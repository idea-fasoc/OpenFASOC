* NGSPICE file created from diff_pair_sample_0225.ext - technology: sky130A

.subckt diff_pair_sample_0225 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t15 w_n2638_n4128# sky130_fd_pr__pfet_01v8 ad=2.607 pd=16.13 as=2.607 ps=16.13 w=15.8 l=1.06
X1 VTAIL.t18 VP.t1 VDD1.t8 w_n2638_n4128# sky130_fd_pr__pfet_01v8 ad=2.607 pd=16.13 as=2.607 ps=16.13 w=15.8 l=1.06
X2 VTAIL.t7 VN.t0 VDD2.t9 w_n2638_n4128# sky130_fd_pr__pfet_01v8 ad=2.607 pd=16.13 as=2.607 ps=16.13 w=15.8 l=1.06
X3 B.t11 B.t9 B.t10 w_n2638_n4128# sky130_fd_pr__pfet_01v8 ad=6.162 pd=32.38 as=0 ps=0 w=15.8 l=1.06
X4 B.t8 B.t6 B.t7 w_n2638_n4128# sky130_fd_pr__pfet_01v8 ad=6.162 pd=32.38 as=0 ps=0 w=15.8 l=1.06
X5 VTAIL.t12 VP.t2 VDD1.t7 w_n2638_n4128# sky130_fd_pr__pfet_01v8 ad=2.607 pd=16.13 as=2.607 ps=16.13 w=15.8 l=1.06
X6 VTAIL.t17 VP.t3 VDD1.t6 w_n2638_n4128# sky130_fd_pr__pfet_01v8 ad=2.607 pd=16.13 as=2.607 ps=16.13 w=15.8 l=1.06
X7 VDD2.t8 VN.t1 VTAIL.t6 w_n2638_n4128# sky130_fd_pr__pfet_01v8 ad=6.162 pd=32.38 as=2.607 ps=16.13 w=15.8 l=1.06
X8 B.t5 B.t3 B.t4 w_n2638_n4128# sky130_fd_pr__pfet_01v8 ad=6.162 pd=32.38 as=0 ps=0 w=15.8 l=1.06
X9 VDD1.t5 VP.t4 VTAIL.t19 w_n2638_n4128# sky130_fd_pr__pfet_01v8 ad=2.607 pd=16.13 as=2.607 ps=16.13 w=15.8 l=1.06
X10 VDD2.t7 VN.t2 VTAIL.t9 w_n2638_n4128# sky130_fd_pr__pfet_01v8 ad=2.607 pd=16.13 as=6.162 ps=32.38 w=15.8 l=1.06
X11 VDD1.t4 VP.t5 VTAIL.t13 w_n2638_n4128# sky130_fd_pr__pfet_01v8 ad=6.162 pd=32.38 as=2.607 ps=16.13 w=15.8 l=1.06
X12 VDD1.t3 VP.t6 VTAIL.t11 w_n2638_n4128# sky130_fd_pr__pfet_01v8 ad=2.607 pd=16.13 as=6.162 ps=32.38 w=15.8 l=1.06
X13 VDD1.t2 VP.t7 VTAIL.t16 w_n2638_n4128# sky130_fd_pr__pfet_01v8 ad=2.607 pd=16.13 as=6.162 ps=32.38 w=15.8 l=1.06
X14 VTAIL.t1 VN.t3 VDD2.t6 w_n2638_n4128# sky130_fd_pr__pfet_01v8 ad=2.607 pd=16.13 as=2.607 ps=16.13 w=15.8 l=1.06
X15 VDD2.t5 VN.t4 VTAIL.t3 w_n2638_n4128# sky130_fd_pr__pfet_01v8 ad=2.607 pd=16.13 as=2.607 ps=16.13 w=15.8 l=1.06
X16 B.t2 B.t0 B.t1 w_n2638_n4128# sky130_fd_pr__pfet_01v8 ad=6.162 pd=32.38 as=0 ps=0 w=15.8 l=1.06
X17 VTAIL.t0 VN.t5 VDD2.t4 w_n2638_n4128# sky130_fd_pr__pfet_01v8 ad=2.607 pd=16.13 as=2.607 ps=16.13 w=15.8 l=1.06
X18 VDD2.t3 VN.t6 VTAIL.t2 w_n2638_n4128# sky130_fd_pr__pfet_01v8 ad=2.607 pd=16.13 as=2.607 ps=16.13 w=15.8 l=1.06
X19 VDD2.t2 VN.t7 VTAIL.t4 w_n2638_n4128# sky130_fd_pr__pfet_01v8 ad=6.162 pd=32.38 as=2.607 ps=16.13 w=15.8 l=1.06
X20 VDD1.t1 VP.t8 VTAIL.t14 w_n2638_n4128# sky130_fd_pr__pfet_01v8 ad=6.162 pd=32.38 as=2.607 ps=16.13 w=15.8 l=1.06
X21 VTAIL.t10 VP.t9 VDD1.t0 w_n2638_n4128# sky130_fd_pr__pfet_01v8 ad=2.607 pd=16.13 as=2.607 ps=16.13 w=15.8 l=1.06
X22 VDD2.t1 VN.t8 VTAIL.t5 w_n2638_n4128# sky130_fd_pr__pfet_01v8 ad=2.607 pd=16.13 as=6.162 ps=32.38 w=15.8 l=1.06
X23 VTAIL.t8 VN.t9 VDD2.t0 w_n2638_n4128# sky130_fd_pr__pfet_01v8 ad=2.607 pd=16.13 as=2.607 ps=16.13 w=15.8 l=1.06
R0 VP.n10 VP.t8 416.486
R1 VP.n5 VP.t5 396.286
R2 VP.n41 VP.t6 396.286
R3 VP.n23 VP.t7 396.286
R4 VP.n34 VP.t0 359.226
R5 VP.n29 VP.t9 359.226
R6 VP.n1 VP.t3 359.226
R7 VP.n16 VP.t4 359.226
R8 VP.n7 VP.t2 359.226
R9 VP.n11 VP.t1 359.226
R10 VP.n13 VP.n12 161.3
R11 VP.n14 VP.n9 161.3
R12 VP.n16 VP.n15 161.3
R13 VP.n17 VP.n8 161.3
R14 VP.n19 VP.n18 161.3
R15 VP.n21 VP.n20 161.3
R16 VP.n22 VP.n6 161.3
R17 VP.n40 VP.n0 161.3
R18 VP.n39 VP.n38 161.3
R19 VP.n37 VP.n36 161.3
R20 VP.n35 VP.n2 161.3
R21 VP.n34 VP.n33 161.3
R22 VP.n32 VP.n3 161.3
R23 VP.n31 VP.n30 161.3
R24 VP.n28 VP.n4 161.3
R25 VP.n27 VP.n26 161.3
R26 VP.n24 VP.n23 80.6037
R27 VP.n42 VP.n41 80.6037
R28 VP.n25 VP.n5 80.6037
R29 VP.n30 VP.n3 56.5617
R30 VP.n36 VP.n35 56.5617
R31 VP.n18 VP.n17 56.5617
R32 VP.n12 VP.n9 56.5617
R33 VP.n25 VP.n24 47.687
R34 VP.n11 VP.n10 38.3612
R35 VP.n27 VP.n5 36.5157
R36 VP.n41 VP.n40 36.5157
R37 VP.n23 VP.n22 36.5157
R38 VP.n28 VP.n27 32.3425
R39 VP.n40 VP.n39 32.3425
R40 VP.n22 VP.n21 32.3425
R41 VP.n13 VP.n10 29.1526
R42 VP.n34 VP.n3 24.5923
R43 VP.n35 VP.n34 24.5923
R44 VP.n16 VP.n9 24.5923
R45 VP.n17 VP.n16 24.5923
R46 VP.n30 VP.n29 19.1821
R47 VP.n36 VP.n1 19.1821
R48 VP.n18 VP.n7 19.1821
R49 VP.n12 VP.n11 19.1821
R50 VP.n29 VP.n28 5.4107
R51 VP.n39 VP.n1 5.4107
R52 VP.n21 VP.n7 5.4107
R53 VP.n24 VP.n6 0.285035
R54 VP.n26 VP.n25 0.285035
R55 VP.n42 VP.n0 0.285035
R56 VP.n14 VP.n13 0.189894
R57 VP.n15 VP.n14 0.189894
R58 VP.n15 VP.n8 0.189894
R59 VP.n19 VP.n8 0.189894
R60 VP.n20 VP.n19 0.189894
R61 VP.n20 VP.n6 0.189894
R62 VP.n26 VP.n4 0.189894
R63 VP.n31 VP.n4 0.189894
R64 VP.n32 VP.n31 0.189894
R65 VP.n33 VP.n32 0.189894
R66 VP.n33 VP.n2 0.189894
R67 VP.n37 VP.n2 0.189894
R68 VP.n38 VP.n37 0.189894
R69 VP.n38 VP.n0 0.189894
R70 VP VP.n42 0.146778
R71 VTAIL.n11 VTAIL.t9 56.9537
R72 VTAIL.n16 VTAIL.t16 56.9536
R73 VTAIL.n17 VTAIL.t5 56.9536
R74 VTAIL.n2 VTAIL.t11 56.9536
R75 VTAIL.n15 VTAIL.n14 54.8965
R76 VTAIL.n13 VTAIL.n12 54.8965
R77 VTAIL.n10 VTAIL.n9 54.8965
R78 VTAIL.n8 VTAIL.n7 54.8965
R79 VTAIL.n19 VTAIL.n18 54.8962
R80 VTAIL.n1 VTAIL.n0 54.8962
R81 VTAIL.n4 VTAIL.n3 54.8962
R82 VTAIL.n6 VTAIL.n5 54.8962
R83 VTAIL.n8 VTAIL.n6 28.3841
R84 VTAIL.n17 VTAIL.n16 27.1858
R85 VTAIL.n18 VTAIL.t3 2.05778
R86 VTAIL.n18 VTAIL.t7 2.05778
R87 VTAIL.n0 VTAIL.t4 2.05778
R88 VTAIL.n0 VTAIL.t1 2.05778
R89 VTAIL.n3 VTAIL.t15 2.05778
R90 VTAIL.n3 VTAIL.t17 2.05778
R91 VTAIL.n5 VTAIL.t13 2.05778
R92 VTAIL.n5 VTAIL.t10 2.05778
R93 VTAIL.n14 VTAIL.t19 2.05778
R94 VTAIL.n14 VTAIL.t12 2.05778
R95 VTAIL.n12 VTAIL.t14 2.05778
R96 VTAIL.n12 VTAIL.t18 2.05778
R97 VTAIL.n9 VTAIL.t2 2.05778
R98 VTAIL.n9 VTAIL.t0 2.05778
R99 VTAIL.n7 VTAIL.t6 2.05778
R100 VTAIL.n7 VTAIL.t8 2.05778
R101 VTAIL.n10 VTAIL.n8 1.19878
R102 VTAIL.n11 VTAIL.n10 1.19878
R103 VTAIL.n15 VTAIL.n13 1.19878
R104 VTAIL.n16 VTAIL.n15 1.19878
R105 VTAIL.n6 VTAIL.n4 1.19878
R106 VTAIL.n4 VTAIL.n2 1.19878
R107 VTAIL.n19 VTAIL.n17 1.19878
R108 VTAIL.n13 VTAIL.n11 1.06947
R109 VTAIL.n2 VTAIL.n1 1.06947
R110 VTAIL VTAIL.n1 0.957397
R111 VTAIL VTAIL.n19 0.241879
R112 VDD1.n1 VDD1.t1 74.8308
R113 VDD1.n3 VDD1.t4 74.8307
R114 VDD1.n5 VDD1.n4 72.4184
R115 VDD1.n1 VDD1.n0 71.5753
R116 VDD1.n7 VDD1.n6 71.5751
R117 VDD1.n3 VDD1.n2 71.575
R118 VDD1.n7 VDD1.n5 44.2099
R119 VDD1.n6 VDD1.t7 2.05778
R120 VDD1.n6 VDD1.t2 2.05778
R121 VDD1.n0 VDD1.t8 2.05778
R122 VDD1.n0 VDD1.t5 2.05778
R123 VDD1.n4 VDD1.t6 2.05778
R124 VDD1.n4 VDD1.t3 2.05778
R125 VDD1.n2 VDD1.t0 2.05778
R126 VDD1.n2 VDD1.t9 2.05778
R127 VDD1 VDD1.n7 0.841017
R128 VDD1 VDD1.n1 0.358259
R129 VDD1.n5 VDD1.n3 0.244723
R130 VN.n4 VN.t7 416.486
R131 VN.n23 VN.t2 416.486
R132 VN.n17 VN.t8 396.286
R133 VN.n36 VN.t1 396.286
R134 VN.n10 VN.t4 359.226
R135 VN.n5 VN.t3 359.226
R136 VN.n1 VN.t0 359.226
R137 VN.n29 VN.t6 359.226
R138 VN.n24 VN.t5 359.226
R139 VN.n20 VN.t9 359.226
R140 VN.n35 VN.n19 161.3
R141 VN.n34 VN.n33 161.3
R142 VN.n32 VN.n31 161.3
R143 VN.n30 VN.n21 161.3
R144 VN.n29 VN.n28 161.3
R145 VN.n27 VN.n22 161.3
R146 VN.n26 VN.n25 161.3
R147 VN.n16 VN.n0 161.3
R148 VN.n15 VN.n14 161.3
R149 VN.n13 VN.n12 161.3
R150 VN.n11 VN.n2 161.3
R151 VN.n10 VN.n9 161.3
R152 VN.n8 VN.n3 161.3
R153 VN.n7 VN.n6 161.3
R154 VN.n37 VN.n36 80.6037
R155 VN.n18 VN.n17 80.6037
R156 VN.n6 VN.n3 56.5617
R157 VN.n12 VN.n11 56.5617
R158 VN.n25 VN.n22 56.5617
R159 VN.n31 VN.n30 56.5617
R160 VN VN.n37 47.9725
R161 VN.n5 VN.n4 38.3612
R162 VN.n24 VN.n23 38.3612
R163 VN.n17 VN.n16 36.5157
R164 VN.n36 VN.n35 36.5157
R165 VN.n16 VN.n15 32.3425
R166 VN.n35 VN.n34 32.3425
R167 VN.n26 VN.n23 29.1526
R168 VN.n7 VN.n4 29.1526
R169 VN.n10 VN.n3 24.5923
R170 VN.n11 VN.n10 24.5923
R171 VN.n30 VN.n29 24.5923
R172 VN.n29 VN.n22 24.5923
R173 VN.n6 VN.n5 19.1821
R174 VN.n12 VN.n1 19.1821
R175 VN.n25 VN.n24 19.1821
R176 VN.n31 VN.n20 19.1821
R177 VN.n15 VN.n1 5.4107
R178 VN.n34 VN.n20 5.4107
R179 VN.n37 VN.n19 0.285035
R180 VN.n18 VN.n0 0.285035
R181 VN.n33 VN.n19 0.189894
R182 VN.n33 VN.n32 0.189894
R183 VN.n32 VN.n21 0.189894
R184 VN.n28 VN.n21 0.189894
R185 VN.n28 VN.n27 0.189894
R186 VN.n27 VN.n26 0.189894
R187 VN.n8 VN.n7 0.189894
R188 VN.n9 VN.n8 0.189894
R189 VN.n9 VN.n2 0.189894
R190 VN.n13 VN.n2 0.189894
R191 VN.n14 VN.n13 0.189894
R192 VN.n14 VN.n0 0.189894
R193 VN VN.n18 0.146778
R194 VDD2.n1 VDD2.t2 74.8307
R195 VDD2.n4 VDD2.t8 73.6325
R196 VDD2.n3 VDD2.n2 72.4184
R197 VDD2 VDD2.n7 72.4156
R198 VDD2.n6 VDD2.n5 71.5753
R199 VDD2.n1 VDD2.n0 71.575
R200 VDD2.n4 VDD2.n3 43.0278
R201 VDD2.n7 VDD2.t4 2.05778
R202 VDD2.n7 VDD2.t7 2.05778
R203 VDD2.n5 VDD2.t0 2.05778
R204 VDD2.n5 VDD2.t3 2.05778
R205 VDD2.n2 VDD2.t9 2.05778
R206 VDD2.n2 VDD2.t1 2.05778
R207 VDD2.n0 VDD2.t6 2.05778
R208 VDD2.n0 VDD2.t5 2.05778
R209 VDD2.n6 VDD2.n4 1.19878
R210 VDD2 VDD2.n6 0.358259
R211 VDD2.n3 VDD2.n1 0.244723
R212 B.n411 B.n410 585
R213 B.n409 B.n114 585
R214 B.n408 B.n407 585
R215 B.n406 B.n115 585
R216 B.n405 B.n404 585
R217 B.n403 B.n116 585
R218 B.n402 B.n401 585
R219 B.n400 B.n117 585
R220 B.n399 B.n398 585
R221 B.n397 B.n118 585
R222 B.n396 B.n395 585
R223 B.n394 B.n119 585
R224 B.n393 B.n392 585
R225 B.n391 B.n120 585
R226 B.n390 B.n389 585
R227 B.n388 B.n121 585
R228 B.n387 B.n386 585
R229 B.n385 B.n122 585
R230 B.n384 B.n383 585
R231 B.n382 B.n123 585
R232 B.n381 B.n380 585
R233 B.n379 B.n124 585
R234 B.n378 B.n377 585
R235 B.n376 B.n125 585
R236 B.n375 B.n374 585
R237 B.n373 B.n126 585
R238 B.n372 B.n371 585
R239 B.n370 B.n127 585
R240 B.n369 B.n368 585
R241 B.n367 B.n128 585
R242 B.n366 B.n365 585
R243 B.n364 B.n129 585
R244 B.n363 B.n362 585
R245 B.n361 B.n130 585
R246 B.n360 B.n359 585
R247 B.n358 B.n131 585
R248 B.n357 B.n356 585
R249 B.n355 B.n132 585
R250 B.n354 B.n353 585
R251 B.n352 B.n133 585
R252 B.n351 B.n350 585
R253 B.n349 B.n134 585
R254 B.n348 B.n347 585
R255 B.n346 B.n135 585
R256 B.n345 B.n344 585
R257 B.n343 B.n136 585
R258 B.n342 B.n341 585
R259 B.n340 B.n137 585
R260 B.n339 B.n338 585
R261 B.n337 B.n138 585
R262 B.n336 B.n335 585
R263 B.n334 B.n139 585
R264 B.n333 B.n332 585
R265 B.n330 B.n140 585
R266 B.n329 B.n328 585
R267 B.n327 B.n143 585
R268 B.n326 B.n325 585
R269 B.n324 B.n144 585
R270 B.n323 B.n322 585
R271 B.n321 B.n145 585
R272 B.n320 B.n319 585
R273 B.n318 B.n146 585
R274 B.n316 B.n315 585
R275 B.n314 B.n149 585
R276 B.n313 B.n312 585
R277 B.n311 B.n150 585
R278 B.n310 B.n309 585
R279 B.n308 B.n151 585
R280 B.n307 B.n306 585
R281 B.n305 B.n152 585
R282 B.n304 B.n303 585
R283 B.n302 B.n153 585
R284 B.n301 B.n300 585
R285 B.n299 B.n154 585
R286 B.n298 B.n297 585
R287 B.n296 B.n155 585
R288 B.n295 B.n294 585
R289 B.n293 B.n156 585
R290 B.n292 B.n291 585
R291 B.n290 B.n157 585
R292 B.n289 B.n288 585
R293 B.n287 B.n158 585
R294 B.n286 B.n285 585
R295 B.n284 B.n159 585
R296 B.n283 B.n282 585
R297 B.n281 B.n160 585
R298 B.n280 B.n279 585
R299 B.n278 B.n161 585
R300 B.n277 B.n276 585
R301 B.n275 B.n162 585
R302 B.n274 B.n273 585
R303 B.n272 B.n163 585
R304 B.n271 B.n270 585
R305 B.n269 B.n164 585
R306 B.n268 B.n267 585
R307 B.n266 B.n165 585
R308 B.n265 B.n264 585
R309 B.n263 B.n166 585
R310 B.n262 B.n261 585
R311 B.n260 B.n167 585
R312 B.n259 B.n258 585
R313 B.n257 B.n168 585
R314 B.n256 B.n255 585
R315 B.n254 B.n169 585
R316 B.n253 B.n252 585
R317 B.n251 B.n170 585
R318 B.n250 B.n249 585
R319 B.n248 B.n171 585
R320 B.n247 B.n246 585
R321 B.n245 B.n172 585
R322 B.n244 B.n243 585
R323 B.n242 B.n173 585
R324 B.n241 B.n240 585
R325 B.n239 B.n174 585
R326 B.n238 B.n237 585
R327 B.n412 B.n113 585
R328 B.n414 B.n413 585
R329 B.n415 B.n112 585
R330 B.n417 B.n416 585
R331 B.n418 B.n111 585
R332 B.n420 B.n419 585
R333 B.n421 B.n110 585
R334 B.n423 B.n422 585
R335 B.n424 B.n109 585
R336 B.n426 B.n425 585
R337 B.n427 B.n108 585
R338 B.n429 B.n428 585
R339 B.n430 B.n107 585
R340 B.n432 B.n431 585
R341 B.n433 B.n106 585
R342 B.n435 B.n434 585
R343 B.n436 B.n105 585
R344 B.n438 B.n437 585
R345 B.n439 B.n104 585
R346 B.n441 B.n440 585
R347 B.n442 B.n103 585
R348 B.n444 B.n443 585
R349 B.n445 B.n102 585
R350 B.n447 B.n446 585
R351 B.n448 B.n101 585
R352 B.n450 B.n449 585
R353 B.n451 B.n100 585
R354 B.n453 B.n452 585
R355 B.n454 B.n99 585
R356 B.n456 B.n455 585
R357 B.n457 B.n98 585
R358 B.n459 B.n458 585
R359 B.n460 B.n97 585
R360 B.n462 B.n461 585
R361 B.n463 B.n96 585
R362 B.n465 B.n464 585
R363 B.n466 B.n95 585
R364 B.n468 B.n467 585
R365 B.n469 B.n94 585
R366 B.n471 B.n470 585
R367 B.n472 B.n93 585
R368 B.n474 B.n473 585
R369 B.n475 B.n92 585
R370 B.n477 B.n476 585
R371 B.n478 B.n91 585
R372 B.n480 B.n479 585
R373 B.n481 B.n90 585
R374 B.n483 B.n482 585
R375 B.n484 B.n89 585
R376 B.n486 B.n485 585
R377 B.n487 B.n88 585
R378 B.n489 B.n488 585
R379 B.n490 B.n87 585
R380 B.n492 B.n491 585
R381 B.n493 B.n86 585
R382 B.n495 B.n494 585
R383 B.n496 B.n85 585
R384 B.n498 B.n497 585
R385 B.n499 B.n84 585
R386 B.n501 B.n500 585
R387 B.n502 B.n83 585
R388 B.n504 B.n503 585
R389 B.n505 B.n82 585
R390 B.n507 B.n506 585
R391 B.n508 B.n81 585
R392 B.n510 B.n509 585
R393 B.n683 B.n18 585
R394 B.n682 B.n681 585
R395 B.n680 B.n19 585
R396 B.n679 B.n678 585
R397 B.n677 B.n20 585
R398 B.n676 B.n675 585
R399 B.n674 B.n21 585
R400 B.n673 B.n672 585
R401 B.n671 B.n22 585
R402 B.n670 B.n669 585
R403 B.n668 B.n23 585
R404 B.n667 B.n666 585
R405 B.n665 B.n24 585
R406 B.n664 B.n663 585
R407 B.n662 B.n25 585
R408 B.n661 B.n660 585
R409 B.n659 B.n26 585
R410 B.n658 B.n657 585
R411 B.n656 B.n27 585
R412 B.n655 B.n654 585
R413 B.n653 B.n28 585
R414 B.n652 B.n651 585
R415 B.n650 B.n29 585
R416 B.n649 B.n648 585
R417 B.n647 B.n30 585
R418 B.n646 B.n645 585
R419 B.n644 B.n31 585
R420 B.n643 B.n642 585
R421 B.n641 B.n32 585
R422 B.n640 B.n639 585
R423 B.n638 B.n33 585
R424 B.n637 B.n636 585
R425 B.n635 B.n34 585
R426 B.n634 B.n633 585
R427 B.n632 B.n35 585
R428 B.n631 B.n630 585
R429 B.n629 B.n36 585
R430 B.n628 B.n627 585
R431 B.n626 B.n37 585
R432 B.n625 B.n624 585
R433 B.n623 B.n38 585
R434 B.n622 B.n621 585
R435 B.n620 B.n39 585
R436 B.n619 B.n618 585
R437 B.n617 B.n40 585
R438 B.n616 B.n615 585
R439 B.n614 B.n41 585
R440 B.n613 B.n612 585
R441 B.n611 B.n42 585
R442 B.n610 B.n609 585
R443 B.n608 B.n43 585
R444 B.n607 B.n606 585
R445 B.n605 B.n44 585
R446 B.n604 B.n603 585
R447 B.n602 B.n45 585
R448 B.n601 B.n600 585
R449 B.n599 B.n49 585
R450 B.n598 B.n597 585
R451 B.n596 B.n50 585
R452 B.n595 B.n594 585
R453 B.n593 B.n51 585
R454 B.n592 B.n591 585
R455 B.n589 B.n52 585
R456 B.n588 B.n587 585
R457 B.n586 B.n55 585
R458 B.n585 B.n584 585
R459 B.n583 B.n56 585
R460 B.n582 B.n581 585
R461 B.n580 B.n57 585
R462 B.n579 B.n578 585
R463 B.n577 B.n58 585
R464 B.n576 B.n575 585
R465 B.n574 B.n59 585
R466 B.n573 B.n572 585
R467 B.n571 B.n60 585
R468 B.n570 B.n569 585
R469 B.n568 B.n61 585
R470 B.n567 B.n566 585
R471 B.n565 B.n62 585
R472 B.n564 B.n563 585
R473 B.n562 B.n63 585
R474 B.n561 B.n560 585
R475 B.n559 B.n64 585
R476 B.n558 B.n557 585
R477 B.n556 B.n65 585
R478 B.n555 B.n554 585
R479 B.n553 B.n66 585
R480 B.n552 B.n551 585
R481 B.n550 B.n67 585
R482 B.n549 B.n548 585
R483 B.n547 B.n68 585
R484 B.n546 B.n545 585
R485 B.n544 B.n69 585
R486 B.n543 B.n542 585
R487 B.n541 B.n70 585
R488 B.n540 B.n539 585
R489 B.n538 B.n71 585
R490 B.n537 B.n536 585
R491 B.n535 B.n72 585
R492 B.n534 B.n533 585
R493 B.n532 B.n73 585
R494 B.n531 B.n530 585
R495 B.n529 B.n74 585
R496 B.n528 B.n527 585
R497 B.n526 B.n75 585
R498 B.n525 B.n524 585
R499 B.n523 B.n76 585
R500 B.n522 B.n521 585
R501 B.n520 B.n77 585
R502 B.n519 B.n518 585
R503 B.n517 B.n78 585
R504 B.n516 B.n515 585
R505 B.n514 B.n79 585
R506 B.n513 B.n512 585
R507 B.n511 B.n80 585
R508 B.n685 B.n684 585
R509 B.n686 B.n17 585
R510 B.n688 B.n687 585
R511 B.n689 B.n16 585
R512 B.n691 B.n690 585
R513 B.n692 B.n15 585
R514 B.n694 B.n693 585
R515 B.n695 B.n14 585
R516 B.n697 B.n696 585
R517 B.n698 B.n13 585
R518 B.n700 B.n699 585
R519 B.n701 B.n12 585
R520 B.n703 B.n702 585
R521 B.n704 B.n11 585
R522 B.n706 B.n705 585
R523 B.n707 B.n10 585
R524 B.n709 B.n708 585
R525 B.n710 B.n9 585
R526 B.n712 B.n711 585
R527 B.n713 B.n8 585
R528 B.n715 B.n714 585
R529 B.n716 B.n7 585
R530 B.n718 B.n717 585
R531 B.n719 B.n6 585
R532 B.n721 B.n720 585
R533 B.n722 B.n5 585
R534 B.n724 B.n723 585
R535 B.n725 B.n4 585
R536 B.n727 B.n726 585
R537 B.n728 B.n3 585
R538 B.n730 B.n729 585
R539 B.n731 B.n0 585
R540 B.n2 B.n1 585
R541 B.n191 B.n190 585
R542 B.n193 B.n192 585
R543 B.n194 B.n189 585
R544 B.n196 B.n195 585
R545 B.n197 B.n188 585
R546 B.n199 B.n198 585
R547 B.n200 B.n187 585
R548 B.n202 B.n201 585
R549 B.n203 B.n186 585
R550 B.n205 B.n204 585
R551 B.n206 B.n185 585
R552 B.n208 B.n207 585
R553 B.n209 B.n184 585
R554 B.n211 B.n210 585
R555 B.n212 B.n183 585
R556 B.n214 B.n213 585
R557 B.n215 B.n182 585
R558 B.n217 B.n216 585
R559 B.n218 B.n181 585
R560 B.n220 B.n219 585
R561 B.n221 B.n180 585
R562 B.n223 B.n222 585
R563 B.n224 B.n179 585
R564 B.n226 B.n225 585
R565 B.n227 B.n178 585
R566 B.n229 B.n228 585
R567 B.n230 B.n177 585
R568 B.n232 B.n231 585
R569 B.n233 B.n176 585
R570 B.n235 B.n234 585
R571 B.n236 B.n175 585
R572 B.n147 B.t3 562.543
R573 B.n141 B.t0 562.543
R574 B.n53 B.t6 562.543
R575 B.n46 B.t9 562.543
R576 B.n237 B.n236 535.745
R577 B.n412 B.n411 535.745
R578 B.n509 B.n80 535.745
R579 B.n684 B.n683 535.745
R580 B.n733 B.n732 256.663
R581 B.n732 B.n731 235.042
R582 B.n732 B.n2 235.042
R583 B.n237 B.n174 163.367
R584 B.n241 B.n174 163.367
R585 B.n242 B.n241 163.367
R586 B.n243 B.n242 163.367
R587 B.n243 B.n172 163.367
R588 B.n247 B.n172 163.367
R589 B.n248 B.n247 163.367
R590 B.n249 B.n248 163.367
R591 B.n249 B.n170 163.367
R592 B.n253 B.n170 163.367
R593 B.n254 B.n253 163.367
R594 B.n255 B.n254 163.367
R595 B.n255 B.n168 163.367
R596 B.n259 B.n168 163.367
R597 B.n260 B.n259 163.367
R598 B.n261 B.n260 163.367
R599 B.n261 B.n166 163.367
R600 B.n265 B.n166 163.367
R601 B.n266 B.n265 163.367
R602 B.n267 B.n266 163.367
R603 B.n267 B.n164 163.367
R604 B.n271 B.n164 163.367
R605 B.n272 B.n271 163.367
R606 B.n273 B.n272 163.367
R607 B.n273 B.n162 163.367
R608 B.n277 B.n162 163.367
R609 B.n278 B.n277 163.367
R610 B.n279 B.n278 163.367
R611 B.n279 B.n160 163.367
R612 B.n283 B.n160 163.367
R613 B.n284 B.n283 163.367
R614 B.n285 B.n284 163.367
R615 B.n285 B.n158 163.367
R616 B.n289 B.n158 163.367
R617 B.n290 B.n289 163.367
R618 B.n291 B.n290 163.367
R619 B.n291 B.n156 163.367
R620 B.n295 B.n156 163.367
R621 B.n296 B.n295 163.367
R622 B.n297 B.n296 163.367
R623 B.n297 B.n154 163.367
R624 B.n301 B.n154 163.367
R625 B.n302 B.n301 163.367
R626 B.n303 B.n302 163.367
R627 B.n303 B.n152 163.367
R628 B.n307 B.n152 163.367
R629 B.n308 B.n307 163.367
R630 B.n309 B.n308 163.367
R631 B.n309 B.n150 163.367
R632 B.n313 B.n150 163.367
R633 B.n314 B.n313 163.367
R634 B.n315 B.n314 163.367
R635 B.n315 B.n146 163.367
R636 B.n320 B.n146 163.367
R637 B.n321 B.n320 163.367
R638 B.n322 B.n321 163.367
R639 B.n322 B.n144 163.367
R640 B.n326 B.n144 163.367
R641 B.n327 B.n326 163.367
R642 B.n328 B.n327 163.367
R643 B.n328 B.n140 163.367
R644 B.n333 B.n140 163.367
R645 B.n334 B.n333 163.367
R646 B.n335 B.n334 163.367
R647 B.n335 B.n138 163.367
R648 B.n339 B.n138 163.367
R649 B.n340 B.n339 163.367
R650 B.n341 B.n340 163.367
R651 B.n341 B.n136 163.367
R652 B.n345 B.n136 163.367
R653 B.n346 B.n345 163.367
R654 B.n347 B.n346 163.367
R655 B.n347 B.n134 163.367
R656 B.n351 B.n134 163.367
R657 B.n352 B.n351 163.367
R658 B.n353 B.n352 163.367
R659 B.n353 B.n132 163.367
R660 B.n357 B.n132 163.367
R661 B.n358 B.n357 163.367
R662 B.n359 B.n358 163.367
R663 B.n359 B.n130 163.367
R664 B.n363 B.n130 163.367
R665 B.n364 B.n363 163.367
R666 B.n365 B.n364 163.367
R667 B.n365 B.n128 163.367
R668 B.n369 B.n128 163.367
R669 B.n370 B.n369 163.367
R670 B.n371 B.n370 163.367
R671 B.n371 B.n126 163.367
R672 B.n375 B.n126 163.367
R673 B.n376 B.n375 163.367
R674 B.n377 B.n376 163.367
R675 B.n377 B.n124 163.367
R676 B.n381 B.n124 163.367
R677 B.n382 B.n381 163.367
R678 B.n383 B.n382 163.367
R679 B.n383 B.n122 163.367
R680 B.n387 B.n122 163.367
R681 B.n388 B.n387 163.367
R682 B.n389 B.n388 163.367
R683 B.n389 B.n120 163.367
R684 B.n393 B.n120 163.367
R685 B.n394 B.n393 163.367
R686 B.n395 B.n394 163.367
R687 B.n395 B.n118 163.367
R688 B.n399 B.n118 163.367
R689 B.n400 B.n399 163.367
R690 B.n401 B.n400 163.367
R691 B.n401 B.n116 163.367
R692 B.n405 B.n116 163.367
R693 B.n406 B.n405 163.367
R694 B.n407 B.n406 163.367
R695 B.n407 B.n114 163.367
R696 B.n411 B.n114 163.367
R697 B.n509 B.n508 163.367
R698 B.n508 B.n507 163.367
R699 B.n507 B.n82 163.367
R700 B.n503 B.n82 163.367
R701 B.n503 B.n502 163.367
R702 B.n502 B.n501 163.367
R703 B.n501 B.n84 163.367
R704 B.n497 B.n84 163.367
R705 B.n497 B.n496 163.367
R706 B.n496 B.n495 163.367
R707 B.n495 B.n86 163.367
R708 B.n491 B.n86 163.367
R709 B.n491 B.n490 163.367
R710 B.n490 B.n489 163.367
R711 B.n489 B.n88 163.367
R712 B.n485 B.n88 163.367
R713 B.n485 B.n484 163.367
R714 B.n484 B.n483 163.367
R715 B.n483 B.n90 163.367
R716 B.n479 B.n90 163.367
R717 B.n479 B.n478 163.367
R718 B.n478 B.n477 163.367
R719 B.n477 B.n92 163.367
R720 B.n473 B.n92 163.367
R721 B.n473 B.n472 163.367
R722 B.n472 B.n471 163.367
R723 B.n471 B.n94 163.367
R724 B.n467 B.n94 163.367
R725 B.n467 B.n466 163.367
R726 B.n466 B.n465 163.367
R727 B.n465 B.n96 163.367
R728 B.n461 B.n96 163.367
R729 B.n461 B.n460 163.367
R730 B.n460 B.n459 163.367
R731 B.n459 B.n98 163.367
R732 B.n455 B.n98 163.367
R733 B.n455 B.n454 163.367
R734 B.n454 B.n453 163.367
R735 B.n453 B.n100 163.367
R736 B.n449 B.n100 163.367
R737 B.n449 B.n448 163.367
R738 B.n448 B.n447 163.367
R739 B.n447 B.n102 163.367
R740 B.n443 B.n102 163.367
R741 B.n443 B.n442 163.367
R742 B.n442 B.n441 163.367
R743 B.n441 B.n104 163.367
R744 B.n437 B.n104 163.367
R745 B.n437 B.n436 163.367
R746 B.n436 B.n435 163.367
R747 B.n435 B.n106 163.367
R748 B.n431 B.n106 163.367
R749 B.n431 B.n430 163.367
R750 B.n430 B.n429 163.367
R751 B.n429 B.n108 163.367
R752 B.n425 B.n108 163.367
R753 B.n425 B.n424 163.367
R754 B.n424 B.n423 163.367
R755 B.n423 B.n110 163.367
R756 B.n419 B.n110 163.367
R757 B.n419 B.n418 163.367
R758 B.n418 B.n417 163.367
R759 B.n417 B.n112 163.367
R760 B.n413 B.n112 163.367
R761 B.n413 B.n412 163.367
R762 B.n683 B.n682 163.367
R763 B.n682 B.n19 163.367
R764 B.n678 B.n19 163.367
R765 B.n678 B.n677 163.367
R766 B.n677 B.n676 163.367
R767 B.n676 B.n21 163.367
R768 B.n672 B.n21 163.367
R769 B.n672 B.n671 163.367
R770 B.n671 B.n670 163.367
R771 B.n670 B.n23 163.367
R772 B.n666 B.n23 163.367
R773 B.n666 B.n665 163.367
R774 B.n665 B.n664 163.367
R775 B.n664 B.n25 163.367
R776 B.n660 B.n25 163.367
R777 B.n660 B.n659 163.367
R778 B.n659 B.n658 163.367
R779 B.n658 B.n27 163.367
R780 B.n654 B.n27 163.367
R781 B.n654 B.n653 163.367
R782 B.n653 B.n652 163.367
R783 B.n652 B.n29 163.367
R784 B.n648 B.n29 163.367
R785 B.n648 B.n647 163.367
R786 B.n647 B.n646 163.367
R787 B.n646 B.n31 163.367
R788 B.n642 B.n31 163.367
R789 B.n642 B.n641 163.367
R790 B.n641 B.n640 163.367
R791 B.n640 B.n33 163.367
R792 B.n636 B.n33 163.367
R793 B.n636 B.n635 163.367
R794 B.n635 B.n634 163.367
R795 B.n634 B.n35 163.367
R796 B.n630 B.n35 163.367
R797 B.n630 B.n629 163.367
R798 B.n629 B.n628 163.367
R799 B.n628 B.n37 163.367
R800 B.n624 B.n37 163.367
R801 B.n624 B.n623 163.367
R802 B.n623 B.n622 163.367
R803 B.n622 B.n39 163.367
R804 B.n618 B.n39 163.367
R805 B.n618 B.n617 163.367
R806 B.n617 B.n616 163.367
R807 B.n616 B.n41 163.367
R808 B.n612 B.n41 163.367
R809 B.n612 B.n611 163.367
R810 B.n611 B.n610 163.367
R811 B.n610 B.n43 163.367
R812 B.n606 B.n43 163.367
R813 B.n606 B.n605 163.367
R814 B.n605 B.n604 163.367
R815 B.n604 B.n45 163.367
R816 B.n600 B.n45 163.367
R817 B.n600 B.n599 163.367
R818 B.n599 B.n598 163.367
R819 B.n598 B.n50 163.367
R820 B.n594 B.n50 163.367
R821 B.n594 B.n593 163.367
R822 B.n593 B.n592 163.367
R823 B.n592 B.n52 163.367
R824 B.n587 B.n52 163.367
R825 B.n587 B.n586 163.367
R826 B.n586 B.n585 163.367
R827 B.n585 B.n56 163.367
R828 B.n581 B.n56 163.367
R829 B.n581 B.n580 163.367
R830 B.n580 B.n579 163.367
R831 B.n579 B.n58 163.367
R832 B.n575 B.n58 163.367
R833 B.n575 B.n574 163.367
R834 B.n574 B.n573 163.367
R835 B.n573 B.n60 163.367
R836 B.n569 B.n60 163.367
R837 B.n569 B.n568 163.367
R838 B.n568 B.n567 163.367
R839 B.n567 B.n62 163.367
R840 B.n563 B.n62 163.367
R841 B.n563 B.n562 163.367
R842 B.n562 B.n561 163.367
R843 B.n561 B.n64 163.367
R844 B.n557 B.n64 163.367
R845 B.n557 B.n556 163.367
R846 B.n556 B.n555 163.367
R847 B.n555 B.n66 163.367
R848 B.n551 B.n66 163.367
R849 B.n551 B.n550 163.367
R850 B.n550 B.n549 163.367
R851 B.n549 B.n68 163.367
R852 B.n545 B.n68 163.367
R853 B.n545 B.n544 163.367
R854 B.n544 B.n543 163.367
R855 B.n543 B.n70 163.367
R856 B.n539 B.n70 163.367
R857 B.n539 B.n538 163.367
R858 B.n538 B.n537 163.367
R859 B.n537 B.n72 163.367
R860 B.n533 B.n72 163.367
R861 B.n533 B.n532 163.367
R862 B.n532 B.n531 163.367
R863 B.n531 B.n74 163.367
R864 B.n527 B.n74 163.367
R865 B.n527 B.n526 163.367
R866 B.n526 B.n525 163.367
R867 B.n525 B.n76 163.367
R868 B.n521 B.n76 163.367
R869 B.n521 B.n520 163.367
R870 B.n520 B.n519 163.367
R871 B.n519 B.n78 163.367
R872 B.n515 B.n78 163.367
R873 B.n515 B.n514 163.367
R874 B.n514 B.n513 163.367
R875 B.n513 B.n80 163.367
R876 B.n684 B.n17 163.367
R877 B.n688 B.n17 163.367
R878 B.n689 B.n688 163.367
R879 B.n690 B.n689 163.367
R880 B.n690 B.n15 163.367
R881 B.n694 B.n15 163.367
R882 B.n695 B.n694 163.367
R883 B.n696 B.n695 163.367
R884 B.n696 B.n13 163.367
R885 B.n700 B.n13 163.367
R886 B.n701 B.n700 163.367
R887 B.n702 B.n701 163.367
R888 B.n702 B.n11 163.367
R889 B.n706 B.n11 163.367
R890 B.n707 B.n706 163.367
R891 B.n708 B.n707 163.367
R892 B.n708 B.n9 163.367
R893 B.n712 B.n9 163.367
R894 B.n713 B.n712 163.367
R895 B.n714 B.n713 163.367
R896 B.n714 B.n7 163.367
R897 B.n718 B.n7 163.367
R898 B.n719 B.n718 163.367
R899 B.n720 B.n719 163.367
R900 B.n720 B.n5 163.367
R901 B.n724 B.n5 163.367
R902 B.n725 B.n724 163.367
R903 B.n726 B.n725 163.367
R904 B.n726 B.n3 163.367
R905 B.n730 B.n3 163.367
R906 B.n731 B.n730 163.367
R907 B.n190 B.n2 163.367
R908 B.n193 B.n190 163.367
R909 B.n194 B.n193 163.367
R910 B.n195 B.n194 163.367
R911 B.n195 B.n188 163.367
R912 B.n199 B.n188 163.367
R913 B.n200 B.n199 163.367
R914 B.n201 B.n200 163.367
R915 B.n201 B.n186 163.367
R916 B.n205 B.n186 163.367
R917 B.n206 B.n205 163.367
R918 B.n207 B.n206 163.367
R919 B.n207 B.n184 163.367
R920 B.n211 B.n184 163.367
R921 B.n212 B.n211 163.367
R922 B.n213 B.n212 163.367
R923 B.n213 B.n182 163.367
R924 B.n217 B.n182 163.367
R925 B.n218 B.n217 163.367
R926 B.n219 B.n218 163.367
R927 B.n219 B.n180 163.367
R928 B.n223 B.n180 163.367
R929 B.n224 B.n223 163.367
R930 B.n225 B.n224 163.367
R931 B.n225 B.n178 163.367
R932 B.n229 B.n178 163.367
R933 B.n230 B.n229 163.367
R934 B.n231 B.n230 163.367
R935 B.n231 B.n176 163.367
R936 B.n235 B.n176 163.367
R937 B.n236 B.n235 163.367
R938 B.n141 B.t1 136.513
R939 B.n53 B.t8 136.513
R940 B.n147 B.t4 136.494
R941 B.n46 B.t11 136.494
R942 B.n142 B.t2 109.555
R943 B.n54 B.t7 109.555
R944 B.n148 B.t5 109.535
R945 B.n47 B.t10 109.535
R946 B.n317 B.n148 59.5399
R947 B.n331 B.n142 59.5399
R948 B.n590 B.n54 59.5399
R949 B.n48 B.n47 59.5399
R950 B.n685 B.n18 34.8103
R951 B.n511 B.n510 34.8103
R952 B.n410 B.n113 34.8103
R953 B.n238 B.n175 34.8103
R954 B.n148 B.n147 26.9581
R955 B.n142 B.n141 26.9581
R956 B.n54 B.n53 26.9581
R957 B.n47 B.n46 26.9581
R958 B B.n733 18.0485
R959 B.n686 B.n685 10.6151
R960 B.n687 B.n686 10.6151
R961 B.n687 B.n16 10.6151
R962 B.n691 B.n16 10.6151
R963 B.n692 B.n691 10.6151
R964 B.n693 B.n692 10.6151
R965 B.n693 B.n14 10.6151
R966 B.n697 B.n14 10.6151
R967 B.n698 B.n697 10.6151
R968 B.n699 B.n698 10.6151
R969 B.n699 B.n12 10.6151
R970 B.n703 B.n12 10.6151
R971 B.n704 B.n703 10.6151
R972 B.n705 B.n704 10.6151
R973 B.n705 B.n10 10.6151
R974 B.n709 B.n10 10.6151
R975 B.n710 B.n709 10.6151
R976 B.n711 B.n710 10.6151
R977 B.n711 B.n8 10.6151
R978 B.n715 B.n8 10.6151
R979 B.n716 B.n715 10.6151
R980 B.n717 B.n716 10.6151
R981 B.n717 B.n6 10.6151
R982 B.n721 B.n6 10.6151
R983 B.n722 B.n721 10.6151
R984 B.n723 B.n722 10.6151
R985 B.n723 B.n4 10.6151
R986 B.n727 B.n4 10.6151
R987 B.n728 B.n727 10.6151
R988 B.n729 B.n728 10.6151
R989 B.n729 B.n0 10.6151
R990 B.n681 B.n18 10.6151
R991 B.n681 B.n680 10.6151
R992 B.n680 B.n679 10.6151
R993 B.n679 B.n20 10.6151
R994 B.n675 B.n20 10.6151
R995 B.n675 B.n674 10.6151
R996 B.n674 B.n673 10.6151
R997 B.n673 B.n22 10.6151
R998 B.n669 B.n22 10.6151
R999 B.n669 B.n668 10.6151
R1000 B.n668 B.n667 10.6151
R1001 B.n667 B.n24 10.6151
R1002 B.n663 B.n24 10.6151
R1003 B.n663 B.n662 10.6151
R1004 B.n662 B.n661 10.6151
R1005 B.n661 B.n26 10.6151
R1006 B.n657 B.n26 10.6151
R1007 B.n657 B.n656 10.6151
R1008 B.n656 B.n655 10.6151
R1009 B.n655 B.n28 10.6151
R1010 B.n651 B.n28 10.6151
R1011 B.n651 B.n650 10.6151
R1012 B.n650 B.n649 10.6151
R1013 B.n649 B.n30 10.6151
R1014 B.n645 B.n30 10.6151
R1015 B.n645 B.n644 10.6151
R1016 B.n644 B.n643 10.6151
R1017 B.n643 B.n32 10.6151
R1018 B.n639 B.n32 10.6151
R1019 B.n639 B.n638 10.6151
R1020 B.n638 B.n637 10.6151
R1021 B.n637 B.n34 10.6151
R1022 B.n633 B.n34 10.6151
R1023 B.n633 B.n632 10.6151
R1024 B.n632 B.n631 10.6151
R1025 B.n631 B.n36 10.6151
R1026 B.n627 B.n36 10.6151
R1027 B.n627 B.n626 10.6151
R1028 B.n626 B.n625 10.6151
R1029 B.n625 B.n38 10.6151
R1030 B.n621 B.n38 10.6151
R1031 B.n621 B.n620 10.6151
R1032 B.n620 B.n619 10.6151
R1033 B.n619 B.n40 10.6151
R1034 B.n615 B.n40 10.6151
R1035 B.n615 B.n614 10.6151
R1036 B.n614 B.n613 10.6151
R1037 B.n613 B.n42 10.6151
R1038 B.n609 B.n42 10.6151
R1039 B.n609 B.n608 10.6151
R1040 B.n608 B.n607 10.6151
R1041 B.n607 B.n44 10.6151
R1042 B.n603 B.n602 10.6151
R1043 B.n602 B.n601 10.6151
R1044 B.n601 B.n49 10.6151
R1045 B.n597 B.n49 10.6151
R1046 B.n597 B.n596 10.6151
R1047 B.n596 B.n595 10.6151
R1048 B.n595 B.n51 10.6151
R1049 B.n591 B.n51 10.6151
R1050 B.n589 B.n588 10.6151
R1051 B.n588 B.n55 10.6151
R1052 B.n584 B.n55 10.6151
R1053 B.n584 B.n583 10.6151
R1054 B.n583 B.n582 10.6151
R1055 B.n582 B.n57 10.6151
R1056 B.n578 B.n57 10.6151
R1057 B.n578 B.n577 10.6151
R1058 B.n577 B.n576 10.6151
R1059 B.n576 B.n59 10.6151
R1060 B.n572 B.n59 10.6151
R1061 B.n572 B.n571 10.6151
R1062 B.n571 B.n570 10.6151
R1063 B.n570 B.n61 10.6151
R1064 B.n566 B.n61 10.6151
R1065 B.n566 B.n565 10.6151
R1066 B.n565 B.n564 10.6151
R1067 B.n564 B.n63 10.6151
R1068 B.n560 B.n63 10.6151
R1069 B.n560 B.n559 10.6151
R1070 B.n559 B.n558 10.6151
R1071 B.n558 B.n65 10.6151
R1072 B.n554 B.n65 10.6151
R1073 B.n554 B.n553 10.6151
R1074 B.n553 B.n552 10.6151
R1075 B.n552 B.n67 10.6151
R1076 B.n548 B.n67 10.6151
R1077 B.n548 B.n547 10.6151
R1078 B.n547 B.n546 10.6151
R1079 B.n546 B.n69 10.6151
R1080 B.n542 B.n69 10.6151
R1081 B.n542 B.n541 10.6151
R1082 B.n541 B.n540 10.6151
R1083 B.n540 B.n71 10.6151
R1084 B.n536 B.n71 10.6151
R1085 B.n536 B.n535 10.6151
R1086 B.n535 B.n534 10.6151
R1087 B.n534 B.n73 10.6151
R1088 B.n530 B.n73 10.6151
R1089 B.n530 B.n529 10.6151
R1090 B.n529 B.n528 10.6151
R1091 B.n528 B.n75 10.6151
R1092 B.n524 B.n75 10.6151
R1093 B.n524 B.n523 10.6151
R1094 B.n523 B.n522 10.6151
R1095 B.n522 B.n77 10.6151
R1096 B.n518 B.n77 10.6151
R1097 B.n518 B.n517 10.6151
R1098 B.n517 B.n516 10.6151
R1099 B.n516 B.n79 10.6151
R1100 B.n512 B.n79 10.6151
R1101 B.n512 B.n511 10.6151
R1102 B.n510 B.n81 10.6151
R1103 B.n506 B.n81 10.6151
R1104 B.n506 B.n505 10.6151
R1105 B.n505 B.n504 10.6151
R1106 B.n504 B.n83 10.6151
R1107 B.n500 B.n83 10.6151
R1108 B.n500 B.n499 10.6151
R1109 B.n499 B.n498 10.6151
R1110 B.n498 B.n85 10.6151
R1111 B.n494 B.n85 10.6151
R1112 B.n494 B.n493 10.6151
R1113 B.n493 B.n492 10.6151
R1114 B.n492 B.n87 10.6151
R1115 B.n488 B.n87 10.6151
R1116 B.n488 B.n487 10.6151
R1117 B.n487 B.n486 10.6151
R1118 B.n486 B.n89 10.6151
R1119 B.n482 B.n89 10.6151
R1120 B.n482 B.n481 10.6151
R1121 B.n481 B.n480 10.6151
R1122 B.n480 B.n91 10.6151
R1123 B.n476 B.n91 10.6151
R1124 B.n476 B.n475 10.6151
R1125 B.n475 B.n474 10.6151
R1126 B.n474 B.n93 10.6151
R1127 B.n470 B.n93 10.6151
R1128 B.n470 B.n469 10.6151
R1129 B.n469 B.n468 10.6151
R1130 B.n468 B.n95 10.6151
R1131 B.n464 B.n95 10.6151
R1132 B.n464 B.n463 10.6151
R1133 B.n463 B.n462 10.6151
R1134 B.n462 B.n97 10.6151
R1135 B.n458 B.n97 10.6151
R1136 B.n458 B.n457 10.6151
R1137 B.n457 B.n456 10.6151
R1138 B.n456 B.n99 10.6151
R1139 B.n452 B.n99 10.6151
R1140 B.n452 B.n451 10.6151
R1141 B.n451 B.n450 10.6151
R1142 B.n450 B.n101 10.6151
R1143 B.n446 B.n101 10.6151
R1144 B.n446 B.n445 10.6151
R1145 B.n445 B.n444 10.6151
R1146 B.n444 B.n103 10.6151
R1147 B.n440 B.n103 10.6151
R1148 B.n440 B.n439 10.6151
R1149 B.n439 B.n438 10.6151
R1150 B.n438 B.n105 10.6151
R1151 B.n434 B.n105 10.6151
R1152 B.n434 B.n433 10.6151
R1153 B.n433 B.n432 10.6151
R1154 B.n432 B.n107 10.6151
R1155 B.n428 B.n107 10.6151
R1156 B.n428 B.n427 10.6151
R1157 B.n427 B.n426 10.6151
R1158 B.n426 B.n109 10.6151
R1159 B.n422 B.n109 10.6151
R1160 B.n422 B.n421 10.6151
R1161 B.n421 B.n420 10.6151
R1162 B.n420 B.n111 10.6151
R1163 B.n416 B.n111 10.6151
R1164 B.n416 B.n415 10.6151
R1165 B.n415 B.n414 10.6151
R1166 B.n414 B.n113 10.6151
R1167 B.n191 B.n1 10.6151
R1168 B.n192 B.n191 10.6151
R1169 B.n192 B.n189 10.6151
R1170 B.n196 B.n189 10.6151
R1171 B.n197 B.n196 10.6151
R1172 B.n198 B.n197 10.6151
R1173 B.n198 B.n187 10.6151
R1174 B.n202 B.n187 10.6151
R1175 B.n203 B.n202 10.6151
R1176 B.n204 B.n203 10.6151
R1177 B.n204 B.n185 10.6151
R1178 B.n208 B.n185 10.6151
R1179 B.n209 B.n208 10.6151
R1180 B.n210 B.n209 10.6151
R1181 B.n210 B.n183 10.6151
R1182 B.n214 B.n183 10.6151
R1183 B.n215 B.n214 10.6151
R1184 B.n216 B.n215 10.6151
R1185 B.n216 B.n181 10.6151
R1186 B.n220 B.n181 10.6151
R1187 B.n221 B.n220 10.6151
R1188 B.n222 B.n221 10.6151
R1189 B.n222 B.n179 10.6151
R1190 B.n226 B.n179 10.6151
R1191 B.n227 B.n226 10.6151
R1192 B.n228 B.n227 10.6151
R1193 B.n228 B.n177 10.6151
R1194 B.n232 B.n177 10.6151
R1195 B.n233 B.n232 10.6151
R1196 B.n234 B.n233 10.6151
R1197 B.n234 B.n175 10.6151
R1198 B.n239 B.n238 10.6151
R1199 B.n240 B.n239 10.6151
R1200 B.n240 B.n173 10.6151
R1201 B.n244 B.n173 10.6151
R1202 B.n245 B.n244 10.6151
R1203 B.n246 B.n245 10.6151
R1204 B.n246 B.n171 10.6151
R1205 B.n250 B.n171 10.6151
R1206 B.n251 B.n250 10.6151
R1207 B.n252 B.n251 10.6151
R1208 B.n252 B.n169 10.6151
R1209 B.n256 B.n169 10.6151
R1210 B.n257 B.n256 10.6151
R1211 B.n258 B.n257 10.6151
R1212 B.n258 B.n167 10.6151
R1213 B.n262 B.n167 10.6151
R1214 B.n263 B.n262 10.6151
R1215 B.n264 B.n263 10.6151
R1216 B.n264 B.n165 10.6151
R1217 B.n268 B.n165 10.6151
R1218 B.n269 B.n268 10.6151
R1219 B.n270 B.n269 10.6151
R1220 B.n270 B.n163 10.6151
R1221 B.n274 B.n163 10.6151
R1222 B.n275 B.n274 10.6151
R1223 B.n276 B.n275 10.6151
R1224 B.n276 B.n161 10.6151
R1225 B.n280 B.n161 10.6151
R1226 B.n281 B.n280 10.6151
R1227 B.n282 B.n281 10.6151
R1228 B.n282 B.n159 10.6151
R1229 B.n286 B.n159 10.6151
R1230 B.n287 B.n286 10.6151
R1231 B.n288 B.n287 10.6151
R1232 B.n288 B.n157 10.6151
R1233 B.n292 B.n157 10.6151
R1234 B.n293 B.n292 10.6151
R1235 B.n294 B.n293 10.6151
R1236 B.n294 B.n155 10.6151
R1237 B.n298 B.n155 10.6151
R1238 B.n299 B.n298 10.6151
R1239 B.n300 B.n299 10.6151
R1240 B.n300 B.n153 10.6151
R1241 B.n304 B.n153 10.6151
R1242 B.n305 B.n304 10.6151
R1243 B.n306 B.n305 10.6151
R1244 B.n306 B.n151 10.6151
R1245 B.n310 B.n151 10.6151
R1246 B.n311 B.n310 10.6151
R1247 B.n312 B.n311 10.6151
R1248 B.n312 B.n149 10.6151
R1249 B.n316 B.n149 10.6151
R1250 B.n319 B.n318 10.6151
R1251 B.n319 B.n145 10.6151
R1252 B.n323 B.n145 10.6151
R1253 B.n324 B.n323 10.6151
R1254 B.n325 B.n324 10.6151
R1255 B.n325 B.n143 10.6151
R1256 B.n329 B.n143 10.6151
R1257 B.n330 B.n329 10.6151
R1258 B.n332 B.n139 10.6151
R1259 B.n336 B.n139 10.6151
R1260 B.n337 B.n336 10.6151
R1261 B.n338 B.n337 10.6151
R1262 B.n338 B.n137 10.6151
R1263 B.n342 B.n137 10.6151
R1264 B.n343 B.n342 10.6151
R1265 B.n344 B.n343 10.6151
R1266 B.n344 B.n135 10.6151
R1267 B.n348 B.n135 10.6151
R1268 B.n349 B.n348 10.6151
R1269 B.n350 B.n349 10.6151
R1270 B.n350 B.n133 10.6151
R1271 B.n354 B.n133 10.6151
R1272 B.n355 B.n354 10.6151
R1273 B.n356 B.n355 10.6151
R1274 B.n356 B.n131 10.6151
R1275 B.n360 B.n131 10.6151
R1276 B.n361 B.n360 10.6151
R1277 B.n362 B.n361 10.6151
R1278 B.n362 B.n129 10.6151
R1279 B.n366 B.n129 10.6151
R1280 B.n367 B.n366 10.6151
R1281 B.n368 B.n367 10.6151
R1282 B.n368 B.n127 10.6151
R1283 B.n372 B.n127 10.6151
R1284 B.n373 B.n372 10.6151
R1285 B.n374 B.n373 10.6151
R1286 B.n374 B.n125 10.6151
R1287 B.n378 B.n125 10.6151
R1288 B.n379 B.n378 10.6151
R1289 B.n380 B.n379 10.6151
R1290 B.n380 B.n123 10.6151
R1291 B.n384 B.n123 10.6151
R1292 B.n385 B.n384 10.6151
R1293 B.n386 B.n385 10.6151
R1294 B.n386 B.n121 10.6151
R1295 B.n390 B.n121 10.6151
R1296 B.n391 B.n390 10.6151
R1297 B.n392 B.n391 10.6151
R1298 B.n392 B.n119 10.6151
R1299 B.n396 B.n119 10.6151
R1300 B.n397 B.n396 10.6151
R1301 B.n398 B.n397 10.6151
R1302 B.n398 B.n117 10.6151
R1303 B.n402 B.n117 10.6151
R1304 B.n403 B.n402 10.6151
R1305 B.n404 B.n403 10.6151
R1306 B.n404 B.n115 10.6151
R1307 B.n408 B.n115 10.6151
R1308 B.n409 B.n408 10.6151
R1309 B.n410 B.n409 10.6151
R1310 B.n733 B.n0 8.11757
R1311 B.n733 B.n1 8.11757
R1312 B.n603 B.n48 6.5566
R1313 B.n591 B.n590 6.5566
R1314 B.n318 B.n317 6.5566
R1315 B.n331 B.n330 6.5566
R1316 B.n48 B.n44 4.05904
R1317 B.n590 B.n589 4.05904
R1318 B.n317 B.n316 4.05904
R1319 B.n332 B.n331 4.05904
C0 VDD2 VDD1 1.2001f
C1 B VDD2 2.1995f
C2 B VDD1 2.1414f
C3 VTAIL VP 10.444099f
C4 VTAIL VN 10.4294f
C5 VN VP 6.83187f
C6 VDD2 w_n2638_n4128# 2.53252f
C7 w_n2638_n4128# VDD1 2.46902f
C8 B w_n2638_n4128# 9.02255f
C9 VTAIL VDD2 14.9861f
C10 VTAIL VDD1 14.95f
C11 VDD2 VP 0.388176f
C12 VDD1 VP 10.809999f
C13 VDD2 VN 10.5775f
C14 VN VDD1 0.150155f
C15 VTAIL B 3.68543f
C16 B VP 1.49925f
C17 B VN 0.938194f
C18 VTAIL w_n2638_n4128# 3.60943f
C19 w_n2638_n4128# VP 5.58674f
C20 VN w_n2638_n4128# 5.24803f
C21 VDD2 VSUBS 1.707074f
C22 VDD1 VSUBS 1.420255f
C23 VTAIL VSUBS 1.022405f
C24 VN VSUBS 5.60146f
C25 VP VSUBS 2.430526f
C26 B VSUBS 3.779438f
C27 w_n2638_n4128# VSUBS 0.13343p
C28 B.n0 VSUBS 0.007815f
C29 B.n1 VSUBS 0.007815f
C30 B.n2 VSUBS 0.011558f
C31 B.n3 VSUBS 0.008857f
C32 B.n4 VSUBS 0.008857f
C33 B.n5 VSUBS 0.008857f
C34 B.n6 VSUBS 0.008857f
C35 B.n7 VSUBS 0.008857f
C36 B.n8 VSUBS 0.008857f
C37 B.n9 VSUBS 0.008857f
C38 B.n10 VSUBS 0.008857f
C39 B.n11 VSUBS 0.008857f
C40 B.n12 VSUBS 0.008857f
C41 B.n13 VSUBS 0.008857f
C42 B.n14 VSUBS 0.008857f
C43 B.n15 VSUBS 0.008857f
C44 B.n16 VSUBS 0.008857f
C45 B.n17 VSUBS 0.008857f
C46 B.n18 VSUBS 0.022136f
C47 B.n19 VSUBS 0.008857f
C48 B.n20 VSUBS 0.008857f
C49 B.n21 VSUBS 0.008857f
C50 B.n22 VSUBS 0.008857f
C51 B.n23 VSUBS 0.008857f
C52 B.n24 VSUBS 0.008857f
C53 B.n25 VSUBS 0.008857f
C54 B.n26 VSUBS 0.008857f
C55 B.n27 VSUBS 0.008857f
C56 B.n28 VSUBS 0.008857f
C57 B.n29 VSUBS 0.008857f
C58 B.n30 VSUBS 0.008857f
C59 B.n31 VSUBS 0.008857f
C60 B.n32 VSUBS 0.008857f
C61 B.n33 VSUBS 0.008857f
C62 B.n34 VSUBS 0.008857f
C63 B.n35 VSUBS 0.008857f
C64 B.n36 VSUBS 0.008857f
C65 B.n37 VSUBS 0.008857f
C66 B.n38 VSUBS 0.008857f
C67 B.n39 VSUBS 0.008857f
C68 B.n40 VSUBS 0.008857f
C69 B.n41 VSUBS 0.008857f
C70 B.n42 VSUBS 0.008857f
C71 B.n43 VSUBS 0.008857f
C72 B.n44 VSUBS 0.006122f
C73 B.n45 VSUBS 0.008857f
C74 B.t10 VSUBS 0.668361f
C75 B.t11 VSUBS 0.682268f
C76 B.t9 VSUBS 0.885266f
C77 B.n46 VSUBS 0.256834f
C78 B.n47 VSUBS 0.083045f
C79 B.n48 VSUBS 0.020521f
C80 B.n49 VSUBS 0.008857f
C81 B.n50 VSUBS 0.008857f
C82 B.n51 VSUBS 0.008857f
C83 B.n52 VSUBS 0.008857f
C84 B.t7 VSUBS 0.668341f
C85 B.t8 VSUBS 0.68225f
C86 B.t6 VSUBS 0.885266f
C87 B.n53 VSUBS 0.256852f
C88 B.n54 VSUBS 0.083065f
C89 B.n55 VSUBS 0.008857f
C90 B.n56 VSUBS 0.008857f
C91 B.n57 VSUBS 0.008857f
C92 B.n58 VSUBS 0.008857f
C93 B.n59 VSUBS 0.008857f
C94 B.n60 VSUBS 0.008857f
C95 B.n61 VSUBS 0.008857f
C96 B.n62 VSUBS 0.008857f
C97 B.n63 VSUBS 0.008857f
C98 B.n64 VSUBS 0.008857f
C99 B.n65 VSUBS 0.008857f
C100 B.n66 VSUBS 0.008857f
C101 B.n67 VSUBS 0.008857f
C102 B.n68 VSUBS 0.008857f
C103 B.n69 VSUBS 0.008857f
C104 B.n70 VSUBS 0.008857f
C105 B.n71 VSUBS 0.008857f
C106 B.n72 VSUBS 0.008857f
C107 B.n73 VSUBS 0.008857f
C108 B.n74 VSUBS 0.008857f
C109 B.n75 VSUBS 0.008857f
C110 B.n76 VSUBS 0.008857f
C111 B.n77 VSUBS 0.008857f
C112 B.n78 VSUBS 0.008857f
C113 B.n79 VSUBS 0.008857f
C114 B.n80 VSUBS 0.022136f
C115 B.n81 VSUBS 0.008857f
C116 B.n82 VSUBS 0.008857f
C117 B.n83 VSUBS 0.008857f
C118 B.n84 VSUBS 0.008857f
C119 B.n85 VSUBS 0.008857f
C120 B.n86 VSUBS 0.008857f
C121 B.n87 VSUBS 0.008857f
C122 B.n88 VSUBS 0.008857f
C123 B.n89 VSUBS 0.008857f
C124 B.n90 VSUBS 0.008857f
C125 B.n91 VSUBS 0.008857f
C126 B.n92 VSUBS 0.008857f
C127 B.n93 VSUBS 0.008857f
C128 B.n94 VSUBS 0.008857f
C129 B.n95 VSUBS 0.008857f
C130 B.n96 VSUBS 0.008857f
C131 B.n97 VSUBS 0.008857f
C132 B.n98 VSUBS 0.008857f
C133 B.n99 VSUBS 0.008857f
C134 B.n100 VSUBS 0.008857f
C135 B.n101 VSUBS 0.008857f
C136 B.n102 VSUBS 0.008857f
C137 B.n103 VSUBS 0.008857f
C138 B.n104 VSUBS 0.008857f
C139 B.n105 VSUBS 0.008857f
C140 B.n106 VSUBS 0.008857f
C141 B.n107 VSUBS 0.008857f
C142 B.n108 VSUBS 0.008857f
C143 B.n109 VSUBS 0.008857f
C144 B.n110 VSUBS 0.008857f
C145 B.n111 VSUBS 0.008857f
C146 B.n112 VSUBS 0.008857f
C147 B.n113 VSUBS 0.022088f
C148 B.n114 VSUBS 0.008857f
C149 B.n115 VSUBS 0.008857f
C150 B.n116 VSUBS 0.008857f
C151 B.n117 VSUBS 0.008857f
C152 B.n118 VSUBS 0.008857f
C153 B.n119 VSUBS 0.008857f
C154 B.n120 VSUBS 0.008857f
C155 B.n121 VSUBS 0.008857f
C156 B.n122 VSUBS 0.008857f
C157 B.n123 VSUBS 0.008857f
C158 B.n124 VSUBS 0.008857f
C159 B.n125 VSUBS 0.008857f
C160 B.n126 VSUBS 0.008857f
C161 B.n127 VSUBS 0.008857f
C162 B.n128 VSUBS 0.008857f
C163 B.n129 VSUBS 0.008857f
C164 B.n130 VSUBS 0.008857f
C165 B.n131 VSUBS 0.008857f
C166 B.n132 VSUBS 0.008857f
C167 B.n133 VSUBS 0.008857f
C168 B.n134 VSUBS 0.008857f
C169 B.n135 VSUBS 0.008857f
C170 B.n136 VSUBS 0.008857f
C171 B.n137 VSUBS 0.008857f
C172 B.n138 VSUBS 0.008857f
C173 B.n139 VSUBS 0.008857f
C174 B.n140 VSUBS 0.008857f
C175 B.t2 VSUBS 0.668341f
C176 B.t1 VSUBS 0.68225f
C177 B.t0 VSUBS 0.885266f
C178 B.n141 VSUBS 0.256852f
C179 B.n142 VSUBS 0.083065f
C180 B.n143 VSUBS 0.008857f
C181 B.n144 VSUBS 0.008857f
C182 B.n145 VSUBS 0.008857f
C183 B.n146 VSUBS 0.008857f
C184 B.t5 VSUBS 0.668361f
C185 B.t4 VSUBS 0.682268f
C186 B.t3 VSUBS 0.885266f
C187 B.n147 VSUBS 0.256834f
C188 B.n148 VSUBS 0.083045f
C189 B.n149 VSUBS 0.008857f
C190 B.n150 VSUBS 0.008857f
C191 B.n151 VSUBS 0.008857f
C192 B.n152 VSUBS 0.008857f
C193 B.n153 VSUBS 0.008857f
C194 B.n154 VSUBS 0.008857f
C195 B.n155 VSUBS 0.008857f
C196 B.n156 VSUBS 0.008857f
C197 B.n157 VSUBS 0.008857f
C198 B.n158 VSUBS 0.008857f
C199 B.n159 VSUBS 0.008857f
C200 B.n160 VSUBS 0.008857f
C201 B.n161 VSUBS 0.008857f
C202 B.n162 VSUBS 0.008857f
C203 B.n163 VSUBS 0.008857f
C204 B.n164 VSUBS 0.008857f
C205 B.n165 VSUBS 0.008857f
C206 B.n166 VSUBS 0.008857f
C207 B.n167 VSUBS 0.008857f
C208 B.n168 VSUBS 0.008857f
C209 B.n169 VSUBS 0.008857f
C210 B.n170 VSUBS 0.008857f
C211 B.n171 VSUBS 0.008857f
C212 B.n172 VSUBS 0.008857f
C213 B.n173 VSUBS 0.008857f
C214 B.n174 VSUBS 0.008857f
C215 B.n175 VSUBS 0.021107f
C216 B.n176 VSUBS 0.008857f
C217 B.n177 VSUBS 0.008857f
C218 B.n178 VSUBS 0.008857f
C219 B.n179 VSUBS 0.008857f
C220 B.n180 VSUBS 0.008857f
C221 B.n181 VSUBS 0.008857f
C222 B.n182 VSUBS 0.008857f
C223 B.n183 VSUBS 0.008857f
C224 B.n184 VSUBS 0.008857f
C225 B.n185 VSUBS 0.008857f
C226 B.n186 VSUBS 0.008857f
C227 B.n187 VSUBS 0.008857f
C228 B.n188 VSUBS 0.008857f
C229 B.n189 VSUBS 0.008857f
C230 B.n190 VSUBS 0.008857f
C231 B.n191 VSUBS 0.008857f
C232 B.n192 VSUBS 0.008857f
C233 B.n193 VSUBS 0.008857f
C234 B.n194 VSUBS 0.008857f
C235 B.n195 VSUBS 0.008857f
C236 B.n196 VSUBS 0.008857f
C237 B.n197 VSUBS 0.008857f
C238 B.n198 VSUBS 0.008857f
C239 B.n199 VSUBS 0.008857f
C240 B.n200 VSUBS 0.008857f
C241 B.n201 VSUBS 0.008857f
C242 B.n202 VSUBS 0.008857f
C243 B.n203 VSUBS 0.008857f
C244 B.n204 VSUBS 0.008857f
C245 B.n205 VSUBS 0.008857f
C246 B.n206 VSUBS 0.008857f
C247 B.n207 VSUBS 0.008857f
C248 B.n208 VSUBS 0.008857f
C249 B.n209 VSUBS 0.008857f
C250 B.n210 VSUBS 0.008857f
C251 B.n211 VSUBS 0.008857f
C252 B.n212 VSUBS 0.008857f
C253 B.n213 VSUBS 0.008857f
C254 B.n214 VSUBS 0.008857f
C255 B.n215 VSUBS 0.008857f
C256 B.n216 VSUBS 0.008857f
C257 B.n217 VSUBS 0.008857f
C258 B.n218 VSUBS 0.008857f
C259 B.n219 VSUBS 0.008857f
C260 B.n220 VSUBS 0.008857f
C261 B.n221 VSUBS 0.008857f
C262 B.n222 VSUBS 0.008857f
C263 B.n223 VSUBS 0.008857f
C264 B.n224 VSUBS 0.008857f
C265 B.n225 VSUBS 0.008857f
C266 B.n226 VSUBS 0.008857f
C267 B.n227 VSUBS 0.008857f
C268 B.n228 VSUBS 0.008857f
C269 B.n229 VSUBS 0.008857f
C270 B.n230 VSUBS 0.008857f
C271 B.n231 VSUBS 0.008857f
C272 B.n232 VSUBS 0.008857f
C273 B.n233 VSUBS 0.008857f
C274 B.n234 VSUBS 0.008857f
C275 B.n235 VSUBS 0.008857f
C276 B.n236 VSUBS 0.021107f
C277 B.n237 VSUBS 0.022136f
C278 B.n238 VSUBS 0.022136f
C279 B.n239 VSUBS 0.008857f
C280 B.n240 VSUBS 0.008857f
C281 B.n241 VSUBS 0.008857f
C282 B.n242 VSUBS 0.008857f
C283 B.n243 VSUBS 0.008857f
C284 B.n244 VSUBS 0.008857f
C285 B.n245 VSUBS 0.008857f
C286 B.n246 VSUBS 0.008857f
C287 B.n247 VSUBS 0.008857f
C288 B.n248 VSUBS 0.008857f
C289 B.n249 VSUBS 0.008857f
C290 B.n250 VSUBS 0.008857f
C291 B.n251 VSUBS 0.008857f
C292 B.n252 VSUBS 0.008857f
C293 B.n253 VSUBS 0.008857f
C294 B.n254 VSUBS 0.008857f
C295 B.n255 VSUBS 0.008857f
C296 B.n256 VSUBS 0.008857f
C297 B.n257 VSUBS 0.008857f
C298 B.n258 VSUBS 0.008857f
C299 B.n259 VSUBS 0.008857f
C300 B.n260 VSUBS 0.008857f
C301 B.n261 VSUBS 0.008857f
C302 B.n262 VSUBS 0.008857f
C303 B.n263 VSUBS 0.008857f
C304 B.n264 VSUBS 0.008857f
C305 B.n265 VSUBS 0.008857f
C306 B.n266 VSUBS 0.008857f
C307 B.n267 VSUBS 0.008857f
C308 B.n268 VSUBS 0.008857f
C309 B.n269 VSUBS 0.008857f
C310 B.n270 VSUBS 0.008857f
C311 B.n271 VSUBS 0.008857f
C312 B.n272 VSUBS 0.008857f
C313 B.n273 VSUBS 0.008857f
C314 B.n274 VSUBS 0.008857f
C315 B.n275 VSUBS 0.008857f
C316 B.n276 VSUBS 0.008857f
C317 B.n277 VSUBS 0.008857f
C318 B.n278 VSUBS 0.008857f
C319 B.n279 VSUBS 0.008857f
C320 B.n280 VSUBS 0.008857f
C321 B.n281 VSUBS 0.008857f
C322 B.n282 VSUBS 0.008857f
C323 B.n283 VSUBS 0.008857f
C324 B.n284 VSUBS 0.008857f
C325 B.n285 VSUBS 0.008857f
C326 B.n286 VSUBS 0.008857f
C327 B.n287 VSUBS 0.008857f
C328 B.n288 VSUBS 0.008857f
C329 B.n289 VSUBS 0.008857f
C330 B.n290 VSUBS 0.008857f
C331 B.n291 VSUBS 0.008857f
C332 B.n292 VSUBS 0.008857f
C333 B.n293 VSUBS 0.008857f
C334 B.n294 VSUBS 0.008857f
C335 B.n295 VSUBS 0.008857f
C336 B.n296 VSUBS 0.008857f
C337 B.n297 VSUBS 0.008857f
C338 B.n298 VSUBS 0.008857f
C339 B.n299 VSUBS 0.008857f
C340 B.n300 VSUBS 0.008857f
C341 B.n301 VSUBS 0.008857f
C342 B.n302 VSUBS 0.008857f
C343 B.n303 VSUBS 0.008857f
C344 B.n304 VSUBS 0.008857f
C345 B.n305 VSUBS 0.008857f
C346 B.n306 VSUBS 0.008857f
C347 B.n307 VSUBS 0.008857f
C348 B.n308 VSUBS 0.008857f
C349 B.n309 VSUBS 0.008857f
C350 B.n310 VSUBS 0.008857f
C351 B.n311 VSUBS 0.008857f
C352 B.n312 VSUBS 0.008857f
C353 B.n313 VSUBS 0.008857f
C354 B.n314 VSUBS 0.008857f
C355 B.n315 VSUBS 0.008857f
C356 B.n316 VSUBS 0.006122f
C357 B.n317 VSUBS 0.020521f
C358 B.n318 VSUBS 0.007164f
C359 B.n319 VSUBS 0.008857f
C360 B.n320 VSUBS 0.008857f
C361 B.n321 VSUBS 0.008857f
C362 B.n322 VSUBS 0.008857f
C363 B.n323 VSUBS 0.008857f
C364 B.n324 VSUBS 0.008857f
C365 B.n325 VSUBS 0.008857f
C366 B.n326 VSUBS 0.008857f
C367 B.n327 VSUBS 0.008857f
C368 B.n328 VSUBS 0.008857f
C369 B.n329 VSUBS 0.008857f
C370 B.n330 VSUBS 0.007164f
C371 B.n331 VSUBS 0.020521f
C372 B.n332 VSUBS 0.006122f
C373 B.n333 VSUBS 0.008857f
C374 B.n334 VSUBS 0.008857f
C375 B.n335 VSUBS 0.008857f
C376 B.n336 VSUBS 0.008857f
C377 B.n337 VSUBS 0.008857f
C378 B.n338 VSUBS 0.008857f
C379 B.n339 VSUBS 0.008857f
C380 B.n340 VSUBS 0.008857f
C381 B.n341 VSUBS 0.008857f
C382 B.n342 VSUBS 0.008857f
C383 B.n343 VSUBS 0.008857f
C384 B.n344 VSUBS 0.008857f
C385 B.n345 VSUBS 0.008857f
C386 B.n346 VSUBS 0.008857f
C387 B.n347 VSUBS 0.008857f
C388 B.n348 VSUBS 0.008857f
C389 B.n349 VSUBS 0.008857f
C390 B.n350 VSUBS 0.008857f
C391 B.n351 VSUBS 0.008857f
C392 B.n352 VSUBS 0.008857f
C393 B.n353 VSUBS 0.008857f
C394 B.n354 VSUBS 0.008857f
C395 B.n355 VSUBS 0.008857f
C396 B.n356 VSUBS 0.008857f
C397 B.n357 VSUBS 0.008857f
C398 B.n358 VSUBS 0.008857f
C399 B.n359 VSUBS 0.008857f
C400 B.n360 VSUBS 0.008857f
C401 B.n361 VSUBS 0.008857f
C402 B.n362 VSUBS 0.008857f
C403 B.n363 VSUBS 0.008857f
C404 B.n364 VSUBS 0.008857f
C405 B.n365 VSUBS 0.008857f
C406 B.n366 VSUBS 0.008857f
C407 B.n367 VSUBS 0.008857f
C408 B.n368 VSUBS 0.008857f
C409 B.n369 VSUBS 0.008857f
C410 B.n370 VSUBS 0.008857f
C411 B.n371 VSUBS 0.008857f
C412 B.n372 VSUBS 0.008857f
C413 B.n373 VSUBS 0.008857f
C414 B.n374 VSUBS 0.008857f
C415 B.n375 VSUBS 0.008857f
C416 B.n376 VSUBS 0.008857f
C417 B.n377 VSUBS 0.008857f
C418 B.n378 VSUBS 0.008857f
C419 B.n379 VSUBS 0.008857f
C420 B.n380 VSUBS 0.008857f
C421 B.n381 VSUBS 0.008857f
C422 B.n382 VSUBS 0.008857f
C423 B.n383 VSUBS 0.008857f
C424 B.n384 VSUBS 0.008857f
C425 B.n385 VSUBS 0.008857f
C426 B.n386 VSUBS 0.008857f
C427 B.n387 VSUBS 0.008857f
C428 B.n388 VSUBS 0.008857f
C429 B.n389 VSUBS 0.008857f
C430 B.n390 VSUBS 0.008857f
C431 B.n391 VSUBS 0.008857f
C432 B.n392 VSUBS 0.008857f
C433 B.n393 VSUBS 0.008857f
C434 B.n394 VSUBS 0.008857f
C435 B.n395 VSUBS 0.008857f
C436 B.n396 VSUBS 0.008857f
C437 B.n397 VSUBS 0.008857f
C438 B.n398 VSUBS 0.008857f
C439 B.n399 VSUBS 0.008857f
C440 B.n400 VSUBS 0.008857f
C441 B.n401 VSUBS 0.008857f
C442 B.n402 VSUBS 0.008857f
C443 B.n403 VSUBS 0.008857f
C444 B.n404 VSUBS 0.008857f
C445 B.n405 VSUBS 0.008857f
C446 B.n406 VSUBS 0.008857f
C447 B.n407 VSUBS 0.008857f
C448 B.n408 VSUBS 0.008857f
C449 B.n409 VSUBS 0.008857f
C450 B.n410 VSUBS 0.021154f
C451 B.n411 VSUBS 0.022136f
C452 B.n412 VSUBS 0.021107f
C453 B.n413 VSUBS 0.008857f
C454 B.n414 VSUBS 0.008857f
C455 B.n415 VSUBS 0.008857f
C456 B.n416 VSUBS 0.008857f
C457 B.n417 VSUBS 0.008857f
C458 B.n418 VSUBS 0.008857f
C459 B.n419 VSUBS 0.008857f
C460 B.n420 VSUBS 0.008857f
C461 B.n421 VSUBS 0.008857f
C462 B.n422 VSUBS 0.008857f
C463 B.n423 VSUBS 0.008857f
C464 B.n424 VSUBS 0.008857f
C465 B.n425 VSUBS 0.008857f
C466 B.n426 VSUBS 0.008857f
C467 B.n427 VSUBS 0.008857f
C468 B.n428 VSUBS 0.008857f
C469 B.n429 VSUBS 0.008857f
C470 B.n430 VSUBS 0.008857f
C471 B.n431 VSUBS 0.008857f
C472 B.n432 VSUBS 0.008857f
C473 B.n433 VSUBS 0.008857f
C474 B.n434 VSUBS 0.008857f
C475 B.n435 VSUBS 0.008857f
C476 B.n436 VSUBS 0.008857f
C477 B.n437 VSUBS 0.008857f
C478 B.n438 VSUBS 0.008857f
C479 B.n439 VSUBS 0.008857f
C480 B.n440 VSUBS 0.008857f
C481 B.n441 VSUBS 0.008857f
C482 B.n442 VSUBS 0.008857f
C483 B.n443 VSUBS 0.008857f
C484 B.n444 VSUBS 0.008857f
C485 B.n445 VSUBS 0.008857f
C486 B.n446 VSUBS 0.008857f
C487 B.n447 VSUBS 0.008857f
C488 B.n448 VSUBS 0.008857f
C489 B.n449 VSUBS 0.008857f
C490 B.n450 VSUBS 0.008857f
C491 B.n451 VSUBS 0.008857f
C492 B.n452 VSUBS 0.008857f
C493 B.n453 VSUBS 0.008857f
C494 B.n454 VSUBS 0.008857f
C495 B.n455 VSUBS 0.008857f
C496 B.n456 VSUBS 0.008857f
C497 B.n457 VSUBS 0.008857f
C498 B.n458 VSUBS 0.008857f
C499 B.n459 VSUBS 0.008857f
C500 B.n460 VSUBS 0.008857f
C501 B.n461 VSUBS 0.008857f
C502 B.n462 VSUBS 0.008857f
C503 B.n463 VSUBS 0.008857f
C504 B.n464 VSUBS 0.008857f
C505 B.n465 VSUBS 0.008857f
C506 B.n466 VSUBS 0.008857f
C507 B.n467 VSUBS 0.008857f
C508 B.n468 VSUBS 0.008857f
C509 B.n469 VSUBS 0.008857f
C510 B.n470 VSUBS 0.008857f
C511 B.n471 VSUBS 0.008857f
C512 B.n472 VSUBS 0.008857f
C513 B.n473 VSUBS 0.008857f
C514 B.n474 VSUBS 0.008857f
C515 B.n475 VSUBS 0.008857f
C516 B.n476 VSUBS 0.008857f
C517 B.n477 VSUBS 0.008857f
C518 B.n478 VSUBS 0.008857f
C519 B.n479 VSUBS 0.008857f
C520 B.n480 VSUBS 0.008857f
C521 B.n481 VSUBS 0.008857f
C522 B.n482 VSUBS 0.008857f
C523 B.n483 VSUBS 0.008857f
C524 B.n484 VSUBS 0.008857f
C525 B.n485 VSUBS 0.008857f
C526 B.n486 VSUBS 0.008857f
C527 B.n487 VSUBS 0.008857f
C528 B.n488 VSUBS 0.008857f
C529 B.n489 VSUBS 0.008857f
C530 B.n490 VSUBS 0.008857f
C531 B.n491 VSUBS 0.008857f
C532 B.n492 VSUBS 0.008857f
C533 B.n493 VSUBS 0.008857f
C534 B.n494 VSUBS 0.008857f
C535 B.n495 VSUBS 0.008857f
C536 B.n496 VSUBS 0.008857f
C537 B.n497 VSUBS 0.008857f
C538 B.n498 VSUBS 0.008857f
C539 B.n499 VSUBS 0.008857f
C540 B.n500 VSUBS 0.008857f
C541 B.n501 VSUBS 0.008857f
C542 B.n502 VSUBS 0.008857f
C543 B.n503 VSUBS 0.008857f
C544 B.n504 VSUBS 0.008857f
C545 B.n505 VSUBS 0.008857f
C546 B.n506 VSUBS 0.008857f
C547 B.n507 VSUBS 0.008857f
C548 B.n508 VSUBS 0.008857f
C549 B.n509 VSUBS 0.021107f
C550 B.n510 VSUBS 0.021107f
C551 B.n511 VSUBS 0.022136f
C552 B.n512 VSUBS 0.008857f
C553 B.n513 VSUBS 0.008857f
C554 B.n514 VSUBS 0.008857f
C555 B.n515 VSUBS 0.008857f
C556 B.n516 VSUBS 0.008857f
C557 B.n517 VSUBS 0.008857f
C558 B.n518 VSUBS 0.008857f
C559 B.n519 VSUBS 0.008857f
C560 B.n520 VSUBS 0.008857f
C561 B.n521 VSUBS 0.008857f
C562 B.n522 VSUBS 0.008857f
C563 B.n523 VSUBS 0.008857f
C564 B.n524 VSUBS 0.008857f
C565 B.n525 VSUBS 0.008857f
C566 B.n526 VSUBS 0.008857f
C567 B.n527 VSUBS 0.008857f
C568 B.n528 VSUBS 0.008857f
C569 B.n529 VSUBS 0.008857f
C570 B.n530 VSUBS 0.008857f
C571 B.n531 VSUBS 0.008857f
C572 B.n532 VSUBS 0.008857f
C573 B.n533 VSUBS 0.008857f
C574 B.n534 VSUBS 0.008857f
C575 B.n535 VSUBS 0.008857f
C576 B.n536 VSUBS 0.008857f
C577 B.n537 VSUBS 0.008857f
C578 B.n538 VSUBS 0.008857f
C579 B.n539 VSUBS 0.008857f
C580 B.n540 VSUBS 0.008857f
C581 B.n541 VSUBS 0.008857f
C582 B.n542 VSUBS 0.008857f
C583 B.n543 VSUBS 0.008857f
C584 B.n544 VSUBS 0.008857f
C585 B.n545 VSUBS 0.008857f
C586 B.n546 VSUBS 0.008857f
C587 B.n547 VSUBS 0.008857f
C588 B.n548 VSUBS 0.008857f
C589 B.n549 VSUBS 0.008857f
C590 B.n550 VSUBS 0.008857f
C591 B.n551 VSUBS 0.008857f
C592 B.n552 VSUBS 0.008857f
C593 B.n553 VSUBS 0.008857f
C594 B.n554 VSUBS 0.008857f
C595 B.n555 VSUBS 0.008857f
C596 B.n556 VSUBS 0.008857f
C597 B.n557 VSUBS 0.008857f
C598 B.n558 VSUBS 0.008857f
C599 B.n559 VSUBS 0.008857f
C600 B.n560 VSUBS 0.008857f
C601 B.n561 VSUBS 0.008857f
C602 B.n562 VSUBS 0.008857f
C603 B.n563 VSUBS 0.008857f
C604 B.n564 VSUBS 0.008857f
C605 B.n565 VSUBS 0.008857f
C606 B.n566 VSUBS 0.008857f
C607 B.n567 VSUBS 0.008857f
C608 B.n568 VSUBS 0.008857f
C609 B.n569 VSUBS 0.008857f
C610 B.n570 VSUBS 0.008857f
C611 B.n571 VSUBS 0.008857f
C612 B.n572 VSUBS 0.008857f
C613 B.n573 VSUBS 0.008857f
C614 B.n574 VSUBS 0.008857f
C615 B.n575 VSUBS 0.008857f
C616 B.n576 VSUBS 0.008857f
C617 B.n577 VSUBS 0.008857f
C618 B.n578 VSUBS 0.008857f
C619 B.n579 VSUBS 0.008857f
C620 B.n580 VSUBS 0.008857f
C621 B.n581 VSUBS 0.008857f
C622 B.n582 VSUBS 0.008857f
C623 B.n583 VSUBS 0.008857f
C624 B.n584 VSUBS 0.008857f
C625 B.n585 VSUBS 0.008857f
C626 B.n586 VSUBS 0.008857f
C627 B.n587 VSUBS 0.008857f
C628 B.n588 VSUBS 0.008857f
C629 B.n589 VSUBS 0.006122f
C630 B.n590 VSUBS 0.020521f
C631 B.n591 VSUBS 0.007164f
C632 B.n592 VSUBS 0.008857f
C633 B.n593 VSUBS 0.008857f
C634 B.n594 VSUBS 0.008857f
C635 B.n595 VSUBS 0.008857f
C636 B.n596 VSUBS 0.008857f
C637 B.n597 VSUBS 0.008857f
C638 B.n598 VSUBS 0.008857f
C639 B.n599 VSUBS 0.008857f
C640 B.n600 VSUBS 0.008857f
C641 B.n601 VSUBS 0.008857f
C642 B.n602 VSUBS 0.008857f
C643 B.n603 VSUBS 0.007164f
C644 B.n604 VSUBS 0.008857f
C645 B.n605 VSUBS 0.008857f
C646 B.n606 VSUBS 0.008857f
C647 B.n607 VSUBS 0.008857f
C648 B.n608 VSUBS 0.008857f
C649 B.n609 VSUBS 0.008857f
C650 B.n610 VSUBS 0.008857f
C651 B.n611 VSUBS 0.008857f
C652 B.n612 VSUBS 0.008857f
C653 B.n613 VSUBS 0.008857f
C654 B.n614 VSUBS 0.008857f
C655 B.n615 VSUBS 0.008857f
C656 B.n616 VSUBS 0.008857f
C657 B.n617 VSUBS 0.008857f
C658 B.n618 VSUBS 0.008857f
C659 B.n619 VSUBS 0.008857f
C660 B.n620 VSUBS 0.008857f
C661 B.n621 VSUBS 0.008857f
C662 B.n622 VSUBS 0.008857f
C663 B.n623 VSUBS 0.008857f
C664 B.n624 VSUBS 0.008857f
C665 B.n625 VSUBS 0.008857f
C666 B.n626 VSUBS 0.008857f
C667 B.n627 VSUBS 0.008857f
C668 B.n628 VSUBS 0.008857f
C669 B.n629 VSUBS 0.008857f
C670 B.n630 VSUBS 0.008857f
C671 B.n631 VSUBS 0.008857f
C672 B.n632 VSUBS 0.008857f
C673 B.n633 VSUBS 0.008857f
C674 B.n634 VSUBS 0.008857f
C675 B.n635 VSUBS 0.008857f
C676 B.n636 VSUBS 0.008857f
C677 B.n637 VSUBS 0.008857f
C678 B.n638 VSUBS 0.008857f
C679 B.n639 VSUBS 0.008857f
C680 B.n640 VSUBS 0.008857f
C681 B.n641 VSUBS 0.008857f
C682 B.n642 VSUBS 0.008857f
C683 B.n643 VSUBS 0.008857f
C684 B.n644 VSUBS 0.008857f
C685 B.n645 VSUBS 0.008857f
C686 B.n646 VSUBS 0.008857f
C687 B.n647 VSUBS 0.008857f
C688 B.n648 VSUBS 0.008857f
C689 B.n649 VSUBS 0.008857f
C690 B.n650 VSUBS 0.008857f
C691 B.n651 VSUBS 0.008857f
C692 B.n652 VSUBS 0.008857f
C693 B.n653 VSUBS 0.008857f
C694 B.n654 VSUBS 0.008857f
C695 B.n655 VSUBS 0.008857f
C696 B.n656 VSUBS 0.008857f
C697 B.n657 VSUBS 0.008857f
C698 B.n658 VSUBS 0.008857f
C699 B.n659 VSUBS 0.008857f
C700 B.n660 VSUBS 0.008857f
C701 B.n661 VSUBS 0.008857f
C702 B.n662 VSUBS 0.008857f
C703 B.n663 VSUBS 0.008857f
C704 B.n664 VSUBS 0.008857f
C705 B.n665 VSUBS 0.008857f
C706 B.n666 VSUBS 0.008857f
C707 B.n667 VSUBS 0.008857f
C708 B.n668 VSUBS 0.008857f
C709 B.n669 VSUBS 0.008857f
C710 B.n670 VSUBS 0.008857f
C711 B.n671 VSUBS 0.008857f
C712 B.n672 VSUBS 0.008857f
C713 B.n673 VSUBS 0.008857f
C714 B.n674 VSUBS 0.008857f
C715 B.n675 VSUBS 0.008857f
C716 B.n676 VSUBS 0.008857f
C717 B.n677 VSUBS 0.008857f
C718 B.n678 VSUBS 0.008857f
C719 B.n679 VSUBS 0.008857f
C720 B.n680 VSUBS 0.008857f
C721 B.n681 VSUBS 0.008857f
C722 B.n682 VSUBS 0.008857f
C723 B.n683 VSUBS 0.022136f
C724 B.n684 VSUBS 0.021107f
C725 B.n685 VSUBS 0.021107f
C726 B.n686 VSUBS 0.008857f
C727 B.n687 VSUBS 0.008857f
C728 B.n688 VSUBS 0.008857f
C729 B.n689 VSUBS 0.008857f
C730 B.n690 VSUBS 0.008857f
C731 B.n691 VSUBS 0.008857f
C732 B.n692 VSUBS 0.008857f
C733 B.n693 VSUBS 0.008857f
C734 B.n694 VSUBS 0.008857f
C735 B.n695 VSUBS 0.008857f
C736 B.n696 VSUBS 0.008857f
C737 B.n697 VSUBS 0.008857f
C738 B.n698 VSUBS 0.008857f
C739 B.n699 VSUBS 0.008857f
C740 B.n700 VSUBS 0.008857f
C741 B.n701 VSUBS 0.008857f
C742 B.n702 VSUBS 0.008857f
C743 B.n703 VSUBS 0.008857f
C744 B.n704 VSUBS 0.008857f
C745 B.n705 VSUBS 0.008857f
C746 B.n706 VSUBS 0.008857f
C747 B.n707 VSUBS 0.008857f
C748 B.n708 VSUBS 0.008857f
C749 B.n709 VSUBS 0.008857f
C750 B.n710 VSUBS 0.008857f
C751 B.n711 VSUBS 0.008857f
C752 B.n712 VSUBS 0.008857f
C753 B.n713 VSUBS 0.008857f
C754 B.n714 VSUBS 0.008857f
C755 B.n715 VSUBS 0.008857f
C756 B.n716 VSUBS 0.008857f
C757 B.n717 VSUBS 0.008857f
C758 B.n718 VSUBS 0.008857f
C759 B.n719 VSUBS 0.008857f
C760 B.n720 VSUBS 0.008857f
C761 B.n721 VSUBS 0.008857f
C762 B.n722 VSUBS 0.008857f
C763 B.n723 VSUBS 0.008857f
C764 B.n724 VSUBS 0.008857f
C765 B.n725 VSUBS 0.008857f
C766 B.n726 VSUBS 0.008857f
C767 B.n727 VSUBS 0.008857f
C768 B.n728 VSUBS 0.008857f
C769 B.n729 VSUBS 0.008857f
C770 B.n730 VSUBS 0.008857f
C771 B.n731 VSUBS 0.011558f
C772 B.n732 VSUBS 0.012312f
C773 B.n733 VSUBS 0.024484f
C774 VDD2.t2 VSUBS 3.64453f
C775 VDD2.t6 VSUBS 0.341433f
C776 VDD2.t5 VSUBS 0.341433f
C777 VDD2.n0 VSUBS 2.79622f
C778 VDD2.n1 VSUBS 1.37347f
C779 VDD2.t9 VSUBS 0.341433f
C780 VDD2.t1 VSUBS 0.341433f
C781 VDD2.n2 VSUBS 2.80453f
C782 VDD2.n3 VSUBS 2.84241f
C783 VDD2.t8 VSUBS 3.63281f
C784 VDD2.n4 VSUBS 3.40447f
C785 VDD2.t0 VSUBS 0.341433f
C786 VDD2.t3 VSUBS 0.341433f
C787 VDD2.n5 VSUBS 2.79622f
C788 VDD2.n6 VSUBS 0.659256f
C789 VDD2.t4 VSUBS 0.341433f
C790 VDD2.t7 VSUBS 0.341433f
C791 VDD2.n7 VSUBS 2.80448f
C792 VN.n0 VSUBS 0.056063f
C793 VN.t0 VSUBS 1.93037f
C794 VN.n1 VSUBS 0.695788f
C795 VN.n2 VSUBS 0.042014f
C796 VN.t4 VSUBS 1.93037f
C797 VN.n3 VSUBS 0.054681f
C798 VN.t7 VSUBS 2.03556f
C799 VN.n4 VSUBS 0.753993f
C800 VN.t3 VSUBS 1.93037f
C801 VN.n5 VSUBS 0.753016f
C802 VN.n6 VSUBS 0.059006f
C803 VN.n7 VSUBS 0.211297f
C804 VN.n8 VSUBS 0.042014f
C805 VN.n9 VSUBS 0.042014f
C806 VN.n10 VSUBS 0.735236f
C807 VN.n11 VSUBS 0.054681f
C808 VN.n12 VSUBS 0.059006f
C809 VN.n13 VSUBS 0.042014f
C810 VN.n14 VSUBS 0.042014f
C811 VN.n15 VSUBS 0.054178f
C812 VN.n16 VSUBS 0.031493f
C813 VN.t8 VSUBS 1.99818f
C814 VN.n17 VSUBS 0.761042f
C815 VN.n18 VSUBS 0.039348f
C816 VN.n19 VSUBS 0.056063f
C817 VN.t9 VSUBS 1.93037f
C818 VN.n20 VSUBS 0.695788f
C819 VN.n21 VSUBS 0.042014f
C820 VN.t6 VSUBS 1.93037f
C821 VN.n22 VSUBS 0.054681f
C822 VN.t2 VSUBS 2.03556f
C823 VN.n23 VSUBS 0.753993f
C824 VN.t5 VSUBS 1.93037f
C825 VN.n24 VSUBS 0.753016f
C826 VN.n25 VSUBS 0.059006f
C827 VN.n26 VSUBS 0.211297f
C828 VN.n27 VSUBS 0.042014f
C829 VN.n28 VSUBS 0.042014f
C830 VN.n29 VSUBS 0.735236f
C831 VN.n30 VSUBS 0.054681f
C832 VN.n31 VSUBS 0.059006f
C833 VN.n32 VSUBS 0.042014f
C834 VN.n33 VSUBS 0.042014f
C835 VN.n34 VSUBS 0.054178f
C836 VN.n35 VSUBS 0.031493f
C837 VN.t1 VSUBS 1.99818f
C838 VN.n36 VSUBS 0.761042f
C839 VN.n37 VSUBS 2.16326f
C840 VDD1.t1 VSUBS 3.63244f
C841 VDD1.t8 VSUBS 0.340299f
C842 VDD1.t5 VSUBS 0.340299f
C843 VDD1.n0 VSUBS 2.78693f
C844 VDD1.n1 VSUBS 1.37627f
C845 VDD1.t4 VSUBS 3.63242f
C846 VDD1.t0 VSUBS 0.340299f
C847 VDD1.t9 VSUBS 0.340299f
C848 VDD1.n2 VSUBS 2.78693f
C849 VDD1.n3 VSUBS 1.36891f
C850 VDD1.t6 VSUBS 0.340299f
C851 VDD1.t3 VSUBS 0.340299f
C852 VDD1.n4 VSUBS 2.79522f
C853 VDD1.n5 VSUBS 2.92777f
C854 VDD1.t7 VSUBS 0.340299f
C855 VDD1.t2 VSUBS 0.340299f
C856 VDD1.n6 VSUBS 2.78692f
C857 VDD1.n7 VSUBS 3.37857f
C858 VTAIL.t4 VSUBS 0.344113f
C859 VTAIL.t1 VSUBS 0.344113f
C860 VTAIL.n0 VSUBS 2.65987f
C861 VTAIL.n1 VSUBS 0.82699f
C862 VTAIL.t11 VSUBS 3.4808f
C863 VTAIL.n2 VSUBS 0.965989f
C864 VTAIL.t15 VSUBS 0.344113f
C865 VTAIL.t17 VSUBS 0.344113f
C866 VTAIL.n3 VSUBS 2.65987f
C867 VTAIL.n4 VSUBS 0.85991f
C868 VTAIL.t13 VSUBS 0.344113f
C869 VTAIL.t10 VSUBS 0.344113f
C870 VTAIL.n5 VSUBS 2.65987f
C871 VTAIL.n6 VSUBS 2.55031f
C872 VTAIL.t6 VSUBS 0.344113f
C873 VTAIL.t8 VSUBS 0.344113f
C874 VTAIL.n7 VSUBS 2.65988f
C875 VTAIL.n8 VSUBS 2.55031f
C876 VTAIL.t2 VSUBS 0.344113f
C877 VTAIL.t0 VSUBS 0.344113f
C878 VTAIL.n9 VSUBS 2.65988f
C879 VTAIL.n10 VSUBS 0.859905f
C880 VTAIL.t9 VSUBS 3.48083f
C881 VTAIL.n11 VSUBS 0.965962f
C882 VTAIL.t14 VSUBS 0.344113f
C883 VTAIL.t18 VSUBS 0.344113f
C884 VTAIL.n12 VSUBS 2.65988f
C885 VTAIL.n13 VSUBS 0.848422f
C886 VTAIL.t19 VSUBS 0.344113f
C887 VTAIL.t12 VSUBS 0.344113f
C888 VTAIL.n14 VSUBS 2.65988f
C889 VTAIL.n15 VSUBS 0.859905f
C890 VTAIL.t16 VSUBS 3.4808f
C891 VTAIL.n16 VSUBS 2.56146f
C892 VTAIL.t5 VSUBS 3.4808f
C893 VTAIL.n17 VSUBS 2.56146f
C894 VTAIL.t3 VSUBS 0.344113f
C895 VTAIL.t7 VSUBS 0.344113f
C896 VTAIL.n18 VSUBS 2.65987f
C897 VTAIL.n19 VSUBS 0.774931f
C898 VP.n0 VSUBS 0.057185f
C899 VP.t3 VSUBS 1.96899f
C900 VP.n1 VSUBS 0.709708f
C901 VP.n2 VSUBS 0.042855f
C902 VP.t0 VSUBS 1.96899f
C903 VP.n3 VSUBS 0.055775f
C904 VP.n4 VSUBS 0.042855f
C905 VP.t9 VSUBS 1.96899f
C906 VP.t5 VSUBS 2.03816f
C907 VP.n5 VSUBS 0.776269f
C908 VP.n6 VSUBS 0.057185f
C909 VP.t7 VSUBS 2.03816f
C910 VP.t2 VSUBS 1.96899f
C911 VP.n7 VSUBS 0.709708f
C912 VP.n8 VSUBS 0.042855f
C913 VP.t4 VSUBS 1.96899f
C914 VP.n9 VSUBS 0.055775f
C915 VP.t8 VSUBS 2.07629f
C916 VP.n10 VSUBS 0.769079f
C917 VP.t1 VSUBS 1.96899f
C918 VP.n11 VSUBS 0.768081f
C919 VP.n12 VSUBS 0.060186f
C920 VP.n13 VSUBS 0.215524f
C921 VP.n14 VSUBS 0.042855f
C922 VP.n15 VSUBS 0.042855f
C923 VP.n16 VSUBS 0.749946f
C924 VP.n17 VSUBS 0.055775f
C925 VP.n18 VSUBS 0.060186f
C926 VP.n19 VSUBS 0.042855f
C927 VP.n20 VSUBS 0.042855f
C928 VP.n21 VSUBS 0.055262f
C929 VP.n22 VSUBS 0.032124f
C930 VP.n23 VSUBS 0.776269f
C931 VP.n24 VSUBS 2.183f
C932 VP.n25 VSUBS 2.2154f
C933 VP.n26 VSUBS 0.057185f
C934 VP.n27 VSUBS 0.032124f
C935 VP.n28 VSUBS 0.055262f
C936 VP.n29 VSUBS 0.709708f
C937 VP.n30 VSUBS 0.060186f
C938 VP.n31 VSUBS 0.042855f
C939 VP.n32 VSUBS 0.042855f
C940 VP.n33 VSUBS 0.042855f
C941 VP.n34 VSUBS 0.749946f
C942 VP.n35 VSUBS 0.055775f
C943 VP.n36 VSUBS 0.060186f
C944 VP.n37 VSUBS 0.042855f
C945 VP.n38 VSUBS 0.042855f
C946 VP.n39 VSUBS 0.055262f
C947 VP.n40 VSUBS 0.032124f
C948 VP.t6 VSUBS 2.03816f
C949 VP.n41 VSUBS 0.776269f
C950 VP.n42 VSUBS 0.040135f
.ends

