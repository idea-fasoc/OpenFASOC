* NGSPICE file created from tg_sample_0008.ext - technology: sky130A

.subckt tg_sample_0008 VIN VGN VGP VSS VCC VOUT
X0 VCC.t18 VCC.t16 VCC.t17 VCC.t6 sky130_fd_pr__pfet_01v8 ad=3.4788 pd=18.62 as=0 ps=0 w=8.92 l=3.54
X1 VCC.t15 VCC.t13 VCC.t14 VCC.t10 sky130_fd_pr__pfet_01v8 ad=3.4788 pd=18.62 as=0 ps=0 w=8.92 l=3.54
X2 VOUT.t33 VOUT.t31 VOUT.t32 VCC.t3 sky130_fd_pr__pfet_01v8 ad=3.4788 pd=18.62 as=0 ps=0 w=8.92 l=3.54
X3 VOUT.t5 VGN.t0 VOUT.t5 VSS.t15 sky130_fd_pr__nfet_01v8 ad=3.15315 pd=19.44 as=0 ps=0 w=19.11 l=0.22
X4 VOUT.t4 VGN.t1 VOUT.t4 VSS.t18 sky130_fd_pr__nfet_01v8 ad=3.15315 pd=19.44 as=0 ps=0 w=19.11 l=0.22
X5 VSS.t13 VSS.t11 VSS.t12 VSS.t8 sky130_fd_pr__nfet_01v8 ad=7.4529 pd=39 as=0 ps=0 w=19.11 l=0.22
X6 VOUT.t3 VGN.t2 VOUT.t2 VSS.t16 sky130_fd_pr__nfet_01v8 ad=7.4529 pd=39 as=0 ps=0 w=19.11 l=0.22
X7 VOUT.t30 VOUT.t29 VOUT.t30 VCC.t0 sky130_fd_pr__pfet_01v8 ad=1.4718 pd=9.25 as=0 ps=0 w=8.92 l=3.54
X8 VCC.t12 VCC.t9 VCC.t11 VCC.t10 sky130_fd_pr__pfet_01v8 ad=3.4788 pd=18.62 as=0 ps=0 w=8.92 l=3.54
X9 VOUT.t1 VGN.t3 VOUT.t1 VSS.t14 sky130_fd_pr__nfet_01v8 ad=3.15315 pd=19.44 as=0 ps=0 w=19.11 l=0.22
X10 VSS.t10 VSS.t7 VSS.t9 VSS.t8 sky130_fd_pr__nfet_01v8 ad=7.4529 pd=39 as=0 ps=0 w=19.11 l=0.22
X11 VOUT.t28 VOUT.t27 VOUT.t28 VCC.t4 sky130_fd_pr__pfet_01v8 ad=1.4718 pd=9.25 as=0 ps=0 w=8.92 l=3.54
X12 VOUT.t6 VGN.t4 VOUT.t6 VSS.t18 sky130_fd_pr__nfet_01v8 ad=3.15315 pd=19.44 as=0 ps=0 w=19.11 l=0.22
X13 VOUT.t26 VOUT.t25 VOUT.t26 VCC.t0 sky130_fd_pr__pfet_01v8 ad=1.4718 pd=9.25 as=0 ps=0 w=8.92 l=3.54
X14 VOUT.t0 VGN.t5 VOUT.t0 VSS.t17 sky130_fd_pr__nfet_01v8 ad=3.15315 pd=19.44 as=0 ps=0 w=19.11 l=0.22
X15 VOUT.t8 VGN.t6 VOUT.t8 VSS.t17 sky130_fd_pr__nfet_01v8 ad=3.15315 pd=19.44 as=0 ps=0 w=19.11 l=0.22
X16 VOUT.t24 VOUT.t23 VOUT.t24 VCC.t4 sky130_fd_pr__pfet_01v8 ad=1.4718 pd=9.25 as=0 ps=0 w=8.92 l=3.54
X17 VOUT.t22 VOUT.t21 VOUT.t22 VCC.t1 sky130_fd_pr__pfet_01v8 ad=1.4718 pd=9.25 as=0 ps=0 w=8.92 l=3.54
X18 VOUT.t20 VOUT.t19 VOUT.t20 VCC.t2 sky130_fd_pr__pfet_01v8 ad=1.4718 pd=9.25 as=0 ps=0 w=8.92 l=3.54
X19 VSS.t6 VSS.t4 VSS.t5 VSS.t1 sky130_fd_pr__nfet_01v8 ad=7.4529 pd=39 as=0 ps=0 w=19.11 l=0.22
X20 VOUT.t11 VGN.t7 VOUT.t10 VSS.t16 sky130_fd_pr__nfet_01v8 ad=7.4529 pd=39 as=0 ps=0 w=19.11 l=0.22
X21 VCC.t8 VCC.t5 VCC.t7 VCC.t6 sky130_fd_pr__pfet_01v8 ad=3.4788 pd=18.62 as=0 ps=0 w=8.92 l=3.54
X22 VSS.t3 VSS.t0 VSS.t2 VSS.t1 sky130_fd_pr__nfet_01v8 ad=7.4529 pd=39 as=0 ps=0 w=19.11 l=0.22
X23 VOUT.t18 VOUT.t16 VOUT.t17 VCC.t3 sky130_fd_pr__pfet_01v8 ad=3.4788 pd=18.62 as=0 ps=0 w=8.92 l=3.54
X24 VOUT.t7 VGN.t8 VOUT.t7 VSS.t15 sky130_fd_pr__nfet_01v8 ad=3.15315 pd=19.44 as=0 ps=0 w=19.11 l=0.22
X25 VOUT.t15 VOUT.t14 VOUT.t15 VCC.t1 sky130_fd_pr__pfet_01v8 ad=1.4718 pd=9.25 as=0 ps=0 w=8.92 l=3.54
X26 VOUT.t13 VOUT.t12 VOUT.t13 VCC.t2 sky130_fd_pr__pfet_01v8 ad=1.4718 pd=9.25 as=0 ps=0 w=8.92 l=3.54
X27 VOUT.t9 VGN.t9 VOUT.t9 VSS.t14 sky130_fd_pr__nfet_01v8 ad=3.15315 pd=19.44 as=0 ps=0 w=19.11 l=0.22
R0 VCC.n717 VCC.n39 357.074
R1 VCC.n715 VCC.n43 357.074
R2 VCC.n346 VCC.n172 357.074
R3 VCC.n344 VCC.n174 357.074
R4 VCC.n579 VCC.t16 269.856
R5 VCC.n646 VCC.t5 269.856
R6 VCC.n196 VCC.t13 269.856
R7 VCC.n177 VCC.t9 269.856
R8 VCC.n715 VCC.n714 185
R9 VCC.n716 VCC.n715 185
R10 VCC.n44 VCC.n42 185
R11 VCC.n42 VCC.n40 185
R12 VCC.n541 VCC.n540 185
R13 VCC.n540 VCC.n539 185
R14 VCC.n47 VCC.n46 185
R15 VCC.n537 VCC.n47 185
R16 VCC.n535 VCC.n534 185
R17 VCC.n536 VCC.n535 185
R18 VCC.n49 VCC.n48 185
R19 VCC.n526 VCC.n48 185
R20 VCC.n530 VCC.n529 185
R21 VCC.n529 VCC.n528 185
R22 VCC.n52 VCC.n51 185
R23 VCC.n525 VCC.n52 185
R24 VCC.n523 VCC.n522 185
R25 VCC.n524 VCC.n523 185
R26 VCC.n55 VCC.n54 185
R27 VCC.n54 VCC.n53 185
R28 VCC.n518 VCC.n517 185
R29 VCC.n517 VCC.n516 185
R30 VCC.n58 VCC.n57 185
R31 VCC.n514 VCC.n58 185
R32 VCC.n512 VCC.n511 185
R33 VCC.n513 VCC.n512 185
R34 VCC.n61 VCC.n60 185
R35 VCC.n60 VCC.n59 185
R36 VCC.n507 VCC.n506 185
R37 VCC.n506 VCC.n505 185
R38 VCC.n64 VCC.n63 185
R39 VCC.n503 VCC.n64 185
R40 VCC.n501 VCC.n500 185
R41 VCC.n502 VCC.n501 185
R42 VCC.n67 VCC.n66 185
R43 VCC.n66 VCC.n65 185
R44 VCC.n496 VCC.n495 185
R45 VCC.n495 VCC.n494 185
R46 VCC.n70 VCC.n69 185
R47 VCC.n492 VCC.n70 185
R48 VCC.n490 VCC.n489 185
R49 VCC.n491 VCC.n490 185
R50 VCC.n73 VCC.n72 185
R51 VCC.n72 VCC.n71 185
R52 VCC.n485 VCC.n484 185
R53 VCC.n484 VCC.n483 185
R54 VCC.n76 VCC.n75 185
R55 VCC.n481 VCC.n76 185
R56 VCC.n479 VCC.n478 185
R57 VCC.n480 VCC.n479 185
R58 VCC.n79 VCC.n78 185
R59 VCC.n78 VCC.n77 185
R60 VCC.n474 VCC.n473 185
R61 VCC.n473 VCC.n472 185
R62 VCC.n82 VCC.n81 185
R63 VCC.n470 VCC.n82 185
R64 VCC.n468 VCC.n467 185
R65 VCC.n469 VCC.n468 185
R66 VCC.n85 VCC.n84 185
R67 VCC.n84 VCC.n83 185
R68 VCC.n463 VCC.n462 185
R69 VCC.n462 VCC.n461 185
R70 VCC.n88 VCC.n87 185
R71 VCC.n89 VCC.n88 185
R72 VCC.n450 VCC.n449 185
R73 VCC.n451 VCC.n450 185
R74 VCC.n97 VCC.n96 185
R75 VCC.n452 VCC.n96 185
R76 VCC.n445 VCC.n444 185
R77 VCC.n444 VCC.n95 185
R78 VCC.n443 VCC.n99 185
R79 VCC.n443 VCC.n442 185
R80 VCC.n109 VCC.n100 185
R81 VCC.n101 VCC.n100 185
R82 VCC.n433 VCC.n432 185
R83 VCC.n434 VCC.n433 185
R84 VCC.n108 VCC.n107 185
R85 VCC.n114 VCC.n107 185
R86 VCC.n427 VCC.n426 185
R87 VCC.n426 VCC.n425 185
R88 VCC.n112 VCC.n111 185
R89 VCC.n113 VCC.n112 185
R90 VCC.n416 VCC.n415 185
R91 VCC.n417 VCC.n416 185
R92 VCC.n122 VCC.n121 185
R93 VCC.n121 VCC.n120 185
R94 VCC.n411 VCC.n410 185
R95 VCC.n410 VCC.n409 185
R96 VCC.n125 VCC.n124 185
R97 VCC.n126 VCC.n125 185
R98 VCC.n400 VCC.n399 185
R99 VCC.n401 VCC.n400 185
R100 VCC.n134 VCC.n133 185
R101 VCC.n133 VCC.n132 185
R102 VCC.n395 VCC.n394 185
R103 VCC.n394 VCC.n393 185
R104 VCC.n137 VCC.n136 185
R105 VCC.n138 VCC.n137 185
R106 VCC.n384 VCC.n383 185
R107 VCC.n385 VCC.n384 185
R108 VCC.n146 VCC.n145 185
R109 VCC.n145 VCC.n144 185
R110 VCC.n379 VCC.n378 185
R111 VCC.n378 VCC.n377 185
R112 VCC.n149 VCC.n148 185
R113 VCC.n150 VCC.n149 185
R114 VCC.n368 VCC.n367 185
R115 VCC.n369 VCC.n368 185
R116 VCC.n158 VCC.n157 185
R117 VCC.n157 VCC.n156 185
R118 VCC.n363 VCC.n362 185
R119 VCC.n362 VCC.n361 185
R120 VCC.n161 VCC.n160 185
R121 VCC.n162 VCC.n161 185
R122 VCC.n352 VCC.n351 185
R123 VCC.n353 VCC.n352 185
R124 VCC.n170 VCC.n169 185
R125 VCC.n169 VCC.n168 185
R126 VCC.n347 VCC.n346 185
R127 VCC.n346 VCC.n345 185
R128 VCC.n344 VCC.n343 185
R129 VCC.n345 VCC.n344 185
R130 VCC.n167 VCC.n166 185
R131 VCC.n168 VCC.n167 185
R132 VCC.n355 VCC.n354 185
R133 VCC.n354 VCC.n353 185
R134 VCC.n164 VCC.n163 185
R135 VCC.n163 VCC.n162 185
R136 VCC.n360 VCC.n359 185
R137 VCC.n361 VCC.n360 185
R138 VCC.n155 VCC.n154 185
R139 VCC.n156 VCC.n155 185
R140 VCC.n371 VCC.n370 185
R141 VCC.n370 VCC.n369 185
R142 VCC.n152 VCC.n151 185
R143 VCC.n151 VCC.n150 185
R144 VCC.n376 VCC.n375 185
R145 VCC.n377 VCC.n376 185
R146 VCC.n143 VCC.n142 185
R147 VCC.n144 VCC.n143 185
R148 VCC.n387 VCC.n386 185
R149 VCC.n386 VCC.n385 185
R150 VCC.n140 VCC.n139 185
R151 VCC.n139 VCC.n138 185
R152 VCC.n392 VCC.n391 185
R153 VCC.n393 VCC.n392 185
R154 VCC.n131 VCC.n130 185
R155 VCC.n132 VCC.n131 185
R156 VCC.n403 VCC.n402 185
R157 VCC.n402 VCC.n401 185
R158 VCC.n128 VCC.n127 185
R159 VCC.n127 VCC.n126 185
R160 VCC.n408 VCC.n407 185
R161 VCC.n409 VCC.n408 185
R162 VCC.n119 VCC.n118 185
R163 VCC.n120 VCC.n119 185
R164 VCC.n419 VCC.n418 185
R165 VCC.n418 VCC.n417 185
R166 VCC.n116 VCC.n115 185
R167 VCC.n115 VCC.n113 185
R168 VCC.n424 VCC.n423 185
R169 VCC.n425 VCC.n424 185
R170 VCC.n106 VCC.n105 185
R171 VCC.n114 VCC.n106 185
R172 VCC.n436 VCC.n435 185
R173 VCC.n435 VCC.n434 185
R174 VCC.n103 VCC.n102 185
R175 VCC.n102 VCC.n101 185
R176 VCC.n441 VCC.n440 185
R177 VCC.n442 VCC.n441 185
R178 VCC.n94 VCC.n93 185
R179 VCC.n95 VCC.n94 185
R180 VCC.n454 VCC.n453 185
R181 VCC.n453 VCC.n452 185
R182 VCC.n91 VCC.n90 185
R183 VCC.n451 VCC.n90 185
R184 VCC.n459 VCC.n458 185
R185 VCC.n459 VCC.n89 185
R186 VCC.n460 VCC.n2 185
R187 VCC.n461 VCC.n460 185
R188 VCC.n761 VCC.n3 185
R189 VCC.n83 VCC.n3 185
R190 VCC.n760 VCC.n4 185
R191 VCC.n469 VCC.n4 185
R192 VCC.n759 VCC.n5 185
R193 VCC.n470 VCC.n5 185
R194 VCC.n471 VCC.n6 185
R195 VCC.n472 VCC.n471 185
R196 VCC.n755 VCC.n8 185
R197 VCC.n77 VCC.n8 185
R198 VCC.n754 VCC.n9 185
R199 VCC.n480 VCC.n9 185
R200 VCC.n753 VCC.n10 185
R201 VCC.n481 VCC.n10 185
R202 VCC.n482 VCC.n11 185
R203 VCC.n483 VCC.n482 185
R204 VCC.n749 VCC.n13 185
R205 VCC.n71 VCC.n13 185
R206 VCC.n748 VCC.n14 185
R207 VCC.n491 VCC.n14 185
R208 VCC.n747 VCC.n15 185
R209 VCC.n492 VCC.n15 185
R210 VCC.n493 VCC.n16 185
R211 VCC.n494 VCC.n493 185
R212 VCC.n743 VCC.n18 185
R213 VCC.n65 VCC.n18 185
R214 VCC.n742 VCC.n19 185
R215 VCC.n502 VCC.n19 185
R216 VCC.n741 VCC.n20 185
R217 VCC.n503 VCC.n20 185
R218 VCC.n504 VCC.n21 185
R219 VCC.n505 VCC.n504 185
R220 VCC.n737 VCC.n23 185
R221 VCC.n59 VCC.n23 185
R222 VCC.n736 VCC.n24 185
R223 VCC.n513 VCC.n24 185
R224 VCC.n735 VCC.n25 185
R225 VCC.n514 VCC.n25 185
R226 VCC.n515 VCC.n26 185
R227 VCC.n516 VCC.n515 185
R228 VCC.n731 VCC.n28 185
R229 VCC.n53 VCC.n28 185
R230 VCC.n730 VCC.n29 185
R231 VCC.n524 VCC.n29 185
R232 VCC.n729 VCC.n30 185
R233 VCC.n525 VCC.n30 185
R234 VCC.n527 VCC.n31 185
R235 VCC.n528 VCC.n527 185
R236 VCC.n725 VCC.n33 185
R237 VCC.n526 VCC.n33 185
R238 VCC.n724 VCC.n34 185
R239 VCC.n536 VCC.n34 185
R240 VCC.n723 VCC.n35 185
R241 VCC.n537 VCC.n35 185
R242 VCC.n538 VCC.n36 185
R243 VCC.n539 VCC.n538 185
R244 VCC.n719 VCC.n38 185
R245 VCC.n40 VCC.n38 185
R246 VCC.n718 VCC.n717 185
R247 VCC.n717 VCC.n716 185
R248 VCC.n712 VCC.n43 185
R249 VCC.n711 VCC.n710 185
R250 VCC.n708 VCC.n544 185
R251 VCC.n706 VCC.n705 185
R252 VCC.n704 VCC.n545 185
R253 VCC.n703 VCC.n702 185
R254 VCC.n700 VCC.n546 185
R255 VCC.n698 VCC.n697 185
R256 VCC.n696 VCC.n547 185
R257 VCC.n695 VCC.n694 185
R258 VCC.n692 VCC.n548 185
R259 VCC.n690 VCC.n689 185
R260 VCC.n688 VCC.n549 185
R261 VCC.n687 VCC.n686 185
R262 VCC.n684 VCC.n550 185
R263 VCC.n682 VCC.n681 185
R264 VCC.n680 VCC.n551 185
R265 VCC.n679 VCC.n678 185
R266 VCC.n676 VCC.n552 185
R267 VCC.n674 VCC.n673 185
R268 VCC.n672 VCC.n553 185
R269 VCC.n671 VCC.n670 185
R270 VCC.n668 VCC.n554 185
R271 VCC.n666 VCC.n665 185
R272 VCC.n664 VCC.n555 185
R273 VCC.n663 VCC.n662 185
R274 VCC.n660 VCC.n556 185
R275 VCC.n658 VCC.n657 185
R276 VCC.n656 VCC.n557 185
R277 VCC.n655 VCC.n654 185
R278 VCC.n652 VCC.n558 185
R279 VCC.n650 VCC.n649 185
R280 VCC.n645 VCC.n559 185
R281 VCC.n644 VCC.n643 185
R282 VCC.n641 VCC.n560 185
R283 VCC.n639 VCC.n638 185
R284 VCC.n637 VCC.n561 185
R285 VCC.n636 VCC.n635 185
R286 VCC.n633 VCC.n562 185
R287 VCC.n631 VCC.n630 185
R288 VCC.n629 VCC.n563 185
R289 VCC.n628 VCC.n627 185
R290 VCC.n625 VCC.n564 185
R291 VCC.n623 VCC.n622 185
R292 VCC.n621 VCC.n565 185
R293 VCC.n620 VCC.n619 185
R294 VCC.n617 VCC.n566 185
R295 VCC.n615 VCC.n614 185
R296 VCC.n613 VCC.n567 185
R297 VCC.n612 VCC.n611 185
R298 VCC.n609 VCC.n568 185
R299 VCC.n607 VCC.n606 185
R300 VCC.n605 VCC.n569 185
R301 VCC.n604 VCC.n603 185
R302 VCC.n601 VCC.n570 185
R303 VCC.n599 VCC.n598 185
R304 VCC.n597 VCC.n571 185
R305 VCC.n596 VCC.n595 185
R306 VCC.n593 VCC.n572 185
R307 VCC.n591 VCC.n590 185
R308 VCC.n589 VCC.n573 185
R309 VCC.n588 VCC.n587 185
R310 VCC.n585 VCC.n574 185
R311 VCC.n583 VCC.n582 185
R312 VCC.n578 VCC.n576 185
R313 VCC.n577 VCC.n39 185
R314 VCC.n341 VCC.n174 185
R315 VCC.n340 VCC.n339 185
R316 VCC.n337 VCC.n175 185
R317 VCC.n337 VCC.n173 185
R318 VCC.n336 VCC.n335 185
R319 VCC.n334 VCC.n333 185
R320 VCC.n332 VCC.n180 185
R321 VCC.n330 VCC.n329 185
R322 VCC.n328 VCC.n181 185
R323 VCC.n327 VCC.n326 185
R324 VCC.n324 VCC.n182 185
R325 VCC.n322 VCC.n321 185
R326 VCC.n320 VCC.n183 185
R327 VCC.n319 VCC.n318 185
R328 VCC.n316 VCC.n184 185
R329 VCC.n314 VCC.n313 185
R330 VCC.n312 VCC.n185 185
R331 VCC.n311 VCC.n310 185
R332 VCC.n308 VCC.n186 185
R333 VCC.n306 VCC.n305 185
R334 VCC.n304 VCC.n187 185
R335 VCC.n303 VCC.n302 185
R336 VCC.n300 VCC.n188 185
R337 VCC.n298 VCC.n297 185
R338 VCC.n296 VCC.n189 185
R339 VCC.n295 VCC.n294 185
R340 VCC.n292 VCC.n190 185
R341 VCC.n290 VCC.n289 185
R342 VCC.n288 VCC.n191 185
R343 VCC.n287 VCC.n286 185
R344 VCC.n284 VCC.n192 185
R345 VCC.n282 VCC.n281 185
R346 VCC.n280 VCC.n193 185
R347 VCC.n279 VCC.n278 185
R348 VCC.n276 VCC.n194 185
R349 VCC.n274 VCC.n273 185
R350 VCC.n271 VCC.n195 185
R351 VCC.n270 VCC.n269 185
R352 VCC.n267 VCC.n198 185
R353 VCC.n265 VCC.n264 185
R354 VCC.n263 VCC.n199 185
R355 VCC.n262 VCC.n261 185
R356 VCC.n259 VCC.n200 185
R357 VCC.n257 VCC.n256 185
R358 VCC.n255 VCC.n201 185
R359 VCC.n254 VCC.n253 185
R360 VCC.n251 VCC.n202 185
R361 VCC.n249 VCC.n248 185
R362 VCC.n247 VCC.n203 185
R363 VCC.n246 VCC.n245 185
R364 VCC.n243 VCC.n204 185
R365 VCC.n241 VCC.n240 185
R366 VCC.n239 VCC.n205 185
R367 VCC.n238 VCC.n237 185
R368 VCC.n235 VCC.n206 185
R369 VCC.n233 VCC.n232 185
R370 VCC.n231 VCC.n207 185
R371 VCC.n230 VCC.n229 185
R372 VCC.n227 VCC.n208 185
R373 VCC.n225 VCC.n224 185
R374 VCC.n223 VCC.n209 185
R375 VCC.n222 VCC.n221 185
R376 VCC.n219 VCC.n210 185
R377 VCC.n217 VCC.n216 185
R378 VCC.n215 VCC.n211 185
R379 VCC.n214 VCC.n213 185
R380 VCC.n172 VCC.n171 185
R381 VCC.n173 VCC.n172 185
R382 VCC.n579 VCC.t17 184.732
R383 VCC.n646 VCC.t7 184.732
R384 VCC.n196 VCC.t15 184.732
R385 VCC.n177 VCC.t12 184.732
R386 VCC.n346 VCC.n169 146.341
R387 VCC.n352 VCC.n169 146.341
R388 VCC.n352 VCC.n161 146.341
R389 VCC.n362 VCC.n161 146.341
R390 VCC.n362 VCC.n157 146.341
R391 VCC.n368 VCC.n157 146.341
R392 VCC.n368 VCC.n149 146.341
R393 VCC.n378 VCC.n149 146.341
R394 VCC.n378 VCC.n145 146.341
R395 VCC.n384 VCC.n145 146.341
R396 VCC.n384 VCC.n137 146.341
R397 VCC.n394 VCC.n137 146.341
R398 VCC.n394 VCC.n133 146.341
R399 VCC.n400 VCC.n133 146.341
R400 VCC.n400 VCC.n125 146.341
R401 VCC.n410 VCC.n125 146.341
R402 VCC.n410 VCC.n121 146.341
R403 VCC.n416 VCC.n121 146.341
R404 VCC.n416 VCC.n112 146.341
R405 VCC.n426 VCC.n112 146.341
R406 VCC.n426 VCC.n107 146.341
R407 VCC.n433 VCC.n107 146.341
R408 VCC.n433 VCC.n100 146.341
R409 VCC.n443 VCC.n100 146.341
R410 VCC.n444 VCC.n443 146.341
R411 VCC.n444 VCC.n96 146.341
R412 VCC.n450 VCC.n96 146.341
R413 VCC.n450 VCC.n88 146.341
R414 VCC.n462 VCC.n88 146.341
R415 VCC.n462 VCC.n84 146.341
R416 VCC.n468 VCC.n84 146.341
R417 VCC.n468 VCC.n82 146.341
R418 VCC.n473 VCC.n82 146.341
R419 VCC.n473 VCC.n78 146.341
R420 VCC.n479 VCC.n78 146.341
R421 VCC.n479 VCC.n76 146.341
R422 VCC.n484 VCC.n76 146.341
R423 VCC.n484 VCC.n72 146.341
R424 VCC.n490 VCC.n72 146.341
R425 VCC.n490 VCC.n70 146.341
R426 VCC.n495 VCC.n70 146.341
R427 VCC.n495 VCC.n66 146.341
R428 VCC.n501 VCC.n66 146.341
R429 VCC.n501 VCC.n64 146.341
R430 VCC.n506 VCC.n64 146.341
R431 VCC.n506 VCC.n60 146.341
R432 VCC.n512 VCC.n60 146.341
R433 VCC.n512 VCC.n58 146.341
R434 VCC.n517 VCC.n58 146.341
R435 VCC.n517 VCC.n54 146.341
R436 VCC.n523 VCC.n54 146.341
R437 VCC.n523 VCC.n52 146.341
R438 VCC.n529 VCC.n52 146.341
R439 VCC.n529 VCC.n48 146.341
R440 VCC.n535 VCC.n48 146.341
R441 VCC.n535 VCC.n47 146.341
R442 VCC.n540 VCC.n47 146.341
R443 VCC.n540 VCC.n42 146.341
R444 VCC.n715 VCC.n42 146.341
R445 VCC.n344 VCC.n167 146.341
R446 VCC.n354 VCC.n167 146.341
R447 VCC.n354 VCC.n163 146.341
R448 VCC.n360 VCC.n163 146.341
R449 VCC.n360 VCC.n155 146.341
R450 VCC.n370 VCC.n155 146.341
R451 VCC.n370 VCC.n151 146.341
R452 VCC.n376 VCC.n151 146.341
R453 VCC.n376 VCC.n143 146.341
R454 VCC.n386 VCC.n143 146.341
R455 VCC.n386 VCC.n139 146.341
R456 VCC.n392 VCC.n139 146.341
R457 VCC.n392 VCC.n131 146.341
R458 VCC.n402 VCC.n131 146.341
R459 VCC.n402 VCC.n127 146.341
R460 VCC.n408 VCC.n127 146.341
R461 VCC.n408 VCC.n119 146.341
R462 VCC.n418 VCC.n119 146.341
R463 VCC.n418 VCC.n115 146.341
R464 VCC.n424 VCC.n115 146.341
R465 VCC.n424 VCC.n106 146.341
R466 VCC.n435 VCC.n106 146.341
R467 VCC.n435 VCC.n102 146.341
R468 VCC.n441 VCC.n102 146.341
R469 VCC.n441 VCC.n94 146.341
R470 VCC.n453 VCC.n94 146.341
R471 VCC.n453 VCC.n90 146.341
R472 VCC.n459 VCC.n90 146.341
R473 VCC.n460 VCC.n459 146.341
R474 VCC.n460 VCC.n3 146.341
R475 VCC.n4 VCC.n3 146.341
R476 VCC.n5 VCC.n4 146.341
R477 VCC.n471 VCC.n5 146.341
R478 VCC.n471 VCC.n8 146.341
R479 VCC.n9 VCC.n8 146.341
R480 VCC.n10 VCC.n9 146.341
R481 VCC.n482 VCC.n10 146.341
R482 VCC.n482 VCC.n13 146.341
R483 VCC.n14 VCC.n13 146.341
R484 VCC.n15 VCC.n14 146.341
R485 VCC.n493 VCC.n15 146.341
R486 VCC.n493 VCC.n18 146.341
R487 VCC.n19 VCC.n18 146.341
R488 VCC.n20 VCC.n19 146.341
R489 VCC.n504 VCC.n20 146.341
R490 VCC.n504 VCC.n23 146.341
R491 VCC.n24 VCC.n23 146.341
R492 VCC.n25 VCC.n24 146.341
R493 VCC.n515 VCC.n25 146.341
R494 VCC.n515 VCC.n28 146.341
R495 VCC.n29 VCC.n28 146.341
R496 VCC.n30 VCC.n29 146.341
R497 VCC.n527 VCC.n30 146.341
R498 VCC.n527 VCC.n33 146.341
R499 VCC.n34 VCC.n33 146.341
R500 VCC.n35 VCC.n34 146.341
R501 VCC.n538 VCC.n35 146.341
R502 VCC.n538 VCC.n38 146.341
R503 VCC.n717 VCC.n38 146.341
R504 VCC.n580 VCC.t18 109.678
R505 VCC.n647 VCC.t8 109.678
R506 VCC.n197 VCC.t14 109.678
R507 VCC.n178 VCC.t11 109.678
R508 VCC.n583 VCC.n576 99.5127
R509 VCC.n587 VCC.n585 99.5127
R510 VCC.n591 VCC.n573 99.5127
R511 VCC.n595 VCC.n593 99.5127
R512 VCC.n599 VCC.n571 99.5127
R513 VCC.n603 VCC.n601 99.5127
R514 VCC.n607 VCC.n569 99.5127
R515 VCC.n611 VCC.n609 99.5127
R516 VCC.n615 VCC.n567 99.5127
R517 VCC.n619 VCC.n617 99.5127
R518 VCC.n623 VCC.n565 99.5127
R519 VCC.n627 VCC.n625 99.5127
R520 VCC.n631 VCC.n563 99.5127
R521 VCC.n635 VCC.n633 99.5127
R522 VCC.n639 VCC.n561 99.5127
R523 VCC.n643 VCC.n641 99.5127
R524 VCC.n650 VCC.n559 99.5127
R525 VCC.n654 VCC.n652 99.5127
R526 VCC.n658 VCC.n557 99.5127
R527 VCC.n662 VCC.n660 99.5127
R528 VCC.n666 VCC.n555 99.5127
R529 VCC.n670 VCC.n668 99.5127
R530 VCC.n674 VCC.n553 99.5127
R531 VCC.n678 VCC.n676 99.5127
R532 VCC.n682 VCC.n551 99.5127
R533 VCC.n686 VCC.n684 99.5127
R534 VCC.n690 VCC.n549 99.5127
R535 VCC.n694 VCC.n692 99.5127
R536 VCC.n698 VCC.n547 99.5127
R537 VCC.n702 VCC.n700 99.5127
R538 VCC.n706 VCC.n545 99.5127
R539 VCC.n710 VCC.n708 99.5127
R540 VCC.n339 VCC.n337 99.5127
R541 VCC.n337 VCC.n336 99.5127
R542 VCC.n333 VCC.n332 99.5127
R543 VCC.n330 VCC.n181 99.5127
R544 VCC.n326 VCC.n324 99.5127
R545 VCC.n322 VCC.n183 99.5127
R546 VCC.n318 VCC.n316 99.5127
R547 VCC.n314 VCC.n185 99.5127
R548 VCC.n310 VCC.n308 99.5127
R549 VCC.n306 VCC.n187 99.5127
R550 VCC.n302 VCC.n300 99.5127
R551 VCC.n298 VCC.n189 99.5127
R552 VCC.n294 VCC.n292 99.5127
R553 VCC.n290 VCC.n191 99.5127
R554 VCC.n286 VCC.n284 99.5127
R555 VCC.n282 VCC.n193 99.5127
R556 VCC.n278 VCC.n276 99.5127
R557 VCC.n274 VCC.n195 99.5127
R558 VCC.n269 VCC.n267 99.5127
R559 VCC.n265 VCC.n199 99.5127
R560 VCC.n261 VCC.n259 99.5127
R561 VCC.n257 VCC.n201 99.5127
R562 VCC.n253 VCC.n251 99.5127
R563 VCC.n249 VCC.n203 99.5127
R564 VCC.n245 VCC.n243 99.5127
R565 VCC.n241 VCC.n205 99.5127
R566 VCC.n237 VCC.n235 99.5127
R567 VCC.n233 VCC.n207 99.5127
R568 VCC.n229 VCC.n227 99.5127
R569 VCC.n225 VCC.n209 99.5127
R570 VCC.n221 VCC.n219 99.5127
R571 VCC.n217 VCC.n211 99.5127
R572 VCC.n213 VCC.n172 99.5127
R573 VCC.n580 VCC.n579 75.0551
R574 VCC.n647 VCC.n646 75.0551
R575 VCC.n197 VCC.n196 75.0551
R576 VCC.n178 VCC.n177 75.0551
R577 VCC.n709 VCC.n41 72.8958
R578 VCC.n707 VCC.n41 72.8958
R579 VCC.n701 VCC.n41 72.8958
R580 VCC.n699 VCC.n41 72.8958
R581 VCC.n693 VCC.n41 72.8958
R582 VCC.n691 VCC.n41 72.8958
R583 VCC.n685 VCC.n41 72.8958
R584 VCC.n683 VCC.n41 72.8958
R585 VCC.n677 VCC.n41 72.8958
R586 VCC.n675 VCC.n41 72.8958
R587 VCC.n669 VCC.n41 72.8958
R588 VCC.n667 VCC.n41 72.8958
R589 VCC.n661 VCC.n41 72.8958
R590 VCC.n659 VCC.n41 72.8958
R591 VCC.n653 VCC.n41 72.8958
R592 VCC.n651 VCC.n41 72.8958
R593 VCC.n642 VCC.n41 72.8958
R594 VCC.n640 VCC.n41 72.8958
R595 VCC.n634 VCC.n41 72.8958
R596 VCC.n632 VCC.n41 72.8958
R597 VCC.n626 VCC.n41 72.8958
R598 VCC.n624 VCC.n41 72.8958
R599 VCC.n618 VCC.n41 72.8958
R600 VCC.n616 VCC.n41 72.8958
R601 VCC.n610 VCC.n41 72.8958
R602 VCC.n608 VCC.n41 72.8958
R603 VCC.n602 VCC.n41 72.8958
R604 VCC.n600 VCC.n41 72.8958
R605 VCC.n594 VCC.n41 72.8958
R606 VCC.n592 VCC.n41 72.8958
R607 VCC.n586 VCC.n41 72.8958
R608 VCC.n584 VCC.n41 72.8958
R609 VCC.n575 VCC.n41 72.8958
R610 VCC.n338 VCC.n173 72.8958
R611 VCC.n176 VCC.n173 72.8958
R612 VCC.n331 VCC.n173 72.8958
R613 VCC.n325 VCC.n173 72.8958
R614 VCC.n323 VCC.n173 72.8958
R615 VCC.n317 VCC.n173 72.8958
R616 VCC.n315 VCC.n173 72.8958
R617 VCC.n309 VCC.n173 72.8958
R618 VCC.n307 VCC.n173 72.8958
R619 VCC.n301 VCC.n173 72.8958
R620 VCC.n299 VCC.n173 72.8958
R621 VCC.n293 VCC.n173 72.8958
R622 VCC.n291 VCC.n173 72.8958
R623 VCC.n285 VCC.n173 72.8958
R624 VCC.n283 VCC.n173 72.8958
R625 VCC.n277 VCC.n173 72.8958
R626 VCC.n275 VCC.n173 72.8958
R627 VCC.n268 VCC.n173 72.8958
R628 VCC.n266 VCC.n173 72.8958
R629 VCC.n260 VCC.n173 72.8958
R630 VCC.n258 VCC.n173 72.8958
R631 VCC.n252 VCC.n173 72.8958
R632 VCC.n250 VCC.n173 72.8958
R633 VCC.n244 VCC.n173 72.8958
R634 VCC.n242 VCC.n173 72.8958
R635 VCC.n236 VCC.n173 72.8958
R636 VCC.n234 VCC.n173 72.8958
R637 VCC.n228 VCC.n173 72.8958
R638 VCC.n226 VCC.n173 72.8958
R639 VCC.n220 VCC.n173 72.8958
R640 VCC.n218 VCC.n173 72.8958
R641 VCC.n212 VCC.n173 72.8958
R642 VCC.n576 VCC.n575 39.2114
R643 VCC.n585 VCC.n584 39.2114
R644 VCC.n586 VCC.n573 39.2114
R645 VCC.n593 VCC.n592 39.2114
R646 VCC.n594 VCC.n571 39.2114
R647 VCC.n601 VCC.n600 39.2114
R648 VCC.n602 VCC.n569 39.2114
R649 VCC.n609 VCC.n608 39.2114
R650 VCC.n610 VCC.n567 39.2114
R651 VCC.n617 VCC.n616 39.2114
R652 VCC.n618 VCC.n565 39.2114
R653 VCC.n625 VCC.n624 39.2114
R654 VCC.n626 VCC.n563 39.2114
R655 VCC.n633 VCC.n632 39.2114
R656 VCC.n634 VCC.n561 39.2114
R657 VCC.n641 VCC.n640 39.2114
R658 VCC.n642 VCC.n559 39.2114
R659 VCC.n652 VCC.n651 39.2114
R660 VCC.n653 VCC.n557 39.2114
R661 VCC.n660 VCC.n659 39.2114
R662 VCC.n661 VCC.n555 39.2114
R663 VCC.n668 VCC.n667 39.2114
R664 VCC.n669 VCC.n553 39.2114
R665 VCC.n676 VCC.n675 39.2114
R666 VCC.n677 VCC.n551 39.2114
R667 VCC.n684 VCC.n683 39.2114
R668 VCC.n685 VCC.n549 39.2114
R669 VCC.n692 VCC.n691 39.2114
R670 VCC.n693 VCC.n547 39.2114
R671 VCC.n700 VCC.n699 39.2114
R672 VCC.n701 VCC.n545 39.2114
R673 VCC.n708 VCC.n707 39.2114
R674 VCC.n709 VCC.n43 39.2114
R675 VCC.n338 VCC.n174 39.2114
R676 VCC.n336 VCC.n176 39.2114
R677 VCC.n332 VCC.n331 39.2114
R678 VCC.n325 VCC.n181 39.2114
R679 VCC.n324 VCC.n323 39.2114
R680 VCC.n317 VCC.n183 39.2114
R681 VCC.n316 VCC.n315 39.2114
R682 VCC.n309 VCC.n185 39.2114
R683 VCC.n308 VCC.n307 39.2114
R684 VCC.n301 VCC.n187 39.2114
R685 VCC.n300 VCC.n299 39.2114
R686 VCC.n293 VCC.n189 39.2114
R687 VCC.n292 VCC.n291 39.2114
R688 VCC.n285 VCC.n191 39.2114
R689 VCC.n284 VCC.n283 39.2114
R690 VCC.n277 VCC.n193 39.2114
R691 VCC.n276 VCC.n275 39.2114
R692 VCC.n268 VCC.n195 39.2114
R693 VCC.n267 VCC.n266 39.2114
R694 VCC.n260 VCC.n199 39.2114
R695 VCC.n259 VCC.n258 39.2114
R696 VCC.n252 VCC.n201 39.2114
R697 VCC.n251 VCC.n250 39.2114
R698 VCC.n244 VCC.n203 39.2114
R699 VCC.n243 VCC.n242 39.2114
R700 VCC.n236 VCC.n205 39.2114
R701 VCC.n235 VCC.n234 39.2114
R702 VCC.n228 VCC.n207 39.2114
R703 VCC.n227 VCC.n226 39.2114
R704 VCC.n220 VCC.n209 39.2114
R705 VCC.n219 VCC.n218 39.2114
R706 VCC.n212 VCC.n211 39.2114
R707 VCC.n710 VCC.n709 39.2114
R708 VCC.n707 VCC.n706 39.2114
R709 VCC.n702 VCC.n701 39.2114
R710 VCC.n699 VCC.n698 39.2114
R711 VCC.n694 VCC.n693 39.2114
R712 VCC.n691 VCC.n690 39.2114
R713 VCC.n686 VCC.n685 39.2114
R714 VCC.n683 VCC.n682 39.2114
R715 VCC.n678 VCC.n677 39.2114
R716 VCC.n675 VCC.n674 39.2114
R717 VCC.n670 VCC.n669 39.2114
R718 VCC.n667 VCC.n666 39.2114
R719 VCC.n662 VCC.n661 39.2114
R720 VCC.n659 VCC.n658 39.2114
R721 VCC.n654 VCC.n653 39.2114
R722 VCC.n651 VCC.n650 39.2114
R723 VCC.n643 VCC.n642 39.2114
R724 VCC.n640 VCC.n639 39.2114
R725 VCC.n635 VCC.n634 39.2114
R726 VCC.n632 VCC.n631 39.2114
R727 VCC.n627 VCC.n626 39.2114
R728 VCC.n624 VCC.n623 39.2114
R729 VCC.n619 VCC.n618 39.2114
R730 VCC.n616 VCC.n615 39.2114
R731 VCC.n611 VCC.n610 39.2114
R732 VCC.n608 VCC.n607 39.2114
R733 VCC.n603 VCC.n602 39.2114
R734 VCC.n600 VCC.n599 39.2114
R735 VCC.n595 VCC.n594 39.2114
R736 VCC.n592 VCC.n591 39.2114
R737 VCC.n587 VCC.n586 39.2114
R738 VCC.n584 VCC.n583 39.2114
R739 VCC.n575 VCC.n39 39.2114
R740 VCC.n339 VCC.n338 39.2114
R741 VCC.n333 VCC.n176 39.2114
R742 VCC.n331 VCC.n330 39.2114
R743 VCC.n326 VCC.n325 39.2114
R744 VCC.n323 VCC.n322 39.2114
R745 VCC.n318 VCC.n317 39.2114
R746 VCC.n315 VCC.n314 39.2114
R747 VCC.n310 VCC.n309 39.2114
R748 VCC.n307 VCC.n306 39.2114
R749 VCC.n302 VCC.n301 39.2114
R750 VCC.n299 VCC.n298 39.2114
R751 VCC.n294 VCC.n293 39.2114
R752 VCC.n291 VCC.n290 39.2114
R753 VCC.n286 VCC.n285 39.2114
R754 VCC.n283 VCC.n282 39.2114
R755 VCC.n278 VCC.n277 39.2114
R756 VCC.n275 VCC.n274 39.2114
R757 VCC.n269 VCC.n268 39.2114
R758 VCC.n266 VCC.n265 39.2114
R759 VCC.n261 VCC.n260 39.2114
R760 VCC.n258 VCC.n257 39.2114
R761 VCC.n253 VCC.n252 39.2114
R762 VCC.n250 VCC.n249 39.2114
R763 VCC.n245 VCC.n244 39.2114
R764 VCC.n242 VCC.n241 39.2114
R765 VCC.n237 VCC.n236 39.2114
R766 VCC.n234 VCC.n233 39.2114
R767 VCC.n229 VCC.n228 39.2114
R768 VCC.n226 VCC.n225 39.2114
R769 VCC.n221 VCC.n220 39.2114
R770 VCC.n218 VCC.n217 39.2114
R771 VCC.n213 VCC.n212 39.2114
R772 VCC.n345 VCC.n173 33.0491
R773 VCC.n716 VCC.n41 33.0491
R774 VCC.n581 VCC.n580 29.2853
R775 VCC.n648 VCC.n647 29.2853
R776 VCC.n272 VCC.n197 29.2853
R777 VCC.n179 VCC.n178 29.2853
R778 VCC.n577 VCC.n37 27.6654
R779 VCC.n713 VCC.n712 27.6654
R780 VCC.n342 VCC.n341 27.6654
R781 VCC.n348 VCC.n171 27.6654
R782 VCC.n345 VCC.n168 19.5559
R783 VCC.n353 VCC.n168 19.5559
R784 VCC.n353 VCC.n162 19.5559
R785 VCC.n361 VCC.n162 19.5559
R786 VCC.n369 VCC.n156 19.5559
R787 VCC.n369 VCC.n150 19.5559
R788 VCC.n377 VCC.n150 19.5559
R789 VCC.n377 VCC.n144 19.5559
R790 VCC.n385 VCC.n144 19.5559
R791 VCC.n385 VCC.n138 19.5559
R792 VCC.n393 VCC.n138 19.5559
R793 VCC.n393 VCC.n132 19.5559
R794 VCC.n401 VCC.n132 19.5559
R795 VCC.n409 VCC.n126 19.5559
R796 VCC.n409 VCC.n120 19.5559
R797 VCC.n417 VCC.n120 19.5559
R798 VCC.n417 VCC.n113 19.5559
R799 VCC.n425 VCC.n113 19.5559
R800 VCC.n425 VCC.n114 19.5559
R801 VCC.n434 VCC.n101 19.5559
R802 VCC.n442 VCC.n101 19.5559
R803 VCC.n442 VCC.n95 19.5559
R804 VCC.n452 VCC.n95 19.5559
R805 VCC.n452 VCC.n451 19.5559
R806 VCC.n451 VCC.n89 19.5559
R807 VCC.n461 VCC.n89 19.5559
R808 VCC.n469 VCC.n83 19.5559
R809 VCC.n470 VCC.n469 19.5559
R810 VCC.n472 VCC.n470 19.5559
R811 VCC.n472 VCC.n77 19.5559
R812 VCC.n480 VCC.n77 19.5559
R813 VCC.n481 VCC.n480 19.5559
R814 VCC.n483 VCC.n481 19.5559
R815 VCC.n491 VCC.n71 19.5559
R816 VCC.n492 VCC.n491 19.5559
R817 VCC.n494 VCC.n492 19.5559
R818 VCC.n494 VCC.n65 19.5559
R819 VCC.n502 VCC.n65 19.5559
R820 VCC.n503 VCC.n502 19.5559
R821 VCC.n505 VCC.n59 19.5559
R822 VCC.n513 VCC.n59 19.5559
R823 VCC.n514 VCC.n513 19.5559
R824 VCC.n516 VCC.n514 19.5559
R825 VCC.n516 VCC.n53 19.5559
R826 VCC.n524 VCC.n53 19.5559
R827 VCC.n525 VCC.n524 19.5559
R828 VCC.n528 VCC.n525 19.5559
R829 VCC.n528 VCC.n526 19.5559
R830 VCC.n537 VCC.n536 19.5559
R831 VCC.n539 VCC.n537 19.5559
R832 VCC.n539 VCC.n40 19.5559
R833 VCC.n716 VCC.n40 19.5559
R834 VCC.n347 VCC.n170 19.3944
R835 VCC.n351 VCC.n170 19.3944
R836 VCC.n351 VCC.n160 19.3944
R837 VCC.n363 VCC.n160 19.3944
R838 VCC.n363 VCC.n158 19.3944
R839 VCC.n367 VCC.n158 19.3944
R840 VCC.n367 VCC.n148 19.3944
R841 VCC.n379 VCC.n148 19.3944
R842 VCC.n379 VCC.n146 19.3944
R843 VCC.n383 VCC.n146 19.3944
R844 VCC.n383 VCC.n136 19.3944
R845 VCC.n395 VCC.n136 19.3944
R846 VCC.n395 VCC.n134 19.3944
R847 VCC.n399 VCC.n134 19.3944
R848 VCC.n399 VCC.n124 19.3944
R849 VCC.n411 VCC.n124 19.3944
R850 VCC.n411 VCC.n122 19.3944
R851 VCC.n415 VCC.n122 19.3944
R852 VCC.n415 VCC.n111 19.3944
R853 VCC.n427 VCC.n111 19.3944
R854 VCC.n427 VCC.n108 19.3944
R855 VCC.n432 VCC.n108 19.3944
R856 VCC.n432 VCC.n109 19.3944
R857 VCC.n109 VCC.n99 19.3944
R858 VCC.n445 VCC.n99 19.3944
R859 VCC.n445 VCC.n97 19.3944
R860 VCC.n449 VCC.n97 19.3944
R861 VCC.n449 VCC.n87 19.3944
R862 VCC.n463 VCC.n87 19.3944
R863 VCC.n463 VCC.n85 19.3944
R864 VCC.n467 VCC.n85 19.3944
R865 VCC.n467 VCC.n81 19.3944
R866 VCC.n474 VCC.n81 19.3944
R867 VCC.n474 VCC.n79 19.3944
R868 VCC.n478 VCC.n79 19.3944
R869 VCC.n478 VCC.n75 19.3944
R870 VCC.n485 VCC.n75 19.3944
R871 VCC.n485 VCC.n73 19.3944
R872 VCC.n489 VCC.n73 19.3944
R873 VCC.n489 VCC.n69 19.3944
R874 VCC.n496 VCC.n69 19.3944
R875 VCC.n496 VCC.n67 19.3944
R876 VCC.n500 VCC.n67 19.3944
R877 VCC.n500 VCC.n63 19.3944
R878 VCC.n507 VCC.n63 19.3944
R879 VCC.n507 VCC.n61 19.3944
R880 VCC.n511 VCC.n61 19.3944
R881 VCC.n511 VCC.n57 19.3944
R882 VCC.n518 VCC.n57 19.3944
R883 VCC.n518 VCC.n55 19.3944
R884 VCC.n522 VCC.n55 19.3944
R885 VCC.n522 VCC.n51 19.3944
R886 VCC.n530 VCC.n51 19.3944
R887 VCC.n530 VCC.n49 19.3944
R888 VCC.n534 VCC.n49 19.3944
R889 VCC.n534 VCC.n46 19.3944
R890 VCC.n541 VCC.n46 19.3944
R891 VCC.n541 VCC.n44 19.3944
R892 VCC.n714 VCC.n44 19.3944
R893 VCC.n343 VCC.n166 19.3944
R894 VCC.n355 VCC.n166 19.3944
R895 VCC.n355 VCC.n164 19.3944
R896 VCC.n359 VCC.n164 19.3944
R897 VCC.n359 VCC.n154 19.3944
R898 VCC.n371 VCC.n154 19.3944
R899 VCC.n371 VCC.n152 19.3944
R900 VCC.n375 VCC.n152 19.3944
R901 VCC.n375 VCC.n142 19.3944
R902 VCC.n387 VCC.n142 19.3944
R903 VCC.n387 VCC.n140 19.3944
R904 VCC.n391 VCC.n140 19.3944
R905 VCC.n391 VCC.n130 19.3944
R906 VCC.n403 VCC.n130 19.3944
R907 VCC.n403 VCC.n128 19.3944
R908 VCC.n407 VCC.n128 19.3944
R909 VCC.n407 VCC.n118 19.3944
R910 VCC.n419 VCC.n118 19.3944
R911 VCC.n419 VCC.n116 19.3944
R912 VCC.n423 VCC.n116 19.3944
R913 VCC.n423 VCC.n105 19.3944
R914 VCC.n436 VCC.n105 19.3944
R915 VCC.n436 VCC.n103 19.3944
R916 VCC.n440 VCC.n103 19.3944
R917 VCC.n440 VCC.n93 19.3944
R918 VCC.n454 VCC.n93 19.3944
R919 VCC.n454 VCC.n91 19.3944
R920 VCC.n458 VCC.n91 19.3944
R921 VCC.n458 VCC.n2 19.3944
R922 VCC.n761 VCC.n2 19.3944
R923 VCC.n761 VCC.n760 19.3944
R924 VCC.n760 VCC.n759 19.3944
R925 VCC.n759 VCC.n6 19.3944
R926 VCC.n755 VCC.n6 19.3944
R927 VCC.n755 VCC.n754 19.3944
R928 VCC.n754 VCC.n753 19.3944
R929 VCC.n753 VCC.n11 19.3944
R930 VCC.n749 VCC.n11 19.3944
R931 VCC.n749 VCC.n748 19.3944
R932 VCC.n748 VCC.n747 19.3944
R933 VCC.n747 VCC.n16 19.3944
R934 VCC.n743 VCC.n16 19.3944
R935 VCC.n743 VCC.n742 19.3944
R936 VCC.n742 VCC.n741 19.3944
R937 VCC.n741 VCC.n21 19.3944
R938 VCC.n737 VCC.n21 19.3944
R939 VCC.n737 VCC.n736 19.3944
R940 VCC.n736 VCC.n735 19.3944
R941 VCC.n735 VCC.n26 19.3944
R942 VCC.n731 VCC.n26 19.3944
R943 VCC.n731 VCC.n730 19.3944
R944 VCC.n730 VCC.n729 19.3944
R945 VCC.n729 VCC.n31 19.3944
R946 VCC.n725 VCC.n31 19.3944
R947 VCC.n725 VCC.n724 19.3944
R948 VCC.n724 VCC.n723 19.3944
R949 VCC.n723 VCC.n36 19.3944
R950 VCC.n719 VCC.n36 19.3944
R951 VCC.n719 VCC.n718 19.3944
R952 VCC.t4 VCC.n126 19.1648
R953 VCC.t3 VCC.n503 19.1648
R954 VCC.t10 VCC.n156 17.6003
R955 VCC.n526 VCC.t6 17.6003
R956 VCC.n114 VCC.t0 14.8626
R957 VCC.t1 VCC.n71 14.8626
R958 VCC.n578 VCC.n577 10.6151
R959 VCC.n582 VCC.n578 10.6151
R960 VCC.n588 VCC.n574 10.6151
R961 VCC.n589 VCC.n588 10.6151
R962 VCC.n590 VCC.n589 10.6151
R963 VCC.n590 VCC.n572 10.6151
R964 VCC.n596 VCC.n572 10.6151
R965 VCC.n597 VCC.n596 10.6151
R966 VCC.n598 VCC.n597 10.6151
R967 VCC.n598 VCC.n570 10.6151
R968 VCC.n604 VCC.n570 10.6151
R969 VCC.n605 VCC.n604 10.6151
R970 VCC.n606 VCC.n605 10.6151
R971 VCC.n606 VCC.n568 10.6151
R972 VCC.n612 VCC.n568 10.6151
R973 VCC.n613 VCC.n612 10.6151
R974 VCC.n614 VCC.n613 10.6151
R975 VCC.n614 VCC.n566 10.6151
R976 VCC.n620 VCC.n566 10.6151
R977 VCC.n621 VCC.n620 10.6151
R978 VCC.n622 VCC.n621 10.6151
R979 VCC.n622 VCC.n564 10.6151
R980 VCC.n628 VCC.n564 10.6151
R981 VCC.n629 VCC.n628 10.6151
R982 VCC.n630 VCC.n629 10.6151
R983 VCC.n630 VCC.n562 10.6151
R984 VCC.n636 VCC.n562 10.6151
R985 VCC.n637 VCC.n636 10.6151
R986 VCC.n638 VCC.n637 10.6151
R987 VCC.n638 VCC.n560 10.6151
R988 VCC.n644 VCC.n560 10.6151
R989 VCC.n645 VCC.n644 10.6151
R990 VCC.n649 VCC.n645 10.6151
R991 VCC.n655 VCC.n558 10.6151
R992 VCC.n656 VCC.n655 10.6151
R993 VCC.n657 VCC.n656 10.6151
R994 VCC.n657 VCC.n556 10.6151
R995 VCC.n663 VCC.n556 10.6151
R996 VCC.n664 VCC.n663 10.6151
R997 VCC.n665 VCC.n664 10.6151
R998 VCC.n665 VCC.n554 10.6151
R999 VCC.n671 VCC.n554 10.6151
R1000 VCC.n672 VCC.n671 10.6151
R1001 VCC.n673 VCC.n672 10.6151
R1002 VCC.n673 VCC.n552 10.6151
R1003 VCC.n679 VCC.n552 10.6151
R1004 VCC.n680 VCC.n679 10.6151
R1005 VCC.n681 VCC.n680 10.6151
R1006 VCC.n681 VCC.n550 10.6151
R1007 VCC.n687 VCC.n550 10.6151
R1008 VCC.n688 VCC.n687 10.6151
R1009 VCC.n689 VCC.n688 10.6151
R1010 VCC.n689 VCC.n548 10.6151
R1011 VCC.n695 VCC.n548 10.6151
R1012 VCC.n696 VCC.n695 10.6151
R1013 VCC.n697 VCC.n696 10.6151
R1014 VCC.n697 VCC.n546 10.6151
R1015 VCC.n703 VCC.n546 10.6151
R1016 VCC.n704 VCC.n703 10.6151
R1017 VCC.n705 VCC.n704 10.6151
R1018 VCC.n705 VCC.n544 10.6151
R1019 VCC.n711 VCC.n544 10.6151
R1020 VCC.n712 VCC.n711 10.6151
R1021 VCC.n341 VCC.n340 10.6151
R1022 VCC.n340 VCC.n175 10.6151
R1023 VCC.n335 VCC.n334 10.6151
R1024 VCC.n334 VCC.n180 10.6151
R1025 VCC.n329 VCC.n180 10.6151
R1026 VCC.n329 VCC.n328 10.6151
R1027 VCC.n328 VCC.n327 10.6151
R1028 VCC.n327 VCC.n182 10.6151
R1029 VCC.n321 VCC.n182 10.6151
R1030 VCC.n321 VCC.n320 10.6151
R1031 VCC.n320 VCC.n319 10.6151
R1032 VCC.n319 VCC.n184 10.6151
R1033 VCC.n313 VCC.n184 10.6151
R1034 VCC.n313 VCC.n312 10.6151
R1035 VCC.n312 VCC.n311 10.6151
R1036 VCC.n311 VCC.n186 10.6151
R1037 VCC.n305 VCC.n186 10.6151
R1038 VCC.n305 VCC.n304 10.6151
R1039 VCC.n304 VCC.n303 10.6151
R1040 VCC.n303 VCC.n188 10.6151
R1041 VCC.n297 VCC.n188 10.6151
R1042 VCC.n297 VCC.n296 10.6151
R1043 VCC.n296 VCC.n295 10.6151
R1044 VCC.n295 VCC.n190 10.6151
R1045 VCC.n289 VCC.n190 10.6151
R1046 VCC.n289 VCC.n288 10.6151
R1047 VCC.n288 VCC.n287 10.6151
R1048 VCC.n287 VCC.n192 10.6151
R1049 VCC.n281 VCC.n192 10.6151
R1050 VCC.n281 VCC.n280 10.6151
R1051 VCC.n280 VCC.n279 10.6151
R1052 VCC.n279 VCC.n194 10.6151
R1053 VCC.n273 VCC.n194 10.6151
R1054 VCC.n271 VCC.n270 10.6151
R1055 VCC.n270 VCC.n198 10.6151
R1056 VCC.n264 VCC.n198 10.6151
R1057 VCC.n264 VCC.n263 10.6151
R1058 VCC.n263 VCC.n262 10.6151
R1059 VCC.n262 VCC.n200 10.6151
R1060 VCC.n256 VCC.n200 10.6151
R1061 VCC.n256 VCC.n255 10.6151
R1062 VCC.n255 VCC.n254 10.6151
R1063 VCC.n254 VCC.n202 10.6151
R1064 VCC.n248 VCC.n202 10.6151
R1065 VCC.n248 VCC.n247 10.6151
R1066 VCC.n247 VCC.n246 10.6151
R1067 VCC.n246 VCC.n204 10.6151
R1068 VCC.n240 VCC.n204 10.6151
R1069 VCC.n240 VCC.n239 10.6151
R1070 VCC.n239 VCC.n238 10.6151
R1071 VCC.n238 VCC.n206 10.6151
R1072 VCC.n232 VCC.n206 10.6151
R1073 VCC.n232 VCC.n231 10.6151
R1074 VCC.n231 VCC.n230 10.6151
R1075 VCC.n230 VCC.n208 10.6151
R1076 VCC.n224 VCC.n208 10.6151
R1077 VCC.n224 VCC.n223 10.6151
R1078 VCC.n223 VCC.n222 10.6151
R1079 VCC.n222 VCC.n210 10.6151
R1080 VCC.n216 VCC.n210 10.6151
R1081 VCC.n216 VCC.n215 10.6151
R1082 VCC.n215 VCC.n214 10.6151
R1083 VCC.n214 VCC.n171 10.6151
R1084 VCC.n581 VCC.n574 10.1468
R1085 VCC.n335 VCC.n179 10.1468
R1086 VCC.n649 VCC.n648 9.83465
R1087 VCC.n273 VCC.n272 9.83465
R1088 VCC.n461 VCC.t2 9.77819
R1089 VCC.t2 VCC.n83 9.77819
R1090 VCC.n760 VCC.n0 9.3005
R1091 VCC.n759 VCC.n758 9.3005
R1092 VCC.n757 VCC.n6 9.3005
R1093 VCC.n756 VCC.n755 9.3005
R1094 VCC.n754 VCC.n7 9.3005
R1095 VCC.n753 VCC.n752 9.3005
R1096 VCC.n751 VCC.n11 9.3005
R1097 VCC.n750 VCC.n749 9.3005
R1098 VCC.n748 VCC.n12 9.3005
R1099 VCC.n747 VCC.n746 9.3005
R1100 VCC.n745 VCC.n16 9.3005
R1101 VCC.n744 VCC.n743 9.3005
R1102 VCC.n742 VCC.n17 9.3005
R1103 VCC.n741 VCC.n740 9.3005
R1104 VCC.n739 VCC.n21 9.3005
R1105 VCC.n738 VCC.n737 9.3005
R1106 VCC.n736 VCC.n22 9.3005
R1107 VCC.n735 VCC.n734 9.3005
R1108 VCC.n733 VCC.n26 9.3005
R1109 VCC.n732 VCC.n731 9.3005
R1110 VCC.n730 VCC.n27 9.3005
R1111 VCC.n729 VCC.n728 9.3005
R1112 VCC.n727 VCC.n31 9.3005
R1113 VCC.n726 VCC.n725 9.3005
R1114 VCC.n724 VCC.n32 9.3005
R1115 VCC.n723 VCC.n722 9.3005
R1116 VCC.n721 VCC.n36 9.3005
R1117 VCC.n720 VCC.n719 9.3005
R1118 VCC.n718 VCC.n37 9.3005
R1119 VCC.n349 VCC.n170 9.3005
R1120 VCC.n351 VCC.n350 9.3005
R1121 VCC.n160 VCC.n159 9.3005
R1122 VCC.n364 VCC.n363 9.3005
R1123 VCC.n365 VCC.n158 9.3005
R1124 VCC.n367 VCC.n366 9.3005
R1125 VCC.n148 VCC.n147 9.3005
R1126 VCC.n380 VCC.n379 9.3005
R1127 VCC.n381 VCC.n146 9.3005
R1128 VCC.n383 VCC.n382 9.3005
R1129 VCC.n136 VCC.n135 9.3005
R1130 VCC.n396 VCC.n395 9.3005
R1131 VCC.n397 VCC.n134 9.3005
R1132 VCC.n399 VCC.n398 9.3005
R1133 VCC.n124 VCC.n123 9.3005
R1134 VCC.n412 VCC.n411 9.3005
R1135 VCC.n413 VCC.n122 9.3005
R1136 VCC.n415 VCC.n414 9.3005
R1137 VCC.n111 VCC.n110 9.3005
R1138 VCC.n428 VCC.n427 9.3005
R1139 VCC.n429 VCC.n108 9.3005
R1140 VCC.n432 VCC.n431 9.3005
R1141 VCC.n430 VCC.n109 9.3005
R1142 VCC.n99 VCC.n98 9.3005
R1143 VCC.n446 VCC.n445 9.3005
R1144 VCC.n447 VCC.n97 9.3005
R1145 VCC.n449 VCC.n448 9.3005
R1146 VCC.n87 VCC.n86 9.3005
R1147 VCC.n464 VCC.n463 9.3005
R1148 VCC.n465 VCC.n85 9.3005
R1149 VCC.n467 VCC.n466 9.3005
R1150 VCC.n81 VCC.n80 9.3005
R1151 VCC.n475 VCC.n474 9.3005
R1152 VCC.n476 VCC.n79 9.3005
R1153 VCC.n478 VCC.n477 9.3005
R1154 VCC.n75 VCC.n74 9.3005
R1155 VCC.n486 VCC.n485 9.3005
R1156 VCC.n487 VCC.n73 9.3005
R1157 VCC.n489 VCC.n488 9.3005
R1158 VCC.n69 VCC.n68 9.3005
R1159 VCC.n497 VCC.n496 9.3005
R1160 VCC.n498 VCC.n67 9.3005
R1161 VCC.n500 VCC.n499 9.3005
R1162 VCC.n63 VCC.n62 9.3005
R1163 VCC.n508 VCC.n507 9.3005
R1164 VCC.n509 VCC.n61 9.3005
R1165 VCC.n511 VCC.n510 9.3005
R1166 VCC.n57 VCC.n56 9.3005
R1167 VCC.n519 VCC.n518 9.3005
R1168 VCC.n520 VCC.n55 9.3005
R1169 VCC.n522 VCC.n521 9.3005
R1170 VCC.n51 VCC.n50 9.3005
R1171 VCC.n531 VCC.n530 9.3005
R1172 VCC.n532 VCC.n49 9.3005
R1173 VCC.n534 VCC.n533 9.3005
R1174 VCC.n46 VCC.n45 9.3005
R1175 VCC.n542 VCC.n541 9.3005
R1176 VCC.n543 VCC.n44 9.3005
R1177 VCC.n714 VCC.n713 9.3005
R1178 VCC.n348 VCC.n347 9.3005
R1179 VCC.n343 VCC.n342 9.3005
R1180 VCC.n166 VCC.n165 9.3005
R1181 VCC.n356 VCC.n355 9.3005
R1182 VCC.n357 VCC.n164 9.3005
R1183 VCC.n359 VCC.n358 9.3005
R1184 VCC.n154 VCC.n153 9.3005
R1185 VCC.n372 VCC.n371 9.3005
R1186 VCC.n373 VCC.n152 9.3005
R1187 VCC.n375 VCC.n374 9.3005
R1188 VCC.n142 VCC.n141 9.3005
R1189 VCC.n388 VCC.n387 9.3005
R1190 VCC.n389 VCC.n140 9.3005
R1191 VCC.n391 VCC.n390 9.3005
R1192 VCC.n130 VCC.n129 9.3005
R1193 VCC.n404 VCC.n403 9.3005
R1194 VCC.n405 VCC.n128 9.3005
R1195 VCC.n407 VCC.n406 9.3005
R1196 VCC.n118 VCC.n117 9.3005
R1197 VCC.n420 VCC.n419 9.3005
R1198 VCC.n421 VCC.n116 9.3005
R1199 VCC.n423 VCC.n422 9.3005
R1200 VCC.n105 VCC.n104 9.3005
R1201 VCC.n437 VCC.n436 9.3005
R1202 VCC.n438 VCC.n103 9.3005
R1203 VCC.n440 VCC.n439 9.3005
R1204 VCC.n93 VCC.n92 9.3005
R1205 VCC.n455 VCC.n454 9.3005
R1206 VCC.n456 VCC.n91 9.3005
R1207 VCC.n458 VCC.n457 9.3005
R1208 VCC.n2 VCC.n1 9.3005
R1209 VCC VCC.n761 9.3005
R1210 VCC.n434 VCC.t0 4.69379
R1211 VCC.n483 VCC.t1 4.69379
R1212 VCC.n361 VCC.t10 1.95604
R1213 VCC.n536 VCC.t6 1.95604
R1214 VCC.n648 VCC.n558 0.780988
R1215 VCC.n272 VCC.n271 0.780988
R1216 VCC.n582 VCC.n581 0.468793
R1217 VCC.n179 VCC.n175 0.468793
R1218 VCC.n401 VCC.t4 0.391607
R1219 VCC.n505 VCC.t3 0.391607
R1220 VCC VCC.n0 0.152939
R1221 VCC.n758 VCC.n0 0.152939
R1222 VCC.n758 VCC.n757 0.152939
R1223 VCC.n757 VCC.n756 0.152939
R1224 VCC.n756 VCC.n7 0.152939
R1225 VCC.n752 VCC.n7 0.152939
R1226 VCC.n752 VCC.n751 0.152939
R1227 VCC.n751 VCC.n750 0.152939
R1228 VCC.n750 VCC.n12 0.152939
R1229 VCC.n746 VCC.n12 0.152939
R1230 VCC.n746 VCC.n745 0.152939
R1231 VCC.n745 VCC.n744 0.152939
R1232 VCC.n744 VCC.n17 0.152939
R1233 VCC.n740 VCC.n17 0.152939
R1234 VCC.n740 VCC.n739 0.152939
R1235 VCC.n739 VCC.n738 0.152939
R1236 VCC.n738 VCC.n22 0.152939
R1237 VCC.n734 VCC.n22 0.152939
R1238 VCC.n734 VCC.n733 0.152939
R1239 VCC.n733 VCC.n732 0.152939
R1240 VCC.n732 VCC.n27 0.152939
R1241 VCC.n728 VCC.n27 0.152939
R1242 VCC.n728 VCC.n727 0.152939
R1243 VCC.n727 VCC.n726 0.152939
R1244 VCC.n726 VCC.n32 0.152939
R1245 VCC.n722 VCC.n32 0.152939
R1246 VCC.n722 VCC.n721 0.152939
R1247 VCC.n721 VCC.n720 0.152939
R1248 VCC.n720 VCC.n37 0.152939
R1249 VCC.n349 VCC.n348 0.152939
R1250 VCC.n350 VCC.n349 0.152939
R1251 VCC.n350 VCC.n159 0.152939
R1252 VCC.n364 VCC.n159 0.152939
R1253 VCC.n365 VCC.n364 0.152939
R1254 VCC.n366 VCC.n365 0.152939
R1255 VCC.n366 VCC.n147 0.152939
R1256 VCC.n380 VCC.n147 0.152939
R1257 VCC.n381 VCC.n380 0.152939
R1258 VCC.n382 VCC.n381 0.152939
R1259 VCC.n382 VCC.n135 0.152939
R1260 VCC.n396 VCC.n135 0.152939
R1261 VCC.n397 VCC.n396 0.152939
R1262 VCC.n398 VCC.n397 0.152939
R1263 VCC.n398 VCC.n123 0.152939
R1264 VCC.n412 VCC.n123 0.152939
R1265 VCC.n413 VCC.n412 0.152939
R1266 VCC.n414 VCC.n413 0.152939
R1267 VCC.n414 VCC.n110 0.152939
R1268 VCC.n428 VCC.n110 0.152939
R1269 VCC.n429 VCC.n428 0.152939
R1270 VCC.n431 VCC.n429 0.152939
R1271 VCC.n431 VCC.n430 0.152939
R1272 VCC.n430 VCC.n98 0.152939
R1273 VCC.n446 VCC.n98 0.152939
R1274 VCC.n447 VCC.n446 0.152939
R1275 VCC.n448 VCC.n447 0.152939
R1276 VCC.n448 VCC.n86 0.152939
R1277 VCC.n464 VCC.n86 0.152939
R1278 VCC.n465 VCC.n464 0.152939
R1279 VCC.n466 VCC.n465 0.152939
R1280 VCC.n466 VCC.n80 0.152939
R1281 VCC.n475 VCC.n80 0.152939
R1282 VCC.n476 VCC.n475 0.152939
R1283 VCC.n477 VCC.n476 0.152939
R1284 VCC.n477 VCC.n74 0.152939
R1285 VCC.n486 VCC.n74 0.152939
R1286 VCC.n487 VCC.n486 0.152939
R1287 VCC.n488 VCC.n487 0.152939
R1288 VCC.n488 VCC.n68 0.152939
R1289 VCC.n497 VCC.n68 0.152939
R1290 VCC.n498 VCC.n497 0.152939
R1291 VCC.n499 VCC.n498 0.152939
R1292 VCC.n499 VCC.n62 0.152939
R1293 VCC.n508 VCC.n62 0.152939
R1294 VCC.n509 VCC.n508 0.152939
R1295 VCC.n510 VCC.n509 0.152939
R1296 VCC.n510 VCC.n56 0.152939
R1297 VCC.n519 VCC.n56 0.152939
R1298 VCC.n520 VCC.n519 0.152939
R1299 VCC.n521 VCC.n520 0.152939
R1300 VCC.n521 VCC.n50 0.152939
R1301 VCC.n531 VCC.n50 0.152939
R1302 VCC.n532 VCC.n531 0.152939
R1303 VCC.n533 VCC.n532 0.152939
R1304 VCC.n533 VCC.n45 0.152939
R1305 VCC.n542 VCC.n45 0.152939
R1306 VCC.n543 VCC.n542 0.152939
R1307 VCC.n713 VCC.n543 0.152939
R1308 VCC.n342 VCC.n165 0.152939
R1309 VCC.n356 VCC.n165 0.152939
R1310 VCC.n357 VCC.n356 0.152939
R1311 VCC.n358 VCC.n357 0.152939
R1312 VCC.n358 VCC.n153 0.152939
R1313 VCC.n372 VCC.n153 0.152939
R1314 VCC.n373 VCC.n372 0.152939
R1315 VCC.n374 VCC.n373 0.152939
R1316 VCC.n374 VCC.n141 0.152939
R1317 VCC.n388 VCC.n141 0.152939
R1318 VCC.n389 VCC.n388 0.152939
R1319 VCC.n390 VCC.n389 0.152939
R1320 VCC.n390 VCC.n129 0.152939
R1321 VCC.n404 VCC.n129 0.152939
R1322 VCC.n405 VCC.n404 0.152939
R1323 VCC.n406 VCC.n405 0.152939
R1324 VCC.n406 VCC.n117 0.152939
R1325 VCC.n420 VCC.n117 0.152939
R1326 VCC.n421 VCC.n420 0.152939
R1327 VCC.n422 VCC.n421 0.152939
R1328 VCC.n422 VCC.n104 0.152939
R1329 VCC.n437 VCC.n104 0.152939
R1330 VCC.n438 VCC.n437 0.152939
R1331 VCC.n439 VCC.n438 0.152939
R1332 VCC.n439 VCC.n92 0.152939
R1333 VCC.n455 VCC.n92 0.152939
R1334 VCC.n456 VCC.n455 0.152939
R1335 VCC.n457 VCC.n456 0.152939
R1336 VCC.n457 VCC.n1 0.152939
R1337 VCC VCC.n1 0.1255
R1338 VOUT.n16 VOUT.n15 161.3
R1339 VOUT.n17 VOUT.n12 161.3
R1340 VOUT.n19 VOUT.n18 161.3
R1341 VOUT.n20 VOUT.n11 161.3
R1342 VOUT.n22 VOUT.n21 161.3
R1343 VOUT.n23 VOUT.n10 161.3
R1344 VOUT.n25 VOUT.n24 161.3
R1345 VOUT.n26 VOUT.n9 161.3
R1346 VOUT.n28 VOUT.n27 161.3
R1347 VOUT.n29 VOUT.n8 161.3
R1348 VOUT.n31 VOUT.n30 161.3
R1349 VOUT.n32 VOUT.n7 161.3
R1350 VOUT.n34 VOUT.n33 161.3
R1351 VOUT.n35 VOUT.n5 161.3
R1352 VOUT.n37 VOUT.n36 161.3
R1353 VOUT.n38 VOUT.n4 161.3
R1354 VOUT.n40 VOUT.n39 161.3
R1355 VOUT.n41 VOUT.n3 161.3
R1356 VOUT.n43 VOUT.n42 161.3
R1357 VOUT.n44 VOUT.n2 161.3
R1358 VOUT.n46 VOUT.n45 161.3
R1359 VOUT.n47 VOUT.n1 161.3
R1360 VOUT.n49 VOUT.n48 161.3
R1361 VOUT.n108 VOUT.n107 161.3
R1362 VOUT.n106 VOUT.n60 161.3
R1363 VOUT.n105 VOUT.n104 161.3
R1364 VOUT.n103 VOUT.n61 161.3
R1365 VOUT.n102 VOUT.n101 161.3
R1366 VOUT.n100 VOUT.n62 161.3
R1367 VOUT.n99 VOUT.n98 161.3
R1368 VOUT.n97 VOUT.n63 161.3
R1369 VOUT.n96 VOUT.n95 161.3
R1370 VOUT.n94 VOUT.n64 161.3
R1371 VOUT.n93 VOUT.n92 161.3
R1372 VOUT.n91 VOUT.n66 161.3
R1373 VOUT.n90 VOUT.n89 161.3
R1374 VOUT.n88 VOUT.n67 161.3
R1375 VOUT.n87 VOUT.n86 161.3
R1376 VOUT.n85 VOUT.n68 161.3
R1377 VOUT.n84 VOUT.n83 161.3
R1378 VOUT.n82 VOUT.n69 161.3
R1379 VOUT.n81 VOUT.n80 161.3
R1380 VOUT.n79 VOUT.n70 161.3
R1381 VOUT.n78 VOUT.n77 161.3
R1382 VOUT.n76 VOUT.n71 161.3
R1383 VOUT.n75 VOUT.n74 161.3
R1384 VOUT.n73 VOUT.t31 94.458
R1385 VOUT.n14 VOUT.t16 94.4578
R1386 VOUT.t24 VOUT.n58 87.1613
R1387 VOUT.n57 VOUT.t28 87.1613
R1388 VOUT.n118 VOUT.n117 80.181
R1389 VOUT.n111 VOUT.n58 80.181
R1390 VOUT.n121 VOUT.n120 80.181
R1391 VOUT.n57 VOUT.n56 80.181
R1392 VOUT.n50 VOUT.n0 78.4415
R1393 VOUT.n109 VOUT.n59 78.4415
R1394 VOUT.n114 VOUT.t33 67.1463
R1395 VOUT.n124 VOUT.t18 67.1463
R1396 VOUT.n123 VOUT.n55 66.8384
R1397 VOUT.t7 VOUT.n126 64.6188
R1398 VOUT.n53 VOUT.t5 64.6188
R1399 VOUT.n116 VOUT.n115 63.5022
R1400 VOUT.n113 VOUT.n112 63.5022
R1401 VOUT.n123 VOUT.n122 63.5022
R1402 VOUT.n134 VOUT.n133 63.1086
R1403 VOUT.n127 VOUT.n126 63.1086
R1404 VOUT.n137 VOUT.n136 63.1086
R1405 VOUT.n139 VOUT.n53 63.1086
R1406 VOUT.n9 VOUT.t19 60.7271
R1407 VOUT.n0 VOUT.t27 60.7271
R1408 VOUT.n6 VOUT.t29 60.7271
R1409 VOUT.n13 VOUT.t21 60.7271
R1410 VOUT.n68 VOUT.t12 60.7271
R1411 VOUT.n72 VOUT.t14 60.7271
R1412 VOUT.n65 VOUT.t25 60.7271
R1413 VOUT.n59 VOUT.t23 60.7271
R1414 VOUT.n14 VOUT.n13 56.6961
R1415 VOUT.n73 VOUT.n72 56.696
R1416 VOUT.n42 VOUT.n2 56.5617
R1417 VOUT.n101 VOUT.n61 56.5617
R1418 VOUT.n129 VOUT.t11 47.4659
R1419 VOUT.n130 VOUT.t3 47.4659
R1420 VOUT.n131 VOUT.n128 46.904
R1421 VOUT.n30 VOUT.n7 46.874
R1422 VOUT.n22 VOUT.n11 46.874
R1423 VOUT.n81 VOUT.n70 46.874
R1424 VOUT.n89 VOUT.n66 46.874
R1425 VOUT.n138 VOUT.n52 46.4298
R1426 VOUT.n141 VOUT.n140 46.4298
R1427 VOUT.n132 VOUT.n131 46.4298
R1428 VOUT.n34 VOUT.n7 34.28
R1429 VOUT.n18 VOUT.n11 34.28
R1430 VOUT.n77 VOUT.n70 34.28
R1431 VOUT.n93 VOUT.n66 34.28
R1432 VOUT.n48 VOUT.n47 24.5923
R1433 VOUT.n47 VOUT.n46 24.5923
R1434 VOUT.n46 VOUT.n2 24.5923
R1435 VOUT.n42 VOUT.n41 24.5923
R1436 VOUT.n41 VOUT.n40 24.5923
R1437 VOUT.n40 VOUT.n4 24.5923
R1438 VOUT.n36 VOUT.n35 24.5923
R1439 VOUT.n35 VOUT.n34 24.5923
R1440 VOUT.n30 VOUT.n29 24.5923
R1441 VOUT.n29 VOUT.n28 24.5923
R1442 VOUT.n28 VOUT.n9 24.5923
R1443 VOUT.n24 VOUT.n9 24.5923
R1444 VOUT.n24 VOUT.n23 24.5923
R1445 VOUT.n23 VOUT.n22 24.5923
R1446 VOUT.n18 VOUT.n17 24.5923
R1447 VOUT.n17 VOUT.n16 24.5923
R1448 VOUT.n77 VOUT.n76 24.5923
R1449 VOUT.n76 VOUT.n75 24.5923
R1450 VOUT.n89 VOUT.n88 24.5923
R1451 VOUT.n88 VOUT.n87 24.5923
R1452 VOUT.n87 VOUT.n68 24.5923
R1453 VOUT.n83 VOUT.n68 24.5923
R1454 VOUT.n83 VOUT.n82 24.5923
R1455 VOUT.n82 VOUT.n81 24.5923
R1456 VOUT.n101 VOUT.n100 24.5923
R1457 VOUT.n100 VOUT.n99 24.5923
R1458 VOUT.n99 VOUT.n63 24.5923
R1459 VOUT.n95 VOUT.n94 24.5923
R1460 VOUT.n94 VOUT.n93 24.5923
R1461 VOUT.n107 VOUT.n106 24.5923
R1462 VOUT.n106 VOUT.n105 24.5923
R1463 VOUT.n105 VOUT.n61 24.5923
R1464 VIN VOUT.n51 23.5393
R1465 VOUT.n135 VOUT.n134 19.2936
R1466 VOUT.n130 VOUT.n129 18.9229
R1467 VOUT.n36 VOUT.n6 18.1985
R1468 VOUT.n16 VOUT.n13 18.1985
R1469 VOUT.n75 VOUT.n72 18.1985
R1470 VOUT.n95 VOUT.n65 18.1985
R1471 VOUT.n135 VOUT.n125 18.1947
R1472 VOUT.n120 VOUT.n119 16.8281
R1473 VOUT.n48 VOUT.n0 11.8046
R1474 VOUT.n107 VOUT.n59 11.8046
R1475 VOUT.n110 VGP 8.58249
R1476 VOUT.n113 VOUT.n110 6.50912
R1477 VOUT.n6 VOUT.n4 6.39438
R1478 VOUT.n65 VOUT.n63 6.39438
R1479 VOUT.n51 VOUT.n50 5.19889
R1480 VOUT.n114 VOUT.n54 5.06539
R1481 VOUT.n125 VOUT.n124 4.88412
R1482 VOUT.n119 VOUT.n54 4.5005
R1483 VOUT.n117 VOUT.t15 3.64456
R1484 VOUT.n117 VOUT.t32 3.64456
R1485 VOUT.t26 VOUT.n111 3.64456
R1486 VOUT.n111 VOUT.t13 3.64456
R1487 VOUT.n116 VOUT.t13 3.64456
R1488 VOUT.t15 VOUT.n116 3.64456
R1489 VOUT.n112 VOUT.t24 3.64456
R1490 VOUT.n112 VOUT.t26 3.64456
R1491 VOUT.n122 VOUT.t20 3.64456
R1492 VOUT.n122 VOUT.t22 3.64456
R1493 VOUT.t28 VOUT.n55 3.64456
R1494 VOUT.t30 VOUT.n55 3.64456
R1495 VOUT.t22 VOUT.n121 3.64456
R1496 VOUT.n121 VOUT.t17 3.64456
R1497 VOUT.n56 VOUT.t30 3.64456
R1498 VOUT.n56 VOUT.t20 3.64456
R1499 VOUT.n125 VOUT.n54 3.38017
R1500 VOUT.n115 VOUT.n113 3.33671
R1501 VOUT.n115 VOUT.n114 3.33671
R1502 VOUT.n124 VOUT.n123 3.33671
R1503 VOUT.n120 VOUT.n57 3.33671
R1504 VOUT.n118 VOUT.n58 3.33671
R1505 VOUT.n74 VOUT.n73 3.08737
R1506 VOUT.n15 VOUT.n14 3.08735
R1507 VOUT VOUT.n118 1.78929
R1508 VOUT.n136 VOUT.n135 1.13843
R1509 VOUT.t4 VOUT.n138 1.03661
R1510 VOUT.n138 VOUT.t9 1.03661
R1511 VOUT.n140 VOUT.t5 1.03661
R1512 VOUT.n140 VOUT.t8 1.03661
R1513 VOUT.n132 VOUT.t6 1.03661
R1514 VOUT.t1 VOUT.n132 1.03661
R1515 VOUT.n128 VOUT.t7 1.03661
R1516 VOUT.n128 VOUT.t0 1.03661
R1517 VOUT.n133 VOUT.t1 1.03661
R1518 VOUT.n133 VOUT.t2 1.03661
R1519 VOUT.t0 VOUT.n127 1.03661
R1520 VOUT.n127 VOUT.t6 1.03661
R1521 VOUT.t9 VOUT.n137 1.03661
R1522 VOUT.n137 VOUT.t10 1.03661
R1523 VOUT.t8 VOUT.n139 1.03661
R1524 VOUT.n139 VOUT.t4 1.03661
R1525 VOUT.n131 VOUT.n130 0.474638
R1526 VOUT.n141 VOUT.n52 0.474638
R1527 VOUT.n129 VOUT.n52 0.474638
R1528 VOUT.n134 VOUT.n126 0.474638
R1529 VOUT.n136 VOUT.n53 0.474638
R1530 VGP VOUT.n109 0.35798
R1531 VOUT.n50 VOUT.n49 0.354861
R1532 VOUT.n109 VOUT.n108 0.354861
R1533 VOUT.n110 VOUT.n51 0.282952
R1534 VIN VOUT.n141 0.241879
R1535 VOUT.n119 VOUT 0.220328
R1536 VOUT.n49 VOUT.n1 0.189894
R1537 VOUT.n45 VOUT.n1 0.189894
R1538 VOUT.n45 VOUT.n44 0.189894
R1539 VOUT.n44 VOUT.n43 0.189894
R1540 VOUT.n43 VOUT.n3 0.189894
R1541 VOUT.n39 VOUT.n3 0.189894
R1542 VOUT.n39 VOUT.n38 0.189894
R1543 VOUT.n38 VOUT.n37 0.189894
R1544 VOUT.n37 VOUT.n5 0.189894
R1545 VOUT.n33 VOUT.n5 0.189894
R1546 VOUT.n33 VOUT.n32 0.189894
R1547 VOUT.n32 VOUT.n31 0.189894
R1548 VOUT.n31 VOUT.n8 0.189894
R1549 VOUT.n27 VOUT.n8 0.189894
R1550 VOUT.n27 VOUT.n26 0.189894
R1551 VOUT.n26 VOUT.n25 0.189894
R1552 VOUT.n25 VOUT.n10 0.189894
R1553 VOUT.n21 VOUT.n10 0.189894
R1554 VOUT.n21 VOUT.n20 0.189894
R1555 VOUT.n20 VOUT.n19 0.189894
R1556 VOUT.n19 VOUT.n12 0.189894
R1557 VOUT.n15 VOUT.n12 0.189894
R1558 VOUT.n108 VOUT.n60 0.189894
R1559 VOUT.n104 VOUT.n60 0.189894
R1560 VOUT.n104 VOUT.n103 0.189894
R1561 VOUT.n103 VOUT.n102 0.189894
R1562 VOUT.n102 VOUT.n62 0.189894
R1563 VOUT.n98 VOUT.n62 0.189894
R1564 VOUT.n98 VOUT.n97 0.189894
R1565 VOUT.n97 VOUT.n96 0.189894
R1566 VOUT.n96 VOUT.n64 0.189894
R1567 VOUT.n92 VOUT.n64 0.189894
R1568 VOUT.n92 VOUT.n91 0.189894
R1569 VOUT.n91 VOUT.n90 0.189894
R1570 VOUT.n90 VOUT.n67 0.189894
R1571 VOUT.n86 VOUT.n67 0.189894
R1572 VOUT.n86 VOUT.n85 0.189894
R1573 VOUT.n85 VOUT.n84 0.189894
R1574 VOUT.n84 VOUT.n69 0.189894
R1575 VOUT.n80 VOUT.n69 0.189894
R1576 VOUT.n80 VOUT.n79 0.189894
R1577 VOUT.n79 VOUT.n78 0.189894
R1578 VOUT.n78 VOUT.n71 0.189894
R1579 VOUT.n74 VOUT.n71 0.189894
R1580 VGN.n18 VGN.t0 2288.04
R1581 VGN.n12 VGN.t7 2288.04
R1582 VGN.n8 VGN.t8 2288.04
R1583 VGN.n2 VGN.t2 2288.04
R1584 VGN.n17 VGN.t6 2236.92
R1585 VGN.n15 VGN.t1 2236.92
R1586 VGN.n11 VGN.t9 2236.92
R1587 VGN.n7 VGN.t5 2236.92
R1588 VGN.n5 VGN.t4 2236.92
R1589 VGN.n1 VGN.t3 2236.92
R1590 VGN.n13 VGN.n12 161.489
R1591 VGN.n3 VGN.n2 161.489
R1592 VGN.n9 VGN.n8 161.3
R1593 VGN.n6 VGN.n0 161.3
R1594 VGN.n4 VGN.n3 161.3
R1595 VGN.n14 VGN.n13 161.3
R1596 VGN.n16 VGN.n10 161.3
R1597 VGN.n19 VGN.n18 161.3
R1598 VGN.n17 VGN.n16 43.8187
R1599 VGN.n14 VGN.n11 43.8187
R1600 VGN.n7 VGN.n6 43.8187
R1601 VGN.n4 VGN.n1 43.8187
R1602 VGN.n16 VGN.n15 36.5157
R1603 VGN.n15 VGN.n14 36.5157
R1604 VGN.n6 VGN.n5 36.5157
R1605 VGN.n5 VGN.n4 36.5157
R1606 VGN.n18 VGN.n17 29.2126
R1607 VGN.n12 VGN.n11 29.2126
R1608 VGN.n8 VGN.n7 29.2126
R1609 VGN.n2 VGN.n1 29.2126
R1610 VGN VGN.n9 17.866
R1611 VGN.n9 VGN.n0 0.189894
R1612 VGN.n3 VGN.n0 0.189894
R1613 VGN.n19 VGN.n10 0.189894
R1614 VGN.n13 VGN.n10 0.189894
R1615 VGN VGN.n19 0.123606
R1616 VSS.n458 VSS.t11 2324.29
R1617 VSS.n508 VSS.t7 2324.29
R1618 VSS.n49 VSS.t4 2324.29
R1619 VSS.n84 VSS.t0 2324.29
R1620 VSS.n371 VSS.n44 622.232
R1621 VSS.n368 VSS.n46 622.232
R1622 VSS.n731 VSS.n17 622.232
R1623 VSS.n734 VSS.n733 622.232
R1624 VSS.n372 VSS.n371 585
R1625 VSS.n371 VSS.n370 585
R1626 VSS.n42 VSS.n41 585
R1627 VSS.n369 VSS.n41 585
R1628 VSS.n377 VSS.n376 585
R1629 VSS.n378 VSS.n377 585
R1630 VSS.n34 VSS.n33 585
R1631 VSS.n35 VSS.n34 585
R1632 VSS.n390 VSS.n389 585
R1633 VSS.n389 VSS.n388 585
R1634 VSS.n31 VSS.n30 585
R1635 VSS.n387 VSS.n30 585
R1636 VSS.n395 VSS.n394 585
R1637 VSS.n396 VSS.n395 585
R1638 VSS.n28 VSS.n27 585
R1639 VSS.n397 VSS.n28 585
R1640 VSS.n400 VSS.n399 585
R1641 VSS.n399 VSS.n398 585
R1642 VSS.n25 VSS.n24 585
R1643 VSS.n24 VSS.n22 585
R1644 VSS.n405 VSS.n404 585
R1645 VSS.n406 VSS.n405 585
R1646 VSS.n21 VSS.n20 585
R1647 VSS.n407 VSS.n21 585
R1648 VSS.n410 VSS.n409 585
R1649 VSS.n409 VSS.n408 585
R1650 VSS.n18 VSS.n16 585
R1651 VSS.n16 VSS.n14 585
R1652 VSS.n731 VSS.n730 585
R1653 VSS.n732 VSS.n731 585
R1654 VSS.n733 VSS.n11 585
R1655 VSS.n733 VSS.n732 585
R1656 VSS.n738 VSS.n10 585
R1657 VSS.n14 VSS.n10 585
R1658 VSS.n739 VSS.n9 585
R1659 VSS.n408 VSS.n9 585
R1660 VSS.n740 VSS.n8 585
R1661 VSS.n407 VSS.n8 585
R1662 VSS.n23 VSS.n6 585
R1663 VSS.n406 VSS.n23 585
R1664 VSS.n744 VSS.n5 585
R1665 VSS.n22 VSS.n5 585
R1666 VSS.n745 VSS.n4 585
R1667 VSS.n398 VSS.n4 585
R1668 VSS.n746 VSS.n3 585
R1669 VSS.n397 VSS.n3 585
R1670 VSS.n29 VSS.n2 585
R1671 VSS.n396 VSS.n29 585
R1672 VSS.n386 VSS.n385 585
R1673 VSS.n387 VSS.n386 585
R1674 VSS.n37 VSS.n36 585
R1675 VSS.n388 VSS.n36 585
R1676 VSS.n381 VSS.n380 585
R1677 VSS.n380 VSS.n35 585
R1678 VSS.n379 VSS.n39 585
R1679 VSS.n379 VSS.n378 585
R1680 VSS.n47 VSS.n40 585
R1681 VSS.n369 VSS.n40 585
R1682 VSS.n368 VSS.n367 585
R1683 VSS.n370 VSS.n368 585
R1684 VSS.n735 VSS.n734 585
R1685 VSS.n507 VSS.n12 585
R1686 VSS.n512 VSS.n511 585
R1687 VSS.n514 VSS.n505 585
R1688 VSS.n516 VSS.n515 585
R1689 VSS.n517 VSS.n504 585
R1690 VSS.n519 VSS.n518 585
R1691 VSS.n521 VSS.n502 585
R1692 VSS.n523 VSS.n522 585
R1693 VSS.n524 VSS.n501 585
R1694 VSS.n526 VSS.n525 585
R1695 VSS.n528 VSS.n499 585
R1696 VSS.n530 VSS.n529 585
R1697 VSS.n531 VSS.n498 585
R1698 VSS.n533 VSS.n532 585
R1699 VSS.n535 VSS.n496 585
R1700 VSS.n537 VSS.n536 585
R1701 VSS.n538 VSS.n495 585
R1702 VSS.n540 VSS.n539 585
R1703 VSS.n542 VSS.n493 585
R1704 VSS.n544 VSS.n543 585
R1705 VSS.n545 VSS.n492 585
R1706 VSS.n547 VSS.n546 585
R1707 VSS.n549 VSS.n490 585
R1708 VSS.n551 VSS.n550 585
R1709 VSS.n552 VSS.n489 585
R1710 VSS.n554 VSS.n553 585
R1711 VSS.n556 VSS.n487 585
R1712 VSS.n558 VSS.n557 585
R1713 VSS.n559 VSS.n486 585
R1714 VSS.n561 VSS.n560 585
R1715 VSS.n563 VSS.n484 585
R1716 VSS.n565 VSS.n564 585
R1717 VSS.n566 VSS.n483 585
R1718 VSS.n568 VSS.n567 585
R1719 VSS.n570 VSS.n481 585
R1720 VSS.n572 VSS.n571 585
R1721 VSS.n573 VSS.n480 585
R1722 VSS.n575 VSS.n574 585
R1723 VSS.n577 VSS.n478 585
R1724 VSS.n579 VSS.n578 585
R1725 VSS.n580 VSS.n477 585
R1726 VSS.n582 VSS.n581 585
R1727 VSS.n584 VSS.n475 585
R1728 VSS.n586 VSS.n585 585
R1729 VSS.n587 VSS.n474 585
R1730 VSS.n589 VSS.n588 585
R1731 VSS.n591 VSS.n472 585
R1732 VSS.n593 VSS.n592 585
R1733 VSS.n594 VSS.n471 585
R1734 VSS.n596 VSS.n595 585
R1735 VSS.n598 VSS.n469 585
R1736 VSS.n600 VSS.n599 585
R1737 VSS.n601 VSS.n468 585
R1738 VSS.n603 VSS.n602 585
R1739 VSS.n605 VSS.n466 585
R1740 VSS.n607 VSS.n606 585
R1741 VSS.n608 VSS.n465 585
R1742 VSS.n610 VSS.n609 585
R1743 VSS.n612 VSS.n463 585
R1744 VSS.n614 VSS.n613 585
R1745 VSS.n615 VSS.n462 585
R1746 VSS.n617 VSS.n616 585
R1747 VSS.n619 VSS.n460 585
R1748 VSS.n621 VSS.n620 585
R1749 VSS.n623 VSS.n457 585
R1750 VSS.n625 VSS.n624 585
R1751 VSS.n627 VSS.n455 585
R1752 VSS.n629 VSS.n628 585
R1753 VSS.n630 VSS.n454 585
R1754 VSS.n632 VSS.n631 585
R1755 VSS.n634 VSS.n452 585
R1756 VSS.n636 VSS.n635 585
R1757 VSS.n637 VSS.n451 585
R1758 VSS.n639 VSS.n638 585
R1759 VSS.n641 VSS.n449 585
R1760 VSS.n643 VSS.n642 585
R1761 VSS.n644 VSS.n448 585
R1762 VSS.n646 VSS.n645 585
R1763 VSS.n648 VSS.n446 585
R1764 VSS.n650 VSS.n649 585
R1765 VSS.n651 VSS.n445 585
R1766 VSS.n653 VSS.n652 585
R1767 VSS.n655 VSS.n443 585
R1768 VSS.n657 VSS.n656 585
R1769 VSS.n658 VSS.n442 585
R1770 VSS.n660 VSS.n659 585
R1771 VSS.n662 VSS.n440 585
R1772 VSS.n664 VSS.n663 585
R1773 VSS.n665 VSS.n439 585
R1774 VSS.n667 VSS.n666 585
R1775 VSS.n669 VSS.n437 585
R1776 VSS.n671 VSS.n670 585
R1777 VSS.n672 VSS.n436 585
R1778 VSS.n674 VSS.n673 585
R1779 VSS.n676 VSS.n434 585
R1780 VSS.n678 VSS.n677 585
R1781 VSS.n679 VSS.n433 585
R1782 VSS.n681 VSS.n680 585
R1783 VSS.n683 VSS.n431 585
R1784 VSS.n685 VSS.n684 585
R1785 VSS.n686 VSS.n430 585
R1786 VSS.n688 VSS.n687 585
R1787 VSS.n690 VSS.n428 585
R1788 VSS.n692 VSS.n691 585
R1789 VSS.n693 VSS.n427 585
R1790 VSS.n695 VSS.n694 585
R1791 VSS.n697 VSS.n425 585
R1792 VSS.n699 VSS.n698 585
R1793 VSS.n700 VSS.n424 585
R1794 VSS.n702 VSS.n701 585
R1795 VSS.n704 VSS.n422 585
R1796 VSS.n706 VSS.n705 585
R1797 VSS.n707 VSS.n421 585
R1798 VSS.n709 VSS.n708 585
R1799 VSS.n711 VSS.n419 585
R1800 VSS.n713 VSS.n712 585
R1801 VSS.n714 VSS.n418 585
R1802 VSS.n716 VSS.n715 585
R1803 VSS.n718 VSS.n416 585
R1804 VSS.n720 VSS.n719 585
R1805 VSS.n721 VSS.n415 585
R1806 VSS.n723 VSS.n722 585
R1807 VSS.n725 VSS.n413 585
R1808 VSS.n727 VSS.n726 585
R1809 VSS.n728 VSS.n17 585
R1810 VSS.n44 VSS.n43 585
R1811 VSS.n117 VSS.n115 585
R1812 VSS.n118 VSS.n114 585
R1813 VSS.n118 VSS.n45 585
R1814 VSS.n121 VSS.n120 585
R1815 VSS.n122 VSS.n113 585
R1816 VSS.n124 VSS.n123 585
R1817 VSS.n126 VSS.n112 585
R1818 VSS.n129 VSS.n128 585
R1819 VSS.n130 VSS.n111 585
R1820 VSS.n132 VSS.n131 585
R1821 VSS.n134 VSS.n110 585
R1822 VSS.n137 VSS.n136 585
R1823 VSS.n138 VSS.n109 585
R1824 VSS.n140 VSS.n139 585
R1825 VSS.n142 VSS.n108 585
R1826 VSS.n145 VSS.n144 585
R1827 VSS.n146 VSS.n107 585
R1828 VSS.n148 VSS.n147 585
R1829 VSS.n150 VSS.n106 585
R1830 VSS.n153 VSS.n152 585
R1831 VSS.n154 VSS.n105 585
R1832 VSS.n156 VSS.n155 585
R1833 VSS.n158 VSS.n104 585
R1834 VSS.n161 VSS.n160 585
R1835 VSS.n162 VSS.n103 585
R1836 VSS.n164 VSS.n163 585
R1837 VSS.n166 VSS.n102 585
R1838 VSS.n169 VSS.n168 585
R1839 VSS.n170 VSS.n101 585
R1840 VSS.n172 VSS.n171 585
R1841 VSS.n174 VSS.n100 585
R1842 VSS.n177 VSS.n176 585
R1843 VSS.n178 VSS.n99 585
R1844 VSS.n180 VSS.n179 585
R1845 VSS.n182 VSS.n98 585
R1846 VSS.n185 VSS.n184 585
R1847 VSS.n186 VSS.n97 585
R1848 VSS.n188 VSS.n187 585
R1849 VSS.n190 VSS.n96 585
R1850 VSS.n193 VSS.n192 585
R1851 VSS.n194 VSS.n95 585
R1852 VSS.n196 VSS.n195 585
R1853 VSS.n198 VSS.n94 585
R1854 VSS.n201 VSS.n200 585
R1855 VSS.n202 VSS.n93 585
R1856 VSS.n204 VSS.n203 585
R1857 VSS.n206 VSS.n92 585
R1858 VSS.n209 VSS.n208 585
R1859 VSS.n210 VSS.n91 585
R1860 VSS.n212 VSS.n211 585
R1861 VSS.n214 VSS.n90 585
R1862 VSS.n217 VSS.n216 585
R1863 VSS.n218 VSS.n89 585
R1864 VSS.n220 VSS.n219 585
R1865 VSS.n222 VSS.n88 585
R1866 VSS.n225 VSS.n224 585
R1867 VSS.n226 VSS.n87 585
R1868 VSS.n228 VSS.n227 585
R1869 VSS.n230 VSS.n86 585
R1870 VSS.n233 VSS.n232 585
R1871 VSS.n234 VSS.n83 585
R1872 VSS.n237 VSS.n236 585
R1873 VSS.n239 VSS.n82 585
R1874 VSS.n242 VSS.n241 585
R1875 VSS.n243 VSS.n81 585
R1876 VSS.n245 VSS.n244 585
R1877 VSS.n247 VSS.n80 585
R1878 VSS.n250 VSS.n249 585
R1879 VSS.n251 VSS.n79 585
R1880 VSS.n253 VSS.n252 585
R1881 VSS.n255 VSS.n78 585
R1882 VSS.n258 VSS.n257 585
R1883 VSS.n259 VSS.n77 585
R1884 VSS.n261 VSS.n260 585
R1885 VSS.n263 VSS.n76 585
R1886 VSS.n266 VSS.n265 585
R1887 VSS.n267 VSS.n75 585
R1888 VSS.n269 VSS.n268 585
R1889 VSS.n271 VSS.n74 585
R1890 VSS.n274 VSS.n273 585
R1891 VSS.n275 VSS.n73 585
R1892 VSS.n277 VSS.n276 585
R1893 VSS.n279 VSS.n72 585
R1894 VSS.n282 VSS.n281 585
R1895 VSS.n283 VSS.n71 585
R1896 VSS.n285 VSS.n284 585
R1897 VSS.n287 VSS.n70 585
R1898 VSS.n290 VSS.n289 585
R1899 VSS.n291 VSS.n69 585
R1900 VSS.n293 VSS.n292 585
R1901 VSS.n295 VSS.n68 585
R1902 VSS.n298 VSS.n297 585
R1903 VSS.n299 VSS.n67 585
R1904 VSS.n301 VSS.n300 585
R1905 VSS.n303 VSS.n66 585
R1906 VSS.n306 VSS.n305 585
R1907 VSS.n307 VSS.n65 585
R1908 VSS.n309 VSS.n308 585
R1909 VSS.n311 VSS.n64 585
R1910 VSS.n314 VSS.n313 585
R1911 VSS.n315 VSS.n63 585
R1912 VSS.n317 VSS.n316 585
R1913 VSS.n319 VSS.n62 585
R1914 VSS.n322 VSS.n321 585
R1915 VSS.n323 VSS.n61 585
R1916 VSS.n325 VSS.n324 585
R1917 VSS.n327 VSS.n60 585
R1918 VSS.n330 VSS.n329 585
R1919 VSS.n331 VSS.n59 585
R1920 VSS.n333 VSS.n332 585
R1921 VSS.n335 VSS.n58 585
R1922 VSS.n338 VSS.n337 585
R1923 VSS.n339 VSS.n57 585
R1924 VSS.n341 VSS.n340 585
R1925 VSS.n343 VSS.n56 585
R1926 VSS.n346 VSS.n345 585
R1927 VSS.n347 VSS.n55 585
R1928 VSS.n349 VSS.n348 585
R1929 VSS.n351 VSS.n54 585
R1930 VSS.n354 VSS.n353 585
R1931 VSS.n355 VSS.n53 585
R1932 VSS.n357 VSS.n356 585
R1933 VSS.n359 VSS.n52 585
R1934 VSS.n360 VSS.n48 585
R1935 VSS.n363 VSS.n362 585
R1936 VSS.n364 VSS.n46 585
R1937 VSS.n46 VSS.n45 585
R1938 VSS.n15 VSS.n13 256.663
R1939 VSS.n513 VSS.n15 256.663
R1940 VSS.n506 VSS.n15 256.663
R1941 VSS.n520 VSS.n15 256.663
R1942 VSS.n503 VSS.n15 256.663
R1943 VSS.n527 VSS.n15 256.663
R1944 VSS.n500 VSS.n15 256.663
R1945 VSS.n534 VSS.n15 256.663
R1946 VSS.n497 VSS.n15 256.663
R1947 VSS.n541 VSS.n15 256.663
R1948 VSS.n494 VSS.n15 256.663
R1949 VSS.n548 VSS.n15 256.663
R1950 VSS.n491 VSS.n15 256.663
R1951 VSS.n555 VSS.n15 256.663
R1952 VSS.n488 VSS.n15 256.663
R1953 VSS.n562 VSS.n15 256.663
R1954 VSS.n485 VSS.n15 256.663
R1955 VSS.n569 VSS.n15 256.663
R1956 VSS.n482 VSS.n15 256.663
R1957 VSS.n576 VSS.n15 256.663
R1958 VSS.n479 VSS.n15 256.663
R1959 VSS.n583 VSS.n15 256.663
R1960 VSS.n476 VSS.n15 256.663
R1961 VSS.n590 VSS.n15 256.663
R1962 VSS.n473 VSS.n15 256.663
R1963 VSS.n597 VSS.n15 256.663
R1964 VSS.n470 VSS.n15 256.663
R1965 VSS.n604 VSS.n15 256.663
R1966 VSS.n467 VSS.n15 256.663
R1967 VSS.n611 VSS.n15 256.663
R1968 VSS.n464 VSS.n15 256.663
R1969 VSS.n618 VSS.n15 256.663
R1970 VSS.n461 VSS.n15 256.663
R1971 VSS.n626 VSS.n15 256.663
R1972 VSS.n456 VSS.n15 256.663
R1973 VSS.n633 VSS.n15 256.663
R1974 VSS.n453 VSS.n15 256.663
R1975 VSS.n640 VSS.n15 256.663
R1976 VSS.n450 VSS.n15 256.663
R1977 VSS.n647 VSS.n15 256.663
R1978 VSS.n447 VSS.n15 256.663
R1979 VSS.n654 VSS.n15 256.663
R1980 VSS.n444 VSS.n15 256.663
R1981 VSS.n661 VSS.n15 256.663
R1982 VSS.n441 VSS.n15 256.663
R1983 VSS.n668 VSS.n15 256.663
R1984 VSS.n438 VSS.n15 256.663
R1985 VSS.n675 VSS.n15 256.663
R1986 VSS.n435 VSS.n15 256.663
R1987 VSS.n682 VSS.n15 256.663
R1988 VSS.n432 VSS.n15 256.663
R1989 VSS.n689 VSS.n15 256.663
R1990 VSS.n429 VSS.n15 256.663
R1991 VSS.n696 VSS.n15 256.663
R1992 VSS.n426 VSS.n15 256.663
R1993 VSS.n703 VSS.n15 256.663
R1994 VSS.n423 VSS.n15 256.663
R1995 VSS.n710 VSS.n15 256.663
R1996 VSS.n420 VSS.n15 256.663
R1997 VSS.n717 VSS.n15 256.663
R1998 VSS.n417 VSS.n15 256.663
R1999 VSS.n724 VSS.n15 256.663
R2000 VSS.n414 VSS.n15 256.663
R2001 VSS.n116 VSS.n45 256.663
R2002 VSS.n119 VSS.n45 256.663
R2003 VSS.n125 VSS.n45 256.663
R2004 VSS.n127 VSS.n45 256.663
R2005 VSS.n133 VSS.n45 256.663
R2006 VSS.n135 VSS.n45 256.663
R2007 VSS.n141 VSS.n45 256.663
R2008 VSS.n143 VSS.n45 256.663
R2009 VSS.n149 VSS.n45 256.663
R2010 VSS.n151 VSS.n45 256.663
R2011 VSS.n157 VSS.n45 256.663
R2012 VSS.n159 VSS.n45 256.663
R2013 VSS.n165 VSS.n45 256.663
R2014 VSS.n167 VSS.n45 256.663
R2015 VSS.n173 VSS.n45 256.663
R2016 VSS.n175 VSS.n45 256.663
R2017 VSS.n181 VSS.n45 256.663
R2018 VSS.n183 VSS.n45 256.663
R2019 VSS.n189 VSS.n45 256.663
R2020 VSS.n191 VSS.n45 256.663
R2021 VSS.n197 VSS.n45 256.663
R2022 VSS.n199 VSS.n45 256.663
R2023 VSS.n205 VSS.n45 256.663
R2024 VSS.n207 VSS.n45 256.663
R2025 VSS.n213 VSS.n45 256.663
R2026 VSS.n215 VSS.n45 256.663
R2027 VSS.n221 VSS.n45 256.663
R2028 VSS.n223 VSS.n45 256.663
R2029 VSS.n229 VSS.n45 256.663
R2030 VSS.n231 VSS.n45 256.663
R2031 VSS.n238 VSS.n45 256.663
R2032 VSS.n240 VSS.n45 256.663
R2033 VSS.n246 VSS.n45 256.663
R2034 VSS.n248 VSS.n45 256.663
R2035 VSS.n254 VSS.n45 256.663
R2036 VSS.n256 VSS.n45 256.663
R2037 VSS.n262 VSS.n45 256.663
R2038 VSS.n264 VSS.n45 256.663
R2039 VSS.n270 VSS.n45 256.663
R2040 VSS.n272 VSS.n45 256.663
R2041 VSS.n278 VSS.n45 256.663
R2042 VSS.n280 VSS.n45 256.663
R2043 VSS.n286 VSS.n45 256.663
R2044 VSS.n288 VSS.n45 256.663
R2045 VSS.n294 VSS.n45 256.663
R2046 VSS.n296 VSS.n45 256.663
R2047 VSS.n302 VSS.n45 256.663
R2048 VSS.n304 VSS.n45 256.663
R2049 VSS.n310 VSS.n45 256.663
R2050 VSS.n312 VSS.n45 256.663
R2051 VSS.n318 VSS.n45 256.663
R2052 VSS.n320 VSS.n45 256.663
R2053 VSS.n326 VSS.n45 256.663
R2054 VSS.n328 VSS.n45 256.663
R2055 VSS.n334 VSS.n45 256.663
R2056 VSS.n336 VSS.n45 256.663
R2057 VSS.n342 VSS.n45 256.663
R2058 VSS.n344 VSS.n45 256.663
R2059 VSS.n350 VSS.n45 256.663
R2060 VSS.n352 VSS.n45 256.663
R2061 VSS.n358 VSS.n45 256.663
R2062 VSS.n361 VSS.n45 256.663
R2063 VSS.n371 VSS.n41 240.244
R2064 VSS.n377 VSS.n41 240.244
R2065 VSS.n377 VSS.n34 240.244
R2066 VSS.n389 VSS.n34 240.244
R2067 VSS.n389 VSS.n30 240.244
R2068 VSS.n395 VSS.n30 240.244
R2069 VSS.n395 VSS.n28 240.244
R2070 VSS.n399 VSS.n28 240.244
R2071 VSS.n399 VSS.n24 240.244
R2072 VSS.n405 VSS.n24 240.244
R2073 VSS.n405 VSS.n21 240.244
R2074 VSS.n409 VSS.n21 240.244
R2075 VSS.n409 VSS.n16 240.244
R2076 VSS.n731 VSS.n16 240.244
R2077 VSS.n368 VSS.n40 240.244
R2078 VSS.n379 VSS.n40 240.244
R2079 VSS.n380 VSS.n379 240.244
R2080 VSS.n380 VSS.n36 240.244
R2081 VSS.n386 VSS.n36 240.244
R2082 VSS.n386 VSS.n29 240.244
R2083 VSS.n29 VSS.n3 240.244
R2084 VSS.n4 VSS.n3 240.244
R2085 VSS.n5 VSS.n4 240.244
R2086 VSS.n23 VSS.n5 240.244
R2087 VSS.n23 VSS.n8 240.244
R2088 VSS.n9 VSS.n8 240.244
R2089 VSS.n10 VSS.n9 240.244
R2090 VSS.n733 VSS.n10 240.244
R2091 VSS.n118 VSS.n117 163.367
R2092 VSS.n120 VSS.n118 163.367
R2093 VSS.n124 VSS.n113 163.367
R2094 VSS.n128 VSS.n126 163.367
R2095 VSS.n132 VSS.n111 163.367
R2096 VSS.n136 VSS.n134 163.367
R2097 VSS.n140 VSS.n109 163.367
R2098 VSS.n144 VSS.n142 163.367
R2099 VSS.n148 VSS.n107 163.367
R2100 VSS.n152 VSS.n150 163.367
R2101 VSS.n156 VSS.n105 163.367
R2102 VSS.n160 VSS.n158 163.367
R2103 VSS.n164 VSS.n103 163.367
R2104 VSS.n168 VSS.n166 163.367
R2105 VSS.n172 VSS.n101 163.367
R2106 VSS.n176 VSS.n174 163.367
R2107 VSS.n180 VSS.n99 163.367
R2108 VSS.n184 VSS.n182 163.367
R2109 VSS.n188 VSS.n97 163.367
R2110 VSS.n192 VSS.n190 163.367
R2111 VSS.n196 VSS.n95 163.367
R2112 VSS.n200 VSS.n198 163.367
R2113 VSS.n204 VSS.n93 163.367
R2114 VSS.n208 VSS.n206 163.367
R2115 VSS.n212 VSS.n91 163.367
R2116 VSS.n216 VSS.n214 163.367
R2117 VSS.n220 VSS.n89 163.367
R2118 VSS.n224 VSS.n222 163.367
R2119 VSS.n228 VSS.n87 163.367
R2120 VSS.n232 VSS.n230 163.367
R2121 VSS.n237 VSS.n83 163.367
R2122 VSS.n241 VSS.n239 163.367
R2123 VSS.n245 VSS.n81 163.367
R2124 VSS.n249 VSS.n247 163.367
R2125 VSS.n253 VSS.n79 163.367
R2126 VSS.n257 VSS.n255 163.367
R2127 VSS.n261 VSS.n77 163.367
R2128 VSS.n265 VSS.n263 163.367
R2129 VSS.n269 VSS.n75 163.367
R2130 VSS.n273 VSS.n271 163.367
R2131 VSS.n277 VSS.n73 163.367
R2132 VSS.n281 VSS.n279 163.367
R2133 VSS.n285 VSS.n71 163.367
R2134 VSS.n289 VSS.n287 163.367
R2135 VSS.n293 VSS.n69 163.367
R2136 VSS.n297 VSS.n295 163.367
R2137 VSS.n301 VSS.n67 163.367
R2138 VSS.n305 VSS.n303 163.367
R2139 VSS.n309 VSS.n65 163.367
R2140 VSS.n313 VSS.n311 163.367
R2141 VSS.n317 VSS.n63 163.367
R2142 VSS.n321 VSS.n319 163.367
R2143 VSS.n325 VSS.n61 163.367
R2144 VSS.n329 VSS.n327 163.367
R2145 VSS.n333 VSS.n59 163.367
R2146 VSS.n337 VSS.n335 163.367
R2147 VSS.n341 VSS.n57 163.367
R2148 VSS.n345 VSS.n343 163.367
R2149 VSS.n349 VSS.n55 163.367
R2150 VSS.n353 VSS.n351 163.367
R2151 VSS.n357 VSS.n53 163.367
R2152 VSS.n360 VSS.n359 163.367
R2153 VSS.n362 VSS.n46 163.367
R2154 VSS.n726 VSS.n725 163.367
R2155 VSS.n723 VSS.n415 163.367
R2156 VSS.n719 VSS.n718 163.367
R2157 VSS.n716 VSS.n418 163.367
R2158 VSS.n712 VSS.n711 163.367
R2159 VSS.n709 VSS.n421 163.367
R2160 VSS.n705 VSS.n704 163.367
R2161 VSS.n702 VSS.n424 163.367
R2162 VSS.n698 VSS.n697 163.367
R2163 VSS.n695 VSS.n427 163.367
R2164 VSS.n691 VSS.n690 163.367
R2165 VSS.n688 VSS.n430 163.367
R2166 VSS.n684 VSS.n683 163.367
R2167 VSS.n681 VSS.n433 163.367
R2168 VSS.n677 VSS.n676 163.367
R2169 VSS.n674 VSS.n436 163.367
R2170 VSS.n670 VSS.n669 163.367
R2171 VSS.n667 VSS.n439 163.367
R2172 VSS.n663 VSS.n662 163.367
R2173 VSS.n660 VSS.n442 163.367
R2174 VSS.n656 VSS.n655 163.367
R2175 VSS.n653 VSS.n445 163.367
R2176 VSS.n649 VSS.n648 163.367
R2177 VSS.n646 VSS.n448 163.367
R2178 VSS.n642 VSS.n641 163.367
R2179 VSS.n639 VSS.n451 163.367
R2180 VSS.n635 VSS.n634 163.367
R2181 VSS.n632 VSS.n454 163.367
R2182 VSS.n628 VSS.n627 163.367
R2183 VSS.n625 VSS.n457 163.367
R2184 VSS.n620 VSS.n619 163.367
R2185 VSS.n617 VSS.n462 163.367
R2186 VSS.n613 VSS.n612 163.367
R2187 VSS.n610 VSS.n465 163.367
R2188 VSS.n606 VSS.n605 163.367
R2189 VSS.n603 VSS.n468 163.367
R2190 VSS.n599 VSS.n598 163.367
R2191 VSS.n596 VSS.n471 163.367
R2192 VSS.n592 VSS.n591 163.367
R2193 VSS.n589 VSS.n474 163.367
R2194 VSS.n585 VSS.n584 163.367
R2195 VSS.n582 VSS.n477 163.367
R2196 VSS.n578 VSS.n577 163.367
R2197 VSS.n575 VSS.n480 163.367
R2198 VSS.n571 VSS.n570 163.367
R2199 VSS.n568 VSS.n483 163.367
R2200 VSS.n564 VSS.n563 163.367
R2201 VSS.n561 VSS.n486 163.367
R2202 VSS.n557 VSS.n556 163.367
R2203 VSS.n554 VSS.n489 163.367
R2204 VSS.n550 VSS.n549 163.367
R2205 VSS.n547 VSS.n492 163.367
R2206 VSS.n543 VSS.n542 163.367
R2207 VSS.n540 VSS.n495 163.367
R2208 VSS.n536 VSS.n535 163.367
R2209 VSS.n533 VSS.n498 163.367
R2210 VSS.n529 VSS.n528 163.367
R2211 VSS.n526 VSS.n501 163.367
R2212 VSS.n522 VSS.n521 163.367
R2213 VSS.n519 VSS.n504 163.367
R2214 VSS.n515 VSS.n514 163.367
R2215 VSS.n512 VSS.n507 163.367
R2216 VSS.n458 VSS.t12 79.185
R2217 VSS.n508 VSS.t9 79.185
R2218 VSS.n49 VSS.t6 79.185
R2219 VSS.n84 VSS.t3 79.185
R2220 VSS.n370 VSS.n45 77.4584
R2221 VSS.n732 VSS.n15 77.4584
R2222 VSS.n116 VSS.n44 71.676
R2223 VSS.n120 VSS.n119 71.676
R2224 VSS.n125 VSS.n124 71.676
R2225 VSS.n128 VSS.n127 71.676
R2226 VSS.n133 VSS.n132 71.676
R2227 VSS.n136 VSS.n135 71.676
R2228 VSS.n141 VSS.n140 71.676
R2229 VSS.n144 VSS.n143 71.676
R2230 VSS.n149 VSS.n148 71.676
R2231 VSS.n152 VSS.n151 71.676
R2232 VSS.n157 VSS.n156 71.676
R2233 VSS.n160 VSS.n159 71.676
R2234 VSS.n165 VSS.n164 71.676
R2235 VSS.n168 VSS.n167 71.676
R2236 VSS.n173 VSS.n172 71.676
R2237 VSS.n176 VSS.n175 71.676
R2238 VSS.n181 VSS.n180 71.676
R2239 VSS.n184 VSS.n183 71.676
R2240 VSS.n189 VSS.n188 71.676
R2241 VSS.n192 VSS.n191 71.676
R2242 VSS.n197 VSS.n196 71.676
R2243 VSS.n200 VSS.n199 71.676
R2244 VSS.n205 VSS.n204 71.676
R2245 VSS.n208 VSS.n207 71.676
R2246 VSS.n213 VSS.n212 71.676
R2247 VSS.n216 VSS.n215 71.676
R2248 VSS.n221 VSS.n220 71.676
R2249 VSS.n224 VSS.n223 71.676
R2250 VSS.n229 VSS.n228 71.676
R2251 VSS.n232 VSS.n231 71.676
R2252 VSS.n238 VSS.n237 71.676
R2253 VSS.n241 VSS.n240 71.676
R2254 VSS.n246 VSS.n245 71.676
R2255 VSS.n249 VSS.n248 71.676
R2256 VSS.n254 VSS.n253 71.676
R2257 VSS.n257 VSS.n256 71.676
R2258 VSS.n262 VSS.n261 71.676
R2259 VSS.n265 VSS.n264 71.676
R2260 VSS.n270 VSS.n269 71.676
R2261 VSS.n273 VSS.n272 71.676
R2262 VSS.n278 VSS.n277 71.676
R2263 VSS.n281 VSS.n280 71.676
R2264 VSS.n286 VSS.n285 71.676
R2265 VSS.n289 VSS.n288 71.676
R2266 VSS.n294 VSS.n293 71.676
R2267 VSS.n297 VSS.n296 71.676
R2268 VSS.n302 VSS.n301 71.676
R2269 VSS.n305 VSS.n304 71.676
R2270 VSS.n310 VSS.n309 71.676
R2271 VSS.n313 VSS.n312 71.676
R2272 VSS.n318 VSS.n317 71.676
R2273 VSS.n321 VSS.n320 71.676
R2274 VSS.n326 VSS.n325 71.676
R2275 VSS.n329 VSS.n328 71.676
R2276 VSS.n334 VSS.n333 71.676
R2277 VSS.n337 VSS.n336 71.676
R2278 VSS.n342 VSS.n341 71.676
R2279 VSS.n345 VSS.n344 71.676
R2280 VSS.n350 VSS.n349 71.676
R2281 VSS.n353 VSS.n352 71.676
R2282 VSS.n358 VSS.n357 71.676
R2283 VSS.n361 VSS.n360 71.676
R2284 VSS.n726 VSS.n414 71.676
R2285 VSS.n724 VSS.n723 71.676
R2286 VSS.n719 VSS.n417 71.676
R2287 VSS.n717 VSS.n716 71.676
R2288 VSS.n712 VSS.n420 71.676
R2289 VSS.n710 VSS.n709 71.676
R2290 VSS.n705 VSS.n423 71.676
R2291 VSS.n703 VSS.n702 71.676
R2292 VSS.n698 VSS.n426 71.676
R2293 VSS.n696 VSS.n695 71.676
R2294 VSS.n691 VSS.n429 71.676
R2295 VSS.n689 VSS.n688 71.676
R2296 VSS.n684 VSS.n432 71.676
R2297 VSS.n682 VSS.n681 71.676
R2298 VSS.n677 VSS.n435 71.676
R2299 VSS.n675 VSS.n674 71.676
R2300 VSS.n670 VSS.n438 71.676
R2301 VSS.n668 VSS.n667 71.676
R2302 VSS.n663 VSS.n441 71.676
R2303 VSS.n661 VSS.n660 71.676
R2304 VSS.n656 VSS.n444 71.676
R2305 VSS.n654 VSS.n653 71.676
R2306 VSS.n649 VSS.n447 71.676
R2307 VSS.n647 VSS.n646 71.676
R2308 VSS.n642 VSS.n450 71.676
R2309 VSS.n640 VSS.n639 71.676
R2310 VSS.n635 VSS.n453 71.676
R2311 VSS.n633 VSS.n632 71.676
R2312 VSS.n628 VSS.n456 71.676
R2313 VSS.n626 VSS.n625 71.676
R2314 VSS.n620 VSS.n461 71.676
R2315 VSS.n618 VSS.n617 71.676
R2316 VSS.n613 VSS.n464 71.676
R2317 VSS.n611 VSS.n610 71.676
R2318 VSS.n606 VSS.n467 71.676
R2319 VSS.n604 VSS.n603 71.676
R2320 VSS.n599 VSS.n470 71.676
R2321 VSS.n597 VSS.n596 71.676
R2322 VSS.n592 VSS.n473 71.676
R2323 VSS.n590 VSS.n589 71.676
R2324 VSS.n585 VSS.n476 71.676
R2325 VSS.n583 VSS.n582 71.676
R2326 VSS.n578 VSS.n479 71.676
R2327 VSS.n576 VSS.n575 71.676
R2328 VSS.n571 VSS.n482 71.676
R2329 VSS.n569 VSS.n568 71.676
R2330 VSS.n564 VSS.n485 71.676
R2331 VSS.n562 VSS.n561 71.676
R2332 VSS.n557 VSS.n488 71.676
R2333 VSS.n555 VSS.n554 71.676
R2334 VSS.n550 VSS.n491 71.676
R2335 VSS.n548 VSS.n547 71.676
R2336 VSS.n543 VSS.n494 71.676
R2337 VSS.n541 VSS.n540 71.676
R2338 VSS.n536 VSS.n497 71.676
R2339 VSS.n534 VSS.n533 71.676
R2340 VSS.n529 VSS.n500 71.676
R2341 VSS.n527 VSS.n526 71.676
R2342 VSS.n522 VSS.n503 71.676
R2343 VSS.n520 VSS.n519 71.676
R2344 VSS.n515 VSS.n506 71.676
R2345 VSS.n513 VSS.n512 71.676
R2346 VSS.n734 VSS.n13 71.676
R2347 VSS.n507 VSS.n13 71.676
R2348 VSS.n514 VSS.n513 71.676
R2349 VSS.n506 VSS.n504 71.676
R2350 VSS.n521 VSS.n520 71.676
R2351 VSS.n503 VSS.n501 71.676
R2352 VSS.n528 VSS.n527 71.676
R2353 VSS.n500 VSS.n498 71.676
R2354 VSS.n535 VSS.n534 71.676
R2355 VSS.n497 VSS.n495 71.676
R2356 VSS.n542 VSS.n541 71.676
R2357 VSS.n494 VSS.n492 71.676
R2358 VSS.n549 VSS.n548 71.676
R2359 VSS.n491 VSS.n489 71.676
R2360 VSS.n556 VSS.n555 71.676
R2361 VSS.n488 VSS.n486 71.676
R2362 VSS.n563 VSS.n562 71.676
R2363 VSS.n485 VSS.n483 71.676
R2364 VSS.n570 VSS.n569 71.676
R2365 VSS.n482 VSS.n480 71.676
R2366 VSS.n577 VSS.n576 71.676
R2367 VSS.n479 VSS.n477 71.676
R2368 VSS.n584 VSS.n583 71.676
R2369 VSS.n476 VSS.n474 71.676
R2370 VSS.n591 VSS.n590 71.676
R2371 VSS.n473 VSS.n471 71.676
R2372 VSS.n598 VSS.n597 71.676
R2373 VSS.n470 VSS.n468 71.676
R2374 VSS.n605 VSS.n604 71.676
R2375 VSS.n467 VSS.n465 71.676
R2376 VSS.n612 VSS.n611 71.676
R2377 VSS.n464 VSS.n462 71.676
R2378 VSS.n619 VSS.n618 71.676
R2379 VSS.n461 VSS.n457 71.676
R2380 VSS.n627 VSS.n626 71.676
R2381 VSS.n456 VSS.n454 71.676
R2382 VSS.n634 VSS.n633 71.676
R2383 VSS.n453 VSS.n451 71.676
R2384 VSS.n641 VSS.n640 71.676
R2385 VSS.n450 VSS.n448 71.676
R2386 VSS.n648 VSS.n647 71.676
R2387 VSS.n447 VSS.n445 71.676
R2388 VSS.n655 VSS.n654 71.676
R2389 VSS.n444 VSS.n442 71.676
R2390 VSS.n662 VSS.n661 71.676
R2391 VSS.n441 VSS.n439 71.676
R2392 VSS.n669 VSS.n668 71.676
R2393 VSS.n438 VSS.n436 71.676
R2394 VSS.n676 VSS.n675 71.676
R2395 VSS.n435 VSS.n433 71.676
R2396 VSS.n683 VSS.n682 71.676
R2397 VSS.n432 VSS.n430 71.676
R2398 VSS.n690 VSS.n689 71.676
R2399 VSS.n429 VSS.n427 71.676
R2400 VSS.n697 VSS.n696 71.676
R2401 VSS.n426 VSS.n424 71.676
R2402 VSS.n704 VSS.n703 71.676
R2403 VSS.n423 VSS.n421 71.676
R2404 VSS.n711 VSS.n710 71.676
R2405 VSS.n420 VSS.n418 71.676
R2406 VSS.n718 VSS.n717 71.676
R2407 VSS.n417 VSS.n415 71.676
R2408 VSS.n725 VSS.n724 71.676
R2409 VSS.n414 VSS.n17 71.676
R2410 VSS.n117 VSS.n116 71.676
R2411 VSS.n119 VSS.n113 71.676
R2412 VSS.n126 VSS.n125 71.676
R2413 VSS.n127 VSS.n111 71.676
R2414 VSS.n134 VSS.n133 71.676
R2415 VSS.n135 VSS.n109 71.676
R2416 VSS.n142 VSS.n141 71.676
R2417 VSS.n143 VSS.n107 71.676
R2418 VSS.n150 VSS.n149 71.676
R2419 VSS.n151 VSS.n105 71.676
R2420 VSS.n158 VSS.n157 71.676
R2421 VSS.n159 VSS.n103 71.676
R2422 VSS.n166 VSS.n165 71.676
R2423 VSS.n167 VSS.n101 71.676
R2424 VSS.n174 VSS.n173 71.676
R2425 VSS.n175 VSS.n99 71.676
R2426 VSS.n182 VSS.n181 71.676
R2427 VSS.n183 VSS.n97 71.676
R2428 VSS.n190 VSS.n189 71.676
R2429 VSS.n191 VSS.n95 71.676
R2430 VSS.n198 VSS.n197 71.676
R2431 VSS.n199 VSS.n93 71.676
R2432 VSS.n206 VSS.n205 71.676
R2433 VSS.n207 VSS.n91 71.676
R2434 VSS.n214 VSS.n213 71.676
R2435 VSS.n215 VSS.n89 71.676
R2436 VSS.n222 VSS.n221 71.676
R2437 VSS.n223 VSS.n87 71.676
R2438 VSS.n230 VSS.n229 71.676
R2439 VSS.n231 VSS.n83 71.676
R2440 VSS.n239 VSS.n238 71.676
R2441 VSS.n240 VSS.n81 71.676
R2442 VSS.n247 VSS.n246 71.676
R2443 VSS.n248 VSS.n79 71.676
R2444 VSS.n255 VSS.n254 71.676
R2445 VSS.n256 VSS.n77 71.676
R2446 VSS.n263 VSS.n262 71.676
R2447 VSS.n264 VSS.n75 71.676
R2448 VSS.n271 VSS.n270 71.676
R2449 VSS.n272 VSS.n73 71.676
R2450 VSS.n279 VSS.n278 71.676
R2451 VSS.n280 VSS.n71 71.676
R2452 VSS.n287 VSS.n286 71.676
R2453 VSS.n288 VSS.n69 71.676
R2454 VSS.n295 VSS.n294 71.676
R2455 VSS.n296 VSS.n67 71.676
R2456 VSS.n303 VSS.n302 71.676
R2457 VSS.n304 VSS.n65 71.676
R2458 VSS.n311 VSS.n310 71.676
R2459 VSS.n312 VSS.n63 71.676
R2460 VSS.n319 VSS.n318 71.676
R2461 VSS.n320 VSS.n61 71.676
R2462 VSS.n327 VSS.n326 71.676
R2463 VSS.n328 VSS.n59 71.676
R2464 VSS.n335 VSS.n334 71.676
R2465 VSS.n336 VSS.n57 71.676
R2466 VSS.n343 VSS.n342 71.676
R2467 VSS.n344 VSS.n55 71.676
R2468 VSS.n351 VSS.n350 71.676
R2469 VSS.n352 VSS.n53 71.676
R2470 VSS.n359 VSS.n358 71.676
R2471 VSS.n362 VSS.n361 71.676
R2472 VSS.n459 VSS.t13 68.5183
R2473 VSS.n509 VSS.t10 68.5183
R2474 VSS.n50 VSS.t5 68.5183
R2475 VSS.n85 VSS.t2 68.5183
R2476 VSS.n622 VSS.n459 49.0672
R2477 VSS.n510 VSS.n509 49.0672
R2478 VSS.n370 VSS.n369 48.7162
R2479 VSS.n378 VSS.n35 48.7162
R2480 VSS.n388 VSS.n35 48.7162
R2481 VSS.n406 VSS.n22 48.7162
R2482 VSS.n407 VSS.n406 48.7162
R2483 VSS.n408 VSS.n407 48.7162
R2484 VSS.n732 VSS.n14 48.7162
R2485 VSS.t8 VSS.n14 43.8446
R2486 VSS.n378 VSS.t1 41.896
R2487 VSS.n398 VSS.t16 39.9474
R2488 VSS.t14 VSS.n397 35.0758
R2489 VSS.n51 VSS.n50 34.3278
R2490 VSS.n235 VSS.n85 34.3278
R2491 VSS.n729 VSS.n728 31.5526
R2492 VSS.n736 VSS.n735 31.5526
R2493 VSS.n373 VSS.n43 31.5526
R2494 VSS.n366 VSS.n364 31.5526
R2495 VSS.t18 VSS.n396 30.2042
R2496 VSS.t15 VSS.n387 28.2556
R2497 VSS.n387 VSS.t17 25.3327
R2498 VSS.n396 VSS.t17 23.384
R2499 VSS.n388 VSS.t15 20.4611
R2500 VSS.n372 VSS.n42 19.3944
R2501 VSS.n376 VSS.n42 19.3944
R2502 VSS.n376 VSS.n33 19.3944
R2503 VSS.n390 VSS.n33 19.3944
R2504 VSS.n390 VSS.n31 19.3944
R2505 VSS.n394 VSS.n31 19.3944
R2506 VSS.n394 VSS.n27 19.3944
R2507 VSS.n400 VSS.n27 19.3944
R2508 VSS.n400 VSS.n25 19.3944
R2509 VSS.n404 VSS.n25 19.3944
R2510 VSS.n404 VSS.n20 19.3944
R2511 VSS.n410 VSS.n20 19.3944
R2512 VSS.n410 VSS.n18 19.3944
R2513 VSS.n730 VSS.n18 19.3944
R2514 VSS.n367 VSS.n47 19.3944
R2515 VSS.n47 VSS.n39 19.3944
R2516 VSS.n381 VSS.n39 19.3944
R2517 VSS.n381 VSS.n37 19.3944
R2518 VSS.n385 VSS.n37 19.3944
R2519 VSS.n385 VSS.n2 19.3944
R2520 VSS.n746 VSS.n2 19.3944
R2521 VSS.n746 VSS.n745 19.3944
R2522 VSS.n745 VSS.n744 19.3944
R2523 VSS.n744 VSS.n6 19.3944
R2524 VSS.n740 VSS.n6 19.3944
R2525 VSS.n740 VSS.n739 19.3944
R2526 VSS.n739 VSS.n738 19.3944
R2527 VSS.n738 VSS.n11 19.3944
R2528 VSS.n397 VSS.t18 18.5125
R2529 VSS.n398 VSS.t14 13.6409
R2530 VSS.n459 VSS.n458 10.6672
R2531 VSS.n509 VSS.n508 10.6672
R2532 VSS.n50 VSS.n49 10.6672
R2533 VSS.n85 VSS.n84 10.6672
R2534 VSS.n728 VSS.n727 10.6151
R2535 VSS.n727 VSS.n413 10.6151
R2536 VSS.n722 VSS.n413 10.6151
R2537 VSS.n722 VSS.n721 10.6151
R2538 VSS.n721 VSS.n720 10.6151
R2539 VSS.n720 VSS.n416 10.6151
R2540 VSS.n715 VSS.n416 10.6151
R2541 VSS.n715 VSS.n714 10.6151
R2542 VSS.n714 VSS.n713 10.6151
R2543 VSS.n713 VSS.n419 10.6151
R2544 VSS.n708 VSS.n419 10.6151
R2545 VSS.n708 VSS.n707 10.6151
R2546 VSS.n707 VSS.n706 10.6151
R2547 VSS.n706 VSS.n422 10.6151
R2548 VSS.n701 VSS.n422 10.6151
R2549 VSS.n701 VSS.n700 10.6151
R2550 VSS.n700 VSS.n699 10.6151
R2551 VSS.n699 VSS.n425 10.6151
R2552 VSS.n694 VSS.n425 10.6151
R2553 VSS.n694 VSS.n693 10.6151
R2554 VSS.n693 VSS.n692 10.6151
R2555 VSS.n692 VSS.n428 10.6151
R2556 VSS.n687 VSS.n428 10.6151
R2557 VSS.n687 VSS.n686 10.6151
R2558 VSS.n686 VSS.n685 10.6151
R2559 VSS.n685 VSS.n431 10.6151
R2560 VSS.n680 VSS.n431 10.6151
R2561 VSS.n680 VSS.n679 10.6151
R2562 VSS.n679 VSS.n678 10.6151
R2563 VSS.n678 VSS.n434 10.6151
R2564 VSS.n673 VSS.n434 10.6151
R2565 VSS.n673 VSS.n672 10.6151
R2566 VSS.n672 VSS.n671 10.6151
R2567 VSS.n671 VSS.n437 10.6151
R2568 VSS.n666 VSS.n437 10.6151
R2569 VSS.n666 VSS.n665 10.6151
R2570 VSS.n665 VSS.n664 10.6151
R2571 VSS.n664 VSS.n440 10.6151
R2572 VSS.n659 VSS.n440 10.6151
R2573 VSS.n659 VSS.n658 10.6151
R2574 VSS.n658 VSS.n657 10.6151
R2575 VSS.n657 VSS.n443 10.6151
R2576 VSS.n652 VSS.n443 10.6151
R2577 VSS.n652 VSS.n651 10.6151
R2578 VSS.n651 VSS.n650 10.6151
R2579 VSS.n650 VSS.n446 10.6151
R2580 VSS.n645 VSS.n446 10.6151
R2581 VSS.n645 VSS.n644 10.6151
R2582 VSS.n644 VSS.n643 10.6151
R2583 VSS.n643 VSS.n449 10.6151
R2584 VSS.n638 VSS.n449 10.6151
R2585 VSS.n638 VSS.n637 10.6151
R2586 VSS.n637 VSS.n636 10.6151
R2587 VSS.n636 VSS.n452 10.6151
R2588 VSS.n631 VSS.n452 10.6151
R2589 VSS.n631 VSS.n630 10.6151
R2590 VSS.n630 VSS.n629 10.6151
R2591 VSS.n629 VSS.n455 10.6151
R2592 VSS.n624 VSS.n455 10.6151
R2593 VSS.n624 VSS.n623 10.6151
R2594 VSS.n621 VSS.n460 10.6151
R2595 VSS.n616 VSS.n460 10.6151
R2596 VSS.n616 VSS.n615 10.6151
R2597 VSS.n615 VSS.n614 10.6151
R2598 VSS.n614 VSS.n463 10.6151
R2599 VSS.n609 VSS.n463 10.6151
R2600 VSS.n609 VSS.n608 10.6151
R2601 VSS.n608 VSS.n607 10.6151
R2602 VSS.n607 VSS.n466 10.6151
R2603 VSS.n602 VSS.n466 10.6151
R2604 VSS.n602 VSS.n601 10.6151
R2605 VSS.n601 VSS.n600 10.6151
R2606 VSS.n600 VSS.n469 10.6151
R2607 VSS.n595 VSS.n469 10.6151
R2608 VSS.n595 VSS.n594 10.6151
R2609 VSS.n594 VSS.n593 10.6151
R2610 VSS.n593 VSS.n472 10.6151
R2611 VSS.n588 VSS.n472 10.6151
R2612 VSS.n588 VSS.n587 10.6151
R2613 VSS.n587 VSS.n586 10.6151
R2614 VSS.n586 VSS.n475 10.6151
R2615 VSS.n581 VSS.n475 10.6151
R2616 VSS.n581 VSS.n580 10.6151
R2617 VSS.n580 VSS.n579 10.6151
R2618 VSS.n579 VSS.n478 10.6151
R2619 VSS.n574 VSS.n478 10.6151
R2620 VSS.n574 VSS.n573 10.6151
R2621 VSS.n573 VSS.n572 10.6151
R2622 VSS.n572 VSS.n481 10.6151
R2623 VSS.n567 VSS.n481 10.6151
R2624 VSS.n567 VSS.n566 10.6151
R2625 VSS.n566 VSS.n565 10.6151
R2626 VSS.n565 VSS.n484 10.6151
R2627 VSS.n560 VSS.n484 10.6151
R2628 VSS.n560 VSS.n559 10.6151
R2629 VSS.n559 VSS.n558 10.6151
R2630 VSS.n558 VSS.n487 10.6151
R2631 VSS.n553 VSS.n487 10.6151
R2632 VSS.n553 VSS.n552 10.6151
R2633 VSS.n552 VSS.n551 10.6151
R2634 VSS.n551 VSS.n490 10.6151
R2635 VSS.n546 VSS.n490 10.6151
R2636 VSS.n546 VSS.n545 10.6151
R2637 VSS.n545 VSS.n544 10.6151
R2638 VSS.n544 VSS.n493 10.6151
R2639 VSS.n539 VSS.n493 10.6151
R2640 VSS.n539 VSS.n538 10.6151
R2641 VSS.n538 VSS.n537 10.6151
R2642 VSS.n537 VSS.n496 10.6151
R2643 VSS.n532 VSS.n496 10.6151
R2644 VSS.n532 VSS.n531 10.6151
R2645 VSS.n531 VSS.n530 10.6151
R2646 VSS.n530 VSS.n499 10.6151
R2647 VSS.n525 VSS.n499 10.6151
R2648 VSS.n525 VSS.n524 10.6151
R2649 VSS.n524 VSS.n523 10.6151
R2650 VSS.n523 VSS.n502 10.6151
R2651 VSS.n518 VSS.n502 10.6151
R2652 VSS.n518 VSS.n517 10.6151
R2653 VSS.n517 VSS.n516 10.6151
R2654 VSS.n516 VSS.n505 10.6151
R2655 VSS.n511 VSS.n12 10.6151
R2656 VSS.n735 VSS.n12 10.6151
R2657 VSS.n115 VSS.n43 10.6151
R2658 VSS.n115 VSS.n114 10.6151
R2659 VSS.n121 VSS.n114 10.6151
R2660 VSS.n122 VSS.n121 10.6151
R2661 VSS.n123 VSS.n122 10.6151
R2662 VSS.n123 VSS.n112 10.6151
R2663 VSS.n129 VSS.n112 10.6151
R2664 VSS.n130 VSS.n129 10.6151
R2665 VSS.n131 VSS.n130 10.6151
R2666 VSS.n131 VSS.n110 10.6151
R2667 VSS.n137 VSS.n110 10.6151
R2668 VSS.n138 VSS.n137 10.6151
R2669 VSS.n139 VSS.n138 10.6151
R2670 VSS.n139 VSS.n108 10.6151
R2671 VSS.n145 VSS.n108 10.6151
R2672 VSS.n146 VSS.n145 10.6151
R2673 VSS.n147 VSS.n146 10.6151
R2674 VSS.n147 VSS.n106 10.6151
R2675 VSS.n153 VSS.n106 10.6151
R2676 VSS.n154 VSS.n153 10.6151
R2677 VSS.n155 VSS.n154 10.6151
R2678 VSS.n155 VSS.n104 10.6151
R2679 VSS.n161 VSS.n104 10.6151
R2680 VSS.n162 VSS.n161 10.6151
R2681 VSS.n163 VSS.n162 10.6151
R2682 VSS.n163 VSS.n102 10.6151
R2683 VSS.n169 VSS.n102 10.6151
R2684 VSS.n170 VSS.n169 10.6151
R2685 VSS.n171 VSS.n170 10.6151
R2686 VSS.n171 VSS.n100 10.6151
R2687 VSS.n177 VSS.n100 10.6151
R2688 VSS.n178 VSS.n177 10.6151
R2689 VSS.n179 VSS.n178 10.6151
R2690 VSS.n179 VSS.n98 10.6151
R2691 VSS.n185 VSS.n98 10.6151
R2692 VSS.n186 VSS.n185 10.6151
R2693 VSS.n187 VSS.n186 10.6151
R2694 VSS.n187 VSS.n96 10.6151
R2695 VSS.n193 VSS.n96 10.6151
R2696 VSS.n194 VSS.n193 10.6151
R2697 VSS.n195 VSS.n194 10.6151
R2698 VSS.n195 VSS.n94 10.6151
R2699 VSS.n201 VSS.n94 10.6151
R2700 VSS.n202 VSS.n201 10.6151
R2701 VSS.n203 VSS.n202 10.6151
R2702 VSS.n203 VSS.n92 10.6151
R2703 VSS.n209 VSS.n92 10.6151
R2704 VSS.n210 VSS.n209 10.6151
R2705 VSS.n211 VSS.n210 10.6151
R2706 VSS.n211 VSS.n90 10.6151
R2707 VSS.n217 VSS.n90 10.6151
R2708 VSS.n218 VSS.n217 10.6151
R2709 VSS.n219 VSS.n218 10.6151
R2710 VSS.n219 VSS.n88 10.6151
R2711 VSS.n225 VSS.n88 10.6151
R2712 VSS.n226 VSS.n225 10.6151
R2713 VSS.n227 VSS.n226 10.6151
R2714 VSS.n227 VSS.n86 10.6151
R2715 VSS.n233 VSS.n86 10.6151
R2716 VSS.n234 VSS.n233 10.6151
R2717 VSS.n236 VSS.n82 10.6151
R2718 VSS.n242 VSS.n82 10.6151
R2719 VSS.n243 VSS.n242 10.6151
R2720 VSS.n244 VSS.n243 10.6151
R2721 VSS.n244 VSS.n80 10.6151
R2722 VSS.n250 VSS.n80 10.6151
R2723 VSS.n251 VSS.n250 10.6151
R2724 VSS.n252 VSS.n251 10.6151
R2725 VSS.n252 VSS.n78 10.6151
R2726 VSS.n258 VSS.n78 10.6151
R2727 VSS.n259 VSS.n258 10.6151
R2728 VSS.n260 VSS.n259 10.6151
R2729 VSS.n260 VSS.n76 10.6151
R2730 VSS.n266 VSS.n76 10.6151
R2731 VSS.n267 VSS.n266 10.6151
R2732 VSS.n268 VSS.n267 10.6151
R2733 VSS.n268 VSS.n74 10.6151
R2734 VSS.n274 VSS.n74 10.6151
R2735 VSS.n275 VSS.n274 10.6151
R2736 VSS.n276 VSS.n275 10.6151
R2737 VSS.n276 VSS.n72 10.6151
R2738 VSS.n282 VSS.n72 10.6151
R2739 VSS.n283 VSS.n282 10.6151
R2740 VSS.n284 VSS.n283 10.6151
R2741 VSS.n284 VSS.n70 10.6151
R2742 VSS.n290 VSS.n70 10.6151
R2743 VSS.n291 VSS.n290 10.6151
R2744 VSS.n292 VSS.n291 10.6151
R2745 VSS.n292 VSS.n68 10.6151
R2746 VSS.n298 VSS.n68 10.6151
R2747 VSS.n299 VSS.n298 10.6151
R2748 VSS.n300 VSS.n299 10.6151
R2749 VSS.n300 VSS.n66 10.6151
R2750 VSS.n306 VSS.n66 10.6151
R2751 VSS.n307 VSS.n306 10.6151
R2752 VSS.n308 VSS.n307 10.6151
R2753 VSS.n308 VSS.n64 10.6151
R2754 VSS.n314 VSS.n64 10.6151
R2755 VSS.n315 VSS.n314 10.6151
R2756 VSS.n316 VSS.n315 10.6151
R2757 VSS.n316 VSS.n62 10.6151
R2758 VSS.n322 VSS.n62 10.6151
R2759 VSS.n323 VSS.n322 10.6151
R2760 VSS.n324 VSS.n323 10.6151
R2761 VSS.n324 VSS.n60 10.6151
R2762 VSS.n330 VSS.n60 10.6151
R2763 VSS.n331 VSS.n330 10.6151
R2764 VSS.n332 VSS.n331 10.6151
R2765 VSS.n332 VSS.n58 10.6151
R2766 VSS.n338 VSS.n58 10.6151
R2767 VSS.n339 VSS.n338 10.6151
R2768 VSS.n340 VSS.n339 10.6151
R2769 VSS.n340 VSS.n56 10.6151
R2770 VSS.n346 VSS.n56 10.6151
R2771 VSS.n347 VSS.n346 10.6151
R2772 VSS.n348 VSS.n347 10.6151
R2773 VSS.n348 VSS.n54 10.6151
R2774 VSS.n354 VSS.n54 10.6151
R2775 VSS.n355 VSS.n354 10.6151
R2776 VSS.n356 VSS.n355 10.6151
R2777 VSS.n356 VSS.n52 10.6151
R2778 VSS.n363 VSS.n48 10.6151
R2779 VSS.n364 VSS.n363 10.6151
R2780 VSS.n622 VSS.n621 9.99074
R2781 VSS.n510 VSS.n505 9.99074
R2782 VSS.n236 VSS.n235 9.99074
R2783 VSS.n52 VSS.n51 9.99074
R2784 VSS.n745 VSS.n0 9.3005
R2785 VSS.n744 VSS.n743 9.3005
R2786 VSS.n742 VSS.n6 9.3005
R2787 VSS.n741 VSS.n740 9.3005
R2788 VSS.n739 VSS.n7 9.3005
R2789 VSS.n738 VSS.n737 9.3005
R2790 VSS.n736 VSS.n11 9.3005
R2791 VSS.n373 VSS.n372 9.3005
R2792 VSS.n374 VSS.n42 9.3005
R2793 VSS.n376 VSS.n375 9.3005
R2794 VSS.n33 VSS.n32 9.3005
R2795 VSS.n391 VSS.n390 9.3005
R2796 VSS.n392 VSS.n31 9.3005
R2797 VSS.n394 VSS.n393 9.3005
R2798 VSS.n27 VSS.n26 9.3005
R2799 VSS.n401 VSS.n400 9.3005
R2800 VSS.n402 VSS.n25 9.3005
R2801 VSS.n404 VSS.n403 9.3005
R2802 VSS.n20 VSS.n19 9.3005
R2803 VSS.n411 VSS.n410 9.3005
R2804 VSS.n412 VSS.n18 9.3005
R2805 VSS.n730 VSS.n729 9.3005
R2806 VSS.n365 VSS.n47 9.3005
R2807 VSS.n39 VSS.n38 9.3005
R2808 VSS.n382 VSS.n381 9.3005
R2809 VSS.n383 VSS.n37 9.3005
R2810 VSS.n385 VSS.n384 9.3005
R2811 VSS.n2 VSS.n1 9.3005
R2812 VSS.n367 VSS.n366 9.3005
R2813 VSS.n747 VSS.n746 9.3005
R2814 VSS.t16 VSS.n22 8.76932
R2815 VSS.n369 VSS.t1 6.82069
R2816 VSS.n408 VSS.t8 4.87207
R2817 VSS.n623 VSS.n622 0.62489
R2818 VSS.n511 VSS.n510 0.62489
R2819 VSS.n235 VSS.n234 0.62489
R2820 VSS.n51 VSS.n48 0.62489
R2821 VSS.n743 VSS.n0 0.152939
R2822 VSS.n743 VSS.n742 0.152939
R2823 VSS.n742 VSS.n741 0.152939
R2824 VSS.n741 VSS.n7 0.152939
R2825 VSS.n737 VSS.n7 0.152939
R2826 VSS.n737 VSS.n736 0.152939
R2827 VSS.n374 VSS.n373 0.152939
R2828 VSS.n375 VSS.n374 0.152939
R2829 VSS.n375 VSS.n32 0.152939
R2830 VSS.n391 VSS.n32 0.152939
R2831 VSS.n392 VSS.n391 0.152939
R2832 VSS.n393 VSS.n392 0.152939
R2833 VSS.n393 VSS.n26 0.152939
R2834 VSS.n401 VSS.n26 0.152939
R2835 VSS.n402 VSS.n401 0.152939
R2836 VSS.n403 VSS.n402 0.152939
R2837 VSS.n403 VSS.n19 0.152939
R2838 VSS.n411 VSS.n19 0.152939
R2839 VSS.n412 VSS.n411 0.152939
R2840 VSS.n729 VSS.n412 0.152939
R2841 VSS.n366 VSS.n365 0.152939
R2842 VSS.n365 VSS.n38 0.152939
R2843 VSS.n382 VSS.n38 0.152939
R2844 VSS.n383 VSS.n382 0.152939
R2845 VSS.n384 VSS.n383 0.152939
R2846 VSS.n384 VSS.n1 0.152939
R2847 VSS.n747 VSS.n1 0.13922
R2848 VSS VSS.n0 0.0767195
R2849 VSS VSS.n747 0.063
C0 VOUT VGN 8.88414f
C1 VOUT VCC 20.099401f
C2 VGN VCC 0.003903f
C3 VGN VSS 4.586157f
C4 VOUT VSS 20.31851f
C5 VGP VSS 0.05975f
C6 VIN VSS 0.223745f
C7 VCC VSS 97.852844f
C8 VGN.n0 VSS 0.043269f
C9 VGN.t8 VSS 0.516948f
C10 VGN.t5 VSS 0.512552f
C11 VGN.t4 VSS 0.512552f
C12 VGN.t3 VSS 0.512552f
C13 VGN.n1 VSS 0.194919f
C14 VGN.t2 VSS 0.516948f
C15 VGN.n2 VSS 0.208141f
C16 VGN.n3 VSS 0.097677f
C17 VGN.n4 VSS 0.015687f
C18 VGN.n5 VSS 0.194919f
C19 VGN.n6 VSS 0.015687f
C20 VGN.n7 VSS 0.194919f
C21 VGN.n8 VSS 0.208077f
C22 VGN.n9 VSS 0.700561f
C23 VGN.n10 VSS 0.043269f
C24 VGN.t0 VSS 0.516948f
C25 VGN.t6 VSS 0.512552f
C26 VGN.t1 VSS 0.512552f
C27 VGN.t9 VSS 0.512552f
C28 VGN.n11 VSS 0.194919f
C29 VGN.t7 VSS 0.516948f
C30 VGN.n12 VSS 0.208141f
C31 VGN.n13 VSS 0.097677f
C32 VGN.n14 VSS 0.015687f
C33 VGN.n15 VSS 0.194919f
C34 VGN.n16 VSS 0.015687f
C35 VGN.n17 VSS 0.194919f
C36 VGN.n18 VSS 0.208077f
C37 VGN.n19 VSS 0.0386f
C38 VOUT.t27 VSS 0.854948f
C39 VOUT.n0 VSS 0.345163f
C40 VOUT.n1 VSS 0.010036f
C41 VOUT.n2 VSS 0.013062f
C42 VOUT.n3 VSS 0.010036f
C43 VOUT.n4 VSS 0.011812f
C44 VOUT.n5 VSS 0.010036f
C45 VOUT.t29 VSS 0.854948f
C46 VOUT.n6 VSS 0.305234f
C47 VOUT.n7 VSS 0.00866f
C48 VOUT.n8 VSS 0.010036f
C49 VOUT.t19 VSS 0.854948f
C50 VOUT.n9 VSS 0.314657f
C51 VOUT.n10 VSS 0.010036f
C52 VOUT.n11 VSS 0.00866f
C53 VOUT.n12 VSS 0.010036f
C54 VOUT.t21 VSS 0.854948f
C55 VOUT.n13 VSS 0.3421f
C56 VOUT.t16 VSS 0.990984f
C57 VOUT.n14 VSS 0.32217f
C58 VOUT.n15 VSS 0.124063f
C59 VOUT.n16 VSS 0.016222f
C60 VOUT.n17 VSS 0.018611f
C61 VOUT.n18 VSS 0.020169f
C62 VOUT.n19 VSS 0.010036f
C63 VOUT.n20 VSS 0.010036f
C64 VOUT.n21 VSS 0.010036f
C65 VOUT.n22 VSS 0.018961f
C66 VOUT.n23 VSS 0.018611f
C67 VOUT.n24 VSS 0.018611f
C68 VOUT.n25 VSS 0.010036f
C69 VOUT.n26 VSS 0.010036f
C70 VOUT.n27 VSS 0.010036f
C71 VOUT.n28 VSS 0.018611f
C72 VOUT.n29 VSS 0.018611f
C73 VOUT.n30 VSS 0.018961f
C74 VOUT.n31 VSS 0.010036f
C75 VOUT.n32 VSS 0.010036f
C76 VOUT.n33 VSS 0.010036f
C77 VOUT.n34 VSS 0.020169f
C78 VOUT.n35 VSS 0.018611f
C79 VOUT.n36 VSS 0.016222f
C80 VOUT.n37 VSS 0.010036f
C81 VOUT.n38 VSS 0.010036f
C82 VOUT.n39 VSS 0.010036f
C83 VOUT.n40 VSS 0.018611f
C84 VOUT.n41 VSS 0.018611f
C85 VOUT.n42 VSS 0.016117f
C86 VOUT.n43 VSS 0.010036f
C87 VOUT.n44 VSS 0.010036f
C88 VOUT.n45 VSS 0.010036f
C89 VOUT.n46 VSS 0.018611f
C90 VOUT.n47 VSS 0.018611f
C91 VOUT.n48 VSS 0.013834f
C92 VOUT.n49 VSS 0.016196f
C93 VOUT.n50 VSS 0.05974f
C94 VOUT.n51 VSS 0.286759f
C95 VOUT.n52 VSS 0.049f
C96 VOUT.t5 VSS 0.751521f
C97 VOUT.n53 VSS 0.092271f
C98 VOUT.n54 VSS 0.090805f
C99 VOUT.n55 VSS 0.194518f
C100 VOUT.t20 VSS 0.055195f
C101 VOUT.t28 VSS 0.300639f
C102 VOUT.t30 VSS 0.055195f
C103 VOUT.n56 VSS 0.204002f
C104 VOUT.n57 VSS 0.271177f
C105 VOUT.n58 VSS 0.271177f
C106 VOUT.t13 VSS 0.055195f
C107 VOUT.t23 VSS 0.854948f
C108 VOUT.n59 VSS 0.345163f
C109 VOUT.n60 VSS 0.010036f
C110 VOUT.n61 VSS 0.013062f
C111 VOUT.n62 VSS 0.010036f
C112 VOUT.n63 VSS 0.011812f
C113 VOUT.n64 VSS 0.010036f
C114 VOUT.t25 VSS 0.854948f
C115 VOUT.n65 VSS 0.305234f
C116 VOUT.n66 VSS 0.00866f
C117 VOUT.n67 VSS 0.010036f
C118 VOUT.t12 VSS 0.854948f
C119 VOUT.n68 VSS 0.314657f
C120 VOUT.n69 VSS 0.010036f
C121 VOUT.n70 VSS 0.00866f
C122 VOUT.n71 VSS 0.010036f
C123 VOUT.t14 VSS 0.854948f
C124 VOUT.n72 VSS 0.3421f
C125 VOUT.t31 VSS 0.990985f
C126 VOUT.n73 VSS 0.322169f
C127 VOUT.n74 VSS 0.124063f
C128 VOUT.n75 VSS 0.016222f
C129 VOUT.n76 VSS 0.018611f
C130 VOUT.n77 VSS 0.020169f
C131 VOUT.n78 VSS 0.010036f
C132 VOUT.n79 VSS 0.010036f
C133 VOUT.n80 VSS 0.010036f
C134 VOUT.n81 VSS 0.018961f
C135 VOUT.n82 VSS 0.018611f
C136 VOUT.n83 VSS 0.018611f
C137 VOUT.n84 VSS 0.010036f
C138 VOUT.n85 VSS 0.010036f
C139 VOUT.n86 VSS 0.010036f
C140 VOUT.n87 VSS 0.018611f
C141 VOUT.n88 VSS 0.018611f
C142 VOUT.n89 VSS 0.018961f
C143 VOUT.n90 VSS 0.010036f
C144 VOUT.n91 VSS 0.010036f
C145 VOUT.n92 VSS 0.010036f
C146 VOUT.n93 VSS 0.020169f
C147 VOUT.n94 VSS 0.018611f
C148 VOUT.n95 VSS 0.016222f
C149 VOUT.n96 VSS 0.010036f
C150 VOUT.n97 VSS 0.010036f
C151 VOUT.n98 VSS 0.010036f
C152 VOUT.n99 VSS 0.018611f
C153 VOUT.n100 VSS 0.018611f
C154 VOUT.n101 VSS 0.016117f
C155 VOUT.n102 VSS 0.010036f
C156 VOUT.n103 VSS 0.010036f
C157 VOUT.n104 VSS 0.010036f
C158 VOUT.n105 VSS 0.018611f
C159 VOUT.n106 VSS 0.018611f
C160 VOUT.n107 VSS 0.013834f
C161 VOUT.n108 VSS 0.016196f
C162 VOUT.n109 VSS 0.031191f
C163 VOUT.n110 VSS 0.12105f
C164 VOUT.t24 VSS 0.300639f
C165 VOUT.n111 VSS 0.204002f
C166 VOUT.t26 VSS 0.055195f
C167 VOUT.n112 VSS 0.186192f
C168 VOUT.n113 VSS 0.169704f
C169 VOUT.t33 VSS 0.248766f
C170 VOUT.n114 VSS 0.150374f
C171 VOUT.n115 VSS 0.16522f
C172 VOUT.n116 VSS 0.186192f
C173 VOUT.t15 VSS 0.055195f
C174 VOUT.t32 VSS 0.027598f
C175 VOUT.n117 VSS 0.204002f
C176 VOUT.n118 VSS 0.133209f
C177 VOUT.n119 VSS 0.103102f
C178 VOUT.n120 VSS 0.232752f
C179 VOUT.t17 VSS 0.027598f
C180 VOUT.n121 VSS 0.204002f
C181 VOUT.t22 VSS 0.055195f
C182 VOUT.n122 VSS 0.186192f
C183 VOUT.n123 VSS 0.32369f
C184 VOUT.t18 VSS 0.248766f
C185 VOUT.n124 VSS 0.150071f
C186 VOUT.n125 VSS 0.280817f
C187 VOUT.n126 VSS 0.092271f
C188 VOUT.t6 VSS 0.118248f
C189 VOUT.t7 VSS 0.751521f
C190 VOUT.n127 VSS 0.541178f
C191 VOUT.t0 VSS 0.118248f
C192 VOUT.n128 VSS 0.530691f
C193 VOUT.t11 VSS 0.677627f
C194 VOUT.n129 VSS 0.192711f
C195 VOUT.t3 VSS 0.677627f
C196 VOUT.n130 VSS 0.192711f
C197 VOUT.n131 VSS 0.099065f
C198 VOUT.n132 VSS 0.53018f
C199 VOUT.t1 VSS 0.118248f
C200 VOUT.t2 VSS 0.059124f
C201 VOUT.n133 VSS 0.541178f
C202 VOUT.n134 VSS 0.183977f
C203 VOUT.n135 VSS 0.303821f
C204 VOUT.n136 VSS 0.05175f
C205 VOUT.t10 VSS 0.059124f
C206 VOUT.n137 VSS 0.541178f
C207 VOUT.t9 VSS 0.118248f
C208 VOUT.n138 VSS 0.53018f
C209 VOUT.t4 VSS 0.118248f
C210 VOUT.n139 VSS 0.541178f
C211 VOUT.t8 VSS 0.118248f
C212 VOUT.n140 VSS 0.53018f
C213 VOUT.n141 VSS 0.046063f
C214 VCC.n0 VSS 0.003824f
C215 VCC.n1 VSS 0.004244f
C216 VCC.n2 VSS 0.003078f
C217 VCC.n3 VSS 0.003824f
C218 VCC.n4 VSS 0.003824f
C219 VCC.n5 VSS 0.003824f
C220 VCC.n6 VSS 0.003078f
C221 VCC.n7 VSS 0.003824f
C222 VCC.n8 VSS 0.003824f
C223 VCC.n9 VSS 0.003824f
C224 VCC.n10 VSS 0.003824f
C225 VCC.n11 VSS 0.003078f
C226 VCC.n12 VSS 0.003824f
C227 VCC.n13 VSS 0.003824f
C228 VCC.n14 VSS 0.003824f
C229 VCC.n15 VSS 0.003824f
C230 VCC.n16 VSS 0.003078f
C231 VCC.n17 VSS 0.003824f
C232 VCC.n18 VSS 0.003824f
C233 VCC.n19 VSS 0.003824f
C234 VCC.n20 VSS 0.003824f
C235 VCC.n21 VSS 0.003078f
C236 VCC.n22 VSS 0.003824f
C237 VCC.n23 VSS 0.003824f
C238 VCC.n24 VSS 0.003824f
C239 VCC.n25 VSS 0.003824f
C240 VCC.n26 VSS 0.003078f
C241 VCC.n27 VSS 0.003824f
C242 VCC.n28 VSS 0.003824f
C243 VCC.n29 VSS 0.003824f
C244 VCC.n30 VSS 0.003824f
C245 VCC.n31 VSS 0.003078f
C246 VCC.n32 VSS 0.003824f
C247 VCC.n33 VSS 0.003824f
C248 VCC.n34 VSS 0.003824f
C249 VCC.n35 VSS 0.003824f
C250 VCC.n36 VSS 0.003078f
C251 VCC.n37 VSS 0.012377f
C252 VCC.n38 VSS 0.003824f
C253 VCC.n39 VSS 0.007052f
C254 VCC.n40 VSS 0.226571f
C255 VCC.n41 VSS 0.42482f
C256 VCC.n42 VSS 0.003824f
C257 VCC.n43 VSS 0.007052f
C258 VCC.n44 VSS 0.003078f
C259 VCC.n45 VSS 0.003824f
C260 VCC.n46 VSS 0.003078f
C261 VCC.n47 VSS 0.003824f
C262 VCC.t6 VSS 0.113285f
C263 VCC.n48 VSS 0.003824f
C264 VCC.n49 VSS 0.003078f
C265 VCC.n50 VSS 0.003824f
C266 VCC.n51 VSS 0.003078f
C267 VCC.n52 VSS 0.003824f
C268 VCC.n53 VSS 0.226571f
C269 VCC.n54 VSS 0.003824f
C270 VCC.n55 VSS 0.003078f
C271 VCC.n56 VSS 0.003824f
C272 VCC.n57 VSS 0.003078f
C273 VCC.n58 VSS 0.003824f
C274 VCC.n59 VSS 0.226571f
C275 VCC.n60 VSS 0.003824f
C276 VCC.n61 VSS 0.003078f
C277 VCC.n62 VSS 0.003824f
C278 VCC.n63 VSS 0.003078f
C279 VCC.n64 VSS 0.003824f
C280 VCC.n65 VSS 0.226571f
C281 VCC.n66 VSS 0.003824f
C282 VCC.n67 VSS 0.003078f
C283 VCC.n68 VSS 0.003824f
C284 VCC.n69 VSS 0.003078f
C285 VCC.n70 VSS 0.003824f
C286 VCC.n71 VSS 0.199382f
C287 VCC.n72 VSS 0.003824f
C288 VCC.n73 VSS 0.003078f
C289 VCC.n74 VSS 0.003824f
C290 VCC.n75 VSS 0.003078f
C291 VCC.n76 VSS 0.003824f
C292 VCC.n77 VSS 0.226571f
C293 VCC.n78 VSS 0.003824f
C294 VCC.n79 VSS 0.003078f
C295 VCC.n80 VSS 0.003824f
C296 VCC.n81 VSS 0.003078f
C297 VCC.n82 VSS 0.003824f
C298 VCC.n83 VSS 0.169928f
C299 VCC.n84 VSS 0.003824f
C300 VCC.n85 VSS 0.003078f
C301 VCC.n86 VSS 0.003824f
C302 VCC.n87 VSS 0.003078f
C303 VCC.n88 VSS 0.003824f
C304 VCC.n89 VSS 0.226571f
C305 VCC.t2 VSS 0.113285f
C306 VCC.n90 VSS 0.003824f
C307 VCC.n91 VSS 0.003078f
C308 VCC.n92 VSS 0.003824f
C309 VCC.n93 VSS 0.003078f
C310 VCC.n94 VSS 0.003824f
C311 VCC.n95 VSS 0.226571f
C312 VCC.n96 VSS 0.003824f
C313 VCC.n97 VSS 0.003078f
C314 VCC.n98 VSS 0.003824f
C315 VCC.n99 VSS 0.003078f
C316 VCC.n100 VSS 0.003824f
C317 VCC.n101 VSS 0.226571f
C318 VCC.n102 VSS 0.003824f
C319 VCC.n103 VSS 0.003078f
C320 VCC.n104 VSS 0.003824f
C321 VCC.n105 VSS 0.003078f
C322 VCC.n106 VSS 0.003824f
C323 VCC.t0 VSS 0.113285f
C324 VCC.n107 VSS 0.003824f
C325 VCC.n108 VSS 0.003078f
C326 VCC.n109 VSS 0.003078f
C327 VCC.n110 VSS 0.003824f
C328 VCC.n111 VSS 0.003078f
C329 VCC.n112 VSS 0.003824f
C330 VCC.n113 VSS 0.226571f
C331 VCC.n114 VSS 0.199382f
C332 VCC.n115 VSS 0.003824f
C333 VCC.n116 VSS 0.003078f
C334 VCC.n117 VSS 0.003824f
C335 VCC.n118 VSS 0.003078f
C336 VCC.n119 VSS 0.003824f
C337 VCC.n120 VSS 0.226571f
C338 VCC.n121 VSS 0.003824f
C339 VCC.n122 VSS 0.003078f
C340 VCC.n123 VSS 0.003824f
C341 VCC.n124 VSS 0.003078f
C342 VCC.n125 VSS 0.003824f
C343 VCC.n126 VSS 0.224305f
C344 VCC.n127 VSS 0.003824f
C345 VCC.n128 VSS 0.003078f
C346 VCC.n129 VSS 0.003824f
C347 VCC.n130 VSS 0.003078f
C348 VCC.n131 VSS 0.003824f
C349 VCC.n132 VSS 0.226571f
C350 VCC.n133 VSS 0.003824f
C351 VCC.n134 VSS 0.003078f
C352 VCC.n135 VSS 0.003824f
C353 VCC.n136 VSS 0.003078f
C354 VCC.n137 VSS 0.003824f
C355 VCC.n138 VSS 0.226571f
C356 VCC.n139 VSS 0.003824f
C357 VCC.n140 VSS 0.003078f
C358 VCC.n141 VSS 0.003824f
C359 VCC.n142 VSS 0.003078f
C360 VCC.n143 VSS 0.003824f
C361 VCC.n144 VSS 0.226571f
C362 VCC.n145 VSS 0.003824f
C363 VCC.n146 VSS 0.003078f
C364 VCC.n147 VSS 0.003824f
C365 VCC.n148 VSS 0.003078f
C366 VCC.n149 VSS 0.003824f
C367 VCC.n150 VSS 0.226571f
C368 VCC.n151 VSS 0.003824f
C369 VCC.n152 VSS 0.003078f
C370 VCC.n153 VSS 0.003824f
C371 VCC.n154 VSS 0.003078f
C372 VCC.n155 VSS 0.003824f
C373 VCC.n156 VSS 0.215242f
C374 VCC.n157 VSS 0.003824f
C375 VCC.n158 VSS 0.003078f
C376 VCC.n159 VSS 0.003824f
C377 VCC.n160 VSS 0.003078f
C378 VCC.n161 VSS 0.003824f
C379 VCC.n162 VSS 0.226571f
C380 VCC.t10 VSS 0.113285f
C381 VCC.n163 VSS 0.003824f
C382 VCC.n164 VSS 0.003078f
C383 VCC.n165 VSS 0.003824f
C384 VCC.n166 VSS 0.003078f
C385 VCC.n167 VSS 0.003824f
C386 VCC.n168 VSS 0.226571f
C387 VCC.n169 VSS 0.003824f
C388 VCC.n170 VSS 0.003078f
C389 VCC.n171 VSS 0.004871f
C390 VCC.n172 VSS 0.007052f
C391 VCC.n173 VSS 0.42482f
C392 VCC.n174 VSS 0.007052f
C393 VCC.n175 VSS 0.001358f
C394 VCC.t11 VSS 0.104021f
C395 VCC.t12 VSS 0.113895f
C396 VCC.t9 VSS 0.55312f
C397 VCC.n177 VSS 0.064333f
C398 VCC.n178 VSS 0.025611f
C399 VCC.n179 VSS 0.003624f
C400 VCC.n180 VSS 0.002601f
C401 VCC.n181 VSS 0.002601f
C402 VCC.n182 VSS 0.002601f
C403 VCC.n183 VSS 0.002601f
C404 VCC.n184 VSS 0.002601f
C405 VCC.n185 VSS 0.002601f
C406 VCC.n186 VSS 0.002601f
C407 VCC.n187 VSS 0.002601f
C408 VCC.n188 VSS 0.002601f
C409 VCC.n189 VSS 0.002601f
C410 VCC.n190 VSS 0.002601f
C411 VCC.n191 VSS 0.002601f
C412 VCC.n192 VSS 0.002601f
C413 VCC.n193 VSS 0.002601f
C414 VCC.n194 VSS 0.002601f
C415 VCC.n195 VSS 0.002601f
C416 VCC.t14 VSS 0.104021f
C417 VCC.t15 VSS 0.113895f
C418 VCC.t13 VSS 0.55312f
C419 VCC.n196 VSS 0.064333f
C420 VCC.n197 VSS 0.025611f
C421 VCC.n198 VSS 0.002601f
C422 VCC.n199 VSS 0.002601f
C423 VCC.n200 VSS 0.002601f
C424 VCC.n201 VSS 0.002601f
C425 VCC.n202 VSS 0.002601f
C426 VCC.n203 VSS 0.002601f
C427 VCC.n204 VSS 0.002601f
C428 VCC.n205 VSS 0.002601f
C429 VCC.n206 VSS 0.002601f
C430 VCC.n207 VSS 0.002601f
C431 VCC.n208 VSS 0.002601f
C432 VCC.n209 VSS 0.002601f
C433 VCC.n210 VSS 0.002601f
C434 VCC.n211 VSS 0.002601f
C435 VCC.n213 VSS 0.002601f
C436 VCC.n214 VSS 0.002601f
C437 VCC.n215 VSS 0.002601f
C438 VCC.n216 VSS 0.002601f
C439 VCC.n217 VSS 0.002601f
C440 VCC.n219 VSS 0.002601f
C441 VCC.n221 VSS 0.002601f
C442 VCC.n222 VSS 0.002601f
C443 VCC.n223 VSS 0.002601f
C444 VCC.n224 VSS 0.002601f
C445 VCC.n225 VSS 0.002601f
C446 VCC.n227 VSS 0.002601f
C447 VCC.n229 VSS 0.002601f
C448 VCC.n230 VSS 0.002601f
C449 VCC.n231 VSS 0.002601f
C450 VCC.n232 VSS 0.002601f
C451 VCC.n233 VSS 0.002601f
C452 VCC.n235 VSS 0.002601f
C453 VCC.n237 VSS 0.002601f
C454 VCC.n238 VSS 0.002601f
C455 VCC.n239 VSS 0.002601f
C456 VCC.n240 VSS 0.002601f
C457 VCC.n241 VSS 0.002601f
C458 VCC.n243 VSS 0.002601f
C459 VCC.n245 VSS 0.002601f
C460 VCC.n246 VSS 0.002601f
C461 VCC.n247 VSS 0.002601f
C462 VCC.n248 VSS 0.002601f
C463 VCC.n249 VSS 0.002601f
C464 VCC.n251 VSS 0.002601f
C465 VCC.n253 VSS 0.002601f
C466 VCC.n254 VSS 0.002601f
C467 VCC.n255 VSS 0.002601f
C468 VCC.n256 VSS 0.002601f
C469 VCC.n257 VSS 0.002601f
C470 VCC.n259 VSS 0.002601f
C471 VCC.n261 VSS 0.002601f
C472 VCC.n262 VSS 0.002601f
C473 VCC.n263 VSS 0.002601f
C474 VCC.n264 VSS 0.002601f
C475 VCC.n265 VSS 0.002601f
C476 VCC.n267 VSS 0.002601f
C477 VCC.n269 VSS 0.002601f
C478 VCC.n270 VSS 0.002601f
C479 VCC.n271 VSS 0.001396f
C480 VCC.n272 VSS 0.003624f
C481 VCC.n273 VSS 0.002505f
C482 VCC.n274 VSS 0.002601f
C483 VCC.n276 VSS 0.002601f
C484 VCC.n278 VSS 0.002601f
C485 VCC.n279 VSS 0.002601f
C486 VCC.n280 VSS 0.002601f
C487 VCC.n281 VSS 0.002601f
C488 VCC.n282 VSS 0.002601f
C489 VCC.n284 VSS 0.002601f
C490 VCC.n286 VSS 0.002601f
C491 VCC.n287 VSS 0.002601f
C492 VCC.n288 VSS 0.002601f
C493 VCC.n289 VSS 0.002601f
C494 VCC.n290 VSS 0.002601f
C495 VCC.n292 VSS 0.002601f
C496 VCC.n294 VSS 0.002601f
C497 VCC.n295 VSS 0.002601f
C498 VCC.n296 VSS 0.002601f
C499 VCC.n297 VSS 0.002601f
C500 VCC.n298 VSS 0.002601f
C501 VCC.n300 VSS 0.002601f
C502 VCC.n302 VSS 0.002601f
C503 VCC.n303 VSS 0.002601f
C504 VCC.n304 VSS 0.002601f
C505 VCC.n305 VSS 0.002601f
C506 VCC.n306 VSS 0.002601f
C507 VCC.n308 VSS 0.002601f
C508 VCC.n310 VSS 0.002601f
C509 VCC.n311 VSS 0.002601f
C510 VCC.n312 VSS 0.002601f
C511 VCC.n313 VSS 0.002601f
C512 VCC.n314 VSS 0.002601f
C513 VCC.n316 VSS 0.002601f
C514 VCC.n318 VSS 0.002601f
C515 VCC.n319 VSS 0.002601f
C516 VCC.n320 VSS 0.002601f
C517 VCC.n321 VSS 0.002601f
C518 VCC.n322 VSS 0.002601f
C519 VCC.n324 VSS 0.002601f
C520 VCC.n326 VSS 0.002601f
C521 VCC.n327 VSS 0.002601f
C522 VCC.n328 VSS 0.002601f
C523 VCC.n329 VSS 0.002601f
C524 VCC.n330 VSS 0.002601f
C525 VCC.n332 VSS 0.002601f
C526 VCC.n333 VSS 0.002601f
C527 VCC.n334 VSS 0.002601f
C528 VCC.n335 VSS 0.002543f
C529 VCC.n336 VSS 0.002601f
C530 VCC.n337 VSS 0.002601f
C531 VCC.n339 VSS 0.002601f
C532 VCC.n340 VSS 0.002601f
C533 VCC.n341 VSS 0.004871f
C534 VCC.n342 VSS 0.012377f
C535 VCC.n343 VSS 0.002555f
C536 VCC.n344 VSS 0.00706f
C537 VCC.n345 VSS 0.304738f
C538 VCC.n346 VSS 0.00706f
C539 VCC.n347 VSS 0.002555f
C540 VCC.n348 VSS 0.012377f
C541 VCC.n349 VSS 0.003824f
C542 VCC.n350 VSS 0.003824f
C543 VCC.n351 VSS 0.003078f
C544 VCC.n352 VSS 0.003824f
C545 VCC.n353 VSS 0.226571f
C546 VCC.n354 VSS 0.003824f
C547 VCC.n355 VSS 0.003078f
C548 VCC.n356 VSS 0.003824f
C549 VCC.n357 VSS 0.003824f
C550 VCC.n358 VSS 0.003824f
C551 VCC.n359 VSS 0.003078f
C552 VCC.n360 VSS 0.003824f
C553 VCC.n361 VSS 0.124614f
C554 VCC.n362 VSS 0.003824f
C555 VCC.n363 VSS 0.003078f
C556 VCC.n364 VSS 0.003824f
C557 VCC.n365 VSS 0.003824f
C558 VCC.n366 VSS 0.003824f
C559 VCC.n367 VSS 0.003078f
C560 VCC.n368 VSS 0.003824f
C561 VCC.n369 VSS 0.226571f
C562 VCC.n370 VSS 0.003824f
C563 VCC.n371 VSS 0.003078f
C564 VCC.n372 VSS 0.003824f
C565 VCC.n373 VSS 0.003824f
C566 VCC.n374 VSS 0.003824f
C567 VCC.n375 VSS 0.003078f
C568 VCC.n376 VSS 0.003824f
C569 VCC.n377 VSS 0.226571f
C570 VCC.n378 VSS 0.003824f
C571 VCC.n379 VSS 0.003078f
C572 VCC.n380 VSS 0.003824f
C573 VCC.n381 VSS 0.003824f
C574 VCC.n382 VSS 0.003824f
C575 VCC.n383 VSS 0.003078f
C576 VCC.n384 VSS 0.003824f
C577 VCC.n385 VSS 0.226571f
C578 VCC.n386 VSS 0.003824f
C579 VCC.n387 VSS 0.003078f
C580 VCC.n388 VSS 0.003824f
C581 VCC.n389 VSS 0.003824f
C582 VCC.n390 VSS 0.003824f
C583 VCC.n391 VSS 0.003078f
C584 VCC.n392 VSS 0.003824f
C585 VCC.n393 VSS 0.226571f
C586 VCC.n394 VSS 0.003824f
C587 VCC.n395 VSS 0.003078f
C588 VCC.n396 VSS 0.003824f
C589 VCC.n397 VSS 0.003824f
C590 VCC.n398 VSS 0.003824f
C591 VCC.n399 VSS 0.003078f
C592 VCC.n400 VSS 0.003824f
C593 VCC.t4 VSS 0.113285f
C594 VCC.n401 VSS 0.115551f
C595 VCC.n402 VSS 0.003824f
C596 VCC.n403 VSS 0.003078f
C597 VCC.n404 VSS 0.003824f
C598 VCC.n405 VSS 0.003824f
C599 VCC.n406 VSS 0.003824f
C600 VCC.n407 VSS 0.003078f
C601 VCC.n408 VSS 0.003824f
C602 VCC.n409 VSS 0.226571f
C603 VCC.n410 VSS 0.003824f
C604 VCC.n411 VSS 0.003078f
C605 VCC.n412 VSS 0.003824f
C606 VCC.n413 VSS 0.003824f
C607 VCC.n414 VSS 0.003824f
C608 VCC.n415 VSS 0.003078f
C609 VCC.n416 VSS 0.003824f
C610 VCC.n417 VSS 0.226571f
C611 VCC.n418 VSS 0.003824f
C612 VCC.n419 VSS 0.003078f
C613 VCC.n420 VSS 0.003824f
C614 VCC.n421 VSS 0.003824f
C615 VCC.n422 VSS 0.003824f
C616 VCC.n423 VSS 0.003078f
C617 VCC.n424 VSS 0.003824f
C618 VCC.n425 VSS 0.226571f
C619 VCC.n426 VSS 0.003824f
C620 VCC.n427 VSS 0.003078f
C621 VCC.n428 VSS 0.003824f
C622 VCC.n429 VSS 0.003824f
C623 VCC.n430 VSS 0.003824f
C624 VCC.n431 VSS 0.003824f
C625 VCC.n432 VSS 0.003078f
C626 VCC.n433 VSS 0.003824f
C627 VCC.n434 VSS 0.140474f
C628 VCC.n435 VSS 0.003824f
C629 VCC.n436 VSS 0.003078f
C630 VCC.n437 VSS 0.003824f
C631 VCC.n438 VSS 0.003824f
C632 VCC.n439 VSS 0.003824f
C633 VCC.n440 VSS 0.003078f
C634 VCC.n441 VSS 0.003824f
C635 VCC.n442 VSS 0.226571f
C636 VCC.n443 VSS 0.003824f
C637 VCC.n444 VSS 0.003824f
C638 VCC.n445 VSS 0.003078f
C639 VCC.n446 VSS 0.003824f
C640 VCC.n447 VSS 0.003824f
C641 VCC.n448 VSS 0.003824f
C642 VCC.n449 VSS 0.003078f
C643 VCC.n450 VSS 0.003824f
C644 VCC.n451 VSS 0.226571f
C645 VCC.n452 VSS 0.226571f
C646 VCC.n453 VSS 0.003824f
C647 VCC.n454 VSS 0.003078f
C648 VCC.n455 VSS 0.003824f
C649 VCC.n456 VSS 0.003824f
C650 VCC.n457 VSS 0.003824f
C651 VCC.n458 VSS 0.003078f
C652 VCC.n459 VSS 0.003824f
C653 VCC.n460 VSS 0.003824f
C654 VCC.n461 VSS 0.169928f
C655 VCC.n462 VSS 0.003824f
C656 VCC.n463 VSS 0.003078f
C657 VCC.n464 VSS 0.003824f
C658 VCC.n465 VSS 0.003824f
C659 VCC.n466 VSS 0.003824f
C660 VCC.n467 VSS 0.003078f
C661 VCC.n468 VSS 0.003824f
C662 VCC.n469 VSS 0.226571f
C663 VCC.n470 VSS 0.226571f
C664 VCC.n471 VSS 0.003824f
C665 VCC.n472 VSS 0.226571f
C666 VCC.n473 VSS 0.003824f
C667 VCC.n474 VSS 0.003078f
C668 VCC.n475 VSS 0.003824f
C669 VCC.n476 VSS 0.003824f
C670 VCC.n477 VSS 0.003824f
C671 VCC.n478 VSS 0.003078f
C672 VCC.n479 VSS 0.003824f
C673 VCC.n480 VSS 0.226571f
C674 VCC.n481 VSS 0.226571f
C675 VCC.t1 VSS 0.113285f
C676 VCC.n482 VSS 0.003824f
C677 VCC.n483 VSS 0.140474f
C678 VCC.n484 VSS 0.003824f
C679 VCC.n485 VSS 0.003078f
C680 VCC.n486 VSS 0.003824f
C681 VCC.n487 VSS 0.003824f
C682 VCC.n488 VSS 0.003824f
C683 VCC.n489 VSS 0.003078f
C684 VCC.n490 VSS 0.003824f
C685 VCC.n491 VSS 0.226571f
C686 VCC.n492 VSS 0.226571f
C687 VCC.n493 VSS 0.003824f
C688 VCC.n494 VSS 0.226571f
C689 VCC.n495 VSS 0.003824f
C690 VCC.n496 VSS 0.003078f
C691 VCC.n497 VSS 0.003824f
C692 VCC.n498 VSS 0.003824f
C693 VCC.n499 VSS 0.003824f
C694 VCC.n500 VSS 0.003078f
C695 VCC.n501 VSS 0.003824f
C696 VCC.n502 VSS 0.226571f
C697 VCC.n503 VSS 0.224305f
C698 VCC.t3 VSS 0.113285f
C699 VCC.n504 VSS 0.003824f
C700 VCC.n505 VSS 0.115551f
C701 VCC.n506 VSS 0.003824f
C702 VCC.n507 VSS 0.003078f
C703 VCC.n508 VSS 0.003824f
C704 VCC.n509 VSS 0.003824f
C705 VCC.n510 VSS 0.003824f
C706 VCC.n511 VSS 0.003078f
C707 VCC.n512 VSS 0.003824f
C708 VCC.n513 VSS 0.226571f
C709 VCC.n514 VSS 0.226571f
C710 VCC.n515 VSS 0.003824f
C711 VCC.n516 VSS 0.226571f
C712 VCC.n517 VSS 0.003824f
C713 VCC.n518 VSS 0.003078f
C714 VCC.n519 VSS 0.003824f
C715 VCC.n520 VSS 0.003824f
C716 VCC.n521 VSS 0.003824f
C717 VCC.n522 VSS 0.003078f
C718 VCC.n523 VSS 0.003824f
C719 VCC.n524 VSS 0.226571f
C720 VCC.n525 VSS 0.226571f
C721 VCC.n526 VSS 0.215242f
C722 VCC.n527 VSS 0.003824f
C723 VCC.n528 VSS 0.226571f
C724 VCC.n529 VSS 0.003824f
C725 VCC.n530 VSS 0.003078f
C726 VCC.n531 VSS 0.003824f
C727 VCC.n532 VSS 0.003824f
C728 VCC.n533 VSS 0.003824f
C729 VCC.n534 VSS 0.003078f
C730 VCC.n535 VSS 0.003824f
C731 VCC.n536 VSS 0.124614f
C732 VCC.n537 VSS 0.226571f
C733 VCC.n538 VSS 0.003824f
C734 VCC.n539 VSS 0.226571f
C735 VCC.n540 VSS 0.003824f
C736 VCC.n541 VSS 0.003078f
C737 VCC.n542 VSS 0.003824f
C738 VCC.n543 VSS 0.003824f
C739 VCC.n544 VSS 0.002601f
C740 VCC.n545 VSS 0.002601f
C741 VCC.n546 VSS 0.002601f
C742 VCC.n547 VSS 0.002601f
C743 VCC.n548 VSS 0.002601f
C744 VCC.n549 VSS 0.002601f
C745 VCC.n550 VSS 0.002601f
C746 VCC.n551 VSS 0.002601f
C747 VCC.n552 VSS 0.002601f
C748 VCC.n553 VSS 0.002601f
C749 VCC.n554 VSS 0.002601f
C750 VCC.n555 VSS 0.002601f
C751 VCC.n556 VSS 0.002601f
C752 VCC.n557 VSS 0.002601f
C753 VCC.n558 VSS 0.001396f
C754 VCC.n559 VSS 0.002601f
C755 VCC.n560 VSS 0.002601f
C756 VCC.n561 VSS 0.002601f
C757 VCC.n562 VSS 0.002601f
C758 VCC.n563 VSS 0.002601f
C759 VCC.n564 VSS 0.002601f
C760 VCC.n565 VSS 0.002601f
C761 VCC.n566 VSS 0.002601f
C762 VCC.n567 VSS 0.002601f
C763 VCC.n568 VSS 0.002601f
C764 VCC.n569 VSS 0.002601f
C765 VCC.n570 VSS 0.002601f
C766 VCC.n571 VSS 0.002601f
C767 VCC.n572 VSS 0.002601f
C768 VCC.n573 VSS 0.002601f
C769 VCC.n574 VSS 0.002543f
C770 VCC.n576 VSS 0.002601f
C771 VCC.n577 VSS 0.004871f
C772 VCC.n578 VSS 0.002601f
C773 VCC.t18 VSS 0.104021f
C774 VCC.t17 VSS 0.113895f
C775 VCC.t16 VSS 0.55312f
C776 VCC.n579 VSS 0.064333f
C777 VCC.n580 VSS 0.025611f
C778 VCC.n581 VSS 0.003624f
C779 VCC.n582 VSS 0.001358f
C780 VCC.n583 VSS 0.002601f
C781 VCC.n585 VSS 0.002601f
C782 VCC.n587 VSS 0.002601f
C783 VCC.n588 VSS 0.002601f
C784 VCC.n589 VSS 0.002601f
C785 VCC.n590 VSS 0.002601f
C786 VCC.n591 VSS 0.002601f
C787 VCC.n593 VSS 0.002601f
C788 VCC.n595 VSS 0.002601f
C789 VCC.n596 VSS 0.002601f
C790 VCC.n597 VSS 0.002601f
C791 VCC.n598 VSS 0.002601f
C792 VCC.n599 VSS 0.002601f
C793 VCC.n601 VSS 0.002601f
C794 VCC.n603 VSS 0.002601f
C795 VCC.n604 VSS 0.002601f
C796 VCC.n605 VSS 0.002601f
C797 VCC.n606 VSS 0.002601f
C798 VCC.n607 VSS 0.002601f
C799 VCC.n609 VSS 0.002601f
C800 VCC.n611 VSS 0.002601f
C801 VCC.n612 VSS 0.002601f
C802 VCC.n613 VSS 0.002601f
C803 VCC.n614 VSS 0.002601f
C804 VCC.n615 VSS 0.002601f
C805 VCC.n617 VSS 0.002601f
C806 VCC.n619 VSS 0.002601f
C807 VCC.n620 VSS 0.002601f
C808 VCC.n621 VSS 0.002601f
C809 VCC.n622 VSS 0.002601f
C810 VCC.n623 VSS 0.002601f
C811 VCC.n625 VSS 0.002601f
C812 VCC.n627 VSS 0.002601f
C813 VCC.n628 VSS 0.002601f
C814 VCC.n629 VSS 0.002601f
C815 VCC.n630 VSS 0.002601f
C816 VCC.n631 VSS 0.002601f
C817 VCC.n633 VSS 0.002601f
C818 VCC.n635 VSS 0.002601f
C819 VCC.n636 VSS 0.002601f
C820 VCC.n637 VSS 0.002601f
C821 VCC.n638 VSS 0.002601f
C822 VCC.n639 VSS 0.002601f
C823 VCC.n641 VSS 0.002601f
C824 VCC.n643 VSS 0.002601f
C825 VCC.n644 VSS 0.002601f
C826 VCC.n645 VSS 0.002601f
C827 VCC.t8 VSS 0.104021f
C828 VCC.t7 VSS 0.113895f
C829 VCC.t5 VSS 0.55312f
C830 VCC.n646 VSS 0.064333f
C831 VCC.n647 VSS 0.025611f
C832 VCC.n648 VSS 0.003624f
C833 VCC.n649 VSS 0.002505f
C834 VCC.n650 VSS 0.002601f
C835 VCC.n652 VSS 0.002601f
C836 VCC.n654 VSS 0.002601f
C837 VCC.n655 VSS 0.002601f
C838 VCC.n656 VSS 0.002601f
C839 VCC.n657 VSS 0.002601f
C840 VCC.n658 VSS 0.002601f
C841 VCC.n660 VSS 0.002601f
C842 VCC.n662 VSS 0.002601f
C843 VCC.n663 VSS 0.002601f
C844 VCC.n664 VSS 0.002601f
C845 VCC.n665 VSS 0.002601f
C846 VCC.n666 VSS 0.002601f
C847 VCC.n668 VSS 0.002601f
C848 VCC.n670 VSS 0.002601f
C849 VCC.n671 VSS 0.002601f
C850 VCC.n672 VSS 0.002601f
C851 VCC.n673 VSS 0.002601f
C852 VCC.n674 VSS 0.002601f
C853 VCC.n676 VSS 0.002601f
C854 VCC.n678 VSS 0.002601f
C855 VCC.n679 VSS 0.002601f
C856 VCC.n680 VSS 0.002601f
C857 VCC.n681 VSS 0.002601f
C858 VCC.n682 VSS 0.002601f
C859 VCC.n684 VSS 0.002601f
C860 VCC.n686 VSS 0.002601f
C861 VCC.n687 VSS 0.002601f
C862 VCC.n688 VSS 0.002601f
C863 VCC.n689 VSS 0.002601f
C864 VCC.n690 VSS 0.002601f
C865 VCC.n692 VSS 0.002601f
C866 VCC.n694 VSS 0.002601f
C867 VCC.n695 VSS 0.002601f
C868 VCC.n696 VSS 0.002601f
C869 VCC.n697 VSS 0.002601f
C870 VCC.n698 VSS 0.002601f
C871 VCC.n700 VSS 0.002601f
C872 VCC.n702 VSS 0.002601f
C873 VCC.n703 VSS 0.002601f
C874 VCC.n704 VSS 0.002601f
C875 VCC.n705 VSS 0.002601f
C876 VCC.n706 VSS 0.002601f
C877 VCC.n708 VSS 0.002601f
C878 VCC.n710 VSS 0.002601f
C879 VCC.n711 VSS 0.002601f
C880 VCC.n712 VSS 0.004871f
C881 VCC.n713 VSS 0.012377f
C882 VCC.n714 VSS 0.002555f
C883 VCC.n715 VSS 0.00706f
C884 VCC.n716 VSS 0.304738f
C885 VCC.n717 VSS 0.00706f
C886 VCC.n718 VSS 0.002555f
C887 VCC.n719 VSS 0.003078f
C888 VCC.n720 VSS 0.003824f
C889 VCC.n721 VSS 0.003824f
C890 VCC.n722 VSS 0.003824f
C891 VCC.n723 VSS 0.003078f
C892 VCC.n724 VSS 0.003078f
C893 VCC.n725 VSS 0.003078f
C894 VCC.n726 VSS 0.003824f
C895 VCC.n727 VSS 0.003824f
C896 VCC.n728 VSS 0.003824f
C897 VCC.n729 VSS 0.003078f
C898 VCC.n730 VSS 0.003078f
C899 VCC.n731 VSS 0.003078f
C900 VCC.n732 VSS 0.003824f
C901 VCC.n733 VSS 0.003824f
C902 VCC.n734 VSS 0.003824f
C903 VCC.n735 VSS 0.003078f
C904 VCC.n736 VSS 0.003078f
C905 VCC.n737 VSS 0.003078f
C906 VCC.n738 VSS 0.003824f
C907 VCC.n739 VSS 0.003824f
C908 VCC.n740 VSS 0.003824f
C909 VCC.n741 VSS 0.003078f
C910 VCC.n742 VSS 0.003078f
C911 VCC.n743 VSS 0.003078f
C912 VCC.n744 VSS 0.003824f
C913 VCC.n745 VSS 0.003824f
C914 VCC.n746 VSS 0.003824f
C915 VCC.n747 VSS 0.003078f
C916 VCC.n748 VSS 0.003078f
C917 VCC.n749 VSS 0.003078f
C918 VCC.n750 VSS 0.003824f
C919 VCC.n751 VSS 0.003824f
C920 VCC.n752 VSS 0.003824f
C921 VCC.n753 VSS 0.003078f
C922 VCC.n754 VSS 0.003078f
C923 VCC.n755 VSS 0.003078f
C924 VCC.n756 VSS 0.003824f
C925 VCC.n757 VSS 0.003824f
C926 VCC.n758 VSS 0.003824f
C927 VCC.n759 VSS 0.003078f
C928 VCC.n760 VSS 0.003078f
C929 VCC.n761 VSS 0.003078f
.ends

