* NGSPICE file created from diff_pair_sample_1343.ext - technology: sky130A

.subckt diff_pair_sample_1343 VTAIL VN VP B VDD2 VDD1
X0 B.t15 B.t13 B.t14 B.t3 sky130_fd_pr__nfet_01v8 ad=1.1193 pd=6.52 as=0 ps=0 w=2.87 l=2.07
X1 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=1.1193 pd=6.52 as=0 ps=0 w=2.87 l=2.07
X2 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=1.1193 pd=6.52 as=0 ps=0 w=2.87 l=2.07
X3 VDD2.t1 VN.t0 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=1.1193 pd=6.52 as=1.1193 ps=6.52 w=2.87 l=2.07
X4 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=1.1193 pd=6.52 as=0 ps=0 w=2.87 l=2.07
X5 VDD2.t0 VN.t1 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=1.1193 pd=6.52 as=1.1193 ps=6.52 w=2.87 l=2.07
X6 VDD1.t1 VP.t0 VTAIL.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=1.1193 pd=6.52 as=1.1193 ps=6.52 w=2.87 l=2.07
X7 VDD1.t0 VP.t1 VTAIL.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=1.1193 pd=6.52 as=1.1193 ps=6.52 w=2.87 l=2.07
R0 B.n308 B.n307 585
R1 B.n308 B.n43 585
R2 B.n311 B.n310 585
R3 B.n312 B.n67 585
R4 B.n314 B.n313 585
R5 B.n316 B.n66 585
R6 B.n319 B.n318 585
R7 B.n320 B.n65 585
R8 B.n322 B.n321 585
R9 B.n324 B.n64 585
R10 B.n327 B.n326 585
R11 B.n328 B.n63 585
R12 B.n330 B.n329 585
R13 B.n332 B.n62 585
R14 B.n335 B.n334 585
R15 B.n336 B.n59 585
R16 B.n339 B.n338 585
R17 B.n341 B.n58 585
R18 B.n344 B.n343 585
R19 B.n345 B.n57 585
R20 B.n347 B.n346 585
R21 B.n349 B.n56 585
R22 B.n352 B.n351 585
R23 B.n353 B.n52 585
R24 B.n355 B.n354 585
R25 B.n357 B.n51 585
R26 B.n360 B.n359 585
R27 B.n361 B.n50 585
R28 B.n363 B.n362 585
R29 B.n365 B.n49 585
R30 B.n368 B.n367 585
R31 B.n369 B.n48 585
R32 B.n371 B.n370 585
R33 B.n373 B.n47 585
R34 B.n376 B.n375 585
R35 B.n377 B.n46 585
R36 B.n379 B.n378 585
R37 B.n381 B.n45 585
R38 B.n384 B.n383 585
R39 B.n385 B.n44 585
R40 B.n306 B.n42 585
R41 B.n388 B.n42 585
R42 B.n305 B.n41 585
R43 B.n389 B.n41 585
R44 B.n304 B.n40 585
R45 B.n390 B.n40 585
R46 B.n303 B.n302 585
R47 B.n302 B.n36 585
R48 B.n301 B.n35 585
R49 B.n396 B.n35 585
R50 B.n300 B.n34 585
R51 B.n397 B.n34 585
R52 B.n299 B.n33 585
R53 B.n398 B.n33 585
R54 B.n298 B.n297 585
R55 B.n297 B.n29 585
R56 B.n296 B.n28 585
R57 B.n404 B.n28 585
R58 B.n295 B.n27 585
R59 B.n405 B.n27 585
R60 B.n294 B.n26 585
R61 B.n406 B.n26 585
R62 B.n293 B.n292 585
R63 B.n292 B.n22 585
R64 B.n291 B.n21 585
R65 B.n412 B.n21 585
R66 B.n290 B.n20 585
R67 B.n413 B.n20 585
R68 B.n289 B.n19 585
R69 B.n414 B.n19 585
R70 B.n288 B.n287 585
R71 B.n287 B.n15 585
R72 B.n286 B.n14 585
R73 B.n420 B.n14 585
R74 B.n285 B.n13 585
R75 B.n421 B.n13 585
R76 B.n284 B.n12 585
R77 B.n422 B.n12 585
R78 B.n283 B.n282 585
R79 B.n282 B.n8 585
R80 B.n281 B.n7 585
R81 B.n428 B.n7 585
R82 B.n280 B.n6 585
R83 B.n429 B.n6 585
R84 B.n279 B.n5 585
R85 B.n430 B.n5 585
R86 B.n278 B.n277 585
R87 B.n277 B.n4 585
R88 B.n276 B.n68 585
R89 B.n276 B.n275 585
R90 B.n266 B.n69 585
R91 B.n70 B.n69 585
R92 B.n268 B.n267 585
R93 B.n269 B.n268 585
R94 B.n265 B.n75 585
R95 B.n75 B.n74 585
R96 B.n264 B.n263 585
R97 B.n263 B.n262 585
R98 B.n77 B.n76 585
R99 B.n78 B.n77 585
R100 B.n255 B.n254 585
R101 B.n256 B.n255 585
R102 B.n253 B.n83 585
R103 B.n83 B.n82 585
R104 B.n252 B.n251 585
R105 B.n251 B.n250 585
R106 B.n85 B.n84 585
R107 B.n86 B.n85 585
R108 B.n243 B.n242 585
R109 B.n244 B.n243 585
R110 B.n241 B.n91 585
R111 B.n91 B.n90 585
R112 B.n240 B.n239 585
R113 B.n239 B.n238 585
R114 B.n93 B.n92 585
R115 B.n94 B.n93 585
R116 B.n231 B.n230 585
R117 B.n232 B.n231 585
R118 B.n229 B.n99 585
R119 B.n99 B.n98 585
R120 B.n228 B.n227 585
R121 B.n227 B.n226 585
R122 B.n101 B.n100 585
R123 B.n102 B.n101 585
R124 B.n219 B.n218 585
R125 B.n220 B.n219 585
R126 B.n217 B.n107 585
R127 B.n107 B.n106 585
R128 B.n216 B.n215 585
R129 B.n215 B.n214 585
R130 B.n211 B.n111 585
R131 B.n210 B.n209 585
R132 B.n207 B.n112 585
R133 B.n207 B.n110 585
R134 B.n206 B.n205 585
R135 B.n204 B.n203 585
R136 B.n202 B.n114 585
R137 B.n200 B.n199 585
R138 B.n198 B.n115 585
R139 B.n197 B.n196 585
R140 B.n194 B.n116 585
R141 B.n192 B.n191 585
R142 B.n190 B.n117 585
R143 B.n189 B.n188 585
R144 B.n186 B.n118 585
R145 B.n184 B.n183 585
R146 B.n181 B.n119 585
R147 B.n180 B.n179 585
R148 B.n177 B.n122 585
R149 B.n175 B.n174 585
R150 B.n173 B.n123 585
R151 B.n172 B.n171 585
R152 B.n169 B.n124 585
R153 B.n167 B.n166 585
R154 B.n165 B.n125 585
R155 B.n163 B.n162 585
R156 B.n160 B.n128 585
R157 B.n158 B.n157 585
R158 B.n156 B.n129 585
R159 B.n155 B.n154 585
R160 B.n152 B.n130 585
R161 B.n150 B.n149 585
R162 B.n148 B.n131 585
R163 B.n147 B.n146 585
R164 B.n144 B.n132 585
R165 B.n142 B.n141 585
R166 B.n140 B.n133 585
R167 B.n139 B.n138 585
R168 B.n136 B.n134 585
R169 B.n109 B.n108 585
R170 B.n213 B.n212 585
R171 B.n214 B.n213 585
R172 B.n105 B.n104 585
R173 B.n106 B.n105 585
R174 B.n222 B.n221 585
R175 B.n221 B.n220 585
R176 B.n223 B.n103 585
R177 B.n103 B.n102 585
R178 B.n225 B.n224 585
R179 B.n226 B.n225 585
R180 B.n97 B.n96 585
R181 B.n98 B.n97 585
R182 B.n234 B.n233 585
R183 B.n233 B.n232 585
R184 B.n235 B.n95 585
R185 B.n95 B.n94 585
R186 B.n237 B.n236 585
R187 B.n238 B.n237 585
R188 B.n89 B.n88 585
R189 B.n90 B.n89 585
R190 B.n246 B.n245 585
R191 B.n245 B.n244 585
R192 B.n247 B.n87 585
R193 B.n87 B.n86 585
R194 B.n249 B.n248 585
R195 B.n250 B.n249 585
R196 B.n81 B.n80 585
R197 B.n82 B.n81 585
R198 B.n258 B.n257 585
R199 B.n257 B.n256 585
R200 B.n259 B.n79 585
R201 B.n79 B.n78 585
R202 B.n261 B.n260 585
R203 B.n262 B.n261 585
R204 B.n73 B.n72 585
R205 B.n74 B.n73 585
R206 B.n271 B.n270 585
R207 B.n270 B.n269 585
R208 B.n272 B.n71 585
R209 B.n71 B.n70 585
R210 B.n274 B.n273 585
R211 B.n275 B.n274 585
R212 B.n2 B.n0 585
R213 B.n4 B.n2 585
R214 B.n3 B.n1 585
R215 B.n429 B.n3 585
R216 B.n427 B.n426 585
R217 B.n428 B.n427 585
R218 B.n425 B.n9 585
R219 B.n9 B.n8 585
R220 B.n424 B.n423 585
R221 B.n423 B.n422 585
R222 B.n11 B.n10 585
R223 B.n421 B.n11 585
R224 B.n419 B.n418 585
R225 B.n420 B.n419 585
R226 B.n417 B.n16 585
R227 B.n16 B.n15 585
R228 B.n416 B.n415 585
R229 B.n415 B.n414 585
R230 B.n18 B.n17 585
R231 B.n413 B.n18 585
R232 B.n411 B.n410 585
R233 B.n412 B.n411 585
R234 B.n409 B.n23 585
R235 B.n23 B.n22 585
R236 B.n408 B.n407 585
R237 B.n407 B.n406 585
R238 B.n25 B.n24 585
R239 B.n405 B.n25 585
R240 B.n403 B.n402 585
R241 B.n404 B.n403 585
R242 B.n401 B.n30 585
R243 B.n30 B.n29 585
R244 B.n400 B.n399 585
R245 B.n399 B.n398 585
R246 B.n32 B.n31 585
R247 B.n397 B.n32 585
R248 B.n395 B.n394 585
R249 B.n396 B.n395 585
R250 B.n393 B.n37 585
R251 B.n37 B.n36 585
R252 B.n392 B.n391 585
R253 B.n391 B.n390 585
R254 B.n39 B.n38 585
R255 B.n389 B.n39 585
R256 B.n387 B.n386 585
R257 B.n388 B.n387 585
R258 B.n432 B.n431 585
R259 B.n431 B.n430 585
R260 B.n213 B.n111 545.355
R261 B.n387 B.n44 545.355
R262 B.n215 B.n109 545.355
R263 B.n308 B.n42 545.355
R264 B.n309 B.n43 256.663
R265 B.n315 B.n43 256.663
R266 B.n317 B.n43 256.663
R267 B.n323 B.n43 256.663
R268 B.n325 B.n43 256.663
R269 B.n331 B.n43 256.663
R270 B.n333 B.n43 256.663
R271 B.n340 B.n43 256.663
R272 B.n342 B.n43 256.663
R273 B.n348 B.n43 256.663
R274 B.n350 B.n43 256.663
R275 B.n356 B.n43 256.663
R276 B.n358 B.n43 256.663
R277 B.n364 B.n43 256.663
R278 B.n366 B.n43 256.663
R279 B.n372 B.n43 256.663
R280 B.n374 B.n43 256.663
R281 B.n380 B.n43 256.663
R282 B.n382 B.n43 256.663
R283 B.n208 B.n110 256.663
R284 B.n113 B.n110 256.663
R285 B.n201 B.n110 256.663
R286 B.n195 B.n110 256.663
R287 B.n193 B.n110 256.663
R288 B.n187 B.n110 256.663
R289 B.n185 B.n110 256.663
R290 B.n178 B.n110 256.663
R291 B.n176 B.n110 256.663
R292 B.n170 B.n110 256.663
R293 B.n168 B.n110 256.663
R294 B.n161 B.n110 256.663
R295 B.n159 B.n110 256.663
R296 B.n153 B.n110 256.663
R297 B.n151 B.n110 256.663
R298 B.n145 B.n110 256.663
R299 B.n143 B.n110 256.663
R300 B.n137 B.n110 256.663
R301 B.n135 B.n110 256.663
R302 B.n126 B.t2 240.492
R303 B.n120 B.t13 240.492
R304 B.n53 B.t10 240.492
R305 B.n60 B.t6 240.492
R306 B.n214 B.n110 187.724
R307 B.n388 B.n43 187.724
R308 B.n213 B.n105 163.367
R309 B.n221 B.n105 163.367
R310 B.n221 B.n103 163.367
R311 B.n225 B.n103 163.367
R312 B.n225 B.n97 163.367
R313 B.n233 B.n97 163.367
R314 B.n233 B.n95 163.367
R315 B.n237 B.n95 163.367
R316 B.n237 B.n89 163.367
R317 B.n245 B.n89 163.367
R318 B.n245 B.n87 163.367
R319 B.n249 B.n87 163.367
R320 B.n249 B.n81 163.367
R321 B.n257 B.n81 163.367
R322 B.n257 B.n79 163.367
R323 B.n261 B.n79 163.367
R324 B.n261 B.n73 163.367
R325 B.n270 B.n73 163.367
R326 B.n270 B.n71 163.367
R327 B.n274 B.n71 163.367
R328 B.n274 B.n2 163.367
R329 B.n431 B.n2 163.367
R330 B.n431 B.n3 163.367
R331 B.n427 B.n3 163.367
R332 B.n427 B.n9 163.367
R333 B.n423 B.n9 163.367
R334 B.n423 B.n11 163.367
R335 B.n419 B.n11 163.367
R336 B.n419 B.n16 163.367
R337 B.n415 B.n16 163.367
R338 B.n415 B.n18 163.367
R339 B.n411 B.n18 163.367
R340 B.n411 B.n23 163.367
R341 B.n407 B.n23 163.367
R342 B.n407 B.n25 163.367
R343 B.n403 B.n25 163.367
R344 B.n403 B.n30 163.367
R345 B.n399 B.n30 163.367
R346 B.n399 B.n32 163.367
R347 B.n395 B.n32 163.367
R348 B.n395 B.n37 163.367
R349 B.n391 B.n37 163.367
R350 B.n391 B.n39 163.367
R351 B.n387 B.n39 163.367
R352 B.n209 B.n207 163.367
R353 B.n207 B.n206 163.367
R354 B.n203 B.n202 163.367
R355 B.n200 B.n115 163.367
R356 B.n196 B.n194 163.367
R357 B.n192 B.n117 163.367
R358 B.n188 B.n186 163.367
R359 B.n184 B.n119 163.367
R360 B.n179 B.n177 163.367
R361 B.n175 B.n123 163.367
R362 B.n171 B.n169 163.367
R363 B.n167 B.n125 163.367
R364 B.n162 B.n160 163.367
R365 B.n158 B.n129 163.367
R366 B.n154 B.n152 163.367
R367 B.n150 B.n131 163.367
R368 B.n146 B.n144 163.367
R369 B.n142 B.n133 163.367
R370 B.n138 B.n136 163.367
R371 B.n215 B.n107 163.367
R372 B.n219 B.n107 163.367
R373 B.n219 B.n101 163.367
R374 B.n227 B.n101 163.367
R375 B.n227 B.n99 163.367
R376 B.n231 B.n99 163.367
R377 B.n231 B.n93 163.367
R378 B.n239 B.n93 163.367
R379 B.n239 B.n91 163.367
R380 B.n243 B.n91 163.367
R381 B.n243 B.n85 163.367
R382 B.n251 B.n85 163.367
R383 B.n251 B.n83 163.367
R384 B.n255 B.n83 163.367
R385 B.n255 B.n77 163.367
R386 B.n263 B.n77 163.367
R387 B.n263 B.n75 163.367
R388 B.n268 B.n75 163.367
R389 B.n268 B.n69 163.367
R390 B.n276 B.n69 163.367
R391 B.n277 B.n276 163.367
R392 B.n277 B.n5 163.367
R393 B.n6 B.n5 163.367
R394 B.n7 B.n6 163.367
R395 B.n282 B.n7 163.367
R396 B.n282 B.n12 163.367
R397 B.n13 B.n12 163.367
R398 B.n14 B.n13 163.367
R399 B.n287 B.n14 163.367
R400 B.n287 B.n19 163.367
R401 B.n20 B.n19 163.367
R402 B.n21 B.n20 163.367
R403 B.n292 B.n21 163.367
R404 B.n292 B.n26 163.367
R405 B.n27 B.n26 163.367
R406 B.n28 B.n27 163.367
R407 B.n297 B.n28 163.367
R408 B.n297 B.n33 163.367
R409 B.n34 B.n33 163.367
R410 B.n35 B.n34 163.367
R411 B.n302 B.n35 163.367
R412 B.n302 B.n40 163.367
R413 B.n41 B.n40 163.367
R414 B.n42 B.n41 163.367
R415 B.n383 B.n381 163.367
R416 B.n379 B.n46 163.367
R417 B.n375 B.n373 163.367
R418 B.n371 B.n48 163.367
R419 B.n367 B.n365 163.367
R420 B.n363 B.n50 163.367
R421 B.n359 B.n357 163.367
R422 B.n355 B.n52 163.367
R423 B.n351 B.n349 163.367
R424 B.n347 B.n57 163.367
R425 B.n343 B.n341 163.367
R426 B.n339 B.n59 163.367
R427 B.n334 B.n332 163.367
R428 B.n330 B.n63 163.367
R429 B.n326 B.n324 163.367
R430 B.n322 B.n65 163.367
R431 B.n318 B.n316 163.367
R432 B.n314 B.n67 163.367
R433 B.n310 B.n308 163.367
R434 B.n126 B.t5 124.939
R435 B.n60 B.t8 124.939
R436 B.n120 B.t15 124.936
R437 B.n53 B.t11 124.936
R438 B.n214 B.n106 91.836
R439 B.n220 B.n106 91.836
R440 B.n220 B.n102 91.836
R441 B.n226 B.n102 91.836
R442 B.n226 B.n98 91.836
R443 B.n232 B.n98 91.836
R444 B.n238 B.n94 91.836
R445 B.n238 B.n90 91.836
R446 B.n244 B.n90 91.836
R447 B.n244 B.n86 91.836
R448 B.n250 B.n86 91.836
R449 B.n250 B.n82 91.836
R450 B.n256 B.n82 91.836
R451 B.n256 B.n78 91.836
R452 B.n262 B.n78 91.836
R453 B.n269 B.n74 91.836
R454 B.n269 B.n70 91.836
R455 B.n275 B.n70 91.836
R456 B.n275 B.n4 91.836
R457 B.n430 B.n4 91.836
R458 B.n430 B.n429 91.836
R459 B.n429 B.n428 91.836
R460 B.n428 B.n8 91.836
R461 B.n422 B.n8 91.836
R462 B.n422 B.n421 91.836
R463 B.n420 B.n15 91.836
R464 B.n414 B.n15 91.836
R465 B.n414 B.n413 91.836
R466 B.n413 B.n412 91.836
R467 B.n412 B.n22 91.836
R468 B.n406 B.n22 91.836
R469 B.n406 B.n405 91.836
R470 B.n405 B.n404 91.836
R471 B.n404 B.n29 91.836
R472 B.n398 B.n397 91.836
R473 B.n397 B.n396 91.836
R474 B.n396 B.n36 91.836
R475 B.n390 B.n36 91.836
R476 B.n390 B.n389 91.836
R477 B.n389 B.n388 91.836
R478 B.n262 B.t1 79.6813
R479 B.t0 B.n420 79.6813
R480 B.n127 B.t4 78.3925
R481 B.n61 B.t9 78.3925
R482 B.n121 B.t14 78.3907
R483 B.n54 B.t12 78.3907
R484 B.n208 B.n111 71.676
R485 B.n206 B.n113 71.676
R486 B.n202 B.n201 71.676
R487 B.n195 B.n115 71.676
R488 B.n194 B.n193 71.676
R489 B.n187 B.n117 71.676
R490 B.n186 B.n185 71.676
R491 B.n178 B.n119 71.676
R492 B.n177 B.n176 71.676
R493 B.n170 B.n123 71.676
R494 B.n169 B.n168 71.676
R495 B.n161 B.n125 71.676
R496 B.n160 B.n159 71.676
R497 B.n153 B.n129 71.676
R498 B.n152 B.n151 71.676
R499 B.n145 B.n131 71.676
R500 B.n144 B.n143 71.676
R501 B.n137 B.n133 71.676
R502 B.n136 B.n135 71.676
R503 B.n382 B.n44 71.676
R504 B.n381 B.n380 71.676
R505 B.n374 B.n46 71.676
R506 B.n373 B.n372 71.676
R507 B.n366 B.n48 71.676
R508 B.n365 B.n364 71.676
R509 B.n358 B.n50 71.676
R510 B.n357 B.n356 71.676
R511 B.n350 B.n52 71.676
R512 B.n349 B.n348 71.676
R513 B.n342 B.n57 71.676
R514 B.n341 B.n340 71.676
R515 B.n333 B.n59 71.676
R516 B.n332 B.n331 71.676
R517 B.n325 B.n63 71.676
R518 B.n324 B.n323 71.676
R519 B.n317 B.n65 71.676
R520 B.n316 B.n315 71.676
R521 B.n309 B.n67 71.676
R522 B.n310 B.n309 71.676
R523 B.n315 B.n314 71.676
R524 B.n318 B.n317 71.676
R525 B.n323 B.n322 71.676
R526 B.n326 B.n325 71.676
R527 B.n331 B.n330 71.676
R528 B.n334 B.n333 71.676
R529 B.n340 B.n339 71.676
R530 B.n343 B.n342 71.676
R531 B.n348 B.n347 71.676
R532 B.n351 B.n350 71.676
R533 B.n356 B.n355 71.676
R534 B.n359 B.n358 71.676
R535 B.n364 B.n363 71.676
R536 B.n367 B.n366 71.676
R537 B.n372 B.n371 71.676
R538 B.n375 B.n374 71.676
R539 B.n380 B.n379 71.676
R540 B.n383 B.n382 71.676
R541 B.n209 B.n208 71.676
R542 B.n203 B.n113 71.676
R543 B.n201 B.n200 71.676
R544 B.n196 B.n195 71.676
R545 B.n193 B.n192 71.676
R546 B.n188 B.n187 71.676
R547 B.n185 B.n184 71.676
R548 B.n179 B.n178 71.676
R549 B.n176 B.n175 71.676
R550 B.n171 B.n170 71.676
R551 B.n168 B.n167 71.676
R552 B.n162 B.n161 71.676
R553 B.n159 B.n158 71.676
R554 B.n154 B.n153 71.676
R555 B.n151 B.n150 71.676
R556 B.n146 B.n145 71.676
R557 B.n143 B.n142 71.676
R558 B.n138 B.n137 71.676
R559 B.n135 B.n109 71.676
R560 B.n164 B.n127 59.5399
R561 B.n182 B.n121 59.5399
R562 B.n55 B.n54 59.5399
R563 B.n337 B.n61 59.5399
R564 B.n232 B.t3 55.3719
R565 B.n398 B.t7 55.3719
R566 B.n127 B.n126 46.546
R567 B.n121 B.n120 46.546
R568 B.n54 B.n53 46.546
R569 B.n61 B.n60 46.546
R570 B.t3 B.n94 36.4646
R571 B.t7 B.n29 36.4646
R572 B.n307 B.n306 35.4346
R573 B.n386 B.n385 35.4346
R574 B.n216 B.n108 35.4346
R575 B.n212 B.n211 35.4346
R576 B B.n432 18.0485
R577 B.t1 B.n74 12.1552
R578 B.n421 B.t0 12.1552
R579 B.n385 B.n384 10.6151
R580 B.n384 B.n45 10.6151
R581 B.n378 B.n45 10.6151
R582 B.n378 B.n377 10.6151
R583 B.n377 B.n376 10.6151
R584 B.n376 B.n47 10.6151
R585 B.n370 B.n47 10.6151
R586 B.n370 B.n369 10.6151
R587 B.n369 B.n368 10.6151
R588 B.n368 B.n49 10.6151
R589 B.n362 B.n49 10.6151
R590 B.n362 B.n361 10.6151
R591 B.n361 B.n360 10.6151
R592 B.n360 B.n51 10.6151
R593 B.n354 B.n353 10.6151
R594 B.n353 B.n352 10.6151
R595 B.n352 B.n56 10.6151
R596 B.n346 B.n56 10.6151
R597 B.n346 B.n345 10.6151
R598 B.n345 B.n344 10.6151
R599 B.n344 B.n58 10.6151
R600 B.n338 B.n58 10.6151
R601 B.n336 B.n335 10.6151
R602 B.n335 B.n62 10.6151
R603 B.n329 B.n62 10.6151
R604 B.n329 B.n328 10.6151
R605 B.n328 B.n327 10.6151
R606 B.n327 B.n64 10.6151
R607 B.n321 B.n64 10.6151
R608 B.n321 B.n320 10.6151
R609 B.n320 B.n319 10.6151
R610 B.n319 B.n66 10.6151
R611 B.n313 B.n66 10.6151
R612 B.n313 B.n312 10.6151
R613 B.n312 B.n311 10.6151
R614 B.n311 B.n307 10.6151
R615 B.n217 B.n216 10.6151
R616 B.n218 B.n217 10.6151
R617 B.n218 B.n100 10.6151
R618 B.n228 B.n100 10.6151
R619 B.n229 B.n228 10.6151
R620 B.n230 B.n229 10.6151
R621 B.n230 B.n92 10.6151
R622 B.n240 B.n92 10.6151
R623 B.n241 B.n240 10.6151
R624 B.n242 B.n241 10.6151
R625 B.n242 B.n84 10.6151
R626 B.n252 B.n84 10.6151
R627 B.n253 B.n252 10.6151
R628 B.n254 B.n253 10.6151
R629 B.n254 B.n76 10.6151
R630 B.n264 B.n76 10.6151
R631 B.n265 B.n264 10.6151
R632 B.n267 B.n265 10.6151
R633 B.n267 B.n266 10.6151
R634 B.n266 B.n68 10.6151
R635 B.n278 B.n68 10.6151
R636 B.n279 B.n278 10.6151
R637 B.n280 B.n279 10.6151
R638 B.n281 B.n280 10.6151
R639 B.n283 B.n281 10.6151
R640 B.n284 B.n283 10.6151
R641 B.n285 B.n284 10.6151
R642 B.n286 B.n285 10.6151
R643 B.n288 B.n286 10.6151
R644 B.n289 B.n288 10.6151
R645 B.n290 B.n289 10.6151
R646 B.n291 B.n290 10.6151
R647 B.n293 B.n291 10.6151
R648 B.n294 B.n293 10.6151
R649 B.n295 B.n294 10.6151
R650 B.n296 B.n295 10.6151
R651 B.n298 B.n296 10.6151
R652 B.n299 B.n298 10.6151
R653 B.n300 B.n299 10.6151
R654 B.n301 B.n300 10.6151
R655 B.n303 B.n301 10.6151
R656 B.n304 B.n303 10.6151
R657 B.n305 B.n304 10.6151
R658 B.n306 B.n305 10.6151
R659 B.n211 B.n210 10.6151
R660 B.n210 B.n112 10.6151
R661 B.n205 B.n112 10.6151
R662 B.n205 B.n204 10.6151
R663 B.n204 B.n114 10.6151
R664 B.n199 B.n114 10.6151
R665 B.n199 B.n198 10.6151
R666 B.n198 B.n197 10.6151
R667 B.n197 B.n116 10.6151
R668 B.n191 B.n116 10.6151
R669 B.n191 B.n190 10.6151
R670 B.n190 B.n189 10.6151
R671 B.n189 B.n118 10.6151
R672 B.n183 B.n118 10.6151
R673 B.n181 B.n180 10.6151
R674 B.n180 B.n122 10.6151
R675 B.n174 B.n122 10.6151
R676 B.n174 B.n173 10.6151
R677 B.n173 B.n172 10.6151
R678 B.n172 B.n124 10.6151
R679 B.n166 B.n124 10.6151
R680 B.n166 B.n165 10.6151
R681 B.n163 B.n128 10.6151
R682 B.n157 B.n128 10.6151
R683 B.n157 B.n156 10.6151
R684 B.n156 B.n155 10.6151
R685 B.n155 B.n130 10.6151
R686 B.n149 B.n130 10.6151
R687 B.n149 B.n148 10.6151
R688 B.n148 B.n147 10.6151
R689 B.n147 B.n132 10.6151
R690 B.n141 B.n132 10.6151
R691 B.n141 B.n140 10.6151
R692 B.n140 B.n139 10.6151
R693 B.n139 B.n134 10.6151
R694 B.n134 B.n108 10.6151
R695 B.n212 B.n104 10.6151
R696 B.n222 B.n104 10.6151
R697 B.n223 B.n222 10.6151
R698 B.n224 B.n223 10.6151
R699 B.n224 B.n96 10.6151
R700 B.n234 B.n96 10.6151
R701 B.n235 B.n234 10.6151
R702 B.n236 B.n235 10.6151
R703 B.n236 B.n88 10.6151
R704 B.n246 B.n88 10.6151
R705 B.n247 B.n246 10.6151
R706 B.n248 B.n247 10.6151
R707 B.n248 B.n80 10.6151
R708 B.n258 B.n80 10.6151
R709 B.n259 B.n258 10.6151
R710 B.n260 B.n259 10.6151
R711 B.n260 B.n72 10.6151
R712 B.n271 B.n72 10.6151
R713 B.n272 B.n271 10.6151
R714 B.n273 B.n272 10.6151
R715 B.n273 B.n0 10.6151
R716 B.n426 B.n1 10.6151
R717 B.n426 B.n425 10.6151
R718 B.n425 B.n424 10.6151
R719 B.n424 B.n10 10.6151
R720 B.n418 B.n10 10.6151
R721 B.n418 B.n417 10.6151
R722 B.n417 B.n416 10.6151
R723 B.n416 B.n17 10.6151
R724 B.n410 B.n17 10.6151
R725 B.n410 B.n409 10.6151
R726 B.n409 B.n408 10.6151
R727 B.n408 B.n24 10.6151
R728 B.n402 B.n24 10.6151
R729 B.n402 B.n401 10.6151
R730 B.n401 B.n400 10.6151
R731 B.n400 B.n31 10.6151
R732 B.n394 B.n31 10.6151
R733 B.n394 B.n393 10.6151
R734 B.n393 B.n392 10.6151
R735 B.n392 B.n38 10.6151
R736 B.n386 B.n38 10.6151
R737 B.n354 B.n55 6.5566
R738 B.n338 B.n337 6.5566
R739 B.n182 B.n181 6.5566
R740 B.n165 B.n164 6.5566
R741 B.n55 B.n51 4.05904
R742 B.n337 B.n336 4.05904
R743 B.n183 B.n182 4.05904
R744 B.n164 B.n163 4.05904
R745 B.n432 B.n0 2.81026
R746 B.n432 B.n1 2.81026
R747 VN VN.t0 128.8
R748 VN VN.t1 92.5164
R749 VTAIL.n1 VTAIL.t3 73.1821
R750 VTAIL.n3 VTAIL.t2 73.1818
R751 VTAIL.n0 VTAIL.t0 73.1818
R752 VTAIL.n2 VTAIL.t1 73.1818
R753 VTAIL.n1 VTAIL.n0 18.9789
R754 VTAIL.n3 VTAIL.n2 16.91
R755 VTAIL.n2 VTAIL.n1 1.50481
R756 VTAIL VTAIL.n0 1.04576
R757 VTAIL VTAIL.n3 0.459552
R758 VDD2.n0 VDD2.t0 120.132
R759 VDD2.n0 VDD2.t1 89.8606
R760 VDD2 VDD2.n0 0.575931
R761 VP.n0 VP.t0 128.609
R762 VP.n0 VP.t1 92.2753
R763 VP VP.n0 0.241678
R764 VDD1 VDD1.t0 121.174
R765 VDD1 VDD1.t1 90.4361
C0 VP VTAIL 0.993522f
C1 VDD1 VDD2 0.610238f
C2 VN VP 3.51934f
C3 VN VTAIL 0.97936f
C4 VP VDD2 0.31573f
C5 VDD2 VTAIL 2.54811f
C6 VN VDD2 0.831138f
C7 VDD1 VP 0.992257f
C8 VDD1 VTAIL 2.49911f
C9 VDD1 VN 0.153108f
C10 VDD2 B 2.566968f
C11 VDD1 B 4.31057f
C12 VTAIL B 3.205231f
C13 VN B 6.94745f
C14 VP B 4.941696f
C15 VDD1.t1 B 0.334155f
C16 VDD1.t0 B 0.526916f
C17 VP.t0 B 0.948334f
C18 VP.t1 B 0.638142f
C19 VP.n0 B 1.86454f
C20 VDD2.t0 B 0.522567f
C21 VDD2.t1 B 0.340919f
C22 VDD2.n0 B 1.55285f
C23 VTAIL.t0 B 0.36779f
C24 VTAIL.n0 B 0.917674f
C25 VTAIL.t3 B 0.367791f
C26 VTAIL.n1 B 0.945965f
C27 VTAIL.t1 B 0.36779f
C28 VTAIL.n2 B 0.818455f
C29 VTAIL.t2 B 0.36779f
C30 VTAIL.n3 B 0.754036f
C31 VN.t1 B 0.631534f
C32 VN.t0 B 0.942732f
.ends

