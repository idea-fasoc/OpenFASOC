* NGSPICE file created from diff_pair_sample_0333.ext - technology: sky130A

.subckt diff_pair_sample_0333 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t11 w_n4474_n1944# sky130_fd_pr__pfet_01v8 ad=0.8052 pd=5.21 as=1.9032 ps=10.54 w=4.88 l=2.59
X1 VDD1.t8 VP.t1 VTAIL.t9 w_n4474_n1944# sky130_fd_pr__pfet_01v8 ad=0.8052 pd=5.21 as=1.9032 ps=10.54 w=4.88 l=2.59
X2 VDD1.t7 VP.t2 VTAIL.t16 w_n4474_n1944# sky130_fd_pr__pfet_01v8 ad=0.8052 pd=5.21 as=0.8052 ps=5.21 w=4.88 l=2.59
X3 VDD1.t6 VP.t3 VTAIL.t7 w_n4474_n1944# sky130_fd_pr__pfet_01v8 ad=1.9032 pd=10.54 as=0.8052 ps=5.21 w=4.88 l=2.59
X4 VTAIL.t14 VP.t4 VDD1.t5 w_n4474_n1944# sky130_fd_pr__pfet_01v8 ad=0.8052 pd=5.21 as=0.8052 ps=5.21 w=4.88 l=2.59
X5 VDD2.t9 VN.t0 VTAIL.t5 w_n4474_n1944# sky130_fd_pr__pfet_01v8 ad=0.8052 pd=5.21 as=0.8052 ps=5.21 w=4.88 l=2.59
X6 B.t11 B.t9 B.t10 w_n4474_n1944# sky130_fd_pr__pfet_01v8 ad=1.9032 pd=10.54 as=0 ps=0 w=4.88 l=2.59
X7 VDD2.t8 VN.t1 VTAIL.t1 w_n4474_n1944# sky130_fd_pr__pfet_01v8 ad=0.8052 pd=5.21 as=1.9032 ps=10.54 w=4.88 l=2.59
X8 VDD2.t7 VN.t2 VTAIL.t18 w_n4474_n1944# sky130_fd_pr__pfet_01v8 ad=1.9032 pd=10.54 as=0.8052 ps=5.21 w=4.88 l=2.59
X9 VDD2.t6 VN.t3 VTAIL.t4 w_n4474_n1944# sky130_fd_pr__pfet_01v8 ad=0.8052 pd=5.21 as=1.9032 ps=10.54 w=4.88 l=2.59
X10 VTAIL.t17 VN.t4 VDD2.t5 w_n4474_n1944# sky130_fd_pr__pfet_01v8 ad=0.8052 pd=5.21 as=0.8052 ps=5.21 w=4.88 l=2.59
X11 B.t8 B.t6 B.t7 w_n4474_n1944# sky130_fd_pr__pfet_01v8 ad=1.9032 pd=10.54 as=0 ps=0 w=4.88 l=2.59
X12 VDD2.t4 VN.t5 VTAIL.t6 w_n4474_n1944# sky130_fd_pr__pfet_01v8 ad=0.8052 pd=5.21 as=0.8052 ps=5.21 w=4.88 l=2.59
X13 VTAIL.t12 VP.t5 VDD1.t4 w_n4474_n1944# sky130_fd_pr__pfet_01v8 ad=0.8052 pd=5.21 as=0.8052 ps=5.21 w=4.88 l=2.59
X14 VDD2.t3 VN.t6 VTAIL.t0 w_n4474_n1944# sky130_fd_pr__pfet_01v8 ad=1.9032 pd=10.54 as=0.8052 ps=5.21 w=4.88 l=2.59
X15 VDD1.t3 VP.t6 VTAIL.t10 w_n4474_n1944# sky130_fd_pr__pfet_01v8 ad=0.8052 pd=5.21 as=0.8052 ps=5.21 w=4.88 l=2.59
X16 B.t5 B.t3 B.t4 w_n4474_n1944# sky130_fd_pr__pfet_01v8 ad=1.9032 pd=10.54 as=0 ps=0 w=4.88 l=2.59
X17 VTAIL.t19 VN.t7 VDD2.t2 w_n4474_n1944# sky130_fd_pr__pfet_01v8 ad=0.8052 pd=5.21 as=0.8052 ps=5.21 w=4.88 l=2.59
X18 VTAIL.t3 VN.t8 VDD2.t1 w_n4474_n1944# sky130_fd_pr__pfet_01v8 ad=0.8052 pd=5.21 as=0.8052 ps=5.21 w=4.88 l=2.59
X19 VTAIL.t13 VP.t7 VDD1.t2 w_n4474_n1944# sky130_fd_pr__pfet_01v8 ad=0.8052 pd=5.21 as=0.8052 ps=5.21 w=4.88 l=2.59
X20 B.t2 B.t0 B.t1 w_n4474_n1944# sky130_fd_pr__pfet_01v8 ad=1.9032 pd=10.54 as=0 ps=0 w=4.88 l=2.59
X21 VTAIL.t15 VP.t8 VDD1.t1 w_n4474_n1944# sky130_fd_pr__pfet_01v8 ad=0.8052 pd=5.21 as=0.8052 ps=5.21 w=4.88 l=2.59
X22 VDD1.t0 VP.t9 VTAIL.t8 w_n4474_n1944# sky130_fd_pr__pfet_01v8 ad=1.9032 pd=10.54 as=0.8052 ps=5.21 w=4.88 l=2.59
X23 VTAIL.t2 VN.t9 VDD2.t0 w_n4474_n1944# sky130_fd_pr__pfet_01v8 ad=0.8052 pd=5.21 as=0.8052 ps=5.21 w=4.88 l=2.59
R0 VP.n25 VP.n22 161.3
R1 VP.n27 VP.n26 161.3
R2 VP.n28 VP.n21 161.3
R3 VP.n30 VP.n29 161.3
R4 VP.n31 VP.n20 161.3
R5 VP.n33 VP.n32 161.3
R6 VP.n35 VP.n19 161.3
R7 VP.n37 VP.n36 161.3
R8 VP.n38 VP.n18 161.3
R9 VP.n40 VP.n39 161.3
R10 VP.n41 VP.n17 161.3
R11 VP.n43 VP.n42 161.3
R12 VP.n45 VP.n44 161.3
R13 VP.n46 VP.n15 161.3
R14 VP.n48 VP.n47 161.3
R15 VP.n49 VP.n14 161.3
R16 VP.n51 VP.n50 161.3
R17 VP.n52 VP.n13 161.3
R18 VP.n94 VP.n0 161.3
R19 VP.n93 VP.n92 161.3
R20 VP.n91 VP.n1 161.3
R21 VP.n90 VP.n89 161.3
R22 VP.n88 VP.n2 161.3
R23 VP.n87 VP.n86 161.3
R24 VP.n85 VP.n84 161.3
R25 VP.n83 VP.n4 161.3
R26 VP.n82 VP.n81 161.3
R27 VP.n80 VP.n5 161.3
R28 VP.n79 VP.n78 161.3
R29 VP.n77 VP.n6 161.3
R30 VP.n75 VP.n74 161.3
R31 VP.n73 VP.n7 161.3
R32 VP.n72 VP.n71 161.3
R33 VP.n70 VP.n8 161.3
R34 VP.n69 VP.n68 161.3
R35 VP.n67 VP.n9 161.3
R36 VP.n66 VP.n65 161.3
R37 VP.n63 VP.n10 161.3
R38 VP.n62 VP.n61 161.3
R39 VP.n60 VP.n11 161.3
R40 VP.n59 VP.n58 161.3
R41 VP.n57 VP.n12 161.3
R42 VP.n56 VP.n55 106.481
R43 VP.n96 VP.n95 106.481
R44 VP.n54 VP.n53 106.481
R45 VP.n24 VP.t9 77.2801
R46 VP.n24 VP.n23 64.3558
R47 VP.n71 VP.n70 56.5617
R48 VP.n82 VP.n5 56.5617
R49 VP.n40 VP.n18 56.5617
R50 VP.n29 VP.n28 56.5617
R51 VP.n62 VP.n11 53.171
R52 VP.n89 VP.n1 53.171
R53 VP.n47 VP.n14 53.171
R54 VP.n55 VP.n54 47.5981
R55 VP.n56 VP.t3 45.409
R56 VP.n64 VP.t5 45.409
R57 VP.n76 VP.t2 45.409
R58 VP.n3 VP.t8 45.409
R59 VP.n95 VP.t1 45.409
R60 VP.n53 VP.t0 45.409
R61 VP.n16 VP.t7 45.409
R62 VP.n34 VP.t6 45.409
R63 VP.n23 VP.t4 45.409
R64 VP.n63 VP.n62 27.983
R65 VP.n89 VP.n88 27.983
R66 VP.n47 VP.n46 27.983
R67 VP.n58 VP.n57 24.5923
R68 VP.n58 VP.n11 24.5923
R69 VP.n65 VP.n63 24.5923
R70 VP.n69 VP.n9 24.5923
R71 VP.n70 VP.n69 24.5923
R72 VP.n71 VP.n7 24.5923
R73 VP.n75 VP.n7 24.5923
R74 VP.n78 VP.n77 24.5923
R75 VP.n78 VP.n5 24.5923
R76 VP.n83 VP.n82 24.5923
R77 VP.n84 VP.n83 24.5923
R78 VP.n88 VP.n87 24.5923
R79 VP.n93 VP.n1 24.5923
R80 VP.n94 VP.n93 24.5923
R81 VP.n51 VP.n14 24.5923
R82 VP.n52 VP.n51 24.5923
R83 VP.n41 VP.n40 24.5923
R84 VP.n42 VP.n41 24.5923
R85 VP.n46 VP.n45 24.5923
R86 VP.n29 VP.n20 24.5923
R87 VP.n33 VP.n20 24.5923
R88 VP.n36 VP.n35 24.5923
R89 VP.n36 VP.n18 24.5923
R90 VP.n27 VP.n22 24.5923
R91 VP.n28 VP.n27 24.5923
R92 VP.n65 VP.n64 16.2311
R93 VP.n87 VP.n3 16.2311
R94 VP.n45 VP.n16 16.2311
R95 VP.n76 VP.n75 12.2964
R96 VP.n77 VP.n76 12.2964
R97 VP.n34 VP.n33 12.2964
R98 VP.n35 VP.n34 12.2964
R99 VP.n64 VP.n9 8.36172
R100 VP.n84 VP.n3 8.36172
R101 VP.n42 VP.n16 8.36172
R102 VP.n23 VP.n22 8.36172
R103 VP.n25 VP.n24 7.1827
R104 VP.n57 VP.n56 4.42703
R105 VP.n95 VP.n94 4.42703
R106 VP.n53 VP.n52 4.42703
R107 VP.n54 VP.n13 0.278335
R108 VP.n55 VP.n12 0.278335
R109 VP.n96 VP.n0 0.278335
R110 VP.n26 VP.n25 0.189894
R111 VP.n26 VP.n21 0.189894
R112 VP.n30 VP.n21 0.189894
R113 VP.n31 VP.n30 0.189894
R114 VP.n32 VP.n31 0.189894
R115 VP.n32 VP.n19 0.189894
R116 VP.n37 VP.n19 0.189894
R117 VP.n38 VP.n37 0.189894
R118 VP.n39 VP.n38 0.189894
R119 VP.n39 VP.n17 0.189894
R120 VP.n43 VP.n17 0.189894
R121 VP.n44 VP.n43 0.189894
R122 VP.n44 VP.n15 0.189894
R123 VP.n48 VP.n15 0.189894
R124 VP.n49 VP.n48 0.189894
R125 VP.n50 VP.n49 0.189894
R126 VP.n50 VP.n13 0.189894
R127 VP.n59 VP.n12 0.189894
R128 VP.n60 VP.n59 0.189894
R129 VP.n61 VP.n60 0.189894
R130 VP.n61 VP.n10 0.189894
R131 VP.n66 VP.n10 0.189894
R132 VP.n67 VP.n66 0.189894
R133 VP.n68 VP.n67 0.189894
R134 VP.n68 VP.n8 0.189894
R135 VP.n72 VP.n8 0.189894
R136 VP.n73 VP.n72 0.189894
R137 VP.n74 VP.n73 0.189894
R138 VP.n74 VP.n6 0.189894
R139 VP.n79 VP.n6 0.189894
R140 VP.n80 VP.n79 0.189894
R141 VP.n81 VP.n80 0.189894
R142 VP.n81 VP.n4 0.189894
R143 VP.n85 VP.n4 0.189894
R144 VP.n86 VP.n85 0.189894
R145 VP.n86 VP.n2 0.189894
R146 VP.n90 VP.n2 0.189894
R147 VP.n91 VP.n90 0.189894
R148 VP.n92 VP.n91 0.189894
R149 VP.n92 VP.n0 0.189894
R150 VP VP.n96 0.153485
R151 VTAIL.n11 VTAIL.t4 89.647
R152 VTAIL.n17 VTAIL.t1 89.647
R153 VTAIL.n2 VTAIL.t9 89.647
R154 VTAIL.n16 VTAIL.t11 89.647
R155 VTAIL.n15 VTAIL.n14 82.9862
R156 VTAIL.n13 VTAIL.n12 82.9862
R157 VTAIL.n10 VTAIL.n9 82.9862
R158 VTAIL.n8 VTAIL.n7 82.9862
R159 VTAIL.n19 VTAIL.n18 82.986
R160 VTAIL.n1 VTAIL.n0 82.986
R161 VTAIL.n4 VTAIL.n3 82.986
R162 VTAIL.n6 VTAIL.n5 82.986
R163 VTAIL.n8 VTAIL.n6 21.6083
R164 VTAIL.n17 VTAIL.n16 19.091
R165 VTAIL.n18 VTAIL.t6 6.66136
R166 VTAIL.n18 VTAIL.t2 6.66136
R167 VTAIL.n0 VTAIL.t18 6.66136
R168 VTAIL.n0 VTAIL.t3 6.66136
R169 VTAIL.n3 VTAIL.t16 6.66136
R170 VTAIL.n3 VTAIL.t15 6.66136
R171 VTAIL.n5 VTAIL.t7 6.66136
R172 VTAIL.n5 VTAIL.t12 6.66136
R173 VTAIL.n14 VTAIL.t10 6.66136
R174 VTAIL.n14 VTAIL.t13 6.66136
R175 VTAIL.n12 VTAIL.t8 6.66136
R176 VTAIL.n12 VTAIL.t14 6.66136
R177 VTAIL.n9 VTAIL.t5 6.66136
R178 VTAIL.n9 VTAIL.t19 6.66136
R179 VTAIL.n7 VTAIL.t0 6.66136
R180 VTAIL.n7 VTAIL.t17 6.66136
R181 VTAIL.n10 VTAIL.n8 2.51774
R182 VTAIL.n11 VTAIL.n10 2.51774
R183 VTAIL.n15 VTAIL.n13 2.51774
R184 VTAIL.n16 VTAIL.n15 2.51774
R185 VTAIL.n6 VTAIL.n4 2.51774
R186 VTAIL.n4 VTAIL.n2 2.51774
R187 VTAIL.n19 VTAIL.n17 2.51774
R188 VTAIL VTAIL.n1 1.94662
R189 VTAIL.n13 VTAIL.n11 1.72895
R190 VTAIL.n2 VTAIL.n1 1.72895
R191 VTAIL VTAIL.n19 0.571621
R192 VDD1.n1 VDD1.t0 108.844
R193 VDD1.n3 VDD1.t6 108.843
R194 VDD1.n5 VDD1.n4 101.498
R195 VDD1.n1 VDD1.n0 99.665
R196 VDD1.n7 VDD1.n6 99.6649
R197 VDD1.n3 VDD1.n2 99.6648
R198 VDD1.n7 VDD1.n5 41.7207
R199 VDD1.n6 VDD1.t2 6.66136
R200 VDD1.n6 VDD1.t9 6.66136
R201 VDD1.n0 VDD1.t5 6.66136
R202 VDD1.n0 VDD1.t3 6.66136
R203 VDD1.n4 VDD1.t1 6.66136
R204 VDD1.n4 VDD1.t8 6.66136
R205 VDD1.n2 VDD1.t4 6.66136
R206 VDD1.n2 VDD1.t7 6.66136
R207 VDD1 VDD1.n7 1.83024
R208 VDD1 VDD1.n1 0.688
R209 VDD1.n5 VDD1.n3 0.574464
R210 VN.n81 VN.n42 161.3
R211 VN.n80 VN.n79 161.3
R212 VN.n78 VN.n43 161.3
R213 VN.n77 VN.n76 161.3
R214 VN.n75 VN.n44 161.3
R215 VN.n74 VN.n73 161.3
R216 VN.n72 VN.n71 161.3
R217 VN.n70 VN.n46 161.3
R218 VN.n69 VN.n68 161.3
R219 VN.n67 VN.n47 161.3
R220 VN.n66 VN.n65 161.3
R221 VN.n64 VN.n48 161.3
R222 VN.n62 VN.n61 161.3
R223 VN.n60 VN.n49 161.3
R224 VN.n59 VN.n58 161.3
R225 VN.n57 VN.n50 161.3
R226 VN.n56 VN.n55 161.3
R227 VN.n54 VN.n51 161.3
R228 VN.n39 VN.n0 161.3
R229 VN.n38 VN.n37 161.3
R230 VN.n36 VN.n1 161.3
R231 VN.n35 VN.n34 161.3
R232 VN.n33 VN.n2 161.3
R233 VN.n32 VN.n31 161.3
R234 VN.n30 VN.n29 161.3
R235 VN.n28 VN.n4 161.3
R236 VN.n27 VN.n26 161.3
R237 VN.n25 VN.n5 161.3
R238 VN.n24 VN.n23 161.3
R239 VN.n22 VN.n6 161.3
R240 VN.n20 VN.n19 161.3
R241 VN.n18 VN.n7 161.3
R242 VN.n17 VN.n16 161.3
R243 VN.n15 VN.n8 161.3
R244 VN.n14 VN.n13 161.3
R245 VN.n12 VN.n9 161.3
R246 VN.n41 VN.n40 106.481
R247 VN.n83 VN.n82 106.481
R248 VN.n11 VN.t2 77.2801
R249 VN.n53 VN.t3 77.2801
R250 VN.n11 VN.n10 64.3558
R251 VN.n53 VN.n52 64.3558
R252 VN.n16 VN.n15 56.5617
R253 VN.n27 VN.n5 56.5617
R254 VN.n58 VN.n57 56.5617
R255 VN.n69 VN.n47 56.5617
R256 VN.n34 VN.n1 53.171
R257 VN.n76 VN.n43 53.171
R258 VN VN.n83 47.877
R259 VN.n10 VN.t8 45.409
R260 VN.n21 VN.t5 45.409
R261 VN.n3 VN.t9 45.409
R262 VN.n40 VN.t1 45.409
R263 VN.n52 VN.t7 45.409
R264 VN.n63 VN.t0 45.409
R265 VN.n45 VN.t4 45.409
R266 VN.n82 VN.t6 45.409
R267 VN.n34 VN.n33 27.983
R268 VN.n76 VN.n75 27.983
R269 VN.n14 VN.n9 24.5923
R270 VN.n15 VN.n14 24.5923
R271 VN.n16 VN.n7 24.5923
R272 VN.n20 VN.n7 24.5923
R273 VN.n23 VN.n22 24.5923
R274 VN.n23 VN.n5 24.5923
R275 VN.n28 VN.n27 24.5923
R276 VN.n29 VN.n28 24.5923
R277 VN.n33 VN.n32 24.5923
R278 VN.n38 VN.n1 24.5923
R279 VN.n39 VN.n38 24.5923
R280 VN.n57 VN.n56 24.5923
R281 VN.n56 VN.n51 24.5923
R282 VN.n65 VN.n47 24.5923
R283 VN.n65 VN.n64 24.5923
R284 VN.n62 VN.n49 24.5923
R285 VN.n58 VN.n49 24.5923
R286 VN.n75 VN.n74 24.5923
R287 VN.n71 VN.n70 24.5923
R288 VN.n70 VN.n69 24.5923
R289 VN.n81 VN.n80 24.5923
R290 VN.n80 VN.n43 24.5923
R291 VN.n32 VN.n3 16.2311
R292 VN.n74 VN.n45 16.2311
R293 VN.n21 VN.n20 12.2964
R294 VN.n22 VN.n21 12.2964
R295 VN.n64 VN.n63 12.2964
R296 VN.n63 VN.n62 12.2964
R297 VN.n10 VN.n9 8.36172
R298 VN.n29 VN.n3 8.36172
R299 VN.n52 VN.n51 8.36172
R300 VN.n71 VN.n45 8.36172
R301 VN.n54 VN.n53 7.1827
R302 VN.n12 VN.n11 7.1827
R303 VN.n40 VN.n39 4.42703
R304 VN.n82 VN.n81 4.42703
R305 VN.n83 VN.n42 0.278335
R306 VN.n41 VN.n0 0.278335
R307 VN.n79 VN.n42 0.189894
R308 VN.n79 VN.n78 0.189894
R309 VN.n78 VN.n77 0.189894
R310 VN.n77 VN.n44 0.189894
R311 VN.n73 VN.n44 0.189894
R312 VN.n73 VN.n72 0.189894
R313 VN.n72 VN.n46 0.189894
R314 VN.n68 VN.n46 0.189894
R315 VN.n68 VN.n67 0.189894
R316 VN.n67 VN.n66 0.189894
R317 VN.n66 VN.n48 0.189894
R318 VN.n61 VN.n48 0.189894
R319 VN.n61 VN.n60 0.189894
R320 VN.n60 VN.n59 0.189894
R321 VN.n59 VN.n50 0.189894
R322 VN.n55 VN.n50 0.189894
R323 VN.n55 VN.n54 0.189894
R324 VN.n13 VN.n12 0.189894
R325 VN.n13 VN.n8 0.189894
R326 VN.n17 VN.n8 0.189894
R327 VN.n18 VN.n17 0.189894
R328 VN.n19 VN.n18 0.189894
R329 VN.n19 VN.n6 0.189894
R330 VN.n24 VN.n6 0.189894
R331 VN.n25 VN.n24 0.189894
R332 VN.n26 VN.n25 0.189894
R333 VN.n26 VN.n4 0.189894
R334 VN.n30 VN.n4 0.189894
R335 VN.n31 VN.n30 0.189894
R336 VN.n31 VN.n2 0.189894
R337 VN.n35 VN.n2 0.189894
R338 VN.n36 VN.n35 0.189894
R339 VN.n37 VN.n36 0.189894
R340 VN.n37 VN.n0 0.189894
R341 VN VN.n41 0.153485
R342 VDD2.n1 VDD2.t7 108.843
R343 VDD2.n4 VDD2.t3 106.326
R344 VDD2.n3 VDD2.n2 101.498
R345 VDD2 VDD2.n7 101.495
R346 VDD2.n6 VDD2.n5 99.665
R347 VDD2.n1 VDD2.n0 99.6648
R348 VDD2.n4 VDD2.n3 39.8791
R349 VDD2.n7 VDD2.t2 6.66136
R350 VDD2.n7 VDD2.t6 6.66136
R351 VDD2.n5 VDD2.t5 6.66136
R352 VDD2.n5 VDD2.t9 6.66136
R353 VDD2.n2 VDD2.t0 6.66136
R354 VDD2.n2 VDD2.t8 6.66136
R355 VDD2.n0 VDD2.t1 6.66136
R356 VDD2.n0 VDD2.t4 6.66136
R357 VDD2.n6 VDD2.n4 2.51774
R358 VDD2 VDD2.n6 0.688
R359 VDD2.n3 VDD2.n1 0.574464
R360 B.n345 B.n344 585
R361 B.n343 B.n122 585
R362 B.n342 B.n341 585
R363 B.n340 B.n123 585
R364 B.n339 B.n338 585
R365 B.n337 B.n124 585
R366 B.n336 B.n335 585
R367 B.n334 B.n125 585
R368 B.n333 B.n332 585
R369 B.n331 B.n126 585
R370 B.n330 B.n329 585
R371 B.n328 B.n127 585
R372 B.n327 B.n326 585
R373 B.n325 B.n128 585
R374 B.n324 B.n323 585
R375 B.n322 B.n129 585
R376 B.n321 B.n320 585
R377 B.n319 B.n130 585
R378 B.n318 B.n317 585
R379 B.n316 B.n131 585
R380 B.n315 B.n314 585
R381 B.n313 B.n312 585
R382 B.n311 B.n135 585
R383 B.n310 B.n309 585
R384 B.n308 B.n136 585
R385 B.n307 B.n306 585
R386 B.n305 B.n137 585
R387 B.n304 B.n303 585
R388 B.n302 B.n138 585
R389 B.n301 B.n300 585
R390 B.n298 B.n139 585
R391 B.n297 B.n296 585
R392 B.n295 B.n142 585
R393 B.n294 B.n293 585
R394 B.n292 B.n143 585
R395 B.n291 B.n290 585
R396 B.n289 B.n144 585
R397 B.n288 B.n287 585
R398 B.n286 B.n145 585
R399 B.n285 B.n284 585
R400 B.n283 B.n146 585
R401 B.n282 B.n281 585
R402 B.n280 B.n147 585
R403 B.n279 B.n278 585
R404 B.n277 B.n148 585
R405 B.n276 B.n275 585
R406 B.n274 B.n149 585
R407 B.n273 B.n272 585
R408 B.n271 B.n150 585
R409 B.n270 B.n269 585
R410 B.n268 B.n151 585
R411 B.n346 B.n121 585
R412 B.n348 B.n347 585
R413 B.n349 B.n120 585
R414 B.n351 B.n350 585
R415 B.n352 B.n119 585
R416 B.n354 B.n353 585
R417 B.n355 B.n118 585
R418 B.n357 B.n356 585
R419 B.n358 B.n117 585
R420 B.n360 B.n359 585
R421 B.n361 B.n116 585
R422 B.n363 B.n362 585
R423 B.n364 B.n115 585
R424 B.n366 B.n365 585
R425 B.n367 B.n114 585
R426 B.n369 B.n368 585
R427 B.n370 B.n113 585
R428 B.n372 B.n371 585
R429 B.n373 B.n112 585
R430 B.n375 B.n374 585
R431 B.n376 B.n111 585
R432 B.n378 B.n377 585
R433 B.n379 B.n110 585
R434 B.n381 B.n380 585
R435 B.n382 B.n109 585
R436 B.n384 B.n383 585
R437 B.n385 B.n108 585
R438 B.n387 B.n386 585
R439 B.n388 B.n107 585
R440 B.n390 B.n389 585
R441 B.n391 B.n106 585
R442 B.n393 B.n392 585
R443 B.n394 B.n105 585
R444 B.n396 B.n395 585
R445 B.n397 B.n104 585
R446 B.n399 B.n398 585
R447 B.n400 B.n103 585
R448 B.n402 B.n401 585
R449 B.n403 B.n102 585
R450 B.n405 B.n404 585
R451 B.n406 B.n101 585
R452 B.n408 B.n407 585
R453 B.n409 B.n100 585
R454 B.n411 B.n410 585
R455 B.n412 B.n99 585
R456 B.n414 B.n413 585
R457 B.n415 B.n98 585
R458 B.n417 B.n416 585
R459 B.n418 B.n97 585
R460 B.n420 B.n419 585
R461 B.n421 B.n96 585
R462 B.n423 B.n422 585
R463 B.n424 B.n95 585
R464 B.n426 B.n425 585
R465 B.n427 B.n94 585
R466 B.n429 B.n428 585
R467 B.n430 B.n93 585
R468 B.n432 B.n431 585
R469 B.n433 B.n92 585
R470 B.n435 B.n434 585
R471 B.n436 B.n91 585
R472 B.n438 B.n437 585
R473 B.n439 B.n90 585
R474 B.n441 B.n440 585
R475 B.n442 B.n89 585
R476 B.n444 B.n443 585
R477 B.n445 B.n88 585
R478 B.n447 B.n446 585
R479 B.n448 B.n87 585
R480 B.n450 B.n449 585
R481 B.n451 B.n86 585
R482 B.n453 B.n452 585
R483 B.n454 B.n85 585
R484 B.n456 B.n455 585
R485 B.n457 B.n84 585
R486 B.n459 B.n458 585
R487 B.n460 B.n83 585
R488 B.n462 B.n461 585
R489 B.n463 B.n82 585
R490 B.n465 B.n464 585
R491 B.n466 B.n81 585
R492 B.n468 B.n467 585
R493 B.n469 B.n80 585
R494 B.n471 B.n470 585
R495 B.n472 B.n79 585
R496 B.n474 B.n473 585
R497 B.n475 B.n78 585
R498 B.n477 B.n476 585
R499 B.n478 B.n77 585
R500 B.n480 B.n479 585
R501 B.n481 B.n76 585
R502 B.n483 B.n482 585
R503 B.n484 B.n75 585
R504 B.n486 B.n485 585
R505 B.n487 B.n74 585
R506 B.n489 B.n488 585
R507 B.n490 B.n73 585
R508 B.n492 B.n491 585
R509 B.n493 B.n72 585
R510 B.n495 B.n494 585
R511 B.n496 B.n71 585
R512 B.n498 B.n497 585
R513 B.n499 B.n70 585
R514 B.n501 B.n500 585
R515 B.n502 B.n69 585
R516 B.n504 B.n503 585
R517 B.n505 B.n68 585
R518 B.n507 B.n506 585
R519 B.n508 B.n67 585
R520 B.n510 B.n509 585
R521 B.n511 B.n66 585
R522 B.n513 B.n512 585
R523 B.n514 B.n65 585
R524 B.n516 B.n515 585
R525 B.n517 B.n64 585
R526 B.n519 B.n518 585
R527 B.n520 B.n63 585
R528 B.n522 B.n521 585
R529 B.n523 B.n62 585
R530 B.n525 B.n524 585
R531 B.n603 B.n602 585
R532 B.n601 B.n32 585
R533 B.n600 B.n599 585
R534 B.n598 B.n33 585
R535 B.n597 B.n596 585
R536 B.n595 B.n34 585
R537 B.n594 B.n593 585
R538 B.n592 B.n35 585
R539 B.n591 B.n590 585
R540 B.n589 B.n36 585
R541 B.n588 B.n587 585
R542 B.n586 B.n37 585
R543 B.n585 B.n584 585
R544 B.n583 B.n38 585
R545 B.n582 B.n581 585
R546 B.n580 B.n39 585
R547 B.n579 B.n578 585
R548 B.n577 B.n40 585
R549 B.n576 B.n575 585
R550 B.n574 B.n41 585
R551 B.n573 B.n572 585
R552 B.n571 B.n570 585
R553 B.n569 B.n45 585
R554 B.n568 B.n567 585
R555 B.n566 B.n46 585
R556 B.n565 B.n564 585
R557 B.n563 B.n47 585
R558 B.n562 B.n561 585
R559 B.n560 B.n48 585
R560 B.n559 B.n558 585
R561 B.n556 B.n49 585
R562 B.n555 B.n554 585
R563 B.n553 B.n52 585
R564 B.n552 B.n551 585
R565 B.n550 B.n53 585
R566 B.n549 B.n548 585
R567 B.n547 B.n54 585
R568 B.n546 B.n545 585
R569 B.n544 B.n55 585
R570 B.n543 B.n542 585
R571 B.n541 B.n56 585
R572 B.n540 B.n539 585
R573 B.n538 B.n57 585
R574 B.n537 B.n536 585
R575 B.n535 B.n58 585
R576 B.n534 B.n533 585
R577 B.n532 B.n59 585
R578 B.n531 B.n530 585
R579 B.n529 B.n60 585
R580 B.n528 B.n527 585
R581 B.n526 B.n61 585
R582 B.n604 B.n31 585
R583 B.n606 B.n605 585
R584 B.n607 B.n30 585
R585 B.n609 B.n608 585
R586 B.n610 B.n29 585
R587 B.n612 B.n611 585
R588 B.n613 B.n28 585
R589 B.n615 B.n614 585
R590 B.n616 B.n27 585
R591 B.n618 B.n617 585
R592 B.n619 B.n26 585
R593 B.n621 B.n620 585
R594 B.n622 B.n25 585
R595 B.n624 B.n623 585
R596 B.n625 B.n24 585
R597 B.n627 B.n626 585
R598 B.n628 B.n23 585
R599 B.n630 B.n629 585
R600 B.n631 B.n22 585
R601 B.n633 B.n632 585
R602 B.n634 B.n21 585
R603 B.n636 B.n635 585
R604 B.n637 B.n20 585
R605 B.n639 B.n638 585
R606 B.n640 B.n19 585
R607 B.n642 B.n641 585
R608 B.n643 B.n18 585
R609 B.n645 B.n644 585
R610 B.n646 B.n17 585
R611 B.n648 B.n647 585
R612 B.n649 B.n16 585
R613 B.n651 B.n650 585
R614 B.n652 B.n15 585
R615 B.n654 B.n653 585
R616 B.n655 B.n14 585
R617 B.n657 B.n656 585
R618 B.n658 B.n13 585
R619 B.n660 B.n659 585
R620 B.n661 B.n12 585
R621 B.n663 B.n662 585
R622 B.n664 B.n11 585
R623 B.n666 B.n665 585
R624 B.n667 B.n10 585
R625 B.n669 B.n668 585
R626 B.n670 B.n9 585
R627 B.n672 B.n671 585
R628 B.n673 B.n8 585
R629 B.n675 B.n674 585
R630 B.n676 B.n7 585
R631 B.n678 B.n677 585
R632 B.n679 B.n6 585
R633 B.n681 B.n680 585
R634 B.n682 B.n5 585
R635 B.n684 B.n683 585
R636 B.n685 B.n4 585
R637 B.n687 B.n686 585
R638 B.n688 B.n3 585
R639 B.n690 B.n689 585
R640 B.n691 B.n0 585
R641 B.n2 B.n1 585
R642 B.n181 B.n180 585
R643 B.n183 B.n182 585
R644 B.n184 B.n179 585
R645 B.n186 B.n185 585
R646 B.n187 B.n178 585
R647 B.n189 B.n188 585
R648 B.n190 B.n177 585
R649 B.n192 B.n191 585
R650 B.n193 B.n176 585
R651 B.n195 B.n194 585
R652 B.n196 B.n175 585
R653 B.n198 B.n197 585
R654 B.n199 B.n174 585
R655 B.n201 B.n200 585
R656 B.n202 B.n173 585
R657 B.n204 B.n203 585
R658 B.n205 B.n172 585
R659 B.n207 B.n206 585
R660 B.n208 B.n171 585
R661 B.n210 B.n209 585
R662 B.n211 B.n170 585
R663 B.n213 B.n212 585
R664 B.n214 B.n169 585
R665 B.n216 B.n215 585
R666 B.n217 B.n168 585
R667 B.n219 B.n218 585
R668 B.n220 B.n167 585
R669 B.n222 B.n221 585
R670 B.n223 B.n166 585
R671 B.n225 B.n224 585
R672 B.n226 B.n165 585
R673 B.n228 B.n227 585
R674 B.n229 B.n164 585
R675 B.n231 B.n230 585
R676 B.n232 B.n163 585
R677 B.n234 B.n233 585
R678 B.n235 B.n162 585
R679 B.n237 B.n236 585
R680 B.n238 B.n161 585
R681 B.n240 B.n239 585
R682 B.n241 B.n160 585
R683 B.n243 B.n242 585
R684 B.n244 B.n159 585
R685 B.n246 B.n245 585
R686 B.n247 B.n158 585
R687 B.n249 B.n248 585
R688 B.n250 B.n157 585
R689 B.n252 B.n251 585
R690 B.n253 B.n156 585
R691 B.n255 B.n254 585
R692 B.n256 B.n155 585
R693 B.n258 B.n257 585
R694 B.n259 B.n154 585
R695 B.n261 B.n260 585
R696 B.n262 B.n153 585
R697 B.n264 B.n263 585
R698 B.n265 B.n152 585
R699 B.n267 B.n266 585
R700 B.n266 B.n151 516.524
R701 B.n344 B.n121 516.524
R702 B.n524 B.n61 516.524
R703 B.n602 B.n31 516.524
R704 B.n693 B.n692 256.663
R705 B.n140 B.t3 253.44
R706 B.n132 B.t0 253.44
R707 B.n50 B.t6 253.44
R708 B.n42 B.t9 253.44
R709 B.n692 B.n691 235.042
R710 B.n692 B.n2 235.042
R711 B.n132 B.t1 173.637
R712 B.n50 B.t8 173.637
R713 B.n140 B.t4 173.632
R714 B.n42 B.t11 173.632
R715 B.n270 B.n151 163.367
R716 B.n271 B.n270 163.367
R717 B.n272 B.n271 163.367
R718 B.n272 B.n149 163.367
R719 B.n276 B.n149 163.367
R720 B.n277 B.n276 163.367
R721 B.n278 B.n277 163.367
R722 B.n278 B.n147 163.367
R723 B.n282 B.n147 163.367
R724 B.n283 B.n282 163.367
R725 B.n284 B.n283 163.367
R726 B.n284 B.n145 163.367
R727 B.n288 B.n145 163.367
R728 B.n289 B.n288 163.367
R729 B.n290 B.n289 163.367
R730 B.n290 B.n143 163.367
R731 B.n294 B.n143 163.367
R732 B.n295 B.n294 163.367
R733 B.n296 B.n295 163.367
R734 B.n296 B.n139 163.367
R735 B.n301 B.n139 163.367
R736 B.n302 B.n301 163.367
R737 B.n303 B.n302 163.367
R738 B.n303 B.n137 163.367
R739 B.n307 B.n137 163.367
R740 B.n308 B.n307 163.367
R741 B.n309 B.n308 163.367
R742 B.n309 B.n135 163.367
R743 B.n313 B.n135 163.367
R744 B.n314 B.n313 163.367
R745 B.n314 B.n131 163.367
R746 B.n318 B.n131 163.367
R747 B.n319 B.n318 163.367
R748 B.n320 B.n319 163.367
R749 B.n320 B.n129 163.367
R750 B.n324 B.n129 163.367
R751 B.n325 B.n324 163.367
R752 B.n326 B.n325 163.367
R753 B.n326 B.n127 163.367
R754 B.n330 B.n127 163.367
R755 B.n331 B.n330 163.367
R756 B.n332 B.n331 163.367
R757 B.n332 B.n125 163.367
R758 B.n336 B.n125 163.367
R759 B.n337 B.n336 163.367
R760 B.n338 B.n337 163.367
R761 B.n338 B.n123 163.367
R762 B.n342 B.n123 163.367
R763 B.n343 B.n342 163.367
R764 B.n344 B.n343 163.367
R765 B.n524 B.n523 163.367
R766 B.n523 B.n522 163.367
R767 B.n522 B.n63 163.367
R768 B.n518 B.n63 163.367
R769 B.n518 B.n517 163.367
R770 B.n517 B.n516 163.367
R771 B.n516 B.n65 163.367
R772 B.n512 B.n65 163.367
R773 B.n512 B.n511 163.367
R774 B.n511 B.n510 163.367
R775 B.n510 B.n67 163.367
R776 B.n506 B.n67 163.367
R777 B.n506 B.n505 163.367
R778 B.n505 B.n504 163.367
R779 B.n504 B.n69 163.367
R780 B.n500 B.n69 163.367
R781 B.n500 B.n499 163.367
R782 B.n499 B.n498 163.367
R783 B.n498 B.n71 163.367
R784 B.n494 B.n71 163.367
R785 B.n494 B.n493 163.367
R786 B.n493 B.n492 163.367
R787 B.n492 B.n73 163.367
R788 B.n488 B.n73 163.367
R789 B.n488 B.n487 163.367
R790 B.n487 B.n486 163.367
R791 B.n486 B.n75 163.367
R792 B.n482 B.n75 163.367
R793 B.n482 B.n481 163.367
R794 B.n481 B.n480 163.367
R795 B.n480 B.n77 163.367
R796 B.n476 B.n77 163.367
R797 B.n476 B.n475 163.367
R798 B.n475 B.n474 163.367
R799 B.n474 B.n79 163.367
R800 B.n470 B.n79 163.367
R801 B.n470 B.n469 163.367
R802 B.n469 B.n468 163.367
R803 B.n468 B.n81 163.367
R804 B.n464 B.n81 163.367
R805 B.n464 B.n463 163.367
R806 B.n463 B.n462 163.367
R807 B.n462 B.n83 163.367
R808 B.n458 B.n83 163.367
R809 B.n458 B.n457 163.367
R810 B.n457 B.n456 163.367
R811 B.n456 B.n85 163.367
R812 B.n452 B.n85 163.367
R813 B.n452 B.n451 163.367
R814 B.n451 B.n450 163.367
R815 B.n450 B.n87 163.367
R816 B.n446 B.n87 163.367
R817 B.n446 B.n445 163.367
R818 B.n445 B.n444 163.367
R819 B.n444 B.n89 163.367
R820 B.n440 B.n89 163.367
R821 B.n440 B.n439 163.367
R822 B.n439 B.n438 163.367
R823 B.n438 B.n91 163.367
R824 B.n434 B.n91 163.367
R825 B.n434 B.n433 163.367
R826 B.n433 B.n432 163.367
R827 B.n432 B.n93 163.367
R828 B.n428 B.n93 163.367
R829 B.n428 B.n427 163.367
R830 B.n427 B.n426 163.367
R831 B.n426 B.n95 163.367
R832 B.n422 B.n95 163.367
R833 B.n422 B.n421 163.367
R834 B.n421 B.n420 163.367
R835 B.n420 B.n97 163.367
R836 B.n416 B.n97 163.367
R837 B.n416 B.n415 163.367
R838 B.n415 B.n414 163.367
R839 B.n414 B.n99 163.367
R840 B.n410 B.n99 163.367
R841 B.n410 B.n409 163.367
R842 B.n409 B.n408 163.367
R843 B.n408 B.n101 163.367
R844 B.n404 B.n101 163.367
R845 B.n404 B.n403 163.367
R846 B.n403 B.n402 163.367
R847 B.n402 B.n103 163.367
R848 B.n398 B.n103 163.367
R849 B.n398 B.n397 163.367
R850 B.n397 B.n396 163.367
R851 B.n396 B.n105 163.367
R852 B.n392 B.n105 163.367
R853 B.n392 B.n391 163.367
R854 B.n391 B.n390 163.367
R855 B.n390 B.n107 163.367
R856 B.n386 B.n107 163.367
R857 B.n386 B.n385 163.367
R858 B.n385 B.n384 163.367
R859 B.n384 B.n109 163.367
R860 B.n380 B.n109 163.367
R861 B.n380 B.n379 163.367
R862 B.n379 B.n378 163.367
R863 B.n378 B.n111 163.367
R864 B.n374 B.n111 163.367
R865 B.n374 B.n373 163.367
R866 B.n373 B.n372 163.367
R867 B.n372 B.n113 163.367
R868 B.n368 B.n113 163.367
R869 B.n368 B.n367 163.367
R870 B.n367 B.n366 163.367
R871 B.n366 B.n115 163.367
R872 B.n362 B.n115 163.367
R873 B.n362 B.n361 163.367
R874 B.n361 B.n360 163.367
R875 B.n360 B.n117 163.367
R876 B.n356 B.n117 163.367
R877 B.n356 B.n355 163.367
R878 B.n355 B.n354 163.367
R879 B.n354 B.n119 163.367
R880 B.n350 B.n119 163.367
R881 B.n350 B.n349 163.367
R882 B.n349 B.n348 163.367
R883 B.n348 B.n121 163.367
R884 B.n602 B.n601 163.367
R885 B.n601 B.n600 163.367
R886 B.n600 B.n33 163.367
R887 B.n596 B.n33 163.367
R888 B.n596 B.n595 163.367
R889 B.n595 B.n594 163.367
R890 B.n594 B.n35 163.367
R891 B.n590 B.n35 163.367
R892 B.n590 B.n589 163.367
R893 B.n589 B.n588 163.367
R894 B.n588 B.n37 163.367
R895 B.n584 B.n37 163.367
R896 B.n584 B.n583 163.367
R897 B.n583 B.n582 163.367
R898 B.n582 B.n39 163.367
R899 B.n578 B.n39 163.367
R900 B.n578 B.n577 163.367
R901 B.n577 B.n576 163.367
R902 B.n576 B.n41 163.367
R903 B.n572 B.n41 163.367
R904 B.n572 B.n571 163.367
R905 B.n571 B.n45 163.367
R906 B.n567 B.n45 163.367
R907 B.n567 B.n566 163.367
R908 B.n566 B.n565 163.367
R909 B.n565 B.n47 163.367
R910 B.n561 B.n47 163.367
R911 B.n561 B.n560 163.367
R912 B.n560 B.n559 163.367
R913 B.n559 B.n49 163.367
R914 B.n554 B.n49 163.367
R915 B.n554 B.n553 163.367
R916 B.n553 B.n552 163.367
R917 B.n552 B.n53 163.367
R918 B.n548 B.n53 163.367
R919 B.n548 B.n547 163.367
R920 B.n547 B.n546 163.367
R921 B.n546 B.n55 163.367
R922 B.n542 B.n55 163.367
R923 B.n542 B.n541 163.367
R924 B.n541 B.n540 163.367
R925 B.n540 B.n57 163.367
R926 B.n536 B.n57 163.367
R927 B.n536 B.n535 163.367
R928 B.n535 B.n534 163.367
R929 B.n534 B.n59 163.367
R930 B.n530 B.n59 163.367
R931 B.n530 B.n529 163.367
R932 B.n529 B.n528 163.367
R933 B.n528 B.n61 163.367
R934 B.n606 B.n31 163.367
R935 B.n607 B.n606 163.367
R936 B.n608 B.n607 163.367
R937 B.n608 B.n29 163.367
R938 B.n612 B.n29 163.367
R939 B.n613 B.n612 163.367
R940 B.n614 B.n613 163.367
R941 B.n614 B.n27 163.367
R942 B.n618 B.n27 163.367
R943 B.n619 B.n618 163.367
R944 B.n620 B.n619 163.367
R945 B.n620 B.n25 163.367
R946 B.n624 B.n25 163.367
R947 B.n625 B.n624 163.367
R948 B.n626 B.n625 163.367
R949 B.n626 B.n23 163.367
R950 B.n630 B.n23 163.367
R951 B.n631 B.n630 163.367
R952 B.n632 B.n631 163.367
R953 B.n632 B.n21 163.367
R954 B.n636 B.n21 163.367
R955 B.n637 B.n636 163.367
R956 B.n638 B.n637 163.367
R957 B.n638 B.n19 163.367
R958 B.n642 B.n19 163.367
R959 B.n643 B.n642 163.367
R960 B.n644 B.n643 163.367
R961 B.n644 B.n17 163.367
R962 B.n648 B.n17 163.367
R963 B.n649 B.n648 163.367
R964 B.n650 B.n649 163.367
R965 B.n650 B.n15 163.367
R966 B.n654 B.n15 163.367
R967 B.n655 B.n654 163.367
R968 B.n656 B.n655 163.367
R969 B.n656 B.n13 163.367
R970 B.n660 B.n13 163.367
R971 B.n661 B.n660 163.367
R972 B.n662 B.n661 163.367
R973 B.n662 B.n11 163.367
R974 B.n666 B.n11 163.367
R975 B.n667 B.n666 163.367
R976 B.n668 B.n667 163.367
R977 B.n668 B.n9 163.367
R978 B.n672 B.n9 163.367
R979 B.n673 B.n672 163.367
R980 B.n674 B.n673 163.367
R981 B.n674 B.n7 163.367
R982 B.n678 B.n7 163.367
R983 B.n679 B.n678 163.367
R984 B.n680 B.n679 163.367
R985 B.n680 B.n5 163.367
R986 B.n684 B.n5 163.367
R987 B.n685 B.n684 163.367
R988 B.n686 B.n685 163.367
R989 B.n686 B.n3 163.367
R990 B.n690 B.n3 163.367
R991 B.n691 B.n690 163.367
R992 B.n181 B.n2 163.367
R993 B.n182 B.n181 163.367
R994 B.n182 B.n179 163.367
R995 B.n186 B.n179 163.367
R996 B.n187 B.n186 163.367
R997 B.n188 B.n187 163.367
R998 B.n188 B.n177 163.367
R999 B.n192 B.n177 163.367
R1000 B.n193 B.n192 163.367
R1001 B.n194 B.n193 163.367
R1002 B.n194 B.n175 163.367
R1003 B.n198 B.n175 163.367
R1004 B.n199 B.n198 163.367
R1005 B.n200 B.n199 163.367
R1006 B.n200 B.n173 163.367
R1007 B.n204 B.n173 163.367
R1008 B.n205 B.n204 163.367
R1009 B.n206 B.n205 163.367
R1010 B.n206 B.n171 163.367
R1011 B.n210 B.n171 163.367
R1012 B.n211 B.n210 163.367
R1013 B.n212 B.n211 163.367
R1014 B.n212 B.n169 163.367
R1015 B.n216 B.n169 163.367
R1016 B.n217 B.n216 163.367
R1017 B.n218 B.n217 163.367
R1018 B.n218 B.n167 163.367
R1019 B.n222 B.n167 163.367
R1020 B.n223 B.n222 163.367
R1021 B.n224 B.n223 163.367
R1022 B.n224 B.n165 163.367
R1023 B.n228 B.n165 163.367
R1024 B.n229 B.n228 163.367
R1025 B.n230 B.n229 163.367
R1026 B.n230 B.n163 163.367
R1027 B.n234 B.n163 163.367
R1028 B.n235 B.n234 163.367
R1029 B.n236 B.n235 163.367
R1030 B.n236 B.n161 163.367
R1031 B.n240 B.n161 163.367
R1032 B.n241 B.n240 163.367
R1033 B.n242 B.n241 163.367
R1034 B.n242 B.n159 163.367
R1035 B.n246 B.n159 163.367
R1036 B.n247 B.n246 163.367
R1037 B.n248 B.n247 163.367
R1038 B.n248 B.n157 163.367
R1039 B.n252 B.n157 163.367
R1040 B.n253 B.n252 163.367
R1041 B.n254 B.n253 163.367
R1042 B.n254 B.n155 163.367
R1043 B.n258 B.n155 163.367
R1044 B.n259 B.n258 163.367
R1045 B.n260 B.n259 163.367
R1046 B.n260 B.n153 163.367
R1047 B.n264 B.n153 163.367
R1048 B.n265 B.n264 163.367
R1049 B.n266 B.n265 163.367
R1050 B.n133 B.t2 117.007
R1051 B.n51 B.t7 117.007
R1052 B.n141 B.t5 117.002
R1053 B.n43 B.t10 117.002
R1054 B.n299 B.n141 59.5399
R1055 B.n134 B.n133 59.5399
R1056 B.n557 B.n51 59.5399
R1057 B.n44 B.n43 59.5399
R1058 B.n141 B.n140 56.6308
R1059 B.n133 B.n132 56.6308
R1060 B.n51 B.n50 56.6308
R1061 B.n43 B.n42 56.6308
R1062 B.n604 B.n603 33.5615
R1063 B.n526 B.n525 33.5615
R1064 B.n346 B.n345 33.5615
R1065 B.n268 B.n267 33.5615
R1066 B B.n693 18.0485
R1067 B.n605 B.n604 10.6151
R1068 B.n605 B.n30 10.6151
R1069 B.n609 B.n30 10.6151
R1070 B.n610 B.n609 10.6151
R1071 B.n611 B.n610 10.6151
R1072 B.n611 B.n28 10.6151
R1073 B.n615 B.n28 10.6151
R1074 B.n616 B.n615 10.6151
R1075 B.n617 B.n616 10.6151
R1076 B.n617 B.n26 10.6151
R1077 B.n621 B.n26 10.6151
R1078 B.n622 B.n621 10.6151
R1079 B.n623 B.n622 10.6151
R1080 B.n623 B.n24 10.6151
R1081 B.n627 B.n24 10.6151
R1082 B.n628 B.n627 10.6151
R1083 B.n629 B.n628 10.6151
R1084 B.n629 B.n22 10.6151
R1085 B.n633 B.n22 10.6151
R1086 B.n634 B.n633 10.6151
R1087 B.n635 B.n634 10.6151
R1088 B.n635 B.n20 10.6151
R1089 B.n639 B.n20 10.6151
R1090 B.n640 B.n639 10.6151
R1091 B.n641 B.n640 10.6151
R1092 B.n641 B.n18 10.6151
R1093 B.n645 B.n18 10.6151
R1094 B.n646 B.n645 10.6151
R1095 B.n647 B.n646 10.6151
R1096 B.n647 B.n16 10.6151
R1097 B.n651 B.n16 10.6151
R1098 B.n652 B.n651 10.6151
R1099 B.n653 B.n652 10.6151
R1100 B.n653 B.n14 10.6151
R1101 B.n657 B.n14 10.6151
R1102 B.n658 B.n657 10.6151
R1103 B.n659 B.n658 10.6151
R1104 B.n659 B.n12 10.6151
R1105 B.n663 B.n12 10.6151
R1106 B.n664 B.n663 10.6151
R1107 B.n665 B.n664 10.6151
R1108 B.n665 B.n10 10.6151
R1109 B.n669 B.n10 10.6151
R1110 B.n670 B.n669 10.6151
R1111 B.n671 B.n670 10.6151
R1112 B.n671 B.n8 10.6151
R1113 B.n675 B.n8 10.6151
R1114 B.n676 B.n675 10.6151
R1115 B.n677 B.n676 10.6151
R1116 B.n677 B.n6 10.6151
R1117 B.n681 B.n6 10.6151
R1118 B.n682 B.n681 10.6151
R1119 B.n683 B.n682 10.6151
R1120 B.n683 B.n4 10.6151
R1121 B.n687 B.n4 10.6151
R1122 B.n688 B.n687 10.6151
R1123 B.n689 B.n688 10.6151
R1124 B.n689 B.n0 10.6151
R1125 B.n603 B.n32 10.6151
R1126 B.n599 B.n32 10.6151
R1127 B.n599 B.n598 10.6151
R1128 B.n598 B.n597 10.6151
R1129 B.n597 B.n34 10.6151
R1130 B.n593 B.n34 10.6151
R1131 B.n593 B.n592 10.6151
R1132 B.n592 B.n591 10.6151
R1133 B.n591 B.n36 10.6151
R1134 B.n587 B.n36 10.6151
R1135 B.n587 B.n586 10.6151
R1136 B.n586 B.n585 10.6151
R1137 B.n585 B.n38 10.6151
R1138 B.n581 B.n38 10.6151
R1139 B.n581 B.n580 10.6151
R1140 B.n580 B.n579 10.6151
R1141 B.n579 B.n40 10.6151
R1142 B.n575 B.n40 10.6151
R1143 B.n575 B.n574 10.6151
R1144 B.n574 B.n573 10.6151
R1145 B.n570 B.n569 10.6151
R1146 B.n569 B.n568 10.6151
R1147 B.n568 B.n46 10.6151
R1148 B.n564 B.n46 10.6151
R1149 B.n564 B.n563 10.6151
R1150 B.n563 B.n562 10.6151
R1151 B.n562 B.n48 10.6151
R1152 B.n558 B.n48 10.6151
R1153 B.n556 B.n555 10.6151
R1154 B.n555 B.n52 10.6151
R1155 B.n551 B.n52 10.6151
R1156 B.n551 B.n550 10.6151
R1157 B.n550 B.n549 10.6151
R1158 B.n549 B.n54 10.6151
R1159 B.n545 B.n54 10.6151
R1160 B.n545 B.n544 10.6151
R1161 B.n544 B.n543 10.6151
R1162 B.n543 B.n56 10.6151
R1163 B.n539 B.n56 10.6151
R1164 B.n539 B.n538 10.6151
R1165 B.n538 B.n537 10.6151
R1166 B.n537 B.n58 10.6151
R1167 B.n533 B.n58 10.6151
R1168 B.n533 B.n532 10.6151
R1169 B.n532 B.n531 10.6151
R1170 B.n531 B.n60 10.6151
R1171 B.n527 B.n60 10.6151
R1172 B.n527 B.n526 10.6151
R1173 B.n525 B.n62 10.6151
R1174 B.n521 B.n62 10.6151
R1175 B.n521 B.n520 10.6151
R1176 B.n520 B.n519 10.6151
R1177 B.n519 B.n64 10.6151
R1178 B.n515 B.n64 10.6151
R1179 B.n515 B.n514 10.6151
R1180 B.n514 B.n513 10.6151
R1181 B.n513 B.n66 10.6151
R1182 B.n509 B.n66 10.6151
R1183 B.n509 B.n508 10.6151
R1184 B.n508 B.n507 10.6151
R1185 B.n507 B.n68 10.6151
R1186 B.n503 B.n68 10.6151
R1187 B.n503 B.n502 10.6151
R1188 B.n502 B.n501 10.6151
R1189 B.n501 B.n70 10.6151
R1190 B.n497 B.n70 10.6151
R1191 B.n497 B.n496 10.6151
R1192 B.n496 B.n495 10.6151
R1193 B.n495 B.n72 10.6151
R1194 B.n491 B.n72 10.6151
R1195 B.n491 B.n490 10.6151
R1196 B.n490 B.n489 10.6151
R1197 B.n489 B.n74 10.6151
R1198 B.n485 B.n74 10.6151
R1199 B.n485 B.n484 10.6151
R1200 B.n484 B.n483 10.6151
R1201 B.n483 B.n76 10.6151
R1202 B.n479 B.n76 10.6151
R1203 B.n479 B.n478 10.6151
R1204 B.n478 B.n477 10.6151
R1205 B.n477 B.n78 10.6151
R1206 B.n473 B.n78 10.6151
R1207 B.n473 B.n472 10.6151
R1208 B.n472 B.n471 10.6151
R1209 B.n471 B.n80 10.6151
R1210 B.n467 B.n80 10.6151
R1211 B.n467 B.n466 10.6151
R1212 B.n466 B.n465 10.6151
R1213 B.n465 B.n82 10.6151
R1214 B.n461 B.n82 10.6151
R1215 B.n461 B.n460 10.6151
R1216 B.n460 B.n459 10.6151
R1217 B.n459 B.n84 10.6151
R1218 B.n455 B.n84 10.6151
R1219 B.n455 B.n454 10.6151
R1220 B.n454 B.n453 10.6151
R1221 B.n453 B.n86 10.6151
R1222 B.n449 B.n86 10.6151
R1223 B.n449 B.n448 10.6151
R1224 B.n448 B.n447 10.6151
R1225 B.n447 B.n88 10.6151
R1226 B.n443 B.n88 10.6151
R1227 B.n443 B.n442 10.6151
R1228 B.n442 B.n441 10.6151
R1229 B.n441 B.n90 10.6151
R1230 B.n437 B.n90 10.6151
R1231 B.n437 B.n436 10.6151
R1232 B.n436 B.n435 10.6151
R1233 B.n435 B.n92 10.6151
R1234 B.n431 B.n92 10.6151
R1235 B.n431 B.n430 10.6151
R1236 B.n430 B.n429 10.6151
R1237 B.n429 B.n94 10.6151
R1238 B.n425 B.n94 10.6151
R1239 B.n425 B.n424 10.6151
R1240 B.n424 B.n423 10.6151
R1241 B.n423 B.n96 10.6151
R1242 B.n419 B.n96 10.6151
R1243 B.n419 B.n418 10.6151
R1244 B.n418 B.n417 10.6151
R1245 B.n417 B.n98 10.6151
R1246 B.n413 B.n98 10.6151
R1247 B.n413 B.n412 10.6151
R1248 B.n412 B.n411 10.6151
R1249 B.n411 B.n100 10.6151
R1250 B.n407 B.n100 10.6151
R1251 B.n407 B.n406 10.6151
R1252 B.n406 B.n405 10.6151
R1253 B.n405 B.n102 10.6151
R1254 B.n401 B.n102 10.6151
R1255 B.n401 B.n400 10.6151
R1256 B.n400 B.n399 10.6151
R1257 B.n399 B.n104 10.6151
R1258 B.n395 B.n104 10.6151
R1259 B.n395 B.n394 10.6151
R1260 B.n394 B.n393 10.6151
R1261 B.n393 B.n106 10.6151
R1262 B.n389 B.n106 10.6151
R1263 B.n389 B.n388 10.6151
R1264 B.n388 B.n387 10.6151
R1265 B.n387 B.n108 10.6151
R1266 B.n383 B.n108 10.6151
R1267 B.n383 B.n382 10.6151
R1268 B.n382 B.n381 10.6151
R1269 B.n381 B.n110 10.6151
R1270 B.n377 B.n110 10.6151
R1271 B.n377 B.n376 10.6151
R1272 B.n376 B.n375 10.6151
R1273 B.n375 B.n112 10.6151
R1274 B.n371 B.n112 10.6151
R1275 B.n371 B.n370 10.6151
R1276 B.n370 B.n369 10.6151
R1277 B.n369 B.n114 10.6151
R1278 B.n365 B.n114 10.6151
R1279 B.n365 B.n364 10.6151
R1280 B.n364 B.n363 10.6151
R1281 B.n363 B.n116 10.6151
R1282 B.n359 B.n116 10.6151
R1283 B.n359 B.n358 10.6151
R1284 B.n358 B.n357 10.6151
R1285 B.n357 B.n118 10.6151
R1286 B.n353 B.n118 10.6151
R1287 B.n353 B.n352 10.6151
R1288 B.n352 B.n351 10.6151
R1289 B.n351 B.n120 10.6151
R1290 B.n347 B.n120 10.6151
R1291 B.n347 B.n346 10.6151
R1292 B.n180 B.n1 10.6151
R1293 B.n183 B.n180 10.6151
R1294 B.n184 B.n183 10.6151
R1295 B.n185 B.n184 10.6151
R1296 B.n185 B.n178 10.6151
R1297 B.n189 B.n178 10.6151
R1298 B.n190 B.n189 10.6151
R1299 B.n191 B.n190 10.6151
R1300 B.n191 B.n176 10.6151
R1301 B.n195 B.n176 10.6151
R1302 B.n196 B.n195 10.6151
R1303 B.n197 B.n196 10.6151
R1304 B.n197 B.n174 10.6151
R1305 B.n201 B.n174 10.6151
R1306 B.n202 B.n201 10.6151
R1307 B.n203 B.n202 10.6151
R1308 B.n203 B.n172 10.6151
R1309 B.n207 B.n172 10.6151
R1310 B.n208 B.n207 10.6151
R1311 B.n209 B.n208 10.6151
R1312 B.n209 B.n170 10.6151
R1313 B.n213 B.n170 10.6151
R1314 B.n214 B.n213 10.6151
R1315 B.n215 B.n214 10.6151
R1316 B.n215 B.n168 10.6151
R1317 B.n219 B.n168 10.6151
R1318 B.n220 B.n219 10.6151
R1319 B.n221 B.n220 10.6151
R1320 B.n221 B.n166 10.6151
R1321 B.n225 B.n166 10.6151
R1322 B.n226 B.n225 10.6151
R1323 B.n227 B.n226 10.6151
R1324 B.n227 B.n164 10.6151
R1325 B.n231 B.n164 10.6151
R1326 B.n232 B.n231 10.6151
R1327 B.n233 B.n232 10.6151
R1328 B.n233 B.n162 10.6151
R1329 B.n237 B.n162 10.6151
R1330 B.n238 B.n237 10.6151
R1331 B.n239 B.n238 10.6151
R1332 B.n239 B.n160 10.6151
R1333 B.n243 B.n160 10.6151
R1334 B.n244 B.n243 10.6151
R1335 B.n245 B.n244 10.6151
R1336 B.n245 B.n158 10.6151
R1337 B.n249 B.n158 10.6151
R1338 B.n250 B.n249 10.6151
R1339 B.n251 B.n250 10.6151
R1340 B.n251 B.n156 10.6151
R1341 B.n255 B.n156 10.6151
R1342 B.n256 B.n255 10.6151
R1343 B.n257 B.n256 10.6151
R1344 B.n257 B.n154 10.6151
R1345 B.n261 B.n154 10.6151
R1346 B.n262 B.n261 10.6151
R1347 B.n263 B.n262 10.6151
R1348 B.n263 B.n152 10.6151
R1349 B.n267 B.n152 10.6151
R1350 B.n269 B.n268 10.6151
R1351 B.n269 B.n150 10.6151
R1352 B.n273 B.n150 10.6151
R1353 B.n274 B.n273 10.6151
R1354 B.n275 B.n274 10.6151
R1355 B.n275 B.n148 10.6151
R1356 B.n279 B.n148 10.6151
R1357 B.n280 B.n279 10.6151
R1358 B.n281 B.n280 10.6151
R1359 B.n281 B.n146 10.6151
R1360 B.n285 B.n146 10.6151
R1361 B.n286 B.n285 10.6151
R1362 B.n287 B.n286 10.6151
R1363 B.n287 B.n144 10.6151
R1364 B.n291 B.n144 10.6151
R1365 B.n292 B.n291 10.6151
R1366 B.n293 B.n292 10.6151
R1367 B.n293 B.n142 10.6151
R1368 B.n297 B.n142 10.6151
R1369 B.n298 B.n297 10.6151
R1370 B.n300 B.n138 10.6151
R1371 B.n304 B.n138 10.6151
R1372 B.n305 B.n304 10.6151
R1373 B.n306 B.n305 10.6151
R1374 B.n306 B.n136 10.6151
R1375 B.n310 B.n136 10.6151
R1376 B.n311 B.n310 10.6151
R1377 B.n312 B.n311 10.6151
R1378 B.n316 B.n315 10.6151
R1379 B.n317 B.n316 10.6151
R1380 B.n317 B.n130 10.6151
R1381 B.n321 B.n130 10.6151
R1382 B.n322 B.n321 10.6151
R1383 B.n323 B.n322 10.6151
R1384 B.n323 B.n128 10.6151
R1385 B.n327 B.n128 10.6151
R1386 B.n328 B.n327 10.6151
R1387 B.n329 B.n328 10.6151
R1388 B.n329 B.n126 10.6151
R1389 B.n333 B.n126 10.6151
R1390 B.n334 B.n333 10.6151
R1391 B.n335 B.n334 10.6151
R1392 B.n335 B.n124 10.6151
R1393 B.n339 B.n124 10.6151
R1394 B.n340 B.n339 10.6151
R1395 B.n341 B.n340 10.6151
R1396 B.n341 B.n122 10.6151
R1397 B.n345 B.n122 10.6151
R1398 B.n693 B.n0 8.11757
R1399 B.n693 B.n1 8.11757
R1400 B.n570 B.n44 6.5566
R1401 B.n558 B.n557 6.5566
R1402 B.n300 B.n299 6.5566
R1403 B.n312 B.n134 6.5566
R1404 B.n573 B.n44 4.05904
R1405 B.n557 B.n556 4.05904
R1406 B.n299 B.n298 4.05904
R1407 B.n315 B.n134 4.05904
C0 B VP 2.22464f
C1 VN VTAIL 5.81515f
C2 B VDD2 2.03145f
C3 B VDD1 1.91381f
C4 w_n4474_n1944# VTAIL 2.20848f
C5 VP VTAIL 5.82933f
C6 VTAIL VDD2 7.15343f
C7 VDD1 VTAIL 7.1009f
C8 w_n4474_n1944# VN 9.43995f
C9 VP VN 7.0611f
C10 VN VDD2 4.64136f
C11 w_n4474_n1944# VP 10.0223f
C12 VDD1 VN 0.157568f
C13 w_n4474_n1944# VDD2 2.43393f
C14 w_n4474_n1944# VDD1 2.29121f
C15 VP VDD2 0.586556f
C16 B VTAIL 2.10992f
C17 VP VDD1 5.06699f
C18 VDD1 VDD2 2.16767f
C19 B VN 1.24534f
C20 B w_n4474_n1944# 8.54696f
C21 VDD2 VSUBS 2.056208f
C22 VDD1 VSUBS 1.75405f
C23 VTAIL VSUBS 0.644776f
C24 VN VSUBS 7.347991f
C25 VP VSUBS 3.664692f
C26 B VSUBS 4.470654f
C27 w_n4474_n1944# VSUBS 0.10904p
C28 B.n0 VSUBS 0.009864f
C29 B.n1 VSUBS 0.009864f
C30 B.n2 VSUBS 0.014589f
C31 B.n3 VSUBS 0.01118f
C32 B.n4 VSUBS 0.01118f
C33 B.n5 VSUBS 0.01118f
C34 B.n6 VSUBS 0.01118f
C35 B.n7 VSUBS 0.01118f
C36 B.n8 VSUBS 0.01118f
C37 B.n9 VSUBS 0.01118f
C38 B.n10 VSUBS 0.01118f
C39 B.n11 VSUBS 0.01118f
C40 B.n12 VSUBS 0.01118f
C41 B.n13 VSUBS 0.01118f
C42 B.n14 VSUBS 0.01118f
C43 B.n15 VSUBS 0.01118f
C44 B.n16 VSUBS 0.01118f
C45 B.n17 VSUBS 0.01118f
C46 B.n18 VSUBS 0.01118f
C47 B.n19 VSUBS 0.01118f
C48 B.n20 VSUBS 0.01118f
C49 B.n21 VSUBS 0.01118f
C50 B.n22 VSUBS 0.01118f
C51 B.n23 VSUBS 0.01118f
C52 B.n24 VSUBS 0.01118f
C53 B.n25 VSUBS 0.01118f
C54 B.n26 VSUBS 0.01118f
C55 B.n27 VSUBS 0.01118f
C56 B.n28 VSUBS 0.01118f
C57 B.n29 VSUBS 0.01118f
C58 B.n30 VSUBS 0.01118f
C59 B.n31 VSUBS 0.025834f
C60 B.n32 VSUBS 0.01118f
C61 B.n33 VSUBS 0.01118f
C62 B.n34 VSUBS 0.01118f
C63 B.n35 VSUBS 0.01118f
C64 B.n36 VSUBS 0.01118f
C65 B.n37 VSUBS 0.01118f
C66 B.n38 VSUBS 0.01118f
C67 B.n39 VSUBS 0.01118f
C68 B.n40 VSUBS 0.01118f
C69 B.n41 VSUBS 0.01118f
C70 B.t10 VSUBS 0.216403f
C71 B.t11 VSUBS 0.247611f
C72 B.t9 VSUBS 0.963384f
C73 B.n42 VSUBS 0.16211f
C74 B.n43 VSUBS 0.11163f
C75 B.n44 VSUBS 0.025902f
C76 B.n45 VSUBS 0.01118f
C77 B.n46 VSUBS 0.01118f
C78 B.n47 VSUBS 0.01118f
C79 B.n48 VSUBS 0.01118f
C80 B.n49 VSUBS 0.01118f
C81 B.t7 VSUBS 0.216403f
C82 B.t8 VSUBS 0.24761f
C83 B.t6 VSUBS 0.963384f
C84 B.n50 VSUBS 0.162111f
C85 B.n51 VSUBS 0.111631f
C86 B.n52 VSUBS 0.01118f
C87 B.n53 VSUBS 0.01118f
C88 B.n54 VSUBS 0.01118f
C89 B.n55 VSUBS 0.01118f
C90 B.n56 VSUBS 0.01118f
C91 B.n57 VSUBS 0.01118f
C92 B.n58 VSUBS 0.01118f
C93 B.n59 VSUBS 0.01118f
C94 B.n60 VSUBS 0.01118f
C95 B.n61 VSUBS 0.027433f
C96 B.n62 VSUBS 0.01118f
C97 B.n63 VSUBS 0.01118f
C98 B.n64 VSUBS 0.01118f
C99 B.n65 VSUBS 0.01118f
C100 B.n66 VSUBS 0.01118f
C101 B.n67 VSUBS 0.01118f
C102 B.n68 VSUBS 0.01118f
C103 B.n69 VSUBS 0.01118f
C104 B.n70 VSUBS 0.01118f
C105 B.n71 VSUBS 0.01118f
C106 B.n72 VSUBS 0.01118f
C107 B.n73 VSUBS 0.01118f
C108 B.n74 VSUBS 0.01118f
C109 B.n75 VSUBS 0.01118f
C110 B.n76 VSUBS 0.01118f
C111 B.n77 VSUBS 0.01118f
C112 B.n78 VSUBS 0.01118f
C113 B.n79 VSUBS 0.01118f
C114 B.n80 VSUBS 0.01118f
C115 B.n81 VSUBS 0.01118f
C116 B.n82 VSUBS 0.01118f
C117 B.n83 VSUBS 0.01118f
C118 B.n84 VSUBS 0.01118f
C119 B.n85 VSUBS 0.01118f
C120 B.n86 VSUBS 0.01118f
C121 B.n87 VSUBS 0.01118f
C122 B.n88 VSUBS 0.01118f
C123 B.n89 VSUBS 0.01118f
C124 B.n90 VSUBS 0.01118f
C125 B.n91 VSUBS 0.01118f
C126 B.n92 VSUBS 0.01118f
C127 B.n93 VSUBS 0.01118f
C128 B.n94 VSUBS 0.01118f
C129 B.n95 VSUBS 0.01118f
C130 B.n96 VSUBS 0.01118f
C131 B.n97 VSUBS 0.01118f
C132 B.n98 VSUBS 0.01118f
C133 B.n99 VSUBS 0.01118f
C134 B.n100 VSUBS 0.01118f
C135 B.n101 VSUBS 0.01118f
C136 B.n102 VSUBS 0.01118f
C137 B.n103 VSUBS 0.01118f
C138 B.n104 VSUBS 0.01118f
C139 B.n105 VSUBS 0.01118f
C140 B.n106 VSUBS 0.01118f
C141 B.n107 VSUBS 0.01118f
C142 B.n108 VSUBS 0.01118f
C143 B.n109 VSUBS 0.01118f
C144 B.n110 VSUBS 0.01118f
C145 B.n111 VSUBS 0.01118f
C146 B.n112 VSUBS 0.01118f
C147 B.n113 VSUBS 0.01118f
C148 B.n114 VSUBS 0.01118f
C149 B.n115 VSUBS 0.01118f
C150 B.n116 VSUBS 0.01118f
C151 B.n117 VSUBS 0.01118f
C152 B.n118 VSUBS 0.01118f
C153 B.n119 VSUBS 0.01118f
C154 B.n120 VSUBS 0.01118f
C155 B.n121 VSUBS 0.025834f
C156 B.n122 VSUBS 0.01118f
C157 B.n123 VSUBS 0.01118f
C158 B.n124 VSUBS 0.01118f
C159 B.n125 VSUBS 0.01118f
C160 B.n126 VSUBS 0.01118f
C161 B.n127 VSUBS 0.01118f
C162 B.n128 VSUBS 0.01118f
C163 B.n129 VSUBS 0.01118f
C164 B.n130 VSUBS 0.01118f
C165 B.n131 VSUBS 0.01118f
C166 B.t2 VSUBS 0.216403f
C167 B.t1 VSUBS 0.24761f
C168 B.t0 VSUBS 0.963384f
C169 B.n132 VSUBS 0.162111f
C170 B.n133 VSUBS 0.111631f
C171 B.n134 VSUBS 0.025902f
C172 B.n135 VSUBS 0.01118f
C173 B.n136 VSUBS 0.01118f
C174 B.n137 VSUBS 0.01118f
C175 B.n138 VSUBS 0.01118f
C176 B.n139 VSUBS 0.01118f
C177 B.t5 VSUBS 0.216403f
C178 B.t4 VSUBS 0.247611f
C179 B.t3 VSUBS 0.963384f
C180 B.n140 VSUBS 0.16211f
C181 B.n141 VSUBS 0.11163f
C182 B.n142 VSUBS 0.01118f
C183 B.n143 VSUBS 0.01118f
C184 B.n144 VSUBS 0.01118f
C185 B.n145 VSUBS 0.01118f
C186 B.n146 VSUBS 0.01118f
C187 B.n147 VSUBS 0.01118f
C188 B.n148 VSUBS 0.01118f
C189 B.n149 VSUBS 0.01118f
C190 B.n150 VSUBS 0.01118f
C191 B.n151 VSUBS 0.027433f
C192 B.n152 VSUBS 0.01118f
C193 B.n153 VSUBS 0.01118f
C194 B.n154 VSUBS 0.01118f
C195 B.n155 VSUBS 0.01118f
C196 B.n156 VSUBS 0.01118f
C197 B.n157 VSUBS 0.01118f
C198 B.n158 VSUBS 0.01118f
C199 B.n159 VSUBS 0.01118f
C200 B.n160 VSUBS 0.01118f
C201 B.n161 VSUBS 0.01118f
C202 B.n162 VSUBS 0.01118f
C203 B.n163 VSUBS 0.01118f
C204 B.n164 VSUBS 0.01118f
C205 B.n165 VSUBS 0.01118f
C206 B.n166 VSUBS 0.01118f
C207 B.n167 VSUBS 0.01118f
C208 B.n168 VSUBS 0.01118f
C209 B.n169 VSUBS 0.01118f
C210 B.n170 VSUBS 0.01118f
C211 B.n171 VSUBS 0.01118f
C212 B.n172 VSUBS 0.01118f
C213 B.n173 VSUBS 0.01118f
C214 B.n174 VSUBS 0.01118f
C215 B.n175 VSUBS 0.01118f
C216 B.n176 VSUBS 0.01118f
C217 B.n177 VSUBS 0.01118f
C218 B.n178 VSUBS 0.01118f
C219 B.n179 VSUBS 0.01118f
C220 B.n180 VSUBS 0.01118f
C221 B.n181 VSUBS 0.01118f
C222 B.n182 VSUBS 0.01118f
C223 B.n183 VSUBS 0.01118f
C224 B.n184 VSUBS 0.01118f
C225 B.n185 VSUBS 0.01118f
C226 B.n186 VSUBS 0.01118f
C227 B.n187 VSUBS 0.01118f
C228 B.n188 VSUBS 0.01118f
C229 B.n189 VSUBS 0.01118f
C230 B.n190 VSUBS 0.01118f
C231 B.n191 VSUBS 0.01118f
C232 B.n192 VSUBS 0.01118f
C233 B.n193 VSUBS 0.01118f
C234 B.n194 VSUBS 0.01118f
C235 B.n195 VSUBS 0.01118f
C236 B.n196 VSUBS 0.01118f
C237 B.n197 VSUBS 0.01118f
C238 B.n198 VSUBS 0.01118f
C239 B.n199 VSUBS 0.01118f
C240 B.n200 VSUBS 0.01118f
C241 B.n201 VSUBS 0.01118f
C242 B.n202 VSUBS 0.01118f
C243 B.n203 VSUBS 0.01118f
C244 B.n204 VSUBS 0.01118f
C245 B.n205 VSUBS 0.01118f
C246 B.n206 VSUBS 0.01118f
C247 B.n207 VSUBS 0.01118f
C248 B.n208 VSUBS 0.01118f
C249 B.n209 VSUBS 0.01118f
C250 B.n210 VSUBS 0.01118f
C251 B.n211 VSUBS 0.01118f
C252 B.n212 VSUBS 0.01118f
C253 B.n213 VSUBS 0.01118f
C254 B.n214 VSUBS 0.01118f
C255 B.n215 VSUBS 0.01118f
C256 B.n216 VSUBS 0.01118f
C257 B.n217 VSUBS 0.01118f
C258 B.n218 VSUBS 0.01118f
C259 B.n219 VSUBS 0.01118f
C260 B.n220 VSUBS 0.01118f
C261 B.n221 VSUBS 0.01118f
C262 B.n222 VSUBS 0.01118f
C263 B.n223 VSUBS 0.01118f
C264 B.n224 VSUBS 0.01118f
C265 B.n225 VSUBS 0.01118f
C266 B.n226 VSUBS 0.01118f
C267 B.n227 VSUBS 0.01118f
C268 B.n228 VSUBS 0.01118f
C269 B.n229 VSUBS 0.01118f
C270 B.n230 VSUBS 0.01118f
C271 B.n231 VSUBS 0.01118f
C272 B.n232 VSUBS 0.01118f
C273 B.n233 VSUBS 0.01118f
C274 B.n234 VSUBS 0.01118f
C275 B.n235 VSUBS 0.01118f
C276 B.n236 VSUBS 0.01118f
C277 B.n237 VSUBS 0.01118f
C278 B.n238 VSUBS 0.01118f
C279 B.n239 VSUBS 0.01118f
C280 B.n240 VSUBS 0.01118f
C281 B.n241 VSUBS 0.01118f
C282 B.n242 VSUBS 0.01118f
C283 B.n243 VSUBS 0.01118f
C284 B.n244 VSUBS 0.01118f
C285 B.n245 VSUBS 0.01118f
C286 B.n246 VSUBS 0.01118f
C287 B.n247 VSUBS 0.01118f
C288 B.n248 VSUBS 0.01118f
C289 B.n249 VSUBS 0.01118f
C290 B.n250 VSUBS 0.01118f
C291 B.n251 VSUBS 0.01118f
C292 B.n252 VSUBS 0.01118f
C293 B.n253 VSUBS 0.01118f
C294 B.n254 VSUBS 0.01118f
C295 B.n255 VSUBS 0.01118f
C296 B.n256 VSUBS 0.01118f
C297 B.n257 VSUBS 0.01118f
C298 B.n258 VSUBS 0.01118f
C299 B.n259 VSUBS 0.01118f
C300 B.n260 VSUBS 0.01118f
C301 B.n261 VSUBS 0.01118f
C302 B.n262 VSUBS 0.01118f
C303 B.n263 VSUBS 0.01118f
C304 B.n264 VSUBS 0.01118f
C305 B.n265 VSUBS 0.01118f
C306 B.n266 VSUBS 0.025834f
C307 B.n267 VSUBS 0.025834f
C308 B.n268 VSUBS 0.027433f
C309 B.n269 VSUBS 0.01118f
C310 B.n270 VSUBS 0.01118f
C311 B.n271 VSUBS 0.01118f
C312 B.n272 VSUBS 0.01118f
C313 B.n273 VSUBS 0.01118f
C314 B.n274 VSUBS 0.01118f
C315 B.n275 VSUBS 0.01118f
C316 B.n276 VSUBS 0.01118f
C317 B.n277 VSUBS 0.01118f
C318 B.n278 VSUBS 0.01118f
C319 B.n279 VSUBS 0.01118f
C320 B.n280 VSUBS 0.01118f
C321 B.n281 VSUBS 0.01118f
C322 B.n282 VSUBS 0.01118f
C323 B.n283 VSUBS 0.01118f
C324 B.n284 VSUBS 0.01118f
C325 B.n285 VSUBS 0.01118f
C326 B.n286 VSUBS 0.01118f
C327 B.n287 VSUBS 0.01118f
C328 B.n288 VSUBS 0.01118f
C329 B.n289 VSUBS 0.01118f
C330 B.n290 VSUBS 0.01118f
C331 B.n291 VSUBS 0.01118f
C332 B.n292 VSUBS 0.01118f
C333 B.n293 VSUBS 0.01118f
C334 B.n294 VSUBS 0.01118f
C335 B.n295 VSUBS 0.01118f
C336 B.n296 VSUBS 0.01118f
C337 B.n297 VSUBS 0.01118f
C338 B.n298 VSUBS 0.007727f
C339 B.n299 VSUBS 0.025902f
C340 B.n300 VSUBS 0.009042f
C341 B.n301 VSUBS 0.01118f
C342 B.n302 VSUBS 0.01118f
C343 B.n303 VSUBS 0.01118f
C344 B.n304 VSUBS 0.01118f
C345 B.n305 VSUBS 0.01118f
C346 B.n306 VSUBS 0.01118f
C347 B.n307 VSUBS 0.01118f
C348 B.n308 VSUBS 0.01118f
C349 B.n309 VSUBS 0.01118f
C350 B.n310 VSUBS 0.01118f
C351 B.n311 VSUBS 0.01118f
C352 B.n312 VSUBS 0.009042f
C353 B.n313 VSUBS 0.01118f
C354 B.n314 VSUBS 0.01118f
C355 B.n315 VSUBS 0.007727f
C356 B.n316 VSUBS 0.01118f
C357 B.n317 VSUBS 0.01118f
C358 B.n318 VSUBS 0.01118f
C359 B.n319 VSUBS 0.01118f
C360 B.n320 VSUBS 0.01118f
C361 B.n321 VSUBS 0.01118f
C362 B.n322 VSUBS 0.01118f
C363 B.n323 VSUBS 0.01118f
C364 B.n324 VSUBS 0.01118f
C365 B.n325 VSUBS 0.01118f
C366 B.n326 VSUBS 0.01118f
C367 B.n327 VSUBS 0.01118f
C368 B.n328 VSUBS 0.01118f
C369 B.n329 VSUBS 0.01118f
C370 B.n330 VSUBS 0.01118f
C371 B.n331 VSUBS 0.01118f
C372 B.n332 VSUBS 0.01118f
C373 B.n333 VSUBS 0.01118f
C374 B.n334 VSUBS 0.01118f
C375 B.n335 VSUBS 0.01118f
C376 B.n336 VSUBS 0.01118f
C377 B.n337 VSUBS 0.01118f
C378 B.n338 VSUBS 0.01118f
C379 B.n339 VSUBS 0.01118f
C380 B.n340 VSUBS 0.01118f
C381 B.n341 VSUBS 0.01118f
C382 B.n342 VSUBS 0.01118f
C383 B.n343 VSUBS 0.01118f
C384 B.n344 VSUBS 0.027433f
C385 B.n345 VSUBS 0.026148f
C386 B.n346 VSUBS 0.02712f
C387 B.n347 VSUBS 0.01118f
C388 B.n348 VSUBS 0.01118f
C389 B.n349 VSUBS 0.01118f
C390 B.n350 VSUBS 0.01118f
C391 B.n351 VSUBS 0.01118f
C392 B.n352 VSUBS 0.01118f
C393 B.n353 VSUBS 0.01118f
C394 B.n354 VSUBS 0.01118f
C395 B.n355 VSUBS 0.01118f
C396 B.n356 VSUBS 0.01118f
C397 B.n357 VSUBS 0.01118f
C398 B.n358 VSUBS 0.01118f
C399 B.n359 VSUBS 0.01118f
C400 B.n360 VSUBS 0.01118f
C401 B.n361 VSUBS 0.01118f
C402 B.n362 VSUBS 0.01118f
C403 B.n363 VSUBS 0.01118f
C404 B.n364 VSUBS 0.01118f
C405 B.n365 VSUBS 0.01118f
C406 B.n366 VSUBS 0.01118f
C407 B.n367 VSUBS 0.01118f
C408 B.n368 VSUBS 0.01118f
C409 B.n369 VSUBS 0.01118f
C410 B.n370 VSUBS 0.01118f
C411 B.n371 VSUBS 0.01118f
C412 B.n372 VSUBS 0.01118f
C413 B.n373 VSUBS 0.01118f
C414 B.n374 VSUBS 0.01118f
C415 B.n375 VSUBS 0.01118f
C416 B.n376 VSUBS 0.01118f
C417 B.n377 VSUBS 0.01118f
C418 B.n378 VSUBS 0.01118f
C419 B.n379 VSUBS 0.01118f
C420 B.n380 VSUBS 0.01118f
C421 B.n381 VSUBS 0.01118f
C422 B.n382 VSUBS 0.01118f
C423 B.n383 VSUBS 0.01118f
C424 B.n384 VSUBS 0.01118f
C425 B.n385 VSUBS 0.01118f
C426 B.n386 VSUBS 0.01118f
C427 B.n387 VSUBS 0.01118f
C428 B.n388 VSUBS 0.01118f
C429 B.n389 VSUBS 0.01118f
C430 B.n390 VSUBS 0.01118f
C431 B.n391 VSUBS 0.01118f
C432 B.n392 VSUBS 0.01118f
C433 B.n393 VSUBS 0.01118f
C434 B.n394 VSUBS 0.01118f
C435 B.n395 VSUBS 0.01118f
C436 B.n396 VSUBS 0.01118f
C437 B.n397 VSUBS 0.01118f
C438 B.n398 VSUBS 0.01118f
C439 B.n399 VSUBS 0.01118f
C440 B.n400 VSUBS 0.01118f
C441 B.n401 VSUBS 0.01118f
C442 B.n402 VSUBS 0.01118f
C443 B.n403 VSUBS 0.01118f
C444 B.n404 VSUBS 0.01118f
C445 B.n405 VSUBS 0.01118f
C446 B.n406 VSUBS 0.01118f
C447 B.n407 VSUBS 0.01118f
C448 B.n408 VSUBS 0.01118f
C449 B.n409 VSUBS 0.01118f
C450 B.n410 VSUBS 0.01118f
C451 B.n411 VSUBS 0.01118f
C452 B.n412 VSUBS 0.01118f
C453 B.n413 VSUBS 0.01118f
C454 B.n414 VSUBS 0.01118f
C455 B.n415 VSUBS 0.01118f
C456 B.n416 VSUBS 0.01118f
C457 B.n417 VSUBS 0.01118f
C458 B.n418 VSUBS 0.01118f
C459 B.n419 VSUBS 0.01118f
C460 B.n420 VSUBS 0.01118f
C461 B.n421 VSUBS 0.01118f
C462 B.n422 VSUBS 0.01118f
C463 B.n423 VSUBS 0.01118f
C464 B.n424 VSUBS 0.01118f
C465 B.n425 VSUBS 0.01118f
C466 B.n426 VSUBS 0.01118f
C467 B.n427 VSUBS 0.01118f
C468 B.n428 VSUBS 0.01118f
C469 B.n429 VSUBS 0.01118f
C470 B.n430 VSUBS 0.01118f
C471 B.n431 VSUBS 0.01118f
C472 B.n432 VSUBS 0.01118f
C473 B.n433 VSUBS 0.01118f
C474 B.n434 VSUBS 0.01118f
C475 B.n435 VSUBS 0.01118f
C476 B.n436 VSUBS 0.01118f
C477 B.n437 VSUBS 0.01118f
C478 B.n438 VSUBS 0.01118f
C479 B.n439 VSUBS 0.01118f
C480 B.n440 VSUBS 0.01118f
C481 B.n441 VSUBS 0.01118f
C482 B.n442 VSUBS 0.01118f
C483 B.n443 VSUBS 0.01118f
C484 B.n444 VSUBS 0.01118f
C485 B.n445 VSUBS 0.01118f
C486 B.n446 VSUBS 0.01118f
C487 B.n447 VSUBS 0.01118f
C488 B.n448 VSUBS 0.01118f
C489 B.n449 VSUBS 0.01118f
C490 B.n450 VSUBS 0.01118f
C491 B.n451 VSUBS 0.01118f
C492 B.n452 VSUBS 0.01118f
C493 B.n453 VSUBS 0.01118f
C494 B.n454 VSUBS 0.01118f
C495 B.n455 VSUBS 0.01118f
C496 B.n456 VSUBS 0.01118f
C497 B.n457 VSUBS 0.01118f
C498 B.n458 VSUBS 0.01118f
C499 B.n459 VSUBS 0.01118f
C500 B.n460 VSUBS 0.01118f
C501 B.n461 VSUBS 0.01118f
C502 B.n462 VSUBS 0.01118f
C503 B.n463 VSUBS 0.01118f
C504 B.n464 VSUBS 0.01118f
C505 B.n465 VSUBS 0.01118f
C506 B.n466 VSUBS 0.01118f
C507 B.n467 VSUBS 0.01118f
C508 B.n468 VSUBS 0.01118f
C509 B.n469 VSUBS 0.01118f
C510 B.n470 VSUBS 0.01118f
C511 B.n471 VSUBS 0.01118f
C512 B.n472 VSUBS 0.01118f
C513 B.n473 VSUBS 0.01118f
C514 B.n474 VSUBS 0.01118f
C515 B.n475 VSUBS 0.01118f
C516 B.n476 VSUBS 0.01118f
C517 B.n477 VSUBS 0.01118f
C518 B.n478 VSUBS 0.01118f
C519 B.n479 VSUBS 0.01118f
C520 B.n480 VSUBS 0.01118f
C521 B.n481 VSUBS 0.01118f
C522 B.n482 VSUBS 0.01118f
C523 B.n483 VSUBS 0.01118f
C524 B.n484 VSUBS 0.01118f
C525 B.n485 VSUBS 0.01118f
C526 B.n486 VSUBS 0.01118f
C527 B.n487 VSUBS 0.01118f
C528 B.n488 VSUBS 0.01118f
C529 B.n489 VSUBS 0.01118f
C530 B.n490 VSUBS 0.01118f
C531 B.n491 VSUBS 0.01118f
C532 B.n492 VSUBS 0.01118f
C533 B.n493 VSUBS 0.01118f
C534 B.n494 VSUBS 0.01118f
C535 B.n495 VSUBS 0.01118f
C536 B.n496 VSUBS 0.01118f
C537 B.n497 VSUBS 0.01118f
C538 B.n498 VSUBS 0.01118f
C539 B.n499 VSUBS 0.01118f
C540 B.n500 VSUBS 0.01118f
C541 B.n501 VSUBS 0.01118f
C542 B.n502 VSUBS 0.01118f
C543 B.n503 VSUBS 0.01118f
C544 B.n504 VSUBS 0.01118f
C545 B.n505 VSUBS 0.01118f
C546 B.n506 VSUBS 0.01118f
C547 B.n507 VSUBS 0.01118f
C548 B.n508 VSUBS 0.01118f
C549 B.n509 VSUBS 0.01118f
C550 B.n510 VSUBS 0.01118f
C551 B.n511 VSUBS 0.01118f
C552 B.n512 VSUBS 0.01118f
C553 B.n513 VSUBS 0.01118f
C554 B.n514 VSUBS 0.01118f
C555 B.n515 VSUBS 0.01118f
C556 B.n516 VSUBS 0.01118f
C557 B.n517 VSUBS 0.01118f
C558 B.n518 VSUBS 0.01118f
C559 B.n519 VSUBS 0.01118f
C560 B.n520 VSUBS 0.01118f
C561 B.n521 VSUBS 0.01118f
C562 B.n522 VSUBS 0.01118f
C563 B.n523 VSUBS 0.01118f
C564 B.n524 VSUBS 0.025834f
C565 B.n525 VSUBS 0.025834f
C566 B.n526 VSUBS 0.027433f
C567 B.n527 VSUBS 0.01118f
C568 B.n528 VSUBS 0.01118f
C569 B.n529 VSUBS 0.01118f
C570 B.n530 VSUBS 0.01118f
C571 B.n531 VSUBS 0.01118f
C572 B.n532 VSUBS 0.01118f
C573 B.n533 VSUBS 0.01118f
C574 B.n534 VSUBS 0.01118f
C575 B.n535 VSUBS 0.01118f
C576 B.n536 VSUBS 0.01118f
C577 B.n537 VSUBS 0.01118f
C578 B.n538 VSUBS 0.01118f
C579 B.n539 VSUBS 0.01118f
C580 B.n540 VSUBS 0.01118f
C581 B.n541 VSUBS 0.01118f
C582 B.n542 VSUBS 0.01118f
C583 B.n543 VSUBS 0.01118f
C584 B.n544 VSUBS 0.01118f
C585 B.n545 VSUBS 0.01118f
C586 B.n546 VSUBS 0.01118f
C587 B.n547 VSUBS 0.01118f
C588 B.n548 VSUBS 0.01118f
C589 B.n549 VSUBS 0.01118f
C590 B.n550 VSUBS 0.01118f
C591 B.n551 VSUBS 0.01118f
C592 B.n552 VSUBS 0.01118f
C593 B.n553 VSUBS 0.01118f
C594 B.n554 VSUBS 0.01118f
C595 B.n555 VSUBS 0.01118f
C596 B.n556 VSUBS 0.007727f
C597 B.n557 VSUBS 0.025902f
C598 B.n558 VSUBS 0.009042f
C599 B.n559 VSUBS 0.01118f
C600 B.n560 VSUBS 0.01118f
C601 B.n561 VSUBS 0.01118f
C602 B.n562 VSUBS 0.01118f
C603 B.n563 VSUBS 0.01118f
C604 B.n564 VSUBS 0.01118f
C605 B.n565 VSUBS 0.01118f
C606 B.n566 VSUBS 0.01118f
C607 B.n567 VSUBS 0.01118f
C608 B.n568 VSUBS 0.01118f
C609 B.n569 VSUBS 0.01118f
C610 B.n570 VSUBS 0.009042f
C611 B.n571 VSUBS 0.01118f
C612 B.n572 VSUBS 0.01118f
C613 B.n573 VSUBS 0.007727f
C614 B.n574 VSUBS 0.01118f
C615 B.n575 VSUBS 0.01118f
C616 B.n576 VSUBS 0.01118f
C617 B.n577 VSUBS 0.01118f
C618 B.n578 VSUBS 0.01118f
C619 B.n579 VSUBS 0.01118f
C620 B.n580 VSUBS 0.01118f
C621 B.n581 VSUBS 0.01118f
C622 B.n582 VSUBS 0.01118f
C623 B.n583 VSUBS 0.01118f
C624 B.n584 VSUBS 0.01118f
C625 B.n585 VSUBS 0.01118f
C626 B.n586 VSUBS 0.01118f
C627 B.n587 VSUBS 0.01118f
C628 B.n588 VSUBS 0.01118f
C629 B.n589 VSUBS 0.01118f
C630 B.n590 VSUBS 0.01118f
C631 B.n591 VSUBS 0.01118f
C632 B.n592 VSUBS 0.01118f
C633 B.n593 VSUBS 0.01118f
C634 B.n594 VSUBS 0.01118f
C635 B.n595 VSUBS 0.01118f
C636 B.n596 VSUBS 0.01118f
C637 B.n597 VSUBS 0.01118f
C638 B.n598 VSUBS 0.01118f
C639 B.n599 VSUBS 0.01118f
C640 B.n600 VSUBS 0.01118f
C641 B.n601 VSUBS 0.01118f
C642 B.n602 VSUBS 0.027433f
C643 B.n603 VSUBS 0.027433f
C644 B.n604 VSUBS 0.025834f
C645 B.n605 VSUBS 0.01118f
C646 B.n606 VSUBS 0.01118f
C647 B.n607 VSUBS 0.01118f
C648 B.n608 VSUBS 0.01118f
C649 B.n609 VSUBS 0.01118f
C650 B.n610 VSUBS 0.01118f
C651 B.n611 VSUBS 0.01118f
C652 B.n612 VSUBS 0.01118f
C653 B.n613 VSUBS 0.01118f
C654 B.n614 VSUBS 0.01118f
C655 B.n615 VSUBS 0.01118f
C656 B.n616 VSUBS 0.01118f
C657 B.n617 VSUBS 0.01118f
C658 B.n618 VSUBS 0.01118f
C659 B.n619 VSUBS 0.01118f
C660 B.n620 VSUBS 0.01118f
C661 B.n621 VSUBS 0.01118f
C662 B.n622 VSUBS 0.01118f
C663 B.n623 VSUBS 0.01118f
C664 B.n624 VSUBS 0.01118f
C665 B.n625 VSUBS 0.01118f
C666 B.n626 VSUBS 0.01118f
C667 B.n627 VSUBS 0.01118f
C668 B.n628 VSUBS 0.01118f
C669 B.n629 VSUBS 0.01118f
C670 B.n630 VSUBS 0.01118f
C671 B.n631 VSUBS 0.01118f
C672 B.n632 VSUBS 0.01118f
C673 B.n633 VSUBS 0.01118f
C674 B.n634 VSUBS 0.01118f
C675 B.n635 VSUBS 0.01118f
C676 B.n636 VSUBS 0.01118f
C677 B.n637 VSUBS 0.01118f
C678 B.n638 VSUBS 0.01118f
C679 B.n639 VSUBS 0.01118f
C680 B.n640 VSUBS 0.01118f
C681 B.n641 VSUBS 0.01118f
C682 B.n642 VSUBS 0.01118f
C683 B.n643 VSUBS 0.01118f
C684 B.n644 VSUBS 0.01118f
C685 B.n645 VSUBS 0.01118f
C686 B.n646 VSUBS 0.01118f
C687 B.n647 VSUBS 0.01118f
C688 B.n648 VSUBS 0.01118f
C689 B.n649 VSUBS 0.01118f
C690 B.n650 VSUBS 0.01118f
C691 B.n651 VSUBS 0.01118f
C692 B.n652 VSUBS 0.01118f
C693 B.n653 VSUBS 0.01118f
C694 B.n654 VSUBS 0.01118f
C695 B.n655 VSUBS 0.01118f
C696 B.n656 VSUBS 0.01118f
C697 B.n657 VSUBS 0.01118f
C698 B.n658 VSUBS 0.01118f
C699 B.n659 VSUBS 0.01118f
C700 B.n660 VSUBS 0.01118f
C701 B.n661 VSUBS 0.01118f
C702 B.n662 VSUBS 0.01118f
C703 B.n663 VSUBS 0.01118f
C704 B.n664 VSUBS 0.01118f
C705 B.n665 VSUBS 0.01118f
C706 B.n666 VSUBS 0.01118f
C707 B.n667 VSUBS 0.01118f
C708 B.n668 VSUBS 0.01118f
C709 B.n669 VSUBS 0.01118f
C710 B.n670 VSUBS 0.01118f
C711 B.n671 VSUBS 0.01118f
C712 B.n672 VSUBS 0.01118f
C713 B.n673 VSUBS 0.01118f
C714 B.n674 VSUBS 0.01118f
C715 B.n675 VSUBS 0.01118f
C716 B.n676 VSUBS 0.01118f
C717 B.n677 VSUBS 0.01118f
C718 B.n678 VSUBS 0.01118f
C719 B.n679 VSUBS 0.01118f
C720 B.n680 VSUBS 0.01118f
C721 B.n681 VSUBS 0.01118f
C722 B.n682 VSUBS 0.01118f
C723 B.n683 VSUBS 0.01118f
C724 B.n684 VSUBS 0.01118f
C725 B.n685 VSUBS 0.01118f
C726 B.n686 VSUBS 0.01118f
C727 B.n687 VSUBS 0.01118f
C728 B.n688 VSUBS 0.01118f
C729 B.n689 VSUBS 0.01118f
C730 B.n690 VSUBS 0.01118f
C731 B.n691 VSUBS 0.014589f
C732 B.n692 VSUBS 0.015541f
C733 B.n693 VSUBS 0.030904f
C734 VDD2.t7 VSUBS 1.17165f
C735 VDD2.t1 VSUBS 0.13607f
C736 VDD2.t4 VSUBS 0.13607f
C737 VDD2.n0 VSUBS 0.847422f
C738 VDD2.n1 VSUBS 1.77434f
C739 VDD2.t0 VSUBS 0.13607f
C740 VDD2.t8 VSUBS 0.13607f
C741 VDD2.n2 VSUBS 0.866314f
C742 VDD2.n3 VSUBS 3.73386f
C743 VDD2.t3 VSUBS 1.15071f
C744 VDD2.n4 VSUBS 3.83912f
C745 VDD2.t5 VSUBS 0.13607f
C746 VDD2.t9 VSUBS 0.13607f
C747 VDD2.n5 VSUBS 0.847426f
C748 VDD2.n6 VSUBS 0.901447f
C749 VDD2.t2 VSUBS 0.13607f
C750 VDD2.t6 VSUBS 0.13607f
C751 VDD2.n7 VSUBS 0.86627f
C752 VN.n0 VSUBS 0.050359f
C753 VN.t1 VSUBS 1.26063f
C754 VN.n1 VSUBS 0.067453f
C755 VN.n2 VSUBS 0.038199f
C756 VN.t9 VSUBS 1.26063f
C757 VN.n3 VSUBS 0.485986f
C758 VN.n4 VSUBS 0.038199f
C759 VN.n5 VSUBS 0.051301f
C760 VN.n6 VSUBS 0.038199f
C761 VN.t5 VSUBS 1.26063f
C762 VN.n7 VSUBS 0.070837f
C763 VN.n8 VSUBS 0.038199f
C764 VN.n9 VSUBS 0.047756f
C765 VN.t2 VSUBS 1.55633f
C766 VN.t8 VSUBS 1.26063f
C767 VN.n10 VSUBS 0.59023f
C768 VN.n11 VSUBS 0.576134f
C769 VN.n12 VSUBS 0.368153f
C770 VN.n13 VSUBS 0.038199f
C771 VN.n14 VSUBS 0.070837f
C772 VN.n15 VSUBS 0.059756f
C773 VN.n16 VSUBS 0.051301f
C774 VN.n17 VSUBS 0.038199f
C775 VN.n18 VSUBS 0.038199f
C776 VN.n19 VSUBS 0.038199f
C777 VN.n20 VSUBS 0.053352f
C778 VN.n21 VSUBS 0.485986f
C779 VN.n22 VSUBS 0.053352f
C780 VN.n23 VSUBS 0.070837f
C781 VN.n24 VSUBS 0.038199f
C782 VN.n25 VSUBS 0.038199f
C783 VN.n26 VSUBS 0.038199f
C784 VN.n27 VSUBS 0.059756f
C785 VN.n28 VSUBS 0.070837f
C786 VN.n29 VSUBS 0.047756f
C787 VN.n30 VSUBS 0.038199f
C788 VN.n31 VSUBS 0.038199f
C789 VN.n32 VSUBS 0.058947f
C790 VN.n33 VSUBS 0.074481f
C791 VN.n34 VSUBS 0.039959f
C792 VN.n35 VSUBS 0.038199f
C793 VN.n36 VSUBS 0.038199f
C794 VN.n37 VSUBS 0.038199f
C795 VN.n38 VSUBS 0.070837f
C796 VN.n39 VSUBS 0.042161f
C797 VN.n40 VSUBS 0.601413f
C798 VN.n41 VSUBS 0.066868f
C799 VN.n42 VSUBS 0.050359f
C800 VN.t6 VSUBS 1.26063f
C801 VN.n43 VSUBS 0.067453f
C802 VN.n44 VSUBS 0.038199f
C803 VN.t4 VSUBS 1.26063f
C804 VN.n45 VSUBS 0.485986f
C805 VN.n46 VSUBS 0.038199f
C806 VN.n47 VSUBS 0.051301f
C807 VN.n48 VSUBS 0.038199f
C808 VN.t0 VSUBS 1.26063f
C809 VN.n49 VSUBS 0.070837f
C810 VN.n50 VSUBS 0.038199f
C811 VN.n51 VSUBS 0.047756f
C812 VN.t3 VSUBS 1.55633f
C813 VN.t7 VSUBS 1.26063f
C814 VN.n52 VSUBS 0.59023f
C815 VN.n53 VSUBS 0.576134f
C816 VN.n54 VSUBS 0.368153f
C817 VN.n55 VSUBS 0.038199f
C818 VN.n56 VSUBS 0.070837f
C819 VN.n57 VSUBS 0.059756f
C820 VN.n58 VSUBS 0.051301f
C821 VN.n59 VSUBS 0.038199f
C822 VN.n60 VSUBS 0.038199f
C823 VN.n61 VSUBS 0.038199f
C824 VN.n62 VSUBS 0.053352f
C825 VN.n63 VSUBS 0.485986f
C826 VN.n64 VSUBS 0.053352f
C827 VN.n65 VSUBS 0.070837f
C828 VN.n66 VSUBS 0.038199f
C829 VN.n67 VSUBS 0.038199f
C830 VN.n68 VSUBS 0.038199f
C831 VN.n69 VSUBS 0.059756f
C832 VN.n70 VSUBS 0.070837f
C833 VN.n71 VSUBS 0.047756f
C834 VN.n72 VSUBS 0.038199f
C835 VN.n73 VSUBS 0.038199f
C836 VN.n74 VSUBS 0.058947f
C837 VN.n75 VSUBS 0.074481f
C838 VN.n76 VSUBS 0.039959f
C839 VN.n77 VSUBS 0.038199f
C840 VN.n78 VSUBS 0.038199f
C841 VN.n79 VSUBS 0.038199f
C842 VN.n80 VSUBS 0.070837f
C843 VN.n81 VSUBS 0.042161f
C844 VN.n82 VSUBS 0.601413f
C845 VN.n83 VSUBS 1.99959f
C846 VDD1.t0 VSUBS 1.05592f
C847 VDD1.t5 VSUBS 0.12263f
C848 VDD1.t3 VSUBS 0.12263f
C849 VDD1.n0 VSUBS 0.763722f
C850 VDD1.n1 VSUBS 1.60942f
C851 VDD1.t6 VSUBS 1.05592f
C852 VDD1.t4 VSUBS 0.12263f
C853 VDD1.t7 VSUBS 0.12263f
C854 VDD1.n2 VSUBS 0.763718f
C855 VDD1.n3 VSUBS 1.59908f
C856 VDD1.t1 VSUBS 0.12263f
C857 VDD1.t8 VSUBS 0.12263f
C858 VDD1.n4 VSUBS 0.780744f
C859 VDD1.n5 VSUBS 3.51619f
C860 VDD1.t2 VSUBS 0.12263f
C861 VDD1.t9 VSUBS 0.12263f
C862 VDD1.n6 VSUBS 0.763718f
C863 VDD1.n7 VSUBS 3.5526f
C864 VTAIL.t18 VSUBS 0.134234f
C865 VTAIL.t3 VSUBS 0.134234f
C866 VTAIL.n0 VSUBS 0.730832f
C867 VTAIL.n1 VSUBS 0.999832f
C868 VTAIL.t9 VSUBS 1.0254f
C869 VTAIL.n2 VSUBS 1.13542f
C870 VTAIL.t16 VSUBS 0.134234f
C871 VTAIL.t15 VSUBS 0.134234f
C872 VTAIL.n3 VSUBS 0.730832f
C873 VTAIL.n4 VSUBS 1.15236f
C874 VTAIL.t7 VSUBS 0.134234f
C875 VTAIL.t12 VSUBS 0.134234f
C876 VTAIL.n5 VSUBS 0.730832f
C877 VTAIL.n6 VSUBS 2.37939f
C878 VTAIL.t0 VSUBS 0.134234f
C879 VTAIL.t17 VSUBS 0.134234f
C880 VTAIL.n7 VSUBS 0.730837f
C881 VTAIL.n8 VSUBS 2.37939f
C882 VTAIL.t5 VSUBS 0.134234f
C883 VTAIL.t19 VSUBS 0.134234f
C884 VTAIL.n9 VSUBS 0.730837f
C885 VTAIL.n10 VSUBS 1.15236f
C886 VTAIL.t4 VSUBS 1.0254f
C887 VTAIL.n11 VSUBS 1.13541f
C888 VTAIL.t8 VSUBS 0.134234f
C889 VTAIL.t14 VSUBS 0.134234f
C890 VTAIL.n12 VSUBS 0.730837f
C891 VTAIL.n13 VSUBS 1.06389f
C892 VTAIL.t10 VSUBS 0.134234f
C893 VTAIL.t13 VSUBS 0.134234f
C894 VTAIL.n14 VSUBS 0.730837f
C895 VTAIL.n15 VSUBS 1.15236f
C896 VTAIL.t11 VSUBS 1.0254f
C897 VTAIL.n16 VSUBS 2.16858f
C898 VTAIL.t1 VSUBS 1.0254f
C899 VTAIL.n17 VSUBS 2.16858f
C900 VTAIL.t6 VSUBS 0.134234f
C901 VTAIL.t2 VSUBS 0.134234f
C902 VTAIL.n18 VSUBS 0.730832f
C903 VTAIL.n19 VSUBS 0.934082f
C904 VP.n0 VSUBS 0.05665f
C905 VP.t1 VSUBS 1.41811f
C906 VP.n1 VSUBS 0.07588f
C907 VP.n2 VSUBS 0.042971f
C908 VP.t8 VSUBS 1.41811f
C909 VP.n3 VSUBS 0.546696f
C910 VP.n4 VSUBS 0.042971f
C911 VP.n5 VSUBS 0.057709f
C912 VP.n6 VSUBS 0.042971f
C913 VP.t2 VSUBS 1.41811f
C914 VP.n7 VSUBS 0.079686f
C915 VP.n8 VSUBS 0.042971f
C916 VP.n9 VSUBS 0.053722f
C917 VP.n10 VSUBS 0.042971f
C918 VP.n11 VSUBS 0.07588f
C919 VP.n12 VSUBS 0.05665f
C920 VP.t3 VSUBS 1.41811f
C921 VP.n13 VSUBS 0.05665f
C922 VP.t0 VSUBS 1.41811f
C923 VP.n14 VSUBS 0.07588f
C924 VP.n15 VSUBS 0.042971f
C925 VP.t7 VSUBS 1.41811f
C926 VP.n16 VSUBS 0.546696f
C927 VP.n17 VSUBS 0.042971f
C928 VP.n18 VSUBS 0.057709f
C929 VP.n19 VSUBS 0.042971f
C930 VP.t6 VSUBS 1.41811f
C931 VP.n20 VSUBS 0.079686f
C932 VP.n21 VSUBS 0.042971f
C933 VP.n22 VSUBS 0.053722f
C934 VP.t9 VSUBS 1.75075f
C935 VP.t4 VSUBS 1.41811f
C936 VP.n23 VSUBS 0.663963f
C937 VP.n24 VSUBS 0.648105f
C938 VP.n25 VSUBS 0.414144f
C939 VP.n26 VSUBS 0.042971f
C940 VP.n27 VSUBS 0.079686f
C941 VP.n28 VSUBS 0.06722f
C942 VP.n29 VSUBS 0.057709f
C943 VP.n30 VSUBS 0.042971f
C944 VP.n31 VSUBS 0.042971f
C945 VP.n32 VSUBS 0.042971f
C946 VP.n33 VSUBS 0.060016f
C947 VP.n34 VSUBS 0.546696f
C948 VP.n35 VSUBS 0.060016f
C949 VP.n36 VSUBS 0.079686f
C950 VP.n37 VSUBS 0.042971f
C951 VP.n38 VSUBS 0.042971f
C952 VP.n39 VSUBS 0.042971f
C953 VP.n40 VSUBS 0.06722f
C954 VP.n41 VSUBS 0.079686f
C955 VP.n42 VSUBS 0.053722f
C956 VP.n43 VSUBS 0.042971f
C957 VP.n44 VSUBS 0.042971f
C958 VP.n45 VSUBS 0.066311f
C959 VP.n46 VSUBS 0.083785f
C960 VP.n47 VSUBS 0.044951f
C961 VP.n48 VSUBS 0.042971f
C962 VP.n49 VSUBS 0.042971f
C963 VP.n50 VSUBS 0.042971f
C964 VP.n51 VSUBS 0.079686f
C965 VP.n52 VSUBS 0.047428f
C966 VP.n53 VSUBS 0.676543f
C967 VP.n54 VSUBS 2.22611f
C968 VP.n55 VSUBS 2.25865f
C969 VP.n56 VSUBS 0.676543f
C970 VP.n57 VSUBS 0.047428f
C971 VP.n58 VSUBS 0.079686f
C972 VP.n59 VSUBS 0.042971f
C973 VP.n60 VSUBS 0.042971f
C974 VP.n61 VSUBS 0.042971f
C975 VP.n62 VSUBS 0.044951f
C976 VP.n63 VSUBS 0.083785f
C977 VP.t5 VSUBS 1.41811f
C978 VP.n64 VSUBS 0.546696f
C979 VP.n65 VSUBS 0.066311f
C980 VP.n66 VSUBS 0.042971f
C981 VP.n67 VSUBS 0.042971f
C982 VP.n68 VSUBS 0.042971f
C983 VP.n69 VSUBS 0.079686f
C984 VP.n70 VSUBS 0.06722f
C985 VP.n71 VSUBS 0.057709f
C986 VP.n72 VSUBS 0.042971f
C987 VP.n73 VSUBS 0.042971f
C988 VP.n74 VSUBS 0.042971f
C989 VP.n75 VSUBS 0.060016f
C990 VP.n76 VSUBS 0.546696f
C991 VP.n77 VSUBS 0.060016f
C992 VP.n78 VSUBS 0.079686f
C993 VP.n79 VSUBS 0.042971f
C994 VP.n80 VSUBS 0.042971f
C995 VP.n81 VSUBS 0.042971f
C996 VP.n82 VSUBS 0.06722f
C997 VP.n83 VSUBS 0.079686f
C998 VP.n84 VSUBS 0.053722f
C999 VP.n85 VSUBS 0.042971f
C1000 VP.n86 VSUBS 0.042971f
C1001 VP.n87 VSUBS 0.066311f
C1002 VP.n88 VSUBS 0.083785f
C1003 VP.n89 VSUBS 0.044951f
C1004 VP.n90 VSUBS 0.042971f
C1005 VP.n91 VSUBS 0.042971f
C1006 VP.n92 VSUBS 0.042971f
C1007 VP.n93 VSUBS 0.079686f
C1008 VP.n94 VSUBS 0.047428f
C1009 VP.n95 VSUBS 0.676543f
C1010 VP.n96 VSUBS 0.075221f
.ends

