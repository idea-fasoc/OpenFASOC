* NGSPICE file created from diff_pair_sample_0608.ext - technology: sky130A

.subckt diff_pair_sample_0608 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t9 B.t0 sky130_fd_pr__nfet_01v8 ad=4.3953 pd=23.32 as=1.85955 ps=11.6 w=11.27 l=2.5
X1 VDD2.t9 VN.t0 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=1.85955 pd=11.6 as=1.85955 ps=11.6 w=11.27 l=2.5
X2 VDD2.t8 VN.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=4.3953 pd=23.32 as=1.85955 ps=11.6 w=11.27 l=2.5
X3 VDD1.t8 VP.t1 VTAIL.t15 B.t9 sky130_fd_pr__nfet_01v8 ad=1.85955 pd=11.6 as=1.85955 ps=11.6 w=11.27 l=2.5
X4 VTAIL.t11 VP.t2 VDD1.t7 B.t1 sky130_fd_pr__nfet_01v8 ad=1.85955 pd=11.6 as=1.85955 ps=11.6 w=11.27 l=2.5
X5 VTAIL.t10 VP.t3 VDD1.t6 B.t4 sky130_fd_pr__nfet_01v8 ad=1.85955 pd=11.6 as=1.85955 ps=11.6 w=11.27 l=2.5
X6 VTAIL.t4 VN.t2 VDD2.t7 B.t4 sky130_fd_pr__nfet_01v8 ad=1.85955 pd=11.6 as=1.85955 ps=11.6 w=11.27 l=2.5
X7 VTAIL.t13 VP.t4 VDD1.t5 B.t8 sky130_fd_pr__nfet_01v8 ad=1.85955 pd=11.6 as=1.85955 ps=11.6 w=11.27 l=2.5
X8 VDD2.t6 VN.t3 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=4.3953 pd=23.32 as=1.85955 ps=11.6 w=11.27 l=2.5
X9 VTAIL.t17 VN.t4 VDD2.t5 B.t8 sky130_fd_pr__nfet_01v8 ad=1.85955 pd=11.6 as=1.85955 ps=11.6 w=11.27 l=2.5
X10 VDD1.t4 VP.t5 VTAIL.t16 B.t6 sky130_fd_pr__nfet_01v8 ad=1.85955 pd=11.6 as=4.3953 ps=23.32 w=11.27 l=2.5
X11 VDD1.t3 VP.t6 VTAIL.t14 B.t7 sky130_fd_pr__nfet_01v8 ad=1.85955 pd=11.6 as=4.3953 ps=23.32 w=11.27 l=2.5
X12 B.t23 B.t21 B.t22 B.t18 sky130_fd_pr__nfet_01v8 ad=4.3953 pd=23.32 as=0 ps=0 w=11.27 l=2.5
X13 B.t20 B.t17 B.t19 B.t18 sky130_fd_pr__nfet_01v8 ad=4.3953 pd=23.32 as=0 ps=0 w=11.27 l=2.5
X14 VDD2.t4 VN.t5 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=1.85955 pd=11.6 as=4.3953 ps=23.32 w=11.27 l=2.5
X15 VDD2.t3 VN.t6 VTAIL.t18 B.t7 sky130_fd_pr__nfet_01v8 ad=1.85955 pd=11.6 as=4.3953 ps=23.32 w=11.27 l=2.5
X16 VDD1.t2 VP.t7 VTAIL.t8 B.t3 sky130_fd_pr__nfet_01v8 ad=4.3953 pd=23.32 as=1.85955 ps=11.6 w=11.27 l=2.5
X17 VTAIL.t1 VN.t7 VDD2.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=1.85955 pd=11.6 as=1.85955 ps=11.6 w=11.27 l=2.5
X18 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=4.3953 pd=23.32 as=0 ps=0 w=11.27 l=2.5
X19 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=4.3953 pd=23.32 as=0 ps=0 w=11.27 l=2.5
X20 VDD2.t1 VN.t8 VTAIL.t19 B.t9 sky130_fd_pr__nfet_01v8 ad=1.85955 pd=11.6 as=1.85955 ps=11.6 w=11.27 l=2.5
X21 VDD1.t1 VP.t8 VTAIL.t7 B.t5 sky130_fd_pr__nfet_01v8 ad=1.85955 pd=11.6 as=1.85955 ps=11.6 w=11.27 l=2.5
X22 VTAIL.t2 VN.t9 VDD2.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=1.85955 pd=11.6 as=1.85955 ps=11.6 w=11.27 l=2.5
X23 VTAIL.t12 VP.t9 VDD1.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=1.85955 pd=11.6 as=1.85955 ps=11.6 w=11.27 l=2.5
R0 VP.n25 VP.n24 161.3
R1 VP.n26 VP.n21 161.3
R2 VP.n28 VP.n27 161.3
R3 VP.n29 VP.n20 161.3
R4 VP.n31 VP.n30 161.3
R5 VP.n32 VP.n19 161.3
R6 VP.n34 VP.n33 161.3
R7 VP.n35 VP.n18 161.3
R8 VP.n37 VP.n36 161.3
R9 VP.n38 VP.n17 161.3
R10 VP.n40 VP.n39 161.3
R11 VP.n42 VP.n41 161.3
R12 VP.n43 VP.n15 161.3
R13 VP.n45 VP.n44 161.3
R14 VP.n46 VP.n14 161.3
R15 VP.n48 VP.n47 161.3
R16 VP.n49 VP.n13 161.3
R17 VP.n88 VP.n0 161.3
R18 VP.n87 VP.n86 161.3
R19 VP.n85 VP.n1 161.3
R20 VP.n84 VP.n83 161.3
R21 VP.n82 VP.n2 161.3
R22 VP.n81 VP.n80 161.3
R23 VP.n79 VP.n78 161.3
R24 VP.n77 VP.n4 161.3
R25 VP.n76 VP.n75 161.3
R26 VP.n74 VP.n5 161.3
R27 VP.n73 VP.n72 161.3
R28 VP.n71 VP.n6 161.3
R29 VP.n70 VP.n69 161.3
R30 VP.n68 VP.n7 161.3
R31 VP.n67 VP.n66 161.3
R32 VP.n65 VP.n8 161.3
R33 VP.n64 VP.n63 161.3
R34 VP.n62 VP.n61 161.3
R35 VP.n60 VP.n10 161.3
R36 VP.n59 VP.n58 161.3
R37 VP.n57 VP.n11 161.3
R38 VP.n56 VP.n55 161.3
R39 VP.n54 VP.n12 161.3
R40 VP.n23 VP.t0 141.612
R41 VP.n71 VP.t8 108.644
R42 VP.n53 VP.t7 108.644
R43 VP.n9 VP.t3 108.644
R44 VP.n3 VP.t9 108.644
R45 VP.n89 VP.t5 108.644
R46 VP.n32 VP.t1 108.644
R47 VP.n50 VP.t6 108.644
R48 VP.n16 VP.t4 108.644
R49 VP.n22 VP.t2 108.644
R50 VP.n53 VP.n52 102.927
R51 VP.n90 VP.n89 102.927
R52 VP.n51 VP.n50 102.927
R53 VP.n59 VP.n11 56.5193
R54 VP.n83 VP.n1 56.5193
R55 VP.n44 VP.n14 56.5193
R56 VP.n23 VP.n22 56.1683
R57 VP.n52 VP.n51 51.9806
R58 VP.n66 VP.n7 48.7492
R59 VP.n76 VP.n5 48.7492
R60 VP.n37 VP.n18 48.7492
R61 VP.n27 VP.n20 48.7492
R62 VP.n66 VP.n65 32.2376
R63 VP.n77 VP.n76 32.2376
R64 VP.n38 VP.n37 32.2376
R65 VP.n27 VP.n26 32.2376
R66 VP.n55 VP.n54 24.4675
R67 VP.n55 VP.n11 24.4675
R68 VP.n60 VP.n59 24.4675
R69 VP.n61 VP.n60 24.4675
R70 VP.n65 VP.n64 24.4675
R71 VP.n70 VP.n7 24.4675
R72 VP.n71 VP.n70 24.4675
R73 VP.n72 VP.n71 24.4675
R74 VP.n72 VP.n5 24.4675
R75 VP.n78 VP.n77 24.4675
R76 VP.n82 VP.n81 24.4675
R77 VP.n83 VP.n82 24.4675
R78 VP.n87 VP.n1 24.4675
R79 VP.n88 VP.n87 24.4675
R80 VP.n48 VP.n14 24.4675
R81 VP.n49 VP.n48 24.4675
R82 VP.n39 VP.n38 24.4675
R83 VP.n43 VP.n42 24.4675
R84 VP.n44 VP.n43 24.4675
R85 VP.n31 VP.n20 24.4675
R86 VP.n32 VP.n31 24.4675
R87 VP.n33 VP.n32 24.4675
R88 VP.n33 VP.n18 24.4675
R89 VP.n26 VP.n25 24.4675
R90 VP.n64 VP.n9 16.1487
R91 VP.n78 VP.n3 16.1487
R92 VP.n39 VP.n16 16.1487
R93 VP.n25 VP.n22 16.1487
R94 VP.n61 VP.n9 8.31928
R95 VP.n81 VP.n3 8.31928
R96 VP.n42 VP.n16 8.31928
R97 VP.n54 VP.n53 7.82994
R98 VP.n89 VP.n88 7.82994
R99 VP.n50 VP.n49 7.82994
R100 VP.n24 VP.n23 6.98649
R101 VP.n51 VP.n13 0.278367
R102 VP.n52 VP.n12 0.278367
R103 VP.n90 VP.n0 0.278367
R104 VP.n24 VP.n21 0.189894
R105 VP.n28 VP.n21 0.189894
R106 VP.n29 VP.n28 0.189894
R107 VP.n30 VP.n29 0.189894
R108 VP.n30 VP.n19 0.189894
R109 VP.n34 VP.n19 0.189894
R110 VP.n35 VP.n34 0.189894
R111 VP.n36 VP.n35 0.189894
R112 VP.n36 VP.n17 0.189894
R113 VP.n40 VP.n17 0.189894
R114 VP.n41 VP.n40 0.189894
R115 VP.n41 VP.n15 0.189894
R116 VP.n45 VP.n15 0.189894
R117 VP.n46 VP.n45 0.189894
R118 VP.n47 VP.n46 0.189894
R119 VP.n47 VP.n13 0.189894
R120 VP.n56 VP.n12 0.189894
R121 VP.n57 VP.n56 0.189894
R122 VP.n58 VP.n57 0.189894
R123 VP.n58 VP.n10 0.189894
R124 VP.n62 VP.n10 0.189894
R125 VP.n63 VP.n62 0.189894
R126 VP.n63 VP.n8 0.189894
R127 VP.n67 VP.n8 0.189894
R128 VP.n68 VP.n67 0.189894
R129 VP.n69 VP.n68 0.189894
R130 VP.n69 VP.n6 0.189894
R131 VP.n73 VP.n6 0.189894
R132 VP.n74 VP.n73 0.189894
R133 VP.n75 VP.n74 0.189894
R134 VP.n75 VP.n4 0.189894
R135 VP.n79 VP.n4 0.189894
R136 VP.n80 VP.n79 0.189894
R137 VP.n80 VP.n2 0.189894
R138 VP.n84 VP.n2 0.189894
R139 VP.n85 VP.n84 0.189894
R140 VP.n86 VP.n85 0.189894
R141 VP.n86 VP.n0 0.189894
R142 VP VP.n90 0.153454
R143 VTAIL.n260 VTAIL.n259 289.615
R144 VTAIL.n62 VTAIL.n61 289.615
R145 VTAIL.n198 VTAIL.n197 289.615
R146 VTAIL.n132 VTAIL.n131 289.615
R147 VTAIL.n221 VTAIL.n220 185
R148 VTAIL.n218 VTAIL.n217 185
R149 VTAIL.n227 VTAIL.n226 185
R150 VTAIL.n229 VTAIL.n228 185
R151 VTAIL.n214 VTAIL.n213 185
R152 VTAIL.n235 VTAIL.n234 185
R153 VTAIL.n237 VTAIL.n236 185
R154 VTAIL.n210 VTAIL.n209 185
R155 VTAIL.n243 VTAIL.n242 185
R156 VTAIL.n245 VTAIL.n244 185
R157 VTAIL.n206 VTAIL.n205 185
R158 VTAIL.n251 VTAIL.n250 185
R159 VTAIL.n253 VTAIL.n252 185
R160 VTAIL.n202 VTAIL.n201 185
R161 VTAIL.n259 VTAIL.n258 185
R162 VTAIL.n23 VTAIL.n22 185
R163 VTAIL.n20 VTAIL.n19 185
R164 VTAIL.n29 VTAIL.n28 185
R165 VTAIL.n31 VTAIL.n30 185
R166 VTAIL.n16 VTAIL.n15 185
R167 VTAIL.n37 VTAIL.n36 185
R168 VTAIL.n39 VTAIL.n38 185
R169 VTAIL.n12 VTAIL.n11 185
R170 VTAIL.n45 VTAIL.n44 185
R171 VTAIL.n47 VTAIL.n46 185
R172 VTAIL.n8 VTAIL.n7 185
R173 VTAIL.n53 VTAIL.n52 185
R174 VTAIL.n55 VTAIL.n54 185
R175 VTAIL.n4 VTAIL.n3 185
R176 VTAIL.n61 VTAIL.n60 185
R177 VTAIL.n197 VTAIL.n196 185
R178 VTAIL.n140 VTAIL.n139 185
R179 VTAIL.n191 VTAIL.n190 185
R180 VTAIL.n189 VTAIL.n188 185
R181 VTAIL.n144 VTAIL.n143 185
R182 VTAIL.n183 VTAIL.n182 185
R183 VTAIL.n181 VTAIL.n180 185
R184 VTAIL.n148 VTAIL.n147 185
R185 VTAIL.n175 VTAIL.n174 185
R186 VTAIL.n173 VTAIL.n172 185
R187 VTAIL.n152 VTAIL.n151 185
R188 VTAIL.n167 VTAIL.n166 185
R189 VTAIL.n165 VTAIL.n164 185
R190 VTAIL.n156 VTAIL.n155 185
R191 VTAIL.n159 VTAIL.n158 185
R192 VTAIL.n131 VTAIL.n130 185
R193 VTAIL.n74 VTAIL.n73 185
R194 VTAIL.n125 VTAIL.n124 185
R195 VTAIL.n123 VTAIL.n122 185
R196 VTAIL.n78 VTAIL.n77 185
R197 VTAIL.n117 VTAIL.n116 185
R198 VTAIL.n115 VTAIL.n114 185
R199 VTAIL.n82 VTAIL.n81 185
R200 VTAIL.n109 VTAIL.n108 185
R201 VTAIL.n107 VTAIL.n106 185
R202 VTAIL.n86 VTAIL.n85 185
R203 VTAIL.n101 VTAIL.n100 185
R204 VTAIL.n99 VTAIL.n98 185
R205 VTAIL.n90 VTAIL.n89 185
R206 VTAIL.n93 VTAIL.n92 185
R207 VTAIL.t18 VTAIL.n219 147.659
R208 VTAIL.t16 VTAIL.n21 147.659
R209 VTAIL.t14 VTAIL.n157 147.659
R210 VTAIL.t6 VTAIL.n91 147.659
R211 VTAIL.n220 VTAIL.n217 104.615
R212 VTAIL.n227 VTAIL.n217 104.615
R213 VTAIL.n228 VTAIL.n227 104.615
R214 VTAIL.n228 VTAIL.n213 104.615
R215 VTAIL.n235 VTAIL.n213 104.615
R216 VTAIL.n236 VTAIL.n235 104.615
R217 VTAIL.n236 VTAIL.n209 104.615
R218 VTAIL.n243 VTAIL.n209 104.615
R219 VTAIL.n244 VTAIL.n243 104.615
R220 VTAIL.n244 VTAIL.n205 104.615
R221 VTAIL.n251 VTAIL.n205 104.615
R222 VTAIL.n252 VTAIL.n251 104.615
R223 VTAIL.n252 VTAIL.n201 104.615
R224 VTAIL.n259 VTAIL.n201 104.615
R225 VTAIL.n22 VTAIL.n19 104.615
R226 VTAIL.n29 VTAIL.n19 104.615
R227 VTAIL.n30 VTAIL.n29 104.615
R228 VTAIL.n30 VTAIL.n15 104.615
R229 VTAIL.n37 VTAIL.n15 104.615
R230 VTAIL.n38 VTAIL.n37 104.615
R231 VTAIL.n38 VTAIL.n11 104.615
R232 VTAIL.n45 VTAIL.n11 104.615
R233 VTAIL.n46 VTAIL.n45 104.615
R234 VTAIL.n46 VTAIL.n7 104.615
R235 VTAIL.n53 VTAIL.n7 104.615
R236 VTAIL.n54 VTAIL.n53 104.615
R237 VTAIL.n54 VTAIL.n3 104.615
R238 VTAIL.n61 VTAIL.n3 104.615
R239 VTAIL.n197 VTAIL.n139 104.615
R240 VTAIL.n190 VTAIL.n139 104.615
R241 VTAIL.n190 VTAIL.n189 104.615
R242 VTAIL.n189 VTAIL.n143 104.615
R243 VTAIL.n182 VTAIL.n143 104.615
R244 VTAIL.n182 VTAIL.n181 104.615
R245 VTAIL.n181 VTAIL.n147 104.615
R246 VTAIL.n174 VTAIL.n147 104.615
R247 VTAIL.n174 VTAIL.n173 104.615
R248 VTAIL.n173 VTAIL.n151 104.615
R249 VTAIL.n166 VTAIL.n151 104.615
R250 VTAIL.n166 VTAIL.n165 104.615
R251 VTAIL.n165 VTAIL.n155 104.615
R252 VTAIL.n158 VTAIL.n155 104.615
R253 VTAIL.n131 VTAIL.n73 104.615
R254 VTAIL.n124 VTAIL.n73 104.615
R255 VTAIL.n124 VTAIL.n123 104.615
R256 VTAIL.n123 VTAIL.n77 104.615
R257 VTAIL.n116 VTAIL.n77 104.615
R258 VTAIL.n116 VTAIL.n115 104.615
R259 VTAIL.n115 VTAIL.n81 104.615
R260 VTAIL.n108 VTAIL.n81 104.615
R261 VTAIL.n108 VTAIL.n107 104.615
R262 VTAIL.n107 VTAIL.n85 104.615
R263 VTAIL.n100 VTAIL.n85 104.615
R264 VTAIL.n100 VTAIL.n99 104.615
R265 VTAIL.n99 VTAIL.n89 104.615
R266 VTAIL.n92 VTAIL.n89 104.615
R267 VTAIL.n220 VTAIL.t18 52.3082
R268 VTAIL.n22 VTAIL.t16 52.3082
R269 VTAIL.n158 VTAIL.t14 52.3082
R270 VTAIL.n92 VTAIL.t6 52.3082
R271 VTAIL.n137 VTAIL.n136 49.1664
R272 VTAIL.n135 VTAIL.n134 49.1664
R273 VTAIL.n71 VTAIL.n70 49.1664
R274 VTAIL.n69 VTAIL.n68 49.1664
R275 VTAIL.n263 VTAIL.n262 49.1662
R276 VTAIL.n1 VTAIL.n0 49.1662
R277 VTAIL.n65 VTAIL.n64 49.1662
R278 VTAIL.n67 VTAIL.n66 49.1662
R279 VTAIL.n261 VTAIL.n260 34.7066
R280 VTAIL.n63 VTAIL.n62 34.7066
R281 VTAIL.n199 VTAIL.n198 34.7066
R282 VTAIL.n133 VTAIL.n132 34.7066
R283 VTAIL.n69 VTAIL.n67 26.9617
R284 VTAIL.n261 VTAIL.n199 24.5221
R285 VTAIL.n221 VTAIL.n219 15.6677
R286 VTAIL.n23 VTAIL.n21 15.6677
R287 VTAIL.n159 VTAIL.n157 15.6677
R288 VTAIL.n93 VTAIL.n91 15.6677
R289 VTAIL.n222 VTAIL.n218 12.8005
R290 VTAIL.n24 VTAIL.n20 12.8005
R291 VTAIL.n160 VTAIL.n156 12.8005
R292 VTAIL.n94 VTAIL.n90 12.8005
R293 VTAIL.n226 VTAIL.n225 12.0247
R294 VTAIL.n28 VTAIL.n27 12.0247
R295 VTAIL.n164 VTAIL.n163 12.0247
R296 VTAIL.n98 VTAIL.n97 12.0247
R297 VTAIL.n229 VTAIL.n216 11.249
R298 VTAIL.n258 VTAIL.n200 11.249
R299 VTAIL.n31 VTAIL.n18 11.249
R300 VTAIL.n60 VTAIL.n2 11.249
R301 VTAIL.n196 VTAIL.n138 11.249
R302 VTAIL.n167 VTAIL.n154 11.249
R303 VTAIL.n130 VTAIL.n72 11.249
R304 VTAIL.n101 VTAIL.n88 11.249
R305 VTAIL.n230 VTAIL.n214 10.4732
R306 VTAIL.n257 VTAIL.n202 10.4732
R307 VTAIL.n32 VTAIL.n16 10.4732
R308 VTAIL.n59 VTAIL.n4 10.4732
R309 VTAIL.n195 VTAIL.n140 10.4732
R310 VTAIL.n168 VTAIL.n152 10.4732
R311 VTAIL.n129 VTAIL.n74 10.4732
R312 VTAIL.n102 VTAIL.n86 10.4732
R313 VTAIL.n234 VTAIL.n233 9.69747
R314 VTAIL.n254 VTAIL.n253 9.69747
R315 VTAIL.n36 VTAIL.n35 9.69747
R316 VTAIL.n56 VTAIL.n55 9.69747
R317 VTAIL.n192 VTAIL.n191 9.69747
R318 VTAIL.n172 VTAIL.n171 9.69747
R319 VTAIL.n126 VTAIL.n125 9.69747
R320 VTAIL.n106 VTAIL.n105 9.69747
R321 VTAIL.n256 VTAIL.n200 9.45567
R322 VTAIL.n58 VTAIL.n2 9.45567
R323 VTAIL.n194 VTAIL.n138 9.45567
R324 VTAIL.n128 VTAIL.n72 9.45567
R325 VTAIL.n208 VTAIL.n207 9.3005
R326 VTAIL.n247 VTAIL.n246 9.3005
R327 VTAIL.n249 VTAIL.n248 9.3005
R328 VTAIL.n204 VTAIL.n203 9.3005
R329 VTAIL.n255 VTAIL.n254 9.3005
R330 VTAIL.n257 VTAIL.n256 9.3005
R331 VTAIL.n239 VTAIL.n238 9.3005
R332 VTAIL.n212 VTAIL.n211 9.3005
R333 VTAIL.n233 VTAIL.n232 9.3005
R334 VTAIL.n231 VTAIL.n230 9.3005
R335 VTAIL.n216 VTAIL.n215 9.3005
R336 VTAIL.n225 VTAIL.n224 9.3005
R337 VTAIL.n223 VTAIL.n222 9.3005
R338 VTAIL.n241 VTAIL.n240 9.3005
R339 VTAIL.n10 VTAIL.n9 9.3005
R340 VTAIL.n49 VTAIL.n48 9.3005
R341 VTAIL.n51 VTAIL.n50 9.3005
R342 VTAIL.n6 VTAIL.n5 9.3005
R343 VTAIL.n57 VTAIL.n56 9.3005
R344 VTAIL.n59 VTAIL.n58 9.3005
R345 VTAIL.n41 VTAIL.n40 9.3005
R346 VTAIL.n14 VTAIL.n13 9.3005
R347 VTAIL.n35 VTAIL.n34 9.3005
R348 VTAIL.n33 VTAIL.n32 9.3005
R349 VTAIL.n18 VTAIL.n17 9.3005
R350 VTAIL.n27 VTAIL.n26 9.3005
R351 VTAIL.n25 VTAIL.n24 9.3005
R352 VTAIL.n43 VTAIL.n42 9.3005
R353 VTAIL.n195 VTAIL.n194 9.3005
R354 VTAIL.n193 VTAIL.n192 9.3005
R355 VTAIL.n142 VTAIL.n141 9.3005
R356 VTAIL.n187 VTAIL.n186 9.3005
R357 VTAIL.n185 VTAIL.n184 9.3005
R358 VTAIL.n146 VTAIL.n145 9.3005
R359 VTAIL.n179 VTAIL.n178 9.3005
R360 VTAIL.n177 VTAIL.n176 9.3005
R361 VTAIL.n150 VTAIL.n149 9.3005
R362 VTAIL.n171 VTAIL.n170 9.3005
R363 VTAIL.n169 VTAIL.n168 9.3005
R364 VTAIL.n154 VTAIL.n153 9.3005
R365 VTAIL.n163 VTAIL.n162 9.3005
R366 VTAIL.n161 VTAIL.n160 9.3005
R367 VTAIL.n119 VTAIL.n118 9.3005
R368 VTAIL.n121 VTAIL.n120 9.3005
R369 VTAIL.n76 VTAIL.n75 9.3005
R370 VTAIL.n127 VTAIL.n126 9.3005
R371 VTAIL.n129 VTAIL.n128 9.3005
R372 VTAIL.n80 VTAIL.n79 9.3005
R373 VTAIL.n113 VTAIL.n112 9.3005
R374 VTAIL.n111 VTAIL.n110 9.3005
R375 VTAIL.n84 VTAIL.n83 9.3005
R376 VTAIL.n105 VTAIL.n104 9.3005
R377 VTAIL.n103 VTAIL.n102 9.3005
R378 VTAIL.n88 VTAIL.n87 9.3005
R379 VTAIL.n97 VTAIL.n96 9.3005
R380 VTAIL.n95 VTAIL.n94 9.3005
R381 VTAIL.n237 VTAIL.n212 8.92171
R382 VTAIL.n250 VTAIL.n204 8.92171
R383 VTAIL.n39 VTAIL.n14 8.92171
R384 VTAIL.n52 VTAIL.n6 8.92171
R385 VTAIL.n188 VTAIL.n142 8.92171
R386 VTAIL.n175 VTAIL.n150 8.92171
R387 VTAIL.n122 VTAIL.n76 8.92171
R388 VTAIL.n109 VTAIL.n84 8.92171
R389 VTAIL.n238 VTAIL.n210 8.14595
R390 VTAIL.n249 VTAIL.n206 8.14595
R391 VTAIL.n40 VTAIL.n12 8.14595
R392 VTAIL.n51 VTAIL.n8 8.14595
R393 VTAIL.n187 VTAIL.n144 8.14595
R394 VTAIL.n176 VTAIL.n148 8.14595
R395 VTAIL.n121 VTAIL.n78 8.14595
R396 VTAIL.n110 VTAIL.n82 8.14595
R397 VTAIL.n242 VTAIL.n241 7.3702
R398 VTAIL.n246 VTAIL.n245 7.3702
R399 VTAIL.n44 VTAIL.n43 7.3702
R400 VTAIL.n48 VTAIL.n47 7.3702
R401 VTAIL.n184 VTAIL.n183 7.3702
R402 VTAIL.n180 VTAIL.n179 7.3702
R403 VTAIL.n118 VTAIL.n117 7.3702
R404 VTAIL.n114 VTAIL.n113 7.3702
R405 VTAIL.n242 VTAIL.n208 6.59444
R406 VTAIL.n245 VTAIL.n208 6.59444
R407 VTAIL.n44 VTAIL.n10 6.59444
R408 VTAIL.n47 VTAIL.n10 6.59444
R409 VTAIL.n183 VTAIL.n146 6.59444
R410 VTAIL.n180 VTAIL.n146 6.59444
R411 VTAIL.n117 VTAIL.n80 6.59444
R412 VTAIL.n114 VTAIL.n80 6.59444
R413 VTAIL.n241 VTAIL.n210 5.81868
R414 VTAIL.n246 VTAIL.n206 5.81868
R415 VTAIL.n43 VTAIL.n12 5.81868
R416 VTAIL.n48 VTAIL.n8 5.81868
R417 VTAIL.n184 VTAIL.n144 5.81868
R418 VTAIL.n179 VTAIL.n148 5.81868
R419 VTAIL.n118 VTAIL.n78 5.81868
R420 VTAIL.n113 VTAIL.n82 5.81868
R421 VTAIL.n238 VTAIL.n237 5.04292
R422 VTAIL.n250 VTAIL.n249 5.04292
R423 VTAIL.n40 VTAIL.n39 5.04292
R424 VTAIL.n52 VTAIL.n51 5.04292
R425 VTAIL.n188 VTAIL.n187 5.04292
R426 VTAIL.n176 VTAIL.n175 5.04292
R427 VTAIL.n122 VTAIL.n121 5.04292
R428 VTAIL.n110 VTAIL.n109 5.04292
R429 VTAIL.n223 VTAIL.n219 4.38563
R430 VTAIL.n25 VTAIL.n21 4.38563
R431 VTAIL.n161 VTAIL.n157 4.38563
R432 VTAIL.n95 VTAIL.n91 4.38563
R433 VTAIL.n234 VTAIL.n212 4.26717
R434 VTAIL.n253 VTAIL.n204 4.26717
R435 VTAIL.n36 VTAIL.n14 4.26717
R436 VTAIL.n55 VTAIL.n6 4.26717
R437 VTAIL.n191 VTAIL.n142 4.26717
R438 VTAIL.n172 VTAIL.n150 4.26717
R439 VTAIL.n125 VTAIL.n76 4.26717
R440 VTAIL.n106 VTAIL.n84 4.26717
R441 VTAIL.n233 VTAIL.n214 3.49141
R442 VTAIL.n254 VTAIL.n202 3.49141
R443 VTAIL.n35 VTAIL.n16 3.49141
R444 VTAIL.n56 VTAIL.n4 3.49141
R445 VTAIL.n192 VTAIL.n140 3.49141
R446 VTAIL.n171 VTAIL.n152 3.49141
R447 VTAIL.n126 VTAIL.n74 3.49141
R448 VTAIL.n105 VTAIL.n86 3.49141
R449 VTAIL.n230 VTAIL.n229 2.71565
R450 VTAIL.n258 VTAIL.n257 2.71565
R451 VTAIL.n32 VTAIL.n31 2.71565
R452 VTAIL.n60 VTAIL.n59 2.71565
R453 VTAIL.n196 VTAIL.n195 2.71565
R454 VTAIL.n168 VTAIL.n167 2.71565
R455 VTAIL.n130 VTAIL.n129 2.71565
R456 VTAIL.n102 VTAIL.n101 2.71565
R457 VTAIL.n71 VTAIL.n69 2.44016
R458 VTAIL.n133 VTAIL.n71 2.44016
R459 VTAIL.n137 VTAIL.n135 2.44016
R460 VTAIL.n199 VTAIL.n137 2.44016
R461 VTAIL.n67 VTAIL.n65 2.44016
R462 VTAIL.n65 VTAIL.n63 2.44016
R463 VTAIL.n263 VTAIL.n261 2.44016
R464 VTAIL.n226 VTAIL.n216 1.93989
R465 VTAIL.n260 VTAIL.n200 1.93989
R466 VTAIL.n28 VTAIL.n18 1.93989
R467 VTAIL.n62 VTAIL.n2 1.93989
R468 VTAIL.n198 VTAIL.n138 1.93989
R469 VTAIL.n164 VTAIL.n154 1.93989
R470 VTAIL.n132 VTAIL.n72 1.93989
R471 VTAIL.n98 VTAIL.n88 1.93989
R472 VTAIL VTAIL.n1 1.88843
R473 VTAIL.n262 VTAIL.t19 1.75738
R474 VTAIL.n262 VTAIL.t17 1.75738
R475 VTAIL.n0 VTAIL.t0 1.75738
R476 VTAIL.n0 VTAIL.t1 1.75738
R477 VTAIL.n64 VTAIL.t7 1.75738
R478 VTAIL.n64 VTAIL.t12 1.75738
R479 VTAIL.n66 VTAIL.t8 1.75738
R480 VTAIL.n66 VTAIL.t10 1.75738
R481 VTAIL.n136 VTAIL.t15 1.75738
R482 VTAIL.n136 VTAIL.t13 1.75738
R483 VTAIL.n134 VTAIL.t9 1.75738
R484 VTAIL.n134 VTAIL.t11 1.75738
R485 VTAIL.n70 VTAIL.t5 1.75738
R486 VTAIL.n70 VTAIL.t2 1.75738
R487 VTAIL.n68 VTAIL.t3 1.75738
R488 VTAIL.n68 VTAIL.t4 1.75738
R489 VTAIL.n135 VTAIL.n133 1.69016
R490 VTAIL.n63 VTAIL.n1 1.69016
R491 VTAIL.n225 VTAIL.n218 1.16414
R492 VTAIL.n27 VTAIL.n20 1.16414
R493 VTAIL.n163 VTAIL.n156 1.16414
R494 VTAIL.n97 VTAIL.n90 1.16414
R495 VTAIL VTAIL.n263 0.552224
R496 VTAIL.n222 VTAIL.n221 0.388379
R497 VTAIL.n24 VTAIL.n23 0.388379
R498 VTAIL.n160 VTAIL.n159 0.388379
R499 VTAIL.n94 VTAIL.n93 0.388379
R500 VTAIL.n224 VTAIL.n223 0.155672
R501 VTAIL.n224 VTAIL.n215 0.155672
R502 VTAIL.n231 VTAIL.n215 0.155672
R503 VTAIL.n232 VTAIL.n231 0.155672
R504 VTAIL.n232 VTAIL.n211 0.155672
R505 VTAIL.n239 VTAIL.n211 0.155672
R506 VTAIL.n240 VTAIL.n239 0.155672
R507 VTAIL.n240 VTAIL.n207 0.155672
R508 VTAIL.n247 VTAIL.n207 0.155672
R509 VTAIL.n248 VTAIL.n247 0.155672
R510 VTAIL.n248 VTAIL.n203 0.155672
R511 VTAIL.n255 VTAIL.n203 0.155672
R512 VTAIL.n256 VTAIL.n255 0.155672
R513 VTAIL.n26 VTAIL.n25 0.155672
R514 VTAIL.n26 VTAIL.n17 0.155672
R515 VTAIL.n33 VTAIL.n17 0.155672
R516 VTAIL.n34 VTAIL.n33 0.155672
R517 VTAIL.n34 VTAIL.n13 0.155672
R518 VTAIL.n41 VTAIL.n13 0.155672
R519 VTAIL.n42 VTAIL.n41 0.155672
R520 VTAIL.n42 VTAIL.n9 0.155672
R521 VTAIL.n49 VTAIL.n9 0.155672
R522 VTAIL.n50 VTAIL.n49 0.155672
R523 VTAIL.n50 VTAIL.n5 0.155672
R524 VTAIL.n57 VTAIL.n5 0.155672
R525 VTAIL.n58 VTAIL.n57 0.155672
R526 VTAIL.n194 VTAIL.n193 0.155672
R527 VTAIL.n193 VTAIL.n141 0.155672
R528 VTAIL.n186 VTAIL.n141 0.155672
R529 VTAIL.n186 VTAIL.n185 0.155672
R530 VTAIL.n185 VTAIL.n145 0.155672
R531 VTAIL.n178 VTAIL.n145 0.155672
R532 VTAIL.n178 VTAIL.n177 0.155672
R533 VTAIL.n177 VTAIL.n149 0.155672
R534 VTAIL.n170 VTAIL.n149 0.155672
R535 VTAIL.n170 VTAIL.n169 0.155672
R536 VTAIL.n169 VTAIL.n153 0.155672
R537 VTAIL.n162 VTAIL.n153 0.155672
R538 VTAIL.n162 VTAIL.n161 0.155672
R539 VTAIL.n128 VTAIL.n127 0.155672
R540 VTAIL.n127 VTAIL.n75 0.155672
R541 VTAIL.n120 VTAIL.n75 0.155672
R542 VTAIL.n120 VTAIL.n119 0.155672
R543 VTAIL.n119 VTAIL.n79 0.155672
R544 VTAIL.n112 VTAIL.n79 0.155672
R545 VTAIL.n112 VTAIL.n111 0.155672
R546 VTAIL.n111 VTAIL.n83 0.155672
R547 VTAIL.n104 VTAIL.n83 0.155672
R548 VTAIL.n104 VTAIL.n103 0.155672
R549 VTAIL.n103 VTAIL.n87 0.155672
R550 VTAIL.n96 VTAIL.n87 0.155672
R551 VTAIL.n96 VTAIL.n95 0.155672
R552 VDD1.n60 VDD1.n59 289.615
R553 VDD1.n123 VDD1.n122 289.615
R554 VDD1.n59 VDD1.n58 185
R555 VDD1.n2 VDD1.n1 185
R556 VDD1.n53 VDD1.n52 185
R557 VDD1.n51 VDD1.n50 185
R558 VDD1.n6 VDD1.n5 185
R559 VDD1.n45 VDD1.n44 185
R560 VDD1.n43 VDD1.n42 185
R561 VDD1.n10 VDD1.n9 185
R562 VDD1.n37 VDD1.n36 185
R563 VDD1.n35 VDD1.n34 185
R564 VDD1.n14 VDD1.n13 185
R565 VDD1.n29 VDD1.n28 185
R566 VDD1.n27 VDD1.n26 185
R567 VDD1.n18 VDD1.n17 185
R568 VDD1.n21 VDD1.n20 185
R569 VDD1.n84 VDD1.n83 185
R570 VDD1.n81 VDD1.n80 185
R571 VDD1.n90 VDD1.n89 185
R572 VDD1.n92 VDD1.n91 185
R573 VDD1.n77 VDD1.n76 185
R574 VDD1.n98 VDD1.n97 185
R575 VDD1.n100 VDD1.n99 185
R576 VDD1.n73 VDD1.n72 185
R577 VDD1.n106 VDD1.n105 185
R578 VDD1.n108 VDD1.n107 185
R579 VDD1.n69 VDD1.n68 185
R580 VDD1.n114 VDD1.n113 185
R581 VDD1.n116 VDD1.n115 185
R582 VDD1.n65 VDD1.n64 185
R583 VDD1.n122 VDD1.n121 185
R584 VDD1.t2 VDD1.n82 147.659
R585 VDD1.t9 VDD1.n19 147.659
R586 VDD1.n59 VDD1.n1 104.615
R587 VDD1.n52 VDD1.n1 104.615
R588 VDD1.n52 VDD1.n51 104.615
R589 VDD1.n51 VDD1.n5 104.615
R590 VDD1.n44 VDD1.n5 104.615
R591 VDD1.n44 VDD1.n43 104.615
R592 VDD1.n43 VDD1.n9 104.615
R593 VDD1.n36 VDD1.n9 104.615
R594 VDD1.n36 VDD1.n35 104.615
R595 VDD1.n35 VDD1.n13 104.615
R596 VDD1.n28 VDD1.n13 104.615
R597 VDD1.n28 VDD1.n27 104.615
R598 VDD1.n27 VDD1.n17 104.615
R599 VDD1.n20 VDD1.n17 104.615
R600 VDD1.n83 VDD1.n80 104.615
R601 VDD1.n90 VDD1.n80 104.615
R602 VDD1.n91 VDD1.n90 104.615
R603 VDD1.n91 VDD1.n76 104.615
R604 VDD1.n98 VDD1.n76 104.615
R605 VDD1.n99 VDD1.n98 104.615
R606 VDD1.n99 VDD1.n72 104.615
R607 VDD1.n106 VDD1.n72 104.615
R608 VDD1.n107 VDD1.n106 104.615
R609 VDD1.n107 VDD1.n68 104.615
R610 VDD1.n114 VDD1.n68 104.615
R611 VDD1.n115 VDD1.n114 104.615
R612 VDD1.n115 VDD1.n64 104.615
R613 VDD1.n122 VDD1.n64 104.615
R614 VDD1.n127 VDD1.n126 67.6194
R615 VDD1.n62 VDD1.n61 65.8451
R616 VDD1.n125 VDD1.n124 65.845
R617 VDD1.n129 VDD1.n128 65.8442
R618 VDD1.n62 VDD1.n60 53.825
R619 VDD1.n125 VDD1.n123 53.825
R620 VDD1.n20 VDD1.t9 52.3082
R621 VDD1.n83 VDD1.t2 52.3082
R622 VDD1.n129 VDD1.n127 46.822
R623 VDD1.n21 VDD1.n19 15.6677
R624 VDD1.n84 VDD1.n82 15.6677
R625 VDD1.n22 VDD1.n18 12.8005
R626 VDD1.n85 VDD1.n81 12.8005
R627 VDD1.n26 VDD1.n25 12.0247
R628 VDD1.n89 VDD1.n88 12.0247
R629 VDD1.n58 VDD1.n0 11.249
R630 VDD1.n29 VDD1.n16 11.249
R631 VDD1.n92 VDD1.n79 11.249
R632 VDD1.n121 VDD1.n63 11.249
R633 VDD1.n57 VDD1.n2 10.4732
R634 VDD1.n30 VDD1.n14 10.4732
R635 VDD1.n93 VDD1.n77 10.4732
R636 VDD1.n120 VDD1.n65 10.4732
R637 VDD1.n54 VDD1.n53 9.69747
R638 VDD1.n34 VDD1.n33 9.69747
R639 VDD1.n97 VDD1.n96 9.69747
R640 VDD1.n117 VDD1.n116 9.69747
R641 VDD1.n56 VDD1.n0 9.45567
R642 VDD1.n119 VDD1.n63 9.45567
R643 VDD1.n47 VDD1.n46 9.3005
R644 VDD1.n49 VDD1.n48 9.3005
R645 VDD1.n4 VDD1.n3 9.3005
R646 VDD1.n55 VDD1.n54 9.3005
R647 VDD1.n57 VDD1.n56 9.3005
R648 VDD1.n8 VDD1.n7 9.3005
R649 VDD1.n41 VDD1.n40 9.3005
R650 VDD1.n39 VDD1.n38 9.3005
R651 VDD1.n12 VDD1.n11 9.3005
R652 VDD1.n33 VDD1.n32 9.3005
R653 VDD1.n31 VDD1.n30 9.3005
R654 VDD1.n16 VDD1.n15 9.3005
R655 VDD1.n25 VDD1.n24 9.3005
R656 VDD1.n23 VDD1.n22 9.3005
R657 VDD1.n71 VDD1.n70 9.3005
R658 VDD1.n110 VDD1.n109 9.3005
R659 VDD1.n112 VDD1.n111 9.3005
R660 VDD1.n67 VDD1.n66 9.3005
R661 VDD1.n118 VDD1.n117 9.3005
R662 VDD1.n120 VDD1.n119 9.3005
R663 VDD1.n102 VDD1.n101 9.3005
R664 VDD1.n75 VDD1.n74 9.3005
R665 VDD1.n96 VDD1.n95 9.3005
R666 VDD1.n94 VDD1.n93 9.3005
R667 VDD1.n79 VDD1.n78 9.3005
R668 VDD1.n88 VDD1.n87 9.3005
R669 VDD1.n86 VDD1.n85 9.3005
R670 VDD1.n104 VDD1.n103 9.3005
R671 VDD1.n50 VDD1.n4 8.92171
R672 VDD1.n37 VDD1.n12 8.92171
R673 VDD1.n100 VDD1.n75 8.92171
R674 VDD1.n113 VDD1.n67 8.92171
R675 VDD1.n49 VDD1.n6 8.14595
R676 VDD1.n38 VDD1.n10 8.14595
R677 VDD1.n101 VDD1.n73 8.14595
R678 VDD1.n112 VDD1.n69 8.14595
R679 VDD1.n46 VDD1.n45 7.3702
R680 VDD1.n42 VDD1.n41 7.3702
R681 VDD1.n105 VDD1.n104 7.3702
R682 VDD1.n109 VDD1.n108 7.3702
R683 VDD1.n45 VDD1.n8 6.59444
R684 VDD1.n42 VDD1.n8 6.59444
R685 VDD1.n105 VDD1.n71 6.59444
R686 VDD1.n108 VDD1.n71 6.59444
R687 VDD1.n46 VDD1.n6 5.81868
R688 VDD1.n41 VDD1.n10 5.81868
R689 VDD1.n104 VDD1.n73 5.81868
R690 VDD1.n109 VDD1.n69 5.81868
R691 VDD1.n50 VDD1.n49 5.04292
R692 VDD1.n38 VDD1.n37 5.04292
R693 VDD1.n101 VDD1.n100 5.04292
R694 VDD1.n113 VDD1.n112 5.04292
R695 VDD1.n86 VDD1.n82 4.38563
R696 VDD1.n23 VDD1.n19 4.38563
R697 VDD1.n53 VDD1.n4 4.26717
R698 VDD1.n34 VDD1.n12 4.26717
R699 VDD1.n97 VDD1.n75 4.26717
R700 VDD1.n116 VDD1.n67 4.26717
R701 VDD1.n54 VDD1.n2 3.49141
R702 VDD1.n33 VDD1.n14 3.49141
R703 VDD1.n96 VDD1.n77 3.49141
R704 VDD1.n117 VDD1.n65 3.49141
R705 VDD1.n58 VDD1.n57 2.71565
R706 VDD1.n30 VDD1.n29 2.71565
R707 VDD1.n93 VDD1.n92 2.71565
R708 VDD1.n121 VDD1.n120 2.71565
R709 VDD1.n60 VDD1.n0 1.93989
R710 VDD1.n26 VDD1.n16 1.93989
R711 VDD1.n89 VDD1.n79 1.93989
R712 VDD1.n123 VDD1.n63 1.93989
R713 VDD1 VDD1.n129 1.77205
R714 VDD1.n128 VDD1.t5 1.75738
R715 VDD1.n128 VDD1.t3 1.75738
R716 VDD1.n61 VDD1.t7 1.75738
R717 VDD1.n61 VDD1.t8 1.75738
R718 VDD1.n126 VDD1.t0 1.75738
R719 VDD1.n126 VDD1.t4 1.75738
R720 VDD1.n124 VDD1.t6 1.75738
R721 VDD1.n124 VDD1.t1 1.75738
R722 VDD1.n25 VDD1.n18 1.16414
R723 VDD1.n88 VDD1.n81 1.16414
R724 VDD1 VDD1.n62 0.668603
R725 VDD1.n127 VDD1.n125 0.555068
R726 VDD1.n22 VDD1.n21 0.388379
R727 VDD1.n85 VDD1.n84 0.388379
R728 VDD1.n56 VDD1.n55 0.155672
R729 VDD1.n55 VDD1.n3 0.155672
R730 VDD1.n48 VDD1.n3 0.155672
R731 VDD1.n48 VDD1.n47 0.155672
R732 VDD1.n47 VDD1.n7 0.155672
R733 VDD1.n40 VDD1.n7 0.155672
R734 VDD1.n40 VDD1.n39 0.155672
R735 VDD1.n39 VDD1.n11 0.155672
R736 VDD1.n32 VDD1.n11 0.155672
R737 VDD1.n32 VDD1.n31 0.155672
R738 VDD1.n31 VDD1.n15 0.155672
R739 VDD1.n24 VDD1.n15 0.155672
R740 VDD1.n24 VDD1.n23 0.155672
R741 VDD1.n87 VDD1.n86 0.155672
R742 VDD1.n87 VDD1.n78 0.155672
R743 VDD1.n94 VDD1.n78 0.155672
R744 VDD1.n95 VDD1.n94 0.155672
R745 VDD1.n95 VDD1.n74 0.155672
R746 VDD1.n102 VDD1.n74 0.155672
R747 VDD1.n103 VDD1.n102 0.155672
R748 VDD1.n103 VDD1.n70 0.155672
R749 VDD1.n110 VDD1.n70 0.155672
R750 VDD1.n111 VDD1.n110 0.155672
R751 VDD1.n111 VDD1.n66 0.155672
R752 VDD1.n118 VDD1.n66 0.155672
R753 VDD1.n119 VDD1.n118 0.155672
R754 B.n745 B.n155 585
R755 B.n155 B.n106 585
R756 B.n747 B.n746 585
R757 B.n749 B.n154 585
R758 B.n752 B.n751 585
R759 B.n753 B.n153 585
R760 B.n755 B.n754 585
R761 B.n757 B.n152 585
R762 B.n760 B.n759 585
R763 B.n761 B.n151 585
R764 B.n763 B.n762 585
R765 B.n765 B.n150 585
R766 B.n768 B.n767 585
R767 B.n769 B.n149 585
R768 B.n771 B.n770 585
R769 B.n773 B.n148 585
R770 B.n776 B.n775 585
R771 B.n777 B.n147 585
R772 B.n779 B.n778 585
R773 B.n781 B.n146 585
R774 B.n784 B.n783 585
R775 B.n785 B.n145 585
R776 B.n787 B.n786 585
R777 B.n789 B.n144 585
R778 B.n792 B.n791 585
R779 B.n793 B.n143 585
R780 B.n795 B.n794 585
R781 B.n797 B.n142 585
R782 B.n800 B.n799 585
R783 B.n801 B.n141 585
R784 B.n803 B.n802 585
R785 B.n805 B.n140 585
R786 B.n808 B.n807 585
R787 B.n809 B.n139 585
R788 B.n811 B.n810 585
R789 B.n813 B.n138 585
R790 B.n816 B.n815 585
R791 B.n817 B.n137 585
R792 B.n819 B.n818 585
R793 B.n821 B.n136 585
R794 B.n824 B.n823 585
R795 B.n826 B.n133 585
R796 B.n828 B.n827 585
R797 B.n830 B.n132 585
R798 B.n833 B.n832 585
R799 B.n834 B.n131 585
R800 B.n836 B.n835 585
R801 B.n838 B.n130 585
R802 B.n841 B.n840 585
R803 B.n842 B.n127 585
R804 B.n845 B.n844 585
R805 B.n847 B.n126 585
R806 B.n850 B.n849 585
R807 B.n851 B.n125 585
R808 B.n853 B.n852 585
R809 B.n855 B.n124 585
R810 B.n858 B.n857 585
R811 B.n859 B.n123 585
R812 B.n861 B.n860 585
R813 B.n863 B.n122 585
R814 B.n866 B.n865 585
R815 B.n867 B.n121 585
R816 B.n869 B.n868 585
R817 B.n871 B.n120 585
R818 B.n874 B.n873 585
R819 B.n875 B.n119 585
R820 B.n877 B.n876 585
R821 B.n879 B.n118 585
R822 B.n882 B.n881 585
R823 B.n883 B.n117 585
R824 B.n885 B.n884 585
R825 B.n887 B.n116 585
R826 B.n890 B.n889 585
R827 B.n891 B.n115 585
R828 B.n893 B.n892 585
R829 B.n895 B.n114 585
R830 B.n898 B.n897 585
R831 B.n899 B.n113 585
R832 B.n901 B.n900 585
R833 B.n903 B.n112 585
R834 B.n906 B.n905 585
R835 B.n907 B.n111 585
R836 B.n909 B.n908 585
R837 B.n911 B.n110 585
R838 B.n914 B.n913 585
R839 B.n915 B.n109 585
R840 B.n917 B.n916 585
R841 B.n919 B.n108 585
R842 B.n922 B.n921 585
R843 B.n923 B.n107 585
R844 B.n744 B.n105 585
R845 B.n926 B.n105 585
R846 B.n743 B.n104 585
R847 B.n927 B.n104 585
R848 B.n742 B.n103 585
R849 B.n928 B.n103 585
R850 B.n741 B.n740 585
R851 B.n740 B.n99 585
R852 B.n739 B.n98 585
R853 B.n934 B.n98 585
R854 B.n738 B.n97 585
R855 B.n935 B.n97 585
R856 B.n737 B.n96 585
R857 B.n936 B.n96 585
R858 B.n736 B.n735 585
R859 B.n735 B.n95 585
R860 B.n734 B.n91 585
R861 B.n942 B.n91 585
R862 B.n733 B.n90 585
R863 B.n943 B.n90 585
R864 B.n732 B.n89 585
R865 B.n944 B.n89 585
R866 B.n731 B.n730 585
R867 B.n730 B.n85 585
R868 B.n729 B.n84 585
R869 B.n950 B.n84 585
R870 B.n728 B.n83 585
R871 B.n951 B.n83 585
R872 B.n727 B.n82 585
R873 B.n952 B.n82 585
R874 B.n726 B.n725 585
R875 B.n725 B.n78 585
R876 B.n724 B.n77 585
R877 B.n958 B.n77 585
R878 B.n723 B.n76 585
R879 B.n959 B.n76 585
R880 B.n722 B.n75 585
R881 B.n960 B.n75 585
R882 B.n721 B.n720 585
R883 B.n720 B.n71 585
R884 B.n719 B.n70 585
R885 B.n966 B.n70 585
R886 B.n718 B.n69 585
R887 B.n967 B.n69 585
R888 B.n717 B.n68 585
R889 B.n968 B.n68 585
R890 B.n716 B.n715 585
R891 B.n715 B.n64 585
R892 B.n714 B.n63 585
R893 B.n974 B.n63 585
R894 B.n713 B.n62 585
R895 B.n975 B.n62 585
R896 B.n712 B.n61 585
R897 B.n976 B.n61 585
R898 B.n711 B.n710 585
R899 B.n710 B.n60 585
R900 B.n709 B.n56 585
R901 B.n982 B.n56 585
R902 B.n708 B.n55 585
R903 B.n983 B.n55 585
R904 B.n707 B.n54 585
R905 B.n984 B.n54 585
R906 B.n706 B.n705 585
R907 B.n705 B.n50 585
R908 B.n704 B.n49 585
R909 B.n990 B.n49 585
R910 B.n703 B.n48 585
R911 B.n991 B.n48 585
R912 B.n702 B.n47 585
R913 B.n992 B.n47 585
R914 B.n701 B.n700 585
R915 B.n700 B.n46 585
R916 B.n699 B.n42 585
R917 B.n998 B.n42 585
R918 B.n698 B.n41 585
R919 B.n999 B.n41 585
R920 B.n697 B.n40 585
R921 B.n1000 B.n40 585
R922 B.n696 B.n695 585
R923 B.n695 B.n36 585
R924 B.n694 B.n35 585
R925 B.n1006 B.n35 585
R926 B.n693 B.n34 585
R927 B.n1007 B.n34 585
R928 B.n692 B.n33 585
R929 B.n1008 B.n33 585
R930 B.n691 B.n690 585
R931 B.n690 B.n32 585
R932 B.n689 B.n28 585
R933 B.n1014 B.n28 585
R934 B.n688 B.n27 585
R935 B.n1015 B.n27 585
R936 B.n687 B.n26 585
R937 B.n1016 B.n26 585
R938 B.n686 B.n685 585
R939 B.n685 B.n22 585
R940 B.n684 B.n21 585
R941 B.n1022 B.n21 585
R942 B.n683 B.n20 585
R943 B.n1023 B.n20 585
R944 B.n682 B.n19 585
R945 B.n1024 B.n19 585
R946 B.n681 B.n680 585
R947 B.n680 B.n15 585
R948 B.n679 B.n14 585
R949 B.n1030 B.n14 585
R950 B.n678 B.n13 585
R951 B.n1031 B.n13 585
R952 B.n677 B.n12 585
R953 B.n1032 B.n12 585
R954 B.n676 B.n675 585
R955 B.n675 B.n8 585
R956 B.n674 B.n7 585
R957 B.n1038 B.n7 585
R958 B.n673 B.n6 585
R959 B.n1039 B.n6 585
R960 B.n672 B.n5 585
R961 B.n1040 B.n5 585
R962 B.n671 B.n670 585
R963 B.n670 B.n4 585
R964 B.n669 B.n156 585
R965 B.n669 B.n668 585
R966 B.n659 B.n157 585
R967 B.n158 B.n157 585
R968 B.n661 B.n660 585
R969 B.n662 B.n661 585
R970 B.n658 B.n163 585
R971 B.n163 B.n162 585
R972 B.n657 B.n656 585
R973 B.n656 B.n655 585
R974 B.n165 B.n164 585
R975 B.n166 B.n165 585
R976 B.n648 B.n647 585
R977 B.n649 B.n648 585
R978 B.n646 B.n171 585
R979 B.n171 B.n170 585
R980 B.n645 B.n644 585
R981 B.n644 B.n643 585
R982 B.n173 B.n172 585
R983 B.n174 B.n173 585
R984 B.n636 B.n635 585
R985 B.n637 B.n636 585
R986 B.n634 B.n179 585
R987 B.n179 B.n178 585
R988 B.n633 B.n632 585
R989 B.n632 B.n631 585
R990 B.n181 B.n180 585
R991 B.n624 B.n181 585
R992 B.n623 B.n622 585
R993 B.n625 B.n623 585
R994 B.n621 B.n186 585
R995 B.n186 B.n185 585
R996 B.n620 B.n619 585
R997 B.n619 B.n618 585
R998 B.n188 B.n187 585
R999 B.n189 B.n188 585
R1000 B.n611 B.n610 585
R1001 B.n612 B.n611 585
R1002 B.n609 B.n194 585
R1003 B.n194 B.n193 585
R1004 B.n608 B.n607 585
R1005 B.n607 B.n606 585
R1006 B.n196 B.n195 585
R1007 B.n599 B.n196 585
R1008 B.n598 B.n597 585
R1009 B.n600 B.n598 585
R1010 B.n596 B.n201 585
R1011 B.n201 B.n200 585
R1012 B.n595 B.n594 585
R1013 B.n594 B.n593 585
R1014 B.n203 B.n202 585
R1015 B.n204 B.n203 585
R1016 B.n586 B.n585 585
R1017 B.n587 B.n586 585
R1018 B.n584 B.n209 585
R1019 B.n209 B.n208 585
R1020 B.n583 B.n582 585
R1021 B.n582 B.n581 585
R1022 B.n211 B.n210 585
R1023 B.n574 B.n211 585
R1024 B.n573 B.n572 585
R1025 B.n575 B.n573 585
R1026 B.n571 B.n216 585
R1027 B.n216 B.n215 585
R1028 B.n570 B.n569 585
R1029 B.n569 B.n568 585
R1030 B.n218 B.n217 585
R1031 B.n219 B.n218 585
R1032 B.n561 B.n560 585
R1033 B.n562 B.n561 585
R1034 B.n559 B.n224 585
R1035 B.n224 B.n223 585
R1036 B.n558 B.n557 585
R1037 B.n557 B.n556 585
R1038 B.n226 B.n225 585
R1039 B.n227 B.n226 585
R1040 B.n549 B.n548 585
R1041 B.n550 B.n549 585
R1042 B.n547 B.n232 585
R1043 B.n232 B.n231 585
R1044 B.n546 B.n545 585
R1045 B.n545 B.n544 585
R1046 B.n234 B.n233 585
R1047 B.n235 B.n234 585
R1048 B.n537 B.n536 585
R1049 B.n538 B.n537 585
R1050 B.n535 B.n240 585
R1051 B.n240 B.n239 585
R1052 B.n534 B.n533 585
R1053 B.n533 B.n532 585
R1054 B.n242 B.n241 585
R1055 B.n243 B.n242 585
R1056 B.n525 B.n524 585
R1057 B.n526 B.n525 585
R1058 B.n523 B.n248 585
R1059 B.n248 B.n247 585
R1060 B.n522 B.n521 585
R1061 B.n521 B.n520 585
R1062 B.n250 B.n249 585
R1063 B.n513 B.n250 585
R1064 B.n512 B.n511 585
R1065 B.n514 B.n512 585
R1066 B.n510 B.n255 585
R1067 B.n255 B.n254 585
R1068 B.n509 B.n508 585
R1069 B.n508 B.n507 585
R1070 B.n257 B.n256 585
R1071 B.n258 B.n257 585
R1072 B.n500 B.n499 585
R1073 B.n501 B.n500 585
R1074 B.n498 B.n263 585
R1075 B.n263 B.n262 585
R1076 B.n497 B.n496 585
R1077 B.n496 B.n495 585
R1078 B.n492 B.n267 585
R1079 B.n491 B.n490 585
R1080 B.n488 B.n268 585
R1081 B.n488 B.n266 585
R1082 B.n487 B.n486 585
R1083 B.n485 B.n484 585
R1084 B.n483 B.n270 585
R1085 B.n481 B.n480 585
R1086 B.n479 B.n271 585
R1087 B.n478 B.n477 585
R1088 B.n475 B.n272 585
R1089 B.n473 B.n472 585
R1090 B.n471 B.n273 585
R1091 B.n470 B.n469 585
R1092 B.n467 B.n274 585
R1093 B.n465 B.n464 585
R1094 B.n463 B.n275 585
R1095 B.n462 B.n461 585
R1096 B.n459 B.n276 585
R1097 B.n457 B.n456 585
R1098 B.n455 B.n277 585
R1099 B.n454 B.n453 585
R1100 B.n451 B.n278 585
R1101 B.n449 B.n448 585
R1102 B.n447 B.n279 585
R1103 B.n446 B.n445 585
R1104 B.n443 B.n280 585
R1105 B.n441 B.n440 585
R1106 B.n439 B.n281 585
R1107 B.n438 B.n437 585
R1108 B.n435 B.n282 585
R1109 B.n433 B.n432 585
R1110 B.n431 B.n283 585
R1111 B.n430 B.n429 585
R1112 B.n427 B.n284 585
R1113 B.n425 B.n424 585
R1114 B.n423 B.n285 585
R1115 B.n422 B.n421 585
R1116 B.n419 B.n286 585
R1117 B.n417 B.n416 585
R1118 B.n415 B.n287 585
R1119 B.n413 B.n412 585
R1120 B.n410 B.n290 585
R1121 B.n408 B.n407 585
R1122 B.n406 B.n291 585
R1123 B.n405 B.n404 585
R1124 B.n402 B.n292 585
R1125 B.n400 B.n399 585
R1126 B.n398 B.n293 585
R1127 B.n397 B.n396 585
R1128 B.n394 B.n393 585
R1129 B.n392 B.n391 585
R1130 B.n390 B.n298 585
R1131 B.n388 B.n387 585
R1132 B.n386 B.n299 585
R1133 B.n385 B.n384 585
R1134 B.n382 B.n300 585
R1135 B.n380 B.n379 585
R1136 B.n378 B.n301 585
R1137 B.n377 B.n376 585
R1138 B.n374 B.n302 585
R1139 B.n372 B.n371 585
R1140 B.n370 B.n303 585
R1141 B.n369 B.n368 585
R1142 B.n366 B.n304 585
R1143 B.n364 B.n363 585
R1144 B.n362 B.n305 585
R1145 B.n361 B.n360 585
R1146 B.n358 B.n306 585
R1147 B.n356 B.n355 585
R1148 B.n354 B.n307 585
R1149 B.n353 B.n352 585
R1150 B.n350 B.n308 585
R1151 B.n348 B.n347 585
R1152 B.n346 B.n309 585
R1153 B.n345 B.n344 585
R1154 B.n342 B.n310 585
R1155 B.n340 B.n339 585
R1156 B.n338 B.n311 585
R1157 B.n337 B.n336 585
R1158 B.n334 B.n312 585
R1159 B.n332 B.n331 585
R1160 B.n330 B.n313 585
R1161 B.n329 B.n328 585
R1162 B.n326 B.n314 585
R1163 B.n324 B.n323 585
R1164 B.n322 B.n315 585
R1165 B.n321 B.n320 585
R1166 B.n318 B.n316 585
R1167 B.n265 B.n264 585
R1168 B.n494 B.n493 585
R1169 B.n495 B.n494 585
R1170 B.n261 B.n260 585
R1171 B.n262 B.n261 585
R1172 B.n503 B.n502 585
R1173 B.n502 B.n501 585
R1174 B.n504 B.n259 585
R1175 B.n259 B.n258 585
R1176 B.n506 B.n505 585
R1177 B.n507 B.n506 585
R1178 B.n253 B.n252 585
R1179 B.n254 B.n253 585
R1180 B.n516 B.n515 585
R1181 B.n515 B.n514 585
R1182 B.n517 B.n251 585
R1183 B.n513 B.n251 585
R1184 B.n519 B.n518 585
R1185 B.n520 B.n519 585
R1186 B.n246 B.n245 585
R1187 B.n247 B.n246 585
R1188 B.n528 B.n527 585
R1189 B.n527 B.n526 585
R1190 B.n529 B.n244 585
R1191 B.n244 B.n243 585
R1192 B.n531 B.n530 585
R1193 B.n532 B.n531 585
R1194 B.n238 B.n237 585
R1195 B.n239 B.n238 585
R1196 B.n540 B.n539 585
R1197 B.n539 B.n538 585
R1198 B.n541 B.n236 585
R1199 B.n236 B.n235 585
R1200 B.n543 B.n542 585
R1201 B.n544 B.n543 585
R1202 B.n230 B.n229 585
R1203 B.n231 B.n230 585
R1204 B.n552 B.n551 585
R1205 B.n551 B.n550 585
R1206 B.n553 B.n228 585
R1207 B.n228 B.n227 585
R1208 B.n555 B.n554 585
R1209 B.n556 B.n555 585
R1210 B.n222 B.n221 585
R1211 B.n223 B.n222 585
R1212 B.n564 B.n563 585
R1213 B.n563 B.n562 585
R1214 B.n565 B.n220 585
R1215 B.n220 B.n219 585
R1216 B.n567 B.n566 585
R1217 B.n568 B.n567 585
R1218 B.n214 B.n213 585
R1219 B.n215 B.n214 585
R1220 B.n577 B.n576 585
R1221 B.n576 B.n575 585
R1222 B.n578 B.n212 585
R1223 B.n574 B.n212 585
R1224 B.n580 B.n579 585
R1225 B.n581 B.n580 585
R1226 B.n207 B.n206 585
R1227 B.n208 B.n207 585
R1228 B.n589 B.n588 585
R1229 B.n588 B.n587 585
R1230 B.n590 B.n205 585
R1231 B.n205 B.n204 585
R1232 B.n592 B.n591 585
R1233 B.n593 B.n592 585
R1234 B.n199 B.n198 585
R1235 B.n200 B.n199 585
R1236 B.n602 B.n601 585
R1237 B.n601 B.n600 585
R1238 B.n603 B.n197 585
R1239 B.n599 B.n197 585
R1240 B.n605 B.n604 585
R1241 B.n606 B.n605 585
R1242 B.n192 B.n191 585
R1243 B.n193 B.n192 585
R1244 B.n614 B.n613 585
R1245 B.n613 B.n612 585
R1246 B.n615 B.n190 585
R1247 B.n190 B.n189 585
R1248 B.n617 B.n616 585
R1249 B.n618 B.n617 585
R1250 B.n184 B.n183 585
R1251 B.n185 B.n184 585
R1252 B.n627 B.n626 585
R1253 B.n626 B.n625 585
R1254 B.n628 B.n182 585
R1255 B.n624 B.n182 585
R1256 B.n630 B.n629 585
R1257 B.n631 B.n630 585
R1258 B.n177 B.n176 585
R1259 B.n178 B.n177 585
R1260 B.n639 B.n638 585
R1261 B.n638 B.n637 585
R1262 B.n640 B.n175 585
R1263 B.n175 B.n174 585
R1264 B.n642 B.n641 585
R1265 B.n643 B.n642 585
R1266 B.n169 B.n168 585
R1267 B.n170 B.n169 585
R1268 B.n651 B.n650 585
R1269 B.n650 B.n649 585
R1270 B.n652 B.n167 585
R1271 B.n167 B.n166 585
R1272 B.n654 B.n653 585
R1273 B.n655 B.n654 585
R1274 B.n161 B.n160 585
R1275 B.n162 B.n161 585
R1276 B.n664 B.n663 585
R1277 B.n663 B.n662 585
R1278 B.n665 B.n159 585
R1279 B.n159 B.n158 585
R1280 B.n667 B.n666 585
R1281 B.n668 B.n667 585
R1282 B.n2 B.n0 585
R1283 B.n4 B.n2 585
R1284 B.n3 B.n1 585
R1285 B.n1039 B.n3 585
R1286 B.n1037 B.n1036 585
R1287 B.n1038 B.n1037 585
R1288 B.n1035 B.n9 585
R1289 B.n9 B.n8 585
R1290 B.n1034 B.n1033 585
R1291 B.n1033 B.n1032 585
R1292 B.n11 B.n10 585
R1293 B.n1031 B.n11 585
R1294 B.n1029 B.n1028 585
R1295 B.n1030 B.n1029 585
R1296 B.n1027 B.n16 585
R1297 B.n16 B.n15 585
R1298 B.n1026 B.n1025 585
R1299 B.n1025 B.n1024 585
R1300 B.n18 B.n17 585
R1301 B.n1023 B.n18 585
R1302 B.n1021 B.n1020 585
R1303 B.n1022 B.n1021 585
R1304 B.n1019 B.n23 585
R1305 B.n23 B.n22 585
R1306 B.n1018 B.n1017 585
R1307 B.n1017 B.n1016 585
R1308 B.n25 B.n24 585
R1309 B.n1015 B.n25 585
R1310 B.n1013 B.n1012 585
R1311 B.n1014 B.n1013 585
R1312 B.n1011 B.n29 585
R1313 B.n32 B.n29 585
R1314 B.n1010 B.n1009 585
R1315 B.n1009 B.n1008 585
R1316 B.n31 B.n30 585
R1317 B.n1007 B.n31 585
R1318 B.n1005 B.n1004 585
R1319 B.n1006 B.n1005 585
R1320 B.n1003 B.n37 585
R1321 B.n37 B.n36 585
R1322 B.n1002 B.n1001 585
R1323 B.n1001 B.n1000 585
R1324 B.n39 B.n38 585
R1325 B.n999 B.n39 585
R1326 B.n997 B.n996 585
R1327 B.n998 B.n997 585
R1328 B.n995 B.n43 585
R1329 B.n46 B.n43 585
R1330 B.n994 B.n993 585
R1331 B.n993 B.n992 585
R1332 B.n45 B.n44 585
R1333 B.n991 B.n45 585
R1334 B.n989 B.n988 585
R1335 B.n990 B.n989 585
R1336 B.n987 B.n51 585
R1337 B.n51 B.n50 585
R1338 B.n986 B.n985 585
R1339 B.n985 B.n984 585
R1340 B.n53 B.n52 585
R1341 B.n983 B.n53 585
R1342 B.n981 B.n980 585
R1343 B.n982 B.n981 585
R1344 B.n979 B.n57 585
R1345 B.n60 B.n57 585
R1346 B.n978 B.n977 585
R1347 B.n977 B.n976 585
R1348 B.n59 B.n58 585
R1349 B.n975 B.n59 585
R1350 B.n973 B.n972 585
R1351 B.n974 B.n973 585
R1352 B.n971 B.n65 585
R1353 B.n65 B.n64 585
R1354 B.n970 B.n969 585
R1355 B.n969 B.n968 585
R1356 B.n67 B.n66 585
R1357 B.n967 B.n67 585
R1358 B.n965 B.n964 585
R1359 B.n966 B.n965 585
R1360 B.n963 B.n72 585
R1361 B.n72 B.n71 585
R1362 B.n962 B.n961 585
R1363 B.n961 B.n960 585
R1364 B.n74 B.n73 585
R1365 B.n959 B.n74 585
R1366 B.n957 B.n956 585
R1367 B.n958 B.n957 585
R1368 B.n955 B.n79 585
R1369 B.n79 B.n78 585
R1370 B.n954 B.n953 585
R1371 B.n953 B.n952 585
R1372 B.n81 B.n80 585
R1373 B.n951 B.n81 585
R1374 B.n949 B.n948 585
R1375 B.n950 B.n949 585
R1376 B.n947 B.n86 585
R1377 B.n86 B.n85 585
R1378 B.n946 B.n945 585
R1379 B.n945 B.n944 585
R1380 B.n88 B.n87 585
R1381 B.n943 B.n88 585
R1382 B.n941 B.n940 585
R1383 B.n942 B.n941 585
R1384 B.n939 B.n92 585
R1385 B.n95 B.n92 585
R1386 B.n938 B.n937 585
R1387 B.n937 B.n936 585
R1388 B.n94 B.n93 585
R1389 B.n935 B.n94 585
R1390 B.n933 B.n932 585
R1391 B.n934 B.n933 585
R1392 B.n931 B.n100 585
R1393 B.n100 B.n99 585
R1394 B.n930 B.n929 585
R1395 B.n929 B.n928 585
R1396 B.n102 B.n101 585
R1397 B.n927 B.n102 585
R1398 B.n925 B.n924 585
R1399 B.n926 B.n925 585
R1400 B.n1042 B.n1041 585
R1401 B.n1041 B.n1040 585
R1402 B.n494 B.n267 468.476
R1403 B.n925 B.n107 468.476
R1404 B.n496 B.n265 468.476
R1405 B.n155 B.n105 468.476
R1406 B.n294 B.t20 324.211
R1407 B.n134 B.t12 324.211
R1408 B.n288 B.t23 324.211
R1409 B.n128 B.t15 324.211
R1410 B.n294 B.t17 316.534
R1411 B.n288 B.t21 316.534
R1412 B.n128 B.t14 316.534
R1413 B.n134 B.t10 316.534
R1414 B.n295 B.t19 269.327
R1415 B.n135 B.t13 269.327
R1416 B.n289 B.t22 269.327
R1417 B.n129 B.t16 269.327
R1418 B.n748 B.n106 256.663
R1419 B.n750 B.n106 256.663
R1420 B.n756 B.n106 256.663
R1421 B.n758 B.n106 256.663
R1422 B.n764 B.n106 256.663
R1423 B.n766 B.n106 256.663
R1424 B.n772 B.n106 256.663
R1425 B.n774 B.n106 256.663
R1426 B.n780 B.n106 256.663
R1427 B.n782 B.n106 256.663
R1428 B.n788 B.n106 256.663
R1429 B.n790 B.n106 256.663
R1430 B.n796 B.n106 256.663
R1431 B.n798 B.n106 256.663
R1432 B.n804 B.n106 256.663
R1433 B.n806 B.n106 256.663
R1434 B.n812 B.n106 256.663
R1435 B.n814 B.n106 256.663
R1436 B.n820 B.n106 256.663
R1437 B.n822 B.n106 256.663
R1438 B.n829 B.n106 256.663
R1439 B.n831 B.n106 256.663
R1440 B.n837 B.n106 256.663
R1441 B.n839 B.n106 256.663
R1442 B.n846 B.n106 256.663
R1443 B.n848 B.n106 256.663
R1444 B.n854 B.n106 256.663
R1445 B.n856 B.n106 256.663
R1446 B.n862 B.n106 256.663
R1447 B.n864 B.n106 256.663
R1448 B.n870 B.n106 256.663
R1449 B.n872 B.n106 256.663
R1450 B.n878 B.n106 256.663
R1451 B.n880 B.n106 256.663
R1452 B.n886 B.n106 256.663
R1453 B.n888 B.n106 256.663
R1454 B.n894 B.n106 256.663
R1455 B.n896 B.n106 256.663
R1456 B.n902 B.n106 256.663
R1457 B.n904 B.n106 256.663
R1458 B.n910 B.n106 256.663
R1459 B.n912 B.n106 256.663
R1460 B.n918 B.n106 256.663
R1461 B.n920 B.n106 256.663
R1462 B.n489 B.n266 256.663
R1463 B.n269 B.n266 256.663
R1464 B.n482 B.n266 256.663
R1465 B.n476 B.n266 256.663
R1466 B.n474 B.n266 256.663
R1467 B.n468 B.n266 256.663
R1468 B.n466 B.n266 256.663
R1469 B.n460 B.n266 256.663
R1470 B.n458 B.n266 256.663
R1471 B.n452 B.n266 256.663
R1472 B.n450 B.n266 256.663
R1473 B.n444 B.n266 256.663
R1474 B.n442 B.n266 256.663
R1475 B.n436 B.n266 256.663
R1476 B.n434 B.n266 256.663
R1477 B.n428 B.n266 256.663
R1478 B.n426 B.n266 256.663
R1479 B.n420 B.n266 256.663
R1480 B.n418 B.n266 256.663
R1481 B.n411 B.n266 256.663
R1482 B.n409 B.n266 256.663
R1483 B.n403 B.n266 256.663
R1484 B.n401 B.n266 256.663
R1485 B.n395 B.n266 256.663
R1486 B.n297 B.n266 256.663
R1487 B.n389 B.n266 256.663
R1488 B.n383 B.n266 256.663
R1489 B.n381 B.n266 256.663
R1490 B.n375 B.n266 256.663
R1491 B.n373 B.n266 256.663
R1492 B.n367 B.n266 256.663
R1493 B.n365 B.n266 256.663
R1494 B.n359 B.n266 256.663
R1495 B.n357 B.n266 256.663
R1496 B.n351 B.n266 256.663
R1497 B.n349 B.n266 256.663
R1498 B.n343 B.n266 256.663
R1499 B.n341 B.n266 256.663
R1500 B.n335 B.n266 256.663
R1501 B.n333 B.n266 256.663
R1502 B.n327 B.n266 256.663
R1503 B.n325 B.n266 256.663
R1504 B.n319 B.n266 256.663
R1505 B.n317 B.n266 256.663
R1506 B.n494 B.n261 163.367
R1507 B.n502 B.n261 163.367
R1508 B.n502 B.n259 163.367
R1509 B.n506 B.n259 163.367
R1510 B.n506 B.n253 163.367
R1511 B.n515 B.n253 163.367
R1512 B.n515 B.n251 163.367
R1513 B.n519 B.n251 163.367
R1514 B.n519 B.n246 163.367
R1515 B.n527 B.n246 163.367
R1516 B.n527 B.n244 163.367
R1517 B.n531 B.n244 163.367
R1518 B.n531 B.n238 163.367
R1519 B.n539 B.n238 163.367
R1520 B.n539 B.n236 163.367
R1521 B.n543 B.n236 163.367
R1522 B.n543 B.n230 163.367
R1523 B.n551 B.n230 163.367
R1524 B.n551 B.n228 163.367
R1525 B.n555 B.n228 163.367
R1526 B.n555 B.n222 163.367
R1527 B.n563 B.n222 163.367
R1528 B.n563 B.n220 163.367
R1529 B.n567 B.n220 163.367
R1530 B.n567 B.n214 163.367
R1531 B.n576 B.n214 163.367
R1532 B.n576 B.n212 163.367
R1533 B.n580 B.n212 163.367
R1534 B.n580 B.n207 163.367
R1535 B.n588 B.n207 163.367
R1536 B.n588 B.n205 163.367
R1537 B.n592 B.n205 163.367
R1538 B.n592 B.n199 163.367
R1539 B.n601 B.n199 163.367
R1540 B.n601 B.n197 163.367
R1541 B.n605 B.n197 163.367
R1542 B.n605 B.n192 163.367
R1543 B.n613 B.n192 163.367
R1544 B.n613 B.n190 163.367
R1545 B.n617 B.n190 163.367
R1546 B.n617 B.n184 163.367
R1547 B.n626 B.n184 163.367
R1548 B.n626 B.n182 163.367
R1549 B.n630 B.n182 163.367
R1550 B.n630 B.n177 163.367
R1551 B.n638 B.n177 163.367
R1552 B.n638 B.n175 163.367
R1553 B.n642 B.n175 163.367
R1554 B.n642 B.n169 163.367
R1555 B.n650 B.n169 163.367
R1556 B.n650 B.n167 163.367
R1557 B.n654 B.n167 163.367
R1558 B.n654 B.n161 163.367
R1559 B.n663 B.n161 163.367
R1560 B.n663 B.n159 163.367
R1561 B.n667 B.n159 163.367
R1562 B.n667 B.n2 163.367
R1563 B.n1041 B.n2 163.367
R1564 B.n1041 B.n3 163.367
R1565 B.n1037 B.n3 163.367
R1566 B.n1037 B.n9 163.367
R1567 B.n1033 B.n9 163.367
R1568 B.n1033 B.n11 163.367
R1569 B.n1029 B.n11 163.367
R1570 B.n1029 B.n16 163.367
R1571 B.n1025 B.n16 163.367
R1572 B.n1025 B.n18 163.367
R1573 B.n1021 B.n18 163.367
R1574 B.n1021 B.n23 163.367
R1575 B.n1017 B.n23 163.367
R1576 B.n1017 B.n25 163.367
R1577 B.n1013 B.n25 163.367
R1578 B.n1013 B.n29 163.367
R1579 B.n1009 B.n29 163.367
R1580 B.n1009 B.n31 163.367
R1581 B.n1005 B.n31 163.367
R1582 B.n1005 B.n37 163.367
R1583 B.n1001 B.n37 163.367
R1584 B.n1001 B.n39 163.367
R1585 B.n997 B.n39 163.367
R1586 B.n997 B.n43 163.367
R1587 B.n993 B.n43 163.367
R1588 B.n993 B.n45 163.367
R1589 B.n989 B.n45 163.367
R1590 B.n989 B.n51 163.367
R1591 B.n985 B.n51 163.367
R1592 B.n985 B.n53 163.367
R1593 B.n981 B.n53 163.367
R1594 B.n981 B.n57 163.367
R1595 B.n977 B.n57 163.367
R1596 B.n977 B.n59 163.367
R1597 B.n973 B.n59 163.367
R1598 B.n973 B.n65 163.367
R1599 B.n969 B.n65 163.367
R1600 B.n969 B.n67 163.367
R1601 B.n965 B.n67 163.367
R1602 B.n965 B.n72 163.367
R1603 B.n961 B.n72 163.367
R1604 B.n961 B.n74 163.367
R1605 B.n957 B.n74 163.367
R1606 B.n957 B.n79 163.367
R1607 B.n953 B.n79 163.367
R1608 B.n953 B.n81 163.367
R1609 B.n949 B.n81 163.367
R1610 B.n949 B.n86 163.367
R1611 B.n945 B.n86 163.367
R1612 B.n945 B.n88 163.367
R1613 B.n941 B.n88 163.367
R1614 B.n941 B.n92 163.367
R1615 B.n937 B.n92 163.367
R1616 B.n937 B.n94 163.367
R1617 B.n933 B.n94 163.367
R1618 B.n933 B.n100 163.367
R1619 B.n929 B.n100 163.367
R1620 B.n929 B.n102 163.367
R1621 B.n925 B.n102 163.367
R1622 B.n490 B.n488 163.367
R1623 B.n488 B.n487 163.367
R1624 B.n484 B.n483 163.367
R1625 B.n481 B.n271 163.367
R1626 B.n477 B.n475 163.367
R1627 B.n473 B.n273 163.367
R1628 B.n469 B.n467 163.367
R1629 B.n465 B.n275 163.367
R1630 B.n461 B.n459 163.367
R1631 B.n457 B.n277 163.367
R1632 B.n453 B.n451 163.367
R1633 B.n449 B.n279 163.367
R1634 B.n445 B.n443 163.367
R1635 B.n441 B.n281 163.367
R1636 B.n437 B.n435 163.367
R1637 B.n433 B.n283 163.367
R1638 B.n429 B.n427 163.367
R1639 B.n425 B.n285 163.367
R1640 B.n421 B.n419 163.367
R1641 B.n417 B.n287 163.367
R1642 B.n412 B.n410 163.367
R1643 B.n408 B.n291 163.367
R1644 B.n404 B.n402 163.367
R1645 B.n400 B.n293 163.367
R1646 B.n396 B.n394 163.367
R1647 B.n391 B.n390 163.367
R1648 B.n388 B.n299 163.367
R1649 B.n384 B.n382 163.367
R1650 B.n380 B.n301 163.367
R1651 B.n376 B.n374 163.367
R1652 B.n372 B.n303 163.367
R1653 B.n368 B.n366 163.367
R1654 B.n364 B.n305 163.367
R1655 B.n360 B.n358 163.367
R1656 B.n356 B.n307 163.367
R1657 B.n352 B.n350 163.367
R1658 B.n348 B.n309 163.367
R1659 B.n344 B.n342 163.367
R1660 B.n340 B.n311 163.367
R1661 B.n336 B.n334 163.367
R1662 B.n332 B.n313 163.367
R1663 B.n328 B.n326 163.367
R1664 B.n324 B.n315 163.367
R1665 B.n320 B.n318 163.367
R1666 B.n496 B.n263 163.367
R1667 B.n500 B.n263 163.367
R1668 B.n500 B.n257 163.367
R1669 B.n508 B.n257 163.367
R1670 B.n508 B.n255 163.367
R1671 B.n512 B.n255 163.367
R1672 B.n512 B.n250 163.367
R1673 B.n521 B.n250 163.367
R1674 B.n521 B.n248 163.367
R1675 B.n525 B.n248 163.367
R1676 B.n525 B.n242 163.367
R1677 B.n533 B.n242 163.367
R1678 B.n533 B.n240 163.367
R1679 B.n537 B.n240 163.367
R1680 B.n537 B.n234 163.367
R1681 B.n545 B.n234 163.367
R1682 B.n545 B.n232 163.367
R1683 B.n549 B.n232 163.367
R1684 B.n549 B.n226 163.367
R1685 B.n557 B.n226 163.367
R1686 B.n557 B.n224 163.367
R1687 B.n561 B.n224 163.367
R1688 B.n561 B.n218 163.367
R1689 B.n569 B.n218 163.367
R1690 B.n569 B.n216 163.367
R1691 B.n573 B.n216 163.367
R1692 B.n573 B.n211 163.367
R1693 B.n582 B.n211 163.367
R1694 B.n582 B.n209 163.367
R1695 B.n586 B.n209 163.367
R1696 B.n586 B.n203 163.367
R1697 B.n594 B.n203 163.367
R1698 B.n594 B.n201 163.367
R1699 B.n598 B.n201 163.367
R1700 B.n598 B.n196 163.367
R1701 B.n607 B.n196 163.367
R1702 B.n607 B.n194 163.367
R1703 B.n611 B.n194 163.367
R1704 B.n611 B.n188 163.367
R1705 B.n619 B.n188 163.367
R1706 B.n619 B.n186 163.367
R1707 B.n623 B.n186 163.367
R1708 B.n623 B.n181 163.367
R1709 B.n632 B.n181 163.367
R1710 B.n632 B.n179 163.367
R1711 B.n636 B.n179 163.367
R1712 B.n636 B.n173 163.367
R1713 B.n644 B.n173 163.367
R1714 B.n644 B.n171 163.367
R1715 B.n648 B.n171 163.367
R1716 B.n648 B.n165 163.367
R1717 B.n656 B.n165 163.367
R1718 B.n656 B.n163 163.367
R1719 B.n661 B.n163 163.367
R1720 B.n661 B.n157 163.367
R1721 B.n669 B.n157 163.367
R1722 B.n670 B.n669 163.367
R1723 B.n670 B.n5 163.367
R1724 B.n6 B.n5 163.367
R1725 B.n7 B.n6 163.367
R1726 B.n675 B.n7 163.367
R1727 B.n675 B.n12 163.367
R1728 B.n13 B.n12 163.367
R1729 B.n14 B.n13 163.367
R1730 B.n680 B.n14 163.367
R1731 B.n680 B.n19 163.367
R1732 B.n20 B.n19 163.367
R1733 B.n21 B.n20 163.367
R1734 B.n685 B.n21 163.367
R1735 B.n685 B.n26 163.367
R1736 B.n27 B.n26 163.367
R1737 B.n28 B.n27 163.367
R1738 B.n690 B.n28 163.367
R1739 B.n690 B.n33 163.367
R1740 B.n34 B.n33 163.367
R1741 B.n35 B.n34 163.367
R1742 B.n695 B.n35 163.367
R1743 B.n695 B.n40 163.367
R1744 B.n41 B.n40 163.367
R1745 B.n42 B.n41 163.367
R1746 B.n700 B.n42 163.367
R1747 B.n700 B.n47 163.367
R1748 B.n48 B.n47 163.367
R1749 B.n49 B.n48 163.367
R1750 B.n705 B.n49 163.367
R1751 B.n705 B.n54 163.367
R1752 B.n55 B.n54 163.367
R1753 B.n56 B.n55 163.367
R1754 B.n710 B.n56 163.367
R1755 B.n710 B.n61 163.367
R1756 B.n62 B.n61 163.367
R1757 B.n63 B.n62 163.367
R1758 B.n715 B.n63 163.367
R1759 B.n715 B.n68 163.367
R1760 B.n69 B.n68 163.367
R1761 B.n70 B.n69 163.367
R1762 B.n720 B.n70 163.367
R1763 B.n720 B.n75 163.367
R1764 B.n76 B.n75 163.367
R1765 B.n77 B.n76 163.367
R1766 B.n725 B.n77 163.367
R1767 B.n725 B.n82 163.367
R1768 B.n83 B.n82 163.367
R1769 B.n84 B.n83 163.367
R1770 B.n730 B.n84 163.367
R1771 B.n730 B.n89 163.367
R1772 B.n90 B.n89 163.367
R1773 B.n91 B.n90 163.367
R1774 B.n735 B.n91 163.367
R1775 B.n735 B.n96 163.367
R1776 B.n97 B.n96 163.367
R1777 B.n98 B.n97 163.367
R1778 B.n740 B.n98 163.367
R1779 B.n740 B.n103 163.367
R1780 B.n104 B.n103 163.367
R1781 B.n105 B.n104 163.367
R1782 B.n921 B.n919 163.367
R1783 B.n917 B.n109 163.367
R1784 B.n913 B.n911 163.367
R1785 B.n909 B.n111 163.367
R1786 B.n905 B.n903 163.367
R1787 B.n901 B.n113 163.367
R1788 B.n897 B.n895 163.367
R1789 B.n893 B.n115 163.367
R1790 B.n889 B.n887 163.367
R1791 B.n885 B.n117 163.367
R1792 B.n881 B.n879 163.367
R1793 B.n877 B.n119 163.367
R1794 B.n873 B.n871 163.367
R1795 B.n869 B.n121 163.367
R1796 B.n865 B.n863 163.367
R1797 B.n861 B.n123 163.367
R1798 B.n857 B.n855 163.367
R1799 B.n853 B.n125 163.367
R1800 B.n849 B.n847 163.367
R1801 B.n845 B.n127 163.367
R1802 B.n840 B.n838 163.367
R1803 B.n836 B.n131 163.367
R1804 B.n832 B.n830 163.367
R1805 B.n828 B.n133 163.367
R1806 B.n823 B.n821 163.367
R1807 B.n819 B.n137 163.367
R1808 B.n815 B.n813 163.367
R1809 B.n811 B.n139 163.367
R1810 B.n807 B.n805 163.367
R1811 B.n803 B.n141 163.367
R1812 B.n799 B.n797 163.367
R1813 B.n795 B.n143 163.367
R1814 B.n791 B.n789 163.367
R1815 B.n787 B.n145 163.367
R1816 B.n783 B.n781 163.367
R1817 B.n779 B.n147 163.367
R1818 B.n775 B.n773 163.367
R1819 B.n771 B.n149 163.367
R1820 B.n767 B.n765 163.367
R1821 B.n763 B.n151 163.367
R1822 B.n759 B.n757 163.367
R1823 B.n755 B.n153 163.367
R1824 B.n751 B.n749 163.367
R1825 B.n747 B.n155 163.367
R1826 B.n495 B.n266 84.4369
R1827 B.n926 B.n106 84.4369
R1828 B.n489 B.n267 71.676
R1829 B.n487 B.n269 71.676
R1830 B.n483 B.n482 71.676
R1831 B.n476 B.n271 71.676
R1832 B.n475 B.n474 71.676
R1833 B.n468 B.n273 71.676
R1834 B.n467 B.n466 71.676
R1835 B.n460 B.n275 71.676
R1836 B.n459 B.n458 71.676
R1837 B.n452 B.n277 71.676
R1838 B.n451 B.n450 71.676
R1839 B.n444 B.n279 71.676
R1840 B.n443 B.n442 71.676
R1841 B.n436 B.n281 71.676
R1842 B.n435 B.n434 71.676
R1843 B.n428 B.n283 71.676
R1844 B.n427 B.n426 71.676
R1845 B.n420 B.n285 71.676
R1846 B.n419 B.n418 71.676
R1847 B.n411 B.n287 71.676
R1848 B.n410 B.n409 71.676
R1849 B.n403 B.n291 71.676
R1850 B.n402 B.n401 71.676
R1851 B.n395 B.n293 71.676
R1852 B.n394 B.n297 71.676
R1853 B.n390 B.n389 71.676
R1854 B.n383 B.n299 71.676
R1855 B.n382 B.n381 71.676
R1856 B.n375 B.n301 71.676
R1857 B.n374 B.n373 71.676
R1858 B.n367 B.n303 71.676
R1859 B.n366 B.n365 71.676
R1860 B.n359 B.n305 71.676
R1861 B.n358 B.n357 71.676
R1862 B.n351 B.n307 71.676
R1863 B.n350 B.n349 71.676
R1864 B.n343 B.n309 71.676
R1865 B.n342 B.n341 71.676
R1866 B.n335 B.n311 71.676
R1867 B.n334 B.n333 71.676
R1868 B.n327 B.n313 71.676
R1869 B.n326 B.n325 71.676
R1870 B.n319 B.n315 71.676
R1871 B.n318 B.n317 71.676
R1872 B.n920 B.n107 71.676
R1873 B.n919 B.n918 71.676
R1874 B.n912 B.n109 71.676
R1875 B.n911 B.n910 71.676
R1876 B.n904 B.n111 71.676
R1877 B.n903 B.n902 71.676
R1878 B.n896 B.n113 71.676
R1879 B.n895 B.n894 71.676
R1880 B.n888 B.n115 71.676
R1881 B.n887 B.n886 71.676
R1882 B.n880 B.n117 71.676
R1883 B.n879 B.n878 71.676
R1884 B.n872 B.n119 71.676
R1885 B.n871 B.n870 71.676
R1886 B.n864 B.n121 71.676
R1887 B.n863 B.n862 71.676
R1888 B.n856 B.n123 71.676
R1889 B.n855 B.n854 71.676
R1890 B.n848 B.n125 71.676
R1891 B.n847 B.n846 71.676
R1892 B.n839 B.n127 71.676
R1893 B.n838 B.n837 71.676
R1894 B.n831 B.n131 71.676
R1895 B.n830 B.n829 71.676
R1896 B.n822 B.n133 71.676
R1897 B.n821 B.n820 71.676
R1898 B.n814 B.n137 71.676
R1899 B.n813 B.n812 71.676
R1900 B.n806 B.n139 71.676
R1901 B.n805 B.n804 71.676
R1902 B.n798 B.n141 71.676
R1903 B.n797 B.n796 71.676
R1904 B.n790 B.n143 71.676
R1905 B.n789 B.n788 71.676
R1906 B.n782 B.n145 71.676
R1907 B.n781 B.n780 71.676
R1908 B.n774 B.n147 71.676
R1909 B.n773 B.n772 71.676
R1910 B.n766 B.n149 71.676
R1911 B.n765 B.n764 71.676
R1912 B.n758 B.n151 71.676
R1913 B.n757 B.n756 71.676
R1914 B.n750 B.n153 71.676
R1915 B.n749 B.n748 71.676
R1916 B.n748 B.n747 71.676
R1917 B.n751 B.n750 71.676
R1918 B.n756 B.n755 71.676
R1919 B.n759 B.n758 71.676
R1920 B.n764 B.n763 71.676
R1921 B.n767 B.n766 71.676
R1922 B.n772 B.n771 71.676
R1923 B.n775 B.n774 71.676
R1924 B.n780 B.n779 71.676
R1925 B.n783 B.n782 71.676
R1926 B.n788 B.n787 71.676
R1927 B.n791 B.n790 71.676
R1928 B.n796 B.n795 71.676
R1929 B.n799 B.n798 71.676
R1930 B.n804 B.n803 71.676
R1931 B.n807 B.n806 71.676
R1932 B.n812 B.n811 71.676
R1933 B.n815 B.n814 71.676
R1934 B.n820 B.n819 71.676
R1935 B.n823 B.n822 71.676
R1936 B.n829 B.n828 71.676
R1937 B.n832 B.n831 71.676
R1938 B.n837 B.n836 71.676
R1939 B.n840 B.n839 71.676
R1940 B.n846 B.n845 71.676
R1941 B.n849 B.n848 71.676
R1942 B.n854 B.n853 71.676
R1943 B.n857 B.n856 71.676
R1944 B.n862 B.n861 71.676
R1945 B.n865 B.n864 71.676
R1946 B.n870 B.n869 71.676
R1947 B.n873 B.n872 71.676
R1948 B.n878 B.n877 71.676
R1949 B.n881 B.n880 71.676
R1950 B.n886 B.n885 71.676
R1951 B.n889 B.n888 71.676
R1952 B.n894 B.n893 71.676
R1953 B.n897 B.n896 71.676
R1954 B.n902 B.n901 71.676
R1955 B.n905 B.n904 71.676
R1956 B.n910 B.n909 71.676
R1957 B.n913 B.n912 71.676
R1958 B.n918 B.n917 71.676
R1959 B.n921 B.n920 71.676
R1960 B.n490 B.n489 71.676
R1961 B.n484 B.n269 71.676
R1962 B.n482 B.n481 71.676
R1963 B.n477 B.n476 71.676
R1964 B.n474 B.n473 71.676
R1965 B.n469 B.n468 71.676
R1966 B.n466 B.n465 71.676
R1967 B.n461 B.n460 71.676
R1968 B.n458 B.n457 71.676
R1969 B.n453 B.n452 71.676
R1970 B.n450 B.n449 71.676
R1971 B.n445 B.n444 71.676
R1972 B.n442 B.n441 71.676
R1973 B.n437 B.n436 71.676
R1974 B.n434 B.n433 71.676
R1975 B.n429 B.n428 71.676
R1976 B.n426 B.n425 71.676
R1977 B.n421 B.n420 71.676
R1978 B.n418 B.n417 71.676
R1979 B.n412 B.n411 71.676
R1980 B.n409 B.n408 71.676
R1981 B.n404 B.n403 71.676
R1982 B.n401 B.n400 71.676
R1983 B.n396 B.n395 71.676
R1984 B.n391 B.n297 71.676
R1985 B.n389 B.n388 71.676
R1986 B.n384 B.n383 71.676
R1987 B.n381 B.n380 71.676
R1988 B.n376 B.n375 71.676
R1989 B.n373 B.n372 71.676
R1990 B.n368 B.n367 71.676
R1991 B.n365 B.n364 71.676
R1992 B.n360 B.n359 71.676
R1993 B.n357 B.n356 71.676
R1994 B.n352 B.n351 71.676
R1995 B.n349 B.n348 71.676
R1996 B.n344 B.n343 71.676
R1997 B.n341 B.n340 71.676
R1998 B.n336 B.n335 71.676
R1999 B.n333 B.n332 71.676
R2000 B.n328 B.n327 71.676
R2001 B.n325 B.n324 71.676
R2002 B.n320 B.n319 71.676
R2003 B.n317 B.n265 71.676
R2004 B.n296 B.n295 59.5399
R2005 B.n414 B.n289 59.5399
R2006 B.n843 B.n129 59.5399
R2007 B.n825 B.n135 59.5399
R2008 B.n295 B.n294 54.8853
R2009 B.n289 B.n288 54.8853
R2010 B.n129 B.n128 54.8853
R2011 B.n135 B.n134 54.8853
R2012 B.n495 B.n262 45.2105
R2013 B.n501 B.n262 45.2105
R2014 B.n501 B.n258 45.2105
R2015 B.n507 B.n258 45.2105
R2016 B.n507 B.n254 45.2105
R2017 B.n514 B.n254 45.2105
R2018 B.n514 B.n513 45.2105
R2019 B.n520 B.n247 45.2105
R2020 B.n526 B.n247 45.2105
R2021 B.n526 B.n243 45.2105
R2022 B.n532 B.n243 45.2105
R2023 B.n532 B.n239 45.2105
R2024 B.n538 B.n239 45.2105
R2025 B.n538 B.n235 45.2105
R2026 B.n544 B.n235 45.2105
R2027 B.n544 B.n231 45.2105
R2028 B.n550 B.n231 45.2105
R2029 B.n556 B.n227 45.2105
R2030 B.n556 B.n223 45.2105
R2031 B.n562 B.n223 45.2105
R2032 B.n562 B.n219 45.2105
R2033 B.n568 B.n219 45.2105
R2034 B.n568 B.n215 45.2105
R2035 B.n575 B.n215 45.2105
R2036 B.n575 B.n574 45.2105
R2037 B.n581 B.n208 45.2105
R2038 B.n587 B.n208 45.2105
R2039 B.n587 B.n204 45.2105
R2040 B.n593 B.n204 45.2105
R2041 B.n593 B.n200 45.2105
R2042 B.n600 B.n200 45.2105
R2043 B.n600 B.n599 45.2105
R2044 B.n606 B.n193 45.2105
R2045 B.n612 B.n193 45.2105
R2046 B.n612 B.n189 45.2105
R2047 B.n618 B.n189 45.2105
R2048 B.n618 B.n185 45.2105
R2049 B.n625 B.n185 45.2105
R2050 B.n625 B.n624 45.2105
R2051 B.n631 B.n178 45.2105
R2052 B.n637 B.n178 45.2105
R2053 B.n637 B.n174 45.2105
R2054 B.n643 B.n174 45.2105
R2055 B.n643 B.n170 45.2105
R2056 B.n649 B.n170 45.2105
R2057 B.n649 B.n166 45.2105
R2058 B.n655 B.n166 45.2105
R2059 B.n662 B.n162 45.2105
R2060 B.n662 B.n158 45.2105
R2061 B.n668 B.n158 45.2105
R2062 B.n668 B.n4 45.2105
R2063 B.n1040 B.n4 45.2105
R2064 B.n1040 B.n1039 45.2105
R2065 B.n1039 B.n1038 45.2105
R2066 B.n1038 B.n8 45.2105
R2067 B.n1032 B.n8 45.2105
R2068 B.n1032 B.n1031 45.2105
R2069 B.n1030 B.n15 45.2105
R2070 B.n1024 B.n15 45.2105
R2071 B.n1024 B.n1023 45.2105
R2072 B.n1023 B.n1022 45.2105
R2073 B.n1022 B.n22 45.2105
R2074 B.n1016 B.n22 45.2105
R2075 B.n1016 B.n1015 45.2105
R2076 B.n1015 B.n1014 45.2105
R2077 B.n1008 B.n32 45.2105
R2078 B.n1008 B.n1007 45.2105
R2079 B.n1007 B.n1006 45.2105
R2080 B.n1006 B.n36 45.2105
R2081 B.n1000 B.n36 45.2105
R2082 B.n1000 B.n999 45.2105
R2083 B.n999 B.n998 45.2105
R2084 B.n992 B.n46 45.2105
R2085 B.n992 B.n991 45.2105
R2086 B.n991 B.n990 45.2105
R2087 B.n990 B.n50 45.2105
R2088 B.n984 B.n50 45.2105
R2089 B.n984 B.n983 45.2105
R2090 B.n983 B.n982 45.2105
R2091 B.n976 B.n60 45.2105
R2092 B.n976 B.n975 45.2105
R2093 B.n975 B.n974 45.2105
R2094 B.n974 B.n64 45.2105
R2095 B.n968 B.n64 45.2105
R2096 B.n968 B.n967 45.2105
R2097 B.n967 B.n966 45.2105
R2098 B.n966 B.n71 45.2105
R2099 B.n960 B.n959 45.2105
R2100 B.n959 B.n958 45.2105
R2101 B.n958 B.n78 45.2105
R2102 B.n952 B.n78 45.2105
R2103 B.n952 B.n951 45.2105
R2104 B.n951 B.n950 45.2105
R2105 B.n950 B.n85 45.2105
R2106 B.n944 B.n85 45.2105
R2107 B.n944 B.n943 45.2105
R2108 B.n943 B.n942 45.2105
R2109 B.n936 B.n95 45.2105
R2110 B.n936 B.n935 45.2105
R2111 B.n935 B.n934 45.2105
R2112 B.n934 B.n99 45.2105
R2113 B.n928 B.n99 45.2105
R2114 B.n928 B.n927 45.2105
R2115 B.n927 B.n926 45.2105
R2116 B.n550 B.t3 42.5511
R2117 B.n960 B.t7 42.5511
R2118 B.n624 B.t2 41.2214
R2119 B.n32 B.t1 41.2214
R2120 B.t6 B.n162 34.5729
R2121 B.n1031 B.t0 34.5729
R2122 B.n581 B.t4 33.2432
R2123 B.n982 B.t8 33.2432
R2124 B.n745 B.n744 30.4395
R2125 B.n924 B.n923 30.4395
R2126 B.n497 B.n264 30.4395
R2127 B.n493 B.n492 30.4395
R2128 B.n520 B.t18 26.5946
R2129 B.n599 B.t5 26.5946
R2130 B.n46 B.t9 26.5946
R2131 B.n942 B.t11 26.5946
R2132 B.n513 B.t18 18.6164
R2133 B.n606 B.t5 18.6164
R2134 B.n998 B.t9 18.6164
R2135 B.n95 B.t11 18.6164
R2136 B B.n1042 18.0485
R2137 B.n574 B.t4 11.9679
R2138 B.n60 B.t8 11.9679
R2139 B.n655 B.t6 10.6382
R2140 B.t0 B.n1030 10.6382
R2141 B.n923 B.n922 10.6151
R2142 B.n922 B.n108 10.6151
R2143 B.n916 B.n108 10.6151
R2144 B.n916 B.n915 10.6151
R2145 B.n915 B.n914 10.6151
R2146 B.n914 B.n110 10.6151
R2147 B.n908 B.n110 10.6151
R2148 B.n908 B.n907 10.6151
R2149 B.n907 B.n906 10.6151
R2150 B.n906 B.n112 10.6151
R2151 B.n900 B.n112 10.6151
R2152 B.n900 B.n899 10.6151
R2153 B.n899 B.n898 10.6151
R2154 B.n898 B.n114 10.6151
R2155 B.n892 B.n114 10.6151
R2156 B.n892 B.n891 10.6151
R2157 B.n891 B.n890 10.6151
R2158 B.n890 B.n116 10.6151
R2159 B.n884 B.n116 10.6151
R2160 B.n884 B.n883 10.6151
R2161 B.n883 B.n882 10.6151
R2162 B.n882 B.n118 10.6151
R2163 B.n876 B.n118 10.6151
R2164 B.n876 B.n875 10.6151
R2165 B.n875 B.n874 10.6151
R2166 B.n874 B.n120 10.6151
R2167 B.n868 B.n120 10.6151
R2168 B.n868 B.n867 10.6151
R2169 B.n867 B.n866 10.6151
R2170 B.n866 B.n122 10.6151
R2171 B.n860 B.n122 10.6151
R2172 B.n860 B.n859 10.6151
R2173 B.n859 B.n858 10.6151
R2174 B.n858 B.n124 10.6151
R2175 B.n852 B.n124 10.6151
R2176 B.n852 B.n851 10.6151
R2177 B.n851 B.n850 10.6151
R2178 B.n850 B.n126 10.6151
R2179 B.n844 B.n126 10.6151
R2180 B.n842 B.n841 10.6151
R2181 B.n841 B.n130 10.6151
R2182 B.n835 B.n130 10.6151
R2183 B.n835 B.n834 10.6151
R2184 B.n834 B.n833 10.6151
R2185 B.n833 B.n132 10.6151
R2186 B.n827 B.n132 10.6151
R2187 B.n827 B.n826 10.6151
R2188 B.n824 B.n136 10.6151
R2189 B.n818 B.n136 10.6151
R2190 B.n818 B.n817 10.6151
R2191 B.n817 B.n816 10.6151
R2192 B.n816 B.n138 10.6151
R2193 B.n810 B.n138 10.6151
R2194 B.n810 B.n809 10.6151
R2195 B.n809 B.n808 10.6151
R2196 B.n808 B.n140 10.6151
R2197 B.n802 B.n140 10.6151
R2198 B.n802 B.n801 10.6151
R2199 B.n801 B.n800 10.6151
R2200 B.n800 B.n142 10.6151
R2201 B.n794 B.n142 10.6151
R2202 B.n794 B.n793 10.6151
R2203 B.n793 B.n792 10.6151
R2204 B.n792 B.n144 10.6151
R2205 B.n786 B.n144 10.6151
R2206 B.n786 B.n785 10.6151
R2207 B.n785 B.n784 10.6151
R2208 B.n784 B.n146 10.6151
R2209 B.n778 B.n146 10.6151
R2210 B.n778 B.n777 10.6151
R2211 B.n777 B.n776 10.6151
R2212 B.n776 B.n148 10.6151
R2213 B.n770 B.n148 10.6151
R2214 B.n770 B.n769 10.6151
R2215 B.n769 B.n768 10.6151
R2216 B.n768 B.n150 10.6151
R2217 B.n762 B.n150 10.6151
R2218 B.n762 B.n761 10.6151
R2219 B.n761 B.n760 10.6151
R2220 B.n760 B.n152 10.6151
R2221 B.n754 B.n152 10.6151
R2222 B.n754 B.n753 10.6151
R2223 B.n753 B.n752 10.6151
R2224 B.n752 B.n154 10.6151
R2225 B.n746 B.n154 10.6151
R2226 B.n746 B.n745 10.6151
R2227 B.n498 B.n497 10.6151
R2228 B.n499 B.n498 10.6151
R2229 B.n499 B.n256 10.6151
R2230 B.n509 B.n256 10.6151
R2231 B.n510 B.n509 10.6151
R2232 B.n511 B.n510 10.6151
R2233 B.n511 B.n249 10.6151
R2234 B.n522 B.n249 10.6151
R2235 B.n523 B.n522 10.6151
R2236 B.n524 B.n523 10.6151
R2237 B.n524 B.n241 10.6151
R2238 B.n534 B.n241 10.6151
R2239 B.n535 B.n534 10.6151
R2240 B.n536 B.n535 10.6151
R2241 B.n536 B.n233 10.6151
R2242 B.n546 B.n233 10.6151
R2243 B.n547 B.n546 10.6151
R2244 B.n548 B.n547 10.6151
R2245 B.n548 B.n225 10.6151
R2246 B.n558 B.n225 10.6151
R2247 B.n559 B.n558 10.6151
R2248 B.n560 B.n559 10.6151
R2249 B.n560 B.n217 10.6151
R2250 B.n570 B.n217 10.6151
R2251 B.n571 B.n570 10.6151
R2252 B.n572 B.n571 10.6151
R2253 B.n572 B.n210 10.6151
R2254 B.n583 B.n210 10.6151
R2255 B.n584 B.n583 10.6151
R2256 B.n585 B.n584 10.6151
R2257 B.n585 B.n202 10.6151
R2258 B.n595 B.n202 10.6151
R2259 B.n596 B.n595 10.6151
R2260 B.n597 B.n596 10.6151
R2261 B.n597 B.n195 10.6151
R2262 B.n608 B.n195 10.6151
R2263 B.n609 B.n608 10.6151
R2264 B.n610 B.n609 10.6151
R2265 B.n610 B.n187 10.6151
R2266 B.n620 B.n187 10.6151
R2267 B.n621 B.n620 10.6151
R2268 B.n622 B.n621 10.6151
R2269 B.n622 B.n180 10.6151
R2270 B.n633 B.n180 10.6151
R2271 B.n634 B.n633 10.6151
R2272 B.n635 B.n634 10.6151
R2273 B.n635 B.n172 10.6151
R2274 B.n645 B.n172 10.6151
R2275 B.n646 B.n645 10.6151
R2276 B.n647 B.n646 10.6151
R2277 B.n647 B.n164 10.6151
R2278 B.n657 B.n164 10.6151
R2279 B.n658 B.n657 10.6151
R2280 B.n660 B.n658 10.6151
R2281 B.n660 B.n659 10.6151
R2282 B.n659 B.n156 10.6151
R2283 B.n671 B.n156 10.6151
R2284 B.n672 B.n671 10.6151
R2285 B.n673 B.n672 10.6151
R2286 B.n674 B.n673 10.6151
R2287 B.n676 B.n674 10.6151
R2288 B.n677 B.n676 10.6151
R2289 B.n678 B.n677 10.6151
R2290 B.n679 B.n678 10.6151
R2291 B.n681 B.n679 10.6151
R2292 B.n682 B.n681 10.6151
R2293 B.n683 B.n682 10.6151
R2294 B.n684 B.n683 10.6151
R2295 B.n686 B.n684 10.6151
R2296 B.n687 B.n686 10.6151
R2297 B.n688 B.n687 10.6151
R2298 B.n689 B.n688 10.6151
R2299 B.n691 B.n689 10.6151
R2300 B.n692 B.n691 10.6151
R2301 B.n693 B.n692 10.6151
R2302 B.n694 B.n693 10.6151
R2303 B.n696 B.n694 10.6151
R2304 B.n697 B.n696 10.6151
R2305 B.n698 B.n697 10.6151
R2306 B.n699 B.n698 10.6151
R2307 B.n701 B.n699 10.6151
R2308 B.n702 B.n701 10.6151
R2309 B.n703 B.n702 10.6151
R2310 B.n704 B.n703 10.6151
R2311 B.n706 B.n704 10.6151
R2312 B.n707 B.n706 10.6151
R2313 B.n708 B.n707 10.6151
R2314 B.n709 B.n708 10.6151
R2315 B.n711 B.n709 10.6151
R2316 B.n712 B.n711 10.6151
R2317 B.n713 B.n712 10.6151
R2318 B.n714 B.n713 10.6151
R2319 B.n716 B.n714 10.6151
R2320 B.n717 B.n716 10.6151
R2321 B.n718 B.n717 10.6151
R2322 B.n719 B.n718 10.6151
R2323 B.n721 B.n719 10.6151
R2324 B.n722 B.n721 10.6151
R2325 B.n723 B.n722 10.6151
R2326 B.n724 B.n723 10.6151
R2327 B.n726 B.n724 10.6151
R2328 B.n727 B.n726 10.6151
R2329 B.n728 B.n727 10.6151
R2330 B.n729 B.n728 10.6151
R2331 B.n731 B.n729 10.6151
R2332 B.n732 B.n731 10.6151
R2333 B.n733 B.n732 10.6151
R2334 B.n734 B.n733 10.6151
R2335 B.n736 B.n734 10.6151
R2336 B.n737 B.n736 10.6151
R2337 B.n738 B.n737 10.6151
R2338 B.n739 B.n738 10.6151
R2339 B.n741 B.n739 10.6151
R2340 B.n742 B.n741 10.6151
R2341 B.n743 B.n742 10.6151
R2342 B.n744 B.n743 10.6151
R2343 B.n492 B.n491 10.6151
R2344 B.n491 B.n268 10.6151
R2345 B.n486 B.n268 10.6151
R2346 B.n486 B.n485 10.6151
R2347 B.n485 B.n270 10.6151
R2348 B.n480 B.n270 10.6151
R2349 B.n480 B.n479 10.6151
R2350 B.n479 B.n478 10.6151
R2351 B.n478 B.n272 10.6151
R2352 B.n472 B.n272 10.6151
R2353 B.n472 B.n471 10.6151
R2354 B.n471 B.n470 10.6151
R2355 B.n470 B.n274 10.6151
R2356 B.n464 B.n274 10.6151
R2357 B.n464 B.n463 10.6151
R2358 B.n463 B.n462 10.6151
R2359 B.n462 B.n276 10.6151
R2360 B.n456 B.n276 10.6151
R2361 B.n456 B.n455 10.6151
R2362 B.n455 B.n454 10.6151
R2363 B.n454 B.n278 10.6151
R2364 B.n448 B.n278 10.6151
R2365 B.n448 B.n447 10.6151
R2366 B.n447 B.n446 10.6151
R2367 B.n446 B.n280 10.6151
R2368 B.n440 B.n280 10.6151
R2369 B.n440 B.n439 10.6151
R2370 B.n439 B.n438 10.6151
R2371 B.n438 B.n282 10.6151
R2372 B.n432 B.n282 10.6151
R2373 B.n432 B.n431 10.6151
R2374 B.n431 B.n430 10.6151
R2375 B.n430 B.n284 10.6151
R2376 B.n424 B.n284 10.6151
R2377 B.n424 B.n423 10.6151
R2378 B.n423 B.n422 10.6151
R2379 B.n422 B.n286 10.6151
R2380 B.n416 B.n286 10.6151
R2381 B.n416 B.n415 10.6151
R2382 B.n413 B.n290 10.6151
R2383 B.n407 B.n290 10.6151
R2384 B.n407 B.n406 10.6151
R2385 B.n406 B.n405 10.6151
R2386 B.n405 B.n292 10.6151
R2387 B.n399 B.n292 10.6151
R2388 B.n399 B.n398 10.6151
R2389 B.n398 B.n397 10.6151
R2390 B.n393 B.n392 10.6151
R2391 B.n392 B.n298 10.6151
R2392 B.n387 B.n298 10.6151
R2393 B.n387 B.n386 10.6151
R2394 B.n386 B.n385 10.6151
R2395 B.n385 B.n300 10.6151
R2396 B.n379 B.n300 10.6151
R2397 B.n379 B.n378 10.6151
R2398 B.n378 B.n377 10.6151
R2399 B.n377 B.n302 10.6151
R2400 B.n371 B.n302 10.6151
R2401 B.n371 B.n370 10.6151
R2402 B.n370 B.n369 10.6151
R2403 B.n369 B.n304 10.6151
R2404 B.n363 B.n304 10.6151
R2405 B.n363 B.n362 10.6151
R2406 B.n362 B.n361 10.6151
R2407 B.n361 B.n306 10.6151
R2408 B.n355 B.n306 10.6151
R2409 B.n355 B.n354 10.6151
R2410 B.n354 B.n353 10.6151
R2411 B.n353 B.n308 10.6151
R2412 B.n347 B.n308 10.6151
R2413 B.n347 B.n346 10.6151
R2414 B.n346 B.n345 10.6151
R2415 B.n345 B.n310 10.6151
R2416 B.n339 B.n310 10.6151
R2417 B.n339 B.n338 10.6151
R2418 B.n338 B.n337 10.6151
R2419 B.n337 B.n312 10.6151
R2420 B.n331 B.n312 10.6151
R2421 B.n331 B.n330 10.6151
R2422 B.n330 B.n329 10.6151
R2423 B.n329 B.n314 10.6151
R2424 B.n323 B.n314 10.6151
R2425 B.n323 B.n322 10.6151
R2426 B.n322 B.n321 10.6151
R2427 B.n321 B.n316 10.6151
R2428 B.n316 B.n264 10.6151
R2429 B.n493 B.n260 10.6151
R2430 B.n503 B.n260 10.6151
R2431 B.n504 B.n503 10.6151
R2432 B.n505 B.n504 10.6151
R2433 B.n505 B.n252 10.6151
R2434 B.n516 B.n252 10.6151
R2435 B.n517 B.n516 10.6151
R2436 B.n518 B.n517 10.6151
R2437 B.n518 B.n245 10.6151
R2438 B.n528 B.n245 10.6151
R2439 B.n529 B.n528 10.6151
R2440 B.n530 B.n529 10.6151
R2441 B.n530 B.n237 10.6151
R2442 B.n540 B.n237 10.6151
R2443 B.n541 B.n540 10.6151
R2444 B.n542 B.n541 10.6151
R2445 B.n542 B.n229 10.6151
R2446 B.n552 B.n229 10.6151
R2447 B.n553 B.n552 10.6151
R2448 B.n554 B.n553 10.6151
R2449 B.n554 B.n221 10.6151
R2450 B.n564 B.n221 10.6151
R2451 B.n565 B.n564 10.6151
R2452 B.n566 B.n565 10.6151
R2453 B.n566 B.n213 10.6151
R2454 B.n577 B.n213 10.6151
R2455 B.n578 B.n577 10.6151
R2456 B.n579 B.n578 10.6151
R2457 B.n579 B.n206 10.6151
R2458 B.n589 B.n206 10.6151
R2459 B.n590 B.n589 10.6151
R2460 B.n591 B.n590 10.6151
R2461 B.n591 B.n198 10.6151
R2462 B.n602 B.n198 10.6151
R2463 B.n603 B.n602 10.6151
R2464 B.n604 B.n603 10.6151
R2465 B.n604 B.n191 10.6151
R2466 B.n614 B.n191 10.6151
R2467 B.n615 B.n614 10.6151
R2468 B.n616 B.n615 10.6151
R2469 B.n616 B.n183 10.6151
R2470 B.n627 B.n183 10.6151
R2471 B.n628 B.n627 10.6151
R2472 B.n629 B.n628 10.6151
R2473 B.n629 B.n176 10.6151
R2474 B.n639 B.n176 10.6151
R2475 B.n640 B.n639 10.6151
R2476 B.n641 B.n640 10.6151
R2477 B.n641 B.n168 10.6151
R2478 B.n651 B.n168 10.6151
R2479 B.n652 B.n651 10.6151
R2480 B.n653 B.n652 10.6151
R2481 B.n653 B.n160 10.6151
R2482 B.n664 B.n160 10.6151
R2483 B.n665 B.n664 10.6151
R2484 B.n666 B.n665 10.6151
R2485 B.n666 B.n0 10.6151
R2486 B.n1036 B.n1 10.6151
R2487 B.n1036 B.n1035 10.6151
R2488 B.n1035 B.n1034 10.6151
R2489 B.n1034 B.n10 10.6151
R2490 B.n1028 B.n10 10.6151
R2491 B.n1028 B.n1027 10.6151
R2492 B.n1027 B.n1026 10.6151
R2493 B.n1026 B.n17 10.6151
R2494 B.n1020 B.n17 10.6151
R2495 B.n1020 B.n1019 10.6151
R2496 B.n1019 B.n1018 10.6151
R2497 B.n1018 B.n24 10.6151
R2498 B.n1012 B.n24 10.6151
R2499 B.n1012 B.n1011 10.6151
R2500 B.n1011 B.n1010 10.6151
R2501 B.n1010 B.n30 10.6151
R2502 B.n1004 B.n30 10.6151
R2503 B.n1004 B.n1003 10.6151
R2504 B.n1003 B.n1002 10.6151
R2505 B.n1002 B.n38 10.6151
R2506 B.n996 B.n38 10.6151
R2507 B.n996 B.n995 10.6151
R2508 B.n995 B.n994 10.6151
R2509 B.n994 B.n44 10.6151
R2510 B.n988 B.n44 10.6151
R2511 B.n988 B.n987 10.6151
R2512 B.n987 B.n986 10.6151
R2513 B.n986 B.n52 10.6151
R2514 B.n980 B.n52 10.6151
R2515 B.n980 B.n979 10.6151
R2516 B.n979 B.n978 10.6151
R2517 B.n978 B.n58 10.6151
R2518 B.n972 B.n58 10.6151
R2519 B.n972 B.n971 10.6151
R2520 B.n971 B.n970 10.6151
R2521 B.n970 B.n66 10.6151
R2522 B.n964 B.n66 10.6151
R2523 B.n964 B.n963 10.6151
R2524 B.n963 B.n962 10.6151
R2525 B.n962 B.n73 10.6151
R2526 B.n956 B.n73 10.6151
R2527 B.n956 B.n955 10.6151
R2528 B.n955 B.n954 10.6151
R2529 B.n954 B.n80 10.6151
R2530 B.n948 B.n80 10.6151
R2531 B.n948 B.n947 10.6151
R2532 B.n947 B.n946 10.6151
R2533 B.n946 B.n87 10.6151
R2534 B.n940 B.n87 10.6151
R2535 B.n940 B.n939 10.6151
R2536 B.n939 B.n938 10.6151
R2537 B.n938 B.n93 10.6151
R2538 B.n932 B.n93 10.6151
R2539 B.n932 B.n931 10.6151
R2540 B.n931 B.n930 10.6151
R2541 B.n930 B.n101 10.6151
R2542 B.n924 B.n101 10.6151
R2543 B.n843 B.n842 6.5566
R2544 B.n826 B.n825 6.5566
R2545 B.n414 B.n413 6.5566
R2546 B.n397 B.n296 6.5566
R2547 B.n844 B.n843 4.05904
R2548 B.n825 B.n824 4.05904
R2549 B.n415 B.n414 4.05904
R2550 B.n393 B.n296 4.05904
R2551 B.n631 B.t2 3.98962
R2552 B.n1014 B.t1 3.98962
R2553 B.n1042 B.n0 2.81026
R2554 B.n1042 B.n1 2.81026
R2555 B.t3 B.n227 2.65991
R2556 B.t7 B.n71 2.65991
R2557 VN.n75 VN.n39 161.3
R2558 VN.n74 VN.n73 161.3
R2559 VN.n72 VN.n40 161.3
R2560 VN.n71 VN.n70 161.3
R2561 VN.n69 VN.n41 161.3
R2562 VN.n68 VN.n67 161.3
R2563 VN.n66 VN.n65 161.3
R2564 VN.n64 VN.n43 161.3
R2565 VN.n63 VN.n62 161.3
R2566 VN.n61 VN.n44 161.3
R2567 VN.n60 VN.n59 161.3
R2568 VN.n58 VN.n45 161.3
R2569 VN.n57 VN.n56 161.3
R2570 VN.n55 VN.n46 161.3
R2571 VN.n54 VN.n53 161.3
R2572 VN.n52 VN.n47 161.3
R2573 VN.n51 VN.n50 161.3
R2574 VN.n36 VN.n0 161.3
R2575 VN.n35 VN.n34 161.3
R2576 VN.n33 VN.n1 161.3
R2577 VN.n32 VN.n31 161.3
R2578 VN.n30 VN.n2 161.3
R2579 VN.n29 VN.n28 161.3
R2580 VN.n27 VN.n26 161.3
R2581 VN.n25 VN.n4 161.3
R2582 VN.n24 VN.n23 161.3
R2583 VN.n22 VN.n5 161.3
R2584 VN.n21 VN.n20 161.3
R2585 VN.n19 VN.n6 161.3
R2586 VN.n18 VN.n17 161.3
R2587 VN.n16 VN.n7 161.3
R2588 VN.n15 VN.n14 161.3
R2589 VN.n13 VN.n8 161.3
R2590 VN.n12 VN.n11 161.3
R2591 VN.n10 VN.t1 141.612
R2592 VN.n49 VN.t5 141.612
R2593 VN.n19 VN.t8 108.644
R2594 VN.n9 VN.t7 108.644
R2595 VN.n3 VN.t4 108.644
R2596 VN.n37 VN.t6 108.644
R2597 VN.n58 VN.t0 108.644
R2598 VN.n48 VN.t9 108.644
R2599 VN.n42 VN.t2 108.644
R2600 VN.n76 VN.t3 108.644
R2601 VN.n38 VN.n37 102.927
R2602 VN.n77 VN.n76 102.927
R2603 VN.n31 VN.n1 56.5193
R2604 VN.n70 VN.n40 56.5193
R2605 VN.n10 VN.n9 56.1683
R2606 VN.n49 VN.n48 56.1683
R2607 VN VN.n77 52.2595
R2608 VN.n14 VN.n7 48.7492
R2609 VN.n24 VN.n5 48.7492
R2610 VN.n53 VN.n46 48.7492
R2611 VN.n63 VN.n44 48.7492
R2612 VN.n14 VN.n13 32.2376
R2613 VN.n25 VN.n24 32.2376
R2614 VN.n53 VN.n52 32.2376
R2615 VN.n64 VN.n63 32.2376
R2616 VN.n13 VN.n12 24.4675
R2617 VN.n18 VN.n7 24.4675
R2618 VN.n19 VN.n18 24.4675
R2619 VN.n20 VN.n19 24.4675
R2620 VN.n20 VN.n5 24.4675
R2621 VN.n26 VN.n25 24.4675
R2622 VN.n30 VN.n29 24.4675
R2623 VN.n31 VN.n30 24.4675
R2624 VN.n35 VN.n1 24.4675
R2625 VN.n36 VN.n35 24.4675
R2626 VN.n52 VN.n51 24.4675
R2627 VN.n59 VN.n44 24.4675
R2628 VN.n59 VN.n58 24.4675
R2629 VN.n58 VN.n57 24.4675
R2630 VN.n57 VN.n46 24.4675
R2631 VN.n70 VN.n69 24.4675
R2632 VN.n69 VN.n68 24.4675
R2633 VN.n65 VN.n64 24.4675
R2634 VN.n75 VN.n74 24.4675
R2635 VN.n74 VN.n40 24.4675
R2636 VN.n12 VN.n9 16.1487
R2637 VN.n26 VN.n3 16.1487
R2638 VN.n51 VN.n48 16.1487
R2639 VN.n65 VN.n42 16.1487
R2640 VN.n29 VN.n3 8.31928
R2641 VN.n68 VN.n42 8.31928
R2642 VN.n37 VN.n36 7.82994
R2643 VN.n76 VN.n75 7.82994
R2644 VN.n50 VN.n49 6.98649
R2645 VN.n11 VN.n10 6.98649
R2646 VN.n77 VN.n39 0.278367
R2647 VN.n38 VN.n0 0.278367
R2648 VN.n73 VN.n39 0.189894
R2649 VN.n73 VN.n72 0.189894
R2650 VN.n72 VN.n71 0.189894
R2651 VN.n71 VN.n41 0.189894
R2652 VN.n67 VN.n41 0.189894
R2653 VN.n67 VN.n66 0.189894
R2654 VN.n66 VN.n43 0.189894
R2655 VN.n62 VN.n43 0.189894
R2656 VN.n62 VN.n61 0.189894
R2657 VN.n61 VN.n60 0.189894
R2658 VN.n60 VN.n45 0.189894
R2659 VN.n56 VN.n45 0.189894
R2660 VN.n56 VN.n55 0.189894
R2661 VN.n55 VN.n54 0.189894
R2662 VN.n54 VN.n47 0.189894
R2663 VN.n50 VN.n47 0.189894
R2664 VN.n11 VN.n8 0.189894
R2665 VN.n15 VN.n8 0.189894
R2666 VN.n16 VN.n15 0.189894
R2667 VN.n17 VN.n16 0.189894
R2668 VN.n17 VN.n6 0.189894
R2669 VN.n21 VN.n6 0.189894
R2670 VN.n22 VN.n21 0.189894
R2671 VN.n23 VN.n22 0.189894
R2672 VN.n23 VN.n4 0.189894
R2673 VN.n27 VN.n4 0.189894
R2674 VN.n28 VN.n27 0.189894
R2675 VN.n28 VN.n2 0.189894
R2676 VN.n32 VN.n2 0.189894
R2677 VN.n33 VN.n32 0.189894
R2678 VN.n34 VN.n33 0.189894
R2679 VN.n34 VN.n0 0.189894
R2680 VN VN.n38 0.153454
R2681 VDD2.n125 VDD2.n124 289.615
R2682 VDD2.n60 VDD2.n59 289.615
R2683 VDD2.n124 VDD2.n123 185
R2684 VDD2.n67 VDD2.n66 185
R2685 VDD2.n118 VDD2.n117 185
R2686 VDD2.n116 VDD2.n115 185
R2687 VDD2.n71 VDD2.n70 185
R2688 VDD2.n110 VDD2.n109 185
R2689 VDD2.n108 VDD2.n107 185
R2690 VDD2.n75 VDD2.n74 185
R2691 VDD2.n102 VDD2.n101 185
R2692 VDD2.n100 VDD2.n99 185
R2693 VDD2.n79 VDD2.n78 185
R2694 VDD2.n94 VDD2.n93 185
R2695 VDD2.n92 VDD2.n91 185
R2696 VDD2.n83 VDD2.n82 185
R2697 VDD2.n86 VDD2.n85 185
R2698 VDD2.n21 VDD2.n20 185
R2699 VDD2.n18 VDD2.n17 185
R2700 VDD2.n27 VDD2.n26 185
R2701 VDD2.n29 VDD2.n28 185
R2702 VDD2.n14 VDD2.n13 185
R2703 VDD2.n35 VDD2.n34 185
R2704 VDD2.n37 VDD2.n36 185
R2705 VDD2.n10 VDD2.n9 185
R2706 VDD2.n43 VDD2.n42 185
R2707 VDD2.n45 VDD2.n44 185
R2708 VDD2.n6 VDD2.n5 185
R2709 VDD2.n51 VDD2.n50 185
R2710 VDD2.n53 VDD2.n52 185
R2711 VDD2.n2 VDD2.n1 185
R2712 VDD2.n59 VDD2.n58 185
R2713 VDD2.t8 VDD2.n19 147.659
R2714 VDD2.t6 VDD2.n84 147.659
R2715 VDD2.n124 VDD2.n66 104.615
R2716 VDD2.n117 VDD2.n66 104.615
R2717 VDD2.n117 VDD2.n116 104.615
R2718 VDD2.n116 VDD2.n70 104.615
R2719 VDD2.n109 VDD2.n70 104.615
R2720 VDD2.n109 VDD2.n108 104.615
R2721 VDD2.n108 VDD2.n74 104.615
R2722 VDD2.n101 VDD2.n74 104.615
R2723 VDD2.n101 VDD2.n100 104.615
R2724 VDD2.n100 VDD2.n78 104.615
R2725 VDD2.n93 VDD2.n78 104.615
R2726 VDD2.n93 VDD2.n92 104.615
R2727 VDD2.n92 VDD2.n82 104.615
R2728 VDD2.n85 VDD2.n82 104.615
R2729 VDD2.n20 VDD2.n17 104.615
R2730 VDD2.n27 VDD2.n17 104.615
R2731 VDD2.n28 VDD2.n27 104.615
R2732 VDD2.n28 VDD2.n13 104.615
R2733 VDD2.n35 VDD2.n13 104.615
R2734 VDD2.n36 VDD2.n35 104.615
R2735 VDD2.n36 VDD2.n9 104.615
R2736 VDD2.n43 VDD2.n9 104.615
R2737 VDD2.n44 VDD2.n43 104.615
R2738 VDD2.n44 VDD2.n5 104.615
R2739 VDD2.n51 VDD2.n5 104.615
R2740 VDD2.n52 VDD2.n51 104.615
R2741 VDD2.n52 VDD2.n1 104.615
R2742 VDD2.n59 VDD2.n1 104.615
R2743 VDD2.n64 VDD2.n63 67.6194
R2744 VDD2 VDD2.n129 67.6157
R2745 VDD2.n128 VDD2.n127 65.8451
R2746 VDD2.n62 VDD2.n61 65.845
R2747 VDD2.n62 VDD2.n60 53.825
R2748 VDD2.n85 VDD2.t6 52.3082
R2749 VDD2.n20 VDD2.t8 52.3082
R2750 VDD2.n126 VDD2.n125 51.3853
R2751 VDD2.n126 VDD2.n64 45.0192
R2752 VDD2.n86 VDD2.n84 15.6677
R2753 VDD2.n21 VDD2.n19 15.6677
R2754 VDD2.n87 VDD2.n83 12.8005
R2755 VDD2.n22 VDD2.n18 12.8005
R2756 VDD2.n91 VDD2.n90 12.0247
R2757 VDD2.n26 VDD2.n25 12.0247
R2758 VDD2.n123 VDD2.n65 11.249
R2759 VDD2.n94 VDD2.n81 11.249
R2760 VDD2.n29 VDD2.n16 11.249
R2761 VDD2.n58 VDD2.n0 11.249
R2762 VDD2.n122 VDD2.n67 10.4732
R2763 VDD2.n95 VDD2.n79 10.4732
R2764 VDD2.n30 VDD2.n14 10.4732
R2765 VDD2.n57 VDD2.n2 10.4732
R2766 VDD2.n119 VDD2.n118 9.69747
R2767 VDD2.n99 VDD2.n98 9.69747
R2768 VDD2.n34 VDD2.n33 9.69747
R2769 VDD2.n54 VDD2.n53 9.69747
R2770 VDD2.n121 VDD2.n65 9.45567
R2771 VDD2.n56 VDD2.n0 9.45567
R2772 VDD2.n112 VDD2.n111 9.3005
R2773 VDD2.n114 VDD2.n113 9.3005
R2774 VDD2.n69 VDD2.n68 9.3005
R2775 VDD2.n120 VDD2.n119 9.3005
R2776 VDD2.n122 VDD2.n121 9.3005
R2777 VDD2.n73 VDD2.n72 9.3005
R2778 VDD2.n106 VDD2.n105 9.3005
R2779 VDD2.n104 VDD2.n103 9.3005
R2780 VDD2.n77 VDD2.n76 9.3005
R2781 VDD2.n98 VDD2.n97 9.3005
R2782 VDD2.n96 VDD2.n95 9.3005
R2783 VDD2.n81 VDD2.n80 9.3005
R2784 VDD2.n90 VDD2.n89 9.3005
R2785 VDD2.n88 VDD2.n87 9.3005
R2786 VDD2.n8 VDD2.n7 9.3005
R2787 VDD2.n47 VDD2.n46 9.3005
R2788 VDD2.n49 VDD2.n48 9.3005
R2789 VDD2.n4 VDD2.n3 9.3005
R2790 VDD2.n55 VDD2.n54 9.3005
R2791 VDD2.n57 VDD2.n56 9.3005
R2792 VDD2.n39 VDD2.n38 9.3005
R2793 VDD2.n12 VDD2.n11 9.3005
R2794 VDD2.n33 VDD2.n32 9.3005
R2795 VDD2.n31 VDD2.n30 9.3005
R2796 VDD2.n16 VDD2.n15 9.3005
R2797 VDD2.n25 VDD2.n24 9.3005
R2798 VDD2.n23 VDD2.n22 9.3005
R2799 VDD2.n41 VDD2.n40 9.3005
R2800 VDD2.n115 VDD2.n69 8.92171
R2801 VDD2.n102 VDD2.n77 8.92171
R2802 VDD2.n37 VDD2.n12 8.92171
R2803 VDD2.n50 VDD2.n4 8.92171
R2804 VDD2.n114 VDD2.n71 8.14595
R2805 VDD2.n103 VDD2.n75 8.14595
R2806 VDD2.n38 VDD2.n10 8.14595
R2807 VDD2.n49 VDD2.n6 8.14595
R2808 VDD2.n111 VDD2.n110 7.3702
R2809 VDD2.n107 VDD2.n106 7.3702
R2810 VDD2.n42 VDD2.n41 7.3702
R2811 VDD2.n46 VDD2.n45 7.3702
R2812 VDD2.n110 VDD2.n73 6.59444
R2813 VDD2.n107 VDD2.n73 6.59444
R2814 VDD2.n42 VDD2.n8 6.59444
R2815 VDD2.n45 VDD2.n8 6.59444
R2816 VDD2.n111 VDD2.n71 5.81868
R2817 VDD2.n106 VDD2.n75 5.81868
R2818 VDD2.n41 VDD2.n10 5.81868
R2819 VDD2.n46 VDD2.n6 5.81868
R2820 VDD2.n115 VDD2.n114 5.04292
R2821 VDD2.n103 VDD2.n102 5.04292
R2822 VDD2.n38 VDD2.n37 5.04292
R2823 VDD2.n50 VDD2.n49 5.04292
R2824 VDD2.n23 VDD2.n19 4.38563
R2825 VDD2.n88 VDD2.n84 4.38563
R2826 VDD2.n118 VDD2.n69 4.26717
R2827 VDD2.n99 VDD2.n77 4.26717
R2828 VDD2.n34 VDD2.n12 4.26717
R2829 VDD2.n53 VDD2.n4 4.26717
R2830 VDD2.n119 VDD2.n67 3.49141
R2831 VDD2.n98 VDD2.n79 3.49141
R2832 VDD2.n33 VDD2.n14 3.49141
R2833 VDD2.n54 VDD2.n2 3.49141
R2834 VDD2.n123 VDD2.n122 2.71565
R2835 VDD2.n95 VDD2.n94 2.71565
R2836 VDD2.n30 VDD2.n29 2.71565
R2837 VDD2.n58 VDD2.n57 2.71565
R2838 VDD2.n128 VDD2.n126 2.44016
R2839 VDD2.n125 VDD2.n65 1.93989
R2840 VDD2.n91 VDD2.n81 1.93989
R2841 VDD2.n26 VDD2.n16 1.93989
R2842 VDD2.n60 VDD2.n0 1.93989
R2843 VDD2.n129 VDD2.t0 1.75738
R2844 VDD2.n129 VDD2.t4 1.75738
R2845 VDD2.n127 VDD2.t7 1.75738
R2846 VDD2.n127 VDD2.t9 1.75738
R2847 VDD2.n63 VDD2.t5 1.75738
R2848 VDD2.n63 VDD2.t3 1.75738
R2849 VDD2.n61 VDD2.t2 1.75738
R2850 VDD2.n61 VDD2.t1 1.75738
R2851 VDD2.n90 VDD2.n83 1.16414
R2852 VDD2.n25 VDD2.n18 1.16414
R2853 VDD2 VDD2.n128 0.668603
R2854 VDD2.n64 VDD2.n62 0.555068
R2855 VDD2.n87 VDD2.n86 0.388379
R2856 VDD2.n22 VDD2.n21 0.388379
R2857 VDD2.n121 VDD2.n120 0.155672
R2858 VDD2.n120 VDD2.n68 0.155672
R2859 VDD2.n113 VDD2.n68 0.155672
R2860 VDD2.n113 VDD2.n112 0.155672
R2861 VDD2.n112 VDD2.n72 0.155672
R2862 VDD2.n105 VDD2.n72 0.155672
R2863 VDD2.n105 VDD2.n104 0.155672
R2864 VDD2.n104 VDD2.n76 0.155672
R2865 VDD2.n97 VDD2.n76 0.155672
R2866 VDD2.n97 VDD2.n96 0.155672
R2867 VDD2.n96 VDD2.n80 0.155672
R2868 VDD2.n89 VDD2.n80 0.155672
R2869 VDD2.n89 VDD2.n88 0.155672
R2870 VDD2.n24 VDD2.n23 0.155672
R2871 VDD2.n24 VDD2.n15 0.155672
R2872 VDD2.n31 VDD2.n15 0.155672
R2873 VDD2.n32 VDD2.n31 0.155672
R2874 VDD2.n32 VDD2.n11 0.155672
R2875 VDD2.n39 VDD2.n11 0.155672
R2876 VDD2.n40 VDD2.n39 0.155672
R2877 VDD2.n40 VDD2.n7 0.155672
R2878 VDD2.n47 VDD2.n7 0.155672
R2879 VDD2.n48 VDD2.n47 0.155672
R2880 VDD2.n48 VDD2.n3 0.155672
R2881 VDD2.n55 VDD2.n3 0.155672
R2882 VDD2.n56 VDD2.n55 0.155672
C0 VN VTAIL 10.600401f
C1 VN VDD1 0.153138f
C2 VP VTAIL 10.6147f
C3 VP VDD1 10.3829f
C4 VN VDD2 9.96895f
C5 VP VDD2 0.570772f
C6 VTAIL VDD1 10.0338f
C7 VTAIL VDD2 10.0841f
C8 VP VN 8.11774f
C9 VDD1 VDD2 2.10928f
C10 VDD2 B 6.975942f
C11 VDD1 B 6.940359f
C12 VTAIL B 7.840959f
C13 VN B 17.60824f
C14 VP B 16.139341f
C15 VDD2.n0 B 0.013796f
C16 VDD2.n1 B 0.031042f
C17 VDD2.n2 B 0.013906f
C18 VDD2.n3 B 0.024441f
C19 VDD2.n4 B 0.013133f
C20 VDD2.n5 B 0.031042f
C21 VDD2.n6 B 0.013906f
C22 VDD2.n7 B 0.024441f
C23 VDD2.n8 B 0.013133f
C24 VDD2.n9 B 0.031042f
C25 VDD2.n10 B 0.013906f
C26 VDD2.n11 B 0.024441f
C27 VDD2.n12 B 0.013133f
C28 VDD2.n13 B 0.031042f
C29 VDD2.n14 B 0.013906f
C30 VDD2.n15 B 0.024441f
C31 VDD2.n16 B 0.013133f
C32 VDD2.n17 B 0.031042f
C33 VDD2.n18 B 0.013906f
C34 VDD2.n19 B 0.136552f
C35 VDD2.t8 B 0.050873f
C36 VDD2.n20 B 0.023282f
C37 VDD2.n21 B 0.018338f
C38 VDD2.n22 B 0.013133f
C39 VDD2.n23 B 1.17234f
C40 VDD2.n24 B 0.024441f
C41 VDD2.n25 B 0.013133f
C42 VDD2.n26 B 0.013906f
C43 VDD2.n27 B 0.031042f
C44 VDD2.n28 B 0.031042f
C45 VDD2.n29 B 0.013906f
C46 VDD2.n30 B 0.013133f
C47 VDD2.n31 B 0.024441f
C48 VDD2.n32 B 0.024441f
C49 VDD2.n33 B 0.013133f
C50 VDD2.n34 B 0.013906f
C51 VDD2.n35 B 0.031042f
C52 VDD2.n36 B 0.031042f
C53 VDD2.n37 B 0.013906f
C54 VDD2.n38 B 0.013133f
C55 VDD2.n39 B 0.024441f
C56 VDD2.n40 B 0.024441f
C57 VDD2.n41 B 0.013133f
C58 VDD2.n42 B 0.013906f
C59 VDD2.n43 B 0.031042f
C60 VDD2.n44 B 0.031042f
C61 VDD2.n45 B 0.013906f
C62 VDD2.n46 B 0.013133f
C63 VDD2.n47 B 0.024441f
C64 VDD2.n48 B 0.024441f
C65 VDD2.n49 B 0.013133f
C66 VDD2.n50 B 0.013906f
C67 VDD2.n51 B 0.031042f
C68 VDD2.n52 B 0.031042f
C69 VDD2.n53 B 0.013906f
C70 VDD2.n54 B 0.013133f
C71 VDD2.n55 B 0.024441f
C72 VDD2.n56 B 0.064173f
C73 VDD2.n57 B 0.013133f
C74 VDD2.n58 B 0.013906f
C75 VDD2.n59 B 0.062245f
C76 VDD2.n60 B 0.081215f
C77 VDD2.t2 B 0.217667f
C78 VDD2.t1 B 0.217667f
C79 VDD2.n61 B 1.94281f
C80 VDD2.n62 B 0.658061f
C81 VDD2.t5 B 0.217667f
C82 VDD2.t3 B 0.217667f
C83 VDD2.n63 B 1.95679f
C84 VDD2.n64 B 2.7356f
C85 VDD2.n65 B 0.013796f
C86 VDD2.n66 B 0.031042f
C87 VDD2.n67 B 0.013906f
C88 VDD2.n68 B 0.024441f
C89 VDD2.n69 B 0.013133f
C90 VDD2.n70 B 0.031042f
C91 VDD2.n71 B 0.013906f
C92 VDD2.n72 B 0.024441f
C93 VDD2.n73 B 0.013133f
C94 VDD2.n74 B 0.031042f
C95 VDD2.n75 B 0.013906f
C96 VDD2.n76 B 0.024441f
C97 VDD2.n77 B 0.013133f
C98 VDD2.n78 B 0.031042f
C99 VDD2.n79 B 0.013906f
C100 VDD2.n80 B 0.024441f
C101 VDD2.n81 B 0.013133f
C102 VDD2.n82 B 0.031042f
C103 VDD2.n83 B 0.013906f
C104 VDD2.n84 B 0.136552f
C105 VDD2.t6 B 0.050873f
C106 VDD2.n85 B 0.023282f
C107 VDD2.n86 B 0.018338f
C108 VDD2.n87 B 0.013133f
C109 VDD2.n88 B 1.17234f
C110 VDD2.n89 B 0.024441f
C111 VDD2.n90 B 0.013133f
C112 VDD2.n91 B 0.013906f
C113 VDD2.n92 B 0.031042f
C114 VDD2.n93 B 0.031042f
C115 VDD2.n94 B 0.013906f
C116 VDD2.n95 B 0.013133f
C117 VDD2.n96 B 0.024441f
C118 VDD2.n97 B 0.024441f
C119 VDD2.n98 B 0.013133f
C120 VDD2.n99 B 0.013906f
C121 VDD2.n100 B 0.031042f
C122 VDD2.n101 B 0.031042f
C123 VDD2.n102 B 0.013906f
C124 VDD2.n103 B 0.013133f
C125 VDD2.n104 B 0.024441f
C126 VDD2.n105 B 0.024441f
C127 VDD2.n106 B 0.013133f
C128 VDD2.n107 B 0.013906f
C129 VDD2.n108 B 0.031042f
C130 VDD2.n109 B 0.031042f
C131 VDD2.n110 B 0.013906f
C132 VDD2.n111 B 0.013133f
C133 VDD2.n112 B 0.024441f
C134 VDD2.n113 B 0.024441f
C135 VDD2.n114 B 0.013133f
C136 VDD2.n115 B 0.013906f
C137 VDD2.n116 B 0.031042f
C138 VDD2.n117 B 0.031042f
C139 VDD2.n118 B 0.013906f
C140 VDD2.n119 B 0.013133f
C141 VDD2.n120 B 0.024441f
C142 VDD2.n121 B 0.064173f
C143 VDD2.n122 B 0.013133f
C144 VDD2.n123 B 0.013906f
C145 VDD2.n124 B 0.062245f
C146 VDD2.n125 B 0.07026f
C147 VDD2.n126 B 2.73493f
C148 VDD2.t7 B 0.217667f
C149 VDD2.t9 B 0.217667f
C150 VDD2.n127 B 1.94282f
C151 VDD2.n128 B 0.435252f
C152 VDD2.t0 B 0.217667f
C153 VDD2.t4 B 0.217667f
C154 VDD2.n129 B 1.95675f
C155 VN.n0 B 0.029218f
C156 VN.t6 B 1.69814f
C157 VN.n1 B 0.032663f
C158 VN.n2 B 0.022162f
C159 VN.t4 B 1.69814f
C160 VN.n3 B 0.60369f
C161 VN.n4 B 0.022162f
C162 VN.n5 B 0.041304f
C163 VN.n6 B 0.022162f
C164 VN.t8 B 1.69814f
C165 VN.n7 B 0.041304f
C166 VN.n8 B 0.022162f
C167 VN.t7 B 1.69814f
C168 VN.n9 B 0.669527f
C169 VN.t1 B 1.86958f
C170 VN.n10 B 0.650104f
C171 VN.n11 B 0.211875f
C172 VN.n12 B 0.034371f
C173 VN.n13 B 0.044647f
C174 VN.n14 B 0.020062f
C175 VN.n15 B 0.022162f
C176 VN.n16 B 0.022162f
C177 VN.n17 B 0.022162f
C178 VN.n18 B 0.041304f
C179 VN.n19 B 0.624602f
C180 VN.n20 B 0.041304f
C181 VN.n21 B 0.022162f
C182 VN.n22 B 0.022162f
C183 VN.n23 B 0.022162f
C184 VN.n24 B 0.020062f
C185 VN.n25 B 0.044647f
C186 VN.n26 B 0.034371f
C187 VN.n27 B 0.022162f
C188 VN.n28 B 0.022162f
C189 VN.n29 B 0.027845f
C190 VN.n30 B 0.041304f
C191 VN.n31 B 0.032046f
C192 VN.n32 B 0.022162f
C193 VN.n33 B 0.022162f
C194 VN.n34 B 0.022162f
C195 VN.n35 B 0.041304f
C196 VN.n36 B 0.027438f
C197 VN.n37 B 0.672415f
C198 VN.n38 B 0.036492f
C199 VN.n39 B 0.029218f
C200 VN.t3 B 1.69814f
C201 VN.n40 B 0.032663f
C202 VN.n41 B 0.022162f
C203 VN.t2 B 1.69814f
C204 VN.n42 B 0.60369f
C205 VN.n43 B 0.022162f
C206 VN.n44 B 0.041304f
C207 VN.n45 B 0.022162f
C208 VN.t0 B 1.69814f
C209 VN.n46 B 0.041304f
C210 VN.n47 B 0.022162f
C211 VN.t9 B 1.69814f
C212 VN.n48 B 0.669527f
C213 VN.t5 B 1.86958f
C214 VN.n49 B 0.650104f
C215 VN.n50 B 0.211875f
C216 VN.n51 B 0.034371f
C217 VN.n52 B 0.044647f
C218 VN.n53 B 0.020062f
C219 VN.n54 B 0.022162f
C220 VN.n55 B 0.022162f
C221 VN.n56 B 0.022162f
C222 VN.n57 B 0.041304f
C223 VN.n58 B 0.624602f
C224 VN.n59 B 0.041304f
C225 VN.n60 B 0.022162f
C226 VN.n61 B 0.022162f
C227 VN.n62 B 0.022162f
C228 VN.n63 B 0.020062f
C229 VN.n64 B 0.044647f
C230 VN.n65 B 0.034371f
C231 VN.n66 B 0.022162f
C232 VN.n67 B 0.022162f
C233 VN.n68 B 0.027845f
C234 VN.n69 B 0.041304f
C235 VN.n70 B 0.032046f
C236 VN.n71 B 0.022162f
C237 VN.n72 B 0.022162f
C238 VN.n73 B 0.022162f
C239 VN.n74 B 0.041304f
C240 VN.n75 B 0.027438f
C241 VN.n76 B 0.672415f
C242 VN.n77 B 1.31663f
C243 VDD1.n0 B 0.013926f
C244 VDD1.n1 B 0.031335f
C245 VDD1.n2 B 0.014037f
C246 VDD1.n3 B 0.024671f
C247 VDD1.n4 B 0.013257f
C248 VDD1.n5 B 0.031335f
C249 VDD1.n6 B 0.014037f
C250 VDD1.n7 B 0.024671f
C251 VDD1.n8 B 0.013257f
C252 VDD1.n9 B 0.031335f
C253 VDD1.n10 B 0.014037f
C254 VDD1.n11 B 0.024671f
C255 VDD1.n12 B 0.013257f
C256 VDD1.n13 B 0.031335f
C257 VDD1.n14 B 0.014037f
C258 VDD1.n15 B 0.024671f
C259 VDD1.n16 B 0.013257f
C260 VDD1.n17 B 0.031335f
C261 VDD1.n18 B 0.014037f
C262 VDD1.n19 B 0.137836f
C263 VDD1.t9 B 0.051352f
C264 VDD1.n20 B 0.023501f
C265 VDD1.n21 B 0.01851f
C266 VDD1.n22 B 0.013257f
C267 VDD1.n23 B 1.18337f
C268 VDD1.n24 B 0.024671f
C269 VDD1.n25 B 0.013257f
C270 VDD1.n26 B 0.014037f
C271 VDD1.n27 B 0.031335f
C272 VDD1.n28 B 0.031335f
C273 VDD1.n29 B 0.014037f
C274 VDD1.n30 B 0.013257f
C275 VDD1.n31 B 0.024671f
C276 VDD1.n32 B 0.024671f
C277 VDD1.n33 B 0.013257f
C278 VDD1.n34 B 0.014037f
C279 VDD1.n35 B 0.031335f
C280 VDD1.n36 B 0.031335f
C281 VDD1.n37 B 0.014037f
C282 VDD1.n38 B 0.013257f
C283 VDD1.n39 B 0.024671f
C284 VDD1.n40 B 0.024671f
C285 VDD1.n41 B 0.013257f
C286 VDD1.n42 B 0.014037f
C287 VDD1.n43 B 0.031335f
C288 VDD1.n44 B 0.031335f
C289 VDD1.n45 B 0.014037f
C290 VDD1.n46 B 0.013257f
C291 VDD1.n47 B 0.024671f
C292 VDD1.n48 B 0.024671f
C293 VDD1.n49 B 0.013257f
C294 VDD1.n50 B 0.014037f
C295 VDD1.n51 B 0.031335f
C296 VDD1.n52 B 0.031335f
C297 VDD1.n53 B 0.014037f
C298 VDD1.n54 B 0.013257f
C299 VDD1.n55 B 0.024671f
C300 VDD1.n56 B 0.064777f
C301 VDD1.n57 B 0.013257f
C302 VDD1.n58 B 0.014037f
C303 VDD1.n59 B 0.06283f
C304 VDD1.n60 B 0.081979f
C305 VDD1.t7 B 0.219715f
C306 VDD1.t8 B 0.219715f
C307 VDD1.n61 B 1.9611f
C308 VDD1.n62 B 0.672243f
C309 VDD1.n63 B 0.013926f
C310 VDD1.n64 B 0.031335f
C311 VDD1.n65 B 0.014037f
C312 VDD1.n66 B 0.024671f
C313 VDD1.n67 B 0.013257f
C314 VDD1.n68 B 0.031335f
C315 VDD1.n69 B 0.014037f
C316 VDD1.n70 B 0.024671f
C317 VDD1.n71 B 0.013257f
C318 VDD1.n72 B 0.031335f
C319 VDD1.n73 B 0.014037f
C320 VDD1.n74 B 0.024671f
C321 VDD1.n75 B 0.013257f
C322 VDD1.n76 B 0.031335f
C323 VDD1.n77 B 0.014037f
C324 VDD1.n78 B 0.024671f
C325 VDD1.n79 B 0.013257f
C326 VDD1.n80 B 0.031335f
C327 VDD1.n81 B 0.014037f
C328 VDD1.n82 B 0.137836f
C329 VDD1.t2 B 0.051352f
C330 VDD1.n83 B 0.023501f
C331 VDD1.n84 B 0.01851f
C332 VDD1.n85 B 0.013257f
C333 VDD1.n86 B 1.18337f
C334 VDD1.n87 B 0.024671f
C335 VDD1.n88 B 0.013257f
C336 VDD1.n89 B 0.014037f
C337 VDD1.n90 B 0.031335f
C338 VDD1.n91 B 0.031335f
C339 VDD1.n92 B 0.014037f
C340 VDD1.n93 B 0.013257f
C341 VDD1.n94 B 0.024671f
C342 VDD1.n95 B 0.024671f
C343 VDD1.n96 B 0.013257f
C344 VDD1.n97 B 0.014037f
C345 VDD1.n98 B 0.031335f
C346 VDD1.n99 B 0.031335f
C347 VDD1.n100 B 0.014037f
C348 VDD1.n101 B 0.013257f
C349 VDD1.n102 B 0.024671f
C350 VDD1.n103 B 0.024671f
C351 VDD1.n104 B 0.013257f
C352 VDD1.n105 B 0.014037f
C353 VDD1.n106 B 0.031335f
C354 VDD1.n107 B 0.031335f
C355 VDD1.n108 B 0.014037f
C356 VDD1.n109 B 0.013257f
C357 VDD1.n110 B 0.024671f
C358 VDD1.n111 B 0.024671f
C359 VDD1.n112 B 0.013257f
C360 VDD1.n113 B 0.014037f
C361 VDD1.n114 B 0.031335f
C362 VDD1.n115 B 0.031335f
C363 VDD1.n116 B 0.014037f
C364 VDD1.n117 B 0.013257f
C365 VDD1.n118 B 0.024671f
C366 VDD1.n119 B 0.064777f
C367 VDD1.n120 B 0.013257f
C368 VDD1.n121 B 0.014037f
C369 VDD1.n122 B 0.06283f
C370 VDD1.n123 B 0.081979f
C371 VDD1.t6 B 0.219715f
C372 VDD1.t1 B 0.219715f
C373 VDD1.n124 B 1.96109f
C374 VDD1.n125 B 0.664253f
C375 VDD1.t0 B 0.219715f
C376 VDD1.t4 B 0.219715f
C377 VDD1.n126 B 1.9752f
C378 VDD1.n127 B 2.88162f
C379 VDD1.t5 B 0.219715f
C380 VDD1.t3 B 0.219715f
C381 VDD1.n128 B 1.96109f
C382 VDD1.n129 B 3.02456f
C383 VTAIL.t0 B 0.223589f
C384 VTAIL.t1 B 0.223589f
C385 VTAIL.n0 B 1.93091f
C386 VTAIL.n1 B 0.515746f
C387 VTAIL.n2 B 0.014172f
C388 VTAIL.n3 B 0.031887f
C389 VTAIL.n4 B 0.014284f
C390 VTAIL.n5 B 0.025106f
C391 VTAIL.n6 B 0.013491f
C392 VTAIL.n7 B 0.031887f
C393 VTAIL.n8 B 0.014284f
C394 VTAIL.n9 B 0.025106f
C395 VTAIL.n10 B 0.013491f
C396 VTAIL.n11 B 0.031887f
C397 VTAIL.n12 B 0.014284f
C398 VTAIL.n13 B 0.025106f
C399 VTAIL.n14 B 0.013491f
C400 VTAIL.n15 B 0.031887f
C401 VTAIL.n16 B 0.014284f
C402 VTAIL.n17 B 0.025106f
C403 VTAIL.n18 B 0.013491f
C404 VTAIL.n19 B 0.031887f
C405 VTAIL.n20 B 0.014284f
C406 VTAIL.n21 B 0.140267f
C407 VTAIL.t16 B 0.052257f
C408 VTAIL.n22 B 0.023915f
C409 VTAIL.n23 B 0.018837f
C410 VTAIL.n24 B 0.013491f
C411 VTAIL.n25 B 1.20424f
C412 VTAIL.n26 B 0.025106f
C413 VTAIL.n27 B 0.013491f
C414 VTAIL.n28 B 0.014284f
C415 VTAIL.n29 B 0.031887f
C416 VTAIL.n30 B 0.031887f
C417 VTAIL.n31 B 0.014284f
C418 VTAIL.n32 B 0.013491f
C419 VTAIL.n33 B 0.025106f
C420 VTAIL.n34 B 0.025106f
C421 VTAIL.n35 B 0.013491f
C422 VTAIL.n36 B 0.014284f
C423 VTAIL.n37 B 0.031887f
C424 VTAIL.n38 B 0.031887f
C425 VTAIL.n39 B 0.014284f
C426 VTAIL.n40 B 0.013491f
C427 VTAIL.n41 B 0.025106f
C428 VTAIL.n42 B 0.025106f
C429 VTAIL.n43 B 0.013491f
C430 VTAIL.n44 B 0.014284f
C431 VTAIL.n45 B 0.031887f
C432 VTAIL.n46 B 0.031887f
C433 VTAIL.n47 B 0.014284f
C434 VTAIL.n48 B 0.013491f
C435 VTAIL.n49 B 0.025106f
C436 VTAIL.n50 B 0.025106f
C437 VTAIL.n51 B 0.013491f
C438 VTAIL.n52 B 0.014284f
C439 VTAIL.n53 B 0.031887f
C440 VTAIL.n54 B 0.031887f
C441 VTAIL.n55 B 0.014284f
C442 VTAIL.n56 B 0.013491f
C443 VTAIL.n57 B 0.025106f
C444 VTAIL.n58 B 0.065919f
C445 VTAIL.n59 B 0.013491f
C446 VTAIL.n60 B 0.014284f
C447 VTAIL.n61 B 0.063938f
C448 VTAIL.n62 B 0.05487f
C449 VTAIL.n63 B 0.358008f
C450 VTAIL.t7 B 0.223589f
C451 VTAIL.t12 B 0.223589f
C452 VTAIL.n64 B 1.93091f
C453 VTAIL.n65 B 0.621051f
C454 VTAIL.t8 B 0.223589f
C455 VTAIL.t10 B 0.223589f
C456 VTAIL.n66 B 1.93091f
C457 VTAIL.n67 B 1.94539f
C458 VTAIL.t3 B 0.223589f
C459 VTAIL.t4 B 0.223589f
C460 VTAIL.n68 B 1.93091f
C461 VTAIL.n69 B 1.94538f
C462 VTAIL.t5 B 0.223589f
C463 VTAIL.t2 B 0.223589f
C464 VTAIL.n70 B 1.93091f
C465 VTAIL.n71 B 0.621045f
C466 VTAIL.n72 B 0.014172f
C467 VTAIL.n73 B 0.031887f
C468 VTAIL.n74 B 0.014284f
C469 VTAIL.n75 B 0.025106f
C470 VTAIL.n76 B 0.013491f
C471 VTAIL.n77 B 0.031887f
C472 VTAIL.n78 B 0.014284f
C473 VTAIL.n79 B 0.025106f
C474 VTAIL.n80 B 0.013491f
C475 VTAIL.n81 B 0.031887f
C476 VTAIL.n82 B 0.014284f
C477 VTAIL.n83 B 0.025106f
C478 VTAIL.n84 B 0.013491f
C479 VTAIL.n85 B 0.031887f
C480 VTAIL.n86 B 0.014284f
C481 VTAIL.n87 B 0.025106f
C482 VTAIL.n88 B 0.013491f
C483 VTAIL.n89 B 0.031887f
C484 VTAIL.n90 B 0.014284f
C485 VTAIL.n91 B 0.140267f
C486 VTAIL.t6 B 0.052257f
C487 VTAIL.n92 B 0.023915f
C488 VTAIL.n93 B 0.018837f
C489 VTAIL.n94 B 0.013491f
C490 VTAIL.n95 B 1.20424f
C491 VTAIL.n96 B 0.025106f
C492 VTAIL.n97 B 0.013491f
C493 VTAIL.n98 B 0.014284f
C494 VTAIL.n99 B 0.031887f
C495 VTAIL.n100 B 0.031887f
C496 VTAIL.n101 B 0.014284f
C497 VTAIL.n102 B 0.013491f
C498 VTAIL.n103 B 0.025106f
C499 VTAIL.n104 B 0.025106f
C500 VTAIL.n105 B 0.013491f
C501 VTAIL.n106 B 0.014284f
C502 VTAIL.n107 B 0.031887f
C503 VTAIL.n108 B 0.031887f
C504 VTAIL.n109 B 0.014284f
C505 VTAIL.n110 B 0.013491f
C506 VTAIL.n111 B 0.025106f
C507 VTAIL.n112 B 0.025106f
C508 VTAIL.n113 B 0.013491f
C509 VTAIL.n114 B 0.014284f
C510 VTAIL.n115 B 0.031887f
C511 VTAIL.n116 B 0.031887f
C512 VTAIL.n117 B 0.014284f
C513 VTAIL.n118 B 0.013491f
C514 VTAIL.n119 B 0.025106f
C515 VTAIL.n120 B 0.025106f
C516 VTAIL.n121 B 0.013491f
C517 VTAIL.n122 B 0.014284f
C518 VTAIL.n123 B 0.031887f
C519 VTAIL.n124 B 0.031887f
C520 VTAIL.n125 B 0.014284f
C521 VTAIL.n126 B 0.013491f
C522 VTAIL.n127 B 0.025106f
C523 VTAIL.n128 B 0.065919f
C524 VTAIL.n129 B 0.013491f
C525 VTAIL.n130 B 0.014284f
C526 VTAIL.n131 B 0.063938f
C527 VTAIL.n132 B 0.05487f
C528 VTAIL.n133 B 0.358008f
C529 VTAIL.t9 B 0.223589f
C530 VTAIL.t11 B 0.223589f
C531 VTAIL.n134 B 1.93091f
C532 VTAIL.n135 B 0.560373f
C533 VTAIL.t15 B 0.223589f
C534 VTAIL.t13 B 0.223589f
C535 VTAIL.n136 B 1.93091f
C536 VTAIL.n137 B 0.621045f
C537 VTAIL.n138 B 0.014172f
C538 VTAIL.n139 B 0.031887f
C539 VTAIL.n140 B 0.014284f
C540 VTAIL.n141 B 0.025106f
C541 VTAIL.n142 B 0.013491f
C542 VTAIL.n143 B 0.031887f
C543 VTAIL.n144 B 0.014284f
C544 VTAIL.n145 B 0.025106f
C545 VTAIL.n146 B 0.013491f
C546 VTAIL.n147 B 0.031887f
C547 VTAIL.n148 B 0.014284f
C548 VTAIL.n149 B 0.025106f
C549 VTAIL.n150 B 0.013491f
C550 VTAIL.n151 B 0.031887f
C551 VTAIL.n152 B 0.014284f
C552 VTAIL.n153 B 0.025106f
C553 VTAIL.n154 B 0.013491f
C554 VTAIL.n155 B 0.031887f
C555 VTAIL.n156 B 0.014284f
C556 VTAIL.n157 B 0.140267f
C557 VTAIL.t14 B 0.052257f
C558 VTAIL.n158 B 0.023915f
C559 VTAIL.n159 B 0.018837f
C560 VTAIL.n160 B 0.013491f
C561 VTAIL.n161 B 1.20424f
C562 VTAIL.n162 B 0.025106f
C563 VTAIL.n163 B 0.013491f
C564 VTAIL.n164 B 0.014284f
C565 VTAIL.n165 B 0.031887f
C566 VTAIL.n166 B 0.031887f
C567 VTAIL.n167 B 0.014284f
C568 VTAIL.n168 B 0.013491f
C569 VTAIL.n169 B 0.025106f
C570 VTAIL.n170 B 0.025106f
C571 VTAIL.n171 B 0.013491f
C572 VTAIL.n172 B 0.014284f
C573 VTAIL.n173 B 0.031887f
C574 VTAIL.n174 B 0.031887f
C575 VTAIL.n175 B 0.014284f
C576 VTAIL.n176 B 0.013491f
C577 VTAIL.n177 B 0.025106f
C578 VTAIL.n178 B 0.025106f
C579 VTAIL.n179 B 0.013491f
C580 VTAIL.n180 B 0.014284f
C581 VTAIL.n181 B 0.031887f
C582 VTAIL.n182 B 0.031887f
C583 VTAIL.n183 B 0.014284f
C584 VTAIL.n184 B 0.013491f
C585 VTAIL.n185 B 0.025106f
C586 VTAIL.n186 B 0.025106f
C587 VTAIL.n187 B 0.013491f
C588 VTAIL.n188 B 0.014284f
C589 VTAIL.n189 B 0.031887f
C590 VTAIL.n190 B 0.031887f
C591 VTAIL.n191 B 0.014284f
C592 VTAIL.n192 B 0.013491f
C593 VTAIL.n193 B 0.025106f
C594 VTAIL.n194 B 0.065919f
C595 VTAIL.n195 B 0.013491f
C596 VTAIL.n196 B 0.014284f
C597 VTAIL.n197 B 0.063938f
C598 VTAIL.n198 B 0.05487f
C599 VTAIL.n199 B 1.54566f
C600 VTAIL.n200 B 0.014172f
C601 VTAIL.n201 B 0.031887f
C602 VTAIL.n202 B 0.014284f
C603 VTAIL.n203 B 0.025106f
C604 VTAIL.n204 B 0.013491f
C605 VTAIL.n205 B 0.031887f
C606 VTAIL.n206 B 0.014284f
C607 VTAIL.n207 B 0.025106f
C608 VTAIL.n208 B 0.013491f
C609 VTAIL.n209 B 0.031887f
C610 VTAIL.n210 B 0.014284f
C611 VTAIL.n211 B 0.025106f
C612 VTAIL.n212 B 0.013491f
C613 VTAIL.n213 B 0.031887f
C614 VTAIL.n214 B 0.014284f
C615 VTAIL.n215 B 0.025106f
C616 VTAIL.n216 B 0.013491f
C617 VTAIL.n217 B 0.031887f
C618 VTAIL.n218 B 0.014284f
C619 VTAIL.n219 B 0.140267f
C620 VTAIL.t18 B 0.052257f
C621 VTAIL.n220 B 0.023915f
C622 VTAIL.n221 B 0.018837f
C623 VTAIL.n222 B 0.013491f
C624 VTAIL.n223 B 1.20424f
C625 VTAIL.n224 B 0.025106f
C626 VTAIL.n225 B 0.013491f
C627 VTAIL.n226 B 0.014284f
C628 VTAIL.n227 B 0.031887f
C629 VTAIL.n228 B 0.031887f
C630 VTAIL.n229 B 0.014284f
C631 VTAIL.n230 B 0.013491f
C632 VTAIL.n231 B 0.025106f
C633 VTAIL.n232 B 0.025106f
C634 VTAIL.n233 B 0.013491f
C635 VTAIL.n234 B 0.014284f
C636 VTAIL.n235 B 0.031887f
C637 VTAIL.n236 B 0.031887f
C638 VTAIL.n237 B 0.014284f
C639 VTAIL.n238 B 0.013491f
C640 VTAIL.n239 B 0.025106f
C641 VTAIL.n240 B 0.025106f
C642 VTAIL.n241 B 0.013491f
C643 VTAIL.n242 B 0.014284f
C644 VTAIL.n243 B 0.031887f
C645 VTAIL.n244 B 0.031887f
C646 VTAIL.n245 B 0.014284f
C647 VTAIL.n246 B 0.013491f
C648 VTAIL.n247 B 0.025106f
C649 VTAIL.n248 B 0.025106f
C650 VTAIL.n249 B 0.013491f
C651 VTAIL.n250 B 0.014284f
C652 VTAIL.n251 B 0.031887f
C653 VTAIL.n252 B 0.031887f
C654 VTAIL.n253 B 0.014284f
C655 VTAIL.n254 B 0.013491f
C656 VTAIL.n255 B 0.025106f
C657 VTAIL.n256 B 0.065919f
C658 VTAIL.n257 B 0.013491f
C659 VTAIL.n258 B 0.014284f
C660 VTAIL.n259 B 0.063938f
C661 VTAIL.n260 B 0.05487f
C662 VTAIL.n261 B 1.54566f
C663 VTAIL.t19 B 0.223589f
C664 VTAIL.t17 B 0.223589f
C665 VTAIL.n262 B 1.93091f
C666 VTAIL.n263 B 0.468324f
C667 VP.n0 B 0.029658f
C668 VP.t5 B 1.72368f
C669 VP.n1 B 0.033154f
C670 VP.n2 B 0.022495f
C671 VP.t9 B 1.72368f
C672 VP.n3 B 0.612769f
C673 VP.n4 B 0.022495f
C674 VP.n5 B 0.041925f
C675 VP.n6 B 0.022495f
C676 VP.t8 B 1.72368f
C677 VP.n7 B 0.041925f
C678 VP.n8 B 0.022495f
C679 VP.t3 B 1.72368f
C680 VP.n9 B 0.612769f
C681 VP.n10 B 0.022495f
C682 VP.n11 B 0.033154f
C683 VP.n12 B 0.029658f
C684 VP.t7 B 1.72368f
C685 VP.n13 B 0.029658f
C686 VP.t6 B 1.72368f
C687 VP.n14 B 0.033154f
C688 VP.n15 B 0.022495f
C689 VP.t4 B 1.72368f
C690 VP.n16 B 0.612769f
C691 VP.n17 B 0.022495f
C692 VP.n18 B 0.041925f
C693 VP.n19 B 0.022495f
C694 VP.t1 B 1.72368f
C695 VP.n20 B 0.041925f
C696 VP.n21 B 0.022495f
C697 VP.t2 B 1.72368f
C698 VP.n22 B 0.679596f
C699 VP.t0 B 1.89769f
C700 VP.n23 B 0.65988f
C701 VP.n24 B 0.215062f
C702 VP.n25 B 0.034888f
C703 VP.n26 B 0.045318f
C704 VP.n27 B 0.020364f
C705 VP.n28 B 0.022495f
C706 VP.n29 B 0.022495f
C707 VP.n30 B 0.022495f
C708 VP.n31 B 0.041925f
C709 VP.n32 B 0.633996f
C710 VP.n33 B 0.041925f
C711 VP.n34 B 0.022495f
C712 VP.n35 B 0.022495f
C713 VP.n36 B 0.022495f
C714 VP.n37 B 0.020364f
C715 VP.n38 B 0.045318f
C716 VP.n39 B 0.034888f
C717 VP.n40 B 0.022495f
C718 VP.n41 B 0.022495f
C719 VP.n42 B 0.028264f
C720 VP.n43 B 0.041925f
C721 VP.n44 B 0.032528f
C722 VP.n45 B 0.022495f
C723 VP.n46 B 0.022495f
C724 VP.n47 B 0.022495f
C725 VP.n48 B 0.041925f
C726 VP.n49 B 0.02785f
C727 VP.n50 B 0.682527f
C728 VP.n51 B 1.32441f
C729 VP.n52 B 1.33997f
C730 VP.n53 B 0.682527f
C731 VP.n54 B 0.02785f
C732 VP.n55 B 0.041925f
C733 VP.n56 B 0.022495f
C734 VP.n57 B 0.022495f
C735 VP.n58 B 0.022495f
C736 VP.n59 B 0.032528f
C737 VP.n60 B 0.041925f
C738 VP.n61 B 0.028264f
C739 VP.n62 B 0.022495f
C740 VP.n63 B 0.022495f
C741 VP.n64 B 0.034888f
C742 VP.n65 B 0.045318f
C743 VP.n66 B 0.020364f
C744 VP.n67 B 0.022495f
C745 VP.n68 B 0.022495f
C746 VP.n69 B 0.022495f
C747 VP.n70 B 0.041925f
C748 VP.n71 B 0.633996f
C749 VP.n72 B 0.041925f
C750 VP.n73 B 0.022495f
C751 VP.n74 B 0.022495f
C752 VP.n75 B 0.022495f
C753 VP.n76 B 0.020364f
C754 VP.n77 B 0.045318f
C755 VP.n78 B 0.034888f
C756 VP.n79 B 0.022495f
C757 VP.n80 B 0.022495f
C758 VP.n81 B 0.028264f
C759 VP.n82 B 0.041925f
C760 VP.n83 B 0.032528f
C761 VP.n84 B 0.022495f
C762 VP.n85 B 0.022495f
C763 VP.n86 B 0.022495f
C764 VP.n87 B 0.041925f
C765 VP.n88 B 0.02785f
C766 VP.n89 B 0.682527f
C767 VP.n90 B 0.037041f
.ends

