* NGSPICE file created from diff_pair_sample_0201.ext - technology: sky130A

.subckt diff_pair_sample_0201 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t1 VN.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.7254 pd=4.5 as=0.7254 ps=4.5 w=1.86 l=0.81
X1 VDD1.t1 VP.t0 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=0.7254 pd=4.5 as=0.7254 ps=4.5 w=1.86 l=0.81
X2 B.t15 B.t13 B.t14 B.t3 sky130_fd_pr__nfet_01v8 ad=0.7254 pd=4.5 as=0 ps=0 w=1.86 l=0.81
X3 VDD2.t0 VN.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.7254 pd=4.5 as=0.7254 ps=4.5 w=1.86 l=0.81
X4 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=0.7254 pd=4.5 as=0 ps=0 w=1.86 l=0.81
X5 VDD1.t0 VP.t1 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=0.7254 pd=4.5 as=0.7254 ps=4.5 w=1.86 l=0.81
X6 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=0.7254 pd=4.5 as=0 ps=0 w=1.86 l=0.81
X7 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=0.7254 pd=4.5 as=0 ps=0 w=1.86 l=0.81
R0 VN VN.t0 298.356
R1 VN VN.t1 265.784
R2 VTAIL.n26 VTAIL.n24 289.615
R3 VTAIL.n2 VTAIL.n0 289.615
R4 VTAIL.n18 VTAIL.n16 289.615
R5 VTAIL.n10 VTAIL.n8 289.615
R6 VTAIL.n27 VTAIL.n26 185
R7 VTAIL.n3 VTAIL.n2 185
R8 VTAIL.n19 VTAIL.n18 185
R9 VTAIL.n11 VTAIL.n10 185
R10 VTAIL.t0 VTAIL.n25 164.876
R11 VTAIL.t3 VTAIL.n1 164.876
R12 VTAIL.t2 VTAIL.n17 164.876
R13 VTAIL.t1 VTAIL.n9 164.876
R14 VTAIL.n26 VTAIL.t0 52.3082
R15 VTAIL.n2 VTAIL.t3 52.3082
R16 VTAIL.n18 VTAIL.t2 52.3082
R17 VTAIL.n10 VTAIL.t1 52.3082
R18 VTAIL.n31 VTAIL.n30 35.6763
R19 VTAIL.n7 VTAIL.n6 35.6763
R20 VTAIL.n23 VTAIL.n22 35.6763
R21 VTAIL.n15 VTAIL.n14 35.6763
R22 VTAIL.n15 VTAIL.n7 15.9531
R23 VTAIL.n31 VTAIL.n23 14.9703
R24 VTAIL.n27 VTAIL.n25 14.7318
R25 VTAIL.n3 VTAIL.n1 14.7318
R26 VTAIL.n19 VTAIL.n17 14.7318
R27 VTAIL.n11 VTAIL.n9 14.7318
R28 VTAIL.n28 VTAIL.n24 12.8005
R29 VTAIL.n4 VTAIL.n0 12.8005
R30 VTAIL.n20 VTAIL.n16 12.8005
R31 VTAIL.n12 VTAIL.n8 12.8005
R32 VTAIL.n30 VTAIL.n29 9.45567
R33 VTAIL.n6 VTAIL.n5 9.45567
R34 VTAIL.n22 VTAIL.n21 9.45567
R35 VTAIL.n14 VTAIL.n13 9.45567
R36 VTAIL.n29 VTAIL.n28 9.3005
R37 VTAIL.n5 VTAIL.n4 9.3005
R38 VTAIL.n21 VTAIL.n20 9.3005
R39 VTAIL.n13 VTAIL.n12 9.3005
R40 VTAIL.n29 VTAIL.n25 5.62509
R41 VTAIL.n5 VTAIL.n1 5.62509
R42 VTAIL.n21 VTAIL.n17 5.62509
R43 VTAIL.n13 VTAIL.n9 5.62509
R44 VTAIL.n30 VTAIL.n24 1.16414
R45 VTAIL.n6 VTAIL.n0 1.16414
R46 VTAIL.n22 VTAIL.n16 1.16414
R47 VTAIL.n14 VTAIL.n8 1.16414
R48 VTAIL.n23 VTAIL.n15 0.961707
R49 VTAIL VTAIL.n7 0.774207
R50 VTAIL.n28 VTAIL.n27 0.388379
R51 VTAIL.n4 VTAIL.n3 0.388379
R52 VTAIL.n20 VTAIL.n19 0.388379
R53 VTAIL.n12 VTAIL.n11 0.388379
R54 VTAIL VTAIL.n31 0.188
R55 VDD2.n9 VDD2.n7 289.615
R56 VDD2.n2 VDD2.n0 289.615
R57 VDD2.n10 VDD2.n9 185
R58 VDD2.n3 VDD2.n2 185
R59 VDD2.t1 VDD2.n8 164.876
R60 VDD2.t0 VDD2.n1 164.876
R61 VDD2.n14 VDD2.n6 79.6007
R62 VDD2.n14 VDD2.n13 52.355
R63 VDD2.n9 VDD2.t1 52.3082
R64 VDD2.n2 VDD2.t0 52.3082
R65 VDD2.n10 VDD2.n8 14.7318
R66 VDD2.n3 VDD2.n1 14.7318
R67 VDD2.n11 VDD2.n7 12.8005
R68 VDD2.n4 VDD2.n0 12.8005
R69 VDD2.n13 VDD2.n12 9.45567
R70 VDD2.n6 VDD2.n5 9.45567
R71 VDD2.n12 VDD2.n11 9.3005
R72 VDD2.n5 VDD2.n4 9.3005
R73 VDD2.n12 VDD2.n8 5.62509
R74 VDD2.n5 VDD2.n1 5.62509
R75 VDD2.n13 VDD2.n7 1.16414
R76 VDD2.n6 VDD2.n0 1.16414
R77 VDD2.n11 VDD2.n10 0.388379
R78 VDD2.n4 VDD2.n3 0.388379
R79 VDD2 VDD2.n14 0.304379
R80 B.n296 B.n295 585
R81 B.n297 B.n296 585
R82 B.n114 B.n48 585
R83 B.n113 B.n112 585
R84 B.n111 B.n110 585
R85 B.n109 B.n108 585
R86 B.n107 B.n106 585
R87 B.n105 B.n104 585
R88 B.n103 B.n102 585
R89 B.n101 B.n100 585
R90 B.n99 B.n98 585
R91 B.n97 B.n96 585
R92 B.n95 B.n94 585
R93 B.n92 B.n91 585
R94 B.n90 B.n89 585
R95 B.n88 B.n87 585
R96 B.n86 B.n85 585
R97 B.n84 B.n83 585
R98 B.n82 B.n81 585
R99 B.n80 B.n79 585
R100 B.n78 B.n77 585
R101 B.n76 B.n75 585
R102 B.n74 B.n73 585
R103 B.n72 B.n71 585
R104 B.n70 B.n69 585
R105 B.n68 B.n67 585
R106 B.n66 B.n65 585
R107 B.n64 B.n63 585
R108 B.n62 B.n61 585
R109 B.n60 B.n59 585
R110 B.n58 B.n57 585
R111 B.n56 B.n55 585
R112 B.n32 B.n31 585
R113 B.n300 B.n299 585
R114 B.n294 B.n49 585
R115 B.n49 B.n29 585
R116 B.n293 B.n28 585
R117 B.n304 B.n28 585
R118 B.n292 B.n27 585
R119 B.n305 B.n27 585
R120 B.n291 B.n26 585
R121 B.n306 B.n26 585
R122 B.n290 B.n289 585
R123 B.n289 B.n22 585
R124 B.n288 B.n21 585
R125 B.n312 B.n21 585
R126 B.n287 B.n20 585
R127 B.n313 B.n20 585
R128 B.n286 B.n19 585
R129 B.n314 B.n19 585
R130 B.n285 B.n284 585
R131 B.n284 B.n15 585
R132 B.n283 B.n14 585
R133 B.n320 B.n14 585
R134 B.n282 B.n13 585
R135 B.n321 B.n13 585
R136 B.n281 B.n12 585
R137 B.n322 B.n12 585
R138 B.n280 B.n279 585
R139 B.n279 B.n8 585
R140 B.n278 B.n7 585
R141 B.n328 B.n7 585
R142 B.n277 B.n6 585
R143 B.n329 B.n6 585
R144 B.n276 B.n5 585
R145 B.n330 B.n5 585
R146 B.n275 B.n274 585
R147 B.n274 B.n4 585
R148 B.n273 B.n115 585
R149 B.n273 B.n272 585
R150 B.n263 B.n116 585
R151 B.n117 B.n116 585
R152 B.n265 B.n264 585
R153 B.n266 B.n265 585
R154 B.n262 B.n122 585
R155 B.n122 B.n121 585
R156 B.n261 B.n260 585
R157 B.n260 B.n259 585
R158 B.n124 B.n123 585
R159 B.n125 B.n124 585
R160 B.n252 B.n251 585
R161 B.n253 B.n252 585
R162 B.n250 B.n130 585
R163 B.n130 B.n129 585
R164 B.n249 B.n248 585
R165 B.n248 B.n247 585
R166 B.n132 B.n131 585
R167 B.n133 B.n132 585
R168 B.n240 B.n239 585
R169 B.n241 B.n240 585
R170 B.n238 B.n138 585
R171 B.n138 B.n137 585
R172 B.n237 B.n236 585
R173 B.n236 B.n235 585
R174 B.n140 B.n139 585
R175 B.n141 B.n140 585
R176 B.n231 B.n230 585
R177 B.n144 B.n143 585
R178 B.n227 B.n226 585
R179 B.n228 B.n227 585
R180 B.n225 B.n160 585
R181 B.n224 B.n223 585
R182 B.n222 B.n221 585
R183 B.n220 B.n219 585
R184 B.n218 B.n217 585
R185 B.n216 B.n215 585
R186 B.n214 B.n213 585
R187 B.n212 B.n211 585
R188 B.n210 B.n209 585
R189 B.n207 B.n206 585
R190 B.n205 B.n204 585
R191 B.n203 B.n202 585
R192 B.n201 B.n200 585
R193 B.n199 B.n198 585
R194 B.n197 B.n196 585
R195 B.n195 B.n194 585
R196 B.n193 B.n192 585
R197 B.n191 B.n190 585
R198 B.n189 B.n188 585
R199 B.n187 B.n186 585
R200 B.n185 B.n184 585
R201 B.n183 B.n182 585
R202 B.n181 B.n180 585
R203 B.n179 B.n178 585
R204 B.n177 B.n176 585
R205 B.n175 B.n174 585
R206 B.n173 B.n172 585
R207 B.n171 B.n170 585
R208 B.n169 B.n168 585
R209 B.n167 B.n166 585
R210 B.n232 B.n142 585
R211 B.n142 B.n141 585
R212 B.n234 B.n233 585
R213 B.n235 B.n234 585
R214 B.n136 B.n135 585
R215 B.n137 B.n136 585
R216 B.n243 B.n242 585
R217 B.n242 B.n241 585
R218 B.n244 B.n134 585
R219 B.n134 B.n133 585
R220 B.n246 B.n245 585
R221 B.n247 B.n246 585
R222 B.n128 B.n127 585
R223 B.n129 B.n128 585
R224 B.n255 B.n254 585
R225 B.n254 B.n253 585
R226 B.n256 B.n126 585
R227 B.n126 B.n125 585
R228 B.n258 B.n257 585
R229 B.n259 B.n258 585
R230 B.n120 B.n119 585
R231 B.n121 B.n120 585
R232 B.n268 B.n267 585
R233 B.n267 B.n266 585
R234 B.n269 B.n118 585
R235 B.n118 B.n117 585
R236 B.n271 B.n270 585
R237 B.n272 B.n271 585
R238 B.n2 B.n0 585
R239 B.n4 B.n2 585
R240 B.n3 B.n1 585
R241 B.n329 B.n3 585
R242 B.n327 B.n326 585
R243 B.n328 B.n327 585
R244 B.n325 B.n9 585
R245 B.n9 B.n8 585
R246 B.n324 B.n323 585
R247 B.n323 B.n322 585
R248 B.n11 B.n10 585
R249 B.n321 B.n11 585
R250 B.n319 B.n318 585
R251 B.n320 B.n319 585
R252 B.n317 B.n16 585
R253 B.n16 B.n15 585
R254 B.n316 B.n315 585
R255 B.n315 B.n314 585
R256 B.n18 B.n17 585
R257 B.n313 B.n18 585
R258 B.n311 B.n310 585
R259 B.n312 B.n311 585
R260 B.n309 B.n23 585
R261 B.n23 B.n22 585
R262 B.n308 B.n307 585
R263 B.n307 B.n306 585
R264 B.n25 B.n24 585
R265 B.n305 B.n25 585
R266 B.n303 B.n302 585
R267 B.n304 B.n303 585
R268 B.n301 B.n30 585
R269 B.n30 B.n29 585
R270 B.n332 B.n331 585
R271 B.n331 B.n330 585
R272 B.n230 B.n142 492.5
R273 B.n299 B.n30 492.5
R274 B.n166 B.n140 492.5
R275 B.n296 B.n49 492.5
R276 B.n163 B.t13 257.868
R277 B.n50 B.t6 257.868
R278 B.n161 B.t2 257.435
R279 B.n52 B.t10 257.435
R280 B.n297 B.n47 256.663
R281 B.n297 B.n46 256.663
R282 B.n297 B.n45 256.663
R283 B.n297 B.n44 256.663
R284 B.n297 B.n43 256.663
R285 B.n297 B.n42 256.663
R286 B.n297 B.n41 256.663
R287 B.n297 B.n40 256.663
R288 B.n297 B.n39 256.663
R289 B.n297 B.n38 256.663
R290 B.n297 B.n37 256.663
R291 B.n297 B.n36 256.663
R292 B.n297 B.n35 256.663
R293 B.n297 B.n34 256.663
R294 B.n297 B.n33 256.663
R295 B.n298 B.n297 256.663
R296 B.n229 B.n228 256.663
R297 B.n228 B.n145 256.663
R298 B.n228 B.n146 256.663
R299 B.n228 B.n147 256.663
R300 B.n228 B.n148 256.663
R301 B.n228 B.n149 256.663
R302 B.n228 B.n150 256.663
R303 B.n228 B.n151 256.663
R304 B.n228 B.n152 256.663
R305 B.n228 B.n153 256.663
R306 B.n228 B.n154 256.663
R307 B.n228 B.n155 256.663
R308 B.n228 B.n156 256.663
R309 B.n228 B.n157 256.663
R310 B.n228 B.n158 256.663
R311 B.n228 B.n159 256.663
R312 B.n228 B.n141 170.65
R313 B.n297 B.n29 170.65
R314 B.n234 B.n142 163.367
R315 B.n234 B.n136 163.367
R316 B.n242 B.n136 163.367
R317 B.n242 B.n134 163.367
R318 B.n246 B.n134 163.367
R319 B.n246 B.n128 163.367
R320 B.n254 B.n128 163.367
R321 B.n254 B.n126 163.367
R322 B.n258 B.n126 163.367
R323 B.n258 B.n120 163.367
R324 B.n267 B.n120 163.367
R325 B.n267 B.n118 163.367
R326 B.n271 B.n118 163.367
R327 B.n271 B.n2 163.367
R328 B.n331 B.n2 163.367
R329 B.n331 B.n3 163.367
R330 B.n327 B.n3 163.367
R331 B.n327 B.n9 163.367
R332 B.n323 B.n9 163.367
R333 B.n323 B.n11 163.367
R334 B.n319 B.n11 163.367
R335 B.n319 B.n16 163.367
R336 B.n315 B.n16 163.367
R337 B.n315 B.n18 163.367
R338 B.n311 B.n18 163.367
R339 B.n311 B.n23 163.367
R340 B.n307 B.n23 163.367
R341 B.n307 B.n25 163.367
R342 B.n303 B.n25 163.367
R343 B.n303 B.n30 163.367
R344 B.n227 B.n144 163.367
R345 B.n227 B.n160 163.367
R346 B.n223 B.n222 163.367
R347 B.n219 B.n218 163.367
R348 B.n215 B.n214 163.367
R349 B.n211 B.n210 163.367
R350 B.n206 B.n205 163.367
R351 B.n202 B.n201 163.367
R352 B.n198 B.n197 163.367
R353 B.n194 B.n193 163.367
R354 B.n190 B.n189 163.367
R355 B.n186 B.n185 163.367
R356 B.n182 B.n181 163.367
R357 B.n178 B.n177 163.367
R358 B.n174 B.n173 163.367
R359 B.n170 B.n169 163.367
R360 B.n236 B.n140 163.367
R361 B.n236 B.n138 163.367
R362 B.n240 B.n138 163.367
R363 B.n240 B.n132 163.367
R364 B.n248 B.n132 163.367
R365 B.n248 B.n130 163.367
R366 B.n252 B.n130 163.367
R367 B.n252 B.n124 163.367
R368 B.n260 B.n124 163.367
R369 B.n260 B.n122 163.367
R370 B.n265 B.n122 163.367
R371 B.n265 B.n116 163.367
R372 B.n273 B.n116 163.367
R373 B.n274 B.n273 163.367
R374 B.n274 B.n5 163.367
R375 B.n6 B.n5 163.367
R376 B.n7 B.n6 163.367
R377 B.n279 B.n7 163.367
R378 B.n279 B.n12 163.367
R379 B.n13 B.n12 163.367
R380 B.n14 B.n13 163.367
R381 B.n284 B.n14 163.367
R382 B.n284 B.n19 163.367
R383 B.n20 B.n19 163.367
R384 B.n21 B.n20 163.367
R385 B.n289 B.n21 163.367
R386 B.n289 B.n26 163.367
R387 B.n27 B.n26 163.367
R388 B.n28 B.n27 163.367
R389 B.n49 B.n28 163.367
R390 B.n55 B.n32 163.367
R391 B.n59 B.n58 163.367
R392 B.n63 B.n62 163.367
R393 B.n67 B.n66 163.367
R394 B.n71 B.n70 163.367
R395 B.n75 B.n74 163.367
R396 B.n79 B.n78 163.367
R397 B.n83 B.n82 163.367
R398 B.n87 B.n86 163.367
R399 B.n91 B.n90 163.367
R400 B.n96 B.n95 163.367
R401 B.n100 B.n99 163.367
R402 B.n104 B.n103 163.367
R403 B.n108 B.n107 163.367
R404 B.n112 B.n111 163.367
R405 B.n296 B.n48 163.367
R406 B.n163 B.t15 142.607
R407 B.n50 B.t8 142.607
R408 B.n161 B.t5 142.607
R409 B.n52 B.t11 142.607
R410 B.n164 B.t14 120.498
R411 B.n51 B.t9 120.498
R412 B.n162 B.t4 120.498
R413 B.n53 B.t12 120.498
R414 B.n235 B.n141 104.543
R415 B.n235 B.n137 104.543
R416 B.n241 B.n137 104.543
R417 B.n241 B.n133 104.543
R418 B.n247 B.n133 104.543
R419 B.n253 B.n129 104.543
R420 B.n253 B.n125 104.543
R421 B.n259 B.n125 104.543
R422 B.n259 B.n121 104.543
R423 B.n266 B.n121 104.543
R424 B.n272 B.n117 104.543
R425 B.n272 B.n4 104.543
R426 B.n330 B.n4 104.543
R427 B.n330 B.n329 104.543
R428 B.n329 B.n328 104.543
R429 B.n328 B.n8 104.543
R430 B.n322 B.n321 104.543
R431 B.n321 B.n320 104.543
R432 B.n320 B.n15 104.543
R433 B.n314 B.n15 104.543
R434 B.n314 B.n313 104.543
R435 B.n312 B.n22 104.543
R436 B.n306 B.n22 104.543
R437 B.n306 B.n305 104.543
R438 B.n305 B.n304 104.543
R439 B.n304 B.n29 104.543
R440 B.t3 B.n129 87.6315
R441 B.n313 B.t7 87.6315
R442 B.n266 B.t1 75.3324
R443 B.n322 B.t0 75.3324
R444 B.n230 B.n229 71.676
R445 B.n160 B.n145 71.676
R446 B.n222 B.n146 71.676
R447 B.n218 B.n147 71.676
R448 B.n214 B.n148 71.676
R449 B.n210 B.n149 71.676
R450 B.n205 B.n150 71.676
R451 B.n201 B.n151 71.676
R452 B.n197 B.n152 71.676
R453 B.n193 B.n153 71.676
R454 B.n189 B.n154 71.676
R455 B.n185 B.n155 71.676
R456 B.n181 B.n156 71.676
R457 B.n177 B.n157 71.676
R458 B.n173 B.n158 71.676
R459 B.n169 B.n159 71.676
R460 B.n299 B.n298 71.676
R461 B.n55 B.n33 71.676
R462 B.n59 B.n34 71.676
R463 B.n63 B.n35 71.676
R464 B.n67 B.n36 71.676
R465 B.n71 B.n37 71.676
R466 B.n75 B.n38 71.676
R467 B.n79 B.n39 71.676
R468 B.n83 B.n40 71.676
R469 B.n87 B.n41 71.676
R470 B.n91 B.n42 71.676
R471 B.n96 B.n43 71.676
R472 B.n100 B.n44 71.676
R473 B.n104 B.n45 71.676
R474 B.n108 B.n46 71.676
R475 B.n112 B.n47 71.676
R476 B.n48 B.n47 71.676
R477 B.n111 B.n46 71.676
R478 B.n107 B.n45 71.676
R479 B.n103 B.n44 71.676
R480 B.n99 B.n43 71.676
R481 B.n95 B.n42 71.676
R482 B.n90 B.n41 71.676
R483 B.n86 B.n40 71.676
R484 B.n82 B.n39 71.676
R485 B.n78 B.n38 71.676
R486 B.n74 B.n37 71.676
R487 B.n70 B.n36 71.676
R488 B.n66 B.n35 71.676
R489 B.n62 B.n34 71.676
R490 B.n58 B.n33 71.676
R491 B.n298 B.n32 71.676
R492 B.n229 B.n144 71.676
R493 B.n223 B.n145 71.676
R494 B.n219 B.n146 71.676
R495 B.n215 B.n147 71.676
R496 B.n211 B.n148 71.676
R497 B.n206 B.n149 71.676
R498 B.n202 B.n150 71.676
R499 B.n198 B.n151 71.676
R500 B.n194 B.n152 71.676
R501 B.n190 B.n153 71.676
R502 B.n186 B.n154 71.676
R503 B.n182 B.n155 71.676
R504 B.n178 B.n156 71.676
R505 B.n174 B.n157 71.676
R506 B.n170 B.n158 71.676
R507 B.n166 B.n159 71.676
R508 B.n165 B.n164 59.5399
R509 B.n208 B.n162 59.5399
R510 B.n54 B.n53 59.5399
R511 B.n93 B.n51 59.5399
R512 B.n301 B.n300 32.0005
R513 B.n295 B.n294 32.0005
R514 B.n167 B.n139 32.0005
R515 B.n232 B.n231 32.0005
R516 B.t1 B.n117 29.2108
R517 B.t0 B.n8 29.2108
R518 B.n164 B.n163 22.1096
R519 B.n162 B.n161 22.1096
R520 B.n53 B.n52 22.1096
R521 B.n51 B.n50 22.1096
R522 B B.n332 18.0485
R523 B.n247 B.t3 16.9117
R524 B.t7 B.n312 16.9117
R525 B.n300 B.n31 10.6151
R526 B.n56 B.n31 10.6151
R527 B.n57 B.n56 10.6151
R528 B.n60 B.n57 10.6151
R529 B.n61 B.n60 10.6151
R530 B.n64 B.n61 10.6151
R531 B.n65 B.n64 10.6151
R532 B.n68 B.n65 10.6151
R533 B.n69 B.n68 10.6151
R534 B.n72 B.n69 10.6151
R535 B.n73 B.n72 10.6151
R536 B.n77 B.n76 10.6151
R537 B.n80 B.n77 10.6151
R538 B.n81 B.n80 10.6151
R539 B.n84 B.n81 10.6151
R540 B.n85 B.n84 10.6151
R541 B.n88 B.n85 10.6151
R542 B.n89 B.n88 10.6151
R543 B.n92 B.n89 10.6151
R544 B.n97 B.n94 10.6151
R545 B.n98 B.n97 10.6151
R546 B.n101 B.n98 10.6151
R547 B.n102 B.n101 10.6151
R548 B.n105 B.n102 10.6151
R549 B.n106 B.n105 10.6151
R550 B.n109 B.n106 10.6151
R551 B.n110 B.n109 10.6151
R552 B.n113 B.n110 10.6151
R553 B.n114 B.n113 10.6151
R554 B.n295 B.n114 10.6151
R555 B.n237 B.n139 10.6151
R556 B.n238 B.n237 10.6151
R557 B.n239 B.n238 10.6151
R558 B.n239 B.n131 10.6151
R559 B.n249 B.n131 10.6151
R560 B.n250 B.n249 10.6151
R561 B.n251 B.n250 10.6151
R562 B.n251 B.n123 10.6151
R563 B.n261 B.n123 10.6151
R564 B.n262 B.n261 10.6151
R565 B.n264 B.n262 10.6151
R566 B.n264 B.n263 10.6151
R567 B.n263 B.n115 10.6151
R568 B.n275 B.n115 10.6151
R569 B.n276 B.n275 10.6151
R570 B.n277 B.n276 10.6151
R571 B.n278 B.n277 10.6151
R572 B.n280 B.n278 10.6151
R573 B.n281 B.n280 10.6151
R574 B.n282 B.n281 10.6151
R575 B.n283 B.n282 10.6151
R576 B.n285 B.n283 10.6151
R577 B.n286 B.n285 10.6151
R578 B.n287 B.n286 10.6151
R579 B.n288 B.n287 10.6151
R580 B.n290 B.n288 10.6151
R581 B.n291 B.n290 10.6151
R582 B.n292 B.n291 10.6151
R583 B.n293 B.n292 10.6151
R584 B.n294 B.n293 10.6151
R585 B.n231 B.n143 10.6151
R586 B.n226 B.n143 10.6151
R587 B.n226 B.n225 10.6151
R588 B.n225 B.n224 10.6151
R589 B.n224 B.n221 10.6151
R590 B.n221 B.n220 10.6151
R591 B.n220 B.n217 10.6151
R592 B.n217 B.n216 10.6151
R593 B.n216 B.n213 10.6151
R594 B.n213 B.n212 10.6151
R595 B.n212 B.n209 10.6151
R596 B.n207 B.n204 10.6151
R597 B.n204 B.n203 10.6151
R598 B.n203 B.n200 10.6151
R599 B.n200 B.n199 10.6151
R600 B.n199 B.n196 10.6151
R601 B.n196 B.n195 10.6151
R602 B.n195 B.n192 10.6151
R603 B.n192 B.n191 10.6151
R604 B.n188 B.n187 10.6151
R605 B.n187 B.n184 10.6151
R606 B.n184 B.n183 10.6151
R607 B.n183 B.n180 10.6151
R608 B.n180 B.n179 10.6151
R609 B.n179 B.n176 10.6151
R610 B.n176 B.n175 10.6151
R611 B.n175 B.n172 10.6151
R612 B.n172 B.n171 10.6151
R613 B.n171 B.n168 10.6151
R614 B.n168 B.n167 10.6151
R615 B.n233 B.n232 10.6151
R616 B.n233 B.n135 10.6151
R617 B.n243 B.n135 10.6151
R618 B.n244 B.n243 10.6151
R619 B.n245 B.n244 10.6151
R620 B.n245 B.n127 10.6151
R621 B.n255 B.n127 10.6151
R622 B.n256 B.n255 10.6151
R623 B.n257 B.n256 10.6151
R624 B.n257 B.n119 10.6151
R625 B.n268 B.n119 10.6151
R626 B.n269 B.n268 10.6151
R627 B.n270 B.n269 10.6151
R628 B.n270 B.n0 10.6151
R629 B.n326 B.n1 10.6151
R630 B.n326 B.n325 10.6151
R631 B.n325 B.n324 10.6151
R632 B.n324 B.n10 10.6151
R633 B.n318 B.n10 10.6151
R634 B.n318 B.n317 10.6151
R635 B.n317 B.n316 10.6151
R636 B.n316 B.n17 10.6151
R637 B.n310 B.n17 10.6151
R638 B.n310 B.n309 10.6151
R639 B.n309 B.n308 10.6151
R640 B.n308 B.n24 10.6151
R641 B.n302 B.n24 10.6151
R642 B.n302 B.n301 10.6151
R643 B.n76 B.n54 7.02489
R644 B.n93 B.n92 7.02489
R645 B.n208 B.n207 7.02489
R646 B.n191 B.n165 7.02489
R647 B.n73 B.n54 3.59074
R648 B.n94 B.n93 3.59074
R649 B.n209 B.n208 3.59074
R650 B.n188 B.n165 3.59074
R651 B.n332 B.n0 2.81026
R652 B.n332 B.n1 2.81026
R653 VP.n0 VP.t1 297.976
R654 VP.n0 VP.t0 265.733
R655 VP VP.n0 0.0516364
R656 VDD1.n2 VDD1.n0 289.615
R657 VDD1.n9 VDD1.n7 289.615
R658 VDD1.n3 VDD1.n2 185
R659 VDD1.n10 VDD1.n9 185
R660 VDD1.t0 VDD1.n1 164.876
R661 VDD1.t1 VDD1.n8 164.876
R662 VDD1 VDD1.n13 80.3712
R663 VDD1 VDD1.n6 52.6589
R664 VDD1.n2 VDD1.t0 52.3082
R665 VDD1.n9 VDD1.t1 52.3082
R666 VDD1.n3 VDD1.n1 14.7318
R667 VDD1.n10 VDD1.n8 14.7318
R668 VDD1.n4 VDD1.n0 12.8005
R669 VDD1.n11 VDD1.n7 12.8005
R670 VDD1.n6 VDD1.n5 9.45567
R671 VDD1.n13 VDD1.n12 9.45567
R672 VDD1.n5 VDD1.n4 9.3005
R673 VDD1.n12 VDD1.n11 9.3005
R674 VDD1.n5 VDD1.n1 5.62509
R675 VDD1.n12 VDD1.n8 5.62509
R676 VDD1.n6 VDD1.n0 1.16414
R677 VDD1.n13 VDD1.n7 1.16414
R678 VDD1.n4 VDD1.n3 0.388379
R679 VDD1.n11 VDD1.n10 0.388379
C0 VP VDD2 0.264938f
C1 VN VP 2.74347f
C2 VDD1 VP 0.635849f
C3 VTAIL VP 0.597253f
C4 VN VDD2 0.527218f
C5 VDD1 VDD2 0.47019f
C6 VTAIL VDD2 1.96168f
C7 VDD1 VN 0.154794f
C8 VTAIL VN 0.583074f
C9 VDD1 VTAIL 1.92136f
C10 VDD2 B 1.89795f
C11 VDD1 B 2.03327f
C12 VTAIL B 2.29328f
C13 VN B 5.503769f
C14 VP B 3.329787f
C15 VP.t1 B 0.379108f
C16 VP.t0 B 0.264023f
C17 VP.n0 B 2.04029f
C18 VN.t1 B 0.258676f
C19 VN.t0 B 0.375446f
.ends

