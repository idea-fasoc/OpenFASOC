* NGSPICE file created from diff_pair_sample_1676.ext - technology: sky130A

.subckt diff_pair_sample_1676 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n4130_n3422# sky130_fd_pr__pfet_01v8 ad=4.7853 pd=25.32 as=0 ps=0 w=12.27 l=2.83
X1 VTAIL.t15 VP.t0 VDD1.t0 w_n4130_n3422# sky130_fd_pr__pfet_01v8 ad=2.02455 pd=12.6 as=2.02455 ps=12.6 w=12.27 l=2.83
X2 VTAIL.t7 VN.t0 VDD2.t7 w_n4130_n3422# sky130_fd_pr__pfet_01v8 ad=2.02455 pd=12.6 as=2.02455 ps=12.6 w=12.27 l=2.83
X3 B.t8 B.t6 B.t7 w_n4130_n3422# sky130_fd_pr__pfet_01v8 ad=4.7853 pd=25.32 as=0 ps=0 w=12.27 l=2.83
X4 VDD1.t4 VP.t1 VTAIL.t14 w_n4130_n3422# sky130_fd_pr__pfet_01v8 ad=2.02455 pd=12.6 as=2.02455 ps=12.6 w=12.27 l=2.83
X5 VDD2.t6 VN.t1 VTAIL.t4 w_n4130_n3422# sky130_fd_pr__pfet_01v8 ad=2.02455 pd=12.6 as=2.02455 ps=12.6 w=12.27 l=2.83
X6 VDD2.t5 VN.t2 VTAIL.t1 w_n4130_n3422# sky130_fd_pr__pfet_01v8 ad=2.02455 pd=12.6 as=4.7853 ps=25.32 w=12.27 l=2.83
X7 VTAIL.t6 VN.t3 VDD2.t4 w_n4130_n3422# sky130_fd_pr__pfet_01v8 ad=2.02455 pd=12.6 as=2.02455 ps=12.6 w=12.27 l=2.83
X8 VTAIL.t5 VN.t4 VDD2.t3 w_n4130_n3422# sky130_fd_pr__pfet_01v8 ad=4.7853 pd=25.32 as=2.02455 ps=12.6 w=12.27 l=2.83
X9 VDD1.t1 VP.t2 VTAIL.t13 w_n4130_n3422# sky130_fd_pr__pfet_01v8 ad=2.02455 pd=12.6 as=4.7853 ps=25.32 w=12.27 l=2.83
X10 VDD2.t2 VN.t5 VTAIL.t3 w_n4130_n3422# sky130_fd_pr__pfet_01v8 ad=2.02455 pd=12.6 as=2.02455 ps=12.6 w=12.27 l=2.83
X11 VTAIL.t12 VP.t3 VDD1.t2 w_n4130_n3422# sky130_fd_pr__pfet_01v8 ad=4.7853 pd=25.32 as=2.02455 ps=12.6 w=12.27 l=2.83
X12 VTAIL.t11 VP.t4 VDD1.t6 w_n4130_n3422# sky130_fd_pr__pfet_01v8 ad=2.02455 pd=12.6 as=2.02455 ps=12.6 w=12.27 l=2.83
X13 B.t5 B.t3 B.t4 w_n4130_n3422# sky130_fd_pr__pfet_01v8 ad=4.7853 pd=25.32 as=0 ps=0 w=12.27 l=2.83
X14 VDD2.t1 VN.t6 VTAIL.t2 w_n4130_n3422# sky130_fd_pr__pfet_01v8 ad=2.02455 pd=12.6 as=4.7853 ps=25.32 w=12.27 l=2.83
X15 VDD1.t5 VP.t5 VTAIL.t10 w_n4130_n3422# sky130_fd_pr__pfet_01v8 ad=2.02455 pd=12.6 as=4.7853 ps=25.32 w=12.27 l=2.83
X16 VTAIL.t0 VN.t7 VDD2.t0 w_n4130_n3422# sky130_fd_pr__pfet_01v8 ad=4.7853 pd=25.32 as=2.02455 ps=12.6 w=12.27 l=2.83
X17 VDD1.t7 VP.t6 VTAIL.t9 w_n4130_n3422# sky130_fd_pr__pfet_01v8 ad=2.02455 pd=12.6 as=2.02455 ps=12.6 w=12.27 l=2.83
X18 B.t2 B.t0 B.t1 w_n4130_n3422# sky130_fd_pr__pfet_01v8 ad=4.7853 pd=25.32 as=0 ps=0 w=12.27 l=2.83
X19 VTAIL.t8 VP.t7 VDD1.t3 w_n4130_n3422# sky130_fd_pr__pfet_01v8 ad=4.7853 pd=25.32 as=2.02455 ps=12.6 w=12.27 l=2.83
R0 B.n435 B.n434 585
R1 B.n433 B.n136 585
R2 B.n432 B.n431 585
R3 B.n430 B.n137 585
R4 B.n429 B.n428 585
R5 B.n427 B.n138 585
R6 B.n426 B.n425 585
R7 B.n424 B.n139 585
R8 B.n423 B.n422 585
R9 B.n421 B.n140 585
R10 B.n420 B.n419 585
R11 B.n418 B.n141 585
R12 B.n417 B.n416 585
R13 B.n415 B.n142 585
R14 B.n414 B.n413 585
R15 B.n412 B.n143 585
R16 B.n411 B.n410 585
R17 B.n409 B.n144 585
R18 B.n408 B.n407 585
R19 B.n406 B.n145 585
R20 B.n405 B.n404 585
R21 B.n403 B.n146 585
R22 B.n402 B.n401 585
R23 B.n400 B.n147 585
R24 B.n399 B.n398 585
R25 B.n397 B.n148 585
R26 B.n396 B.n395 585
R27 B.n394 B.n149 585
R28 B.n393 B.n392 585
R29 B.n391 B.n150 585
R30 B.n390 B.n389 585
R31 B.n388 B.n151 585
R32 B.n387 B.n386 585
R33 B.n385 B.n152 585
R34 B.n384 B.n383 585
R35 B.n382 B.n153 585
R36 B.n381 B.n380 585
R37 B.n379 B.n154 585
R38 B.n378 B.n377 585
R39 B.n376 B.n155 585
R40 B.n375 B.n374 585
R41 B.n373 B.n156 585
R42 B.n372 B.n371 585
R43 B.n367 B.n157 585
R44 B.n366 B.n365 585
R45 B.n364 B.n158 585
R46 B.n363 B.n362 585
R47 B.n361 B.n159 585
R48 B.n360 B.n359 585
R49 B.n358 B.n160 585
R50 B.n357 B.n356 585
R51 B.n355 B.n161 585
R52 B.n353 B.n352 585
R53 B.n351 B.n164 585
R54 B.n350 B.n349 585
R55 B.n348 B.n165 585
R56 B.n347 B.n346 585
R57 B.n345 B.n166 585
R58 B.n344 B.n343 585
R59 B.n342 B.n167 585
R60 B.n341 B.n340 585
R61 B.n339 B.n168 585
R62 B.n338 B.n337 585
R63 B.n336 B.n169 585
R64 B.n335 B.n334 585
R65 B.n333 B.n170 585
R66 B.n332 B.n331 585
R67 B.n330 B.n171 585
R68 B.n329 B.n328 585
R69 B.n327 B.n172 585
R70 B.n326 B.n325 585
R71 B.n324 B.n173 585
R72 B.n323 B.n322 585
R73 B.n321 B.n174 585
R74 B.n320 B.n319 585
R75 B.n318 B.n175 585
R76 B.n317 B.n316 585
R77 B.n315 B.n176 585
R78 B.n314 B.n313 585
R79 B.n312 B.n177 585
R80 B.n311 B.n310 585
R81 B.n309 B.n178 585
R82 B.n308 B.n307 585
R83 B.n306 B.n179 585
R84 B.n305 B.n304 585
R85 B.n303 B.n180 585
R86 B.n302 B.n301 585
R87 B.n300 B.n181 585
R88 B.n299 B.n298 585
R89 B.n297 B.n182 585
R90 B.n296 B.n295 585
R91 B.n294 B.n183 585
R92 B.n293 B.n292 585
R93 B.n291 B.n184 585
R94 B.n436 B.n135 585
R95 B.n438 B.n437 585
R96 B.n439 B.n134 585
R97 B.n441 B.n440 585
R98 B.n442 B.n133 585
R99 B.n444 B.n443 585
R100 B.n445 B.n132 585
R101 B.n447 B.n446 585
R102 B.n448 B.n131 585
R103 B.n450 B.n449 585
R104 B.n451 B.n130 585
R105 B.n453 B.n452 585
R106 B.n454 B.n129 585
R107 B.n456 B.n455 585
R108 B.n457 B.n128 585
R109 B.n459 B.n458 585
R110 B.n460 B.n127 585
R111 B.n462 B.n461 585
R112 B.n463 B.n126 585
R113 B.n465 B.n464 585
R114 B.n466 B.n125 585
R115 B.n468 B.n467 585
R116 B.n469 B.n124 585
R117 B.n471 B.n470 585
R118 B.n472 B.n123 585
R119 B.n474 B.n473 585
R120 B.n475 B.n122 585
R121 B.n477 B.n476 585
R122 B.n478 B.n121 585
R123 B.n480 B.n479 585
R124 B.n481 B.n120 585
R125 B.n483 B.n482 585
R126 B.n484 B.n119 585
R127 B.n486 B.n485 585
R128 B.n487 B.n118 585
R129 B.n489 B.n488 585
R130 B.n490 B.n117 585
R131 B.n492 B.n491 585
R132 B.n493 B.n116 585
R133 B.n495 B.n494 585
R134 B.n496 B.n115 585
R135 B.n498 B.n497 585
R136 B.n499 B.n114 585
R137 B.n501 B.n500 585
R138 B.n502 B.n113 585
R139 B.n504 B.n503 585
R140 B.n505 B.n112 585
R141 B.n507 B.n506 585
R142 B.n508 B.n111 585
R143 B.n510 B.n509 585
R144 B.n511 B.n110 585
R145 B.n513 B.n512 585
R146 B.n514 B.n109 585
R147 B.n516 B.n515 585
R148 B.n517 B.n108 585
R149 B.n519 B.n518 585
R150 B.n520 B.n107 585
R151 B.n522 B.n521 585
R152 B.n523 B.n106 585
R153 B.n525 B.n524 585
R154 B.n526 B.n105 585
R155 B.n528 B.n527 585
R156 B.n529 B.n104 585
R157 B.n531 B.n530 585
R158 B.n532 B.n103 585
R159 B.n534 B.n533 585
R160 B.n535 B.n102 585
R161 B.n537 B.n536 585
R162 B.n538 B.n101 585
R163 B.n540 B.n539 585
R164 B.n541 B.n100 585
R165 B.n543 B.n542 585
R166 B.n544 B.n99 585
R167 B.n546 B.n545 585
R168 B.n547 B.n98 585
R169 B.n549 B.n548 585
R170 B.n550 B.n97 585
R171 B.n552 B.n551 585
R172 B.n553 B.n96 585
R173 B.n555 B.n554 585
R174 B.n556 B.n95 585
R175 B.n558 B.n557 585
R176 B.n559 B.n94 585
R177 B.n561 B.n560 585
R178 B.n562 B.n93 585
R179 B.n564 B.n563 585
R180 B.n565 B.n92 585
R181 B.n567 B.n566 585
R182 B.n568 B.n91 585
R183 B.n570 B.n569 585
R184 B.n571 B.n90 585
R185 B.n573 B.n572 585
R186 B.n574 B.n89 585
R187 B.n576 B.n575 585
R188 B.n577 B.n88 585
R189 B.n579 B.n578 585
R190 B.n580 B.n87 585
R191 B.n582 B.n581 585
R192 B.n583 B.n86 585
R193 B.n585 B.n584 585
R194 B.n586 B.n85 585
R195 B.n588 B.n587 585
R196 B.n589 B.n84 585
R197 B.n591 B.n590 585
R198 B.n592 B.n83 585
R199 B.n594 B.n593 585
R200 B.n595 B.n82 585
R201 B.n597 B.n596 585
R202 B.n598 B.n81 585
R203 B.n600 B.n599 585
R204 B.n742 B.n29 585
R205 B.n741 B.n740 585
R206 B.n739 B.n30 585
R207 B.n738 B.n737 585
R208 B.n736 B.n31 585
R209 B.n735 B.n734 585
R210 B.n733 B.n32 585
R211 B.n732 B.n731 585
R212 B.n730 B.n33 585
R213 B.n729 B.n728 585
R214 B.n727 B.n34 585
R215 B.n726 B.n725 585
R216 B.n724 B.n35 585
R217 B.n723 B.n722 585
R218 B.n721 B.n36 585
R219 B.n720 B.n719 585
R220 B.n718 B.n37 585
R221 B.n717 B.n716 585
R222 B.n715 B.n38 585
R223 B.n714 B.n713 585
R224 B.n712 B.n39 585
R225 B.n711 B.n710 585
R226 B.n709 B.n40 585
R227 B.n708 B.n707 585
R228 B.n706 B.n41 585
R229 B.n705 B.n704 585
R230 B.n703 B.n42 585
R231 B.n702 B.n701 585
R232 B.n700 B.n43 585
R233 B.n699 B.n698 585
R234 B.n697 B.n44 585
R235 B.n696 B.n695 585
R236 B.n694 B.n45 585
R237 B.n693 B.n692 585
R238 B.n691 B.n46 585
R239 B.n690 B.n689 585
R240 B.n688 B.n47 585
R241 B.n687 B.n686 585
R242 B.n685 B.n48 585
R243 B.n684 B.n683 585
R244 B.n682 B.n49 585
R245 B.n681 B.n680 585
R246 B.n679 B.n678 585
R247 B.n677 B.n53 585
R248 B.n676 B.n675 585
R249 B.n674 B.n54 585
R250 B.n673 B.n672 585
R251 B.n671 B.n55 585
R252 B.n670 B.n669 585
R253 B.n668 B.n56 585
R254 B.n667 B.n666 585
R255 B.n665 B.n57 585
R256 B.n663 B.n662 585
R257 B.n661 B.n60 585
R258 B.n660 B.n659 585
R259 B.n658 B.n61 585
R260 B.n657 B.n656 585
R261 B.n655 B.n62 585
R262 B.n654 B.n653 585
R263 B.n652 B.n63 585
R264 B.n651 B.n650 585
R265 B.n649 B.n64 585
R266 B.n648 B.n647 585
R267 B.n646 B.n65 585
R268 B.n645 B.n644 585
R269 B.n643 B.n66 585
R270 B.n642 B.n641 585
R271 B.n640 B.n67 585
R272 B.n639 B.n638 585
R273 B.n637 B.n68 585
R274 B.n636 B.n635 585
R275 B.n634 B.n69 585
R276 B.n633 B.n632 585
R277 B.n631 B.n70 585
R278 B.n630 B.n629 585
R279 B.n628 B.n71 585
R280 B.n627 B.n626 585
R281 B.n625 B.n72 585
R282 B.n624 B.n623 585
R283 B.n622 B.n73 585
R284 B.n621 B.n620 585
R285 B.n619 B.n74 585
R286 B.n618 B.n617 585
R287 B.n616 B.n75 585
R288 B.n615 B.n614 585
R289 B.n613 B.n76 585
R290 B.n612 B.n611 585
R291 B.n610 B.n77 585
R292 B.n609 B.n608 585
R293 B.n607 B.n78 585
R294 B.n606 B.n605 585
R295 B.n604 B.n79 585
R296 B.n603 B.n602 585
R297 B.n601 B.n80 585
R298 B.n744 B.n743 585
R299 B.n745 B.n28 585
R300 B.n747 B.n746 585
R301 B.n748 B.n27 585
R302 B.n750 B.n749 585
R303 B.n751 B.n26 585
R304 B.n753 B.n752 585
R305 B.n754 B.n25 585
R306 B.n756 B.n755 585
R307 B.n757 B.n24 585
R308 B.n759 B.n758 585
R309 B.n760 B.n23 585
R310 B.n762 B.n761 585
R311 B.n763 B.n22 585
R312 B.n765 B.n764 585
R313 B.n766 B.n21 585
R314 B.n768 B.n767 585
R315 B.n769 B.n20 585
R316 B.n771 B.n770 585
R317 B.n772 B.n19 585
R318 B.n774 B.n773 585
R319 B.n775 B.n18 585
R320 B.n777 B.n776 585
R321 B.n778 B.n17 585
R322 B.n780 B.n779 585
R323 B.n781 B.n16 585
R324 B.n783 B.n782 585
R325 B.n784 B.n15 585
R326 B.n786 B.n785 585
R327 B.n787 B.n14 585
R328 B.n789 B.n788 585
R329 B.n790 B.n13 585
R330 B.n792 B.n791 585
R331 B.n793 B.n12 585
R332 B.n795 B.n794 585
R333 B.n796 B.n11 585
R334 B.n798 B.n797 585
R335 B.n799 B.n10 585
R336 B.n801 B.n800 585
R337 B.n802 B.n9 585
R338 B.n804 B.n803 585
R339 B.n805 B.n8 585
R340 B.n807 B.n806 585
R341 B.n808 B.n7 585
R342 B.n810 B.n809 585
R343 B.n811 B.n6 585
R344 B.n813 B.n812 585
R345 B.n814 B.n5 585
R346 B.n816 B.n815 585
R347 B.n817 B.n4 585
R348 B.n819 B.n818 585
R349 B.n820 B.n3 585
R350 B.n822 B.n821 585
R351 B.n823 B.n0 585
R352 B.n2 B.n1 585
R353 B.n212 B.n211 585
R354 B.n213 B.n210 585
R355 B.n215 B.n214 585
R356 B.n216 B.n209 585
R357 B.n218 B.n217 585
R358 B.n219 B.n208 585
R359 B.n221 B.n220 585
R360 B.n222 B.n207 585
R361 B.n224 B.n223 585
R362 B.n225 B.n206 585
R363 B.n227 B.n226 585
R364 B.n228 B.n205 585
R365 B.n230 B.n229 585
R366 B.n231 B.n204 585
R367 B.n233 B.n232 585
R368 B.n234 B.n203 585
R369 B.n236 B.n235 585
R370 B.n237 B.n202 585
R371 B.n239 B.n238 585
R372 B.n240 B.n201 585
R373 B.n242 B.n241 585
R374 B.n243 B.n200 585
R375 B.n245 B.n244 585
R376 B.n246 B.n199 585
R377 B.n248 B.n247 585
R378 B.n249 B.n198 585
R379 B.n251 B.n250 585
R380 B.n252 B.n197 585
R381 B.n254 B.n253 585
R382 B.n255 B.n196 585
R383 B.n257 B.n256 585
R384 B.n258 B.n195 585
R385 B.n260 B.n259 585
R386 B.n261 B.n194 585
R387 B.n263 B.n262 585
R388 B.n264 B.n193 585
R389 B.n266 B.n265 585
R390 B.n267 B.n192 585
R391 B.n269 B.n268 585
R392 B.n270 B.n191 585
R393 B.n272 B.n271 585
R394 B.n273 B.n190 585
R395 B.n275 B.n274 585
R396 B.n276 B.n189 585
R397 B.n278 B.n277 585
R398 B.n279 B.n188 585
R399 B.n281 B.n280 585
R400 B.n282 B.n187 585
R401 B.n284 B.n283 585
R402 B.n285 B.n186 585
R403 B.n287 B.n286 585
R404 B.n288 B.n185 585
R405 B.n290 B.n289 585
R406 B.n291 B.n290 545.355
R407 B.n434 B.n135 545.355
R408 B.n601 B.n600 545.355
R409 B.n744 B.n29 545.355
R410 B.n162 B.t0 312.86
R411 B.n368 B.t3 312.86
R412 B.n58 B.t9 312.86
R413 B.n50 B.t6 312.86
R414 B.n825 B.n824 256.663
R415 B.n824 B.n823 235.042
R416 B.n824 B.n2 235.042
R417 B.n368 B.t4 168.911
R418 B.n58 B.t11 168.911
R419 B.n162 B.t1 168.895
R420 B.n50 B.t8 168.895
R421 B.n292 B.n291 163.367
R422 B.n292 B.n183 163.367
R423 B.n296 B.n183 163.367
R424 B.n297 B.n296 163.367
R425 B.n298 B.n297 163.367
R426 B.n298 B.n181 163.367
R427 B.n302 B.n181 163.367
R428 B.n303 B.n302 163.367
R429 B.n304 B.n303 163.367
R430 B.n304 B.n179 163.367
R431 B.n308 B.n179 163.367
R432 B.n309 B.n308 163.367
R433 B.n310 B.n309 163.367
R434 B.n310 B.n177 163.367
R435 B.n314 B.n177 163.367
R436 B.n315 B.n314 163.367
R437 B.n316 B.n315 163.367
R438 B.n316 B.n175 163.367
R439 B.n320 B.n175 163.367
R440 B.n321 B.n320 163.367
R441 B.n322 B.n321 163.367
R442 B.n322 B.n173 163.367
R443 B.n326 B.n173 163.367
R444 B.n327 B.n326 163.367
R445 B.n328 B.n327 163.367
R446 B.n328 B.n171 163.367
R447 B.n332 B.n171 163.367
R448 B.n333 B.n332 163.367
R449 B.n334 B.n333 163.367
R450 B.n334 B.n169 163.367
R451 B.n338 B.n169 163.367
R452 B.n339 B.n338 163.367
R453 B.n340 B.n339 163.367
R454 B.n340 B.n167 163.367
R455 B.n344 B.n167 163.367
R456 B.n345 B.n344 163.367
R457 B.n346 B.n345 163.367
R458 B.n346 B.n165 163.367
R459 B.n350 B.n165 163.367
R460 B.n351 B.n350 163.367
R461 B.n352 B.n351 163.367
R462 B.n352 B.n161 163.367
R463 B.n357 B.n161 163.367
R464 B.n358 B.n357 163.367
R465 B.n359 B.n358 163.367
R466 B.n359 B.n159 163.367
R467 B.n363 B.n159 163.367
R468 B.n364 B.n363 163.367
R469 B.n365 B.n364 163.367
R470 B.n365 B.n157 163.367
R471 B.n372 B.n157 163.367
R472 B.n373 B.n372 163.367
R473 B.n374 B.n373 163.367
R474 B.n374 B.n155 163.367
R475 B.n378 B.n155 163.367
R476 B.n379 B.n378 163.367
R477 B.n380 B.n379 163.367
R478 B.n380 B.n153 163.367
R479 B.n384 B.n153 163.367
R480 B.n385 B.n384 163.367
R481 B.n386 B.n385 163.367
R482 B.n386 B.n151 163.367
R483 B.n390 B.n151 163.367
R484 B.n391 B.n390 163.367
R485 B.n392 B.n391 163.367
R486 B.n392 B.n149 163.367
R487 B.n396 B.n149 163.367
R488 B.n397 B.n396 163.367
R489 B.n398 B.n397 163.367
R490 B.n398 B.n147 163.367
R491 B.n402 B.n147 163.367
R492 B.n403 B.n402 163.367
R493 B.n404 B.n403 163.367
R494 B.n404 B.n145 163.367
R495 B.n408 B.n145 163.367
R496 B.n409 B.n408 163.367
R497 B.n410 B.n409 163.367
R498 B.n410 B.n143 163.367
R499 B.n414 B.n143 163.367
R500 B.n415 B.n414 163.367
R501 B.n416 B.n415 163.367
R502 B.n416 B.n141 163.367
R503 B.n420 B.n141 163.367
R504 B.n421 B.n420 163.367
R505 B.n422 B.n421 163.367
R506 B.n422 B.n139 163.367
R507 B.n426 B.n139 163.367
R508 B.n427 B.n426 163.367
R509 B.n428 B.n427 163.367
R510 B.n428 B.n137 163.367
R511 B.n432 B.n137 163.367
R512 B.n433 B.n432 163.367
R513 B.n434 B.n433 163.367
R514 B.n600 B.n81 163.367
R515 B.n596 B.n81 163.367
R516 B.n596 B.n595 163.367
R517 B.n595 B.n594 163.367
R518 B.n594 B.n83 163.367
R519 B.n590 B.n83 163.367
R520 B.n590 B.n589 163.367
R521 B.n589 B.n588 163.367
R522 B.n588 B.n85 163.367
R523 B.n584 B.n85 163.367
R524 B.n584 B.n583 163.367
R525 B.n583 B.n582 163.367
R526 B.n582 B.n87 163.367
R527 B.n578 B.n87 163.367
R528 B.n578 B.n577 163.367
R529 B.n577 B.n576 163.367
R530 B.n576 B.n89 163.367
R531 B.n572 B.n89 163.367
R532 B.n572 B.n571 163.367
R533 B.n571 B.n570 163.367
R534 B.n570 B.n91 163.367
R535 B.n566 B.n91 163.367
R536 B.n566 B.n565 163.367
R537 B.n565 B.n564 163.367
R538 B.n564 B.n93 163.367
R539 B.n560 B.n93 163.367
R540 B.n560 B.n559 163.367
R541 B.n559 B.n558 163.367
R542 B.n558 B.n95 163.367
R543 B.n554 B.n95 163.367
R544 B.n554 B.n553 163.367
R545 B.n553 B.n552 163.367
R546 B.n552 B.n97 163.367
R547 B.n548 B.n97 163.367
R548 B.n548 B.n547 163.367
R549 B.n547 B.n546 163.367
R550 B.n546 B.n99 163.367
R551 B.n542 B.n99 163.367
R552 B.n542 B.n541 163.367
R553 B.n541 B.n540 163.367
R554 B.n540 B.n101 163.367
R555 B.n536 B.n101 163.367
R556 B.n536 B.n535 163.367
R557 B.n535 B.n534 163.367
R558 B.n534 B.n103 163.367
R559 B.n530 B.n103 163.367
R560 B.n530 B.n529 163.367
R561 B.n529 B.n528 163.367
R562 B.n528 B.n105 163.367
R563 B.n524 B.n105 163.367
R564 B.n524 B.n523 163.367
R565 B.n523 B.n522 163.367
R566 B.n522 B.n107 163.367
R567 B.n518 B.n107 163.367
R568 B.n518 B.n517 163.367
R569 B.n517 B.n516 163.367
R570 B.n516 B.n109 163.367
R571 B.n512 B.n109 163.367
R572 B.n512 B.n511 163.367
R573 B.n511 B.n510 163.367
R574 B.n510 B.n111 163.367
R575 B.n506 B.n111 163.367
R576 B.n506 B.n505 163.367
R577 B.n505 B.n504 163.367
R578 B.n504 B.n113 163.367
R579 B.n500 B.n113 163.367
R580 B.n500 B.n499 163.367
R581 B.n499 B.n498 163.367
R582 B.n498 B.n115 163.367
R583 B.n494 B.n115 163.367
R584 B.n494 B.n493 163.367
R585 B.n493 B.n492 163.367
R586 B.n492 B.n117 163.367
R587 B.n488 B.n117 163.367
R588 B.n488 B.n487 163.367
R589 B.n487 B.n486 163.367
R590 B.n486 B.n119 163.367
R591 B.n482 B.n119 163.367
R592 B.n482 B.n481 163.367
R593 B.n481 B.n480 163.367
R594 B.n480 B.n121 163.367
R595 B.n476 B.n121 163.367
R596 B.n476 B.n475 163.367
R597 B.n475 B.n474 163.367
R598 B.n474 B.n123 163.367
R599 B.n470 B.n123 163.367
R600 B.n470 B.n469 163.367
R601 B.n469 B.n468 163.367
R602 B.n468 B.n125 163.367
R603 B.n464 B.n125 163.367
R604 B.n464 B.n463 163.367
R605 B.n463 B.n462 163.367
R606 B.n462 B.n127 163.367
R607 B.n458 B.n127 163.367
R608 B.n458 B.n457 163.367
R609 B.n457 B.n456 163.367
R610 B.n456 B.n129 163.367
R611 B.n452 B.n129 163.367
R612 B.n452 B.n451 163.367
R613 B.n451 B.n450 163.367
R614 B.n450 B.n131 163.367
R615 B.n446 B.n131 163.367
R616 B.n446 B.n445 163.367
R617 B.n445 B.n444 163.367
R618 B.n444 B.n133 163.367
R619 B.n440 B.n133 163.367
R620 B.n440 B.n439 163.367
R621 B.n439 B.n438 163.367
R622 B.n438 B.n135 163.367
R623 B.n740 B.n29 163.367
R624 B.n740 B.n739 163.367
R625 B.n739 B.n738 163.367
R626 B.n738 B.n31 163.367
R627 B.n734 B.n31 163.367
R628 B.n734 B.n733 163.367
R629 B.n733 B.n732 163.367
R630 B.n732 B.n33 163.367
R631 B.n728 B.n33 163.367
R632 B.n728 B.n727 163.367
R633 B.n727 B.n726 163.367
R634 B.n726 B.n35 163.367
R635 B.n722 B.n35 163.367
R636 B.n722 B.n721 163.367
R637 B.n721 B.n720 163.367
R638 B.n720 B.n37 163.367
R639 B.n716 B.n37 163.367
R640 B.n716 B.n715 163.367
R641 B.n715 B.n714 163.367
R642 B.n714 B.n39 163.367
R643 B.n710 B.n39 163.367
R644 B.n710 B.n709 163.367
R645 B.n709 B.n708 163.367
R646 B.n708 B.n41 163.367
R647 B.n704 B.n41 163.367
R648 B.n704 B.n703 163.367
R649 B.n703 B.n702 163.367
R650 B.n702 B.n43 163.367
R651 B.n698 B.n43 163.367
R652 B.n698 B.n697 163.367
R653 B.n697 B.n696 163.367
R654 B.n696 B.n45 163.367
R655 B.n692 B.n45 163.367
R656 B.n692 B.n691 163.367
R657 B.n691 B.n690 163.367
R658 B.n690 B.n47 163.367
R659 B.n686 B.n47 163.367
R660 B.n686 B.n685 163.367
R661 B.n685 B.n684 163.367
R662 B.n684 B.n49 163.367
R663 B.n680 B.n49 163.367
R664 B.n680 B.n679 163.367
R665 B.n679 B.n53 163.367
R666 B.n675 B.n53 163.367
R667 B.n675 B.n674 163.367
R668 B.n674 B.n673 163.367
R669 B.n673 B.n55 163.367
R670 B.n669 B.n55 163.367
R671 B.n669 B.n668 163.367
R672 B.n668 B.n667 163.367
R673 B.n667 B.n57 163.367
R674 B.n662 B.n57 163.367
R675 B.n662 B.n661 163.367
R676 B.n661 B.n660 163.367
R677 B.n660 B.n61 163.367
R678 B.n656 B.n61 163.367
R679 B.n656 B.n655 163.367
R680 B.n655 B.n654 163.367
R681 B.n654 B.n63 163.367
R682 B.n650 B.n63 163.367
R683 B.n650 B.n649 163.367
R684 B.n649 B.n648 163.367
R685 B.n648 B.n65 163.367
R686 B.n644 B.n65 163.367
R687 B.n644 B.n643 163.367
R688 B.n643 B.n642 163.367
R689 B.n642 B.n67 163.367
R690 B.n638 B.n67 163.367
R691 B.n638 B.n637 163.367
R692 B.n637 B.n636 163.367
R693 B.n636 B.n69 163.367
R694 B.n632 B.n69 163.367
R695 B.n632 B.n631 163.367
R696 B.n631 B.n630 163.367
R697 B.n630 B.n71 163.367
R698 B.n626 B.n71 163.367
R699 B.n626 B.n625 163.367
R700 B.n625 B.n624 163.367
R701 B.n624 B.n73 163.367
R702 B.n620 B.n73 163.367
R703 B.n620 B.n619 163.367
R704 B.n619 B.n618 163.367
R705 B.n618 B.n75 163.367
R706 B.n614 B.n75 163.367
R707 B.n614 B.n613 163.367
R708 B.n613 B.n612 163.367
R709 B.n612 B.n77 163.367
R710 B.n608 B.n77 163.367
R711 B.n608 B.n607 163.367
R712 B.n607 B.n606 163.367
R713 B.n606 B.n79 163.367
R714 B.n602 B.n79 163.367
R715 B.n602 B.n601 163.367
R716 B.n745 B.n744 163.367
R717 B.n746 B.n745 163.367
R718 B.n746 B.n27 163.367
R719 B.n750 B.n27 163.367
R720 B.n751 B.n750 163.367
R721 B.n752 B.n751 163.367
R722 B.n752 B.n25 163.367
R723 B.n756 B.n25 163.367
R724 B.n757 B.n756 163.367
R725 B.n758 B.n757 163.367
R726 B.n758 B.n23 163.367
R727 B.n762 B.n23 163.367
R728 B.n763 B.n762 163.367
R729 B.n764 B.n763 163.367
R730 B.n764 B.n21 163.367
R731 B.n768 B.n21 163.367
R732 B.n769 B.n768 163.367
R733 B.n770 B.n769 163.367
R734 B.n770 B.n19 163.367
R735 B.n774 B.n19 163.367
R736 B.n775 B.n774 163.367
R737 B.n776 B.n775 163.367
R738 B.n776 B.n17 163.367
R739 B.n780 B.n17 163.367
R740 B.n781 B.n780 163.367
R741 B.n782 B.n781 163.367
R742 B.n782 B.n15 163.367
R743 B.n786 B.n15 163.367
R744 B.n787 B.n786 163.367
R745 B.n788 B.n787 163.367
R746 B.n788 B.n13 163.367
R747 B.n792 B.n13 163.367
R748 B.n793 B.n792 163.367
R749 B.n794 B.n793 163.367
R750 B.n794 B.n11 163.367
R751 B.n798 B.n11 163.367
R752 B.n799 B.n798 163.367
R753 B.n800 B.n799 163.367
R754 B.n800 B.n9 163.367
R755 B.n804 B.n9 163.367
R756 B.n805 B.n804 163.367
R757 B.n806 B.n805 163.367
R758 B.n806 B.n7 163.367
R759 B.n810 B.n7 163.367
R760 B.n811 B.n810 163.367
R761 B.n812 B.n811 163.367
R762 B.n812 B.n5 163.367
R763 B.n816 B.n5 163.367
R764 B.n817 B.n816 163.367
R765 B.n818 B.n817 163.367
R766 B.n818 B.n3 163.367
R767 B.n822 B.n3 163.367
R768 B.n823 B.n822 163.367
R769 B.n212 B.n2 163.367
R770 B.n213 B.n212 163.367
R771 B.n214 B.n213 163.367
R772 B.n214 B.n209 163.367
R773 B.n218 B.n209 163.367
R774 B.n219 B.n218 163.367
R775 B.n220 B.n219 163.367
R776 B.n220 B.n207 163.367
R777 B.n224 B.n207 163.367
R778 B.n225 B.n224 163.367
R779 B.n226 B.n225 163.367
R780 B.n226 B.n205 163.367
R781 B.n230 B.n205 163.367
R782 B.n231 B.n230 163.367
R783 B.n232 B.n231 163.367
R784 B.n232 B.n203 163.367
R785 B.n236 B.n203 163.367
R786 B.n237 B.n236 163.367
R787 B.n238 B.n237 163.367
R788 B.n238 B.n201 163.367
R789 B.n242 B.n201 163.367
R790 B.n243 B.n242 163.367
R791 B.n244 B.n243 163.367
R792 B.n244 B.n199 163.367
R793 B.n248 B.n199 163.367
R794 B.n249 B.n248 163.367
R795 B.n250 B.n249 163.367
R796 B.n250 B.n197 163.367
R797 B.n254 B.n197 163.367
R798 B.n255 B.n254 163.367
R799 B.n256 B.n255 163.367
R800 B.n256 B.n195 163.367
R801 B.n260 B.n195 163.367
R802 B.n261 B.n260 163.367
R803 B.n262 B.n261 163.367
R804 B.n262 B.n193 163.367
R805 B.n266 B.n193 163.367
R806 B.n267 B.n266 163.367
R807 B.n268 B.n267 163.367
R808 B.n268 B.n191 163.367
R809 B.n272 B.n191 163.367
R810 B.n273 B.n272 163.367
R811 B.n274 B.n273 163.367
R812 B.n274 B.n189 163.367
R813 B.n278 B.n189 163.367
R814 B.n279 B.n278 163.367
R815 B.n280 B.n279 163.367
R816 B.n280 B.n187 163.367
R817 B.n284 B.n187 163.367
R818 B.n285 B.n284 163.367
R819 B.n286 B.n285 163.367
R820 B.n286 B.n185 163.367
R821 B.n290 B.n185 163.367
R822 B.n369 B.t5 107.626
R823 B.n59 B.t10 107.626
R824 B.n163 B.t2 107.611
R825 B.n51 B.t7 107.611
R826 B.n163 B.n162 61.2853
R827 B.n369 B.n368 61.2853
R828 B.n59 B.n58 61.2853
R829 B.n51 B.n50 61.2853
R830 B.n354 B.n163 59.5399
R831 B.n370 B.n369 59.5399
R832 B.n664 B.n59 59.5399
R833 B.n52 B.n51 59.5399
R834 B.n743 B.n742 35.4346
R835 B.n599 B.n80 35.4346
R836 B.n289 B.n184 35.4346
R837 B.n436 B.n435 35.4346
R838 B B.n825 18.0485
R839 B.n743 B.n28 10.6151
R840 B.n747 B.n28 10.6151
R841 B.n748 B.n747 10.6151
R842 B.n749 B.n748 10.6151
R843 B.n749 B.n26 10.6151
R844 B.n753 B.n26 10.6151
R845 B.n754 B.n753 10.6151
R846 B.n755 B.n754 10.6151
R847 B.n755 B.n24 10.6151
R848 B.n759 B.n24 10.6151
R849 B.n760 B.n759 10.6151
R850 B.n761 B.n760 10.6151
R851 B.n761 B.n22 10.6151
R852 B.n765 B.n22 10.6151
R853 B.n766 B.n765 10.6151
R854 B.n767 B.n766 10.6151
R855 B.n767 B.n20 10.6151
R856 B.n771 B.n20 10.6151
R857 B.n772 B.n771 10.6151
R858 B.n773 B.n772 10.6151
R859 B.n773 B.n18 10.6151
R860 B.n777 B.n18 10.6151
R861 B.n778 B.n777 10.6151
R862 B.n779 B.n778 10.6151
R863 B.n779 B.n16 10.6151
R864 B.n783 B.n16 10.6151
R865 B.n784 B.n783 10.6151
R866 B.n785 B.n784 10.6151
R867 B.n785 B.n14 10.6151
R868 B.n789 B.n14 10.6151
R869 B.n790 B.n789 10.6151
R870 B.n791 B.n790 10.6151
R871 B.n791 B.n12 10.6151
R872 B.n795 B.n12 10.6151
R873 B.n796 B.n795 10.6151
R874 B.n797 B.n796 10.6151
R875 B.n797 B.n10 10.6151
R876 B.n801 B.n10 10.6151
R877 B.n802 B.n801 10.6151
R878 B.n803 B.n802 10.6151
R879 B.n803 B.n8 10.6151
R880 B.n807 B.n8 10.6151
R881 B.n808 B.n807 10.6151
R882 B.n809 B.n808 10.6151
R883 B.n809 B.n6 10.6151
R884 B.n813 B.n6 10.6151
R885 B.n814 B.n813 10.6151
R886 B.n815 B.n814 10.6151
R887 B.n815 B.n4 10.6151
R888 B.n819 B.n4 10.6151
R889 B.n820 B.n819 10.6151
R890 B.n821 B.n820 10.6151
R891 B.n821 B.n0 10.6151
R892 B.n742 B.n741 10.6151
R893 B.n741 B.n30 10.6151
R894 B.n737 B.n30 10.6151
R895 B.n737 B.n736 10.6151
R896 B.n736 B.n735 10.6151
R897 B.n735 B.n32 10.6151
R898 B.n731 B.n32 10.6151
R899 B.n731 B.n730 10.6151
R900 B.n730 B.n729 10.6151
R901 B.n729 B.n34 10.6151
R902 B.n725 B.n34 10.6151
R903 B.n725 B.n724 10.6151
R904 B.n724 B.n723 10.6151
R905 B.n723 B.n36 10.6151
R906 B.n719 B.n36 10.6151
R907 B.n719 B.n718 10.6151
R908 B.n718 B.n717 10.6151
R909 B.n717 B.n38 10.6151
R910 B.n713 B.n38 10.6151
R911 B.n713 B.n712 10.6151
R912 B.n712 B.n711 10.6151
R913 B.n711 B.n40 10.6151
R914 B.n707 B.n40 10.6151
R915 B.n707 B.n706 10.6151
R916 B.n706 B.n705 10.6151
R917 B.n705 B.n42 10.6151
R918 B.n701 B.n42 10.6151
R919 B.n701 B.n700 10.6151
R920 B.n700 B.n699 10.6151
R921 B.n699 B.n44 10.6151
R922 B.n695 B.n44 10.6151
R923 B.n695 B.n694 10.6151
R924 B.n694 B.n693 10.6151
R925 B.n693 B.n46 10.6151
R926 B.n689 B.n46 10.6151
R927 B.n689 B.n688 10.6151
R928 B.n688 B.n687 10.6151
R929 B.n687 B.n48 10.6151
R930 B.n683 B.n48 10.6151
R931 B.n683 B.n682 10.6151
R932 B.n682 B.n681 10.6151
R933 B.n678 B.n677 10.6151
R934 B.n677 B.n676 10.6151
R935 B.n676 B.n54 10.6151
R936 B.n672 B.n54 10.6151
R937 B.n672 B.n671 10.6151
R938 B.n671 B.n670 10.6151
R939 B.n670 B.n56 10.6151
R940 B.n666 B.n56 10.6151
R941 B.n666 B.n665 10.6151
R942 B.n663 B.n60 10.6151
R943 B.n659 B.n60 10.6151
R944 B.n659 B.n658 10.6151
R945 B.n658 B.n657 10.6151
R946 B.n657 B.n62 10.6151
R947 B.n653 B.n62 10.6151
R948 B.n653 B.n652 10.6151
R949 B.n652 B.n651 10.6151
R950 B.n651 B.n64 10.6151
R951 B.n647 B.n64 10.6151
R952 B.n647 B.n646 10.6151
R953 B.n646 B.n645 10.6151
R954 B.n645 B.n66 10.6151
R955 B.n641 B.n66 10.6151
R956 B.n641 B.n640 10.6151
R957 B.n640 B.n639 10.6151
R958 B.n639 B.n68 10.6151
R959 B.n635 B.n68 10.6151
R960 B.n635 B.n634 10.6151
R961 B.n634 B.n633 10.6151
R962 B.n633 B.n70 10.6151
R963 B.n629 B.n70 10.6151
R964 B.n629 B.n628 10.6151
R965 B.n628 B.n627 10.6151
R966 B.n627 B.n72 10.6151
R967 B.n623 B.n72 10.6151
R968 B.n623 B.n622 10.6151
R969 B.n622 B.n621 10.6151
R970 B.n621 B.n74 10.6151
R971 B.n617 B.n74 10.6151
R972 B.n617 B.n616 10.6151
R973 B.n616 B.n615 10.6151
R974 B.n615 B.n76 10.6151
R975 B.n611 B.n76 10.6151
R976 B.n611 B.n610 10.6151
R977 B.n610 B.n609 10.6151
R978 B.n609 B.n78 10.6151
R979 B.n605 B.n78 10.6151
R980 B.n605 B.n604 10.6151
R981 B.n604 B.n603 10.6151
R982 B.n603 B.n80 10.6151
R983 B.n599 B.n598 10.6151
R984 B.n598 B.n597 10.6151
R985 B.n597 B.n82 10.6151
R986 B.n593 B.n82 10.6151
R987 B.n593 B.n592 10.6151
R988 B.n592 B.n591 10.6151
R989 B.n591 B.n84 10.6151
R990 B.n587 B.n84 10.6151
R991 B.n587 B.n586 10.6151
R992 B.n586 B.n585 10.6151
R993 B.n585 B.n86 10.6151
R994 B.n581 B.n86 10.6151
R995 B.n581 B.n580 10.6151
R996 B.n580 B.n579 10.6151
R997 B.n579 B.n88 10.6151
R998 B.n575 B.n88 10.6151
R999 B.n575 B.n574 10.6151
R1000 B.n574 B.n573 10.6151
R1001 B.n573 B.n90 10.6151
R1002 B.n569 B.n90 10.6151
R1003 B.n569 B.n568 10.6151
R1004 B.n568 B.n567 10.6151
R1005 B.n567 B.n92 10.6151
R1006 B.n563 B.n92 10.6151
R1007 B.n563 B.n562 10.6151
R1008 B.n562 B.n561 10.6151
R1009 B.n561 B.n94 10.6151
R1010 B.n557 B.n94 10.6151
R1011 B.n557 B.n556 10.6151
R1012 B.n556 B.n555 10.6151
R1013 B.n555 B.n96 10.6151
R1014 B.n551 B.n96 10.6151
R1015 B.n551 B.n550 10.6151
R1016 B.n550 B.n549 10.6151
R1017 B.n549 B.n98 10.6151
R1018 B.n545 B.n98 10.6151
R1019 B.n545 B.n544 10.6151
R1020 B.n544 B.n543 10.6151
R1021 B.n543 B.n100 10.6151
R1022 B.n539 B.n100 10.6151
R1023 B.n539 B.n538 10.6151
R1024 B.n538 B.n537 10.6151
R1025 B.n537 B.n102 10.6151
R1026 B.n533 B.n102 10.6151
R1027 B.n533 B.n532 10.6151
R1028 B.n532 B.n531 10.6151
R1029 B.n531 B.n104 10.6151
R1030 B.n527 B.n104 10.6151
R1031 B.n527 B.n526 10.6151
R1032 B.n526 B.n525 10.6151
R1033 B.n525 B.n106 10.6151
R1034 B.n521 B.n106 10.6151
R1035 B.n521 B.n520 10.6151
R1036 B.n520 B.n519 10.6151
R1037 B.n519 B.n108 10.6151
R1038 B.n515 B.n108 10.6151
R1039 B.n515 B.n514 10.6151
R1040 B.n514 B.n513 10.6151
R1041 B.n513 B.n110 10.6151
R1042 B.n509 B.n110 10.6151
R1043 B.n509 B.n508 10.6151
R1044 B.n508 B.n507 10.6151
R1045 B.n507 B.n112 10.6151
R1046 B.n503 B.n112 10.6151
R1047 B.n503 B.n502 10.6151
R1048 B.n502 B.n501 10.6151
R1049 B.n501 B.n114 10.6151
R1050 B.n497 B.n114 10.6151
R1051 B.n497 B.n496 10.6151
R1052 B.n496 B.n495 10.6151
R1053 B.n495 B.n116 10.6151
R1054 B.n491 B.n116 10.6151
R1055 B.n491 B.n490 10.6151
R1056 B.n490 B.n489 10.6151
R1057 B.n489 B.n118 10.6151
R1058 B.n485 B.n118 10.6151
R1059 B.n485 B.n484 10.6151
R1060 B.n484 B.n483 10.6151
R1061 B.n483 B.n120 10.6151
R1062 B.n479 B.n120 10.6151
R1063 B.n479 B.n478 10.6151
R1064 B.n478 B.n477 10.6151
R1065 B.n477 B.n122 10.6151
R1066 B.n473 B.n122 10.6151
R1067 B.n473 B.n472 10.6151
R1068 B.n472 B.n471 10.6151
R1069 B.n471 B.n124 10.6151
R1070 B.n467 B.n124 10.6151
R1071 B.n467 B.n466 10.6151
R1072 B.n466 B.n465 10.6151
R1073 B.n465 B.n126 10.6151
R1074 B.n461 B.n126 10.6151
R1075 B.n461 B.n460 10.6151
R1076 B.n460 B.n459 10.6151
R1077 B.n459 B.n128 10.6151
R1078 B.n455 B.n128 10.6151
R1079 B.n455 B.n454 10.6151
R1080 B.n454 B.n453 10.6151
R1081 B.n453 B.n130 10.6151
R1082 B.n449 B.n130 10.6151
R1083 B.n449 B.n448 10.6151
R1084 B.n448 B.n447 10.6151
R1085 B.n447 B.n132 10.6151
R1086 B.n443 B.n132 10.6151
R1087 B.n443 B.n442 10.6151
R1088 B.n442 B.n441 10.6151
R1089 B.n441 B.n134 10.6151
R1090 B.n437 B.n134 10.6151
R1091 B.n437 B.n436 10.6151
R1092 B.n211 B.n1 10.6151
R1093 B.n211 B.n210 10.6151
R1094 B.n215 B.n210 10.6151
R1095 B.n216 B.n215 10.6151
R1096 B.n217 B.n216 10.6151
R1097 B.n217 B.n208 10.6151
R1098 B.n221 B.n208 10.6151
R1099 B.n222 B.n221 10.6151
R1100 B.n223 B.n222 10.6151
R1101 B.n223 B.n206 10.6151
R1102 B.n227 B.n206 10.6151
R1103 B.n228 B.n227 10.6151
R1104 B.n229 B.n228 10.6151
R1105 B.n229 B.n204 10.6151
R1106 B.n233 B.n204 10.6151
R1107 B.n234 B.n233 10.6151
R1108 B.n235 B.n234 10.6151
R1109 B.n235 B.n202 10.6151
R1110 B.n239 B.n202 10.6151
R1111 B.n240 B.n239 10.6151
R1112 B.n241 B.n240 10.6151
R1113 B.n241 B.n200 10.6151
R1114 B.n245 B.n200 10.6151
R1115 B.n246 B.n245 10.6151
R1116 B.n247 B.n246 10.6151
R1117 B.n247 B.n198 10.6151
R1118 B.n251 B.n198 10.6151
R1119 B.n252 B.n251 10.6151
R1120 B.n253 B.n252 10.6151
R1121 B.n253 B.n196 10.6151
R1122 B.n257 B.n196 10.6151
R1123 B.n258 B.n257 10.6151
R1124 B.n259 B.n258 10.6151
R1125 B.n259 B.n194 10.6151
R1126 B.n263 B.n194 10.6151
R1127 B.n264 B.n263 10.6151
R1128 B.n265 B.n264 10.6151
R1129 B.n265 B.n192 10.6151
R1130 B.n269 B.n192 10.6151
R1131 B.n270 B.n269 10.6151
R1132 B.n271 B.n270 10.6151
R1133 B.n271 B.n190 10.6151
R1134 B.n275 B.n190 10.6151
R1135 B.n276 B.n275 10.6151
R1136 B.n277 B.n276 10.6151
R1137 B.n277 B.n188 10.6151
R1138 B.n281 B.n188 10.6151
R1139 B.n282 B.n281 10.6151
R1140 B.n283 B.n282 10.6151
R1141 B.n283 B.n186 10.6151
R1142 B.n287 B.n186 10.6151
R1143 B.n288 B.n287 10.6151
R1144 B.n289 B.n288 10.6151
R1145 B.n293 B.n184 10.6151
R1146 B.n294 B.n293 10.6151
R1147 B.n295 B.n294 10.6151
R1148 B.n295 B.n182 10.6151
R1149 B.n299 B.n182 10.6151
R1150 B.n300 B.n299 10.6151
R1151 B.n301 B.n300 10.6151
R1152 B.n301 B.n180 10.6151
R1153 B.n305 B.n180 10.6151
R1154 B.n306 B.n305 10.6151
R1155 B.n307 B.n306 10.6151
R1156 B.n307 B.n178 10.6151
R1157 B.n311 B.n178 10.6151
R1158 B.n312 B.n311 10.6151
R1159 B.n313 B.n312 10.6151
R1160 B.n313 B.n176 10.6151
R1161 B.n317 B.n176 10.6151
R1162 B.n318 B.n317 10.6151
R1163 B.n319 B.n318 10.6151
R1164 B.n319 B.n174 10.6151
R1165 B.n323 B.n174 10.6151
R1166 B.n324 B.n323 10.6151
R1167 B.n325 B.n324 10.6151
R1168 B.n325 B.n172 10.6151
R1169 B.n329 B.n172 10.6151
R1170 B.n330 B.n329 10.6151
R1171 B.n331 B.n330 10.6151
R1172 B.n331 B.n170 10.6151
R1173 B.n335 B.n170 10.6151
R1174 B.n336 B.n335 10.6151
R1175 B.n337 B.n336 10.6151
R1176 B.n337 B.n168 10.6151
R1177 B.n341 B.n168 10.6151
R1178 B.n342 B.n341 10.6151
R1179 B.n343 B.n342 10.6151
R1180 B.n343 B.n166 10.6151
R1181 B.n347 B.n166 10.6151
R1182 B.n348 B.n347 10.6151
R1183 B.n349 B.n348 10.6151
R1184 B.n349 B.n164 10.6151
R1185 B.n353 B.n164 10.6151
R1186 B.n356 B.n355 10.6151
R1187 B.n356 B.n160 10.6151
R1188 B.n360 B.n160 10.6151
R1189 B.n361 B.n360 10.6151
R1190 B.n362 B.n361 10.6151
R1191 B.n362 B.n158 10.6151
R1192 B.n366 B.n158 10.6151
R1193 B.n367 B.n366 10.6151
R1194 B.n371 B.n367 10.6151
R1195 B.n375 B.n156 10.6151
R1196 B.n376 B.n375 10.6151
R1197 B.n377 B.n376 10.6151
R1198 B.n377 B.n154 10.6151
R1199 B.n381 B.n154 10.6151
R1200 B.n382 B.n381 10.6151
R1201 B.n383 B.n382 10.6151
R1202 B.n383 B.n152 10.6151
R1203 B.n387 B.n152 10.6151
R1204 B.n388 B.n387 10.6151
R1205 B.n389 B.n388 10.6151
R1206 B.n389 B.n150 10.6151
R1207 B.n393 B.n150 10.6151
R1208 B.n394 B.n393 10.6151
R1209 B.n395 B.n394 10.6151
R1210 B.n395 B.n148 10.6151
R1211 B.n399 B.n148 10.6151
R1212 B.n400 B.n399 10.6151
R1213 B.n401 B.n400 10.6151
R1214 B.n401 B.n146 10.6151
R1215 B.n405 B.n146 10.6151
R1216 B.n406 B.n405 10.6151
R1217 B.n407 B.n406 10.6151
R1218 B.n407 B.n144 10.6151
R1219 B.n411 B.n144 10.6151
R1220 B.n412 B.n411 10.6151
R1221 B.n413 B.n412 10.6151
R1222 B.n413 B.n142 10.6151
R1223 B.n417 B.n142 10.6151
R1224 B.n418 B.n417 10.6151
R1225 B.n419 B.n418 10.6151
R1226 B.n419 B.n140 10.6151
R1227 B.n423 B.n140 10.6151
R1228 B.n424 B.n423 10.6151
R1229 B.n425 B.n424 10.6151
R1230 B.n425 B.n138 10.6151
R1231 B.n429 B.n138 10.6151
R1232 B.n430 B.n429 10.6151
R1233 B.n431 B.n430 10.6151
R1234 B.n431 B.n136 10.6151
R1235 B.n435 B.n136 10.6151
R1236 B.n681 B.n52 9.36635
R1237 B.n664 B.n663 9.36635
R1238 B.n354 B.n353 9.36635
R1239 B.n370 B.n156 9.36635
R1240 B.n825 B.n0 8.11757
R1241 B.n825 B.n1 8.11757
R1242 B.n678 B.n52 1.24928
R1243 B.n665 B.n664 1.24928
R1244 B.n355 B.n354 1.24928
R1245 B.n371 B.n370 1.24928
R1246 VP.n19 VP.n16 161.3
R1247 VP.n21 VP.n20 161.3
R1248 VP.n22 VP.n15 161.3
R1249 VP.n24 VP.n23 161.3
R1250 VP.n25 VP.n14 161.3
R1251 VP.n27 VP.n26 161.3
R1252 VP.n29 VP.n13 161.3
R1253 VP.n31 VP.n30 161.3
R1254 VP.n32 VP.n12 161.3
R1255 VP.n34 VP.n33 161.3
R1256 VP.n35 VP.n11 161.3
R1257 VP.n37 VP.n36 161.3
R1258 VP.n69 VP.n68 161.3
R1259 VP.n67 VP.n1 161.3
R1260 VP.n66 VP.n65 161.3
R1261 VP.n64 VP.n2 161.3
R1262 VP.n63 VP.n62 161.3
R1263 VP.n61 VP.n3 161.3
R1264 VP.n59 VP.n58 161.3
R1265 VP.n57 VP.n4 161.3
R1266 VP.n56 VP.n55 161.3
R1267 VP.n54 VP.n5 161.3
R1268 VP.n53 VP.n52 161.3
R1269 VP.n51 VP.n6 161.3
R1270 VP.n50 VP.n49 161.3
R1271 VP.n47 VP.n7 161.3
R1272 VP.n46 VP.n45 161.3
R1273 VP.n44 VP.n8 161.3
R1274 VP.n43 VP.n42 161.3
R1275 VP.n41 VP.n9 161.3
R1276 VP.n18 VP.t3 136.45
R1277 VP.n40 VP.t7 104.49
R1278 VP.n48 VP.t6 104.49
R1279 VP.n60 VP.t4 104.49
R1280 VP.n0 VP.t2 104.49
R1281 VP.n10 VP.t5 104.49
R1282 VP.n28 VP.t0 104.49
R1283 VP.n17 VP.t1 104.49
R1284 VP.n40 VP.n39 66.0897
R1285 VP.n70 VP.n0 66.0897
R1286 VP.n38 VP.n10 66.0897
R1287 VP.n18 VP.n17 57.5527
R1288 VP.n55 VP.n54 56.5193
R1289 VP.n23 VP.n22 56.5193
R1290 VP.n39 VP.n38 52.3175
R1291 VP.n46 VP.n8 49.2348
R1292 VP.n66 VP.n2 49.2348
R1293 VP.n34 VP.n12 49.2348
R1294 VP.n42 VP.n8 31.752
R1295 VP.n67 VP.n66 31.752
R1296 VP.n35 VP.n34 31.752
R1297 VP.n42 VP.n41 24.4675
R1298 VP.n47 VP.n46 24.4675
R1299 VP.n49 VP.n47 24.4675
R1300 VP.n53 VP.n6 24.4675
R1301 VP.n54 VP.n53 24.4675
R1302 VP.n55 VP.n4 24.4675
R1303 VP.n59 VP.n4 24.4675
R1304 VP.n62 VP.n61 24.4675
R1305 VP.n62 VP.n2 24.4675
R1306 VP.n68 VP.n67 24.4675
R1307 VP.n36 VP.n35 24.4675
R1308 VP.n23 VP.n14 24.4675
R1309 VP.n27 VP.n14 24.4675
R1310 VP.n30 VP.n29 24.4675
R1311 VP.n30 VP.n12 24.4675
R1312 VP.n21 VP.n16 24.4675
R1313 VP.n22 VP.n21 24.4675
R1314 VP.n41 VP.n40 23.9782
R1315 VP.n68 VP.n0 23.9782
R1316 VP.n36 VP.n10 23.9782
R1317 VP.n48 VP.n6 16.1487
R1318 VP.n60 VP.n59 16.1487
R1319 VP.n28 VP.n27 16.1487
R1320 VP.n17 VP.n16 16.1487
R1321 VP.n49 VP.n48 8.31928
R1322 VP.n61 VP.n60 8.31928
R1323 VP.n29 VP.n28 8.31928
R1324 VP.n19 VP.n18 5.24057
R1325 VP.n38 VP.n37 0.354971
R1326 VP.n39 VP.n9 0.354971
R1327 VP.n70 VP.n69 0.354971
R1328 VP VP.n70 0.26696
R1329 VP.n20 VP.n19 0.189894
R1330 VP.n20 VP.n15 0.189894
R1331 VP.n24 VP.n15 0.189894
R1332 VP.n25 VP.n24 0.189894
R1333 VP.n26 VP.n25 0.189894
R1334 VP.n26 VP.n13 0.189894
R1335 VP.n31 VP.n13 0.189894
R1336 VP.n32 VP.n31 0.189894
R1337 VP.n33 VP.n32 0.189894
R1338 VP.n33 VP.n11 0.189894
R1339 VP.n37 VP.n11 0.189894
R1340 VP.n43 VP.n9 0.189894
R1341 VP.n44 VP.n43 0.189894
R1342 VP.n45 VP.n44 0.189894
R1343 VP.n45 VP.n7 0.189894
R1344 VP.n50 VP.n7 0.189894
R1345 VP.n51 VP.n50 0.189894
R1346 VP.n52 VP.n51 0.189894
R1347 VP.n52 VP.n5 0.189894
R1348 VP.n56 VP.n5 0.189894
R1349 VP.n57 VP.n56 0.189894
R1350 VP.n58 VP.n57 0.189894
R1351 VP.n58 VP.n3 0.189894
R1352 VP.n63 VP.n3 0.189894
R1353 VP.n64 VP.n63 0.189894
R1354 VP.n65 VP.n64 0.189894
R1355 VP.n65 VP.n1 0.189894
R1356 VP.n69 VP.n1 0.189894
R1357 VDD1 VDD1.n0 77.3527
R1358 VDD1.n3 VDD1.n2 77.239
R1359 VDD1.n3 VDD1.n1 77.239
R1360 VDD1.n5 VDD1.n4 75.9313
R1361 VDD1.n5 VDD1.n3 47.1345
R1362 VDD1.n4 VDD1.t0 2.64964
R1363 VDD1.n4 VDD1.t5 2.64964
R1364 VDD1.n0 VDD1.t2 2.64964
R1365 VDD1.n0 VDD1.t4 2.64964
R1366 VDD1.n2 VDD1.t6 2.64964
R1367 VDD1.n2 VDD1.t1 2.64964
R1368 VDD1.n1 VDD1.t3 2.64964
R1369 VDD1.n1 VDD1.t7 2.64964
R1370 VDD1 VDD1.n5 1.30438
R1371 VTAIL.n11 VTAIL.t12 61.9028
R1372 VTAIL.n10 VTAIL.t1 61.9028
R1373 VTAIL.n7 VTAIL.t0 61.9028
R1374 VTAIL.n15 VTAIL.t2 61.9018
R1375 VTAIL.n2 VTAIL.t5 61.9018
R1376 VTAIL.n3 VTAIL.t13 61.9018
R1377 VTAIL.n6 VTAIL.t8 61.9018
R1378 VTAIL.n14 VTAIL.t10 61.9016
R1379 VTAIL.n13 VTAIL.n12 59.2537
R1380 VTAIL.n9 VTAIL.n8 59.2537
R1381 VTAIL.n1 VTAIL.n0 59.2535
R1382 VTAIL.n5 VTAIL.n4 59.2535
R1383 VTAIL.n15 VTAIL.n14 25.6686
R1384 VTAIL.n7 VTAIL.n6 25.6686
R1385 VTAIL.n9 VTAIL.n7 2.72464
R1386 VTAIL.n10 VTAIL.n9 2.72464
R1387 VTAIL.n13 VTAIL.n11 2.72464
R1388 VTAIL.n14 VTAIL.n13 2.72464
R1389 VTAIL.n6 VTAIL.n5 2.72464
R1390 VTAIL.n5 VTAIL.n3 2.72464
R1391 VTAIL.n2 VTAIL.n1 2.72464
R1392 VTAIL VTAIL.n15 2.66645
R1393 VTAIL.n0 VTAIL.t3 2.64964
R1394 VTAIL.n0 VTAIL.t6 2.64964
R1395 VTAIL.n4 VTAIL.t9 2.64964
R1396 VTAIL.n4 VTAIL.t11 2.64964
R1397 VTAIL.n12 VTAIL.t14 2.64964
R1398 VTAIL.n12 VTAIL.t15 2.64964
R1399 VTAIL.n8 VTAIL.t4 2.64964
R1400 VTAIL.n8 VTAIL.t7 2.64964
R1401 VTAIL.n11 VTAIL.n10 0.470328
R1402 VTAIL.n3 VTAIL.n2 0.470328
R1403 VTAIL VTAIL.n1 0.0586897
R1404 VN.n56 VN.n55 161.3
R1405 VN.n54 VN.n30 161.3
R1406 VN.n53 VN.n52 161.3
R1407 VN.n51 VN.n31 161.3
R1408 VN.n50 VN.n49 161.3
R1409 VN.n48 VN.n32 161.3
R1410 VN.n46 VN.n45 161.3
R1411 VN.n44 VN.n33 161.3
R1412 VN.n43 VN.n42 161.3
R1413 VN.n41 VN.n34 161.3
R1414 VN.n40 VN.n39 161.3
R1415 VN.n38 VN.n35 161.3
R1416 VN.n27 VN.n26 161.3
R1417 VN.n25 VN.n1 161.3
R1418 VN.n24 VN.n23 161.3
R1419 VN.n22 VN.n2 161.3
R1420 VN.n21 VN.n20 161.3
R1421 VN.n19 VN.n3 161.3
R1422 VN.n17 VN.n16 161.3
R1423 VN.n15 VN.n4 161.3
R1424 VN.n14 VN.n13 161.3
R1425 VN.n12 VN.n5 161.3
R1426 VN.n11 VN.n10 161.3
R1427 VN.n9 VN.n6 161.3
R1428 VN.n37 VN.t2 136.45
R1429 VN.n8 VN.t4 136.45
R1430 VN.n7 VN.t5 104.49
R1431 VN.n18 VN.t3 104.49
R1432 VN.n0 VN.t6 104.49
R1433 VN.n36 VN.t0 104.49
R1434 VN.n47 VN.t1 104.49
R1435 VN.n29 VN.t7 104.49
R1436 VN.n28 VN.n0 66.0897
R1437 VN.n57 VN.n29 66.0897
R1438 VN.n8 VN.n7 57.5527
R1439 VN.n37 VN.n36 57.5527
R1440 VN.n13 VN.n12 56.5193
R1441 VN.n42 VN.n41 56.5193
R1442 VN VN.n57 52.4829
R1443 VN.n24 VN.n2 49.2348
R1444 VN.n53 VN.n31 49.2348
R1445 VN.n25 VN.n24 31.752
R1446 VN.n54 VN.n53 31.752
R1447 VN.n11 VN.n6 24.4675
R1448 VN.n12 VN.n11 24.4675
R1449 VN.n13 VN.n4 24.4675
R1450 VN.n17 VN.n4 24.4675
R1451 VN.n20 VN.n19 24.4675
R1452 VN.n20 VN.n2 24.4675
R1453 VN.n26 VN.n25 24.4675
R1454 VN.n41 VN.n40 24.4675
R1455 VN.n40 VN.n35 24.4675
R1456 VN.n49 VN.n31 24.4675
R1457 VN.n49 VN.n48 24.4675
R1458 VN.n46 VN.n33 24.4675
R1459 VN.n42 VN.n33 24.4675
R1460 VN.n55 VN.n54 24.4675
R1461 VN.n26 VN.n0 23.9782
R1462 VN.n55 VN.n29 23.9782
R1463 VN.n7 VN.n6 16.1487
R1464 VN.n18 VN.n17 16.1487
R1465 VN.n36 VN.n35 16.1487
R1466 VN.n47 VN.n46 16.1487
R1467 VN.n19 VN.n18 8.31928
R1468 VN.n48 VN.n47 8.31928
R1469 VN.n38 VN.n37 5.2406
R1470 VN.n9 VN.n8 5.2406
R1471 VN.n57 VN.n56 0.354971
R1472 VN.n28 VN.n27 0.354971
R1473 VN VN.n28 0.26696
R1474 VN.n56 VN.n30 0.189894
R1475 VN.n52 VN.n30 0.189894
R1476 VN.n52 VN.n51 0.189894
R1477 VN.n51 VN.n50 0.189894
R1478 VN.n50 VN.n32 0.189894
R1479 VN.n45 VN.n32 0.189894
R1480 VN.n45 VN.n44 0.189894
R1481 VN.n44 VN.n43 0.189894
R1482 VN.n43 VN.n34 0.189894
R1483 VN.n39 VN.n34 0.189894
R1484 VN.n39 VN.n38 0.189894
R1485 VN.n10 VN.n9 0.189894
R1486 VN.n10 VN.n5 0.189894
R1487 VN.n14 VN.n5 0.189894
R1488 VN.n15 VN.n14 0.189894
R1489 VN.n16 VN.n15 0.189894
R1490 VN.n16 VN.n3 0.189894
R1491 VN.n21 VN.n3 0.189894
R1492 VN.n22 VN.n21 0.189894
R1493 VN.n23 VN.n22 0.189894
R1494 VN.n23 VN.n1 0.189894
R1495 VN.n27 VN.n1 0.189894
R1496 VDD2.n2 VDD2.n1 77.239
R1497 VDD2.n2 VDD2.n0 77.239
R1498 VDD2 VDD2.n5 77.2352
R1499 VDD2.n4 VDD2.n3 75.9325
R1500 VDD2.n4 VDD2.n2 46.5515
R1501 VDD2.n5 VDD2.t7 2.64964
R1502 VDD2.n5 VDD2.t5 2.64964
R1503 VDD2.n3 VDD2.t0 2.64964
R1504 VDD2.n3 VDD2.t6 2.64964
R1505 VDD2.n1 VDD2.t4 2.64964
R1506 VDD2.n1 VDD2.t1 2.64964
R1507 VDD2.n0 VDD2.t3 2.64964
R1508 VDD2.n0 VDD2.t2 2.64964
R1509 VDD2 VDD2.n4 1.42076
C0 VDD2 B 1.82926f
C1 w_n4130_n3422# B 10.543599f
C2 VP VTAIL 9.49461f
C3 VDD1 VP 9.414889f
C4 VDD1 VTAIL 8.22136f
C5 VDD2 VN 9.0244f
C6 w_n4130_n3422# VN 8.478629f
C7 B VP 2.18306f
C8 B VTAIL 5.17576f
C9 B VDD1 1.726f
C10 VDD2 w_n4130_n3422# 2.15862f
C11 VN VP 7.99614f
C12 VN VTAIL 9.4805f
C13 VN VDD1 0.151975f
C14 VDD2 VP 0.543976f
C15 w_n4130_n3422# VP 9.01547f
C16 VDD2 VTAIL 8.27732f
C17 B VN 1.28191f
C18 w_n4130_n3422# VTAIL 4.29277f
C19 VDD2 VDD1 1.89599f
C20 w_n4130_n3422# VDD1 2.03427f
C21 VDD2 VSUBS 1.952843f
C22 VDD1 VSUBS 2.63302f
C23 VTAIL VSUBS 1.389408f
C24 VN VSUBS 7.06508f
C25 VP VSUBS 3.846992f
C26 B VSUBS 5.284576f
C27 w_n4130_n3422# VSUBS 0.173906p
C28 VDD2.t3 VSUBS 0.264707f
C29 VDD2.t2 VSUBS 0.264707f
C30 VDD2.n0 VSUBS 2.10978f
C31 VDD2.t4 VSUBS 0.264707f
C32 VDD2.t1 VSUBS 0.264707f
C33 VDD2.n1 VSUBS 2.10978f
C34 VDD2.n2 VSUBS 4.27501f
C35 VDD2.t0 VSUBS 0.264707f
C36 VDD2.t6 VSUBS 0.264707f
C37 VDD2.n3 VSUBS 2.09525f
C38 VDD2.n4 VSUBS 3.59938f
C39 VDD2.t7 VSUBS 0.264707f
C40 VDD2.t5 VSUBS 0.264707f
C41 VDD2.n5 VSUBS 2.10973f
C42 VN.t6 VSUBS 2.6149f
C43 VN.n0 VSUBS 1.03272f
C44 VN.n1 VSUBS 0.027621f
C45 VN.n2 VSUBS 0.051221f
C46 VN.n3 VSUBS 0.027621f
C47 VN.t3 VSUBS 2.6149f
C48 VN.n4 VSUBS 0.051479f
C49 VN.n5 VSUBS 0.027621f
C50 VN.n6 VSUBS 0.042838f
C51 VN.t5 VSUBS 2.6149f
C52 VN.n7 VSUBS 1.01074f
C53 VN.t4 VSUBS 2.87373f
C54 VN.n8 VSUBS 0.978168f
C55 VN.n9 VSUBS 0.291097f
C56 VN.n10 VSUBS 0.027621f
C57 VN.n11 VSUBS 0.051479f
C58 VN.n12 VSUBS 0.040322f
C59 VN.n13 VSUBS 0.040322f
C60 VN.n14 VSUBS 0.027621f
C61 VN.n15 VSUBS 0.027621f
C62 VN.n16 VSUBS 0.027621f
C63 VN.n17 VSUBS 0.042838f
C64 VN.n18 VSUBS 0.92139f
C65 VN.n19 VSUBS 0.034705f
C66 VN.n20 VSUBS 0.051479f
C67 VN.n21 VSUBS 0.027621f
C68 VN.n22 VSUBS 0.027621f
C69 VN.n23 VSUBS 0.027621f
C70 VN.n24 VSUBS 0.025343f
C71 VN.n25 VSUBS 0.055559f
C72 VN.n26 VSUBS 0.050971f
C73 VN.n27 VSUBS 0.04458f
C74 VN.n28 VSUBS 0.050833f
C75 VN.t7 VSUBS 2.6149f
C76 VN.n29 VSUBS 1.03272f
C77 VN.n30 VSUBS 0.027621f
C78 VN.n31 VSUBS 0.051221f
C79 VN.n32 VSUBS 0.027621f
C80 VN.t1 VSUBS 2.6149f
C81 VN.n33 VSUBS 0.051479f
C82 VN.n34 VSUBS 0.027621f
C83 VN.n35 VSUBS 0.042838f
C84 VN.t2 VSUBS 2.87373f
C85 VN.t0 VSUBS 2.6149f
C86 VN.n36 VSUBS 1.01074f
C87 VN.n37 VSUBS 0.978168f
C88 VN.n38 VSUBS 0.291097f
C89 VN.n39 VSUBS 0.027621f
C90 VN.n40 VSUBS 0.051479f
C91 VN.n41 VSUBS 0.040322f
C92 VN.n42 VSUBS 0.040322f
C93 VN.n43 VSUBS 0.027621f
C94 VN.n44 VSUBS 0.027621f
C95 VN.n45 VSUBS 0.027621f
C96 VN.n46 VSUBS 0.042838f
C97 VN.n47 VSUBS 0.92139f
C98 VN.n48 VSUBS 0.034705f
C99 VN.n49 VSUBS 0.051479f
C100 VN.n50 VSUBS 0.027621f
C101 VN.n51 VSUBS 0.027621f
C102 VN.n52 VSUBS 0.027621f
C103 VN.n53 VSUBS 0.025343f
C104 VN.n54 VSUBS 0.055559f
C105 VN.n55 VSUBS 0.050971f
C106 VN.n56 VSUBS 0.04458f
C107 VN.n57 VSUBS 1.67032f
C108 VTAIL.t3 VSUBS 0.244749f
C109 VTAIL.t6 VSUBS 0.244749f
C110 VTAIL.n0 VSUBS 1.81033f
C111 VTAIL.n1 VSUBS 0.774721f
C112 VTAIL.t5 VSUBS 2.38226f
C113 VTAIL.n2 VSUBS 0.903764f
C114 VTAIL.t13 VSUBS 2.38226f
C115 VTAIL.n3 VSUBS 0.903764f
C116 VTAIL.t9 VSUBS 0.244749f
C117 VTAIL.t11 VSUBS 0.244749f
C118 VTAIL.n4 VSUBS 1.81033f
C119 VTAIL.n5 VSUBS 0.991557f
C120 VTAIL.t8 VSUBS 2.38226f
C121 VTAIL.n6 VSUBS 2.29033f
C122 VTAIL.t0 VSUBS 2.38226f
C123 VTAIL.n7 VSUBS 2.29033f
C124 VTAIL.t4 VSUBS 0.244749f
C125 VTAIL.t7 VSUBS 0.244749f
C126 VTAIL.n8 VSUBS 1.81033f
C127 VTAIL.n9 VSUBS 0.991549f
C128 VTAIL.t1 VSUBS 2.38226f
C129 VTAIL.n10 VSUBS 0.90376f
C130 VTAIL.t12 VSUBS 2.38226f
C131 VTAIL.n11 VSUBS 0.90376f
C132 VTAIL.t14 VSUBS 0.244749f
C133 VTAIL.t15 VSUBS 0.244749f
C134 VTAIL.n12 VSUBS 1.81033f
C135 VTAIL.n13 VSUBS 0.991549f
C136 VTAIL.t10 VSUBS 2.38225f
C137 VTAIL.n14 VSUBS 2.29034f
C138 VTAIL.t2 VSUBS 2.38226f
C139 VTAIL.n15 VSUBS 2.2856f
C140 VDD1.t2 VSUBS 0.264696f
C141 VDD1.t4 VSUBS 0.264696f
C142 VDD1.n0 VSUBS 2.1111f
C143 VDD1.t3 VSUBS 0.264696f
C144 VDD1.t7 VSUBS 0.264696f
C145 VDD1.n1 VSUBS 2.10969f
C146 VDD1.t6 VSUBS 0.264696f
C147 VDD1.t1 VSUBS 0.264696f
C148 VDD1.n2 VSUBS 2.10969f
C149 VDD1.n3 VSUBS 4.33154f
C150 VDD1.t0 VSUBS 0.264696f
C151 VDD1.t5 VSUBS 0.264696f
C152 VDD1.n4 VSUBS 2.09515f
C153 VDD1.n5 VSUBS 3.63311f
C154 VP.t2 VSUBS 2.84967f
C155 VP.n0 VSUBS 1.12544f
C156 VP.n1 VSUBS 0.030101f
C157 VP.n2 VSUBS 0.05582f
C158 VP.n3 VSUBS 0.030101f
C159 VP.t4 VSUBS 2.84967f
C160 VP.n4 VSUBS 0.056101f
C161 VP.n5 VSUBS 0.030101f
C162 VP.n6 VSUBS 0.046684f
C163 VP.n7 VSUBS 0.030101f
C164 VP.n8 VSUBS 0.027618f
C165 VP.n9 VSUBS 0.048583f
C166 VP.t7 VSUBS 2.84967f
C167 VP.t5 VSUBS 2.84967f
C168 VP.n10 VSUBS 1.12544f
C169 VP.n11 VSUBS 0.030101f
C170 VP.n12 VSUBS 0.05582f
C171 VP.n13 VSUBS 0.030101f
C172 VP.t0 VSUBS 2.84967f
C173 VP.n14 VSUBS 0.056101f
C174 VP.n15 VSUBS 0.030101f
C175 VP.n16 VSUBS 0.046684f
C176 VP.t3 VSUBS 3.13173f
C177 VP.t1 VSUBS 2.84967f
C178 VP.n17 VSUBS 1.10149f
C179 VP.n18 VSUBS 1.06599f
C180 VP.n19 VSUBS 0.317232f
C181 VP.n20 VSUBS 0.030101f
C182 VP.n21 VSUBS 0.056101f
C183 VP.n22 VSUBS 0.043942f
C184 VP.n23 VSUBS 0.043942f
C185 VP.n24 VSUBS 0.030101f
C186 VP.n25 VSUBS 0.030101f
C187 VP.n26 VSUBS 0.030101f
C188 VP.n27 VSUBS 0.046684f
C189 VP.n28 VSUBS 1.00411f
C190 VP.n29 VSUBS 0.037821f
C191 VP.n30 VSUBS 0.056101f
C192 VP.n31 VSUBS 0.030101f
C193 VP.n32 VSUBS 0.030101f
C194 VP.n33 VSUBS 0.030101f
C195 VP.n34 VSUBS 0.027618f
C196 VP.n35 VSUBS 0.060547f
C197 VP.n36 VSUBS 0.055547f
C198 VP.n37 VSUBS 0.048583f
C199 VP.n38 VSUBS 1.80816f
C200 VP.n39 VSUBS 1.82884f
C201 VP.n40 VSUBS 1.12544f
C202 VP.n41 VSUBS 0.055547f
C203 VP.n42 VSUBS 0.060547f
C204 VP.n43 VSUBS 0.030101f
C205 VP.n44 VSUBS 0.030101f
C206 VP.n45 VSUBS 0.030101f
C207 VP.n46 VSUBS 0.05582f
C208 VP.n47 VSUBS 0.056101f
C209 VP.t6 VSUBS 2.84967f
C210 VP.n48 VSUBS 1.00411f
C211 VP.n49 VSUBS 0.037821f
C212 VP.n50 VSUBS 0.030101f
C213 VP.n51 VSUBS 0.030101f
C214 VP.n52 VSUBS 0.030101f
C215 VP.n53 VSUBS 0.056101f
C216 VP.n54 VSUBS 0.043942f
C217 VP.n55 VSUBS 0.043942f
C218 VP.n56 VSUBS 0.030101f
C219 VP.n57 VSUBS 0.030101f
C220 VP.n58 VSUBS 0.030101f
C221 VP.n59 VSUBS 0.046684f
C222 VP.n60 VSUBS 1.00411f
C223 VP.n61 VSUBS 0.037821f
C224 VP.n62 VSUBS 0.056101f
C225 VP.n63 VSUBS 0.030101f
C226 VP.n64 VSUBS 0.030101f
C227 VP.n65 VSUBS 0.030101f
C228 VP.n66 VSUBS 0.027618f
C229 VP.n67 VSUBS 0.060547f
C230 VP.n68 VSUBS 0.055547f
C231 VP.n69 VSUBS 0.048583f
C232 VP.n70 VSUBS 0.055397f
C233 B.n0 VSUBS 0.006585f
C234 B.n1 VSUBS 0.006585f
C235 B.n2 VSUBS 0.009738f
C236 B.n3 VSUBS 0.007463f
C237 B.n4 VSUBS 0.007463f
C238 B.n5 VSUBS 0.007463f
C239 B.n6 VSUBS 0.007463f
C240 B.n7 VSUBS 0.007463f
C241 B.n8 VSUBS 0.007463f
C242 B.n9 VSUBS 0.007463f
C243 B.n10 VSUBS 0.007463f
C244 B.n11 VSUBS 0.007463f
C245 B.n12 VSUBS 0.007463f
C246 B.n13 VSUBS 0.007463f
C247 B.n14 VSUBS 0.007463f
C248 B.n15 VSUBS 0.007463f
C249 B.n16 VSUBS 0.007463f
C250 B.n17 VSUBS 0.007463f
C251 B.n18 VSUBS 0.007463f
C252 B.n19 VSUBS 0.007463f
C253 B.n20 VSUBS 0.007463f
C254 B.n21 VSUBS 0.007463f
C255 B.n22 VSUBS 0.007463f
C256 B.n23 VSUBS 0.007463f
C257 B.n24 VSUBS 0.007463f
C258 B.n25 VSUBS 0.007463f
C259 B.n26 VSUBS 0.007463f
C260 B.n27 VSUBS 0.007463f
C261 B.n28 VSUBS 0.007463f
C262 B.n29 VSUBS 0.018745f
C263 B.n30 VSUBS 0.007463f
C264 B.n31 VSUBS 0.007463f
C265 B.n32 VSUBS 0.007463f
C266 B.n33 VSUBS 0.007463f
C267 B.n34 VSUBS 0.007463f
C268 B.n35 VSUBS 0.007463f
C269 B.n36 VSUBS 0.007463f
C270 B.n37 VSUBS 0.007463f
C271 B.n38 VSUBS 0.007463f
C272 B.n39 VSUBS 0.007463f
C273 B.n40 VSUBS 0.007463f
C274 B.n41 VSUBS 0.007463f
C275 B.n42 VSUBS 0.007463f
C276 B.n43 VSUBS 0.007463f
C277 B.n44 VSUBS 0.007463f
C278 B.n45 VSUBS 0.007463f
C279 B.n46 VSUBS 0.007463f
C280 B.n47 VSUBS 0.007463f
C281 B.n48 VSUBS 0.007463f
C282 B.n49 VSUBS 0.007463f
C283 B.t7 VSUBS 0.427279f
C284 B.t8 VSUBS 0.451574f
C285 B.t6 VSUBS 1.69344f
C286 B.n50 VSUBS 0.241911f
C287 B.n51 VSUBS 0.0776f
C288 B.n52 VSUBS 0.01729f
C289 B.n53 VSUBS 0.007463f
C290 B.n54 VSUBS 0.007463f
C291 B.n55 VSUBS 0.007463f
C292 B.n56 VSUBS 0.007463f
C293 B.n57 VSUBS 0.007463f
C294 B.t10 VSUBS 0.42727f
C295 B.t11 VSUBS 0.451566f
C296 B.t9 VSUBS 1.69344f
C297 B.n58 VSUBS 0.241918f
C298 B.n59 VSUBS 0.077609f
C299 B.n60 VSUBS 0.007463f
C300 B.n61 VSUBS 0.007463f
C301 B.n62 VSUBS 0.007463f
C302 B.n63 VSUBS 0.007463f
C303 B.n64 VSUBS 0.007463f
C304 B.n65 VSUBS 0.007463f
C305 B.n66 VSUBS 0.007463f
C306 B.n67 VSUBS 0.007463f
C307 B.n68 VSUBS 0.007463f
C308 B.n69 VSUBS 0.007463f
C309 B.n70 VSUBS 0.007463f
C310 B.n71 VSUBS 0.007463f
C311 B.n72 VSUBS 0.007463f
C312 B.n73 VSUBS 0.007463f
C313 B.n74 VSUBS 0.007463f
C314 B.n75 VSUBS 0.007463f
C315 B.n76 VSUBS 0.007463f
C316 B.n77 VSUBS 0.007463f
C317 B.n78 VSUBS 0.007463f
C318 B.n79 VSUBS 0.007463f
C319 B.n80 VSUBS 0.018745f
C320 B.n81 VSUBS 0.007463f
C321 B.n82 VSUBS 0.007463f
C322 B.n83 VSUBS 0.007463f
C323 B.n84 VSUBS 0.007463f
C324 B.n85 VSUBS 0.007463f
C325 B.n86 VSUBS 0.007463f
C326 B.n87 VSUBS 0.007463f
C327 B.n88 VSUBS 0.007463f
C328 B.n89 VSUBS 0.007463f
C329 B.n90 VSUBS 0.007463f
C330 B.n91 VSUBS 0.007463f
C331 B.n92 VSUBS 0.007463f
C332 B.n93 VSUBS 0.007463f
C333 B.n94 VSUBS 0.007463f
C334 B.n95 VSUBS 0.007463f
C335 B.n96 VSUBS 0.007463f
C336 B.n97 VSUBS 0.007463f
C337 B.n98 VSUBS 0.007463f
C338 B.n99 VSUBS 0.007463f
C339 B.n100 VSUBS 0.007463f
C340 B.n101 VSUBS 0.007463f
C341 B.n102 VSUBS 0.007463f
C342 B.n103 VSUBS 0.007463f
C343 B.n104 VSUBS 0.007463f
C344 B.n105 VSUBS 0.007463f
C345 B.n106 VSUBS 0.007463f
C346 B.n107 VSUBS 0.007463f
C347 B.n108 VSUBS 0.007463f
C348 B.n109 VSUBS 0.007463f
C349 B.n110 VSUBS 0.007463f
C350 B.n111 VSUBS 0.007463f
C351 B.n112 VSUBS 0.007463f
C352 B.n113 VSUBS 0.007463f
C353 B.n114 VSUBS 0.007463f
C354 B.n115 VSUBS 0.007463f
C355 B.n116 VSUBS 0.007463f
C356 B.n117 VSUBS 0.007463f
C357 B.n118 VSUBS 0.007463f
C358 B.n119 VSUBS 0.007463f
C359 B.n120 VSUBS 0.007463f
C360 B.n121 VSUBS 0.007463f
C361 B.n122 VSUBS 0.007463f
C362 B.n123 VSUBS 0.007463f
C363 B.n124 VSUBS 0.007463f
C364 B.n125 VSUBS 0.007463f
C365 B.n126 VSUBS 0.007463f
C366 B.n127 VSUBS 0.007463f
C367 B.n128 VSUBS 0.007463f
C368 B.n129 VSUBS 0.007463f
C369 B.n130 VSUBS 0.007463f
C370 B.n131 VSUBS 0.007463f
C371 B.n132 VSUBS 0.007463f
C372 B.n133 VSUBS 0.007463f
C373 B.n134 VSUBS 0.007463f
C374 B.n135 VSUBS 0.01813f
C375 B.n136 VSUBS 0.007463f
C376 B.n137 VSUBS 0.007463f
C377 B.n138 VSUBS 0.007463f
C378 B.n139 VSUBS 0.007463f
C379 B.n140 VSUBS 0.007463f
C380 B.n141 VSUBS 0.007463f
C381 B.n142 VSUBS 0.007463f
C382 B.n143 VSUBS 0.007463f
C383 B.n144 VSUBS 0.007463f
C384 B.n145 VSUBS 0.007463f
C385 B.n146 VSUBS 0.007463f
C386 B.n147 VSUBS 0.007463f
C387 B.n148 VSUBS 0.007463f
C388 B.n149 VSUBS 0.007463f
C389 B.n150 VSUBS 0.007463f
C390 B.n151 VSUBS 0.007463f
C391 B.n152 VSUBS 0.007463f
C392 B.n153 VSUBS 0.007463f
C393 B.n154 VSUBS 0.007463f
C394 B.n155 VSUBS 0.007463f
C395 B.n156 VSUBS 0.007024f
C396 B.n157 VSUBS 0.007463f
C397 B.n158 VSUBS 0.007463f
C398 B.n159 VSUBS 0.007463f
C399 B.n160 VSUBS 0.007463f
C400 B.n161 VSUBS 0.007463f
C401 B.t2 VSUBS 0.427279f
C402 B.t1 VSUBS 0.451574f
C403 B.t0 VSUBS 1.69344f
C404 B.n162 VSUBS 0.241911f
C405 B.n163 VSUBS 0.0776f
C406 B.n164 VSUBS 0.007463f
C407 B.n165 VSUBS 0.007463f
C408 B.n166 VSUBS 0.007463f
C409 B.n167 VSUBS 0.007463f
C410 B.n168 VSUBS 0.007463f
C411 B.n169 VSUBS 0.007463f
C412 B.n170 VSUBS 0.007463f
C413 B.n171 VSUBS 0.007463f
C414 B.n172 VSUBS 0.007463f
C415 B.n173 VSUBS 0.007463f
C416 B.n174 VSUBS 0.007463f
C417 B.n175 VSUBS 0.007463f
C418 B.n176 VSUBS 0.007463f
C419 B.n177 VSUBS 0.007463f
C420 B.n178 VSUBS 0.007463f
C421 B.n179 VSUBS 0.007463f
C422 B.n180 VSUBS 0.007463f
C423 B.n181 VSUBS 0.007463f
C424 B.n182 VSUBS 0.007463f
C425 B.n183 VSUBS 0.007463f
C426 B.n184 VSUBS 0.018745f
C427 B.n185 VSUBS 0.007463f
C428 B.n186 VSUBS 0.007463f
C429 B.n187 VSUBS 0.007463f
C430 B.n188 VSUBS 0.007463f
C431 B.n189 VSUBS 0.007463f
C432 B.n190 VSUBS 0.007463f
C433 B.n191 VSUBS 0.007463f
C434 B.n192 VSUBS 0.007463f
C435 B.n193 VSUBS 0.007463f
C436 B.n194 VSUBS 0.007463f
C437 B.n195 VSUBS 0.007463f
C438 B.n196 VSUBS 0.007463f
C439 B.n197 VSUBS 0.007463f
C440 B.n198 VSUBS 0.007463f
C441 B.n199 VSUBS 0.007463f
C442 B.n200 VSUBS 0.007463f
C443 B.n201 VSUBS 0.007463f
C444 B.n202 VSUBS 0.007463f
C445 B.n203 VSUBS 0.007463f
C446 B.n204 VSUBS 0.007463f
C447 B.n205 VSUBS 0.007463f
C448 B.n206 VSUBS 0.007463f
C449 B.n207 VSUBS 0.007463f
C450 B.n208 VSUBS 0.007463f
C451 B.n209 VSUBS 0.007463f
C452 B.n210 VSUBS 0.007463f
C453 B.n211 VSUBS 0.007463f
C454 B.n212 VSUBS 0.007463f
C455 B.n213 VSUBS 0.007463f
C456 B.n214 VSUBS 0.007463f
C457 B.n215 VSUBS 0.007463f
C458 B.n216 VSUBS 0.007463f
C459 B.n217 VSUBS 0.007463f
C460 B.n218 VSUBS 0.007463f
C461 B.n219 VSUBS 0.007463f
C462 B.n220 VSUBS 0.007463f
C463 B.n221 VSUBS 0.007463f
C464 B.n222 VSUBS 0.007463f
C465 B.n223 VSUBS 0.007463f
C466 B.n224 VSUBS 0.007463f
C467 B.n225 VSUBS 0.007463f
C468 B.n226 VSUBS 0.007463f
C469 B.n227 VSUBS 0.007463f
C470 B.n228 VSUBS 0.007463f
C471 B.n229 VSUBS 0.007463f
C472 B.n230 VSUBS 0.007463f
C473 B.n231 VSUBS 0.007463f
C474 B.n232 VSUBS 0.007463f
C475 B.n233 VSUBS 0.007463f
C476 B.n234 VSUBS 0.007463f
C477 B.n235 VSUBS 0.007463f
C478 B.n236 VSUBS 0.007463f
C479 B.n237 VSUBS 0.007463f
C480 B.n238 VSUBS 0.007463f
C481 B.n239 VSUBS 0.007463f
C482 B.n240 VSUBS 0.007463f
C483 B.n241 VSUBS 0.007463f
C484 B.n242 VSUBS 0.007463f
C485 B.n243 VSUBS 0.007463f
C486 B.n244 VSUBS 0.007463f
C487 B.n245 VSUBS 0.007463f
C488 B.n246 VSUBS 0.007463f
C489 B.n247 VSUBS 0.007463f
C490 B.n248 VSUBS 0.007463f
C491 B.n249 VSUBS 0.007463f
C492 B.n250 VSUBS 0.007463f
C493 B.n251 VSUBS 0.007463f
C494 B.n252 VSUBS 0.007463f
C495 B.n253 VSUBS 0.007463f
C496 B.n254 VSUBS 0.007463f
C497 B.n255 VSUBS 0.007463f
C498 B.n256 VSUBS 0.007463f
C499 B.n257 VSUBS 0.007463f
C500 B.n258 VSUBS 0.007463f
C501 B.n259 VSUBS 0.007463f
C502 B.n260 VSUBS 0.007463f
C503 B.n261 VSUBS 0.007463f
C504 B.n262 VSUBS 0.007463f
C505 B.n263 VSUBS 0.007463f
C506 B.n264 VSUBS 0.007463f
C507 B.n265 VSUBS 0.007463f
C508 B.n266 VSUBS 0.007463f
C509 B.n267 VSUBS 0.007463f
C510 B.n268 VSUBS 0.007463f
C511 B.n269 VSUBS 0.007463f
C512 B.n270 VSUBS 0.007463f
C513 B.n271 VSUBS 0.007463f
C514 B.n272 VSUBS 0.007463f
C515 B.n273 VSUBS 0.007463f
C516 B.n274 VSUBS 0.007463f
C517 B.n275 VSUBS 0.007463f
C518 B.n276 VSUBS 0.007463f
C519 B.n277 VSUBS 0.007463f
C520 B.n278 VSUBS 0.007463f
C521 B.n279 VSUBS 0.007463f
C522 B.n280 VSUBS 0.007463f
C523 B.n281 VSUBS 0.007463f
C524 B.n282 VSUBS 0.007463f
C525 B.n283 VSUBS 0.007463f
C526 B.n284 VSUBS 0.007463f
C527 B.n285 VSUBS 0.007463f
C528 B.n286 VSUBS 0.007463f
C529 B.n287 VSUBS 0.007463f
C530 B.n288 VSUBS 0.007463f
C531 B.n289 VSUBS 0.01813f
C532 B.n290 VSUBS 0.01813f
C533 B.n291 VSUBS 0.018745f
C534 B.n292 VSUBS 0.007463f
C535 B.n293 VSUBS 0.007463f
C536 B.n294 VSUBS 0.007463f
C537 B.n295 VSUBS 0.007463f
C538 B.n296 VSUBS 0.007463f
C539 B.n297 VSUBS 0.007463f
C540 B.n298 VSUBS 0.007463f
C541 B.n299 VSUBS 0.007463f
C542 B.n300 VSUBS 0.007463f
C543 B.n301 VSUBS 0.007463f
C544 B.n302 VSUBS 0.007463f
C545 B.n303 VSUBS 0.007463f
C546 B.n304 VSUBS 0.007463f
C547 B.n305 VSUBS 0.007463f
C548 B.n306 VSUBS 0.007463f
C549 B.n307 VSUBS 0.007463f
C550 B.n308 VSUBS 0.007463f
C551 B.n309 VSUBS 0.007463f
C552 B.n310 VSUBS 0.007463f
C553 B.n311 VSUBS 0.007463f
C554 B.n312 VSUBS 0.007463f
C555 B.n313 VSUBS 0.007463f
C556 B.n314 VSUBS 0.007463f
C557 B.n315 VSUBS 0.007463f
C558 B.n316 VSUBS 0.007463f
C559 B.n317 VSUBS 0.007463f
C560 B.n318 VSUBS 0.007463f
C561 B.n319 VSUBS 0.007463f
C562 B.n320 VSUBS 0.007463f
C563 B.n321 VSUBS 0.007463f
C564 B.n322 VSUBS 0.007463f
C565 B.n323 VSUBS 0.007463f
C566 B.n324 VSUBS 0.007463f
C567 B.n325 VSUBS 0.007463f
C568 B.n326 VSUBS 0.007463f
C569 B.n327 VSUBS 0.007463f
C570 B.n328 VSUBS 0.007463f
C571 B.n329 VSUBS 0.007463f
C572 B.n330 VSUBS 0.007463f
C573 B.n331 VSUBS 0.007463f
C574 B.n332 VSUBS 0.007463f
C575 B.n333 VSUBS 0.007463f
C576 B.n334 VSUBS 0.007463f
C577 B.n335 VSUBS 0.007463f
C578 B.n336 VSUBS 0.007463f
C579 B.n337 VSUBS 0.007463f
C580 B.n338 VSUBS 0.007463f
C581 B.n339 VSUBS 0.007463f
C582 B.n340 VSUBS 0.007463f
C583 B.n341 VSUBS 0.007463f
C584 B.n342 VSUBS 0.007463f
C585 B.n343 VSUBS 0.007463f
C586 B.n344 VSUBS 0.007463f
C587 B.n345 VSUBS 0.007463f
C588 B.n346 VSUBS 0.007463f
C589 B.n347 VSUBS 0.007463f
C590 B.n348 VSUBS 0.007463f
C591 B.n349 VSUBS 0.007463f
C592 B.n350 VSUBS 0.007463f
C593 B.n351 VSUBS 0.007463f
C594 B.n352 VSUBS 0.007463f
C595 B.n353 VSUBS 0.007024f
C596 B.n354 VSUBS 0.01729f
C597 B.n355 VSUBS 0.00417f
C598 B.n356 VSUBS 0.007463f
C599 B.n357 VSUBS 0.007463f
C600 B.n358 VSUBS 0.007463f
C601 B.n359 VSUBS 0.007463f
C602 B.n360 VSUBS 0.007463f
C603 B.n361 VSUBS 0.007463f
C604 B.n362 VSUBS 0.007463f
C605 B.n363 VSUBS 0.007463f
C606 B.n364 VSUBS 0.007463f
C607 B.n365 VSUBS 0.007463f
C608 B.n366 VSUBS 0.007463f
C609 B.n367 VSUBS 0.007463f
C610 B.t5 VSUBS 0.42727f
C611 B.t4 VSUBS 0.451566f
C612 B.t3 VSUBS 1.69344f
C613 B.n368 VSUBS 0.241918f
C614 B.n369 VSUBS 0.077609f
C615 B.n370 VSUBS 0.01729f
C616 B.n371 VSUBS 0.00417f
C617 B.n372 VSUBS 0.007463f
C618 B.n373 VSUBS 0.007463f
C619 B.n374 VSUBS 0.007463f
C620 B.n375 VSUBS 0.007463f
C621 B.n376 VSUBS 0.007463f
C622 B.n377 VSUBS 0.007463f
C623 B.n378 VSUBS 0.007463f
C624 B.n379 VSUBS 0.007463f
C625 B.n380 VSUBS 0.007463f
C626 B.n381 VSUBS 0.007463f
C627 B.n382 VSUBS 0.007463f
C628 B.n383 VSUBS 0.007463f
C629 B.n384 VSUBS 0.007463f
C630 B.n385 VSUBS 0.007463f
C631 B.n386 VSUBS 0.007463f
C632 B.n387 VSUBS 0.007463f
C633 B.n388 VSUBS 0.007463f
C634 B.n389 VSUBS 0.007463f
C635 B.n390 VSUBS 0.007463f
C636 B.n391 VSUBS 0.007463f
C637 B.n392 VSUBS 0.007463f
C638 B.n393 VSUBS 0.007463f
C639 B.n394 VSUBS 0.007463f
C640 B.n395 VSUBS 0.007463f
C641 B.n396 VSUBS 0.007463f
C642 B.n397 VSUBS 0.007463f
C643 B.n398 VSUBS 0.007463f
C644 B.n399 VSUBS 0.007463f
C645 B.n400 VSUBS 0.007463f
C646 B.n401 VSUBS 0.007463f
C647 B.n402 VSUBS 0.007463f
C648 B.n403 VSUBS 0.007463f
C649 B.n404 VSUBS 0.007463f
C650 B.n405 VSUBS 0.007463f
C651 B.n406 VSUBS 0.007463f
C652 B.n407 VSUBS 0.007463f
C653 B.n408 VSUBS 0.007463f
C654 B.n409 VSUBS 0.007463f
C655 B.n410 VSUBS 0.007463f
C656 B.n411 VSUBS 0.007463f
C657 B.n412 VSUBS 0.007463f
C658 B.n413 VSUBS 0.007463f
C659 B.n414 VSUBS 0.007463f
C660 B.n415 VSUBS 0.007463f
C661 B.n416 VSUBS 0.007463f
C662 B.n417 VSUBS 0.007463f
C663 B.n418 VSUBS 0.007463f
C664 B.n419 VSUBS 0.007463f
C665 B.n420 VSUBS 0.007463f
C666 B.n421 VSUBS 0.007463f
C667 B.n422 VSUBS 0.007463f
C668 B.n423 VSUBS 0.007463f
C669 B.n424 VSUBS 0.007463f
C670 B.n425 VSUBS 0.007463f
C671 B.n426 VSUBS 0.007463f
C672 B.n427 VSUBS 0.007463f
C673 B.n428 VSUBS 0.007463f
C674 B.n429 VSUBS 0.007463f
C675 B.n430 VSUBS 0.007463f
C676 B.n431 VSUBS 0.007463f
C677 B.n432 VSUBS 0.007463f
C678 B.n433 VSUBS 0.007463f
C679 B.n434 VSUBS 0.018745f
C680 B.n435 VSUBS 0.017932f
C681 B.n436 VSUBS 0.018943f
C682 B.n437 VSUBS 0.007463f
C683 B.n438 VSUBS 0.007463f
C684 B.n439 VSUBS 0.007463f
C685 B.n440 VSUBS 0.007463f
C686 B.n441 VSUBS 0.007463f
C687 B.n442 VSUBS 0.007463f
C688 B.n443 VSUBS 0.007463f
C689 B.n444 VSUBS 0.007463f
C690 B.n445 VSUBS 0.007463f
C691 B.n446 VSUBS 0.007463f
C692 B.n447 VSUBS 0.007463f
C693 B.n448 VSUBS 0.007463f
C694 B.n449 VSUBS 0.007463f
C695 B.n450 VSUBS 0.007463f
C696 B.n451 VSUBS 0.007463f
C697 B.n452 VSUBS 0.007463f
C698 B.n453 VSUBS 0.007463f
C699 B.n454 VSUBS 0.007463f
C700 B.n455 VSUBS 0.007463f
C701 B.n456 VSUBS 0.007463f
C702 B.n457 VSUBS 0.007463f
C703 B.n458 VSUBS 0.007463f
C704 B.n459 VSUBS 0.007463f
C705 B.n460 VSUBS 0.007463f
C706 B.n461 VSUBS 0.007463f
C707 B.n462 VSUBS 0.007463f
C708 B.n463 VSUBS 0.007463f
C709 B.n464 VSUBS 0.007463f
C710 B.n465 VSUBS 0.007463f
C711 B.n466 VSUBS 0.007463f
C712 B.n467 VSUBS 0.007463f
C713 B.n468 VSUBS 0.007463f
C714 B.n469 VSUBS 0.007463f
C715 B.n470 VSUBS 0.007463f
C716 B.n471 VSUBS 0.007463f
C717 B.n472 VSUBS 0.007463f
C718 B.n473 VSUBS 0.007463f
C719 B.n474 VSUBS 0.007463f
C720 B.n475 VSUBS 0.007463f
C721 B.n476 VSUBS 0.007463f
C722 B.n477 VSUBS 0.007463f
C723 B.n478 VSUBS 0.007463f
C724 B.n479 VSUBS 0.007463f
C725 B.n480 VSUBS 0.007463f
C726 B.n481 VSUBS 0.007463f
C727 B.n482 VSUBS 0.007463f
C728 B.n483 VSUBS 0.007463f
C729 B.n484 VSUBS 0.007463f
C730 B.n485 VSUBS 0.007463f
C731 B.n486 VSUBS 0.007463f
C732 B.n487 VSUBS 0.007463f
C733 B.n488 VSUBS 0.007463f
C734 B.n489 VSUBS 0.007463f
C735 B.n490 VSUBS 0.007463f
C736 B.n491 VSUBS 0.007463f
C737 B.n492 VSUBS 0.007463f
C738 B.n493 VSUBS 0.007463f
C739 B.n494 VSUBS 0.007463f
C740 B.n495 VSUBS 0.007463f
C741 B.n496 VSUBS 0.007463f
C742 B.n497 VSUBS 0.007463f
C743 B.n498 VSUBS 0.007463f
C744 B.n499 VSUBS 0.007463f
C745 B.n500 VSUBS 0.007463f
C746 B.n501 VSUBS 0.007463f
C747 B.n502 VSUBS 0.007463f
C748 B.n503 VSUBS 0.007463f
C749 B.n504 VSUBS 0.007463f
C750 B.n505 VSUBS 0.007463f
C751 B.n506 VSUBS 0.007463f
C752 B.n507 VSUBS 0.007463f
C753 B.n508 VSUBS 0.007463f
C754 B.n509 VSUBS 0.007463f
C755 B.n510 VSUBS 0.007463f
C756 B.n511 VSUBS 0.007463f
C757 B.n512 VSUBS 0.007463f
C758 B.n513 VSUBS 0.007463f
C759 B.n514 VSUBS 0.007463f
C760 B.n515 VSUBS 0.007463f
C761 B.n516 VSUBS 0.007463f
C762 B.n517 VSUBS 0.007463f
C763 B.n518 VSUBS 0.007463f
C764 B.n519 VSUBS 0.007463f
C765 B.n520 VSUBS 0.007463f
C766 B.n521 VSUBS 0.007463f
C767 B.n522 VSUBS 0.007463f
C768 B.n523 VSUBS 0.007463f
C769 B.n524 VSUBS 0.007463f
C770 B.n525 VSUBS 0.007463f
C771 B.n526 VSUBS 0.007463f
C772 B.n527 VSUBS 0.007463f
C773 B.n528 VSUBS 0.007463f
C774 B.n529 VSUBS 0.007463f
C775 B.n530 VSUBS 0.007463f
C776 B.n531 VSUBS 0.007463f
C777 B.n532 VSUBS 0.007463f
C778 B.n533 VSUBS 0.007463f
C779 B.n534 VSUBS 0.007463f
C780 B.n535 VSUBS 0.007463f
C781 B.n536 VSUBS 0.007463f
C782 B.n537 VSUBS 0.007463f
C783 B.n538 VSUBS 0.007463f
C784 B.n539 VSUBS 0.007463f
C785 B.n540 VSUBS 0.007463f
C786 B.n541 VSUBS 0.007463f
C787 B.n542 VSUBS 0.007463f
C788 B.n543 VSUBS 0.007463f
C789 B.n544 VSUBS 0.007463f
C790 B.n545 VSUBS 0.007463f
C791 B.n546 VSUBS 0.007463f
C792 B.n547 VSUBS 0.007463f
C793 B.n548 VSUBS 0.007463f
C794 B.n549 VSUBS 0.007463f
C795 B.n550 VSUBS 0.007463f
C796 B.n551 VSUBS 0.007463f
C797 B.n552 VSUBS 0.007463f
C798 B.n553 VSUBS 0.007463f
C799 B.n554 VSUBS 0.007463f
C800 B.n555 VSUBS 0.007463f
C801 B.n556 VSUBS 0.007463f
C802 B.n557 VSUBS 0.007463f
C803 B.n558 VSUBS 0.007463f
C804 B.n559 VSUBS 0.007463f
C805 B.n560 VSUBS 0.007463f
C806 B.n561 VSUBS 0.007463f
C807 B.n562 VSUBS 0.007463f
C808 B.n563 VSUBS 0.007463f
C809 B.n564 VSUBS 0.007463f
C810 B.n565 VSUBS 0.007463f
C811 B.n566 VSUBS 0.007463f
C812 B.n567 VSUBS 0.007463f
C813 B.n568 VSUBS 0.007463f
C814 B.n569 VSUBS 0.007463f
C815 B.n570 VSUBS 0.007463f
C816 B.n571 VSUBS 0.007463f
C817 B.n572 VSUBS 0.007463f
C818 B.n573 VSUBS 0.007463f
C819 B.n574 VSUBS 0.007463f
C820 B.n575 VSUBS 0.007463f
C821 B.n576 VSUBS 0.007463f
C822 B.n577 VSUBS 0.007463f
C823 B.n578 VSUBS 0.007463f
C824 B.n579 VSUBS 0.007463f
C825 B.n580 VSUBS 0.007463f
C826 B.n581 VSUBS 0.007463f
C827 B.n582 VSUBS 0.007463f
C828 B.n583 VSUBS 0.007463f
C829 B.n584 VSUBS 0.007463f
C830 B.n585 VSUBS 0.007463f
C831 B.n586 VSUBS 0.007463f
C832 B.n587 VSUBS 0.007463f
C833 B.n588 VSUBS 0.007463f
C834 B.n589 VSUBS 0.007463f
C835 B.n590 VSUBS 0.007463f
C836 B.n591 VSUBS 0.007463f
C837 B.n592 VSUBS 0.007463f
C838 B.n593 VSUBS 0.007463f
C839 B.n594 VSUBS 0.007463f
C840 B.n595 VSUBS 0.007463f
C841 B.n596 VSUBS 0.007463f
C842 B.n597 VSUBS 0.007463f
C843 B.n598 VSUBS 0.007463f
C844 B.n599 VSUBS 0.01813f
C845 B.n600 VSUBS 0.01813f
C846 B.n601 VSUBS 0.018745f
C847 B.n602 VSUBS 0.007463f
C848 B.n603 VSUBS 0.007463f
C849 B.n604 VSUBS 0.007463f
C850 B.n605 VSUBS 0.007463f
C851 B.n606 VSUBS 0.007463f
C852 B.n607 VSUBS 0.007463f
C853 B.n608 VSUBS 0.007463f
C854 B.n609 VSUBS 0.007463f
C855 B.n610 VSUBS 0.007463f
C856 B.n611 VSUBS 0.007463f
C857 B.n612 VSUBS 0.007463f
C858 B.n613 VSUBS 0.007463f
C859 B.n614 VSUBS 0.007463f
C860 B.n615 VSUBS 0.007463f
C861 B.n616 VSUBS 0.007463f
C862 B.n617 VSUBS 0.007463f
C863 B.n618 VSUBS 0.007463f
C864 B.n619 VSUBS 0.007463f
C865 B.n620 VSUBS 0.007463f
C866 B.n621 VSUBS 0.007463f
C867 B.n622 VSUBS 0.007463f
C868 B.n623 VSUBS 0.007463f
C869 B.n624 VSUBS 0.007463f
C870 B.n625 VSUBS 0.007463f
C871 B.n626 VSUBS 0.007463f
C872 B.n627 VSUBS 0.007463f
C873 B.n628 VSUBS 0.007463f
C874 B.n629 VSUBS 0.007463f
C875 B.n630 VSUBS 0.007463f
C876 B.n631 VSUBS 0.007463f
C877 B.n632 VSUBS 0.007463f
C878 B.n633 VSUBS 0.007463f
C879 B.n634 VSUBS 0.007463f
C880 B.n635 VSUBS 0.007463f
C881 B.n636 VSUBS 0.007463f
C882 B.n637 VSUBS 0.007463f
C883 B.n638 VSUBS 0.007463f
C884 B.n639 VSUBS 0.007463f
C885 B.n640 VSUBS 0.007463f
C886 B.n641 VSUBS 0.007463f
C887 B.n642 VSUBS 0.007463f
C888 B.n643 VSUBS 0.007463f
C889 B.n644 VSUBS 0.007463f
C890 B.n645 VSUBS 0.007463f
C891 B.n646 VSUBS 0.007463f
C892 B.n647 VSUBS 0.007463f
C893 B.n648 VSUBS 0.007463f
C894 B.n649 VSUBS 0.007463f
C895 B.n650 VSUBS 0.007463f
C896 B.n651 VSUBS 0.007463f
C897 B.n652 VSUBS 0.007463f
C898 B.n653 VSUBS 0.007463f
C899 B.n654 VSUBS 0.007463f
C900 B.n655 VSUBS 0.007463f
C901 B.n656 VSUBS 0.007463f
C902 B.n657 VSUBS 0.007463f
C903 B.n658 VSUBS 0.007463f
C904 B.n659 VSUBS 0.007463f
C905 B.n660 VSUBS 0.007463f
C906 B.n661 VSUBS 0.007463f
C907 B.n662 VSUBS 0.007463f
C908 B.n663 VSUBS 0.007024f
C909 B.n664 VSUBS 0.01729f
C910 B.n665 VSUBS 0.00417f
C911 B.n666 VSUBS 0.007463f
C912 B.n667 VSUBS 0.007463f
C913 B.n668 VSUBS 0.007463f
C914 B.n669 VSUBS 0.007463f
C915 B.n670 VSUBS 0.007463f
C916 B.n671 VSUBS 0.007463f
C917 B.n672 VSUBS 0.007463f
C918 B.n673 VSUBS 0.007463f
C919 B.n674 VSUBS 0.007463f
C920 B.n675 VSUBS 0.007463f
C921 B.n676 VSUBS 0.007463f
C922 B.n677 VSUBS 0.007463f
C923 B.n678 VSUBS 0.00417f
C924 B.n679 VSUBS 0.007463f
C925 B.n680 VSUBS 0.007463f
C926 B.n681 VSUBS 0.007024f
C927 B.n682 VSUBS 0.007463f
C928 B.n683 VSUBS 0.007463f
C929 B.n684 VSUBS 0.007463f
C930 B.n685 VSUBS 0.007463f
C931 B.n686 VSUBS 0.007463f
C932 B.n687 VSUBS 0.007463f
C933 B.n688 VSUBS 0.007463f
C934 B.n689 VSUBS 0.007463f
C935 B.n690 VSUBS 0.007463f
C936 B.n691 VSUBS 0.007463f
C937 B.n692 VSUBS 0.007463f
C938 B.n693 VSUBS 0.007463f
C939 B.n694 VSUBS 0.007463f
C940 B.n695 VSUBS 0.007463f
C941 B.n696 VSUBS 0.007463f
C942 B.n697 VSUBS 0.007463f
C943 B.n698 VSUBS 0.007463f
C944 B.n699 VSUBS 0.007463f
C945 B.n700 VSUBS 0.007463f
C946 B.n701 VSUBS 0.007463f
C947 B.n702 VSUBS 0.007463f
C948 B.n703 VSUBS 0.007463f
C949 B.n704 VSUBS 0.007463f
C950 B.n705 VSUBS 0.007463f
C951 B.n706 VSUBS 0.007463f
C952 B.n707 VSUBS 0.007463f
C953 B.n708 VSUBS 0.007463f
C954 B.n709 VSUBS 0.007463f
C955 B.n710 VSUBS 0.007463f
C956 B.n711 VSUBS 0.007463f
C957 B.n712 VSUBS 0.007463f
C958 B.n713 VSUBS 0.007463f
C959 B.n714 VSUBS 0.007463f
C960 B.n715 VSUBS 0.007463f
C961 B.n716 VSUBS 0.007463f
C962 B.n717 VSUBS 0.007463f
C963 B.n718 VSUBS 0.007463f
C964 B.n719 VSUBS 0.007463f
C965 B.n720 VSUBS 0.007463f
C966 B.n721 VSUBS 0.007463f
C967 B.n722 VSUBS 0.007463f
C968 B.n723 VSUBS 0.007463f
C969 B.n724 VSUBS 0.007463f
C970 B.n725 VSUBS 0.007463f
C971 B.n726 VSUBS 0.007463f
C972 B.n727 VSUBS 0.007463f
C973 B.n728 VSUBS 0.007463f
C974 B.n729 VSUBS 0.007463f
C975 B.n730 VSUBS 0.007463f
C976 B.n731 VSUBS 0.007463f
C977 B.n732 VSUBS 0.007463f
C978 B.n733 VSUBS 0.007463f
C979 B.n734 VSUBS 0.007463f
C980 B.n735 VSUBS 0.007463f
C981 B.n736 VSUBS 0.007463f
C982 B.n737 VSUBS 0.007463f
C983 B.n738 VSUBS 0.007463f
C984 B.n739 VSUBS 0.007463f
C985 B.n740 VSUBS 0.007463f
C986 B.n741 VSUBS 0.007463f
C987 B.n742 VSUBS 0.018745f
C988 B.n743 VSUBS 0.01813f
C989 B.n744 VSUBS 0.01813f
C990 B.n745 VSUBS 0.007463f
C991 B.n746 VSUBS 0.007463f
C992 B.n747 VSUBS 0.007463f
C993 B.n748 VSUBS 0.007463f
C994 B.n749 VSUBS 0.007463f
C995 B.n750 VSUBS 0.007463f
C996 B.n751 VSUBS 0.007463f
C997 B.n752 VSUBS 0.007463f
C998 B.n753 VSUBS 0.007463f
C999 B.n754 VSUBS 0.007463f
C1000 B.n755 VSUBS 0.007463f
C1001 B.n756 VSUBS 0.007463f
C1002 B.n757 VSUBS 0.007463f
C1003 B.n758 VSUBS 0.007463f
C1004 B.n759 VSUBS 0.007463f
C1005 B.n760 VSUBS 0.007463f
C1006 B.n761 VSUBS 0.007463f
C1007 B.n762 VSUBS 0.007463f
C1008 B.n763 VSUBS 0.007463f
C1009 B.n764 VSUBS 0.007463f
C1010 B.n765 VSUBS 0.007463f
C1011 B.n766 VSUBS 0.007463f
C1012 B.n767 VSUBS 0.007463f
C1013 B.n768 VSUBS 0.007463f
C1014 B.n769 VSUBS 0.007463f
C1015 B.n770 VSUBS 0.007463f
C1016 B.n771 VSUBS 0.007463f
C1017 B.n772 VSUBS 0.007463f
C1018 B.n773 VSUBS 0.007463f
C1019 B.n774 VSUBS 0.007463f
C1020 B.n775 VSUBS 0.007463f
C1021 B.n776 VSUBS 0.007463f
C1022 B.n777 VSUBS 0.007463f
C1023 B.n778 VSUBS 0.007463f
C1024 B.n779 VSUBS 0.007463f
C1025 B.n780 VSUBS 0.007463f
C1026 B.n781 VSUBS 0.007463f
C1027 B.n782 VSUBS 0.007463f
C1028 B.n783 VSUBS 0.007463f
C1029 B.n784 VSUBS 0.007463f
C1030 B.n785 VSUBS 0.007463f
C1031 B.n786 VSUBS 0.007463f
C1032 B.n787 VSUBS 0.007463f
C1033 B.n788 VSUBS 0.007463f
C1034 B.n789 VSUBS 0.007463f
C1035 B.n790 VSUBS 0.007463f
C1036 B.n791 VSUBS 0.007463f
C1037 B.n792 VSUBS 0.007463f
C1038 B.n793 VSUBS 0.007463f
C1039 B.n794 VSUBS 0.007463f
C1040 B.n795 VSUBS 0.007463f
C1041 B.n796 VSUBS 0.007463f
C1042 B.n797 VSUBS 0.007463f
C1043 B.n798 VSUBS 0.007463f
C1044 B.n799 VSUBS 0.007463f
C1045 B.n800 VSUBS 0.007463f
C1046 B.n801 VSUBS 0.007463f
C1047 B.n802 VSUBS 0.007463f
C1048 B.n803 VSUBS 0.007463f
C1049 B.n804 VSUBS 0.007463f
C1050 B.n805 VSUBS 0.007463f
C1051 B.n806 VSUBS 0.007463f
C1052 B.n807 VSUBS 0.007463f
C1053 B.n808 VSUBS 0.007463f
C1054 B.n809 VSUBS 0.007463f
C1055 B.n810 VSUBS 0.007463f
C1056 B.n811 VSUBS 0.007463f
C1057 B.n812 VSUBS 0.007463f
C1058 B.n813 VSUBS 0.007463f
C1059 B.n814 VSUBS 0.007463f
C1060 B.n815 VSUBS 0.007463f
C1061 B.n816 VSUBS 0.007463f
C1062 B.n817 VSUBS 0.007463f
C1063 B.n818 VSUBS 0.007463f
C1064 B.n819 VSUBS 0.007463f
C1065 B.n820 VSUBS 0.007463f
C1066 B.n821 VSUBS 0.007463f
C1067 B.n822 VSUBS 0.007463f
C1068 B.n823 VSUBS 0.009738f
C1069 B.n824 VSUBS 0.010374f
C1070 B.n825 VSUBS 0.02063f
.ends

