* NGSPICE file created from diff_pair_sample_1455.ext - technology: sky130A

.subckt diff_pair_sample_1455 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n3400_n1070# sky130_fd_pr__pfet_01v8 ad=0.1989 pd=1.8 as=0 ps=0 w=0.51 l=3.72
X1 VTAIL.t7 VP.t0 VDD1.t3 w_n3400_n1070# sky130_fd_pr__pfet_01v8 ad=0.1989 pd=1.8 as=0.08415 ps=0.84 w=0.51 l=3.72
X2 VDD1.t2 VP.t1 VTAIL.t6 w_n3400_n1070# sky130_fd_pr__pfet_01v8 ad=0.08415 pd=0.84 as=0.1989 ps=1.8 w=0.51 l=3.72
X3 B.t8 B.t6 B.t7 w_n3400_n1070# sky130_fd_pr__pfet_01v8 ad=0.1989 pd=1.8 as=0 ps=0 w=0.51 l=3.72
X4 VDD1.t1 VP.t2 VTAIL.t5 w_n3400_n1070# sky130_fd_pr__pfet_01v8 ad=0.08415 pd=0.84 as=0.1989 ps=1.8 w=0.51 l=3.72
X5 VDD2.t3 VN.t0 VTAIL.t2 w_n3400_n1070# sky130_fd_pr__pfet_01v8 ad=0.08415 pd=0.84 as=0.1989 ps=1.8 w=0.51 l=3.72
X6 VDD2.t2 VN.t1 VTAIL.t3 w_n3400_n1070# sky130_fd_pr__pfet_01v8 ad=0.08415 pd=0.84 as=0.1989 ps=1.8 w=0.51 l=3.72
X7 VTAIL.t1 VN.t2 VDD2.t1 w_n3400_n1070# sky130_fd_pr__pfet_01v8 ad=0.1989 pd=1.8 as=0.08415 ps=0.84 w=0.51 l=3.72
X8 B.t5 B.t3 B.t4 w_n3400_n1070# sky130_fd_pr__pfet_01v8 ad=0.1989 pd=1.8 as=0 ps=0 w=0.51 l=3.72
X9 B.t2 B.t0 B.t1 w_n3400_n1070# sky130_fd_pr__pfet_01v8 ad=0.1989 pd=1.8 as=0 ps=0 w=0.51 l=3.72
X10 VTAIL.t0 VN.t3 VDD2.t0 w_n3400_n1070# sky130_fd_pr__pfet_01v8 ad=0.1989 pd=1.8 as=0.08415 ps=0.84 w=0.51 l=3.72
X11 VTAIL.t4 VP.t3 VDD1.t0 w_n3400_n1070# sky130_fd_pr__pfet_01v8 ad=0.1989 pd=1.8 as=0.08415 ps=0.84 w=0.51 l=3.72
R0 B.n90 B.t8 746.87
R1 B.n96 B.t2 746.87
R2 B.n28 B.t10 746.87
R3 B.n36 B.t4 746.87
R4 B.n91 B.t7 668.323
R5 B.n97 B.t1 668.323
R6 B.n29 B.t11 668.323
R7 B.n37 B.t5 668.323
R8 B.n362 B.n361 585
R9 B.n363 B.n40 585
R10 B.n365 B.n364 585
R11 B.n366 B.n39 585
R12 B.n368 B.n367 585
R13 B.n369 B.n38 585
R14 B.n371 B.n370 585
R15 B.n372 B.n35 585
R16 B.n375 B.n374 585
R17 B.n376 B.n34 585
R18 B.n378 B.n377 585
R19 B.n379 B.n33 585
R20 B.n381 B.n380 585
R21 B.n382 B.n32 585
R22 B.n384 B.n383 585
R23 B.n385 B.n31 585
R24 B.n387 B.n386 585
R25 B.n389 B.n388 585
R26 B.n390 B.n27 585
R27 B.n392 B.n391 585
R28 B.n393 B.n26 585
R29 B.n395 B.n394 585
R30 B.n396 B.n25 585
R31 B.n398 B.n397 585
R32 B.n399 B.n24 585
R33 B.n360 B.n41 585
R34 B.n359 B.n358 585
R35 B.n357 B.n42 585
R36 B.n356 B.n355 585
R37 B.n354 B.n43 585
R38 B.n353 B.n352 585
R39 B.n351 B.n44 585
R40 B.n350 B.n349 585
R41 B.n348 B.n45 585
R42 B.n347 B.n346 585
R43 B.n345 B.n46 585
R44 B.n344 B.n343 585
R45 B.n342 B.n47 585
R46 B.n341 B.n340 585
R47 B.n339 B.n48 585
R48 B.n338 B.n337 585
R49 B.n336 B.n49 585
R50 B.n335 B.n334 585
R51 B.n333 B.n50 585
R52 B.n332 B.n331 585
R53 B.n330 B.n51 585
R54 B.n329 B.n328 585
R55 B.n327 B.n52 585
R56 B.n326 B.n325 585
R57 B.n324 B.n53 585
R58 B.n323 B.n322 585
R59 B.n321 B.n54 585
R60 B.n320 B.n319 585
R61 B.n318 B.n55 585
R62 B.n317 B.n316 585
R63 B.n315 B.n56 585
R64 B.n314 B.n313 585
R65 B.n312 B.n57 585
R66 B.n311 B.n310 585
R67 B.n309 B.n58 585
R68 B.n308 B.n307 585
R69 B.n306 B.n59 585
R70 B.n305 B.n304 585
R71 B.n303 B.n60 585
R72 B.n302 B.n301 585
R73 B.n300 B.n61 585
R74 B.n299 B.n298 585
R75 B.n297 B.n62 585
R76 B.n296 B.n295 585
R77 B.n294 B.n63 585
R78 B.n293 B.n292 585
R79 B.n291 B.n64 585
R80 B.n290 B.n289 585
R81 B.n288 B.n65 585
R82 B.n287 B.n286 585
R83 B.n285 B.n66 585
R84 B.n284 B.n283 585
R85 B.n282 B.n67 585
R86 B.n281 B.n280 585
R87 B.n279 B.n68 585
R88 B.n278 B.n277 585
R89 B.n276 B.n69 585
R90 B.n275 B.n274 585
R91 B.n273 B.n70 585
R92 B.n272 B.n271 585
R93 B.n270 B.n71 585
R94 B.n269 B.n268 585
R95 B.n267 B.n72 585
R96 B.n266 B.n265 585
R97 B.n264 B.n73 585
R98 B.n263 B.n262 585
R99 B.n261 B.n74 585
R100 B.n260 B.n259 585
R101 B.n258 B.n75 585
R102 B.n257 B.n256 585
R103 B.n255 B.n76 585
R104 B.n254 B.n253 585
R105 B.n252 B.n77 585
R106 B.n251 B.n250 585
R107 B.n249 B.n78 585
R108 B.n248 B.n247 585
R109 B.n246 B.n79 585
R110 B.n245 B.n244 585
R111 B.n243 B.n80 585
R112 B.n242 B.n241 585
R113 B.n240 B.n81 585
R114 B.n239 B.n238 585
R115 B.n237 B.n82 585
R116 B.n236 B.n235 585
R117 B.n234 B.n83 585
R118 B.n233 B.n232 585
R119 B.n231 B.n84 585
R120 B.n230 B.n229 585
R121 B.n228 B.n85 585
R122 B.n189 B.n102 585
R123 B.n191 B.n190 585
R124 B.n192 B.n101 585
R125 B.n194 B.n193 585
R126 B.n195 B.n100 585
R127 B.n197 B.n196 585
R128 B.n198 B.n99 585
R129 B.n200 B.n199 585
R130 B.n202 B.n201 585
R131 B.n203 B.n95 585
R132 B.n205 B.n204 585
R133 B.n206 B.n94 585
R134 B.n208 B.n207 585
R135 B.n209 B.n93 585
R136 B.n211 B.n210 585
R137 B.n212 B.n92 585
R138 B.n214 B.n213 585
R139 B.n216 B.n89 585
R140 B.n218 B.n217 585
R141 B.n219 B.n88 585
R142 B.n221 B.n220 585
R143 B.n222 B.n87 585
R144 B.n224 B.n223 585
R145 B.n225 B.n86 585
R146 B.n227 B.n226 585
R147 B.n188 B.n187 585
R148 B.n186 B.n103 585
R149 B.n185 B.n184 585
R150 B.n183 B.n104 585
R151 B.n182 B.n181 585
R152 B.n180 B.n105 585
R153 B.n179 B.n178 585
R154 B.n177 B.n106 585
R155 B.n176 B.n175 585
R156 B.n174 B.n107 585
R157 B.n173 B.n172 585
R158 B.n171 B.n108 585
R159 B.n170 B.n169 585
R160 B.n168 B.n109 585
R161 B.n167 B.n166 585
R162 B.n165 B.n110 585
R163 B.n164 B.n163 585
R164 B.n162 B.n111 585
R165 B.n161 B.n160 585
R166 B.n159 B.n112 585
R167 B.n158 B.n157 585
R168 B.n156 B.n113 585
R169 B.n155 B.n154 585
R170 B.n153 B.n114 585
R171 B.n152 B.n151 585
R172 B.n150 B.n115 585
R173 B.n149 B.n148 585
R174 B.n147 B.n116 585
R175 B.n146 B.n145 585
R176 B.n144 B.n117 585
R177 B.n143 B.n142 585
R178 B.n141 B.n118 585
R179 B.n140 B.n139 585
R180 B.n138 B.n119 585
R181 B.n137 B.n136 585
R182 B.n135 B.n120 585
R183 B.n134 B.n133 585
R184 B.n132 B.n121 585
R185 B.n131 B.n130 585
R186 B.n129 B.n122 585
R187 B.n128 B.n127 585
R188 B.n126 B.n123 585
R189 B.n125 B.n124 585
R190 B.n2 B.n0 585
R191 B.n465 B.n1 585
R192 B.n464 B.n463 585
R193 B.n462 B.n3 585
R194 B.n461 B.n460 585
R195 B.n459 B.n4 585
R196 B.n458 B.n457 585
R197 B.n456 B.n5 585
R198 B.n455 B.n454 585
R199 B.n453 B.n6 585
R200 B.n452 B.n451 585
R201 B.n450 B.n7 585
R202 B.n449 B.n448 585
R203 B.n447 B.n8 585
R204 B.n446 B.n445 585
R205 B.n444 B.n9 585
R206 B.n443 B.n442 585
R207 B.n441 B.n10 585
R208 B.n440 B.n439 585
R209 B.n438 B.n11 585
R210 B.n437 B.n436 585
R211 B.n435 B.n12 585
R212 B.n434 B.n433 585
R213 B.n432 B.n13 585
R214 B.n431 B.n430 585
R215 B.n429 B.n14 585
R216 B.n428 B.n427 585
R217 B.n426 B.n15 585
R218 B.n425 B.n424 585
R219 B.n423 B.n16 585
R220 B.n422 B.n421 585
R221 B.n420 B.n17 585
R222 B.n419 B.n418 585
R223 B.n417 B.n18 585
R224 B.n416 B.n415 585
R225 B.n414 B.n19 585
R226 B.n413 B.n412 585
R227 B.n411 B.n20 585
R228 B.n410 B.n409 585
R229 B.n408 B.n21 585
R230 B.n407 B.n406 585
R231 B.n405 B.n22 585
R232 B.n404 B.n403 585
R233 B.n402 B.n23 585
R234 B.n401 B.n400 585
R235 B.n467 B.n466 585
R236 B.n189 B.n188 492.5
R237 B.n400 B.n399 492.5
R238 B.n226 B.n85 492.5
R239 B.n362 B.n41 492.5
R240 B.n90 B.t6 210.361
R241 B.n96 B.t0 210.361
R242 B.n28 B.t9 210.361
R243 B.n36 B.t3 210.361
R244 B.n188 B.n103 163.367
R245 B.n184 B.n103 163.367
R246 B.n184 B.n183 163.367
R247 B.n183 B.n182 163.367
R248 B.n182 B.n105 163.367
R249 B.n178 B.n105 163.367
R250 B.n178 B.n177 163.367
R251 B.n177 B.n176 163.367
R252 B.n176 B.n107 163.367
R253 B.n172 B.n107 163.367
R254 B.n172 B.n171 163.367
R255 B.n171 B.n170 163.367
R256 B.n170 B.n109 163.367
R257 B.n166 B.n109 163.367
R258 B.n166 B.n165 163.367
R259 B.n165 B.n164 163.367
R260 B.n164 B.n111 163.367
R261 B.n160 B.n111 163.367
R262 B.n160 B.n159 163.367
R263 B.n159 B.n158 163.367
R264 B.n158 B.n113 163.367
R265 B.n154 B.n113 163.367
R266 B.n154 B.n153 163.367
R267 B.n153 B.n152 163.367
R268 B.n152 B.n115 163.367
R269 B.n148 B.n115 163.367
R270 B.n148 B.n147 163.367
R271 B.n147 B.n146 163.367
R272 B.n146 B.n117 163.367
R273 B.n142 B.n117 163.367
R274 B.n142 B.n141 163.367
R275 B.n141 B.n140 163.367
R276 B.n140 B.n119 163.367
R277 B.n136 B.n119 163.367
R278 B.n136 B.n135 163.367
R279 B.n135 B.n134 163.367
R280 B.n134 B.n121 163.367
R281 B.n130 B.n121 163.367
R282 B.n130 B.n129 163.367
R283 B.n129 B.n128 163.367
R284 B.n128 B.n123 163.367
R285 B.n124 B.n123 163.367
R286 B.n124 B.n2 163.367
R287 B.n466 B.n2 163.367
R288 B.n466 B.n465 163.367
R289 B.n465 B.n464 163.367
R290 B.n464 B.n3 163.367
R291 B.n460 B.n3 163.367
R292 B.n460 B.n459 163.367
R293 B.n459 B.n458 163.367
R294 B.n458 B.n5 163.367
R295 B.n454 B.n5 163.367
R296 B.n454 B.n453 163.367
R297 B.n453 B.n452 163.367
R298 B.n452 B.n7 163.367
R299 B.n448 B.n7 163.367
R300 B.n448 B.n447 163.367
R301 B.n447 B.n446 163.367
R302 B.n446 B.n9 163.367
R303 B.n442 B.n9 163.367
R304 B.n442 B.n441 163.367
R305 B.n441 B.n440 163.367
R306 B.n440 B.n11 163.367
R307 B.n436 B.n11 163.367
R308 B.n436 B.n435 163.367
R309 B.n435 B.n434 163.367
R310 B.n434 B.n13 163.367
R311 B.n430 B.n13 163.367
R312 B.n430 B.n429 163.367
R313 B.n429 B.n428 163.367
R314 B.n428 B.n15 163.367
R315 B.n424 B.n15 163.367
R316 B.n424 B.n423 163.367
R317 B.n423 B.n422 163.367
R318 B.n422 B.n17 163.367
R319 B.n418 B.n17 163.367
R320 B.n418 B.n417 163.367
R321 B.n417 B.n416 163.367
R322 B.n416 B.n19 163.367
R323 B.n412 B.n19 163.367
R324 B.n412 B.n411 163.367
R325 B.n411 B.n410 163.367
R326 B.n410 B.n21 163.367
R327 B.n406 B.n21 163.367
R328 B.n406 B.n405 163.367
R329 B.n405 B.n404 163.367
R330 B.n404 B.n23 163.367
R331 B.n400 B.n23 163.367
R332 B.n190 B.n189 163.367
R333 B.n190 B.n101 163.367
R334 B.n194 B.n101 163.367
R335 B.n195 B.n194 163.367
R336 B.n196 B.n195 163.367
R337 B.n196 B.n99 163.367
R338 B.n200 B.n99 163.367
R339 B.n201 B.n200 163.367
R340 B.n201 B.n95 163.367
R341 B.n205 B.n95 163.367
R342 B.n206 B.n205 163.367
R343 B.n207 B.n206 163.367
R344 B.n207 B.n93 163.367
R345 B.n211 B.n93 163.367
R346 B.n212 B.n211 163.367
R347 B.n213 B.n212 163.367
R348 B.n213 B.n89 163.367
R349 B.n218 B.n89 163.367
R350 B.n219 B.n218 163.367
R351 B.n220 B.n219 163.367
R352 B.n220 B.n87 163.367
R353 B.n224 B.n87 163.367
R354 B.n225 B.n224 163.367
R355 B.n226 B.n225 163.367
R356 B.n230 B.n85 163.367
R357 B.n231 B.n230 163.367
R358 B.n232 B.n231 163.367
R359 B.n232 B.n83 163.367
R360 B.n236 B.n83 163.367
R361 B.n237 B.n236 163.367
R362 B.n238 B.n237 163.367
R363 B.n238 B.n81 163.367
R364 B.n242 B.n81 163.367
R365 B.n243 B.n242 163.367
R366 B.n244 B.n243 163.367
R367 B.n244 B.n79 163.367
R368 B.n248 B.n79 163.367
R369 B.n249 B.n248 163.367
R370 B.n250 B.n249 163.367
R371 B.n250 B.n77 163.367
R372 B.n254 B.n77 163.367
R373 B.n255 B.n254 163.367
R374 B.n256 B.n255 163.367
R375 B.n256 B.n75 163.367
R376 B.n260 B.n75 163.367
R377 B.n261 B.n260 163.367
R378 B.n262 B.n261 163.367
R379 B.n262 B.n73 163.367
R380 B.n266 B.n73 163.367
R381 B.n267 B.n266 163.367
R382 B.n268 B.n267 163.367
R383 B.n268 B.n71 163.367
R384 B.n272 B.n71 163.367
R385 B.n273 B.n272 163.367
R386 B.n274 B.n273 163.367
R387 B.n274 B.n69 163.367
R388 B.n278 B.n69 163.367
R389 B.n279 B.n278 163.367
R390 B.n280 B.n279 163.367
R391 B.n280 B.n67 163.367
R392 B.n284 B.n67 163.367
R393 B.n285 B.n284 163.367
R394 B.n286 B.n285 163.367
R395 B.n286 B.n65 163.367
R396 B.n290 B.n65 163.367
R397 B.n291 B.n290 163.367
R398 B.n292 B.n291 163.367
R399 B.n292 B.n63 163.367
R400 B.n296 B.n63 163.367
R401 B.n297 B.n296 163.367
R402 B.n298 B.n297 163.367
R403 B.n298 B.n61 163.367
R404 B.n302 B.n61 163.367
R405 B.n303 B.n302 163.367
R406 B.n304 B.n303 163.367
R407 B.n304 B.n59 163.367
R408 B.n308 B.n59 163.367
R409 B.n309 B.n308 163.367
R410 B.n310 B.n309 163.367
R411 B.n310 B.n57 163.367
R412 B.n314 B.n57 163.367
R413 B.n315 B.n314 163.367
R414 B.n316 B.n315 163.367
R415 B.n316 B.n55 163.367
R416 B.n320 B.n55 163.367
R417 B.n321 B.n320 163.367
R418 B.n322 B.n321 163.367
R419 B.n322 B.n53 163.367
R420 B.n326 B.n53 163.367
R421 B.n327 B.n326 163.367
R422 B.n328 B.n327 163.367
R423 B.n328 B.n51 163.367
R424 B.n332 B.n51 163.367
R425 B.n333 B.n332 163.367
R426 B.n334 B.n333 163.367
R427 B.n334 B.n49 163.367
R428 B.n338 B.n49 163.367
R429 B.n339 B.n338 163.367
R430 B.n340 B.n339 163.367
R431 B.n340 B.n47 163.367
R432 B.n344 B.n47 163.367
R433 B.n345 B.n344 163.367
R434 B.n346 B.n345 163.367
R435 B.n346 B.n45 163.367
R436 B.n350 B.n45 163.367
R437 B.n351 B.n350 163.367
R438 B.n352 B.n351 163.367
R439 B.n352 B.n43 163.367
R440 B.n356 B.n43 163.367
R441 B.n357 B.n356 163.367
R442 B.n358 B.n357 163.367
R443 B.n358 B.n41 163.367
R444 B.n399 B.n398 163.367
R445 B.n398 B.n25 163.367
R446 B.n394 B.n25 163.367
R447 B.n394 B.n393 163.367
R448 B.n393 B.n392 163.367
R449 B.n392 B.n27 163.367
R450 B.n388 B.n27 163.367
R451 B.n388 B.n387 163.367
R452 B.n387 B.n31 163.367
R453 B.n383 B.n31 163.367
R454 B.n383 B.n382 163.367
R455 B.n382 B.n381 163.367
R456 B.n381 B.n33 163.367
R457 B.n377 B.n33 163.367
R458 B.n377 B.n376 163.367
R459 B.n376 B.n375 163.367
R460 B.n375 B.n35 163.367
R461 B.n370 B.n35 163.367
R462 B.n370 B.n369 163.367
R463 B.n369 B.n368 163.367
R464 B.n368 B.n39 163.367
R465 B.n364 B.n39 163.367
R466 B.n364 B.n363 163.367
R467 B.n363 B.n362 163.367
R468 B.n91 B.n90 78.546
R469 B.n97 B.n96 78.546
R470 B.n29 B.n28 78.546
R471 B.n37 B.n36 78.546
R472 B.n215 B.n91 59.5399
R473 B.n98 B.n97 59.5399
R474 B.n30 B.n29 59.5399
R475 B.n373 B.n37 59.5399
R476 B.n401 B.n24 32.0005
R477 B.n361 B.n360 32.0005
R478 B.n228 B.n227 32.0005
R479 B.n187 B.n102 32.0005
R480 B B.n467 18.0485
R481 B.n397 B.n24 10.6151
R482 B.n397 B.n396 10.6151
R483 B.n396 B.n395 10.6151
R484 B.n395 B.n26 10.6151
R485 B.n391 B.n26 10.6151
R486 B.n391 B.n390 10.6151
R487 B.n390 B.n389 10.6151
R488 B.n386 B.n385 10.6151
R489 B.n385 B.n384 10.6151
R490 B.n384 B.n32 10.6151
R491 B.n380 B.n32 10.6151
R492 B.n380 B.n379 10.6151
R493 B.n379 B.n378 10.6151
R494 B.n378 B.n34 10.6151
R495 B.n374 B.n34 10.6151
R496 B.n372 B.n371 10.6151
R497 B.n371 B.n38 10.6151
R498 B.n367 B.n38 10.6151
R499 B.n367 B.n366 10.6151
R500 B.n366 B.n365 10.6151
R501 B.n365 B.n40 10.6151
R502 B.n361 B.n40 10.6151
R503 B.n229 B.n228 10.6151
R504 B.n229 B.n84 10.6151
R505 B.n233 B.n84 10.6151
R506 B.n234 B.n233 10.6151
R507 B.n235 B.n234 10.6151
R508 B.n235 B.n82 10.6151
R509 B.n239 B.n82 10.6151
R510 B.n240 B.n239 10.6151
R511 B.n241 B.n240 10.6151
R512 B.n241 B.n80 10.6151
R513 B.n245 B.n80 10.6151
R514 B.n246 B.n245 10.6151
R515 B.n247 B.n246 10.6151
R516 B.n247 B.n78 10.6151
R517 B.n251 B.n78 10.6151
R518 B.n252 B.n251 10.6151
R519 B.n253 B.n252 10.6151
R520 B.n253 B.n76 10.6151
R521 B.n257 B.n76 10.6151
R522 B.n258 B.n257 10.6151
R523 B.n259 B.n258 10.6151
R524 B.n259 B.n74 10.6151
R525 B.n263 B.n74 10.6151
R526 B.n264 B.n263 10.6151
R527 B.n265 B.n264 10.6151
R528 B.n265 B.n72 10.6151
R529 B.n269 B.n72 10.6151
R530 B.n270 B.n269 10.6151
R531 B.n271 B.n270 10.6151
R532 B.n271 B.n70 10.6151
R533 B.n275 B.n70 10.6151
R534 B.n276 B.n275 10.6151
R535 B.n277 B.n276 10.6151
R536 B.n277 B.n68 10.6151
R537 B.n281 B.n68 10.6151
R538 B.n282 B.n281 10.6151
R539 B.n283 B.n282 10.6151
R540 B.n283 B.n66 10.6151
R541 B.n287 B.n66 10.6151
R542 B.n288 B.n287 10.6151
R543 B.n289 B.n288 10.6151
R544 B.n289 B.n64 10.6151
R545 B.n293 B.n64 10.6151
R546 B.n294 B.n293 10.6151
R547 B.n295 B.n294 10.6151
R548 B.n295 B.n62 10.6151
R549 B.n299 B.n62 10.6151
R550 B.n300 B.n299 10.6151
R551 B.n301 B.n300 10.6151
R552 B.n301 B.n60 10.6151
R553 B.n305 B.n60 10.6151
R554 B.n306 B.n305 10.6151
R555 B.n307 B.n306 10.6151
R556 B.n307 B.n58 10.6151
R557 B.n311 B.n58 10.6151
R558 B.n312 B.n311 10.6151
R559 B.n313 B.n312 10.6151
R560 B.n313 B.n56 10.6151
R561 B.n317 B.n56 10.6151
R562 B.n318 B.n317 10.6151
R563 B.n319 B.n318 10.6151
R564 B.n319 B.n54 10.6151
R565 B.n323 B.n54 10.6151
R566 B.n324 B.n323 10.6151
R567 B.n325 B.n324 10.6151
R568 B.n325 B.n52 10.6151
R569 B.n329 B.n52 10.6151
R570 B.n330 B.n329 10.6151
R571 B.n331 B.n330 10.6151
R572 B.n331 B.n50 10.6151
R573 B.n335 B.n50 10.6151
R574 B.n336 B.n335 10.6151
R575 B.n337 B.n336 10.6151
R576 B.n337 B.n48 10.6151
R577 B.n341 B.n48 10.6151
R578 B.n342 B.n341 10.6151
R579 B.n343 B.n342 10.6151
R580 B.n343 B.n46 10.6151
R581 B.n347 B.n46 10.6151
R582 B.n348 B.n347 10.6151
R583 B.n349 B.n348 10.6151
R584 B.n349 B.n44 10.6151
R585 B.n353 B.n44 10.6151
R586 B.n354 B.n353 10.6151
R587 B.n355 B.n354 10.6151
R588 B.n355 B.n42 10.6151
R589 B.n359 B.n42 10.6151
R590 B.n360 B.n359 10.6151
R591 B.n191 B.n102 10.6151
R592 B.n192 B.n191 10.6151
R593 B.n193 B.n192 10.6151
R594 B.n193 B.n100 10.6151
R595 B.n197 B.n100 10.6151
R596 B.n198 B.n197 10.6151
R597 B.n199 B.n198 10.6151
R598 B.n203 B.n202 10.6151
R599 B.n204 B.n203 10.6151
R600 B.n204 B.n94 10.6151
R601 B.n208 B.n94 10.6151
R602 B.n209 B.n208 10.6151
R603 B.n210 B.n209 10.6151
R604 B.n210 B.n92 10.6151
R605 B.n214 B.n92 10.6151
R606 B.n217 B.n216 10.6151
R607 B.n217 B.n88 10.6151
R608 B.n221 B.n88 10.6151
R609 B.n222 B.n221 10.6151
R610 B.n223 B.n222 10.6151
R611 B.n223 B.n86 10.6151
R612 B.n227 B.n86 10.6151
R613 B.n187 B.n186 10.6151
R614 B.n186 B.n185 10.6151
R615 B.n185 B.n104 10.6151
R616 B.n181 B.n104 10.6151
R617 B.n181 B.n180 10.6151
R618 B.n180 B.n179 10.6151
R619 B.n179 B.n106 10.6151
R620 B.n175 B.n106 10.6151
R621 B.n175 B.n174 10.6151
R622 B.n174 B.n173 10.6151
R623 B.n173 B.n108 10.6151
R624 B.n169 B.n108 10.6151
R625 B.n169 B.n168 10.6151
R626 B.n168 B.n167 10.6151
R627 B.n167 B.n110 10.6151
R628 B.n163 B.n110 10.6151
R629 B.n163 B.n162 10.6151
R630 B.n162 B.n161 10.6151
R631 B.n161 B.n112 10.6151
R632 B.n157 B.n112 10.6151
R633 B.n157 B.n156 10.6151
R634 B.n156 B.n155 10.6151
R635 B.n155 B.n114 10.6151
R636 B.n151 B.n114 10.6151
R637 B.n151 B.n150 10.6151
R638 B.n150 B.n149 10.6151
R639 B.n149 B.n116 10.6151
R640 B.n145 B.n116 10.6151
R641 B.n145 B.n144 10.6151
R642 B.n144 B.n143 10.6151
R643 B.n143 B.n118 10.6151
R644 B.n139 B.n118 10.6151
R645 B.n139 B.n138 10.6151
R646 B.n138 B.n137 10.6151
R647 B.n137 B.n120 10.6151
R648 B.n133 B.n120 10.6151
R649 B.n133 B.n132 10.6151
R650 B.n132 B.n131 10.6151
R651 B.n131 B.n122 10.6151
R652 B.n127 B.n122 10.6151
R653 B.n127 B.n126 10.6151
R654 B.n126 B.n125 10.6151
R655 B.n125 B.n0 10.6151
R656 B.n463 B.n1 10.6151
R657 B.n463 B.n462 10.6151
R658 B.n462 B.n461 10.6151
R659 B.n461 B.n4 10.6151
R660 B.n457 B.n4 10.6151
R661 B.n457 B.n456 10.6151
R662 B.n456 B.n455 10.6151
R663 B.n455 B.n6 10.6151
R664 B.n451 B.n6 10.6151
R665 B.n451 B.n450 10.6151
R666 B.n450 B.n449 10.6151
R667 B.n449 B.n8 10.6151
R668 B.n445 B.n8 10.6151
R669 B.n445 B.n444 10.6151
R670 B.n444 B.n443 10.6151
R671 B.n443 B.n10 10.6151
R672 B.n439 B.n10 10.6151
R673 B.n439 B.n438 10.6151
R674 B.n438 B.n437 10.6151
R675 B.n437 B.n12 10.6151
R676 B.n433 B.n12 10.6151
R677 B.n433 B.n432 10.6151
R678 B.n432 B.n431 10.6151
R679 B.n431 B.n14 10.6151
R680 B.n427 B.n14 10.6151
R681 B.n427 B.n426 10.6151
R682 B.n426 B.n425 10.6151
R683 B.n425 B.n16 10.6151
R684 B.n421 B.n16 10.6151
R685 B.n421 B.n420 10.6151
R686 B.n420 B.n419 10.6151
R687 B.n419 B.n18 10.6151
R688 B.n415 B.n18 10.6151
R689 B.n415 B.n414 10.6151
R690 B.n414 B.n413 10.6151
R691 B.n413 B.n20 10.6151
R692 B.n409 B.n20 10.6151
R693 B.n409 B.n408 10.6151
R694 B.n408 B.n407 10.6151
R695 B.n407 B.n22 10.6151
R696 B.n403 B.n22 10.6151
R697 B.n403 B.n402 10.6151
R698 B.n402 B.n401 10.6151
R699 B.n386 B.n30 6.5566
R700 B.n374 B.n373 6.5566
R701 B.n202 B.n98 6.5566
R702 B.n215 B.n214 6.5566
R703 B.n389 B.n30 4.05904
R704 B.n373 B.n372 4.05904
R705 B.n199 B.n98 4.05904
R706 B.n216 B.n215 4.05904
R707 B.n467 B.n0 2.81026
R708 B.n467 B.n1 2.81026
R709 VP.n21 VP.n20 161.3
R710 VP.n19 VP.n1 161.3
R711 VP.n18 VP.n17 161.3
R712 VP.n16 VP.n2 161.3
R713 VP.n15 VP.n14 161.3
R714 VP.n13 VP.n3 161.3
R715 VP.n12 VP.n11 161.3
R716 VP.n10 VP.n4 161.3
R717 VP.n9 VP.n8 161.3
R718 VP.n7 VP.n6 88.8441
R719 VP.n22 VP.n0 88.8441
R720 VP.n6 VP.n5 42.9554
R721 VP.n14 VP.n13 40.4934
R722 VP.n14 VP.n2 40.4934
R723 VP.n5 VP.t3 36.7201
R724 VP.n5 VP.t1 35.3897
R725 VP.n8 VP.n4 24.4675
R726 VP.n12 VP.n4 24.4675
R727 VP.n13 VP.n12 24.4675
R728 VP.n18 VP.n2 24.4675
R729 VP.n19 VP.n18 24.4675
R730 VP.n20 VP.n19 24.4675
R731 VP.n7 VP.t0 3.30453
R732 VP.n0 VP.t2 3.30453
R733 VP.n8 VP.n7 1.22385
R734 VP.n20 VP.n0 1.22385
R735 VP.n9 VP.n6 0.354971
R736 VP.n22 VP.n21 0.354971
R737 VP VP.n22 0.26696
R738 VP.n10 VP.n9 0.189894
R739 VP.n11 VP.n10 0.189894
R740 VP.n11 VP.n3 0.189894
R741 VP.n15 VP.n3 0.189894
R742 VP.n16 VP.n15 0.189894
R743 VP.n17 VP.n16 0.189894
R744 VP.n17 VP.n1 0.189894
R745 VP.n21 VP.n1 0.189894
R746 VDD1 VDD1.n1 667.273
R747 VDD1 VDD1.n0 632.177
R748 VDD1.n0 VDD1.t0 63.7358
R749 VDD1.n0 VDD1.t2 63.7358
R750 VDD1.n1 VDD1.t3 63.7358
R751 VDD1.n1 VDD1.t1 63.7358
R752 VTAIL.n7 VTAIL.t2 679.176
R753 VTAIL.n0 VTAIL.t1 679.176
R754 VTAIL.n1 VTAIL.t5 679.176
R755 VTAIL.n2 VTAIL.t7 679.176
R756 VTAIL.n6 VTAIL.t6 679.176
R757 VTAIL.n5 VTAIL.t4 679.176
R758 VTAIL.n4 VTAIL.t3 679.176
R759 VTAIL.n3 VTAIL.t0 679.176
R760 VTAIL.n7 VTAIL.n6 16.2979
R761 VTAIL.n3 VTAIL.n2 16.2979
R762 VTAIL.n4 VTAIL.n3 3.49188
R763 VTAIL.n6 VTAIL.n5 3.49188
R764 VTAIL.n2 VTAIL.n1 3.49188
R765 VTAIL VTAIL.n0 1.80438
R766 VTAIL VTAIL.n7 1.688
R767 VTAIL.n5 VTAIL.n4 0.470328
R768 VTAIL.n1 VTAIL.n0 0.470328
R769 VN VN.n1 43.1208
R770 VN.n1 VN.t1 36.7202
R771 VN.n0 VN.t2 36.7202
R772 VN.n0 VN.t0 35.3897
R773 VN.n1 VN.t3 35.3897
R774 VN VN.n0 1.92
R775 VDD2.n2 VDD2.n0 666.747
R776 VDD2.n2 VDD2.n1 632.119
R777 VDD2.n1 VDD2.t0 63.7358
R778 VDD2.n1 VDD2.t2 63.7358
R779 VDD2.n0 VDD2.t1 63.7358
R780 VDD2.n0 VDD2.t3 63.7358
R781 VDD2 VDD2.n2 0.0586897
C0 VDD2 B 1.22477f
C1 VDD2 VN 0.550193f
C2 w_n3400_n1070# B 7.56127f
C3 VTAIL VDD2 3.37097f
C4 w_n3400_n1070# VN 5.76363f
C5 w_n3400_n1070# VTAIL 1.41285f
C6 VDD2 VDD1 1.29726f
C7 VP VDD2 0.475422f
C8 w_n3400_n1070# VDD1 1.34078f
C9 w_n3400_n1070# VP 6.19394f
C10 VN B 1.07067f
C11 VTAIL B 1.15523f
C12 VTAIL VN 1.66493f
C13 B VDD1 1.15298f
C14 VP B 1.8043f
C15 w_n3400_n1070# VDD2 1.42019f
C16 VN VDD1 0.157735f
C17 VTAIL VDD1 3.30926f
C18 VP VN 4.88344f
C19 VTAIL VP 1.67904f
C20 VP VDD1 0.864322f
C21 VDD2 VSUBS 0.868274f
C22 VDD1 VSUBS 4.18106f
C23 VTAIL VSUBS 0.526162f
C24 VN VSUBS 6.87435f
C25 VP VSUBS 2.27521f
C26 B VSUBS 4.017826f
C27 w_n3400_n1070# VSUBS 47.2056f
C28 VDD2.t1 VSUBS 0.011667f
C29 VDD2.t3 VSUBS 0.011667f
C30 VDD2.n0 VSUBS 0.073355f
C31 VDD2.t0 VSUBS 0.011667f
C32 VDD2.t2 VSUBS 0.011667f
C33 VDD2.n1 VSUBS 0.026113f
C34 VDD2.n2 VSUBS 2.92194f
C35 VN.t0 VSUBS 0.664927f
C36 VN.t2 VSUBS 0.695245f
C37 VN.n0 VSUBS 0.786086f
C38 VN.t3 VSUBS 0.664927f
C39 VN.t1 VSUBS 0.695245f
C40 VN.n1 VSUBS 3.82247f
C41 VTAIL.t1 VSUBS 0.052779f
C42 VTAIL.n0 VSUBS 0.259972f
C43 VTAIL.t5 VSUBS 0.052779f
C44 VTAIL.n1 VSUBS 0.420219f
C45 VTAIL.t7 VSUBS 0.052779f
C46 VTAIL.n2 VSUBS 1.14922f
C47 VTAIL.t0 VSUBS 0.052779f
C48 VTAIL.n3 VSUBS 1.14922f
C49 VTAIL.t3 VSUBS 0.052779f
C50 VTAIL.n4 VSUBS 0.420219f
C51 VTAIL.t4 VSUBS 0.052779f
C52 VTAIL.n5 VSUBS 0.420219f
C53 VTAIL.t6 VSUBS 0.052779f
C54 VTAIL.n6 VSUBS 1.14922f
C55 VTAIL.t2 VSUBS 0.052779f
C56 VTAIL.n7 VSUBS 0.977924f
C57 VDD1.t0 VSUBS 0.010979f
C58 VDD1.t2 VSUBS 0.010979f
C59 VDD1.n0 VSUBS 0.024608f
C60 VDD1.t3 VSUBS 0.010979f
C61 VDD1.t1 VSUBS 0.010979f
C62 VDD1.n1 VSUBS 0.072549f
C63 VP.t2 VSUBS 0.114333f
C64 VP.n0 VSUBS 0.390201f
C65 VP.n1 VSUBS 0.062077f
C66 VP.n2 VSUBS 0.123378f
C67 VP.n3 VSUBS 0.062077f
C68 VP.n4 VSUBS 0.115696f
C69 VP.t3 VSUBS 0.726903f
C70 VP.t1 VSUBS 0.695207f
C71 VP.n5 VSUBS 3.96983f
C72 VP.n6 VSUBS 2.87103f
C73 VP.t0 VSUBS 0.114333f
C74 VP.n7 VSUBS 0.390201f
C75 VP.n8 VSUBS 0.06143f
C76 VP.n9 VSUBS 0.100191f
C77 VP.n10 VSUBS 0.062077f
C78 VP.n11 VSUBS 0.062077f
C79 VP.n12 VSUBS 0.115696f
C80 VP.n13 VSUBS 0.123378f
C81 VP.n14 VSUBS 0.050184f
C82 VP.n15 VSUBS 0.062077f
C83 VP.n16 VSUBS 0.062077f
C84 VP.n17 VSUBS 0.062077f
C85 VP.n18 VSUBS 0.115696f
C86 VP.n19 VSUBS 0.115696f
C87 VP.n20 VSUBS 0.06143f
C88 VP.n21 VSUBS 0.100191f
C89 VP.n22 VSUBS 0.190798f
C90 B.n0 VSUBS 0.007795f
C91 B.n1 VSUBS 0.007795f
C92 B.n2 VSUBS 0.012327f
C93 B.n3 VSUBS 0.012327f
C94 B.n4 VSUBS 0.012327f
C95 B.n5 VSUBS 0.012327f
C96 B.n6 VSUBS 0.012327f
C97 B.n7 VSUBS 0.012327f
C98 B.n8 VSUBS 0.012327f
C99 B.n9 VSUBS 0.012327f
C100 B.n10 VSUBS 0.012327f
C101 B.n11 VSUBS 0.012327f
C102 B.n12 VSUBS 0.012327f
C103 B.n13 VSUBS 0.012327f
C104 B.n14 VSUBS 0.012327f
C105 B.n15 VSUBS 0.012327f
C106 B.n16 VSUBS 0.012327f
C107 B.n17 VSUBS 0.012327f
C108 B.n18 VSUBS 0.012327f
C109 B.n19 VSUBS 0.012327f
C110 B.n20 VSUBS 0.012327f
C111 B.n21 VSUBS 0.012327f
C112 B.n22 VSUBS 0.012327f
C113 B.n23 VSUBS 0.012327f
C114 B.n24 VSUBS 0.028841f
C115 B.n25 VSUBS 0.012327f
C116 B.n26 VSUBS 0.012327f
C117 B.n27 VSUBS 0.012327f
C118 B.t11 VSUBS 0.016699f
C119 B.t10 VSUBS 0.022739f
C120 B.t9 VSUBS 0.167986f
C121 B.n28 VSUBS 0.119882f
C122 B.n29 VSUBS 0.075007f
C123 B.n30 VSUBS 0.028559f
C124 B.n31 VSUBS 0.012327f
C125 B.n32 VSUBS 0.012327f
C126 B.n33 VSUBS 0.012327f
C127 B.n34 VSUBS 0.012327f
C128 B.n35 VSUBS 0.012327f
C129 B.t5 VSUBS 0.016699f
C130 B.t4 VSUBS 0.022739f
C131 B.t3 VSUBS 0.167986f
C132 B.n36 VSUBS 0.119882f
C133 B.n37 VSUBS 0.075007f
C134 B.n38 VSUBS 0.012327f
C135 B.n39 VSUBS 0.012327f
C136 B.n40 VSUBS 0.012327f
C137 B.n41 VSUBS 0.028079f
C138 B.n42 VSUBS 0.012327f
C139 B.n43 VSUBS 0.012327f
C140 B.n44 VSUBS 0.012327f
C141 B.n45 VSUBS 0.012327f
C142 B.n46 VSUBS 0.012327f
C143 B.n47 VSUBS 0.012327f
C144 B.n48 VSUBS 0.012327f
C145 B.n49 VSUBS 0.012327f
C146 B.n50 VSUBS 0.012327f
C147 B.n51 VSUBS 0.012327f
C148 B.n52 VSUBS 0.012327f
C149 B.n53 VSUBS 0.012327f
C150 B.n54 VSUBS 0.012327f
C151 B.n55 VSUBS 0.012327f
C152 B.n56 VSUBS 0.012327f
C153 B.n57 VSUBS 0.012327f
C154 B.n58 VSUBS 0.012327f
C155 B.n59 VSUBS 0.012327f
C156 B.n60 VSUBS 0.012327f
C157 B.n61 VSUBS 0.012327f
C158 B.n62 VSUBS 0.012327f
C159 B.n63 VSUBS 0.012327f
C160 B.n64 VSUBS 0.012327f
C161 B.n65 VSUBS 0.012327f
C162 B.n66 VSUBS 0.012327f
C163 B.n67 VSUBS 0.012327f
C164 B.n68 VSUBS 0.012327f
C165 B.n69 VSUBS 0.012327f
C166 B.n70 VSUBS 0.012327f
C167 B.n71 VSUBS 0.012327f
C168 B.n72 VSUBS 0.012327f
C169 B.n73 VSUBS 0.012327f
C170 B.n74 VSUBS 0.012327f
C171 B.n75 VSUBS 0.012327f
C172 B.n76 VSUBS 0.012327f
C173 B.n77 VSUBS 0.012327f
C174 B.n78 VSUBS 0.012327f
C175 B.n79 VSUBS 0.012327f
C176 B.n80 VSUBS 0.012327f
C177 B.n81 VSUBS 0.012327f
C178 B.n82 VSUBS 0.012327f
C179 B.n83 VSUBS 0.012327f
C180 B.n84 VSUBS 0.012327f
C181 B.n85 VSUBS 0.028079f
C182 B.n86 VSUBS 0.012327f
C183 B.n87 VSUBS 0.012327f
C184 B.n88 VSUBS 0.012327f
C185 B.n89 VSUBS 0.012327f
C186 B.t7 VSUBS 0.016699f
C187 B.t8 VSUBS 0.022739f
C188 B.t6 VSUBS 0.167986f
C189 B.n90 VSUBS 0.119882f
C190 B.n91 VSUBS 0.075007f
C191 B.n92 VSUBS 0.012327f
C192 B.n93 VSUBS 0.012327f
C193 B.n94 VSUBS 0.012327f
C194 B.n95 VSUBS 0.012327f
C195 B.t1 VSUBS 0.016699f
C196 B.t2 VSUBS 0.022739f
C197 B.t0 VSUBS 0.167986f
C198 B.n96 VSUBS 0.119882f
C199 B.n97 VSUBS 0.075007f
C200 B.n98 VSUBS 0.028559f
C201 B.n99 VSUBS 0.012327f
C202 B.n100 VSUBS 0.012327f
C203 B.n101 VSUBS 0.012327f
C204 B.n102 VSUBS 0.028841f
C205 B.n103 VSUBS 0.012327f
C206 B.n104 VSUBS 0.012327f
C207 B.n105 VSUBS 0.012327f
C208 B.n106 VSUBS 0.012327f
C209 B.n107 VSUBS 0.012327f
C210 B.n108 VSUBS 0.012327f
C211 B.n109 VSUBS 0.012327f
C212 B.n110 VSUBS 0.012327f
C213 B.n111 VSUBS 0.012327f
C214 B.n112 VSUBS 0.012327f
C215 B.n113 VSUBS 0.012327f
C216 B.n114 VSUBS 0.012327f
C217 B.n115 VSUBS 0.012327f
C218 B.n116 VSUBS 0.012327f
C219 B.n117 VSUBS 0.012327f
C220 B.n118 VSUBS 0.012327f
C221 B.n119 VSUBS 0.012327f
C222 B.n120 VSUBS 0.012327f
C223 B.n121 VSUBS 0.012327f
C224 B.n122 VSUBS 0.012327f
C225 B.n123 VSUBS 0.012327f
C226 B.n124 VSUBS 0.012327f
C227 B.n125 VSUBS 0.012327f
C228 B.n126 VSUBS 0.012327f
C229 B.n127 VSUBS 0.012327f
C230 B.n128 VSUBS 0.012327f
C231 B.n129 VSUBS 0.012327f
C232 B.n130 VSUBS 0.012327f
C233 B.n131 VSUBS 0.012327f
C234 B.n132 VSUBS 0.012327f
C235 B.n133 VSUBS 0.012327f
C236 B.n134 VSUBS 0.012327f
C237 B.n135 VSUBS 0.012327f
C238 B.n136 VSUBS 0.012327f
C239 B.n137 VSUBS 0.012327f
C240 B.n138 VSUBS 0.012327f
C241 B.n139 VSUBS 0.012327f
C242 B.n140 VSUBS 0.012327f
C243 B.n141 VSUBS 0.012327f
C244 B.n142 VSUBS 0.012327f
C245 B.n143 VSUBS 0.012327f
C246 B.n144 VSUBS 0.012327f
C247 B.n145 VSUBS 0.012327f
C248 B.n146 VSUBS 0.012327f
C249 B.n147 VSUBS 0.012327f
C250 B.n148 VSUBS 0.012327f
C251 B.n149 VSUBS 0.012327f
C252 B.n150 VSUBS 0.012327f
C253 B.n151 VSUBS 0.012327f
C254 B.n152 VSUBS 0.012327f
C255 B.n153 VSUBS 0.012327f
C256 B.n154 VSUBS 0.012327f
C257 B.n155 VSUBS 0.012327f
C258 B.n156 VSUBS 0.012327f
C259 B.n157 VSUBS 0.012327f
C260 B.n158 VSUBS 0.012327f
C261 B.n159 VSUBS 0.012327f
C262 B.n160 VSUBS 0.012327f
C263 B.n161 VSUBS 0.012327f
C264 B.n162 VSUBS 0.012327f
C265 B.n163 VSUBS 0.012327f
C266 B.n164 VSUBS 0.012327f
C267 B.n165 VSUBS 0.012327f
C268 B.n166 VSUBS 0.012327f
C269 B.n167 VSUBS 0.012327f
C270 B.n168 VSUBS 0.012327f
C271 B.n169 VSUBS 0.012327f
C272 B.n170 VSUBS 0.012327f
C273 B.n171 VSUBS 0.012327f
C274 B.n172 VSUBS 0.012327f
C275 B.n173 VSUBS 0.012327f
C276 B.n174 VSUBS 0.012327f
C277 B.n175 VSUBS 0.012327f
C278 B.n176 VSUBS 0.012327f
C279 B.n177 VSUBS 0.012327f
C280 B.n178 VSUBS 0.012327f
C281 B.n179 VSUBS 0.012327f
C282 B.n180 VSUBS 0.012327f
C283 B.n181 VSUBS 0.012327f
C284 B.n182 VSUBS 0.012327f
C285 B.n183 VSUBS 0.012327f
C286 B.n184 VSUBS 0.012327f
C287 B.n185 VSUBS 0.012327f
C288 B.n186 VSUBS 0.012327f
C289 B.n187 VSUBS 0.028079f
C290 B.n188 VSUBS 0.028079f
C291 B.n189 VSUBS 0.028841f
C292 B.n190 VSUBS 0.012327f
C293 B.n191 VSUBS 0.012327f
C294 B.n192 VSUBS 0.012327f
C295 B.n193 VSUBS 0.012327f
C296 B.n194 VSUBS 0.012327f
C297 B.n195 VSUBS 0.012327f
C298 B.n196 VSUBS 0.012327f
C299 B.n197 VSUBS 0.012327f
C300 B.n198 VSUBS 0.012327f
C301 B.n199 VSUBS 0.00852f
C302 B.n200 VSUBS 0.012327f
C303 B.n201 VSUBS 0.012327f
C304 B.n202 VSUBS 0.00997f
C305 B.n203 VSUBS 0.012327f
C306 B.n204 VSUBS 0.012327f
C307 B.n205 VSUBS 0.012327f
C308 B.n206 VSUBS 0.012327f
C309 B.n207 VSUBS 0.012327f
C310 B.n208 VSUBS 0.012327f
C311 B.n209 VSUBS 0.012327f
C312 B.n210 VSUBS 0.012327f
C313 B.n211 VSUBS 0.012327f
C314 B.n212 VSUBS 0.012327f
C315 B.n213 VSUBS 0.012327f
C316 B.n214 VSUBS 0.00997f
C317 B.n215 VSUBS 0.028559f
C318 B.n216 VSUBS 0.00852f
C319 B.n217 VSUBS 0.012327f
C320 B.n218 VSUBS 0.012327f
C321 B.n219 VSUBS 0.012327f
C322 B.n220 VSUBS 0.012327f
C323 B.n221 VSUBS 0.012327f
C324 B.n222 VSUBS 0.012327f
C325 B.n223 VSUBS 0.012327f
C326 B.n224 VSUBS 0.012327f
C327 B.n225 VSUBS 0.012327f
C328 B.n226 VSUBS 0.028841f
C329 B.n227 VSUBS 0.028841f
C330 B.n228 VSUBS 0.028079f
C331 B.n229 VSUBS 0.012327f
C332 B.n230 VSUBS 0.012327f
C333 B.n231 VSUBS 0.012327f
C334 B.n232 VSUBS 0.012327f
C335 B.n233 VSUBS 0.012327f
C336 B.n234 VSUBS 0.012327f
C337 B.n235 VSUBS 0.012327f
C338 B.n236 VSUBS 0.012327f
C339 B.n237 VSUBS 0.012327f
C340 B.n238 VSUBS 0.012327f
C341 B.n239 VSUBS 0.012327f
C342 B.n240 VSUBS 0.012327f
C343 B.n241 VSUBS 0.012327f
C344 B.n242 VSUBS 0.012327f
C345 B.n243 VSUBS 0.012327f
C346 B.n244 VSUBS 0.012327f
C347 B.n245 VSUBS 0.012327f
C348 B.n246 VSUBS 0.012327f
C349 B.n247 VSUBS 0.012327f
C350 B.n248 VSUBS 0.012327f
C351 B.n249 VSUBS 0.012327f
C352 B.n250 VSUBS 0.012327f
C353 B.n251 VSUBS 0.012327f
C354 B.n252 VSUBS 0.012327f
C355 B.n253 VSUBS 0.012327f
C356 B.n254 VSUBS 0.012327f
C357 B.n255 VSUBS 0.012327f
C358 B.n256 VSUBS 0.012327f
C359 B.n257 VSUBS 0.012327f
C360 B.n258 VSUBS 0.012327f
C361 B.n259 VSUBS 0.012327f
C362 B.n260 VSUBS 0.012327f
C363 B.n261 VSUBS 0.012327f
C364 B.n262 VSUBS 0.012327f
C365 B.n263 VSUBS 0.012327f
C366 B.n264 VSUBS 0.012327f
C367 B.n265 VSUBS 0.012327f
C368 B.n266 VSUBS 0.012327f
C369 B.n267 VSUBS 0.012327f
C370 B.n268 VSUBS 0.012327f
C371 B.n269 VSUBS 0.012327f
C372 B.n270 VSUBS 0.012327f
C373 B.n271 VSUBS 0.012327f
C374 B.n272 VSUBS 0.012327f
C375 B.n273 VSUBS 0.012327f
C376 B.n274 VSUBS 0.012327f
C377 B.n275 VSUBS 0.012327f
C378 B.n276 VSUBS 0.012327f
C379 B.n277 VSUBS 0.012327f
C380 B.n278 VSUBS 0.012327f
C381 B.n279 VSUBS 0.012327f
C382 B.n280 VSUBS 0.012327f
C383 B.n281 VSUBS 0.012327f
C384 B.n282 VSUBS 0.012327f
C385 B.n283 VSUBS 0.012327f
C386 B.n284 VSUBS 0.012327f
C387 B.n285 VSUBS 0.012327f
C388 B.n286 VSUBS 0.012327f
C389 B.n287 VSUBS 0.012327f
C390 B.n288 VSUBS 0.012327f
C391 B.n289 VSUBS 0.012327f
C392 B.n290 VSUBS 0.012327f
C393 B.n291 VSUBS 0.012327f
C394 B.n292 VSUBS 0.012327f
C395 B.n293 VSUBS 0.012327f
C396 B.n294 VSUBS 0.012327f
C397 B.n295 VSUBS 0.012327f
C398 B.n296 VSUBS 0.012327f
C399 B.n297 VSUBS 0.012327f
C400 B.n298 VSUBS 0.012327f
C401 B.n299 VSUBS 0.012327f
C402 B.n300 VSUBS 0.012327f
C403 B.n301 VSUBS 0.012327f
C404 B.n302 VSUBS 0.012327f
C405 B.n303 VSUBS 0.012327f
C406 B.n304 VSUBS 0.012327f
C407 B.n305 VSUBS 0.012327f
C408 B.n306 VSUBS 0.012327f
C409 B.n307 VSUBS 0.012327f
C410 B.n308 VSUBS 0.012327f
C411 B.n309 VSUBS 0.012327f
C412 B.n310 VSUBS 0.012327f
C413 B.n311 VSUBS 0.012327f
C414 B.n312 VSUBS 0.012327f
C415 B.n313 VSUBS 0.012327f
C416 B.n314 VSUBS 0.012327f
C417 B.n315 VSUBS 0.012327f
C418 B.n316 VSUBS 0.012327f
C419 B.n317 VSUBS 0.012327f
C420 B.n318 VSUBS 0.012327f
C421 B.n319 VSUBS 0.012327f
C422 B.n320 VSUBS 0.012327f
C423 B.n321 VSUBS 0.012327f
C424 B.n322 VSUBS 0.012327f
C425 B.n323 VSUBS 0.012327f
C426 B.n324 VSUBS 0.012327f
C427 B.n325 VSUBS 0.012327f
C428 B.n326 VSUBS 0.012327f
C429 B.n327 VSUBS 0.012327f
C430 B.n328 VSUBS 0.012327f
C431 B.n329 VSUBS 0.012327f
C432 B.n330 VSUBS 0.012327f
C433 B.n331 VSUBS 0.012327f
C434 B.n332 VSUBS 0.012327f
C435 B.n333 VSUBS 0.012327f
C436 B.n334 VSUBS 0.012327f
C437 B.n335 VSUBS 0.012327f
C438 B.n336 VSUBS 0.012327f
C439 B.n337 VSUBS 0.012327f
C440 B.n338 VSUBS 0.012327f
C441 B.n339 VSUBS 0.012327f
C442 B.n340 VSUBS 0.012327f
C443 B.n341 VSUBS 0.012327f
C444 B.n342 VSUBS 0.012327f
C445 B.n343 VSUBS 0.012327f
C446 B.n344 VSUBS 0.012327f
C447 B.n345 VSUBS 0.012327f
C448 B.n346 VSUBS 0.012327f
C449 B.n347 VSUBS 0.012327f
C450 B.n348 VSUBS 0.012327f
C451 B.n349 VSUBS 0.012327f
C452 B.n350 VSUBS 0.012327f
C453 B.n351 VSUBS 0.012327f
C454 B.n352 VSUBS 0.012327f
C455 B.n353 VSUBS 0.012327f
C456 B.n354 VSUBS 0.012327f
C457 B.n355 VSUBS 0.012327f
C458 B.n356 VSUBS 0.012327f
C459 B.n357 VSUBS 0.012327f
C460 B.n358 VSUBS 0.012327f
C461 B.n359 VSUBS 0.012327f
C462 B.n360 VSUBS 0.029566f
C463 B.n361 VSUBS 0.027354f
C464 B.n362 VSUBS 0.028841f
C465 B.n363 VSUBS 0.012327f
C466 B.n364 VSUBS 0.012327f
C467 B.n365 VSUBS 0.012327f
C468 B.n366 VSUBS 0.012327f
C469 B.n367 VSUBS 0.012327f
C470 B.n368 VSUBS 0.012327f
C471 B.n369 VSUBS 0.012327f
C472 B.n370 VSUBS 0.012327f
C473 B.n371 VSUBS 0.012327f
C474 B.n372 VSUBS 0.00852f
C475 B.n373 VSUBS 0.028559f
C476 B.n374 VSUBS 0.00997f
C477 B.n375 VSUBS 0.012327f
C478 B.n376 VSUBS 0.012327f
C479 B.n377 VSUBS 0.012327f
C480 B.n378 VSUBS 0.012327f
C481 B.n379 VSUBS 0.012327f
C482 B.n380 VSUBS 0.012327f
C483 B.n381 VSUBS 0.012327f
C484 B.n382 VSUBS 0.012327f
C485 B.n383 VSUBS 0.012327f
C486 B.n384 VSUBS 0.012327f
C487 B.n385 VSUBS 0.012327f
C488 B.n386 VSUBS 0.00997f
C489 B.n387 VSUBS 0.012327f
C490 B.n388 VSUBS 0.012327f
C491 B.n389 VSUBS 0.00852f
C492 B.n390 VSUBS 0.012327f
C493 B.n391 VSUBS 0.012327f
C494 B.n392 VSUBS 0.012327f
C495 B.n393 VSUBS 0.012327f
C496 B.n394 VSUBS 0.012327f
C497 B.n395 VSUBS 0.012327f
C498 B.n396 VSUBS 0.012327f
C499 B.n397 VSUBS 0.012327f
C500 B.n398 VSUBS 0.012327f
C501 B.n399 VSUBS 0.028841f
C502 B.n400 VSUBS 0.028079f
C503 B.n401 VSUBS 0.028079f
C504 B.n402 VSUBS 0.012327f
C505 B.n403 VSUBS 0.012327f
C506 B.n404 VSUBS 0.012327f
C507 B.n405 VSUBS 0.012327f
C508 B.n406 VSUBS 0.012327f
C509 B.n407 VSUBS 0.012327f
C510 B.n408 VSUBS 0.012327f
C511 B.n409 VSUBS 0.012327f
C512 B.n410 VSUBS 0.012327f
C513 B.n411 VSUBS 0.012327f
C514 B.n412 VSUBS 0.012327f
C515 B.n413 VSUBS 0.012327f
C516 B.n414 VSUBS 0.012327f
C517 B.n415 VSUBS 0.012327f
C518 B.n416 VSUBS 0.012327f
C519 B.n417 VSUBS 0.012327f
C520 B.n418 VSUBS 0.012327f
C521 B.n419 VSUBS 0.012327f
C522 B.n420 VSUBS 0.012327f
C523 B.n421 VSUBS 0.012327f
C524 B.n422 VSUBS 0.012327f
C525 B.n423 VSUBS 0.012327f
C526 B.n424 VSUBS 0.012327f
C527 B.n425 VSUBS 0.012327f
C528 B.n426 VSUBS 0.012327f
C529 B.n427 VSUBS 0.012327f
C530 B.n428 VSUBS 0.012327f
C531 B.n429 VSUBS 0.012327f
C532 B.n430 VSUBS 0.012327f
C533 B.n431 VSUBS 0.012327f
C534 B.n432 VSUBS 0.012327f
C535 B.n433 VSUBS 0.012327f
C536 B.n434 VSUBS 0.012327f
C537 B.n435 VSUBS 0.012327f
C538 B.n436 VSUBS 0.012327f
C539 B.n437 VSUBS 0.012327f
C540 B.n438 VSUBS 0.012327f
C541 B.n439 VSUBS 0.012327f
C542 B.n440 VSUBS 0.012327f
C543 B.n441 VSUBS 0.012327f
C544 B.n442 VSUBS 0.012327f
C545 B.n443 VSUBS 0.012327f
C546 B.n444 VSUBS 0.012327f
C547 B.n445 VSUBS 0.012327f
C548 B.n446 VSUBS 0.012327f
C549 B.n447 VSUBS 0.012327f
C550 B.n448 VSUBS 0.012327f
C551 B.n449 VSUBS 0.012327f
C552 B.n450 VSUBS 0.012327f
C553 B.n451 VSUBS 0.012327f
C554 B.n452 VSUBS 0.012327f
C555 B.n453 VSUBS 0.012327f
C556 B.n454 VSUBS 0.012327f
C557 B.n455 VSUBS 0.012327f
C558 B.n456 VSUBS 0.012327f
C559 B.n457 VSUBS 0.012327f
C560 B.n458 VSUBS 0.012327f
C561 B.n459 VSUBS 0.012327f
C562 B.n460 VSUBS 0.012327f
C563 B.n461 VSUBS 0.012327f
C564 B.n462 VSUBS 0.012327f
C565 B.n463 VSUBS 0.012327f
C566 B.n464 VSUBS 0.012327f
C567 B.n465 VSUBS 0.012327f
C568 B.n466 VSUBS 0.012327f
C569 B.n467 VSUBS 0.027912f
.ends

