* NGSPICE file created from diff_pair_sample_0659.ext - technology: sky130A

.subckt diff_pair_sample_0659 VTAIL VN VP B VDD2 VDD1
X0 B.t17 B.t15 B.t16 B.t12 sky130_fd_pr__nfet_01v8 ad=4.1184 pd=21.9 as=0 ps=0 w=10.56 l=3.36
X1 B.t14 B.t11 B.t13 B.t12 sky130_fd_pr__nfet_01v8 ad=4.1184 pd=21.9 as=0 ps=0 w=10.56 l=3.36
X2 VTAIL.t5 VN.t0 VDD2.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=4.1184 pd=21.9 as=1.7424 ps=10.89 w=10.56 l=3.36
X3 B.t10 B.t8 B.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=4.1184 pd=21.9 as=0 ps=0 w=10.56 l=3.36
X4 VTAIL.t7 VP.t0 VDD1.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=4.1184 pd=21.9 as=1.7424 ps=10.89 w=10.56 l=3.36
X5 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=4.1184 pd=21.9 as=0 ps=0 w=10.56 l=3.36
X6 VDD2.t2 VN.t1 VTAIL.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=1.7424 pd=10.89 as=4.1184 ps=21.9 w=10.56 l=3.36
X7 VDD2.t0 VN.t2 VTAIL.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=1.7424 pd=10.89 as=4.1184 ps=21.9 w=10.56 l=3.36
X8 VTAIL.t2 VN.t3 VDD2.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=4.1184 pd=21.9 as=1.7424 ps=10.89 w=10.56 l=3.36
X9 VDD1.t2 VP.t1 VTAIL.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=1.7424 pd=10.89 as=4.1184 ps=21.9 w=10.56 l=3.36
X10 VTAIL.t0 VP.t2 VDD1.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=4.1184 pd=21.9 as=1.7424 ps=10.89 w=10.56 l=3.36
X11 VDD1.t0 VP.t3 VTAIL.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=1.7424 pd=10.89 as=4.1184 ps=21.9 w=10.56 l=3.36
R0 B.n755 B.n754 585
R1 B.n287 B.n118 585
R2 B.n286 B.n285 585
R3 B.n284 B.n283 585
R4 B.n282 B.n281 585
R5 B.n280 B.n279 585
R6 B.n278 B.n277 585
R7 B.n276 B.n275 585
R8 B.n274 B.n273 585
R9 B.n272 B.n271 585
R10 B.n270 B.n269 585
R11 B.n268 B.n267 585
R12 B.n266 B.n265 585
R13 B.n264 B.n263 585
R14 B.n262 B.n261 585
R15 B.n260 B.n259 585
R16 B.n258 B.n257 585
R17 B.n256 B.n255 585
R18 B.n254 B.n253 585
R19 B.n252 B.n251 585
R20 B.n250 B.n249 585
R21 B.n248 B.n247 585
R22 B.n246 B.n245 585
R23 B.n244 B.n243 585
R24 B.n242 B.n241 585
R25 B.n240 B.n239 585
R26 B.n238 B.n237 585
R27 B.n236 B.n235 585
R28 B.n234 B.n233 585
R29 B.n232 B.n231 585
R30 B.n230 B.n229 585
R31 B.n228 B.n227 585
R32 B.n226 B.n225 585
R33 B.n224 B.n223 585
R34 B.n222 B.n221 585
R35 B.n220 B.n219 585
R36 B.n218 B.n217 585
R37 B.n215 B.n214 585
R38 B.n213 B.n212 585
R39 B.n211 B.n210 585
R40 B.n209 B.n208 585
R41 B.n207 B.n206 585
R42 B.n205 B.n204 585
R43 B.n203 B.n202 585
R44 B.n201 B.n200 585
R45 B.n199 B.n198 585
R46 B.n197 B.n196 585
R47 B.n194 B.n193 585
R48 B.n192 B.n191 585
R49 B.n190 B.n189 585
R50 B.n188 B.n187 585
R51 B.n186 B.n185 585
R52 B.n184 B.n183 585
R53 B.n182 B.n181 585
R54 B.n180 B.n179 585
R55 B.n178 B.n177 585
R56 B.n176 B.n175 585
R57 B.n174 B.n173 585
R58 B.n172 B.n171 585
R59 B.n170 B.n169 585
R60 B.n168 B.n167 585
R61 B.n166 B.n165 585
R62 B.n164 B.n163 585
R63 B.n162 B.n161 585
R64 B.n160 B.n159 585
R65 B.n158 B.n157 585
R66 B.n156 B.n155 585
R67 B.n154 B.n153 585
R68 B.n152 B.n151 585
R69 B.n150 B.n149 585
R70 B.n148 B.n147 585
R71 B.n146 B.n145 585
R72 B.n144 B.n143 585
R73 B.n142 B.n141 585
R74 B.n140 B.n139 585
R75 B.n138 B.n137 585
R76 B.n136 B.n135 585
R77 B.n134 B.n133 585
R78 B.n132 B.n131 585
R79 B.n130 B.n129 585
R80 B.n128 B.n127 585
R81 B.n126 B.n125 585
R82 B.n124 B.n123 585
R83 B.n75 B.n74 585
R84 B.n753 B.n76 585
R85 B.n758 B.n76 585
R86 B.n752 B.n751 585
R87 B.n751 B.n72 585
R88 B.n750 B.n71 585
R89 B.n764 B.n71 585
R90 B.n749 B.n70 585
R91 B.n765 B.n70 585
R92 B.n748 B.n69 585
R93 B.n766 B.n69 585
R94 B.n747 B.n746 585
R95 B.n746 B.n65 585
R96 B.n745 B.n64 585
R97 B.n772 B.n64 585
R98 B.n744 B.n63 585
R99 B.n773 B.n63 585
R100 B.n743 B.n62 585
R101 B.n774 B.n62 585
R102 B.n742 B.n741 585
R103 B.n741 B.n58 585
R104 B.n740 B.n57 585
R105 B.n780 B.n57 585
R106 B.n739 B.n56 585
R107 B.n781 B.n56 585
R108 B.n738 B.n55 585
R109 B.n782 B.n55 585
R110 B.n737 B.n736 585
R111 B.n736 B.n51 585
R112 B.n735 B.n50 585
R113 B.n788 B.n50 585
R114 B.n734 B.n49 585
R115 B.n789 B.n49 585
R116 B.n733 B.n48 585
R117 B.n790 B.n48 585
R118 B.n732 B.n731 585
R119 B.n731 B.n44 585
R120 B.n730 B.n43 585
R121 B.n796 B.n43 585
R122 B.n729 B.n42 585
R123 B.n797 B.n42 585
R124 B.n728 B.n41 585
R125 B.n798 B.n41 585
R126 B.n727 B.n726 585
R127 B.n726 B.n37 585
R128 B.n725 B.n36 585
R129 B.n804 B.n36 585
R130 B.n724 B.n35 585
R131 B.n805 B.n35 585
R132 B.n723 B.n34 585
R133 B.n806 B.n34 585
R134 B.n722 B.n721 585
R135 B.n721 B.n30 585
R136 B.n720 B.n29 585
R137 B.n812 B.n29 585
R138 B.n719 B.n28 585
R139 B.n813 B.n28 585
R140 B.n718 B.n27 585
R141 B.n814 B.n27 585
R142 B.n717 B.n716 585
R143 B.n716 B.n23 585
R144 B.n715 B.n22 585
R145 B.n820 B.n22 585
R146 B.n714 B.n21 585
R147 B.n821 B.n21 585
R148 B.n713 B.n20 585
R149 B.n822 B.n20 585
R150 B.n712 B.n711 585
R151 B.n711 B.n19 585
R152 B.n710 B.n15 585
R153 B.n828 B.n15 585
R154 B.n709 B.n14 585
R155 B.n829 B.n14 585
R156 B.n708 B.n13 585
R157 B.n830 B.n13 585
R158 B.n707 B.n706 585
R159 B.n706 B.n12 585
R160 B.n705 B.n704 585
R161 B.n705 B.n8 585
R162 B.n703 B.n7 585
R163 B.n837 B.n7 585
R164 B.n702 B.n6 585
R165 B.n838 B.n6 585
R166 B.n701 B.n5 585
R167 B.n839 B.n5 585
R168 B.n700 B.n699 585
R169 B.n699 B.n4 585
R170 B.n698 B.n288 585
R171 B.n698 B.n697 585
R172 B.n688 B.n289 585
R173 B.n290 B.n289 585
R174 B.n690 B.n689 585
R175 B.n691 B.n690 585
R176 B.n687 B.n295 585
R177 B.n295 B.n294 585
R178 B.n686 B.n685 585
R179 B.n685 B.n684 585
R180 B.n297 B.n296 585
R181 B.n677 B.n297 585
R182 B.n676 B.n675 585
R183 B.n678 B.n676 585
R184 B.n674 B.n302 585
R185 B.n302 B.n301 585
R186 B.n673 B.n672 585
R187 B.n672 B.n671 585
R188 B.n304 B.n303 585
R189 B.n305 B.n304 585
R190 B.n664 B.n663 585
R191 B.n665 B.n664 585
R192 B.n662 B.n310 585
R193 B.n310 B.n309 585
R194 B.n661 B.n660 585
R195 B.n660 B.n659 585
R196 B.n312 B.n311 585
R197 B.n313 B.n312 585
R198 B.n652 B.n651 585
R199 B.n653 B.n652 585
R200 B.n650 B.n318 585
R201 B.n318 B.n317 585
R202 B.n649 B.n648 585
R203 B.n648 B.n647 585
R204 B.n320 B.n319 585
R205 B.n321 B.n320 585
R206 B.n640 B.n639 585
R207 B.n641 B.n640 585
R208 B.n638 B.n326 585
R209 B.n326 B.n325 585
R210 B.n637 B.n636 585
R211 B.n636 B.n635 585
R212 B.n328 B.n327 585
R213 B.n329 B.n328 585
R214 B.n628 B.n627 585
R215 B.n629 B.n628 585
R216 B.n626 B.n334 585
R217 B.n334 B.n333 585
R218 B.n625 B.n624 585
R219 B.n624 B.n623 585
R220 B.n336 B.n335 585
R221 B.n337 B.n336 585
R222 B.n616 B.n615 585
R223 B.n617 B.n616 585
R224 B.n614 B.n342 585
R225 B.n342 B.n341 585
R226 B.n613 B.n612 585
R227 B.n612 B.n611 585
R228 B.n344 B.n343 585
R229 B.n345 B.n344 585
R230 B.n604 B.n603 585
R231 B.n605 B.n604 585
R232 B.n602 B.n350 585
R233 B.n350 B.n349 585
R234 B.n601 B.n600 585
R235 B.n600 B.n599 585
R236 B.n352 B.n351 585
R237 B.n353 B.n352 585
R238 B.n592 B.n591 585
R239 B.n593 B.n592 585
R240 B.n590 B.n358 585
R241 B.n358 B.n357 585
R242 B.n589 B.n588 585
R243 B.n588 B.n587 585
R244 B.n360 B.n359 585
R245 B.n361 B.n360 585
R246 B.n580 B.n579 585
R247 B.n581 B.n580 585
R248 B.n364 B.n363 585
R249 B.n415 B.n414 585
R250 B.n416 B.n412 585
R251 B.n412 B.n365 585
R252 B.n418 B.n417 585
R253 B.n420 B.n411 585
R254 B.n423 B.n422 585
R255 B.n424 B.n410 585
R256 B.n426 B.n425 585
R257 B.n428 B.n409 585
R258 B.n431 B.n430 585
R259 B.n432 B.n408 585
R260 B.n434 B.n433 585
R261 B.n436 B.n407 585
R262 B.n439 B.n438 585
R263 B.n440 B.n406 585
R264 B.n442 B.n441 585
R265 B.n444 B.n405 585
R266 B.n447 B.n446 585
R267 B.n448 B.n404 585
R268 B.n450 B.n449 585
R269 B.n452 B.n403 585
R270 B.n455 B.n454 585
R271 B.n456 B.n402 585
R272 B.n458 B.n457 585
R273 B.n460 B.n401 585
R274 B.n463 B.n462 585
R275 B.n464 B.n400 585
R276 B.n466 B.n465 585
R277 B.n468 B.n399 585
R278 B.n471 B.n470 585
R279 B.n472 B.n398 585
R280 B.n474 B.n473 585
R281 B.n476 B.n397 585
R282 B.n479 B.n478 585
R283 B.n480 B.n396 585
R284 B.n482 B.n481 585
R285 B.n484 B.n395 585
R286 B.n487 B.n486 585
R287 B.n488 B.n391 585
R288 B.n490 B.n489 585
R289 B.n492 B.n390 585
R290 B.n495 B.n494 585
R291 B.n496 B.n389 585
R292 B.n498 B.n497 585
R293 B.n500 B.n388 585
R294 B.n503 B.n502 585
R295 B.n504 B.n385 585
R296 B.n507 B.n506 585
R297 B.n509 B.n384 585
R298 B.n512 B.n511 585
R299 B.n513 B.n383 585
R300 B.n515 B.n514 585
R301 B.n517 B.n382 585
R302 B.n520 B.n519 585
R303 B.n521 B.n381 585
R304 B.n523 B.n522 585
R305 B.n525 B.n380 585
R306 B.n528 B.n527 585
R307 B.n529 B.n379 585
R308 B.n531 B.n530 585
R309 B.n533 B.n378 585
R310 B.n536 B.n535 585
R311 B.n537 B.n377 585
R312 B.n539 B.n538 585
R313 B.n541 B.n376 585
R314 B.n544 B.n543 585
R315 B.n545 B.n375 585
R316 B.n547 B.n546 585
R317 B.n549 B.n374 585
R318 B.n552 B.n551 585
R319 B.n553 B.n373 585
R320 B.n555 B.n554 585
R321 B.n557 B.n372 585
R322 B.n560 B.n559 585
R323 B.n561 B.n371 585
R324 B.n563 B.n562 585
R325 B.n565 B.n370 585
R326 B.n568 B.n567 585
R327 B.n569 B.n369 585
R328 B.n571 B.n570 585
R329 B.n573 B.n368 585
R330 B.n574 B.n367 585
R331 B.n577 B.n576 585
R332 B.n578 B.n366 585
R333 B.n366 B.n365 585
R334 B.n583 B.n582 585
R335 B.n582 B.n581 585
R336 B.n584 B.n362 585
R337 B.n362 B.n361 585
R338 B.n586 B.n585 585
R339 B.n587 B.n586 585
R340 B.n356 B.n355 585
R341 B.n357 B.n356 585
R342 B.n595 B.n594 585
R343 B.n594 B.n593 585
R344 B.n596 B.n354 585
R345 B.n354 B.n353 585
R346 B.n598 B.n597 585
R347 B.n599 B.n598 585
R348 B.n348 B.n347 585
R349 B.n349 B.n348 585
R350 B.n607 B.n606 585
R351 B.n606 B.n605 585
R352 B.n608 B.n346 585
R353 B.n346 B.n345 585
R354 B.n610 B.n609 585
R355 B.n611 B.n610 585
R356 B.n340 B.n339 585
R357 B.n341 B.n340 585
R358 B.n619 B.n618 585
R359 B.n618 B.n617 585
R360 B.n620 B.n338 585
R361 B.n338 B.n337 585
R362 B.n622 B.n621 585
R363 B.n623 B.n622 585
R364 B.n332 B.n331 585
R365 B.n333 B.n332 585
R366 B.n631 B.n630 585
R367 B.n630 B.n629 585
R368 B.n632 B.n330 585
R369 B.n330 B.n329 585
R370 B.n634 B.n633 585
R371 B.n635 B.n634 585
R372 B.n324 B.n323 585
R373 B.n325 B.n324 585
R374 B.n643 B.n642 585
R375 B.n642 B.n641 585
R376 B.n644 B.n322 585
R377 B.n322 B.n321 585
R378 B.n646 B.n645 585
R379 B.n647 B.n646 585
R380 B.n316 B.n315 585
R381 B.n317 B.n316 585
R382 B.n655 B.n654 585
R383 B.n654 B.n653 585
R384 B.n656 B.n314 585
R385 B.n314 B.n313 585
R386 B.n658 B.n657 585
R387 B.n659 B.n658 585
R388 B.n308 B.n307 585
R389 B.n309 B.n308 585
R390 B.n667 B.n666 585
R391 B.n666 B.n665 585
R392 B.n668 B.n306 585
R393 B.n306 B.n305 585
R394 B.n670 B.n669 585
R395 B.n671 B.n670 585
R396 B.n300 B.n299 585
R397 B.n301 B.n300 585
R398 B.n680 B.n679 585
R399 B.n679 B.n678 585
R400 B.n681 B.n298 585
R401 B.n677 B.n298 585
R402 B.n683 B.n682 585
R403 B.n684 B.n683 585
R404 B.n293 B.n292 585
R405 B.n294 B.n293 585
R406 B.n693 B.n692 585
R407 B.n692 B.n691 585
R408 B.n694 B.n291 585
R409 B.n291 B.n290 585
R410 B.n696 B.n695 585
R411 B.n697 B.n696 585
R412 B.n3 B.n0 585
R413 B.n4 B.n3 585
R414 B.n836 B.n1 585
R415 B.n837 B.n836 585
R416 B.n835 B.n834 585
R417 B.n835 B.n8 585
R418 B.n833 B.n9 585
R419 B.n12 B.n9 585
R420 B.n832 B.n831 585
R421 B.n831 B.n830 585
R422 B.n11 B.n10 585
R423 B.n829 B.n11 585
R424 B.n827 B.n826 585
R425 B.n828 B.n827 585
R426 B.n825 B.n16 585
R427 B.n19 B.n16 585
R428 B.n824 B.n823 585
R429 B.n823 B.n822 585
R430 B.n18 B.n17 585
R431 B.n821 B.n18 585
R432 B.n819 B.n818 585
R433 B.n820 B.n819 585
R434 B.n817 B.n24 585
R435 B.n24 B.n23 585
R436 B.n816 B.n815 585
R437 B.n815 B.n814 585
R438 B.n26 B.n25 585
R439 B.n813 B.n26 585
R440 B.n811 B.n810 585
R441 B.n812 B.n811 585
R442 B.n809 B.n31 585
R443 B.n31 B.n30 585
R444 B.n808 B.n807 585
R445 B.n807 B.n806 585
R446 B.n33 B.n32 585
R447 B.n805 B.n33 585
R448 B.n803 B.n802 585
R449 B.n804 B.n803 585
R450 B.n801 B.n38 585
R451 B.n38 B.n37 585
R452 B.n800 B.n799 585
R453 B.n799 B.n798 585
R454 B.n40 B.n39 585
R455 B.n797 B.n40 585
R456 B.n795 B.n794 585
R457 B.n796 B.n795 585
R458 B.n793 B.n45 585
R459 B.n45 B.n44 585
R460 B.n792 B.n791 585
R461 B.n791 B.n790 585
R462 B.n47 B.n46 585
R463 B.n789 B.n47 585
R464 B.n787 B.n786 585
R465 B.n788 B.n787 585
R466 B.n785 B.n52 585
R467 B.n52 B.n51 585
R468 B.n784 B.n783 585
R469 B.n783 B.n782 585
R470 B.n54 B.n53 585
R471 B.n781 B.n54 585
R472 B.n779 B.n778 585
R473 B.n780 B.n779 585
R474 B.n777 B.n59 585
R475 B.n59 B.n58 585
R476 B.n776 B.n775 585
R477 B.n775 B.n774 585
R478 B.n61 B.n60 585
R479 B.n773 B.n61 585
R480 B.n771 B.n770 585
R481 B.n772 B.n771 585
R482 B.n769 B.n66 585
R483 B.n66 B.n65 585
R484 B.n768 B.n767 585
R485 B.n767 B.n766 585
R486 B.n68 B.n67 585
R487 B.n765 B.n68 585
R488 B.n763 B.n762 585
R489 B.n764 B.n763 585
R490 B.n761 B.n73 585
R491 B.n73 B.n72 585
R492 B.n760 B.n759 585
R493 B.n759 B.n758 585
R494 B.n840 B.n839 585
R495 B.n838 B.n2 585
R496 B.n759 B.n75 554.963
R497 B.n755 B.n76 554.963
R498 B.n580 B.n366 554.963
R499 B.n582 B.n364 554.963
R500 B.n119 B.t16 328.596
R501 B.n386 B.t10 328.596
R502 B.n121 B.t13 328.596
R503 B.n392 B.t7 328.596
R504 B.n121 B.t11 284.707
R505 B.n119 B.t15 284.707
R506 B.n386 B.t8 284.707
R507 B.n392 B.t4 284.707
R508 B.n120 B.t17 257.033
R509 B.n387 B.t9 257.033
R510 B.n122 B.t14 257.031
R511 B.n393 B.t6 257.031
R512 B.n757 B.n756 256.663
R513 B.n757 B.n117 256.663
R514 B.n757 B.n116 256.663
R515 B.n757 B.n115 256.663
R516 B.n757 B.n114 256.663
R517 B.n757 B.n113 256.663
R518 B.n757 B.n112 256.663
R519 B.n757 B.n111 256.663
R520 B.n757 B.n110 256.663
R521 B.n757 B.n109 256.663
R522 B.n757 B.n108 256.663
R523 B.n757 B.n107 256.663
R524 B.n757 B.n106 256.663
R525 B.n757 B.n105 256.663
R526 B.n757 B.n104 256.663
R527 B.n757 B.n103 256.663
R528 B.n757 B.n102 256.663
R529 B.n757 B.n101 256.663
R530 B.n757 B.n100 256.663
R531 B.n757 B.n99 256.663
R532 B.n757 B.n98 256.663
R533 B.n757 B.n97 256.663
R534 B.n757 B.n96 256.663
R535 B.n757 B.n95 256.663
R536 B.n757 B.n94 256.663
R537 B.n757 B.n93 256.663
R538 B.n757 B.n92 256.663
R539 B.n757 B.n91 256.663
R540 B.n757 B.n90 256.663
R541 B.n757 B.n89 256.663
R542 B.n757 B.n88 256.663
R543 B.n757 B.n87 256.663
R544 B.n757 B.n86 256.663
R545 B.n757 B.n85 256.663
R546 B.n757 B.n84 256.663
R547 B.n757 B.n83 256.663
R548 B.n757 B.n82 256.663
R549 B.n757 B.n81 256.663
R550 B.n757 B.n80 256.663
R551 B.n757 B.n79 256.663
R552 B.n757 B.n78 256.663
R553 B.n757 B.n77 256.663
R554 B.n413 B.n365 256.663
R555 B.n419 B.n365 256.663
R556 B.n421 B.n365 256.663
R557 B.n427 B.n365 256.663
R558 B.n429 B.n365 256.663
R559 B.n435 B.n365 256.663
R560 B.n437 B.n365 256.663
R561 B.n443 B.n365 256.663
R562 B.n445 B.n365 256.663
R563 B.n451 B.n365 256.663
R564 B.n453 B.n365 256.663
R565 B.n459 B.n365 256.663
R566 B.n461 B.n365 256.663
R567 B.n467 B.n365 256.663
R568 B.n469 B.n365 256.663
R569 B.n475 B.n365 256.663
R570 B.n477 B.n365 256.663
R571 B.n483 B.n365 256.663
R572 B.n485 B.n365 256.663
R573 B.n491 B.n365 256.663
R574 B.n493 B.n365 256.663
R575 B.n499 B.n365 256.663
R576 B.n501 B.n365 256.663
R577 B.n508 B.n365 256.663
R578 B.n510 B.n365 256.663
R579 B.n516 B.n365 256.663
R580 B.n518 B.n365 256.663
R581 B.n524 B.n365 256.663
R582 B.n526 B.n365 256.663
R583 B.n532 B.n365 256.663
R584 B.n534 B.n365 256.663
R585 B.n540 B.n365 256.663
R586 B.n542 B.n365 256.663
R587 B.n548 B.n365 256.663
R588 B.n550 B.n365 256.663
R589 B.n556 B.n365 256.663
R590 B.n558 B.n365 256.663
R591 B.n564 B.n365 256.663
R592 B.n566 B.n365 256.663
R593 B.n572 B.n365 256.663
R594 B.n575 B.n365 256.663
R595 B.n842 B.n841 256.663
R596 B.n125 B.n124 163.367
R597 B.n129 B.n128 163.367
R598 B.n133 B.n132 163.367
R599 B.n137 B.n136 163.367
R600 B.n141 B.n140 163.367
R601 B.n145 B.n144 163.367
R602 B.n149 B.n148 163.367
R603 B.n153 B.n152 163.367
R604 B.n157 B.n156 163.367
R605 B.n161 B.n160 163.367
R606 B.n165 B.n164 163.367
R607 B.n169 B.n168 163.367
R608 B.n173 B.n172 163.367
R609 B.n177 B.n176 163.367
R610 B.n181 B.n180 163.367
R611 B.n185 B.n184 163.367
R612 B.n189 B.n188 163.367
R613 B.n193 B.n192 163.367
R614 B.n198 B.n197 163.367
R615 B.n202 B.n201 163.367
R616 B.n206 B.n205 163.367
R617 B.n210 B.n209 163.367
R618 B.n214 B.n213 163.367
R619 B.n219 B.n218 163.367
R620 B.n223 B.n222 163.367
R621 B.n227 B.n226 163.367
R622 B.n231 B.n230 163.367
R623 B.n235 B.n234 163.367
R624 B.n239 B.n238 163.367
R625 B.n243 B.n242 163.367
R626 B.n247 B.n246 163.367
R627 B.n251 B.n250 163.367
R628 B.n255 B.n254 163.367
R629 B.n259 B.n258 163.367
R630 B.n263 B.n262 163.367
R631 B.n267 B.n266 163.367
R632 B.n271 B.n270 163.367
R633 B.n275 B.n274 163.367
R634 B.n279 B.n278 163.367
R635 B.n283 B.n282 163.367
R636 B.n285 B.n118 163.367
R637 B.n580 B.n360 163.367
R638 B.n588 B.n360 163.367
R639 B.n588 B.n358 163.367
R640 B.n592 B.n358 163.367
R641 B.n592 B.n352 163.367
R642 B.n600 B.n352 163.367
R643 B.n600 B.n350 163.367
R644 B.n604 B.n350 163.367
R645 B.n604 B.n344 163.367
R646 B.n612 B.n344 163.367
R647 B.n612 B.n342 163.367
R648 B.n616 B.n342 163.367
R649 B.n616 B.n336 163.367
R650 B.n624 B.n336 163.367
R651 B.n624 B.n334 163.367
R652 B.n628 B.n334 163.367
R653 B.n628 B.n328 163.367
R654 B.n636 B.n328 163.367
R655 B.n636 B.n326 163.367
R656 B.n640 B.n326 163.367
R657 B.n640 B.n320 163.367
R658 B.n648 B.n320 163.367
R659 B.n648 B.n318 163.367
R660 B.n652 B.n318 163.367
R661 B.n652 B.n312 163.367
R662 B.n660 B.n312 163.367
R663 B.n660 B.n310 163.367
R664 B.n664 B.n310 163.367
R665 B.n664 B.n304 163.367
R666 B.n672 B.n304 163.367
R667 B.n672 B.n302 163.367
R668 B.n676 B.n302 163.367
R669 B.n676 B.n297 163.367
R670 B.n685 B.n297 163.367
R671 B.n685 B.n295 163.367
R672 B.n690 B.n295 163.367
R673 B.n690 B.n289 163.367
R674 B.n698 B.n289 163.367
R675 B.n699 B.n698 163.367
R676 B.n699 B.n5 163.367
R677 B.n6 B.n5 163.367
R678 B.n7 B.n6 163.367
R679 B.n705 B.n7 163.367
R680 B.n706 B.n705 163.367
R681 B.n706 B.n13 163.367
R682 B.n14 B.n13 163.367
R683 B.n15 B.n14 163.367
R684 B.n711 B.n15 163.367
R685 B.n711 B.n20 163.367
R686 B.n21 B.n20 163.367
R687 B.n22 B.n21 163.367
R688 B.n716 B.n22 163.367
R689 B.n716 B.n27 163.367
R690 B.n28 B.n27 163.367
R691 B.n29 B.n28 163.367
R692 B.n721 B.n29 163.367
R693 B.n721 B.n34 163.367
R694 B.n35 B.n34 163.367
R695 B.n36 B.n35 163.367
R696 B.n726 B.n36 163.367
R697 B.n726 B.n41 163.367
R698 B.n42 B.n41 163.367
R699 B.n43 B.n42 163.367
R700 B.n731 B.n43 163.367
R701 B.n731 B.n48 163.367
R702 B.n49 B.n48 163.367
R703 B.n50 B.n49 163.367
R704 B.n736 B.n50 163.367
R705 B.n736 B.n55 163.367
R706 B.n56 B.n55 163.367
R707 B.n57 B.n56 163.367
R708 B.n741 B.n57 163.367
R709 B.n741 B.n62 163.367
R710 B.n63 B.n62 163.367
R711 B.n64 B.n63 163.367
R712 B.n746 B.n64 163.367
R713 B.n746 B.n69 163.367
R714 B.n70 B.n69 163.367
R715 B.n71 B.n70 163.367
R716 B.n751 B.n71 163.367
R717 B.n751 B.n76 163.367
R718 B.n414 B.n412 163.367
R719 B.n418 B.n412 163.367
R720 B.n422 B.n420 163.367
R721 B.n426 B.n410 163.367
R722 B.n430 B.n428 163.367
R723 B.n434 B.n408 163.367
R724 B.n438 B.n436 163.367
R725 B.n442 B.n406 163.367
R726 B.n446 B.n444 163.367
R727 B.n450 B.n404 163.367
R728 B.n454 B.n452 163.367
R729 B.n458 B.n402 163.367
R730 B.n462 B.n460 163.367
R731 B.n466 B.n400 163.367
R732 B.n470 B.n468 163.367
R733 B.n474 B.n398 163.367
R734 B.n478 B.n476 163.367
R735 B.n482 B.n396 163.367
R736 B.n486 B.n484 163.367
R737 B.n490 B.n391 163.367
R738 B.n494 B.n492 163.367
R739 B.n498 B.n389 163.367
R740 B.n502 B.n500 163.367
R741 B.n507 B.n385 163.367
R742 B.n511 B.n509 163.367
R743 B.n515 B.n383 163.367
R744 B.n519 B.n517 163.367
R745 B.n523 B.n381 163.367
R746 B.n527 B.n525 163.367
R747 B.n531 B.n379 163.367
R748 B.n535 B.n533 163.367
R749 B.n539 B.n377 163.367
R750 B.n543 B.n541 163.367
R751 B.n547 B.n375 163.367
R752 B.n551 B.n549 163.367
R753 B.n555 B.n373 163.367
R754 B.n559 B.n557 163.367
R755 B.n563 B.n371 163.367
R756 B.n567 B.n565 163.367
R757 B.n571 B.n369 163.367
R758 B.n574 B.n573 163.367
R759 B.n576 B.n366 163.367
R760 B.n582 B.n362 163.367
R761 B.n586 B.n362 163.367
R762 B.n586 B.n356 163.367
R763 B.n594 B.n356 163.367
R764 B.n594 B.n354 163.367
R765 B.n598 B.n354 163.367
R766 B.n598 B.n348 163.367
R767 B.n606 B.n348 163.367
R768 B.n606 B.n346 163.367
R769 B.n610 B.n346 163.367
R770 B.n610 B.n340 163.367
R771 B.n618 B.n340 163.367
R772 B.n618 B.n338 163.367
R773 B.n622 B.n338 163.367
R774 B.n622 B.n332 163.367
R775 B.n630 B.n332 163.367
R776 B.n630 B.n330 163.367
R777 B.n634 B.n330 163.367
R778 B.n634 B.n324 163.367
R779 B.n642 B.n324 163.367
R780 B.n642 B.n322 163.367
R781 B.n646 B.n322 163.367
R782 B.n646 B.n316 163.367
R783 B.n654 B.n316 163.367
R784 B.n654 B.n314 163.367
R785 B.n658 B.n314 163.367
R786 B.n658 B.n308 163.367
R787 B.n666 B.n308 163.367
R788 B.n666 B.n306 163.367
R789 B.n670 B.n306 163.367
R790 B.n670 B.n300 163.367
R791 B.n679 B.n300 163.367
R792 B.n679 B.n298 163.367
R793 B.n683 B.n298 163.367
R794 B.n683 B.n293 163.367
R795 B.n692 B.n293 163.367
R796 B.n692 B.n291 163.367
R797 B.n696 B.n291 163.367
R798 B.n696 B.n3 163.367
R799 B.n840 B.n3 163.367
R800 B.n836 B.n2 163.367
R801 B.n836 B.n835 163.367
R802 B.n835 B.n9 163.367
R803 B.n831 B.n9 163.367
R804 B.n831 B.n11 163.367
R805 B.n827 B.n11 163.367
R806 B.n827 B.n16 163.367
R807 B.n823 B.n16 163.367
R808 B.n823 B.n18 163.367
R809 B.n819 B.n18 163.367
R810 B.n819 B.n24 163.367
R811 B.n815 B.n24 163.367
R812 B.n815 B.n26 163.367
R813 B.n811 B.n26 163.367
R814 B.n811 B.n31 163.367
R815 B.n807 B.n31 163.367
R816 B.n807 B.n33 163.367
R817 B.n803 B.n33 163.367
R818 B.n803 B.n38 163.367
R819 B.n799 B.n38 163.367
R820 B.n799 B.n40 163.367
R821 B.n795 B.n40 163.367
R822 B.n795 B.n45 163.367
R823 B.n791 B.n45 163.367
R824 B.n791 B.n47 163.367
R825 B.n787 B.n47 163.367
R826 B.n787 B.n52 163.367
R827 B.n783 B.n52 163.367
R828 B.n783 B.n54 163.367
R829 B.n779 B.n54 163.367
R830 B.n779 B.n59 163.367
R831 B.n775 B.n59 163.367
R832 B.n775 B.n61 163.367
R833 B.n771 B.n61 163.367
R834 B.n771 B.n66 163.367
R835 B.n767 B.n66 163.367
R836 B.n767 B.n68 163.367
R837 B.n763 B.n68 163.367
R838 B.n763 B.n73 163.367
R839 B.n759 B.n73 163.367
R840 B.n581 B.n365 93.7801
R841 B.n758 B.n757 93.7801
R842 B.n77 B.n75 71.676
R843 B.n125 B.n78 71.676
R844 B.n129 B.n79 71.676
R845 B.n133 B.n80 71.676
R846 B.n137 B.n81 71.676
R847 B.n141 B.n82 71.676
R848 B.n145 B.n83 71.676
R849 B.n149 B.n84 71.676
R850 B.n153 B.n85 71.676
R851 B.n157 B.n86 71.676
R852 B.n161 B.n87 71.676
R853 B.n165 B.n88 71.676
R854 B.n169 B.n89 71.676
R855 B.n173 B.n90 71.676
R856 B.n177 B.n91 71.676
R857 B.n181 B.n92 71.676
R858 B.n185 B.n93 71.676
R859 B.n189 B.n94 71.676
R860 B.n193 B.n95 71.676
R861 B.n198 B.n96 71.676
R862 B.n202 B.n97 71.676
R863 B.n206 B.n98 71.676
R864 B.n210 B.n99 71.676
R865 B.n214 B.n100 71.676
R866 B.n219 B.n101 71.676
R867 B.n223 B.n102 71.676
R868 B.n227 B.n103 71.676
R869 B.n231 B.n104 71.676
R870 B.n235 B.n105 71.676
R871 B.n239 B.n106 71.676
R872 B.n243 B.n107 71.676
R873 B.n247 B.n108 71.676
R874 B.n251 B.n109 71.676
R875 B.n255 B.n110 71.676
R876 B.n259 B.n111 71.676
R877 B.n263 B.n112 71.676
R878 B.n267 B.n113 71.676
R879 B.n271 B.n114 71.676
R880 B.n275 B.n115 71.676
R881 B.n279 B.n116 71.676
R882 B.n283 B.n117 71.676
R883 B.n756 B.n118 71.676
R884 B.n756 B.n755 71.676
R885 B.n285 B.n117 71.676
R886 B.n282 B.n116 71.676
R887 B.n278 B.n115 71.676
R888 B.n274 B.n114 71.676
R889 B.n270 B.n113 71.676
R890 B.n266 B.n112 71.676
R891 B.n262 B.n111 71.676
R892 B.n258 B.n110 71.676
R893 B.n254 B.n109 71.676
R894 B.n250 B.n108 71.676
R895 B.n246 B.n107 71.676
R896 B.n242 B.n106 71.676
R897 B.n238 B.n105 71.676
R898 B.n234 B.n104 71.676
R899 B.n230 B.n103 71.676
R900 B.n226 B.n102 71.676
R901 B.n222 B.n101 71.676
R902 B.n218 B.n100 71.676
R903 B.n213 B.n99 71.676
R904 B.n209 B.n98 71.676
R905 B.n205 B.n97 71.676
R906 B.n201 B.n96 71.676
R907 B.n197 B.n95 71.676
R908 B.n192 B.n94 71.676
R909 B.n188 B.n93 71.676
R910 B.n184 B.n92 71.676
R911 B.n180 B.n91 71.676
R912 B.n176 B.n90 71.676
R913 B.n172 B.n89 71.676
R914 B.n168 B.n88 71.676
R915 B.n164 B.n87 71.676
R916 B.n160 B.n86 71.676
R917 B.n156 B.n85 71.676
R918 B.n152 B.n84 71.676
R919 B.n148 B.n83 71.676
R920 B.n144 B.n82 71.676
R921 B.n140 B.n81 71.676
R922 B.n136 B.n80 71.676
R923 B.n132 B.n79 71.676
R924 B.n128 B.n78 71.676
R925 B.n124 B.n77 71.676
R926 B.n413 B.n364 71.676
R927 B.n419 B.n418 71.676
R928 B.n422 B.n421 71.676
R929 B.n427 B.n426 71.676
R930 B.n430 B.n429 71.676
R931 B.n435 B.n434 71.676
R932 B.n438 B.n437 71.676
R933 B.n443 B.n442 71.676
R934 B.n446 B.n445 71.676
R935 B.n451 B.n450 71.676
R936 B.n454 B.n453 71.676
R937 B.n459 B.n458 71.676
R938 B.n462 B.n461 71.676
R939 B.n467 B.n466 71.676
R940 B.n470 B.n469 71.676
R941 B.n475 B.n474 71.676
R942 B.n478 B.n477 71.676
R943 B.n483 B.n482 71.676
R944 B.n486 B.n485 71.676
R945 B.n491 B.n490 71.676
R946 B.n494 B.n493 71.676
R947 B.n499 B.n498 71.676
R948 B.n502 B.n501 71.676
R949 B.n508 B.n507 71.676
R950 B.n511 B.n510 71.676
R951 B.n516 B.n515 71.676
R952 B.n519 B.n518 71.676
R953 B.n524 B.n523 71.676
R954 B.n527 B.n526 71.676
R955 B.n532 B.n531 71.676
R956 B.n535 B.n534 71.676
R957 B.n540 B.n539 71.676
R958 B.n543 B.n542 71.676
R959 B.n548 B.n547 71.676
R960 B.n551 B.n550 71.676
R961 B.n556 B.n555 71.676
R962 B.n559 B.n558 71.676
R963 B.n564 B.n563 71.676
R964 B.n567 B.n566 71.676
R965 B.n572 B.n571 71.676
R966 B.n575 B.n574 71.676
R967 B.n414 B.n413 71.676
R968 B.n420 B.n419 71.676
R969 B.n421 B.n410 71.676
R970 B.n428 B.n427 71.676
R971 B.n429 B.n408 71.676
R972 B.n436 B.n435 71.676
R973 B.n437 B.n406 71.676
R974 B.n444 B.n443 71.676
R975 B.n445 B.n404 71.676
R976 B.n452 B.n451 71.676
R977 B.n453 B.n402 71.676
R978 B.n460 B.n459 71.676
R979 B.n461 B.n400 71.676
R980 B.n468 B.n467 71.676
R981 B.n469 B.n398 71.676
R982 B.n476 B.n475 71.676
R983 B.n477 B.n396 71.676
R984 B.n484 B.n483 71.676
R985 B.n485 B.n391 71.676
R986 B.n492 B.n491 71.676
R987 B.n493 B.n389 71.676
R988 B.n500 B.n499 71.676
R989 B.n501 B.n385 71.676
R990 B.n509 B.n508 71.676
R991 B.n510 B.n383 71.676
R992 B.n517 B.n516 71.676
R993 B.n518 B.n381 71.676
R994 B.n525 B.n524 71.676
R995 B.n526 B.n379 71.676
R996 B.n533 B.n532 71.676
R997 B.n534 B.n377 71.676
R998 B.n541 B.n540 71.676
R999 B.n542 B.n375 71.676
R1000 B.n549 B.n548 71.676
R1001 B.n550 B.n373 71.676
R1002 B.n557 B.n556 71.676
R1003 B.n558 B.n371 71.676
R1004 B.n565 B.n564 71.676
R1005 B.n566 B.n369 71.676
R1006 B.n573 B.n572 71.676
R1007 B.n576 B.n575 71.676
R1008 B.n841 B.n840 71.676
R1009 B.n841 B.n2 71.676
R1010 B.n122 B.n121 71.5641
R1011 B.n120 B.n119 71.5641
R1012 B.n387 B.n386 71.5641
R1013 B.n393 B.n392 71.5641
R1014 B.n195 B.n122 59.5399
R1015 B.n216 B.n120 59.5399
R1016 B.n505 B.n387 59.5399
R1017 B.n394 B.n393 59.5399
R1018 B.n581 B.n361 47.2376
R1019 B.n587 B.n361 47.2376
R1020 B.n587 B.n357 47.2376
R1021 B.n593 B.n357 47.2376
R1022 B.n593 B.n353 47.2376
R1023 B.n599 B.n353 47.2376
R1024 B.n599 B.n349 47.2376
R1025 B.n605 B.n349 47.2376
R1026 B.n611 B.n345 47.2376
R1027 B.n611 B.n341 47.2376
R1028 B.n617 B.n341 47.2376
R1029 B.n617 B.n337 47.2376
R1030 B.n623 B.n337 47.2376
R1031 B.n623 B.n333 47.2376
R1032 B.n629 B.n333 47.2376
R1033 B.n629 B.n329 47.2376
R1034 B.n635 B.n329 47.2376
R1035 B.n635 B.n325 47.2376
R1036 B.n641 B.n325 47.2376
R1037 B.n641 B.n321 47.2376
R1038 B.n647 B.n321 47.2376
R1039 B.n653 B.n317 47.2376
R1040 B.n653 B.n313 47.2376
R1041 B.n659 B.n313 47.2376
R1042 B.n659 B.n309 47.2376
R1043 B.n665 B.n309 47.2376
R1044 B.n665 B.n305 47.2376
R1045 B.n671 B.n305 47.2376
R1046 B.n671 B.n301 47.2376
R1047 B.n678 B.n301 47.2376
R1048 B.n678 B.n677 47.2376
R1049 B.n684 B.n294 47.2376
R1050 B.n691 B.n294 47.2376
R1051 B.n691 B.n290 47.2376
R1052 B.n697 B.n290 47.2376
R1053 B.n697 B.n4 47.2376
R1054 B.n839 B.n4 47.2376
R1055 B.n839 B.n838 47.2376
R1056 B.n838 B.n837 47.2376
R1057 B.n837 B.n8 47.2376
R1058 B.n12 B.n8 47.2376
R1059 B.n830 B.n12 47.2376
R1060 B.n830 B.n829 47.2376
R1061 B.n829 B.n828 47.2376
R1062 B.n822 B.n19 47.2376
R1063 B.n822 B.n821 47.2376
R1064 B.n821 B.n820 47.2376
R1065 B.n820 B.n23 47.2376
R1066 B.n814 B.n23 47.2376
R1067 B.n814 B.n813 47.2376
R1068 B.n813 B.n812 47.2376
R1069 B.n812 B.n30 47.2376
R1070 B.n806 B.n30 47.2376
R1071 B.n806 B.n805 47.2376
R1072 B.n804 B.n37 47.2376
R1073 B.n798 B.n37 47.2376
R1074 B.n798 B.n797 47.2376
R1075 B.n797 B.n796 47.2376
R1076 B.n796 B.n44 47.2376
R1077 B.n790 B.n44 47.2376
R1078 B.n790 B.n789 47.2376
R1079 B.n789 B.n788 47.2376
R1080 B.n788 B.n51 47.2376
R1081 B.n782 B.n51 47.2376
R1082 B.n782 B.n781 47.2376
R1083 B.n781 B.n780 47.2376
R1084 B.n780 B.n58 47.2376
R1085 B.n774 B.n773 47.2376
R1086 B.n773 B.n772 47.2376
R1087 B.n772 B.n65 47.2376
R1088 B.n766 B.n65 47.2376
R1089 B.n766 B.n765 47.2376
R1090 B.n765 B.n764 47.2376
R1091 B.n764 B.n72 47.2376
R1092 B.n758 B.n72 47.2376
R1093 B.n583 B.n363 36.059
R1094 B.n579 B.n578 36.059
R1095 B.n754 B.n753 36.059
R1096 B.n760 B.n74 36.059
R1097 B.n647 B.t0 29.1764
R1098 B.t2 B.n804 29.1764
R1099 B.n605 B.t5 26.3977
R1100 B.n774 B.t12 26.3977
R1101 B.n684 B.t3 25.0084
R1102 B.n828 B.t1 25.0084
R1103 B.n677 B.t3 22.2297
R1104 B.n19 B.t1 22.2297
R1105 B.t5 B.n345 20.8404
R1106 B.t12 B.n58 20.8404
R1107 B.t0 B.n317 18.0618
R1108 B.n805 B.t2 18.0618
R1109 B B.n842 18.0485
R1110 B.n584 B.n583 10.6151
R1111 B.n585 B.n584 10.6151
R1112 B.n585 B.n355 10.6151
R1113 B.n595 B.n355 10.6151
R1114 B.n596 B.n595 10.6151
R1115 B.n597 B.n596 10.6151
R1116 B.n597 B.n347 10.6151
R1117 B.n607 B.n347 10.6151
R1118 B.n608 B.n607 10.6151
R1119 B.n609 B.n608 10.6151
R1120 B.n609 B.n339 10.6151
R1121 B.n619 B.n339 10.6151
R1122 B.n620 B.n619 10.6151
R1123 B.n621 B.n620 10.6151
R1124 B.n621 B.n331 10.6151
R1125 B.n631 B.n331 10.6151
R1126 B.n632 B.n631 10.6151
R1127 B.n633 B.n632 10.6151
R1128 B.n633 B.n323 10.6151
R1129 B.n643 B.n323 10.6151
R1130 B.n644 B.n643 10.6151
R1131 B.n645 B.n644 10.6151
R1132 B.n645 B.n315 10.6151
R1133 B.n655 B.n315 10.6151
R1134 B.n656 B.n655 10.6151
R1135 B.n657 B.n656 10.6151
R1136 B.n657 B.n307 10.6151
R1137 B.n667 B.n307 10.6151
R1138 B.n668 B.n667 10.6151
R1139 B.n669 B.n668 10.6151
R1140 B.n669 B.n299 10.6151
R1141 B.n680 B.n299 10.6151
R1142 B.n681 B.n680 10.6151
R1143 B.n682 B.n681 10.6151
R1144 B.n682 B.n292 10.6151
R1145 B.n693 B.n292 10.6151
R1146 B.n694 B.n693 10.6151
R1147 B.n695 B.n694 10.6151
R1148 B.n695 B.n0 10.6151
R1149 B.n415 B.n363 10.6151
R1150 B.n416 B.n415 10.6151
R1151 B.n417 B.n416 10.6151
R1152 B.n417 B.n411 10.6151
R1153 B.n423 B.n411 10.6151
R1154 B.n424 B.n423 10.6151
R1155 B.n425 B.n424 10.6151
R1156 B.n425 B.n409 10.6151
R1157 B.n431 B.n409 10.6151
R1158 B.n432 B.n431 10.6151
R1159 B.n433 B.n432 10.6151
R1160 B.n433 B.n407 10.6151
R1161 B.n439 B.n407 10.6151
R1162 B.n440 B.n439 10.6151
R1163 B.n441 B.n440 10.6151
R1164 B.n441 B.n405 10.6151
R1165 B.n447 B.n405 10.6151
R1166 B.n448 B.n447 10.6151
R1167 B.n449 B.n448 10.6151
R1168 B.n449 B.n403 10.6151
R1169 B.n455 B.n403 10.6151
R1170 B.n456 B.n455 10.6151
R1171 B.n457 B.n456 10.6151
R1172 B.n457 B.n401 10.6151
R1173 B.n463 B.n401 10.6151
R1174 B.n464 B.n463 10.6151
R1175 B.n465 B.n464 10.6151
R1176 B.n465 B.n399 10.6151
R1177 B.n471 B.n399 10.6151
R1178 B.n472 B.n471 10.6151
R1179 B.n473 B.n472 10.6151
R1180 B.n473 B.n397 10.6151
R1181 B.n479 B.n397 10.6151
R1182 B.n480 B.n479 10.6151
R1183 B.n481 B.n480 10.6151
R1184 B.n481 B.n395 10.6151
R1185 B.n488 B.n487 10.6151
R1186 B.n489 B.n488 10.6151
R1187 B.n489 B.n390 10.6151
R1188 B.n495 B.n390 10.6151
R1189 B.n496 B.n495 10.6151
R1190 B.n497 B.n496 10.6151
R1191 B.n497 B.n388 10.6151
R1192 B.n503 B.n388 10.6151
R1193 B.n504 B.n503 10.6151
R1194 B.n506 B.n384 10.6151
R1195 B.n512 B.n384 10.6151
R1196 B.n513 B.n512 10.6151
R1197 B.n514 B.n513 10.6151
R1198 B.n514 B.n382 10.6151
R1199 B.n520 B.n382 10.6151
R1200 B.n521 B.n520 10.6151
R1201 B.n522 B.n521 10.6151
R1202 B.n522 B.n380 10.6151
R1203 B.n528 B.n380 10.6151
R1204 B.n529 B.n528 10.6151
R1205 B.n530 B.n529 10.6151
R1206 B.n530 B.n378 10.6151
R1207 B.n536 B.n378 10.6151
R1208 B.n537 B.n536 10.6151
R1209 B.n538 B.n537 10.6151
R1210 B.n538 B.n376 10.6151
R1211 B.n544 B.n376 10.6151
R1212 B.n545 B.n544 10.6151
R1213 B.n546 B.n545 10.6151
R1214 B.n546 B.n374 10.6151
R1215 B.n552 B.n374 10.6151
R1216 B.n553 B.n552 10.6151
R1217 B.n554 B.n553 10.6151
R1218 B.n554 B.n372 10.6151
R1219 B.n560 B.n372 10.6151
R1220 B.n561 B.n560 10.6151
R1221 B.n562 B.n561 10.6151
R1222 B.n562 B.n370 10.6151
R1223 B.n568 B.n370 10.6151
R1224 B.n569 B.n568 10.6151
R1225 B.n570 B.n569 10.6151
R1226 B.n570 B.n368 10.6151
R1227 B.n368 B.n367 10.6151
R1228 B.n577 B.n367 10.6151
R1229 B.n578 B.n577 10.6151
R1230 B.n579 B.n359 10.6151
R1231 B.n589 B.n359 10.6151
R1232 B.n590 B.n589 10.6151
R1233 B.n591 B.n590 10.6151
R1234 B.n591 B.n351 10.6151
R1235 B.n601 B.n351 10.6151
R1236 B.n602 B.n601 10.6151
R1237 B.n603 B.n602 10.6151
R1238 B.n603 B.n343 10.6151
R1239 B.n613 B.n343 10.6151
R1240 B.n614 B.n613 10.6151
R1241 B.n615 B.n614 10.6151
R1242 B.n615 B.n335 10.6151
R1243 B.n625 B.n335 10.6151
R1244 B.n626 B.n625 10.6151
R1245 B.n627 B.n626 10.6151
R1246 B.n627 B.n327 10.6151
R1247 B.n637 B.n327 10.6151
R1248 B.n638 B.n637 10.6151
R1249 B.n639 B.n638 10.6151
R1250 B.n639 B.n319 10.6151
R1251 B.n649 B.n319 10.6151
R1252 B.n650 B.n649 10.6151
R1253 B.n651 B.n650 10.6151
R1254 B.n651 B.n311 10.6151
R1255 B.n661 B.n311 10.6151
R1256 B.n662 B.n661 10.6151
R1257 B.n663 B.n662 10.6151
R1258 B.n663 B.n303 10.6151
R1259 B.n673 B.n303 10.6151
R1260 B.n674 B.n673 10.6151
R1261 B.n675 B.n674 10.6151
R1262 B.n675 B.n296 10.6151
R1263 B.n686 B.n296 10.6151
R1264 B.n687 B.n686 10.6151
R1265 B.n689 B.n687 10.6151
R1266 B.n689 B.n688 10.6151
R1267 B.n688 B.n288 10.6151
R1268 B.n700 B.n288 10.6151
R1269 B.n701 B.n700 10.6151
R1270 B.n702 B.n701 10.6151
R1271 B.n703 B.n702 10.6151
R1272 B.n704 B.n703 10.6151
R1273 B.n707 B.n704 10.6151
R1274 B.n708 B.n707 10.6151
R1275 B.n709 B.n708 10.6151
R1276 B.n710 B.n709 10.6151
R1277 B.n712 B.n710 10.6151
R1278 B.n713 B.n712 10.6151
R1279 B.n714 B.n713 10.6151
R1280 B.n715 B.n714 10.6151
R1281 B.n717 B.n715 10.6151
R1282 B.n718 B.n717 10.6151
R1283 B.n719 B.n718 10.6151
R1284 B.n720 B.n719 10.6151
R1285 B.n722 B.n720 10.6151
R1286 B.n723 B.n722 10.6151
R1287 B.n724 B.n723 10.6151
R1288 B.n725 B.n724 10.6151
R1289 B.n727 B.n725 10.6151
R1290 B.n728 B.n727 10.6151
R1291 B.n729 B.n728 10.6151
R1292 B.n730 B.n729 10.6151
R1293 B.n732 B.n730 10.6151
R1294 B.n733 B.n732 10.6151
R1295 B.n734 B.n733 10.6151
R1296 B.n735 B.n734 10.6151
R1297 B.n737 B.n735 10.6151
R1298 B.n738 B.n737 10.6151
R1299 B.n739 B.n738 10.6151
R1300 B.n740 B.n739 10.6151
R1301 B.n742 B.n740 10.6151
R1302 B.n743 B.n742 10.6151
R1303 B.n744 B.n743 10.6151
R1304 B.n745 B.n744 10.6151
R1305 B.n747 B.n745 10.6151
R1306 B.n748 B.n747 10.6151
R1307 B.n749 B.n748 10.6151
R1308 B.n750 B.n749 10.6151
R1309 B.n752 B.n750 10.6151
R1310 B.n753 B.n752 10.6151
R1311 B.n834 B.n1 10.6151
R1312 B.n834 B.n833 10.6151
R1313 B.n833 B.n832 10.6151
R1314 B.n832 B.n10 10.6151
R1315 B.n826 B.n10 10.6151
R1316 B.n826 B.n825 10.6151
R1317 B.n825 B.n824 10.6151
R1318 B.n824 B.n17 10.6151
R1319 B.n818 B.n17 10.6151
R1320 B.n818 B.n817 10.6151
R1321 B.n817 B.n816 10.6151
R1322 B.n816 B.n25 10.6151
R1323 B.n810 B.n25 10.6151
R1324 B.n810 B.n809 10.6151
R1325 B.n809 B.n808 10.6151
R1326 B.n808 B.n32 10.6151
R1327 B.n802 B.n32 10.6151
R1328 B.n802 B.n801 10.6151
R1329 B.n801 B.n800 10.6151
R1330 B.n800 B.n39 10.6151
R1331 B.n794 B.n39 10.6151
R1332 B.n794 B.n793 10.6151
R1333 B.n793 B.n792 10.6151
R1334 B.n792 B.n46 10.6151
R1335 B.n786 B.n46 10.6151
R1336 B.n786 B.n785 10.6151
R1337 B.n785 B.n784 10.6151
R1338 B.n784 B.n53 10.6151
R1339 B.n778 B.n53 10.6151
R1340 B.n778 B.n777 10.6151
R1341 B.n777 B.n776 10.6151
R1342 B.n776 B.n60 10.6151
R1343 B.n770 B.n60 10.6151
R1344 B.n770 B.n769 10.6151
R1345 B.n769 B.n768 10.6151
R1346 B.n768 B.n67 10.6151
R1347 B.n762 B.n67 10.6151
R1348 B.n762 B.n761 10.6151
R1349 B.n761 B.n760 10.6151
R1350 B.n123 B.n74 10.6151
R1351 B.n126 B.n123 10.6151
R1352 B.n127 B.n126 10.6151
R1353 B.n130 B.n127 10.6151
R1354 B.n131 B.n130 10.6151
R1355 B.n134 B.n131 10.6151
R1356 B.n135 B.n134 10.6151
R1357 B.n138 B.n135 10.6151
R1358 B.n139 B.n138 10.6151
R1359 B.n142 B.n139 10.6151
R1360 B.n143 B.n142 10.6151
R1361 B.n146 B.n143 10.6151
R1362 B.n147 B.n146 10.6151
R1363 B.n150 B.n147 10.6151
R1364 B.n151 B.n150 10.6151
R1365 B.n154 B.n151 10.6151
R1366 B.n155 B.n154 10.6151
R1367 B.n158 B.n155 10.6151
R1368 B.n159 B.n158 10.6151
R1369 B.n162 B.n159 10.6151
R1370 B.n163 B.n162 10.6151
R1371 B.n166 B.n163 10.6151
R1372 B.n167 B.n166 10.6151
R1373 B.n170 B.n167 10.6151
R1374 B.n171 B.n170 10.6151
R1375 B.n174 B.n171 10.6151
R1376 B.n175 B.n174 10.6151
R1377 B.n178 B.n175 10.6151
R1378 B.n179 B.n178 10.6151
R1379 B.n182 B.n179 10.6151
R1380 B.n183 B.n182 10.6151
R1381 B.n186 B.n183 10.6151
R1382 B.n187 B.n186 10.6151
R1383 B.n190 B.n187 10.6151
R1384 B.n191 B.n190 10.6151
R1385 B.n194 B.n191 10.6151
R1386 B.n199 B.n196 10.6151
R1387 B.n200 B.n199 10.6151
R1388 B.n203 B.n200 10.6151
R1389 B.n204 B.n203 10.6151
R1390 B.n207 B.n204 10.6151
R1391 B.n208 B.n207 10.6151
R1392 B.n211 B.n208 10.6151
R1393 B.n212 B.n211 10.6151
R1394 B.n215 B.n212 10.6151
R1395 B.n220 B.n217 10.6151
R1396 B.n221 B.n220 10.6151
R1397 B.n224 B.n221 10.6151
R1398 B.n225 B.n224 10.6151
R1399 B.n228 B.n225 10.6151
R1400 B.n229 B.n228 10.6151
R1401 B.n232 B.n229 10.6151
R1402 B.n233 B.n232 10.6151
R1403 B.n236 B.n233 10.6151
R1404 B.n237 B.n236 10.6151
R1405 B.n240 B.n237 10.6151
R1406 B.n241 B.n240 10.6151
R1407 B.n244 B.n241 10.6151
R1408 B.n245 B.n244 10.6151
R1409 B.n248 B.n245 10.6151
R1410 B.n249 B.n248 10.6151
R1411 B.n252 B.n249 10.6151
R1412 B.n253 B.n252 10.6151
R1413 B.n256 B.n253 10.6151
R1414 B.n257 B.n256 10.6151
R1415 B.n260 B.n257 10.6151
R1416 B.n261 B.n260 10.6151
R1417 B.n264 B.n261 10.6151
R1418 B.n265 B.n264 10.6151
R1419 B.n268 B.n265 10.6151
R1420 B.n269 B.n268 10.6151
R1421 B.n272 B.n269 10.6151
R1422 B.n273 B.n272 10.6151
R1423 B.n276 B.n273 10.6151
R1424 B.n277 B.n276 10.6151
R1425 B.n280 B.n277 10.6151
R1426 B.n281 B.n280 10.6151
R1427 B.n284 B.n281 10.6151
R1428 B.n286 B.n284 10.6151
R1429 B.n287 B.n286 10.6151
R1430 B.n754 B.n287 10.6151
R1431 B.n395 B.n394 9.36635
R1432 B.n506 B.n505 9.36635
R1433 B.n195 B.n194 9.36635
R1434 B.n217 B.n216 9.36635
R1435 B.n842 B.n0 8.11757
R1436 B.n842 B.n1 8.11757
R1437 B.n487 B.n394 1.24928
R1438 B.n505 B.n504 1.24928
R1439 B.n196 B.n195 1.24928
R1440 B.n216 B.n215 1.24928
R1441 VN.n1 VN.t1 110.731
R1442 VN.n0 VN.t3 110.731
R1443 VN.n0 VN.t2 109.599
R1444 VN.n1 VN.t0 109.599
R1445 VN VN.n1 50.2451
R1446 VN VN.n0 2.41559
R1447 VDD2.n2 VDD2.n0 102.374
R1448 VDD2.n2 VDD2.n1 60.0128
R1449 VDD2.n1 VDD2.t1 1.8755
R1450 VDD2.n1 VDD2.t2 1.8755
R1451 VDD2.n0 VDD2.t3 1.8755
R1452 VDD2.n0 VDD2.t0 1.8755
R1453 VDD2 VDD2.n2 0.0586897
R1454 VTAIL.n458 VTAIL.n406 289.615
R1455 VTAIL.n52 VTAIL.n0 289.615
R1456 VTAIL.n110 VTAIL.n58 289.615
R1457 VTAIL.n168 VTAIL.n116 289.615
R1458 VTAIL.n400 VTAIL.n348 289.615
R1459 VTAIL.n342 VTAIL.n290 289.615
R1460 VTAIL.n284 VTAIL.n232 289.615
R1461 VTAIL.n226 VTAIL.n174 289.615
R1462 VTAIL.n425 VTAIL.n424 185
R1463 VTAIL.n422 VTAIL.n421 185
R1464 VTAIL.n431 VTAIL.n430 185
R1465 VTAIL.n433 VTAIL.n432 185
R1466 VTAIL.n418 VTAIL.n417 185
R1467 VTAIL.n439 VTAIL.n438 185
R1468 VTAIL.n442 VTAIL.n441 185
R1469 VTAIL.n440 VTAIL.n414 185
R1470 VTAIL.n447 VTAIL.n413 185
R1471 VTAIL.n449 VTAIL.n448 185
R1472 VTAIL.n451 VTAIL.n450 185
R1473 VTAIL.n410 VTAIL.n409 185
R1474 VTAIL.n457 VTAIL.n456 185
R1475 VTAIL.n459 VTAIL.n458 185
R1476 VTAIL.n19 VTAIL.n18 185
R1477 VTAIL.n16 VTAIL.n15 185
R1478 VTAIL.n25 VTAIL.n24 185
R1479 VTAIL.n27 VTAIL.n26 185
R1480 VTAIL.n12 VTAIL.n11 185
R1481 VTAIL.n33 VTAIL.n32 185
R1482 VTAIL.n36 VTAIL.n35 185
R1483 VTAIL.n34 VTAIL.n8 185
R1484 VTAIL.n41 VTAIL.n7 185
R1485 VTAIL.n43 VTAIL.n42 185
R1486 VTAIL.n45 VTAIL.n44 185
R1487 VTAIL.n4 VTAIL.n3 185
R1488 VTAIL.n51 VTAIL.n50 185
R1489 VTAIL.n53 VTAIL.n52 185
R1490 VTAIL.n77 VTAIL.n76 185
R1491 VTAIL.n74 VTAIL.n73 185
R1492 VTAIL.n83 VTAIL.n82 185
R1493 VTAIL.n85 VTAIL.n84 185
R1494 VTAIL.n70 VTAIL.n69 185
R1495 VTAIL.n91 VTAIL.n90 185
R1496 VTAIL.n94 VTAIL.n93 185
R1497 VTAIL.n92 VTAIL.n66 185
R1498 VTAIL.n99 VTAIL.n65 185
R1499 VTAIL.n101 VTAIL.n100 185
R1500 VTAIL.n103 VTAIL.n102 185
R1501 VTAIL.n62 VTAIL.n61 185
R1502 VTAIL.n109 VTAIL.n108 185
R1503 VTAIL.n111 VTAIL.n110 185
R1504 VTAIL.n135 VTAIL.n134 185
R1505 VTAIL.n132 VTAIL.n131 185
R1506 VTAIL.n141 VTAIL.n140 185
R1507 VTAIL.n143 VTAIL.n142 185
R1508 VTAIL.n128 VTAIL.n127 185
R1509 VTAIL.n149 VTAIL.n148 185
R1510 VTAIL.n152 VTAIL.n151 185
R1511 VTAIL.n150 VTAIL.n124 185
R1512 VTAIL.n157 VTAIL.n123 185
R1513 VTAIL.n159 VTAIL.n158 185
R1514 VTAIL.n161 VTAIL.n160 185
R1515 VTAIL.n120 VTAIL.n119 185
R1516 VTAIL.n167 VTAIL.n166 185
R1517 VTAIL.n169 VTAIL.n168 185
R1518 VTAIL.n401 VTAIL.n400 185
R1519 VTAIL.n399 VTAIL.n398 185
R1520 VTAIL.n352 VTAIL.n351 185
R1521 VTAIL.n393 VTAIL.n392 185
R1522 VTAIL.n391 VTAIL.n390 185
R1523 VTAIL.n389 VTAIL.n355 185
R1524 VTAIL.n359 VTAIL.n356 185
R1525 VTAIL.n384 VTAIL.n383 185
R1526 VTAIL.n382 VTAIL.n381 185
R1527 VTAIL.n361 VTAIL.n360 185
R1528 VTAIL.n376 VTAIL.n375 185
R1529 VTAIL.n374 VTAIL.n373 185
R1530 VTAIL.n365 VTAIL.n364 185
R1531 VTAIL.n368 VTAIL.n367 185
R1532 VTAIL.n343 VTAIL.n342 185
R1533 VTAIL.n341 VTAIL.n340 185
R1534 VTAIL.n294 VTAIL.n293 185
R1535 VTAIL.n335 VTAIL.n334 185
R1536 VTAIL.n333 VTAIL.n332 185
R1537 VTAIL.n331 VTAIL.n297 185
R1538 VTAIL.n301 VTAIL.n298 185
R1539 VTAIL.n326 VTAIL.n325 185
R1540 VTAIL.n324 VTAIL.n323 185
R1541 VTAIL.n303 VTAIL.n302 185
R1542 VTAIL.n318 VTAIL.n317 185
R1543 VTAIL.n316 VTAIL.n315 185
R1544 VTAIL.n307 VTAIL.n306 185
R1545 VTAIL.n310 VTAIL.n309 185
R1546 VTAIL.n285 VTAIL.n284 185
R1547 VTAIL.n283 VTAIL.n282 185
R1548 VTAIL.n236 VTAIL.n235 185
R1549 VTAIL.n277 VTAIL.n276 185
R1550 VTAIL.n275 VTAIL.n274 185
R1551 VTAIL.n273 VTAIL.n239 185
R1552 VTAIL.n243 VTAIL.n240 185
R1553 VTAIL.n268 VTAIL.n267 185
R1554 VTAIL.n266 VTAIL.n265 185
R1555 VTAIL.n245 VTAIL.n244 185
R1556 VTAIL.n260 VTAIL.n259 185
R1557 VTAIL.n258 VTAIL.n257 185
R1558 VTAIL.n249 VTAIL.n248 185
R1559 VTAIL.n252 VTAIL.n251 185
R1560 VTAIL.n227 VTAIL.n226 185
R1561 VTAIL.n225 VTAIL.n224 185
R1562 VTAIL.n178 VTAIL.n177 185
R1563 VTAIL.n219 VTAIL.n218 185
R1564 VTAIL.n217 VTAIL.n216 185
R1565 VTAIL.n215 VTAIL.n181 185
R1566 VTAIL.n185 VTAIL.n182 185
R1567 VTAIL.n210 VTAIL.n209 185
R1568 VTAIL.n208 VTAIL.n207 185
R1569 VTAIL.n187 VTAIL.n186 185
R1570 VTAIL.n202 VTAIL.n201 185
R1571 VTAIL.n200 VTAIL.n199 185
R1572 VTAIL.n191 VTAIL.n190 185
R1573 VTAIL.n194 VTAIL.n193 185
R1574 VTAIL.t3 VTAIL.n423 149.524
R1575 VTAIL.t2 VTAIL.n17 149.524
R1576 VTAIL.t6 VTAIL.n75 149.524
R1577 VTAIL.t0 VTAIL.n133 149.524
R1578 VTAIL.t1 VTAIL.n366 149.524
R1579 VTAIL.t7 VTAIL.n308 149.524
R1580 VTAIL.t4 VTAIL.n250 149.524
R1581 VTAIL.t5 VTAIL.n192 149.524
R1582 VTAIL.n424 VTAIL.n421 104.615
R1583 VTAIL.n431 VTAIL.n421 104.615
R1584 VTAIL.n432 VTAIL.n431 104.615
R1585 VTAIL.n432 VTAIL.n417 104.615
R1586 VTAIL.n439 VTAIL.n417 104.615
R1587 VTAIL.n441 VTAIL.n439 104.615
R1588 VTAIL.n441 VTAIL.n440 104.615
R1589 VTAIL.n440 VTAIL.n413 104.615
R1590 VTAIL.n449 VTAIL.n413 104.615
R1591 VTAIL.n450 VTAIL.n449 104.615
R1592 VTAIL.n450 VTAIL.n409 104.615
R1593 VTAIL.n457 VTAIL.n409 104.615
R1594 VTAIL.n458 VTAIL.n457 104.615
R1595 VTAIL.n18 VTAIL.n15 104.615
R1596 VTAIL.n25 VTAIL.n15 104.615
R1597 VTAIL.n26 VTAIL.n25 104.615
R1598 VTAIL.n26 VTAIL.n11 104.615
R1599 VTAIL.n33 VTAIL.n11 104.615
R1600 VTAIL.n35 VTAIL.n33 104.615
R1601 VTAIL.n35 VTAIL.n34 104.615
R1602 VTAIL.n34 VTAIL.n7 104.615
R1603 VTAIL.n43 VTAIL.n7 104.615
R1604 VTAIL.n44 VTAIL.n43 104.615
R1605 VTAIL.n44 VTAIL.n3 104.615
R1606 VTAIL.n51 VTAIL.n3 104.615
R1607 VTAIL.n52 VTAIL.n51 104.615
R1608 VTAIL.n76 VTAIL.n73 104.615
R1609 VTAIL.n83 VTAIL.n73 104.615
R1610 VTAIL.n84 VTAIL.n83 104.615
R1611 VTAIL.n84 VTAIL.n69 104.615
R1612 VTAIL.n91 VTAIL.n69 104.615
R1613 VTAIL.n93 VTAIL.n91 104.615
R1614 VTAIL.n93 VTAIL.n92 104.615
R1615 VTAIL.n92 VTAIL.n65 104.615
R1616 VTAIL.n101 VTAIL.n65 104.615
R1617 VTAIL.n102 VTAIL.n101 104.615
R1618 VTAIL.n102 VTAIL.n61 104.615
R1619 VTAIL.n109 VTAIL.n61 104.615
R1620 VTAIL.n110 VTAIL.n109 104.615
R1621 VTAIL.n134 VTAIL.n131 104.615
R1622 VTAIL.n141 VTAIL.n131 104.615
R1623 VTAIL.n142 VTAIL.n141 104.615
R1624 VTAIL.n142 VTAIL.n127 104.615
R1625 VTAIL.n149 VTAIL.n127 104.615
R1626 VTAIL.n151 VTAIL.n149 104.615
R1627 VTAIL.n151 VTAIL.n150 104.615
R1628 VTAIL.n150 VTAIL.n123 104.615
R1629 VTAIL.n159 VTAIL.n123 104.615
R1630 VTAIL.n160 VTAIL.n159 104.615
R1631 VTAIL.n160 VTAIL.n119 104.615
R1632 VTAIL.n167 VTAIL.n119 104.615
R1633 VTAIL.n168 VTAIL.n167 104.615
R1634 VTAIL.n400 VTAIL.n399 104.615
R1635 VTAIL.n399 VTAIL.n351 104.615
R1636 VTAIL.n392 VTAIL.n351 104.615
R1637 VTAIL.n392 VTAIL.n391 104.615
R1638 VTAIL.n391 VTAIL.n355 104.615
R1639 VTAIL.n359 VTAIL.n355 104.615
R1640 VTAIL.n383 VTAIL.n359 104.615
R1641 VTAIL.n383 VTAIL.n382 104.615
R1642 VTAIL.n382 VTAIL.n360 104.615
R1643 VTAIL.n375 VTAIL.n360 104.615
R1644 VTAIL.n375 VTAIL.n374 104.615
R1645 VTAIL.n374 VTAIL.n364 104.615
R1646 VTAIL.n367 VTAIL.n364 104.615
R1647 VTAIL.n342 VTAIL.n341 104.615
R1648 VTAIL.n341 VTAIL.n293 104.615
R1649 VTAIL.n334 VTAIL.n293 104.615
R1650 VTAIL.n334 VTAIL.n333 104.615
R1651 VTAIL.n333 VTAIL.n297 104.615
R1652 VTAIL.n301 VTAIL.n297 104.615
R1653 VTAIL.n325 VTAIL.n301 104.615
R1654 VTAIL.n325 VTAIL.n324 104.615
R1655 VTAIL.n324 VTAIL.n302 104.615
R1656 VTAIL.n317 VTAIL.n302 104.615
R1657 VTAIL.n317 VTAIL.n316 104.615
R1658 VTAIL.n316 VTAIL.n306 104.615
R1659 VTAIL.n309 VTAIL.n306 104.615
R1660 VTAIL.n284 VTAIL.n283 104.615
R1661 VTAIL.n283 VTAIL.n235 104.615
R1662 VTAIL.n276 VTAIL.n235 104.615
R1663 VTAIL.n276 VTAIL.n275 104.615
R1664 VTAIL.n275 VTAIL.n239 104.615
R1665 VTAIL.n243 VTAIL.n239 104.615
R1666 VTAIL.n267 VTAIL.n243 104.615
R1667 VTAIL.n267 VTAIL.n266 104.615
R1668 VTAIL.n266 VTAIL.n244 104.615
R1669 VTAIL.n259 VTAIL.n244 104.615
R1670 VTAIL.n259 VTAIL.n258 104.615
R1671 VTAIL.n258 VTAIL.n248 104.615
R1672 VTAIL.n251 VTAIL.n248 104.615
R1673 VTAIL.n226 VTAIL.n225 104.615
R1674 VTAIL.n225 VTAIL.n177 104.615
R1675 VTAIL.n218 VTAIL.n177 104.615
R1676 VTAIL.n218 VTAIL.n217 104.615
R1677 VTAIL.n217 VTAIL.n181 104.615
R1678 VTAIL.n185 VTAIL.n181 104.615
R1679 VTAIL.n209 VTAIL.n185 104.615
R1680 VTAIL.n209 VTAIL.n208 104.615
R1681 VTAIL.n208 VTAIL.n186 104.615
R1682 VTAIL.n201 VTAIL.n186 104.615
R1683 VTAIL.n201 VTAIL.n200 104.615
R1684 VTAIL.n200 VTAIL.n190 104.615
R1685 VTAIL.n193 VTAIL.n190 104.615
R1686 VTAIL.n424 VTAIL.t3 52.3082
R1687 VTAIL.n18 VTAIL.t2 52.3082
R1688 VTAIL.n76 VTAIL.t6 52.3082
R1689 VTAIL.n134 VTAIL.t0 52.3082
R1690 VTAIL.n367 VTAIL.t1 52.3082
R1691 VTAIL.n309 VTAIL.t7 52.3082
R1692 VTAIL.n251 VTAIL.t4 52.3082
R1693 VTAIL.n193 VTAIL.t5 52.3082
R1694 VTAIL.n463 VTAIL.n462 29.8581
R1695 VTAIL.n57 VTAIL.n56 29.8581
R1696 VTAIL.n115 VTAIL.n114 29.8581
R1697 VTAIL.n173 VTAIL.n172 29.8581
R1698 VTAIL.n405 VTAIL.n404 29.8581
R1699 VTAIL.n347 VTAIL.n346 29.8581
R1700 VTAIL.n289 VTAIL.n288 29.8581
R1701 VTAIL.n231 VTAIL.n230 29.8581
R1702 VTAIL.n463 VTAIL.n405 24.6514
R1703 VTAIL.n231 VTAIL.n173 24.6514
R1704 VTAIL.n448 VTAIL.n447 13.1884
R1705 VTAIL.n42 VTAIL.n41 13.1884
R1706 VTAIL.n100 VTAIL.n99 13.1884
R1707 VTAIL.n158 VTAIL.n157 13.1884
R1708 VTAIL.n390 VTAIL.n389 13.1884
R1709 VTAIL.n332 VTAIL.n331 13.1884
R1710 VTAIL.n274 VTAIL.n273 13.1884
R1711 VTAIL.n216 VTAIL.n215 13.1884
R1712 VTAIL.n446 VTAIL.n414 12.8005
R1713 VTAIL.n451 VTAIL.n412 12.8005
R1714 VTAIL.n40 VTAIL.n8 12.8005
R1715 VTAIL.n45 VTAIL.n6 12.8005
R1716 VTAIL.n98 VTAIL.n66 12.8005
R1717 VTAIL.n103 VTAIL.n64 12.8005
R1718 VTAIL.n156 VTAIL.n124 12.8005
R1719 VTAIL.n161 VTAIL.n122 12.8005
R1720 VTAIL.n393 VTAIL.n354 12.8005
R1721 VTAIL.n388 VTAIL.n356 12.8005
R1722 VTAIL.n335 VTAIL.n296 12.8005
R1723 VTAIL.n330 VTAIL.n298 12.8005
R1724 VTAIL.n277 VTAIL.n238 12.8005
R1725 VTAIL.n272 VTAIL.n240 12.8005
R1726 VTAIL.n219 VTAIL.n180 12.8005
R1727 VTAIL.n214 VTAIL.n182 12.8005
R1728 VTAIL.n443 VTAIL.n442 12.0247
R1729 VTAIL.n452 VTAIL.n410 12.0247
R1730 VTAIL.n37 VTAIL.n36 12.0247
R1731 VTAIL.n46 VTAIL.n4 12.0247
R1732 VTAIL.n95 VTAIL.n94 12.0247
R1733 VTAIL.n104 VTAIL.n62 12.0247
R1734 VTAIL.n153 VTAIL.n152 12.0247
R1735 VTAIL.n162 VTAIL.n120 12.0247
R1736 VTAIL.n394 VTAIL.n352 12.0247
R1737 VTAIL.n385 VTAIL.n384 12.0247
R1738 VTAIL.n336 VTAIL.n294 12.0247
R1739 VTAIL.n327 VTAIL.n326 12.0247
R1740 VTAIL.n278 VTAIL.n236 12.0247
R1741 VTAIL.n269 VTAIL.n268 12.0247
R1742 VTAIL.n220 VTAIL.n178 12.0247
R1743 VTAIL.n211 VTAIL.n210 12.0247
R1744 VTAIL.n438 VTAIL.n416 11.249
R1745 VTAIL.n456 VTAIL.n455 11.249
R1746 VTAIL.n32 VTAIL.n10 11.249
R1747 VTAIL.n50 VTAIL.n49 11.249
R1748 VTAIL.n90 VTAIL.n68 11.249
R1749 VTAIL.n108 VTAIL.n107 11.249
R1750 VTAIL.n148 VTAIL.n126 11.249
R1751 VTAIL.n166 VTAIL.n165 11.249
R1752 VTAIL.n398 VTAIL.n397 11.249
R1753 VTAIL.n381 VTAIL.n358 11.249
R1754 VTAIL.n340 VTAIL.n339 11.249
R1755 VTAIL.n323 VTAIL.n300 11.249
R1756 VTAIL.n282 VTAIL.n281 11.249
R1757 VTAIL.n265 VTAIL.n242 11.249
R1758 VTAIL.n224 VTAIL.n223 11.249
R1759 VTAIL.n207 VTAIL.n184 11.249
R1760 VTAIL.n437 VTAIL.n418 10.4732
R1761 VTAIL.n459 VTAIL.n408 10.4732
R1762 VTAIL.n31 VTAIL.n12 10.4732
R1763 VTAIL.n53 VTAIL.n2 10.4732
R1764 VTAIL.n89 VTAIL.n70 10.4732
R1765 VTAIL.n111 VTAIL.n60 10.4732
R1766 VTAIL.n147 VTAIL.n128 10.4732
R1767 VTAIL.n169 VTAIL.n118 10.4732
R1768 VTAIL.n401 VTAIL.n350 10.4732
R1769 VTAIL.n380 VTAIL.n361 10.4732
R1770 VTAIL.n343 VTAIL.n292 10.4732
R1771 VTAIL.n322 VTAIL.n303 10.4732
R1772 VTAIL.n285 VTAIL.n234 10.4732
R1773 VTAIL.n264 VTAIL.n245 10.4732
R1774 VTAIL.n227 VTAIL.n176 10.4732
R1775 VTAIL.n206 VTAIL.n187 10.4732
R1776 VTAIL.n425 VTAIL.n423 10.2747
R1777 VTAIL.n19 VTAIL.n17 10.2747
R1778 VTAIL.n77 VTAIL.n75 10.2747
R1779 VTAIL.n135 VTAIL.n133 10.2747
R1780 VTAIL.n368 VTAIL.n366 10.2747
R1781 VTAIL.n310 VTAIL.n308 10.2747
R1782 VTAIL.n252 VTAIL.n250 10.2747
R1783 VTAIL.n194 VTAIL.n192 10.2747
R1784 VTAIL.n434 VTAIL.n433 9.69747
R1785 VTAIL.n460 VTAIL.n406 9.69747
R1786 VTAIL.n28 VTAIL.n27 9.69747
R1787 VTAIL.n54 VTAIL.n0 9.69747
R1788 VTAIL.n86 VTAIL.n85 9.69747
R1789 VTAIL.n112 VTAIL.n58 9.69747
R1790 VTAIL.n144 VTAIL.n143 9.69747
R1791 VTAIL.n170 VTAIL.n116 9.69747
R1792 VTAIL.n402 VTAIL.n348 9.69747
R1793 VTAIL.n377 VTAIL.n376 9.69747
R1794 VTAIL.n344 VTAIL.n290 9.69747
R1795 VTAIL.n319 VTAIL.n318 9.69747
R1796 VTAIL.n286 VTAIL.n232 9.69747
R1797 VTAIL.n261 VTAIL.n260 9.69747
R1798 VTAIL.n228 VTAIL.n174 9.69747
R1799 VTAIL.n203 VTAIL.n202 9.69747
R1800 VTAIL.n462 VTAIL.n461 9.45567
R1801 VTAIL.n56 VTAIL.n55 9.45567
R1802 VTAIL.n114 VTAIL.n113 9.45567
R1803 VTAIL.n172 VTAIL.n171 9.45567
R1804 VTAIL.n404 VTAIL.n403 9.45567
R1805 VTAIL.n346 VTAIL.n345 9.45567
R1806 VTAIL.n288 VTAIL.n287 9.45567
R1807 VTAIL.n230 VTAIL.n229 9.45567
R1808 VTAIL.n461 VTAIL.n460 9.3005
R1809 VTAIL.n408 VTAIL.n407 9.3005
R1810 VTAIL.n455 VTAIL.n454 9.3005
R1811 VTAIL.n453 VTAIL.n452 9.3005
R1812 VTAIL.n412 VTAIL.n411 9.3005
R1813 VTAIL.n427 VTAIL.n426 9.3005
R1814 VTAIL.n429 VTAIL.n428 9.3005
R1815 VTAIL.n420 VTAIL.n419 9.3005
R1816 VTAIL.n435 VTAIL.n434 9.3005
R1817 VTAIL.n437 VTAIL.n436 9.3005
R1818 VTAIL.n416 VTAIL.n415 9.3005
R1819 VTAIL.n444 VTAIL.n443 9.3005
R1820 VTAIL.n446 VTAIL.n445 9.3005
R1821 VTAIL.n55 VTAIL.n54 9.3005
R1822 VTAIL.n2 VTAIL.n1 9.3005
R1823 VTAIL.n49 VTAIL.n48 9.3005
R1824 VTAIL.n47 VTAIL.n46 9.3005
R1825 VTAIL.n6 VTAIL.n5 9.3005
R1826 VTAIL.n21 VTAIL.n20 9.3005
R1827 VTAIL.n23 VTAIL.n22 9.3005
R1828 VTAIL.n14 VTAIL.n13 9.3005
R1829 VTAIL.n29 VTAIL.n28 9.3005
R1830 VTAIL.n31 VTAIL.n30 9.3005
R1831 VTAIL.n10 VTAIL.n9 9.3005
R1832 VTAIL.n38 VTAIL.n37 9.3005
R1833 VTAIL.n40 VTAIL.n39 9.3005
R1834 VTAIL.n113 VTAIL.n112 9.3005
R1835 VTAIL.n60 VTAIL.n59 9.3005
R1836 VTAIL.n107 VTAIL.n106 9.3005
R1837 VTAIL.n105 VTAIL.n104 9.3005
R1838 VTAIL.n64 VTAIL.n63 9.3005
R1839 VTAIL.n79 VTAIL.n78 9.3005
R1840 VTAIL.n81 VTAIL.n80 9.3005
R1841 VTAIL.n72 VTAIL.n71 9.3005
R1842 VTAIL.n87 VTAIL.n86 9.3005
R1843 VTAIL.n89 VTAIL.n88 9.3005
R1844 VTAIL.n68 VTAIL.n67 9.3005
R1845 VTAIL.n96 VTAIL.n95 9.3005
R1846 VTAIL.n98 VTAIL.n97 9.3005
R1847 VTAIL.n171 VTAIL.n170 9.3005
R1848 VTAIL.n118 VTAIL.n117 9.3005
R1849 VTAIL.n165 VTAIL.n164 9.3005
R1850 VTAIL.n163 VTAIL.n162 9.3005
R1851 VTAIL.n122 VTAIL.n121 9.3005
R1852 VTAIL.n137 VTAIL.n136 9.3005
R1853 VTAIL.n139 VTAIL.n138 9.3005
R1854 VTAIL.n130 VTAIL.n129 9.3005
R1855 VTAIL.n145 VTAIL.n144 9.3005
R1856 VTAIL.n147 VTAIL.n146 9.3005
R1857 VTAIL.n126 VTAIL.n125 9.3005
R1858 VTAIL.n154 VTAIL.n153 9.3005
R1859 VTAIL.n156 VTAIL.n155 9.3005
R1860 VTAIL.n370 VTAIL.n369 9.3005
R1861 VTAIL.n372 VTAIL.n371 9.3005
R1862 VTAIL.n363 VTAIL.n362 9.3005
R1863 VTAIL.n378 VTAIL.n377 9.3005
R1864 VTAIL.n380 VTAIL.n379 9.3005
R1865 VTAIL.n358 VTAIL.n357 9.3005
R1866 VTAIL.n386 VTAIL.n385 9.3005
R1867 VTAIL.n388 VTAIL.n387 9.3005
R1868 VTAIL.n403 VTAIL.n402 9.3005
R1869 VTAIL.n350 VTAIL.n349 9.3005
R1870 VTAIL.n397 VTAIL.n396 9.3005
R1871 VTAIL.n395 VTAIL.n394 9.3005
R1872 VTAIL.n354 VTAIL.n353 9.3005
R1873 VTAIL.n312 VTAIL.n311 9.3005
R1874 VTAIL.n314 VTAIL.n313 9.3005
R1875 VTAIL.n305 VTAIL.n304 9.3005
R1876 VTAIL.n320 VTAIL.n319 9.3005
R1877 VTAIL.n322 VTAIL.n321 9.3005
R1878 VTAIL.n300 VTAIL.n299 9.3005
R1879 VTAIL.n328 VTAIL.n327 9.3005
R1880 VTAIL.n330 VTAIL.n329 9.3005
R1881 VTAIL.n345 VTAIL.n344 9.3005
R1882 VTAIL.n292 VTAIL.n291 9.3005
R1883 VTAIL.n339 VTAIL.n338 9.3005
R1884 VTAIL.n337 VTAIL.n336 9.3005
R1885 VTAIL.n296 VTAIL.n295 9.3005
R1886 VTAIL.n254 VTAIL.n253 9.3005
R1887 VTAIL.n256 VTAIL.n255 9.3005
R1888 VTAIL.n247 VTAIL.n246 9.3005
R1889 VTAIL.n262 VTAIL.n261 9.3005
R1890 VTAIL.n264 VTAIL.n263 9.3005
R1891 VTAIL.n242 VTAIL.n241 9.3005
R1892 VTAIL.n270 VTAIL.n269 9.3005
R1893 VTAIL.n272 VTAIL.n271 9.3005
R1894 VTAIL.n287 VTAIL.n286 9.3005
R1895 VTAIL.n234 VTAIL.n233 9.3005
R1896 VTAIL.n281 VTAIL.n280 9.3005
R1897 VTAIL.n279 VTAIL.n278 9.3005
R1898 VTAIL.n238 VTAIL.n237 9.3005
R1899 VTAIL.n196 VTAIL.n195 9.3005
R1900 VTAIL.n198 VTAIL.n197 9.3005
R1901 VTAIL.n189 VTAIL.n188 9.3005
R1902 VTAIL.n204 VTAIL.n203 9.3005
R1903 VTAIL.n206 VTAIL.n205 9.3005
R1904 VTAIL.n184 VTAIL.n183 9.3005
R1905 VTAIL.n212 VTAIL.n211 9.3005
R1906 VTAIL.n214 VTAIL.n213 9.3005
R1907 VTAIL.n229 VTAIL.n228 9.3005
R1908 VTAIL.n176 VTAIL.n175 9.3005
R1909 VTAIL.n223 VTAIL.n222 9.3005
R1910 VTAIL.n221 VTAIL.n220 9.3005
R1911 VTAIL.n180 VTAIL.n179 9.3005
R1912 VTAIL.n430 VTAIL.n420 8.92171
R1913 VTAIL.n24 VTAIL.n14 8.92171
R1914 VTAIL.n82 VTAIL.n72 8.92171
R1915 VTAIL.n140 VTAIL.n130 8.92171
R1916 VTAIL.n373 VTAIL.n363 8.92171
R1917 VTAIL.n315 VTAIL.n305 8.92171
R1918 VTAIL.n257 VTAIL.n247 8.92171
R1919 VTAIL.n199 VTAIL.n189 8.92171
R1920 VTAIL.n429 VTAIL.n422 8.14595
R1921 VTAIL.n23 VTAIL.n16 8.14595
R1922 VTAIL.n81 VTAIL.n74 8.14595
R1923 VTAIL.n139 VTAIL.n132 8.14595
R1924 VTAIL.n372 VTAIL.n365 8.14595
R1925 VTAIL.n314 VTAIL.n307 8.14595
R1926 VTAIL.n256 VTAIL.n249 8.14595
R1927 VTAIL.n198 VTAIL.n191 8.14595
R1928 VTAIL.n426 VTAIL.n425 7.3702
R1929 VTAIL.n20 VTAIL.n19 7.3702
R1930 VTAIL.n78 VTAIL.n77 7.3702
R1931 VTAIL.n136 VTAIL.n135 7.3702
R1932 VTAIL.n369 VTAIL.n368 7.3702
R1933 VTAIL.n311 VTAIL.n310 7.3702
R1934 VTAIL.n253 VTAIL.n252 7.3702
R1935 VTAIL.n195 VTAIL.n194 7.3702
R1936 VTAIL.n426 VTAIL.n422 5.81868
R1937 VTAIL.n20 VTAIL.n16 5.81868
R1938 VTAIL.n78 VTAIL.n74 5.81868
R1939 VTAIL.n136 VTAIL.n132 5.81868
R1940 VTAIL.n369 VTAIL.n365 5.81868
R1941 VTAIL.n311 VTAIL.n307 5.81868
R1942 VTAIL.n253 VTAIL.n249 5.81868
R1943 VTAIL.n195 VTAIL.n191 5.81868
R1944 VTAIL.n430 VTAIL.n429 5.04292
R1945 VTAIL.n24 VTAIL.n23 5.04292
R1946 VTAIL.n82 VTAIL.n81 5.04292
R1947 VTAIL.n140 VTAIL.n139 5.04292
R1948 VTAIL.n373 VTAIL.n372 5.04292
R1949 VTAIL.n315 VTAIL.n314 5.04292
R1950 VTAIL.n257 VTAIL.n256 5.04292
R1951 VTAIL.n199 VTAIL.n198 5.04292
R1952 VTAIL.n433 VTAIL.n420 4.26717
R1953 VTAIL.n462 VTAIL.n406 4.26717
R1954 VTAIL.n27 VTAIL.n14 4.26717
R1955 VTAIL.n56 VTAIL.n0 4.26717
R1956 VTAIL.n85 VTAIL.n72 4.26717
R1957 VTAIL.n114 VTAIL.n58 4.26717
R1958 VTAIL.n143 VTAIL.n130 4.26717
R1959 VTAIL.n172 VTAIL.n116 4.26717
R1960 VTAIL.n404 VTAIL.n348 4.26717
R1961 VTAIL.n376 VTAIL.n363 4.26717
R1962 VTAIL.n346 VTAIL.n290 4.26717
R1963 VTAIL.n318 VTAIL.n305 4.26717
R1964 VTAIL.n288 VTAIL.n232 4.26717
R1965 VTAIL.n260 VTAIL.n247 4.26717
R1966 VTAIL.n230 VTAIL.n174 4.26717
R1967 VTAIL.n202 VTAIL.n189 4.26717
R1968 VTAIL.n434 VTAIL.n418 3.49141
R1969 VTAIL.n460 VTAIL.n459 3.49141
R1970 VTAIL.n28 VTAIL.n12 3.49141
R1971 VTAIL.n54 VTAIL.n53 3.49141
R1972 VTAIL.n86 VTAIL.n70 3.49141
R1973 VTAIL.n112 VTAIL.n111 3.49141
R1974 VTAIL.n144 VTAIL.n128 3.49141
R1975 VTAIL.n170 VTAIL.n169 3.49141
R1976 VTAIL.n402 VTAIL.n401 3.49141
R1977 VTAIL.n377 VTAIL.n361 3.49141
R1978 VTAIL.n344 VTAIL.n343 3.49141
R1979 VTAIL.n319 VTAIL.n303 3.49141
R1980 VTAIL.n286 VTAIL.n285 3.49141
R1981 VTAIL.n261 VTAIL.n245 3.49141
R1982 VTAIL.n228 VTAIL.n227 3.49141
R1983 VTAIL.n203 VTAIL.n187 3.49141
R1984 VTAIL.n289 VTAIL.n231 3.18153
R1985 VTAIL.n405 VTAIL.n347 3.18153
R1986 VTAIL.n173 VTAIL.n115 3.18153
R1987 VTAIL.n427 VTAIL.n423 2.84303
R1988 VTAIL.n21 VTAIL.n17 2.84303
R1989 VTAIL.n79 VTAIL.n75 2.84303
R1990 VTAIL.n137 VTAIL.n133 2.84303
R1991 VTAIL.n370 VTAIL.n366 2.84303
R1992 VTAIL.n312 VTAIL.n308 2.84303
R1993 VTAIL.n254 VTAIL.n250 2.84303
R1994 VTAIL.n196 VTAIL.n192 2.84303
R1995 VTAIL.n438 VTAIL.n437 2.71565
R1996 VTAIL.n456 VTAIL.n408 2.71565
R1997 VTAIL.n32 VTAIL.n31 2.71565
R1998 VTAIL.n50 VTAIL.n2 2.71565
R1999 VTAIL.n90 VTAIL.n89 2.71565
R2000 VTAIL.n108 VTAIL.n60 2.71565
R2001 VTAIL.n148 VTAIL.n147 2.71565
R2002 VTAIL.n166 VTAIL.n118 2.71565
R2003 VTAIL.n398 VTAIL.n350 2.71565
R2004 VTAIL.n381 VTAIL.n380 2.71565
R2005 VTAIL.n340 VTAIL.n292 2.71565
R2006 VTAIL.n323 VTAIL.n322 2.71565
R2007 VTAIL.n282 VTAIL.n234 2.71565
R2008 VTAIL.n265 VTAIL.n264 2.71565
R2009 VTAIL.n224 VTAIL.n176 2.71565
R2010 VTAIL.n207 VTAIL.n206 2.71565
R2011 VTAIL.n442 VTAIL.n416 1.93989
R2012 VTAIL.n455 VTAIL.n410 1.93989
R2013 VTAIL.n36 VTAIL.n10 1.93989
R2014 VTAIL.n49 VTAIL.n4 1.93989
R2015 VTAIL.n94 VTAIL.n68 1.93989
R2016 VTAIL.n107 VTAIL.n62 1.93989
R2017 VTAIL.n152 VTAIL.n126 1.93989
R2018 VTAIL.n165 VTAIL.n120 1.93989
R2019 VTAIL.n397 VTAIL.n352 1.93989
R2020 VTAIL.n384 VTAIL.n358 1.93989
R2021 VTAIL.n339 VTAIL.n294 1.93989
R2022 VTAIL.n326 VTAIL.n300 1.93989
R2023 VTAIL.n281 VTAIL.n236 1.93989
R2024 VTAIL.n268 VTAIL.n242 1.93989
R2025 VTAIL.n223 VTAIL.n178 1.93989
R2026 VTAIL.n210 VTAIL.n184 1.93989
R2027 VTAIL VTAIL.n57 1.64921
R2028 VTAIL VTAIL.n463 1.53283
R2029 VTAIL.n443 VTAIL.n414 1.16414
R2030 VTAIL.n452 VTAIL.n451 1.16414
R2031 VTAIL.n37 VTAIL.n8 1.16414
R2032 VTAIL.n46 VTAIL.n45 1.16414
R2033 VTAIL.n95 VTAIL.n66 1.16414
R2034 VTAIL.n104 VTAIL.n103 1.16414
R2035 VTAIL.n153 VTAIL.n124 1.16414
R2036 VTAIL.n162 VTAIL.n161 1.16414
R2037 VTAIL.n394 VTAIL.n393 1.16414
R2038 VTAIL.n385 VTAIL.n356 1.16414
R2039 VTAIL.n336 VTAIL.n335 1.16414
R2040 VTAIL.n327 VTAIL.n298 1.16414
R2041 VTAIL.n278 VTAIL.n277 1.16414
R2042 VTAIL.n269 VTAIL.n240 1.16414
R2043 VTAIL.n220 VTAIL.n219 1.16414
R2044 VTAIL.n211 VTAIL.n182 1.16414
R2045 VTAIL.n347 VTAIL.n289 0.470328
R2046 VTAIL.n115 VTAIL.n57 0.470328
R2047 VTAIL.n447 VTAIL.n446 0.388379
R2048 VTAIL.n448 VTAIL.n412 0.388379
R2049 VTAIL.n41 VTAIL.n40 0.388379
R2050 VTAIL.n42 VTAIL.n6 0.388379
R2051 VTAIL.n99 VTAIL.n98 0.388379
R2052 VTAIL.n100 VTAIL.n64 0.388379
R2053 VTAIL.n157 VTAIL.n156 0.388379
R2054 VTAIL.n158 VTAIL.n122 0.388379
R2055 VTAIL.n390 VTAIL.n354 0.388379
R2056 VTAIL.n389 VTAIL.n388 0.388379
R2057 VTAIL.n332 VTAIL.n296 0.388379
R2058 VTAIL.n331 VTAIL.n330 0.388379
R2059 VTAIL.n274 VTAIL.n238 0.388379
R2060 VTAIL.n273 VTAIL.n272 0.388379
R2061 VTAIL.n216 VTAIL.n180 0.388379
R2062 VTAIL.n215 VTAIL.n214 0.388379
R2063 VTAIL.n428 VTAIL.n427 0.155672
R2064 VTAIL.n428 VTAIL.n419 0.155672
R2065 VTAIL.n435 VTAIL.n419 0.155672
R2066 VTAIL.n436 VTAIL.n435 0.155672
R2067 VTAIL.n436 VTAIL.n415 0.155672
R2068 VTAIL.n444 VTAIL.n415 0.155672
R2069 VTAIL.n445 VTAIL.n444 0.155672
R2070 VTAIL.n445 VTAIL.n411 0.155672
R2071 VTAIL.n453 VTAIL.n411 0.155672
R2072 VTAIL.n454 VTAIL.n453 0.155672
R2073 VTAIL.n454 VTAIL.n407 0.155672
R2074 VTAIL.n461 VTAIL.n407 0.155672
R2075 VTAIL.n22 VTAIL.n21 0.155672
R2076 VTAIL.n22 VTAIL.n13 0.155672
R2077 VTAIL.n29 VTAIL.n13 0.155672
R2078 VTAIL.n30 VTAIL.n29 0.155672
R2079 VTAIL.n30 VTAIL.n9 0.155672
R2080 VTAIL.n38 VTAIL.n9 0.155672
R2081 VTAIL.n39 VTAIL.n38 0.155672
R2082 VTAIL.n39 VTAIL.n5 0.155672
R2083 VTAIL.n47 VTAIL.n5 0.155672
R2084 VTAIL.n48 VTAIL.n47 0.155672
R2085 VTAIL.n48 VTAIL.n1 0.155672
R2086 VTAIL.n55 VTAIL.n1 0.155672
R2087 VTAIL.n80 VTAIL.n79 0.155672
R2088 VTAIL.n80 VTAIL.n71 0.155672
R2089 VTAIL.n87 VTAIL.n71 0.155672
R2090 VTAIL.n88 VTAIL.n87 0.155672
R2091 VTAIL.n88 VTAIL.n67 0.155672
R2092 VTAIL.n96 VTAIL.n67 0.155672
R2093 VTAIL.n97 VTAIL.n96 0.155672
R2094 VTAIL.n97 VTAIL.n63 0.155672
R2095 VTAIL.n105 VTAIL.n63 0.155672
R2096 VTAIL.n106 VTAIL.n105 0.155672
R2097 VTAIL.n106 VTAIL.n59 0.155672
R2098 VTAIL.n113 VTAIL.n59 0.155672
R2099 VTAIL.n138 VTAIL.n137 0.155672
R2100 VTAIL.n138 VTAIL.n129 0.155672
R2101 VTAIL.n145 VTAIL.n129 0.155672
R2102 VTAIL.n146 VTAIL.n145 0.155672
R2103 VTAIL.n146 VTAIL.n125 0.155672
R2104 VTAIL.n154 VTAIL.n125 0.155672
R2105 VTAIL.n155 VTAIL.n154 0.155672
R2106 VTAIL.n155 VTAIL.n121 0.155672
R2107 VTAIL.n163 VTAIL.n121 0.155672
R2108 VTAIL.n164 VTAIL.n163 0.155672
R2109 VTAIL.n164 VTAIL.n117 0.155672
R2110 VTAIL.n171 VTAIL.n117 0.155672
R2111 VTAIL.n403 VTAIL.n349 0.155672
R2112 VTAIL.n396 VTAIL.n349 0.155672
R2113 VTAIL.n396 VTAIL.n395 0.155672
R2114 VTAIL.n395 VTAIL.n353 0.155672
R2115 VTAIL.n387 VTAIL.n353 0.155672
R2116 VTAIL.n387 VTAIL.n386 0.155672
R2117 VTAIL.n386 VTAIL.n357 0.155672
R2118 VTAIL.n379 VTAIL.n357 0.155672
R2119 VTAIL.n379 VTAIL.n378 0.155672
R2120 VTAIL.n378 VTAIL.n362 0.155672
R2121 VTAIL.n371 VTAIL.n362 0.155672
R2122 VTAIL.n371 VTAIL.n370 0.155672
R2123 VTAIL.n345 VTAIL.n291 0.155672
R2124 VTAIL.n338 VTAIL.n291 0.155672
R2125 VTAIL.n338 VTAIL.n337 0.155672
R2126 VTAIL.n337 VTAIL.n295 0.155672
R2127 VTAIL.n329 VTAIL.n295 0.155672
R2128 VTAIL.n329 VTAIL.n328 0.155672
R2129 VTAIL.n328 VTAIL.n299 0.155672
R2130 VTAIL.n321 VTAIL.n299 0.155672
R2131 VTAIL.n321 VTAIL.n320 0.155672
R2132 VTAIL.n320 VTAIL.n304 0.155672
R2133 VTAIL.n313 VTAIL.n304 0.155672
R2134 VTAIL.n313 VTAIL.n312 0.155672
R2135 VTAIL.n287 VTAIL.n233 0.155672
R2136 VTAIL.n280 VTAIL.n233 0.155672
R2137 VTAIL.n280 VTAIL.n279 0.155672
R2138 VTAIL.n279 VTAIL.n237 0.155672
R2139 VTAIL.n271 VTAIL.n237 0.155672
R2140 VTAIL.n271 VTAIL.n270 0.155672
R2141 VTAIL.n270 VTAIL.n241 0.155672
R2142 VTAIL.n263 VTAIL.n241 0.155672
R2143 VTAIL.n263 VTAIL.n262 0.155672
R2144 VTAIL.n262 VTAIL.n246 0.155672
R2145 VTAIL.n255 VTAIL.n246 0.155672
R2146 VTAIL.n255 VTAIL.n254 0.155672
R2147 VTAIL.n229 VTAIL.n175 0.155672
R2148 VTAIL.n222 VTAIL.n175 0.155672
R2149 VTAIL.n222 VTAIL.n221 0.155672
R2150 VTAIL.n221 VTAIL.n179 0.155672
R2151 VTAIL.n213 VTAIL.n179 0.155672
R2152 VTAIL.n213 VTAIL.n212 0.155672
R2153 VTAIL.n212 VTAIL.n183 0.155672
R2154 VTAIL.n205 VTAIL.n183 0.155672
R2155 VTAIL.n205 VTAIL.n204 0.155672
R2156 VTAIL.n204 VTAIL.n188 0.155672
R2157 VTAIL.n197 VTAIL.n188 0.155672
R2158 VTAIL.n197 VTAIL.n196 0.155672
R2159 VP.n17 VP.n16 161.3
R2160 VP.n15 VP.n1 161.3
R2161 VP.n14 VP.n13 161.3
R2162 VP.n12 VP.n2 161.3
R2163 VP.n11 VP.n10 161.3
R2164 VP.n9 VP.n3 161.3
R2165 VP.n8 VP.n7 161.3
R2166 VP.n5 VP.t0 110.731
R2167 VP.n5 VP.t3 109.599
R2168 VP.n4 VP.t2 75.7434
R2169 VP.n0 VP.t1 75.7434
R2170 VP.n6 VP.n4 73.094
R2171 VP.n18 VP.n0 73.094
R2172 VP.n6 VP.n5 50.0797
R2173 VP.n10 VP.n2 40.4106
R2174 VP.n14 VP.n2 40.4106
R2175 VP.n9 VP.n8 24.3439
R2176 VP.n10 VP.n9 24.3439
R2177 VP.n15 VP.n14 24.3439
R2178 VP.n16 VP.n15 24.3439
R2179 VP.n8 VP.n4 16.7975
R2180 VP.n16 VP.n0 16.7975
R2181 VP.n7 VP.n6 0.355081
R2182 VP.n18 VP.n17 0.355081
R2183 VP VP.n18 0.26685
R2184 VP.n7 VP.n3 0.189894
R2185 VP.n11 VP.n3 0.189894
R2186 VP.n12 VP.n11 0.189894
R2187 VP.n13 VP.n12 0.189894
R2188 VP.n13 VP.n1 0.189894
R2189 VP.n17 VP.n1 0.189894
R2190 VDD1 VDD1.n1 102.9
R2191 VDD1 VDD1.n0 60.071
R2192 VDD1.n0 VDD1.t3 1.8755
R2193 VDD1.n0 VDD1.t0 1.8755
R2194 VDD1.n1 VDD1.t1 1.8755
R2195 VDD1.n1 VDD1.t2 1.8755
C0 VDD1 VDD2 1.20298f
C1 VTAIL VP 4.49861f
C2 VN VDD2 4.39852f
C3 VDD1 VN 0.1492f
C4 VP VDD2 0.442178f
C5 VDD1 VP 4.69057f
C6 VP VN 6.47499f
C7 VTAIL VDD2 5.34179f
C8 VDD1 VTAIL 5.28249f
C9 VTAIL VN 4.484509f
C10 VDD2 B 4.092903f
C11 VDD1 B 8.386981f
C12 VTAIL B 9.624362f
C13 VN B 12.05771f
C14 VP B 10.461353f
C15 VDD1.t3 B 0.231453f
C16 VDD1.t0 B 0.231453f
C17 VDD1.n0 B 2.04338f
C18 VDD1.t1 B 0.231453f
C19 VDD1.t2 B 0.231453f
C20 VDD1.n1 B 2.76733f
C21 VP.t1 B 2.17564f
C22 VP.n0 B 0.864047f
C23 VP.n1 B 0.022593f
C24 VP.n2 B 0.018283f
C25 VP.n3 B 0.022593f
C26 VP.t2 B 2.17564f
C27 VP.n4 B 0.864047f
C28 VP.t0 B 2.47431f
C29 VP.t3 B 2.46509f
C30 VP.n5 B 2.8397f
C31 VP.n6 B 1.28794f
C32 VP.n7 B 0.03647f
C33 VP.n8 B 0.035841f
C34 VP.n9 B 0.042319f
C35 VP.n10 B 0.045143f
C36 VP.n11 B 0.022593f
C37 VP.n12 B 0.022593f
C38 VP.n13 B 0.022593f
C39 VP.n14 B 0.045143f
C40 VP.n15 B 0.042319f
C41 VP.n16 B 0.035841f
C42 VP.n17 B 0.03647f
C43 VP.n18 B 0.053131f
C44 VTAIL.n0 B 0.022089f
C45 VTAIL.n1 B 0.017384f
C46 VTAIL.n2 B 0.009341f
C47 VTAIL.n3 B 0.022079f
C48 VTAIL.n4 B 0.009891f
C49 VTAIL.n5 B 0.017384f
C50 VTAIL.n6 B 0.009341f
C51 VTAIL.n7 B 0.022079f
C52 VTAIL.n8 B 0.009891f
C53 VTAIL.n9 B 0.017384f
C54 VTAIL.n10 B 0.009341f
C55 VTAIL.n11 B 0.022079f
C56 VTAIL.n12 B 0.009891f
C57 VTAIL.n13 B 0.017384f
C58 VTAIL.n14 B 0.009341f
C59 VTAIL.n15 B 0.022079f
C60 VTAIL.n16 B 0.009891f
C61 VTAIL.n17 B 0.115724f
C62 VTAIL.t2 B 0.037156f
C63 VTAIL.n18 B 0.016559f
C64 VTAIL.n19 B 0.015608f
C65 VTAIL.n20 B 0.009341f
C66 VTAIL.n21 B 0.765634f
C67 VTAIL.n22 B 0.017384f
C68 VTAIL.n23 B 0.009341f
C69 VTAIL.n24 B 0.009891f
C70 VTAIL.n25 B 0.022079f
C71 VTAIL.n26 B 0.022079f
C72 VTAIL.n27 B 0.009891f
C73 VTAIL.n28 B 0.009341f
C74 VTAIL.n29 B 0.017384f
C75 VTAIL.n30 B 0.017384f
C76 VTAIL.n31 B 0.009341f
C77 VTAIL.n32 B 0.009891f
C78 VTAIL.n33 B 0.022079f
C79 VTAIL.n34 B 0.022079f
C80 VTAIL.n35 B 0.022079f
C81 VTAIL.n36 B 0.009891f
C82 VTAIL.n37 B 0.009341f
C83 VTAIL.n38 B 0.017384f
C84 VTAIL.n39 B 0.017384f
C85 VTAIL.n40 B 0.009341f
C86 VTAIL.n41 B 0.009616f
C87 VTAIL.n42 B 0.009616f
C88 VTAIL.n43 B 0.022079f
C89 VTAIL.n44 B 0.022079f
C90 VTAIL.n45 B 0.009891f
C91 VTAIL.n46 B 0.009341f
C92 VTAIL.n47 B 0.017384f
C93 VTAIL.n48 B 0.017384f
C94 VTAIL.n49 B 0.009341f
C95 VTAIL.n50 B 0.009891f
C96 VTAIL.n51 B 0.022079f
C97 VTAIL.n52 B 0.04365f
C98 VTAIL.n53 B 0.009891f
C99 VTAIL.n54 B 0.009341f
C100 VTAIL.n55 B 0.037332f
C101 VTAIL.n56 B 0.023907f
C102 VTAIL.n57 B 0.131909f
C103 VTAIL.n58 B 0.022089f
C104 VTAIL.n59 B 0.017384f
C105 VTAIL.n60 B 0.009341f
C106 VTAIL.n61 B 0.022079f
C107 VTAIL.n62 B 0.009891f
C108 VTAIL.n63 B 0.017384f
C109 VTAIL.n64 B 0.009341f
C110 VTAIL.n65 B 0.022079f
C111 VTAIL.n66 B 0.009891f
C112 VTAIL.n67 B 0.017384f
C113 VTAIL.n68 B 0.009341f
C114 VTAIL.n69 B 0.022079f
C115 VTAIL.n70 B 0.009891f
C116 VTAIL.n71 B 0.017384f
C117 VTAIL.n72 B 0.009341f
C118 VTAIL.n73 B 0.022079f
C119 VTAIL.n74 B 0.009891f
C120 VTAIL.n75 B 0.115724f
C121 VTAIL.t6 B 0.037156f
C122 VTAIL.n76 B 0.016559f
C123 VTAIL.n77 B 0.015608f
C124 VTAIL.n78 B 0.009341f
C125 VTAIL.n79 B 0.765634f
C126 VTAIL.n80 B 0.017384f
C127 VTAIL.n81 B 0.009341f
C128 VTAIL.n82 B 0.009891f
C129 VTAIL.n83 B 0.022079f
C130 VTAIL.n84 B 0.022079f
C131 VTAIL.n85 B 0.009891f
C132 VTAIL.n86 B 0.009341f
C133 VTAIL.n87 B 0.017384f
C134 VTAIL.n88 B 0.017384f
C135 VTAIL.n89 B 0.009341f
C136 VTAIL.n90 B 0.009891f
C137 VTAIL.n91 B 0.022079f
C138 VTAIL.n92 B 0.022079f
C139 VTAIL.n93 B 0.022079f
C140 VTAIL.n94 B 0.009891f
C141 VTAIL.n95 B 0.009341f
C142 VTAIL.n96 B 0.017384f
C143 VTAIL.n97 B 0.017384f
C144 VTAIL.n98 B 0.009341f
C145 VTAIL.n99 B 0.009616f
C146 VTAIL.n100 B 0.009616f
C147 VTAIL.n101 B 0.022079f
C148 VTAIL.n102 B 0.022079f
C149 VTAIL.n103 B 0.009891f
C150 VTAIL.n104 B 0.009341f
C151 VTAIL.n105 B 0.017384f
C152 VTAIL.n106 B 0.017384f
C153 VTAIL.n107 B 0.009341f
C154 VTAIL.n108 B 0.009891f
C155 VTAIL.n109 B 0.022079f
C156 VTAIL.n110 B 0.04365f
C157 VTAIL.n111 B 0.009891f
C158 VTAIL.n112 B 0.009341f
C159 VTAIL.n113 B 0.037332f
C160 VTAIL.n114 B 0.023907f
C161 VTAIL.n115 B 0.217741f
C162 VTAIL.n116 B 0.022089f
C163 VTAIL.n117 B 0.017384f
C164 VTAIL.n118 B 0.009341f
C165 VTAIL.n119 B 0.022079f
C166 VTAIL.n120 B 0.009891f
C167 VTAIL.n121 B 0.017384f
C168 VTAIL.n122 B 0.009341f
C169 VTAIL.n123 B 0.022079f
C170 VTAIL.n124 B 0.009891f
C171 VTAIL.n125 B 0.017384f
C172 VTAIL.n126 B 0.009341f
C173 VTAIL.n127 B 0.022079f
C174 VTAIL.n128 B 0.009891f
C175 VTAIL.n129 B 0.017384f
C176 VTAIL.n130 B 0.009341f
C177 VTAIL.n131 B 0.022079f
C178 VTAIL.n132 B 0.009891f
C179 VTAIL.n133 B 0.115724f
C180 VTAIL.t0 B 0.037156f
C181 VTAIL.n134 B 0.016559f
C182 VTAIL.n135 B 0.015608f
C183 VTAIL.n136 B 0.009341f
C184 VTAIL.n137 B 0.765634f
C185 VTAIL.n138 B 0.017384f
C186 VTAIL.n139 B 0.009341f
C187 VTAIL.n140 B 0.009891f
C188 VTAIL.n141 B 0.022079f
C189 VTAIL.n142 B 0.022079f
C190 VTAIL.n143 B 0.009891f
C191 VTAIL.n144 B 0.009341f
C192 VTAIL.n145 B 0.017384f
C193 VTAIL.n146 B 0.017384f
C194 VTAIL.n147 B 0.009341f
C195 VTAIL.n148 B 0.009891f
C196 VTAIL.n149 B 0.022079f
C197 VTAIL.n150 B 0.022079f
C198 VTAIL.n151 B 0.022079f
C199 VTAIL.n152 B 0.009891f
C200 VTAIL.n153 B 0.009341f
C201 VTAIL.n154 B 0.017384f
C202 VTAIL.n155 B 0.017384f
C203 VTAIL.n156 B 0.009341f
C204 VTAIL.n157 B 0.009616f
C205 VTAIL.n158 B 0.009616f
C206 VTAIL.n159 B 0.022079f
C207 VTAIL.n160 B 0.022079f
C208 VTAIL.n161 B 0.009891f
C209 VTAIL.n162 B 0.009341f
C210 VTAIL.n163 B 0.017384f
C211 VTAIL.n164 B 0.017384f
C212 VTAIL.n165 B 0.009341f
C213 VTAIL.n166 B 0.009891f
C214 VTAIL.n167 B 0.022079f
C215 VTAIL.n168 B 0.04365f
C216 VTAIL.n169 B 0.009891f
C217 VTAIL.n170 B 0.009341f
C218 VTAIL.n171 B 0.037332f
C219 VTAIL.n172 B 0.023907f
C220 VTAIL.n173 B 1.11566f
C221 VTAIL.n174 B 0.022089f
C222 VTAIL.n175 B 0.017384f
C223 VTAIL.n176 B 0.009341f
C224 VTAIL.n177 B 0.022079f
C225 VTAIL.n178 B 0.009891f
C226 VTAIL.n179 B 0.017384f
C227 VTAIL.n180 B 0.009341f
C228 VTAIL.n181 B 0.022079f
C229 VTAIL.n182 B 0.009891f
C230 VTAIL.n183 B 0.017384f
C231 VTAIL.n184 B 0.009341f
C232 VTAIL.n185 B 0.022079f
C233 VTAIL.n186 B 0.022079f
C234 VTAIL.n187 B 0.009891f
C235 VTAIL.n188 B 0.017384f
C236 VTAIL.n189 B 0.009341f
C237 VTAIL.n190 B 0.022079f
C238 VTAIL.n191 B 0.009891f
C239 VTAIL.n192 B 0.115724f
C240 VTAIL.t5 B 0.037156f
C241 VTAIL.n193 B 0.016559f
C242 VTAIL.n194 B 0.015608f
C243 VTAIL.n195 B 0.009341f
C244 VTAIL.n196 B 0.765634f
C245 VTAIL.n197 B 0.017384f
C246 VTAIL.n198 B 0.009341f
C247 VTAIL.n199 B 0.009891f
C248 VTAIL.n200 B 0.022079f
C249 VTAIL.n201 B 0.022079f
C250 VTAIL.n202 B 0.009891f
C251 VTAIL.n203 B 0.009341f
C252 VTAIL.n204 B 0.017384f
C253 VTAIL.n205 B 0.017384f
C254 VTAIL.n206 B 0.009341f
C255 VTAIL.n207 B 0.009891f
C256 VTAIL.n208 B 0.022079f
C257 VTAIL.n209 B 0.022079f
C258 VTAIL.n210 B 0.009891f
C259 VTAIL.n211 B 0.009341f
C260 VTAIL.n212 B 0.017384f
C261 VTAIL.n213 B 0.017384f
C262 VTAIL.n214 B 0.009341f
C263 VTAIL.n215 B 0.009616f
C264 VTAIL.n216 B 0.009616f
C265 VTAIL.n217 B 0.022079f
C266 VTAIL.n218 B 0.022079f
C267 VTAIL.n219 B 0.009891f
C268 VTAIL.n220 B 0.009341f
C269 VTAIL.n221 B 0.017384f
C270 VTAIL.n222 B 0.017384f
C271 VTAIL.n223 B 0.009341f
C272 VTAIL.n224 B 0.009891f
C273 VTAIL.n225 B 0.022079f
C274 VTAIL.n226 B 0.04365f
C275 VTAIL.n227 B 0.009891f
C276 VTAIL.n228 B 0.009341f
C277 VTAIL.n229 B 0.037332f
C278 VTAIL.n230 B 0.023907f
C279 VTAIL.n231 B 1.11566f
C280 VTAIL.n232 B 0.022089f
C281 VTAIL.n233 B 0.017384f
C282 VTAIL.n234 B 0.009341f
C283 VTAIL.n235 B 0.022079f
C284 VTAIL.n236 B 0.009891f
C285 VTAIL.n237 B 0.017384f
C286 VTAIL.n238 B 0.009341f
C287 VTAIL.n239 B 0.022079f
C288 VTAIL.n240 B 0.009891f
C289 VTAIL.n241 B 0.017384f
C290 VTAIL.n242 B 0.009341f
C291 VTAIL.n243 B 0.022079f
C292 VTAIL.n244 B 0.022079f
C293 VTAIL.n245 B 0.009891f
C294 VTAIL.n246 B 0.017384f
C295 VTAIL.n247 B 0.009341f
C296 VTAIL.n248 B 0.022079f
C297 VTAIL.n249 B 0.009891f
C298 VTAIL.n250 B 0.115724f
C299 VTAIL.t4 B 0.037156f
C300 VTAIL.n251 B 0.016559f
C301 VTAIL.n252 B 0.015608f
C302 VTAIL.n253 B 0.009341f
C303 VTAIL.n254 B 0.765634f
C304 VTAIL.n255 B 0.017384f
C305 VTAIL.n256 B 0.009341f
C306 VTAIL.n257 B 0.009891f
C307 VTAIL.n258 B 0.022079f
C308 VTAIL.n259 B 0.022079f
C309 VTAIL.n260 B 0.009891f
C310 VTAIL.n261 B 0.009341f
C311 VTAIL.n262 B 0.017384f
C312 VTAIL.n263 B 0.017384f
C313 VTAIL.n264 B 0.009341f
C314 VTAIL.n265 B 0.009891f
C315 VTAIL.n266 B 0.022079f
C316 VTAIL.n267 B 0.022079f
C317 VTAIL.n268 B 0.009891f
C318 VTAIL.n269 B 0.009341f
C319 VTAIL.n270 B 0.017384f
C320 VTAIL.n271 B 0.017384f
C321 VTAIL.n272 B 0.009341f
C322 VTAIL.n273 B 0.009616f
C323 VTAIL.n274 B 0.009616f
C324 VTAIL.n275 B 0.022079f
C325 VTAIL.n276 B 0.022079f
C326 VTAIL.n277 B 0.009891f
C327 VTAIL.n278 B 0.009341f
C328 VTAIL.n279 B 0.017384f
C329 VTAIL.n280 B 0.017384f
C330 VTAIL.n281 B 0.009341f
C331 VTAIL.n282 B 0.009891f
C332 VTAIL.n283 B 0.022079f
C333 VTAIL.n284 B 0.04365f
C334 VTAIL.n285 B 0.009891f
C335 VTAIL.n286 B 0.009341f
C336 VTAIL.n287 B 0.037332f
C337 VTAIL.n288 B 0.023907f
C338 VTAIL.n289 B 0.217741f
C339 VTAIL.n290 B 0.022089f
C340 VTAIL.n291 B 0.017384f
C341 VTAIL.n292 B 0.009341f
C342 VTAIL.n293 B 0.022079f
C343 VTAIL.n294 B 0.009891f
C344 VTAIL.n295 B 0.017384f
C345 VTAIL.n296 B 0.009341f
C346 VTAIL.n297 B 0.022079f
C347 VTAIL.n298 B 0.009891f
C348 VTAIL.n299 B 0.017384f
C349 VTAIL.n300 B 0.009341f
C350 VTAIL.n301 B 0.022079f
C351 VTAIL.n302 B 0.022079f
C352 VTAIL.n303 B 0.009891f
C353 VTAIL.n304 B 0.017384f
C354 VTAIL.n305 B 0.009341f
C355 VTAIL.n306 B 0.022079f
C356 VTAIL.n307 B 0.009891f
C357 VTAIL.n308 B 0.115724f
C358 VTAIL.t7 B 0.037156f
C359 VTAIL.n309 B 0.016559f
C360 VTAIL.n310 B 0.015608f
C361 VTAIL.n311 B 0.009341f
C362 VTAIL.n312 B 0.765634f
C363 VTAIL.n313 B 0.017384f
C364 VTAIL.n314 B 0.009341f
C365 VTAIL.n315 B 0.009891f
C366 VTAIL.n316 B 0.022079f
C367 VTAIL.n317 B 0.022079f
C368 VTAIL.n318 B 0.009891f
C369 VTAIL.n319 B 0.009341f
C370 VTAIL.n320 B 0.017384f
C371 VTAIL.n321 B 0.017384f
C372 VTAIL.n322 B 0.009341f
C373 VTAIL.n323 B 0.009891f
C374 VTAIL.n324 B 0.022079f
C375 VTAIL.n325 B 0.022079f
C376 VTAIL.n326 B 0.009891f
C377 VTAIL.n327 B 0.009341f
C378 VTAIL.n328 B 0.017384f
C379 VTAIL.n329 B 0.017384f
C380 VTAIL.n330 B 0.009341f
C381 VTAIL.n331 B 0.009616f
C382 VTAIL.n332 B 0.009616f
C383 VTAIL.n333 B 0.022079f
C384 VTAIL.n334 B 0.022079f
C385 VTAIL.n335 B 0.009891f
C386 VTAIL.n336 B 0.009341f
C387 VTAIL.n337 B 0.017384f
C388 VTAIL.n338 B 0.017384f
C389 VTAIL.n339 B 0.009341f
C390 VTAIL.n340 B 0.009891f
C391 VTAIL.n341 B 0.022079f
C392 VTAIL.n342 B 0.04365f
C393 VTAIL.n343 B 0.009891f
C394 VTAIL.n344 B 0.009341f
C395 VTAIL.n345 B 0.037332f
C396 VTAIL.n346 B 0.023907f
C397 VTAIL.n347 B 0.217741f
C398 VTAIL.n348 B 0.022089f
C399 VTAIL.n349 B 0.017384f
C400 VTAIL.n350 B 0.009341f
C401 VTAIL.n351 B 0.022079f
C402 VTAIL.n352 B 0.009891f
C403 VTAIL.n353 B 0.017384f
C404 VTAIL.n354 B 0.009341f
C405 VTAIL.n355 B 0.022079f
C406 VTAIL.n356 B 0.009891f
C407 VTAIL.n357 B 0.017384f
C408 VTAIL.n358 B 0.009341f
C409 VTAIL.n359 B 0.022079f
C410 VTAIL.n360 B 0.022079f
C411 VTAIL.n361 B 0.009891f
C412 VTAIL.n362 B 0.017384f
C413 VTAIL.n363 B 0.009341f
C414 VTAIL.n364 B 0.022079f
C415 VTAIL.n365 B 0.009891f
C416 VTAIL.n366 B 0.115724f
C417 VTAIL.t1 B 0.037156f
C418 VTAIL.n367 B 0.016559f
C419 VTAIL.n368 B 0.015608f
C420 VTAIL.n369 B 0.009341f
C421 VTAIL.n370 B 0.765634f
C422 VTAIL.n371 B 0.017384f
C423 VTAIL.n372 B 0.009341f
C424 VTAIL.n373 B 0.009891f
C425 VTAIL.n374 B 0.022079f
C426 VTAIL.n375 B 0.022079f
C427 VTAIL.n376 B 0.009891f
C428 VTAIL.n377 B 0.009341f
C429 VTAIL.n378 B 0.017384f
C430 VTAIL.n379 B 0.017384f
C431 VTAIL.n380 B 0.009341f
C432 VTAIL.n381 B 0.009891f
C433 VTAIL.n382 B 0.022079f
C434 VTAIL.n383 B 0.022079f
C435 VTAIL.n384 B 0.009891f
C436 VTAIL.n385 B 0.009341f
C437 VTAIL.n386 B 0.017384f
C438 VTAIL.n387 B 0.017384f
C439 VTAIL.n388 B 0.009341f
C440 VTAIL.n389 B 0.009616f
C441 VTAIL.n390 B 0.009616f
C442 VTAIL.n391 B 0.022079f
C443 VTAIL.n392 B 0.022079f
C444 VTAIL.n393 B 0.009891f
C445 VTAIL.n394 B 0.009341f
C446 VTAIL.n395 B 0.017384f
C447 VTAIL.n396 B 0.017384f
C448 VTAIL.n397 B 0.009341f
C449 VTAIL.n398 B 0.009891f
C450 VTAIL.n399 B 0.022079f
C451 VTAIL.n400 B 0.04365f
C452 VTAIL.n401 B 0.009891f
C453 VTAIL.n402 B 0.009341f
C454 VTAIL.n403 B 0.037332f
C455 VTAIL.n404 B 0.023907f
C456 VTAIL.n405 B 1.11566f
C457 VTAIL.n406 B 0.022089f
C458 VTAIL.n407 B 0.017384f
C459 VTAIL.n408 B 0.009341f
C460 VTAIL.n409 B 0.022079f
C461 VTAIL.n410 B 0.009891f
C462 VTAIL.n411 B 0.017384f
C463 VTAIL.n412 B 0.009341f
C464 VTAIL.n413 B 0.022079f
C465 VTAIL.n414 B 0.009891f
C466 VTAIL.n415 B 0.017384f
C467 VTAIL.n416 B 0.009341f
C468 VTAIL.n417 B 0.022079f
C469 VTAIL.n418 B 0.009891f
C470 VTAIL.n419 B 0.017384f
C471 VTAIL.n420 B 0.009341f
C472 VTAIL.n421 B 0.022079f
C473 VTAIL.n422 B 0.009891f
C474 VTAIL.n423 B 0.115724f
C475 VTAIL.t3 B 0.037156f
C476 VTAIL.n424 B 0.016559f
C477 VTAIL.n425 B 0.015608f
C478 VTAIL.n426 B 0.009341f
C479 VTAIL.n427 B 0.765634f
C480 VTAIL.n428 B 0.017384f
C481 VTAIL.n429 B 0.009341f
C482 VTAIL.n430 B 0.009891f
C483 VTAIL.n431 B 0.022079f
C484 VTAIL.n432 B 0.022079f
C485 VTAIL.n433 B 0.009891f
C486 VTAIL.n434 B 0.009341f
C487 VTAIL.n435 B 0.017384f
C488 VTAIL.n436 B 0.017384f
C489 VTAIL.n437 B 0.009341f
C490 VTAIL.n438 B 0.009891f
C491 VTAIL.n439 B 0.022079f
C492 VTAIL.n440 B 0.022079f
C493 VTAIL.n441 B 0.022079f
C494 VTAIL.n442 B 0.009891f
C495 VTAIL.n443 B 0.009341f
C496 VTAIL.n444 B 0.017384f
C497 VTAIL.n445 B 0.017384f
C498 VTAIL.n446 B 0.009341f
C499 VTAIL.n447 B 0.009616f
C500 VTAIL.n448 B 0.009616f
C501 VTAIL.n449 B 0.022079f
C502 VTAIL.n450 B 0.022079f
C503 VTAIL.n451 B 0.009891f
C504 VTAIL.n452 B 0.009341f
C505 VTAIL.n453 B 0.017384f
C506 VTAIL.n454 B 0.017384f
C507 VTAIL.n455 B 0.009341f
C508 VTAIL.n456 B 0.009891f
C509 VTAIL.n457 B 0.022079f
C510 VTAIL.n458 B 0.04365f
C511 VTAIL.n459 B 0.009891f
C512 VTAIL.n460 B 0.009341f
C513 VTAIL.n461 B 0.037332f
C514 VTAIL.n462 B 0.023907f
C515 VTAIL.n463 B 1.02331f
C516 VDD2.t3 B 0.226834f
C517 VDD2.t0 B 0.226834f
C518 VDD2.n0 B 2.68472f
C519 VDD2.t1 B 0.226834f
C520 VDD2.t2 B 0.226834f
C521 VDD2.n1 B 2.00209f
C522 VDD2.n2 B 3.82139f
C523 VN.t2 B 2.41311f
C524 VN.t3 B 2.42213f
C525 VN.n0 B 1.44852f
C526 VN.t0 B 2.41311f
C527 VN.t1 B 2.42213f
C528 VN.n1 B 2.7888f
.ends

