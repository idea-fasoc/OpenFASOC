* NGSPICE file created from diff_pair_sample_0468.ext - technology: sky130A

.subckt diff_pair_sample_0468 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t16 VP.t0 VDD1.t1 B.t5 sky130_fd_pr__nfet_01v8 ad=1.7325 pd=10.83 as=1.7325 ps=10.83 w=10.5 l=0.61
X1 VTAIL.t15 VP.t1 VDD1.t0 B.t4 sky130_fd_pr__nfet_01v8 ad=1.7325 pd=10.83 as=1.7325 ps=10.83 w=10.5 l=0.61
X2 B.t20 B.t18 B.t19 B.t12 sky130_fd_pr__nfet_01v8 ad=4.095 pd=21.78 as=0 ps=0 w=10.5 l=0.61
X3 VDD1.t5 VP.t2 VTAIL.t14 B.t2 sky130_fd_pr__nfet_01v8 ad=4.095 pd=21.78 as=1.7325 ps=10.83 w=10.5 l=0.61
X4 B.t17 B.t15 B.t16 B.t8 sky130_fd_pr__nfet_01v8 ad=4.095 pd=21.78 as=0 ps=0 w=10.5 l=0.61
X5 VTAIL.t5 VN.t0 VDD2.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=1.7325 pd=10.83 as=1.7325 ps=10.83 w=10.5 l=0.61
X6 VDD1.t3 VP.t3 VTAIL.t13 B.t23 sky130_fd_pr__nfet_01v8 ad=1.7325 pd=10.83 as=4.095 ps=21.78 w=10.5 l=0.61
X7 VDD2.t8 VN.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.7325 pd=10.83 as=1.7325 ps=10.83 w=10.5 l=0.61
X8 VDD1.t8 VP.t4 VTAIL.t12 B.t6 sky130_fd_pr__nfet_01v8 ad=4.095 pd=21.78 as=1.7325 ps=10.83 w=10.5 l=0.61
X9 VTAIL.t11 VP.t5 VDD1.t7 B.t22 sky130_fd_pr__nfet_01v8 ad=1.7325 pd=10.83 as=1.7325 ps=10.83 w=10.5 l=0.61
X10 B.t14 B.t11 B.t13 B.t12 sky130_fd_pr__nfet_01v8 ad=4.095 pd=21.78 as=0 ps=0 w=10.5 l=0.61
X11 VDD1.t6 VP.t6 VTAIL.t10 B.t1 sky130_fd_pr__nfet_01v8 ad=1.7325 pd=10.83 as=1.7325 ps=10.83 w=10.5 l=0.61
X12 VTAIL.t9 VP.t7 VDD1.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=1.7325 pd=10.83 as=1.7325 ps=10.83 w=10.5 l=0.61
X13 VDD2.t7 VN.t2 VTAIL.t18 B.t21 sky130_fd_pr__nfet_01v8 ad=1.7325 pd=10.83 as=1.7325 ps=10.83 w=10.5 l=0.61
X14 VTAIL.t4 VN.t3 VDD2.t6 B.t4 sky130_fd_pr__nfet_01v8 ad=1.7325 pd=10.83 as=1.7325 ps=10.83 w=10.5 l=0.61
X15 VTAIL.t17 VN.t4 VDD2.t5 B.t22 sky130_fd_pr__nfet_01v8 ad=1.7325 pd=10.83 as=1.7325 ps=10.83 w=10.5 l=0.61
X16 VDD2.t4 VN.t5 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=4.095 pd=21.78 as=1.7325 ps=10.83 w=10.5 l=0.61
X17 VDD2.t3 VN.t6 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.7325 pd=10.83 as=4.095 ps=21.78 w=10.5 l=0.61
X18 VDD1.t9 VP.t8 VTAIL.t8 B.t21 sky130_fd_pr__nfet_01v8 ad=1.7325 pd=10.83 as=1.7325 ps=10.83 w=10.5 l=0.61
X19 VDD2.t2 VN.t7 VTAIL.t19 B.t23 sky130_fd_pr__nfet_01v8 ad=1.7325 pd=10.83 as=4.095 ps=21.78 w=10.5 l=0.61
X20 B.t10 B.t7 B.t9 B.t8 sky130_fd_pr__nfet_01v8 ad=4.095 pd=21.78 as=0 ps=0 w=10.5 l=0.61
X21 VDD1.t4 VP.t9 VTAIL.t7 B.t0 sky130_fd_pr__nfet_01v8 ad=1.7325 pd=10.83 as=4.095 ps=21.78 w=10.5 l=0.61
X22 VTAIL.t3 VN.t8 VDD2.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=1.7325 pd=10.83 as=1.7325 ps=10.83 w=10.5 l=0.61
X23 VDD2.t0 VN.t9 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=4.095 pd=21.78 as=1.7325 ps=10.83 w=10.5 l=0.61
R0 VP.n6 VP.t2 505.904
R1 VP.n14 VP.t4 479.235
R2 VP.n16 VP.t1 479.235
R3 VP.n1 VP.t6 479.235
R4 VP.n20 VP.t7 479.235
R5 VP.n22 VP.t9 479.235
R6 VP.n11 VP.t3 479.235
R7 VP.n9 VP.t0 479.235
R8 VP.n8 VP.t8 479.235
R9 VP.n7 VP.t5 479.235
R10 VP.n23 VP.n22 161.3
R11 VP.n9 VP.n4 161.3
R12 VP.n10 VP.n3 161.3
R13 VP.n12 VP.n11 161.3
R14 VP.n21 VP.n0 161.3
R15 VP.n20 VP.n19 161.3
R16 VP.n17 VP.n16 161.3
R17 VP.n15 VP.n2 161.3
R18 VP.n14 VP.n13 161.3
R19 VP.n8 VP.n5 80.6037
R20 VP.n18 VP.n1 80.6037
R21 VP.n16 VP.n1 48.2005
R22 VP.n20 VP.n1 48.2005
R23 VP.n9 VP.n8 48.2005
R24 VP.n8 VP.n7 48.2005
R25 VP.n15 VP.n14 47.4702
R26 VP.n22 VP.n21 47.4702
R27 VP.n11 VP.n10 47.4702
R28 VP.n6 VP.n5 45.2144
R29 VP.n13 VP.n12 41.1899
R30 VP.n7 VP.n6 13.6377
R31 VP.n16 VP.n15 0.730803
R32 VP.n21 VP.n20 0.730803
R33 VP.n10 VP.n9 0.730803
R34 VP.n5 VP.n4 0.285035
R35 VP.n18 VP.n17 0.285035
R36 VP.n19 VP.n18 0.285035
R37 VP.n4 VP.n3 0.189894
R38 VP.n12 VP.n3 0.189894
R39 VP.n13 VP.n2 0.189894
R40 VP.n17 VP.n2 0.189894
R41 VP.n19 VP.n0 0.189894
R42 VP.n23 VP.n0 0.189894
R43 VP VP.n23 0.0516364
R44 VDD1.n1 VDD1.t5 68.67
R45 VDD1.n3 VDD1.t8 68.6697
R46 VDD1.n5 VDD1.n4 66.5261
R47 VDD1.n1 VDD1.n0 65.9739
R48 VDD1.n7 VDD1.n6 65.9737
R49 VDD1.n3 VDD1.n2 65.9737
R50 VDD1.n7 VDD1.n5 37.6043
R51 VDD1.n6 VDD1.t1 1.88621
R52 VDD1.n6 VDD1.t3 1.88621
R53 VDD1.n0 VDD1.t7 1.88621
R54 VDD1.n0 VDD1.t9 1.88621
R55 VDD1.n4 VDD1.t2 1.88621
R56 VDD1.n4 VDD1.t4 1.88621
R57 VDD1.n2 VDD1.t0 1.88621
R58 VDD1.n2 VDD1.t6 1.88621
R59 VDD1 VDD1.n7 0.550069
R60 VDD1 VDD1.n1 0.261276
R61 VDD1.n5 VDD1.n3 0.14774
R62 VTAIL.n11 VTAIL.t0 51.1808
R63 VTAIL.n17 VTAIL.t19 51.1806
R64 VTAIL.n2 VTAIL.t7 51.1806
R65 VTAIL.n16 VTAIL.t13 51.1806
R66 VTAIL.n15 VTAIL.n14 49.2951
R67 VTAIL.n13 VTAIL.n12 49.2951
R68 VTAIL.n10 VTAIL.n9 49.2951
R69 VTAIL.n8 VTAIL.n7 49.2951
R70 VTAIL.n19 VTAIL.n18 49.2949
R71 VTAIL.n1 VTAIL.n0 49.2949
R72 VTAIL.n4 VTAIL.n3 49.2949
R73 VTAIL.n6 VTAIL.n5 49.2949
R74 VTAIL.n8 VTAIL.n6 23.0393
R75 VTAIL.n17 VTAIL.n16 22.2289
R76 VTAIL.n18 VTAIL.t18 1.88621
R77 VTAIL.n18 VTAIL.t5 1.88621
R78 VTAIL.n0 VTAIL.t2 1.88621
R79 VTAIL.n0 VTAIL.t17 1.88621
R80 VTAIL.n3 VTAIL.t10 1.88621
R81 VTAIL.n3 VTAIL.t9 1.88621
R82 VTAIL.n5 VTAIL.t12 1.88621
R83 VTAIL.n5 VTAIL.t15 1.88621
R84 VTAIL.n14 VTAIL.t8 1.88621
R85 VTAIL.n14 VTAIL.t16 1.88621
R86 VTAIL.n12 VTAIL.t14 1.88621
R87 VTAIL.n12 VTAIL.t11 1.88621
R88 VTAIL.n9 VTAIL.t1 1.88621
R89 VTAIL.n9 VTAIL.t3 1.88621
R90 VTAIL.n7 VTAIL.t6 1.88621
R91 VTAIL.n7 VTAIL.t4 1.88621
R92 VTAIL.n13 VTAIL.n11 0.8755
R93 VTAIL.n2 VTAIL.n1 0.8755
R94 VTAIL.n10 VTAIL.n8 0.810845
R95 VTAIL.n11 VTAIL.n10 0.810845
R96 VTAIL.n15 VTAIL.n13 0.810845
R97 VTAIL.n16 VTAIL.n15 0.810845
R98 VTAIL.n6 VTAIL.n4 0.810845
R99 VTAIL.n4 VTAIL.n2 0.810845
R100 VTAIL.n19 VTAIL.n17 0.810845
R101 VTAIL VTAIL.n1 0.666448
R102 VTAIL VTAIL.n19 0.144897
R103 B.n93 B.t18 619.072
R104 B.n91 B.t11 619.072
R105 B.n325 B.t15 619.072
R106 B.n331 B.t7 619.072
R107 B.n627 B.n626 585
R108 B.n259 B.n90 585
R109 B.n258 B.n257 585
R110 B.n256 B.n255 585
R111 B.n254 B.n253 585
R112 B.n252 B.n251 585
R113 B.n250 B.n249 585
R114 B.n248 B.n247 585
R115 B.n246 B.n245 585
R116 B.n244 B.n243 585
R117 B.n242 B.n241 585
R118 B.n240 B.n239 585
R119 B.n238 B.n237 585
R120 B.n236 B.n235 585
R121 B.n234 B.n233 585
R122 B.n232 B.n231 585
R123 B.n230 B.n229 585
R124 B.n228 B.n227 585
R125 B.n226 B.n225 585
R126 B.n224 B.n223 585
R127 B.n222 B.n221 585
R128 B.n220 B.n219 585
R129 B.n218 B.n217 585
R130 B.n216 B.n215 585
R131 B.n214 B.n213 585
R132 B.n212 B.n211 585
R133 B.n210 B.n209 585
R134 B.n208 B.n207 585
R135 B.n206 B.n205 585
R136 B.n204 B.n203 585
R137 B.n202 B.n201 585
R138 B.n200 B.n199 585
R139 B.n198 B.n197 585
R140 B.n196 B.n195 585
R141 B.n194 B.n193 585
R142 B.n192 B.n191 585
R143 B.n190 B.n189 585
R144 B.n187 B.n186 585
R145 B.n185 B.n184 585
R146 B.n183 B.n182 585
R147 B.n181 B.n180 585
R148 B.n179 B.n178 585
R149 B.n177 B.n176 585
R150 B.n175 B.n174 585
R151 B.n173 B.n172 585
R152 B.n171 B.n170 585
R153 B.n169 B.n168 585
R154 B.n166 B.n165 585
R155 B.n164 B.n163 585
R156 B.n162 B.n161 585
R157 B.n160 B.n159 585
R158 B.n158 B.n157 585
R159 B.n156 B.n155 585
R160 B.n154 B.n153 585
R161 B.n152 B.n151 585
R162 B.n150 B.n149 585
R163 B.n148 B.n147 585
R164 B.n146 B.n145 585
R165 B.n144 B.n143 585
R166 B.n142 B.n141 585
R167 B.n140 B.n139 585
R168 B.n138 B.n137 585
R169 B.n136 B.n135 585
R170 B.n134 B.n133 585
R171 B.n132 B.n131 585
R172 B.n130 B.n129 585
R173 B.n128 B.n127 585
R174 B.n126 B.n125 585
R175 B.n124 B.n123 585
R176 B.n122 B.n121 585
R177 B.n120 B.n119 585
R178 B.n118 B.n117 585
R179 B.n116 B.n115 585
R180 B.n114 B.n113 585
R181 B.n112 B.n111 585
R182 B.n110 B.n109 585
R183 B.n108 B.n107 585
R184 B.n106 B.n105 585
R185 B.n104 B.n103 585
R186 B.n102 B.n101 585
R187 B.n100 B.n99 585
R188 B.n98 B.n97 585
R189 B.n96 B.n95 585
R190 B.n47 B.n46 585
R191 B.n625 B.n48 585
R192 B.n630 B.n48 585
R193 B.n624 B.n623 585
R194 B.n623 B.n44 585
R195 B.n622 B.n43 585
R196 B.n636 B.n43 585
R197 B.n621 B.n42 585
R198 B.n637 B.n42 585
R199 B.n620 B.n41 585
R200 B.n638 B.n41 585
R201 B.n619 B.n618 585
R202 B.n618 B.n37 585
R203 B.n617 B.n36 585
R204 B.n644 B.n36 585
R205 B.n616 B.n35 585
R206 B.n645 B.n35 585
R207 B.n615 B.n34 585
R208 B.n646 B.n34 585
R209 B.n614 B.n613 585
R210 B.n613 B.n30 585
R211 B.n612 B.n29 585
R212 B.n652 B.n29 585
R213 B.n611 B.n28 585
R214 B.n653 B.n28 585
R215 B.n610 B.n27 585
R216 B.n654 B.n27 585
R217 B.n609 B.n608 585
R218 B.n608 B.n26 585
R219 B.n607 B.n22 585
R220 B.n660 B.n22 585
R221 B.n606 B.n21 585
R222 B.n661 B.n21 585
R223 B.n605 B.n20 585
R224 B.n662 B.n20 585
R225 B.n604 B.n603 585
R226 B.n603 B.n16 585
R227 B.n602 B.n15 585
R228 B.n668 B.n15 585
R229 B.n601 B.n14 585
R230 B.n669 B.n14 585
R231 B.n600 B.n13 585
R232 B.n670 B.n13 585
R233 B.n599 B.n598 585
R234 B.n598 B.n12 585
R235 B.n597 B.n596 585
R236 B.n597 B.n8 585
R237 B.n595 B.n7 585
R238 B.n677 B.n7 585
R239 B.n594 B.n6 585
R240 B.n678 B.n6 585
R241 B.n593 B.n5 585
R242 B.n679 B.n5 585
R243 B.n592 B.n591 585
R244 B.n591 B.n4 585
R245 B.n590 B.n260 585
R246 B.n590 B.n589 585
R247 B.n579 B.n261 585
R248 B.n582 B.n261 585
R249 B.n581 B.n580 585
R250 B.n583 B.n581 585
R251 B.n578 B.n266 585
R252 B.n266 B.n265 585
R253 B.n577 B.n576 585
R254 B.n576 B.n575 585
R255 B.n268 B.n267 585
R256 B.n269 B.n268 585
R257 B.n568 B.n567 585
R258 B.n569 B.n568 585
R259 B.n566 B.n273 585
R260 B.n276 B.n273 585
R261 B.n565 B.n564 585
R262 B.n564 B.n563 585
R263 B.n275 B.n274 585
R264 B.n556 B.n275 585
R265 B.n555 B.n554 585
R266 B.n557 B.n555 585
R267 B.n553 B.n281 585
R268 B.n281 B.n280 585
R269 B.n552 B.n551 585
R270 B.n551 B.n550 585
R271 B.n283 B.n282 585
R272 B.n284 B.n283 585
R273 B.n543 B.n542 585
R274 B.n544 B.n543 585
R275 B.n541 B.n289 585
R276 B.n289 B.n288 585
R277 B.n540 B.n539 585
R278 B.n539 B.n538 585
R279 B.n291 B.n290 585
R280 B.n292 B.n291 585
R281 B.n531 B.n530 585
R282 B.n532 B.n531 585
R283 B.n529 B.n297 585
R284 B.n297 B.n296 585
R285 B.n528 B.n527 585
R286 B.n527 B.n526 585
R287 B.n299 B.n298 585
R288 B.n300 B.n299 585
R289 B.n519 B.n518 585
R290 B.n520 B.n519 585
R291 B.n303 B.n302 585
R292 B.n354 B.n353 585
R293 B.n355 B.n351 585
R294 B.n351 B.n304 585
R295 B.n357 B.n356 585
R296 B.n359 B.n350 585
R297 B.n362 B.n361 585
R298 B.n363 B.n349 585
R299 B.n365 B.n364 585
R300 B.n367 B.n348 585
R301 B.n370 B.n369 585
R302 B.n371 B.n347 585
R303 B.n373 B.n372 585
R304 B.n375 B.n346 585
R305 B.n378 B.n377 585
R306 B.n379 B.n345 585
R307 B.n381 B.n380 585
R308 B.n383 B.n344 585
R309 B.n386 B.n385 585
R310 B.n387 B.n343 585
R311 B.n389 B.n388 585
R312 B.n391 B.n342 585
R313 B.n394 B.n393 585
R314 B.n395 B.n341 585
R315 B.n397 B.n396 585
R316 B.n399 B.n340 585
R317 B.n402 B.n401 585
R318 B.n403 B.n339 585
R319 B.n405 B.n404 585
R320 B.n407 B.n338 585
R321 B.n410 B.n409 585
R322 B.n411 B.n337 585
R323 B.n413 B.n412 585
R324 B.n415 B.n336 585
R325 B.n418 B.n417 585
R326 B.n419 B.n335 585
R327 B.n421 B.n420 585
R328 B.n423 B.n334 585
R329 B.n426 B.n425 585
R330 B.n427 B.n330 585
R331 B.n429 B.n428 585
R332 B.n431 B.n329 585
R333 B.n434 B.n433 585
R334 B.n435 B.n328 585
R335 B.n437 B.n436 585
R336 B.n439 B.n327 585
R337 B.n442 B.n441 585
R338 B.n443 B.n324 585
R339 B.n446 B.n445 585
R340 B.n448 B.n323 585
R341 B.n451 B.n450 585
R342 B.n452 B.n322 585
R343 B.n454 B.n453 585
R344 B.n456 B.n321 585
R345 B.n459 B.n458 585
R346 B.n460 B.n320 585
R347 B.n462 B.n461 585
R348 B.n464 B.n319 585
R349 B.n467 B.n466 585
R350 B.n468 B.n318 585
R351 B.n470 B.n469 585
R352 B.n472 B.n317 585
R353 B.n475 B.n474 585
R354 B.n476 B.n316 585
R355 B.n478 B.n477 585
R356 B.n480 B.n315 585
R357 B.n483 B.n482 585
R358 B.n484 B.n314 585
R359 B.n486 B.n485 585
R360 B.n488 B.n313 585
R361 B.n491 B.n490 585
R362 B.n492 B.n312 585
R363 B.n494 B.n493 585
R364 B.n496 B.n311 585
R365 B.n499 B.n498 585
R366 B.n500 B.n310 585
R367 B.n502 B.n501 585
R368 B.n504 B.n309 585
R369 B.n507 B.n506 585
R370 B.n508 B.n308 585
R371 B.n510 B.n509 585
R372 B.n512 B.n307 585
R373 B.n513 B.n306 585
R374 B.n516 B.n515 585
R375 B.n517 B.n305 585
R376 B.n305 B.n304 585
R377 B.n522 B.n521 585
R378 B.n521 B.n520 585
R379 B.n523 B.n301 585
R380 B.n301 B.n300 585
R381 B.n525 B.n524 585
R382 B.n526 B.n525 585
R383 B.n295 B.n294 585
R384 B.n296 B.n295 585
R385 B.n534 B.n533 585
R386 B.n533 B.n532 585
R387 B.n535 B.n293 585
R388 B.n293 B.n292 585
R389 B.n537 B.n536 585
R390 B.n538 B.n537 585
R391 B.n287 B.n286 585
R392 B.n288 B.n287 585
R393 B.n546 B.n545 585
R394 B.n545 B.n544 585
R395 B.n547 B.n285 585
R396 B.n285 B.n284 585
R397 B.n549 B.n548 585
R398 B.n550 B.n549 585
R399 B.n279 B.n278 585
R400 B.n280 B.n279 585
R401 B.n559 B.n558 585
R402 B.n558 B.n557 585
R403 B.n560 B.n277 585
R404 B.n556 B.n277 585
R405 B.n562 B.n561 585
R406 B.n563 B.n562 585
R407 B.n272 B.n271 585
R408 B.n276 B.n272 585
R409 B.n571 B.n570 585
R410 B.n570 B.n569 585
R411 B.n572 B.n270 585
R412 B.n270 B.n269 585
R413 B.n574 B.n573 585
R414 B.n575 B.n574 585
R415 B.n264 B.n263 585
R416 B.n265 B.n264 585
R417 B.n585 B.n584 585
R418 B.n584 B.n583 585
R419 B.n586 B.n262 585
R420 B.n582 B.n262 585
R421 B.n588 B.n587 585
R422 B.n589 B.n588 585
R423 B.n3 B.n0 585
R424 B.n4 B.n3 585
R425 B.n676 B.n1 585
R426 B.n677 B.n676 585
R427 B.n675 B.n674 585
R428 B.n675 B.n8 585
R429 B.n673 B.n9 585
R430 B.n12 B.n9 585
R431 B.n672 B.n671 585
R432 B.n671 B.n670 585
R433 B.n11 B.n10 585
R434 B.n669 B.n11 585
R435 B.n667 B.n666 585
R436 B.n668 B.n667 585
R437 B.n665 B.n17 585
R438 B.n17 B.n16 585
R439 B.n664 B.n663 585
R440 B.n663 B.n662 585
R441 B.n19 B.n18 585
R442 B.n661 B.n19 585
R443 B.n659 B.n658 585
R444 B.n660 B.n659 585
R445 B.n657 B.n23 585
R446 B.n26 B.n23 585
R447 B.n656 B.n655 585
R448 B.n655 B.n654 585
R449 B.n25 B.n24 585
R450 B.n653 B.n25 585
R451 B.n651 B.n650 585
R452 B.n652 B.n651 585
R453 B.n649 B.n31 585
R454 B.n31 B.n30 585
R455 B.n648 B.n647 585
R456 B.n647 B.n646 585
R457 B.n33 B.n32 585
R458 B.n645 B.n33 585
R459 B.n643 B.n642 585
R460 B.n644 B.n643 585
R461 B.n641 B.n38 585
R462 B.n38 B.n37 585
R463 B.n640 B.n639 585
R464 B.n639 B.n638 585
R465 B.n40 B.n39 585
R466 B.n637 B.n40 585
R467 B.n635 B.n634 585
R468 B.n636 B.n635 585
R469 B.n633 B.n45 585
R470 B.n45 B.n44 585
R471 B.n632 B.n631 585
R472 B.n631 B.n630 585
R473 B.n680 B.n679 585
R474 B.n678 B.n2 585
R475 B.n631 B.n47 530.939
R476 B.n627 B.n48 530.939
R477 B.n519 B.n305 530.939
R478 B.n521 B.n303 530.939
R479 B.n629 B.n628 256.663
R480 B.n629 B.n89 256.663
R481 B.n629 B.n88 256.663
R482 B.n629 B.n87 256.663
R483 B.n629 B.n86 256.663
R484 B.n629 B.n85 256.663
R485 B.n629 B.n84 256.663
R486 B.n629 B.n83 256.663
R487 B.n629 B.n82 256.663
R488 B.n629 B.n81 256.663
R489 B.n629 B.n80 256.663
R490 B.n629 B.n79 256.663
R491 B.n629 B.n78 256.663
R492 B.n629 B.n77 256.663
R493 B.n629 B.n76 256.663
R494 B.n629 B.n75 256.663
R495 B.n629 B.n74 256.663
R496 B.n629 B.n73 256.663
R497 B.n629 B.n72 256.663
R498 B.n629 B.n71 256.663
R499 B.n629 B.n70 256.663
R500 B.n629 B.n69 256.663
R501 B.n629 B.n68 256.663
R502 B.n629 B.n67 256.663
R503 B.n629 B.n66 256.663
R504 B.n629 B.n65 256.663
R505 B.n629 B.n64 256.663
R506 B.n629 B.n63 256.663
R507 B.n629 B.n62 256.663
R508 B.n629 B.n61 256.663
R509 B.n629 B.n60 256.663
R510 B.n629 B.n59 256.663
R511 B.n629 B.n58 256.663
R512 B.n629 B.n57 256.663
R513 B.n629 B.n56 256.663
R514 B.n629 B.n55 256.663
R515 B.n629 B.n54 256.663
R516 B.n629 B.n53 256.663
R517 B.n629 B.n52 256.663
R518 B.n629 B.n51 256.663
R519 B.n629 B.n50 256.663
R520 B.n629 B.n49 256.663
R521 B.n352 B.n304 256.663
R522 B.n358 B.n304 256.663
R523 B.n360 B.n304 256.663
R524 B.n366 B.n304 256.663
R525 B.n368 B.n304 256.663
R526 B.n374 B.n304 256.663
R527 B.n376 B.n304 256.663
R528 B.n382 B.n304 256.663
R529 B.n384 B.n304 256.663
R530 B.n390 B.n304 256.663
R531 B.n392 B.n304 256.663
R532 B.n398 B.n304 256.663
R533 B.n400 B.n304 256.663
R534 B.n406 B.n304 256.663
R535 B.n408 B.n304 256.663
R536 B.n414 B.n304 256.663
R537 B.n416 B.n304 256.663
R538 B.n422 B.n304 256.663
R539 B.n424 B.n304 256.663
R540 B.n430 B.n304 256.663
R541 B.n432 B.n304 256.663
R542 B.n438 B.n304 256.663
R543 B.n440 B.n304 256.663
R544 B.n447 B.n304 256.663
R545 B.n449 B.n304 256.663
R546 B.n455 B.n304 256.663
R547 B.n457 B.n304 256.663
R548 B.n463 B.n304 256.663
R549 B.n465 B.n304 256.663
R550 B.n471 B.n304 256.663
R551 B.n473 B.n304 256.663
R552 B.n479 B.n304 256.663
R553 B.n481 B.n304 256.663
R554 B.n487 B.n304 256.663
R555 B.n489 B.n304 256.663
R556 B.n495 B.n304 256.663
R557 B.n497 B.n304 256.663
R558 B.n503 B.n304 256.663
R559 B.n505 B.n304 256.663
R560 B.n511 B.n304 256.663
R561 B.n514 B.n304 256.663
R562 B.n682 B.n681 256.663
R563 B.n97 B.n96 163.367
R564 B.n101 B.n100 163.367
R565 B.n105 B.n104 163.367
R566 B.n109 B.n108 163.367
R567 B.n113 B.n112 163.367
R568 B.n117 B.n116 163.367
R569 B.n121 B.n120 163.367
R570 B.n125 B.n124 163.367
R571 B.n129 B.n128 163.367
R572 B.n133 B.n132 163.367
R573 B.n137 B.n136 163.367
R574 B.n141 B.n140 163.367
R575 B.n145 B.n144 163.367
R576 B.n149 B.n148 163.367
R577 B.n153 B.n152 163.367
R578 B.n157 B.n156 163.367
R579 B.n161 B.n160 163.367
R580 B.n165 B.n164 163.367
R581 B.n170 B.n169 163.367
R582 B.n174 B.n173 163.367
R583 B.n178 B.n177 163.367
R584 B.n182 B.n181 163.367
R585 B.n186 B.n185 163.367
R586 B.n191 B.n190 163.367
R587 B.n195 B.n194 163.367
R588 B.n199 B.n198 163.367
R589 B.n203 B.n202 163.367
R590 B.n207 B.n206 163.367
R591 B.n211 B.n210 163.367
R592 B.n215 B.n214 163.367
R593 B.n219 B.n218 163.367
R594 B.n223 B.n222 163.367
R595 B.n227 B.n226 163.367
R596 B.n231 B.n230 163.367
R597 B.n235 B.n234 163.367
R598 B.n239 B.n238 163.367
R599 B.n243 B.n242 163.367
R600 B.n247 B.n246 163.367
R601 B.n251 B.n250 163.367
R602 B.n255 B.n254 163.367
R603 B.n257 B.n90 163.367
R604 B.n519 B.n299 163.367
R605 B.n527 B.n299 163.367
R606 B.n527 B.n297 163.367
R607 B.n531 B.n297 163.367
R608 B.n531 B.n291 163.367
R609 B.n539 B.n291 163.367
R610 B.n539 B.n289 163.367
R611 B.n543 B.n289 163.367
R612 B.n543 B.n283 163.367
R613 B.n551 B.n283 163.367
R614 B.n551 B.n281 163.367
R615 B.n555 B.n281 163.367
R616 B.n555 B.n275 163.367
R617 B.n564 B.n275 163.367
R618 B.n564 B.n273 163.367
R619 B.n568 B.n273 163.367
R620 B.n568 B.n268 163.367
R621 B.n576 B.n268 163.367
R622 B.n576 B.n266 163.367
R623 B.n581 B.n266 163.367
R624 B.n581 B.n261 163.367
R625 B.n590 B.n261 163.367
R626 B.n591 B.n590 163.367
R627 B.n591 B.n5 163.367
R628 B.n6 B.n5 163.367
R629 B.n7 B.n6 163.367
R630 B.n597 B.n7 163.367
R631 B.n598 B.n597 163.367
R632 B.n598 B.n13 163.367
R633 B.n14 B.n13 163.367
R634 B.n15 B.n14 163.367
R635 B.n603 B.n15 163.367
R636 B.n603 B.n20 163.367
R637 B.n21 B.n20 163.367
R638 B.n22 B.n21 163.367
R639 B.n608 B.n22 163.367
R640 B.n608 B.n27 163.367
R641 B.n28 B.n27 163.367
R642 B.n29 B.n28 163.367
R643 B.n613 B.n29 163.367
R644 B.n613 B.n34 163.367
R645 B.n35 B.n34 163.367
R646 B.n36 B.n35 163.367
R647 B.n618 B.n36 163.367
R648 B.n618 B.n41 163.367
R649 B.n42 B.n41 163.367
R650 B.n43 B.n42 163.367
R651 B.n623 B.n43 163.367
R652 B.n623 B.n48 163.367
R653 B.n353 B.n351 163.367
R654 B.n357 B.n351 163.367
R655 B.n361 B.n359 163.367
R656 B.n365 B.n349 163.367
R657 B.n369 B.n367 163.367
R658 B.n373 B.n347 163.367
R659 B.n377 B.n375 163.367
R660 B.n381 B.n345 163.367
R661 B.n385 B.n383 163.367
R662 B.n389 B.n343 163.367
R663 B.n393 B.n391 163.367
R664 B.n397 B.n341 163.367
R665 B.n401 B.n399 163.367
R666 B.n405 B.n339 163.367
R667 B.n409 B.n407 163.367
R668 B.n413 B.n337 163.367
R669 B.n417 B.n415 163.367
R670 B.n421 B.n335 163.367
R671 B.n425 B.n423 163.367
R672 B.n429 B.n330 163.367
R673 B.n433 B.n431 163.367
R674 B.n437 B.n328 163.367
R675 B.n441 B.n439 163.367
R676 B.n446 B.n324 163.367
R677 B.n450 B.n448 163.367
R678 B.n454 B.n322 163.367
R679 B.n458 B.n456 163.367
R680 B.n462 B.n320 163.367
R681 B.n466 B.n464 163.367
R682 B.n470 B.n318 163.367
R683 B.n474 B.n472 163.367
R684 B.n478 B.n316 163.367
R685 B.n482 B.n480 163.367
R686 B.n486 B.n314 163.367
R687 B.n490 B.n488 163.367
R688 B.n494 B.n312 163.367
R689 B.n498 B.n496 163.367
R690 B.n502 B.n310 163.367
R691 B.n506 B.n504 163.367
R692 B.n510 B.n308 163.367
R693 B.n513 B.n512 163.367
R694 B.n515 B.n305 163.367
R695 B.n521 B.n301 163.367
R696 B.n525 B.n301 163.367
R697 B.n525 B.n295 163.367
R698 B.n533 B.n295 163.367
R699 B.n533 B.n293 163.367
R700 B.n537 B.n293 163.367
R701 B.n537 B.n287 163.367
R702 B.n545 B.n287 163.367
R703 B.n545 B.n285 163.367
R704 B.n549 B.n285 163.367
R705 B.n549 B.n279 163.367
R706 B.n558 B.n279 163.367
R707 B.n558 B.n277 163.367
R708 B.n562 B.n277 163.367
R709 B.n562 B.n272 163.367
R710 B.n570 B.n272 163.367
R711 B.n570 B.n270 163.367
R712 B.n574 B.n270 163.367
R713 B.n574 B.n264 163.367
R714 B.n584 B.n264 163.367
R715 B.n584 B.n262 163.367
R716 B.n588 B.n262 163.367
R717 B.n588 B.n3 163.367
R718 B.n680 B.n3 163.367
R719 B.n676 B.n2 163.367
R720 B.n676 B.n675 163.367
R721 B.n675 B.n9 163.367
R722 B.n671 B.n9 163.367
R723 B.n671 B.n11 163.367
R724 B.n667 B.n11 163.367
R725 B.n667 B.n17 163.367
R726 B.n663 B.n17 163.367
R727 B.n663 B.n19 163.367
R728 B.n659 B.n19 163.367
R729 B.n659 B.n23 163.367
R730 B.n655 B.n23 163.367
R731 B.n655 B.n25 163.367
R732 B.n651 B.n25 163.367
R733 B.n651 B.n31 163.367
R734 B.n647 B.n31 163.367
R735 B.n647 B.n33 163.367
R736 B.n643 B.n33 163.367
R737 B.n643 B.n38 163.367
R738 B.n639 B.n38 163.367
R739 B.n639 B.n40 163.367
R740 B.n635 B.n40 163.367
R741 B.n635 B.n45 163.367
R742 B.n631 B.n45 163.367
R743 B.n520 B.n304 95.5314
R744 B.n630 B.n629 95.5314
R745 B.n91 B.t13 92.0716
R746 B.n325 B.t17 92.0716
R747 B.n93 B.t19 92.0589
R748 B.n331 B.t10 92.0589
R749 B.n92 B.t14 73.8413
R750 B.n326 B.t16 73.8413
R751 B.n94 B.t20 73.8286
R752 B.n332 B.t9 73.8286
R753 B.n49 B.n47 71.676
R754 B.n97 B.n50 71.676
R755 B.n101 B.n51 71.676
R756 B.n105 B.n52 71.676
R757 B.n109 B.n53 71.676
R758 B.n113 B.n54 71.676
R759 B.n117 B.n55 71.676
R760 B.n121 B.n56 71.676
R761 B.n125 B.n57 71.676
R762 B.n129 B.n58 71.676
R763 B.n133 B.n59 71.676
R764 B.n137 B.n60 71.676
R765 B.n141 B.n61 71.676
R766 B.n145 B.n62 71.676
R767 B.n149 B.n63 71.676
R768 B.n153 B.n64 71.676
R769 B.n157 B.n65 71.676
R770 B.n161 B.n66 71.676
R771 B.n165 B.n67 71.676
R772 B.n170 B.n68 71.676
R773 B.n174 B.n69 71.676
R774 B.n178 B.n70 71.676
R775 B.n182 B.n71 71.676
R776 B.n186 B.n72 71.676
R777 B.n191 B.n73 71.676
R778 B.n195 B.n74 71.676
R779 B.n199 B.n75 71.676
R780 B.n203 B.n76 71.676
R781 B.n207 B.n77 71.676
R782 B.n211 B.n78 71.676
R783 B.n215 B.n79 71.676
R784 B.n219 B.n80 71.676
R785 B.n223 B.n81 71.676
R786 B.n227 B.n82 71.676
R787 B.n231 B.n83 71.676
R788 B.n235 B.n84 71.676
R789 B.n239 B.n85 71.676
R790 B.n243 B.n86 71.676
R791 B.n247 B.n87 71.676
R792 B.n251 B.n88 71.676
R793 B.n255 B.n89 71.676
R794 B.n628 B.n90 71.676
R795 B.n628 B.n627 71.676
R796 B.n257 B.n89 71.676
R797 B.n254 B.n88 71.676
R798 B.n250 B.n87 71.676
R799 B.n246 B.n86 71.676
R800 B.n242 B.n85 71.676
R801 B.n238 B.n84 71.676
R802 B.n234 B.n83 71.676
R803 B.n230 B.n82 71.676
R804 B.n226 B.n81 71.676
R805 B.n222 B.n80 71.676
R806 B.n218 B.n79 71.676
R807 B.n214 B.n78 71.676
R808 B.n210 B.n77 71.676
R809 B.n206 B.n76 71.676
R810 B.n202 B.n75 71.676
R811 B.n198 B.n74 71.676
R812 B.n194 B.n73 71.676
R813 B.n190 B.n72 71.676
R814 B.n185 B.n71 71.676
R815 B.n181 B.n70 71.676
R816 B.n177 B.n69 71.676
R817 B.n173 B.n68 71.676
R818 B.n169 B.n67 71.676
R819 B.n164 B.n66 71.676
R820 B.n160 B.n65 71.676
R821 B.n156 B.n64 71.676
R822 B.n152 B.n63 71.676
R823 B.n148 B.n62 71.676
R824 B.n144 B.n61 71.676
R825 B.n140 B.n60 71.676
R826 B.n136 B.n59 71.676
R827 B.n132 B.n58 71.676
R828 B.n128 B.n57 71.676
R829 B.n124 B.n56 71.676
R830 B.n120 B.n55 71.676
R831 B.n116 B.n54 71.676
R832 B.n112 B.n53 71.676
R833 B.n108 B.n52 71.676
R834 B.n104 B.n51 71.676
R835 B.n100 B.n50 71.676
R836 B.n96 B.n49 71.676
R837 B.n352 B.n303 71.676
R838 B.n358 B.n357 71.676
R839 B.n361 B.n360 71.676
R840 B.n366 B.n365 71.676
R841 B.n369 B.n368 71.676
R842 B.n374 B.n373 71.676
R843 B.n377 B.n376 71.676
R844 B.n382 B.n381 71.676
R845 B.n385 B.n384 71.676
R846 B.n390 B.n389 71.676
R847 B.n393 B.n392 71.676
R848 B.n398 B.n397 71.676
R849 B.n401 B.n400 71.676
R850 B.n406 B.n405 71.676
R851 B.n409 B.n408 71.676
R852 B.n414 B.n413 71.676
R853 B.n417 B.n416 71.676
R854 B.n422 B.n421 71.676
R855 B.n425 B.n424 71.676
R856 B.n430 B.n429 71.676
R857 B.n433 B.n432 71.676
R858 B.n438 B.n437 71.676
R859 B.n441 B.n440 71.676
R860 B.n447 B.n446 71.676
R861 B.n450 B.n449 71.676
R862 B.n455 B.n454 71.676
R863 B.n458 B.n457 71.676
R864 B.n463 B.n462 71.676
R865 B.n466 B.n465 71.676
R866 B.n471 B.n470 71.676
R867 B.n474 B.n473 71.676
R868 B.n479 B.n478 71.676
R869 B.n482 B.n481 71.676
R870 B.n487 B.n486 71.676
R871 B.n490 B.n489 71.676
R872 B.n495 B.n494 71.676
R873 B.n498 B.n497 71.676
R874 B.n503 B.n502 71.676
R875 B.n506 B.n505 71.676
R876 B.n511 B.n510 71.676
R877 B.n514 B.n513 71.676
R878 B.n353 B.n352 71.676
R879 B.n359 B.n358 71.676
R880 B.n360 B.n349 71.676
R881 B.n367 B.n366 71.676
R882 B.n368 B.n347 71.676
R883 B.n375 B.n374 71.676
R884 B.n376 B.n345 71.676
R885 B.n383 B.n382 71.676
R886 B.n384 B.n343 71.676
R887 B.n391 B.n390 71.676
R888 B.n392 B.n341 71.676
R889 B.n399 B.n398 71.676
R890 B.n400 B.n339 71.676
R891 B.n407 B.n406 71.676
R892 B.n408 B.n337 71.676
R893 B.n415 B.n414 71.676
R894 B.n416 B.n335 71.676
R895 B.n423 B.n422 71.676
R896 B.n424 B.n330 71.676
R897 B.n431 B.n430 71.676
R898 B.n432 B.n328 71.676
R899 B.n439 B.n438 71.676
R900 B.n440 B.n324 71.676
R901 B.n448 B.n447 71.676
R902 B.n449 B.n322 71.676
R903 B.n456 B.n455 71.676
R904 B.n457 B.n320 71.676
R905 B.n464 B.n463 71.676
R906 B.n465 B.n318 71.676
R907 B.n472 B.n471 71.676
R908 B.n473 B.n316 71.676
R909 B.n480 B.n479 71.676
R910 B.n481 B.n314 71.676
R911 B.n488 B.n487 71.676
R912 B.n489 B.n312 71.676
R913 B.n496 B.n495 71.676
R914 B.n497 B.n310 71.676
R915 B.n504 B.n503 71.676
R916 B.n505 B.n308 71.676
R917 B.n512 B.n511 71.676
R918 B.n515 B.n514 71.676
R919 B.n681 B.n680 71.676
R920 B.n681 B.n2 71.676
R921 B.n167 B.n94 59.5399
R922 B.n188 B.n92 59.5399
R923 B.n444 B.n326 59.5399
R924 B.n333 B.n332 59.5399
R925 B.n520 B.n300 47.4173
R926 B.n526 B.n300 47.4173
R927 B.n526 B.n296 47.4173
R928 B.n532 B.n296 47.4173
R929 B.n538 B.n292 47.4173
R930 B.n538 B.n288 47.4173
R931 B.n544 B.n288 47.4173
R932 B.n544 B.n284 47.4173
R933 B.n550 B.n284 47.4173
R934 B.n557 B.n280 47.4173
R935 B.n557 B.n556 47.4173
R936 B.n563 B.n276 47.4173
R937 B.n569 B.n269 47.4173
R938 B.n575 B.n269 47.4173
R939 B.n583 B.n265 47.4173
R940 B.n583 B.n582 47.4173
R941 B.n589 B.n4 47.4173
R942 B.n679 B.n4 47.4173
R943 B.n679 B.n678 47.4173
R944 B.n678 B.n677 47.4173
R945 B.n677 B.n8 47.4173
R946 B.n670 B.n12 47.4173
R947 B.n670 B.n669 47.4173
R948 B.n668 B.n16 47.4173
R949 B.n662 B.n16 47.4173
R950 B.n661 B.n660 47.4173
R951 B.n654 B.n26 47.4173
R952 B.n654 B.n653 47.4173
R953 B.n652 B.n30 47.4173
R954 B.n646 B.n30 47.4173
R955 B.n646 B.n645 47.4173
R956 B.n645 B.n644 47.4173
R957 B.n644 B.n37 47.4173
R958 B.n638 B.n637 47.4173
R959 B.n637 B.n636 47.4173
R960 B.n636 B.n44 47.4173
R961 B.n630 B.n44 47.4173
R962 B.n276 B.t1 46.72
R963 B.t21 B.n661 46.72
R964 B.n563 B.t4 36.9577
R965 B.n660 B.t5 36.9577
R966 B.n575 B.t3 35.5631
R967 B.t22 B.n668 35.5631
R968 B.n522 B.n302 34.4981
R969 B.n518 B.n517 34.4981
R970 B.n626 B.n625 34.4981
R971 B.n632 B.n46 34.4981
R972 B.t6 B.n280 25.8008
R973 B.n653 B.t23 25.8008
R974 B.t8 B.n292 24.4062
R975 B.n582 B.t0 24.4062
R976 B.n12 B.t2 24.4062
R977 B.t12 B.n37 24.4062
R978 B.n532 B.t8 23.0116
R979 B.n589 B.t0 23.0116
R980 B.t2 B.n8 23.0116
R981 B.n638 B.t12 23.0116
R982 B.n550 B.t6 21.617
R983 B.t23 B.n652 21.617
R984 B.n94 B.n93 18.2308
R985 B.n92 B.n91 18.2308
R986 B.n326 B.n325 18.2308
R987 B.n332 B.n331 18.2308
R988 B B.n682 18.0485
R989 B.t3 B.n265 11.8547
R990 B.n669 B.t22 11.8547
R991 B.n523 B.n522 10.6151
R992 B.n524 B.n523 10.6151
R993 B.n524 B.n294 10.6151
R994 B.n534 B.n294 10.6151
R995 B.n535 B.n534 10.6151
R996 B.n536 B.n535 10.6151
R997 B.n536 B.n286 10.6151
R998 B.n546 B.n286 10.6151
R999 B.n547 B.n546 10.6151
R1000 B.n548 B.n547 10.6151
R1001 B.n548 B.n278 10.6151
R1002 B.n559 B.n278 10.6151
R1003 B.n560 B.n559 10.6151
R1004 B.n561 B.n560 10.6151
R1005 B.n561 B.n271 10.6151
R1006 B.n571 B.n271 10.6151
R1007 B.n572 B.n571 10.6151
R1008 B.n573 B.n572 10.6151
R1009 B.n573 B.n263 10.6151
R1010 B.n585 B.n263 10.6151
R1011 B.n586 B.n585 10.6151
R1012 B.n587 B.n586 10.6151
R1013 B.n587 B.n0 10.6151
R1014 B.n354 B.n302 10.6151
R1015 B.n355 B.n354 10.6151
R1016 B.n356 B.n355 10.6151
R1017 B.n356 B.n350 10.6151
R1018 B.n362 B.n350 10.6151
R1019 B.n363 B.n362 10.6151
R1020 B.n364 B.n363 10.6151
R1021 B.n364 B.n348 10.6151
R1022 B.n370 B.n348 10.6151
R1023 B.n371 B.n370 10.6151
R1024 B.n372 B.n371 10.6151
R1025 B.n372 B.n346 10.6151
R1026 B.n378 B.n346 10.6151
R1027 B.n379 B.n378 10.6151
R1028 B.n380 B.n379 10.6151
R1029 B.n380 B.n344 10.6151
R1030 B.n386 B.n344 10.6151
R1031 B.n387 B.n386 10.6151
R1032 B.n388 B.n387 10.6151
R1033 B.n388 B.n342 10.6151
R1034 B.n394 B.n342 10.6151
R1035 B.n395 B.n394 10.6151
R1036 B.n396 B.n395 10.6151
R1037 B.n396 B.n340 10.6151
R1038 B.n402 B.n340 10.6151
R1039 B.n403 B.n402 10.6151
R1040 B.n404 B.n403 10.6151
R1041 B.n404 B.n338 10.6151
R1042 B.n410 B.n338 10.6151
R1043 B.n411 B.n410 10.6151
R1044 B.n412 B.n411 10.6151
R1045 B.n412 B.n336 10.6151
R1046 B.n418 B.n336 10.6151
R1047 B.n419 B.n418 10.6151
R1048 B.n420 B.n419 10.6151
R1049 B.n420 B.n334 10.6151
R1050 B.n427 B.n426 10.6151
R1051 B.n428 B.n427 10.6151
R1052 B.n428 B.n329 10.6151
R1053 B.n434 B.n329 10.6151
R1054 B.n435 B.n434 10.6151
R1055 B.n436 B.n435 10.6151
R1056 B.n436 B.n327 10.6151
R1057 B.n442 B.n327 10.6151
R1058 B.n443 B.n442 10.6151
R1059 B.n445 B.n323 10.6151
R1060 B.n451 B.n323 10.6151
R1061 B.n452 B.n451 10.6151
R1062 B.n453 B.n452 10.6151
R1063 B.n453 B.n321 10.6151
R1064 B.n459 B.n321 10.6151
R1065 B.n460 B.n459 10.6151
R1066 B.n461 B.n460 10.6151
R1067 B.n461 B.n319 10.6151
R1068 B.n467 B.n319 10.6151
R1069 B.n468 B.n467 10.6151
R1070 B.n469 B.n468 10.6151
R1071 B.n469 B.n317 10.6151
R1072 B.n475 B.n317 10.6151
R1073 B.n476 B.n475 10.6151
R1074 B.n477 B.n476 10.6151
R1075 B.n477 B.n315 10.6151
R1076 B.n483 B.n315 10.6151
R1077 B.n484 B.n483 10.6151
R1078 B.n485 B.n484 10.6151
R1079 B.n485 B.n313 10.6151
R1080 B.n491 B.n313 10.6151
R1081 B.n492 B.n491 10.6151
R1082 B.n493 B.n492 10.6151
R1083 B.n493 B.n311 10.6151
R1084 B.n499 B.n311 10.6151
R1085 B.n500 B.n499 10.6151
R1086 B.n501 B.n500 10.6151
R1087 B.n501 B.n309 10.6151
R1088 B.n507 B.n309 10.6151
R1089 B.n508 B.n507 10.6151
R1090 B.n509 B.n508 10.6151
R1091 B.n509 B.n307 10.6151
R1092 B.n307 B.n306 10.6151
R1093 B.n516 B.n306 10.6151
R1094 B.n517 B.n516 10.6151
R1095 B.n518 B.n298 10.6151
R1096 B.n528 B.n298 10.6151
R1097 B.n529 B.n528 10.6151
R1098 B.n530 B.n529 10.6151
R1099 B.n530 B.n290 10.6151
R1100 B.n540 B.n290 10.6151
R1101 B.n541 B.n540 10.6151
R1102 B.n542 B.n541 10.6151
R1103 B.n542 B.n282 10.6151
R1104 B.n552 B.n282 10.6151
R1105 B.n553 B.n552 10.6151
R1106 B.n554 B.n553 10.6151
R1107 B.n554 B.n274 10.6151
R1108 B.n565 B.n274 10.6151
R1109 B.n566 B.n565 10.6151
R1110 B.n567 B.n566 10.6151
R1111 B.n567 B.n267 10.6151
R1112 B.n577 B.n267 10.6151
R1113 B.n578 B.n577 10.6151
R1114 B.n580 B.n578 10.6151
R1115 B.n580 B.n579 10.6151
R1116 B.n579 B.n260 10.6151
R1117 B.n592 B.n260 10.6151
R1118 B.n593 B.n592 10.6151
R1119 B.n594 B.n593 10.6151
R1120 B.n595 B.n594 10.6151
R1121 B.n596 B.n595 10.6151
R1122 B.n599 B.n596 10.6151
R1123 B.n600 B.n599 10.6151
R1124 B.n601 B.n600 10.6151
R1125 B.n602 B.n601 10.6151
R1126 B.n604 B.n602 10.6151
R1127 B.n605 B.n604 10.6151
R1128 B.n606 B.n605 10.6151
R1129 B.n607 B.n606 10.6151
R1130 B.n609 B.n607 10.6151
R1131 B.n610 B.n609 10.6151
R1132 B.n611 B.n610 10.6151
R1133 B.n612 B.n611 10.6151
R1134 B.n614 B.n612 10.6151
R1135 B.n615 B.n614 10.6151
R1136 B.n616 B.n615 10.6151
R1137 B.n617 B.n616 10.6151
R1138 B.n619 B.n617 10.6151
R1139 B.n620 B.n619 10.6151
R1140 B.n621 B.n620 10.6151
R1141 B.n622 B.n621 10.6151
R1142 B.n624 B.n622 10.6151
R1143 B.n625 B.n624 10.6151
R1144 B.n674 B.n1 10.6151
R1145 B.n674 B.n673 10.6151
R1146 B.n673 B.n672 10.6151
R1147 B.n672 B.n10 10.6151
R1148 B.n666 B.n10 10.6151
R1149 B.n666 B.n665 10.6151
R1150 B.n665 B.n664 10.6151
R1151 B.n664 B.n18 10.6151
R1152 B.n658 B.n18 10.6151
R1153 B.n658 B.n657 10.6151
R1154 B.n657 B.n656 10.6151
R1155 B.n656 B.n24 10.6151
R1156 B.n650 B.n24 10.6151
R1157 B.n650 B.n649 10.6151
R1158 B.n649 B.n648 10.6151
R1159 B.n648 B.n32 10.6151
R1160 B.n642 B.n32 10.6151
R1161 B.n642 B.n641 10.6151
R1162 B.n641 B.n640 10.6151
R1163 B.n640 B.n39 10.6151
R1164 B.n634 B.n39 10.6151
R1165 B.n634 B.n633 10.6151
R1166 B.n633 B.n632 10.6151
R1167 B.n95 B.n46 10.6151
R1168 B.n98 B.n95 10.6151
R1169 B.n99 B.n98 10.6151
R1170 B.n102 B.n99 10.6151
R1171 B.n103 B.n102 10.6151
R1172 B.n106 B.n103 10.6151
R1173 B.n107 B.n106 10.6151
R1174 B.n110 B.n107 10.6151
R1175 B.n111 B.n110 10.6151
R1176 B.n114 B.n111 10.6151
R1177 B.n115 B.n114 10.6151
R1178 B.n118 B.n115 10.6151
R1179 B.n119 B.n118 10.6151
R1180 B.n122 B.n119 10.6151
R1181 B.n123 B.n122 10.6151
R1182 B.n126 B.n123 10.6151
R1183 B.n127 B.n126 10.6151
R1184 B.n130 B.n127 10.6151
R1185 B.n131 B.n130 10.6151
R1186 B.n134 B.n131 10.6151
R1187 B.n135 B.n134 10.6151
R1188 B.n138 B.n135 10.6151
R1189 B.n139 B.n138 10.6151
R1190 B.n142 B.n139 10.6151
R1191 B.n143 B.n142 10.6151
R1192 B.n146 B.n143 10.6151
R1193 B.n147 B.n146 10.6151
R1194 B.n150 B.n147 10.6151
R1195 B.n151 B.n150 10.6151
R1196 B.n154 B.n151 10.6151
R1197 B.n155 B.n154 10.6151
R1198 B.n158 B.n155 10.6151
R1199 B.n159 B.n158 10.6151
R1200 B.n162 B.n159 10.6151
R1201 B.n163 B.n162 10.6151
R1202 B.n166 B.n163 10.6151
R1203 B.n171 B.n168 10.6151
R1204 B.n172 B.n171 10.6151
R1205 B.n175 B.n172 10.6151
R1206 B.n176 B.n175 10.6151
R1207 B.n179 B.n176 10.6151
R1208 B.n180 B.n179 10.6151
R1209 B.n183 B.n180 10.6151
R1210 B.n184 B.n183 10.6151
R1211 B.n187 B.n184 10.6151
R1212 B.n192 B.n189 10.6151
R1213 B.n193 B.n192 10.6151
R1214 B.n196 B.n193 10.6151
R1215 B.n197 B.n196 10.6151
R1216 B.n200 B.n197 10.6151
R1217 B.n201 B.n200 10.6151
R1218 B.n204 B.n201 10.6151
R1219 B.n205 B.n204 10.6151
R1220 B.n208 B.n205 10.6151
R1221 B.n209 B.n208 10.6151
R1222 B.n212 B.n209 10.6151
R1223 B.n213 B.n212 10.6151
R1224 B.n216 B.n213 10.6151
R1225 B.n217 B.n216 10.6151
R1226 B.n220 B.n217 10.6151
R1227 B.n221 B.n220 10.6151
R1228 B.n224 B.n221 10.6151
R1229 B.n225 B.n224 10.6151
R1230 B.n228 B.n225 10.6151
R1231 B.n229 B.n228 10.6151
R1232 B.n232 B.n229 10.6151
R1233 B.n233 B.n232 10.6151
R1234 B.n236 B.n233 10.6151
R1235 B.n237 B.n236 10.6151
R1236 B.n240 B.n237 10.6151
R1237 B.n241 B.n240 10.6151
R1238 B.n244 B.n241 10.6151
R1239 B.n245 B.n244 10.6151
R1240 B.n248 B.n245 10.6151
R1241 B.n249 B.n248 10.6151
R1242 B.n252 B.n249 10.6151
R1243 B.n253 B.n252 10.6151
R1244 B.n256 B.n253 10.6151
R1245 B.n258 B.n256 10.6151
R1246 B.n259 B.n258 10.6151
R1247 B.n626 B.n259 10.6151
R1248 B.n556 B.t4 10.4601
R1249 B.n26 B.t5 10.4601
R1250 B.n334 B.n333 9.36635
R1251 B.n445 B.n444 9.36635
R1252 B.n167 B.n166 9.36635
R1253 B.n189 B.n188 9.36635
R1254 B.n682 B.n0 8.11757
R1255 B.n682 B.n1 8.11757
R1256 B.n426 B.n333 1.24928
R1257 B.n444 B.n443 1.24928
R1258 B.n168 B.n167 1.24928
R1259 B.n188 B.n187 1.24928
R1260 B.n569 B.t1 0.697806
R1261 B.n662 B.t21 0.697806
R1262 VN.n3 VN.t9 505.904
R1263 VN.n13 VN.t6 505.904
R1264 VN.n2 VN.t4 479.235
R1265 VN.n1 VN.t2 479.235
R1266 VN.n6 VN.t0 479.235
R1267 VN.n8 VN.t7 479.235
R1268 VN.n12 VN.t8 479.235
R1269 VN.n11 VN.t1 479.235
R1270 VN.n16 VN.t3 479.235
R1271 VN.n18 VN.t5 479.235
R1272 VN.n9 VN.n8 161.3
R1273 VN.n19 VN.n18 161.3
R1274 VN.n17 VN.n10 161.3
R1275 VN.n16 VN.n15 161.3
R1276 VN.n7 VN.n0 161.3
R1277 VN.n6 VN.n5 161.3
R1278 VN.n14 VN.n11 80.6037
R1279 VN.n4 VN.n1 80.6037
R1280 VN.n2 VN.n1 48.2005
R1281 VN.n6 VN.n1 48.2005
R1282 VN.n12 VN.n11 48.2005
R1283 VN.n16 VN.n11 48.2005
R1284 VN.n8 VN.n7 47.4702
R1285 VN.n18 VN.n17 47.4702
R1286 VN.n14 VN.n13 45.2144
R1287 VN.n4 VN.n3 45.2144
R1288 VN VN.n19 41.5706
R1289 VN.n3 VN.n2 13.6377
R1290 VN.n13 VN.n12 13.6377
R1291 VN.n7 VN.n6 0.730803
R1292 VN.n17 VN.n16 0.730803
R1293 VN.n15 VN.n14 0.285035
R1294 VN.n5 VN.n4 0.285035
R1295 VN.n19 VN.n10 0.189894
R1296 VN.n15 VN.n10 0.189894
R1297 VN.n5 VN.n0 0.189894
R1298 VN.n9 VN.n0 0.189894
R1299 VN VN.n9 0.0516364
R1300 VDD2.n1 VDD2.t0 68.6697
R1301 VDD2.n4 VDD2.t4 67.8596
R1302 VDD2.n3 VDD2.n2 66.5261
R1303 VDD2 VDD2.n7 66.5233
R1304 VDD2.n6 VDD2.n5 65.9739
R1305 VDD2.n1 VDD2.n0 65.9737
R1306 VDD2.n4 VDD2.n3 36.6162
R1307 VDD2.n7 VDD2.t1 1.88621
R1308 VDD2.n7 VDD2.t3 1.88621
R1309 VDD2.n5 VDD2.t6 1.88621
R1310 VDD2.n5 VDD2.t8 1.88621
R1311 VDD2.n2 VDD2.t9 1.88621
R1312 VDD2.n2 VDD2.t2 1.88621
R1313 VDD2.n0 VDD2.t5 1.88621
R1314 VDD2.n0 VDD2.t7 1.88621
R1315 VDD2.n6 VDD2.n4 0.810845
R1316 VDD2 VDD2.n6 0.261276
R1317 VDD2.n3 VDD2.n1 0.14774
C0 VTAIL VP 5.337029f
C1 VDD2 VN 5.47646f
C2 VDD1 VP 5.65329f
C3 VTAIL VN 5.32246f
C4 VDD2 VTAIL 13.5547f
C5 VDD1 VN 0.149252f
C6 VDD2 VDD1 0.916707f
C7 VDD1 VTAIL 13.5206f
C8 VN VP 5.18343f
C9 VDD2 VP 0.330345f
C10 VDD2 B 4.606632f
C11 VDD1 B 4.524714f
C12 VTAIL B 5.892758f
C13 VN B 8.89049f
C14 VP B 6.95894f
C15 VDD2.t0 B 2.36056f
C16 VDD2.t5 B 0.208873f
C17 VDD2.t7 B 0.208873f
C18 VDD2.n0 B 1.84828f
C19 VDD2.n1 B 0.621345f
C20 VDD2.t9 B 0.208873f
C21 VDD2.t2 B 0.208873f
C22 VDD2.n2 B 1.85098f
C23 VDD2.n3 B 1.77267f
C24 VDD2.t4 B 2.35655f
C25 VDD2.n4 B 2.24255f
C26 VDD2.t6 B 0.208873f
C27 VDD2.t8 B 0.208873f
C28 VDD2.n5 B 1.84828f
C29 VDD2.n6 B 0.290114f
C30 VDD2.t1 B 0.208873f
C31 VDD2.t3 B 0.208873f
C32 VDD2.n7 B 1.85095f
C33 VN.n0 B 0.044914f
C34 VN.t2 B 0.822324f
C35 VN.n1 B 0.347727f
C36 VN.t9 B 0.840121f
C37 VN.t4 B 0.822324f
C38 VN.n2 B 0.347518f
C39 VN.n3 B 0.321286f
C40 VN.n4 B 0.21846f
C41 VN.n5 B 0.059932f
C42 VN.t0 B 0.822324f
C43 VN.n6 B 0.337673f
C44 VN.n7 B 0.010192f
C45 VN.t7 B 0.822324f
C46 VN.n8 B 0.337396f
C47 VN.n9 B 0.034807f
C48 VN.n10 B 0.044914f
C49 VN.t1 B 0.822324f
C50 VN.n11 B 0.347727f
C51 VN.t3 B 0.822324f
C52 VN.t6 B 0.840121f
C53 VN.t8 B 0.822324f
C54 VN.n12 B 0.347518f
C55 VN.n13 B 0.321286f
C56 VN.n14 B 0.21846f
C57 VN.n15 B 0.059932f
C58 VN.n16 B 0.337673f
C59 VN.n17 B 0.010192f
C60 VN.t5 B 0.822324f
C61 VN.n18 B 0.337396f
C62 VN.n19 B 1.82378f
C63 VTAIL.t2 B 0.219573f
C64 VTAIL.t17 B 0.219573f
C65 VTAIL.n0 B 1.87238f
C66 VTAIL.n1 B 0.379656f
C67 VTAIL.t7 B 2.38826f
C68 VTAIL.n2 B 0.47493f
C69 VTAIL.t10 B 0.219573f
C70 VTAIL.t9 B 0.219573f
C71 VTAIL.n3 B 1.87238f
C72 VTAIL.n4 B 0.386455f
C73 VTAIL.t12 B 0.219573f
C74 VTAIL.t15 B 0.219573f
C75 VTAIL.n5 B 1.87238f
C76 VTAIL.n6 B 1.58685f
C77 VTAIL.t6 B 0.219573f
C78 VTAIL.t4 B 0.219573f
C79 VTAIL.n7 B 1.87239f
C80 VTAIL.n8 B 1.58685f
C81 VTAIL.t1 B 0.219573f
C82 VTAIL.t3 B 0.219573f
C83 VTAIL.n9 B 1.87239f
C84 VTAIL.n10 B 0.38645f
C85 VTAIL.t0 B 2.38826f
C86 VTAIL.n11 B 0.474924f
C87 VTAIL.t14 B 0.219573f
C88 VTAIL.t11 B 0.219573f
C89 VTAIL.n12 B 1.87239f
C90 VTAIL.n13 B 0.391963f
C91 VTAIL.t8 B 0.219573f
C92 VTAIL.t16 B 0.219573f
C93 VTAIL.n14 B 1.87239f
C94 VTAIL.n15 B 0.38645f
C95 VTAIL.t13 B 2.38826f
C96 VTAIL.n16 B 1.60072f
C97 VTAIL.t19 B 2.38826f
C98 VTAIL.n17 B 1.60072f
C99 VTAIL.t18 B 0.219573f
C100 VTAIL.t5 B 0.219573f
C101 VTAIL.n18 B 1.87238f
C102 VTAIL.n19 B 0.329671f
C103 VDD1.t5 B 2.36143f
C104 VDD1.t7 B 0.208949f
C105 VDD1.t9 B 0.208949f
C106 VDD1.n0 B 1.84896f
C107 VDD1.n1 B 0.626812f
C108 VDD1.t8 B 2.36143f
C109 VDD1.t0 B 0.208949f
C110 VDD1.t6 B 0.208949f
C111 VDD1.n2 B 1.84895f
C112 VDD1.n3 B 0.621572f
C113 VDD1.t2 B 0.208949f
C114 VDD1.t4 B 0.208949f
C115 VDD1.n4 B 1.85165f
C116 VDD1.n5 B 1.8483f
C117 VDD1.t1 B 0.208949f
C118 VDD1.t3 B 0.208949f
C119 VDD1.n6 B 1.84895f
C120 VDD1.n7 B 2.24459f
C121 VP.n0 B 0.045656f
C122 VP.t6 B 0.835902f
C123 VP.n1 B 0.353468f
C124 VP.n2 B 0.045656f
C125 VP.n3 B 0.045656f
C126 VP.t3 B 0.835902f
C127 VP.t0 B 0.835902f
C128 VP.n4 B 0.060922f
C129 VP.t8 B 0.835902f
C130 VP.n5 B 0.222067f
C131 VP.t5 B 0.835902f
C132 VP.t2 B 0.853992f
C133 VP.n6 B 0.32659f
C134 VP.n7 B 0.353256f
C135 VP.n8 B 0.353468f
C136 VP.n9 B 0.343249f
C137 VP.n10 B 0.01036f
C138 VP.n11 B 0.342967f
C139 VP.n12 B 1.82388f
C140 VP.n13 B 1.86384f
C141 VP.t4 B 0.835902f
C142 VP.n14 B 0.342967f
C143 VP.n15 B 0.01036f
C144 VP.t1 B 0.835902f
C145 VP.n16 B 0.343249f
C146 VP.n17 B 0.060922f
C147 VP.n18 B 0.060779f
C148 VP.n19 B 0.060922f
C149 VP.t7 B 0.835902f
C150 VP.n20 B 0.343249f
C151 VP.n21 B 0.01036f
C152 VP.t9 B 0.835902f
C153 VP.n22 B 0.342967f
C154 VP.n23 B 0.035381f
.ends

