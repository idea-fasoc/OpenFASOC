* NGSPICE file created from diff_pair_sample_0545.ext - technology: sky130A

.subckt diff_pair_sample_0545 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t19 VP.t0 VDD1.t7 B.t1 sky130_fd_pr__nfet_01v8 ad=2.41395 pd=14.96 as=2.41395 ps=14.96 w=14.63 l=1.54
X1 VDD1.t6 VP.t1 VTAIL.t18 B.t7 sky130_fd_pr__nfet_01v8 ad=5.7057 pd=30.04 as=2.41395 ps=14.96 w=14.63 l=1.54
X2 B.t23 B.t21 B.t22 B.t11 sky130_fd_pr__nfet_01v8 ad=5.7057 pd=30.04 as=0 ps=0 w=14.63 l=1.54
X3 VTAIL.t3 VN.t0 VDD2.t9 B.t3 sky130_fd_pr__nfet_01v8 ad=2.41395 pd=14.96 as=2.41395 ps=14.96 w=14.63 l=1.54
X4 VDD2.t8 VN.t1 VTAIL.t8 B.t8 sky130_fd_pr__nfet_01v8 ad=2.41395 pd=14.96 as=2.41395 ps=14.96 w=14.63 l=1.54
X5 VDD1.t3 VP.t2 VTAIL.t17 B.t8 sky130_fd_pr__nfet_01v8 ad=2.41395 pd=14.96 as=2.41395 ps=14.96 w=14.63 l=1.54
X6 VTAIL.t2 VN.t2 VDD2.t7 B.t2 sky130_fd_pr__nfet_01v8 ad=2.41395 pd=14.96 as=2.41395 ps=14.96 w=14.63 l=1.54
X7 B.t20 B.t18 B.t19 B.t15 sky130_fd_pr__nfet_01v8 ad=5.7057 pd=30.04 as=0 ps=0 w=14.63 l=1.54
X8 VTAIL.t16 VP.t3 VDD1.t2 B.t4 sky130_fd_pr__nfet_01v8 ad=2.41395 pd=14.96 as=2.41395 ps=14.96 w=14.63 l=1.54
X9 VDD2.t6 VN.t3 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.41395 pd=14.96 as=5.7057 ps=30.04 w=14.63 l=1.54
X10 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=5.7057 pd=30.04 as=0 ps=0 w=14.63 l=1.54
X11 VTAIL.t4 VN.t4 VDD2.t5 B.t4 sky130_fd_pr__nfet_01v8 ad=2.41395 pd=14.96 as=2.41395 ps=14.96 w=14.63 l=1.54
X12 VTAIL.t15 VP.t4 VDD1.t9 B.t3 sky130_fd_pr__nfet_01v8 ad=2.41395 pd=14.96 as=2.41395 ps=14.96 w=14.63 l=1.54
X13 VDD2.t4 VN.t5 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=5.7057 pd=30.04 as=2.41395 ps=14.96 w=14.63 l=1.54
X14 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=5.7057 pd=30.04 as=0 ps=0 w=14.63 l=1.54
X15 VDD2.t3 VN.t6 VTAIL.t9 B.t9 sky130_fd_pr__nfet_01v8 ad=5.7057 pd=30.04 as=2.41395 ps=14.96 w=14.63 l=1.54
X16 VTAIL.t14 VP.t5 VDD1.t8 B.t2 sky130_fd_pr__nfet_01v8 ad=2.41395 pd=14.96 as=2.41395 ps=14.96 w=14.63 l=1.54
X17 VDD1.t5 VP.t6 VTAIL.t13 B.t5 sky130_fd_pr__nfet_01v8 ad=2.41395 pd=14.96 as=2.41395 ps=14.96 w=14.63 l=1.54
X18 VDD2.t2 VN.t7 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=2.41395 pd=14.96 as=5.7057 ps=30.04 w=14.63 l=1.54
X19 VDD1.t4 VP.t7 VTAIL.t12 B.t9 sky130_fd_pr__nfet_01v8 ad=5.7057 pd=30.04 as=2.41395 ps=14.96 w=14.63 l=1.54
X20 VDD1.t1 VP.t8 VTAIL.t11 B.t0 sky130_fd_pr__nfet_01v8 ad=2.41395 pd=14.96 as=5.7057 ps=30.04 w=14.63 l=1.54
X21 VDD1.t0 VP.t9 VTAIL.t10 B.t6 sky130_fd_pr__nfet_01v8 ad=2.41395 pd=14.96 as=5.7057 ps=30.04 w=14.63 l=1.54
X22 VDD2.t1 VN.t8 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=2.41395 pd=14.96 as=2.41395 ps=14.96 w=14.63 l=1.54
X23 VTAIL.t1 VN.t9 VDD2.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=2.41395 pd=14.96 as=2.41395 ps=14.96 w=14.63 l=1.54
R0 VP.n15 VP.t1 263.575
R1 VP.n48 VP.t6 228.951
R2 VP.n35 VP.t7 228.951
R3 VP.n41 VP.t5 228.951
R4 VP.n54 VP.t0 228.951
R5 VP.n61 VP.t9 228.951
R6 VP.n20 VP.t2 228.951
R7 VP.n33 VP.t8 228.951
R8 VP.n26 VP.t4 228.951
R9 VP.n14 VP.t3 228.951
R10 VP.n36 VP.n35 174.024
R11 VP.n62 VP.n61 174.024
R12 VP.n34 VP.n33 174.024
R13 VP.n16 VP.n13 161.3
R14 VP.n18 VP.n17 161.3
R15 VP.n19 VP.n12 161.3
R16 VP.n21 VP.n20 161.3
R17 VP.n22 VP.n11 161.3
R18 VP.n24 VP.n23 161.3
R19 VP.n25 VP.n10 161.3
R20 VP.n28 VP.n27 161.3
R21 VP.n29 VP.n9 161.3
R22 VP.n31 VP.n30 161.3
R23 VP.n32 VP.n8 161.3
R24 VP.n60 VP.n0 161.3
R25 VP.n59 VP.n58 161.3
R26 VP.n57 VP.n1 161.3
R27 VP.n56 VP.n55 161.3
R28 VP.n53 VP.n2 161.3
R29 VP.n52 VP.n51 161.3
R30 VP.n50 VP.n3 161.3
R31 VP.n49 VP.n48 161.3
R32 VP.n47 VP.n4 161.3
R33 VP.n46 VP.n45 161.3
R34 VP.n44 VP.n5 161.3
R35 VP.n43 VP.n42 161.3
R36 VP.n40 VP.n6 161.3
R37 VP.n39 VP.n38 161.3
R38 VP.n37 VP.n7 161.3
R39 VP.n40 VP.n39 56.5193
R40 VP.n59 VP.n1 56.5193
R41 VP.n31 VP.n9 56.5193
R42 VP.n36 VP.n34 49.3073
R43 VP.n15 VP.n14 48.4385
R44 VP.n47 VP.n46 46.8066
R45 VP.n52 VP.n3 46.8066
R46 VP.n24 VP.n11 46.8066
R47 VP.n19 VP.n18 46.8066
R48 VP.n46 VP.n5 34.1802
R49 VP.n53 VP.n52 34.1802
R50 VP.n25 VP.n24 34.1802
R51 VP.n18 VP.n13 34.1802
R52 VP.n39 VP.n7 24.4675
R53 VP.n42 VP.n40 24.4675
R54 VP.n48 VP.n47 24.4675
R55 VP.n48 VP.n3 24.4675
R56 VP.n55 VP.n1 24.4675
R57 VP.n60 VP.n59 24.4675
R58 VP.n32 VP.n31 24.4675
R59 VP.n27 VP.n9 24.4675
R60 VP.n20 VP.n19 24.4675
R61 VP.n20 VP.n11 24.4675
R62 VP.n41 VP.n5 18.1061
R63 VP.n54 VP.n53 18.1061
R64 VP.n26 VP.n25 18.1061
R65 VP.n14 VP.n13 18.1061
R66 VP.n16 VP.n15 17.6128
R67 VP.n35 VP.n7 11.7447
R68 VP.n61 VP.n60 11.7447
R69 VP.n33 VP.n32 11.7447
R70 VP.n42 VP.n41 6.36192
R71 VP.n55 VP.n54 6.36192
R72 VP.n27 VP.n26 6.36192
R73 VP.n17 VP.n16 0.189894
R74 VP.n17 VP.n12 0.189894
R75 VP.n21 VP.n12 0.189894
R76 VP.n22 VP.n21 0.189894
R77 VP.n23 VP.n22 0.189894
R78 VP.n23 VP.n10 0.189894
R79 VP.n28 VP.n10 0.189894
R80 VP.n29 VP.n28 0.189894
R81 VP.n30 VP.n29 0.189894
R82 VP.n30 VP.n8 0.189894
R83 VP.n34 VP.n8 0.189894
R84 VP.n37 VP.n36 0.189894
R85 VP.n38 VP.n37 0.189894
R86 VP.n38 VP.n6 0.189894
R87 VP.n43 VP.n6 0.189894
R88 VP.n44 VP.n43 0.189894
R89 VP.n45 VP.n44 0.189894
R90 VP.n45 VP.n4 0.189894
R91 VP.n49 VP.n4 0.189894
R92 VP.n50 VP.n49 0.189894
R93 VP.n51 VP.n50 0.189894
R94 VP.n51 VP.n2 0.189894
R95 VP.n56 VP.n2 0.189894
R96 VP.n57 VP.n56 0.189894
R97 VP.n58 VP.n57 0.189894
R98 VP.n58 VP.n0 0.189894
R99 VP.n62 VP.n0 0.189894
R100 VP VP.n62 0.0516364
R101 VDD1.n76 VDD1.n0 289.615
R102 VDD1.n159 VDD1.n83 289.615
R103 VDD1.n77 VDD1.n76 185
R104 VDD1.n75 VDD1.n74 185
R105 VDD1.n73 VDD1.n3 185
R106 VDD1.n7 VDD1.n4 185
R107 VDD1.n68 VDD1.n67 185
R108 VDD1.n66 VDD1.n65 185
R109 VDD1.n9 VDD1.n8 185
R110 VDD1.n60 VDD1.n59 185
R111 VDD1.n58 VDD1.n57 185
R112 VDD1.n13 VDD1.n12 185
R113 VDD1.n52 VDD1.n51 185
R114 VDD1.n50 VDD1.n49 185
R115 VDD1.n17 VDD1.n16 185
R116 VDD1.n44 VDD1.n43 185
R117 VDD1.n42 VDD1.n41 185
R118 VDD1.n21 VDD1.n20 185
R119 VDD1.n36 VDD1.n35 185
R120 VDD1.n34 VDD1.n33 185
R121 VDD1.n25 VDD1.n24 185
R122 VDD1.n28 VDD1.n27 185
R123 VDD1.n110 VDD1.n109 185
R124 VDD1.n107 VDD1.n106 185
R125 VDD1.n116 VDD1.n115 185
R126 VDD1.n118 VDD1.n117 185
R127 VDD1.n103 VDD1.n102 185
R128 VDD1.n124 VDD1.n123 185
R129 VDD1.n126 VDD1.n125 185
R130 VDD1.n99 VDD1.n98 185
R131 VDD1.n132 VDD1.n131 185
R132 VDD1.n134 VDD1.n133 185
R133 VDD1.n95 VDD1.n94 185
R134 VDD1.n140 VDD1.n139 185
R135 VDD1.n142 VDD1.n141 185
R136 VDD1.n91 VDD1.n90 185
R137 VDD1.n148 VDD1.n147 185
R138 VDD1.n151 VDD1.n150 185
R139 VDD1.n149 VDD1.n87 185
R140 VDD1.n156 VDD1.n86 185
R141 VDD1.n158 VDD1.n157 185
R142 VDD1.n160 VDD1.n159 185
R143 VDD1.t6 VDD1.n26 147.659
R144 VDD1.t4 VDD1.n108 147.659
R145 VDD1.n76 VDD1.n75 104.615
R146 VDD1.n75 VDD1.n3 104.615
R147 VDD1.n7 VDD1.n3 104.615
R148 VDD1.n67 VDD1.n7 104.615
R149 VDD1.n67 VDD1.n66 104.615
R150 VDD1.n66 VDD1.n8 104.615
R151 VDD1.n59 VDD1.n8 104.615
R152 VDD1.n59 VDD1.n58 104.615
R153 VDD1.n58 VDD1.n12 104.615
R154 VDD1.n51 VDD1.n12 104.615
R155 VDD1.n51 VDD1.n50 104.615
R156 VDD1.n50 VDD1.n16 104.615
R157 VDD1.n43 VDD1.n16 104.615
R158 VDD1.n43 VDD1.n42 104.615
R159 VDD1.n42 VDD1.n20 104.615
R160 VDD1.n35 VDD1.n20 104.615
R161 VDD1.n35 VDD1.n34 104.615
R162 VDD1.n34 VDD1.n24 104.615
R163 VDD1.n27 VDD1.n24 104.615
R164 VDD1.n109 VDD1.n106 104.615
R165 VDD1.n116 VDD1.n106 104.615
R166 VDD1.n117 VDD1.n116 104.615
R167 VDD1.n117 VDD1.n102 104.615
R168 VDD1.n124 VDD1.n102 104.615
R169 VDD1.n125 VDD1.n124 104.615
R170 VDD1.n125 VDD1.n98 104.615
R171 VDD1.n132 VDD1.n98 104.615
R172 VDD1.n133 VDD1.n132 104.615
R173 VDD1.n133 VDD1.n94 104.615
R174 VDD1.n140 VDD1.n94 104.615
R175 VDD1.n141 VDD1.n140 104.615
R176 VDD1.n141 VDD1.n90 104.615
R177 VDD1.n148 VDD1.n90 104.615
R178 VDD1.n150 VDD1.n148 104.615
R179 VDD1.n150 VDD1.n149 104.615
R180 VDD1.n149 VDD1.n86 104.615
R181 VDD1.n158 VDD1.n86 104.615
R182 VDD1.n159 VDD1.n158 104.615
R183 VDD1.n167 VDD1.n166 61.8807
R184 VDD1.n82 VDD1.n81 60.7272
R185 VDD1.n169 VDD1.n168 60.727
R186 VDD1.n165 VDD1.n164 60.727
R187 VDD1.n27 VDD1.t6 52.3082
R188 VDD1.n109 VDD1.t4 52.3082
R189 VDD1.n82 VDD1.n80 50.2823
R190 VDD1.n165 VDD1.n163 50.2823
R191 VDD1.n169 VDD1.n167 45.3737
R192 VDD1.n28 VDD1.n26 15.6677
R193 VDD1.n110 VDD1.n108 15.6677
R194 VDD1.n74 VDD1.n73 13.1884
R195 VDD1.n157 VDD1.n156 13.1884
R196 VDD1.n77 VDD1.n2 12.8005
R197 VDD1.n72 VDD1.n4 12.8005
R198 VDD1.n29 VDD1.n25 12.8005
R199 VDD1.n111 VDD1.n107 12.8005
R200 VDD1.n155 VDD1.n87 12.8005
R201 VDD1.n160 VDD1.n85 12.8005
R202 VDD1.n78 VDD1.n0 12.0247
R203 VDD1.n69 VDD1.n68 12.0247
R204 VDD1.n33 VDD1.n32 12.0247
R205 VDD1.n115 VDD1.n114 12.0247
R206 VDD1.n152 VDD1.n151 12.0247
R207 VDD1.n161 VDD1.n83 12.0247
R208 VDD1.n65 VDD1.n6 11.249
R209 VDD1.n36 VDD1.n23 11.249
R210 VDD1.n118 VDD1.n105 11.249
R211 VDD1.n147 VDD1.n89 11.249
R212 VDD1.n64 VDD1.n9 10.4732
R213 VDD1.n37 VDD1.n21 10.4732
R214 VDD1.n119 VDD1.n103 10.4732
R215 VDD1.n146 VDD1.n91 10.4732
R216 VDD1.n61 VDD1.n60 9.69747
R217 VDD1.n41 VDD1.n40 9.69747
R218 VDD1.n123 VDD1.n122 9.69747
R219 VDD1.n143 VDD1.n142 9.69747
R220 VDD1.n80 VDD1.n79 9.45567
R221 VDD1.n163 VDD1.n162 9.45567
R222 VDD1.n54 VDD1.n53 9.3005
R223 VDD1.n56 VDD1.n55 9.3005
R224 VDD1.n11 VDD1.n10 9.3005
R225 VDD1.n62 VDD1.n61 9.3005
R226 VDD1.n64 VDD1.n63 9.3005
R227 VDD1.n6 VDD1.n5 9.3005
R228 VDD1.n70 VDD1.n69 9.3005
R229 VDD1.n72 VDD1.n71 9.3005
R230 VDD1.n79 VDD1.n78 9.3005
R231 VDD1.n2 VDD1.n1 9.3005
R232 VDD1.n15 VDD1.n14 9.3005
R233 VDD1.n48 VDD1.n47 9.3005
R234 VDD1.n46 VDD1.n45 9.3005
R235 VDD1.n19 VDD1.n18 9.3005
R236 VDD1.n40 VDD1.n39 9.3005
R237 VDD1.n38 VDD1.n37 9.3005
R238 VDD1.n23 VDD1.n22 9.3005
R239 VDD1.n32 VDD1.n31 9.3005
R240 VDD1.n30 VDD1.n29 9.3005
R241 VDD1.n162 VDD1.n161 9.3005
R242 VDD1.n85 VDD1.n84 9.3005
R243 VDD1.n130 VDD1.n129 9.3005
R244 VDD1.n128 VDD1.n127 9.3005
R245 VDD1.n101 VDD1.n100 9.3005
R246 VDD1.n122 VDD1.n121 9.3005
R247 VDD1.n120 VDD1.n119 9.3005
R248 VDD1.n105 VDD1.n104 9.3005
R249 VDD1.n114 VDD1.n113 9.3005
R250 VDD1.n112 VDD1.n111 9.3005
R251 VDD1.n97 VDD1.n96 9.3005
R252 VDD1.n136 VDD1.n135 9.3005
R253 VDD1.n138 VDD1.n137 9.3005
R254 VDD1.n93 VDD1.n92 9.3005
R255 VDD1.n144 VDD1.n143 9.3005
R256 VDD1.n146 VDD1.n145 9.3005
R257 VDD1.n89 VDD1.n88 9.3005
R258 VDD1.n153 VDD1.n152 9.3005
R259 VDD1.n155 VDD1.n154 9.3005
R260 VDD1.n57 VDD1.n11 8.92171
R261 VDD1.n44 VDD1.n19 8.92171
R262 VDD1.n126 VDD1.n101 8.92171
R263 VDD1.n139 VDD1.n93 8.92171
R264 VDD1.n56 VDD1.n13 8.14595
R265 VDD1.n45 VDD1.n17 8.14595
R266 VDD1.n127 VDD1.n99 8.14595
R267 VDD1.n138 VDD1.n95 8.14595
R268 VDD1.n53 VDD1.n52 7.3702
R269 VDD1.n49 VDD1.n48 7.3702
R270 VDD1.n131 VDD1.n130 7.3702
R271 VDD1.n135 VDD1.n134 7.3702
R272 VDD1.n52 VDD1.n15 6.59444
R273 VDD1.n49 VDD1.n15 6.59444
R274 VDD1.n131 VDD1.n97 6.59444
R275 VDD1.n134 VDD1.n97 6.59444
R276 VDD1.n53 VDD1.n13 5.81868
R277 VDD1.n48 VDD1.n17 5.81868
R278 VDD1.n130 VDD1.n99 5.81868
R279 VDD1.n135 VDD1.n95 5.81868
R280 VDD1.n57 VDD1.n56 5.04292
R281 VDD1.n45 VDD1.n44 5.04292
R282 VDD1.n127 VDD1.n126 5.04292
R283 VDD1.n139 VDD1.n138 5.04292
R284 VDD1.n30 VDD1.n26 4.38563
R285 VDD1.n112 VDD1.n108 4.38563
R286 VDD1.n60 VDD1.n11 4.26717
R287 VDD1.n41 VDD1.n19 4.26717
R288 VDD1.n123 VDD1.n101 4.26717
R289 VDD1.n142 VDD1.n93 4.26717
R290 VDD1.n61 VDD1.n9 3.49141
R291 VDD1.n40 VDD1.n21 3.49141
R292 VDD1.n122 VDD1.n103 3.49141
R293 VDD1.n143 VDD1.n91 3.49141
R294 VDD1.n65 VDD1.n64 2.71565
R295 VDD1.n37 VDD1.n36 2.71565
R296 VDD1.n119 VDD1.n118 2.71565
R297 VDD1.n147 VDD1.n146 2.71565
R298 VDD1.n80 VDD1.n0 1.93989
R299 VDD1.n68 VDD1.n6 1.93989
R300 VDD1.n33 VDD1.n23 1.93989
R301 VDD1.n115 VDD1.n105 1.93989
R302 VDD1.n151 VDD1.n89 1.93989
R303 VDD1.n163 VDD1.n83 1.93989
R304 VDD1.n168 VDD1.t9 1.35388
R305 VDD1.n168 VDD1.t1 1.35388
R306 VDD1.n81 VDD1.t2 1.35388
R307 VDD1.n81 VDD1.t3 1.35388
R308 VDD1.n166 VDD1.t7 1.35388
R309 VDD1.n166 VDD1.t0 1.35388
R310 VDD1.n164 VDD1.t8 1.35388
R311 VDD1.n164 VDD1.t5 1.35388
R312 VDD1.n78 VDD1.n77 1.16414
R313 VDD1.n69 VDD1.n4 1.16414
R314 VDD1.n32 VDD1.n25 1.16414
R315 VDD1.n114 VDD1.n107 1.16414
R316 VDD1.n152 VDD1.n87 1.16414
R317 VDD1.n161 VDD1.n160 1.16414
R318 VDD1 VDD1.n169 1.15136
R319 VDD1 VDD1.n82 0.461707
R320 VDD1.n74 VDD1.n2 0.388379
R321 VDD1.n73 VDD1.n72 0.388379
R322 VDD1.n29 VDD1.n28 0.388379
R323 VDD1.n111 VDD1.n110 0.388379
R324 VDD1.n156 VDD1.n155 0.388379
R325 VDD1.n157 VDD1.n85 0.388379
R326 VDD1.n167 VDD1.n165 0.348171
R327 VDD1.n79 VDD1.n1 0.155672
R328 VDD1.n71 VDD1.n1 0.155672
R329 VDD1.n71 VDD1.n70 0.155672
R330 VDD1.n70 VDD1.n5 0.155672
R331 VDD1.n63 VDD1.n5 0.155672
R332 VDD1.n63 VDD1.n62 0.155672
R333 VDD1.n62 VDD1.n10 0.155672
R334 VDD1.n55 VDD1.n10 0.155672
R335 VDD1.n55 VDD1.n54 0.155672
R336 VDD1.n54 VDD1.n14 0.155672
R337 VDD1.n47 VDD1.n14 0.155672
R338 VDD1.n47 VDD1.n46 0.155672
R339 VDD1.n46 VDD1.n18 0.155672
R340 VDD1.n39 VDD1.n18 0.155672
R341 VDD1.n39 VDD1.n38 0.155672
R342 VDD1.n38 VDD1.n22 0.155672
R343 VDD1.n31 VDD1.n22 0.155672
R344 VDD1.n31 VDD1.n30 0.155672
R345 VDD1.n113 VDD1.n112 0.155672
R346 VDD1.n113 VDD1.n104 0.155672
R347 VDD1.n120 VDD1.n104 0.155672
R348 VDD1.n121 VDD1.n120 0.155672
R349 VDD1.n121 VDD1.n100 0.155672
R350 VDD1.n128 VDD1.n100 0.155672
R351 VDD1.n129 VDD1.n128 0.155672
R352 VDD1.n129 VDD1.n96 0.155672
R353 VDD1.n136 VDD1.n96 0.155672
R354 VDD1.n137 VDD1.n136 0.155672
R355 VDD1.n137 VDD1.n92 0.155672
R356 VDD1.n144 VDD1.n92 0.155672
R357 VDD1.n145 VDD1.n144 0.155672
R358 VDD1.n145 VDD1.n88 0.155672
R359 VDD1.n153 VDD1.n88 0.155672
R360 VDD1.n154 VDD1.n153 0.155672
R361 VDD1.n154 VDD1.n84 0.155672
R362 VDD1.n162 VDD1.n84 0.155672
R363 VTAIL.n336 VTAIL.n260 289.615
R364 VTAIL.n78 VTAIL.n2 289.615
R365 VTAIL.n254 VTAIL.n178 289.615
R366 VTAIL.n168 VTAIL.n92 289.615
R367 VTAIL.n287 VTAIL.n286 185
R368 VTAIL.n284 VTAIL.n283 185
R369 VTAIL.n293 VTAIL.n292 185
R370 VTAIL.n295 VTAIL.n294 185
R371 VTAIL.n280 VTAIL.n279 185
R372 VTAIL.n301 VTAIL.n300 185
R373 VTAIL.n303 VTAIL.n302 185
R374 VTAIL.n276 VTAIL.n275 185
R375 VTAIL.n309 VTAIL.n308 185
R376 VTAIL.n311 VTAIL.n310 185
R377 VTAIL.n272 VTAIL.n271 185
R378 VTAIL.n317 VTAIL.n316 185
R379 VTAIL.n319 VTAIL.n318 185
R380 VTAIL.n268 VTAIL.n267 185
R381 VTAIL.n325 VTAIL.n324 185
R382 VTAIL.n328 VTAIL.n327 185
R383 VTAIL.n326 VTAIL.n264 185
R384 VTAIL.n333 VTAIL.n263 185
R385 VTAIL.n335 VTAIL.n334 185
R386 VTAIL.n337 VTAIL.n336 185
R387 VTAIL.n29 VTAIL.n28 185
R388 VTAIL.n26 VTAIL.n25 185
R389 VTAIL.n35 VTAIL.n34 185
R390 VTAIL.n37 VTAIL.n36 185
R391 VTAIL.n22 VTAIL.n21 185
R392 VTAIL.n43 VTAIL.n42 185
R393 VTAIL.n45 VTAIL.n44 185
R394 VTAIL.n18 VTAIL.n17 185
R395 VTAIL.n51 VTAIL.n50 185
R396 VTAIL.n53 VTAIL.n52 185
R397 VTAIL.n14 VTAIL.n13 185
R398 VTAIL.n59 VTAIL.n58 185
R399 VTAIL.n61 VTAIL.n60 185
R400 VTAIL.n10 VTAIL.n9 185
R401 VTAIL.n67 VTAIL.n66 185
R402 VTAIL.n70 VTAIL.n69 185
R403 VTAIL.n68 VTAIL.n6 185
R404 VTAIL.n75 VTAIL.n5 185
R405 VTAIL.n77 VTAIL.n76 185
R406 VTAIL.n79 VTAIL.n78 185
R407 VTAIL.n255 VTAIL.n254 185
R408 VTAIL.n253 VTAIL.n252 185
R409 VTAIL.n251 VTAIL.n181 185
R410 VTAIL.n185 VTAIL.n182 185
R411 VTAIL.n246 VTAIL.n245 185
R412 VTAIL.n244 VTAIL.n243 185
R413 VTAIL.n187 VTAIL.n186 185
R414 VTAIL.n238 VTAIL.n237 185
R415 VTAIL.n236 VTAIL.n235 185
R416 VTAIL.n191 VTAIL.n190 185
R417 VTAIL.n230 VTAIL.n229 185
R418 VTAIL.n228 VTAIL.n227 185
R419 VTAIL.n195 VTAIL.n194 185
R420 VTAIL.n222 VTAIL.n221 185
R421 VTAIL.n220 VTAIL.n219 185
R422 VTAIL.n199 VTAIL.n198 185
R423 VTAIL.n214 VTAIL.n213 185
R424 VTAIL.n212 VTAIL.n211 185
R425 VTAIL.n203 VTAIL.n202 185
R426 VTAIL.n206 VTAIL.n205 185
R427 VTAIL.n169 VTAIL.n168 185
R428 VTAIL.n167 VTAIL.n166 185
R429 VTAIL.n165 VTAIL.n95 185
R430 VTAIL.n99 VTAIL.n96 185
R431 VTAIL.n160 VTAIL.n159 185
R432 VTAIL.n158 VTAIL.n157 185
R433 VTAIL.n101 VTAIL.n100 185
R434 VTAIL.n152 VTAIL.n151 185
R435 VTAIL.n150 VTAIL.n149 185
R436 VTAIL.n105 VTAIL.n104 185
R437 VTAIL.n144 VTAIL.n143 185
R438 VTAIL.n142 VTAIL.n141 185
R439 VTAIL.n109 VTAIL.n108 185
R440 VTAIL.n136 VTAIL.n135 185
R441 VTAIL.n134 VTAIL.n133 185
R442 VTAIL.n113 VTAIL.n112 185
R443 VTAIL.n128 VTAIL.n127 185
R444 VTAIL.n126 VTAIL.n125 185
R445 VTAIL.n117 VTAIL.n116 185
R446 VTAIL.n120 VTAIL.n119 185
R447 VTAIL.t11 VTAIL.n204 147.659
R448 VTAIL.t6 VTAIL.n118 147.659
R449 VTAIL.t0 VTAIL.n285 147.659
R450 VTAIL.t10 VTAIL.n27 147.659
R451 VTAIL.n286 VTAIL.n283 104.615
R452 VTAIL.n293 VTAIL.n283 104.615
R453 VTAIL.n294 VTAIL.n293 104.615
R454 VTAIL.n294 VTAIL.n279 104.615
R455 VTAIL.n301 VTAIL.n279 104.615
R456 VTAIL.n302 VTAIL.n301 104.615
R457 VTAIL.n302 VTAIL.n275 104.615
R458 VTAIL.n309 VTAIL.n275 104.615
R459 VTAIL.n310 VTAIL.n309 104.615
R460 VTAIL.n310 VTAIL.n271 104.615
R461 VTAIL.n317 VTAIL.n271 104.615
R462 VTAIL.n318 VTAIL.n317 104.615
R463 VTAIL.n318 VTAIL.n267 104.615
R464 VTAIL.n325 VTAIL.n267 104.615
R465 VTAIL.n327 VTAIL.n325 104.615
R466 VTAIL.n327 VTAIL.n326 104.615
R467 VTAIL.n326 VTAIL.n263 104.615
R468 VTAIL.n335 VTAIL.n263 104.615
R469 VTAIL.n336 VTAIL.n335 104.615
R470 VTAIL.n28 VTAIL.n25 104.615
R471 VTAIL.n35 VTAIL.n25 104.615
R472 VTAIL.n36 VTAIL.n35 104.615
R473 VTAIL.n36 VTAIL.n21 104.615
R474 VTAIL.n43 VTAIL.n21 104.615
R475 VTAIL.n44 VTAIL.n43 104.615
R476 VTAIL.n44 VTAIL.n17 104.615
R477 VTAIL.n51 VTAIL.n17 104.615
R478 VTAIL.n52 VTAIL.n51 104.615
R479 VTAIL.n52 VTAIL.n13 104.615
R480 VTAIL.n59 VTAIL.n13 104.615
R481 VTAIL.n60 VTAIL.n59 104.615
R482 VTAIL.n60 VTAIL.n9 104.615
R483 VTAIL.n67 VTAIL.n9 104.615
R484 VTAIL.n69 VTAIL.n67 104.615
R485 VTAIL.n69 VTAIL.n68 104.615
R486 VTAIL.n68 VTAIL.n5 104.615
R487 VTAIL.n77 VTAIL.n5 104.615
R488 VTAIL.n78 VTAIL.n77 104.615
R489 VTAIL.n254 VTAIL.n253 104.615
R490 VTAIL.n253 VTAIL.n181 104.615
R491 VTAIL.n185 VTAIL.n181 104.615
R492 VTAIL.n245 VTAIL.n185 104.615
R493 VTAIL.n245 VTAIL.n244 104.615
R494 VTAIL.n244 VTAIL.n186 104.615
R495 VTAIL.n237 VTAIL.n186 104.615
R496 VTAIL.n237 VTAIL.n236 104.615
R497 VTAIL.n236 VTAIL.n190 104.615
R498 VTAIL.n229 VTAIL.n190 104.615
R499 VTAIL.n229 VTAIL.n228 104.615
R500 VTAIL.n228 VTAIL.n194 104.615
R501 VTAIL.n221 VTAIL.n194 104.615
R502 VTAIL.n221 VTAIL.n220 104.615
R503 VTAIL.n220 VTAIL.n198 104.615
R504 VTAIL.n213 VTAIL.n198 104.615
R505 VTAIL.n213 VTAIL.n212 104.615
R506 VTAIL.n212 VTAIL.n202 104.615
R507 VTAIL.n205 VTAIL.n202 104.615
R508 VTAIL.n168 VTAIL.n167 104.615
R509 VTAIL.n167 VTAIL.n95 104.615
R510 VTAIL.n99 VTAIL.n95 104.615
R511 VTAIL.n159 VTAIL.n99 104.615
R512 VTAIL.n159 VTAIL.n158 104.615
R513 VTAIL.n158 VTAIL.n100 104.615
R514 VTAIL.n151 VTAIL.n100 104.615
R515 VTAIL.n151 VTAIL.n150 104.615
R516 VTAIL.n150 VTAIL.n104 104.615
R517 VTAIL.n143 VTAIL.n104 104.615
R518 VTAIL.n143 VTAIL.n142 104.615
R519 VTAIL.n142 VTAIL.n108 104.615
R520 VTAIL.n135 VTAIL.n108 104.615
R521 VTAIL.n135 VTAIL.n134 104.615
R522 VTAIL.n134 VTAIL.n112 104.615
R523 VTAIL.n127 VTAIL.n112 104.615
R524 VTAIL.n127 VTAIL.n126 104.615
R525 VTAIL.n126 VTAIL.n116 104.615
R526 VTAIL.n119 VTAIL.n116 104.615
R527 VTAIL.n286 VTAIL.t0 52.3082
R528 VTAIL.n28 VTAIL.t10 52.3082
R529 VTAIL.n205 VTAIL.t11 52.3082
R530 VTAIL.n119 VTAIL.t6 52.3082
R531 VTAIL.n177 VTAIL.n176 44.0484
R532 VTAIL.n175 VTAIL.n174 44.0484
R533 VTAIL.n91 VTAIL.n90 44.0484
R534 VTAIL.n89 VTAIL.n88 44.0484
R535 VTAIL.n343 VTAIL.n342 44.0482
R536 VTAIL.n1 VTAIL.n0 44.0482
R537 VTAIL.n85 VTAIL.n84 44.0482
R538 VTAIL.n87 VTAIL.n86 44.0482
R539 VTAIL.n341 VTAIL.n340 31.9914
R540 VTAIL.n83 VTAIL.n82 31.9914
R541 VTAIL.n259 VTAIL.n258 31.9914
R542 VTAIL.n173 VTAIL.n172 31.9914
R543 VTAIL.n89 VTAIL.n87 28.2031
R544 VTAIL.n341 VTAIL.n259 26.591
R545 VTAIL.n287 VTAIL.n285 15.6677
R546 VTAIL.n29 VTAIL.n27 15.6677
R547 VTAIL.n206 VTAIL.n204 15.6677
R548 VTAIL.n120 VTAIL.n118 15.6677
R549 VTAIL.n334 VTAIL.n333 13.1884
R550 VTAIL.n76 VTAIL.n75 13.1884
R551 VTAIL.n252 VTAIL.n251 13.1884
R552 VTAIL.n166 VTAIL.n165 13.1884
R553 VTAIL.n288 VTAIL.n284 12.8005
R554 VTAIL.n332 VTAIL.n264 12.8005
R555 VTAIL.n337 VTAIL.n262 12.8005
R556 VTAIL.n30 VTAIL.n26 12.8005
R557 VTAIL.n74 VTAIL.n6 12.8005
R558 VTAIL.n79 VTAIL.n4 12.8005
R559 VTAIL.n255 VTAIL.n180 12.8005
R560 VTAIL.n250 VTAIL.n182 12.8005
R561 VTAIL.n207 VTAIL.n203 12.8005
R562 VTAIL.n169 VTAIL.n94 12.8005
R563 VTAIL.n164 VTAIL.n96 12.8005
R564 VTAIL.n121 VTAIL.n117 12.8005
R565 VTAIL.n292 VTAIL.n291 12.0247
R566 VTAIL.n329 VTAIL.n328 12.0247
R567 VTAIL.n338 VTAIL.n260 12.0247
R568 VTAIL.n34 VTAIL.n33 12.0247
R569 VTAIL.n71 VTAIL.n70 12.0247
R570 VTAIL.n80 VTAIL.n2 12.0247
R571 VTAIL.n256 VTAIL.n178 12.0247
R572 VTAIL.n247 VTAIL.n246 12.0247
R573 VTAIL.n211 VTAIL.n210 12.0247
R574 VTAIL.n170 VTAIL.n92 12.0247
R575 VTAIL.n161 VTAIL.n160 12.0247
R576 VTAIL.n125 VTAIL.n124 12.0247
R577 VTAIL.n295 VTAIL.n282 11.249
R578 VTAIL.n324 VTAIL.n266 11.249
R579 VTAIL.n37 VTAIL.n24 11.249
R580 VTAIL.n66 VTAIL.n8 11.249
R581 VTAIL.n243 VTAIL.n184 11.249
R582 VTAIL.n214 VTAIL.n201 11.249
R583 VTAIL.n157 VTAIL.n98 11.249
R584 VTAIL.n128 VTAIL.n115 11.249
R585 VTAIL.n296 VTAIL.n280 10.4732
R586 VTAIL.n323 VTAIL.n268 10.4732
R587 VTAIL.n38 VTAIL.n22 10.4732
R588 VTAIL.n65 VTAIL.n10 10.4732
R589 VTAIL.n242 VTAIL.n187 10.4732
R590 VTAIL.n215 VTAIL.n199 10.4732
R591 VTAIL.n156 VTAIL.n101 10.4732
R592 VTAIL.n129 VTAIL.n113 10.4732
R593 VTAIL.n300 VTAIL.n299 9.69747
R594 VTAIL.n320 VTAIL.n319 9.69747
R595 VTAIL.n42 VTAIL.n41 9.69747
R596 VTAIL.n62 VTAIL.n61 9.69747
R597 VTAIL.n239 VTAIL.n238 9.69747
R598 VTAIL.n219 VTAIL.n218 9.69747
R599 VTAIL.n153 VTAIL.n152 9.69747
R600 VTAIL.n133 VTAIL.n132 9.69747
R601 VTAIL.n340 VTAIL.n339 9.45567
R602 VTAIL.n82 VTAIL.n81 9.45567
R603 VTAIL.n258 VTAIL.n257 9.45567
R604 VTAIL.n172 VTAIL.n171 9.45567
R605 VTAIL.n339 VTAIL.n338 9.3005
R606 VTAIL.n262 VTAIL.n261 9.3005
R607 VTAIL.n307 VTAIL.n306 9.3005
R608 VTAIL.n305 VTAIL.n304 9.3005
R609 VTAIL.n278 VTAIL.n277 9.3005
R610 VTAIL.n299 VTAIL.n298 9.3005
R611 VTAIL.n297 VTAIL.n296 9.3005
R612 VTAIL.n282 VTAIL.n281 9.3005
R613 VTAIL.n291 VTAIL.n290 9.3005
R614 VTAIL.n289 VTAIL.n288 9.3005
R615 VTAIL.n274 VTAIL.n273 9.3005
R616 VTAIL.n313 VTAIL.n312 9.3005
R617 VTAIL.n315 VTAIL.n314 9.3005
R618 VTAIL.n270 VTAIL.n269 9.3005
R619 VTAIL.n321 VTAIL.n320 9.3005
R620 VTAIL.n323 VTAIL.n322 9.3005
R621 VTAIL.n266 VTAIL.n265 9.3005
R622 VTAIL.n330 VTAIL.n329 9.3005
R623 VTAIL.n332 VTAIL.n331 9.3005
R624 VTAIL.n81 VTAIL.n80 9.3005
R625 VTAIL.n4 VTAIL.n3 9.3005
R626 VTAIL.n49 VTAIL.n48 9.3005
R627 VTAIL.n47 VTAIL.n46 9.3005
R628 VTAIL.n20 VTAIL.n19 9.3005
R629 VTAIL.n41 VTAIL.n40 9.3005
R630 VTAIL.n39 VTAIL.n38 9.3005
R631 VTAIL.n24 VTAIL.n23 9.3005
R632 VTAIL.n33 VTAIL.n32 9.3005
R633 VTAIL.n31 VTAIL.n30 9.3005
R634 VTAIL.n16 VTAIL.n15 9.3005
R635 VTAIL.n55 VTAIL.n54 9.3005
R636 VTAIL.n57 VTAIL.n56 9.3005
R637 VTAIL.n12 VTAIL.n11 9.3005
R638 VTAIL.n63 VTAIL.n62 9.3005
R639 VTAIL.n65 VTAIL.n64 9.3005
R640 VTAIL.n8 VTAIL.n7 9.3005
R641 VTAIL.n72 VTAIL.n71 9.3005
R642 VTAIL.n74 VTAIL.n73 9.3005
R643 VTAIL.n232 VTAIL.n231 9.3005
R644 VTAIL.n234 VTAIL.n233 9.3005
R645 VTAIL.n189 VTAIL.n188 9.3005
R646 VTAIL.n240 VTAIL.n239 9.3005
R647 VTAIL.n242 VTAIL.n241 9.3005
R648 VTAIL.n184 VTAIL.n183 9.3005
R649 VTAIL.n248 VTAIL.n247 9.3005
R650 VTAIL.n250 VTAIL.n249 9.3005
R651 VTAIL.n257 VTAIL.n256 9.3005
R652 VTAIL.n180 VTAIL.n179 9.3005
R653 VTAIL.n193 VTAIL.n192 9.3005
R654 VTAIL.n226 VTAIL.n225 9.3005
R655 VTAIL.n224 VTAIL.n223 9.3005
R656 VTAIL.n197 VTAIL.n196 9.3005
R657 VTAIL.n218 VTAIL.n217 9.3005
R658 VTAIL.n216 VTAIL.n215 9.3005
R659 VTAIL.n201 VTAIL.n200 9.3005
R660 VTAIL.n210 VTAIL.n209 9.3005
R661 VTAIL.n208 VTAIL.n207 9.3005
R662 VTAIL.n146 VTAIL.n145 9.3005
R663 VTAIL.n148 VTAIL.n147 9.3005
R664 VTAIL.n103 VTAIL.n102 9.3005
R665 VTAIL.n154 VTAIL.n153 9.3005
R666 VTAIL.n156 VTAIL.n155 9.3005
R667 VTAIL.n98 VTAIL.n97 9.3005
R668 VTAIL.n162 VTAIL.n161 9.3005
R669 VTAIL.n164 VTAIL.n163 9.3005
R670 VTAIL.n171 VTAIL.n170 9.3005
R671 VTAIL.n94 VTAIL.n93 9.3005
R672 VTAIL.n107 VTAIL.n106 9.3005
R673 VTAIL.n140 VTAIL.n139 9.3005
R674 VTAIL.n138 VTAIL.n137 9.3005
R675 VTAIL.n111 VTAIL.n110 9.3005
R676 VTAIL.n132 VTAIL.n131 9.3005
R677 VTAIL.n130 VTAIL.n129 9.3005
R678 VTAIL.n115 VTAIL.n114 9.3005
R679 VTAIL.n124 VTAIL.n123 9.3005
R680 VTAIL.n122 VTAIL.n121 9.3005
R681 VTAIL.n303 VTAIL.n278 8.92171
R682 VTAIL.n316 VTAIL.n270 8.92171
R683 VTAIL.n45 VTAIL.n20 8.92171
R684 VTAIL.n58 VTAIL.n12 8.92171
R685 VTAIL.n235 VTAIL.n189 8.92171
R686 VTAIL.n222 VTAIL.n197 8.92171
R687 VTAIL.n149 VTAIL.n103 8.92171
R688 VTAIL.n136 VTAIL.n111 8.92171
R689 VTAIL.n304 VTAIL.n276 8.14595
R690 VTAIL.n315 VTAIL.n272 8.14595
R691 VTAIL.n46 VTAIL.n18 8.14595
R692 VTAIL.n57 VTAIL.n14 8.14595
R693 VTAIL.n234 VTAIL.n191 8.14595
R694 VTAIL.n223 VTAIL.n195 8.14595
R695 VTAIL.n148 VTAIL.n105 8.14595
R696 VTAIL.n137 VTAIL.n109 8.14595
R697 VTAIL.n308 VTAIL.n307 7.3702
R698 VTAIL.n312 VTAIL.n311 7.3702
R699 VTAIL.n50 VTAIL.n49 7.3702
R700 VTAIL.n54 VTAIL.n53 7.3702
R701 VTAIL.n231 VTAIL.n230 7.3702
R702 VTAIL.n227 VTAIL.n226 7.3702
R703 VTAIL.n145 VTAIL.n144 7.3702
R704 VTAIL.n141 VTAIL.n140 7.3702
R705 VTAIL.n308 VTAIL.n274 6.59444
R706 VTAIL.n311 VTAIL.n274 6.59444
R707 VTAIL.n50 VTAIL.n16 6.59444
R708 VTAIL.n53 VTAIL.n16 6.59444
R709 VTAIL.n230 VTAIL.n193 6.59444
R710 VTAIL.n227 VTAIL.n193 6.59444
R711 VTAIL.n144 VTAIL.n107 6.59444
R712 VTAIL.n141 VTAIL.n107 6.59444
R713 VTAIL.n307 VTAIL.n276 5.81868
R714 VTAIL.n312 VTAIL.n272 5.81868
R715 VTAIL.n49 VTAIL.n18 5.81868
R716 VTAIL.n54 VTAIL.n14 5.81868
R717 VTAIL.n231 VTAIL.n191 5.81868
R718 VTAIL.n226 VTAIL.n195 5.81868
R719 VTAIL.n145 VTAIL.n105 5.81868
R720 VTAIL.n140 VTAIL.n109 5.81868
R721 VTAIL.n304 VTAIL.n303 5.04292
R722 VTAIL.n316 VTAIL.n315 5.04292
R723 VTAIL.n46 VTAIL.n45 5.04292
R724 VTAIL.n58 VTAIL.n57 5.04292
R725 VTAIL.n235 VTAIL.n234 5.04292
R726 VTAIL.n223 VTAIL.n222 5.04292
R727 VTAIL.n149 VTAIL.n148 5.04292
R728 VTAIL.n137 VTAIL.n136 5.04292
R729 VTAIL.n208 VTAIL.n204 4.38563
R730 VTAIL.n122 VTAIL.n118 4.38563
R731 VTAIL.n289 VTAIL.n285 4.38563
R732 VTAIL.n31 VTAIL.n27 4.38563
R733 VTAIL.n300 VTAIL.n278 4.26717
R734 VTAIL.n319 VTAIL.n270 4.26717
R735 VTAIL.n42 VTAIL.n20 4.26717
R736 VTAIL.n61 VTAIL.n12 4.26717
R737 VTAIL.n238 VTAIL.n189 4.26717
R738 VTAIL.n219 VTAIL.n197 4.26717
R739 VTAIL.n152 VTAIL.n103 4.26717
R740 VTAIL.n133 VTAIL.n111 4.26717
R741 VTAIL.n299 VTAIL.n280 3.49141
R742 VTAIL.n320 VTAIL.n268 3.49141
R743 VTAIL.n41 VTAIL.n22 3.49141
R744 VTAIL.n62 VTAIL.n10 3.49141
R745 VTAIL.n239 VTAIL.n187 3.49141
R746 VTAIL.n218 VTAIL.n199 3.49141
R747 VTAIL.n153 VTAIL.n101 3.49141
R748 VTAIL.n132 VTAIL.n113 3.49141
R749 VTAIL.n296 VTAIL.n295 2.71565
R750 VTAIL.n324 VTAIL.n323 2.71565
R751 VTAIL.n38 VTAIL.n37 2.71565
R752 VTAIL.n66 VTAIL.n65 2.71565
R753 VTAIL.n243 VTAIL.n242 2.71565
R754 VTAIL.n215 VTAIL.n214 2.71565
R755 VTAIL.n157 VTAIL.n156 2.71565
R756 VTAIL.n129 VTAIL.n128 2.71565
R757 VTAIL.n292 VTAIL.n282 1.93989
R758 VTAIL.n328 VTAIL.n266 1.93989
R759 VTAIL.n340 VTAIL.n260 1.93989
R760 VTAIL.n34 VTAIL.n24 1.93989
R761 VTAIL.n70 VTAIL.n8 1.93989
R762 VTAIL.n82 VTAIL.n2 1.93989
R763 VTAIL.n258 VTAIL.n178 1.93989
R764 VTAIL.n246 VTAIL.n184 1.93989
R765 VTAIL.n211 VTAIL.n201 1.93989
R766 VTAIL.n172 VTAIL.n92 1.93989
R767 VTAIL.n160 VTAIL.n98 1.93989
R768 VTAIL.n125 VTAIL.n115 1.93989
R769 VTAIL.n91 VTAIL.n89 1.61257
R770 VTAIL.n173 VTAIL.n91 1.61257
R771 VTAIL.n177 VTAIL.n175 1.61257
R772 VTAIL.n259 VTAIL.n177 1.61257
R773 VTAIL.n87 VTAIL.n85 1.61257
R774 VTAIL.n85 VTAIL.n83 1.61257
R775 VTAIL.n343 VTAIL.n341 1.61257
R776 VTAIL.n342 VTAIL.t8 1.35388
R777 VTAIL.n342 VTAIL.t3 1.35388
R778 VTAIL.n0 VTAIL.t7 1.35388
R779 VTAIL.n0 VTAIL.t4 1.35388
R780 VTAIL.n84 VTAIL.t13 1.35388
R781 VTAIL.n84 VTAIL.t19 1.35388
R782 VTAIL.n86 VTAIL.t12 1.35388
R783 VTAIL.n86 VTAIL.t14 1.35388
R784 VTAIL.n176 VTAIL.t17 1.35388
R785 VTAIL.n176 VTAIL.t15 1.35388
R786 VTAIL.n174 VTAIL.t18 1.35388
R787 VTAIL.n174 VTAIL.t16 1.35388
R788 VTAIL.n90 VTAIL.t5 1.35388
R789 VTAIL.n90 VTAIL.t1 1.35388
R790 VTAIL.n88 VTAIL.t9 1.35388
R791 VTAIL.n88 VTAIL.t2 1.35388
R792 VTAIL.n175 VTAIL.n173 1.27636
R793 VTAIL.n83 VTAIL.n1 1.27636
R794 VTAIL VTAIL.n1 1.26774
R795 VTAIL.n291 VTAIL.n284 1.16414
R796 VTAIL.n329 VTAIL.n264 1.16414
R797 VTAIL.n338 VTAIL.n337 1.16414
R798 VTAIL.n33 VTAIL.n26 1.16414
R799 VTAIL.n71 VTAIL.n6 1.16414
R800 VTAIL.n80 VTAIL.n79 1.16414
R801 VTAIL.n256 VTAIL.n255 1.16414
R802 VTAIL.n247 VTAIL.n182 1.16414
R803 VTAIL.n210 VTAIL.n203 1.16414
R804 VTAIL.n170 VTAIL.n169 1.16414
R805 VTAIL.n161 VTAIL.n96 1.16414
R806 VTAIL.n124 VTAIL.n117 1.16414
R807 VTAIL.n288 VTAIL.n287 0.388379
R808 VTAIL.n333 VTAIL.n332 0.388379
R809 VTAIL.n334 VTAIL.n262 0.388379
R810 VTAIL.n30 VTAIL.n29 0.388379
R811 VTAIL.n75 VTAIL.n74 0.388379
R812 VTAIL.n76 VTAIL.n4 0.388379
R813 VTAIL.n252 VTAIL.n180 0.388379
R814 VTAIL.n251 VTAIL.n250 0.388379
R815 VTAIL.n207 VTAIL.n206 0.388379
R816 VTAIL.n166 VTAIL.n94 0.388379
R817 VTAIL.n165 VTAIL.n164 0.388379
R818 VTAIL.n121 VTAIL.n120 0.388379
R819 VTAIL VTAIL.n343 0.345328
R820 VTAIL.n290 VTAIL.n289 0.155672
R821 VTAIL.n290 VTAIL.n281 0.155672
R822 VTAIL.n297 VTAIL.n281 0.155672
R823 VTAIL.n298 VTAIL.n297 0.155672
R824 VTAIL.n298 VTAIL.n277 0.155672
R825 VTAIL.n305 VTAIL.n277 0.155672
R826 VTAIL.n306 VTAIL.n305 0.155672
R827 VTAIL.n306 VTAIL.n273 0.155672
R828 VTAIL.n313 VTAIL.n273 0.155672
R829 VTAIL.n314 VTAIL.n313 0.155672
R830 VTAIL.n314 VTAIL.n269 0.155672
R831 VTAIL.n321 VTAIL.n269 0.155672
R832 VTAIL.n322 VTAIL.n321 0.155672
R833 VTAIL.n322 VTAIL.n265 0.155672
R834 VTAIL.n330 VTAIL.n265 0.155672
R835 VTAIL.n331 VTAIL.n330 0.155672
R836 VTAIL.n331 VTAIL.n261 0.155672
R837 VTAIL.n339 VTAIL.n261 0.155672
R838 VTAIL.n32 VTAIL.n31 0.155672
R839 VTAIL.n32 VTAIL.n23 0.155672
R840 VTAIL.n39 VTAIL.n23 0.155672
R841 VTAIL.n40 VTAIL.n39 0.155672
R842 VTAIL.n40 VTAIL.n19 0.155672
R843 VTAIL.n47 VTAIL.n19 0.155672
R844 VTAIL.n48 VTAIL.n47 0.155672
R845 VTAIL.n48 VTAIL.n15 0.155672
R846 VTAIL.n55 VTAIL.n15 0.155672
R847 VTAIL.n56 VTAIL.n55 0.155672
R848 VTAIL.n56 VTAIL.n11 0.155672
R849 VTAIL.n63 VTAIL.n11 0.155672
R850 VTAIL.n64 VTAIL.n63 0.155672
R851 VTAIL.n64 VTAIL.n7 0.155672
R852 VTAIL.n72 VTAIL.n7 0.155672
R853 VTAIL.n73 VTAIL.n72 0.155672
R854 VTAIL.n73 VTAIL.n3 0.155672
R855 VTAIL.n81 VTAIL.n3 0.155672
R856 VTAIL.n257 VTAIL.n179 0.155672
R857 VTAIL.n249 VTAIL.n179 0.155672
R858 VTAIL.n249 VTAIL.n248 0.155672
R859 VTAIL.n248 VTAIL.n183 0.155672
R860 VTAIL.n241 VTAIL.n183 0.155672
R861 VTAIL.n241 VTAIL.n240 0.155672
R862 VTAIL.n240 VTAIL.n188 0.155672
R863 VTAIL.n233 VTAIL.n188 0.155672
R864 VTAIL.n233 VTAIL.n232 0.155672
R865 VTAIL.n232 VTAIL.n192 0.155672
R866 VTAIL.n225 VTAIL.n192 0.155672
R867 VTAIL.n225 VTAIL.n224 0.155672
R868 VTAIL.n224 VTAIL.n196 0.155672
R869 VTAIL.n217 VTAIL.n196 0.155672
R870 VTAIL.n217 VTAIL.n216 0.155672
R871 VTAIL.n216 VTAIL.n200 0.155672
R872 VTAIL.n209 VTAIL.n200 0.155672
R873 VTAIL.n209 VTAIL.n208 0.155672
R874 VTAIL.n171 VTAIL.n93 0.155672
R875 VTAIL.n163 VTAIL.n93 0.155672
R876 VTAIL.n163 VTAIL.n162 0.155672
R877 VTAIL.n162 VTAIL.n97 0.155672
R878 VTAIL.n155 VTAIL.n97 0.155672
R879 VTAIL.n155 VTAIL.n154 0.155672
R880 VTAIL.n154 VTAIL.n102 0.155672
R881 VTAIL.n147 VTAIL.n102 0.155672
R882 VTAIL.n147 VTAIL.n146 0.155672
R883 VTAIL.n146 VTAIL.n106 0.155672
R884 VTAIL.n139 VTAIL.n106 0.155672
R885 VTAIL.n139 VTAIL.n138 0.155672
R886 VTAIL.n138 VTAIL.n110 0.155672
R887 VTAIL.n131 VTAIL.n110 0.155672
R888 VTAIL.n131 VTAIL.n130 0.155672
R889 VTAIL.n130 VTAIL.n114 0.155672
R890 VTAIL.n123 VTAIL.n114 0.155672
R891 VTAIL.n123 VTAIL.n122 0.155672
R892 B.n881 B.n880 585
R893 B.n349 B.n130 585
R894 B.n348 B.n347 585
R895 B.n346 B.n345 585
R896 B.n344 B.n343 585
R897 B.n342 B.n341 585
R898 B.n340 B.n339 585
R899 B.n338 B.n337 585
R900 B.n336 B.n335 585
R901 B.n334 B.n333 585
R902 B.n332 B.n331 585
R903 B.n330 B.n329 585
R904 B.n328 B.n327 585
R905 B.n326 B.n325 585
R906 B.n324 B.n323 585
R907 B.n322 B.n321 585
R908 B.n320 B.n319 585
R909 B.n318 B.n317 585
R910 B.n316 B.n315 585
R911 B.n314 B.n313 585
R912 B.n312 B.n311 585
R913 B.n310 B.n309 585
R914 B.n308 B.n307 585
R915 B.n306 B.n305 585
R916 B.n304 B.n303 585
R917 B.n302 B.n301 585
R918 B.n300 B.n299 585
R919 B.n298 B.n297 585
R920 B.n296 B.n295 585
R921 B.n294 B.n293 585
R922 B.n292 B.n291 585
R923 B.n290 B.n289 585
R924 B.n288 B.n287 585
R925 B.n286 B.n285 585
R926 B.n284 B.n283 585
R927 B.n282 B.n281 585
R928 B.n280 B.n279 585
R929 B.n278 B.n277 585
R930 B.n276 B.n275 585
R931 B.n274 B.n273 585
R932 B.n272 B.n271 585
R933 B.n270 B.n269 585
R934 B.n268 B.n267 585
R935 B.n266 B.n265 585
R936 B.n264 B.n263 585
R937 B.n262 B.n261 585
R938 B.n260 B.n259 585
R939 B.n258 B.n257 585
R940 B.n256 B.n255 585
R941 B.n253 B.n252 585
R942 B.n251 B.n250 585
R943 B.n249 B.n248 585
R944 B.n247 B.n246 585
R945 B.n245 B.n244 585
R946 B.n243 B.n242 585
R947 B.n241 B.n240 585
R948 B.n239 B.n238 585
R949 B.n237 B.n236 585
R950 B.n235 B.n234 585
R951 B.n232 B.n231 585
R952 B.n230 B.n229 585
R953 B.n228 B.n227 585
R954 B.n226 B.n225 585
R955 B.n224 B.n223 585
R956 B.n222 B.n221 585
R957 B.n220 B.n219 585
R958 B.n218 B.n217 585
R959 B.n216 B.n215 585
R960 B.n214 B.n213 585
R961 B.n212 B.n211 585
R962 B.n210 B.n209 585
R963 B.n208 B.n207 585
R964 B.n206 B.n205 585
R965 B.n204 B.n203 585
R966 B.n202 B.n201 585
R967 B.n200 B.n199 585
R968 B.n198 B.n197 585
R969 B.n196 B.n195 585
R970 B.n194 B.n193 585
R971 B.n192 B.n191 585
R972 B.n190 B.n189 585
R973 B.n188 B.n187 585
R974 B.n186 B.n185 585
R975 B.n184 B.n183 585
R976 B.n182 B.n181 585
R977 B.n180 B.n179 585
R978 B.n178 B.n177 585
R979 B.n176 B.n175 585
R980 B.n174 B.n173 585
R981 B.n172 B.n171 585
R982 B.n170 B.n169 585
R983 B.n168 B.n167 585
R984 B.n166 B.n165 585
R985 B.n164 B.n163 585
R986 B.n162 B.n161 585
R987 B.n160 B.n159 585
R988 B.n158 B.n157 585
R989 B.n156 B.n155 585
R990 B.n154 B.n153 585
R991 B.n152 B.n151 585
R992 B.n150 B.n149 585
R993 B.n148 B.n147 585
R994 B.n146 B.n145 585
R995 B.n144 B.n143 585
R996 B.n142 B.n141 585
R997 B.n140 B.n139 585
R998 B.n138 B.n137 585
R999 B.n136 B.n135 585
R1000 B.n879 B.n76 585
R1001 B.n884 B.n76 585
R1002 B.n878 B.n75 585
R1003 B.n885 B.n75 585
R1004 B.n877 B.n876 585
R1005 B.n876 B.n71 585
R1006 B.n875 B.n70 585
R1007 B.n891 B.n70 585
R1008 B.n874 B.n69 585
R1009 B.n892 B.n69 585
R1010 B.n873 B.n68 585
R1011 B.n893 B.n68 585
R1012 B.n872 B.n871 585
R1013 B.n871 B.n64 585
R1014 B.n870 B.n63 585
R1015 B.n899 B.n63 585
R1016 B.n869 B.n62 585
R1017 B.n900 B.n62 585
R1018 B.n868 B.n61 585
R1019 B.n901 B.n61 585
R1020 B.n867 B.n866 585
R1021 B.n866 B.n57 585
R1022 B.n865 B.n56 585
R1023 B.n907 B.n56 585
R1024 B.n864 B.n55 585
R1025 B.n908 B.n55 585
R1026 B.n863 B.n54 585
R1027 B.n909 B.n54 585
R1028 B.n862 B.n861 585
R1029 B.n861 B.n53 585
R1030 B.n860 B.n49 585
R1031 B.n915 B.n49 585
R1032 B.n859 B.n48 585
R1033 B.n916 B.n48 585
R1034 B.n858 B.n47 585
R1035 B.n917 B.n47 585
R1036 B.n857 B.n856 585
R1037 B.n856 B.n43 585
R1038 B.n855 B.n42 585
R1039 B.n923 B.n42 585
R1040 B.n854 B.n41 585
R1041 B.n924 B.n41 585
R1042 B.n853 B.n40 585
R1043 B.n925 B.n40 585
R1044 B.n852 B.n851 585
R1045 B.n851 B.n36 585
R1046 B.n850 B.n35 585
R1047 B.n931 B.n35 585
R1048 B.n849 B.n34 585
R1049 B.n932 B.n34 585
R1050 B.n848 B.n33 585
R1051 B.n933 B.n33 585
R1052 B.n847 B.n846 585
R1053 B.n846 B.n29 585
R1054 B.n845 B.n28 585
R1055 B.n939 B.n28 585
R1056 B.n844 B.n27 585
R1057 B.n940 B.n27 585
R1058 B.n843 B.n26 585
R1059 B.n941 B.n26 585
R1060 B.n842 B.n841 585
R1061 B.n841 B.n22 585
R1062 B.n840 B.n21 585
R1063 B.n947 B.n21 585
R1064 B.n839 B.n20 585
R1065 B.n948 B.n20 585
R1066 B.n838 B.n19 585
R1067 B.n949 B.n19 585
R1068 B.n837 B.n836 585
R1069 B.n836 B.n15 585
R1070 B.n835 B.n14 585
R1071 B.n955 B.n14 585
R1072 B.n834 B.n13 585
R1073 B.n956 B.n13 585
R1074 B.n833 B.n12 585
R1075 B.n957 B.n12 585
R1076 B.n832 B.n831 585
R1077 B.n831 B.n8 585
R1078 B.n830 B.n7 585
R1079 B.n963 B.n7 585
R1080 B.n829 B.n6 585
R1081 B.n964 B.n6 585
R1082 B.n828 B.n5 585
R1083 B.n965 B.n5 585
R1084 B.n827 B.n826 585
R1085 B.n826 B.n4 585
R1086 B.n825 B.n350 585
R1087 B.n825 B.n824 585
R1088 B.n815 B.n351 585
R1089 B.n352 B.n351 585
R1090 B.n817 B.n816 585
R1091 B.n818 B.n817 585
R1092 B.n814 B.n356 585
R1093 B.n360 B.n356 585
R1094 B.n813 B.n812 585
R1095 B.n812 B.n811 585
R1096 B.n358 B.n357 585
R1097 B.n359 B.n358 585
R1098 B.n804 B.n803 585
R1099 B.n805 B.n804 585
R1100 B.n802 B.n365 585
R1101 B.n365 B.n364 585
R1102 B.n801 B.n800 585
R1103 B.n800 B.n799 585
R1104 B.n367 B.n366 585
R1105 B.n368 B.n367 585
R1106 B.n792 B.n791 585
R1107 B.n793 B.n792 585
R1108 B.n790 B.n373 585
R1109 B.n373 B.n372 585
R1110 B.n789 B.n788 585
R1111 B.n788 B.n787 585
R1112 B.n375 B.n374 585
R1113 B.n376 B.n375 585
R1114 B.n780 B.n779 585
R1115 B.n781 B.n780 585
R1116 B.n778 B.n381 585
R1117 B.n381 B.n380 585
R1118 B.n777 B.n776 585
R1119 B.n776 B.n775 585
R1120 B.n383 B.n382 585
R1121 B.n384 B.n383 585
R1122 B.n768 B.n767 585
R1123 B.n769 B.n768 585
R1124 B.n766 B.n388 585
R1125 B.n392 B.n388 585
R1126 B.n765 B.n764 585
R1127 B.n764 B.n763 585
R1128 B.n390 B.n389 585
R1129 B.n391 B.n390 585
R1130 B.n756 B.n755 585
R1131 B.n757 B.n756 585
R1132 B.n754 B.n397 585
R1133 B.n397 B.n396 585
R1134 B.n753 B.n752 585
R1135 B.n752 B.n751 585
R1136 B.n399 B.n398 585
R1137 B.n744 B.n399 585
R1138 B.n743 B.n742 585
R1139 B.n745 B.n743 585
R1140 B.n741 B.n404 585
R1141 B.n404 B.n403 585
R1142 B.n740 B.n739 585
R1143 B.n739 B.n738 585
R1144 B.n406 B.n405 585
R1145 B.n407 B.n406 585
R1146 B.n731 B.n730 585
R1147 B.n732 B.n731 585
R1148 B.n729 B.n412 585
R1149 B.n412 B.n411 585
R1150 B.n728 B.n727 585
R1151 B.n727 B.n726 585
R1152 B.n414 B.n413 585
R1153 B.n415 B.n414 585
R1154 B.n719 B.n718 585
R1155 B.n720 B.n719 585
R1156 B.n717 B.n420 585
R1157 B.n420 B.n419 585
R1158 B.n716 B.n715 585
R1159 B.n715 B.n714 585
R1160 B.n422 B.n421 585
R1161 B.n423 B.n422 585
R1162 B.n707 B.n706 585
R1163 B.n708 B.n707 585
R1164 B.n705 B.n428 585
R1165 B.n428 B.n427 585
R1166 B.n700 B.n699 585
R1167 B.n698 B.n484 585
R1168 B.n697 B.n483 585
R1169 B.n702 B.n483 585
R1170 B.n696 B.n695 585
R1171 B.n694 B.n693 585
R1172 B.n692 B.n691 585
R1173 B.n690 B.n689 585
R1174 B.n688 B.n687 585
R1175 B.n686 B.n685 585
R1176 B.n684 B.n683 585
R1177 B.n682 B.n681 585
R1178 B.n680 B.n679 585
R1179 B.n678 B.n677 585
R1180 B.n676 B.n675 585
R1181 B.n674 B.n673 585
R1182 B.n672 B.n671 585
R1183 B.n670 B.n669 585
R1184 B.n668 B.n667 585
R1185 B.n666 B.n665 585
R1186 B.n664 B.n663 585
R1187 B.n662 B.n661 585
R1188 B.n660 B.n659 585
R1189 B.n658 B.n657 585
R1190 B.n656 B.n655 585
R1191 B.n654 B.n653 585
R1192 B.n652 B.n651 585
R1193 B.n650 B.n649 585
R1194 B.n648 B.n647 585
R1195 B.n646 B.n645 585
R1196 B.n644 B.n643 585
R1197 B.n642 B.n641 585
R1198 B.n640 B.n639 585
R1199 B.n638 B.n637 585
R1200 B.n636 B.n635 585
R1201 B.n634 B.n633 585
R1202 B.n632 B.n631 585
R1203 B.n630 B.n629 585
R1204 B.n628 B.n627 585
R1205 B.n626 B.n625 585
R1206 B.n624 B.n623 585
R1207 B.n622 B.n621 585
R1208 B.n620 B.n619 585
R1209 B.n618 B.n617 585
R1210 B.n616 B.n615 585
R1211 B.n614 B.n613 585
R1212 B.n612 B.n611 585
R1213 B.n610 B.n609 585
R1214 B.n608 B.n607 585
R1215 B.n606 B.n605 585
R1216 B.n604 B.n603 585
R1217 B.n602 B.n601 585
R1218 B.n600 B.n599 585
R1219 B.n598 B.n597 585
R1220 B.n596 B.n595 585
R1221 B.n594 B.n593 585
R1222 B.n592 B.n591 585
R1223 B.n590 B.n589 585
R1224 B.n588 B.n587 585
R1225 B.n586 B.n585 585
R1226 B.n584 B.n583 585
R1227 B.n582 B.n581 585
R1228 B.n580 B.n579 585
R1229 B.n578 B.n577 585
R1230 B.n576 B.n575 585
R1231 B.n574 B.n573 585
R1232 B.n572 B.n571 585
R1233 B.n570 B.n569 585
R1234 B.n568 B.n567 585
R1235 B.n566 B.n565 585
R1236 B.n564 B.n563 585
R1237 B.n562 B.n561 585
R1238 B.n560 B.n559 585
R1239 B.n558 B.n557 585
R1240 B.n556 B.n555 585
R1241 B.n554 B.n553 585
R1242 B.n552 B.n551 585
R1243 B.n550 B.n549 585
R1244 B.n548 B.n547 585
R1245 B.n546 B.n545 585
R1246 B.n544 B.n543 585
R1247 B.n542 B.n541 585
R1248 B.n540 B.n539 585
R1249 B.n538 B.n537 585
R1250 B.n536 B.n535 585
R1251 B.n534 B.n533 585
R1252 B.n532 B.n531 585
R1253 B.n530 B.n529 585
R1254 B.n528 B.n527 585
R1255 B.n526 B.n525 585
R1256 B.n524 B.n523 585
R1257 B.n522 B.n521 585
R1258 B.n520 B.n519 585
R1259 B.n518 B.n517 585
R1260 B.n516 B.n515 585
R1261 B.n514 B.n513 585
R1262 B.n512 B.n511 585
R1263 B.n510 B.n509 585
R1264 B.n508 B.n507 585
R1265 B.n506 B.n505 585
R1266 B.n504 B.n503 585
R1267 B.n502 B.n501 585
R1268 B.n500 B.n499 585
R1269 B.n498 B.n497 585
R1270 B.n496 B.n495 585
R1271 B.n494 B.n493 585
R1272 B.n492 B.n491 585
R1273 B.n430 B.n429 585
R1274 B.n704 B.n703 585
R1275 B.n703 B.n702 585
R1276 B.n426 B.n425 585
R1277 B.n427 B.n426 585
R1278 B.n710 B.n709 585
R1279 B.n709 B.n708 585
R1280 B.n711 B.n424 585
R1281 B.n424 B.n423 585
R1282 B.n713 B.n712 585
R1283 B.n714 B.n713 585
R1284 B.n418 B.n417 585
R1285 B.n419 B.n418 585
R1286 B.n722 B.n721 585
R1287 B.n721 B.n720 585
R1288 B.n723 B.n416 585
R1289 B.n416 B.n415 585
R1290 B.n725 B.n724 585
R1291 B.n726 B.n725 585
R1292 B.n410 B.n409 585
R1293 B.n411 B.n410 585
R1294 B.n734 B.n733 585
R1295 B.n733 B.n732 585
R1296 B.n735 B.n408 585
R1297 B.n408 B.n407 585
R1298 B.n737 B.n736 585
R1299 B.n738 B.n737 585
R1300 B.n402 B.n401 585
R1301 B.n403 B.n402 585
R1302 B.n747 B.n746 585
R1303 B.n746 B.n745 585
R1304 B.n748 B.n400 585
R1305 B.n744 B.n400 585
R1306 B.n750 B.n749 585
R1307 B.n751 B.n750 585
R1308 B.n395 B.n394 585
R1309 B.n396 B.n395 585
R1310 B.n759 B.n758 585
R1311 B.n758 B.n757 585
R1312 B.n760 B.n393 585
R1313 B.n393 B.n391 585
R1314 B.n762 B.n761 585
R1315 B.n763 B.n762 585
R1316 B.n387 B.n386 585
R1317 B.n392 B.n387 585
R1318 B.n771 B.n770 585
R1319 B.n770 B.n769 585
R1320 B.n772 B.n385 585
R1321 B.n385 B.n384 585
R1322 B.n774 B.n773 585
R1323 B.n775 B.n774 585
R1324 B.n379 B.n378 585
R1325 B.n380 B.n379 585
R1326 B.n783 B.n782 585
R1327 B.n782 B.n781 585
R1328 B.n784 B.n377 585
R1329 B.n377 B.n376 585
R1330 B.n786 B.n785 585
R1331 B.n787 B.n786 585
R1332 B.n371 B.n370 585
R1333 B.n372 B.n371 585
R1334 B.n795 B.n794 585
R1335 B.n794 B.n793 585
R1336 B.n796 B.n369 585
R1337 B.n369 B.n368 585
R1338 B.n798 B.n797 585
R1339 B.n799 B.n798 585
R1340 B.n363 B.n362 585
R1341 B.n364 B.n363 585
R1342 B.n807 B.n806 585
R1343 B.n806 B.n805 585
R1344 B.n808 B.n361 585
R1345 B.n361 B.n359 585
R1346 B.n810 B.n809 585
R1347 B.n811 B.n810 585
R1348 B.n355 B.n354 585
R1349 B.n360 B.n355 585
R1350 B.n820 B.n819 585
R1351 B.n819 B.n818 585
R1352 B.n821 B.n353 585
R1353 B.n353 B.n352 585
R1354 B.n823 B.n822 585
R1355 B.n824 B.n823 585
R1356 B.n2 B.n0 585
R1357 B.n4 B.n2 585
R1358 B.n3 B.n1 585
R1359 B.n964 B.n3 585
R1360 B.n962 B.n961 585
R1361 B.n963 B.n962 585
R1362 B.n960 B.n9 585
R1363 B.n9 B.n8 585
R1364 B.n959 B.n958 585
R1365 B.n958 B.n957 585
R1366 B.n11 B.n10 585
R1367 B.n956 B.n11 585
R1368 B.n954 B.n953 585
R1369 B.n955 B.n954 585
R1370 B.n952 B.n16 585
R1371 B.n16 B.n15 585
R1372 B.n951 B.n950 585
R1373 B.n950 B.n949 585
R1374 B.n18 B.n17 585
R1375 B.n948 B.n18 585
R1376 B.n946 B.n945 585
R1377 B.n947 B.n946 585
R1378 B.n944 B.n23 585
R1379 B.n23 B.n22 585
R1380 B.n943 B.n942 585
R1381 B.n942 B.n941 585
R1382 B.n25 B.n24 585
R1383 B.n940 B.n25 585
R1384 B.n938 B.n937 585
R1385 B.n939 B.n938 585
R1386 B.n936 B.n30 585
R1387 B.n30 B.n29 585
R1388 B.n935 B.n934 585
R1389 B.n934 B.n933 585
R1390 B.n32 B.n31 585
R1391 B.n932 B.n32 585
R1392 B.n930 B.n929 585
R1393 B.n931 B.n930 585
R1394 B.n928 B.n37 585
R1395 B.n37 B.n36 585
R1396 B.n927 B.n926 585
R1397 B.n926 B.n925 585
R1398 B.n39 B.n38 585
R1399 B.n924 B.n39 585
R1400 B.n922 B.n921 585
R1401 B.n923 B.n922 585
R1402 B.n920 B.n44 585
R1403 B.n44 B.n43 585
R1404 B.n919 B.n918 585
R1405 B.n918 B.n917 585
R1406 B.n46 B.n45 585
R1407 B.n916 B.n46 585
R1408 B.n914 B.n913 585
R1409 B.n915 B.n914 585
R1410 B.n912 B.n50 585
R1411 B.n53 B.n50 585
R1412 B.n911 B.n910 585
R1413 B.n910 B.n909 585
R1414 B.n52 B.n51 585
R1415 B.n908 B.n52 585
R1416 B.n906 B.n905 585
R1417 B.n907 B.n906 585
R1418 B.n904 B.n58 585
R1419 B.n58 B.n57 585
R1420 B.n903 B.n902 585
R1421 B.n902 B.n901 585
R1422 B.n60 B.n59 585
R1423 B.n900 B.n60 585
R1424 B.n898 B.n897 585
R1425 B.n899 B.n898 585
R1426 B.n896 B.n65 585
R1427 B.n65 B.n64 585
R1428 B.n895 B.n894 585
R1429 B.n894 B.n893 585
R1430 B.n67 B.n66 585
R1431 B.n892 B.n67 585
R1432 B.n890 B.n889 585
R1433 B.n891 B.n890 585
R1434 B.n888 B.n72 585
R1435 B.n72 B.n71 585
R1436 B.n887 B.n886 585
R1437 B.n886 B.n885 585
R1438 B.n74 B.n73 585
R1439 B.n884 B.n74 585
R1440 B.n967 B.n966 585
R1441 B.n966 B.n965 585
R1442 B.n700 B.n426 540.549
R1443 B.n135 B.n74 540.549
R1444 B.n703 B.n428 540.549
R1445 B.n881 B.n76 540.549
R1446 B.n488 B.t10 434.536
R1447 B.n485 B.t21 434.536
R1448 B.n133 B.t14 434.536
R1449 B.n131 B.t18 434.536
R1450 B.n488 B.t13 363.378
R1451 B.n485 B.t23 363.378
R1452 B.n133 B.t16 363.378
R1453 B.n131 B.t19 363.378
R1454 B.n489 B.t12 327.113
R1455 B.n132 B.t20 327.113
R1456 B.n486 B.t22 327.113
R1457 B.n134 B.t17 327.113
R1458 B.n883 B.n882 256.663
R1459 B.n883 B.n129 256.663
R1460 B.n883 B.n128 256.663
R1461 B.n883 B.n127 256.663
R1462 B.n883 B.n126 256.663
R1463 B.n883 B.n125 256.663
R1464 B.n883 B.n124 256.663
R1465 B.n883 B.n123 256.663
R1466 B.n883 B.n122 256.663
R1467 B.n883 B.n121 256.663
R1468 B.n883 B.n120 256.663
R1469 B.n883 B.n119 256.663
R1470 B.n883 B.n118 256.663
R1471 B.n883 B.n117 256.663
R1472 B.n883 B.n116 256.663
R1473 B.n883 B.n115 256.663
R1474 B.n883 B.n114 256.663
R1475 B.n883 B.n113 256.663
R1476 B.n883 B.n112 256.663
R1477 B.n883 B.n111 256.663
R1478 B.n883 B.n110 256.663
R1479 B.n883 B.n109 256.663
R1480 B.n883 B.n108 256.663
R1481 B.n883 B.n107 256.663
R1482 B.n883 B.n106 256.663
R1483 B.n883 B.n105 256.663
R1484 B.n883 B.n104 256.663
R1485 B.n883 B.n103 256.663
R1486 B.n883 B.n102 256.663
R1487 B.n883 B.n101 256.663
R1488 B.n883 B.n100 256.663
R1489 B.n883 B.n99 256.663
R1490 B.n883 B.n98 256.663
R1491 B.n883 B.n97 256.663
R1492 B.n883 B.n96 256.663
R1493 B.n883 B.n95 256.663
R1494 B.n883 B.n94 256.663
R1495 B.n883 B.n93 256.663
R1496 B.n883 B.n92 256.663
R1497 B.n883 B.n91 256.663
R1498 B.n883 B.n90 256.663
R1499 B.n883 B.n89 256.663
R1500 B.n883 B.n88 256.663
R1501 B.n883 B.n87 256.663
R1502 B.n883 B.n86 256.663
R1503 B.n883 B.n85 256.663
R1504 B.n883 B.n84 256.663
R1505 B.n883 B.n83 256.663
R1506 B.n883 B.n82 256.663
R1507 B.n883 B.n81 256.663
R1508 B.n883 B.n80 256.663
R1509 B.n883 B.n79 256.663
R1510 B.n883 B.n78 256.663
R1511 B.n883 B.n77 256.663
R1512 B.n702 B.n701 256.663
R1513 B.n702 B.n431 256.663
R1514 B.n702 B.n432 256.663
R1515 B.n702 B.n433 256.663
R1516 B.n702 B.n434 256.663
R1517 B.n702 B.n435 256.663
R1518 B.n702 B.n436 256.663
R1519 B.n702 B.n437 256.663
R1520 B.n702 B.n438 256.663
R1521 B.n702 B.n439 256.663
R1522 B.n702 B.n440 256.663
R1523 B.n702 B.n441 256.663
R1524 B.n702 B.n442 256.663
R1525 B.n702 B.n443 256.663
R1526 B.n702 B.n444 256.663
R1527 B.n702 B.n445 256.663
R1528 B.n702 B.n446 256.663
R1529 B.n702 B.n447 256.663
R1530 B.n702 B.n448 256.663
R1531 B.n702 B.n449 256.663
R1532 B.n702 B.n450 256.663
R1533 B.n702 B.n451 256.663
R1534 B.n702 B.n452 256.663
R1535 B.n702 B.n453 256.663
R1536 B.n702 B.n454 256.663
R1537 B.n702 B.n455 256.663
R1538 B.n702 B.n456 256.663
R1539 B.n702 B.n457 256.663
R1540 B.n702 B.n458 256.663
R1541 B.n702 B.n459 256.663
R1542 B.n702 B.n460 256.663
R1543 B.n702 B.n461 256.663
R1544 B.n702 B.n462 256.663
R1545 B.n702 B.n463 256.663
R1546 B.n702 B.n464 256.663
R1547 B.n702 B.n465 256.663
R1548 B.n702 B.n466 256.663
R1549 B.n702 B.n467 256.663
R1550 B.n702 B.n468 256.663
R1551 B.n702 B.n469 256.663
R1552 B.n702 B.n470 256.663
R1553 B.n702 B.n471 256.663
R1554 B.n702 B.n472 256.663
R1555 B.n702 B.n473 256.663
R1556 B.n702 B.n474 256.663
R1557 B.n702 B.n475 256.663
R1558 B.n702 B.n476 256.663
R1559 B.n702 B.n477 256.663
R1560 B.n702 B.n478 256.663
R1561 B.n702 B.n479 256.663
R1562 B.n702 B.n480 256.663
R1563 B.n702 B.n481 256.663
R1564 B.n702 B.n482 256.663
R1565 B.n709 B.n426 163.367
R1566 B.n709 B.n424 163.367
R1567 B.n713 B.n424 163.367
R1568 B.n713 B.n418 163.367
R1569 B.n721 B.n418 163.367
R1570 B.n721 B.n416 163.367
R1571 B.n725 B.n416 163.367
R1572 B.n725 B.n410 163.367
R1573 B.n733 B.n410 163.367
R1574 B.n733 B.n408 163.367
R1575 B.n737 B.n408 163.367
R1576 B.n737 B.n402 163.367
R1577 B.n746 B.n402 163.367
R1578 B.n746 B.n400 163.367
R1579 B.n750 B.n400 163.367
R1580 B.n750 B.n395 163.367
R1581 B.n758 B.n395 163.367
R1582 B.n758 B.n393 163.367
R1583 B.n762 B.n393 163.367
R1584 B.n762 B.n387 163.367
R1585 B.n770 B.n387 163.367
R1586 B.n770 B.n385 163.367
R1587 B.n774 B.n385 163.367
R1588 B.n774 B.n379 163.367
R1589 B.n782 B.n379 163.367
R1590 B.n782 B.n377 163.367
R1591 B.n786 B.n377 163.367
R1592 B.n786 B.n371 163.367
R1593 B.n794 B.n371 163.367
R1594 B.n794 B.n369 163.367
R1595 B.n798 B.n369 163.367
R1596 B.n798 B.n363 163.367
R1597 B.n806 B.n363 163.367
R1598 B.n806 B.n361 163.367
R1599 B.n810 B.n361 163.367
R1600 B.n810 B.n355 163.367
R1601 B.n819 B.n355 163.367
R1602 B.n819 B.n353 163.367
R1603 B.n823 B.n353 163.367
R1604 B.n823 B.n2 163.367
R1605 B.n966 B.n2 163.367
R1606 B.n966 B.n3 163.367
R1607 B.n962 B.n3 163.367
R1608 B.n962 B.n9 163.367
R1609 B.n958 B.n9 163.367
R1610 B.n958 B.n11 163.367
R1611 B.n954 B.n11 163.367
R1612 B.n954 B.n16 163.367
R1613 B.n950 B.n16 163.367
R1614 B.n950 B.n18 163.367
R1615 B.n946 B.n18 163.367
R1616 B.n946 B.n23 163.367
R1617 B.n942 B.n23 163.367
R1618 B.n942 B.n25 163.367
R1619 B.n938 B.n25 163.367
R1620 B.n938 B.n30 163.367
R1621 B.n934 B.n30 163.367
R1622 B.n934 B.n32 163.367
R1623 B.n930 B.n32 163.367
R1624 B.n930 B.n37 163.367
R1625 B.n926 B.n37 163.367
R1626 B.n926 B.n39 163.367
R1627 B.n922 B.n39 163.367
R1628 B.n922 B.n44 163.367
R1629 B.n918 B.n44 163.367
R1630 B.n918 B.n46 163.367
R1631 B.n914 B.n46 163.367
R1632 B.n914 B.n50 163.367
R1633 B.n910 B.n50 163.367
R1634 B.n910 B.n52 163.367
R1635 B.n906 B.n52 163.367
R1636 B.n906 B.n58 163.367
R1637 B.n902 B.n58 163.367
R1638 B.n902 B.n60 163.367
R1639 B.n898 B.n60 163.367
R1640 B.n898 B.n65 163.367
R1641 B.n894 B.n65 163.367
R1642 B.n894 B.n67 163.367
R1643 B.n890 B.n67 163.367
R1644 B.n890 B.n72 163.367
R1645 B.n886 B.n72 163.367
R1646 B.n886 B.n74 163.367
R1647 B.n484 B.n483 163.367
R1648 B.n695 B.n483 163.367
R1649 B.n693 B.n692 163.367
R1650 B.n689 B.n688 163.367
R1651 B.n685 B.n684 163.367
R1652 B.n681 B.n680 163.367
R1653 B.n677 B.n676 163.367
R1654 B.n673 B.n672 163.367
R1655 B.n669 B.n668 163.367
R1656 B.n665 B.n664 163.367
R1657 B.n661 B.n660 163.367
R1658 B.n657 B.n656 163.367
R1659 B.n653 B.n652 163.367
R1660 B.n649 B.n648 163.367
R1661 B.n645 B.n644 163.367
R1662 B.n641 B.n640 163.367
R1663 B.n637 B.n636 163.367
R1664 B.n633 B.n632 163.367
R1665 B.n629 B.n628 163.367
R1666 B.n625 B.n624 163.367
R1667 B.n621 B.n620 163.367
R1668 B.n617 B.n616 163.367
R1669 B.n613 B.n612 163.367
R1670 B.n609 B.n608 163.367
R1671 B.n605 B.n604 163.367
R1672 B.n601 B.n600 163.367
R1673 B.n597 B.n596 163.367
R1674 B.n593 B.n592 163.367
R1675 B.n589 B.n588 163.367
R1676 B.n585 B.n584 163.367
R1677 B.n581 B.n580 163.367
R1678 B.n577 B.n576 163.367
R1679 B.n573 B.n572 163.367
R1680 B.n569 B.n568 163.367
R1681 B.n565 B.n564 163.367
R1682 B.n561 B.n560 163.367
R1683 B.n557 B.n556 163.367
R1684 B.n553 B.n552 163.367
R1685 B.n549 B.n548 163.367
R1686 B.n545 B.n544 163.367
R1687 B.n541 B.n540 163.367
R1688 B.n537 B.n536 163.367
R1689 B.n533 B.n532 163.367
R1690 B.n529 B.n528 163.367
R1691 B.n525 B.n524 163.367
R1692 B.n521 B.n520 163.367
R1693 B.n517 B.n516 163.367
R1694 B.n513 B.n512 163.367
R1695 B.n509 B.n508 163.367
R1696 B.n505 B.n504 163.367
R1697 B.n501 B.n500 163.367
R1698 B.n497 B.n496 163.367
R1699 B.n493 B.n492 163.367
R1700 B.n703 B.n430 163.367
R1701 B.n707 B.n428 163.367
R1702 B.n707 B.n422 163.367
R1703 B.n715 B.n422 163.367
R1704 B.n715 B.n420 163.367
R1705 B.n719 B.n420 163.367
R1706 B.n719 B.n414 163.367
R1707 B.n727 B.n414 163.367
R1708 B.n727 B.n412 163.367
R1709 B.n731 B.n412 163.367
R1710 B.n731 B.n406 163.367
R1711 B.n739 B.n406 163.367
R1712 B.n739 B.n404 163.367
R1713 B.n743 B.n404 163.367
R1714 B.n743 B.n399 163.367
R1715 B.n752 B.n399 163.367
R1716 B.n752 B.n397 163.367
R1717 B.n756 B.n397 163.367
R1718 B.n756 B.n390 163.367
R1719 B.n764 B.n390 163.367
R1720 B.n764 B.n388 163.367
R1721 B.n768 B.n388 163.367
R1722 B.n768 B.n383 163.367
R1723 B.n776 B.n383 163.367
R1724 B.n776 B.n381 163.367
R1725 B.n780 B.n381 163.367
R1726 B.n780 B.n375 163.367
R1727 B.n788 B.n375 163.367
R1728 B.n788 B.n373 163.367
R1729 B.n792 B.n373 163.367
R1730 B.n792 B.n367 163.367
R1731 B.n800 B.n367 163.367
R1732 B.n800 B.n365 163.367
R1733 B.n804 B.n365 163.367
R1734 B.n804 B.n358 163.367
R1735 B.n812 B.n358 163.367
R1736 B.n812 B.n356 163.367
R1737 B.n817 B.n356 163.367
R1738 B.n817 B.n351 163.367
R1739 B.n825 B.n351 163.367
R1740 B.n826 B.n825 163.367
R1741 B.n826 B.n5 163.367
R1742 B.n6 B.n5 163.367
R1743 B.n7 B.n6 163.367
R1744 B.n831 B.n7 163.367
R1745 B.n831 B.n12 163.367
R1746 B.n13 B.n12 163.367
R1747 B.n14 B.n13 163.367
R1748 B.n836 B.n14 163.367
R1749 B.n836 B.n19 163.367
R1750 B.n20 B.n19 163.367
R1751 B.n21 B.n20 163.367
R1752 B.n841 B.n21 163.367
R1753 B.n841 B.n26 163.367
R1754 B.n27 B.n26 163.367
R1755 B.n28 B.n27 163.367
R1756 B.n846 B.n28 163.367
R1757 B.n846 B.n33 163.367
R1758 B.n34 B.n33 163.367
R1759 B.n35 B.n34 163.367
R1760 B.n851 B.n35 163.367
R1761 B.n851 B.n40 163.367
R1762 B.n41 B.n40 163.367
R1763 B.n42 B.n41 163.367
R1764 B.n856 B.n42 163.367
R1765 B.n856 B.n47 163.367
R1766 B.n48 B.n47 163.367
R1767 B.n49 B.n48 163.367
R1768 B.n861 B.n49 163.367
R1769 B.n861 B.n54 163.367
R1770 B.n55 B.n54 163.367
R1771 B.n56 B.n55 163.367
R1772 B.n866 B.n56 163.367
R1773 B.n866 B.n61 163.367
R1774 B.n62 B.n61 163.367
R1775 B.n63 B.n62 163.367
R1776 B.n871 B.n63 163.367
R1777 B.n871 B.n68 163.367
R1778 B.n69 B.n68 163.367
R1779 B.n70 B.n69 163.367
R1780 B.n876 B.n70 163.367
R1781 B.n876 B.n75 163.367
R1782 B.n76 B.n75 163.367
R1783 B.n139 B.n138 163.367
R1784 B.n143 B.n142 163.367
R1785 B.n147 B.n146 163.367
R1786 B.n151 B.n150 163.367
R1787 B.n155 B.n154 163.367
R1788 B.n159 B.n158 163.367
R1789 B.n163 B.n162 163.367
R1790 B.n167 B.n166 163.367
R1791 B.n171 B.n170 163.367
R1792 B.n175 B.n174 163.367
R1793 B.n179 B.n178 163.367
R1794 B.n183 B.n182 163.367
R1795 B.n187 B.n186 163.367
R1796 B.n191 B.n190 163.367
R1797 B.n195 B.n194 163.367
R1798 B.n199 B.n198 163.367
R1799 B.n203 B.n202 163.367
R1800 B.n207 B.n206 163.367
R1801 B.n211 B.n210 163.367
R1802 B.n215 B.n214 163.367
R1803 B.n219 B.n218 163.367
R1804 B.n223 B.n222 163.367
R1805 B.n227 B.n226 163.367
R1806 B.n231 B.n230 163.367
R1807 B.n236 B.n235 163.367
R1808 B.n240 B.n239 163.367
R1809 B.n244 B.n243 163.367
R1810 B.n248 B.n247 163.367
R1811 B.n252 B.n251 163.367
R1812 B.n257 B.n256 163.367
R1813 B.n261 B.n260 163.367
R1814 B.n265 B.n264 163.367
R1815 B.n269 B.n268 163.367
R1816 B.n273 B.n272 163.367
R1817 B.n277 B.n276 163.367
R1818 B.n281 B.n280 163.367
R1819 B.n285 B.n284 163.367
R1820 B.n289 B.n288 163.367
R1821 B.n293 B.n292 163.367
R1822 B.n297 B.n296 163.367
R1823 B.n301 B.n300 163.367
R1824 B.n305 B.n304 163.367
R1825 B.n309 B.n308 163.367
R1826 B.n313 B.n312 163.367
R1827 B.n317 B.n316 163.367
R1828 B.n321 B.n320 163.367
R1829 B.n325 B.n324 163.367
R1830 B.n329 B.n328 163.367
R1831 B.n333 B.n332 163.367
R1832 B.n337 B.n336 163.367
R1833 B.n341 B.n340 163.367
R1834 B.n345 B.n344 163.367
R1835 B.n347 B.n130 163.367
R1836 B.n702 B.n427 72.3944
R1837 B.n884 B.n883 72.3944
R1838 B.n701 B.n700 71.676
R1839 B.n695 B.n431 71.676
R1840 B.n692 B.n432 71.676
R1841 B.n688 B.n433 71.676
R1842 B.n684 B.n434 71.676
R1843 B.n680 B.n435 71.676
R1844 B.n676 B.n436 71.676
R1845 B.n672 B.n437 71.676
R1846 B.n668 B.n438 71.676
R1847 B.n664 B.n439 71.676
R1848 B.n660 B.n440 71.676
R1849 B.n656 B.n441 71.676
R1850 B.n652 B.n442 71.676
R1851 B.n648 B.n443 71.676
R1852 B.n644 B.n444 71.676
R1853 B.n640 B.n445 71.676
R1854 B.n636 B.n446 71.676
R1855 B.n632 B.n447 71.676
R1856 B.n628 B.n448 71.676
R1857 B.n624 B.n449 71.676
R1858 B.n620 B.n450 71.676
R1859 B.n616 B.n451 71.676
R1860 B.n612 B.n452 71.676
R1861 B.n608 B.n453 71.676
R1862 B.n604 B.n454 71.676
R1863 B.n600 B.n455 71.676
R1864 B.n596 B.n456 71.676
R1865 B.n592 B.n457 71.676
R1866 B.n588 B.n458 71.676
R1867 B.n584 B.n459 71.676
R1868 B.n580 B.n460 71.676
R1869 B.n576 B.n461 71.676
R1870 B.n572 B.n462 71.676
R1871 B.n568 B.n463 71.676
R1872 B.n564 B.n464 71.676
R1873 B.n560 B.n465 71.676
R1874 B.n556 B.n466 71.676
R1875 B.n552 B.n467 71.676
R1876 B.n548 B.n468 71.676
R1877 B.n544 B.n469 71.676
R1878 B.n540 B.n470 71.676
R1879 B.n536 B.n471 71.676
R1880 B.n532 B.n472 71.676
R1881 B.n528 B.n473 71.676
R1882 B.n524 B.n474 71.676
R1883 B.n520 B.n475 71.676
R1884 B.n516 B.n476 71.676
R1885 B.n512 B.n477 71.676
R1886 B.n508 B.n478 71.676
R1887 B.n504 B.n479 71.676
R1888 B.n500 B.n480 71.676
R1889 B.n496 B.n481 71.676
R1890 B.n492 B.n482 71.676
R1891 B.n135 B.n77 71.676
R1892 B.n139 B.n78 71.676
R1893 B.n143 B.n79 71.676
R1894 B.n147 B.n80 71.676
R1895 B.n151 B.n81 71.676
R1896 B.n155 B.n82 71.676
R1897 B.n159 B.n83 71.676
R1898 B.n163 B.n84 71.676
R1899 B.n167 B.n85 71.676
R1900 B.n171 B.n86 71.676
R1901 B.n175 B.n87 71.676
R1902 B.n179 B.n88 71.676
R1903 B.n183 B.n89 71.676
R1904 B.n187 B.n90 71.676
R1905 B.n191 B.n91 71.676
R1906 B.n195 B.n92 71.676
R1907 B.n199 B.n93 71.676
R1908 B.n203 B.n94 71.676
R1909 B.n207 B.n95 71.676
R1910 B.n211 B.n96 71.676
R1911 B.n215 B.n97 71.676
R1912 B.n219 B.n98 71.676
R1913 B.n223 B.n99 71.676
R1914 B.n227 B.n100 71.676
R1915 B.n231 B.n101 71.676
R1916 B.n236 B.n102 71.676
R1917 B.n240 B.n103 71.676
R1918 B.n244 B.n104 71.676
R1919 B.n248 B.n105 71.676
R1920 B.n252 B.n106 71.676
R1921 B.n257 B.n107 71.676
R1922 B.n261 B.n108 71.676
R1923 B.n265 B.n109 71.676
R1924 B.n269 B.n110 71.676
R1925 B.n273 B.n111 71.676
R1926 B.n277 B.n112 71.676
R1927 B.n281 B.n113 71.676
R1928 B.n285 B.n114 71.676
R1929 B.n289 B.n115 71.676
R1930 B.n293 B.n116 71.676
R1931 B.n297 B.n117 71.676
R1932 B.n301 B.n118 71.676
R1933 B.n305 B.n119 71.676
R1934 B.n309 B.n120 71.676
R1935 B.n313 B.n121 71.676
R1936 B.n317 B.n122 71.676
R1937 B.n321 B.n123 71.676
R1938 B.n325 B.n124 71.676
R1939 B.n329 B.n125 71.676
R1940 B.n333 B.n126 71.676
R1941 B.n337 B.n127 71.676
R1942 B.n341 B.n128 71.676
R1943 B.n345 B.n129 71.676
R1944 B.n882 B.n130 71.676
R1945 B.n882 B.n881 71.676
R1946 B.n347 B.n129 71.676
R1947 B.n344 B.n128 71.676
R1948 B.n340 B.n127 71.676
R1949 B.n336 B.n126 71.676
R1950 B.n332 B.n125 71.676
R1951 B.n328 B.n124 71.676
R1952 B.n324 B.n123 71.676
R1953 B.n320 B.n122 71.676
R1954 B.n316 B.n121 71.676
R1955 B.n312 B.n120 71.676
R1956 B.n308 B.n119 71.676
R1957 B.n304 B.n118 71.676
R1958 B.n300 B.n117 71.676
R1959 B.n296 B.n116 71.676
R1960 B.n292 B.n115 71.676
R1961 B.n288 B.n114 71.676
R1962 B.n284 B.n113 71.676
R1963 B.n280 B.n112 71.676
R1964 B.n276 B.n111 71.676
R1965 B.n272 B.n110 71.676
R1966 B.n268 B.n109 71.676
R1967 B.n264 B.n108 71.676
R1968 B.n260 B.n107 71.676
R1969 B.n256 B.n106 71.676
R1970 B.n251 B.n105 71.676
R1971 B.n247 B.n104 71.676
R1972 B.n243 B.n103 71.676
R1973 B.n239 B.n102 71.676
R1974 B.n235 B.n101 71.676
R1975 B.n230 B.n100 71.676
R1976 B.n226 B.n99 71.676
R1977 B.n222 B.n98 71.676
R1978 B.n218 B.n97 71.676
R1979 B.n214 B.n96 71.676
R1980 B.n210 B.n95 71.676
R1981 B.n206 B.n94 71.676
R1982 B.n202 B.n93 71.676
R1983 B.n198 B.n92 71.676
R1984 B.n194 B.n91 71.676
R1985 B.n190 B.n90 71.676
R1986 B.n186 B.n89 71.676
R1987 B.n182 B.n88 71.676
R1988 B.n178 B.n87 71.676
R1989 B.n174 B.n86 71.676
R1990 B.n170 B.n85 71.676
R1991 B.n166 B.n84 71.676
R1992 B.n162 B.n83 71.676
R1993 B.n158 B.n82 71.676
R1994 B.n154 B.n81 71.676
R1995 B.n150 B.n80 71.676
R1996 B.n146 B.n79 71.676
R1997 B.n142 B.n78 71.676
R1998 B.n138 B.n77 71.676
R1999 B.n701 B.n484 71.676
R2000 B.n693 B.n431 71.676
R2001 B.n689 B.n432 71.676
R2002 B.n685 B.n433 71.676
R2003 B.n681 B.n434 71.676
R2004 B.n677 B.n435 71.676
R2005 B.n673 B.n436 71.676
R2006 B.n669 B.n437 71.676
R2007 B.n665 B.n438 71.676
R2008 B.n661 B.n439 71.676
R2009 B.n657 B.n440 71.676
R2010 B.n653 B.n441 71.676
R2011 B.n649 B.n442 71.676
R2012 B.n645 B.n443 71.676
R2013 B.n641 B.n444 71.676
R2014 B.n637 B.n445 71.676
R2015 B.n633 B.n446 71.676
R2016 B.n629 B.n447 71.676
R2017 B.n625 B.n448 71.676
R2018 B.n621 B.n449 71.676
R2019 B.n617 B.n450 71.676
R2020 B.n613 B.n451 71.676
R2021 B.n609 B.n452 71.676
R2022 B.n605 B.n453 71.676
R2023 B.n601 B.n454 71.676
R2024 B.n597 B.n455 71.676
R2025 B.n593 B.n456 71.676
R2026 B.n589 B.n457 71.676
R2027 B.n585 B.n458 71.676
R2028 B.n581 B.n459 71.676
R2029 B.n577 B.n460 71.676
R2030 B.n573 B.n461 71.676
R2031 B.n569 B.n462 71.676
R2032 B.n565 B.n463 71.676
R2033 B.n561 B.n464 71.676
R2034 B.n557 B.n465 71.676
R2035 B.n553 B.n466 71.676
R2036 B.n549 B.n467 71.676
R2037 B.n545 B.n468 71.676
R2038 B.n541 B.n469 71.676
R2039 B.n537 B.n470 71.676
R2040 B.n533 B.n471 71.676
R2041 B.n529 B.n472 71.676
R2042 B.n525 B.n473 71.676
R2043 B.n521 B.n474 71.676
R2044 B.n517 B.n475 71.676
R2045 B.n513 B.n476 71.676
R2046 B.n509 B.n477 71.676
R2047 B.n505 B.n478 71.676
R2048 B.n501 B.n479 71.676
R2049 B.n497 B.n480 71.676
R2050 B.n493 B.n481 71.676
R2051 B.n482 B.n430 71.676
R2052 B.n490 B.n489 59.5399
R2053 B.n487 B.n486 59.5399
R2054 B.n233 B.n134 59.5399
R2055 B.n254 B.n132 59.5399
R2056 B.n708 B.n427 37.579
R2057 B.n708 B.n423 37.579
R2058 B.n714 B.n423 37.579
R2059 B.n714 B.n419 37.579
R2060 B.n720 B.n419 37.579
R2061 B.n726 B.n415 37.579
R2062 B.n726 B.n411 37.579
R2063 B.n732 B.n411 37.579
R2064 B.n732 B.n407 37.579
R2065 B.n738 B.n407 37.579
R2066 B.n738 B.n403 37.579
R2067 B.n745 B.n403 37.579
R2068 B.n745 B.n744 37.579
R2069 B.n751 B.n396 37.579
R2070 B.n757 B.n396 37.579
R2071 B.n757 B.n391 37.579
R2072 B.n763 B.n391 37.579
R2073 B.n763 B.n392 37.579
R2074 B.n769 B.n384 37.579
R2075 B.n775 B.n384 37.579
R2076 B.n775 B.n380 37.579
R2077 B.n781 B.n380 37.579
R2078 B.n787 B.n376 37.579
R2079 B.n787 B.n372 37.579
R2080 B.n793 B.n372 37.579
R2081 B.n793 B.n368 37.579
R2082 B.n799 B.n368 37.579
R2083 B.n805 B.n364 37.579
R2084 B.n805 B.n359 37.579
R2085 B.n811 B.n359 37.579
R2086 B.n811 B.n360 37.579
R2087 B.n818 B.n352 37.579
R2088 B.n824 B.n352 37.579
R2089 B.n824 B.n4 37.579
R2090 B.n965 B.n4 37.579
R2091 B.n965 B.n964 37.579
R2092 B.n964 B.n963 37.579
R2093 B.n963 B.n8 37.579
R2094 B.n957 B.n8 37.579
R2095 B.n956 B.n955 37.579
R2096 B.n955 B.n15 37.579
R2097 B.n949 B.n15 37.579
R2098 B.n949 B.n948 37.579
R2099 B.n947 B.n22 37.579
R2100 B.n941 B.n22 37.579
R2101 B.n941 B.n940 37.579
R2102 B.n940 B.n939 37.579
R2103 B.n939 B.n29 37.579
R2104 B.n933 B.n932 37.579
R2105 B.n932 B.n931 37.579
R2106 B.n931 B.n36 37.579
R2107 B.n925 B.n36 37.579
R2108 B.n924 B.n923 37.579
R2109 B.n923 B.n43 37.579
R2110 B.n917 B.n43 37.579
R2111 B.n917 B.n916 37.579
R2112 B.n916 B.n915 37.579
R2113 B.n909 B.n53 37.579
R2114 B.n909 B.n908 37.579
R2115 B.n908 B.n907 37.579
R2116 B.n907 B.n57 37.579
R2117 B.n901 B.n57 37.579
R2118 B.n901 B.n900 37.579
R2119 B.n900 B.n899 37.579
R2120 B.n899 B.n64 37.579
R2121 B.n893 B.n892 37.579
R2122 B.n892 B.n891 37.579
R2123 B.n891 B.n71 37.579
R2124 B.n885 B.n71 37.579
R2125 B.n885 B.n884 37.579
R2126 B.n489 B.n488 36.2672
R2127 B.n486 B.n485 36.2672
R2128 B.n134 B.n133 36.2672
R2129 B.n132 B.n131 36.2672
R2130 B.n720 B.t11 35.3685
R2131 B.n893 B.t15 35.3685
R2132 B.n136 B.n73 35.1225
R2133 B.n705 B.n704 35.1225
R2134 B.n699 B.n425 35.1225
R2135 B.n880 B.n879 35.1224
R2136 B.n769 B.t2 32.0527
R2137 B.t1 B.n364 32.0527
R2138 B.n948 B.t4 32.0527
R2139 B.n925 B.t3 32.0527
R2140 B.n744 B.t9 24.316
R2141 B.n781 B.t5 24.316
R2142 B.n360 B.t6 24.316
R2143 B.t7 B.n956 24.316
R2144 B.n933 B.t8 24.316
R2145 B.n53 B.t0 24.316
R2146 B B.n967 18.0485
R2147 B.n751 B.t9 13.2635
R2148 B.t5 B.n376 13.2635
R2149 B.n818 B.t6 13.2635
R2150 B.n957 B.t7 13.2635
R2151 B.t8 B.n29 13.2635
R2152 B.n915 B.t0 13.2635
R2153 B.n137 B.n136 10.6151
R2154 B.n140 B.n137 10.6151
R2155 B.n141 B.n140 10.6151
R2156 B.n144 B.n141 10.6151
R2157 B.n145 B.n144 10.6151
R2158 B.n148 B.n145 10.6151
R2159 B.n149 B.n148 10.6151
R2160 B.n152 B.n149 10.6151
R2161 B.n153 B.n152 10.6151
R2162 B.n156 B.n153 10.6151
R2163 B.n157 B.n156 10.6151
R2164 B.n160 B.n157 10.6151
R2165 B.n161 B.n160 10.6151
R2166 B.n164 B.n161 10.6151
R2167 B.n165 B.n164 10.6151
R2168 B.n168 B.n165 10.6151
R2169 B.n169 B.n168 10.6151
R2170 B.n172 B.n169 10.6151
R2171 B.n173 B.n172 10.6151
R2172 B.n176 B.n173 10.6151
R2173 B.n177 B.n176 10.6151
R2174 B.n180 B.n177 10.6151
R2175 B.n181 B.n180 10.6151
R2176 B.n184 B.n181 10.6151
R2177 B.n185 B.n184 10.6151
R2178 B.n188 B.n185 10.6151
R2179 B.n189 B.n188 10.6151
R2180 B.n192 B.n189 10.6151
R2181 B.n193 B.n192 10.6151
R2182 B.n196 B.n193 10.6151
R2183 B.n197 B.n196 10.6151
R2184 B.n200 B.n197 10.6151
R2185 B.n201 B.n200 10.6151
R2186 B.n204 B.n201 10.6151
R2187 B.n205 B.n204 10.6151
R2188 B.n208 B.n205 10.6151
R2189 B.n209 B.n208 10.6151
R2190 B.n212 B.n209 10.6151
R2191 B.n213 B.n212 10.6151
R2192 B.n216 B.n213 10.6151
R2193 B.n217 B.n216 10.6151
R2194 B.n220 B.n217 10.6151
R2195 B.n221 B.n220 10.6151
R2196 B.n224 B.n221 10.6151
R2197 B.n225 B.n224 10.6151
R2198 B.n228 B.n225 10.6151
R2199 B.n229 B.n228 10.6151
R2200 B.n232 B.n229 10.6151
R2201 B.n237 B.n234 10.6151
R2202 B.n238 B.n237 10.6151
R2203 B.n241 B.n238 10.6151
R2204 B.n242 B.n241 10.6151
R2205 B.n245 B.n242 10.6151
R2206 B.n246 B.n245 10.6151
R2207 B.n249 B.n246 10.6151
R2208 B.n250 B.n249 10.6151
R2209 B.n253 B.n250 10.6151
R2210 B.n258 B.n255 10.6151
R2211 B.n259 B.n258 10.6151
R2212 B.n262 B.n259 10.6151
R2213 B.n263 B.n262 10.6151
R2214 B.n266 B.n263 10.6151
R2215 B.n267 B.n266 10.6151
R2216 B.n270 B.n267 10.6151
R2217 B.n271 B.n270 10.6151
R2218 B.n274 B.n271 10.6151
R2219 B.n275 B.n274 10.6151
R2220 B.n278 B.n275 10.6151
R2221 B.n279 B.n278 10.6151
R2222 B.n282 B.n279 10.6151
R2223 B.n283 B.n282 10.6151
R2224 B.n286 B.n283 10.6151
R2225 B.n287 B.n286 10.6151
R2226 B.n290 B.n287 10.6151
R2227 B.n291 B.n290 10.6151
R2228 B.n294 B.n291 10.6151
R2229 B.n295 B.n294 10.6151
R2230 B.n298 B.n295 10.6151
R2231 B.n299 B.n298 10.6151
R2232 B.n302 B.n299 10.6151
R2233 B.n303 B.n302 10.6151
R2234 B.n306 B.n303 10.6151
R2235 B.n307 B.n306 10.6151
R2236 B.n310 B.n307 10.6151
R2237 B.n311 B.n310 10.6151
R2238 B.n314 B.n311 10.6151
R2239 B.n315 B.n314 10.6151
R2240 B.n318 B.n315 10.6151
R2241 B.n319 B.n318 10.6151
R2242 B.n322 B.n319 10.6151
R2243 B.n323 B.n322 10.6151
R2244 B.n326 B.n323 10.6151
R2245 B.n327 B.n326 10.6151
R2246 B.n330 B.n327 10.6151
R2247 B.n331 B.n330 10.6151
R2248 B.n334 B.n331 10.6151
R2249 B.n335 B.n334 10.6151
R2250 B.n338 B.n335 10.6151
R2251 B.n339 B.n338 10.6151
R2252 B.n342 B.n339 10.6151
R2253 B.n343 B.n342 10.6151
R2254 B.n346 B.n343 10.6151
R2255 B.n348 B.n346 10.6151
R2256 B.n349 B.n348 10.6151
R2257 B.n880 B.n349 10.6151
R2258 B.n706 B.n705 10.6151
R2259 B.n706 B.n421 10.6151
R2260 B.n716 B.n421 10.6151
R2261 B.n717 B.n716 10.6151
R2262 B.n718 B.n717 10.6151
R2263 B.n718 B.n413 10.6151
R2264 B.n728 B.n413 10.6151
R2265 B.n729 B.n728 10.6151
R2266 B.n730 B.n729 10.6151
R2267 B.n730 B.n405 10.6151
R2268 B.n740 B.n405 10.6151
R2269 B.n741 B.n740 10.6151
R2270 B.n742 B.n741 10.6151
R2271 B.n742 B.n398 10.6151
R2272 B.n753 B.n398 10.6151
R2273 B.n754 B.n753 10.6151
R2274 B.n755 B.n754 10.6151
R2275 B.n755 B.n389 10.6151
R2276 B.n765 B.n389 10.6151
R2277 B.n766 B.n765 10.6151
R2278 B.n767 B.n766 10.6151
R2279 B.n767 B.n382 10.6151
R2280 B.n777 B.n382 10.6151
R2281 B.n778 B.n777 10.6151
R2282 B.n779 B.n778 10.6151
R2283 B.n779 B.n374 10.6151
R2284 B.n789 B.n374 10.6151
R2285 B.n790 B.n789 10.6151
R2286 B.n791 B.n790 10.6151
R2287 B.n791 B.n366 10.6151
R2288 B.n801 B.n366 10.6151
R2289 B.n802 B.n801 10.6151
R2290 B.n803 B.n802 10.6151
R2291 B.n803 B.n357 10.6151
R2292 B.n813 B.n357 10.6151
R2293 B.n814 B.n813 10.6151
R2294 B.n816 B.n814 10.6151
R2295 B.n816 B.n815 10.6151
R2296 B.n815 B.n350 10.6151
R2297 B.n827 B.n350 10.6151
R2298 B.n828 B.n827 10.6151
R2299 B.n829 B.n828 10.6151
R2300 B.n830 B.n829 10.6151
R2301 B.n832 B.n830 10.6151
R2302 B.n833 B.n832 10.6151
R2303 B.n834 B.n833 10.6151
R2304 B.n835 B.n834 10.6151
R2305 B.n837 B.n835 10.6151
R2306 B.n838 B.n837 10.6151
R2307 B.n839 B.n838 10.6151
R2308 B.n840 B.n839 10.6151
R2309 B.n842 B.n840 10.6151
R2310 B.n843 B.n842 10.6151
R2311 B.n844 B.n843 10.6151
R2312 B.n845 B.n844 10.6151
R2313 B.n847 B.n845 10.6151
R2314 B.n848 B.n847 10.6151
R2315 B.n849 B.n848 10.6151
R2316 B.n850 B.n849 10.6151
R2317 B.n852 B.n850 10.6151
R2318 B.n853 B.n852 10.6151
R2319 B.n854 B.n853 10.6151
R2320 B.n855 B.n854 10.6151
R2321 B.n857 B.n855 10.6151
R2322 B.n858 B.n857 10.6151
R2323 B.n859 B.n858 10.6151
R2324 B.n860 B.n859 10.6151
R2325 B.n862 B.n860 10.6151
R2326 B.n863 B.n862 10.6151
R2327 B.n864 B.n863 10.6151
R2328 B.n865 B.n864 10.6151
R2329 B.n867 B.n865 10.6151
R2330 B.n868 B.n867 10.6151
R2331 B.n869 B.n868 10.6151
R2332 B.n870 B.n869 10.6151
R2333 B.n872 B.n870 10.6151
R2334 B.n873 B.n872 10.6151
R2335 B.n874 B.n873 10.6151
R2336 B.n875 B.n874 10.6151
R2337 B.n877 B.n875 10.6151
R2338 B.n878 B.n877 10.6151
R2339 B.n879 B.n878 10.6151
R2340 B.n699 B.n698 10.6151
R2341 B.n698 B.n697 10.6151
R2342 B.n697 B.n696 10.6151
R2343 B.n696 B.n694 10.6151
R2344 B.n694 B.n691 10.6151
R2345 B.n691 B.n690 10.6151
R2346 B.n690 B.n687 10.6151
R2347 B.n687 B.n686 10.6151
R2348 B.n686 B.n683 10.6151
R2349 B.n683 B.n682 10.6151
R2350 B.n682 B.n679 10.6151
R2351 B.n679 B.n678 10.6151
R2352 B.n678 B.n675 10.6151
R2353 B.n675 B.n674 10.6151
R2354 B.n674 B.n671 10.6151
R2355 B.n671 B.n670 10.6151
R2356 B.n670 B.n667 10.6151
R2357 B.n667 B.n666 10.6151
R2358 B.n666 B.n663 10.6151
R2359 B.n663 B.n662 10.6151
R2360 B.n662 B.n659 10.6151
R2361 B.n659 B.n658 10.6151
R2362 B.n658 B.n655 10.6151
R2363 B.n655 B.n654 10.6151
R2364 B.n654 B.n651 10.6151
R2365 B.n651 B.n650 10.6151
R2366 B.n650 B.n647 10.6151
R2367 B.n647 B.n646 10.6151
R2368 B.n646 B.n643 10.6151
R2369 B.n643 B.n642 10.6151
R2370 B.n642 B.n639 10.6151
R2371 B.n639 B.n638 10.6151
R2372 B.n638 B.n635 10.6151
R2373 B.n635 B.n634 10.6151
R2374 B.n634 B.n631 10.6151
R2375 B.n631 B.n630 10.6151
R2376 B.n630 B.n627 10.6151
R2377 B.n627 B.n626 10.6151
R2378 B.n626 B.n623 10.6151
R2379 B.n623 B.n622 10.6151
R2380 B.n622 B.n619 10.6151
R2381 B.n619 B.n618 10.6151
R2382 B.n618 B.n615 10.6151
R2383 B.n615 B.n614 10.6151
R2384 B.n614 B.n611 10.6151
R2385 B.n611 B.n610 10.6151
R2386 B.n610 B.n607 10.6151
R2387 B.n607 B.n606 10.6151
R2388 B.n603 B.n602 10.6151
R2389 B.n602 B.n599 10.6151
R2390 B.n599 B.n598 10.6151
R2391 B.n598 B.n595 10.6151
R2392 B.n595 B.n594 10.6151
R2393 B.n594 B.n591 10.6151
R2394 B.n591 B.n590 10.6151
R2395 B.n590 B.n587 10.6151
R2396 B.n587 B.n586 10.6151
R2397 B.n583 B.n582 10.6151
R2398 B.n582 B.n579 10.6151
R2399 B.n579 B.n578 10.6151
R2400 B.n578 B.n575 10.6151
R2401 B.n575 B.n574 10.6151
R2402 B.n574 B.n571 10.6151
R2403 B.n571 B.n570 10.6151
R2404 B.n570 B.n567 10.6151
R2405 B.n567 B.n566 10.6151
R2406 B.n566 B.n563 10.6151
R2407 B.n563 B.n562 10.6151
R2408 B.n562 B.n559 10.6151
R2409 B.n559 B.n558 10.6151
R2410 B.n558 B.n555 10.6151
R2411 B.n555 B.n554 10.6151
R2412 B.n554 B.n551 10.6151
R2413 B.n551 B.n550 10.6151
R2414 B.n550 B.n547 10.6151
R2415 B.n547 B.n546 10.6151
R2416 B.n546 B.n543 10.6151
R2417 B.n543 B.n542 10.6151
R2418 B.n542 B.n539 10.6151
R2419 B.n539 B.n538 10.6151
R2420 B.n538 B.n535 10.6151
R2421 B.n535 B.n534 10.6151
R2422 B.n534 B.n531 10.6151
R2423 B.n531 B.n530 10.6151
R2424 B.n530 B.n527 10.6151
R2425 B.n527 B.n526 10.6151
R2426 B.n526 B.n523 10.6151
R2427 B.n523 B.n522 10.6151
R2428 B.n522 B.n519 10.6151
R2429 B.n519 B.n518 10.6151
R2430 B.n518 B.n515 10.6151
R2431 B.n515 B.n514 10.6151
R2432 B.n514 B.n511 10.6151
R2433 B.n511 B.n510 10.6151
R2434 B.n510 B.n507 10.6151
R2435 B.n507 B.n506 10.6151
R2436 B.n506 B.n503 10.6151
R2437 B.n503 B.n502 10.6151
R2438 B.n502 B.n499 10.6151
R2439 B.n499 B.n498 10.6151
R2440 B.n498 B.n495 10.6151
R2441 B.n495 B.n494 10.6151
R2442 B.n494 B.n491 10.6151
R2443 B.n491 B.n429 10.6151
R2444 B.n704 B.n429 10.6151
R2445 B.n710 B.n425 10.6151
R2446 B.n711 B.n710 10.6151
R2447 B.n712 B.n711 10.6151
R2448 B.n712 B.n417 10.6151
R2449 B.n722 B.n417 10.6151
R2450 B.n723 B.n722 10.6151
R2451 B.n724 B.n723 10.6151
R2452 B.n724 B.n409 10.6151
R2453 B.n734 B.n409 10.6151
R2454 B.n735 B.n734 10.6151
R2455 B.n736 B.n735 10.6151
R2456 B.n736 B.n401 10.6151
R2457 B.n747 B.n401 10.6151
R2458 B.n748 B.n747 10.6151
R2459 B.n749 B.n748 10.6151
R2460 B.n749 B.n394 10.6151
R2461 B.n759 B.n394 10.6151
R2462 B.n760 B.n759 10.6151
R2463 B.n761 B.n760 10.6151
R2464 B.n761 B.n386 10.6151
R2465 B.n771 B.n386 10.6151
R2466 B.n772 B.n771 10.6151
R2467 B.n773 B.n772 10.6151
R2468 B.n773 B.n378 10.6151
R2469 B.n783 B.n378 10.6151
R2470 B.n784 B.n783 10.6151
R2471 B.n785 B.n784 10.6151
R2472 B.n785 B.n370 10.6151
R2473 B.n795 B.n370 10.6151
R2474 B.n796 B.n795 10.6151
R2475 B.n797 B.n796 10.6151
R2476 B.n797 B.n362 10.6151
R2477 B.n807 B.n362 10.6151
R2478 B.n808 B.n807 10.6151
R2479 B.n809 B.n808 10.6151
R2480 B.n809 B.n354 10.6151
R2481 B.n820 B.n354 10.6151
R2482 B.n821 B.n820 10.6151
R2483 B.n822 B.n821 10.6151
R2484 B.n822 B.n0 10.6151
R2485 B.n961 B.n1 10.6151
R2486 B.n961 B.n960 10.6151
R2487 B.n960 B.n959 10.6151
R2488 B.n959 B.n10 10.6151
R2489 B.n953 B.n10 10.6151
R2490 B.n953 B.n952 10.6151
R2491 B.n952 B.n951 10.6151
R2492 B.n951 B.n17 10.6151
R2493 B.n945 B.n17 10.6151
R2494 B.n945 B.n944 10.6151
R2495 B.n944 B.n943 10.6151
R2496 B.n943 B.n24 10.6151
R2497 B.n937 B.n24 10.6151
R2498 B.n937 B.n936 10.6151
R2499 B.n936 B.n935 10.6151
R2500 B.n935 B.n31 10.6151
R2501 B.n929 B.n31 10.6151
R2502 B.n929 B.n928 10.6151
R2503 B.n928 B.n927 10.6151
R2504 B.n927 B.n38 10.6151
R2505 B.n921 B.n38 10.6151
R2506 B.n921 B.n920 10.6151
R2507 B.n920 B.n919 10.6151
R2508 B.n919 B.n45 10.6151
R2509 B.n913 B.n45 10.6151
R2510 B.n913 B.n912 10.6151
R2511 B.n912 B.n911 10.6151
R2512 B.n911 B.n51 10.6151
R2513 B.n905 B.n51 10.6151
R2514 B.n905 B.n904 10.6151
R2515 B.n904 B.n903 10.6151
R2516 B.n903 B.n59 10.6151
R2517 B.n897 B.n59 10.6151
R2518 B.n897 B.n896 10.6151
R2519 B.n896 B.n895 10.6151
R2520 B.n895 B.n66 10.6151
R2521 B.n889 B.n66 10.6151
R2522 B.n889 B.n888 10.6151
R2523 B.n888 B.n887 10.6151
R2524 B.n887 B.n73 10.6151
R2525 B.n233 B.n232 9.36635
R2526 B.n255 B.n254 9.36635
R2527 B.n606 B.n487 9.36635
R2528 B.n583 B.n490 9.36635
R2529 B.n392 B.t2 5.52675
R2530 B.n799 B.t1 5.52675
R2531 B.t4 B.n947 5.52675
R2532 B.t3 B.n924 5.52675
R2533 B.n967 B.n0 2.81026
R2534 B.n967 B.n1 2.81026
R2535 B.t11 B.n415 2.211
R2536 B.t15 B.n64 2.211
R2537 B.n234 B.n233 1.24928
R2538 B.n254 B.n253 1.24928
R2539 B.n603 B.n487 1.24928
R2540 B.n586 B.n490 1.24928
R2541 VN.n7 VN.t5 263.575
R2542 VN.n34 VN.t7 263.575
R2543 VN.n12 VN.t1 228.951
R2544 VN.n6 VN.t4 228.951
R2545 VN.n18 VN.t0 228.951
R2546 VN.n25 VN.t3 228.951
R2547 VN.n39 VN.t8 228.951
R2548 VN.n33 VN.t9 228.951
R2549 VN.n45 VN.t2 228.951
R2550 VN.n52 VN.t6 228.951
R2551 VN.n26 VN.n25 174.024
R2552 VN.n53 VN.n52 174.024
R2553 VN.n51 VN.n27 161.3
R2554 VN.n50 VN.n49 161.3
R2555 VN.n48 VN.n28 161.3
R2556 VN.n47 VN.n46 161.3
R2557 VN.n44 VN.n29 161.3
R2558 VN.n43 VN.n42 161.3
R2559 VN.n41 VN.n30 161.3
R2560 VN.n40 VN.n39 161.3
R2561 VN.n38 VN.n31 161.3
R2562 VN.n37 VN.n36 161.3
R2563 VN.n35 VN.n32 161.3
R2564 VN.n24 VN.n0 161.3
R2565 VN.n23 VN.n22 161.3
R2566 VN.n21 VN.n1 161.3
R2567 VN.n20 VN.n19 161.3
R2568 VN.n17 VN.n2 161.3
R2569 VN.n16 VN.n15 161.3
R2570 VN.n14 VN.n3 161.3
R2571 VN.n13 VN.n12 161.3
R2572 VN.n11 VN.n4 161.3
R2573 VN.n10 VN.n9 161.3
R2574 VN.n8 VN.n5 161.3
R2575 VN.n23 VN.n1 56.5193
R2576 VN.n50 VN.n28 56.5193
R2577 VN VN.n53 49.688
R2578 VN.n7 VN.n6 48.4385
R2579 VN.n34 VN.n33 48.4385
R2580 VN.n11 VN.n10 46.8066
R2581 VN.n16 VN.n3 46.8066
R2582 VN.n38 VN.n37 46.8066
R2583 VN.n43 VN.n30 46.8066
R2584 VN.n10 VN.n5 34.1802
R2585 VN.n17 VN.n16 34.1802
R2586 VN.n37 VN.n32 34.1802
R2587 VN.n44 VN.n43 34.1802
R2588 VN.n12 VN.n11 24.4675
R2589 VN.n12 VN.n3 24.4675
R2590 VN.n19 VN.n1 24.4675
R2591 VN.n24 VN.n23 24.4675
R2592 VN.n39 VN.n30 24.4675
R2593 VN.n39 VN.n38 24.4675
R2594 VN.n46 VN.n28 24.4675
R2595 VN.n51 VN.n50 24.4675
R2596 VN.n6 VN.n5 18.1061
R2597 VN.n18 VN.n17 18.1061
R2598 VN.n33 VN.n32 18.1061
R2599 VN.n45 VN.n44 18.1061
R2600 VN.n35 VN.n34 17.6128
R2601 VN.n8 VN.n7 17.6128
R2602 VN.n25 VN.n24 11.7447
R2603 VN.n52 VN.n51 11.7447
R2604 VN.n19 VN.n18 6.36192
R2605 VN.n46 VN.n45 6.36192
R2606 VN.n53 VN.n27 0.189894
R2607 VN.n49 VN.n27 0.189894
R2608 VN.n49 VN.n48 0.189894
R2609 VN.n48 VN.n47 0.189894
R2610 VN.n47 VN.n29 0.189894
R2611 VN.n42 VN.n29 0.189894
R2612 VN.n42 VN.n41 0.189894
R2613 VN.n41 VN.n40 0.189894
R2614 VN.n40 VN.n31 0.189894
R2615 VN.n36 VN.n31 0.189894
R2616 VN.n36 VN.n35 0.189894
R2617 VN.n9 VN.n8 0.189894
R2618 VN.n9 VN.n4 0.189894
R2619 VN.n13 VN.n4 0.189894
R2620 VN.n14 VN.n13 0.189894
R2621 VN.n15 VN.n14 0.189894
R2622 VN.n15 VN.n2 0.189894
R2623 VN.n20 VN.n2 0.189894
R2624 VN.n21 VN.n20 0.189894
R2625 VN.n22 VN.n21 0.189894
R2626 VN.n22 VN.n0 0.189894
R2627 VN.n26 VN.n0 0.189894
R2628 VN VN.n26 0.0516364
R2629 VDD2.n161 VDD2.n85 289.615
R2630 VDD2.n76 VDD2.n0 289.615
R2631 VDD2.n162 VDD2.n161 185
R2632 VDD2.n160 VDD2.n159 185
R2633 VDD2.n158 VDD2.n88 185
R2634 VDD2.n92 VDD2.n89 185
R2635 VDD2.n153 VDD2.n152 185
R2636 VDD2.n151 VDD2.n150 185
R2637 VDD2.n94 VDD2.n93 185
R2638 VDD2.n145 VDD2.n144 185
R2639 VDD2.n143 VDD2.n142 185
R2640 VDD2.n98 VDD2.n97 185
R2641 VDD2.n137 VDD2.n136 185
R2642 VDD2.n135 VDD2.n134 185
R2643 VDD2.n102 VDD2.n101 185
R2644 VDD2.n129 VDD2.n128 185
R2645 VDD2.n127 VDD2.n126 185
R2646 VDD2.n106 VDD2.n105 185
R2647 VDD2.n121 VDD2.n120 185
R2648 VDD2.n119 VDD2.n118 185
R2649 VDD2.n110 VDD2.n109 185
R2650 VDD2.n113 VDD2.n112 185
R2651 VDD2.n27 VDD2.n26 185
R2652 VDD2.n24 VDD2.n23 185
R2653 VDD2.n33 VDD2.n32 185
R2654 VDD2.n35 VDD2.n34 185
R2655 VDD2.n20 VDD2.n19 185
R2656 VDD2.n41 VDD2.n40 185
R2657 VDD2.n43 VDD2.n42 185
R2658 VDD2.n16 VDD2.n15 185
R2659 VDD2.n49 VDD2.n48 185
R2660 VDD2.n51 VDD2.n50 185
R2661 VDD2.n12 VDD2.n11 185
R2662 VDD2.n57 VDD2.n56 185
R2663 VDD2.n59 VDD2.n58 185
R2664 VDD2.n8 VDD2.n7 185
R2665 VDD2.n65 VDD2.n64 185
R2666 VDD2.n68 VDD2.n67 185
R2667 VDD2.n66 VDD2.n4 185
R2668 VDD2.n73 VDD2.n3 185
R2669 VDD2.n75 VDD2.n74 185
R2670 VDD2.n77 VDD2.n76 185
R2671 VDD2.t3 VDD2.n111 147.659
R2672 VDD2.t4 VDD2.n25 147.659
R2673 VDD2.n161 VDD2.n160 104.615
R2674 VDD2.n160 VDD2.n88 104.615
R2675 VDD2.n92 VDD2.n88 104.615
R2676 VDD2.n152 VDD2.n92 104.615
R2677 VDD2.n152 VDD2.n151 104.615
R2678 VDD2.n151 VDD2.n93 104.615
R2679 VDD2.n144 VDD2.n93 104.615
R2680 VDD2.n144 VDD2.n143 104.615
R2681 VDD2.n143 VDD2.n97 104.615
R2682 VDD2.n136 VDD2.n97 104.615
R2683 VDD2.n136 VDD2.n135 104.615
R2684 VDD2.n135 VDD2.n101 104.615
R2685 VDD2.n128 VDD2.n101 104.615
R2686 VDD2.n128 VDD2.n127 104.615
R2687 VDD2.n127 VDD2.n105 104.615
R2688 VDD2.n120 VDD2.n105 104.615
R2689 VDD2.n120 VDD2.n119 104.615
R2690 VDD2.n119 VDD2.n109 104.615
R2691 VDD2.n112 VDD2.n109 104.615
R2692 VDD2.n26 VDD2.n23 104.615
R2693 VDD2.n33 VDD2.n23 104.615
R2694 VDD2.n34 VDD2.n33 104.615
R2695 VDD2.n34 VDD2.n19 104.615
R2696 VDD2.n41 VDD2.n19 104.615
R2697 VDD2.n42 VDD2.n41 104.615
R2698 VDD2.n42 VDD2.n15 104.615
R2699 VDD2.n49 VDD2.n15 104.615
R2700 VDD2.n50 VDD2.n49 104.615
R2701 VDD2.n50 VDD2.n11 104.615
R2702 VDD2.n57 VDD2.n11 104.615
R2703 VDD2.n58 VDD2.n57 104.615
R2704 VDD2.n58 VDD2.n7 104.615
R2705 VDD2.n65 VDD2.n7 104.615
R2706 VDD2.n67 VDD2.n65 104.615
R2707 VDD2.n67 VDD2.n66 104.615
R2708 VDD2.n66 VDD2.n3 104.615
R2709 VDD2.n75 VDD2.n3 104.615
R2710 VDD2.n76 VDD2.n75 104.615
R2711 VDD2.n84 VDD2.n83 61.8807
R2712 VDD2 VDD2.n169 61.8778
R2713 VDD2.n168 VDD2.n167 60.7272
R2714 VDD2.n82 VDD2.n81 60.727
R2715 VDD2.n112 VDD2.t3 52.3082
R2716 VDD2.n26 VDD2.t4 52.3082
R2717 VDD2.n82 VDD2.n80 50.2823
R2718 VDD2.n166 VDD2.n165 48.6702
R2719 VDD2.n166 VDD2.n84 43.9847
R2720 VDD2.n113 VDD2.n111 15.6677
R2721 VDD2.n27 VDD2.n25 15.6677
R2722 VDD2.n159 VDD2.n158 13.1884
R2723 VDD2.n74 VDD2.n73 13.1884
R2724 VDD2.n162 VDD2.n87 12.8005
R2725 VDD2.n157 VDD2.n89 12.8005
R2726 VDD2.n114 VDD2.n110 12.8005
R2727 VDD2.n28 VDD2.n24 12.8005
R2728 VDD2.n72 VDD2.n4 12.8005
R2729 VDD2.n77 VDD2.n2 12.8005
R2730 VDD2.n163 VDD2.n85 12.0247
R2731 VDD2.n154 VDD2.n153 12.0247
R2732 VDD2.n118 VDD2.n117 12.0247
R2733 VDD2.n32 VDD2.n31 12.0247
R2734 VDD2.n69 VDD2.n68 12.0247
R2735 VDD2.n78 VDD2.n0 12.0247
R2736 VDD2.n150 VDD2.n91 11.249
R2737 VDD2.n121 VDD2.n108 11.249
R2738 VDD2.n35 VDD2.n22 11.249
R2739 VDD2.n64 VDD2.n6 11.249
R2740 VDD2.n149 VDD2.n94 10.4732
R2741 VDD2.n122 VDD2.n106 10.4732
R2742 VDD2.n36 VDD2.n20 10.4732
R2743 VDD2.n63 VDD2.n8 10.4732
R2744 VDD2.n146 VDD2.n145 9.69747
R2745 VDD2.n126 VDD2.n125 9.69747
R2746 VDD2.n40 VDD2.n39 9.69747
R2747 VDD2.n60 VDD2.n59 9.69747
R2748 VDD2.n165 VDD2.n164 9.45567
R2749 VDD2.n80 VDD2.n79 9.45567
R2750 VDD2.n139 VDD2.n138 9.3005
R2751 VDD2.n141 VDD2.n140 9.3005
R2752 VDD2.n96 VDD2.n95 9.3005
R2753 VDD2.n147 VDD2.n146 9.3005
R2754 VDD2.n149 VDD2.n148 9.3005
R2755 VDD2.n91 VDD2.n90 9.3005
R2756 VDD2.n155 VDD2.n154 9.3005
R2757 VDD2.n157 VDD2.n156 9.3005
R2758 VDD2.n164 VDD2.n163 9.3005
R2759 VDD2.n87 VDD2.n86 9.3005
R2760 VDD2.n100 VDD2.n99 9.3005
R2761 VDD2.n133 VDD2.n132 9.3005
R2762 VDD2.n131 VDD2.n130 9.3005
R2763 VDD2.n104 VDD2.n103 9.3005
R2764 VDD2.n125 VDD2.n124 9.3005
R2765 VDD2.n123 VDD2.n122 9.3005
R2766 VDD2.n108 VDD2.n107 9.3005
R2767 VDD2.n117 VDD2.n116 9.3005
R2768 VDD2.n115 VDD2.n114 9.3005
R2769 VDD2.n79 VDD2.n78 9.3005
R2770 VDD2.n2 VDD2.n1 9.3005
R2771 VDD2.n47 VDD2.n46 9.3005
R2772 VDD2.n45 VDD2.n44 9.3005
R2773 VDD2.n18 VDD2.n17 9.3005
R2774 VDD2.n39 VDD2.n38 9.3005
R2775 VDD2.n37 VDD2.n36 9.3005
R2776 VDD2.n22 VDD2.n21 9.3005
R2777 VDD2.n31 VDD2.n30 9.3005
R2778 VDD2.n29 VDD2.n28 9.3005
R2779 VDD2.n14 VDD2.n13 9.3005
R2780 VDD2.n53 VDD2.n52 9.3005
R2781 VDD2.n55 VDD2.n54 9.3005
R2782 VDD2.n10 VDD2.n9 9.3005
R2783 VDD2.n61 VDD2.n60 9.3005
R2784 VDD2.n63 VDD2.n62 9.3005
R2785 VDD2.n6 VDD2.n5 9.3005
R2786 VDD2.n70 VDD2.n69 9.3005
R2787 VDD2.n72 VDD2.n71 9.3005
R2788 VDD2.n142 VDD2.n96 8.92171
R2789 VDD2.n129 VDD2.n104 8.92171
R2790 VDD2.n43 VDD2.n18 8.92171
R2791 VDD2.n56 VDD2.n10 8.92171
R2792 VDD2.n141 VDD2.n98 8.14595
R2793 VDD2.n130 VDD2.n102 8.14595
R2794 VDD2.n44 VDD2.n16 8.14595
R2795 VDD2.n55 VDD2.n12 8.14595
R2796 VDD2.n138 VDD2.n137 7.3702
R2797 VDD2.n134 VDD2.n133 7.3702
R2798 VDD2.n48 VDD2.n47 7.3702
R2799 VDD2.n52 VDD2.n51 7.3702
R2800 VDD2.n137 VDD2.n100 6.59444
R2801 VDD2.n134 VDD2.n100 6.59444
R2802 VDD2.n48 VDD2.n14 6.59444
R2803 VDD2.n51 VDD2.n14 6.59444
R2804 VDD2.n138 VDD2.n98 5.81868
R2805 VDD2.n133 VDD2.n102 5.81868
R2806 VDD2.n47 VDD2.n16 5.81868
R2807 VDD2.n52 VDD2.n12 5.81868
R2808 VDD2.n142 VDD2.n141 5.04292
R2809 VDD2.n130 VDD2.n129 5.04292
R2810 VDD2.n44 VDD2.n43 5.04292
R2811 VDD2.n56 VDD2.n55 5.04292
R2812 VDD2.n115 VDD2.n111 4.38563
R2813 VDD2.n29 VDD2.n25 4.38563
R2814 VDD2.n145 VDD2.n96 4.26717
R2815 VDD2.n126 VDD2.n104 4.26717
R2816 VDD2.n40 VDD2.n18 4.26717
R2817 VDD2.n59 VDD2.n10 4.26717
R2818 VDD2.n146 VDD2.n94 3.49141
R2819 VDD2.n125 VDD2.n106 3.49141
R2820 VDD2.n39 VDD2.n20 3.49141
R2821 VDD2.n60 VDD2.n8 3.49141
R2822 VDD2.n150 VDD2.n149 2.71565
R2823 VDD2.n122 VDD2.n121 2.71565
R2824 VDD2.n36 VDD2.n35 2.71565
R2825 VDD2.n64 VDD2.n63 2.71565
R2826 VDD2.n165 VDD2.n85 1.93989
R2827 VDD2.n153 VDD2.n91 1.93989
R2828 VDD2.n118 VDD2.n108 1.93989
R2829 VDD2.n32 VDD2.n22 1.93989
R2830 VDD2.n68 VDD2.n6 1.93989
R2831 VDD2.n80 VDD2.n0 1.93989
R2832 VDD2.n168 VDD2.n166 1.61257
R2833 VDD2.n169 VDD2.t0 1.35388
R2834 VDD2.n169 VDD2.t2 1.35388
R2835 VDD2.n167 VDD2.t7 1.35388
R2836 VDD2.n167 VDD2.t1 1.35388
R2837 VDD2.n83 VDD2.t9 1.35388
R2838 VDD2.n83 VDD2.t6 1.35388
R2839 VDD2.n81 VDD2.t5 1.35388
R2840 VDD2.n81 VDD2.t8 1.35388
R2841 VDD2.n163 VDD2.n162 1.16414
R2842 VDD2.n154 VDD2.n89 1.16414
R2843 VDD2.n117 VDD2.n110 1.16414
R2844 VDD2.n31 VDD2.n24 1.16414
R2845 VDD2.n69 VDD2.n4 1.16414
R2846 VDD2.n78 VDD2.n77 1.16414
R2847 VDD2 VDD2.n168 0.461707
R2848 VDD2.n159 VDD2.n87 0.388379
R2849 VDD2.n158 VDD2.n157 0.388379
R2850 VDD2.n114 VDD2.n113 0.388379
R2851 VDD2.n28 VDD2.n27 0.388379
R2852 VDD2.n73 VDD2.n72 0.388379
R2853 VDD2.n74 VDD2.n2 0.388379
R2854 VDD2.n84 VDD2.n82 0.348171
R2855 VDD2.n164 VDD2.n86 0.155672
R2856 VDD2.n156 VDD2.n86 0.155672
R2857 VDD2.n156 VDD2.n155 0.155672
R2858 VDD2.n155 VDD2.n90 0.155672
R2859 VDD2.n148 VDD2.n90 0.155672
R2860 VDD2.n148 VDD2.n147 0.155672
R2861 VDD2.n147 VDD2.n95 0.155672
R2862 VDD2.n140 VDD2.n95 0.155672
R2863 VDD2.n140 VDD2.n139 0.155672
R2864 VDD2.n139 VDD2.n99 0.155672
R2865 VDD2.n132 VDD2.n99 0.155672
R2866 VDD2.n132 VDD2.n131 0.155672
R2867 VDD2.n131 VDD2.n103 0.155672
R2868 VDD2.n124 VDD2.n103 0.155672
R2869 VDD2.n124 VDD2.n123 0.155672
R2870 VDD2.n123 VDD2.n107 0.155672
R2871 VDD2.n116 VDD2.n107 0.155672
R2872 VDD2.n116 VDD2.n115 0.155672
R2873 VDD2.n30 VDD2.n29 0.155672
R2874 VDD2.n30 VDD2.n21 0.155672
R2875 VDD2.n37 VDD2.n21 0.155672
R2876 VDD2.n38 VDD2.n37 0.155672
R2877 VDD2.n38 VDD2.n17 0.155672
R2878 VDD2.n45 VDD2.n17 0.155672
R2879 VDD2.n46 VDD2.n45 0.155672
R2880 VDD2.n46 VDD2.n13 0.155672
R2881 VDD2.n53 VDD2.n13 0.155672
R2882 VDD2.n54 VDD2.n53 0.155672
R2883 VDD2.n54 VDD2.n9 0.155672
R2884 VDD2.n61 VDD2.n9 0.155672
R2885 VDD2.n62 VDD2.n61 0.155672
R2886 VDD2.n62 VDD2.n5 0.155672
R2887 VDD2.n70 VDD2.n5 0.155672
R2888 VDD2.n71 VDD2.n70 0.155672
R2889 VDD2.n71 VDD2.n1 0.155672
R2890 VDD2.n79 VDD2.n1 0.155672
C0 VDD2 VP 0.448712f
C1 VP VN 7.32071f
C2 VDD2 VN 11.276401f
C3 VP VTAIL 11.3834f
C4 VDD2 VTAIL 12.509099f
C5 VN VTAIL 11.368999f
C6 VP VDD1 11.5695f
C7 VDD2 VDD1 1.48537f
C8 VN VDD1 0.150892f
C9 VTAIL VDD1 12.4678f
C10 VDD2 B 6.430647f
C11 VDD1 B 6.405116f
C12 VTAIL B 8.342573f
C13 VN B 13.43029f
C14 VP B 11.719082f
C15 VDD2.n0 B 0.028317f
C16 VDD2.n1 B 0.022404f
C17 VDD2.n2 B 0.012039f
C18 VDD2.n3 B 0.028456f
C19 VDD2.n4 B 0.012747f
C20 VDD2.n5 B 0.022404f
C21 VDD2.n6 B 0.012039f
C22 VDD2.n7 B 0.028456f
C23 VDD2.n8 B 0.012747f
C24 VDD2.n9 B 0.022404f
C25 VDD2.n10 B 0.012039f
C26 VDD2.n11 B 0.028456f
C27 VDD2.n12 B 0.012747f
C28 VDD2.n13 B 0.022404f
C29 VDD2.n14 B 0.012039f
C30 VDD2.n15 B 0.028456f
C31 VDD2.n16 B 0.012747f
C32 VDD2.n17 B 0.022404f
C33 VDD2.n18 B 0.012039f
C34 VDD2.n19 B 0.028456f
C35 VDD2.n20 B 0.012747f
C36 VDD2.n21 B 0.022404f
C37 VDD2.n22 B 0.012039f
C38 VDD2.n23 B 0.028456f
C39 VDD2.n24 B 0.012747f
C40 VDD2.n25 B 0.144047f
C41 VDD2.t4 B 0.046892f
C42 VDD2.n26 B 0.021342f
C43 VDD2.n27 B 0.01681f
C44 VDD2.n28 B 0.012039f
C45 VDD2.n29 B 1.41966f
C46 VDD2.n30 B 0.022404f
C47 VDD2.n31 B 0.012039f
C48 VDD2.n32 B 0.012747f
C49 VDD2.n33 B 0.028456f
C50 VDD2.n34 B 0.028456f
C51 VDD2.n35 B 0.012747f
C52 VDD2.n36 B 0.012039f
C53 VDD2.n37 B 0.022404f
C54 VDD2.n38 B 0.022404f
C55 VDD2.n39 B 0.012039f
C56 VDD2.n40 B 0.012747f
C57 VDD2.n41 B 0.028456f
C58 VDD2.n42 B 0.028456f
C59 VDD2.n43 B 0.012747f
C60 VDD2.n44 B 0.012039f
C61 VDD2.n45 B 0.022404f
C62 VDD2.n46 B 0.022404f
C63 VDD2.n47 B 0.012039f
C64 VDD2.n48 B 0.012747f
C65 VDD2.n49 B 0.028456f
C66 VDD2.n50 B 0.028456f
C67 VDD2.n51 B 0.012747f
C68 VDD2.n52 B 0.012039f
C69 VDD2.n53 B 0.022404f
C70 VDD2.n54 B 0.022404f
C71 VDD2.n55 B 0.012039f
C72 VDD2.n56 B 0.012747f
C73 VDD2.n57 B 0.028456f
C74 VDD2.n58 B 0.028456f
C75 VDD2.n59 B 0.012747f
C76 VDD2.n60 B 0.012039f
C77 VDD2.n61 B 0.022404f
C78 VDD2.n62 B 0.022404f
C79 VDD2.n63 B 0.012039f
C80 VDD2.n64 B 0.012747f
C81 VDD2.n65 B 0.028456f
C82 VDD2.n66 B 0.028456f
C83 VDD2.n67 B 0.028456f
C84 VDD2.n68 B 0.012747f
C85 VDD2.n69 B 0.012039f
C86 VDD2.n70 B 0.022404f
C87 VDD2.n71 B 0.022404f
C88 VDD2.n72 B 0.012039f
C89 VDD2.n73 B 0.012393f
C90 VDD2.n74 B 0.012393f
C91 VDD2.n75 B 0.028456f
C92 VDD2.n76 B 0.055989f
C93 VDD2.n77 B 0.012747f
C94 VDD2.n78 B 0.012039f
C95 VDD2.n79 B 0.05148f
C96 VDD2.n80 B 0.051322f
C97 VDD2.t5 B 0.259017f
C98 VDD2.t8 B 0.259017f
C99 VDD2.n81 B 2.33828f
C100 VDD2.n82 B 0.480528f
C101 VDD2.t9 B 0.259017f
C102 VDD2.t6 B 0.259017f
C103 VDD2.n83 B 2.34559f
C104 VDD2.n84 B 2.24943f
C105 VDD2.n85 B 0.028317f
C106 VDD2.n86 B 0.022404f
C107 VDD2.n87 B 0.012039f
C108 VDD2.n88 B 0.028456f
C109 VDD2.n89 B 0.012747f
C110 VDD2.n90 B 0.022404f
C111 VDD2.n91 B 0.012039f
C112 VDD2.n92 B 0.028456f
C113 VDD2.n93 B 0.028456f
C114 VDD2.n94 B 0.012747f
C115 VDD2.n95 B 0.022404f
C116 VDD2.n96 B 0.012039f
C117 VDD2.n97 B 0.028456f
C118 VDD2.n98 B 0.012747f
C119 VDD2.n99 B 0.022404f
C120 VDD2.n100 B 0.012039f
C121 VDD2.n101 B 0.028456f
C122 VDD2.n102 B 0.012747f
C123 VDD2.n103 B 0.022404f
C124 VDD2.n104 B 0.012039f
C125 VDD2.n105 B 0.028456f
C126 VDD2.n106 B 0.012747f
C127 VDD2.n107 B 0.022404f
C128 VDD2.n108 B 0.012039f
C129 VDD2.n109 B 0.028456f
C130 VDD2.n110 B 0.012747f
C131 VDD2.n111 B 0.144047f
C132 VDD2.t3 B 0.046892f
C133 VDD2.n112 B 0.021342f
C134 VDD2.n113 B 0.01681f
C135 VDD2.n114 B 0.012039f
C136 VDD2.n115 B 1.41966f
C137 VDD2.n116 B 0.022404f
C138 VDD2.n117 B 0.012039f
C139 VDD2.n118 B 0.012747f
C140 VDD2.n119 B 0.028456f
C141 VDD2.n120 B 0.028456f
C142 VDD2.n121 B 0.012747f
C143 VDD2.n122 B 0.012039f
C144 VDD2.n123 B 0.022404f
C145 VDD2.n124 B 0.022404f
C146 VDD2.n125 B 0.012039f
C147 VDD2.n126 B 0.012747f
C148 VDD2.n127 B 0.028456f
C149 VDD2.n128 B 0.028456f
C150 VDD2.n129 B 0.012747f
C151 VDD2.n130 B 0.012039f
C152 VDD2.n131 B 0.022404f
C153 VDD2.n132 B 0.022404f
C154 VDD2.n133 B 0.012039f
C155 VDD2.n134 B 0.012747f
C156 VDD2.n135 B 0.028456f
C157 VDD2.n136 B 0.028456f
C158 VDD2.n137 B 0.012747f
C159 VDD2.n138 B 0.012039f
C160 VDD2.n139 B 0.022404f
C161 VDD2.n140 B 0.022404f
C162 VDD2.n141 B 0.012039f
C163 VDD2.n142 B 0.012747f
C164 VDD2.n143 B 0.028456f
C165 VDD2.n144 B 0.028456f
C166 VDD2.n145 B 0.012747f
C167 VDD2.n146 B 0.012039f
C168 VDD2.n147 B 0.022404f
C169 VDD2.n148 B 0.022404f
C170 VDD2.n149 B 0.012039f
C171 VDD2.n150 B 0.012747f
C172 VDD2.n151 B 0.028456f
C173 VDD2.n152 B 0.028456f
C174 VDD2.n153 B 0.012747f
C175 VDD2.n154 B 0.012039f
C176 VDD2.n155 B 0.022404f
C177 VDD2.n156 B 0.022404f
C178 VDD2.n157 B 0.012039f
C179 VDD2.n158 B 0.012393f
C180 VDD2.n159 B 0.012393f
C181 VDD2.n160 B 0.028456f
C182 VDD2.n161 B 0.055989f
C183 VDD2.n162 B 0.012747f
C184 VDD2.n163 B 0.012039f
C185 VDD2.n164 B 0.05148f
C186 VDD2.n165 B 0.046214f
C187 VDD2.n166 B 2.40306f
C188 VDD2.t7 B 0.259017f
C189 VDD2.t1 B 0.259017f
C190 VDD2.n167 B 2.33829f
C191 VDD2.n168 B 0.332987f
C192 VDD2.t0 B 0.259017f
C193 VDD2.t2 B 0.259017f
C194 VDD2.n169 B 2.34556f
C195 VN.n0 B 0.029142f
C196 VN.t3 B 1.79807f
C197 VN.n1 B 0.04701f
C198 VN.n2 B 0.029142f
C199 VN.t0 B 1.79807f
C200 VN.n3 B 0.055336f
C201 VN.n4 B 0.029142f
C202 VN.t1 B 1.79807f
C203 VN.n5 B 0.051912f
C204 VN.t5 B 1.89747f
C205 VN.t4 B 1.79807f
C206 VN.n6 B 0.701903f
C207 VN.n7 B 0.706397f
C208 VN.n8 B 0.186044f
C209 VN.n9 B 0.029142f
C210 VN.n10 B 0.02518f
C211 VN.n11 B 0.055336f
C212 VN.n12 B 0.667645f
C213 VN.n13 B 0.029142f
C214 VN.n14 B 0.029142f
C215 VN.n15 B 0.029142f
C216 VN.n16 B 0.02518f
C217 VN.n17 B 0.051912f
C218 VN.n18 B 0.640146f
C219 VN.n19 B 0.03447f
C220 VN.n20 B 0.029142f
C221 VN.n21 B 0.029142f
C222 VN.n22 B 0.029142f
C223 VN.n23 B 0.038078f
C224 VN.n24 B 0.040369f
C225 VN.n25 B 0.704406f
C226 VN.n26 B 0.027652f
C227 VN.n27 B 0.029142f
C228 VN.t6 B 1.79807f
C229 VN.n28 B 0.04701f
C230 VN.n29 B 0.029142f
C231 VN.t2 B 1.79807f
C232 VN.n30 B 0.055336f
C233 VN.n31 B 0.029142f
C234 VN.t8 B 1.79807f
C235 VN.n32 B 0.051912f
C236 VN.t7 B 1.89747f
C237 VN.t9 B 1.79807f
C238 VN.n33 B 0.701903f
C239 VN.n34 B 0.706397f
C240 VN.n35 B 0.186044f
C241 VN.n36 B 0.029142f
C242 VN.n37 B 0.02518f
C243 VN.n38 B 0.055336f
C244 VN.n39 B 0.667645f
C245 VN.n40 B 0.029142f
C246 VN.n41 B 0.029142f
C247 VN.n42 B 0.029142f
C248 VN.n43 B 0.02518f
C249 VN.n44 B 0.051912f
C250 VN.n45 B 0.640146f
C251 VN.n46 B 0.03447f
C252 VN.n47 B 0.029142f
C253 VN.n48 B 0.029142f
C254 VN.n49 B 0.029142f
C255 VN.n50 B 0.038078f
C256 VN.n51 B 0.040369f
C257 VN.n52 B 0.704406f
C258 VN.n53 B 1.57535f
C259 VTAIL.t7 B 0.27728f
C260 VTAIL.t4 B 0.27728f
C261 VTAIL.n0 B 2.43056f
C262 VTAIL.n1 B 0.432765f
C263 VTAIL.n2 B 0.030313f
C264 VTAIL.n3 B 0.023984f
C265 VTAIL.n4 B 0.012888f
C266 VTAIL.n5 B 0.030462f
C267 VTAIL.n6 B 0.013646f
C268 VTAIL.n7 B 0.023984f
C269 VTAIL.n8 B 0.012888f
C270 VTAIL.n9 B 0.030462f
C271 VTAIL.n10 B 0.013646f
C272 VTAIL.n11 B 0.023984f
C273 VTAIL.n12 B 0.012888f
C274 VTAIL.n13 B 0.030462f
C275 VTAIL.n14 B 0.013646f
C276 VTAIL.n15 B 0.023984f
C277 VTAIL.n16 B 0.012888f
C278 VTAIL.n17 B 0.030462f
C279 VTAIL.n18 B 0.013646f
C280 VTAIL.n19 B 0.023984f
C281 VTAIL.n20 B 0.012888f
C282 VTAIL.n21 B 0.030462f
C283 VTAIL.n22 B 0.013646f
C284 VTAIL.n23 B 0.023984f
C285 VTAIL.n24 B 0.012888f
C286 VTAIL.n25 B 0.030462f
C287 VTAIL.n26 B 0.013646f
C288 VTAIL.n27 B 0.154204f
C289 VTAIL.t10 B 0.050198f
C290 VTAIL.n28 B 0.022847f
C291 VTAIL.n29 B 0.017995f
C292 VTAIL.n30 B 0.012888f
C293 VTAIL.n31 B 1.51976f
C294 VTAIL.n32 B 0.023984f
C295 VTAIL.n33 B 0.012888f
C296 VTAIL.n34 B 0.013646f
C297 VTAIL.n35 B 0.030462f
C298 VTAIL.n36 B 0.030462f
C299 VTAIL.n37 B 0.013646f
C300 VTAIL.n38 B 0.012888f
C301 VTAIL.n39 B 0.023984f
C302 VTAIL.n40 B 0.023984f
C303 VTAIL.n41 B 0.012888f
C304 VTAIL.n42 B 0.013646f
C305 VTAIL.n43 B 0.030462f
C306 VTAIL.n44 B 0.030462f
C307 VTAIL.n45 B 0.013646f
C308 VTAIL.n46 B 0.012888f
C309 VTAIL.n47 B 0.023984f
C310 VTAIL.n48 B 0.023984f
C311 VTAIL.n49 B 0.012888f
C312 VTAIL.n50 B 0.013646f
C313 VTAIL.n51 B 0.030462f
C314 VTAIL.n52 B 0.030462f
C315 VTAIL.n53 B 0.013646f
C316 VTAIL.n54 B 0.012888f
C317 VTAIL.n55 B 0.023984f
C318 VTAIL.n56 B 0.023984f
C319 VTAIL.n57 B 0.012888f
C320 VTAIL.n58 B 0.013646f
C321 VTAIL.n59 B 0.030462f
C322 VTAIL.n60 B 0.030462f
C323 VTAIL.n61 B 0.013646f
C324 VTAIL.n62 B 0.012888f
C325 VTAIL.n63 B 0.023984f
C326 VTAIL.n64 B 0.023984f
C327 VTAIL.n65 B 0.012888f
C328 VTAIL.n66 B 0.013646f
C329 VTAIL.n67 B 0.030462f
C330 VTAIL.n68 B 0.030462f
C331 VTAIL.n69 B 0.030462f
C332 VTAIL.n70 B 0.013646f
C333 VTAIL.n71 B 0.012888f
C334 VTAIL.n72 B 0.023984f
C335 VTAIL.n73 B 0.023984f
C336 VTAIL.n74 B 0.012888f
C337 VTAIL.n75 B 0.013267f
C338 VTAIL.n76 B 0.013267f
C339 VTAIL.n77 B 0.030462f
C340 VTAIL.n78 B 0.059937f
C341 VTAIL.n79 B 0.013646f
C342 VTAIL.n80 B 0.012888f
C343 VTAIL.n81 B 0.05511f
C344 VTAIL.n82 B 0.032909f
C345 VTAIL.n83 B 0.243483f
C346 VTAIL.t13 B 0.27728f
C347 VTAIL.t19 B 0.27728f
C348 VTAIL.n84 B 2.43056f
C349 VTAIL.n85 B 0.485397f
C350 VTAIL.t12 B 0.27728f
C351 VTAIL.t14 B 0.27728f
C352 VTAIL.n86 B 2.43056f
C353 VTAIL.n87 B 1.91046f
C354 VTAIL.t9 B 0.27728f
C355 VTAIL.t2 B 0.27728f
C356 VTAIL.n88 B 2.43058f
C357 VTAIL.n89 B 1.91044f
C358 VTAIL.t5 B 0.27728f
C359 VTAIL.t1 B 0.27728f
C360 VTAIL.n90 B 2.43058f
C361 VTAIL.n91 B 0.485384f
C362 VTAIL.n92 B 0.030313f
C363 VTAIL.n93 B 0.023984f
C364 VTAIL.n94 B 0.012888f
C365 VTAIL.n95 B 0.030462f
C366 VTAIL.n96 B 0.013646f
C367 VTAIL.n97 B 0.023984f
C368 VTAIL.n98 B 0.012888f
C369 VTAIL.n99 B 0.030462f
C370 VTAIL.n100 B 0.030462f
C371 VTAIL.n101 B 0.013646f
C372 VTAIL.n102 B 0.023984f
C373 VTAIL.n103 B 0.012888f
C374 VTAIL.n104 B 0.030462f
C375 VTAIL.n105 B 0.013646f
C376 VTAIL.n106 B 0.023984f
C377 VTAIL.n107 B 0.012888f
C378 VTAIL.n108 B 0.030462f
C379 VTAIL.n109 B 0.013646f
C380 VTAIL.n110 B 0.023984f
C381 VTAIL.n111 B 0.012888f
C382 VTAIL.n112 B 0.030462f
C383 VTAIL.n113 B 0.013646f
C384 VTAIL.n114 B 0.023984f
C385 VTAIL.n115 B 0.012888f
C386 VTAIL.n116 B 0.030462f
C387 VTAIL.n117 B 0.013646f
C388 VTAIL.n118 B 0.154204f
C389 VTAIL.t6 B 0.050198f
C390 VTAIL.n119 B 0.022847f
C391 VTAIL.n120 B 0.017995f
C392 VTAIL.n121 B 0.012888f
C393 VTAIL.n122 B 1.51976f
C394 VTAIL.n123 B 0.023984f
C395 VTAIL.n124 B 0.012888f
C396 VTAIL.n125 B 0.013646f
C397 VTAIL.n126 B 0.030462f
C398 VTAIL.n127 B 0.030462f
C399 VTAIL.n128 B 0.013646f
C400 VTAIL.n129 B 0.012888f
C401 VTAIL.n130 B 0.023984f
C402 VTAIL.n131 B 0.023984f
C403 VTAIL.n132 B 0.012888f
C404 VTAIL.n133 B 0.013646f
C405 VTAIL.n134 B 0.030462f
C406 VTAIL.n135 B 0.030462f
C407 VTAIL.n136 B 0.013646f
C408 VTAIL.n137 B 0.012888f
C409 VTAIL.n138 B 0.023984f
C410 VTAIL.n139 B 0.023984f
C411 VTAIL.n140 B 0.012888f
C412 VTAIL.n141 B 0.013646f
C413 VTAIL.n142 B 0.030462f
C414 VTAIL.n143 B 0.030462f
C415 VTAIL.n144 B 0.013646f
C416 VTAIL.n145 B 0.012888f
C417 VTAIL.n146 B 0.023984f
C418 VTAIL.n147 B 0.023984f
C419 VTAIL.n148 B 0.012888f
C420 VTAIL.n149 B 0.013646f
C421 VTAIL.n150 B 0.030462f
C422 VTAIL.n151 B 0.030462f
C423 VTAIL.n152 B 0.013646f
C424 VTAIL.n153 B 0.012888f
C425 VTAIL.n154 B 0.023984f
C426 VTAIL.n155 B 0.023984f
C427 VTAIL.n156 B 0.012888f
C428 VTAIL.n157 B 0.013646f
C429 VTAIL.n158 B 0.030462f
C430 VTAIL.n159 B 0.030462f
C431 VTAIL.n160 B 0.013646f
C432 VTAIL.n161 B 0.012888f
C433 VTAIL.n162 B 0.023984f
C434 VTAIL.n163 B 0.023984f
C435 VTAIL.n164 B 0.012888f
C436 VTAIL.n165 B 0.013267f
C437 VTAIL.n166 B 0.013267f
C438 VTAIL.n167 B 0.030462f
C439 VTAIL.n168 B 0.059937f
C440 VTAIL.n169 B 0.013646f
C441 VTAIL.n170 B 0.012888f
C442 VTAIL.n171 B 0.05511f
C443 VTAIL.n172 B 0.032909f
C444 VTAIL.n173 B 0.243483f
C445 VTAIL.t18 B 0.27728f
C446 VTAIL.t16 B 0.27728f
C447 VTAIL.n174 B 2.43058f
C448 VTAIL.n175 B 0.459401f
C449 VTAIL.t17 B 0.27728f
C450 VTAIL.t15 B 0.27728f
C451 VTAIL.n176 B 2.43058f
C452 VTAIL.n177 B 0.485384f
C453 VTAIL.n178 B 0.030313f
C454 VTAIL.n179 B 0.023984f
C455 VTAIL.n180 B 0.012888f
C456 VTAIL.n181 B 0.030462f
C457 VTAIL.n182 B 0.013646f
C458 VTAIL.n183 B 0.023984f
C459 VTAIL.n184 B 0.012888f
C460 VTAIL.n185 B 0.030462f
C461 VTAIL.n186 B 0.030462f
C462 VTAIL.n187 B 0.013646f
C463 VTAIL.n188 B 0.023984f
C464 VTAIL.n189 B 0.012888f
C465 VTAIL.n190 B 0.030462f
C466 VTAIL.n191 B 0.013646f
C467 VTAIL.n192 B 0.023984f
C468 VTAIL.n193 B 0.012888f
C469 VTAIL.n194 B 0.030462f
C470 VTAIL.n195 B 0.013646f
C471 VTAIL.n196 B 0.023984f
C472 VTAIL.n197 B 0.012888f
C473 VTAIL.n198 B 0.030462f
C474 VTAIL.n199 B 0.013646f
C475 VTAIL.n200 B 0.023984f
C476 VTAIL.n201 B 0.012888f
C477 VTAIL.n202 B 0.030462f
C478 VTAIL.n203 B 0.013646f
C479 VTAIL.n204 B 0.154204f
C480 VTAIL.t11 B 0.050198f
C481 VTAIL.n205 B 0.022847f
C482 VTAIL.n206 B 0.017995f
C483 VTAIL.n207 B 0.012888f
C484 VTAIL.n208 B 1.51976f
C485 VTAIL.n209 B 0.023984f
C486 VTAIL.n210 B 0.012888f
C487 VTAIL.n211 B 0.013646f
C488 VTAIL.n212 B 0.030462f
C489 VTAIL.n213 B 0.030462f
C490 VTAIL.n214 B 0.013646f
C491 VTAIL.n215 B 0.012888f
C492 VTAIL.n216 B 0.023984f
C493 VTAIL.n217 B 0.023984f
C494 VTAIL.n218 B 0.012888f
C495 VTAIL.n219 B 0.013646f
C496 VTAIL.n220 B 0.030462f
C497 VTAIL.n221 B 0.030462f
C498 VTAIL.n222 B 0.013646f
C499 VTAIL.n223 B 0.012888f
C500 VTAIL.n224 B 0.023984f
C501 VTAIL.n225 B 0.023984f
C502 VTAIL.n226 B 0.012888f
C503 VTAIL.n227 B 0.013646f
C504 VTAIL.n228 B 0.030462f
C505 VTAIL.n229 B 0.030462f
C506 VTAIL.n230 B 0.013646f
C507 VTAIL.n231 B 0.012888f
C508 VTAIL.n232 B 0.023984f
C509 VTAIL.n233 B 0.023984f
C510 VTAIL.n234 B 0.012888f
C511 VTAIL.n235 B 0.013646f
C512 VTAIL.n236 B 0.030462f
C513 VTAIL.n237 B 0.030462f
C514 VTAIL.n238 B 0.013646f
C515 VTAIL.n239 B 0.012888f
C516 VTAIL.n240 B 0.023984f
C517 VTAIL.n241 B 0.023984f
C518 VTAIL.n242 B 0.012888f
C519 VTAIL.n243 B 0.013646f
C520 VTAIL.n244 B 0.030462f
C521 VTAIL.n245 B 0.030462f
C522 VTAIL.n246 B 0.013646f
C523 VTAIL.n247 B 0.012888f
C524 VTAIL.n248 B 0.023984f
C525 VTAIL.n249 B 0.023984f
C526 VTAIL.n250 B 0.012888f
C527 VTAIL.n251 B 0.013267f
C528 VTAIL.n252 B 0.013267f
C529 VTAIL.n253 B 0.030462f
C530 VTAIL.n254 B 0.059937f
C531 VTAIL.n255 B 0.013646f
C532 VTAIL.n256 B 0.012888f
C533 VTAIL.n257 B 0.05511f
C534 VTAIL.n258 B 0.032909f
C535 VTAIL.n259 B 1.56994f
C536 VTAIL.n260 B 0.030313f
C537 VTAIL.n261 B 0.023984f
C538 VTAIL.n262 B 0.012888f
C539 VTAIL.n263 B 0.030462f
C540 VTAIL.n264 B 0.013646f
C541 VTAIL.n265 B 0.023984f
C542 VTAIL.n266 B 0.012888f
C543 VTAIL.n267 B 0.030462f
C544 VTAIL.n268 B 0.013646f
C545 VTAIL.n269 B 0.023984f
C546 VTAIL.n270 B 0.012888f
C547 VTAIL.n271 B 0.030462f
C548 VTAIL.n272 B 0.013646f
C549 VTAIL.n273 B 0.023984f
C550 VTAIL.n274 B 0.012888f
C551 VTAIL.n275 B 0.030462f
C552 VTAIL.n276 B 0.013646f
C553 VTAIL.n277 B 0.023984f
C554 VTAIL.n278 B 0.012888f
C555 VTAIL.n279 B 0.030462f
C556 VTAIL.n280 B 0.013646f
C557 VTAIL.n281 B 0.023984f
C558 VTAIL.n282 B 0.012888f
C559 VTAIL.n283 B 0.030462f
C560 VTAIL.n284 B 0.013646f
C561 VTAIL.n285 B 0.154204f
C562 VTAIL.t0 B 0.050198f
C563 VTAIL.n286 B 0.022847f
C564 VTAIL.n287 B 0.017995f
C565 VTAIL.n288 B 0.012888f
C566 VTAIL.n289 B 1.51976f
C567 VTAIL.n290 B 0.023984f
C568 VTAIL.n291 B 0.012888f
C569 VTAIL.n292 B 0.013646f
C570 VTAIL.n293 B 0.030462f
C571 VTAIL.n294 B 0.030462f
C572 VTAIL.n295 B 0.013646f
C573 VTAIL.n296 B 0.012888f
C574 VTAIL.n297 B 0.023984f
C575 VTAIL.n298 B 0.023984f
C576 VTAIL.n299 B 0.012888f
C577 VTAIL.n300 B 0.013646f
C578 VTAIL.n301 B 0.030462f
C579 VTAIL.n302 B 0.030462f
C580 VTAIL.n303 B 0.013646f
C581 VTAIL.n304 B 0.012888f
C582 VTAIL.n305 B 0.023984f
C583 VTAIL.n306 B 0.023984f
C584 VTAIL.n307 B 0.012888f
C585 VTAIL.n308 B 0.013646f
C586 VTAIL.n309 B 0.030462f
C587 VTAIL.n310 B 0.030462f
C588 VTAIL.n311 B 0.013646f
C589 VTAIL.n312 B 0.012888f
C590 VTAIL.n313 B 0.023984f
C591 VTAIL.n314 B 0.023984f
C592 VTAIL.n315 B 0.012888f
C593 VTAIL.n316 B 0.013646f
C594 VTAIL.n317 B 0.030462f
C595 VTAIL.n318 B 0.030462f
C596 VTAIL.n319 B 0.013646f
C597 VTAIL.n320 B 0.012888f
C598 VTAIL.n321 B 0.023984f
C599 VTAIL.n322 B 0.023984f
C600 VTAIL.n323 B 0.012888f
C601 VTAIL.n324 B 0.013646f
C602 VTAIL.n325 B 0.030462f
C603 VTAIL.n326 B 0.030462f
C604 VTAIL.n327 B 0.030462f
C605 VTAIL.n328 B 0.013646f
C606 VTAIL.n329 B 0.012888f
C607 VTAIL.n330 B 0.023984f
C608 VTAIL.n331 B 0.023984f
C609 VTAIL.n332 B 0.012888f
C610 VTAIL.n333 B 0.013267f
C611 VTAIL.n334 B 0.013267f
C612 VTAIL.n335 B 0.030462f
C613 VTAIL.n336 B 0.059937f
C614 VTAIL.n337 B 0.013646f
C615 VTAIL.n338 B 0.012888f
C616 VTAIL.n339 B 0.05511f
C617 VTAIL.n340 B 0.032909f
C618 VTAIL.n341 B 1.56994f
C619 VTAIL.t8 B 0.27728f
C620 VTAIL.t3 B 0.27728f
C621 VTAIL.n342 B 2.43056f
C622 VTAIL.n343 B 0.387462f
C623 VDD1.n0 B 0.028574f
C624 VDD1.n1 B 0.022608f
C625 VDD1.n2 B 0.012149f
C626 VDD1.n3 B 0.028715f
C627 VDD1.n4 B 0.012863f
C628 VDD1.n5 B 0.022608f
C629 VDD1.n6 B 0.012149f
C630 VDD1.n7 B 0.028715f
C631 VDD1.n8 B 0.028715f
C632 VDD1.n9 B 0.012863f
C633 VDD1.n10 B 0.022608f
C634 VDD1.n11 B 0.012149f
C635 VDD1.n12 B 0.028715f
C636 VDD1.n13 B 0.012863f
C637 VDD1.n14 B 0.022608f
C638 VDD1.n15 B 0.012149f
C639 VDD1.n16 B 0.028715f
C640 VDD1.n17 B 0.012863f
C641 VDD1.n18 B 0.022608f
C642 VDD1.n19 B 0.012149f
C643 VDD1.n20 B 0.028715f
C644 VDD1.n21 B 0.012863f
C645 VDD1.n22 B 0.022608f
C646 VDD1.n23 B 0.012149f
C647 VDD1.n24 B 0.028715f
C648 VDD1.n25 B 0.012863f
C649 VDD1.n26 B 0.145357f
C650 VDD1.t6 B 0.047319f
C651 VDD1.n27 B 0.021536f
C652 VDD1.n28 B 0.016963f
C653 VDD1.n29 B 0.012149f
C654 VDD1.n30 B 1.43258f
C655 VDD1.n31 B 0.022608f
C656 VDD1.n32 B 0.012149f
C657 VDD1.n33 B 0.012863f
C658 VDD1.n34 B 0.028715f
C659 VDD1.n35 B 0.028715f
C660 VDD1.n36 B 0.012863f
C661 VDD1.n37 B 0.012149f
C662 VDD1.n38 B 0.022608f
C663 VDD1.n39 B 0.022608f
C664 VDD1.n40 B 0.012149f
C665 VDD1.n41 B 0.012863f
C666 VDD1.n42 B 0.028715f
C667 VDD1.n43 B 0.028715f
C668 VDD1.n44 B 0.012863f
C669 VDD1.n45 B 0.012149f
C670 VDD1.n46 B 0.022608f
C671 VDD1.n47 B 0.022608f
C672 VDD1.n48 B 0.012149f
C673 VDD1.n49 B 0.012863f
C674 VDD1.n50 B 0.028715f
C675 VDD1.n51 B 0.028715f
C676 VDD1.n52 B 0.012863f
C677 VDD1.n53 B 0.012149f
C678 VDD1.n54 B 0.022608f
C679 VDD1.n55 B 0.022608f
C680 VDD1.n56 B 0.012149f
C681 VDD1.n57 B 0.012863f
C682 VDD1.n58 B 0.028715f
C683 VDD1.n59 B 0.028715f
C684 VDD1.n60 B 0.012863f
C685 VDD1.n61 B 0.012149f
C686 VDD1.n62 B 0.022608f
C687 VDD1.n63 B 0.022608f
C688 VDD1.n64 B 0.012149f
C689 VDD1.n65 B 0.012863f
C690 VDD1.n66 B 0.028715f
C691 VDD1.n67 B 0.028715f
C692 VDD1.n68 B 0.012863f
C693 VDD1.n69 B 0.012149f
C694 VDD1.n70 B 0.022608f
C695 VDD1.n71 B 0.022608f
C696 VDD1.n72 B 0.012149f
C697 VDD1.n73 B 0.012506f
C698 VDD1.n74 B 0.012506f
C699 VDD1.n75 B 0.028715f
C700 VDD1.n76 B 0.056498f
C701 VDD1.n77 B 0.012863f
C702 VDD1.n78 B 0.012149f
C703 VDD1.n79 B 0.051949f
C704 VDD1.n80 B 0.051789f
C705 VDD1.t2 B 0.261374f
C706 VDD1.t3 B 0.261374f
C707 VDD1.n81 B 2.35956f
C708 VDD1.n82 B 0.491654f
C709 VDD1.n83 B 0.028574f
C710 VDD1.n84 B 0.022608f
C711 VDD1.n85 B 0.012149f
C712 VDD1.n86 B 0.028715f
C713 VDD1.n87 B 0.012863f
C714 VDD1.n88 B 0.022608f
C715 VDD1.n89 B 0.012149f
C716 VDD1.n90 B 0.028715f
C717 VDD1.n91 B 0.012863f
C718 VDD1.n92 B 0.022608f
C719 VDD1.n93 B 0.012149f
C720 VDD1.n94 B 0.028715f
C721 VDD1.n95 B 0.012863f
C722 VDD1.n96 B 0.022608f
C723 VDD1.n97 B 0.012149f
C724 VDD1.n98 B 0.028715f
C725 VDD1.n99 B 0.012863f
C726 VDD1.n100 B 0.022608f
C727 VDD1.n101 B 0.012149f
C728 VDD1.n102 B 0.028715f
C729 VDD1.n103 B 0.012863f
C730 VDD1.n104 B 0.022608f
C731 VDD1.n105 B 0.012149f
C732 VDD1.n106 B 0.028715f
C733 VDD1.n107 B 0.012863f
C734 VDD1.n108 B 0.145357f
C735 VDD1.t4 B 0.047319f
C736 VDD1.n109 B 0.021536f
C737 VDD1.n110 B 0.016963f
C738 VDD1.n111 B 0.012149f
C739 VDD1.n112 B 1.43258f
C740 VDD1.n113 B 0.022608f
C741 VDD1.n114 B 0.012149f
C742 VDD1.n115 B 0.012863f
C743 VDD1.n116 B 0.028715f
C744 VDD1.n117 B 0.028715f
C745 VDD1.n118 B 0.012863f
C746 VDD1.n119 B 0.012149f
C747 VDD1.n120 B 0.022608f
C748 VDD1.n121 B 0.022608f
C749 VDD1.n122 B 0.012149f
C750 VDD1.n123 B 0.012863f
C751 VDD1.n124 B 0.028715f
C752 VDD1.n125 B 0.028715f
C753 VDD1.n126 B 0.012863f
C754 VDD1.n127 B 0.012149f
C755 VDD1.n128 B 0.022608f
C756 VDD1.n129 B 0.022608f
C757 VDD1.n130 B 0.012149f
C758 VDD1.n131 B 0.012863f
C759 VDD1.n132 B 0.028715f
C760 VDD1.n133 B 0.028715f
C761 VDD1.n134 B 0.012863f
C762 VDD1.n135 B 0.012149f
C763 VDD1.n136 B 0.022608f
C764 VDD1.n137 B 0.022608f
C765 VDD1.n138 B 0.012149f
C766 VDD1.n139 B 0.012863f
C767 VDD1.n140 B 0.028715f
C768 VDD1.n141 B 0.028715f
C769 VDD1.n142 B 0.012863f
C770 VDD1.n143 B 0.012149f
C771 VDD1.n144 B 0.022608f
C772 VDD1.n145 B 0.022608f
C773 VDD1.n146 B 0.012149f
C774 VDD1.n147 B 0.012863f
C775 VDD1.n148 B 0.028715f
C776 VDD1.n149 B 0.028715f
C777 VDD1.n150 B 0.028715f
C778 VDD1.n151 B 0.012863f
C779 VDD1.n152 B 0.012149f
C780 VDD1.n153 B 0.022608f
C781 VDD1.n154 B 0.022608f
C782 VDD1.n155 B 0.012149f
C783 VDD1.n156 B 0.012506f
C784 VDD1.n157 B 0.012506f
C785 VDD1.n158 B 0.028715f
C786 VDD1.n159 B 0.056498f
C787 VDD1.n160 B 0.012863f
C788 VDD1.n161 B 0.012149f
C789 VDD1.n162 B 0.051949f
C790 VDD1.n163 B 0.051789f
C791 VDD1.t8 B 0.261374f
C792 VDD1.t5 B 0.261374f
C793 VDD1.n164 B 2.35955f
C794 VDD1.n165 B 0.484899f
C795 VDD1.t7 B 0.261374f
C796 VDD1.t0 B 0.261374f
C797 VDD1.n166 B 2.36693f
C798 VDD1.n167 B 2.35915f
C799 VDD1.t9 B 0.261374f
C800 VDD1.t1 B 0.261374f
C801 VDD1.n168 B 2.35955f
C802 VDD1.n169 B 2.65374f
C803 VP.n0 B 0.029473f
C804 VP.t9 B 1.81854f
C805 VP.n1 B 0.047545f
C806 VP.n2 B 0.029473f
C807 VP.t0 B 1.81854f
C808 VP.n3 B 0.055966f
C809 VP.n4 B 0.029473f
C810 VP.t6 B 1.81854f
C811 VP.n5 B 0.052503f
C812 VP.n6 B 0.029473f
C813 VP.n7 B 0.040828f
C814 VP.n8 B 0.029473f
C815 VP.t8 B 1.81854f
C816 VP.n9 B 0.047545f
C817 VP.n10 B 0.029473f
C818 VP.t4 B 1.81854f
C819 VP.n11 B 0.055966f
C820 VP.n12 B 0.029473f
C821 VP.t2 B 1.81854f
C822 VP.n13 B 0.052503f
C823 VP.t1 B 1.91906f
C824 VP.t3 B 1.81854f
C825 VP.n14 B 0.709892f
C826 VP.n15 B 0.714437f
C827 VP.n16 B 0.188162f
C828 VP.n17 B 0.029473f
C829 VP.n18 B 0.025467f
C830 VP.n19 B 0.055966f
C831 VP.n20 B 0.675243f
C832 VP.n21 B 0.029473f
C833 VP.n22 B 0.029473f
C834 VP.n23 B 0.029473f
C835 VP.n24 B 0.025467f
C836 VP.n25 B 0.052503f
C837 VP.n26 B 0.647432f
C838 VP.n27 B 0.034862f
C839 VP.n28 B 0.029473f
C840 VP.n29 B 0.029473f
C841 VP.n30 B 0.029473f
C842 VP.n31 B 0.038511f
C843 VP.n32 B 0.040828f
C844 VP.n33 B 0.712423f
C845 VP.n34 B 1.57411f
C846 VP.t7 B 1.81854f
C847 VP.n35 B 0.712423f
C848 VP.n36 B 1.59559f
C849 VP.n37 B 0.029473f
C850 VP.n38 B 0.029473f
C851 VP.n39 B 0.038511f
C852 VP.n40 B 0.047545f
C853 VP.t5 B 1.81854f
C854 VP.n41 B 0.647432f
C855 VP.n42 B 0.034862f
C856 VP.n43 B 0.029473f
C857 VP.n44 B 0.029473f
C858 VP.n45 B 0.029473f
C859 VP.n46 B 0.025467f
C860 VP.n47 B 0.055966f
C861 VP.n48 B 0.675243f
C862 VP.n49 B 0.029473f
C863 VP.n50 B 0.029473f
C864 VP.n51 B 0.029473f
C865 VP.n52 B 0.025467f
C866 VP.n53 B 0.052503f
C867 VP.n54 B 0.647432f
C868 VP.n55 B 0.034862f
C869 VP.n56 B 0.029473f
C870 VP.n57 B 0.029473f
C871 VP.n58 B 0.029473f
C872 VP.n59 B 0.038511f
C873 VP.n60 B 0.040828f
C874 VP.n61 B 0.712423f
C875 VP.n62 B 0.027967f
.ends

