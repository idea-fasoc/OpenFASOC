* NGSPICE file created from diff_pair_sample_0723.ext - technology: sky130A

.subckt diff_pair_sample_0723 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t7 VP.t0 VDD1.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=6.5988 pd=34.62 as=2.7918 ps=17.25 w=16.92 l=1.06
X1 B.t17 B.t15 B.t16 B.t12 sky130_fd_pr__nfet_01v8 ad=6.5988 pd=34.62 as=0 ps=0 w=16.92 l=1.06
X2 VDD1.t0 VP.t1 VTAIL.t6 B.t0 sky130_fd_pr__nfet_01v8 ad=2.7918 pd=17.25 as=6.5988 ps=34.62 w=16.92 l=1.06
X3 B.t14 B.t11 B.t13 B.t12 sky130_fd_pr__nfet_01v8 ad=6.5988 pd=34.62 as=0 ps=0 w=16.92 l=1.06
X4 VDD2.t3 VN.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.7918 pd=17.25 as=6.5988 ps=34.62 w=16.92 l=1.06
X5 VDD1.t3 VP.t2 VTAIL.t5 B.t1 sky130_fd_pr__nfet_01v8 ad=2.7918 pd=17.25 as=6.5988 ps=34.62 w=16.92 l=1.06
X6 VTAIL.t2 VN.t1 VDD2.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=6.5988 pd=34.62 as=2.7918 ps=17.25 w=16.92 l=1.06
X7 VDD2.t1 VN.t2 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.7918 pd=17.25 as=6.5988 ps=34.62 w=16.92 l=1.06
X8 B.t10 B.t8 B.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=6.5988 pd=34.62 as=0 ps=0 w=16.92 l=1.06
X9 VTAIL.t3 VN.t3 VDD2.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=6.5988 pd=34.62 as=2.7918 ps=17.25 w=16.92 l=1.06
X10 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=6.5988 pd=34.62 as=0 ps=0 w=16.92 l=1.06
X11 VTAIL.t4 VP.t3 VDD1.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=6.5988 pd=34.62 as=2.7918 ps=17.25 w=16.92 l=1.06
R0 VP.n0 VP.t0 440.812
R1 VP.n0 VP.t2 440.724
R2 VP.n2 VP.t3 422.205
R3 VP.n3 VP.t1 422.205
R4 VP.n4 VP.n3 80.6037
R5 VP.n2 VP.n1 80.6037
R6 VP.n1 VP.n0 76.6168
R7 VP.n3 VP.n2 48.2005
R8 VP.n4 VP.n1 0.380177
R9 VP VP.n4 0.146778
R10 VDD1 VDD1.n1 105.472
R11 VDD1 VDD1.n0 63.1101
R12 VDD1.n0 VDD1.t1 1.17071
R13 VDD1.n0 VDD1.t3 1.17071
R14 VDD1.n1 VDD1.t2 1.17071
R15 VDD1.n1 VDD1.t0 1.17071
R16 VTAIL.n746 VTAIL.n658 289.615
R17 VTAIL.n88 VTAIL.n0 289.615
R18 VTAIL.n182 VTAIL.n94 289.615
R19 VTAIL.n276 VTAIL.n188 289.615
R20 VTAIL.n652 VTAIL.n564 289.615
R21 VTAIL.n558 VTAIL.n470 289.615
R22 VTAIL.n464 VTAIL.n376 289.615
R23 VTAIL.n370 VTAIL.n282 289.615
R24 VTAIL.n689 VTAIL.n688 185
R25 VTAIL.n686 VTAIL.n685 185
R26 VTAIL.n695 VTAIL.n694 185
R27 VTAIL.n697 VTAIL.n696 185
R28 VTAIL.n682 VTAIL.n681 185
R29 VTAIL.n703 VTAIL.n702 185
R30 VTAIL.n705 VTAIL.n704 185
R31 VTAIL.n678 VTAIL.n677 185
R32 VTAIL.n711 VTAIL.n710 185
R33 VTAIL.n713 VTAIL.n712 185
R34 VTAIL.n674 VTAIL.n673 185
R35 VTAIL.n719 VTAIL.n718 185
R36 VTAIL.n721 VTAIL.n720 185
R37 VTAIL.n670 VTAIL.n669 185
R38 VTAIL.n727 VTAIL.n726 185
R39 VTAIL.n730 VTAIL.n729 185
R40 VTAIL.n728 VTAIL.n666 185
R41 VTAIL.n735 VTAIL.n665 185
R42 VTAIL.n737 VTAIL.n736 185
R43 VTAIL.n739 VTAIL.n738 185
R44 VTAIL.n662 VTAIL.n661 185
R45 VTAIL.n745 VTAIL.n744 185
R46 VTAIL.n747 VTAIL.n746 185
R47 VTAIL.n31 VTAIL.n30 185
R48 VTAIL.n28 VTAIL.n27 185
R49 VTAIL.n37 VTAIL.n36 185
R50 VTAIL.n39 VTAIL.n38 185
R51 VTAIL.n24 VTAIL.n23 185
R52 VTAIL.n45 VTAIL.n44 185
R53 VTAIL.n47 VTAIL.n46 185
R54 VTAIL.n20 VTAIL.n19 185
R55 VTAIL.n53 VTAIL.n52 185
R56 VTAIL.n55 VTAIL.n54 185
R57 VTAIL.n16 VTAIL.n15 185
R58 VTAIL.n61 VTAIL.n60 185
R59 VTAIL.n63 VTAIL.n62 185
R60 VTAIL.n12 VTAIL.n11 185
R61 VTAIL.n69 VTAIL.n68 185
R62 VTAIL.n72 VTAIL.n71 185
R63 VTAIL.n70 VTAIL.n8 185
R64 VTAIL.n77 VTAIL.n7 185
R65 VTAIL.n79 VTAIL.n78 185
R66 VTAIL.n81 VTAIL.n80 185
R67 VTAIL.n4 VTAIL.n3 185
R68 VTAIL.n87 VTAIL.n86 185
R69 VTAIL.n89 VTAIL.n88 185
R70 VTAIL.n125 VTAIL.n124 185
R71 VTAIL.n122 VTAIL.n121 185
R72 VTAIL.n131 VTAIL.n130 185
R73 VTAIL.n133 VTAIL.n132 185
R74 VTAIL.n118 VTAIL.n117 185
R75 VTAIL.n139 VTAIL.n138 185
R76 VTAIL.n141 VTAIL.n140 185
R77 VTAIL.n114 VTAIL.n113 185
R78 VTAIL.n147 VTAIL.n146 185
R79 VTAIL.n149 VTAIL.n148 185
R80 VTAIL.n110 VTAIL.n109 185
R81 VTAIL.n155 VTAIL.n154 185
R82 VTAIL.n157 VTAIL.n156 185
R83 VTAIL.n106 VTAIL.n105 185
R84 VTAIL.n163 VTAIL.n162 185
R85 VTAIL.n166 VTAIL.n165 185
R86 VTAIL.n164 VTAIL.n102 185
R87 VTAIL.n171 VTAIL.n101 185
R88 VTAIL.n173 VTAIL.n172 185
R89 VTAIL.n175 VTAIL.n174 185
R90 VTAIL.n98 VTAIL.n97 185
R91 VTAIL.n181 VTAIL.n180 185
R92 VTAIL.n183 VTAIL.n182 185
R93 VTAIL.n219 VTAIL.n218 185
R94 VTAIL.n216 VTAIL.n215 185
R95 VTAIL.n225 VTAIL.n224 185
R96 VTAIL.n227 VTAIL.n226 185
R97 VTAIL.n212 VTAIL.n211 185
R98 VTAIL.n233 VTAIL.n232 185
R99 VTAIL.n235 VTAIL.n234 185
R100 VTAIL.n208 VTAIL.n207 185
R101 VTAIL.n241 VTAIL.n240 185
R102 VTAIL.n243 VTAIL.n242 185
R103 VTAIL.n204 VTAIL.n203 185
R104 VTAIL.n249 VTAIL.n248 185
R105 VTAIL.n251 VTAIL.n250 185
R106 VTAIL.n200 VTAIL.n199 185
R107 VTAIL.n257 VTAIL.n256 185
R108 VTAIL.n260 VTAIL.n259 185
R109 VTAIL.n258 VTAIL.n196 185
R110 VTAIL.n265 VTAIL.n195 185
R111 VTAIL.n267 VTAIL.n266 185
R112 VTAIL.n269 VTAIL.n268 185
R113 VTAIL.n192 VTAIL.n191 185
R114 VTAIL.n275 VTAIL.n274 185
R115 VTAIL.n277 VTAIL.n276 185
R116 VTAIL.n653 VTAIL.n652 185
R117 VTAIL.n651 VTAIL.n650 185
R118 VTAIL.n568 VTAIL.n567 185
R119 VTAIL.n645 VTAIL.n644 185
R120 VTAIL.n643 VTAIL.n642 185
R121 VTAIL.n641 VTAIL.n571 185
R122 VTAIL.n575 VTAIL.n572 185
R123 VTAIL.n636 VTAIL.n635 185
R124 VTAIL.n634 VTAIL.n633 185
R125 VTAIL.n577 VTAIL.n576 185
R126 VTAIL.n628 VTAIL.n627 185
R127 VTAIL.n626 VTAIL.n625 185
R128 VTAIL.n581 VTAIL.n580 185
R129 VTAIL.n620 VTAIL.n619 185
R130 VTAIL.n618 VTAIL.n617 185
R131 VTAIL.n585 VTAIL.n584 185
R132 VTAIL.n612 VTAIL.n611 185
R133 VTAIL.n610 VTAIL.n609 185
R134 VTAIL.n589 VTAIL.n588 185
R135 VTAIL.n604 VTAIL.n603 185
R136 VTAIL.n602 VTAIL.n601 185
R137 VTAIL.n593 VTAIL.n592 185
R138 VTAIL.n596 VTAIL.n595 185
R139 VTAIL.n559 VTAIL.n558 185
R140 VTAIL.n557 VTAIL.n556 185
R141 VTAIL.n474 VTAIL.n473 185
R142 VTAIL.n551 VTAIL.n550 185
R143 VTAIL.n549 VTAIL.n548 185
R144 VTAIL.n547 VTAIL.n477 185
R145 VTAIL.n481 VTAIL.n478 185
R146 VTAIL.n542 VTAIL.n541 185
R147 VTAIL.n540 VTAIL.n539 185
R148 VTAIL.n483 VTAIL.n482 185
R149 VTAIL.n534 VTAIL.n533 185
R150 VTAIL.n532 VTAIL.n531 185
R151 VTAIL.n487 VTAIL.n486 185
R152 VTAIL.n526 VTAIL.n525 185
R153 VTAIL.n524 VTAIL.n523 185
R154 VTAIL.n491 VTAIL.n490 185
R155 VTAIL.n518 VTAIL.n517 185
R156 VTAIL.n516 VTAIL.n515 185
R157 VTAIL.n495 VTAIL.n494 185
R158 VTAIL.n510 VTAIL.n509 185
R159 VTAIL.n508 VTAIL.n507 185
R160 VTAIL.n499 VTAIL.n498 185
R161 VTAIL.n502 VTAIL.n501 185
R162 VTAIL.n465 VTAIL.n464 185
R163 VTAIL.n463 VTAIL.n462 185
R164 VTAIL.n380 VTAIL.n379 185
R165 VTAIL.n457 VTAIL.n456 185
R166 VTAIL.n455 VTAIL.n454 185
R167 VTAIL.n453 VTAIL.n383 185
R168 VTAIL.n387 VTAIL.n384 185
R169 VTAIL.n448 VTAIL.n447 185
R170 VTAIL.n446 VTAIL.n445 185
R171 VTAIL.n389 VTAIL.n388 185
R172 VTAIL.n440 VTAIL.n439 185
R173 VTAIL.n438 VTAIL.n437 185
R174 VTAIL.n393 VTAIL.n392 185
R175 VTAIL.n432 VTAIL.n431 185
R176 VTAIL.n430 VTAIL.n429 185
R177 VTAIL.n397 VTAIL.n396 185
R178 VTAIL.n424 VTAIL.n423 185
R179 VTAIL.n422 VTAIL.n421 185
R180 VTAIL.n401 VTAIL.n400 185
R181 VTAIL.n416 VTAIL.n415 185
R182 VTAIL.n414 VTAIL.n413 185
R183 VTAIL.n405 VTAIL.n404 185
R184 VTAIL.n408 VTAIL.n407 185
R185 VTAIL.n371 VTAIL.n370 185
R186 VTAIL.n369 VTAIL.n368 185
R187 VTAIL.n286 VTAIL.n285 185
R188 VTAIL.n363 VTAIL.n362 185
R189 VTAIL.n361 VTAIL.n360 185
R190 VTAIL.n359 VTAIL.n289 185
R191 VTAIL.n293 VTAIL.n290 185
R192 VTAIL.n354 VTAIL.n353 185
R193 VTAIL.n352 VTAIL.n351 185
R194 VTAIL.n295 VTAIL.n294 185
R195 VTAIL.n346 VTAIL.n345 185
R196 VTAIL.n344 VTAIL.n343 185
R197 VTAIL.n299 VTAIL.n298 185
R198 VTAIL.n338 VTAIL.n337 185
R199 VTAIL.n336 VTAIL.n335 185
R200 VTAIL.n303 VTAIL.n302 185
R201 VTAIL.n330 VTAIL.n329 185
R202 VTAIL.n328 VTAIL.n327 185
R203 VTAIL.n307 VTAIL.n306 185
R204 VTAIL.n322 VTAIL.n321 185
R205 VTAIL.n320 VTAIL.n319 185
R206 VTAIL.n311 VTAIL.n310 185
R207 VTAIL.n314 VTAIL.n313 185
R208 VTAIL.t5 VTAIL.n594 147.659
R209 VTAIL.t7 VTAIL.n500 147.659
R210 VTAIL.t0 VTAIL.n406 147.659
R211 VTAIL.t3 VTAIL.n312 147.659
R212 VTAIL.t1 VTAIL.n687 147.659
R213 VTAIL.t2 VTAIL.n29 147.659
R214 VTAIL.t6 VTAIL.n123 147.659
R215 VTAIL.t4 VTAIL.n217 147.659
R216 VTAIL.n688 VTAIL.n685 104.615
R217 VTAIL.n695 VTAIL.n685 104.615
R218 VTAIL.n696 VTAIL.n695 104.615
R219 VTAIL.n696 VTAIL.n681 104.615
R220 VTAIL.n703 VTAIL.n681 104.615
R221 VTAIL.n704 VTAIL.n703 104.615
R222 VTAIL.n704 VTAIL.n677 104.615
R223 VTAIL.n711 VTAIL.n677 104.615
R224 VTAIL.n712 VTAIL.n711 104.615
R225 VTAIL.n712 VTAIL.n673 104.615
R226 VTAIL.n719 VTAIL.n673 104.615
R227 VTAIL.n720 VTAIL.n719 104.615
R228 VTAIL.n720 VTAIL.n669 104.615
R229 VTAIL.n727 VTAIL.n669 104.615
R230 VTAIL.n729 VTAIL.n727 104.615
R231 VTAIL.n729 VTAIL.n728 104.615
R232 VTAIL.n728 VTAIL.n665 104.615
R233 VTAIL.n737 VTAIL.n665 104.615
R234 VTAIL.n738 VTAIL.n737 104.615
R235 VTAIL.n738 VTAIL.n661 104.615
R236 VTAIL.n745 VTAIL.n661 104.615
R237 VTAIL.n746 VTAIL.n745 104.615
R238 VTAIL.n30 VTAIL.n27 104.615
R239 VTAIL.n37 VTAIL.n27 104.615
R240 VTAIL.n38 VTAIL.n37 104.615
R241 VTAIL.n38 VTAIL.n23 104.615
R242 VTAIL.n45 VTAIL.n23 104.615
R243 VTAIL.n46 VTAIL.n45 104.615
R244 VTAIL.n46 VTAIL.n19 104.615
R245 VTAIL.n53 VTAIL.n19 104.615
R246 VTAIL.n54 VTAIL.n53 104.615
R247 VTAIL.n54 VTAIL.n15 104.615
R248 VTAIL.n61 VTAIL.n15 104.615
R249 VTAIL.n62 VTAIL.n61 104.615
R250 VTAIL.n62 VTAIL.n11 104.615
R251 VTAIL.n69 VTAIL.n11 104.615
R252 VTAIL.n71 VTAIL.n69 104.615
R253 VTAIL.n71 VTAIL.n70 104.615
R254 VTAIL.n70 VTAIL.n7 104.615
R255 VTAIL.n79 VTAIL.n7 104.615
R256 VTAIL.n80 VTAIL.n79 104.615
R257 VTAIL.n80 VTAIL.n3 104.615
R258 VTAIL.n87 VTAIL.n3 104.615
R259 VTAIL.n88 VTAIL.n87 104.615
R260 VTAIL.n124 VTAIL.n121 104.615
R261 VTAIL.n131 VTAIL.n121 104.615
R262 VTAIL.n132 VTAIL.n131 104.615
R263 VTAIL.n132 VTAIL.n117 104.615
R264 VTAIL.n139 VTAIL.n117 104.615
R265 VTAIL.n140 VTAIL.n139 104.615
R266 VTAIL.n140 VTAIL.n113 104.615
R267 VTAIL.n147 VTAIL.n113 104.615
R268 VTAIL.n148 VTAIL.n147 104.615
R269 VTAIL.n148 VTAIL.n109 104.615
R270 VTAIL.n155 VTAIL.n109 104.615
R271 VTAIL.n156 VTAIL.n155 104.615
R272 VTAIL.n156 VTAIL.n105 104.615
R273 VTAIL.n163 VTAIL.n105 104.615
R274 VTAIL.n165 VTAIL.n163 104.615
R275 VTAIL.n165 VTAIL.n164 104.615
R276 VTAIL.n164 VTAIL.n101 104.615
R277 VTAIL.n173 VTAIL.n101 104.615
R278 VTAIL.n174 VTAIL.n173 104.615
R279 VTAIL.n174 VTAIL.n97 104.615
R280 VTAIL.n181 VTAIL.n97 104.615
R281 VTAIL.n182 VTAIL.n181 104.615
R282 VTAIL.n218 VTAIL.n215 104.615
R283 VTAIL.n225 VTAIL.n215 104.615
R284 VTAIL.n226 VTAIL.n225 104.615
R285 VTAIL.n226 VTAIL.n211 104.615
R286 VTAIL.n233 VTAIL.n211 104.615
R287 VTAIL.n234 VTAIL.n233 104.615
R288 VTAIL.n234 VTAIL.n207 104.615
R289 VTAIL.n241 VTAIL.n207 104.615
R290 VTAIL.n242 VTAIL.n241 104.615
R291 VTAIL.n242 VTAIL.n203 104.615
R292 VTAIL.n249 VTAIL.n203 104.615
R293 VTAIL.n250 VTAIL.n249 104.615
R294 VTAIL.n250 VTAIL.n199 104.615
R295 VTAIL.n257 VTAIL.n199 104.615
R296 VTAIL.n259 VTAIL.n257 104.615
R297 VTAIL.n259 VTAIL.n258 104.615
R298 VTAIL.n258 VTAIL.n195 104.615
R299 VTAIL.n267 VTAIL.n195 104.615
R300 VTAIL.n268 VTAIL.n267 104.615
R301 VTAIL.n268 VTAIL.n191 104.615
R302 VTAIL.n275 VTAIL.n191 104.615
R303 VTAIL.n276 VTAIL.n275 104.615
R304 VTAIL.n652 VTAIL.n651 104.615
R305 VTAIL.n651 VTAIL.n567 104.615
R306 VTAIL.n644 VTAIL.n567 104.615
R307 VTAIL.n644 VTAIL.n643 104.615
R308 VTAIL.n643 VTAIL.n571 104.615
R309 VTAIL.n575 VTAIL.n571 104.615
R310 VTAIL.n635 VTAIL.n575 104.615
R311 VTAIL.n635 VTAIL.n634 104.615
R312 VTAIL.n634 VTAIL.n576 104.615
R313 VTAIL.n627 VTAIL.n576 104.615
R314 VTAIL.n627 VTAIL.n626 104.615
R315 VTAIL.n626 VTAIL.n580 104.615
R316 VTAIL.n619 VTAIL.n580 104.615
R317 VTAIL.n619 VTAIL.n618 104.615
R318 VTAIL.n618 VTAIL.n584 104.615
R319 VTAIL.n611 VTAIL.n584 104.615
R320 VTAIL.n611 VTAIL.n610 104.615
R321 VTAIL.n610 VTAIL.n588 104.615
R322 VTAIL.n603 VTAIL.n588 104.615
R323 VTAIL.n603 VTAIL.n602 104.615
R324 VTAIL.n602 VTAIL.n592 104.615
R325 VTAIL.n595 VTAIL.n592 104.615
R326 VTAIL.n558 VTAIL.n557 104.615
R327 VTAIL.n557 VTAIL.n473 104.615
R328 VTAIL.n550 VTAIL.n473 104.615
R329 VTAIL.n550 VTAIL.n549 104.615
R330 VTAIL.n549 VTAIL.n477 104.615
R331 VTAIL.n481 VTAIL.n477 104.615
R332 VTAIL.n541 VTAIL.n481 104.615
R333 VTAIL.n541 VTAIL.n540 104.615
R334 VTAIL.n540 VTAIL.n482 104.615
R335 VTAIL.n533 VTAIL.n482 104.615
R336 VTAIL.n533 VTAIL.n532 104.615
R337 VTAIL.n532 VTAIL.n486 104.615
R338 VTAIL.n525 VTAIL.n486 104.615
R339 VTAIL.n525 VTAIL.n524 104.615
R340 VTAIL.n524 VTAIL.n490 104.615
R341 VTAIL.n517 VTAIL.n490 104.615
R342 VTAIL.n517 VTAIL.n516 104.615
R343 VTAIL.n516 VTAIL.n494 104.615
R344 VTAIL.n509 VTAIL.n494 104.615
R345 VTAIL.n509 VTAIL.n508 104.615
R346 VTAIL.n508 VTAIL.n498 104.615
R347 VTAIL.n501 VTAIL.n498 104.615
R348 VTAIL.n464 VTAIL.n463 104.615
R349 VTAIL.n463 VTAIL.n379 104.615
R350 VTAIL.n456 VTAIL.n379 104.615
R351 VTAIL.n456 VTAIL.n455 104.615
R352 VTAIL.n455 VTAIL.n383 104.615
R353 VTAIL.n387 VTAIL.n383 104.615
R354 VTAIL.n447 VTAIL.n387 104.615
R355 VTAIL.n447 VTAIL.n446 104.615
R356 VTAIL.n446 VTAIL.n388 104.615
R357 VTAIL.n439 VTAIL.n388 104.615
R358 VTAIL.n439 VTAIL.n438 104.615
R359 VTAIL.n438 VTAIL.n392 104.615
R360 VTAIL.n431 VTAIL.n392 104.615
R361 VTAIL.n431 VTAIL.n430 104.615
R362 VTAIL.n430 VTAIL.n396 104.615
R363 VTAIL.n423 VTAIL.n396 104.615
R364 VTAIL.n423 VTAIL.n422 104.615
R365 VTAIL.n422 VTAIL.n400 104.615
R366 VTAIL.n415 VTAIL.n400 104.615
R367 VTAIL.n415 VTAIL.n414 104.615
R368 VTAIL.n414 VTAIL.n404 104.615
R369 VTAIL.n407 VTAIL.n404 104.615
R370 VTAIL.n370 VTAIL.n369 104.615
R371 VTAIL.n369 VTAIL.n285 104.615
R372 VTAIL.n362 VTAIL.n285 104.615
R373 VTAIL.n362 VTAIL.n361 104.615
R374 VTAIL.n361 VTAIL.n289 104.615
R375 VTAIL.n293 VTAIL.n289 104.615
R376 VTAIL.n353 VTAIL.n293 104.615
R377 VTAIL.n353 VTAIL.n352 104.615
R378 VTAIL.n352 VTAIL.n294 104.615
R379 VTAIL.n345 VTAIL.n294 104.615
R380 VTAIL.n345 VTAIL.n344 104.615
R381 VTAIL.n344 VTAIL.n298 104.615
R382 VTAIL.n337 VTAIL.n298 104.615
R383 VTAIL.n337 VTAIL.n336 104.615
R384 VTAIL.n336 VTAIL.n302 104.615
R385 VTAIL.n329 VTAIL.n302 104.615
R386 VTAIL.n329 VTAIL.n328 104.615
R387 VTAIL.n328 VTAIL.n306 104.615
R388 VTAIL.n321 VTAIL.n306 104.615
R389 VTAIL.n321 VTAIL.n320 104.615
R390 VTAIL.n320 VTAIL.n310 104.615
R391 VTAIL.n313 VTAIL.n310 104.615
R392 VTAIL.n688 VTAIL.t1 52.3082
R393 VTAIL.n30 VTAIL.t2 52.3082
R394 VTAIL.n124 VTAIL.t6 52.3082
R395 VTAIL.n218 VTAIL.t4 52.3082
R396 VTAIL.n595 VTAIL.t5 52.3082
R397 VTAIL.n501 VTAIL.t7 52.3082
R398 VTAIL.n407 VTAIL.t0 52.3082
R399 VTAIL.n313 VTAIL.t3 52.3082
R400 VTAIL.n751 VTAIL.n750 34.5126
R401 VTAIL.n93 VTAIL.n92 34.5126
R402 VTAIL.n187 VTAIL.n186 34.5126
R403 VTAIL.n281 VTAIL.n280 34.5126
R404 VTAIL.n657 VTAIL.n656 34.5126
R405 VTAIL.n563 VTAIL.n562 34.5126
R406 VTAIL.n469 VTAIL.n468 34.5126
R407 VTAIL.n375 VTAIL.n374 34.5126
R408 VTAIL.n751 VTAIL.n657 28.1514
R409 VTAIL.n375 VTAIL.n281 28.1514
R410 VTAIL.n689 VTAIL.n687 15.6677
R411 VTAIL.n31 VTAIL.n29 15.6677
R412 VTAIL.n125 VTAIL.n123 15.6677
R413 VTAIL.n219 VTAIL.n217 15.6677
R414 VTAIL.n596 VTAIL.n594 15.6677
R415 VTAIL.n502 VTAIL.n500 15.6677
R416 VTAIL.n408 VTAIL.n406 15.6677
R417 VTAIL.n314 VTAIL.n312 15.6677
R418 VTAIL.n736 VTAIL.n735 13.1884
R419 VTAIL.n78 VTAIL.n77 13.1884
R420 VTAIL.n172 VTAIL.n171 13.1884
R421 VTAIL.n266 VTAIL.n265 13.1884
R422 VTAIL.n642 VTAIL.n641 13.1884
R423 VTAIL.n548 VTAIL.n547 13.1884
R424 VTAIL.n454 VTAIL.n453 13.1884
R425 VTAIL.n360 VTAIL.n359 13.1884
R426 VTAIL.n690 VTAIL.n686 12.8005
R427 VTAIL.n734 VTAIL.n666 12.8005
R428 VTAIL.n739 VTAIL.n664 12.8005
R429 VTAIL.n32 VTAIL.n28 12.8005
R430 VTAIL.n76 VTAIL.n8 12.8005
R431 VTAIL.n81 VTAIL.n6 12.8005
R432 VTAIL.n126 VTAIL.n122 12.8005
R433 VTAIL.n170 VTAIL.n102 12.8005
R434 VTAIL.n175 VTAIL.n100 12.8005
R435 VTAIL.n220 VTAIL.n216 12.8005
R436 VTAIL.n264 VTAIL.n196 12.8005
R437 VTAIL.n269 VTAIL.n194 12.8005
R438 VTAIL.n645 VTAIL.n570 12.8005
R439 VTAIL.n640 VTAIL.n572 12.8005
R440 VTAIL.n597 VTAIL.n593 12.8005
R441 VTAIL.n551 VTAIL.n476 12.8005
R442 VTAIL.n546 VTAIL.n478 12.8005
R443 VTAIL.n503 VTAIL.n499 12.8005
R444 VTAIL.n457 VTAIL.n382 12.8005
R445 VTAIL.n452 VTAIL.n384 12.8005
R446 VTAIL.n409 VTAIL.n405 12.8005
R447 VTAIL.n363 VTAIL.n288 12.8005
R448 VTAIL.n358 VTAIL.n290 12.8005
R449 VTAIL.n315 VTAIL.n311 12.8005
R450 VTAIL.n694 VTAIL.n693 12.0247
R451 VTAIL.n731 VTAIL.n730 12.0247
R452 VTAIL.n740 VTAIL.n662 12.0247
R453 VTAIL.n36 VTAIL.n35 12.0247
R454 VTAIL.n73 VTAIL.n72 12.0247
R455 VTAIL.n82 VTAIL.n4 12.0247
R456 VTAIL.n130 VTAIL.n129 12.0247
R457 VTAIL.n167 VTAIL.n166 12.0247
R458 VTAIL.n176 VTAIL.n98 12.0247
R459 VTAIL.n224 VTAIL.n223 12.0247
R460 VTAIL.n261 VTAIL.n260 12.0247
R461 VTAIL.n270 VTAIL.n192 12.0247
R462 VTAIL.n646 VTAIL.n568 12.0247
R463 VTAIL.n637 VTAIL.n636 12.0247
R464 VTAIL.n601 VTAIL.n600 12.0247
R465 VTAIL.n552 VTAIL.n474 12.0247
R466 VTAIL.n543 VTAIL.n542 12.0247
R467 VTAIL.n507 VTAIL.n506 12.0247
R468 VTAIL.n458 VTAIL.n380 12.0247
R469 VTAIL.n449 VTAIL.n448 12.0247
R470 VTAIL.n413 VTAIL.n412 12.0247
R471 VTAIL.n364 VTAIL.n286 12.0247
R472 VTAIL.n355 VTAIL.n354 12.0247
R473 VTAIL.n319 VTAIL.n318 12.0247
R474 VTAIL.n697 VTAIL.n684 11.249
R475 VTAIL.n726 VTAIL.n668 11.249
R476 VTAIL.n744 VTAIL.n743 11.249
R477 VTAIL.n39 VTAIL.n26 11.249
R478 VTAIL.n68 VTAIL.n10 11.249
R479 VTAIL.n86 VTAIL.n85 11.249
R480 VTAIL.n133 VTAIL.n120 11.249
R481 VTAIL.n162 VTAIL.n104 11.249
R482 VTAIL.n180 VTAIL.n179 11.249
R483 VTAIL.n227 VTAIL.n214 11.249
R484 VTAIL.n256 VTAIL.n198 11.249
R485 VTAIL.n274 VTAIL.n273 11.249
R486 VTAIL.n650 VTAIL.n649 11.249
R487 VTAIL.n633 VTAIL.n574 11.249
R488 VTAIL.n604 VTAIL.n591 11.249
R489 VTAIL.n556 VTAIL.n555 11.249
R490 VTAIL.n539 VTAIL.n480 11.249
R491 VTAIL.n510 VTAIL.n497 11.249
R492 VTAIL.n462 VTAIL.n461 11.249
R493 VTAIL.n445 VTAIL.n386 11.249
R494 VTAIL.n416 VTAIL.n403 11.249
R495 VTAIL.n368 VTAIL.n367 11.249
R496 VTAIL.n351 VTAIL.n292 11.249
R497 VTAIL.n322 VTAIL.n309 11.249
R498 VTAIL.n698 VTAIL.n682 10.4732
R499 VTAIL.n725 VTAIL.n670 10.4732
R500 VTAIL.n747 VTAIL.n660 10.4732
R501 VTAIL.n40 VTAIL.n24 10.4732
R502 VTAIL.n67 VTAIL.n12 10.4732
R503 VTAIL.n89 VTAIL.n2 10.4732
R504 VTAIL.n134 VTAIL.n118 10.4732
R505 VTAIL.n161 VTAIL.n106 10.4732
R506 VTAIL.n183 VTAIL.n96 10.4732
R507 VTAIL.n228 VTAIL.n212 10.4732
R508 VTAIL.n255 VTAIL.n200 10.4732
R509 VTAIL.n277 VTAIL.n190 10.4732
R510 VTAIL.n653 VTAIL.n566 10.4732
R511 VTAIL.n632 VTAIL.n577 10.4732
R512 VTAIL.n605 VTAIL.n589 10.4732
R513 VTAIL.n559 VTAIL.n472 10.4732
R514 VTAIL.n538 VTAIL.n483 10.4732
R515 VTAIL.n511 VTAIL.n495 10.4732
R516 VTAIL.n465 VTAIL.n378 10.4732
R517 VTAIL.n444 VTAIL.n389 10.4732
R518 VTAIL.n417 VTAIL.n401 10.4732
R519 VTAIL.n371 VTAIL.n284 10.4732
R520 VTAIL.n350 VTAIL.n295 10.4732
R521 VTAIL.n323 VTAIL.n307 10.4732
R522 VTAIL.n702 VTAIL.n701 9.69747
R523 VTAIL.n722 VTAIL.n721 9.69747
R524 VTAIL.n748 VTAIL.n658 9.69747
R525 VTAIL.n44 VTAIL.n43 9.69747
R526 VTAIL.n64 VTAIL.n63 9.69747
R527 VTAIL.n90 VTAIL.n0 9.69747
R528 VTAIL.n138 VTAIL.n137 9.69747
R529 VTAIL.n158 VTAIL.n157 9.69747
R530 VTAIL.n184 VTAIL.n94 9.69747
R531 VTAIL.n232 VTAIL.n231 9.69747
R532 VTAIL.n252 VTAIL.n251 9.69747
R533 VTAIL.n278 VTAIL.n188 9.69747
R534 VTAIL.n654 VTAIL.n564 9.69747
R535 VTAIL.n629 VTAIL.n628 9.69747
R536 VTAIL.n609 VTAIL.n608 9.69747
R537 VTAIL.n560 VTAIL.n470 9.69747
R538 VTAIL.n535 VTAIL.n534 9.69747
R539 VTAIL.n515 VTAIL.n514 9.69747
R540 VTAIL.n466 VTAIL.n376 9.69747
R541 VTAIL.n441 VTAIL.n440 9.69747
R542 VTAIL.n421 VTAIL.n420 9.69747
R543 VTAIL.n372 VTAIL.n282 9.69747
R544 VTAIL.n347 VTAIL.n346 9.69747
R545 VTAIL.n327 VTAIL.n326 9.69747
R546 VTAIL.n750 VTAIL.n749 9.45567
R547 VTAIL.n92 VTAIL.n91 9.45567
R548 VTAIL.n186 VTAIL.n185 9.45567
R549 VTAIL.n280 VTAIL.n279 9.45567
R550 VTAIL.n656 VTAIL.n655 9.45567
R551 VTAIL.n562 VTAIL.n561 9.45567
R552 VTAIL.n468 VTAIL.n467 9.45567
R553 VTAIL.n374 VTAIL.n373 9.45567
R554 VTAIL.n749 VTAIL.n748 9.3005
R555 VTAIL.n660 VTAIL.n659 9.3005
R556 VTAIL.n743 VTAIL.n742 9.3005
R557 VTAIL.n741 VTAIL.n740 9.3005
R558 VTAIL.n664 VTAIL.n663 9.3005
R559 VTAIL.n709 VTAIL.n708 9.3005
R560 VTAIL.n707 VTAIL.n706 9.3005
R561 VTAIL.n680 VTAIL.n679 9.3005
R562 VTAIL.n701 VTAIL.n700 9.3005
R563 VTAIL.n699 VTAIL.n698 9.3005
R564 VTAIL.n684 VTAIL.n683 9.3005
R565 VTAIL.n693 VTAIL.n692 9.3005
R566 VTAIL.n691 VTAIL.n690 9.3005
R567 VTAIL.n676 VTAIL.n675 9.3005
R568 VTAIL.n715 VTAIL.n714 9.3005
R569 VTAIL.n717 VTAIL.n716 9.3005
R570 VTAIL.n672 VTAIL.n671 9.3005
R571 VTAIL.n723 VTAIL.n722 9.3005
R572 VTAIL.n725 VTAIL.n724 9.3005
R573 VTAIL.n668 VTAIL.n667 9.3005
R574 VTAIL.n732 VTAIL.n731 9.3005
R575 VTAIL.n734 VTAIL.n733 9.3005
R576 VTAIL.n91 VTAIL.n90 9.3005
R577 VTAIL.n2 VTAIL.n1 9.3005
R578 VTAIL.n85 VTAIL.n84 9.3005
R579 VTAIL.n83 VTAIL.n82 9.3005
R580 VTAIL.n6 VTAIL.n5 9.3005
R581 VTAIL.n51 VTAIL.n50 9.3005
R582 VTAIL.n49 VTAIL.n48 9.3005
R583 VTAIL.n22 VTAIL.n21 9.3005
R584 VTAIL.n43 VTAIL.n42 9.3005
R585 VTAIL.n41 VTAIL.n40 9.3005
R586 VTAIL.n26 VTAIL.n25 9.3005
R587 VTAIL.n35 VTAIL.n34 9.3005
R588 VTAIL.n33 VTAIL.n32 9.3005
R589 VTAIL.n18 VTAIL.n17 9.3005
R590 VTAIL.n57 VTAIL.n56 9.3005
R591 VTAIL.n59 VTAIL.n58 9.3005
R592 VTAIL.n14 VTAIL.n13 9.3005
R593 VTAIL.n65 VTAIL.n64 9.3005
R594 VTAIL.n67 VTAIL.n66 9.3005
R595 VTAIL.n10 VTAIL.n9 9.3005
R596 VTAIL.n74 VTAIL.n73 9.3005
R597 VTAIL.n76 VTAIL.n75 9.3005
R598 VTAIL.n185 VTAIL.n184 9.3005
R599 VTAIL.n96 VTAIL.n95 9.3005
R600 VTAIL.n179 VTAIL.n178 9.3005
R601 VTAIL.n177 VTAIL.n176 9.3005
R602 VTAIL.n100 VTAIL.n99 9.3005
R603 VTAIL.n145 VTAIL.n144 9.3005
R604 VTAIL.n143 VTAIL.n142 9.3005
R605 VTAIL.n116 VTAIL.n115 9.3005
R606 VTAIL.n137 VTAIL.n136 9.3005
R607 VTAIL.n135 VTAIL.n134 9.3005
R608 VTAIL.n120 VTAIL.n119 9.3005
R609 VTAIL.n129 VTAIL.n128 9.3005
R610 VTAIL.n127 VTAIL.n126 9.3005
R611 VTAIL.n112 VTAIL.n111 9.3005
R612 VTAIL.n151 VTAIL.n150 9.3005
R613 VTAIL.n153 VTAIL.n152 9.3005
R614 VTAIL.n108 VTAIL.n107 9.3005
R615 VTAIL.n159 VTAIL.n158 9.3005
R616 VTAIL.n161 VTAIL.n160 9.3005
R617 VTAIL.n104 VTAIL.n103 9.3005
R618 VTAIL.n168 VTAIL.n167 9.3005
R619 VTAIL.n170 VTAIL.n169 9.3005
R620 VTAIL.n279 VTAIL.n278 9.3005
R621 VTAIL.n190 VTAIL.n189 9.3005
R622 VTAIL.n273 VTAIL.n272 9.3005
R623 VTAIL.n271 VTAIL.n270 9.3005
R624 VTAIL.n194 VTAIL.n193 9.3005
R625 VTAIL.n239 VTAIL.n238 9.3005
R626 VTAIL.n237 VTAIL.n236 9.3005
R627 VTAIL.n210 VTAIL.n209 9.3005
R628 VTAIL.n231 VTAIL.n230 9.3005
R629 VTAIL.n229 VTAIL.n228 9.3005
R630 VTAIL.n214 VTAIL.n213 9.3005
R631 VTAIL.n223 VTAIL.n222 9.3005
R632 VTAIL.n221 VTAIL.n220 9.3005
R633 VTAIL.n206 VTAIL.n205 9.3005
R634 VTAIL.n245 VTAIL.n244 9.3005
R635 VTAIL.n247 VTAIL.n246 9.3005
R636 VTAIL.n202 VTAIL.n201 9.3005
R637 VTAIL.n253 VTAIL.n252 9.3005
R638 VTAIL.n255 VTAIL.n254 9.3005
R639 VTAIL.n198 VTAIL.n197 9.3005
R640 VTAIL.n262 VTAIL.n261 9.3005
R641 VTAIL.n264 VTAIL.n263 9.3005
R642 VTAIL.n622 VTAIL.n621 9.3005
R643 VTAIL.n624 VTAIL.n623 9.3005
R644 VTAIL.n579 VTAIL.n578 9.3005
R645 VTAIL.n630 VTAIL.n629 9.3005
R646 VTAIL.n632 VTAIL.n631 9.3005
R647 VTAIL.n574 VTAIL.n573 9.3005
R648 VTAIL.n638 VTAIL.n637 9.3005
R649 VTAIL.n640 VTAIL.n639 9.3005
R650 VTAIL.n655 VTAIL.n654 9.3005
R651 VTAIL.n566 VTAIL.n565 9.3005
R652 VTAIL.n649 VTAIL.n648 9.3005
R653 VTAIL.n647 VTAIL.n646 9.3005
R654 VTAIL.n570 VTAIL.n569 9.3005
R655 VTAIL.n583 VTAIL.n582 9.3005
R656 VTAIL.n616 VTAIL.n615 9.3005
R657 VTAIL.n614 VTAIL.n613 9.3005
R658 VTAIL.n587 VTAIL.n586 9.3005
R659 VTAIL.n608 VTAIL.n607 9.3005
R660 VTAIL.n606 VTAIL.n605 9.3005
R661 VTAIL.n591 VTAIL.n590 9.3005
R662 VTAIL.n600 VTAIL.n599 9.3005
R663 VTAIL.n598 VTAIL.n597 9.3005
R664 VTAIL.n528 VTAIL.n527 9.3005
R665 VTAIL.n530 VTAIL.n529 9.3005
R666 VTAIL.n485 VTAIL.n484 9.3005
R667 VTAIL.n536 VTAIL.n535 9.3005
R668 VTAIL.n538 VTAIL.n537 9.3005
R669 VTAIL.n480 VTAIL.n479 9.3005
R670 VTAIL.n544 VTAIL.n543 9.3005
R671 VTAIL.n546 VTAIL.n545 9.3005
R672 VTAIL.n561 VTAIL.n560 9.3005
R673 VTAIL.n472 VTAIL.n471 9.3005
R674 VTAIL.n555 VTAIL.n554 9.3005
R675 VTAIL.n553 VTAIL.n552 9.3005
R676 VTAIL.n476 VTAIL.n475 9.3005
R677 VTAIL.n489 VTAIL.n488 9.3005
R678 VTAIL.n522 VTAIL.n521 9.3005
R679 VTAIL.n520 VTAIL.n519 9.3005
R680 VTAIL.n493 VTAIL.n492 9.3005
R681 VTAIL.n514 VTAIL.n513 9.3005
R682 VTAIL.n512 VTAIL.n511 9.3005
R683 VTAIL.n497 VTAIL.n496 9.3005
R684 VTAIL.n506 VTAIL.n505 9.3005
R685 VTAIL.n504 VTAIL.n503 9.3005
R686 VTAIL.n434 VTAIL.n433 9.3005
R687 VTAIL.n436 VTAIL.n435 9.3005
R688 VTAIL.n391 VTAIL.n390 9.3005
R689 VTAIL.n442 VTAIL.n441 9.3005
R690 VTAIL.n444 VTAIL.n443 9.3005
R691 VTAIL.n386 VTAIL.n385 9.3005
R692 VTAIL.n450 VTAIL.n449 9.3005
R693 VTAIL.n452 VTAIL.n451 9.3005
R694 VTAIL.n467 VTAIL.n466 9.3005
R695 VTAIL.n378 VTAIL.n377 9.3005
R696 VTAIL.n461 VTAIL.n460 9.3005
R697 VTAIL.n459 VTAIL.n458 9.3005
R698 VTAIL.n382 VTAIL.n381 9.3005
R699 VTAIL.n395 VTAIL.n394 9.3005
R700 VTAIL.n428 VTAIL.n427 9.3005
R701 VTAIL.n426 VTAIL.n425 9.3005
R702 VTAIL.n399 VTAIL.n398 9.3005
R703 VTAIL.n420 VTAIL.n419 9.3005
R704 VTAIL.n418 VTAIL.n417 9.3005
R705 VTAIL.n403 VTAIL.n402 9.3005
R706 VTAIL.n412 VTAIL.n411 9.3005
R707 VTAIL.n410 VTAIL.n409 9.3005
R708 VTAIL.n340 VTAIL.n339 9.3005
R709 VTAIL.n342 VTAIL.n341 9.3005
R710 VTAIL.n297 VTAIL.n296 9.3005
R711 VTAIL.n348 VTAIL.n347 9.3005
R712 VTAIL.n350 VTAIL.n349 9.3005
R713 VTAIL.n292 VTAIL.n291 9.3005
R714 VTAIL.n356 VTAIL.n355 9.3005
R715 VTAIL.n358 VTAIL.n357 9.3005
R716 VTAIL.n373 VTAIL.n372 9.3005
R717 VTAIL.n284 VTAIL.n283 9.3005
R718 VTAIL.n367 VTAIL.n366 9.3005
R719 VTAIL.n365 VTAIL.n364 9.3005
R720 VTAIL.n288 VTAIL.n287 9.3005
R721 VTAIL.n301 VTAIL.n300 9.3005
R722 VTAIL.n334 VTAIL.n333 9.3005
R723 VTAIL.n332 VTAIL.n331 9.3005
R724 VTAIL.n305 VTAIL.n304 9.3005
R725 VTAIL.n326 VTAIL.n325 9.3005
R726 VTAIL.n324 VTAIL.n323 9.3005
R727 VTAIL.n309 VTAIL.n308 9.3005
R728 VTAIL.n318 VTAIL.n317 9.3005
R729 VTAIL.n316 VTAIL.n315 9.3005
R730 VTAIL.n705 VTAIL.n680 8.92171
R731 VTAIL.n718 VTAIL.n672 8.92171
R732 VTAIL.n47 VTAIL.n22 8.92171
R733 VTAIL.n60 VTAIL.n14 8.92171
R734 VTAIL.n141 VTAIL.n116 8.92171
R735 VTAIL.n154 VTAIL.n108 8.92171
R736 VTAIL.n235 VTAIL.n210 8.92171
R737 VTAIL.n248 VTAIL.n202 8.92171
R738 VTAIL.n625 VTAIL.n579 8.92171
R739 VTAIL.n612 VTAIL.n587 8.92171
R740 VTAIL.n531 VTAIL.n485 8.92171
R741 VTAIL.n518 VTAIL.n493 8.92171
R742 VTAIL.n437 VTAIL.n391 8.92171
R743 VTAIL.n424 VTAIL.n399 8.92171
R744 VTAIL.n343 VTAIL.n297 8.92171
R745 VTAIL.n330 VTAIL.n305 8.92171
R746 VTAIL.n706 VTAIL.n678 8.14595
R747 VTAIL.n717 VTAIL.n674 8.14595
R748 VTAIL.n48 VTAIL.n20 8.14595
R749 VTAIL.n59 VTAIL.n16 8.14595
R750 VTAIL.n142 VTAIL.n114 8.14595
R751 VTAIL.n153 VTAIL.n110 8.14595
R752 VTAIL.n236 VTAIL.n208 8.14595
R753 VTAIL.n247 VTAIL.n204 8.14595
R754 VTAIL.n624 VTAIL.n581 8.14595
R755 VTAIL.n613 VTAIL.n585 8.14595
R756 VTAIL.n530 VTAIL.n487 8.14595
R757 VTAIL.n519 VTAIL.n491 8.14595
R758 VTAIL.n436 VTAIL.n393 8.14595
R759 VTAIL.n425 VTAIL.n397 8.14595
R760 VTAIL.n342 VTAIL.n299 8.14595
R761 VTAIL.n331 VTAIL.n303 8.14595
R762 VTAIL.n710 VTAIL.n709 7.3702
R763 VTAIL.n714 VTAIL.n713 7.3702
R764 VTAIL.n52 VTAIL.n51 7.3702
R765 VTAIL.n56 VTAIL.n55 7.3702
R766 VTAIL.n146 VTAIL.n145 7.3702
R767 VTAIL.n150 VTAIL.n149 7.3702
R768 VTAIL.n240 VTAIL.n239 7.3702
R769 VTAIL.n244 VTAIL.n243 7.3702
R770 VTAIL.n621 VTAIL.n620 7.3702
R771 VTAIL.n617 VTAIL.n616 7.3702
R772 VTAIL.n527 VTAIL.n526 7.3702
R773 VTAIL.n523 VTAIL.n522 7.3702
R774 VTAIL.n433 VTAIL.n432 7.3702
R775 VTAIL.n429 VTAIL.n428 7.3702
R776 VTAIL.n339 VTAIL.n338 7.3702
R777 VTAIL.n335 VTAIL.n334 7.3702
R778 VTAIL.n710 VTAIL.n676 6.59444
R779 VTAIL.n713 VTAIL.n676 6.59444
R780 VTAIL.n52 VTAIL.n18 6.59444
R781 VTAIL.n55 VTAIL.n18 6.59444
R782 VTAIL.n146 VTAIL.n112 6.59444
R783 VTAIL.n149 VTAIL.n112 6.59444
R784 VTAIL.n240 VTAIL.n206 6.59444
R785 VTAIL.n243 VTAIL.n206 6.59444
R786 VTAIL.n620 VTAIL.n583 6.59444
R787 VTAIL.n617 VTAIL.n583 6.59444
R788 VTAIL.n526 VTAIL.n489 6.59444
R789 VTAIL.n523 VTAIL.n489 6.59444
R790 VTAIL.n432 VTAIL.n395 6.59444
R791 VTAIL.n429 VTAIL.n395 6.59444
R792 VTAIL.n338 VTAIL.n301 6.59444
R793 VTAIL.n335 VTAIL.n301 6.59444
R794 VTAIL.n709 VTAIL.n678 5.81868
R795 VTAIL.n714 VTAIL.n674 5.81868
R796 VTAIL.n51 VTAIL.n20 5.81868
R797 VTAIL.n56 VTAIL.n16 5.81868
R798 VTAIL.n145 VTAIL.n114 5.81868
R799 VTAIL.n150 VTAIL.n110 5.81868
R800 VTAIL.n239 VTAIL.n208 5.81868
R801 VTAIL.n244 VTAIL.n204 5.81868
R802 VTAIL.n621 VTAIL.n581 5.81868
R803 VTAIL.n616 VTAIL.n585 5.81868
R804 VTAIL.n527 VTAIL.n487 5.81868
R805 VTAIL.n522 VTAIL.n491 5.81868
R806 VTAIL.n433 VTAIL.n393 5.81868
R807 VTAIL.n428 VTAIL.n397 5.81868
R808 VTAIL.n339 VTAIL.n299 5.81868
R809 VTAIL.n334 VTAIL.n303 5.81868
R810 VTAIL.n706 VTAIL.n705 5.04292
R811 VTAIL.n718 VTAIL.n717 5.04292
R812 VTAIL.n48 VTAIL.n47 5.04292
R813 VTAIL.n60 VTAIL.n59 5.04292
R814 VTAIL.n142 VTAIL.n141 5.04292
R815 VTAIL.n154 VTAIL.n153 5.04292
R816 VTAIL.n236 VTAIL.n235 5.04292
R817 VTAIL.n248 VTAIL.n247 5.04292
R818 VTAIL.n625 VTAIL.n624 5.04292
R819 VTAIL.n613 VTAIL.n612 5.04292
R820 VTAIL.n531 VTAIL.n530 5.04292
R821 VTAIL.n519 VTAIL.n518 5.04292
R822 VTAIL.n437 VTAIL.n436 5.04292
R823 VTAIL.n425 VTAIL.n424 5.04292
R824 VTAIL.n343 VTAIL.n342 5.04292
R825 VTAIL.n331 VTAIL.n330 5.04292
R826 VTAIL.n598 VTAIL.n594 4.38563
R827 VTAIL.n504 VTAIL.n500 4.38563
R828 VTAIL.n410 VTAIL.n406 4.38563
R829 VTAIL.n316 VTAIL.n312 4.38563
R830 VTAIL.n691 VTAIL.n687 4.38563
R831 VTAIL.n33 VTAIL.n29 4.38563
R832 VTAIL.n127 VTAIL.n123 4.38563
R833 VTAIL.n221 VTAIL.n217 4.38563
R834 VTAIL.n702 VTAIL.n680 4.26717
R835 VTAIL.n721 VTAIL.n672 4.26717
R836 VTAIL.n750 VTAIL.n658 4.26717
R837 VTAIL.n44 VTAIL.n22 4.26717
R838 VTAIL.n63 VTAIL.n14 4.26717
R839 VTAIL.n92 VTAIL.n0 4.26717
R840 VTAIL.n138 VTAIL.n116 4.26717
R841 VTAIL.n157 VTAIL.n108 4.26717
R842 VTAIL.n186 VTAIL.n94 4.26717
R843 VTAIL.n232 VTAIL.n210 4.26717
R844 VTAIL.n251 VTAIL.n202 4.26717
R845 VTAIL.n280 VTAIL.n188 4.26717
R846 VTAIL.n656 VTAIL.n564 4.26717
R847 VTAIL.n628 VTAIL.n579 4.26717
R848 VTAIL.n609 VTAIL.n587 4.26717
R849 VTAIL.n562 VTAIL.n470 4.26717
R850 VTAIL.n534 VTAIL.n485 4.26717
R851 VTAIL.n515 VTAIL.n493 4.26717
R852 VTAIL.n468 VTAIL.n376 4.26717
R853 VTAIL.n440 VTAIL.n391 4.26717
R854 VTAIL.n421 VTAIL.n399 4.26717
R855 VTAIL.n374 VTAIL.n282 4.26717
R856 VTAIL.n346 VTAIL.n297 4.26717
R857 VTAIL.n327 VTAIL.n305 4.26717
R858 VTAIL.n701 VTAIL.n682 3.49141
R859 VTAIL.n722 VTAIL.n670 3.49141
R860 VTAIL.n748 VTAIL.n747 3.49141
R861 VTAIL.n43 VTAIL.n24 3.49141
R862 VTAIL.n64 VTAIL.n12 3.49141
R863 VTAIL.n90 VTAIL.n89 3.49141
R864 VTAIL.n137 VTAIL.n118 3.49141
R865 VTAIL.n158 VTAIL.n106 3.49141
R866 VTAIL.n184 VTAIL.n183 3.49141
R867 VTAIL.n231 VTAIL.n212 3.49141
R868 VTAIL.n252 VTAIL.n200 3.49141
R869 VTAIL.n278 VTAIL.n277 3.49141
R870 VTAIL.n654 VTAIL.n653 3.49141
R871 VTAIL.n629 VTAIL.n577 3.49141
R872 VTAIL.n608 VTAIL.n589 3.49141
R873 VTAIL.n560 VTAIL.n559 3.49141
R874 VTAIL.n535 VTAIL.n483 3.49141
R875 VTAIL.n514 VTAIL.n495 3.49141
R876 VTAIL.n466 VTAIL.n465 3.49141
R877 VTAIL.n441 VTAIL.n389 3.49141
R878 VTAIL.n420 VTAIL.n401 3.49141
R879 VTAIL.n372 VTAIL.n371 3.49141
R880 VTAIL.n347 VTAIL.n295 3.49141
R881 VTAIL.n326 VTAIL.n307 3.49141
R882 VTAIL.n698 VTAIL.n697 2.71565
R883 VTAIL.n726 VTAIL.n725 2.71565
R884 VTAIL.n744 VTAIL.n660 2.71565
R885 VTAIL.n40 VTAIL.n39 2.71565
R886 VTAIL.n68 VTAIL.n67 2.71565
R887 VTAIL.n86 VTAIL.n2 2.71565
R888 VTAIL.n134 VTAIL.n133 2.71565
R889 VTAIL.n162 VTAIL.n161 2.71565
R890 VTAIL.n180 VTAIL.n96 2.71565
R891 VTAIL.n228 VTAIL.n227 2.71565
R892 VTAIL.n256 VTAIL.n255 2.71565
R893 VTAIL.n274 VTAIL.n190 2.71565
R894 VTAIL.n650 VTAIL.n566 2.71565
R895 VTAIL.n633 VTAIL.n632 2.71565
R896 VTAIL.n605 VTAIL.n604 2.71565
R897 VTAIL.n556 VTAIL.n472 2.71565
R898 VTAIL.n539 VTAIL.n538 2.71565
R899 VTAIL.n511 VTAIL.n510 2.71565
R900 VTAIL.n462 VTAIL.n378 2.71565
R901 VTAIL.n445 VTAIL.n444 2.71565
R902 VTAIL.n417 VTAIL.n416 2.71565
R903 VTAIL.n368 VTAIL.n284 2.71565
R904 VTAIL.n351 VTAIL.n350 2.71565
R905 VTAIL.n323 VTAIL.n322 2.71565
R906 VTAIL.n694 VTAIL.n684 1.93989
R907 VTAIL.n730 VTAIL.n668 1.93989
R908 VTAIL.n743 VTAIL.n662 1.93989
R909 VTAIL.n36 VTAIL.n26 1.93989
R910 VTAIL.n72 VTAIL.n10 1.93989
R911 VTAIL.n85 VTAIL.n4 1.93989
R912 VTAIL.n130 VTAIL.n120 1.93989
R913 VTAIL.n166 VTAIL.n104 1.93989
R914 VTAIL.n179 VTAIL.n98 1.93989
R915 VTAIL.n224 VTAIL.n214 1.93989
R916 VTAIL.n260 VTAIL.n198 1.93989
R917 VTAIL.n273 VTAIL.n192 1.93989
R918 VTAIL.n649 VTAIL.n568 1.93989
R919 VTAIL.n636 VTAIL.n574 1.93989
R920 VTAIL.n601 VTAIL.n591 1.93989
R921 VTAIL.n555 VTAIL.n474 1.93989
R922 VTAIL.n542 VTAIL.n480 1.93989
R923 VTAIL.n507 VTAIL.n497 1.93989
R924 VTAIL.n461 VTAIL.n380 1.93989
R925 VTAIL.n448 VTAIL.n386 1.93989
R926 VTAIL.n413 VTAIL.n403 1.93989
R927 VTAIL.n367 VTAIL.n286 1.93989
R928 VTAIL.n354 VTAIL.n292 1.93989
R929 VTAIL.n319 VTAIL.n309 1.93989
R930 VTAIL.n469 VTAIL.n375 1.19878
R931 VTAIL.n657 VTAIL.n563 1.19878
R932 VTAIL.n281 VTAIL.n187 1.19878
R933 VTAIL.n693 VTAIL.n686 1.16414
R934 VTAIL.n731 VTAIL.n666 1.16414
R935 VTAIL.n740 VTAIL.n739 1.16414
R936 VTAIL.n35 VTAIL.n28 1.16414
R937 VTAIL.n73 VTAIL.n8 1.16414
R938 VTAIL.n82 VTAIL.n81 1.16414
R939 VTAIL.n129 VTAIL.n122 1.16414
R940 VTAIL.n167 VTAIL.n102 1.16414
R941 VTAIL.n176 VTAIL.n175 1.16414
R942 VTAIL.n223 VTAIL.n216 1.16414
R943 VTAIL.n261 VTAIL.n196 1.16414
R944 VTAIL.n270 VTAIL.n269 1.16414
R945 VTAIL.n646 VTAIL.n645 1.16414
R946 VTAIL.n637 VTAIL.n572 1.16414
R947 VTAIL.n600 VTAIL.n593 1.16414
R948 VTAIL.n552 VTAIL.n551 1.16414
R949 VTAIL.n543 VTAIL.n478 1.16414
R950 VTAIL.n506 VTAIL.n499 1.16414
R951 VTAIL.n458 VTAIL.n457 1.16414
R952 VTAIL.n449 VTAIL.n384 1.16414
R953 VTAIL.n412 VTAIL.n405 1.16414
R954 VTAIL.n364 VTAIL.n363 1.16414
R955 VTAIL.n355 VTAIL.n290 1.16414
R956 VTAIL.n318 VTAIL.n311 1.16414
R957 VTAIL VTAIL.n93 0.657828
R958 VTAIL VTAIL.n751 0.541448
R959 VTAIL.n563 VTAIL.n469 0.470328
R960 VTAIL.n187 VTAIL.n93 0.470328
R961 VTAIL.n690 VTAIL.n689 0.388379
R962 VTAIL.n735 VTAIL.n734 0.388379
R963 VTAIL.n736 VTAIL.n664 0.388379
R964 VTAIL.n32 VTAIL.n31 0.388379
R965 VTAIL.n77 VTAIL.n76 0.388379
R966 VTAIL.n78 VTAIL.n6 0.388379
R967 VTAIL.n126 VTAIL.n125 0.388379
R968 VTAIL.n171 VTAIL.n170 0.388379
R969 VTAIL.n172 VTAIL.n100 0.388379
R970 VTAIL.n220 VTAIL.n219 0.388379
R971 VTAIL.n265 VTAIL.n264 0.388379
R972 VTAIL.n266 VTAIL.n194 0.388379
R973 VTAIL.n642 VTAIL.n570 0.388379
R974 VTAIL.n641 VTAIL.n640 0.388379
R975 VTAIL.n597 VTAIL.n596 0.388379
R976 VTAIL.n548 VTAIL.n476 0.388379
R977 VTAIL.n547 VTAIL.n546 0.388379
R978 VTAIL.n503 VTAIL.n502 0.388379
R979 VTAIL.n454 VTAIL.n382 0.388379
R980 VTAIL.n453 VTAIL.n452 0.388379
R981 VTAIL.n409 VTAIL.n408 0.388379
R982 VTAIL.n360 VTAIL.n288 0.388379
R983 VTAIL.n359 VTAIL.n358 0.388379
R984 VTAIL.n315 VTAIL.n314 0.388379
R985 VTAIL.n692 VTAIL.n691 0.155672
R986 VTAIL.n692 VTAIL.n683 0.155672
R987 VTAIL.n699 VTAIL.n683 0.155672
R988 VTAIL.n700 VTAIL.n699 0.155672
R989 VTAIL.n700 VTAIL.n679 0.155672
R990 VTAIL.n707 VTAIL.n679 0.155672
R991 VTAIL.n708 VTAIL.n707 0.155672
R992 VTAIL.n708 VTAIL.n675 0.155672
R993 VTAIL.n715 VTAIL.n675 0.155672
R994 VTAIL.n716 VTAIL.n715 0.155672
R995 VTAIL.n716 VTAIL.n671 0.155672
R996 VTAIL.n723 VTAIL.n671 0.155672
R997 VTAIL.n724 VTAIL.n723 0.155672
R998 VTAIL.n724 VTAIL.n667 0.155672
R999 VTAIL.n732 VTAIL.n667 0.155672
R1000 VTAIL.n733 VTAIL.n732 0.155672
R1001 VTAIL.n733 VTAIL.n663 0.155672
R1002 VTAIL.n741 VTAIL.n663 0.155672
R1003 VTAIL.n742 VTAIL.n741 0.155672
R1004 VTAIL.n742 VTAIL.n659 0.155672
R1005 VTAIL.n749 VTAIL.n659 0.155672
R1006 VTAIL.n34 VTAIL.n33 0.155672
R1007 VTAIL.n34 VTAIL.n25 0.155672
R1008 VTAIL.n41 VTAIL.n25 0.155672
R1009 VTAIL.n42 VTAIL.n41 0.155672
R1010 VTAIL.n42 VTAIL.n21 0.155672
R1011 VTAIL.n49 VTAIL.n21 0.155672
R1012 VTAIL.n50 VTAIL.n49 0.155672
R1013 VTAIL.n50 VTAIL.n17 0.155672
R1014 VTAIL.n57 VTAIL.n17 0.155672
R1015 VTAIL.n58 VTAIL.n57 0.155672
R1016 VTAIL.n58 VTAIL.n13 0.155672
R1017 VTAIL.n65 VTAIL.n13 0.155672
R1018 VTAIL.n66 VTAIL.n65 0.155672
R1019 VTAIL.n66 VTAIL.n9 0.155672
R1020 VTAIL.n74 VTAIL.n9 0.155672
R1021 VTAIL.n75 VTAIL.n74 0.155672
R1022 VTAIL.n75 VTAIL.n5 0.155672
R1023 VTAIL.n83 VTAIL.n5 0.155672
R1024 VTAIL.n84 VTAIL.n83 0.155672
R1025 VTAIL.n84 VTAIL.n1 0.155672
R1026 VTAIL.n91 VTAIL.n1 0.155672
R1027 VTAIL.n128 VTAIL.n127 0.155672
R1028 VTAIL.n128 VTAIL.n119 0.155672
R1029 VTAIL.n135 VTAIL.n119 0.155672
R1030 VTAIL.n136 VTAIL.n135 0.155672
R1031 VTAIL.n136 VTAIL.n115 0.155672
R1032 VTAIL.n143 VTAIL.n115 0.155672
R1033 VTAIL.n144 VTAIL.n143 0.155672
R1034 VTAIL.n144 VTAIL.n111 0.155672
R1035 VTAIL.n151 VTAIL.n111 0.155672
R1036 VTAIL.n152 VTAIL.n151 0.155672
R1037 VTAIL.n152 VTAIL.n107 0.155672
R1038 VTAIL.n159 VTAIL.n107 0.155672
R1039 VTAIL.n160 VTAIL.n159 0.155672
R1040 VTAIL.n160 VTAIL.n103 0.155672
R1041 VTAIL.n168 VTAIL.n103 0.155672
R1042 VTAIL.n169 VTAIL.n168 0.155672
R1043 VTAIL.n169 VTAIL.n99 0.155672
R1044 VTAIL.n177 VTAIL.n99 0.155672
R1045 VTAIL.n178 VTAIL.n177 0.155672
R1046 VTAIL.n178 VTAIL.n95 0.155672
R1047 VTAIL.n185 VTAIL.n95 0.155672
R1048 VTAIL.n222 VTAIL.n221 0.155672
R1049 VTAIL.n222 VTAIL.n213 0.155672
R1050 VTAIL.n229 VTAIL.n213 0.155672
R1051 VTAIL.n230 VTAIL.n229 0.155672
R1052 VTAIL.n230 VTAIL.n209 0.155672
R1053 VTAIL.n237 VTAIL.n209 0.155672
R1054 VTAIL.n238 VTAIL.n237 0.155672
R1055 VTAIL.n238 VTAIL.n205 0.155672
R1056 VTAIL.n245 VTAIL.n205 0.155672
R1057 VTAIL.n246 VTAIL.n245 0.155672
R1058 VTAIL.n246 VTAIL.n201 0.155672
R1059 VTAIL.n253 VTAIL.n201 0.155672
R1060 VTAIL.n254 VTAIL.n253 0.155672
R1061 VTAIL.n254 VTAIL.n197 0.155672
R1062 VTAIL.n262 VTAIL.n197 0.155672
R1063 VTAIL.n263 VTAIL.n262 0.155672
R1064 VTAIL.n263 VTAIL.n193 0.155672
R1065 VTAIL.n271 VTAIL.n193 0.155672
R1066 VTAIL.n272 VTAIL.n271 0.155672
R1067 VTAIL.n272 VTAIL.n189 0.155672
R1068 VTAIL.n279 VTAIL.n189 0.155672
R1069 VTAIL.n655 VTAIL.n565 0.155672
R1070 VTAIL.n648 VTAIL.n565 0.155672
R1071 VTAIL.n648 VTAIL.n647 0.155672
R1072 VTAIL.n647 VTAIL.n569 0.155672
R1073 VTAIL.n639 VTAIL.n569 0.155672
R1074 VTAIL.n639 VTAIL.n638 0.155672
R1075 VTAIL.n638 VTAIL.n573 0.155672
R1076 VTAIL.n631 VTAIL.n573 0.155672
R1077 VTAIL.n631 VTAIL.n630 0.155672
R1078 VTAIL.n630 VTAIL.n578 0.155672
R1079 VTAIL.n623 VTAIL.n578 0.155672
R1080 VTAIL.n623 VTAIL.n622 0.155672
R1081 VTAIL.n622 VTAIL.n582 0.155672
R1082 VTAIL.n615 VTAIL.n582 0.155672
R1083 VTAIL.n615 VTAIL.n614 0.155672
R1084 VTAIL.n614 VTAIL.n586 0.155672
R1085 VTAIL.n607 VTAIL.n586 0.155672
R1086 VTAIL.n607 VTAIL.n606 0.155672
R1087 VTAIL.n606 VTAIL.n590 0.155672
R1088 VTAIL.n599 VTAIL.n590 0.155672
R1089 VTAIL.n599 VTAIL.n598 0.155672
R1090 VTAIL.n561 VTAIL.n471 0.155672
R1091 VTAIL.n554 VTAIL.n471 0.155672
R1092 VTAIL.n554 VTAIL.n553 0.155672
R1093 VTAIL.n553 VTAIL.n475 0.155672
R1094 VTAIL.n545 VTAIL.n475 0.155672
R1095 VTAIL.n545 VTAIL.n544 0.155672
R1096 VTAIL.n544 VTAIL.n479 0.155672
R1097 VTAIL.n537 VTAIL.n479 0.155672
R1098 VTAIL.n537 VTAIL.n536 0.155672
R1099 VTAIL.n536 VTAIL.n484 0.155672
R1100 VTAIL.n529 VTAIL.n484 0.155672
R1101 VTAIL.n529 VTAIL.n528 0.155672
R1102 VTAIL.n528 VTAIL.n488 0.155672
R1103 VTAIL.n521 VTAIL.n488 0.155672
R1104 VTAIL.n521 VTAIL.n520 0.155672
R1105 VTAIL.n520 VTAIL.n492 0.155672
R1106 VTAIL.n513 VTAIL.n492 0.155672
R1107 VTAIL.n513 VTAIL.n512 0.155672
R1108 VTAIL.n512 VTAIL.n496 0.155672
R1109 VTAIL.n505 VTAIL.n496 0.155672
R1110 VTAIL.n505 VTAIL.n504 0.155672
R1111 VTAIL.n467 VTAIL.n377 0.155672
R1112 VTAIL.n460 VTAIL.n377 0.155672
R1113 VTAIL.n460 VTAIL.n459 0.155672
R1114 VTAIL.n459 VTAIL.n381 0.155672
R1115 VTAIL.n451 VTAIL.n381 0.155672
R1116 VTAIL.n451 VTAIL.n450 0.155672
R1117 VTAIL.n450 VTAIL.n385 0.155672
R1118 VTAIL.n443 VTAIL.n385 0.155672
R1119 VTAIL.n443 VTAIL.n442 0.155672
R1120 VTAIL.n442 VTAIL.n390 0.155672
R1121 VTAIL.n435 VTAIL.n390 0.155672
R1122 VTAIL.n435 VTAIL.n434 0.155672
R1123 VTAIL.n434 VTAIL.n394 0.155672
R1124 VTAIL.n427 VTAIL.n394 0.155672
R1125 VTAIL.n427 VTAIL.n426 0.155672
R1126 VTAIL.n426 VTAIL.n398 0.155672
R1127 VTAIL.n419 VTAIL.n398 0.155672
R1128 VTAIL.n419 VTAIL.n418 0.155672
R1129 VTAIL.n418 VTAIL.n402 0.155672
R1130 VTAIL.n411 VTAIL.n402 0.155672
R1131 VTAIL.n411 VTAIL.n410 0.155672
R1132 VTAIL.n373 VTAIL.n283 0.155672
R1133 VTAIL.n366 VTAIL.n283 0.155672
R1134 VTAIL.n366 VTAIL.n365 0.155672
R1135 VTAIL.n365 VTAIL.n287 0.155672
R1136 VTAIL.n357 VTAIL.n287 0.155672
R1137 VTAIL.n357 VTAIL.n356 0.155672
R1138 VTAIL.n356 VTAIL.n291 0.155672
R1139 VTAIL.n349 VTAIL.n291 0.155672
R1140 VTAIL.n349 VTAIL.n348 0.155672
R1141 VTAIL.n348 VTAIL.n296 0.155672
R1142 VTAIL.n341 VTAIL.n296 0.155672
R1143 VTAIL.n341 VTAIL.n340 0.155672
R1144 VTAIL.n340 VTAIL.n300 0.155672
R1145 VTAIL.n333 VTAIL.n300 0.155672
R1146 VTAIL.n333 VTAIL.n332 0.155672
R1147 VTAIL.n332 VTAIL.n304 0.155672
R1148 VTAIL.n325 VTAIL.n304 0.155672
R1149 VTAIL.n325 VTAIL.n324 0.155672
R1150 VTAIL.n324 VTAIL.n308 0.155672
R1151 VTAIL.n317 VTAIL.n308 0.155672
R1152 VTAIL.n317 VTAIL.n316 0.155672
R1153 B.n105 B.t15 588.008
R1154 B.n102 B.t11 588.008
R1155 B.n577 B.t4 588.008
R1156 B.n419 B.t8 588.008
R1157 B.n785 B.n784 585
R1158 B.n346 B.n101 585
R1159 B.n345 B.n344 585
R1160 B.n343 B.n342 585
R1161 B.n341 B.n340 585
R1162 B.n339 B.n338 585
R1163 B.n337 B.n336 585
R1164 B.n335 B.n334 585
R1165 B.n333 B.n332 585
R1166 B.n331 B.n330 585
R1167 B.n329 B.n328 585
R1168 B.n327 B.n326 585
R1169 B.n325 B.n324 585
R1170 B.n323 B.n322 585
R1171 B.n321 B.n320 585
R1172 B.n319 B.n318 585
R1173 B.n317 B.n316 585
R1174 B.n315 B.n314 585
R1175 B.n313 B.n312 585
R1176 B.n311 B.n310 585
R1177 B.n309 B.n308 585
R1178 B.n307 B.n306 585
R1179 B.n305 B.n304 585
R1180 B.n303 B.n302 585
R1181 B.n301 B.n300 585
R1182 B.n299 B.n298 585
R1183 B.n297 B.n296 585
R1184 B.n295 B.n294 585
R1185 B.n293 B.n292 585
R1186 B.n291 B.n290 585
R1187 B.n289 B.n288 585
R1188 B.n287 B.n286 585
R1189 B.n285 B.n284 585
R1190 B.n283 B.n282 585
R1191 B.n281 B.n280 585
R1192 B.n279 B.n278 585
R1193 B.n277 B.n276 585
R1194 B.n275 B.n274 585
R1195 B.n273 B.n272 585
R1196 B.n271 B.n270 585
R1197 B.n269 B.n268 585
R1198 B.n267 B.n266 585
R1199 B.n265 B.n264 585
R1200 B.n263 B.n262 585
R1201 B.n261 B.n260 585
R1202 B.n259 B.n258 585
R1203 B.n257 B.n256 585
R1204 B.n255 B.n254 585
R1205 B.n253 B.n252 585
R1206 B.n251 B.n250 585
R1207 B.n249 B.n248 585
R1208 B.n247 B.n246 585
R1209 B.n245 B.n244 585
R1210 B.n243 B.n242 585
R1211 B.n241 B.n240 585
R1212 B.n239 B.n238 585
R1213 B.n237 B.n236 585
R1214 B.n235 B.n234 585
R1215 B.n233 B.n232 585
R1216 B.n231 B.n230 585
R1217 B.n229 B.n228 585
R1218 B.n227 B.n226 585
R1219 B.n225 B.n224 585
R1220 B.n223 B.n222 585
R1221 B.n221 B.n220 585
R1222 B.n219 B.n218 585
R1223 B.n217 B.n216 585
R1224 B.n215 B.n214 585
R1225 B.n213 B.n212 585
R1226 B.n211 B.n210 585
R1227 B.n209 B.n208 585
R1228 B.n207 B.n206 585
R1229 B.n205 B.n204 585
R1230 B.n203 B.n202 585
R1231 B.n201 B.n200 585
R1232 B.n199 B.n198 585
R1233 B.n197 B.n196 585
R1234 B.n195 B.n194 585
R1235 B.n193 B.n192 585
R1236 B.n191 B.n190 585
R1237 B.n189 B.n188 585
R1238 B.n187 B.n186 585
R1239 B.n185 B.n184 585
R1240 B.n183 B.n182 585
R1241 B.n181 B.n180 585
R1242 B.n179 B.n178 585
R1243 B.n177 B.n176 585
R1244 B.n175 B.n174 585
R1245 B.n173 B.n172 585
R1246 B.n171 B.n170 585
R1247 B.n169 B.n168 585
R1248 B.n167 B.n166 585
R1249 B.n165 B.n164 585
R1250 B.n163 B.n162 585
R1251 B.n161 B.n160 585
R1252 B.n159 B.n158 585
R1253 B.n157 B.n156 585
R1254 B.n155 B.n154 585
R1255 B.n153 B.n152 585
R1256 B.n151 B.n150 585
R1257 B.n149 B.n148 585
R1258 B.n147 B.n146 585
R1259 B.n145 B.n144 585
R1260 B.n143 B.n142 585
R1261 B.n141 B.n140 585
R1262 B.n139 B.n138 585
R1263 B.n137 B.n136 585
R1264 B.n135 B.n134 585
R1265 B.n133 B.n132 585
R1266 B.n131 B.n130 585
R1267 B.n129 B.n128 585
R1268 B.n127 B.n126 585
R1269 B.n125 B.n124 585
R1270 B.n123 B.n122 585
R1271 B.n121 B.n120 585
R1272 B.n119 B.n118 585
R1273 B.n117 B.n116 585
R1274 B.n115 B.n114 585
R1275 B.n113 B.n112 585
R1276 B.n111 B.n110 585
R1277 B.n109 B.n108 585
R1278 B.n39 B.n38 585
R1279 B.n783 B.n40 585
R1280 B.n788 B.n40 585
R1281 B.n782 B.n781 585
R1282 B.n781 B.n36 585
R1283 B.n780 B.n35 585
R1284 B.n794 B.n35 585
R1285 B.n779 B.n34 585
R1286 B.n795 B.n34 585
R1287 B.n778 B.n33 585
R1288 B.n796 B.n33 585
R1289 B.n777 B.n776 585
R1290 B.n776 B.n32 585
R1291 B.n775 B.n28 585
R1292 B.n802 B.n28 585
R1293 B.n774 B.n27 585
R1294 B.n803 B.n27 585
R1295 B.n773 B.n26 585
R1296 B.n804 B.n26 585
R1297 B.n772 B.n771 585
R1298 B.n771 B.n22 585
R1299 B.n770 B.n21 585
R1300 B.n810 B.n21 585
R1301 B.n769 B.n20 585
R1302 B.n811 B.n20 585
R1303 B.n768 B.n19 585
R1304 B.n812 B.n19 585
R1305 B.n767 B.n766 585
R1306 B.n766 B.n15 585
R1307 B.n765 B.n14 585
R1308 B.n818 B.n14 585
R1309 B.n764 B.n13 585
R1310 B.n819 B.n13 585
R1311 B.n763 B.n12 585
R1312 B.n820 B.n12 585
R1313 B.n762 B.n761 585
R1314 B.n761 B.n760 585
R1315 B.n759 B.n758 585
R1316 B.n759 B.n8 585
R1317 B.n757 B.n7 585
R1318 B.n827 B.n7 585
R1319 B.n756 B.n6 585
R1320 B.n828 B.n6 585
R1321 B.n755 B.n5 585
R1322 B.n829 B.n5 585
R1323 B.n754 B.n753 585
R1324 B.n753 B.n4 585
R1325 B.n752 B.n347 585
R1326 B.n752 B.n751 585
R1327 B.n742 B.n348 585
R1328 B.n349 B.n348 585
R1329 B.n744 B.n743 585
R1330 B.n745 B.n744 585
R1331 B.n741 B.n354 585
R1332 B.n354 B.n353 585
R1333 B.n740 B.n739 585
R1334 B.n739 B.n738 585
R1335 B.n356 B.n355 585
R1336 B.n357 B.n356 585
R1337 B.n731 B.n730 585
R1338 B.n732 B.n731 585
R1339 B.n729 B.n362 585
R1340 B.n362 B.n361 585
R1341 B.n728 B.n727 585
R1342 B.n727 B.n726 585
R1343 B.n364 B.n363 585
R1344 B.n365 B.n364 585
R1345 B.n719 B.n718 585
R1346 B.n720 B.n719 585
R1347 B.n717 B.n370 585
R1348 B.n370 B.n369 585
R1349 B.n716 B.n715 585
R1350 B.n715 B.n714 585
R1351 B.n372 B.n371 585
R1352 B.n707 B.n372 585
R1353 B.n706 B.n705 585
R1354 B.n708 B.n706 585
R1355 B.n704 B.n377 585
R1356 B.n377 B.n376 585
R1357 B.n703 B.n702 585
R1358 B.n702 B.n701 585
R1359 B.n379 B.n378 585
R1360 B.n380 B.n379 585
R1361 B.n694 B.n693 585
R1362 B.n695 B.n694 585
R1363 B.n383 B.n382 585
R1364 B.n450 B.n448 585
R1365 B.n451 B.n447 585
R1366 B.n451 B.n384 585
R1367 B.n454 B.n453 585
R1368 B.n455 B.n446 585
R1369 B.n457 B.n456 585
R1370 B.n459 B.n445 585
R1371 B.n462 B.n461 585
R1372 B.n463 B.n444 585
R1373 B.n465 B.n464 585
R1374 B.n467 B.n443 585
R1375 B.n470 B.n469 585
R1376 B.n471 B.n442 585
R1377 B.n473 B.n472 585
R1378 B.n475 B.n441 585
R1379 B.n478 B.n477 585
R1380 B.n479 B.n440 585
R1381 B.n481 B.n480 585
R1382 B.n483 B.n439 585
R1383 B.n486 B.n485 585
R1384 B.n487 B.n438 585
R1385 B.n489 B.n488 585
R1386 B.n491 B.n437 585
R1387 B.n494 B.n493 585
R1388 B.n495 B.n436 585
R1389 B.n497 B.n496 585
R1390 B.n499 B.n435 585
R1391 B.n502 B.n501 585
R1392 B.n503 B.n434 585
R1393 B.n505 B.n504 585
R1394 B.n507 B.n433 585
R1395 B.n510 B.n509 585
R1396 B.n511 B.n432 585
R1397 B.n513 B.n512 585
R1398 B.n515 B.n431 585
R1399 B.n518 B.n517 585
R1400 B.n519 B.n430 585
R1401 B.n521 B.n520 585
R1402 B.n523 B.n429 585
R1403 B.n526 B.n525 585
R1404 B.n527 B.n428 585
R1405 B.n529 B.n528 585
R1406 B.n531 B.n427 585
R1407 B.n534 B.n533 585
R1408 B.n535 B.n426 585
R1409 B.n537 B.n536 585
R1410 B.n539 B.n425 585
R1411 B.n542 B.n541 585
R1412 B.n543 B.n424 585
R1413 B.n545 B.n544 585
R1414 B.n547 B.n423 585
R1415 B.n550 B.n549 585
R1416 B.n551 B.n422 585
R1417 B.n553 B.n552 585
R1418 B.n555 B.n421 585
R1419 B.n558 B.n557 585
R1420 B.n560 B.n418 585
R1421 B.n562 B.n561 585
R1422 B.n564 B.n417 585
R1423 B.n567 B.n566 585
R1424 B.n568 B.n416 585
R1425 B.n570 B.n569 585
R1426 B.n572 B.n415 585
R1427 B.n575 B.n574 585
R1428 B.n576 B.n414 585
R1429 B.n581 B.n580 585
R1430 B.n583 B.n413 585
R1431 B.n586 B.n585 585
R1432 B.n587 B.n412 585
R1433 B.n589 B.n588 585
R1434 B.n591 B.n411 585
R1435 B.n594 B.n593 585
R1436 B.n595 B.n410 585
R1437 B.n597 B.n596 585
R1438 B.n599 B.n409 585
R1439 B.n602 B.n601 585
R1440 B.n603 B.n408 585
R1441 B.n605 B.n604 585
R1442 B.n607 B.n407 585
R1443 B.n610 B.n609 585
R1444 B.n611 B.n406 585
R1445 B.n613 B.n612 585
R1446 B.n615 B.n405 585
R1447 B.n618 B.n617 585
R1448 B.n619 B.n404 585
R1449 B.n621 B.n620 585
R1450 B.n623 B.n403 585
R1451 B.n626 B.n625 585
R1452 B.n627 B.n402 585
R1453 B.n629 B.n628 585
R1454 B.n631 B.n401 585
R1455 B.n634 B.n633 585
R1456 B.n635 B.n400 585
R1457 B.n637 B.n636 585
R1458 B.n639 B.n399 585
R1459 B.n642 B.n641 585
R1460 B.n643 B.n398 585
R1461 B.n645 B.n644 585
R1462 B.n647 B.n397 585
R1463 B.n650 B.n649 585
R1464 B.n651 B.n396 585
R1465 B.n653 B.n652 585
R1466 B.n655 B.n395 585
R1467 B.n658 B.n657 585
R1468 B.n659 B.n394 585
R1469 B.n661 B.n660 585
R1470 B.n663 B.n393 585
R1471 B.n666 B.n665 585
R1472 B.n667 B.n392 585
R1473 B.n669 B.n668 585
R1474 B.n671 B.n391 585
R1475 B.n674 B.n673 585
R1476 B.n675 B.n390 585
R1477 B.n677 B.n676 585
R1478 B.n679 B.n389 585
R1479 B.n682 B.n681 585
R1480 B.n683 B.n388 585
R1481 B.n685 B.n684 585
R1482 B.n687 B.n387 585
R1483 B.n688 B.n386 585
R1484 B.n691 B.n690 585
R1485 B.n692 B.n385 585
R1486 B.n385 B.n384 585
R1487 B.n697 B.n696 585
R1488 B.n696 B.n695 585
R1489 B.n698 B.n381 585
R1490 B.n381 B.n380 585
R1491 B.n700 B.n699 585
R1492 B.n701 B.n700 585
R1493 B.n375 B.n374 585
R1494 B.n376 B.n375 585
R1495 B.n710 B.n709 585
R1496 B.n709 B.n708 585
R1497 B.n711 B.n373 585
R1498 B.n707 B.n373 585
R1499 B.n713 B.n712 585
R1500 B.n714 B.n713 585
R1501 B.n368 B.n367 585
R1502 B.n369 B.n368 585
R1503 B.n722 B.n721 585
R1504 B.n721 B.n720 585
R1505 B.n723 B.n366 585
R1506 B.n366 B.n365 585
R1507 B.n725 B.n724 585
R1508 B.n726 B.n725 585
R1509 B.n360 B.n359 585
R1510 B.n361 B.n360 585
R1511 B.n734 B.n733 585
R1512 B.n733 B.n732 585
R1513 B.n735 B.n358 585
R1514 B.n358 B.n357 585
R1515 B.n737 B.n736 585
R1516 B.n738 B.n737 585
R1517 B.n352 B.n351 585
R1518 B.n353 B.n352 585
R1519 B.n747 B.n746 585
R1520 B.n746 B.n745 585
R1521 B.n748 B.n350 585
R1522 B.n350 B.n349 585
R1523 B.n750 B.n749 585
R1524 B.n751 B.n750 585
R1525 B.n3 B.n0 585
R1526 B.n4 B.n3 585
R1527 B.n826 B.n1 585
R1528 B.n827 B.n826 585
R1529 B.n825 B.n824 585
R1530 B.n825 B.n8 585
R1531 B.n823 B.n9 585
R1532 B.n760 B.n9 585
R1533 B.n822 B.n821 585
R1534 B.n821 B.n820 585
R1535 B.n11 B.n10 585
R1536 B.n819 B.n11 585
R1537 B.n817 B.n816 585
R1538 B.n818 B.n817 585
R1539 B.n815 B.n16 585
R1540 B.n16 B.n15 585
R1541 B.n814 B.n813 585
R1542 B.n813 B.n812 585
R1543 B.n18 B.n17 585
R1544 B.n811 B.n18 585
R1545 B.n809 B.n808 585
R1546 B.n810 B.n809 585
R1547 B.n807 B.n23 585
R1548 B.n23 B.n22 585
R1549 B.n806 B.n805 585
R1550 B.n805 B.n804 585
R1551 B.n25 B.n24 585
R1552 B.n803 B.n25 585
R1553 B.n801 B.n800 585
R1554 B.n802 B.n801 585
R1555 B.n799 B.n29 585
R1556 B.n32 B.n29 585
R1557 B.n798 B.n797 585
R1558 B.n797 B.n796 585
R1559 B.n31 B.n30 585
R1560 B.n795 B.n31 585
R1561 B.n793 B.n792 585
R1562 B.n794 B.n793 585
R1563 B.n791 B.n37 585
R1564 B.n37 B.n36 585
R1565 B.n790 B.n789 585
R1566 B.n789 B.n788 585
R1567 B.n830 B.n829 585
R1568 B.n828 B.n2 585
R1569 B.n789 B.n39 458.866
R1570 B.n785 B.n40 458.866
R1571 B.n694 B.n385 458.866
R1572 B.n696 B.n383 458.866
R1573 B.n102 B.t13 394.055
R1574 B.n577 B.t7 394.055
R1575 B.n105 B.t16 394.055
R1576 B.n419 B.t10 394.055
R1577 B.n103 B.t14 367.099
R1578 B.n578 B.t6 367.099
R1579 B.n106 B.t17 367.099
R1580 B.n420 B.t9 367.099
R1581 B.n787 B.n786 256.663
R1582 B.n787 B.n100 256.663
R1583 B.n787 B.n99 256.663
R1584 B.n787 B.n98 256.663
R1585 B.n787 B.n97 256.663
R1586 B.n787 B.n96 256.663
R1587 B.n787 B.n95 256.663
R1588 B.n787 B.n94 256.663
R1589 B.n787 B.n93 256.663
R1590 B.n787 B.n92 256.663
R1591 B.n787 B.n91 256.663
R1592 B.n787 B.n90 256.663
R1593 B.n787 B.n89 256.663
R1594 B.n787 B.n88 256.663
R1595 B.n787 B.n87 256.663
R1596 B.n787 B.n86 256.663
R1597 B.n787 B.n85 256.663
R1598 B.n787 B.n84 256.663
R1599 B.n787 B.n83 256.663
R1600 B.n787 B.n82 256.663
R1601 B.n787 B.n81 256.663
R1602 B.n787 B.n80 256.663
R1603 B.n787 B.n79 256.663
R1604 B.n787 B.n78 256.663
R1605 B.n787 B.n77 256.663
R1606 B.n787 B.n76 256.663
R1607 B.n787 B.n75 256.663
R1608 B.n787 B.n74 256.663
R1609 B.n787 B.n73 256.663
R1610 B.n787 B.n72 256.663
R1611 B.n787 B.n71 256.663
R1612 B.n787 B.n70 256.663
R1613 B.n787 B.n69 256.663
R1614 B.n787 B.n68 256.663
R1615 B.n787 B.n67 256.663
R1616 B.n787 B.n66 256.663
R1617 B.n787 B.n65 256.663
R1618 B.n787 B.n64 256.663
R1619 B.n787 B.n63 256.663
R1620 B.n787 B.n62 256.663
R1621 B.n787 B.n61 256.663
R1622 B.n787 B.n60 256.663
R1623 B.n787 B.n59 256.663
R1624 B.n787 B.n58 256.663
R1625 B.n787 B.n57 256.663
R1626 B.n787 B.n56 256.663
R1627 B.n787 B.n55 256.663
R1628 B.n787 B.n54 256.663
R1629 B.n787 B.n53 256.663
R1630 B.n787 B.n52 256.663
R1631 B.n787 B.n51 256.663
R1632 B.n787 B.n50 256.663
R1633 B.n787 B.n49 256.663
R1634 B.n787 B.n48 256.663
R1635 B.n787 B.n47 256.663
R1636 B.n787 B.n46 256.663
R1637 B.n787 B.n45 256.663
R1638 B.n787 B.n44 256.663
R1639 B.n787 B.n43 256.663
R1640 B.n787 B.n42 256.663
R1641 B.n787 B.n41 256.663
R1642 B.n449 B.n384 256.663
R1643 B.n452 B.n384 256.663
R1644 B.n458 B.n384 256.663
R1645 B.n460 B.n384 256.663
R1646 B.n466 B.n384 256.663
R1647 B.n468 B.n384 256.663
R1648 B.n474 B.n384 256.663
R1649 B.n476 B.n384 256.663
R1650 B.n482 B.n384 256.663
R1651 B.n484 B.n384 256.663
R1652 B.n490 B.n384 256.663
R1653 B.n492 B.n384 256.663
R1654 B.n498 B.n384 256.663
R1655 B.n500 B.n384 256.663
R1656 B.n506 B.n384 256.663
R1657 B.n508 B.n384 256.663
R1658 B.n514 B.n384 256.663
R1659 B.n516 B.n384 256.663
R1660 B.n522 B.n384 256.663
R1661 B.n524 B.n384 256.663
R1662 B.n530 B.n384 256.663
R1663 B.n532 B.n384 256.663
R1664 B.n538 B.n384 256.663
R1665 B.n540 B.n384 256.663
R1666 B.n546 B.n384 256.663
R1667 B.n548 B.n384 256.663
R1668 B.n554 B.n384 256.663
R1669 B.n556 B.n384 256.663
R1670 B.n563 B.n384 256.663
R1671 B.n565 B.n384 256.663
R1672 B.n571 B.n384 256.663
R1673 B.n573 B.n384 256.663
R1674 B.n582 B.n384 256.663
R1675 B.n584 B.n384 256.663
R1676 B.n590 B.n384 256.663
R1677 B.n592 B.n384 256.663
R1678 B.n598 B.n384 256.663
R1679 B.n600 B.n384 256.663
R1680 B.n606 B.n384 256.663
R1681 B.n608 B.n384 256.663
R1682 B.n614 B.n384 256.663
R1683 B.n616 B.n384 256.663
R1684 B.n622 B.n384 256.663
R1685 B.n624 B.n384 256.663
R1686 B.n630 B.n384 256.663
R1687 B.n632 B.n384 256.663
R1688 B.n638 B.n384 256.663
R1689 B.n640 B.n384 256.663
R1690 B.n646 B.n384 256.663
R1691 B.n648 B.n384 256.663
R1692 B.n654 B.n384 256.663
R1693 B.n656 B.n384 256.663
R1694 B.n662 B.n384 256.663
R1695 B.n664 B.n384 256.663
R1696 B.n670 B.n384 256.663
R1697 B.n672 B.n384 256.663
R1698 B.n678 B.n384 256.663
R1699 B.n680 B.n384 256.663
R1700 B.n686 B.n384 256.663
R1701 B.n689 B.n384 256.663
R1702 B.n832 B.n831 256.663
R1703 B.n110 B.n109 163.367
R1704 B.n114 B.n113 163.367
R1705 B.n118 B.n117 163.367
R1706 B.n122 B.n121 163.367
R1707 B.n126 B.n125 163.367
R1708 B.n130 B.n129 163.367
R1709 B.n134 B.n133 163.367
R1710 B.n138 B.n137 163.367
R1711 B.n142 B.n141 163.367
R1712 B.n146 B.n145 163.367
R1713 B.n150 B.n149 163.367
R1714 B.n154 B.n153 163.367
R1715 B.n158 B.n157 163.367
R1716 B.n162 B.n161 163.367
R1717 B.n166 B.n165 163.367
R1718 B.n170 B.n169 163.367
R1719 B.n174 B.n173 163.367
R1720 B.n178 B.n177 163.367
R1721 B.n182 B.n181 163.367
R1722 B.n186 B.n185 163.367
R1723 B.n190 B.n189 163.367
R1724 B.n194 B.n193 163.367
R1725 B.n198 B.n197 163.367
R1726 B.n202 B.n201 163.367
R1727 B.n206 B.n205 163.367
R1728 B.n210 B.n209 163.367
R1729 B.n214 B.n213 163.367
R1730 B.n218 B.n217 163.367
R1731 B.n222 B.n221 163.367
R1732 B.n226 B.n225 163.367
R1733 B.n230 B.n229 163.367
R1734 B.n234 B.n233 163.367
R1735 B.n238 B.n237 163.367
R1736 B.n242 B.n241 163.367
R1737 B.n246 B.n245 163.367
R1738 B.n250 B.n249 163.367
R1739 B.n254 B.n253 163.367
R1740 B.n258 B.n257 163.367
R1741 B.n262 B.n261 163.367
R1742 B.n266 B.n265 163.367
R1743 B.n270 B.n269 163.367
R1744 B.n274 B.n273 163.367
R1745 B.n278 B.n277 163.367
R1746 B.n282 B.n281 163.367
R1747 B.n286 B.n285 163.367
R1748 B.n290 B.n289 163.367
R1749 B.n294 B.n293 163.367
R1750 B.n298 B.n297 163.367
R1751 B.n302 B.n301 163.367
R1752 B.n306 B.n305 163.367
R1753 B.n310 B.n309 163.367
R1754 B.n314 B.n313 163.367
R1755 B.n318 B.n317 163.367
R1756 B.n322 B.n321 163.367
R1757 B.n326 B.n325 163.367
R1758 B.n330 B.n329 163.367
R1759 B.n334 B.n333 163.367
R1760 B.n338 B.n337 163.367
R1761 B.n342 B.n341 163.367
R1762 B.n344 B.n101 163.367
R1763 B.n694 B.n379 163.367
R1764 B.n702 B.n379 163.367
R1765 B.n702 B.n377 163.367
R1766 B.n706 B.n377 163.367
R1767 B.n706 B.n372 163.367
R1768 B.n715 B.n372 163.367
R1769 B.n715 B.n370 163.367
R1770 B.n719 B.n370 163.367
R1771 B.n719 B.n364 163.367
R1772 B.n727 B.n364 163.367
R1773 B.n727 B.n362 163.367
R1774 B.n731 B.n362 163.367
R1775 B.n731 B.n356 163.367
R1776 B.n739 B.n356 163.367
R1777 B.n739 B.n354 163.367
R1778 B.n744 B.n354 163.367
R1779 B.n744 B.n348 163.367
R1780 B.n752 B.n348 163.367
R1781 B.n753 B.n752 163.367
R1782 B.n753 B.n5 163.367
R1783 B.n6 B.n5 163.367
R1784 B.n7 B.n6 163.367
R1785 B.n759 B.n7 163.367
R1786 B.n761 B.n759 163.367
R1787 B.n761 B.n12 163.367
R1788 B.n13 B.n12 163.367
R1789 B.n14 B.n13 163.367
R1790 B.n766 B.n14 163.367
R1791 B.n766 B.n19 163.367
R1792 B.n20 B.n19 163.367
R1793 B.n21 B.n20 163.367
R1794 B.n771 B.n21 163.367
R1795 B.n771 B.n26 163.367
R1796 B.n27 B.n26 163.367
R1797 B.n28 B.n27 163.367
R1798 B.n776 B.n28 163.367
R1799 B.n776 B.n33 163.367
R1800 B.n34 B.n33 163.367
R1801 B.n35 B.n34 163.367
R1802 B.n781 B.n35 163.367
R1803 B.n781 B.n40 163.367
R1804 B.n451 B.n450 163.367
R1805 B.n453 B.n451 163.367
R1806 B.n457 B.n446 163.367
R1807 B.n461 B.n459 163.367
R1808 B.n465 B.n444 163.367
R1809 B.n469 B.n467 163.367
R1810 B.n473 B.n442 163.367
R1811 B.n477 B.n475 163.367
R1812 B.n481 B.n440 163.367
R1813 B.n485 B.n483 163.367
R1814 B.n489 B.n438 163.367
R1815 B.n493 B.n491 163.367
R1816 B.n497 B.n436 163.367
R1817 B.n501 B.n499 163.367
R1818 B.n505 B.n434 163.367
R1819 B.n509 B.n507 163.367
R1820 B.n513 B.n432 163.367
R1821 B.n517 B.n515 163.367
R1822 B.n521 B.n430 163.367
R1823 B.n525 B.n523 163.367
R1824 B.n529 B.n428 163.367
R1825 B.n533 B.n531 163.367
R1826 B.n537 B.n426 163.367
R1827 B.n541 B.n539 163.367
R1828 B.n545 B.n424 163.367
R1829 B.n549 B.n547 163.367
R1830 B.n553 B.n422 163.367
R1831 B.n557 B.n555 163.367
R1832 B.n562 B.n418 163.367
R1833 B.n566 B.n564 163.367
R1834 B.n570 B.n416 163.367
R1835 B.n574 B.n572 163.367
R1836 B.n581 B.n414 163.367
R1837 B.n585 B.n583 163.367
R1838 B.n589 B.n412 163.367
R1839 B.n593 B.n591 163.367
R1840 B.n597 B.n410 163.367
R1841 B.n601 B.n599 163.367
R1842 B.n605 B.n408 163.367
R1843 B.n609 B.n607 163.367
R1844 B.n613 B.n406 163.367
R1845 B.n617 B.n615 163.367
R1846 B.n621 B.n404 163.367
R1847 B.n625 B.n623 163.367
R1848 B.n629 B.n402 163.367
R1849 B.n633 B.n631 163.367
R1850 B.n637 B.n400 163.367
R1851 B.n641 B.n639 163.367
R1852 B.n645 B.n398 163.367
R1853 B.n649 B.n647 163.367
R1854 B.n653 B.n396 163.367
R1855 B.n657 B.n655 163.367
R1856 B.n661 B.n394 163.367
R1857 B.n665 B.n663 163.367
R1858 B.n669 B.n392 163.367
R1859 B.n673 B.n671 163.367
R1860 B.n677 B.n390 163.367
R1861 B.n681 B.n679 163.367
R1862 B.n685 B.n388 163.367
R1863 B.n688 B.n687 163.367
R1864 B.n690 B.n385 163.367
R1865 B.n696 B.n381 163.367
R1866 B.n700 B.n381 163.367
R1867 B.n700 B.n375 163.367
R1868 B.n709 B.n375 163.367
R1869 B.n709 B.n373 163.367
R1870 B.n713 B.n373 163.367
R1871 B.n713 B.n368 163.367
R1872 B.n721 B.n368 163.367
R1873 B.n721 B.n366 163.367
R1874 B.n725 B.n366 163.367
R1875 B.n725 B.n360 163.367
R1876 B.n733 B.n360 163.367
R1877 B.n733 B.n358 163.367
R1878 B.n737 B.n358 163.367
R1879 B.n737 B.n352 163.367
R1880 B.n746 B.n352 163.367
R1881 B.n746 B.n350 163.367
R1882 B.n750 B.n350 163.367
R1883 B.n750 B.n3 163.367
R1884 B.n830 B.n3 163.367
R1885 B.n826 B.n2 163.367
R1886 B.n826 B.n825 163.367
R1887 B.n825 B.n9 163.367
R1888 B.n821 B.n9 163.367
R1889 B.n821 B.n11 163.367
R1890 B.n817 B.n11 163.367
R1891 B.n817 B.n16 163.367
R1892 B.n813 B.n16 163.367
R1893 B.n813 B.n18 163.367
R1894 B.n809 B.n18 163.367
R1895 B.n809 B.n23 163.367
R1896 B.n805 B.n23 163.367
R1897 B.n805 B.n25 163.367
R1898 B.n801 B.n25 163.367
R1899 B.n801 B.n29 163.367
R1900 B.n797 B.n29 163.367
R1901 B.n797 B.n31 163.367
R1902 B.n793 B.n31 163.367
R1903 B.n793 B.n37 163.367
R1904 B.n789 B.n37 163.367
R1905 B.n41 B.n39 71.676
R1906 B.n110 B.n42 71.676
R1907 B.n114 B.n43 71.676
R1908 B.n118 B.n44 71.676
R1909 B.n122 B.n45 71.676
R1910 B.n126 B.n46 71.676
R1911 B.n130 B.n47 71.676
R1912 B.n134 B.n48 71.676
R1913 B.n138 B.n49 71.676
R1914 B.n142 B.n50 71.676
R1915 B.n146 B.n51 71.676
R1916 B.n150 B.n52 71.676
R1917 B.n154 B.n53 71.676
R1918 B.n158 B.n54 71.676
R1919 B.n162 B.n55 71.676
R1920 B.n166 B.n56 71.676
R1921 B.n170 B.n57 71.676
R1922 B.n174 B.n58 71.676
R1923 B.n178 B.n59 71.676
R1924 B.n182 B.n60 71.676
R1925 B.n186 B.n61 71.676
R1926 B.n190 B.n62 71.676
R1927 B.n194 B.n63 71.676
R1928 B.n198 B.n64 71.676
R1929 B.n202 B.n65 71.676
R1930 B.n206 B.n66 71.676
R1931 B.n210 B.n67 71.676
R1932 B.n214 B.n68 71.676
R1933 B.n218 B.n69 71.676
R1934 B.n222 B.n70 71.676
R1935 B.n226 B.n71 71.676
R1936 B.n230 B.n72 71.676
R1937 B.n234 B.n73 71.676
R1938 B.n238 B.n74 71.676
R1939 B.n242 B.n75 71.676
R1940 B.n246 B.n76 71.676
R1941 B.n250 B.n77 71.676
R1942 B.n254 B.n78 71.676
R1943 B.n258 B.n79 71.676
R1944 B.n262 B.n80 71.676
R1945 B.n266 B.n81 71.676
R1946 B.n270 B.n82 71.676
R1947 B.n274 B.n83 71.676
R1948 B.n278 B.n84 71.676
R1949 B.n282 B.n85 71.676
R1950 B.n286 B.n86 71.676
R1951 B.n290 B.n87 71.676
R1952 B.n294 B.n88 71.676
R1953 B.n298 B.n89 71.676
R1954 B.n302 B.n90 71.676
R1955 B.n306 B.n91 71.676
R1956 B.n310 B.n92 71.676
R1957 B.n314 B.n93 71.676
R1958 B.n318 B.n94 71.676
R1959 B.n322 B.n95 71.676
R1960 B.n326 B.n96 71.676
R1961 B.n330 B.n97 71.676
R1962 B.n334 B.n98 71.676
R1963 B.n338 B.n99 71.676
R1964 B.n342 B.n100 71.676
R1965 B.n786 B.n101 71.676
R1966 B.n786 B.n785 71.676
R1967 B.n344 B.n100 71.676
R1968 B.n341 B.n99 71.676
R1969 B.n337 B.n98 71.676
R1970 B.n333 B.n97 71.676
R1971 B.n329 B.n96 71.676
R1972 B.n325 B.n95 71.676
R1973 B.n321 B.n94 71.676
R1974 B.n317 B.n93 71.676
R1975 B.n313 B.n92 71.676
R1976 B.n309 B.n91 71.676
R1977 B.n305 B.n90 71.676
R1978 B.n301 B.n89 71.676
R1979 B.n297 B.n88 71.676
R1980 B.n293 B.n87 71.676
R1981 B.n289 B.n86 71.676
R1982 B.n285 B.n85 71.676
R1983 B.n281 B.n84 71.676
R1984 B.n277 B.n83 71.676
R1985 B.n273 B.n82 71.676
R1986 B.n269 B.n81 71.676
R1987 B.n265 B.n80 71.676
R1988 B.n261 B.n79 71.676
R1989 B.n257 B.n78 71.676
R1990 B.n253 B.n77 71.676
R1991 B.n249 B.n76 71.676
R1992 B.n245 B.n75 71.676
R1993 B.n241 B.n74 71.676
R1994 B.n237 B.n73 71.676
R1995 B.n233 B.n72 71.676
R1996 B.n229 B.n71 71.676
R1997 B.n225 B.n70 71.676
R1998 B.n221 B.n69 71.676
R1999 B.n217 B.n68 71.676
R2000 B.n213 B.n67 71.676
R2001 B.n209 B.n66 71.676
R2002 B.n205 B.n65 71.676
R2003 B.n201 B.n64 71.676
R2004 B.n197 B.n63 71.676
R2005 B.n193 B.n62 71.676
R2006 B.n189 B.n61 71.676
R2007 B.n185 B.n60 71.676
R2008 B.n181 B.n59 71.676
R2009 B.n177 B.n58 71.676
R2010 B.n173 B.n57 71.676
R2011 B.n169 B.n56 71.676
R2012 B.n165 B.n55 71.676
R2013 B.n161 B.n54 71.676
R2014 B.n157 B.n53 71.676
R2015 B.n153 B.n52 71.676
R2016 B.n149 B.n51 71.676
R2017 B.n145 B.n50 71.676
R2018 B.n141 B.n49 71.676
R2019 B.n137 B.n48 71.676
R2020 B.n133 B.n47 71.676
R2021 B.n129 B.n46 71.676
R2022 B.n125 B.n45 71.676
R2023 B.n121 B.n44 71.676
R2024 B.n117 B.n43 71.676
R2025 B.n113 B.n42 71.676
R2026 B.n109 B.n41 71.676
R2027 B.n449 B.n383 71.676
R2028 B.n453 B.n452 71.676
R2029 B.n458 B.n457 71.676
R2030 B.n461 B.n460 71.676
R2031 B.n466 B.n465 71.676
R2032 B.n469 B.n468 71.676
R2033 B.n474 B.n473 71.676
R2034 B.n477 B.n476 71.676
R2035 B.n482 B.n481 71.676
R2036 B.n485 B.n484 71.676
R2037 B.n490 B.n489 71.676
R2038 B.n493 B.n492 71.676
R2039 B.n498 B.n497 71.676
R2040 B.n501 B.n500 71.676
R2041 B.n506 B.n505 71.676
R2042 B.n509 B.n508 71.676
R2043 B.n514 B.n513 71.676
R2044 B.n517 B.n516 71.676
R2045 B.n522 B.n521 71.676
R2046 B.n525 B.n524 71.676
R2047 B.n530 B.n529 71.676
R2048 B.n533 B.n532 71.676
R2049 B.n538 B.n537 71.676
R2050 B.n541 B.n540 71.676
R2051 B.n546 B.n545 71.676
R2052 B.n549 B.n548 71.676
R2053 B.n554 B.n553 71.676
R2054 B.n557 B.n556 71.676
R2055 B.n563 B.n562 71.676
R2056 B.n566 B.n565 71.676
R2057 B.n571 B.n570 71.676
R2058 B.n574 B.n573 71.676
R2059 B.n582 B.n581 71.676
R2060 B.n585 B.n584 71.676
R2061 B.n590 B.n589 71.676
R2062 B.n593 B.n592 71.676
R2063 B.n598 B.n597 71.676
R2064 B.n601 B.n600 71.676
R2065 B.n606 B.n605 71.676
R2066 B.n609 B.n608 71.676
R2067 B.n614 B.n613 71.676
R2068 B.n617 B.n616 71.676
R2069 B.n622 B.n621 71.676
R2070 B.n625 B.n624 71.676
R2071 B.n630 B.n629 71.676
R2072 B.n633 B.n632 71.676
R2073 B.n638 B.n637 71.676
R2074 B.n641 B.n640 71.676
R2075 B.n646 B.n645 71.676
R2076 B.n649 B.n648 71.676
R2077 B.n654 B.n653 71.676
R2078 B.n657 B.n656 71.676
R2079 B.n662 B.n661 71.676
R2080 B.n665 B.n664 71.676
R2081 B.n670 B.n669 71.676
R2082 B.n673 B.n672 71.676
R2083 B.n678 B.n677 71.676
R2084 B.n681 B.n680 71.676
R2085 B.n686 B.n685 71.676
R2086 B.n689 B.n688 71.676
R2087 B.n450 B.n449 71.676
R2088 B.n452 B.n446 71.676
R2089 B.n459 B.n458 71.676
R2090 B.n460 B.n444 71.676
R2091 B.n467 B.n466 71.676
R2092 B.n468 B.n442 71.676
R2093 B.n475 B.n474 71.676
R2094 B.n476 B.n440 71.676
R2095 B.n483 B.n482 71.676
R2096 B.n484 B.n438 71.676
R2097 B.n491 B.n490 71.676
R2098 B.n492 B.n436 71.676
R2099 B.n499 B.n498 71.676
R2100 B.n500 B.n434 71.676
R2101 B.n507 B.n506 71.676
R2102 B.n508 B.n432 71.676
R2103 B.n515 B.n514 71.676
R2104 B.n516 B.n430 71.676
R2105 B.n523 B.n522 71.676
R2106 B.n524 B.n428 71.676
R2107 B.n531 B.n530 71.676
R2108 B.n532 B.n426 71.676
R2109 B.n539 B.n538 71.676
R2110 B.n540 B.n424 71.676
R2111 B.n547 B.n546 71.676
R2112 B.n548 B.n422 71.676
R2113 B.n555 B.n554 71.676
R2114 B.n556 B.n418 71.676
R2115 B.n564 B.n563 71.676
R2116 B.n565 B.n416 71.676
R2117 B.n572 B.n571 71.676
R2118 B.n573 B.n414 71.676
R2119 B.n583 B.n582 71.676
R2120 B.n584 B.n412 71.676
R2121 B.n591 B.n590 71.676
R2122 B.n592 B.n410 71.676
R2123 B.n599 B.n598 71.676
R2124 B.n600 B.n408 71.676
R2125 B.n607 B.n606 71.676
R2126 B.n608 B.n406 71.676
R2127 B.n615 B.n614 71.676
R2128 B.n616 B.n404 71.676
R2129 B.n623 B.n622 71.676
R2130 B.n624 B.n402 71.676
R2131 B.n631 B.n630 71.676
R2132 B.n632 B.n400 71.676
R2133 B.n639 B.n638 71.676
R2134 B.n640 B.n398 71.676
R2135 B.n647 B.n646 71.676
R2136 B.n648 B.n396 71.676
R2137 B.n655 B.n654 71.676
R2138 B.n656 B.n394 71.676
R2139 B.n663 B.n662 71.676
R2140 B.n664 B.n392 71.676
R2141 B.n671 B.n670 71.676
R2142 B.n672 B.n390 71.676
R2143 B.n679 B.n678 71.676
R2144 B.n680 B.n388 71.676
R2145 B.n687 B.n686 71.676
R2146 B.n690 B.n689 71.676
R2147 B.n831 B.n830 71.676
R2148 B.n831 B.n2 71.676
R2149 B.n107 B.n106 59.5399
R2150 B.n104 B.n103 59.5399
R2151 B.n579 B.n578 59.5399
R2152 B.n559 B.n420 59.5399
R2153 B.n695 B.n384 56.9953
R2154 B.n788 B.n787 56.9953
R2155 B.n695 B.n380 33.7018
R2156 B.n701 B.n380 33.7018
R2157 B.n701 B.n376 33.7018
R2158 B.n708 B.n376 33.7018
R2159 B.n708 B.n707 33.7018
R2160 B.n714 B.n369 33.7018
R2161 B.n720 B.n369 33.7018
R2162 B.n720 B.n365 33.7018
R2163 B.n726 B.n365 33.7018
R2164 B.n726 B.n361 33.7018
R2165 B.n732 B.n361 33.7018
R2166 B.n738 B.n357 33.7018
R2167 B.n738 B.n353 33.7018
R2168 B.n745 B.n353 33.7018
R2169 B.n751 B.n349 33.7018
R2170 B.n751 B.n4 33.7018
R2171 B.n829 B.n4 33.7018
R2172 B.n829 B.n828 33.7018
R2173 B.n828 B.n827 33.7018
R2174 B.n827 B.n8 33.7018
R2175 B.n760 B.n8 33.7018
R2176 B.n820 B.n819 33.7018
R2177 B.n819 B.n818 33.7018
R2178 B.n818 B.n15 33.7018
R2179 B.n812 B.n811 33.7018
R2180 B.n811 B.n810 33.7018
R2181 B.n810 B.n22 33.7018
R2182 B.n804 B.n22 33.7018
R2183 B.n804 B.n803 33.7018
R2184 B.n803 B.n802 33.7018
R2185 B.n796 B.n32 33.7018
R2186 B.n796 B.n795 33.7018
R2187 B.n795 B.n794 33.7018
R2188 B.n794 B.n36 33.7018
R2189 B.n788 B.n36 33.7018
R2190 B.n697 B.n382 29.8151
R2191 B.n693 B.n692 29.8151
R2192 B.n784 B.n783 29.8151
R2193 B.n790 B.n38 29.8151
R2194 B.n745 B.t0 28.7457
R2195 B.n820 B.t2 28.7457
R2196 B.n106 B.n105 26.9581
R2197 B.n103 B.n102 26.9581
R2198 B.n578 B.n577 26.9581
R2199 B.n420 B.n419 26.9581
R2200 B.n732 B.t3 25.7721
R2201 B.n812 B.t1 25.7721
R2202 B B.n832 18.0485
R2203 B.n714 B.t5 17.8424
R2204 B.n802 B.t12 17.8424
R2205 B.n707 B.t5 15.8599
R2206 B.n32 B.t12 15.8599
R2207 B.n698 B.n697 10.6151
R2208 B.n699 B.n698 10.6151
R2209 B.n699 B.n374 10.6151
R2210 B.n710 B.n374 10.6151
R2211 B.n711 B.n710 10.6151
R2212 B.n712 B.n711 10.6151
R2213 B.n712 B.n367 10.6151
R2214 B.n722 B.n367 10.6151
R2215 B.n723 B.n722 10.6151
R2216 B.n724 B.n723 10.6151
R2217 B.n724 B.n359 10.6151
R2218 B.n734 B.n359 10.6151
R2219 B.n735 B.n734 10.6151
R2220 B.n736 B.n735 10.6151
R2221 B.n736 B.n351 10.6151
R2222 B.n747 B.n351 10.6151
R2223 B.n748 B.n747 10.6151
R2224 B.n749 B.n748 10.6151
R2225 B.n749 B.n0 10.6151
R2226 B.n448 B.n382 10.6151
R2227 B.n448 B.n447 10.6151
R2228 B.n454 B.n447 10.6151
R2229 B.n455 B.n454 10.6151
R2230 B.n456 B.n455 10.6151
R2231 B.n456 B.n445 10.6151
R2232 B.n462 B.n445 10.6151
R2233 B.n463 B.n462 10.6151
R2234 B.n464 B.n463 10.6151
R2235 B.n464 B.n443 10.6151
R2236 B.n470 B.n443 10.6151
R2237 B.n471 B.n470 10.6151
R2238 B.n472 B.n471 10.6151
R2239 B.n472 B.n441 10.6151
R2240 B.n478 B.n441 10.6151
R2241 B.n479 B.n478 10.6151
R2242 B.n480 B.n479 10.6151
R2243 B.n480 B.n439 10.6151
R2244 B.n486 B.n439 10.6151
R2245 B.n487 B.n486 10.6151
R2246 B.n488 B.n487 10.6151
R2247 B.n488 B.n437 10.6151
R2248 B.n494 B.n437 10.6151
R2249 B.n495 B.n494 10.6151
R2250 B.n496 B.n495 10.6151
R2251 B.n496 B.n435 10.6151
R2252 B.n502 B.n435 10.6151
R2253 B.n503 B.n502 10.6151
R2254 B.n504 B.n503 10.6151
R2255 B.n504 B.n433 10.6151
R2256 B.n510 B.n433 10.6151
R2257 B.n511 B.n510 10.6151
R2258 B.n512 B.n511 10.6151
R2259 B.n512 B.n431 10.6151
R2260 B.n518 B.n431 10.6151
R2261 B.n519 B.n518 10.6151
R2262 B.n520 B.n519 10.6151
R2263 B.n520 B.n429 10.6151
R2264 B.n526 B.n429 10.6151
R2265 B.n527 B.n526 10.6151
R2266 B.n528 B.n527 10.6151
R2267 B.n528 B.n427 10.6151
R2268 B.n534 B.n427 10.6151
R2269 B.n535 B.n534 10.6151
R2270 B.n536 B.n535 10.6151
R2271 B.n536 B.n425 10.6151
R2272 B.n542 B.n425 10.6151
R2273 B.n543 B.n542 10.6151
R2274 B.n544 B.n543 10.6151
R2275 B.n544 B.n423 10.6151
R2276 B.n550 B.n423 10.6151
R2277 B.n551 B.n550 10.6151
R2278 B.n552 B.n551 10.6151
R2279 B.n552 B.n421 10.6151
R2280 B.n558 B.n421 10.6151
R2281 B.n561 B.n560 10.6151
R2282 B.n561 B.n417 10.6151
R2283 B.n567 B.n417 10.6151
R2284 B.n568 B.n567 10.6151
R2285 B.n569 B.n568 10.6151
R2286 B.n569 B.n415 10.6151
R2287 B.n575 B.n415 10.6151
R2288 B.n576 B.n575 10.6151
R2289 B.n580 B.n576 10.6151
R2290 B.n586 B.n413 10.6151
R2291 B.n587 B.n586 10.6151
R2292 B.n588 B.n587 10.6151
R2293 B.n588 B.n411 10.6151
R2294 B.n594 B.n411 10.6151
R2295 B.n595 B.n594 10.6151
R2296 B.n596 B.n595 10.6151
R2297 B.n596 B.n409 10.6151
R2298 B.n602 B.n409 10.6151
R2299 B.n603 B.n602 10.6151
R2300 B.n604 B.n603 10.6151
R2301 B.n604 B.n407 10.6151
R2302 B.n610 B.n407 10.6151
R2303 B.n611 B.n610 10.6151
R2304 B.n612 B.n611 10.6151
R2305 B.n612 B.n405 10.6151
R2306 B.n618 B.n405 10.6151
R2307 B.n619 B.n618 10.6151
R2308 B.n620 B.n619 10.6151
R2309 B.n620 B.n403 10.6151
R2310 B.n626 B.n403 10.6151
R2311 B.n627 B.n626 10.6151
R2312 B.n628 B.n627 10.6151
R2313 B.n628 B.n401 10.6151
R2314 B.n634 B.n401 10.6151
R2315 B.n635 B.n634 10.6151
R2316 B.n636 B.n635 10.6151
R2317 B.n636 B.n399 10.6151
R2318 B.n642 B.n399 10.6151
R2319 B.n643 B.n642 10.6151
R2320 B.n644 B.n643 10.6151
R2321 B.n644 B.n397 10.6151
R2322 B.n650 B.n397 10.6151
R2323 B.n651 B.n650 10.6151
R2324 B.n652 B.n651 10.6151
R2325 B.n652 B.n395 10.6151
R2326 B.n658 B.n395 10.6151
R2327 B.n659 B.n658 10.6151
R2328 B.n660 B.n659 10.6151
R2329 B.n660 B.n393 10.6151
R2330 B.n666 B.n393 10.6151
R2331 B.n667 B.n666 10.6151
R2332 B.n668 B.n667 10.6151
R2333 B.n668 B.n391 10.6151
R2334 B.n674 B.n391 10.6151
R2335 B.n675 B.n674 10.6151
R2336 B.n676 B.n675 10.6151
R2337 B.n676 B.n389 10.6151
R2338 B.n682 B.n389 10.6151
R2339 B.n683 B.n682 10.6151
R2340 B.n684 B.n683 10.6151
R2341 B.n684 B.n387 10.6151
R2342 B.n387 B.n386 10.6151
R2343 B.n691 B.n386 10.6151
R2344 B.n692 B.n691 10.6151
R2345 B.n693 B.n378 10.6151
R2346 B.n703 B.n378 10.6151
R2347 B.n704 B.n703 10.6151
R2348 B.n705 B.n704 10.6151
R2349 B.n705 B.n371 10.6151
R2350 B.n716 B.n371 10.6151
R2351 B.n717 B.n716 10.6151
R2352 B.n718 B.n717 10.6151
R2353 B.n718 B.n363 10.6151
R2354 B.n728 B.n363 10.6151
R2355 B.n729 B.n728 10.6151
R2356 B.n730 B.n729 10.6151
R2357 B.n730 B.n355 10.6151
R2358 B.n740 B.n355 10.6151
R2359 B.n741 B.n740 10.6151
R2360 B.n743 B.n741 10.6151
R2361 B.n743 B.n742 10.6151
R2362 B.n742 B.n347 10.6151
R2363 B.n754 B.n347 10.6151
R2364 B.n755 B.n754 10.6151
R2365 B.n756 B.n755 10.6151
R2366 B.n757 B.n756 10.6151
R2367 B.n758 B.n757 10.6151
R2368 B.n762 B.n758 10.6151
R2369 B.n763 B.n762 10.6151
R2370 B.n764 B.n763 10.6151
R2371 B.n765 B.n764 10.6151
R2372 B.n767 B.n765 10.6151
R2373 B.n768 B.n767 10.6151
R2374 B.n769 B.n768 10.6151
R2375 B.n770 B.n769 10.6151
R2376 B.n772 B.n770 10.6151
R2377 B.n773 B.n772 10.6151
R2378 B.n774 B.n773 10.6151
R2379 B.n775 B.n774 10.6151
R2380 B.n777 B.n775 10.6151
R2381 B.n778 B.n777 10.6151
R2382 B.n779 B.n778 10.6151
R2383 B.n780 B.n779 10.6151
R2384 B.n782 B.n780 10.6151
R2385 B.n783 B.n782 10.6151
R2386 B.n824 B.n1 10.6151
R2387 B.n824 B.n823 10.6151
R2388 B.n823 B.n822 10.6151
R2389 B.n822 B.n10 10.6151
R2390 B.n816 B.n10 10.6151
R2391 B.n816 B.n815 10.6151
R2392 B.n815 B.n814 10.6151
R2393 B.n814 B.n17 10.6151
R2394 B.n808 B.n17 10.6151
R2395 B.n808 B.n807 10.6151
R2396 B.n807 B.n806 10.6151
R2397 B.n806 B.n24 10.6151
R2398 B.n800 B.n24 10.6151
R2399 B.n800 B.n799 10.6151
R2400 B.n799 B.n798 10.6151
R2401 B.n798 B.n30 10.6151
R2402 B.n792 B.n30 10.6151
R2403 B.n792 B.n791 10.6151
R2404 B.n791 B.n790 10.6151
R2405 B.n108 B.n38 10.6151
R2406 B.n111 B.n108 10.6151
R2407 B.n112 B.n111 10.6151
R2408 B.n115 B.n112 10.6151
R2409 B.n116 B.n115 10.6151
R2410 B.n119 B.n116 10.6151
R2411 B.n120 B.n119 10.6151
R2412 B.n123 B.n120 10.6151
R2413 B.n124 B.n123 10.6151
R2414 B.n127 B.n124 10.6151
R2415 B.n128 B.n127 10.6151
R2416 B.n131 B.n128 10.6151
R2417 B.n132 B.n131 10.6151
R2418 B.n135 B.n132 10.6151
R2419 B.n136 B.n135 10.6151
R2420 B.n139 B.n136 10.6151
R2421 B.n140 B.n139 10.6151
R2422 B.n143 B.n140 10.6151
R2423 B.n144 B.n143 10.6151
R2424 B.n147 B.n144 10.6151
R2425 B.n148 B.n147 10.6151
R2426 B.n151 B.n148 10.6151
R2427 B.n152 B.n151 10.6151
R2428 B.n155 B.n152 10.6151
R2429 B.n156 B.n155 10.6151
R2430 B.n159 B.n156 10.6151
R2431 B.n160 B.n159 10.6151
R2432 B.n163 B.n160 10.6151
R2433 B.n164 B.n163 10.6151
R2434 B.n167 B.n164 10.6151
R2435 B.n168 B.n167 10.6151
R2436 B.n171 B.n168 10.6151
R2437 B.n172 B.n171 10.6151
R2438 B.n175 B.n172 10.6151
R2439 B.n176 B.n175 10.6151
R2440 B.n179 B.n176 10.6151
R2441 B.n180 B.n179 10.6151
R2442 B.n183 B.n180 10.6151
R2443 B.n184 B.n183 10.6151
R2444 B.n187 B.n184 10.6151
R2445 B.n188 B.n187 10.6151
R2446 B.n191 B.n188 10.6151
R2447 B.n192 B.n191 10.6151
R2448 B.n195 B.n192 10.6151
R2449 B.n196 B.n195 10.6151
R2450 B.n199 B.n196 10.6151
R2451 B.n200 B.n199 10.6151
R2452 B.n203 B.n200 10.6151
R2453 B.n204 B.n203 10.6151
R2454 B.n207 B.n204 10.6151
R2455 B.n208 B.n207 10.6151
R2456 B.n211 B.n208 10.6151
R2457 B.n212 B.n211 10.6151
R2458 B.n215 B.n212 10.6151
R2459 B.n216 B.n215 10.6151
R2460 B.n220 B.n219 10.6151
R2461 B.n223 B.n220 10.6151
R2462 B.n224 B.n223 10.6151
R2463 B.n227 B.n224 10.6151
R2464 B.n228 B.n227 10.6151
R2465 B.n231 B.n228 10.6151
R2466 B.n232 B.n231 10.6151
R2467 B.n235 B.n232 10.6151
R2468 B.n236 B.n235 10.6151
R2469 B.n240 B.n239 10.6151
R2470 B.n243 B.n240 10.6151
R2471 B.n244 B.n243 10.6151
R2472 B.n247 B.n244 10.6151
R2473 B.n248 B.n247 10.6151
R2474 B.n251 B.n248 10.6151
R2475 B.n252 B.n251 10.6151
R2476 B.n255 B.n252 10.6151
R2477 B.n256 B.n255 10.6151
R2478 B.n259 B.n256 10.6151
R2479 B.n260 B.n259 10.6151
R2480 B.n263 B.n260 10.6151
R2481 B.n264 B.n263 10.6151
R2482 B.n267 B.n264 10.6151
R2483 B.n268 B.n267 10.6151
R2484 B.n271 B.n268 10.6151
R2485 B.n272 B.n271 10.6151
R2486 B.n275 B.n272 10.6151
R2487 B.n276 B.n275 10.6151
R2488 B.n279 B.n276 10.6151
R2489 B.n280 B.n279 10.6151
R2490 B.n283 B.n280 10.6151
R2491 B.n284 B.n283 10.6151
R2492 B.n287 B.n284 10.6151
R2493 B.n288 B.n287 10.6151
R2494 B.n291 B.n288 10.6151
R2495 B.n292 B.n291 10.6151
R2496 B.n295 B.n292 10.6151
R2497 B.n296 B.n295 10.6151
R2498 B.n299 B.n296 10.6151
R2499 B.n300 B.n299 10.6151
R2500 B.n303 B.n300 10.6151
R2501 B.n304 B.n303 10.6151
R2502 B.n307 B.n304 10.6151
R2503 B.n308 B.n307 10.6151
R2504 B.n311 B.n308 10.6151
R2505 B.n312 B.n311 10.6151
R2506 B.n315 B.n312 10.6151
R2507 B.n316 B.n315 10.6151
R2508 B.n319 B.n316 10.6151
R2509 B.n320 B.n319 10.6151
R2510 B.n323 B.n320 10.6151
R2511 B.n324 B.n323 10.6151
R2512 B.n327 B.n324 10.6151
R2513 B.n328 B.n327 10.6151
R2514 B.n331 B.n328 10.6151
R2515 B.n332 B.n331 10.6151
R2516 B.n335 B.n332 10.6151
R2517 B.n336 B.n335 10.6151
R2518 B.n339 B.n336 10.6151
R2519 B.n340 B.n339 10.6151
R2520 B.n343 B.n340 10.6151
R2521 B.n345 B.n343 10.6151
R2522 B.n346 B.n345 10.6151
R2523 B.n784 B.n346 10.6151
R2524 B.n559 B.n558 9.36635
R2525 B.n579 B.n413 9.36635
R2526 B.n216 B.n107 9.36635
R2527 B.n239 B.n104 9.36635
R2528 B.n832 B.n0 8.11757
R2529 B.n832 B.n1 8.11757
R2530 B.t3 B.n357 7.93021
R2531 B.t1 B.n15 7.93021
R2532 B.t0 B.n349 4.95657
R2533 B.n760 B.t2 4.95657
R2534 B.n560 B.n559 1.24928
R2535 B.n580 B.n579 1.24928
R2536 B.n219 B.n107 1.24928
R2537 B.n236 B.n104 1.24928
R2538 VN.n0 VN.t1 440.812
R2539 VN.n1 VN.t2 440.812
R2540 VN.n1 VN.t3 440.724
R2541 VN.n0 VN.t0 440.724
R2542 VN VN.n1 76.9023
R2543 VN VN.n0 31.2622
R2544 VDD2.n2 VDD2.n0 104.948
R2545 VDD2.n2 VDD2.n1 63.0519
R2546 VDD2.n1 VDD2.t0 1.17071
R2547 VDD2.n1 VDD2.t1 1.17071
R2548 VDD2.n0 VDD2.t2 1.17071
R2549 VDD2.n0 VDD2.t3 1.17071
R2550 VDD2 VDD2.n2 0.0586897
C0 VDD1 VDD2 0.65288f
C1 VP VN 5.99385f
C2 VN VTAIL 4.63084f
C3 VP VTAIL 4.64494f
C4 VDD2 VN 5.15118f
C5 VP VDD2 0.296091f
C6 VDD2 VTAIL 7.75613f
C7 VDD1 VN 0.147387f
C8 VP VDD1 5.29954f
C9 VDD1 VTAIL 7.71225f
C10 VDD2 B 3.291714f
C11 VDD1 B 7.539269f
C12 VTAIL B 11.909898f
C13 VN B 9.047919f
C14 VP B 6.007596f
C15 VDD2.t2 B 0.365179f
C16 VDD2.t3 B 0.365179f
C17 VDD2.n0 B 4.09259f
C18 VDD2.t0 B 0.365179f
C19 VDD2.t1 B 0.365179f
C20 VDD2.n1 B 3.32119f
C21 VDD2.n2 B 4.01417f
C22 VN.t1 B 2.13399f
C23 VN.t0 B 2.13382f
C24 VN.n0 B 1.52601f
C25 VN.t2 B 2.13399f
C26 VN.t3 B 2.13382f
C27 VN.n1 B 2.76639f
C28 VTAIL.n0 B 0.021927f
C29 VTAIL.n1 B 0.015306f
C30 VTAIL.n2 B 0.008225f
C31 VTAIL.n3 B 0.019441f
C32 VTAIL.n4 B 0.008709f
C33 VTAIL.n5 B 0.015306f
C34 VTAIL.n6 B 0.008225f
C35 VTAIL.n7 B 0.019441f
C36 VTAIL.n8 B 0.008709f
C37 VTAIL.n9 B 0.015306f
C38 VTAIL.n10 B 0.008225f
C39 VTAIL.n11 B 0.019441f
C40 VTAIL.n12 B 0.008709f
C41 VTAIL.n13 B 0.015306f
C42 VTAIL.n14 B 0.008225f
C43 VTAIL.n15 B 0.019441f
C44 VTAIL.n16 B 0.008709f
C45 VTAIL.n17 B 0.015306f
C46 VTAIL.n18 B 0.008225f
C47 VTAIL.n19 B 0.019441f
C48 VTAIL.n20 B 0.008709f
C49 VTAIL.n21 B 0.015306f
C50 VTAIL.n22 B 0.008225f
C51 VTAIL.n23 B 0.019441f
C52 VTAIL.n24 B 0.008709f
C53 VTAIL.n25 B 0.015306f
C54 VTAIL.n26 B 0.008225f
C55 VTAIL.n27 B 0.019441f
C56 VTAIL.n28 B 0.008709f
C57 VTAIL.n29 B 0.107199f
C58 VTAIL.t2 B 0.032156f
C59 VTAIL.n30 B 0.01458f
C60 VTAIL.n31 B 0.011484f
C61 VTAIL.n32 B 0.008225f
C62 VTAIL.n33 B 1.13053f
C63 VTAIL.n34 B 0.015306f
C64 VTAIL.n35 B 0.008225f
C65 VTAIL.n36 B 0.008709f
C66 VTAIL.n37 B 0.019441f
C67 VTAIL.n38 B 0.019441f
C68 VTAIL.n39 B 0.008709f
C69 VTAIL.n40 B 0.008225f
C70 VTAIL.n41 B 0.015306f
C71 VTAIL.n42 B 0.015306f
C72 VTAIL.n43 B 0.008225f
C73 VTAIL.n44 B 0.008709f
C74 VTAIL.n45 B 0.019441f
C75 VTAIL.n46 B 0.019441f
C76 VTAIL.n47 B 0.008709f
C77 VTAIL.n48 B 0.008225f
C78 VTAIL.n49 B 0.015306f
C79 VTAIL.n50 B 0.015306f
C80 VTAIL.n51 B 0.008225f
C81 VTAIL.n52 B 0.008709f
C82 VTAIL.n53 B 0.019441f
C83 VTAIL.n54 B 0.019441f
C84 VTAIL.n55 B 0.008709f
C85 VTAIL.n56 B 0.008225f
C86 VTAIL.n57 B 0.015306f
C87 VTAIL.n58 B 0.015306f
C88 VTAIL.n59 B 0.008225f
C89 VTAIL.n60 B 0.008709f
C90 VTAIL.n61 B 0.019441f
C91 VTAIL.n62 B 0.019441f
C92 VTAIL.n63 B 0.008709f
C93 VTAIL.n64 B 0.008225f
C94 VTAIL.n65 B 0.015306f
C95 VTAIL.n66 B 0.015306f
C96 VTAIL.n67 B 0.008225f
C97 VTAIL.n68 B 0.008709f
C98 VTAIL.n69 B 0.019441f
C99 VTAIL.n70 B 0.019441f
C100 VTAIL.n71 B 0.019441f
C101 VTAIL.n72 B 0.008709f
C102 VTAIL.n73 B 0.008225f
C103 VTAIL.n74 B 0.015306f
C104 VTAIL.n75 B 0.015306f
C105 VTAIL.n76 B 0.008225f
C106 VTAIL.n77 B 0.008467f
C107 VTAIL.n78 B 0.008467f
C108 VTAIL.n79 B 0.019441f
C109 VTAIL.n80 B 0.019441f
C110 VTAIL.n81 B 0.008709f
C111 VTAIL.n82 B 0.008225f
C112 VTAIL.n83 B 0.015306f
C113 VTAIL.n84 B 0.015306f
C114 VTAIL.n85 B 0.008225f
C115 VTAIL.n86 B 0.008709f
C116 VTAIL.n87 B 0.019441f
C117 VTAIL.n88 B 0.042816f
C118 VTAIL.n89 B 0.008709f
C119 VTAIL.n90 B 0.008225f
C120 VTAIL.n91 B 0.037889f
C121 VTAIL.n92 B 0.024107f
C122 VTAIL.n93 B 0.070082f
C123 VTAIL.n94 B 0.021927f
C124 VTAIL.n95 B 0.015306f
C125 VTAIL.n96 B 0.008225f
C126 VTAIL.n97 B 0.019441f
C127 VTAIL.n98 B 0.008709f
C128 VTAIL.n99 B 0.015306f
C129 VTAIL.n100 B 0.008225f
C130 VTAIL.n101 B 0.019441f
C131 VTAIL.n102 B 0.008709f
C132 VTAIL.n103 B 0.015306f
C133 VTAIL.n104 B 0.008225f
C134 VTAIL.n105 B 0.019441f
C135 VTAIL.n106 B 0.008709f
C136 VTAIL.n107 B 0.015306f
C137 VTAIL.n108 B 0.008225f
C138 VTAIL.n109 B 0.019441f
C139 VTAIL.n110 B 0.008709f
C140 VTAIL.n111 B 0.015306f
C141 VTAIL.n112 B 0.008225f
C142 VTAIL.n113 B 0.019441f
C143 VTAIL.n114 B 0.008709f
C144 VTAIL.n115 B 0.015306f
C145 VTAIL.n116 B 0.008225f
C146 VTAIL.n117 B 0.019441f
C147 VTAIL.n118 B 0.008709f
C148 VTAIL.n119 B 0.015306f
C149 VTAIL.n120 B 0.008225f
C150 VTAIL.n121 B 0.019441f
C151 VTAIL.n122 B 0.008709f
C152 VTAIL.n123 B 0.107199f
C153 VTAIL.t6 B 0.032156f
C154 VTAIL.n124 B 0.01458f
C155 VTAIL.n125 B 0.011484f
C156 VTAIL.n126 B 0.008225f
C157 VTAIL.n127 B 1.13053f
C158 VTAIL.n128 B 0.015306f
C159 VTAIL.n129 B 0.008225f
C160 VTAIL.n130 B 0.008709f
C161 VTAIL.n131 B 0.019441f
C162 VTAIL.n132 B 0.019441f
C163 VTAIL.n133 B 0.008709f
C164 VTAIL.n134 B 0.008225f
C165 VTAIL.n135 B 0.015306f
C166 VTAIL.n136 B 0.015306f
C167 VTAIL.n137 B 0.008225f
C168 VTAIL.n138 B 0.008709f
C169 VTAIL.n139 B 0.019441f
C170 VTAIL.n140 B 0.019441f
C171 VTAIL.n141 B 0.008709f
C172 VTAIL.n142 B 0.008225f
C173 VTAIL.n143 B 0.015306f
C174 VTAIL.n144 B 0.015306f
C175 VTAIL.n145 B 0.008225f
C176 VTAIL.n146 B 0.008709f
C177 VTAIL.n147 B 0.019441f
C178 VTAIL.n148 B 0.019441f
C179 VTAIL.n149 B 0.008709f
C180 VTAIL.n150 B 0.008225f
C181 VTAIL.n151 B 0.015306f
C182 VTAIL.n152 B 0.015306f
C183 VTAIL.n153 B 0.008225f
C184 VTAIL.n154 B 0.008709f
C185 VTAIL.n155 B 0.019441f
C186 VTAIL.n156 B 0.019441f
C187 VTAIL.n157 B 0.008709f
C188 VTAIL.n158 B 0.008225f
C189 VTAIL.n159 B 0.015306f
C190 VTAIL.n160 B 0.015306f
C191 VTAIL.n161 B 0.008225f
C192 VTAIL.n162 B 0.008709f
C193 VTAIL.n163 B 0.019441f
C194 VTAIL.n164 B 0.019441f
C195 VTAIL.n165 B 0.019441f
C196 VTAIL.n166 B 0.008709f
C197 VTAIL.n167 B 0.008225f
C198 VTAIL.n168 B 0.015306f
C199 VTAIL.n169 B 0.015306f
C200 VTAIL.n170 B 0.008225f
C201 VTAIL.n171 B 0.008467f
C202 VTAIL.n172 B 0.008467f
C203 VTAIL.n173 B 0.019441f
C204 VTAIL.n174 B 0.019441f
C205 VTAIL.n175 B 0.008709f
C206 VTAIL.n176 B 0.008225f
C207 VTAIL.n177 B 0.015306f
C208 VTAIL.n178 B 0.015306f
C209 VTAIL.n179 B 0.008225f
C210 VTAIL.n180 B 0.008709f
C211 VTAIL.n181 B 0.019441f
C212 VTAIL.n182 B 0.042816f
C213 VTAIL.n183 B 0.008709f
C214 VTAIL.n184 B 0.008225f
C215 VTAIL.n185 B 0.037889f
C216 VTAIL.n186 B 0.024107f
C217 VTAIL.n187 B 0.096762f
C218 VTAIL.n188 B 0.021927f
C219 VTAIL.n189 B 0.015306f
C220 VTAIL.n190 B 0.008225f
C221 VTAIL.n191 B 0.019441f
C222 VTAIL.n192 B 0.008709f
C223 VTAIL.n193 B 0.015306f
C224 VTAIL.n194 B 0.008225f
C225 VTAIL.n195 B 0.019441f
C226 VTAIL.n196 B 0.008709f
C227 VTAIL.n197 B 0.015306f
C228 VTAIL.n198 B 0.008225f
C229 VTAIL.n199 B 0.019441f
C230 VTAIL.n200 B 0.008709f
C231 VTAIL.n201 B 0.015306f
C232 VTAIL.n202 B 0.008225f
C233 VTAIL.n203 B 0.019441f
C234 VTAIL.n204 B 0.008709f
C235 VTAIL.n205 B 0.015306f
C236 VTAIL.n206 B 0.008225f
C237 VTAIL.n207 B 0.019441f
C238 VTAIL.n208 B 0.008709f
C239 VTAIL.n209 B 0.015306f
C240 VTAIL.n210 B 0.008225f
C241 VTAIL.n211 B 0.019441f
C242 VTAIL.n212 B 0.008709f
C243 VTAIL.n213 B 0.015306f
C244 VTAIL.n214 B 0.008225f
C245 VTAIL.n215 B 0.019441f
C246 VTAIL.n216 B 0.008709f
C247 VTAIL.n217 B 0.107199f
C248 VTAIL.t4 B 0.032156f
C249 VTAIL.n218 B 0.01458f
C250 VTAIL.n219 B 0.011484f
C251 VTAIL.n220 B 0.008225f
C252 VTAIL.n221 B 1.13053f
C253 VTAIL.n222 B 0.015306f
C254 VTAIL.n223 B 0.008225f
C255 VTAIL.n224 B 0.008709f
C256 VTAIL.n225 B 0.019441f
C257 VTAIL.n226 B 0.019441f
C258 VTAIL.n227 B 0.008709f
C259 VTAIL.n228 B 0.008225f
C260 VTAIL.n229 B 0.015306f
C261 VTAIL.n230 B 0.015306f
C262 VTAIL.n231 B 0.008225f
C263 VTAIL.n232 B 0.008709f
C264 VTAIL.n233 B 0.019441f
C265 VTAIL.n234 B 0.019441f
C266 VTAIL.n235 B 0.008709f
C267 VTAIL.n236 B 0.008225f
C268 VTAIL.n237 B 0.015306f
C269 VTAIL.n238 B 0.015306f
C270 VTAIL.n239 B 0.008225f
C271 VTAIL.n240 B 0.008709f
C272 VTAIL.n241 B 0.019441f
C273 VTAIL.n242 B 0.019441f
C274 VTAIL.n243 B 0.008709f
C275 VTAIL.n244 B 0.008225f
C276 VTAIL.n245 B 0.015306f
C277 VTAIL.n246 B 0.015306f
C278 VTAIL.n247 B 0.008225f
C279 VTAIL.n248 B 0.008709f
C280 VTAIL.n249 B 0.019441f
C281 VTAIL.n250 B 0.019441f
C282 VTAIL.n251 B 0.008709f
C283 VTAIL.n252 B 0.008225f
C284 VTAIL.n253 B 0.015306f
C285 VTAIL.n254 B 0.015306f
C286 VTAIL.n255 B 0.008225f
C287 VTAIL.n256 B 0.008709f
C288 VTAIL.n257 B 0.019441f
C289 VTAIL.n258 B 0.019441f
C290 VTAIL.n259 B 0.019441f
C291 VTAIL.n260 B 0.008709f
C292 VTAIL.n261 B 0.008225f
C293 VTAIL.n262 B 0.015306f
C294 VTAIL.n263 B 0.015306f
C295 VTAIL.n264 B 0.008225f
C296 VTAIL.n265 B 0.008467f
C297 VTAIL.n266 B 0.008467f
C298 VTAIL.n267 B 0.019441f
C299 VTAIL.n268 B 0.019441f
C300 VTAIL.n269 B 0.008709f
C301 VTAIL.n270 B 0.008225f
C302 VTAIL.n271 B 0.015306f
C303 VTAIL.n272 B 0.015306f
C304 VTAIL.n273 B 0.008225f
C305 VTAIL.n274 B 0.008709f
C306 VTAIL.n275 B 0.019441f
C307 VTAIL.n276 B 0.042816f
C308 VTAIL.n277 B 0.008709f
C309 VTAIL.n278 B 0.008225f
C310 VTAIL.n279 B 0.037889f
C311 VTAIL.n280 B 0.024107f
C312 VTAIL.n281 B 1.06f
C313 VTAIL.n282 B 0.021927f
C314 VTAIL.n283 B 0.015306f
C315 VTAIL.n284 B 0.008225f
C316 VTAIL.n285 B 0.019441f
C317 VTAIL.n286 B 0.008709f
C318 VTAIL.n287 B 0.015306f
C319 VTAIL.n288 B 0.008225f
C320 VTAIL.n289 B 0.019441f
C321 VTAIL.n290 B 0.008709f
C322 VTAIL.n291 B 0.015306f
C323 VTAIL.n292 B 0.008225f
C324 VTAIL.n293 B 0.019441f
C325 VTAIL.n294 B 0.019441f
C326 VTAIL.n295 B 0.008709f
C327 VTAIL.n296 B 0.015306f
C328 VTAIL.n297 B 0.008225f
C329 VTAIL.n298 B 0.019441f
C330 VTAIL.n299 B 0.008709f
C331 VTAIL.n300 B 0.015306f
C332 VTAIL.n301 B 0.008225f
C333 VTAIL.n302 B 0.019441f
C334 VTAIL.n303 B 0.008709f
C335 VTAIL.n304 B 0.015306f
C336 VTAIL.n305 B 0.008225f
C337 VTAIL.n306 B 0.019441f
C338 VTAIL.n307 B 0.008709f
C339 VTAIL.n308 B 0.015306f
C340 VTAIL.n309 B 0.008225f
C341 VTAIL.n310 B 0.019441f
C342 VTAIL.n311 B 0.008709f
C343 VTAIL.n312 B 0.107199f
C344 VTAIL.t3 B 0.032156f
C345 VTAIL.n313 B 0.01458f
C346 VTAIL.n314 B 0.011484f
C347 VTAIL.n315 B 0.008225f
C348 VTAIL.n316 B 1.13053f
C349 VTAIL.n317 B 0.015306f
C350 VTAIL.n318 B 0.008225f
C351 VTAIL.n319 B 0.008709f
C352 VTAIL.n320 B 0.019441f
C353 VTAIL.n321 B 0.019441f
C354 VTAIL.n322 B 0.008709f
C355 VTAIL.n323 B 0.008225f
C356 VTAIL.n324 B 0.015306f
C357 VTAIL.n325 B 0.015306f
C358 VTAIL.n326 B 0.008225f
C359 VTAIL.n327 B 0.008709f
C360 VTAIL.n328 B 0.019441f
C361 VTAIL.n329 B 0.019441f
C362 VTAIL.n330 B 0.008709f
C363 VTAIL.n331 B 0.008225f
C364 VTAIL.n332 B 0.015306f
C365 VTAIL.n333 B 0.015306f
C366 VTAIL.n334 B 0.008225f
C367 VTAIL.n335 B 0.008709f
C368 VTAIL.n336 B 0.019441f
C369 VTAIL.n337 B 0.019441f
C370 VTAIL.n338 B 0.008709f
C371 VTAIL.n339 B 0.008225f
C372 VTAIL.n340 B 0.015306f
C373 VTAIL.n341 B 0.015306f
C374 VTAIL.n342 B 0.008225f
C375 VTAIL.n343 B 0.008709f
C376 VTAIL.n344 B 0.019441f
C377 VTAIL.n345 B 0.019441f
C378 VTAIL.n346 B 0.008709f
C379 VTAIL.n347 B 0.008225f
C380 VTAIL.n348 B 0.015306f
C381 VTAIL.n349 B 0.015306f
C382 VTAIL.n350 B 0.008225f
C383 VTAIL.n351 B 0.008709f
C384 VTAIL.n352 B 0.019441f
C385 VTAIL.n353 B 0.019441f
C386 VTAIL.n354 B 0.008709f
C387 VTAIL.n355 B 0.008225f
C388 VTAIL.n356 B 0.015306f
C389 VTAIL.n357 B 0.015306f
C390 VTAIL.n358 B 0.008225f
C391 VTAIL.n359 B 0.008467f
C392 VTAIL.n360 B 0.008467f
C393 VTAIL.n361 B 0.019441f
C394 VTAIL.n362 B 0.019441f
C395 VTAIL.n363 B 0.008709f
C396 VTAIL.n364 B 0.008225f
C397 VTAIL.n365 B 0.015306f
C398 VTAIL.n366 B 0.015306f
C399 VTAIL.n367 B 0.008225f
C400 VTAIL.n368 B 0.008709f
C401 VTAIL.n369 B 0.019441f
C402 VTAIL.n370 B 0.042816f
C403 VTAIL.n371 B 0.008709f
C404 VTAIL.n372 B 0.008225f
C405 VTAIL.n373 B 0.037889f
C406 VTAIL.n374 B 0.024107f
C407 VTAIL.n375 B 1.06f
C408 VTAIL.n376 B 0.021927f
C409 VTAIL.n377 B 0.015306f
C410 VTAIL.n378 B 0.008225f
C411 VTAIL.n379 B 0.019441f
C412 VTAIL.n380 B 0.008709f
C413 VTAIL.n381 B 0.015306f
C414 VTAIL.n382 B 0.008225f
C415 VTAIL.n383 B 0.019441f
C416 VTAIL.n384 B 0.008709f
C417 VTAIL.n385 B 0.015306f
C418 VTAIL.n386 B 0.008225f
C419 VTAIL.n387 B 0.019441f
C420 VTAIL.n388 B 0.019441f
C421 VTAIL.n389 B 0.008709f
C422 VTAIL.n390 B 0.015306f
C423 VTAIL.n391 B 0.008225f
C424 VTAIL.n392 B 0.019441f
C425 VTAIL.n393 B 0.008709f
C426 VTAIL.n394 B 0.015306f
C427 VTAIL.n395 B 0.008225f
C428 VTAIL.n396 B 0.019441f
C429 VTAIL.n397 B 0.008709f
C430 VTAIL.n398 B 0.015306f
C431 VTAIL.n399 B 0.008225f
C432 VTAIL.n400 B 0.019441f
C433 VTAIL.n401 B 0.008709f
C434 VTAIL.n402 B 0.015306f
C435 VTAIL.n403 B 0.008225f
C436 VTAIL.n404 B 0.019441f
C437 VTAIL.n405 B 0.008709f
C438 VTAIL.n406 B 0.107199f
C439 VTAIL.t0 B 0.032156f
C440 VTAIL.n407 B 0.01458f
C441 VTAIL.n408 B 0.011484f
C442 VTAIL.n409 B 0.008225f
C443 VTAIL.n410 B 1.13053f
C444 VTAIL.n411 B 0.015306f
C445 VTAIL.n412 B 0.008225f
C446 VTAIL.n413 B 0.008709f
C447 VTAIL.n414 B 0.019441f
C448 VTAIL.n415 B 0.019441f
C449 VTAIL.n416 B 0.008709f
C450 VTAIL.n417 B 0.008225f
C451 VTAIL.n418 B 0.015306f
C452 VTAIL.n419 B 0.015306f
C453 VTAIL.n420 B 0.008225f
C454 VTAIL.n421 B 0.008709f
C455 VTAIL.n422 B 0.019441f
C456 VTAIL.n423 B 0.019441f
C457 VTAIL.n424 B 0.008709f
C458 VTAIL.n425 B 0.008225f
C459 VTAIL.n426 B 0.015306f
C460 VTAIL.n427 B 0.015306f
C461 VTAIL.n428 B 0.008225f
C462 VTAIL.n429 B 0.008709f
C463 VTAIL.n430 B 0.019441f
C464 VTAIL.n431 B 0.019441f
C465 VTAIL.n432 B 0.008709f
C466 VTAIL.n433 B 0.008225f
C467 VTAIL.n434 B 0.015306f
C468 VTAIL.n435 B 0.015306f
C469 VTAIL.n436 B 0.008225f
C470 VTAIL.n437 B 0.008709f
C471 VTAIL.n438 B 0.019441f
C472 VTAIL.n439 B 0.019441f
C473 VTAIL.n440 B 0.008709f
C474 VTAIL.n441 B 0.008225f
C475 VTAIL.n442 B 0.015306f
C476 VTAIL.n443 B 0.015306f
C477 VTAIL.n444 B 0.008225f
C478 VTAIL.n445 B 0.008709f
C479 VTAIL.n446 B 0.019441f
C480 VTAIL.n447 B 0.019441f
C481 VTAIL.n448 B 0.008709f
C482 VTAIL.n449 B 0.008225f
C483 VTAIL.n450 B 0.015306f
C484 VTAIL.n451 B 0.015306f
C485 VTAIL.n452 B 0.008225f
C486 VTAIL.n453 B 0.008467f
C487 VTAIL.n454 B 0.008467f
C488 VTAIL.n455 B 0.019441f
C489 VTAIL.n456 B 0.019441f
C490 VTAIL.n457 B 0.008709f
C491 VTAIL.n458 B 0.008225f
C492 VTAIL.n459 B 0.015306f
C493 VTAIL.n460 B 0.015306f
C494 VTAIL.n461 B 0.008225f
C495 VTAIL.n462 B 0.008709f
C496 VTAIL.n463 B 0.019441f
C497 VTAIL.n464 B 0.042816f
C498 VTAIL.n465 B 0.008709f
C499 VTAIL.n466 B 0.008225f
C500 VTAIL.n467 B 0.037889f
C501 VTAIL.n468 B 0.024107f
C502 VTAIL.n469 B 0.096762f
C503 VTAIL.n470 B 0.021927f
C504 VTAIL.n471 B 0.015306f
C505 VTAIL.n472 B 0.008225f
C506 VTAIL.n473 B 0.019441f
C507 VTAIL.n474 B 0.008709f
C508 VTAIL.n475 B 0.015306f
C509 VTAIL.n476 B 0.008225f
C510 VTAIL.n477 B 0.019441f
C511 VTAIL.n478 B 0.008709f
C512 VTAIL.n479 B 0.015306f
C513 VTAIL.n480 B 0.008225f
C514 VTAIL.n481 B 0.019441f
C515 VTAIL.n482 B 0.019441f
C516 VTAIL.n483 B 0.008709f
C517 VTAIL.n484 B 0.015306f
C518 VTAIL.n485 B 0.008225f
C519 VTAIL.n486 B 0.019441f
C520 VTAIL.n487 B 0.008709f
C521 VTAIL.n488 B 0.015306f
C522 VTAIL.n489 B 0.008225f
C523 VTAIL.n490 B 0.019441f
C524 VTAIL.n491 B 0.008709f
C525 VTAIL.n492 B 0.015306f
C526 VTAIL.n493 B 0.008225f
C527 VTAIL.n494 B 0.019441f
C528 VTAIL.n495 B 0.008709f
C529 VTAIL.n496 B 0.015306f
C530 VTAIL.n497 B 0.008225f
C531 VTAIL.n498 B 0.019441f
C532 VTAIL.n499 B 0.008709f
C533 VTAIL.n500 B 0.107199f
C534 VTAIL.t7 B 0.032156f
C535 VTAIL.n501 B 0.01458f
C536 VTAIL.n502 B 0.011484f
C537 VTAIL.n503 B 0.008225f
C538 VTAIL.n504 B 1.13053f
C539 VTAIL.n505 B 0.015306f
C540 VTAIL.n506 B 0.008225f
C541 VTAIL.n507 B 0.008709f
C542 VTAIL.n508 B 0.019441f
C543 VTAIL.n509 B 0.019441f
C544 VTAIL.n510 B 0.008709f
C545 VTAIL.n511 B 0.008225f
C546 VTAIL.n512 B 0.015306f
C547 VTAIL.n513 B 0.015306f
C548 VTAIL.n514 B 0.008225f
C549 VTAIL.n515 B 0.008709f
C550 VTAIL.n516 B 0.019441f
C551 VTAIL.n517 B 0.019441f
C552 VTAIL.n518 B 0.008709f
C553 VTAIL.n519 B 0.008225f
C554 VTAIL.n520 B 0.015306f
C555 VTAIL.n521 B 0.015306f
C556 VTAIL.n522 B 0.008225f
C557 VTAIL.n523 B 0.008709f
C558 VTAIL.n524 B 0.019441f
C559 VTAIL.n525 B 0.019441f
C560 VTAIL.n526 B 0.008709f
C561 VTAIL.n527 B 0.008225f
C562 VTAIL.n528 B 0.015306f
C563 VTAIL.n529 B 0.015306f
C564 VTAIL.n530 B 0.008225f
C565 VTAIL.n531 B 0.008709f
C566 VTAIL.n532 B 0.019441f
C567 VTAIL.n533 B 0.019441f
C568 VTAIL.n534 B 0.008709f
C569 VTAIL.n535 B 0.008225f
C570 VTAIL.n536 B 0.015306f
C571 VTAIL.n537 B 0.015306f
C572 VTAIL.n538 B 0.008225f
C573 VTAIL.n539 B 0.008709f
C574 VTAIL.n540 B 0.019441f
C575 VTAIL.n541 B 0.019441f
C576 VTAIL.n542 B 0.008709f
C577 VTAIL.n543 B 0.008225f
C578 VTAIL.n544 B 0.015306f
C579 VTAIL.n545 B 0.015306f
C580 VTAIL.n546 B 0.008225f
C581 VTAIL.n547 B 0.008467f
C582 VTAIL.n548 B 0.008467f
C583 VTAIL.n549 B 0.019441f
C584 VTAIL.n550 B 0.019441f
C585 VTAIL.n551 B 0.008709f
C586 VTAIL.n552 B 0.008225f
C587 VTAIL.n553 B 0.015306f
C588 VTAIL.n554 B 0.015306f
C589 VTAIL.n555 B 0.008225f
C590 VTAIL.n556 B 0.008709f
C591 VTAIL.n557 B 0.019441f
C592 VTAIL.n558 B 0.042816f
C593 VTAIL.n559 B 0.008709f
C594 VTAIL.n560 B 0.008225f
C595 VTAIL.n561 B 0.037889f
C596 VTAIL.n562 B 0.024107f
C597 VTAIL.n563 B 0.096762f
C598 VTAIL.n564 B 0.021927f
C599 VTAIL.n565 B 0.015306f
C600 VTAIL.n566 B 0.008225f
C601 VTAIL.n567 B 0.019441f
C602 VTAIL.n568 B 0.008709f
C603 VTAIL.n569 B 0.015306f
C604 VTAIL.n570 B 0.008225f
C605 VTAIL.n571 B 0.019441f
C606 VTAIL.n572 B 0.008709f
C607 VTAIL.n573 B 0.015306f
C608 VTAIL.n574 B 0.008225f
C609 VTAIL.n575 B 0.019441f
C610 VTAIL.n576 B 0.019441f
C611 VTAIL.n577 B 0.008709f
C612 VTAIL.n578 B 0.015306f
C613 VTAIL.n579 B 0.008225f
C614 VTAIL.n580 B 0.019441f
C615 VTAIL.n581 B 0.008709f
C616 VTAIL.n582 B 0.015306f
C617 VTAIL.n583 B 0.008225f
C618 VTAIL.n584 B 0.019441f
C619 VTAIL.n585 B 0.008709f
C620 VTAIL.n586 B 0.015306f
C621 VTAIL.n587 B 0.008225f
C622 VTAIL.n588 B 0.019441f
C623 VTAIL.n589 B 0.008709f
C624 VTAIL.n590 B 0.015306f
C625 VTAIL.n591 B 0.008225f
C626 VTAIL.n592 B 0.019441f
C627 VTAIL.n593 B 0.008709f
C628 VTAIL.n594 B 0.107199f
C629 VTAIL.t5 B 0.032156f
C630 VTAIL.n595 B 0.01458f
C631 VTAIL.n596 B 0.011484f
C632 VTAIL.n597 B 0.008225f
C633 VTAIL.n598 B 1.13053f
C634 VTAIL.n599 B 0.015306f
C635 VTAIL.n600 B 0.008225f
C636 VTAIL.n601 B 0.008709f
C637 VTAIL.n602 B 0.019441f
C638 VTAIL.n603 B 0.019441f
C639 VTAIL.n604 B 0.008709f
C640 VTAIL.n605 B 0.008225f
C641 VTAIL.n606 B 0.015306f
C642 VTAIL.n607 B 0.015306f
C643 VTAIL.n608 B 0.008225f
C644 VTAIL.n609 B 0.008709f
C645 VTAIL.n610 B 0.019441f
C646 VTAIL.n611 B 0.019441f
C647 VTAIL.n612 B 0.008709f
C648 VTAIL.n613 B 0.008225f
C649 VTAIL.n614 B 0.015306f
C650 VTAIL.n615 B 0.015306f
C651 VTAIL.n616 B 0.008225f
C652 VTAIL.n617 B 0.008709f
C653 VTAIL.n618 B 0.019441f
C654 VTAIL.n619 B 0.019441f
C655 VTAIL.n620 B 0.008709f
C656 VTAIL.n621 B 0.008225f
C657 VTAIL.n622 B 0.015306f
C658 VTAIL.n623 B 0.015306f
C659 VTAIL.n624 B 0.008225f
C660 VTAIL.n625 B 0.008709f
C661 VTAIL.n626 B 0.019441f
C662 VTAIL.n627 B 0.019441f
C663 VTAIL.n628 B 0.008709f
C664 VTAIL.n629 B 0.008225f
C665 VTAIL.n630 B 0.015306f
C666 VTAIL.n631 B 0.015306f
C667 VTAIL.n632 B 0.008225f
C668 VTAIL.n633 B 0.008709f
C669 VTAIL.n634 B 0.019441f
C670 VTAIL.n635 B 0.019441f
C671 VTAIL.n636 B 0.008709f
C672 VTAIL.n637 B 0.008225f
C673 VTAIL.n638 B 0.015306f
C674 VTAIL.n639 B 0.015306f
C675 VTAIL.n640 B 0.008225f
C676 VTAIL.n641 B 0.008467f
C677 VTAIL.n642 B 0.008467f
C678 VTAIL.n643 B 0.019441f
C679 VTAIL.n644 B 0.019441f
C680 VTAIL.n645 B 0.008709f
C681 VTAIL.n646 B 0.008225f
C682 VTAIL.n647 B 0.015306f
C683 VTAIL.n648 B 0.015306f
C684 VTAIL.n649 B 0.008225f
C685 VTAIL.n650 B 0.008709f
C686 VTAIL.n651 B 0.019441f
C687 VTAIL.n652 B 0.042816f
C688 VTAIL.n653 B 0.008709f
C689 VTAIL.n654 B 0.008225f
C690 VTAIL.n655 B 0.037889f
C691 VTAIL.n656 B 0.024107f
C692 VTAIL.n657 B 1.06f
C693 VTAIL.n658 B 0.021927f
C694 VTAIL.n659 B 0.015306f
C695 VTAIL.n660 B 0.008225f
C696 VTAIL.n661 B 0.019441f
C697 VTAIL.n662 B 0.008709f
C698 VTAIL.n663 B 0.015306f
C699 VTAIL.n664 B 0.008225f
C700 VTAIL.n665 B 0.019441f
C701 VTAIL.n666 B 0.008709f
C702 VTAIL.n667 B 0.015306f
C703 VTAIL.n668 B 0.008225f
C704 VTAIL.n669 B 0.019441f
C705 VTAIL.n670 B 0.008709f
C706 VTAIL.n671 B 0.015306f
C707 VTAIL.n672 B 0.008225f
C708 VTAIL.n673 B 0.019441f
C709 VTAIL.n674 B 0.008709f
C710 VTAIL.n675 B 0.015306f
C711 VTAIL.n676 B 0.008225f
C712 VTAIL.n677 B 0.019441f
C713 VTAIL.n678 B 0.008709f
C714 VTAIL.n679 B 0.015306f
C715 VTAIL.n680 B 0.008225f
C716 VTAIL.n681 B 0.019441f
C717 VTAIL.n682 B 0.008709f
C718 VTAIL.n683 B 0.015306f
C719 VTAIL.n684 B 0.008225f
C720 VTAIL.n685 B 0.019441f
C721 VTAIL.n686 B 0.008709f
C722 VTAIL.n687 B 0.107199f
C723 VTAIL.t1 B 0.032156f
C724 VTAIL.n688 B 0.01458f
C725 VTAIL.n689 B 0.011484f
C726 VTAIL.n690 B 0.008225f
C727 VTAIL.n691 B 1.13053f
C728 VTAIL.n692 B 0.015306f
C729 VTAIL.n693 B 0.008225f
C730 VTAIL.n694 B 0.008709f
C731 VTAIL.n695 B 0.019441f
C732 VTAIL.n696 B 0.019441f
C733 VTAIL.n697 B 0.008709f
C734 VTAIL.n698 B 0.008225f
C735 VTAIL.n699 B 0.015306f
C736 VTAIL.n700 B 0.015306f
C737 VTAIL.n701 B 0.008225f
C738 VTAIL.n702 B 0.008709f
C739 VTAIL.n703 B 0.019441f
C740 VTAIL.n704 B 0.019441f
C741 VTAIL.n705 B 0.008709f
C742 VTAIL.n706 B 0.008225f
C743 VTAIL.n707 B 0.015306f
C744 VTAIL.n708 B 0.015306f
C745 VTAIL.n709 B 0.008225f
C746 VTAIL.n710 B 0.008709f
C747 VTAIL.n711 B 0.019441f
C748 VTAIL.n712 B 0.019441f
C749 VTAIL.n713 B 0.008709f
C750 VTAIL.n714 B 0.008225f
C751 VTAIL.n715 B 0.015306f
C752 VTAIL.n716 B 0.015306f
C753 VTAIL.n717 B 0.008225f
C754 VTAIL.n718 B 0.008709f
C755 VTAIL.n719 B 0.019441f
C756 VTAIL.n720 B 0.019441f
C757 VTAIL.n721 B 0.008709f
C758 VTAIL.n722 B 0.008225f
C759 VTAIL.n723 B 0.015306f
C760 VTAIL.n724 B 0.015306f
C761 VTAIL.n725 B 0.008225f
C762 VTAIL.n726 B 0.008709f
C763 VTAIL.n727 B 0.019441f
C764 VTAIL.n728 B 0.019441f
C765 VTAIL.n729 B 0.019441f
C766 VTAIL.n730 B 0.008709f
C767 VTAIL.n731 B 0.008225f
C768 VTAIL.n732 B 0.015306f
C769 VTAIL.n733 B 0.015306f
C770 VTAIL.n734 B 0.008225f
C771 VTAIL.n735 B 0.008467f
C772 VTAIL.n736 B 0.008467f
C773 VTAIL.n737 B 0.019441f
C774 VTAIL.n738 B 0.019441f
C775 VTAIL.n739 B 0.008709f
C776 VTAIL.n740 B 0.008225f
C777 VTAIL.n741 B 0.015306f
C778 VTAIL.n742 B 0.015306f
C779 VTAIL.n743 B 0.008225f
C780 VTAIL.n744 B 0.008709f
C781 VTAIL.n745 B 0.019441f
C782 VTAIL.n746 B 0.042816f
C783 VTAIL.n747 B 0.008709f
C784 VTAIL.n748 B 0.008225f
C785 VTAIL.n749 B 0.037889f
C786 VTAIL.n750 B 0.024107f
C787 VTAIL.n751 B 1.02758f
C788 VDD1.t1 B 0.362367f
C789 VDD1.t3 B 0.362367f
C790 VDD1.n0 B 3.29593f
C791 VDD1.t2 B 0.362367f
C792 VDD1.t0 B 0.362367f
C793 VDD1.n1 B 4.08859f
C794 VP.t2 B 2.15523f
C795 VP.t0 B 2.15541f
C796 VP.n0 B 2.77728f
C797 VP.n1 B 2.86634f
C798 VP.t3 B 2.12145f
C799 VP.n2 B 0.803967f
C800 VP.t1 B 2.12145f
C801 VP.n3 B 0.803967f
C802 VP.n4 B 0.052964f
.ends

