* NGSPICE file created from diff_pair_sample_1443.ext - technology: sky130A

.subckt diff_pair_sample_1443 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VP.t0 VDD1.t7 w_n2660_n3676# sky130_fd_pr__pfet_01v8 ad=5.2806 pd=27.86 as=2.2341 ps=13.87 w=13.54 l=1.36
X1 VDD2.t7 VN.t0 VTAIL.t2 w_n2660_n3676# sky130_fd_pr__pfet_01v8 ad=2.2341 pd=13.87 as=2.2341 ps=13.87 w=13.54 l=1.36
X2 VTAIL.t4 VN.t1 VDD2.t6 w_n2660_n3676# sky130_fd_pr__pfet_01v8 ad=2.2341 pd=13.87 as=2.2341 ps=13.87 w=13.54 l=1.36
X3 VDD2.t5 VN.t2 VTAIL.t7 w_n2660_n3676# sky130_fd_pr__pfet_01v8 ad=2.2341 pd=13.87 as=2.2341 ps=13.87 w=13.54 l=1.36
X4 B.t11 B.t9 B.t10 w_n2660_n3676# sky130_fd_pr__pfet_01v8 ad=5.2806 pd=27.86 as=0 ps=0 w=13.54 l=1.36
X5 VDD1.t3 VP.t1 VTAIL.t14 w_n2660_n3676# sky130_fd_pr__pfet_01v8 ad=2.2341 pd=13.87 as=2.2341 ps=13.87 w=13.54 l=1.36
X6 VDD2.t4 VN.t3 VTAIL.t1 w_n2660_n3676# sky130_fd_pr__pfet_01v8 ad=2.2341 pd=13.87 as=5.2806 ps=27.86 w=13.54 l=1.36
X7 VDD2.t3 VN.t4 VTAIL.t3 w_n2660_n3676# sky130_fd_pr__pfet_01v8 ad=2.2341 pd=13.87 as=5.2806 ps=27.86 w=13.54 l=1.36
X8 B.t8 B.t6 B.t7 w_n2660_n3676# sky130_fd_pr__pfet_01v8 ad=5.2806 pd=27.86 as=0 ps=0 w=13.54 l=1.36
X9 VTAIL.t13 VP.t2 VDD1.t2 w_n2660_n3676# sky130_fd_pr__pfet_01v8 ad=5.2806 pd=27.86 as=2.2341 ps=13.87 w=13.54 l=1.36
X10 VDD1.t4 VP.t3 VTAIL.t12 w_n2660_n3676# sky130_fd_pr__pfet_01v8 ad=2.2341 pd=13.87 as=5.2806 ps=27.86 w=13.54 l=1.36
X11 B.t5 B.t3 B.t4 w_n2660_n3676# sky130_fd_pr__pfet_01v8 ad=5.2806 pd=27.86 as=0 ps=0 w=13.54 l=1.36
X12 VTAIL.t5 VN.t5 VDD2.t2 w_n2660_n3676# sky130_fd_pr__pfet_01v8 ad=2.2341 pd=13.87 as=2.2341 ps=13.87 w=13.54 l=1.36
X13 B.t2 B.t0 B.t1 w_n2660_n3676# sky130_fd_pr__pfet_01v8 ad=5.2806 pd=27.86 as=0 ps=0 w=13.54 l=1.36
X14 VTAIL.t0 VN.t6 VDD2.t1 w_n2660_n3676# sky130_fd_pr__pfet_01v8 ad=5.2806 pd=27.86 as=2.2341 ps=13.87 w=13.54 l=1.36
X15 VDD1.t6 VP.t4 VTAIL.t11 w_n2660_n3676# sky130_fd_pr__pfet_01v8 ad=2.2341 pd=13.87 as=2.2341 ps=13.87 w=13.54 l=1.36
X16 VTAIL.t10 VP.t5 VDD1.t5 w_n2660_n3676# sky130_fd_pr__pfet_01v8 ad=2.2341 pd=13.87 as=2.2341 ps=13.87 w=13.54 l=1.36
X17 VDD1.t0 VP.t6 VTAIL.t9 w_n2660_n3676# sky130_fd_pr__pfet_01v8 ad=2.2341 pd=13.87 as=5.2806 ps=27.86 w=13.54 l=1.36
X18 VTAIL.t8 VP.t7 VDD1.t1 w_n2660_n3676# sky130_fd_pr__pfet_01v8 ad=2.2341 pd=13.87 as=2.2341 ps=13.87 w=13.54 l=1.36
X19 VTAIL.t6 VN.t7 VDD2.t0 w_n2660_n3676# sky130_fd_pr__pfet_01v8 ad=5.2806 pd=27.86 as=2.2341 ps=13.87 w=13.54 l=1.36
R0 VP.n11 VP.t2 270.158
R1 VP.n5 VP.t0 239.938
R2 VP.n29 VP.t4 239.938
R3 VP.n36 VP.t5 239.938
R4 VP.n43 VP.t3 239.938
R5 VP.n23 VP.t6 239.938
R6 VP.n16 VP.t7 239.938
R7 VP.n10 VP.t1 239.938
R8 VP.n25 VP.n5 171.875
R9 VP.n44 VP.n43 171.875
R10 VP.n24 VP.n23 171.875
R11 VP.n12 VP.n9 161.3
R12 VP.n14 VP.n13 161.3
R13 VP.n15 VP.n8 161.3
R14 VP.n18 VP.n17 161.3
R15 VP.n19 VP.n7 161.3
R16 VP.n21 VP.n20 161.3
R17 VP.n22 VP.n6 161.3
R18 VP.n42 VP.n0 161.3
R19 VP.n41 VP.n40 161.3
R20 VP.n39 VP.n1 161.3
R21 VP.n38 VP.n37 161.3
R22 VP.n35 VP.n2 161.3
R23 VP.n34 VP.n33 161.3
R24 VP.n32 VP.n3 161.3
R25 VP.n31 VP.n30 161.3
R26 VP.n28 VP.n4 161.3
R27 VP.n27 VP.n26 161.3
R28 VP.n11 VP.n10 60.629
R29 VP.n35 VP.n34 56.5617
R30 VP.n15 VP.n14 56.5617
R31 VP.n30 VP.n28 46.3896
R32 VP.n41 VP.n1 46.3896
R33 VP.n21 VP.n7 46.3896
R34 VP.n25 VP.n24 46.2126
R35 VP.n28 VP.n27 34.7644
R36 VP.n42 VP.n41 34.7644
R37 VP.n22 VP.n21 34.7644
R38 VP.n12 VP.n11 26.9001
R39 VP.n34 VP.n3 24.5923
R40 VP.n37 VP.n35 24.5923
R41 VP.n17 VP.n15 24.5923
R42 VP.n14 VP.n9 24.5923
R43 VP.n30 VP.n29 19.9199
R44 VP.n36 VP.n1 19.9199
R45 VP.n16 VP.n7 19.9199
R46 VP.n27 VP.n5 14.0178
R47 VP.n43 VP.n42 14.0178
R48 VP.n23 VP.n22 14.0178
R49 VP.n29 VP.n3 4.67295
R50 VP.n37 VP.n36 4.67295
R51 VP.n17 VP.n16 4.67295
R52 VP.n10 VP.n9 4.67295
R53 VP.n13 VP.n12 0.189894
R54 VP.n13 VP.n8 0.189894
R55 VP.n18 VP.n8 0.189894
R56 VP.n19 VP.n18 0.189894
R57 VP.n20 VP.n19 0.189894
R58 VP.n20 VP.n6 0.189894
R59 VP.n24 VP.n6 0.189894
R60 VP.n26 VP.n25 0.189894
R61 VP.n26 VP.n4 0.189894
R62 VP.n31 VP.n4 0.189894
R63 VP.n32 VP.n31 0.189894
R64 VP.n33 VP.n32 0.189894
R65 VP.n33 VP.n2 0.189894
R66 VP.n38 VP.n2 0.189894
R67 VP.n39 VP.n38 0.189894
R68 VP.n40 VP.n39 0.189894
R69 VP.n40 VP.n0 0.189894
R70 VP.n44 VP.n0 0.189894
R71 VP VP.n44 0.0516364
R72 VDD1 VDD1.n0 72.6796
R73 VDD1.n3 VDD1.n2 72.5659
R74 VDD1.n3 VDD1.n1 72.5659
R75 VDD1.n5 VDD1.n4 71.8928
R76 VDD1.n5 VDD1.n3 42.5268
R77 VDD1.n4 VDD1.t1 2.40116
R78 VDD1.n4 VDD1.t0 2.40116
R79 VDD1.n0 VDD1.t2 2.40116
R80 VDD1.n0 VDD1.t3 2.40116
R81 VDD1.n2 VDD1.t5 2.40116
R82 VDD1.n2 VDD1.t4 2.40116
R83 VDD1.n1 VDD1.t7 2.40116
R84 VDD1.n1 VDD1.t6 2.40116
R85 VDD1 VDD1.n5 0.670759
R86 VTAIL.n594 VTAIL.n526 756.745
R87 VTAIL.n70 VTAIL.n2 756.745
R88 VTAIL.n144 VTAIL.n76 756.745
R89 VTAIL.n220 VTAIL.n152 756.745
R90 VTAIL.n520 VTAIL.n452 756.745
R91 VTAIL.n444 VTAIL.n376 756.745
R92 VTAIL.n370 VTAIL.n302 756.745
R93 VTAIL.n294 VTAIL.n226 756.745
R94 VTAIL.n551 VTAIL.n550 585
R95 VTAIL.n553 VTAIL.n552 585
R96 VTAIL.n546 VTAIL.n545 585
R97 VTAIL.n559 VTAIL.n558 585
R98 VTAIL.n561 VTAIL.n560 585
R99 VTAIL.n542 VTAIL.n541 585
R100 VTAIL.n568 VTAIL.n567 585
R101 VTAIL.n569 VTAIL.n540 585
R102 VTAIL.n571 VTAIL.n570 585
R103 VTAIL.n538 VTAIL.n537 585
R104 VTAIL.n577 VTAIL.n576 585
R105 VTAIL.n579 VTAIL.n578 585
R106 VTAIL.n534 VTAIL.n533 585
R107 VTAIL.n585 VTAIL.n584 585
R108 VTAIL.n587 VTAIL.n586 585
R109 VTAIL.n530 VTAIL.n529 585
R110 VTAIL.n593 VTAIL.n592 585
R111 VTAIL.n595 VTAIL.n594 585
R112 VTAIL.n27 VTAIL.n26 585
R113 VTAIL.n29 VTAIL.n28 585
R114 VTAIL.n22 VTAIL.n21 585
R115 VTAIL.n35 VTAIL.n34 585
R116 VTAIL.n37 VTAIL.n36 585
R117 VTAIL.n18 VTAIL.n17 585
R118 VTAIL.n44 VTAIL.n43 585
R119 VTAIL.n45 VTAIL.n16 585
R120 VTAIL.n47 VTAIL.n46 585
R121 VTAIL.n14 VTAIL.n13 585
R122 VTAIL.n53 VTAIL.n52 585
R123 VTAIL.n55 VTAIL.n54 585
R124 VTAIL.n10 VTAIL.n9 585
R125 VTAIL.n61 VTAIL.n60 585
R126 VTAIL.n63 VTAIL.n62 585
R127 VTAIL.n6 VTAIL.n5 585
R128 VTAIL.n69 VTAIL.n68 585
R129 VTAIL.n71 VTAIL.n70 585
R130 VTAIL.n101 VTAIL.n100 585
R131 VTAIL.n103 VTAIL.n102 585
R132 VTAIL.n96 VTAIL.n95 585
R133 VTAIL.n109 VTAIL.n108 585
R134 VTAIL.n111 VTAIL.n110 585
R135 VTAIL.n92 VTAIL.n91 585
R136 VTAIL.n118 VTAIL.n117 585
R137 VTAIL.n119 VTAIL.n90 585
R138 VTAIL.n121 VTAIL.n120 585
R139 VTAIL.n88 VTAIL.n87 585
R140 VTAIL.n127 VTAIL.n126 585
R141 VTAIL.n129 VTAIL.n128 585
R142 VTAIL.n84 VTAIL.n83 585
R143 VTAIL.n135 VTAIL.n134 585
R144 VTAIL.n137 VTAIL.n136 585
R145 VTAIL.n80 VTAIL.n79 585
R146 VTAIL.n143 VTAIL.n142 585
R147 VTAIL.n145 VTAIL.n144 585
R148 VTAIL.n177 VTAIL.n176 585
R149 VTAIL.n179 VTAIL.n178 585
R150 VTAIL.n172 VTAIL.n171 585
R151 VTAIL.n185 VTAIL.n184 585
R152 VTAIL.n187 VTAIL.n186 585
R153 VTAIL.n168 VTAIL.n167 585
R154 VTAIL.n194 VTAIL.n193 585
R155 VTAIL.n195 VTAIL.n166 585
R156 VTAIL.n197 VTAIL.n196 585
R157 VTAIL.n164 VTAIL.n163 585
R158 VTAIL.n203 VTAIL.n202 585
R159 VTAIL.n205 VTAIL.n204 585
R160 VTAIL.n160 VTAIL.n159 585
R161 VTAIL.n211 VTAIL.n210 585
R162 VTAIL.n213 VTAIL.n212 585
R163 VTAIL.n156 VTAIL.n155 585
R164 VTAIL.n219 VTAIL.n218 585
R165 VTAIL.n221 VTAIL.n220 585
R166 VTAIL.n521 VTAIL.n520 585
R167 VTAIL.n519 VTAIL.n518 585
R168 VTAIL.n456 VTAIL.n455 585
R169 VTAIL.n513 VTAIL.n512 585
R170 VTAIL.n511 VTAIL.n510 585
R171 VTAIL.n460 VTAIL.n459 585
R172 VTAIL.n505 VTAIL.n504 585
R173 VTAIL.n503 VTAIL.n502 585
R174 VTAIL.n464 VTAIL.n463 585
R175 VTAIL.n468 VTAIL.n466 585
R176 VTAIL.n497 VTAIL.n496 585
R177 VTAIL.n495 VTAIL.n494 585
R178 VTAIL.n470 VTAIL.n469 585
R179 VTAIL.n489 VTAIL.n488 585
R180 VTAIL.n487 VTAIL.n486 585
R181 VTAIL.n474 VTAIL.n473 585
R182 VTAIL.n481 VTAIL.n480 585
R183 VTAIL.n479 VTAIL.n478 585
R184 VTAIL.n445 VTAIL.n444 585
R185 VTAIL.n443 VTAIL.n442 585
R186 VTAIL.n380 VTAIL.n379 585
R187 VTAIL.n437 VTAIL.n436 585
R188 VTAIL.n435 VTAIL.n434 585
R189 VTAIL.n384 VTAIL.n383 585
R190 VTAIL.n429 VTAIL.n428 585
R191 VTAIL.n427 VTAIL.n426 585
R192 VTAIL.n388 VTAIL.n387 585
R193 VTAIL.n392 VTAIL.n390 585
R194 VTAIL.n421 VTAIL.n420 585
R195 VTAIL.n419 VTAIL.n418 585
R196 VTAIL.n394 VTAIL.n393 585
R197 VTAIL.n413 VTAIL.n412 585
R198 VTAIL.n411 VTAIL.n410 585
R199 VTAIL.n398 VTAIL.n397 585
R200 VTAIL.n405 VTAIL.n404 585
R201 VTAIL.n403 VTAIL.n402 585
R202 VTAIL.n371 VTAIL.n370 585
R203 VTAIL.n369 VTAIL.n368 585
R204 VTAIL.n306 VTAIL.n305 585
R205 VTAIL.n363 VTAIL.n362 585
R206 VTAIL.n361 VTAIL.n360 585
R207 VTAIL.n310 VTAIL.n309 585
R208 VTAIL.n355 VTAIL.n354 585
R209 VTAIL.n353 VTAIL.n352 585
R210 VTAIL.n314 VTAIL.n313 585
R211 VTAIL.n318 VTAIL.n316 585
R212 VTAIL.n347 VTAIL.n346 585
R213 VTAIL.n345 VTAIL.n344 585
R214 VTAIL.n320 VTAIL.n319 585
R215 VTAIL.n339 VTAIL.n338 585
R216 VTAIL.n337 VTAIL.n336 585
R217 VTAIL.n324 VTAIL.n323 585
R218 VTAIL.n331 VTAIL.n330 585
R219 VTAIL.n329 VTAIL.n328 585
R220 VTAIL.n295 VTAIL.n294 585
R221 VTAIL.n293 VTAIL.n292 585
R222 VTAIL.n230 VTAIL.n229 585
R223 VTAIL.n287 VTAIL.n286 585
R224 VTAIL.n285 VTAIL.n284 585
R225 VTAIL.n234 VTAIL.n233 585
R226 VTAIL.n279 VTAIL.n278 585
R227 VTAIL.n277 VTAIL.n276 585
R228 VTAIL.n238 VTAIL.n237 585
R229 VTAIL.n242 VTAIL.n240 585
R230 VTAIL.n271 VTAIL.n270 585
R231 VTAIL.n269 VTAIL.n268 585
R232 VTAIL.n244 VTAIL.n243 585
R233 VTAIL.n263 VTAIL.n262 585
R234 VTAIL.n261 VTAIL.n260 585
R235 VTAIL.n248 VTAIL.n247 585
R236 VTAIL.n255 VTAIL.n254 585
R237 VTAIL.n253 VTAIL.n252 585
R238 VTAIL.n549 VTAIL.t1 329.036
R239 VTAIL.n25 VTAIL.t0 329.036
R240 VTAIL.n99 VTAIL.t12 329.036
R241 VTAIL.n175 VTAIL.t15 329.036
R242 VTAIL.n477 VTAIL.t9 329.036
R243 VTAIL.n401 VTAIL.t13 329.036
R244 VTAIL.n327 VTAIL.t3 329.036
R245 VTAIL.n251 VTAIL.t6 329.036
R246 VTAIL.n552 VTAIL.n551 171.744
R247 VTAIL.n552 VTAIL.n545 171.744
R248 VTAIL.n559 VTAIL.n545 171.744
R249 VTAIL.n560 VTAIL.n559 171.744
R250 VTAIL.n560 VTAIL.n541 171.744
R251 VTAIL.n568 VTAIL.n541 171.744
R252 VTAIL.n569 VTAIL.n568 171.744
R253 VTAIL.n570 VTAIL.n569 171.744
R254 VTAIL.n570 VTAIL.n537 171.744
R255 VTAIL.n577 VTAIL.n537 171.744
R256 VTAIL.n578 VTAIL.n577 171.744
R257 VTAIL.n578 VTAIL.n533 171.744
R258 VTAIL.n585 VTAIL.n533 171.744
R259 VTAIL.n586 VTAIL.n585 171.744
R260 VTAIL.n586 VTAIL.n529 171.744
R261 VTAIL.n593 VTAIL.n529 171.744
R262 VTAIL.n594 VTAIL.n593 171.744
R263 VTAIL.n28 VTAIL.n27 171.744
R264 VTAIL.n28 VTAIL.n21 171.744
R265 VTAIL.n35 VTAIL.n21 171.744
R266 VTAIL.n36 VTAIL.n35 171.744
R267 VTAIL.n36 VTAIL.n17 171.744
R268 VTAIL.n44 VTAIL.n17 171.744
R269 VTAIL.n45 VTAIL.n44 171.744
R270 VTAIL.n46 VTAIL.n45 171.744
R271 VTAIL.n46 VTAIL.n13 171.744
R272 VTAIL.n53 VTAIL.n13 171.744
R273 VTAIL.n54 VTAIL.n53 171.744
R274 VTAIL.n54 VTAIL.n9 171.744
R275 VTAIL.n61 VTAIL.n9 171.744
R276 VTAIL.n62 VTAIL.n61 171.744
R277 VTAIL.n62 VTAIL.n5 171.744
R278 VTAIL.n69 VTAIL.n5 171.744
R279 VTAIL.n70 VTAIL.n69 171.744
R280 VTAIL.n102 VTAIL.n101 171.744
R281 VTAIL.n102 VTAIL.n95 171.744
R282 VTAIL.n109 VTAIL.n95 171.744
R283 VTAIL.n110 VTAIL.n109 171.744
R284 VTAIL.n110 VTAIL.n91 171.744
R285 VTAIL.n118 VTAIL.n91 171.744
R286 VTAIL.n119 VTAIL.n118 171.744
R287 VTAIL.n120 VTAIL.n119 171.744
R288 VTAIL.n120 VTAIL.n87 171.744
R289 VTAIL.n127 VTAIL.n87 171.744
R290 VTAIL.n128 VTAIL.n127 171.744
R291 VTAIL.n128 VTAIL.n83 171.744
R292 VTAIL.n135 VTAIL.n83 171.744
R293 VTAIL.n136 VTAIL.n135 171.744
R294 VTAIL.n136 VTAIL.n79 171.744
R295 VTAIL.n143 VTAIL.n79 171.744
R296 VTAIL.n144 VTAIL.n143 171.744
R297 VTAIL.n178 VTAIL.n177 171.744
R298 VTAIL.n178 VTAIL.n171 171.744
R299 VTAIL.n185 VTAIL.n171 171.744
R300 VTAIL.n186 VTAIL.n185 171.744
R301 VTAIL.n186 VTAIL.n167 171.744
R302 VTAIL.n194 VTAIL.n167 171.744
R303 VTAIL.n195 VTAIL.n194 171.744
R304 VTAIL.n196 VTAIL.n195 171.744
R305 VTAIL.n196 VTAIL.n163 171.744
R306 VTAIL.n203 VTAIL.n163 171.744
R307 VTAIL.n204 VTAIL.n203 171.744
R308 VTAIL.n204 VTAIL.n159 171.744
R309 VTAIL.n211 VTAIL.n159 171.744
R310 VTAIL.n212 VTAIL.n211 171.744
R311 VTAIL.n212 VTAIL.n155 171.744
R312 VTAIL.n219 VTAIL.n155 171.744
R313 VTAIL.n220 VTAIL.n219 171.744
R314 VTAIL.n520 VTAIL.n519 171.744
R315 VTAIL.n519 VTAIL.n455 171.744
R316 VTAIL.n512 VTAIL.n455 171.744
R317 VTAIL.n512 VTAIL.n511 171.744
R318 VTAIL.n511 VTAIL.n459 171.744
R319 VTAIL.n504 VTAIL.n459 171.744
R320 VTAIL.n504 VTAIL.n503 171.744
R321 VTAIL.n503 VTAIL.n463 171.744
R322 VTAIL.n468 VTAIL.n463 171.744
R323 VTAIL.n496 VTAIL.n468 171.744
R324 VTAIL.n496 VTAIL.n495 171.744
R325 VTAIL.n495 VTAIL.n469 171.744
R326 VTAIL.n488 VTAIL.n469 171.744
R327 VTAIL.n488 VTAIL.n487 171.744
R328 VTAIL.n487 VTAIL.n473 171.744
R329 VTAIL.n480 VTAIL.n473 171.744
R330 VTAIL.n480 VTAIL.n479 171.744
R331 VTAIL.n444 VTAIL.n443 171.744
R332 VTAIL.n443 VTAIL.n379 171.744
R333 VTAIL.n436 VTAIL.n379 171.744
R334 VTAIL.n436 VTAIL.n435 171.744
R335 VTAIL.n435 VTAIL.n383 171.744
R336 VTAIL.n428 VTAIL.n383 171.744
R337 VTAIL.n428 VTAIL.n427 171.744
R338 VTAIL.n427 VTAIL.n387 171.744
R339 VTAIL.n392 VTAIL.n387 171.744
R340 VTAIL.n420 VTAIL.n392 171.744
R341 VTAIL.n420 VTAIL.n419 171.744
R342 VTAIL.n419 VTAIL.n393 171.744
R343 VTAIL.n412 VTAIL.n393 171.744
R344 VTAIL.n412 VTAIL.n411 171.744
R345 VTAIL.n411 VTAIL.n397 171.744
R346 VTAIL.n404 VTAIL.n397 171.744
R347 VTAIL.n404 VTAIL.n403 171.744
R348 VTAIL.n370 VTAIL.n369 171.744
R349 VTAIL.n369 VTAIL.n305 171.744
R350 VTAIL.n362 VTAIL.n305 171.744
R351 VTAIL.n362 VTAIL.n361 171.744
R352 VTAIL.n361 VTAIL.n309 171.744
R353 VTAIL.n354 VTAIL.n309 171.744
R354 VTAIL.n354 VTAIL.n353 171.744
R355 VTAIL.n353 VTAIL.n313 171.744
R356 VTAIL.n318 VTAIL.n313 171.744
R357 VTAIL.n346 VTAIL.n318 171.744
R358 VTAIL.n346 VTAIL.n345 171.744
R359 VTAIL.n345 VTAIL.n319 171.744
R360 VTAIL.n338 VTAIL.n319 171.744
R361 VTAIL.n338 VTAIL.n337 171.744
R362 VTAIL.n337 VTAIL.n323 171.744
R363 VTAIL.n330 VTAIL.n323 171.744
R364 VTAIL.n330 VTAIL.n329 171.744
R365 VTAIL.n294 VTAIL.n293 171.744
R366 VTAIL.n293 VTAIL.n229 171.744
R367 VTAIL.n286 VTAIL.n229 171.744
R368 VTAIL.n286 VTAIL.n285 171.744
R369 VTAIL.n285 VTAIL.n233 171.744
R370 VTAIL.n278 VTAIL.n233 171.744
R371 VTAIL.n278 VTAIL.n277 171.744
R372 VTAIL.n277 VTAIL.n237 171.744
R373 VTAIL.n242 VTAIL.n237 171.744
R374 VTAIL.n270 VTAIL.n242 171.744
R375 VTAIL.n270 VTAIL.n269 171.744
R376 VTAIL.n269 VTAIL.n243 171.744
R377 VTAIL.n262 VTAIL.n243 171.744
R378 VTAIL.n262 VTAIL.n261 171.744
R379 VTAIL.n261 VTAIL.n247 171.744
R380 VTAIL.n254 VTAIL.n247 171.744
R381 VTAIL.n254 VTAIL.n253 171.744
R382 VTAIL.n551 VTAIL.t1 85.8723
R383 VTAIL.n27 VTAIL.t0 85.8723
R384 VTAIL.n101 VTAIL.t12 85.8723
R385 VTAIL.n177 VTAIL.t15 85.8723
R386 VTAIL.n479 VTAIL.t9 85.8723
R387 VTAIL.n403 VTAIL.t13 85.8723
R388 VTAIL.n329 VTAIL.t3 85.8723
R389 VTAIL.n253 VTAIL.t6 85.8723
R390 VTAIL.n451 VTAIL.n450 55.2142
R391 VTAIL.n301 VTAIL.n300 55.2142
R392 VTAIL.n1 VTAIL.n0 55.214
R393 VTAIL.n151 VTAIL.n150 55.214
R394 VTAIL.n599 VTAIL.n598 31.7975
R395 VTAIL.n75 VTAIL.n74 31.7975
R396 VTAIL.n149 VTAIL.n148 31.7975
R397 VTAIL.n225 VTAIL.n224 31.7975
R398 VTAIL.n525 VTAIL.n524 31.7975
R399 VTAIL.n449 VTAIL.n448 31.7975
R400 VTAIL.n375 VTAIL.n374 31.7975
R401 VTAIL.n299 VTAIL.n298 31.7975
R402 VTAIL.n599 VTAIL.n525 25.4962
R403 VTAIL.n299 VTAIL.n225 25.4962
R404 VTAIL.n571 VTAIL.n538 13.1884
R405 VTAIL.n47 VTAIL.n14 13.1884
R406 VTAIL.n121 VTAIL.n88 13.1884
R407 VTAIL.n197 VTAIL.n164 13.1884
R408 VTAIL.n466 VTAIL.n464 13.1884
R409 VTAIL.n390 VTAIL.n388 13.1884
R410 VTAIL.n316 VTAIL.n314 13.1884
R411 VTAIL.n240 VTAIL.n238 13.1884
R412 VTAIL.n572 VTAIL.n540 12.8005
R413 VTAIL.n576 VTAIL.n575 12.8005
R414 VTAIL.n48 VTAIL.n16 12.8005
R415 VTAIL.n52 VTAIL.n51 12.8005
R416 VTAIL.n122 VTAIL.n90 12.8005
R417 VTAIL.n126 VTAIL.n125 12.8005
R418 VTAIL.n198 VTAIL.n166 12.8005
R419 VTAIL.n202 VTAIL.n201 12.8005
R420 VTAIL.n502 VTAIL.n501 12.8005
R421 VTAIL.n498 VTAIL.n497 12.8005
R422 VTAIL.n426 VTAIL.n425 12.8005
R423 VTAIL.n422 VTAIL.n421 12.8005
R424 VTAIL.n352 VTAIL.n351 12.8005
R425 VTAIL.n348 VTAIL.n347 12.8005
R426 VTAIL.n276 VTAIL.n275 12.8005
R427 VTAIL.n272 VTAIL.n271 12.8005
R428 VTAIL.n567 VTAIL.n566 12.0247
R429 VTAIL.n579 VTAIL.n536 12.0247
R430 VTAIL.n43 VTAIL.n42 12.0247
R431 VTAIL.n55 VTAIL.n12 12.0247
R432 VTAIL.n117 VTAIL.n116 12.0247
R433 VTAIL.n129 VTAIL.n86 12.0247
R434 VTAIL.n193 VTAIL.n192 12.0247
R435 VTAIL.n205 VTAIL.n162 12.0247
R436 VTAIL.n505 VTAIL.n462 12.0247
R437 VTAIL.n494 VTAIL.n467 12.0247
R438 VTAIL.n429 VTAIL.n386 12.0247
R439 VTAIL.n418 VTAIL.n391 12.0247
R440 VTAIL.n355 VTAIL.n312 12.0247
R441 VTAIL.n344 VTAIL.n317 12.0247
R442 VTAIL.n279 VTAIL.n236 12.0247
R443 VTAIL.n268 VTAIL.n241 12.0247
R444 VTAIL.n565 VTAIL.n542 11.249
R445 VTAIL.n580 VTAIL.n534 11.249
R446 VTAIL.n41 VTAIL.n18 11.249
R447 VTAIL.n56 VTAIL.n10 11.249
R448 VTAIL.n115 VTAIL.n92 11.249
R449 VTAIL.n130 VTAIL.n84 11.249
R450 VTAIL.n191 VTAIL.n168 11.249
R451 VTAIL.n206 VTAIL.n160 11.249
R452 VTAIL.n506 VTAIL.n460 11.249
R453 VTAIL.n493 VTAIL.n470 11.249
R454 VTAIL.n430 VTAIL.n384 11.249
R455 VTAIL.n417 VTAIL.n394 11.249
R456 VTAIL.n356 VTAIL.n310 11.249
R457 VTAIL.n343 VTAIL.n320 11.249
R458 VTAIL.n280 VTAIL.n234 11.249
R459 VTAIL.n267 VTAIL.n244 11.249
R460 VTAIL.n550 VTAIL.n549 10.7239
R461 VTAIL.n26 VTAIL.n25 10.7239
R462 VTAIL.n100 VTAIL.n99 10.7239
R463 VTAIL.n176 VTAIL.n175 10.7239
R464 VTAIL.n478 VTAIL.n477 10.7239
R465 VTAIL.n402 VTAIL.n401 10.7239
R466 VTAIL.n328 VTAIL.n327 10.7239
R467 VTAIL.n252 VTAIL.n251 10.7239
R468 VTAIL.n562 VTAIL.n561 10.4732
R469 VTAIL.n584 VTAIL.n583 10.4732
R470 VTAIL.n38 VTAIL.n37 10.4732
R471 VTAIL.n60 VTAIL.n59 10.4732
R472 VTAIL.n112 VTAIL.n111 10.4732
R473 VTAIL.n134 VTAIL.n133 10.4732
R474 VTAIL.n188 VTAIL.n187 10.4732
R475 VTAIL.n210 VTAIL.n209 10.4732
R476 VTAIL.n510 VTAIL.n509 10.4732
R477 VTAIL.n490 VTAIL.n489 10.4732
R478 VTAIL.n434 VTAIL.n433 10.4732
R479 VTAIL.n414 VTAIL.n413 10.4732
R480 VTAIL.n360 VTAIL.n359 10.4732
R481 VTAIL.n340 VTAIL.n339 10.4732
R482 VTAIL.n284 VTAIL.n283 10.4732
R483 VTAIL.n264 VTAIL.n263 10.4732
R484 VTAIL.n558 VTAIL.n544 9.69747
R485 VTAIL.n587 VTAIL.n532 9.69747
R486 VTAIL.n34 VTAIL.n20 9.69747
R487 VTAIL.n63 VTAIL.n8 9.69747
R488 VTAIL.n108 VTAIL.n94 9.69747
R489 VTAIL.n137 VTAIL.n82 9.69747
R490 VTAIL.n184 VTAIL.n170 9.69747
R491 VTAIL.n213 VTAIL.n158 9.69747
R492 VTAIL.n513 VTAIL.n458 9.69747
R493 VTAIL.n486 VTAIL.n472 9.69747
R494 VTAIL.n437 VTAIL.n382 9.69747
R495 VTAIL.n410 VTAIL.n396 9.69747
R496 VTAIL.n363 VTAIL.n308 9.69747
R497 VTAIL.n336 VTAIL.n322 9.69747
R498 VTAIL.n287 VTAIL.n232 9.69747
R499 VTAIL.n260 VTAIL.n246 9.69747
R500 VTAIL.n598 VTAIL.n597 9.45567
R501 VTAIL.n74 VTAIL.n73 9.45567
R502 VTAIL.n148 VTAIL.n147 9.45567
R503 VTAIL.n224 VTAIL.n223 9.45567
R504 VTAIL.n524 VTAIL.n523 9.45567
R505 VTAIL.n448 VTAIL.n447 9.45567
R506 VTAIL.n374 VTAIL.n373 9.45567
R507 VTAIL.n298 VTAIL.n297 9.45567
R508 VTAIL.n597 VTAIL.n596 9.3005
R509 VTAIL.n591 VTAIL.n590 9.3005
R510 VTAIL.n589 VTAIL.n588 9.3005
R511 VTAIL.n532 VTAIL.n531 9.3005
R512 VTAIL.n583 VTAIL.n582 9.3005
R513 VTAIL.n581 VTAIL.n580 9.3005
R514 VTAIL.n536 VTAIL.n535 9.3005
R515 VTAIL.n575 VTAIL.n574 9.3005
R516 VTAIL.n548 VTAIL.n547 9.3005
R517 VTAIL.n555 VTAIL.n554 9.3005
R518 VTAIL.n557 VTAIL.n556 9.3005
R519 VTAIL.n544 VTAIL.n543 9.3005
R520 VTAIL.n563 VTAIL.n562 9.3005
R521 VTAIL.n565 VTAIL.n564 9.3005
R522 VTAIL.n566 VTAIL.n539 9.3005
R523 VTAIL.n573 VTAIL.n572 9.3005
R524 VTAIL.n528 VTAIL.n527 9.3005
R525 VTAIL.n73 VTAIL.n72 9.3005
R526 VTAIL.n67 VTAIL.n66 9.3005
R527 VTAIL.n65 VTAIL.n64 9.3005
R528 VTAIL.n8 VTAIL.n7 9.3005
R529 VTAIL.n59 VTAIL.n58 9.3005
R530 VTAIL.n57 VTAIL.n56 9.3005
R531 VTAIL.n12 VTAIL.n11 9.3005
R532 VTAIL.n51 VTAIL.n50 9.3005
R533 VTAIL.n24 VTAIL.n23 9.3005
R534 VTAIL.n31 VTAIL.n30 9.3005
R535 VTAIL.n33 VTAIL.n32 9.3005
R536 VTAIL.n20 VTAIL.n19 9.3005
R537 VTAIL.n39 VTAIL.n38 9.3005
R538 VTAIL.n41 VTAIL.n40 9.3005
R539 VTAIL.n42 VTAIL.n15 9.3005
R540 VTAIL.n49 VTAIL.n48 9.3005
R541 VTAIL.n4 VTAIL.n3 9.3005
R542 VTAIL.n147 VTAIL.n146 9.3005
R543 VTAIL.n141 VTAIL.n140 9.3005
R544 VTAIL.n139 VTAIL.n138 9.3005
R545 VTAIL.n82 VTAIL.n81 9.3005
R546 VTAIL.n133 VTAIL.n132 9.3005
R547 VTAIL.n131 VTAIL.n130 9.3005
R548 VTAIL.n86 VTAIL.n85 9.3005
R549 VTAIL.n125 VTAIL.n124 9.3005
R550 VTAIL.n98 VTAIL.n97 9.3005
R551 VTAIL.n105 VTAIL.n104 9.3005
R552 VTAIL.n107 VTAIL.n106 9.3005
R553 VTAIL.n94 VTAIL.n93 9.3005
R554 VTAIL.n113 VTAIL.n112 9.3005
R555 VTAIL.n115 VTAIL.n114 9.3005
R556 VTAIL.n116 VTAIL.n89 9.3005
R557 VTAIL.n123 VTAIL.n122 9.3005
R558 VTAIL.n78 VTAIL.n77 9.3005
R559 VTAIL.n223 VTAIL.n222 9.3005
R560 VTAIL.n217 VTAIL.n216 9.3005
R561 VTAIL.n215 VTAIL.n214 9.3005
R562 VTAIL.n158 VTAIL.n157 9.3005
R563 VTAIL.n209 VTAIL.n208 9.3005
R564 VTAIL.n207 VTAIL.n206 9.3005
R565 VTAIL.n162 VTAIL.n161 9.3005
R566 VTAIL.n201 VTAIL.n200 9.3005
R567 VTAIL.n174 VTAIL.n173 9.3005
R568 VTAIL.n181 VTAIL.n180 9.3005
R569 VTAIL.n183 VTAIL.n182 9.3005
R570 VTAIL.n170 VTAIL.n169 9.3005
R571 VTAIL.n189 VTAIL.n188 9.3005
R572 VTAIL.n191 VTAIL.n190 9.3005
R573 VTAIL.n192 VTAIL.n165 9.3005
R574 VTAIL.n199 VTAIL.n198 9.3005
R575 VTAIL.n154 VTAIL.n153 9.3005
R576 VTAIL.n476 VTAIL.n475 9.3005
R577 VTAIL.n483 VTAIL.n482 9.3005
R578 VTAIL.n485 VTAIL.n484 9.3005
R579 VTAIL.n472 VTAIL.n471 9.3005
R580 VTAIL.n491 VTAIL.n490 9.3005
R581 VTAIL.n493 VTAIL.n492 9.3005
R582 VTAIL.n467 VTAIL.n465 9.3005
R583 VTAIL.n499 VTAIL.n498 9.3005
R584 VTAIL.n523 VTAIL.n522 9.3005
R585 VTAIL.n454 VTAIL.n453 9.3005
R586 VTAIL.n517 VTAIL.n516 9.3005
R587 VTAIL.n515 VTAIL.n514 9.3005
R588 VTAIL.n458 VTAIL.n457 9.3005
R589 VTAIL.n509 VTAIL.n508 9.3005
R590 VTAIL.n507 VTAIL.n506 9.3005
R591 VTAIL.n462 VTAIL.n461 9.3005
R592 VTAIL.n501 VTAIL.n500 9.3005
R593 VTAIL.n400 VTAIL.n399 9.3005
R594 VTAIL.n407 VTAIL.n406 9.3005
R595 VTAIL.n409 VTAIL.n408 9.3005
R596 VTAIL.n396 VTAIL.n395 9.3005
R597 VTAIL.n415 VTAIL.n414 9.3005
R598 VTAIL.n417 VTAIL.n416 9.3005
R599 VTAIL.n391 VTAIL.n389 9.3005
R600 VTAIL.n423 VTAIL.n422 9.3005
R601 VTAIL.n447 VTAIL.n446 9.3005
R602 VTAIL.n378 VTAIL.n377 9.3005
R603 VTAIL.n441 VTAIL.n440 9.3005
R604 VTAIL.n439 VTAIL.n438 9.3005
R605 VTAIL.n382 VTAIL.n381 9.3005
R606 VTAIL.n433 VTAIL.n432 9.3005
R607 VTAIL.n431 VTAIL.n430 9.3005
R608 VTAIL.n386 VTAIL.n385 9.3005
R609 VTAIL.n425 VTAIL.n424 9.3005
R610 VTAIL.n326 VTAIL.n325 9.3005
R611 VTAIL.n333 VTAIL.n332 9.3005
R612 VTAIL.n335 VTAIL.n334 9.3005
R613 VTAIL.n322 VTAIL.n321 9.3005
R614 VTAIL.n341 VTAIL.n340 9.3005
R615 VTAIL.n343 VTAIL.n342 9.3005
R616 VTAIL.n317 VTAIL.n315 9.3005
R617 VTAIL.n349 VTAIL.n348 9.3005
R618 VTAIL.n373 VTAIL.n372 9.3005
R619 VTAIL.n304 VTAIL.n303 9.3005
R620 VTAIL.n367 VTAIL.n366 9.3005
R621 VTAIL.n365 VTAIL.n364 9.3005
R622 VTAIL.n308 VTAIL.n307 9.3005
R623 VTAIL.n359 VTAIL.n358 9.3005
R624 VTAIL.n357 VTAIL.n356 9.3005
R625 VTAIL.n312 VTAIL.n311 9.3005
R626 VTAIL.n351 VTAIL.n350 9.3005
R627 VTAIL.n250 VTAIL.n249 9.3005
R628 VTAIL.n257 VTAIL.n256 9.3005
R629 VTAIL.n259 VTAIL.n258 9.3005
R630 VTAIL.n246 VTAIL.n245 9.3005
R631 VTAIL.n265 VTAIL.n264 9.3005
R632 VTAIL.n267 VTAIL.n266 9.3005
R633 VTAIL.n241 VTAIL.n239 9.3005
R634 VTAIL.n273 VTAIL.n272 9.3005
R635 VTAIL.n297 VTAIL.n296 9.3005
R636 VTAIL.n228 VTAIL.n227 9.3005
R637 VTAIL.n291 VTAIL.n290 9.3005
R638 VTAIL.n289 VTAIL.n288 9.3005
R639 VTAIL.n232 VTAIL.n231 9.3005
R640 VTAIL.n283 VTAIL.n282 9.3005
R641 VTAIL.n281 VTAIL.n280 9.3005
R642 VTAIL.n236 VTAIL.n235 9.3005
R643 VTAIL.n275 VTAIL.n274 9.3005
R644 VTAIL.n557 VTAIL.n546 8.92171
R645 VTAIL.n588 VTAIL.n530 8.92171
R646 VTAIL.n33 VTAIL.n22 8.92171
R647 VTAIL.n64 VTAIL.n6 8.92171
R648 VTAIL.n107 VTAIL.n96 8.92171
R649 VTAIL.n138 VTAIL.n80 8.92171
R650 VTAIL.n183 VTAIL.n172 8.92171
R651 VTAIL.n214 VTAIL.n156 8.92171
R652 VTAIL.n514 VTAIL.n456 8.92171
R653 VTAIL.n485 VTAIL.n474 8.92171
R654 VTAIL.n438 VTAIL.n380 8.92171
R655 VTAIL.n409 VTAIL.n398 8.92171
R656 VTAIL.n364 VTAIL.n306 8.92171
R657 VTAIL.n335 VTAIL.n324 8.92171
R658 VTAIL.n288 VTAIL.n230 8.92171
R659 VTAIL.n259 VTAIL.n248 8.92171
R660 VTAIL.n554 VTAIL.n553 8.14595
R661 VTAIL.n592 VTAIL.n591 8.14595
R662 VTAIL.n30 VTAIL.n29 8.14595
R663 VTAIL.n68 VTAIL.n67 8.14595
R664 VTAIL.n104 VTAIL.n103 8.14595
R665 VTAIL.n142 VTAIL.n141 8.14595
R666 VTAIL.n180 VTAIL.n179 8.14595
R667 VTAIL.n218 VTAIL.n217 8.14595
R668 VTAIL.n518 VTAIL.n517 8.14595
R669 VTAIL.n482 VTAIL.n481 8.14595
R670 VTAIL.n442 VTAIL.n441 8.14595
R671 VTAIL.n406 VTAIL.n405 8.14595
R672 VTAIL.n368 VTAIL.n367 8.14595
R673 VTAIL.n332 VTAIL.n331 8.14595
R674 VTAIL.n292 VTAIL.n291 8.14595
R675 VTAIL.n256 VTAIL.n255 8.14595
R676 VTAIL.n550 VTAIL.n548 7.3702
R677 VTAIL.n595 VTAIL.n528 7.3702
R678 VTAIL.n598 VTAIL.n526 7.3702
R679 VTAIL.n26 VTAIL.n24 7.3702
R680 VTAIL.n71 VTAIL.n4 7.3702
R681 VTAIL.n74 VTAIL.n2 7.3702
R682 VTAIL.n100 VTAIL.n98 7.3702
R683 VTAIL.n145 VTAIL.n78 7.3702
R684 VTAIL.n148 VTAIL.n76 7.3702
R685 VTAIL.n176 VTAIL.n174 7.3702
R686 VTAIL.n221 VTAIL.n154 7.3702
R687 VTAIL.n224 VTAIL.n152 7.3702
R688 VTAIL.n524 VTAIL.n452 7.3702
R689 VTAIL.n521 VTAIL.n454 7.3702
R690 VTAIL.n478 VTAIL.n476 7.3702
R691 VTAIL.n448 VTAIL.n376 7.3702
R692 VTAIL.n445 VTAIL.n378 7.3702
R693 VTAIL.n402 VTAIL.n400 7.3702
R694 VTAIL.n374 VTAIL.n302 7.3702
R695 VTAIL.n371 VTAIL.n304 7.3702
R696 VTAIL.n328 VTAIL.n326 7.3702
R697 VTAIL.n298 VTAIL.n226 7.3702
R698 VTAIL.n295 VTAIL.n228 7.3702
R699 VTAIL.n252 VTAIL.n250 7.3702
R700 VTAIL.n596 VTAIL.n595 6.59444
R701 VTAIL.n596 VTAIL.n526 6.59444
R702 VTAIL.n72 VTAIL.n71 6.59444
R703 VTAIL.n72 VTAIL.n2 6.59444
R704 VTAIL.n146 VTAIL.n145 6.59444
R705 VTAIL.n146 VTAIL.n76 6.59444
R706 VTAIL.n222 VTAIL.n221 6.59444
R707 VTAIL.n222 VTAIL.n152 6.59444
R708 VTAIL.n522 VTAIL.n452 6.59444
R709 VTAIL.n522 VTAIL.n521 6.59444
R710 VTAIL.n446 VTAIL.n376 6.59444
R711 VTAIL.n446 VTAIL.n445 6.59444
R712 VTAIL.n372 VTAIL.n302 6.59444
R713 VTAIL.n372 VTAIL.n371 6.59444
R714 VTAIL.n296 VTAIL.n226 6.59444
R715 VTAIL.n296 VTAIL.n295 6.59444
R716 VTAIL.n553 VTAIL.n548 5.81868
R717 VTAIL.n592 VTAIL.n528 5.81868
R718 VTAIL.n29 VTAIL.n24 5.81868
R719 VTAIL.n68 VTAIL.n4 5.81868
R720 VTAIL.n103 VTAIL.n98 5.81868
R721 VTAIL.n142 VTAIL.n78 5.81868
R722 VTAIL.n179 VTAIL.n174 5.81868
R723 VTAIL.n218 VTAIL.n154 5.81868
R724 VTAIL.n518 VTAIL.n454 5.81868
R725 VTAIL.n481 VTAIL.n476 5.81868
R726 VTAIL.n442 VTAIL.n378 5.81868
R727 VTAIL.n405 VTAIL.n400 5.81868
R728 VTAIL.n368 VTAIL.n304 5.81868
R729 VTAIL.n331 VTAIL.n326 5.81868
R730 VTAIL.n292 VTAIL.n228 5.81868
R731 VTAIL.n255 VTAIL.n250 5.81868
R732 VTAIL.n554 VTAIL.n546 5.04292
R733 VTAIL.n591 VTAIL.n530 5.04292
R734 VTAIL.n30 VTAIL.n22 5.04292
R735 VTAIL.n67 VTAIL.n6 5.04292
R736 VTAIL.n104 VTAIL.n96 5.04292
R737 VTAIL.n141 VTAIL.n80 5.04292
R738 VTAIL.n180 VTAIL.n172 5.04292
R739 VTAIL.n217 VTAIL.n156 5.04292
R740 VTAIL.n517 VTAIL.n456 5.04292
R741 VTAIL.n482 VTAIL.n474 5.04292
R742 VTAIL.n441 VTAIL.n380 5.04292
R743 VTAIL.n406 VTAIL.n398 5.04292
R744 VTAIL.n367 VTAIL.n306 5.04292
R745 VTAIL.n332 VTAIL.n324 5.04292
R746 VTAIL.n291 VTAIL.n230 5.04292
R747 VTAIL.n256 VTAIL.n248 5.04292
R748 VTAIL.n558 VTAIL.n557 4.26717
R749 VTAIL.n588 VTAIL.n587 4.26717
R750 VTAIL.n34 VTAIL.n33 4.26717
R751 VTAIL.n64 VTAIL.n63 4.26717
R752 VTAIL.n108 VTAIL.n107 4.26717
R753 VTAIL.n138 VTAIL.n137 4.26717
R754 VTAIL.n184 VTAIL.n183 4.26717
R755 VTAIL.n214 VTAIL.n213 4.26717
R756 VTAIL.n514 VTAIL.n513 4.26717
R757 VTAIL.n486 VTAIL.n485 4.26717
R758 VTAIL.n438 VTAIL.n437 4.26717
R759 VTAIL.n410 VTAIL.n409 4.26717
R760 VTAIL.n364 VTAIL.n363 4.26717
R761 VTAIL.n336 VTAIL.n335 4.26717
R762 VTAIL.n288 VTAIL.n287 4.26717
R763 VTAIL.n260 VTAIL.n259 4.26717
R764 VTAIL.n561 VTAIL.n544 3.49141
R765 VTAIL.n584 VTAIL.n532 3.49141
R766 VTAIL.n37 VTAIL.n20 3.49141
R767 VTAIL.n60 VTAIL.n8 3.49141
R768 VTAIL.n111 VTAIL.n94 3.49141
R769 VTAIL.n134 VTAIL.n82 3.49141
R770 VTAIL.n187 VTAIL.n170 3.49141
R771 VTAIL.n210 VTAIL.n158 3.49141
R772 VTAIL.n510 VTAIL.n458 3.49141
R773 VTAIL.n489 VTAIL.n472 3.49141
R774 VTAIL.n434 VTAIL.n382 3.49141
R775 VTAIL.n413 VTAIL.n396 3.49141
R776 VTAIL.n360 VTAIL.n308 3.49141
R777 VTAIL.n339 VTAIL.n322 3.49141
R778 VTAIL.n284 VTAIL.n232 3.49141
R779 VTAIL.n263 VTAIL.n246 3.49141
R780 VTAIL.n562 VTAIL.n542 2.71565
R781 VTAIL.n583 VTAIL.n534 2.71565
R782 VTAIL.n38 VTAIL.n18 2.71565
R783 VTAIL.n59 VTAIL.n10 2.71565
R784 VTAIL.n112 VTAIL.n92 2.71565
R785 VTAIL.n133 VTAIL.n84 2.71565
R786 VTAIL.n188 VTAIL.n168 2.71565
R787 VTAIL.n209 VTAIL.n160 2.71565
R788 VTAIL.n509 VTAIL.n460 2.71565
R789 VTAIL.n490 VTAIL.n470 2.71565
R790 VTAIL.n433 VTAIL.n384 2.71565
R791 VTAIL.n414 VTAIL.n394 2.71565
R792 VTAIL.n359 VTAIL.n310 2.71565
R793 VTAIL.n340 VTAIL.n320 2.71565
R794 VTAIL.n283 VTAIL.n234 2.71565
R795 VTAIL.n264 VTAIL.n244 2.71565
R796 VTAIL.n549 VTAIL.n547 2.41282
R797 VTAIL.n25 VTAIL.n23 2.41282
R798 VTAIL.n99 VTAIL.n97 2.41282
R799 VTAIL.n175 VTAIL.n173 2.41282
R800 VTAIL.n477 VTAIL.n475 2.41282
R801 VTAIL.n401 VTAIL.n399 2.41282
R802 VTAIL.n327 VTAIL.n325 2.41282
R803 VTAIL.n251 VTAIL.n249 2.41282
R804 VTAIL.n0 VTAIL.t2 2.40116
R805 VTAIL.n0 VTAIL.t5 2.40116
R806 VTAIL.n150 VTAIL.t11 2.40116
R807 VTAIL.n150 VTAIL.t10 2.40116
R808 VTAIL.n450 VTAIL.t14 2.40116
R809 VTAIL.n450 VTAIL.t8 2.40116
R810 VTAIL.n300 VTAIL.t7 2.40116
R811 VTAIL.n300 VTAIL.t4 2.40116
R812 VTAIL.n567 VTAIL.n565 1.93989
R813 VTAIL.n580 VTAIL.n579 1.93989
R814 VTAIL.n43 VTAIL.n41 1.93989
R815 VTAIL.n56 VTAIL.n55 1.93989
R816 VTAIL.n117 VTAIL.n115 1.93989
R817 VTAIL.n130 VTAIL.n129 1.93989
R818 VTAIL.n193 VTAIL.n191 1.93989
R819 VTAIL.n206 VTAIL.n205 1.93989
R820 VTAIL.n506 VTAIL.n505 1.93989
R821 VTAIL.n494 VTAIL.n493 1.93989
R822 VTAIL.n430 VTAIL.n429 1.93989
R823 VTAIL.n418 VTAIL.n417 1.93989
R824 VTAIL.n356 VTAIL.n355 1.93989
R825 VTAIL.n344 VTAIL.n343 1.93989
R826 VTAIL.n280 VTAIL.n279 1.93989
R827 VTAIL.n268 VTAIL.n267 1.93989
R828 VTAIL.n301 VTAIL.n299 1.4574
R829 VTAIL.n375 VTAIL.n301 1.4574
R830 VTAIL.n451 VTAIL.n449 1.4574
R831 VTAIL.n525 VTAIL.n451 1.4574
R832 VTAIL.n225 VTAIL.n151 1.4574
R833 VTAIL.n151 VTAIL.n149 1.4574
R834 VTAIL.n75 VTAIL.n1 1.4574
R835 VTAIL VTAIL.n599 1.39921
R836 VTAIL.n566 VTAIL.n540 1.16414
R837 VTAIL.n576 VTAIL.n536 1.16414
R838 VTAIL.n42 VTAIL.n16 1.16414
R839 VTAIL.n52 VTAIL.n12 1.16414
R840 VTAIL.n116 VTAIL.n90 1.16414
R841 VTAIL.n126 VTAIL.n86 1.16414
R842 VTAIL.n192 VTAIL.n166 1.16414
R843 VTAIL.n202 VTAIL.n162 1.16414
R844 VTAIL.n502 VTAIL.n462 1.16414
R845 VTAIL.n497 VTAIL.n467 1.16414
R846 VTAIL.n426 VTAIL.n386 1.16414
R847 VTAIL.n421 VTAIL.n391 1.16414
R848 VTAIL.n352 VTAIL.n312 1.16414
R849 VTAIL.n347 VTAIL.n317 1.16414
R850 VTAIL.n276 VTAIL.n236 1.16414
R851 VTAIL.n271 VTAIL.n241 1.16414
R852 VTAIL.n449 VTAIL.n375 0.470328
R853 VTAIL.n149 VTAIL.n75 0.470328
R854 VTAIL.n572 VTAIL.n571 0.388379
R855 VTAIL.n575 VTAIL.n538 0.388379
R856 VTAIL.n48 VTAIL.n47 0.388379
R857 VTAIL.n51 VTAIL.n14 0.388379
R858 VTAIL.n122 VTAIL.n121 0.388379
R859 VTAIL.n125 VTAIL.n88 0.388379
R860 VTAIL.n198 VTAIL.n197 0.388379
R861 VTAIL.n201 VTAIL.n164 0.388379
R862 VTAIL.n501 VTAIL.n464 0.388379
R863 VTAIL.n498 VTAIL.n466 0.388379
R864 VTAIL.n425 VTAIL.n388 0.388379
R865 VTAIL.n422 VTAIL.n390 0.388379
R866 VTAIL.n351 VTAIL.n314 0.388379
R867 VTAIL.n348 VTAIL.n316 0.388379
R868 VTAIL.n275 VTAIL.n238 0.388379
R869 VTAIL.n272 VTAIL.n240 0.388379
R870 VTAIL.n555 VTAIL.n547 0.155672
R871 VTAIL.n556 VTAIL.n555 0.155672
R872 VTAIL.n556 VTAIL.n543 0.155672
R873 VTAIL.n563 VTAIL.n543 0.155672
R874 VTAIL.n564 VTAIL.n563 0.155672
R875 VTAIL.n564 VTAIL.n539 0.155672
R876 VTAIL.n573 VTAIL.n539 0.155672
R877 VTAIL.n574 VTAIL.n573 0.155672
R878 VTAIL.n574 VTAIL.n535 0.155672
R879 VTAIL.n581 VTAIL.n535 0.155672
R880 VTAIL.n582 VTAIL.n581 0.155672
R881 VTAIL.n582 VTAIL.n531 0.155672
R882 VTAIL.n589 VTAIL.n531 0.155672
R883 VTAIL.n590 VTAIL.n589 0.155672
R884 VTAIL.n590 VTAIL.n527 0.155672
R885 VTAIL.n597 VTAIL.n527 0.155672
R886 VTAIL.n31 VTAIL.n23 0.155672
R887 VTAIL.n32 VTAIL.n31 0.155672
R888 VTAIL.n32 VTAIL.n19 0.155672
R889 VTAIL.n39 VTAIL.n19 0.155672
R890 VTAIL.n40 VTAIL.n39 0.155672
R891 VTAIL.n40 VTAIL.n15 0.155672
R892 VTAIL.n49 VTAIL.n15 0.155672
R893 VTAIL.n50 VTAIL.n49 0.155672
R894 VTAIL.n50 VTAIL.n11 0.155672
R895 VTAIL.n57 VTAIL.n11 0.155672
R896 VTAIL.n58 VTAIL.n57 0.155672
R897 VTAIL.n58 VTAIL.n7 0.155672
R898 VTAIL.n65 VTAIL.n7 0.155672
R899 VTAIL.n66 VTAIL.n65 0.155672
R900 VTAIL.n66 VTAIL.n3 0.155672
R901 VTAIL.n73 VTAIL.n3 0.155672
R902 VTAIL.n105 VTAIL.n97 0.155672
R903 VTAIL.n106 VTAIL.n105 0.155672
R904 VTAIL.n106 VTAIL.n93 0.155672
R905 VTAIL.n113 VTAIL.n93 0.155672
R906 VTAIL.n114 VTAIL.n113 0.155672
R907 VTAIL.n114 VTAIL.n89 0.155672
R908 VTAIL.n123 VTAIL.n89 0.155672
R909 VTAIL.n124 VTAIL.n123 0.155672
R910 VTAIL.n124 VTAIL.n85 0.155672
R911 VTAIL.n131 VTAIL.n85 0.155672
R912 VTAIL.n132 VTAIL.n131 0.155672
R913 VTAIL.n132 VTAIL.n81 0.155672
R914 VTAIL.n139 VTAIL.n81 0.155672
R915 VTAIL.n140 VTAIL.n139 0.155672
R916 VTAIL.n140 VTAIL.n77 0.155672
R917 VTAIL.n147 VTAIL.n77 0.155672
R918 VTAIL.n181 VTAIL.n173 0.155672
R919 VTAIL.n182 VTAIL.n181 0.155672
R920 VTAIL.n182 VTAIL.n169 0.155672
R921 VTAIL.n189 VTAIL.n169 0.155672
R922 VTAIL.n190 VTAIL.n189 0.155672
R923 VTAIL.n190 VTAIL.n165 0.155672
R924 VTAIL.n199 VTAIL.n165 0.155672
R925 VTAIL.n200 VTAIL.n199 0.155672
R926 VTAIL.n200 VTAIL.n161 0.155672
R927 VTAIL.n207 VTAIL.n161 0.155672
R928 VTAIL.n208 VTAIL.n207 0.155672
R929 VTAIL.n208 VTAIL.n157 0.155672
R930 VTAIL.n215 VTAIL.n157 0.155672
R931 VTAIL.n216 VTAIL.n215 0.155672
R932 VTAIL.n216 VTAIL.n153 0.155672
R933 VTAIL.n223 VTAIL.n153 0.155672
R934 VTAIL.n523 VTAIL.n453 0.155672
R935 VTAIL.n516 VTAIL.n453 0.155672
R936 VTAIL.n516 VTAIL.n515 0.155672
R937 VTAIL.n515 VTAIL.n457 0.155672
R938 VTAIL.n508 VTAIL.n457 0.155672
R939 VTAIL.n508 VTAIL.n507 0.155672
R940 VTAIL.n507 VTAIL.n461 0.155672
R941 VTAIL.n500 VTAIL.n461 0.155672
R942 VTAIL.n500 VTAIL.n499 0.155672
R943 VTAIL.n499 VTAIL.n465 0.155672
R944 VTAIL.n492 VTAIL.n465 0.155672
R945 VTAIL.n492 VTAIL.n491 0.155672
R946 VTAIL.n491 VTAIL.n471 0.155672
R947 VTAIL.n484 VTAIL.n471 0.155672
R948 VTAIL.n484 VTAIL.n483 0.155672
R949 VTAIL.n483 VTAIL.n475 0.155672
R950 VTAIL.n447 VTAIL.n377 0.155672
R951 VTAIL.n440 VTAIL.n377 0.155672
R952 VTAIL.n440 VTAIL.n439 0.155672
R953 VTAIL.n439 VTAIL.n381 0.155672
R954 VTAIL.n432 VTAIL.n381 0.155672
R955 VTAIL.n432 VTAIL.n431 0.155672
R956 VTAIL.n431 VTAIL.n385 0.155672
R957 VTAIL.n424 VTAIL.n385 0.155672
R958 VTAIL.n424 VTAIL.n423 0.155672
R959 VTAIL.n423 VTAIL.n389 0.155672
R960 VTAIL.n416 VTAIL.n389 0.155672
R961 VTAIL.n416 VTAIL.n415 0.155672
R962 VTAIL.n415 VTAIL.n395 0.155672
R963 VTAIL.n408 VTAIL.n395 0.155672
R964 VTAIL.n408 VTAIL.n407 0.155672
R965 VTAIL.n407 VTAIL.n399 0.155672
R966 VTAIL.n373 VTAIL.n303 0.155672
R967 VTAIL.n366 VTAIL.n303 0.155672
R968 VTAIL.n366 VTAIL.n365 0.155672
R969 VTAIL.n365 VTAIL.n307 0.155672
R970 VTAIL.n358 VTAIL.n307 0.155672
R971 VTAIL.n358 VTAIL.n357 0.155672
R972 VTAIL.n357 VTAIL.n311 0.155672
R973 VTAIL.n350 VTAIL.n311 0.155672
R974 VTAIL.n350 VTAIL.n349 0.155672
R975 VTAIL.n349 VTAIL.n315 0.155672
R976 VTAIL.n342 VTAIL.n315 0.155672
R977 VTAIL.n342 VTAIL.n341 0.155672
R978 VTAIL.n341 VTAIL.n321 0.155672
R979 VTAIL.n334 VTAIL.n321 0.155672
R980 VTAIL.n334 VTAIL.n333 0.155672
R981 VTAIL.n333 VTAIL.n325 0.155672
R982 VTAIL.n297 VTAIL.n227 0.155672
R983 VTAIL.n290 VTAIL.n227 0.155672
R984 VTAIL.n290 VTAIL.n289 0.155672
R985 VTAIL.n289 VTAIL.n231 0.155672
R986 VTAIL.n282 VTAIL.n231 0.155672
R987 VTAIL.n282 VTAIL.n281 0.155672
R988 VTAIL.n281 VTAIL.n235 0.155672
R989 VTAIL.n274 VTAIL.n235 0.155672
R990 VTAIL.n274 VTAIL.n273 0.155672
R991 VTAIL.n273 VTAIL.n239 0.155672
R992 VTAIL.n266 VTAIL.n239 0.155672
R993 VTAIL.n266 VTAIL.n265 0.155672
R994 VTAIL.n265 VTAIL.n245 0.155672
R995 VTAIL.n258 VTAIL.n245 0.155672
R996 VTAIL.n258 VTAIL.n257 0.155672
R997 VTAIL.n257 VTAIL.n249 0.155672
R998 VTAIL VTAIL.n1 0.0586897
R999 VN.n5 VN.t6 270.158
R1000 VN.n25 VN.t4 270.158
R1001 VN.n4 VN.t0 239.938
R1002 VN.n10 VN.t5 239.938
R1003 VN.n17 VN.t3 239.938
R1004 VN.n24 VN.t1 239.938
R1005 VN.n22 VN.t2 239.938
R1006 VN.n36 VN.t7 239.938
R1007 VN.n18 VN.n17 171.875
R1008 VN.n37 VN.n36 171.875
R1009 VN.n35 VN.n19 161.3
R1010 VN.n34 VN.n33 161.3
R1011 VN.n32 VN.n20 161.3
R1012 VN.n31 VN.n30 161.3
R1013 VN.n29 VN.n21 161.3
R1014 VN.n28 VN.n27 161.3
R1015 VN.n26 VN.n23 161.3
R1016 VN.n16 VN.n0 161.3
R1017 VN.n15 VN.n14 161.3
R1018 VN.n13 VN.n1 161.3
R1019 VN.n12 VN.n11 161.3
R1020 VN.n9 VN.n2 161.3
R1021 VN.n8 VN.n7 161.3
R1022 VN.n6 VN.n3 161.3
R1023 VN.n5 VN.n4 60.629
R1024 VN.n25 VN.n24 60.629
R1025 VN.n9 VN.n8 56.5617
R1026 VN.n29 VN.n28 56.5617
R1027 VN VN.n37 46.5933
R1028 VN.n15 VN.n1 46.3896
R1029 VN.n34 VN.n20 46.3896
R1030 VN.n16 VN.n15 34.7644
R1031 VN.n35 VN.n34 34.7644
R1032 VN.n26 VN.n25 26.9001
R1033 VN.n6 VN.n5 26.9001
R1034 VN.n8 VN.n3 24.5923
R1035 VN.n11 VN.n9 24.5923
R1036 VN.n28 VN.n23 24.5923
R1037 VN.n30 VN.n29 24.5923
R1038 VN.n10 VN.n1 19.9199
R1039 VN.n22 VN.n20 19.9199
R1040 VN.n17 VN.n16 14.0178
R1041 VN.n36 VN.n35 14.0178
R1042 VN.n4 VN.n3 4.67295
R1043 VN.n11 VN.n10 4.67295
R1044 VN.n24 VN.n23 4.67295
R1045 VN.n30 VN.n22 4.67295
R1046 VN.n37 VN.n19 0.189894
R1047 VN.n33 VN.n19 0.189894
R1048 VN.n33 VN.n32 0.189894
R1049 VN.n32 VN.n31 0.189894
R1050 VN.n31 VN.n21 0.189894
R1051 VN.n27 VN.n21 0.189894
R1052 VN.n27 VN.n26 0.189894
R1053 VN.n7 VN.n6 0.189894
R1054 VN.n7 VN.n2 0.189894
R1055 VN.n12 VN.n2 0.189894
R1056 VN.n13 VN.n12 0.189894
R1057 VN.n14 VN.n13 0.189894
R1058 VN.n14 VN.n0 0.189894
R1059 VN.n18 VN.n0 0.189894
R1060 VN VN.n18 0.0516364
R1061 VDD2.n2 VDD2.n1 72.5659
R1062 VDD2.n2 VDD2.n0 72.5659
R1063 VDD2 VDD2.n5 72.5631
R1064 VDD2.n4 VDD2.n3 71.893
R1065 VDD2.n4 VDD2.n2 41.9437
R1066 VDD2.n5 VDD2.t6 2.40116
R1067 VDD2.n5 VDD2.t3 2.40116
R1068 VDD2.n3 VDD2.t0 2.40116
R1069 VDD2.n3 VDD2.t5 2.40116
R1070 VDD2.n1 VDD2.t2 2.40116
R1071 VDD2.n1 VDD2.t4 2.40116
R1072 VDD2.n0 VDD2.t1 2.40116
R1073 VDD2.n0 VDD2.t7 2.40116
R1074 VDD2 VDD2.n4 0.787138
R1075 B.n483 B.n74 585
R1076 B.n485 B.n484 585
R1077 B.n486 B.n73 585
R1078 B.n488 B.n487 585
R1079 B.n489 B.n72 585
R1080 B.n491 B.n490 585
R1081 B.n492 B.n71 585
R1082 B.n494 B.n493 585
R1083 B.n495 B.n70 585
R1084 B.n497 B.n496 585
R1085 B.n498 B.n69 585
R1086 B.n500 B.n499 585
R1087 B.n501 B.n68 585
R1088 B.n503 B.n502 585
R1089 B.n504 B.n67 585
R1090 B.n506 B.n505 585
R1091 B.n507 B.n66 585
R1092 B.n509 B.n508 585
R1093 B.n510 B.n65 585
R1094 B.n512 B.n511 585
R1095 B.n513 B.n64 585
R1096 B.n515 B.n514 585
R1097 B.n516 B.n63 585
R1098 B.n518 B.n517 585
R1099 B.n519 B.n62 585
R1100 B.n521 B.n520 585
R1101 B.n522 B.n61 585
R1102 B.n524 B.n523 585
R1103 B.n525 B.n60 585
R1104 B.n527 B.n526 585
R1105 B.n528 B.n59 585
R1106 B.n530 B.n529 585
R1107 B.n531 B.n58 585
R1108 B.n533 B.n532 585
R1109 B.n534 B.n57 585
R1110 B.n536 B.n535 585
R1111 B.n537 B.n56 585
R1112 B.n539 B.n538 585
R1113 B.n540 B.n55 585
R1114 B.n542 B.n541 585
R1115 B.n543 B.n54 585
R1116 B.n545 B.n544 585
R1117 B.n546 B.n53 585
R1118 B.n548 B.n547 585
R1119 B.n549 B.n49 585
R1120 B.n551 B.n550 585
R1121 B.n552 B.n48 585
R1122 B.n554 B.n553 585
R1123 B.n555 B.n47 585
R1124 B.n557 B.n556 585
R1125 B.n558 B.n46 585
R1126 B.n560 B.n559 585
R1127 B.n561 B.n45 585
R1128 B.n563 B.n562 585
R1129 B.n564 B.n44 585
R1130 B.n566 B.n565 585
R1131 B.n568 B.n41 585
R1132 B.n570 B.n569 585
R1133 B.n571 B.n40 585
R1134 B.n573 B.n572 585
R1135 B.n574 B.n39 585
R1136 B.n576 B.n575 585
R1137 B.n577 B.n38 585
R1138 B.n579 B.n578 585
R1139 B.n580 B.n37 585
R1140 B.n582 B.n581 585
R1141 B.n583 B.n36 585
R1142 B.n585 B.n584 585
R1143 B.n586 B.n35 585
R1144 B.n588 B.n587 585
R1145 B.n589 B.n34 585
R1146 B.n591 B.n590 585
R1147 B.n592 B.n33 585
R1148 B.n594 B.n593 585
R1149 B.n595 B.n32 585
R1150 B.n597 B.n596 585
R1151 B.n598 B.n31 585
R1152 B.n600 B.n599 585
R1153 B.n601 B.n30 585
R1154 B.n603 B.n602 585
R1155 B.n604 B.n29 585
R1156 B.n606 B.n605 585
R1157 B.n607 B.n28 585
R1158 B.n609 B.n608 585
R1159 B.n610 B.n27 585
R1160 B.n612 B.n611 585
R1161 B.n613 B.n26 585
R1162 B.n615 B.n614 585
R1163 B.n616 B.n25 585
R1164 B.n618 B.n617 585
R1165 B.n619 B.n24 585
R1166 B.n621 B.n620 585
R1167 B.n622 B.n23 585
R1168 B.n624 B.n623 585
R1169 B.n625 B.n22 585
R1170 B.n627 B.n626 585
R1171 B.n628 B.n21 585
R1172 B.n630 B.n629 585
R1173 B.n631 B.n20 585
R1174 B.n633 B.n632 585
R1175 B.n634 B.n19 585
R1176 B.n636 B.n635 585
R1177 B.n482 B.n481 585
R1178 B.n480 B.n75 585
R1179 B.n479 B.n478 585
R1180 B.n477 B.n76 585
R1181 B.n476 B.n475 585
R1182 B.n474 B.n77 585
R1183 B.n473 B.n472 585
R1184 B.n471 B.n78 585
R1185 B.n470 B.n469 585
R1186 B.n468 B.n79 585
R1187 B.n467 B.n466 585
R1188 B.n465 B.n80 585
R1189 B.n464 B.n463 585
R1190 B.n462 B.n81 585
R1191 B.n461 B.n460 585
R1192 B.n459 B.n82 585
R1193 B.n458 B.n457 585
R1194 B.n456 B.n83 585
R1195 B.n455 B.n454 585
R1196 B.n453 B.n84 585
R1197 B.n452 B.n451 585
R1198 B.n450 B.n85 585
R1199 B.n449 B.n448 585
R1200 B.n447 B.n86 585
R1201 B.n446 B.n445 585
R1202 B.n444 B.n87 585
R1203 B.n443 B.n442 585
R1204 B.n441 B.n88 585
R1205 B.n440 B.n439 585
R1206 B.n438 B.n89 585
R1207 B.n437 B.n436 585
R1208 B.n435 B.n90 585
R1209 B.n434 B.n433 585
R1210 B.n432 B.n91 585
R1211 B.n431 B.n430 585
R1212 B.n429 B.n92 585
R1213 B.n428 B.n427 585
R1214 B.n426 B.n93 585
R1215 B.n425 B.n424 585
R1216 B.n423 B.n94 585
R1217 B.n422 B.n421 585
R1218 B.n420 B.n95 585
R1219 B.n419 B.n418 585
R1220 B.n417 B.n96 585
R1221 B.n416 B.n415 585
R1222 B.n414 B.n97 585
R1223 B.n413 B.n412 585
R1224 B.n411 B.n98 585
R1225 B.n410 B.n409 585
R1226 B.n408 B.n99 585
R1227 B.n407 B.n406 585
R1228 B.n405 B.n100 585
R1229 B.n404 B.n403 585
R1230 B.n402 B.n101 585
R1231 B.n401 B.n400 585
R1232 B.n399 B.n102 585
R1233 B.n398 B.n397 585
R1234 B.n396 B.n103 585
R1235 B.n395 B.n394 585
R1236 B.n393 B.n104 585
R1237 B.n392 B.n391 585
R1238 B.n390 B.n105 585
R1239 B.n389 B.n388 585
R1240 B.n387 B.n106 585
R1241 B.n386 B.n385 585
R1242 B.n384 B.n107 585
R1243 B.n383 B.n382 585
R1244 B.n228 B.n163 585
R1245 B.n230 B.n229 585
R1246 B.n231 B.n162 585
R1247 B.n233 B.n232 585
R1248 B.n234 B.n161 585
R1249 B.n236 B.n235 585
R1250 B.n237 B.n160 585
R1251 B.n239 B.n238 585
R1252 B.n240 B.n159 585
R1253 B.n242 B.n241 585
R1254 B.n243 B.n158 585
R1255 B.n245 B.n244 585
R1256 B.n246 B.n157 585
R1257 B.n248 B.n247 585
R1258 B.n249 B.n156 585
R1259 B.n251 B.n250 585
R1260 B.n252 B.n155 585
R1261 B.n254 B.n253 585
R1262 B.n255 B.n154 585
R1263 B.n257 B.n256 585
R1264 B.n258 B.n153 585
R1265 B.n260 B.n259 585
R1266 B.n261 B.n152 585
R1267 B.n263 B.n262 585
R1268 B.n264 B.n151 585
R1269 B.n266 B.n265 585
R1270 B.n267 B.n150 585
R1271 B.n269 B.n268 585
R1272 B.n270 B.n149 585
R1273 B.n272 B.n271 585
R1274 B.n273 B.n148 585
R1275 B.n275 B.n274 585
R1276 B.n276 B.n147 585
R1277 B.n278 B.n277 585
R1278 B.n279 B.n146 585
R1279 B.n281 B.n280 585
R1280 B.n282 B.n145 585
R1281 B.n284 B.n283 585
R1282 B.n285 B.n144 585
R1283 B.n287 B.n286 585
R1284 B.n288 B.n143 585
R1285 B.n290 B.n289 585
R1286 B.n291 B.n142 585
R1287 B.n293 B.n292 585
R1288 B.n294 B.n141 585
R1289 B.n296 B.n295 585
R1290 B.n298 B.n138 585
R1291 B.n300 B.n299 585
R1292 B.n301 B.n137 585
R1293 B.n303 B.n302 585
R1294 B.n304 B.n136 585
R1295 B.n306 B.n305 585
R1296 B.n307 B.n135 585
R1297 B.n309 B.n308 585
R1298 B.n310 B.n134 585
R1299 B.n312 B.n311 585
R1300 B.n314 B.n313 585
R1301 B.n315 B.n130 585
R1302 B.n317 B.n316 585
R1303 B.n318 B.n129 585
R1304 B.n320 B.n319 585
R1305 B.n321 B.n128 585
R1306 B.n323 B.n322 585
R1307 B.n324 B.n127 585
R1308 B.n326 B.n325 585
R1309 B.n327 B.n126 585
R1310 B.n329 B.n328 585
R1311 B.n330 B.n125 585
R1312 B.n332 B.n331 585
R1313 B.n333 B.n124 585
R1314 B.n335 B.n334 585
R1315 B.n336 B.n123 585
R1316 B.n338 B.n337 585
R1317 B.n339 B.n122 585
R1318 B.n341 B.n340 585
R1319 B.n342 B.n121 585
R1320 B.n344 B.n343 585
R1321 B.n345 B.n120 585
R1322 B.n347 B.n346 585
R1323 B.n348 B.n119 585
R1324 B.n350 B.n349 585
R1325 B.n351 B.n118 585
R1326 B.n353 B.n352 585
R1327 B.n354 B.n117 585
R1328 B.n356 B.n355 585
R1329 B.n357 B.n116 585
R1330 B.n359 B.n358 585
R1331 B.n360 B.n115 585
R1332 B.n362 B.n361 585
R1333 B.n363 B.n114 585
R1334 B.n365 B.n364 585
R1335 B.n366 B.n113 585
R1336 B.n368 B.n367 585
R1337 B.n369 B.n112 585
R1338 B.n371 B.n370 585
R1339 B.n372 B.n111 585
R1340 B.n374 B.n373 585
R1341 B.n375 B.n110 585
R1342 B.n377 B.n376 585
R1343 B.n378 B.n109 585
R1344 B.n380 B.n379 585
R1345 B.n381 B.n108 585
R1346 B.n227 B.n226 585
R1347 B.n225 B.n164 585
R1348 B.n224 B.n223 585
R1349 B.n222 B.n165 585
R1350 B.n221 B.n220 585
R1351 B.n219 B.n166 585
R1352 B.n218 B.n217 585
R1353 B.n216 B.n167 585
R1354 B.n215 B.n214 585
R1355 B.n213 B.n168 585
R1356 B.n212 B.n211 585
R1357 B.n210 B.n169 585
R1358 B.n209 B.n208 585
R1359 B.n207 B.n170 585
R1360 B.n206 B.n205 585
R1361 B.n204 B.n171 585
R1362 B.n203 B.n202 585
R1363 B.n201 B.n172 585
R1364 B.n200 B.n199 585
R1365 B.n198 B.n173 585
R1366 B.n197 B.n196 585
R1367 B.n195 B.n174 585
R1368 B.n194 B.n193 585
R1369 B.n192 B.n175 585
R1370 B.n191 B.n190 585
R1371 B.n189 B.n176 585
R1372 B.n188 B.n187 585
R1373 B.n186 B.n177 585
R1374 B.n185 B.n184 585
R1375 B.n183 B.n178 585
R1376 B.n182 B.n181 585
R1377 B.n180 B.n179 585
R1378 B.n2 B.n0 585
R1379 B.n685 B.n1 585
R1380 B.n684 B.n683 585
R1381 B.n682 B.n3 585
R1382 B.n681 B.n680 585
R1383 B.n679 B.n4 585
R1384 B.n678 B.n677 585
R1385 B.n676 B.n5 585
R1386 B.n675 B.n674 585
R1387 B.n673 B.n6 585
R1388 B.n672 B.n671 585
R1389 B.n670 B.n7 585
R1390 B.n669 B.n668 585
R1391 B.n667 B.n8 585
R1392 B.n666 B.n665 585
R1393 B.n664 B.n9 585
R1394 B.n663 B.n662 585
R1395 B.n661 B.n10 585
R1396 B.n660 B.n659 585
R1397 B.n658 B.n11 585
R1398 B.n657 B.n656 585
R1399 B.n655 B.n12 585
R1400 B.n654 B.n653 585
R1401 B.n652 B.n13 585
R1402 B.n651 B.n650 585
R1403 B.n649 B.n14 585
R1404 B.n648 B.n647 585
R1405 B.n646 B.n15 585
R1406 B.n645 B.n644 585
R1407 B.n643 B.n16 585
R1408 B.n642 B.n641 585
R1409 B.n640 B.n17 585
R1410 B.n639 B.n638 585
R1411 B.n637 B.n18 585
R1412 B.n687 B.n686 585
R1413 B.n228 B.n227 482.89
R1414 B.n637 B.n636 482.89
R1415 B.n383 B.n108 482.89
R1416 B.n481 B.n74 482.89
R1417 B.n131 B.t0 444.815
R1418 B.n139 B.t6 444.815
R1419 B.n42 B.t9 444.815
R1420 B.n50 B.t3 444.815
R1421 B.n131 B.t2 436.291
R1422 B.n50 B.t4 436.291
R1423 B.n139 B.t8 436.291
R1424 B.n42 B.t10 436.291
R1425 B.n132 B.t1 403.515
R1426 B.n51 B.t5 403.515
R1427 B.n140 B.t7 403.515
R1428 B.n43 B.t11 403.515
R1429 B.n227 B.n164 163.367
R1430 B.n223 B.n164 163.367
R1431 B.n223 B.n222 163.367
R1432 B.n222 B.n221 163.367
R1433 B.n221 B.n166 163.367
R1434 B.n217 B.n166 163.367
R1435 B.n217 B.n216 163.367
R1436 B.n216 B.n215 163.367
R1437 B.n215 B.n168 163.367
R1438 B.n211 B.n168 163.367
R1439 B.n211 B.n210 163.367
R1440 B.n210 B.n209 163.367
R1441 B.n209 B.n170 163.367
R1442 B.n205 B.n170 163.367
R1443 B.n205 B.n204 163.367
R1444 B.n204 B.n203 163.367
R1445 B.n203 B.n172 163.367
R1446 B.n199 B.n172 163.367
R1447 B.n199 B.n198 163.367
R1448 B.n198 B.n197 163.367
R1449 B.n197 B.n174 163.367
R1450 B.n193 B.n174 163.367
R1451 B.n193 B.n192 163.367
R1452 B.n192 B.n191 163.367
R1453 B.n191 B.n176 163.367
R1454 B.n187 B.n176 163.367
R1455 B.n187 B.n186 163.367
R1456 B.n186 B.n185 163.367
R1457 B.n185 B.n178 163.367
R1458 B.n181 B.n178 163.367
R1459 B.n181 B.n180 163.367
R1460 B.n180 B.n2 163.367
R1461 B.n686 B.n2 163.367
R1462 B.n686 B.n685 163.367
R1463 B.n685 B.n684 163.367
R1464 B.n684 B.n3 163.367
R1465 B.n680 B.n3 163.367
R1466 B.n680 B.n679 163.367
R1467 B.n679 B.n678 163.367
R1468 B.n678 B.n5 163.367
R1469 B.n674 B.n5 163.367
R1470 B.n674 B.n673 163.367
R1471 B.n673 B.n672 163.367
R1472 B.n672 B.n7 163.367
R1473 B.n668 B.n7 163.367
R1474 B.n668 B.n667 163.367
R1475 B.n667 B.n666 163.367
R1476 B.n666 B.n9 163.367
R1477 B.n662 B.n9 163.367
R1478 B.n662 B.n661 163.367
R1479 B.n661 B.n660 163.367
R1480 B.n660 B.n11 163.367
R1481 B.n656 B.n11 163.367
R1482 B.n656 B.n655 163.367
R1483 B.n655 B.n654 163.367
R1484 B.n654 B.n13 163.367
R1485 B.n650 B.n13 163.367
R1486 B.n650 B.n649 163.367
R1487 B.n649 B.n648 163.367
R1488 B.n648 B.n15 163.367
R1489 B.n644 B.n15 163.367
R1490 B.n644 B.n643 163.367
R1491 B.n643 B.n642 163.367
R1492 B.n642 B.n17 163.367
R1493 B.n638 B.n17 163.367
R1494 B.n638 B.n637 163.367
R1495 B.n229 B.n228 163.367
R1496 B.n229 B.n162 163.367
R1497 B.n233 B.n162 163.367
R1498 B.n234 B.n233 163.367
R1499 B.n235 B.n234 163.367
R1500 B.n235 B.n160 163.367
R1501 B.n239 B.n160 163.367
R1502 B.n240 B.n239 163.367
R1503 B.n241 B.n240 163.367
R1504 B.n241 B.n158 163.367
R1505 B.n245 B.n158 163.367
R1506 B.n246 B.n245 163.367
R1507 B.n247 B.n246 163.367
R1508 B.n247 B.n156 163.367
R1509 B.n251 B.n156 163.367
R1510 B.n252 B.n251 163.367
R1511 B.n253 B.n252 163.367
R1512 B.n253 B.n154 163.367
R1513 B.n257 B.n154 163.367
R1514 B.n258 B.n257 163.367
R1515 B.n259 B.n258 163.367
R1516 B.n259 B.n152 163.367
R1517 B.n263 B.n152 163.367
R1518 B.n264 B.n263 163.367
R1519 B.n265 B.n264 163.367
R1520 B.n265 B.n150 163.367
R1521 B.n269 B.n150 163.367
R1522 B.n270 B.n269 163.367
R1523 B.n271 B.n270 163.367
R1524 B.n271 B.n148 163.367
R1525 B.n275 B.n148 163.367
R1526 B.n276 B.n275 163.367
R1527 B.n277 B.n276 163.367
R1528 B.n277 B.n146 163.367
R1529 B.n281 B.n146 163.367
R1530 B.n282 B.n281 163.367
R1531 B.n283 B.n282 163.367
R1532 B.n283 B.n144 163.367
R1533 B.n287 B.n144 163.367
R1534 B.n288 B.n287 163.367
R1535 B.n289 B.n288 163.367
R1536 B.n289 B.n142 163.367
R1537 B.n293 B.n142 163.367
R1538 B.n294 B.n293 163.367
R1539 B.n295 B.n294 163.367
R1540 B.n295 B.n138 163.367
R1541 B.n300 B.n138 163.367
R1542 B.n301 B.n300 163.367
R1543 B.n302 B.n301 163.367
R1544 B.n302 B.n136 163.367
R1545 B.n306 B.n136 163.367
R1546 B.n307 B.n306 163.367
R1547 B.n308 B.n307 163.367
R1548 B.n308 B.n134 163.367
R1549 B.n312 B.n134 163.367
R1550 B.n313 B.n312 163.367
R1551 B.n313 B.n130 163.367
R1552 B.n317 B.n130 163.367
R1553 B.n318 B.n317 163.367
R1554 B.n319 B.n318 163.367
R1555 B.n319 B.n128 163.367
R1556 B.n323 B.n128 163.367
R1557 B.n324 B.n323 163.367
R1558 B.n325 B.n324 163.367
R1559 B.n325 B.n126 163.367
R1560 B.n329 B.n126 163.367
R1561 B.n330 B.n329 163.367
R1562 B.n331 B.n330 163.367
R1563 B.n331 B.n124 163.367
R1564 B.n335 B.n124 163.367
R1565 B.n336 B.n335 163.367
R1566 B.n337 B.n336 163.367
R1567 B.n337 B.n122 163.367
R1568 B.n341 B.n122 163.367
R1569 B.n342 B.n341 163.367
R1570 B.n343 B.n342 163.367
R1571 B.n343 B.n120 163.367
R1572 B.n347 B.n120 163.367
R1573 B.n348 B.n347 163.367
R1574 B.n349 B.n348 163.367
R1575 B.n349 B.n118 163.367
R1576 B.n353 B.n118 163.367
R1577 B.n354 B.n353 163.367
R1578 B.n355 B.n354 163.367
R1579 B.n355 B.n116 163.367
R1580 B.n359 B.n116 163.367
R1581 B.n360 B.n359 163.367
R1582 B.n361 B.n360 163.367
R1583 B.n361 B.n114 163.367
R1584 B.n365 B.n114 163.367
R1585 B.n366 B.n365 163.367
R1586 B.n367 B.n366 163.367
R1587 B.n367 B.n112 163.367
R1588 B.n371 B.n112 163.367
R1589 B.n372 B.n371 163.367
R1590 B.n373 B.n372 163.367
R1591 B.n373 B.n110 163.367
R1592 B.n377 B.n110 163.367
R1593 B.n378 B.n377 163.367
R1594 B.n379 B.n378 163.367
R1595 B.n379 B.n108 163.367
R1596 B.n384 B.n383 163.367
R1597 B.n385 B.n384 163.367
R1598 B.n385 B.n106 163.367
R1599 B.n389 B.n106 163.367
R1600 B.n390 B.n389 163.367
R1601 B.n391 B.n390 163.367
R1602 B.n391 B.n104 163.367
R1603 B.n395 B.n104 163.367
R1604 B.n396 B.n395 163.367
R1605 B.n397 B.n396 163.367
R1606 B.n397 B.n102 163.367
R1607 B.n401 B.n102 163.367
R1608 B.n402 B.n401 163.367
R1609 B.n403 B.n402 163.367
R1610 B.n403 B.n100 163.367
R1611 B.n407 B.n100 163.367
R1612 B.n408 B.n407 163.367
R1613 B.n409 B.n408 163.367
R1614 B.n409 B.n98 163.367
R1615 B.n413 B.n98 163.367
R1616 B.n414 B.n413 163.367
R1617 B.n415 B.n414 163.367
R1618 B.n415 B.n96 163.367
R1619 B.n419 B.n96 163.367
R1620 B.n420 B.n419 163.367
R1621 B.n421 B.n420 163.367
R1622 B.n421 B.n94 163.367
R1623 B.n425 B.n94 163.367
R1624 B.n426 B.n425 163.367
R1625 B.n427 B.n426 163.367
R1626 B.n427 B.n92 163.367
R1627 B.n431 B.n92 163.367
R1628 B.n432 B.n431 163.367
R1629 B.n433 B.n432 163.367
R1630 B.n433 B.n90 163.367
R1631 B.n437 B.n90 163.367
R1632 B.n438 B.n437 163.367
R1633 B.n439 B.n438 163.367
R1634 B.n439 B.n88 163.367
R1635 B.n443 B.n88 163.367
R1636 B.n444 B.n443 163.367
R1637 B.n445 B.n444 163.367
R1638 B.n445 B.n86 163.367
R1639 B.n449 B.n86 163.367
R1640 B.n450 B.n449 163.367
R1641 B.n451 B.n450 163.367
R1642 B.n451 B.n84 163.367
R1643 B.n455 B.n84 163.367
R1644 B.n456 B.n455 163.367
R1645 B.n457 B.n456 163.367
R1646 B.n457 B.n82 163.367
R1647 B.n461 B.n82 163.367
R1648 B.n462 B.n461 163.367
R1649 B.n463 B.n462 163.367
R1650 B.n463 B.n80 163.367
R1651 B.n467 B.n80 163.367
R1652 B.n468 B.n467 163.367
R1653 B.n469 B.n468 163.367
R1654 B.n469 B.n78 163.367
R1655 B.n473 B.n78 163.367
R1656 B.n474 B.n473 163.367
R1657 B.n475 B.n474 163.367
R1658 B.n475 B.n76 163.367
R1659 B.n479 B.n76 163.367
R1660 B.n480 B.n479 163.367
R1661 B.n481 B.n480 163.367
R1662 B.n636 B.n19 163.367
R1663 B.n632 B.n19 163.367
R1664 B.n632 B.n631 163.367
R1665 B.n631 B.n630 163.367
R1666 B.n630 B.n21 163.367
R1667 B.n626 B.n21 163.367
R1668 B.n626 B.n625 163.367
R1669 B.n625 B.n624 163.367
R1670 B.n624 B.n23 163.367
R1671 B.n620 B.n23 163.367
R1672 B.n620 B.n619 163.367
R1673 B.n619 B.n618 163.367
R1674 B.n618 B.n25 163.367
R1675 B.n614 B.n25 163.367
R1676 B.n614 B.n613 163.367
R1677 B.n613 B.n612 163.367
R1678 B.n612 B.n27 163.367
R1679 B.n608 B.n27 163.367
R1680 B.n608 B.n607 163.367
R1681 B.n607 B.n606 163.367
R1682 B.n606 B.n29 163.367
R1683 B.n602 B.n29 163.367
R1684 B.n602 B.n601 163.367
R1685 B.n601 B.n600 163.367
R1686 B.n600 B.n31 163.367
R1687 B.n596 B.n31 163.367
R1688 B.n596 B.n595 163.367
R1689 B.n595 B.n594 163.367
R1690 B.n594 B.n33 163.367
R1691 B.n590 B.n33 163.367
R1692 B.n590 B.n589 163.367
R1693 B.n589 B.n588 163.367
R1694 B.n588 B.n35 163.367
R1695 B.n584 B.n35 163.367
R1696 B.n584 B.n583 163.367
R1697 B.n583 B.n582 163.367
R1698 B.n582 B.n37 163.367
R1699 B.n578 B.n37 163.367
R1700 B.n578 B.n577 163.367
R1701 B.n577 B.n576 163.367
R1702 B.n576 B.n39 163.367
R1703 B.n572 B.n39 163.367
R1704 B.n572 B.n571 163.367
R1705 B.n571 B.n570 163.367
R1706 B.n570 B.n41 163.367
R1707 B.n565 B.n41 163.367
R1708 B.n565 B.n564 163.367
R1709 B.n564 B.n563 163.367
R1710 B.n563 B.n45 163.367
R1711 B.n559 B.n45 163.367
R1712 B.n559 B.n558 163.367
R1713 B.n558 B.n557 163.367
R1714 B.n557 B.n47 163.367
R1715 B.n553 B.n47 163.367
R1716 B.n553 B.n552 163.367
R1717 B.n552 B.n551 163.367
R1718 B.n551 B.n49 163.367
R1719 B.n547 B.n49 163.367
R1720 B.n547 B.n546 163.367
R1721 B.n546 B.n545 163.367
R1722 B.n545 B.n54 163.367
R1723 B.n541 B.n54 163.367
R1724 B.n541 B.n540 163.367
R1725 B.n540 B.n539 163.367
R1726 B.n539 B.n56 163.367
R1727 B.n535 B.n56 163.367
R1728 B.n535 B.n534 163.367
R1729 B.n534 B.n533 163.367
R1730 B.n533 B.n58 163.367
R1731 B.n529 B.n58 163.367
R1732 B.n529 B.n528 163.367
R1733 B.n528 B.n527 163.367
R1734 B.n527 B.n60 163.367
R1735 B.n523 B.n60 163.367
R1736 B.n523 B.n522 163.367
R1737 B.n522 B.n521 163.367
R1738 B.n521 B.n62 163.367
R1739 B.n517 B.n62 163.367
R1740 B.n517 B.n516 163.367
R1741 B.n516 B.n515 163.367
R1742 B.n515 B.n64 163.367
R1743 B.n511 B.n64 163.367
R1744 B.n511 B.n510 163.367
R1745 B.n510 B.n509 163.367
R1746 B.n509 B.n66 163.367
R1747 B.n505 B.n66 163.367
R1748 B.n505 B.n504 163.367
R1749 B.n504 B.n503 163.367
R1750 B.n503 B.n68 163.367
R1751 B.n499 B.n68 163.367
R1752 B.n499 B.n498 163.367
R1753 B.n498 B.n497 163.367
R1754 B.n497 B.n70 163.367
R1755 B.n493 B.n70 163.367
R1756 B.n493 B.n492 163.367
R1757 B.n492 B.n491 163.367
R1758 B.n491 B.n72 163.367
R1759 B.n487 B.n72 163.367
R1760 B.n487 B.n486 163.367
R1761 B.n486 B.n485 163.367
R1762 B.n485 B.n74 163.367
R1763 B.n133 B.n132 59.5399
R1764 B.n297 B.n140 59.5399
R1765 B.n567 B.n43 59.5399
R1766 B.n52 B.n51 59.5399
R1767 B.n132 B.n131 32.7763
R1768 B.n140 B.n139 32.7763
R1769 B.n43 B.n42 32.7763
R1770 B.n51 B.n50 32.7763
R1771 B.n635 B.n18 31.3761
R1772 B.n483 B.n482 31.3761
R1773 B.n382 B.n381 31.3761
R1774 B.n226 B.n163 31.3761
R1775 B B.n687 18.0485
R1776 B.n635 B.n634 10.6151
R1777 B.n634 B.n633 10.6151
R1778 B.n633 B.n20 10.6151
R1779 B.n629 B.n20 10.6151
R1780 B.n629 B.n628 10.6151
R1781 B.n628 B.n627 10.6151
R1782 B.n627 B.n22 10.6151
R1783 B.n623 B.n22 10.6151
R1784 B.n623 B.n622 10.6151
R1785 B.n622 B.n621 10.6151
R1786 B.n621 B.n24 10.6151
R1787 B.n617 B.n24 10.6151
R1788 B.n617 B.n616 10.6151
R1789 B.n616 B.n615 10.6151
R1790 B.n615 B.n26 10.6151
R1791 B.n611 B.n26 10.6151
R1792 B.n611 B.n610 10.6151
R1793 B.n610 B.n609 10.6151
R1794 B.n609 B.n28 10.6151
R1795 B.n605 B.n28 10.6151
R1796 B.n605 B.n604 10.6151
R1797 B.n604 B.n603 10.6151
R1798 B.n603 B.n30 10.6151
R1799 B.n599 B.n30 10.6151
R1800 B.n599 B.n598 10.6151
R1801 B.n598 B.n597 10.6151
R1802 B.n597 B.n32 10.6151
R1803 B.n593 B.n32 10.6151
R1804 B.n593 B.n592 10.6151
R1805 B.n592 B.n591 10.6151
R1806 B.n591 B.n34 10.6151
R1807 B.n587 B.n34 10.6151
R1808 B.n587 B.n586 10.6151
R1809 B.n586 B.n585 10.6151
R1810 B.n585 B.n36 10.6151
R1811 B.n581 B.n36 10.6151
R1812 B.n581 B.n580 10.6151
R1813 B.n580 B.n579 10.6151
R1814 B.n579 B.n38 10.6151
R1815 B.n575 B.n38 10.6151
R1816 B.n575 B.n574 10.6151
R1817 B.n574 B.n573 10.6151
R1818 B.n573 B.n40 10.6151
R1819 B.n569 B.n40 10.6151
R1820 B.n569 B.n568 10.6151
R1821 B.n566 B.n44 10.6151
R1822 B.n562 B.n44 10.6151
R1823 B.n562 B.n561 10.6151
R1824 B.n561 B.n560 10.6151
R1825 B.n560 B.n46 10.6151
R1826 B.n556 B.n46 10.6151
R1827 B.n556 B.n555 10.6151
R1828 B.n555 B.n554 10.6151
R1829 B.n554 B.n48 10.6151
R1830 B.n550 B.n549 10.6151
R1831 B.n549 B.n548 10.6151
R1832 B.n548 B.n53 10.6151
R1833 B.n544 B.n53 10.6151
R1834 B.n544 B.n543 10.6151
R1835 B.n543 B.n542 10.6151
R1836 B.n542 B.n55 10.6151
R1837 B.n538 B.n55 10.6151
R1838 B.n538 B.n537 10.6151
R1839 B.n537 B.n536 10.6151
R1840 B.n536 B.n57 10.6151
R1841 B.n532 B.n57 10.6151
R1842 B.n532 B.n531 10.6151
R1843 B.n531 B.n530 10.6151
R1844 B.n530 B.n59 10.6151
R1845 B.n526 B.n59 10.6151
R1846 B.n526 B.n525 10.6151
R1847 B.n525 B.n524 10.6151
R1848 B.n524 B.n61 10.6151
R1849 B.n520 B.n61 10.6151
R1850 B.n520 B.n519 10.6151
R1851 B.n519 B.n518 10.6151
R1852 B.n518 B.n63 10.6151
R1853 B.n514 B.n63 10.6151
R1854 B.n514 B.n513 10.6151
R1855 B.n513 B.n512 10.6151
R1856 B.n512 B.n65 10.6151
R1857 B.n508 B.n65 10.6151
R1858 B.n508 B.n507 10.6151
R1859 B.n507 B.n506 10.6151
R1860 B.n506 B.n67 10.6151
R1861 B.n502 B.n67 10.6151
R1862 B.n502 B.n501 10.6151
R1863 B.n501 B.n500 10.6151
R1864 B.n500 B.n69 10.6151
R1865 B.n496 B.n69 10.6151
R1866 B.n496 B.n495 10.6151
R1867 B.n495 B.n494 10.6151
R1868 B.n494 B.n71 10.6151
R1869 B.n490 B.n71 10.6151
R1870 B.n490 B.n489 10.6151
R1871 B.n489 B.n488 10.6151
R1872 B.n488 B.n73 10.6151
R1873 B.n484 B.n73 10.6151
R1874 B.n484 B.n483 10.6151
R1875 B.n382 B.n107 10.6151
R1876 B.n386 B.n107 10.6151
R1877 B.n387 B.n386 10.6151
R1878 B.n388 B.n387 10.6151
R1879 B.n388 B.n105 10.6151
R1880 B.n392 B.n105 10.6151
R1881 B.n393 B.n392 10.6151
R1882 B.n394 B.n393 10.6151
R1883 B.n394 B.n103 10.6151
R1884 B.n398 B.n103 10.6151
R1885 B.n399 B.n398 10.6151
R1886 B.n400 B.n399 10.6151
R1887 B.n400 B.n101 10.6151
R1888 B.n404 B.n101 10.6151
R1889 B.n405 B.n404 10.6151
R1890 B.n406 B.n405 10.6151
R1891 B.n406 B.n99 10.6151
R1892 B.n410 B.n99 10.6151
R1893 B.n411 B.n410 10.6151
R1894 B.n412 B.n411 10.6151
R1895 B.n412 B.n97 10.6151
R1896 B.n416 B.n97 10.6151
R1897 B.n417 B.n416 10.6151
R1898 B.n418 B.n417 10.6151
R1899 B.n418 B.n95 10.6151
R1900 B.n422 B.n95 10.6151
R1901 B.n423 B.n422 10.6151
R1902 B.n424 B.n423 10.6151
R1903 B.n424 B.n93 10.6151
R1904 B.n428 B.n93 10.6151
R1905 B.n429 B.n428 10.6151
R1906 B.n430 B.n429 10.6151
R1907 B.n430 B.n91 10.6151
R1908 B.n434 B.n91 10.6151
R1909 B.n435 B.n434 10.6151
R1910 B.n436 B.n435 10.6151
R1911 B.n436 B.n89 10.6151
R1912 B.n440 B.n89 10.6151
R1913 B.n441 B.n440 10.6151
R1914 B.n442 B.n441 10.6151
R1915 B.n442 B.n87 10.6151
R1916 B.n446 B.n87 10.6151
R1917 B.n447 B.n446 10.6151
R1918 B.n448 B.n447 10.6151
R1919 B.n448 B.n85 10.6151
R1920 B.n452 B.n85 10.6151
R1921 B.n453 B.n452 10.6151
R1922 B.n454 B.n453 10.6151
R1923 B.n454 B.n83 10.6151
R1924 B.n458 B.n83 10.6151
R1925 B.n459 B.n458 10.6151
R1926 B.n460 B.n459 10.6151
R1927 B.n460 B.n81 10.6151
R1928 B.n464 B.n81 10.6151
R1929 B.n465 B.n464 10.6151
R1930 B.n466 B.n465 10.6151
R1931 B.n466 B.n79 10.6151
R1932 B.n470 B.n79 10.6151
R1933 B.n471 B.n470 10.6151
R1934 B.n472 B.n471 10.6151
R1935 B.n472 B.n77 10.6151
R1936 B.n476 B.n77 10.6151
R1937 B.n477 B.n476 10.6151
R1938 B.n478 B.n477 10.6151
R1939 B.n478 B.n75 10.6151
R1940 B.n482 B.n75 10.6151
R1941 B.n230 B.n163 10.6151
R1942 B.n231 B.n230 10.6151
R1943 B.n232 B.n231 10.6151
R1944 B.n232 B.n161 10.6151
R1945 B.n236 B.n161 10.6151
R1946 B.n237 B.n236 10.6151
R1947 B.n238 B.n237 10.6151
R1948 B.n238 B.n159 10.6151
R1949 B.n242 B.n159 10.6151
R1950 B.n243 B.n242 10.6151
R1951 B.n244 B.n243 10.6151
R1952 B.n244 B.n157 10.6151
R1953 B.n248 B.n157 10.6151
R1954 B.n249 B.n248 10.6151
R1955 B.n250 B.n249 10.6151
R1956 B.n250 B.n155 10.6151
R1957 B.n254 B.n155 10.6151
R1958 B.n255 B.n254 10.6151
R1959 B.n256 B.n255 10.6151
R1960 B.n256 B.n153 10.6151
R1961 B.n260 B.n153 10.6151
R1962 B.n261 B.n260 10.6151
R1963 B.n262 B.n261 10.6151
R1964 B.n262 B.n151 10.6151
R1965 B.n266 B.n151 10.6151
R1966 B.n267 B.n266 10.6151
R1967 B.n268 B.n267 10.6151
R1968 B.n268 B.n149 10.6151
R1969 B.n272 B.n149 10.6151
R1970 B.n273 B.n272 10.6151
R1971 B.n274 B.n273 10.6151
R1972 B.n274 B.n147 10.6151
R1973 B.n278 B.n147 10.6151
R1974 B.n279 B.n278 10.6151
R1975 B.n280 B.n279 10.6151
R1976 B.n280 B.n145 10.6151
R1977 B.n284 B.n145 10.6151
R1978 B.n285 B.n284 10.6151
R1979 B.n286 B.n285 10.6151
R1980 B.n286 B.n143 10.6151
R1981 B.n290 B.n143 10.6151
R1982 B.n291 B.n290 10.6151
R1983 B.n292 B.n291 10.6151
R1984 B.n292 B.n141 10.6151
R1985 B.n296 B.n141 10.6151
R1986 B.n299 B.n298 10.6151
R1987 B.n299 B.n137 10.6151
R1988 B.n303 B.n137 10.6151
R1989 B.n304 B.n303 10.6151
R1990 B.n305 B.n304 10.6151
R1991 B.n305 B.n135 10.6151
R1992 B.n309 B.n135 10.6151
R1993 B.n310 B.n309 10.6151
R1994 B.n311 B.n310 10.6151
R1995 B.n315 B.n314 10.6151
R1996 B.n316 B.n315 10.6151
R1997 B.n316 B.n129 10.6151
R1998 B.n320 B.n129 10.6151
R1999 B.n321 B.n320 10.6151
R2000 B.n322 B.n321 10.6151
R2001 B.n322 B.n127 10.6151
R2002 B.n326 B.n127 10.6151
R2003 B.n327 B.n326 10.6151
R2004 B.n328 B.n327 10.6151
R2005 B.n328 B.n125 10.6151
R2006 B.n332 B.n125 10.6151
R2007 B.n333 B.n332 10.6151
R2008 B.n334 B.n333 10.6151
R2009 B.n334 B.n123 10.6151
R2010 B.n338 B.n123 10.6151
R2011 B.n339 B.n338 10.6151
R2012 B.n340 B.n339 10.6151
R2013 B.n340 B.n121 10.6151
R2014 B.n344 B.n121 10.6151
R2015 B.n345 B.n344 10.6151
R2016 B.n346 B.n345 10.6151
R2017 B.n346 B.n119 10.6151
R2018 B.n350 B.n119 10.6151
R2019 B.n351 B.n350 10.6151
R2020 B.n352 B.n351 10.6151
R2021 B.n352 B.n117 10.6151
R2022 B.n356 B.n117 10.6151
R2023 B.n357 B.n356 10.6151
R2024 B.n358 B.n357 10.6151
R2025 B.n358 B.n115 10.6151
R2026 B.n362 B.n115 10.6151
R2027 B.n363 B.n362 10.6151
R2028 B.n364 B.n363 10.6151
R2029 B.n364 B.n113 10.6151
R2030 B.n368 B.n113 10.6151
R2031 B.n369 B.n368 10.6151
R2032 B.n370 B.n369 10.6151
R2033 B.n370 B.n111 10.6151
R2034 B.n374 B.n111 10.6151
R2035 B.n375 B.n374 10.6151
R2036 B.n376 B.n375 10.6151
R2037 B.n376 B.n109 10.6151
R2038 B.n380 B.n109 10.6151
R2039 B.n381 B.n380 10.6151
R2040 B.n226 B.n225 10.6151
R2041 B.n225 B.n224 10.6151
R2042 B.n224 B.n165 10.6151
R2043 B.n220 B.n165 10.6151
R2044 B.n220 B.n219 10.6151
R2045 B.n219 B.n218 10.6151
R2046 B.n218 B.n167 10.6151
R2047 B.n214 B.n167 10.6151
R2048 B.n214 B.n213 10.6151
R2049 B.n213 B.n212 10.6151
R2050 B.n212 B.n169 10.6151
R2051 B.n208 B.n169 10.6151
R2052 B.n208 B.n207 10.6151
R2053 B.n207 B.n206 10.6151
R2054 B.n206 B.n171 10.6151
R2055 B.n202 B.n171 10.6151
R2056 B.n202 B.n201 10.6151
R2057 B.n201 B.n200 10.6151
R2058 B.n200 B.n173 10.6151
R2059 B.n196 B.n173 10.6151
R2060 B.n196 B.n195 10.6151
R2061 B.n195 B.n194 10.6151
R2062 B.n194 B.n175 10.6151
R2063 B.n190 B.n175 10.6151
R2064 B.n190 B.n189 10.6151
R2065 B.n189 B.n188 10.6151
R2066 B.n188 B.n177 10.6151
R2067 B.n184 B.n177 10.6151
R2068 B.n184 B.n183 10.6151
R2069 B.n183 B.n182 10.6151
R2070 B.n182 B.n179 10.6151
R2071 B.n179 B.n0 10.6151
R2072 B.n683 B.n1 10.6151
R2073 B.n683 B.n682 10.6151
R2074 B.n682 B.n681 10.6151
R2075 B.n681 B.n4 10.6151
R2076 B.n677 B.n4 10.6151
R2077 B.n677 B.n676 10.6151
R2078 B.n676 B.n675 10.6151
R2079 B.n675 B.n6 10.6151
R2080 B.n671 B.n6 10.6151
R2081 B.n671 B.n670 10.6151
R2082 B.n670 B.n669 10.6151
R2083 B.n669 B.n8 10.6151
R2084 B.n665 B.n8 10.6151
R2085 B.n665 B.n664 10.6151
R2086 B.n664 B.n663 10.6151
R2087 B.n663 B.n10 10.6151
R2088 B.n659 B.n10 10.6151
R2089 B.n659 B.n658 10.6151
R2090 B.n658 B.n657 10.6151
R2091 B.n657 B.n12 10.6151
R2092 B.n653 B.n12 10.6151
R2093 B.n653 B.n652 10.6151
R2094 B.n652 B.n651 10.6151
R2095 B.n651 B.n14 10.6151
R2096 B.n647 B.n14 10.6151
R2097 B.n647 B.n646 10.6151
R2098 B.n646 B.n645 10.6151
R2099 B.n645 B.n16 10.6151
R2100 B.n641 B.n16 10.6151
R2101 B.n641 B.n640 10.6151
R2102 B.n640 B.n639 10.6151
R2103 B.n639 B.n18 10.6151
R2104 B.n568 B.n567 9.36635
R2105 B.n550 B.n52 9.36635
R2106 B.n297 B.n296 9.36635
R2107 B.n314 B.n133 9.36635
R2108 B.n687 B.n0 2.81026
R2109 B.n687 B.n1 2.81026
R2110 B.n567 B.n566 1.24928
R2111 B.n52 B.n48 1.24928
R2112 B.n298 B.n297 1.24928
R2113 B.n311 B.n133 1.24928
C0 VDD2 VTAIL 9.47776f
C1 VDD2 VDD1 1.15548f
C2 VN B 0.957206f
C3 w_n2660_n3676# B 8.64834f
C4 B VP 1.52335f
C5 VN w_n2660_n3676# 5.08905f
C6 VN VP 6.42645f
C7 VTAIL B 4.7718f
C8 VTAIL VN 8.14622f
C9 B VDD1 1.31326f
C10 VN VDD1 0.149494f
C11 VDD2 B 1.37039f
C12 VDD2 VN 8.21713f
C13 w_n2660_n3676# VP 5.43072f
C14 VTAIL w_n2660_n3676# 4.52542f
C15 VTAIL VP 8.16033f
C16 w_n2660_n3676# VDD1 1.5792f
C17 VDD1 VP 8.454599f
C18 VTAIL VDD1 9.431661f
C19 VDD2 w_n2660_n3676# 1.64183f
C20 VDD2 VP 0.38773f
C21 VDD2 VSUBS 1.506725f
C22 VDD1 VSUBS 1.931826f
C23 VTAIL VSUBS 1.156341f
C24 VN VSUBS 5.32276f
C25 VP VSUBS 2.365627f
C26 B VSUBS 3.750108f
C27 w_n2660_n3676# VSUBS 0.120115p
C28 B.n0 VSUBS 0.00464f
C29 B.n1 VSUBS 0.00464f
C30 B.n2 VSUBS 0.007338f
C31 B.n3 VSUBS 0.007338f
C32 B.n4 VSUBS 0.007338f
C33 B.n5 VSUBS 0.007338f
C34 B.n6 VSUBS 0.007338f
C35 B.n7 VSUBS 0.007338f
C36 B.n8 VSUBS 0.007338f
C37 B.n9 VSUBS 0.007338f
C38 B.n10 VSUBS 0.007338f
C39 B.n11 VSUBS 0.007338f
C40 B.n12 VSUBS 0.007338f
C41 B.n13 VSUBS 0.007338f
C42 B.n14 VSUBS 0.007338f
C43 B.n15 VSUBS 0.007338f
C44 B.n16 VSUBS 0.007338f
C45 B.n17 VSUBS 0.007338f
C46 B.n18 VSUBS 0.016275f
C47 B.n19 VSUBS 0.007338f
C48 B.n20 VSUBS 0.007338f
C49 B.n21 VSUBS 0.007338f
C50 B.n22 VSUBS 0.007338f
C51 B.n23 VSUBS 0.007338f
C52 B.n24 VSUBS 0.007338f
C53 B.n25 VSUBS 0.007338f
C54 B.n26 VSUBS 0.007338f
C55 B.n27 VSUBS 0.007338f
C56 B.n28 VSUBS 0.007338f
C57 B.n29 VSUBS 0.007338f
C58 B.n30 VSUBS 0.007338f
C59 B.n31 VSUBS 0.007338f
C60 B.n32 VSUBS 0.007338f
C61 B.n33 VSUBS 0.007338f
C62 B.n34 VSUBS 0.007338f
C63 B.n35 VSUBS 0.007338f
C64 B.n36 VSUBS 0.007338f
C65 B.n37 VSUBS 0.007338f
C66 B.n38 VSUBS 0.007338f
C67 B.n39 VSUBS 0.007338f
C68 B.n40 VSUBS 0.007338f
C69 B.n41 VSUBS 0.007338f
C70 B.t11 VSUBS 0.25786f
C71 B.t10 VSUBS 0.278133f
C72 B.t9 VSUBS 0.830807f
C73 B.n42 VSUBS 0.408547f
C74 B.n43 VSUBS 0.280338f
C75 B.n44 VSUBS 0.007338f
C76 B.n45 VSUBS 0.007338f
C77 B.n46 VSUBS 0.007338f
C78 B.n47 VSUBS 0.007338f
C79 B.n48 VSUBS 0.004101f
C80 B.n49 VSUBS 0.007338f
C81 B.t5 VSUBS 0.257863f
C82 B.t4 VSUBS 0.278136f
C83 B.t3 VSUBS 0.830807f
C84 B.n50 VSUBS 0.408544f
C85 B.n51 VSUBS 0.280335f
C86 B.n52 VSUBS 0.017002f
C87 B.n53 VSUBS 0.007338f
C88 B.n54 VSUBS 0.007338f
C89 B.n55 VSUBS 0.007338f
C90 B.n56 VSUBS 0.007338f
C91 B.n57 VSUBS 0.007338f
C92 B.n58 VSUBS 0.007338f
C93 B.n59 VSUBS 0.007338f
C94 B.n60 VSUBS 0.007338f
C95 B.n61 VSUBS 0.007338f
C96 B.n62 VSUBS 0.007338f
C97 B.n63 VSUBS 0.007338f
C98 B.n64 VSUBS 0.007338f
C99 B.n65 VSUBS 0.007338f
C100 B.n66 VSUBS 0.007338f
C101 B.n67 VSUBS 0.007338f
C102 B.n68 VSUBS 0.007338f
C103 B.n69 VSUBS 0.007338f
C104 B.n70 VSUBS 0.007338f
C105 B.n71 VSUBS 0.007338f
C106 B.n72 VSUBS 0.007338f
C107 B.n73 VSUBS 0.007338f
C108 B.n74 VSUBS 0.017178f
C109 B.n75 VSUBS 0.007338f
C110 B.n76 VSUBS 0.007338f
C111 B.n77 VSUBS 0.007338f
C112 B.n78 VSUBS 0.007338f
C113 B.n79 VSUBS 0.007338f
C114 B.n80 VSUBS 0.007338f
C115 B.n81 VSUBS 0.007338f
C116 B.n82 VSUBS 0.007338f
C117 B.n83 VSUBS 0.007338f
C118 B.n84 VSUBS 0.007338f
C119 B.n85 VSUBS 0.007338f
C120 B.n86 VSUBS 0.007338f
C121 B.n87 VSUBS 0.007338f
C122 B.n88 VSUBS 0.007338f
C123 B.n89 VSUBS 0.007338f
C124 B.n90 VSUBS 0.007338f
C125 B.n91 VSUBS 0.007338f
C126 B.n92 VSUBS 0.007338f
C127 B.n93 VSUBS 0.007338f
C128 B.n94 VSUBS 0.007338f
C129 B.n95 VSUBS 0.007338f
C130 B.n96 VSUBS 0.007338f
C131 B.n97 VSUBS 0.007338f
C132 B.n98 VSUBS 0.007338f
C133 B.n99 VSUBS 0.007338f
C134 B.n100 VSUBS 0.007338f
C135 B.n101 VSUBS 0.007338f
C136 B.n102 VSUBS 0.007338f
C137 B.n103 VSUBS 0.007338f
C138 B.n104 VSUBS 0.007338f
C139 B.n105 VSUBS 0.007338f
C140 B.n106 VSUBS 0.007338f
C141 B.n107 VSUBS 0.007338f
C142 B.n108 VSUBS 0.017178f
C143 B.n109 VSUBS 0.007338f
C144 B.n110 VSUBS 0.007338f
C145 B.n111 VSUBS 0.007338f
C146 B.n112 VSUBS 0.007338f
C147 B.n113 VSUBS 0.007338f
C148 B.n114 VSUBS 0.007338f
C149 B.n115 VSUBS 0.007338f
C150 B.n116 VSUBS 0.007338f
C151 B.n117 VSUBS 0.007338f
C152 B.n118 VSUBS 0.007338f
C153 B.n119 VSUBS 0.007338f
C154 B.n120 VSUBS 0.007338f
C155 B.n121 VSUBS 0.007338f
C156 B.n122 VSUBS 0.007338f
C157 B.n123 VSUBS 0.007338f
C158 B.n124 VSUBS 0.007338f
C159 B.n125 VSUBS 0.007338f
C160 B.n126 VSUBS 0.007338f
C161 B.n127 VSUBS 0.007338f
C162 B.n128 VSUBS 0.007338f
C163 B.n129 VSUBS 0.007338f
C164 B.n130 VSUBS 0.007338f
C165 B.t1 VSUBS 0.257863f
C166 B.t2 VSUBS 0.278136f
C167 B.t0 VSUBS 0.830807f
C168 B.n131 VSUBS 0.408544f
C169 B.n132 VSUBS 0.280335f
C170 B.n133 VSUBS 0.017002f
C171 B.n134 VSUBS 0.007338f
C172 B.n135 VSUBS 0.007338f
C173 B.n136 VSUBS 0.007338f
C174 B.n137 VSUBS 0.007338f
C175 B.n138 VSUBS 0.007338f
C176 B.t7 VSUBS 0.25786f
C177 B.t8 VSUBS 0.278133f
C178 B.t6 VSUBS 0.830807f
C179 B.n139 VSUBS 0.408547f
C180 B.n140 VSUBS 0.280338f
C181 B.n141 VSUBS 0.007338f
C182 B.n142 VSUBS 0.007338f
C183 B.n143 VSUBS 0.007338f
C184 B.n144 VSUBS 0.007338f
C185 B.n145 VSUBS 0.007338f
C186 B.n146 VSUBS 0.007338f
C187 B.n147 VSUBS 0.007338f
C188 B.n148 VSUBS 0.007338f
C189 B.n149 VSUBS 0.007338f
C190 B.n150 VSUBS 0.007338f
C191 B.n151 VSUBS 0.007338f
C192 B.n152 VSUBS 0.007338f
C193 B.n153 VSUBS 0.007338f
C194 B.n154 VSUBS 0.007338f
C195 B.n155 VSUBS 0.007338f
C196 B.n156 VSUBS 0.007338f
C197 B.n157 VSUBS 0.007338f
C198 B.n158 VSUBS 0.007338f
C199 B.n159 VSUBS 0.007338f
C200 B.n160 VSUBS 0.007338f
C201 B.n161 VSUBS 0.007338f
C202 B.n162 VSUBS 0.007338f
C203 B.n163 VSUBS 0.017178f
C204 B.n164 VSUBS 0.007338f
C205 B.n165 VSUBS 0.007338f
C206 B.n166 VSUBS 0.007338f
C207 B.n167 VSUBS 0.007338f
C208 B.n168 VSUBS 0.007338f
C209 B.n169 VSUBS 0.007338f
C210 B.n170 VSUBS 0.007338f
C211 B.n171 VSUBS 0.007338f
C212 B.n172 VSUBS 0.007338f
C213 B.n173 VSUBS 0.007338f
C214 B.n174 VSUBS 0.007338f
C215 B.n175 VSUBS 0.007338f
C216 B.n176 VSUBS 0.007338f
C217 B.n177 VSUBS 0.007338f
C218 B.n178 VSUBS 0.007338f
C219 B.n179 VSUBS 0.007338f
C220 B.n180 VSUBS 0.007338f
C221 B.n181 VSUBS 0.007338f
C222 B.n182 VSUBS 0.007338f
C223 B.n183 VSUBS 0.007338f
C224 B.n184 VSUBS 0.007338f
C225 B.n185 VSUBS 0.007338f
C226 B.n186 VSUBS 0.007338f
C227 B.n187 VSUBS 0.007338f
C228 B.n188 VSUBS 0.007338f
C229 B.n189 VSUBS 0.007338f
C230 B.n190 VSUBS 0.007338f
C231 B.n191 VSUBS 0.007338f
C232 B.n192 VSUBS 0.007338f
C233 B.n193 VSUBS 0.007338f
C234 B.n194 VSUBS 0.007338f
C235 B.n195 VSUBS 0.007338f
C236 B.n196 VSUBS 0.007338f
C237 B.n197 VSUBS 0.007338f
C238 B.n198 VSUBS 0.007338f
C239 B.n199 VSUBS 0.007338f
C240 B.n200 VSUBS 0.007338f
C241 B.n201 VSUBS 0.007338f
C242 B.n202 VSUBS 0.007338f
C243 B.n203 VSUBS 0.007338f
C244 B.n204 VSUBS 0.007338f
C245 B.n205 VSUBS 0.007338f
C246 B.n206 VSUBS 0.007338f
C247 B.n207 VSUBS 0.007338f
C248 B.n208 VSUBS 0.007338f
C249 B.n209 VSUBS 0.007338f
C250 B.n210 VSUBS 0.007338f
C251 B.n211 VSUBS 0.007338f
C252 B.n212 VSUBS 0.007338f
C253 B.n213 VSUBS 0.007338f
C254 B.n214 VSUBS 0.007338f
C255 B.n215 VSUBS 0.007338f
C256 B.n216 VSUBS 0.007338f
C257 B.n217 VSUBS 0.007338f
C258 B.n218 VSUBS 0.007338f
C259 B.n219 VSUBS 0.007338f
C260 B.n220 VSUBS 0.007338f
C261 B.n221 VSUBS 0.007338f
C262 B.n222 VSUBS 0.007338f
C263 B.n223 VSUBS 0.007338f
C264 B.n224 VSUBS 0.007338f
C265 B.n225 VSUBS 0.007338f
C266 B.n226 VSUBS 0.016275f
C267 B.n227 VSUBS 0.016275f
C268 B.n228 VSUBS 0.017178f
C269 B.n229 VSUBS 0.007338f
C270 B.n230 VSUBS 0.007338f
C271 B.n231 VSUBS 0.007338f
C272 B.n232 VSUBS 0.007338f
C273 B.n233 VSUBS 0.007338f
C274 B.n234 VSUBS 0.007338f
C275 B.n235 VSUBS 0.007338f
C276 B.n236 VSUBS 0.007338f
C277 B.n237 VSUBS 0.007338f
C278 B.n238 VSUBS 0.007338f
C279 B.n239 VSUBS 0.007338f
C280 B.n240 VSUBS 0.007338f
C281 B.n241 VSUBS 0.007338f
C282 B.n242 VSUBS 0.007338f
C283 B.n243 VSUBS 0.007338f
C284 B.n244 VSUBS 0.007338f
C285 B.n245 VSUBS 0.007338f
C286 B.n246 VSUBS 0.007338f
C287 B.n247 VSUBS 0.007338f
C288 B.n248 VSUBS 0.007338f
C289 B.n249 VSUBS 0.007338f
C290 B.n250 VSUBS 0.007338f
C291 B.n251 VSUBS 0.007338f
C292 B.n252 VSUBS 0.007338f
C293 B.n253 VSUBS 0.007338f
C294 B.n254 VSUBS 0.007338f
C295 B.n255 VSUBS 0.007338f
C296 B.n256 VSUBS 0.007338f
C297 B.n257 VSUBS 0.007338f
C298 B.n258 VSUBS 0.007338f
C299 B.n259 VSUBS 0.007338f
C300 B.n260 VSUBS 0.007338f
C301 B.n261 VSUBS 0.007338f
C302 B.n262 VSUBS 0.007338f
C303 B.n263 VSUBS 0.007338f
C304 B.n264 VSUBS 0.007338f
C305 B.n265 VSUBS 0.007338f
C306 B.n266 VSUBS 0.007338f
C307 B.n267 VSUBS 0.007338f
C308 B.n268 VSUBS 0.007338f
C309 B.n269 VSUBS 0.007338f
C310 B.n270 VSUBS 0.007338f
C311 B.n271 VSUBS 0.007338f
C312 B.n272 VSUBS 0.007338f
C313 B.n273 VSUBS 0.007338f
C314 B.n274 VSUBS 0.007338f
C315 B.n275 VSUBS 0.007338f
C316 B.n276 VSUBS 0.007338f
C317 B.n277 VSUBS 0.007338f
C318 B.n278 VSUBS 0.007338f
C319 B.n279 VSUBS 0.007338f
C320 B.n280 VSUBS 0.007338f
C321 B.n281 VSUBS 0.007338f
C322 B.n282 VSUBS 0.007338f
C323 B.n283 VSUBS 0.007338f
C324 B.n284 VSUBS 0.007338f
C325 B.n285 VSUBS 0.007338f
C326 B.n286 VSUBS 0.007338f
C327 B.n287 VSUBS 0.007338f
C328 B.n288 VSUBS 0.007338f
C329 B.n289 VSUBS 0.007338f
C330 B.n290 VSUBS 0.007338f
C331 B.n291 VSUBS 0.007338f
C332 B.n292 VSUBS 0.007338f
C333 B.n293 VSUBS 0.007338f
C334 B.n294 VSUBS 0.007338f
C335 B.n295 VSUBS 0.007338f
C336 B.n296 VSUBS 0.006906f
C337 B.n297 VSUBS 0.017002f
C338 B.n298 VSUBS 0.004101f
C339 B.n299 VSUBS 0.007338f
C340 B.n300 VSUBS 0.007338f
C341 B.n301 VSUBS 0.007338f
C342 B.n302 VSUBS 0.007338f
C343 B.n303 VSUBS 0.007338f
C344 B.n304 VSUBS 0.007338f
C345 B.n305 VSUBS 0.007338f
C346 B.n306 VSUBS 0.007338f
C347 B.n307 VSUBS 0.007338f
C348 B.n308 VSUBS 0.007338f
C349 B.n309 VSUBS 0.007338f
C350 B.n310 VSUBS 0.007338f
C351 B.n311 VSUBS 0.004101f
C352 B.n312 VSUBS 0.007338f
C353 B.n313 VSUBS 0.007338f
C354 B.n314 VSUBS 0.006906f
C355 B.n315 VSUBS 0.007338f
C356 B.n316 VSUBS 0.007338f
C357 B.n317 VSUBS 0.007338f
C358 B.n318 VSUBS 0.007338f
C359 B.n319 VSUBS 0.007338f
C360 B.n320 VSUBS 0.007338f
C361 B.n321 VSUBS 0.007338f
C362 B.n322 VSUBS 0.007338f
C363 B.n323 VSUBS 0.007338f
C364 B.n324 VSUBS 0.007338f
C365 B.n325 VSUBS 0.007338f
C366 B.n326 VSUBS 0.007338f
C367 B.n327 VSUBS 0.007338f
C368 B.n328 VSUBS 0.007338f
C369 B.n329 VSUBS 0.007338f
C370 B.n330 VSUBS 0.007338f
C371 B.n331 VSUBS 0.007338f
C372 B.n332 VSUBS 0.007338f
C373 B.n333 VSUBS 0.007338f
C374 B.n334 VSUBS 0.007338f
C375 B.n335 VSUBS 0.007338f
C376 B.n336 VSUBS 0.007338f
C377 B.n337 VSUBS 0.007338f
C378 B.n338 VSUBS 0.007338f
C379 B.n339 VSUBS 0.007338f
C380 B.n340 VSUBS 0.007338f
C381 B.n341 VSUBS 0.007338f
C382 B.n342 VSUBS 0.007338f
C383 B.n343 VSUBS 0.007338f
C384 B.n344 VSUBS 0.007338f
C385 B.n345 VSUBS 0.007338f
C386 B.n346 VSUBS 0.007338f
C387 B.n347 VSUBS 0.007338f
C388 B.n348 VSUBS 0.007338f
C389 B.n349 VSUBS 0.007338f
C390 B.n350 VSUBS 0.007338f
C391 B.n351 VSUBS 0.007338f
C392 B.n352 VSUBS 0.007338f
C393 B.n353 VSUBS 0.007338f
C394 B.n354 VSUBS 0.007338f
C395 B.n355 VSUBS 0.007338f
C396 B.n356 VSUBS 0.007338f
C397 B.n357 VSUBS 0.007338f
C398 B.n358 VSUBS 0.007338f
C399 B.n359 VSUBS 0.007338f
C400 B.n360 VSUBS 0.007338f
C401 B.n361 VSUBS 0.007338f
C402 B.n362 VSUBS 0.007338f
C403 B.n363 VSUBS 0.007338f
C404 B.n364 VSUBS 0.007338f
C405 B.n365 VSUBS 0.007338f
C406 B.n366 VSUBS 0.007338f
C407 B.n367 VSUBS 0.007338f
C408 B.n368 VSUBS 0.007338f
C409 B.n369 VSUBS 0.007338f
C410 B.n370 VSUBS 0.007338f
C411 B.n371 VSUBS 0.007338f
C412 B.n372 VSUBS 0.007338f
C413 B.n373 VSUBS 0.007338f
C414 B.n374 VSUBS 0.007338f
C415 B.n375 VSUBS 0.007338f
C416 B.n376 VSUBS 0.007338f
C417 B.n377 VSUBS 0.007338f
C418 B.n378 VSUBS 0.007338f
C419 B.n379 VSUBS 0.007338f
C420 B.n380 VSUBS 0.007338f
C421 B.n381 VSUBS 0.017178f
C422 B.n382 VSUBS 0.016275f
C423 B.n383 VSUBS 0.016275f
C424 B.n384 VSUBS 0.007338f
C425 B.n385 VSUBS 0.007338f
C426 B.n386 VSUBS 0.007338f
C427 B.n387 VSUBS 0.007338f
C428 B.n388 VSUBS 0.007338f
C429 B.n389 VSUBS 0.007338f
C430 B.n390 VSUBS 0.007338f
C431 B.n391 VSUBS 0.007338f
C432 B.n392 VSUBS 0.007338f
C433 B.n393 VSUBS 0.007338f
C434 B.n394 VSUBS 0.007338f
C435 B.n395 VSUBS 0.007338f
C436 B.n396 VSUBS 0.007338f
C437 B.n397 VSUBS 0.007338f
C438 B.n398 VSUBS 0.007338f
C439 B.n399 VSUBS 0.007338f
C440 B.n400 VSUBS 0.007338f
C441 B.n401 VSUBS 0.007338f
C442 B.n402 VSUBS 0.007338f
C443 B.n403 VSUBS 0.007338f
C444 B.n404 VSUBS 0.007338f
C445 B.n405 VSUBS 0.007338f
C446 B.n406 VSUBS 0.007338f
C447 B.n407 VSUBS 0.007338f
C448 B.n408 VSUBS 0.007338f
C449 B.n409 VSUBS 0.007338f
C450 B.n410 VSUBS 0.007338f
C451 B.n411 VSUBS 0.007338f
C452 B.n412 VSUBS 0.007338f
C453 B.n413 VSUBS 0.007338f
C454 B.n414 VSUBS 0.007338f
C455 B.n415 VSUBS 0.007338f
C456 B.n416 VSUBS 0.007338f
C457 B.n417 VSUBS 0.007338f
C458 B.n418 VSUBS 0.007338f
C459 B.n419 VSUBS 0.007338f
C460 B.n420 VSUBS 0.007338f
C461 B.n421 VSUBS 0.007338f
C462 B.n422 VSUBS 0.007338f
C463 B.n423 VSUBS 0.007338f
C464 B.n424 VSUBS 0.007338f
C465 B.n425 VSUBS 0.007338f
C466 B.n426 VSUBS 0.007338f
C467 B.n427 VSUBS 0.007338f
C468 B.n428 VSUBS 0.007338f
C469 B.n429 VSUBS 0.007338f
C470 B.n430 VSUBS 0.007338f
C471 B.n431 VSUBS 0.007338f
C472 B.n432 VSUBS 0.007338f
C473 B.n433 VSUBS 0.007338f
C474 B.n434 VSUBS 0.007338f
C475 B.n435 VSUBS 0.007338f
C476 B.n436 VSUBS 0.007338f
C477 B.n437 VSUBS 0.007338f
C478 B.n438 VSUBS 0.007338f
C479 B.n439 VSUBS 0.007338f
C480 B.n440 VSUBS 0.007338f
C481 B.n441 VSUBS 0.007338f
C482 B.n442 VSUBS 0.007338f
C483 B.n443 VSUBS 0.007338f
C484 B.n444 VSUBS 0.007338f
C485 B.n445 VSUBS 0.007338f
C486 B.n446 VSUBS 0.007338f
C487 B.n447 VSUBS 0.007338f
C488 B.n448 VSUBS 0.007338f
C489 B.n449 VSUBS 0.007338f
C490 B.n450 VSUBS 0.007338f
C491 B.n451 VSUBS 0.007338f
C492 B.n452 VSUBS 0.007338f
C493 B.n453 VSUBS 0.007338f
C494 B.n454 VSUBS 0.007338f
C495 B.n455 VSUBS 0.007338f
C496 B.n456 VSUBS 0.007338f
C497 B.n457 VSUBS 0.007338f
C498 B.n458 VSUBS 0.007338f
C499 B.n459 VSUBS 0.007338f
C500 B.n460 VSUBS 0.007338f
C501 B.n461 VSUBS 0.007338f
C502 B.n462 VSUBS 0.007338f
C503 B.n463 VSUBS 0.007338f
C504 B.n464 VSUBS 0.007338f
C505 B.n465 VSUBS 0.007338f
C506 B.n466 VSUBS 0.007338f
C507 B.n467 VSUBS 0.007338f
C508 B.n468 VSUBS 0.007338f
C509 B.n469 VSUBS 0.007338f
C510 B.n470 VSUBS 0.007338f
C511 B.n471 VSUBS 0.007338f
C512 B.n472 VSUBS 0.007338f
C513 B.n473 VSUBS 0.007338f
C514 B.n474 VSUBS 0.007338f
C515 B.n475 VSUBS 0.007338f
C516 B.n476 VSUBS 0.007338f
C517 B.n477 VSUBS 0.007338f
C518 B.n478 VSUBS 0.007338f
C519 B.n479 VSUBS 0.007338f
C520 B.n480 VSUBS 0.007338f
C521 B.n481 VSUBS 0.016275f
C522 B.n482 VSUBS 0.017178f
C523 B.n483 VSUBS 0.016275f
C524 B.n484 VSUBS 0.007338f
C525 B.n485 VSUBS 0.007338f
C526 B.n486 VSUBS 0.007338f
C527 B.n487 VSUBS 0.007338f
C528 B.n488 VSUBS 0.007338f
C529 B.n489 VSUBS 0.007338f
C530 B.n490 VSUBS 0.007338f
C531 B.n491 VSUBS 0.007338f
C532 B.n492 VSUBS 0.007338f
C533 B.n493 VSUBS 0.007338f
C534 B.n494 VSUBS 0.007338f
C535 B.n495 VSUBS 0.007338f
C536 B.n496 VSUBS 0.007338f
C537 B.n497 VSUBS 0.007338f
C538 B.n498 VSUBS 0.007338f
C539 B.n499 VSUBS 0.007338f
C540 B.n500 VSUBS 0.007338f
C541 B.n501 VSUBS 0.007338f
C542 B.n502 VSUBS 0.007338f
C543 B.n503 VSUBS 0.007338f
C544 B.n504 VSUBS 0.007338f
C545 B.n505 VSUBS 0.007338f
C546 B.n506 VSUBS 0.007338f
C547 B.n507 VSUBS 0.007338f
C548 B.n508 VSUBS 0.007338f
C549 B.n509 VSUBS 0.007338f
C550 B.n510 VSUBS 0.007338f
C551 B.n511 VSUBS 0.007338f
C552 B.n512 VSUBS 0.007338f
C553 B.n513 VSUBS 0.007338f
C554 B.n514 VSUBS 0.007338f
C555 B.n515 VSUBS 0.007338f
C556 B.n516 VSUBS 0.007338f
C557 B.n517 VSUBS 0.007338f
C558 B.n518 VSUBS 0.007338f
C559 B.n519 VSUBS 0.007338f
C560 B.n520 VSUBS 0.007338f
C561 B.n521 VSUBS 0.007338f
C562 B.n522 VSUBS 0.007338f
C563 B.n523 VSUBS 0.007338f
C564 B.n524 VSUBS 0.007338f
C565 B.n525 VSUBS 0.007338f
C566 B.n526 VSUBS 0.007338f
C567 B.n527 VSUBS 0.007338f
C568 B.n528 VSUBS 0.007338f
C569 B.n529 VSUBS 0.007338f
C570 B.n530 VSUBS 0.007338f
C571 B.n531 VSUBS 0.007338f
C572 B.n532 VSUBS 0.007338f
C573 B.n533 VSUBS 0.007338f
C574 B.n534 VSUBS 0.007338f
C575 B.n535 VSUBS 0.007338f
C576 B.n536 VSUBS 0.007338f
C577 B.n537 VSUBS 0.007338f
C578 B.n538 VSUBS 0.007338f
C579 B.n539 VSUBS 0.007338f
C580 B.n540 VSUBS 0.007338f
C581 B.n541 VSUBS 0.007338f
C582 B.n542 VSUBS 0.007338f
C583 B.n543 VSUBS 0.007338f
C584 B.n544 VSUBS 0.007338f
C585 B.n545 VSUBS 0.007338f
C586 B.n546 VSUBS 0.007338f
C587 B.n547 VSUBS 0.007338f
C588 B.n548 VSUBS 0.007338f
C589 B.n549 VSUBS 0.007338f
C590 B.n550 VSUBS 0.006906f
C591 B.n551 VSUBS 0.007338f
C592 B.n552 VSUBS 0.007338f
C593 B.n553 VSUBS 0.007338f
C594 B.n554 VSUBS 0.007338f
C595 B.n555 VSUBS 0.007338f
C596 B.n556 VSUBS 0.007338f
C597 B.n557 VSUBS 0.007338f
C598 B.n558 VSUBS 0.007338f
C599 B.n559 VSUBS 0.007338f
C600 B.n560 VSUBS 0.007338f
C601 B.n561 VSUBS 0.007338f
C602 B.n562 VSUBS 0.007338f
C603 B.n563 VSUBS 0.007338f
C604 B.n564 VSUBS 0.007338f
C605 B.n565 VSUBS 0.007338f
C606 B.n566 VSUBS 0.004101f
C607 B.n567 VSUBS 0.017002f
C608 B.n568 VSUBS 0.006906f
C609 B.n569 VSUBS 0.007338f
C610 B.n570 VSUBS 0.007338f
C611 B.n571 VSUBS 0.007338f
C612 B.n572 VSUBS 0.007338f
C613 B.n573 VSUBS 0.007338f
C614 B.n574 VSUBS 0.007338f
C615 B.n575 VSUBS 0.007338f
C616 B.n576 VSUBS 0.007338f
C617 B.n577 VSUBS 0.007338f
C618 B.n578 VSUBS 0.007338f
C619 B.n579 VSUBS 0.007338f
C620 B.n580 VSUBS 0.007338f
C621 B.n581 VSUBS 0.007338f
C622 B.n582 VSUBS 0.007338f
C623 B.n583 VSUBS 0.007338f
C624 B.n584 VSUBS 0.007338f
C625 B.n585 VSUBS 0.007338f
C626 B.n586 VSUBS 0.007338f
C627 B.n587 VSUBS 0.007338f
C628 B.n588 VSUBS 0.007338f
C629 B.n589 VSUBS 0.007338f
C630 B.n590 VSUBS 0.007338f
C631 B.n591 VSUBS 0.007338f
C632 B.n592 VSUBS 0.007338f
C633 B.n593 VSUBS 0.007338f
C634 B.n594 VSUBS 0.007338f
C635 B.n595 VSUBS 0.007338f
C636 B.n596 VSUBS 0.007338f
C637 B.n597 VSUBS 0.007338f
C638 B.n598 VSUBS 0.007338f
C639 B.n599 VSUBS 0.007338f
C640 B.n600 VSUBS 0.007338f
C641 B.n601 VSUBS 0.007338f
C642 B.n602 VSUBS 0.007338f
C643 B.n603 VSUBS 0.007338f
C644 B.n604 VSUBS 0.007338f
C645 B.n605 VSUBS 0.007338f
C646 B.n606 VSUBS 0.007338f
C647 B.n607 VSUBS 0.007338f
C648 B.n608 VSUBS 0.007338f
C649 B.n609 VSUBS 0.007338f
C650 B.n610 VSUBS 0.007338f
C651 B.n611 VSUBS 0.007338f
C652 B.n612 VSUBS 0.007338f
C653 B.n613 VSUBS 0.007338f
C654 B.n614 VSUBS 0.007338f
C655 B.n615 VSUBS 0.007338f
C656 B.n616 VSUBS 0.007338f
C657 B.n617 VSUBS 0.007338f
C658 B.n618 VSUBS 0.007338f
C659 B.n619 VSUBS 0.007338f
C660 B.n620 VSUBS 0.007338f
C661 B.n621 VSUBS 0.007338f
C662 B.n622 VSUBS 0.007338f
C663 B.n623 VSUBS 0.007338f
C664 B.n624 VSUBS 0.007338f
C665 B.n625 VSUBS 0.007338f
C666 B.n626 VSUBS 0.007338f
C667 B.n627 VSUBS 0.007338f
C668 B.n628 VSUBS 0.007338f
C669 B.n629 VSUBS 0.007338f
C670 B.n630 VSUBS 0.007338f
C671 B.n631 VSUBS 0.007338f
C672 B.n632 VSUBS 0.007338f
C673 B.n633 VSUBS 0.007338f
C674 B.n634 VSUBS 0.007338f
C675 B.n635 VSUBS 0.017178f
C676 B.n636 VSUBS 0.017178f
C677 B.n637 VSUBS 0.016275f
C678 B.n638 VSUBS 0.007338f
C679 B.n639 VSUBS 0.007338f
C680 B.n640 VSUBS 0.007338f
C681 B.n641 VSUBS 0.007338f
C682 B.n642 VSUBS 0.007338f
C683 B.n643 VSUBS 0.007338f
C684 B.n644 VSUBS 0.007338f
C685 B.n645 VSUBS 0.007338f
C686 B.n646 VSUBS 0.007338f
C687 B.n647 VSUBS 0.007338f
C688 B.n648 VSUBS 0.007338f
C689 B.n649 VSUBS 0.007338f
C690 B.n650 VSUBS 0.007338f
C691 B.n651 VSUBS 0.007338f
C692 B.n652 VSUBS 0.007338f
C693 B.n653 VSUBS 0.007338f
C694 B.n654 VSUBS 0.007338f
C695 B.n655 VSUBS 0.007338f
C696 B.n656 VSUBS 0.007338f
C697 B.n657 VSUBS 0.007338f
C698 B.n658 VSUBS 0.007338f
C699 B.n659 VSUBS 0.007338f
C700 B.n660 VSUBS 0.007338f
C701 B.n661 VSUBS 0.007338f
C702 B.n662 VSUBS 0.007338f
C703 B.n663 VSUBS 0.007338f
C704 B.n664 VSUBS 0.007338f
C705 B.n665 VSUBS 0.007338f
C706 B.n666 VSUBS 0.007338f
C707 B.n667 VSUBS 0.007338f
C708 B.n668 VSUBS 0.007338f
C709 B.n669 VSUBS 0.007338f
C710 B.n670 VSUBS 0.007338f
C711 B.n671 VSUBS 0.007338f
C712 B.n672 VSUBS 0.007338f
C713 B.n673 VSUBS 0.007338f
C714 B.n674 VSUBS 0.007338f
C715 B.n675 VSUBS 0.007338f
C716 B.n676 VSUBS 0.007338f
C717 B.n677 VSUBS 0.007338f
C718 B.n678 VSUBS 0.007338f
C719 B.n679 VSUBS 0.007338f
C720 B.n680 VSUBS 0.007338f
C721 B.n681 VSUBS 0.007338f
C722 B.n682 VSUBS 0.007338f
C723 B.n683 VSUBS 0.007338f
C724 B.n684 VSUBS 0.007338f
C725 B.n685 VSUBS 0.007338f
C726 B.n686 VSUBS 0.007338f
C727 B.n687 VSUBS 0.016616f
C728 VDD2.t1 VSUBS 0.269692f
C729 VDD2.t7 VSUBS 0.269692f
C730 VDD2.n0 VSUBS 2.15028f
C731 VDD2.t2 VSUBS 0.269692f
C732 VDD2.t4 VSUBS 0.269692f
C733 VDD2.n1 VSUBS 2.15028f
C734 VDD2.n2 VSUBS 3.22789f
C735 VDD2.t0 VSUBS 0.269692f
C736 VDD2.t5 VSUBS 0.269692f
C737 VDD2.n3 VSUBS 2.14408f
C738 VDD2.n4 VSUBS 2.93839f
C739 VDD2.t6 VSUBS 0.269692f
C740 VDD2.t3 VSUBS 0.269692f
C741 VDD2.n5 VSUBS 2.15025f
C742 VN.n0 VSUBS 0.039477f
C743 VN.t3 VSUBS 1.9871f
C744 VN.n1 VSUBS 0.068038f
C745 VN.n2 VSUBS 0.039477f
C746 VN.n3 VSUBS 0.043933f
C747 VN.t6 VSUBS 2.08182f
C748 VN.t0 VSUBS 1.9871f
C749 VN.n4 VSUBS 0.770812f
C750 VN.n5 VSUBS 0.811084f
C751 VN.n6 VSUBS 0.210949f
C752 VN.n7 VSUBS 0.039477f
C753 VN.n8 VSUBS 0.057386f
C754 VN.n9 VSUBS 0.057386f
C755 VN.t5 VSUBS 1.9871f
C756 VN.n10 VSUBS 0.715225f
C757 VN.n11 VSUBS 0.043933f
C758 VN.n12 VSUBS 0.039477f
C759 VN.n13 VSUBS 0.039477f
C760 VN.n14 VSUBS 0.039477f
C761 VN.n15 VSUBS 0.033734f
C762 VN.n16 VSUBS 0.0638f
C763 VN.n17 VSUBS 0.793764f
C764 VN.n18 VSUBS 0.035742f
C765 VN.n19 VSUBS 0.039477f
C766 VN.t7 VSUBS 1.9871f
C767 VN.n20 VSUBS 0.068038f
C768 VN.n21 VSUBS 0.039477f
C769 VN.t2 VSUBS 1.9871f
C770 VN.n22 VSUBS 0.715225f
C771 VN.n23 VSUBS 0.043933f
C772 VN.t4 VSUBS 2.08182f
C773 VN.t1 VSUBS 1.9871f
C774 VN.n24 VSUBS 0.770812f
C775 VN.n25 VSUBS 0.811084f
C776 VN.n26 VSUBS 0.210949f
C777 VN.n27 VSUBS 0.039477f
C778 VN.n28 VSUBS 0.057386f
C779 VN.n29 VSUBS 0.057386f
C780 VN.n30 VSUBS 0.043933f
C781 VN.n31 VSUBS 0.039477f
C782 VN.n32 VSUBS 0.039477f
C783 VN.n33 VSUBS 0.039477f
C784 VN.n34 VSUBS 0.033734f
C785 VN.n35 VSUBS 0.0638f
C786 VN.n36 VSUBS 0.793764f
C787 VN.n37 VSUBS 1.9326f
C788 VTAIL.t2 VSUBS 0.256028f
C789 VTAIL.t5 VSUBS 0.256028f
C790 VTAIL.n0 VSUBS 1.89737f
C791 VTAIL.n1 VSUBS 0.683955f
C792 VTAIL.n2 VSUBS 0.026801f
C793 VTAIL.n3 VSUBS 0.023928f
C794 VTAIL.n4 VSUBS 0.012858f
C795 VTAIL.n5 VSUBS 0.030392f
C796 VTAIL.n6 VSUBS 0.013614f
C797 VTAIL.n7 VSUBS 0.023928f
C798 VTAIL.n8 VSUBS 0.012858f
C799 VTAIL.n9 VSUBS 0.030392f
C800 VTAIL.n10 VSUBS 0.013614f
C801 VTAIL.n11 VSUBS 0.023928f
C802 VTAIL.n12 VSUBS 0.012858f
C803 VTAIL.n13 VSUBS 0.030392f
C804 VTAIL.n14 VSUBS 0.013236f
C805 VTAIL.n15 VSUBS 0.023928f
C806 VTAIL.n16 VSUBS 0.013614f
C807 VTAIL.n17 VSUBS 0.030392f
C808 VTAIL.n18 VSUBS 0.013614f
C809 VTAIL.n19 VSUBS 0.023928f
C810 VTAIL.n20 VSUBS 0.012858f
C811 VTAIL.n21 VSUBS 0.030392f
C812 VTAIL.n22 VSUBS 0.013614f
C813 VTAIL.n23 VSUBS 1.33715f
C814 VTAIL.n24 VSUBS 0.012858f
C815 VTAIL.t0 VSUBS 0.065613f
C816 VTAIL.n25 VSUBS 0.205111f
C817 VTAIL.n26 VSUBS 0.022862f
C818 VTAIL.n27 VSUBS 0.022794f
C819 VTAIL.n28 VSUBS 0.030392f
C820 VTAIL.n29 VSUBS 0.013614f
C821 VTAIL.n30 VSUBS 0.012858f
C822 VTAIL.n31 VSUBS 0.023928f
C823 VTAIL.n32 VSUBS 0.023928f
C824 VTAIL.n33 VSUBS 0.012858f
C825 VTAIL.n34 VSUBS 0.013614f
C826 VTAIL.n35 VSUBS 0.030392f
C827 VTAIL.n36 VSUBS 0.030392f
C828 VTAIL.n37 VSUBS 0.013614f
C829 VTAIL.n38 VSUBS 0.012858f
C830 VTAIL.n39 VSUBS 0.023928f
C831 VTAIL.n40 VSUBS 0.023928f
C832 VTAIL.n41 VSUBS 0.012858f
C833 VTAIL.n42 VSUBS 0.012858f
C834 VTAIL.n43 VSUBS 0.013614f
C835 VTAIL.n44 VSUBS 0.030392f
C836 VTAIL.n45 VSUBS 0.030392f
C837 VTAIL.n46 VSUBS 0.030392f
C838 VTAIL.n47 VSUBS 0.013236f
C839 VTAIL.n48 VSUBS 0.012858f
C840 VTAIL.n49 VSUBS 0.023928f
C841 VTAIL.n50 VSUBS 0.023928f
C842 VTAIL.n51 VSUBS 0.012858f
C843 VTAIL.n52 VSUBS 0.013614f
C844 VTAIL.n53 VSUBS 0.030392f
C845 VTAIL.n54 VSUBS 0.030392f
C846 VTAIL.n55 VSUBS 0.013614f
C847 VTAIL.n56 VSUBS 0.012858f
C848 VTAIL.n57 VSUBS 0.023928f
C849 VTAIL.n58 VSUBS 0.023928f
C850 VTAIL.n59 VSUBS 0.012858f
C851 VTAIL.n60 VSUBS 0.013614f
C852 VTAIL.n61 VSUBS 0.030392f
C853 VTAIL.n62 VSUBS 0.030392f
C854 VTAIL.n63 VSUBS 0.013614f
C855 VTAIL.n64 VSUBS 0.012858f
C856 VTAIL.n65 VSUBS 0.023928f
C857 VTAIL.n66 VSUBS 0.023928f
C858 VTAIL.n67 VSUBS 0.012858f
C859 VTAIL.n68 VSUBS 0.013614f
C860 VTAIL.n69 VSUBS 0.030392f
C861 VTAIL.n70 VSUBS 0.075308f
C862 VTAIL.n71 VSUBS 0.013614f
C863 VTAIL.n72 VSUBS 0.012858f
C864 VTAIL.n73 VSUBS 0.054656f
C865 VTAIL.n74 VSUBS 0.037928f
C866 VTAIL.n75 VSUBS 0.168624f
C867 VTAIL.n76 VSUBS 0.026801f
C868 VTAIL.n77 VSUBS 0.023928f
C869 VTAIL.n78 VSUBS 0.012858f
C870 VTAIL.n79 VSUBS 0.030392f
C871 VTAIL.n80 VSUBS 0.013614f
C872 VTAIL.n81 VSUBS 0.023928f
C873 VTAIL.n82 VSUBS 0.012858f
C874 VTAIL.n83 VSUBS 0.030392f
C875 VTAIL.n84 VSUBS 0.013614f
C876 VTAIL.n85 VSUBS 0.023928f
C877 VTAIL.n86 VSUBS 0.012858f
C878 VTAIL.n87 VSUBS 0.030392f
C879 VTAIL.n88 VSUBS 0.013236f
C880 VTAIL.n89 VSUBS 0.023928f
C881 VTAIL.n90 VSUBS 0.013614f
C882 VTAIL.n91 VSUBS 0.030392f
C883 VTAIL.n92 VSUBS 0.013614f
C884 VTAIL.n93 VSUBS 0.023928f
C885 VTAIL.n94 VSUBS 0.012858f
C886 VTAIL.n95 VSUBS 0.030392f
C887 VTAIL.n96 VSUBS 0.013614f
C888 VTAIL.n97 VSUBS 1.33715f
C889 VTAIL.n98 VSUBS 0.012858f
C890 VTAIL.t12 VSUBS 0.065613f
C891 VTAIL.n99 VSUBS 0.205111f
C892 VTAIL.n100 VSUBS 0.022862f
C893 VTAIL.n101 VSUBS 0.022794f
C894 VTAIL.n102 VSUBS 0.030392f
C895 VTAIL.n103 VSUBS 0.013614f
C896 VTAIL.n104 VSUBS 0.012858f
C897 VTAIL.n105 VSUBS 0.023928f
C898 VTAIL.n106 VSUBS 0.023928f
C899 VTAIL.n107 VSUBS 0.012858f
C900 VTAIL.n108 VSUBS 0.013614f
C901 VTAIL.n109 VSUBS 0.030392f
C902 VTAIL.n110 VSUBS 0.030392f
C903 VTAIL.n111 VSUBS 0.013614f
C904 VTAIL.n112 VSUBS 0.012858f
C905 VTAIL.n113 VSUBS 0.023928f
C906 VTAIL.n114 VSUBS 0.023928f
C907 VTAIL.n115 VSUBS 0.012858f
C908 VTAIL.n116 VSUBS 0.012858f
C909 VTAIL.n117 VSUBS 0.013614f
C910 VTAIL.n118 VSUBS 0.030392f
C911 VTAIL.n119 VSUBS 0.030392f
C912 VTAIL.n120 VSUBS 0.030392f
C913 VTAIL.n121 VSUBS 0.013236f
C914 VTAIL.n122 VSUBS 0.012858f
C915 VTAIL.n123 VSUBS 0.023928f
C916 VTAIL.n124 VSUBS 0.023928f
C917 VTAIL.n125 VSUBS 0.012858f
C918 VTAIL.n126 VSUBS 0.013614f
C919 VTAIL.n127 VSUBS 0.030392f
C920 VTAIL.n128 VSUBS 0.030392f
C921 VTAIL.n129 VSUBS 0.013614f
C922 VTAIL.n130 VSUBS 0.012858f
C923 VTAIL.n131 VSUBS 0.023928f
C924 VTAIL.n132 VSUBS 0.023928f
C925 VTAIL.n133 VSUBS 0.012858f
C926 VTAIL.n134 VSUBS 0.013614f
C927 VTAIL.n135 VSUBS 0.030392f
C928 VTAIL.n136 VSUBS 0.030392f
C929 VTAIL.n137 VSUBS 0.013614f
C930 VTAIL.n138 VSUBS 0.012858f
C931 VTAIL.n139 VSUBS 0.023928f
C932 VTAIL.n140 VSUBS 0.023928f
C933 VTAIL.n141 VSUBS 0.012858f
C934 VTAIL.n142 VSUBS 0.013614f
C935 VTAIL.n143 VSUBS 0.030392f
C936 VTAIL.n144 VSUBS 0.075308f
C937 VTAIL.n145 VSUBS 0.013614f
C938 VTAIL.n146 VSUBS 0.012858f
C939 VTAIL.n147 VSUBS 0.054656f
C940 VTAIL.n148 VSUBS 0.037928f
C941 VTAIL.n149 VSUBS 0.168624f
C942 VTAIL.t11 VSUBS 0.256028f
C943 VTAIL.t10 VSUBS 0.256028f
C944 VTAIL.n150 VSUBS 1.89737f
C945 VTAIL.n151 VSUBS 0.791799f
C946 VTAIL.n152 VSUBS 0.026801f
C947 VTAIL.n153 VSUBS 0.023928f
C948 VTAIL.n154 VSUBS 0.012858f
C949 VTAIL.n155 VSUBS 0.030392f
C950 VTAIL.n156 VSUBS 0.013614f
C951 VTAIL.n157 VSUBS 0.023928f
C952 VTAIL.n158 VSUBS 0.012858f
C953 VTAIL.n159 VSUBS 0.030392f
C954 VTAIL.n160 VSUBS 0.013614f
C955 VTAIL.n161 VSUBS 0.023928f
C956 VTAIL.n162 VSUBS 0.012858f
C957 VTAIL.n163 VSUBS 0.030392f
C958 VTAIL.n164 VSUBS 0.013236f
C959 VTAIL.n165 VSUBS 0.023928f
C960 VTAIL.n166 VSUBS 0.013614f
C961 VTAIL.n167 VSUBS 0.030392f
C962 VTAIL.n168 VSUBS 0.013614f
C963 VTAIL.n169 VSUBS 0.023928f
C964 VTAIL.n170 VSUBS 0.012858f
C965 VTAIL.n171 VSUBS 0.030392f
C966 VTAIL.n172 VSUBS 0.013614f
C967 VTAIL.n173 VSUBS 1.33715f
C968 VTAIL.n174 VSUBS 0.012858f
C969 VTAIL.t15 VSUBS 0.065613f
C970 VTAIL.n175 VSUBS 0.205111f
C971 VTAIL.n176 VSUBS 0.022862f
C972 VTAIL.n177 VSUBS 0.022794f
C973 VTAIL.n178 VSUBS 0.030392f
C974 VTAIL.n179 VSUBS 0.013614f
C975 VTAIL.n180 VSUBS 0.012858f
C976 VTAIL.n181 VSUBS 0.023928f
C977 VTAIL.n182 VSUBS 0.023928f
C978 VTAIL.n183 VSUBS 0.012858f
C979 VTAIL.n184 VSUBS 0.013614f
C980 VTAIL.n185 VSUBS 0.030392f
C981 VTAIL.n186 VSUBS 0.030392f
C982 VTAIL.n187 VSUBS 0.013614f
C983 VTAIL.n188 VSUBS 0.012858f
C984 VTAIL.n189 VSUBS 0.023928f
C985 VTAIL.n190 VSUBS 0.023928f
C986 VTAIL.n191 VSUBS 0.012858f
C987 VTAIL.n192 VSUBS 0.012858f
C988 VTAIL.n193 VSUBS 0.013614f
C989 VTAIL.n194 VSUBS 0.030392f
C990 VTAIL.n195 VSUBS 0.030392f
C991 VTAIL.n196 VSUBS 0.030392f
C992 VTAIL.n197 VSUBS 0.013236f
C993 VTAIL.n198 VSUBS 0.012858f
C994 VTAIL.n199 VSUBS 0.023928f
C995 VTAIL.n200 VSUBS 0.023928f
C996 VTAIL.n201 VSUBS 0.012858f
C997 VTAIL.n202 VSUBS 0.013614f
C998 VTAIL.n203 VSUBS 0.030392f
C999 VTAIL.n204 VSUBS 0.030392f
C1000 VTAIL.n205 VSUBS 0.013614f
C1001 VTAIL.n206 VSUBS 0.012858f
C1002 VTAIL.n207 VSUBS 0.023928f
C1003 VTAIL.n208 VSUBS 0.023928f
C1004 VTAIL.n209 VSUBS 0.012858f
C1005 VTAIL.n210 VSUBS 0.013614f
C1006 VTAIL.n211 VSUBS 0.030392f
C1007 VTAIL.n212 VSUBS 0.030392f
C1008 VTAIL.n213 VSUBS 0.013614f
C1009 VTAIL.n214 VSUBS 0.012858f
C1010 VTAIL.n215 VSUBS 0.023928f
C1011 VTAIL.n216 VSUBS 0.023928f
C1012 VTAIL.n217 VSUBS 0.012858f
C1013 VTAIL.n218 VSUBS 0.013614f
C1014 VTAIL.n219 VSUBS 0.030392f
C1015 VTAIL.n220 VSUBS 0.075308f
C1016 VTAIL.n221 VSUBS 0.013614f
C1017 VTAIL.n222 VSUBS 0.012858f
C1018 VTAIL.n223 VSUBS 0.054656f
C1019 VTAIL.n224 VSUBS 0.037928f
C1020 VTAIL.n225 VSUBS 1.46975f
C1021 VTAIL.n226 VSUBS 0.026801f
C1022 VTAIL.n227 VSUBS 0.023928f
C1023 VTAIL.n228 VSUBS 0.012858f
C1024 VTAIL.n229 VSUBS 0.030392f
C1025 VTAIL.n230 VSUBS 0.013614f
C1026 VTAIL.n231 VSUBS 0.023928f
C1027 VTAIL.n232 VSUBS 0.012858f
C1028 VTAIL.n233 VSUBS 0.030392f
C1029 VTAIL.n234 VSUBS 0.013614f
C1030 VTAIL.n235 VSUBS 0.023928f
C1031 VTAIL.n236 VSUBS 0.012858f
C1032 VTAIL.n237 VSUBS 0.030392f
C1033 VTAIL.n238 VSUBS 0.013236f
C1034 VTAIL.n239 VSUBS 0.023928f
C1035 VTAIL.n240 VSUBS 0.013236f
C1036 VTAIL.n241 VSUBS 0.012858f
C1037 VTAIL.n242 VSUBS 0.030392f
C1038 VTAIL.n243 VSUBS 0.030392f
C1039 VTAIL.n244 VSUBS 0.013614f
C1040 VTAIL.n245 VSUBS 0.023928f
C1041 VTAIL.n246 VSUBS 0.012858f
C1042 VTAIL.n247 VSUBS 0.030392f
C1043 VTAIL.n248 VSUBS 0.013614f
C1044 VTAIL.n249 VSUBS 1.33715f
C1045 VTAIL.n250 VSUBS 0.012858f
C1046 VTAIL.t6 VSUBS 0.065613f
C1047 VTAIL.n251 VSUBS 0.205111f
C1048 VTAIL.n252 VSUBS 0.022862f
C1049 VTAIL.n253 VSUBS 0.022794f
C1050 VTAIL.n254 VSUBS 0.030392f
C1051 VTAIL.n255 VSUBS 0.013614f
C1052 VTAIL.n256 VSUBS 0.012858f
C1053 VTAIL.n257 VSUBS 0.023928f
C1054 VTAIL.n258 VSUBS 0.023928f
C1055 VTAIL.n259 VSUBS 0.012858f
C1056 VTAIL.n260 VSUBS 0.013614f
C1057 VTAIL.n261 VSUBS 0.030392f
C1058 VTAIL.n262 VSUBS 0.030392f
C1059 VTAIL.n263 VSUBS 0.013614f
C1060 VTAIL.n264 VSUBS 0.012858f
C1061 VTAIL.n265 VSUBS 0.023928f
C1062 VTAIL.n266 VSUBS 0.023928f
C1063 VTAIL.n267 VSUBS 0.012858f
C1064 VTAIL.n268 VSUBS 0.013614f
C1065 VTAIL.n269 VSUBS 0.030392f
C1066 VTAIL.n270 VSUBS 0.030392f
C1067 VTAIL.n271 VSUBS 0.013614f
C1068 VTAIL.n272 VSUBS 0.012858f
C1069 VTAIL.n273 VSUBS 0.023928f
C1070 VTAIL.n274 VSUBS 0.023928f
C1071 VTAIL.n275 VSUBS 0.012858f
C1072 VTAIL.n276 VSUBS 0.013614f
C1073 VTAIL.n277 VSUBS 0.030392f
C1074 VTAIL.n278 VSUBS 0.030392f
C1075 VTAIL.n279 VSUBS 0.013614f
C1076 VTAIL.n280 VSUBS 0.012858f
C1077 VTAIL.n281 VSUBS 0.023928f
C1078 VTAIL.n282 VSUBS 0.023928f
C1079 VTAIL.n283 VSUBS 0.012858f
C1080 VTAIL.n284 VSUBS 0.013614f
C1081 VTAIL.n285 VSUBS 0.030392f
C1082 VTAIL.n286 VSUBS 0.030392f
C1083 VTAIL.n287 VSUBS 0.013614f
C1084 VTAIL.n288 VSUBS 0.012858f
C1085 VTAIL.n289 VSUBS 0.023928f
C1086 VTAIL.n290 VSUBS 0.023928f
C1087 VTAIL.n291 VSUBS 0.012858f
C1088 VTAIL.n292 VSUBS 0.013614f
C1089 VTAIL.n293 VSUBS 0.030392f
C1090 VTAIL.n294 VSUBS 0.075308f
C1091 VTAIL.n295 VSUBS 0.013614f
C1092 VTAIL.n296 VSUBS 0.012858f
C1093 VTAIL.n297 VSUBS 0.054656f
C1094 VTAIL.n298 VSUBS 0.037928f
C1095 VTAIL.n299 VSUBS 1.46975f
C1096 VTAIL.t7 VSUBS 0.256028f
C1097 VTAIL.t4 VSUBS 0.256028f
C1098 VTAIL.n300 VSUBS 1.89739f
C1099 VTAIL.n301 VSUBS 0.791787f
C1100 VTAIL.n302 VSUBS 0.026801f
C1101 VTAIL.n303 VSUBS 0.023928f
C1102 VTAIL.n304 VSUBS 0.012858f
C1103 VTAIL.n305 VSUBS 0.030392f
C1104 VTAIL.n306 VSUBS 0.013614f
C1105 VTAIL.n307 VSUBS 0.023928f
C1106 VTAIL.n308 VSUBS 0.012858f
C1107 VTAIL.n309 VSUBS 0.030392f
C1108 VTAIL.n310 VSUBS 0.013614f
C1109 VTAIL.n311 VSUBS 0.023928f
C1110 VTAIL.n312 VSUBS 0.012858f
C1111 VTAIL.n313 VSUBS 0.030392f
C1112 VTAIL.n314 VSUBS 0.013236f
C1113 VTAIL.n315 VSUBS 0.023928f
C1114 VTAIL.n316 VSUBS 0.013236f
C1115 VTAIL.n317 VSUBS 0.012858f
C1116 VTAIL.n318 VSUBS 0.030392f
C1117 VTAIL.n319 VSUBS 0.030392f
C1118 VTAIL.n320 VSUBS 0.013614f
C1119 VTAIL.n321 VSUBS 0.023928f
C1120 VTAIL.n322 VSUBS 0.012858f
C1121 VTAIL.n323 VSUBS 0.030392f
C1122 VTAIL.n324 VSUBS 0.013614f
C1123 VTAIL.n325 VSUBS 1.33715f
C1124 VTAIL.n326 VSUBS 0.012858f
C1125 VTAIL.t3 VSUBS 0.065613f
C1126 VTAIL.n327 VSUBS 0.205111f
C1127 VTAIL.n328 VSUBS 0.022862f
C1128 VTAIL.n329 VSUBS 0.022794f
C1129 VTAIL.n330 VSUBS 0.030392f
C1130 VTAIL.n331 VSUBS 0.013614f
C1131 VTAIL.n332 VSUBS 0.012858f
C1132 VTAIL.n333 VSUBS 0.023928f
C1133 VTAIL.n334 VSUBS 0.023928f
C1134 VTAIL.n335 VSUBS 0.012858f
C1135 VTAIL.n336 VSUBS 0.013614f
C1136 VTAIL.n337 VSUBS 0.030392f
C1137 VTAIL.n338 VSUBS 0.030392f
C1138 VTAIL.n339 VSUBS 0.013614f
C1139 VTAIL.n340 VSUBS 0.012858f
C1140 VTAIL.n341 VSUBS 0.023928f
C1141 VTAIL.n342 VSUBS 0.023928f
C1142 VTAIL.n343 VSUBS 0.012858f
C1143 VTAIL.n344 VSUBS 0.013614f
C1144 VTAIL.n345 VSUBS 0.030392f
C1145 VTAIL.n346 VSUBS 0.030392f
C1146 VTAIL.n347 VSUBS 0.013614f
C1147 VTAIL.n348 VSUBS 0.012858f
C1148 VTAIL.n349 VSUBS 0.023928f
C1149 VTAIL.n350 VSUBS 0.023928f
C1150 VTAIL.n351 VSUBS 0.012858f
C1151 VTAIL.n352 VSUBS 0.013614f
C1152 VTAIL.n353 VSUBS 0.030392f
C1153 VTAIL.n354 VSUBS 0.030392f
C1154 VTAIL.n355 VSUBS 0.013614f
C1155 VTAIL.n356 VSUBS 0.012858f
C1156 VTAIL.n357 VSUBS 0.023928f
C1157 VTAIL.n358 VSUBS 0.023928f
C1158 VTAIL.n359 VSUBS 0.012858f
C1159 VTAIL.n360 VSUBS 0.013614f
C1160 VTAIL.n361 VSUBS 0.030392f
C1161 VTAIL.n362 VSUBS 0.030392f
C1162 VTAIL.n363 VSUBS 0.013614f
C1163 VTAIL.n364 VSUBS 0.012858f
C1164 VTAIL.n365 VSUBS 0.023928f
C1165 VTAIL.n366 VSUBS 0.023928f
C1166 VTAIL.n367 VSUBS 0.012858f
C1167 VTAIL.n368 VSUBS 0.013614f
C1168 VTAIL.n369 VSUBS 0.030392f
C1169 VTAIL.n370 VSUBS 0.075308f
C1170 VTAIL.n371 VSUBS 0.013614f
C1171 VTAIL.n372 VSUBS 0.012858f
C1172 VTAIL.n373 VSUBS 0.054656f
C1173 VTAIL.n374 VSUBS 0.037928f
C1174 VTAIL.n375 VSUBS 0.168624f
C1175 VTAIL.n376 VSUBS 0.026801f
C1176 VTAIL.n377 VSUBS 0.023928f
C1177 VTAIL.n378 VSUBS 0.012858f
C1178 VTAIL.n379 VSUBS 0.030392f
C1179 VTAIL.n380 VSUBS 0.013614f
C1180 VTAIL.n381 VSUBS 0.023928f
C1181 VTAIL.n382 VSUBS 0.012858f
C1182 VTAIL.n383 VSUBS 0.030392f
C1183 VTAIL.n384 VSUBS 0.013614f
C1184 VTAIL.n385 VSUBS 0.023928f
C1185 VTAIL.n386 VSUBS 0.012858f
C1186 VTAIL.n387 VSUBS 0.030392f
C1187 VTAIL.n388 VSUBS 0.013236f
C1188 VTAIL.n389 VSUBS 0.023928f
C1189 VTAIL.n390 VSUBS 0.013236f
C1190 VTAIL.n391 VSUBS 0.012858f
C1191 VTAIL.n392 VSUBS 0.030392f
C1192 VTAIL.n393 VSUBS 0.030392f
C1193 VTAIL.n394 VSUBS 0.013614f
C1194 VTAIL.n395 VSUBS 0.023928f
C1195 VTAIL.n396 VSUBS 0.012858f
C1196 VTAIL.n397 VSUBS 0.030392f
C1197 VTAIL.n398 VSUBS 0.013614f
C1198 VTAIL.n399 VSUBS 1.33715f
C1199 VTAIL.n400 VSUBS 0.012858f
C1200 VTAIL.t13 VSUBS 0.065613f
C1201 VTAIL.n401 VSUBS 0.205111f
C1202 VTAIL.n402 VSUBS 0.022862f
C1203 VTAIL.n403 VSUBS 0.022794f
C1204 VTAIL.n404 VSUBS 0.030392f
C1205 VTAIL.n405 VSUBS 0.013614f
C1206 VTAIL.n406 VSUBS 0.012858f
C1207 VTAIL.n407 VSUBS 0.023928f
C1208 VTAIL.n408 VSUBS 0.023928f
C1209 VTAIL.n409 VSUBS 0.012858f
C1210 VTAIL.n410 VSUBS 0.013614f
C1211 VTAIL.n411 VSUBS 0.030392f
C1212 VTAIL.n412 VSUBS 0.030392f
C1213 VTAIL.n413 VSUBS 0.013614f
C1214 VTAIL.n414 VSUBS 0.012858f
C1215 VTAIL.n415 VSUBS 0.023928f
C1216 VTAIL.n416 VSUBS 0.023928f
C1217 VTAIL.n417 VSUBS 0.012858f
C1218 VTAIL.n418 VSUBS 0.013614f
C1219 VTAIL.n419 VSUBS 0.030392f
C1220 VTAIL.n420 VSUBS 0.030392f
C1221 VTAIL.n421 VSUBS 0.013614f
C1222 VTAIL.n422 VSUBS 0.012858f
C1223 VTAIL.n423 VSUBS 0.023928f
C1224 VTAIL.n424 VSUBS 0.023928f
C1225 VTAIL.n425 VSUBS 0.012858f
C1226 VTAIL.n426 VSUBS 0.013614f
C1227 VTAIL.n427 VSUBS 0.030392f
C1228 VTAIL.n428 VSUBS 0.030392f
C1229 VTAIL.n429 VSUBS 0.013614f
C1230 VTAIL.n430 VSUBS 0.012858f
C1231 VTAIL.n431 VSUBS 0.023928f
C1232 VTAIL.n432 VSUBS 0.023928f
C1233 VTAIL.n433 VSUBS 0.012858f
C1234 VTAIL.n434 VSUBS 0.013614f
C1235 VTAIL.n435 VSUBS 0.030392f
C1236 VTAIL.n436 VSUBS 0.030392f
C1237 VTAIL.n437 VSUBS 0.013614f
C1238 VTAIL.n438 VSUBS 0.012858f
C1239 VTAIL.n439 VSUBS 0.023928f
C1240 VTAIL.n440 VSUBS 0.023928f
C1241 VTAIL.n441 VSUBS 0.012858f
C1242 VTAIL.n442 VSUBS 0.013614f
C1243 VTAIL.n443 VSUBS 0.030392f
C1244 VTAIL.n444 VSUBS 0.075308f
C1245 VTAIL.n445 VSUBS 0.013614f
C1246 VTAIL.n446 VSUBS 0.012858f
C1247 VTAIL.n447 VSUBS 0.054656f
C1248 VTAIL.n448 VSUBS 0.037928f
C1249 VTAIL.n449 VSUBS 0.168624f
C1250 VTAIL.t14 VSUBS 0.256028f
C1251 VTAIL.t8 VSUBS 0.256028f
C1252 VTAIL.n450 VSUBS 1.89739f
C1253 VTAIL.n451 VSUBS 0.791787f
C1254 VTAIL.n452 VSUBS 0.026801f
C1255 VTAIL.n453 VSUBS 0.023928f
C1256 VTAIL.n454 VSUBS 0.012858f
C1257 VTAIL.n455 VSUBS 0.030392f
C1258 VTAIL.n456 VSUBS 0.013614f
C1259 VTAIL.n457 VSUBS 0.023928f
C1260 VTAIL.n458 VSUBS 0.012858f
C1261 VTAIL.n459 VSUBS 0.030392f
C1262 VTAIL.n460 VSUBS 0.013614f
C1263 VTAIL.n461 VSUBS 0.023928f
C1264 VTAIL.n462 VSUBS 0.012858f
C1265 VTAIL.n463 VSUBS 0.030392f
C1266 VTAIL.n464 VSUBS 0.013236f
C1267 VTAIL.n465 VSUBS 0.023928f
C1268 VTAIL.n466 VSUBS 0.013236f
C1269 VTAIL.n467 VSUBS 0.012858f
C1270 VTAIL.n468 VSUBS 0.030392f
C1271 VTAIL.n469 VSUBS 0.030392f
C1272 VTAIL.n470 VSUBS 0.013614f
C1273 VTAIL.n471 VSUBS 0.023928f
C1274 VTAIL.n472 VSUBS 0.012858f
C1275 VTAIL.n473 VSUBS 0.030392f
C1276 VTAIL.n474 VSUBS 0.013614f
C1277 VTAIL.n475 VSUBS 1.33715f
C1278 VTAIL.n476 VSUBS 0.012858f
C1279 VTAIL.t9 VSUBS 0.065613f
C1280 VTAIL.n477 VSUBS 0.205111f
C1281 VTAIL.n478 VSUBS 0.022862f
C1282 VTAIL.n479 VSUBS 0.022794f
C1283 VTAIL.n480 VSUBS 0.030392f
C1284 VTAIL.n481 VSUBS 0.013614f
C1285 VTAIL.n482 VSUBS 0.012858f
C1286 VTAIL.n483 VSUBS 0.023928f
C1287 VTAIL.n484 VSUBS 0.023928f
C1288 VTAIL.n485 VSUBS 0.012858f
C1289 VTAIL.n486 VSUBS 0.013614f
C1290 VTAIL.n487 VSUBS 0.030392f
C1291 VTAIL.n488 VSUBS 0.030392f
C1292 VTAIL.n489 VSUBS 0.013614f
C1293 VTAIL.n490 VSUBS 0.012858f
C1294 VTAIL.n491 VSUBS 0.023928f
C1295 VTAIL.n492 VSUBS 0.023928f
C1296 VTAIL.n493 VSUBS 0.012858f
C1297 VTAIL.n494 VSUBS 0.013614f
C1298 VTAIL.n495 VSUBS 0.030392f
C1299 VTAIL.n496 VSUBS 0.030392f
C1300 VTAIL.n497 VSUBS 0.013614f
C1301 VTAIL.n498 VSUBS 0.012858f
C1302 VTAIL.n499 VSUBS 0.023928f
C1303 VTAIL.n500 VSUBS 0.023928f
C1304 VTAIL.n501 VSUBS 0.012858f
C1305 VTAIL.n502 VSUBS 0.013614f
C1306 VTAIL.n503 VSUBS 0.030392f
C1307 VTAIL.n504 VSUBS 0.030392f
C1308 VTAIL.n505 VSUBS 0.013614f
C1309 VTAIL.n506 VSUBS 0.012858f
C1310 VTAIL.n507 VSUBS 0.023928f
C1311 VTAIL.n508 VSUBS 0.023928f
C1312 VTAIL.n509 VSUBS 0.012858f
C1313 VTAIL.n510 VSUBS 0.013614f
C1314 VTAIL.n511 VSUBS 0.030392f
C1315 VTAIL.n512 VSUBS 0.030392f
C1316 VTAIL.n513 VSUBS 0.013614f
C1317 VTAIL.n514 VSUBS 0.012858f
C1318 VTAIL.n515 VSUBS 0.023928f
C1319 VTAIL.n516 VSUBS 0.023928f
C1320 VTAIL.n517 VSUBS 0.012858f
C1321 VTAIL.n518 VSUBS 0.013614f
C1322 VTAIL.n519 VSUBS 0.030392f
C1323 VTAIL.n520 VSUBS 0.075308f
C1324 VTAIL.n521 VSUBS 0.013614f
C1325 VTAIL.n522 VSUBS 0.012858f
C1326 VTAIL.n523 VSUBS 0.054656f
C1327 VTAIL.n524 VSUBS 0.037928f
C1328 VTAIL.n525 VSUBS 1.46975f
C1329 VTAIL.n526 VSUBS 0.026801f
C1330 VTAIL.n527 VSUBS 0.023928f
C1331 VTAIL.n528 VSUBS 0.012858f
C1332 VTAIL.n529 VSUBS 0.030392f
C1333 VTAIL.n530 VSUBS 0.013614f
C1334 VTAIL.n531 VSUBS 0.023928f
C1335 VTAIL.n532 VSUBS 0.012858f
C1336 VTAIL.n533 VSUBS 0.030392f
C1337 VTAIL.n534 VSUBS 0.013614f
C1338 VTAIL.n535 VSUBS 0.023928f
C1339 VTAIL.n536 VSUBS 0.012858f
C1340 VTAIL.n537 VSUBS 0.030392f
C1341 VTAIL.n538 VSUBS 0.013236f
C1342 VTAIL.n539 VSUBS 0.023928f
C1343 VTAIL.n540 VSUBS 0.013614f
C1344 VTAIL.n541 VSUBS 0.030392f
C1345 VTAIL.n542 VSUBS 0.013614f
C1346 VTAIL.n543 VSUBS 0.023928f
C1347 VTAIL.n544 VSUBS 0.012858f
C1348 VTAIL.n545 VSUBS 0.030392f
C1349 VTAIL.n546 VSUBS 0.013614f
C1350 VTAIL.n547 VSUBS 1.33715f
C1351 VTAIL.n548 VSUBS 0.012858f
C1352 VTAIL.t1 VSUBS 0.065613f
C1353 VTAIL.n549 VSUBS 0.205111f
C1354 VTAIL.n550 VSUBS 0.022862f
C1355 VTAIL.n551 VSUBS 0.022794f
C1356 VTAIL.n552 VSUBS 0.030392f
C1357 VTAIL.n553 VSUBS 0.013614f
C1358 VTAIL.n554 VSUBS 0.012858f
C1359 VTAIL.n555 VSUBS 0.023928f
C1360 VTAIL.n556 VSUBS 0.023928f
C1361 VTAIL.n557 VSUBS 0.012858f
C1362 VTAIL.n558 VSUBS 0.013614f
C1363 VTAIL.n559 VSUBS 0.030392f
C1364 VTAIL.n560 VSUBS 0.030392f
C1365 VTAIL.n561 VSUBS 0.013614f
C1366 VTAIL.n562 VSUBS 0.012858f
C1367 VTAIL.n563 VSUBS 0.023928f
C1368 VTAIL.n564 VSUBS 0.023928f
C1369 VTAIL.n565 VSUBS 0.012858f
C1370 VTAIL.n566 VSUBS 0.012858f
C1371 VTAIL.n567 VSUBS 0.013614f
C1372 VTAIL.n568 VSUBS 0.030392f
C1373 VTAIL.n569 VSUBS 0.030392f
C1374 VTAIL.n570 VSUBS 0.030392f
C1375 VTAIL.n571 VSUBS 0.013236f
C1376 VTAIL.n572 VSUBS 0.012858f
C1377 VTAIL.n573 VSUBS 0.023928f
C1378 VTAIL.n574 VSUBS 0.023928f
C1379 VTAIL.n575 VSUBS 0.012858f
C1380 VTAIL.n576 VSUBS 0.013614f
C1381 VTAIL.n577 VSUBS 0.030392f
C1382 VTAIL.n578 VSUBS 0.030392f
C1383 VTAIL.n579 VSUBS 0.013614f
C1384 VTAIL.n580 VSUBS 0.012858f
C1385 VTAIL.n581 VSUBS 0.023928f
C1386 VTAIL.n582 VSUBS 0.023928f
C1387 VTAIL.n583 VSUBS 0.012858f
C1388 VTAIL.n584 VSUBS 0.013614f
C1389 VTAIL.n585 VSUBS 0.030392f
C1390 VTAIL.n586 VSUBS 0.030392f
C1391 VTAIL.n587 VSUBS 0.013614f
C1392 VTAIL.n588 VSUBS 0.012858f
C1393 VTAIL.n589 VSUBS 0.023928f
C1394 VTAIL.n590 VSUBS 0.023928f
C1395 VTAIL.n591 VSUBS 0.012858f
C1396 VTAIL.n592 VSUBS 0.013614f
C1397 VTAIL.n593 VSUBS 0.030392f
C1398 VTAIL.n594 VSUBS 0.075308f
C1399 VTAIL.n595 VSUBS 0.013614f
C1400 VTAIL.n596 VSUBS 0.012858f
C1401 VTAIL.n597 VSUBS 0.054656f
C1402 VTAIL.n598 VSUBS 0.037928f
C1403 VTAIL.n599 VSUBS 1.46526f
C1404 VDD1.t2 VSUBS 0.271313f
C1405 VDD1.t3 VSUBS 0.271313f
C1406 VDD1.n0 VSUBS 2.16435f
C1407 VDD1.t7 VSUBS 0.271313f
C1408 VDD1.t6 VSUBS 0.271313f
C1409 VDD1.n1 VSUBS 2.1632f
C1410 VDD1.t5 VSUBS 0.271313f
C1411 VDD1.t4 VSUBS 0.271313f
C1412 VDD1.n2 VSUBS 2.1632f
C1413 VDD1.n3 VSUBS 3.30082f
C1414 VDD1.t1 VSUBS 0.271313f
C1415 VDD1.t0 VSUBS 0.271313f
C1416 VDD1.n4 VSUBS 2.15695f
C1417 VDD1.n5 VSUBS 2.98667f
C1418 VP.n0 VSUBS 0.040552f
C1419 VP.t3 VSUBS 2.04121f
C1420 VP.n1 VSUBS 0.069891f
C1421 VP.n2 VSUBS 0.040552f
C1422 VP.n3 VSUBS 0.04513f
C1423 VP.n4 VSUBS 0.040552f
C1424 VP.t0 VSUBS 2.04121f
C1425 VP.n5 VSUBS 0.815378f
C1426 VP.n6 VSUBS 0.040552f
C1427 VP.t6 VSUBS 2.04121f
C1428 VP.n7 VSUBS 0.069891f
C1429 VP.n8 VSUBS 0.040552f
C1430 VP.n9 VSUBS 0.04513f
C1431 VP.t2 VSUBS 2.1385f
C1432 VP.t1 VSUBS 2.04121f
C1433 VP.n10 VSUBS 0.791802f
C1434 VP.n11 VSUBS 0.83317f
C1435 VP.n12 VSUBS 0.216693f
C1436 VP.n13 VSUBS 0.040552f
C1437 VP.n14 VSUBS 0.058949f
C1438 VP.n15 VSUBS 0.058949f
C1439 VP.t7 VSUBS 2.04121f
C1440 VP.n16 VSUBS 0.734701f
C1441 VP.n17 VSUBS 0.04513f
C1442 VP.n18 VSUBS 0.040552f
C1443 VP.n19 VSUBS 0.040552f
C1444 VP.n20 VSUBS 0.040552f
C1445 VP.n21 VSUBS 0.034653f
C1446 VP.n22 VSUBS 0.065537f
C1447 VP.n23 VSUBS 0.815378f
C1448 VP.n24 VSUBS 1.95875f
C1449 VP.n25 VSUBS 1.99039f
C1450 VP.n26 VSUBS 0.040552f
C1451 VP.n27 VSUBS 0.065537f
C1452 VP.n28 VSUBS 0.034653f
C1453 VP.t4 VSUBS 2.04121f
C1454 VP.n29 VSUBS 0.734701f
C1455 VP.n30 VSUBS 0.069891f
C1456 VP.n31 VSUBS 0.040552f
C1457 VP.n32 VSUBS 0.040552f
C1458 VP.n33 VSUBS 0.040552f
C1459 VP.n34 VSUBS 0.058949f
C1460 VP.n35 VSUBS 0.058949f
C1461 VP.t5 VSUBS 2.04121f
C1462 VP.n36 VSUBS 0.734701f
C1463 VP.n37 VSUBS 0.04513f
C1464 VP.n38 VSUBS 0.040552f
C1465 VP.n39 VSUBS 0.040552f
C1466 VP.n40 VSUBS 0.040552f
C1467 VP.n41 VSUBS 0.034653f
C1468 VP.n42 VSUBS 0.065537f
C1469 VP.n43 VSUBS 0.815378f
C1470 VP.n44 VSUBS 0.036716f
.ends

