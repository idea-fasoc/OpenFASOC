* NGSPICE file created from diff_pair_sample_0153.ext - technology: sky130A

.subckt diff_pair_sample_0153 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n3626_n1764# sky130_fd_pr__pfet_01v8 ad=1.5522 pd=8.74 as=0 ps=0 w=3.98 l=2.99
X1 VTAIL.t8 VN.t0 VDD2.t3 w_n3626_n1764# sky130_fd_pr__pfet_01v8 ad=0.6567 pd=4.31 as=0.6567 ps=4.31 w=3.98 l=2.99
X2 VDD1.t5 VP.t0 VTAIL.t9 w_n3626_n1764# sky130_fd_pr__pfet_01v8 ad=1.5522 pd=8.74 as=0.6567 ps=4.31 w=3.98 l=2.99
X3 VDD1.t4 VP.t1 VTAIL.t11 w_n3626_n1764# sky130_fd_pr__pfet_01v8 ad=0.6567 pd=4.31 as=1.5522 ps=8.74 w=3.98 l=2.99
X4 VTAIL.t10 VP.t2 VDD1.t3 w_n3626_n1764# sky130_fd_pr__pfet_01v8 ad=0.6567 pd=4.31 as=0.6567 ps=4.31 w=3.98 l=2.99
X5 VDD2.t4 VN.t1 VTAIL.t7 w_n3626_n1764# sky130_fd_pr__pfet_01v8 ad=0.6567 pd=4.31 as=1.5522 ps=8.74 w=3.98 l=2.99
X6 VDD2.t1 VN.t2 VTAIL.t6 w_n3626_n1764# sky130_fd_pr__pfet_01v8 ad=0.6567 pd=4.31 as=1.5522 ps=8.74 w=3.98 l=2.99
X7 B.t8 B.t6 B.t7 w_n3626_n1764# sky130_fd_pr__pfet_01v8 ad=1.5522 pd=8.74 as=0 ps=0 w=3.98 l=2.99
X8 B.t5 B.t3 B.t4 w_n3626_n1764# sky130_fd_pr__pfet_01v8 ad=1.5522 pd=8.74 as=0 ps=0 w=3.98 l=2.99
X9 VDD2.t5 VN.t3 VTAIL.t5 w_n3626_n1764# sky130_fd_pr__pfet_01v8 ad=1.5522 pd=8.74 as=0.6567 ps=4.31 w=3.98 l=2.99
X10 B.t2 B.t0 B.t1 w_n3626_n1764# sky130_fd_pr__pfet_01v8 ad=1.5522 pd=8.74 as=0 ps=0 w=3.98 l=2.99
X11 VTAIL.t4 VN.t4 VDD2.t0 w_n3626_n1764# sky130_fd_pr__pfet_01v8 ad=0.6567 pd=4.31 as=0.6567 ps=4.31 w=3.98 l=2.99
X12 VDD1.t2 VP.t3 VTAIL.t2 w_n3626_n1764# sky130_fd_pr__pfet_01v8 ad=1.5522 pd=8.74 as=0.6567 ps=4.31 w=3.98 l=2.99
X13 VTAIL.t1 VP.t4 VDD1.t1 w_n3626_n1764# sky130_fd_pr__pfet_01v8 ad=0.6567 pd=4.31 as=0.6567 ps=4.31 w=3.98 l=2.99
X14 VDD2.t2 VN.t5 VTAIL.t3 w_n3626_n1764# sky130_fd_pr__pfet_01v8 ad=1.5522 pd=8.74 as=0.6567 ps=4.31 w=3.98 l=2.99
X15 VDD1.t0 VP.t5 VTAIL.t0 w_n3626_n1764# sky130_fd_pr__pfet_01v8 ad=0.6567 pd=4.31 as=1.5522 ps=8.74 w=3.98 l=2.99
R0 B.n434 B.n53 585
R1 B.n436 B.n435 585
R2 B.n437 B.n52 585
R3 B.n439 B.n438 585
R4 B.n440 B.n51 585
R5 B.n442 B.n441 585
R6 B.n443 B.n50 585
R7 B.n445 B.n444 585
R8 B.n446 B.n49 585
R9 B.n448 B.n447 585
R10 B.n449 B.n48 585
R11 B.n451 B.n450 585
R12 B.n452 B.n47 585
R13 B.n454 B.n453 585
R14 B.n455 B.n46 585
R15 B.n457 B.n456 585
R16 B.n458 B.n45 585
R17 B.n460 B.n459 585
R18 B.n462 B.n42 585
R19 B.n464 B.n463 585
R20 B.n465 B.n41 585
R21 B.n467 B.n466 585
R22 B.n468 B.n40 585
R23 B.n470 B.n469 585
R24 B.n471 B.n39 585
R25 B.n473 B.n472 585
R26 B.n474 B.n35 585
R27 B.n476 B.n475 585
R28 B.n477 B.n34 585
R29 B.n479 B.n478 585
R30 B.n480 B.n33 585
R31 B.n482 B.n481 585
R32 B.n483 B.n32 585
R33 B.n485 B.n484 585
R34 B.n486 B.n31 585
R35 B.n488 B.n487 585
R36 B.n489 B.n30 585
R37 B.n491 B.n490 585
R38 B.n492 B.n29 585
R39 B.n494 B.n493 585
R40 B.n495 B.n28 585
R41 B.n497 B.n496 585
R42 B.n498 B.n27 585
R43 B.n500 B.n499 585
R44 B.n501 B.n26 585
R45 B.n503 B.n502 585
R46 B.n433 B.n432 585
R47 B.n431 B.n54 585
R48 B.n430 B.n429 585
R49 B.n428 B.n55 585
R50 B.n427 B.n426 585
R51 B.n425 B.n56 585
R52 B.n424 B.n423 585
R53 B.n422 B.n57 585
R54 B.n421 B.n420 585
R55 B.n419 B.n58 585
R56 B.n418 B.n417 585
R57 B.n416 B.n59 585
R58 B.n415 B.n414 585
R59 B.n413 B.n60 585
R60 B.n412 B.n411 585
R61 B.n410 B.n61 585
R62 B.n409 B.n408 585
R63 B.n407 B.n62 585
R64 B.n406 B.n405 585
R65 B.n404 B.n63 585
R66 B.n403 B.n402 585
R67 B.n401 B.n64 585
R68 B.n400 B.n399 585
R69 B.n398 B.n65 585
R70 B.n397 B.n396 585
R71 B.n395 B.n66 585
R72 B.n394 B.n393 585
R73 B.n392 B.n67 585
R74 B.n391 B.n390 585
R75 B.n389 B.n68 585
R76 B.n388 B.n387 585
R77 B.n386 B.n69 585
R78 B.n385 B.n384 585
R79 B.n383 B.n70 585
R80 B.n382 B.n381 585
R81 B.n380 B.n71 585
R82 B.n379 B.n378 585
R83 B.n377 B.n72 585
R84 B.n376 B.n375 585
R85 B.n374 B.n73 585
R86 B.n373 B.n372 585
R87 B.n371 B.n74 585
R88 B.n370 B.n369 585
R89 B.n368 B.n75 585
R90 B.n367 B.n366 585
R91 B.n365 B.n76 585
R92 B.n364 B.n363 585
R93 B.n362 B.n77 585
R94 B.n361 B.n360 585
R95 B.n359 B.n78 585
R96 B.n358 B.n357 585
R97 B.n356 B.n79 585
R98 B.n355 B.n354 585
R99 B.n353 B.n80 585
R100 B.n352 B.n351 585
R101 B.n350 B.n81 585
R102 B.n349 B.n348 585
R103 B.n347 B.n82 585
R104 B.n346 B.n345 585
R105 B.n344 B.n83 585
R106 B.n343 B.n342 585
R107 B.n341 B.n84 585
R108 B.n340 B.n339 585
R109 B.n338 B.n85 585
R110 B.n337 B.n336 585
R111 B.n335 B.n86 585
R112 B.n334 B.n333 585
R113 B.n332 B.n87 585
R114 B.n331 B.n330 585
R115 B.n329 B.n88 585
R116 B.n328 B.n327 585
R117 B.n326 B.n89 585
R118 B.n325 B.n324 585
R119 B.n323 B.n90 585
R120 B.n322 B.n321 585
R121 B.n320 B.n91 585
R122 B.n319 B.n318 585
R123 B.n317 B.n92 585
R124 B.n316 B.n315 585
R125 B.n314 B.n93 585
R126 B.n313 B.n312 585
R127 B.n311 B.n94 585
R128 B.n310 B.n309 585
R129 B.n308 B.n95 585
R130 B.n307 B.n306 585
R131 B.n305 B.n96 585
R132 B.n304 B.n303 585
R133 B.n302 B.n97 585
R134 B.n301 B.n300 585
R135 B.n299 B.n98 585
R136 B.n298 B.n297 585
R137 B.n296 B.n99 585
R138 B.n295 B.n294 585
R139 B.n293 B.n100 585
R140 B.n292 B.n291 585
R141 B.n221 B.n128 585
R142 B.n223 B.n222 585
R143 B.n224 B.n127 585
R144 B.n226 B.n225 585
R145 B.n227 B.n126 585
R146 B.n229 B.n228 585
R147 B.n230 B.n125 585
R148 B.n232 B.n231 585
R149 B.n233 B.n124 585
R150 B.n235 B.n234 585
R151 B.n236 B.n123 585
R152 B.n238 B.n237 585
R153 B.n239 B.n122 585
R154 B.n241 B.n240 585
R155 B.n242 B.n121 585
R156 B.n244 B.n243 585
R157 B.n245 B.n120 585
R158 B.n247 B.n246 585
R159 B.n249 B.n248 585
R160 B.n250 B.n116 585
R161 B.n252 B.n251 585
R162 B.n253 B.n115 585
R163 B.n255 B.n254 585
R164 B.n256 B.n114 585
R165 B.n258 B.n257 585
R166 B.n259 B.n113 585
R167 B.n261 B.n260 585
R168 B.n262 B.n110 585
R169 B.n265 B.n264 585
R170 B.n266 B.n109 585
R171 B.n268 B.n267 585
R172 B.n269 B.n108 585
R173 B.n271 B.n270 585
R174 B.n272 B.n107 585
R175 B.n274 B.n273 585
R176 B.n275 B.n106 585
R177 B.n277 B.n276 585
R178 B.n278 B.n105 585
R179 B.n280 B.n279 585
R180 B.n281 B.n104 585
R181 B.n283 B.n282 585
R182 B.n284 B.n103 585
R183 B.n286 B.n285 585
R184 B.n287 B.n102 585
R185 B.n289 B.n288 585
R186 B.n290 B.n101 585
R187 B.n220 B.n219 585
R188 B.n218 B.n129 585
R189 B.n217 B.n216 585
R190 B.n215 B.n130 585
R191 B.n214 B.n213 585
R192 B.n212 B.n131 585
R193 B.n211 B.n210 585
R194 B.n209 B.n132 585
R195 B.n208 B.n207 585
R196 B.n206 B.n133 585
R197 B.n205 B.n204 585
R198 B.n203 B.n134 585
R199 B.n202 B.n201 585
R200 B.n200 B.n135 585
R201 B.n199 B.n198 585
R202 B.n197 B.n136 585
R203 B.n196 B.n195 585
R204 B.n194 B.n137 585
R205 B.n193 B.n192 585
R206 B.n191 B.n138 585
R207 B.n190 B.n189 585
R208 B.n188 B.n139 585
R209 B.n187 B.n186 585
R210 B.n185 B.n140 585
R211 B.n184 B.n183 585
R212 B.n182 B.n141 585
R213 B.n181 B.n180 585
R214 B.n179 B.n142 585
R215 B.n178 B.n177 585
R216 B.n176 B.n143 585
R217 B.n175 B.n174 585
R218 B.n173 B.n144 585
R219 B.n172 B.n171 585
R220 B.n170 B.n145 585
R221 B.n169 B.n168 585
R222 B.n167 B.n146 585
R223 B.n166 B.n165 585
R224 B.n164 B.n147 585
R225 B.n163 B.n162 585
R226 B.n161 B.n148 585
R227 B.n160 B.n159 585
R228 B.n158 B.n149 585
R229 B.n157 B.n156 585
R230 B.n155 B.n150 585
R231 B.n154 B.n153 585
R232 B.n152 B.n151 585
R233 B.n2 B.n0 585
R234 B.n573 B.n1 585
R235 B.n572 B.n571 585
R236 B.n570 B.n3 585
R237 B.n569 B.n568 585
R238 B.n567 B.n4 585
R239 B.n566 B.n565 585
R240 B.n564 B.n5 585
R241 B.n563 B.n562 585
R242 B.n561 B.n6 585
R243 B.n560 B.n559 585
R244 B.n558 B.n7 585
R245 B.n557 B.n556 585
R246 B.n555 B.n8 585
R247 B.n554 B.n553 585
R248 B.n552 B.n9 585
R249 B.n551 B.n550 585
R250 B.n549 B.n10 585
R251 B.n548 B.n547 585
R252 B.n546 B.n11 585
R253 B.n545 B.n544 585
R254 B.n543 B.n12 585
R255 B.n542 B.n541 585
R256 B.n540 B.n13 585
R257 B.n539 B.n538 585
R258 B.n537 B.n14 585
R259 B.n536 B.n535 585
R260 B.n534 B.n15 585
R261 B.n533 B.n532 585
R262 B.n531 B.n16 585
R263 B.n530 B.n529 585
R264 B.n528 B.n17 585
R265 B.n527 B.n526 585
R266 B.n525 B.n18 585
R267 B.n524 B.n523 585
R268 B.n522 B.n19 585
R269 B.n521 B.n520 585
R270 B.n519 B.n20 585
R271 B.n518 B.n517 585
R272 B.n516 B.n21 585
R273 B.n515 B.n514 585
R274 B.n513 B.n22 585
R275 B.n512 B.n511 585
R276 B.n510 B.n23 585
R277 B.n509 B.n508 585
R278 B.n507 B.n24 585
R279 B.n506 B.n505 585
R280 B.n504 B.n25 585
R281 B.n575 B.n574 585
R282 B.n219 B.n128 497.305
R283 B.n502 B.n25 497.305
R284 B.n291 B.n290 497.305
R285 B.n434 B.n433 497.305
R286 B.n111 B.t2 299.63
R287 B.n43 B.t4 299.63
R288 B.n117 B.t8 299.63
R289 B.n36 B.t10 299.63
R290 B.n111 B.t0 240.649
R291 B.n117 B.t6 240.649
R292 B.n36 B.t9 240.649
R293 B.n43 B.t3 240.649
R294 B.n112 B.t1 235.242
R295 B.n44 B.t5 235.242
R296 B.n118 B.t7 235.242
R297 B.n37 B.t11 235.242
R298 B.n219 B.n218 163.367
R299 B.n218 B.n217 163.367
R300 B.n217 B.n130 163.367
R301 B.n213 B.n130 163.367
R302 B.n213 B.n212 163.367
R303 B.n212 B.n211 163.367
R304 B.n211 B.n132 163.367
R305 B.n207 B.n132 163.367
R306 B.n207 B.n206 163.367
R307 B.n206 B.n205 163.367
R308 B.n205 B.n134 163.367
R309 B.n201 B.n134 163.367
R310 B.n201 B.n200 163.367
R311 B.n200 B.n199 163.367
R312 B.n199 B.n136 163.367
R313 B.n195 B.n136 163.367
R314 B.n195 B.n194 163.367
R315 B.n194 B.n193 163.367
R316 B.n193 B.n138 163.367
R317 B.n189 B.n138 163.367
R318 B.n189 B.n188 163.367
R319 B.n188 B.n187 163.367
R320 B.n187 B.n140 163.367
R321 B.n183 B.n140 163.367
R322 B.n183 B.n182 163.367
R323 B.n182 B.n181 163.367
R324 B.n181 B.n142 163.367
R325 B.n177 B.n142 163.367
R326 B.n177 B.n176 163.367
R327 B.n176 B.n175 163.367
R328 B.n175 B.n144 163.367
R329 B.n171 B.n144 163.367
R330 B.n171 B.n170 163.367
R331 B.n170 B.n169 163.367
R332 B.n169 B.n146 163.367
R333 B.n165 B.n146 163.367
R334 B.n165 B.n164 163.367
R335 B.n164 B.n163 163.367
R336 B.n163 B.n148 163.367
R337 B.n159 B.n148 163.367
R338 B.n159 B.n158 163.367
R339 B.n158 B.n157 163.367
R340 B.n157 B.n150 163.367
R341 B.n153 B.n150 163.367
R342 B.n153 B.n152 163.367
R343 B.n152 B.n2 163.367
R344 B.n574 B.n2 163.367
R345 B.n574 B.n573 163.367
R346 B.n573 B.n572 163.367
R347 B.n572 B.n3 163.367
R348 B.n568 B.n3 163.367
R349 B.n568 B.n567 163.367
R350 B.n567 B.n566 163.367
R351 B.n566 B.n5 163.367
R352 B.n562 B.n5 163.367
R353 B.n562 B.n561 163.367
R354 B.n561 B.n560 163.367
R355 B.n560 B.n7 163.367
R356 B.n556 B.n7 163.367
R357 B.n556 B.n555 163.367
R358 B.n555 B.n554 163.367
R359 B.n554 B.n9 163.367
R360 B.n550 B.n9 163.367
R361 B.n550 B.n549 163.367
R362 B.n549 B.n548 163.367
R363 B.n548 B.n11 163.367
R364 B.n544 B.n11 163.367
R365 B.n544 B.n543 163.367
R366 B.n543 B.n542 163.367
R367 B.n542 B.n13 163.367
R368 B.n538 B.n13 163.367
R369 B.n538 B.n537 163.367
R370 B.n537 B.n536 163.367
R371 B.n536 B.n15 163.367
R372 B.n532 B.n15 163.367
R373 B.n532 B.n531 163.367
R374 B.n531 B.n530 163.367
R375 B.n530 B.n17 163.367
R376 B.n526 B.n17 163.367
R377 B.n526 B.n525 163.367
R378 B.n525 B.n524 163.367
R379 B.n524 B.n19 163.367
R380 B.n520 B.n19 163.367
R381 B.n520 B.n519 163.367
R382 B.n519 B.n518 163.367
R383 B.n518 B.n21 163.367
R384 B.n514 B.n21 163.367
R385 B.n514 B.n513 163.367
R386 B.n513 B.n512 163.367
R387 B.n512 B.n23 163.367
R388 B.n508 B.n23 163.367
R389 B.n508 B.n507 163.367
R390 B.n507 B.n506 163.367
R391 B.n506 B.n25 163.367
R392 B.n223 B.n128 163.367
R393 B.n224 B.n223 163.367
R394 B.n225 B.n224 163.367
R395 B.n225 B.n126 163.367
R396 B.n229 B.n126 163.367
R397 B.n230 B.n229 163.367
R398 B.n231 B.n230 163.367
R399 B.n231 B.n124 163.367
R400 B.n235 B.n124 163.367
R401 B.n236 B.n235 163.367
R402 B.n237 B.n236 163.367
R403 B.n237 B.n122 163.367
R404 B.n241 B.n122 163.367
R405 B.n242 B.n241 163.367
R406 B.n243 B.n242 163.367
R407 B.n243 B.n120 163.367
R408 B.n247 B.n120 163.367
R409 B.n248 B.n247 163.367
R410 B.n248 B.n116 163.367
R411 B.n252 B.n116 163.367
R412 B.n253 B.n252 163.367
R413 B.n254 B.n253 163.367
R414 B.n254 B.n114 163.367
R415 B.n258 B.n114 163.367
R416 B.n259 B.n258 163.367
R417 B.n260 B.n259 163.367
R418 B.n260 B.n110 163.367
R419 B.n265 B.n110 163.367
R420 B.n266 B.n265 163.367
R421 B.n267 B.n266 163.367
R422 B.n267 B.n108 163.367
R423 B.n271 B.n108 163.367
R424 B.n272 B.n271 163.367
R425 B.n273 B.n272 163.367
R426 B.n273 B.n106 163.367
R427 B.n277 B.n106 163.367
R428 B.n278 B.n277 163.367
R429 B.n279 B.n278 163.367
R430 B.n279 B.n104 163.367
R431 B.n283 B.n104 163.367
R432 B.n284 B.n283 163.367
R433 B.n285 B.n284 163.367
R434 B.n285 B.n102 163.367
R435 B.n289 B.n102 163.367
R436 B.n290 B.n289 163.367
R437 B.n291 B.n100 163.367
R438 B.n295 B.n100 163.367
R439 B.n296 B.n295 163.367
R440 B.n297 B.n296 163.367
R441 B.n297 B.n98 163.367
R442 B.n301 B.n98 163.367
R443 B.n302 B.n301 163.367
R444 B.n303 B.n302 163.367
R445 B.n303 B.n96 163.367
R446 B.n307 B.n96 163.367
R447 B.n308 B.n307 163.367
R448 B.n309 B.n308 163.367
R449 B.n309 B.n94 163.367
R450 B.n313 B.n94 163.367
R451 B.n314 B.n313 163.367
R452 B.n315 B.n314 163.367
R453 B.n315 B.n92 163.367
R454 B.n319 B.n92 163.367
R455 B.n320 B.n319 163.367
R456 B.n321 B.n320 163.367
R457 B.n321 B.n90 163.367
R458 B.n325 B.n90 163.367
R459 B.n326 B.n325 163.367
R460 B.n327 B.n326 163.367
R461 B.n327 B.n88 163.367
R462 B.n331 B.n88 163.367
R463 B.n332 B.n331 163.367
R464 B.n333 B.n332 163.367
R465 B.n333 B.n86 163.367
R466 B.n337 B.n86 163.367
R467 B.n338 B.n337 163.367
R468 B.n339 B.n338 163.367
R469 B.n339 B.n84 163.367
R470 B.n343 B.n84 163.367
R471 B.n344 B.n343 163.367
R472 B.n345 B.n344 163.367
R473 B.n345 B.n82 163.367
R474 B.n349 B.n82 163.367
R475 B.n350 B.n349 163.367
R476 B.n351 B.n350 163.367
R477 B.n351 B.n80 163.367
R478 B.n355 B.n80 163.367
R479 B.n356 B.n355 163.367
R480 B.n357 B.n356 163.367
R481 B.n357 B.n78 163.367
R482 B.n361 B.n78 163.367
R483 B.n362 B.n361 163.367
R484 B.n363 B.n362 163.367
R485 B.n363 B.n76 163.367
R486 B.n367 B.n76 163.367
R487 B.n368 B.n367 163.367
R488 B.n369 B.n368 163.367
R489 B.n369 B.n74 163.367
R490 B.n373 B.n74 163.367
R491 B.n374 B.n373 163.367
R492 B.n375 B.n374 163.367
R493 B.n375 B.n72 163.367
R494 B.n379 B.n72 163.367
R495 B.n380 B.n379 163.367
R496 B.n381 B.n380 163.367
R497 B.n381 B.n70 163.367
R498 B.n385 B.n70 163.367
R499 B.n386 B.n385 163.367
R500 B.n387 B.n386 163.367
R501 B.n387 B.n68 163.367
R502 B.n391 B.n68 163.367
R503 B.n392 B.n391 163.367
R504 B.n393 B.n392 163.367
R505 B.n393 B.n66 163.367
R506 B.n397 B.n66 163.367
R507 B.n398 B.n397 163.367
R508 B.n399 B.n398 163.367
R509 B.n399 B.n64 163.367
R510 B.n403 B.n64 163.367
R511 B.n404 B.n403 163.367
R512 B.n405 B.n404 163.367
R513 B.n405 B.n62 163.367
R514 B.n409 B.n62 163.367
R515 B.n410 B.n409 163.367
R516 B.n411 B.n410 163.367
R517 B.n411 B.n60 163.367
R518 B.n415 B.n60 163.367
R519 B.n416 B.n415 163.367
R520 B.n417 B.n416 163.367
R521 B.n417 B.n58 163.367
R522 B.n421 B.n58 163.367
R523 B.n422 B.n421 163.367
R524 B.n423 B.n422 163.367
R525 B.n423 B.n56 163.367
R526 B.n427 B.n56 163.367
R527 B.n428 B.n427 163.367
R528 B.n429 B.n428 163.367
R529 B.n429 B.n54 163.367
R530 B.n433 B.n54 163.367
R531 B.n502 B.n501 163.367
R532 B.n501 B.n500 163.367
R533 B.n500 B.n27 163.367
R534 B.n496 B.n27 163.367
R535 B.n496 B.n495 163.367
R536 B.n495 B.n494 163.367
R537 B.n494 B.n29 163.367
R538 B.n490 B.n29 163.367
R539 B.n490 B.n489 163.367
R540 B.n489 B.n488 163.367
R541 B.n488 B.n31 163.367
R542 B.n484 B.n31 163.367
R543 B.n484 B.n483 163.367
R544 B.n483 B.n482 163.367
R545 B.n482 B.n33 163.367
R546 B.n478 B.n33 163.367
R547 B.n478 B.n477 163.367
R548 B.n477 B.n476 163.367
R549 B.n476 B.n35 163.367
R550 B.n472 B.n35 163.367
R551 B.n472 B.n471 163.367
R552 B.n471 B.n470 163.367
R553 B.n470 B.n40 163.367
R554 B.n466 B.n40 163.367
R555 B.n466 B.n465 163.367
R556 B.n465 B.n464 163.367
R557 B.n464 B.n42 163.367
R558 B.n459 B.n42 163.367
R559 B.n459 B.n458 163.367
R560 B.n458 B.n457 163.367
R561 B.n457 B.n46 163.367
R562 B.n453 B.n46 163.367
R563 B.n453 B.n452 163.367
R564 B.n452 B.n451 163.367
R565 B.n451 B.n48 163.367
R566 B.n447 B.n48 163.367
R567 B.n447 B.n446 163.367
R568 B.n446 B.n445 163.367
R569 B.n445 B.n50 163.367
R570 B.n441 B.n50 163.367
R571 B.n441 B.n440 163.367
R572 B.n440 B.n439 163.367
R573 B.n439 B.n52 163.367
R574 B.n435 B.n52 163.367
R575 B.n435 B.n434 163.367
R576 B.n112 B.n111 64.3884
R577 B.n118 B.n117 64.3884
R578 B.n37 B.n36 64.3884
R579 B.n44 B.n43 64.3884
R580 B.n263 B.n112 59.5399
R581 B.n119 B.n118 59.5399
R582 B.n38 B.n37 59.5399
R583 B.n461 B.n44 59.5399
R584 B.n504 B.n503 32.3127
R585 B.n432 B.n53 32.3127
R586 B.n292 B.n101 32.3127
R587 B.n221 B.n220 32.3127
R588 B B.n575 18.0485
R589 B.n503 B.n26 10.6151
R590 B.n499 B.n26 10.6151
R591 B.n499 B.n498 10.6151
R592 B.n498 B.n497 10.6151
R593 B.n497 B.n28 10.6151
R594 B.n493 B.n28 10.6151
R595 B.n493 B.n492 10.6151
R596 B.n492 B.n491 10.6151
R597 B.n491 B.n30 10.6151
R598 B.n487 B.n30 10.6151
R599 B.n487 B.n486 10.6151
R600 B.n486 B.n485 10.6151
R601 B.n485 B.n32 10.6151
R602 B.n481 B.n32 10.6151
R603 B.n481 B.n480 10.6151
R604 B.n480 B.n479 10.6151
R605 B.n479 B.n34 10.6151
R606 B.n475 B.n474 10.6151
R607 B.n474 B.n473 10.6151
R608 B.n473 B.n39 10.6151
R609 B.n469 B.n39 10.6151
R610 B.n469 B.n468 10.6151
R611 B.n468 B.n467 10.6151
R612 B.n467 B.n41 10.6151
R613 B.n463 B.n41 10.6151
R614 B.n463 B.n462 10.6151
R615 B.n460 B.n45 10.6151
R616 B.n456 B.n45 10.6151
R617 B.n456 B.n455 10.6151
R618 B.n455 B.n454 10.6151
R619 B.n454 B.n47 10.6151
R620 B.n450 B.n47 10.6151
R621 B.n450 B.n449 10.6151
R622 B.n449 B.n448 10.6151
R623 B.n448 B.n49 10.6151
R624 B.n444 B.n49 10.6151
R625 B.n444 B.n443 10.6151
R626 B.n443 B.n442 10.6151
R627 B.n442 B.n51 10.6151
R628 B.n438 B.n51 10.6151
R629 B.n438 B.n437 10.6151
R630 B.n437 B.n436 10.6151
R631 B.n436 B.n53 10.6151
R632 B.n293 B.n292 10.6151
R633 B.n294 B.n293 10.6151
R634 B.n294 B.n99 10.6151
R635 B.n298 B.n99 10.6151
R636 B.n299 B.n298 10.6151
R637 B.n300 B.n299 10.6151
R638 B.n300 B.n97 10.6151
R639 B.n304 B.n97 10.6151
R640 B.n305 B.n304 10.6151
R641 B.n306 B.n305 10.6151
R642 B.n306 B.n95 10.6151
R643 B.n310 B.n95 10.6151
R644 B.n311 B.n310 10.6151
R645 B.n312 B.n311 10.6151
R646 B.n312 B.n93 10.6151
R647 B.n316 B.n93 10.6151
R648 B.n317 B.n316 10.6151
R649 B.n318 B.n317 10.6151
R650 B.n318 B.n91 10.6151
R651 B.n322 B.n91 10.6151
R652 B.n323 B.n322 10.6151
R653 B.n324 B.n323 10.6151
R654 B.n324 B.n89 10.6151
R655 B.n328 B.n89 10.6151
R656 B.n329 B.n328 10.6151
R657 B.n330 B.n329 10.6151
R658 B.n330 B.n87 10.6151
R659 B.n334 B.n87 10.6151
R660 B.n335 B.n334 10.6151
R661 B.n336 B.n335 10.6151
R662 B.n336 B.n85 10.6151
R663 B.n340 B.n85 10.6151
R664 B.n341 B.n340 10.6151
R665 B.n342 B.n341 10.6151
R666 B.n342 B.n83 10.6151
R667 B.n346 B.n83 10.6151
R668 B.n347 B.n346 10.6151
R669 B.n348 B.n347 10.6151
R670 B.n348 B.n81 10.6151
R671 B.n352 B.n81 10.6151
R672 B.n353 B.n352 10.6151
R673 B.n354 B.n353 10.6151
R674 B.n354 B.n79 10.6151
R675 B.n358 B.n79 10.6151
R676 B.n359 B.n358 10.6151
R677 B.n360 B.n359 10.6151
R678 B.n360 B.n77 10.6151
R679 B.n364 B.n77 10.6151
R680 B.n365 B.n364 10.6151
R681 B.n366 B.n365 10.6151
R682 B.n366 B.n75 10.6151
R683 B.n370 B.n75 10.6151
R684 B.n371 B.n370 10.6151
R685 B.n372 B.n371 10.6151
R686 B.n372 B.n73 10.6151
R687 B.n376 B.n73 10.6151
R688 B.n377 B.n376 10.6151
R689 B.n378 B.n377 10.6151
R690 B.n378 B.n71 10.6151
R691 B.n382 B.n71 10.6151
R692 B.n383 B.n382 10.6151
R693 B.n384 B.n383 10.6151
R694 B.n384 B.n69 10.6151
R695 B.n388 B.n69 10.6151
R696 B.n389 B.n388 10.6151
R697 B.n390 B.n389 10.6151
R698 B.n390 B.n67 10.6151
R699 B.n394 B.n67 10.6151
R700 B.n395 B.n394 10.6151
R701 B.n396 B.n395 10.6151
R702 B.n396 B.n65 10.6151
R703 B.n400 B.n65 10.6151
R704 B.n401 B.n400 10.6151
R705 B.n402 B.n401 10.6151
R706 B.n402 B.n63 10.6151
R707 B.n406 B.n63 10.6151
R708 B.n407 B.n406 10.6151
R709 B.n408 B.n407 10.6151
R710 B.n408 B.n61 10.6151
R711 B.n412 B.n61 10.6151
R712 B.n413 B.n412 10.6151
R713 B.n414 B.n413 10.6151
R714 B.n414 B.n59 10.6151
R715 B.n418 B.n59 10.6151
R716 B.n419 B.n418 10.6151
R717 B.n420 B.n419 10.6151
R718 B.n420 B.n57 10.6151
R719 B.n424 B.n57 10.6151
R720 B.n425 B.n424 10.6151
R721 B.n426 B.n425 10.6151
R722 B.n426 B.n55 10.6151
R723 B.n430 B.n55 10.6151
R724 B.n431 B.n430 10.6151
R725 B.n432 B.n431 10.6151
R726 B.n222 B.n221 10.6151
R727 B.n222 B.n127 10.6151
R728 B.n226 B.n127 10.6151
R729 B.n227 B.n226 10.6151
R730 B.n228 B.n227 10.6151
R731 B.n228 B.n125 10.6151
R732 B.n232 B.n125 10.6151
R733 B.n233 B.n232 10.6151
R734 B.n234 B.n233 10.6151
R735 B.n234 B.n123 10.6151
R736 B.n238 B.n123 10.6151
R737 B.n239 B.n238 10.6151
R738 B.n240 B.n239 10.6151
R739 B.n240 B.n121 10.6151
R740 B.n244 B.n121 10.6151
R741 B.n245 B.n244 10.6151
R742 B.n246 B.n245 10.6151
R743 B.n250 B.n249 10.6151
R744 B.n251 B.n250 10.6151
R745 B.n251 B.n115 10.6151
R746 B.n255 B.n115 10.6151
R747 B.n256 B.n255 10.6151
R748 B.n257 B.n256 10.6151
R749 B.n257 B.n113 10.6151
R750 B.n261 B.n113 10.6151
R751 B.n262 B.n261 10.6151
R752 B.n264 B.n109 10.6151
R753 B.n268 B.n109 10.6151
R754 B.n269 B.n268 10.6151
R755 B.n270 B.n269 10.6151
R756 B.n270 B.n107 10.6151
R757 B.n274 B.n107 10.6151
R758 B.n275 B.n274 10.6151
R759 B.n276 B.n275 10.6151
R760 B.n276 B.n105 10.6151
R761 B.n280 B.n105 10.6151
R762 B.n281 B.n280 10.6151
R763 B.n282 B.n281 10.6151
R764 B.n282 B.n103 10.6151
R765 B.n286 B.n103 10.6151
R766 B.n287 B.n286 10.6151
R767 B.n288 B.n287 10.6151
R768 B.n288 B.n101 10.6151
R769 B.n220 B.n129 10.6151
R770 B.n216 B.n129 10.6151
R771 B.n216 B.n215 10.6151
R772 B.n215 B.n214 10.6151
R773 B.n214 B.n131 10.6151
R774 B.n210 B.n131 10.6151
R775 B.n210 B.n209 10.6151
R776 B.n209 B.n208 10.6151
R777 B.n208 B.n133 10.6151
R778 B.n204 B.n133 10.6151
R779 B.n204 B.n203 10.6151
R780 B.n203 B.n202 10.6151
R781 B.n202 B.n135 10.6151
R782 B.n198 B.n135 10.6151
R783 B.n198 B.n197 10.6151
R784 B.n197 B.n196 10.6151
R785 B.n196 B.n137 10.6151
R786 B.n192 B.n137 10.6151
R787 B.n192 B.n191 10.6151
R788 B.n191 B.n190 10.6151
R789 B.n190 B.n139 10.6151
R790 B.n186 B.n139 10.6151
R791 B.n186 B.n185 10.6151
R792 B.n185 B.n184 10.6151
R793 B.n184 B.n141 10.6151
R794 B.n180 B.n141 10.6151
R795 B.n180 B.n179 10.6151
R796 B.n179 B.n178 10.6151
R797 B.n178 B.n143 10.6151
R798 B.n174 B.n143 10.6151
R799 B.n174 B.n173 10.6151
R800 B.n173 B.n172 10.6151
R801 B.n172 B.n145 10.6151
R802 B.n168 B.n145 10.6151
R803 B.n168 B.n167 10.6151
R804 B.n167 B.n166 10.6151
R805 B.n166 B.n147 10.6151
R806 B.n162 B.n147 10.6151
R807 B.n162 B.n161 10.6151
R808 B.n161 B.n160 10.6151
R809 B.n160 B.n149 10.6151
R810 B.n156 B.n149 10.6151
R811 B.n156 B.n155 10.6151
R812 B.n155 B.n154 10.6151
R813 B.n154 B.n151 10.6151
R814 B.n151 B.n0 10.6151
R815 B.n571 B.n1 10.6151
R816 B.n571 B.n570 10.6151
R817 B.n570 B.n569 10.6151
R818 B.n569 B.n4 10.6151
R819 B.n565 B.n4 10.6151
R820 B.n565 B.n564 10.6151
R821 B.n564 B.n563 10.6151
R822 B.n563 B.n6 10.6151
R823 B.n559 B.n6 10.6151
R824 B.n559 B.n558 10.6151
R825 B.n558 B.n557 10.6151
R826 B.n557 B.n8 10.6151
R827 B.n553 B.n8 10.6151
R828 B.n553 B.n552 10.6151
R829 B.n552 B.n551 10.6151
R830 B.n551 B.n10 10.6151
R831 B.n547 B.n10 10.6151
R832 B.n547 B.n546 10.6151
R833 B.n546 B.n545 10.6151
R834 B.n545 B.n12 10.6151
R835 B.n541 B.n12 10.6151
R836 B.n541 B.n540 10.6151
R837 B.n540 B.n539 10.6151
R838 B.n539 B.n14 10.6151
R839 B.n535 B.n14 10.6151
R840 B.n535 B.n534 10.6151
R841 B.n534 B.n533 10.6151
R842 B.n533 B.n16 10.6151
R843 B.n529 B.n16 10.6151
R844 B.n529 B.n528 10.6151
R845 B.n528 B.n527 10.6151
R846 B.n527 B.n18 10.6151
R847 B.n523 B.n18 10.6151
R848 B.n523 B.n522 10.6151
R849 B.n522 B.n521 10.6151
R850 B.n521 B.n20 10.6151
R851 B.n517 B.n20 10.6151
R852 B.n517 B.n516 10.6151
R853 B.n516 B.n515 10.6151
R854 B.n515 B.n22 10.6151
R855 B.n511 B.n22 10.6151
R856 B.n511 B.n510 10.6151
R857 B.n510 B.n509 10.6151
R858 B.n509 B.n24 10.6151
R859 B.n505 B.n24 10.6151
R860 B.n505 B.n504 10.6151
R861 B.n38 B.n34 9.36635
R862 B.n461 B.n460 9.36635
R863 B.n246 B.n119 9.36635
R864 B.n264 B.n263 9.36635
R865 B.n575 B.n0 2.81026
R866 B.n575 B.n1 2.81026
R867 B.n475 B.n38 1.24928
R868 B.n462 B.n461 1.24928
R869 B.n249 B.n119 1.24928
R870 B.n263 B.n262 1.24928
R871 VN.n30 VN.n29 161.3
R872 VN.n28 VN.n17 161.3
R873 VN.n27 VN.n26 161.3
R874 VN.n25 VN.n18 161.3
R875 VN.n24 VN.n23 161.3
R876 VN.n22 VN.n19 161.3
R877 VN.n14 VN.n13 161.3
R878 VN.n12 VN.n1 161.3
R879 VN.n11 VN.n10 161.3
R880 VN.n9 VN.n2 161.3
R881 VN.n8 VN.n7 161.3
R882 VN.n6 VN.n3 161.3
R883 VN.n15 VN.n0 74.5068
R884 VN.n31 VN.n16 74.5068
R885 VN.n20 VN.t2 65.3335
R886 VN.n4 VN.t5 65.3335
R887 VN.n11 VN.n2 56.0773
R888 VN.n27 VN.n18 56.0773
R889 VN.n5 VN.n4 49.3258
R890 VN.n21 VN.n20 49.3258
R891 VN VN.n31 44.3466
R892 VN.n5 VN.t4 32.0801
R893 VN.n0 VN.t1 32.0801
R894 VN.n21 VN.t0 32.0801
R895 VN.n16 VN.t3 32.0801
R896 VN.n7 VN.n2 25.0767
R897 VN.n23 VN.n18 25.0767
R898 VN.n6 VN.n5 24.5923
R899 VN.n7 VN.n6 24.5923
R900 VN.n12 VN.n11 24.5923
R901 VN.n13 VN.n12 24.5923
R902 VN.n23 VN.n22 24.5923
R903 VN.n22 VN.n21 24.5923
R904 VN.n29 VN.n28 24.5923
R905 VN.n28 VN.n27 24.5923
R906 VN.n13 VN.n0 15.7393
R907 VN.n29 VN.n16 15.7393
R908 VN.n4 VN.n3 4.10787
R909 VN.n20 VN.n19 4.10787
R910 VN.n31 VN.n30 0.354861
R911 VN.n15 VN.n14 0.354861
R912 VN VN.n15 0.267071
R913 VN.n30 VN.n17 0.189894
R914 VN.n26 VN.n17 0.189894
R915 VN.n26 VN.n25 0.189894
R916 VN.n25 VN.n24 0.189894
R917 VN.n24 VN.n19 0.189894
R918 VN.n8 VN.n3 0.189894
R919 VN.n9 VN.n8 0.189894
R920 VN.n10 VN.n9 0.189894
R921 VN.n10 VN.n1 0.189894
R922 VN.n14 VN.n1 0.189894
R923 VDD2.n35 VDD2.n21 756.745
R924 VDD2.n14 VDD2.n0 756.745
R925 VDD2.n36 VDD2.n35 585
R926 VDD2.n34 VDD2.n33 585
R927 VDD2.n25 VDD2.n24 585
R928 VDD2.n28 VDD2.n27 585
R929 VDD2.n7 VDD2.n6 585
R930 VDD2.n4 VDD2.n3 585
R931 VDD2.n13 VDD2.n12 585
R932 VDD2.n15 VDD2.n14 585
R933 VDD2.t5 VDD2.n26 330.707
R934 VDD2.t2 VDD2.n5 330.707
R935 VDD2.n35 VDD2.n34 171.744
R936 VDD2.n34 VDD2.n24 171.744
R937 VDD2.n27 VDD2.n24 171.744
R938 VDD2.n6 VDD2.n3 171.744
R939 VDD2.n13 VDD2.n3 171.744
R940 VDD2.n14 VDD2.n13 171.744
R941 VDD2.n20 VDD2.n19 116.944
R942 VDD2 VDD2.n41 116.941
R943 VDD2.n27 VDD2.t5 85.8723
R944 VDD2.n6 VDD2.t2 85.8723
R945 VDD2.n20 VDD2.n18 53.6705
R946 VDD2.n40 VDD2.n39 51.5793
R947 VDD2.n40 VDD2.n20 36.4481
R948 VDD2.n28 VDD2.n26 16.3201
R949 VDD2.n7 VDD2.n5 16.3201
R950 VDD2.n29 VDD2.n25 12.8005
R951 VDD2.n8 VDD2.n4 12.8005
R952 VDD2.n33 VDD2.n32 12.0247
R953 VDD2.n12 VDD2.n11 12.0247
R954 VDD2.n36 VDD2.n23 11.249
R955 VDD2.n15 VDD2.n2 11.249
R956 VDD2.n37 VDD2.n21 10.4732
R957 VDD2.n16 VDD2.n0 10.4732
R958 VDD2.n39 VDD2.n38 9.45567
R959 VDD2.n18 VDD2.n17 9.45567
R960 VDD2.n38 VDD2.n37 9.3005
R961 VDD2.n23 VDD2.n22 9.3005
R962 VDD2.n32 VDD2.n31 9.3005
R963 VDD2.n30 VDD2.n29 9.3005
R964 VDD2.n17 VDD2.n16 9.3005
R965 VDD2.n2 VDD2.n1 9.3005
R966 VDD2.n11 VDD2.n10 9.3005
R967 VDD2.n9 VDD2.n8 9.3005
R968 VDD2.n41 VDD2.t3 8.16759
R969 VDD2.n41 VDD2.t1 8.16759
R970 VDD2.n19 VDD2.t0 8.16759
R971 VDD2.n19 VDD2.t4 8.16759
R972 VDD2.n30 VDD2.n26 3.78097
R973 VDD2.n9 VDD2.n5 3.78097
R974 VDD2.n39 VDD2.n21 3.49141
R975 VDD2.n18 VDD2.n0 3.49141
R976 VDD2.n37 VDD2.n36 2.71565
R977 VDD2.n16 VDD2.n15 2.71565
R978 VDD2 VDD2.n40 2.20524
R979 VDD2.n33 VDD2.n23 1.93989
R980 VDD2.n12 VDD2.n2 1.93989
R981 VDD2.n32 VDD2.n25 1.16414
R982 VDD2.n11 VDD2.n4 1.16414
R983 VDD2.n29 VDD2.n28 0.388379
R984 VDD2.n8 VDD2.n7 0.388379
R985 VDD2.n38 VDD2.n22 0.155672
R986 VDD2.n31 VDD2.n22 0.155672
R987 VDD2.n31 VDD2.n30 0.155672
R988 VDD2.n10 VDD2.n9 0.155672
R989 VDD2.n10 VDD2.n1 0.155672
R990 VDD2.n17 VDD2.n1 0.155672
R991 VTAIL.n82 VTAIL.n68 756.745
R992 VTAIL.n16 VTAIL.n2 756.745
R993 VTAIL.n62 VTAIL.n48 756.745
R994 VTAIL.n40 VTAIL.n26 756.745
R995 VTAIL.n75 VTAIL.n74 585
R996 VTAIL.n72 VTAIL.n71 585
R997 VTAIL.n81 VTAIL.n80 585
R998 VTAIL.n83 VTAIL.n82 585
R999 VTAIL.n9 VTAIL.n8 585
R1000 VTAIL.n6 VTAIL.n5 585
R1001 VTAIL.n15 VTAIL.n14 585
R1002 VTAIL.n17 VTAIL.n16 585
R1003 VTAIL.n63 VTAIL.n62 585
R1004 VTAIL.n61 VTAIL.n60 585
R1005 VTAIL.n52 VTAIL.n51 585
R1006 VTAIL.n55 VTAIL.n54 585
R1007 VTAIL.n41 VTAIL.n40 585
R1008 VTAIL.n39 VTAIL.n38 585
R1009 VTAIL.n30 VTAIL.n29 585
R1010 VTAIL.n33 VTAIL.n32 585
R1011 VTAIL.t7 VTAIL.n73 330.707
R1012 VTAIL.t11 VTAIL.n7 330.707
R1013 VTAIL.t0 VTAIL.n53 330.707
R1014 VTAIL.t6 VTAIL.n31 330.707
R1015 VTAIL.n74 VTAIL.n71 171.744
R1016 VTAIL.n81 VTAIL.n71 171.744
R1017 VTAIL.n82 VTAIL.n81 171.744
R1018 VTAIL.n8 VTAIL.n5 171.744
R1019 VTAIL.n15 VTAIL.n5 171.744
R1020 VTAIL.n16 VTAIL.n15 171.744
R1021 VTAIL.n62 VTAIL.n61 171.744
R1022 VTAIL.n61 VTAIL.n51 171.744
R1023 VTAIL.n54 VTAIL.n51 171.744
R1024 VTAIL.n40 VTAIL.n39 171.744
R1025 VTAIL.n39 VTAIL.n29 171.744
R1026 VTAIL.n32 VTAIL.n29 171.744
R1027 VTAIL.n47 VTAIL.n46 99.6047
R1028 VTAIL.n25 VTAIL.n24 99.6047
R1029 VTAIL.n1 VTAIL.n0 99.6045
R1030 VTAIL.n23 VTAIL.n22 99.6045
R1031 VTAIL.n74 VTAIL.t7 85.8723
R1032 VTAIL.n8 VTAIL.t11 85.8723
R1033 VTAIL.n54 VTAIL.t0 85.8723
R1034 VTAIL.n32 VTAIL.t6 85.8723
R1035 VTAIL.n87 VTAIL.n86 34.9005
R1036 VTAIL.n21 VTAIL.n20 34.9005
R1037 VTAIL.n67 VTAIL.n66 34.9005
R1038 VTAIL.n45 VTAIL.n44 34.9005
R1039 VTAIL.n25 VTAIL.n23 21.5221
R1040 VTAIL.n87 VTAIL.n67 18.66
R1041 VTAIL.n75 VTAIL.n73 16.3201
R1042 VTAIL.n9 VTAIL.n7 16.3201
R1043 VTAIL.n55 VTAIL.n53 16.3201
R1044 VTAIL.n33 VTAIL.n31 16.3201
R1045 VTAIL.n76 VTAIL.n72 12.8005
R1046 VTAIL.n10 VTAIL.n6 12.8005
R1047 VTAIL.n56 VTAIL.n52 12.8005
R1048 VTAIL.n34 VTAIL.n30 12.8005
R1049 VTAIL.n80 VTAIL.n79 12.0247
R1050 VTAIL.n14 VTAIL.n13 12.0247
R1051 VTAIL.n60 VTAIL.n59 12.0247
R1052 VTAIL.n38 VTAIL.n37 12.0247
R1053 VTAIL.n83 VTAIL.n70 11.249
R1054 VTAIL.n17 VTAIL.n4 11.249
R1055 VTAIL.n63 VTAIL.n50 11.249
R1056 VTAIL.n41 VTAIL.n28 11.249
R1057 VTAIL.n84 VTAIL.n68 10.4732
R1058 VTAIL.n18 VTAIL.n2 10.4732
R1059 VTAIL.n64 VTAIL.n48 10.4732
R1060 VTAIL.n42 VTAIL.n26 10.4732
R1061 VTAIL.n86 VTAIL.n85 9.45567
R1062 VTAIL.n20 VTAIL.n19 9.45567
R1063 VTAIL.n66 VTAIL.n65 9.45567
R1064 VTAIL.n44 VTAIL.n43 9.45567
R1065 VTAIL.n85 VTAIL.n84 9.3005
R1066 VTAIL.n70 VTAIL.n69 9.3005
R1067 VTAIL.n79 VTAIL.n78 9.3005
R1068 VTAIL.n77 VTAIL.n76 9.3005
R1069 VTAIL.n19 VTAIL.n18 9.3005
R1070 VTAIL.n4 VTAIL.n3 9.3005
R1071 VTAIL.n13 VTAIL.n12 9.3005
R1072 VTAIL.n11 VTAIL.n10 9.3005
R1073 VTAIL.n65 VTAIL.n64 9.3005
R1074 VTAIL.n50 VTAIL.n49 9.3005
R1075 VTAIL.n59 VTAIL.n58 9.3005
R1076 VTAIL.n57 VTAIL.n56 9.3005
R1077 VTAIL.n43 VTAIL.n42 9.3005
R1078 VTAIL.n28 VTAIL.n27 9.3005
R1079 VTAIL.n37 VTAIL.n36 9.3005
R1080 VTAIL.n35 VTAIL.n34 9.3005
R1081 VTAIL.n0 VTAIL.t3 8.16759
R1082 VTAIL.n0 VTAIL.t4 8.16759
R1083 VTAIL.n22 VTAIL.t2 8.16759
R1084 VTAIL.n22 VTAIL.t10 8.16759
R1085 VTAIL.n46 VTAIL.t9 8.16759
R1086 VTAIL.n46 VTAIL.t1 8.16759
R1087 VTAIL.n24 VTAIL.t5 8.16759
R1088 VTAIL.n24 VTAIL.t8 8.16759
R1089 VTAIL.n77 VTAIL.n73 3.78097
R1090 VTAIL.n11 VTAIL.n7 3.78097
R1091 VTAIL.n57 VTAIL.n53 3.78097
R1092 VTAIL.n35 VTAIL.n31 3.78097
R1093 VTAIL.n86 VTAIL.n68 3.49141
R1094 VTAIL.n20 VTAIL.n2 3.49141
R1095 VTAIL.n66 VTAIL.n48 3.49141
R1096 VTAIL.n44 VTAIL.n26 3.49141
R1097 VTAIL.n45 VTAIL.n25 2.86257
R1098 VTAIL.n67 VTAIL.n47 2.86257
R1099 VTAIL.n23 VTAIL.n21 2.86257
R1100 VTAIL.n84 VTAIL.n83 2.71565
R1101 VTAIL.n18 VTAIL.n17 2.71565
R1102 VTAIL.n64 VTAIL.n63 2.71565
R1103 VTAIL.n42 VTAIL.n41 2.71565
R1104 VTAIL VTAIL.n87 2.08886
R1105 VTAIL.n80 VTAIL.n70 1.93989
R1106 VTAIL.n14 VTAIL.n4 1.93989
R1107 VTAIL.n60 VTAIL.n50 1.93989
R1108 VTAIL.n38 VTAIL.n28 1.93989
R1109 VTAIL.n47 VTAIL.n45 1.90136
R1110 VTAIL.n21 VTAIL.n1 1.90136
R1111 VTAIL.n79 VTAIL.n72 1.16414
R1112 VTAIL.n13 VTAIL.n6 1.16414
R1113 VTAIL.n59 VTAIL.n52 1.16414
R1114 VTAIL.n37 VTAIL.n30 1.16414
R1115 VTAIL VTAIL.n1 0.774207
R1116 VTAIL.n76 VTAIL.n75 0.388379
R1117 VTAIL.n10 VTAIL.n9 0.388379
R1118 VTAIL.n56 VTAIL.n55 0.388379
R1119 VTAIL.n34 VTAIL.n33 0.388379
R1120 VTAIL.n78 VTAIL.n77 0.155672
R1121 VTAIL.n78 VTAIL.n69 0.155672
R1122 VTAIL.n85 VTAIL.n69 0.155672
R1123 VTAIL.n12 VTAIL.n11 0.155672
R1124 VTAIL.n12 VTAIL.n3 0.155672
R1125 VTAIL.n19 VTAIL.n3 0.155672
R1126 VTAIL.n65 VTAIL.n49 0.155672
R1127 VTAIL.n58 VTAIL.n49 0.155672
R1128 VTAIL.n58 VTAIL.n57 0.155672
R1129 VTAIL.n43 VTAIL.n27 0.155672
R1130 VTAIL.n36 VTAIL.n27 0.155672
R1131 VTAIL.n36 VTAIL.n35 0.155672
R1132 VP.n13 VP.n10 161.3
R1133 VP.n15 VP.n14 161.3
R1134 VP.n16 VP.n9 161.3
R1135 VP.n18 VP.n17 161.3
R1136 VP.n19 VP.n8 161.3
R1137 VP.n21 VP.n20 161.3
R1138 VP.n44 VP.n43 161.3
R1139 VP.n42 VP.n1 161.3
R1140 VP.n41 VP.n40 161.3
R1141 VP.n39 VP.n2 161.3
R1142 VP.n38 VP.n37 161.3
R1143 VP.n36 VP.n3 161.3
R1144 VP.n35 VP.n34 161.3
R1145 VP.n33 VP.n4 161.3
R1146 VP.n32 VP.n31 161.3
R1147 VP.n30 VP.n5 161.3
R1148 VP.n29 VP.n28 161.3
R1149 VP.n27 VP.n6 161.3
R1150 VP.n26 VP.n25 161.3
R1151 VP.n24 VP.n23 74.5068
R1152 VP.n45 VP.n0 74.5068
R1153 VP.n22 VP.n7 74.5068
R1154 VP.n11 VP.t0 65.3333
R1155 VP.n30 VP.n29 56.0773
R1156 VP.n41 VP.n2 56.0773
R1157 VP.n18 VP.n9 56.0773
R1158 VP.n12 VP.n11 49.3258
R1159 VP.n23 VP.n22 44.1814
R1160 VP.n35 VP.t2 32.0801
R1161 VP.n24 VP.t3 32.0801
R1162 VP.n0 VP.t1 32.0801
R1163 VP.n12 VP.t4 32.0801
R1164 VP.n7 VP.t5 32.0801
R1165 VP.n31 VP.n30 25.0767
R1166 VP.n37 VP.n2 25.0767
R1167 VP.n14 VP.n9 25.0767
R1168 VP.n25 VP.n6 24.5923
R1169 VP.n29 VP.n6 24.5923
R1170 VP.n31 VP.n4 24.5923
R1171 VP.n35 VP.n4 24.5923
R1172 VP.n36 VP.n35 24.5923
R1173 VP.n37 VP.n36 24.5923
R1174 VP.n42 VP.n41 24.5923
R1175 VP.n43 VP.n42 24.5923
R1176 VP.n19 VP.n18 24.5923
R1177 VP.n20 VP.n19 24.5923
R1178 VP.n13 VP.n12 24.5923
R1179 VP.n14 VP.n13 24.5923
R1180 VP.n25 VP.n24 15.7393
R1181 VP.n43 VP.n0 15.7393
R1182 VP.n20 VP.n7 15.7393
R1183 VP.n11 VP.n10 4.10785
R1184 VP.n22 VP.n21 0.354861
R1185 VP.n26 VP.n23 0.354861
R1186 VP.n45 VP.n44 0.354861
R1187 VP VP.n45 0.267071
R1188 VP.n15 VP.n10 0.189894
R1189 VP.n16 VP.n15 0.189894
R1190 VP.n17 VP.n16 0.189894
R1191 VP.n17 VP.n8 0.189894
R1192 VP.n21 VP.n8 0.189894
R1193 VP.n27 VP.n26 0.189894
R1194 VP.n28 VP.n27 0.189894
R1195 VP.n28 VP.n5 0.189894
R1196 VP.n32 VP.n5 0.189894
R1197 VP.n33 VP.n32 0.189894
R1198 VP.n34 VP.n33 0.189894
R1199 VP.n34 VP.n3 0.189894
R1200 VP.n38 VP.n3 0.189894
R1201 VP.n39 VP.n38 0.189894
R1202 VP.n40 VP.n39 0.189894
R1203 VP.n40 VP.n1 0.189894
R1204 VP.n44 VP.n1 0.189894
R1205 VDD1.n14 VDD1.n0 756.745
R1206 VDD1.n33 VDD1.n19 756.745
R1207 VDD1.n15 VDD1.n14 585
R1208 VDD1.n13 VDD1.n12 585
R1209 VDD1.n4 VDD1.n3 585
R1210 VDD1.n7 VDD1.n6 585
R1211 VDD1.n26 VDD1.n25 585
R1212 VDD1.n23 VDD1.n22 585
R1213 VDD1.n32 VDD1.n31 585
R1214 VDD1.n34 VDD1.n33 585
R1215 VDD1.t5 VDD1.n5 330.707
R1216 VDD1.t2 VDD1.n24 330.707
R1217 VDD1.n14 VDD1.n13 171.744
R1218 VDD1.n13 VDD1.n3 171.744
R1219 VDD1.n6 VDD1.n3 171.744
R1220 VDD1.n25 VDD1.n22 171.744
R1221 VDD1.n32 VDD1.n22 171.744
R1222 VDD1.n33 VDD1.n32 171.744
R1223 VDD1.n39 VDD1.n38 116.944
R1224 VDD1.n41 VDD1.n40 116.284
R1225 VDD1.n6 VDD1.t5 85.8723
R1226 VDD1.n25 VDD1.t2 85.8723
R1227 VDD1 VDD1.n18 53.784
R1228 VDD1.n39 VDD1.n37 53.6705
R1229 VDD1.n41 VDD1.n39 38.4621
R1230 VDD1.n7 VDD1.n5 16.3201
R1231 VDD1.n26 VDD1.n24 16.3201
R1232 VDD1.n8 VDD1.n4 12.8005
R1233 VDD1.n27 VDD1.n23 12.8005
R1234 VDD1.n12 VDD1.n11 12.0247
R1235 VDD1.n31 VDD1.n30 12.0247
R1236 VDD1.n15 VDD1.n2 11.249
R1237 VDD1.n34 VDD1.n21 11.249
R1238 VDD1.n16 VDD1.n0 10.4732
R1239 VDD1.n35 VDD1.n19 10.4732
R1240 VDD1.n18 VDD1.n17 9.45567
R1241 VDD1.n37 VDD1.n36 9.45567
R1242 VDD1.n17 VDD1.n16 9.3005
R1243 VDD1.n2 VDD1.n1 9.3005
R1244 VDD1.n11 VDD1.n10 9.3005
R1245 VDD1.n9 VDD1.n8 9.3005
R1246 VDD1.n36 VDD1.n35 9.3005
R1247 VDD1.n21 VDD1.n20 9.3005
R1248 VDD1.n30 VDD1.n29 9.3005
R1249 VDD1.n28 VDD1.n27 9.3005
R1250 VDD1.n40 VDD1.t1 8.16759
R1251 VDD1.n40 VDD1.t0 8.16759
R1252 VDD1.n38 VDD1.t3 8.16759
R1253 VDD1.n38 VDD1.t4 8.16759
R1254 VDD1.n9 VDD1.n5 3.78097
R1255 VDD1.n28 VDD1.n24 3.78097
R1256 VDD1.n18 VDD1.n0 3.49141
R1257 VDD1.n37 VDD1.n19 3.49141
R1258 VDD1.n16 VDD1.n15 2.71565
R1259 VDD1.n35 VDD1.n34 2.71565
R1260 VDD1.n12 VDD1.n2 1.93989
R1261 VDD1.n31 VDD1.n21 1.93989
R1262 VDD1.n11 VDD1.n4 1.16414
R1263 VDD1.n30 VDD1.n23 1.16414
R1264 VDD1 VDD1.n41 0.657828
R1265 VDD1.n8 VDD1.n7 0.388379
R1266 VDD1.n27 VDD1.n26 0.388379
R1267 VDD1.n17 VDD1.n1 0.155672
R1268 VDD1.n10 VDD1.n1 0.155672
R1269 VDD1.n10 VDD1.n9 0.155672
R1270 VDD1.n29 VDD1.n28 0.155672
R1271 VDD1.n29 VDD1.n20 0.155672
R1272 VDD1.n36 VDD1.n20 0.155672
C0 VN VP 5.825991f
C1 VDD1 VN 0.15597f
C2 VP VTAIL 3.37922f
C3 VN w_n3626_n1764# 6.82365f
C4 VDD1 VTAIL 5.06189f
C5 VN VDD2 2.54893f
C6 w_n3626_n1764# VTAIL 1.88606f
C7 VN B 1.17805f
C8 VDD2 VTAIL 5.11734f
C9 VTAIL B 1.96405f
C10 VDD1 VP 2.88649f
C11 VP w_n3626_n1764# 7.292601f
C12 VP VDD2 0.496077f
C13 VDD1 w_n3626_n1764# 1.83188f
C14 VDD1 VDD2 1.55874f
C15 VN VTAIL 3.36506f
C16 VP B 1.96433f
C17 VDD1 B 1.55574f
C18 w_n3626_n1764# VDD2 1.92902f
C19 w_n3626_n1764# B 7.988379f
C20 VDD2 B 1.63936f
C21 VDD2 VSUBS 1.421904f
C22 VDD1 VSUBS 1.625281f
C23 VTAIL VSUBS 0.614649f
C24 VN VSUBS 6.01419f
C25 VP VSUBS 2.716431f
C26 B VSUBS 4.089189f
C27 w_n3626_n1764# VSUBS 80.5407f
C28 VDD1.n0 VSUBS 0.025244f
C29 VDD1.n1 VSUBS 0.022885f
C30 VDD1.n2 VSUBS 0.012297f
C31 VDD1.n3 VSUBS 0.029066f
C32 VDD1.n4 VSUBS 0.013021f
C33 VDD1.n5 VSUBS 0.08914f
C34 VDD1.t5 VSUBS 0.064495f
C35 VDD1.n6 VSUBS 0.021799f
C36 VDD1.n7 VSUBS 0.018282f
C37 VDD1.n8 VSUBS 0.012297f
C38 VDD1.n9 VSUBS 0.311464f
C39 VDD1.n10 VSUBS 0.022885f
C40 VDD1.n11 VSUBS 0.012297f
C41 VDD1.n12 VSUBS 0.013021f
C42 VDD1.n13 VSUBS 0.029066f
C43 VDD1.n14 VSUBS 0.070701f
C44 VDD1.n15 VSUBS 0.013021f
C45 VDD1.n16 VSUBS 0.012297f
C46 VDD1.n17 VSUBS 0.057273f
C47 VDD1.n18 VSUBS 0.060043f
C48 VDD1.n19 VSUBS 0.025244f
C49 VDD1.n20 VSUBS 0.022885f
C50 VDD1.n21 VSUBS 0.012297f
C51 VDD1.n22 VSUBS 0.029066f
C52 VDD1.n23 VSUBS 0.013021f
C53 VDD1.n24 VSUBS 0.08914f
C54 VDD1.t2 VSUBS 0.064495f
C55 VDD1.n25 VSUBS 0.021799f
C56 VDD1.n26 VSUBS 0.018282f
C57 VDD1.n27 VSUBS 0.012297f
C58 VDD1.n28 VSUBS 0.311464f
C59 VDD1.n29 VSUBS 0.022885f
C60 VDD1.n30 VSUBS 0.012297f
C61 VDD1.n31 VSUBS 0.013021f
C62 VDD1.n32 VSUBS 0.029066f
C63 VDD1.n33 VSUBS 0.070701f
C64 VDD1.n34 VSUBS 0.013021f
C65 VDD1.n35 VSUBS 0.012297f
C66 VDD1.n36 VSUBS 0.057273f
C67 VDD1.n37 VSUBS 0.059302f
C68 VDD1.t3 VSUBS 0.071975f
C69 VDD1.t4 VSUBS 0.071975f
C70 VDD1.n38 VSUBS 0.423436f
C71 VDD1.n39 VSUBS 2.41645f
C72 VDD1.t1 VSUBS 0.071975f
C73 VDD1.t0 VSUBS 0.071975f
C74 VDD1.n40 VSUBS 0.42009f
C75 VDD1.n41 VSUBS 2.22006f
C76 VP.t1 VSUBS 1.33658f
C77 VP.n0 VSUBS 0.685276f
C78 VP.n1 VSUBS 0.043741f
C79 VP.n2 VSUBS 0.052042f
C80 VP.n3 VSUBS 0.043741f
C81 VP.t2 VSUBS 1.33658f
C82 VP.n4 VSUBS 0.081113f
C83 VP.n5 VSUBS 0.043741f
C84 VP.n6 VSUBS 0.081113f
C85 VP.t5 VSUBS 1.33658f
C86 VP.n7 VSUBS 0.685276f
C87 VP.n8 VSUBS 0.043741f
C88 VP.n9 VSUBS 0.052042f
C89 VP.n10 VSUBS 0.496567f
C90 VP.t4 VSUBS 1.33658f
C91 VP.t0 VSUBS 1.75463f
C92 VP.n11 VSUBS 0.642124f
C93 VP.n12 VSUBS 0.686893f
C94 VP.n13 VSUBS 0.081113f
C95 VP.n14 VSUBS 0.081871f
C96 VP.n15 VSUBS 0.043741f
C97 VP.n16 VSUBS 0.043741f
C98 VP.n17 VSUBS 0.043741f
C99 VP.n18 VSUBS 0.074368f
C100 VP.n19 VSUBS 0.081113f
C101 VP.n20 VSUBS 0.066698f
C102 VP.n21 VSUBS 0.070585f
C103 VP.n22 VSUBS 2.06076f
C104 VP.n23 VSUBS 2.09645f
C105 VP.t3 VSUBS 1.33658f
C106 VP.n24 VSUBS 0.685276f
C107 VP.n25 VSUBS 0.066698f
C108 VP.n26 VSUBS 0.070585f
C109 VP.n27 VSUBS 0.043741f
C110 VP.n28 VSUBS 0.043741f
C111 VP.n29 VSUBS 0.074368f
C112 VP.n30 VSUBS 0.052042f
C113 VP.n31 VSUBS 0.081871f
C114 VP.n32 VSUBS 0.043741f
C115 VP.n33 VSUBS 0.043741f
C116 VP.n34 VSUBS 0.043741f
C117 VP.n35 VSUBS 0.567363f
C118 VP.n36 VSUBS 0.081113f
C119 VP.n37 VSUBS 0.081871f
C120 VP.n38 VSUBS 0.043741f
C121 VP.n39 VSUBS 0.043741f
C122 VP.n40 VSUBS 0.043741f
C123 VP.n41 VSUBS 0.074368f
C124 VP.n42 VSUBS 0.081113f
C125 VP.n43 VSUBS 0.066698f
C126 VP.n44 VSUBS 0.070585f
C127 VP.n45 VSUBS 0.098623f
C128 VTAIL.t3 VSUBS 0.095386f
C129 VTAIL.t4 VSUBS 0.095386f
C130 VTAIL.n0 VSUBS 0.486024f
C131 VTAIL.n1 VSUBS 0.718909f
C132 VTAIL.n2 VSUBS 0.033455f
C133 VTAIL.n3 VSUBS 0.030328f
C134 VTAIL.n4 VSUBS 0.016297f
C135 VTAIL.n5 VSUBS 0.03852f
C136 VTAIL.n6 VSUBS 0.017256f
C137 VTAIL.n7 VSUBS 0.118135f
C138 VTAIL.t11 VSUBS 0.085474f
C139 VTAIL.n8 VSUBS 0.02889f
C140 VTAIL.n9 VSUBS 0.024229f
C141 VTAIL.n10 VSUBS 0.016297f
C142 VTAIL.n11 VSUBS 0.412775f
C143 VTAIL.n12 VSUBS 0.030328f
C144 VTAIL.n13 VSUBS 0.016297f
C145 VTAIL.n14 VSUBS 0.017256f
C146 VTAIL.n15 VSUBS 0.03852f
C147 VTAIL.n16 VSUBS 0.093698f
C148 VTAIL.n17 VSUBS 0.017256f
C149 VTAIL.n18 VSUBS 0.016297f
C150 VTAIL.n19 VSUBS 0.075903f
C151 VTAIL.n20 VSUBS 0.047311f
C152 VTAIL.n21 VSUBS 0.494638f
C153 VTAIL.t2 VSUBS 0.095386f
C154 VTAIL.t10 VSUBS 0.095386f
C155 VTAIL.n22 VSUBS 0.486024f
C156 VTAIL.n23 VSUBS 2.04389f
C157 VTAIL.t5 VSUBS 0.095386f
C158 VTAIL.t8 VSUBS 0.095386f
C159 VTAIL.n24 VSUBS 0.486027f
C160 VTAIL.n25 VSUBS 2.04389f
C161 VTAIL.n26 VSUBS 0.033455f
C162 VTAIL.n27 VSUBS 0.030328f
C163 VTAIL.n28 VSUBS 0.016297f
C164 VTAIL.n29 VSUBS 0.03852f
C165 VTAIL.n30 VSUBS 0.017256f
C166 VTAIL.n31 VSUBS 0.118135f
C167 VTAIL.t6 VSUBS 0.085474f
C168 VTAIL.n32 VSUBS 0.02889f
C169 VTAIL.n33 VSUBS 0.024229f
C170 VTAIL.n34 VSUBS 0.016297f
C171 VTAIL.n35 VSUBS 0.412775f
C172 VTAIL.n36 VSUBS 0.030328f
C173 VTAIL.n37 VSUBS 0.016297f
C174 VTAIL.n38 VSUBS 0.017256f
C175 VTAIL.n39 VSUBS 0.03852f
C176 VTAIL.n40 VSUBS 0.093698f
C177 VTAIL.n41 VSUBS 0.017256f
C178 VTAIL.n42 VSUBS 0.016297f
C179 VTAIL.n43 VSUBS 0.075903f
C180 VTAIL.n44 VSUBS 0.047311f
C181 VTAIL.n45 VSUBS 0.494638f
C182 VTAIL.t9 VSUBS 0.095386f
C183 VTAIL.t1 VSUBS 0.095386f
C184 VTAIL.n46 VSUBS 0.486027f
C185 VTAIL.n47 VSUBS 0.92299f
C186 VTAIL.n48 VSUBS 0.033455f
C187 VTAIL.n49 VSUBS 0.030328f
C188 VTAIL.n50 VSUBS 0.016297f
C189 VTAIL.n51 VSUBS 0.03852f
C190 VTAIL.n52 VSUBS 0.017256f
C191 VTAIL.n53 VSUBS 0.118135f
C192 VTAIL.t0 VSUBS 0.085474f
C193 VTAIL.n54 VSUBS 0.02889f
C194 VTAIL.n55 VSUBS 0.024229f
C195 VTAIL.n56 VSUBS 0.016297f
C196 VTAIL.n57 VSUBS 0.412775f
C197 VTAIL.n58 VSUBS 0.030328f
C198 VTAIL.n59 VSUBS 0.016297f
C199 VTAIL.n60 VSUBS 0.017256f
C200 VTAIL.n61 VSUBS 0.03852f
C201 VTAIL.n62 VSUBS 0.093698f
C202 VTAIL.n63 VSUBS 0.017256f
C203 VTAIL.n64 VSUBS 0.016297f
C204 VTAIL.n65 VSUBS 0.075903f
C205 VTAIL.n66 VSUBS 0.047311f
C206 VTAIL.n67 VSUBS 1.33584f
C207 VTAIL.n68 VSUBS 0.033455f
C208 VTAIL.n69 VSUBS 0.030328f
C209 VTAIL.n70 VSUBS 0.016297f
C210 VTAIL.n71 VSUBS 0.03852f
C211 VTAIL.n72 VSUBS 0.017256f
C212 VTAIL.n73 VSUBS 0.118135f
C213 VTAIL.t7 VSUBS 0.085474f
C214 VTAIL.n74 VSUBS 0.02889f
C215 VTAIL.n75 VSUBS 0.024229f
C216 VTAIL.n76 VSUBS 0.016297f
C217 VTAIL.n77 VSUBS 0.412775f
C218 VTAIL.n78 VSUBS 0.030328f
C219 VTAIL.n79 VSUBS 0.016297f
C220 VTAIL.n80 VSUBS 0.017256f
C221 VTAIL.n81 VSUBS 0.03852f
C222 VTAIL.n82 VSUBS 0.093698f
C223 VTAIL.n83 VSUBS 0.017256f
C224 VTAIL.n84 VSUBS 0.016297f
C225 VTAIL.n85 VSUBS 0.075903f
C226 VTAIL.n86 VSUBS 0.047311f
C227 VTAIL.n87 VSUBS 1.26023f
C228 VDD2.n0 VSUBS 0.024237f
C229 VDD2.n1 VSUBS 0.021972f
C230 VDD2.n2 VSUBS 0.011807f
C231 VDD2.n3 VSUBS 0.027908f
C232 VDD2.n4 VSUBS 0.012502f
C233 VDD2.n5 VSUBS 0.085588f
C234 VDD2.t2 VSUBS 0.061925f
C235 VDD2.n6 VSUBS 0.020931f
C236 VDD2.n7 VSUBS 0.017553f
C237 VDD2.n8 VSUBS 0.011807f
C238 VDD2.n9 VSUBS 0.299051f
C239 VDD2.n10 VSUBS 0.021972f
C240 VDD2.n11 VSUBS 0.011807f
C241 VDD2.n12 VSUBS 0.012502f
C242 VDD2.n13 VSUBS 0.027908f
C243 VDD2.n14 VSUBS 0.067883f
C244 VDD2.n15 VSUBS 0.012502f
C245 VDD2.n16 VSUBS 0.011807f
C246 VDD2.n17 VSUBS 0.054991f
C247 VDD2.n18 VSUBS 0.056938f
C248 VDD2.t0 VSUBS 0.069106f
C249 VDD2.t4 VSUBS 0.069106f
C250 VDD2.n19 VSUBS 0.40656f
C251 VDD2.n20 VSUBS 2.20955f
C252 VDD2.n21 VSUBS 0.024237f
C253 VDD2.n22 VSUBS 0.021972f
C254 VDD2.n23 VSUBS 0.011807f
C255 VDD2.n24 VSUBS 0.027908f
C256 VDD2.n25 VSUBS 0.012502f
C257 VDD2.n26 VSUBS 0.085588f
C258 VDD2.t5 VSUBS 0.061925f
C259 VDD2.n27 VSUBS 0.020931f
C260 VDD2.n28 VSUBS 0.017553f
C261 VDD2.n29 VSUBS 0.011807f
C262 VDD2.n30 VSUBS 0.299051f
C263 VDD2.n31 VSUBS 0.021972f
C264 VDD2.n32 VSUBS 0.011807f
C265 VDD2.n33 VSUBS 0.012502f
C266 VDD2.n34 VSUBS 0.027908f
C267 VDD2.n35 VSUBS 0.067883f
C268 VDD2.n36 VSUBS 0.012502f
C269 VDD2.n37 VSUBS 0.011807f
C270 VDD2.n38 VSUBS 0.054991f
C271 VDD2.n39 VSUBS 0.049418f
C272 VDD2.n40 VSUBS 1.79368f
C273 VDD2.t3 VSUBS 0.069106f
C274 VDD2.t1 VSUBS 0.069106f
C275 VDD2.n41 VSUBS 0.406541f
C276 VN.t1 VSUBS 1.27054f
C277 VN.n0 VSUBS 0.65142f
C278 VN.n1 VSUBS 0.04158f
C279 VN.n2 VSUBS 0.04947f
C280 VN.n3 VSUBS 0.472034f
C281 VN.t4 VSUBS 1.27054f
C282 VN.t5 VSUBS 1.66795f
C283 VN.n4 VSUBS 0.610399f
C284 VN.n5 VSUBS 0.652957f
C285 VN.n6 VSUBS 0.077106f
C286 VN.n7 VSUBS 0.077826f
C287 VN.n8 VSUBS 0.04158f
C288 VN.n9 VSUBS 0.04158f
C289 VN.n10 VSUBS 0.04158f
C290 VN.n11 VSUBS 0.070694f
C291 VN.n12 VSUBS 0.077106f
C292 VN.n13 VSUBS 0.063402f
C293 VN.n14 VSUBS 0.067098f
C294 VN.n15 VSUBS 0.09375f
C295 VN.t3 VSUBS 1.27054f
C296 VN.n16 VSUBS 0.65142f
C297 VN.n17 VSUBS 0.04158f
C298 VN.n18 VSUBS 0.04947f
C299 VN.n19 VSUBS 0.472034f
C300 VN.t0 VSUBS 1.27054f
C301 VN.t2 VSUBS 1.66795f
C302 VN.n20 VSUBS 0.610399f
C303 VN.n21 VSUBS 0.652957f
C304 VN.n22 VSUBS 0.077106f
C305 VN.n23 VSUBS 0.077826f
C306 VN.n24 VSUBS 0.04158f
C307 VN.n25 VSUBS 0.04158f
C308 VN.n26 VSUBS 0.04158f
C309 VN.n27 VSUBS 0.070694f
C310 VN.n28 VSUBS 0.077106f
C311 VN.n29 VSUBS 0.063402f
C312 VN.n30 VSUBS 0.067098f
C313 VN.n31 VSUBS 1.97675f
C314 B.n0 VSUBS 0.004406f
C315 B.n1 VSUBS 0.004406f
C316 B.n2 VSUBS 0.006967f
C317 B.n3 VSUBS 0.006967f
C318 B.n4 VSUBS 0.006967f
C319 B.n5 VSUBS 0.006967f
C320 B.n6 VSUBS 0.006967f
C321 B.n7 VSUBS 0.006967f
C322 B.n8 VSUBS 0.006967f
C323 B.n9 VSUBS 0.006967f
C324 B.n10 VSUBS 0.006967f
C325 B.n11 VSUBS 0.006967f
C326 B.n12 VSUBS 0.006967f
C327 B.n13 VSUBS 0.006967f
C328 B.n14 VSUBS 0.006967f
C329 B.n15 VSUBS 0.006967f
C330 B.n16 VSUBS 0.006967f
C331 B.n17 VSUBS 0.006967f
C332 B.n18 VSUBS 0.006967f
C333 B.n19 VSUBS 0.006967f
C334 B.n20 VSUBS 0.006967f
C335 B.n21 VSUBS 0.006967f
C336 B.n22 VSUBS 0.006967f
C337 B.n23 VSUBS 0.006967f
C338 B.n24 VSUBS 0.006967f
C339 B.n25 VSUBS 0.015549f
C340 B.n26 VSUBS 0.006967f
C341 B.n27 VSUBS 0.006967f
C342 B.n28 VSUBS 0.006967f
C343 B.n29 VSUBS 0.006967f
C344 B.n30 VSUBS 0.006967f
C345 B.n31 VSUBS 0.006967f
C346 B.n32 VSUBS 0.006967f
C347 B.n33 VSUBS 0.006967f
C348 B.n34 VSUBS 0.006557f
C349 B.n35 VSUBS 0.006967f
C350 B.t11 VSUBS 0.057463f
C351 B.t10 VSUBS 0.080303f
C352 B.t9 VSUBS 0.572767f
C353 B.n36 VSUBS 0.138245f
C354 B.n37 VSUBS 0.116224f
C355 B.n38 VSUBS 0.016142f
C356 B.n39 VSUBS 0.006967f
C357 B.n40 VSUBS 0.006967f
C358 B.n41 VSUBS 0.006967f
C359 B.n42 VSUBS 0.006967f
C360 B.t5 VSUBS 0.057464f
C361 B.t4 VSUBS 0.080304f
C362 B.t3 VSUBS 0.572767f
C363 B.n43 VSUBS 0.138245f
C364 B.n44 VSUBS 0.116223f
C365 B.n45 VSUBS 0.006967f
C366 B.n46 VSUBS 0.006967f
C367 B.n47 VSUBS 0.006967f
C368 B.n48 VSUBS 0.006967f
C369 B.n49 VSUBS 0.006967f
C370 B.n50 VSUBS 0.006967f
C371 B.n51 VSUBS 0.006967f
C372 B.n52 VSUBS 0.006967f
C373 B.n53 VSUBS 0.015995f
C374 B.n54 VSUBS 0.006967f
C375 B.n55 VSUBS 0.006967f
C376 B.n56 VSUBS 0.006967f
C377 B.n57 VSUBS 0.006967f
C378 B.n58 VSUBS 0.006967f
C379 B.n59 VSUBS 0.006967f
C380 B.n60 VSUBS 0.006967f
C381 B.n61 VSUBS 0.006967f
C382 B.n62 VSUBS 0.006967f
C383 B.n63 VSUBS 0.006967f
C384 B.n64 VSUBS 0.006967f
C385 B.n65 VSUBS 0.006967f
C386 B.n66 VSUBS 0.006967f
C387 B.n67 VSUBS 0.006967f
C388 B.n68 VSUBS 0.006967f
C389 B.n69 VSUBS 0.006967f
C390 B.n70 VSUBS 0.006967f
C391 B.n71 VSUBS 0.006967f
C392 B.n72 VSUBS 0.006967f
C393 B.n73 VSUBS 0.006967f
C394 B.n74 VSUBS 0.006967f
C395 B.n75 VSUBS 0.006967f
C396 B.n76 VSUBS 0.006967f
C397 B.n77 VSUBS 0.006967f
C398 B.n78 VSUBS 0.006967f
C399 B.n79 VSUBS 0.006967f
C400 B.n80 VSUBS 0.006967f
C401 B.n81 VSUBS 0.006967f
C402 B.n82 VSUBS 0.006967f
C403 B.n83 VSUBS 0.006967f
C404 B.n84 VSUBS 0.006967f
C405 B.n85 VSUBS 0.006967f
C406 B.n86 VSUBS 0.006967f
C407 B.n87 VSUBS 0.006967f
C408 B.n88 VSUBS 0.006967f
C409 B.n89 VSUBS 0.006967f
C410 B.n90 VSUBS 0.006967f
C411 B.n91 VSUBS 0.006967f
C412 B.n92 VSUBS 0.006967f
C413 B.n93 VSUBS 0.006967f
C414 B.n94 VSUBS 0.006967f
C415 B.n95 VSUBS 0.006967f
C416 B.n96 VSUBS 0.006967f
C417 B.n97 VSUBS 0.006967f
C418 B.n98 VSUBS 0.006967f
C419 B.n99 VSUBS 0.006967f
C420 B.n100 VSUBS 0.006967f
C421 B.n101 VSUBS 0.016827f
C422 B.n102 VSUBS 0.006967f
C423 B.n103 VSUBS 0.006967f
C424 B.n104 VSUBS 0.006967f
C425 B.n105 VSUBS 0.006967f
C426 B.n106 VSUBS 0.006967f
C427 B.n107 VSUBS 0.006967f
C428 B.n108 VSUBS 0.006967f
C429 B.n109 VSUBS 0.006967f
C430 B.n110 VSUBS 0.006967f
C431 B.t1 VSUBS 0.057464f
C432 B.t2 VSUBS 0.080304f
C433 B.t0 VSUBS 0.572767f
C434 B.n111 VSUBS 0.138245f
C435 B.n112 VSUBS 0.116223f
C436 B.n113 VSUBS 0.006967f
C437 B.n114 VSUBS 0.006967f
C438 B.n115 VSUBS 0.006967f
C439 B.n116 VSUBS 0.006967f
C440 B.t7 VSUBS 0.057463f
C441 B.t8 VSUBS 0.080303f
C442 B.t6 VSUBS 0.572767f
C443 B.n117 VSUBS 0.138245f
C444 B.n118 VSUBS 0.116224f
C445 B.n119 VSUBS 0.016142f
C446 B.n120 VSUBS 0.006967f
C447 B.n121 VSUBS 0.006967f
C448 B.n122 VSUBS 0.006967f
C449 B.n123 VSUBS 0.006967f
C450 B.n124 VSUBS 0.006967f
C451 B.n125 VSUBS 0.006967f
C452 B.n126 VSUBS 0.006967f
C453 B.n127 VSUBS 0.006967f
C454 B.n128 VSUBS 0.016827f
C455 B.n129 VSUBS 0.006967f
C456 B.n130 VSUBS 0.006967f
C457 B.n131 VSUBS 0.006967f
C458 B.n132 VSUBS 0.006967f
C459 B.n133 VSUBS 0.006967f
C460 B.n134 VSUBS 0.006967f
C461 B.n135 VSUBS 0.006967f
C462 B.n136 VSUBS 0.006967f
C463 B.n137 VSUBS 0.006967f
C464 B.n138 VSUBS 0.006967f
C465 B.n139 VSUBS 0.006967f
C466 B.n140 VSUBS 0.006967f
C467 B.n141 VSUBS 0.006967f
C468 B.n142 VSUBS 0.006967f
C469 B.n143 VSUBS 0.006967f
C470 B.n144 VSUBS 0.006967f
C471 B.n145 VSUBS 0.006967f
C472 B.n146 VSUBS 0.006967f
C473 B.n147 VSUBS 0.006967f
C474 B.n148 VSUBS 0.006967f
C475 B.n149 VSUBS 0.006967f
C476 B.n150 VSUBS 0.006967f
C477 B.n151 VSUBS 0.006967f
C478 B.n152 VSUBS 0.006967f
C479 B.n153 VSUBS 0.006967f
C480 B.n154 VSUBS 0.006967f
C481 B.n155 VSUBS 0.006967f
C482 B.n156 VSUBS 0.006967f
C483 B.n157 VSUBS 0.006967f
C484 B.n158 VSUBS 0.006967f
C485 B.n159 VSUBS 0.006967f
C486 B.n160 VSUBS 0.006967f
C487 B.n161 VSUBS 0.006967f
C488 B.n162 VSUBS 0.006967f
C489 B.n163 VSUBS 0.006967f
C490 B.n164 VSUBS 0.006967f
C491 B.n165 VSUBS 0.006967f
C492 B.n166 VSUBS 0.006967f
C493 B.n167 VSUBS 0.006967f
C494 B.n168 VSUBS 0.006967f
C495 B.n169 VSUBS 0.006967f
C496 B.n170 VSUBS 0.006967f
C497 B.n171 VSUBS 0.006967f
C498 B.n172 VSUBS 0.006967f
C499 B.n173 VSUBS 0.006967f
C500 B.n174 VSUBS 0.006967f
C501 B.n175 VSUBS 0.006967f
C502 B.n176 VSUBS 0.006967f
C503 B.n177 VSUBS 0.006967f
C504 B.n178 VSUBS 0.006967f
C505 B.n179 VSUBS 0.006967f
C506 B.n180 VSUBS 0.006967f
C507 B.n181 VSUBS 0.006967f
C508 B.n182 VSUBS 0.006967f
C509 B.n183 VSUBS 0.006967f
C510 B.n184 VSUBS 0.006967f
C511 B.n185 VSUBS 0.006967f
C512 B.n186 VSUBS 0.006967f
C513 B.n187 VSUBS 0.006967f
C514 B.n188 VSUBS 0.006967f
C515 B.n189 VSUBS 0.006967f
C516 B.n190 VSUBS 0.006967f
C517 B.n191 VSUBS 0.006967f
C518 B.n192 VSUBS 0.006967f
C519 B.n193 VSUBS 0.006967f
C520 B.n194 VSUBS 0.006967f
C521 B.n195 VSUBS 0.006967f
C522 B.n196 VSUBS 0.006967f
C523 B.n197 VSUBS 0.006967f
C524 B.n198 VSUBS 0.006967f
C525 B.n199 VSUBS 0.006967f
C526 B.n200 VSUBS 0.006967f
C527 B.n201 VSUBS 0.006967f
C528 B.n202 VSUBS 0.006967f
C529 B.n203 VSUBS 0.006967f
C530 B.n204 VSUBS 0.006967f
C531 B.n205 VSUBS 0.006967f
C532 B.n206 VSUBS 0.006967f
C533 B.n207 VSUBS 0.006967f
C534 B.n208 VSUBS 0.006967f
C535 B.n209 VSUBS 0.006967f
C536 B.n210 VSUBS 0.006967f
C537 B.n211 VSUBS 0.006967f
C538 B.n212 VSUBS 0.006967f
C539 B.n213 VSUBS 0.006967f
C540 B.n214 VSUBS 0.006967f
C541 B.n215 VSUBS 0.006967f
C542 B.n216 VSUBS 0.006967f
C543 B.n217 VSUBS 0.006967f
C544 B.n218 VSUBS 0.006967f
C545 B.n219 VSUBS 0.015549f
C546 B.n220 VSUBS 0.015549f
C547 B.n221 VSUBS 0.016827f
C548 B.n222 VSUBS 0.006967f
C549 B.n223 VSUBS 0.006967f
C550 B.n224 VSUBS 0.006967f
C551 B.n225 VSUBS 0.006967f
C552 B.n226 VSUBS 0.006967f
C553 B.n227 VSUBS 0.006967f
C554 B.n228 VSUBS 0.006967f
C555 B.n229 VSUBS 0.006967f
C556 B.n230 VSUBS 0.006967f
C557 B.n231 VSUBS 0.006967f
C558 B.n232 VSUBS 0.006967f
C559 B.n233 VSUBS 0.006967f
C560 B.n234 VSUBS 0.006967f
C561 B.n235 VSUBS 0.006967f
C562 B.n236 VSUBS 0.006967f
C563 B.n237 VSUBS 0.006967f
C564 B.n238 VSUBS 0.006967f
C565 B.n239 VSUBS 0.006967f
C566 B.n240 VSUBS 0.006967f
C567 B.n241 VSUBS 0.006967f
C568 B.n242 VSUBS 0.006967f
C569 B.n243 VSUBS 0.006967f
C570 B.n244 VSUBS 0.006967f
C571 B.n245 VSUBS 0.006967f
C572 B.n246 VSUBS 0.006557f
C573 B.n247 VSUBS 0.006967f
C574 B.n248 VSUBS 0.006967f
C575 B.n249 VSUBS 0.003893f
C576 B.n250 VSUBS 0.006967f
C577 B.n251 VSUBS 0.006967f
C578 B.n252 VSUBS 0.006967f
C579 B.n253 VSUBS 0.006967f
C580 B.n254 VSUBS 0.006967f
C581 B.n255 VSUBS 0.006967f
C582 B.n256 VSUBS 0.006967f
C583 B.n257 VSUBS 0.006967f
C584 B.n258 VSUBS 0.006967f
C585 B.n259 VSUBS 0.006967f
C586 B.n260 VSUBS 0.006967f
C587 B.n261 VSUBS 0.006967f
C588 B.n262 VSUBS 0.003893f
C589 B.n263 VSUBS 0.016142f
C590 B.n264 VSUBS 0.006557f
C591 B.n265 VSUBS 0.006967f
C592 B.n266 VSUBS 0.006967f
C593 B.n267 VSUBS 0.006967f
C594 B.n268 VSUBS 0.006967f
C595 B.n269 VSUBS 0.006967f
C596 B.n270 VSUBS 0.006967f
C597 B.n271 VSUBS 0.006967f
C598 B.n272 VSUBS 0.006967f
C599 B.n273 VSUBS 0.006967f
C600 B.n274 VSUBS 0.006967f
C601 B.n275 VSUBS 0.006967f
C602 B.n276 VSUBS 0.006967f
C603 B.n277 VSUBS 0.006967f
C604 B.n278 VSUBS 0.006967f
C605 B.n279 VSUBS 0.006967f
C606 B.n280 VSUBS 0.006967f
C607 B.n281 VSUBS 0.006967f
C608 B.n282 VSUBS 0.006967f
C609 B.n283 VSUBS 0.006967f
C610 B.n284 VSUBS 0.006967f
C611 B.n285 VSUBS 0.006967f
C612 B.n286 VSUBS 0.006967f
C613 B.n287 VSUBS 0.006967f
C614 B.n288 VSUBS 0.006967f
C615 B.n289 VSUBS 0.006967f
C616 B.n290 VSUBS 0.016827f
C617 B.n291 VSUBS 0.015549f
C618 B.n292 VSUBS 0.015549f
C619 B.n293 VSUBS 0.006967f
C620 B.n294 VSUBS 0.006967f
C621 B.n295 VSUBS 0.006967f
C622 B.n296 VSUBS 0.006967f
C623 B.n297 VSUBS 0.006967f
C624 B.n298 VSUBS 0.006967f
C625 B.n299 VSUBS 0.006967f
C626 B.n300 VSUBS 0.006967f
C627 B.n301 VSUBS 0.006967f
C628 B.n302 VSUBS 0.006967f
C629 B.n303 VSUBS 0.006967f
C630 B.n304 VSUBS 0.006967f
C631 B.n305 VSUBS 0.006967f
C632 B.n306 VSUBS 0.006967f
C633 B.n307 VSUBS 0.006967f
C634 B.n308 VSUBS 0.006967f
C635 B.n309 VSUBS 0.006967f
C636 B.n310 VSUBS 0.006967f
C637 B.n311 VSUBS 0.006967f
C638 B.n312 VSUBS 0.006967f
C639 B.n313 VSUBS 0.006967f
C640 B.n314 VSUBS 0.006967f
C641 B.n315 VSUBS 0.006967f
C642 B.n316 VSUBS 0.006967f
C643 B.n317 VSUBS 0.006967f
C644 B.n318 VSUBS 0.006967f
C645 B.n319 VSUBS 0.006967f
C646 B.n320 VSUBS 0.006967f
C647 B.n321 VSUBS 0.006967f
C648 B.n322 VSUBS 0.006967f
C649 B.n323 VSUBS 0.006967f
C650 B.n324 VSUBS 0.006967f
C651 B.n325 VSUBS 0.006967f
C652 B.n326 VSUBS 0.006967f
C653 B.n327 VSUBS 0.006967f
C654 B.n328 VSUBS 0.006967f
C655 B.n329 VSUBS 0.006967f
C656 B.n330 VSUBS 0.006967f
C657 B.n331 VSUBS 0.006967f
C658 B.n332 VSUBS 0.006967f
C659 B.n333 VSUBS 0.006967f
C660 B.n334 VSUBS 0.006967f
C661 B.n335 VSUBS 0.006967f
C662 B.n336 VSUBS 0.006967f
C663 B.n337 VSUBS 0.006967f
C664 B.n338 VSUBS 0.006967f
C665 B.n339 VSUBS 0.006967f
C666 B.n340 VSUBS 0.006967f
C667 B.n341 VSUBS 0.006967f
C668 B.n342 VSUBS 0.006967f
C669 B.n343 VSUBS 0.006967f
C670 B.n344 VSUBS 0.006967f
C671 B.n345 VSUBS 0.006967f
C672 B.n346 VSUBS 0.006967f
C673 B.n347 VSUBS 0.006967f
C674 B.n348 VSUBS 0.006967f
C675 B.n349 VSUBS 0.006967f
C676 B.n350 VSUBS 0.006967f
C677 B.n351 VSUBS 0.006967f
C678 B.n352 VSUBS 0.006967f
C679 B.n353 VSUBS 0.006967f
C680 B.n354 VSUBS 0.006967f
C681 B.n355 VSUBS 0.006967f
C682 B.n356 VSUBS 0.006967f
C683 B.n357 VSUBS 0.006967f
C684 B.n358 VSUBS 0.006967f
C685 B.n359 VSUBS 0.006967f
C686 B.n360 VSUBS 0.006967f
C687 B.n361 VSUBS 0.006967f
C688 B.n362 VSUBS 0.006967f
C689 B.n363 VSUBS 0.006967f
C690 B.n364 VSUBS 0.006967f
C691 B.n365 VSUBS 0.006967f
C692 B.n366 VSUBS 0.006967f
C693 B.n367 VSUBS 0.006967f
C694 B.n368 VSUBS 0.006967f
C695 B.n369 VSUBS 0.006967f
C696 B.n370 VSUBS 0.006967f
C697 B.n371 VSUBS 0.006967f
C698 B.n372 VSUBS 0.006967f
C699 B.n373 VSUBS 0.006967f
C700 B.n374 VSUBS 0.006967f
C701 B.n375 VSUBS 0.006967f
C702 B.n376 VSUBS 0.006967f
C703 B.n377 VSUBS 0.006967f
C704 B.n378 VSUBS 0.006967f
C705 B.n379 VSUBS 0.006967f
C706 B.n380 VSUBS 0.006967f
C707 B.n381 VSUBS 0.006967f
C708 B.n382 VSUBS 0.006967f
C709 B.n383 VSUBS 0.006967f
C710 B.n384 VSUBS 0.006967f
C711 B.n385 VSUBS 0.006967f
C712 B.n386 VSUBS 0.006967f
C713 B.n387 VSUBS 0.006967f
C714 B.n388 VSUBS 0.006967f
C715 B.n389 VSUBS 0.006967f
C716 B.n390 VSUBS 0.006967f
C717 B.n391 VSUBS 0.006967f
C718 B.n392 VSUBS 0.006967f
C719 B.n393 VSUBS 0.006967f
C720 B.n394 VSUBS 0.006967f
C721 B.n395 VSUBS 0.006967f
C722 B.n396 VSUBS 0.006967f
C723 B.n397 VSUBS 0.006967f
C724 B.n398 VSUBS 0.006967f
C725 B.n399 VSUBS 0.006967f
C726 B.n400 VSUBS 0.006967f
C727 B.n401 VSUBS 0.006967f
C728 B.n402 VSUBS 0.006967f
C729 B.n403 VSUBS 0.006967f
C730 B.n404 VSUBS 0.006967f
C731 B.n405 VSUBS 0.006967f
C732 B.n406 VSUBS 0.006967f
C733 B.n407 VSUBS 0.006967f
C734 B.n408 VSUBS 0.006967f
C735 B.n409 VSUBS 0.006967f
C736 B.n410 VSUBS 0.006967f
C737 B.n411 VSUBS 0.006967f
C738 B.n412 VSUBS 0.006967f
C739 B.n413 VSUBS 0.006967f
C740 B.n414 VSUBS 0.006967f
C741 B.n415 VSUBS 0.006967f
C742 B.n416 VSUBS 0.006967f
C743 B.n417 VSUBS 0.006967f
C744 B.n418 VSUBS 0.006967f
C745 B.n419 VSUBS 0.006967f
C746 B.n420 VSUBS 0.006967f
C747 B.n421 VSUBS 0.006967f
C748 B.n422 VSUBS 0.006967f
C749 B.n423 VSUBS 0.006967f
C750 B.n424 VSUBS 0.006967f
C751 B.n425 VSUBS 0.006967f
C752 B.n426 VSUBS 0.006967f
C753 B.n427 VSUBS 0.006967f
C754 B.n428 VSUBS 0.006967f
C755 B.n429 VSUBS 0.006967f
C756 B.n430 VSUBS 0.006967f
C757 B.n431 VSUBS 0.006967f
C758 B.n432 VSUBS 0.016381f
C759 B.n433 VSUBS 0.015549f
C760 B.n434 VSUBS 0.016827f
C761 B.n435 VSUBS 0.006967f
C762 B.n436 VSUBS 0.006967f
C763 B.n437 VSUBS 0.006967f
C764 B.n438 VSUBS 0.006967f
C765 B.n439 VSUBS 0.006967f
C766 B.n440 VSUBS 0.006967f
C767 B.n441 VSUBS 0.006967f
C768 B.n442 VSUBS 0.006967f
C769 B.n443 VSUBS 0.006967f
C770 B.n444 VSUBS 0.006967f
C771 B.n445 VSUBS 0.006967f
C772 B.n446 VSUBS 0.006967f
C773 B.n447 VSUBS 0.006967f
C774 B.n448 VSUBS 0.006967f
C775 B.n449 VSUBS 0.006967f
C776 B.n450 VSUBS 0.006967f
C777 B.n451 VSUBS 0.006967f
C778 B.n452 VSUBS 0.006967f
C779 B.n453 VSUBS 0.006967f
C780 B.n454 VSUBS 0.006967f
C781 B.n455 VSUBS 0.006967f
C782 B.n456 VSUBS 0.006967f
C783 B.n457 VSUBS 0.006967f
C784 B.n458 VSUBS 0.006967f
C785 B.n459 VSUBS 0.006967f
C786 B.n460 VSUBS 0.006557f
C787 B.n461 VSUBS 0.016142f
C788 B.n462 VSUBS 0.003893f
C789 B.n463 VSUBS 0.006967f
C790 B.n464 VSUBS 0.006967f
C791 B.n465 VSUBS 0.006967f
C792 B.n466 VSUBS 0.006967f
C793 B.n467 VSUBS 0.006967f
C794 B.n468 VSUBS 0.006967f
C795 B.n469 VSUBS 0.006967f
C796 B.n470 VSUBS 0.006967f
C797 B.n471 VSUBS 0.006967f
C798 B.n472 VSUBS 0.006967f
C799 B.n473 VSUBS 0.006967f
C800 B.n474 VSUBS 0.006967f
C801 B.n475 VSUBS 0.003893f
C802 B.n476 VSUBS 0.006967f
C803 B.n477 VSUBS 0.006967f
C804 B.n478 VSUBS 0.006967f
C805 B.n479 VSUBS 0.006967f
C806 B.n480 VSUBS 0.006967f
C807 B.n481 VSUBS 0.006967f
C808 B.n482 VSUBS 0.006967f
C809 B.n483 VSUBS 0.006967f
C810 B.n484 VSUBS 0.006967f
C811 B.n485 VSUBS 0.006967f
C812 B.n486 VSUBS 0.006967f
C813 B.n487 VSUBS 0.006967f
C814 B.n488 VSUBS 0.006967f
C815 B.n489 VSUBS 0.006967f
C816 B.n490 VSUBS 0.006967f
C817 B.n491 VSUBS 0.006967f
C818 B.n492 VSUBS 0.006967f
C819 B.n493 VSUBS 0.006967f
C820 B.n494 VSUBS 0.006967f
C821 B.n495 VSUBS 0.006967f
C822 B.n496 VSUBS 0.006967f
C823 B.n497 VSUBS 0.006967f
C824 B.n498 VSUBS 0.006967f
C825 B.n499 VSUBS 0.006967f
C826 B.n500 VSUBS 0.006967f
C827 B.n501 VSUBS 0.006967f
C828 B.n502 VSUBS 0.016827f
C829 B.n503 VSUBS 0.016827f
C830 B.n504 VSUBS 0.015549f
C831 B.n505 VSUBS 0.006967f
C832 B.n506 VSUBS 0.006967f
C833 B.n507 VSUBS 0.006967f
C834 B.n508 VSUBS 0.006967f
C835 B.n509 VSUBS 0.006967f
C836 B.n510 VSUBS 0.006967f
C837 B.n511 VSUBS 0.006967f
C838 B.n512 VSUBS 0.006967f
C839 B.n513 VSUBS 0.006967f
C840 B.n514 VSUBS 0.006967f
C841 B.n515 VSUBS 0.006967f
C842 B.n516 VSUBS 0.006967f
C843 B.n517 VSUBS 0.006967f
C844 B.n518 VSUBS 0.006967f
C845 B.n519 VSUBS 0.006967f
C846 B.n520 VSUBS 0.006967f
C847 B.n521 VSUBS 0.006967f
C848 B.n522 VSUBS 0.006967f
C849 B.n523 VSUBS 0.006967f
C850 B.n524 VSUBS 0.006967f
C851 B.n525 VSUBS 0.006967f
C852 B.n526 VSUBS 0.006967f
C853 B.n527 VSUBS 0.006967f
C854 B.n528 VSUBS 0.006967f
C855 B.n529 VSUBS 0.006967f
C856 B.n530 VSUBS 0.006967f
C857 B.n531 VSUBS 0.006967f
C858 B.n532 VSUBS 0.006967f
C859 B.n533 VSUBS 0.006967f
C860 B.n534 VSUBS 0.006967f
C861 B.n535 VSUBS 0.006967f
C862 B.n536 VSUBS 0.006967f
C863 B.n537 VSUBS 0.006967f
C864 B.n538 VSUBS 0.006967f
C865 B.n539 VSUBS 0.006967f
C866 B.n540 VSUBS 0.006967f
C867 B.n541 VSUBS 0.006967f
C868 B.n542 VSUBS 0.006967f
C869 B.n543 VSUBS 0.006967f
C870 B.n544 VSUBS 0.006967f
C871 B.n545 VSUBS 0.006967f
C872 B.n546 VSUBS 0.006967f
C873 B.n547 VSUBS 0.006967f
C874 B.n548 VSUBS 0.006967f
C875 B.n549 VSUBS 0.006967f
C876 B.n550 VSUBS 0.006967f
C877 B.n551 VSUBS 0.006967f
C878 B.n552 VSUBS 0.006967f
C879 B.n553 VSUBS 0.006967f
C880 B.n554 VSUBS 0.006967f
C881 B.n555 VSUBS 0.006967f
C882 B.n556 VSUBS 0.006967f
C883 B.n557 VSUBS 0.006967f
C884 B.n558 VSUBS 0.006967f
C885 B.n559 VSUBS 0.006967f
C886 B.n560 VSUBS 0.006967f
C887 B.n561 VSUBS 0.006967f
C888 B.n562 VSUBS 0.006967f
C889 B.n563 VSUBS 0.006967f
C890 B.n564 VSUBS 0.006967f
C891 B.n565 VSUBS 0.006967f
C892 B.n566 VSUBS 0.006967f
C893 B.n567 VSUBS 0.006967f
C894 B.n568 VSUBS 0.006967f
C895 B.n569 VSUBS 0.006967f
C896 B.n570 VSUBS 0.006967f
C897 B.n571 VSUBS 0.006967f
C898 B.n572 VSUBS 0.006967f
C899 B.n573 VSUBS 0.006967f
C900 B.n574 VSUBS 0.006967f
C901 B.n575 VSUBS 0.015775f
.ends

