* NGSPICE file created from opamp_sample_0013.ext - technology: sky130A

.subckt opamp_sample_0013 GND VOUT VDD VN VP CS_BIAS DIFFPAIR_BIAS
X0 VOUT.t44 GND.t128 VDD.t165 VDD.t86 sky130_fd_pr__pfet_01v8 ad=0.6138 pd=4.05 as=1.4508 ps=8.22 w=3.72 l=2.01
X1 GND.t123 GND.t121 GND.t122 GND.t73 sky130_fd_pr__nfet_01v8 ad=1.0101 pd=5.96 as=0 ps=0 w=2.59 l=4.93
X2 VOUT.t43 GND.t129 VDD.t164 VDD.t82 sky130_fd_pr__pfet_01v8 ad=1.4508 pd=8.22 as=0.6138 ps=4.05 w=3.72 l=2.01
X3 VOUT.t47 CS_BIAS.t8 GND.t127 GND.t29 sky130_fd_pr__nfet_01v8 ad=0.42735 pd=2.92 as=1.0101 ps=5.96 w=2.59 l=4.93
X4 CS_BIAS.t7 CS_BIAS.t6 GND.t31 GND.t29 sky130_fd_pr__nfet_01v8 ad=0.42735 pd=2.92 as=1.0101 ps=5.96 w=2.59 l=4.93
X5 VDD.t163 GND.t130 a_n2040_7754.t8 VDD.t162 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=1.95 ps=10.78 w=5 l=2.71
X6 VOUT.t42 GND.t131 VDD.t161 VDD.t130 sky130_fd_pr__pfet_01v8 ad=0.6138 pd=4.05 as=0.6138 ps=4.05 w=3.72 l=2.01
X7 GND.t120 GND.t118 GND.t119 GND.t37 sky130_fd_pr__nfet_01v8 ad=1.0101 pd=5.96 as=0 ps=0 w=2.59 l=4.93
X8 VDD.t80 VDD.t78 VDD.t79 VDD.t25 sky130_fd_pr__pfet_01v8 ad=1.4508 pd=8.22 as=0 ps=0 w=3.72 l=2.01
X9 VDD.t160 GND.t132 a_n5586_9514.t7 VDD.t159 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=1.95 ps=10.78 w=5 l=2.71
X10 a_n1816_n673.t10 VP.t3 GND.t15 GND.t14 sky130_fd_pr__nfet_01v8 ad=1.06755 pd=6.8 as=1.06755 ps=6.8 w=6.47 l=2.44
X11 VDD.t77 VDD.t75 VDD.t76 VDD.t69 sky130_fd_pr__pfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=2.71
X12 VDD.t74 VDD.t72 VDD.t73 VDD.t25 sky130_fd_pr__pfet_01v8 ad=1.4508 pd=8.22 as=0 ps=0 w=3.72 l=2.01
X13 VOUT.t41 GND.t133 VDD.t158 VDD.t108 sky130_fd_pr__pfet_01v8 ad=0.6138 pd=4.05 as=1.4508 ps=8.22 w=3.72 l=2.01
X14 VDD.t71 VDD.t68 VDD.t70 VDD.t69 sky130_fd_pr__pfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=2.71
X15 VDD.t67 VDD.t65 VDD.t66 VDD.t21 sky130_fd_pr__pfet_01v8 ad=1.4508 pd=8.22 as=0 ps=0 w=3.72 l=2.01
X16 GND.t117 GND.t115 GND.t116 GND.t61 sky130_fd_pr__nfet_01v8 ad=2.5233 pd=13.72 as=0 ps=0 w=6.47 l=2.44
X17 VOUT.t40 GND.t134 VDD.t157 VDD.t108 sky130_fd_pr__pfet_01v8 ad=0.6138 pd=4.05 as=1.4508 ps=8.22 w=3.72 l=2.01
X18 VDD.t156 GND.t135 VOUT.t39 VDD.t100 sky130_fd_pr__pfet_01v8 ad=0.6138 pd=4.05 as=0.6138 ps=4.05 w=3.72 l=2.01
X19 VOUT.t38 GND.t136 VDD.t155 VDD.t130 sky130_fd_pr__pfet_01v8 ad=0.6138 pd=4.05 as=0.6138 ps=4.05 w=3.72 l=2.01
X20 VOUT.t1 CS_BIAS.t9 GND.t18 GND.t10 sky130_fd_pr__nfet_01v8 ad=0.42735 pd=2.92 as=1.0101 ps=5.96 w=2.59 l=4.93
X21 VOUT.t48 a_n2040_7754.t0 sky130_fd_pr__cap_mim_m3_1 l=8.2 w=5.36
X22 VOUT.t0 CS_BIAS.t10 GND.t11 GND.t10 sky130_fd_pr__nfet_01v8 ad=0.42735 pd=2.92 as=1.0101 ps=5.96 w=2.59 l=4.93
X23 GND.t114 GND.t113 a_n2040_7754.t10 VDD.t121 sky130_fd_pr__pfet_01v8 ad=1.95 pd=10.78 as=1.95 ps=10.78 w=5 l=2.71
X24 VDD.t154 GND.t137 VOUT.t37 VDD.t100 sky130_fd_pr__pfet_01v8 ad=0.6138 pd=4.05 as=0.6138 ps=4.05 w=3.72 l=2.01
X25 VDD.t64 VDD.t62 VDD.t63 VDD.t17 sky130_fd_pr__pfet_01v8 ad=1.4508 pd=8.22 as=0 ps=0 w=3.72 l=2.01
X26 GND.t109 GND.t108 a_n2040_7754.t9 VDD.t102 sky130_fd_pr__pfet_01v8 ad=1.95 pd=10.78 as=1.95 ps=10.78 w=5 l=2.71
X27 VDD.t153 GND.t138 a_n5586_9514.t6 VDD.t152 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=2.71
X28 GND.t112 GND.t110 GND.t111 GND.t96 sky130_fd_pr__nfet_01v8 ad=1.0101 pd=5.96 as=0 ps=0 w=2.59 l=4.93
X29 GND.t107 GND.t105 GND.t106 GND.t96 sky130_fd_pr__nfet_01v8 ad=1.0101 pd=5.96 as=0 ps=0 w=2.59 l=4.93
X30 GND.t104 GND.t102 VN.t2 GND.t103 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X31 DIFFPAIR_BIAS.t1 DIFFPAIR_BIAS.t0 a_n1945_n3383.t2 GND.t4 sky130_fd_pr__nfet_01v8 ad=2.3088 pd=12.62 as=2.3088 ps=12.62 w=5.92 l=2.02
X32 VP.t2 GND.t99 GND.t101 GND.t100 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X33 GND.t98 GND.t95 GND.t97 GND.t96 sky130_fd_pr__nfet_01v8 ad=1.0101 pd=5.96 as=0 ps=0 w=2.59 l=4.93
X34 VDD.t151 GND.t139 VOUT.t36 VDD.t90 sky130_fd_pr__pfet_01v8 ad=0.6138 pd=4.05 as=0.6138 ps=4.05 w=3.72 l=2.01
X35 VDD.t150 GND.t140 VOUT.t35 VDD.t94 sky130_fd_pr__pfet_01v8 ad=0.6138 pd=4.05 as=0.6138 ps=4.05 w=3.72 l=2.01
X36 VOUT.t34 GND.t141 VDD.t149 VDD.t82 sky130_fd_pr__pfet_01v8 ad=1.4508 pd=8.22 as=0.6138 ps=4.05 w=3.72 l=2.01
X37 GND.t13 VN.t3 a_n1816_n673.t1 GND.t12 sky130_fd_pr__nfet_01v8 ad=2.5233 pd=13.72 as=1.06755 ps=6.8 w=6.47 l=2.44
X38 VDD.t61 VDD.t59 VDD.t60 VDD.t10 sky130_fd_pr__pfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=2.71
X39 a_n5586_9514.t5 GND.t142 VDD.t148 VDD.t147 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=2.71
X40 GND.t94 GND.t92 GND.t93 GND.t55 sky130_fd_pr__nfet_01v8 ad=1.0101 pd=5.96 as=0 ps=0 w=2.59 l=4.93
X41 a_n6412_9514# a_n6412_9514# a_n6412_9514# VDD.t81 sky130_fd_pr__pfet_01v8 ad=1.95 pd=10.78 as=3.9 ps=21.56 w=5 l=2.71
X42 GND.t6 VP.t4 a_n1816_n673.t9 GND.t5 sky130_fd_pr__nfet_01v8 ad=2.5233 pd=13.72 as=1.06755 ps=6.8 w=6.47 l=2.44
X43 VDD.t58 VDD.t56 VDD.t57 VDD.t6 sky130_fd_pr__pfet_01v8 ad=1.4508 pd=8.22 as=0 ps=0 w=3.72 l=2.01
X44 VOUT.t33 GND.t143 VDD.t146 VDD.t82 sky130_fd_pr__pfet_01v8 ad=1.4508 pd=8.22 as=0.6138 ps=4.05 w=3.72 l=2.01
X45 VDD.t140 GND.t144 VOUT.t32 VDD.t90 sky130_fd_pr__pfet_01v8 ad=0.6138 pd=4.05 as=0.6138 ps=4.05 w=3.72 l=2.01
X46 GND.t91 GND.t89 GND.t90 GND.t77 sky130_fd_pr__nfet_01v8 ad=2.5233 pd=13.72 as=0 ps=0 w=6.47 l=2.44
X47 a_n5586_9514.t4 GND.t145 VDD.t145 VDD.t144 sky130_fd_pr__pfet_01v8 ad=1.95 pd=10.78 as=0.825 ps=5.33 w=5 l=2.71
X48 VOUT.t31 GND.t146 VDD.t143 VDD.t86 sky130_fd_pr__pfet_01v8 ad=0.6138 pd=4.05 as=1.4508 ps=8.22 w=3.72 l=2.01
X49 GND.t126 CS_BIAS.t11 VOUT.t46 GND.t20 sky130_fd_pr__nfet_01v8 ad=1.0101 pd=5.96 as=0.42735 ps=2.92 w=2.59 l=4.93
X50 GND.t24 CS_BIAS.t12 VOUT.t2 GND.t20 sky130_fd_pr__nfet_01v8 ad=1.0101 pd=5.96 as=0.42735 ps=2.92 w=2.59 l=4.93
X51 VOUT.t30 GND.t147 VDD.t142 VDD.t88 sky130_fd_pr__pfet_01v8 ad=0.6138 pd=4.05 as=0.6138 ps=4.05 w=3.72 l=2.01
X52 VOUT.t29 GND.t148 VDD.t141 VDD.t108 sky130_fd_pr__pfet_01v8 ad=0.6138 pd=4.05 as=1.4508 ps=8.22 w=3.72 l=2.01
X53 a_n2040_7754.t7 GND.t149 VDD.t139 VDD.t138 sky130_fd_pr__pfet_01v8 ad=1.95 pd=10.78 as=0.825 ps=5.33 w=5 l=2.71
X54 a_n5586_9514.t3 GND.t150 VDD.t137 VDD.t136 sky130_fd_pr__pfet_01v8 ad=1.95 pd=10.78 as=0.825 ps=5.33 w=5 l=2.71
X55 CS_BIAS.t5 CS_BIAS.t4 GND.t27 GND.t10 sky130_fd_pr__nfet_01v8 ad=0.42735 pd=2.92 as=1.0101 ps=5.96 w=2.59 l=4.93
X56 GND.t88 GND.t86 VN.t1 GND.t87 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X57 VOUT.t28 GND.t151 VDD.t135 VDD.t130 sky130_fd_pr__pfet_01v8 ad=0.6138 pd=4.05 as=0.6138 ps=4.05 w=3.72 l=2.01
X58 VOUT.t27 GND.t152 VDD.t134 VDD.t96 sky130_fd_pr__pfet_01v8 ad=1.4508 pd=8.22 as=0.6138 ps=4.05 w=3.72 l=2.01
X59 VDD.t55 VDD.t53 VDD.t54 VDD.t44 sky130_fd_pr__pfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=2.71
X60 VDD.t133 GND.t153 a_n2040_7754.t6 VDD.t132 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=1.95 ps=10.78 w=5 l=2.71
X61 VOUT.t26 GND.t154 VDD.t131 VDD.t130 sky130_fd_pr__pfet_01v8 ad=0.6138 pd=4.05 as=0.6138 ps=4.05 w=3.72 l=2.01
X62 VDD.t129 GND.t155 VOUT.t25 VDD.t98 sky130_fd_pr__pfet_01v8 ad=0.6138 pd=4.05 as=0.6138 ps=4.05 w=3.72 l=2.01
X63 GND.t85 GND.t83 GND.t84 GND.t37 sky130_fd_pr__nfet_01v8 ad=1.0101 pd=5.96 as=0 ps=0 w=2.59 l=4.93
X64 VDD.t52 VDD.t50 VDD.t51 VDD.t17 sky130_fd_pr__pfet_01v8 ad=1.4508 pd=8.22 as=0 ps=0 w=3.72 l=2.01
X65 VDD.t128 GND.t156 a_n5586_9514.t2 VDD.t127 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=2.71
X66 VDD.t49 VDD.t47 VDD.t48 VDD.t21 sky130_fd_pr__pfet_01v8 ad=1.4508 pd=8.22 as=0 ps=0 w=3.72 l=2.01
X67 GND.t25 VN.t4 a_n1816_n673.t4 GND.t0 sky130_fd_pr__nfet_01v8 ad=1.06755 pd=6.8 as=2.5233 ps=13.72 w=6.47 l=2.44
X68 VOUT.t24 GND.t157 VDD.t126 VDD.t96 sky130_fd_pr__pfet_01v8 ad=1.4508 pd=8.22 as=0.6138 ps=4.05 w=3.72 l=2.01
X69 VDD.t46 VDD.t43 VDD.t45 VDD.t44 sky130_fd_pr__pfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=2.71
X70 VDD.t42 VDD.t40 VDD.t41 VDD.t21 sky130_fd_pr__pfet_01v8 ad=1.4508 pd=8.22 as=0 ps=0 w=3.72 l=2.01
X71 GND.t21 CS_BIAS.t2 CS_BIAS.t3 GND.t20 sky130_fd_pr__nfet_01v8 ad=1.0101 pd=5.96 as=0.42735 ps=2.92 w=2.59 l=4.93
X72 a_n1816_n673.t3 DIFFPAIR_BIAS.t6 a_n1279_n3383.t2 GND.t19 sky130_fd_pr__nfet_01v8 ad=2.3088 pd=12.62 as=2.3088 ps=12.62 w=5.92 l=2.02
X73 a_n1816_n673.t11 DIFFPAIR_BIAS.t7 a_n1279_n3383.t1 GND.t32 sky130_fd_pr__nfet_01v8 ad=2.3088 pd=12.62 as=2.3088 ps=12.62 w=5.92 l=2.02
X74 VOUT.t49 a_n2040_7754.t0 sky130_fd_pr__cap_mim_m3_1 l=8.2 w=5.36
X75 a_n1816_n673.t8 VP.t5 GND.t9 GND.t8 sky130_fd_pr__nfet_01v8 ad=1.06755 pd=6.8 as=1.06755 ps=6.8 w=6.47 l=2.44
X76 GND.t82 GND.t80 GND.t81 GND.t73 sky130_fd_pr__nfet_01v8 ad=1.0101 pd=5.96 as=0 ps=0 w=2.59 l=4.93
X77 VOUT.t23 GND.t158 VDD.t125 VDD.t88 sky130_fd_pr__pfet_01v8 ad=0.6138 pd=4.05 as=0.6138 ps=4.05 w=3.72 l=2.01
X78 GND.t28 VP.t6 a_n1816_n673.t7 GND.t16 sky130_fd_pr__nfet_01v8 ad=1.06755 pd=6.8 as=2.5233 ps=13.72 w=6.47 l=2.44
X79 VDD.t124 GND.t159 VOUT.t22 VDD.t98 sky130_fd_pr__pfet_01v8 ad=0.6138 pd=4.05 as=0.6138 ps=4.05 w=3.72 l=2.01
X80 VOUT.t50 a_n2040_7754.t0 sky130_fd_pr__cap_mim_m3_1 l=8.2 w=5.36
X81 VDD.t123 GND.t160 VOUT.t21 VDD.t94 sky130_fd_pr__pfet_01v8 ad=0.6138 pd=4.05 as=0.6138 ps=4.05 w=3.72 l=2.01
X82 VDD.t122 GND.t161 VOUT.t20 VDD.t90 sky130_fd_pr__pfet_01v8 ad=0.6138 pd=4.05 as=0.6138 ps=4.05 w=3.72 l=2.01
X83 GND.t26 CS_BIAS.t13 VOUT.t3 GND.t22 sky130_fd_pr__nfet_01v8 ad=1.0101 pd=5.96 as=0.42735 ps=2.92 w=2.59 l=4.93
X84 a_n5586_9514.t9 GND.t64 GND.t65 VDD.t121 sky130_fd_pr__pfet_01v8 ad=1.95 pd=10.78 as=1.95 ps=10.78 w=5 l=2.71
X85 VDD.t120 GND.t162 a_n2040_7754.t5 VDD.t119 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=2.71
X86 VDD.t118 GND.t163 a_n2040_7754.t4 VDD.t117 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=2.71
X87 VDD.t116 GND.t164 VOUT.t19 VDD.t94 sky130_fd_pr__pfet_01v8 ad=0.6138 pd=4.05 as=0.6138 ps=4.05 w=3.72 l=2.01
X88 VOUT.t18 GND.t165 VDD.t115 VDD.t88 sky130_fd_pr__pfet_01v8 ad=0.6138 pd=4.05 as=0.6138 ps=4.05 w=3.72 l=2.01
X89 VOUT.t17 GND.t166 VDD.t114 VDD.t86 sky130_fd_pr__pfet_01v8 ad=0.6138 pd=4.05 as=1.4508 ps=8.22 w=3.72 l=2.01
X90 VDD.t39 VDD.t37 VDD.t38 VDD.t25 sky130_fd_pr__pfet_01v8 ad=1.4508 pd=8.22 as=0 ps=0 w=3.72 l=2.01
X91 VDD.t36 VDD.t34 VDD.t35 VDD.t6 sky130_fd_pr__pfet_01v8 ad=1.4508 pd=8.22 as=0 ps=0 w=3.72 l=2.01
X92 GND.t79 GND.t76 GND.t78 GND.t77 sky130_fd_pr__nfet_01v8 ad=2.5233 pd=13.72 as=0 ps=0 w=6.47 l=2.44
X93 GND.t75 GND.t72 GND.t74 GND.t73 sky130_fd_pr__nfet_01v8 ad=1.0101 pd=5.96 as=0 ps=0 w=2.59 l=4.93
X94 VDD.t33 VDD.t31 VDD.t32 VDD.t6 sky130_fd_pr__pfet_01v8 ad=1.4508 pd=8.22 as=0 ps=0 w=3.72 l=2.01
X95 GND.t71 GND.t69 VP.t1 GND.t70 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X96 VOUT.t16 GND.t167 VDD.t113 VDD.t96 sky130_fd_pr__pfet_01v8 ad=1.4508 pd=8.22 as=0.6138 ps=4.05 w=3.72 l=2.01
X97 GND.t68 GND.t66 GND.t67 GND.t55 sky130_fd_pr__nfet_01v8 ad=1.0101 pd=5.96 as=0 ps=0 w=2.59 l=4.93
X98 VOUT.t51 a_n2040_7754.t0 sky130_fd_pr__cap_mim_m3_1 l=8.2 w=5.36
X99 VOUT.t52 a_n2040_7754.t0 sky130_fd_pr__cap_mim_m3_1 l=8.2 w=5.36
X100 a_n2040_7754.t3 GND.t168 VDD.t112 VDD.t111 sky130_fd_pr__pfet_01v8 ad=1.95 pd=10.78 as=0.825 ps=5.33 w=5 l=2.71
X101 DIFFPAIR_BIAS.t5 DIFFPAIR_BIAS.t4 a_n1945_n3383.t1 GND.t2 sky130_fd_pr__nfet_01v8 ad=2.3088 pd=12.62 as=2.3088 ps=12.62 w=5.92 l=2.02
X102 DIFFPAIR_BIAS.t3 DIFFPAIR_BIAS.t2 a_n1945_n3383.t0 GND.t3 sky130_fd_pr__nfet_01v8 ad=2.3088 pd=12.62 as=2.3088 ps=12.62 w=5.92 l=2.02
X103 a_n1816_n673.t13 VN.t5 GND.t35 GND.t14 sky130_fd_pr__nfet_01v8 ad=1.06755 pd=6.8 as=1.06755 ps=6.8 w=6.47 l=2.44
X104 VDD.t30 VDD.t28 VDD.t29 VDD.t17 sky130_fd_pr__pfet_01v8 ad=1.4508 pd=8.22 as=0 ps=0 w=3.72 l=2.01
X105 VOUT.t15 GND.t169 VDD.t109 VDD.t108 sky130_fd_pr__pfet_01v8 ad=0.6138 pd=4.05 as=1.4508 ps=8.22 w=3.72 l=2.01
X106 GND.t63 GND.t60 GND.t62 GND.t61 sky130_fd_pr__nfet_01v8 ad=2.5233 pd=13.72 as=0 ps=0 w=6.47 l=2.44
X107 VDD.t110 GND.t170 VOUT.t14 VDD.t100 sky130_fd_pr__pfet_01v8 ad=0.6138 pd=4.05 as=0.6138 ps=4.05 w=3.72 l=2.01
X108 VDD.t107 GND.t171 VOUT.t13 VDD.t98 sky130_fd_pr__pfet_01v8 ad=0.6138 pd=4.05 as=0.6138 ps=4.05 w=3.72 l=2.01
X109 VDD.t27 VDD.t24 VDD.t26 VDD.t25 sky130_fd_pr__pfet_01v8 ad=1.4508 pd=8.22 as=0 ps=0 w=3.72 l=2.01
X110 VDD.t106 GND.t172 a_n5586_9514.t1 VDD.t105 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=1.95 ps=10.78 w=5 l=2.71
X111 a_n2040_7754.t2 GND.t173 VDD.t104 VDD.t103 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=2.71
X112 GND.t124 CS_BIAS.t14 VOUT.t45 GND.t22 sky130_fd_pr__nfet_01v8 ad=1.0101 pd=5.96 as=0.42735 ps=2.92 w=2.59 l=4.93
X113 GND.t1 VP.t7 a_n1816_n673.t6 GND.t0 sky130_fd_pr__nfet_01v8 ad=1.06755 pd=6.8 as=2.5233 ps=13.72 w=6.47 l=2.44
X114 VDD.t23 VDD.t20 VDD.t22 VDD.t21 sky130_fd_pr__pfet_01v8 ad=1.4508 pd=8.22 as=0 ps=0 w=3.72 l=2.01
X115 VDD.t19 VDD.t16 VDD.t18 VDD.t17 sky130_fd_pr__pfet_01v8 ad=1.4508 pd=8.22 as=0 ps=0 w=3.72 l=2.01
X116 GND.t57 GND.t54 GND.t56 GND.t55 sky130_fd_pr__nfet_01v8 ad=1.0101 pd=5.96 as=0 ps=0 w=2.59 l=4.93
X117 a_n5586_9514.t8 GND.t58 GND.t59 VDD.t102 sky130_fd_pr__pfet_01v8 ad=1.95 pd=10.78 as=1.95 ps=10.78 w=5 l=2.71
X118 GND.t53 GND.t50 GND.t52 GND.t51 sky130_fd_pr__nfet_01v8 ad=2.3088 pd=12.62 as=0 ps=0 w=5.92 l=2.02
X119 VN.t0 GND.t47 GND.t49 GND.t48 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X120 a_n1816_n673.t0 DIFFPAIR_BIAS.t8 a_n1279_n3383.t0 GND.t7 sky130_fd_pr__nfet_01v8 ad=2.3088 pd=12.62 as=2.3088 ps=12.62 w=5.92 l=2.02
X121 GND.t46 GND.t44 VP.t0 GND.t45 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X122 VDD.t101 GND.t174 VOUT.t12 VDD.t100 sky130_fd_pr__pfet_01v8 ad=0.6138 pd=4.05 as=0.6138 ps=4.05 w=3.72 l=2.01
X123 VDD.t99 GND.t175 VOUT.t11 VDD.t98 sky130_fd_pr__pfet_01v8 ad=0.6138 pd=4.05 as=0.6138 ps=4.05 w=3.72 l=2.01
X124 VOUT.t4 CS_BIAS.t15 GND.t30 GND.t29 sky130_fd_pr__nfet_01v8 ad=0.42735 pd=2.92 as=1.0101 ps=5.96 w=2.59 l=4.93
X125 VOUT.t10 GND.t176 VDD.t97 VDD.t96 sky130_fd_pr__pfet_01v8 ad=1.4508 pd=8.22 as=0.6138 ps=4.05 w=3.72 l=2.01
X126 VDD.t95 GND.t177 VOUT.t9 VDD.t94 sky130_fd_pr__pfet_01v8 ad=0.6138 pd=4.05 as=0.6138 ps=4.05 w=3.72 l=2.01
X127 VDD.t15 VDD.t13 VDD.t14 VDD.t2 sky130_fd_pr__pfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=2.71
X128 a_n1816_n673.t14 VN.t6 GND.t125 GND.t8 sky130_fd_pr__nfet_01v8 ad=1.06755 pd=6.8 as=1.06755 ps=6.8 w=6.47 l=2.44
X129 a_n2040_7754.t1 GND.t178 VDD.t93 VDD.t92 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=2.71
X130 GND.t23 CS_BIAS.t0 CS_BIAS.t1 GND.t22 sky130_fd_pr__nfet_01v8 ad=1.0101 pd=5.96 as=0.42735 ps=2.92 w=2.59 l=4.93
X131 GND.t17 VN.t7 a_n1816_n673.t2 GND.t16 sky130_fd_pr__nfet_01v8 ad=1.06755 pd=6.8 as=2.5233 ps=13.72 w=6.47 l=2.44
X132 a_5714_9514# a_5714_9514# a_5714_9514# VDD.t0 sky130_fd_pr__pfet_01v8 ad=1.95 pd=10.78 as=3.9 ps=21.56 w=5 l=2.71
X133 VDD.t91 GND.t179 VOUT.t8 VDD.t90 sky130_fd_pr__pfet_01v8 ad=0.6138 pd=4.05 as=0.6138 ps=4.05 w=3.72 l=2.01
X134 VOUT.t7 GND.t180 VDD.t89 VDD.t88 sky130_fd_pr__pfet_01v8 ad=0.6138 pd=4.05 as=0.6138 ps=4.05 w=3.72 l=2.01
X135 VDD.t12 VDD.t9 VDD.t11 VDD.t10 sky130_fd_pr__pfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=2.71
X136 GND.t43 GND.t40 GND.t42 GND.t41 sky130_fd_pr__nfet_01v8 ad=2.3088 pd=12.62 as=0 ps=0 w=5.92 l=2.02
X137 GND.t39 GND.t36 GND.t38 GND.t37 sky130_fd_pr__nfet_01v8 ad=1.0101 pd=5.96 as=0 ps=0 w=2.59 l=4.93
X138 VOUT.t6 GND.t181 VDD.t87 VDD.t86 sky130_fd_pr__pfet_01v8 ad=0.6138 pd=4.05 as=1.4508 ps=8.22 w=3.72 l=2.01
X139 a_n5586_9514.t0 GND.t182 VDD.t85 VDD.t84 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=2.71
X140 VOUT.t5 GND.t183 VDD.t83 VDD.t82 sky130_fd_pr__pfet_01v8 ad=1.4508 pd=8.22 as=0.6138 ps=4.05 w=3.72 l=2.01
X141 GND.t33 VP.t8 a_n1816_n673.t5 GND.t12 sky130_fd_pr__nfet_01v8 ad=2.5233 pd=13.72 as=1.06755 ps=6.8 w=6.47 l=2.44
X142 VDD.t8 VDD.t5 VDD.t7 VDD.t6 sky130_fd_pr__pfet_01v8 ad=1.4508 pd=8.22 as=0 ps=0 w=3.72 l=2.01
X143 VDD.t4 VDD.t1 VDD.t3 VDD.t2 sky130_fd_pr__pfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=2.71
X144 VOUT.t53 a_n2040_7754.t0 sky130_fd_pr__cap_mim_m3_1 l=8.2 w=5.36
X145 GND.t34 VN.t8 a_n1816_n673.t12 GND.t5 sky130_fd_pr__nfet_01v8 ad=2.5233 pd=13.72 as=1.06755 ps=6.8 w=6.47 l=2.44
R0 GND.n5542 GND.n453 2347.19
R1 GND.n4866 GND.n904 924.168
R2 GND.n4973 GND.n799 826.439
R3 GND.n5543 GND.n454 826.439
R4 GND.n5685 GND.n374 826.439
R5 GND.n4859 GND.n905 826.439
R6 GND.n273 GND.n261 821.635
R7 GND.n4242 GND.n309 821.635
R8 GND.n4426 GND.n2381 821.635
R9 GND.n4388 GND.n2802 821.635
R10 GND.n4799 GND.n981 821.635
R11 GND.n4781 GND.n4780 821.635
R12 GND.n1206 GND.n1174 821.635
R13 GND.n4652 GND.n1171 821.635
R14 GND.n5791 GND.n266 807.22
R15 GND.n5749 GND.n308 807.22
R16 GND.n4391 GND.n4390 807.22
R17 GND.n4423 GND.n2398 807.22
R18 GND.n4699 GND.n1176 807.22
R19 GND.n4701 GND.n1169 807.22
R20 GND.n995 GND.n975 807.22
R21 GND.n4778 GND.n997 807.22
R22 GND.n4972 GND.n4971 804.557
R23 GND.n3880 GND.n2371 706.317
R24 GND.n3889 GND.n3091 706.317
R25 GND.n3281 GND.n3280 706.317
R26 GND.n3276 GND.n2073 706.317
R27 GND.n802 GND.n799 585
R28 GND.n4971 GND.n799 585
R29 GND.n4969 GND.n4968 585
R30 GND.n4970 GND.n4969 585
R31 GND.n4967 GND.n801 585
R32 GND.n801 GND.n800 585
R33 GND.n4966 GND.n4965 585
R34 GND.n4965 GND.n4964 585
R35 GND.n807 GND.n806 585
R36 GND.n4963 GND.n807 585
R37 GND.n4961 GND.n4960 585
R38 GND.n4962 GND.n4961 585
R39 GND.n4959 GND.n809 585
R40 GND.n809 GND.n808 585
R41 GND.n4958 GND.n4957 585
R42 GND.n4957 GND.n4956 585
R43 GND.n815 GND.n814 585
R44 GND.n4955 GND.n815 585
R45 GND.n4953 GND.n4952 585
R46 GND.n4954 GND.n4953 585
R47 GND.n4951 GND.n817 585
R48 GND.n817 GND.n816 585
R49 GND.n4950 GND.n4949 585
R50 GND.n4949 GND.n4948 585
R51 GND.n823 GND.n822 585
R52 GND.n4947 GND.n823 585
R53 GND.n4945 GND.n4944 585
R54 GND.n4946 GND.n4945 585
R55 GND.n4943 GND.n825 585
R56 GND.n825 GND.n824 585
R57 GND.n4942 GND.n4941 585
R58 GND.n4941 GND.n4940 585
R59 GND.n831 GND.n830 585
R60 GND.n4939 GND.n831 585
R61 GND.n4937 GND.n4936 585
R62 GND.n4938 GND.n4937 585
R63 GND.n4935 GND.n833 585
R64 GND.n833 GND.n832 585
R65 GND.n4934 GND.n4933 585
R66 GND.n4933 GND.n4932 585
R67 GND.n839 GND.n838 585
R68 GND.n4931 GND.n839 585
R69 GND.n4929 GND.n4928 585
R70 GND.n4930 GND.n4929 585
R71 GND.n4927 GND.n841 585
R72 GND.n841 GND.n840 585
R73 GND.n4926 GND.n4925 585
R74 GND.n4925 GND.n4924 585
R75 GND.n847 GND.n846 585
R76 GND.n4923 GND.n847 585
R77 GND.n4921 GND.n4920 585
R78 GND.n4922 GND.n4921 585
R79 GND.n4919 GND.n849 585
R80 GND.n849 GND.n848 585
R81 GND.n4918 GND.n4917 585
R82 GND.n4917 GND.n4916 585
R83 GND.n855 GND.n854 585
R84 GND.n4915 GND.n855 585
R85 GND.n4913 GND.n4912 585
R86 GND.n4914 GND.n4913 585
R87 GND.n4911 GND.n857 585
R88 GND.n857 GND.n856 585
R89 GND.n4910 GND.n4909 585
R90 GND.n4909 GND.n4908 585
R91 GND.n863 GND.n862 585
R92 GND.n4907 GND.n863 585
R93 GND.n4905 GND.n4904 585
R94 GND.n4906 GND.n4905 585
R95 GND.n4903 GND.n865 585
R96 GND.n865 GND.n864 585
R97 GND.n4902 GND.n4901 585
R98 GND.n4901 GND.n4900 585
R99 GND.n871 GND.n870 585
R100 GND.n4899 GND.n871 585
R101 GND.n4897 GND.n4896 585
R102 GND.n4898 GND.n4897 585
R103 GND.n4895 GND.n873 585
R104 GND.n873 GND.n872 585
R105 GND.n4894 GND.n4893 585
R106 GND.n4893 GND.n4892 585
R107 GND.n879 GND.n878 585
R108 GND.n4891 GND.n879 585
R109 GND.n4889 GND.n4888 585
R110 GND.n4890 GND.n4889 585
R111 GND.n4887 GND.n881 585
R112 GND.n881 GND.n880 585
R113 GND.n4886 GND.n4885 585
R114 GND.n4885 GND.n4884 585
R115 GND.n887 GND.n886 585
R116 GND.n4883 GND.n887 585
R117 GND.n4881 GND.n4880 585
R118 GND.n4882 GND.n4881 585
R119 GND.n4879 GND.n889 585
R120 GND.n889 GND.n888 585
R121 GND.n4878 GND.n4877 585
R122 GND.n4877 GND.n4876 585
R123 GND.n895 GND.n894 585
R124 GND.n4875 GND.n895 585
R125 GND.n4873 GND.n4872 585
R126 GND.n4874 GND.n4873 585
R127 GND.n4871 GND.n897 585
R128 GND.n897 GND.n896 585
R129 GND.n4870 GND.n4869 585
R130 GND.n4869 GND.n4868 585
R131 GND.n903 GND.n902 585
R132 GND.n4867 GND.n903 585
R133 GND.n4865 GND.n4864 585
R134 GND.n4866 GND.n4865 585
R135 GND.n4974 GND.n4973 585
R136 GND.n4973 GND.n4972 585
R137 GND.n797 GND.n796 585
R138 GND.n796 GND.n795 585
R139 GND.n4979 GND.n4978 585
R140 GND.n4980 GND.n4979 585
R141 GND.n794 GND.n793 585
R142 GND.n4981 GND.n794 585
R143 GND.n4984 GND.n4983 585
R144 GND.n4983 GND.n4982 585
R145 GND.n791 GND.n790 585
R146 GND.n790 GND.n789 585
R147 GND.n4989 GND.n4988 585
R148 GND.n4990 GND.n4989 585
R149 GND.n788 GND.n787 585
R150 GND.n4991 GND.n788 585
R151 GND.n4994 GND.n4993 585
R152 GND.n4993 GND.n4992 585
R153 GND.n785 GND.n784 585
R154 GND.n784 GND.n783 585
R155 GND.n4999 GND.n4998 585
R156 GND.n5000 GND.n4999 585
R157 GND.n782 GND.n781 585
R158 GND.n5001 GND.n782 585
R159 GND.n5004 GND.n5003 585
R160 GND.n5003 GND.n5002 585
R161 GND.n779 GND.n778 585
R162 GND.n778 GND.n777 585
R163 GND.n5009 GND.n5008 585
R164 GND.n5010 GND.n5009 585
R165 GND.n776 GND.n775 585
R166 GND.n5011 GND.n776 585
R167 GND.n5014 GND.n5013 585
R168 GND.n5013 GND.n5012 585
R169 GND.n773 GND.n772 585
R170 GND.n772 GND.n771 585
R171 GND.n5019 GND.n5018 585
R172 GND.n5020 GND.n5019 585
R173 GND.n770 GND.n769 585
R174 GND.n5021 GND.n770 585
R175 GND.n5024 GND.n5023 585
R176 GND.n5023 GND.n5022 585
R177 GND.n767 GND.n766 585
R178 GND.n766 GND.n765 585
R179 GND.n5029 GND.n5028 585
R180 GND.n5030 GND.n5029 585
R181 GND.n764 GND.n763 585
R182 GND.n5031 GND.n764 585
R183 GND.n5034 GND.n5033 585
R184 GND.n5033 GND.n5032 585
R185 GND.n761 GND.n760 585
R186 GND.n760 GND.n759 585
R187 GND.n5039 GND.n5038 585
R188 GND.n5040 GND.n5039 585
R189 GND.n758 GND.n757 585
R190 GND.n5041 GND.n758 585
R191 GND.n5044 GND.n5043 585
R192 GND.n5043 GND.n5042 585
R193 GND.n755 GND.n754 585
R194 GND.n754 GND.n753 585
R195 GND.n5049 GND.n5048 585
R196 GND.n5050 GND.n5049 585
R197 GND.n752 GND.n751 585
R198 GND.n5051 GND.n752 585
R199 GND.n5054 GND.n5053 585
R200 GND.n5053 GND.n5052 585
R201 GND.n749 GND.n748 585
R202 GND.n748 GND.n747 585
R203 GND.n5059 GND.n5058 585
R204 GND.n5060 GND.n5059 585
R205 GND.n746 GND.n745 585
R206 GND.n5061 GND.n746 585
R207 GND.n5064 GND.n5063 585
R208 GND.n5063 GND.n5062 585
R209 GND.n743 GND.n742 585
R210 GND.n742 GND.n741 585
R211 GND.n5069 GND.n5068 585
R212 GND.n5070 GND.n5069 585
R213 GND.n740 GND.n739 585
R214 GND.n5071 GND.n740 585
R215 GND.n5074 GND.n5073 585
R216 GND.n5073 GND.n5072 585
R217 GND.n737 GND.n736 585
R218 GND.n736 GND.n735 585
R219 GND.n5079 GND.n5078 585
R220 GND.n5080 GND.n5079 585
R221 GND.n734 GND.n733 585
R222 GND.n5081 GND.n734 585
R223 GND.n5084 GND.n5083 585
R224 GND.n5083 GND.n5082 585
R225 GND.n731 GND.n730 585
R226 GND.n730 GND.n729 585
R227 GND.n5089 GND.n5088 585
R228 GND.n5090 GND.n5089 585
R229 GND.n728 GND.n727 585
R230 GND.n5091 GND.n728 585
R231 GND.n5094 GND.n5093 585
R232 GND.n5093 GND.n5092 585
R233 GND.n725 GND.n724 585
R234 GND.n724 GND.n723 585
R235 GND.n5099 GND.n5098 585
R236 GND.n5100 GND.n5099 585
R237 GND.n722 GND.n721 585
R238 GND.n5101 GND.n722 585
R239 GND.n5104 GND.n5103 585
R240 GND.n5103 GND.n5102 585
R241 GND.n719 GND.n718 585
R242 GND.n718 GND.n717 585
R243 GND.n5109 GND.n5108 585
R244 GND.n5110 GND.n5109 585
R245 GND.n716 GND.n715 585
R246 GND.n5111 GND.n716 585
R247 GND.n5114 GND.n5113 585
R248 GND.n5113 GND.n5112 585
R249 GND.n713 GND.n712 585
R250 GND.n712 GND.n711 585
R251 GND.n5119 GND.n5118 585
R252 GND.n5120 GND.n5119 585
R253 GND.n710 GND.n709 585
R254 GND.n5121 GND.n710 585
R255 GND.n5124 GND.n5123 585
R256 GND.n5123 GND.n5122 585
R257 GND.n707 GND.n706 585
R258 GND.n706 GND.n705 585
R259 GND.n5129 GND.n5128 585
R260 GND.n5130 GND.n5129 585
R261 GND.n704 GND.n703 585
R262 GND.n5131 GND.n704 585
R263 GND.n5134 GND.n5133 585
R264 GND.n5133 GND.n5132 585
R265 GND.n701 GND.n700 585
R266 GND.n700 GND.n699 585
R267 GND.n5139 GND.n5138 585
R268 GND.n5140 GND.n5139 585
R269 GND.n698 GND.n697 585
R270 GND.n5141 GND.n698 585
R271 GND.n5144 GND.n5143 585
R272 GND.n5143 GND.n5142 585
R273 GND.n695 GND.n694 585
R274 GND.n694 GND.n693 585
R275 GND.n5149 GND.n5148 585
R276 GND.n5150 GND.n5149 585
R277 GND.n692 GND.n691 585
R278 GND.n5151 GND.n692 585
R279 GND.n5154 GND.n5153 585
R280 GND.n5153 GND.n5152 585
R281 GND.n689 GND.n688 585
R282 GND.n688 GND.n687 585
R283 GND.n5159 GND.n5158 585
R284 GND.n5160 GND.n5159 585
R285 GND.n686 GND.n685 585
R286 GND.n5161 GND.n686 585
R287 GND.n5164 GND.n5163 585
R288 GND.n5163 GND.n5162 585
R289 GND.n683 GND.n682 585
R290 GND.n682 GND.n681 585
R291 GND.n5169 GND.n5168 585
R292 GND.n5170 GND.n5169 585
R293 GND.n680 GND.n679 585
R294 GND.n5171 GND.n680 585
R295 GND.n5174 GND.n5173 585
R296 GND.n5173 GND.n5172 585
R297 GND.n677 GND.n676 585
R298 GND.n676 GND.n675 585
R299 GND.n5179 GND.n5178 585
R300 GND.n5180 GND.n5179 585
R301 GND.n674 GND.n673 585
R302 GND.n5181 GND.n674 585
R303 GND.n5184 GND.n5183 585
R304 GND.n5183 GND.n5182 585
R305 GND.n671 GND.n670 585
R306 GND.n670 GND.n669 585
R307 GND.n5189 GND.n5188 585
R308 GND.n5190 GND.n5189 585
R309 GND.n668 GND.n667 585
R310 GND.n5191 GND.n668 585
R311 GND.n5194 GND.n5193 585
R312 GND.n5193 GND.n5192 585
R313 GND.n665 GND.n664 585
R314 GND.n664 GND.n663 585
R315 GND.n5199 GND.n5198 585
R316 GND.n5200 GND.n5199 585
R317 GND.n662 GND.n661 585
R318 GND.n5201 GND.n662 585
R319 GND.n5204 GND.n5203 585
R320 GND.n5203 GND.n5202 585
R321 GND.n659 GND.n658 585
R322 GND.n658 GND.n657 585
R323 GND.n5209 GND.n5208 585
R324 GND.n5210 GND.n5209 585
R325 GND.n656 GND.n655 585
R326 GND.n5211 GND.n656 585
R327 GND.n5214 GND.n5213 585
R328 GND.n5213 GND.n5212 585
R329 GND.n653 GND.n652 585
R330 GND.n652 GND.n651 585
R331 GND.n5219 GND.n5218 585
R332 GND.n5220 GND.n5219 585
R333 GND.n650 GND.n649 585
R334 GND.n5221 GND.n650 585
R335 GND.n5224 GND.n5223 585
R336 GND.n5223 GND.n5222 585
R337 GND.n647 GND.n646 585
R338 GND.n646 GND.n645 585
R339 GND.n5229 GND.n5228 585
R340 GND.n5230 GND.n5229 585
R341 GND.n644 GND.n643 585
R342 GND.n5231 GND.n644 585
R343 GND.n5234 GND.n5233 585
R344 GND.n5233 GND.n5232 585
R345 GND.n641 GND.n640 585
R346 GND.n640 GND.n639 585
R347 GND.n5239 GND.n5238 585
R348 GND.n5240 GND.n5239 585
R349 GND.n638 GND.n637 585
R350 GND.n5241 GND.n638 585
R351 GND.n5244 GND.n5243 585
R352 GND.n5243 GND.n5242 585
R353 GND.n635 GND.n634 585
R354 GND.n634 GND.n633 585
R355 GND.n5249 GND.n5248 585
R356 GND.n5250 GND.n5249 585
R357 GND.n632 GND.n631 585
R358 GND.n5251 GND.n632 585
R359 GND.n5254 GND.n5253 585
R360 GND.n5253 GND.n5252 585
R361 GND.n629 GND.n628 585
R362 GND.n628 GND.n627 585
R363 GND.n5259 GND.n5258 585
R364 GND.n5260 GND.n5259 585
R365 GND.n626 GND.n625 585
R366 GND.n5261 GND.n626 585
R367 GND.n5264 GND.n5263 585
R368 GND.n5263 GND.n5262 585
R369 GND.n623 GND.n622 585
R370 GND.n622 GND.n621 585
R371 GND.n5269 GND.n5268 585
R372 GND.n5270 GND.n5269 585
R373 GND.n620 GND.n619 585
R374 GND.n5271 GND.n620 585
R375 GND.n5274 GND.n5273 585
R376 GND.n5273 GND.n5272 585
R377 GND.n617 GND.n616 585
R378 GND.n616 GND.n615 585
R379 GND.n5279 GND.n5278 585
R380 GND.n5280 GND.n5279 585
R381 GND.n614 GND.n613 585
R382 GND.n5281 GND.n614 585
R383 GND.n5284 GND.n5283 585
R384 GND.n5283 GND.n5282 585
R385 GND.n611 GND.n610 585
R386 GND.n610 GND.n609 585
R387 GND.n5289 GND.n5288 585
R388 GND.n5290 GND.n5289 585
R389 GND.n608 GND.n607 585
R390 GND.n5291 GND.n608 585
R391 GND.n5294 GND.n5293 585
R392 GND.n5293 GND.n5292 585
R393 GND.n605 GND.n604 585
R394 GND.n604 GND.n603 585
R395 GND.n5299 GND.n5298 585
R396 GND.n5300 GND.n5299 585
R397 GND.n602 GND.n601 585
R398 GND.n5301 GND.n602 585
R399 GND.n5304 GND.n5303 585
R400 GND.n5303 GND.n5302 585
R401 GND.n599 GND.n598 585
R402 GND.n598 GND.n597 585
R403 GND.n5309 GND.n5308 585
R404 GND.n5310 GND.n5309 585
R405 GND.n596 GND.n595 585
R406 GND.n5311 GND.n596 585
R407 GND.n5314 GND.n5313 585
R408 GND.n5313 GND.n5312 585
R409 GND.n593 GND.n592 585
R410 GND.n592 GND.n591 585
R411 GND.n5319 GND.n5318 585
R412 GND.n5320 GND.n5319 585
R413 GND.n590 GND.n589 585
R414 GND.n5321 GND.n590 585
R415 GND.n5324 GND.n5323 585
R416 GND.n5323 GND.n5322 585
R417 GND.n587 GND.n586 585
R418 GND.n586 GND.n585 585
R419 GND.n5329 GND.n5328 585
R420 GND.n5330 GND.n5329 585
R421 GND.n584 GND.n583 585
R422 GND.n5331 GND.n584 585
R423 GND.n5334 GND.n5333 585
R424 GND.n5333 GND.n5332 585
R425 GND.n581 GND.n580 585
R426 GND.n580 GND.n579 585
R427 GND.n5339 GND.n5338 585
R428 GND.n5340 GND.n5339 585
R429 GND.n578 GND.n577 585
R430 GND.n5341 GND.n578 585
R431 GND.n5344 GND.n5343 585
R432 GND.n5343 GND.n5342 585
R433 GND.n575 GND.n574 585
R434 GND.n574 GND.n573 585
R435 GND.n5349 GND.n5348 585
R436 GND.n5350 GND.n5349 585
R437 GND.n572 GND.n571 585
R438 GND.n5351 GND.n572 585
R439 GND.n5354 GND.n5353 585
R440 GND.n5353 GND.n5352 585
R441 GND.n569 GND.n568 585
R442 GND.n568 GND.n567 585
R443 GND.n5359 GND.n5358 585
R444 GND.n5360 GND.n5359 585
R445 GND.n566 GND.n565 585
R446 GND.n5361 GND.n566 585
R447 GND.n5364 GND.n5363 585
R448 GND.n5363 GND.n5362 585
R449 GND.n563 GND.n562 585
R450 GND.n562 GND.n561 585
R451 GND.n5369 GND.n5368 585
R452 GND.n5370 GND.n5369 585
R453 GND.n560 GND.n559 585
R454 GND.n5371 GND.n560 585
R455 GND.n5374 GND.n5373 585
R456 GND.n5373 GND.n5372 585
R457 GND.n557 GND.n556 585
R458 GND.n556 GND.n555 585
R459 GND.n5379 GND.n5378 585
R460 GND.n5380 GND.n5379 585
R461 GND.n554 GND.n553 585
R462 GND.n5381 GND.n554 585
R463 GND.n5384 GND.n5383 585
R464 GND.n5383 GND.n5382 585
R465 GND.n551 GND.n550 585
R466 GND.n550 GND.n549 585
R467 GND.n5389 GND.n5388 585
R468 GND.n5390 GND.n5389 585
R469 GND.n548 GND.n547 585
R470 GND.n5391 GND.n548 585
R471 GND.n5394 GND.n5393 585
R472 GND.n5393 GND.n5392 585
R473 GND.n545 GND.n544 585
R474 GND.n544 GND.n543 585
R475 GND.n5399 GND.n5398 585
R476 GND.n5400 GND.n5399 585
R477 GND.n542 GND.n541 585
R478 GND.n5401 GND.n542 585
R479 GND.n5404 GND.n5403 585
R480 GND.n5403 GND.n5402 585
R481 GND.n539 GND.n538 585
R482 GND.n538 GND.n537 585
R483 GND.n5409 GND.n5408 585
R484 GND.n5410 GND.n5409 585
R485 GND.n536 GND.n535 585
R486 GND.n5411 GND.n536 585
R487 GND.n5414 GND.n5413 585
R488 GND.n5413 GND.n5412 585
R489 GND.n533 GND.n532 585
R490 GND.n532 GND.n531 585
R491 GND.n5419 GND.n5418 585
R492 GND.n5420 GND.n5419 585
R493 GND.n530 GND.n529 585
R494 GND.n5421 GND.n530 585
R495 GND.n5424 GND.n5423 585
R496 GND.n5423 GND.n5422 585
R497 GND.n527 GND.n526 585
R498 GND.n526 GND.n525 585
R499 GND.n5429 GND.n5428 585
R500 GND.n5430 GND.n5429 585
R501 GND.n524 GND.n523 585
R502 GND.n5431 GND.n524 585
R503 GND.n5434 GND.n5433 585
R504 GND.n5433 GND.n5432 585
R505 GND.n521 GND.n520 585
R506 GND.n520 GND.n519 585
R507 GND.n5439 GND.n5438 585
R508 GND.n5440 GND.n5439 585
R509 GND.n518 GND.n517 585
R510 GND.n5441 GND.n518 585
R511 GND.n5444 GND.n5443 585
R512 GND.n5443 GND.n5442 585
R513 GND.n515 GND.n514 585
R514 GND.n514 GND.n513 585
R515 GND.n5449 GND.n5448 585
R516 GND.n5450 GND.n5449 585
R517 GND.n512 GND.n511 585
R518 GND.n5451 GND.n512 585
R519 GND.n5454 GND.n5453 585
R520 GND.n5453 GND.n5452 585
R521 GND.n509 GND.n508 585
R522 GND.n508 GND.n507 585
R523 GND.n5459 GND.n5458 585
R524 GND.n5460 GND.n5459 585
R525 GND.n506 GND.n505 585
R526 GND.n5461 GND.n506 585
R527 GND.n5464 GND.n5463 585
R528 GND.n5463 GND.n5462 585
R529 GND.n503 GND.n502 585
R530 GND.n502 GND.n501 585
R531 GND.n5469 GND.n5468 585
R532 GND.n5470 GND.n5469 585
R533 GND.n500 GND.n499 585
R534 GND.n5471 GND.n500 585
R535 GND.n5474 GND.n5473 585
R536 GND.n5473 GND.n5472 585
R537 GND.n497 GND.n496 585
R538 GND.n496 GND.n495 585
R539 GND.n5479 GND.n5478 585
R540 GND.n5480 GND.n5479 585
R541 GND.n494 GND.n493 585
R542 GND.n5481 GND.n494 585
R543 GND.n5484 GND.n5483 585
R544 GND.n5483 GND.n5482 585
R545 GND.n491 GND.n490 585
R546 GND.n490 GND.n489 585
R547 GND.n5489 GND.n5488 585
R548 GND.n5490 GND.n5489 585
R549 GND.n488 GND.n487 585
R550 GND.n5491 GND.n488 585
R551 GND.n5494 GND.n5493 585
R552 GND.n5493 GND.n5492 585
R553 GND.n485 GND.n484 585
R554 GND.n484 GND.n483 585
R555 GND.n5499 GND.n5498 585
R556 GND.n5500 GND.n5499 585
R557 GND.n482 GND.n481 585
R558 GND.n5501 GND.n482 585
R559 GND.n5504 GND.n5503 585
R560 GND.n5503 GND.n5502 585
R561 GND.n479 GND.n478 585
R562 GND.n478 GND.n477 585
R563 GND.n5509 GND.n5508 585
R564 GND.n5510 GND.n5509 585
R565 GND.n476 GND.n475 585
R566 GND.n5511 GND.n476 585
R567 GND.n5514 GND.n5513 585
R568 GND.n5513 GND.n5512 585
R569 GND.n473 GND.n472 585
R570 GND.n472 GND.n471 585
R571 GND.n5519 GND.n5518 585
R572 GND.n5520 GND.n5519 585
R573 GND.n470 GND.n469 585
R574 GND.n5521 GND.n470 585
R575 GND.n5524 GND.n5523 585
R576 GND.n5523 GND.n5522 585
R577 GND.n467 GND.n466 585
R578 GND.n466 GND.n465 585
R579 GND.n5529 GND.n5528 585
R580 GND.n5530 GND.n5529 585
R581 GND.n464 GND.n463 585
R582 GND.n5531 GND.n464 585
R583 GND.n5534 GND.n5533 585
R584 GND.n5533 GND.n5532 585
R585 GND.n461 GND.n460 585
R586 GND.n460 GND.n459 585
R587 GND.n5539 GND.n5538 585
R588 GND.n5540 GND.n5539 585
R589 GND.n458 GND.n457 585
R590 GND.n5541 GND.n458 585
R591 GND.n5544 GND.n5543 585
R592 GND.n5543 GND.n5542 585
R593 GND.n5681 GND.n5680 585
R594 GND.n5682 GND.n5681 585
R595 GND.n377 GND.n376 585
R596 GND.n376 GND.n375 585
R597 GND.n5674 GND.n5673 585
R598 GND.n5673 GND.n5672 585
R599 GND.n380 GND.n379 585
R600 GND.n5671 GND.n380 585
R601 GND.n5669 GND.n5668 585
R602 GND.n5670 GND.n5669 585
R603 GND.n383 GND.n382 585
R604 GND.n382 GND.n381 585
R605 GND.n5664 GND.n5663 585
R606 GND.n5663 GND.n5662 585
R607 GND.n386 GND.n385 585
R608 GND.n5661 GND.n386 585
R609 GND.n5659 GND.n5658 585
R610 GND.n5660 GND.n5659 585
R611 GND.n389 GND.n388 585
R612 GND.n388 GND.n387 585
R613 GND.n5654 GND.n5653 585
R614 GND.n5653 GND.n5652 585
R615 GND.n392 GND.n391 585
R616 GND.n5651 GND.n392 585
R617 GND.n5649 GND.n5648 585
R618 GND.n5650 GND.n5649 585
R619 GND.n395 GND.n394 585
R620 GND.n394 GND.n393 585
R621 GND.n5644 GND.n5643 585
R622 GND.n5643 GND.n5642 585
R623 GND.n398 GND.n397 585
R624 GND.n5641 GND.n398 585
R625 GND.n5639 GND.n5638 585
R626 GND.n5640 GND.n5639 585
R627 GND.n401 GND.n400 585
R628 GND.n400 GND.n399 585
R629 GND.n5634 GND.n5633 585
R630 GND.n5633 GND.n5632 585
R631 GND.n404 GND.n403 585
R632 GND.n5631 GND.n404 585
R633 GND.n5629 GND.n5628 585
R634 GND.n5630 GND.n5629 585
R635 GND.n407 GND.n406 585
R636 GND.n406 GND.n405 585
R637 GND.n5624 GND.n5623 585
R638 GND.n5623 GND.n5622 585
R639 GND.n410 GND.n409 585
R640 GND.n5621 GND.n410 585
R641 GND.n5619 GND.n5618 585
R642 GND.n5620 GND.n5619 585
R643 GND.n413 GND.n412 585
R644 GND.n412 GND.n411 585
R645 GND.n5614 GND.n5613 585
R646 GND.n5613 GND.n5612 585
R647 GND.n416 GND.n415 585
R648 GND.n5611 GND.n416 585
R649 GND.n5609 GND.n5608 585
R650 GND.n5610 GND.n5609 585
R651 GND.n419 GND.n418 585
R652 GND.n418 GND.n417 585
R653 GND.n5604 GND.n5603 585
R654 GND.n5603 GND.n5602 585
R655 GND.n422 GND.n421 585
R656 GND.n5601 GND.n422 585
R657 GND.n5599 GND.n5598 585
R658 GND.n5600 GND.n5599 585
R659 GND.n425 GND.n424 585
R660 GND.n424 GND.n423 585
R661 GND.n5594 GND.n5593 585
R662 GND.n5593 GND.n5592 585
R663 GND.n428 GND.n427 585
R664 GND.n5591 GND.n428 585
R665 GND.n5589 GND.n5588 585
R666 GND.n5590 GND.n5589 585
R667 GND.n431 GND.n430 585
R668 GND.n430 GND.n429 585
R669 GND.n5584 GND.n5583 585
R670 GND.n5583 GND.n5582 585
R671 GND.n434 GND.n433 585
R672 GND.n5581 GND.n434 585
R673 GND.n5579 GND.n5578 585
R674 GND.n5580 GND.n5579 585
R675 GND.n437 GND.n436 585
R676 GND.n436 GND.n435 585
R677 GND.n5574 GND.n5573 585
R678 GND.n5573 GND.n5572 585
R679 GND.n440 GND.n439 585
R680 GND.n5571 GND.n440 585
R681 GND.n5569 GND.n5568 585
R682 GND.n5570 GND.n5569 585
R683 GND.n443 GND.n442 585
R684 GND.n442 GND.n441 585
R685 GND.n5564 GND.n5563 585
R686 GND.n5563 GND.n5562 585
R687 GND.n446 GND.n445 585
R688 GND.n5561 GND.n446 585
R689 GND.n5559 GND.n5558 585
R690 GND.n5560 GND.n5559 585
R691 GND.n449 GND.n448 585
R692 GND.n448 GND.n447 585
R693 GND.n5554 GND.n5553 585
R694 GND.n5553 GND.n5552 585
R695 GND.n452 GND.n451 585
R696 GND.n5551 GND.n452 585
R697 GND.n5549 GND.n5548 585
R698 GND.n5550 GND.n5549 585
R699 GND.n455 GND.n454 585
R700 GND.n454 GND.n453 585
R701 GND.n4431 GND.n2371 585
R702 GND.n3890 GND.n2371 585
R703 GND.n4433 GND.n4432 585
R704 GND.n4434 GND.n4433 585
R705 GND.n2372 GND.n2370 585
R706 GND.n2370 GND.n2361 585
R707 GND.n3798 GND.n3797 585
R708 GND.n3799 GND.n3798 585
R709 GND.n2343 GND.n2342 585
R710 GND.n3772 GND.n2343 585
R711 GND.n4450 GND.n4449 585
R712 GND.n4449 GND.n4448 585
R713 GND.n4451 GND.n2329 585
R714 GND.n3768 GND.n2329 585
R715 GND.n4453 GND.n4452 585
R716 GND.n4454 GND.n4453 585
R717 GND.n2330 GND.n2328 585
R718 GND.n2328 GND.n2318 585
R719 GND.n2336 GND.n2335 585
R720 GND.n2335 GND.n2316 585
R721 GND.n2334 GND.n2333 585
R722 GND.n2334 GND.n2302 585
R723 GND.n2291 GND.n2290 585
R724 GND.n2300 GND.n2291 585
R725 GND.n4478 GND.n4477 585
R726 GND.n4477 GND.n4476 585
R727 GND.n4479 GND.n2280 585
R728 GND.n3747 GND.n2280 585
R729 GND.n4481 GND.n4480 585
R730 GND.n4482 GND.n4481 585
R731 GND.n2281 GND.n2279 585
R732 GND.n3710 GND.n2279 585
R733 GND.n2284 GND.n2283 585
R734 GND.n2283 GND.n2259 585
R735 GND.n2247 GND.n2246 585
R736 GND.n2257 GND.n2247 585
R737 GND.n4498 GND.n4497 585
R738 GND.n4497 GND.n4496 585
R739 GND.n4499 GND.n2236 585
R740 GND.n3698 GND.n2236 585
R741 GND.n4501 GND.n4500 585
R742 GND.n4502 GND.n4501 585
R743 GND.n2237 GND.n2235 585
R744 GND.n2235 GND.n2225 585
R745 GND.n2240 GND.n2239 585
R746 GND.n2239 GND.n2223 585
R747 GND.n2211 GND.n2210 585
R748 GND.n3126 GND.n2211 585
R749 GND.n4519 GND.n4518 585
R750 GND.n4518 GND.n4517 585
R751 GND.n4520 GND.n2205 585
R752 GND.n3129 GND.n2205 585
R753 GND.n4522 GND.n4521 585
R754 GND.n4523 GND.n4522 585
R755 GND.n2191 GND.n2190 585
R756 GND.n3659 GND.n2191 585
R757 GND.n4533 GND.n4532 585
R758 GND.n4532 GND.n4531 585
R759 GND.n4534 GND.n2185 585
R760 GND.n3634 GND.n2185 585
R761 GND.n4536 GND.n4535 585
R762 GND.n4537 GND.n4536 585
R763 GND.n2173 GND.n2172 585
R764 GND.n3145 GND.n2173 585
R765 GND.n4547 GND.n4546 585
R766 GND.n4546 GND.n4545 585
R767 GND.n4548 GND.n2167 585
R768 GND.n3148 GND.n2167 585
R769 GND.n4550 GND.n4549 585
R770 GND.n4551 GND.n4550 585
R771 GND.n2153 GND.n2152 585
R772 GND.n3578 GND.n2153 585
R773 GND.n4561 GND.n4560 585
R774 GND.n4560 GND.n4559 585
R775 GND.n4562 GND.n2147 585
R776 GND.n3584 GND.n2147 585
R777 GND.n4564 GND.n4563 585
R778 GND.n4565 GND.n4564 585
R779 GND.n2133 GND.n2132 585
R780 GND.n3563 GND.n2133 585
R781 GND.n4575 GND.n4574 585
R782 GND.n4574 GND.n4573 585
R783 GND.n4576 GND.n2127 585
R784 GND.n3554 GND.n2127 585
R785 GND.n4578 GND.n4577 585
R786 GND.n4579 GND.n4578 585
R787 GND.n2113 GND.n2112 585
R788 GND.n3515 GND.n2113 585
R789 GND.n4589 GND.n4588 585
R790 GND.n4588 GND.n4587 585
R791 GND.n4590 GND.n2103 585
R792 GND.n3507 GND.n2103 585
R793 GND.n4592 GND.n4591 585
R794 GND.n4593 GND.n4592 585
R795 GND.n2104 GND.n2102 585
R796 GND.n3489 GND.n2102 585
R797 GND.n2106 GND.n2105 585
R798 GND.n2105 GND.n2090 585
R799 GND.n2079 GND.n2078 585
R800 GND.n2088 GND.n2079 585
R801 GND.n4610 GND.n4609 585
R802 GND.n4609 GND.n4608 585
R803 GND.n2076 GND.n2074 585
R804 GND.n3478 GND.n2074 585
R805 GND.n4615 GND.n4614 585
R806 GND.n4616 GND.n4615 585
R807 GND.n2075 GND.n2073 585
R808 GND.n2073 GND.n2063 585
R809 GND.n3276 GND.n3275 585
R810 GND.n3274 GND.n3211 585
R811 GND.n3273 GND.n3210 585
R812 GND.n3278 GND.n3210 585
R813 GND.n3272 GND.n3271 585
R814 GND.n3270 GND.n3269 585
R815 GND.n3268 GND.n3267 585
R816 GND.n3266 GND.n3265 585
R817 GND.n3264 GND.n3263 585
R818 GND.n3262 GND.n3261 585
R819 GND.n3260 GND.n3259 585
R820 GND.n3258 GND.n3257 585
R821 GND.n3256 GND.n3255 585
R822 GND.n3254 GND.n3253 585
R823 GND.n3252 GND.n3251 585
R824 GND.n3250 GND.n3249 585
R825 GND.n3248 GND.n3247 585
R826 GND.n3246 GND.n3245 585
R827 GND.n3244 GND.n3243 585
R828 GND.n3242 GND.n3241 585
R829 GND.n3240 GND.n3239 585
R830 GND.n3238 GND.n3237 585
R831 GND.n3236 GND.n3199 585
R832 GND.n3280 GND.n3198 585
R833 GND.n3885 GND.n3091 585
R834 GND.n3884 GND.n3883 585
R835 GND.n3807 GND.n3806 585
R836 GND.n3841 GND.n3840 585
R837 GND.n3843 GND.n3842 585
R838 GND.n3845 GND.n3844 585
R839 GND.n3847 GND.n3846 585
R840 GND.n3849 GND.n3848 585
R841 GND.n3851 GND.n3850 585
R842 GND.n3853 GND.n3852 585
R843 GND.n3855 GND.n3854 585
R844 GND.n3857 GND.n3856 585
R845 GND.n3859 GND.n3858 585
R846 GND.n3861 GND.n3860 585
R847 GND.n3863 GND.n3862 585
R848 GND.n3865 GND.n3864 585
R849 GND.n3867 GND.n3866 585
R850 GND.n3869 GND.n3868 585
R851 GND.n3871 GND.n3870 585
R852 GND.n3874 GND.n3873 585
R853 GND.n3872 GND.n3819 585
R854 GND.n3878 GND.n3818 585
R855 GND.n3880 GND.n3879 585
R856 GND.n3881 GND.n3880 585
R857 GND.n3889 GND.n3888 585
R858 GND.n3890 GND.n3889 585
R859 GND.n3092 GND.n2369 585
R860 GND.n4434 GND.n2369 585
R861 GND.n3802 GND.n3801 585
R862 GND.n3801 GND.n2361 585
R863 GND.n3800 GND.n3094 585
R864 GND.n3800 GND.n3799 585
R865 GND.n3764 GND.n3095 585
R866 GND.n3772 GND.n3095 585
R867 GND.n3765 GND.n2345 585
R868 GND.n4448 GND.n2345 585
R869 GND.n3767 GND.n3766 585
R870 GND.n3768 GND.n3767 585
R871 GND.n3102 GND.n2326 585
R872 GND.n4454 GND.n2326 585
R873 GND.n3758 GND.n3757 585
R874 GND.n3757 GND.n2318 585
R875 GND.n3756 GND.n3104 585
R876 GND.n3756 GND.n2316 585
R877 GND.n3755 GND.n3754 585
R878 GND.n3755 GND.n2302 585
R879 GND.n3106 GND.n3105 585
R880 GND.n3105 GND.n2300 585
R881 GND.n3750 GND.n2293 585
R882 GND.n4476 GND.n2293 585
R883 GND.n3749 GND.n3748 585
R884 GND.n3748 GND.n3747 585
R885 GND.n3108 GND.n2277 585
R886 GND.n4482 GND.n2277 585
R887 GND.n3709 GND.n3708 585
R888 GND.n3710 GND.n3709 585
R889 GND.n3118 GND.n3117 585
R890 GND.n3117 GND.n2259 585
R891 GND.n3703 GND.n3702 585
R892 GND.n3702 GND.n2257 585
R893 GND.n3701 GND.n2250 585
R894 GND.n4496 GND.n2250 585
R895 GND.n3700 GND.n3699 585
R896 GND.n3699 GND.n3698 585
R897 GND.n3120 GND.n2233 585
R898 GND.n4502 GND.n2233 585
R899 GND.n3649 GND.n3648 585
R900 GND.n3649 GND.n2225 585
R901 GND.n3650 GND.n3644 585
R902 GND.n3650 GND.n2223 585
R903 GND.n3652 GND.n3651 585
R904 GND.n3651 GND.n3126 585
R905 GND.n3653 GND.n2213 585
R906 GND.n4517 GND.n2213 585
R907 GND.n3655 GND.n3654 585
R908 GND.n3654 GND.n3129 585
R909 GND.n3656 GND.n2203 585
R910 GND.n4523 GND.n2203 585
R911 GND.n3658 GND.n3657 585
R912 GND.n3659 GND.n3658 585
R913 GND.n3134 GND.n2193 585
R914 GND.n4531 GND.n2193 585
R915 GND.n3636 GND.n3635 585
R916 GND.n3635 GND.n3634 585
R917 GND.n3136 GND.n2184 585
R918 GND.n4537 GND.n2184 585
R919 GND.n3169 GND.n3168 585
R920 GND.n3168 GND.n3145 585
R921 GND.n3170 GND.n2175 585
R922 GND.n4545 GND.n2175 585
R923 GND.n3172 GND.n3171 585
R924 GND.n3171 GND.n3148 585
R925 GND.n3173 GND.n2165 585
R926 GND.n4551 GND.n2165 585
R927 GND.n3580 GND.n3579 585
R928 GND.n3579 GND.n3578 585
R929 GND.n3581 GND.n2155 585
R930 GND.n4559 GND.n2155 585
R931 GND.n3583 GND.n3582 585
R932 GND.n3584 GND.n3583 585
R933 GND.n3160 GND.n2145 585
R934 GND.n4565 GND.n2145 585
R935 GND.n3562 GND.n3561 585
R936 GND.n3563 GND.n3562 585
R937 GND.n3176 GND.n2135 585
R938 GND.n4573 GND.n2135 585
R939 GND.n3556 GND.n3555 585
R940 GND.n3555 GND.n3554 585
R941 GND.n3178 GND.n2125 585
R942 GND.n4579 GND.n2125 585
R943 GND.n3514 GND.n3513 585
R944 GND.n3515 GND.n3514 585
R945 GND.n3182 GND.n2115 585
R946 GND.n4587 GND.n2115 585
R947 GND.n3509 GND.n3508 585
R948 GND.n3508 GND.n3507 585
R949 GND.n3184 GND.n2100 585
R950 GND.n4593 GND.n2100 585
R951 GND.n3488 GND.n3487 585
R952 GND.n3489 GND.n3488 585
R953 GND.n3194 GND.n3193 585
R954 GND.n3193 GND.n2090 585
R955 GND.n3483 GND.n3482 585
R956 GND.n3482 GND.n2088 585
R957 GND.n3481 GND.n2080 585
R958 GND.n4608 GND.n2080 585
R959 GND.n3480 GND.n3479 585
R960 GND.n3479 GND.n3478 585
R961 GND.n3196 GND.n2071 585
R962 GND.n4616 GND.n2071 585
R963 GND.n3282 GND.n3281 585
R964 GND.n3281 GND.n2063 585
R965 GND.n4699 GND.n4698 585
R966 GND.n4700 GND.n4699 585
R967 GND.n1177 GND.n1175 585
R968 GND.n2040 GND.n1175 585
R969 GND.n2033 GND.n1501 585
R970 GND.n1501 GND.n1493 585
R971 GND.n2035 GND.n2034 585
R972 GND.n2036 GND.n2035 585
R973 GND.n1502 GND.n1500 585
R974 GND.n2008 GND.n1500 585
R975 GND.n2028 GND.n2027 585
R976 GND.n2027 GND.n2026 585
R977 GND.n1505 GND.n1504 585
R978 GND.n2023 GND.n1505 585
R979 GND.n1999 GND.n1524 585
R980 GND.n1524 GND.n1523 585
R981 GND.n2001 GND.n2000 585
R982 GND.n2002 GND.n2001 585
R983 GND.n1525 GND.n1522 585
R984 GND.n1989 GND.n1522 585
R985 GND.n1994 GND.n1993 585
R986 GND.n1993 GND.n1992 585
R987 GND.n1528 GND.n1527 585
R988 GND.n1987 GND.n1528 585
R989 GND.n1975 GND.n1547 585
R990 GND.n1547 GND.n1546 585
R991 GND.n1977 GND.n1976 585
R992 GND.n1978 GND.n1977 585
R993 GND.n1548 GND.n1545 585
R994 GND.n1965 GND.n1545 585
R995 GND.n1970 GND.n1969 585
R996 GND.n1969 GND.n1968 585
R997 GND.n1551 GND.n1550 585
R998 GND.n1962 GND.n1551 585
R999 GND.n1950 GND.n1569 585
R1000 GND.n1569 GND.n1568 585
R1001 GND.n1952 GND.n1951 585
R1002 GND.n1953 GND.n1952 585
R1003 GND.n1570 GND.n1567 585
R1004 GND.n1913 GND.n1567 585
R1005 GND.n1907 GND.n1906 585
R1006 GND.n1908 GND.n1907 585
R1007 GND.n1905 GND.n1904 585
R1008 GND.n1905 GND.n1610 585
R1009 GND.n1903 GND.n1604 585
R1010 GND.n1922 GND.n1604 585
R1011 GND.n1927 GND.n1926 585
R1012 GND.n1926 GND.n1925 585
R1013 GND.n1929 GND.n1928 585
R1014 GND.n1930 GND.n1929 585
R1015 GND.n1603 GND.n1602 585
R1016 GND.n1603 GND.n1595 585
R1017 GND.n1601 GND.n1576 585
R1018 GND.n1601 GND.n1588 585
R1019 GND.n1580 GND.n1577 585
R1020 GND.n1939 GND.n1580 585
R1021 GND.n1945 GND.n1944 585
R1022 GND.n1944 GND.n1943 585
R1023 GND.n1579 GND.n1578 585
R1024 GND.n1680 GND.n1579 585
R1025 GND.n1879 GND.n1878 585
R1026 GND.n1880 GND.n1879 585
R1027 GND.n1684 GND.n1683 585
R1028 GND.n1868 GND.n1683 585
R1029 GND.n1874 GND.n1873 585
R1030 GND.n1873 GND.n1872 585
R1031 GND.n1687 GND.n1686 585
R1032 GND.n1866 GND.n1687 585
R1033 GND.n1854 GND.n1705 585
R1034 GND.n1705 GND.n1704 585
R1035 GND.n1856 GND.n1855 585
R1036 GND.n1857 GND.n1856 585
R1037 GND.n1706 GND.n1702 585
R1038 GND.n1844 GND.n1702 585
R1039 GND.n1849 GND.n1848 585
R1040 GND.n1848 GND.n1847 585
R1041 GND.n1709 GND.n1708 585
R1042 GND.n1841 GND.n1709 585
R1043 GND.n1829 GND.n1728 585
R1044 GND.n1728 GND.n1727 585
R1045 GND.n1831 GND.n1830 585
R1046 GND.n1832 GND.n1831 585
R1047 GND.n1729 GND.n1726 585
R1048 GND.n1819 GND.n1726 585
R1049 GND.n1824 GND.n1823 585
R1050 GND.n1823 GND.n1822 585
R1051 GND.n1733 GND.n1732 585
R1052 GND.n1771 GND.n1733 585
R1053 GND.n1003 GND.n1002 585
R1054 GND.n1757 GND.n1003 585
R1055 GND.n4775 GND.n4774 585
R1056 GND.n4774 GND.n4773 585
R1057 GND.n4776 GND.n998 585
R1058 GND.n1078 GND.n998 585
R1059 GND.n4778 GND.n4777 585
R1060 GND.n4779 GND.n4778 585
R1061 GND.n1032 GND.n997 585
R1062 GND.n1035 GND.n1034 585
R1063 GND.n1033 GND.n1030 585
R1064 GND.n1040 GND.n1039 585
R1065 GND.n1042 GND.n1041 585
R1066 GND.n1045 GND.n1044 585
R1067 GND.n1043 GND.n1028 585
R1068 GND.n1050 GND.n1049 585
R1069 GND.n1052 GND.n1051 585
R1070 GND.n1054 GND.n1053 585
R1071 GND.n1056 GND.n1055 585
R1072 GND.n1060 GND.n1022 585
R1073 GND.n1062 GND.n1061 585
R1074 GND.n1064 GND.n1063 585
R1075 GND.n1066 GND.n1065 585
R1076 GND.n1019 GND.n1018 585
R1077 GND.n1070 GND.n1020 585
R1078 GND.n1071 GND.n1015 585
R1079 GND.n1072 GND.n975 585
R1080 GND.n4800 GND.n975 585
R1081 GND.n4670 GND.n1169 585
R1082 GND.n4638 GND.n1204 585
R1083 GND.n4674 GND.n1201 585
R1084 GND.n4675 GND.n1200 585
R1085 GND.n4676 GND.n1199 585
R1086 GND.n4641 GND.n1197 585
R1087 GND.n4680 GND.n1196 585
R1088 GND.n4681 GND.n1195 585
R1089 GND.n4682 GND.n1194 585
R1090 GND.n4644 GND.n1192 585
R1091 GND.n4686 GND.n1191 585
R1092 GND.n4688 GND.n1185 585
R1093 GND.n4689 GND.n1184 585
R1094 GND.n4648 GND.n1182 585
R1095 GND.n4693 GND.n1181 585
R1096 GND.n4694 GND.n1180 585
R1097 GND.n4695 GND.n1176 585
R1098 GND.n4651 GND.n1176 585
R1099 GND.n4702 GND.n4701 585
R1100 GND.n4701 GND.n4700 585
R1101 GND.n4703 GND.n1168 585
R1102 GND.n2040 GND.n1168 585
R1103 GND.n1492 GND.n1163 585
R1104 GND.n1493 GND.n1492 585
R1105 GND.n4707 GND.n1162 585
R1106 GND.n2036 GND.n1162 585
R1107 GND.n4708 GND.n1161 585
R1108 GND.n2008 GND.n1161 585
R1109 GND.n4709 GND.n1160 585
R1110 GND.n2026 GND.n1160 585
R1111 GND.n1511 GND.n1155 585
R1112 GND.n2023 GND.n1511 585
R1113 GND.n4713 GND.n1154 585
R1114 GND.n1523 GND.n1154 585
R1115 GND.n4714 GND.n1153 585
R1116 GND.n2002 GND.n1153 585
R1117 GND.n4715 GND.n1152 585
R1118 GND.n1989 GND.n1152 585
R1119 GND.n1530 GND.n1147 585
R1120 GND.n1992 GND.n1530 585
R1121 GND.n4719 GND.n1146 585
R1122 GND.n1987 GND.n1146 585
R1123 GND.n4720 GND.n1145 585
R1124 GND.n1546 GND.n1145 585
R1125 GND.n4721 GND.n1144 585
R1126 GND.n1978 GND.n1144 585
R1127 GND.n1964 GND.n1139 585
R1128 GND.n1965 GND.n1964 585
R1129 GND.n4725 GND.n1138 585
R1130 GND.n1968 GND.n1138 585
R1131 GND.n4726 GND.n1137 585
R1132 GND.n1962 GND.n1137 585
R1133 GND.n4727 GND.n1136 585
R1134 GND.n1568 GND.n1136 585
R1135 GND.n1564 GND.n1131 585
R1136 GND.n1953 GND.n1564 585
R1137 GND.n4731 GND.n1130 585
R1138 GND.n1913 GND.n1130 585
R1139 GND.n4732 GND.n1129 585
R1140 GND.n1908 GND.n1129 585
R1141 GND.n4733 GND.n1128 585
R1142 GND.n1610 GND.n1128 585
R1143 GND.n1608 GND.n1123 585
R1144 GND.n1922 GND.n1608 585
R1145 GND.n4737 GND.n1122 585
R1146 GND.n1925 GND.n1122 585
R1147 GND.n4738 GND.n1121 585
R1148 GND.n1930 GND.n1121 585
R1149 GND.n4739 GND.n1120 585
R1150 GND.n1595 GND.n1120 585
R1151 GND.n1587 GND.n1115 585
R1152 GND.n1588 GND.n1587 585
R1153 GND.n4743 GND.n1114 585
R1154 GND.n1939 GND.n1114 585
R1155 GND.n4744 GND.n1113 585
R1156 GND.n1943 GND.n1113 585
R1157 GND.n4745 GND.n1112 585
R1158 GND.n1680 GND.n1112 585
R1159 GND.n1679 GND.n1107 585
R1160 GND.n1880 GND.n1679 585
R1161 GND.n4749 GND.n1106 585
R1162 GND.n1868 GND.n1106 585
R1163 GND.n4750 GND.n1105 585
R1164 GND.n1872 GND.n1105 585
R1165 GND.n4751 GND.n1104 585
R1166 GND.n1866 GND.n1104 585
R1167 GND.n1703 GND.n1099 585
R1168 GND.n1704 GND.n1703 585
R1169 GND.n4755 GND.n1098 585
R1170 GND.n1857 GND.n1098 585
R1171 GND.n4756 GND.n1097 585
R1172 GND.n1844 GND.n1097 585
R1173 GND.n4757 GND.n1096 585
R1174 GND.n1847 GND.n1096 585
R1175 GND.n1715 GND.n1091 585
R1176 GND.n1841 GND.n1715 585
R1177 GND.n4761 GND.n1090 585
R1178 GND.n1727 GND.n1090 585
R1179 GND.n4762 GND.n1089 585
R1180 GND.n1832 GND.n1089 585
R1181 GND.n4763 GND.n1088 585
R1182 GND.n1819 GND.n1088 585
R1183 GND.n1735 GND.n1083 585
R1184 GND.n1822 GND.n1735 585
R1185 GND.n4767 GND.n1082 585
R1186 GND.n1771 GND.n1082 585
R1187 GND.n4768 GND.n1081 585
R1188 GND.n1757 GND.n1081 585
R1189 GND.n4769 GND.n1005 585
R1190 GND.n4773 GND.n1005 585
R1191 GND.n1080 GND.n1079 585
R1192 GND.n1079 GND.n1078 585
R1193 GND.n1077 GND.n995 585
R1194 GND.n4779 GND.n995 585
R1195 GND.n261 GND.n260 585
R1196 GND.n5748 GND.n261 585
R1197 GND.n5800 GND.n5799 585
R1198 GND.n5799 GND.n5798 585
R1199 GND.n5801 GND.n256 585
R1200 GND.n4250 GND.n256 585
R1201 GND.n5803 GND.n5802 585
R1202 GND.n5804 GND.n5803 585
R1203 GND.n241 GND.n240 585
R1204 GND.n4256 GND.n241 585
R1205 GND.n5812 GND.n5811 585
R1206 GND.n5811 GND.n5810 585
R1207 GND.n5813 GND.n236 585
R1208 GND.n4262 GND.n236 585
R1209 GND.n5815 GND.n5814 585
R1210 GND.n5816 GND.n5815 585
R1211 GND.n220 GND.n219 585
R1212 GND.n4208 GND.n220 585
R1213 GND.n5824 GND.n5823 585
R1214 GND.n5823 GND.n5822 585
R1215 GND.n5825 GND.n215 585
R1216 GND.n4199 GND.n215 585
R1217 GND.n5827 GND.n5826 585
R1218 GND.n5828 GND.n5827 585
R1219 GND.n199 GND.n198 585
R1220 GND.n4193 GND.n199 585
R1221 GND.n5836 GND.n5835 585
R1222 GND.n5835 GND.n5834 585
R1223 GND.n5837 GND.n194 585
R1224 GND.n4185 GND.n194 585
R1225 GND.n5839 GND.n5838 585
R1226 GND.n5840 GND.n5839 585
R1227 GND.n179 GND.n178 585
R1228 GND.n4179 GND.n179 585
R1229 GND.n5848 GND.n5847 585
R1230 GND.n5847 GND.n5846 585
R1231 GND.n5849 GND.n173 585
R1232 GND.n4171 GND.n173 585
R1233 GND.n5851 GND.n5850 585
R1234 GND.n5852 GND.n5851 585
R1235 GND.n174 GND.n172 585
R1236 GND.n4165 GND.n172 585
R1237 GND.n2927 GND.n2926 585
R1238 GND.n2931 GND.n2927 585
R1239 GND.n4311 GND.n4310 585
R1240 GND.n4310 GND.n4309 585
R1241 GND.n4312 GND.n152 585
R1242 GND.n5859 GND.n152 585
R1243 GND.n4313 GND.n2920 585
R1244 GND.n4149 GND.n2920 585
R1245 GND.n4315 GND.n4314 585
R1246 GND.n4319 GND.n4315 585
R1247 GND.n2921 GND.n2919 585
R1248 GND.n2919 GND.n2915 585
R1249 GND.n4142 GND.n4141 585
R1250 GND.n4141 GND.n2908 585
R1251 GND.n2899 GND.n2898 585
R1252 GND.n4328 GND.n2899 585
R1253 GND.n4335 GND.n4334 585
R1254 GND.n4334 GND.n4333 585
R1255 GND.n4336 GND.n2894 585
R1256 GND.n4135 GND.n2894 585
R1257 GND.n4338 GND.n4337 585
R1258 GND.n4339 GND.n4338 585
R1259 GND.n2877 GND.n2876 585
R1260 GND.n4115 GND.n2877 585
R1261 GND.n4347 GND.n4346 585
R1262 GND.n4346 GND.n4345 585
R1263 GND.n4348 GND.n2872 585
R1264 GND.n4108 GND.n2872 585
R1265 GND.n4350 GND.n4349 585
R1266 GND.n4351 GND.n4350 585
R1267 GND.n2856 GND.n2855 585
R1268 GND.n4100 GND.n2856 585
R1269 GND.n4359 GND.n4358 585
R1270 GND.n4358 GND.n4357 585
R1271 GND.n4360 GND.n2851 585
R1272 GND.n4093 GND.n2851 585
R1273 GND.n4362 GND.n4361 585
R1274 GND.n4363 GND.n4362 585
R1275 GND.n2836 GND.n2835 585
R1276 GND.n4085 GND.n2836 585
R1277 GND.n4371 GND.n4370 585
R1278 GND.n4370 GND.n4369 585
R1279 GND.n4372 GND.n2829 585
R1280 GND.n4078 GND.n2829 585
R1281 GND.n4374 GND.n4373 585
R1282 GND.n4375 GND.n4374 585
R1283 GND.n2830 GND.n2828 585
R1284 GND.n2999 GND.n2828 585
R1285 GND.n2812 GND.n2805 585
R1286 GND.n4381 GND.n2812 585
R1287 GND.n4386 GND.n2803 585
R1288 GND.n2994 GND.n2803 585
R1289 GND.n4388 GND.n4387 585
R1290 GND.n4389 GND.n4388 585
R1291 GND.n2802 GND.n2801 585
R1292 GND.n2800 GND.n2799 585
R1293 GND.n2798 GND.n2797 585
R1294 GND.n2796 GND.n2795 585
R1295 GND.n2794 GND.n2793 585
R1296 GND.n2792 GND.n2791 585
R1297 GND.n2790 GND.n2789 585
R1298 GND.n2380 GND.n2379 585
R1299 GND.n4427 GND.n4426 585
R1300 GND.n4426 GND.n4425 585
R1301 GND.n4243 GND.n4242 585
R1302 GND.n4241 GND.n4221 585
R1303 GND.n4240 GND.n4239 585
R1304 GND.n4233 GND.n4222 585
R1305 GND.n4235 GND.n4234 585
R1306 GND.n4232 GND.n4231 585
R1307 GND.n4230 GND.n4229 585
R1308 GND.n4226 GND.n4225 585
R1309 GND.n4224 GND.n273 585
R1310 GND.n5790 GND.n273 585
R1311 GND.n4246 GND.n309 585
R1312 GND.n5748 GND.n309 585
R1313 GND.n4247 GND.n264 585
R1314 GND.n5798 GND.n264 585
R1315 GND.n4249 GND.n4248 585
R1316 GND.n4250 GND.n4249 585
R1317 GND.n2961 GND.n254 585
R1318 GND.n5804 GND.n254 585
R1319 GND.n4258 GND.n4257 585
R1320 GND.n4257 GND.n4256 585
R1321 GND.n4259 GND.n243 585
R1322 GND.n5810 GND.n243 585
R1323 GND.n4261 GND.n4260 585
R1324 GND.n4262 GND.n4261 585
R1325 GND.n2957 GND.n234 585
R1326 GND.n5816 GND.n234 585
R1327 GND.n4207 GND.n4206 585
R1328 GND.n4208 GND.n4207 585
R1329 GND.n2964 GND.n223 585
R1330 GND.n5822 GND.n223 585
R1331 GND.n4201 GND.n4200 585
R1332 GND.n4200 GND.n4199 585
R1333 GND.n2966 GND.n213 585
R1334 GND.n5828 GND.n213 585
R1335 GND.n4192 GND.n4191 585
R1336 GND.n4193 GND.n4192 585
R1337 GND.n2969 GND.n202 585
R1338 GND.n5834 GND.n202 585
R1339 GND.n4187 GND.n4186 585
R1340 GND.n4186 GND.n4185 585
R1341 GND.n2971 GND.n192 585
R1342 GND.n5840 GND.n192 585
R1343 GND.n4178 GND.n4177 585
R1344 GND.n4179 GND.n4178 585
R1345 GND.n2974 GND.n182 585
R1346 GND.n5846 GND.n182 585
R1347 GND.n4173 GND.n4172 585
R1348 GND.n4172 GND.n4171 585
R1349 GND.n2976 GND.n170 585
R1350 GND.n5852 GND.n170 585
R1351 GND.n4164 GND.n4163 585
R1352 GND.n4165 GND.n4164 585
R1353 GND.n4160 GND.n4159 585
R1354 GND.n4159 GND.n2931 585
R1355 GND.n148 GND.n146 585
R1356 GND.n4309 GND.n148 585
R1357 GND.n5861 GND.n5860 585
R1358 GND.n5860 GND.n5859 585
R1359 GND.n147 GND.n145 585
R1360 GND.n4149 GND.n147 585
R1361 GND.n4126 GND.n2917 585
R1362 GND.n4319 GND.n2917 585
R1363 GND.n4128 GND.n4127 585
R1364 GND.n4128 GND.n2915 585
R1365 GND.n4130 GND.n4129 585
R1366 GND.n4129 GND.n2908 585
R1367 GND.n4131 GND.n2907 585
R1368 GND.n4328 GND.n2907 585
R1369 GND.n4132 GND.n2902 585
R1370 GND.n4333 GND.n2902 585
R1371 GND.n4134 GND.n4133 585
R1372 GND.n4135 GND.n4134 585
R1373 GND.n2979 GND.n2892 585
R1374 GND.n4339 GND.n2892 585
R1375 GND.n4117 GND.n4116 585
R1376 GND.n4116 GND.n4115 585
R1377 GND.n2981 GND.n2880 585
R1378 GND.n4345 GND.n2880 585
R1379 GND.n4107 GND.n4106 585
R1380 GND.n4108 GND.n4107 585
R1381 GND.n2983 GND.n2870 585
R1382 GND.n4351 GND.n2870 585
R1383 GND.n4102 GND.n4101 585
R1384 GND.n4101 GND.n4100 585
R1385 GND.n2985 GND.n2859 585
R1386 GND.n4357 GND.n2859 585
R1387 GND.n4092 GND.n4091 585
R1388 GND.n4093 GND.n4092 585
R1389 GND.n2987 GND.n2849 585
R1390 GND.n4363 GND.n2849 585
R1391 GND.n4087 GND.n4086 585
R1392 GND.n4086 GND.n4085 585
R1393 GND.n2989 GND.n2838 585
R1394 GND.n4369 GND.n2838 585
R1395 GND.n3006 GND.n3005 585
R1396 GND.n4078 GND.n3006 585
R1397 GND.n2991 GND.n2826 585
R1398 GND.n4375 GND.n2826 585
R1399 GND.n3001 GND.n3000 585
R1400 GND.n3000 GND.n2999 585
R1401 GND.n2998 GND.n2810 585
R1402 GND.n4381 GND.n2810 585
R1403 GND.n2997 GND.n2995 585
R1404 GND.n2995 GND.n2994 585
R1405 GND.n2993 GND.n2381 585
R1406 GND.n4389 GND.n2381 585
R1407 GND.n5795 GND.n266 585
R1408 GND.n5748 GND.n266 585
R1409 GND.n5797 GND.n5796 585
R1410 GND.n5798 GND.n5797 585
R1411 GND.n251 GND.n250 585
R1412 GND.n4250 GND.n251 585
R1413 GND.n5806 GND.n5805 585
R1414 GND.n5805 GND.n5804 585
R1415 GND.n5807 GND.n245 585
R1416 GND.n4256 GND.n245 585
R1417 GND.n5809 GND.n5808 585
R1418 GND.n5810 GND.n5809 585
R1419 GND.n231 GND.n230 585
R1420 GND.n4262 GND.n231 585
R1421 GND.n5818 GND.n5817 585
R1422 GND.n5817 GND.n5816 585
R1423 GND.n5819 GND.n225 585
R1424 GND.n4208 GND.n225 585
R1425 GND.n5821 GND.n5820 585
R1426 GND.n5822 GND.n5821 585
R1427 GND.n210 GND.n209 585
R1428 GND.n4199 GND.n210 585
R1429 GND.n5830 GND.n5829 585
R1430 GND.n5829 GND.n5828 585
R1431 GND.n5831 GND.n204 585
R1432 GND.n4193 GND.n204 585
R1433 GND.n5833 GND.n5832 585
R1434 GND.n5834 GND.n5833 585
R1435 GND.n189 GND.n188 585
R1436 GND.n4185 GND.n189 585
R1437 GND.n5842 GND.n5841 585
R1438 GND.n5841 GND.n5840 585
R1439 GND.n5843 GND.n184 585
R1440 GND.n4179 GND.n184 585
R1441 GND.n5845 GND.n5844 585
R1442 GND.n5846 GND.n5845 585
R1443 GND.n167 GND.n165 585
R1444 GND.n4171 GND.n167 585
R1445 GND.n5854 GND.n5853 585
R1446 GND.n5853 GND.n5852 585
R1447 GND.n166 GND.n164 585
R1448 GND.n4165 GND.n166 585
R1449 GND.n2930 GND.n2929 585
R1450 GND.n2931 GND.n2930 585
R1451 GND.n156 GND.n154 585
R1452 GND.n4309 GND.n154 585
R1453 GND.n5858 GND.n5857 585
R1454 GND.n5859 GND.n5858 585
R1455 GND.n155 GND.n153 585
R1456 GND.n4149 GND.n153 585
R1457 GND.n4318 GND.n4317 585
R1458 GND.n4319 GND.n4318 585
R1459 GND.n4316 GND.n162 585
R1460 GND.n4316 GND.n2915 585
R1461 GND.n2904 GND.n2903 585
R1462 GND.n2908 GND.n2904 585
R1463 GND.n4330 GND.n4329 585
R1464 GND.n4329 GND.n4328 585
R1465 GND.n4332 GND.n4331 585
R1466 GND.n4333 GND.n4332 585
R1467 GND.n2889 GND.n2888 585
R1468 GND.n4135 GND.n2889 585
R1469 GND.n4341 GND.n4340 585
R1470 GND.n4340 GND.n4339 585
R1471 GND.n4342 GND.n2882 585
R1472 GND.n4115 GND.n2882 585
R1473 GND.n4344 GND.n4343 585
R1474 GND.n4345 GND.n4344 585
R1475 GND.n2867 GND.n2866 585
R1476 GND.n4108 GND.n2867 585
R1477 GND.n4353 GND.n4352 585
R1478 GND.n4352 GND.n4351 585
R1479 GND.n4354 GND.n2861 585
R1480 GND.n4100 GND.n2861 585
R1481 GND.n4356 GND.n4355 585
R1482 GND.n4357 GND.n4356 585
R1483 GND.n2846 GND.n2845 585
R1484 GND.n4093 GND.n2846 585
R1485 GND.n4365 GND.n4364 585
R1486 GND.n4364 GND.n4363 585
R1487 GND.n4366 GND.n2840 585
R1488 GND.n4085 GND.n2840 585
R1489 GND.n4368 GND.n4367 585
R1490 GND.n4369 GND.n4368 585
R1491 GND.n2823 GND.n2822 585
R1492 GND.n4078 GND.n2823 585
R1493 GND.n4377 GND.n4376 585
R1494 GND.n4376 GND.n4375 585
R1495 GND.n4378 GND.n2814 585
R1496 GND.n2999 GND.n2814 585
R1497 GND.n4380 GND.n4379 585
R1498 GND.n4381 GND.n4380 585
R1499 GND.n2815 GND.n2813 585
R1500 GND.n2994 GND.n2813 585
R1501 GND.n2816 GND.n2398 585
R1502 GND.n4389 GND.n2398 585
R1503 GND.n4423 GND.n4422 585
R1504 GND.n4421 GND.n2397 585
R1505 GND.n4420 GND.n2396 585
R1506 GND.n4425 GND.n2396 585
R1507 GND.n4419 GND.n4418 585
R1508 GND.n4417 GND.n4416 585
R1509 GND.n4415 GND.n4414 585
R1510 GND.n4412 GND.n4411 585
R1511 GND.n4410 GND.n4409 585
R1512 GND.n4408 GND.n4407 585
R1513 GND.n4406 GND.n4405 585
R1514 GND.n4404 GND.n4403 585
R1515 GND.n4402 GND.n4401 585
R1516 GND.n4400 GND.n4399 585
R1517 GND.n4398 GND.n4397 585
R1518 GND.n4396 GND.n2418 585
R1519 GND.n2422 GND.n2419 585
R1520 GND.n4392 GND.n4391 585
R1521 GND.n308 GND.n303 585
R1522 GND.n5756 GND.n5755 585
R1523 GND.n5758 GND.n5757 585
R1524 GND.n5760 GND.n5759 585
R1525 GND.n5762 GND.n5761 585
R1526 GND.n5764 GND.n5763 585
R1527 GND.n5766 GND.n5765 585
R1528 GND.n5768 GND.n5767 585
R1529 GND.n5770 GND.n5769 585
R1530 GND.n5772 GND.n5771 585
R1531 GND.n5774 GND.n5773 585
R1532 GND.n5779 GND.n5778 585
R1533 GND.n5781 GND.n5780 585
R1534 GND.n5783 GND.n5782 585
R1535 GND.n5785 GND.n5784 585
R1536 GND.n5786 GND.n287 585
R1537 GND.n5788 GND.n5787 585
R1538 GND.n271 GND.n270 585
R1539 GND.n5792 GND.n5791 585
R1540 GND.n5791 GND.n5790 585
R1541 GND.n5750 GND.n5749 585
R1542 GND.n5749 GND.n5748 585
R1543 GND.n307 GND.n263 585
R1544 GND.n5798 GND.n263 585
R1545 GND.n4252 GND.n4251 585
R1546 GND.n4251 GND.n4250 585
R1547 GND.n4253 GND.n253 585
R1548 GND.n5804 GND.n253 585
R1549 GND.n4255 GND.n4254 585
R1550 GND.n4256 GND.n4255 585
R1551 GND.n4213 GND.n242 585
R1552 GND.n5810 GND.n242 585
R1553 GND.n4212 GND.n2956 585
R1554 GND.n4262 GND.n2956 585
R1555 GND.n4211 GND.n233 585
R1556 GND.n5816 GND.n233 585
R1557 GND.n4210 GND.n4209 585
R1558 GND.n4209 GND.n4208 585
R1559 GND.n2962 GND.n222 585
R1560 GND.n5822 GND.n222 585
R1561 GND.n4198 GND.n4197 585
R1562 GND.n4199 GND.n4198 585
R1563 GND.n4196 GND.n212 585
R1564 GND.n5828 GND.n212 585
R1565 GND.n4195 GND.n4194 585
R1566 GND.n4194 GND.n4193 585
R1567 GND.n2967 GND.n201 585
R1568 GND.n5834 GND.n201 585
R1569 GND.n4184 GND.n4183 585
R1570 GND.n4185 GND.n4184 585
R1571 GND.n4182 GND.n191 585
R1572 GND.n5840 GND.n191 585
R1573 GND.n4181 GND.n4180 585
R1574 GND.n4180 GND.n4179 585
R1575 GND.n2972 GND.n181 585
R1576 GND.n5846 GND.n181 585
R1577 GND.n4170 GND.n4169 585
R1578 GND.n4171 GND.n4170 585
R1579 GND.n4168 GND.n169 585
R1580 GND.n5852 GND.n169 585
R1581 GND.n4167 GND.n4166 585
R1582 GND.n4166 GND.n4165 585
R1583 GND.n4157 GND.n4154 585
R1584 GND.n4157 GND.n2931 585
R1585 GND.n4153 GND.n2928 585
R1586 GND.n4309 GND.n2928 585
R1587 GND.n4152 GND.n150 585
R1588 GND.n5859 GND.n150 585
R1589 GND.n4151 GND.n4150 585
R1590 GND.n4150 GND.n4149 585
R1591 GND.n4148 GND.n2916 585
R1592 GND.n4319 GND.n2916 585
R1593 GND.n4147 GND.n4146 585
R1594 GND.n4146 GND.n2915 585
R1595 GND.n4145 GND.n2977 585
R1596 GND.n4145 GND.n2908 585
R1597 GND.n4139 GND.n2906 585
R1598 GND.n4328 GND.n2906 585
R1599 GND.n4138 GND.n2901 585
R1600 GND.n4333 GND.n2901 585
R1601 GND.n4137 GND.n4136 585
R1602 GND.n4136 GND.n4135 585
R1603 GND.n2978 GND.n2891 585
R1604 GND.n4339 GND.n2891 585
R1605 GND.n4114 GND.n4113 585
R1606 GND.n4115 GND.n4114 585
R1607 GND.n4111 GND.n2879 585
R1608 GND.n4345 GND.n2879 585
R1609 GND.n4110 GND.n4109 585
R1610 GND.n4109 GND.n4108 585
R1611 GND.n2982 GND.n2869 585
R1612 GND.n4351 GND.n2869 585
R1613 GND.n4099 GND.n4098 585
R1614 GND.n4100 GND.n4099 585
R1615 GND.n4096 GND.n2858 585
R1616 GND.n4357 GND.n2858 585
R1617 GND.n4095 GND.n4094 585
R1618 GND.n4094 GND.n4093 585
R1619 GND.n2986 GND.n2848 585
R1620 GND.n4363 GND.n2848 585
R1621 GND.n4084 GND.n4083 585
R1622 GND.n4085 GND.n4084 585
R1623 GND.n4081 GND.n2837 585
R1624 GND.n4369 GND.n2837 585
R1625 GND.n4080 GND.n4079 585
R1626 GND.n4079 GND.n4078 585
R1627 GND.n2990 GND.n2825 585
R1628 GND.n4375 GND.n2825 585
R1629 GND.n2808 GND.n2807 585
R1630 GND.n2999 GND.n2808 585
R1631 GND.n4383 GND.n4382 585
R1632 GND.n4382 GND.n4381 585
R1633 GND.n4384 GND.n2424 585
R1634 GND.n2994 GND.n2424 585
R1635 GND.n4390 GND.n2425 585
R1636 GND.n4390 GND.n4389 585
R1637 GND.n4004 GND.n4003 585
R1638 GND.n4005 GND.n4004 585
R1639 GND.n3033 GND.n3031 585
R1640 GND.n3031 GND.n3028 585
R1641 GND.n2366 GND.n2365 585
R1642 GND.n3891 GND.n2366 585
R1643 GND.n4436 GND.n4435 585
R1644 GND.n4435 GND.n4434 585
R1645 GND.n4437 GND.n2363 585
R1646 GND.n3787 GND.n2363 585
R1647 GND.n4439 GND.n4438 585
R1648 GND.n4440 GND.n4439 585
R1649 GND.n2364 GND.n2362 585
R1650 GND.n3793 GND.n2362 585
R1651 GND.n3774 GND.n3771 585
R1652 GND.n3774 GND.n3773 585
R1653 GND.n3776 GND.n3775 585
R1654 GND.n3775 GND.n2346 585
R1655 GND.n3777 GND.n3770 585
R1656 GND.n3770 GND.n2344 585
R1657 GND.n3779 GND.n3778 585
R1658 GND.n3780 GND.n3779 585
R1659 GND.n2323 GND.n2322 585
R1660 GND.n3101 GND.n2323 585
R1661 GND.n4457 GND.n4456 585
R1662 GND.n4456 GND.n4455 585
R1663 GND.n4458 GND.n2320 585
R1664 GND.n3727 GND.n2320 585
R1665 GND.n4460 GND.n4459 585
R1666 GND.n4461 GND.n4460 585
R1667 GND.n2321 GND.n2319 585
R1668 GND.n3733 GND.n2319 585
R1669 GND.n2299 GND.n2298 585
R1670 GND.n3735 GND.n2299 585
R1671 GND.n4471 GND.n4470 585
R1672 GND.n4470 GND.n4469 585
R1673 GND.n4472 GND.n2296 585
R1674 GND.n3740 GND.n2296 585
R1675 GND.n4474 GND.n4473 585
R1676 GND.n4475 GND.n4474 585
R1677 GND.n2297 GND.n2295 585
R1678 GND.n3746 GND.n2295 585
R1679 GND.n3713 GND.n3712 585
R1680 GND.n3713 GND.n3110 585
R1681 GND.n3715 GND.n3714 585
R1682 GND.n3714 GND.n2278 585
R1683 GND.n3716 GND.n3711 585
R1684 GND.n3711 GND.n2276 585
R1685 GND.n3718 GND.n3717 585
R1686 GND.n3719 GND.n3718 585
R1687 GND.n2256 GND.n2255 585
R1688 GND.n3115 GND.n2256 585
R1689 GND.n4492 GND.n4491 585
R1690 GND.n4491 GND.n4490 585
R1691 GND.n4493 GND.n2253 585
R1692 GND.n3691 GND.n2253 585
R1693 GND.n4495 GND.n4494 585
R1694 GND.n4496 GND.n4495 585
R1695 GND.n2254 GND.n2252 585
R1696 GND.n3697 GND.n2252 585
R1697 GND.n2230 GND.n2229 585
R1698 GND.n3122 GND.n2230 585
R1699 GND.n4505 GND.n4504 585
R1700 GND.n4504 GND.n4503 585
R1701 GND.n4506 GND.n2227 585
R1702 GND.n3684 GND.n2227 585
R1703 GND.n4508 GND.n4507 585
R1704 GND.n4509 GND.n4508 585
R1705 GND.n2228 GND.n2226 585
R1706 GND.n3680 GND.n2226 585
R1707 GND.n3677 GND.n3676 585
R1708 GND.n3678 GND.n3677 585
R1709 GND.n3675 GND.n3127 585
R1710 GND.n3127 GND.n2214 585
R1711 GND.n3674 GND.n3673 585
R1712 GND.n3673 GND.n2212 585
R1713 GND.n3672 GND.n3128 585
R1714 GND.n3672 GND.n3671 585
R1715 GND.n2200 GND.n2199 585
R1716 GND.n3130 GND.n2200 585
R1717 GND.n4526 GND.n4525 585
R1718 GND.n4525 GND.n4524 585
R1719 GND.n4527 GND.n2197 585
R1720 GND.n3660 GND.n2197 585
R1721 GND.n4529 GND.n4528 585
R1722 GND.n4530 GND.n4529 585
R1723 GND.n2198 GND.n2196 585
R1724 GND.n2196 GND.n2192 585
R1725 GND.n3632 GND.n3631 585
R1726 GND.n3633 GND.n3632 585
R1727 GND.n2182 GND.n2181 585
R1728 GND.n3606 GND.n2182 585
R1729 GND.n4540 GND.n4539 585
R1730 GND.n4539 GND.n4538 585
R1731 GND.n4541 GND.n2179 585
R1732 GND.n3612 GND.n2179 585
R1733 GND.n4543 GND.n4542 585
R1734 GND.n4544 GND.n4543 585
R1735 GND.n2180 GND.n2178 585
R1736 GND.n2178 GND.n2174 585
R1737 GND.n3597 GND.n3596 585
R1738 GND.n3598 GND.n3597 585
R1739 GND.n2162 GND.n2161 585
R1740 GND.n2166 GND.n2162 585
R1741 GND.n4554 GND.n4553 585
R1742 GND.n4553 GND.n4552 585
R1743 GND.n4555 GND.n2159 585
R1744 GND.n3578 GND.n2159 585
R1745 GND.n4557 GND.n4556 585
R1746 GND.n4558 GND.n4557 585
R1747 GND.n2160 GND.n2158 585
R1748 GND.n2158 GND.n2154 585
R1749 GND.n3158 GND.n3157 585
R1750 GND.n3159 GND.n3158 585
R1751 GND.n2142 GND.n2141 585
R1752 GND.n2146 GND.n2142 585
R1753 GND.n4568 GND.n4567 585
R1754 GND.n4567 GND.n4566 585
R1755 GND.n4569 GND.n2139 585
R1756 GND.n3564 GND.n2139 585
R1757 GND.n4571 GND.n4570 585
R1758 GND.n4572 GND.n4571 585
R1759 GND.n2140 GND.n2138 585
R1760 GND.n2138 GND.n2134 585
R1761 GND.n3525 GND.n3524 585
R1762 GND.n3526 GND.n3525 585
R1763 GND.n2122 GND.n2121 585
R1764 GND.n2126 GND.n2122 585
R1765 GND.n4582 GND.n4581 585
R1766 GND.n4581 GND.n4580 585
R1767 GND.n4583 GND.n2119 585
R1768 GND.n3516 GND.n2119 585
R1769 GND.n4585 GND.n4584 585
R1770 GND.n4586 GND.n4585 585
R1771 GND.n2120 GND.n2118 585
R1772 GND.n3506 GND.n2118 585
R1773 GND.n3492 GND.n3491 585
R1774 GND.n3492 GND.n3186 585
R1775 GND.n3494 GND.n3493 585
R1776 GND.n3493 GND.n2101 585
R1777 GND.n3495 GND.n3490 585
R1778 GND.n3490 GND.n2099 585
R1779 GND.n3497 GND.n3496 585
R1780 GND.n3498 GND.n3497 585
R1781 GND.n2087 GND.n2086 585
R1782 GND.n3191 GND.n2087 585
R1783 GND.n4603 GND.n4602 585
R1784 GND.n4602 GND.n4601 585
R1785 GND.n4604 GND.n2084 585
R1786 GND.n3462 GND.n2084 585
R1787 GND.n4606 GND.n4605 585
R1788 GND.n4607 GND.n4606 585
R1789 GND.n2085 GND.n2083 585
R1790 GND.n3477 GND.n2083 585
R1791 GND.n2068 GND.n2067 585
R1792 GND.n3286 GND.n2068 585
R1793 GND.n4618 GND.n4617 585
R1794 GND.n4617 GND.n4616 585
R1795 GND.n4619 GND.n2065 585
R1796 GND.n3455 GND.n2065 585
R1797 GND.n4621 GND.n4620 585
R1798 GND.n4622 GND.n4621 585
R1799 GND.n2066 GND.n2064 585
R1800 GND.n2064 GND.n2061 585
R1801 GND.n3335 GND.n3334 585
R1802 GND.n3338 GND.n3337 585
R1803 GND.n3339 GND.n3322 585
R1804 GND.n3322 GND.n2053 585
R1805 GND.n3341 GND.n3340 585
R1806 GND.n3343 GND.n3321 585
R1807 GND.n3346 GND.n3345 585
R1808 GND.n3347 GND.n3320 585
R1809 GND.n3349 GND.n3348 585
R1810 GND.n3351 GND.n3319 585
R1811 GND.n3354 GND.n3353 585
R1812 GND.n3355 GND.n3318 585
R1813 GND.n3357 GND.n3356 585
R1814 GND.n3359 GND.n3317 585
R1815 GND.n3362 GND.n3361 585
R1816 GND.n3363 GND.n3316 585
R1817 GND.n3365 GND.n3364 585
R1818 GND.n3367 GND.n3315 585
R1819 GND.n3370 GND.n3369 585
R1820 GND.n3371 GND.n3314 585
R1821 GND.n3373 GND.n3372 585
R1822 GND.n3375 GND.n3313 585
R1823 GND.n3378 GND.n3377 585
R1824 GND.n3379 GND.n3312 585
R1825 GND.n3381 GND.n3380 585
R1826 GND.n3383 GND.n3311 585
R1827 GND.n3386 GND.n3385 585
R1828 GND.n3387 GND.n3307 585
R1829 GND.n3389 GND.n3388 585
R1830 GND.n3391 GND.n3306 585
R1831 GND.n3392 GND.n1190 585
R1832 GND.n3394 GND.n1190 585
R1833 GND.n3397 GND.n3396 585
R1834 GND.n3398 GND.n3305 585
R1835 GND.n3400 GND.n3399 585
R1836 GND.n3402 GND.n3304 585
R1837 GND.n3405 GND.n3404 585
R1838 GND.n3406 GND.n3300 585
R1839 GND.n3408 GND.n3407 585
R1840 GND.n3410 GND.n3299 585
R1841 GND.n3413 GND.n3412 585
R1842 GND.n3414 GND.n3298 585
R1843 GND.n3416 GND.n3415 585
R1844 GND.n3418 GND.n3297 585
R1845 GND.n3421 GND.n3420 585
R1846 GND.n3422 GND.n3296 585
R1847 GND.n3424 GND.n3423 585
R1848 GND.n3426 GND.n3295 585
R1849 GND.n3429 GND.n3428 585
R1850 GND.n3430 GND.n3294 585
R1851 GND.n3432 GND.n3431 585
R1852 GND.n3434 GND.n3293 585
R1853 GND.n3437 GND.n3436 585
R1854 GND.n3438 GND.n3292 585
R1855 GND.n3440 GND.n3439 585
R1856 GND.n3442 GND.n3291 585
R1857 GND.n3445 GND.n3444 585
R1858 GND.n3446 GND.n3290 585
R1859 GND.n3448 GND.n3447 585
R1860 GND.n3450 GND.n3289 585
R1861 GND.n3451 GND.n3288 585
R1862 GND.n3451 GND.n2053 585
R1863 GND.n3897 GND.n3896 585
R1864 GND.n3899 GND.n3087 585
R1865 GND.n3901 GND.n3900 585
R1866 GND.n3902 GND.n3086 585
R1867 GND.n3904 GND.n3903 585
R1868 GND.n3906 GND.n3084 585
R1869 GND.n3908 GND.n3907 585
R1870 GND.n3909 GND.n3083 585
R1871 GND.n3911 GND.n3910 585
R1872 GND.n3913 GND.n3081 585
R1873 GND.n3915 GND.n3914 585
R1874 GND.n3916 GND.n3080 585
R1875 GND.n3918 GND.n3917 585
R1876 GND.n3920 GND.n3078 585
R1877 GND.n3922 GND.n3921 585
R1878 GND.n3923 GND.n3077 585
R1879 GND.n3925 GND.n3924 585
R1880 GND.n3927 GND.n3075 585
R1881 GND.n3929 GND.n3928 585
R1882 GND.n3930 GND.n3074 585
R1883 GND.n3932 GND.n3931 585
R1884 GND.n3934 GND.n3072 585
R1885 GND.n3936 GND.n3935 585
R1886 GND.n3937 GND.n3068 585
R1887 GND.n3939 GND.n3938 585
R1888 GND.n3941 GND.n3066 585
R1889 GND.n3943 GND.n3942 585
R1890 GND.n3944 GND.n3065 585
R1891 GND.n3946 GND.n3945 585
R1892 GND.n3951 GND.n3950 585
R1893 GND.n3953 GND.n3952 585
R1894 GND.n3955 GND.n3063 585
R1895 GND.n3957 GND.n3956 585
R1896 GND.n3959 GND.n3060 585
R1897 GND.n3961 GND.n3960 585
R1898 GND.n3963 GND.n3058 585
R1899 GND.n3965 GND.n3964 585
R1900 GND.n3966 GND.n3057 585
R1901 GND.n3968 GND.n3967 585
R1902 GND.n3970 GND.n3055 585
R1903 GND.n3972 GND.n3971 585
R1904 GND.n3973 GND.n3054 585
R1905 GND.n3975 GND.n3974 585
R1906 GND.n3977 GND.n3052 585
R1907 GND.n3979 GND.n3978 585
R1908 GND.n3980 GND.n3051 585
R1909 GND.n3982 GND.n3981 585
R1910 GND.n3984 GND.n3049 585
R1911 GND.n3986 GND.n3985 585
R1912 GND.n3987 GND.n3048 585
R1913 GND.n3989 GND.n3988 585
R1914 GND.n3991 GND.n3046 585
R1915 GND.n3993 GND.n3992 585
R1916 GND.n3994 GND.n3045 585
R1917 GND.n3996 GND.n3995 585
R1918 GND.n3998 GND.n3043 585
R1919 GND.n4000 GND.n3999 585
R1920 GND.n4001 GND.n3032 585
R1921 GND.n3895 GND.n3029 585
R1922 GND.n4005 GND.n3029 585
R1923 GND.n3894 GND.n3893 585
R1924 GND.n3893 GND.n3028 585
R1925 GND.n3892 GND.n3089 585
R1926 GND.n3892 GND.n3891 585
R1927 GND.n3786 GND.n2368 585
R1928 GND.n4434 GND.n2368 585
R1929 GND.n3789 GND.n3788 585
R1930 GND.n3788 GND.n3787 585
R1931 GND.n3790 GND.n2360 585
R1932 GND.n4440 GND.n2360 585
R1933 GND.n3792 GND.n3791 585
R1934 GND.n3793 GND.n3792 585
R1935 GND.n3785 GND.n3097 585
R1936 GND.n3773 GND.n3097 585
R1937 GND.n3784 GND.n3783 585
R1938 GND.n3783 GND.n2346 585
R1939 GND.n3782 GND.n3098 585
R1940 GND.n3782 GND.n2344 585
R1941 GND.n3781 GND.n3100 585
R1942 GND.n3781 GND.n3780 585
R1943 GND.n3725 GND.n3099 585
R1944 GND.n3101 GND.n3099 585
R1945 GND.n3726 GND.n2325 585
R1946 GND.n4455 GND.n2325 585
R1947 GND.n3729 GND.n3728 585
R1948 GND.n3728 GND.n3727 585
R1949 GND.n3730 GND.n2317 585
R1950 GND.n4461 GND.n2317 585
R1951 GND.n3732 GND.n3731 585
R1952 GND.n3733 GND.n3732 585
R1953 GND.n3737 GND.n3736 585
R1954 GND.n3736 GND.n3735 585
R1955 GND.n3738 GND.n2301 585
R1956 GND.n4469 GND.n2301 585
R1957 GND.n3742 GND.n3741 585
R1958 GND.n3741 GND.n3740 585
R1959 GND.n3743 GND.n2294 585
R1960 GND.n4475 GND.n2294 585
R1961 GND.n3745 GND.n3744 585
R1962 GND.n3746 GND.n3745 585
R1963 GND.n3724 GND.n3111 585
R1964 GND.n3111 GND.n3110 585
R1965 GND.n3723 GND.n3722 585
R1966 GND.n3722 GND.n2278 585
R1967 GND.n3721 GND.n3112 585
R1968 GND.n3721 GND.n2276 585
R1969 GND.n3720 GND.n3114 585
R1970 GND.n3720 GND.n3719 585
R1971 GND.n3689 GND.n3113 585
R1972 GND.n3115 GND.n3113 585
R1973 GND.n3690 GND.n2258 585
R1974 GND.n4490 GND.n2258 585
R1975 GND.n3693 GND.n3692 585
R1976 GND.n3692 GND.n3691 585
R1977 GND.n3694 GND.n2249 585
R1978 GND.n4496 GND.n2249 585
R1979 GND.n3696 GND.n3695 585
R1980 GND.n3697 GND.n3696 585
R1981 GND.n3688 GND.n3123 585
R1982 GND.n3123 GND.n3122 585
R1983 GND.n3687 GND.n2232 585
R1984 GND.n4503 GND.n2232 585
R1985 GND.n3686 GND.n3685 585
R1986 GND.n3685 GND.n3684 585
R1987 GND.n3683 GND.n2224 585
R1988 GND.n4509 GND.n2224 585
R1989 GND.n3682 GND.n3681 585
R1990 GND.n3681 GND.n3680 585
R1991 GND.n3125 GND.n3124 585
R1992 GND.n3678 GND.n3125 585
R1993 GND.n3666 GND.n3665 585
R1994 GND.n3665 GND.n2214 585
R1995 GND.n3667 GND.n3132 585
R1996 GND.n3132 GND.n2212 585
R1997 GND.n3669 GND.n3668 585
R1998 GND.n3671 GND.n3669 585
R1999 GND.n3664 GND.n3131 585
R2000 GND.n3131 GND.n3130 585
R2001 GND.n3663 GND.n2202 585
R2002 GND.n4524 GND.n2202 585
R2003 GND.n3662 GND.n3661 585
R2004 GND.n3661 GND.n3660 585
R2005 GND.n3133 GND.n2194 585
R2006 GND.n4530 GND.n2194 585
R2007 GND.n3604 GND.n3603 585
R2008 GND.n3603 GND.n2192 585
R2009 GND.n3605 GND.n3138 585
R2010 GND.n3633 GND.n3138 585
R2011 GND.n3608 GND.n3607 585
R2012 GND.n3607 GND.n3606 585
R2013 GND.n3609 GND.n2183 585
R2014 GND.n4538 GND.n2183 585
R2015 GND.n3611 GND.n3610 585
R2016 GND.n3612 GND.n3611 585
R2017 GND.n3602 GND.n2176 585
R2018 GND.n4544 GND.n2176 585
R2019 GND.n3601 GND.n3600 585
R2020 GND.n3600 GND.n2174 585
R2021 GND.n3599 GND.n3146 585
R2022 GND.n3599 GND.n3598 585
R2023 GND.n3574 GND.n3147 585
R2024 GND.n3147 GND.n2166 585
R2025 GND.n3575 GND.n2164 585
R2026 GND.n4552 GND.n2164 585
R2027 GND.n3577 GND.n3576 585
R2028 GND.n3578 GND.n3577 585
R2029 GND.n3573 GND.n2156 585
R2030 GND.n4558 GND.n2156 585
R2031 GND.n3572 GND.n3571 585
R2032 GND.n3571 GND.n2154 585
R2033 GND.n3570 GND.n3174 585
R2034 GND.n3570 GND.n3159 585
R2035 GND.n3569 GND.n3568 585
R2036 GND.n3569 GND.n2146 585
R2037 GND.n3567 GND.n2144 585
R2038 GND.n4566 GND.n2144 585
R2039 GND.n3566 GND.n3565 585
R2040 GND.n3565 GND.n3564 585
R2041 GND.n3175 GND.n2136 585
R2042 GND.n4572 GND.n2136 585
R2043 GND.n3521 GND.n3180 585
R2044 GND.n3180 GND.n2134 585
R2045 GND.n3523 GND.n3522 585
R2046 GND.n3526 GND.n3523 585
R2047 GND.n3520 GND.n3179 585
R2048 GND.n3179 GND.n2126 585
R2049 GND.n3519 GND.n2124 585
R2050 GND.n4580 GND.n2124 585
R2051 GND.n3518 GND.n3517 585
R2052 GND.n3517 GND.n3516 585
R2053 GND.n3181 GND.n2116 585
R2054 GND.n4586 GND.n2116 585
R2055 GND.n3505 GND.n3504 585
R2056 GND.n3506 GND.n3505 585
R2057 GND.n3503 GND.n3187 585
R2058 GND.n3187 GND.n3186 585
R2059 GND.n3502 GND.n3501 585
R2060 GND.n3501 GND.n2101 585
R2061 GND.n3500 GND.n3188 585
R2062 GND.n3500 GND.n2099 585
R2063 GND.n3499 GND.n3190 585
R2064 GND.n3499 GND.n3498 585
R2065 GND.n3460 GND.n3189 585
R2066 GND.n3191 GND.n3189 585
R2067 GND.n3461 GND.n2089 585
R2068 GND.n4601 GND.n2089 585
R2069 GND.n3464 GND.n3463 585
R2070 GND.n3463 GND.n3462 585
R2071 GND.n3465 GND.n2081 585
R2072 GND.n4607 GND.n2081 585
R2073 GND.n3467 GND.n3466 585
R2074 GND.n3477 GND.n3467 585
R2075 GND.n3459 GND.n3287 585
R2076 GND.n3287 GND.n3286 585
R2077 GND.n3458 GND.n2070 585
R2078 GND.n4616 GND.n2070 585
R2079 GND.n3457 GND.n3456 585
R2080 GND.n3456 GND.n3455 585
R2081 GND.n3454 GND.n2062 585
R2082 GND.n4622 GND.n2062 585
R2083 GND.n3453 GND.n3452 585
R2084 GND.n3452 GND.n2061 585
R2085 GND.n4863 GND.n905 585
R2086 GND.n905 GND.n904 585
R2087 GND.n5679 GND.n374 585
R2088 GND.n5683 GND.n374 585
R2089 GND.n5686 GND.n5685 585
R2090 GND.n5685 GND.n5684 585
R2091 GND.n5687 GND.n369 585
R2092 GND.n369 GND.n368 585
R2093 GND.n5689 GND.n5688 585
R2094 GND.n5690 GND.n5689 585
R2095 GND.n367 GND.n366 585
R2096 GND.n5691 GND.n367 585
R2097 GND.n5694 GND.n5693 585
R2098 GND.n5693 GND.n5692 585
R2099 GND.n5695 GND.n361 585
R2100 GND.n361 GND.n360 585
R2101 GND.n5697 GND.n5696 585
R2102 GND.n5698 GND.n5697 585
R2103 GND.n359 GND.n358 585
R2104 GND.n5699 GND.n359 585
R2105 GND.n5702 GND.n5701 585
R2106 GND.n5701 GND.n5700 585
R2107 GND.n5703 GND.n353 585
R2108 GND.n353 GND.n352 585
R2109 GND.n5705 GND.n5704 585
R2110 GND.n5706 GND.n5705 585
R2111 GND.n351 GND.n350 585
R2112 GND.n5707 GND.n351 585
R2113 GND.n5710 GND.n5709 585
R2114 GND.n5709 GND.n5708 585
R2115 GND.n5711 GND.n345 585
R2116 GND.n345 GND.n344 585
R2117 GND.n5713 GND.n5712 585
R2118 GND.n5714 GND.n5713 585
R2119 GND.n343 GND.n342 585
R2120 GND.n5715 GND.n343 585
R2121 GND.n5718 GND.n5717 585
R2122 GND.n5717 GND.n5716 585
R2123 GND.n5719 GND.n337 585
R2124 GND.n337 GND.n336 585
R2125 GND.n5721 GND.n5720 585
R2126 GND.n5722 GND.n5721 585
R2127 GND.n335 GND.n334 585
R2128 GND.n5723 GND.n335 585
R2129 GND.n5726 GND.n5725 585
R2130 GND.n5725 GND.n5724 585
R2131 GND.n5727 GND.n329 585
R2132 GND.n329 GND.n328 585
R2133 GND.n5729 GND.n5728 585
R2134 GND.n5730 GND.n5729 585
R2135 GND.n327 GND.n326 585
R2136 GND.n5731 GND.n327 585
R2137 GND.n5734 GND.n5733 585
R2138 GND.n5733 GND.n5732 585
R2139 GND.n5735 GND.n319 585
R2140 GND.n319 GND.n318 585
R2141 GND.n5737 GND.n5736 585
R2142 GND.n5738 GND.n5737 585
R2143 GND.n320 GND.n317 585
R2144 GND.n5739 GND.n317 585
R2145 GND.n5741 GND.n316 585
R2146 GND.n5741 GND.n5740 585
R2147 GND.n5743 GND.n5742 585
R2148 GND.n5742 GND.n278 585
R2149 GND.n5744 GND.n311 585
R2150 GND.n311 GND.n272 585
R2151 GND.n5746 GND.n5745 585
R2152 GND.n5747 GND.n5746 585
R2153 GND.n312 GND.n310 585
R2154 GND.n310 GND.n265 585
R2155 GND.n4275 GND.n4270 585
R2156 GND.n4270 GND.n262 585
R2157 GND.n4277 GND.n4276 585
R2158 GND.n4277 GND.n255 585
R2159 GND.n4278 GND.n4269 585
R2160 GND.n4278 GND.n252 585
R2161 GND.n4280 GND.n4279 585
R2162 GND.n4279 GND.n244 585
R2163 GND.n4281 GND.n4264 585
R2164 GND.n4264 GND.n4263 585
R2165 GND.n4283 GND.n4282 585
R2166 GND.n4283 GND.n235 585
R2167 GND.n4284 GND.n2955 585
R2168 GND.n4284 GND.n232 585
R2169 GND.n4286 GND.n4285 585
R2170 GND.n4285 GND.n224 585
R2171 GND.n4287 GND.n2950 585
R2172 GND.n2950 GND.n221 585
R2173 GND.n4289 GND.n4288 585
R2174 GND.n4289 GND.n214 585
R2175 GND.n4290 GND.n2949 585
R2176 GND.n4290 GND.n211 585
R2177 GND.n4292 GND.n4291 585
R2178 GND.n4291 GND.n203 585
R2179 GND.n4293 GND.n2944 585
R2180 GND.n2944 GND.n200 585
R2181 GND.n4295 GND.n4294 585
R2182 GND.n4295 GND.n193 585
R2183 GND.n4296 GND.n2943 585
R2184 GND.n4296 GND.n190 585
R2185 GND.n4298 GND.n4297 585
R2186 GND.n4297 GND.n183 585
R2187 GND.n4299 GND.n2940 585
R2188 GND.n2940 GND.n180 585
R2189 GND.n4301 GND.n4300 585
R2190 GND.n4301 GND.n171 585
R2191 GND.n4303 GND.n4302 585
R2192 GND.n4302 GND.n168 585
R2193 GND.n4304 GND.n2933 585
R2194 GND.n4158 GND.n2933 585
R2195 GND.n4307 GND.n4306 585
R2196 GND.n4308 GND.n4307 585
R2197 GND.n2938 GND.n2932 585
R2198 GND.n2932 GND.n151 585
R2199 GND.n2936 GND.n2935 585
R2200 GND.n2935 GND.n149 585
R2201 GND.n2934 GND.n2913 585
R2202 GND.n2918 GND.n2913 585
R2203 GND.n4322 GND.n4321 585
R2204 GND.n4321 GND.n4320 585
R2205 GND.n4323 GND.n2910 585
R2206 GND.n2914 GND.n2910 585
R2207 GND.n4326 GND.n4325 585
R2208 GND.n4327 GND.n4326 585
R2209 GND.n2911 GND.n2909 585
R2210 GND.n2909 GND.n2905 585
R2211 GND.n4058 GND.n4057 585
R2212 GND.n4058 GND.n2900 585
R2213 GND.n4059 GND.n4053 585
R2214 GND.n4059 GND.n2893 585
R2215 GND.n4061 GND.n4060 585
R2216 GND.n4060 GND.n2890 585
R2217 GND.n4062 GND.n4048 585
R2218 GND.n4048 GND.n2881 585
R2219 GND.n4064 GND.n4063 585
R2220 GND.n4064 GND.n2878 585
R2221 GND.n4065 GND.n4047 585
R2222 GND.n4065 GND.n2871 585
R2223 GND.n4067 GND.n4066 585
R2224 GND.n4066 GND.n2868 585
R2225 GND.n4068 GND.n4042 585
R2226 GND.n4042 GND.n2860 585
R2227 GND.n4070 GND.n4069 585
R2228 GND.n4070 GND.n2857 585
R2229 GND.n4071 GND.n4041 585
R2230 GND.n4071 GND.n2850 585
R2231 GND.n4073 GND.n4072 585
R2232 GND.n4072 GND.n2847 585
R2233 GND.n4074 GND.n3008 585
R2234 GND.n3008 GND.n2839 585
R2235 GND.n4076 GND.n4075 585
R2236 GND.n4077 GND.n4076 585
R2237 GND.n3009 GND.n3007 585
R2238 GND.n3007 GND.n2827 585
R2239 GND.n4035 GND.n4034 585
R2240 GND.n4034 GND.n2824 585
R2241 GND.n4033 GND.n3011 585
R2242 GND.n4033 GND.n2811 585
R2243 GND.n4032 GND.n4031 585
R2244 GND.n4032 GND.n2809 585
R2245 GND.n3013 GND.n3012 585
R2246 GND.n3012 GND.n2427 585
R2247 GND.n4027 GND.n4026 585
R2248 GND.n4026 GND.n2426 585
R2249 GND.n4025 GND.n3015 585
R2250 GND.n4025 GND.n2395 585
R2251 GND.n4024 GND.n4023 585
R2252 GND.n4024 GND.n2382 585
R2253 GND.n3017 GND.n3016 585
R2254 GND.n4016 GND.n3016 585
R2255 GND.n4019 GND.n4018 585
R2256 GND.n4018 GND.n4017 585
R2257 GND.n3020 GND.n3019 585
R2258 GND.n4015 GND.n3020 585
R2259 GND.n4013 GND.n4012 585
R2260 GND.n4014 GND.n4013 585
R2261 GND.n3023 GND.n3022 585
R2262 GND.n3030 GND.n3022 585
R2263 GND.n4008 GND.n4007 585
R2264 GND.n4007 GND.n4006 585
R2265 GND.n3027 GND.n3026 585
R2266 GND.n3090 GND.n3027 585
R2267 GND.n2359 GND.n2358 585
R2268 GND.n2367 GND.n2359 585
R2269 GND.n4443 GND.n4442 585
R2270 GND.n4442 GND.n4441 585
R2271 GND.n4444 GND.n2348 585
R2272 GND.n3096 GND.n2348 585
R2273 GND.n4446 GND.n4445 585
R2274 GND.n4447 GND.n4446 585
R2275 GND.n2349 GND.n2347 585
R2276 GND.n3769 GND.n2347 585
R2277 GND.n2352 GND.n2351 585
R2278 GND.n2351 GND.n2327 585
R2279 GND.n2315 GND.n2314 585
R2280 GND.n2324 GND.n2315 585
R2281 GND.n4464 GND.n4463 585
R2282 GND.n4463 GND.n4462 585
R2283 GND.n4465 GND.n2304 585
R2284 GND.n3734 GND.n2304 585
R2285 GND.n4467 GND.n4466 585
R2286 GND.n4468 GND.n4467 585
R2287 GND.n2305 GND.n2303 585
R2288 GND.n3739 GND.n2303 585
R2289 GND.n2308 GND.n2307 585
R2290 GND.n2307 GND.n2292 585
R2291 GND.n2275 GND.n2274 585
R2292 GND.n3109 GND.n2275 585
R2293 GND.n4485 GND.n4484 585
R2294 GND.n4484 GND.n4483 585
R2295 GND.n4486 GND.n2261 585
R2296 GND.n3116 GND.n2261 585
R2297 GND.n4488 GND.n4487 585
R2298 GND.n4489 GND.n4488 585
R2299 GND.n2262 GND.n2260 585
R2300 GND.n2260 GND.n2251 585
R2301 GND.n2268 GND.n2267 585
R2302 GND.n2267 GND.n2248 585
R2303 GND.n2266 GND.n2265 585
R2304 GND.n2266 GND.n2234 585
R2305 GND.n2222 GND.n2221 585
R2306 GND.n2231 GND.n2222 585
R2307 GND.n4512 GND.n4511 585
R2308 GND.n4511 GND.n4510 585
R2309 GND.n4513 GND.n2216 585
R2310 GND.n3679 GND.n2216 585
R2311 GND.n4515 GND.n4514 585
R2312 GND.n4516 GND.n4515 585
R2313 GND.n2217 GND.n2215 585
R2314 GND.n3670 GND.n2215 585
R2315 GND.n3624 GND.n3623 585
R2316 GND.n3624 GND.n2204 585
R2317 GND.n3626 GND.n3625 585
R2318 GND.n3625 GND.n2201 585
R2319 GND.n3627 GND.n3140 585
R2320 GND.n3140 GND.n2195 585
R2321 GND.n3629 GND.n3628 585
R2322 GND.n3630 GND.n3629 585
R2323 GND.n3141 GND.n3139 585
R2324 GND.n3139 GND.n3137 585
R2325 GND.n3615 GND.n3614 585
R2326 GND.n3614 GND.n3613 585
R2327 GND.n3144 GND.n3143 585
R2328 GND.n3144 GND.n2177 585
R2329 GND.n3594 GND.n3593 585
R2330 GND.n3595 GND.n3594 585
R2331 GND.n3151 GND.n3150 585
R2332 GND.n3150 GND.n3149 585
R2333 GND.n3589 GND.n3588 585
R2334 GND.n3588 GND.n2163 585
R2335 GND.n3587 GND.n3153 585
R2336 GND.n3587 GND.n2157 585
R2337 GND.n3586 GND.n3155 585
R2338 GND.n3586 GND.n3585 585
R2339 GND.n3547 GND.n3154 585
R2340 GND.n3156 GND.n3154 585
R2341 GND.n3549 GND.n3548 585
R2342 GND.n3548 GND.n2143 585
R2343 GND.n3550 GND.n3529 585
R2344 GND.n3529 GND.n2137 585
R2345 GND.n3552 GND.n3551 585
R2346 GND.n3553 GND.n3552 585
R2347 GND.n3530 GND.n3528 585
R2348 GND.n3528 GND.n3527 585
R2349 GND.n3539 GND.n3538 585
R2350 GND.n3538 GND.n2123 585
R2351 GND.n3537 GND.n3532 585
R2352 GND.n3537 GND.n2117 585
R2353 GND.n3536 GND.n3535 585
R2354 GND.n3536 GND.n2114 585
R2355 GND.n2098 GND.n2097 585
R2356 GND.n3185 GND.n2098 585
R2357 GND.n4596 GND.n4595 585
R2358 GND.n4595 GND.n4594 585
R2359 GND.n4597 GND.n2092 585
R2360 GND.n3192 GND.n2092 585
R2361 GND.n4599 GND.n4598 585
R2362 GND.n4600 GND.n4599 585
R2363 GND.n2093 GND.n2091 585
R2364 GND.n2091 GND.n2082 585
R2365 GND.n3475 GND.n3474 585
R2366 GND.n3476 GND.n3475 585
R2367 GND.n3469 GND.n3468 585
R2368 GND.n3468 GND.n2072 585
R2369 GND.n2060 GND.n2059 585
R2370 GND.n2069 GND.n2060 585
R2371 GND.n4625 GND.n4624 585
R2372 GND.n4624 GND.n4623 585
R2373 GND.n4626 GND.n2054 585
R2374 GND.n3209 GND.n2054 585
R2375 GND.n4628 GND.n4627 585
R2376 GND.n4629 GND.n4628 585
R2377 GND.n2052 GND.n2051 585
R2378 GND.n4630 GND.n2052 585
R2379 GND.n4633 GND.n4632 585
R2380 GND.n4632 GND.n4631 585
R2381 GND.n4634 GND.n1486 585
R2382 GND.n1486 GND.n1484 585
R2383 GND.n4636 GND.n4635 585
R2384 GND.n4637 GND.n4636 585
R2385 GND.n1487 GND.n1485 585
R2386 GND.n1485 GND.n1478 585
R2387 GND.n2045 GND.n2044 585
R2388 GND.n2044 GND.n1172 585
R2389 GND.n2043 GND.n1489 585
R2390 GND.n2043 GND.n1170 585
R2391 GND.n2042 GND.n1491 585
R2392 GND.n2042 GND.n2041 585
R2393 GND.n1642 GND.n1490 585
R2394 GND.n1499 GND.n1490 585
R2395 GND.n1644 GND.n1643 585
R2396 GND.n1643 GND.n1497 585
R2397 GND.n1645 GND.n1635 585
R2398 GND.n1635 GND.n1508 585
R2399 GND.n1647 GND.n1646 585
R2400 GND.n1647 GND.n1506 585
R2401 GND.n1648 GND.n1634 585
R2402 GND.n1648 GND.n1510 585
R2403 GND.n1650 GND.n1649 585
R2404 GND.n1649 GND.n1519 585
R2405 GND.n1651 GND.n1629 585
R2406 GND.n1629 GND.n1518 585
R2407 GND.n1653 GND.n1652 585
R2408 GND.n1653 GND.n1532 585
R2409 GND.n1654 GND.n1628 585
R2410 GND.n1654 GND.n1529 585
R2411 GND.n1656 GND.n1655 585
R2412 GND.n1655 GND.n1535 585
R2413 GND.n1657 GND.n1623 585
R2414 GND.n1623 GND.n1543 585
R2415 GND.n1659 GND.n1658 585
R2416 GND.n1659 GND.n1542 585
R2417 GND.n1660 GND.n1622 585
R2418 GND.n1660 GND.n1554 585
R2419 GND.n1662 GND.n1661 585
R2420 GND.n1661 GND.n1552 585
R2421 GND.n1663 GND.n1617 585
R2422 GND.n1617 GND.n1557 585
R2423 GND.n1665 GND.n1664 585
R2424 GND.n1665 GND.n1565 585
R2425 GND.n1666 GND.n1616 585
R2426 GND.n1909 GND.n1666 585
R2427 GND.n1916 GND.n1915 585
R2428 GND.n1915 GND.n1914 585
R2429 GND.n1918 GND.n1612 585
R2430 GND.n1667 GND.n1612 585
R2431 GND.n1920 GND.n1919 585
R2432 GND.n1921 GND.n1920 585
R2433 GND.n1614 GND.n1611 585
R2434 GND.n1611 GND.n1606 585
R2435 GND.n1613 GND.n1593 585
R2436 GND.n1597 GND.n1593 585
R2437 GND.n1933 GND.n1932 585
R2438 GND.n1932 GND.n1931 585
R2439 GND.n1934 GND.n1590 585
R2440 GND.n1594 GND.n1590 585
R2441 GND.n1937 GND.n1936 585
R2442 GND.n1938 GND.n1937 585
R2443 GND.n1591 GND.n1589 585
R2444 GND.n1589 GND.n1583 585
R2445 GND.n1797 GND.n1793 585
R2446 GND.n1793 GND.n1581 585
R2447 GND.n1799 GND.n1798 585
R2448 GND.n1799 GND.n1681 585
R2449 GND.n1800 GND.n1792 585
R2450 GND.n1800 GND.n1678 585
R2451 GND.n1802 GND.n1801 585
R2452 GND.n1801 GND.n1690 585
R2453 GND.n1803 GND.n1787 585
R2454 GND.n1787 GND.n1688 585
R2455 GND.n1805 GND.n1804 585
R2456 GND.n1805 GND.n1692 585
R2457 GND.n1806 GND.n1786 585
R2458 GND.n1806 GND.n1700 585
R2459 GND.n1808 GND.n1807 585
R2460 GND.n1807 GND.n1699 585
R2461 GND.n1809 GND.n1781 585
R2462 GND.n1781 GND.n1712 585
R2463 GND.n1811 GND.n1810 585
R2464 GND.n1811 GND.n1710 585
R2465 GND.n1812 GND.n1780 585
R2466 GND.n1812 GND.n1714 585
R2467 GND.n1814 GND.n1813 585
R2468 GND.n1813 GND.n1723 585
R2469 GND.n1815 GND.n1739 585
R2470 GND.n1739 GND.n1722 585
R2471 GND.n1817 GND.n1816 585
R2472 GND.n1818 GND.n1817 585
R2473 GND.n1740 GND.n1738 585
R2474 GND.n1738 GND.n1734 585
R2475 GND.n1774 GND.n1773 585
R2476 GND.n1773 GND.n1772 585
R2477 GND.n1756 GND.n1742 585
R2478 GND.n1756 GND.n1007 585
R2479 GND.n1755 GND.n1754 585
R2480 GND.n1755 GND.n1004 585
R2481 GND.n1744 GND.n1743 585
R2482 GND.n1743 GND.n996 585
R2483 GND.n1750 GND.n1749 585
R2484 GND.n1749 GND.n994 585
R2485 GND.n1748 GND.n1747 585
R2486 GND.n1748 GND.n980 585
R2487 GND.n965 GND.n964 585
R2488 GND.n4801 GND.n965 585
R2489 GND.n4804 GND.n4803 585
R2490 GND.n4803 GND.n4802 585
R2491 GND.n4805 GND.n959 585
R2492 GND.n959 GND.n958 585
R2493 GND.n4807 GND.n4806 585
R2494 GND.n4808 GND.n4807 585
R2495 GND.n957 GND.n956 585
R2496 GND.n4809 GND.n957 585
R2497 GND.n4812 GND.n4811 585
R2498 GND.n4811 GND.n4810 585
R2499 GND.n4813 GND.n951 585
R2500 GND.n951 GND.n950 585
R2501 GND.n4815 GND.n4814 585
R2502 GND.n4816 GND.n4815 585
R2503 GND.n949 GND.n948 585
R2504 GND.n4817 GND.n949 585
R2505 GND.n4820 GND.n4819 585
R2506 GND.n4819 GND.n4818 585
R2507 GND.n4821 GND.n943 585
R2508 GND.n943 GND.n942 585
R2509 GND.n4823 GND.n4822 585
R2510 GND.n4824 GND.n4823 585
R2511 GND.n941 GND.n940 585
R2512 GND.n4825 GND.n941 585
R2513 GND.n4828 GND.n4827 585
R2514 GND.n4827 GND.n4826 585
R2515 GND.n4829 GND.n935 585
R2516 GND.n935 GND.n934 585
R2517 GND.n4831 GND.n4830 585
R2518 GND.n4832 GND.n4831 585
R2519 GND.n933 GND.n932 585
R2520 GND.n4833 GND.n933 585
R2521 GND.n4836 GND.n4835 585
R2522 GND.n4835 GND.n4834 585
R2523 GND.n4837 GND.n927 585
R2524 GND.n927 GND.n926 585
R2525 GND.n4839 GND.n4838 585
R2526 GND.n4840 GND.n4839 585
R2527 GND.n925 GND.n924 585
R2528 GND.n4841 GND.n925 585
R2529 GND.n4844 GND.n4843 585
R2530 GND.n4843 GND.n4842 585
R2531 GND.n4845 GND.n919 585
R2532 GND.n919 GND.n918 585
R2533 GND.n4847 GND.n4846 585
R2534 GND.n4848 GND.n4847 585
R2535 GND.n917 GND.n916 585
R2536 GND.n4849 GND.n917 585
R2537 GND.n4852 GND.n4851 585
R2538 GND.n4851 GND.n4850 585
R2539 GND.n4853 GND.n912 585
R2540 GND.n912 GND.n911 585
R2541 GND.n4855 GND.n4854 585
R2542 GND.n4856 GND.n4855 585
R2543 GND.n910 GND.n909 585
R2544 GND.n4857 GND.n910 585
R2545 GND.n4860 GND.n4859 585
R2546 GND.n4859 GND.n4858 585
R2547 GND.n4799 GND.n4798 585
R2548 GND.n4800 GND.n4799 585
R2549 GND.n4797 GND.n982 585
R2550 GND.n986 GND.n984 585
R2551 GND.n4793 GND.n987 585
R2552 GND.n4792 GND.n988 585
R2553 GND.n4791 GND.n989 585
R2554 GND.n4783 GND.n990 585
R2555 GND.n4787 GND.n4784 585
R2556 GND.n4782 GND.n4781 585
R2557 GND.n1174 GND.n1173 585
R2558 GND.n4700 GND.n1174 585
R2559 GND.n2039 GND.n1166 585
R2560 GND.n2040 GND.n2039 585
R2561 GND.n2038 GND.n1165 585
R2562 GND.n2038 GND.n1493 585
R2563 GND.n2037 GND.n1164 585
R2564 GND.n2037 GND.n2036 585
R2565 GND.n1496 GND.n1495 585
R2566 GND.n2008 GND.n1496 585
R2567 GND.n2025 GND.n1158 585
R2568 GND.n2026 GND.n2025 585
R2569 GND.n2024 GND.n1157 585
R2570 GND.n2024 GND.n2023 585
R2571 GND.n1509 GND.n1156 585
R2572 GND.n1523 GND.n1509 585
R2573 GND.n1521 GND.n1520 585
R2574 GND.n2002 GND.n1521 585
R2575 GND.n1990 GND.n1150 585
R2576 GND.n1990 GND.n1989 585
R2577 GND.n1991 GND.n1149 585
R2578 GND.n1992 GND.n1991 585
R2579 GND.n1988 GND.n1148 585
R2580 GND.n1988 GND.n1987 585
R2581 GND.n1534 GND.n1533 585
R2582 GND.n1546 GND.n1534 585
R2583 GND.n1544 GND.n1142 585
R2584 GND.n1978 GND.n1544 585
R2585 GND.n1966 GND.n1141 585
R2586 GND.n1966 GND.n1965 585
R2587 GND.n1967 GND.n1140 585
R2588 GND.n1968 GND.n1967 585
R2589 GND.n1963 GND.n1556 585
R2590 GND.n1963 GND.n1962 585
R2591 GND.n1555 GND.n1134 585
R2592 GND.n1568 GND.n1555 585
R2593 GND.n1566 GND.n1133 585
R2594 GND.n1953 GND.n1566 585
R2595 GND.n1912 GND.n1132 585
R2596 GND.n1913 GND.n1912 585
R2597 GND.n1911 GND.n1910 585
R2598 GND.n1911 GND.n1908 585
R2599 GND.n1607 GND.n1126 585
R2600 GND.n1610 GND.n1607 585
R2601 GND.n1923 GND.n1125 585
R2602 GND.n1923 GND.n1922 585
R2603 GND.n1924 GND.n1124 585
R2604 GND.n1925 GND.n1924 585
R2605 GND.n1600 GND.n1599 585
R2606 GND.n1930 GND.n1600 585
R2607 GND.n1598 GND.n1118 585
R2608 GND.n1598 GND.n1595 585
R2609 GND.n1585 GND.n1117 585
R2610 GND.n1588 GND.n1585 585
R2611 GND.n1940 GND.n1116 585
R2612 GND.n1940 GND.n1939 585
R2613 GND.n1942 GND.n1941 585
R2614 GND.n1943 GND.n1942 585
R2615 GND.n1584 GND.n1110 585
R2616 GND.n1680 GND.n1584 585
R2617 GND.n1682 GND.n1109 585
R2618 GND.n1880 GND.n1682 585
R2619 GND.n1869 GND.n1108 585
R2620 GND.n1869 GND.n1868 585
R2621 GND.n1871 GND.n1870 585
R2622 GND.n1872 GND.n1871 585
R2623 GND.n1867 GND.n1102 585
R2624 GND.n1867 GND.n1866 585
R2625 GND.n1691 GND.n1101 585
R2626 GND.n1704 GND.n1691 585
R2627 GND.n1701 GND.n1100 585
R2628 GND.n1857 GND.n1701 585
R2629 GND.n1845 GND.n1843 585
R2630 GND.n1845 GND.n1844 585
R2631 GND.n1846 GND.n1094 585
R2632 GND.n1847 GND.n1846 585
R2633 GND.n1842 GND.n1093 585
R2634 GND.n1842 GND.n1841 585
R2635 GND.n1713 GND.n1092 585
R2636 GND.n1727 GND.n1713 585
R2637 GND.n1725 GND.n1724 585
R2638 GND.n1832 GND.n1725 585
R2639 GND.n1820 GND.n1086 585
R2640 GND.n1820 GND.n1819 585
R2641 GND.n1821 GND.n1085 585
R2642 GND.n1822 GND.n1821 585
R2643 GND.n1737 GND.n1084 585
R2644 GND.n1771 GND.n1737 585
R2645 GND.n1011 GND.n1009 585
R2646 GND.n1757 GND.n1009 585
R2647 GND.n4772 GND.n4771 585
R2648 GND.n4773 GND.n4772 585
R2649 GND.n1010 GND.n1008 585
R2650 GND.n1078 GND.n1008 585
R2651 GND.n1075 GND.n981 585
R2652 GND.n4779 GND.n981 585
R2653 GND.n4653 GND.n4652 585
R2654 GND.n4652 GND.n4651 585
R2655 GND.n1477 GND.n1473 585
R2656 GND.n4658 GND.n1470 585
R2657 GND.n4659 GND.n1469 585
R2658 GND.n4660 GND.n1468 585
R2659 GND.n1480 GND.n1209 585
R2660 GND.n4665 GND.n1208 585
R2661 GND.n4666 GND.n1207 585
R2662 GND.n4667 GND.n1206 585
R2663 GND.n2011 GND.n1171 585
R2664 GND.n4700 GND.n1171 585
R2665 GND.n2012 GND.n1494 585
R2666 GND.n2040 GND.n1494 585
R2667 GND.n2015 GND.n2010 585
R2668 GND.n2010 GND.n1493 585
R2669 GND.n2016 GND.n1498 585
R2670 GND.n2036 GND.n1498 585
R2671 GND.n2017 GND.n2009 585
R2672 GND.n2009 GND.n2008 585
R2673 GND.n1514 GND.n1507 585
R2674 GND.n2026 GND.n1507 585
R2675 GND.n2022 GND.n2021 585
R2676 GND.n2023 GND.n2022 585
R2677 GND.n1513 GND.n1512 585
R2678 GND.n1523 GND.n1512 585
R2679 GND.n2004 GND.n2003 585
R2680 GND.n2003 GND.n2002 585
R2681 GND.n1517 GND.n1516 585
R2682 GND.n1989 GND.n1517 585
R2683 GND.n1538 GND.n1531 585
R2684 GND.n1992 GND.n1531 585
R2685 GND.n1986 GND.n1985 585
R2686 GND.n1987 GND.n1986 585
R2687 GND.n1537 GND.n1536 585
R2688 GND.n1546 GND.n1536 585
R2689 GND.n1980 GND.n1979 585
R2690 GND.n1979 GND.n1978 585
R2691 GND.n1541 GND.n1540 585
R2692 GND.n1965 GND.n1541 585
R2693 GND.n1560 GND.n1553 585
R2694 GND.n1968 GND.n1553 585
R2695 GND.n1961 GND.n1960 585
R2696 GND.n1962 GND.n1961 585
R2697 GND.n1559 GND.n1558 585
R2698 GND.n1568 GND.n1558 585
R2699 GND.n1955 GND.n1954 585
R2700 GND.n1954 GND.n1953 585
R2701 GND.n1563 GND.n1562 585
R2702 GND.n1913 GND.n1563 585
R2703 GND.n1902 GND.n1901 585
R2704 GND.n1908 GND.n1902 585
R2705 GND.n1669 GND.n1668 585
R2706 GND.n1668 GND.n1610 585
R2707 GND.n1897 GND.n1609 585
R2708 GND.n1922 GND.n1609 585
R2709 GND.n1896 GND.n1605 585
R2710 GND.n1925 GND.n1605 585
R2711 GND.n1895 GND.n1596 585
R2712 GND.n1930 GND.n1596 585
R2713 GND.n1888 GND.n1671 585
R2714 GND.n1888 GND.n1595 585
R2715 GND.n1890 GND.n1889 585
R2716 GND.n1889 GND.n1588 585
R2717 GND.n1887 GND.n1586 585
R2718 GND.n1939 GND.n1586 585
R2719 GND.n1886 GND.n1582 585
R2720 GND.n1943 GND.n1582 585
R2721 GND.n1677 GND.n1673 585
R2722 GND.n1680 GND.n1677 585
R2723 GND.n1882 GND.n1881 585
R2724 GND.n1881 GND.n1880 585
R2725 GND.n1676 GND.n1675 585
R2726 GND.n1868 GND.n1676 585
R2727 GND.n1695 GND.n1689 585
R2728 GND.n1872 GND.n1689 585
R2729 GND.n1865 GND.n1864 585
R2730 GND.n1866 GND.n1865 585
R2731 GND.n1694 GND.n1693 585
R2732 GND.n1704 GND.n1693 585
R2733 GND.n1859 GND.n1858 585
R2734 GND.n1858 GND.n1857 585
R2735 GND.n1698 GND.n1697 585
R2736 GND.n1844 GND.n1698 585
R2737 GND.n1718 GND.n1711 585
R2738 GND.n1847 GND.n1711 585
R2739 GND.n1840 GND.n1839 585
R2740 GND.n1841 GND.n1840 585
R2741 GND.n1717 GND.n1716 585
R2742 GND.n1727 GND.n1716 585
R2743 GND.n1834 GND.n1833 585
R2744 GND.n1833 GND.n1832 585
R2745 GND.n1721 GND.n1720 585
R2746 GND.n1819 GND.n1721 585
R2747 GND.n1760 GND.n1736 585
R2748 GND.n1822 GND.n1736 585
R2749 GND.n1770 GND.n1769 585
R2750 GND.n1771 GND.n1770 585
R2751 GND.n1759 GND.n1758 585
R2752 GND.n1758 GND.n1757 585
R2753 GND.n1764 GND.n1006 585
R2754 GND.n4773 GND.n1006 585
R2755 GND.n1763 GND.n992 585
R2756 GND.n1078 GND.n992 585
R2757 GND.n4780 GND.n993 585
R2758 GND.n4780 GND.n4779 585
R2759 GND.n4004 GND.n3032 554.963
R2760 GND.n3897 GND.n3029 554.963
R2761 GND.n3452 GND.n3451 554.963
R2762 GND.n3335 GND.n2064 554.963
R2763 GND.n5683 GND.n5682 326.649
R2764 GND.n3326 GND.t104 314.291
R2765 GND.n3036 GND.t46 314.291
R2766 GND.n5550 GND.n453 301.784
R2767 GND.n5551 GND.n5550 301.784
R2768 GND.n5552 GND.n5551 301.784
R2769 GND.n5552 GND.n447 301.784
R2770 GND.n5560 GND.n447 301.784
R2771 GND.n5561 GND.n5560 301.784
R2772 GND.n5562 GND.n5561 301.784
R2773 GND.n5562 GND.n441 301.784
R2774 GND.n5570 GND.n441 301.784
R2775 GND.n5571 GND.n5570 301.784
R2776 GND.n5572 GND.n5571 301.784
R2777 GND.n5572 GND.n435 301.784
R2778 GND.n5580 GND.n435 301.784
R2779 GND.n5581 GND.n5580 301.784
R2780 GND.n5582 GND.n5581 301.784
R2781 GND.n5582 GND.n429 301.784
R2782 GND.n5590 GND.n429 301.784
R2783 GND.n5591 GND.n5590 301.784
R2784 GND.n5592 GND.n5591 301.784
R2785 GND.n5592 GND.n423 301.784
R2786 GND.n5600 GND.n423 301.784
R2787 GND.n5601 GND.n5600 301.784
R2788 GND.n5602 GND.n5601 301.784
R2789 GND.n5602 GND.n417 301.784
R2790 GND.n5610 GND.n417 301.784
R2791 GND.n5611 GND.n5610 301.784
R2792 GND.n5612 GND.n5611 301.784
R2793 GND.n5612 GND.n411 301.784
R2794 GND.n5620 GND.n411 301.784
R2795 GND.n5621 GND.n5620 301.784
R2796 GND.n5622 GND.n5621 301.784
R2797 GND.n5622 GND.n405 301.784
R2798 GND.n5630 GND.n405 301.784
R2799 GND.n5631 GND.n5630 301.784
R2800 GND.n5632 GND.n5631 301.784
R2801 GND.n5632 GND.n399 301.784
R2802 GND.n5640 GND.n399 301.784
R2803 GND.n5641 GND.n5640 301.784
R2804 GND.n5642 GND.n5641 301.784
R2805 GND.n5642 GND.n393 301.784
R2806 GND.n5650 GND.n393 301.784
R2807 GND.n5651 GND.n5650 301.784
R2808 GND.n5652 GND.n5651 301.784
R2809 GND.n5652 GND.n387 301.784
R2810 GND.n5660 GND.n387 301.784
R2811 GND.n5661 GND.n5660 301.784
R2812 GND.n5662 GND.n5661 301.784
R2813 GND.n5662 GND.n381 301.784
R2814 GND.n5670 GND.n381 301.784
R2815 GND.n5671 GND.n5670 301.784
R2816 GND.n5672 GND.n5671 301.784
R2817 GND.n5672 GND.n375 301.784
R2818 GND.n5682 GND.n375 301.784
R2819 GND.n53 GND.n47 289.615
R2820 GND.n64 GND.n58 289.615
R2821 GND.n29 GND.n23 289.615
R2822 GND.n40 GND.n34 289.615
R2823 GND.n6 GND.n0 289.615
R2824 GND.n17 GND.n11 289.615
R2825 GND.n1464 GND.n1463 289.615
R2826 GND.n1242 GND.n1241 289.615
R2827 GND.n136 GND.n130 289.615
R2828 GND.n125 GND.n119 289.615
R2829 GND.n112 GND.n106 289.615
R2830 GND.n101 GND.n95 289.615
R2831 GND.n89 GND.n83 289.615
R2832 GND.n78 GND.n72 289.615
R2833 GND.n2500 GND.n2499 289.615
R2834 GND.n2465 GND.n2464 289.615
R2835 GND.n4972 GND.n795 280.613
R2836 GND.n4980 GND.n795 280.613
R2837 GND.n4981 GND.n4980 280.613
R2838 GND.n4982 GND.n4981 280.613
R2839 GND.n4982 GND.n789 280.613
R2840 GND.n4990 GND.n789 280.613
R2841 GND.n4991 GND.n4990 280.613
R2842 GND.n4992 GND.n4991 280.613
R2843 GND.n4992 GND.n783 280.613
R2844 GND.n5000 GND.n783 280.613
R2845 GND.n5001 GND.n5000 280.613
R2846 GND.n5002 GND.n5001 280.613
R2847 GND.n5002 GND.n777 280.613
R2848 GND.n5010 GND.n777 280.613
R2849 GND.n5011 GND.n5010 280.613
R2850 GND.n5012 GND.n5011 280.613
R2851 GND.n5012 GND.n771 280.613
R2852 GND.n5020 GND.n771 280.613
R2853 GND.n5021 GND.n5020 280.613
R2854 GND.n5022 GND.n5021 280.613
R2855 GND.n5022 GND.n765 280.613
R2856 GND.n5030 GND.n765 280.613
R2857 GND.n5031 GND.n5030 280.613
R2858 GND.n5032 GND.n5031 280.613
R2859 GND.n5032 GND.n759 280.613
R2860 GND.n5040 GND.n759 280.613
R2861 GND.n5041 GND.n5040 280.613
R2862 GND.n5042 GND.n5041 280.613
R2863 GND.n5042 GND.n753 280.613
R2864 GND.n5050 GND.n753 280.613
R2865 GND.n5051 GND.n5050 280.613
R2866 GND.n5052 GND.n5051 280.613
R2867 GND.n5052 GND.n747 280.613
R2868 GND.n5060 GND.n747 280.613
R2869 GND.n5061 GND.n5060 280.613
R2870 GND.n5062 GND.n5061 280.613
R2871 GND.n5062 GND.n741 280.613
R2872 GND.n5070 GND.n741 280.613
R2873 GND.n5071 GND.n5070 280.613
R2874 GND.n5072 GND.n5071 280.613
R2875 GND.n5072 GND.n735 280.613
R2876 GND.n5080 GND.n735 280.613
R2877 GND.n5081 GND.n5080 280.613
R2878 GND.n5082 GND.n5081 280.613
R2879 GND.n5082 GND.n729 280.613
R2880 GND.n5090 GND.n729 280.613
R2881 GND.n5091 GND.n5090 280.613
R2882 GND.n5092 GND.n5091 280.613
R2883 GND.n5092 GND.n723 280.613
R2884 GND.n5100 GND.n723 280.613
R2885 GND.n5101 GND.n5100 280.613
R2886 GND.n5102 GND.n5101 280.613
R2887 GND.n5102 GND.n717 280.613
R2888 GND.n5110 GND.n717 280.613
R2889 GND.n5111 GND.n5110 280.613
R2890 GND.n5112 GND.n5111 280.613
R2891 GND.n5112 GND.n711 280.613
R2892 GND.n5120 GND.n711 280.613
R2893 GND.n5121 GND.n5120 280.613
R2894 GND.n5122 GND.n5121 280.613
R2895 GND.n5122 GND.n705 280.613
R2896 GND.n5130 GND.n705 280.613
R2897 GND.n5131 GND.n5130 280.613
R2898 GND.n5132 GND.n5131 280.613
R2899 GND.n5132 GND.n699 280.613
R2900 GND.n5140 GND.n699 280.613
R2901 GND.n5141 GND.n5140 280.613
R2902 GND.n5142 GND.n5141 280.613
R2903 GND.n5142 GND.n693 280.613
R2904 GND.n5150 GND.n693 280.613
R2905 GND.n5151 GND.n5150 280.613
R2906 GND.n5152 GND.n5151 280.613
R2907 GND.n5152 GND.n687 280.613
R2908 GND.n5160 GND.n687 280.613
R2909 GND.n5161 GND.n5160 280.613
R2910 GND.n5162 GND.n5161 280.613
R2911 GND.n5162 GND.n681 280.613
R2912 GND.n5170 GND.n681 280.613
R2913 GND.n5171 GND.n5170 280.613
R2914 GND.n5172 GND.n5171 280.613
R2915 GND.n5172 GND.n675 280.613
R2916 GND.n5180 GND.n675 280.613
R2917 GND.n5181 GND.n5180 280.613
R2918 GND.n5182 GND.n5181 280.613
R2919 GND.n5182 GND.n669 280.613
R2920 GND.n5190 GND.n669 280.613
R2921 GND.n5191 GND.n5190 280.613
R2922 GND.n5192 GND.n5191 280.613
R2923 GND.n5192 GND.n663 280.613
R2924 GND.n5200 GND.n663 280.613
R2925 GND.n5201 GND.n5200 280.613
R2926 GND.n5202 GND.n5201 280.613
R2927 GND.n5202 GND.n657 280.613
R2928 GND.n5210 GND.n657 280.613
R2929 GND.n5211 GND.n5210 280.613
R2930 GND.n5212 GND.n5211 280.613
R2931 GND.n5212 GND.n651 280.613
R2932 GND.n5220 GND.n651 280.613
R2933 GND.n5221 GND.n5220 280.613
R2934 GND.n5222 GND.n5221 280.613
R2935 GND.n5222 GND.n645 280.613
R2936 GND.n5230 GND.n645 280.613
R2937 GND.n5231 GND.n5230 280.613
R2938 GND.n5232 GND.n5231 280.613
R2939 GND.n5232 GND.n639 280.613
R2940 GND.n5240 GND.n639 280.613
R2941 GND.n5241 GND.n5240 280.613
R2942 GND.n5242 GND.n5241 280.613
R2943 GND.n5242 GND.n633 280.613
R2944 GND.n5250 GND.n633 280.613
R2945 GND.n5251 GND.n5250 280.613
R2946 GND.n5252 GND.n5251 280.613
R2947 GND.n5252 GND.n627 280.613
R2948 GND.n5260 GND.n627 280.613
R2949 GND.n5261 GND.n5260 280.613
R2950 GND.n5262 GND.n5261 280.613
R2951 GND.n5262 GND.n621 280.613
R2952 GND.n5270 GND.n621 280.613
R2953 GND.n5271 GND.n5270 280.613
R2954 GND.n5272 GND.n5271 280.613
R2955 GND.n5272 GND.n615 280.613
R2956 GND.n5280 GND.n615 280.613
R2957 GND.n5281 GND.n5280 280.613
R2958 GND.n5282 GND.n5281 280.613
R2959 GND.n5282 GND.n609 280.613
R2960 GND.n5290 GND.n609 280.613
R2961 GND.n5291 GND.n5290 280.613
R2962 GND.n5292 GND.n5291 280.613
R2963 GND.n5292 GND.n603 280.613
R2964 GND.n5300 GND.n603 280.613
R2965 GND.n5301 GND.n5300 280.613
R2966 GND.n5302 GND.n5301 280.613
R2967 GND.n5302 GND.n597 280.613
R2968 GND.n5310 GND.n597 280.613
R2969 GND.n5311 GND.n5310 280.613
R2970 GND.n5312 GND.n5311 280.613
R2971 GND.n5312 GND.n591 280.613
R2972 GND.n5320 GND.n591 280.613
R2973 GND.n5321 GND.n5320 280.613
R2974 GND.n5322 GND.n5321 280.613
R2975 GND.n5322 GND.n585 280.613
R2976 GND.n5330 GND.n585 280.613
R2977 GND.n5331 GND.n5330 280.613
R2978 GND.n5332 GND.n5331 280.613
R2979 GND.n5332 GND.n579 280.613
R2980 GND.n5340 GND.n579 280.613
R2981 GND.n5341 GND.n5340 280.613
R2982 GND.n5342 GND.n5341 280.613
R2983 GND.n5342 GND.n573 280.613
R2984 GND.n5350 GND.n573 280.613
R2985 GND.n5351 GND.n5350 280.613
R2986 GND.n5352 GND.n5351 280.613
R2987 GND.n5352 GND.n567 280.613
R2988 GND.n5360 GND.n567 280.613
R2989 GND.n5361 GND.n5360 280.613
R2990 GND.n5362 GND.n5361 280.613
R2991 GND.n5362 GND.n561 280.613
R2992 GND.n5370 GND.n561 280.613
R2993 GND.n5371 GND.n5370 280.613
R2994 GND.n5372 GND.n5371 280.613
R2995 GND.n5372 GND.n555 280.613
R2996 GND.n5380 GND.n555 280.613
R2997 GND.n5381 GND.n5380 280.613
R2998 GND.n5382 GND.n5381 280.613
R2999 GND.n5382 GND.n549 280.613
R3000 GND.n5390 GND.n549 280.613
R3001 GND.n5391 GND.n5390 280.613
R3002 GND.n5392 GND.n5391 280.613
R3003 GND.n5392 GND.n543 280.613
R3004 GND.n5400 GND.n543 280.613
R3005 GND.n5401 GND.n5400 280.613
R3006 GND.n5402 GND.n5401 280.613
R3007 GND.n5402 GND.n537 280.613
R3008 GND.n5410 GND.n537 280.613
R3009 GND.n5411 GND.n5410 280.613
R3010 GND.n5412 GND.n5411 280.613
R3011 GND.n5412 GND.n531 280.613
R3012 GND.n5420 GND.n531 280.613
R3013 GND.n5421 GND.n5420 280.613
R3014 GND.n5422 GND.n5421 280.613
R3015 GND.n5422 GND.n525 280.613
R3016 GND.n5430 GND.n525 280.613
R3017 GND.n5431 GND.n5430 280.613
R3018 GND.n5432 GND.n5431 280.613
R3019 GND.n5432 GND.n519 280.613
R3020 GND.n5440 GND.n519 280.613
R3021 GND.n5441 GND.n5440 280.613
R3022 GND.n5442 GND.n5441 280.613
R3023 GND.n5442 GND.n513 280.613
R3024 GND.n5450 GND.n513 280.613
R3025 GND.n5451 GND.n5450 280.613
R3026 GND.n5452 GND.n5451 280.613
R3027 GND.n5452 GND.n507 280.613
R3028 GND.n5460 GND.n507 280.613
R3029 GND.n5461 GND.n5460 280.613
R3030 GND.n5462 GND.n5461 280.613
R3031 GND.n5462 GND.n501 280.613
R3032 GND.n5470 GND.n501 280.613
R3033 GND.n5471 GND.n5470 280.613
R3034 GND.n5472 GND.n5471 280.613
R3035 GND.n5472 GND.n495 280.613
R3036 GND.n5480 GND.n495 280.613
R3037 GND.n5481 GND.n5480 280.613
R3038 GND.n5482 GND.n5481 280.613
R3039 GND.n5482 GND.n489 280.613
R3040 GND.n5490 GND.n489 280.613
R3041 GND.n5491 GND.n5490 280.613
R3042 GND.n5492 GND.n5491 280.613
R3043 GND.n5492 GND.n483 280.613
R3044 GND.n5500 GND.n483 280.613
R3045 GND.n5501 GND.n5500 280.613
R3046 GND.n5502 GND.n5501 280.613
R3047 GND.n5502 GND.n477 280.613
R3048 GND.n5510 GND.n477 280.613
R3049 GND.n5511 GND.n5510 280.613
R3050 GND.n5512 GND.n5511 280.613
R3051 GND.n5512 GND.n471 280.613
R3052 GND.n5520 GND.n471 280.613
R3053 GND.n5521 GND.n5520 280.613
R3054 GND.n5522 GND.n5521 280.613
R3055 GND.n5522 GND.n465 280.613
R3056 GND.n5530 GND.n465 280.613
R3057 GND.n5531 GND.n5530 280.613
R3058 GND.n5532 GND.n5531 280.613
R3059 GND.n5532 GND.n459 280.613
R3060 GND.n5540 GND.n459 280.613
R3061 GND.n5541 GND.n5540 280.613
R3062 GND.n5542 GND.n5541 280.613
R3063 GND.n3835 GND.t50 277.594
R3064 GND.n3230 GND.t40 277.594
R3065 GND.n3301 GND.t60 271.697
R3066 GND.n3069 GND.t89 271.697
R3067 GND.n3308 GND.t115 271.697
R3068 GND.n3061 GND.t76 271.697
R3069 GND.n3336 GND.n2053 256.663
R3070 GND.n3342 GND.n2053 256.663
R3071 GND.n3344 GND.n2053 256.663
R3072 GND.n3350 GND.n2053 256.663
R3073 GND.n3352 GND.n2053 256.663
R3074 GND.n3358 GND.n2053 256.663
R3075 GND.n3360 GND.n2053 256.663
R3076 GND.n3366 GND.n2053 256.663
R3077 GND.n3368 GND.n2053 256.663
R3078 GND.n3374 GND.n2053 256.663
R3079 GND.n3376 GND.n2053 256.663
R3080 GND.n3382 GND.n2053 256.663
R3081 GND.n3384 GND.n2053 256.663
R3082 GND.n3390 GND.n2053 256.663
R3083 GND.n3393 GND.n2053 256.663
R3084 GND.n3395 GND.n2053 256.663
R3085 GND.n3401 GND.n2053 256.663
R3086 GND.n3403 GND.n2053 256.663
R3087 GND.n3409 GND.n2053 256.663
R3088 GND.n3411 GND.n2053 256.663
R3089 GND.n3417 GND.n2053 256.663
R3090 GND.n3419 GND.n2053 256.663
R3091 GND.n3425 GND.n2053 256.663
R3092 GND.n3427 GND.n2053 256.663
R3093 GND.n3433 GND.n2053 256.663
R3094 GND.n3435 GND.n2053 256.663
R3095 GND.n3441 GND.n2053 256.663
R3096 GND.n3443 GND.n2053 256.663
R3097 GND.n3449 GND.n2053 256.663
R3098 GND.n3898 GND.n3021 256.663
R3099 GND.n3088 GND.n3021 256.663
R3100 GND.n3905 GND.n3021 256.663
R3101 GND.n3085 GND.n3021 256.663
R3102 GND.n3912 GND.n3021 256.663
R3103 GND.n3082 GND.n3021 256.663
R3104 GND.n3919 GND.n3021 256.663
R3105 GND.n3079 GND.n3021 256.663
R3106 GND.n3926 GND.n3021 256.663
R3107 GND.n3076 GND.n3021 256.663
R3108 GND.n3933 GND.n3021 256.663
R3109 GND.n3073 GND.n3021 256.663
R3110 GND.n3940 GND.n3021 256.663
R3111 GND.n3067 GND.n3021 256.663
R3112 GND.n3947 GND.n3021 256.663
R3113 GND.n3948 GND.n2405 256.663
R3114 GND.n3949 GND.n3021 256.663
R3115 GND.n3954 GND.n3021 256.663
R3116 GND.n3064 GND.n3021 256.663
R3117 GND.n3962 GND.n3021 256.663
R3118 GND.n3059 GND.n3021 256.663
R3119 GND.n3969 GND.n3021 256.663
R3120 GND.n3056 GND.n3021 256.663
R3121 GND.n3976 GND.n3021 256.663
R3122 GND.n3053 GND.n3021 256.663
R3123 GND.n3983 GND.n3021 256.663
R3124 GND.n3050 GND.n3021 256.663
R3125 GND.n3990 GND.n3021 256.663
R3126 GND.n3047 GND.n3021 256.663
R3127 GND.n3997 GND.n3021 256.663
R3128 GND.n3044 GND.n3021 256.663
R3129 GND.n3278 GND.n3277 242.672
R3130 GND.n3278 GND.n3200 242.672
R3131 GND.n3278 GND.n3201 242.672
R3132 GND.n3278 GND.n3202 242.672
R3133 GND.n3278 GND.n3203 242.672
R3134 GND.n3278 GND.n3204 242.672
R3135 GND.n3278 GND.n3205 242.672
R3136 GND.n3278 GND.n3206 242.672
R3137 GND.n3278 GND.n3207 242.672
R3138 GND.n3278 GND.n3208 242.672
R3139 GND.n3279 GND.n3278 242.672
R3140 GND.n3882 GND.n3881 242.672
R3141 GND.n3881 GND.n3808 242.672
R3142 GND.n3881 GND.n3809 242.672
R3143 GND.n3881 GND.n3810 242.672
R3144 GND.n3881 GND.n3811 242.672
R3145 GND.n3881 GND.n3812 242.672
R3146 GND.n3881 GND.n3813 242.672
R3147 GND.n3881 GND.n3814 242.672
R3148 GND.n3881 GND.n3815 242.672
R3149 GND.n3881 GND.n3816 242.672
R3150 GND.n3881 GND.n3817 242.672
R3151 GND.n4800 GND.n966 242.672
R3152 GND.n4800 GND.n967 242.672
R3153 GND.n4800 GND.n968 242.672
R3154 GND.n4800 GND.n969 242.672
R3155 GND.n4800 GND.n970 242.672
R3156 GND.n4800 GND.n971 242.672
R3157 GND.n4800 GND.n972 242.672
R3158 GND.n4800 GND.n973 242.672
R3159 GND.n4800 GND.n974 242.672
R3160 GND.n4651 GND.n4639 242.672
R3161 GND.n4651 GND.n4640 242.672
R3162 GND.n4651 GND.n4642 242.672
R3163 GND.n4651 GND.n4643 242.672
R3164 GND.n4651 GND.n4645 242.672
R3165 GND.n4651 GND.n4646 242.672
R3166 GND.n4687 GND.n1189 242.672
R3167 GND.n4651 GND.n4647 242.672
R3168 GND.n4651 GND.n4649 242.672
R3169 GND.n4651 GND.n4650 242.672
R3170 GND.n4425 GND.n2391 242.672
R3171 GND.n4425 GND.n2392 242.672
R3172 GND.n4425 GND.n2393 242.672
R3173 GND.n4425 GND.n2394 242.672
R3174 GND.n5790 GND.n277 242.672
R3175 GND.n5790 GND.n276 242.672
R3176 GND.n5790 GND.n275 242.672
R3177 GND.n5790 GND.n274 242.672
R3178 GND.n4425 GND.n4424 242.672
R3179 GND.n4425 GND.n2383 242.672
R3180 GND.n4425 GND.n2384 242.672
R3181 GND.n4413 GND.n2406 242.672
R3182 GND.n4425 GND.n2385 242.672
R3183 GND.n4425 GND.n2386 242.672
R3184 GND.n4425 GND.n2387 242.672
R3185 GND.n4425 GND.n2388 242.672
R3186 GND.n4425 GND.n2389 242.672
R3187 GND.n4425 GND.n2390 242.672
R3188 GND.n5790 GND.n279 242.672
R3189 GND.n5790 GND.n280 242.672
R3190 GND.n5790 GND.n281 242.672
R3191 GND.n5790 GND.n282 242.672
R3192 GND.n5790 GND.n283 242.672
R3193 GND.n5790 GND.n284 242.672
R3194 GND.n5790 GND.n285 242.672
R3195 GND.n5790 GND.n286 242.672
R3196 GND.n5790 GND.n5789 242.672
R3197 GND.n4800 GND.n976 242.672
R3198 GND.n4800 GND.n977 242.672
R3199 GND.n4800 GND.n978 242.672
R3200 GND.n4800 GND.n979 242.672
R3201 GND.n4651 GND.n1483 242.672
R3202 GND.n4651 GND.n1482 242.672
R3203 GND.n4651 GND.n1481 242.672
R3204 GND.n4651 GND.n1479 242.672
R3205 GND.n3301 GND.t63 240.314
R3206 GND.n3069 GND.t90 240.314
R3207 GND.n3308 GND.t117 240.314
R3208 GND.n3061 GND.t78 240.314
R3209 GND.n5791 GND.n271 240.244
R3210 GND.n5788 GND.n287 240.244
R3211 GND.n5784 GND.n5783 240.244
R3212 GND.n5780 GND.n5779 240.244
R3213 GND.n5773 GND.n5772 240.244
R3214 GND.n5769 GND.n5768 240.244
R3215 GND.n5765 GND.n5764 240.244
R3216 GND.n5761 GND.n5760 240.244
R3217 GND.n5757 GND.n5756 240.244
R3218 GND.n4390 GND.n2424 240.244
R3219 GND.n4382 GND.n2424 240.244
R3220 GND.n4382 GND.n2808 240.244
R3221 GND.n2825 GND.n2808 240.244
R3222 GND.n4079 GND.n2825 240.244
R3223 GND.n4079 GND.n2837 240.244
R3224 GND.n4084 GND.n2837 240.244
R3225 GND.n4084 GND.n2848 240.244
R3226 GND.n4094 GND.n2848 240.244
R3227 GND.n4094 GND.n2858 240.244
R3228 GND.n4099 GND.n2858 240.244
R3229 GND.n4099 GND.n2869 240.244
R3230 GND.n4109 GND.n2869 240.244
R3231 GND.n4109 GND.n2879 240.244
R3232 GND.n4114 GND.n2879 240.244
R3233 GND.n4114 GND.n2891 240.244
R3234 GND.n4136 GND.n2891 240.244
R3235 GND.n4136 GND.n2901 240.244
R3236 GND.n2906 GND.n2901 240.244
R3237 GND.n4145 GND.n2906 240.244
R3238 GND.n4146 GND.n4145 240.244
R3239 GND.n4146 GND.n2916 240.244
R3240 GND.n4150 GND.n2916 240.244
R3241 GND.n4150 GND.n150 240.244
R3242 GND.n2928 GND.n150 240.244
R3243 GND.n4157 GND.n2928 240.244
R3244 GND.n4166 GND.n4157 240.244
R3245 GND.n4166 GND.n169 240.244
R3246 GND.n4170 GND.n169 240.244
R3247 GND.n4170 GND.n181 240.244
R3248 GND.n4180 GND.n181 240.244
R3249 GND.n4180 GND.n191 240.244
R3250 GND.n4184 GND.n191 240.244
R3251 GND.n4184 GND.n201 240.244
R3252 GND.n4194 GND.n201 240.244
R3253 GND.n4194 GND.n212 240.244
R3254 GND.n4198 GND.n212 240.244
R3255 GND.n4198 GND.n222 240.244
R3256 GND.n4209 GND.n222 240.244
R3257 GND.n4209 GND.n233 240.244
R3258 GND.n2956 GND.n233 240.244
R3259 GND.n2956 GND.n242 240.244
R3260 GND.n4255 GND.n242 240.244
R3261 GND.n4255 GND.n253 240.244
R3262 GND.n4251 GND.n253 240.244
R3263 GND.n4251 GND.n263 240.244
R3264 GND.n5749 GND.n263 240.244
R3265 GND.n2397 GND.n2396 240.244
R3266 GND.n4418 GND.n2396 240.244
R3267 GND.n4416 GND.n4415 240.244
R3268 GND.n4411 GND.n4410 240.244
R3269 GND.n4407 GND.n4406 240.244
R3270 GND.n4403 GND.n4402 240.244
R3271 GND.n4399 GND.n4398 240.244
R3272 GND.n2419 GND.n2418 240.244
R3273 GND.n2813 GND.n2398 240.244
R3274 GND.n4380 GND.n2813 240.244
R3275 GND.n4380 GND.n2814 240.244
R3276 GND.n4376 GND.n2814 240.244
R3277 GND.n4376 GND.n2823 240.244
R3278 GND.n4368 GND.n2823 240.244
R3279 GND.n4368 GND.n2840 240.244
R3280 GND.n4364 GND.n2840 240.244
R3281 GND.n4364 GND.n2846 240.244
R3282 GND.n4356 GND.n2846 240.244
R3283 GND.n4356 GND.n2861 240.244
R3284 GND.n4352 GND.n2861 240.244
R3285 GND.n4352 GND.n2867 240.244
R3286 GND.n4344 GND.n2867 240.244
R3287 GND.n4344 GND.n2882 240.244
R3288 GND.n4340 GND.n2882 240.244
R3289 GND.n4340 GND.n2889 240.244
R3290 GND.n4332 GND.n2889 240.244
R3291 GND.n4332 GND.n4329 240.244
R3292 GND.n4329 GND.n2904 240.244
R3293 GND.n4316 GND.n2904 240.244
R3294 GND.n4318 GND.n4316 240.244
R3295 GND.n4318 GND.n153 240.244
R3296 GND.n5858 GND.n153 240.244
R3297 GND.n5858 GND.n154 240.244
R3298 GND.n2930 GND.n154 240.244
R3299 GND.n2930 GND.n166 240.244
R3300 GND.n5853 GND.n166 240.244
R3301 GND.n5853 GND.n167 240.244
R3302 GND.n5845 GND.n167 240.244
R3303 GND.n5845 GND.n184 240.244
R3304 GND.n5841 GND.n184 240.244
R3305 GND.n5841 GND.n189 240.244
R3306 GND.n5833 GND.n189 240.244
R3307 GND.n5833 GND.n204 240.244
R3308 GND.n5829 GND.n204 240.244
R3309 GND.n5829 GND.n210 240.244
R3310 GND.n5821 GND.n210 240.244
R3311 GND.n5821 GND.n225 240.244
R3312 GND.n5817 GND.n225 240.244
R3313 GND.n5817 GND.n231 240.244
R3314 GND.n5809 GND.n231 240.244
R3315 GND.n5809 GND.n245 240.244
R3316 GND.n5805 GND.n245 240.244
R3317 GND.n5805 GND.n251 240.244
R3318 GND.n5797 GND.n251 240.244
R3319 GND.n5797 GND.n266 240.244
R3320 GND.n4225 GND.n273 240.244
R3321 GND.n4231 GND.n4230 240.244
R3322 GND.n4234 GND.n4233 240.244
R3323 GND.n4239 GND.n4221 240.244
R3324 GND.n2995 GND.n2381 240.244
R3325 GND.n2995 GND.n2810 240.244
R3326 GND.n3000 GND.n2810 240.244
R3327 GND.n3000 GND.n2826 240.244
R3328 GND.n3006 GND.n2826 240.244
R3329 GND.n3006 GND.n2838 240.244
R3330 GND.n4086 GND.n2838 240.244
R3331 GND.n4086 GND.n2849 240.244
R3332 GND.n4092 GND.n2849 240.244
R3333 GND.n4092 GND.n2859 240.244
R3334 GND.n4101 GND.n2859 240.244
R3335 GND.n4101 GND.n2870 240.244
R3336 GND.n4107 GND.n2870 240.244
R3337 GND.n4107 GND.n2880 240.244
R3338 GND.n4116 GND.n2880 240.244
R3339 GND.n4116 GND.n2892 240.244
R3340 GND.n4134 GND.n2892 240.244
R3341 GND.n4134 GND.n2902 240.244
R3342 GND.n2907 GND.n2902 240.244
R3343 GND.n4129 GND.n2907 240.244
R3344 GND.n4129 GND.n4128 240.244
R3345 GND.n4128 GND.n2917 240.244
R3346 GND.n2917 GND.n147 240.244
R3347 GND.n5860 GND.n147 240.244
R3348 GND.n5860 GND.n148 240.244
R3349 GND.n4159 GND.n148 240.244
R3350 GND.n4164 GND.n4159 240.244
R3351 GND.n4164 GND.n170 240.244
R3352 GND.n4172 GND.n170 240.244
R3353 GND.n4172 GND.n182 240.244
R3354 GND.n4178 GND.n182 240.244
R3355 GND.n4178 GND.n192 240.244
R3356 GND.n4186 GND.n192 240.244
R3357 GND.n4186 GND.n202 240.244
R3358 GND.n4192 GND.n202 240.244
R3359 GND.n4192 GND.n213 240.244
R3360 GND.n4200 GND.n213 240.244
R3361 GND.n4200 GND.n223 240.244
R3362 GND.n4207 GND.n223 240.244
R3363 GND.n4207 GND.n234 240.244
R3364 GND.n4261 GND.n234 240.244
R3365 GND.n4261 GND.n243 240.244
R3366 GND.n4257 GND.n243 240.244
R3367 GND.n4257 GND.n254 240.244
R3368 GND.n4249 GND.n254 240.244
R3369 GND.n4249 GND.n264 240.244
R3370 GND.n309 GND.n264 240.244
R3371 GND.n2799 GND.n2798 240.244
R3372 GND.n2795 GND.n2794 240.244
R3373 GND.n2791 GND.n2790 240.244
R3374 GND.n4426 GND.n2380 240.244
R3375 GND.n4388 GND.n2803 240.244
R3376 GND.n2812 GND.n2803 240.244
R3377 GND.n2828 GND.n2812 240.244
R3378 GND.n4374 GND.n2828 240.244
R3379 GND.n4374 GND.n2829 240.244
R3380 GND.n4370 GND.n2829 240.244
R3381 GND.n4370 GND.n2836 240.244
R3382 GND.n4362 GND.n2836 240.244
R3383 GND.n4362 GND.n2851 240.244
R3384 GND.n4358 GND.n2851 240.244
R3385 GND.n4358 GND.n2856 240.244
R3386 GND.n4350 GND.n2856 240.244
R3387 GND.n4350 GND.n2872 240.244
R3388 GND.n4346 GND.n2872 240.244
R3389 GND.n4346 GND.n2877 240.244
R3390 GND.n4338 GND.n2877 240.244
R3391 GND.n4338 GND.n2894 240.244
R3392 GND.n4334 GND.n2894 240.244
R3393 GND.n4334 GND.n2899 240.244
R3394 GND.n4141 GND.n2899 240.244
R3395 GND.n4141 GND.n2919 240.244
R3396 GND.n4315 GND.n2919 240.244
R3397 GND.n4315 GND.n2920 240.244
R3398 GND.n2920 GND.n152 240.244
R3399 GND.n4310 GND.n152 240.244
R3400 GND.n4310 GND.n2927 240.244
R3401 GND.n2927 GND.n172 240.244
R3402 GND.n5851 GND.n172 240.244
R3403 GND.n5851 GND.n173 240.244
R3404 GND.n5847 GND.n173 240.244
R3405 GND.n5847 GND.n179 240.244
R3406 GND.n5839 GND.n179 240.244
R3407 GND.n5839 GND.n194 240.244
R3408 GND.n5835 GND.n194 240.244
R3409 GND.n5835 GND.n199 240.244
R3410 GND.n5827 GND.n199 240.244
R3411 GND.n5827 GND.n215 240.244
R3412 GND.n5823 GND.n215 240.244
R3413 GND.n5823 GND.n220 240.244
R3414 GND.n5815 GND.n220 240.244
R3415 GND.n5815 GND.n236 240.244
R3416 GND.n5811 GND.n236 240.244
R3417 GND.n5811 GND.n241 240.244
R3418 GND.n5803 GND.n241 240.244
R3419 GND.n5803 GND.n256 240.244
R3420 GND.n5799 GND.n256 240.244
R3421 GND.n5799 GND.n261 240.244
R3422 GND.n1180 GND.n1176 240.244
R3423 GND.n4648 GND.n1181 240.244
R3424 GND.n1185 GND.n1184 240.244
R3425 GND.n4644 GND.n1191 240.244
R3426 GND.n1195 GND.n1194 240.244
R3427 GND.n4641 GND.n1196 240.244
R3428 GND.n1200 GND.n1199 240.244
R3429 GND.n4638 GND.n1201 240.244
R3430 GND.n1079 GND.n995 240.244
R3431 GND.n1079 GND.n1005 240.244
R3432 GND.n1081 GND.n1005 240.244
R3433 GND.n1082 GND.n1081 240.244
R3434 GND.n1735 GND.n1082 240.244
R3435 GND.n1735 GND.n1088 240.244
R3436 GND.n1089 GND.n1088 240.244
R3437 GND.n1090 GND.n1089 240.244
R3438 GND.n1715 GND.n1090 240.244
R3439 GND.n1715 GND.n1096 240.244
R3440 GND.n1097 GND.n1096 240.244
R3441 GND.n1098 GND.n1097 240.244
R3442 GND.n1703 GND.n1098 240.244
R3443 GND.n1703 GND.n1104 240.244
R3444 GND.n1105 GND.n1104 240.244
R3445 GND.n1106 GND.n1105 240.244
R3446 GND.n1679 GND.n1106 240.244
R3447 GND.n1679 GND.n1112 240.244
R3448 GND.n1113 GND.n1112 240.244
R3449 GND.n1114 GND.n1113 240.244
R3450 GND.n1587 GND.n1114 240.244
R3451 GND.n1587 GND.n1120 240.244
R3452 GND.n1121 GND.n1120 240.244
R3453 GND.n1122 GND.n1121 240.244
R3454 GND.n1608 GND.n1122 240.244
R3455 GND.n1608 GND.n1128 240.244
R3456 GND.n1129 GND.n1128 240.244
R3457 GND.n1130 GND.n1129 240.244
R3458 GND.n1564 GND.n1130 240.244
R3459 GND.n1564 GND.n1136 240.244
R3460 GND.n1137 GND.n1136 240.244
R3461 GND.n1138 GND.n1137 240.244
R3462 GND.n1964 GND.n1138 240.244
R3463 GND.n1964 GND.n1144 240.244
R3464 GND.n1145 GND.n1144 240.244
R3465 GND.n1146 GND.n1145 240.244
R3466 GND.n1530 GND.n1146 240.244
R3467 GND.n1530 GND.n1152 240.244
R3468 GND.n1153 GND.n1152 240.244
R3469 GND.n1154 GND.n1153 240.244
R3470 GND.n1511 GND.n1154 240.244
R3471 GND.n1511 GND.n1160 240.244
R3472 GND.n1161 GND.n1160 240.244
R3473 GND.n1162 GND.n1161 240.244
R3474 GND.n1492 GND.n1162 240.244
R3475 GND.n1492 GND.n1168 240.244
R3476 GND.n4701 GND.n1168 240.244
R3477 GND.n1034 GND.n1033 240.244
R3478 GND.n1041 GND.n1040 240.244
R3479 GND.n1044 GND.n1043 240.244
R3480 GND.n1051 GND.n1050 240.244
R3481 GND.n1055 GND.n1054 240.244
R3482 GND.n1061 GND.n1060 240.244
R3483 GND.n1065 GND.n1064 240.244
R3484 GND.n1020 GND.n1019 240.244
R3485 GND.n1015 GND.n975 240.244
R3486 GND.n4778 GND.n998 240.244
R3487 GND.n4774 GND.n998 240.244
R3488 GND.n4774 GND.n1003 240.244
R3489 GND.n1733 GND.n1003 240.244
R3490 GND.n1823 GND.n1733 240.244
R3491 GND.n1823 GND.n1726 240.244
R3492 GND.n1831 GND.n1726 240.244
R3493 GND.n1831 GND.n1728 240.244
R3494 GND.n1728 GND.n1709 240.244
R3495 GND.n1848 GND.n1709 240.244
R3496 GND.n1848 GND.n1702 240.244
R3497 GND.n1856 GND.n1702 240.244
R3498 GND.n1856 GND.n1705 240.244
R3499 GND.n1705 GND.n1687 240.244
R3500 GND.n1873 GND.n1687 240.244
R3501 GND.n1873 GND.n1683 240.244
R3502 GND.n1879 GND.n1683 240.244
R3503 GND.n1879 GND.n1579 240.244
R3504 GND.n1944 GND.n1579 240.244
R3505 GND.n1944 GND.n1580 240.244
R3506 GND.n1601 GND.n1580 240.244
R3507 GND.n1603 GND.n1601 240.244
R3508 GND.n1929 GND.n1603 240.244
R3509 GND.n1929 GND.n1926 240.244
R3510 GND.n1926 GND.n1604 240.244
R3511 GND.n1905 GND.n1604 240.244
R3512 GND.n1907 GND.n1905 240.244
R3513 GND.n1907 GND.n1567 240.244
R3514 GND.n1952 GND.n1567 240.244
R3515 GND.n1952 GND.n1569 240.244
R3516 GND.n1569 GND.n1551 240.244
R3517 GND.n1969 GND.n1551 240.244
R3518 GND.n1969 GND.n1545 240.244
R3519 GND.n1977 GND.n1545 240.244
R3520 GND.n1977 GND.n1547 240.244
R3521 GND.n1547 GND.n1528 240.244
R3522 GND.n1993 GND.n1528 240.244
R3523 GND.n1993 GND.n1522 240.244
R3524 GND.n2001 GND.n1522 240.244
R3525 GND.n2001 GND.n1524 240.244
R3526 GND.n1524 GND.n1505 240.244
R3527 GND.n2027 GND.n1505 240.244
R3528 GND.n2027 GND.n1500 240.244
R3529 GND.n2035 GND.n1500 240.244
R3530 GND.n2035 GND.n1501 240.244
R3531 GND.n1501 GND.n1175 240.244
R3532 GND.n4699 GND.n1175 240.244
R3533 GND.n3880 GND.n3818 240.244
R3534 GND.n3873 GND.n3872 240.244
R3535 GND.n3870 GND.n3869 240.244
R3536 GND.n3866 GND.n3865 240.244
R3537 GND.n3862 GND.n3861 240.244
R3538 GND.n3858 GND.n3857 240.244
R3539 GND.n3854 GND.n3853 240.244
R3540 GND.n3850 GND.n3849 240.244
R3541 GND.n3846 GND.n3845 240.244
R3542 GND.n3842 GND.n3841 240.244
R3543 GND.n3883 GND.n3807 240.244
R3544 GND.n3281 GND.n2071 240.244
R3545 GND.n3479 GND.n2071 240.244
R3546 GND.n3479 GND.n2080 240.244
R3547 GND.n3482 GND.n2080 240.244
R3548 GND.n3482 GND.n3193 240.244
R3549 GND.n3488 GND.n3193 240.244
R3550 GND.n3488 GND.n2100 240.244
R3551 GND.n3508 GND.n2100 240.244
R3552 GND.n3508 GND.n2115 240.244
R3553 GND.n3514 GND.n2115 240.244
R3554 GND.n3514 GND.n2125 240.244
R3555 GND.n3555 GND.n2125 240.244
R3556 GND.n3555 GND.n2135 240.244
R3557 GND.n3562 GND.n2135 240.244
R3558 GND.n3562 GND.n2145 240.244
R3559 GND.n3583 GND.n2145 240.244
R3560 GND.n3583 GND.n2155 240.244
R3561 GND.n3579 GND.n2155 240.244
R3562 GND.n3579 GND.n2165 240.244
R3563 GND.n3171 GND.n2165 240.244
R3564 GND.n3171 GND.n2175 240.244
R3565 GND.n3168 GND.n2175 240.244
R3566 GND.n3168 GND.n2184 240.244
R3567 GND.n3635 GND.n2184 240.244
R3568 GND.n3635 GND.n2193 240.244
R3569 GND.n3658 GND.n2193 240.244
R3570 GND.n3658 GND.n2203 240.244
R3571 GND.n3654 GND.n2203 240.244
R3572 GND.n3654 GND.n2213 240.244
R3573 GND.n3651 GND.n2213 240.244
R3574 GND.n3651 GND.n3650 240.244
R3575 GND.n3650 GND.n3649 240.244
R3576 GND.n3649 GND.n2233 240.244
R3577 GND.n3699 GND.n2233 240.244
R3578 GND.n3699 GND.n2250 240.244
R3579 GND.n3702 GND.n2250 240.244
R3580 GND.n3702 GND.n3117 240.244
R3581 GND.n3709 GND.n3117 240.244
R3582 GND.n3709 GND.n2277 240.244
R3583 GND.n3748 GND.n2277 240.244
R3584 GND.n3748 GND.n2293 240.244
R3585 GND.n3105 GND.n2293 240.244
R3586 GND.n3755 GND.n3105 240.244
R3587 GND.n3756 GND.n3755 240.244
R3588 GND.n3757 GND.n3756 240.244
R3589 GND.n3757 GND.n2326 240.244
R3590 GND.n3767 GND.n2326 240.244
R3591 GND.n3767 GND.n2345 240.244
R3592 GND.n3095 GND.n2345 240.244
R3593 GND.n3800 GND.n3095 240.244
R3594 GND.n3801 GND.n3800 240.244
R3595 GND.n3801 GND.n2369 240.244
R3596 GND.n3889 GND.n2369 240.244
R3597 GND.n3211 GND.n3210 240.244
R3598 GND.n3271 GND.n3210 240.244
R3599 GND.n3269 GND.n3268 240.244
R3600 GND.n3265 GND.n3264 240.244
R3601 GND.n3261 GND.n3260 240.244
R3602 GND.n3257 GND.n3256 240.244
R3603 GND.n3253 GND.n3252 240.244
R3604 GND.n3249 GND.n3248 240.244
R3605 GND.n3245 GND.n3244 240.244
R3606 GND.n3241 GND.n3240 240.244
R3607 GND.n3237 GND.n3199 240.244
R3608 GND.n4615 GND.n2073 240.244
R3609 GND.n4615 GND.n2074 240.244
R3610 GND.n4609 GND.n2074 240.244
R3611 GND.n4609 GND.n2079 240.244
R3612 GND.n2105 GND.n2079 240.244
R3613 GND.n2105 GND.n2102 240.244
R3614 GND.n4592 GND.n2102 240.244
R3615 GND.n4592 GND.n2103 240.244
R3616 GND.n4588 GND.n2103 240.244
R3617 GND.n4588 GND.n2113 240.244
R3618 GND.n4578 GND.n2113 240.244
R3619 GND.n4578 GND.n2127 240.244
R3620 GND.n4574 GND.n2127 240.244
R3621 GND.n4574 GND.n2133 240.244
R3622 GND.n4564 GND.n2133 240.244
R3623 GND.n4564 GND.n2147 240.244
R3624 GND.n4560 GND.n2147 240.244
R3625 GND.n4560 GND.n2153 240.244
R3626 GND.n4550 GND.n2153 240.244
R3627 GND.n4550 GND.n2167 240.244
R3628 GND.n4546 GND.n2167 240.244
R3629 GND.n4546 GND.n2173 240.244
R3630 GND.n4536 GND.n2173 240.244
R3631 GND.n4536 GND.n2185 240.244
R3632 GND.n4532 GND.n2185 240.244
R3633 GND.n4532 GND.n2191 240.244
R3634 GND.n4522 GND.n2191 240.244
R3635 GND.n4522 GND.n2205 240.244
R3636 GND.n4518 GND.n2205 240.244
R3637 GND.n4518 GND.n2211 240.244
R3638 GND.n2239 GND.n2211 240.244
R3639 GND.n2239 GND.n2235 240.244
R3640 GND.n4501 GND.n2235 240.244
R3641 GND.n4501 GND.n2236 240.244
R3642 GND.n4497 GND.n2236 240.244
R3643 GND.n4497 GND.n2247 240.244
R3644 GND.n2283 GND.n2247 240.244
R3645 GND.n2283 GND.n2279 240.244
R3646 GND.n4481 GND.n2279 240.244
R3647 GND.n4481 GND.n2280 240.244
R3648 GND.n4477 GND.n2280 240.244
R3649 GND.n4477 GND.n2291 240.244
R3650 GND.n2334 GND.n2291 240.244
R3651 GND.n2335 GND.n2334 240.244
R3652 GND.n2335 GND.n2328 240.244
R3653 GND.n4453 GND.n2328 240.244
R3654 GND.n4453 GND.n2329 240.244
R3655 GND.n4449 GND.n2329 240.244
R3656 GND.n4449 GND.n2343 240.244
R3657 GND.n3798 GND.n2343 240.244
R3658 GND.n3798 GND.n2370 240.244
R3659 GND.n4433 GND.n2370 240.244
R3660 GND.n4433 GND.n2371 240.244
R3661 GND.n4973 GND.n796 240.244
R3662 GND.n4979 GND.n796 240.244
R3663 GND.n4979 GND.n794 240.244
R3664 GND.n4983 GND.n794 240.244
R3665 GND.n4983 GND.n790 240.244
R3666 GND.n4989 GND.n790 240.244
R3667 GND.n4989 GND.n788 240.244
R3668 GND.n4993 GND.n788 240.244
R3669 GND.n4993 GND.n784 240.244
R3670 GND.n4999 GND.n784 240.244
R3671 GND.n4999 GND.n782 240.244
R3672 GND.n5003 GND.n782 240.244
R3673 GND.n5003 GND.n778 240.244
R3674 GND.n5009 GND.n778 240.244
R3675 GND.n5009 GND.n776 240.244
R3676 GND.n5013 GND.n776 240.244
R3677 GND.n5013 GND.n772 240.244
R3678 GND.n5019 GND.n772 240.244
R3679 GND.n5019 GND.n770 240.244
R3680 GND.n5023 GND.n770 240.244
R3681 GND.n5023 GND.n766 240.244
R3682 GND.n5029 GND.n766 240.244
R3683 GND.n5029 GND.n764 240.244
R3684 GND.n5033 GND.n764 240.244
R3685 GND.n5033 GND.n760 240.244
R3686 GND.n5039 GND.n760 240.244
R3687 GND.n5039 GND.n758 240.244
R3688 GND.n5043 GND.n758 240.244
R3689 GND.n5043 GND.n754 240.244
R3690 GND.n5049 GND.n754 240.244
R3691 GND.n5049 GND.n752 240.244
R3692 GND.n5053 GND.n752 240.244
R3693 GND.n5053 GND.n748 240.244
R3694 GND.n5059 GND.n748 240.244
R3695 GND.n5059 GND.n746 240.244
R3696 GND.n5063 GND.n746 240.244
R3697 GND.n5063 GND.n742 240.244
R3698 GND.n5069 GND.n742 240.244
R3699 GND.n5069 GND.n740 240.244
R3700 GND.n5073 GND.n740 240.244
R3701 GND.n5073 GND.n736 240.244
R3702 GND.n5079 GND.n736 240.244
R3703 GND.n5079 GND.n734 240.244
R3704 GND.n5083 GND.n734 240.244
R3705 GND.n5083 GND.n730 240.244
R3706 GND.n5089 GND.n730 240.244
R3707 GND.n5089 GND.n728 240.244
R3708 GND.n5093 GND.n728 240.244
R3709 GND.n5093 GND.n724 240.244
R3710 GND.n5099 GND.n724 240.244
R3711 GND.n5099 GND.n722 240.244
R3712 GND.n5103 GND.n722 240.244
R3713 GND.n5103 GND.n718 240.244
R3714 GND.n5109 GND.n718 240.244
R3715 GND.n5109 GND.n716 240.244
R3716 GND.n5113 GND.n716 240.244
R3717 GND.n5113 GND.n712 240.244
R3718 GND.n5119 GND.n712 240.244
R3719 GND.n5119 GND.n710 240.244
R3720 GND.n5123 GND.n710 240.244
R3721 GND.n5123 GND.n706 240.244
R3722 GND.n5129 GND.n706 240.244
R3723 GND.n5129 GND.n704 240.244
R3724 GND.n5133 GND.n704 240.244
R3725 GND.n5133 GND.n700 240.244
R3726 GND.n5139 GND.n700 240.244
R3727 GND.n5139 GND.n698 240.244
R3728 GND.n5143 GND.n698 240.244
R3729 GND.n5143 GND.n694 240.244
R3730 GND.n5149 GND.n694 240.244
R3731 GND.n5149 GND.n692 240.244
R3732 GND.n5153 GND.n692 240.244
R3733 GND.n5153 GND.n688 240.244
R3734 GND.n5159 GND.n688 240.244
R3735 GND.n5159 GND.n686 240.244
R3736 GND.n5163 GND.n686 240.244
R3737 GND.n5163 GND.n682 240.244
R3738 GND.n5169 GND.n682 240.244
R3739 GND.n5169 GND.n680 240.244
R3740 GND.n5173 GND.n680 240.244
R3741 GND.n5173 GND.n676 240.244
R3742 GND.n5179 GND.n676 240.244
R3743 GND.n5179 GND.n674 240.244
R3744 GND.n5183 GND.n674 240.244
R3745 GND.n5183 GND.n670 240.244
R3746 GND.n5189 GND.n670 240.244
R3747 GND.n5189 GND.n668 240.244
R3748 GND.n5193 GND.n668 240.244
R3749 GND.n5193 GND.n664 240.244
R3750 GND.n5199 GND.n664 240.244
R3751 GND.n5199 GND.n662 240.244
R3752 GND.n5203 GND.n662 240.244
R3753 GND.n5203 GND.n658 240.244
R3754 GND.n5209 GND.n658 240.244
R3755 GND.n5209 GND.n656 240.244
R3756 GND.n5213 GND.n656 240.244
R3757 GND.n5213 GND.n652 240.244
R3758 GND.n5219 GND.n652 240.244
R3759 GND.n5219 GND.n650 240.244
R3760 GND.n5223 GND.n650 240.244
R3761 GND.n5223 GND.n646 240.244
R3762 GND.n5229 GND.n646 240.244
R3763 GND.n5229 GND.n644 240.244
R3764 GND.n5233 GND.n644 240.244
R3765 GND.n5233 GND.n640 240.244
R3766 GND.n5239 GND.n640 240.244
R3767 GND.n5239 GND.n638 240.244
R3768 GND.n5243 GND.n638 240.244
R3769 GND.n5243 GND.n634 240.244
R3770 GND.n5249 GND.n634 240.244
R3771 GND.n5249 GND.n632 240.244
R3772 GND.n5253 GND.n632 240.244
R3773 GND.n5253 GND.n628 240.244
R3774 GND.n5259 GND.n628 240.244
R3775 GND.n5259 GND.n626 240.244
R3776 GND.n5263 GND.n626 240.244
R3777 GND.n5263 GND.n622 240.244
R3778 GND.n5269 GND.n622 240.244
R3779 GND.n5269 GND.n620 240.244
R3780 GND.n5273 GND.n620 240.244
R3781 GND.n5273 GND.n616 240.244
R3782 GND.n5279 GND.n616 240.244
R3783 GND.n5279 GND.n614 240.244
R3784 GND.n5283 GND.n614 240.244
R3785 GND.n5283 GND.n610 240.244
R3786 GND.n5289 GND.n610 240.244
R3787 GND.n5289 GND.n608 240.244
R3788 GND.n5293 GND.n608 240.244
R3789 GND.n5293 GND.n604 240.244
R3790 GND.n5299 GND.n604 240.244
R3791 GND.n5299 GND.n602 240.244
R3792 GND.n5303 GND.n602 240.244
R3793 GND.n5303 GND.n598 240.244
R3794 GND.n5309 GND.n598 240.244
R3795 GND.n5309 GND.n596 240.244
R3796 GND.n5313 GND.n596 240.244
R3797 GND.n5313 GND.n592 240.244
R3798 GND.n5319 GND.n592 240.244
R3799 GND.n5319 GND.n590 240.244
R3800 GND.n5323 GND.n590 240.244
R3801 GND.n5323 GND.n586 240.244
R3802 GND.n5329 GND.n586 240.244
R3803 GND.n5329 GND.n584 240.244
R3804 GND.n5333 GND.n584 240.244
R3805 GND.n5333 GND.n580 240.244
R3806 GND.n5339 GND.n580 240.244
R3807 GND.n5339 GND.n578 240.244
R3808 GND.n5343 GND.n578 240.244
R3809 GND.n5343 GND.n574 240.244
R3810 GND.n5349 GND.n574 240.244
R3811 GND.n5349 GND.n572 240.244
R3812 GND.n5353 GND.n572 240.244
R3813 GND.n5353 GND.n568 240.244
R3814 GND.n5359 GND.n568 240.244
R3815 GND.n5359 GND.n566 240.244
R3816 GND.n5363 GND.n566 240.244
R3817 GND.n5363 GND.n562 240.244
R3818 GND.n5369 GND.n562 240.244
R3819 GND.n5369 GND.n560 240.244
R3820 GND.n5373 GND.n560 240.244
R3821 GND.n5373 GND.n556 240.244
R3822 GND.n5379 GND.n556 240.244
R3823 GND.n5379 GND.n554 240.244
R3824 GND.n5383 GND.n554 240.244
R3825 GND.n5383 GND.n550 240.244
R3826 GND.n5389 GND.n550 240.244
R3827 GND.n5389 GND.n548 240.244
R3828 GND.n5393 GND.n548 240.244
R3829 GND.n5393 GND.n544 240.244
R3830 GND.n5399 GND.n544 240.244
R3831 GND.n5399 GND.n542 240.244
R3832 GND.n5403 GND.n542 240.244
R3833 GND.n5403 GND.n538 240.244
R3834 GND.n5409 GND.n538 240.244
R3835 GND.n5409 GND.n536 240.244
R3836 GND.n5413 GND.n536 240.244
R3837 GND.n5413 GND.n532 240.244
R3838 GND.n5419 GND.n532 240.244
R3839 GND.n5419 GND.n530 240.244
R3840 GND.n5423 GND.n530 240.244
R3841 GND.n5423 GND.n526 240.244
R3842 GND.n5429 GND.n526 240.244
R3843 GND.n5429 GND.n524 240.244
R3844 GND.n5433 GND.n524 240.244
R3845 GND.n5433 GND.n520 240.244
R3846 GND.n5439 GND.n520 240.244
R3847 GND.n5439 GND.n518 240.244
R3848 GND.n5443 GND.n518 240.244
R3849 GND.n5443 GND.n514 240.244
R3850 GND.n5449 GND.n514 240.244
R3851 GND.n5449 GND.n512 240.244
R3852 GND.n5453 GND.n512 240.244
R3853 GND.n5453 GND.n508 240.244
R3854 GND.n5459 GND.n508 240.244
R3855 GND.n5459 GND.n506 240.244
R3856 GND.n5463 GND.n506 240.244
R3857 GND.n5463 GND.n502 240.244
R3858 GND.n5469 GND.n502 240.244
R3859 GND.n5469 GND.n500 240.244
R3860 GND.n5473 GND.n500 240.244
R3861 GND.n5473 GND.n496 240.244
R3862 GND.n5479 GND.n496 240.244
R3863 GND.n5479 GND.n494 240.244
R3864 GND.n5483 GND.n494 240.244
R3865 GND.n5483 GND.n490 240.244
R3866 GND.n5489 GND.n490 240.244
R3867 GND.n5489 GND.n488 240.244
R3868 GND.n5493 GND.n488 240.244
R3869 GND.n5493 GND.n484 240.244
R3870 GND.n5499 GND.n484 240.244
R3871 GND.n5499 GND.n482 240.244
R3872 GND.n5503 GND.n482 240.244
R3873 GND.n5503 GND.n478 240.244
R3874 GND.n5509 GND.n478 240.244
R3875 GND.n5509 GND.n476 240.244
R3876 GND.n5513 GND.n476 240.244
R3877 GND.n5513 GND.n472 240.244
R3878 GND.n5519 GND.n472 240.244
R3879 GND.n5519 GND.n470 240.244
R3880 GND.n5523 GND.n470 240.244
R3881 GND.n5523 GND.n466 240.244
R3882 GND.n5529 GND.n466 240.244
R3883 GND.n5529 GND.n464 240.244
R3884 GND.n5533 GND.n464 240.244
R3885 GND.n5533 GND.n460 240.244
R3886 GND.n5539 GND.n460 240.244
R3887 GND.n5539 GND.n458 240.244
R3888 GND.n5543 GND.n458 240.244
R3889 GND.n5549 GND.n454 240.244
R3890 GND.n5549 GND.n452 240.244
R3891 GND.n5553 GND.n452 240.244
R3892 GND.n5553 GND.n448 240.244
R3893 GND.n5559 GND.n448 240.244
R3894 GND.n5559 GND.n446 240.244
R3895 GND.n5563 GND.n446 240.244
R3896 GND.n5563 GND.n442 240.244
R3897 GND.n5569 GND.n442 240.244
R3898 GND.n5569 GND.n440 240.244
R3899 GND.n5573 GND.n440 240.244
R3900 GND.n5573 GND.n436 240.244
R3901 GND.n5579 GND.n436 240.244
R3902 GND.n5579 GND.n434 240.244
R3903 GND.n5583 GND.n434 240.244
R3904 GND.n5583 GND.n430 240.244
R3905 GND.n5589 GND.n430 240.244
R3906 GND.n5589 GND.n428 240.244
R3907 GND.n5593 GND.n428 240.244
R3908 GND.n5593 GND.n424 240.244
R3909 GND.n5599 GND.n424 240.244
R3910 GND.n5599 GND.n422 240.244
R3911 GND.n5603 GND.n422 240.244
R3912 GND.n5603 GND.n418 240.244
R3913 GND.n5609 GND.n418 240.244
R3914 GND.n5609 GND.n416 240.244
R3915 GND.n5613 GND.n416 240.244
R3916 GND.n5613 GND.n412 240.244
R3917 GND.n5619 GND.n412 240.244
R3918 GND.n5619 GND.n410 240.244
R3919 GND.n5623 GND.n410 240.244
R3920 GND.n5623 GND.n406 240.244
R3921 GND.n5629 GND.n406 240.244
R3922 GND.n5629 GND.n404 240.244
R3923 GND.n5633 GND.n404 240.244
R3924 GND.n5633 GND.n400 240.244
R3925 GND.n5639 GND.n400 240.244
R3926 GND.n5639 GND.n398 240.244
R3927 GND.n5643 GND.n398 240.244
R3928 GND.n5643 GND.n394 240.244
R3929 GND.n5649 GND.n394 240.244
R3930 GND.n5649 GND.n392 240.244
R3931 GND.n5653 GND.n392 240.244
R3932 GND.n5653 GND.n388 240.244
R3933 GND.n5659 GND.n388 240.244
R3934 GND.n5659 GND.n386 240.244
R3935 GND.n5663 GND.n386 240.244
R3936 GND.n5663 GND.n382 240.244
R3937 GND.n5669 GND.n382 240.244
R3938 GND.n5669 GND.n380 240.244
R3939 GND.n5673 GND.n380 240.244
R3940 GND.n5673 GND.n376 240.244
R3941 GND.n5681 GND.n376 240.244
R3942 GND.n5681 GND.n374 240.244
R3943 GND.n4859 GND.n910 240.244
R3944 GND.n4855 GND.n910 240.244
R3945 GND.n4855 GND.n912 240.244
R3946 GND.n4851 GND.n912 240.244
R3947 GND.n4851 GND.n917 240.244
R3948 GND.n4847 GND.n917 240.244
R3949 GND.n4847 GND.n919 240.244
R3950 GND.n4843 GND.n919 240.244
R3951 GND.n4843 GND.n925 240.244
R3952 GND.n4839 GND.n925 240.244
R3953 GND.n4839 GND.n927 240.244
R3954 GND.n4835 GND.n927 240.244
R3955 GND.n4835 GND.n933 240.244
R3956 GND.n4831 GND.n933 240.244
R3957 GND.n4831 GND.n935 240.244
R3958 GND.n4827 GND.n935 240.244
R3959 GND.n4827 GND.n941 240.244
R3960 GND.n4823 GND.n941 240.244
R3961 GND.n4823 GND.n943 240.244
R3962 GND.n4819 GND.n943 240.244
R3963 GND.n4819 GND.n949 240.244
R3964 GND.n4815 GND.n949 240.244
R3965 GND.n4815 GND.n951 240.244
R3966 GND.n4811 GND.n951 240.244
R3967 GND.n4811 GND.n957 240.244
R3968 GND.n4807 GND.n957 240.244
R3969 GND.n4807 GND.n959 240.244
R3970 GND.n4803 GND.n959 240.244
R3971 GND.n4803 GND.n965 240.244
R3972 GND.n1748 GND.n965 240.244
R3973 GND.n1749 GND.n1748 240.244
R3974 GND.n1749 GND.n1743 240.244
R3975 GND.n1755 GND.n1743 240.244
R3976 GND.n1756 GND.n1755 240.244
R3977 GND.n1773 GND.n1756 240.244
R3978 GND.n1773 GND.n1738 240.244
R3979 GND.n1817 GND.n1738 240.244
R3980 GND.n1817 GND.n1739 240.244
R3981 GND.n1813 GND.n1739 240.244
R3982 GND.n1813 GND.n1812 240.244
R3983 GND.n1812 GND.n1811 240.244
R3984 GND.n1811 GND.n1781 240.244
R3985 GND.n1807 GND.n1781 240.244
R3986 GND.n1807 GND.n1806 240.244
R3987 GND.n1806 GND.n1805 240.244
R3988 GND.n1805 GND.n1787 240.244
R3989 GND.n1801 GND.n1787 240.244
R3990 GND.n1801 GND.n1800 240.244
R3991 GND.n1800 GND.n1799 240.244
R3992 GND.n1799 GND.n1793 240.244
R3993 GND.n1793 GND.n1589 240.244
R3994 GND.n1937 GND.n1589 240.244
R3995 GND.n1937 GND.n1590 240.244
R3996 GND.n1932 GND.n1590 240.244
R3997 GND.n1932 GND.n1593 240.244
R3998 GND.n1611 GND.n1593 240.244
R3999 GND.n1920 GND.n1611 240.244
R4000 GND.n1920 GND.n1612 240.244
R4001 GND.n1915 GND.n1612 240.244
R4002 GND.n1915 GND.n1666 240.244
R4003 GND.n1666 GND.n1665 240.244
R4004 GND.n1665 GND.n1617 240.244
R4005 GND.n1661 GND.n1617 240.244
R4006 GND.n1661 GND.n1660 240.244
R4007 GND.n1660 GND.n1659 240.244
R4008 GND.n1659 GND.n1623 240.244
R4009 GND.n1655 GND.n1623 240.244
R4010 GND.n1655 GND.n1654 240.244
R4011 GND.n1654 GND.n1653 240.244
R4012 GND.n1653 GND.n1629 240.244
R4013 GND.n1649 GND.n1629 240.244
R4014 GND.n1649 GND.n1648 240.244
R4015 GND.n1648 GND.n1647 240.244
R4016 GND.n1647 GND.n1635 240.244
R4017 GND.n1643 GND.n1635 240.244
R4018 GND.n1643 GND.n1490 240.244
R4019 GND.n2042 GND.n1490 240.244
R4020 GND.n2043 GND.n2042 240.244
R4021 GND.n2044 GND.n2043 240.244
R4022 GND.n2044 GND.n1485 240.244
R4023 GND.n4636 GND.n1485 240.244
R4024 GND.n4636 GND.n1486 240.244
R4025 GND.n4632 GND.n1486 240.244
R4026 GND.n4632 GND.n2052 240.244
R4027 GND.n4628 GND.n2052 240.244
R4028 GND.n4628 GND.n2054 240.244
R4029 GND.n4624 GND.n2054 240.244
R4030 GND.n4624 GND.n2060 240.244
R4031 GND.n3468 GND.n2060 240.244
R4032 GND.n3475 GND.n3468 240.244
R4033 GND.n3475 GND.n2091 240.244
R4034 GND.n4599 GND.n2091 240.244
R4035 GND.n4599 GND.n2092 240.244
R4036 GND.n4595 GND.n2092 240.244
R4037 GND.n4595 GND.n2098 240.244
R4038 GND.n3536 GND.n2098 240.244
R4039 GND.n3537 GND.n3536 240.244
R4040 GND.n3538 GND.n3537 240.244
R4041 GND.n3538 GND.n3528 240.244
R4042 GND.n3552 GND.n3528 240.244
R4043 GND.n3552 GND.n3529 240.244
R4044 GND.n3548 GND.n3529 240.244
R4045 GND.n3548 GND.n3154 240.244
R4046 GND.n3586 GND.n3154 240.244
R4047 GND.n3587 GND.n3586 240.244
R4048 GND.n3588 GND.n3587 240.244
R4049 GND.n3588 GND.n3150 240.244
R4050 GND.n3594 GND.n3150 240.244
R4051 GND.n3594 GND.n3144 240.244
R4052 GND.n3614 GND.n3144 240.244
R4053 GND.n3614 GND.n3139 240.244
R4054 GND.n3629 GND.n3139 240.244
R4055 GND.n3629 GND.n3140 240.244
R4056 GND.n3625 GND.n3140 240.244
R4057 GND.n3625 GND.n3624 240.244
R4058 GND.n3624 GND.n2215 240.244
R4059 GND.n4515 GND.n2215 240.244
R4060 GND.n4515 GND.n2216 240.244
R4061 GND.n4511 GND.n2216 240.244
R4062 GND.n4511 GND.n2222 240.244
R4063 GND.n2266 GND.n2222 240.244
R4064 GND.n2267 GND.n2266 240.244
R4065 GND.n2267 GND.n2260 240.244
R4066 GND.n4488 GND.n2260 240.244
R4067 GND.n4488 GND.n2261 240.244
R4068 GND.n4484 GND.n2261 240.244
R4069 GND.n4484 GND.n2275 240.244
R4070 GND.n2307 GND.n2275 240.244
R4071 GND.n2307 GND.n2303 240.244
R4072 GND.n4467 GND.n2303 240.244
R4073 GND.n4467 GND.n2304 240.244
R4074 GND.n4463 GND.n2304 240.244
R4075 GND.n4463 GND.n2315 240.244
R4076 GND.n2351 GND.n2315 240.244
R4077 GND.n2351 GND.n2347 240.244
R4078 GND.n4446 GND.n2347 240.244
R4079 GND.n4446 GND.n2348 240.244
R4080 GND.n4442 GND.n2348 240.244
R4081 GND.n4442 GND.n2359 240.244
R4082 GND.n3027 GND.n2359 240.244
R4083 GND.n4007 GND.n3027 240.244
R4084 GND.n4007 GND.n3022 240.244
R4085 GND.n4013 GND.n3022 240.244
R4086 GND.n4013 GND.n3020 240.244
R4087 GND.n4018 GND.n3020 240.244
R4088 GND.n4018 GND.n3016 240.244
R4089 GND.n4024 GND.n3016 240.244
R4090 GND.n4025 GND.n4024 240.244
R4091 GND.n4026 GND.n4025 240.244
R4092 GND.n4026 GND.n3012 240.244
R4093 GND.n4032 GND.n3012 240.244
R4094 GND.n4033 GND.n4032 240.244
R4095 GND.n4034 GND.n4033 240.244
R4096 GND.n4034 GND.n3007 240.244
R4097 GND.n4076 GND.n3007 240.244
R4098 GND.n4076 GND.n3008 240.244
R4099 GND.n4072 GND.n3008 240.244
R4100 GND.n4072 GND.n4071 240.244
R4101 GND.n4071 GND.n4070 240.244
R4102 GND.n4070 GND.n4042 240.244
R4103 GND.n4066 GND.n4042 240.244
R4104 GND.n4066 GND.n4065 240.244
R4105 GND.n4065 GND.n4064 240.244
R4106 GND.n4064 GND.n4048 240.244
R4107 GND.n4060 GND.n4048 240.244
R4108 GND.n4060 GND.n4059 240.244
R4109 GND.n4059 GND.n4058 240.244
R4110 GND.n4058 GND.n2909 240.244
R4111 GND.n4326 GND.n2909 240.244
R4112 GND.n4326 GND.n2910 240.244
R4113 GND.n4321 GND.n2910 240.244
R4114 GND.n4321 GND.n2913 240.244
R4115 GND.n2935 GND.n2913 240.244
R4116 GND.n2935 GND.n2932 240.244
R4117 GND.n4307 GND.n2932 240.244
R4118 GND.n4307 GND.n2933 240.244
R4119 GND.n4302 GND.n2933 240.244
R4120 GND.n4302 GND.n4301 240.244
R4121 GND.n4301 GND.n2940 240.244
R4122 GND.n4297 GND.n2940 240.244
R4123 GND.n4297 GND.n4296 240.244
R4124 GND.n4296 GND.n4295 240.244
R4125 GND.n4295 GND.n2944 240.244
R4126 GND.n4291 GND.n2944 240.244
R4127 GND.n4291 GND.n4290 240.244
R4128 GND.n4290 GND.n4289 240.244
R4129 GND.n4289 GND.n2950 240.244
R4130 GND.n4285 GND.n2950 240.244
R4131 GND.n4285 GND.n4284 240.244
R4132 GND.n4284 GND.n4283 240.244
R4133 GND.n4283 GND.n4264 240.244
R4134 GND.n4279 GND.n4264 240.244
R4135 GND.n4279 GND.n4278 240.244
R4136 GND.n4278 GND.n4277 240.244
R4137 GND.n4277 GND.n4270 240.244
R4138 GND.n4270 GND.n310 240.244
R4139 GND.n5746 GND.n310 240.244
R4140 GND.n5746 GND.n311 240.244
R4141 GND.n5742 GND.n311 240.244
R4142 GND.n5742 GND.n5741 240.244
R4143 GND.n5741 GND.n317 240.244
R4144 GND.n5737 GND.n317 240.244
R4145 GND.n5737 GND.n319 240.244
R4146 GND.n5733 GND.n319 240.244
R4147 GND.n5733 GND.n327 240.244
R4148 GND.n5729 GND.n327 240.244
R4149 GND.n5729 GND.n329 240.244
R4150 GND.n5725 GND.n329 240.244
R4151 GND.n5725 GND.n335 240.244
R4152 GND.n5721 GND.n335 240.244
R4153 GND.n5721 GND.n337 240.244
R4154 GND.n5717 GND.n337 240.244
R4155 GND.n5717 GND.n343 240.244
R4156 GND.n5713 GND.n343 240.244
R4157 GND.n5713 GND.n345 240.244
R4158 GND.n5709 GND.n345 240.244
R4159 GND.n5709 GND.n351 240.244
R4160 GND.n5705 GND.n351 240.244
R4161 GND.n5705 GND.n353 240.244
R4162 GND.n5701 GND.n353 240.244
R4163 GND.n5701 GND.n359 240.244
R4164 GND.n5697 GND.n359 240.244
R4165 GND.n5697 GND.n361 240.244
R4166 GND.n5693 GND.n361 240.244
R4167 GND.n5693 GND.n367 240.244
R4168 GND.n5689 GND.n367 240.244
R4169 GND.n5689 GND.n369 240.244
R4170 GND.n5685 GND.n369 240.244
R4171 GND.n4969 GND.n799 240.244
R4172 GND.n4969 GND.n801 240.244
R4173 GND.n4965 GND.n801 240.244
R4174 GND.n4965 GND.n807 240.244
R4175 GND.n4961 GND.n807 240.244
R4176 GND.n4961 GND.n809 240.244
R4177 GND.n4957 GND.n809 240.244
R4178 GND.n4957 GND.n815 240.244
R4179 GND.n4953 GND.n815 240.244
R4180 GND.n4953 GND.n817 240.244
R4181 GND.n4949 GND.n817 240.244
R4182 GND.n4949 GND.n823 240.244
R4183 GND.n4945 GND.n823 240.244
R4184 GND.n4945 GND.n825 240.244
R4185 GND.n4941 GND.n825 240.244
R4186 GND.n4941 GND.n831 240.244
R4187 GND.n4937 GND.n831 240.244
R4188 GND.n4937 GND.n833 240.244
R4189 GND.n4933 GND.n833 240.244
R4190 GND.n4933 GND.n839 240.244
R4191 GND.n4929 GND.n839 240.244
R4192 GND.n4929 GND.n841 240.244
R4193 GND.n4925 GND.n841 240.244
R4194 GND.n4925 GND.n847 240.244
R4195 GND.n4921 GND.n847 240.244
R4196 GND.n4921 GND.n849 240.244
R4197 GND.n4917 GND.n849 240.244
R4198 GND.n4917 GND.n855 240.244
R4199 GND.n4913 GND.n855 240.244
R4200 GND.n4913 GND.n857 240.244
R4201 GND.n4909 GND.n857 240.244
R4202 GND.n4909 GND.n863 240.244
R4203 GND.n4905 GND.n863 240.244
R4204 GND.n4905 GND.n865 240.244
R4205 GND.n4901 GND.n865 240.244
R4206 GND.n4901 GND.n871 240.244
R4207 GND.n4897 GND.n871 240.244
R4208 GND.n4897 GND.n873 240.244
R4209 GND.n4893 GND.n873 240.244
R4210 GND.n4893 GND.n879 240.244
R4211 GND.n4889 GND.n879 240.244
R4212 GND.n4889 GND.n881 240.244
R4213 GND.n4885 GND.n881 240.244
R4214 GND.n4885 GND.n887 240.244
R4215 GND.n4881 GND.n887 240.244
R4216 GND.n4881 GND.n889 240.244
R4217 GND.n4877 GND.n889 240.244
R4218 GND.n4877 GND.n895 240.244
R4219 GND.n4873 GND.n895 240.244
R4220 GND.n4873 GND.n897 240.244
R4221 GND.n4869 GND.n897 240.244
R4222 GND.n4869 GND.n903 240.244
R4223 GND.n4865 GND.n903 240.244
R4224 GND.n4865 GND.n905 240.244
R4225 GND.n4799 GND.n982 240.244
R4226 GND.n987 GND.n986 240.244
R4227 GND.n989 GND.n988 240.244
R4228 GND.n4784 GND.n4783 240.244
R4229 GND.n1008 GND.n981 240.244
R4230 GND.n4772 GND.n1008 240.244
R4231 GND.n4772 GND.n1009 240.244
R4232 GND.n1737 GND.n1009 240.244
R4233 GND.n1821 GND.n1737 240.244
R4234 GND.n1821 GND.n1820 240.244
R4235 GND.n1820 GND.n1725 240.244
R4236 GND.n1725 GND.n1713 240.244
R4237 GND.n1842 GND.n1713 240.244
R4238 GND.n1846 GND.n1842 240.244
R4239 GND.n1846 GND.n1845 240.244
R4240 GND.n1845 GND.n1701 240.244
R4241 GND.n1701 GND.n1691 240.244
R4242 GND.n1867 GND.n1691 240.244
R4243 GND.n1871 GND.n1867 240.244
R4244 GND.n1871 GND.n1869 240.244
R4245 GND.n1869 GND.n1682 240.244
R4246 GND.n1682 GND.n1584 240.244
R4247 GND.n1942 GND.n1584 240.244
R4248 GND.n1942 GND.n1940 240.244
R4249 GND.n1940 GND.n1585 240.244
R4250 GND.n1598 GND.n1585 240.244
R4251 GND.n1600 GND.n1598 240.244
R4252 GND.n1924 GND.n1600 240.244
R4253 GND.n1924 GND.n1923 240.244
R4254 GND.n1923 GND.n1607 240.244
R4255 GND.n1911 GND.n1607 240.244
R4256 GND.n1912 GND.n1911 240.244
R4257 GND.n1912 GND.n1566 240.244
R4258 GND.n1566 GND.n1555 240.244
R4259 GND.n1963 GND.n1555 240.244
R4260 GND.n1967 GND.n1963 240.244
R4261 GND.n1967 GND.n1966 240.244
R4262 GND.n1966 GND.n1544 240.244
R4263 GND.n1544 GND.n1534 240.244
R4264 GND.n1988 GND.n1534 240.244
R4265 GND.n1991 GND.n1988 240.244
R4266 GND.n1991 GND.n1990 240.244
R4267 GND.n1990 GND.n1521 240.244
R4268 GND.n1521 GND.n1509 240.244
R4269 GND.n2024 GND.n1509 240.244
R4270 GND.n2025 GND.n2024 240.244
R4271 GND.n2025 GND.n1496 240.244
R4272 GND.n2037 GND.n1496 240.244
R4273 GND.n2038 GND.n2037 240.244
R4274 GND.n2039 GND.n2038 240.244
R4275 GND.n2039 GND.n1174 240.244
R4276 GND.n1208 GND.n1207 240.244
R4277 GND.n1480 GND.n1468 240.244
R4278 GND.n1470 GND.n1469 240.244
R4279 GND.n4652 GND.n1477 240.244
R4280 GND.n4780 GND.n992 240.244
R4281 GND.n1006 GND.n992 240.244
R4282 GND.n1758 GND.n1006 240.244
R4283 GND.n1770 GND.n1758 240.244
R4284 GND.n1770 GND.n1736 240.244
R4285 GND.n1736 GND.n1721 240.244
R4286 GND.n1833 GND.n1721 240.244
R4287 GND.n1833 GND.n1716 240.244
R4288 GND.n1840 GND.n1716 240.244
R4289 GND.n1840 GND.n1711 240.244
R4290 GND.n1711 GND.n1698 240.244
R4291 GND.n1858 GND.n1698 240.244
R4292 GND.n1858 GND.n1693 240.244
R4293 GND.n1865 GND.n1693 240.244
R4294 GND.n1865 GND.n1689 240.244
R4295 GND.n1689 GND.n1676 240.244
R4296 GND.n1881 GND.n1676 240.244
R4297 GND.n1881 GND.n1677 240.244
R4298 GND.n1677 GND.n1582 240.244
R4299 GND.n1586 GND.n1582 240.244
R4300 GND.n1889 GND.n1586 240.244
R4301 GND.n1889 GND.n1888 240.244
R4302 GND.n1888 GND.n1596 240.244
R4303 GND.n1605 GND.n1596 240.244
R4304 GND.n1609 GND.n1605 240.244
R4305 GND.n1668 GND.n1609 240.244
R4306 GND.n1902 GND.n1668 240.244
R4307 GND.n1902 GND.n1563 240.244
R4308 GND.n1954 GND.n1563 240.244
R4309 GND.n1954 GND.n1558 240.244
R4310 GND.n1961 GND.n1558 240.244
R4311 GND.n1961 GND.n1553 240.244
R4312 GND.n1553 GND.n1541 240.244
R4313 GND.n1979 GND.n1541 240.244
R4314 GND.n1979 GND.n1536 240.244
R4315 GND.n1986 GND.n1536 240.244
R4316 GND.n1986 GND.n1531 240.244
R4317 GND.n1531 GND.n1517 240.244
R4318 GND.n2003 GND.n1517 240.244
R4319 GND.n2003 GND.n1512 240.244
R4320 GND.n2022 GND.n1512 240.244
R4321 GND.n2022 GND.n1507 240.244
R4322 GND.n2009 GND.n1507 240.244
R4323 GND.n2009 GND.n1498 240.244
R4324 GND.n2010 GND.n1498 240.244
R4325 GND.n2010 GND.n1494 240.244
R4326 GND.n1494 GND.n1171 240.244
R4327 GND.n1471 GND.t93 226.457
R4328 GND.n1186 GND.t56 226.457
R4329 GND.n1202 GND.t67 226.457
R4330 GND.n2408 GND.t120 226.457
R4331 GND.n2420 GND.t39 226.457
R4332 GND.n304 GND.t81 226.457
R4333 GND.n5775 GND.t74 226.457
R4334 GND.n4219 GND.t122 226.457
R4335 GND.n2377 GND.t85 226.457
R4336 GND.n1024 GND.t107 226.457
R4337 GND.n1016 GND.t98 226.457
R4338 GND.n4785 GND.t112 226.457
R4339 GND.n3835 GND.t52 223.011
R4340 GND.n3230 GND.t43 223.011
R4341 GND.n1471 GND.t92 210.257
R4342 GND.n1186 GND.t54 210.257
R4343 GND.n1202 GND.t66 210.257
R4344 GND.n2408 GND.t118 210.257
R4345 GND.n2420 GND.t36 210.257
R4346 GND.n304 GND.t80 210.257
R4347 GND.n5775 GND.t72 210.257
R4348 GND.n4219 GND.t121 210.257
R4349 GND.n2377 GND.t83 210.257
R4350 GND.n1024 GND.t105 210.257
R4351 GND.n1016 GND.t95 210.257
R4352 GND.n4785 GND.t110 210.257
R4353 GND.n2406 GND.n2384 199.319
R4354 GND.n2406 GND.n2385 199.319
R4355 GND.n4647 GND.n1189 199.319
R4356 GND.n4646 GND.n1189 199.319
R4357 GND.n3302 GND.t62 186.593
R4358 GND.n3070 GND.t91 186.593
R4359 GND.n3309 GND.t116 186.593
R4360 GND.n3062 GND.t79 186.593
R4361 GND.n3326 GND.n3325 186.49
R4362 GND.n3036 GND.n3035 186.49
R4363 GND.n54 GND.n53 185
R4364 GND.n52 GND.n51 185
R4365 GND.n65 GND.n64 185
R4366 GND.n63 GND.n62 185
R4367 GND.n30 GND.n29 185
R4368 GND.n28 GND.n27 185
R4369 GND.n41 GND.n40 185
R4370 GND.n39 GND.n38 185
R4371 GND.n7 GND.n6 185
R4372 GND.n5 GND.n4 185
R4373 GND.n18 GND.n17 185
R4374 GND.n16 GND.n15 185
R4375 GND.n1463 GND.n1462 185
R4376 GND.n1434 GND.n1433 185
R4377 GND.n1457 GND.n1456 185
R4378 GND.n1455 GND.n1454 185
R4379 GND.n1438 GND.n1437 185
R4380 GND.n1449 GND.n1448 185
R4381 GND.n1447 GND.n1446 185
R4382 GND.n1442 GND.n1441 185
R4383 GND.n1220 GND.n1219 185
R4384 GND.n1225 GND.n1224 185
R4385 GND.n1227 GND.n1226 185
R4386 GND.n1216 GND.n1215 185
R4387 GND.n1233 GND.n1232 185
R4388 GND.n1235 GND.n1234 185
R4389 GND.n1212 GND.n1211 185
R4390 GND.n1241 GND.n1240 185
R4391 GND.n137 GND.n136 185
R4392 GND.n135 GND.n134 185
R4393 GND.n126 GND.n125 185
R4394 GND.n124 GND.n123 185
R4395 GND.n113 GND.n112 185
R4396 GND.n111 GND.n110 185
R4397 GND.n102 GND.n101 185
R4398 GND.n100 GND.n99 185
R4399 GND.n90 GND.n89 185
R4400 GND.n88 GND.n87 185
R4401 GND.n79 GND.n78 185
R4402 GND.n77 GND.n76 185
R4403 GND.n2499 GND.n2498 185
R4404 GND.n2470 GND.n2469 185
R4405 GND.n2493 GND.n2492 185
R4406 GND.n2491 GND.n2490 185
R4407 GND.n2474 GND.n2473 185
R4408 GND.n2485 GND.n2484 185
R4409 GND.n2483 GND.n2482 185
R4410 GND.n2478 GND.n2477 185
R4411 GND.n2443 GND.n2442 185
R4412 GND.n2448 GND.n2447 185
R4413 GND.n2450 GND.n2449 185
R4414 GND.n2439 GND.n2438 185
R4415 GND.n2456 GND.n2455 185
R4416 GND.n2458 GND.n2457 185
R4417 GND.n2435 GND.n2434 185
R4418 GND.n2464 GND.n2463 185
R4419 GND.n3836 GND.t53 177.435
R4420 GND.n3231 GND.t42 177.435
R4421 GND.n3999 GND.n3998 163.367
R4422 GND.n3996 GND.n3045 163.367
R4423 GND.n3992 GND.n3991 163.367
R4424 GND.n3989 GND.n3048 163.367
R4425 GND.n3985 GND.n3984 163.367
R4426 GND.n3982 GND.n3051 163.367
R4427 GND.n3978 GND.n3977 163.367
R4428 GND.n3975 GND.n3054 163.367
R4429 GND.n3971 GND.n3970 163.367
R4430 GND.n3968 GND.n3057 163.367
R4431 GND.n3964 GND.n3963 163.367
R4432 GND.n3961 GND.n3060 163.367
R4433 GND.n3956 GND.n3955 163.367
R4434 GND.n3953 GND.n3950 163.367
R4435 GND.n3946 GND.n3065 163.367
R4436 GND.n3942 GND.n3941 163.367
R4437 GND.n3939 GND.n3068 163.367
R4438 GND.n3935 GND.n3934 163.367
R4439 GND.n3932 GND.n3074 163.367
R4440 GND.n3928 GND.n3927 163.367
R4441 GND.n3925 GND.n3077 163.367
R4442 GND.n3921 GND.n3920 163.367
R4443 GND.n3918 GND.n3080 163.367
R4444 GND.n3914 GND.n3913 163.367
R4445 GND.n3911 GND.n3083 163.367
R4446 GND.n3907 GND.n3906 163.367
R4447 GND.n3904 GND.n3086 163.367
R4448 GND.n3900 GND.n3899 163.367
R4449 GND.n3452 GND.n2062 163.367
R4450 GND.n3456 GND.n2062 163.367
R4451 GND.n3456 GND.n2070 163.367
R4452 GND.n3287 GND.n2070 163.367
R4453 GND.n3467 GND.n3287 163.367
R4454 GND.n3467 GND.n2081 163.367
R4455 GND.n3463 GND.n2081 163.367
R4456 GND.n3463 GND.n2089 163.367
R4457 GND.n3189 GND.n2089 163.367
R4458 GND.n3499 GND.n3189 163.367
R4459 GND.n3500 GND.n3499 163.367
R4460 GND.n3501 GND.n3500 163.367
R4461 GND.n3501 GND.n3187 163.367
R4462 GND.n3505 GND.n3187 163.367
R4463 GND.n3505 GND.n2116 163.367
R4464 GND.n3517 GND.n2116 163.367
R4465 GND.n3517 GND.n2124 163.367
R4466 GND.n3179 GND.n2124 163.367
R4467 GND.n3523 GND.n3179 163.367
R4468 GND.n3523 GND.n3180 163.367
R4469 GND.n3180 GND.n2136 163.367
R4470 GND.n3565 GND.n2136 163.367
R4471 GND.n3565 GND.n2144 163.367
R4472 GND.n3569 GND.n2144 163.367
R4473 GND.n3570 GND.n3569 163.367
R4474 GND.n3571 GND.n3570 163.367
R4475 GND.n3571 GND.n2156 163.367
R4476 GND.n3577 GND.n2156 163.367
R4477 GND.n3577 GND.n2164 163.367
R4478 GND.n3147 GND.n2164 163.367
R4479 GND.n3599 GND.n3147 163.367
R4480 GND.n3600 GND.n3599 163.367
R4481 GND.n3600 GND.n2176 163.367
R4482 GND.n3611 GND.n2176 163.367
R4483 GND.n3611 GND.n2183 163.367
R4484 GND.n3607 GND.n2183 163.367
R4485 GND.n3607 GND.n3138 163.367
R4486 GND.n3603 GND.n3138 163.367
R4487 GND.n3603 GND.n2194 163.367
R4488 GND.n3661 GND.n2194 163.367
R4489 GND.n3661 GND.n2202 163.367
R4490 GND.n3131 GND.n2202 163.367
R4491 GND.n3669 GND.n3131 163.367
R4492 GND.n3669 GND.n3132 163.367
R4493 GND.n3665 GND.n3132 163.367
R4494 GND.n3665 GND.n3125 163.367
R4495 GND.n3681 GND.n3125 163.367
R4496 GND.n3681 GND.n2224 163.367
R4497 GND.n3685 GND.n2224 163.367
R4498 GND.n3685 GND.n2232 163.367
R4499 GND.n3123 GND.n2232 163.367
R4500 GND.n3696 GND.n3123 163.367
R4501 GND.n3696 GND.n2249 163.367
R4502 GND.n3692 GND.n2249 163.367
R4503 GND.n3692 GND.n2258 163.367
R4504 GND.n3113 GND.n2258 163.367
R4505 GND.n3720 GND.n3113 163.367
R4506 GND.n3721 GND.n3720 163.367
R4507 GND.n3722 GND.n3721 163.367
R4508 GND.n3722 GND.n3111 163.367
R4509 GND.n3745 GND.n3111 163.367
R4510 GND.n3745 GND.n2294 163.367
R4511 GND.n3741 GND.n2294 163.367
R4512 GND.n3741 GND.n2301 163.367
R4513 GND.n3736 GND.n2301 163.367
R4514 GND.n3736 GND.n3732 163.367
R4515 GND.n3732 GND.n2317 163.367
R4516 GND.n3728 GND.n2317 163.367
R4517 GND.n3728 GND.n2325 163.367
R4518 GND.n3099 GND.n2325 163.367
R4519 GND.n3781 GND.n3099 163.367
R4520 GND.n3782 GND.n3781 163.367
R4521 GND.n3783 GND.n3782 163.367
R4522 GND.n3783 GND.n3097 163.367
R4523 GND.n3792 GND.n3097 163.367
R4524 GND.n3792 GND.n2360 163.367
R4525 GND.n3788 GND.n2360 163.367
R4526 GND.n3788 GND.n2368 163.367
R4527 GND.n3892 GND.n2368 163.367
R4528 GND.n3893 GND.n3892 163.367
R4529 GND.n3893 GND.n3029 163.367
R4530 GND.n3337 GND.n3322 163.367
R4531 GND.n3341 GND.n3322 163.367
R4532 GND.n3345 GND.n3343 163.367
R4533 GND.n3349 GND.n3320 163.367
R4534 GND.n3353 GND.n3351 163.367
R4535 GND.n3357 GND.n3318 163.367
R4536 GND.n3361 GND.n3359 163.367
R4537 GND.n3365 GND.n3316 163.367
R4538 GND.n3369 GND.n3367 163.367
R4539 GND.n3373 GND.n3314 163.367
R4540 GND.n3377 GND.n3375 163.367
R4541 GND.n3381 GND.n3312 163.367
R4542 GND.n3385 GND.n3383 163.367
R4543 GND.n3389 GND.n3307 163.367
R4544 GND.n3392 GND.n3391 163.367
R4545 GND.n3396 GND.n3394 163.367
R4546 GND.n3400 GND.n3305 163.367
R4547 GND.n3404 GND.n3402 163.367
R4548 GND.n3408 GND.n3300 163.367
R4549 GND.n3412 GND.n3410 163.367
R4550 GND.n3416 GND.n3298 163.367
R4551 GND.n3420 GND.n3418 163.367
R4552 GND.n3424 GND.n3296 163.367
R4553 GND.n3428 GND.n3426 163.367
R4554 GND.n3432 GND.n3294 163.367
R4555 GND.n3436 GND.n3434 163.367
R4556 GND.n3440 GND.n3292 163.367
R4557 GND.n3444 GND.n3442 163.367
R4558 GND.n3448 GND.n3290 163.367
R4559 GND.n3451 GND.n3450 163.367
R4560 GND.n4621 GND.n2064 163.367
R4561 GND.n4621 GND.n2065 163.367
R4562 GND.n4617 GND.n2065 163.367
R4563 GND.n4617 GND.n2068 163.367
R4564 GND.n2083 GND.n2068 163.367
R4565 GND.n4606 GND.n2083 163.367
R4566 GND.n4606 GND.n2084 163.367
R4567 GND.n4602 GND.n2084 163.367
R4568 GND.n4602 GND.n2087 163.367
R4569 GND.n3497 GND.n2087 163.367
R4570 GND.n3497 GND.n3490 163.367
R4571 GND.n3493 GND.n3490 163.367
R4572 GND.n3493 GND.n3492 163.367
R4573 GND.n3492 GND.n2118 163.367
R4574 GND.n4585 GND.n2118 163.367
R4575 GND.n4585 GND.n2119 163.367
R4576 GND.n4581 GND.n2119 163.367
R4577 GND.n4581 GND.n2122 163.367
R4578 GND.n3525 GND.n2122 163.367
R4579 GND.n3525 GND.n2138 163.367
R4580 GND.n4571 GND.n2138 163.367
R4581 GND.n4571 GND.n2139 163.367
R4582 GND.n4567 GND.n2139 163.367
R4583 GND.n4567 GND.n2142 163.367
R4584 GND.n3158 GND.n2142 163.367
R4585 GND.n3158 GND.n2158 163.367
R4586 GND.n4557 GND.n2158 163.367
R4587 GND.n4557 GND.n2159 163.367
R4588 GND.n4553 GND.n2159 163.367
R4589 GND.n4553 GND.n2162 163.367
R4590 GND.n3597 GND.n2162 163.367
R4591 GND.n3597 GND.n2178 163.367
R4592 GND.n4543 GND.n2178 163.367
R4593 GND.n4543 GND.n2179 163.367
R4594 GND.n4539 GND.n2179 163.367
R4595 GND.n4539 GND.n2182 163.367
R4596 GND.n3632 GND.n2182 163.367
R4597 GND.n3632 GND.n2196 163.367
R4598 GND.n4529 GND.n2196 163.367
R4599 GND.n4529 GND.n2197 163.367
R4600 GND.n4525 GND.n2197 163.367
R4601 GND.n4525 GND.n2200 163.367
R4602 GND.n3672 GND.n2200 163.367
R4603 GND.n3673 GND.n3672 163.367
R4604 GND.n3673 GND.n3127 163.367
R4605 GND.n3677 GND.n3127 163.367
R4606 GND.n3677 GND.n2226 163.367
R4607 GND.n4508 GND.n2226 163.367
R4608 GND.n4508 GND.n2227 163.367
R4609 GND.n4504 GND.n2227 163.367
R4610 GND.n4504 GND.n2230 163.367
R4611 GND.n2252 GND.n2230 163.367
R4612 GND.n4495 GND.n2252 163.367
R4613 GND.n4495 GND.n2253 163.367
R4614 GND.n4491 GND.n2253 163.367
R4615 GND.n4491 GND.n2256 163.367
R4616 GND.n3718 GND.n2256 163.367
R4617 GND.n3718 GND.n3711 163.367
R4618 GND.n3714 GND.n3711 163.367
R4619 GND.n3714 GND.n3713 163.367
R4620 GND.n3713 GND.n2295 163.367
R4621 GND.n4474 GND.n2295 163.367
R4622 GND.n4474 GND.n2296 163.367
R4623 GND.n4470 GND.n2296 163.367
R4624 GND.n4470 GND.n2299 163.367
R4625 GND.n2319 GND.n2299 163.367
R4626 GND.n4460 GND.n2319 163.367
R4627 GND.n4460 GND.n2320 163.367
R4628 GND.n4456 GND.n2320 163.367
R4629 GND.n4456 GND.n2323 163.367
R4630 GND.n3779 GND.n2323 163.367
R4631 GND.n3779 GND.n3770 163.367
R4632 GND.n3775 GND.n3770 163.367
R4633 GND.n3775 GND.n3774 163.367
R4634 GND.n3774 GND.n2362 163.367
R4635 GND.n4439 GND.n2362 163.367
R4636 GND.n4439 GND.n2363 163.367
R4637 GND.n4435 GND.n2363 163.367
R4638 GND.n4435 GND.n2366 163.367
R4639 GND.n3031 GND.n2366 163.367
R4640 GND.n4004 GND.n3031 163.367
R4641 GND.n1326 GND.n1281 161.3
R4642 GND.n1325 GND.n1324 161.3
R4643 GND.n1323 GND.n1282 161.3
R4644 GND.n1322 GND.n1321 161.3
R4645 GND.n1320 GND.n1283 161.3
R4646 GND.n1319 GND.n1318 161.3
R4647 GND.n1317 GND.n1316 161.3
R4648 GND.n1315 GND.n1285 161.3
R4649 GND.n1314 GND.n1313 161.3
R4650 GND.n1312 GND.n1286 161.3
R4651 GND.n1311 GND.n1310 161.3
R4652 GND.n1309 GND.n1287 161.3
R4653 GND.n1308 GND.n1307 161.3
R4654 GND.n1306 GND.n1305 161.3
R4655 GND.n1304 GND.n1289 161.3
R4656 GND.n1303 GND.n1302 161.3
R4657 GND.n1301 GND.n1290 161.3
R4658 GND.n1300 GND.n1299 161.3
R4659 GND.n1298 GND.n1291 161.3
R4660 GND.n1359 GND.n1270 161.3
R4661 GND.n1358 GND.n1357 161.3
R4662 GND.n1356 GND.n1271 161.3
R4663 GND.n1355 GND.n1354 161.3
R4664 GND.n1353 GND.n1272 161.3
R4665 GND.n1352 GND.n1351 161.3
R4666 GND.n1350 GND.n1349 161.3
R4667 GND.n1348 GND.n1274 161.3
R4668 GND.n1347 GND.n1346 161.3
R4669 GND.n1345 GND.n1275 161.3
R4670 GND.n1344 GND.n1343 161.3
R4671 GND.n1342 GND.n1276 161.3
R4672 GND.n1341 GND.n1340 161.3
R4673 GND.n1339 GND.n1338 161.3
R4674 GND.n1337 GND.n1278 161.3
R4675 GND.n1336 GND.n1335 161.3
R4676 GND.n1334 GND.n1279 161.3
R4677 GND.n1333 GND.n1332 161.3
R4678 GND.n1331 GND.n1280 161.3
R4679 GND.n1392 GND.n1259 161.3
R4680 GND.n1391 GND.n1390 161.3
R4681 GND.n1389 GND.n1260 161.3
R4682 GND.n1388 GND.n1387 161.3
R4683 GND.n1386 GND.n1261 161.3
R4684 GND.n1385 GND.n1384 161.3
R4685 GND.n1383 GND.n1382 161.3
R4686 GND.n1381 GND.n1263 161.3
R4687 GND.n1380 GND.n1379 161.3
R4688 GND.n1378 GND.n1264 161.3
R4689 GND.n1377 GND.n1376 161.3
R4690 GND.n1375 GND.n1265 161.3
R4691 GND.n1374 GND.n1373 161.3
R4692 GND.n1372 GND.n1371 161.3
R4693 GND.n1370 GND.n1267 161.3
R4694 GND.n1369 GND.n1368 161.3
R4695 GND.n1367 GND.n1268 161.3
R4696 GND.n1366 GND.n1365 161.3
R4697 GND.n1364 GND.n1269 161.3
R4698 GND.n1425 GND.n1248 161.3
R4699 GND.n1424 GND.n1423 161.3
R4700 GND.n1422 GND.n1249 161.3
R4701 GND.n1421 GND.n1420 161.3
R4702 GND.n1419 GND.n1250 161.3
R4703 GND.n1418 GND.n1417 161.3
R4704 GND.n1416 GND.n1415 161.3
R4705 GND.n1414 GND.n1252 161.3
R4706 GND.n1413 GND.n1412 161.3
R4707 GND.n1411 GND.n1253 161.3
R4708 GND.n1410 GND.n1409 161.3
R4709 GND.n1408 GND.n1254 161.3
R4710 GND.n1407 GND.n1406 161.3
R4711 GND.n1405 GND.n1404 161.3
R4712 GND.n1403 GND.n1256 161.3
R4713 GND.n1402 GND.n1401 161.3
R4714 GND.n1400 GND.n1257 161.3
R4715 GND.n1399 GND.n1398 161.3
R4716 GND.n1397 GND.n1258 161.3
R4717 GND.n2755 GND.n2754 161.3
R4718 GND.n2756 GND.n2751 161.3
R4719 GND.n2758 GND.n2757 161.3
R4720 GND.n2759 GND.n2750 161.3
R4721 GND.n2761 GND.n2760 161.3
R4722 GND.n2763 GND.n2749 161.3
R4723 GND.n2765 GND.n2764 161.3
R4724 GND.n2766 GND.n2748 161.3
R4725 GND.n2768 GND.n2767 161.3
R4726 GND.n2769 GND.n2747 161.3
R4727 GND.n2772 GND.n2771 161.3
R4728 GND.n2773 GND.n2746 161.3
R4729 GND.n2775 GND.n2774 161.3
R4730 GND.n2776 GND.n2745 161.3
R4731 GND.n2720 GND.n2719 161.3
R4732 GND.n2721 GND.n2716 161.3
R4733 GND.n2723 GND.n2722 161.3
R4734 GND.n2724 GND.n2715 161.3
R4735 GND.n2726 GND.n2725 161.3
R4736 GND.n2728 GND.n2714 161.3
R4737 GND.n2730 GND.n2729 161.3
R4738 GND.n2731 GND.n2713 161.3
R4739 GND.n2733 GND.n2732 161.3
R4740 GND.n2734 GND.n2712 161.3
R4741 GND.n2737 GND.n2736 161.3
R4742 GND.n2738 GND.n2711 161.3
R4743 GND.n2740 GND.n2739 161.3
R4744 GND.n2741 GND.n2710 161.3
R4745 GND.n2685 GND.n2684 161.3
R4746 GND.n2686 GND.n2681 161.3
R4747 GND.n2688 GND.n2687 161.3
R4748 GND.n2689 GND.n2680 161.3
R4749 GND.n2691 GND.n2690 161.3
R4750 GND.n2693 GND.n2679 161.3
R4751 GND.n2695 GND.n2694 161.3
R4752 GND.n2696 GND.n2678 161.3
R4753 GND.n2698 GND.n2697 161.3
R4754 GND.n2699 GND.n2677 161.3
R4755 GND.n2702 GND.n2701 161.3
R4756 GND.n2703 GND.n2676 161.3
R4757 GND.n2705 GND.n2704 161.3
R4758 GND.n2706 GND.n2675 161.3
R4759 GND.n2651 GND.n2650 161.3
R4760 GND.n2652 GND.n2647 161.3
R4761 GND.n2654 GND.n2653 161.3
R4762 GND.n2655 GND.n2646 161.3
R4763 GND.n2657 GND.n2656 161.3
R4764 GND.n2659 GND.n2645 161.3
R4765 GND.n2661 GND.n2660 161.3
R4766 GND.n2662 GND.n2644 161.3
R4767 GND.n2664 GND.n2663 161.3
R4768 GND.n2665 GND.n2643 161.3
R4769 GND.n2668 GND.n2667 161.3
R4770 GND.n2669 GND.n2642 161.3
R4771 GND.n2671 GND.n2670 161.3
R4772 GND.n2672 GND.n2641 161.3
R4773 GND.n2637 GND.n2606 161.3
R4774 GND.n2636 GND.n2635 161.3
R4775 GND.n2634 GND.n2607 161.3
R4776 GND.n2633 GND.n2632 161.3
R4777 GND.n2630 GND.n2608 161.3
R4778 GND.n2629 GND.n2628 161.3
R4779 GND.n2627 GND.n2609 161.3
R4780 GND.n2626 GND.n2625 161.3
R4781 GND.n2624 GND.n2610 161.3
R4782 GND.n2622 GND.n2621 161.3
R4783 GND.n2620 GND.n2611 161.3
R4784 GND.n2619 GND.n2618 161.3
R4785 GND.n2617 GND.n2612 161.3
R4786 GND.n2616 GND.n2615 161.3
R4787 GND.n2602 GND.n2571 161.3
R4788 GND.n2601 GND.n2600 161.3
R4789 GND.n2599 GND.n2572 161.3
R4790 GND.n2598 GND.n2597 161.3
R4791 GND.n2595 GND.n2573 161.3
R4792 GND.n2594 GND.n2593 161.3
R4793 GND.n2592 GND.n2574 161.3
R4794 GND.n2591 GND.n2590 161.3
R4795 GND.n2589 GND.n2575 161.3
R4796 GND.n2587 GND.n2586 161.3
R4797 GND.n2585 GND.n2576 161.3
R4798 GND.n2584 GND.n2583 161.3
R4799 GND.n2582 GND.n2577 161.3
R4800 GND.n2581 GND.n2580 161.3
R4801 GND.n2567 GND.n2536 161.3
R4802 GND.n2566 GND.n2565 161.3
R4803 GND.n2564 GND.n2537 161.3
R4804 GND.n2563 GND.n2562 161.3
R4805 GND.n2560 GND.n2538 161.3
R4806 GND.n2559 GND.n2558 161.3
R4807 GND.n2557 GND.n2539 161.3
R4808 GND.n2556 GND.n2555 161.3
R4809 GND.n2554 GND.n2540 161.3
R4810 GND.n2552 GND.n2551 161.3
R4811 GND.n2550 GND.n2541 161.3
R4812 GND.n2549 GND.n2548 161.3
R4813 GND.n2547 GND.n2542 161.3
R4814 GND.n2546 GND.n2545 161.3
R4815 GND.n2533 GND.n2502 161.3
R4816 GND.n2532 GND.n2531 161.3
R4817 GND.n2530 GND.n2503 161.3
R4818 GND.n2529 GND.n2528 161.3
R4819 GND.n2526 GND.n2504 161.3
R4820 GND.n2525 GND.n2524 161.3
R4821 GND.n2523 GND.n2505 161.3
R4822 GND.n2522 GND.n2521 161.3
R4823 GND.n2520 GND.n2506 161.3
R4824 GND.n2518 GND.n2517 161.3
R4825 GND.n2516 GND.n2507 161.3
R4826 GND.n2515 GND.n2514 161.3
R4827 GND.n2513 GND.n2508 161.3
R4828 GND.n2512 GND.n2511 161.3
R4829 GND.n3042 GND.n3041 155.685
R4830 GND.n2501 GND.t109 154.006
R4831 GND.n3330 GND.n3323 152
R4832 GND.n3332 GND.n3331 152
R4833 GND.n3040 GND.n3034 152
R4834 GND.n50 GND.t27 151.613
R4835 GND.n61 GND.t23 151.613
R4836 GND.n26 GND.t18 151.613
R4837 GND.n37 GND.t26 151.613
R4838 GND.n3 GND.t11 151.613
R4839 GND.n14 GND.t124 151.613
R4840 GND.n133 GND.t31 151.613
R4841 GND.n122 GND.t21 151.613
R4842 GND.n109 GND.t30 151.613
R4843 GND.n98 GND.t126 151.613
R4844 GND.n86 GND.t127 151.613
R4845 GND.n75 GND.t24 151.613
R4846 GND.n3038 GND.t44 151.333
R4847 GND.n1443 GND.t6 149.525
R4848 GND.n2479 GND.t13 149.525
R4849 GND.n1221 GND.t33 149.525
R4850 GND.n2444 GND.t34 149.525
R4851 GND.n2501 GND.t114 144.651
R4852 GND.n3949 GND.n3948 143.351
R4853 GND.n3948 GND.n3947 143.351
R4854 GND.n3328 GND.t86 131.925
R4855 GND.n3331 GND.t102 126.766
R4856 GND.n3329 GND.t47 126.766
R4857 GND.n3039 GND.t99 126.766
R4858 GND.n3041 GND.t69 126.766
R4859 GND.n1472 GND.t94 124.445
R4860 GND.n1187 GND.t57 124.445
R4861 GND.n1203 GND.t68 124.445
R4862 GND.n2409 GND.t119 124.445
R4863 GND.n2421 GND.t38 124.445
R4864 GND.n305 GND.t82 124.445
R4865 GND.n5776 GND.t75 124.445
R4866 GND.n4220 GND.t123 124.445
R4867 GND.n2378 GND.t84 124.445
R4868 GND.n1025 GND.t106 124.445
R4869 GND.n1017 GND.t97 124.445
R4870 GND.n4786 GND.t111 124.445
R4871 GND.n1247 GND.t65 108.153
R4872 GND.n1396 GND.n1395 107.957
R4873 GND.n1427 GND.n1426 107.957
R4874 GND.n1363 GND.n1362 107.957
R4875 GND.n1394 GND.n1393 107.957
R4876 GND.n1330 GND.n1329 107.957
R4877 GND.n1361 GND.n1360 107.957
R4878 GND.n1297 GND.n1296 107.957
R4879 GND.n1328 GND.n1327 107.957
R4880 GND.n1294 GND.t59 107.198
R4881 GND.n53 GND.n52 104.615
R4882 GND.n64 GND.n63 104.615
R4883 GND.n29 GND.n28 104.615
R4884 GND.n40 GND.n39 104.615
R4885 GND.n6 GND.n5 104.615
R4886 GND.n17 GND.n16 104.615
R4887 GND.n1463 GND.n1433 104.615
R4888 GND.n1456 GND.n1433 104.615
R4889 GND.n1456 GND.n1455 104.615
R4890 GND.n1455 GND.n1437 104.615
R4891 GND.n1448 GND.n1437 104.615
R4892 GND.n1448 GND.n1447 104.615
R4893 GND.n1447 GND.n1441 104.615
R4894 GND.n1225 GND.n1219 104.615
R4895 GND.n1226 GND.n1225 104.615
R4896 GND.n1226 GND.n1215 104.615
R4897 GND.n1233 GND.n1215 104.615
R4898 GND.n1234 GND.n1233 104.615
R4899 GND.n1234 GND.n1211 104.615
R4900 GND.n1241 GND.n1211 104.615
R4901 GND.n136 GND.n135 104.615
R4902 GND.n125 GND.n124 104.615
R4903 GND.n112 GND.n111 104.615
R4904 GND.n101 GND.n100 104.615
R4905 GND.n89 GND.n88 104.615
R4906 GND.n78 GND.n77 104.615
R4907 GND.n2499 GND.n2469 104.615
R4908 GND.n2492 GND.n2469 104.615
R4909 GND.n2492 GND.n2491 104.615
R4910 GND.n2491 GND.n2473 104.615
R4911 GND.n2484 GND.n2473 104.615
R4912 GND.n2484 GND.n2483 104.615
R4913 GND.n2483 GND.n2477 104.615
R4914 GND.n2448 GND.n2442 104.615
R4915 GND.n2449 GND.n2448 104.615
R4916 GND.n2449 GND.n2438 104.615
R4917 GND.n2456 GND.n2438 104.615
R4918 GND.n2457 GND.n2456 104.615
R4919 GND.n2457 GND.n2434 104.615
R4920 GND.n2464 GND.n2434 104.615
R4921 GND.n1472 GND.n1471 102.013
R4922 GND.n1187 GND.n1186 102.013
R4923 GND.n1203 GND.n1202 102.013
R4924 GND.n2409 GND.n2408 102.013
R4925 GND.n2421 GND.n2420 102.013
R4926 GND.n305 GND.n304 102.013
R4927 GND.n5776 GND.n5775 102.013
R4928 GND.n4220 GND.n4219 102.013
R4929 GND.n2378 GND.n2377 102.013
R4930 GND.n1025 GND.n1024 102.013
R4931 GND.n1017 GND.n1016 102.013
R4932 GND.n4786 GND.n4785 102.013
R4933 GND.n5789 GND.n5788 99.6594
R4934 GND.n5784 GND.n286 99.6594
R4935 GND.n5780 GND.n285 99.6594
R4936 GND.n5773 GND.n284 99.6594
R4937 GND.n5769 GND.n283 99.6594
R4938 GND.n5765 GND.n282 99.6594
R4939 GND.n5761 GND.n281 99.6594
R4940 GND.n5757 GND.n280 99.6594
R4941 GND.n308 GND.n279 99.6594
R4942 GND.n4424 GND.n4423 99.6594
R4943 GND.n4418 GND.n2383 99.6594
R4944 GND.n4415 GND.n2384 99.6594
R4945 GND.n4410 GND.n2386 99.6594
R4946 GND.n4406 GND.n2387 99.6594
R4947 GND.n4402 GND.n2388 99.6594
R4948 GND.n4398 GND.n2389 99.6594
R4949 GND.n2419 GND.n2390 99.6594
R4950 GND.n4230 GND.n274 99.6594
R4951 GND.n4234 GND.n275 99.6594
R4952 GND.n4239 GND.n276 99.6594
R4953 GND.n4242 GND.n277 99.6594
R4954 GND.n2802 GND.n2391 99.6594
R4955 GND.n2798 GND.n2392 99.6594
R4956 GND.n2794 GND.n2393 99.6594
R4957 GND.n2790 GND.n2394 99.6594
R4958 GND.n4650 GND.n1181 99.6594
R4959 GND.n4649 GND.n1184 99.6594
R4960 GND.n4646 GND.n1191 99.6594
R4961 GND.n4645 GND.n1194 99.6594
R4962 GND.n4643 GND.n1196 99.6594
R4963 GND.n4642 GND.n1199 99.6594
R4964 GND.n4640 GND.n1201 99.6594
R4965 GND.n4639 GND.n1169 99.6594
R4966 GND.n997 GND.n966 99.6594
R4967 GND.n1033 GND.n967 99.6594
R4968 GND.n1041 GND.n968 99.6594
R4969 GND.n1043 GND.n969 99.6594
R4970 GND.n1051 GND.n970 99.6594
R4971 GND.n1055 GND.n971 99.6594
R4972 GND.n1061 GND.n972 99.6594
R4973 GND.n1065 GND.n973 99.6594
R4974 GND.n1020 GND.n974 99.6594
R4975 GND.n3872 GND.n3817 99.6594
R4976 GND.n3870 GND.n3816 99.6594
R4977 GND.n3866 GND.n3815 99.6594
R4978 GND.n3862 GND.n3814 99.6594
R4979 GND.n3858 GND.n3813 99.6594
R4980 GND.n3854 GND.n3812 99.6594
R4981 GND.n3850 GND.n3811 99.6594
R4982 GND.n3846 GND.n3810 99.6594
R4983 GND.n3842 GND.n3809 99.6594
R4984 GND.n3808 GND.n3807 99.6594
R4985 GND.n3882 GND.n3091 99.6594
R4986 GND.n3277 GND.n3276 99.6594
R4987 GND.n3271 GND.n3200 99.6594
R4988 GND.n3268 GND.n3201 99.6594
R4989 GND.n3264 GND.n3202 99.6594
R4990 GND.n3260 GND.n3203 99.6594
R4991 GND.n3256 GND.n3204 99.6594
R4992 GND.n3252 GND.n3205 99.6594
R4993 GND.n3248 GND.n3206 99.6594
R4994 GND.n3244 GND.n3207 99.6594
R4995 GND.n3240 GND.n3208 99.6594
R4996 GND.n3279 GND.n3199 99.6594
R4997 GND.n3277 GND.n3211 99.6594
R4998 GND.n3269 GND.n3200 99.6594
R4999 GND.n3265 GND.n3201 99.6594
R5000 GND.n3261 GND.n3202 99.6594
R5001 GND.n3257 GND.n3203 99.6594
R5002 GND.n3253 GND.n3204 99.6594
R5003 GND.n3249 GND.n3205 99.6594
R5004 GND.n3245 GND.n3206 99.6594
R5005 GND.n3241 GND.n3207 99.6594
R5006 GND.n3237 GND.n3208 99.6594
R5007 GND.n3280 GND.n3279 99.6594
R5008 GND.n3883 GND.n3882 99.6594
R5009 GND.n3841 GND.n3808 99.6594
R5010 GND.n3845 GND.n3809 99.6594
R5011 GND.n3849 GND.n3810 99.6594
R5012 GND.n3853 GND.n3811 99.6594
R5013 GND.n3857 GND.n3812 99.6594
R5014 GND.n3861 GND.n3813 99.6594
R5015 GND.n3865 GND.n3814 99.6594
R5016 GND.n3869 GND.n3815 99.6594
R5017 GND.n3873 GND.n3816 99.6594
R5018 GND.n3818 GND.n3817 99.6594
R5019 GND.n1034 GND.n966 99.6594
R5020 GND.n1040 GND.n967 99.6594
R5021 GND.n1044 GND.n968 99.6594
R5022 GND.n1050 GND.n969 99.6594
R5023 GND.n1054 GND.n970 99.6594
R5024 GND.n1060 GND.n971 99.6594
R5025 GND.n1064 GND.n972 99.6594
R5026 GND.n1019 GND.n973 99.6594
R5027 GND.n1015 GND.n974 99.6594
R5028 GND.n4639 GND.n4638 99.6594
R5029 GND.n4640 GND.n1200 99.6594
R5030 GND.n4642 GND.n4641 99.6594
R5031 GND.n4643 GND.n1195 99.6594
R5032 GND.n4645 GND.n4644 99.6594
R5033 GND.n4647 GND.n1185 99.6594
R5034 GND.n4649 GND.n4648 99.6594
R5035 GND.n4650 GND.n1180 99.6594
R5036 GND.n2799 GND.n2391 99.6594
R5037 GND.n2795 GND.n2392 99.6594
R5038 GND.n2791 GND.n2393 99.6594
R5039 GND.n2394 GND.n2380 99.6594
R5040 GND.n4221 GND.n277 99.6594
R5041 GND.n4233 GND.n276 99.6594
R5042 GND.n4231 GND.n275 99.6594
R5043 GND.n4225 GND.n274 99.6594
R5044 GND.n4424 GND.n2397 99.6594
R5045 GND.n4416 GND.n2383 99.6594
R5046 GND.n4411 GND.n2385 99.6594
R5047 GND.n4407 GND.n2386 99.6594
R5048 GND.n4403 GND.n2387 99.6594
R5049 GND.n4399 GND.n2388 99.6594
R5050 GND.n2418 GND.n2389 99.6594
R5051 GND.n4391 GND.n2390 99.6594
R5052 GND.n5756 GND.n279 99.6594
R5053 GND.n5760 GND.n280 99.6594
R5054 GND.n5764 GND.n281 99.6594
R5055 GND.n5768 GND.n282 99.6594
R5056 GND.n5772 GND.n283 99.6594
R5057 GND.n5779 GND.n284 99.6594
R5058 GND.n5783 GND.n285 99.6594
R5059 GND.n287 GND.n286 99.6594
R5060 GND.n5789 GND.n271 99.6594
R5061 GND.n982 GND.n976 99.6594
R5062 GND.n987 GND.n977 99.6594
R5063 GND.n989 GND.n978 99.6594
R5064 GND.n4784 GND.n979 99.6594
R5065 GND.n986 GND.n976 99.6594
R5066 GND.n988 GND.n977 99.6594
R5067 GND.n4783 GND.n978 99.6594
R5068 GND.n4781 GND.n979 99.6594
R5069 GND.n1479 GND.n1206 99.6594
R5070 GND.n1481 GND.n1208 99.6594
R5071 GND.n1482 GND.n1468 99.6594
R5072 GND.n1483 GND.n1470 99.6594
R5073 GND.n1483 GND.n1477 99.6594
R5074 GND.n1482 GND.n1469 99.6594
R5075 GND.n1481 GND.n1480 99.6594
R5076 GND.n1479 GND.n1207 99.6594
R5077 GND.n2778 GND.n2777 89.6708
R5078 GND.n2743 GND.n2742 89.6708
R5079 GND.n2708 GND.n2707 89.6708
R5080 GND.n2674 GND.n2673 89.6708
R5081 GND.n2639 GND.n2638 89.6708
R5082 GND.n2604 GND.n2603 89.6708
R5083 GND.n2569 GND.n2568 89.6708
R5084 GND.n2535 GND.n2534 89.6708
R5085 GND.n1246 GND.t58 85.6032
R5086 GND.n1292 GND.t64 85.6032
R5087 GND.n1293 GND.t108 85.6032
R5088 GND.n1429 GND.t113 85.6032
R5089 GND.n4971 GND.n4970 80.7937
R5090 GND.n4970 GND.n800 80.7937
R5091 GND.n4964 GND.n800 80.7937
R5092 GND.n4964 GND.n4963 80.7937
R5093 GND.n4963 GND.n4962 80.7937
R5094 GND.n4962 GND.n808 80.7937
R5095 GND.n4956 GND.n808 80.7937
R5096 GND.n4956 GND.n4955 80.7937
R5097 GND.n4955 GND.n4954 80.7937
R5098 GND.n4954 GND.n816 80.7937
R5099 GND.n4948 GND.n816 80.7937
R5100 GND.n4948 GND.n4947 80.7937
R5101 GND.n4947 GND.n4946 80.7937
R5102 GND.n4946 GND.n824 80.7937
R5103 GND.n4940 GND.n824 80.7937
R5104 GND.n4940 GND.n4939 80.7937
R5105 GND.n4939 GND.n4938 80.7937
R5106 GND.n4938 GND.n832 80.7937
R5107 GND.n4932 GND.n832 80.7937
R5108 GND.n4932 GND.n4931 80.7937
R5109 GND.n4931 GND.n4930 80.7937
R5110 GND.n4930 GND.n840 80.7937
R5111 GND.n4924 GND.n840 80.7937
R5112 GND.n4924 GND.n4923 80.7937
R5113 GND.n4923 GND.n4922 80.7937
R5114 GND.n4922 GND.n848 80.7937
R5115 GND.n4916 GND.n848 80.7937
R5116 GND.n4916 GND.n4915 80.7937
R5117 GND.n4915 GND.n4914 80.7937
R5118 GND.n4914 GND.n856 80.7937
R5119 GND.n4908 GND.n856 80.7937
R5120 GND.n4908 GND.n4907 80.7937
R5121 GND.n4907 GND.n4906 80.7937
R5122 GND.n4906 GND.n864 80.7937
R5123 GND.n4900 GND.n864 80.7937
R5124 GND.n4900 GND.n4899 80.7937
R5125 GND.n4899 GND.n4898 80.7937
R5126 GND.n4898 GND.n872 80.7937
R5127 GND.n4892 GND.n872 80.7937
R5128 GND.n4892 GND.n4891 80.7937
R5129 GND.n4891 GND.n4890 80.7937
R5130 GND.n4890 GND.n880 80.7937
R5131 GND.n4884 GND.n880 80.7937
R5132 GND.n4884 GND.n4883 80.7937
R5133 GND.n4883 GND.n4882 80.7937
R5134 GND.n4882 GND.n888 80.7937
R5135 GND.n4876 GND.n888 80.7937
R5136 GND.n4876 GND.n4875 80.7937
R5137 GND.n4875 GND.n4874 80.7937
R5138 GND.n4874 GND.n896 80.7937
R5139 GND.n4868 GND.n896 80.7937
R5140 GND.n4868 GND.n4867 80.7937
R5141 GND.n4867 GND.n4866 80.7937
R5142 GND.n3328 GND.n3327 80.3738
R5143 GND.n2753 GND.t148 75.0788
R5144 GND.n2718 GND.t133 75.0788
R5145 GND.n2683 GND.t169 75.0788
R5146 GND.n2649 GND.t134 75.0788
R5147 GND.n2614 GND.t141 75.0788
R5148 GND.n2579 GND.t129 75.0788
R5149 GND.n2544 GND.t183 75.0788
R5150 GND.n2510 GND.t143 75.0788
R5151 GND.n3329 GND.n3324 72.8411
R5152 GND.n3999 GND.n3044 71.676
R5153 GND.n3997 GND.n3996 71.676
R5154 GND.n3992 GND.n3047 71.676
R5155 GND.n3990 GND.n3989 71.676
R5156 GND.n3985 GND.n3050 71.676
R5157 GND.n3983 GND.n3982 71.676
R5158 GND.n3978 GND.n3053 71.676
R5159 GND.n3976 GND.n3975 71.676
R5160 GND.n3971 GND.n3056 71.676
R5161 GND.n3969 GND.n3968 71.676
R5162 GND.n3964 GND.n3059 71.676
R5163 GND.n3962 GND.n3961 71.676
R5164 GND.n3956 GND.n3064 71.676
R5165 GND.n3954 GND.n3953 71.676
R5166 GND.n3947 GND.n3946 71.676
R5167 GND.n3942 GND.n3067 71.676
R5168 GND.n3940 GND.n3939 71.676
R5169 GND.n3935 GND.n3073 71.676
R5170 GND.n3933 GND.n3932 71.676
R5171 GND.n3928 GND.n3076 71.676
R5172 GND.n3926 GND.n3925 71.676
R5173 GND.n3921 GND.n3079 71.676
R5174 GND.n3919 GND.n3918 71.676
R5175 GND.n3914 GND.n3082 71.676
R5176 GND.n3912 GND.n3911 71.676
R5177 GND.n3907 GND.n3085 71.676
R5178 GND.n3905 GND.n3904 71.676
R5179 GND.n3900 GND.n3088 71.676
R5180 GND.n3898 GND.n3897 71.676
R5181 GND.n3336 GND.n3335 71.676
R5182 GND.n3342 GND.n3341 71.676
R5183 GND.n3345 GND.n3344 71.676
R5184 GND.n3350 GND.n3349 71.676
R5185 GND.n3353 GND.n3352 71.676
R5186 GND.n3358 GND.n3357 71.676
R5187 GND.n3361 GND.n3360 71.676
R5188 GND.n3366 GND.n3365 71.676
R5189 GND.n3369 GND.n3368 71.676
R5190 GND.n3374 GND.n3373 71.676
R5191 GND.n3377 GND.n3376 71.676
R5192 GND.n3382 GND.n3381 71.676
R5193 GND.n3385 GND.n3384 71.676
R5194 GND.n3390 GND.n3389 71.676
R5195 GND.n3393 GND.n3392 71.676
R5196 GND.n3396 GND.n3395 71.676
R5197 GND.n3401 GND.n3400 71.676
R5198 GND.n3404 GND.n3403 71.676
R5199 GND.n3409 GND.n3408 71.676
R5200 GND.n3412 GND.n3411 71.676
R5201 GND.n3417 GND.n3416 71.676
R5202 GND.n3420 GND.n3419 71.676
R5203 GND.n3425 GND.n3424 71.676
R5204 GND.n3428 GND.n3427 71.676
R5205 GND.n3433 GND.n3432 71.676
R5206 GND.n3436 GND.n3435 71.676
R5207 GND.n3441 GND.n3440 71.676
R5208 GND.n3444 GND.n3443 71.676
R5209 GND.n3449 GND.n3448 71.676
R5210 GND.n3337 GND.n3336 71.676
R5211 GND.n3343 GND.n3342 71.676
R5212 GND.n3344 GND.n3320 71.676
R5213 GND.n3351 GND.n3350 71.676
R5214 GND.n3352 GND.n3318 71.676
R5215 GND.n3359 GND.n3358 71.676
R5216 GND.n3360 GND.n3316 71.676
R5217 GND.n3367 GND.n3366 71.676
R5218 GND.n3368 GND.n3314 71.676
R5219 GND.n3375 GND.n3374 71.676
R5220 GND.n3376 GND.n3312 71.676
R5221 GND.n3383 GND.n3382 71.676
R5222 GND.n3384 GND.n3307 71.676
R5223 GND.n3391 GND.n3390 71.676
R5224 GND.n3394 GND.n3393 71.676
R5225 GND.n3395 GND.n3305 71.676
R5226 GND.n3402 GND.n3401 71.676
R5227 GND.n3403 GND.n3300 71.676
R5228 GND.n3410 GND.n3409 71.676
R5229 GND.n3411 GND.n3298 71.676
R5230 GND.n3418 GND.n3417 71.676
R5231 GND.n3419 GND.n3296 71.676
R5232 GND.n3426 GND.n3425 71.676
R5233 GND.n3427 GND.n3294 71.676
R5234 GND.n3434 GND.n3433 71.676
R5235 GND.n3435 GND.n3292 71.676
R5236 GND.n3442 GND.n3441 71.676
R5237 GND.n3443 GND.n3290 71.676
R5238 GND.n3450 GND.n3449 71.676
R5239 GND.n3899 GND.n3898 71.676
R5240 GND.n3088 GND.n3086 71.676
R5241 GND.n3906 GND.n3905 71.676
R5242 GND.n3085 GND.n3083 71.676
R5243 GND.n3913 GND.n3912 71.676
R5244 GND.n3082 GND.n3080 71.676
R5245 GND.n3920 GND.n3919 71.676
R5246 GND.n3079 GND.n3077 71.676
R5247 GND.n3927 GND.n3926 71.676
R5248 GND.n3076 GND.n3074 71.676
R5249 GND.n3934 GND.n3933 71.676
R5250 GND.n3073 GND.n3068 71.676
R5251 GND.n3941 GND.n3940 71.676
R5252 GND.n3067 GND.n3065 71.676
R5253 GND.n3950 GND.n3949 71.676
R5254 GND.n3955 GND.n3954 71.676
R5255 GND.n3064 GND.n3060 71.676
R5256 GND.n3963 GND.n3962 71.676
R5257 GND.n3059 GND.n3057 71.676
R5258 GND.n3970 GND.n3969 71.676
R5259 GND.n3056 GND.n3054 71.676
R5260 GND.n3977 GND.n3976 71.676
R5261 GND.n3053 GND.n3051 71.676
R5262 GND.n3984 GND.n3983 71.676
R5263 GND.n3050 GND.n3048 71.676
R5264 GND.n3991 GND.n3990 71.676
R5265 GND.n3047 GND.n3045 71.676
R5266 GND.n3998 GND.n3997 71.676
R5267 GND.n3044 GND.n3032 71.676
R5268 GND.n1431 GND.n1245 68.1049
R5269 GND.n1244 GND.n1243 68.088
R5270 GND.n2467 GND.n2466 68.088
R5271 GND.n2784 GND.n2783 67.5474
R5272 GND.n2753 GND.n2752 65.3586
R5273 GND.n2718 GND.n2717 65.3586
R5274 GND.n2683 GND.n2682 65.3586
R5275 GND.n2649 GND.n2648 65.3586
R5276 GND.n2614 GND.n2613 65.3586
R5277 GND.n2579 GND.n2578 65.3586
R5278 GND.n2544 GND.n2543 65.3586
R5279 GND.n2510 GND.n2509 65.3586
R5280 GND.n4858 GND.n904 63.8436
R5281 GND.n5684 GND.n5683 63.8436
R5282 GND.n3333 GND.n3332 59.9562
R5283 GND.n3303 GND.n3302 59.5399
R5284 GND.n3071 GND.n3070 59.5399
R5285 GND.n3310 GND.n3309 59.5399
R5286 GND.n3958 GND.n3062 59.5399
R5287 GND.n2775 GND.n2746 56.4773
R5288 GND.n2740 GND.n2711 56.4773
R5289 GND.n2705 GND.n2676 56.4773
R5290 GND.n2671 GND.n2642 56.4773
R5291 GND.n2636 GND.n2607 56.4773
R5292 GND.n2601 GND.n2572 56.4773
R5293 GND.n2566 GND.n2537 56.4773
R5294 GND.n2532 GND.n2503 56.4773
R5295 GND.n3302 GND.n3301 53.7217
R5296 GND.n3070 GND.n3069 53.7217
R5297 GND.n3309 GND.n3308 53.7217
R5298 GND.n3062 GND.n3061 53.7217
R5299 GND.n2782 GND.n2500 52.3611
R5300 GND.n1244 GND.n1242 52.3452
R5301 GND.n2467 GND.n2465 52.3452
R5302 GND.n52 GND.t27 52.3082
R5303 GND.n63 GND.t23 52.3082
R5304 GND.n28 GND.t18 52.3082
R5305 GND.n39 GND.t26 52.3082
R5306 GND.n5 GND.t11 52.3082
R5307 GND.n16 GND.t124 52.3082
R5308 GND.t6 GND.n1441 52.3082
R5309 GND.t33 GND.n1219 52.3082
R5310 GND.n135 GND.t31 52.3082
R5311 GND.n124 GND.t21 52.3082
R5312 GND.n111 GND.t30 52.3082
R5313 GND.n100 GND.t126 52.3082
R5314 GND.n88 GND.t127 52.3082
R5315 GND.n77 GND.t24 52.3082
R5316 GND.t13 GND.n2477 52.3082
R5317 GND.t34 GND.n2442 52.3082
R5318 GND.n1465 GND.n1464 50.6096
R5319 GND.n3038 GND.n3037 48.9137
R5320 GND.n2764 GND.n2748 48.2005
R5321 GND.n2757 GND.n2750 48.2005
R5322 GND.n2729 GND.n2713 48.2005
R5323 GND.n2722 GND.n2715 48.2005
R5324 GND.n2694 GND.n2678 48.2005
R5325 GND.n2687 GND.n2680 48.2005
R5326 GND.n2660 GND.n2644 48.2005
R5327 GND.n2653 GND.n2646 48.2005
R5328 GND.n2618 GND.n2611 48.2005
R5329 GND.n2625 GND.n2609 48.2005
R5330 GND.n2583 GND.n2576 48.2005
R5331 GND.n2590 GND.n2574 48.2005
R5332 GND.n2548 GND.n2541 48.2005
R5333 GND.n2555 GND.n2539 48.2005
R5334 GND.n2514 GND.n2507 48.2005
R5335 GND.n2521 GND.n2505 48.2005
R5336 GND.n3836 GND.n3835 45.5763
R5337 GND.n3231 GND.n3230 45.5763
R5338 GND.n2777 GND.t167 44.6035
R5339 GND.n2770 GND.t177 44.6035
R5340 GND.n2762 GND.t154 44.6035
R5341 GND.n2752 GND.t161 44.6035
R5342 GND.n2742 GND.t152 44.6035
R5343 GND.n2735 GND.t160 44.6035
R5344 GND.n2727 GND.t136 44.6035
R5345 GND.n2717 GND.t144 44.6035
R5346 GND.n2707 GND.t157 44.6035
R5347 GND.n2700 GND.t140 44.6035
R5348 GND.n2692 GND.t131 44.6035
R5349 GND.n2682 GND.t179 44.6035
R5350 GND.n2673 GND.t176 44.6035
R5351 GND.n2666 GND.t164 44.6035
R5352 GND.n2658 GND.t151 44.6035
R5353 GND.n2648 GND.t139 44.6035
R5354 GND.n2613 GND.t175 44.6035
R5355 GND.n2623 GND.t165 44.6035
R5356 GND.n2631 GND.t135 44.6035
R5357 GND.n2638 GND.t181 44.6035
R5358 GND.n2578 GND.t159 44.6035
R5359 GND.n2588 GND.t147 44.6035
R5360 GND.n2596 GND.t174 44.6035
R5361 GND.n2603 GND.t166 44.6035
R5362 GND.n2543 GND.t155 44.6035
R5363 GND.n2553 GND.t158 44.6035
R5364 GND.n2561 GND.t170 44.6035
R5365 GND.n2568 GND.t128 44.6035
R5366 GND.n2509 GND.t171 44.6035
R5367 GND.n2519 GND.t180 44.6035
R5368 GND.n2527 GND.t137 44.6035
R5369 GND.n2534 GND.t146 44.6035
R5370 GND.n1396 GND.t145 44.4654
R5371 GND.n1255 GND.t156 44.4654
R5372 GND.n1251 GND.t182 44.4654
R5373 GND.n1426 GND.t172 44.4654
R5374 GND.n1363 GND.t150 44.4654
R5375 GND.n1266 GND.t138 44.4654
R5376 GND.n1262 GND.t142 44.4654
R5377 GND.n1393 GND.t132 44.4654
R5378 GND.n1330 GND.t168 44.4654
R5379 GND.n1277 GND.t163 44.4654
R5380 GND.n1273 GND.t178 44.4654
R5381 GND.n1360 GND.t153 44.4654
R5382 GND.n1297 GND.t149 44.4654
R5383 GND.n1288 GND.t162 44.4654
R5384 GND.n1284 GND.t173 44.4654
R5385 GND.n1327 GND.t130 44.4654
R5386 GND.n1402 GND.n1257 44.4521
R5387 GND.n1420 GND.n1249 44.4521
R5388 GND.n1369 GND.n1268 44.4521
R5389 GND.n1387 GND.n1260 44.4521
R5390 GND.n1336 GND.n1279 44.4521
R5391 GND.n1354 GND.n1271 44.4521
R5392 GND.n1303 GND.n1290 44.4521
R5393 GND.n1321 GND.n1282 44.4521
R5394 GND.n4002 GND.n3042 44.3322
R5395 GND.n3329 GND.n3328 42.7233
R5396 GND.n1473 GND.n1472 42.2793
R5397 GND.n1204 GND.n1203 42.2793
R5398 GND.n2422 GND.n2421 42.2793
R5399 GND.n5755 GND.n305 42.2793
R5400 GND.n5777 GND.n5776 42.2793
R5401 GND.n4241 GND.n4220 42.2793
R5402 GND.n2379 GND.n2378 42.2793
R5403 GND.n3837 GND.n3836 42.2793
R5404 GND.n3232 GND.n3231 42.2793
R5405 GND.n1026 GND.n1025 42.2793
R5406 GND.n1071 GND.n1017 42.2793
R5407 GND.n4787 GND.n4786 42.2793
R5408 GND.n3327 GND.n3326 41.6274
R5409 GND.n3037 GND.n3036 41.6274
R5410 GND.n1409 GND.n1253 40.577
R5411 GND.n1413 GND.n1253 40.577
R5412 GND.n1376 GND.n1264 40.577
R5413 GND.n1380 GND.n1264 40.577
R5414 GND.n1343 GND.n1275 40.577
R5415 GND.n1347 GND.n1275 40.577
R5416 GND.n1310 GND.n1286 40.577
R5417 GND.n1314 GND.n1286 40.577
R5418 GND.n69 GND.n57 40.4047
R5419 GND.n45 GND.n33 40.4047
R5420 GND.n22 GND.n10 40.4047
R5421 GND.n141 GND.n129 40.4047
R5422 GND.n117 GND.n105 40.4047
R5423 GND.n94 GND.n82 40.4047
R5424 GND.n3330 GND.n3329 37.9763
R5425 GND.n3040 GND.n3039 37.9763
R5426 GND.n4687 GND.n1187 36.9518
R5427 GND.n4413 GND.n2409 36.9518
R5428 GND.n1403 GND.n1402 36.702
R5429 GND.n1420 GND.n1419 36.702
R5430 GND.n1370 GND.n1369 36.702
R5431 GND.n1387 GND.n1386 36.702
R5432 GND.n1337 GND.n1336 36.702
R5433 GND.n1354 GND.n1353 36.702
R5434 GND.n1304 GND.n1303 36.702
R5435 GND.n1321 GND.n1320 36.702
R5436 GND.n3896 GND.n3895 36.059
R5437 GND.n3453 GND.n3288 36.059
R5438 GND.n69 GND.n68 35.8702
R5439 GND.n45 GND.n44 35.8702
R5440 GND.n22 GND.n21 35.8702
R5441 GND.n141 GND.n140 35.8702
R5442 GND.n117 GND.n116 35.8702
R5443 GND.n94 GND.n93 35.8702
R5444 GND.n4858 GND.n4857 34.5103
R5445 GND.n4857 GND.n4856 34.5103
R5446 GND.n4856 GND.n911 34.5103
R5447 GND.n4850 GND.n911 34.5103
R5448 GND.n4850 GND.n4849 34.5103
R5449 GND.n4849 GND.n4848 34.5103
R5450 GND.n4848 GND.n918 34.5103
R5451 GND.n4842 GND.n918 34.5103
R5452 GND.n4842 GND.n4841 34.5103
R5453 GND.n4841 GND.n4840 34.5103
R5454 GND.n4840 GND.n926 34.5103
R5455 GND.n4834 GND.n926 34.5103
R5456 GND.n4834 GND.n4833 34.5103
R5457 GND.n4833 GND.n4832 34.5103
R5458 GND.n4832 GND.n934 34.5103
R5459 GND.n4826 GND.n934 34.5103
R5460 GND.n4826 GND.n4825 34.5103
R5461 GND.n4825 GND.n4824 34.5103
R5462 GND.n4824 GND.n942 34.5103
R5463 GND.n4818 GND.n942 34.5103
R5464 GND.n4818 GND.n4817 34.5103
R5465 GND.n4817 GND.n4816 34.5103
R5466 GND.n4816 GND.n950 34.5103
R5467 GND.n4810 GND.n950 34.5103
R5468 GND.n4810 GND.n4809 34.5103
R5469 GND.n4809 GND.n4808 34.5103
R5470 GND.n4808 GND.n958 34.5103
R5471 GND.n4802 GND.n958 34.5103
R5472 GND.n4802 GND.n4801 34.5103
R5473 GND.n994 GND.n980 34.5103
R5474 GND.n1478 GND.n1172 34.5103
R5475 GND.n4637 GND.n1484 34.5103
R5476 GND.n4631 GND.n1484 34.5103
R5477 GND.n4631 GND.n4630 34.5103
R5478 GND.n4630 GND.n4629 34.5103
R5479 GND.n4017 GND.n4015 34.5103
R5480 GND.n4017 GND.n4016 34.5103
R5481 GND.n4016 GND.n2382 34.5103
R5482 GND.n2426 GND.n2395 34.5103
R5483 GND.n5747 GND.n272 34.5103
R5484 GND.n5740 GND.n278 34.5103
R5485 GND.n5740 GND.n5739 34.5103
R5486 GND.n5739 GND.n5738 34.5103
R5487 GND.n5738 GND.n318 34.5103
R5488 GND.n5732 GND.n318 34.5103
R5489 GND.n5732 GND.n5731 34.5103
R5490 GND.n5731 GND.n5730 34.5103
R5491 GND.n5730 GND.n328 34.5103
R5492 GND.n5724 GND.n328 34.5103
R5493 GND.n5724 GND.n5723 34.5103
R5494 GND.n5723 GND.n5722 34.5103
R5495 GND.n5722 GND.n336 34.5103
R5496 GND.n5716 GND.n336 34.5103
R5497 GND.n5716 GND.n5715 34.5103
R5498 GND.n5715 GND.n5714 34.5103
R5499 GND.n5714 GND.n344 34.5103
R5500 GND.n5708 GND.n344 34.5103
R5501 GND.n5708 GND.n5707 34.5103
R5502 GND.n5707 GND.n5706 34.5103
R5503 GND.n5706 GND.n352 34.5103
R5504 GND.n5700 GND.n352 34.5103
R5505 GND.n5700 GND.n5699 34.5103
R5506 GND.n5699 GND.n5698 34.5103
R5507 GND.n5698 GND.n360 34.5103
R5508 GND.n5692 GND.n360 34.5103
R5509 GND.n5692 GND.n5691 34.5103
R5510 GND.n5691 GND.n5690 34.5103
R5511 GND.n5690 GND.n368 34.5103
R5512 GND.n5684 GND.n368 34.5103
R5513 GND.n2768 GND.n2748 32.6207
R5514 GND.n2757 GND.n2756 32.6207
R5515 GND.n2733 GND.n2713 32.6207
R5516 GND.n2722 GND.n2721 32.6207
R5517 GND.n2698 GND.n2678 32.6207
R5518 GND.n2687 GND.n2686 32.6207
R5519 GND.n2664 GND.n2644 32.6207
R5520 GND.n2653 GND.n2652 32.6207
R5521 GND.n2618 GND.n2617 32.6207
R5522 GND.n2629 GND.n2609 32.6207
R5523 GND.n2583 GND.n2582 32.6207
R5524 GND.n2594 GND.n2574 32.6207
R5525 GND.n2548 GND.n2547 32.6207
R5526 GND.n2559 GND.n2539 32.6207
R5527 GND.n2514 GND.n2513 32.6207
R5528 GND.n2525 GND.n2505 32.6207
R5529 GND.n4015 GND.t70 32.4397
R5530 GND.n4687 GND.n1190 30.6565
R5531 GND.n4413 GND.n2405 30.6565
R5532 GND.n3278 GND.n2053 29.3338
R5533 GND.n3881 GND.n3021 29.3338
R5534 GND.n1398 GND.n1397 24.5923
R5535 GND.n1398 GND.n1257 24.5923
R5536 GND.n1404 GND.n1403 24.5923
R5537 GND.n1408 GND.n1407 24.5923
R5538 GND.n1409 GND.n1408 24.5923
R5539 GND.n1414 GND.n1413 24.5923
R5540 GND.n1415 GND.n1414 24.5923
R5541 GND.n1419 GND.n1418 24.5923
R5542 GND.n1424 GND.n1249 24.5923
R5543 GND.n1425 GND.n1424 24.5923
R5544 GND.n1365 GND.n1364 24.5923
R5545 GND.n1365 GND.n1268 24.5923
R5546 GND.n1371 GND.n1370 24.5923
R5547 GND.n1375 GND.n1374 24.5923
R5548 GND.n1376 GND.n1375 24.5923
R5549 GND.n1381 GND.n1380 24.5923
R5550 GND.n1382 GND.n1381 24.5923
R5551 GND.n1386 GND.n1385 24.5923
R5552 GND.n1391 GND.n1260 24.5923
R5553 GND.n1392 GND.n1391 24.5923
R5554 GND.n1332 GND.n1331 24.5923
R5555 GND.n1332 GND.n1279 24.5923
R5556 GND.n1338 GND.n1337 24.5923
R5557 GND.n1342 GND.n1341 24.5923
R5558 GND.n1343 GND.n1342 24.5923
R5559 GND.n1348 GND.n1347 24.5923
R5560 GND.n1349 GND.n1348 24.5923
R5561 GND.n1353 GND.n1352 24.5923
R5562 GND.n1358 GND.n1271 24.5923
R5563 GND.n1359 GND.n1358 24.5923
R5564 GND.n1299 GND.n1298 24.5923
R5565 GND.n1299 GND.n1290 24.5923
R5566 GND.n1305 GND.n1304 24.5923
R5567 GND.n1309 GND.n1308 24.5923
R5568 GND.n1310 GND.n1309 24.5923
R5569 GND.n1315 GND.n1314 24.5923
R5570 GND.n1316 GND.n1315 24.5923
R5571 GND.n1320 GND.n1319 24.5923
R5572 GND.n1325 GND.n1282 24.5923
R5573 GND.n1326 GND.n1325 24.5923
R5574 GND.n2776 GND.n2775 24.3439
R5575 GND.n2771 GND.n2746 24.3439
R5576 GND.n2769 GND.n2768 24.3439
R5577 GND.n2764 GND.n2763 24.3439
R5578 GND.n2761 GND.n2750 24.3439
R5579 GND.n2756 GND.n2755 24.3439
R5580 GND.n2741 GND.n2740 24.3439
R5581 GND.n2736 GND.n2711 24.3439
R5582 GND.n2734 GND.n2733 24.3439
R5583 GND.n2729 GND.n2728 24.3439
R5584 GND.n2726 GND.n2715 24.3439
R5585 GND.n2721 GND.n2720 24.3439
R5586 GND.n2706 GND.n2705 24.3439
R5587 GND.n2701 GND.n2676 24.3439
R5588 GND.n2699 GND.n2698 24.3439
R5589 GND.n2694 GND.n2693 24.3439
R5590 GND.n2691 GND.n2680 24.3439
R5591 GND.n2686 GND.n2685 24.3439
R5592 GND.n2672 GND.n2671 24.3439
R5593 GND.n2667 GND.n2642 24.3439
R5594 GND.n2665 GND.n2664 24.3439
R5595 GND.n2660 GND.n2659 24.3439
R5596 GND.n2657 GND.n2646 24.3439
R5597 GND.n2652 GND.n2651 24.3439
R5598 GND.n2617 GND.n2616 24.3439
R5599 GND.n2622 GND.n2611 24.3439
R5600 GND.n2625 GND.n2624 24.3439
R5601 GND.n2630 GND.n2629 24.3439
R5602 GND.n2632 GND.n2607 24.3439
R5603 GND.n2637 GND.n2636 24.3439
R5604 GND.n2582 GND.n2581 24.3439
R5605 GND.n2587 GND.n2576 24.3439
R5606 GND.n2590 GND.n2589 24.3439
R5607 GND.n2595 GND.n2594 24.3439
R5608 GND.n2597 GND.n2572 24.3439
R5609 GND.n2602 GND.n2601 24.3439
R5610 GND.n2547 GND.n2546 24.3439
R5611 GND.n2552 GND.n2541 24.3439
R5612 GND.n2555 GND.n2554 24.3439
R5613 GND.n2560 GND.n2559 24.3439
R5614 GND.n2562 GND.n2537 24.3439
R5615 GND.n2567 GND.n2566 24.3439
R5616 GND.n2513 GND.n2512 24.3439
R5617 GND.n2518 GND.n2507 24.3439
R5618 GND.n2521 GND.n2520 24.3439
R5619 GND.n2526 GND.n2525 24.3439
R5620 GND.n2528 GND.n2503 24.3439
R5621 GND.n2533 GND.n2532 24.3439
R5622 GND.n4651 GND.n4637 24.1574
R5623 GND.n4425 GND.n2382 24.1574
R5624 GND.n1431 GND.n1430 23.886
R5625 GND.n1404 GND.n1255 23.6087
R5626 GND.n1418 GND.n1251 23.6087
R5627 GND.n1371 GND.n1266 23.6087
R5628 GND.n1385 GND.n1262 23.6087
R5629 GND.n1338 GND.n1277 23.6087
R5630 GND.n1352 GND.n1273 23.6087
R5631 GND.n1305 GND.n1288 23.6087
R5632 GND.n1319 GND.n1284 23.6087
R5633 GND.n3333 GND.n2066 21.3859
R5634 GND.n4003 GND.n4002 21.3859
R5635 GND.n2777 GND.n2776 20.9359
R5636 GND.n2742 GND.n2741 20.9359
R5637 GND.n2707 GND.n2706 20.9359
R5638 GND.n2673 GND.n2672 20.9359
R5639 GND.n2638 GND.n2637 20.9359
R5640 GND.n2603 GND.n2602 20.9359
R5641 GND.n2568 GND.n2567 20.9359
R5642 GND.n2534 GND.n2533 20.9359
R5643 GND.n4779 GND.n996 20.7064
R5644 GND.n1078 GND.n1004 20.7064
R5645 GND.n4773 GND.n1007 20.7064
R5646 GND.n1772 GND.n1757 20.7064
R5647 GND.n1771 GND.n1734 20.7064
R5648 GND.n1819 GND.n1722 20.7064
R5649 GND.n1832 GND.n1723 20.7064
R5650 GND.n1727 GND.n1714 20.7064
R5651 GND.n1841 GND.n1710 20.7064
R5652 GND.n1847 GND.n1712 20.7064
R5653 GND.n1844 GND.n1699 20.7064
R5654 GND.n1857 GND.n1700 20.7064
R5655 GND.n1704 GND.n1692 20.7064
R5656 GND.n1866 GND.n1688 20.7064
R5657 GND.n1872 GND.n1690 20.7064
R5658 GND.n1868 GND.n1678 20.7064
R5659 GND.n1880 GND.n1681 20.7064
R5660 GND.n1943 GND.n1583 20.7064
R5661 GND.n1939 GND.n1938 20.7064
R5662 GND.n1594 GND.n1588 20.7064
R5663 GND.n1931 GND.n1595 20.7064
R5664 GND.n1930 GND.n1597 20.7064
R5665 GND.n1925 GND.n1606 20.7064
R5666 GND.n1922 GND.n1921 20.7064
R5667 GND.n1667 GND.n1610 20.7064
R5668 GND.n1914 GND.n1908 20.7064
R5669 GND.n1913 GND.n1909 20.7064
R5670 GND.n1953 GND.n1565 20.7064
R5671 GND.n1568 GND.n1557 20.7064
R5672 GND.n1962 GND.n1552 20.7064
R5673 GND.n1968 GND.n1554 20.7064
R5674 GND.n1965 GND.n1542 20.7064
R5675 GND.n1978 GND.n1543 20.7064
R5676 GND.n1546 GND.n1535 20.7064
R5677 GND.n1987 GND.n1529 20.7064
R5678 GND.n1992 GND.n1532 20.7064
R5679 GND.n1989 GND.n1518 20.7064
R5680 GND.n2002 GND.n1519 20.7064
R5681 GND.n1523 GND.n1510 20.7064
R5682 GND.n2026 GND.n1508 20.7064
R5683 GND.n2008 GND.n1497 20.7064
R5684 GND.n2036 GND.n1499 20.7064
R5685 GND.n2041 GND.n1493 20.7064
R5686 GND.n2040 GND.n1170 20.7064
R5687 GND.n4700 GND.n1172 20.7064
R5688 GND.n4389 GND.n2426 20.7064
R5689 GND.n2994 GND.n2427 20.7064
R5690 GND.n4381 GND.n2809 20.7064
R5691 GND.n2999 GND.n2811 20.7064
R5692 GND.n4375 GND.n2824 20.7064
R5693 GND.n4078 GND.n2827 20.7064
R5694 GND.n4085 GND.n2839 20.7064
R5695 GND.n4363 GND.n2847 20.7064
R5696 GND.n4093 GND.n2850 20.7064
R5697 GND.n4357 GND.n2857 20.7064
R5698 GND.n4100 GND.n2860 20.7064
R5699 GND.n4351 GND.n2868 20.7064
R5700 GND.n4108 GND.n2871 20.7064
R5701 GND.n4345 GND.n2878 20.7064
R5702 GND.n4115 GND.n2881 20.7064
R5703 GND.n4339 GND.n2890 20.7064
R5704 GND.n4135 GND.n2893 20.7064
R5705 GND.n4333 GND.n2900 20.7064
R5706 GND.n4328 GND.n2905 20.7064
R5707 GND.n4327 GND.n2908 20.7064
R5708 GND.n2915 GND.n2914 20.7064
R5709 GND.n4320 GND.n4319 20.7064
R5710 GND.n4149 GND.n2918 20.7064
R5711 GND.n5859 GND.n149 20.7064
R5712 GND.n4309 GND.n151 20.7064
R5713 GND.n4308 GND.n2931 20.7064
R5714 GND.n4165 GND.n4158 20.7064
R5715 GND.n5852 GND.n168 20.7064
R5716 GND.n5846 GND.n180 20.7064
R5717 GND.n4179 GND.n183 20.7064
R5718 GND.n5840 GND.n190 20.7064
R5719 GND.n4185 GND.n193 20.7064
R5720 GND.n5834 GND.n200 20.7064
R5721 GND.n4193 GND.n203 20.7064
R5722 GND.n5828 GND.n211 20.7064
R5723 GND.n4199 GND.n214 20.7064
R5724 GND.n5822 GND.n221 20.7064
R5725 GND.n4208 GND.n224 20.7064
R5726 GND.n5816 GND.n232 20.7064
R5727 GND.n4262 GND.n235 20.7064
R5728 GND.n4256 GND.n244 20.7064
R5729 GND.n5804 GND.n252 20.7064
R5730 GND.n4250 GND.n255 20.7064
R5731 GND.n5798 GND.n262 20.7064
R5732 GND.n5748 GND.n265 20.7064
R5733 GND.n2785 GND.n2784 20.1619
R5734 GND.n2771 GND.n2770 19.9621
R5735 GND.n2736 GND.n2735 19.9621
R5736 GND.n2701 GND.n2700 19.9621
R5737 GND.n2667 GND.n2666 19.9621
R5738 GND.n2632 GND.n2631 19.9621
R5739 GND.n2597 GND.n2596 19.9621
R5740 GND.n2562 GND.n2561 19.9621
R5741 GND.n2528 GND.n2527 19.9621
R5742 GND.n3325 GND.t49 19.8005
R5743 GND.n3325 GND.t88 19.8005
R5744 GND.n3035 GND.t101 19.8005
R5745 GND.n3035 GND.t71 19.8005
R5746 GND.n3324 GND.n3323 19.5087
R5747 GND.n4667 GND.n4666 19.3944
R5748 GND.n4666 GND.n4665 19.3944
R5749 GND.n4665 GND.n1209 19.3944
R5750 GND.n4660 GND.n1209 19.3944
R5751 GND.n4660 GND.n4659 19.3944
R5752 GND.n4659 GND.n4658 19.3944
R5753 GND.n1075 GND.n1010 19.3944
R5754 GND.n4771 GND.n1010 19.3944
R5755 GND.n4771 GND.n1011 19.3944
R5756 GND.n1084 GND.n1011 19.3944
R5757 GND.n1085 GND.n1084 19.3944
R5758 GND.n1086 GND.n1085 19.3944
R5759 GND.n1724 GND.n1086 19.3944
R5760 GND.n1724 GND.n1092 19.3944
R5761 GND.n1093 GND.n1092 19.3944
R5762 GND.n1094 GND.n1093 19.3944
R5763 GND.n1843 GND.n1094 19.3944
R5764 GND.n1843 GND.n1100 19.3944
R5765 GND.n1101 GND.n1100 19.3944
R5766 GND.n1102 GND.n1101 19.3944
R5767 GND.n1870 GND.n1102 19.3944
R5768 GND.n1870 GND.n1108 19.3944
R5769 GND.n1109 GND.n1108 19.3944
R5770 GND.n1110 GND.n1109 19.3944
R5771 GND.n1941 GND.n1110 19.3944
R5772 GND.n1941 GND.n1116 19.3944
R5773 GND.n1117 GND.n1116 19.3944
R5774 GND.n1118 GND.n1117 19.3944
R5775 GND.n1599 GND.n1118 19.3944
R5776 GND.n1599 GND.n1124 19.3944
R5777 GND.n1125 GND.n1124 19.3944
R5778 GND.n1126 GND.n1125 19.3944
R5779 GND.n1910 GND.n1126 19.3944
R5780 GND.n1910 GND.n1132 19.3944
R5781 GND.n1133 GND.n1132 19.3944
R5782 GND.n1134 GND.n1133 19.3944
R5783 GND.n1556 GND.n1134 19.3944
R5784 GND.n1556 GND.n1140 19.3944
R5785 GND.n1141 GND.n1140 19.3944
R5786 GND.n1142 GND.n1141 19.3944
R5787 GND.n1533 GND.n1142 19.3944
R5788 GND.n1533 GND.n1148 19.3944
R5789 GND.n1149 GND.n1148 19.3944
R5790 GND.n1150 GND.n1149 19.3944
R5791 GND.n1520 GND.n1150 19.3944
R5792 GND.n1520 GND.n1156 19.3944
R5793 GND.n1157 GND.n1156 19.3944
R5794 GND.n1158 GND.n1157 19.3944
R5795 GND.n1495 GND.n1158 19.3944
R5796 GND.n1495 GND.n1164 19.3944
R5797 GND.n1165 GND.n1164 19.3944
R5798 GND.n1166 GND.n1165 19.3944
R5799 GND.n1173 GND.n1166 19.3944
R5800 GND.n1080 GND.n1077 19.3944
R5801 GND.n4769 GND.n1080 19.3944
R5802 GND.n4769 GND.n4768 19.3944
R5803 GND.n4768 GND.n4767 19.3944
R5804 GND.n4767 GND.n1083 19.3944
R5805 GND.n4763 GND.n1083 19.3944
R5806 GND.n4763 GND.n4762 19.3944
R5807 GND.n4762 GND.n4761 19.3944
R5808 GND.n4761 GND.n1091 19.3944
R5809 GND.n4757 GND.n1091 19.3944
R5810 GND.n4757 GND.n4756 19.3944
R5811 GND.n4756 GND.n4755 19.3944
R5812 GND.n4755 GND.n1099 19.3944
R5813 GND.n4751 GND.n1099 19.3944
R5814 GND.n4751 GND.n4750 19.3944
R5815 GND.n4750 GND.n4749 19.3944
R5816 GND.n4749 GND.n1107 19.3944
R5817 GND.n4745 GND.n1107 19.3944
R5818 GND.n4745 GND.n4744 19.3944
R5819 GND.n4744 GND.n4743 19.3944
R5820 GND.n4743 GND.n1115 19.3944
R5821 GND.n4739 GND.n1115 19.3944
R5822 GND.n4739 GND.n4738 19.3944
R5823 GND.n4738 GND.n4737 19.3944
R5824 GND.n4737 GND.n1123 19.3944
R5825 GND.n4733 GND.n1123 19.3944
R5826 GND.n4733 GND.n4732 19.3944
R5827 GND.n4732 GND.n4731 19.3944
R5828 GND.n4731 GND.n1131 19.3944
R5829 GND.n4727 GND.n1131 19.3944
R5830 GND.n4727 GND.n4726 19.3944
R5831 GND.n4726 GND.n4725 19.3944
R5832 GND.n4725 GND.n1139 19.3944
R5833 GND.n4721 GND.n1139 19.3944
R5834 GND.n4721 GND.n4720 19.3944
R5835 GND.n4720 GND.n4719 19.3944
R5836 GND.n4719 GND.n1147 19.3944
R5837 GND.n4715 GND.n1147 19.3944
R5838 GND.n4715 GND.n4714 19.3944
R5839 GND.n4714 GND.n4713 19.3944
R5840 GND.n4713 GND.n1155 19.3944
R5841 GND.n4709 GND.n1155 19.3944
R5842 GND.n4709 GND.n4708 19.3944
R5843 GND.n4708 GND.n4707 19.3944
R5844 GND.n4707 GND.n1163 19.3944
R5845 GND.n4703 GND.n1163 19.3944
R5846 GND.n4703 GND.n4702 19.3944
R5847 GND.n4695 GND.n4694 19.3944
R5848 GND.n4694 GND.n4693 19.3944
R5849 GND.n4693 GND.n1182 19.3944
R5850 GND.n4689 GND.n1182 19.3944
R5851 GND.n4689 GND.n4688 19.3944
R5852 GND.n4686 GND.n1192 19.3944
R5853 GND.n4682 GND.n1192 19.3944
R5854 GND.n4682 GND.n4681 19.3944
R5855 GND.n4681 GND.n4680 19.3944
R5856 GND.n4680 GND.n1197 19.3944
R5857 GND.n4676 GND.n1197 19.3944
R5858 GND.n4676 GND.n4675 19.3944
R5859 GND.n4675 GND.n4674 19.3944
R5860 GND.n5548 GND.n455 19.3944
R5861 GND.n5548 GND.n451 19.3944
R5862 GND.n5554 GND.n451 19.3944
R5863 GND.n5554 GND.n449 19.3944
R5864 GND.n5558 GND.n449 19.3944
R5865 GND.n5558 GND.n445 19.3944
R5866 GND.n5564 GND.n445 19.3944
R5867 GND.n5564 GND.n443 19.3944
R5868 GND.n5568 GND.n443 19.3944
R5869 GND.n5568 GND.n439 19.3944
R5870 GND.n5574 GND.n439 19.3944
R5871 GND.n5574 GND.n437 19.3944
R5872 GND.n5578 GND.n437 19.3944
R5873 GND.n5578 GND.n433 19.3944
R5874 GND.n5584 GND.n433 19.3944
R5875 GND.n5584 GND.n431 19.3944
R5876 GND.n5588 GND.n431 19.3944
R5877 GND.n5588 GND.n427 19.3944
R5878 GND.n5594 GND.n427 19.3944
R5879 GND.n5594 GND.n425 19.3944
R5880 GND.n5598 GND.n425 19.3944
R5881 GND.n5598 GND.n421 19.3944
R5882 GND.n5604 GND.n421 19.3944
R5883 GND.n5604 GND.n419 19.3944
R5884 GND.n5608 GND.n419 19.3944
R5885 GND.n5608 GND.n415 19.3944
R5886 GND.n5614 GND.n415 19.3944
R5887 GND.n5614 GND.n413 19.3944
R5888 GND.n5618 GND.n413 19.3944
R5889 GND.n5618 GND.n409 19.3944
R5890 GND.n5624 GND.n409 19.3944
R5891 GND.n5624 GND.n407 19.3944
R5892 GND.n5628 GND.n407 19.3944
R5893 GND.n5628 GND.n403 19.3944
R5894 GND.n5634 GND.n403 19.3944
R5895 GND.n5634 GND.n401 19.3944
R5896 GND.n5638 GND.n401 19.3944
R5897 GND.n5638 GND.n397 19.3944
R5898 GND.n5644 GND.n397 19.3944
R5899 GND.n5644 GND.n395 19.3944
R5900 GND.n5648 GND.n395 19.3944
R5901 GND.n5648 GND.n391 19.3944
R5902 GND.n5654 GND.n391 19.3944
R5903 GND.n5654 GND.n389 19.3944
R5904 GND.n5658 GND.n389 19.3944
R5905 GND.n5658 GND.n385 19.3944
R5906 GND.n5664 GND.n385 19.3944
R5907 GND.n5664 GND.n383 19.3944
R5908 GND.n5668 GND.n383 19.3944
R5909 GND.n5668 GND.n379 19.3944
R5910 GND.n5674 GND.n379 19.3944
R5911 GND.n5674 GND.n377 19.3944
R5912 GND.n5680 GND.n377 19.3944
R5913 GND.n5680 GND.n5679 19.3944
R5914 GND.n4974 GND.n797 19.3944
R5915 GND.n4978 GND.n797 19.3944
R5916 GND.n4978 GND.n793 19.3944
R5917 GND.n4984 GND.n793 19.3944
R5918 GND.n4984 GND.n791 19.3944
R5919 GND.n4988 GND.n791 19.3944
R5920 GND.n4988 GND.n787 19.3944
R5921 GND.n4994 GND.n787 19.3944
R5922 GND.n4994 GND.n785 19.3944
R5923 GND.n4998 GND.n785 19.3944
R5924 GND.n4998 GND.n781 19.3944
R5925 GND.n5004 GND.n781 19.3944
R5926 GND.n5004 GND.n779 19.3944
R5927 GND.n5008 GND.n779 19.3944
R5928 GND.n5008 GND.n775 19.3944
R5929 GND.n5014 GND.n775 19.3944
R5930 GND.n5014 GND.n773 19.3944
R5931 GND.n5018 GND.n773 19.3944
R5932 GND.n5018 GND.n769 19.3944
R5933 GND.n5024 GND.n769 19.3944
R5934 GND.n5024 GND.n767 19.3944
R5935 GND.n5028 GND.n767 19.3944
R5936 GND.n5028 GND.n763 19.3944
R5937 GND.n5034 GND.n763 19.3944
R5938 GND.n5034 GND.n761 19.3944
R5939 GND.n5038 GND.n761 19.3944
R5940 GND.n5038 GND.n757 19.3944
R5941 GND.n5044 GND.n757 19.3944
R5942 GND.n5044 GND.n755 19.3944
R5943 GND.n5048 GND.n755 19.3944
R5944 GND.n5048 GND.n751 19.3944
R5945 GND.n5054 GND.n751 19.3944
R5946 GND.n5054 GND.n749 19.3944
R5947 GND.n5058 GND.n749 19.3944
R5948 GND.n5058 GND.n745 19.3944
R5949 GND.n5064 GND.n745 19.3944
R5950 GND.n5064 GND.n743 19.3944
R5951 GND.n5068 GND.n743 19.3944
R5952 GND.n5068 GND.n739 19.3944
R5953 GND.n5074 GND.n739 19.3944
R5954 GND.n5074 GND.n737 19.3944
R5955 GND.n5078 GND.n737 19.3944
R5956 GND.n5078 GND.n733 19.3944
R5957 GND.n5084 GND.n733 19.3944
R5958 GND.n5084 GND.n731 19.3944
R5959 GND.n5088 GND.n731 19.3944
R5960 GND.n5088 GND.n727 19.3944
R5961 GND.n5094 GND.n727 19.3944
R5962 GND.n5094 GND.n725 19.3944
R5963 GND.n5098 GND.n725 19.3944
R5964 GND.n5098 GND.n721 19.3944
R5965 GND.n5104 GND.n721 19.3944
R5966 GND.n5104 GND.n719 19.3944
R5967 GND.n5108 GND.n719 19.3944
R5968 GND.n5108 GND.n715 19.3944
R5969 GND.n5114 GND.n715 19.3944
R5970 GND.n5114 GND.n713 19.3944
R5971 GND.n5118 GND.n713 19.3944
R5972 GND.n5118 GND.n709 19.3944
R5973 GND.n5124 GND.n709 19.3944
R5974 GND.n5124 GND.n707 19.3944
R5975 GND.n5128 GND.n707 19.3944
R5976 GND.n5128 GND.n703 19.3944
R5977 GND.n5134 GND.n703 19.3944
R5978 GND.n5134 GND.n701 19.3944
R5979 GND.n5138 GND.n701 19.3944
R5980 GND.n5138 GND.n697 19.3944
R5981 GND.n5144 GND.n697 19.3944
R5982 GND.n5144 GND.n695 19.3944
R5983 GND.n5148 GND.n695 19.3944
R5984 GND.n5148 GND.n691 19.3944
R5985 GND.n5154 GND.n691 19.3944
R5986 GND.n5154 GND.n689 19.3944
R5987 GND.n5158 GND.n689 19.3944
R5988 GND.n5158 GND.n685 19.3944
R5989 GND.n5164 GND.n685 19.3944
R5990 GND.n5164 GND.n683 19.3944
R5991 GND.n5168 GND.n683 19.3944
R5992 GND.n5168 GND.n679 19.3944
R5993 GND.n5174 GND.n679 19.3944
R5994 GND.n5174 GND.n677 19.3944
R5995 GND.n5178 GND.n677 19.3944
R5996 GND.n5178 GND.n673 19.3944
R5997 GND.n5184 GND.n673 19.3944
R5998 GND.n5184 GND.n671 19.3944
R5999 GND.n5188 GND.n671 19.3944
R6000 GND.n5188 GND.n667 19.3944
R6001 GND.n5194 GND.n667 19.3944
R6002 GND.n5194 GND.n665 19.3944
R6003 GND.n5198 GND.n665 19.3944
R6004 GND.n5198 GND.n661 19.3944
R6005 GND.n5204 GND.n661 19.3944
R6006 GND.n5204 GND.n659 19.3944
R6007 GND.n5208 GND.n659 19.3944
R6008 GND.n5208 GND.n655 19.3944
R6009 GND.n5214 GND.n655 19.3944
R6010 GND.n5214 GND.n653 19.3944
R6011 GND.n5218 GND.n653 19.3944
R6012 GND.n5218 GND.n649 19.3944
R6013 GND.n5224 GND.n649 19.3944
R6014 GND.n5224 GND.n647 19.3944
R6015 GND.n5228 GND.n647 19.3944
R6016 GND.n5228 GND.n643 19.3944
R6017 GND.n5234 GND.n643 19.3944
R6018 GND.n5234 GND.n641 19.3944
R6019 GND.n5238 GND.n641 19.3944
R6020 GND.n5238 GND.n637 19.3944
R6021 GND.n5244 GND.n637 19.3944
R6022 GND.n5244 GND.n635 19.3944
R6023 GND.n5248 GND.n635 19.3944
R6024 GND.n5248 GND.n631 19.3944
R6025 GND.n5254 GND.n631 19.3944
R6026 GND.n5254 GND.n629 19.3944
R6027 GND.n5258 GND.n629 19.3944
R6028 GND.n5258 GND.n625 19.3944
R6029 GND.n5264 GND.n625 19.3944
R6030 GND.n5264 GND.n623 19.3944
R6031 GND.n5268 GND.n623 19.3944
R6032 GND.n5268 GND.n619 19.3944
R6033 GND.n5274 GND.n619 19.3944
R6034 GND.n5274 GND.n617 19.3944
R6035 GND.n5278 GND.n617 19.3944
R6036 GND.n5278 GND.n613 19.3944
R6037 GND.n5284 GND.n613 19.3944
R6038 GND.n5284 GND.n611 19.3944
R6039 GND.n5288 GND.n611 19.3944
R6040 GND.n5288 GND.n607 19.3944
R6041 GND.n5294 GND.n607 19.3944
R6042 GND.n5294 GND.n605 19.3944
R6043 GND.n5298 GND.n605 19.3944
R6044 GND.n5298 GND.n601 19.3944
R6045 GND.n5304 GND.n601 19.3944
R6046 GND.n5304 GND.n599 19.3944
R6047 GND.n5308 GND.n599 19.3944
R6048 GND.n5308 GND.n595 19.3944
R6049 GND.n5314 GND.n595 19.3944
R6050 GND.n5314 GND.n593 19.3944
R6051 GND.n5318 GND.n593 19.3944
R6052 GND.n5318 GND.n589 19.3944
R6053 GND.n5324 GND.n589 19.3944
R6054 GND.n5324 GND.n587 19.3944
R6055 GND.n5328 GND.n587 19.3944
R6056 GND.n5328 GND.n583 19.3944
R6057 GND.n5334 GND.n583 19.3944
R6058 GND.n5334 GND.n581 19.3944
R6059 GND.n5338 GND.n581 19.3944
R6060 GND.n5338 GND.n577 19.3944
R6061 GND.n5344 GND.n577 19.3944
R6062 GND.n5344 GND.n575 19.3944
R6063 GND.n5348 GND.n575 19.3944
R6064 GND.n5348 GND.n571 19.3944
R6065 GND.n5354 GND.n571 19.3944
R6066 GND.n5354 GND.n569 19.3944
R6067 GND.n5358 GND.n569 19.3944
R6068 GND.n5358 GND.n565 19.3944
R6069 GND.n5364 GND.n565 19.3944
R6070 GND.n5364 GND.n563 19.3944
R6071 GND.n5368 GND.n563 19.3944
R6072 GND.n5368 GND.n559 19.3944
R6073 GND.n5374 GND.n559 19.3944
R6074 GND.n5374 GND.n557 19.3944
R6075 GND.n5378 GND.n557 19.3944
R6076 GND.n5378 GND.n553 19.3944
R6077 GND.n5384 GND.n553 19.3944
R6078 GND.n5384 GND.n551 19.3944
R6079 GND.n5388 GND.n551 19.3944
R6080 GND.n5388 GND.n547 19.3944
R6081 GND.n5394 GND.n547 19.3944
R6082 GND.n5394 GND.n545 19.3944
R6083 GND.n5398 GND.n545 19.3944
R6084 GND.n5398 GND.n541 19.3944
R6085 GND.n5404 GND.n541 19.3944
R6086 GND.n5404 GND.n539 19.3944
R6087 GND.n5408 GND.n539 19.3944
R6088 GND.n5408 GND.n535 19.3944
R6089 GND.n5414 GND.n535 19.3944
R6090 GND.n5414 GND.n533 19.3944
R6091 GND.n5418 GND.n533 19.3944
R6092 GND.n5418 GND.n529 19.3944
R6093 GND.n5424 GND.n529 19.3944
R6094 GND.n5424 GND.n527 19.3944
R6095 GND.n5428 GND.n527 19.3944
R6096 GND.n5428 GND.n523 19.3944
R6097 GND.n5434 GND.n523 19.3944
R6098 GND.n5434 GND.n521 19.3944
R6099 GND.n5438 GND.n521 19.3944
R6100 GND.n5438 GND.n517 19.3944
R6101 GND.n5444 GND.n517 19.3944
R6102 GND.n5444 GND.n515 19.3944
R6103 GND.n5448 GND.n515 19.3944
R6104 GND.n5448 GND.n511 19.3944
R6105 GND.n5454 GND.n511 19.3944
R6106 GND.n5454 GND.n509 19.3944
R6107 GND.n5458 GND.n509 19.3944
R6108 GND.n5458 GND.n505 19.3944
R6109 GND.n5464 GND.n505 19.3944
R6110 GND.n5464 GND.n503 19.3944
R6111 GND.n5468 GND.n503 19.3944
R6112 GND.n5468 GND.n499 19.3944
R6113 GND.n5474 GND.n499 19.3944
R6114 GND.n5474 GND.n497 19.3944
R6115 GND.n5478 GND.n497 19.3944
R6116 GND.n5478 GND.n493 19.3944
R6117 GND.n5484 GND.n493 19.3944
R6118 GND.n5484 GND.n491 19.3944
R6119 GND.n5488 GND.n491 19.3944
R6120 GND.n5488 GND.n487 19.3944
R6121 GND.n5494 GND.n487 19.3944
R6122 GND.n5494 GND.n485 19.3944
R6123 GND.n5498 GND.n485 19.3944
R6124 GND.n5498 GND.n481 19.3944
R6125 GND.n5504 GND.n481 19.3944
R6126 GND.n5504 GND.n479 19.3944
R6127 GND.n5508 GND.n479 19.3944
R6128 GND.n5508 GND.n475 19.3944
R6129 GND.n5514 GND.n475 19.3944
R6130 GND.n5514 GND.n473 19.3944
R6131 GND.n5518 GND.n473 19.3944
R6132 GND.n5518 GND.n469 19.3944
R6133 GND.n5524 GND.n469 19.3944
R6134 GND.n5524 GND.n467 19.3944
R6135 GND.n5528 GND.n467 19.3944
R6136 GND.n5528 GND.n463 19.3944
R6137 GND.n5534 GND.n463 19.3944
R6138 GND.n5534 GND.n461 19.3944
R6139 GND.n5538 GND.n461 19.3944
R6140 GND.n5538 GND.n457 19.3944
R6141 GND.n5544 GND.n457 19.3944
R6142 GND.n4422 GND.n4421 19.3944
R6143 GND.n4421 GND.n4420 19.3944
R6144 GND.n4420 GND.n4419 19.3944
R6145 GND.n4419 GND.n4417 19.3944
R6146 GND.n4417 GND.n4414 19.3944
R6147 GND.n4412 GND.n4409 19.3944
R6148 GND.n4409 GND.n4408 19.3944
R6149 GND.n4408 GND.n4405 19.3944
R6150 GND.n4405 GND.n4404 19.3944
R6151 GND.n4404 GND.n4401 19.3944
R6152 GND.n4401 GND.n4400 19.3944
R6153 GND.n4400 GND.n4397 19.3944
R6154 GND.n4397 GND.n4396 19.3944
R6155 GND.n4384 GND.n2425 19.3944
R6156 GND.n4384 GND.n4383 19.3944
R6157 GND.n4383 GND.n2807 19.3944
R6158 GND.n2990 GND.n2807 19.3944
R6159 GND.n4080 GND.n2990 19.3944
R6160 GND.n4081 GND.n4080 19.3944
R6161 GND.n4083 GND.n4081 19.3944
R6162 GND.n4083 GND.n2986 19.3944
R6163 GND.n4095 GND.n2986 19.3944
R6164 GND.n4096 GND.n4095 19.3944
R6165 GND.n4098 GND.n4096 19.3944
R6166 GND.n4098 GND.n2982 19.3944
R6167 GND.n4110 GND.n2982 19.3944
R6168 GND.n4111 GND.n4110 19.3944
R6169 GND.n4113 GND.n4111 19.3944
R6170 GND.n4113 GND.n2978 19.3944
R6171 GND.n4137 GND.n2978 19.3944
R6172 GND.n4138 GND.n4137 19.3944
R6173 GND.n4139 GND.n4138 19.3944
R6174 GND.n4139 GND.n2977 19.3944
R6175 GND.n4147 GND.n2977 19.3944
R6176 GND.n4148 GND.n4147 19.3944
R6177 GND.n4151 GND.n4148 19.3944
R6178 GND.n4152 GND.n4151 19.3944
R6179 GND.n4153 GND.n4152 19.3944
R6180 GND.n4154 GND.n4153 19.3944
R6181 GND.n4167 GND.n4154 19.3944
R6182 GND.n4168 GND.n4167 19.3944
R6183 GND.n4169 GND.n4168 19.3944
R6184 GND.n4169 GND.n2972 19.3944
R6185 GND.n4181 GND.n2972 19.3944
R6186 GND.n4182 GND.n4181 19.3944
R6187 GND.n4183 GND.n4182 19.3944
R6188 GND.n4183 GND.n2967 19.3944
R6189 GND.n4195 GND.n2967 19.3944
R6190 GND.n4196 GND.n4195 19.3944
R6191 GND.n4197 GND.n4196 19.3944
R6192 GND.n4197 GND.n2962 19.3944
R6193 GND.n4210 GND.n2962 19.3944
R6194 GND.n4211 GND.n4210 19.3944
R6195 GND.n4212 GND.n4211 19.3944
R6196 GND.n4213 GND.n4212 19.3944
R6197 GND.n4254 GND.n4213 19.3944
R6198 GND.n4254 GND.n4253 19.3944
R6199 GND.n4253 GND.n4252 19.3944
R6200 GND.n4252 GND.n307 19.3944
R6201 GND.n5750 GND.n307 19.3944
R6202 GND.n4387 GND.n4386 19.3944
R6203 GND.n4386 GND.n2805 19.3944
R6204 GND.n2830 GND.n2805 19.3944
R6205 GND.n4373 GND.n2830 19.3944
R6206 GND.n4373 GND.n4372 19.3944
R6207 GND.n4372 GND.n4371 19.3944
R6208 GND.n4371 GND.n2835 19.3944
R6209 GND.n4361 GND.n2835 19.3944
R6210 GND.n4361 GND.n4360 19.3944
R6211 GND.n4360 GND.n4359 19.3944
R6212 GND.n4359 GND.n2855 19.3944
R6213 GND.n4349 GND.n2855 19.3944
R6214 GND.n4349 GND.n4348 19.3944
R6215 GND.n4348 GND.n4347 19.3944
R6216 GND.n4347 GND.n2876 19.3944
R6217 GND.n4337 GND.n2876 19.3944
R6218 GND.n4337 GND.n4336 19.3944
R6219 GND.n4336 GND.n4335 19.3944
R6220 GND.n4335 GND.n2898 19.3944
R6221 GND.n4142 GND.n2898 19.3944
R6222 GND.n4142 GND.n2921 19.3944
R6223 GND.n4314 GND.n2921 19.3944
R6224 GND.n4314 GND.n4313 19.3944
R6225 GND.n4313 GND.n4312 19.3944
R6226 GND.n4312 GND.n4311 19.3944
R6227 GND.n4311 GND.n2926 19.3944
R6228 GND.n2926 GND.n174 19.3944
R6229 GND.n5850 GND.n174 19.3944
R6230 GND.n5850 GND.n5849 19.3944
R6231 GND.n5849 GND.n5848 19.3944
R6232 GND.n5848 GND.n178 19.3944
R6233 GND.n5838 GND.n178 19.3944
R6234 GND.n5838 GND.n5837 19.3944
R6235 GND.n5837 GND.n5836 19.3944
R6236 GND.n5836 GND.n198 19.3944
R6237 GND.n5826 GND.n198 19.3944
R6238 GND.n5826 GND.n5825 19.3944
R6239 GND.n5825 GND.n5824 19.3944
R6240 GND.n5824 GND.n219 19.3944
R6241 GND.n5814 GND.n219 19.3944
R6242 GND.n5814 GND.n5813 19.3944
R6243 GND.n5813 GND.n5812 19.3944
R6244 GND.n5812 GND.n240 19.3944
R6245 GND.n5802 GND.n240 19.3944
R6246 GND.n5802 GND.n5801 19.3944
R6247 GND.n5801 GND.n5800 19.3944
R6248 GND.n5800 GND.n260 19.3944
R6249 GND.n5774 GND.n5771 19.3944
R6250 GND.n5771 GND.n5770 19.3944
R6251 GND.n5770 GND.n5767 19.3944
R6252 GND.n5767 GND.n5766 19.3944
R6253 GND.n5766 GND.n5763 19.3944
R6254 GND.n5763 GND.n5762 19.3944
R6255 GND.n5762 GND.n5759 19.3944
R6256 GND.n5759 GND.n5758 19.3944
R6257 GND.n5792 GND.n270 19.3944
R6258 GND.n5787 GND.n270 19.3944
R6259 GND.n5787 GND.n5786 19.3944
R6260 GND.n5786 GND.n5785 19.3944
R6261 GND.n5785 GND.n5782 19.3944
R6262 GND.n5782 GND.n5781 19.3944
R6263 GND.n5781 GND.n5778 19.3944
R6264 GND.n4226 GND.n4224 19.3944
R6265 GND.n4229 GND.n4226 19.3944
R6266 GND.n4232 GND.n4229 19.3944
R6267 GND.n4235 GND.n4232 19.3944
R6268 GND.n4235 GND.n4222 19.3944
R6269 GND.n4240 GND.n4222 19.3944
R6270 GND.n2997 GND.n2993 19.3944
R6271 GND.n2998 GND.n2997 19.3944
R6272 GND.n3001 GND.n2998 19.3944
R6273 GND.n3001 GND.n2991 19.3944
R6274 GND.n3005 GND.n2991 19.3944
R6275 GND.n3005 GND.n2989 19.3944
R6276 GND.n4087 GND.n2989 19.3944
R6277 GND.n4087 GND.n2987 19.3944
R6278 GND.n4091 GND.n2987 19.3944
R6279 GND.n4091 GND.n2985 19.3944
R6280 GND.n4102 GND.n2985 19.3944
R6281 GND.n4102 GND.n2983 19.3944
R6282 GND.n4106 GND.n2983 19.3944
R6283 GND.n4106 GND.n2981 19.3944
R6284 GND.n4117 GND.n2981 19.3944
R6285 GND.n4117 GND.n2979 19.3944
R6286 GND.n4133 GND.n2979 19.3944
R6287 GND.n4133 GND.n4132 19.3944
R6288 GND.n4132 GND.n4131 19.3944
R6289 GND.n4131 GND.n4130 19.3944
R6290 GND.n4130 GND.n4127 19.3944
R6291 GND.n4127 GND.n4126 19.3944
R6292 GND.n4126 GND.n145 19.3944
R6293 GND.n5861 GND.n145 19.3944
R6294 GND.n5861 GND.n146 19.3944
R6295 GND.n4160 GND.n146 19.3944
R6296 GND.n4163 GND.n4160 19.3944
R6297 GND.n4163 GND.n2976 19.3944
R6298 GND.n4173 GND.n2976 19.3944
R6299 GND.n4173 GND.n2974 19.3944
R6300 GND.n4177 GND.n2974 19.3944
R6301 GND.n4177 GND.n2971 19.3944
R6302 GND.n4187 GND.n2971 19.3944
R6303 GND.n4187 GND.n2969 19.3944
R6304 GND.n4191 GND.n2969 19.3944
R6305 GND.n4191 GND.n2966 19.3944
R6306 GND.n4201 GND.n2966 19.3944
R6307 GND.n4201 GND.n2964 19.3944
R6308 GND.n4206 GND.n2964 19.3944
R6309 GND.n4206 GND.n2957 19.3944
R6310 GND.n4260 GND.n2957 19.3944
R6311 GND.n4260 GND.n4259 19.3944
R6312 GND.n4259 GND.n4258 19.3944
R6313 GND.n4258 GND.n2961 19.3944
R6314 GND.n4248 GND.n2961 19.3944
R6315 GND.n4248 GND.n4247 19.3944
R6316 GND.n4247 GND.n4246 19.3944
R6317 GND.n2801 GND.n2800 19.3944
R6318 GND.n2800 GND.n2797 19.3944
R6319 GND.n2797 GND.n2796 19.3944
R6320 GND.n2796 GND.n2793 19.3944
R6321 GND.n2793 GND.n2792 19.3944
R6322 GND.n2792 GND.n2789 19.3944
R6323 GND.n3840 GND.n3806 19.3944
R6324 GND.n3884 GND.n3806 19.3944
R6325 GND.n3885 GND.n3884 19.3944
R6326 GND.n3879 GND.n3878 19.3944
R6327 GND.n3878 GND.n3819 19.3944
R6328 GND.n3874 GND.n3819 19.3944
R6329 GND.n3874 GND.n3871 19.3944
R6330 GND.n3871 GND.n3868 19.3944
R6331 GND.n3868 GND.n3867 19.3944
R6332 GND.n3867 GND.n3864 19.3944
R6333 GND.n3864 GND.n3863 19.3944
R6334 GND.n3863 GND.n3860 19.3944
R6335 GND.n3860 GND.n3859 19.3944
R6336 GND.n3859 GND.n3856 19.3944
R6337 GND.n3856 GND.n3855 19.3944
R6338 GND.n3855 GND.n3852 19.3944
R6339 GND.n3852 GND.n3851 19.3944
R6340 GND.n3851 GND.n3848 19.3944
R6341 GND.n3848 GND.n3847 19.3944
R6342 GND.n3847 GND.n3844 19.3944
R6343 GND.n3844 GND.n3843 19.3944
R6344 GND.n3282 GND.n3196 19.3944
R6345 GND.n3480 GND.n3196 19.3944
R6346 GND.n3481 GND.n3480 19.3944
R6347 GND.n3483 GND.n3481 19.3944
R6348 GND.n3483 GND.n3194 19.3944
R6349 GND.n3487 GND.n3194 19.3944
R6350 GND.n3487 GND.n3184 19.3944
R6351 GND.n3509 GND.n3184 19.3944
R6352 GND.n3509 GND.n3182 19.3944
R6353 GND.n3513 GND.n3182 19.3944
R6354 GND.n3513 GND.n3178 19.3944
R6355 GND.n3556 GND.n3178 19.3944
R6356 GND.n3556 GND.n3176 19.3944
R6357 GND.n3561 GND.n3176 19.3944
R6358 GND.n3561 GND.n3160 19.3944
R6359 GND.n3582 GND.n3160 19.3944
R6360 GND.n3582 GND.n3581 19.3944
R6361 GND.n3581 GND.n3580 19.3944
R6362 GND.n3580 GND.n3173 19.3944
R6363 GND.n3173 GND.n3172 19.3944
R6364 GND.n3172 GND.n3170 19.3944
R6365 GND.n3170 GND.n3169 19.3944
R6366 GND.n3169 GND.n3136 19.3944
R6367 GND.n3636 GND.n3136 19.3944
R6368 GND.n3636 GND.n3134 19.3944
R6369 GND.n3657 GND.n3134 19.3944
R6370 GND.n3657 GND.n3656 19.3944
R6371 GND.n3656 GND.n3655 19.3944
R6372 GND.n3655 GND.n3653 19.3944
R6373 GND.n3653 GND.n3652 19.3944
R6374 GND.n3652 GND.n3644 19.3944
R6375 GND.n3648 GND.n3644 19.3944
R6376 GND.n3648 GND.n3120 19.3944
R6377 GND.n3700 GND.n3120 19.3944
R6378 GND.n3701 GND.n3700 19.3944
R6379 GND.n3703 GND.n3701 19.3944
R6380 GND.n3703 GND.n3118 19.3944
R6381 GND.n3708 GND.n3118 19.3944
R6382 GND.n3708 GND.n3108 19.3944
R6383 GND.n3749 GND.n3108 19.3944
R6384 GND.n3750 GND.n3749 19.3944
R6385 GND.n3750 GND.n3106 19.3944
R6386 GND.n3754 GND.n3106 19.3944
R6387 GND.n3754 GND.n3104 19.3944
R6388 GND.n3758 GND.n3104 19.3944
R6389 GND.n3758 GND.n3102 19.3944
R6390 GND.n3766 GND.n3102 19.3944
R6391 GND.n3766 GND.n3765 19.3944
R6392 GND.n3765 GND.n3764 19.3944
R6393 GND.n3764 GND.n3094 19.3944
R6394 GND.n3802 GND.n3094 19.3944
R6395 GND.n3802 GND.n3092 19.3944
R6396 GND.n3888 GND.n3092 19.3944
R6397 GND.n3275 GND.n3274 19.3944
R6398 GND.n3274 GND.n3273 19.3944
R6399 GND.n3273 GND.n3272 19.3944
R6400 GND.n3272 GND.n3270 19.3944
R6401 GND.n3270 GND.n3267 19.3944
R6402 GND.n3267 GND.n3266 19.3944
R6403 GND.n3266 GND.n3263 19.3944
R6404 GND.n3263 GND.n3262 19.3944
R6405 GND.n3262 GND.n3259 19.3944
R6406 GND.n3259 GND.n3258 19.3944
R6407 GND.n3258 GND.n3255 19.3944
R6408 GND.n3255 GND.n3254 19.3944
R6409 GND.n3254 GND.n3251 19.3944
R6410 GND.n3251 GND.n3250 19.3944
R6411 GND.n3250 GND.n3247 19.3944
R6412 GND.n3247 GND.n3246 19.3944
R6413 GND.n3246 GND.n3243 19.3944
R6414 GND.n3243 GND.n3242 19.3944
R6415 GND.n3239 GND.n3238 19.3944
R6416 GND.n3238 GND.n3236 19.3944
R6417 GND.n3236 GND.n3198 19.3944
R6418 GND.n4614 GND.n2075 19.3944
R6419 GND.n4614 GND.n2076 19.3944
R6420 GND.n4610 GND.n2076 19.3944
R6421 GND.n4610 GND.n2078 19.3944
R6422 GND.n2106 GND.n2078 19.3944
R6423 GND.n2106 GND.n2104 19.3944
R6424 GND.n4591 GND.n2104 19.3944
R6425 GND.n4591 GND.n4590 19.3944
R6426 GND.n4590 GND.n4589 19.3944
R6427 GND.n4589 GND.n2112 19.3944
R6428 GND.n4577 GND.n2112 19.3944
R6429 GND.n4577 GND.n4576 19.3944
R6430 GND.n4576 GND.n4575 19.3944
R6431 GND.n4575 GND.n2132 19.3944
R6432 GND.n4563 GND.n2132 19.3944
R6433 GND.n4563 GND.n4562 19.3944
R6434 GND.n4562 GND.n4561 19.3944
R6435 GND.n4561 GND.n2152 19.3944
R6436 GND.n4549 GND.n2152 19.3944
R6437 GND.n4549 GND.n4548 19.3944
R6438 GND.n4548 GND.n4547 19.3944
R6439 GND.n4547 GND.n2172 19.3944
R6440 GND.n4535 GND.n2172 19.3944
R6441 GND.n4535 GND.n4534 19.3944
R6442 GND.n4534 GND.n4533 19.3944
R6443 GND.n4533 GND.n2190 19.3944
R6444 GND.n4521 GND.n2190 19.3944
R6445 GND.n4521 GND.n4520 19.3944
R6446 GND.n4520 GND.n4519 19.3944
R6447 GND.n4519 GND.n2210 19.3944
R6448 GND.n2240 GND.n2210 19.3944
R6449 GND.n2240 GND.n2237 19.3944
R6450 GND.n4500 GND.n2237 19.3944
R6451 GND.n4500 GND.n4499 19.3944
R6452 GND.n4499 GND.n4498 19.3944
R6453 GND.n4498 GND.n2246 19.3944
R6454 GND.n2284 GND.n2246 19.3944
R6455 GND.n2284 GND.n2281 19.3944
R6456 GND.n4480 GND.n2281 19.3944
R6457 GND.n4480 GND.n4479 19.3944
R6458 GND.n4479 GND.n4478 19.3944
R6459 GND.n4478 GND.n2290 19.3944
R6460 GND.n2333 GND.n2290 19.3944
R6461 GND.n2336 GND.n2333 19.3944
R6462 GND.n2336 GND.n2330 19.3944
R6463 GND.n4452 GND.n2330 19.3944
R6464 GND.n4452 GND.n4451 19.3944
R6465 GND.n4451 GND.n4450 19.3944
R6466 GND.n4450 GND.n2342 19.3944
R6467 GND.n3797 GND.n2342 19.3944
R6468 GND.n3797 GND.n2372 19.3944
R6469 GND.n4432 GND.n2372 19.3944
R6470 GND.n4432 GND.n4431 19.3944
R6471 GND.n2816 GND.n2815 19.3944
R6472 GND.n4379 GND.n2815 19.3944
R6473 GND.n4379 GND.n4378 19.3944
R6474 GND.n4378 GND.n4377 19.3944
R6475 GND.n4377 GND.n2822 19.3944
R6476 GND.n4367 GND.n2822 19.3944
R6477 GND.n4367 GND.n4366 19.3944
R6478 GND.n4366 GND.n4365 19.3944
R6479 GND.n4365 GND.n2845 19.3944
R6480 GND.n4355 GND.n2845 19.3944
R6481 GND.n4355 GND.n4354 19.3944
R6482 GND.n4354 GND.n4353 19.3944
R6483 GND.n4353 GND.n2866 19.3944
R6484 GND.n4343 GND.n2866 19.3944
R6485 GND.n4343 GND.n4342 19.3944
R6486 GND.n4342 GND.n4341 19.3944
R6487 GND.n4341 GND.n2888 19.3944
R6488 GND.n4331 GND.n2888 19.3944
R6489 GND.n4331 GND.n4330 19.3944
R6490 GND.n2903 GND.n162 19.3944
R6491 GND.n4317 GND.n162 19.3944
R6492 GND.n5857 GND.n155 19.3944
R6493 GND.n2929 GND.n156 19.3944
R6494 GND.n5854 GND.n164 19.3944
R6495 GND.n5854 GND.n165 19.3944
R6496 GND.n5844 GND.n165 19.3944
R6497 GND.n5844 GND.n5843 19.3944
R6498 GND.n5843 GND.n5842 19.3944
R6499 GND.n5842 GND.n188 19.3944
R6500 GND.n5832 GND.n188 19.3944
R6501 GND.n5832 GND.n5831 19.3944
R6502 GND.n5831 GND.n5830 19.3944
R6503 GND.n5830 GND.n209 19.3944
R6504 GND.n5820 GND.n209 19.3944
R6505 GND.n5820 GND.n5819 19.3944
R6506 GND.n5819 GND.n5818 19.3944
R6507 GND.n5818 GND.n230 19.3944
R6508 GND.n5808 GND.n230 19.3944
R6509 GND.n5808 GND.n5807 19.3944
R6510 GND.n5807 GND.n5806 19.3944
R6511 GND.n5806 GND.n250 19.3944
R6512 GND.n5796 GND.n250 19.3944
R6513 GND.n5796 GND.n5795 19.3944
R6514 GND.n4860 GND.n909 19.3944
R6515 GND.n4854 GND.n909 19.3944
R6516 GND.n4854 GND.n4853 19.3944
R6517 GND.n4853 GND.n4852 19.3944
R6518 GND.n4852 GND.n916 19.3944
R6519 GND.n4846 GND.n916 19.3944
R6520 GND.n4846 GND.n4845 19.3944
R6521 GND.n4845 GND.n4844 19.3944
R6522 GND.n4844 GND.n924 19.3944
R6523 GND.n4838 GND.n924 19.3944
R6524 GND.n4838 GND.n4837 19.3944
R6525 GND.n4837 GND.n4836 19.3944
R6526 GND.n4836 GND.n932 19.3944
R6527 GND.n4830 GND.n932 19.3944
R6528 GND.n4830 GND.n4829 19.3944
R6529 GND.n4829 GND.n4828 19.3944
R6530 GND.n4828 GND.n940 19.3944
R6531 GND.n4822 GND.n940 19.3944
R6532 GND.n4822 GND.n4821 19.3944
R6533 GND.n4821 GND.n4820 19.3944
R6534 GND.n4820 GND.n948 19.3944
R6535 GND.n4814 GND.n948 19.3944
R6536 GND.n4814 GND.n4813 19.3944
R6537 GND.n4813 GND.n4812 19.3944
R6538 GND.n4812 GND.n956 19.3944
R6539 GND.n4806 GND.n956 19.3944
R6540 GND.n4806 GND.n4805 19.3944
R6541 GND.n4805 GND.n4804 19.3944
R6542 GND.n4804 GND.n964 19.3944
R6543 GND.n1747 GND.n964 19.3944
R6544 GND.n1750 GND.n1747 19.3944
R6545 GND.n1750 GND.n1744 19.3944
R6546 GND.n1754 GND.n1744 19.3944
R6547 GND.n1754 GND.n1742 19.3944
R6548 GND.n1774 GND.n1742 19.3944
R6549 GND.n1774 GND.n1740 19.3944
R6550 GND.n1816 GND.n1740 19.3944
R6551 GND.n1816 GND.n1815 19.3944
R6552 GND.n1815 GND.n1814 19.3944
R6553 GND.n1814 GND.n1780 19.3944
R6554 GND.n1810 GND.n1780 19.3944
R6555 GND.n1810 GND.n1809 19.3944
R6556 GND.n1809 GND.n1808 19.3944
R6557 GND.n1808 GND.n1786 19.3944
R6558 GND.n1804 GND.n1786 19.3944
R6559 GND.n1804 GND.n1803 19.3944
R6560 GND.n1803 GND.n1802 19.3944
R6561 GND.n1802 GND.n1792 19.3944
R6562 GND.n1798 GND.n1792 19.3944
R6563 GND.n1798 GND.n1797 19.3944
R6564 GND.n1936 GND.n1591 19.3944
R6565 GND.n1934 GND.n1933 19.3944
R6566 GND.n1614 GND.n1613 19.3944
R6567 GND.n1919 GND.n1918 19.3944
R6568 GND.n1916 GND.n1616 19.3944
R6569 GND.n1664 GND.n1616 19.3944
R6570 GND.n1664 GND.n1663 19.3944
R6571 GND.n1663 GND.n1662 19.3944
R6572 GND.n1662 GND.n1622 19.3944
R6573 GND.n1658 GND.n1622 19.3944
R6574 GND.n1658 GND.n1657 19.3944
R6575 GND.n1657 GND.n1656 19.3944
R6576 GND.n1656 GND.n1628 19.3944
R6577 GND.n1652 GND.n1628 19.3944
R6578 GND.n1652 GND.n1651 19.3944
R6579 GND.n1651 GND.n1650 19.3944
R6580 GND.n1650 GND.n1634 19.3944
R6581 GND.n1646 GND.n1634 19.3944
R6582 GND.n1646 GND.n1645 19.3944
R6583 GND.n1645 GND.n1644 19.3944
R6584 GND.n1644 GND.n1642 19.3944
R6585 GND.n1642 GND.n1491 19.3944
R6586 GND.n1491 GND.n1489 19.3944
R6587 GND.n2045 GND.n1489 19.3944
R6588 GND.n2045 GND.n1487 19.3944
R6589 GND.n4635 GND.n1487 19.3944
R6590 GND.n4635 GND.n4634 19.3944
R6591 GND.n4634 GND.n4633 19.3944
R6592 GND.n4633 GND.n2051 19.3944
R6593 GND.n4627 GND.n2051 19.3944
R6594 GND.n4627 GND.n4626 19.3944
R6595 GND.n4626 GND.n4625 19.3944
R6596 GND.n4625 GND.n2059 19.3944
R6597 GND.n3469 GND.n2059 19.3944
R6598 GND.n3474 GND.n3469 19.3944
R6599 GND.n3474 GND.n2093 19.3944
R6600 GND.n4598 GND.n2093 19.3944
R6601 GND.n4598 GND.n4597 19.3944
R6602 GND.n4597 GND.n4596 19.3944
R6603 GND.n4596 GND.n2097 19.3944
R6604 GND.n3535 GND.n2097 19.3944
R6605 GND.n3535 GND.n3532 19.3944
R6606 GND.n3539 GND.n3532 19.3944
R6607 GND.n3539 GND.n3530 19.3944
R6608 GND.n3551 GND.n3530 19.3944
R6609 GND.n3551 GND.n3550 19.3944
R6610 GND.n3550 GND.n3549 19.3944
R6611 GND.n3549 GND.n3547 19.3944
R6612 GND.n3547 GND.n3155 19.3944
R6613 GND.n3155 GND.n3153 19.3944
R6614 GND.n3589 GND.n3153 19.3944
R6615 GND.n3589 GND.n3151 19.3944
R6616 GND.n3593 GND.n3151 19.3944
R6617 GND.n3593 GND.n3143 19.3944
R6618 GND.n3615 GND.n3143 19.3944
R6619 GND.n3615 GND.n3141 19.3944
R6620 GND.n3628 GND.n3141 19.3944
R6621 GND.n3628 GND.n3627 19.3944
R6622 GND.n3627 GND.n3626 19.3944
R6623 GND.n3626 GND.n3623 19.3944
R6624 GND.n3623 GND.n2217 19.3944
R6625 GND.n4514 GND.n2217 19.3944
R6626 GND.n4514 GND.n4513 19.3944
R6627 GND.n4513 GND.n4512 19.3944
R6628 GND.n4512 GND.n2221 19.3944
R6629 GND.n2265 GND.n2221 19.3944
R6630 GND.n2268 GND.n2265 19.3944
R6631 GND.n2268 GND.n2262 19.3944
R6632 GND.n4487 GND.n2262 19.3944
R6633 GND.n4487 GND.n4486 19.3944
R6634 GND.n4486 GND.n4485 19.3944
R6635 GND.n4485 GND.n2274 19.3944
R6636 GND.n2308 GND.n2274 19.3944
R6637 GND.n2308 GND.n2305 19.3944
R6638 GND.n4466 GND.n2305 19.3944
R6639 GND.n4466 GND.n4465 19.3944
R6640 GND.n4465 GND.n4464 19.3944
R6641 GND.n4464 GND.n2314 19.3944
R6642 GND.n2352 GND.n2314 19.3944
R6643 GND.n2352 GND.n2349 19.3944
R6644 GND.n4445 GND.n2349 19.3944
R6645 GND.n4445 GND.n4444 19.3944
R6646 GND.n4444 GND.n4443 19.3944
R6647 GND.n4443 GND.n2358 19.3944
R6648 GND.n3026 GND.n2358 19.3944
R6649 GND.n4008 GND.n3026 19.3944
R6650 GND.n4008 GND.n3023 19.3944
R6651 GND.n4012 GND.n3023 19.3944
R6652 GND.n4012 GND.n3019 19.3944
R6653 GND.n4019 GND.n3019 19.3944
R6654 GND.n4019 GND.n3017 19.3944
R6655 GND.n4023 GND.n3017 19.3944
R6656 GND.n4023 GND.n3015 19.3944
R6657 GND.n4027 GND.n3015 19.3944
R6658 GND.n4027 GND.n3013 19.3944
R6659 GND.n4031 GND.n3013 19.3944
R6660 GND.n4031 GND.n3011 19.3944
R6661 GND.n4035 GND.n3011 19.3944
R6662 GND.n4035 GND.n3009 19.3944
R6663 GND.n4075 GND.n3009 19.3944
R6664 GND.n4075 GND.n4074 19.3944
R6665 GND.n4074 GND.n4073 19.3944
R6666 GND.n4073 GND.n4041 19.3944
R6667 GND.n4069 GND.n4041 19.3944
R6668 GND.n4069 GND.n4068 19.3944
R6669 GND.n4068 GND.n4067 19.3944
R6670 GND.n4067 GND.n4047 19.3944
R6671 GND.n4063 GND.n4047 19.3944
R6672 GND.n4063 GND.n4062 19.3944
R6673 GND.n4062 GND.n4061 19.3944
R6674 GND.n4061 GND.n4053 19.3944
R6675 GND.n4057 GND.n4053 19.3944
R6676 GND.n4057 GND.n2911 19.3944
R6677 GND.n4325 GND.n2911 19.3944
R6678 GND.n4323 GND.n4322 19.3944
R6679 GND.n2936 GND.n2934 19.3944
R6680 GND.n4306 GND.n2938 19.3944
R6681 GND.n4304 GND.n4303 19.3944
R6682 GND.n4300 GND.n4299 19.3944
R6683 GND.n4299 GND.n4298 19.3944
R6684 GND.n4298 GND.n2943 19.3944
R6685 GND.n4294 GND.n2943 19.3944
R6686 GND.n4294 GND.n4293 19.3944
R6687 GND.n4293 GND.n4292 19.3944
R6688 GND.n4292 GND.n2949 19.3944
R6689 GND.n4288 GND.n2949 19.3944
R6690 GND.n4288 GND.n4287 19.3944
R6691 GND.n4287 GND.n4286 19.3944
R6692 GND.n4286 GND.n2955 19.3944
R6693 GND.n4282 GND.n2955 19.3944
R6694 GND.n4282 GND.n4281 19.3944
R6695 GND.n4281 GND.n4280 19.3944
R6696 GND.n4280 GND.n4269 19.3944
R6697 GND.n4276 GND.n4269 19.3944
R6698 GND.n4276 GND.n4275 19.3944
R6699 GND.n4275 GND.n312 19.3944
R6700 GND.n5745 GND.n312 19.3944
R6701 GND.n5745 GND.n5744 19.3944
R6702 GND.n5744 GND.n5743 19.3944
R6703 GND.n5743 GND.n316 19.3944
R6704 GND.n320 GND.n316 19.3944
R6705 GND.n5736 GND.n320 19.3944
R6706 GND.n5736 GND.n5735 19.3944
R6707 GND.n5735 GND.n5734 19.3944
R6708 GND.n5734 GND.n326 19.3944
R6709 GND.n5728 GND.n326 19.3944
R6710 GND.n5728 GND.n5727 19.3944
R6711 GND.n5727 GND.n5726 19.3944
R6712 GND.n5726 GND.n334 19.3944
R6713 GND.n5720 GND.n334 19.3944
R6714 GND.n5720 GND.n5719 19.3944
R6715 GND.n5719 GND.n5718 19.3944
R6716 GND.n5718 GND.n342 19.3944
R6717 GND.n5712 GND.n342 19.3944
R6718 GND.n5712 GND.n5711 19.3944
R6719 GND.n5711 GND.n5710 19.3944
R6720 GND.n5710 GND.n350 19.3944
R6721 GND.n5704 GND.n350 19.3944
R6722 GND.n5704 GND.n5703 19.3944
R6723 GND.n5703 GND.n5702 19.3944
R6724 GND.n5702 GND.n358 19.3944
R6725 GND.n5696 GND.n358 19.3944
R6726 GND.n5696 GND.n5695 19.3944
R6727 GND.n5695 GND.n5694 19.3944
R6728 GND.n5694 GND.n366 19.3944
R6729 GND.n5688 GND.n366 19.3944
R6730 GND.n5688 GND.n5687 19.3944
R6731 GND.n5687 GND.n5686 19.3944
R6732 GND.n1035 GND.n1032 19.3944
R6733 GND.n1035 GND.n1030 19.3944
R6734 GND.n1039 GND.n1030 19.3944
R6735 GND.n1042 GND.n1039 19.3944
R6736 GND.n1045 GND.n1042 19.3944
R6737 GND.n1045 GND.n1028 19.3944
R6738 GND.n1049 GND.n1028 19.3944
R6739 GND.n1053 GND.n1052 19.3944
R6740 GND.n1056 GND.n1053 19.3944
R6741 GND.n1056 GND.n1022 19.3944
R6742 GND.n1062 GND.n1022 19.3944
R6743 GND.n1063 GND.n1062 19.3944
R6744 GND.n1066 GND.n1063 19.3944
R6745 GND.n1066 GND.n1018 19.3944
R6746 GND.n1070 GND.n1018 19.3944
R6747 GND.n4777 GND.n4776 19.3944
R6748 GND.n4776 GND.n4775 19.3944
R6749 GND.n4775 GND.n1002 19.3944
R6750 GND.n1732 GND.n1002 19.3944
R6751 GND.n1824 GND.n1732 19.3944
R6752 GND.n1824 GND.n1729 19.3944
R6753 GND.n1830 GND.n1729 19.3944
R6754 GND.n1830 GND.n1829 19.3944
R6755 GND.n1829 GND.n1708 19.3944
R6756 GND.n1849 GND.n1708 19.3944
R6757 GND.n1849 GND.n1706 19.3944
R6758 GND.n1855 GND.n1706 19.3944
R6759 GND.n1855 GND.n1854 19.3944
R6760 GND.n1854 GND.n1686 19.3944
R6761 GND.n1874 GND.n1686 19.3944
R6762 GND.n1874 GND.n1684 19.3944
R6763 GND.n1878 GND.n1684 19.3944
R6764 GND.n1878 GND.n1578 19.3944
R6765 GND.n1945 GND.n1578 19.3944
R6766 GND.n1577 GND.n1576 19.3944
R6767 GND.n1602 GND.n1576 19.3944
R6768 GND.n1928 GND.n1927 19.3944
R6769 GND.n1904 GND.n1903 19.3944
R6770 GND.n1906 GND.n1570 19.3944
R6771 GND.n1951 GND.n1570 19.3944
R6772 GND.n1951 GND.n1950 19.3944
R6773 GND.n1950 GND.n1550 19.3944
R6774 GND.n1970 GND.n1550 19.3944
R6775 GND.n1970 GND.n1548 19.3944
R6776 GND.n1976 GND.n1548 19.3944
R6777 GND.n1976 GND.n1975 19.3944
R6778 GND.n1975 GND.n1527 19.3944
R6779 GND.n1994 GND.n1527 19.3944
R6780 GND.n1994 GND.n1525 19.3944
R6781 GND.n2000 GND.n1525 19.3944
R6782 GND.n2000 GND.n1999 19.3944
R6783 GND.n1999 GND.n1504 19.3944
R6784 GND.n2028 GND.n1504 19.3944
R6785 GND.n2028 GND.n1502 19.3944
R6786 GND.n2034 GND.n1502 19.3944
R6787 GND.n2034 GND.n2033 19.3944
R6788 GND.n2033 GND.n1177 19.3944
R6789 GND.n4698 GND.n1177 19.3944
R6790 GND.n4968 GND.n802 19.3944
R6791 GND.n4968 GND.n4967 19.3944
R6792 GND.n4967 GND.n4966 19.3944
R6793 GND.n4966 GND.n806 19.3944
R6794 GND.n4960 GND.n806 19.3944
R6795 GND.n4960 GND.n4959 19.3944
R6796 GND.n4959 GND.n4958 19.3944
R6797 GND.n4958 GND.n814 19.3944
R6798 GND.n4952 GND.n814 19.3944
R6799 GND.n4952 GND.n4951 19.3944
R6800 GND.n4951 GND.n4950 19.3944
R6801 GND.n4950 GND.n822 19.3944
R6802 GND.n4944 GND.n822 19.3944
R6803 GND.n4944 GND.n4943 19.3944
R6804 GND.n4943 GND.n4942 19.3944
R6805 GND.n4942 GND.n830 19.3944
R6806 GND.n4936 GND.n830 19.3944
R6807 GND.n4936 GND.n4935 19.3944
R6808 GND.n4935 GND.n4934 19.3944
R6809 GND.n4934 GND.n838 19.3944
R6810 GND.n4928 GND.n838 19.3944
R6811 GND.n4928 GND.n4927 19.3944
R6812 GND.n4927 GND.n4926 19.3944
R6813 GND.n4926 GND.n846 19.3944
R6814 GND.n4920 GND.n846 19.3944
R6815 GND.n4920 GND.n4919 19.3944
R6816 GND.n4919 GND.n4918 19.3944
R6817 GND.n4918 GND.n854 19.3944
R6818 GND.n4912 GND.n854 19.3944
R6819 GND.n4912 GND.n4911 19.3944
R6820 GND.n4911 GND.n4910 19.3944
R6821 GND.n4910 GND.n862 19.3944
R6822 GND.n4904 GND.n862 19.3944
R6823 GND.n4904 GND.n4903 19.3944
R6824 GND.n4903 GND.n4902 19.3944
R6825 GND.n4902 GND.n870 19.3944
R6826 GND.n4896 GND.n870 19.3944
R6827 GND.n4896 GND.n4895 19.3944
R6828 GND.n4895 GND.n4894 19.3944
R6829 GND.n4894 GND.n878 19.3944
R6830 GND.n4888 GND.n878 19.3944
R6831 GND.n4888 GND.n4887 19.3944
R6832 GND.n4887 GND.n4886 19.3944
R6833 GND.n4886 GND.n886 19.3944
R6834 GND.n4880 GND.n886 19.3944
R6835 GND.n4880 GND.n4879 19.3944
R6836 GND.n4879 GND.n4878 19.3944
R6837 GND.n4878 GND.n894 19.3944
R6838 GND.n4872 GND.n894 19.3944
R6839 GND.n4872 GND.n4871 19.3944
R6840 GND.n4871 GND.n4870 19.3944
R6841 GND.n4870 GND.n902 19.3944
R6842 GND.n4864 GND.n902 19.3944
R6843 GND.n4864 GND.n4863 19.3944
R6844 GND.n4798 GND.n4797 19.3944
R6845 GND.n4797 GND.n984 19.3944
R6846 GND.n4793 GND.n984 19.3944
R6847 GND.n4793 GND.n4792 19.3944
R6848 GND.n4792 GND.n4791 19.3944
R6849 GND.n4791 GND.n990 19.3944
R6850 GND.n1763 GND.n993 19.3944
R6851 GND.n1764 GND.n1763 19.3944
R6852 GND.n1764 GND.n1759 19.3944
R6853 GND.n1769 GND.n1759 19.3944
R6854 GND.n1769 GND.n1760 19.3944
R6855 GND.n1760 GND.n1720 19.3944
R6856 GND.n1834 GND.n1720 19.3944
R6857 GND.n1834 GND.n1717 19.3944
R6858 GND.n1839 GND.n1717 19.3944
R6859 GND.n1839 GND.n1718 19.3944
R6860 GND.n1718 GND.n1697 19.3944
R6861 GND.n1859 GND.n1697 19.3944
R6862 GND.n1859 GND.n1694 19.3944
R6863 GND.n1864 GND.n1694 19.3944
R6864 GND.n1864 GND.n1695 19.3944
R6865 GND.n1695 GND.n1675 19.3944
R6866 GND.n1882 GND.n1675 19.3944
R6867 GND.n1882 GND.n1673 19.3944
R6868 GND.n1886 GND.n1673 19.3944
R6869 GND.n1887 GND.n1886 19.3944
R6870 GND.n1890 GND.n1887 19.3944
R6871 GND.n1890 GND.n1671 19.3944
R6872 GND.n1895 GND.n1671 19.3944
R6873 GND.n1896 GND.n1895 19.3944
R6874 GND.n1897 GND.n1896 19.3944
R6875 GND.n1897 GND.n1669 19.3944
R6876 GND.n1901 GND.n1669 19.3944
R6877 GND.n1901 GND.n1562 19.3944
R6878 GND.n1955 GND.n1562 19.3944
R6879 GND.n1955 GND.n1559 19.3944
R6880 GND.n1960 GND.n1559 19.3944
R6881 GND.n1960 GND.n1560 19.3944
R6882 GND.n1560 GND.n1540 19.3944
R6883 GND.n1980 GND.n1540 19.3944
R6884 GND.n1980 GND.n1537 19.3944
R6885 GND.n1985 GND.n1537 19.3944
R6886 GND.n1985 GND.n1538 19.3944
R6887 GND.n1538 GND.n1516 19.3944
R6888 GND.n2004 GND.n1516 19.3944
R6889 GND.n2004 GND.n1513 19.3944
R6890 GND.n2021 GND.n1513 19.3944
R6891 GND.n2021 GND.n1514 19.3944
R6892 GND.n2017 GND.n1514 19.3944
R6893 GND.n2017 GND.n2016 19.3944
R6894 GND.n2016 GND.n2015 19.3944
R6895 GND.n2015 GND.n2012 19.3944
R6896 GND.n2012 GND.n2011 19.3944
R6897 GND.n1466 GND.n1465 18.7521
R6898 GND.n1822 GND.t96 18.6358
R6899 GND.n4623 GND.n2061 18.6358
R6900 GND.n5810 GND.t73 18.6358
R6901 GND.n4688 GND.n4687 18.6187
R6902 GND.n4414 GND.n4413 18.6187
R6903 GND.n4658 GND.n1473 18.4247
R6904 GND.n4241 GND.n4240 18.4247
R6905 GND.n2789 GND.n2379 18.4247
R6906 GND.n4787 GND.n990 18.4247
R6907 GND.n2785 GND.n2467 17.6668
R6908 GND.n1466 GND.n1244 17.3295
R6909 GND.n4801 GND.n4800 17.2554
R6910 GND.n4800 GND.n980 17.2554
R6911 GND.n4616 GND.n2069 17.2554
R6912 GND.n4616 GND.n2072 17.2554
R6913 GND.n4600 GND.n2090 17.2554
R6914 GND.n4594 GND.n4593 17.2554
R6915 GND.n4587 GND.n2114 17.2554
R6916 GND.n3515 GND.n2123 17.2554
R6917 GND.n3554 GND.n3553 17.2554
R6918 GND.n3563 GND.n2143 17.2554
R6919 GND.n3585 GND.n3584 17.2554
R6920 GND.n3578 GND.n2157 17.2554
R6921 GND.n3578 GND.n2163 17.2554
R6922 GND.n3149 GND.n3148 17.2554
R6923 GND.n3145 GND.n2177 17.2554
R6924 GND.n3634 GND.n3137 17.2554
R6925 GND.n3659 GND.n2195 17.2554
R6926 GND.n4523 GND.n2204 17.2554
R6927 GND.n4517 GND.n4516 17.2554
R6928 GND.n4510 GND.n2223 17.2554
R6929 GND.n4502 GND.n2234 17.2554
R6930 GND.n4496 GND.n2248 17.2554
R6931 GND.n4496 GND.n2251 17.2554
R6932 GND.n4489 GND.n2259 17.2554
R6933 GND.n4483 GND.n4482 17.2554
R6934 GND.n4476 GND.n2292 17.2554
R6935 GND.n4468 GND.n2302 17.2554
R6936 GND.n4462 GND.n2316 17.2554
R6937 GND.n4454 GND.n2327 17.2554
R6938 GND.n4448 GND.n4447 17.2554
R6939 GND.n4434 GND.n2367 17.2554
R6940 GND.n5790 GND.n272 17.2554
R6941 GND.n5790 GND.n278 17.2554
R6942 GND.n1429 GND.n1428 16.7936
R6943 GND.n1295 GND.n1293 16.778
R6944 GND.n3507 GND.n3506 16.5652
R6945 GND.n4580 GND.n4579 16.5652
R6946 GND.n4531 GND.n4530 16.5652
R6947 GND.n3130 GND.n3129 16.5652
R6948 GND.n4469 GND.n2300 16.5652
R6949 GND.n4461 GND.n2318 16.5652
R6950 GND.n3476 GND.t41 16.2201
R6951 GND.n4441 GND.t51 16.2201
R6952 GND.n2023 GND.t55 15.875
R6953 GND.n4607 GND.n2082 15.875
R6954 GND.n3159 GND.n3156 15.875
R6955 GND.n3598 GND.n3595 15.875
R6956 GND.n4503 GND.n2231 15.875
R6957 GND.n3116 GND.n3115 15.875
R6958 GND.n3793 GND.n3096 15.875
R6959 GND.n4005 GND.n3030 15.875
R6960 GND.n4369 GND.t37 15.875
R6961 GND.n3327 GND.n3324 15.8238
R6962 GND.n1294 GND.n1246 15.7648
R6963 GND.n51 GND.n50 15.3979
R6964 GND.n62 GND.n61 15.3979
R6965 GND.n27 GND.n26 15.3979
R6966 GND.n38 GND.n37 15.3979
R6967 GND.n4 GND.n3 15.3979
R6968 GND.n15 GND.n14 15.3979
R6969 GND.n134 GND.n133 15.3979
R6970 GND.n123 GND.n122 15.3979
R6971 GND.n110 GND.n109 15.3979
R6972 GND.n99 GND.n98 15.3979
R6973 GND.n87 GND.n86 15.3979
R6974 GND.n76 GND.n75 15.3979
R6975 GND.n3489 GND.n2099 15.1848
R6976 GND.n4573 GND.n2134 15.1848
R6977 GND.n3747 GND.n3746 15.1848
R6978 GND.n3768 GND.n3101 15.1848
R6979 GND.n3039 GND.n3038 14.6967
R6980 GND.n3334 GND.n3333 14.6737
R6981 GND.n4002 GND.n4001 14.6737
R6982 GND.n3192 GND.n3191 14.4946
R6983 GND.n3564 GND.n2137 14.4946
R6984 GND.n3613 GND.n3612 14.4946
R6985 GND.n3680 GND.n3679 14.4946
R6986 GND.n3109 GND.n2278 14.4946
R6987 GND.n3769 GND.n2344 14.4946
R6988 GND.n4674 GND.n1204 14.1581
R6989 GND.n4396 GND.n2422 14.1581
R6990 GND.n5758 GND.n5755 14.1581
R6991 GND.n1071 GND.n1070 14.1581
R6992 GND.n4779 GND.n994 13.8044
R6993 GND.n1078 GND.n996 13.8044
R6994 GND.n4773 GND.n1004 13.8044
R6995 GND.n1757 GND.n1007 13.8044
R6996 GND.n1772 GND.n1771 13.8044
R6997 GND.n1822 GND.n1734 13.8044
R6998 GND.n1819 GND.n1818 13.8044
R6999 GND.n1832 GND.n1722 13.8044
R7000 GND.n1727 GND.n1723 13.8044
R7001 GND.n1841 GND.n1714 13.8044
R7002 GND.n1847 GND.n1710 13.8044
R7003 GND.n1844 GND.n1712 13.8044
R7004 GND.n1857 GND.n1699 13.8044
R7005 GND.n1704 GND.n1700 13.8044
R7006 GND.n1866 GND.n1692 13.8044
R7007 GND.n1872 GND.n1688 13.8044
R7008 GND.n1868 GND.n1690 13.8044
R7009 GND.n1880 GND.n1678 13.8044
R7010 GND.n1681 GND.n1680 13.8044
R7011 GND.n1943 GND.n1581 13.8044
R7012 GND.n1939 GND.n1583 13.8044
R7013 GND.n1938 GND.n1588 13.8044
R7014 GND.n1595 GND.n1594 13.8044
R7015 GND.n1931 GND.n1930 13.8044
R7016 GND.n1925 GND.n1597 13.8044
R7017 GND.n1922 GND.n1606 13.8044
R7018 GND.n1921 GND.n1610 13.8044
R7019 GND.n1908 GND.n1667 13.8044
R7020 GND.n1914 GND.n1913 13.8044
R7021 GND.n1568 GND.n1565 13.8044
R7022 GND.n1962 GND.n1557 13.8044
R7023 GND.n1968 GND.n1552 13.8044
R7024 GND.n1965 GND.n1554 13.8044
R7025 GND.n1978 GND.n1542 13.8044
R7026 GND.n1546 GND.n1543 13.8044
R7027 GND.n1987 GND.n1535 13.8044
R7028 GND.n1992 GND.n1529 13.8044
R7029 GND.n1989 GND.n1532 13.8044
R7030 GND.n2002 GND.n1518 13.8044
R7031 GND.n1523 GND.n1519 13.8044
R7032 GND.n2023 GND.n1510 13.8044
R7033 GND.n2026 GND.n1506 13.8044
R7034 GND.n2008 GND.n1508 13.8044
R7035 GND.n2036 GND.n1497 13.8044
R7036 GND.n1499 GND.n1493 13.8044
R7037 GND.n2041 GND.n2040 13.8044
R7038 GND.n4700 GND.n1170 13.8044
R7039 GND.n4601 GND.n2088 13.8044
R7040 GND.n4566 GND.n4565 13.8044
R7041 GND.n4545 GND.n4544 13.8044
R7042 GND.n4509 GND.n2225 13.8044
R7043 GND.n3710 GND.n2276 13.8044
R7044 GND.n3772 GND.n2346 13.8044
R7045 GND.n4006 GND.t100 13.8044
R7046 GND.n4389 GND.n2427 13.8044
R7047 GND.n2994 GND.n2809 13.8044
R7048 GND.n4381 GND.n2811 13.8044
R7049 GND.n2999 GND.n2824 13.8044
R7050 GND.n4375 GND.n2827 13.8044
R7051 GND.n4078 GND.n4077 13.8044
R7052 GND.n4369 GND.n2839 13.8044
R7053 GND.n4085 GND.n2847 13.8044
R7054 GND.n4363 GND.n2850 13.8044
R7055 GND.n4093 GND.n2857 13.8044
R7056 GND.n4357 GND.n2860 13.8044
R7057 GND.n4100 GND.n2868 13.8044
R7058 GND.n4351 GND.n2871 13.8044
R7059 GND.n4108 GND.n2878 13.8044
R7060 GND.n4345 GND.n2881 13.8044
R7061 GND.n4115 GND.n2890 13.8044
R7062 GND.n4339 GND.n2893 13.8044
R7063 GND.n4135 GND.n2900 13.8044
R7064 GND.n4328 GND.n4327 13.8044
R7065 GND.n2914 GND.n2908 13.8044
R7066 GND.n4320 GND.n2915 13.8044
R7067 GND.n4319 GND.n2918 13.8044
R7068 GND.n4149 GND.n149 13.8044
R7069 GND.n5859 GND.n151 13.8044
R7070 GND.n4309 GND.n4308 13.8044
R7071 GND.n4158 GND.n2931 13.8044
R7072 GND.n4165 GND.n168 13.8044
R7073 GND.n5852 GND.n171 13.8044
R7074 GND.n4171 GND.n180 13.8044
R7075 GND.n5846 GND.n183 13.8044
R7076 GND.n4179 GND.n190 13.8044
R7077 GND.n5840 GND.n193 13.8044
R7078 GND.n4185 GND.n200 13.8044
R7079 GND.n5834 GND.n203 13.8044
R7080 GND.n4193 GND.n211 13.8044
R7081 GND.n5828 GND.n214 13.8044
R7082 GND.n4199 GND.n221 13.8044
R7083 GND.n5822 GND.n224 13.8044
R7084 GND.n4208 GND.n232 13.8044
R7085 GND.n5816 GND.n235 13.8044
R7086 GND.n4263 GND.n4262 13.8044
R7087 GND.n5810 GND.n244 13.8044
R7088 GND.n4256 GND.n252 13.8044
R7089 GND.n5804 GND.n255 13.8044
R7090 GND.n4250 GND.n262 13.8044
R7091 GND.n5798 GND.n265 13.8044
R7092 GND.n5748 GND.n5747 13.8044
R7093 GND.n1292 GND.n1247 13.4981
R7094 GND.n3332 GND.n3323 13.1884
R7095 GND.n2754 GND.n2753 13.1807
R7096 GND.n2719 GND.n2718 13.1807
R7097 GND.n2684 GND.n2683 13.1807
R7098 GND.n2650 GND.n2649 13.1807
R7099 GND.n2615 GND.n2614 13.1807
R7100 GND.n2580 GND.n2579 13.1807
R7101 GND.n2545 GND.n2544 13.1807
R7102 GND.n2511 GND.n2510 13.1807
R7103 GND.t103 GND.n2061 13.1142
R7104 GND.n3185 GND.n2101 13.1142
R7105 GND.n3633 GND.n3630 13.1142
R7106 GND.n3670 GND.n2212 13.1142
R7107 GND.n4455 GND.n2324 13.1142
R7108 GND.n54 GND.n49 12.8005
R7109 GND.n65 GND.n60 12.8005
R7110 GND.n30 GND.n25 12.8005
R7111 GND.n41 GND.n36 12.8005
R7112 GND.n7 GND.n2 12.8005
R7113 GND.n18 GND.n13 12.8005
R7114 GND.n1462 GND.n1432 12.8005
R7115 GND.n1240 GND.n1210 12.8005
R7116 GND.n137 GND.n132 12.8005
R7117 GND.n126 GND.n121 12.8005
R7118 GND.n113 GND.n108 12.8005
R7119 GND.n102 GND.n97 12.8005
R7120 GND.n90 GND.n85 12.8005
R7121 GND.n79 GND.n74 12.8005
R7122 GND.n2498 GND.n2468 12.8005
R7123 GND.n2463 GND.n2433 12.8005
R7124 GND.t22 GND.n1581 12.424
R7125 GND.n4622 GND.n2063 12.424
R7126 GND.n3478 GND.n3477 12.424
R7127 GND.n4559 GND.n2154 12.424
R7128 GND.n4551 GND.n2166 12.424
R7129 GND.n3698 GND.n3122 12.424
R7130 GND.n4490 GND.n2257 12.424
R7131 GND.n4440 GND.n2361 12.424
R7132 GND.n3890 GND.n3028 12.424
R7133 GND.t29 GND.n171 12.424
R7134 GND.n2782 GND.n2781 12.3289
R7135 GND.n2763 GND.n2762 12.1722
R7136 GND.n2762 GND.n2761 12.1722
R7137 GND.n2728 GND.n2727 12.1722
R7138 GND.n2727 GND.n2726 12.1722
R7139 GND.n2693 GND.n2692 12.1722
R7140 GND.n2692 GND.n2691 12.1722
R7141 GND.n2659 GND.n2658 12.1722
R7142 GND.n2658 GND.n2657 12.1722
R7143 GND.n2623 GND.n2622 12.1722
R7144 GND.n2624 GND.n2623 12.1722
R7145 GND.n2588 GND.n2587 12.1722
R7146 GND.n2589 GND.n2588 12.1722
R7147 GND.n2553 GND.n2552 12.1722
R7148 GND.n2554 GND.n2553 12.1722
R7149 GND.n2519 GND.n2518 12.1722
R7150 GND.n2520 GND.n2519 12.1722
R7151 GND.n55 GND.n47 12.0247
R7152 GND.n66 GND.n58 12.0247
R7153 GND.n31 GND.n23 12.0247
R7154 GND.n42 GND.n34 12.0247
R7155 GND.n8 GND.n0 12.0247
R7156 GND.n19 GND.n11 12.0247
R7157 GND.n1461 GND.n1434 12.0247
R7158 GND.n1239 GND.n1212 12.0247
R7159 GND.n138 GND.n130 12.0247
R7160 GND.n127 GND.n119 12.0247
R7161 GND.n114 GND.n106 12.0247
R7162 GND.n103 GND.n95 12.0247
R7163 GND.n91 GND.n83 12.0247
R7164 GND.n80 GND.n72 12.0247
R7165 GND.n2497 GND.n2470 12.0247
R7166 GND.n2462 GND.n2435 12.0247
R7167 GND.n4670 GND.n1204 11.8308
R7168 GND.n4392 GND.n2422 11.8308
R7169 GND.n5755 GND.n303 11.8308
R7170 GND.n1072 GND.n1071 11.8308
R7171 GND.n4586 GND.n2117 11.7338
R7172 GND.n3516 GND.n2117 11.7338
R7173 GND.n3660 GND.n2201 11.7338
R7174 GND.n4524 GND.n2201 11.7338
R7175 GND.n3735 GND.n3734 11.7338
R7176 GND.n3734 GND.n3733 11.7338
R7177 GND.n2781 GND.n2501 11.4887
R7178 GND.n1458 GND.n1457 11.249
R7179 GND.n1236 GND.n1235 11.249
R7180 GND.n2494 GND.n2493 11.249
R7181 GND.n2459 GND.n2458 11.249
R7182 GND.t5 GND.n3526 11.0436
R7183 GND.n4552 GND.n4551 11.0436
R7184 GND.n3698 GND.n3697 11.0436
R7185 GND.n4475 GND.t16 11.0436
R7186 GND.n3787 GND.n2361 11.0436
R7187 GND.n3891 GND.n3890 11.0436
R7188 GND.n71 GND.n70 10.833
R7189 GND.n5864 GND.n142 10.833
R7190 GND.n3945 GND.n3944 10.6151
R7191 GND.n3944 GND.n3943 10.6151
R7192 GND.n3943 GND.n3066 10.6151
R7193 GND.n3938 GND.n3937 10.6151
R7194 GND.n3937 GND.n3936 10.6151
R7195 GND.n3936 GND.n3072 10.6151
R7196 GND.n3931 GND.n3072 10.6151
R7197 GND.n3931 GND.n3930 10.6151
R7198 GND.n3930 GND.n3929 10.6151
R7199 GND.n3929 GND.n3075 10.6151
R7200 GND.n3924 GND.n3075 10.6151
R7201 GND.n3924 GND.n3923 10.6151
R7202 GND.n3923 GND.n3922 10.6151
R7203 GND.n3922 GND.n3078 10.6151
R7204 GND.n3917 GND.n3078 10.6151
R7205 GND.n3917 GND.n3916 10.6151
R7206 GND.n3916 GND.n3915 10.6151
R7207 GND.n3915 GND.n3081 10.6151
R7208 GND.n3910 GND.n3081 10.6151
R7209 GND.n3910 GND.n3909 10.6151
R7210 GND.n3909 GND.n3908 10.6151
R7211 GND.n3908 GND.n3084 10.6151
R7212 GND.n3903 GND.n3084 10.6151
R7213 GND.n3903 GND.n3902 10.6151
R7214 GND.n3902 GND.n3901 10.6151
R7215 GND.n3901 GND.n3087 10.6151
R7216 GND.n3896 GND.n3087 10.6151
R7217 GND.n3454 GND.n3453 10.6151
R7218 GND.n3457 GND.n3454 10.6151
R7219 GND.n3458 GND.n3457 10.6151
R7220 GND.n3459 GND.n3458 10.6151
R7221 GND.n3466 GND.n3459 10.6151
R7222 GND.n3466 GND.n3465 10.6151
R7223 GND.n3465 GND.n3464 10.6151
R7224 GND.n3464 GND.n3461 10.6151
R7225 GND.n3461 GND.n3460 10.6151
R7226 GND.n3460 GND.n3190 10.6151
R7227 GND.n3190 GND.n3188 10.6151
R7228 GND.n3502 GND.n3188 10.6151
R7229 GND.n3503 GND.n3502 10.6151
R7230 GND.n3504 GND.n3503 10.6151
R7231 GND.n3504 GND.n3181 10.6151
R7232 GND.n3518 GND.n3181 10.6151
R7233 GND.n3519 GND.n3518 10.6151
R7234 GND.n3520 GND.n3519 10.6151
R7235 GND.n3522 GND.n3520 10.6151
R7236 GND.n3522 GND.n3521 10.6151
R7237 GND.n3521 GND.n3175 10.6151
R7238 GND.n3566 GND.n3175 10.6151
R7239 GND.n3567 GND.n3566 10.6151
R7240 GND.n3568 GND.n3567 10.6151
R7241 GND.n3568 GND.n3174 10.6151
R7242 GND.n3572 GND.n3174 10.6151
R7243 GND.n3573 GND.n3572 10.6151
R7244 GND.n3576 GND.n3573 10.6151
R7245 GND.n3576 GND.n3575 10.6151
R7246 GND.n3575 GND.n3574 10.6151
R7247 GND.n3574 GND.n3146 10.6151
R7248 GND.n3601 GND.n3146 10.6151
R7249 GND.n3602 GND.n3601 10.6151
R7250 GND.n3610 GND.n3602 10.6151
R7251 GND.n3610 GND.n3609 10.6151
R7252 GND.n3609 GND.n3608 10.6151
R7253 GND.n3608 GND.n3605 10.6151
R7254 GND.n3605 GND.n3604 10.6151
R7255 GND.n3604 GND.n3133 10.6151
R7256 GND.n3662 GND.n3133 10.6151
R7257 GND.n3663 GND.n3662 10.6151
R7258 GND.n3664 GND.n3663 10.6151
R7259 GND.n3668 GND.n3664 10.6151
R7260 GND.n3668 GND.n3667 10.6151
R7261 GND.n3667 GND.n3666 10.6151
R7262 GND.n3666 GND.n3124 10.6151
R7263 GND.n3682 GND.n3124 10.6151
R7264 GND.n3683 GND.n3682 10.6151
R7265 GND.n3686 GND.n3683 10.6151
R7266 GND.n3687 GND.n3686 10.6151
R7267 GND.n3688 GND.n3687 10.6151
R7268 GND.n3695 GND.n3688 10.6151
R7269 GND.n3695 GND.n3694 10.6151
R7270 GND.n3694 GND.n3693 10.6151
R7271 GND.n3693 GND.n3690 10.6151
R7272 GND.n3690 GND.n3689 10.6151
R7273 GND.n3689 GND.n3114 10.6151
R7274 GND.n3114 GND.n3112 10.6151
R7275 GND.n3723 GND.n3112 10.6151
R7276 GND.n3724 GND.n3723 10.6151
R7277 GND.n3744 GND.n3724 10.6151
R7278 GND.n3744 GND.n3743 10.6151
R7279 GND.n3743 GND.n3742 10.6151
R7280 GND.n3742 GND.n3738 10.6151
R7281 GND.n3738 GND.n3737 10.6151
R7282 GND.n3737 GND.n3731 10.6151
R7283 GND.n3731 GND.n3730 10.6151
R7284 GND.n3730 GND.n3729 10.6151
R7285 GND.n3729 GND.n3726 10.6151
R7286 GND.n3726 GND.n3725 10.6151
R7287 GND.n3725 GND.n3100 10.6151
R7288 GND.n3100 GND.n3098 10.6151
R7289 GND.n3784 GND.n3098 10.6151
R7290 GND.n3785 GND.n3784 10.6151
R7291 GND.n3791 GND.n3785 10.6151
R7292 GND.n3791 GND.n3790 10.6151
R7293 GND.n3790 GND.n3789 10.6151
R7294 GND.n3789 GND.n3786 10.6151
R7295 GND.n3786 GND.n3089 10.6151
R7296 GND.n3894 GND.n3089 10.6151
R7297 GND.n3895 GND.n3894 10.6151
R7298 GND.n3398 GND.n3397 10.6151
R7299 GND.n3399 GND.n3398 10.6151
R7300 GND.n3399 GND.n3304 10.6151
R7301 GND.n3406 GND.n3405 10.6151
R7302 GND.n3407 GND.n3406 10.6151
R7303 GND.n3407 GND.n3299 10.6151
R7304 GND.n3413 GND.n3299 10.6151
R7305 GND.n3414 GND.n3413 10.6151
R7306 GND.n3415 GND.n3414 10.6151
R7307 GND.n3415 GND.n3297 10.6151
R7308 GND.n3421 GND.n3297 10.6151
R7309 GND.n3422 GND.n3421 10.6151
R7310 GND.n3423 GND.n3422 10.6151
R7311 GND.n3423 GND.n3295 10.6151
R7312 GND.n3429 GND.n3295 10.6151
R7313 GND.n3430 GND.n3429 10.6151
R7314 GND.n3431 GND.n3430 10.6151
R7315 GND.n3431 GND.n3293 10.6151
R7316 GND.n3437 GND.n3293 10.6151
R7317 GND.n3438 GND.n3437 10.6151
R7318 GND.n3439 GND.n3438 10.6151
R7319 GND.n3439 GND.n3291 10.6151
R7320 GND.n3445 GND.n3291 10.6151
R7321 GND.n3446 GND.n3445 10.6151
R7322 GND.n3447 GND.n3446 10.6151
R7323 GND.n3447 GND.n3289 10.6151
R7324 GND.n3289 GND.n3288 10.6151
R7325 GND.n3338 GND.n3334 10.6151
R7326 GND.n3339 GND.n3338 10.6151
R7327 GND.n3340 GND.n3339 10.6151
R7328 GND.n3340 GND.n3321 10.6151
R7329 GND.n3346 GND.n3321 10.6151
R7330 GND.n3347 GND.n3346 10.6151
R7331 GND.n3348 GND.n3347 10.6151
R7332 GND.n3348 GND.n3319 10.6151
R7333 GND.n3354 GND.n3319 10.6151
R7334 GND.n3355 GND.n3354 10.6151
R7335 GND.n3356 GND.n3355 10.6151
R7336 GND.n3356 GND.n3317 10.6151
R7337 GND.n3362 GND.n3317 10.6151
R7338 GND.n3363 GND.n3362 10.6151
R7339 GND.n3364 GND.n3363 10.6151
R7340 GND.n3364 GND.n3315 10.6151
R7341 GND.n3370 GND.n3315 10.6151
R7342 GND.n3371 GND.n3370 10.6151
R7343 GND.n3372 GND.n3371 10.6151
R7344 GND.n3372 GND.n3313 10.6151
R7345 GND.n3378 GND.n3313 10.6151
R7346 GND.n3379 GND.n3378 10.6151
R7347 GND.n3380 GND.n3379 10.6151
R7348 GND.n3380 GND.n3311 10.6151
R7349 GND.n3387 GND.n3386 10.6151
R7350 GND.n3388 GND.n3387 10.6151
R7351 GND.n3388 GND.n3306 10.6151
R7352 GND.n4001 GND.n4000 10.6151
R7353 GND.n4000 GND.n3043 10.6151
R7354 GND.n3995 GND.n3043 10.6151
R7355 GND.n3995 GND.n3994 10.6151
R7356 GND.n3994 GND.n3993 10.6151
R7357 GND.n3993 GND.n3046 10.6151
R7358 GND.n3988 GND.n3046 10.6151
R7359 GND.n3988 GND.n3987 10.6151
R7360 GND.n3987 GND.n3986 10.6151
R7361 GND.n3986 GND.n3049 10.6151
R7362 GND.n3981 GND.n3049 10.6151
R7363 GND.n3981 GND.n3980 10.6151
R7364 GND.n3980 GND.n3979 10.6151
R7365 GND.n3979 GND.n3052 10.6151
R7366 GND.n3974 GND.n3052 10.6151
R7367 GND.n3974 GND.n3973 10.6151
R7368 GND.n3973 GND.n3972 10.6151
R7369 GND.n3972 GND.n3055 10.6151
R7370 GND.n3967 GND.n3055 10.6151
R7371 GND.n3967 GND.n3966 10.6151
R7372 GND.n3966 GND.n3965 10.6151
R7373 GND.n3965 GND.n3058 10.6151
R7374 GND.n3960 GND.n3058 10.6151
R7375 GND.n3960 GND.n3959 10.6151
R7376 GND.n3957 GND.n3063 10.6151
R7377 GND.n3952 GND.n3063 10.6151
R7378 GND.n3952 GND.n3951 10.6151
R7379 GND.n4620 GND.n2066 10.6151
R7380 GND.n4620 GND.n4619 10.6151
R7381 GND.n4619 GND.n4618 10.6151
R7382 GND.n4618 GND.n2067 10.6151
R7383 GND.n2085 GND.n2067 10.6151
R7384 GND.n4605 GND.n2085 10.6151
R7385 GND.n4605 GND.n4604 10.6151
R7386 GND.n4604 GND.n4603 10.6151
R7387 GND.n4603 GND.n2086 10.6151
R7388 GND.n3496 GND.n2086 10.6151
R7389 GND.n3496 GND.n3495 10.6151
R7390 GND.n3495 GND.n3494 10.6151
R7391 GND.n3494 GND.n3491 10.6151
R7392 GND.n3491 GND.n2120 10.6151
R7393 GND.n4584 GND.n2120 10.6151
R7394 GND.n4584 GND.n4583 10.6151
R7395 GND.n4583 GND.n4582 10.6151
R7396 GND.n4582 GND.n2121 10.6151
R7397 GND.n3524 GND.n2121 10.6151
R7398 GND.n3524 GND.n2140 10.6151
R7399 GND.n4570 GND.n2140 10.6151
R7400 GND.n4570 GND.n4569 10.6151
R7401 GND.n4569 GND.n4568 10.6151
R7402 GND.n4568 GND.n2141 10.6151
R7403 GND.n3157 GND.n2141 10.6151
R7404 GND.n3157 GND.n2160 10.6151
R7405 GND.n4556 GND.n2160 10.6151
R7406 GND.n4556 GND.n4555 10.6151
R7407 GND.n4555 GND.n4554 10.6151
R7408 GND.n4554 GND.n2161 10.6151
R7409 GND.n3596 GND.n2161 10.6151
R7410 GND.n3596 GND.n2180 10.6151
R7411 GND.n4542 GND.n2180 10.6151
R7412 GND.n4542 GND.n4541 10.6151
R7413 GND.n4541 GND.n4540 10.6151
R7414 GND.n4540 GND.n2181 10.6151
R7415 GND.n3631 GND.n2181 10.6151
R7416 GND.n3631 GND.n2198 10.6151
R7417 GND.n4528 GND.n2198 10.6151
R7418 GND.n4528 GND.n4527 10.6151
R7419 GND.n4527 GND.n4526 10.6151
R7420 GND.n4526 GND.n2199 10.6151
R7421 GND.n3128 GND.n2199 10.6151
R7422 GND.n3674 GND.n3128 10.6151
R7423 GND.n3675 GND.n3674 10.6151
R7424 GND.n3676 GND.n3675 10.6151
R7425 GND.n3676 GND.n2228 10.6151
R7426 GND.n4507 GND.n2228 10.6151
R7427 GND.n4507 GND.n4506 10.6151
R7428 GND.n4506 GND.n4505 10.6151
R7429 GND.n4505 GND.n2229 10.6151
R7430 GND.n2254 GND.n2229 10.6151
R7431 GND.n4494 GND.n2254 10.6151
R7432 GND.n4494 GND.n4493 10.6151
R7433 GND.n4493 GND.n4492 10.6151
R7434 GND.n4492 GND.n2255 10.6151
R7435 GND.n3717 GND.n2255 10.6151
R7436 GND.n3717 GND.n3716 10.6151
R7437 GND.n3716 GND.n3715 10.6151
R7438 GND.n3715 GND.n3712 10.6151
R7439 GND.n3712 GND.n2297 10.6151
R7440 GND.n4473 GND.n2297 10.6151
R7441 GND.n4473 GND.n4472 10.6151
R7442 GND.n4472 GND.n4471 10.6151
R7443 GND.n4471 GND.n2298 10.6151
R7444 GND.n2321 GND.n2298 10.6151
R7445 GND.n4459 GND.n2321 10.6151
R7446 GND.n4459 GND.n4458 10.6151
R7447 GND.n4458 GND.n4457 10.6151
R7448 GND.n4457 GND.n2322 10.6151
R7449 GND.n3778 GND.n2322 10.6151
R7450 GND.n3778 GND.n3777 10.6151
R7451 GND.n3777 GND.n3776 10.6151
R7452 GND.n3776 GND.n3771 10.6151
R7453 GND.n3771 GND.n2364 10.6151
R7454 GND.n4438 GND.n2364 10.6151
R7455 GND.n4438 GND.n4437 10.6151
R7456 GND.n4437 GND.n4436 10.6151
R7457 GND.n4436 GND.n2365 10.6151
R7458 GND.n3033 GND.n2365 10.6151
R7459 GND.n4003 GND.n3033 10.6151
R7460 GND.n1454 GND.n1436 10.4732
R7461 GND.n1232 GND.n1214 10.4732
R7462 GND.n2490 GND.n2472 10.4732
R7463 GND.n2455 GND.n2437 10.4732
R7464 GND.n4651 GND.n1478 10.3534
R7465 GND.n3186 GND.n3185 10.3534
R7466 GND.n3527 GND.n2126 10.3534
R7467 GND.n3630 GND.n2192 10.3534
R7468 GND.n3671 GND.n3670 10.3534
R7469 GND.n3740 GND.n3739 10.3534
R7470 GND.n3727 GND.n2324 10.3534
R7471 GND.n4425 GND.n2395 10.3534
R7472 GND.n1443 GND.n1442 10.2746
R7473 GND.n1221 GND.n1220 10.2746
R7474 GND.n2479 GND.n2478 10.2746
R7475 GND.n2444 GND.n2443 10.2746
R7476 GND.n3331 GND.n3330 10.2247
R7477 GND.n3041 GND.n3040 10.2247
R7478 GND.n1453 GND.n1438 9.69747
R7479 GND.n1231 GND.n1216 9.69747
R7480 GND.n2489 GND.n2474 9.69747
R7481 GND.n2454 GND.n2439 9.69747
R7482 GND.n4565 GND.n2146 9.66325
R7483 GND.n4545 GND.n2174 9.66325
R7484 GND.n3684 GND.n2225 9.66325
R7485 GND.n3719 GND.n3710 9.66325
R7486 GND.n3042 GND.n3034 9.50353
R7487 GND.n57 GND.n56 9.45567
R7488 GND.n68 GND.n67 9.45567
R7489 GND.n33 GND.n32 9.45567
R7490 GND.n44 GND.n43 9.45567
R7491 GND.n10 GND.n9 9.45567
R7492 GND.n21 GND.n20 9.45567
R7493 GND.n1460 GND.n1432 9.45567
R7494 GND.n1238 GND.n1210 9.45567
R7495 GND.n140 GND.n139 9.45567
R7496 GND.n129 GND.n128 9.45567
R7497 GND.n116 GND.n115 9.45567
R7498 GND.n105 GND.n104 9.45567
R7499 GND.n93 GND.n92 9.45567
R7500 GND.n82 GND.n81 9.45567
R7501 GND.n2496 GND.n2468 9.45567
R7502 GND.n2461 GND.n2433 9.45567
R7503 GND.n3938 GND.n3071 9.36635
R7504 GND.n3405 GND.n3303 9.36635
R7505 GND.n3311 GND.n3310 9.36635
R7506 GND.n3959 GND.n3958 9.36635
R7507 GND.n3606 GND.t32 9.31815
R7508 GND.t4 GND.n2214 9.31815
R7509 GND.n56 GND.n55 9.3005
R7510 GND.n49 GND.n48 9.3005
R7511 GND.n67 GND.n66 9.3005
R7512 GND.n60 GND.n59 9.3005
R7513 GND.n32 GND.n31 9.3005
R7514 GND.n25 GND.n24 9.3005
R7515 GND.n43 GND.n42 9.3005
R7516 GND.n36 GND.n35 9.3005
R7517 GND.n9 GND.n8 9.3005
R7518 GND.n2 GND.n1 9.3005
R7519 GND.n20 GND.n19 9.3005
R7520 GND.n13 GND.n12 9.3005
R7521 GND.n1440 GND.n1439 9.3005
R7522 GND.n1451 GND.n1450 9.3005
R7523 GND.n1453 GND.n1452 9.3005
R7524 GND.n1436 GND.n1435 9.3005
R7525 GND.n1459 GND.n1458 9.3005
R7526 GND.n1461 GND.n1460 9.3005
R7527 GND.n1445 GND.n1444 9.3005
R7528 GND.n1223 GND.n1222 9.3005
R7529 GND.n1218 GND.n1217 9.3005
R7530 GND.n1229 GND.n1228 9.3005
R7531 GND.n1231 GND.n1230 9.3005
R7532 GND.n1214 GND.n1213 9.3005
R7533 GND.n1237 GND.n1236 9.3005
R7534 GND.n1239 GND.n1238 9.3005
R7535 GND.n4975 GND.n4974 9.3005
R7536 GND.n4976 GND.n797 9.3005
R7537 GND.n4978 GND.n4977 9.3005
R7538 GND.n793 GND.n792 9.3005
R7539 GND.n4985 GND.n4984 9.3005
R7540 GND.n4986 GND.n791 9.3005
R7541 GND.n4988 GND.n4987 9.3005
R7542 GND.n787 GND.n786 9.3005
R7543 GND.n4995 GND.n4994 9.3005
R7544 GND.n4996 GND.n785 9.3005
R7545 GND.n4998 GND.n4997 9.3005
R7546 GND.n781 GND.n780 9.3005
R7547 GND.n5005 GND.n5004 9.3005
R7548 GND.n5006 GND.n779 9.3005
R7549 GND.n5008 GND.n5007 9.3005
R7550 GND.n775 GND.n774 9.3005
R7551 GND.n5015 GND.n5014 9.3005
R7552 GND.n5016 GND.n773 9.3005
R7553 GND.n5018 GND.n5017 9.3005
R7554 GND.n769 GND.n768 9.3005
R7555 GND.n5025 GND.n5024 9.3005
R7556 GND.n5026 GND.n767 9.3005
R7557 GND.n5028 GND.n5027 9.3005
R7558 GND.n763 GND.n762 9.3005
R7559 GND.n5035 GND.n5034 9.3005
R7560 GND.n5036 GND.n761 9.3005
R7561 GND.n5038 GND.n5037 9.3005
R7562 GND.n757 GND.n756 9.3005
R7563 GND.n5045 GND.n5044 9.3005
R7564 GND.n5046 GND.n755 9.3005
R7565 GND.n5048 GND.n5047 9.3005
R7566 GND.n751 GND.n750 9.3005
R7567 GND.n5055 GND.n5054 9.3005
R7568 GND.n5056 GND.n749 9.3005
R7569 GND.n5058 GND.n5057 9.3005
R7570 GND.n745 GND.n744 9.3005
R7571 GND.n5065 GND.n5064 9.3005
R7572 GND.n5066 GND.n743 9.3005
R7573 GND.n5068 GND.n5067 9.3005
R7574 GND.n739 GND.n738 9.3005
R7575 GND.n5075 GND.n5074 9.3005
R7576 GND.n5076 GND.n737 9.3005
R7577 GND.n5078 GND.n5077 9.3005
R7578 GND.n733 GND.n732 9.3005
R7579 GND.n5085 GND.n5084 9.3005
R7580 GND.n5086 GND.n731 9.3005
R7581 GND.n5088 GND.n5087 9.3005
R7582 GND.n727 GND.n726 9.3005
R7583 GND.n5095 GND.n5094 9.3005
R7584 GND.n5096 GND.n725 9.3005
R7585 GND.n5098 GND.n5097 9.3005
R7586 GND.n721 GND.n720 9.3005
R7587 GND.n5105 GND.n5104 9.3005
R7588 GND.n5106 GND.n719 9.3005
R7589 GND.n5108 GND.n5107 9.3005
R7590 GND.n715 GND.n714 9.3005
R7591 GND.n5115 GND.n5114 9.3005
R7592 GND.n5116 GND.n713 9.3005
R7593 GND.n5118 GND.n5117 9.3005
R7594 GND.n709 GND.n708 9.3005
R7595 GND.n5125 GND.n5124 9.3005
R7596 GND.n5126 GND.n707 9.3005
R7597 GND.n5128 GND.n5127 9.3005
R7598 GND.n703 GND.n702 9.3005
R7599 GND.n5135 GND.n5134 9.3005
R7600 GND.n5136 GND.n701 9.3005
R7601 GND.n5138 GND.n5137 9.3005
R7602 GND.n697 GND.n696 9.3005
R7603 GND.n5145 GND.n5144 9.3005
R7604 GND.n5146 GND.n695 9.3005
R7605 GND.n5148 GND.n5147 9.3005
R7606 GND.n691 GND.n690 9.3005
R7607 GND.n5155 GND.n5154 9.3005
R7608 GND.n5156 GND.n689 9.3005
R7609 GND.n5158 GND.n5157 9.3005
R7610 GND.n685 GND.n684 9.3005
R7611 GND.n5165 GND.n5164 9.3005
R7612 GND.n5166 GND.n683 9.3005
R7613 GND.n5168 GND.n5167 9.3005
R7614 GND.n679 GND.n678 9.3005
R7615 GND.n5175 GND.n5174 9.3005
R7616 GND.n5176 GND.n677 9.3005
R7617 GND.n5178 GND.n5177 9.3005
R7618 GND.n673 GND.n672 9.3005
R7619 GND.n5185 GND.n5184 9.3005
R7620 GND.n5186 GND.n671 9.3005
R7621 GND.n5188 GND.n5187 9.3005
R7622 GND.n667 GND.n666 9.3005
R7623 GND.n5195 GND.n5194 9.3005
R7624 GND.n5196 GND.n665 9.3005
R7625 GND.n5198 GND.n5197 9.3005
R7626 GND.n661 GND.n660 9.3005
R7627 GND.n5205 GND.n5204 9.3005
R7628 GND.n5206 GND.n659 9.3005
R7629 GND.n5208 GND.n5207 9.3005
R7630 GND.n655 GND.n654 9.3005
R7631 GND.n5215 GND.n5214 9.3005
R7632 GND.n5216 GND.n653 9.3005
R7633 GND.n5218 GND.n5217 9.3005
R7634 GND.n649 GND.n648 9.3005
R7635 GND.n5225 GND.n5224 9.3005
R7636 GND.n5226 GND.n647 9.3005
R7637 GND.n5228 GND.n5227 9.3005
R7638 GND.n643 GND.n642 9.3005
R7639 GND.n5235 GND.n5234 9.3005
R7640 GND.n5236 GND.n641 9.3005
R7641 GND.n5238 GND.n5237 9.3005
R7642 GND.n637 GND.n636 9.3005
R7643 GND.n5245 GND.n5244 9.3005
R7644 GND.n5246 GND.n635 9.3005
R7645 GND.n5248 GND.n5247 9.3005
R7646 GND.n631 GND.n630 9.3005
R7647 GND.n5255 GND.n5254 9.3005
R7648 GND.n5256 GND.n629 9.3005
R7649 GND.n5258 GND.n5257 9.3005
R7650 GND.n625 GND.n624 9.3005
R7651 GND.n5265 GND.n5264 9.3005
R7652 GND.n5266 GND.n623 9.3005
R7653 GND.n5268 GND.n5267 9.3005
R7654 GND.n619 GND.n618 9.3005
R7655 GND.n5275 GND.n5274 9.3005
R7656 GND.n5276 GND.n617 9.3005
R7657 GND.n5278 GND.n5277 9.3005
R7658 GND.n613 GND.n612 9.3005
R7659 GND.n5285 GND.n5284 9.3005
R7660 GND.n5286 GND.n611 9.3005
R7661 GND.n5288 GND.n5287 9.3005
R7662 GND.n607 GND.n606 9.3005
R7663 GND.n5295 GND.n5294 9.3005
R7664 GND.n5296 GND.n605 9.3005
R7665 GND.n5298 GND.n5297 9.3005
R7666 GND.n601 GND.n600 9.3005
R7667 GND.n5305 GND.n5304 9.3005
R7668 GND.n5306 GND.n599 9.3005
R7669 GND.n5308 GND.n5307 9.3005
R7670 GND.n595 GND.n594 9.3005
R7671 GND.n5315 GND.n5314 9.3005
R7672 GND.n5316 GND.n593 9.3005
R7673 GND.n5318 GND.n5317 9.3005
R7674 GND.n589 GND.n588 9.3005
R7675 GND.n5325 GND.n5324 9.3005
R7676 GND.n5326 GND.n587 9.3005
R7677 GND.n5328 GND.n5327 9.3005
R7678 GND.n583 GND.n582 9.3005
R7679 GND.n5335 GND.n5334 9.3005
R7680 GND.n5336 GND.n581 9.3005
R7681 GND.n5338 GND.n5337 9.3005
R7682 GND.n577 GND.n576 9.3005
R7683 GND.n5345 GND.n5344 9.3005
R7684 GND.n5346 GND.n575 9.3005
R7685 GND.n5348 GND.n5347 9.3005
R7686 GND.n571 GND.n570 9.3005
R7687 GND.n5355 GND.n5354 9.3005
R7688 GND.n5356 GND.n569 9.3005
R7689 GND.n5358 GND.n5357 9.3005
R7690 GND.n565 GND.n564 9.3005
R7691 GND.n5365 GND.n5364 9.3005
R7692 GND.n5366 GND.n563 9.3005
R7693 GND.n5368 GND.n5367 9.3005
R7694 GND.n559 GND.n558 9.3005
R7695 GND.n5375 GND.n5374 9.3005
R7696 GND.n5376 GND.n557 9.3005
R7697 GND.n5378 GND.n5377 9.3005
R7698 GND.n553 GND.n552 9.3005
R7699 GND.n5385 GND.n5384 9.3005
R7700 GND.n5386 GND.n551 9.3005
R7701 GND.n5388 GND.n5387 9.3005
R7702 GND.n547 GND.n546 9.3005
R7703 GND.n5395 GND.n5394 9.3005
R7704 GND.n5396 GND.n545 9.3005
R7705 GND.n5398 GND.n5397 9.3005
R7706 GND.n541 GND.n540 9.3005
R7707 GND.n5405 GND.n5404 9.3005
R7708 GND.n5406 GND.n539 9.3005
R7709 GND.n5408 GND.n5407 9.3005
R7710 GND.n535 GND.n534 9.3005
R7711 GND.n5415 GND.n5414 9.3005
R7712 GND.n5416 GND.n533 9.3005
R7713 GND.n5418 GND.n5417 9.3005
R7714 GND.n529 GND.n528 9.3005
R7715 GND.n5425 GND.n5424 9.3005
R7716 GND.n5426 GND.n527 9.3005
R7717 GND.n5428 GND.n5427 9.3005
R7718 GND.n523 GND.n522 9.3005
R7719 GND.n5435 GND.n5434 9.3005
R7720 GND.n5436 GND.n521 9.3005
R7721 GND.n5438 GND.n5437 9.3005
R7722 GND.n517 GND.n516 9.3005
R7723 GND.n5445 GND.n5444 9.3005
R7724 GND.n5446 GND.n515 9.3005
R7725 GND.n5448 GND.n5447 9.3005
R7726 GND.n511 GND.n510 9.3005
R7727 GND.n5455 GND.n5454 9.3005
R7728 GND.n5456 GND.n509 9.3005
R7729 GND.n5458 GND.n5457 9.3005
R7730 GND.n505 GND.n504 9.3005
R7731 GND.n5465 GND.n5464 9.3005
R7732 GND.n5466 GND.n503 9.3005
R7733 GND.n5468 GND.n5467 9.3005
R7734 GND.n499 GND.n498 9.3005
R7735 GND.n5475 GND.n5474 9.3005
R7736 GND.n5476 GND.n497 9.3005
R7737 GND.n5478 GND.n5477 9.3005
R7738 GND.n493 GND.n492 9.3005
R7739 GND.n5485 GND.n5484 9.3005
R7740 GND.n5486 GND.n491 9.3005
R7741 GND.n5488 GND.n5487 9.3005
R7742 GND.n487 GND.n486 9.3005
R7743 GND.n5495 GND.n5494 9.3005
R7744 GND.n5496 GND.n485 9.3005
R7745 GND.n5498 GND.n5497 9.3005
R7746 GND.n481 GND.n480 9.3005
R7747 GND.n5505 GND.n5504 9.3005
R7748 GND.n5506 GND.n479 9.3005
R7749 GND.n5508 GND.n5507 9.3005
R7750 GND.n475 GND.n474 9.3005
R7751 GND.n5515 GND.n5514 9.3005
R7752 GND.n5516 GND.n473 9.3005
R7753 GND.n5518 GND.n5517 9.3005
R7754 GND.n469 GND.n468 9.3005
R7755 GND.n5525 GND.n5524 9.3005
R7756 GND.n5526 GND.n467 9.3005
R7757 GND.n5528 GND.n5527 9.3005
R7758 GND.n463 GND.n462 9.3005
R7759 GND.n5535 GND.n5534 9.3005
R7760 GND.n5536 GND.n461 9.3005
R7761 GND.n5538 GND.n5537 9.3005
R7762 GND.n457 GND.n456 9.3005
R7763 GND.n5545 GND.n5544 9.3005
R7764 GND.n5548 GND.n5547 9.3005
R7765 GND.n451 GND.n450 9.3005
R7766 GND.n5555 GND.n5554 9.3005
R7767 GND.n5556 GND.n449 9.3005
R7768 GND.n5558 GND.n5557 9.3005
R7769 GND.n445 GND.n444 9.3005
R7770 GND.n5565 GND.n5564 9.3005
R7771 GND.n5566 GND.n443 9.3005
R7772 GND.n5568 GND.n5567 9.3005
R7773 GND.n439 GND.n438 9.3005
R7774 GND.n5575 GND.n5574 9.3005
R7775 GND.n5576 GND.n437 9.3005
R7776 GND.n5578 GND.n5577 9.3005
R7777 GND.n433 GND.n432 9.3005
R7778 GND.n5585 GND.n5584 9.3005
R7779 GND.n5586 GND.n431 9.3005
R7780 GND.n5588 GND.n5587 9.3005
R7781 GND.n427 GND.n426 9.3005
R7782 GND.n5595 GND.n5594 9.3005
R7783 GND.n5596 GND.n425 9.3005
R7784 GND.n5598 GND.n5597 9.3005
R7785 GND.n421 GND.n420 9.3005
R7786 GND.n5605 GND.n5604 9.3005
R7787 GND.n5606 GND.n419 9.3005
R7788 GND.n5608 GND.n5607 9.3005
R7789 GND.n415 GND.n414 9.3005
R7790 GND.n5615 GND.n5614 9.3005
R7791 GND.n5616 GND.n413 9.3005
R7792 GND.n5618 GND.n5617 9.3005
R7793 GND.n409 GND.n408 9.3005
R7794 GND.n5625 GND.n5624 9.3005
R7795 GND.n5626 GND.n407 9.3005
R7796 GND.n5628 GND.n5627 9.3005
R7797 GND.n403 GND.n402 9.3005
R7798 GND.n5635 GND.n5634 9.3005
R7799 GND.n5636 GND.n401 9.3005
R7800 GND.n5638 GND.n5637 9.3005
R7801 GND.n397 GND.n396 9.3005
R7802 GND.n5645 GND.n5644 9.3005
R7803 GND.n5646 GND.n395 9.3005
R7804 GND.n5648 GND.n5647 9.3005
R7805 GND.n391 GND.n390 9.3005
R7806 GND.n5655 GND.n5654 9.3005
R7807 GND.n5656 GND.n389 9.3005
R7808 GND.n5658 GND.n5657 9.3005
R7809 GND.n385 GND.n384 9.3005
R7810 GND.n5665 GND.n5664 9.3005
R7811 GND.n5666 GND.n383 9.3005
R7812 GND.n5668 GND.n5667 9.3005
R7813 GND.n379 GND.n378 9.3005
R7814 GND.n5675 GND.n5674 9.3005
R7815 GND.n5676 GND.n377 9.3005
R7816 GND.n5680 GND.n5677 9.3005
R7817 GND.n5679 GND.n5678 9.3005
R7818 GND.n5546 GND.n455 9.3005
R7819 GND.n139 GND.n138 9.3005
R7820 GND.n132 GND.n131 9.3005
R7821 GND.n128 GND.n127 9.3005
R7822 GND.n121 GND.n120 9.3005
R7823 GND.n115 GND.n114 9.3005
R7824 GND.n108 GND.n107 9.3005
R7825 GND.n104 GND.n103 9.3005
R7826 GND.n97 GND.n96 9.3005
R7827 GND.n92 GND.n91 9.3005
R7828 GND.n85 GND.n84 9.3005
R7829 GND.n81 GND.n80 9.3005
R7830 GND.n74 GND.n73 9.3005
R7831 GND.n2476 GND.n2475 9.3005
R7832 GND.n2487 GND.n2486 9.3005
R7833 GND.n2489 GND.n2488 9.3005
R7834 GND.n2472 GND.n2471 9.3005
R7835 GND.n2495 GND.n2494 9.3005
R7836 GND.n2497 GND.n2496 9.3005
R7837 GND.n2481 GND.n2480 9.3005
R7838 GND.n2446 GND.n2445 9.3005
R7839 GND.n2441 GND.n2440 9.3005
R7840 GND.n2452 GND.n2451 9.3005
R7841 GND.n2454 GND.n2453 9.3005
R7842 GND.n2437 GND.n2436 9.3005
R7843 GND.n2460 GND.n2459 9.3005
R7844 GND.n2462 GND.n2461 9.3005
R7845 GND.n4614 GND.n4613 9.3005
R7846 GND.n4612 GND.n2076 9.3005
R7847 GND.n4611 GND.n4610 9.3005
R7848 GND.n2078 GND.n2077 9.3005
R7849 GND.n2107 GND.n2106 9.3005
R7850 GND.n2108 GND.n2104 9.3005
R7851 GND.n4591 GND.n2109 9.3005
R7852 GND.n4590 GND.n2110 9.3005
R7853 GND.n4589 GND.n2111 9.3005
R7854 GND.n2128 GND.n2112 9.3005
R7855 GND.n4577 GND.n2129 9.3005
R7856 GND.n4576 GND.n2130 9.3005
R7857 GND.n4575 GND.n2131 9.3005
R7858 GND.n2148 GND.n2132 9.3005
R7859 GND.n4563 GND.n2149 9.3005
R7860 GND.n4562 GND.n2150 9.3005
R7861 GND.n4561 GND.n2151 9.3005
R7862 GND.n2168 GND.n2152 9.3005
R7863 GND.n4549 GND.n2169 9.3005
R7864 GND.n4548 GND.n2170 9.3005
R7865 GND.n4547 GND.n2171 9.3005
R7866 GND.n2186 GND.n2172 9.3005
R7867 GND.n4535 GND.n2187 9.3005
R7868 GND.n4534 GND.n2188 9.3005
R7869 GND.n4533 GND.n2189 9.3005
R7870 GND.n2206 GND.n2190 9.3005
R7871 GND.n4521 GND.n2207 9.3005
R7872 GND.n4520 GND.n2208 9.3005
R7873 GND.n4519 GND.n2209 9.3005
R7874 GND.n2238 GND.n2210 9.3005
R7875 GND.n2241 GND.n2240 9.3005
R7876 GND.n2242 GND.n2237 9.3005
R7877 GND.n4500 GND.n2243 9.3005
R7878 GND.n4499 GND.n2244 9.3005
R7879 GND.n4498 GND.n2245 9.3005
R7880 GND.n2282 GND.n2246 9.3005
R7881 GND.n2285 GND.n2284 9.3005
R7882 GND.n2286 GND.n2281 9.3005
R7883 GND.n4480 GND.n2287 9.3005
R7884 GND.n4479 GND.n2288 9.3005
R7885 GND.n4478 GND.n2289 9.3005
R7886 GND.n2331 GND.n2290 9.3005
R7887 GND.n2333 GND.n2332 9.3005
R7888 GND.n2337 GND.n2336 9.3005
R7889 GND.n2338 GND.n2330 9.3005
R7890 GND.n4452 GND.n2339 9.3005
R7891 GND.n4451 GND.n2340 9.3005
R7892 GND.n4450 GND.n2341 9.3005
R7893 GND.n3794 GND.n2342 9.3005
R7894 GND.n3797 GND.n3796 9.3005
R7895 GND.n3795 GND.n2372 9.3005
R7896 GND.n4432 GND.n2373 9.3005
R7897 GND.n4431 GND.n4430 9.3005
R7898 GND.n2075 GND.n1474 9.3005
R7899 GND.n3236 GND.n3235 9.3005
R7900 GND.n3238 GND.n3234 9.3005
R7901 GND.n3239 GND.n3233 9.3005
R7902 GND.n3242 GND.n3229 9.3005
R7903 GND.n3243 GND.n3228 9.3005
R7904 GND.n3246 GND.n3227 9.3005
R7905 GND.n3247 GND.n3226 9.3005
R7906 GND.n3250 GND.n3225 9.3005
R7907 GND.n3251 GND.n3224 9.3005
R7908 GND.n3254 GND.n3223 9.3005
R7909 GND.n3255 GND.n3222 9.3005
R7910 GND.n3258 GND.n3221 9.3005
R7911 GND.n3259 GND.n3220 9.3005
R7912 GND.n3262 GND.n3219 9.3005
R7913 GND.n3263 GND.n3218 9.3005
R7914 GND.n3266 GND.n3217 9.3005
R7915 GND.n3267 GND.n3216 9.3005
R7916 GND.n3270 GND.n3215 9.3005
R7917 GND.n3272 GND.n3214 9.3005
R7918 GND.n3273 GND.n3213 9.3005
R7919 GND.n3274 GND.n3212 9.3005
R7920 GND.n3275 GND.n1475 9.3005
R7921 GND.n3198 GND.n3197 9.3005
R7922 GND.n3284 GND.n3196 9.3005
R7923 GND.n3480 GND.n3285 9.3005
R7924 GND.n3481 GND.n3195 9.3005
R7925 GND.n3484 GND.n3483 9.3005
R7926 GND.n3485 GND.n3194 9.3005
R7927 GND.n3487 GND.n3486 9.3005
R7928 GND.n3184 GND.n3183 9.3005
R7929 GND.n3510 GND.n3509 9.3005
R7930 GND.n3511 GND.n3182 9.3005
R7931 GND.n3513 GND.n3512 9.3005
R7932 GND.n3178 GND.n3177 9.3005
R7933 GND.n3557 GND.n3556 9.3005
R7934 GND.n3558 GND.n3176 9.3005
R7935 GND.n3561 GND.n3560 9.3005
R7936 GND.n3559 GND.n3160 9.3005
R7937 GND.n3582 GND.n3161 9.3005
R7938 GND.n3581 GND.n3162 9.3005
R7939 GND.n3580 GND.n3163 9.3005
R7940 GND.n3173 GND.n3164 9.3005
R7941 GND.n3172 GND.n3165 9.3005
R7942 GND.n3170 GND.n3166 9.3005
R7943 GND.n3169 GND.n3167 9.3005
R7944 GND.n3136 GND.n3135 9.3005
R7945 GND.n3637 GND.n3636 9.3005
R7946 GND.n3638 GND.n3134 9.3005
R7947 GND.n3657 GND.n3639 9.3005
R7948 GND.n3656 GND.n3640 9.3005
R7949 GND.n3655 GND.n3641 9.3005
R7950 GND.n3653 GND.n3642 9.3005
R7951 GND.n3652 GND.n3643 9.3005
R7952 GND.n3645 GND.n3644 9.3005
R7953 GND.n3648 GND.n3647 9.3005
R7954 GND.n3646 GND.n3120 9.3005
R7955 GND.n3700 GND.n3121 9.3005
R7956 GND.n3701 GND.n3119 9.3005
R7957 GND.n3704 GND.n3703 9.3005
R7958 GND.n3705 GND.n3118 9.3005
R7959 GND.n3708 GND.n3707 9.3005
R7960 GND.n3706 GND.n3108 9.3005
R7961 GND.n3749 GND.n3107 9.3005
R7962 GND.n3751 GND.n3750 9.3005
R7963 GND.n3752 GND.n3106 9.3005
R7964 GND.n3754 GND.n3753 9.3005
R7965 GND.n3104 GND.n3103 9.3005
R7966 GND.n3759 GND.n3758 9.3005
R7967 GND.n3760 GND.n3102 9.3005
R7968 GND.n3766 GND.n3761 9.3005
R7969 GND.n3765 GND.n3762 9.3005
R7970 GND.n3764 GND.n3763 9.3005
R7971 GND.n3094 GND.n3093 9.3005
R7972 GND.n3803 GND.n3802 9.3005
R7973 GND.n3804 GND.n3092 9.3005
R7974 GND.n3888 GND.n3887 9.3005
R7975 GND.n3283 GND.n3282 9.3005
R7976 GND.n3878 GND.n3877 9.3005
R7977 GND.n3876 GND.n3819 9.3005
R7978 GND.n3875 GND.n3874 9.3005
R7979 GND.n3871 GND.n3820 9.3005
R7980 GND.n3868 GND.n3821 9.3005
R7981 GND.n3867 GND.n3822 9.3005
R7982 GND.n3864 GND.n3823 9.3005
R7983 GND.n3863 GND.n3824 9.3005
R7984 GND.n3860 GND.n3825 9.3005
R7985 GND.n3859 GND.n3826 9.3005
R7986 GND.n3856 GND.n3827 9.3005
R7987 GND.n3855 GND.n3828 9.3005
R7988 GND.n3852 GND.n3829 9.3005
R7989 GND.n3851 GND.n3830 9.3005
R7990 GND.n3848 GND.n3831 9.3005
R7991 GND.n3847 GND.n3832 9.3005
R7992 GND.n3844 GND.n3833 9.3005
R7993 GND.n3843 GND.n3834 9.3005
R7994 GND.n3840 GND.n3839 9.3005
R7995 GND.n3838 GND.n3806 9.3005
R7996 GND.n3884 GND.n3805 9.3005
R7997 GND.n3886 GND.n3885 9.3005
R7998 GND.n3879 GND.n2374 9.3005
R7999 GND.n2789 GND.n2788 9.3005
R8000 GND.n2792 GND.n2787 9.3005
R8001 GND.n2793 GND.n2432 9.3005
R8002 GND.n2796 GND.n2431 9.3005
R8003 GND.n2797 GND.n2430 9.3005
R8004 GND.n2800 GND.n2429 9.3005
R8005 GND.n2801 GND.n2428 9.3005
R8006 GND.n2379 GND.n2375 9.3005
R8007 GND.n4428 GND.n4427 9.3005
R8008 GND.n2997 GND.n2996 9.3005
R8009 GND.n2998 GND.n2992 9.3005
R8010 GND.n3002 GND.n3001 9.3005
R8011 GND.n3003 GND.n2991 9.3005
R8012 GND.n3005 GND.n3004 9.3005
R8013 GND.n2989 GND.n2988 9.3005
R8014 GND.n4088 GND.n4087 9.3005
R8015 GND.n4089 GND.n2987 9.3005
R8016 GND.n4091 GND.n4090 9.3005
R8017 GND.n2985 GND.n2984 9.3005
R8018 GND.n4103 GND.n4102 9.3005
R8019 GND.n4104 GND.n2983 9.3005
R8020 GND.n4106 GND.n4105 9.3005
R8021 GND.n2981 GND.n2980 9.3005
R8022 GND.n4118 GND.n4117 9.3005
R8023 GND.n4119 GND.n2979 9.3005
R8024 GND.n4133 GND.n4120 9.3005
R8025 GND.n4132 GND.n4121 9.3005
R8026 GND.n4131 GND.n4122 9.3005
R8027 GND.n4130 GND.n4123 9.3005
R8028 GND.n4127 GND.n4124 9.3005
R8029 GND.n4126 GND.n4125 9.3005
R8030 GND.n145 GND.n143 9.3005
R8031 GND.n2993 GND.n2376 9.3005
R8032 GND.n5862 GND.n5861 9.3005
R8033 GND.n146 GND.n144 9.3005
R8034 GND.n4161 GND.n4160 9.3005
R8035 GND.n4163 GND.n4162 9.3005
R8036 GND.n2976 GND.n2975 9.3005
R8037 GND.n4174 GND.n4173 9.3005
R8038 GND.n4175 GND.n2974 9.3005
R8039 GND.n4177 GND.n4176 9.3005
R8040 GND.n2971 GND.n2970 9.3005
R8041 GND.n4188 GND.n4187 9.3005
R8042 GND.n4189 GND.n2969 9.3005
R8043 GND.n4191 GND.n4190 9.3005
R8044 GND.n2966 GND.n2965 9.3005
R8045 GND.n4202 GND.n4201 9.3005
R8046 GND.n4203 GND.n2964 9.3005
R8047 GND.n4206 GND.n4205 9.3005
R8048 GND.n4204 GND.n2957 9.3005
R8049 GND.n4260 GND.n2958 9.3005
R8050 GND.n4259 GND.n2959 9.3005
R8051 GND.n4258 GND.n2960 9.3005
R8052 GND.n4215 GND.n2961 9.3005
R8053 GND.n4248 GND.n4216 9.3005
R8054 GND.n4247 GND.n4217 9.3005
R8055 GND.n4246 GND.n4245 9.3005
R8056 GND.n4227 GND.n4226 9.3005
R8057 GND.n4229 GND.n4228 9.3005
R8058 GND.n4232 GND.n4223 9.3005
R8059 GND.n4236 GND.n4235 9.3005
R8060 GND.n4237 GND.n4222 9.3005
R8061 GND.n4240 GND.n4238 9.3005
R8062 GND.n4241 GND.n4218 9.3005
R8063 GND.n4244 GND.n4243 9.3005
R8064 GND.n4224 GND.n306 9.3005
R8065 GND.n270 GND.n269 9.3005
R8066 GND.n5787 GND.n288 9.3005
R8067 GND.n5786 GND.n289 9.3005
R8068 GND.n5785 GND.n290 9.3005
R8069 GND.n5782 GND.n291 9.3005
R8070 GND.n5781 GND.n292 9.3005
R8071 GND.n5778 GND.n293 9.3005
R8072 GND.n5774 GND.n294 9.3005
R8073 GND.n5771 GND.n295 9.3005
R8074 GND.n5770 GND.n296 9.3005
R8075 GND.n5767 GND.n297 9.3005
R8076 GND.n5766 GND.n298 9.3005
R8077 GND.n5763 GND.n299 9.3005
R8078 GND.n5762 GND.n300 9.3005
R8079 GND.n5759 GND.n301 9.3005
R8080 GND.n5758 GND.n302 9.3005
R8081 GND.n5755 GND.n5754 9.3005
R8082 GND.n5753 GND.n303 9.3005
R8083 GND.n5793 GND.n5792 9.3005
R8084 GND.n4386 GND.n4385 9.3005
R8085 GND.n2806 GND.n2805 9.3005
R8086 GND.n2831 GND.n2830 9.3005
R8087 GND.n4373 GND.n2832 9.3005
R8088 GND.n4372 GND.n2833 9.3005
R8089 GND.n4371 GND.n2834 9.3005
R8090 GND.n4082 GND.n2835 9.3005
R8091 GND.n4361 GND.n2852 9.3005
R8092 GND.n4360 GND.n2853 9.3005
R8093 GND.n4359 GND.n2854 9.3005
R8094 GND.n4097 GND.n2855 9.3005
R8095 GND.n4349 GND.n2873 9.3005
R8096 GND.n4348 GND.n2874 9.3005
R8097 GND.n4347 GND.n2875 9.3005
R8098 GND.n4112 GND.n2876 9.3005
R8099 GND.n4337 GND.n2895 9.3005
R8100 GND.n4336 GND.n2896 9.3005
R8101 GND.n4335 GND.n2897 9.3005
R8102 GND.n4140 GND.n2898 9.3005
R8103 GND.n4143 GND.n4142 9.3005
R8104 GND.n4144 GND.n2921 9.3005
R8105 GND.n4314 GND.n2922 9.3005
R8106 GND.n4313 GND.n2923 9.3005
R8107 GND.n4312 GND.n2924 9.3005
R8108 GND.n4311 GND.n2925 9.3005
R8109 GND.n4155 GND.n2926 9.3005
R8110 GND.n4156 GND.n174 9.3005
R8111 GND.n5850 GND.n175 9.3005
R8112 GND.n5849 GND.n176 9.3005
R8113 GND.n5848 GND.n177 9.3005
R8114 GND.n2973 GND.n178 9.3005
R8115 GND.n5838 GND.n195 9.3005
R8116 GND.n5837 GND.n196 9.3005
R8117 GND.n5836 GND.n197 9.3005
R8118 GND.n2968 GND.n198 9.3005
R8119 GND.n5826 GND.n216 9.3005
R8120 GND.n5825 GND.n217 9.3005
R8121 GND.n5824 GND.n218 9.3005
R8122 GND.n2963 GND.n219 9.3005
R8123 GND.n5814 GND.n237 9.3005
R8124 GND.n5813 GND.n238 9.3005
R8125 GND.n5812 GND.n239 9.3005
R8126 GND.n4214 GND.n240 9.3005
R8127 GND.n5802 GND.n257 9.3005
R8128 GND.n5801 GND.n258 9.3005
R8129 GND.n5800 GND.n259 9.3005
R8130 GND.n5751 GND.n260 9.3005
R8131 GND.n4387 GND.n2804 9.3005
R8132 GND.n4385 GND.n4384 9.3005
R8133 GND.n4383 GND.n2806 9.3005
R8134 GND.n2831 GND.n2807 9.3005
R8135 GND.n2990 GND.n2832 9.3005
R8136 GND.n4080 GND.n2833 9.3005
R8137 GND.n4081 GND.n2834 9.3005
R8138 GND.n4083 GND.n4082 9.3005
R8139 GND.n2986 GND.n2852 9.3005
R8140 GND.n4095 GND.n2853 9.3005
R8141 GND.n4096 GND.n2854 9.3005
R8142 GND.n4098 GND.n4097 9.3005
R8143 GND.n2982 GND.n2873 9.3005
R8144 GND.n4110 GND.n2874 9.3005
R8145 GND.n4111 GND.n2875 9.3005
R8146 GND.n4113 GND.n4112 9.3005
R8147 GND.n2978 GND.n2895 9.3005
R8148 GND.n4137 GND.n2896 9.3005
R8149 GND.n4138 GND.n2897 9.3005
R8150 GND.n4140 GND.n4139 9.3005
R8151 GND.n4143 GND.n2977 9.3005
R8152 GND.n4147 GND.n4144 9.3005
R8153 GND.n4148 GND.n2922 9.3005
R8154 GND.n4151 GND.n2923 9.3005
R8155 GND.n4152 GND.n2924 9.3005
R8156 GND.n4153 GND.n2925 9.3005
R8157 GND.n4155 GND.n4154 9.3005
R8158 GND.n4167 GND.n4156 9.3005
R8159 GND.n4168 GND.n175 9.3005
R8160 GND.n4169 GND.n176 9.3005
R8161 GND.n2972 GND.n177 9.3005
R8162 GND.n4181 GND.n2973 9.3005
R8163 GND.n4182 GND.n195 9.3005
R8164 GND.n4183 GND.n196 9.3005
R8165 GND.n2967 GND.n197 9.3005
R8166 GND.n4195 GND.n2968 9.3005
R8167 GND.n4196 GND.n216 9.3005
R8168 GND.n4197 GND.n217 9.3005
R8169 GND.n2962 GND.n218 9.3005
R8170 GND.n4210 GND.n2963 9.3005
R8171 GND.n4211 GND.n237 9.3005
R8172 GND.n4212 GND.n238 9.3005
R8173 GND.n4213 GND.n239 9.3005
R8174 GND.n4254 GND.n4214 9.3005
R8175 GND.n4253 GND.n257 9.3005
R8176 GND.n4252 GND.n258 9.3005
R8177 GND.n307 GND.n259 9.3005
R8178 GND.n5751 GND.n5750 9.3005
R8179 GND.n2804 GND.n2425 9.3005
R8180 GND.n4396 GND.n4395 9.3005
R8181 GND.n4397 GND.n2417 9.3005
R8182 GND.n4400 GND.n2416 9.3005
R8183 GND.n4401 GND.n2415 9.3005
R8184 GND.n4404 GND.n2414 9.3005
R8185 GND.n4405 GND.n2413 9.3005
R8186 GND.n4408 GND.n2412 9.3005
R8187 GND.n4409 GND.n2411 9.3005
R8188 GND.n4412 GND.n2410 9.3005
R8189 GND.n4414 GND.n2404 9.3005
R8190 GND.n4417 GND.n2403 9.3005
R8191 GND.n4419 GND.n2402 9.3005
R8192 GND.n4420 GND.n2401 9.3005
R8193 GND.n4421 GND.n2400 9.3005
R8194 GND.n4422 GND.n2399 9.3005
R8195 GND.n4394 GND.n2422 9.3005
R8196 GND.n4393 GND.n4392 9.3005
R8197 GND.n2818 GND.n2815 9.3005
R8198 GND.n4379 GND.n2819 9.3005
R8199 GND.n4378 GND.n2820 9.3005
R8200 GND.n4377 GND.n2821 9.3005
R8201 GND.n2841 GND.n2822 9.3005
R8202 GND.n4367 GND.n2842 9.3005
R8203 GND.n4366 GND.n2843 9.3005
R8204 GND.n4365 GND.n2844 9.3005
R8205 GND.n2862 GND.n2845 9.3005
R8206 GND.n4355 GND.n2863 9.3005
R8207 GND.n4354 GND.n2864 9.3005
R8208 GND.n4353 GND.n2865 9.3005
R8209 GND.n2883 GND.n2866 9.3005
R8210 GND.n4343 GND.n2884 9.3005
R8211 GND.n4342 GND.n2885 9.3005
R8212 GND.n4341 GND.n2886 9.3005
R8213 GND.n2888 GND.n2887 9.3005
R8214 GND.n4331 GND.n158 9.3005
R8215 GND.n165 GND.n157 9.3005
R8216 GND.n5844 GND.n185 9.3005
R8217 GND.n5843 GND.n186 9.3005
R8218 GND.n5842 GND.n187 9.3005
R8219 GND.n205 GND.n188 9.3005
R8220 GND.n5832 GND.n206 9.3005
R8221 GND.n5831 GND.n207 9.3005
R8222 GND.n5830 GND.n208 9.3005
R8223 GND.n226 GND.n209 9.3005
R8224 GND.n5820 GND.n227 9.3005
R8225 GND.n5819 GND.n228 9.3005
R8226 GND.n5818 GND.n229 9.3005
R8227 GND.n246 GND.n230 9.3005
R8228 GND.n5808 GND.n247 9.3005
R8229 GND.n5807 GND.n248 9.3005
R8230 GND.n5806 GND.n249 9.3005
R8231 GND.n267 GND.n250 9.3005
R8232 GND.n5796 GND.n268 9.3005
R8233 GND.n5795 GND.n5794 9.3005
R8234 GND.n2817 GND.n2816 9.3005
R8235 GND.n5855 GND.n162 9.3005
R8236 GND.n5855 GND.n5854 9.3005
R8237 GND.n1618 GND.n1616 9.3005
R8238 GND.n1664 GND.n1619 9.3005
R8239 GND.n1663 GND.n1620 9.3005
R8240 GND.n1662 GND.n1621 9.3005
R8241 GND.n1624 GND.n1622 9.3005
R8242 GND.n1658 GND.n1625 9.3005
R8243 GND.n1657 GND.n1626 9.3005
R8244 GND.n1656 GND.n1627 9.3005
R8245 GND.n1630 GND.n1628 9.3005
R8246 GND.n1652 GND.n1631 9.3005
R8247 GND.n1651 GND.n1632 9.3005
R8248 GND.n1650 GND.n1633 9.3005
R8249 GND.n1636 GND.n1634 9.3005
R8250 GND.n1646 GND.n1637 9.3005
R8251 GND.n1645 GND.n1638 9.3005
R8252 GND.n1644 GND.n1639 9.3005
R8253 GND.n1642 GND.n1641 9.3005
R8254 GND.n1640 GND.n1491 9.3005
R8255 GND.n1489 GND.n1488 9.3005
R8256 GND.n2046 GND.n2045 9.3005
R8257 GND.n2047 GND.n1487 9.3005
R8258 GND.n4635 GND.n2048 9.3005
R8259 GND.n4634 GND.n2049 9.3005
R8260 GND.n4633 GND.n2050 9.3005
R8261 GND.n2055 GND.n2051 9.3005
R8262 GND.n4627 GND.n2056 9.3005
R8263 GND.n4626 GND.n2057 9.3005
R8264 GND.n4625 GND.n2058 9.3005
R8265 GND.n3470 GND.n2059 9.3005
R8266 GND.n3471 GND.n3469 9.3005
R8267 GND.n3474 GND.n3473 9.3005
R8268 GND.n3472 GND.n2093 9.3005
R8269 GND.n4598 GND.n2094 9.3005
R8270 GND.n4597 GND.n2095 9.3005
R8271 GND.n4596 GND.n2096 9.3005
R8272 GND.n3533 GND.n2097 9.3005
R8273 GND.n3535 GND.n3534 9.3005
R8274 GND.n3532 GND.n3531 9.3005
R8275 GND.n3540 GND.n3539 9.3005
R8276 GND.n3541 GND.n3530 9.3005
R8277 GND.n3551 GND.n3542 9.3005
R8278 GND.n3550 GND.n3543 9.3005
R8279 GND.n3549 GND.n3544 9.3005
R8280 GND.n3547 GND.n3546 9.3005
R8281 GND.n3545 GND.n3155 9.3005
R8282 GND.n3153 GND.n3152 9.3005
R8283 GND.n3590 GND.n3589 9.3005
R8284 GND.n3591 GND.n3151 9.3005
R8285 GND.n3593 GND.n3592 9.3005
R8286 GND.n3143 GND.n3142 9.3005
R8287 GND.n3616 GND.n3615 9.3005
R8288 GND.n3617 GND.n3141 9.3005
R8289 GND.n3628 GND.n3618 9.3005
R8290 GND.n3627 GND.n3619 9.3005
R8291 GND.n3626 GND.n3620 9.3005
R8292 GND.n3623 GND.n3622 9.3005
R8293 GND.n3621 GND.n2217 9.3005
R8294 GND.n4514 GND.n2218 9.3005
R8295 GND.n4513 GND.n2219 9.3005
R8296 GND.n4512 GND.n2220 9.3005
R8297 GND.n2263 GND.n2221 9.3005
R8298 GND.n2265 GND.n2264 9.3005
R8299 GND.n2269 GND.n2268 9.3005
R8300 GND.n2270 GND.n2262 9.3005
R8301 GND.n4487 GND.n2271 9.3005
R8302 GND.n4486 GND.n2272 9.3005
R8303 GND.n4485 GND.n2273 9.3005
R8304 GND.n2306 GND.n2274 9.3005
R8305 GND.n2309 GND.n2308 9.3005
R8306 GND.n2310 GND.n2305 9.3005
R8307 GND.n4466 GND.n2311 9.3005
R8308 GND.n4465 GND.n2312 9.3005
R8309 GND.n4464 GND.n2313 9.3005
R8310 GND.n2350 GND.n2314 9.3005
R8311 GND.n2353 GND.n2352 9.3005
R8312 GND.n2354 GND.n2349 9.3005
R8313 GND.n4445 GND.n2355 9.3005
R8314 GND.n4444 GND.n2356 9.3005
R8315 GND.n4443 GND.n2357 9.3005
R8316 GND.n3024 GND.n2358 9.3005
R8317 GND.n3026 GND.n3025 9.3005
R8318 GND.n4009 GND.n4008 9.3005
R8319 GND.n4010 GND.n3023 9.3005
R8320 GND.n4012 GND.n4011 9.3005
R8321 GND.n3019 GND.n3018 9.3005
R8322 GND.n4020 GND.n4019 9.3005
R8323 GND.n4021 GND.n3017 9.3005
R8324 GND.n4023 GND.n4022 9.3005
R8325 GND.n3015 GND.n3014 9.3005
R8326 GND.n4028 GND.n4027 9.3005
R8327 GND.n4029 GND.n3013 9.3005
R8328 GND.n4031 GND.n4030 9.3005
R8329 GND.n3011 GND.n3010 9.3005
R8330 GND.n4036 GND.n4035 9.3005
R8331 GND.n4037 GND.n3009 9.3005
R8332 GND.n4075 GND.n4038 9.3005
R8333 GND.n4074 GND.n4039 9.3005
R8334 GND.n4073 GND.n4040 9.3005
R8335 GND.n4043 GND.n4041 9.3005
R8336 GND.n4069 GND.n4044 9.3005
R8337 GND.n4068 GND.n4045 9.3005
R8338 GND.n4067 GND.n4046 9.3005
R8339 GND.n4049 GND.n4047 9.3005
R8340 GND.n4063 GND.n4050 9.3005
R8341 GND.n4062 GND.n4051 9.3005
R8342 GND.n4061 GND.n4052 9.3005
R8343 GND.n4054 GND.n4053 9.3005
R8344 GND.n4057 GND.n4056 9.3005
R8345 GND.n4055 GND.n2911 9.3005
R8346 GND.n4299 GND.n2941 9.3005
R8347 GND.n4298 GND.n2942 9.3005
R8348 GND.n2945 GND.n2943 9.3005
R8349 GND.n4294 GND.n2946 9.3005
R8350 GND.n4293 GND.n2947 9.3005
R8351 GND.n4292 GND.n2948 9.3005
R8352 GND.n2951 GND.n2949 9.3005
R8353 GND.n4288 GND.n2952 9.3005
R8354 GND.n4287 GND.n2953 9.3005
R8355 GND.n4286 GND.n2954 9.3005
R8356 GND.n4265 GND.n2955 9.3005
R8357 GND.n4282 GND.n4266 9.3005
R8358 GND.n4281 GND.n4267 9.3005
R8359 GND.n4280 GND.n4268 9.3005
R8360 GND.n4271 GND.n4269 9.3005
R8361 GND.n4276 GND.n4272 9.3005
R8362 GND.n4275 GND.n4274 9.3005
R8363 GND.n4273 GND.n312 9.3005
R8364 GND.n5745 GND.n313 9.3005
R8365 GND.n5744 GND.n314 9.3005
R8366 GND.n5743 GND.n315 9.3005
R8367 GND.n321 GND.n316 9.3005
R8368 GND.n322 GND.n320 9.3005
R8369 GND.n5736 GND.n323 9.3005
R8370 GND.n5735 GND.n324 9.3005
R8371 GND.n5734 GND.n325 9.3005
R8372 GND.n330 GND.n326 9.3005
R8373 GND.n5728 GND.n331 9.3005
R8374 GND.n5727 GND.n332 9.3005
R8375 GND.n5726 GND.n333 9.3005
R8376 GND.n338 GND.n334 9.3005
R8377 GND.n5720 GND.n339 9.3005
R8378 GND.n5719 GND.n340 9.3005
R8379 GND.n5718 GND.n341 9.3005
R8380 GND.n346 GND.n342 9.3005
R8381 GND.n5712 GND.n347 9.3005
R8382 GND.n5711 GND.n348 9.3005
R8383 GND.n5710 GND.n349 9.3005
R8384 GND.n354 GND.n350 9.3005
R8385 GND.n5704 GND.n355 9.3005
R8386 GND.n5703 GND.n356 9.3005
R8387 GND.n5702 GND.n357 9.3005
R8388 GND.n362 GND.n358 9.3005
R8389 GND.n5696 GND.n363 9.3005
R8390 GND.n5695 GND.n364 9.3005
R8391 GND.n5694 GND.n365 9.3005
R8392 GND.n370 GND.n366 9.3005
R8393 GND.n5688 GND.n371 9.3005
R8394 GND.n5687 GND.n372 9.3005
R8395 GND.n5686 GND.n373 9.3005
R8396 GND.n1070 GND.n1069 9.3005
R8397 GND.n1068 GND.n1018 9.3005
R8398 GND.n1067 GND.n1066 9.3005
R8399 GND.n1063 GND.n1021 9.3005
R8400 GND.n1062 GND.n1059 9.3005
R8401 GND.n1058 GND.n1022 9.3005
R8402 GND.n1057 GND.n1056 9.3005
R8403 GND.n1053 GND.n1023 9.3005
R8404 GND.n1052 GND.n1027 9.3005
R8405 GND.n1047 GND.n1028 9.3005
R8406 GND.n1046 GND.n1045 9.3005
R8407 GND.n1042 GND.n1029 9.3005
R8408 GND.n1039 GND.n1038 9.3005
R8409 GND.n1037 GND.n1030 9.3005
R8410 GND.n1036 GND.n1035 9.3005
R8411 GND.n1032 GND.n1031 9.3005
R8412 GND.n1049 GND.n1048 9.3005
R8413 GND.n1071 GND.n1014 9.3005
R8414 GND.n1073 GND.n1072 9.3005
R8415 GND.n4776 GND.n1000 9.3005
R8416 GND.n4775 GND.n1001 9.3005
R8417 GND.n1730 GND.n1002 9.3005
R8418 GND.n1732 GND.n1731 9.3005
R8419 GND.n1825 GND.n1824 9.3005
R8420 GND.n1826 GND.n1729 9.3005
R8421 GND.n1830 GND.n1827 9.3005
R8422 GND.n1829 GND.n1828 9.3005
R8423 GND.n1708 GND.n1707 9.3005
R8424 GND.n1850 GND.n1849 9.3005
R8425 GND.n1851 GND.n1706 9.3005
R8426 GND.n1855 GND.n1852 9.3005
R8427 GND.n1854 GND.n1853 9.3005
R8428 GND.n1686 GND.n1685 9.3005
R8429 GND.n1875 GND.n1874 9.3005
R8430 GND.n1876 GND.n1684 9.3005
R8431 GND.n1878 GND.n1877 9.3005
R8432 GND.n1578 GND.n1571 9.3005
R8433 GND.n1951 GND.n1948 9.3005
R8434 GND.n1950 GND.n1949 9.3005
R8435 GND.n1550 GND.n1549 9.3005
R8436 GND.n1971 GND.n1970 9.3005
R8437 GND.n1972 GND.n1548 9.3005
R8438 GND.n1976 GND.n1973 9.3005
R8439 GND.n1975 GND.n1974 9.3005
R8440 GND.n1527 GND.n1526 9.3005
R8441 GND.n1995 GND.n1994 9.3005
R8442 GND.n1996 GND.n1525 9.3005
R8443 GND.n2000 GND.n1997 9.3005
R8444 GND.n1999 GND.n1998 9.3005
R8445 GND.n1504 GND.n1503 9.3005
R8446 GND.n2029 GND.n2028 9.3005
R8447 GND.n2030 GND.n1502 9.3005
R8448 GND.n2034 GND.n2031 9.3005
R8449 GND.n2033 GND.n2032 9.3005
R8450 GND.n1178 GND.n1177 9.3005
R8451 GND.n4698 GND.n4697 9.3005
R8452 GND.n4777 GND.n999 9.3005
R8453 GND.n1947 GND.n1576 9.3005
R8454 GND.n1947 GND.n1570 9.3005
R8455 GND.n909 GND.n908 9.3005
R8456 GND.n4854 GND.n913 9.3005
R8457 GND.n4853 GND.n914 9.3005
R8458 GND.n4852 GND.n915 9.3005
R8459 GND.n920 GND.n916 9.3005
R8460 GND.n4846 GND.n921 9.3005
R8461 GND.n4845 GND.n922 9.3005
R8462 GND.n4844 GND.n923 9.3005
R8463 GND.n928 GND.n924 9.3005
R8464 GND.n4838 GND.n929 9.3005
R8465 GND.n4837 GND.n930 9.3005
R8466 GND.n4836 GND.n931 9.3005
R8467 GND.n936 GND.n932 9.3005
R8468 GND.n4830 GND.n937 9.3005
R8469 GND.n4829 GND.n938 9.3005
R8470 GND.n4828 GND.n939 9.3005
R8471 GND.n944 GND.n940 9.3005
R8472 GND.n4822 GND.n945 9.3005
R8473 GND.n4821 GND.n946 9.3005
R8474 GND.n4820 GND.n947 9.3005
R8475 GND.n952 GND.n948 9.3005
R8476 GND.n4814 GND.n953 9.3005
R8477 GND.n4813 GND.n954 9.3005
R8478 GND.n4812 GND.n955 9.3005
R8479 GND.n960 GND.n956 9.3005
R8480 GND.n4806 GND.n961 9.3005
R8481 GND.n4805 GND.n962 9.3005
R8482 GND.n4804 GND.n963 9.3005
R8483 GND.n1745 GND.n964 9.3005
R8484 GND.n1747 GND.n1746 9.3005
R8485 GND.n1751 GND.n1750 9.3005
R8486 GND.n1752 GND.n1744 9.3005
R8487 GND.n1754 GND.n1753 9.3005
R8488 GND.n1742 GND.n1741 9.3005
R8489 GND.n1775 GND.n1774 9.3005
R8490 GND.n1776 GND.n1740 9.3005
R8491 GND.n1816 GND.n1777 9.3005
R8492 GND.n1815 GND.n1778 9.3005
R8493 GND.n1814 GND.n1779 9.3005
R8494 GND.n1782 GND.n1780 9.3005
R8495 GND.n1810 GND.n1783 9.3005
R8496 GND.n1809 GND.n1784 9.3005
R8497 GND.n1808 GND.n1785 9.3005
R8498 GND.n1788 GND.n1786 9.3005
R8499 GND.n1804 GND.n1789 9.3005
R8500 GND.n1803 GND.n1790 9.3005
R8501 GND.n1802 GND.n1791 9.3005
R8502 GND.n1794 GND.n1792 9.3005
R8503 GND.n1798 GND.n1795 9.3005
R8504 GND.n4861 GND.n4860 9.3005
R8505 GND.n4864 GND.n907 9.3005
R8506 GND.n906 GND.n902 9.3005
R8507 GND.n4870 GND.n901 9.3005
R8508 GND.n4871 GND.n900 9.3005
R8509 GND.n4872 GND.n899 9.3005
R8510 GND.n898 GND.n894 9.3005
R8511 GND.n4878 GND.n893 9.3005
R8512 GND.n4879 GND.n892 9.3005
R8513 GND.n4880 GND.n891 9.3005
R8514 GND.n890 GND.n886 9.3005
R8515 GND.n4886 GND.n885 9.3005
R8516 GND.n4887 GND.n884 9.3005
R8517 GND.n4888 GND.n883 9.3005
R8518 GND.n882 GND.n878 9.3005
R8519 GND.n4894 GND.n877 9.3005
R8520 GND.n4895 GND.n876 9.3005
R8521 GND.n4896 GND.n875 9.3005
R8522 GND.n874 GND.n870 9.3005
R8523 GND.n4902 GND.n869 9.3005
R8524 GND.n4903 GND.n868 9.3005
R8525 GND.n4904 GND.n867 9.3005
R8526 GND.n866 GND.n862 9.3005
R8527 GND.n4910 GND.n861 9.3005
R8528 GND.n4911 GND.n860 9.3005
R8529 GND.n4912 GND.n859 9.3005
R8530 GND.n858 GND.n854 9.3005
R8531 GND.n4918 GND.n853 9.3005
R8532 GND.n4919 GND.n852 9.3005
R8533 GND.n4920 GND.n851 9.3005
R8534 GND.n850 GND.n846 9.3005
R8535 GND.n4926 GND.n845 9.3005
R8536 GND.n4927 GND.n844 9.3005
R8537 GND.n4928 GND.n843 9.3005
R8538 GND.n842 GND.n838 9.3005
R8539 GND.n4934 GND.n837 9.3005
R8540 GND.n4935 GND.n836 9.3005
R8541 GND.n4936 GND.n835 9.3005
R8542 GND.n834 GND.n830 9.3005
R8543 GND.n4942 GND.n829 9.3005
R8544 GND.n4943 GND.n828 9.3005
R8545 GND.n4944 GND.n827 9.3005
R8546 GND.n826 GND.n822 9.3005
R8547 GND.n4950 GND.n821 9.3005
R8548 GND.n4951 GND.n820 9.3005
R8549 GND.n4952 GND.n819 9.3005
R8550 GND.n818 GND.n814 9.3005
R8551 GND.n4958 GND.n813 9.3005
R8552 GND.n4959 GND.n812 9.3005
R8553 GND.n4960 GND.n811 9.3005
R8554 GND.n810 GND.n806 9.3005
R8555 GND.n4966 GND.n805 9.3005
R8556 GND.n4967 GND.n804 9.3005
R8557 GND.n4968 GND.n803 9.3005
R8558 GND.n802 GND.n798 9.3005
R8559 GND.n4863 GND.n4862 9.3005
R8560 GND.n1896 GND.n1670 9.3005
R8561 GND.n1898 GND.n1897 9.3005
R8562 GND.n1899 GND.n1669 9.3005
R8563 GND.n1901 GND.n1900 9.3005
R8564 GND.n1562 GND.n1561 9.3005
R8565 GND.n1956 GND.n1955 9.3005
R8566 GND.n1957 GND.n1559 9.3005
R8567 GND.n1960 GND.n1959 9.3005
R8568 GND.n1958 GND.n1560 9.3005
R8569 GND.n1540 GND.n1539 9.3005
R8570 GND.n1981 GND.n1980 9.3005
R8571 GND.n1982 GND.n1537 9.3005
R8572 GND.n1985 GND.n1984 9.3005
R8573 GND.n1983 GND.n1538 9.3005
R8574 GND.n1516 GND.n1515 9.3005
R8575 GND.n2005 GND.n2004 9.3005
R8576 GND.n2006 GND.n1513 9.3005
R8577 GND.n2021 GND.n2020 9.3005
R8578 GND.n2019 GND.n1514 9.3005
R8579 GND.n2018 GND.n2017 9.3005
R8580 GND.n2016 GND.n2007 9.3005
R8581 GND.n2015 GND.n2014 9.3005
R8582 GND.n2013 GND.n2012 9.3005
R8583 GND.n2011 GND.n1476 9.3005
R8584 GND.n4666 GND.n1205 9.3005
R8585 GND.n4665 GND.n4664 9.3005
R8586 GND.n4663 GND.n1209 9.3005
R8587 GND.n4661 GND.n4660 9.3005
R8588 GND.n4659 GND.n1467 9.3005
R8589 GND.n4658 GND.n4657 9.3005
R8590 GND.n4656 GND.n1473 9.3005
R8591 GND.n4654 GND.n4653 9.3005
R8592 GND.n4668 GND.n4667 9.3005
R8593 GND.n4688 GND.n1183 9.3005
R8594 GND.n4690 GND.n4689 9.3005
R8595 GND.n4691 GND.n1182 9.3005
R8596 GND.n4693 GND.n4692 9.3005
R8597 GND.n4694 GND.n1179 9.3005
R8598 GND.n4696 GND.n4695 9.3005
R8599 GND.n4686 GND.n4685 9.3005
R8600 GND.n4684 GND.n1192 9.3005
R8601 GND.n4683 GND.n4682 9.3005
R8602 GND.n4681 GND.n1193 9.3005
R8603 GND.n4680 GND.n4679 9.3005
R8604 GND.n4678 GND.n1197 9.3005
R8605 GND.n4677 GND.n4676 9.3005
R8606 GND.n4675 GND.n1198 9.3005
R8607 GND.n4674 GND.n4673 9.3005
R8608 GND.n4672 GND.n1204 9.3005
R8609 GND.n4671 GND.n4670 9.3005
R8610 GND.n1012 GND.n1010 9.3005
R8611 GND.n4771 GND.n4770 9.3005
R8612 GND.n1013 GND.n1011 9.3005
R8613 GND.n4766 GND.n1084 9.3005
R8614 GND.n4765 GND.n1085 9.3005
R8615 GND.n4764 GND.n1086 9.3005
R8616 GND.n1724 GND.n1087 9.3005
R8617 GND.n4760 GND.n1092 9.3005
R8618 GND.n4759 GND.n1093 9.3005
R8619 GND.n4758 GND.n1094 9.3005
R8620 GND.n1843 GND.n1095 9.3005
R8621 GND.n4754 GND.n1100 9.3005
R8622 GND.n4753 GND.n1101 9.3005
R8623 GND.n4752 GND.n1102 9.3005
R8624 GND.n1870 GND.n1103 9.3005
R8625 GND.n4748 GND.n1108 9.3005
R8626 GND.n4747 GND.n1109 9.3005
R8627 GND.n4746 GND.n1110 9.3005
R8628 GND.n1941 GND.n1111 9.3005
R8629 GND.n4742 GND.n1116 9.3005
R8630 GND.n4741 GND.n1117 9.3005
R8631 GND.n4740 GND.n1118 9.3005
R8632 GND.n1599 GND.n1119 9.3005
R8633 GND.n4736 GND.n1124 9.3005
R8634 GND.n4735 GND.n1125 9.3005
R8635 GND.n4734 GND.n1126 9.3005
R8636 GND.n1910 GND.n1127 9.3005
R8637 GND.n4730 GND.n1132 9.3005
R8638 GND.n4729 GND.n1133 9.3005
R8639 GND.n4728 GND.n1134 9.3005
R8640 GND.n1556 GND.n1135 9.3005
R8641 GND.n4724 GND.n1140 9.3005
R8642 GND.n4723 GND.n1141 9.3005
R8643 GND.n4722 GND.n1142 9.3005
R8644 GND.n1533 GND.n1143 9.3005
R8645 GND.n4718 GND.n1148 9.3005
R8646 GND.n4717 GND.n1149 9.3005
R8647 GND.n4716 GND.n1150 9.3005
R8648 GND.n1520 GND.n1151 9.3005
R8649 GND.n4712 GND.n1156 9.3005
R8650 GND.n4711 GND.n1157 9.3005
R8651 GND.n4710 GND.n1158 9.3005
R8652 GND.n1495 GND.n1159 9.3005
R8653 GND.n4706 GND.n1164 9.3005
R8654 GND.n4705 GND.n1165 9.3005
R8655 GND.n4704 GND.n1166 9.3005
R8656 GND.n1173 GND.n1167 9.3005
R8657 GND.n1076 GND.n1075 9.3005
R8658 GND.n1080 GND.n1012 9.3005
R8659 GND.n4770 GND.n4769 9.3005
R8660 GND.n4768 GND.n1013 9.3005
R8661 GND.n4767 GND.n4766 9.3005
R8662 GND.n4765 GND.n1083 9.3005
R8663 GND.n4764 GND.n4763 9.3005
R8664 GND.n4762 GND.n1087 9.3005
R8665 GND.n4761 GND.n4760 9.3005
R8666 GND.n4759 GND.n1091 9.3005
R8667 GND.n4758 GND.n4757 9.3005
R8668 GND.n4756 GND.n1095 9.3005
R8669 GND.n4755 GND.n4754 9.3005
R8670 GND.n4753 GND.n1099 9.3005
R8671 GND.n4752 GND.n4751 9.3005
R8672 GND.n4750 GND.n1103 9.3005
R8673 GND.n4749 GND.n4748 9.3005
R8674 GND.n4747 GND.n1107 9.3005
R8675 GND.n4746 GND.n4745 9.3005
R8676 GND.n4744 GND.n1111 9.3005
R8677 GND.n4743 GND.n4742 9.3005
R8678 GND.n4741 GND.n1115 9.3005
R8679 GND.n4740 GND.n4739 9.3005
R8680 GND.n4738 GND.n1119 9.3005
R8681 GND.n4737 GND.n4736 9.3005
R8682 GND.n4735 GND.n1123 9.3005
R8683 GND.n4734 GND.n4733 9.3005
R8684 GND.n4732 GND.n1127 9.3005
R8685 GND.n4731 GND.n4730 9.3005
R8686 GND.n4729 GND.n1131 9.3005
R8687 GND.n4728 GND.n4727 9.3005
R8688 GND.n4726 GND.n1135 9.3005
R8689 GND.n4725 GND.n4724 9.3005
R8690 GND.n4723 GND.n1139 9.3005
R8691 GND.n4722 GND.n4721 9.3005
R8692 GND.n4720 GND.n1143 9.3005
R8693 GND.n4719 GND.n4718 9.3005
R8694 GND.n4717 GND.n1147 9.3005
R8695 GND.n4716 GND.n4715 9.3005
R8696 GND.n4714 GND.n1151 9.3005
R8697 GND.n4713 GND.n4712 9.3005
R8698 GND.n4711 GND.n1155 9.3005
R8699 GND.n4710 GND.n4709 9.3005
R8700 GND.n4708 GND.n1159 9.3005
R8701 GND.n4707 GND.n4706 9.3005
R8702 GND.n4705 GND.n1163 9.3005
R8703 GND.n4704 GND.n4703 9.3005
R8704 GND.n4702 GND.n1167 9.3005
R8705 GND.n1077 GND.n1076 9.3005
R8706 GND.n4789 GND.n990 9.3005
R8707 GND.n4791 GND.n4790 9.3005
R8708 GND.n4792 GND.n985 9.3005
R8709 GND.n4794 GND.n4793 9.3005
R8710 GND.n4795 GND.n984 9.3005
R8711 GND.n4797 GND.n4796 9.3005
R8712 GND.n4798 GND.n983 9.3005
R8713 GND.n4788 GND.n4787 9.3005
R8714 GND.n4782 GND.n991 9.3005
R8715 GND.n1763 GND.n1762 9.3005
R8716 GND.n1765 GND.n1764 9.3005
R8717 GND.n1766 GND.n1759 9.3005
R8718 GND.n1769 GND.n1768 9.3005
R8719 GND.n1767 GND.n1760 9.3005
R8720 GND.n1720 GND.n1719 9.3005
R8721 GND.n1835 GND.n1834 9.3005
R8722 GND.n1836 GND.n1717 9.3005
R8723 GND.n1839 GND.n1838 9.3005
R8724 GND.n1837 GND.n1718 9.3005
R8725 GND.n1697 GND.n1696 9.3005
R8726 GND.n1860 GND.n1859 9.3005
R8727 GND.n1861 GND.n1694 9.3005
R8728 GND.n1864 GND.n1863 9.3005
R8729 GND.n1862 GND.n1695 9.3005
R8730 GND.n1675 GND.n1674 9.3005
R8731 GND.n1883 GND.n1882 9.3005
R8732 GND.n1884 GND.n1673 9.3005
R8733 GND.n1886 GND.n1885 9.3005
R8734 GND.n1887 GND.n1672 9.3005
R8735 GND.n1891 GND.n1890 9.3005
R8736 GND.n1892 GND.n1671 9.3005
R8737 GND.n1895 GND.n1894 9.3005
R8738 GND.n1761 GND.n993 9.3005
R8739 GND.n3498 GND.n3192 8.97305
R8740 GND.n4572 GND.n2137 8.97305
R8741 GND.n3110 GND.n3109 8.97305
R8742 GND.n3780 GND.n3769 8.97305
R8743 GND.n3090 GND.t45 8.97305
R8744 GND.n1450 GND.n1449 8.92171
R8745 GND.n1228 GND.n1227 8.92171
R8746 GND.n2486 GND.n2485 8.92171
R8747 GND.n2451 GND.n2450 8.92171
R8748 GND.n5864 GND.n5863 8.76487
R8749 GND.n1893 GND.n71 8.76487
R8750 GND.n1680 GND.t22 8.28285
R8751 GND.n1953 GND.t10 8.28285
R8752 GND.t48 GND.n2063 8.28285
R8753 GND.n3498 GND.n3489 8.28285
R8754 GND.n4573 GND.n4572 8.28285
R8755 GND.n4538 GND.n4537 8.28285
R8756 GND.n3678 GND.n3126 8.28285
R8757 GND.n3747 GND.n3110 8.28285
R8758 GND.n3780 GND.n3768 8.28285
R8759 GND.n4434 GND.t45 8.28285
R8760 GND.n4333 GND.t20 8.28285
R8761 GND.n4171 GND.t29 8.28285
R8762 GND.n1446 GND.n1440 8.14595
R8763 GND.n1224 GND.n1218 8.14595
R8764 GND.n2482 GND.n2476 8.14595
R8765 GND.n2447 GND.n2441 8.14595
R8766 GND.n3286 GND.t87 7.59266
R8767 GND.n3462 GND.n2082 7.59266
R8768 GND.n3156 GND.n2146 7.59266
R8769 GND.t14 GND.n4558 7.59266
R8770 GND.n3595 GND.n2174 7.59266
R8771 GND.n3684 GND.n2231 7.59266
R8772 GND.n3691 GND.t8 7.59266
R8773 GND.n3719 GND.n3116 7.59266
R8774 GND.n3773 GND.n3096 7.59266
R8775 GND.n4653 GND.n1473 7.56414
R8776 GND.n4243 GND.n4241 7.56414
R8777 GND.n4427 GND.n2379 7.56414
R8778 GND.n4787 GND.n4782 7.56414
R8779 GND.n1445 GND.n1442 7.3702
R8780 GND.n1223 GND.n1220 7.3702
R8781 GND.n2481 GND.n2478 7.3702
R8782 GND.n2446 GND.n2443 7.3702
R8783 GND.n2709 GND.n2674 7.28789
R8784 GND.n2570 GND.n2535 7.28789
R8785 GND.n46 GND.n22 6.9186
R8786 GND.n118 GND.n94 6.9186
R8787 GND.n3507 GND.n3186 6.90246
R8788 GND.n4579 GND.n2126 6.90246
R8789 GND.n4531 GND.n2192 6.90246
R8790 GND.n3671 GND.n3129 6.90246
R8791 GND.n3740 GND.n2300 6.90246
R8792 GND.n3727 GND.n2318 6.90246
R8793 GND.n1296 GND.n1295 6.52659
R8794 GND.n1428 GND.n1427 6.52659
R8795 GND.n1293 GND.n1292 6.40821
R8796 GND.n5777 GND.n5774 6.4005
R8797 GND.n1052 GND.n1026 6.4005
R8798 GND.n2780 GND.n2640 6.31255
R8799 GND.n3455 GND.n2069 6.21226
R8800 GND.n3286 GND.n2072 6.21226
R8801 GND.n4558 GND.n2157 6.21226
R8802 GND.n4552 GND.n2163 6.21226
R8803 GND.n3697 GND.n2248 6.21226
R8804 GND.n3691 GND.n2251 6.21226
R8805 GND.n3787 GND.n2367 6.21226
R8806 GND.n3891 GND.n3090 6.21226
R8807 GND.n2780 GND.n2779 6.01802
R8808 GND.n4537 GND.t32 5.86717
R8809 GND.n3126 GND.t4 5.86717
R8810 GND.n1446 GND.n1445 5.81868
R8811 GND.n1224 GND.n1223 5.81868
R8812 GND.n2482 GND.n2481 5.81868
R8813 GND.n2447 GND.n2446 5.81868
R8814 GND.n1909 GND.t10 5.52207
R8815 GND.t61 GND.n2088 5.52207
R8816 GND.n4587 GND.n4586 5.52207
R8817 GND.n3660 GND.n3659 5.52207
R8818 GND.n4524 GND.n4523 5.52207
R8819 GND.n3733 GND.n2316 5.52207
R8820 GND.t77 GND.n3772 5.52207
R8821 GND.n2905 GND.t20 5.52207
R8822 GND.t7 GND.n3515 5.17697
R8823 GND.t3 GND.n2302 5.17697
R8824 GND.n2779 GND.n2778 5.05683
R8825 GND.n2744 GND.n2743 5.05683
R8826 GND.n2709 GND.n2708 5.05683
R8827 GND.n2640 GND.n2639 5.05683
R8828 GND.n2605 GND.n2604 5.05683
R8829 GND.n2570 GND.n2569 5.05683
R8830 GND.n1449 GND.n1440 5.04292
R8831 GND.n1227 GND.n1218 5.04292
R8832 GND.n2485 GND.n2476 5.04292
R8833 GND.n2450 GND.n2441 5.04292
R8834 GND.n3843 GND.n3837 5.04292
R8835 GND.n3242 GND.n3232 5.04292
R8836 GND.n1430 GND.n1429 4.96553
R8837 GND.n70 GND.n69 4.94662
R8838 GND.n142 GND.n141 4.94662
R8839 GND.n46 GND.n45 4.88412
R8840 GND.n118 GND.n117 4.88412
R8841 GND.t55 GND.n1506 4.83187
R8842 GND.n4623 GND.n4622 4.83187
R8843 GND.n3477 GND.n3476 4.83187
R8844 GND.n3149 GND.n2166 4.83187
R8845 GND.n3613 GND.t0 4.83187
R8846 GND.n3679 GND.t12 4.83187
R8847 GND.n3122 GND.n2234 4.83187
R8848 GND.n4441 GND.n4440 4.83187
R8849 GND.n4006 GND.n3028 4.83187
R8850 GND.t100 GND.n4005 4.83187
R8851 GND.n4077 GND.t37 4.83187
R8852 GND.n4330 GND.n163 4.74817
R8853 GND.n161 GND.n155 4.74817
R8854 GND.n5856 GND.n156 4.74817
R8855 GND.n164 GND.n160 4.74817
R8856 GND.n2903 GND.n163 4.74817
R8857 GND.n4317 GND.n161 4.74817
R8858 GND.n5857 GND.n5856 4.74817
R8859 GND.n2929 GND.n160 4.74817
R8860 GND.n1797 GND.n1796 4.74817
R8861 GND.n1935 GND.n1934 4.74817
R8862 GND.n1613 GND.n1592 4.74817
R8863 GND.n1919 GND.n1615 4.74817
R8864 GND.n1917 GND.n1916 4.74817
R8865 GND.n4324 GND.n4323 4.74817
R8866 GND.n2934 GND.n2912 4.74817
R8867 GND.n2938 GND.n2937 4.74817
R8868 GND.n4305 GND.n4304 4.74817
R8869 GND.n4300 GND.n2939 4.74817
R8870 GND.n4325 GND.n4324 4.74817
R8871 GND.n4322 GND.n2912 4.74817
R8872 GND.n2937 GND.n2936 4.74817
R8873 GND.n4306 GND.n4305 4.74817
R8874 GND.n4303 GND.n2939 4.74817
R8875 GND.n1946 GND.n1945 4.74817
R8876 GND.n1928 GND.n1575 4.74817
R8877 GND.n1903 GND.n1574 4.74817
R8878 GND.n1906 GND.n1573 4.74817
R8879 GND.n1946 GND.n1577 4.74817
R8880 GND.n1602 GND.n1575 4.74817
R8881 GND.n1927 GND.n1574 4.74817
R8882 GND.n1904 GND.n1573 4.74817
R8883 GND.n1796 GND.n1591 4.74817
R8884 GND.n1936 GND.n1935 4.74817
R8885 GND.n1933 GND.n1592 4.74817
R8886 GND.n1615 GND.n1614 4.74817
R8887 GND.n1918 GND.n1917 4.74817
R8888 GND.n50 GND.n48 4.69785
R8889 GND.n61 GND.n59 4.69785
R8890 GND.n26 GND.n24 4.69785
R8891 GND.n37 GND.n35 4.69785
R8892 GND.n3 GND.n1 4.69785
R8893 GND.n14 GND.n12 4.69785
R8894 GND.n133 GND.n131 4.69785
R8895 GND.n122 GND.n120 4.69785
R8896 GND.n109 GND.n107 4.69785
R8897 GND.n98 GND.n96 4.69785
R8898 GND.n86 GND.n84 4.69785
R8899 GND.n75 GND.n73 4.69785
R8900 GND.n4413 GND.n2407 4.6132
R8901 GND.n4687 GND.n1188 4.6132
R8902 GND.t2 GND.n2154 4.48677
R8903 GND.n4490 GND.t19 4.48677
R8904 GND.n2770 GND.n2769 4.38232
R8905 GND.n2755 GND.n2752 4.38232
R8906 GND.n2735 GND.n2734 4.38232
R8907 GND.n2720 GND.n2717 4.38232
R8908 GND.n2700 GND.n2699 4.38232
R8909 GND.n2685 GND.n2682 4.38232
R8910 GND.n2666 GND.n2665 4.38232
R8911 GND.n2651 GND.n2648 4.38232
R8912 GND.n2616 GND.n2613 4.38232
R8913 GND.n2631 GND.n2630 4.38232
R8914 GND.n2581 GND.n2578 4.38232
R8915 GND.n2596 GND.n2595 4.38232
R8916 GND.n2546 GND.n2543 4.38232
R8917 GND.n2561 GND.n2560 4.38232
R8918 GND.n2512 GND.n2509 4.38232
R8919 GND.n2527 GND.n2526 4.38232
R8920 GND.n1450 GND.n1438 4.26717
R8921 GND.n1228 GND.n1216 4.26717
R8922 GND.n2486 GND.n2474 4.26717
R8923 GND.n2451 GND.n2439 4.26717
R8924 GND.n3462 GND.t61 4.14168
R8925 GND.n4593 GND.n2101 4.14168
R8926 GND.n3554 GND.n3526 4.14168
R8927 GND.n4538 GND.t0 4.14168
R8928 GND.n3634 GND.n3633 4.14168
R8929 GND.n4517 GND.n2212 4.14168
R8930 GND.t12 GND.n3678 4.14168
R8931 GND.n4476 GND.n4475 4.14168
R8932 GND.n4455 GND.n4454 4.14168
R8933 GND.n3773 GND.t77 4.14168
R8934 GND.n3037 GND.n3034 3.68535
R8935 GND.n1454 GND.n1453 3.49141
R8936 GND.n1232 GND.n1231 3.49141
R8937 GND.n2490 GND.n2489 3.49141
R8938 GND.n2455 GND.n2454 3.49141
R8939 GND.n3478 GND.t87 3.45148
R8940 GND.n4601 GND.n4600 3.45148
R8941 GND.n4566 GND.n2143 3.45148
R8942 GND.n4559 GND.t14 3.45148
R8943 GND.n4544 GND.n2177 3.45148
R8944 GND.n4510 GND.n4509 3.45148
R8945 GND.t8 GND.n2257 3.45148
R8946 GND.n4483 GND.n2276 3.45148
R8947 GND.n4447 GND.n2346 3.45148
R8948 GND.n2781 GND.n2780 3.4105
R8949 GND.n1428 GND.n1247 3.2808
R8950 GND.n70 GND.n46 3.12126
R8951 GND.n142 GND.n118 3.12126
R8952 GND.n4629 GND.n2053 3.10638
R8953 GND.n4014 GND.n3021 3.10638
R8954 GND.n1245 GND.t15 3.06078
R8955 GND.n1245 GND.t1 3.06078
R8956 GND.n1243 GND.t9 3.06078
R8957 GND.n1243 GND.t28 3.06078
R8958 GND.n2783 GND.t125 3.06078
R8959 GND.n2783 GND.t17 3.06078
R8960 GND.n2466 GND.t35 3.06078
R8961 GND.n2466 GND.t25 3.06078
R8962 GND.n1397 GND.n1396 2.95152
R8963 GND.n1426 GND.n1425 2.95152
R8964 GND.n1364 GND.n1363 2.95152
R8965 GND.n1393 GND.n1392 2.95152
R8966 GND.n1331 GND.n1330 2.95152
R8967 GND.n1360 GND.n1359 2.95152
R8968 GND.n1298 GND.n1297 2.95152
R8969 GND.n1327 GND.n1326 2.95152
R8970 GND.n1444 GND.n1443 2.84308
R8971 GND.n2480 GND.n2479 2.84308
R8972 GND.n1222 GND.n1221 2.84308
R8973 GND.n2445 GND.n2444 2.84308
R8974 GND.n3209 GND.t103 2.76128
R8975 GND.n3455 GND.t48 2.76128
R8976 GND.n3191 GND.n2090 2.76128
R8977 GND.n3564 GND.n3563 2.76128
R8978 GND.n3612 GND.n3145 2.76128
R8979 GND.n3680 GND.n2223 2.76128
R8980 GND.n4482 GND.n2278 2.76128
R8981 GND.n4448 GND.n2344 2.76128
R8982 GND.n1457 GND.n1436 2.71565
R8983 GND.n1235 GND.n1214 2.71565
R8984 GND.n2493 GND.n2472 2.71565
R8985 GND.n2458 GND.n2437 2.71565
R8986 GND.n5855 GND.n163 2.27742
R8987 GND.n5855 GND.n161 2.27742
R8988 GND.n5856 GND.n5855 2.27742
R8989 GND.n5855 GND.n160 2.27742
R8990 GND.n4324 GND.n159 2.27742
R8991 GND.n2912 GND.n159 2.27742
R8992 GND.n2937 GND.n159 2.27742
R8993 GND.n4305 GND.n159 2.27742
R8994 GND.n2939 GND.n159 2.27742
R8995 GND.n1947 GND.n1946 2.27742
R8996 GND.n1947 GND.n1575 2.27742
R8997 GND.n1947 GND.n1574 2.27742
R8998 GND.n1947 GND.n1573 2.27742
R8999 GND.n1796 GND.n1572 2.27742
R9000 GND.n1935 GND.n1572 2.27742
R9001 GND.n1592 GND.n1572 2.27742
R9002 GND.n1615 GND.n1572 2.27742
R9003 GND.n1917 GND.n1572 2.27742
R9004 GND.n2744 GND.n2709 2.23535
R9005 GND.n2605 GND.n2570 2.23535
R9006 GND.n2779 GND.n2744 2.23156
R9007 GND.n2640 GND.n2605 2.23156
R9008 GND.n1818 GND.t96 2.07109
R9009 GND.n3278 GND.n3209 2.07109
R9010 GND.n4594 GND.n2099 2.07109
R9011 GND.n3527 GND.t5 2.07109
R9012 GND.n3553 GND.n2134 2.07109
R9013 GND.n3606 GND.n3137 2.07109
R9014 GND.n4516 GND.n2214 2.07109
R9015 GND.n3746 GND.n2292 2.07109
R9016 GND.n3739 GND.t16 2.07109
R9017 GND.n3101 GND.n2327 2.07109
R9018 GND.n3881 GND.n3030 2.07109
R9019 GND.t70 GND.n4014 2.07109
R9020 GND.n4263 GND.t73 2.07109
R9021 GND.n1362 GND.n1361 2.02238
R9022 GND.n57 GND.n47 1.93989
R9023 GND.n68 GND.n58 1.93989
R9024 GND.n33 GND.n23 1.93989
R9025 GND.n44 GND.n34 1.93989
R9026 GND.n10 GND.n0 1.93989
R9027 GND.n21 GND.n11 1.93989
R9028 GND.n1458 GND.n1434 1.93989
R9029 GND.n1236 GND.n1212 1.93989
R9030 GND.n140 GND.n130 1.93989
R9031 GND.n129 GND.n119 1.93989
R9032 GND.n116 GND.n106 1.93989
R9033 GND.n105 GND.n95 1.93989
R9034 GND.n93 GND.n83 1.93989
R9035 GND.n82 GND.n72 1.93989
R9036 GND.n2494 GND.n2470 1.93989
R9037 GND.n2459 GND.n2435 1.93989
R9038 GND.n1465 GND.n1431 1.75199
R9039 GND.n3840 GND.n3837 1.55202
R9040 GND.n3239 GND.n3232 1.55202
R9041 GND.n1430 GND.n1246 1.4053
R9042 GND.n4608 GND.n4607 1.38089
R9043 GND.n3584 GND.n3159 1.38089
R9044 GND.n3598 GND.n3148 1.38089
R9045 GND.n4503 GND.n4502 1.38089
R9046 GND.n3115 GND.n2259 1.38089
R9047 GND.n3799 GND.n3793 1.38089
R9048 GND.n3071 GND.n3066 1.24928
R9049 GND.n3304 GND.n3303 1.24928
R9050 GND.n3386 GND.n3310 1.24928
R9051 GND.n3958 GND.n3957 1.24928
R9052 GND.n1329 GND.n1328 1.2364
R9053 GND.n1395 GND.n1394 1.2364
R9054 GND.n55 GND.n54 1.16414
R9055 GND.n66 GND.n65 1.16414
R9056 GND.n31 GND.n30 1.16414
R9057 GND.n42 GND.n41 1.16414
R9058 GND.n8 GND.n7 1.16414
R9059 GND.n19 GND.n18 1.16414
R9060 GND.n1462 GND.n1461 1.16414
R9061 GND.n1240 GND.n1239 1.16414
R9062 GND.n138 GND.n137 1.16414
R9063 GND.n127 GND.n126 1.16414
R9064 GND.n114 GND.n113 1.16414
R9065 GND.n103 GND.n102 1.16414
R9066 GND.n91 GND.n90 1.16414
R9067 GND.n80 GND.n79 1.16414
R9068 GND.n2498 GND.n2497 1.16414
R9069 GND.n2463 GND.n2462 1.16414
R9070 GND.n4608 GND.t41 1.03579
R9071 GND.n3799 GND.t51 1.03579
R9072 GND.n1295 GND.n1294 1.02891
R9073 GND.n1407 GND.n1255 0.984173
R9074 GND.n1415 GND.n1251 0.984173
R9075 GND.n1374 GND.n1266 0.984173
R9076 GND.n1382 GND.n1262 0.984173
R9077 GND.n1341 GND.n1277 0.984173
R9078 GND.n1349 GND.n1273 0.984173
R9079 GND.n1308 GND.n1288 0.984173
R9080 GND.n1316 GND.n1284 0.984173
R9081 GND GND.n71 0.9029
R9082 GND.n4687 GND.n4686 0.776258
R9083 GND.n4413 GND.n4412 0.776258
R9084 GND GND.n5864 0.745215
R9085 GND.n3506 GND.n2114 0.690696
R9086 GND.n4580 GND.n2123 0.690696
R9087 GND.n4530 GND.n2195 0.690696
R9088 GND.n3130 GND.n2204 0.690696
R9089 GND.n4469 GND.n4468 0.690696
R9090 GND.n4462 GND.n4461 0.690696
R9091 GND.n5855 GND.n159 0.643
R9092 GND.n1947 GND.n1572 0.643
R9093 GND.n2784 GND.n2782 0.558028
R9094 GND.n4975 GND.n798 0.52489
R9095 GND.n5546 GND.n5545 0.52489
R9096 GND.n5678 GND.n373 0.52489
R9097 GND.n4862 GND.n4861 0.52489
R9098 GND.n1761 GND.n991 0.521842
R9099 GND.n4245 GND.n4244 0.521841
R9100 GND.n5794 GND.n5793 0.512695
R9101 GND.n2817 GND.n2399 0.512695
R9102 GND.n4697 GND.n4696 0.512695
R9103 GND.n1031 GND.n999 0.512695
R9104 GND.n3283 GND.n3197 0.448671
R9105 GND.n3887 GND.n3886 0.448671
R9106 GND.n51 GND.n49 0.388379
R9107 GND.n62 GND.n60 0.388379
R9108 GND.n27 GND.n25 0.388379
R9109 GND.n38 GND.n36 0.388379
R9110 GND.n4 GND.n2 0.388379
R9111 GND.n15 GND.n13 0.388379
R9112 GND.n1464 GND.n1432 0.388379
R9113 GND.n1242 GND.n1210 0.388379
R9114 GND.n134 GND.n132 0.388379
R9115 GND.n123 GND.n121 0.388379
R9116 GND.n110 GND.n108 0.388379
R9117 GND.n99 GND.n97 0.388379
R9118 GND.n87 GND.n85 0.388379
R9119 GND.n76 GND.n74 0.388379
R9120 GND.n2500 GND.n2468 0.388379
R9121 GND.n2465 GND.n2433 0.388379
R9122 GND.n4655 GND.n1474 0.355683
R9123 GND.n4430 GND.n4429 0.355683
R9124 GND.n3516 GND.t7 0.345598
R9125 GND.n3585 GND.t2 0.345598
R9126 GND.t19 GND.n4489 0.345598
R9127 GND.n3735 GND.t3 0.345598
R9128 GND.n4428 GND.n2376 0.323822
R9129 GND.n4654 GND.n1476 0.323822
R9130 GND.n3945 GND.n2405 0.312695
R9131 GND.n3397 GND.n1190 0.312695
R9132 GND.n3306 GND.n1190 0.312695
R9133 GND.n3951 GND.n2405 0.312695
R9134 GND.n5752 GND.n306 0.294707
R9135 GND.n1074 GND.n983 0.294707
R9136 GND.n5753 GND.n5752 0.285561
R9137 GND.n4393 GND.n2423 0.285561
R9138 GND.n1074 GND.n1073 0.285561
R9139 GND.n4671 GND.n4669 0.285561
R9140 GND.n2778 GND.n2745 0.278398
R9141 GND.n2743 GND.n2710 0.278398
R9142 GND.n2708 GND.n2675 0.278398
R9143 GND.n2674 GND.n2641 0.278398
R9144 GND.n2639 GND.n2606 0.278398
R9145 GND.n2604 GND.n2571 0.278398
R9146 GND.n2569 GND.n2536 0.278398
R9147 GND.n2535 GND.n2502 0.278398
R9148 GND.n1296 GND.n1291 0.278335
R9149 GND.n1328 GND.n1281 0.278335
R9150 GND.n1329 GND.n1280 0.278335
R9151 GND.n1361 GND.n1270 0.278335
R9152 GND.n1362 GND.n1269 0.278335
R9153 GND.n1394 GND.n1259 0.278335
R9154 GND.n1395 GND.n1258 0.278335
R9155 GND.n1427 GND.n1248 0.278335
R9156 GND.n2407 GND.n2404 0.229039
R9157 GND.n2410 GND.n2407 0.229039
R9158 GND.n1188 GND.n1183 0.229039
R9159 GND.n4685 GND.n1188 0.229039
R9160 GND.n5778 GND.n5777 0.194439
R9161 GND.n1049 GND.n1026 0.194439
R9162 GND.n1300 GND.n1291 0.189894
R9163 GND.n1301 GND.n1300 0.189894
R9164 GND.n1302 GND.n1301 0.189894
R9165 GND.n1302 GND.n1289 0.189894
R9166 GND.n1306 GND.n1289 0.189894
R9167 GND.n1307 GND.n1306 0.189894
R9168 GND.n1307 GND.n1287 0.189894
R9169 GND.n1311 GND.n1287 0.189894
R9170 GND.n1312 GND.n1311 0.189894
R9171 GND.n1313 GND.n1312 0.189894
R9172 GND.n1313 GND.n1285 0.189894
R9173 GND.n1317 GND.n1285 0.189894
R9174 GND.n1318 GND.n1317 0.189894
R9175 GND.n1318 GND.n1283 0.189894
R9176 GND.n1322 GND.n1283 0.189894
R9177 GND.n1323 GND.n1322 0.189894
R9178 GND.n1324 GND.n1323 0.189894
R9179 GND.n1324 GND.n1281 0.189894
R9180 GND.n1333 GND.n1280 0.189894
R9181 GND.n1334 GND.n1333 0.189894
R9182 GND.n1335 GND.n1334 0.189894
R9183 GND.n1335 GND.n1278 0.189894
R9184 GND.n1339 GND.n1278 0.189894
R9185 GND.n1340 GND.n1339 0.189894
R9186 GND.n1340 GND.n1276 0.189894
R9187 GND.n1344 GND.n1276 0.189894
R9188 GND.n1345 GND.n1344 0.189894
R9189 GND.n1346 GND.n1345 0.189894
R9190 GND.n1346 GND.n1274 0.189894
R9191 GND.n1350 GND.n1274 0.189894
R9192 GND.n1351 GND.n1350 0.189894
R9193 GND.n1351 GND.n1272 0.189894
R9194 GND.n1355 GND.n1272 0.189894
R9195 GND.n1356 GND.n1355 0.189894
R9196 GND.n1357 GND.n1356 0.189894
R9197 GND.n1357 GND.n1270 0.189894
R9198 GND.n1366 GND.n1269 0.189894
R9199 GND.n1367 GND.n1366 0.189894
R9200 GND.n1368 GND.n1367 0.189894
R9201 GND.n1368 GND.n1267 0.189894
R9202 GND.n1372 GND.n1267 0.189894
R9203 GND.n1373 GND.n1372 0.189894
R9204 GND.n1373 GND.n1265 0.189894
R9205 GND.n1377 GND.n1265 0.189894
R9206 GND.n1378 GND.n1377 0.189894
R9207 GND.n1379 GND.n1378 0.189894
R9208 GND.n1379 GND.n1263 0.189894
R9209 GND.n1383 GND.n1263 0.189894
R9210 GND.n1384 GND.n1383 0.189894
R9211 GND.n1384 GND.n1261 0.189894
R9212 GND.n1388 GND.n1261 0.189894
R9213 GND.n1389 GND.n1388 0.189894
R9214 GND.n1390 GND.n1389 0.189894
R9215 GND.n1390 GND.n1259 0.189894
R9216 GND.n1399 GND.n1258 0.189894
R9217 GND.n1400 GND.n1399 0.189894
R9218 GND.n1401 GND.n1400 0.189894
R9219 GND.n1401 GND.n1256 0.189894
R9220 GND.n1405 GND.n1256 0.189894
R9221 GND.n1406 GND.n1405 0.189894
R9222 GND.n1406 GND.n1254 0.189894
R9223 GND.n1410 GND.n1254 0.189894
R9224 GND.n1411 GND.n1410 0.189894
R9225 GND.n1412 GND.n1411 0.189894
R9226 GND.n1412 GND.n1252 0.189894
R9227 GND.n1416 GND.n1252 0.189894
R9228 GND.n1417 GND.n1416 0.189894
R9229 GND.n1417 GND.n1250 0.189894
R9230 GND.n1421 GND.n1250 0.189894
R9231 GND.n1422 GND.n1421 0.189894
R9232 GND.n1423 GND.n1422 0.189894
R9233 GND.n1423 GND.n1248 0.189894
R9234 GND.n2774 GND.n2745 0.189894
R9235 GND.n2774 GND.n2773 0.189894
R9236 GND.n2773 GND.n2772 0.189894
R9237 GND.n2772 GND.n2747 0.189894
R9238 GND.n2767 GND.n2747 0.189894
R9239 GND.n2767 GND.n2766 0.189894
R9240 GND.n2766 GND.n2765 0.189894
R9241 GND.n2765 GND.n2749 0.189894
R9242 GND.n2760 GND.n2749 0.189894
R9243 GND.n2760 GND.n2759 0.189894
R9244 GND.n2759 GND.n2758 0.189894
R9245 GND.n2758 GND.n2751 0.189894
R9246 GND.n2754 GND.n2751 0.189894
R9247 GND.n2739 GND.n2710 0.189894
R9248 GND.n2739 GND.n2738 0.189894
R9249 GND.n2738 GND.n2737 0.189894
R9250 GND.n2737 GND.n2712 0.189894
R9251 GND.n2732 GND.n2712 0.189894
R9252 GND.n2732 GND.n2731 0.189894
R9253 GND.n2731 GND.n2730 0.189894
R9254 GND.n2730 GND.n2714 0.189894
R9255 GND.n2725 GND.n2714 0.189894
R9256 GND.n2725 GND.n2724 0.189894
R9257 GND.n2724 GND.n2723 0.189894
R9258 GND.n2723 GND.n2716 0.189894
R9259 GND.n2719 GND.n2716 0.189894
R9260 GND.n2704 GND.n2675 0.189894
R9261 GND.n2704 GND.n2703 0.189894
R9262 GND.n2703 GND.n2702 0.189894
R9263 GND.n2702 GND.n2677 0.189894
R9264 GND.n2697 GND.n2677 0.189894
R9265 GND.n2697 GND.n2696 0.189894
R9266 GND.n2696 GND.n2695 0.189894
R9267 GND.n2695 GND.n2679 0.189894
R9268 GND.n2690 GND.n2679 0.189894
R9269 GND.n2690 GND.n2689 0.189894
R9270 GND.n2689 GND.n2688 0.189894
R9271 GND.n2688 GND.n2681 0.189894
R9272 GND.n2684 GND.n2681 0.189894
R9273 GND.n2670 GND.n2641 0.189894
R9274 GND.n2670 GND.n2669 0.189894
R9275 GND.n2669 GND.n2668 0.189894
R9276 GND.n2668 GND.n2643 0.189894
R9277 GND.n2663 GND.n2643 0.189894
R9278 GND.n2663 GND.n2662 0.189894
R9279 GND.n2662 GND.n2661 0.189894
R9280 GND.n2661 GND.n2645 0.189894
R9281 GND.n2656 GND.n2645 0.189894
R9282 GND.n2656 GND.n2655 0.189894
R9283 GND.n2655 GND.n2654 0.189894
R9284 GND.n2654 GND.n2647 0.189894
R9285 GND.n2650 GND.n2647 0.189894
R9286 GND.n2615 GND.n2612 0.189894
R9287 GND.n2619 GND.n2612 0.189894
R9288 GND.n2620 GND.n2619 0.189894
R9289 GND.n2621 GND.n2620 0.189894
R9290 GND.n2621 GND.n2610 0.189894
R9291 GND.n2626 GND.n2610 0.189894
R9292 GND.n2627 GND.n2626 0.189894
R9293 GND.n2628 GND.n2627 0.189894
R9294 GND.n2628 GND.n2608 0.189894
R9295 GND.n2633 GND.n2608 0.189894
R9296 GND.n2634 GND.n2633 0.189894
R9297 GND.n2635 GND.n2634 0.189894
R9298 GND.n2635 GND.n2606 0.189894
R9299 GND.n2580 GND.n2577 0.189894
R9300 GND.n2584 GND.n2577 0.189894
R9301 GND.n2585 GND.n2584 0.189894
R9302 GND.n2586 GND.n2585 0.189894
R9303 GND.n2586 GND.n2575 0.189894
R9304 GND.n2591 GND.n2575 0.189894
R9305 GND.n2592 GND.n2591 0.189894
R9306 GND.n2593 GND.n2592 0.189894
R9307 GND.n2593 GND.n2573 0.189894
R9308 GND.n2598 GND.n2573 0.189894
R9309 GND.n2599 GND.n2598 0.189894
R9310 GND.n2600 GND.n2599 0.189894
R9311 GND.n2600 GND.n2571 0.189894
R9312 GND.n2545 GND.n2542 0.189894
R9313 GND.n2549 GND.n2542 0.189894
R9314 GND.n2550 GND.n2549 0.189894
R9315 GND.n2551 GND.n2550 0.189894
R9316 GND.n2551 GND.n2540 0.189894
R9317 GND.n2556 GND.n2540 0.189894
R9318 GND.n2557 GND.n2556 0.189894
R9319 GND.n2558 GND.n2557 0.189894
R9320 GND.n2558 GND.n2538 0.189894
R9321 GND.n2563 GND.n2538 0.189894
R9322 GND.n2564 GND.n2563 0.189894
R9323 GND.n2565 GND.n2564 0.189894
R9324 GND.n2565 GND.n2536 0.189894
R9325 GND.n2511 GND.n2508 0.189894
R9326 GND.n2515 GND.n2508 0.189894
R9327 GND.n2516 GND.n2515 0.189894
R9328 GND.n2517 GND.n2516 0.189894
R9329 GND.n2517 GND.n2506 0.189894
R9330 GND.n2522 GND.n2506 0.189894
R9331 GND.n2523 GND.n2522 0.189894
R9332 GND.n2524 GND.n2523 0.189894
R9333 GND.n2524 GND.n2504 0.189894
R9334 GND.n2529 GND.n2504 0.189894
R9335 GND.n2530 GND.n2529 0.189894
R9336 GND.n2531 GND.n2530 0.189894
R9337 GND.n2531 GND.n2502 0.189894
R9338 GND.n56 GND.n48 0.155672
R9339 GND.n67 GND.n59 0.155672
R9340 GND.n32 GND.n24 0.155672
R9341 GND.n43 GND.n35 0.155672
R9342 GND.n9 GND.n1 0.155672
R9343 GND.n20 GND.n12 0.155672
R9344 GND.n1460 GND.n1459 0.155672
R9345 GND.n1459 GND.n1435 0.155672
R9346 GND.n1452 GND.n1435 0.155672
R9347 GND.n1452 GND.n1451 0.155672
R9348 GND.n1451 GND.n1439 0.155672
R9349 GND.n1444 GND.n1439 0.155672
R9350 GND.n1222 GND.n1217 0.155672
R9351 GND.n1229 GND.n1217 0.155672
R9352 GND.n1230 GND.n1229 0.155672
R9353 GND.n1230 GND.n1213 0.155672
R9354 GND.n1237 GND.n1213 0.155672
R9355 GND.n1238 GND.n1237 0.155672
R9356 GND.n139 GND.n131 0.155672
R9357 GND.n128 GND.n120 0.155672
R9358 GND.n115 GND.n107 0.155672
R9359 GND.n104 GND.n96 0.155672
R9360 GND.n92 GND.n84 0.155672
R9361 GND.n81 GND.n73 0.155672
R9362 GND.n2496 GND.n2495 0.155672
R9363 GND.n2495 GND.n2471 0.155672
R9364 GND.n2488 GND.n2471 0.155672
R9365 GND.n2488 GND.n2487 0.155672
R9366 GND.n2487 GND.n2475 0.155672
R9367 GND.n2480 GND.n2475 0.155672
R9368 GND.n2445 GND.n2440 0.155672
R9369 GND.n2452 GND.n2440 0.155672
R9370 GND.n2453 GND.n2452 0.155672
R9371 GND.n2453 GND.n2436 0.155672
R9372 GND.n2460 GND.n2436 0.155672
R9373 GND.n2461 GND.n2460 0.155672
R9374 GND.n4976 GND.n4975 0.152939
R9375 GND.n4977 GND.n4976 0.152939
R9376 GND.n4977 GND.n792 0.152939
R9377 GND.n4985 GND.n792 0.152939
R9378 GND.n4986 GND.n4985 0.152939
R9379 GND.n4987 GND.n4986 0.152939
R9380 GND.n4987 GND.n786 0.152939
R9381 GND.n4995 GND.n786 0.152939
R9382 GND.n4996 GND.n4995 0.152939
R9383 GND.n4997 GND.n4996 0.152939
R9384 GND.n4997 GND.n780 0.152939
R9385 GND.n5005 GND.n780 0.152939
R9386 GND.n5006 GND.n5005 0.152939
R9387 GND.n5007 GND.n5006 0.152939
R9388 GND.n5007 GND.n774 0.152939
R9389 GND.n5015 GND.n774 0.152939
R9390 GND.n5016 GND.n5015 0.152939
R9391 GND.n5017 GND.n5016 0.152939
R9392 GND.n5017 GND.n768 0.152939
R9393 GND.n5025 GND.n768 0.152939
R9394 GND.n5026 GND.n5025 0.152939
R9395 GND.n5027 GND.n5026 0.152939
R9396 GND.n5027 GND.n762 0.152939
R9397 GND.n5035 GND.n762 0.152939
R9398 GND.n5036 GND.n5035 0.152939
R9399 GND.n5037 GND.n5036 0.152939
R9400 GND.n5037 GND.n756 0.152939
R9401 GND.n5045 GND.n756 0.152939
R9402 GND.n5046 GND.n5045 0.152939
R9403 GND.n5047 GND.n5046 0.152939
R9404 GND.n5047 GND.n750 0.152939
R9405 GND.n5055 GND.n750 0.152939
R9406 GND.n5056 GND.n5055 0.152939
R9407 GND.n5057 GND.n5056 0.152939
R9408 GND.n5057 GND.n744 0.152939
R9409 GND.n5065 GND.n744 0.152939
R9410 GND.n5066 GND.n5065 0.152939
R9411 GND.n5067 GND.n5066 0.152939
R9412 GND.n5067 GND.n738 0.152939
R9413 GND.n5075 GND.n738 0.152939
R9414 GND.n5076 GND.n5075 0.152939
R9415 GND.n5077 GND.n5076 0.152939
R9416 GND.n5077 GND.n732 0.152939
R9417 GND.n5085 GND.n732 0.152939
R9418 GND.n5086 GND.n5085 0.152939
R9419 GND.n5087 GND.n5086 0.152939
R9420 GND.n5087 GND.n726 0.152939
R9421 GND.n5095 GND.n726 0.152939
R9422 GND.n5096 GND.n5095 0.152939
R9423 GND.n5097 GND.n5096 0.152939
R9424 GND.n5097 GND.n720 0.152939
R9425 GND.n5105 GND.n720 0.152939
R9426 GND.n5106 GND.n5105 0.152939
R9427 GND.n5107 GND.n5106 0.152939
R9428 GND.n5107 GND.n714 0.152939
R9429 GND.n5115 GND.n714 0.152939
R9430 GND.n5116 GND.n5115 0.152939
R9431 GND.n5117 GND.n5116 0.152939
R9432 GND.n5117 GND.n708 0.152939
R9433 GND.n5125 GND.n708 0.152939
R9434 GND.n5126 GND.n5125 0.152939
R9435 GND.n5127 GND.n5126 0.152939
R9436 GND.n5127 GND.n702 0.152939
R9437 GND.n5135 GND.n702 0.152939
R9438 GND.n5136 GND.n5135 0.152939
R9439 GND.n5137 GND.n5136 0.152939
R9440 GND.n5137 GND.n696 0.152939
R9441 GND.n5145 GND.n696 0.152939
R9442 GND.n5146 GND.n5145 0.152939
R9443 GND.n5147 GND.n5146 0.152939
R9444 GND.n5147 GND.n690 0.152939
R9445 GND.n5155 GND.n690 0.152939
R9446 GND.n5156 GND.n5155 0.152939
R9447 GND.n5157 GND.n5156 0.152939
R9448 GND.n5157 GND.n684 0.152939
R9449 GND.n5165 GND.n684 0.152939
R9450 GND.n5166 GND.n5165 0.152939
R9451 GND.n5167 GND.n5166 0.152939
R9452 GND.n5167 GND.n678 0.152939
R9453 GND.n5175 GND.n678 0.152939
R9454 GND.n5176 GND.n5175 0.152939
R9455 GND.n5177 GND.n5176 0.152939
R9456 GND.n5177 GND.n672 0.152939
R9457 GND.n5185 GND.n672 0.152939
R9458 GND.n5186 GND.n5185 0.152939
R9459 GND.n5187 GND.n5186 0.152939
R9460 GND.n5187 GND.n666 0.152939
R9461 GND.n5195 GND.n666 0.152939
R9462 GND.n5196 GND.n5195 0.152939
R9463 GND.n5197 GND.n5196 0.152939
R9464 GND.n5197 GND.n660 0.152939
R9465 GND.n5205 GND.n660 0.152939
R9466 GND.n5206 GND.n5205 0.152939
R9467 GND.n5207 GND.n5206 0.152939
R9468 GND.n5207 GND.n654 0.152939
R9469 GND.n5215 GND.n654 0.152939
R9470 GND.n5216 GND.n5215 0.152939
R9471 GND.n5217 GND.n5216 0.152939
R9472 GND.n5217 GND.n648 0.152939
R9473 GND.n5225 GND.n648 0.152939
R9474 GND.n5226 GND.n5225 0.152939
R9475 GND.n5227 GND.n5226 0.152939
R9476 GND.n5227 GND.n642 0.152939
R9477 GND.n5235 GND.n642 0.152939
R9478 GND.n5236 GND.n5235 0.152939
R9479 GND.n5237 GND.n5236 0.152939
R9480 GND.n5237 GND.n636 0.152939
R9481 GND.n5245 GND.n636 0.152939
R9482 GND.n5246 GND.n5245 0.152939
R9483 GND.n5247 GND.n5246 0.152939
R9484 GND.n5247 GND.n630 0.152939
R9485 GND.n5255 GND.n630 0.152939
R9486 GND.n5256 GND.n5255 0.152939
R9487 GND.n5257 GND.n5256 0.152939
R9488 GND.n5257 GND.n624 0.152939
R9489 GND.n5265 GND.n624 0.152939
R9490 GND.n5266 GND.n5265 0.152939
R9491 GND.n5267 GND.n5266 0.152939
R9492 GND.n5267 GND.n618 0.152939
R9493 GND.n5275 GND.n618 0.152939
R9494 GND.n5276 GND.n5275 0.152939
R9495 GND.n5277 GND.n5276 0.152939
R9496 GND.n5277 GND.n612 0.152939
R9497 GND.n5285 GND.n612 0.152939
R9498 GND.n5286 GND.n5285 0.152939
R9499 GND.n5287 GND.n5286 0.152939
R9500 GND.n5287 GND.n606 0.152939
R9501 GND.n5295 GND.n606 0.152939
R9502 GND.n5296 GND.n5295 0.152939
R9503 GND.n5297 GND.n5296 0.152939
R9504 GND.n5297 GND.n600 0.152939
R9505 GND.n5305 GND.n600 0.152939
R9506 GND.n5306 GND.n5305 0.152939
R9507 GND.n5307 GND.n5306 0.152939
R9508 GND.n5307 GND.n594 0.152939
R9509 GND.n5315 GND.n594 0.152939
R9510 GND.n5316 GND.n5315 0.152939
R9511 GND.n5317 GND.n5316 0.152939
R9512 GND.n5317 GND.n588 0.152939
R9513 GND.n5325 GND.n588 0.152939
R9514 GND.n5326 GND.n5325 0.152939
R9515 GND.n5327 GND.n5326 0.152939
R9516 GND.n5327 GND.n582 0.152939
R9517 GND.n5335 GND.n582 0.152939
R9518 GND.n5336 GND.n5335 0.152939
R9519 GND.n5337 GND.n5336 0.152939
R9520 GND.n5337 GND.n576 0.152939
R9521 GND.n5345 GND.n576 0.152939
R9522 GND.n5346 GND.n5345 0.152939
R9523 GND.n5347 GND.n5346 0.152939
R9524 GND.n5347 GND.n570 0.152939
R9525 GND.n5355 GND.n570 0.152939
R9526 GND.n5356 GND.n5355 0.152939
R9527 GND.n5357 GND.n5356 0.152939
R9528 GND.n5357 GND.n564 0.152939
R9529 GND.n5365 GND.n564 0.152939
R9530 GND.n5366 GND.n5365 0.152939
R9531 GND.n5367 GND.n5366 0.152939
R9532 GND.n5367 GND.n558 0.152939
R9533 GND.n5375 GND.n558 0.152939
R9534 GND.n5376 GND.n5375 0.152939
R9535 GND.n5377 GND.n5376 0.152939
R9536 GND.n5377 GND.n552 0.152939
R9537 GND.n5385 GND.n552 0.152939
R9538 GND.n5386 GND.n5385 0.152939
R9539 GND.n5387 GND.n5386 0.152939
R9540 GND.n5387 GND.n546 0.152939
R9541 GND.n5395 GND.n546 0.152939
R9542 GND.n5396 GND.n5395 0.152939
R9543 GND.n5397 GND.n5396 0.152939
R9544 GND.n5397 GND.n540 0.152939
R9545 GND.n5405 GND.n540 0.152939
R9546 GND.n5406 GND.n5405 0.152939
R9547 GND.n5407 GND.n5406 0.152939
R9548 GND.n5407 GND.n534 0.152939
R9549 GND.n5415 GND.n534 0.152939
R9550 GND.n5416 GND.n5415 0.152939
R9551 GND.n5417 GND.n5416 0.152939
R9552 GND.n5417 GND.n528 0.152939
R9553 GND.n5425 GND.n528 0.152939
R9554 GND.n5426 GND.n5425 0.152939
R9555 GND.n5427 GND.n5426 0.152939
R9556 GND.n5427 GND.n522 0.152939
R9557 GND.n5435 GND.n522 0.152939
R9558 GND.n5436 GND.n5435 0.152939
R9559 GND.n5437 GND.n5436 0.152939
R9560 GND.n5437 GND.n516 0.152939
R9561 GND.n5445 GND.n516 0.152939
R9562 GND.n5446 GND.n5445 0.152939
R9563 GND.n5447 GND.n5446 0.152939
R9564 GND.n5447 GND.n510 0.152939
R9565 GND.n5455 GND.n510 0.152939
R9566 GND.n5456 GND.n5455 0.152939
R9567 GND.n5457 GND.n5456 0.152939
R9568 GND.n5457 GND.n504 0.152939
R9569 GND.n5465 GND.n504 0.152939
R9570 GND.n5466 GND.n5465 0.152939
R9571 GND.n5467 GND.n5466 0.152939
R9572 GND.n5467 GND.n498 0.152939
R9573 GND.n5475 GND.n498 0.152939
R9574 GND.n5476 GND.n5475 0.152939
R9575 GND.n5477 GND.n5476 0.152939
R9576 GND.n5477 GND.n492 0.152939
R9577 GND.n5485 GND.n492 0.152939
R9578 GND.n5486 GND.n5485 0.152939
R9579 GND.n5487 GND.n5486 0.152939
R9580 GND.n5487 GND.n486 0.152939
R9581 GND.n5495 GND.n486 0.152939
R9582 GND.n5496 GND.n5495 0.152939
R9583 GND.n5497 GND.n5496 0.152939
R9584 GND.n5497 GND.n480 0.152939
R9585 GND.n5505 GND.n480 0.152939
R9586 GND.n5506 GND.n5505 0.152939
R9587 GND.n5507 GND.n5506 0.152939
R9588 GND.n5507 GND.n474 0.152939
R9589 GND.n5515 GND.n474 0.152939
R9590 GND.n5516 GND.n5515 0.152939
R9591 GND.n5517 GND.n5516 0.152939
R9592 GND.n5517 GND.n468 0.152939
R9593 GND.n5525 GND.n468 0.152939
R9594 GND.n5526 GND.n5525 0.152939
R9595 GND.n5527 GND.n5526 0.152939
R9596 GND.n5527 GND.n462 0.152939
R9597 GND.n5535 GND.n462 0.152939
R9598 GND.n5536 GND.n5535 0.152939
R9599 GND.n5537 GND.n5536 0.152939
R9600 GND.n5537 GND.n456 0.152939
R9601 GND.n5545 GND.n456 0.152939
R9602 GND.n5547 GND.n5546 0.152939
R9603 GND.n5547 GND.n450 0.152939
R9604 GND.n5555 GND.n450 0.152939
R9605 GND.n5556 GND.n5555 0.152939
R9606 GND.n5557 GND.n5556 0.152939
R9607 GND.n5557 GND.n444 0.152939
R9608 GND.n5565 GND.n444 0.152939
R9609 GND.n5566 GND.n5565 0.152939
R9610 GND.n5567 GND.n5566 0.152939
R9611 GND.n5567 GND.n438 0.152939
R9612 GND.n5575 GND.n438 0.152939
R9613 GND.n5576 GND.n5575 0.152939
R9614 GND.n5577 GND.n5576 0.152939
R9615 GND.n5577 GND.n432 0.152939
R9616 GND.n5585 GND.n432 0.152939
R9617 GND.n5586 GND.n5585 0.152939
R9618 GND.n5587 GND.n5586 0.152939
R9619 GND.n5587 GND.n426 0.152939
R9620 GND.n5595 GND.n426 0.152939
R9621 GND.n5596 GND.n5595 0.152939
R9622 GND.n5597 GND.n5596 0.152939
R9623 GND.n5597 GND.n420 0.152939
R9624 GND.n5605 GND.n420 0.152939
R9625 GND.n5606 GND.n5605 0.152939
R9626 GND.n5607 GND.n5606 0.152939
R9627 GND.n5607 GND.n414 0.152939
R9628 GND.n5615 GND.n414 0.152939
R9629 GND.n5616 GND.n5615 0.152939
R9630 GND.n5617 GND.n5616 0.152939
R9631 GND.n5617 GND.n408 0.152939
R9632 GND.n5625 GND.n408 0.152939
R9633 GND.n5626 GND.n5625 0.152939
R9634 GND.n5627 GND.n5626 0.152939
R9635 GND.n5627 GND.n402 0.152939
R9636 GND.n5635 GND.n402 0.152939
R9637 GND.n5636 GND.n5635 0.152939
R9638 GND.n5637 GND.n5636 0.152939
R9639 GND.n5637 GND.n396 0.152939
R9640 GND.n5645 GND.n396 0.152939
R9641 GND.n5646 GND.n5645 0.152939
R9642 GND.n5647 GND.n5646 0.152939
R9643 GND.n5647 GND.n390 0.152939
R9644 GND.n5655 GND.n390 0.152939
R9645 GND.n5656 GND.n5655 0.152939
R9646 GND.n5657 GND.n5656 0.152939
R9647 GND.n5657 GND.n384 0.152939
R9648 GND.n5665 GND.n384 0.152939
R9649 GND.n5666 GND.n5665 0.152939
R9650 GND.n5667 GND.n5666 0.152939
R9651 GND.n5667 GND.n378 0.152939
R9652 GND.n5675 GND.n378 0.152939
R9653 GND.n5676 GND.n5675 0.152939
R9654 GND.n5677 GND.n5676 0.152939
R9655 GND.n5678 GND.n5677 0.152939
R9656 GND.n2942 GND.n2941 0.152939
R9657 GND.n2945 GND.n2942 0.152939
R9658 GND.n2946 GND.n2945 0.152939
R9659 GND.n2947 GND.n2946 0.152939
R9660 GND.n2948 GND.n2947 0.152939
R9661 GND.n2951 GND.n2948 0.152939
R9662 GND.n2952 GND.n2951 0.152939
R9663 GND.n2953 GND.n2952 0.152939
R9664 GND.n2954 GND.n2953 0.152939
R9665 GND.n4265 GND.n2954 0.152939
R9666 GND.n4266 GND.n4265 0.152939
R9667 GND.n4267 GND.n4266 0.152939
R9668 GND.n4268 GND.n4267 0.152939
R9669 GND.n4271 GND.n4268 0.152939
R9670 GND.n4272 GND.n4271 0.152939
R9671 GND.n4274 GND.n4272 0.152939
R9672 GND.n4274 GND.n4273 0.152939
R9673 GND.n4273 GND.n313 0.152939
R9674 GND.n314 GND.n313 0.152939
R9675 GND.n315 GND.n314 0.152939
R9676 GND.n321 GND.n315 0.152939
R9677 GND.n322 GND.n321 0.152939
R9678 GND.n323 GND.n322 0.152939
R9679 GND.n324 GND.n323 0.152939
R9680 GND.n325 GND.n324 0.152939
R9681 GND.n330 GND.n325 0.152939
R9682 GND.n331 GND.n330 0.152939
R9683 GND.n332 GND.n331 0.152939
R9684 GND.n333 GND.n332 0.152939
R9685 GND.n338 GND.n333 0.152939
R9686 GND.n339 GND.n338 0.152939
R9687 GND.n340 GND.n339 0.152939
R9688 GND.n341 GND.n340 0.152939
R9689 GND.n346 GND.n341 0.152939
R9690 GND.n347 GND.n346 0.152939
R9691 GND.n348 GND.n347 0.152939
R9692 GND.n349 GND.n348 0.152939
R9693 GND.n354 GND.n349 0.152939
R9694 GND.n355 GND.n354 0.152939
R9695 GND.n356 GND.n355 0.152939
R9696 GND.n357 GND.n356 0.152939
R9697 GND.n362 GND.n357 0.152939
R9698 GND.n363 GND.n362 0.152939
R9699 GND.n364 GND.n363 0.152939
R9700 GND.n365 GND.n364 0.152939
R9701 GND.n370 GND.n365 0.152939
R9702 GND.n371 GND.n370 0.152939
R9703 GND.n372 GND.n371 0.152939
R9704 GND.n373 GND.n372 0.152939
R9705 GND.n185 GND.n157 0.152939
R9706 GND.n186 GND.n185 0.152939
R9707 GND.n187 GND.n186 0.152939
R9708 GND.n205 GND.n187 0.152939
R9709 GND.n206 GND.n205 0.152939
R9710 GND.n207 GND.n206 0.152939
R9711 GND.n208 GND.n207 0.152939
R9712 GND.n226 GND.n208 0.152939
R9713 GND.n227 GND.n226 0.152939
R9714 GND.n228 GND.n227 0.152939
R9715 GND.n229 GND.n228 0.152939
R9716 GND.n246 GND.n229 0.152939
R9717 GND.n247 GND.n246 0.152939
R9718 GND.n248 GND.n247 0.152939
R9719 GND.n249 GND.n248 0.152939
R9720 GND.n267 GND.n249 0.152939
R9721 GND.n268 GND.n267 0.152939
R9722 GND.n5794 GND.n268 0.152939
R9723 GND.n4613 GND.n1474 0.152939
R9724 GND.n4613 GND.n4612 0.152939
R9725 GND.n4612 GND.n4611 0.152939
R9726 GND.n4611 GND.n2077 0.152939
R9727 GND.n2107 GND.n2077 0.152939
R9728 GND.n2108 GND.n2107 0.152939
R9729 GND.n2109 GND.n2108 0.152939
R9730 GND.n2110 GND.n2109 0.152939
R9731 GND.n2111 GND.n2110 0.152939
R9732 GND.n2128 GND.n2111 0.152939
R9733 GND.n2129 GND.n2128 0.152939
R9734 GND.n2130 GND.n2129 0.152939
R9735 GND.n2131 GND.n2130 0.152939
R9736 GND.n2148 GND.n2131 0.152939
R9737 GND.n2149 GND.n2148 0.152939
R9738 GND.n2150 GND.n2149 0.152939
R9739 GND.n2151 GND.n2150 0.152939
R9740 GND.n2168 GND.n2151 0.152939
R9741 GND.n2169 GND.n2168 0.152939
R9742 GND.n2170 GND.n2169 0.152939
R9743 GND.n2171 GND.n2170 0.152939
R9744 GND.n2186 GND.n2171 0.152939
R9745 GND.n2187 GND.n2186 0.152939
R9746 GND.n2188 GND.n2187 0.152939
R9747 GND.n2189 GND.n2188 0.152939
R9748 GND.n2206 GND.n2189 0.152939
R9749 GND.n2207 GND.n2206 0.152939
R9750 GND.n2208 GND.n2207 0.152939
R9751 GND.n2209 GND.n2208 0.152939
R9752 GND.n2238 GND.n2209 0.152939
R9753 GND.n2241 GND.n2238 0.152939
R9754 GND.n2242 GND.n2241 0.152939
R9755 GND.n2243 GND.n2242 0.152939
R9756 GND.n2244 GND.n2243 0.152939
R9757 GND.n2245 GND.n2244 0.152939
R9758 GND.n2282 GND.n2245 0.152939
R9759 GND.n2285 GND.n2282 0.152939
R9760 GND.n2286 GND.n2285 0.152939
R9761 GND.n2287 GND.n2286 0.152939
R9762 GND.n2288 GND.n2287 0.152939
R9763 GND.n2289 GND.n2288 0.152939
R9764 GND.n2331 GND.n2289 0.152939
R9765 GND.n2332 GND.n2331 0.152939
R9766 GND.n2337 GND.n2332 0.152939
R9767 GND.n2338 GND.n2337 0.152939
R9768 GND.n2339 GND.n2338 0.152939
R9769 GND.n2340 GND.n2339 0.152939
R9770 GND.n2341 GND.n2340 0.152939
R9771 GND.n3794 GND.n2341 0.152939
R9772 GND.n3796 GND.n3794 0.152939
R9773 GND.n3796 GND.n3795 0.152939
R9774 GND.n3795 GND.n2373 0.152939
R9775 GND.n4430 GND.n2373 0.152939
R9776 GND.n3212 GND.n1475 0.152939
R9777 GND.n3213 GND.n3212 0.152939
R9778 GND.n3214 GND.n3213 0.152939
R9779 GND.n3215 GND.n3214 0.152939
R9780 GND.n3216 GND.n3215 0.152939
R9781 GND.n3217 GND.n3216 0.152939
R9782 GND.n3218 GND.n3217 0.152939
R9783 GND.n3219 GND.n3218 0.152939
R9784 GND.n3220 GND.n3219 0.152939
R9785 GND.n3221 GND.n3220 0.152939
R9786 GND.n3222 GND.n3221 0.152939
R9787 GND.n3223 GND.n3222 0.152939
R9788 GND.n3224 GND.n3223 0.152939
R9789 GND.n3225 GND.n3224 0.152939
R9790 GND.n3226 GND.n3225 0.152939
R9791 GND.n3227 GND.n3226 0.152939
R9792 GND.n3228 GND.n3227 0.152939
R9793 GND.n3229 GND.n3228 0.152939
R9794 GND.n3233 GND.n3229 0.152939
R9795 GND.n3234 GND.n3233 0.152939
R9796 GND.n3235 GND.n3234 0.152939
R9797 GND.n3235 GND.n3197 0.152939
R9798 GND.n3284 GND.n3283 0.152939
R9799 GND.n3285 GND.n3284 0.152939
R9800 GND.n3285 GND.n3195 0.152939
R9801 GND.n3484 GND.n3195 0.152939
R9802 GND.n3485 GND.n3484 0.152939
R9803 GND.n3486 GND.n3485 0.152939
R9804 GND.n3486 GND.n3183 0.152939
R9805 GND.n3510 GND.n3183 0.152939
R9806 GND.n3511 GND.n3510 0.152939
R9807 GND.n3512 GND.n3511 0.152939
R9808 GND.n3512 GND.n3177 0.152939
R9809 GND.n3557 GND.n3177 0.152939
R9810 GND.n3558 GND.n3557 0.152939
R9811 GND.n3560 GND.n3558 0.152939
R9812 GND.n3560 GND.n3559 0.152939
R9813 GND.n3559 GND.n3161 0.152939
R9814 GND.n3162 GND.n3161 0.152939
R9815 GND.n3163 GND.n3162 0.152939
R9816 GND.n3164 GND.n3163 0.152939
R9817 GND.n3165 GND.n3164 0.152939
R9818 GND.n3166 GND.n3165 0.152939
R9819 GND.n3167 GND.n3166 0.152939
R9820 GND.n3167 GND.n3135 0.152939
R9821 GND.n3637 GND.n3135 0.152939
R9822 GND.n3638 GND.n3637 0.152939
R9823 GND.n3639 GND.n3638 0.152939
R9824 GND.n3640 GND.n3639 0.152939
R9825 GND.n3641 GND.n3640 0.152939
R9826 GND.n3642 GND.n3641 0.152939
R9827 GND.n3643 GND.n3642 0.152939
R9828 GND.n3645 GND.n3643 0.152939
R9829 GND.n3647 GND.n3645 0.152939
R9830 GND.n3647 GND.n3646 0.152939
R9831 GND.n3646 GND.n3121 0.152939
R9832 GND.n3121 GND.n3119 0.152939
R9833 GND.n3704 GND.n3119 0.152939
R9834 GND.n3705 GND.n3704 0.152939
R9835 GND.n3707 GND.n3705 0.152939
R9836 GND.n3707 GND.n3706 0.152939
R9837 GND.n3706 GND.n3107 0.152939
R9838 GND.n3751 GND.n3107 0.152939
R9839 GND.n3752 GND.n3751 0.152939
R9840 GND.n3753 GND.n3752 0.152939
R9841 GND.n3753 GND.n3103 0.152939
R9842 GND.n3759 GND.n3103 0.152939
R9843 GND.n3760 GND.n3759 0.152939
R9844 GND.n3761 GND.n3760 0.152939
R9845 GND.n3762 GND.n3761 0.152939
R9846 GND.n3763 GND.n3762 0.152939
R9847 GND.n3763 GND.n3093 0.152939
R9848 GND.n3803 GND.n3093 0.152939
R9849 GND.n3804 GND.n3803 0.152939
R9850 GND.n3887 GND.n3804 0.152939
R9851 GND.n3877 GND.n2374 0.152939
R9852 GND.n3877 GND.n3876 0.152939
R9853 GND.n3876 GND.n3875 0.152939
R9854 GND.n3875 GND.n3820 0.152939
R9855 GND.n3821 GND.n3820 0.152939
R9856 GND.n3822 GND.n3821 0.152939
R9857 GND.n3823 GND.n3822 0.152939
R9858 GND.n3824 GND.n3823 0.152939
R9859 GND.n3825 GND.n3824 0.152939
R9860 GND.n3826 GND.n3825 0.152939
R9861 GND.n3827 GND.n3826 0.152939
R9862 GND.n3828 GND.n3827 0.152939
R9863 GND.n3829 GND.n3828 0.152939
R9864 GND.n3830 GND.n3829 0.152939
R9865 GND.n3831 GND.n3830 0.152939
R9866 GND.n3832 GND.n3831 0.152939
R9867 GND.n3833 GND.n3832 0.152939
R9868 GND.n3834 GND.n3833 0.152939
R9869 GND.n3839 GND.n3834 0.152939
R9870 GND.n3839 GND.n3838 0.152939
R9871 GND.n3838 GND.n3805 0.152939
R9872 GND.n3886 GND.n3805 0.152939
R9873 GND.n2996 GND.n2376 0.152939
R9874 GND.n2996 GND.n2992 0.152939
R9875 GND.n3002 GND.n2992 0.152939
R9876 GND.n3003 GND.n3002 0.152939
R9877 GND.n3004 GND.n3003 0.152939
R9878 GND.n3004 GND.n2988 0.152939
R9879 GND.n4088 GND.n2988 0.152939
R9880 GND.n4089 GND.n4088 0.152939
R9881 GND.n4090 GND.n4089 0.152939
R9882 GND.n4090 GND.n2984 0.152939
R9883 GND.n4103 GND.n2984 0.152939
R9884 GND.n4104 GND.n4103 0.152939
R9885 GND.n4105 GND.n4104 0.152939
R9886 GND.n4105 GND.n2980 0.152939
R9887 GND.n4118 GND.n2980 0.152939
R9888 GND.n4119 GND.n4118 0.152939
R9889 GND.n4120 GND.n4119 0.152939
R9890 GND.n4121 GND.n4120 0.152939
R9891 GND.n4122 GND.n4121 0.152939
R9892 GND.n4123 GND.n4122 0.152939
R9893 GND.n4124 GND.n4123 0.152939
R9894 GND.n4125 GND.n4124 0.152939
R9895 GND.n4125 GND.n143 0.152939
R9896 GND.n5862 GND.n144 0.152939
R9897 GND.n4161 GND.n144 0.152939
R9898 GND.n4162 GND.n4161 0.152939
R9899 GND.n4162 GND.n2975 0.152939
R9900 GND.n4174 GND.n2975 0.152939
R9901 GND.n4175 GND.n4174 0.152939
R9902 GND.n4176 GND.n4175 0.152939
R9903 GND.n4176 GND.n2970 0.152939
R9904 GND.n4188 GND.n2970 0.152939
R9905 GND.n4189 GND.n4188 0.152939
R9906 GND.n4190 GND.n4189 0.152939
R9907 GND.n4190 GND.n2965 0.152939
R9908 GND.n4202 GND.n2965 0.152939
R9909 GND.n4203 GND.n4202 0.152939
R9910 GND.n4205 GND.n4203 0.152939
R9911 GND.n4205 GND.n4204 0.152939
R9912 GND.n4204 GND.n2958 0.152939
R9913 GND.n2959 GND.n2958 0.152939
R9914 GND.n2960 GND.n2959 0.152939
R9915 GND.n4215 GND.n2960 0.152939
R9916 GND.n4216 GND.n4215 0.152939
R9917 GND.n4217 GND.n4216 0.152939
R9918 GND.n4245 GND.n4217 0.152939
R9919 GND.n4227 GND.n306 0.152939
R9920 GND.n4228 GND.n4227 0.152939
R9921 GND.n4228 GND.n4223 0.152939
R9922 GND.n4236 GND.n4223 0.152939
R9923 GND.n4237 GND.n4236 0.152939
R9924 GND.n4238 GND.n4237 0.152939
R9925 GND.n4238 GND.n4218 0.152939
R9926 GND.n4244 GND.n4218 0.152939
R9927 GND.n5793 GND.n269 0.152939
R9928 GND.n288 GND.n269 0.152939
R9929 GND.n289 GND.n288 0.152939
R9930 GND.n290 GND.n289 0.152939
R9931 GND.n291 GND.n290 0.152939
R9932 GND.n292 GND.n291 0.152939
R9933 GND.n293 GND.n292 0.152939
R9934 GND.n294 GND.n293 0.152939
R9935 GND.n295 GND.n294 0.152939
R9936 GND.n296 GND.n295 0.152939
R9937 GND.n297 GND.n296 0.152939
R9938 GND.n298 GND.n297 0.152939
R9939 GND.n299 GND.n298 0.152939
R9940 GND.n300 GND.n299 0.152939
R9941 GND.n301 GND.n300 0.152939
R9942 GND.n302 GND.n301 0.152939
R9943 GND.n5754 GND.n302 0.152939
R9944 GND.n5754 GND.n5753 0.152939
R9945 GND.n2400 GND.n2399 0.152939
R9946 GND.n2401 GND.n2400 0.152939
R9947 GND.n2402 GND.n2401 0.152939
R9948 GND.n2403 GND.n2402 0.152939
R9949 GND.n2404 GND.n2403 0.152939
R9950 GND.n2411 GND.n2410 0.152939
R9951 GND.n2412 GND.n2411 0.152939
R9952 GND.n2413 GND.n2412 0.152939
R9953 GND.n2414 GND.n2413 0.152939
R9954 GND.n2415 GND.n2414 0.152939
R9955 GND.n2416 GND.n2415 0.152939
R9956 GND.n2417 GND.n2416 0.152939
R9957 GND.n4395 GND.n2417 0.152939
R9958 GND.n4395 GND.n4394 0.152939
R9959 GND.n4394 GND.n4393 0.152939
R9960 GND.n2818 GND.n2817 0.152939
R9961 GND.n2819 GND.n2818 0.152939
R9962 GND.n2820 GND.n2819 0.152939
R9963 GND.n2821 GND.n2820 0.152939
R9964 GND.n2841 GND.n2821 0.152939
R9965 GND.n2842 GND.n2841 0.152939
R9966 GND.n2843 GND.n2842 0.152939
R9967 GND.n2844 GND.n2843 0.152939
R9968 GND.n2862 GND.n2844 0.152939
R9969 GND.n2863 GND.n2862 0.152939
R9970 GND.n2864 GND.n2863 0.152939
R9971 GND.n2865 GND.n2864 0.152939
R9972 GND.n2883 GND.n2865 0.152939
R9973 GND.n2884 GND.n2883 0.152939
R9974 GND.n2885 GND.n2884 0.152939
R9975 GND.n2886 GND.n2885 0.152939
R9976 GND.n2887 GND.n2886 0.152939
R9977 GND.n2887 GND.n158 0.152939
R9978 GND.n1619 GND.n1618 0.152939
R9979 GND.n1620 GND.n1619 0.152939
R9980 GND.n1621 GND.n1620 0.152939
R9981 GND.n1624 GND.n1621 0.152939
R9982 GND.n1625 GND.n1624 0.152939
R9983 GND.n1626 GND.n1625 0.152939
R9984 GND.n1627 GND.n1626 0.152939
R9985 GND.n1630 GND.n1627 0.152939
R9986 GND.n1631 GND.n1630 0.152939
R9987 GND.n1632 GND.n1631 0.152939
R9988 GND.n1633 GND.n1632 0.152939
R9989 GND.n1636 GND.n1633 0.152939
R9990 GND.n1637 GND.n1636 0.152939
R9991 GND.n1638 GND.n1637 0.152939
R9992 GND.n1639 GND.n1638 0.152939
R9993 GND.n1641 GND.n1639 0.152939
R9994 GND.n1641 GND.n1640 0.152939
R9995 GND.n1640 GND.n1488 0.152939
R9996 GND.n2046 GND.n1488 0.152939
R9997 GND.n2047 GND.n2046 0.152939
R9998 GND.n2048 GND.n2047 0.152939
R9999 GND.n2049 GND.n2048 0.152939
R10000 GND.n2050 GND.n2049 0.152939
R10001 GND.n2055 GND.n2050 0.152939
R10002 GND.n2056 GND.n2055 0.152939
R10003 GND.n2057 GND.n2056 0.152939
R10004 GND.n2058 GND.n2057 0.152939
R10005 GND.n3470 GND.n2058 0.152939
R10006 GND.n3471 GND.n3470 0.152939
R10007 GND.n3473 GND.n3471 0.152939
R10008 GND.n3473 GND.n3472 0.152939
R10009 GND.n3472 GND.n2094 0.152939
R10010 GND.n2095 GND.n2094 0.152939
R10011 GND.n2096 GND.n2095 0.152939
R10012 GND.n3533 GND.n2096 0.152939
R10013 GND.n3534 GND.n3533 0.152939
R10014 GND.n3534 GND.n3531 0.152939
R10015 GND.n3540 GND.n3531 0.152939
R10016 GND.n3541 GND.n3540 0.152939
R10017 GND.n3542 GND.n3541 0.152939
R10018 GND.n3543 GND.n3542 0.152939
R10019 GND.n3544 GND.n3543 0.152939
R10020 GND.n3546 GND.n3544 0.152939
R10021 GND.n3546 GND.n3545 0.152939
R10022 GND.n3545 GND.n3152 0.152939
R10023 GND.n3590 GND.n3152 0.152939
R10024 GND.n3591 GND.n3590 0.152939
R10025 GND.n3592 GND.n3591 0.152939
R10026 GND.n3592 GND.n3142 0.152939
R10027 GND.n3616 GND.n3142 0.152939
R10028 GND.n3617 GND.n3616 0.152939
R10029 GND.n3618 GND.n3617 0.152939
R10030 GND.n3619 GND.n3618 0.152939
R10031 GND.n3620 GND.n3619 0.152939
R10032 GND.n3622 GND.n3620 0.152939
R10033 GND.n3622 GND.n3621 0.152939
R10034 GND.n3621 GND.n2218 0.152939
R10035 GND.n2219 GND.n2218 0.152939
R10036 GND.n2220 GND.n2219 0.152939
R10037 GND.n2263 GND.n2220 0.152939
R10038 GND.n2264 GND.n2263 0.152939
R10039 GND.n2269 GND.n2264 0.152939
R10040 GND.n2270 GND.n2269 0.152939
R10041 GND.n2271 GND.n2270 0.152939
R10042 GND.n2272 GND.n2271 0.152939
R10043 GND.n2273 GND.n2272 0.152939
R10044 GND.n2306 GND.n2273 0.152939
R10045 GND.n2309 GND.n2306 0.152939
R10046 GND.n2310 GND.n2309 0.152939
R10047 GND.n2311 GND.n2310 0.152939
R10048 GND.n2312 GND.n2311 0.152939
R10049 GND.n2313 GND.n2312 0.152939
R10050 GND.n2350 GND.n2313 0.152939
R10051 GND.n2353 GND.n2350 0.152939
R10052 GND.n2354 GND.n2353 0.152939
R10053 GND.n2355 GND.n2354 0.152939
R10054 GND.n2356 GND.n2355 0.152939
R10055 GND.n2357 GND.n2356 0.152939
R10056 GND.n3024 GND.n2357 0.152939
R10057 GND.n3025 GND.n3024 0.152939
R10058 GND.n4009 GND.n3025 0.152939
R10059 GND.n4010 GND.n4009 0.152939
R10060 GND.n4011 GND.n4010 0.152939
R10061 GND.n4011 GND.n3018 0.152939
R10062 GND.n4020 GND.n3018 0.152939
R10063 GND.n4021 GND.n4020 0.152939
R10064 GND.n4022 GND.n4021 0.152939
R10065 GND.n4022 GND.n3014 0.152939
R10066 GND.n4028 GND.n3014 0.152939
R10067 GND.n4029 GND.n4028 0.152939
R10068 GND.n4030 GND.n4029 0.152939
R10069 GND.n4030 GND.n3010 0.152939
R10070 GND.n4036 GND.n3010 0.152939
R10071 GND.n4037 GND.n4036 0.152939
R10072 GND.n4038 GND.n4037 0.152939
R10073 GND.n4039 GND.n4038 0.152939
R10074 GND.n4040 GND.n4039 0.152939
R10075 GND.n4043 GND.n4040 0.152939
R10076 GND.n4044 GND.n4043 0.152939
R10077 GND.n4045 GND.n4044 0.152939
R10078 GND.n4046 GND.n4045 0.152939
R10079 GND.n4049 GND.n4046 0.152939
R10080 GND.n4050 GND.n4049 0.152939
R10081 GND.n4051 GND.n4050 0.152939
R10082 GND.n4052 GND.n4051 0.152939
R10083 GND.n4054 GND.n4052 0.152939
R10084 GND.n4056 GND.n4054 0.152939
R10085 GND.n4056 GND.n4055 0.152939
R10086 GND.n1949 GND.n1948 0.152939
R10087 GND.n1949 GND.n1549 0.152939
R10088 GND.n1971 GND.n1549 0.152939
R10089 GND.n1972 GND.n1971 0.152939
R10090 GND.n1973 GND.n1972 0.152939
R10091 GND.n1974 GND.n1973 0.152939
R10092 GND.n1974 GND.n1526 0.152939
R10093 GND.n1995 GND.n1526 0.152939
R10094 GND.n1996 GND.n1995 0.152939
R10095 GND.n1997 GND.n1996 0.152939
R10096 GND.n1998 GND.n1997 0.152939
R10097 GND.n1998 GND.n1503 0.152939
R10098 GND.n2029 GND.n1503 0.152939
R10099 GND.n2030 GND.n2029 0.152939
R10100 GND.n2031 GND.n2030 0.152939
R10101 GND.n2032 GND.n2031 0.152939
R10102 GND.n2032 GND.n1178 0.152939
R10103 GND.n4697 GND.n1178 0.152939
R10104 GND.n1036 GND.n1031 0.152939
R10105 GND.n1037 GND.n1036 0.152939
R10106 GND.n1038 GND.n1037 0.152939
R10107 GND.n1038 GND.n1029 0.152939
R10108 GND.n1046 GND.n1029 0.152939
R10109 GND.n1047 GND.n1046 0.152939
R10110 GND.n1048 GND.n1047 0.152939
R10111 GND.n1048 GND.n1027 0.152939
R10112 GND.n1027 GND.n1023 0.152939
R10113 GND.n1057 GND.n1023 0.152939
R10114 GND.n1058 GND.n1057 0.152939
R10115 GND.n1059 GND.n1058 0.152939
R10116 GND.n1059 GND.n1021 0.152939
R10117 GND.n1067 GND.n1021 0.152939
R10118 GND.n1068 GND.n1067 0.152939
R10119 GND.n1069 GND.n1068 0.152939
R10120 GND.n1069 GND.n1014 0.152939
R10121 GND.n1073 GND.n1014 0.152939
R10122 GND.n1000 GND.n999 0.152939
R10123 GND.n1001 GND.n1000 0.152939
R10124 GND.n1730 GND.n1001 0.152939
R10125 GND.n1731 GND.n1730 0.152939
R10126 GND.n1825 GND.n1731 0.152939
R10127 GND.n1826 GND.n1825 0.152939
R10128 GND.n1827 GND.n1826 0.152939
R10129 GND.n1828 GND.n1827 0.152939
R10130 GND.n1828 GND.n1707 0.152939
R10131 GND.n1850 GND.n1707 0.152939
R10132 GND.n1851 GND.n1850 0.152939
R10133 GND.n1852 GND.n1851 0.152939
R10134 GND.n1853 GND.n1852 0.152939
R10135 GND.n1853 GND.n1685 0.152939
R10136 GND.n1875 GND.n1685 0.152939
R10137 GND.n1876 GND.n1875 0.152939
R10138 GND.n1877 GND.n1876 0.152939
R10139 GND.n1877 GND.n1571 0.152939
R10140 GND.n4861 GND.n908 0.152939
R10141 GND.n913 GND.n908 0.152939
R10142 GND.n914 GND.n913 0.152939
R10143 GND.n915 GND.n914 0.152939
R10144 GND.n920 GND.n915 0.152939
R10145 GND.n921 GND.n920 0.152939
R10146 GND.n922 GND.n921 0.152939
R10147 GND.n923 GND.n922 0.152939
R10148 GND.n928 GND.n923 0.152939
R10149 GND.n929 GND.n928 0.152939
R10150 GND.n930 GND.n929 0.152939
R10151 GND.n931 GND.n930 0.152939
R10152 GND.n936 GND.n931 0.152939
R10153 GND.n937 GND.n936 0.152939
R10154 GND.n938 GND.n937 0.152939
R10155 GND.n939 GND.n938 0.152939
R10156 GND.n944 GND.n939 0.152939
R10157 GND.n945 GND.n944 0.152939
R10158 GND.n946 GND.n945 0.152939
R10159 GND.n947 GND.n946 0.152939
R10160 GND.n952 GND.n947 0.152939
R10161 GND.n953 GND.n952 0.152939
R10162 GND.n954 GND.n953 0.152939
R10163 GND.n955 GND.n954 0.152939
R10164 GND.n960 GND.n955 0.152939
R10165 GND.n961 GND.n960 0.152939
R10166 GND.n962 GND.n961 0.152939
R10167 GND.n963 GND.n962 0.152939
R10168 GND.n1745 GND.n963 0.152939
R10169 GND.n1746 GND.n1745 0.152939
R10170 GND.n1751 GND.n1746 0.152939
R10171 GND.n1752 GND.n1751 0.152939
R10172 GND.n1753 GND.n1752 0.152939
R10173 GND.n1753 GND.n1741 0.152939
R10174 GND.n1775 GND.n1741 0.152939
R10175 GND.n1776 GND.n1775 0.152939
R10176 GND.n1777 GND.n1776 0.152939
R10177 GND.n1778 GND.n1777 0.152939
R10178 GND.n1779 GND.n1778 0.152939
R10179 GND.n1782 GND.n1779 0.152939
R10180 GND.n1783 GND.n1782 0.152939
R10181 GND.n1784 GND.n1783 0.152939
R10182 GND.n1785 GND.n1784 0.152939
R10183 GND.n1788 GND.n1785 0.152939
R10184 GND.n1789 GND.n1788 0.152939
R10185 GND.n1790 GND.n1789 0.152939
R10186 GND.n1791 GND.n1790 0.152939
R10187 GND.n1794 GND.n1791 0.152939
R10188 GND.n1795 GND.n1794 0.152939
R10189 GND.n803 GND.n798 0.152939
R10190 GND.n804 GND.n803 0.152939
R10191 GND.n805 GND.n804 0.152939
R10192 GND.n810 GND.n805 0.152939
R10193 GND.n811 GND.n810 0.152939
R10194 GND.n812 GND.n811 0.152939
R10195 GND.n813 GND.n812 0.152939
R10196 GND.n818 GND.n813 0.152939
R10197 GND.n819 GND.n818 0.152939
R10198 GND.n820 GND.n819 0.152939
R10199 GND.n821 GND.n820 0.152939
R10200 GND.n826 GND.n821 0.152939
R10201 GND.n827 GND.n826 0.152939
R10202 GND.n828 GND.n827 0.152939
R10203 GND.n829 GND.n828 0.152939
R10204 GND.n834 GND.n829 0.152939
R10205 GND.n835 GND.n834 0.152939
R10206 GND.n836 GND.n835 0.152939
R10207 GND.n837 GND.n836 0.152939
R10208 GND.n842 GND.n837 0.152939
R10209 GND.n843 GND.n842 0.152939
R10210 GND.n844 GND.n843 0.152939
R10211 GND.n845 GND.n844 0.152939
R10212 GND.n850 GND.n845 0.152939
R10213 GND.n851 GND.n850 0.152939
R10214 GND.n852 GND.n851 0.152939
R10215 GND.n853 GND.n852 0.152939
R10216 GND.n858 GND.n853 0.152939
R10217 GND.n859 GND.n858 0.152939
R10218 GND.n860 GND.n859 0.152939
R10219 GND.n861 GND.n860 0.152939
R10220 GND.n866 GND.n861 0.152939
R10221 GND.n867 GND.n866 0.152939
R10222 GND.n868 GND.n867 0.152939
R10223 GND.n869 GND.n868 0.152939
R10224 GND.n874 GND.n869 0.152939
R10225 GND.n875 GND.n874 0.152939
R10226 GND.n876 GND.n875 0.152939
R10227 GND.n877 GND.n876 0.152939
R10228 GND.n882 GND.n877 0.152939
R10229 GND.n883 GND.n882 0.152939
R10230 GND.n884 GND.n883 0.152939
R10231 GND.n885 GND.n884 0.152939
R10232 GND.n890 GND.n885 0.152939
R10233 GND.n891 GND.n890 0.152939
R10234 GND.n892 GND.n891 0.152939
R10235 GND.n893 GND.n892 0.152939
R10236 GND.n898 GND.n893 0.152939
R10237 GND.n899 GND.n898 0.152939
R10238 GND.n900 GND.n899 0.152939
R10239 GND.n901 GND.n900 0.152939
R10240 GND.n906 GND.n901 0.152939
R10241 GND.n907 GND.n906 0.152939
R10242 GND.n4862 GND.n907 0.152939
R10243 GND.n1898 GND.n1670 0.152939
R10244 GND.n1899 GND.n1898 0.152939
R10245 GND.n1900 GND.n1899 0.152939
R10246 GND.n1900 GND.n1561 0.152939
R10247 GND.n1956 GND.n1561 0.152939
R10248 GND.n1957 GND.n1956 0.152939
R10249 GND.n1959 GND.n1957 0.152939
R10250 GND.n1959 GND.n1958 0.152939
R10251 GND.n1958 GND.n1539 0.152939
R10252 GND.n1981 GND.n1539 0.152939
R10253 GND.n1982 GND.n1981 0.152939
R10254 GND.n1984 GND.n1982 0.152939
R10255 GND.n1984 GND.n1983 0.152939
R10256 GND.n1983 GND.n1515 0.152939
R10257 GND.n2005 GND.n1515 0.152939
R10258 GND.n2006 GND.n2005 0.152939
R10259 GND.n2020 GND.n2006 0.152939
R10260 GND.n2020 GND.n2019 0.152939
R10261 GND.n2019 GND.n2018 0.152939
R10262 GND.n2018 GND.n2007 0.152939
R10263 GND.n2014 GND.n2007 0.152939
R10264 GND.n2014 GND.n2013 0.152939
R10265 GND.n2013 GND.n1476 0.152939
R10266 GND.n4696 GND.n1179 0.152939
R10267 GND.n4692 GND.n1179 0.152939
R10268 GND.n4692 GND.n4691 0.152939
R10269 GND.n4691 GND.n4690 0.152939
R10270 GND.n4690 GND.n1183 0.152939
R10271 GND.n4685 GND.n4684 0.152939
R10272 GND.n4684 GND.n4683 0.152939
R10273 GND.n4683 GND.n1193 0.152939
R10274 GND.n4679 GND.n1193 0.152939
R10275 GND.n4679 GND.n4678 0.152939
R10276 GND.n4678 GND.n4677 0.152939
R10277 GND.n4677 GND.n1198 0.152939
R10278 GND.n4673 GND.n1198 0.152939
R10279 GND.n4673 GND.n4672 0.152939
R10280 GND.n4672 GND.n4671 0.152939
R10281 GND.n4796 GND.n983 0.152939
R10282 GND.n4796 GND.n4795 0.152939
R10283 GND.n4795 GND.n4794 0.152939
R10284 GND.n4794 GND.n985 0.152939
R10285 GND.n4790 GND.n985 0.152939
R10286 GND.n4790 GND.n4789 0.152939
R10287 GND.n4789 GND.n4788 0.152939
R10288 GND.n4788 GND.n991 0.152939
R10289 GND.n1762 GND.n1761 0.152939
R10290 GND.n1765 GND.n1762 0.152939
R10291 GND.n1766 GND.n1765 0.152939
R10292 GND.n1768 GND.n1766 0.152939
R10293 GND.n1768 GND.n1767 0.152939
R10294 GND.n1767 GND.n1719 0.152939
R10295 GND.n1835 GND.n1719 0.152939
R10296 GND.n1836 GND.n1835 0.152939
R10297 GND.n1838 GND.n1836 0.152939
R10298 GND.n1838 GND.n1837 0.152939
R10299 GND.n1837 GND.n1696 0.152939
R10300 GND.n1860 GND.n1696 0.152939
R10301 GND.n1861 GND.n1860 0.152939
R10302 GND.n1863 GND.n1861 0.152939
R10303 GND.n1863 GND.n1862 0.152939
R10304 GND.n1862 GND.n1674 0.152939
R10305 GND.n1883 GND.n1674 0.152939
R10306 GND.n1884 GND.n1883 0.152939
R10307 GND.n1885 GND.n1884 0.152939
R10308 GND.n1885 GND.n1672 0.152939
R10309 GND.n1891 GND.n1672 0.152939
R10310 GND.n1892 GND.n1891 0.152939
R10311 GND.n1894 GND.n1892 0.152939
R10312 GND.n2941 GND.n159 0.137695
R10313 GND.n1795 GND.n1572 0.137695
R10314 GND.n2428 GND.n2423 0.0966879
R10315 GND.n4669 GND.n4668 0.0966879
R10316 GND.n4655 GND.n1475 0.0934878
R10317 GND.n4429 GND.n2374 0.0934878
R10318 GND.n5855 GND.n157 0.0767195
R10319 GND.n5855 GND.n158 0.0767195
R10320 GND.n1948 GND.n1947 0.0767195
R10321 GND.n1947 GND.n1571 0.0767195
R10322 GND.n5863 GND.n143 0.0695946
R10323 GND.n5863 GND.n5862 0.0695946
R10324 GND.n1893 GND.n1670 0.0695946
R10325 GND.n1894 GND.n1893 0.0695946
R10326 GND.n2804 GND.n2423 0.0511114
R10327 GND.n5752 GND.n5751 0.0511114
R10328 GND.n1076 GND.n1074 0.0511114
R10329 GND.n4669 GND.n1167 0.0511114
R10330 GND.n4385 GND.n2804 0.0344674
R10331 GND.n4385 GND.n2806 0.0344674
R10332 GND.n2831 GND.n2806 0.0344674
R10333 GND.n2832 GND.n2831 0.0344674
R10334 GND.n2833 GND.n2832 0.0344674
R10335 GND.n2834 GND.n2833 0.0344674
R10336 GND.n4082 GND.n2834 0.0344674
R10337 GND.n4082 GND.n2852 0.0344674
R10338 GND.n2853 GND.n2852 0.0344674
R10339 GND.n2854 GND.n2853 0.0344674
R10340 GND.n4097 GND.n2854 0.0344674
R10341 GND.n4097 GND.n2873 0.0344674
R10342 GND.n2874 GND.n2873 0.0344674
R10343 GND.n2875 GND.n2874 0.0344674
R10344 GND.n4112 GND.n2875 0.0344674
R10345 GND.n4112 GND.n2895 0.0344674
R10346 GND.n2896 GND.n2895 0.0344674
R10347 GND.n2897 GND.n2896 0.0344674
R10348 GND.n4140 GND.n2897 0.0344674
R10349 GND.n4143 GND.n4140 0.0344674
R10350 GND.n4144 GND.n4143 0.0344674
R10351 GND.n4144 GND.n2922 0.0344674
R10352 GND.n2923 GND.n2922 0.0344674
R10353 GND.n2924 GND.n2923 0.0344674
R10354 GND.n2925 GND.n2924 0.0344674
R10355 GND.n4155 GND.n2925 0.0344674
R10356 GND.n4156 GND.n4155 0.0344674
R10357 GND.n4156 GND.n175 0.0344674
R10358 GND.n176 GND.n175 0.0344674
R10359 GND.n177 GND.n176 0.0344674
R10360 GND.n2973 GND.n177 0.0344674
R10361 GND.n2973 GND.n195 0.0344674
R10362 GND.n196 GND.n195 0.0344674
R10363 GND.n197 GND.n196 0.0344674
R10364 GND.n2968 GND.n197 0.0344674
R10365 GND.n2968 GND.n216 0.0344674
R10366 GND.n217 GND.n216 0.0344674
R10367 GND.n218 GND.n217 0.0344674
R10368 GND.n2963 GND.n218 0.0344674
R10369 GND.n2963 GND.n237 0.0344674
R10370 GND.n238 GND.n237 0.0344674
R10371 GND.n239 GND.n238 0.0344674
R10372 GND.n4214 GND.n239 0.0344674
R10373 GND.n4214 GND.n257 0.0344674
R10374 GND.n258 GND.n257 0.0344674
R10375 GND.n259 GND.n258 0.0344674
R10376 GND.n5751 GND.n259 0.0344674
R10377 GND.n1076 GND.n1012 0.0344674
R10378 GND.n4770 GND.n1012 0.0344674
R10379 GND.n4770 GND.n1013 0.0344674
R10380 GND.n4766 GND.n1013 0.0344674
R10381 GND.n4766 GND.n4765 0.0344674
R10382 GND.n4765 GND.n4764 0.0344674
R10383 GND.n4764 GND.n1087 0.0344674
R10384 GND.n4760 GND.n1087 0.0344674
R10385 GND.n4760 GND.n4759 0.0344674
R10386 GND.n4759 GND.n4758 0.0344674
R10387 GND.n4758 GND.n1095 0.0344674
R10388 GND.n4754 GND.n1095 0.0344674
R10389 GND.n4754 GND.n4753 0.0344674
R10390 GND.n4753 GND.n4752 0.0344674
R10391 GND.n4752 GND.n1103 0.0344674
R10392 GND.n4748 GND.n1103 0.0344674
R10393 GND.n4748 GND.n4747 0.0344674
R10394 GND.n4747 GND.n4746 0.0344674
R10395 GND.n4746 GND.n1111 0.0344674
R10396 GND.n4742 GND.n1111 0.0344674
R10397 GND.n4742 GND.n4741 0.0344674
R10398 GND.n4741 GND.n4740 0.0344674
R10399 GND.n4740 GND.n1119 0.0344674
R10400 GND.n4736 GND.n1119 0.0344674
R10401 GND.n4736 GND.n4735 0.0344674
R10402 GND.n4735 GND.n4734 0.0344674
R10403 GND.n4734 GND.n1127 0.0344674
R10404 GND.n4730 GND.n1127 0.0344674
R10405 GND.n4730 GND.n4729 0.0344674
R10406 GND.n4729 GND.n4728 0.0344674
R10407 GND.n4728 GND.n1135 0.0344674
R10408 GND.n4724 GND.n1135 0.0344674
R10409 GND.n4724 GND.n4723 0.0344674
R10410 GND.n4723 GND.n4722 0.0344674
R10411 GND.n4722 GND.n1143 0.0344674
R10412 GND.n4718 GND.n1143 0.0344674
R10413 GND.n4718 GND.n4717 0.0344674
R10414 GND.n4717 GND.n4716 0.0344674
R10415 GND.n4716 GND.n1151 0.0344674
R10416 GND.n4712 GND.n1151 0.0344674
R10417 GND.n4712 GND.n4711 0.0344674
R10418 GND.n4711 GND.n4710 0.0344674
R10419 GND.n4710 GND.n1159 0.0344674
R10420 GND.n4706 GND.n1159 0.0344674
R10421 GND.n4706 GND.n4705 0.0344674
R10422 GND.n4705 GND.n4704 0.0344674
R10423 GND.n4704 GND.n1167 0.0344674
R10424 GND.n2429 GND.n2428 0.0226631
R10425 GND.n2430 GND.n2429 0.0226631
R10426 GND.n2431 GND.n2430 0.0226631
R10427 GND.n2432 GND.n2431 0.0226631
R10428 GND.n2788 GND.n2787 0.0226631
R10429 GND.n2788 GND.n2375 0.0226631
R10430 GND.n4668 GND.n1205 0.0226631
R10431 GND.n4664 GND.n1205 0.0226631
R10432 GND.n4664 GND.n4663 0.0226631
R10433 GND.n4661 GND.n1467 0.0226631
R10434 GND.n4657 GND.n1467 0.0226631
R10435 GND.n4657 GND.n4656 0.0226631
R10436 GND.n4429 GND.n2375 0.0213333
R10437 GND.n4656 GND.n4655 0.0213333
R10438 GND.n4662 GND.n1466 0.0179419
R10439 GND.n2786 GND.n2785 0.0179419
R10440 GND.n1618 GND.n1572 0.0157439
R10441 GND.n4055 GND.n159 0.0157439
R10442 GND.n4662 GND.n4661 0.014906
R10443 GND.n2787 GND.n2786 0.0118032
R10444 GND.n2786 GND.n2432 0.0113599
R10445 GND.n4663 GND.n4662 0.00825709
R10446 GND.n4429 GND.n4428 0.00182979
R10447 GND.n4655 GND.n4654 0.00182979
R10448 VDD.n2341 VDD.n88 501.952
R10449 VDD.n169 VDD.n86 501.952
R10450 VDD.n2041 VDD.n238 501.952
R10451 VDD.n2143 VDD.n241 501.952
R10452 VDD.n1319 VDD.n607 501.952
R10453 VDD.n1322 VDD.n1321 501.952
R10454 VDD.n827 VDD.n733 501.952
R10455 VDD.n911 VDD.n736 501.952
R10456 VDD.n1835 VDD.n1732 338.05
R10457 VDD.n2007 VDD.n327 338.05
R10458 VDD.n1970 VDD.n1969 338.05
R10459 VDD.n1793 VDD.n1628 338.05
R10460 VDD.n1625 VDD.n466 338.05
R10461 VDD.n1585 VDD.n1584 338.05
R10462 VDD.n1282 VDD.n583 338.05
R10463 VDD.n1427 VDD.n581 338.05
R10464 VDD.n1947 VDD.n1946 338.05
R10465 VDD.n2017 VDD.n319 338.05
R10466 VDD.n1731 VDD.n1629 338.05
R10467 VDD.n1837 VDD.n443 338.05
R10468 VDD.n1570 VDD.n1569 338.05
R10469 VDD.n1526 VDD.n455 338.05
R10470 VDD.n1335 VDD.n584 338.05
R10471 VDD.n1425 VDD.n585 338.05
R10472 VDD.n1336 VDD.t68 252.673
R10473 VDD.n487 VDD.t9 252.673
R10474 VDD.n1228 VDD.t75 252.673
R10475 VDD.n469 VDD.t59 252.673
R10476 VDD.n1631 VDD.t1 252.673
R10477 VDD.n343 VDD.t43 252.673
R10478 VDD.n1743 VDD.t13 252.673
R10479 VDD.n314 VDD.t53 252.673
R10480 VDD.n831 VDD.t20 251.804
R10481 VDD.n851 VDD.t40 251.804
R10482 VDD.n872 VDD.t65 251.804
R10483 VDD.n893 VDD.t47 251.804
R10484 VDD.n598 VDD.t5 251.804
R10485 VDD.n1141 VDD.t31 251.804
R10486 VDD.n1165 VDD.t56 251.804
R10487 VDD.n1189 VDD.t34 251.804
R10488 VDD.n171 VDD.t72 251.804
R10489 VDD.n2271 VDD.t24 251.804
R10490 VDD.n2295 VDD.t37 251.804
R10491 VDD.n2319 VDD.t78 251.804
R10492 VDD.n2069 VDD.t50 251.804
R10493 VDD.n2096 VDD.t16 251.804
R10494 VDD.n2123 VDD.t62 251.804
R10495 VDD.n2045 VDD.t28 251.804
R10496 VDD.n602 VDD.t0 201.612
R10497 VDD.n2141 VDD.t81 201.612
R10498 VDD.n1948 VDD.n1947 185
R10499 VDD.n1947 VDD.n324 185
R10500 VDD.n1949 VDD.n325 185
R10501 VDD.n2012 VDD.n325 185
R10502 VDD.n1951 VDD.n1950 185
R10503 VDD.n1950 VDD.n322 185
R10504 VDD.n1952 VDD.n349 185
R10505 VDD.n1962 VDD.n349 185
R10506 VDD.n1953 VDD.n356 185
R10507 VDD.n356 VDD.n347 185
R10508 VDD.n1955 VDD.n1954 185
R10509 VDD.n1956 VDD.n1955 185
R10510 VDD.n1923 VDD.n355 185
R10511 VDD.n362 VDD.n355 185
R10512 VDD.n1922 VDD.n1921 185
R10513 VDD.n1921 VDD.n1920 185
R10514 VDD.n358 VDD.n357 185
R10515 VDD.n359 VDD.n358 185
R10516 VDD.n1913 VDD.n1912 185
R10517 VDD.n1914 VDD.n1913 185
R10518 VDD.n1911 VDD.n369 185
R10519 VDD.n369 VDD.n366 185
R10520 VDD.n1910 VDD.n1909 185
R10521 VDD.n1909 VDD.n1908 185
R10522 VDD.n371 VDD.n370 185
R10523 VDD.n372 VDD.n371 185
R10524 VDD.n1901 VDD.n1900 185
R10525 VDD.n1902 VDD.n1901 185
R10526 VDD.n1899 VDD.n381 185
R10527 VDD.n381 VDD.n378 185
R10528 VDD.n1898 VDD.n1897 185
R10529 VDD.n1897 VDD.n1896 185
R10530 VDD.n383 VDD.n382 185
R10531 VDD.n384 VDD.n383 185
R10532 VDD.n1889 VDD.n1888 185
R10533 VDD.n1890 VDD.n1889 185
R10534 VDD.n1887 VDD.n392 185
R10535 VDD.n398 VDD.n392 185
R10536 VDD.n1886 VDD.n1885 185
R10537 VDD.n1885 VDD.n1884 185
R10538 VDD.n394 VDD.n393 185
R10539 VDD.n395 VDD.n394 185
R10540 VDD.n1877 VDD.n1876 185
R10541 VDD.n1878 VDD.n1877 185
R10542 VDD.n1875 VDD.n405 185
R10543 VDD.n405 VDD.n402 185
R10544 VDD.n1874 VDD.n1873 185
R10545 VDD.n1873 VDD.n1872 185
R10546 VDD.n407 VDD.n406 185
R10547 VDD.n416 VDD.n407 185
R10548 VDD.n1865 VDD.n1864 185
R10549 VDD.n1866 VDD.n1865 185
R10550 VDD.n1863 VDD.n417 185
R10551 VDD.n417 VDD.n413 185
R10552 VDD.n1862 VDD.n1861 185
R10553 VDD.n1861 VDD.n1860 185
R10554 VDD.n419 VDD.n418 185
R10555 VDD.n420 VDD.n419 185
R10556 VDD.n1853 VDD.n1852 185
R10557 VDD.n1854 VDD.n1853 185
R10558 VDD.n1851 VDD.n428 185
R10559 VDD.n434 VDD.n428 185
R10560 VDD.n1850 VDD.n1849 185
R10561 VDD.n1849 VDD.n1848 185
R10562 VDD.n430 VDD.n429 185
R10563 VDD.n431 VDD.n430 185
R10564 VDD.n1841 VDD.n1840 185
R10565 VDD.n1842 VDD.n1841 185
R10566 VDD.n1839 VDD.n441 185
R10567 VDD.n441 VDD.n438 185
R10568 VDD.n1838 VDD.n1837 185
R10569 VDD.n1837 VDD.n1836 185
R10570 VDD.n443 VDD.n442 185
R10571 VDD.n1644 VDD.n1643 185
R10572 VDD.n1646 VDD.n1645 185
R10573 VDD.n1648 VDD.n1641 185
R10574 VDD.n1651 VDD.n1650 185
R10575 VDD.n1652 VDD.n1640 185
R10576 VDD.n1654 VDD.n1653 185
R10577 VDD.n1656 VDD.n1639 185
R10578 VDD.n1659 VDD.n1658 185
R10579 VDD.n1660 VDD.n1638 185
R10580 VDD.n1662 VDD.n1661 185
R10581 VDD.n1664 VDD.n1637 185
R10582 VDD.n1667 VDD.n1666 185
R10583 VDD.n1668 VDD.n1636 185
R10584 VDD.n1670 VDD.n1669 185
R10585 VDD.n1672 VDD.n1635 185
R10586 VDD.n1675 VDD.n1674 185
R10587 VDD.n1676 VDD.n1634 185
R10588 VDD.n1678 VDD.n1677 185
R10589 VDD.n1681 VDD.n1680 185
R10590 VDD.n1682 VDD.n1629 185
R10591 VDD.n1629 VDD.n1627 185
R10592 VDD.n2017 VDD.n2016 185
R10593 VDD.n2019 VDD.n318 185
R10594 VDD.n2021 VDD.n2020 185
R10595 VDD.n2022 VDD.n313 185
R10596 VDD.n2024 VDD.n2023 185
R10597 VDD.n2026 VDD.n311 185
R10598 VDD.n2028 VDD.n2027 185
R10599 VDD.n2029 VDD.n310 185
R10600 VDD.n2031 VDD.n2030 185
R10601 VDD.n2033 VDD.n307 185
R10602 VDD.n2035 VDD.n2034 185
R10603 VDD.n1931 VDD.n306 185
R10604 VDD.n1933 VDD.n1932 185
R10605 VDD.n1934 VDD.n1929 185
R10606 VDD.n1936 VDD.n1935 185
R10607 VDD.n1938 VDD.n1927 185
R10608 VDD.n1940 VDD.n1939 185
R10609 VDD.n1941 VDD.n1926 185
R10610 VDD.n1943 VDD.n1942 185
R10611 VDD.n1945 VDD.n1925 185
R10612 VDD.n1946 VDD.n1924 185
R10613 VDD.n1946 VDD.n309 185
R10614 VDD.n2015 VDD.n319 185
R10615 VDD.n324 VDD.n319 185
R10616 VDD.n2014 VDD.n2013 185
R10617 VDD.n2013 VDD.n2012 185
R10618 VDD.n321 VDD.n320 185
R10619 VDD.n322 VDD.n321 185
R10620 VDD.n1683 VDD.n348 185
R10621 VDD.n1962 VDD.n348 185
R10622 VDD.n1685 VDD.n1684 185
R10623 VDD.n1684 VDD.n347 185
R10624 VDD.n1686 VDD.n354 185
R10625 VDD.n1956 VDD.n354 185
R10626 VDD.n1688 VDD.n1687 185
R10627 VDD.n1687 VDD.n362 185
R10628 VDD.n1689 VDD.n361 185
R10629 VDD.n1920 VDD.n361 185
R10630 VDD.n1691 VDD.n1690 185
R10631 VDD.n1690 VDD.n359 185
R10632 VDD.n1692 VDD.n368 185
R10633 VDD.n1914 VDD.n368 185
R10634 VDD.n1694 VDD.n1693 185
R10635 VDD.n1693 VDD.n366 185
R10636 VDD.n1695 VDD.n374 185
R10637 VDD.n1908 VDD.n374 185
R10638 VDD.n1697 VDD.n1696 185
R10639 VDD.n1696 VDD.n372 185
R10640 VDD.n1698 VDD.n380 185
R10641 VDD.n1902 VDD.n380 185
R10642 VDD.n1700 VDD.n1699 185
R10643 VDD.n1699 VDD.n378 185
R10644 VDD.n1701 VDD.n386 185
R10645 VDD.n1896 VDD.n386 185
R10646 VDD.n1703 VDD.n1702 185
R10647 VDD.n1702 VDD.n384 185
R10648 VDD.n1704 VDD.n391 185
R10649 VDD.n1890 VDD.n391 185
R10650 VDD.n1706 VDD.n1705 185
R10651 VDD.n1705 VDD.n398 185
R10652 VDD.n1707 VDD.n397 185
R10653 VDD.n1884 VDD.n397 185
R10654 VDD.n1709 VDD.n1708 185
R10655 VDD.n1708 VDD.n395 185
R10656 VDD.n1710 VDD.n404 185
R10657 VDD.n1878 VDD.n404 185
R10658 VDD.n1712 VDD.n1711 185
R10659 VDD.n1711 VDD.n402 185
R10660 VDD.n1713 VDD.n409 185
R10661 VDD.n1872 VDD.n409 185
R10662 VDD.n1715 VDD.n1714 185
R10663 VDD.n1714 VDD.n416 185
R10664 VDD.n1716 VDD.n415 185
R10665 VDD.n1866 VDD.n415 185
R10666 VDD.n1718 VDD.n1717 185
R10667 VDD.n1717 VDD.n413 185
R10668 VDD.n1719 VDD.n422 185
R10669 VDD.n1860 VDD.n422 185
R10670 VDD.n1721 VDD.n1720 185
R10671 VDD.n1720 VDD.n420 185
R10672 VDD.n1722 VDD.n427 185
R10673 VDD.n1854 VDD.n427 185
R10674 VDD.n1724 VDD.n1723 185
R10675 VDD.n1723 VDD.n434 185
R10676 VDD.n1725 VDD.n433 185
R10677 VDD.n1848 VDD.n433 185
R10678 VDD.n1727 VDD.n1726 185
R10679 VDD.n1726 VDD.n431 185
R10680 VDD.n1728 VDD.n440 185
R10681 VDD.n1842 VDD.n440 185
R10682 VDD.n1729 VDD.n1630 185
R10683 VDD.n1630 VDD.n438 185
R10684 VDD.n1731 VDD.n1730 185
R10685 VDD.n1836 VDD.n1731 185
R10686 VDD.n1319 VDD.n1318 185
R10687 VDD.n1320 VDD.n1319 185
R10688 VDD.n608 VDD.n606 185
R10689 VDD.n606 VDD.n605 185
R10690 VDD.n1060 VDD.n1059 185
R10691 VDD.n1059 VDD.n1058 185
R10692 VDD.n611 VDD.n610 185
R10693 VDD.n619 VDD.n611 185
R10694 VDD.n1046 VDD.n1045 185
R10695 VDD.n1047 VDD.n1046 185
R10696 VDD.n621 VDD.n620 185
R10697 VDD.n620 VDD.n618 185
R10698 VDD.n1041 VDD.n1040 185
R10699 VDD.n1040 VDD.n1039 185
R10700 VDD.n624 VDD.n623 185
R10701 VDD.n625 VDD.n624 185
R10702 VDD.n1030 VDD.n1029 185
R10703 VDD.n1031 VDD.n1030 185
R10704 VDD.n633 VDD.n632 185
R10705 VDD.n632 VDD.n631 185
R10706 VDD.n1025 VDD.n1024 185
R10707 VDD.n1024 VDD.n1023 185
R10708 VDD.n636 VDD.n635 185
R10709 VDD.n637 VDD.n636 185
R10710 VDD.n1014 VDD.n1013 185
R10711 VDD.n1015 VDD.n1014 185
R10712 VDD.n645 VDD.n644 185
R10713 VDD.n644 VDD.n643 185
R10714 VDD.n1009 VDD.n1008 185
R10715 VDD.n1008 VDD.n1007 185
R10716 VDD.n648 VDD.n647 185
R10717 VDD.n649 VDD.n648 185
R10718 VDD.n998 VDD.n997 185
R10719 VDD.n999 VDD.n998 185
R10720 VDD.n657 VDD.n656 185
R10721 VDD.n656 VDD.n655 185
R10722 VDD.n993 VDD.n992 185
R10723 VDD.n992 VDD.n991 185
R10724 VDD.n680 VDD.n679 185
R10725 VDD.n687 VDD.n680 185
R10726 VDD.n982 VDD.n981 185
R10727 VDD.n983 VDD.n982 185
R10728 VDD.n689 VDD.n688 185
R10729 VDD.n688 VDD.n686 185
R10730 VDD.n976 VDD.n975 185
R10731 VDD.n975 VDD.n974 185
R10732 VDD.n692 VDD.n691 185
R10733 VDD.n693 VDD.n692 185
R10734 VDD.n965 VDD.n964 185
R10735 VDD.n966 VDD.n965 185
R10736 VDD.n701 VDD.n700 185
R10737 VDD.n700 VDD.n699 185
R10738 VDD.n960 VDD.n959 185
R10739 VDD.n959 VDD.n958 185
R10740 VDD.n704 VDD.n703 185
R10741 VDD.n705 VDD.n704 185
R10742 VDD.n949 VDD.n948 185
R10743 VDD.n950 VDD.n949 185
R10744 VDD.n713 VDD.n712 185
R10745 VDD.n712 VDD.n711 185
R10746 VDD.n944 VDD.n943 185
R10747 VDD.n943 VDD.n942 185
R10748 VDD.n716 VDD.n715 185
R10749 VDD.n717 VDD.n716 185
R10750 VDD.n933 VDD.n932 185
R10751 VDD.n934 VDD.n933 185
R10752 VDD.n725 VDD.n724 185
R10753 VDD.n724 VDD.n723 185
R10754 VDD.n928 VDD.n927 185
R10755 VDD.n927 VDD.n926 185
R10756 VDD.n728 VDD.n727 185
R10757 VDD.n735 VDD.n728 185
R10758 VDD.n917 VDD.n916 185
R10759 VDD.n918 VDD.n917 185
R10760 VDD.n737 VDD.n736 185
R10761 VDD.n736 VDD.n734 185
R10762 VDD.n912 VDD.n911 185
R10763 VDD.n740 VDD.n739 185
R10764 VDD.n908 VDD.n907 185
R10765 VDD.n909 VDD.n908 185
R10766 VDD.n764 VDD.n763 185
R10767 VDD.n903 VDD.n766 185
R10768 VDD.n902 VDD.n767 185
R10769 VDD.n901 VDD.n768 185
R10770 VDD.n770 VDD.n769 185
R10771 VDD.n897 VDD.n772 185
R10772 VDD.n896 VDD.n773 185
R10773 VDD.n892 VDD.n774 185
R10774 VDD.n776 VDD.n775 185
R10775 VDD.n888 VDD.n778 185
R10776 VDD.n887 VDD.n779 185
R10777 VDD.n886 VDD.n780 185
R10778 VDD.n782 VDD.n781 185
R10779 VDD.n882 VDD.n784 185
R10780 VDD.n881 VDD.n785 185
R10781 VDD.n880 VDD.n786 185
R10782 VDD.n788 VDD.n787 185
R10783 VDD.n876 VDD.n790 185
R10784 VDD.n875 VDD.n791 185
R10785 VDD.n871 VDD.n792 185
R10786 VDD.n794 VDD.n793 185
R10787 VDD.n867 VDD.n796 185
R10788 VDD.n866 VDD.n797 185
R10789 VDD.n865 VDD.n798 185
R10790 VDD.n800 VDD.n799 185
R10791 VDD.n861 VDD.n802 185
R10792 VDD.n860 VDD.n803 185
R10793 VDD.n859 VDD.n804 185
R10794 VDD.n806 VDD.n805 185
R10795 VDD.n855 VDD.n808 185
R10796 VDD.n854 VDD.n809 185
R10797 VDD.n850 VDD.n810 185
R10798 VDD.n812 VDD.n811 185
R10799 VDD.n846 VDD.n814 185
R10800 VDD.n845 VDD.n815 185
R10801 VDD.n844 VDD.n816 185
R10802 VDD.n818 VDD.n817 185
R10803 VDD.n840 VDD.n820 185
R10804 VDD.n839 VDD.n821 185
R10805 VDD.n838 VDD.n822 185
R10806 VDD.n824 VDD.n823 185
R10807 VDD.n834 VDD.n826 185
R10808 VDD.n833 VDD.n830 185
R10809 VDD.n829 VDD.n827 185
R10810 VDD.n1322 VDD.n597 185
R10811 VDD.n1325 VDD.n1324 185
R10812 VDD.n1326 VDD.n596 185
R10813 VDD.n1327 VDD.n595 185
R10814 VDD.n1124 VDD.n594 185
R10815 VDD.n1127 VDD.n1126 185
R10816 VDD.n1129 VDD.n1128 185
R10817 VDD.n1131 VDD.n1122 185
R10818 VDD.n1133 VDD.n1132 185
R10819 VDD.n1134 VDD.n1118 185
R10820 VDD.n1136 VDD.n1135 185
R10821 VDD.n1138 VDD.n1116 185
R10822 VDD.n1140 VDD.n1139 185
R10823 VDD.n1144 VDD.n1111 185
R10824 VDD.n1146 VDD.n1145 185
R10825 VDD.n1148 VDD.n1109 185
R10826 VDD.n1150 VDD.n1149 185
R10827 VDD.n1151 VDD.n1104 185
R10828 VDD.n1153 VDD.n1152 185
R10829 VDD.n1155 VDD.n1102 185
R10830 VDD.n1157 VDD.n1156 185
R10831 VDD.n1158 VDD.n1097 185
R10832 VDD.n1160 VDD.n1159 185
R10833 VDD.n1162 VDD.n1095 185
R10834 VDD.n1164 VDD.n1163 185
R10835 VDD.n1168 VDD.n1090 185
R10836 VDD.n1170 VDD.n1169 185
R10837 VDD.n1172 VDD.n1088 185
R10838 VDD.n1174 VDD.n1173 185
R10839 VDD.n1175 VDD.n1083 185
R10840 VDD.n1177 VDD.n1176 185
R10841 VDD.n1179 VDD.n1081 185
R10842 VDD.n1181 VDD.n1180 185
R10843 VDD.n1182 VDD.n1076 185
R10844 VDD.n1184 VDD.n1183 185
R10845 VDD.n1186 VDD.n1074 185
R10846 VDD.n1188 VDD.n1187 185
R10847 VDD.n1192 VDD.n1071 185
R10848 VDD.n1194 VDD.n1193 185
R10849 VDD.n1196 VDD.n1069 185
R10850 VDD.n1198 VDD.n1197 185
R10851 VDD.n1067 VDD.n1066 185
R10852 VDD.n1308 VDD.n1307 185
R10853 VDD.n1310 VDD.n1065 185
R10854 VDD.n1311 VDD.n1064 185
R10855 VDD.n1314 VDD.n1313 185
R10856 VDD.n1315 VDD.n607 185
R10857 VDD.n607 VDD.n602 185
R10858 VDD.n1321 VDD.n604 185
R10859 VDD.n1321 VDD.n1320 185
R10860 VDD.n614 VDD.n603 185
R10861 VDD.n605 VDD.n603 185
R10862 VDD.n1057 VDD.n1056 185
R10863 VDD.n1058 VDD.n1057 185
R10864 VDD.n613 VDD.n612 185
R10865 VDD.n619 VDD.n612 185
R10866 VDD.n1049 VDD.n1048 185
R10867 VDD.n1048 VDD.n1047 185
R10868 VDD.n617 VDD.n616 185
R10869 VDD.n618 VDD.n617 185
R10870 VDD.n1038 VDD.n1037 185
R10871 VDD.n1039 VDD.n1038 185
R10872 VDD.n627 VDD.n626 185
R10873 VDD.n626 VDD.n625 185
R10874 VDD.n1033 VDD.n1032 185
R10875 VDD.n1032 VDD.n1031 185
R10876 VDD.n630 VDD.n629 185
R10877 VDD.n631 VDD.n630 185
R10878 VDD.n1022 VDD.n1021 185
R10879 VDD.n1023 VDD.n1022 185
R10880 VDD.n639 VDD.n638 185
R10881 VDD.n638 VDD.n637 185
R10882 VDD.n1017 VDD.n1016 185
R10883 VDD.n1016 VDD.n1015 185
R10884 VDD.n642 VDD.n641 185
R10885 VDD.n643 VDD.n642 185
R10886 VDD.n1006 VDD.n1005 185
R10887 VDD.n1007 VDD.n1006 185
R10888 VDD.n651 VDD.n650 185
R10889 VDD.n650 VDD.n649 185
R10890 VDD.n1001 VDD.n1000 185
R10891 VDD.n1000 VDD.n999 185
R10892 VDD.n654 VDD.n653 185
R10893 VDD.n655 VDD.n654 185
R10894 VDD.n990 VDD.n989 185
R10895 VDD.n991 VDD.n990 185
R10896 VDD.n682 VDD.n681 185
R10897 VDD.n687 VDD.n681 185
R10898 VDD.n985 VDD.n984 185
R10899 VDD.n984 VDD.n983 185
R10900 VDD.n685 VDD.n684 185
R10901 VDD.n686 VDD.n685 185
R10902 VDD.n973 VDD.n972 185
R10903 VDD.n974 VDD.n973 185
R10904 VDD.n695 VDD.n694 185
R10905 VDD.n694 VDD.n693 185
R10906 VDD.n968 VDD.n967 185
R10907 VDD.n967 VDD.n966 185
R10908 VDD.n698 VDD.n697 185
R10909 VDD.n699 VDD.n698 185
R10910 VDD.n957 VDD.n956 185
R10911 VDD.n958 VDD.n957 185
R10912 VDD.n707 VDD.n706 185
R10913 VDD.n706 VDD.n705 185
R10914 VDD.n952 VDD.n951 185
R10915 VDD.n951 VDD.n950 185
R10916 VDD.n710 VDD.n709 185
R10917 VDD.n711 VDD.n710 185
R10918 VDD.n941 VDD.n940 185
R10919 VDD.n942 VDD.n941 185
R10920 VDD.n719 VDD.n718 185
R10921 VDD.n718 VDD.n717 185
R10922 VDD.n936 VDD.n935 185
R10923 VDD.n935 VDD.n934 185
R10924 VDD.n722 VDD.n721 185
R10925 VDD.n723 VDD.n722 185
R10926 VDD.n925 VDD.n924 185
R10927 VDD.n926 VDD.n925 185
R10928 VDD.n730 VDD.n729 185
R10929 VDD.n735 VDD.n729 185
R10930 VDD.n920 VDD.n919 185
R10931 VDD.n919 VDD.n918 185
R10932 VDD.n733 VDD.n732 185
R10933 VDD.n734 VDD.n733 185
R10934 VDD.n468 VDD.n466 185
R10935 VDD.n466 VDD.n444 185
R10936 VDD.n1581 VDD.n1580 185
R10937 VDD.n1582 VDD.n1581 185
R10938 VDD.n1579 VDD.n478 185
R10939 VDD.n478 VDD.n475 185
R10940 VDD.n1578 VDD.n1577 185
R10941 VDD.n1577 VDD.n1576 185
R10942 VDD.n480 VDD.n479 185
R10943 VDD.n481 VDD.n480 185
R10944 VDD.n1517 VDD.n1516 185
R10945 VDD.n1518 VDD.n1517 185
R10946 VDD.n1515 VDD.n493 185
R10947 VDD.n499 VDD.n493 185
R10948 VDD.n1514 VDD.n1513 185
R10949 VDD.n1513 VDD.n1512 185
R10950 VDD.n495 VDD.n494 185
R10951 VDD.n496 VDD.n495 185
R10952 VDD.n1503 VDD.n1502 185
R10953 VDD.n1504 VDD.n1503 185
R10954 VDD.n1501 VDD.n507 185
R10955 VDD.n507 VDD.n504 185
R10956 VDD.n1500 VDD.n1499 185
R10957 VDD.n1499 VDD.n1498 185
R10958 VDD.n509 VDD.n508 185
R10959 VDD.n518 VDD.n509 185
R10960 VDD.n1491 VDD.n1490 185
R10961 VDD.n1492 VDD.n1491 185
R10962 VDD.n1489 VDD.n519 185
R10963 VDD.n519 VDD.n515 185
R10964 VDD.n1488 VDD.n1487 185
R10965 VDD.n1487 VDD.n1486 185
R10966 VDD.n521 VDD.n520 185
R10967 VDD.n522 VDD.n521 185
R10968 VDD.n1479 VDD.n1478 185
R10969 VDD.n1480 VDD.n1479 185
R10970 VDD.n1477 VDD.n530 185
R10971 VDD.n536 VDD.n530 185
R10972 VDD.n1476 VDD.n1475 185
R10973 VDD.n1475 VDD.n1474 185
R10974 VDD.n532 VDD.n531 185
R10975 VDD.n533 VDD.n532 185
R10976 VDD.n1467 VDD.n1466 185
R10977 VDD.n1468 VDD.n1467 185
R10978 VDD.n1465 VDD.n543 185
R10979 VDD.n543 VDD.n540 185
R10980 VDD.n1464 VDD.n1463 185
R10981 VDD.n1463 VDD.n1462 185
R10982 VDD.n545 VDD.n544 185
R10983 VDD.n546 VDD.n545 185
R10984 VDD.n1455 VDD.n1454 185
R10985 VDD.n1456 VDD.n1455 185
R10986 VDD.n1453 VDD.n555 185
R10987 VDD.n555 VDD.n552 185
R10988 VDD.n1452 VDD.n1451 185
R10989 VDD.n1451 VDD.n1450 185
R10990 VDD.n557 VDD.n556 185
R10991 VDD.n558 VDD.n557 185
R10992 VDD.n1443 VDD.n1442 185
R10993 VDD.n1444 VDD.n1443 185
R10994 VDD.n1441 VDD.n566 185
R10995 VDD.n572 VDD.n566 185
R10996 VDD.n1440 VDD.n1439 185
R10997 VDD.n1439 VDD.n1438 185
R10998 VDD.n568 VDD.n567 185
R10999 VDD.n569 VDD.n568 185
R11000 VDD.n1431 VDD.n1430 185
R11001 VDD.n1432 VDD.n1431 185
R11002 VDD.n1429 VDD.n579 185
R11003 VDD.n579 VDD.n576 185
R11004 VDD.n1428 VDD.n1427 185
R11005 VDD.n1427 VDD.n1426 185
R11006 VDD.n581 VDD.n580 185
R11007 VDD.n1207 VDD.n1206 185
R11008 VDD.n1208 VDD.n1204 185
R11009 VDD.n1204 VDD.n582 185
R11010 VDD.n1210 VDD.n1209 185
R11011 VDD.n1212 VDD.n1203 185
R11012 VDD.n1215 VDD.n1214 185
R11013 VDD.n1216 VDD.n1202 185
R11014 VDD.n1218 VDD.n1217 185
R11015 VDD.n1220 VDD.n1201 185
R11016 VDD.n1221 VDD.n1200 185
R11017 VDD.n1302 VDD.n1223 185
R11018 VDD.n1301 VDD.n1300 185
R11019 VDD.n1298 VDD.n1224 185
R11020 VDD.n1297 VDD.n1296 185
R11021 VDD.n1295 VDD.n1294 185
R11022 VDD.n1293 VDD.n1226 185
R11023 VDD.n1291 VDD.n1290 185
R11024 VDD.n1289 VDD.n1227 185
R11025 VDD.n1288 VDD.n1287 185
R11026 VDD.n1285 VDD.n1284 185
R11027 VDD.n1283 VDD.n1282 185
R11028 VDD.n1586 VDD.n1585 185
R11029 VDD.n1588 VDD.n1587 185
R11030 VDD.n1590 VDD.n1589 185
R11031 VDD.n1592 VDD.n1591 185
R11032 VDD.n1594 VDD.n1593 185
R11033 VDD.n1596 VDD.n1595 185
R11034 VDD.n1598 VDD.n1597 185
R11035 VDD.n1600 VDD.n1599 185
R11036 VDD.n1602 VDD.n1601 185
R11037 VDD.n1604 VDD.n1603 185
R11038 VDD.n1606 VDD.n1605 185
R11039 VDD.n1608 VDD.n1607 185
R11040 VDD.n1610 VDD.n1609 185
R11041 VDD.n1612 VDD.n1611 185
R11042 VDD.n1614 VDD.n1613 185
R11043 VDD.n1616 VDD.n1615 185
R11044 VDD.n1618 VDD.n1617 185
R11045 VDD.n1620 VDD.n1619 185
R11046 VDD.n1622 VDD.n1621 185
R11047 VDD.n1623 VDD.n467 185
R11048 VDD.n1625 VDD.n1624 185
R11049 VDD.n1626 VDD.n1625 185
R11050 VDD.n1584 VDD.n472 185
R11051 VDD.n1584 VDD.n444 185
R11052 VDD.n1583 VDD.n474 185
R11053 VDD.n1583 VDD.n1582 185
R11054 VDD.n1232 VDD.n473 185
R11055 VDD.n475 VDD.n473 185
R11056 VDD.n1233 VDD.n482 185
R11057 VDD.n1576 VDD.n482 185
R11058 VDD.n1235 VDD.n1234 185
R11059 VDD.n1234 VDD.n481 185
R11060 VDD.n1236 VDD.n491 185
R11061 VDD.n1518 VDD.n491 185
R11062 VDD.n1238 VDD.n1237 185
R11063 VDD.n1237 VDD.n499 185
R11064 VDD.n1239 VDD.n497 185
R11065 VDD.n1512 VDD.n497 185
R11066 VDD.n1241 VDD.n1240 185
R11067 VDD.n1240 VDD.n496 185
R11068 VDD.n1242 VDD.n505 185
R11069 VDD.n1504 VDD.n505 185
R11070 VDD.n1244 VDD.n1243 185
R11071 VDD.n1243 VDD.n504 185
R11072 VDD.n1245 VDD.n510 185
R11073 VDD.n1498 VDD.n510 185
R11074 VDD.n1247 VDD.n1246 185
R11075 VDD.n1246 VDD.n518 185
R11076 VDD.n1248 VDD.n516 185
R11077 VDD.n1492 VDD.n516 185
R11078 VDD.n1250 VDD.n1249 185
R11079 VDD.n1249 VDD.n515 185
R11080 VDD.n1251 VDD.n523 185
R11081 VDD.n1486 VDD.n523 185
R11082 VDD.n1253 VDD.n1252 185
R11083 VDD.n1252 VDD.n522 185
R11084 VDD.n1254 VDD.n528 185
R11085 VDD.n1480 VDD.n528 185
R11086 VDD.n1256 VDD.n1255 185
R11087 VDD.n1255 VDD.n536 185
R11088 VDD.n1257 VDD.n534 185
R11089 VDD.n1474 VDD.n534 185
R11090 VDD.n1259 VDD.n1258 185
R11091 VDD.n1258 VDD.n533 185
R11092 VDD.n1260 VDD.n541 185
R11093 VDD.n1468 VDD.n541 185
R11094 VDD.n1262 VDD.n1261 185
R11095 VDD.n1261 VDD.n540 185
R11096 VDD.n1263 VDD.n547 185
R11097 VDD.n1462 VDD.n547 185
R11098 VDD.n1265 VDD.n1264 185
R11099 VDD.n1264 VDD.n546 185
R11100 VDD.n1266 VDD.n553 185
R11101 VDD.n1456 VDD.n553 185
R11102 VDD.n1268 VDD.n1267 185
R11103 VDD.n1267 VDD.n552 185
R11104 VDD.n1269 VDD.n559 185
R11105 VDD.n1450 VDD.n559 185
R11106 VDD.n1271 VDD.n1270 185
R11107 VDD.n1270 VDD.n558 185
R11108 VDD.n1272 VDD.n564 185
R11109 VDD.n1444 VDD.n564 185
R11110 VDD.n1274 VDD.n1273 185
R11111 VDD.n1273 VDD.n572 185
R11112 VDD.n1275 VDD.n570 185
R11113 VDD.n1438 VDD.n570 185
R11114 VDD.n1277 VDD.n1276 185
R11115 VDD.n1276 VDD.n569 185
R11116 VDD.n1278 VDD.n577 185
R11117 VDD.n1432 VDD.n577 185
R11118 VDD.n1280 VDD.n1279 185
R11119 VDD.n1279 VDD.n576 185
R11120 VDD.n1281 VDD.n583 185
R11121 VDD.n1426 VDD.n583 185
R11122 VDD.n2341 VDD.n2340 185
R11123 VDD.n2342 VDD.n2341 185
R11124 VDD.n83 VDD.n82 185
R11125 VDD.n2343 VDD.n83 185
R11126 VDD.n2346 VDD.n2345 185
R11127 VDD.n2345 VDD.n2344 185
R11128 VDD.n2347 VDD.n77 185
R11129 VDD.n77 VDD.n76 185
R11130 VDD.n2349 VDD.n2348 185
R11131 VDD.n2350 VDD.n2349 185
R11132 VDD.n72 VDD.n71 185
R11133 VDD.n2351 VDD.n72 185
R11134 VDD.n2354 VDD.n2353 185
R11135 VDD.n2353 VDD.n2352 185
R11136 VDD.n2355 VDD.n66 185
R11137 VDD.n66 VDD.n65 185
R11138 VDD.n2357 VDD.n2356 185
R11139 VDD.n2358 VDD.n2357 185
R11140 VDD.n61 VDD.n60 185
R11141 VDD.n2359 VDD.n61 185
R11142 VDD.n2362 VDD.n2361 185
R11143 VDD.n2361 VDD.n2360 185
R11144 VDD.n2363 VDD.n55 185
R11145 VDD.n55 VDD.n54 185
R11146 VDD.n2365 VDD.n2364 185
R11147 VDD.n2366 VDD.n2365 185
R11148 VDD.n50 VDD.n49 185
R11149 VDD.n2367 VDD.n50 185
R11150 VDD.n2370 VDD.n2369 185
R11151 VDD.n2369 VDD.n2368 185
R11152 VDD.n2371 VDD.n45 185
R11153 VDD.n45 VDD.n44 185
R11154 VDD.n2373 VDD.n2372 185
R11155 VDD.n2374 VDD.n2373 185
R11156 VDD.n40 VDD.n38 185
R11157 VDD.n2375 VDD.n40 185
R11158 VDD.n2378 VDD.n2377 185
R11159 VDD.n2377 VDD.n2376 185
R11160 VDD.n39 VDD.n37 185
R11161 VDD.n192 VDD.n39 185
R11162 VDD.n2213 VDD.n2212 185
R11163 VDD.n2214 VDD.n2213 185
R11164 VDD.n194 VDD.n193 185
R11165 VDD.n193 VDD.n191 185
R11166 VDD.n2208 VDD.n2207 185
R11167 VDD.n2207 VDD.n2206 185
R11168 VDD.n197 VDD.n196 185
R11169 VDD.n198 VDD.n197 185
R11170 VDD.n2197 VDD.n2196 185
R11171 VDD.n2198 VDD.n2197 185
R11172 VDD.n206 VDD.n205 185
R11173 VDD.n205 VDD.n204 185
R11174 VDD.n2192 VDD.n2191 185
R11175 VDD.n2191 VDD.n2190 185
R11176 VDD.n209 VDD.n208 185
R11177 VDD.n210 VDD.n209 185
R11178 VDD.n2181 VDD.n2180 185
R11179 VDD.n2182 VDD.n2181 185
R11180 VDD.n218 VDD.n217 185
R11181 VDD.n217 VDD.n216 185
R11182 VDD.n2176 VDD.n2175 185
R11183 VDD.n2175 VDD.n2174 185
R11184 VDD.n221 VDD.n220 185
R11185 VDD.n222 VDD.n221 185
R11186 VDD.n2165 VDD.n2164 185
R11187 VDD.n2166 VDD.n2165 185
R11188 VDD.n230 VDD.n229 185
R11189 VDD.n229 VDD.n228 185
R11190 VDD.n2160 VDD.n2159 185
R11191 VDD.n2159 VDD.n2158 185
R11192 VDD.n233 VDD.n232 185
R11193 VDD.n240 VDD.n233 185
R11194 VDD.n2149 VDD.n2148 185
R11195 VDD.n2150 VDD.n2149 185
R11196 VDD.n242 VDD.n241 185
R11197 VDD.n241 VDD.n239 185
R11198 VDD.n2144 VDD.n2143 185
R11199 VDD.n245 VDD.n244 185
R11200 VDD.n2140 VDD.n2139 185
R11201 VDD.n2141 VDD.n2140 185
R11202 VDD.n2138 VDD.n268 185
R11203 VDD.n2137 VDD.n2136 185
R11204 VDD.n2135 VDD.n2134 185
R11205 VDD.n2133 VDD.n2132 185
R11206 VDD.n2131 VDD.n2130 185
R11207 VDD.n2129 VDD.n2128 185
R11208 VDD.n2127 VDD.n2126 185
R11209 VDD.n2122 VDD.n2121 185
R11210 VDD.n2120 VDD.n2119 185
R11211 VDD.n2118 VDD.n2117 185
R11212 VDD.n2116 VDD.n2115 185
R11213 VDD.n2114 VDD.n2113 185
R11214 VDD.n2112 VDD.n2111 185
R11215 VDD.n2110 VDD.n2109 185
R11216 VDD.n2108 VDD.n2107 185
R11217 VDD.n2106 VDD.n2105 185
R11218 VDD.n2104 VDD.n2103 185
R11219 VDD.n2102 VDD.n2101 185
R11220 VDD.n2100 VDD.n2099 185
R11221 VDD.n2095 VDD.n2094 185
R11222 VDD.n2093 VDD.n2092 185
R11223 VDD.n2091 VDD.n2090 185
R11224 VDD.n2089 VDD.n2088 185
R11225 VDD.n2087 VDD.n2086 185
R11226 VDD.n2085 VDD.n2084 185
R11227 VDD.n2083 VDD.n2082 185
R11228 VDD.n2081 VDD.n2080 185
R11229 VDD.n2079 VDD.n2078 185
R11230 VDD.n2077 VDD.n2076 185
R11231 VDD.n2075 VDD.n2074 185
R11232 VDD.n2073 VDD.n2072 185
R11233 VDD.n2068 VDD.n2067 185
R11234 VDD.n2066 VDD.n2065 185
R11235 VDD.n2064 VDD.n2063 185
R11236 VDD.n2062 VDD.n2061 185
R11237 VDD.n2060 VDD.n2059 185
R11238 VDD.n2058 VDD.n2057 185
R11239 VDD.n2036 VDD.n304 185
R11240 VDD.n2038 VDD.n2037 185
R11241 VDD.n2053 VDD.n2039 185
R11242 VDD.n2052 VDD.n2051 185
R11243 VDD.n2050 VDD.n2049 185
R11244 VDD.n2048 VDD.n2047 185
R11245 VDD.n2042 VDD.n2041 185
R11246 VDD.n170 VDD.n169 185
R11247 VDD.n2250 VDD.n165 185
R11248 VDD.n2252 VDD.n2251 185
R11249 VDD.n2254 VDD.n163 185
R11250 VDD.n2256 VDD.n2255 185
R11251 VDD.n2257 VDD.n158 185
R11252 VDD.n2259 VDD.n2258 185
R11253 VDD.n2261 VDD.n156 185
R11254 VDD.n2263 VDD.n2262 185
R11255 VDD.n2264 VDD.n151 185
R11256 VDD.n2266 VDD.n2265 185
R11257 VDD.n2268 VDD.n149 185
R11258 VDD.n2270 VDD.n2269 185
R11259 VDD.n2274 VDD.n144 185
R11260 VDD.n2276 VDD.n2275 185
R11261 VDD.n2278 VDD.n142 185
R11262 VDD.n2280 VDD.n2279 185
R11263 VDD.n2281 VDD.n137 185
R11264 VDD.n2283 VDD.n2282 185
R11265 VDD.n2285 VDD.n135 185
R11266 VDD.n2287 VDD.n2286 185
R11267 VDD.n2288 VDD.n130 185
R11268 VDD.n2290 VDD.n2289 185
R11269 VDD.n2292 VDD.n128 185
R11270 VDD.n2294 VDD.n2293 185
R11271 VDD.n2298 VDD.n123 185
R11272 VDD.n2300 VDD.n2299 185
R11273 VDD.n2302 VDD.n121 185
R11274 VDD.n2304 VDD.n2303 185
R11275 VDD.n2305 VDD.n116 185
R11276 VDD.n2307 VDD.n2306 185
R11277 VDD.n2309 VDD.n114 185
R11278 VDD.n2311 VDD.n2310 185
R11279 VDD.n2312 VDD.n109 185
R11280 VDD.n2314 VDD.n2313 185
R11281 VDD.n2316 VDD.n107 185
R11282 VDD.n2318 VDD.n2317 185
R11283 VDD.n2322 VDD.n102 185
R11284 VDD.n2324 VDD.n2323 185
R11285 VDD.n2326 VDD.n100 185
R11286 VDD.n2328 VDD.n2327 185
R11287 VDD.n2329 VDD.n95 185
R11288 VDD.n2331 VDD.n2330 185
R11289 VDD.n2333 VDD.n93 185
R11290 VDD.n2335 VDD.n2334 185
R11291 VDD.n2336 VDD.n91 185
R11292 VDD.n2337 VDD.n88 185
R11293 VDD.n88 VDD.n87 185
R11294 VDD.n2246 VDD.n86 185
R11295 VDD.n2342 VDD.n86 185
R11296 VDD.n2245 VDD.n85 185
R11297 VDD.n2343 VDD.n85 185
R11298 VDD.n2244 VDD.n84 185
R11299 VDD.n2344 VDD.n84 185
R11300 VDD.n175 VDD.n174 185
R11301 VDD.n174 VDD.n76 185
R11302 VDD.n2240 VDD.n75 185
R11303 VDD.n2350 VDD.n75 185
R11304 VDD.n2239 VDD.n74 185
R11305 VDD.n2351 VDD.n74 185
R11306 VDD.n2238 VDD.n73 185
R11307 VDD.n2352 VDD.n73 185
R11308 VDD.n178 VDD.n177 185
R11309 VDD.n177 VDD.n65 185
R11310 VDD.n2234 VDD.n64 185
R11311 VDD.n2358 VDD.n64 185
R11312 VDD.n2233 VDD.n63 185
R11313 VDD.n2359 VDD.n63 185
R11314 VDD.n2232 VDD.n62 185
R11315 VDD.n2360 VDD.n62 185
R11316 VDD.n181 VDD.n180 185
R11317 VDD.n180 VDD.n54 185
R11318 VDD.n2228 VDD.n53 185
R11319 VDD.n2366 VDD.n53 185
R11320 VDD.n2227 VDD.n52 185
R11321 VDD.n2367 VDD.n52 185
R11322 VDD.n2226 VDD.n51 185
R11323 VDD.n2368 VDD.n51 185
R11324 VDD.n184 VDD.n183 185
R11325 VDD.n183 VDD.n44 185
R11326 VDD.n2222 VDD.n43 185
R11327 VDD.n2374 VDD.n43 185
R11328 VDD.n2221 VDD.n42 185
R11329 VDD.n2375 VDD.n42 185
R11330 VDD.n2220 VDD.n41 185
R11331 VDD.n2376 VDD.n41 185
R11332 VDD.n190 VDD.n186 185
R11333 VDD.n192 VDD.n190 185
R11334 VDD.n2216 VDD.n2215 185
R11335 VDD.n2215 VDD.n2214 185
R11336 VDD.n189 VDD.n188 185
R11337 VDD.n191 VDD.n189 185
R11338 VDD.n2205 VDD.n2204 185
R11339 VDD.n2206 VDD.n2205 185
R11340 VDD.n200 VDD.n199 185
R11341 VDD.n199 VDD.n198 185
R11342 VDD.n2200 VDD.n2199 185
R11343 VDD.n2199 VDD.n2198 185
R11344 VDD.n203 VDD.n202 185
R11345 VDD.n204 VDD.n203 185
R11346 VDD.n2189 VDD.n2188 185
R11347 VDD.n2190 VDD.n2189 185
R11348 VDD.n212 VDD.n211 185
R11349 VDD.n211 VDD.n210 185
R11350 VDD.n2184 VDD.n2183 185
R11351 VDD.n2183 VDD.n2182 185
R11352 VDD.n215 VDD.n214 185
R11353 VDD.n216 VDD.n215 185
R11354 VDD.n2173 VDD.n2172 185
R11355 VDD.n2174 VDD.n2173 185
R11356 VDD.n224 VDD.n223 185
R11357 VDD.n223 VDD.n222 185
R11358 VDD.n2168 VDD.n2167 185
R11359 VDD.n2167 VDD.n2166 185
R11360 VDD.n227 VDD.n226 185
R11361 VDD.n228 VDD.n227 185
R11362 VDD.n2157 VDD.n2156 185
R11363 VDD.n2158 VDD.n2157 185
R11364 VDD.n235 VDD.n234 185
R11365 VDD.n240 VDD.n234 185
R11366 VDD.n2152 VDD.n2151 185
R11367 VDD.n2151 VDD.n2150 185
R11368 VDD.n238 VDD.n237 185
R11369 VDD.n239 VDD.n238 185
R11370 VDD.n1833 VDD.n1732 185
R11371 VDD.n1832 VDD.n1831 185
R11372 VDD.n1829 VDD.n1733 185
R11373 VDD.n1829 VDD.n1627 185
R11374 VDD.n1828 VDD.n1827 185
R11375 VDD.n1826 VDD.n1825 185
R11376 VDD.n1824 VDD.n1735 185
R11377 VDD.n1822 VDD.n1821 185
R11378 VDD.n1820 VDD.n1736 185
R11379 VDD.n1819 VDD.n1818 185
R11380 VDD.n1816 VDD.n1737 185
R11381 VDD.n1814 VDD.n1813 185
R11382 VDD.n1812 VDD.n1738 185
R11383 VDD.n1811 VDD.n1810 185
R11384 VDD.n1808 VDD.n1739 185
R11385 VDD.n1806 VDD.n1805 185
R11386 VDD.n1804 VDD.n1740 185
R11387 VDD.n1803 VDD.n1802 185
R11388 VDD.n1800 VDD.n1741 185
R11389 VDD.n1798 VDD.n1797 185
R11390 VDD.n1795 VDD.n1742 185
R11391 VDD.n1794 VDD.n1793 185
R11392 VDD.n1971 VDD.n1970 185
R11393 VDD.n1972 VDD.n342 185
R11394 VDD.n1975 VDD.n1974 185
R11395 VDD.n1977 VDD.n340 185
R11396 VDD.n1979 VDD.n1978 185
R11397 VDD.n1980 VDD.n339 185
R11398 VDD.n1982 VDD.n1981 185
R11399 VDD.n1984 VDD.n337 185
R11400 VDD.n1986 VDD.n1985 185
R11401 VDD.n1987 VDD.n336 185
R11402 VDD.n1990 VDD.n1989 185
R11403 VDD.n1992 VDD.n334 185
R11404 VDD.n1994 VDD.n1993 185
R11405 VDD.n1995 VDD.n333 185
R11406 VDD.n1997 VDD.n1996 185
R11407 VDD.n1999 VDD.n331 185
R11408 VDD.n2001 VDD.n2000 185
R11409 VDD.n2002 VDD.n330 185
R11410 VDD.n2004 VDD.n2003 185
R11411 VDD.n2006 VDD.n329 185
R11412 VDD.n2008 VDD.n2007 185
R11413 VDD.n2007 VDD.n309 185
R11414 VDD.n1969 VDD.n1967 185
R11415 VDD.n1969 VDD.n324 185
R11416 VDD.n1966 VDD.n323 185
R11417 VDD.n2012 VDD.n323 185
R11418 VDD.n1965 VDD.n1964 185
R11419 VDD.n1964 VDD.n322 185
R11420 VDD.n1963 VDD.n345 185
R11421 VDD.n1963 VDD.n1962 185
R11422 VDD.n1745 VDD.n346 185
R11423 VDD.n347 VDD.n346 185
R11424 VDD.n1746 VDD.n353 185
R11425 VDD.n1956 VDD.n353 185
R11426 VDD.n1748 VDD.n1747 185
R11427 VDD.n1747 VDD.n362 185
R11428 VDD.n1749 VDD.n360 185
R11429 VDD.n1920 VDD.n360 185
R11430 VDD.n1751 VDD.n1750 185
R11431 VDD.n1750 VDD.n359 185
R11432 VDD.n1752 VDD.n367 185
R11433 VDD.n1914 VDD.n367 185
R11434 VDD.n1754 VDD.n1753 185
R11435 VDD.n1753 VDD.n366 185
R11436 VDD.n1755 VDD.n373 185
R11437 VDD.n1908 VDD.n373 185
R11438 VDD.n1757 VDD.n1756 185
R11439 VDD.n1756 VDD.n372 185
R11440 VDD.n1758 VDD.n379 185
R11441 VDD.n1902 VDD.n379 185
R11442 VDD.n1760 VDD.n1759 185
R11443 VDD.n1759 VDD.n378 185
R11444 VDD.n1761 VDD.n385 185
R11445 VDD.n1896 VDD.n385 185
R11446 VDD.n1763 VDD.n1762 185
R11447 VDD.n1762 VDD.n384 185
R11448 VDD.n1764 VDD.n390 185
R11449 VDD.n1890 VDD.n390 185
R11450 VDD.n1766 VDD.n1765 185
R11451 VDD.n1765 VDD.n398 185
R11452 VDD.n1767 VDD.n396 185
R11453 VDD.n1884 VDD.n396 185
R11454 VDD.n1769 VDD.n1768 185
R11455 VDD.n1768 VDD.n395 185
R11456 VDD.n1770 VDD.n403 185
R11457 VDD.n1878 VDD.n403 185
R11458 VDD.n1772 VDD.n1771 185
R11459 VDD.n1771 VDD.n402 185
R11460 VDD.n1773 VDD.n408 185
R11461 VDD.n1872 VDD.n408 185
R11462 VDD.n1775 VDD.n1774 185
R11463 VDD.n1774 VDD.n416 185
R11464 VDD.n1776 VDD.n414 185
R11465 VDD.n1866 VDD.n414 185
R11466 VDD.n1778 VDD.n1777 185
R11467 VDD.n1777 VDD.n413 185
R11468 VDD.n1779 VDD.n421 185
R11469 VDD.n1860 VDD.n421 185
R11470 VDD.n1781 VDD.n1780 185
R11471 VDD.n1780 VDD.n420 185
R11472 VDD.n1782 VDD.n426 185
R11473 VDD.n1854 VDD.n426 185
R11474 VDD.n1784 VDD.n1783 185
R11475 VDD.n1783 VDD.n434 185
R11476 VDD.n1785 VDD.n432 185
R11477 VDD.n1848 VDD.n432 185
R11478 VDD.n1787 VDD.n1786 185
R11479 VDD.n1786 VDD.n431 185
R11480 VDD.n1788 VDD.n439 185
R11481 VDD.n1842 VDD.n439 185
R11482 VDD.n1790 VDD.n1789 185
R11483 VDD.n1789 VDD.n438 185
R11484 VDD.n1791 VDD.n1628 185
R11485 VDD.n1836 VDD.n1628 185
R11486 VDD.n1835 VDD.n1834 185
R11487 VDD.n1836 VDD.n1835 185
R11488 VDD.n437 VDD.n436 185
R11489 VDD.n438 VDD.n437 185
R11490 VDD.n1844 VDD.n1843 185
R11491 VDD.n1843 VDD.n1842 185
R11492 VDD.n1845 VDD.n435 185
R11493 VDD.n435 VDD.n431 185
R11494 VDD.n1847 VDD.n1846 185
R11495 VDD.n1848 VDD.n1847 185
R11496 VDD.n425 VDD.n424 185
R11497 VDD.n434 VDD.n425 185
R11498 VDD.n1856 VDD.n1855 185
R11499 VDD.n1855 VDD.n1854 185
R11500 VDD.n1857 VDD.n423 185
R11501 VDD.n423 VDD.n420 185
R11502 VDD.n1859 VDD.n1858 185
R11503 VDD.n1860 VDD.n1859 185
R11504 VDD.n412 VDD.n411 185
R11505 VDD.n413 VDD.n412 185
R11506 VDD.n1868 VDD.n1867 185
R11507 VDD.n1867 VDD.n1866 185
R11508 VDD.n1869 VDD.n410 185
R11509 VDD.n416 VDD.n410 185
R11510 VDD.n1871 VDD.n1870 185
R11511 VDD.n1872 VDD.n1871 185
R11512 VDD.n401 VDD.n400 185
R11513 VDD.n402 VDD.n401 185
R11514 VDD.n1880 VDD.n1879 185
R11515 VDD.n1879 VDD.n1878 185
R11516 VDD.n1881 VDD.n399 185
R11517 VDD.n399 VDD.n395 185
R11518 VDD.n1883 VDD.n1882 185
R11519 VDD.n1884 VDD.n1883 185
R11520 VDD.n389 VDD.n388 185
R11521 VDD.n398 VDD.n389 185
R11522 VDD.n1892 VDD.n1891 185
R11523 VDD.n1891 VDD.n1890 185
R11524 VDD.n1893 VDD.n387 185
R11525 VDD.n387 VDD.n384 185
R11526 VDD.n1895 VDD.n1894 185
R11527 VDD.n1896 VDD.n1895 185
R11528 VDD.n377 VDD.n376 185
R11529 VDD.n378 VDD.n377 185
R11530 VDD.n1904 VDD.n1903 185
R11531 VDD.n1903 VDD.n1902 185
R11532 VDD.n1905 VDD.n375 185
R11533 VDD.n375 VDD.n372 185
R11534 VDD.n1907 VDD.n1906 185
R11535 VDD.n1908 VDD.n1907 185
R11536 VDD.n365 VDD.n364 185
R11537 VDD.n366 VDD.n365 185
R11538 VDD.n1916 VDD.n1915 185
R11539 VDD.n1915 VDD.n1914 185
R11540 VDD.n1917 VDD.n363 185
R11541 VDD.n363 VDD.n359 185
R11542 VDD.n1919 VDD.n1918 185
R11543 VDD.n1920 VDD.n1919 185
R11544 VDD.n352 VDD.n351 185
R11545 VDD.n362 VDD.n352 185
R11546 VDD.n1958 VDD.n1957 185
R11547 VDD.n1957 VDD.n1956 185
R11548 VDD.n1959 VDD.n350 185
R11549 VDD.n350 VDD.n347 185
R11550 VDD.n1961 VDD.n1960 185
R11551 VDD.n1962 VDD.n1961 185
R11552 VDD.n328 VDD.n326 185
R11553 VDD.n326 VDD.n322 185
R11554 VDD.n2011 VDD.n2010 185
R11555 VDD.n2012 VDD.n2011 185
R11556 VDD.n2009 VDD.n327 185
R11557 VDD.n327 VDD.n324 185
R11558 VDD.n1571 VDD.n1570 185
R11559 VDD.n1570 VDD.n444 185
R11560 VDD.n1572 VDD.n477 185
R11561 VDD.n1582 VDD.n477 185
R11562 VDD.n1573 VDD.n485 185
R11563 VDD.n485 VDD.n475 185
R11564 VDD.n1575 VDD.n1574 185
R11565 VDD.n1576 VDD.n1575 185
R11566 VDD.n486 VDD.n484 185
R11567 VDD.n484 VDD.n481 185
R11568 VDD.n1508 VDD.n492 185
R11569 VDD.n1518 VDD.n492 185
R11570 VDD.n1509 VDD.n501 185
R11571 VDD.n501 VDD.n499 185
R11572 VDD.n1511 VDD.n1510 185
R11573 VDD.n1512 VDD.n1511 185
R11574 VDD.n1507 VDD.n500 185
R11575 VDD.n500 VDD.n496 185
R11576 VDD.n1506 VDD.n1505 185
R11577 VDD.n1505 VDD.n1504 185
R11578 VDD.n503 VDD.n502 185
R11579 VDD.n504 VDD.n503 185
R11580 VDD.n1497 VDD.n1496 185
R11581 VDD.n1498 VDD.n1497 185
R11582 VDD.n1495 VDD.n512 185
R11583 VDD.n518 VDD.n512 185
R11584 VDD.n1494 VDD.n1493 185
R11585 VDD.n1493 VDD.n1492 185
R11586 VDD.n514 VDD.n513 185
R11587 VDD.n515 VDD.n514 185
R11588 VDD.n1485 VDD.n1484 185
R11589 VDD.n1486 VDD.n1485 185
R11590 VDD.n1483 VDD.n525 185
R11591 VDD.n525 VDD.n522 185
R11592 VDD.n1482 VDD.n1481 185
R11593 VDD.n1481 VDD.n1480 185
R11594 VDD.n527 VDD.n526 185
R11595 VDD.n536 VDD.n527 185
R11596 VDD.n1473 VDD.n1472 185
R11597 VDD.n1474 VDD.n1473 185
R11598 VDD.n1471 VDD.n537 185
R11599 VDD.n537 VDD.n533 185
R11600 VDD.n1470 VDD.n1469 185
R11601 VDD.n1469 VDD.n1468 185
R11602 VDD.n539 VDD.n538 185
R11603 VDD.n540 VDD.n539 185
R11604 VDD.n1461 VDD.n1460 185
R11605 VDD.n1462 VDD.n1461 185
R11606 VDD.n1459 VDD.n549 185
R11607 VDD.n549 VDD.n546 185
R11608 VDD.n1458 VDD.n1457 185
R11609 VDD.n1457 VDD.n1456 185
R11610 VDD.n551 VDD.n550 185
R11611 VDD.n552 VDD.n551 185
R11612 VDD.n1449 VDD.n1448 185
R11613 VDD.n1450 VDD.n1449 185
R11614 VDD.n1447 VDD.n561 185
R11615 VDD.n561 VDD.n558 185
R11616 VDD.n1446 VDD.n1445 185
R11617 VDD.n1445 VDD.n1444 185
R11618 VDD.n563 VDD.n562 185
R11619 VDD.n572 VDD.n563 185
R11620 VDD.n1437 VDD.n1436 185
R11621 VDD.n1438 VDD.n1437 185
R11622 VDD.n1435 VDD.n573 185
R11623 VDD.n573 VDD.n569 185
R11624 VDD.n1434 VDD.n1433 185
R11625 VDD.n1433 VDD.n1432 185
R11626 VDD.n575 VDD.n574 185
R11627 VDD.n576 VDD.n575 185
R11628 VDD.n1425 VDD.n1424 185
R11629 VDD.n1426 VDD.n1425 185
R11630 VDD.n1528 VDD.n455 185
R11631 VDD.n1626 VDD.n455 185
R11632 VDD.n1530 VDD.n1529 185
R11633 VDD.n1533 VDD.n1532 185
R11634 VDD.n1535 VDD.n1534 185
R11635 VDD.n1537 VDD.n1536 185
R11636 VDD.n1539 VDD.n1538 185
R11637 VDD.n1541 VDD.n1540 185
R11638 VDD.n1543 VDD.n1542 185
R11639 VDD.n1545 VDD.n1544 185
R11640 VDD.n1547 VDD.n1546 185
R11641 VDD.n1549 VDD.n1548 185
R11642 VDD.n1551 VDD.n1550 185
R11643 VDD.n1553 VDD.n1552 185
R11644 VDD.n1555 VDD.n1554 185
R11645 VDD.n1557 VDD.n1556 185
R11646 VDD.n1559 VDD.n1558 185
R11647 VDD.n1561 VDD.n1560 185
R11648 VDD.n1563 VDD.n1562 185
R11649 VDD.n1565 VDD.n1564 185
R11650 VDD.n1567 VDD.n1566 185
R11651 VDD.n1569 VDD.n1568 185
R11652 VDD.n1527 VDD.n1526 185
R11653 VDD.n1526 VDD.n444 185
R11654 VDD.n1525 VDD.n476 185
R11655 VDD.n1582 VDD.n476 185
R11656 VDD.n1524 VDD.n1523 185
R11657 VDD.n1523 VDD.n475 185
R11658 VDD.n1522 VDD.n483 185
R11659 VDD.n1576 VDD.n483 185
R11660 VDD.n1521 VDD.n1520 185
R11661 VDD.n1520 VDD.n481 185
R11662 VDD.n1519 VDD.n489 185
R11663 VDD.n1519 VDD.n1518 185
R11664 VDD.n1339 VDD.n490 185
R11665 VDD.n499 VDD.n490 185
R11666 VDD.n1340 VDD.n498 185
R11667 VDD.n1512 VDD.n498 185
R11668 VDD.n1342 VDD.n1341 185
R11669 VDD.n1341 VDD.n496 185
R11670 VDD.n1343 VDD.n506 185
R11671 VDD.n1504 VDD.n506 185
R11672 VDD.n1345 VDD.n1344 185
R11673 VDD.n1344 VDD.n504 185
R11674 VDD.n1346 VDD.n511 185
R11675 VDD.n1498 VDD.n511 185
R11676 VDD.n1348 VDD.n1347 185
R11677 VDD.n1347 VDD.n518 185
R11678 VDD.n1349 VDD.n517 185
R11679 VDD.n1492 VDD.n517 185
R11680 VDD.n1351 VDD.n1350 185
R11681 VDD.n1350 VDD.n515 185
R11682 VDD.n1352 VDD.n524 185
R11683 VDD.n1486 VDD.n524 185
R11684 VDD.n1354 VDD.n1353 185
R11685 VDD.n1353 VDD.n522 185
R11686 VDD.n1355 VDD.n529 185
R11687 VDD.n1480 VDD.n529 185
R11688 VDD.n1357 VDD.n1356 185
R11689 VDD.n1356 VDD.n536 185
R11690 VDD.n1358 VDD.n535 185
R11691 VDD.n1474 VDD.n535 185
R11692 VDD.n1360 VDD.n1359 185
R11693 VDD.n1359 VDD.n533 185
R11694 VDD.n1361 VDD.n542 185
R11695 VDD.n1468 VDD.n542 185
R11696 VDD.n1363 VDD.n1362 185
R11697 VDD.n1362 VDD.n540 185
R11698 VDD.n1364 VDD.n548 185
R11699 VDD.n1462 VDD.n548 185
R11700 VDD.n1366 VDD.n1365 185
R11701 VDD.n1365 VDD.n546 185
R11702 VDD.n1367 VDD.n554 185
R11703 VDD.n1456 VDD.n554 185
R11704 VDD.n1369 VDD.n1368 185
R11705 VDD.n1368 VDD.n552 185
R11706 VDD.n1370 VDD.n560 185
R11707 VDD.n1450 VDD.n560 185
R11708 VDD.n1372 VDD.n1371 185
R11709 VDD.n1371 VDD.n558 185
R11710 VDD.n1373 VDD.n565 185
R11711 VDD.n1444 VDD.n565 185
R11712 VDD.n1375 VDD.n1374 185
R11713 VDD.n1374 VDD.n572 185
R11714 VDD.n1376 VDD.n571 185
R11715 VDD.n1438 VDD.n571 185
R11716 VDD.n1378 VDD.n1377 185
R11717 VDD.n1377 VDD.n569 185
R11718 VDD.n1379 VDD.n578 185
R11719 VDD.n1432 VDD.n578 185
R11720 VDD.n1381 VDD.n1380 185
R11721 VDD.n1380 VDD.n576 185
R11722 VDD.n1382 VDD.n584 185
R11723 VDD.n1426 VDD.n584 185
R11724 VDD.n1423 VDD.n585 185
R11725 VDD.n1422 VDD.n1421 185
R11726 VDD.n1419 VDD.n586 185
R11727 VDD.n1417 VDD.n1416 185
R11728 VDD.n1415 VDD.n587 185
R11729 VDD.n1414 VDD.n1413 185
R11730 VDD.n1411 VDD.n588 185
R11731 VDD.n1409 VDD.n1408 185
R11732 VDD.n1407 VDD.n589 185
R11733 VDD.n1406 VDD.n1405 185
R11734 VDD.n1403 VDD.n1330 185
R11735 VDD.n1401 VDD.n1400 185
R11736 VDD.n1399 VDD.n1331 185
R11737 VDD.n1398 VDD.n1397 185
R11738 VDD.n1395 VDD.n1332 185
R11739 VDD.n1393 VDD.n1392 185
R11740 VDD.n1391 VDD.n1333 185
R11741 VDD.n1390 VDD.n1389 185
R11742 VDD.n1387 VDD.n1334 185
R11743 VDD.n1385 VDD.n1384 185
R11744 VDD.n1383 VDD.n1335 185
R11745 VDD.n1335 VDD.n582 185
R11746 VDD.n1336 VDD.t71 178.127
R11747 VDD.n487 VDD.t11 178.127
R11748 VDD.n1228 VDD.t77 178.127
R11749 VDD.n469 VDD.t60 178.127
R11750 VDD.n1631 VDD.t4 178.127
R11751 VDD.n343 VDD.t45 178.127
R11752 VDD.n1743 VDD.t15 178.127
R11753 VDD.n314 VDD.t54 178.127
R11754 VDD.n831 VDD.t23 177.585
R11755 VDD.n851 VDD.t42 177.585
R11756 VDD.n872 VDD.t67 177.585
R11757 VDD.n893 VDD.t49 177.585
R11758 VDD.n598 VDD.t7 177.585
R11759 VDD.n1141 VDD.t32 177.585
R11760 VDD.n1165 VDD.t57 177.585
R11761 VDD.n1189 VDD.t35 177.585
R11762 VDD.n171 VDD.t73 177.585
R11763 VDD.n2271 VDD.t26 177.585
R11764 VDD.n2295 VDD.t38 177.585
R11765 VDD.n2319 VDD.t79 177.585
R11766 VDD.n2069 VDD.t52 177.585
R11767 VDD.n2096 VDD.t19 177.585
R11768 VDD.n2123 VDD.t64 177.585
R11769 VDD.n2045 VDD.t30 177.585
R11770 VDD.n91 VDD.n88 146.341
R11771 VDD.n2334 VDD.n2333 146.341
R11772 VDD.n2331 VDD.n95 146.341
R11773 VDD.n2327 VDD.n2326 146.341
R11774 VDD.n2324 VDD.n102 146.341
R11775 VDD.n2317 VDD.n2316 146.341
R11776 VDD.n2314 VDD.n109 146.341
R11777 VDD.n2310 VDD.n2309 146.341
R11778 VDD.n2307 VDD.n116 146.341
R11779 VDD.n2303 VDD.n2302 146.341
R11780 VDD.n2300 VDD.n123 146.341
R11781 VDD.n2293 VDD.n2292 146.341
R11782 VDD.n2290 VDD.n130 146.341
R11783 VDD.n2286 VDD.n2285 146.341
R11784 VDD.n2283 VDD.n137 146.341
R11785 VDD.n2279 VDD.n2278 146.341
R11786 VDD.n2276 VDD.n144 146.341
R11787 VDD.n2269 VDD.n2268 146.341
R11788 VDD.n2266 VDD.n151 146.341
R11789 VDD.n2262 VDD.n2261 146.341
R11790 VDD.n2259 VDD.n158 146.341
R11791 VDD.n2255 VDD.n2254 146.341
R11792 VDD.n2252 VDD.n165 146.341
R11793 VDD.n2151 VDD.n238 146.341
R11794 VDD.n2151 VDD.n234 146.341
R11795 VDD.n2157 VDD.n234 146.341
R11796 VDD.n2157 VDD.n227 146.341
R11797 VDD.n2167 VDD.n227 146.341
R11798 VDD.n2167 VDD.n223 146.341
R11799 VDD.n2173 VDD.n223 146.341
R11800 VDD.n2173 VDD.n215 146.341
R11801 VDD.n2183 VDD.n215 146.341
R11802 VDD.n2183 VDD.n211 146.341
R11803 VDD.n2189 VDD.n211 146.341
R11804 VDD.n2189 VDD.n203 146.341
R11805 VDD.n2199 VDD.n203 146.341
R11806 VDD.n2199 VDD.n199 146.341
R11807 VDD.n2205 VDD.n199 146.341
R11808 VDD.n2205 VDD.n189 146.341
R11809 VDD.n2215 VDD.n189 146.341
R11810 VDD.n2215 VDD.n190 146.341
R11811 VDD.n190 VDD.n41 146.341
R11812 VDD.n42 VDD.n41 146.341
R11813 VDD.n43 VDD.n42 146.341
R11814 VDD.n183 VDD.n43 146.341
R11815 VDD.n183 VDD.n51 146.341
R11816 VDD.n52 VDD.n51 146.341
R11817 VDD.n53 VDD.n52 146.341
R11818 VDD.n180 VDD.n53 146.341
R11819 VDD.n180 VDD.n62 146.341
R11820 VDD.n63 VDD.n62 146.341
R11821 VDD.n64 VDD.n63 146.341
R11822 VDD.n177 VDD.n64 146.341
R11823 VDD.n177 VDD.n73 146.341
R11824 VDD.n74 VDD.n73 146.341
R11825 VDD.n75 VDD.n74 146.341
R11826 VDD.n174 VDD.n75 146.341
R11827 VDD.n174 VDD.n84 146.341
R11828 VDD.n85 VDD.n84 146.341
R11829 VDD.n86 VDD.n85 146.341
R11830 VDD.n2140 VDD.n245 146.341
R11831 VDD.n2140 VDD.n268 146.341
R11832 VDD.n2136 VDD.n2135 146.341
R11833 VDD.n2132 VDD.n2131 146.341
R11834 VDD.n2128 VDD.n2127 146.341
R11835 VDD.n2121 VDD.n2120 146.341
R11836 VDD.n2117 VDD.n2116 146.341
R11837 VDD.n2113 VDD.n2112 146.341
R11838 VDD.n2109 VDD.n2108 146.341
R11839 VDD.n2105 VDD.n2104 146.341
R11840 VDD.n2101 VDD.n2100 146.341
R11841 VDD.n2094 VDD.n2093 146.341
R11842 VDD.n2090 VDD.n2089 146.341
R11843 VDD.n2086 VDD.n2085 146.341
R11844 VDD.n2082 VDD.n2081 146.341
R11845 VDD.n2078 VDD.n2077 146.341
R11846 VDD.n2074 VDD.n2073 146.341
R11847 VDD.n2067 VDD.n2066 146.341
R11848 VDD.n2063 VDD.n2062 146.341
R11849 VDD.n2059 VDD.n2058 146.341
R11850 VDD.n2037 VDD.n2036 146.341
R11851 VDD.n2051 VDD.n2039 146.341
R11852 VDD.n2049 VDD.n2048 146.341
R11853 VDD.n2149 VDD.n241 146.341
R11854 VDD.n2149 VDD.n233 146.341
R11855 VDD.n2159 VDD.n233 146.341
R11856 VDD.n2159 VDD.n229 146.341
R11857 VDD.n2165 VDD.n229 146.341
R11858 VDD.n2165 VDD.n221 146.341
R11859 VDD.n2175 VDD.n221 146.341
R11860 VDD.n2175 VDD.n217 146.341
R11861 VDD.n2181 VDD.n217 146.341
R11862 VDD.n2181 VDD.n209 146.341
R11863 VDD.n2191 VDD.n209 146.341
R11864 VDD.n2191 VDD.n205 146.341
R11865 VDD.n2197 VDD.n205 146.341
R11866 VDD.n2197 VDD.n197 146.341
R11867 VDD.n2207 VDD.n197 146.341
R11868 VDD.n2207 VDD.n193 146.341
R11869 VDD.n2213 VDD.n193 146.341
R11870 VDD.n2213 VDD.n39 146.341
R11871 VDD.n2377 VDD.n39 146.341
R11872 VDD.n2377 VDD.n40 146.341
R11873 VDD.n2373 VDD.n40 146.341
R11874 VDD.n2373 VDD.n45 146.341
R11875 VDD.n2369 VDD.n45 146.341
R11876 VDD.n2369 VDD.n50 146.341
R11877 VDD.n2365 VDD.n50 146.341
R11878 VDD.n2365 VDD.n55 146.341
R11879 VDD.n2361 VDD.n55 146.341
R11880 VDD.n2361 VDD.n61 146.341
R11881 VDD.n2357 VDD.n61 146.341
R11882 VDD.n2357 VDD.n66 146.341
R11883 VDD.n2353 VDD.n66 146.341
R11884 VDD.n2353 VDD.n72 146.341
R11885 VDD.n2349 VDD.n72 146.341
R11886 VDD.n2349 VDD.n77 146.341
R11887 VDD.n2345 VDD.n77 146.341
R11888 VDD.n2345 VDD.n83 146.341
R11889 VDD.n2341 VDD.n83 146.341
R11890 VDD.n1313 VDD.n607 146.341
R11891 VDD.n1311 VDD.n1310 146.341
R11892 VDD.n1308 VDD.n1066 146.341
R11893 VDD.n1197 VDD.n1196 146.341
R11894 VDD.n1194 VDD.n1071 146.341
R11895 VDD.n1187 VDD.n1186 146.341
R11896 VDD.n1184 VDD.n1076 146.341
R11897 VDD.n1180 VDD.n1179 146.341
R11898 VDD.n1177 VDD.n1083 146.341
R11899 VDD.n1173 VDD.n1172 146.341
R11900 VDD.n1170 VDD.n1090 146.341
R11901 VDD.n1163 VDD.n1162 146.341
R11902 VDD.n1160 VDD.n1097 146.341
R11903 VDD.n1156 VDD.n1155 146.341
R11904 VDD.n1153 VDD.n1104 146.341
R11905 VDD.n1149 VDD.n1148 146.341
R11906 VDD.n1146 VDD.n1111 146.341
R11907 VDD.n1139 VDD.n1138 146.341
R11908 VDD.n1136 VDD.n1118 146.341
R11909 VDD.n1132 VDD.n1131 146.341
R11910 VDD.n1129 VDD.n1126 146.341
R11911 VDD.n1124 VDD.n595 146.341
R11912 VDD.n1324 VDD.n596 146.341
R11913 VDD.n919 VDD.n733 146.341
R11914 VDD.n919 VDD.n729 146.341
R11915 VDD.n925 VDD.n729 146.341
R11916 VDD.n925 VDD.n722 146.341
R11917 VDD.n935 VDD.n722 146.341
R11918 VDD.n935 VDD.n718 146.341
R11919 VDD.n941 VDD.n718 146.341
R11920 VDD.n941 VDD.n710 146.341
R11921 VDD.n951 VDD.n710 146.341
R11922 VDD.n951 VDD.n706 146.341
R11923 VDD.n957 VDD.n706 146.341
R11924 VDD.n957 VDD.n698 146.341
R11925 VDD.n967 VDD.n698 146.341
R11926 VDD.n967 VDD.n694 146.341
R11927 VDD.n973 VDD.n694 146.341
R11928 VDD.n973 VDD.n685 146.341
R11929 VDD.n984 VDD.n685 146.341
R11930 VDD.n984 VDD.n681 146.341
R11931 VDD.n990 VDD.n681 146.341
R11932 VDD.n990 VDD.n654 146.341
R11933 VDD.n1000 VDD.n654 146.341
R11934 VDD.n1000 VDD.n650 146.341
R11935 VDD.n1006 VDD.n650 146.341
R11936 VDD.n1006 VDD.n642 146.341
R11937 VDD.n1016 VDD.n642 146.341
R11938 VDD.n1016 VDD.n638 146.341
R11939 VDD.n1022 VDD.n638 146.341
R11940 VDD.n1022 VDD.n630 146.341
R11941 VDD.n1032 VDD.n630 146.341
R11942 VDD.n1032 VDD.n626 146.341
R11943 VDD.n1038 VDD.n626 146.341
R11944 VDD.n1038 VDD.n617 146.341
R11945 VDD.n1048 VDD.n617 146.341
R11946 VDD.n1048 VDD.n612 146.341
R11947 VDD.n1057 VDD.n612 146.341
R11948 VDD.n1057 VDD.n603 146.341
R11949 VDD.n1321 VDD.n603 146.341
R11950 VDD.n908 VDD.n740 146.341
R11951 VDD.n908 VDD.n763 146.341
R11952 VDD.n767 VDD.n766 146.341
R11953 VDD.n769 VDD.n768 146.341
R11954 VDD.n773 VDD.n772 146.341
R11955 VDD.n775 VDD.n774 146.341
R11956 VDD.n779 VDD.n778 146.341
R11957 VDD.n781 VDD.n780 146.341
R11958 VDD.n785 VDD.n784 146.341
R11959 VDD.n787 VDD.n786 146.341
R11960 VDD.n791 VDD.n790 146.341
R11961 VDD.n793 VDD.n792 146.341
R11962 VDD.n797 VDD.n796 146.341
R11963 VDD.n799 VDD.n798 146.341
R11964 VDD.n803 VDD.n802 146.341
R11965 VDD.n805 VDD.n804 146.341
R11966 VDD.n809 VDD.n808 146.341
R11967 VDD.n811 VDD.n810 146.341
R11968 VDD.n815 VDD.n814 146.341
R11969 VDD.n817 VDD.n816 146.341
R11970 VDD.n821 VDD.n820 146.341
R11971 VDD.n823 VDD.n822 146.341
R11972 VDD.n830 VDD.n826 146.341
R11973 VDD.n917 VDD.n736 146.341
R11974 VDD.n917 VDD.n728 146.341
R11975 VDD.n927 VDD.n728 146.341
R11976 VDD.n927 VDD.n724 146.341
R11977 VDD.n933 VDD.n724 146.341
R11978 VDD.n933 VDD.n716 146.341
R11979 VDD.n943 VDD.n716 146.341
R11980 VDD.n943 VDD.n712 146.341
R11981 VDD.n949 VDD.n712 146.341
R11982 VDD.n949 VDD.n704 146.341
R11983 VDD.n959 VDD.n704 146.341
R11984 VDD.n959 VDD.n700 146.341
R11985 VDD.n965 VDD.n700 146.341
R11986 VDD.n965 VDD.n692 146.341
R11987 VDD.n975 VDD.n692 146.341
R11988 VDD.n975 VDD.n688 146.341
R11989 VDD.n982 VDD.n688 146.341
R11990 VDD.n982 VDD.n680 146.341
R11991 VDD.n992 VDD.n680 146.341
R11992 VDD.n992 VDD.n656 146.341
R11993 VDD.n998 VDD.n656 146.341
R11994 VDD.n998 VDD.n648 146.341
R11995 VDD.n1008 VDD.n648 146.341
R11996 VDD.n1008 VDD.n644 146.341
R11997 VDD.n1014 VDD.n644 146.341
R11998 VDD.n1014 VDD.n636 146.341
R11999 VDD.n1024 VDD.n636 146.341
R12000 VDD.n1024 VDD.n632 146.341
R12001 VDD.n1030 VDD.n632 146.341
R12002 VDD.n1030 VDD.n624 146.341
R12003 VDD.n1040 VDD.n624 146.341
R12004 VDD.n1040 VDD.n620 146.341
R12005 VDD.n1046 VDD.n620 146.341
R12006 VDD.n1046 VDD.n611 146.341
R12007 VDD.n1059 VDD.n611 146.341
R12008 VDD.n1059 VDD.n606 146.341
R12009 VDD.n1319 VDD.n606 146.341
R12010 VDD.t0 VDD.t138 145.315
R12011 VDD.t105 VDD.t81 145.315
R12012 VDD.n832 VDD.t22 132.203
R12013 VDD.n852 VDD.t41 132.203
R12014 VDD.n873 VDD.t66 132.203
R12015 VDD.n894 VDD.t48 132.203
R12016 VDD.n599 VDD.t8 132.203
R12017 VDD.n1142 VDD.t33 132.203
R12018 VDD.n1166 VDD.t58 132.203
R12019 VDD.n1190 VDD.t36 132.203
R12020 VDD.n172 VDD.t74 132.203
R12021 VDD.n2272 VDD.t27 132.203
R12022 VDD.n2296 VDD.t39 132.203
R12023 VDD.n2320 VDD.t80 132.203
R12024 VDD.n2070 VDD.t51 132.203
R12025 VDD.n2097 VDD.t18 132.203
R12026 VDD.n2124 VDD.t63 132.203
R12027 VDD.n2046 VDD.t29 132.203
R12028 VDD.n1627 VDD.n1626 127.722
R12029 VDD.n1337 VDD.t70 119.169
R12030 VDD.n488 VDD.t12 119.169
R12031 VDD.n1229 VDD.t76 119.169
R12032 VDD.n470 VDD.t61 119.169
R12033 VDD.n1632 VDD.t3 119.169
R12034 VDD.n344 VDD.t46 119.169
R12035 VDD.n1744 VDD.t14 119.169
R12036 VDD.n315 VDD.t55 119.169
R12037 VDD.n673 VDD.t143 112.609
R12038 VDD.n668 VDD.t165 112.609
R12039 VDD.n663 VDD.t114 112.609
R12040 VDD.n659 VDD.t87 112.609
R12041 VDD.n33 VDD.t157 110.591
R12042 VDD.n28 VDD.t109 110.591
R12043 VDD.n23 VDD.t158 110.591
R12044 VDD.n19 VDD.t141 110.591
R12045 VDD.t138 VDD.t119 106.963
R12046 VDD.t119 VDD.t103 106.963
R12047 VDD.t103 VDD.t162 106.963
R12048 VDD.t144 VDD.t127 106.963
R12049 VDD.t127 VDD.t84 106.963
R12050 VDD.t84 VDD.t105 106.963
R12051 VDD.n9 VDD.n7 104.614
R12052 VDD.n2 VDD.n0 104.614
R12053 VDD.n32 VDD.n30 103.871
R12054 VDD.n27 VDD.n25 103.871
R12055 VDD.n22 VDD.n20 103.871
R12056 VDD.n18 VDD.n16 103.871
R12057 VDD.n9 VDD.n8 101.993
R12058 VDD.n11 VDD.n10 101.993
R12059 VDD.n13 VDD.n12 101.993
R12060 VDD.n6 VDD.n5 101.993
R12061 VDD.n4 VDD.n3 101.993
R12062 VDD.n2 VDD.n1 101.993
R12063 VDD.n32 VDD.n31 101.853
R12064 VDD.n27 VDD.n26 101.853
R12065 VDD.n22 VDD.n21 101.853
R12066 VDD.n18 VDD.n17 101.853
R12067 VDD.n673 VDD.n672 101.853
R12068 VDD.n675 VDD.n674 101.853
R12069 VDD.n668 VDD.n667 101.853
R12070 VDD.n670 VDD.n669 101.853
R12071 VDD.n663 VDD.n662 101.853
R12072 VDD.n665 VDD.n664 101.853
R12073 VDD.n659 VDD.n658 101.853
R12074 VDD.n661 VDD.n660 101.853
R12075 VDD.n1835 VDD.n437 99.5127
R12076 VDD.n1843 VDD.n437 99.5127
R12077 VDD.n1843 VDD.n435 99.5127
R12078 VDD.n1847 VDD.n435 99.5127
R12079 VDD.n1847 VDD.n425 99.5127
R12080 VDD.n1855 VDD.n425 99.5127
R12081 VDD.n1855 VDD.n423 99.5127
R12082 VDD.n1859 VDD.n423 99.5127
R12083 VDD.n1859 VDD.n412 99.5127
R12084 VDD.n1867 VDD.n412 99.5127
R12085 VDD.n1867 VDD.n410 99.5127
R12086 VDD.n1871 VDD.n410 99.5127
R12087 VDD.n1871 VDD.n401 99.5127
R12088 VDD.n1879 VDD.n401 99.5127
R12089 VDD.n1879 VDD.n399 99.5127
R12090 VDD.n1883 VDD.n399 99.5127
R12091 VDD.n1883 VDD.n389 99.5127
R12092 VDD.n1891 VDD.n389 99.5127
R12093 VDD.n1891 VDD.n387 99.5127
R12094 VDD.n1895 VDD.n387 99.5127
R12095 VDD.n1895 VDD.n377 99.5127
R12096 VDD.n1903 VDD.n377 99.5127
R12097 VDD.n1903 VDD.n375 99.5127
R12098 VDD.n1907 VDD.n375 99.5127
R12099 VDD.n1907 VDD.n365 99.5127
R12100 VDD.n1915 VDD.n365 99.5127
R12101 VDD.n1915 VDD.n363 99.5127
R12102 VDD.n1919 VDD.n363 99.5127
R12103 VDD.n1919 VDD.n352 99.5127
R12104 VDD.n1957 VDD.n352 99.5127
R12105 VDD.n1957 VDD.n350 99.5127
R12106 VDD.n1961 VDD.n350 99.5127
R12107 VDD.n1961 VDD.n326 99.5127
R12108 VDD.n2011 VDD.n326 99.5127
R12109 VDD.n2011 VDD.n327 99.5127
R12110 VDD.n2007 VDD.n2006 99.5127
R12111 VDD.n2004 VDD.n330 99.5127
R12112 VDD.n2000 VDD.n1999 99.5127
R12113 VDD.n1997 VDD.n333 99.5127
R12114 VDD.n1993 VDD.n1992 99.5127
R12115 VDD.n1990 VDD.n336 99.5127
R12116 VDD.n1985 VDD.n1984 99.5127
R12117 VDD.n1982 VDD.n339 99.5127
R12118 VDD.n1978 VDD.n1977 99.5127
R12119 VDD.n1975 VDD.n342 99.5127
R12120 VDD.n1789 VDD.n1628 99.5127
R12121 VDD.n1789 VDD.n439 99.5127
R12122 VDD.n1786 VDD.n439 99.5127
R12123 VDD.n1786 VDD.n432 99.5127
R12124 VDD.n1783 VDD.n432 99.5127
R12125 VDD.n1783 VDD.n426 99.5127
R12126 VDD.n1780 VDD.n426 99.5127
R12127 VDD.n1780 VDD.n421 99.5127
R12128 VDD.n1777 VDD.n421 99.5127
R12129 VDD.n1777 VDD.n414 99.5127
R12130 VDD.n1774 VDD.n414 99.5127
R12131 VDD.n1774 VDD.n408 99.5127
R12132 VDD.n1771 VDD.n408 99.5127
R12133 VDD.n1771 VDD.n403 99.5127
R12134 VDD.n1768 VDD.n403 99.5127
R12135 VDD.n1768 VDD.n396 99.5127
R12136 VDD.n1765 VDD.n396 99.5127
R12137 VDD.n1765 VDD.n390 99.5127
R12138 VDD.n1762 VDD.n390 99.5127
R12139 VDD.n1762 VDD.n385 99.5127
R12140 VDD.n1759 VDD.n385 99.5127
R12141 VDD.n1759 VDD.n379 99.5127
R12142 VDD.n1756 VDD.n379 99.5127
R12143 VDD.n1756 VDD.n373 99.5127
R12144 VDD.n1753 VDD.n373 99.5127
R12145 VDD.n1753 VDD.n367 99.5127
R12146 VDD.n1750 VDD.n367 99.5127
R12147 VDD.n1750 VDD.n360 99.5127
R12148 VDD.n1747 VDD.n360 99.5127
R12149 VDD.n1747 VDD.n353 99.5127
R12150 VDD.n353 VDD.n346 99.5127
R12151 VDD.n1963 VDD.n346 99.5127
R12152 VDD.n1964 VDD.n1963 99.5127
R12153 VDD.n1964 VDD.n323 99.5127
R12154 VDD.n1969 VDD.n323 99.5127
R12155 VDD.n1831 VDD.n1829 99.5127
R12156 VDD.n1829 VDD.n1828 99.5127
R12157 VDD.n1825 VDD.n1824 99.5127
R12158 VDD.n1822 VDD.n1736 99.5127
R12159 VDD.n1818 VDD.n1816 99.5127
R12160 VDD.n1814 VDD.n1738 99.5127
R12161 VDD.n1810 VDD.n1808 99.5127
R12162 VDD.n1806 VDD.n1740 99.5127
R12163 VDD.n1802 VDD.n1800 99.5127
R12164 VDD.n1798 VDD.n1742 99.5127
R12165 VDD.n1625 VDD.n467 99.5127
R12166 VDD.n1621 VDD.n1620 99.5127
R12167 VDD.n1617 VDD.n1616 99.5127
R12168 VDD.n1613 VDD.n1612 99.5127
R12169 VDD.n1609 VDD.n1608 99.5127
R12170 VDD.n1605 VDD.n1604 99.5127
R12171 VDD.n1601 VDD.n1600 99.5127
R12172 VDD.n1597 VDD.n1596 99.5127
R12173 VDD.n1593 VDD.n1592 99.5127
R12174 VDD.n1589 VDD.n1588 99.5127
R12175 VDD.n1279 VDD.n583 99.5127
R12176 VDD.n1279 VDD.n577 99.5127
R12177 VDD.n1276 VDD.n577 99.5127
R12178 VDD.n1276 VDD.n570 99.5127
R12179 VDD.n1273 VDD.n570 99.5127
R12180 VDD.n1273 VDD.n564 99.5127
R12181 VDD.n1270 VDD.n564 99.5127
R12182 VDD.n1270 VDD.n559 99.5127
R12183 VDD.n1267 VDD.n559 99.5127
R12184 VDD.n1267 VDD.n553 99.5127
R12185 VDD.n1264 VDD.n553 99.5127
R12186 VDD.n1264 VDD.n547 99.5127
R12187 VDD.n1261 VDD.n547 99.5127
R12188 VDD.n1261 VDD.n541 99.5127
R12189 VDD.n1258 VDD.n541 99.5127
R12190 VDD.n1258 VDD.n534 99.5127
R12191 VDD.n1255 VDD.n534 99.5127
R12192 VDD.n1255 VDD.n528 99.5127
R12193 VDD.n1252 VDD.n528 99.5127
R12194 VDD.n1252 VDD.n523 99.5127
R12195 VDD.n1249 VDD.n523 99.5127
R12196 VDD.n1249 VDD.n516 99.5127
R12197 VDD.n1246 VDD.n516 99.5127
R12198 VDD.n1246 VDD.n510 99.5127
R12199 VDD.n1243 VDD.n510 99.5127
R12200 VDD.n1243 VDD.n505 99.5127
R12201 VDD.n1240 VDD.n505 99.5127
R12202 VDD.n1240 VDD.n497 99.5127
R12203 VDD.n1237 VDD.n497 99.5127
R12204 VDD.n1237 VDD.n491 99.5127
R12205 VDD.n1234 VDD.n491 99.5127
R12206 VDD.n1234 VDD.n482 99.5127
R12207 VDD.n482 VDD.n473 99.5127
R12208 VDD.n1583 VDD.n473 99.5127
R12209 VDD.n1584 VDD.n1583 99.5127
R12210 VDD.n1206 VDD.n1204 99.5127
R12211 VDD.n1210 VDD.n1204 99.5127
R12212 VDD.n1214 VDD.n1212 99.5127
R12213 VDD.n1218 VDD.n1202 99.5127
R12214 VDD.n1221 VDD.n1220 99.5127
R12215 VDD.n1300 VDD.n1223 99.5127
R12216 VDD.n1298 VDD.n1297 99.5127
R12217 VDD.n1294 VDD.n1293 99.5127
R12218 VDD.n1291 VDD.n1227 99.5127
R12219 VDD.n1287 VDD.n1285 99.5127
R12220 VDD.n1427 VDD.n579 99.5127
R12221 VDD.n1431 VDD.n579 99.5127
R12222 VDD.n1431 VDD.n568 99.5127
R12223 VDD.n1439 VDD.n568 99.5127
R12224 VDD.n1439 VDD.n566 99.5127
R12225 VDD.n1443 VDD.n566 99.5127
R12226 VDD.n1443 VDD.n557 99.5127
R12227 VDD.n1451 VDD.n557 99.5127
R12228 VDD.n1451 VDD.n555 99.5127
R12229 VDD.n1455 VDD.n555 99.5127
R12230 VDD.n1455 VDD.n545 99.5127
R12231 VDD.n1463 VDD.n545 99.5127
R12232 VDD.n1463 VDD.n543 99.5127
R12233 VDD.n1467 VDD.n543 99.5127
R12234 VDD.n1467 VDD.n532 99.5127
R12235 VDD.n1475 VDD.n532 99.5127
R12236 VDD.n1475 VDD.n530 99.5127
R12237 VDD.n1479 VDD.n530 99.5127
R12238 VDD.n1479 VDD.n521 99.5127
R12239 VDD.n1487 VDD.n521 99.5127
R12240 VDD.n1487 VDD.n519 99.5127
R12241 VDD.n1491 VDD.n519 99.5127
R12242 VDD.n1491 VDD.n509 99.5127
R12243 VDD.n1499 VDD.n509 99.5127
R12244 VDD.n1499 VDD.n507 99.5127
R12245 VDD.n1503 VDD.n507 99.5127
R12246 VDD.n1503 VDD.n495 99.5127
R12247 VDD.n1513 VDD.n495 99.5127
R12248 VDD.n1513 VDD.n493 99.5127
R12249 VDD.n1517 VDD.n493 99.5127
R12250 VDD.n1517 VDD.n480 99.5127
R12251 VDD.n1577 VDD.n480 99.5127
R12252 VDD.n1577 VDD.n478 99.5127
R12253 VDD.n1581 VDD.n478 99.5127
R12254 VDD.n1581 VDD.n466 99.5127
R12255 VDD.n1946 VDD.n1945 99.5127
R12256 VDD.n1943 VDD.n1926 99.5127
R12257 VDD.n1939 VDD.n1938 99.5127
R12258 VDD.n1936 VDD.n1929 99.5127
R12259 VDD.n1932 VDD.n1931 99.5127
R12260 VDD.n2034 VDD.n2033 99.5127
R12261 VDD.n2031 VDD.n310 99.5127
R12262 VDD.n2027 VDD.n2026 99.5127
R12263 VDD.n2024 VDD.n313 99.5127
R12264 VDD.n2020 VDD.n2019 99.5127
R12265 VDD.n1731 VDD.n1630 99.5127
R12266 VDD.n1630 VDD.n440 99.5127
R12267 VDD.n1726 VDD.n440 99.5127
R12268 VDD.n1726 VDD.n433 99.5127
R12269 VDD.n1723 VDD.n433 99.5127
R12270 VDD.n1723 VDD.n427 99.5127
R12271 VDD.n1720 VDD.n427 99.5127
R12272 VDD.n1720 VDD.n422 99.5127
R12273 VDD.n1717 VDD.n422 99.5127
R12274 VDD.n1717 VDD.n415 99.5127
R12275 VDD.n1714 VDD.n415 99.5127
R12276 VDD.n1714 VDD.n409 99.5127
R12277 VDD.n1711 VDD.n409 99.5127
R12278 VDD.n1711 VDD.n404 99.5127
R12279 VDD.n1708 VDD.n404 99.5127
R12280 VDD.n1708 VDD.n397 99.5127
R12281 VDD.n1705 VDD.n397 99.5127
R12282 VDD.n1705 VDD.n391 99.5127
R12283 VDD.n1702 VDD.n391 99.5127
R12284 VDD.n1702 VDD.n386 99.5127
R12285 VDD.n1699 VDD.n386 99.5127
R12286 VDD.n1699 VDD.n380 99.5127
R12287 VDD.n1696 VDD.n380 99.5127
R12288 VDD.n1696 VDD.n374 99.5127
R12289 VDD.n1693 VDD.n374 99.5127
R12290 VDD.n1693 VDD.n368 99.5127
R12291 VDD.n1690 VDD.n368 99.5127
R12292 VDD.n1690 VDD.n361 99.5127
R12293 VDD.n1687 VDD.n361 99.5127
R12294 VDD.n1687 VDD.n354 99.5127
R12295 VDD.n1684 VDD.n354 99.5127
R12296 VDD.n1684 VDD.n348 99.5127
R12297 VDD.n348 VDD.n321 99.5127
R12298 VDD.n2013 VDD.n321 99.5127
R12299 VDD.n2013 VDD.n319 99.5127
R12300 VDD.n1646 VDD.n1643 99.5127
R12301 VDD.n1650 VDD.n1648 99.5127
R12302 VDD.n1654 VDD.n1640 99.5127
R12303 VDD.n1658 VDD.n1656 99.5127
R12304 VDD.n1662 VDD.n1638 99.5127
R12305 VDD.n1666 VDD.n1664 99.5127
R12306 VDD.n1670 VDD.n1636 99.5127
R12307 VDD.n1674 VDD.n1672 99.5127
R12308 VDD.n1678 VDD.n1634 99.5127
R12309 VDD.n1680 VDD.n1629 99.5127
R12310 VDD.n1837 VDD.n441 99.5127
R12311 VDD.n1841 VDD.n441 99.5127
R12312 VDD.n1841 VDD.n430 99.5127
R12313 VDD.n1849 VDD.n430 99.5127
R12314 VDD.n1849 VDD.n428 99.5127
R12315 VDD.n1853 VDD.n428 99.5127
R12316 VDD.n1853 VDD.n419 99.5127
R12317 VDD.n1861 VDD.n419 99.5127
R12318 VDD.n1861 VDD.n417 99.5127
R12319 VDD.n1865 VDD.n417 99.5127
R12320 VDD.n1865 VDD.n407 99.5127
R12321 VDD.n1873 VDD.n407 99.5127
R12322 VDD.n1873 VDD.n405 99.5127
R12323 VDD.n1877 VDD.n405 99.5127
R12324 VDD.n1877 VDD.n394 99.5127
R12325 VDD.n1885 VDD.n394 99.5127
R12326 VDD.n1885 VDD.n392 99.5127
R12327 VDD.n1889 VDD.n392 99.5127
R12328 VDD.n1889 VDD.n383 99.5127
R12329 VDD.n1897 VDD.n383 99.5127
R12330 VDD.n1897 VDD.n381 99.5127
R12331 VDD.n1901 VDD.n381 99.5127
R12332 VDD.n1901 VDD.n371 99.5127
R12333 VDD.n1909 VDD.n371 99.5127
R12334 VDD.n1909 VDD.n369 99.5127
R12335 VDD.n1913 VDD.n369 99.5127
R12336 VDD.n1913 VDD.n358 99.5127
R12337 VDD.n1921 VDD.n358 99.5127
R12338 VDD.n1921 VDD.n355 99.5127
R12339 VDD.n1955 VDD.n355 99.5127
R12340 VDD.n1955 VDD.n356 99.5127
R12341 VDD.n356 VDD.n349 99.5127
R12342 VDD.n1950 VDD.n349 99.5127
R12343 VDD.n1950 VDD.n325 99.5127
R12344 VDD.n1947 VDD.n325 99.5127
R12345 VDD.n1566 VDD.n1565 99.5127
R12346 VDD.n1562 VDD.n1561 99.5127
R12347 VDD.n1558 VDD.n1557 99.5127
R12348 VDD.n1554 VDD.n1553 99.5127
R12349 VDD.n1550 VDD.n1549 99.5127
R12350 VDD.n1546 VDD.n1545 99.5127
R12351 VDD.n1542 VDD.n1541 99.5127
R12352 VDD.n1538 VDD.n1537 99.5127
R12353 VDD.n1534 VDD.n1533 99.5127
R12354 VDD.n1529 VDD.n455 99.5127
R12355 VDD.n1380 VDD.n584 99.5127
R12356 VDD.n1380 VDD.n578 99.5127
R12357 VDD.n1377 VDD.n578 99.5127
R12358 VDD.n1377 VDD.n571 99.5127
R12359 VDD.n1374 VDD.n571 99.5127
R12360 VDD.n1374 VDD.n565 99.5127
R12361 VDD.n1371 VDD.n565 99.5127
R12362 VDD.n1371 VDD.n560 99.5127
R12363 VDD.n1368 VDD.n560 99.5127
R12364 VDD.n1368 VDD.n554 99.5127
R12365 VDD.n1365 VDD.n554 99.5127
R12366 VDD.n1365 VDD.n548 99.5127
R12367 VDD.n1362 VDD.n548 99.5127
R12368 VDD.n1362 VDD.n542 99.5127
R12369 VDD.n1359 VDD.n542 99.5127
R12370 VDD.n1359 VDD.n535 99.5127
R12371 VDD.n1356 VDD.n535 99.5127
R12372 VDD.n1356 VDD.n529 99.5127
R12373 VDD.n1353 VDD.n529 99.5127
R12374 VDD.n1353 VDD.n524 99.5127
R12375 VDD.n1350 VDD.n524 99.5127
R12376 VDD.n1350 VDD.n517 99.5127
R12377 VDD.n1347 VDD.n517 99.5127
R12378 VDD.n1347 VDD.n511 99.5127
R12379 VDD.n1344 VDD.n511 99.5127
R12380 VDD.n1344 VDD.n506 99.5127
R12381 VDD.n1341 VDD.n506 99.5127
R12382 VDD.n1341 VDD.n498 99.5127
R12383 VDD.n498 VDD.n490 99.5127
R12384 VDD.n1519 VDD.n490 99.5127
R12385 VDD.n1520 VDD.n1519 99.5127
R12386 VDD.n1520 VDD.n483 99.5127
R12387 VDD.n1523 VDD.n483 99.5127
R12388 VDD.n1523 VDD.n476 99.5127
R12389 VDD.n1526 VDD.n476 99.5127
R12390 VDD.n1421 VDD.n1419 99.5127
R12391 VDD.n1417 VDD.n587 99.5127
R12392 VDD.n1413 VDD.n1411 99.5127
R12393 VDD.n1409 VDD.n589 99.5127
R12394 VDD.n1405 VDD.n1403 99.5127
R12395 VDD.n1401 VDD.n1331 99.5127
R12396 VDD.n1397 VDD.n1395 99.5127
R12397 VDD.n1393 VDD.n1333 99.5127
R12398 VDD.n1389 VDD.n1387 99.5127
R12399 VDD.n1385 VDD.n1335 99.5127
R12400 VDD.n1425 VDD.n575 99.5127
R12401 VDD.n1433 VDD.n575 99.5127
R12402 VDD.n1433 VDD.n573 99.5127
R12403 VDD.n1437 VDD.n573 99.5127
R12404 VDD.n1437 VDD.n563 99.5127
R12405 VDD.n1445 VDD.n563 99.5127
R12406 VDD.n1445 VDD.n561 99.5127
R12407 VDD.n1449 VDD.n561 99.5127
R12408 VDD.n1449 VDD.n551 99.5127
R12409 VDD.n1457 VDD.n551 99.5127
R12410 VDD.n1457 VDD.n549 99.5127
R12411 VDD.n1461 VDD.n549 99.5127
R12412 VDD.n1461 VDD.n539 99.5127
R12413 VDD.n1469 VDD.n539 99.5127
R12414 VDD.n1469 VDD.n537 99.5127
R12415 VDD.n1473 VDD.n537 99.5127
R12416 VDD.n1473 VDD.n527 99.5127
R12417 VDD.n1481 VDD.n527 99.5127
R12418 VDD.n1481 VDD.n525 99.5127
R12419 VDD.n1485 VDD.n525 99.5127
R12420 VDD.n1485 VDD.n514 99.5127
R12421 VDD.n1493 VDD.n514 99.5127
R12422 VDD.n1493 VDD.n512 99.5127
R12423 VDD.n1497 VDD.n512 99.5127
R12424 VDD.n1497 VDD.n503 99.5127
R12425 VDD.n1505 VDD.n503 99.5127
R12426 VDD.n1505 VDD.n500 99.5127
R12427 VDD.n1511 VDD.n500 99.5127
R12428 VDD.n1511 VDD.n501 99.5127
R12429 VDD.n501 VDD.n492 99.5127
R12430 VDD.n492 VDD.n484 99.5127
R12431 VDD.n1575 VDD.n484 99.5127
R12432 VDD.n1575 VDD.n485 99.5127
R12433 VDD.n485 VDD.n477 99.5127
R12434 VDD.n1570 VDD.n477 99.5127
R12435 VDD.n1642 VDD.n1627 72.8958
R12436 VDD.n1647 VDD.n1627 72.8958
R12437 VDD.n1649 VDD.n1627 72.8958
R12438 VDD.n1655 VDD.n1627 72.8958
R12439 VDD.n1657 VDD.n1627 72.8958
R12440 VDD.n1663 VDD.n1627 72.8958
R12441 VDD.n1665 VDD.n1627 72.8958
R12442 VDD.n1671 VDD.n1627 72.8958
R12443 VDD.n1673 VDD.n1627 72.8958
R12444 VDD.n1679 VDD.n1627 72.8958
R12445 VDD.n2018 VDD.n309 72.8958
R12446 VDD.n317 VDD.n309 72.8958
R12447 VDD.n2025 VDD.n309 72.8958
R12448 VDD.n312 VDD.n309 72.8958
R12449 VDD.n2032 VDD.n309 72.8958
R12450 VDD.n309 VDD.n308 72.8958
R12451 VDD.n1930 VDD.n309 72.8958
R12452 VDD.n1937 VDD.n309 72.8958
R12453 VDD.n1928 VDD.n309 72.8958
R12454 VDD.n1944 VDD.n309 72.8958
R12455 VDD.n1205 VDD.n582 72.8958
R12456 VDD.n1211 VDD.n582 72.8958
R12457 VDD.n1213 VDD.n582 72.8958
R12458 VDD.n1219 VDD.n582 72.8958
R12459 VDD.n1222 VDD.n582 72.8958
R12460 VDD.n1299 VDD.n582 72.8958
R12461 VDD.n1225 VDD.n582 72.8958
R12462 VDD.n1292 VDD.n582 72.8958
R12463 VDD.n1286 VDD.n582 72.8958
R12464 VDD.n1231 VDD.n582 72.8958
R12465 VDD.n1626 VDD.n456 72.8958
R12466 VDD.n1626 VDD.n457 72.8958
R12467 VDD.n1626 VDD.n458 72.8958
R12468 VDD.n1626 VDD.n459 72.8958
R12469 VDD.n1626 VDD.n460 72.8958
R12470 VDD.n1626 VDD.n461 72.8958
R12471 VDD.n1626 VDD.n462 72.8958
R12472 VDD.n1626 VDD.n463 72.8958
R12473 VDD.n1626 VDD.n464 72.8958
R12474 VDD.n1626 VDD.n465 72.8958
R12475 VDD.n1830 VDD.n1627 72.8958
R12476 VDD.n1734 VDD.n1627 72.8958
R12477 VDD.n1823 VDD.n1627 72.8958
R12478 VDD.n1817 VDD.n1627 72.8958
R12479 VDD.n1815 VDD.n1627 72.8958
R12480 VDD.n1809 VDD.n1627 72.8958
R12481 VDD.n1807 VDD.n1627 72.8958
R12482 VDD.n1801 VDD.n1627 72.8958
R12483 VDD.n1799 VDD.n1627 72.8958
R12484 VDD.n1792 VDD.n1627 72.8958
R12485 VDD.n1968 VDD.n309 72.8958
R12486 VDD.n1976 VDD.n309 72.8958
R12487 VDD.n341 VDD.n309 72.8958
R12488 VDD.n1983 VDD.n309 72.8958
R12489 VDD.n338 VDD.n309 72.8958
R12490 VDD.n1991 VDD.n309 72.8958
R12491 VDD.n335 VDD.n309 72.8958
R12492 VDD.n1998 VDD.n309 72.8958
R12493 VDD.n332 VDD.n309 72.8958
R12494 VDD.n2005 VDD.n309 72.8958
R12495 VDD.n1626 VDD.n454 72.8958
R12496 VDD.n1626 VDD.n453 72.8958
R12497 VDD.n1626 VDD.n452 72.8958
R12498 VDD.n1626 VDD.n451 72.8958
R12499 VDD.n1626 VDD.n450 72.8958
R12500 VDD.n1626 VDD.n449 72.8958
R12501 VDD.n1626 VDD.n448 72.8958
R12502 VDD.n1626 VDD.n447 72.8958
R12503 VDD.n1626 VDD.n446 72.8958
R12504 VDD.n1626 VDD.n445 72.8958
R12505 VDD.n1420 VDD.n582 72.8958
R12506 VDD.n1418 VDD.n582 72.8958
R12507 VDD.n1412 VDD.n582 72.8958
R12508 VDD.n1410 VDD.n582 72.8958
R12509 VDD.n1404 VDD.n582 72.8958
R12510 VDD.n1402 VDD.n582 72.8958
R12511 VDD.n1396 VDD.n582 72.8958
R12512 VDD.n1394 VDD.n582 72.8958
R12513 VDD.n1388 VDD.n582 72.8958
R12514 VDD.n1386 VDD.n582 72.8958
R12515 VDD.t162 VDD.n582 69.3153
R12516 VDD.n309 VDD.t144 69.3153
R12517 VDD.n910 VDD.n909 66.2847
R12518 VDD.n909 VDD.n741 66.2847
R12519 VDD.n909 VDD.n742 66.2847
R12520 VDD.n909 VDD.n743 66.2847
R12521 VDD.n909 VDD.n744 66.2847
R12522 VDD.n909 VDD.n745 66.2847
R12523 VDD.n909 VDD.n746 66.2847
R12524 VDD.n909 VDD.n747 66.2847
R12525 VDD.n909 VDD.n748 66.2847
R12526 VDD.n909 VDD.n749 66.2847
R12527 VDD.n909 VDD.n750 66.2847
R12528 VDD.n909 VDD.n751 66.2847
R12529 VDD.n909 VDD.n752 66.2847
R12530 VDD.n909 VDD.n753 66.2847
R12531 VDD.n909 VDD.n754 66.2847
R12532 VDD.n909 VDD.n755 66.2847
R12533 VDD.n909 VDD.n756 66.2847
R12534 VDD.n909 VDD.n757 66.2847
R12535 VDD.n909 VDD.n758 66.2847
R12536 VDD.n909 VDD.n759 66.2847
R12537 VDD.n909 VDD.n760 66.2847
R12538 VDD.n909 VDD.n761 66.2847
R12539 VDD.n909 VDD.n762 66.2847
R12540 VDD.n1323 VDD.n602 66.2847
R12541 VDD.n602 VDD.n601 66.2847
R12542 VDD.n1125 VDD.n602 66.2847
R12543 VDD.n1130 VDD.n602 66.2847
R12544 VDD.n1123 VDD.n602 66.2847
R12545 VDD.n1137 VDD.n602 66.2847
R12546 VDD.n1117 VDD.n602 66.2847
R12547 VDD.n1147 VDD.n602 66.2847
R12548 VDD.n1110 VDD.n602 66.2847
R12549 VDD.n1154 VDD.n602 66.2847
R12550 VDD.n1103 VDD.n602 66.2847
R12551 VDD.n1161 VDD.n602 66.2847
R12552 VDD.n1096 VDD.n602 66.2847
R12553 VDD.n1171 VDD.n602 66.2847
R12554 VDD.n1089 VDD.n602 66.2847
R12555 VDD.n1178 VDD.n602 66.2847
R12556 VDD.n1082 VDD.n602 66.2847
R12557 VDD.n1185 VDD.n602 66.2847
R12558 VDD.n1075 VDD.n602 66.2847
R12559 VDD.n1195 VDD.n602 66.2847
R12560 VDD.n1070 VDD.n602 66.2847
R12561 VDD.n1309 VDD.n602 66.2847
R12562 VDD.n1312 VDD.n602 66.2847
R12563 VDD.n2142 VDD.n2141 66.2847
R12564 VDD.n2141 VDD.n246 66.2847
R12565 VDD.n2141 VDD.n247 66.2847
R12566 VDD.n2141 VDD.n248 66.2847
R12567 VDD.n2141 VDD.n249 66.2847
R12568 VDD.n2141 VDD.n250 66.2847
R12569 VDD.n2141 VDD.n251 66.2847
R12570 VDD.n2141 VDD.n252 66.2847
R12571 VDD.n2141 VDD.n253 66.2847
R12572 VDD.n2141 VDD.n254 66.2847
R12573 VDD.n2141 VDD.n255 66.2847
R12574 VDD.n2141 VDD.n256 66.2847
R12575 VDD.n2141 VDD.n257 66.2847
R12576 VDD.n2141 VDD.n258 66.2847
R12577 VDD.n2141 VDD.n259 66.2847
R12578 VDD.n2141 VDD.n260 66.2847
R12579 VDD.n2141 VDD.n261 66.2847
R12580 VDD.n2141 VDD.n262 66.2847
R12581 VDD.n2141 VDD.n263 66.2847
R12582 VDD.n2141 VDD.n264 66.2847
R12583 VDD.n2141 VDD.n265 66.2847
R12584 VDD.n2141 VDD.n266 66.2847
R12585 VDD.n2141 VDD.n267 66.2847
R12586 VDD.n168 VDD.n87 66.2847
R12587 VDD.n2253 VDD.n87 66.2847
R12588 VDD.n164 VDD.n87 66.2847
R12589 VDD.n2260 VDD.n87 66.2847
R12590 VDD.n157 VDD.n87 66.2847
R12591 VDD.n2267 VDD.n87 66.2847
R12592 VDD.n150 VDD.n87 66.2847
R12593 VDD.n2277 VDD.n87 66.2847
R12594 VDD.n143 VDD.n87 66.2847
R12595 VDD.n2284 VDD.n87 66.2847
R12596 VDD.n136 VDD.n87 66.2847
R12597 VDD.n2291 VDD.n87 66.2847
R12598 VDD.n129 VDD.n87 66.2847
R12599 VDD.n2301 VDD.n87 66.2847
R12600 VDD.n122 VDD.n87 66.2847
R12601 VDD.n2308 VDD.n87 66.2847
R12602 VDD.n115 VDD.n87 66.2847
R12603 VDD.n2315 VDD.n87 66.2847
R12604 VDD.n108 VDD.n87 66.2847
R12605 VDD.n2325 VDD.n87 66.2847
R12606 VDD.n101 VDD.n87 66.2847
R12607 VDD.n2332 VDD.n87 66.2847
R12608 VDD.n94 VDD.n87 66.2847
R12609 VDD.n1337 VDD.n1336 58.9581
R12610 VDD.n488 VDD.n487 58.9581
R12611 VDD.n1229 VDD.n1228 58.9581
R12612 VDD.n470 VDD.n469 58.9581
R12613 VDD.n1632 VDD.n1631 58.9581
R12614 VDD.n344 VDD.n343 58.9581
R12615 VDD.n1744 VDD.n1743 58.9581
R12616 VDD.n315 VDD.n314 58.9581
R12617 VDD.n2334 VDD.n94 52.4337
R12618 VDD.n2332 VDD.n2331 52.4337
R12619 VDD.n2327 VDD.n101 52.4337
R12620 VDD.n2325 VDD.n2324 52.4337
R12621 VDD.n2317 VDD.n108 52.4337
R12622 VDD.n2315 VDD.n2314 52.4337
R12623 VDD.n2310 VDD.n115 52.4337
R12624 VDD.n2308 VDD.n2307 52.4337
R12625 VDD.n2303 VDD.n122 52.4337
R12626 VDD.n2301 VDD.n2300 52.4337
R12627 VDD.n2293 VDD.n129 52.4337
R12628 VDD.n2291 VDD.n2290 52.4337
R12629 VDD.n2286 VDD.n136 52.4337
R12630 VDD.n2284 VDD.n2283 52.4337
R12631 VDD.n2279 VDD.n143 52.4337
R12632 VDD.n2277 VDD.n2276 52.4337
R12633 VDD.n2269 VDD.n150 52.4337
R12634 VDD.n2267 VDD.n2266 52.4337
R12635 VDD.n2262 VDD.n157 52.4337
R12636 VDD.n2260 VDD.n2259 52.4337
R12637 VDD.n2255 VDD.n164 52.4337
R12638 VDD.n2253 VDD.n2252 52.4337
R12639 VDD.n169 VDD.n168 52.4337
R12640 VDD.n2143 VDD.n2142 52.4337
R12641 VDD.n268 VDD.n246 52.4337
R12642 VDD.n2135 VDD.n247 52.4337
R12643 VDD.n2131 VDD.n248 52.4337
R12644 VDD.n2127 VDD.n249 52.4337
R12645 VDD.n2120 VDD.n250 52.4337
R12646 VDD.n2116 VDD.n251 52.4337
R12647 VDD.n2112 VDD.n252 52.4337
R12648 VDD.n2108 VDD.n253 52.4337
R12649 VDD.n2104 VDD.n254 52.4337
R12650 VDD.n2100 VDD.n255 52.4337
R12651 VDD.n2093 VDD.n256 52.4337
R12652 VDD.n2089 VDD.n257 52.4337
R12653 VDD.n2085 VDD.n258 52.4337
R12654 VDD.n2081 VDD.n259 52.4337
R12655 VDD.n2077 VDD.n260 52.4337
R12656 VDD.n2073 VDD.n261 52.4337
R12657 VDD.n2066 VDD.n262 52.4337
R12658 VDD.n2062 VDD.n263 52.4337
R12659 VDD.n2058 VDD.n264 52.4337
R12660 VDD.n2037 VDD.n265 52.4337
R12661 VDD.n2051 VDD.n266 52.4337
R12662 VDD.n2048 VDD.n267 52.4337
R12663 VDD.n1312 VDD.n1311 52.4337
R12664 VDD.n1309 VDD.n1308 52.4337
R12665 VDD.n1197 VDD.n1070 52.4337
R12666 VDD.n1195 VDD.n1194 52.4337
R12667 VDD.n1187 VDD.n1075 52.4337
R12668 VDD.n1185 VDD.n1184 52.4337
R12669 VDD.n1180 VDD.n1082 52.4337
R12670 VDD.n1178 VDD.n1177 52.4337
R12671 VDD.n1173 VDD.n1089 52.4337
R12672 VDD.n1171 VDD.n1170 52.4337
R12673 VDD.n1163 VDD.n1096 52.4337
R12674 VDD.n1161 VDD.n1160 52.4337
R12675 VDD.n1156 VDD.n1103 52.4337
R12676 VDD.n1154 VDD.n1153 52.4337
R12677 VDD.n1149 VDD.n1110 52.4337
R12678 VDD.n1147 VDD.n1146 52.4337
R12679 VDD.n1139 VDD.n1117 52.4337
R12680 VDD.n1137 VDD.n1136 52.4337
R12681 VDD.n1132 VDD.n1123 52.4337
R12682 VDD.n1130 VDD.n1129 52.4337
R12683 VDD.n1125 VDD.n1124 52.4337
R12684 VDD.n601 VDD.n596 52.4337
R12685 VDD.n1323 VDD.n1322 52.4337
R12686 VDD.n911 VDD.n910 52.4337
R12687 VDD.n763 VDD.n741 52.4337
R12688 VDD.n767 VDD.n742 52.4337
R12689 VDD.n769 VDD.n743 52.4337
R12690 VDD.n773 VDD.n744 52.4337
R12691 VDD.n775 VDD.n745 52.4337
R12692 VDD.n779 VDD.n746 52.4337
R12693 VDD.n781 VDD.n747 52.4337
R12694 VDD.n785 VDD.n748 52.4337
R12695 VDD.n787 VDD.n749 52.4337
R12696 VDD.n791 VDD.n750 52.4337
R12697 VDD.n793 VDD.n751 52.4337
R12698 VDD.n797 VDD.n752 52.4337
R12699 VDD.n799 VDD.n753 52.4337
R12700 VDD.n803 VDD.n754 52.4337
R12701 VDD.n805 VDD.n755 52.4337
R12702 VDD.n809 VDD.n756 52.4337
R12703 VDD.n811 VDD.n757 52.4337
R12704 VDD.n815 VDD.n758 52.4337
R12705 VDD.n817 VDD.n759 52.4337
R12706 VDD.n821 VDD.n760 52.4337
R12707 VDD.n823 VDD.n761 52.4337
R12708 VDD.n830 VDD.n762 52.4337
R12709 VDD.n910 VDD.n740 52.4337
R12710 VDD.n766 VDD.n741 52.4337
R12711 VDD.n768 VDD.n742 52.4337
R12712 VDD.n772 VDD.n743 52.4337
R12713 VDD.n774 VDD.n744 52.4337
R12714 VDD.n778 VDD.n745 52.4337
R12715 VDD.n780 VDD.n746 52.4337
R12716 VDD.n784 VDD.n747 52.4337
R12717 VDD.n786 VDD.n748 52.4337
R12718 VDD.n790 VDD.n749 52.4337
R12719 VDD.n792 VDD.n750 52.4337
R12720 VDD.n796 VDD.n751 52.4337
R12721 VDD.n798 VDD.n752 52.4337
R12722 VDD.n802 VDD.n753 52.4337
R12723 VDD.n804 VDD.n754 52.4337
R12724 VDD.n808 VDD.n755 52.4337
R12725 VDD.n810 VDD.n756 52.4337
R12726 VDD.n814 VDD.n757 52.4337
R12727 VDD.n816 VDD.n758 52.4337
R12728 VDD.n820 VDD.n759 52.4337
R12729 VDD.n822 VDD.n760 52.4337
R12730 VDD.n826 VDD.n761 52.4337
R12731 VDD.n827 VDD.n762 52.4337
R12732 VDD.n1324 VDD.n1323 52.4337
R12733 VDD.n601 VDD.n595 52.4337
R12734 VDD.n1126 VDD.n1125 52.4337
R12735 VDD.n1131 VDD.n1130 52.4337
R12736 VDD.n1123 VDD.n1118 52.4337
R12737 VDD.n1138 VDD.n1137 52.4337
R12738 VDD.n1117 VDD.n1111 52.4337
R12739 VDD.n1148 VDD.n1147 52.4337
R12740 VDD.n1110 VDD.n1104 52.4337
R12741 VDD.n1155 VDD.n1154 52.4337
R12742 VDD.n1103 VDD.n1097 52.4337
R12743 VDD.n1162 VDD.n1161 52.4337
R12744 VDD.n1096 VDD.n1090 52.4337
R12745 VDD.n1172 VDD.n1171 52.4337
R12746 VDD.n1089 VDD.n1083 52.4337
R12747 VDD.n1179 VDD.n1178 52.4337
R12748 VDD.n1082 VDD.n1076 52.4337
R12749 VDD.n1186 VDD.n1185 52.4337
R12750 VDD.n1075 VDD.n1071 52.4337
R12751 VDD.n1196 VDD.n1195 52.4337
R12752 VDD.n1070 VDD.n1066 52.4337
R12753 VDD.n1310 VDD.n1309 52.4337
R12754 VDD.n1313 VDD.n1312 52.4337
R12755 VDD.n2142 VDD.n245 52.4337
R12756 VDD.n2136 VDD.n246 52.4337
R12757 VDD.n2132 VDD.n247 52.4337
R12758 VDD.n2128 VDD.n248 52.4337
R12759 VDD.n2121 VDD.n249 52.4337
R12760 VDD.n2117 VDD.n250 52.4337
R12761 VDD.n2113 VDD.n251 52.4337
R12762 VDD.n2109 VDD.n252 52.4337
R12763 VDD.n2105 VDD.n253 52.4337
R12764 VDD.n2101 VDD.n254 52.4337
R12765 VDD.n2094 VDD.n255 52.4337
R12766 VDD.n2090 VDD.n256 52.4337
R12767 VDD.n2086 VDD.n257 52.4337
R12768 VDD.n2082 VDD.n258 52.4337
R12769 VDD.n2078 VDD.n259 52.4337
R12770 VDD.n2074 VDD.n260 52.4337
R12771 VDD.n2067 VDD.n261 52.4337
R12772 VDD.n2063 VDD.n262 52.4337
R12773 VDD.n2059 VDD.n263 52.4337
R12774 VDD.n2036 VDD.n264 52.4337
R12775 VDD.n2039 VDD.n265 52.4337
R12776 VDD.n2049 VDD.n266 52.4337
R12777 VDD.n2041 VDD.n267 52.4337
R12778 VDD.n168 VDD.n165 52.4337
R12779 VDD.n2254 VDD.n2253 52.4337
R12780 VDD.n164 VDD.n158 52.4337
R12781 VDD.n2261 VDD.n2260 52.4337
R12782 VDD.n157 VDD.n151 52.4337
R12783 VDD.n2268 VDD.n2267 52.4337
R12784 VDD.n150 VDD.n144 52.4337
R12785 VDD.n2278 VDD.n2277 52.4337
R12786 VDD.n143 VDD.n137 52.4337
R12787 VDD.n2285 VDD.n2284 52.4337
R12788 VDD.n136 VDD.n130 52.4337
R12789 VDD.n2292 VDD.n2291 52.4337
R12790 VDD.n129 VDD.n123 52.4337
R12791 VDD.n2302 VDD.n2301 52.4337
R12792 VDD.n122 VDD.n116 52.4337
R12793 VDD.n2309 VDD.n2308 52.4337
R12794 VDD.n115 VDD.n109 52.4337
R12795 VDD.n2316 VDD.n2315 52.4337
R12796 VDD.n108 VDD.n102 52.4337
R12797 VDD.n2326 VDD.n2325 52.4337
R12798 VDD.n101 VDD.n95 52.4337
R12799 VDD.n2333 VDD.n2332 52.4337
R12800 VDD.n94 VDD.n91 52.4337
R12801 VDD.n832 VDD.n831 45.3823
R12802 VDD.n852 VDD.n851 45.3823
R12803 VDD.n873 VDD.n872 45.3823
R12804 VDD.n894 VDD.n893 45.3823
R12805 VDD.n599 VDD.n598 45.3823
R12806 VDD.n1142 VDD.n1141 45.3823
R12807 VDD.n1166 VDD.n1165 45.3823
R12808 VDD.n1190 VDD.n1189 45.3823
R12809 VDD.n172 VDD.n171 45.3823
R12810 VDD.n2272 VDD.n2271 45.3823
R12811 VDD.n2296 VDD.n2295 45.3823
R12812 VDD.n2320 VDD.n2319 45.3823
R12813 VDD.n2070 VDD.n2069 45.3823
R12814 VDD.n2097 VDD.n2096 45.3823
R12815 VDD.n2124 VDD.n2123 45.3823
R12816 VDD.n2046 VDD.n2045 45.3823
R12817 VDD.n2005 VDD.n2004 39.2114
R12818 VDD.n2000 VDD.n332 39.2114
R12819 VDD.n1998 VDD.n1997 39.2114
R12820 VDD.n1993 VDD.n335 39.2114
R12821 VDD.n1991 VDD.n1990 39.2114
R12822 VDD.n1985 VDD.n338 39.2114
R12823 VDD.n1983 VDD.n1982 39.2114
R12824 VDD.n1978 VDD.n341 39.2114
R12825 VDD.n1976 VDD.n1975 39.2114
R12826 VDD.n1970 VDD.n1968 39.2114
R12827 VDD.n1830 VDD.n1732 39.2114
R12828 VDD.n1828 VDD.n1734 39.2114
R12829 VDD.n1824 VDD.n1823 39.2114
R12830 VDD.n1817 VDD.n1736 39.2114
R12831 VDD.n1816 VDD.n1815 39.2114
R12832 VDD.n1809 VDD.n1738 39.2114
R12833 VDD.n1808 VDD.n1807 39.2114
R12834 VDD.n1801 VDD.n1740 39.2114
R12835 VDD.n1800 VDD.n1799 39.2114
R12836 VDD.n1792 VDD.n1742 39.2114
R12837 VDD.n1621 VDD.n465 39.2114
R12838 VDD.n1617 VDD.n464 39.2114
R12839 VDD.n1613 VDD.n463 39.2114
R12840 VDD.n1609 VDD.n462 39.2114
R12841 VDD.n1605 VDD.n461 39.2114
R12842 VDD.n1601 VDD.n460 39.2114
R12843 VDD.n1597 VDD.n459 39.2114
R12844 VDD.n1593 VDD.n458 39.2114
R12845 VDD.n1589 VDD.n457 39.2114
R12846 VDD.n1585 VDD.n456 39.2114
R12847 VDD.n1205 VDD.n581 39.2114
R12848 VDD.n1211 VDD.n1210 39.2114
R12849 VDD.n1214 VDD.n1213 39.2114
R12850 VDD.n1219 VDD.n1218 39.2114
R12851 VDD.n1222 VDD.n1221 39.2114
R12852 VDD.n1300 VDD.n1299 39.2114
R12853 VDD.n1297 VDD.n1225 39.2114
R12854 VDD.n1293 VDD.n1292 39.2114
R12855 VDD.n1286 VDD.n1227 39.2114
R12856 VDD.n1285 VDD.n1231 39.2114
R12857 VDD.n1944 VDD.n1943 39.2114
R12858 VDD.n1939 VDD.n1928 39.2114
R12859 VDD.n1937 VDD.n1936 39.2114
R12860 VDD.n1932 VDD.n1930 39.2114
R12861 VDD.n2034 VDD.n308 39.2114
R12862 VDD.n2032 VDD.n2031 39.2114
R12863 VDD.n2027 VDD.n312 39.2114
R12864 VDD.n2025 VDD.n2024 39.2114
R12865 VDD.n2020 VDD.n317 39.2114
R12866 VDD.n2018 VDD.n2017 39.2114
R12867 VDD.n1642 VDD.n443 39.2114
R12868 VDD.n1647 VDD.n1646 39.2114
R12869 VDD.n1650 VDD.n1649 39.2114
R12870 VDD.n1655 VDD.n1654 39.2114
R12871 VDD.n1658 VDD.n1657 39.2114
R12872 VDD.n1663 VDD.n1662 39.2114
R12873 VDD.n1666 VDD.n1665 39.2114
R12874 VDD.n1671 VDD.n1670 39.2114
R12875 VDD.n1674 VDD.n1673 39.2114
R12876 VDD.n1679 VDD.n1678 39.2114
R12877 VDD.n1643 VDD.n1642 39.2114
R12878 VDD.n1648 VDD.n1647 39.2114
R12879 VDD.n1649 VDD.n1640 39.2114
R12880 VDD.n1656 VDD.n1655 39.2114
R12881 VDD.n1657 VDD.n1638 39.2114
R12882 VDD.n1664 VDD.n1663 39.2114
R12883 VDD.n1665 VDD.n1636 39.2114
R12884 VDD.n1672 VDD.n1671 39.2114
R12885 VDD.n1673 VDD.n1634 39.2114
R12886 VDD.n1680 VDD.n1679 39.2114
R12887 VDD.n2019 VDD.n2018 39.2114
R12888 VDD.n317 VDD.n313 39.2114
R12889 VDD.n2026 VDD.n2025 39.2114
R12890 VDD.n312 VDD.n310 39.2114
R12891 VDD.n2033 VDD.n2032 39.2114
R12892 VDD.n1931 VDD.n308 39.2114
R12893 VDD.n1930 VDD.n1929 39.2114
R12894 VDD.n1938 VDD.n1937 39.2114
R12895 VDD.n1928 VDD.n1926 39.2114
R12896 VDD.n1945 VDD.n1944 39.2114
R12897 VDD.n1206 VDD.n1205 39.2114
R12898 VDD.n1212 VDD.n1211 39.2114
R12899 VDD.n1213 VDD.n1202 39.2114
R12900 VDD.n1220 VDD.n1219 39.2114
R12901 VDD.n1223 VDD.n1222 39.2114
R12902 VDD.n1299 VDD.n1298 39.2114
R12903 VDD.n1294 VDD.n1225 39.2114
R12904 VDD.n1292 VDD.n1291 39.2114
R12905 VDD.n1287 VDD.n1286 39.2114
R12906 VDD.n1282 VDD.n1231 39.2114
R12907 VDD.n1588 VDD.n456 39.2114
R12908 VDD.n1592 VDD.n457 39.2114
R12909 VDD.n1596 VDD.n458 39.2114
R12910 VDD.n1600 VDD.n459 39.2114
R12911 VDD.n1604 VDD.n460 39.2114
R12912 VDD.n1608 VDD.n461 39.2114
R12913 VDD.n1612 VDD.n462 39.2114
R12914 VDD.n1616 VDD.n463 39.2114
R12915 VDD.n1620 VDD.n464 39.2114
R12916 VDD.n467 VDD.n465 39.2114
R12917 VDD.n1831 VDD.n1830 39.2114
R12918 VDD.n1825 VDD.n1734 39.2114
R12919 VDD.n1823 VDD.n1822 39.2114
R12920 VDD.n1818 VDD.n1817 39.2114
R12921 VDD.n1815 VDD.n1814 39.2114
R12922 VDD.n1810 VDD.n1809 39.2114
R12923 VDD.n1807 VDD.n1806 39.2114
R12924 VDD.n1802 VDD.n1801 39.2114
R12925 VDD.n1799 VDD.n1798 39.2114
R12926 VDD.n1793 VDD.n1792 39.2114
R12927 VDD.n1968 VDD.n342 39.2114
R12928 VDD.n1977 VDD.n1976 39.2114
R12929 VDD.n341 VDD.n339 39.2114
R12930 VDD.n1984 VDD.n1983 39.2114
R12931 VDD.n338 VDD.n336 39.2114
R12932 VDD.n1992 VDD.n1991 39.2114
R12933 VDD.n335 VDD.n333 39.2114
R12934 VDD.n1999 VDD.n1998 39.2114
R12935 VDD.n332 VDD.n330 39.2114
R12936 VDD.n2006 VDD.n2005 39.2114
R12937 VDD.n1569 VDD.n445 39.2114
R12938 VDD.n1565 VDD.n446 39.2114
R12939 VDD.n1561 VDD.n447 39.2114
R12940 VDD.n1557 VDD.n448 39.2114
R12941 VDD.n1553 VDD.n449 39.2114
R12942 VDD.n1549 VDD.n450 39.2114
R12943 VDD.n1545 VDD.n451 39.2114
R12944 VDD.n1541 VDD.n452 39.2114
R12945 VDD.n1537 VDD.n453 39.2114
R12946 VDD.n1533 VDD.n454 39.2114
R12947 VDD.n1420 VDD.n585 39.2114
R12948 VDD.n1419 VDD.n1418 39.2114
R12949 VDD.n1412 VDD.n587 39.2114
R12950 VDD.n1411 VDD.n1410 39.2114
R12951 VDD.n1404 VDD.n589 39.2114
R12952 VDD.n1403 VDD.n1402 39.2114
R12953 VDD.n1396 VDD.n1331 39.2114
R12954 VDD.n1395 VDD.n1394 39.2114
R12955 VDD.n1388 VDD.n1333 39.2114
R12956 VDD.n1387 VDD.n1386 39.2114
R12957 VDD.n1529 VDD.n454 39.2114
R12958 VDD.n1534 VDD.n453 39.2114
R12959 VDD.n1538 VDD.n452 39.2114
R12960 VDD.n1542 VDD.n451 39.2114
R12961 VDD.n1546 VDD.n450 39.2114
R12962 VDD.n1550 VDD.n449 39.2114
R12963 VDD.n1554 VDD.n448 39.2114
R12964 VDD.n1558 VDD.n447 39.2114
R12965 VDD.n1562 VDD.n446 39.2114
R12966 VDD.n1566 VDD.n445 39.2114
R12967 VDD.n1421 VDD.n1420 39.2114
R12968 VDD.n1418 VDD.n1417 39.2114
R12969 VDD.n1413 VDD.n1412 39.2114
R12970 VDD.n1410 VDD.n1409 39.2114
R12971 VDD.n1405 VDD.n1404 39.2114
R12972 VDD.n1402 VDD.n1401 39.2114
R12973 VDD.n1397 VDD.n1396 39.2114
R12974 VDD.n1394 VDD.n1393 39.2114
R12975 VDD.n1389 VDD.n1388 39.2114
R12976 VDD.n1386 VDD.n1385 39.2114
R12977 VDD.n833 VDD.n832 37.2369
R12978 VDD.n853 VDD.n852 37.2369
R12979 VDD.n874 VDD.n873 37.2369
R12980 VDD.n895 VDD.n894 37.2369
R12981 VDD.n1325 VDD.n599 37.2369
R12982 VDD.n1143 VDD.n1142 37.2369
R12983 VDD.n1167 VDD.n1166 37.2369
R12984 VDD.n1191 VDD.n1190 37.2369
R12985 VDD.n2250 VDD.n172 37.2369
R12986 VDD.n2273 VDD.n2272 37.2369
R12987 VDD.n2297 VDD.n2296 37.2369
R12988 VDD.n2321 VDD.n2320 37.2369
R12989 VDD.n2071 VDD.n2070 37.2369
R12990 VDD.n2098 VDD.n2097 37.2369
R12991 VDD.n2125 VDD.n2124 37.2369
R12992 VDD.n2047 VDD.n2046 37.2369
R12993 VDD.n1428 VDD.n580 36.059
R12994 VDD.n1624 VDD.n468 36.059
R12995 VDD.n1586 VDD.n472 36.059
R12996 VDD.n1283 VDD.n1281 36.059
R12997 VDD.n1794 VDD.n1791 36.059
R12998 VDD.n1971 VDD.n1967 36.059
R12999 VDD.n1834 VDD.n1833 36.059
R13000 VDD.n2009 VDD.n2008 36.059
R13001 VDD.n1948 VDD.n1924 36.059
R13002 VDD.n2016 VDD.n2015 36.059
R13003 VDD.n1730 VDD.n1682 36.059
R13004 VDD.n1838 VDD.n442 36.059
R13005 VDD.n1424 VDD.n1423 36.059
R13006 VDD.n1571 VDD.n1568 36.059
R13007 VDD.n1528 VDD.n1527 36.059
R13008 VDD.n1383 VDD.n1382 36.059
R13009 VDD.n909 VDD.n734 34.8338
R13010 VDD.n1320 VDD.n602 34.8338
R13011 VDD.n2141 VDD.n239 34.8338
R13012 VDD.n2342 VDD.n87 34.8338
R13013 VDD.n1338 VDD.n1337 30.449
R13014 VDD.n1531 VDD.n488 30.449
R13015 VDD.n1230 VDD.n1229 30.449
R13016 VDD.n471 VDD.n470 30.449
R13017 VDD.n1633 VDD.n1632 30.449
R13018 VDD.n1973 VDD.n344 30.449
R13019 VDD.n1796 VDD.n1744 30.449
R13020 VDD.n316 VDD.n315 30.449
R13021 VDD.n1426 VDD.n582 24.2783
R13022 VDD.n1626 VDD.n444 24.2783
R13023 VDD.n1836 VDD.n1627 24.2783
R13024 VDD.n324 VDD.n309 24.2783
R13025 VDD.n920 VDD.n732 19.3944
R13026 VDD.n920 VDD.n730 19.3944
R13027 VDD.n924 VDD.n730 19.3944
R13028 VDD.n924 VDD.n721 19.3944
R13029 VDD.n936 VDD.n721 19.3944
R13030 VDD.n936 VDD.n719 19.3944
R13031 VDD.n940 VDD.n719 19.3944
R13032 VDD.n940 VDD.n709 19.3944
R13033 VDD.n952 VDD.n709 19.3944
R13034 VDD.n952 VDD.n707 19.3944
R13035 VDD.n956 VDD.n707 19.3944
R13036 VDD.n956 VDD.n697 19.3944
R13037 VDD.n968 VDD.n697 19.3944
R13038 VDD.n968 VDD.n695 19.3944
R13039 VDD.n972 VDD.n695 19.3944
R13040 VDD.n972 VDD.n684 19.3944
R13041 VDD.n985 VDD.n684 19.3944
R13042 VDD.n985 VDD.n682 19.3944
R13043 VDD.n989 VDD.n682 19.3944
R13044 VDD.n989 VDD.n653 19.3944
R13045 VDD.n1001 VDD.n653 19.3944
R13046 VDD.n1001 VDD.n651 19.3944
R13047 VDD.n1005 VDD.n651 19.3944
R13048 VDD.n1005 VDD.n641 19.3944
R13049 VDD.n1017 VDD.n641 19.3944
R13050 VDD.n1017 VDD.n639 19.3944
R13051 VDD.n1021 VDD.n639 19.3944
R13052 VDD.n1021 VDD.n629 19.3944
R13053 VDD.n1033 VDD.n629 19.3944
R13054 VDD.n1033 VDD.n627 19.3944
R13055 VDD.n1037 VDD.n627 19.3944
R13056 VDD.n1037 VDD.n616 19.3944
R13057 VDD.n1049 VDD.n616 19.3944
R13058 VDD.n1049 VDD.n613 19.3944
R13059 VDD.n1056 VDD.n613 19.3944
R13060 VDD.n1056 VDD.n614 19.3944
R13061 VDD.n614 VDD.n604 19.3944
R13062 VDD.n850 VDD.n812 19.3944
R13063 VDD.n846 VDD.n812 19.3944
R13064 VDD.n846 VDD.n845 19.3944
R13065 VDD.n845 VDD.n844 19.3944
R13066 VDD.n844 VDD.n818 19.3944
R13067 VDD.n840 VDD.n818 19.3944
R13068 VDD.n840 VDD.n839 19.3944
R13069 VDD.n839 VDD.n838 19.3944
R13070 VDD.n838 VDD.n824 19.3944
R13071 VDD.n834 VDD.n824 19.3944
R13072 VDD.n871 VDD.n794 19.3944
R13073 VDD.n867 VDD.n794 19.3944
R13074 VDD.n867 VDD.n866 19.3944
R13075 VDD.n866 VDD.n865 19.3944
R13076 VDD.n865 VDD.n800 19.3944
R13077 VDD.n861 VDD.n800 19.3944
R13078 VDD.n861 VDD.n860 19.3944
R13079 VDD.n860 VDD.n859 19.3944
R13080 VDD.n859 VDD.n806 19.3944
R13081 VDD.n855 VDD.n806 19.3944
R13082 VDD.n855 VDD.n854 19.3944
R13083 VDD.n892 VDD.n776 19.3944
R13084 VDD.n888 VDD.n776 19.3944
R13085 VDD.n888 VDD.n887 19.3944
R13086 VDD.n887 VDD.n886 19.3944
R13087 VDD.n886 VDD.n782 19.3944
R13088 VDD.n882 VDD.n782 19.3944
R13089 VDD.n882 VDD.n881 19.3944
R13090 VDD.n881 VDD.n880 19.3944
R13091 VDD.n880 VDD.n788 19.3944
R13092 VDD.n876 VDD.n788 19.3944
R13093 VDD.n876 VDD.n875 19.3944
R13094 VDD.n912 VDD.n739 19.3944
R13095 VDD.n907 VDD.n739 19.3944
R13096 VDD.n907 VDD.n764 19.3944
R13097 VDD.n903 VDD.n764 19.3944
R13098 VDD.n903 VDD.n902 19.3944
R13099 VDD.n902 VDD.n901 19.3944
R13100 VDD.n901 VDD.n770 19.3944
R13101 VDD.n897 VDD.n770 19.3944
R13102 VDD.n897 VDD.n896 19.3944
R13103 VDD.n1140 VDD.n1116 19.3944
R13104 VDD.n1135 VDD.n1116 19.3944
R13105 VDD.n1135 VDD.n1134 19.3944
R13106 VDD.n1134 VDD.n1133 19.3944
R13107 VDD.n1133 VDD.n1122 19.3944
R13108 VDD.n1128 VDD.n1127 19.3944
R13109 VDD.n1327 VDD.n594 19.3944
R13110 VDD.n1327 VDD.n1326 19.3944
R13111 VDD.n1164 VDD.n1095 19.3944
R13112 VDD.n1159 VDD.n1095 19.3944
R13113 VDD.n1159 VDD.n1158 19.3944
R13114 VDD.n1158 VDD.n1157 19.3944
R13115 VDD.n1157 VDD.n1102 19.3944
R13116 VDD.n1152 VDD.n1102 19.3944
R13117 VDD.n1152 VDD.n1151 19.3944
R13118 VDD.n1151 VDD.n1150 19.3944
R13119 VDD.n1150 VDD.n1109 19.3944
R13120 VDD.n1145 VDD.n1109 19.3944
R13121 VDD.n1145 VDD.n1144 19.3944
R13122 VDD.n1188 VDD.n1074 19.3944
R13123 VDD.n1183 VDD.n1074 19.3944
R13124 VDD.n1183 VDD.n1182 19.3944
R13125 VDD.n1182 VDD.n1181 19.3944
R13126 VDD.n1181 VDD.n1081 19.3944
R13127 VDD.n1176 VDD.n1081 19.3944
R13128 VDD.n1176 VDD.n1175 19.3944
R13129 VDD.n1175 VDD.n1174 19.3944
R13130 VDD.n1174 VDD.n1088 19.3944
R13131 VDD.n1169 VDD.n1088 19.3944
R13132 VDD.n1169 VDD.n1168 19.3944
R13133 VDD.n1315 VDD.n1314 19.3944
R13134 VDD.n1314 VDD.n1064 19.3944
R13135 VDD.n1065 VDD.n1064 19.3944
R13136 VDD.n1307 VDD.n1065 19.3944
R13137 VDD.n1198 VDD.n1067 19.3944
R13138 VDD.n1193 VDD.n1069 19.3944
R13139 VDD.n1193 VDD.n1192 19.3944
R13140 VDD.n916 VDD.n737 19.3944
R13141 VDD.n916 VDD.n727 19.3944
R13142 VDD.n928 VDD.n727 19.3944
R13143 VDD.n928 VDD.n725 19.3944
R13144 VDD.n932 VDD.n725 19.3944
R13145 VDD.n932 VDD.n715 19.3944
R13146 VDD.n944 VDD.n715 19.3944
R13147 VDD.n944 VDD.n713 19.3944
R13148 VDD.n948 VDD.n713 19.3944
R13149 VDD.n948 VDD.n703 19.3944
R13150 VDD.n960 VDD.n703 19.3944
R13151 VDD.n960 VDD.n701 19.3944
R13152 VDD.n964 VDD.n701 19.3944
R13153 VDD.n964 VDD.n691 19.3944
R13154 VDD.n976 VDD.n691 19.3944
R13155 VDD.n976 VDD.n689 19.3944
R13156 VDD.n981 VDD.n689 19.3944
R13157 VDD.n981 VDD.n679 19.3944
R13158 VDD.n993 VDD.n679 19.3944
R13159 VDD.n993 VDD.n657 19.3944
R13160 VDD.n997 VDD.n657 19.3944
R13161 VDD.n997 VDD.n647 19.3944
R13162 VDD.n1009 VDD.n647 19.3944
R13163 VDD.n1009 VDD.n645 19.3944
R13164 VDD.n1013 VDD.n645 19.3944
R13165 VDD.n1013 VDD.n635 19.3944
R13166 VDD.n1025 VDD.n635 19.3944
R13167 VDD.n1025 VDD.n633 19.3944
R13168 VDD.n1029 VDD.n633 19.3944
R13169 VDD.n1029 VDD.n623 19.3944
R13170 VDD.n1041 VDD.n623 19.3944
R13171 VDD.n1041 VDD.n621 19.3944
R13172 VDD.n1045 VDD.n621 19.3944
R13173 VDD.n1045 VDD.n610 19.3944
R13174 VDD.n1060 VDD.n610 19.3944
R13175 VDD.n1060 VDD.n608 19.3944
R13176 VDD.n1318 VDD.n608 19.3944
R13177 VDD.n2152 VDD.n237 19.3944
R13178 VDD.n2152 VDD.n235 19.3944
R13179 VDD.n2156 VDD.n235 19.3944
R13180 VDD.n2156 VDD.n226 19.3944
R13181 VDD.n2168 VDD.n226 19.3944
R13182 VDD.n2168 VDD.n224 19.3944
R13183 VDD.n2172 VDD.n224 19.3944
R13184 VDD.n2172 VDD.n214 19.3944
R13185 VDD.n2184 VDD.n214 19.3944
R13186 VDD.n2184 VDD.n212 19.3944
R13187 VDD.n2188 VDD.n212 19.3944
R13188 VDD.n2188 VDD.n202 19.3944
R13189 VDD.n2200 VDD.n202 19.3944
R13190 VDD.n2200 VDD.n200 19.3944
R13191 VDD.n2204 VDD.n200 19.3944
R13192 VDD.n2204 VDD.n188 19.3944
R13193 VDD.n2216 VDD.n188 19.3944
R13194 VDD.n2216 VDD.n186 19.3944
R13195 VDD.n2220 VDD.n186 19.3944
R13196 VDD.n2221 VDD.n2220 19.3944
R13197 VDD.n2222 VDD.n2221 19.3944
R13198 VDD.n2222 VDD.n184 19.3944
R13199 VDD.n2226 VDD.n184 19.3944
R13200 VDD.n2227 VDD.n2226 19.3944
R13201 VDD.n2228 VDD.n2227 19.3944
R13202 VDD.n2228 VDD.n181 19.3944
R13203 VDD.n2232 VDD.n181 19.3944
R13204 VDD.n2233 VDD.n2232 19.3944
R13205 VDD.n2234 VDD.n2233 19.3944
R13206 VDD.n2234 VDD.n178 19.3944
R13207 VDD.n2238 VDD.n178 19.3944
R13208 VDD.n2239 VDD.n2238 19.3944
R13209 VDD.n2240 VDD.n2239 19.3944
R13210 VDD.n2240 VDD.n175 19.3944
R13211 VDD.n2244 VDD.n175 19.3944
R13212 VDD.n2245 VDD.n2244 19.3944
R13213 VDD.n2246 VDD.n2245 19.3944
R13214 VDD.n2270 VDD.n149 19.3944
R13215 VDD.n2265 VDD.n149 19.3944
R13216 VDD.n2265 VDD.n2264 19.3944
R13217 VDD.n2264 VDD.n2263 19.3944
R13218 VDD.n2263 VDD.n156 19.3944
R13219 VDD.n2258 VDD.n156 19.3944
R13220 VDD.n2258 VDD.n2257 19.3944
R13221 VDD.n2257 VDD.n2256 19.3944
R13222 VDD.n2256 VDD.n163 19.3944
R13223 VDD.n2251 VDD.n163 19.3944
R13224 VDD.n2294 VDD.n128 19.3944
R13225 VDD.n2289 VDD.n128 19.3944
R13226 VDD.n2289 VDD.n2288 19.3944
R13227 VDD.n2288 VDD.n2287 19.3944
R13228 VDD.n2287 VDD.n135 19.3944
R13229 VDD.n2282 VDD.n135 19.3944
R13230 VDD.n2282 VDD.n2281 19.3944
R13231 VDD.n2281 VDD.n2280 19.3944
R13232 VDD.n2280 VDD.n142 19.3944
R13233 VDD.n2275 VDD.n142 19.3944
R13234 VDD.n2275 VDD.n2274 19.3944
R13235 VDD.n2318 VDD.n107 19.3944
R13236 VDD.n2313 VDD.n107 19.3944
R13237 VDD.n2313 VDD.n2312 19.3944
R13238 VDD.n2312 VDD.n2311 19.3944
R13239 VDD.n2311 VDD.n114 19.3944
R13240 VDD.n2306 VDD.n114 19.3944
R13241 VDD.n2306 VDD.n2305 19.3944
R13242 VDD.n2305 VDD.n2304 19.3944
R13243 VDD.n2304 VDD.n121 19.3944
R13244 VDD.n2299 VDD.n121 19.3944
R13245 VDD.n2299 VDD.n2298 19.3944
R13246 VDD.n2337 VDD.n2336 19.3944
R13247 VDD.n2336 VDD.n2335 19.3944
R13248 VDD.n2335 VDD.n93 19.3944
R13249 VDD.n2330 VDD.n93 19.3944
R13250 VDD.n2330 VDD.n2329 19.3944
R13251 VDD.n2329 VDD.n2328 19.3944
R13252 VDD.n2328 VDD.n100 19.3944
R13253 VDD.n2323 VDD.n100 19.3944
R13254 VDD.n2323 VDD.n2322 19.3944
R13255 VDD.n2148 VDD.n242 19.3944
R13256 VDD.n2148 VDD.n232 19.3944
R13257 VDD.n2160 VDD.n232 19.3944
R13258 VDD.n2160 VDD.n230 19.3944
R13259 VDD.n2164 VDD.n230 19.3944
R13260 VDD.n2164 VDD.n220 19.3944
R13261 VDD.n2176 VDD.n220 19.3944
R13262 VDD.n2176 VDD.n218 19.3944
R13263 VDD.n2180 VDD.n218 19.3944
R13264 VDD.n2180 VDD.n208 19.3944
R13265 VDD.n2192 VDD.n208 19.3944
R13266 VDD.n2192 VDD.n206 19.3944
R13267 VDD.n2196 VDD.n206 19.3944
R13268 VDD.n2196 VDD.n196 19.3944
R13269 VDD.n2208 VDD.n196 19.3944
R13270 VDD.n2208 VDD.n194 19.3944
R13271 VDD.n2212 VDD.n194 19.3944
R13272 VDD.n2212 VDD.n37 19.3944
R13273 VDD.n2378 VDD.n37 19.3944
R13274 VDD.n2378 VDD.n38 19.3944
R13275 VDD.n2372 VDD.n38 19.3944
R13276 VDD.n2372 VDD.n2371 19.3944
R13277 VDD.n2371 VDD.n2370 19.3944
R13278 VDD.n2370 VDD.n49 19.3944
R13279 VDD.n2364 VDD.n49 19.3944
R13280 VDD.n2364 VDD.n2363 19.3944
R13281 VDD.n2363 VDD.n2362 19.3944
R13282 VDD.n2362 VDD.n60 19.3944
R13283 VDD.n2356 VDD.n60 19.3944
R13284 VDD.n2356 VDD.n2355 19.3944
R13285 VDD.n2355 VDD.n2354 19.3944
R13286 VDD.n2354 VDD.n71 19.3944
R13287 VDD.n2348 VDD.n71 19.3944
R13288 VDD.n2348 VDD.n2347 19.3944
R13289 VDD.n2347 VDD.n2346 19.3944
R13290 VDD.n2346 VDD.n82 19.3944
R13291 VDD.n2340 VDD.n82 19.3944
R13292 VDD.n2095 VDD.n2092 19.3944
R13293 VDD.n2092 VDD.n2091 19.3944
R13294 VDD.n2091 VDD.n2088 19.3944
R13295 VDD.n2088 VDD.n2087 19.3944
R13296 VDD.n2087 VDD.n2084 19.3944
R13297 VDD.n2084 VDD.n2083 19.3944
R13298 VDD.n2083 VDD.n2080 19.3944
R13299 VDD.n2080 VDD.n2079 19.3944
R13300 VDD.n2079 VDD.n2076 19.3944
R13301 VDD.n2076 VDD.n2075 19.3944
R13302 VDD.n2075 VDD.n2072 19.3944
R13303 VDD.n2122 VDD.n2119 19.3944
R13304 VDD.n2119 VDD.n2118 19.3944
R13305 VDD.n2118 VDD.n2115 19.3944
R13306 VDD.n2115 VDD.n2114 19.3944
R13307 VDD.n2114 VDD.n2111 19.3944
R13308 VDD.n2111 VDD.n2110 19.3944
R13309 VDD.n2110 VDD.n2107 19.3944
R13310 VDD.n2107 VDD.n2106 19.3944
R13311 VDD.n2106 VDD.n2103 19.3944
R13312 VDD.n2103 VDD.n2102 19.3944
R13313 VDD.n2102 VDD.n2099 19.3944
R13314 VDD.n2144 VDD.n244 19.3944
R13315 VDD.n2139 VDD.n244 19.3944
R13316 VDD.n2139 VDD.n2138 19.3944
R13317 VDD.n2138 VDD.n2137 19.3944
R13318 VDD.n2134 VDD.n2133 19.3944
R13319 VDD.n2130 VDD.n2129 19.3944
R13320 VDD.n2129 VDD.n2126 19.3944
R13321 VDD.n2068 VDD.n2065 19.3944
R13322 VDD.n2065 VDD.n2064 19.3944
R13323 VDD.n2064 VDD.n2061 19.3944
R13324 VDD.n2061 VDD.n2060 19.3944
R13325 VDD.n2060 VDD.n2057 19.3944
R13326 VDD.n2038 VDD.n304 19.3944
R13327 VDD.n2053 VDD.n2052 19.3944
R13328 VDD.n2052 VDD.n2050 19.3944
R13329 VDD.n834 VDD.n833 19.2005
R13330 VDD.n1326 VDD.n1325 19.2005
R13331 VDD.n2251 VDD.n2250 19.2005
R13332 VDD.n2050 VDD.n2047 19.2005
R13333 VDD.n918 VDD.n734 17.5931
R13334 VDD.n918 VDD.n735 17.5931
R13335 VDD.n926 VDD.n723 17.5931
R13336 VDD.n934 VDD.n723 17.5931
R13337 VDD.n934 VDD.n717 17.5931
R13338 VDD.n942 VDD.n717 17.5931
R13339 VDD.n942 VDD.n711 17.5931
R13340 VDD.n950 VDD.n711 17.5931
R13341 VDD.n958 VDD.n705 17.5931
R13342 VDD.n958 VDD.n699 17.5931
R13343 VDD.n966 VDD.n699 17.5931
R13344 VDD.n974 VDD.n693 17.5931
R13345 VDD.n974 VDD.n686 17.5931
R13346 VDD.n983 VDD.n686 17.5931
R13347 VDD.n983 VDD.n687 17.5931
R13348 VDD.n991 VDD.n655 17.5931
R13349 VDD.n999 VDD.n655 17.5931
R13350 VDD.n999 VDD.n649 17.5931
R13351 VDD.n1007 VDD.n649 17.5931
R13352 VDD.n1015 VDD.n643 17.5931
R13353 VDD.n1015 VDD.n637 17.5931
R13354 VDD.n1023 VDD.n637 17.5931
R13355 VDD.n1031 VDD.n631 17.5931
R13356 VDD.n1031 VDD.n625 17.5931
R13357 VDD.n1039 VDD.n625 17.5931
R13358 VDD.n1039 VDD.n618 17.5931
R13359 VDD.n1047 VDD.n618 17.5931
R13360 VDD.n1047 VDD.n619 17.5931
R13361 VDD.n1058 VDD.n605 17.5931
R13362 VDD.n1320 VDD.n605 17.5931
R13363 VDD.n2150 VDD.n239 17.5931
R13364 VDD.n2150 VDD.n240 17.5931
R13365 VDD.n2158 VDD.n228 17.5931
R13366 VDD.n2166 VDD.n228 17.5931
R13367 VDD.n2166 VDD.n222 17.5931
R13368 VDD.n2174 VDD.n222 17.5931
R13369 VDD.n2174 VDD.n216 17.5931
R13370 VDD.n2182 VDD.n216 17.5931
R13371 VDD.n2190 VDD.n210 17.5931
R13372 VDD.n2190 VDD.n204 17.5931
R13373 VDD.n2198 VDD.n204 17.5931
R13374 VDD.n2206 VDD.n198 17.5931
R13375 VDD.n2206 VDD.n191 17.5931
R13376 VDD.n2214 VDD.n191 17.5931
R13377 VDD.n2214 VDD.n192 17.5931
R13378 VDD.n2376 VDD.n2375 17.5931
R13379 VDD.n2375 VDD.n2374 17.5931
R13380 VDD.n2374 VDD.n44 17.5931
R13381 VDD.n2368 VDD.n44 17.5931
R13382 VDD.n2367 VDD.n2366 17.5931
R13383 VDD.n2366 VDD.n54 17.5931
R13384 VDD.n2360 VDD.n54 17.5931
R13385 VDD.n2359 VDD.n2358 17.5931
R13386 VDD.n2358 VDD.n65 17.5931
R13387 VDD.n2352 VDD.n65 17.5931
R13388 VDD.n2352 VDD.n2351 17.5931
R13389 VDD.n2351 VDD.n2350 17.5931
R13390 VDD.n2350 VDD.n76 17.5931
R13391 VDD.n2344 VDD.n2343 17.5931
R13392 VDD.n2343 VDD.n2342 17.5931
R13393 VDD.t82 VDD.n705 15.1301
R13394 VDD.n1023 VDD.t86 15.1301
R13395 VDD.t96 VDD.n210 15.1301
R13396 VDD.n2360 VDD.t108 15.1301
R13397 VDD.n966 VDD.t98 14.4264
R13398 VDD.t100 VDD.n643 14.4264
R13399 VDD.n2198 VDD.t94 14.4264
R13400 VDD.t90 VDD.n2367 14.4264
R13401 VDD.n926 VDD.t21 12.6672
R13402 VDD.n619 VDD.t6 12.6672
R13403 VDD.n2158 VDD.t17 12.6672
R13404 VDD.t25 VDD.n76 12.6672
R13405 VDD.n1426 VDD.n576 11.9635
R13406 VDD.n1432 VDD.n576 11.9635
R13407 VDD.n1432 VDD.n569 11.9635
R13408 VDD.n1438 VDD.n569 11.9635
R13409 VDD.n1438 VDD.n572 11.9635
R13410 VDD.n1444 VDD.n558 11.9635
R13411 VDD.n1450 VDD.n558 11.9635
R13412 VDD.n1450 VDD.n552 11.9635
R13413 VDD.n1456 VDD.n552 11.9635
R13414 VDD.n1456 VDD.n546 11.9635
R13415 VDD.n1462 VDD.n546 11.9635
R13416 VDD.n1462 VDD.n540 11.9635
R13417 VDD.n1468 VDD.n540 11.9635
R13418 VDD.n1474 VDD.n533 11.9635
R13419 VDD.n1474 VDD.n536 11.9635
R13420 VDD.n1480 VDD.n522 11.9635
R13421 VDD.n1486 VDD.n522 11.9635
R13422 VDD.n1486 VDD.n515 11.9635
R13423 VDD.n1492 VDD.n515 11.9635
R13424 VDD.n1492 VDD.n518 11.9635
R13425 VDD.n1498 VDD.n504 11.9635
R13426 VDD.n1504 VDD.n504 11.9635
R13427 VDD.n1504 VDD.n496 11.9635
R13428 VDD.n1512 VDD.n496 11.9635
R13429 VDD.n1512 VDD.n499 11.9635
R13430 VDD.n1518 VDD.n481 11.9635
R13431 VDD.n1576 VDD.n481 11.9635
R13432 VDD.n1582 VDD.n475 11.9635
R13433 VDD.n1582 VDD.n444 11.9635
R13434 VDD.n1836 VDD.n438 11.9635
R13435 VDD.n1842 VDD.n438 11.9635
R13436 VDD.n1848 VDD.n431 11.9635
R13437 VDD.n1848 VDD.n434 11.9635
R13438 VDD.n1854 VDD.n420 11.9635
R13439 VDD.n1860 VDD.n420 11.9635
R13440 VDD.n1860 VDD.n413 11.9635
R13441 VDD.n1866 VDD.n413 11.9635
R13442 VDD.n1866 VDD.n416 11.9635
R13443 VDD.n1872 VDD.n402 11.9635
R13444 VDD.n1878 VDD.n402 11.9635
R13445 VDD.n1878 VDD.n395 11.9635
R13446 VDD.n1884 VDD.n395 11.9635
R13447 VDD.n1884 VDD.n398 11.9635
R13448 VDD.n1890 VDD.n384 11.9635
R13449 VDD.n1896 VDD.n384 11.9635
R13450 VDD.n1902 VDD.n378 11.9635
R13451 VDD.n1902 VDD.n372 11.9635
R13452 VDD.n1908 VDD.n372 11.9635
R13453 VDD.n1908 VDD.n366 11.9635
R13454 VDD.n1914 VDD.n366 11.9635
R13455 VDD.n1914 VDD.n359 11.9635
R13456 VDD.n1920 VDD.n359 11.9635
R13457 VDD.n1920 VDD.n362 11.9635
R13458 VDD.n1956 VDD.n347 11.9635
R13459 VDD.n1962 VDD.n347 11.9635
R13460 VDD.n1962 VDD.n322 11.9635
R13461 VDD.n2012 VDD.n322 11.9635
R13462 VDD.n2012 VDD.n324 11.9635
R13463 VDD.n1429 VDD.n1428 10.6151
R13464 VDD.n1430 VDD.n1429 10.6151
R13465 VDD.n1430 VDD.n567 10.6151
R13466 VDD.n1440 VDD.n567 10.6151
R13467 VDD.n1441 VDD.n1440 10.6151
R13468 VDD.n1442 VDD.n1441 10.6151
R13469 VDD.n1442 VDD.n556 10.6151
R13470 VDD.n1452 VDD.n556 10.6151
R13471 VDD.n1453 VDD.n1452 10.6151
R13472 VDD.n1454 VDD.n1453 10.6151
R13473 VDD.n1454 VDD.n544 10.6151
R13474 VDD.n1464 VDD.n544 10.6151
R13475 VDD.n1465 VDD.n1464 10.6151
R13476 VDD.n1466 VDD.n1465 10.6151
R13477 VDD.n1466 VDD.n531 10.6151
R13478 VDD.n1476 VDD.n531 10.6151
R13479 VDD.n1477 VDD.n1476 10.6151
R13480 VDD.n1478 VDD.n1477 10.6151
R13481 VDD.n1478 VDD.n520 10.6151
R13482 VDD.n1488 VDD.n520 10.6151
R13483 VDD.n1489 VDD.n1488 10.6151
R13484 VDD.n1490 VDD.n1489 10.6151
R13485 VDD.n1490 VDD.n508 10.6151
R13486 VDD.n1500 VDD.n508 10.6151
R13487 VDD.n1501 VDD.n1500 10.6151
R13488 VDD.n1502 VDD.n1501 10.6151
R13489 VDD.n1502 VDD.n494 10.6151
R13490 VDD.n1514 VDD.n494 10.6151
R13491 VDD.n1515 VDD.n1514 10.6151
R13492 VDD.n1516 VDD.n1515 10.6151
R13493 VDD.n1516 VDD.n479 10.6151
R13494 VDD.n1578 VDD.n479 10.6151
R13495 VDD.n1579 VDD.n1578 10.6151
R13496 VDD.n1580 VDD.n1579 10.6151
R13497 VDD.n1580 VDD.n468 10.6151
R13498 VDD.n1624 VDD.n1623 10.6151
R13499 VDD.n1623 VDD.n1622 10.6151
R13500 VDD.n1622 VDD.n1619 10.6151
R13501 VDD.n1619 VDD.n1618 10.6151
R13502 VDD.n1618 VDD.n1615 10.6151
R13503 VDD.n1615 VDD.n1614 10.6151
R13504 VDD.n1614 VDD.n1611 10.6151
R13505 VDD.n1611 VDD.n1610 10.6151
R13506 VDD.n1610 VDD.n1607 10.6151
R13507 VDD.n1607 VDD.n1606 10.6151
R13508 VDD.n1606 VDD.n1603 10.6151
R13509 VDD.n1603 VDD.n1602 10.6151
R13510 VDD.n1602 VDD.n1599 10.6151
R13511 VDD.n1599 VDD.n1598 10.6151
R13512 VDD.n1598 VDD.n1595 10.6151
R13513 VDD.n1595 VDD.n1594 10.6151
R13514 VDD.n1594 VDD.n1591 10.6151
R13515 VDD.n1591 VDD.n1590 10.6151
R13516 VDD.n1587 VDD.n1586 10.6151
R13517 VDD.n1281 VDD.n1280 10.6151
R13518 VDD.n1280 VDD.n1278 10.6151
R13519 VDD.n1278 VDD.n1277 10.6151
R13520 VDD.n1277 VDD.n1275 10.6151
R13521 VDD.n1275 VDD.n1274 10.6151
R13522 VDD.n1274 VDD.n1272 10.6151
R13523 VDD.n1272 VDD.n1271 10.6151
R13524 VDD.n1271 VDD.n1269 10.6151
R13525 VDD.n1269 VDD.n1268 10.6151
R13526 VDD.n1268 VDD.n1266 10.6151
R13527 VDD.n1266 VDD.n1265 10.6151
R13528 VDD.n1265 VDD.n1263 10.6151
R13529 VDD.n1263 VDD.n1262 10.6151
R13530 VDD.n1262 VDD.n1260 10.6151
R13531 VDD.n1260 VDD.n1259 10.6151
R13532 VDD.n1259 VDD.n1257 10.6151
R13533 VDD.n1257 VDD.n1256 10.6151
R13534 VDD.n1256 VDD.n1254 10.6151
R13535 VDD.n1254 VDD.n1253 10.6151
R13536 VDD.n1253 VDD.n1251 10.6151
R13537 VDD.n1251 VDD.n1250 10.6151
R13538 VDD.n1250 VDD.n1248 10.6151
R13539 VDD.n1248 VDD.n1247 10.6151
R13540 VDD.n1247 VDD.n1245 10.6151
R13541 VDD.n1245 VDD.n1244 10.6151
R13542 VDD.n1244 VDD.n1242 10.6151
R13543 VDD.n1242 VDD.n1241 10.6151
R13544 VDD.n1241 VDD.n1239 10.6151
R13545 VDD.n1239 VDD.n1238 10.6151
R13546 VDD.n1238 VDD.n1236 10.6151
R13547 VDD.n1236 VDD.n1235 10.6151
R13548 VDD.n1235 VDD.n1233 10.6151
R13549 VDD.n1233 VDD.n1232 10.6151
R13550 VDD.n1232 VDD.n474 10.6151
R13551 VDD.n474 VDD.n472 10.6151
R13552 VDD.n1207 VDD.n580 10.6151
R13553 VDD.n1208 VDD.n1207 10.6151
R13554 VDD.n1209 VDD.n1208 10.6151
R13555 VDD.n1209 VDD.n1203 10.6151
R13556 VDD.n1215 VDD.n1203 10.6151
R13557 VDD.n1216 VDD.n1215 10.6151
R13558 VDD.n1217 VDD.n1216 10.6151
R13559 VDD.n1217 VDD.n1201 10.6151
R13560 VDD.n1201 VDD.n1200 10.6151
R13561 VDD.n1302 VDD.n1200 10.6151
R13562 VDD.n1302 VDD.n1301 10.6151
R13563 VDD.n1301 VDD.n1224 10.6151
R13564 VDD.n1296 VDD.n1224 10.6151
R13565 VDD.n1296 VDD.n1295 10.6151
R13566 VDD.n1295 VDD.n1226 10.6151
R13567 VDD.n1290 VDD.n1226 10.6151
R13568 VDD.n1290 VDD.n1289 10.6151
R13569 VDD.n1289 VDD.n1288 10.6151
R13570 VDD.n1284 VDD.n1283 10.6151
R13571 VDD.n1791 VDD.n1790 10.6151
R13572 VDD.n1790 VDD.n1788 10.6151
R13573 VDD.n1788 VDD.n1787 10.6151
R13574 VDD.n1787 VDD.n1785 10.6151
R13575 VDD.n1785 VDD.n1784 10.6151
R13576 VDD.n1784 VDD.n1782 10.6151
R13577 VDD.n1782 VDD.n1781 10.6151
R13578 VDD.n1781 VDD.n1779 10.6151
R13579 VDD.n1779 VDD.n1778 10.6151
R13580 VDD.n1778 VDD.n1776 10.6151
R13581 VDD.n1776 VDD.n1775 10.6151
R13582 VDD.n1775 VDD.n1773 10.6151
R13583 VDD.n1773 VDD.n1772 10.6151
R13584 VDD.n1772 VDD.n1770 10.6151
R13585 VDD.n1770 VDD.n1769 10.6151
R13586 VDD.n1769 VDD.n1767 10.6151
R13587 VDD.n1767 VDD.n1766 10.6151
R13588 VDD.n1766 VDD.n1764 10.6151
R13589 VDD.n1764 VDD.n1763 10.6151
R13590 VDD.n1763 VDD.n1761 10.6151
R13591 VDD.n1761 VDD.n1760 10.6151
R13592 VDD.n1760 VDD.n1758 10.6151
R13593 VDD.n1758 VDD.n1757 10.6151
R13594 VDD.n1757 VDD.n1755 10.6151
R13595 VDD.n1755 VDD.n1754 10.6151
R13596 VDD.n1754 VDD.n1752 10.6151
R13597 VDD.n1752 VDD.n1751 10.6151
R13598 VDD.n1751 VDD.n1749 10.6151
R13599 VDD.n1749 VDD.n1748 10.6151
R13600 VDD.n1748 VDD.n1746 10.6151
R13601 VDD.n1746 VDD.n1745 10.6151
R13602 VDD.n1745 VDD.n345 10.6151
R13603 VDD.n1965 VDD.n345 10.6151
R13604 VDD.n1966 VDD.n1965 10.6151
R13605 VDD.n1967 VDD.n1966 10.6151
R13606 VDD.n1833 VDD.n1832 10.6151
R13607 VDD.n1832 VDD.n1733 10.6151
R13608 VDD.n1827 VDD.n1733 10.6151
R13609 VDD.n1827 VDD.n1826 10.6151
R13610 VDD.n1826 VDD.n1735 10.6151
R13611 VDD.n1821 VDD.n1735 10.6151
R13612 VDD.n1821 VDD.n1820 10.6151
R13613 VDD.n1820 VDD.n1819 10.6151
R13614 VDD.n1819 VDD.n1737 10.6151
R13615 VDD.n1813 VDD.n1737 10.6151
R13616 VDD.n1813 VDD.n1812 10.6151
R13617 VDD.n1812 VDD.n1811 10.6151
R13618 VDD.n1811 VDD.n1739 10.6151
R13619 VDD.n1805 VDD.n1739 10.6151
R13620 VDD.n1805 VDD.n1804 10.6151
R13621 VDD.n1804 VDD.n1803 10.6151
R13622 VDD.n1803 VDD.n1741 10.6151
R13623 VDD.n1797 VDD.n1741 10.6151
R13624 VDD.n1795 VDD.n1794 10.6151
R13625 VDD.n1834 VDD.n436 10.6151
R13626 VDD.n1844 VDD.n436 10.6151
R13627 VDD.n1845 VDD.n1844 10.6151
R13628 VDD.n1846 VDD.n1845 10.6151
R13629 VDD.n1846 VDD.n424 10.6151
R13630 VDD.n1856 VDD.n424 10.6151
R13631 VDD.n1857 VDD.n1856 10.6151
R13632 VDD.n1858 VDD.n1857 10.6151
R13633 VDD.n1858 VDD.n411 10.6151
R13634 VDD.n1868 VDD.n411 10.6151
R13635 VDD.n1869 VDD.n1868 10.6151
R13636 VDD.n1870 VDD.n1869 10.6151
R13637 VDD.n1870 VDD.n400 10.6151
R13638 VDD.n1880 VDD.n400 10.6151
R13639 VDD.n1881 VDD.n1880 10.6151
R13640 VDD.n1882 VDD.n1881 10.6151
R13641 VDD.n1882 VDD.n388 10.6151
R13642 VDD.n1892 VDD.n388 10.6151
R13643 VDD.n1893 VDD.n1892 10.6151
R13644 VDD.n1894 VDD.n1893 10.6151
R13645 VDD.n1894 VDD.n376 10.6151
R13646 VDD.n1904 VDD.n376 10.6151
R13647 VDD.n1905 VDD.n1904 10.6151
R13648 VDD.n1906 VDD.n1905 10.6151
R13649 VDD.n1906 VDD.n364 10.6151
R13650 VDD.n1916 VDD.n364 10.6151
R13651 VDD.n1917 VDD.n1916 10.6151
R13652 VDD.n1918 VDD.n1917 10.6151
R13653 VDD.n1918 VDD.n351 10.6151
R13654 VDD.n1958 VDD.n351 10.6151
R13655 VDD.n1959 VDD.n1958 10.6151
R13656 VDD.n1960 VDD.n1959 10.6151
R13657 VDD.n1960 VDD.n328 10.6151
R13658 VDD.n2010 VDD.n328 10.6151
R13659 VDD.n2010 VDD.n2009 10.6151
R13660 VDD.n2008 VDD.n329 10.6151
R13661 VDD.n2003 VDD.n329 10.6151
R13662 VDD.n2003 VDD.n2002 10.6151
R13663 VDD.n2002 VDD.n2001 10.6151
R13664 VDD.n2001 VDD.n331 10.6151
R13665 VDD.n1996 VDD.n331 10.6151
R13666 VDD.n1996 VDD.n1995 10.6151
R13667 VDD.n1995 VDD.n1994 10.6151
R13668 VDD.n1994 VDD.n334 10.6151
R13669 VDD.n1989 VDD.n334 10.6151
R13670 VDD.n1989 VDD.n1987 10.6151
R13671 VDD.n1987 VDD.n1986 10.6151
R13672 VDD.n1986 VDD.n337 10.6151
R13673 VDD.n1981 VDD.n337 10.6151
R13674 VDD.n1981 VDD.n1980 10.6151
R13675 VDD.n1980 VDD.n1979 10.6151
R13676 VDD.n1979 VDD.n340 10.6151
R13677 VDD.n1974 VDD.n340 10.6151
R13678 VDD.n1972 VDD.n1971 10.6151
R13679 VDD.n1925 VDD.n1924 10.6151
R13680 VDD.n1942 VDD.n1925 10.6151
R13681 VDD.n1942 VDD.n1941 10.6151
R13682 VDD.n1941 VDD.n1940 10.6151
R13683 VDD.n1940 VDD.n1927 10.6151
R13684 VDD.n1935 VDD.n1927 10.6151
R13685 VDD.n1935 VDD.n1934 10.6151
R13686 VDD.n1934 VDD.n1933 10.6151
R13687 VDD.n1933 VDD.n306 10.6151
R13688 VDD.n2035 VDD.n306 10.6151
R13689 VDD.n2035 VDD.n307 10.6151
R13690 VDD.n2030 VDD.n307 10.6151
R13691 VDD.n2030 VDD.n2029 10.6151
R13692 VDD.n2029 VDD.n2028 10.6151
R13693 VDD.n2028 VDD.n311 10.6151
R13694 VDD.n2023 VDD.n311 10.6151
R13695 VDD.n2023 VDD.n2022 10.6151
R13696 VDD.n2022 VDD.n2021 10.6151
R13697 VDD.n2016 VDD.n318 10.6151
R13698 VDD.n1730 VDD.n1729 10.6151
R13699 VDD.n1729 VDD.n1728 10.6151
R13700 VDD.n1728 VDD.n1727 10.6151
R13701 VDD.n1727 VDD.n1725 10.6151
R13702 VDD.n1725 VDD.n1724 10.6151
R13703 VDD.n1724 VDD.n1722 10.6151
R13704 VDD.n1722 VDD.n1721 10.6151
R13705 VDD.n1721 VDD.n1719 10.6151
R13706 VDD.n1719 VDD.n1718 10.6151
R13707 VDD.n1718 VDD.n1716 10.6151
R13708 VDD.n1716 VDD.n1715 10.6151
R13709 VDD.n1715 VDD.n1713 10.6151
R13710 VDD.n1713 VDD.n1712 10.6151
R13711 VDD.n1712 VDD.n1710 10.6151
R13712 VDD.n1710 VDD.n1709 10.6151
R13713 VDD.n1709 VDD.n1707 10.6151
R13714 VDD.n1707 VDD.n1706 10.6151
R13715 VDD.n1706 VDD.n1704 10.6151
R13716 VDD.n1704 VDD.n1703 10.6151
R13717 VDD.n1703 VDD.n1701 10.6151
R13718 VDD.n1701 VDD.n1700 10.6151
R13719 VDD.n1700 VDD.n1698 10.6151
R13720 VDD.n1698 VDD.n1697 10.6151
R13721 VDD.n1697 VDD.n1695 10.6151
R13722 VDD.n1695 VDD.n1694 10.6151
R13723 VDD.n1694 VDD.n1692 10.6151
R13724 VDD.n1692 VDD.n1691 10.6151
R13725 VDD.n1691 VDD.n1689 10.6151
R13726 VDD.n1689 VDD.n1688 10.6151
R13727 VDD.n1688 VDD.n1686 10.6151
R13728 VDD.n1686 VDD.n1685 10.6151
R13729 VDD.n1685 VDD.n1683 10.6151
R13730 VDD.n1683 VDD.n320 10.6151
R13731 VDD.n2014 VDD.n320 10.6151
R13732 VDD.n2015 VDD.n2014 10.6151
R13733 VDD.n1644 VDD.n442 10.6151
R13734 VDD.n1645 VDD.n1644 10.6151
R13735 VDD.n1645 VDD.n1641 10.6151
R13736 VDD.n1651 VDD.n1641 10.6151
R13737 VDD.n1652 VDD.n1651 10.6151
R13738 VDD.n1653 VDD.n1652 10.6151
R13739 VDD.n1653 VDD.n1639 10.6151
R13740 VDD.n1659 VDD.n1639 10.6151
R13741 VDD.n1660 VDD.n1659 10.6151
R13742 VDD.n1661 VDD.n1660 10.6151
R13743 VDD.n1661 VDD.n1637 10.6151
R13744 VDD.n1667 VDD.n1637 10.6151
R13745 VDD.n1668 VDD.n1667 10.6151
R13746 VDD.n1669 VDD.n1668 10.6151
R13747 VDD.n1669 VDD.n1635 10.6151
R13748 VDD.n1675 VDD.n1635 10.6151
R13749 VDD.n1676 VDD.n1675 10.6151
R13750 VDD.n1677 VDD.n1676 10.6151
R13751 VDD.n1682 VDD.n1681 10.6151
R13752 VDD.n1839 VDD.n1838 10.6151
R13753 VDD.n1840 VDD.n1839 10.6151
R13754 VDD.n1840 VDD.n429 10.6151
R13755 VDD.n1850 VDD.n429 10.6151
R13756 VDD.n1851 VDD.n1850 10.6151
R13757 VDD.n1852 VDD.n1851 10.6151
R13758 VDD.n1852 VDD.n418 10.6151
R13759 VDD.n1862 VDD.n418 10.6151
R13760 VDD.n1863 VDD.n1862 10.6151
R13761 VDD.n1864 VDD.n1863 10.6151
R13762 VDD.n1864 VDD.n406 10.6151
R13763 VDD.n1874 VDD.n406 10.6151
R13764 VDD.n1875 VDD.n1874 10.6151
R13765 VDD.n1876 VDD.n1875 10.6151
R13766 VDD.n1876 VDD.n393 10.6151
R13767 VDD.n1886 VDD.n393 10.6151
R13768 VDD.n1887 VDD.n1886 10.6151
R13769 VDD.n1888 VDD.n1887 10.6151
R13770 VDD.n1888 VDD.n382 10.6151
R13771 VDD.n1898 VDD.n382 10.6151
R13772 VDD.n1899 VDD.n1898 10.6151
R13773 VDD.n1900 VDD.n1899 10.6151
R13774 VDD.n1900 VDD.n370 10.6151
R13775 VDD.n1910 VDD.n370 10.6151
R13776 VDD.n1911 VDD.n1910 10.6151
R13777 VDD.n1912 VDD.n1911 10.6151
R13778 VDD.n1912 VDD.n357 10.6151
R13779 VDD.n1922 VDD.n357 10.6151
R13780 VDD.n1923 VDD.n1922 10.6151
R13781 VDD.n1954 VDD.n1923 10.6151
R13782 VDD.n1954 VDD.n1953 10.6151
R13783 VDD.n1953 VDD.n1952 10.6151
R13784 VDD.n1952 VDD.n1951 10.6151
R13785 VDD.n1951 VDD.n1949 10.6151
R13786 VDD.n1949 VDD.n1948 10.6151
R13787 VDD.n1424 VDD.n574 10.6151
R13788 VDD.n1434 VDD.n574 10.6151
R13789 VDD.n1435 VDD.n1434 10.6151
R13790 VDD.n1436 VDD.n1435 10.6151
R13791 VDD.n1436 VDD.n562 10.6151
R13792 VDD.n1446 VDD.n562 10.6151
R13793 VDD.n1447 VDD.n1446 10.6151
R13794 VDD.n1448 VDD.n1447 10.6151
R13795 VDD.n1448 VDD.n550 10.6151
R13796 VDD.n1458 VDD.n550 10.6151
R13797 VDD.n1459 VDD.n1458 10.6151
R13798 VDD.n1460 VDD.n1459 10.6151
R13799 VDD.n1460 VDD.n538 10.6151
R13800 VDD.n1470 VDD.n538 10.6151
R13801 VDD.n1471 VDD.n1470 10.6151
R13802 VDD.n1472 VDD.n1471 10.6151
R13803 VDD.n1472 VDD.n526 10.6151
R13804 VDD.n1482 VDD.n526 10.6151
R13805 VDD.n1483 VDD.n1482 10.6151
R13806 VDD.n1484 VDD.n1483 10.6151
R13807 VDD.n1484 VDD.n513 10.6151
R13808 VDD.n1494 VDD.n513 10.6151
R13809 VDD.n1495 VDD.n1494 10.6151
R13810 VDD.n1496 VDD.n1495 10.6151
R13811 VDD.n1496 VDD.n502 10.6151
R13812 VDD.n1506 VDD.n502 10.6151
R13813 VDD.n1507 VDD.n1506 10.6151
R13814 VDD.n1510 VDD.n1507 10.6151
R13815 VDD.n1510 VDD.n1509 10.6151
R13816 VDD.n1509 VDD.n1508 10.6151
R13817 VDD.n1508 VDD.n486 10.6151
R13818 VDD.n1574 VDD.n486 10.6151
R13819 VDD.n1574 VDD.n1573 10.6151
R13820 VDD.n1573 VDD.n1572 10.6151
R13821 VDD.n1572 VDD.n1571 10.6151
R13822 VDD.n1568 VDD.n1567 10.6151
R13823 VDD.n1567 VDD.n1564 10.6151
R13824 VDD.n1564 VDD.n1563 10.6151
R13825 VDD.n1563 VDD.n1560 10.6151
R13826 VDD.n1560 VDD.n1559 10.6151
R13827 VDD.n1559 VDD.n1556 10.6151
R13828 VDD.n1556 VDD.n1555 10.6151
R13829 VDD.n1555 VDD.n1552 10.6151
R13830 VDD.n1552 VDD.n1551 10.6151
R13831 VDD.n1551 VDD.n1548 10.6151
R13832 VDD.n1548 VDD.n1547 10.6151
R13833 VDD.n1547 VDD.n1544 10.6151
R13834 VDD.n1544 VDD.n1543 10.6151
R13835 VDD.n1543 VDD.n1540 10.6151
R13836 VDD.n1540 VDD.n1539 10.6151
R13837 VDD.n1539 VDD.n1536 10.6151
R13838 VDD.n1536 VDD.n1535 10.6151
R13839 VDD.n1535 VDD.n1532 10.6151
R13840 VDD.n1530 VDD.n1528 10.6151
R13841 VDD.n1382 VDD.n1381 10.6151
R13842 VDD.n1381 VDD.n1379 10.6151
R13843 VDD.n1379 VDD.n1378 10.6151
R13844 VDD.n1378 VDD.n1376 10.6151
R13845 VDD.n1376 VDD.n1375 10.6151
R13846 VDD.n1375 VDD.n1373 10.6151
R13847 VDD.n1373 VDD.n1372 10.6151
R13848 VDD.n1372 VDD.n1370 10.6151
R13849 VDD.n1370 VDD.n1369 10.6151
R13850 VDD.n1369 VDD.n1367 10.6151
R13851 VDD.n1367 VDD.n1366 10.6151
R13852 VDD.n1366 VDD.n1364 10.6151
R13853 VDD.n1364 VDD.n1363 10.6151
R13854 VDD.n1363 VDD.n1361 10.6151
R13855 VDD.n1361 VDD.n1360 10.6151
R13856 VDD.n1360 VDD.n1358 10.6151
R13857 VDD.n1358 VDD.n1357 10.6151
R13858 VDD.n1357 VDD.n1355 10.6151
R13859 VDD.n1355 VDD.n1354 10.6151
R13860 VDD.n1354 VDD.n1352 10.6151
R13861 VDD.n1352 VDD.n1351 10.6151
R13862 VDD.n1351 VDD.n1349 10.6151
R13863 VDD.n1349 VDD.n1348 10.6151
R13864 VDD.n1348 VDD.n1346 10.6151
R13865 VDD.n1346 VDD.n1345 10.6151
R13866 VDD.n1345 VDD.n1343 10.6151
R13867 VDD.n1343 VDD.n1342 10.6151
R13868 VDD.n1342 VDD.n1340 10.6151
R13869 VDD.n1340 VDD.n1339 10.6151
R13870 VDD.n1339 VDD.n489 10.6151
R13871 VDD.n1521 VDD.n489 10.6151
R13872 VDD.n1522 VDD.n1521 10.6151
R13873 VDD.n1524 VDD.n1522 10.6151
R13874 VDD.n1525 VDD.n1524 10.6151
R13875 VDD.n1527 VDD.n1525 10.6151
R13876 VDD.n1423 VDD.n1422 10.6151
R13877 VDD.n1422 VDD.n586 10.6151
R13878 VDD.n1416 VDD.n586 10.6151
R13879 VDD.n1416 VDD.n1415 10.6151
R13880 VDD.n1415 VDD.n1414 10.6151
R13881 VDD.n1414 VDD.n588 10.6151
R13882 VDD.n1408 VDD.n588 10.6151
R13883 VDD.n1408 VDD.n1407 10.6151
R13884 VDD.n1407 VDD.n1406 10.6151
R13885 VDD.n1406 VDD.n1330 10.6151
R13886 VDD.n1400 VDD.n1330 10.6151
R13887 VDD.n1400 VDD.n1399 10.6151
R13888 VDD.n1399 VDD.n1398 10.6151
R13889 VDD.n1398 VDD.n1332 10.6151
R13890 VDD.n1392 VDD.n1332 10.6151
R13891 VDD.n1392 VDD.n1391 10.6151
R13892 VDD.n1391 VDD.n1390 10.6151
R13893 VDD.n1390 VDD.n1334 10.6151
R13894 VDD.n1384 VDD.n1383 10.6151
R13895 VDD.n1305 VDD.n1302 10.5971
R13896 VDD.n1989 VDD.n1988 10.5971
R13897 VDD.n2055 VDD.n2035 10.5971
R13898 VDD.n1330 VDD.n1329 10.5971
R13899 VDD.n1140 VDD.n1115 9.3005
R13900 VDD.n1119 VDD.n1116 9.3005
R13901 VDD.n1135 VDD.n1120 9.3005
R13902 VDD.n1134 VDD.n1121 9.3005
R13903 VDD.n1133 VDD.n590 9.3005
R13904 VDD.n1164 VDD.n1094 9.3005
R13905 VDD.n1098 VDD.n1095 9.3005
R13906 VDD.n1159 VDD.n1099 9.3005
R13907 VDD.n1158 VDD.n1100 9.3005
R13908 VDD.n1157 VDD.n1101 9.3005
R13909 VDD.n1105 VDD.n1102 9.3005
R13910 VDD.n1152 VDD.n1106 9.3005
R13911 VDD.n1151 VDD.n1107 9.3005
R13912 VDD.n1150 VDD.n1108 9.3005
R13913 VDD.n1112 VDD.n1109 9.3005
R13914 VDD.n1145 VDD.n1113 9.3005
R13915 VDD.n1144 VDD.n1114 9.3005
R13916 VDD.n1188 VDD.n1073 9.3005
R13917 VDD.n1077 VDD.n1074 9.3005
R13918 VDD.n1183 VDD.n1078 9.3005
R13919 VDD.n1182 VDD.n1079 9.3005
R13920 VDD.n1181 VDD.n1080 9.3005
R13921 VDD.n1084 VDD.n1081 9.3005
R13922 VDD.n1176 VDD.n1085 9.3005
R13923 VDD.n1175 VDD.n1086 9.3005
R13924 VDD.n1174 VDD.n1087 9.3005
R13925 VDD.n1091 VDD.n1088 9.3005
R13926 VDD.n1169 VDD.n1092 9.3005
R13927 VDD.n1168 VDD.n1093 9.3005
R13928 VDD.n1193 VDD.n1068 9.3005
R13929 VDD.n1192 VDD.n1072 9.3005
R13930 VDD.n1314 VDD.n1063 9.3005
R13931 VDD.n1303 VDD.n1064 9.3005
R13932 VDD.n1304 VDD.n1065 9.3005
R13933 VDD.n1316 VDD.n1315 9.3005
R13934 VDD.n994 VDD.n993 9.3005
R13935 VDD.n995 VDD.n657 9.3005
R13936 VDD.n997 VDD.n996 9.3005
R13937 VDD.n647 VDD.n646 9.3005
R13938 VDD.n1010 VDD.n1009 9.3005
R13939 VDD.n1011 VDD.n645 9.3005
R13940 VDD.n1013 VDD.n1012 9.3005
R13941 VDD.n635 VDD.n634 9.3005
R13942 VDD.n1026 VDD.n1025 9.3005
R13943 VDD.n1027 VDD.n633 9.3005
R13944 VDD.n1029 VDD.n1028 9.3005
R13945 VDD.n623 VDD.n622 9.3005
R13946 VDD.n1042 VDD.n1041 9.3005
R13947 VDD.n1043 VDD.n621 9.3005
R13948 VDD.n1045 VDD.n1044 9.3005
R13949 VDD.n610 VDD.n609 9.3005
R13950 VDD.n1061 VDD.n1060 9.3005
R13951 VDD.n1062 VDD.n608 9.3005
R13952 VDD.n1318 VDD.n1317 9.3005
R13953 VDD.n2075 VDD.n297 9.3005
R13954 VDD.n2076 VDD.n296 9.3005
R13955 VDD.n2079 VDD.n295 9.3005
R13956 VDD.n2080 VDD.n294 9.3005
R13957 VDD.n2083 VDD.n293 9.3005
R13958 VDD.n2084 VDD.n292 9.3005
R13959 VDD.n2087 VDD.n291 9.3005
R13960 VDD.n2088 VDD.n290 9.3005
R13961 VDD.n2091 VDD.n289 9.3005
R13962 VDD.n2092 VDD.n288 9.3005
R13963 VDD.n2095 VDD.n287 9.3005
R13964 VDD.n2072 VDD.n298 9.3005
R13965 VDD.n2102 VDD.n285 9.3005
R13966 VDD.n2103 VDD.n284 9.3005
R13967 VDD.n2106 VDD.n283 9.3005
R13968 VDD.n2107 VDD.n282 9.3005
R13969 VDD.n2110 VDD.n281 9.3005
R13970 VDD.n2111 VDD.n280 9.3005
R13971 VDD.n2114 VDD.n279 9.3005
R13972 VDD.n2115 VDD.n278 9.3005
R13973 VDD.n2118 VDD.n277 9.3005
R13974 VDD.n2119 VDD.n276 9.3005
R13975 VDD.n2122 VDD.n275 9.3005
R13976 VDD.n2099 VDD.n286 9.3005
R13977 VDD.n2126 VDD.n274 9.3005
R13978 VDD.n2129 VDD.n273 9.3005
R13979 VDD.n2138 VDD.n270 9.3005
R13980 VDD.n2139 VDD.n269 9.3005
R13981 VDD.n244 VDD.n243 9.3005
R13982 VDD.n2145 VDD.n2144 9.3005
R13983 VDD.n2148 VDD.n2147 9.3005
R13984 VDD.n232 VDD.n231 9.3005
R13985 VDD.n2161 VDD.n2160 9.3005
R13986 VDD.n2162 VDD.n230 9.3005
R13987 VDD.n2164 VDD.n2163 9.3005
R13988 VDD.n220 VDD.n219 9.3005
R13989 VDD.n2177 VDD.n2176 9.3005
R13990 VDD.n2178 VDD.n218 9.3005
R13991 VDD.n2180 VDD.n2179 9.3005
R13992 VDD.n208 VDD.n207 9.3005
R13993 VDD.n2193 VDD.n2192 9.3005
R13994 VDD.n2194 VDD.n206 9.3005
R13995 VDD.n2196 VDD.n2195 9.3005
R13996 VDD.n196 VDD.n195 9.3005
R13997 VDD.n2209 VDD.n2208 9.3005
R13998 VDD.n2210 VDD.n194 9.3005
R13999 VDD.n2212 VDD.n2211 9.3005
R14000 VDD.n37 VDD.n35 9.3005
R14001 VDD.n2146 VDD.n242 9.3005
R14002 VDD.n2379 VDD.n2378 9.3005
R14003 VDD.n38 VDD.n36 9.3005
R14004 VDD.n2372 VDD.n46 9.3005
R14005 VDD.n2371 VDD.n47 9.3005
R14006 VDD.n2370 VDD.n48 9.3005
R14007 VDD.n56 VDD.n49 9.3005
R14008 VDD.n2364 VDD.n57 9.3005
R14009 VDD.n2363 VDD.n58 9.3005
R14010 VDD.n2362 VDD.n59 9.3005
R14011 VDD.n67 VDD.n60 9.3005
R14012 VDD.n2356 VDD.n68 9.3005
R14013 VDD.n2355 VDD.n69 9.3005
R14014 VDD.n2354 VDD.n70 9.3005
R14015 VDD.n78 VDD.n71 9.3005
R14016 VDD.n2348 VDD.n79 9.3005
R14017 VDD.n2347 VDD.n80 9.3005
R14018 VDD.n2346 VDD.n81 9.3005
R14019 VDD.n89 VDD.n82 9.3005
R14020 VDD.n2340 VDD.n2339 9.3005
R14021 VDD.n2336 VDD.n90 9.3005
R14022 VDD.n2335 VDD.n92 9.3005
R14023 VDD.n96 VDD.n93 9.3005
R14024 VDD.n2330 VDD.n97 9.3005
R14025 VDD.n2329 VDD.n98 9.3005
R14026 VDD.n2328 VDD.n99 9.3005
R14027 VDD.n103 VDD.n100 9.3005
R14028 VDD.n2323 VDD.n104 9.3005
R14029 VDD.n2322 VDD.n105 9.3005
R14030 VDD.n2318 VDD.n106 9.3005
R14031 VDD.n110 VDD.n107 9.3005
R14032 VDD.n2313 VDD.n111 9.3005
R14033 VDD.n2312 VDD.n112 9.3005
R14034 VDD.n2311 VDD.n113 9.3005
R14035 VDD.n117 VDD.n114 9.3005
R14036 VDD.n2306 VDD.n118 9.3005
R14037 VDD.n2305 VDD.n119 9.3005
R14038 VDD.n2304 VDD.n120 9.3005
R14039 VDD.n124 VDD.n121 9.3005
R14040 VDD.n2299 VDD.n125 9.3005
R14041 VDD.n2298 VDD.n126 9.3005
R14042 VDD.n2294 VDD.n127 9.3005
R14043 VDD.n131 VDD.n128 9.3005
R14044 VDD.n2289 VDD.n132 9.3005
R14045 VDD.n2288 VDD.n133 9.3005
R14046 VDD.n2287 VDD.n134 9.3005
R14047 VDD.n138 VDD.n135 9.3005
R14048 VDD.n2282 VDD.n139 9.3005
R14049 VDD.n2281 VDD.n140 9.3005
R14050 VDD.n2280 VDD.n141 9.3005
R14051 VDD.n145 VDD.n142 9.3005
R14052 VDD.n2275 VDD.n146 9.3005
R14053 VDD.n2274 VDD.n147 9.3005
R14054 VDD.n2270 VDD.n148 9.3005
R14055 VDD.n152 VDD.n149 9.3005
R14056 VDD.n2265 VDD.n153 9.3005
R14057 VDD.n2264 VDD.n154 9.3005
R14058 VDD.n2263 VDD.n155 9.3005
R14059 VDD.n159 VDD.n156 9.3005
R14060 VDD.n2258 VDD.n160 9.3005
R14061 VDD.n2257 VDD.n161 9.3005
R14062 VDD.n2256 VDD.n162 9.3005
R14063 VDD.n166 VDD.n163 9.3005
R14064 VDD.n2251 VDD.n167 9.3005
R14065 VDD.n2250 VDD.n2249 9.3005
R14066 VDD.n2248 VDD.n170 9.3005
R14067 VDD.n2338 VDD.n2337 9.3005
R14068 VDD.n2153 VDD.n2152 9.3005
R14069 VDD.n2154 VDD.n235 9.3005
R14070 VDD.n2156 VDD.n2155 9.3005
R14071 VDD.n226 VDD.n225 9.3005
R14072 VDD.n2169 VDD.n2168 9.3005
R14073 VDD.n2170 VDD.n224 9.3005
R14074 VDD.n2172 VDD.n2171 9.3005
R14075 VDD.n214 VDD.n213 9.3005
R14076 VDD.n2185 VDD.n2184 9.3005
R14077 VDD.n2186 VDD.n212 9.3005
R14078 VDD.n2188 VDD.n2187 9.3005
R14079 VDD.n202 VDD.n201 9.3005
R14080 VDD.n2201 VDD.n2200 9.3005
R14081 VDD.n2202 VDD.n200 9.3005
R14082 VDD.n2204 VDD.n2203 9.3005
R14083 VDD.n188 VDD.n187 9.3005
R14084 VDD.n2217 VDD.n2216 9.3005
R14085 VDD.n2218 VDD.n186 9.3005
R14086 VDD.n2220 VDD.n2219 9.3005
R14087 VDD.n2221 VDD.n185 9.3005
R14088 VDD.n2223 VDD.n2222 9.3005
R14089 VDD.n2224 VDD.n184 9.3005
R14090 VDD.n2226 VDD.n2225 9.3005
R14091 VDD.n2227 VDD.n182 9.3005
R14092 VDD.n2229 VDD.n2228 9.3005
R14093 VDD.n2230 VDD.n181 9.3005
R14094 VDD.n2232 VDD.n2231 9.3005
R14095 VDD.n2233 VDD.n179 9.3005
R14096 VDD.n2235 VDD.n2234 9.3005
R14097 VDD.n2236 VDD.n178 9.3005
R14098 VDD.n2238 VDD.n2237 9.3005
R14099 VDD.n2239 VDD.n176 9.3005
R14100 VDD.n2241 VDD.n2240 9.3005
R14101 VDD.n2242 VDD.n175 9.3005
R14102 VDD.n2244 VDD.n2243 9.3005
R14103 VDD.n2245 VDD.n173 9.3005
R14104 VDD.n2247 VDD.n2246 9.3005
R14105 VDD.n237 VDD.n236 9.3005
R14106 VDD.n2043 VDD.n2042 9.3005
R14107 VDD.n2047 VDD.n2044 9.3005
R14108 VDD.n2050 VDD.n2040 9.3005
R14109 VDD.n2052 VDD.n305 9.3005
R14110 VDD.n2060 VDD.n303 9.3005
R14111 VDD.n2061 VDD.n302 9.3005
R14112 VDD.n2064 VDD.n301 9.3005
R14113 VDD.n2065 VDD.n300 9.3005
R14114 VDD.n2068 VDD.n299 9.3005
R14115 VDD.n1328 VDD.n1327 9.3005
R14116 VDD.n1326 VDD.n593 9.3005
R14117 VDD.n1325 VDD.n600 9.3005
R14118 VDD.n1052 VDD.n597 9.3005
R14119 VDD.n921 VDD.n920 9.3005
R14120 VDD.n922 VDD.n730 9.3005
R14121 VDD.n924 VDD.n923 9.3005
R14122 VDD.n721 VDD.n720 9.3005
R14123 VDD.n937 VDD.n936 9.3005
R14124 VDD.n938 VDD.n719 9.3005
R14125 VDD.n940 VDD.n939 9.3005
R14126 VDD.n709 VDD.n708 9.3005
R14127 VDD.n953 VDD.n952 9.3005
R14128 VDD.n954 VDD.n707 9.3005
R14129 VDD.n956 VDD.n955 9.3005
R14130 VDD.n697 VDD.n696 9.3005
R14131 VDD.n969 VDD.n968 9.3005
R14132 VDD.n970 VDD.n695 9.3005
R14133 VDD.n972 VDD.n971 9.3005
R14134 VDD.n684 VDD.n683 9.3005
R14135 VDD.n986 VDD.n985 9.3005
R14136 VDD.n987 VDD.n682 9.3005
R14137 VDD.n989 VDD.n988 9.3005
R14138 VDD.n653 VDD.n652 9.3005
R14139 VDD.n1002 VDD.n1001 9.3005
R14140 VDD.n1003 VDD.n651 9.3005
R14141 VDD.n1005 VDD.n1004 9.3005
R14142 VDD.n641 VDD.n640 9.3005
R14143 VDD.n1018 VDD.n1017 9.3005
R14144 VDD.n1019 VDD.n639 9.3005
R14145 VDD.n1021 VDD.n1020 9.3005
R14146 VDD.n629 VDD.n628 9.3005
R14147 VDD.n1034 VDD.n1033 9.3005
R14148 VDD.n1035 VDD.n627 9.3005
R14149 VDD.n1037 VDD.n1036 9.3005
R14150 VDD.n616 VDD.n615 9.3005
R14151 VDD.n1050 VDD.n1049 9.3005
R14152 VDD.n1051 VDD.n613 9.3005
R14153 VDD.n1056 VDD.n1055 9.3005
R14154 VDD.n1054 VDD.n614 9.3005
R14155 VDD.n1053 VDD.n604 9.3005
R14156 VDD.n732 VDD.n731 9.3005
R14157 VDD.n835 VDD.n834 9.3005
R14158 VDD.n836 VDD.n824 9.3005
R14159 VDD.n838 VDD.n837 9.3005
R14160 VDD.n839 VDD.n819 9.3005
R14161 VDD.n841 VDD.n840 9.3005
R14162 VDD.n842 VDD.n818 9.3005
R14163 VDD.n844 VDD.n843 9.3005
R14164 VDD.n845 VDD.n813 9.3005
R14165 VDD.n847 VDD.n846 9.3005
R14166 VDD.n848 VDD.n812 9.3005
R14167 VDD.n850 VDD.n849 9.3005
R14168 VDD.n856 VDD.n855 9.3005
R14169 VDD.n857 VDD.n806 9.3005
R14170 VDD.n859 VDD.n858 9.3005
R14171 VDD.n860 VDD.n801 9.3005
R14172 VDD.n862 VDD.n861 9.3005
R14173 VDD.n863 VDD.n800 9.3005
R14174 VDD.n865 VDD.n864 9.3005
R14175 VDD.n866 VDD.n795 9.3005
R14176 VDD.n868 VDD.n867 9.3005
R14177 VDD.n869 VDD.n794 9.3005
R14178 VDD.n871 VDD.n870 9.3005
R14179 VDD.n877 VDD.n876 9.3005
R14180 VDD.n878 VDD.n788 9.3005
R14181 VDD.n880 VDD.n879 9.3005
R14182 VDD.n881 VDD.n783 9.3005
R14183 VDD.n883 VDD.n882 9.3005
R14184 VDD.n884 VDD.n782 9.3005
R14185 VDD.n886 VDD.n885 9.3005
R14186 VDD.n887 VDD.n777 9.3005
R14187 VDD.n889 VDD.n888 9.3005
R14188 VDD.n890 VDD.n776 9.3005
R14189 VDD.n892 VDD.n891 9.3005
R14190 VDD.n896 VDD.n771 9.3005
R14191 VDD.n898 VDD.n897 9.3005
R14192 VDD.n899 VDD.n770 9.3005
R14193 VDD.n901 VDD.n900 9.3005
R14194 VDD.n902 VDD.n765 9.3005
R14195 VDD.n904 VDD.n903 9.3005
R14196 VDD.n905 VDD.n764 9.3005
R14197 VDD.n907 VDD.n906 9.3005
R14198 VDD.n739 VDD.n738 9.3005
R14199 VDD.n913 VDD.n912 9.3005
R14200 VDD.n875 VDD.n789 9.3005
R14201 VDD.n854 VDD.n807 9.3005
R14202 VDD.n833 VDD.n825 9.3005
R14203 VDD.n829 VDD.n828 9.3005
R14204 VDD.n916 VDD.n915 9.3005
R14205 VDD.n727 VDD.n726 9.3005
R14206 VDD.n929 VDD.n928 9.3005
R14207 VDD.n930 VDD.n725 9.3005
R14208 VDD.n932 VDD.n931 9.3005
R14209 VDD.n715 VDD.n714 9.3005
R14210 VDD.n945 VDD.n944 9.3005
R14211 VDD.n946 VDD.n713 9.3005
R14212 VDD.n948 VDD.n947 9.3005
R14213 VDD.n703 VDD.n702 9.3005
R14214 VDD.n961 VDD.n960 9.3005
R14215 VDD.n962 VDD.n701 9.3005
R14216 VDD.n964 VDD.n963 9.3005
R14217 VDD.n691 VDD.n690 9.3005
R14218 VDD.n977 VDD.n976 9.3005
R14219 VDD.n978 VDD.n689 9.3005
R14220 VDD.n981 VDD.n980 9.3005
R14221 VDD.n979 VDD.n679 9.3005
R14222 VDD.n914 VDD.n737 9.3005
R14223 VDD.n687 VDD.t88 8.7968
R14224 VDD.n991 VDD.t88 8.7968
R14225 VDD.n192 VDD.t130 8.7968
R14226 VDD.n2376 VDD.t130 8.7968
R14227 VDD.n31 VDD.t135 8.7384
R14228 VDD.n31 VDD.t151 8.7384
R14229 VDD.n30 VDD.t97 8.7384
R14230 VDD.n30 VDD.t116 8.7384
R14231 VDD.n26 VDD.t161 8.7384
R14232 VDD.n26 VDD.t91 8.7384
R14233 VDD.n25 VDD.t126 8.7384
R14234 VDD.n25 VDD.t150 8.7384
R14235 VDD.n21 VDD.t155 8.7384
R14236 VDD.n21 VDD.t140 8.7384
R14237 VDD.n20 VDD.t134 8.7384
R14238 VDD.n20 VDD.t123 8.7384
R14239 VDD.n17 VDD.t131 8.7384
R14240 VDD.n17 VDD.t122 8.7384
R14241 VDD.n16 VDD.t113 8.7384
R14242 VDD.n16 VDD.t95 8.7384
R14243 VDD.n672 VDD.t89 8.7384
R14244 VDD.n672 VDD.t154 8.7384
R14245 VDD.n674 VDD.t146 8.7384
R14246 VDD.n674 VDD.t107 8.7384
R14247 VDD.n667 VDD.t125 8.7384
R14248 VDD.n667 VDD.t110 8.7384
R14249 VDD.n669 VDD.t83 8.7384
R14250 VDD.n669 VDD.t129 8.7384
R14251 VDD.n662 VDD.t142 8.7384
R14252 VDD.n662 VDD.t101 8.7384
R14253 VDD.n664 VDD.t164 8.7384
R14254 VDD.n664 VDD.t124 8.7384
R14255 VDD.n658 VDD.t115 8.7384
R14256 VDD.n658 VDD.t156 8.7384
R14257 VDD.n660 VDD.t149 8.7384
R14258 VDD.n660 VDD.t99 8.7384
R14259 VDD.n666 VDD.n661 8.41429
R14260 VDD.n15 VDD.n14 8.25626
R14261 VDD.n2381 VDD.n2380 8.08313
R14262 VDD.n678 VDD.n677 8.08313
R14263 VDD.n1468 VDD.t117 7.91717
R14264 VDD.t147 VDD.n378 7.91717
R14265 VDD.n499 VDD.t10 7.74124
R14266 VDD.n1854 VDD.t2 7.74124
R14267 VDD.n24 VDD.n19 7.40567
R14268 VDD.n518 VDD.t92 7.21346
R14269 VDD.n1872 VDD.t152 7.21346
R14270 VDD.n833 VDD.n829 6.78838
R14271 VDD.n1325 VDD.n597 6.78838
R14272 VDD.n2047 VDD.n2042 6.78838
R14273 VDD.n2250 VDD.n170 6.78838
R14274 VDD.n1576 VDD.t132 6.50976
R14275 VDD.t136 VDD.n431 6.50976
R14276 VDD.n7 VDD.t85 6.5015
R14277 VDD.n7 VDD.t106 6.5015
R14278 VDD.n8 VDD.t145 6.5015
R14279 VDD.n8 VDD.t128 6.5015
R14280 VDD.n10 VDD.t148 6.5015
R14281 VDD.n10 VDD.t160 6.5015
R14282 VDD.n12 VDD.t137 6.5015
R14283 VDD.n12 VDD.t153 6.5015
R14284 VDD.n5 VDD.t93 6.5015
R14285 VDD.n5 VDD.t133 6.5015
R14286 VDD.n3 VDD.t112 6.5015
R14287 VDD.n3 VDD.t118 6.5015
R14288 VDD.n1 VDD.t104 6.5015
R14289 VDD.n1 VDD.t163 6.5015
R14290 VDD.n0 VDD.t139 6.5015
R14291 VDD.n0 VDD.t120 6.5015
R14292 VDD.n853 VDD.n850 6.4005
R14293 VDD.n874 VDD.n871 6.4005
R14294 VDD.n1143 VDD.n1140 6.4005
R14295 VDD.n1167 VDD.n1164 6.4005
R14296 VDD.n2273 VDD.n2270 6.4005
R14297 VDD.n2297 VDD.n2294 6.4005
R14298 VDD.n2098 VDD.n2095 6.4005
R14299 VDD.n2071 VDD.n2068 6.4005
R14300 VDD.n1590 VDD.n471 6.0883
R14301 VDD.n1288 VDD.n1230 6.0883
R14302 VDD.n1797 VDD.n1796 6.0883
R14303 VDD.n1974 VDD.n1973 6.0883
R14304 VDD.n2021 VDD.n316 6.0883
R14305 VDD.n1677 VDD.n1633 6.0883
R14306 VDD.n1532 VDD.n1531 6.0883
R14307 VDD.n1338 VDD.n1334 6.0883
R14308 VDD.n895 VDD.n892 6.01262
R14309 VDD.n1191 VDD.n1188 6.01262
R14310 VDD.n2321 VDD.n2318 6.01262
R14311 VDD.n2125 VDD.n2122 6.01262
R14312 VDD.n536 VDD.t102 5.98198
R14313 VDD.n1480 VDD.t102 5.98198
R14314 VDD.n398 VDD.t121 5.98198
R14315 VDD.n1890 VDD.t121 5.98198
R14316 VDD.n676 VDD.n675 5.89274
R14317 VDD.n671 VDD.n670 5.89274
R14318 VDD.n666 VDD.n665 5.89274
R14319 VDD.t132 VDD.n475 5.4542
R14320 VDD.n1842 VDD.t136 5.4542
R14321 VDD.n2381 VDD.n34 5.08553
R14322 VDD.n677 VDD.n676 5.08553
R14323 VDD.n735 VDD.t21 4.92643
R14324 VDD.n1058 VDD.t6 4.92643
R14325 VDD.n240 VDD.t17 4.92643
R14326 VDD.n2344 VDD.t25 4.92643
R14327 VDD.n34 VDD.n33 4.88412
R14328 VDD.n29 VDD.n28 4.88412
R14329 VDD.n24 VDD.n23 4.88412
R14330 VDD.n1498 VDD.t92 4.7505
R14331 VDD.n416 VDD.t152 4.7505
R14332 VDD.n1122 VDD.n591 4.74817
R14333 VDD.n1127 VDD.n592 4.74817
R14334 VDD.n1307 VDD.n1306 4.74817
R14335 VDD.n1199 VDD.n1069 4.74817
R14336 VDD.n1306 VDD.n1067 4.74817
R14337 VDD.n1199 VDD.n1198 4.74817
R14338 VDD.n2137 VDD.n271 4.74817
R14339 VDD.n2130 VDD.n272 4.74817
R14340 VDD.n2133 VDD.n272 4.74817
R14341 VDD.n2134 VDD.n271 4.74817
R14342 VDD.n2056 VDD.n304 4.74817
R14343 VDD.n2054 VDD.n2053 4.74817
R14344 VDD.n2054 VDD.n2038 4.74817
R14345 VDD.n2057 VDD.n2056 4.74817
R14346 VDD.n1128 VDD.n591 4.74817
R14347 VDD.n594 VDD.n592 4.74817
R14348 VDD.n1587 VDD.n471 4.52733
R14349 VDD.n1284 VDD.n1230 4.52733
R14350 VDD.n1796 VDD.n1795 4.52733
R14351 VDD.n1973 VDD.n1972 4.52733
R14352 VDD.n318 VDD.n316 4.52733
R14353 VDD.n1681 VDD.n1633 4.52733
R14354 VDD.n1531 VDD.n1530 4.52733
R14355 VDD.n1384 VDD.n1338 4.52733
R14356 VDD.t69 VDD.t111 4.39865
R14357 VDD.t159 VDD.t44 4.39865
R14358 VDD.n572 VDD.t69 4.22272
R14359 VDD.n1518 VDD.t10 4.22272
R14360 VDD.n434 VDD.t2 4.22272
R14361 VDD.n1956 VDD.t44 4.22272
R14362 VDD.t117 VDD.n533 4.0468
R14363 VDD.n1896 VDD.t147 4.0468
R14364 VDD.n1444 VDD.t111 3.34309
R14365 VDD.n362 VDD.t159 3.34309
R14366 VDD.n11 VDD.n9 3.29576
R14367 VDD.n4 VDD.n2 3.29576
R14368 VDD.t98 VDD.n693 3.16717
R14369 VDD.n1007 VDD.t100 3.16717
R14370 VDD.t94 VDD.n198 3.16717
R14371 VDD.n2368 VDD.t90 3.16717
R14372 VDD.n13 VDD.n11 2.62119
R14373 VDD.n6 VDD.n4 2.62119
R14374 VDD.n29 VDD.n24 2.52636
R14375 VDD.n671 VDD.n666 2.52636
R14376 VDD.n34 VDD.n29 2.52205
R14377 VDD.n676 VDD.n671 2.52205
R14378 VDD.n950 VDD.t82 2.46346
R14379 VDD.t86 VDD.n631 2.46346
R14380 VDD.n2182 VDD.t96 2.46346
R14381 VDD.t108 VDD.n2359 2.46346
R14382 VDD.n1306 VDD.n1305 2.27742
R14383 VDD.n1305 VDD.n1199 2.27742
R14384 VDD.n1988 VDD.n272 2.27742
R14385 VDD.n1988 VDD.n271 2.27742
R14386 VDD.n2055 VDD.n2054 2.27742
R14387 VDD.n2056 VDD.n2055 2.27742
R14388 VDD.n1329 VDD.n591 2.27742
R14389 VDD.n1329 VDD.n592 2.27742
R14390 VDD.n14 VDD.n13 2.04939
R14391 VDD.n14 VDD.n6 2.04939
R14392 VDD.n33 VDD.n32 2.01774
R14393 VDD.n28 VDD.n27 2.01774
R14394 VDD.n23 VDD.n22 2.01774
R14395 VDD.n19 VDD.n18 2.01774
R14396 VDD.n675 VDD.n673 2.01774
R14397 VDD.n670 VDD.n668 2.01774
R14398 VDD.n665 VDD.n663 2.01774
R14399 VDD.n661 VDD.n659 2.01774
R14400 VDD.n677 VDD.n15 1.4116
R14401 VDD VDD.n2381 1.40376
R14402 VDD.n896 VDD.n895 0.582318
R14403 VDD.n1192 VDD.n1191 0.582318
R14404 VDD.n2322 VDD.n2321 0.582318
R14405 VDD.n2126 VDD.n2125 0.582318
R14406 VDD.n1317 VDD.n1316 0.523366
R14407 VDD.n2146 VDD.n2145 0.523366
R14408 VDD.n2339 VDD.n2338 0.523366
R14409 VDD.n2248 VDD.n2247 0.523366
R14410 VDD.n2043 VDD.n236 0.523366
R14411 VDD.n1053 VDD.n1052 0.523366
R14412 VDD.n828 VDD.n731 0.523366
R14413 VDD.n914 VDD.n913 0.523366
R14414 VDD.n854 VDD.n853 0.194439
R14415 VDD.n875 VDD.n874 0.194439
R14416 VDD.n1144 VDD.n1143 0.194439
R14417 VDD.n1168 VDD.n1167 0.194439
R14418 VDD.n2274 VDD.n2273 0.194439
R14419 VDD.n2298 VDD.n2297 0.194439
R14420 VDD.n2072 VDD.n2071 0.194439
R14421 VDD.n2099 VDD.n2098 0.194439
R14422 VDD.n1072 VDD.n1068 0.152939
R14423 VDD.n1073 VDD.n1072 0.152939
R14424 VDD.n1077 VDD.n1073 0.152939
R14425 VDD.n1078 VDD.n1077 0.152939
R14426 VDD.n1079 VDD.n1078 0.152939
R14427 VDD.n1080 VDD.n1079 0.152939
R14428 VDD.n1084 VDD.n1080 0.152939
R14429 VDD.n1085 VDD.n1084 0.152939
R14430 VDD.n1086 VDD.n1085 0.152939
R14431 VDD.n1087 VDD.n1086 0.152939
R14432 VDD.n1091 VDD.n1087 0.152939
R14433 VDD.n1092 VDD.n1091 0.152939
R14434 VDD.n1093 VDD.n1092 0.152939
R14435 VDD.n1094 VDD.n1093 0.152939
R14436 VDD.n1098 VDD.n1094 0.152939
R14437 VDD.n1099 VDD.n1098 0.152939
R14438 VDD.n1100 VDD.n1099 0.152939
R14439 VDD.n1101 VDD.n1100 0.152939
R14440 VDD.n1105 VDD.n1101 0.152939
R14441 VDD.n1106 VDD.n1105 0.152939
R14442 VDD.n1107 VDD.n1106 0.152939
R14443 VDD.n1108 VDD.n1107 0.152939
R14444 VDD.n1112 VDD.n1108 0.152939
R14445 VDD.n1113 VDD.n1112 0.152939
R14446 VDD.n1114 VDD.n1113 0.152939
R14447 VDD.n1115 VDD.n1114 0.152939
R14448 VDD.n1119 VDD.n1115 0.152939
R14449 VDD.n1120 VDD.n1119 0.152939
R14450 VDD.n1121 VDD.n1120 0.152939
R14451 VDD.n1121 VDD.n590 0.152939
R14452 VDD.n1316 VDD.n1063 0.152939
R14453 VDD.n1303 VDD.n1063 0.152939
R14454 VDD.n1304 VDD.n1303 0.152939
R14455 VDD.n995 VDD.n994 0.152939
R14456 VDD.n996 VDD.n995 0.152939
R14457 VDD.n996 VDD.n646 0.152939
R14458 VDD.n1010 VDD.n646 0.152939
R14459 VDD.n1011 VDD.n1010 0.152939
R14460 VDD.n1012 VDD.n1011 0.152939
R14461 VDD.n1012 VDD.n634 0.152939
R14462 VDD.n1026 VDD.n634 0.152939
R14463 VDD.n1027 VDD.n1026 0.152939
R14464 VDD.n1028 VDD.n1027 0.152939
R14465 VDD.n1028 VDD.n622 0.152939
R14466 VDD.n1042 VDD.n622 0.152939
R14467 VDD.n1043 VDD.n1042 0.152939
R14468 VDD.n1044 VDD.n1043 0.152939
R14469 VDD.n1044 VDD.n609 0.152939
R14470 VDD.n1061 VDD.n609 0.152939
R14471 VDD.n1062 VDD.n1061 0.152939
R14472 VDD.n1317 VDD.n1062 0.152939
R14473 VDD.n274 VDD.n273 0.152939
R14474 VDD.n275 VDD.n274 0.152939
R14475 VDD.n276 VDD.n275 0.152939
R14476 VDD.n277 VDD.n276 0.152939
R14477 VDD.n278 VDD.n277 0.152939
R14478 VDD.n279 VDD.n278 0.152939
R14479 VDD.n280 VDD.n279 0.152939
R14480 VDD.n281 VDD.n280 0.152939
R14481 VDD.n282 VDD.n281 0.152939
R14482 VDD.n283 VDD.n282 0.152939
R14483 VDD.n284 VDD.n283 0.152939
R14484 VDD.n285 VDD.n284 0.152939
R14485 VDD.n286 VDD.n285 0.152939
R14486 VDD.n287 VDD.n286 0.152939
R14487 VDD.n288 VDD.n287 0.152939
R14488 VDD.n289 VDD.n288 0.152939
R14489 VDD.n290 VDD.n289 0.152939
R14490 VDD.n291 VDD.n290 0.152939
R14491 VDD.n292 VDD.n291 0.152939
R14492 VDD.n293 VDD.n292 0.152939
R14493 VDD.n294 VDD.n293 0.152939
R14494 VDD.n295 VDD.n294 0.152939
R14495 VDD.n296 VDD.n295 0.152939
R14496 VDD.n297 VDD.n296 0.152939
R14497 VDD.n298 VDD.n297 0.152939
R14498 VDD.n299 VDD.n298 0.152939
R14499 VDD.n300 VDD.n299 0.152939
R14500 VDD.n301 VDD.n300 0.152939
R14501 VDD.n302 VDD.n301 0.152939
R14502 VDD.n303 VDD.n302 0.152939
R14503 VDD.n2145 VDD.n243 0.152939
R14504 VDD.n269 VDD.n243 0.152939
R14505 VDD.n270 VDD.n269 0.152939
R14506 VDD.n2147 VDD.n2146 0.152939
R14507 VDD.n2147 VDD.n231 0.152939
R14508 VDD.n2161 VDD.n231 0.152939
R14509 VDD.n2162 VDD.n2161 0.152939
R14510 VDD.n2163 VDD.n2162 0.152939
R14511 VDD.n2163 VDD.n219 0.152939
R14512 VDD.n2177 VDD.n219 0.152939
R14513 VDD.n2178 VDD.n2177 0.152939
R14514 VDD.n2179 VDD.n2178 0.152939
R14515 VDD.n2179 VDD.n207 0.152939
R14516 VDD.n2193 VDD.n207 0.152939
R14517 VDD.n2194 VDD.n2193 0.152939
R14518 VDD.n2195 VDD.n2194 0.152939
R14519 VDD.n2195 VDD.n195 0.152939
R14520 VDD.n2209 VDD.n195 0.152939
R14521 VDD.n2210 VDD.n2209 0.152939
R14522 VDD.n2211 VDD.n2210 0.152939
R14523 VDD.n2211 VDD.n35 0.152939
R14524 VDD.n2379 VDD.n36 0.152939
R14525 VDD.n46 VDD.n36 0.152939
R14526 VDD.n47 VDD.n46 0.152939
R14527 VDD.n48 VDD.n47 0.152939
R14528 VDD.n56 VDD.n48 0.152939
R14529 VDD.n57 VDD.n56 0.152939
R14530 VDD.n58 VDD.n57 0.152939
R14531 VDD.n59 VDD.n58 0.152939
R14532 VDD.n67 VDD.n59 0.152939
R14533 VDD.n68 VDD.n67 0.152939
R14534 VDD.n69 VDD.n68 0.152939
R14535 VDD.n70 VDD.n69 0.152939
R14536 VDD.n78 VDD.n70 0.152939
R14537 VDD.n79 VDD.n78 0.152939
R14538 VDD.n80 VDD.n79 0.152939
R14539 VDD.n81 VDD.n80 0.152939
R14540 VDD.n89 VDD.n81 0.152939
R14541 VDD.n2339 VDD.n89 0.152939
R14542 VDD.n2338 VDD.n90 0.152939
R14543 VDD.n92 VDD.n90 0.152939
R14544 VDD.n96 VDD.n92 0.152939
R14545 VDD.n97 VDD.n96 0.152939
R14546 VDD.n98 VDD.n97 0.152939
R14547 VDD.n99 VDD.n98 0.152939
R14548 VDD.n103 VDD.n99 0.152939
R14549 VDD.n104 VDD.n103 0.152939
R14550 VDD.n105 VDD.n104 0.152939
R14551 VDD.n106 VDD.n105 0.152939
R14552 VDD.n110 VDD.n106 0.152939
R14553 VDD.n111 VDD.n110 0.152939
R14554 VDD.n112 VDD.n111 0.152939
R14555 VDD.n113 VDD.n112 0.152939
R14556 VDD.n117 VDD.n113 0.152939
R14557 VDD.n118 VDD.n117 0.152939
R14558 VDD.n119 VDD.n118 0.152939
R14559 VDD.n120 VDD.n119 0.152939
R14560 VDD.n124 VDD.n120 0.152939
R14561 VDD.n125 VDD.n124 0.152939
R14562 VDD.n126 VDD.n125 0.152939
R14563 VDD.n127 VDD.n126 0.152939
R14564 VDD.n131 VDD.n127 0.152939
R14565 VDD.n132 VDD.n131 0.152939
R14566 VDD.n133 VDD.n132 0.152939
R14567 VDD.n134 VDD.n133 0.152939
R14568 VDD.n138 VDD.n134 0.152939
R14569 VDD.n139 VDD.n138 0.152939
R14570 VDD.n140 VDD.n139 0.152939
R14571 VDD.n141 VDD.n140 0.152939
R14572 VDD.n145 VDD.n141 0.152939
R14573 VDD.n146 VDD.n145 0.152939
R14574 VDD.n147 VDD.n146 0.152939
R14575 VDD.n148 VDD.n147 0.152939
R14576 VDD.n152 VDD.n148 0.152939
R14577 VDD.n153 VDD.n152 0.152939
R14578 VDD.n154 VDD.n153 0.152939
R14579 VDD.n155 VDD.n154 0.152939
R14580 VDD.n159 VDD.n155 0.152939
R14581 VDD.n160 VDD.n159 0.152939
R14582 VDD.n161 VDD.n160 0.152939
R14583 VDD.n162 VDD.n161 0.152939
R14584 VDD.n166 VDD.n162 0.152939
R14585 VDD.n167 VDD.n166 0.152939
R14586 VDD.n2249 VDD.n167 0.152939
R14587 VDD.n2249 VDD.n2248 0.152939
R14588 VDD.n2153 VDD.n236 0.152939
R14589 VDD.n2154 VDD.n2153 0.152939
R14590 VDD.n2155 VDD.n2154 0.152939
R14591 VDD.n2155 VDD.n225 0.152939
R14592 VDD.n2169 VDD.n225 0.152939
R14593 VDD.n2170 VDD.n2169 0.152939
R14594 VDD.n2171 VDD.n2170 0.152939
R14595 VDD.n2171 VDD.n213 0.152939
R14596 VDD.n2185 VDD.n213 0.152939
R14597 VDD.n2186 VDD.n2185 0.152939
R14598 VDD.n2187 VDD.n2186 0.152939
R14599 VDD.n2187 VDD.n201 0.152939
R14600 VDD.n2201 VDD.n201 0.152939
R14601 VDD.n2202 VDD.n2201 0.152939
R14602 VDD.n2203 VDD.n2202 0.152939
R14603 VDD.n2203 VDD.n187 0.152939
R14604 VDD.n2217 VDD.n187 0.152939
R14605 VDD.n2218 VDD.n2217 0.152939
R14606 VDD.n2219 VDD.n2218 0.152939
R14607 VDD.n2219 VDD.n185 0.152939
R14608 VDD.n2223 VDD.n185 0.152939
R14609 VDD.n2224 VDD.n2223 0.152939
R14610 VDD.n2225 VDD.n2224 0.152939
R14611 VDD.n2225 VDD.n182 0.152939
R14612 VDD.n2229 VDD.n182 0.152939
R14613 VDD.n2230 VDD.n2229 0.152939
R14614 VDD.n2231 VDD.n2230 0.152939
R14615 VDD.n2231 VDD.n179 0.152939
R14616 VDD.n2235 VDD.n179 0.152939
R14617 VDD.n2236 VDD.n2235 0.152939
R14618 VDD.n2237 VDD.n2236 0.152939
R14619 VDD.n2237 VDD.n176 0.152939
R14620 VDD.n2241 VDD.n176 0.152939
R14621 VDD.n2242 VDD.n2241 0.152939
R14622 VDD.n2243 VDD.n2242 0.152939
R14623 VDD.n2243 VDD.n173 0.152939
R14624 VDD.n2247 VDD.n173 0.152939
R14625 VDD.n2040 VDD.n305 0.152939
R14626 VDD.n2044 VDD.n2040 0.152939
R14627 VDD.n2044 VDD.n2043 0.152939
R14628 VDD.n1328 VDD.n593 0.152939
R14629 VDD.n600 VDD.n593 0.152939
R14630 VDD.n1052 VDD.n600 0.152939
R14631 VDD.n921 VDD.n731 0.152939
R14632 VDD.n922 VDD.n921 0.152939
R14633 VDD.n923 VDD.n922 0.152939
R14634 VDD.n923 VDD.n720 0.152939
R14635 VDD.n937 VDD.n720 0.152939
R14636 VDD.n938 VDD.n937 0.152939
R14637 VDD.n939 VDD.n938 0.152939
R14638 VDD.n939 VDD.n708 0.152939
R14639 VDD.n953 VDD.n708 0.152939
R14640 VDD.n954 VDD.n953 0.152939
R14641 VDD.n955 VDD.n954 0.152939
R14642 VDD.n955 VDD.n696 0.152939
R14643 VDD.n969 VDD.n696 0.152939
R14644 VDD.n970 VDD.n969 0.152939
R14645 VDD.n971 VDD.n970 0.152939
R14646 VDD.n971 VDD.n683 0.152939
R14647 VDD.n986 VDD.n683 0.152939
R14648 VDD.n987 VDD.n986 0.152939
R14649 VDD.n988 VDD.n987 0.152939
R14650 VDD.n988 VDD.n652 0.152939
R14651 VDD.n1002 VDD.n652 0.152939
R14652 VDD.n1003 VDD.n1002 0.152939
R14653 VDD.n1004 VDD.n1003 0.152939
R14654 VDD.n1004 VDD.n640 0.152939
R14655 VDD.n1018 VDD.n640 0.152939
R14656 VDD.n1019 VDD.n1018 0.152939
R14657 VDD.n1020 VDD.n1019 0.152939
R14658 VDD.n1020 VDD.n628 0.152939
R14659 VDD.n1034 VDD.n628 0.152939
R14660 VDD.n1035 VDD.n1034 0.152939
R14661 VDD.n1036 VDD.n1035 0.152939
R14662 VDD.n1036 VDD.n615 0.152939
R14663 VDD.n1050 VDD.n615 0.152939
R14664 VDD.n1051 VDD.n1050 0.152939
R14665 VDD.n1055 VDD.n1051 0.152939
R14666 VDD.n1055 VDD.n1054 0.152939
R14667 VDD.n1054 VDD.n1053 0.152939
R14668 VDD.n913 VDD.n738 0.152939
R14669 VDD.n906 VDD.n738 0.152939
R14670 VDD.n906 VDD.n905 0.152939
R14671 VDD.n905 VDD.n904 0.152939
R14672 VDD.n904 VDD.n765 0.152939
R14673 VDD.n900 VDD.n765 0.152939
R14674 VDD.n900 VDD.n899 0.152939
R14675 VDD.n899 VDD.n898 0.152939
R14676 VDD.n898 VDD.n771 0.152939
R14677 VDD.n891 VDD.n771 0.152939
R14678 VDD.n891 VDD.n890 0.152939
R14679 VDD.n890 VDD.n889 0.152939
R14680 VDD.n889 VDD.n777 0.152939
R14681 VDD.n885 VDD.n777 0.152939
R14682 VDD.n885 VDD.n884 0.152939
R14683 VDD.n884 VDD.n883 0.152939
R14684 VDD.n883 VDD.n783 0.152939
R14685 VDD.n879 VDD.n783 0.152939
R14686 VDD.n879 VDD.n878 0.152939
R14687 VDD.n878 VDD.n877 0.152939
R14688 VDD.n877 VDD.n789 0.152939
R14689 VDD.n870 VDD.n789 0.152939
R14690 VDD.n870 VDD.n869 0.152939
R14691 VDD.n869 VDD.n868 0.152939
R14692 VDD.n868 VDD.n795 0.152939
R14693 VDD.n864 VDD.n795 0.152939
R14694 VDD.n864 VDD.n863 0.152939
R14695 VDD.n863 VDD.n862 0.152939
R14696 VDD.n862 VDD.n801 0.152939
R14697 VDD.n858 VDD.n801 0.152939
R14698 VDD.n858 VDD.n857 0.152939
R14699 VDD.n857 VDD.n856 0.152939
R14700 VDD.n856 VDD.n807 0.152939
R14701 VDD.n849 VDD.n807 0.152939
R14702 VDD.n849 VDD.n848 0.152939
R14703 VDD.n848 VDD.n847 0.152939
R14704 VDD.n847 VDD.n813 0.152939
R14705 VDD.n843 VDD.n813 0.152939
R14706 VDD.n843 VDD.n842 0.152939
R14707 VDD.n842 VDD.n841 0.152939
R14708 VDD.n841 VDD.n819 0.152939
R14709 VDD.n837 VDD.n819 0.152939
R14710 VDD.n837 VDD.n836 0.152939
R14711 VDD.n836 VDD.n835 0.152939
R14712 VDD.n835 VDD.n825 0.152939
R14713 VDD.n828 VDD.n825 0.152939
R14714 VDD.n915 VDD.n914 0.152939
R14715 VDD.n915 VDD.n726 0.152939
R14716 VDD.n929 VDD.n726 0.152939
R14717 VDD.n930 VDD.n929 0.152939
R14718 VDD.n931 VDD.n930 0.152939
R14719 VDD.n931 VDD.n714 0.152939
R14720 VDD.n945 VDD.n714 0.152939
R14721 VDD.n946 VDD.n945 0.152939
R14722 VDD.n947 VDD.n946 0.152939
R14723 VDD.n947 VDD.n702 0.152939
R14724 VDD.n961 VDD.n702 0.152939
R14725 VDD.n962 VDD.n961 0.152939
R14726 VDD.n963 VDD.n962 0.152939
R14727 VDD.n963 VDD.n690 0.152939
R14728 VDD.n977 VDD.n690 0.152939
R14729 VDD.n978 VDD.n977 0.152939
R14730 VDD.n980 VDD.n978 0.152939
R14731 VDD.n980 VDD.n979 0.152939
R14732 VDD.n1305 VDD.n1304 0.0828171
R14733 VDD.n1988 VDD.n270 0.0828171
R14734 VDD.n2055 VDD.n305 0.0828171
R14735 VDD.n1329 VDD.n1328 0.0828171
R14736 VDD.n1305 VDD.n1068 0.070622
R14737 VDD.n1329 VDD.n590 0.070622
R14738 VDD.n1988 VDD.n273 0.070622
R14739 VDD.n2055 VDD.n303 0.070622
R14740 VDD.n994 VDD.n678 0.0695946
R14741 VDD.n2380 VDD.n35 0.0695946
R14742 VDD.n2380 VDD.n2379 0.0695946
R14743 VDD.n979 VDD.n678 0.0695946
R14744 VDD VDD.n15 0.00833333
R14745 VOUT.n48 VOUT.t10 129.287
R14746 VOUT.n43 VOUT.t24 129.287
R14747 VOUT.n38 VOUT.t27 129.287
R14748 VOUT.n34 VOUT.t16 129.287
R14749 VOUT.n17 VOUT.t33 127.27
R14750 VOUT.n12 VOUT.t5 127.27
R14751 VOUT.n7 VOUT.t43 127.27
R14752 VOUT.n3 VOUT.t34 127.27
R14753 VOUT.n16 VOUT.n14 120.549
R14754 VOUT.n11 VOUT.n9 120.549
R14755 VOUT.n6 VOUT.n4 120.549
R14756 VOUT.n2 VOUT.n0 120.549
R14757 VOUT.n50 VOUT.n49 118.532
R14758 VOUT.n48 VOUT.n47 118.532
R14759 VOUT.n45 VOUT.n44 118.532
R14760 VOUT.n43 VOUT.n42 118.532
R14761 VOUT.n40 VOUT.n39 118.532
R14762 VOUT.n38 VOUT.n37 118.532
R14763 VOUT.n36 VOUT.n35 118.532
R14764 VOUT.n34 VOUT.n33 118.532
R14765 VOUT.n16 VOUT.n15 118.532
R14766 VOUT.n11 VOUT.n10 118.532
R14767 VOUT.n6 VOUT.n5 118.532
R14768 VOUT.n2 VOUT.n1 118.532
R14769 VOUT.n55 VOUT.n53 98.3467
R14770 VOUT.n59 VOUT.n57 98.3467
R14771 VOUT.n55 VOUT.n54 96.3122
R14772 VOUT.n59 VOUT.n58 96.3122
R14773 VOUT.n56 VOUT.n55 10.0764
R14774 VOUT.n60 VOUT.n59 10.0764
R14775 VOUT.n41 VOUT.n36 8.93153
R14776 VOUT.n56 VOUT.n52 8.81804
R14777 VOUT.n49 VOUT.t36 8.7384
R14778 VOUT.n49 VOUT.t40 8.7384
R14779 VOUT.n47 VOUT.t19 8.7384
R14780 VOUT.n47 VOUT.t28 8.7384
R14781 VOUT.n44 VOUT.t8 8.7384
R14782 VOUT.n44 VOUT.t15 8.7384
R14783 VOUT.n42 VOUT.t35 8.7384
R14784 VOUT.n42 VOUT.t42 8.7384
R14785 VOUT.n39 VOUT.t32 8.7384
R14786 VOUT.n39 VOUT.t41 8.7384
R14787 VOUT.n37 VOUT.t21 8.7384
R14788 VOUT.n37 VOUT.t38 8.7384
R14789 VOUT.n35 VOUT.t20 8.7384
R14790 VOUT.n35 VOUT.t29 8.7384
R14791 VOUT.n33 VOUT.t9 8.7384
R14792 VOUT.n33 VOUT.t26 8.7384
R14793 VOUT.n14 VOUT.t37 8.7384
R14794 VOUT.n14 VOUT.t31 8.7384
R14795 VOUT.n15 VOUT.t13 8.7384
R14796 VOUT.n15 VOUT.t7 8.7384
R14797 VOUT.n9 VOUT.t14 8.7384
R14798 VOUT.n9 VOUT.t44 8.7384
R14799 VOUT.n10 VOUT.t25 8.7384
R14800 VOUT.n10 VOUT.t23 8.7384
R14801 VOUT.n4 VOUT.t12 8.7384
R14802 VOUT.n4 VOUT.t17 8.7384
R14803 VOUT.n5 VOUT.t22 8.7384
R14804 VOUT.n5 VOUT.t30 8.7384
R14805 VOUT.n0 VOUT.t39 8.7384
R14806 VOUT.n0 VOUT.t6 8.7384
R14807 VOUT.n1 VOUT.t11 8.7384
R14808 VOUT.n1 VOUT.t18 8.7384
R14809 VOUT.n8 VOUT.n3 7.92291
R14810 VOUT.n54 VOUT.t2 7.64529
R14811 VOUT.n54 VOUT.t47 7.64529
R14812 VOUT.n53 VOUT.t46 7.64529
R14813 VOUT.n53 VOUT.t4 7.64529
R14814 VOUT.n58 VOUT.t45 7.64529
R14815 VOUT.n58 VOUT.t0 7.64529
R14816 VOUT.n57 VOUT.t3 7.64529
R14817 VOUT.n57 VOUT.t1 7.64529
R14818 VOUT.n51 VOUT.n50 6.40998
R14819 VOUT.n46 VOUT.n45 6.40998
R14820 VOUT.n41 VOUT.n40 6.40998
R14821 VOUT.n52 VOUT.n51 6.17128
R14822 VOUT.n19 VOUT.n18 6.17128
R14823 VOUT.n18 VOUT.n17 5.40136
R14824 VOUT.n13 VOUT.n12 5.40136
R14825 VOUT.n8 VOUT.n7 5.40136
R14826 VOUT.n61 VOUT.n19 4.61632
R14827 VOUT.n61 VOUT.n60 4.18271
R14828 VOUT.n52 VOUT.n19 3.4409
R14829 VOUT.n32 VOUT 2.9333
R14830 VOUT.n46 VOUT.n41 2.52636
R14831 VOUT.n13 VOUT.n8 2.52636
R14832 VOUT.n51 VOUT.n46 2.52205
R14833 VOUT.n18 VOUT.n13 2.52205
R14834 VOUT.n60 VOUT.n56 2.27937
R14835 VOUT.n50 VOUT.n48 2.01774
R14836 VOUT.n45 VOUT.n43 2.01774
R14837 VOUT.n40 VOUT.n38 2.01774
R14838 VOUT.n36 VOUT.n34 2.01774
R14839 VOUT.n17 VOUT.n16 2.01774
R14840 VOUT.n12 VOUT.n11 2.01774
R14841 VOUT.n7 VOUT.n6 2.01774
R14842 VOUT.n3 VOUT.n2 2.01774
R14843 VOUT.n32 VOUT.n31 0.335243
R14844 VOUT.n61 VOUT.n32 0.28438
R14845 VOUT.n23 VOUT.t50 0.221979
R14846 VOUT.n29 VOUT.t53 0.221979
R14847 VOUT.n31 VOUT.t49 0.221979
R14848 VOUT.n25 VOUT.t50 0.175863
R14849 VOUT.t53 VOUT.n28 0.175863
R14850 VOUT.t49 VOUT.n30 0.175863
R14851 VOUT.n26 VOUT.t51 0.099351
R14852 VOUT.n27 VOUT.t52 0.0991714
R14853 VOUT.n22 VOUT.t48 0.098698
R14854 VOUT.n26 VOUT.n25 0.0952941
R14855 VOUT.n28 VOUT.n27 0.0936984
R14856 VOUT.n23 VOUT.n22 0.0910262
R14857 VOUT.n30 VOUT.n29 0.0844497
R14858 VOUT.n27 VOUT.n26 0.0619976
R14859 VOUT.n22 VOUT.n20 0.0479372
R14860 VOUT.n24 VOUT.n21 0.0391444
R14861 VOUT.n24 VOUT.n23 0.0193427
R14862 VOUT.n29 VOUT.n21 0.0193427
R14863 VOUT.n31 VOUT.n20 0.0193427
R14864 VOUT.n25 VOUT.n24 0.015385
R14865 VOUT.n28 VOUT.n21 0.015385
R14866 VOUT.n30 VOUT.n20 0.015385
R14867 VOUT VOUT.n61 0.0099
R14868 CS_BIAS.n9 CS_BIAS.n8 161.3
R14869 CS_BIAS.n10 CS_BIAS.n2 161.3
R14870 CS_BIAS.n12 CS_BIAS.n11 161.3
R14871 CS_BIAS.n13 CS_BIAS.n1 161.3
R14872 CS_BIAS.n15 CS_BIAS.n14 161.3
R14873 CS_BIAS.n34 CS_BIAS.n33 161.3
R14874 CS_BIAS.n32 CS_BIAS.n20 161.3
R14875 CS_BIAS.n31 CS_BIAS.n30 161.3
R14876 CS_BIAS.n29 CS_BIAS.n21 161.3
R14877 CS_BIAS.n28 CS_BIAS.n27 161.3
R14878 CS_BIAS.n8 CS_BIAS.n7 99.6671
R14879 CS_BIAS.n27 CS_BIAS.n26 99.667
R14880 CS_BIAS.n5 CS_BIAS.n4 88.6441
R14881 CS_BIAS.n24 CS_BIAS.n22 88.6441
R14882 CS_BIAS.n16 CS_BIAS.n0 60.223
R14883 CS_BIAS.n35 CS_BIAS.n19 60.223
R14884 CS_BIAS.n17 CS_BIAS.t8 46.3887
R14885 CS_BIAS.n36 CS_BIAS.t14 46.3887
R14886 CS_BIAS.n23 CS_BIAS.t0 46.3887
R14887 CS_BIAS.n3 CS_BIAS.t6 46.3885
R14888 CS_BIAS.n17 CS_BIAS.t12 44.527
R14889 CS_BIAS.n3 CS_BIAS.t2 44.527
R14890 CS_BIAS.n36 CS_BIAS.t10 44.527
R14891 CS_BIAS.n23 CS_BIAS.t4 44.527
R14892 CS_BIAS.n26 CS_BIAS.t13 37.5179
R14893 CS_BIAS.n7 CS_BIAS.t15 37.5178
R14894 CS_BIAS.n14 CS_BIAS.n13 24.4675
R14895 CS_BIAS.n13 CS_BIAS.n12 24.4675
R14896 CS_BIAS.n12 CS_BIAS.n2 24.4675
R14897 CS_BIAS.n8 CS_BIAS.n2 24.4675
R14898 CS_BIAS.n27 CS_BIAS.n21 24.4675
R14899 CS_BIAS.n31 CS_BIAS.n21 24.4675
R14900 CS_BIAS.n32 CS_BIAS.n31 24.4675
R14901 CS_BIAS.n33 CS_BIAS.n32 24.4675
R14902 CS_BIAS.n14 CS_BIAS.n0 18.5954
R14903 CS_BIAS.n33 CS_BIAS.n19 18.5954
R14904 CS_BIAS.n24 CS_BIAS.n23 14.8586
R14905 CS_BIAS.n5 CS_BIAS.n3 14.8586
R14906 CS_BIAS.n0 CS_BIAS.t11 12.6616
R14907 CS_BIAS.n19 CS_BIAS.t9 12.6616
R14908 CS_BIAS.n38 CS_BIAS.n18 11.4116
R14909 CS_BIAS.n38 CS_BIAS.n37 9.89345
R14910 CS_BIAS.n6 CS_BIAS.n5 9.503
R14911 CS_BIAS.n25 CS_BIAS.n24 9.503
R14912 CS_BIAS.n26 CS_BIAS.n25 8.9142
R14913 CS_BIAS.n7 CS_BIAS.n6 8.91415
R14914 CS_BIAS.n4 CS_BIAS.t3 7.64529
R14915 CS_BIAS.n4 CS_BIAS.t7 7.64529
R14916 CS_BIAS.n22 CS_BIAS.t1 7.64529
R14917 CS_BIAS.n22 CS_BIAS.t5 7.64529
R14918 CS_BIAS.n18 CS_BIAS.n16 7.20766
R14919 CS_BIAS.n37 CS_BIAS.n35 7.20766
R14920 CS_BIAS.n18 CS_BIAS.n17 6.23401
R14921 CS_BIAS.n37 CS_BIAS.n36 6.23401
R14922 CS_BIAS CS_BIAS.n38 4.18569
R14923 CS_BIAS.n16 CS_BIAS.n15 0.466196
R14924 CS_BIAS.n35 CS_BIAS.n34 0.466196
R14925 CS_BIAS.n15 CS_BIAS.n1 0.189894
R14926 CS_BIAS.n11 CS_BIAS.n1 0.189894
R14927 CS_BIAS.n11 CS_BIAS.n10 0.189894
R14928 CS_BIAS.n10 CS_BIAS.n9 0.189894
R14929 CS_BIAS.n29 CS_BIAS.n28 0.189894
R14930 CS_BIAS.n30 CS_BIAS.n29 0.189894
R14931 CS_BIAS.n30 CS_BIAS.n20 0.189894
R14932 CS_BIAS.n34 CS_BIAS.n20 0.189894
R14933 CS_BIAS.n9 CS_BIAS.n6 0.0762576
R14934 CS_BIAS.n28 CS_BIAS.n25 0.0762576
R14935 a_n2040_7754.n2 a_n2040_7754.t10 127.13
R14936 a_n2040_7754.n1 a_n2040_7754.t9 107.555
R14937 a_n2040_7754.n7 a_n2040_7754.t6 94.4351
R14938 a_n2040_7754.n0 a_n2040_7754.t3 91.8144
R14939 a_n2040_7754.n3 a_n2040_7754.t7 91.8144
R14940 a_n2040_7754.t8 a_n2040_7754.n0 91.8144
R14941 a_n2040_7754.n7 a_n2040_7754.n6 85.3135
R14942 a_n2040_7754.n5 a_n2040_7754.n4 85.3135
R14943 a_n2040_7754.n1 a_n2040_7754.t0 9.01154
R14944 a_n2040_7754.n3 a_n2040_7754.n2 6.78929
R14945 a_n2040_7754.n6 a_n2040_7754.t4 6.5015
R14946 a_n2040_7754.n6 a_n2040_7754.t1 6.5015
R14947 a_n2040_7754.n4 a_n2040_7754.t5 6.5015
R14948 a_n2040_7754.n4 a_n2040_7754.t2 6.5015
R14949 a_n2040_7754.n0 a_n2040_7754.n5 3.29576
R14950 a_n2040_7754.n2 a_n2040_7754.n1 3.2808
R14951 a_n2040_7754.n5 a_n2040_7754.n3 2.62119
R14952 a_n2040_7754.n0 a_n2040_7754.n7 2.62119
R14953 a_n5586_9514.n3 a_n5586_9514.t8 133.567
R14954 a_n5586_9514.n3 a_n5586_9514.t9 127.624
R14955 a_n5586_9514.n2 a_n5586_9514.t3 94.4351
R14956 a_n5586_9514.n4 a_n5586_9514.t1 91.8144
R14957 a_n5586_9514.n0 a_n5586_9514.t4 91.8144
R14958 a_n5586_9514.t7 a_n5586_9514.n0 91.8144
R14959 a_n5586_9514.n6 a_n5586_9514.n5 85.3135
R14960 a_n5586_9514.n2 a_n5586_9514.n1 85.3135
R14961 a_n5586_9514.n4 a_n5586_9514.n3 6.78929
R14962 a_n5586_9514.n5 a_n5586_9514.t2 6.5015
R14963 a_n5586_9514.n5 a_n5586_9514.t0 6.5015
R14964 a_n5586_9514.n1 a_n5586_9514.t6 6.5015
R14965 a_n5586_9514.n1 a_n5586_9514.t5 6.5015
R14966 a_n5586_9514.n0 a_n5586_9514.n2 3.29576
R14967 a_n5586_9514.n0 a_n5586_9514.n6 2.62119
R14968 a_n5586_9514.n6 a_n5586_9514.n4 2.62119
R14969 VP.n30 VP.t1 243.255
R14970 VP.n30 VP.n29 224.169
R14971 VP.n19 VP.n16 161.3
R14972 VP.n21 VP.n20 161.3
R14973 VP.n22 VP.n15 161.3
R14974 VP.n24 VP.n23 161.3
R14975 VP.n25 VP.n14 161.3
R14976 VP.n11 VP.n0 161.3
R14977 VP.n10 VP.n9 161.3
R14978 VP.n8 VP.n1 161.3
R14979 VP.n7 VP.n6 161.3
R14980 VP.n5 VP.n2 161.3
R14981 VP.n17 VP.t7 98.5691
R14982 VP.n3 VP.t8 98.5691
R14983 VP.n27 VP.n26 97.5443
R14984 VP.n13 VP.n12 97.5443
R14985 VP.n18 VP.t3 63.905
R14986 VP.n26 VP.t4 63.905
R14987 VP.n4 VP.t5 63.905
R14988 VP.n12 VP.t6 63.905
R14989 VP.n20 VP.n15 51.663
R14990 VP.n6 VP.n1 51.663
R14991 VP.n18 VP.n17 48.034
R14992 VP.n4 VP.n3 48.034
R14993 VP.n28 VP.n27 31.9754
R14994 VP.n24 VP.n15 29.3238
R14995 VP.n10 VP.n1 29.3238
R14996 VP.n25 VP.n24 24.4675
R14997 VP.n20 VP.n19 24.4675
R14998 VP.n19 VP.n18 24.4675
R14999 VP.n5 VP.n4 24.4675
R15000 VP.n6 VP.n5 24.4675
R15001 VP.n11 VP.n10 24.4675
R15002 VP.n29 VP.t0 19.8005
R15003 VP.n29 VP.t2 19.8005
R15004 VP.n26 VP.n25 13.2127
R15005 VP.n12 VP.n11 13.2127
R15006 VP.n28 VP.n13 12.4224
R15007 VP VP.n31 11.9627
R15008 VP.n17 VP.n16 6.62503
R15009 VP.n3 VP.n2 6.62503
R15010 VP.n31 VP.n30 4.80222
R15011 VP.n31 VP.n28 0.972091
R15012 VP.n27 VP.n14 0.278367
R15013 VP.n13 VP.n0 0.278367
R15014 VP.n23 VP.n14 0.189894
R15015 VP.n23 VP.n22 0.189894
R15016 VP.n22 VP.n21 0.189894
R15017 VP.n21 VP.n16 0.189894
R15018 VP.n7 VP.n2 0.189894
R15019 VP.n8 VP.n7 0.189894
R15020 VP.n9 VP.n8 0.189894
R15021 VP.n9 VP.n0 0.189894
R15022 a_n1816_n673.n0 a_n1816_n673.n1 7.60658
R15023 a_n1816_n673.n2 a_n1816_n673.n3 7.60658
R15024 a_n1816_n673.n90 a_n1816_n673.n74 289.615
R15025 a_n1816_n673.n69 a_n1816_n673.n53 289.615
R15026 a_n1816_n673.n48 a_n1816_n673.n32 289.615
R15027 a_n1816_n673.n13 a_n1816_n673.n14 7.60658
R15028 a_n1816_n673.n15 a_n1816_n673.n16 7.60658
R15029 a_n1816_n673.n147 a_n1816_n673.n146 185
R15030 a_n1816_n673.n165 a_n1816_n673.n164 185
R15031 a_n1816_n673.n163 a_n1816_n673.n162 185
R15032 a_n1816_n673.n150 a_n1816_n673.n149 185
R15033 a_n1816_n673.n159 a_n1816_n673.n158 185
R15034 a_n1816_n673.n157 a_n1816_n673.n156 185
R15035 a_n1816_n673.n153 a_n1816_n673.n152 185
R15036 a_n1816_n673.n172 a_n1816_n673.n171 185
R15037 a_n1816_n673.n190 a_n1816_n673.n189 185
R15038 a_n1816_n673.n188 a_n1816_n673.n187 185
R15039 a_n1816_n673.n175 a_n1816_n673.n174 185
R15040 a_n1816_n673.n184 a_n1816_n673.n183 185
R15041 a_n1816_n673.n182 a_n1816_n673.n181 185
R15042 a_n1816_n673.n178 a_n1816_n673.n177 185
R15043 a_n1816_n673.n91 a_n1816_n673.n90 185
R15044 a_n1816_n673.n89 a_n1816_n673.n88 185
R15045 a_n1816_n673.n77 a_n1816_n673.n76 185
R15046 a_n1816_n673.n85 a_n1816_n673.n84 185
R15047 a_n1816_n673.n83 a_n1816_n673.n82 185
R15048 a_n1816_n673.n5 a_n1816_n673.n79 185
R15049 a_n1816_n673.n6 a_n1816_n673.n80 185
R15050 a_n1816_n673.n70 a_n1816_n673.n69 185
R15051 a_n1816_n673.n68 a_n1816_n673.n67 185
R15052 a_n1816_n673.n56 a_n1816_n673.n55 185
R15053 a_n1816_n673.n64 a_n1816_n673.n63 185
R15054 a_n1816_n673.n62 a_n1816_n673.n61 185
R15055 a_n1816_n673.n8 a_n1816_n673.n58 185
R15056 a_n1816_n673.n9 a_n1816_n673.n59 185
R15057 a_n1816_n673.n49 a_n1816_n673.n48 185
R15058 a_n1816_n673.n47 a_n1816_n673.n46 185
R15059 a_n1816_n673.n35 a_n1816_n673.n34 185
R15060 a_n1816_n673.n43 a_n1816_n673.n42 185
R15061 a_n1816_n673.n41 a_n1816_n673.n40 185
R15062 a_n1816_n673.n11 a_n1816_n673.n37 185
R15063 a_n1816_n673.n12 a_n1816_n673.n38 185
R15064 a_n1816_n673.n129 a_n1816_n673.n128 185
R15065 a_n1816_n673.n133 a_n1816_n673.n132 185
R15066 a_n1816_n673.n135 a_n1816_n673.n134 185
R15067 a_n1816_n673.n126 a_n1816_n673.n125 185
R15068 a_n1816_n673.n139 a_n1816_n673.n138 185
R15069 a_n1816_n673.n141 a_n1816_n673.n140 185
R15070 a_n1816_n673.n123 a_n1816_n673.n122 185
R15071 a_n1816_n673.n104 a_n1816_n673.n103 185
R15072 a_n1816_n673.n108 a_n1816_n673.n107 185
R15073 a_n1816_n673.n110 a_n1816_n673.n109 185
R15074 a_n1816_n673.n101 a_n1816_n673.n100 185
R15075 a_n1816_n673.n114 a_n1816_n673.n113 185
R15076 a_n1816_n673.n116 a_n1816_n673.n115 185
R15077 a_n1816_n673.n98 a_n1816_n673.n97 185
R15078 a_n1816_n673.n179 a_n1816_n673.t6 149.525
R15079 a_n1816_n673.n154 a_n1816_n673.t2 149.525
R15080 a_n1816_n673.n130 a_n1816_n673.t7 149.525
R15081 a_n1816_n673.n105 a_n1816_n673.t4 149.525
R15082 a_n1816_n673.n94 a_n1816_n673.n93 136.37
R15083 a_n1816_n673.n73 a_n1816_n673.n72 136.37
R15084 a_n1816_n673.n52 a_n1816_n673.n51 136.37
R15085 a_n1816_n673.n1 a_n1816_n673.n146 214.541
R15086 a_n1816_n673.n164 a_n1816_n673.n146 104.615
R15087 a_n1816_n673.n164 a_n1816_n673.n163 104.615
R15088 a_n1816_n673.n163 a_n1816_n673.n149 104.615
R15089 a_n1816_n673.n158 a_n1816_n673.n149 104.615
R15090 a_n1816_n673.n158 a_n1816_n673.n157 104.615
R15091 a_n1816_n673.n157 a_n1816_n673.n152 104.615
R15092 a_n1816_n673.n3 a_n1816_n673.n171 214.541
R15093 a_n1816_n673.n189 a_n1816_n673.n171 104.615
R15094 a_n1816_n673.n189 a_n1816_n673.n188 104.615
R15095 a_n1816_n673.n188 a_n1816_n673.n174 104.615
R15096 a_n1816_n673.n183 a_n1816_n673.n174 104.615
R15097 a_n1816_n673.n183 a_n1816_n673.n182 104.615
R15098 a_n1816_n673.n182 a_n1816_n673.n177 104.615
R15099 a_n1816_n673.n90 a_n1816_n673.n89 104.615
R15100 a_n1816_n673.n89 a_n1816_n673.n76 104.615
R15101 a_n1816_n673.n84 a_n1816_n673.n76 104.615
R15102 a_n1816_n673.n84 a_n1816_n673.n83 104.615
R15103 a_n1816_n673.n83 a_n1816_n673.n79 104.615
R15104 a_n1816_n673.n80 a_n1816_n673.n79 104.615
R15105 a_n1816_n673.n69 a_n1816_n673.n68 104.615
R15106 a_n1816_n673.n68 a_n1816_n673.n55 104.615
R15107 a_n1816_n673.n63 a_n1816_n673.n55 104.615
R15108 a_n1816_n673.n63 a_n1816_n673.n62 104.615
R15109 a_n1816_n673.n62 a_n1816_n673.n58 104.615
R15110 a_n1816_n673.n59 a_n1816_n673.n58 104.615
R15111 a_n1816_n673.n48 a_n1816_n673.n47 104.615
R15112 a_n1816_n673.n47 a_n1816_n673.n34 104.615
R15113 a_n1816_n673.n42 a_n1816_n673.n34 104.615
R15114 a_n1816_n673.n42 a_n1816_n673.n41 104.615
R15115 a_n1816_n673.n41 a_n1816_n673.n37 104.615
R15116 a_n1816_n673.n38 a_n1816_n673.n37 104.615
R15117 a_n1816_n673.n133 a_n1816_n673.n128 104.615
R15118 a_n1816_n673.n134 a_n1816_n673.n133 104.615
R15119 a_n1816_n673.n134 a_n1816_n673.n125 104.615
R15120 a_n1816_n673.n139 a_n1816_n673.n125 104.615
R15121 a_n1816_n673.n140 a_n1816_n673.n139 104.615
R15122 a_n1816_n673.n140 a_n1816_n673.n122 104.615
R15123 a_n1816_n673.n14 a_n1816_n673.n122 214.541
R15124 a_n1816_n673.n108 a_n1816_n673.n103 104.615
R15125 a_n1816_n673.n109 a_n1816_n673.n108 104.615
R15126 a_n1816_n673.n109 a_n1816_n673.n100 104.615
R15127 a_n1816_n673.n114 a_n1816_n673.n100 104.615
R15128 a_n1816_n673.n115 a_n1816_n673.n114 104.615
R15129 a_n1816_n673.n115 a_n1816_n673.n97 104.615
R15130 a_n1816_n673.n16 a_n1816_n673.n97 214.541
R15131 a_n1816_n673.t2 a_n1816_n673.n152 52.3082
R15132 a_n1816_n673.t6 a_n1816_n673.n177 52.3082
R15133 a_n1816_n673.n80 a_n1816_n673.t3 52.3082
R15134 a_n1816_n673.n59 a_n1816_n673.t11 52.3082
R15135 a_n1816_n673.n38 a_n1816_n673.t0 52.3082
R15136 a_n1816_n673.t7 a_n1816_n673.n128 52.3082
R15137 a_n1816_n673.t4 a_n1816_n673.n103 52.3082
R15138 a_n1816_n673.n170 a_n1816_n673.n169 50.8686
R15139 a_n1816_n673.n195 a_n1816_n673.n194 50.8686
R15140 a_n1816_n673.n121 a_n1816_n673.n120 50.8676
R15141 a_n1816_n673.n96 a_n1816_n673.n95 50.8676
R15142 a_n1816_n673.n168 a_n1816_n673.n0 33.9308
R15143 a_n1816_n673.n193 a_n1816_n673.n2 33.9308
R15144 a_n1816_n673.n144 a_n1816_n673.n13 33.9308
R15145 a_n1816_n673.n119 a_n1816_n673.n15 33.9308
R15146 a_n1816_n673.n6 a_n1816_n673.n4 5.10449
R15147 a_n1816_n673.n9 a_n1816_n673.n7 5.10449
R15148 a_n1816_n673.n12 a_n1816_n673.n10 5.10449
R15149 a_n1816_n673.n194 a_n1816_n673.n31 14.2233
R15150 a_n1816_n673.n168 a_n1816_n673.n145 13.0294
R15151 a_n1816_n673.n167 a_n1816_n673.n1 6.02292
R15152 a_n1816_n673.n192 a_n1816_n673.n3 6.02292
R15153 a_n1816_n673.n6 a_n1816_n673.n5 12.8005
R15154 a_n1816_n673.n9 a_n1816_n673.n8 12.8005
R15155 a_n1816_n673.n12 a_n1816_n673.n11 12.8005
R15156 a_n1816_n673.n167 a_n1816_n673.n147 12.0247
R15157 a_n1816_n673.n192 a_n1816_n673.n172 12.0247
R15158 a_n1816_n673.n82 a_n1816_n673.n81 12.0247
R15159 a_n1816_n673.n61 a_n1816_n673.n60 12.0247
R15160 a_n1816_n673.n40 a_n1816_n673.n39 12.0247
R15161 a_n1816_n673.n143 a_n1816_n673.n123 12.0247
R15162 a_n1816_n673.n118 a_n1816_n673.n98 12.0247
R15163 a_n1816_n673.n166 a_n1816_n673.n165 11.249
R15164 a_n1816_n673.n191 a_n1816_n673.n190 11.249
R15165 a_n1816_n673.n85 a_n1816_n673.n78 11.249
R15166 a_n1816_n673.n64 a_n1816_n673.n57 11.249
R15167 a_n1816_n673.n43 a_n1816_n673.n36 11.249
R15168 a_n1816_n673.n142 a_n1816_n673.n141 11.249
R15169 a_n1816_n673.n117 a_n1816_n673.n116 11.249
R15170 a_n1816_n673.n162 a_n1816_n673.n148 10.4732
R15171 a_n1816_n673.n187 a_n1816_n673.n173 10.4732
R15172 a_n1816_n673.n86 a_n1816_n673.n77 10.4732
R15173 a_n1816_n673.n65 a_n1816_n673.n56 10.4732
R15174 a_n1816_n673.n44 a_n1816_n673.n35 10.4732
R15175 a_n1816_n673.n138 a_n1816_n673.n124 10.4732
R15176 a_n1816_n673.n113 a_n1816_n673.n99 10.4732
R15177 a_n1816_n673.n154 a_n1816_n673.n153 10.2746
R15178 a_n1816_n673.n179 a_n1816_n673.n178 10.2746
R15179 a_n1816_n673.n130 a_n1816_n673.n129 10.2746
R15180 a_n1816_n673.n105 a_n1816_n673.n104 10.2746
R15181 a_n1816_n673.n18 a_n1816_n673.n15 9.84355
R15182 a_n1816_n673.n20 a_n1816_n673.n13 9.84355
R15183 a_n1816_n673.n161 a_n1816_n673.n150 9.69747
R15184 a_n1816_n673.n186 a_n1816_n673.n175 9.69747
R15185 a_n1816_n673.n88 a_n1816_n673.n87 9.69747
R15186 a_n1816_n673.n67 a_n1816_n673.n66 9.69747
R15187 a_n1816_n673.n46 a_n1816_n673.n45 9.69747
R15188 a_n1816_n673.n137 a_n1816_n673.n126 9.69747
R15189 a_n1816_n673.n112 a_n1816_n673.n101 9.69747
R15190 a_n1816_n673.n21 a_n1816_n673.n10 1.42956
R15191 a_n1816_n673.n93 a_n1816_n673.n26 9.45567
R15192 a_n1816_n673.n72 a_n1816_n673.n24 9.45567
R15193 a_n1816_n673.n51 a_n1816_n673.n22 9.45567
R15194 a_n1816_n673.n167 a_n1816_n673.n29 9.3005
R15195 a_n1816_n673.n29 a_n1816_n673.n166 9.3005
R15196 a_n1816_n673.n148 a_n1816_n673.n29 9.3005
R15197 a_n1816_n673.n161 a_n1816_n673.n30 9.3005
R15198 a_n1816_n673.n30 a_n1816_n673.n160 9.3005
R15199 a_n1816_n673.n151 a_n1816_n673.n30 9.3005
R15200 a_n1816_n673.n155 a_n1816_n673.n30 9.3005
R15201 a_n1816_n673.n176 a_n1816_n673.n28 9.3005
R15202 a_n1816_n673.n28 a_n1816_n673.n185 9.3005
R15203 a_n1816_n673.n186 a_n1816_n673.n28 9.3005
R15204 a_n1816_n673.n173 a_n1816_n673.n27 9.3005
R15205 a_n1816_n673.n27 a_n1816_n673.n191 9.3005
R15206 a_n1816_n673.n192 a_n1816_n673.n27 9.3005
R15207 a_n1816_n673.n180 a_n1816_n673.n28 9.3005
R15208 a_n1816_n673.n26 a_n1816_n673.n92 9.3005
R15209 a_n1816_n673.n75 a_n1816_n673.n26 9.3005
R15210 a_n1816_n673.n87 a_n1816_n673.n26 9.3005
R15211 a_n1816_n673.n25 a_n1816_n673.n86 9.3005
R15212 a_n1816_n673.n78 a_n1816_n673.n25 9.3005
R15213 a_n1816_n673.n81 a_n1816_n673.n25 9.3005
R15214 a_n1816_n673.n24 a_n1816_n673.n71 9.3005
R15215 a_n1816_n673.n54 a_n1816_n673.n24 9.3005
R15216 a_n1816_n673.n66 a_n1816_n673.n24 9.3005
R15217 a_n1816_n673.n23 a_n1816_n673.n65 9.3005
R15218 a_n1816_n673.n57 a_n1816_n673.n23 9.3005
R15219 a_n1816_n673.n60 a_n1816_n673.n23 9.3005
R15220 a_n1816_n673.n22 a_n1816_n673.n50 9.3005
R15221 a_n1816_n673.n33 a_n1816_n673.n22 9.3005
R15222 a_n1816_n673.n45 a_n1816_n673.n22 9.3005
R15223 a_n1816_n673.n21 a_n1816_n673.n44 9.3005
R15224 a_n1816_n673.n36 a_n1816_n673.n21 9.3005
R15225 a_n1816_n673.n39 a_n1816_n673.n21 9.3005
R15226 a_n1816_n673.n131 a_n1816_n673.n19 9.3005
R15227 a_n1816_n673.n127 a_n1816_n673.n19 9.3005
R15228 a_n1816_n673.n19 a_n1816_n673.n136 9.3005
R15229 a_n1816_n673.n137 a_n1816_n673.n20 9.3005
R15230 a_n1816_n673.n124 a_n1816_n673.n20 9.3005
R15231 a_n1816_n673.n20 a_n1816_n673.n142 9.3005
R15232 a_n1816_n673.n143 a_n1816_n673.n20 9.3005
R15233 a_n1816_n673.n106 a_n1816_n673.n17 9.3005
R15234 a_n1816_n673.n102 a_n1816_n673.n17 9.3005
R15235 a_n1816_n673.n17 a_n1816_n673.n111 9.3005
R15236 a_n1816_n673.n112 a_n1816_n673.n18 9.3005
R15237 a_n1816_n673.n99 a_n1816_n673.n18 9.3005
R15238 a_n1816_n673.n18 a_n1816_n673.n117 9.3005
R15239 a_n1816_n673.n118 a_n1816_n673.n18 9.3005
R15240 a_n1816_n673.n160 a_n1816_n673.n159 8.92171
R15241 a_n1816_n673.n185 a_n1816_n673.n184 8.92171
R15242 a_n1816_n673.n91 a_n1816_n673.n75 8.92171
R15243 a_n1816_n673.n70 a_n1816_n673.n54 8.92171
R15244 a_n1816_n673.n49 a_n1816_n673.n33 8.92171
R15245 a_n1816_n673.n136 a_n1816_n673.n135 8.92171
R15246 a_n1816_n673.n111 a_n1816_n673.n110 8.92171
R15247 a_n1816_n673.n156 a_n1816_n673.n151 8.14595
R15248 a_n1816_n673.n181 a_n1816_n673.n176 8.14595
R15249 a_n1816_n673.n92 a_n1816_n673.n74 8.14595
R15250 a_n1816_n673.n71 a_n1816_n673.n53 8.14595
R15251 a_n1816_n673.n50 a_n1816_n673.n32 8.14595
R15252 a_n1816_n673.n132 a_n1816_n673.n127 8.14595
R15253 a_n1816_n673.n107 a_n1816_n673.n102 8.14595
R15254 a_n1816_n673.n96 a_n1816_n673.n31 7.65136
R15255 a_n1816_n673.n155 a_n1816_n673.n153 7.3702
R15256 a_n1816_n673.n180 a_n1816_n673.n178 7.3702
R15257 a_n1816_n673.n131 a_n1816_n673.n129 7.3702
R15258 a_n1816_n673.n106 a_n1816_n673.n104 7.3702
R15259 a_n1816_n673.n145 a_n1816_n673.n144 6.4574
R15260 a_n1816_n673.n156 a_n1816_n673.n155 5.81868
R15261 a_n1816_n673.n181 a_n1816_n673.n180 5.81868
R15262 a_n1816_n673.n93 a_n1816_n673.n74 5.81868
R15263 a_n1816_n673.n72 a_n1816_n673.n53 5.81868
R15264 a_n1816_n673.n51 a_n1816_n673.n32 5.81868
R15265 a_n1816_n673.n132 a_n1816_n673.n131 5.81868
R15266 a_n1816_n673.n107 a_n1816_n673.n106 5.81868
R15267 a_n1816_n673.n159 a_n1816_n673.n151 5.04292
R15268 a_n1816_n673.n184 a_n1816_n673.n176 5.04292
R15269 a_n1816_n673.n92 a_n1816_n673.n91 5.04292
R15270 a_n1816_n673.n71 a_n1816_n673.n70 5.04292
R15271 a_n1816_n673.n50 a_n1816_n673.n49 5.04292
R15272 a_n1816_n673.n135 a_n1816_n673.n127 5.04292
R15273 a_n1816_n673.n110 a_n1816_n673.n102 5.04292
R15274 a_n1816_n673.n145 a_n1816_n673.n94 4.43117
R15275 a_n1816_n673.n4 a_n1816_n673.t3 149.972
R15276 a_n1816_n673.n7 a_n1816_n673.t11 149.972
R15277 a_n1816_n673.n10 a_n1816_n673.t0 149.972
R15278 a_n1816_n673.n27 a_n1816_n673.n2 9.84355
R15279 a_n1816_n673.n29 a_n1816_n673.n0 9.84355
R15280 a_n1816_n673.n25 a_n1816_n673.n4 1.42956
R15281 a_n1816_n673.n23 a_n1816_n673.n7 1.42956
R15282 a_n1816_n673.n160 a_n1816_n673.n150 4.26717
R15283 a_n1816_n673.n185 a_n1816_n673.n175 4.26717
R15284 a_n1816_n673.n88 a_n1816_n673.n75 4.26717
R15285 a_n1816_n673.n67 a_n1816_n673.n54 4.26717
R15286 a_n1816_n673.n46 a_n1816_n673.n33 4.26717
R15287 a_n1816_n673.n136 a_n1816_n673.n126 4.26717
R15288 a_n1816_n673.n111 a_n1816_n673.n101 4.26717
R15289 a_n1816_n673.n162 a_n1816_n673.n161 3.49141
R15290 a_n1816_n673.n187 a_n1816_n673.n186 3.49141
R15291 a_n1816_n673.n87 a_n1816_n673.n77 3.49141
R15292 a_n1816_n673.n66 a_n1816_n673.n56 3.49141
R15293 a_n1816_n673.n45 a_n1816_n673.n35 3.49141
R15294 a_n1816_n673.n138 a_n1816_n673.n137 3.49141
R15295 a_n1816_n673.n113 a_n1816_n673.n112 3.49141
R15296 a_n1816_n673.n169 a_n1816_n673.t1 3.06078
R15297 a_n1816_n673.n169 a_n1816_n673.t14 3.06078
R15298 a_n1816_n673.n120 a_n1816_n673.t5 3.06078
R15299 a_n1816_n673.n120 a_n1816_n673.t8 3.06078
R15300 a_n1816_n673.n95 a_n1816_n673.t12 3.06078
R15301 a_n1816_n673.n95 a_n1816_n673.t13 3.06078
R15302 a_n1816_n673.n195 a_n1816_n673.t9 3.06078
R15303 a_n1816_n673.t10 a_n1816_n673.n195 3.06078
R15304 a_n1816_n673.n28 a_n1816_n673.n179 2.84308
R15305 a_n1816_n673.n30 a_n1816_n673.n154 2.84308
R15306 a_n1816_n673.n19 a_n1816_n673.n130 2.84308
R15307 a_n1816_n673.n17 a_n1816_n673.n105 2.84308
R15308 a_n1816_n673.n52 a_n1816_n673.n31 2.78001
R15309 a_n1816_n673.n165 a_n1816_n673.n148 2.71565
R15310 a_n1816_n673.n190 a_n1816_n673.n173 2.71565
R15311 a_n1816_n673.n86 a_n1816_n673.n85 2.71565
R15312 a_n1816_n673.n65 a_n1816_n673.n64 2.71565
R15313 a_n1816_n673.n44 a_n1816_n673.n43 2.71565
R15314 a_n1816_n673.n141 a_n1816_n673.n124 2.71565
R15315 a_n1816_n673.n116 a_n1816_n673.n99 2.71565
R15316 a_n1816_n673.n119 a_n1816_n673.n96 2.38843
R15317 a_n1816_n673.n144 a_n1816_n673.n121 2.38843
R15318 a_n1816_n673.n194 a_n1816_n673.n193 2.38843
R15319 a_n1816_n673.n170 a_n1816_n673.n168 2.38843
R15320 a_n1816_n673.n166 a_n1816_n673.n147 1.93989
R15321 a_n1816_n673.n191 a_n1816_n673.n172 1.93989
R15322 a_n1816_n673.n82 a_n1816_n673.n78 1.93989
R15323 a_n1816_n673.n61 a_n1816_n673.n57 1.93989
R15324 a_n1816_n673.n40 a_n1816_n673.n36 1.93989
R15325 a_n1816_n673.n142 a_n1816_n673.n123 1.93989
R15326 a_n1816_n673.n117 a_n1816_n673.n98 1.93989
R15327 a_n1816_n673.n73 a_n1816_n673.n52 1.93655
R15328 a_n1816_n673.n94 a_n1816_n673.n73 1.93655
R15329 a_n1816_n673.n121 a_n1816_n673.n119 1.66429
R15330 a_n1816_n673.n193 a_n1816_n673.n170 1.66429
R15331 a_n1816_n673.n81 a_n1816_n673.n5 1.16414
R15332 a_n1816_n673.n60 a_n1816_n673.n8 1.16414
R15333 a_n1816_n673.n39 a_n1816_n673.n11 1.16414
R15334 a_n1816_n673.n14 a_n1816_n673.n143 6.02292
R15335 a_n1816_n673.n16 a_n1816_n673.n118 6.02292
R15336 a_n1816_n673.n30 a_n1816_n673.n29 0.931534
R15337 a_n1816_n673.n28 a_n1816_n673.n27 0.931534
R15338 a_n1816_n673.n26 a_n1816_n673.n25 0.931534
R15339 a_n1816_n673.n24 a_n1816_n673.n23 0.931534
R15340 a_n1816_n673.n22 a_n1816_n673.n21 0.931534
R15341 a_n1816_n673.n20 a_n1816_n673.n19 0.931534
R15342 a_n1816_n673.n18 a_n1816_n673.n17 0.931534
R15343 VN.n30 VN.t1 243.97
R15344 VN.n30 VN.n29 223.454
R15345 VN.n25 VN.n14 161.3
R15346 VN.n24 VN.n23 161.3
R15347 VN.n22 VN.n15 161.3
R15348 VN.n21 VN.n20 161.3
R15349 VN.n19 VN.n16 161.3
R15350 VN.n5 VN.n2 161.3
R15351 VN.n7 VN.n6 161.3
R15352 VN.n8 VN.n1 161.3
R15353 VN.n10 VN.n9 161.3
R15354 VN.n11 VN.n0 161.3
R15355 VN.n17 VN.t3 98.5691
R15356 VN.n3 VN.t4 98.5691
R15357 VN.n27 VN.n26 97.5443
R15358 VN.n13 VN.n12 97.5443
R15359 VN.n18 VN.t6 63.905
R15360 VN.n26 VN.t7 63.905
R15361 VN.n4 VN.t5 63.905
R15362 VN.n12 VN.t8 63.905
R15363 VN.n20 VN.n15 51.663
R15364 VN.n6 VN.n1 51.663
R15365 VN.n18 VN.n17 48.034
R15366 VN.n4 VN.n3 48.034
R15367 VN.n28 VN.n27 31.7595
R15368 VN.n24 VN.n15 29.3238
R15369 VN.n10 VN.n1 29.3238
R15370 VN.n19 VN.n18 24.4675
R15371 VN.n20 VN.n19 24.4675
R15372 VN.n25 VN.n24 24.4675
R15373 VN.n11 VN.n10 24.4675
R15374 VN.n6 VN.n5 24.4675
R15375 VN.n5 VN.n4 24.4675
R15376 VN.n29 VN.t2 19.8005
R15377 VN.n29 VN.t0 19.8005
R15378 VN VN.n31 14.8362
R15379 VN.n26 VN.n25 13.2127
R15380 VN.n12 VN.n11 13.2127
R15381 VN.n28 VN.n13 12.2065
R15382 VN.n17 VN.n16 6.62503
R15383 VN.n3 VN.n2 6.62503
R15384 VN.n31 VN.n30 5.40567
R15385 VN.n31 VN.n28 1.188
R15386 VN.n27 VN.n14 0.278367
R15387 VN.n13 VN.n0 0.278367
R15388 VN.n21 VN.n16 0.189894
R15389 VN.n22 VN.n21 0.189894
R15390 VN.n23 VN.n22 0.189894
R15391 VN.n23 VN.n14 0.189894
R15392 VN.n9 VN.n0 0.189894
R15393 VN.n9 VN.n8 0.189894
R15394 VN.n8 VN.n7 0.189894
R15395 VN.n7 VN.n2 0.189894
R15396 DIFFPAIR_BIAS.n26 DIFFPAIR_BIAS.n0 289.615
R15397 DIFFPAIR_BIAS.n57 DIFFPAIR_BIAS.n31 289.615
R15398 DIFFPAIR_BIAS.n89 DIFFPAIR_BIAS.n63 289.615
R15399 DIFFPAIR_BIAS.n27 DIFFPAIR_BIAS.n26 185
R15400 DIFFPAIR_BIAS.n25 DIFFPAIR_BIAS.n24 185
R15401 DIFFPAIR_BIAS.n4 DIFFPAIR_BIAS.n3 185
R15402 DIFFPAIR_BIAS.n19 DIFFPAIR_BIAS.n18 185
R15403 DIFFPAIR_BIAS.n17 DIFFPAIR_BIAS.n16 185
R15404 DIFFPAIR_BIAS.n8 DIFFPAIR_BIAS.n7 185
R15405 DIFFPAIR_BIAS.n11 DIFFPAIR_BIAS.n10 185
R15406 DIFFPAIR_BIAS.n58 DIFFPAIR_BIAS.n57 185
R15407 DIFFPAIR_BIAS.n56 DIFFPAIR_BIAS.n55 185
R15408 DIFFPAIR_BIAS.n35 DIFFPAIR_BIAS.n34 185
R15409 DIFFPAIR_BIAS.n50 DIFFPAIR_BIAS.n49 185
R15410 DIFFPAIR_BIAS.n48 DIFFPAIR_BIAS.n47 185
R15411 DIFFPAIR_BIAS.n39 DIFFPAIR_BIAS.n38 185
R15412 DIFFPAIR_BIAS.n42 DIFFPAIR_BIAS.n41 185
R15413 DIFFPAIR_BIAS.n90 DIFFPAIR_BIAS.n89 185
R15414 DIFFPAIR_BIAS.n88 DIFFPAIR_BIAS.n87 185
R15415 DIFFPAIR_BIAS.n67 DIFFPAIR_BIAS.n66 185
R15416 DIFFPAIR_BIAS.n82 DIFFPAIR_BIAS.n81 185
R15417 DIFFPAIR_BIAS.n80 DIFFPAIR_BIAS.n79 185
R15418 DIFFPAIR_BIAS.n71 DIFFPAIR_BIAS.n70 185
R15419 DIFFPAIR_BIAS.n74 DIFFPAIR_BIAS.n73 185
R15420 DIFFPAIR_BIAS.n100 DIFFPAIR_BIAS.t6 176.166
R15421 DIFFPAIR_BIAS.n99 DIFFPAIR_BIAS.t7 174.857
R15422 DIFFPAIR_BIAS.n98 DIFFPAIR_BIAS.t8 174.857
R15423 DIFFPAIR_BIAS.t3 DIFFPAIR_BIAS.n9 147.661
R15424 DIFFPAIR_BIAS.t1 DIFFPAIR_BIAS.n40 147.661
R15425 DIFFPAIR_BIAS.t5 DIFFPAIR_BIAS.n72 147.661
R15426 DIFFPAIR_BIAS.n95 DIFFPAIR_BIAS.t2 130.703
R15427 DIFFPAIR_BIAS.n95 DIFFPAIR_BIAS.t0 128.767
R15428 DIFFPAIR_BIAS.n96 DIFFPAIR_BIAS.t4 128.767
R15429 DIFFPAIR_BIAS.n26 DIFFPAIR_BIAS.n25 104.615
R15430 DIFFPAIR_BIAS.n25 DIFFPAIR_BIAS.n3 104.615
R15431 DIFFPAIR_BIAS.n18 DIFFPAIR_BIAS.n3 104.615
R15432 DIFFPAIR_BIAS.n18 DIFFPAIR_BIAS.n17 104.615
R15433 DIFFPAIR_BIAS.n17 DIFFPAIR_BIAS.n7 104.615
R15434 DIFFPAIR_BIAS.n10 DIFFPAIR_BIAS.n7 104.615
R15435 DIFFPAIR_BIAS.n57 DIFFPAIR_BIAS.n56 104.615
R15436 DIFFPAIR_BIAS.n56 DIFFPAIR_BIAS.n34 104.615
R15437 DIFFPAIR_BIAS.n49 DIFFPAIR_BIAS.n34 104.615
R15438 DIFFPAIR_BIAS.n49 DIFFPAIR_BIAS.n48 104.615
R15439 DIFFPAIR_BIAS.n48 DIFFPAIR_BIAS.n38 104.615
R15440 DIFFPAIR_BIAS.n41 DIFFPAIR_BIAS.n38 104.615
R15441 DIFFPAIR_BIAS.n89 DIFFPAIR_BIAS.n88 104.615
R15442 DIFFPAIR_BIAS.n88 DIFFPAIR_BIAS.n66 104.615
R15443 DIFFPAIR_BIAS.n81 DIFFPAIR_BIAS.n66 104.615
R15444 DIFFPAIR_BIAS.n81 DIFFPAIR_BIAS.n80 104.615
R15445 DIFFPAIR_BIAS.n80 DIFFPAIR_BIAS.n70 104.615
R15446 DIFFPAIR_BIAS.n73 DIFFPAIR_BIAS.n70 104.615
R15447 DIFFPAIR_BIAS.n62 DIFFPAIR_BIAS.n30 70.0396
R15448 DIFFPAIR_BIAS.n62 DIFFPAIR_BIAS.n61 68.1035
R15449 DIFFPAIR_BIAS.n94 DIFFPAIR_BIAS.n93 68.1035
R15450 DIFFPAIR_BIAS.n10 DIFFPAIR_BIAS.t3 52.3082
R15451 DIFFPAIR_BIAS.n41 DIFFPAIR_BIAS.t1 52.3082
R15452 DIFFPAIR_BIAS.n73 DIFFPAIR_BIAS.t5 52.3082
R15453 DIFFPAIR_BIAS.n11 DIFFPAIR_BIAS.n9 15.6674
R15454 DIFFPAIR_BIAS.n42 DIFFPAIR_BIAS.n40 15.6674
R15455 DIFFPAIR_BIAS.n74 DIFFPAIR_BIAS.n72 15.6674
R15456 DIFFPAIR_BIAS.n12 DIFFPAIR_BIAS.n8 12.8005
R15457 DIFFPAIR_BIAS.n43 DIFFPAIR_BIAS.n39 12.8005
R15458 DIFFPAIR_BIAS.n75 DIFFPAIR_BIAS.n71 12.8005
R15459 DIFFPAIR_BIAS.n16 DIFFPAIR_BIAS.n15 12.0247
R15460 DIFFPAIR_BIAS.n47 DIFFPAIR_BIAS.n46 12.0247
R15461 DIFFPAIR_BIAS.n79 DIFFPAIR_BIAS.n78 12.0247
R15462 DIFFPAIR_BIAS.n19 DIFFPAIR_BIAS.n6 11.249
R15463 DIFFPAIR_BIAS.n50 DIFFPAIR_BIAS.n37 11.249
R15464 DIFFPAIR_BIAS.n82 DIFFPAIR_BIAS.n69 11.249
R15465 DIFFPAIR_BIAS.n20 DIFFPAIR_BIAS.n4 10.4732
R15466 DIFFPAIR_BIAS.n51 DIFFPAIR_BIAS.n35 10.4732
R15467 DIFFPAIR_BIAS.n83 DIFFPAIR_BIAS.n67 10.4732
R15468 DIFFPAIR_BIAS.n24 DIFFPAIR_BIAS.n23 9.69747
R15469 DIFFPAIR_BIAS.n55 DIFFPAIR_BIAS.n54 9.69747
R15470 DIFFPAIR_BIAS.n87 DIFFPAIR_BIAS.n86 9.69747
R15471 DIFFPAIR_BIAS.n30 DIFFPAIR_BIAS.n29 9.45567
R15472 DIFFPAIR_BIAS.n61 DIFFPAIR_BIAS.n60 9.45567
R15473 DIFFPAIR_BIAS.n93 DIFFPAIR_BIAS.n92 9.45567
R15474 DIFFPAIR_BIAS.n29 DIFFPAIR_BIAS.n28 9.3005
R15475 DIFFPAIR_BIAS.n2 DIFFPAIR_BIAS.n1 9.3005
R15476 DIFFPAIR_BIAS.n23 DIFFPAIR_BIAS.n22 9.3005
R15477 DIFFPAIR_BIAS.n21 DIFFPAIR_BIAS.n20 9.3005
R15478 DIFFPAIR_BIAS.n6 DIFFPAIR_BIAS.n5 9.3005
R15479 DIFFPAIR_BIAS.n15 DIFFPAIR_BIAS.n14 9.3005
R15480 DIFFPAIR_BIAS.n13 DIFFPAIR_BIAS.n12 9.3005
R15481 DIFFPAIR_BIAS.n60 DIFFPAIR_BIAS.n59 9.3005
R15482 DIFFPAIR_BIAS.n33 DIFFPAIR_BIAS.n32 9.3005
R15483 DIFFPAIR_BIAS.n54 DIFFPAIR_BIAS.n53 9.3005
R15484 DIFFPAIR_BIAS.n52 DIFFPAIR_BIAS.n51 9.3005
R15485 DIFFPAIR_BIAS.n37 DIFFPAIR_BIAS.n36 9.3005
R15486 DIFFPAIR_BIAS.n46 DIFFPAIR_BIAS.n45 9.3005
R15487 DIFFPAIR_BIAS.n44 DIFFPAIR_BIAS.n43 9.3005
R15488 DIFFPAIR_BIAS.n92 DIFFPAIR_BIAS.n91 9.3005
R15489 DIFFPAIR_BIAS.n65 DIFFPAIR_BIAS.n64 9.3005
R15490 DIFFPAIR_BIAS.n86 DIFFPAIR_BIAS.n85 9.3005
R15491 DIFFPAIR_BIAS.n84 DIFFPAIR_BIAS.n83 9.3005
R15492 DIFFPAIR_BIAS.n69 DIFFPAIR_BIAS.n68 9.3005
R15493 DIFFPAIR_BIAS.n78 DIFFPAIR_BIAS.n77 9.3005
R15494 DIFFPAIR_BIAS.n76 DIFFPAIR_BIAS.n75 9.3005
R15495 DIFFPAIR_BIAS.n27 DIFFPAIR_BIAS.n2 8.92171
R15496 DIFFPAIR_BIAS.n58 DIFFPAIR_BIAS.n33 8.92171
R15497 DIFFPAIR_BIAS.n90 DIFFPAIR_BIAS.n65 8.92171
R15498 DIFFPAIR_BIAS.n28 DIFFPAIR_BIAS.n0 8.14595
R15499 DIFFPAIR_BIAS.n59 DIFFPAIR_BIAS.n31 8.14595
R15500 DIFFPAIR_BIAS.n91 DIFFPAIR_BIAS.n63 8.14595
R15501 DIFFPAIR_BIAS.n30 DIFFPAIR_BIAS.n0 5.81868
R15502 DIFFPAIR_BIAS.n61 DIFFPAIR_BIAS.n31 5.81868
R15503 DIFFPAIR_BIAS.n93 DIFFPAIR_BIAS.n63 5.81868
R15504 DIFFPAIR_BIAS.n97 DIFFPAIR_BIAS.n96 5.21819
R15505 DIFFPAIR_BIAS.n97 DIFFPAIR_BIAS.n94 5.12393
R15506 DIFFPAIR_BIAS.n28 DIFFPAIR_BIAS.n27 5.04292
R15507 DIFFPAIR_BIAS.n59 DIFFPAIR_BIAS.n58 5.04292
R15508 DIFFPAIR_BIAS.n91 DIFFPAIR_BIAS.n90 5.04292
R15509 DIFFPAIR_BIAS.n13 DIFFPAIR_BIAS.n9 4.38594
R15510 DIFFPAIR_BIAS.n44 DIFFPAIR_BIAS.n40 4.38594
R15511 DIFFPAIR_BIAS.n76 DIFFPAIR_BIAS.n72 4.38594
R15512 DIFFPAIR_BIAS.n98 DIFFPAIR_BIAS.n97 4.28744
R15513 DIFFPAIR_BIAS.n24 DIFFPAIR_BIAS.n2 4.26717
R15514 DIFFPAIR_BIAS.n55 DIFFPAIR_BIAS.n33 4.26717
R15515 DIFFPAIR_BIAS.n87 DIFFPAIR_BIAS.n65 4.26717
R15516 DIFFPAIR_BIAS.n23 DIFFPAIR_BIAS.n4 3.49141
R15517 DIFFPAIR_BIAS.n54 DIFFPAIR_BIAS.n35 3.49141
R15518 DIFFPAIR_BIAS.n86 DIFFPAIR_BIAS.n67 3.49141
R15519 DIFFPAIR_BIAS.n20 DIFFPAIR_BIAS.n19 2.71565
R15520 DIFFPAIR_BIAS.n51 DIFFPAIR_BIAS.n50 2.71565
R15521 DIFFPAIR_BIAS.n83 DIFFPAIR_BIAS.n82 2.71565
R15522 DIFFPAIR_BIAS.n16 DIFFPAIR_BIAS.n6 1.93989
R15523 DIFFPAIR_BIAS.n47 DIFFPAIR_BIAS.n37 1.93989
R15524 DIFFPAIR_BIAS.n79 DIFFPAIR_BIAS.n69 1.93989
R15525 DIFFPAIR_BIAS.n96 DIFFPAIR_BIAS.n95 1.93823
R15526 DIFFPAIR_BIAS.n99 DIFFPAIR_BIAS.n98 1.9382
R15527 DIFFPAIR_BIAS.n94 DIFFPAIR_BIAS.n62 1.93655
R15528 DIFFPAIR_BIAS.n15 DIFFPAIR_BIAS.n8 1.16414
R15529 DIFFPAIR_BIAS.n46 DIFFPAIR_BIAS.n39 1.16414
R15530 DIFFPAIR_BIAS.n78 DIFFPAIR_BIAS.n71 1.16414
R15531 DIFFPAIR_BIAS DIFFPAIR_BIAS.n100 0.6855
R15532 DIFFPAIR_BIAS.n12 DIFFPAIR_BIAS.n11 0.388379
R15533 DIFFPAIR_BIAS.n43 DIFFPAIR_BIAS.n42 0.388379
R15534 DIFFPAIR_BIAS.n75 DIFFPAIR_BIAS.n74 0.388379
R15535 DIFFPAIR_BIAS.n100 DIFFPAIR_BIAS.n99 0.339824
R15536 DIFFPAIR_BIAS.n29 DIFFPAIR_BIAS.n1 0.155672
R15537 DIFFPAIR_BIAS.n22 DIFFPAIR_BIAS.n1 0.155672
R15538 DIFFPAIR_BIAS.n22 DIFFPAIR_BIAS.n21 0.155672
R15539 DIFFPAIR_BIAS.n21 DIFFPAIR_BIAS.n5 0.155672
R15540 DIFFPAIR_BIAS.n14 DIFFPAIR_BIAS.n5 0.155672
R15541 DIFFPAIR_BIAS.n14 DIFFPAIR_BIAS.n13 0.155672
R15542 DIFFPAIR_BIAS.n60 DIFFPAIR_BIAS.n32 0.155672
R15543 DIFFPAIR_BIAS.n53 DIFFPAIR_BIAS.n32 0.155672
R15544 DIFFPAIR_BIAS.n53 DIFFPAIR_BIAS.n52 0.155672
R15545 DIFFPAIR_BIAS.n52 DIFFPAIR_BIAS.n36 0.155672
R15546 DIFFPAIR_BIAS.n45 DIFFPAIR_BIAS.n36 0.155672
R15547 DIFFPAIR_BIAS.n45 DIFFPAIR_BIAS.n44 0.155672
R15548 DIFFPAIR_BIAS.n92 DIFFPAIR_BIAS.n64 0.155672
R15549 DIFFPAIR_BIAS.n85 DIFFPAIR_BIAS.n64 0.155672
R15550 DIFFPAIR_BIAS.n85 DIFFPAIR_BIAS.n84 0.155672
R15551 DIFFPAIR_BIAS.n84 DIFFPAIR_BIAS.n68 0.155672
R15552 DIFFPAIR_BIAS.n77 DIFFPAIR_BIAS.n68 0.155672
R15553 DIFFPAIR_BIAS.n77 DIFFPAIR_BIAS.n76 0.155672
R15554 a_n1945_n3383.n34 a_n1945_n3383.n18 289.615
R15555 a_n1945_n3383.n54 a_n1945_n3383.n38 289.615
R15556 a_n1945_n3383.n60 a_n1945_n3383.n16 289.615
R15557 a_n1945_n3383.n35 a_n1945_n3383.n34 185
R15558 a_n1945_n3383.n33 a_n1945_n3383.n32 185
R15559 a_n1945_n3383.n21 a_n1945_n3383.n20 185
R15560 a_n1945_n3383.n29 a_n1945_n3383.n28 185
R15561 a_n1945_n3383.n27 a_n1945_n3383.n26 185
R15562 a_n1945_n3383.n4 a_n1945_n3383.n23 185
R15563 a_n1945_n3383.n5 a_n1945_n3383.n24 185
R15564 a_n1945_n3383.n55 a_n1945_n3383.n54 185
R15565 a_n1945_n3383.n53 a_n1945_n3383.n52 185
R15566 a_n1945_n3383.n41 a_n1945_n3383.n40 185
R15567 a_n1945_n3383.n49 a_n1945_n3383.n48 185
R15568 a_n1945_n3383.n47 a_n1945_n3383.n46 185
R15569 a_n1945_n3383.n7 a_n1945_n3383.n43 185
R15570 a_n1945_n3383.n8 a_n1945_n3383.n44 185
R15571 a_n1945_n3383.n17 a_n1945_n3383.n16 185
R15572 a_n1945_n3383.n64 a_n1945_n3383.n63 185
R15573 a_n1945_n3383.n66 a_n1945_n3383.n65 185
R15574 a_n1945_n3383.n14 a_n1945_n3383.n13 185
R15575 a_n1945_n3383.n70 a_n1945_n3383.n69 185
R15576 a_n1945_n3383.n72 a_n1945_n3383.n71 185
R15577 a_n1945_n3383.n10 a_n1945_n3383.n9 185
R15578 a_n1945_n3383.n34 a_n1945_n3383.n33 104.615
R15579 a_n1945_n3383.n33 a_n1945_n3383.n20 104.615
R15580 a_n1945_n3383.n28 a_n1945_n3383.n20 104.615
R15581 a_n1945_n3383.n28 a_n1945_n3383.n27 104.615
R15582 a_n1945_n3383.n27 a_n1945_n3383.n23 104.615
R15583 a_n1945_n3383.n24 a_n1945_n3383.n23 104.615
R15584 a_n1945_n3383.n54 a_n1945_n3383.n53 104.615
R15585 a_n1945_n3383.n53 a_n1945_n3383.n40 104.615
R15586 a_n1945_n3383.n48 a_n1945_n3383.n40 104.615
R15587 a_n1945_n3383.n48 a_n1945_n3383.n47 104.615
R15588 a_n1945_n3383.n47 a_n1945_n3383.n43 104.615
R15589 a_n1945_n3383.n44 a_n1945_n3383.n43 104.615
R15590 a_n1945_n3383.n64 a_n1945_n3383.n16 104.615
R15591 a_n1945_n3383.n65 a_n1945_n3383.n64 104.615
R15592 a_n1945_n3383.n65 a_n1945_n3383.n13 104.615
R15593 a_n1945_n3383.n70 a_n1945_n3383.n13 104.615
R15594 a_n1945_n3383.n71 a_n1945_n3383.n70 104.615
R15595 a_n1945_n3383.n71 a_n1945_n3383.n9 104.615
R15596 a_n1945_n3383.n24 a_n1945_n3383.t0 52.3082
R15597 a_n1945_n3383.n44 a_n1945_n3383.t2 52.3082
R15598 a_n1945_n3383.t1 a_n1945_n3383.n9 52.3082
R15599 a_n1945_n3383.n58 a_n1945_n3383.n37 42.5002
R15600 a_n1945_n3383.n59 a_n1945_n3383.n58 42.5002
R15601 a_n1945_n3383.n58 a_n1945_n3383.n57 40.5641
R15602 a_n1945_n3383.n5 a_n1945_n3383.n3 5.10449
R15603 a_n1945_n3383.n8 a_n1945_n3383.n6 5.10449
R15604 a_n1945_n3383.n11 a_n1945_n3383.n10 5.10449
R15605 a_n1945_n3383.n5 a_n1945_n3383.n4 12.8005
R15606 a_n1945_n3383.n8 a_n1945_n3383.n7 12.8005
R15607 a_n1945_n3383.n10 a_n1945_n3383.n72 12.8005
R15608 a_n1945_n3383.n26 a_n1945_n3383.n25 12.0247
R15609 a_n1945_n3383.n46 a_n1945_n3383.n45 12.0247
R15610 a_n1945_n3383.n69 a_n1945_n3383.n12 12.0247
R15611 a_n1945_n3383.n29 a_n1945_n3383.n22 11.249
R15612 a_n1945_n3383.n49 a_n1945_n3383.n42 11.249
R15613 a_n1945_n3383.n68 a_n1945_n3383.n14 11.249
R15614 a_n1945_n3383.n30 a_n1945_n3383.n21 10.4732
R15615 a_n1945_n3383.n50 a_n1945_n3383.n41 10.4732
R15616 a_n1945_n3383.n67 a_n1945_n3383.n66 10.4732
R15617 a_n1945_n3383.n32 a_n1945_n3383.n31 9.69747
R15618 a_n1945_n3383.n52 a_n1945_n3383.n51 9.69747
R15619 a_n1945_n3383.n63 a_n1945_n3383.n15 9.69747
R15620 a_n1945_n3383.n37 a_n1945_n3383.n0 9.45567
R15621 a_n1945_n3383.n57 a_n1945_n3383.n1 9.45567
R15622 a_n1945_n3383.n2 a_n1945_n3383.n59 9.45567
R15623 a_n1945_n3383.n0 a_n1945_n3383.n36 9.3005
R15624 a_n1945_n3383.n19 a_n1945_n3383.n0 9.3005
R15625 a_n1945_n3383.n31 a_n1945_n3383.n0 9.3005
R15626 a_n1945_n3383.n0 a_n1945_n3383.n30 9.3005
R15627 a_n1945_n3383.n22 a_n1945_n3383.n0 9.3005
R15628 a_n1945_n3383.n25 a_n1945_n3383.n0 9.3005
R15629 a_n1945_n3383.n1 a_n1945_n3383.n56 9.3005
R15630 a_n1945_n3383.n39 a_n1945_n3383.n1 9.3005
R15631 a_n1945_n3383.n51 a_n1945_n3383.n1 9.3005
R15632 a_n1945_n3383.n1 a_n1945_n3383.n50 9.3005
R15633 a_n1945_n3383.n42 a_n1945_n3383.n1 9.3005
R15634 a_n1945_n3383.n45 a_n1945_n3383.n1 9.3005
R15635 a_n1945_n3383.n2 a_n1945_n3383.n61 9.3005
R15636 a_n1945_n3383.n62 a_n1945_n3383.n2 9.3005
R15637 a_n1945_n3383.n15 a_n1945_n3383.n2 9.3005
R15638 a_n1945_n3383.n2 a_n1945_n3383.n67 9.3005
R15639 a_n1945_n3383.n68 a_n1945_n3383.n2 9.3005
R15640 a_n1945_n3383.n2 a_n1945_n3383.n12 9.3005
R15641 a_n1945_n3383.n35 a_n1945_n3383.n19 8.92171
R15642 a_n1945_n3383.n55 a_n1945_n3383.n39 8.92171
R15643 a_n1945_n3383.n62 a_n1945_n3383.n17 8.92171
R15644 a_n1945_n3383.n36 a_n1945_n3383.n18 8.14595
R15645 a_n1945_n3383.n56 a_n1945_n3383.n38 8.14595
R15646 a_n1945_n3383.n61 a_n1945_n3383.n60 8.14595
R15647 a_n1945_n3383.n37 a_n1945_n3383.n18 5.81868
R15648 a_n1945_n3383.n57 a_n1945_n3383.n38 5.81868
R15649 a_n1945_n3383.n60 a_n1945_n3383.n59 5.81868
R15650 a_n1945_n3383.n36 a_n1945_n3383.n35 5.04292
R15651 a_n1945_n3383.n56 a_n1945_n3383.n55 5.04292
R15652 a_n1945_n3383.n61 a_n1945_n3383.n17 5.04292
R15653 a_n1945_n3383.n3 a_n1945_n3383.t0 149.972
R15654 a_n1945_n3383.n6 a_n1945_n3383.t2 149.972
R15655 a_n1945_n3383.t1 a_n1945_n3383.n11 149.972
R15656 a_n1945_n3383.n32 a_n1945_n3383.n19 4.26717
R15657 a_n1945_n3383.n52 a_n1945_n3383.n39 4.26717
R15658 a_n1945_n3383.n63 a_n1945_n3383.n62 4.26717
R15659 a_n1945_n3383.n31 a_n1945_n3383.n21 3.49141
R15660 a_n1945_n3383.n51 a_n1945_n3383.n41 3.49141
R15661 a_n1945_n3383.n66 a_n1945_n3383.n15 3.49141
R15662 a_n1945_n3383.n30 a_n1945_n3383.n29 2.71565
R15663 a_n1945_n3383.n50 a_n1945_n3383.n49 2.71565
R15664 a_n1945_n3383.n67 a_n1945_n3383.n14 2.71565
R15665 a_n1945_n3383.n11 a_n1945_n3383.n2 2.36059
R15666 a_n1945_n3383.n1 a_n1945_n3383.n6 2.36059
R15667 a_n1945_n3383.n0 a_n1945_n3383.n3 2.36059
R15668 a_n1945_n3383.n26 a_n1945_n3383.n22 1.93989
R15669 a_n1945_n3383.n46 a_n1945_n3383.n42 1.93989
R15670 a_n1945_n3383.n69 a_n1945_n3383.n68 1.93989
R15671 a_n1945_n3383.n25 a_n1945_n3383.n4 1.16414
R15672 a_n1945_n3383.n45 a_n1945_n3383.n7 1.16414
R15673 a_n1945_n3383.n72 a_n1945_n3383.n12 1.16414
R15674 a_n1279_n3383.n54 a_n1279_n3383.n38 289.615
R15675 a_n1279_n3383.n34 a_n1279_n3383.n18 289.615
R15676 a_n1279_n3383.n60 a_n1279_n3383.n16 289.615
R15677 a_n1279_n3383.n55 a_n1279_n3383.n54 185
R15678 a_n1279_n3383.n53 a_n1279_n3383.n52 185
R15679 a_n1279_n3383.n41 a_n1279_n3383.n40 185
R15680 a_n1279_n3383.n49 a_n1279_n3383.n48 185
R15681 a_n1279_n3383.n47 a_n1279_n3383.n46 185
R15682 a_n1279_n3383.n4 a_n1279_n3383.n43 185
R15683 a_n1279_n3383.n5 a_n1279_n3383.n44 185
R15684 a_n1279_n3383.n35 a_n1279_n3383.n34 185
R15685 a_n1279_n3383.n33 a_n1279_n3383.n32 185
R15686 a_n1279_n3383.n21 a_n1279_n3383.n20 185
R15687 a_n1279_n3383.n29 a_n1279_n3383.n28 185
R15688 a_n1279_n3383.n27 a_n1279_n3383.n26 185
R15689 a_n1279_n3383.n7 a_n1279_n3383.n23 185
R15690 a_n1279_n3383.n8 a_n1279_n3383.n24 185
R15691 a_n1279_n3383.n17 a_n1279_n3383.n16 185
R15692 a_n1279_n3383.n64 a_n1279_n3383.n63 185
R15693 a_n1279_n3383.n66 a_n1279_n3383.n65 185
R15694 a_n1279_n3383.n14 a_n1279_n3383.n13 185
R15695 a_n1279_n3383.n70 a_n1279_n3383.n69 185
R15696 a_n1279_n3383.n72 a_n1279_n3383.n71 185
R15697 a_n1279_n3383.n10 a_n1279_n3383.n9 185
R15698 a_n1279_n3383.n58 a_n1279_n3383.n57 110.766
R15699 a_n1279_n3383.n58 a_n1279_n3383.n37 110.766
R15700 a_n1279_n3383.n59 a_n1279_n3383.n58 108.831
R15701 a_n1279_n3383.n54 a_n1279_n3383.n53 104.615
R15702 a_n1279_n3383.n53 a_n1279_n3383.n40 104.615
R15703 a_n1279_n3383.n48 a_n1279_n3383.n40 104.615
R15704 a_n1279_n3383.n48 a_n1279_n3383.n47 104.615
R15705 a_n1279_n3383.n47 a_n1279_n3383.n43 104.615
R15706 a_n1279_n3383.n44 a_n1279_n3383.n43 104.615
R15707 a_n1279_n3383.n34 a_n1279_n3383.n33 104.615
R15708 a_n1279_n3383.n33 a_n1279_n3383.n20 104.615
R15709 a_n1279_n3383.n28 a_n1279_n3383.n20 104.615
R15710 a_n1279_n3383.n28 a_n1279_n3383.n27 104.615
R15711 a_n1279_n3383.n27 a_n1279_n3383.n23 104.615
R15712 a_n1279_n3383.n24 a_n1279_n3383.n23 104.615
R15713 a_n1279_n3383.n64 a_n1279_n3383.n16 104.615
R15714 a_n1279_n3383.n65 a_n1279_n3383.n64 104.615
R15715 a_n1279_n3383.n65 a_n1279_n3383.n13 104.615
R15716 a_n1279_n3383.n70 a_n1279_n3383.n13 104.615
R15717 a_n1279_n3383.n71 a_n1279_n3383.n70 104.615
R15718 a_n1279_n3383.n71 a_n1279_n3383.n9 104.615
R15719 a_n1279_n3383.n44 a_n1279_n3383.t2 52.3082
R15720 a_n1279_n3383.n24 a_n1279_n3383.t0 52.3082
R15721 a_n1279_n3383.t1 a_n1279_n3383.n9 52.3082
R15722 a_n1279_n3383.n5 a_n1279_n3383.n3 5.10449
R15723 a_n1279_n3383.n8 a_n1279_n3383.n6 5.10449
R15724 a_n1279_n3383.n11 a_n1279_n3383.n10 5.10449
R15725 a_n1279_n3383.n5 a_n1279_n3383.n4 12.8005
R15726 a_n1279_n3383.n8 a_n1279_n3383.n7 12.8005
R15727 a_n1279_n3383.n10 a_n1279_n3383.n72 12.8005
R15728 a_n1279_n3383.n46 a_n1279_n3383.n45 12.0247
R15729 a_n1279_n3383.n26 a_n1279_n3383.n25 12.0247
R15730 a_n1279_n3383.n69 a_n1279_n3383.n12 12.0247
R15731 a_n1279_n3383.n49 a_n1279_n3383.n42 11.249
R15732 a_n1279_n3383.n29 a_n1279_n3383.n22 11.249
R15733 a_n1279_n3383.n68 a_n1279_n3383.n14 11.249
R15734 a_n1279_n3383.n50 a_n1279_n3383.n41 10.4732
R15735 a_n1279_n3383.n30 a_n1279_n3383.n21 10.4732
R15736 a_n1279_n3383.n67 a_n1279_n3383.n66 10.4732
R15737 a_n1279_n3383.n52 a_n1279_n3383.n51 9.69747
R15738 a_n1279_n3383.n32 a_n1279_n3383.n31 9.69747
R15739 a_n1279_n3383.n63 a_n1279_n3383.n15 9.69747
R15740 a_n1279_n3383.n57 a_n1279_n3383.n0 9.45567
R15741 a_n1279_n3383.n37 a_n1279_n3383.n1 9.45567
R15742 a_n1279_n3383.n2 a_n1279_n3383.n59 9.45567
R15743 a_n1279_n3383.n0 a_n1279_n3383.n56 9.3005
R15744 a_n1279_n3383.n39 a_n1279_n3383.n0 9.3005
R15745 a_n1279_n3383.n51 a_n1279_n3383.n0 9.3005
R15746 a_n1279_n3383.n0 a_n1279_n3383.n50 9.3005
R15747 a_n1279_n3383.n42 a_n1279_n3383.n0 9.3005
R15748 a_n1279_n3383.n45 a_n1279_n3383.n0 9.3005
R15749 a_n1279_n3383.n1 a_n1279_n3383.n36 9.3005
R15750 a_n1279_n3383.n19 a_n1279_n3383.n1 9.3005
R15751 a_n1279_n3383.n31 a_n1279_n3383.n1 9.3005
R15752 a_n1279_n3383.n1 a_n1279_n3383.n30 9.3005
R15753 a_n1279_n3383.n22 a_n1279_n3383.n1 9.3005
R15754 a_n1279_n3383.n25 a_n1279_n3383.n1 9.3005
R15755 a_n1279_n3383.n2 a_n1279_n3383.n61 9.3005
R15756 a_n1279_n3383.n62 a_n1279_n3383.n2 9.3005
R15757 a_n1279_n3383.n15 a_n1279_n3383.n2 9.3005
R15758 a_n1279_n3383.n2 a_n1279_n3383.n67 9.3005
R15759 a_n1279_n3383.n68 a_n1279_n3383.n2 9.3005
R15760 a_n1279_n3383.n2 a_n1279_n3383.n12 9.3005
R15761 a_n1279_n3383.n55 a_n1279_n3383.n39 8.92171
R15762 a_n1279_n3383.n35 a_n1279_n3383.n19 8.92171
R15763 a_n1279_n3383.n62 a_n1279_n3383.n17 8.92171
R15764 a_n1279_n3383.n56 a_n1279_n3383.n38 8.14595
R15765 a_n1279_n3383.n36 a_n1279_n3383.n18 8.14595
R15766 a_n1279_n3383.n61 a_n1279_n3383.n60 8.14595
R15767 a_n1279_n3383.n57 a_n1279_n3383.n38 5.81868
R15768 a_n1279_n3383.n37 a_n1279_n3383.n18 5.81868
R15769 a_n1279_n3383.n60 a_n1279_n3383.n59 5.81868
R15770 a_n1279_n3383.n56 a_n1279_n3383.n55 5.04292
R15771 a_n1279_n3383.n36 a_n1279_n3383.n35 5.04292
R15772 a_n1279_n3383.n61 a_n1279_n3383.n17 5.04292
R15773 a_n1279_n3383.n3 a_n1279_n3383.t2 149.972
R15774 a_n1279_n3383.n6 a_n1279_n3383.t0 149.972
R15775 a_n1279_n3383.t1 a_n1279_n3383.n11 149.972
R15776 a_n1279_n3383.n52 a_n1279_n3383.n39 4.26717
R15777 a_n1279_n3383.n32 a_n1279_n3383.n19 4.26717
R15778 a_n1279_n3383.n63 a_n1279_n3383.n62 4.26717
R15779 a_n1279_n3383.n51 a_n1279_n3383.n41 3.49141
R15780 a_n1279_n3383.n31 a_n1279_n3383.n21 3.49141
R15781 a_n1279_n3383.n66 a_n1279_n3383.n15 3.49141
R15782 a_n1279_n3383.n50 a_n1279_n3383.n49 2.71565
R15783 a_n1279_n3383.n30 a_n1279_n3383.n29 2.71565
R15784 a_n1279_n3383.n67 a_n1279_n3383.n14 2.71565
R15785 a_n1279_n3383.n11 a_n1279_n3383.n2 2.36059
R15786 a_n1279_n3383.n1 a_n1279_n3383.n6 2.36059
R15787 a_n1279_n3383.n0 a_n1279_n3383.n3 2.36059
R15788 a_n1279_n3383.n46 a_n1279_n3383.n42 1.93989
R15789 a_n1279_n3383.n26 a_n1279_n3383.n22 1.93989
R15790 a_n1279_n3383.n69 a_n1279_n3383.n68 1.93989
R15791 a_n1279_n3383.n45 a_n1279_n3383.n4 1.16414
R15792 a_n1279_n3383.n25 a_n1279_n3383.n7 1.16414
R15793 a_n1279_n3383.n72 a_n1279_n3383.n12 1.16414
C0 VN DIFFPAIR_BIAS 0.012812f
C1 a_5714_9514# VDD 1.18258f
C2 VDD VOUT 36.1872f
C3 a_n6412_9514# VDD 1.18304f
C4 VOUT VP 3.11141f
C5 VDD VN 0.093182f
C6 VOUT VN 0.881137f
C7 VP VN 9.36455f
C8 VOUT CS_BIAS 8.9821f
C9 VP CS_BIAS 0.441231f
C10 VN CS_BIAS 0.395109f
C11 VP DIFFPAIR_BIAS 0.013013f
C12 DIFFPAIR_BIAS GND 16.627352f
C13 CS_BIAS GND 59.813557f
C14 VN GND 33.28204f
C15 VP GND 27.987982f
C16 VOUT GND 64.13233f
C17 VDD GND 0.472657p
C18 a_5714_9514# GND 0.847588f
C19 a_n6412_9514# GND 0.845641f
C20 a_n1279_n3383.n0 GND 0.734167f
C21 a_n1279_n3383.n1 GND 0.734167f
C22 a_n1279_n3383.n2 GND 0.734167f
C23 a_n1279_n3383.n3 GND 0.100457f
C24 a_n1279_n3383.n4 GND 0.013636f
C25 a_n1279_n3383.n5 GND 0.03086f
C26 a_n1279_n3383.n6 GND 0.100457f
C27 a_n1279_n3383.n7 GND 0.013636f
C28 a_n1279_n3383.n8 GND 0.03086f
C29 a_n1279_n3383.n9 GND 0.02283f
C30 a_n1279_n3383.n10 GND 0.03086f
C31 a_n1279_n3383.n11 GND 0.100457f
C32 a_n1279_n3383.n12 GND 0.012879f
C33 a_n1279_n3383.n13 GND 0.030441f
C34 a_n1279_n3383.n14 GND 0.013636f
C35 a_n1279_n3383.n15 GND 0.012879f
C36 a_n1279_n3383.n16 GND 0.063611f
C37 a_n1279_n3383.n17 GND 0.013636f
C38 a_n1279_n3383.n18 GND 0.032394f
C39 a_n1279_n3383.n19 GND 0.012879f
C40 a_n1279_n3383.n20 GND 0.030441f
C41 a_n1279_n3383.n21 GND 0.013636f
C42 a_n1279_n3383.n22 GND 0.012879f
C43 a_n1279_n3383.n23 GND 0.030441f
C44 a_n1279_n3383.t0 GND 0.051155f
C45 a_n1279_n3383.n24 GND 0.02283f
C46 a_n1279_n3383.n25 GND 0.012879f
C47 a_n1279_n3383.n26 GND 0.013636f
C48 a_n1279_n3383.n27 GND 0.030441f
C49 a_n1279_n3383.n28 GND 0.030441f
C50 a_n1279_n3383.n29 GND 0.013636f
C51 a_n1279_n3383.n30 GND 0.012879f
C52 a_n1279_n3383.n31 GND 0.012879f
C53 a_n1279_n3383.n32 GND 0.013636f
C54 a_n1279_n3383.n33 GND 0.030441f
C55 a_n1279_n3383.n34 GND 0.063611f
C56 a_n1279_n3383.n35 GND 0.013636f
C57 a_n1279_n3383.n36 GND 0.012879f
C58 a_n1279_n3383.n37 GND 0.132341f
C59 a_n1279_n3383.n38 GND 0.032394f
C60 a_n1279_n3383.n39 GND 0.012879f
C61 a_n1279_n3383.n40 GND 0.030441f
C62 a_n1279_n3383.n41 GND 0.013636f
C63 a_n1279_n3383.n42 GND 0.012879f
C64 a_n1279_n3383.n43 GND 0.030441f
C65 a_n1279_n3383.t2 GND 0.051155f
C66 a_n1279_n3383.n44 GND 0.02283f
C67 a_n1279_n3383.n45 GND 0.012879f
C68 a_n1279_n3383.n46 GND 0.013636f
C69 a_n1279_n3383.n47 GND 0.030441f
C70 a_n1279_n3383.n48 GND 0.030441f
C71 a_n1279_n3383.n49 GND 0.013636f
C72 a_n1279_n3383.n50 GND 0.012879f
C73 a_n1279_n3383.n51 GND 0.012879f
C74 a_n1279_n3383.n52 GND 0.013636f
C75 a_n1279_n3383.n53 GND 0.030441f
C76 a_n1279_n3383.n54 GND 0.063611f
C77 a_n1279_n3383.n55 GND 0.013636f
C78 a_n1279_n3383.n56 GND 0.012879f
C79 a_n1279_n3383.n57 GND 0.137311f
C80 a_n1279_n3383.n58 GND 2.57074f
C81 a_n1279_n3383.n59 GND 0.119308f
C82 a_n1279_n3383.n60 GND 0.032394f
C83 a_n1279_n3383.n61 GND 0.012879f
C84 a_n1279_n3383.n62 GND 0.012879f
C85 a_n1279_n3383.n63 GND 0.013636f
C86 a_n1279_n3383.n64 GND 0.030441f
C87 a_n1279_n3383.n65 GND 0.030441f
C88 a_n1279_n3383.n66 GND 0.013636f
C89 a_n1279_n3383.n67 GND 0.012879f
C90 a_n1279_n3383.n68 GND 0.012879f
C91 a_n1279_n3383.n69 GND 0.013636f
C92 a_n1279_n3383.n70 GND 0.030441f
C93 a_n1279_n3383.n71 GND 0.030441f
C94 a_n1279_n3383.n72 GND 0.013636f
C95 a_n1279_n3383.t1 GND 0.051155f
C96 a_n1945_n3383.n0 GND 0.471965f
C97 a_n1945_n3383.n1 GND 0.471965f
C98 a_n1945_n3383.n2 GND 0.471965f
C99 a_n1945_n3383.n3 GND 0.06458f
C100 a_n1945_n3383.n4 GND 0.008766f
C101 a_n1945_n3383.n5 GND 0.019838f
C102 a_n1945_n3383.n6 GND 0.06458f
C103 a_n1945_n3383.n7 GND 0.008766f
C104 a_n1945_n3383.n8 GND 0.019838f
C105 a_n1945_n3383.n9 GND 0.014677f
C106 a_n1945_n3383.n10 GND 0.019838f
C107 a_n1945_n3383.n11 GND 0.06458f
C108 a_n1945_n3383.n12 GND 0.008279f
C109 a_n1945_n3383.n13 GND 0.019569f
C110 a_n1945_n3383.n14 GND 0.008766f
C111 a_n1945_n3383.n15 GND 0.008279f
C112 a_n1945_n3383.n16 GND 0.040893f
C113 a_n1945_n3383.n17 GND 0.008766f
C114 a_n1945_n3383.n18 GND 0.020825f
C115 a_n1945_n3383.n19 GND 0.008279f
C116 a_n1945_n3383.n20 GND 0.019569f
C117 a_n1945_n3383.n21 GND 0.008766f
C118 a_n1945_n3383.n22 GND 0.008279f
C119 a_n1945_n3383.n23 GND 0.019569f
C120 a_n1945_n3383.t0 GND 0.032885f
C121 a_n1945_n3383.n24 GND 0.014677f
C122 a_n1945_n3383.n25 GND 0.008279f
C123 a_n1945_n3383.n26 GND 0.008766f
C124 a_n1945_n3383.n27 GND 0.019569f
C125 a_n1945_n3383.n28 GND 0.019569f
C126 a_n1945_n3383.n29 GND 0.008766f
C127 a_n1945_n3383.n30 GND 0.008279f
C128 a_n1945_n3383.n31 GND 0.008279f
C129 a_n1945_n3383.n32 GND 0.008766f
C130 a_n1945_n3383.n33 GND 0.019569f
C131 a_n1945_n3383.n34 GND 0.040893f
C132 a_n1945_n3383.n35 GND 0.008766f
C133 a_n1945_n3383.n36 GND 0.008279f
C134 a_n1945_n3383.n37 GND 0.091252f
C135 a_n1945_n3383.n38 GND 0.020825f
C136 a_n1945_n3383.n39 GND 0.008279f
C137 a_n1945_n3383.n40 GND 0.019569f
C138 a_n1945_n3383.n41 GND 0.008766f
C139 a_n1945_n3383.n42 GND 0.008279f
C140 a_n1945_n3383.n43 GND 0.019569f
C141 a_n1945_n3383.t2 GND 0.032885f
C142 a_n1945_n3383.n44 GND 0.014677f
C143 a_n1945_n3383.n45 GND 0.008279f
C144 a_n1945_n3383.n46 GND 0.008766f
C145 a_n1945_n3383.n47 GND 0.019569f
C146 a_n1945_n3383.n48 GND 0.019569f
C147 a_n1945_n3383.n49 GND 0.008766f
C148 a_n1945_n3383.n50 GND 0.008279f
C149 a_n1945_n3383.n51 GND 0.008279f
C150 a_n1945_n3383.n52 GND 0.008766f
C151 a_n1945_n3383.n53 GND 0.019569f
C152 a_n1945_n3383.n54 GND 0.040893f
C153 a_n1945_n3383.n55 GND 0.008766f
C154 a_n1945_n3383.n56 GND 0.008279f
C155 a_n1945_n3383.n57 GND 0.070431f
C156 a_n1945_n3383.n58 GND 1.6388f
C157 a_n1945_n3383.n59 GND 0.10218f
C158 a_n1945_n3383.n60 GND 0.020825f
C159 a_n1945_n3383.n61 GND 0.008279f
C160 a_n1945_n3383.n62 GND 0.008279f
C161 a_n1945_n3383.n63 GND 0.008766f
C162 a_n1945_n3383.n64 GND 0.019569f
C163 a_n1945_n3383.n65 GND 0.019569f
C164 a_n1945_n3383.n66 GND 0.008766f
C165 a_n1945_n3383.n67 GND 0.008279f
C166 a_n1945_n3383.n68 GND 0.008279f
C167 a_n1945_n3383.n69 GND 0.008766f
C168 a_n1945_n3383.n70 GND 0.019569f
C169 a_n1945_n3383.n71 GND 0.019569f
C170 a_n1945_n3383.n72 GND 0.008766f
C171 a_n1945_n3383.t1 GND 0.032885f
C172 DIFFPAIR_BIAS.t6 GND 0.595909f
C173 DIFFPAIR_BIAS.n0 GND 0.006812f
C174 DIFFPAIR_BIAS.n1 GND 0.00504f
C175 DIFFPAIR_BIAS.n2 GND 0.002708f
C176 DIFFPAIR_BIAS.n3 GND 0.006402f
C177 DIFFPAIR_BIAS.n4 GND 0.002868f
C178 DIFFPAIR_BIAS.n5 GND 0.00504f
C179 DIFFPAIR_BIAS.n6 GND 0.002708f
C180 DIFFPAIR_BIAS.n7 GND 0.006402f
C181 DIFFPAIR_BIAS.n8 GND 0.002868f
C182 DIFFPAIR_BIAS.n9 GND 0.021456f
C183 DIFFPAIR_BIAS.t3 GND 0.010427f
C184 DIFFPAIR_BIAS.n10 GND 0.004801f
C185 DIFFPAIR_BIAS.n11 GND 0.003781f
C186 DIFFPAIR_BIAS.n12 GND 0.002708f
C187 DIFFPAIR_BIAS.n13 GND 0.118093f
C188 DIFFPAIR_BIAS.n14 GND 0.00504f
C189 DIFFPAIR_BIAS.n15 GND 0.002708f
C190 DIFFPAIR_BIAS.n16 GND 0.002868f
C191 DIFFPAIR_BIAS.n17 GND 0.006402f
C192 DIFFPAIR_BIAS.n18 GND 0.006402f
C193 DIFFPAIR_BIAS.n19 GND 0.002868f
C194 DIFFPAIR_BIAS.n20 GND 0.002708f
C195 DIFFPAIR_BIAS.n21 GND 0.00504f
C196 DIFFPAIR_BIAS.n22 GND 0.00504f
C197 DIFFPAIR_BIAS.n23 GND 0.002708f
C198 DIFFPAIR_BIAS.n24 GND 0.002868f
C199 DIFFPAIR_BIAS.n25 GND 0.006402f
C200 DIFFPAIR_BIAS.n26 GND 0.013377f
C201 DIFFPAIR_BIAS.n27 GND 0.002868f
C202 DIFFPAIR_BIAS.n28 GND 0.002708f
C203 DIFFPAIR_BIAS.n29 GND 0.011099f
C204 DIFFPAIR_BIAS.n30 GND 0.025428f
C205 DIFFPAIR_BIAS.n31 GND 0.006812f
C206 DIFFPAIR_BIAS.n32 GND 0.00504f
C207 DIFFPAIR_BIAS.n33 GND 0.002708f
C208 DIFFPAIR_BIAS.n34 GND 0.006402f
C209 DIFFPAIR_BIAS.n35 GND 0.002868f
C210 DIFFPAIR_BIAS.n36 GND 0.00504f
C211 DIFFPAIR_BIAS.n37 GND 0.002708f
C212 DIFFPAIR_BIAS.n38 GND 0.006402f
C213 DIFFPAIR_BIAS.n39 GND 0.002868f
C214 DIFFPAIR_BIAS.n40 GND 0.021456f
C215 DIFFPAIR_BIAS.t1 GND 0.010427f
C216 DIFFPAIR_BIAS.n41 GND 0.004801f
C217 DIFFPAIR_BIAS.n42 GND 0.003781f
C218 DIFFPAIR_BIAS.n43 GND 0.002708f
C219 DIFFPAIR_BIAS.n44 GND 0.118093f
C220 DIFFPAIR_BIAS.n45 GND 0.00504f
C221 DIFFPAIR_BIAS.n46 GND 0.002708f
C222 DIFFPAIR_BIAS.n47 GND 0.002868f
C223 DIFFPAIR_BIAS.n48 GND 0.006402f
C224 DIFFPAIR_BIAS.n49 GND 0.006402f
C225 DIFFPAIR_BIAS.n50 GND 0.002868f
C226 DIFFPAIR_BIAS.n51 GND 0.002708f
C227 DIFFPAIR_BIAS.n52 GND 0.00504f
C228 DIFFPAIR_BIAS.n53 GND 0.00504f
C229 DIFFPAIR_BIAS.n54 GND 0.002708f
C230 DIFFPAIR_BIAS.n55 GND 0.002868f
C231 DIFFPAIR_BIAS.n56 GND 0.006402f
C232 DIFFPAIR_BIAS.n57 GND 0.013377f
C233 DIFFPAIR_BIAS.n58 GND 0.002868f
C234 DIFFPAIR_BIAS.n59 GND 0.002708f
C235 DIFFPAIR_BIAS.n60 GND 0.011099f
C236 DIFFPAIR_BIAS.n61 GND 0.020979f
C237 DIFFPAIR_BIAS.n62 GND 0.334318f
C238 DIFFPAIR_BIAS.n63 GND 0.006812f
C239 DIFFPAIR_BIAS.n64 GND 0.00504f
C240 DIFFPAIR_BIAS.n65 GND 0.002708f
C241 DIFFPAIR_BIAS.n66 GND 0.006402f
C242 DIFFPAIR_BIAS.n67 GND 0.002868f
C243 DIFFPAIR_BIAS.n68 GND 0.00504f
C244 DIFFPAIR_BIAS.n69 GND 0.002708f
C245 DIFFPAIR_BIAS.n70 GND 0.006402f
C246 DIFFPAIR_BIAS.n71 GND 0.002868f
C247 DIFFPAIR_BIAS.n72 GND 0.021456f
C248 DIFFPAIR_BIAS.t5 GND 0.010427f
C249 DIFFPAIR_BIAS.n73 GND 0.004801f
C250 DIFFPAIR_BIAS.n74 GND 0.003781f
C251 DIFFPAIR_BIAS.n75 GND 0.002708f
C252 DIFFPAIR_BIAS.n76 GND 0.118093f
C253 DIFFPAIR_BIAS.n77 GND 0.00504f
C254 DIFFPAIR_BIAS.n78 GND 0.002708f
C255 DIFFPAIR_BIAS.n79 GND 0.002868f
C256 DIFFPAIR_BIAS.n80 GND 0.006402f
C257 DIFFPAIR_BIAS.n81 GND 0.006402f
C258 DIFFPAIR_BIAS.n82 GND 0.002868f
C259 DIFFPAIR_BIAS.n83 GND 0.002708f
C260 DIFFPAIR_BIAS.n84 GND 0.00504f
C261 DIFFPAIR_BIAS.n85 GND 0.00504f
C262 DIFFPAIR_BIAS.n86 GND 0.002708f
C263 DIFFPAIR_BIAS.n87 GND 0.002868f
C264 DIFFPAIR_BIAS.n88 GND 0.006402f
C265 DIFFPAIR_BIAS.n89 GND 0.013377f
C266 DIFFPAIR_BIAS.n90 GND 0.002868f
C267 DIFFPAIR_BIAS.n91 GND 0.002708f
C268 DIFFPAIR_BIAS.n92 GND 0.011099f
C269 DIFFPAIR_BIAS.n93 GND 0.020979f
C270 DIFFPAIR_BIAS.n94 GND 0.216534f
C271 DIFFPAIR_BIAS.t4 GND 0.560233f
C272 DIFFPAIR_BIAS.t0 GND 0.560233f
C273 DIFFPAIR_BIAS.t2 GND 0.565062f
C274 DIFFPAIR_BIAS.n95 GND 0.694826f
C275 DIFFPAIR_BIAS.n96 GND 0.412047f
C276 DIFFPAIR_BIAS.n97 GND 0.798027f
C277 DIFFPAIR_BIAS.t8 GND 0.593255f
C278 DIFFPAIR_BIAS.n98 GND 0.348556f
C279 DIFFPAIR_BIAS.t7 GND 0.593255f
C280 DIFFPAIR_BIAS.n99 GND 0.293801f
C281 DIFFPAIR_BIAS.n100 GND 0.574347f
C282 VN.n0 GND 0.015828f
C283 VN.t8 GND 0.503775f
C284 VN.n1 GND 0.011913f
C285 VN.n2 GND 0.114089f
C286 VN.t5 GND 0.503775f
C287 VN.t4 GND 0.595388f
C288 VN.n3 GND 0.211948f
C289 VN.n4 GND 0.22795f
C290 VN.n5 GND 0.022375f
C291 VN.n6 GND 0.021677f
C292 VN.n7 GND 0.012005f
C293 VN.n8 GND 0.012005f
C294 VN.n9 GND 0.012005f
C295 VN.n10 GND 0.023838f
C296 VN.n11 GND 0.017293f
C297 VN.n12 GND 0.227941f
C298 VN.n13 GND 0.164642f
C299 VN.n14 GND 0.015828f
C300 VN.t7 GND 0.503775f
C301 VN.n15 GND 0.011913f
C302 VN.n16 GND 0.114089f
C303 VN.t6 GND 0.503775f
C304 VN.t3 GND 0.595388f
C305 VN.n17 GND 0.211948f
C306 VN.n18 GND 0.22795f
C307 VN.n19 GND 0.022375f
C308 VN.n20 GND 0.021677f
C309 VN.n21 GND 0.012005f
C310 VN.n22 GND 0.012005f
C311 VN.n23 GND 0.012005f
C312 VN.n24 GND 0.023838f
C313 VN.n25 GND 0.017293f
C314 VN.n26 GND 0.227941f
C315 VN.n27 GND 0.392505f
C316 VN.n28 GND 0.555641f
C317 VN.t1 GND 0.020725f
C318 VN.t2 GND 0.003701f
C319 VN.t0 GND 0.003701f
C320 VN.n29 GND 0.012003f
C321 VN.n30 GND 0.112759f
C322 VN.n31 GND 1.50307f
C323 a_n1816_n673.n0 GND 0.026598f
C324 a_n1816_n673.n1 GND 0.013462f
C325 a_n1816_n673.n2 GND 0.026598f
C326 a_n1816_n673.n3 GND 0.013462f
C327 a_n1816_n673.n4 GND 0.042474f
C328 a_n1816_n673.n5 GND 0.005766f
C329 a_n1816_n673.n6 GND 0.013048f
C330 a_n1816_n673.n7 GND 0.042474f
C331 a_n1816_n673.n8 GND 0.005766f
C332 a_n1816_n673.n9 GND 0.013048f
C333 a_n1816_n673.n10 GND 0.042474f
C334 a_n1816_n673.n11 GND 0.005766f
C335 a_n1816_n673.n12 GND 0.013048f
C336 a_n1816_n673.n13 GND 0.026598f
C337 a_n1816_n673.n14 GND 0.013462f
C338 a_n1816_n673.n15 GND 0.026598f
C339 a_n1816_n673.n16 GND 0.013462f
C340 a_n1816_n673.n17 GND 0.282168f
C341 a_n1816_n673.n18 GND 0.055346f
C342 a_n1816_n673.n19 GND 0.282168f
C343 a_n1816_n673.n20 GND 0.055346f
C344 a_n1816_n673.n21 GND 0.267832f
C345 a_n1816_n673.n22 GND 0.042582f
C346 a_n1816_n673.n23 GND 0.267832f
C347 a_n1816_n673.n24 GND 0.042582f
C348 a_n1816_n673.n25 GND 0.267832f
C349 a_n1816_n673.n26 GND 0.042582f
C350 a_n1816_n673.n27 GND 0.045213f
C351 a_n1816_n673.n28 GND 0.292302f
C352 a_n1816_n673.n29 GND 0.045213f
C353 a_n1816_n673.n30 GND 0.292302f
C354 a_n1816_n673.t9 GND 0.05181f
C355 a_n1816_n673.n31 GND 0.638579f
C356 a_n1816_n673.n32 GND 0.013696f
C357 a_n1816_n673.n33 GND 0.005445f
C358 a_n1816_n673.n34 GND 0.012871f
C359 a_n1816_n673.n35 GND 0.005766f
C360 a_n1816_n673.n36 GND 0.005445f
C361 a_n1816_n673.n37 GND 0.012871f
C362 a_n1816_n673.t0 GND 0.021629f
C363 a_n1816_n673.n38 GND 0.009653f
C364 a_n1816_n673.n39 GND 0.005445f
C365 a_n1816_n673.n40 GND 0.005766f
C366 a_n1816_n673.n41 GND 0.012871f
C367 a_n1816_n673.n42 GND 0.012871f
C368 a_n1816_n673.n43 GND 0.005766f
C369 a_n1816_n673.n44 GND 0.005445f
C370 a_n1816_n673.n45 GND 0.005445f
C371 a_n1816_n673.n46 GND 0.005766f
C372 a_n1816_n673.n47 GND 0.012871f
C373 a_n1816_n673.n48 GND 0.026895f
C374 a_n1816_n673.n49 GND 0.005766f
C375 a_n1816_n673.n50 GND 0.005445f
C376 a_n1816_n673.n51 GND 0.059204f
C377 a_n1816_n673.n52 GND 0.379744f
C378 a_n1816_n673.n53 GND 0.013696f
C379 a_n1816_n673.n54 GND 0.005445f
C380 a_n1816_n673.n55 GND 0.012871f
C381 a_n1816_n673.n56 GND 0.005766f
C382 a_n1816_n673.n57 GND 0.005445f
C383 a_n1816_n673.n58 GND 0.012871f
C384 a_n1816_n673.t11 GND 0.021629f
C385 a_n1816_n673.n59 GND 0.009653f
C386 a_n1816_n673.n60 GND 0.005445f
C387 a_n1816_n673.n61 GND 0.005766f
C388 a_n1816_n673.n62 GND 0.012871f
C389 a_n1816_n673.n63 GND 0.012871f
C390 a_n1816_n673.n64 GND 0.005766f
C391 a_n1816_n673.n65 GND 0.005445f
C392 a_n1816_n673.n66 GND 0.005445f
C393 a_n1816_n673.n67 GND 0.005766f
C394 a_n1816_n673.n68 GND 0.012871f
C395 a_n1816_n673.n69 GND 0.026895f
C396 a_n1816_n673.n70 GND 0.005766f
C397 a_n1816_n673.n71 GND 0.005445f
C398 a_n1816_n673.n72 GND 0.059204f
C399 a_n1816_n673.n73 GND 0.34326f
C400 a_n1816_n673.n74 GND 0.013696f
C401 a_n1816_n673.n75 GND 0.005445f
C402 a_n1816_n673.n76 GND 0.012871f
C403 a_n1816_n673.n77 GND 0.005766f
C404 a_n1816_n673.n78 GND 0.005445f
C405 a_n1816_n673.n79 GND 0.012871f
C406 a_n1816_n673.t3 GND 0.021629f
C407 a_n1816_n673.n80 GND 0.009653f
C408 a_n1816_n673.n81 GND 0.005445f
C409 a_n1816_n673.n82 GND 0.005766f
C410 a_n1816_n673.n83 GND 0.012871f
C411 a_n1816_n673.n84 GND 0.012871f
C412 a_n1816_n673.n85 GND 0.005766f
C413 a_n1816_n673.n86 GND 0.005445f
C414 a_n1816_n673.n87 GND 0.005445f
C415 a_n1816_n673.n88 GND 0.005766f
C416 a_n1816_n673.n89 GND 0.012871f
C417 a_n1816_n673.n90 GND 0.026895f
C418 a_n1816_n673.n91 GND 0.005766f
C419 a_n1816_n673.n92 GND 0.005445f
C420 a_n1816_n673.n93 GND 0.059204f
C421 a_n1816_n673.n94 GND 0.507247f
C422 a_n1816_n673.t12 GND 0.05181f
C423 a_n1816_n673.t13 GND 0.05181f
C424 a_n1816_n673.n95 GND 0.41486f
C425 a_n1816_n673.n96 GND 0.339674f
C426 a_n1816_n673.n97 GND 0.025846f
C427 a_n1816_n673.n98 GND 0.005766f
C428 a_n1816_n673.n99 GND 0.005445f
C429 a_n1816_n673.n100 GND 0.012871f
C430 a_n1816_n673.n101 GND 0.005766f
C431 a_n1816_n673.n102 GND 0.005445f
C432 a_n1816_n673.n103 GND 0.009653f
C433 a_n1816_n673.n104 GND 0.009098f
C434 a_n1816_n673.t4 GND 0.021459f
C435 a_n1816_n673.n105 GND 0.051588f
C436 a_n1816_n673.n106 GND 0.005445f
C437 a_n1816_n673.n107 GND 0.005766f
C438 a_n1816_n673.n108 GND 0.012871f
C439 a_n1816_n673.n109 GND 0.012871f
C440 a_n1816_n673.n110 GND 0.005766f
C441 a_n1816_n673.n111 GND 0.005445f
C442 a_n1816_n673.n112 GND 0.005445f
C443 a_n1816_n673.n113 GND 0.005766f
C444 a_n1816_n673.n114 GND 0.012871f
C445 a_n1816_n673.n115 GND 0.012871f
C446 a_n1816_n673.n116 GND 0.005766f
C447 a_n1816_n673.n117 GND 0.005445f
C448 a_n1816_n673.n118 GND 0.010097f
C449 a_n1816_n673.n119 GND 0.141656f
C450 a_n1816_n673.t5 GND 0.05181f
C451 a_n1816_n673.t8 GND 0.05181f
C452 a_n1816_n673.n120 GND 0.41486f
C453 a_n1816_n673.n121 GND 0.222431f
C454 a_n1816_n673.n122 GND 0.025846f
C455 a_n1816_n673.n123 GND 0.005766f
C456 a_n1816_n673.n124 GND 0.005445f
C457 a_n1816_n673.n125 GND 0.012871f
C458 a_n1816_n673.n126 GND 0.005766f
C459 a_n1816_n673.n127 GND 0.005445f
C460 a_n1816_n673.n128 GND 0.009653f
C461 a_n1816_n673.n129 GND 0.009098f
C462 a_n1816_n673.t7 GND 0.021459f
C463 a_n1816_n673.n130 GND 0.051588f
C464 a_n1816_n673.n131 GND 0.005445f
C465 a_n1816_n673.n132 GND 0.005766f
C466 a_n1816_n673.n133 GND 0.012871f
C467 a_n1816_n673.n134 GND 0.012871f
C468 a_n1816_n673.n135 GND 0.005766f
C469 a_n1816_n673.n136 GND 0.005445f
C470 a_n1816_n673.n137 GND 0.005445f
C471 a_n1816_n673.n138 GND 0.005766f
C472 a_n1816_n673.n139 GND 0.012871f
C473 a_n1816_n673.n140 GND 0.012871f
C474 a_n1816_n673.n141 GND 0.005766f
C475 a_n1816_n673.n142 GND 0.005445f
C476 a_n1816_n673.n143 GND 0.010097f
C477 a_n1816_n673.n144 GND 0.205446f
C478 a_n1816_n673.n145 GND 0.697452f
C479 a_n1816_n673.n146 GND 0.025846f
C480 a_n1816_n673.n147 GND 0.005766f
C481 a_n1816_n673.n148 GND 0.005445f
C482 a_n1816_n673.n149 GND 0.012871f
C483 a_n1816_n673.n150 GND 0.005766f
C484 a_n1816_n673.n151 GND 0.005445f
C485 a_n1816_n673.n152 GND 0.009653f
C486 a_n1816_n673.n153 GND 0.009098f
C487 a_n1816_n673.t2 GND 0.021459f
C488 a_n1816_n673.n154 GND 0.051588f
C489 a_n1816_n673.n155 GND 0.005445f
C490 a_n1816_n673.n156 GND 0.005766f
C491 a_n1816_n673.n157 GND 0.012871f
C492 a_n1816_n673.n158 GND 0.012871f
C493 a_n1816_n673.n159 GND 0.005766f
C494 a_n1816_n673.n160 GND 0.005445f
C495 a_n1816_n673.n161 GND 0.005445f
C496 a_n1816_n673.n162 GND 0.005766f
C497 a_n1816_n673.n163 GND 0.012871f
C498 a_n1816_n673.n164 GND 0.012871f
C499 a_n1816_n673.n165 GND 0.005766f
C500 a_n1816_n673.n166 GND 0.005445f
C501 a_n1816_n673.n167 GND 0.010097f
C502 a_n1816_n673.n168 GND 0.360149f
C503 a_n1816_n673.t1 GND 0.05181f
C504 a_n1816_n673.t14 GND 0.05181f
C505 a_n1816_n673.n169 GND 0.414859f
C506 a_n1816_n673.n170 GND 0.222431f
C507 a_n1816_n673.n171 GND 0.025846f
C508 a_n1816_n673.n172 GND 0.005766f
C509 a_n1816_n673.n173 GND 0.005445f
C510 a_n1816_n673.n174 GND 0.012871f
C511 a_n1816_n673.n175 GND 0.005766f
C512 a_n1816_n673.n176 GND 0.005445f
C513 a_n1816_n673.n177 GND 0.009653f
C514 a_n1816_n673.n178 GND 0.009098f
C515 a_n1816_n673.t6 GND 0.021459f
C516 a_n1816_n673.n179 GND 0.051588f
C517 a_n1816_n673.n180 GND 0.005445f
C518 a_n1816_n673.n181 GND 0.005766f
C519 a_n1816_n673.n182 GND 0.012871f
C520 a_n1816_n673.n183 GND 0.012871f
C521 a_n1816_n673.n184 GND 0.005766f
C522 a_n1816_n673.n185 GND 0.005445f
C523 a_n1816_n673.n186 GND 0.005445f
C524 a_n1816_n673.n187 GND 0.005766f
C525 a_n1816_n673.n188 GND 0.012871f
C526 a_n1816_n673.n189 GND 0.012871f
C527 a_n1816_n673.n190 GND 0.005766f
C528 a_n1816_n673.n191 GND 0.005445f
C529 a_n1816_n673.n192 GND 0.010097f
C530 a_n1816_n673.n193 GND 0.141656f
C531 a_n1816_n673.n194 GND 0.49272f
C532 a_n1816_n673.n195 GND 0.414859f
C533 a_n1816_n673.t10 GND 0.05181f
C534 VP.n0 GND 0.024517f
C535 VP.t6 GND 0.780352f
C536 VP.n1 GND 0.018453f
C537 VP.n2 GND 0.176725f
C538 VP.t5 GND 0.780352f
C539 VP.t8 GND 0.922262f
C540 VP.n3 GND 0.32831f
C541 VP.n4 GND 0.353096f
C542 VP.n5 GND 0.034659f
C543 VP.n6 GND 0.033578f
C544 VP.n7 GND 0.018596f
C545 VP.n8 GND 0.018596f
C546 VP.n9 GND 0.018596f
C547 VP.n10 GND 0.036926f
C548 VP.n11 GND 0.026788f
C549 VP.n12 GND 0.353083f
C550 VP.n13 GND 0.259638f
C551 VP.n14 GND 0.024517f
C552 VP.t4 GND 0.780352f
C553 VP.n15 GND 0.018453f
C554 VP.n16 GND 0.176725f
C555 VP.t3 GND 0.780352f
C556 VP.t7 GND 0.922262f
C557 VP.n17 GND 0.32831f
C558 VP.n18 GND 0.353096f
C559 VP.n19 GND 0.034659f
C560 VP.n20 GND 0.033578f
C561 VP.n21 GND 0.018596f
C562 VP.n22 GND 0.018596f
C563 VP.n23 GND 0.018596f
C564 VP.n24 GND 0.036926f
C565 VP.n25 GND 0.026788f
C566 VP.n26 GND 0.353083f
C567 VP.n27 GND 0.615393f
C568 VP.n28 GND 0.868294f
C569 VP.t0 GND 0.005733f
C570 VP.t2 GND 0.005733f
C571 VP.n29 GND 0.01885f
C572 VP.t1 GND 0.031907f
C573 VP.n30 GND 0.167257f
C574 VP.n31 GND 1.34703f
C575 a_n5586_9514.n0 GND 0.858862f
C576 a_n5586_9514.t3 GND 0.456993f
C577 a_n5586_9514.t6 GND 0.057468f
C578 a_n5586_9514.t5 GND 0.057468f
C579 a_n5586_9514.n1 GND 0.318651f
C580 a_n5586_9514.n2 GND 0.88352f
C581 a_n5586_9514.t9 GND 0.647459f
C582 a_n5586_9514.t8 GND 0.808438f
C583 a_n5586_9514.n3 GND 3.95972f
C584 a_n5586_9514.t1 GND 0.445791f
C585 a_n5586_9514.n4 GND 0.58941f
C586 a_n5586_9514.t2 GND 0.057468f
C587 a_n5586_9514.t0 GND 0.057468f
C588 a_n5586_9514.n5 GND 0.318651f
C589 a_n5586_9514.n6 GND 0.491047f
C590 a_n5586_9514.t4 GND 0.445791f
C591 a_n5586_9514.t7 GND 0.445791f
C592 a_n2040_7754.n0 GND 0.539339f
C593 a_n2040_7754.t0 GND 31.4708f
C594 a_n2040_7754.t9 GND 0.36854f
C595 a_n2040_7754.n1 GND 2.31657f
C596 a_n2040_7754.t10 GND 0.500768f
C597 a_n2040_7754.n2 GND 1.49935f
C598 a_n2040_7754.t7 GND 0.279943f
C599 a_n2040_7754.n3 GND 0.370131f
C600 a_n2040_7754.t5 GND 0.036088f
C601 a_n2040_7754.t2 GND 0.036088f
C602 a_n2040_7754.n4 GND 0.200103f
C603 a_n2040_7754.n5 GND 0.308363f
C604 a_n2040_7754.t6 GND 0.286978f
C605 a_n2040_7754.t4 GND 0.036088f
C606 a_n2040_7754.t1 GND 0.036088f
C607 a_n2040_7754.n6 GND 0.200103f
C608 a_n2040_7754.n7 GND 0.554823f
C609 a_n2040_7754.t3 GND 0.279943f
C610 a_n2040_7754.t8 GND 0.279943f
C611 CS_BIAS.t11 GND 0.144704f
C612 CS_BIAS.n0 GND 0.080302f
C613 CS_BIAS.n1 GND 0.004641f
C614 CS_BIAS.n2 GND 0.00865f
C615 CS_BIAS.t6 GND 0.219205f
C616 CS_BIAS.t2 GND 0.214449f
C617 CS_BIAS.n3 GND 0.248811f
C618 CS_BIAS.t3 GND 0.003706f
C619 CS_BIAS.t7 GND 0.003706f
C620 CS_BIAS.n4 GND 0.026378f
C621 CS_BIAS.n5 GND 0.065559f
C622 CS_BIAS.n6 GND 0.094397f
C623 CS_BIAS.t15 GND 0.20525f
C624 CS_BIAS.n7 GND 0.055586f
C625 CS_BIAS.n8 GND 0.014216f
C626 CS_BIAS.n9 GND 0.004055f
C627 CS_BIAS.n10 GND 0.004641f
C628 CS_BIAS.n11 GND 0.004641f
C629 CS_BIAS.n12 GND 0.00865f
C630 CS_BIAS.n13 GND 0.00865f
C631 CS_BIAS.n14 GND 0.007625f
C632 CS_BIAS.n15 GND 0.009821f
C633 CS_BIAS.n16 GND 0.048007f
C634 CS_BIAS.t8 GND 0.219205f
C635 CS_BIAS.t12 GND 0.214449f
C636 CS_BIAS.n17 GND 0.22352f
C637 CS_BIAS.n18 GND 0.21803f
C638 CS_BIAS.t9 GND 0.144704f
C639 CS_BIAS.n19 GND 0.080302f
C640 CS_BIAS.n20 GND 0.004641f
C641 CS_BIAS.n21 GND 0.00865f
C642 CS_BIAS.t1 GND 0.003706f
C643 CS_BIAS.t5 GND 0.003706f
C644 CS_BIAS.n22 GND 0.026378f
C645 CS_BIAS.t4 GND 0.214449f
C646 CS_BIAS.t0 GND 0.219205f
C647 CS_BIAS.n23 GND 0.248811f
C648 CS_BIAS.n24 GND 0.065559f
C649 CS_BIAS.n25 GND 0.094397f
C650 CS_BIAS.t13 GND 0.205251f
C651 CS_BIAS.n26 GND 0.055586f
C652 CS_BIAS.n27 GND 0.014216f
C653 CS_BIAS.n28 GND 0.004055f
C654 CS_BIAS.n29 GND 0.004641f
C655 CS_BIAS.n30 GND 0.004641f
C656 CS_BIAS.n31 GND 0.00865f
C657 CS_BIAS.n32 GND 0.00865f
C658 CS_BIAS.n33 GND 0.007625f
C659 CS_BIAS.n34 GND 0.009821f
C660 CS_BIAS.n35 GND 0.048007f
C661 CS_BIAS.t10 GND 0.214449f
C662 CS_BIAS.t14 GND 0.219205f
C663 CS_BIAS.n36 GND 0.22352f
C664 CS_BIAS.n37 GND 0.124016f
C665 CS_BIAS.n38 GND 2.49715f
C666 VOUT.t39 GND 0.017634f
C667 VOUT.t6 GND 0.017634f
C668 VOUT.n0 GND 0.099644f
C669 VOUT.t11 GND 0.017634f
C670 VOUT.t18 GND 0.017634f
C671 VOUT.n1 GND 0.096857f
C672 VOUT.n2 GND 0.327978f
C673 VOUT.t34 GND 0.136207f
C674 VOUT.n3 GND 0.192181f
C675 VOUT.t12 GND 0.017634f
C676 VOUT.t17 GND 0.017634f
C677 VOUT.n4 GND 0.099644f
C678 VOUT.t22 GND 0.017634f
C679 VOUT.t30 GND 0.017634f
C680 VOUT.n5 GND 0.096857f
C681 VOUT.n6 GND 0.327978f
C682 VOUT.t43 GND 0.136207f
C683 VOUT.n7 GND 0.172701f
C684 VOUT.n8 GND 0.149331f
C685 VOUT.t14 GND 0.017634f
C686 VOUT.t44 GND 0.017634f
C687 VOUT.n9 GND 0.099644f
C688 VOUT.t25 GND 0.017634f
C689 VOUT.t23 GND 0.017634f
C690 VOUT.n10 GND 0.096857f
C691 VOUT.n11 GND 0.327978f
C692 VOUT.t5 GND 0.136207f
C693 VOUT.n12 GND 0.172701f
C694 VOUT.n13 GND 0.107608f
C695 VOUT.t37 GND 0.017634f
C696 VOUT.t31 GND 0.017634f
C697 VOUT.n14 GND 0.099644f
C698 VOUT.t13 GND 0.017634f
C699 VOUT.t7 GND 0.017634f
C700 VOUT.n15 GND 0.096857f
C701 VOUT.n16 GND 0.327978f
C702 VOUT.t33 GND 0.136207f
C703 VOUT.n17 GND 0.172701f
C704 VOUT.n18 GND 0.212042f
C705 VOUT.n19 GND 5.93891f
C706 VOUT.n20 GND 1.13521f
C707 VOUT.n21 GND 0.829208f
C708 VOUT.t51 GND 2.58989f
C709 VOUT.t50 GND 2.52537f
C710 VOUT.t48 GND 2.59424f
C711 VOUT.n22 GND 2.18311f
C712 VOUT.n23 GND 1.08754f
C713 VOUT.n24 GND 0.829208f
C714 VOUT.n25 GND 1.02965f
C715 VOUT.n26 GND 2.47205f
C716 VOUT.t52 GND 2.58989f
C717 VOUT.n27 GND 2.63422f
C718 VOUT.n28 GND 1.00924f
C719 VOUT.t53 GND 2.52537f
C720 VOUT.n29 GND 1.02187f
C721 VOUT.n30 GND 0.903885f
C722 VOUT.t49 GND 2.52537f
C723 VOUT.n31 GND 2.3922f
C724 VOUT.n32 GND 1.67477f
C725 VOUT.t16 GND 0.138335f
C726 VOUT.t9 GND 0.017634f
C727 VOUT.t26 GND 0.017634f
C728 VOUT.n33 GND 0.096857f
C729 VOUT.n34 GND 0.298389f
C730 VOUT.t20 GND 0.017634f
C731 VOUT.t29 GND 0.017634f
C732 VOUT.n35 GND 0.096857f
C733 VOUT.n36 GND 0.21365f
C734 VOUT.t27 GND 0.138335f
C735 VOUT.t21 GND 0.017634f
C736 VOUT.t38 GND 0.017634f
C737 VOUT.n37 GND 0.096857f
C738 VOUT.n38 GND 0.298389f
C739 VOUT.t32 GND 0.017634f
C740 VOUT.t41 GND 0.017634f
C741 VOUT.n39 GND 0.096857f
C742 VOUT.n40 GND 0.193781f
C743 VOUT.n41 GND 0.167282f
C744 VOUT.t24 GND 0.138335f
C745 VOUT.t35 GND 0.017634f
C746 VOUT.t42 GND 0.017634f
C747 VOUT.n42 GND 0.096857f
C748 VOUT.n43 GND 0.298389f
C749 VOUT.t8 GND 0.017634f
C750 VOUT.t15 GND 0.017634f
C751 VOUT.n44 GND 0.096857f
C752 VOUT.n45 GND 0.193781f
C753 VOUT.n46 GND 0.116778f
C754 VOUT.t10 GND 0.138335f
C755 VOUT.t19 GND 0.017634f
C756 VOUT.t28 GND 0.017634f
C757 VOUT.n47 GND 0.096857f
C758 VOUT.n48 GND 0.298389f
C759 VOUT.t36 GND 0.017634f
C760 VOUT.t40 GND 0.017634f
C761 VOUT.n49 GND 0.096857f
C762 VOUT.n50 GND 0.193781f
C763 VOUT.n51 GND 0.221212f
C764 VOUT.n52 GND 8.20988f
C765 VOUT.t46 GND 0.012277f
C766 VOUT.t4 GND 0.012277f
C767 VOUT.n53 GND 0.112326f
C768 VOUT.t2 GND 0.012277f
C769 VOUT.t47 GND 0.012277f
C770 VOUT.n54 GND 0.106242f
C771 VOUT.n55 GND 0.795291f
C772 VOUT.n56 GND 7.77987f
C773 VOUT.t3 GND 0.012277f
C774 VOUT.t1 GND 0.012277f
C775 VOUT.n57 GND 0.112326f
C776 VOUT.t45 GND 0.012277f
C777 VOUT.t0 GND 0.012277f
C778 VOUT.n58 GND 0.106242f
C779 VOUT.n59 GND 0.795291f
C780 VOUT.n60 GND 5.2838f
C781 VOUT.n61 GND 4.83139f
C782 VDD.t139 GND 0.005427f
C783 VDD.t120 GND 0.005427f
C784 VDD.n0 GND 0.035266f
C785 VDD.t104 GND 0.005427f
C786 VDD.t163 GND 0.005427f
C787 VDD.n1 GND 0.034145f
C788 VDD.n2 GND 0.090794f
C789 VDD.t112 GND 0.005427f
C790 VDD.t118 GND 0.005427f
C791 VDD.n3 GND 0.034145f
C792 VDD.n4 GND 0.047173f
C793 VDD.t93 GND 0.005427f
C794 VDD.t133 GND 0.005427f
C795 VDD.n5 GND 0.034145f
C796 VDD.n6 GND 0.041671f
C797 VDD.t85 GND 0.005427f
C798 VDD.t106 GND 0.005427f
C799 VDD.n7 GND 0.035266f
C800 VDD.t145 GND 0.005427f
C801 VDD.t128 GND 0.005427f
C802 VDD.n8 GND 0.034145f
C803 VDD.n9 GND 0.090794f
C804 VDD.t148 GND 0.005427f
C805 VDD.t160 GND 0.005427f
C806 VDD.n10 GND 0.034145f
C807 VDD.n11 GND 0.047173f
C808 VDD.t137 GND 0.005427f
C809 VDD.t153 GND 0.005427f
C810 VDD.n12 GND 0.034145f
C811 VDD.n13 GND 0.041671f
C812 VDD.n14 GND 0.027727f
C813 VDD.n15 GND 0.75704f
C814 VDD.t113 GND 0.004038f
C815 VDD.t95 GND 0.004038f
C816 VDD.n16 GND 0.019756f
C817 VDD.t131 GND 0.004038f
C818 VDD.t122 GND 0.004038f
C819 VDD.n17 GND 0.018989f
C820 VDD.n18 GND 0.077617f
C821 VDD.t141 GND 0.02795f
C822 VDD.n19 GND 0.041571f
C823 VDD.t134 GND 0.004038f
C824 VDD.t123 GND 0.004038f
C825 VDD.n20 GND 0.019756f
C826 VDD.t155 GND 0.004038f
C827 VDD.t140 GND 0.004038f
C828 VDD.n21 GND 0.018989f
C829 VDD.n22 GND 0.077617f
C830 VDD.t158 GND 0.02795f
C831 VDD.n23 GND 0.037037f
C832 VDD.n24 GND 0.032724f
C833 VDD.t126 GND 0.004038f
C834 VDD.t150 GND 0.004038f
C835 VDD.n25 GND 0.019756f
C836 VDD.t161 GND 0.004038f
C837 VDD.t91 GND 0.004038f
C838 VDD.n26 GND 0.018989f
C839 VDD.n27 GND 0.077617f
C840 VDD.t109 GND 0.02795f
C841 VDD.n28 GND 0.037037f
C842 VDD.n29 GND 0.023942f
C843 VDD.t97 GND 0.004038f
C844 VDD.t116 GND 0.004038f
C845 VDD.n30 GND 0.019756f
C846 VDD.t135 GND 0.004038f
C847 VDD.t151 GND 0.004038f
C848 VDD.n31 GND 0.018989f
C849 VDD.n32 GND 0.077617f
C850 VDD.t157 GND 0.02795f
C851 VDD.n33 GND 0.037037f
C852 VDD.n34 GND 0.047543f
C853 VDD.n35 GND 0.002073f
C854 VDD.n36 GND 0.002697f
C855 VDD.n37 GND 0.002171f
C856 VDD.n38 GND 0.002171f
C857 VDD.n39 GND 0.002697f
C858 VDD.n40 GND 0.002697f
C859 VDD.t130 GND 0.088808f
C860 VDD.n41 GND 0.002697f
C861 VDD.n42 GND 0.002697f
C862 VDD.n43 GND 0.002697f
C863 VDD.n44 GND 0.177615f
C864 VDD.n45 GND 0.002697f
C865 VDD.n46 GND 0.002697f
C866 VDD.n47 GND 0.002697f
C867 VDD.n48 GND 0.002697f
C868 VDD.n49 GND 0.002171f
C869 VDD.n50 GND 0.002697f
C870 VDD.n51 GND 0.002697f
C871 VDD.n52 GND 0.002697f
C872 VDD.n53 GND 0.002697f
C873 VDD.n54 GND 0.177615f
C874 VDD.n55 GND 0.002697f
C875 VDD.n56 GND 0.002697f
C876 VDD.n57 GND 0.002697f
C877 VDD.n58 GND 0.002697f
C878 VDD.n59 GND 0.002697f
C879 VDD.n60 GND 0.002171f
C880 VDD.n61 GND 0.002697f
C881 VDD.n62 GND 0.002697f
C882 VDD.n63 GND 0.002697f
C883 VDD.n64 GND 0.002697f
C884 VDD.n65 GND 0.177615f
C885 VDD.n66 GND 0.002697f
C886 VDD.n67 GND 0.002697f
C887 VDD.n68 GND 0.002697f
C888 VDD.n69 GND 0.002697f
C889 VDD.n70 GND 0.002697f
C890 VDD.n71 GND 0.002171f
C891 VDD.n72 GND 0.002697f
C892 VDD.n73 GND 0.002697f
C893 VDD.n74 GND 0.002697f
C894 VDD.n75 GND 0.002697f
C895 VDD.n76 GND 0.152749f
C896 VDD.n77 GND 0.002697f
C897 VDD.n78 GND 0.002697f
C898 VDD.n79 GND 0.002697f
C899 VDD.n80 GND 0.002697f
C900 VDD.n81 GND 0.002697f
C901 VDD.n82 GND 0.002171f
C902 VDD.n83 GND 0.002697f
C903 VDD.t25 GND 0.088808f
C904 VDD.n84 GND 0.002697f
C905 VDD.n85 GND 0.002697f
C906 VDD.n86 GND 0.006442f
C907 VDD.n87 GND 0.422724f
C908 VDD.n88 GND 0.006612f
C909 VDD.n89 GND 0.002697f
C910 VDD.n90 GND 0.002697f
C911 VDD.n91 GND 0.002697f
C912 VDD.n92 GND 0.002697f
C913 VDD.n93 GND 0.002171f
C914 VDD.n95 GND 0.002697f
C915 VDD.n96 GND 0.002697f
C916 VDD.n97 GND 0.002697f
C917 VDD.n98 GND 0.002697f
C918 VDD.n99 GND 0.002697f
C919 VDD.n100 GND 0.002171f
C920 VDD.n102 GND 0.002697f
C921 VDD.n103 GND 0.002697f
C922 VDD.n104 GND 0.002697f
C923 VDD.n105 GND 0.002697f
C924 VDD.n106 GND 0.002697f
C925 VDD.n107 GND 0.002171f
C926 VDD.n109 GND 0.002697f
C927 VDD.n110 GND 0.002697f
C928 VDD.n111 GND 0.002697f
C929 VDD.n112 GND 0.002697f
C930 VDD.n113 GND 0.002697f
C931 VDD.n114 GND 0.002171f
C932 VDD.n116 GND 0.002697f
C933 VDD.n117 GND 0.002697f
C934 VDD.n118 GND 0.002697f
C935 VDD.n119 GND 0.002697f
C936 VDD.n120 GND 0.002697f
C937 VDD.n121 GND 0.002171f
C938 VDD.n123 GND 0.002697f
C939 VDD.n124 GND 0.002697f
C940 VDD.n125 GND 0.002697f
C941 VDD.n126 GND 0.002697f
C942 VDD.n127 GND 0.002697f
C943 VDD.n128 GND 0.002171f
C944 VDD.n130 GND 0.002697f
C945 VDD.n131 GND 0.002697f
C946 VDD.n132 GND 0.002697f
C947 VDD.n133 GND 0.002697f
C948 VDD.n134 GND 0.002697f
C949 VDD.n135 GND 0.002171f
C950 VDD.n137 GND 0.002697f
C951 VDD.n138 GND 0.002697f
C952 VDD.n139 GND 0.002697f
C953 VDD.n140 GND 0.002697f
C954 VDD.n141 GND 0.002697f
C955 VDD.n142 GND 0.002171f
C956 VDD.n144 GND 0.002697f
C957 VDD.n145 GND 0.002697f
C958 VDD.n146 GND 0.002697f
C959 VDD.n147 GND 0.002697f
C960 VDD.n148 GND 0.002697f
C961 VDD.n149 GND 0.002171f
C962 VDD.n151 GND 0.002697f
C963 VDD.n152 GND 0.002697f
C964 VDD.n153 GND 0.002697f
C965 VDD.n154 GND 0.002697f
C966 VDD.n155 GND 0.002697f
C967 VDD.n156 GND 0.002171f
C968 VDD.n158 GND 0.002697f
C969 VDD.n159 GND 0.002697f
C970 VDD.n160 GND 0.002697f
C971 VDD.n161 GND 0.002697f
C972 VDD.n162 GND 0.002697f
C973 VDD.n163 GND 0.002171f
C974 VDD.n165 GND 0.002697f
C975 VDD.n166 GND 0.002697f
C976 VDD.n167 GND 0.002697f
C977 VDD.n169 GND 0.006612f
C978 VDD.n170 GND 0.001096f
C979 VDD.t74 GND 0.024975f
C980 VDD.t73 GND 0.028713f
C981 VDD.t72 GND 0.09359f
C982 VDD.n171 GND 0.022187f
C983 VDD.n172 GND 0.015995f
C984 VDD.n173 GND 0.002697f
C985 VDD.n174 GND 0.002697f
C986 VDD.n175 GND 0.002171f
C987 VDD.n176 GND 0.002697f
C988 VDD.n177 GND 0.002697f
C989 VDD.n178 GND 0.002171f
C990 VDD.n179 GND 0.002697f
C991 VDD.n180 GND 0.002697f
C992 VDD.n181 GND 0.002171f
C993 VDD.n182 GND 0.002697f
C994 VDD.n183 GND 0.002697f
C995 VDD.n184 GND 0.002171f
C996 VDD.n185 GND 0.002697f
C997 VDD.n186 GND 0.002171f
C998 VDD.n187 GND 0.002697f
C999 VDD.n188 GND 0.002171f
C1000 VDD.n189 GND 0.002697f
C1001 VDD.n190 GND 0.002697f
C1002 VDD.n191 GND 0.177615f
C1003 VDD.n192 GND 0.133211f
C1004 VDD.n193 GND 0.002697f
C1005 VDD.n194 GND 0.002171f
C1006 VDD.n195 GND 0.002697f
C1007 VDD.n196 GND 0.002171f
C1008 VDD.n197 GND 0.002697f
C1009 VDD.n198 GND 0.104793f
C1010 VDD.n199 GND 0.002697f
C1011 VDD.n200 GND 0.002171f
C1012 VDD.n201 GND 0.002697f
C1013 VDD.n202 GND 0.002171f
C1014 VDD.n203 GND 0.002697f
C1015 VDD.n204 GND 0.177615f
C1016 VDD.t94 GND 0.088808f
C1017 VDD.n205 GND 0.002697f
C1018 VDD.n206 GND 0.002171f
C1019 VDD.n207 GND 0.002697f
C1020 VDD.n208 GND 0.002171f
C1021 VDD.n209 GND 0.002697f
C1022 VDD.n210 GND 0.165182f
C1023 VDD.n211 GND 0.002697f
C1024 VDD.n212 GND 0.002171f
C1025 VDD.n213 GND 0.002697f
C1026 VDD.n214 GND 0.002171f
C1027 VDD.n215 GND 0.002697f
C1028 VDD.n216 GND 0.177615f
C1029 VDD.t96 GND 0.088808f
C1030 VDD.n217 GND 0.002697f
C1031 VDD.n218 GND 0.002171f
C1032 VDD.n219 GND 0.002697f
C1033 VDD.n220 GND 0.002171f
C1034 VDD.n221 GND 0.002697f
C1035 VDD.n222 GND 0.177615f
C1036 VDD.n223 GND 0.002697f
C1037 VDD.n224 GND 0.002171f
C1038 VDD.n225 GND 0.002697f
C1039 VDD.n226 GND 0.002171f
C1040 VDD.n227 GND 0.002697f
C1041 VDD.n228 GND 0.177615f
C1042 VDD.n229 GND 0.002697f
C1043 VDD.n230 GND 0.002171f
C1044 VDD.n231 GND 0.002697f
C1045 VDD.n232 GND 0.002171f
C1046 VDD.n233 GND 0.002697f
C1047 VDD.t17 GND 0.088808f
C1048 VDD.n234 GND 0.002697f
C1049 VDD.n235 GND 0.002171f
C1050 VDD.n236 GND 0.006442f
C1051 VDD.n237 GND 0.001802f
C1052 VDD.n238 GND 0.006442f
C1053 VDD.n239 GND 0.264647f
C1054 VDD.n240 GND 0.113674f
C1055 VDD.n241 GND 0.006442f
C1056 VDD.n242 GND 0.001802f
C1057 VDD.n243 GND 0.002697f
C1058 VDD.n244 GND 0.002171f
C1059 VDD.n245 GND 0.002697f
C1060 VDD.t81 GND 1.75129f
C1061 VDD.n268 GND 0.002697f
C1062 VDD.n269 GND 0.002697f
C1063 VDD.n270 GND 0.002077f
C1064 VDD.n273 GND 0.001969f
C1065 VDD.n274 GND 0.002697f
C1066 VDD.n275 GND 0.002697f
C1067 VDD.n276 GND 0.002697f
C1068 VDD.n277 GND 0.002697f
C1069 VDD.n278 GND 0.002697f
C1070 VDD.n279 GND 0.002697f
C1071 VDD.n280 GND 0.002697f
C1072 VDD.n281 GND 0.002697f
C1073 VDD.n282 GND 0.002697f
C1074 VDD.n283 GND 0.002697f
C1075 VDD.n284 GND 0.002697f
C1076 VDD.n285 GND 0.002697f
C1077 VDD.n286 GND 0.002697f
C1078 VDD.n287 GND 0.002697f
C1079 VDD.n288 GND 0.002697f
C1080 VDD.n289 GND 0.002697f
C1081 VDD.n290 GND 0.002697f
C1082 VDD.n291 GND 0.002697f
C1083 VDD.n292 GND 0.002697f
C1084 VDD.n293 GND 0.002697f
C1085 VDD.n294 GND 0.002697f
C1086 VDD.n295 GND 0.002697f
C1087 VDD.n296 GND 0.002697f
C1088 VDD.n297 GND 0.002697f
C1089 VDD.n298 GND 0.002697f
C1090 VDD.n299 GND 0.002697f
C1091 VDD.n300 GND 0.002697f
C1092 VDD.n301 GND 0.002697f
C1093 VDD.n302 GND 0.002697f
C1094 VDD.n303 GND 0.001969f
C1095 VDD.n304 GND 0.002171f
C1096 VDD.n305 GND 0.002077f
C1097 VDD.n306 GND 0.001834f
C1098 VDD.n307 GND 0.001834f
C1099 VDD.t105 GND 1.2735f
C1100 VDD.t84 GND 1.0799f
C1101 VDD.t127 GND 1.0799f
C1102 VDD.t144 GND 0.889852f
C1103 VDD.n309 GND 0.472457f
C1104 VDD.n310 GND 0.001834f
C1105 VDD.n311 GND 0.001834f
C1106 VDD.n313 GND 0.001834f
C1107 VDD.t55 GND 0.036555f
C1108 VDD.t54 GND 0.041821f
C1109 VDD.t53 GND 0.169586f
C1110 VDD.n314 GND 0.027364f
C1111 VDD.n315 GND 0.016899f
C1112 VDD.n316 GND 0.002621f
C1113 VDD.n318 GND 0.001308f
C1114 VDD.n319 GND 0.004477f
C1115 VDD.n320 GND 0.001834f
C1116 VDD.n321 GND 0.001834f
C1117 VDD.n322 GND 0.120778f
C1118 VDD.n323 GND 0.001834f
C1119 VDD.n324 GND 0.182944f
C1120 VDD.n325 GND 0.001834f
C1121 VDD.n326 GND 0.001834f
C1122 VDD.n327 GND 0.004477f
C1123 VDD.n328 GND 0.001834f
C1124 VDD.n329 GND 0.001834f
C1125 VDD.n330 GND 0.001834f
C1126 VDD.n331 GND 0.001834f
C1127 VDD.n333 GND 0.001834f
C1128 VDD.n334 GND 0.001834f
C1129 VDD.n336 GND 0.001834f
C1130 VDD.n337 GND 0.001834f
C1131 VDD.n339 GND 0.001834f
C1132 VDD.n340 GND 0.001834f
C1133 VDD.n342 GND 0.001834f
C1134 VDD.t46 GND 0.036555f
C1135 VDD.t45 GND 0.041821f
C1136 VDD.t43 GND 0.169586f
C1137 VDD.n343 GND 0.027364f
C1138 VDD.n344 GND 0.016899f
C1139 VDD.n345 GND 0.001834f
C1140 VDD.n346 GND 0.001834f
C1141 VDD.n347 GND 0.120778f
C1142 VDD.n348 GND 0.001834f
C1143 VDD.n349 GND 0.001834f
C1144 VDD.n350 GND 0.001834f
C1145 VDD.n351 GND 0.001834f
C1146 VDD.n352 GND 0.001834f
C1147 VDD.t44 GND 0.043516f
C1148 VDD.n353 GND 0.001834f
C1149 VDD.n354 GND 0.001834f
C1150 VDD.n355 GND 0.001834f
C1151 VDD.n356 GND 0.001834f
C1152 VDD.n357 GND 0.001834f
C1153 VDD.n358 GND 0.001834f
C1154 VDD.n359 GND 0.120778f
C1155 VDD.n360 GND 0.001834f
C1156 VDD.n361 GND 0.001834f
C1157 VDD.t159 GND 0.039075f
C1158 VDD.n362 GND 0.077263f
C1159 VDD.n363 GND 0.001834f
C1160 VDD.n364 GND 0.001834f
C1161 VDD.n365 GND 0.001834f
C1162 VDD.n366 GND 0.120778f
C1163 VDD.n367 GND 0.001834f
C1164 VDD.n368 GND 0.001834f
C1165 VDD.n369 GND 0.001834f
C1166 VDD.n370 GND 0.001834f
C1167 VDD.n371 GND 0.001834f
C1168 VDD.n372 GND 0.120778f
C1169 VDD.n373 GND 0.001834f
C1170 VDD.n374 GND 0.001834f
C1171 VDD.n375 GND 0.001834f
C1172 VDD.n376 GND 0.001834f
C1173 VDD.n377 GND 0.001834f
C1174 VDD.n378 GND 0.100353f
C1175 VDD.n379 GND 0.001834f
C1176 VDD.n380 GND 0.001834f
C1177 VDD.n381 GND 0.001834f
C1178 VDD.n382 GND 0.001834f
C1179 VDD.n383 GND 0.001834f
C1180 VDD.n384 GND 0.120778f
C1181 VDD.n385 GND 0.001834f
C1182 VDD.n386 GND 0.001834f
C1183 VDD.t147 GND 0.060389f
C1184 VDD.n387 GND 0.001834f
C1185 VDD.n388 GND 0.001834f
C1186 VDD.n389 GND 0.001834f
C1187 VDD.t121 GND 0.060389f
C1188 VDD.n390 GND 0.001834f
C1189 VDD.n391 GND 0.001834f
C1190 VDD.n392 GND 0.001834f
C1191 VDD.n393 GND 0.001834f
C1192 VDD.n394 GND 0.001834f
C1193 VDD.n395 GND 0.120778f
C1194 VDD.n396 GND 0.001834f
C1195 VDD.n397 GND 0.001834f
C1196 VDD.n398 GND 0.090584f
C1197 VDD.n399 GND 0.001834f
C1198 VDD.n400 GND 0.001834f
C1199 VDD.n401 GND 0.001834f
C1200 VDD.n402 GND 0.120778f
C1201 VDD.n403 GND 0.001834f
C1202 VDD.n404 GND 0.001834f
C1203 VDD.n405 GND 0.001834f
C1204 VDD.n406 GND 0.001834f
C1205 VDD.n407 GND 0.001834f
C1206 VDD.t152 GND 0.060389f
C1207 VDD.n408 GND 0.001834f
C1208 VDD.n409 GND 0.001834f
C1209 VDD.n410 GND 0.001834f
C1210 VDD.n411 GND 0.001834f
C1211 VDD.n412 GND 0.001834f
C1212 VDD.n413 GND 0.120778f
C1213 VDD.n414 GND 0.001834f
C1214 VDD.n415 GND 0.001834f
C1215 VDD.n416 GND 0.084367f
C1216 VDD.n417 GND 0.001834f
C1217 VDD.n418 GND 0.001834f
C1218 VDD.n419 GND 0.001834f
C1219 VDD.n420 GND 0.120778f
C1220 VDD.n421 GND 0.001834f
C1221 VDD.n422 GND 0.001834f
C1222 VDD.n423 GND 0.001834f
C1223 VDD.n424 GND 0.001834f
C1224 VDD.n425 GND 0.001834f
C1225 VDD.t2 GND 0.060389f
C1226 VDD.n426 GND 0.001834f
C1227 VDD.n427 GND 0.001834f
C1228 VDD.n428 GND 0.001834f
C1229 VDD.n429 GND 0.001834f
C1230 VDD.n430 GND 0.001834f
C1231 VDD.n431 GND 0.093248f
C1232 VDD.n432 GND 0.001834f
C1233 VDD.n433 GND 0.001834f
C1234 VDD.n434 GND 0.081703f
C1235 VDD.n435 GND 0.001834f
C1236 VDD.n436 GND 0.001834f
C1237 VDD.n437 GND 0.001834f
C1238 VDD.n438 GND 0.120778f
C1239 VDD.n439 GND 0.001834f
C1240 VDD.n440 GND 0.001834f
C1241 VDD.t136 GND 0.060389f
C1242 VDD.n441 GND 0.001834f
C1243 VDD.n442 GND 0.004693f
C1244 VDD.n443 GND 0.004693f
C1245 VDD.n444 GND 0.182944f
C1246 VDD.n455 GND 0.004693f
C1247 VDD.n466 GND 0.004477f
C1248 VDD.n467 GND 0.001834f
C1249 VDD.n468 GND 0.004477f
C1250 VDD.t61 GND 0.036555f
C1251 VDD.t60 GND 0.041821f
C1252 VDD.t59 GND 0.169586f
C1253 VDD.n469 GND 0.027364f
C1254 VDD.n470 GND 0.016899f
C1255 VDD.n471 GND 0.002621f
C1256 VDD.n472 GND 0.004674f
C1257 VDD.n473 GND 0.001834f
C1258 VDD.n474 GND 0.001834f
C1259 VDD.n475 GND 0.08792f
C1260 VDD.n476 GND 0.001834f
C1261 VDD.n477 GND 0.001834f
C1262 VDD.n478 GND 0.001834f
C1263 VDD.n479 GND 0.001834f
C1264 VDD.n480 GND 0.001834f
C1265 VDD.n481 GND 0.120778f
C1266 VDD.n482 GND 0.001834f
C1267 VDD.n483 GND 0.001834f
C1268 VDD.t132 GND 0.060389f
C1269 VDD.n484 GND 0.001834f
C1270 VDD.n485 GND 0.001834f
C1271 VDD.n486 GND 0.001834f
C1272 VDD.t12 GND 0.036555f
C1273 VDD.t11 GND 0.041821f
C1274 VDD.t9 GND 0.169586f
C1275 VDD.n487 GND 0.027364f
C1276 VDD.n488 GND 0.016899f
C1277 VDD.n489 GND 0.001834f
C1278 VDD.n490 GND 0.001834f
C1279 VDD.t10 GND 0.060389f
C1280 VDD.n491 GND 0.001834f
C1281 VDD.n492 GND 0.001834f
C1282 VDD.n493 GND 0.001834f
C1283 VDD.n494 GND 0.001834f
C1284 VDD.n495 GND 0.001834f
C1285 VDD.n496 GND 0.120778f
C1286 VDD.n497 GND 0.001834f
C1287 VDD.n498 GND 0.001834f
C1288 VDD.n499 GND 0.099464f
C1289 VDD.n500 GND 0.001834f
C1290 VDD.n501 GND 0.001834f
C1291 VDD.n502 GND 0.001834f
C1292 VDD.n503 GND 0.001834f
C1293 VDD.n504 GND 0.120778f
C1294 VDD.n505 GND 0.001834f
C1295 VDD.n506 GND 0.001834f
C1296 VDD.n507 GND 0.001834f
C1297 VDD.n508 GND 0.001834f
C1298 VDD.n509 GND 0.001834f
C1299 VDD.t92 GND 0.060389f
C1300 VDD.n510 GND 0.001834f
C1301 VDD.n511 GND 0.001834f
C1302 VDD.n512 GND 0.001834f
C1303 VDD.n513 GND 0.001834f
C1304 VDD.n514 GND 0.001834f
C1305 VDD.n515 GND 0.120778f
C1306 VDD.n516 GND 0.001834f
C1307 VDD.n517 GND 0.001834f
C1308 VDD.n518 GND 0.0968f
C1309 VDD.n519 GND 0.001834f
C1310 VDD.n520 GND 0.001834f
C1311 VDD.n521 GND 0.001834f
C1312 VDD.n522 GND 0.120778f
C1313 VDD.n523 GND 0.001834f
C1314 VDD.n524 GND 0.001834f
C1315 VDD.n525 GND 0.001834f
C1316 VDD.n526 GND 0.001834f
C1317 VDD.n527 GND 0.001834f
C1318 VDD.t102 GND 0.060389f
C1319 VDD.n528 GND 0.001834f
C1320 VDD.n529 GND 0.001834f
C1321 VDD.n530 GND 0.001834f
C1322 VDD.n531 GND 0.001834f
C1323 VDD.n532 GND 0.001834f
C1324 VDD.n533 GND 0.080815f
C1325 VDD.n534 GND 0.001834f
C1326 VDD.n535 GND 0.001834f
C1327 VDD.n536 GND 0.090584f
C1328 VDD.n537 GND 0.001834f
C1329 VDD.n538 GND 0.001834f
C1330 VDD.n539 GND 0.001834f
C1331 VDD.n540 GND 0.120778f
C1332 VDD.n541 GND 0.001834f
C1333 VDD.n542 GND 0.001834f
C1334 VDD.t117 GND 0.060389f
C1335 VDD.n543 GND 0.001834f
C1336 VDD.n544 GND 0.001834f
C1337 VDD.n545 GND 0.001834f
C1338 VDD.n546 GND 0.120778f
C1339 VDD.n547 GND 0.001834f
C1340 VDD.n548 GND 0.001834f
C1341 VDD.n549 GND 0.001834f
C1342 VDD.n550 GND 0.001834f
C1343 VDD.n551 GND 0.001834f
C1344 VDD.n552 GND 0.120778f
C1345 VDD.n553 GND 0.001834f
C1346 VDD.n554 GND 0.001834f
C1347 VDD.n555 GND 0.001834f
C1348 VDD.n556 GND 0.001834f
C1349 VDD.n557 GND 0.001834f
C1350 VDD.n558 GND 0.120778f
C1351 VDD.n559 GND 0.001834f
C1352 VDD.n560 GND 0.001834f
C1353 VDD.n561 GND 0.001834f
C1354 VDD.n562 GND 0.001834f
C1355 VDD.n563 GND 0.001834f
C1356 VDD.t111 GND 0.039075f
C1357 VDD.n564 GND 0.001834f
C1358 VDD.n565 GND 0.001834f
C1359 VDD.n566 GND 0.001834f
C1360 VDD.n567 GND 0.001834f
C1361 VDD.n568 GND 0.001834f
C1362 VDD.n569 GND 0.120778f
C1363 VDD.n570 GND 0.001834f
C1364 VDD.n571 GND 0.001834f
C1365 VDD.t69 GND 0.043516f
C1366 VDD.n572 GND 0.081703f
C1367 VDD.n573 GND 0.001834f
C1368 VDD.n574 GND 0.001834f
C1369 VDD.n575 GND 0.001834f
C1370 VDD.n576 GND 0.120778f
C1371 VDD.n577 GND 0.001834f
C1372 VDD.n578 GND 0.001834f
C1373 VDD.n579 GND 0.001834f
C1374 VDD.n580 GND 0.004693f
C1375 VDD.n581 GND 0.004693f
C1376 VDD.n582 GND 0.472457f
C1377 VDD.n583 GND 0.004477f
C1378 VDD.n584 GND 0.004477f
C1379 VDD.n585 GND 0.004693f
C1380 VDD.n586 GND 0.001834f
C1381 VDD.n587 GND 0.001834f
C1382 VDD.n588 GND 0.001834f
C1383 VDD.n589 GND 0.001834f
C1384 VDD.n590 GND 0.001969f
C1385 VDD.n593 GND 0.002697f
C1386 VDD.n594 GND 0.002171f
C1387 VDD.n595 GND 0.002697f
C1388 VDD.n596 GND 0.002697f
C1389 VDD.n597 GND 0.001096f
C1390 VDD.t8 GND 0.024975f
C1391 VDD.t7 GND 0.028713f
C1392 VDD.t5 GND 0.09359f
C1393 VDD.n598 GND 0.022187f
C1394 VDD.n599 GND 0.015995f
C1395 VDD.n600 GND 0.002697f
C1396 VDD.t162 GND 0.889852f
C1397 VDD.t103 GND 1.0799f
C1398 VDD.t119 GND 1.0799f
C1399 VDD.t138 GND 1.2735f
C1400 VDD.t0 GND 1.75129f
C1401 VDD.n602 GND 1.19357f
C1402 VDD.n603 GND 0.002697f
C1403 VDD.n604 GND 0.001802f
C1404 VDD.n605 GND 0.177615f
C1405 VDD.n606 GND 0.002697f
C1406 VDD.n607 GND 0.006612f
C1407 VDD.n608 GND 0.002171f
C1408 VDD.n609 GND 0.002697f
C1409 VDD.n610 GND 0.002171f
C1410 VDD.n611 GND 0.002697f
C1411 VDD.t6 GND 0.088808f
C1412 VDD.n612 GND 0.002697f
C1413 VDD.n613 GND 0.002171f
C1414 VDD.n614 GND 0.002171f
C1415 VDD.n615 GND 0.002697f
C1416 VDD.n616 GND 0.002171f
C1417 VDD.n617 GND 0.002697f
C1418 VDD.n618 GND 0.177615f
C1419 VDD.n619 GND 0.152749f
C1420 VDD.n620 GND 0.002697f
C1421 VDD.n621 GND 0.002171f
C1422 VDD.n622 GND 0.002697f
C1423 VDD.n623 GND 0.002171f
C1424 VDD.n624 GND 0.002697f
C1425 VDD.n625 GND 0.177615f
C1426 VDD.n626 GND 0.002697f
C1427 VDD.n627 GND 0.002171f
C1428 VDD.n628 GND 0.002697f
C1429 VDD.n629 GND 0.002171f
C1430 VDD.n630 GND 0.002697f
C1431 VDD.n631 GND 0.101241f
C1432 VDD.n632 GND 0.002697f
C1433 VDD.n633 GND 0.002171f
C1434 VDD.n634 GND 0.002697f
C1435 VDD.n635 GND 0.002171f
C1436 VDD.n636 GND 0.002697f
C1437 VDD.n637 GND 0.177615f
C1438 VDD.n638 GND 0.002697f
C1439 VDD.n639 GND 0.002171f
C1440 VDD.n640 GND 0.002697f
C1441 VDD.n641 GND 0.002171f
C1442 VDD.n642 GND 0.002697f
C1443 VDD.n643 GND 0.16163f
C1444 VDD.n644 GND 0.002697f
C1445 VDD.n645 GND 0.002171f
C1446 VDD.n646 GND 0.002697f
C1447 VDD.n647 GND 0.002171f
C1448 VDD.n648 GND 0.002697f
C1449 VDD.n649 GND 0.177615f
C1450 VDD.n650 GND 0.002697f
C1451 VDD.n651 GND 0.002171f
C1452 VDD.n652 GND 0.002697f
C1453 VDD.n653 GND 0.002171f
C1454 VDD.n654 GND 0.002697f
C1455 VDD.n655 GND 0.177615f
C1456 VDD.n656 GND 0.002697f
C1457 VDD.n657 GND 0.002171f
C1458 VDD.t87 GND 0.028534f
C1459 VDD.t115 GND 0.004038f
C1460 VDD.t156 GND 0.004038f
C1461 VDD.n658 GND 0.018989f
C1462 VDD.n659 GND 0.070923f
C1463 VDD.t149 GND 0.004038f
C1464 VDD.t99 GND 0.004038f
C1465 VDD.n660 GND 0.018989f
C1466 VDD.n661 GND 0.04677f
C1467 VDD.t114 GND 0.028534f
C1468 VDD.t142 GND 0.004038f
C1469 VDD.t101 GND 0.004038f
C1470 VDD.n662 GND 0.018989f
C1471 VDD.n663 GND 0.070923f
C1472 VDD.t164 GND 0.004038f
C1473 VDD.t124 GND 0.004038f
C1474 VDD.n664 GND 0.018989f
C1475 VDD.n665 GND 0.042294f
C1476 VDD.n666 GND 0.036022f
C1477 VDD.t165 GND 0.028534f
C1478 VDD.t125 GND 0.004038f
C1479 VDD.t110 GND 0.004038f
C1480 VDD.n667 GND 0.018989f
C1481 VDD.n668 GND 0.070923f
C1482 VDD.t83 GND 0.004038f
C1483 VDD.t129 GND 0.004038f
C1484 VDD.n669 GND 0.018989f
C1485 VDD.n670 GND 0.042294f
C1486 VDD.n671 GND 0.025562f
C1487 VDD.t143 GND 0.028534f
C1488 VDD.t89 GND 0.004038f
C1489 VDD.t154 GND 0.004038f
C1490 VDD.n672 GND 0.018989f
C1491 VDD.n673 GND 0.070923f
C1492 VDD.t146 GND 0.004038f
C1493 VDD.t107 GND 0.004038f
C1494 VDD.n674 GND 0.018989f
C1495 VDD.n675 GND 0.042294f
C1496 VDD.n676 GND 0.049162f
C1497 VDD.n677 GND 0.679009f
C1498 VDD.n678 GND 0.068919f
C1499 VDD.n679 GND 0.002171f
C1500 VDD.n680 GND 0.002697f
C1501 VDD.t88 GND 0.088808f
C1502 VDD.n681 GND 0.002697f
C1503 VDD.n682 GND 0.002171f
C1504 VDD.n683 GND 0.002697f
C1505 VDD.n684 GND 0.002171f
C1506 VDD.n685 GND 0.002697f
C1507 VDD.n686 GND 0.177615f
C1508 VDD.n687 GND 0.133211f
C1509 VDD.n688 GND 0.002697f
C1510 VDD.n689 GND 0.002171f
C1511 VDD.n690 GND 0.002697f
C1512 VDD.n691 GND 0.002171f
C1513 VDD.n692 GND 0.002697f
C1514 VDD.n693 GND 0.104793f
C1515 VDD.n694 GND 0.002697f
C1516 VDD.n695 GND 0.002171f
C1517 VDD.n696 GND 0.002697f
C1518 VDD.n697 GND 0.002171f
C1519 VDD.n698 GND 0.002697f
C1520 VDD.n699 GND 0.177615f
C1521 VDD.t98 GND 0.088808f
C1522 VDD.n700 GND 0.002697f
C1523 VDD.n701 GND 0.002171f
C1524 VDD.n702 GND 0.002697f
C1525 VDD.n703 GND 0.002171f
C1526 VDD.n704 GND 0.002697f
C1527 VDD.n705 GND 0.165182f
C1528 VDD.n706 GND 0.002697f
C1529 VDD.n707 GND 0.002171f
C1530 VDD.n708 GND 0.002697f
C1531 VDD.n709 GND 0.002171f
C1532 VDD.n710 GND 0.002697f
C1533 VDD.n711 GND 0.177615f
C1534 VDD.t82 GND 0.088808f
C1535 VDD.n712 GND 0.002697f
C1536 VDD.n713 GND 0.002171f
C1537 VDD.n714 GND 0.002697f
C1538 VDD.n715 GND 0.002171f
C1539 VDD.n716 GND 0.002697f
C1540 VDD.n717 GND 0.177615f
C1541 VDD.n718 GND 0.002697f
C1542 VDD.n719 GND 0.002171f
C1543 VDD.n720 GND 0.002697f
C1544 VDD.n721 GND 0.002171f
C1545 VDD.n722 GND 0.002697f
C1546 VDD.n723 GND 0.177615f
C1547 VDD.n724 GND 0.002697f
C1548 VDD.n725 GND 0.002171f
C1549 VDD.n726 GND 0.002697f
C1550 VDD.n727 GND 0.002171f
C1551 VDD.n728 GND 0.002697f
C1552 VDD.t21 GND 0.088808f
C1553 VDD.n729 GND 0.002697f
C1554 VDD.n730 GND 0.002171f
C1555 VDD.n731 GND 0.006442f
C1556 VDD.n732 GND 0.001802f
C1557 VDD.n733 GND 0.006442f
C1558 VDD.n734 GND 0.264647f
C1559 VDD.n735 GND 0.113674f
C1560 VDD.n736 GND 0.006442f
C1561 VDD.n737 GND 0.001802f
C1562 VDD.n738 GND 0.002697f
C1563 VDD.n739 GND 0.002171f
C1564 VDD.n740 GND 0.002697f
C1565 VDD.n763 GND 0.002697f
C1566 VDD.n764 GND 0.002171f
C1567 VDD.n765 GND 0.002697f
C1568 VDD.n766 GND 0.002697f
C1569 VDD.n767 GND 0.002697f
C1570 VDD.n768 GND 0.002697f
C1571 VDD.n769 GND 0.002697f
C1572 VDD.n770 GND 0.002171f
C1573 VDD.n771 GND 0.002697f
C1574 VDD.n772 GND 0.002697f
C1575 VDD.n773 GND 0.002697f
C1576 VDD.n774 GND 0.002697f
C1577 VDD.n775 GND 0.002697f
C1578 VDD.n776 GND 0.002171f
C1579 VDD.n777 GND 0.002697f
C1580 VDD.n778 GND 0.002697f
C1581 VDD.n779 GND 0.002697f
C1582 VDD.n780 GND 0.002697f
C1583 VDD.n781 GND 0.002697f
C1584 VDD.n782 GND 0.002171f
C1585 VDD.n783 GND 0.002697f
C1586 VDD.n784 GND 0.002697f
C1587 VDD.n785 GND 0.002697f
C1588 VDD.n786 GND 0.002697f
C1589 VDD.n787 GND 0.002697f
C1590 VDD.n788 GND 0.002171f
C1591 VDD.n789 GND 0.002697f
C1592 VDD.n790 GND 0.002697f
C1593 VDD.n791 GND 0.002697f
C1594 VDD.n792 GND 0.002697f
C1595 VDD.n793 GND 0.002697f
C1596 VDD.n794 GND 0.002171f
C1597 VDD.n795 GND 0.002697f
C1598 VDD.n796 GND 0.002697f
C1599 VDD.n797 GND 0.002697f
C1600 VDD.n798 GND 0.002697f
C1601 VDD.n799 GND 0.002697f
C1602 VDD.n800 GND 0.002171f
C1603 VDD.n801 GND 0.002697f
C1604 VDD.n802 GND 0.002697f
C1605 VDD.n803 GND 0.002697f
C1606 VDD.n804 GND 0.002697f
C1607 VDD.n805 GND 0.002697f
C1608 VDD.n806 GND 0.002171f
C1609 VDD.n807 GND 0.002697f
C1610 VDD.n808 GND 0.002697f
C1611 VDD.n809 GND 0.002697f
C1612 VDD.n810 GND 0.002697f
C1613 VDD.n811 GND 0.002697f
C1614 VDD.n812 GND 0.002171f
C1615 VDD.n813 GND 0.002697f
C1616 VDD.n814 GND 0.002697f
C1617 VDD.n815 GND 0.002697f
C1618 VDD.n816 GND 0.002697f
C1619 VDD.n817 GND 0.002697f
C1620 VDD.n818 GND 0.002171f
C1621 VDD.n819 GND 0.002697f
C1622 VDD.n820 GND 0.002697f
C1623 VDD.n821 GND 0.002697f
C1624 VDD.n822 GND 0.002697f
C1625 VDD.n823 GND 0.002697f
C1626 VDD.n824 GND 0.002171f
C1627 VDD.n825 GND 0.002697f
C1628 VDD.n826 GND 0.002697f
C1629 VDD.n827 GND 0.006612f
C1630 VDD.n828 GND 0.006612f
C1631 VDD.n829 GND 0.001096f
C1632 VDD.n830 GND 0.002697f
C1633 VDD.t22 GND 0.024975f
C1634 VDD.t23 GND 0.028713f
C1635 VDD.t20 GND 0.09359f
C1636 VDD.n831 GND 0.022187f
C1637 VDD.n832 GND 0.015995f
C1638 VDD.n833 GND 0.004429f
C1639 VDD.n834 GND 0.00216f
C1640 VDD.n835 GND 0.002697f
C1641 VDD.n836 GND 0.002697f
C1642 VDD.n837 GND 0.002697f
C1643 VDD.n838 GND 0.002171f
C1644 VDD.n839 GND 0.002171f
C1645 VDD.n840 GND 0.002171f
C1646 VDD.n841 GND 0.002697f
C1647 VDD.n842 GND 0.002697f
C1648 VDD.n843 GND 0.002697f
C1649 VDD.n844 GND 0.002171f
C1650 VDD.n845 GND 0.002171f
C1651 VDD.n846 GND 0.002171f
C1652 VDD.n847 GND 0.002697f
C1653 VDD.n848 GND 0.002697f
C1654 VDD.n849 GND 0.002697f
C1655 VDD.n850 GND 0.001444f
C1656 VDD.t41 GND 0.024975f
C1657 VDD.t42 GND 0.028713f
C1658 VDD.t40 GND 0.09359f
C1659 VDD.n851 GND 0.022187f
C1660 VDD.n852 GND 0.015995f
C1661 VDD.n853 GND 0.003343f
C1662 VDD.n854 GND 0.001096f
C1663 VDD.n855 GND 0.002171f
C1664 VDD.n856 GND 0.002697f
C1665 VDD.n857 GND 0.002697f
C1666 VDD.n858 GND 0.002697f
C1667 VDD.n859 GND 0.002171f
C1668 VDD.n860 GND 0.002171f
C1669 VDD.n861 GND 0.002171f
C1670 VDD.n862 GND 0.002697f
C1671 VDD.n863 GND 0.002697f
C1672 VDD.n864 GND 0.002697f
C1673 VDD.n865 GND 0.002171f
C1674 VDD.n866 GND 0.002171f
C1675 VDD.n867 GND 0.002171f
C1676 VDD.n868 GND 0.002697f
C1677 VDD.n869 GND 0.002697f
C1678 VDD.n870 GND 0.002697f
C1679 VDD.n871 GND 0.001444f
C1680 VDD.t66 GND 0.024975f
C1681 VDD.t67 GND 0.028713f
C1682 VDD.t65 GND 0.09359f
C1683 VDD.n872 GND 0.022187f
C1684 VDD.n873 GND 0.015995f
C1685 VDD.n874 GND 0.003343f
C1686 VDD.n875 GND 0.001096f
C1687 VDD.n876 GND 0.002171f
C1688 VDD.n877 GND 0.002697f
C1689 VDD.n878 GND 0.002697f
C1690 VDD.n879 GND 0.002697f
C1691 VDD.n880 GND 0.002171f
C1692 VDD.n881 GND 0.002171f
C1693 VDD.n882 GND 0.002171f
C1694 VDD.n883 GND 0.002697f
C1695 VDD.n884 GND 0.002697f
C1696 VDD.n885 GND 0.002697f
C1697 VDD.n886 GND 0.002171f
C1698 VDD.n887 GND 0.002171f
C1699 VDD.n888 GND 0.002171f
C1700 VDD.n889 GND 0.002697f
C1701 VDD.n890 GND 0.002697f
C1702 VDD.n891 GND 0.002697f
C1703 VDD.n892 GND 0.001422f
C1704 VDD.t48 GND 0.024975f
C1705 VDD.t49 GND 0.028713f
C1706 VDD.t47 GND 0.09359f
C1707 VDD.n893 GND 0.022187f
C1708 VDD.n894 GND 0.015995f
C1709 VDD.n895 GND 0.003343f
C1710 VDD.n896 GND 0.001118f
C1711 VDD.n897 GND 0.002171f
C1712 VDD.n898 GND 0.002697f
C1713 VDD.n899 GND 0.002697f
C1714 VDD.n900 GND 0.002697f
C1715 VDD.n901 GND 0.002171f
C1716 VDD.n902 GND 0.002171f
C1717 VDD.n903 GND 0.002171f
C1718 VDD.n904 GND 0.002697f
C1719 VDD.n905 GND 0.002697f
C1720 VDD.n906 GND 0.002697f
C1721 VDD.n907 GND 0.002171f
C1722 VDD.n908 GND 0.002697f
C1723 VDD.n909 GND 0.422724f
C1724 VDD.n911 GND 0.006612f
C1725 VDD.n912 GND 0.001802f
C1726 VDD.n913 GND 0.006612f
C1727 VDD.n914 GND 0.006442f
C1728 VDD.n915 GND 0.002697f
C1729 VDD.n916 GND 0.002171f
C1730 VDD.n917 GND 0.002697f
C1731 VDD.n918 GND 0.177615f
C1732 VDD.n919 GND 0.002697f
C1733 VDD.n920 GND 0.002171f
C1734 VDD.n921 GND 0.002697f
C1735 VDD.n922 GND 0.002697f
C1736 VDD.n923 GND 0.002697f
C1737 VDD.n924 GND 0.002171f
C1738 VDD.n925 GND 0.002697f
C1739 VDD.n926 GND 0.152749f
C1740 VDD.n927 GND 0.002697f
C1741 VDD.n928 GND 0.002171f
C1742 VDD.n929 GND 0.002697f
C1743 VDD.n930 GND 0.002697f
C1744 VDD.n931 GND 0.002697f
C1745 VDD.n932 GND 0.002171f
C1746 VDD.n933 GND 0.002697f
C1747 VDD.n934 GND 0.177615f
C1748 VDD.n935 GND 0.002697f
C1749 VDD.n936 GND 0.002171f
C1750 VDD.n937 GND 0.002697f
C1751 VDD.n938 GND 0.002697f
C1752 VDD.n939 GND 0.002697f
C1753 VDD.n940 GND 0.002171f
C1754 VDD.n941 GND 0.002697f
C1755 VDD.n942 GND 0.177615f
C1756 VDD.n943 GND 0.002697f
C1757 VDD.n944 GND 0.002171f
C1758 VDD.n945 GND 0.002697f
C1759 VDD.n946 GND 0.002697f
C1760 VDD.n947 GND 0.002697f
C1761 VDD.n948 GND 0.002171f
C1762 VDD.n949 GND 0.002697f
C1763 VDD.n950 GND 0.101241f
C1764 VDD.n951 GND 0.002697f
C1765 VDD.n952 GND 0.002171f
C1766 VDD.n953 GND 0.002697f
C1767 VDD.n954 GND 0.002697f
C1768 VDD.n955 GND 0.002697f
C1769 VDD.n956 GND 0.002171f
C1770 VDD.n957 GND 0.002697f
C1771 VDD.n958 GND 0.177615f
C1772 VDD.n959 GND 0.002697f
C1773 VDD.n960 GND 0.002171f
C1774 VDD.n961 GND 0.002697f
C1775 VDD.n962 GND 0.002697f
C1776 VDD.n963 GND 0.002697f
C1777 VDD.n964 GND 0.002171f
C1778 VDD.n965 GND 0.002697f
C1779 VDD.n966 GND 0.16163f
C1780 VDD.n967 GND 0.002697f
C1781 VDD.n968 GND 0.002171f
C1782 VDD.n969 GND 0.002697f
C1783 VDD.n970 GND 0.002697f
C1784 VDD.n971 GND 0.002697f
C1785 VDD.n972 GND 0.002171f
C1786 VDD.n973 GND 0.002697f
C1787 VDD.n974 GND 0.177615f
C1788 VDD.n975 GND 0.002697f
C1789 VDD.n976 GND 0.002171f
C1790 VDD.n977 GND 0.002697f
C1791 VDD.n978 GND 0.002697f
C1792 VDD.n979 GND 0.002073f
C1793 VDD.n980 GND 0.002697f
C1794 VDD.n981 GND 0.002171f
C1795 VDD.n982 GND 0.002697f
C1796 VDD.n983 GND 0.177615f
C1797 VDD.n984 GND 0.002697f
C1798 VDD.n985 GND 0.002171f
C1799 VDD.n986 GND 0.002697f
C1800 VDD.n987 GND 0.002697f
C1801 VDD.n988 GND 0.002697f
C1802 VDD.n989 GND 0.002171f
C1803 VDD.n990 GND 0.002697f
C1804 VDD.n991 GND 0.133211f
C1805 VDD.n992 GND 0.002697f
C1806 VDD.n993 GND 0.002171f
C1807 VDD.n994 GND 0.002073f
C1808 VDD.n995 GND 0.002697f
C1809 VDD.n996 GND 0.002697f
C1810 VDD.n997 GND 0.002171f
C1811 VDD.n998 GND 0.002697f
C1812 VDD.n999 GND 0.177615f
C1813 VDD.n1000 GND 0.002697f
C1814 VDD.n1001 GND 0.002171f
C1815 VDD.n1002 GND 0.002697f
C1816 VDD.n1003 GND 0.002697f
C1817 VDD.n1004 GND 0.002697f
C1818 VDD.n1005 GND 0.002171f
C1819 VDD.n1006 GND 0.002697f
C1820 VDD.t100 GND 0.088808f
C1821 VDD.n1007 GND 0.104793f
C1822 VDD.n1008 GND 0.002697f
C1823 VDD.n1009 GND 0.002171f
C1824 VDD.n1010 GND 0.002697f
C1825 VDD.n1011 GND 0.002697f
C1826 VDD.n1012 GND 0.002697f
C1827 VDD.n1013 GND 0.002171f
C1828 VDD.n1014 GND 0.002697f
C1829 VDD.n1015 GND 0.177615f
C1830 VDD.n1016 GND 0.002697f
C1831 VDD.n1017 GND 0.002171f
C1832 VDD.n1018 GND 0.002697f
C1833 VDD.n1019 GND 0.002697f
C1834 VDD.n1020 GND 0.002697f
C1835 VDD.n1021 GND 0.002171f
C1836 VDD.n1022 GND 0.002697f
C1837 VDD.t86 GND 0.088808f
C1838 VDD.n1023 GND 0.165182f
C1839 VDD.n1024 GND 0.002697f
C1840 VDD.n1025 GND 0.002171f
C1841 VDD.n1026 GND 0.002697f
C1842 VDD.n1027 GND 0.002697f
C1843 VDD.n1028 GND 0.002697f
C1844 VDD.n1029 GND 0.002171f
C1845 VDD.n1030 GND 0.002697f
C1846 VDD.n1031 GND 0.177615f
C1847 VDD.n1032 GND 0.002697f
C1848 VDD.n1033 GND 0.002171f
C1849 VDD.n1034 GND 0.002697f
C1850 VDD.n1035 GND 0.002697f
C1851 VDD.n1036 GND 0.002697f
C1852 VDD.n1037 GND 0.002171f
C1853 VDD.n1038 GND 0.002697f
C1854 VDD.n1039 GND 0.177615f
C1855 VDD.n1040 GND 0.002697f
C1856 VDD.n1041 GND 0.002171f
C1857 VDD.n1042 GND 0.002697f
C1858 VDD.n1043 GND 0.002697f
C1859 VDD.n1044 GND 0.002697f
C1860 VDD.n1045 GND 0.002171f
C1861 VDD.n1046 GND 0.002697f
C1862 VDD.n1047 GND 0.177615f
C1863 VDD.n1048 GND 0.002697f
C1864 VDD.n1049 GND 0.002171f
C1865 VDD.n1050 GND 0.002697f
C1866 VDD.n1051 GND 0.002697f
C1867 VDD.n1052 GND 0.006612f
C1868 VDD.n1053 GND 0.006442f
C1869 VDD.n1054 GND 0.002697f
C1870 VDD.n1055 GND 0.002697f
C1871 VDD.n1056 GND 0.002171f
C1872 VDD.n1057 GND 0.002697f
C1873 VDD.n1058 GND 0.113674f
C1874 VDD.n1059 GND 0.002697f
C1875 VDD.n1060 GND 0.002171f
C1876 VDD.n1061 GND 0.002697f
C1877 VDD.n1062 GND 0.002697f
C1878 VDD.n1063 GND 0.002697f
C1879 VDD.n1064 GND 0.002171f
C1880 VDD.n1065 GND 0.002171f
C1881 VDD.n1066 GND 0.002697f
C1882 VDD.n1067 GND 0.002171f
C1883 VDD.n1068 GND 0.001969f
C1884 VDD.n1069 GND 0.002171f
C1885 VDD.n1071 GND 0.002697f
C1886 VDD.n1072 GND 0.002697f
C1887 VDD.n1073 GND 0.002697f
C1888 VDD.n1074 GND 0.002171f
C1889 VDD.n1076 GND 0.002697f
C1890 VDD.n1077 GND 0.002697f
C1891 VDD.n1078 GND 0.002697f
C1892 VDD.n1079 GND 0.002697f
C1893 VDD.n1080 GND 0.002697f
C1894 VDD.n1081 GND 0.002171f
C1895 VDD.n1083 GND 0.002697f
C1896 VDD.n1084 GND 0.002697f
C1897 VDD.n1085 GND 0.002697f
C1898 VDD.n1086 GND 0.002697f
C1899 VDD.n1087 GND 0.002697f
C1900 VDD.n1088 GND 0.002171f
C1901 VDD.n1090 GND 0.002697f
C1902 VDD.n1091 GND 0.002697f
C1903 VDD.n1092 GND 0.002697f
C1904 VDD.n1093 GND 0.002697f
C1905 VDD.n1094 GND 0.002697f
C1906 VDD.n1095 GND 0.002171f
C1907 VDD.n1097 GND 0.002697f
C1908 VDD.n1098 GND 0.002697f
C1909 VDD.n1099 GND 0.002697f
C1910 VDD.n1100 GND 0.002697f
C1911 VDD.n1101 GND 0.002697f
C1912 VDD.n1102 GND 0.002171f
C1913 VDD.n1104 GND 0.002697f
C1914 VDD.n1105 GND 0.002697f
C1915 VDD.n1106 GND 0.002697f
C1916 VDD.n1107 GND 0.002697f
C1917 VDD.n1108 GND 0.002697f
C1918 VDD.n1109 GND 0.002171f
C1919 VDD.n1111 GND 0.002697f
C1920 VDD.n1112 GND 0.002697f
C1921 VDD.n1113 GND 0.002697f
C1922 VDD.n1114 GND 0.002697f
C1923 VDD.n1115 GND 0.002697f
C1924 VDD.n1116 GND 0.002171f
C1925 VDD.n1118 GND 0.002697f
C1926 VDD.n1119 GND 0.002697f
C1927 VDD.n1120 GND 0.002697f
C1928 VDD.n1121 GND 0.002697f
C1929 VDD.n1122 GND 0.002171f
C1930 VDD.n1124 GND 0.002697f
C1931 VDD.n1126 GND 0.002697f
C1932 VDD.n1127 GND 0.002171f
C1933 VDD.n1128 GND 0.002171f
C1934 VDD.n1129 GND 0.002697f
C1935 VDD.n1131 GND 0.002697f
C1936 VDD.n1132 GND 0.002697f
C1937 VDD.n1133 GND 0.002171f
C1938 VDD.n1134 GND 0.002171f
C1939 VDD.n1135 GND 0.002171f
C1940 VDD.n1136 GND 0.002697f
C1941 VDD.n1138 GND 0.002697f
C1942 VDD.n1139 GND 0.002697f
C1943 VDD.n1140 GND 0.001444f
C1944 VDD.t33 GND 0.024975f
C1945 VDD.t32 GND 0.028713f
C1946 VDD.t31 GND 0.09359f
C1947 VDD.n1141 GND 0.022187f
C1948 VDD.n1142 GND 0.015995f
C1949 VDD.n1143 GND 0.003343f
C1950 VDD.n1144 GND 0.001096f
C1951 VDD.n1145 GND 0.002171f
C1952 VDD.n1146 GND 0.002697f
C1953 VDD.n1148 GND 0.002697f
C1954 VDD.n1149 GND 0.002697f
C1955 VDD.n1150 GND 0.002171f
C1956 VDD.n1151 GND 0.002171f
C1957 VDD.n1152 GND 0.002171f
C1958 VDD.n1153 GND 0.002697f
C1959 VDD.n1155 GND 0.002697f
C1960 VDD.n1156 GND 0.002697f
C1961 VDD.n1157 GND 0.002171f
C1962 VDD.n1158 GND 0.002171f
C1963 VDD.n1159 GND 0.002171f
C1964 VDD.n1160 GND 0.002697f
C1965 VDD.n1162 GND 0.002697f
C1966 VDD.n1163 GND 0.002697f
C1967 VDD.n1164 GND 0.001444f
C1968 VDD.t58 GND 0.024975f
C1969 VDD.t57 GND 0.028713f
C1970 VDD.t56 GND 0.09359f
C1971 VDD.n1165 GND 0.022187f
C1972 VDD.n1166 GND 0.015995f
C1973 VDD.n1167 GND 0.003343f
C1974 VDD.n1168 GND 0.001096f
C1975 VDD.n1169 GND 0.002171f
C1976 VDD.n1170 GND 0.002697f
C1977 VDD.n1172 GND 0.002697f
C1978 VDD.n1173 GND 0.002697f
C1979 VDD.n1174 GND 0.002171f
C1980 VDD.n1175 GND 0.002171f
C1981 VDD.n1176 GND 0.002171f
C1982 VDD.n1177 GND 0.002697f
C1983 VDD.n1179 GND 0.002697f
C1984 VDD.n1180 GND 0.002697f
C1985 VDD.n1181 GND 0.002171f
C1986 VDD.n1182 GND 0.002171f
C1987 VDD.n1183 GND 0.002171f
C1988 VDD.n1184 GND 0.002697f
C1989 VDD.n1186 GND 0.002697f
C1990 VDD.n1187 GND 0.002697f
C1991 VDD.n1188 GND 0.001422f
C1992 VDD.t36 GND 0.024975f
C1993 VDD.t35 GND 0.028713f
C1994 VDD.t34 GND 0.09359f
C1995 VDD.n1189 GND 0.022187f
C1996 VDD.n1190 GND 0.015995f
C1997 VDD.n1191 GND 0.003343f
C1998 VDD.n1192 GND 0.001118f
C1999 VDD.n1193 GND 0.002171f
C2000 VDD.n1194 GND 0.002697f
C2001 VDD.n1196 GND 0.002697f
C2002 VDD.n1197 GND 0.002697f
C2003 VDD.n1198 GND 0.002171f
C2004 VDD.n1200 GND 0.001834f
C2005 VDD.n1201 GND 0.001834f
C2006 VDD.n1202 GND 0.001834f
C2007 VDD.n1203 GND 0.001834f
C2008 VDD.n1204 GND 0.001834f
C2009 VDD.n1206 GND 0.001834f
C2010 VDD.n1207 GND 0.001834f
C2011 VDD.n1208 GND 0.001834f
C2012 VDD.n1209 GND 0.001834f
C2013 VDD.n1210 GND 0.001834f
C2014 VDD.n1212 GND 0.001834f
C2015 VDD.n1214 GND 0.001834f
C2016 VDD.n1215 GND 0.001834f
C2017 VDD.n1216 GND 0.001834f
C2018 VDD.n1217 GND 0.001834f
C2019 VDD.n1218 GND 0.001834f
C2020 VDD.n1220 GND 0.001834f
C2021 VDD.n1221 GND 0.001834f
C2022 VDD.n1223 GND 0.001834f
C2023 VDD.n1224 GND 0.001834f
C2024 VDD.n1226 GND 0.001834f
C2025 VDD.n1227 GND 0.001834f
C2026 VDD.t76 GND 0.036555f
C2027 VDD.t77 GND 0.041821f
C2028 VDD.t75 GND 0.169586f
C2029 VDD.n1228 GND 0.027364f
C2030 VDD.n1229 GND 0.016899f
C2031 VDD.n1230 GND 0.002621f
C2032 VDD.n1232 GND 0.001834f
C2033 VDD.n1233 GND 0.001834f
C2034 VDD.n1234 GND 0.001834f
C2035 VDD.n1235 GND 0.001834f
C2036 VDD.n1236 GND 0.001834f
C2037 VDD.n1237 GND 0.001834f
C2038 VDD.n1238 GND 0.001834f
C2039 VDD.n1239 GND 0.001834f
C2040 VDD.n1240 GND 0.001834f
C2041 VDD.n1241 GND 0.001834f
C2042 VDD.n1242 GND 0.001834f
C2043 VDD.n1243 GND 0.001834f
C2044 VDD.n1244 GND 0.001834f
C2045 VDD.n1245 GND 0.001834f
C2046 VDD.n1246 GND 0.001834f
C2047 VDD.n1247 GND 0.001834f
C2048 VDD.n1248 GND 0.001834f
C2049 VDD.n1249 GND 0.001834f
C2050 VDD.n1250 GND 0.001834f
C2051 VDD.n1251 GND 0.001834f
C2052 VDD.n1252 GND 0.001834f
C2053 VDD.n1253 GND 0.001834f
C2054 VDD.n1254 GND 0.001834f
C2055 VDD.n1255 GND 0.001834f
C2056 VDD.n1256 GND 0.001834f
C2057 VDD.n1257 GND 0.001834f
C2058 VDD.n1258 GND 0.001834f
C2059 VDD.n1259 GND 0.001834f
C2060 VDD.n1260 GND 0.001834f
C2061 VDD.n1261 GND 0.001834f
C2062 VDD.n1262 GND 0.001834f
C2063 VDD.n1263 GND 0.001834f
C2064 VDD.n1264 GND 0.001834f
C2065 VDD.n1265 GND 0.001834f
C2066 VDD.n1266 GND 0.001834f
C2067 VDD.n1267 GND 0.001834f
C2068 VDD.n1268 GND 0.001834f
C2069 VDD.n1269 GND 0.001834f
C2070 VDD.n1270 GND 0.001834f
C2071 VDD.n1271 GND 0.001834f
C2072 VDD.n1272 GND 0.001834f
C2073 VDD.n1273 GND 0.001834f
C2074 VDD.n1274 GND 0.001834f
C2075 VDD.n1275 GND 0.001834f
C2076 VDD.n1276 GND 0.001834f
C2077 VDD.n1277 GND 0.001834f
C2078 VDD.n1278 GND 0.001834f
C2079 VDD.n1279 GND 0.001834f
C2080 VDD.n1280 GND 0.001834f
C2081 VDD.n1281 GND 0.004477f
C2082 VDD.n1282 GND 0.004693f
C2083 VDD.n1283 GND 0.004693f
C2084 VDD.n1284 GND 0.001308f
C2085 VDD.n1285 GND 0.001834f
C2086 VDD.n1287 GND 0.001834f
C2087 VDD.n1288 GND 0.001443f
C2088 VDD.n1289 GND 0.001834f
C2089 VDD.n1290 GND 0.001834f
C2090 VDD.n1291 GND 0.001834f
C2091 VDD.n1293 GND 0.001834f
C2092 VDD.n1294 GND 0.001834f
C2093 VDD.n1295 GND 0.001834f
C2094 VDD.n1296 GND 0.001834f
C2095 VDD.n1297 GND 0.001834f
C2096 VDD.n1298 GND 0.001834f
C2097 VDD.n1300 GND 0.001834f
C2098 VDD.n1301 GND 0.001834f
C2099 VDD.n1302 GND 0.035715f
C2100 VDD.n1303 GND 0.002697f
C2101 VDD.n1304 GND 0.002077f
C2102 VDD.n1305 GND 0.518733f
C2103 VDD.n1307 GND 0.002171f
C2104 VDD.n1308 GND 0.002697f
C2105 VDD.n1310 GND 0.002697f
C2106 VDD.n1311 GND 0.002697f
C2107 VDD.n1313 GND 0.002697f
C2108 VDD.n1314 GND 0.002171f
C2109 VDD.n1315 GND 0.001802f
C2110 VDD.n1316 GND 0.006612f
C2111 VDD.n1317 GND 0.006442f
C2112 VDD.n1318 GND 0.001802f
C2113 VDD.n1319 GND 0.006442f
C2114 VDD.n1320 GND 0.264647f
C2115 VDD.n1321 GND 0.006442f
C2116 VDD.n1322 GND 0.006612f
C2117 VDD.n1324 GND 0.002697f
C2118 VDD.n1325 GND 0.004429f
C2119 VDD.n1326 GND 0.00216f
C2120 VDD.n1327 GND 0.002171f
C2121 VDD.n1328 GND 0.002077f
C2122 VDD.n1329 GND 0.518733f
C2123 VDD.n1330 GND 0.035715f
C2124 VDD.n1331 GND 0.001834f
C2125 VDD.n1332 GND 0.001834f
C2126 VDD.n1333 GND 0.001834f
C2127 VDD.n1334 GND 0.001443f
C2128 VDD.n1335 GND 0.004693f
C2129 VDD.t70 GND 0.036555f
C2130 VDD.t71 GND 0.041821f
C2131 VDD.t68 GND 0.169586f
C2132 VDD.n1336 GND 0.027364f
C2133 VDD.n1337 GND 0.016899f
C2134 VDD.n1338 GND 0.002621f
C2135 VDD.n1339 GND 0.001834f
C2136 VDD.n1340 GND 0.001834f
C2137 VDD.n1341 GND 0.001834f
C2138 VDD.n1342 GND 0.001834f
C2139 VDD.n1343 GND 0.001834f
C2140 VDD.n1344 GND 0.001834f
C2141 VDD.n1345 GND 0.001834f
C2142 VDD.n1346 GND 0.001834f
C2143 VDD.n1347 GND 0.001834f
C2144 VDD.n1348 GND 0.001834f
C2145 VDD.n1349 GND 0.001834f
C2146 VDD.n1350 GND 0.001834f
C2147 VDD.n1351 GND 0.001834f
C2148 VDD.n1352 GND 0.001834f
C2149 VDD.n1353 GND 0.001834f
C2150 VDD.n1354 GND 0.001834f
C2151 VDD.n1355 GND 0.001834f
C2152 VDD.n1356 GND 0.001834f
C2153 VDD.n1357 GND 0.001834f
C2154 VDD.n1358 GND 0.001834f
C2155 VDD.n1359 GND 0.001834f
C2156 VDD.n1360 GND 0.001834f
C2157 VDD.n1361 GND 0.001834f
C2158 VDD.n1362 GND 0.001834f
C2159 VDD.n1363 GND 0.001834f
C2160 VDD.n1364 GND 0.001834f
C2161 VDD.n1365 GND 0.001834f
C2162 VDD.n1366 GND 0.001834f
C2163 VDD.n1367 GND 0.001834f
C2164 VDD.n1368 GND 0.001834f
C2165 VDD.n1369 GND 0.001834f
C2166 VDD.n1370 GND 0.001834f
C2167 VDD.n1371 GND 0.001834f
C2168 VDD.n1372 GND 0.001834f
C2169 VDD.n1373 GND 0.001834f
C2170 VDD.n1374 GND 0.001834f
C2171 VDD.n1375 GND 0.001834f
C2172 VDD.n1376 GND 0.001834f
C2173 VDD.n1377 GND 0.001834f
C2174 VDD.n1378 GND 0.001834f
C2175 VDD.n1379 GND 0.001834f
C2176 VDD.n1380 GND 0.001834f
C2177 VDD.n1381 GND 0.001834f
C2178 VDD.n1382 GND 0.004477f
C2179 VDD.n1383 GND 0.004693f
C2180 VDD.n1384 GND 0.001308f
C2181 VDD.n1385 GND 0.001834f
C2182 VDD.n1387 GND 0.001834f
C2183 VDD.n1389 GND 0.001834f
C2184 VDD.n1390 GND 0.001834f
C2185 VDD.n1391 GND 0.001834f
C2186 VDD.n1392 GND 0.001834f
C2187 VDD.n1393 GND 0.001834f
C2188 VDD.n1395 GND 0.001834f
C2189 VDD.n1397 GND 0.001834f
C2190 VDD.n1398 GND 0.001834f
C2191 VDD.n1399 GND 0.001834f
C2192 VDD.n1400 GND 0.001834f
C2193 VDD.n1401 GND 0.001834f
C2194 VDD.n1403 GND 0.001834f
C2195 VDD.n1405 GND 0.001834f
C2196 VDD.n1406 GND 0.001834f
C2197 VDD.n1407 GND 0.001834f
C2198 VDD.n1408 GND 0.001834f
C2199 VDD.n1409 GND 0.001834f
C2200 VDD.n1411 GND 0.001834f
C2201 VDD.n1413 GND 0.001834f
C2202 VDD.n1414 GND 0.001834f
C2203 VDD.n1415 GND 0.001834f
C2204 VDD.n1416 GND 0.001834f
C2205 VDD.n1417 GND 0.001834f
C2206 VDD.n1419 GND 0.001834f
C2207 VDD.n1421 GND 0.001834f
C2208 VDD.n1422 GND 0.001834f
C2209 VDD.n1423 GND 0.004693f
C2210 VDD.n1424 GND 0.004477f
C2211 VDD.n1425 GND 0.004477f
C2212 VDD.n1426 GND 0.182944f
C2213 VDD.n1427 GND 0.004477f
C2214 VDD.n1428 GND 0.004477f
C2215 VDD.n1429 GND 0.001834f
C2216 VDD.n1430 GND 0.001834f
C2217 VDD.n1431 GND 0.001834f
C2218 VDD.n1432 GND 0.120778f
C2219 VDD.n1433 GND 0.001834f
C2220 VDD.n1434 GND 0.001834f
C2221 VDD.n1435 GND 0.001834f
C2222 VDD.n1436 GND 0.001834f
C2223 VDD.n1437 GND 0.001834f
C2224 VDD.n1438 GND 0.120778f
C2225 VDD.n1439 GND 0.001834f
C2226 VDD.n1440 GND 0.001834f
C2227 VDD.n1441 GND 0.001834f
C2228 VDD.n1442 GND 0.001834f
C2229 VDD.n1443 GND 0.001834f
C2230 VDD.n1444 GND 0.077263f
C2231 VDD.n1445 GND 0.001834f
C2232 VDD.n1446 GND 0.001834f
C2233 VDD.n1447 GND 0.001834f
C2234 VDD.n1448 GND 0.001834f
C2235 VDD.n1449 GND 0.001834f
C2236 VDD.n1450 GND 0.120778f
C2237 VDD.n1451 GND 0.001834f
C2238 VDD.n1452 GND 0.001834f
C2239 VDD.n1453 GND 0.001834f
C2240 VDD.n1454 GND 0.001834f
C2241 VDD.n1455 GND 0.001834f
C2242 VDD.n1456 GND 0.120778f
C2243 VDD.n1457 GND 0.001834f
C2244 VDD.n1458 GND 0.001834f
C2245 VDD.n1459 GND 0.001834f
C2246 VDD.n1460 GND 0.001834f
C2247 VDD.n1461 GND 0.001834f
C2248 VDD.n1462 GND 0.120778f
C2249 VDD.n1463 GND 0.001834f
C2250 VDD.n1464 GND 0.001834f
C2251 VDD.n1465 GND 0.001834f
C2252 VDD.n1466 GND 0.001834f
C2253 VDD.n1467 GND 0.001834f
C2254 VDD.n1468 GND 0.100353f
C2255 VDD.n1469 GND 0.001834f
C2256 VDD.n1470 GND 0.001834f
C2257 VDD.n1471 GND 0.001834f
C2258 VDD.n1472 GND 0.001834f
C2259 VDD.n1473 GND 0.001834f
C2260 VDD.n1474 GND 0.120778f
C2261 VDD.n1475 GND 0.001834f
C2262 VDD.n1476 GND 0.001834f
C2263 VDD.n1477 GND 0.001834f
C2264 VDD.n1478 GND 0.001834f
C2265 VDD.n1479 GND 0.001834f
C2266 VDD.n1480 GND 0.090584f
C2267 VDD.n1481 GND 0.001834f
C2268 VDD.n1482 GND 0.001834f
C2269 VDD.n1483 GND 0.001834f
C2270 VDD.n1484 GND 0.001834f
C2271 VDD.n1485 GND 0.001834f
C2272 VDD.n1486 GND 0.120778f
C2273 VDD.n1487 GND 0.001834f
C2274 VDD.n1488 GND 0.001834f
C2275 VDD.n1489 GND 0.001834f
C2276 VDD.n1490 GND 0.001834f
C2277 VDD.n1491 GND 0.001834f
C2278 VDD.n1492 GND 0.120778f
C2279 VDD.n1493 GND 0.001834f
C2280 VDD.n1494 GND 0.001834f
C2281 VDD.n1495 GND 0.001834f
C2282 VDD.n1496 GND 0.001834f
C2283 VDD.n1497 GND 0.001834f
C2284 VDD.n1498 GND 0.084367f
C2285 VDD.n1499 GND 0.001834f
C2286 VDD.n1500 GND 0.001834f
C2287 VDD.n1501 GND 0.001834f
C2288 VDD.n1502 GND 0.001834f
C2289 VDD.n1503 GND 0.001834f
C2290 VDD.n1504 GND 0.120778f
C2291 VDD.n1505 GND 0.001834f
C2292 VDD.n1506 GND 0.001834f
C2293 VDD.n1507 GND 0.001834f
C2294 VDD.n1508 GND 0.001834f
C2295 VDD.n1509 GND 0.001834f
C2296 VDD.n1510 GND 0.001834f
C2297 VDD.n1511 GND 0.001834f
C2298 VDD.n1512 GND 0.120778f
C2299 VDD.n1513 GND 0.001834f
C2300 VDD.n1514 GND 0.001834f
C2301 VDD.n1515 GND 0.001834f
C2302 VDD.n1516 GND 0.001834f
C2303 VDD.n1517 GND 0.001834f
C2304 VDD.n1518 GND 0.081703f
C2305 VDD.n1519 GND 0.001834f
C2306 VDD.n1520 GND 0.001834f
C2307 VDD.n1521 GND 0.001834f
C2308 VDD.n1522 GND 0.001834f
C2309 VDD.n1523 GND 0.001834f
C2310 VDD.n1524 GND 0.001834f
C2311 VDD.n1525 GND 0.001834f
C2312 VDD.n1526 GND 0.004477f
C2313 VDD.n1527 GND 0.004674f
C2314 VDD.n1528 GND 0.004497f
C2315 VDD.n1529 GND 0.001834f
C2316 VDD.n1530 GND 0.001308f
C2317 VDD.n1531 GND 0.002621f
C2318 VDD.n1532 GND 0.001443f
C2319 VDD.n1533 GND 0.001834f
C2320 VDD.n1534 GND 0.001834f
C2321 VDD.n1535 GND 0.001834f
C2322 VDD.n1536 GND 0.001834f
C2323 VDD.n1537 GND 0.001834f
C2324 VDD.n1538 GND 0.001834f
C2325 VDD.n1539 GND 0.001834f
C2326 VDD.n1540 GND 0.001834f
C2327 VDD.n1541 GND 0.001834f
C2328 VDD.n1542 GND 0.001834f
C2329 VDD.n1543 GND 0.001834f
C2330 VDD.n1544 GND 0.001834f
C2331 VDD.n1545 GND 0.001834f
C2332 VDD.n1546 GND 0.001834f
C2333 VDD.n1547 GND 0.001834f
C2334 VDD.n1548 GND 0.001834f
C2335 VDD.n1549 GND 0.001834f
C2336 VDD.n1550 GND 0.001834f
C2337 VDD.n1551 GND 0.001834f
C2338 VDD.n1552 GND 0.001834f
C2339 VDD.n1553 GND 0.001834f
C2340 VDD.n1554 GND 0.001834f
C2341 VDD.n1555 GND 0.001834f
C2342 VDD.n1556 GND 0.001834f
C2343 VDD.n1557 GND 0.001834f
C2344 VDD.n1558 GND 0.001834f
C2345 VDD.n1559 GND 0.001834f
C2346 VDD.n1560 GND 0.001834f
C2347 VDD.n1561 GND 0.001834f
C2348 VDD.n1562 GND 0.001834f
C2349 VDD.n1563 GND 0.001834f
C2350 VDD.n1564 GND 0.001834f
C2351 VDD.n1565 GND 0.001834f
C2352 VDD.n1566 GND 0.001834f
C2353 VDD.n1567 GND 0.001834f
C2354 VDD.n1568 GND 0.004693f
C2355 VDD.n1569 GND 0.004693f
C2356 VDD.n1570 GND 0.004477f
C2357 VDD.n1571 GND 0.004477f
C2358 VDD.n1572 GND 0.001834f
C2359 VDD.n1573 GND 0.001834f
C2360 VDD.n1574 GND 0.001834f
C2361 VDD.n1575 GND 0.001834f
C2362 VDD.n1576 GND 0.093248f
C2363 VDD.n1577 GND 0.001834f
C2364 VDD.n1578 GND 0.001834f
C2365 VDD.n1579 GND 0.001834f
C2366 VDD.n1580 GND 0.001834f
C2367 VDD.n1581 GND 0.001834f
C2368 VDD.n1582 GND 0.120778f
C2369 VDD.n1583 GND 0.001834f
C2370 VDD.n1584 GND 0.004477f
C2371 VDD.n1585 GND 0.004693f
C2372 VDD.n1586 GND 0.004497f
C2373 VDD.n1587 GND 0.001308f
C2374 VDD.n1588 GND 0.001834f
C2375 VDD.n1589 GND 0.001834f
C2376 VDD.n1590 GND 0.001443f
C2377 VDD.n1591 GND 0.001834f
C2378 VDD.n1592 GND 0.001834f
C2379 VDD.n1593 GND 0.001834f
C2380 VDD.n1594 GND 0.001834f
C2381 VDD.n1595 GND 0.001834f
C2382 VDD.n1596 GND 0.001834f
C2383 VDD.n1597 GND 0.001834f
C2384 VDD.n1598 GND 0.001834f
C2385 VDD.n1599 GND 0.001834f
C2386 VDD.n1600 GND 0.001834f
C2387 VDD.n1601 GND 0.001834f
C2388 VDD.n1602 GND 0.001834f
C2389 VDD.n1603 GND 0.001834f
C2390 VDD.n1604 GND 0.001834f
C2391 VDD.n1605 GND 0.001834f
C2392 VDD.n1606 GND 0.001834f
C2393 VDD.n1607 GND 0.001834f
C2394 VDD.n1608 GND 0.001834f
C2395 VDD.n1609 GND 0.001834f
C2396 VDD.n1610 GND 0.001834f
C2397 VDD.n1611 GND 0.001834f
C2398 VDD.n1612 GND 0.001834f
C2399 VDD.n1613 GND 0.001834f
C2400 VDD.n1614 GND 0.001834f
C2401 VDD.n1615 GND 0.001834f
C2402 VDD.n1616 GND 0.001834f
C2403 VDD.n1617 GND 0.001834f
C2404 VDD.n1618 GND 0.001834f
C2405 VDD.n1619 GND 0.001834f
C2406 VDD.n1620 GND 0.001834f
C2407 VDD.n1621 GND 0.001834f
C2408 VDD.n1622 GND 0.001834f
C2409 VDD.n1623 GND 0.001834f
C2410 VDD.n1624 GND 0.004693f
C2411 VDD.n1625 GND 0.004693f
C2412 VDD.n1626 GND 0.767298f
C2413 VDD.n1627 GND 0.767298f
C2414 VDD.n1628 GND 0.004477f
C2415 VDD.n1629 GND 0.004693f
C2416 VDD.n1630 GND 0.001834f
C2417 VDD.t3 GND 0.036555f
C2418 VDD.t4 GND 0.041821f
C2419 VDD.t1 GND 0.169586f
C2420 VDD.n1631 GND 0.027364f
C2421 VDD.n1632 GND 0.016899f
C2422 VDD.n1633 GND 0.002621f
C2423 VDD.n1634 GND 0.001834f
C2424 VDD.n1635 GND 0.001834f
C2425 VDD.n1636 GND 0.001834f
C2426 VDD.n1637 GND 0.001834f
C2427 VDD.n1638 GND 0.001834f
C2428 VDD.n1639 GND 0.001834f
C2429 VDD.n1640 GND 0.001834f
C2430 VDD.n1641 GND 0.001834f
C2431 VDD.n1643 GND 0.001834f
C2432 VDD.n1644 GND 0.001834f
C2433 VDD.n1645 GND 0.001834f
C2434 VDD.n1646 GND 0.001834f
C2435 VDD.n1648 GND 0.001834f
C2436 VDD.n1650 GND 0.001834f
C2437 VDD.n1651 GND 0.001834f
C2438 VDD.n1652 GND 0.001834f
C2439 VDD.n1653 GND 0.001834f
C2440 VDD.n1654 GND 0.001834f
C2441 VDD.n1656 GND 0.001834f
C2442 VDD.n1658 GND 0.001834f
C2443 VDD.n1659 GND 0.001834f
C2444 VDD.n1660 GND 0.001834f
C2445 VDD.n1661 GND 0.001834f
C2446 VDD.n1662 GND 0.001834f
C2447 VDD.n1664 GND 0.001834f
C2448 VDD.n1666 GND 0.001834f
C2449 VDD.n1667 GND 0.001834f
C2450 VDD.n1668 GND 0.001834f
C2451 VDD.n1669 GND 0.001834f
C2452 VDD.n1670 GND 0.001834f
C2453 VDD.n1672 GND 0.001834f
C2454 VDD.n1674 GND 0.001834f
C2455 VDD.n1675 GND 0.001834f
C2456 VDD.n1676 GND 0.001834f
C2457 VDD.n1677 GND 0.001443f
C2458 VDD.n1678 GND 0.001834f
C2459 VDD.n1680 GND 0.001834f
C2460 VDD.n1681 GND 0.001308f
C2461 VDD.n1682 GND 0.004693f
C2462 VDD.n1683 GND 0.001834f
C2463 VDD.n1684 GND 0.001834f
C2464 VDD.n1685 GND 0.001834f
C2465 VDD.n1686 GND 0.001834f
C2466 VDD.n1687 GND 0.001834f
C2467 VDD.n1688 GND 0.001834f
C2468 VDD.n1689 GND 0.001834f
C2469 VDD.n1690 GND 0.001834f
C2470 VDD.n1691 GND 0.001834f
C2471 VDD.n1692 GND 0.001834f
C2472 VDD.n1693 GND 0.001834f
C2473 VDD.n1694 GND 0.001834f
C2474 VDD.n1695 GND 0.001834f
C2475 VDD.n1696 GND 0.001834f
C2476 VDD.n1697 GND 0.001834f
C2477 VDD.n1698 GND 0.001834f
C2478 VDD.n1699 GND 0.001834f
C2479 VDD.n1700 GND 0.001834f
C2480 VDD.n1701 GND 0.001834f
C2481 VDD.n1702 GND 0.001834f
C2482 VDD.n1703 GND 0.001834f
C2483 VDD.n1704 GND 0.001834f
C2484 VDD.n1705 GND 0.001834f
C2485 VDD.n1706 GND 0.001834f
C2486 VDD.n1707 GND 0.001834f
C2487 VDD.n1708 GND 0.001834f
C2488 VDD.n1709 GND 0.001834f
C2489 VDD.n1710 GND 0.001834f
C2490 VDD.n1711 GND 0.001834f
C2491 VDD.n1712 GND 0.001834f
C2492 VDD.n1713 GND 0.001834f
C2493 VDD.n1714 GND 0.001834f
C2494 VDD.n1715 GND 0.001834f
C2495 VDD.n1716 GND 0.001834f
C2496 VDD.n1717 GND 0.001834f
C2497 VDD.n1718 GND 0.001834f
C2498 VDD.n1719 GND 0.001834f
C2499 VDD.n1720 GND 0.001834f
C2500 VDD.n1721 GND 0.001834f
C2501 VDD.n1722 GND 0.001834f
C2502 VDD.n1723 GND 0.001834f
C2503 VDD.n1724 GND 0.001834f
C2504 VDD.n1725 GND 0.001834f
C2505 VDD.n1726 GND 0.001834f
C2506 VDD.n1727 GND 0.001834f
C2507 VDD.n1728 GND 0.001834f
C2508 VDD.n1729 GND 0.001834f
C2509 VDD.n1730 GND 0.004477f
C2510 VDD.n1731 GND 0.004477f
C2511 VDD.n1732 GND 0.004693f
C2512 VDD.n1733 GND 0.001834f
C2513 VDD.n1735 GND 0.001834f
C2514 VDD.n1736 GND 0.001834f
C2515 VDD.n1737 GND 0.001834f
C2516 VDD.n1738 GND 0.001834f
C2517 VDD.n1739 GND 0.001834f
C2518 VDD.n1740 GND 0.001834f
C2519 VDD.n1741 GND 0.001834f
C2520 VDD.n1742 GND 0.001834f
C2521 VDD.t14 GND 0.036555f
C2522 VDD.t15 GND 0.041821f
C2523 VDD.t13 GND 0.169586f
C2524 VDD.n1743 GND 0.027364f
C2525 VDD.n1744 GND 0.016899f
C2526 VDD.n1745 GND 0.001834f
C2527 VDD.n1746 GND 0.001834f
C2528 VDD.n1747 GND 0.001834f
C2529 VDD.n1748 GND 0.001834f
C2530 VDD.n1749 GND 0.001834f
C2531 VDD.n1750 GND 0.001834f
C2532 VDD.n1751 GND 0.001834f
C2533 VDD.n1752 GND 0.001834f
C2534 VDD.n1753 GND 0.001834f
C2535 VDD.n1754 GND 0.001834f
C2536 VDD.n1755 GND 0.001834f
C2537 VDD.n1756 GND 0.001834f
C2538 VDD.n1757 GND 0.001834f
C2539 VDD.n1758 GND 0.001834f
C2540 VDD.n1759 GND 0.001834f
C2541 VDD.n1760 GND 0.001834f
C2542 VDD.n1761 GND 0.001834f
C2543 VDD.n1762 GND 0.001834f
C2544 VDD.n1763 GND 0.001834f
C2545 VDD.n1764 GND 0.001834f
C2546 VDD.n1765 GND 0.001834f
C2547 VDD.n1766 GND 0.001834f
C2548 VDD.n1767 GND 0.001834f
C2549 VDD.n1768 GND 0.001834f
C2550 VDD.n1769 GND 0.001834f
C2551 VDD.n1770 GND 0.001834f
C2552 VDD.n1771 GND 0.001834f
C2553 VDD.n1772 GND 0.001834f
C2554 VDD.n1773 GND 0.001834f
C2555 VDD.n1774 GND 0.001834f
C2556 VDD.n1775 GND 0.001834f
C2557 VDD.n1776 GND 0.001834f
C2558 VDD.n1777 GND 0.001834f
C2559 VDD.n1778 GND 0.001834f
C2560 VDD.n1779 GND 0.001834f
C2561 VDD.n1780 GND 0.001834f
C2562 VDD.n1781 GND 0.001834f
C2563 VDD.n1782 GND 0.001834f
C2564 VDD.n1783 GND 0.001834f
C2565 VDD.n1784 GND 0.001834f
C2566 VDD.n1785 GND 0.001834f
C2567 VDD.n1786 GND 0.001834f
C2568 VDD.n1787 GND 0.001834f
C2569 VDD.n1788 GND 0.001834f
C2570 VDD.n1789 GND 0.001834f
C2571 VDD.n1790 GND 0.001834f
C2572 VDD.n1791 GND 0.004477f
C2573 VDD.n1793 GND 0.004693f
C2574 VDD.n1794 GND 0.004693f
C2575 VDD.n1795 GND 0.001308f
C2576 VDD.n1796 GND 0.002621f
C2577 VDD.n1797 GND 0.001443f
C2578 VDD.n1798 GND 0.001834f
C2579 VDD.n1800 GND 0.001834f
C2580 VDD.n1802 GND 0.001834f
C2581 VDD.n1803 GND 0.001834f
C2582 VDD.n1804 GND 0.001834f
C2583 VDD.n1805 GND 0.001834f
C2584 VDD.n1806 GND 0.001834f
C2585 VDD.n1808 GND 0.001834f
C2586 VDD.n1810 GND 0.001834f
C2587 VDD.n1811 GND 0.001834f
C2588 VDD.n1812 GND 0.001834f
C2589 VDD.n1813 GND 0.001834f
C2590 VDD.n1814 GND 0.001834f
C2591 VDD.n1816 GND 0.001834f
C2592 VDD.n1818 GND 0.001834f
C2593 VDD.n1819 GND 0.001834f
C2594 VDD.n1820 GND 0.001834f
C2595 VDD.n1821 GND 0.001834f
C2596 VDD.n1822 GND 0.001834f
C2597 VDD.n1824 GND 0.001834f
C2598 VDD.n1825 GND 0.001834f
C2599 VDD.n1826 GND 0.001834f
C2600 VDD.n1827 GND 0.001834f
C2601 VDD.n1828 GND 0.001834f
C2602 VDD.n1829 GND 0.001834f
C2603 VDD.n1831 GND 0.001834f
C2604 VDD.n1832 GND 0.001834f
C2605 VDD.n1833 GND 0.004693f
C2606 VDD.n1834 GND 0.004477f
C2607 VDD.n1835 GND 0.004477f
C2608 VDD.n1836 GND 0.182944f
C2609 VDD.n1837 GND 0.004477f
C2610 VDD.n1838 GND 0.004477f
C2611 VDD.n1839 GND 0.001834f
C2612 VDD.n1840 GND 0.001834f
C2613 VDD.n1841 GND 0.001834f
C2614 VDD.n1842 GND 0.08792f
C2615 VDD.n1843 GND 0.001834f
C2616 VDD.n1844 GND 0.001834f
C2617 VDD.n1845 GND 0.001834f
C2618 VDD.n1846 GND 0.001834f
C2619 VDD.n1847 GND 0.001834f
C2620 VDD.n1848 GND 0.120778f
C2621 VDD.n1849 GND 0.001834f
C2622 VDD.n1850 GND 0.001834f
C2623 VDD.n1851 GND 0.001834f
C2624 VDD.n1852 GND 0.001834f
C2625 VDD.n1853 GND 0.001834f
C2626 VDD.n1854 GND 0.099464f
C2627 VDD.n1855 GND 0.001834f
C2628 VDD.n1856 GND 0.001834f
C2629 VDD.n1857 GND 0.001834f
C2630 VDD.n1858 GND 0.001834f
C2631 VDD.n1859 GND 0.001834f
C2632 VDD.n1860 GND 0.120778f
C2633 VDD.n1861 GND 0.001834f
C2634 VDD.n1862 GND 0.001834f
C2635 VDD.n1863 GND 0.001834f
C2636 VDD.n1864 GND 0.001834f
C2637 VDD.n1865 GND 0.001834f
C2638 VDD.n1866 GND 0.120778f
C2639 VDD.n1867 GND 0.001834f
C2640 VDD.n1868 GND 0.001834f
C2641 VDD.n1869 GND 0.001834f
C2642 VDD.n1870 GND 0.001834f
C2643 VDD.n1871 GND 0.001834f
C2644 VDD.n1872 GND 0.0968f
C2645 VDD.n1873 GND 0.001834f
C2646 VDD.n1874 GND 0.001834f
C2647 VDD.n1875 GND 0.001834f
C2648 VDD.n1876 GND 0.001834f
C2649 VDD.n1877 GND 0.001834f
C2650 VDD.n1878 GND 0.120778f
C2651 VDD.n1879 GND 0.001834f
C2652 VDD.n1880 GND 0.001834f
C2653 VDD.n1881 GND 0.001834f
C2654 VDD.n1882 GND 0.001834f
C2655 VDD.n1883 GND 0.001834f
C2656 VDD.n1884 GND 0.120778f
C2657 VDD.n1885 GND 0.001834f
C2658 VDD.n1886 GND 0.001834f
C2659 VDD.n1887 GND 0.001834f
C2660 VDD.n1888 GND 0.001834f
C2661 VDD.n1889 GND 0.001834f
C2662 VDD.n1890 GND 0.090584f
C2663 VDD.n1891 GND 0.001834f
C2664 VDD.n1892 GND 0.001834f
C2665 VDD.n1893 GND 0.001834f
C2666 VDD.n1894 GND 0.001834f
C2667 VDD.n1895 GND 0.001834f
C2668 VDD.n1896 GND 0.080815f
C2669 VDD.n1897 GND 0.001834f
C2670 VDD.n1898 GND 0.001834f
C2671 VDD.n1899 GND 0.001834f
C2672 VDD.n1900 GND 0.001834f
C2673 VDD.n1901 GND 0.001834f
C2674 VDD.n1902 GND 0.120778f
C2675 VDD.n1903 GND 0.001834f
C2676 VDD.n1904 GND 0.001834f
C2677 VDD.n1905 GND 0.001834f
C2678 VDD.n1906 GND 0.001834f
C2679 VDD.n1907 GND 0.001834f
C2680 VDD.n1908 GND 0.120778f
C2681 VDD.n1909 GND 0.001834f
C2682 VDD.n1910 GND 0.001834f
C2683 VDD.n1911 GND 0.001834f
C2684 VDD.n1912 GND 0.001834f
C2685 VDD.n1913 GND 0.001834f
C2686 VDD.n1914 GND 0.120778f
C2687 VDD.n1915 GND 0.001834f
C2688 VDD.n1916 GND 0.001834f
C2689 VDD.n1917 GND 0.001834f
C2690 VDD.n1918 GND 0.001834f
C2691 VDD.n1919 GND 0.001834f
C2692 VDD.n1920 GND 0.120778f
C2693 VDD.n1921 GND 0.001834f
C2694 VDD.n1922 GND 0.001834f
C2695 VDD.n1923 GND 0.001834f
C2696 VDD.n1924 GND 0.004693f
C2697 VDD.n1925 GND 0.001834f
C2698 VDD.n1926 GND 0.001834f
C2699 VDD.n1927 GND 0.001834f
C2700 VDD.n1929 GND 0.001834f
C2701 VDD.n1931 GND 0.001834f
C2702 VDD.n1932 GND 0.001834f
C2703 VDD.n1933 GND 0.001834f
C2704 VDD.n1934 GND 0.001834f
C2705 VDD.n1935 GND 0.001834f
C2706 VDD.n1936 GND 0.001834f
C2707 VDD.n1938 GND 0.001834f
C2708 VDD.n1939 GND 0.001834f
C2709 VDD.n1940 GND 0.001834f
C2710 VDD.n1941 GND 0.001834f
C2711 VDD.n1942 GND 0.001834f
C2712 VDD.n1943 GND 0.001834f
C2713 VDD.n1945 GND 0.001834f
C2714 VDD.n1946 GND 0.004693f
C2715 VDD.n1947 GND 0.004477f
C2716 VDD.n1948 GND 0.004477f
C2717 VDD.n1949 GND 0.001834f
C2718 VDD.n1950 GND 0.001834f
C2719 VDD.n1951 GND 0.001834f
C2720 VDD.n1952 GND 0.001834f
C2721 VDD.n1953 GND 0.001834f
C2722 VDD.n1954 GND 0.001834f
C2723 VDD.n1955 GND 0.001834f
C2724 VDD.n1956 GND 0.081703f
C2725 VDD.n1957 GND 0.001834f
C2726 VDD.n1958 GND 0.001834f
C2727 VDD.n1959 GND 0.001834f
C2728 VDD.n1960 GND 0.001834f
C2729 VDD.n1961 GND 0.001834f
C2730 VDD.n1962 GND 0.120778f
C2731 VDD.n1963 GND 0.001834f
C2732 VDD.n1964 GND 0.001834f
C2733 VDD.n1965 GND 0.001834f
C2734 VDD.n1966 GND 0.001834f
C2735 VDD.n1967 GND 0.004674f
C2736 VDD.n1969 GND 0.004477f
C2737 VDD.n1970 GND 0.004693f
C2738 VDD.n1971 GND 0.004497f
C2739 VDD.n1972 GND 0.001308f
C2740 VDD.n1973 GND 0.002621f
C2741 VDD.n1974 GND 0.001443f
C2742 VDD.n1975 GND 0.001834f
C2743 VDD.n1977 GND 0.001834f
C2744 VDD.n1978 GND 0.001834f
C2745 VDD.n1979 GND 0.001834f
C2746 VDD.n1980 GND 0.001834f
C2747 VDD.n1981 GND 0.001834f
C2748 VDD.n1982 GND 0.001834f
C2749 VDD.n1984 GND 0.001834f
C2750 VDD.n1985 GND 0.001834f
C2751 VDD.n1986 GND 0.001834f
C2752 VDD.n1987 GND 0.001834f
C2753 VDD.n1988 GND 0.519704f
C2754 VDD.n1989 GND 0.034744f
C2755 VDD.n1990 GND 0.001834f
C2756 VDD.n1992 GND 0.001834f
C2757 VDD.n1993 GND 0.001834f
C2758 VDD.n1994 GND 0.001834f
C2759 VDD.n1995 GND 0.001834f
C2760 VDD.n1996 GND 0.001834f
C2761 VDD.n1997 GND 0.001834f
C2762 VDD.n1999 GND 0.001834f
C2763 VDD.n2000 GND 0.001834f
C2764 VDD.n2001 GND 0.001834f
C2765 VDD.n2002 GND 0.001834f
C2766 VDD.n2003 GND 0.001834f
C2767 VDD.n2004 GND 0.001834f
C2768 VDD.n2006 GND 0.001834f
C2769 VDD.n2007 GND 0.004693f
C2770 VDD.n2008 GND 0.004693f
C2771 VDD.n2009 GND 0.004477f
C2772 VDD.n2010 GND 0.001834f
C2773 VDD.n2011 GND 0.001834f
C2774 VDD.n2012 GND 0.120778f
C2775 VDD.n2013 GND 0.001834f
C2776 VDD.n2014 GND 0.001834f
C2777 VDD.n2015 GND 0.004674f
C2778 VDD.n2016 GND 0.004497f
C2779 VDD.n2017 GND 0.004693f
C2780 VDD.n2019 GND 0.001834f
C2781 VDD.n2020 GND 0.001834f
C2782 VDD.n2021 GND 0.001443f
C2783 VDD.n2022 GND 0.001834f
C2784 VDD.n2023 GND 0.001834f
C2785 VDD.n2024 GND 0.001834f
C2786 VDD.n2026 GND 0.001834f
C2787 VDD.n2027 GND 0.001834f
C2788 VDD.n2028 GND 0.001834f
C2789 VDD.n2029 GND 0.001834f
C2790 VDD.n2030 GND 0.001834f
C2791 VDD.n2031 GND 0.001834f
C2792 VDD.n2033 GND 0.001834f
C2793 VDD.n2034 GND 0.001834f
C2794 VDD.n2035 GND 0.034744f
C2795 VDD.n2036 GND 0.002697f
C2796 VDD.n2037 GND 0.002697f
C2797 VDD.n2038 GND 0.002171f
C2798 VDD.n2039 GND 0.002697f
C2799 VDD.n2040 GND 0.002697f
C2800 VDD.n2041 GND 0.006612f
C2801 VDD.n2042 GND 0.001096f
C2802 VDD.n2043 GND 0.006612f
C2803 VDD.n2044 GND 0.002697f
C2804 VDD.t29 GND 0.024975f
C2805 VDD.t30 GND 0.028713f
C2806 VDD.t28 GND 0.09359f
C2807 VDD.n2045 GND 0.022187f
C2808 VDD.n2046 GND 0.015995f
C2809 VDD.n2047 GND 0.004429f
C2810 VDD.n2048 GND 0.002697f
C2811 VDD.n2049 GND 0.002697f
C2812 VDD.n2050 GND 0.00216f
C2813 VDD.n2051 GND 0.002697f
C2814 VDD.n2052 GND 0.002171f
C2815 VDD.n2053 GND 0.002171f
C2816 VDD.n2055 GND 0.519704f
C2817 VDD.n2057 GND 0.002171f
C2818 VDD.n2058 GND 0.002697f
C2819 VDD.n2059 GND 0.002697f
C2820 VDD.n2060 GND 0.002171f
C2821 VDD.n2061 GND 0.002171f
C2822 VDD.n2062 GND 0.002697f
C2823 VDD.n2063 GND 0.002697f
C2824 VDD.n2064 GND 0.002171f
C2825 VDD.n2065 GND 0.002171f
C2826 VDD.n2066 GND 0.002697f
C2827 VDD.n2067 GND 0.002697f
C2828 VDD.n2068 GND 0.001444f
C2829 VDD.t51 GND 0.024975f
C2830 VDD.t52 GND 0.028713f
C2831 VDD.t50 GND 0.09359f
C2832 VDD.n2069 GND 0.022187f
C2833 VDD.n2070 GND 0.015995f
C2834 VDD.n2071 GND 0.003343f
C2835 VDD.n2072 GND 0.001096f
C2836 VDD.n2073 GND 0.002697f
C2837 VDD.n2074 GND 0.002697f
C2838 VDD.n2075 GND 0.002171f
C2839 VDD.n2076 GND 0.002171f
C2840 VDD.n2077 GND 0.002697f
C2841 VDD.n2078 GND 0.002697f
C2842 VDD.n2079 GND 0.002171f
C2843 VDD.n2080 GND 0.002171f
C2844 VDD.n2081 GND 0.002697f
C2845 VDD.n2082 GND 0.002697f
C2846 VDD.n2083 GND 0.002171f
C2847 VDD.n2084 GND 0.002171f
C2848 VDD.n2085 GND 0.002697f
C2849 VDD.n2086 GND 0.002697f
C2850 VDD.n2087 GND 0.002171f
C2851 VDD.n2088 GND 0.002171f
C2852 VDD.n2089 GND 0.002697f
C2853 VDD.n2090 GND 0.002697f
C2854 VDD.n2091 GND 0.002171f
C2855 VDD.n2092 GND 0.002171f
C2856 VDD.n2093 GND 0.002697f
C2857 VDD.n2094 GND 0.002697f
C2858 VDD.n2095 GND 0.001444f
C2859 VDD.t18 GND 0.024975f
C2860 VDD.t19 GND 0.028713f
C2861 VDD.t16 GND 0.09359f
C2862 VDD.n2096 GND 0.022187f
C2863 VDD.n2097 GND 0.015995f
C2864 VDD.n2098 GND 0.003343f
C2865 VDD.n2099 GND 0.001096f
C2866 VDD.n2100 GND 0.002697f
C2867 VDD.n2101 GND 0.002697f
C2868 VDD.n2102 GND 0.002171f
C2869 VDD.n2103 GND 0.002171f
C2870 VDD.n2104 GND 0.002697f
C2871 VDD.n2105 GND 0.002697f
C2872 VDD.n2106 GND 0.002171f
C2873 VDD.n2107 GND 0.002171f
C2874 VDD.n2108 GND 0.002697f
C2875 VDD.n2109 GND 0.002697f
C2876 VDD.n2110 GND 0.002171f
C2877 VDD.n2111 GND 0.002171f
C2878 VDD.n2112 GND 0.002697f
C2879 VDD.n2113 GND 0.002697f
C2880 VDD.n2114 GND 0.002171f
C2881 VDD.n2115 GND 0.002171f
C2882 VDD.n2116 GND 0.002697f
C2883 VDD.n2117 GND 0.002697f
C2884 VDD.n2118 GND 0.002171f
C2885 VDD.n2119 GND 0.002171f
C2886 VDD.n2120 GND 0.002697f
C2887 VDD.n2121 GND 0.002697f
C2888 VDD.n2122 GND 0.001422f
C2889 VDD.t63 GND 0.024975f
C2890 VDD.t64 GND 0.028713f
C2891 VDD.t62 GND 0.09359f
C2892 VDD.n2123 GND 0.022187f
C2893 VDD.n2124 GND 0.015995f
C2894 VDD.n2125 GND 0.003343f
C2895 VDD.n2126 GND 0.001118f
C2896 VDD.n2127 GND 0.002697f
C2897 VDD.n2128 GND 0.002697f
C2898 VDD.n2129 GND 0.002171f
C2899 VDD.n2130 GND 0.002171f
C2900 VDD.n2131 GND 0.002697f
C2901 VDD.n2132 GND 0.002697f
C2902 VDD.n2133 GND 0.002171f
C2903 VDD.n2134 GND 0.002171f
C2904 VDD.n2135 GND 0.002697f
C2905 VDD.n2136 GND 0.002697f
C2906 VDD.n2137 GND 0.002171f
C2907 VDD.n2138 GND 0.002171f
C2908 VDD.n2139 GND 0.002171f
C2909 VDD.n2140 GND 0.002697f
C2910 VDD.n2141 GND 1.19357f
C2911 VDD.n2143 GND 0.006612f
C2912 VDD.n2144 GND 0.001802f
C2913 VDD.n2145 GND 0.006612f
C2914 VDD.n2146 GND 0.006442f
C2915 VDD.n2147 GND 0.002697f
C2916 VDD.n2148 GND 0.002171f
C2917 VDD.n2149 GND 0.002697f
C2918 VDD.n2150 GND 0.177615f
C2919 VDD.n2151 GND 0.002697f
C2920 VDD.n2152 GND 0.002171f
C2921 VDD.n2153 GND 0.002697f
C2922 VDD.n2154 GND 0.002697f
C2923 VDD.n2155 GND 0.002697f
C2924 VDD.n2156 GND 0.002171f
C2925 VDD.n2157 GND 0.002697f
C2926 VDD.n2158 GND 0.152749f
C2927 VDD.n2159 GND 0.002697f
C2928 VDD.n2160 GND 0.002171f
C2929 VDD.n2161 GND 0.002697f
C2930 VDD.n2162 GND 0.002697f
C2931 VDD.n2163 GND 0.002697f
C2932 VDD.n2164 GND 0.002171f
C2933 VDD.n2165 GND 0.002697f
C2934 VDD.n2166 GND 0.177615f
C2935 VDD.n2167 GND 0.002697f
C2936 VDD.n2168 GND 0.002171f
C2937 VDD.n2169 GND 0.002697f
C2938 VDD.n2170 GND 0.002697f
C2939 VDD.n2171 GND 0.002697f
C2940 VDD.n2172 GND 0.002171f
C2941 VDD.n2173 GND 0.002697f
C2942 VDD.n2174 GND 0.177615f
C2943 VDD.n2175 GND 0.002697f
C2944 VDD.n2176 GND 0.002171f
C2945 VDD.n2177 GND 0.002697f
C2946 VDD.n2178 GND 0.002697f
C2947 VDD.n2179 GND 0.002697f
C2948 VDD.n2180 GND 0.002171f
C2949 VDD.n2181 GND 0.002697f
C2950 VDD.n2182 GND 0.101241f
C2951 VDD.n2183 GND 0.002697f
C2952 VDD.n2184 GND 0.002171f
C2953 VDD.n2185 GND 0.002697f
C2954 VDD.n2186 GND 0.002697f
C2955 VDD.n2187 GND 0.002697f
C2956 VDD.n2188 GND 0.002171f
C2957 VDD.n2189 GND 0.002697f
C2958 VDD.n2190 GND 0.177615f
C2959 VDD.n2191 GND 0.002697f
C2960 VDD.n2192 GND 0.002171f
C2961 VDD.n2193 GND 0.002697f
C2962 VDD.n2194 GND 0.002697f
C2963 VDD.n2195 GND 0.002697f
C2964 VDD.n2196 GND 0.002171f
C2965 VDD.n2197 GND 0.002697f
C2966 VDD.n2198 GND 0.16163f
C2967 VDD.n2199 GND 0.002697f
C2968 VDD.n2200 GND 0.002171f
C2969 VDD.n2201 GND 0.002697f
C2970 VDD.n2202 GND 0.002697f
C2971 VDD.n2203 GND 0.002697f
C2972 VDD.n2204 GND 0.002171f
C2973 VDD.n2205 GND 0.002697f
C2974 VDD.n2206 GND 0.177615f
C2975 VDD.n2207 GND 0.002697f
C2976 VDD.n2208 GND 0.002171f
C2977 VDD.n2209 GND 0.002697f
C2978 VDD.n2210 GND 0.002697f
C2979 VDD.n2211 GND 0.002697f
C2980 VDD.n2212 GND 0.002171f
C2981 VDD.n2213 GND 0.002697f
C2982 VDD.n2214 GND 0.177615f
C2983 VDD.n2215 GND 0.002697f
C2984 VDD.n2216 GND 0.002171f
C2985 VDD.n2217 GND 0.002697f
C2986 VDD.n2218 GND 0.002697f
C2987 VDD.n2219 GND 0.002697f
C2988 VDD.n2220 GND 0.002171f
C2989 VDD.n2221 GND 0.002171f
C2990 VDD.n2222 GND 0.002171f
C2991 VDD.n2223 GND 0.002697f
C2992 VDD.n2224 GND 0.002697f
C2993 VDD.n2225 GND 0.002697f
C2994 VDD.n2226 GND 0.002171f
C2995 VDD.n2227 GND 0.002171f
C2996 VDD.n2228 GND 0.002171f
C2997 VDD.n2229 GND 0.002697f
C2998 VDD.n2230 GND 0.002697f
C2999 VDD.n2231 GND 0.002697f
C3000 VDD.n2232 GND 0.002171f
C3001 VDD.n2233 GND 0.002171f
C3002 VDD.n2234 GND 0.002171f
C3003 VDD.n2235 GND 0.002697f
C3004 VDD.n2236 GND 0.002697f
C3005 VDD.n2237 GND 0.002697f
C3006 VDD.n2238 GND 0.002171f
C3007 VDD.n2239 GND 0.002171f
C3008 VDD.n2240 GND 0.002171f
C3009 VDD.n2241 GND 0.002697f
C3010 VDD.n2242 GND 0.002697f
C3011 VDD.n2243 GND 0.002697f
C3012 VDD.n2244 GND 0.002171f
C3013 VDD.n2245 GND 0.002171f
C3014 VDD.n2246 GND 0.001802f
C3015 VDD.n2247 GND 0.006442f
C3016 VDD.n2248 GND 0.006612f
C3017 VDD.n2249 GND 0.002697f
C3018 VDD.n2250 GND 0.004429f
C3019 VDD.n2251 GND 0.00216f
C3020 VDD.n2252 GND 0.002697f
C3021 VDD.n2254 GND 0.002697f
C3022 VDD.n2255 GND 0.002697f
C3023 VDD.n2256 GND 0.002171f
C3024 VDD.n2257 GND 0.002171f
C3025 VDD.n2258 GND 0.002171f
C3026 VDD.n2259 GND 0.002697f
C3027 VDD.n2261 GND 0.002697f
C3028 VDD.n2262 GND 0.002697f
C3029 VDD.n2263 GND 0.002171f
C3030 VDD.n2264 GND 0.002171f
C3031 VDD.n2265 GND 0.002171f
C3032 VDD.n2266 GND 0.002697f
C3033 VDD.n2268 GND 0.002697f
C3034 VDD.n2269 GND 0.002697f
C3035 VDD.n2270 GND 0.001444f
C3036 VDD.t27 GND 0.024975f
C3037 VDD.t26 GND 0.028713f
C3038 VDD.t24 GND 0.09359f
C3039 VDD.n2271 GND 0.022187f
C3040 VDD.n2272 GND 0.015995f
C3041 VDD.n2273 GND 0.003343f
C3042 VDD.n2274 GND 0.001096f
C3043 VDD.n2275 GND 0.002171f
C3044 VDD.n2276 GND 0.002697f
C3045 VDD.n2278 GND 0.002697f
C3046 VDD.n2279 GND 0.002697f
C3047 VDD.n2280 GND 0.002171f
C3048 VDD.n2281 GND 0.002171f
C3049 VDD.n2282 GND 0.002171f
C3050 VDD.n2283 GND 0.002697f
C3051 VDD.n2285 GND 0.002697f
C3052 VDD.n2286 GND 0.002697f
C3053 VDD.n2287 GND 0.002171f
C3054 VDD.n2288 GND 0.002171f
C3055 VDD.n2289 GND 0.002171f
C3056 VDD.n2290 GND 0.002697f
C3057 VDD.n2292 GND 0.002697f
C3058 VDD.n2293 GND 0.002697f
C3059 VDD.n2294 GND 0.001444f
C3060 VDD.t39 GND 0.024975f
C3061 VDD.t38 GND 0.028713f
C3062 VDD.t37 GND 0.09359f
C3063 VDD.n2295 GND 0.022187f
C3064 VDD.n2296 GND 0.015995f
C3065 VDD.n2297 GND 0.003343f
C3066 VDD.n2298 GND 0.001096f
C3067 VDD.n2299 GND 0.002171f
C3068 VDD.n2300 GND 0.002697f
C3069 VDD.n2302 GND 0.002697f
C3070 VDD.n2303 GND 0.002697f
C3071 VDD.n2304 GND 0.002171f
C3072 VDD.n2305 GND 0.002171f
C3073 VDD.n2306 GND 0.002171f
C3074 VDD.n2307 GND 0.002697f
C3075 VDD.n2309 GND 0.002697f
C3076 VDD.n2310 GND 0.002697f
C3077 VDD.n2311 GND 0.002171f
C3078 VDD.n2312 GND 0.002171f
C3079 VDD.n2313 GND 0.002171f
C3080 VDD.n2314 GND 0.002697f
C3081 VDD.n2316 GND 0.002697f
C3082 VDD.n2317 GND 0.002697f
C3083 VDD.n2318 GND 0.001422f
C3084 VDD.t80 GND 0.024975f
C3085 VDD.t79 GND 0.028713f
C3086 VDD.t78 GND 0.09359f
C3087 VDD.n2319 GND 0.022187f
C3088 VDD.n2320 GND 0.015995f
C3089 VDD.n2321 GND 0.003343f
C3090 VDD.n2322 GND 0.001118f
C3091 VDD.n2323 GND 0.002171f
C3092 VDD.n2324 GND 0.002697f
C3093 VDD.n2326 GND 0.002697f
C3094 VDD.n2327 GND 0.002697f
C3095 VDD.n2328 GND 0.002171f
C3096 VDD.n2329 GND 0.002171f
C3097 VDD.n2330 GND 0.002171f
C3098 VDD.n2331 GND 0.002697f
C3099 VDD.n2333 GND 0.002697f
C3100 VDD.n2334 GND 0.002697f
C3101 VDD.n2335 GND 0.002171f
C3102 VDD.n2336 GND 0.002171f
C3103 VDD.n2337 GND 0.001802f
C3104 VDD.n2338 GND 0.006612f
C3105 VDD.n2339 GND 0.006442f
C3106 VDD.n2340 GND 0.001802f
C3107 VDD.n2341 GND 0.006442f
C3108 VDD.n2342 GND 0.264647f
C3109 VDD.n2343 GND 0.177615f
C3110 VDD.n2344 GND 0.113674f
C3111 VDD.n2345 GND 0.002697f
C3112 VDD.n2346 GND 0.002171f
C3113 VDD.n2347 GND 0.002171f
C3114 VDD.n2348 GND 0.002171f
C3115 VDD.n2349 GND 0.002697f
C3116 VDD.n2350 GND 0.177615f
C3117 VDD.n2351 GND 0.177615f
C3118 VDD.n2352 GND 0.177615f
C3119 VDD.n2353 GND 0.002697f
C3120 VDD.n2354 GND 0.002171f
C3121 VDD.n2355 GND 0.002171f
C3122 VDD.n2356 GND 0.002171f
C3123 VDD.n2357 GND 0.002697f
C3124 VDD.n2358 GND 0.177615f
C3125 VDD.n2359 GND 0.101241f
C3126 VDD.t108 GND 0.088808f
C3127 VDD.n2360 GND 0.165182f
C3128 VDD.n2361 GND 0.002697f
C3129 VDD.n2362 GND 0.002171f
C3130 VDD.n2363 GND 0.002171f
C3131 VDD.n2364 GND 0.002171f
C3132 VDD.n2365 GND 0.002697f
C3133 VDD.n2366 GND 0.177615f
C3134 VDD.n2367 GND 0.16163f
C3135 VDD.t90 GND 0.088808f
C3136 VDD.n2368 GND 0.104793f
C3137 VDD.n2369 GND 0.002697f
C3138 VDD.n2370 GND 0.002171f
C3139 VDD.n2371 GND 0.002171f
C3140 VDD.n2372 GND 0.002171f
C3141 VDD.n2373 GND 0.002697f
C3142 VDD.n2374 GND 0.177615f
C3143 VDD.n2375 GND 0.177615f
C3144 VDD.n2376 GND 0.133211f
C3145 VDD.n2377 GND 0.002697f
C3146 VDD.n2378 GND 0.002171f
C3147 VDD.n2379 GND 0.002073f
C3148 VDD.n2380 GND 0.068919f
C3149 VDD.n2381 GND 0.676176f
.ends

