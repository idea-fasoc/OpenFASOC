* NGSPICE file created from diff_pair_sample_0475.ext - technology: sky130A

.subckt diff_pair_sample_0475 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t15 w_n1966_n1882# sky130_fd_pr__pfet_01v8 ad=1.7823 pd=9.92 as=0.75405 ps=4.9 w=4.57 l=0.5
X1 VDD2.t9 VN.t0 VTAIL.t7 w_n1966_n1882# sky130_fd_pr__pfet_01v8 ad=1.7823 pd=9.92 as=0.75405 ps=4.9 w=4.57 l=0.5
X2 VDD2.t8 VN.t1 VTAIL.t9 w_n1966_n1882# sky130_fd_pr__pfet_01v8 ad=0.75405 pd=4.9 as=0.75405 ps=4.9 w=4.57 l=0.5
X3 VTAIL.t10 VP.t1 VDD1.t8 w_n1966_n1882# sky130_fd_pr__pfet_01v8 ad=0.75405 pd=4.9 as=0.75405 ps=4.9 w=4.57 l=0.5
X4 B.t11 B.t9 B.t10 w_n1966_n1882# sky130_fd_pr__pfet_01v8 ad=1.7823 pd=9.92 as=0 ps=0 w=4.57 l=0.5
X5 B.t8 B.t6 B.t7 w_n1966_n1882# sky130_fd_pr__pfet_01v8 ad=1.7823 pd=9.92 as=0 ps=0 w=4.57 l=0.5
X6 VDD1.t7 VP.t2 VTAIL.t13 w_n1966_n1882# sky130_fd_pr__pfet_01v8 ad=0.75405 pd=4.9 as=1.7823 ps=9.92 w=4.57 l=0.5
X7 VTAIL.t18 VP.t3 VDD1.t6 w_n1966_n1882# sky130_fd_pr__pfet_01v8 ad=0.75405 pd=4.9 as=0.75405 ps=4.9 w=4.57 l=0.5
X8 VDD2.t7 VN.t2 VTAIL.t8 w_n1966_n1882# sky130_fd_pr__pfet_01v8 ad=0.75405 pd=4.9 as=1.7823 ps=9.92 w=4.57 l=0.5
X9 VDD1.t5 VP.t4 VTAIL.t16 w_n1966_n1882# sky130_fd_pr__pfet_01v8 ad=1.7823 pd=9.92 as=0.75405 ps=4.9 w=4.57 l=0.5
X10 VTAIL.t19 VP.t5 VDD1.t4 w_n1966_n1882# sky130_fd_pr__pfet_01v8 ad=0.75405 pd=4.9 as=0.75405 ps=4.9 w=4.57 l=0.5
X11 VTAIL.t17 VP.t6 VDD1.t3 w_n1966_n1882# sky130_fd_pr__pfet_01v8 ad=0.75405 pd=4.9 as=0.75405 ps=4.9 w=4.57 l=0.5
X12 VTAIL.t3 VN.t3 VDD2.t6 w_n1966_n1882# sky130_fd_pr__pfet_01v8 ad=0.75405 pd=4.9 as=0.75405 ps=4.9 w=4.57 l=0.5
X13 VDD2.t5 VN.t4 VTAIL.t5 w_n1966_n1882# sky130_fd_pr__pfet_01v8 ad=1.7823 pd=9.92 as=0.75405 ps=4.9 w=4.57 l=0.5
X14 VTAIL.t6 VN.t5 VDD2.t4 w_n1966_n1882# sky130_fd_pr__pfet_01v8 ad=0.75405 pd=4.9 as=0.75405 ps=4.9 w=4.57 l=0.5
X15 B.t5 B.t3 B.t4 w_n1966_n1882# sky130_fd_pr__pfet_01v8 ad=1.7823 pd=9.92 as=0 ps=0 w=4.57 l=0.5
X16 VDD1.t2 VP.t7 VTAIL.t12 w_n1966_n1882# sky130_fd_pr__pfet_01v8 ad=0.75405 pd=4.9 as=1.7823 ps=9.92 w=4.57 l=0.5
X17 VDD1.t1 VP.t8 VTAIL.t14 w_n1966_n1882# sky130_fd_pr__pfet_01v8 ad=0.75405 pd=4.9 as=0.75405 ps=4.9 w=4.57 l=0.5
X18 VDD2.t3 VN.t6 VTAIL.t0 w_n1966_n1882# sky130_fd_pr__pfet_01v8 ad=0.75405 pd=4.9 as=1.7823 ps=9.92 w=4.57 l=0.5
X19 VDD1.t0 VP.t9 VTAIL.t11 w_n1966_n1882# sky130_fd_pr__pfet_01v8 ad=0.75405 pd=4.9 as=0.75405 ps=4.9 w=4.57 l=0.5
X20 B.t2 B.t0 B.t1 w_n1966_n1882# sky130_fd_pr__pfet_01v8 ad=1.7823 pd=9.92 as=0 ps=0 w=4.57 l=0.5
X21 VTAIL.t1 VN.t7 VDD2.t2 w_n1966_n1882# sky130_fd_pr__pfet_01v8 ad=0.75405 pd=4.9 as=0.75405 ps=4.9 w=4.57 l=0.5
X22 VTAIL.t2 VN.t8 VDD2.t1 w_n1966_n1882# sky130_fd_pr__pfet_01v8 ad=0.75405 pd=4.9 as=0.75405 ps=4.9 w=4.57 l=0.5
X23 VDD2.t0 VN.t9 VTAIL.t4 w_n1966_n1882# sky130_fd_pr__pfet_01v8 ad=0.75405 pd=4.9 as=0.75405 ps=4.9 w=4.57 l=0.5
R0 VP.n5 VP.t0 320.305
R1 VP.n16 VP.t4 299.322
R2 VP.n17 VP.t6 299.322
R3 VP.n1 VP.t9 299.322
R4 VP.n23 VP.t3 299.322
R5 VP.n24 VP.t2 299.322
R6 VP.n13 VP.t7 299.322
R7 VP.n12 VP.t1 299.322
R8 VP.n4 VP.t8 299.322
R9 VP.n6 VP.t5 299.322
R10 VP.n25 VP.n24 161.3
R11 VP.n8 VP.n7 161.3
R12 VP.n9 VP.n4 161.3
R13 VP.n11 VP.n10 161.3
R14 VP.n12 VP.n3 161.3
R15 VP.n14 VP.n13 161.3
R16 VP.n23 VP.n0 161.3
R17 VP.n22 VP.n21 161.3
R18 VP.n20 VP.n1 161.3
R19 VP.n19 VP.n18 161.3
R20 VP.n17 VP.n2 161.3
R21 VP.n16 VP.n15 161.3
R22 VP.n8 VP.n5 70.4033
R23 VP.n17 VP.n16 48.2005
R24 VP.n24 VP.n23 48.2005
R25 VP.n13 VP.n12 48.2005
R26 VP.n18 VP.n1 36.5157
R27 VP.n22 VP.n1 36.5157
R28 VP.n11 VP.n4 36.5157
R29 VP.n7 VP.n4 36.5157
R30 VP.n15 VP.n14 36.0952
R31 VP.n6 VP.n5 20.9576
R32 VP.n18 VP.n17 11.6853
R33 VP.n23 VP.n22 11.6853
R34 VP.n12 VP.n11 11.6853
R35 VP.n7 VP.n6 11.6853
R36 VP.n9 VP.n8 0.189894
R37 VP.n10 VP.n9 0.189894
R38 VP.n10 VP.n3 0.189894
R39 VP.n14 VP.n3 0.189894
R40 VP.n15 VP.n2 0.189894
R41 VP.n19 VP.n2 0.189894
R42 VP.n20 VP.n19 0.189894
R43 VP.n21 VP.n20 0.189894
R44 VP.n21 VP.n0 0.189894
R45 VP.n25 VP.n0 0.189894
R46 VP VP.n25 0.0516364
R47 VTAIL.n104 VTAIL.n86 756.745
R48 VTAIL.n20 VTAIL.n2 756.745
R49 VTAIL.n80 VTAIL.n62 756.745
R50 VTAIL.n52 VTAIL.n34 756.745
R51 VTAIL.n95 VTAIL.n94 585
R52 VTAIL.n97 VTAIL.n96 585
R53 VTAIL.n90 VTAIL.n89 585
R54 VTAIL.n103 VTAIL.n102 585
R55 VTAIL.n105 VTAIL.n104 585
R56 VTAIL.n11 VTAIL.n10 585
R57 VTAIL.n13 VTAIL.n12 585
R58 VTAIL.n6 VTAIL.n5 585
R59 VTAIL.n19 VTAIL.n18 585
R60 VTAIL.n21 VTAIL.n20 585
R61 VTAIL.n81 VTAIL.n80 585
R62 VTAIL.n79 VTAIL.n78 585
R63 VTAIL.n66 VTAIL.n65 585
R64 VTAIL.n73 VTAIL.n72 585
R65 VTAIL.n71 VTAIL.n70 585
R66 VTAIL.n53 VTAIL.n52 585
R67 VTAIL.n51 VTAIL.n50 585
R68 VTAIL.n38 VTAIL.n37 585
R69 VTAIL.n45 VTAIL.n44 585
R70 VTAIL.n43 VTAIL.n42 585
R71 VTAIL.n93 VTAIL.t0 328.587
R72 VTAIL.n9 VTAIL.t13 328.587
R73 VTAIL.n69 VTAIL.t12 328.587
R74 VTAIL.n41 VTAIL.t8 328.587
R75 VTAIL.n96 VTAIL.n95 171.744
R76 VTAIL.n96 VTAIL.n89 171.744
R77 VTAIL.n103 VTAIL.n89 171.744
R78 VTAIL.n104 VTAIL.n103 171.744
R79 VTAIL.n12 VTAIL.n11 171.744
R80 VTAIL.n12 VTAIL.n5 171.744
R81 VTAIL.n19 VTAIL.n5 171.744
R82 VTAIL.n20 VTAIL.n19 171.744
R83 VTAIL.n80 VTAIL.n79 171.744
R84 VTAIL.n79 VTAIL.n65 171.744
R85 VTAIL.n72 VTAIL.n65 171.744
R86 VTAIL.n72 VTAIL.n71 171.744
R87 VTAIL.n52 VTAIL.n51 171.744
R88 VTAIL.n51 VTAIL.n37 171.744
R89 VTAIL.n44 VTAIL.n37 171.744
R90 VTAIL.n44 VTAIL.n43 171.744
R91 VTAIL.n61 VTAIL.n60 87.595
R92 VTAIL.n59 VTAIL.n58 87.595
R93 VTAIL.n33 VTAIL.n32 87.595
R94 VTAIL.n31 VTAIL.n30 87.595
R95 VTAIL.n111 VTAIL.n110 87.5948
R96 VTAIL.n1 VTAIL.n0 87.5948
R97 VTAIL.n27 VTAIL.n26 87.5948
R98 VTAIL.n29 VTAIL.n28 87.5948
R99 VTAIL.n95 VTAIL.t0 85.8723
R100 VTAIL.n11 VTAIL.t13 85.8723
R101 VTAIL.n71 VTAIL.t12 85.8723
R102 VTAIL.n43 VTAIL.t8 85.8723
R103 VTAIL.n109 VTAIL.n108 32.3793
R104 VTAIL.n25 VTAIL.n24 32.3793
R105 VTAIL.n85 VTAIL.n84 32.3793
R106 VTAIL.n57 VTAIL.n56 32.3793
R107 VTAIL.n31 VTAIL.n29 17.7376
R108 VTAIL.n109 VTAIL.n85 17.0221
R109 VTAIL.n94 VTAIL.n93 16.3651
R110 VTAIL.n10 VTAIL.n9 16.3651
R111 VTAIL.n70 VTAIL.n69 16.3651
R112 VTAIL.n42 VTAIL.n41 16.3651
R113 VTAIL.n97 VTAIL.n92 12.8005
R114 VTAIL.n13 VTAIL.n8 12.8005
R115 VTAIL.n73 VTAIL.n68 12.8005
R116 VTAIL.n45 VTAIL.n40 12.8005
R117 VTAIL.n98 VTAIL.n90 12.0247
R118 VTAIL.n14 VTAIL.n6 12.0247
R119 VTAIL.n74 VTAIL.n66 12.0247
R120 VTAIL.n46 VTAIL.n38 12.0247
R121 VTAIL.n102 VTAIL.n101 11.249
R122 VTAIL.n18 VTAIL.n17 11.249
R123 VTAIL.n78 VTAIL.n77 11.249
R124 VTAIL.n50 VTAIL.n49 11.249
R125 VTAIL.n105 VTAIL.n88 10.4732
R126 VTAIL.n21 VTAIL.n4 10.4732
R127 VTAIL.n81 VTAIL.n64 10.4732
R128 VTAIL.n53 VTAIL.n36 10.4732
R129 VTAIL.n106 VTAIL.n86 9.69747
R130 VTAIL.n22 VTAIL.n2 9.69747
R131 VTAIL.n82 VTAIL.n62 9.69747
R132 VTAIL.n54 VTAIL.n34 9.69747
R133 VTAIL.n108 VTAIL.n107 9.45567
R134 VTAIL.n24 VTAIL.n23 9.45567
R135 VTAIL.n84 VTAIL.n83 9.45567
R136 VTAIL.n56 VTAIL.n55 9.45567
R137 VTAIL.n107 VTAIL.n106 9.3005
R138 VTAIL.n88 VTAIL.n87 9.3005
R139 VTAIL.n101 VTAIL.n100 9.3005
R140 VTAIL.n99 VTAIL.n98 9.3005
R141 VTAIL.n92 VTAIL.n91 9.3005
R142 VTAIL.n23 VTAIL.n22 9.3005
R143 VTAIL.n4 VTAIL.n3 9.3005
R144 VTAIL.n17 VTAIL.n16 9.3005
R145 VTAIL.n15 VTAIL.n14 9.3005
R146 VTAIL.n8 VTAIL.n7 9.3005
R147 VTAIL.n83 VTAIL.n82 9.3005
R148 VTAIL.n64 VTAIL.n63 9.3005
R149 VTAIL.n77 VTAIL.n76 9.3005
R150 VTAIL.n75 VTAIL.n74 9.3005
R151 VTAIL.n68 VTAIL.n67 9.3005
R152 VTAIL.n55 VTAIL.n54 9.3005
R153 VTAIL.n36 VTAIL.n35 9.3005
R154 VTAIL.n49 VTAIL.n48 9.3005
R155 VTAIL.n47 VTAIL.n46 9.3005
R156 VTAIL.n40 VTAIL.n39 9.3005
R157 VTAIL.n110 VTAIL.t4 7.11319
R158 VTAIL.n110 VTAIL.t2 7.11319
R159 VTAIL.n0 VTAIL.t5 7.11319
R160 VTAIL.n0 VTAIL.t3 7.11319
R161 VTAIL.n26 VTAIL.t11 7.11319
R162 VTAIL.n26 VTAIL.t18 7.11319
R163 VTAIL.n28 VTAIL.t16 7.11319
R164 VTAIL.n28 VTAIL.t17 7.11319
R165 VTAIL.n60 VTAIL.t14 7.11319
R166 VTAIL.n60 VTAIL.t10 7.11319
R167 VTAIL.n58 VTAIL.t15 7.11319
R168 VTAIL.n58 VTAIL.t19 7.11319
R169 VTAIL.n32 VTAIL.t9 7.11319
R170 VTAIL.n32 VTAIL.t1 7.11319
R171 VTAIL.n30 VTAIL.t7 7.11319
R172 VTAIL.n30 VTAIL.t6 7.11319
R173 VTAIL.n108 VTAIL.n86 4.26717
R174 VTAIL.n24 VTAIL.n2 4.26717
R175 VTAIL.n84 VTAIL.n62 4.26717
R176 VTAIL.n56 VTAIL.n34 4.26717
R177 VTAIL.n93 VTAIL.n91 3.73474
R178 VTAIL.n9 VTAIL.n7 3.73474
R179 VTAIL.n69 VTAIL.n67 3.73474
R180 VTAIL.n41 VTAIL.n39 3.73474
R181 VTAIL.n106 VTAIL.n105 3.49141
R182 VTAIL.n22 VTAIL.n21 3.49141
R183 VTAIL.n82 VTAIL.n81 3.49141
R184 VTAIL.n54 VTAIL.n53 3.49141
R185 VTAIL.n102 VTAIL.n88 2.71565
R186 VTAIL.n18 VTAIL.n4 2.71565
R187 VTAIL.n78 VTAIL.n64 2.71565
R188 VTAIL.n50 VTAIL.n36 2.71565
R189 VTAIL.n101 VTAIL.n90 1.93989
R190 VTAIL.n17 VTAIL.n6 1.93989
R191 VTAIL.n77 VTAIL.n66 1.93989
R192 VTAIL.n49 VTAIL.n38 1.93989
R193 VTAIL.n98 VTAIL.n97 1.16414
R194 VTAIL.n14 VTAIL.n13 1.16414
R195 VTAIL.n74 VTAIL.n73 1.16414
R196 VTAIL.n46 VTAIL.n45 1.16414
R197 VTAIL.n59 VTAIL.n57 0.828086
R198 VTAIL.n25 VTAIL.n1 0.828086
R199 VTAIL.n33 VTAIL.n31 0.716017
R200 VTAIL.n57 VTAIL.n33 0.716017
R201 VTAIL.n61 VTAIL.n59 0.716017
R202 VTAIL.n85 VTAIL.n61 0.716017
R203 VTAIL.n29 VTAIL.n27 0.716017
R204 VTAIL.n27 VTAIL.n25 0.716017
R205 VTAIL.n111 VTAIL.n109 0.716017
R206 VTAIL VTAIL.n1 0.595328
R207 VTAIL.n94 VTAIL.n92 0.388379
R208 VTAIL.n10 VTAIL.n8 0.388379
R209 VTAIL.n70 VTAIL.n68 0.388379
R210 VTAIL.n42 VTAIL.n40 0.388379
R211 VTAIL.n99 VTAIL.n91 0.155672
R212 VTAIL.n100 VTAIL.n99 0.155672
R213 VTAIL.n100 VTAIL.n87 0.155672
R214 VTAIL.n107 VTAIL.n87 0.155672
R215 VTAIL.n15 VTAIL.n7 0.155672
R216 VTAIL.n16 VTAIL.n15 0.155672
R217 VTAIL.n16 VTAIL.n3 0.155672
R218 VTAIL.n23 VTAIL.n3 0.155672
R219 VTAIL.n83 VTAIL.n63 0.155672
R220 VTAIL.n76 VTAIL.n63 0.155672
R221 VTAIL.n76 VTAIL.n75 0.155672
R222 VTAIL.n75 VTAIL.n67 0.155672
R223 VTAIL.n55 VTAIL.n35 0.155672
R224 VTAIL.n48 VTAIL.n35 0.155672
R225 VTAIL.n48 VTAIL.n47 0.155672
R226 VTAIL.n47 VTAIL.n39 0.155672
R227 VTAIL VTAIL.n111 0.12119
R228 VDD1.n18 VDD1.n0 756.745
R229 VDD1.n43 VDD1.n25 756.745
R230 VDD1.n19 VDD1.n18 585
R231 VDD1.n17 VDD1.n16 585
R232 VDD1.n4 VDD1.n3 585
R233 VDD1.n11 VDD1.n10 585
R234 VDD1.n9 VDD1.n8 585
R235 VDD1.n34 VDD1.n33 585
R236 VDD1.n36 VDD1.n35 585
R237 VDD1.n29 VDD1.n28 585
R238 VDD1.n42 VDD1.n41 585
R239 VDD1.n44 VDD1.n43 585
R240 VDD1.n7 VDD1.t9 328.587
R241 VDD1.n32 VDD1.t5 328.587
R242 VDD1.n18 VDD1.n17 171.744
R243 VDD1.n17 VDD1.n3 171.744
R244 VDD1.n10 VDD1.n3 171.744
R245 VDD1.n10 VDD1.n9 171.744
R246 VDD1.n35 VDD1.n34 171.744
R247 VDD1.n35 VDD1.n28 171.744
R248 VDD1.n42 VDD1.n28 171.744
R249 VDD1.n43 VDD1.n42 171.744
R250 VDD1.n51 VDD1.n50 104.754
R251 VDD1.n24 VDD1.n23 104.273
R252 VDD1.n53 VDD1.n52 104.273
R253 VDD1.n49 VDD1.n48 104.273
R254 VDD1.n9 VDD1.t9 85.8723
R255 VDD1.n34 VDD1.t5 85.8723
R256 VDD1.n24 VDD1.n22 49.7736
R257 VDD1.n49 VDD1.n47 49.7736
R258 VDD1.n53 VDD1.n51 31.9944
R259 VDD1.n8 VDD1.n7 16.3651
R260 VDD1.n33 VDD1.n32 16.3651
R261 VDD1.n11 VDD1.n6 12.8005
R262 VDD1.n36 VDD1.n31 12.8005
R263 VDD1.n12 VDD1.n4 12.0247
R264 VDD1.n37 VDD1.n29 12.0247
R265 VDD1.n16 VDD1.n15 11.249
R266 VDD1.n41 VDD1.n40 11.249
R267 VDD1.n19 VDD1.n2 10.4732
R268 VDD1.n44 VDD1.n27 10.4732
R269 VDD1.n20 VDD1.n0 9.69747
R270 VDD1.n45 VDD1.n25 9.69747
R271 VDD1.n22 VDD1.n21 9.45567
R272 VDD1.n47 VDD1.n46 9.45567
R273 VDD1.n21 VDD1.n20 9.3005
R274 VDD1.n2 VDD1.n1 9.3005
R275 VDD1.n15 VDD1.n14 9.3005
R276 VDD1.n13 VDD1.n12 9.3005
R277 VDD1.n6 VDD1.n5 9.3005
R278 VDD1.n46 VDD1.n45 9.3005
R279 VDD1.n27 VDD1.n26 9.3005
R280 VDD1.n40 VDD1.n39 9.3005
R281 VDD1.n38 VDD1.n37 9.3005
R282 VDD1.n31 VDD1.n30 9.3005
R283 VDD1.n52 VDD1.t8 7.11319
R284 VDD1.n52 VDD1.t2 7.11319
R285 VDD1.n23 VDD1.t4 7.11319
R286 VDD1.n23 VDD1.t1 7.11319
R287 VDD1.n50 VDD1.t6 7.11319
R288 VDD1.n50 VDD1.t7 7.11319
R289 VDD1.n48 VDD1.t3 7.11319
R290 VDD1.n48 VDD1.t0 7.11319
R291 VDD1.n22 VDD1.n0 4.26717
R292 VDD1.n47 VDD1.n25 4.26717
R293 VDD1.n7 VDD1.n5 3.73474
R294 VDD1.n32 VDD1.n30 3.73474
R295 VDD1.n20 VDD1.n19 3.49141
R296 VDD1.n45 VDD1.n44 3.49141
R297 VDD1.n16 VDD1.n2 2.71565
R298 VDD1.n41 VDD1.n27 2.71565
R299 VDD1.n15 VDD1.n4 1.93989
R300 VDD1.n40 VDD1.n29 1.93989
R301 VDD1.n12 VDD1.n11 1.16414
R302 VDD1.n37 VDD1.n36 1.16414
R303 VDD1 VDD1.n53 0.478948
R304 VDD1.n8 VDD1.n6 0.388379
R305 VDD1.n33 VDD1.n31 0.388379
R306 VDD1 VDD1.n24 0.237569
R307 VDD1.n21 VDD1.n1 0.155672
R308 VDD1.n14 VDD1.n1 0.155672
R309 VDD1.n14 VDD1.n13 0.155672
R310 VDD1.n13 VDD1.n5 0.155672
R311 VDD1.n38 VDD1.n30 0.155672
R312 VDD1.n39 VDD1.n38 0.155672
R313 VDD1.n39 VDD1.n26 0.155672
R314 VDD1.n46 VDD1.n26 0.155672
R315 VDD1.n51 VDD1.n49 0.124033
R316 VN.n2 VN.t4 320.305
R317 VN.n14 VN.t2 320.305
R318 VN.n3 VN.t3 299.322
R319 VN.n1 VN.t9 299.322
R320 VN.n9 VN.t8 299.322
R321 VN.n10 VN.t6 299.322
R322 VN.n15 VN.t7 299.322
R323 VN.n13 VN.t1 299.322
R324 VN.n21 VN.t5 299.322
R325 VN.n22 VN.t0 299.322
R326 VN.n11 VN.n10 161.3
R327 VN.n23 VN.n22 161.3
R328 VN.n21 VN.n12 161.3
R329 VN.n20 VN.n19 161.3
R330 VN.n18 VN.n13 161.3
R331 VN.n17 VN.n16 161.3
R332 VN.n9 VN.n0 161.3
R333 VN.n8 VN.n7 161.3
R334 VN.n6 VN.n1 161.3
R335 VN.n5 VN.n4 161.3
R336 VN.n17 VN.n14 70.4033
R337 VN.n5 VN.n2 70.4033
R338 VN.n10 VN.n9 48.2005
R339 VN.n22 VN.n21 48.2005
R340 VN.n4 VN.n1 36.5157
R341 VN.n8 VN.n1 36.5157
R342 VN.n16 VN.n13 36.5157
R343 VN.n20 VN.n13 36.5157
R344 VN VN.n23 36.4759
R345 VN.n15 VN.n14 20.9576
R346 VN.n3 VN.n2 20.9576
R347 VN.n4 VN.n3 11.6853
R348 VN.n9 VN.n8 11.6853
R349 VN.n16 VN.n15 11.6853
R350 VN.n21 VN.n20 11.6853
R351 VN.n23 VN.n12 0.189894
R352 VN.n19 VN.n12 0.189894
R353 VN.n19 VN.n18 0.189894
R354 VN.n18 VN.n17 0.189894
R355 VN.n6 VN.n5 0.189894
R356 VN.n7 VN.n6 0.189894
R357 VN.n7 VN.n0 0.189894
R358 VN.n11 VN.n0 0.189894
R359 VN VN.n11 0.0516364
R360 VDD2.n45 VDD2.n27 756.745
R361 VDD2.n18 VDD2.n0 756.745
R362 VDD2.n46 VDD2.n45 585
R363 VDD2.n44 VDD2.n43 585
R364 VDD2.n31 VDD2.n30 585
R365 VDD2.n38 VDD2.n37 585
R366 VDD2.n36 VDD2.n35 585
R367 VDD2.n9 VDD2.n8 585
R368 VDD2.n11 VDD2.n10 585
R369 VDD2.n4 VDD2.n3 585
R370 VDD2.n17 VDD2.n16 585
R371 VDD2.n19 VDD2.n18 585
R372 VDD2.n34 VDD2.t9 328.587
R373 VDD2.n7 VDD2.t5 328.587
R374 VDD2.n45 VDD2.n44 171.744
R375 VDD2.n44 VDD2.n30 171.744
R376 VDD2.n37 VDD2.n30 171.744
R377 VDD2.n37 VDD2.n36 171.744
R378 VDD2.n10 VDD2.n9 171.744
R379 VDD2.n10 VDD2.n3 171.744
R380 VDD2.n17 VDD2.n3 171.744
R381 VDD2.n18 VDD2.n17 171.744
R382 VDD2.n26 VDD2.n25 104.754
R383 VDD2 VDD2.n53 104.752
R384 VDD2.n52 VDD2.n51 104.273
R385 VDD2.n24 VDD2.n23 104.273
R386 VDD2.n36 VDD2.t9 85.8723
R387 VDD2.n9 VDD2.t5 85.8723
R388 VDD2.n24 VDD2.n22 49.7736
R389 VDD2.n50 VDD2.n49 49.0581
R390 VDD2.n50 VDD2.n26 31.0537
R391 VDD2.n35 VDD2.n34 16.3651
R392 VDD2.n8 VDD2.n7 16.3651
R393 VDD2.n38 VDD2.n33 12.8005
R394 VDD2.n11 VDD2.n6 12.8005
R395 VDD2.n39 VDD2.n31 12.0247
R396 VDD2.n12 VDD2.n4 12.0247
R397 VDD2.n43 VDD2.n42 11.249
R398 VDD2.n16 VDD2.n15 11.249
R399 VDD2.n46 VDD2.n29 10.4732
R400 VDD2.n19 VDD2.n2 10.4732
R401 VDD2.n47 VDD2.n27 9.69747
R402 VDD2.n20 VDD2.n0 9.69747
R403 VDD2.n49 VDD2.n48 9.45567
R404 VDD2.n22 VDD2.n21 9.45567
R405 VDD2.n48 VDD2.n47 9.3005
R406 VDD2.n29 VDD2.n28 9.3005
R407 VDD2.n42 VDD2.n41 9.3005
R408 VDD2.n40 VDD2.n39 9.3005
R409 VDD2.n33 VDD2.n32 9.3005
R410 VDD2.n21 VDD2.n20 9.3005
R411 VDD2.n2 VDD2.n1 9.3005
R412 VDD2.n15 VDD2.n14 9.3005
R413 VDD2.n13 VDD2.n12 9.3005
R414 VDD2.n6 VDD2.n5 9.3005
R415 VDD2.n53 VDD2.t2 7.11319
R416 VDD2.n53 VDD2.t7 7.11319
R417 VDD2.n51 VDD2.t4 7.11319
R418 VDD2.n51 VDD2.t8 7.11319
R419 VDD2.n25 VDD2.t1 7.11319
R420 VDD2.n25 VDD2.t3 7.11319
R421 VDD2.n23 VDD2.t6 7.11319
R422 VDD2.n23 VDD2.t0 7.11319
R423 VDD2.n49 VDD2.n27 4.26717
R424 VDD2.n22 VDD2.n0 4.26717
R425 VDD2.n34 VDD2.n32 3.73474
R426 VDD2.n7 VDD2.n5 3.73474
R427 VDD2.n47 VDD2.n46 3.49141
R428 VDD2.n20 VDD2.n19 3.49141
R429 VDD2.n43 VDD2.n29 2.71565
R430 VDD2.n16 VDD2.n2 2.71565
R431 VDD2.n42 VDD2.n31 1.93989
R432 VDD2.n15 VDD2.n4 1.93989
R433 VDD2.n39 VDD2.n38 1.16414
R434 VDD2.n12 VDD2.n11 1.16414
R435 VDD2.n52 VDD2.n50 0.716017
R436 VDD2.n35 VDD2.n33 0.388379
R437 VDD2.n8 VDD2.n6 0.388379
R438 VDD2 VDD2.n52 0.237569
R439 VDD2.n48 VDD2.n28 0.155672
R440 VDD2.n41 VDD2.n28 0.155672
R441 VDD2.n41 VDD2.n40 0.155672
R442 VDD2.n40 VDD2.n32 0.155672
R443 VDD2.n13 VDD2.n5 0.155672
R444 VDD2.n14 VDD2.n13 0.155672
R445 VDD2.n14 VDD2.n1 0.155672
R446 VDD2.n21 VDD2.n1 0.155672
R447 VDD2.n26 VDD2.n24 0.124033
R448 B.n210 B.n209 585
R449 B.n208 B.n65 585
R450 B.n207 B.n206 585
R451 B.n205 B.n66 585
R452 B.n204 B.n203 585
R453 B.n202 B.n67 585
R454 B.n201 B.n200 585
R455 B.n199 B.n68 585
R456 B.n198 B.n197 585
R457 B.n196 B.n69 585
R458 B.n195 B.n194 585
R459 B.n193 B.n70 585
R460 B.n192 B.n191 585
R461 B.n190 B.n71 585
R462 B.n189 B.n188 585
R463 B.n187 B.n72 585
R464 B.n186 B.n185 585
R465 B.n184 B.n73 585
R466 B.n183 B.n182 585
R467 B.n181 B.n74 585
R468 B.n180 B.n179 585
R469 B.n175 B.n75 585
R470 B.n174 B.n173 585
R471 B.n172 B.n76 585
R472 B.n171 B.n170 585
R473 B.n169 B.n77 585
R474 B.n168 B.n167 585
R475 B.n166 B.n78 585
R476 B.n165 B.n164 585
R477 B.n162 B.n79 585
R478 B.n161 B.n160 585
R479 B.n159 B.n82 585
R480 B.n158 B.n157 585
R481 B.n156 B.n83 585
R482 B.n155 B.n154 585
R483 B.n153 B.n84 585
R484 B.n152 B.n151 585
R485 B.n150 B.n85 585
R486 B.n149 B.n148 585
R487 B.n147 B.n86 585
R488 B.n146 B.n145 585
R489 B.n144 B.n87 585
R490 B.n143 B.n142 585
R491 B.n141 B.n88 585
R492 B.n140 B.n139 585
R493 B.n138 B.n89 585
R494 B.n137 B.n136 585
R495 B.n135 B.n90 585
R496 B.n134 B.n133 585
R497 B.n211 B.n64 585
R498 B.n213 B.n212 585
R499 B.n214 B.n63 585
R500 B.n216 B.n215 585
R501 B.n217 B.n62 585
R502 B.n219 B.n218 585
R503 B.n220 B.n61 585
R504 B.n222 B.n221 585
R505 B.n223 B.n60 585
R506 B.n225 B.n224 585
R507 B.n226 B.n59 585
R508 B.n228 B.n227 585
R509 B.n229 B.n58 585
R510 B.n231 B.n230 585
R511 B.n232 B.n57 585
R512 B.n234 B.n233 585
R513 B.n235 B.n56 585
R514 B.n237 B.n236 585
R515 B.n238 B.n55 585
R516 B.n240 B.n239 585
R517 B.n241 B.n54 585
R518 B.n243 B.n242 585
R519 B.n244 B.n53 585
R520 B.n246 B.n245 585
R521 B.n247 B.n52 585
R522 B.n249 B.n248 585
R523 B.n250 B.n51 585
R524 B.n252 B.n251 585
R525 B.n253 B.n50 585
R526 B.n255 B.n254 585
R527 B.n256 B.n49 585
R528 B.n258 B.n257 585
R529 B.n259 B.n48 585
R530 B.n261 B.n260 585
R531 B.n262 B.n47 585
R532 B.n264 B.n263 585
R533 B.n265 B.n46 585
R534 B.n267 B.n266 585
R535 B.n268 B.n45 585
R536 B.n270 B.n269 585
R537 B.n271 B.n44 585
R538 B.n273 B.n272 585
R539 B.n274 B.n43 585
R540 B.n276 B.n275 585
R541 B.n277 B.n42 585
R542 B.n279 B.n278 585
R543 B.n354 B.n13 585
R544 B.n353 B.n352 585
R545 B.n351 B.n14 585
R546 B.n350 B.n349 585
R547 B.n348 B.n15 585
R548 B.n347 B.n346 585
R549 B.n345 B.n16 585
R550 B.n344 B.n343 585
R551 B.n342 B.n17 585
R552 B.n341 B.n340 585
R553 B.n339 B.n18 585
R554 B.n338 B.n337 585
R555 B.n336 B.n19 585
R556 B.n335 B.n334 585
R557 B.n333 B.n20 585
R558 B.n332 B.n331 585
R559 B.n330 B.n21 585
R560 B.n329 B.n328 585
R561 B.n327 B.n22 585
R562 B.n326 B.n325 585
R563 B.n323 B.n23 585
R564 B.n322 B.n321 585
R565 B.n320 B.n26 585
R566 B.n319 B.n318 585
R567 B.n317 B.n27 585
R568 B.n316 B.n315 585
R569 B.n314 B.n28 585
R570 B.n313 B.n312 585
R571 B.n311 B.n29 585
R572 B.n309 B.n308 585
R573 B.n307 B.n32 585
R574 B.n306 B.n305 585
R575 B.n304 B.n33 585
R576 B.n303 B.n302 585
R577 B.n301 B.n34 585
R578 B.n300 B.n299 585
R579 B.n298 B.n35 585
R580 B.n297 B.n296 585
R581 B.n295 B.n36 585
R582 B.n294 B.n293 585
R583 B.n292 B.n37 585
R584 B.n291 B.n290 585
R585 B.n289 B.n38 585
R586 B.n288 B.n287 585
R587 B.n286 B.n39 585
R588 B.n285 B.n284 585
R589 B.n283 B.n40 585
R590 B.n282 B.n281 585
R591 B.n280 B.n41 585
R592 B.n356 B.n355 585
R593 B.n357 B.n12 585
R594 B.n359 B.n358 585
R595 B.n360 B.n11 585
R596 B.n362 B.n361 585
R597 B.n363 B.n10 585
R598 B.n365 B.n364 585
R599 B.n366 B.n9 585
R600 B.n368 B.n367 585
R601 B.n369 B.n8 585
R602 B.n371 B.n370 585
R603 B.n372 B.n7 585
R604 B.n374 B.n373 585
R605 B.n375 B.n6 585
R606 B.n377 B.n376 585
R607 B.n378 B.n5 585
R608 B.n380 B.n379 585
R609 B.n381 B.n4 585
R610 B.n383 B.n382 585
R611 B.n384 B.n3 585
R612 B.n386 B.n385 585
R613 B.n387 B.n0 585
R614 B.n2 B.n1 585
R615 B.n102 B.n101 585
R616 B.n104 B.n103 585
R617 B.n105 B.n100 585
R618 B.n107 B.n106 585
R619 B.n108 B.n99 585
R620 B.n110 B.n109 585
R621 B.n111 B.n98 585
R622 B.n113 B.n112 585
R623 B.n114 B.n97 585
R624 B.n116 B.n115 585
R625 B.n117 B.n96 585
R626 B.n119 B.n118 585
R627 B.n120 B.n95 585
R628 B.n122 B.n121 585
R629 B.n123 B.n94 585
R630 B.n125 B.n124 585
R631 B.n126 B.n93 585
R632 B.n128 B.n127 585
R633 B.n129 B.n92 585
R634 B.n131 B.n130 585
R635 B.n132 B.n91 585
R636 B.n134 B.n91 550.159
R637 B.n211 B.n210 550.159
R638 B.n278 B.n41 550.159
R639 B.n356 B.n13 550.159
R640 B.n80 B.t6 426.683
R641 B.n176 B.t9 426.683
R642 B.n30 B.t3 426.683
R643 B.n24 B.t0 426.683
R644 B.n176 B.t10 259.86
R645 B.n30 B.t5 259.86
R646 B.n80 B.t7 259.86
R647 B.n24 B.t2 259.86
R648 B.n389 B.n388 256.663
R649 B.n177 B.t11 243.762
R650 B.n31 B.t4 243.762
R651 B.n81 B.t8 243.762
R652 B.n25 B.t1 243.762
R653 B.n388 B.n387 235.042
R654 B.n388 B.n2 235.042
R655 B.n135 B.n134 163.367
R656 B.n136 B.n135 163.367
R657 B.n136 B.n89 163.367
R658 B.n140 B.n89 163.367
R659 B.n141 B.n140 163.367
R660 B.n142 B.n141 163.367
R661 B.n142 B.n87 163.367
R662 B.n146 B.n87 163.367
R663 B.n147 B.n146 163.367
R664 B.n148 B.n147 163.367
R665 B.n148 B.n85 163.367
R666 B.n152 B.n85 163.367
R667 B.n153 B.n152 163.367
R668 B.n154 B.n153 163.367
R669 B.n154 B.n83 163.367
R670 B.n158 B.n83 163.367
R671 B.n159 B.n158 163.367
R672 B.n160 B.n159 163.367
R673 B.n160 B.n79 163.367
R674 B.n165 B.n79 163.367
R675 B.n166 B.n165 163.367
R676 B.n167 B.n166 163.367
R677 B.n167 B.n77 163.367
R678 B.n171 B.n77 163.367
R679 B.n172 B.n171 163.367
R680 B.n173 B.n172 163.367
R681 B.n173 B.n75 163.367
R682 B.n180 B.n75 163.367
R683 B.n181 B.n180 163.367
R684 B.n182 B.n181 163.367
R685 B.n182 B.n73 163.367
R686 B.n186 B.n73 163.367
R687 B.n187 B.n186 163.367
R688 B.n188 B.n187 163.367
R689 B.n188 B.n71 163.367
R690 B.n192 B.n71 163.367
R691 B.n193 B.n192 163.367
R692 B.n194 B.n193 163.367
R693 B.n194 B.n69 163.367
R694 B.n198 B.n69 163.367
R695 B.n199 B.n198 163.367
R696 B.n200 B.n199 163.367
R697 B.n200 B.n67 163.367
R698 B.n204 B.n67 163.367
R699 B.n205 B.n204 163.367
R700 B.n206 B.n205 163.367
R701 B.n206 B.n65 163.367
R702 B.n210 B.n65 163.367
R703 B.n278 B.n277 163.367
R704 B.n277 B.n276 163.367
R705 B.n276 B.n43 163.367
R706 B.n272 B.n43 163.367
R707 B.n272 B.n271 163.367
R708 B.n271 B.n270 163.367
R709 B.n270 B.n45 163.367
R710 B.n266 B.n45 163.367
R711 B.n266 B.n265 163.367
R712 B.n265 B.n264 163.367
R713 B.n264 B.n47 163.367
R714 B.n260 B.n47 163.367
R715 B.n260 B.n259 163.367
R716 B.n259 B.n258 163.367
R717 B.n258 B.n49 163.367
R718 B.n254 B.n49 163.367
R719 B.n254 B.n253 163.367
R720 B.n253 B.n252 163.367
R721 B.n252 B.n51 163.367
R722 B.n248 B.n51 163.367
R723 B.n248 B.n247 163.367
R724 B.n247 B.n246 163.367
R725 B.n246 B.n53 163.367
R726 B.n242 B.n53 163.367
R727 B.n242 B.n241 163.367
R728 B.n241 B.n240 163.367
R729 B.n240 B.n55 163.367
R730 B.n236 B.n55 163.367
R731 B.n236 B.n235 163.367
R732 B.n235 B.n234 163.367
R733 B.n234 B.n57 163.367
R734 B.n230 B.n57 163.367
R735 B.n230 B.n229 163.367
R736 B.n229 B.n228 163.367
R737 B.n228 B.n59 163.367
R738 B.n224 B.n59 163.367
R739 B.n224 B.n223 163.367
R740 B.n223 B.n222 163.367
R741 B.n222 B.n61 163.367
R742 B.n218 B.n61 163.367
R743 B.n218 B.n217 163.367
R744 B.n217 B.n216 163.367
R745 B.n216 B.n63 163.367
R746 B.n212 B.n63 163.367
R747 B.n212 B.n211 163.367
R748 B.n352 B.n13 163.367
R749 B.n352 B.n351 163.367
R750 B.n351 B.n350 163.367
R751 B.n350 B.n15 163.367
R752 B.n346 B.n15 163.367
R753 B.n346 B.n345 163.367
R754 B.n345 B.n344 163.367
R755 B.n344 B.n17 163.367
R756 B.n340 B.n17 163.367
R757 B.n340 B.n339 163.367
R758 B.n339 B.n338 163.367
R759 B.n338 B.n19 163.367
R760 B.n334 B.n19 163.367
R761 B.n334 B.n333 163.367
R762 B.n333 B.n332 163.367
R763 B.n332 B.n21 163.367
R764 B.n328 B.n21 163.367
R765 B.n328 B.n327 163.367
R766 B.n327 B.n326 163.367
R767 B.n326 B.n23 163.367
R768 B.n321 B.n23 163.367
R769 B.n321 B.n320 163.367
R770 B.n320 B.n319 163.367
R771 B.n319 B.n27 163.367
R772 B.n315 B.n27 163.367
R773 B.n315 B.n314 163.367
R774 B.n314 B.n313 163.367
R775 B.n313 B.n29 163.367
R776 B.n308 B.n29 163.367
R777 B.n308 B.n307 163.367
R778 B.n307 B.n306 163.367
R779 B.n306 B.n33 163.367
R780 B.n302 B.n33 163.367
R781 B.n302 B.n301 163.367
R782 B.n301 B.n300 163.367
R783 B.n300 B.n35 163.367
R784 B.n296 B.n35 163.367
R785 B.n296 B.n295 163.367
R786 B.n295 B.n294 163.367
R787 B.n294 B.n37 163.367
R788 B.n290 B.n37 163.367
R789 B.n290 B.n289 163.367
R790 B.n289 B.n288 163.367
R791 B.n288 B.n39 163.367
R792 B.n284 B.n39 163.367
R793 B.n284 B.n283 163.367
R794 B.n283 B.n282 163.367
R795 B.n282 B.n41 163.367
R796 B.n357 B.n356 163.367
R797 B.n358 B.n357 163.367
R798 B.n358 B.n11 163.367
R799 B.n362 B.n11 163.367
R800 B.n363 B.n362 163.367
R801 B.n364 B.n363 163.367
R802 B.n364 B.n9 163.367
R803 B.n368 B.n9 163.367
R804 B.n369 B.n368 163.367
R805 B.n370 B.n369 163.367
R806 B.n370 B.n7 163.367
R807 B.n374 B.n7 163.367
R808 B.n375 B.n374 163.367
R809 B.n376 B.n375 163.367
R810 B.n376 B.n5 163.367
R811 B.n380 B.n5 163.367
R812 B.n381 B.n380 163.367
R813 B.n382 B.n381 163.367
R814 B.n382 B.n3 163.367
R815 B.n386 B.n3 163.367
R816 B.n387 B.n386 163.367
R817 B.n101 B.n2 163.367
R818 B.n104 B.n101 163.367
R819 B.n105 B.n104 163.367
R820 B.n106 B.n105 163.367
R821 B.n106 B.n99 163.367
R822 B.n110 B.n99 163.367
R823 B.n111 B.n110 163.367
R824 B.n112 B.n111 163.367
R825 B.n112 B.n97 163.367
R826 B.n116 B.n97 163.367
R827 B.n117 B.n116 163.367
R828 B.n118 B.n117 163.367
R829 B.n118 B.n95 163.367
R830 B.n122 B.n95 163.367
R831 B.n123 B.n122 163.367
R832 B.n124 B.n123 163.367
R833 B.n124 B.n93 163.367
R834 B.n128 B.n93 163.367
R835 B.n129 B.n128 163.367
R836 B.n130 B.n129 163.367
R837 B.n130 B.n91 163.367
R838 B.n163 B.n81 59.5399
R839 B.n178 B.n177 59.5399
R840 B.n310 B.n31 59.5399
R841 B.n324 B.n25 59.5399
R842 B.n209 B.n64 35.7468
R843 B.n355 B.n354 35.7468
R844 B.n280 B.n279 35.7468
R845 B.n133 B.n132 35.7468
R846 B B.n389 18.0485
R847 B.n81 B.n80 16.0975
R848 B.n177 B.n176 16.0975
R849 B.n31 B.n30 16.0975
R850 B.n25 B.n24 16.0975
R851 B.n355 B.n12 10.6151
R852 B.n359 B.n12 10.6151
R853 B.n360 B.n359 10.6151
R854 B.n361 B.n360 10.6151
R855 B.n361 B.n10 10.6151
R856 B.n365 B.n10 10.6151
R857 B.n366 B.n365 10.6151
R858 B.n367 B.n366 10.6151
R859 B.n367 B.n8 10.6151
R860 B.n371 B.n8 10.6151
R861 B.n372 B.n371 10.6151
R862 B.n373 B.n372 10.6151
R863 B.n373 B.n6 10.6151
R864 B.n377 B.n6 10.6151
R865 B.n378 B.n377 10.6151
R866 B.n379 B.n378 10.6151
R867 B.n379 B.n4 10.6151
R868 B.n383 B.n4 10.6151
R869 B.n384 B.n383 10.6151
R870 B.n385 B.n384 10.6151
R871 B.n385 B.n0 10.6151
R872 B.n354 B.n353 10.6151
R873 B.n353 B.n14 10.6151
R874 B.n349 B.n14 10.6151
R875 B.n349 B.n348 10.6151
R876 B.n348 B.n347 10.6151
R877 B.n347 B.n16 10.6151
R878 B.n343 B.n16 10.6151
R879 B.n343 B.n342 10.6151
R880 B.n342 B.n341 10.6151
R881 B.n341 B.n18 10.6151
R882 B.n337 B.n18 10.6151
R883 B.n337 B.n336 10.6151
R884 B.n336 B.n335 10.6151
R885 B.n335 B.n20 10.6151
R886 B.n331 B.n20 10.6151
R887 B.n331 B.n330 10.6151
R888 B.n330 B.n329 10.6151
R889 B.n329 B.n22 10.6151
R890 B.n325 B.n22 10.6151
R891 B.n323 B.n322 10.6151
R892 B.n322 B.n26 10.6151
R893 B.n318 B.n26 10.6151
R894 B.n318 B.n317 10.6151
R895 B.n317 B.n316 10.6151
R896 B.n316 B.n28 10.6151
R897 B.n312 B.n28 10.6151
R898 B.n312 B.n311 10.6151
R899 B.n309 B.n32 10.6151
R900 B.n305 B.n32 10.6151
R901 B.n305 B.n304 10.6151
R902 B.n304 B.n303 10.6151
R903 B.n303 B.n34 10.6151
R904 B.n299 B.n34 10.6151
R905 B.n299 B.n298 10.6151
R906 B.n298 B.n297 10.6151
R907 B.n297 B.n36 10.6151
R908 B.n293 B.n36 10.6151
R909 B.n293 B.n292 10.6151
R910 B.n292 B.n291 10.6151
R911 B.n291 B.n38 10.6151
R912 B.n287 B.n38 10.6151
R913 B.n287 B.n286 10.6151
R914 B.n286 B.n285 10.6151
R915 B.n285 B.n40 10.6151
R916 B.n281 B.n40 10.6151
R917 B.n281 B.n280 10.6151
R918 B.n279 B.n42 10.6151
R919 B.n275 B.n42 10.6151
R920 B.n275 B.n274 10.6151
R921 B.n274 B.n273 10.6151
R922 B.n273 B.n44 10.6151
R923 B.n269 B.n44 10.6151
R924 B.n269 B.n268 10.6151
R925 B.n268 B.n267 10.6151
R926 B.n267 B.n46 10.6151
R927 B.n263 B.n46 10.6151
R928 B.n263 B.n262 10.6151
R929 B.n262 B.n261 10.6151
R930 B.n261 B.n48 10.6151
R931 B.n257 B.n48 10.6151
R932 B.n257 B.n256 10.6151
R933 B.n256 B.n255 10.6151
R934 B.n255 B.n50 10.6151
R935 B.n251 B.n50 10.6151
R936 B.n251 B.n250 10.6151
R937 B.n250 B.n249 10.6151
R938 B.n249 B.n52 10.6151
R939 B.n245 B.n52 10.6151
R940 B.n245 B.n244 10.6151
R941 B.n244 B.n243 10.6151
R942 B.n243 B.n54 10.6151
R943 B.n239 B.n54 10.6151
R944 B.n239 B.n238 10.6151
R945 B.n238 B.n237 10.6151
R946 B.n237 B.n56 10.6151
R947 B.n233 B.n56 10.6151
R948 B.n233 B.n232 10.6151
R949 B.n232 B.n231 10.6151
R950 B.n231 B.n58 10.6151
R951 B.n227 B.n58 10.6151
R952 B.n227 B.n226 10.6151
R953 B.n226 B.n225 10.6151
R954 B.n225 B.n60 10.6151
R955 B.n221 B.n60 10.6151
R956 B.n221 B.n220 10.6151
R957 B.n220 B.n219 10.6151
R958 B.n219 B.n62 10.6151
R959 B.n215 B.n62 10.6151
R960 B.n215 B.n214 10.6151
R961 B.n214 B.n213 10.6151
R962 B.n213 B.n64 10.6151
R963 B.n102 B.n1 10.6151
R964 B.n103 B.n102 10.6151
R965 B.n103 B.n100 10.6151
R966 B.n107 B.n100 10.6151
R967 B.n108 B.n107 10.6151
R968 B.n109 B.n108 10.6151
R969 B.n109 B.n98 10.6151
R970 B.n113 B.n98 10.6151
R971 B.n114 B.n113 10.6151
R972 B.n115 B.n114 10.6151
R973 B.n115 B.n96 10.6151
R974 B.n119 B.n96 10.6151
R975 B.n120 B.n119 10.6151
R976 B.n121 B.n120 10.6151
R977 B.n121 B.n94 10.6151
R978 B.n125 B.n94 10.6151
R979 B.n126 B.n125 10.6151
R980 B.n127 B.n126 10.6151
R981 B.n127 B.n92 10.6151
R982 B.n131 B.n92 10.6151
R983 B.n132 B.n131 10.6151
R984 B.n133 B.n90 10.6151
R985 B.n137 B.n90 10.6151
R986 B.n138 B.n137 10.6151
R987 B.n139 B.n138 10.6151
R988 B.n139 B.n88 10.6151
R989 B.n143 B.n88 10.6151
R990 B.n144 B.n143 10.6151
R991 B.n145 B.n144 10.6151
R992 B.n145 B.n86 10.6151
R993 B.n149 B.n86 10.6151
R994 B.n150 B.n149 10.6151
R995 B.n151 B.n150 10.6151
R996 B.n151 B.n84 10.6151
R997 B.n155 B.n84 10.6151
R998 B.n156 B.n155 10.6151
R999 B.n157 B.n156 10.6151
R1000 B.n157 B.n82 10.6151
R1001 B.n161 B.n82 10.6151
R1002 B.n162 B.n161 10.6151
R1003 B.n164 B.n78 10.6151
R1004 B.n168 B.n78 10.6151
R1005 B.n169 B.n168 10.6151
R1006 B.n170 B.n169 10.6151
R1007 B.n170 B.n76 10.6151
R1008 B.n174 B.n76 10.6151
R1009 B.n175 B.n174 10.6151
R1010 B.n179 B.n175 10.6151
R1011 B.n183 B.n74 10.6151
R1012 B.n184 B.n183 10.6151
R1013 B.n185 B.n184 10.6151
R1014 B.n185 B.n72 10.6151
R1015 B.n189 B.n72 10.6151
R1016 B.n190 B.n189 10.6151
R1017 B.n191 B.n190 10.6151
R1018 B.n191 B.n70 10.6151
R1019 B.n195 B.n70 10.6151
R1020 B.n196 B.n195 10.6151
R1021 B.n197 B.n196 10.6151
R1022 B.n197 B.n68 10.6151
R1023 B.n201 B.n68 10.6151
R1024 B.n202 B.n201 10.6151
R1025 B.n203 B.n202 10.6151
R1026 B.n203 B.n66 10.6151
R1027 B.n207 B.n66 10.6151
R1028 B.n208 B.n207 10.6151
R1029 B.n209 B.n208 10.6151
R1030 B.n389 B.n0 8.11757
R1031 B.n389 B.n1 8.11757
R1032 B.n324 B.n323 6.5566
R1033 B.n311 B.n310 6.5566
R1034 B.n164 B.n163 6.5566
R1035 B.n179 B.n178 6.5566
R1036 B.n325 B.n324 4.05904
R1037 B.n310 B.n309 4.05904
R1038 B.n163 B.n162 4.05904
R1039 B.n178 B.n74 4.05904
C0 VDD2 VTAIL 7.7585f
C1 w_n1966_n1882# VN 3.42251f
C2 VDD1 VN 0.152548f
C3 VP B 1.07278f
C4 VDD2 w_n1966_n1882# 1.43024f
C5 VDD2 VDD1 0.845709f
C6 VDD2 VN 2.35961f
C7 VP VTAIL 2.46411f
C8 w_n1966_n1882# VP 3.67184f
C9 VTAIL B 1.31408f
C10 VDD1 VP 2.52383f
C11 VP VN 3.93238f
C12 w_n1966_n1882# B 4.93526f
C13 VDD1 B 1.08302f
C14 VDD2 VP 0.319248f
C15 VN B 0.664938f
C16 VDD2 B 1.11968f
C17 w_n1966_n1882# VTAIL 1.836f
C18 VDD1 VTAIL 7.72187f
C19 VN VTAIL 2.44978f
C20 w_n1966_n1882# VDD1 1.39613f
C21 VDD2 VSUBS 1.043014f
C22 VDD1 VSUBS 0.840236f
C23 VTAIL VSUBS 0.365167f
C24 VN VSUBS 4.12766f
C25 VP VSUBS 1.190292f
C26 B VSUBS 2.034056f
C27 w_n1966_n1882# VSUBS 46.452602f
C28 B.n0 VSUBS 0.00625f
C29 B.n1 VSUBS 0.00625f
C30 B.n2 VSUBS 0.009243f
C31 B.n3 VSUBS 0.007083f
C32 B.n4 VSUBS 0.007083f
C33 B.n5 VSUBS 0.007083f
C34 B.n6 VSUBS 0.007083f
C35 B.n7 VSUBS 0.007083f
C36 B.n8 VSUBS 0.007083f
C37 B.n9 VSUBS 0.007083f
C38 B.n10 VSUBS 0.007083f
C39 B.n11 VSUBS 0.007083f
C40 B.n12 VSUBS 0.007083f
C41 B.n13 VSUBS 0.018098f
C42 B.n14 VSUBS 0.007083f
C43 B.n15 VSUBS 0.007083f
C44 B.n16 VSUBS 0.007083f
C45 B.n17 VSUBS 0.007083f
C46 B.n18 VSUBS 0.007083f
C47 B.n19 VSUBS 0.007083f
C48 B.n20 VSUBS 0.007083f
C49 B.n21 VSUBS 0.007083f
C50 B.n22 VSUBS 0.007083f
C51 B.n23 VSUBS 0.007083f
C52 B.t1 VSUBS 0.066783f
C53 B.t2 VSUBS 0.07365f
C54 B.t0 VSUBS 0.099711f
C55 B.n24 VSUBS 0.132867f
C56 B.n25 VSUBS 0.120951f
C57 B.n26 VSUBS 0.007083f
C58 B.n27 VSUBS 0.007083f
C59 B.n28 VSUBS 0.007083f
C60 B.n29 VSUBS 0.007083f
C61 B.t4 VSUBS 0.066785f
C62 B.t5 VSUBS 0.073651f
C63 B.t3 VSUBS 0.099711f
C64 B.n30 VSUBS 0.132866f
C65 B.n31 VSUBS 0.12095f
C66 B.n32 VSUBS 0.007083f
C67 B.n33 VSUBS 0.007083f
C68 B.n34 VSUBS 0.007083f
C69 B.n35 VSUBS 0.007083f
C70 B.n36 VSUBS 0.007083f
C71 B.n37 VSUBS 0.007083f
C72 B.n38 VSUBS 0.007083f
C73 B.n39 VSUBS 0.007083f
C74 B.n40 VSUBS 0.007083f
C75 B.n41 VSUBS 0.018098f
C76 B.n42 VSUBS 0.007083f
C77 B.n43 VSUBS 0.007083f
C78 B.n44 VSUBS 0.007083f
C79 B.n45 VSUBS 0.007083f
C80 B.n46 VSUBS 0.007083f
C81 B.n47 VSUBS 0.007083f
C82 B.n48 VSUBS 0.007083f
C83 B.n49 VSUBS 0.007083f
C84 B.n50 VSUBS 0.007083f
C85 B.n51 VSUBS 0.007083f
C86 B.n52 VSUBS 0.007083f
C87 B.n53 VSUBS 0.007083f
C88 B.n54 VSUBS 0.007083f
C89 B.n55 VSUBS 0.007083f
C90 B.n56 VSUBS 0.007083f
C91 B.n57 VSUBS 0.007083f
C92 B.n58 VSUBS 0.007083f
C93 B.n59 VSUBS 0.007083f
C94 B.n60 VSUBS 0.007083f
C95 B.n61 VSUBS 0.007083f
C96 B.n62 VSUBS 0.007083f
C97 B.n63 VSUBS 0.007083f
C98 B.n64 VSUBS 0.017874f
C99 B.n65 VSUBS 0.007083f
C100 B.n66 VSUBS 0.007083f
C101 B.n67 VSUBS 0.007083f
C102 B.n68 VSUBS 0.007083f
C103 B.n69 VSUBS 0.007083f
C104 B.n70 VSUBS 0.007083f
C105 B.n71 VSUBS 0.007083f
C106 B.n72 VSUBS 0.007083f
C107 B.n73 VSUBS 0.007083f
C108 B.n74 VSUBS 0.004896f
C109 B.n75 VSUBS 0.007083f
C110 B.n76 VSUBS 0.007083f
C111 B.n77 VSUBS 0.007083f
C112 B.n78 VSUBS 0.007083f
C113 B.n79 VSUBS 0.007083f
C114 B.t8 VSUBS 0.066783f
C115 B.t7 VSUBS 0.07365f
C116 B.t6 VSUBS 0.099711f
C117 B.n80 VSUBS 0.132867f
C118 B.n81 VSUBS 0.120951f
C119 B.n82 VSUBS 0.007083f
C120 B.n83 VSUBS 0.007083f
C121 B.n84 VSUBS 0.007083f
C122 B.n85 VSUBS 0.007083f
C123 B.n86 VSUBS 0.007083f
C124 B.n87 VSUBS 0.007083f
C125 B.n88 VSUBS 0.007083f
C126 B.n89 VSUBS 0.007083f
C127 B.n90 VSUBS 0.007083f
C128 B.n91 VSUBS 0.01711f
C129 B.n92 VSUBS 0.007083f
C130 B.n93 VSUBS 0.007083f
C131 B.n94 VSUBS 0.007083f
C132 B.n95 VSUBS 0.007083f
C133 B.n96 VSUBS 0.007083f
C134 B.n97 VSUBS 0.007083f
C135 B.n98 VSUBS 0.007083f
C136 B.n99 VSUBS 0.007083f
C137 B.n100 VSUBS 0.007083f
C138 B.n101 VSUBS 0.007083f
C139 B.n102 VSUBS 0.007083f
C140 B.n103 VSUBS 0.007083f
C141 B.n104 VSUBS 0.007083f
C142 B.n105 VSUBS 0.007083f
C143 B.n106 VSUBS 0.007083f
C144 B.n107 VSUBS 0.007083f
C145 B.n108 VSUBS 0.007083f
C146 B.n109 VSUBS 0.007083f
C147 B.n110 VSUBS 0.007083f
C148 B.n111 VSUBS 0.007083f
C149 B.n112 VSUBS 0.007083f
C150 B.n113 VSUBS 0.007083f
C151 B.n114 VSUBS 0.007083f
C152 B.n115 VSUBS 0.007083f
C153 B.n116 VSUBS 0.007083f
C154 B.n117 VSUBS 0.007083f
C155 B.n118 VSUBS 0.007083f
C156 B.n119 VSUBS 0.007083f
C157 B.n120 VSUBS 0.007083f
C158 B.n121 VSUBS 0.007083f
C159 B.n122 VSUBS 0.007083f
C160 B.n123 VSUBS 0.007083f
C161 B.n124 VSUBS 0.007083f
C162 B.n125 VSUBS 0.007083f
C163 B.n126 VSUBS 0.007083f
C164 B.n127 VSUBS 0.007083f
C165 B.n128 VSUBS 0.007083f
C166 B.n129 VSUBS 0.007083f
C167 B.n130 VSUBS 0.007083f
C168 B.n131 VSUBS 0.007083f
C169 B.n132 VSUBS 0.01711f
C170 B.n133 VSUBS 0.018098f
C171 B.n134 VSUBS 0.018098f
C172 B.n135 VSUBS 0.007083f
C173 B.n136 VSUBS 0.007083f
C174 B.n137 VSUBS 0.007083f
C175 B.n138 VSUBS 0.007083f
C176 B.n139 VSUBS 0.007083f
C177 B.n140 VSUBS 0.007083f
C178 B.n141 VSUBS 0.007083f
C179 B.n142 VSUBS 0.007083f
C180 B.n143 VSUBS 0.007083f
C181 B.n144 VSUBS 0.007083f
C182 B.n145 VSUBS 0.007083f
C183 B.n146 VSUBS 0.007083f
C184 B.n147 VSUBS 0.007083f
C185 B.n148 VSUBS 0.007083f
C186 B.n149 VSUBS 0.007083f
C187 B.n150 VSUBS 0.007083f
C188 B.n151 VSUBS 0.007083f
C189 B.n152 VSUBS 0.007083f
C190 B.n153 VSUBS 0.007083f
C191 B.n154 VSUBS 0.007083f
C192 B.n155 VSUBS 0.007083f
C193 B.n156 VSUBS 0.007083f
C194 B.n157 VSUBS 0.007083f
C195 B.n158 VSUBS 0.007083f
C196 B.n159 VSUBS 0.007083f
C197 B.n160 VSUBS 0.007083f
C198 B.n161 VSUBS 0.007083f
C199 B.n162 VSUBS 0.004896f
C200 B.n163 VSUBS 0.016411f
C201 B.n164 VSUBS 0.005729f
C202 B.n165 VSUBS 0.007083f
C203 B.n166 VSUBS 0.007083f
C204 B.n167 VSUBS 0.007083f
C205 B.n168 VSUBS 0.007083f
C206 B.n169 VSUBS 0.007083f
C207 B.n170 VSUBS 0.007083f
C208 B.n171 VSUBS 0.007083f
C209 B.n172 VSUBS 0.007083f
C210 B.n173 VSUBS 0.007083f
C211 B.n174 VSUBS 0.007083f
C212 B.n175 VSUBS 0.007083f
C213 B.t11 VSUBS 0.066785f
C214 B.t10 VSUBS 0.073651f
C215 B.t9 VSUBS 0.099711f
C216 B.n176 VSUBS 0.132866f
C217 B.n177 VSUBS 0.12095f
C218 B.n178 VSUBS 0.016411f
C219 B.n179 VSUBS 0.005729f
C220 B.n180 VSUBS 0.007083f
C221 B.n181 VSUBS 0.007083f
C222 B.n182 VSUBS 0.007083f
C223 B.n183 VSUBS 0.007083f
C224 B.n184 VSUBS 0.007083f
C225 B.n185 VSUBS 0.007083f
C226 B.n186 VSUBS 0.007083f
C227 B.n187 VSUBS 0.007083f
C228 B.n188 VSUBS 0.007083f
C229 B.n189 VSUBS 0.007083f
C230 B.n190 VSUBS 0.007083f
C231 B.n191 VSUBS 0.007083f
C232 B.n192 VSUBS 0.007083f
C233 B.n193 VSUBS 0.007083f
C234 B.n194 VSUBS 0.007083f
C235 B.n195 VSUBS 0.007083f
C236 B.n196 VSUBS 0.007083f
C237 B.n197 VSUBS 0.007083f
C238 B.n198 VSUBS 0.007083f
C239 B.n199 VSUBS 0.007083f
C240 B.n200 VSUBS 0.007083f
C241 B.n201 VSUBS 0.007083f
C242 B.n202 VSUBS 0.007083f
C243 B.n203 VSUBS 0.007083f
C244 B.n204 VSUBS 0.007083f
C245 B.n205 VSUBS 0.007083f
C246 B.n206 VSUBS 0.007083f
C247 B.n207 VSUBS 0.007083f
C248 B.n208 VSUBS 0.007083f
C249 B.n209 VSUBS 0.017334f
C250 B.n210 VSUBS 0.018098f
C251 B.n211 VSUBS 0.01711f
C252 B.n212 VSUBS 0.007083f
C253 B.n213 VSUBS 0.007083f
C254 B.n214 VSUBS 0.007083f
C255 B.n215 VSUBS 0.007083f
C256 B.n216 VSUBS 0.007083f
C257 B.n217 VSUBS 0.007083f
C258 B.n218 VSUBS 0.007083f
C259 B.n219 VSUBS 0.007083f
C260 B.n220 VSUBS 0.007083f
C261 B.n221 VSUBS 0.007083f
C262 B.n222 VSUBS 0.007083f
C263 B.n223 VSUBS 0.007083f
C264 B.n224 VSUBS 0.007083f
C265 B.n225 VSUBS 0.007083f
C266 B.n226 VSUBS 0.007083f
C267 B.n227 VSUBS 0.007083f
C268 B.n228 VSUBS 0.007083f
C269 B.n229 VSUBS 0.007083f
C270 B.n230 VSUBS 0.007083f
C271 B.n231 VSUBS 0.007083f
C272 B.n232 VSUBS 0.007083f
C273 B.n233 VSUBS 0.007083f
C274 B.n234 VSUBS 0.007083f
C275 B.n235 VSUBS 0.007083f
C276 B.n236 VSUBS 0.007083f
C277 B.n237 VSUBS 0.007083f
C278 B.n238 VSUBS 0.007083f
C279 B.n239 VSUBS 0.007083f
C280 B.n240 VSUBS 0.007083f
C281 B.n241 VSUBS 0.007083f
C282 B.n242 VSUBS 0.007083f
C283 B.n243 VSUBS 0.007083f
C284 B.n244 VSUBS 0.007083f
C285 B.n245 VSUBS 0.007083f
C286 B.n246 VSUBS 0.007083f
C287 B.n247 VSUBS 0.007083f
C288 B.n248 VSUBS 0.007083f
C289 B.n249 VSUBS 0.007083f
C290 B.n250 VSUBS 0.007083f
C291 B.n251 VSUBS 0.007083f
C292 B.n252 VSUBS 0.007083f
C293 B.n253 VSUBS 0.007083f
C294 B.n254 VSUBS 0.007083f
C295 B.n255 VSUBS 0.007083f
C296 B.n256 VSUBS 0.007083f
C297 B.n257 VSUBS 0.007083f
C298 B.n258 VSUBS 0.007083f
C299 B.n259 VSUBS 0.007083f
C300 B.n260 VSUBS 0.007083f
C301 B.n261 VSUBS 0.007083f
C302 B.n262 VSUBS 0.007083f
C303 B.n263 VSUBS 0.007083f
C304 B.n264 VSUBS 0.007083f
C305 B.n265 VSUBS 0.007083f
C306 B.n266 VSUBS 0.007083f
C307 B.n267 VSUBS 0.007083f
C308 B.n268 VSUBS 0.007083f
C309 B.n269 VSUBS 0.007083f
C310 B.n270 VSUBS 0.007083f
C311 B.n271 VSUBS 0.007083f
C312 B.n272 VSUBS 0.007083f
C313 B.n273 VSUBS 0.007083f
C314 B.n274 VSUBS 0.007083f
C315 B.n275 VSUBS 0.007083f
C316 B.n276 VSUBS 0.007083f
C317 B.n277 VSUBS 0.007083f
C318 B.n278 VSUBS 0.01711f
C319 B.n279 VSUBS 0.01711f
C320 B.n280 VSUBS 0.018098f
C321 B.n281 VSUBS 0.007083f
C322 B.n282 VSUBS 0.007083f
C323 B.n283 VSUBS 0.007083f
C324 B.n284 VSUBS 0.007083f
C325 B.n285 VSUBS 0.007083f
C326 B.n286 VSUBS 0.007083f
C327 B.n287 VSUBS 0.007083f
C328 B.n288 VSUBS 0.007083f
C329 B.n289 VSUBS 0.007083f
C330 B.n290 VSUBS 0.007083f
C331 B.n291 VSUBS 0.007083f
C332 B.n292 VSUBS 0.007083f
C333 B.n293 VSUBS 0.007083f
C334 B.n294 VSUBS 0.007083f
C335 B.n295 VSUBS 0.007083f
C336 B.n296 VSUBS 0.007083f
C337 B.n297 VSUBS 0.007083f
C338 B.n298 VSUBS 0.007083f
C339 B.n299 VSUBS 0.007083f
C340 B.n300 VSUBS 0.007083f
C341 B.n301 VSUBS 0.007083f
C342 B.n302 VSUBS 0.007083f
C343 B.n303 VSUBS 0.007083f
C344 B.n304 VSUBS 0.007083f
C345 B.n305 VSUBS 0.007083f
C346 B.n306 VSUBS 0.007083f
C347 B.n307 VSUBS 0.007083f
C348 B.n308 VSUBS 0.007083f
C349 B.n309 VSUBS 0.004896f
C350 B.n310 VSUBS 0.016411f
C351 B.n311 VSUBS 0.005729f
C352 B.n312 VSUBS 0.007083f
C353 B.n313 VSUBS 0.007083f
C354 B.n314 VSUBS 0.007083f
C355 B.n315 VSUBS 0.007083f
C356 B.n316 VSUBS 0.007083f
C357 B.n317 VSUBS 0.007083f
C358 B.n318 VSUBS 0.007083f
C359 B.n319 VSUBS 0.007083f
C360 B.n320 VSUBS 0.007083f
C361 B.n321 VSUBS 0.007083f
C362 B.n322 VSUBS 0.007083f
C363 B.n323 VSUBS 0.005729f
C364 B.n324 VSUBS 0.016411f
C365 B.n325 VSUBS 0.004896f
C366 B.n326 VSUBS 0.007083f
C367 B.n327 VSUBS 0.007083f
C368 B.n328 VSUBS 0.007083f
C369 B.n329 VSUBS 0.007083f
C370 B.n330 VSUBS 0.007083f
C371 B.n331 VSUBS 0.007083f
C372 B.n332 VSUBS 0.007083f
C373 B.n333 VSUBS 0.007083f
C374 B.n334 VSUBS 0.007083f
C375 B.n335 VSUBS 0.007083f
C376 B.n336 VSUBS 0.007083f
C377 B.n337 VSUBS 0.007083f
C378 B.n338 VSUBS 0.007083f
C379 B.n339 VSUBS 0.007083f
C380 B.n340 VSUBS 0.007083f
C381 B.n341 VSUBS 0.007083f
C382 B.n342 VSUBS 0.007083f
C383 B.n343 VSUBS 0.007083f
C384 B.n344 VSUBS 0.007083f
C385 B.n345 VSUBS 0.007083f
C386 B.n346 VSUBS 0.007083f
C387 B.n347 VSUBS 0.007083f
C388 B.n348 VSUBS 0.007083f
C389 B.n349 VSUBS 0.007083f
C390 B.n350 VSUBS 0.007083f
C391 B.n351 VSUBS 0.007083f
C392 B.n352 VSUBS 0.007083f
C393 B.n353 VSUBS 0.007083f
C394 B.n354 VSUBS 0.018098f
C395 B.n355 VSUBS 0.01711f
C396 B.n356 VSUBS 0.01711f
C397 B.n357 VSUBS 0.007083f
C398 B.n358 VSUBS 0.007083f
C399 B.n359 VSUBS 0.007083f
C400 B.n360 VSUBS 0.007083f
C401 B.n361 VSUBS 0.007083f
C402 B.n362 VSUBS 0.007083f
C403 B.n363 VSUBS 0.007083f
C404 B.n364 VSUBS 0.007083f
C405 B.n365 VSUBS 0.007083f
C406 B.n366 VSUBS 0.007083f
C407 B.n367 VSUBS 0.007083f
C408 B.n368 VSUBS 0.007083f
C409 B.n369 VSUBS 0.007083f
C410 B.n370 VSUBS 0.007083f
C411 B.n371 VSUBS 0.007083f
C412 B.n372 VSUBS 0.007083f
C413 B.n373 VSUBS 0.007083f
C414 B.n374 VSUBS 0.007083f
C415 B.n375 VSUBS 0.007083f
C416 B.n376 VSUBS 0.007083f
C417 B.n377 VSUBS 0.007083f
C418 B.n378 VSUBS 0.007083f
C419 B.n379 VSUBS 0.007083f
C420 B.n380 VSUBS 0.007083f
C421 B.n381 VSUBS 0.007083f
C422 B.n382 VSUBS 0.007083f
C423 B.n383 VSUBS 0.007083f
C424 B.n384 VSUBS 0.007083f
C425 B.n385 VSUBS 0.007083f
C426 B.n386 VSUBS 0.007083f
C427 B.n387 VSUBS 0.009243f
C428 B.n388 VSUBS 0.009846f
C429 B.n389 VSUBS 0.019581f
C430 VDD2.n0 VSUBS 0.027905f
C431 VDD2.n1 VSUBS 0.026204f
C432 VDD2.n2 VSUBS 0.014081f
C433 VDD2.n3 VSUBS 0.033282f
C434 VDD2.n4 VSUBS 0.014909f
C435 VDD2.n5 VSUBS 0.429344f
C436 VDD2.n6 VSUBS 0.014081f
C437 VDD2.t5 VSUBS 0.072312f
C438 VDD2.n7 VSUBS 0.105534f
C439 VDD2.n8 VSUBS 0.021084f
C440 VDD2.n9 VSUBS 0.024961f
C441 VDD2.n10 VSUBS 0.033282f
C442 VDD2.n11 VSUBS 0.014909f
C443 VDD2.n12 VSUBS 0.014081f
C444 VDD2.n13 VSUBS 0.026204f
C445 VDD2.n14 VSUBS 0.026204f
C446 VDD2.n15 VSUBS 0.014081f
C447 VDD2.n16 VSUBS 0.014909f
C448 VDD2.n17 VSUBS 0.033282f
C449 VDD2.n18 VSUBS 0.07755f
C450 VDD2.n19 VSUBS 0.014909f
C451 VDD2.n20 VSUBS 0.014081f
C452 VDD2.n21 VSUBS 0.060926f
C453 VDD2.n22 VSUBS 0.058563f
C454 VDD2.t6 VSUBS 0.094631f
C455 VDD2.t0 VSUBS 0.094631f
C456 VDD2.n23 VSUBS 0.577975f
C457 VDD2.n24 VSUBS 0.574368f
C458 VDD2.t1 VSUBS 0.094631f
C459 VDD2.t3 VSUBS 0.094631f
C460 VDD2.n25 VSUBS 0.580282f
C461 VDD2.n26 VSUBS 1.59692f
C462 VDD2.n27 VSUBS 0.027905f
C463 VDD2.n28 VSUBS 0.026204f
C464 VDD2.n29 VSUBS 0.014081f
C465 VDD2.n30 VSUBS 0.033282f
C466 VDD2.n31 VSUBS 0.014909f
C467 VDD2.n32 VSUBS 0.429344f
C468 VDD2.n33 VSUBS 0.014081f
C469 VDD2.t9 VSUBS 0.072312f
C470 VDD2.n34 VSUBS 0.105534f
C471 VDD2.n35 VSUBS 0.021084f
C472 VDD2.n36 VSUBS 0.024961f
C473 VDD2.n37 VSUBS 0.033282f
C474 VDD2.n38 VSUBS 0.014909f
C475 VDD2.n39 VSUBS 0.014081f
C476 VDD2.n40 VSUBS 0.026204f
C477 VDD2.n41 VSUBS 0.026204f
C478 VDD2.n42 VSUBS 0.014081f
C479 VDD2.n43 VSUBS 0.014909f
C480 VDD2.n44 VSUBS 0.033282f
C481 VDD2.n45 VSUBS 0.07755f
C482 VDD2.n46 VSUBS 0.014909f
C483 VDD2.n47 VSUBS 0.014081f
C484 VDD2.n48 VSUBS 0.060926f
C485 VDD2.n49 VSUBS 0.056966f
C486 VDD2.n50 VSUBS 1.55524f
C487 VDD2.t4 VSUBS 0.094631f
C488 VDD2.t8 VSUBS 0.094631f
C489 VDD2.n51 VSUBS 0.577978f
C490 VDD2.n52 VSUBS 0.469555f
C491 VDD2.t2 VSUBS 0.094631f
C492 VDD2.t7 VSUBS 0.094631f
C493 VDD2.n53 VSUBS 0.580261f
C494 VN.n0 VSUBS 0.066967f
C495 VN.t9 VSUBS 0.448852f
C496 VN.n1 VSUBS 0.237101f
C497 VN.t4 VSUBS 0.46393f
C498 VN.n2 VSUBS 0.215494f
C499 VN.t3 VSUBS 0.448852f
C500 VN.n3 VSUBS 0.233385f
C501 VN.n4 VSUBS 0.015196f
C502 VN.n5 VSUBS 0.213624f
C503 VN.n6 VSUBS 0.066967f
C504 VN.n7 VSUBS 0.066967f
C505 VN.n8 VSUBS 0.015196f
C506 VN.t8 VSUBS 0.448852f
C507 VN.n9 VSUBS 0.233385f
C508 VN.t6 VSUBS 0.448852f
C509 VN.n10 VSUBS 0.230082f
C510 VN.n11 VSUBS 0.051897f
C511 VN.n12 VSUBS 0.066967f
C512 VN.t1 VSUBS 0.448852f
C513 VN.n13 VSUBS 0.237101f
C514 VN.t2 VSUBS 0.46393f
C515 VN.n14 VSUBS 0.215494f
C516 VN.t7 VSUBS 0.448852f
C517 VN.n15 VSUBS 0.233385f
C518 VN.n16 VSUBS 0.015196f
C519 VN.n17 VSUBS 0.213624f
C520 VN.n18 VSUBS 0.066967f
C521 VN.n19 VSUBS 0.066967f
C522 VN.n20 VSUBS 0.015196f
C523 VN.t5 VSUBS 0.448852f
C524 VN.n21 VSUBS 0.233385f
C525 VN.t0 VSUBS 0.448852f
C526 VN.n22 VSUBS 0.230082f
C527 VN.n23 VSUBS 2.16029f
C528 VDD1.n0 VSUBS 0.027643f
C529 VDD1.n1 VSUBS 0.025957f
C530 VDD1.n2 VSUBS 0.013948f
C531 VDD1.n3 VSUBS 0.032969f
C532 VDD1.n4 VSUBS 0.014769f
C533 VDD1.n5 VSUBS 0.425309f
C534 VDD1.n6 VSUBS 0.013948f
C535 VDD1.t9 VSUBS 0.071632f
C536 VDD1.n7 VSUBS 0.104542f
C537 VDD1.n8 VSUBS 0.020886f
C538 VDD1.n9 VSUBS 0.024727f
C539 VDD1.n10 VSUBS 0.032969f
C540 VDD1.n11 VSUBS 0.014769f
C541 VDD1.n12 VSUBS 0.013948f
C542 VDD1.n13 VSUBS 0.025957f
C543 VDD1.n14 VSUBS 0.025957f
C544 VDD1.n15 VSUBS 0.013948f
C545 VDD1.n16 VSUBS 0.014769f
C546 VDD1.n17 VSUBS 0.032969f
C547 VDD1.n18 VSUBS 0.076821f
C548 VDD1.n19 VSUBS 0.014769f
C549 VDD1.n20 VSUBS 0.013948f
C550 VDD1.n21 VSUBS 0.060354f
C551 VDD1.n22 VSUBS 0.058012f
C552 VDD1.t4 VSUBS 0.093741f
C553 VDD1.t1 VSUBS 0.093741f
C554 VDD1.n23 VSUBS 0.572546f
C555 VDD1.n24 VSUBS 0.573591f
C556 VDD1.n25 VSUBS 0.027643f
C557 VDD1.n26 VSUBS 0.025957f
C558 VDD1.n27 VSUBS 0.013948f
C559 VDD1.n28 VSUBS 0.032969f
C560 VDD1.n29 VSUBS 0.014769f
C561 VDD1.n30 VSUBS 0.425309f
C562 VDD1.n31 VSUBS 0.013948f
C563 VDD1.t5 VSUBS 0.071632f
C564 VDD1.n32 VSUBS 0.104542f
C565 VDD1.n33 VSUBS 0.020886f
C566 VDD1.n34 VSUBS 0.024727f
C567 VDD1.n35 VSUBS 0.032969f
C568 VDD1.n36 VSUBS 0.014769f
C569 VDD1.n37 VSUBS 0.013948f
C570 VDD1.n38 VSUBS 0.025957f
C571 VDD1.n39 VSUBS 0.025957f
C572 VDD1.n40 VSUBS 0.013948f
C573 VDD1.n41 VSUBS 0.014769f
C574 VDD1.n42 VSUBS 0.032969f
C575 VDD1.n43 VSUBS 0.076821f
C576 VDD1.n44 VSUBS 0.014769f
C577 VDD1.n45 VSUBS 0.013948f
C578 VDD1.n46 VSUBS 0.060354f
C579 VDD1.n47 VSUBS 0.058012f
C580 VDD1.t3 VSUBS 0.093741f
C581 VDD1.t0 VSUBS 0.093741f
C582 VDD1.n48 VSUBS 0.572543f
C583 VDD1.n49 VSUBS 0.568969f
C584 VDD1.t6 VSUBS 0.093741f
C585 VDD1.t7 VSUBS 0.093741f
C586 VDD1.n50 VSUBS 0.574827f
C587 VDD1.n51 VSUBS 1.65427f
C588 VDD1.t8 VSUBS 0.093741f
C589 VDD1.t2 VSUBS 0.093741f
C590 VDD1.n52 VSUBS 0.572543f
C591 VDD1.n53 VSUBS 1.94989f
C592 VTAIL.t5 VSUBS 0.106731f
C593 VTAIL.t3 VSUBS 0.106731f
C594 VTAIL.n0 VSUBS 0.569384f
C595 VTAIL.n1 VSUBS 0.616667f
C596 VTAIL.n2 VSUBS 0.031473f
C597 VTAIL.n3 VSUBS 0.029554f
C598 VTAIL.n4 VSUBS 0.015881f
C599 VTAIL.n5 VSUBS 0.037537f
C600 VTAIL.n6 VSUBS 0.016815f
C601 VTAIL.n7 VSUBS 0.484243f
C602 VTAIL.n8 VSUBS 0.015881f
C603 VTAIL.t13 VSUBS 0.081558f
C604 VTAIL.n9 VSUBS 0.119028f
C605 VTAIL.n10 VSUBS 0.02378f
C606 VTAIL.n11 VSUBS 0.028153f
C607 VTAIL.n12 VSUBS 0.037537f
C608 VTAIL.n13 VSUBS 0.016815f
C609 VTAIL.n14 VSUBS 0.015881f
C610 VTAIL.n15 VSUBS 0.029554f
C611 VTAIL.n16 VSUBS 0.029554f
C612 VTAIL.n17 VSUBS 0.015881f
C613 VTAIL.n18 VSUBS 0.016815f
C614 VTAIL.n19 VSUBS 0.037537f
C615 VTAIL.n20 VSUBS 0.087466f
C616 VTAIL.n21 VSUBS 0.016815f
C617 VTAIL.n22 VSUBS 0.015881f
C618 VTAIL.n23 VSUBS 0.068717f
C619 VTAIL.n24 VSUBS 0.043847f
C620 VTAIL.n25 VSUBS 0.17242f
C621 VTAIL.t11 VSUBS 0.106731f
C622 VTAIL.t18 VSUBS 0.106731f
C623 VTAIL.n26 VSUBS 0.569384f
C624 VTAIL.n27 VSUBS 0.617488f
C625 VTAIL.t16 VSUBS 0.106731f
C626 VTAIL.t17 VSUBS 0.106731f
C627 VTAIL.n28 VSUBS 0.569384f
C628 VTAIL.n29 VSUBS 1.46226f
C629 VTAIL.t7 VSUBS 0.106731f
C630 VTAIL.t6 VSUBS 0.106731f
C631 VTAIL.n30 VSUBS 0.569388f
C632 VTAIL.n31 VSUBS 1.46226f
C633 VTAIL.t9 VSUBS 0.106731f
C634 VTAIL.t1 VSUBS 0.106731f
C635 VTAIL.n32 VSUBS 0.569388f
C636 VTAIL.n33 VSUBS 0.617484f
C637 VTAIL.n34 VSUBS 0.031473f
C638 VTAIL.n35 VSUBS 0.029554f
C639 VTAIL.n36 VSUBS 0.015881f
C640 VTAIL.n37 VSUBS 0.037537f
C641 VTAIL.n38 VSUBS 0.016815f
C642 VTAIL.n39 VSUBS 0.484243f
C643 VTAIL.n40 VSUBS 0.015881f
C644 VTAIL.t8 VSUBS 0.081558f
C645 VTAIL.n41 VSUBS 0.119028f
C646 VTAIL.n42 VSUBS 0.02378f
C647 VTAIL.n43 VSUBS 0.028153f
C648 VTAIL.n44 VSUBS 0.037537f
C649 VTAIL.n45 VSUBS 0.016815f
C650 VTAIL.n46 VSUBS 0.015881f
C651 VTAIL.n47 VSUBS 0.029554f
C652 VTAIL.n48 VSUBS 0.029554f
C653 VTAIL.n49 VSUBS 0.015881f
C654 VTAIL.n50 VSUBS 0.016815f
C655 VTAIL.n51 VSUBS 0.037537f
C656 VTAIL.n52 VSUBS 0.087466f
C657 VTAIL.n53 VSUBS 0.016815f
C658 VTAIL.n54 VSUBS 0.015881f
C659 VTAIL.n55 VSUBS 0.068717f
C660 VTAIL.n56 VSUBS 0.043847f
C661 VTAIL.n57 VSUBS 0.17242f
C662 VTAIL.t15 VSUBS 0.106731f
C663 VTAIL.t19 VSUBS 0.106731f
C664 VTAIL.n58 VSUBS 0.569388f
C665 VTAIL.n59 VSUBS 0.628156f
C666 VTAIL.t14 VSUBS 0.106731f
C667 VTAIL.t10 VSUBS 0.106731f
C668 VTAIL.n60 VSUBS 0.569388f
C669 VTAIL.n61 VSUBS 0.617484f
C670 VTAIL.n62 VSUBS 0.031473f
C671 VTAIL.n63 VSUBS 0.029554f
C672 VTAIL.n64 VSUBS 0.015881f
C673 VTAIL.n65 VSUBS 0.037537f
C674 VTAIL.n66 VSUBS 0.016815f
C675 VTAIL.n67 VSUBS 0.484243f
C676 VTAIL.n68 VSUBS 0.015881f
C677 VTAIL.t12 VSUBS 0.081558f
C678 VTAIL.n69 VSUBS 0.119028f
C679 VTAIL.n70 VSUBS 0.02378f
C680 VTAIL.n71 VSUBS 0.028153f
C681 VTAIL.n72 VSUBS 0.037537f
C682 VTAIL.n73 VSUBS 0.016815f
C683 VTAIL.n74 VSUBS 0.015881f
C684 VTAIL.n75 VSUBS 0.029554f
C685 VTAIL.n76 VSUBS 0.029554f
C686 VTAIL.n77 VSUBS 0.015881f
C687 VTAIL.n78 VSUBS 0.016815f
C688 VTAIL.n79 VSUBS 0.037537f
C689 VTAIL.n80 VSUBS 0.087466f
C690 VTAIL.n81 VSUBS 0.016815f
C691 VTAIL.n82 VSUBS 0.015881f
C692 VTAIL.n83 VSUBS 0.068717f
C693 VTAIL.n84 VSUBS 0.043847f
C694 VTAIL.n85 VSUBS 0.938383f
C695 VTAIL.n86 VSUBS 0.031473f
C696 VTAIL.n87 VSUBS 0.029554f
C697 VTAIL.n88 VSUBS 0.015881f
C698 VTAIL.n89 VSUBS 0.037537f
C699 VTAIL.n90 VSUBS 0.016815f
C700 VTAIL.n91 VSUBS 0.484243f
C701 VTAIL.n92 VSUBS 0.015881f
C702 VTAIL.t0 VSUBS 0.081558f
C703 VTAIL.n93 VSUBS 0.119028f
C704 VTAIL.n94 VSUBS 0.02378f
C705 VTAIL.n95 VSUBS 0.028153f
C706 VTAIL.n96 VSUBS 0.037537f
C707 VTAIL.n97 VSUBS 0.016815f
C708 VTAIL.n98 VSUBS 0.015881f
C709 VTAIL.n99 VSUBS 0.029554f
C710 VTAIL.n100 VSUBS 0.029554f
C711 VTAIL.n101 VSUBS 0.015881f
C712 VTAIL.n102 VSUBS 0.016815f
C713 VTAIL.n103 VSUBS 0.037537f
C714 VTAIL.n104 VSUBS 0.087466f
C715 VTAIL.n105 VSUBS 0.016815f
C716 VTAIL.n106 VSUBS 0.015881f
C717 VTAIL.n107 VSUBS 0.068717f
C718 VTAIL.n108 VSUBS 0.043847f
C719 VTAIL.n109 VSUBS 0.938383f
C720 VTAIL.t4 VSUBS 0.106731f
C721 VTAIL.t2 VSUBS 0.106731f
C722 VTAIL.n110 VSUBS 0.569384f
C723 VTAIL.n111 VSUBS 0.560842f
C724 VP.n0 VSUBS 0.070281f
C725 VP.t9 VSUBS 0.471065f
C726 VP.n1 VSUBS 0.248835f
C727 VP.n2 VSUBS 0.070281f
C728 VP.n3 VSUBS 0.070281f
C729 VP.t7 VSUBS 0.471065f
C730 VP.t1 VSUBS 0.471065f
C731 VP.t8 VSUBS 0.471065f
C732 VP.n4 VSUBS 0.248835f
C733 VP.t0 VSUBS 0.486888f
C734 VP.n5 VSUBS 0.226158f
C735 VP.t5 VSUBS 0.471065f
C736 VP.n6 VSUBS 0.244935f
C737 VP.n7 VSUBS 0.015948f
C738 VP.n8 VSUBS 0.224196f
C739 VP.n9 VSUBS 0.070281f
C740 VP.n10 VSUBS 0.070281f
C741 VP.n11 VSUBS 0.015948f
C742 VP.n12 VSUBS 0.244935f
C743 VP.n13 VSUBS 0.241468f
C744 VP.n14 VSUBS 2.22059f
C745 VP.n15 VSUBS 2.29058f
C746 VP.t4 VSUBS 0.471065f
C747 VP.n16 VSUBS 0.241468f
C748 VP.t6 VSUBS 0.471065f
C749 VP.n17 VSUBS 0.244935f
C750 VP.n18 VSUBS 0.015948f
C751 VP.n19 VSUBS 0.070281f
C752 VP.n20 VSUBS 0.070281f
C753 VP.n21 VSUBS 0.070281f
C754 VP.n22 VSUBS 0.015948f
C755 VP.t3 VSUBS 0.471065f
C756 VP.n23 VSUBS 0.244935f
C757 VP.t2 VSUBS 0.471065f
C758 VP.n24 VSUBS 0.241468f
C759 VP.n25 VSUBS 0.054465f
.ends

