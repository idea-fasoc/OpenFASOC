* NGSPICE file created from diff_pair_sample_1436.ext - technology: sky130A

.subckt diff_pair_sample_1436 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VP.t0 VDD1.t6 w_n1480_n4314# sky130_fd_pr__pfet_01v8 ad=2.76045 pd=17.06 as=2.76045 ps=17.06 w=16.73 l=0.18
X1 B.t11 B.t9 B.t10 w_n1480_n4314# sky130_fd_pr__pfet_01v8 ad=6.5247 pd=34.24 as=0 ps=0 w=16.73 l=0.18
X2 VDD2.t7 VN.t0 VTAIL.t5 w_n1480_n4314# sky130_fd_pr__pfet_01v8 ad=2.76045 pd=17.06 as=6.5247 ps=34.24 w=16.73 l=0.18
X3 VDD2.t6 VN.t1 VTAIL.t1 w_n1480_n4314# sky130_fd_pr__pfet_01v8 ad=2.76045 pd=17.06 as=6.5247 ps=34.24 w=16.73 l=0.18
X4 VDD1.t5 VP.t1 VTAIL.t14 w_n1480_n4314# sky130_fd_pr__pfet_01v8 ad=2.76045 pd=17.06 as=2.76045 ps=17.06 w=16.73 l=0.18
X5 VTAIL.t6 VN.t2 VDD2.t5 w_n1480_n4314# sky130_fd_pr__pfet_01v8 ad=2.76045 pd=17.06 as=2.76045 ps=17.06 w=16.73 l=0.18
X6 VDD2.t4 VN.t3 VTAIL.t4 w_n1480_n4314# sky130_fd_pr__pfet_01v8 ad=2.76045 pd=17.06 as=2.76045 ps=17.06 w=16.73 l=0.18
X7 VTAIL.t0 VN.t4 VDD2.t3 w_n1480_n4314# sky130_fd_pr__pfet_01v8 ad=6.5247 pd=34.24 as=2.76045 ps=17.06 w=16.73 l=0.18
X8 B.t8 B.t6 B.t7 w_n1480_n4314# sky130_fd_pr__pfet_01v8 ad=6.5247 pd=34.24 as=0 ps=0 w=16.73 l=0.18
X9 VTAIL.t7 VN.t5 VDD2.t2 w_n1480_n4314# sky130_fd_pr__pfet_01v8 ad=6.5247 pd=34.24 as=2.76045 ps=17.06 w=16.73 l=0.18
X10 VTAIL.t13 VP.t2 VDD1.t3 w_n1480_n4314# sky130_fd_pr__pfet_01v8 ad=6.5247 pd=34.24 as=2.76045 ps=17.06 w=16.73 l=0.18
X11 VDD1.t2 VP.t3 VTAIL.t12 w_n1480_n4314# sky130_fd_pr__pfet_01v8 ad=2.76045 pd=17.06 as=2.76045 ps=17.06 w=16.73 l=0.18
X12 VTAIL.t11 VP.t4 VDD1.t0 w_n1480_n4314# sky130_fd_pr__pfet_01v8 ad=2.76045 pd=17.06 as=2.76045 ps=17.06 w=16.73 l=0.18
X13 VTAIL.t10 VP.t5 VDD1.t7 w_n1480_n4314# sky130_fd_pr__pfet_01v8 ad=6.5247 pd=34.24 as=2.76045 ps=17.06 w=16.73 l=0.18
X14 VDD1.t1 VP.t6 VTAIL.t9 w_n1480_n4314# sky130_fd_pr__pfet_01v8 ad=2.76045 pd=17.06 as=6.5247 ps=34.24 w=16.73 l=0.18
X15 B.t5 B.t3 B.t4 w_n1480_n4314# sky130_fd_pr__pfet_01v8 ad=6.5247 pd=34.24 as=0 ps=0 w=16.73 l=0.18
X16 VDD1.t4 VP.t7 VTAIL.t8 w_n1480_n4314# sky130_fd_pr__pfet_01v8 ad=2.76045 pd=17.06 as=6.5247 ps=34.24 w=16.73 l=0.18
X17 VDD2.t1 VN.t6 VTAIL.t2 w_n1480_n4314# sky130_fd_pr__pfet_01v8 ad=2.76045 pd=17.06 as=2.76045 ps=17.06 w=16.73 l=0.18
X18 VTAIL.t3 VN.t7 VDD2.t0 w_n1480_n4314# sky130_fd_pr__pfet_01v8 ad=2.76045 pd=17.06 as=2.76045 ps=17.06 w=16.73 l=0.18
X19 B.t2 B.t0 B.t1 w_n1480_n4314# sky130_fd_pr__pfet_01v8 ad=6.5247 pd=34.24 as=0 ps=0 w=16.73 l=0.18
R0 VP.n13 VP.t7 2454.06
R1 VP.n9 VP.t5 2454.06
R2 VP.n2 VP.t2 2454.06
R3 VP.n6 VP.t6 2454.06
R4 VP.n12 VP.t0 2415.36
R5 VP.n10 VP.t1 2415.36
R6 VP.n3 VP.t3 2415.36
R7 VP.n5 VP.t4 2415.36
R8 VP.n2 VP.n1 161.489
R9 VP.n14 VP.n13 161.3
R10 VP.n4 VP.n1 161.3
R11 VP.n7 VP.n6 161.3
R12 VP.n11 VP.n0 161.3
R13 VP.n9 VP.n8 161.3
R14 VP.n8 VP.n7 43.1823
R15 VP.n11 VP.n10 37.246
R16 VP.n12 VP.n11 37.246
R17 VP.n4 VP.n3 37.246
R18 VP.n5 VP.n4 37.246
R19 VP.n10 VP.n9 35.7853
R20 VP.n13 VP.n12 35.7853
R21 VP.n3 VP.n2 35.7853
R22 VP.n6 VP.n5 35.7853
R23 VP.n7 VP.n1 0.189894
R24 VP.n8 VP.n0 0.189894
R25 VP.n14 VP.n0 0.189894
R26 VP VP.n14 0.0516364
R27 VDD1 VDD1.n0 68.3125
R28 VDD1.n3 VDD1.n2 68.1987
R29 VDD1.n3 VDD1.n1 68.1987
R30 VDD1.n5 VDD1.n4 68.0343
R31 VDD1.n5 VDD1.n3 40.6992
R32 VDD1.n4 VDD1.t0 1.94342
R33 VDD1.n4 VDD1.t1 1.94342
R34 VDD1.n0 VDD1.t3 1.94342
R35 VDD1.n0 VDD1.t2 1.94342
R36 VDD1.n2 VDD1.t6 1.94342
R37 VDD1.n2 VDD1.t4 1.94342
R38 VDD1.n1 VDD1.t7 1.94342
R39 VDD1.n1 VDD1.t5 1.94342
R40 VDD1 VDD1.n5 0.162138
R41 VTAIL.n754 VTAIL.n666 756.745
R42 VTAIL.n90 VTAIL.n2 756.745
R43 VTAIL.n184 VTAIL.n96 756.745
R44 VTAIL.n280 VTAIL.n192 756.745
R45 VTAIL.n660 VTAIL.n572 756.745
R46 VTAIL.n564 VTAIL.n476 756.745
R47 VTAIL.n470 VTAIL.n382 756.745
R48 VTAIL.n374 VTAIL.n286 756.745
R49 VTAIL.n697 VTAIL.n696 585
R50 VTAIL.n694 VTAIL.n693 585
R51 VTAIL.n703 VTAIL.n702 585
R52 VTAIL.n705 VTAIL.n704 585
R53 VTAIL.n690 VTAIL.n689 585
R54 VTAIL.n711 VTAIL.n710 585
R55 VTAIL.n713 VTAIL.n712 585
R56 VTAIL.n686 VTAIL.n685 585
R57 VTAIL.n719 VTAIL.n718 585
R58 VTAIL.n721 VTAIL.n720 585
R59 VTAIL.n682 VTAIL.n681 585
R60 VTAIL.n727 VTAIL.n726 585
R61 VTAIL.n729 VTAIL.n728 585
R62 VTAIL.n678 VTAIL.n677 585
R63 VTAIL.n735 VTAIL.n734 585
R64 VTAIL.n738 VTAIL.n737 585
R65 VTAIL.n736 VTAIL.n674 585
R66 VTAIL.n743 VTAIL.n673 585
R67 VTAIL.n745 VTAIL.n744 585
R68 VTAIL.n747 VTAIL.n746 585
R69 VTAIL.n670 VTAIL.n669 585
R70 VTAIL.n753 VTAIL.n752 585
R71 VTAIL.n755 VTAIL.n754 585
R72 VTAIL.n33 VTAIL.n32 585
R73 VTAIL.n30 VTAIL.n29 585
R74 VTAIL.n39 VTAIL.n38 585
R75 VTAIL.n41 VTAIL.n40 585
R76 VTAIL.n26 VTAIL.n25 585
R77 VTAIL.n47 VTAIL.n46 585
R78 VTAIL.n49 VTAIL.n48 585
R79 VTAIL.n22 VTAIL.n21 585
R80 VTAIL.n55 VTAIL.n54 585
R81 VTAIL.n57 VTAIL.n56 585
R82 VTAIL.n18 VTAIL.n17 585
R83 VTAIL.n63 VTAIL.n62 585
R84 VTAIL.n65 VTAIL.n64 585
R85 VTAIL.n14 VTAIL.n13 585
R86 VTAIL.n71 VTAIL.n70 585
R87 VTAIL.n74 VTAIL.n73 585
R88 VTAIL.n72 VTAIL.n10 585
R89 VTAIL.n79 VTAIL.n9 585
R90 VTAIL.n81 VTAIL.n80 585
R91 VTAIL.n83 VTAIL.n82 585
R92 VTAIL.n6 VTAIL.n5 585
R93 VTAIL.n89 VTAIL.n88 585
R94 VTAIL.n91 VTAIL.n90 585
R95 VTAIL.n127 VTAIL.n126 585
R96 VTAIL.n124 VTAIL.n123 585
R97 VTAIL.n133 VTAIL.n132 585
R98 VTAIL.n135 VTAIL.n134 585
R99 VTAIL.n120 VTAIL.n119 585
R100 VTAIL.n141 VTAIL.n140 585
R101 VTAIL.n143 VTAIL.n142 585
R102 VTAIL.n116 VTAIL.n115 585
R103 VTAIL.n149 VTAIL.n148 585
R104 VTAIL.n151 VTAIL.n150 585
R105 VTAIL.n112 VTAIL.n111 585
R106 VTAIL.n157 VTAIL.n156 585
R107 VTAIL.n159 VTAIL.n158 585
R108 VTAIL.n108 VTAIL.n107 585
R109 VTAIL.n165 VTAIL.n164 585
R110 VTAIL.n168 VTAIL.n167 585
R111 VTAIL.n166 VTAIL.n104 585
R112 VTAIL.n173 VTAIL.n103 585
R113 VTAIL.n175 VTAIL.n174 585
R114 VTAIL.n177 VTAIL.n176 585
R115 VTAIL.n100 VTAIL.n99 585
R116 VTAIL.n183 VTAIL.n182 585
R117 VTAIL.n185 VTAIL.n184 585
R118 VTAIL.n223 VTAIL.n222 585
R119 VTAIL.n220 VTAIL.n219 585
R120 VTAIL.n229 VTAIL.n228 585
R121 VTAIL.n231 VTAIL.n230 585
R122 VTAIL.n216 VTAIL.n215 585
R123 VTAIL.n237 VTAIL.n236 585
R124 VTAIL.n239 VTAIL.n238 585
R125 VTAIL.n212 VTAIL.n211 585
R126 VTAIL.n245 VTAIL.n244 585
R127 VTAIL.n247 VTAIL.n246 585
R128 VTAIL.n208 VTAIL.n207 585
R129 VTAIL.n253 VTAIL.n252 585
R130 VTAIL.n255 VTAIL.n254 585
R131 VTAIL.n204 VTAIL.n203 585
R132 VTAIL.n261 VTAIL.n260 585
R133 VTAIL.n264 VTAIL.n263 585
R134 VTAIL.n262 VTAIL.n200 585
R135 VTAIL.n269 VTAIL.n199 585
R136 VTAIL.n271 VTAIL.n270 585
R137 VTAIL.n273 VTAIL.n272 585
R138 VTAIL.n196 VTAIL.n195 585
R139 VTAIL.n279 VTAIL.n278 585
R140 VTAIL.n281 VTAIL.n280 585
R141 VTAIL.n661 VTAIL.n660 585
R142 VTAIL.n659 VTAIL.n658 585
R143 VTAIL.n576 VTAIL.n575 585
R144 VTAIL.n653 VTAIL.n652 585
R145 VTAIL.n651 VTAIL.n650 585
R146 VTAIL.n649 VTAIL.n579 585
R147 VTAIL.n583 VTAIL.n580 585
R148 VTAIL.n644 VTAIL.n643 585
R149 VTAIL.n642 VTAIL.n641 585
R150 VTAIL.n585 VTAIL.n584 585
R151 VTAIL.n636 VTAIL.n635 585
R152 VTAIL.n634 VTAIL.n633 585
R153 VTAIL.n589 VTAIL.n588 585
R154 VTAIL.n628 VTAIL.n627 585
R155 VTAIL.n626 VTAIL.n625 585
R156 VTAIL.n593 VTAIL.n592 585
R157 VTAIL.n620 VTAIL.n619 585
R158 VTAIL.n618 VTAIL.n617 585
R159 VTAIL.n597 VTAIL.n596 585
R160 VTAIL.n612 VTAIL.n611 585
R161 VTAIL.n610 VTAIL.n609 585
R162 VTAIL.n601 VTAIL.n600 585
R163 VTAIL.n604 VTAIL.n603 585
R164 VTAIL.n565 VTAIL.n564 585
R165 VTAIL.n563 VTAIL.n562 585
R166 VTAIL.n480 VTAIL.n479 585
R167 VTAIL.n557 VTAIL.n556 585
R168 VTAIL.n555 VTAIL.n554 585
R169 VTAIL.n553 VTAIL.n483 585
R170 VTAIL.n487 VTAIL.n484 585
R171 VTAIL.n548 VTAIL.n547 585
R172 VTAIL.n546 VTAIL.n545 585
R173 VTAIL.n489 VTAIL.n488 585
R174 VTAIL.n540 VTAIL.n539 585
R175 VTAIL.n538 VTAIL.n537 585
R176 VTAIL.n493 VTAIL.n492 585
R177 VTAIL.n532 VTAIL.n531 585
R178 VTAIL.n530 VTAIL.n529 585
R179 VTAIL.n497 VTAIL.n496 585
R180 VTAIL.n524 VTAIL.n523 585
R181 VTAIL.n522 VTAIL.n521 585
R182 VTAIL.n501 VTAIL.n500 585
R183 VTAIL.n516 VTAIL.n515 585
R184 VTAIL.n514 VTAIL.n513 585
R185 VTAIL.n505 VTAIL.n504 585
R186 VTAIL.n508 VTAIL.n507 585
R187 VTAIL.n471 VTAIL.n470 585
R188 VTAIL.n469 VTAIL.n468 585
R189 VTAIL.n386 VTAIL.n385 585
R190 VTAIL.n463 VTAIL.n462 585
R191 VTAIL.n461 VTAIL.n460 585
R192 VTAIL.n459 VTAIL.n389 585
R193 VTAIL.n393 VTAIL.n390 585
R194 VTAIL.n454 VTAIL.n453 585
R195 VTAIL.n452 VTAIL.n451 585
R196 VTAIL.n395 VTAIL.n394 585
R197 VTAIL.n446 VTAIL.n445 585
R198 VTAIL.n444 VTAIL.n443 585
R199 VTAIL.n399 VTAIL.n398 585
R200 VTAIL.n438 VTAIL.n437 585
R201 VTAIL.n436 VTAIL.n435 585
R202 VTAIL.n403 VTAIL.n402 585
R203 VTAIL.n430 VTAIL.n429 585
R204 VTAIL.n428 VTAIL.n427 585
R205 VTAIL.n407 VTAIL.n406 585
R206 VTAIL.n422 VTAIL.n421 585
R207 VTAIL.n420 VTAIL.n419 585
R208 VTAIL.n411 VTAIL.n410 585
R209 VTAIL.n414 VTAIL.n413 585
R210 VTAIL.n375 VTAIL.n374 585
R211 VTAIL.n373 VTAIL.n372 585
R212 VTAIL.n290 VTAIL.n289 585
R213 VTAIL.n367 VTAIL.n366 585
R214 VTAIL.n365 VTAIL.n364 585
R215 VTAIL.n363 VTAIL.n293 585
R216 VTAIL.n297 VTAIL.n294 585
R217 VTAIL.n358 VTAIL.n357 585
R218 VTAIL.n356 VTAIL.n355 585
R219 VTAIL.n299 VTAIL.n298 585
R220 VTAIL.n350 VTAIL.n349 585
R221 VTAIL.n348 VTAIL.n347 585
R222 VTAIL.n303 VTAIL.n302 585
R223 VTAIL.n342 VTAIL.n341 585
R224 VTAIL.n340 VTAIL.n339 585
R225 VTAIL.n307 VTAIL.n306 585
R226 VTAIL.n334 VTAIL.n333 585
R227 VTAIL.n332 VTAIL.n331 585
R228 VTAIL.n311 VTAIL.n310 585
R229 VTAIL.n326 VTAIL.n325 585
R230 VTAIL.n324 VTAIL.n323 585
R231 VTAIL.n315 VTAIL.n314 585
R232 VTAIL.n318 VTAIL.n317 585
R233 VTAIL.t9 VTAIL.n602 327.466
R234 VTAIL.t13 VTAIL.n506 327.466
R235 VTAIL.t1 VTAIL.n412 327.466
R236 VTAIL.t7 VTAIL.n316 327.466
R237 VTAIL.t5 VTAIL.n695 327.466
R238 VTAIL.t0 VTAIL.n31 327.466
R239 VTAIL.t8 VTAIL.n125 327.466
R240 VTAIL.t10 VTAIL.n221 327.466
R241 VTAIL.n696 VTAIL.n693 171.744
R242 VTAIL.n703 VTAIL.n693 171.744
R243 VTAIL.n704 VTAIL.n703 171.744
R244 VTAIL.n704 VTAIL.n689 171.744
R245 VTAIL.n711 VTAIL.n689 171.744
R246 VTAIL.n712 VTAIL.n711 171.744
R247 VTAIL.n712 VTAIL.n685 171.744
R248 VTAIL.n719 VTAIL.n685 171.744
R249 VTAIL.n720 VTAIL.n719 171.744
R250 VTAIL.n720 VTAIL.n681 171.744
R251 VTAIL.n727 VTAIL.n681 171.744
R252 VTAIL.n728 VTAIL.n727 171.744
R253 VTAIL.n728 VTAIL.n677 171.744
R254 VTAIL.n735 VTAIL.n677 171.744
R255 VTAIL.n737 VTAIL.n735 171.744
R256 VTAIL.n737 VTAIL.n736 171.744
R257 VTAIL.n736 VTAIL.n673 171.744
R258 VTAIL.n745 VTAIL.n673 171.744
R259 VTAIL.n746 VTAIL.n745 171.744
R260 VTAIL.n746 VTAIL.n669 171.744
R261 VTAIL.n753 VTAIL.n669 171.744
R262 VTAIL.n754 VTAIL.n753 171.744
R263 VTAIL.n32 VTAIL.n29 171.744
R264 VTAIL.n39 VTAIL.n29 171.744
R265 VTAIL.n40 VTAIL.n39 171.744
R266 VTAIL.n40 VTAIL.n25 171.744
R267 VTAIL.n47 VTAIL.n25 171.744
R268 VTAIL.n48 VTAIL.n47 171.744
R269 VTAIL.n48 VTAIL.n21 171.744
R270 VTAIL.n55 VTAIL.n21 171.744
R271 VTAIL.n56 VTAIL.n55 171.744
R272 VTAIL.n56 VTAIL.n17 171.744
R273 VTAIL.n63 VTAIL.n17 171.744
R274 VTAIL.n64 VTAIL.n63 171.744
R275 VTAIL.n64 VTAIL.n13 171.744
R276 VTAIL.n71 VTAIL.n13 171.744
R277 VTAIL.n73 VTAIL.n71 171.744
R278 VTAIL.n73 VTAIL.n72 171.744
R279 VTAIL.n72 VTAIL.n9 171.744
R280 VTAIL.n81 VTAIL.n9 171.744
R281 VTAIL.n82 VTAIL.n81 171.744
R282 VTAIL.n82 VTAIL.n5 171.744
R283 VTAIL.n89 VTAIL.n5 171.744
R284 VTAIL.n90 VTAIL.n89 171.744
R285 VTAIL.n126 VTAIL.n123 171.744
R286 VTAIL.n133 VTAIL.n123 171.744
R287 VTAIL.n134 VTAIL.n133 171.744
R288 VTAIL.n134 VTAIL.n119 171.744
R289 VTAIL.n141 VTAIL.n119 171.744
R290 VTAIL.n142 VTAIL.n141 171.744
R291 VTAIL.n142 VTAIL.n115 171.744
R292 VTAIL.n149 VTAIL.n115 171.744
R293 VTAIL.n150 VTAIL.n149 171.744
R294 VTAIL.n150 VTAIL.n111 171.744
R295 VTAIL.n157 VTAIL.n111 171.744
R296 VTAIL.n158 VTAIL.n157 171.744
R297 VTAIL.n158 VTAIL.n107 171.744
R298 VTAIL.n165 VTAIL.n107 171.744
R299 VTAIL.n167 VTAIL.n165 171.744
R300 VTAIL.n167 VTAIL.n166 171.744
R301 VTAIL.n166 VTAIL.n103 171.744
R302 VTAIL.n175 VTAIL.n103 171.744
R303 VTAIL.n176 VTAIL.n175 171.744
R304 VTAIL.n176 VTAIL.n99 171.744
R305 VTAIL.n183 VTAIL.n99 171.744
R306 VTAIL.n184 VTAIL.n183 171.744
R307 VTAIL.n222 VTAIL.n219 171.744
R308 VTAIL.n229 VTAIL.n219 171.744
R309 VTAIL.n230 VTAIL.n229 171.744
R310 VTAIL.n230 VTAIL.n215 171.744
R311 VTAIL.n237 VTAIL.n215 171.744
R312 VTAIL.n238 VTAIL.n237 171.744
R313 VTAIL.n238 VTAIL.n211 171.744
R314 VTAIL.n245 VTAIL.n211 171.744
R315 VTAIL.n246 VTAIL.n245 171.744
R316 VTAIL.n246 VTAIL.n207 171.744
R317 VTAIL.n253 VTAIL.n207 171.744
R318 VTAIL.n254 VTAIL.n253 171.744
R319 VTAIL.n254 VTAIL.n203 171.744
R320 VTAIL.n261 VTAIL.n203 171.744
R321 VTAIL.n263 VTAIL.n261 171.744
R322 VTAIL.n263 VTAIL.n262 171.744
R323 VTAIL.n262 VTAIL.n199 171.744
R324 VTAIL.n271 VTAIL.n199 171.744
R325 VTAIL.n272 VTAIL.n271 171.744
R326 VTAIL.n272 VTAIL.n195 171.744
R327 VTAIL.n279 VTAIL.n195 171.744
R328 VTAIL.n280 VTAIL.n279 171.744
R329 VTAIL.n660 VTAIL.n659 171.744
R330 VTAIL.n659 VTAIL.n575 171.744
R331 VTAIL.n652 VTAIL.n575 171.744
R332 VTAIL.n652 VTAIL.n651 171.744
R333 VTAIL.n651 VTAIL.n579 171.744
R334 VTAIL.n583 VTAIL.n579 171.744
R335 VTAIL.n643 VTAIL.n583 171.744
R336 VTAIL.n643 VTAIL.n642 171.744
R337 VTAIL.n642 VTAIL.n584 171.744
R338 VTAIL.n635 VTAIL.n584 171.744
R339 VTAIL.n635 VTAIL.n634 171.744
R340 VTAIL.n634 VTAIL.n588 171.744
R341 VTAIL.n627 VTAIL.n588 171.744
R342 VTAIL.n627 VTAIL.n626 171.744
R343 VTAIL.n626 VTAIL.n592 171.744
R344 VTAIL.n619 VTAIL.n592 171.744
R345 VTAIL.n619 VTAIL.n618 171.744
R346 VTAIL.n618 VTAIL.n596 171.744
R347 VTAIL.n611 VTAIL.n596 171.744
R348 VTAIL.n611 VTAIL.n610 171.744
R349 VTAIL.n610 VTAIL.n600 171.744
R350 VTAIL.n603 VTAIL.n600 171.744
R351 VTAIL.n564 VTAIL.n563 171.744
R352 VTAIL.n563 VTAIL.n479 171.744
R353 VTAIL.n556 VTAIL.n479 171.744
R354 VTAIL.n556 VTAIL.n555 171.744
R355 VTAIL.n555 VTAIL.n483 171.744
R356 VTAIL.n487 VTAIL.n483 171.744
R357 VTAIL.n547 VTAIL.n487 171.744
R358 VTAIL.n547 VTAIL.n546 171.744
R359 VTAIL.n546 VTAIL.n488 171.744
R360 VTAIL.n539 VTAIL.n488 171.744
R361 VTAIL.n539 VTAIL.n538 171.744
R362 VTAIL.n538 VTAIL.n492 171.744
R363 VTAIL.n531 VTAIL.n492 171.744
R364 VTAIL.n531 VTAIL.n530 171.744
R365 VTAIL.n530 VTAIL.n496 171.744
R366 VTAIL.n523 VTAIL.n496 171.744
R367 VTAIL.n523 VTAIL.n522 171.744
R368 VTAIL.n522 VTAIL.n500 171.744
R369 VTAIL.n515 VTAIL.n500 171.744
R370 VTAIL.n515 VTAIL.n514 171.744
R371 VTAIL.n514 VTAIL.n504 171.744
R372 VTAIL.n507 VTAIL.n504 171.744
R373 VTAIL.n470 VTAIL.n469 171.744
R374 VTAIL.n469 VTAIL.n385 171.744
R375 VTAIL.n462 VTAIL.n385 171.744
R376 VTAIL.n462 VTAIL.n461 171.744
R377 VTAIL.n461 VTAIL.n389 171.744
R378 VTAIL.n393 VTAIL.n389 171.744
R379 VTAIL.n453 VTAIL.n393 171.744
R380 VTAIL.n453 VTAIL.n452 171.744
R381 VTAIL.n452 VTAIL.n394 171.744
R382 VTAIL.n445 VTAIL.n394 171.744
R383 VTAIL.n445 VTAIL.n444 171.744
R384 VTAIL.n444 VTAIL.n398 171.744
R385 VTAIL.n437 VTAIL.n398 171.744
R386 VTAIL.n437 VTAIL.n436 171.744
R387 VTAIL.n436 VTAIL.n402 171.744
R388 VTAIL.n429 VTAIL.n402 171.744
R389 VTAIL.n429 VTAIL.n428 171.744
R390 VTAIL.n428 VTAIL.n406 171.744
R391 VTAIL.n421 VTAIL.n406 171.744
R392 VTAIL.n421 VTAIL.n420 171.744
R393 VTAIL.n420 VTAIL.n410 171.744
R394 VTAIL.n413 VTAIL.n410 171.744
R395 VTAIL.n374 VTAIL.n373 171.744
R396 VTAIL.n373 VTAIL.n289 171.744
R397 VTAIL.n366 VTAIL.n289 171.744
R398 VTAIL.n366 VTAIL.n365 171.744
R399 VTAIL.n365 VTAIL.n293 171.744
R400 VTAIL.n297 VTAIL.n293 171.744
R401 VTAIL.n357 VTAIL.n297 171.744
R402 VTAIL.n357 VTAIL.n356 171.744
R403 VTAIL.n356 VTAIL.n298 171.744
R404 VTAIL.n349 VTAIL.n298 171.744
R405 VTAIL.n349 VTAIL.n348 171.744
R406 VTAIL.n348 VTAIL.n302 171.744
R407 VTAIL.n341 VTAIL.n302 171.744
R408 VTAIL.n341 VTAIL.n340 171.744
R409 VTAIL.n340 VTAIL.n306 171.744
R410 VTAIL.n333 VTAIL.n306 171.744
R411 VTAIL.n333 VTAIL.n332 171.744
R412 VTAIL.n332 VTAIL.n310 171.744
R413 VTAIL.n325 VTAIL.n310 171.744
R414 VTAIL.n325 VTAIL.n324 171.744
R415 VTAIL.n324 VTAIL.n314 171.744
R416 VTAIL.n317 VTAIL.n314 171.744
R417 VTAIL.n696 VTAIL.t5 85.8723
R418 VTAIL.n32 VTAIL.t0 85.8723
R419 VTAIL.n126 VTAIL.t8 85.8723
R420 VTAIL.n222 VTAIL.t10 85.8723
R421 VTAIL.n603 VTAIL.t9 85.8723
R422 VTAIL.n507 VTAIL.t13 85.8723
R423 VTAIL.n413 VTAIL.t1 85.8723
R424 VTAIL.n317 VTAIL.t7 85.8723
R425 VTAIL.n571 VTAIL.n570 51.3557
R426 VTAIL.n381 VTAIL.n380 51.3557
R427 VTAIL.n1 VTAIL.n0 51.3555
R428 VTAIL.n191 VTAIL.n190 51.3555
R429 VTAIL.n759 VTAIL.n758 30.8278
R430 VTAIL.n95 VTAIL.n94 30.8278
R431 VTAIL.n189 VTAIL.n188 30.8278
R432 VTAIL.n285 VTAIL.n284 30.8278
R433 VTAIL.n665 VTAIL.n664 30.8278
R434 VTAIL.n569 VTAIL.n568 30.8278
R435 VTAIL.n475 VTAIL.n474 30.8278
R436 VTAIL.n379 VTAIL.n378 30.8278
R437 VTAIL.n759 VTAIL.n665 27.2289
R438 VTAIL.n379 VTAIL.n285 27.2289
R439 VTAIL.n697 VTAIL.n695 16.3895
R440 VTAIL.n33 VTAIL.n31 16.3895
R441 VTAIL.n127 VTAIL.n125 16.3895
R442 VTAIL.n223 VTAIL.n221 16.3895
R443 VTAIL.n604 VTAIL.n602 16.3895
R444 VTAIL.n508 VTAIL.n506 16.3895
R445 VTAIL.n414 VTAIL.n412 16.3895
R446 VTAIL.n318 VTAIL.n316 16.3895
R447 VTAIL.n744 VTAIL.n743 13.1884
R448 VTAIL.n80 VTAIL.n79 13.1884
R449 VTAIL.n174 VTAIL.n173 13.1884
R450 VTAIL.n270 VTAIL.n269 13.1884
R451 VTAIL.n650 VTAIL.n649 13.1884
R452 VTAIL.n554 VTAIL.n553 13.1884
R453 VTAIL.n460 VTAIL.n459 13.1884
R454 VTAIL.n364 VTAIL.n363 13.1884
R455 VTAIL.n698 VTAIL.n694 12.8005
R456 VTAIL.n742 VTAIL.n674 12.8005
R457 VTAIL.n747 VTAIL.n672 12.8005
R458 VTAIL.n34 VTAIL.n30 12.8005
R459 VTAIL.n78 VTAIL.n10 12.8005
R460 VTAIL.n83 VTAIL.n8 12.8005
R461 VTAIL.n128 VTAIL.n124 12.8005
R462 VTAIL.n172 VTAIL.n104 12.8005
R463 VTAIL.n177 VTAIL.n102 12.8005
R464 VTAIL.n224 VTAIL.n220 12.8005
R465 VTAIL.n268 VTAIL.n200 12.8005
R466 VTAIL.n273 VTAIL.n198 12.8005
R467 VTAIL.n653 VTAIL.n578 12.8005
R468 VTAIL.n648 VTAIL.n580 12.8005
R469 VTAIL.n605 VTAIL.n601 12.8005
R470 VTAIL.n557 VTAIL.n482 12.8005
R471 VTAIL.n552 VTAIL.n484 12.8005
R472 VTAIL.n509 VTAIL.n505 12.8005
R473 VTAIL.n463 VTAIL.n388 12.8005
R474 VTAIL.n458 VTAIL.n390 12.8005
R475 VTAIL.n415 VTAIL.n411 12.8005
R476 VTAIL.n367 VTAIL.n292 12.8005
R477 VTAIL.n362 VTAIL.n294 12.8005
R478 VTAIL.n319 VTAIL.n315 12.8005
R479 VTAIL.n702 VTAIL.n701 12.0247
R480 VTAIL.n739 VTAIL.n738 12.0247
R481 VTAIL.n748 VTAIL.n670 12.0247
R482 VTAIL.n38 VTAIL.n37 12.0247
R483 VTAIL.n75 VTAIL.n74 12.0247
R484 VTAIL.n84 VTAIL.n6 12.0247
R485 VTAIL.n132 VTAIL.n131 12.0247
R486 VTAIL.n169 VTAIL.n168 12.0247
R487 VTAIL.n178 VTAIL.n100 12.0247
R488 VTAIL.n228 VTAIL.n227 12.0247
R489 VTAIL.n265 VTAIL.n264 12.0247
R490 VTAIL.n274 VTAIL.n196 12.0247
R491 VTAIL.n654 VTAIL.n576 12.0247
R492 VTAIL.n645 VTAIL.n644 12.0247
R493 VTAIL.n609 VTAIL.n608 12.0247
R494 VTAIL.n558 VTAIL.n480 12.0247
R495 VTAIL.n549 VTAIL.n548 12.0247
R496 VTAIL.n513 VTAIL.n512 12.0247
R497 VTAIL.n464 VTAIL.n386 12.0247
R498 VTAIL.n455 VTAIL.n454 12.0247
R499 VTAIL.n419 VTAIL.n418 12.0247
R500 VTAIL.n368 VTAIL.n290 12.0247
R501 VTAIL.n359 VTAIL.n358 12.0247
R502 VTAIL.n323 VTAIL.n322 12.0247
R503 VTAIL.n705 VTAIL.n692 11.249
R504 VTAIL.n734 VTAIL.n676 11.249
R505 VTAIL.n752 VTAIL.n751 11.249
R506 VTAIL.n41 VTAIL.n28 11.249
R507 VTAIL.n70 VTAIL.n12 11.249
R508 VTAIL.n88 VTAIL.n87 11.249
R509 VTAIL.n135 VTAIL.n122 11.249
R510 VTAIL.n164 VTAIL.n106 11.249
R511 VTAIL.n182 VTAIL.n181 11.249
R512 VTAIL.n231 VTAIL.n218 11.249
R513 VTAIL.n260 VTAIL.n202 11.249
R514 VTAIL.n278 VTAIL.n277 11.249
R515 VTAIL.n658 VTAIL.n657 11.249
R516 VTAIL.n641 VTAIL.n582 11.249
R517 VTAIL.n612 VTAIL.n599 11.249
R518 VTAIL.n562 VTAIL.n561 11.249
R519 VTAIL.n545 VTAIL.n486 11.249
R520 VTAIL.n516 VTAIL.n503 11.249
R521 VTAIL.n468 VTAIL.n467 11.249
R522 VTAIL.n451 VTAIL.n392 11.249
R523 VTAIL.n422 VTAIL.n409 11.249
R524 VTAIL.n372 VTAIL.n371 11.249
R525 VTAIL.n355 VTAIL.n296 11.249
R526 VTAIL.n326 VTAIL.n313 11.249
R527 VTAIL.n706 VTAIL.n690 10.4732
R528 VTAIL.n733 VTAIL.n678 10.4732
R529 VTAIL.n755 VTAIL.n668 10.4732
R530 VTAIL.n42 VTAIL.n26 10.4732
R531 VTAIL.n69 VTAIL.n14 10.4732
R532 VTAIL.n91 VTAIL.n4 10.4732
R533 VTAIL.n136 VTAIL.n120 10.4732
R534 VTAIL.n163 VTAIL.n108 10.4732
R535 VTAIL.n185 VTAIL.n98 10.4732
R536 VTAIL.n232 VTAIL.n216 10.4732
R537 VTAIL.n259 VTAIL.n204 10.4732
R538 VTAIL.n281 VTAIL.n194 10.4732
R539 VTAIL.n661 VTAIL.n574 10.4732
R540 VTAIL.n640 VTAIL.n585 10.4732
R541 VTAIL.n613 VTAIL.n597 10.4732
R542 VTAIL.n565 VTAIL.n478 10.4732
R543 VTAIL.n544 VTAIL.n489 10.4732
R544 VTAIL.n517 VTAIL.n501 10.4732
R545 VTAIL.n471 VTAIL.n384 10.4732
R546 VTAIL.n450 VTAIL.n395 10.4732
R547 VTAIL.n423 VTAIL.n407 10.4732
R548 VTAIL.n375 VTAIL.n288 10.4732
R549 VTAIL.n354 VTAIL.n299 10.4732
R550 VTAIL.n327 VTAIL.n311 10.4732
R551 VTAIL.n710 VTAIL.n709 9.69747
R552 VTAIL.n730 VTAIL.n729 9.69747
R553 VTAIL.n756 VTAIL.n666 9.69747
R554 VTAIL.n46 VTAIL.n45 9.69747
R555 VTAIL.n66 VTAIL.n65 9.69747
R556 VTAIL.n92 VTAIL.n2 9.69747
R557 VTAIL.n140 VTAIL.n139 9.69747
R558 VTAIL.n160 VTAIL.n159 9.69747
R559 VTAIL.n186 VTAIL.n96 9.69747
R560 VTAIL.n236 VTAIL.n235 9.69747
R561 VTAIL.n256 VTAIL.n255 9.69747
R562 VTAIL.n282 VTAIL.n192 9.69747
R563 VTAIL.n662 VTAIL.n572 9.69747
R564 VTAIL.n637 VTAIL.n636 9.69747
R565 VTAIL.n617 VTAIL.n616 9.69747
R566 VTAIL.n566 VTAIL.n476 9.69747
R567 VTAIL.n541 VTAIL.n540 9.69747
R568 VTAIL.n521 VTAIL.n520 9.69747
R569 VTAIL.n472 VTAIL.n382 9.69747
R570 VTAIL.n447 VTAIL.n446 9.69747
R571 VTAIL.n427 VTAIL.n426 9.69747
R572 VTAIL.n376 VTAIL.n286 9.69747
R573 VTAIL.n351 VTAIL.n350 9.69747
R574 VTAIL.n331 VTAIL.n330 9.69747
R575 VTAIL.n758 VTAIL.n757 9.45567
R576 VTAIL.n94 VTAIL.n93 9.45567
R577 VTAIL.n188 VTAIL.n187 9.45567
R578 VTAIL.n284 VTAIL.n283 9.45567
R579 VTAIL.n664 VTAIL.n663 9.45567
R580 VTAIL.n568 VTAIL.n567 9.45567
R581 VTAIL.n474 VTAIL.n473 9.45567
R582 VTAIL.n378 VTAIL.n377 9.45567
R583 VTAIL.n757 VTAIL.n756 9.3005
R584 VTAIL.n668 VTAIL.n667 9.3005
R585 VTAIL.n751 VTAIL.n750 9.3005
R586 VTAIL.n749 VTAIL.n748 9.3005
R587 VTAIL.n672 VTAIL.n671 9.3005
R588 VTAIL.n717 VTAIL.n716 9.3005
R589 VTAIL.n715 VTAIL.n714 9.3005
R590 VTAIL.n688 VTAIL.n687 9.3005
R591 VTAIL.n709 VTAIL.n708 9.3005
R592 VTAIL.n707 VTAIL.n706 9.3005
R593 VTAIL.n692 VTAIL.n691 9.3005
R594 VTAIL.n701 VTAIL.n700 9.3005
R595 VTAIL.n699 VTAIL.n698 9.3005
R596 VTAIL.n684 VTAIL.n683 9.3005
R597 VTAIL.n723 VTAIL.n722 9.3005
R598 VTAIL.n725 VTAIL.n724 9.3005
R599 VTAIL.n680 VTAIL.n679 9.3005
R600 VTAIL.n731 VTAIL.n730 9.3005
R601 VTAIL.n733 VTAIL.n732 9.3005
R602 VTAIL.n676 VTAIL.n675 9.3005
R603 VTAIL.n740 VTAIL.n739 9.3005
R604 VTAIL.n742 VTAIL.n741 9.3005
R605 VTAIL.n93 VTAIL.n92 9.3005
R606 VTAIL.n4 VTAIL.n3 9.3005
R607 VTAIL.n87 VTAIL.n86 9.3005
R608 VTAIL.n85 VTAIL.n84 9.3005
R609 VTAIL.n8 VTAIL.n7 9.3005
R610 VTAIL.n53 VTAIL.n52 9.3005
R611 VTAIL.n51 VTAIL.n50 9.3005
R612 VTAIL.n24 VTAIL.n23 9.3005
R613 VTAIL.n45 VTAIL.n44 9.3005
R614 VTAIL.n43 VTAIL.n42 9.3005
R615 VTAIL.n28 VTAIL.n27 9.3005
R616 VTAIL.n37 VTAIL.n36 9.3005
R617 VTAIL.n35 VTAIL.n34 9.3005
R618 VTAIL.n20 VTAIL.n19 9.3005
R619 VTAIL.n59 VTAIL.n58 9.3005
R620 VTAIL.n61 VTAIL.n60 9.3005
R621 VTAIL.n16 VTAIL.n15 9.3005
R622 VTAIL.n67 VTAIL.n66 9.3005
R623 VTAIL.n69 VTAIL.n68 9.3005
R624 VTAIL.n12 VTAIL.n11 9.3005
R625 VTAIL.n76 VTAIL.n75 9.3005
R626 VTAIL.n78 VTAIL.n77 9.3005
R627 VTAIL.n187 VTAIL.n186 9.3005
R628 VTAIL.n98 VTAIL.n97 9.3005
R629 VTAIL.n181 VTAIL.n180 9.3005
R630 VTAIL.n179 VTAIL.n178 9.3005
R631 VTAIL.n102 VTAIL.n101 9.3005
R632 VTAIL.n147 VTAIL.n146 9.3005
R633 VTAIL.n145 VTAIL.n144 9.3005
R634 VTAIL.n118 VTAIL.n117 9.3005
R635 VTAIL.n139 VTAIL.n138 9.3005
R636 VTAIL.n137 VTAIL.n136 9.3005
R637 VTAIL.n122 VTAIL.n121 9.3005
R638 VTAIL.n131 VTAIL.n130 9.3005
R639 VTAIL.n129 VTAIL.n128 9.3005
R640 VTAIL.n114 VTAIL.n113 9.3005
R641 VTAIL.n153 VTAIL.n152 9.3005
R642 VTAIL.n155 VTAIL.n154 9.3005
R643 VTAIL.n110 VTAIL.n109 9.3005
R644 VTAIL.n161 VTAIL.n160 9.3005
R645 VTAIL.n163 VTAIL.n162 9.3005
R646 VTAIL.n106 VTAIL.n105 9.3005
R647 VTAIL.n170 VTAIL.n169 9.3005
R648 VTAIL.n172 VTAIL.n171 9.3005
R649 VTAIL.n283 VTAIL.n282 9.3005
R650 VTAIL.n194 VTAIL.n193 9.3005
R651 VTAIL.n277 VTAIL.n276 9.3005
R652 VTAIL.n275 VTAIL.n274 9.3005
R653 VTAIL.n198 VTAIL.n197 9.3005
R654 VTAIL.n243 VTAIL.n242 9.3005
R655 VTAIL.n241 VTAIL.n240 9.3005
R656 VTAIL.n214 VTAIL.n213 9.3005
R657 VTAIL.n235 VTAIL.n234 9.3005
R658 VTAIL.n233 VTAIL.n232 9.3005
R659 VTAIL.n218 VTAIL.n217 9.3005
R660 VTAIL.n227 VTAIL.n226 9.3005
R661 VTAIL.n225 VTAIL.n224 9.3005
R662 VTAIL.n210 VTAIL.n209 9.3005
R663 VTAIL.n249 VTAIL.n248 9.3005
R664 VTAIL.n251 VTAIL.n250 9.3005
R665 VTAIL.n206 VTAIL.n205 9.3005
R666 VTAIL.n257 VTAIL.n256 9.3005
R667 VTAIL.n259 VTAIL.n258 9.3005
R668 VTAIL.n202 VTAIL.n201 9.3005
R669 VTAIL.n266 VTAIL.n265 9.3005
R670 VTAIL.n268 VTAIL.n267 9.3005
R671 VTAIL.n630 VTAIL.n629 9.3005
R672 VTAIL.n632 VTAIL.n631 9.3005
R673 VTAIL.n587 VTAIL.n586 9.3005
R674 VTAIL.n638 VTAIL.n637 9.3005
R675 VTAIL.n640 VTAIL.n639 9.3005
R676 VTAIL.n582 VTAIL.n581 9.3005
R677 VTAIL.n646 VTAIL.n645 9.3005
R678 VTAIL.n648 VTAIL.n647 9.3005
R679 VTAIL.n663 VTAIL.n662 9.3005
R680 VTAIL.n574 VTAIL.n573 9.3005
R681 VTAIL.n657 VTAIL.n656 9.3005
R682 VTAIL.n655 VTAIL.n654 9.3005
R683 VTAIL.n578 VTAIL.n577 9.3005
R684 VTAIL.n591 VTAIL.n590 9.3005
R685 VTAIL.n624 VTAIL.n623 9.3005
R686 VTAIL.n622 VTAIL.n621 9.3005
R687 VTAIL.n595 VTAIL.n594 9.3005
R688 VTAIL.n616 VTAIL.n615 9.3005
R689 VTAIL.n614 VTAIL.n613 9.3005
R690 VTAIL.n599 VTAIL.n598 9.3005
R691 VTAIL.n608 VTAIL.n607 9.3005
R692 VTAIL.n606 VTAIL.n605 9.3005
R693 VTAIL.n534 VTAIL.n533 9.3005
R694 VTAIL.n536 VTAIL.n535 9.3005
R695 VTAIL.n491 VTAIL.n490 9.3005
R696 VTAIL.n542 VTAIL.n541 9.3005
R697 VTAIL.n544 VTAIL.n543 9.3005
R698 VTAIL.n486 VTAIL.n485 9.3005
R699 VTAIL.n550 VTAIL.n549 9.3005
R700 VTAIL.n552 VTAIL.n551 9.3005
R701 VTAIL.n567 VTAIL.n566 9.3005
R702 VTAIL.n478 VTAIL.n477 9.3005
R703 VTAIL.n561 VTAIL.n560 9.3005
R704 VTAIL.n559 VTAIL.n558 9.3005
R705 VTAIL.n482 VTAIL.n481 9.3005
R706 VTAIL.n495 VTAIL.n494 9.3005
R707 VTAIL.n528 VTAIL.n527 9.3005
R708 VTAIL.n526 VTAIL.n525 9.3005
R709 VTAIL.n499 VTAIL.n498 9.3005
R710 VTAIL.n520 VTAIL.n519 9.3005
R711 VTAIL.n518 VTAIL.n517 9.3005
R712 VTAIL.n503 VTAIL.n502 9.3005
R713 VTAIL.n512 VTAIL.n511 9.3005
R714 VTAIL.n510 VTAIL.n509 9.3005
R715 VTAIL.n440 VTAIL.n439 9.3005
R716 VTAIL.n442 VTAIL.n441 9.3005
R717 VTAIL.n397 VTAIL.n396 9.3005
R718 VTAIL.n448 VTAIL.n447 9.3005
R719 VTAIL.n450 VTAIL.n449 9.3005
R720 VTAIL.n392 VTAIL.n391 9.3005
R721 VTAIL.n456 VTAIL.n455 9.3005
R722 VTAIL.n458 VTAIL.n457 9.3005
R723 VTAIL.n473 VTAIL.n472 9.3005
R724 VTAIL.n384 VTAIL.n383 9.3005
R725 VTAIL.n467 VTAIL.n466 9.3005
R726 VTAIL.n465 VTAIL.n464 9.3005
R727 VTAIL.n388 VTAIL.n387 9.3005
R728 VTAIL.n401 VTAIL.n400 9.3005
R729 VTAIL.n434 VTAIL.n433 9.3005
R730 VTAIL.n432 VTAIL.n431 9.3005
R731 VTAIL.n405 VTAIL.n404 9.3005
R732 VTAIL.n426 VTAIL.n425 9.3005
R733 VTAIL.n424 VTAIL.n423 9.3005
R734 VTAIL.n409 VTAIL.n408 9.3005
R735 VTAIL.n418 VTAIL.n417 9.3005
R736 VTAIL.n416 VTAIL.n415 9.3005
R737 VTAIL.n344 VTAIL.n343 9.3005
R738 VTAIL.n346 VTAIL.n345 9.3005
R739 VTAIL.n301 VTAIL.n300 9.3005
R740 VTAIL.n352 VTAIL.n351 9.3005
R741 VTAIL.n354 VTAIL.n353 9.3005
R742 VTAIL.n296 VTAIL.n295 9.3005
R743 VTAIL.n360 VTAIL.n359 9.3005
R744 VTAIL.n362 VTAIL.n361 9.3005
R745 VTAIL.n377 VTAIL.n376 9.3005
R746 VTAIL.n288 VTAIL.n287 9.3005
R747 VTAIL.n371 VTAIL.n370 9.3005
R748 VTAIL.n369 VTAIL.n368 9.3005
R749 VTAIL.n292 VTAIL.n291 9.3005
R750 VTAIL.n305 VTAIL.n304 9.3005
R751 VTAIL.n338 VTAIL.n337 9.3005
R752 VTAIL.n336 VTAIL.n335 9.3005
R753 VTAIL.n309 VTAIL.n308 9.3005
R754 VTAIL.n330 VTAIL.n329 9.3005
R755 VTAIL.n328 VTAIL.n327 9.3005
R756 VTAIL.n313 VTAIL.n312 9.3005
R757 VTAIL.n322 VTAIL.n321 9.3005
R758 VTAIL.n320 VTAIL.n319 9.3005
R759 VTAIL.n713 VTAIL.n688 8.92171
R760 VTAIL.n726 VTAIL.n680 8.92171
R761 VTAIL.n49 VTAIL.n24 8.92171
R762 VTAIL.n62 VTAIL.n16 8.92171
R763 VTAIL.n143 VTAIL.n118 8.92171
R764 VTAIL.n156 VTAIL.n110 8.92171
R765 VTAIL.n239 VTAIL.n214 8.92171
R766 VTAIL.n252 VTAIL.n206 8.92171
R767 VTAIL.n633 VTAIL.n587 8.92171
R768 VTAIL.n620 VTAIL.n595 8.92171
R769 VTAIL.n537 VTAIL.n491 8.92171
R770 VTAIL.n524 VTAIL.n499 8.92171
R771 VTAIL.n443 VTAIL.n397 8.92171
R772 VTAIL.n430 VTAIL.n405 8.92171
R773 VTAIL.n347 VTAIL.n301 8.92171
R774 VTAIL.n334 VTAIL.n309 8.92171
R775 VTAIL.n714 VTAIL.n686 8.14595
R776 VTAIL.n725 VTAIL.n682 8.14595
R777 VTAIL.n50 VTAIL.n22 8.14595
R778 VTAIL.n61 VTAIL.n18 8.14595
R779 VTAIL.n144 VTAIL.n116 8.14595
R780 VTAIL.n155 VTAIL.n112 8.14595
R781 VTAIL.n240 VTAIL.n212 8.14595
R782 VTAIL.n251 VTAIL.n208 8.14595
R783 VTAIL.n632 VTAIL.n589 8.14595
R784 VTAIL.n621 VTAIL.n593 8.14595
R785 VTAIL.n536 VTAIL.n493 8.14595
R786 VTAIL.n525 VTAIL.n497 8.14595
R787 VTAIL.n442 VTAIL.n399 8.14595
R788 VTAIL.n431 VTAIL.n403 8.14595
R789 VTAIL.n346 VTAIL.n303 8.14595
R790 VTAIL.n335 VTAIL.n307 8.14595
R791 VTAIL.n718 VTAIL.n717 7.3702
R792 VTAIL.n722 VTAIL.n721 7.3702
R793 VTAIL.n54 VTAIL.n53 7.3702
R794 VTAIL.n58 VTAIL.n57 7.3702
R795 VTAIL.n148 VTAIL.n147 7.3702
R796 VTAIL.n152 VTAIL.n151 7.3702
R797 VTAIL.n244 VTAIL.n243 7.3702
R798 VTAIL.n248 VTAIL.n247 7.3702
R799 VTAIL.n629 VTAIL.n628 7.3702
R800 VTAIL.n625 VTAIL.n624 7.3702
R801 VTAIL.n533 VTAIL.n532 7.3702
R802 VTAIL.n529 VTAIL.n528 7.3702
R803 VTAIL.n439 VTAIL.n438 7.3702
R804 VTAIL.n435 VTAIL.n434 7.3702
R805 VTAIL.n343 VTAIL.n342 7.3702
R806 VTAIL.n339 VTAIL.n338 7.3702
R807 VTAIL.n718 VTAIL.n684 6.59444
R808 VTAIL.n721 VTAIL.n684 6.59444
R809 VTAIL.n54 VTAIL.n20 6.59444
R810 VTAIL.n57 VTAIL.n20 6.59444
R811 VTAIL.n148 VTAIL.n114 6.59444
R812 VTAIL.n151 VTAIL.n114 6.59444
R813 VTAIL.n244 VTAIL.n210 6.59444
R814 VTAIL.n247 VTAIL.n210 6.59444
R815 VTAIL.n628 VTAIL.n591 6.59444
R816 VTAIL.n625 VTAIL.n591 6.59444
R817 VTAIL.n532 VTAIL.n495 6.59444
R818 VTAIL.n529 VTAIL.n495 6.59444
R819 VTAIL.n438 VTAIL.n401 6.59444
R820 VTAIL.n435 VTAIL.n401 6.59444
R821 VTAIL.n342 VTAIL.n305 6.59444
R822 VTAIL.n339 VTAIL.n305 6.59444
R823 VTAIL.n717 VTAIL.n686 5.81868
R824 VTAIL.n722 VTAIL.n682 5.81868
R825 VTAIL.n53 VTAIL.n22 5.81868
R826 VTAIL.n58 VTAIL.n18 5.81868
R827 VTAIL.n147 VTAIL.n116 5.81868
R828 VTAIL.n152 VTAIL.n112 5.81868
R829 VTAIL.n243 VTAIL.n212 5.81868
R830 VTAIL.n248 VTAIL.n208 5.81868
R831 VTAIL.n629 VTAIL.n589 5.81868
R832 VTAIL.n624 VTAIL.n593 5.81868
R833 VTAIL.n533 VTAIL.n493 5.81868
R834 VTAIL.n528 VTAIL.n497 5.81868
R835 VTAIL.n439 VTAIL.n399 5.81868
R836 VTAIL.n434 VTAIL.n403 5.81868
R837 VTAIL.n343 VTAIL.n303 5.81868
R838 VTAIL.n338 VTAIL.n307 5.81868
R839 VTAIL.n714 VTAIL.n713 5.04292
R840 VTAIL.n726 VTAIL.n725 5.04292
R841 VTAIL.n50 VTAIL.n49 5.04292
R842 VTAIL.n62 VTAIL.n61 5.04292
R843 VTAIL.n144 VTAIL.n143 5.04292
R844 VTAIL.n156 VTAIL.n155 5.04292
R845 VTAIL.n240 VTAIL.n239 5.04292
R846 VTAIL.n252 VTAIL.n251 5.04292
R847 VTAIL.n633 VTAIL.n632 5.04292
R848 VTAIL.n621 VTAIL.n620 5.04292
R849 VTAIL.n537 VTAIL.n536 5.04292
R850 VTAIL.n525 VTAIL.n524 5.04292
R851 VTAIL.n443 VTAIL.n442 5.04292
R852 VTAIL.n431 VTAIL.n430 5.04292
R853 VTAIL.n347 VTAIL.n346 5.04292
R854 VTAIL.n335 VTAIL.n334 5.04292
R855 VTAIL.n710 VTAIL.n688 4.26717
R856 VTAIL.n729 VTAIL.n680 4.26717
R857 VTAIL.n758 VTAIL.n666 4.26717
R858 VTAIL.n46 VTAIL.n24 4.26717
R859 VTAIL.n65 VTAIL.n16 4.26717
R860 VTAIL.n94 VTAIL.n2 4.26717
R861 VTAIL.n140 VTAIL.n118 4.26717
R862 VTAIL.n159 VTAIL.n110 4.26717
R863 VTAIL.n188 VTAIL.n96 4.26717
R864 VTAIL.n236 VTAIL.n214 4.26717
R865 VTAIL.n255 VTAIL.n206 4.26717
R866 VTAIL.n284 VTAIL.n192 4.26717
R867 VTAIL.n664 VTAIL.n572 4.26717
R868 VTAIL.n636 VTAIL.n587 4.26717
R869 VTAIL.n617 VTAIL.n595 4.26717
R870 VTAIL.n568 VTAIL.n476 4.26717
R871 VTAIL.n540 VTAIL.n491 4.26717
R872 VTAIL.n521 VTAIL.n499 4.26717
R873 VTAIL.n474 VTAIL.n382 4.26717
R874 VTAIL.n446 VTAIL.n397 4.26717
R875 VTAIL.n427 VTAIL.n405 4.26717
R876 VTAIL.n378 VTAIL.n286 4.26717
R877 VTAIL.n350 VTAIL.n301 4.26717
R878 VTAIL.n331 VTAIL.n309 4.26717
R879 VTAIL.n699 VTAIL.n695 3.70982
R880 VTAIL.n35 VTAIL.n31 3.70982
R881 VTAIL.n129 VTAIL.n125 3.70982
R882 VTAIL.n225 VTAIL.n221 3.70982
R883 VTAIL.n606 VTAIL.n602 3.70982
R884 VTAIL.n510 VTAIL.n506 3.70982
R885 VTAIL.n416 VTAIL.n412 3.70982
R886 VTAIL.n320 VTAIL.n316 3.70982
R887 VTAIL.n709 VTAIL.n690 3.49141
R888 VTAIL.n730 VTAIL.n678 3.49141
R889 VTAIL.n756 VTAIL.n755 3.49141
R890 VTAIL.n45 VTAIL.n26 3.49141
R891 VTAIL.n66 VTAIL.n14 3.49141
R892 VTAIL.n92 VTAIL.n91 3.49141
R893 VTAIL.n139 VTAIL.n120 3.49141
R894 VTAIL.n160 VTAIL.n108 3.49141
R895 VTAIL.n186 VTAIL.n185 3.49141
R896 VTAIL.n235 VTAIL.n216 3.49141
R897 VTAIL.n256 VTAIL.n204 3.49141
R898 VTAIL.n282 VTAIL.n281 3.49141
R899 VTAIL.n662 VTAIL.n661 3.49141
R900 VTAIL.n637 VTAIL.n585 3.49141
R901 VTAIL.n616 VTAIL.n597 3.49141
R902 VTAIL.n566 VTAIL.n565 3.49141
R903 VTAIL.n541 VTAIL.n489 3.49141
R904 VTAIL.n520 VTAIL.n501 3.49141
R905 VTAIL.n472 VTAIL.n471 3.49141
R906 VTAIL.n447 VTAIL.n395 3.49141
R907 VTAIL.n426 VTAIL.n407 3.49141
R908 VTAIL.n376 VTAIL.n375 3.49141
R909 VTAIL.n351 VTAIL.n299 3.49141
R910 VTAIL.n330 VTAIL.n311 3.49141
R911 VTAIL.n706 VTAIL.n705 2.71565
R912 VTAIL.n734 VTAIL.n733 2.71565
R913 VTAIL.n752 VTAIL.n668 2.71565
R914 VTAIL.n42 VTAIL.n41 2.71565
R915 VTAIL.n70 VTAIL.n69 2.71565
R916 VTAIL.n88 VTAIL.n4 2.71565
R917 VTAIL.n136 VTAIL.n135 2.71565
R918 VTAIL.n164 VTAIL.n163 2.71565
R919 VTAIL.n182 VTAIL.n98 2.71565
R920 VTAIL.n232 VTAIL.n231 2.71565
R921 VTAIL.n260 VTAIL.n259 2.71565
R922 VTAIL.n278 VTAIL.n194 2.71565
R923 VTAIL.n658 VTAIL.n574 2.71565
R924 VTAIL.n641 VTAIL.n640 2.71565
R925 VTAIL.n613 VTAIL.n612 2.71565
R926 VTAIL.n562 VTAIL.n478 2.71565
R927 VTAIL.n545 VTAIL.n544 2.71565
R928 VTAIL.n517 VTAIL.n516 2.71565
R929 VTAIL.n468 VTAIL.n384 2.71565
R930 VTAIL.n451 VTAIL.n450 2.71565
R931 VTAIL.n423 VTAIL.n422 2.71565
R932 VTAIL.n372 VTAIL.n288 2.71565
R933 VTAIL.n355 VTAIL.n354 2.71565
R934 VTAIL.n327 VTAIL.n326 2.71565
R935 VTAIL.n0 VTAIL.t2 1.94342
R936 VTAIL.n0 VTAIL.t3 1.94342
R937 VTAIL.n190 VTAIL.t14 1.94342
R938 VTAIL.n190 VTAIL.t15 1.94342
R939 VTAIL.n570 VTAIL.t12 1.94342
R940 VTAIL.n570 VTAIL.t11 1.94342
R941 VTAIL.n380 VTAIL.t4 1.94342
R942 VTAIL.n380 VTAIL.t6 1.94342
R943 VTAIL.n702 VTAIL.n692 1.93989
R944 VTAIL.n738 VTAIL.n676 1.93989
R945 VTAIL.n751 VTAIL.n670 1.93989
R946 VTAIL.n38 VTAIL.n28 1.93989
R947 VTAIL.n74 VTAIL.n12 1.93989
R948 VTAIL.n87 VTAIL.n6 1.93989
R949 VTAIL.n132 VTAIL.n122 1.93989
R950 VTAIL.n168 VTAIL.n106 1.93989
R951 VTAIL.n181 VTAIL.n100 1.93989
R952 VTAIL.n228 VTAIL.n218 1.93989
R953 VTAIL.n264 VTAIL.n202 1.93989
R954 VTAIL.n277 VTAIL.n196 1.93989
R955 VTAIL.n657 VTAIL.n576 1.93989
R956 VTAIL.n644 VTAIL.n582 1.93989
R957 VTAIL.n609 VTAIL.n599 1.93989
R958 VTAIL.n561 VTAIL.n480 1.93989
R959 VTAIL.n548 VTAIL.n486 1.93989
R960 VTAIL.n513 VTAIL.n503 1.93989
R961 VTAIL.n467 VTAIL.n386 1.93989
R962 VTAIL.n454 VTAIL.n392 1.93989
R963 VTAIL.n419 VTAIL.n409 1.93989
R964 VTAIL.n371 VTAIL.n290 1.93989
R965 VTAIL.n358 VTAIL.n296 1.93989
R966 VTAIL.n323 VTAIL.n313 1.93989
R967 VTAIL.n701 VTAIL.n694 1.16414
R968 VTAIL.n739 VTAIL.n674 1.16414
R969 VTAIL.n748 VTAIL.n747 1.16414
R970 VTAIL.n37 VTAIL.n30 1.16414
R971 VTAIL.n75 VTAIL.n10 1.16414
R972 VTAIL.n84 VTAIL.n83 1.16414
R973 VTAIL.n131 VTAIL.n124 1.16414
R974 VTAIL.n169 VTAIL.n104 1.16414
R975 VTAIL.n178 VTAIL.n177 1.16414
R976 VTAIL.n227 VTAIL.n220 1.16414
R977 VTAIL.n265 VTAIL.n200 1.16414
R978 VTAIL.n274 VTAIL.n273 1.16414
R979 VTAIL.n654 VTAIL.n653 1.16414
R980 VTAIL.n645 VTAIL.n580 1.16414
R981 VTAIL.n608 VTAIL.n601 1.16414
R982 VTAIL.n558 VTAIL.n557 1.16414
R983 VTAIL.n549 VTAIL.n484 1.16414
R984 VTAIL.n512 VTAIL.n505 1.16414
R985 VTAIL.n464 VTAIL.n463 1.16414
R986 VTAIL.n455 VTAIL.n390 1.16414
R987 VTAIL.n418 VTAIL.n411 1.16414
R988 VTAIL.n368 VTAIL.n367 1.16414
R989 VTAIL.n359 VTAIL.n294 1.16414
R990 VTAIL.n322 VTAIL.n315 1.16414
R991 VTAIL.n569 VTAIL.n475 0.470328
R992 VTAIL.n189 VTAIL.n95 0.470328
R993 VTAIL.n381 VTAIL.n379 0.440155
R994 VTAIL.n475 VTAIL.n381 0.440155
R995 VTAIL.n571 VTAIL.n569 0.440155
R996 VTAIL.n665 VTAIL.n571 0.440155
R997 VTAIL.n285 VTAIL.n191 0.440155
R998 VTAIL.n191 VTAIL.n189 0.440155
R999 VTAIL.n95 VTAIL.n1 0.440155
R1000 VTAIL.n698 VTAIL.n697 0.388379
R1001 VTAIL.n743 VTAIL.n742 0.388379
R1002 VTAIL.n744 VTAIL.n672 0.388379
R1003 VTAIL.n34 VTAIL.n33 0.388379
R1004 VTAIL.n79 VTAIL.n78 0.388379
R1005 VTAIL.n80 VTAIL.n8 0.388379
R1006 VTAIL.n128 VTAIL.n127 0.388379
R1007 VTAIL.n173 VTAIL.n172 0.388379
R1008 VTAIL.n174 VTAIL.n102 0.388379
R1009 VTAIL.n224 VTAIL.n223 0.388379
R1010 VTAIL.n269 VTAIL.n268 0.388379
R1011 VTAIL.n270 VTAIL.n198 0.388379
R1012 VTAIL.n650 VTAIL.n578 0.388379
R1013 VTAIL.n649 VTAIL.n648 0.388379
R1014 VTAIL.n605 VTAIL.n604 0.388379
R1015 VTAIL.n554 VTAIL.n482 0.388379
R1016 VTAIL.n553 VTAIL.n552 0.388379
R1017 VTAIL.n509 VTAIL.n508 0.388379
R1018 VTAIL.n460 VTAIL.n388 0.388379
R1019 VTAIL.n459 VTAIL.n458 0.388379
R1020 VTAIL.n415 VTAIL.n414 0.388379
R1021 VTAIL.n364 VTAIL.n292 0.388379
R1022 VTAIL.n363 VTAIL.n362 0.388379
R1023 VTAIL.n319 VTAIL.n318 0.388379
R1024 VTAIL VTAIL.n759 0.381966
R1025 VTAIL.n700 VTAIL.n699 0.155672
R1026 VTAIL.n700 VTAIL.n691 0.155672
R1027 VTAIL.n707 VTAIL.n691 0.155672
R1028 VTAIL.n708 VTAIL.n707 0.155672
R1029 VTAIL.n708 VTAIL.n687 0.155672
R1030 VTAIL.n715 VTAIL.n687 0.155672
R1031 VTAIL.n716 VTAIL.n715 0.155672
R1032 VTAIL.n716 VTAIL.n683 0.155672
R1033 VTAIL.n723 VTAIL.n683 0.155672
R1034 VTAIL.n724 VTAIL.n723 0.155672
R1035 VTAIL.n724 VTAIL.n679 0.155672
R1036 VTAIL.n731 VTAIL.n679 0.155672
R1037 VTAIL.n732 VTAIL.n731 0.155672
R1038 VTAIL.n732 VTAIL.n675 0.155672
R1039 VTAIL.n740 VTAIL.n675 0.155672
R1040 VTAIL.n741 VTAIL.n740 0.155672
R1041 VTAIL.n741 VTAIL.n671 0.155672
R1042 VTAIL.n749 VTAIL.n671 0.155672
R1043 VTAIL.n750 VTAIL.n749 0.155672
R1044 VTAIL.n750 VTAIL.n667 0.155672
R1045 VTAIL.n757 VTAIL.n667 0.155672
R1046 VTAIL.n36 VTAIL.n35 0.155672
R1047 VTAIL.n36 VTAIL.n27 0.155672
R1048 VTAIL.n43 VTAIL.n27 0.155672
R1049 VTAIL.n44 VTAIL.n43 0.155672
R1050 VTAIL.n44 VTAIL.n23 0.155672
R1051 VTAIL.n51 VTAIL.n23 0.155672
R1052 VTAIL.n52 VTAIL.n51 0.155672
R1053 VTAIL.n52 VTAIL.n19 0.155672
R1054 VTAIL.n59 VTAIL.n19 0.155672
R1055 VTAIL.n60 VTAIL.n59 0.155672
R1056 VTAIL.n60 VTAIL.n15 0.155672
R1057 VTAIL.n67 VTAIL.n15 0.155672
R1058 VTAIL.n68 VTAIL.n67 0.155672
R1059 VTAIL.n68 VTAIL.n11 0.155672
R1060 VTAIL.n76 VTAIL.n11 0.155672
R1061 VTAIL.n77 VTAIL.n76 0.155672
R1062 VTAIL.n77 VTAIL.n7 0.155672
R1063 VTAIL.n85 VTAIL.n7 0.155672
R1064 VTAIL.n86 VTAIL.n85 0.155672
R1065 VTAIL.n86 VTAIL.n3 0.155672
R1066 VTAIL.n93 VTAIL.n3 0.155672
R1067 VTAIL.n130 VTAIL.n129 0.155672
R1068 VTAIL.n130 VTAIL.n121 0.155672
R1069 VTAIL.n137 VTAIL.n121 0.155672
R1070 VTAIL.n138 VTAIL.n137 0.155672
R1071 VTAIL.n138 VTAIL.n117 0.155672
R1072 VTAIL.n145 VTAIL.n117 0.155672
R1073 VTAIL.n146 VTAIL.n145 0.155672
R1074 VTAIL.n146 VTAIL.n113 0.155672
R1075 VTAIL.n153 VTAIL.n113 0.155672
R1076 VTAIL.n154 VTAIL.n153 0.155672
R1077 VTAIL.n154 VTAIL.n109 0.155672
R1078 VTAIL.n161 VTAIL.n109 0.155672
R1079 VTAIL.n162 VTAIL.n161 0.155672
R1080 VTAIL.n162 VTAIL.n105 0.155672
R1081 VTAIL.n170 VTAIL.n105 0.155672
R1082 VTAIL.n171 VTAIL.n170 0.155672
R1083 VTAIL.n171 VTAIL.n101 0.155672
R1084 VTAIL.n179 VTAIL.n101 0.155672
R1085 VTAIL.n180 VTAIL.n179 0.155672
R1086 VTAIL.n180 VTAIL.n97 0.155672
R1087 VTAIL.n187 VTAIL.n97 0.155672
R1088 VTAIL.n226 VTAIL.n225 0.155672
R1089 VTAIL.n226 VTAIL.n217 0.155672
R1090 VTAIL.n233 VTAIL.n217 0.155672
R1091 VTAIL.n234 VTAIL.n233 0.155672
R1092 VTAIL.n234 VTAIL.n213 0.155672
R1093 VTAIL.n241 VTAIL.n213 0.155672
R1094 VTAIL.n242 VTAIL.n241 0.155672
R1095 VTAIL.n242 VTAIL.n209 0.155672
R1096 VTAIL.n249 VTAIL.n209 0.155672
R1097 VTAIL.n250 VTAIL.n249 0.155672
R1098 VTAIL.n250 VTAIL.n205 0.155672
R1099 VTAIL.n257 VTAIL.n205 0.155672
R1100 VTAIL.n258 VTAIL.n257 0.155672
R1101 VTAIL.n258 VTAIL.n201 0.155672
R1102 VTAIL.n266 VTAIL.n201 0.155672
R1103 VTAIL.n267 VTAIL.n266 0.155672
R1104 VTAIL.n267 VTAIL.n197 0.155672
R1105 VTAIL.n275 VTAIL.n197 0.155672
R1106 VTAIL.n276 VTAIL.n275 0.155672
R1107 VTAIL.n276 VTAIL.n193 0.155672
R1108 VTAIL.n283 VTAIL.n193 0.155672
R1109 VTAIL.n663 VTAIL.n573 0.155672
R1110 VTAIL.n656 VTAIL.n573 0.155672
R1111 VTAIL.n656 VTAIL.n655 0.155672
R1112 VTAIL.n655 VTAIL.n577 0.155672
R1113 VTAIL.n647 VTAIL.n577 0.155672
R1114 VTAIL.n647 VTAIL.n646 0.155672
R1115 VTAIL.n646 VTAIL.n581 0.155672
R1116 VTAIL.n639 VTAIL.n581 0.155672
R1117 VTAIL.n639 VTAIL.n638 0.155672
R1118 VTAIL.n638 VTAIL.n586 0.155672
R1119 VTAIL.n631 VTAIL.n586 0.155672
R1120 VTAIL.n631 VTAIL.n630 0.155672
R1121 VTAIL.n630 VTAIL.n590 0.155672
R1122 VTAIL.n623 VTAIL.n590 0.155672
R1123 VTAIL.n623 VTAIL.n622 0.155672
R1124 VTAIL.n622 VTAIL.n594 0.155672
R1125 VTAIL.n615 VTAIL.n594 0.155672
R1126 VTAIL.n615 VTAIL.n614 0.155672
R1127 VTAIL.n614 VTAIL.n598 0.155672
R1128 VTAIL.n607 VTAIL.n598 0.155672
R1129 VTAIL.n607 VTAIL.n606 0.155672
R1130 VTAIL.n567 VTAIL.n477 0.155672
R1131 VTAIL.n560 VTAIL.n477 0.155672
R1132 VTAIL.n560 VTAIL.n559 0.155672
R1133 VTAIL.n559 VTAIL.n481 0.155672
R1134 VTAIL.n551 VTAIL.n481 0.155672
R1135 VTAIL.n551 VTAIL.n550 0.155672
R1136 VTAIL.n550 VTAIL.n485 0.155672
R1137 VTAIL.n543 VTAIL.n485 0.155672
R1138 VTAIL.n543 VTAIL.n542 0.155672
R1139 VTAIL.n542 VTAIL.n490 0.155672
R1140 VTAIL.n535 VTAIL.n490 0.155672
R1141 VTAIL.n535 VTAIL.n534 0.155672
R1142 VTAIL.n534 VTAIL.n494 0.155672
R1143 VTAIL.n527 VTAIL.n494 0.155672
R1144 VTAIL.n527 VTAIL.n526 0.155672
R1145 VTAIL.n526 VTAIL.n498 0.155672
R1146 VTAIL.n519 VTAIL.n498 0.155672
R1147 VTAIL.n519 VTAIL.n518 0.155672
R1148 VTAIL.n518 VTAIL.n502 0.155672
R1149 VTAIL.n511 VTAIL.n502 0.155672
R1150 VTAIL.n511 VTAIL.n510 0.155672
R1151 VTAIL.n473 VTAIL.n383 0.155672
R1152 VTAIL.n466 VTAIL.n383 0.155672
R1153 VTAIL.n466 VTAIL.n465 0.155672
R1154 VTAIL.n465 VTAIL.n387 0.155672
R1155 VTAIL.n457 VTAIL.n387 0.155672
R1156 VTAIL.n457 VTAIL.n456 0.155672
R1157 VTAIL.n456 VTAIL.n391 0.155672
R1158 VTAIL.n449 VTAIL.n391 0.155672
R1159 VTAIL.n449 VTAIL.n448 0.155672
R1160 VTAIL.n448 VTAIL.n396 0.155672
R1161 VTAIL.n441 VTAIL.n396 0.155672
R1162 VTAIL.n441 VTAIL.n440 0.155672
R1163 VTAIL.n440 VTAIL.n400 0.155672
R1164 VTAIL.n433 VTAIL.n400 0.155672
R1165 VTAIL.n433 VTAIL.n432 0.155672
R1166 VTAIL.n432 VTAIL.n404 0.155672
R1167 VTAIL.n425 VTAIL.n404 0.155672
R1168 VTAIL.n425 VTAIL.n424 0.155672
R1169 VTAIL.n424 VTAIL.n408 0.155672
R1170 VTAIL.n417 VTAIL.n408 0.155672
R1171 VTAIL.n417 VTAIL.n416 0.155672
R1172 VTAIL.n377 VTAIL.n287 0.155672
R1173 VTAIL.n370 VTAIL.n287 0.155672
R1174 VTAIL.n370 VTAIL.n369 0.155672
R1175 VTAIL.n369 VTAIL.n291 0.155672
R1176 VTAIL.n361 VTAIL.n291 0.155672
R1177 VTAIL.n361 VTAIL.n360 0.155672
R1178 VTAIL.n360 VTAIL.n295 0.155672
R1179 VTAIL.n353 VTAIL.n295 0.155672
R1180 VTAIL.n353 VTAIL.n352 0.155672
R1181 VTAIL.n352 VTAIL.n300 0.155672
R1182 VTAIL.n345 VTAIL.n300 0.155672
R1183 VTAIL.n345 VTAIL.n344 0.155672
R1184 VTAIL.n344 VTAIL.n304 0.155672
R1185 VTAIL.n337 VTAIL.n304 0.155672
R1186 VTAIL.n337 VTAIL.n336 0.155672
R1187 VTAIL.n336 VTAIL.n308 0.155672
R1188 VTAIL.n329 VTAIL.n308 0.155672
R1189 VTAIL.n329 VTAIL.n328 0.155672
R1190 VTAIL.n328 VTAIL.n312 0.155672
R1191 VTAIL.n321 VTAIL.n312 0.155672
R1192 VTAIL.n321 VTAIL.n320 0.155672
R1193 VTAIL VTAIL.n1 0.0586897
R1194 B.n124 B.t6 2483.01
R1195 B.n278 B.t3 2483.01
R1196 B.n44 B.t0 2483.01
R1197 B.n38 B.t9 2483.01
R1198 B.n366 B.n365 585
R1199 B.n364 B.n91 585
R1200 B.n363 B.n362 585
R1201 B.n361 B.n92 585
R1202 B.n360 B.n359 585
R1203 B.n358 B.n93 585
R1204 B.n357 B.n356 585
R1205 B.n355 B.n94 585
R1206 B.n354 B.n353 585
R1207 B.n352 B.n95 585
R1208 B.n351 B.n350 585
R1209 B.n349 B.n96 585
R1210 B.n348 B.n347 585
R1211 B.n346 B.n97 585
R1212 B.n345 B.n344 585
R1213 B.n343 B.n98 585
R1214 B.n342 B.n341 585
R1215 B.n340 B.n99 585
R1216 B.n339 B.n338 585
R1217 B.n337 B.n100 585
R1218 B.n336 B.n335 585
R1219 B.n334 B.n101 585
R1220 B.n333 B.n332 585
R1221 B.n331 B.n102 585
R1222 B.n330 B.n329 585
R1223 B.n328 B.n103 585
R1224 B.n327 B.n326 585
R1225 B.n325 B.n104 585
R1226 B.n324 B.n323 585
R1227 B.n322 B.n105 585
R1228 B.n321 B.n320 585
R1229 B.n319 B.n106 585
R1230 B.n318 B.n317 585
R1231 B.n316 B.n107 585
R1232 B.n315 B.n314 585
R1233 B.n313 B.n108 585
R1234 B.n312 B.n311 585
R1235 B.n310 B.n109 585
R1236 B.n309 B.n308 585
R1237 B.n307 B.n110 585
R1238 B.n306 B.n305 585
R1239 B.n304 B.n111 585
R1240 B.n303 B.n302 585
R1241 B.n301 B.n112 585
R1242 B.n300 B.n299 585
R1243 B.n298 B.n113 585
R1244 B.n297 B.n296 585
R1245 B.n295 B.n114 585
R1246 B.n294 B.n293 585
R1247 B.n292 B.n115 585
R1248 B.n291 B.n290 585
R1249 B.n289 B.n116 585
R1250 B.n288 B.n287 585
R1251 B.n286 B.n117 585
R1252 B.n285 B.n284 585
R1253 B.n283 B.n118 585
R1254 B.n282 B.n281 585
R1255 B.n277 B.n119 585
R1256 B.n276 B.n275 585
R1257 B.n274 B.n120 585
R1258 B.n273 B.n272 585
R1259 B.n271 B.n121 585
R1260 B.n270 B.n269 585
R1261 B.n268 B.n122 585
R1262 B.n267 B.n266 585
R1263 B.n264 B.n123 585
R1264 B.n263 B.n262 585
R1265 B.n261 B.n126 585
R1266 B.n260 B.n259 585
R1267 B.n258 B.n127 585
R1268 B.n257 B.n256 585
R1269 B.n255 B.n128 585
R1270 B.n254 B.n253 585
R1271 B.n252 B.n129 585
R1272 B.n251 B.n250 585
R1273 B.n249 B.n130 585
R1274 B.n248 B.n247 585
R1275 B.n246 B.n131 585
R1276 B.n245 B.n244 585
R1277 B.n243 B.n132 585
R1278 B.n242 B.n241 585
R1279 B.n240 B.n133 585
R1280 B.n239 B.n238 585
R1281 B.n237 B.n134 585
R1282 B.n236 B.n235 585
R1283 B.n234 B.n135 585
R1284 B.n233 B.n232 585
R1285 B.n231 B.n136 585
R1286 B.n230 B.n229 585
R1287 B.n228 B.n137 585
R1288 B.n227 B.n226 585
R1289 B.n225 B.n138 585
R1290 B.n224 B.n223 585
R1291 B.n222 B.n139 585
R1292 B.n221 B.n220 585
R1293 B.n219 B.n140 585
R1294 B.n218 B.n217 585
R1295 B.n216 B.n141 585
R1296 B.n215 B.n214 585
R1297 B.n213 B.n142 585
R1298 B.n212 B.n211 585
R1299 B.n210 B.n143 585
R1300 B.n209 B.n208 585
R1301 B.n207 B.n144 585
R1302 B.n206 B.n205 585
R1303 B.n204 B.n145 585
R1304 B.n203 B.n202 585
R1305 B.n201 B.n146 585
R1306 B.n200 B.n199 585
R1307 B.n198 B.n147 585
R1308 B.n197 B.n196 585
R1309 B.n195 B.n148 585
R1310 B.n194 B.n193 585
R1311 B.n192 B.n149 585
R1312 B.n191 B.n190 585
R1313 B.n189 B.n150 585
R1314 B.n188 B.n187 585
R1315 B.n186 B.n151 585
R1316 B.n185 B.n184 585
R1317 B.n183 B.n152 585
R1318 B.n182 B.n181 585
R1319 B.n367 B.n90 585
R1320 B.n369 B.n368 585
R1321 B.n370 B.n89 585
R1322 B.n372 B.n371 585
R1323 B.n373 B.n88 585
R1324 B.n375 B.n374 585
R1325 B.n376 B.n87 585
R1326 B.n378 B.n377 585
R1327 B.n379 B.n86 585
R1328 B.n381 B.n380 585
R1329 B.n382 B.n85 585
R1330 B.n384 B.n383 585
R1331 B.n385 B.n84 585
R1332 B.n387 B.n386 585
R1333 B.n388 B.n83 585
R1334 B.n390 B.n389 585
R1335 B.n391 B.n82 585
R1336 B.n393 B.n392 585
R1337 B.n394 B.n81 585
R1338 B.n396 B.n395 585
R1339 B.n397 B.n80 585
R1340 B.n399 B.n398 585
R1341 B.n400 B.n79 585
R1342 B.n402 B.n401 585
R1343 B.n403 B.n78 585
R1344 B.n405 B.n404 585
R1345 B.n406 B.n77 585
R1346 B.n408 B.n407 585
R1347 B.n409 B.n76 585
R1348 B.n411 B.n410 585
R1349 B.n412 B.n75 585
R1350 B.n414 B.n413 585
R1351 B.n597 B.n596 585
R1352 B.n595 B.n10 585
R1353 B.n594 B.n593 585
R1354 B.n592 B.n11 585
R1355 B.n591 B.n590 585
R1356 B.n589 B.n12 585
R1357 B.n588 B.n587 585
R1358 B.n586 B.n13 585
R1359 B.n585 B.n584 585
R1360 B.n583 B.n14 585
R1361 B.n582 B.n581 585
R1362 B.n580 B.n15 585
R1363 B.n579 B.n578 585
R1364 B.n577 B.n16 585
R1365 B.n576 B.n575 585
R1366 B.n574 B.n17 585
R1367 B.n573 B.n572 585
R1368 B.n571 B.n18 585
R1369 B.n570 B.n569 585
R1370 B.n568 B.n19 585
R1371 B.n567 B.n566 585
R1372 B.n565 B.n20 585
R1373 B.n564 B.n563 585
R1374 B.n562 B.n21 585
R1375 B.n561 B.n560 585
R1376 B.n559 B.n22 585
R1377 B.n558 B.n557 585
R1378 B.n556 B.n23 585
R1379 B.n555 B.n554 585
R1380 B.n553 B.n24 585
R1381 B.n552 B.n551 585
R1382 B.n550 B.n25 585
R1383 B.n549 B.n548 585
R1384 B.n547 B.n26 585
R1385 B.n546 B.n545 585
R1386 B.n544 B.n27 585
R1387 B.n543 B.n542 585
R1388 B.n541 B.n28 585
R1389 B.n540 B.n539 585
R1390 B.n538 B.n29 585
R1391 B.n537 B.n536 585
R1392 B.n535 B.n30 585
R1393 B.n534 B.n533 585
R1394 B.n532 B.n31 585
R1395 B.n531 B.n530 585
R1396 B.n529 B.n32 585
R1397 B.n528 B.n527 585
R1398 B.n526 B.n33 585
R1399 B.n525 B.n524 585
R1400 B.n523 B.n34 585
R1401 B.n522 B.n521 585
R1402 B.n520 B.n35 585
R1403 B.n519 B.n518 585
R1404 B.n517 B.n36 585
R1405 B.n516 B.n515 585
R1406 B.n514 B.n37 585
R1407 B.n512 B.n511 585
R1408 B.n510 B.n40 585
R1409 B.n509 B.n508 585
R1410 B.n507 B.n41 585
R1411 B.n506 B.n505 585
R1412 B.n504 B.n42 585
R1413 B.n503 B.n502 585
R1414 B.n501 B.n43 585
R1415 B.n500 B.n499 585
R1416 B.n498 B.n497 585
R1417 B.n496 B.n47 585
R1418 B.n495 B.n494 585
R1419 B.n493 B.n48 585
R1420 B.n492 B.n491 585
R1421 B.n490 B.n49 585
R1422 B.n489 B.n488 585
R1423 B.n487 B.n50 585
R1424 B.n486 B.n485 585
R1425 B.n484 B.n51 585
R1426 B.n483 B.n482 585
R1427 B.n481 B.n52 585
R1428 B.n480 B.n479 585
R1429 B.n478 B.n53 585
R1430 B.n477 B.n476 585
R1431 B.n475 B.n54 585
R1432 B.n474 B.n473 585
R1433 B.n472 B.n55 585
R1434 B.n471 B.n470 585
R1435 B.n469 B.n56 585
R1436 B.n468 B.n467 585
R1437 B.n466 B.n57 585
R1438 B.n465 B.n464 585
R1439 B.n463 B.n58 585
R1440 B.n462 B.n461 585
R1441 B.n460 B.n59 585
R1442 B.n459 B.n458 585
R1443 B.n457 B.n60 585
R1444 B.n456 B.n455 585
R1445 B.n454 B.n61 585
R1446 B.n453 B.n452 585
R1447 B.n451 B.n62 585
R1448 B.n450 B.n449 585
R1449 B.n448 B.n63 585
R1450 B.n447 B.n446 585
R1451 B.n445 B.n64 585
R1452 B.n444 B.n443 585
R1453 B.n442 B.n65 585
R1454 B.n441 B.n440 585
R1455 B.n439 B.n66 585
R1456 B.n438 B.n437 585
R1457 B.n436 B.n67 585
R1458 B.n435 B.n434 585
R1459 B.n433 B.n68 585
R1460 B.n432 B.n431 585
R1461 B.n430 B.n69 585
R1462 B.n429 B.n428 585
R1463 B.n427 B.n70 585
R1464 B.n426 B.n425 585
R1465 B.n424 B.n71 585
R1466 B.n423 B.n422 585
R1467 B.n421 B.n72 585
R1468 B.n420 B.n419 585
R1469 B.n418 B.n73 585
R1470 B.n417 B.n416 585
R1471 B.n415 B.n74 585
R1472 B.n598 B.n9 585
R1473 B.n600 B.n599 585
R1474 B.n601 B.n8 585
R1475 B.n603 B.n602 585
R1476 B.n604 B.n7 585
R1477 B.n606 B.n605 585
R1478 B.n607 B.n6 585
R1479 B.n609 B.n608 585
R1480 B.n610 B.n5 585
R1481 B.n612 B.n611 585
R1482 B.n613 B.n4 585
R1483 B.n615 B.n614 585
R1484 B.n616 B.n3 585
R1485 B.n618 B.n617 585
R1486 B.n619 B.n0 585
R1487 B.n2 B.n1 585
R1488 B.n161 B.n160 585
R1489 B.n162 B.n159 585
R1490 B.n164 B.n163 585
R1491 B.n165 B.n158 585
R1492 B.n167 B.n166 585
R1493 B.n168 B.n157 585
R1494 B.n170 B.n169 585
R1495 B.n171 B.n156 585
R1496 B.n173 B.n172 585
R1497 B.n174 B.n155 585
R1498 B.n176 B.n175 585
R1499 B.n177 B.n154 585
R1500 B.n179 B.n178 585
R1501 B.n180 B.n153 585
R1502 B.n182 B.n153 487.695
R1503 B.n367 B.n366 487.695
R1504 B.n415 B.n414 487.695
R1505 B.n596 B.n9 487.695
R1506 B.n278 B.t4 470.575
R1507 B.n44 B.t2 470.575
R1508 B.n124 B.t7 470.574
R1509 B.n38 B.t11 470.574
R1510 B.n279 B.t5 460.683
R1511 B.n45 B.t1 460.683
R1512 B.n125 B.t8 460.683
R1513 B.n39 B.t10 460.683
R1514 B.n621 B.n620 256.663
R1515 B.n620 B.n619 235.042
R1516 B.n620 B.n2 235.042
R1517 B.n183 B.n182 163.367
R1518 B.n184 B.n183 163.367
R1519 B.n184 B.n151 163.367
R1520 B.n188 B.n151 163.367
R1521 B.n189 B.n188 163.367
R1522 B.n190 B.n189 163.367
R1523 B.n190 B.n149 163.367
R1524 B.n194 B.n149 163.367
R1525 B.n195 B.n194 163.367
R1526 B.n196 B.n195 163.367
R1527 B.n196 B.n147 163.367
R1528 B.n200 B.n147 163.367
R1529 B.n201 B.n200 163.367
R1530 B.n202 B.n201 163.367
R1531 B.n202 B.n145 163.367
R1532 B.n206 B.n145 163.367
R1533 B.n207 B.n206 163.367
R1534 B.n208 B.n207 163.367
R1535 B.n208 B.n143 163.367
R1536 B.n212 B.n143 163.367
R1537 B.n213 B.n212 163.367
R1538 B.n214 B.n213 163.367
R1539 B.n214 B.n141 163.367
R1540 B.n218 B.n141 163.367
R1541 B.n219 B.n218 163.367
R1542 B.n220 B.n219 163.367
R1543 B.n220 B.n139 163.367
R1544 B.n224 B.n139 163.367
R1545 B.n225 B.n224 163.367
R1546 B.n226 B.n225 163.367
R1547 B.n226 B.n137 163.367
R1548 B.n230 B.n137 163.367
R1549 B.n231 B.n230 163.367
R1550 B.n232 B.n231 163.367
R1551 B.n232 B.n135 163.367
R1552 B.n236 B.n135 163.367
R1553 B.n237 B.n236 163.367
R1554 B.n238 B.n237 163.367
R1555 B.n238 B.n133 163.367
R1556 B.n242 B.n133 163.367
R1557 B.n243 B.n242 163.367
R1558 B.n244 B.n243 163.367
R1559 B.n244 B.n131 163.367
R1560 B.n248 B.n131 163.367
R1561 B.n249 B.n248 163.367
R1562 B.n250 B.n249 163.367
R1563 B.n250 B.n129 163.367
R1564 B.n254 B.n129 163.367
R1565 B.n255 B.n254 163.367
R1566 B.n256 B.n255 163.367
R1567 B.n256 B.n127 163.367
R1568 B.n260 B.n127 163.367
R1569 B.n261 B.n260 163.367
R1570 B.n262 B.n261 163.367
R1571 B.n262 B.n123 163.367
R1572 B.n267 B.n123 163.367
R1573 B.n268 B.n267 163.367
R1574 B.n269 B.n268 163.367
R1575 B.n269 B.n121 163.367
R1576 B.n273 B.n121 163.367
R1577 B.n274 B.n273 163.367
R1578 B.n275 B.n274 163.367
R1579 B.n275 B.n119 163.367
R1580 B.n282 B.n119 163.367
R1581 B.n283 B.n282 163.367
R1582 B.n284 B.n283 163.367
R1583 B.n284 B.n117 163.367
R1584 B.n288 B.n117 163.367
R1585 B.n289 B.n288 163.367
R1586 B.n290 B.n289 163.367
R1587 B.n290 B.n115 163.367
R1588 B.n294 B.n115 163.367
R1589 B.n295 B.n294 163.367
R1590 B.n296 B.n295 163.367
R1591 B.n296 B.n113 163.367
R1592 B.n300 B.n113 163.367
R1593 B.n301 B.n300 163.367
R1594 B.n302 B.n301 163.367
R1595 B.n302 B.n111 163.367
R1596 B.n306 B.n111 163.367
R1597 B.n307 B.n306 163.367
R1598 B.n308 B.n307 163.367
R1599 B.n308 B.n109 163.367
R1600 B.n312 B.n109 163.367
R1601 B.n313 B.n312 163.367
R1602 B.n314 B.n313 163.367
R1603 B.n314 B.n107 163.367
R1604 B.n318 B.n107 163.367
R1605 B.n319 B.n318 163.367
R1606 B.n320 B.n319 163.367
R1607 B.n320 B.n105 163.367
R1608 B.n324 B.n105 163.367
R1609 B.n325 B.n324 163.367
R1610 B.n326 B.n325 163.367
R1611 B.n326 B.n103 163.367
R1612 B.n330 B.n103 163.367
R1613 B.n331 B.n330 163.367
R1614 B.n332 B.n331 163.367
R1615 B.n332 B.n101 163.367
R1616 B.n336 B.n101 163.367
R1617 B.n337 B.n336 163.367
R1618 B.n338 B.n337 163.367
R1619 B.n338 B.n99 163.367
R1620 B.n342 B.n99 163.367
R1621 B.n343 B.n342 163.367
R1622 B.n344 B.n343 163.367
R1623 B.n344 B.n97 163.367
R1624 B.n348 B.n97 163.367
R1625 B.n349 B.n348 163.367
R1626 B.n350 B.n349 163.367
R1627 B.n350 B.n95 163.367
R1628 B.n354 B.n95 163.367
R1629 B.n355 B.n354 163.367
R1630 B.n356 B.n355 163.367
R1631 B.n356 B.n93 163.367
R1632 B.n360 B.n93 163.367
R1633 B.n361 B.n360 163.367
R1634 B.n362 B.n361 163.367
R1635 B.n362 B.n91 163.367
R1636 B.n366 B.n91 163.367
R1637 B.n414 B.n75 163.367
R1638 B.n410 B.n75 163.367
R1639 B.n410 B.n409 163.367
R1640 B.n409 B.n408 163.367
R1641 B.n408 B.n77 163.367
R1642 B.n404 B.n77 163.367
R1643 B.n404 B.n403 163.367
R1644 B.n403 B.n402 163.367
R1645 B.n402 B.n79 163.367
R1646 B.n398 B.n79 163.367
R1647 B.n398 B.n397 163.367
R1648 B.n397 B.n396 163.367
R1649 B.n396 B.n81 163.367
R1650 B.n392 B.n81 163.367
R1651 B.n392 B.n391 163.367
R1652 B.n391 B.n390 163.367
R1653 B.n390 B.n83 163.367
R1654 B.n386 B.n83 163.367
R1655 B.n386 B.n385 163.367
R1656 B.n385 B.n384 163.367
R1657 B.n384 B.n85 163.367
R1658 B.n380 B.n85 163.367
R1659 B.n380 B.n379 163.367
R1660 B.n379 B.n378 163.367
R1661 B.n378 B.n87 163.367
R1662 B.n374 B.n87 163.367
R1663 B.n374 B.n373 163.367
R1664 B.n373 B.n372 163.367
R1665 B.n372 B.n89 163.367
R1666 B.n368 B.n89 163.367
R1667 B.n368 B.n367 163.367
R1668 B.n596 B.n595 163.367
R1669 B.n595 B.n594 163.367
R1670 B.n594 B.n11 163.367
R1671 B.n590 B.n11 163.367
R1672 B.n590 B.n589 163.367
R1673 B.n589 B.n588 163.367
R1674 B.n588 B.n13 163.367
R1675 B.n584 B.n13 163.367
R1676 B.n584 B.n583 163.367
R1677 B.n583 B.n582 163.367
R1678 B.n582 B.n15 163.367
R1679 B.n578 B.n15 163.367
R1680 B.n578 B.n577 163.367
R1681 B.n577 B.n576 163.367
R1682 B.n576 B.n17 163.367
R1683 B.n572 B.n17 163.367
R1684 B.n572 B.n571 163.367
R1685 B.n571 B.n570 163.367
R1686 B.n570 B.n19 163.367
R1687 B.n566 B.n19 163.367
R1688 B.n566 B.n565 163.367
R1689 B.n565 B.n564 163.367
R1690 B.n564 B.n21 163.367
R1691 B.n560 B.n21 163.367
R1692 B.n560 B.n559 163.367
R1693 B.n559 B.n558 163.367
R1694 B.n558 B.n23 163.367
R1695 B.n554 B.n23 163.367
R1696 B.n554 B.n553 163.367
R1697 B.n553 B.n552 163.367
R1698 B.n552 B.n25 163.367
R1699 B.n548 B.n25 163.367
R1700 B.n548 B.n547 163.367
R1701 B.n547 B.n546 163.367
R1702 B.n546 B.n27 163.367
R1703 B.n542 B.n27 163.367
R1704 B.n542 B.n541 163.367
R1705 B.n541 B.n540 163.367
R1706 B.n540 B.n29 163.367
R1707 B.n536 B.n29 163.367
R1708 B.n536 B.n535 163.367
R1709 B.n535 B.n534 163.367
R1710 B.n534 B.n31 163.367
R1711 B.n530 B.n31 163.367
R1712 B.n530 B.n529 163.367
R1713 B.n529 B.n528 163.367
R1714 B.n528 B.n33 163.367
R1715 B.n524 B.n33 163.367
R1716 B.n524 B.n523 163.367
R1717 B.n523 B.n522 163.367
R1718 B.n522 B.n35 163.367
R1719 B.n518 B.n35 163.367
R1720 B.n518 B.n517 163.367
R1721 B.n517 B.n516 163.367
R1722 B.n516 B.n37 163.367
R1723 B.n511 B.n37 163.367
R1724 B.n511 B.n510 163.367
R1725 B.n510 B.n509 163.367
R1726 B.n509 B.n41 163.367
R1727 B.n505 B.n41 163.367
R1728 B.n505 B.n504 163.367
R1729 B.n504 B.n503 163.367
R1730 B.n503 B.n43 163.367
R1731 B.n499 B.n43 163.367
R1732 B.n499 B.n498 163.367
R1733 B.n498 B.n47 163.367
R1734 B.n494 B.n47 163.367
R1735 B.n494 B.n493 163.367
R1736 B.n493 B.n492 163.367
R1737 B.n492 B.n49 163.367
R1738 B.n488 B.n49 163.367
R1739 B.n488 B.n487 163.367
R1740 B.n487 B.n486 163.367
R1741 B.n486 B.n51 163.367
R1742 B.n482 B.n51 163.367
R1743 B.n482 B.n481 163.367
R1744 B.n481 B.n480 163.367
R1745 B.n480 B.n53 163.367
R1746 B.n476 B.n53 163.367
R1747 B.n476 B.n475 163.367
R1748 B.n475 B.n474 163.367
R1749 B.n474 B.n55 163.367
R1750 B.n470 B.n55 163.367
R1751 B.n470 B.n469 163.367
R1752 B.n469 B.n468 163.367
R1753 B.n468 B.n57 163.367
R1754 B.n464 B.n57 163.367
R1755 B.n464 B.n463 163.367
R1756 B.n463 B.n462 163.367
R1757 B.n462 B.n59 163.367
R1758 B.n458 B.n59 163.367
R1759 B.n458 B.n457 163.367
R1760 B.n457 B.n456 163.367
R1761 B.n456 B.n61 163.367
R1762 B.n452 B.n61 163.367
R1763 B.n452 B.n451 163.367
R1764 B.n451 B.n450 163.367
R1765 B.n450 B.n63 163.367
R1766 B.n446 B.n63 163.367
R1767 B.n446 B.n445 163.367
R1768 B.n445 B.n444 163.367
R1769 B.n444 B.n65 163.367
R1770 B.n440 B.n65 163.367
R1771 B.n440 B.n439 163.367
R1772 B.n439 B.n438 163.367
R1773 B.n438 B.n67 163.367
R1774 B.n434 B.n67 163.367
R1775 B.n434 B.n433 163.367
R1776 B.n433 B.n432 163.367
R1777 B.n432 B.n69 163.367
R1778 B.n428 B.n69 163.367
R1779 B.n428 B.n427 163.367
R1780 B.n427 B.n426 163.367
R1781 B.n426 B.n71 163.367
R1782 B.n422 B.n71 163.367
R1783 B.n422 B.n421 163.367
R1784 B.n421 B.n420 163.367
R1785 B.n420 B.n73 163.367
R1786 B.n416 B.n73 163.367
R1787 B.n416 B.n415 163.367
R1788 B.n600 B.n9 163.367
R1789 B.n601 B.n600 163.367
R1790 B.n602 B.n601 163.367
R1791 B.n602 B.n7 163.367
R1792 B.n606 B.n7 163.367
R1793 B.n607 B.n606 163.367
R1794 B.n608 B.n607 163.367
R1795 B.n608 B.n5 163.367
R1796 B.n612 B.n5 163.367
R1797 B.n613 B.n612 163.367
R1798 B.n614 B.n613 163.367
R1799 B.n614 B.n3 163.367
R1800 B.n618 B.n3 163.367
R1801 B.n619 B.n618 163.367
R1802 B.n160 B.n2 163.367
R1803 B.n160 B.n159 163.367
R1804 B.n164 B.n159 163.367
R1805 B.n165 B.n164 163.367
R1806 B.n166 B.n165 163.367
R1807 B.n166 B.n157 163.367
R1808 B.n170 B.n157 163.367
R1809 B.n171 B.n170 163.367
R1810 B.n172 B.n171 163.367
R1811 B.n172 B.n155 163.367
R1812 B.n176 B.n155 163.367
R1813 B.n177 B.n176 163.367
R1814 B.n178 B.n177 163.367
R1815 B.n178 B.n153 163.367
R1816 B.n265 B.n125 59.5399
R1817 B.n280 B.n279 59.5399
R1818 B.n46 B.n45 59.5399
R1819 B.n513 B.n39 59.5399
R1820 B.n598 B.n597 31.6883
R1821 B.n413 B.n74 31.6883
R1822 B.n365 B.n90 31.6883
R1823 B.n181 B.n180 31.6883
R1824 B B.n621 18.0485
R1825 B.n599 B.n598 10.6151
R1826 B.n599 B.n8 10.6151
R1827 B.n603 B.n8 10.6151
R1828 B.n604 B.n603 10.6151
R1829 B.n605 B.n604 10.6151
R1830 B.n605 B.n6 10.6151
R1831 B.n609 B.n6 10.6151
R1832 B.n610 B.n609 10.6151
R1833 B.n611 B.n610 10.6151
R1834 B.n611 B.n4 10.6151
R1835 B.n615 B.n4 10.6151
R1836 B.n616 B.n615 10.6151
R1837 B.n617 B.n616 10.6151
R1838 B.n617 B.n0 10.6151
R1839 B.n597 B.n10 10.6151
R1840 B.n593 B.n10 10.6151
R1841 B.n593 B.n592 10.6151
R1842 B.n592 B.n591 10.6151
R1843 B.n591 B.n12 10.6151
R1844 B.n587 B.n12 10.6151
R1845 B.n587 B.n586 10.6151
R1846 B.n586 B.n585 10.6151
R1847 B.n585 B.n14 10.6151
R1848 B.n581 B.n14 10.6151
R1849 B.n581 B.n580 10.6151
R1850 B.n580 B.n579 10.6151
R1851 B.n579 B.n16 10.6151
R1852 B.n575 B.n16 10.6151
R1853 B.n575 B.n574 10.6151
R1854 B.n574 B.n573 10.6151
R1855 B.n573 B.n18 10.6151
R1856 B.n569 B.n18 10.6151
R1857 B.n569 B.n568 10.6151
R1858 B.n568 B.n567 10.6151
R1859 B.n567 B.n20 10.6151
R1860 B.n563 B.n20 10.6151
R1861 B.n563 B.n562 10.6151
R1862 B.n562 B.n561 10.6151
R1863 B.n561 B.n22 10.6151
R1864 B.n557 B.n22 10.6151
R1865 B.n557 B.n556 10.6151
R1866 B.n556 B.n555 10.6151
R1867 B.n555 B.n24 10.6151
R1868 B.n551 B.n24 10.6151
R1869 B.n551 B.n550 10.6151
R1870 B.n550 B.n549 10.6151
R1871 B.n549 B.n26 10.6151
R1872 B.n545 B.n26 10.6151
R1873 B.n545 B.n544 10.6151
R1874 B.n544 B.n543 10.6151
R1875 B.n543 B.n28 10.6151
R1876 B.n539 B.n28 10.6151
R1877 B.n539 B.n538 10.6151
R1878 B.n538 B.n537 10.6151
R1879 B.n537 B.n30 10.6151
R1880 B.n533 B.n30 10.6151
R1881 B.n533 B.n532 10.6151
R1882 B.n532 B.n531 10.6151
R1883 B.n531 B.n32 10.6151
R1884 B.n527 B.n32 10.6151
R1885 B.n527 B.n526 10.6151
R1886 B.n526 B.n525 10.6151
R1887 B.n525 B.n34 10.6151
R1888 B.n521 B.n34 10.6151
R1889 B.n521 B.n520 10.6151
R1890 B.n520 B.n519 10.6151
R1891 B.n519 B.n36 10.6151
R1892 B.n515 B.n36 10.6151
R1893 B.n515 B.n514 10.6151
R1894 B.n512 B.n40 10.6151
R1895 B.n508 B.n40 10.6151
R1896 B.n508 B.n507 10.6151
R1897 B.n507 B.n506 10.6151
R1898 B.n506 B.n42 10.6151
R1899 B.n502 B.n42 10.6151
R1900 B.n502 B.n501 10.6151
R1901 B.n501 B.n500 10.6151
R1902 B.n497 B.n496 10.6151
R1903 B.n496 B.n495 10.6151
R1904 B.n495 B.n48 10.6151
R1905 B.n491 B.n48 10.6151
R1906 B.n491 B.n490 10.6151
R1907 B.n490 B.n489 10.6151
R1908 B.n489 B.n50 10.6151
R1909 B.n485 B.n50 10.6151
R1910 B.n485 B.n484 10.6151
R1911 B.n484 B.n483 10.6151
R1912 B.n483 B.n52 10.6151
R1913 B.n479 B.n52 10.6151
R1914 B.n479 B.n478 10.6151
R1915 B.n478 B.n477 10.6151
R1916 B.n477 B.n54 10.6151
R1917 B.n473 B.n54 10.6151
R1918 B.n473 B.n472 10.6151
R1919 B.n472 B.n471 10.6151
R1920 B.n471 B.n56 10.6151
R1921 B.n467 B.n56 10.6151
R1922 B.n467 B.n466 10.6151
R1923 B.n466 B.n465 10.6151
R1924 B.n465 B.n58 10.6151
R1925 B.n461 B.n58 10.6151
R1926 B.n461 B.n460 10.6151
R1927 B.n460 B.n459 10.6151
R1928 B.n459 B.n60 10.6151
R1929 B.n455 B.n60 10.6151
R1930 B.n455 B.n454 10.6151
R1931 B.n454 B.n453 10.6151
R1932 B.n453 B.n62 10.6151
R1933 B.n449 B.n62 10.6151
R1934 B.n449 B.n448 10.6151
R1935 B.n448 B.n447 10.6151
R1936 B.n447 B.n64 10.6151
R1937 B.n443 B.n64 10.6151
R1938 B.n443 B.n442 10.6151
R1939 B.n442 B.n441 10.6151
R1940 B.n441 B.n66 10.6151
R1941 B.n437 B.n66 10.6151
R1942 B.n437 B.n436 10.6151
R1943 B.n436 B.n435 10.6151
R1944 B.n435 B.n68 10.6151
R1945 B.n431 B.n68 10.6151
R1946 B.n431 B.n430 10.6151
R1947 B.n430 B.n429 10.6151
R1948 B.n429 B.n70 10.6151
R1949 B.n425 B.n70 10.6151
R1950 B.n425 B.n424 10.6151
R1951 B.n424 B.n423 10.6151
R1952 B.n423 B.n72 10.6151
R1953 B.n419 B.n72 10.6151
R1954 B.n419 B.n418 10.6151
R1955 B.n418 B.n417 10.6151
R1956 B.n417 B.n74 10.6151
R1957 B.n413 B.n412 10.6151
R1958 B.n412 B.n411 10.6151
R1959 B.n411 B.n76 10.6151
R1960 B.n407 B.n76 10.6151
R1961 B.n407 B.n406 10.6151
R1962 B.n406 B.n405 10.6151
R1963 B.n405 B.n78 10.6151
R1964 B.n401 B.n78 10.6151
R1965 B.n401 B.n400 10.6151
R1966 B.n400 B.n399 10.6151
R1967 B.n399 B.n80 10.6151
R1968 B.n395 B.n80 10.6151
R1969 B.n395 B.n394 10.6151
R1970 B.n394 B.n393 10.6151
R1971 B.n393 B.n82 10.6151
R1972 B.n389 B.n82 10.6151
R1973 B.n389 B.n388 10.6151
R1974 B.n388 B.n387 10.6151
R1975 B.n387 B.n84 10.6151
R1976 B.n383 B.n84 10.6151
R1977 B.n383 B.n382 10.6151
R1978 B.n382 B.n381 10.6151
R1979 B.n381 B.n86 10.6151
R1980 B.n377 B.n86 10.6151
R1981 B.n377 B.n376 10.6151
R1982 B.n376 B.n375 10.6151
R1983 B.n375 B.n88 10.6151
R1984 B.n371 B.n88 10.6151
R1985 B.n371 B.n370 10.6151
R1986 B.n370 B.n369 10.6151
R1987 B.n369 B.n90 10.6151
R1988 B.n161 B.n1 10.6151
R1989 B.n162 B.n161 10.6151
R1990 B.n163 B.n162 10.6151
R1991 B.n163 B.n158 10.6151
R1992 B.n167 B.n158 10.6151
R1993 B.n168 B.n167 10.6151
R1994 B.n169 B.n168 10.6151
R1995 B.n169 B.n156 10.6151
R1996 B.n173 B.n156 10.6151
R1997 B.n174 B.n173 10.6151
R1998 B.n175 B.n174 10.6151
R1999 B.n175 B.n154 10.6151
R2000 B.n179 B.n154 10.6151
R2001 B.n180 B.n179 10.6151
R2002 B.n181 B.n152 10.6151
R2003 B.n185 B.n152 10.6151
R2004 B.n186 B.n185 10.6151
R2005 B.n187 B.n186 10.6151
R2006 B.n187 B.n150 10.6151
R2007 B.n191 B.n150 10.6151
R2008 B.n192 B.n191 10.6151
R2009 B.n193 B.n192 10.6151
R2010 B.n193 B.n148 10.6151
R2011 B.n197 B.n148 10.6151
R2012 B.n198 B.n197 10.6151
R2013 B.n199 B.n198 10.6151
R2014 B.n199 B.n146 10.6151
R2015 B.n203 B.n146 10.6151
R2016 B.n204 B.n203 10.6151
R2017 B.n205 B.n204 10.6151
R2018 B.n205 B.n144 10.6151
R2019 B.n209 B.n144 10.6151
R2020 B.n210 B.n209 10.6151
R2021 B.n211 B.n210 10.6151
R2022 B.n211 B.n142 10.6151
R2023 B.n215 B.n142 10.6151
R2024 B.n216 B.n215 10.6151
R2025 B.n217 B.n216 10.6151
R2026 B.n217 B.n140 10.6151
R2027 B.n221 B.n140 10.6151
R2028 B.n222 B.n221 10.6151
R2029 B.n223 B.n222 10.6151
R2030 B.n223 B.n138 10.6151
R2031 B.n227 B.n138 10.6151
R2032 B.n228 B.n227 10.6151
R2033 B.n229 B.n228 10.6151
R2034 B.n229 B.n136 10.6151
R2035 B.n233 B.n136 10.6151
R2036 B.n234 B.n233 10.6151
R2037 B.n235 B.n234 10.6151
R2038 B.n235 B.n134 10.6151
R2039 B.n239 B.n134 10.6151
R2040 B.n240 B.n239 10.6151
R2041 B.n241 B.n240 10.6151
R2042 B.n241 B.n132 10.6151
R2043 B.n245 B.n132 10.6151
R2044 B.n246 B.n245 10.6151
R2045 B.n247 B.n246 10.6151
R2046 B.n247 B.n130 10.6151
R2047 B.n251 B.n130 10.6151
R2048 B.n252 B.n251 10.6151
R2049 B.n253 B.n252 10.6151
R2050 B.n253 B.n128 10.6151
R2051 B.n257 B.n128 10.6151
R2052 B.n258 B.n257 10.6151
R2053 B.n259 B.n258 10.6151
R2054 B.n259 B.n126 10.6151
R2055 B.n263 B.n126 10.6151
R2056 B.n264 B.n263 10.6151
R2057 B.n266 B.n122 10.6151
R2058 B.n270 B.n122 10.6151
R2059 B.n271 B.n270 10.6151
R2060 B.n272 B.n271 10.6151
R2061 B.n272 B.n120 10.6151
R2062 B.n276 B.n120 10.6151
R2063 B.n277 B.n276 10.6151
R2064 B.n281 B.n277 10.6151
R2065 B.n285 B.n118 10.6151
R2066 B.n286 B.n285 10.6151
R2067 B.n287 B.n286 10.6151
R2068 B.n287 B.n116 10.6151
R2069 B.n291 B.n116 10.6151
R2070 B.n292 B.n291 10.6151
R2071 B.n293 B.n292 10.6151
R2072 B.n293 B.n114 10.6151
R2073 B.n297 B.n114 10.6151
R2074 B.n298 B.n297 10.6151
R2075 B.n299 B.n298 10.6151
R2076 B.n299 B.n112 10.6151
R2077 B.n303 B.n112 10.6151
R2078 B.n304 B.n303 10.6151
R2079 B.n305 B.n304 10.6151
R2080 B.n305 B.n110 10.6151
R2081 B.n309 B.n110 10.6151
R2082 B.n310 B.n309 10.6151
R2083 B.n311 B.n310 10.6151
R2084 B.n311 B.n108 10.6151
R2085 B.n315 B.n108 10.6151
R2086 B.n316 B.n315 10.6151
R2087 B.n317 B.n316 10.6151
R2088 B.n317 B.n106 10.6151
R2089 B.n321 B.n106 10.6151
R2090 B.n322 B.n321 10.6151
R2091 B.n323 B.n322 10.6151
R2092 B.n323 B.n104 10.6151
R2093 B.n327 B.n104 10.6151
R2094 B.n328 B.n327 10.6151
R2095 B.n329 B.n328 10.6151
R2096 B.n329 B.n102 10.6151
R2097 B.n333 B.n102 10.6151
R2098 B.n334 B.n333 10.6151
R2099 B.n335 B.n334 10.6151
R2100 B.n335 B.n100 10.6151
R2101 B.n339 B.n100 10.6151
R2102 B.n340 B.n339 10.6151
R2103 B.n341 B.n340 10.6151
R2104 B.n341 B.n98 10.6151
R2105 B.n345 B.n98 10.6151
R2106 B.n346 B.n345 10.6151
R2107 B.n347 B.n346 10.6151
R2108 B.n347 B.n96 10.6151
R2109 B.n351 B.n96 10.6151
R2110 B.n352 B.n351 10.6151
R2111 B.n353 B.n352 10.6151
R2112 B.n353 B.n94 10.6151
R2113 B.n357 B.n94 10.6151
R2114 B.n358 B.n357 10.6151
R2115 B.n359 B.n358 10.6151
R2116 B.n359 B.n92 10.6151
R2117 B.n363 B.n92 10.6151
R2118 B.n364 B.n363 10.6151
R2119 B.n365 B.n364 10.6151
R2120 B.n125 B.n124 9.89141
R2121 B.n279 B.n278 9.89141
R2122 B.n45 B.n44 9.89141
R2123 B.n39 B.n38 9.89141
R2124 B.n621 B.n0 8.11757
R2125 B.n621 B.n1 8.11757
R2126 B.n513 B.n512 6.5566
R2127 B.n500 B.n46 6.5566
R2128 B.n266 B.n265 6.5566
R2129 B.n281 B.n280 6.5566
R2130 B.n514 B.n513 4.05904
R2131 B.n497 B.n46 4.05904
R2132 B.n265 B.n264 4.05904
R2133 B.n280 B.n118 4.05904
R2134 VN.n5 VN.t0 2454.06
R2135 VN.n1 VN.t4 2454.06
R2136 VN.n12 VN.t5 2454.06
R2137 VN.n8 VN.t1 2454.06
R2138 VN.n4 VN.t7 2415.36
R2139 VN.n2 VN.t6 2415.36
R2140 VN.n11 VN.t3 2415.36
R2141 VN.n9 VN.t2 2415.36
R2142 VN.n8 VN.n7 161.489
R2143 VN.n1 VN.n0 161.489
R2144 VN.n6 VN.n5 161.3
R2145 VN.n13 VN.n12 161.3
R2146 VN.n10 VN.n7 161.3
R2147 VN.n3 VN.n0 161.3
R2148 VN VN.n13 43.563
R2149 VN.n3 VN.n2 37.246
R2150 VN.n4 VN.n3 37.246
R2151 VN.n11 VN.n10 37.246
R2152 VN.n10 VN.n9 37.246
R2153 VN.n2 VN.n1 35.7853
R2154 VN.n5 VN.n4 35.7853
R2155 VN.n12 VN.n11 35.7853
R2156 VN.n9 VN.n8 35.7853
R2157 VN.n13 VN.n7 0.189894
R2158 VN.n6 VN.n0 0.189894
R2159 VN VN.n6 0.0516364
R2160 VDD2.n2 VDD2.n1 68.1987
R2161 VDD2.n2 VDD2.n0 68.1987
R2162 VDD2 VDD2.n5 68.1959
R2163 VDD2.n4 VDD2.n3 68.0345
R2164 VDD2.n4 VDD2.n2 40.1162
R2165 VDD2.n5 VDD2.t5 1.94342
R2166 VDD2.n5 VDD2.t6 1.94342
R2167 VDD2.n3 VDD2.t2 1.94342
R2168 VDD2.n3 VDD2.t4 1.94342
R2169 VDD2.n1 VDD2.t0 1.94342
R2170 VDD2.n1 VDD2.t7 1.94342
R2171 VDD2.n0 VDD2.t3 1.94342
R2172 VDD2.n0 VDD2.t1 1.94342
R2173 VDD2 VDD2.n4 0.278517
C0 VP w_n1480_n4314# 2.62145f
C1 VDD1 VDD2 0.572911f
C2 VN VTAIL 2.56607f
C3 B VDD2 1.05957f
C4 VTAIL VDD1 27.664598f
C5 B VTAIL 4.52358f
C6 VTAIL VDD2 27.7028f
C7 VN w_n1480_n4314# 2.43645f
C8 VDD1 w_n1480_n4314# 1.20118f
C9 B w_n1480_n4314# 7.80689f
C10 VDD2 w_n1480_n4314# 1.21501f
C11 VTAIL w_n1480_n4314# 5.58016f
C12 VP VN 5.581f
C13 VP VDD1 3.40191f
C14 B VP 1.0092f
C15 VP VDD2 0.261618f
C16 VP VTAIL 2.58018f
C17 VN VDD1 0.146814f
C18 B VN 0.711973f
C19 B VDD1 1.03841f
C20 VN VDD2 3.28728f
C21 VDD2 VSUBS 1.619883f
C22 VDD1 VSUBS 1.821097f
C23 VTAIL VSUBS 0.752624f
C24 VN VSUBS 5.08069f
C25 VP VSUBS 1.295766f
C26 B VSUBS 2.692472f
C27 w_n1480_n4314# VSUBS 78.1618f
C28 VDD2.t3 VSUBS 0.523008f
C29 VDD2.t1 VSUBS 0.523008f
C30 VDD2.n0 VSUBS 4.29677f
C31 VDD2.t0 VSUBS 0.523008f
C32 VDD2.t7 VSUBS 0.523008f
C33 VDD2.n1 VSUBS 4.29677f
C34 VDD2.n2 VSUBS 4.32817f
C35 VDD2.t2 VSUBS 0.523008f
C36 VDD2.t4 VSUBS 0.523008f
C37 VDD2.n3 VSUBS 4.294661f
C38 VDD2.n4 VSUBS 4.37378f
C39 VDD2.t5 VSUBS 0.523008f
C40 VDD2.t6 VSUBS 0.523008f
C41 VDD2.n5 VSUBS 4.296721f
C42 VN.n0 VSUBS 0.156118f
C43 VN.t7 VSUBS 0.622923f
C44 VN.t6 VSUBS 0.622923f
C45 VN.t4 VSUBS 0.62675f
C46 VN.n1 VSUBS 0.26371f
C47 VN.n2 VSUBS 0.24514f
C48 VN.n3 VSUBS 0.024788f
C49 VN.n4 VSUBS 0.24514f
C50 VN.t0 VSUBS 0.62675f
C51 VN.n5 VSUBS 0.263613f
C52 VN.n6 VSUBS 0.05685f
C53 VN.n7 VSUBS 0.156118f
C54 VN.t5 VSUBS 0.62675f
C55 VN.t3 VSUBS 0.622923f
C56 VN.t2 VSUBS 0.622923f
C57 VN.t1 VSUBS 0.62675f
C58 VN.n8 VSUBS 0.26371f
C59 VN.n9 VSUBS 0.24514f
C60 VN.n10 VSUBS 0.024788f
C61 VN.n11 VSUBS 0.24514f
C62 VN.n12 VSUBS 0.263613f
C63 VN.n13 VSUBS 3.21813f
C64 B.n0 VSUBS 0.007532f
C65 B.n1 VSUBS 0.007532f
C66 B.n2 VSUBS 0.011139f
C67 B.n3 VSUBS 0.008536f
C68 B.n4 VSUBS 0.008536f
C69 B.n5 VSUBS 0.008536f
C70 B.n6 VSUBS 0.008536f
C71 B.n7 VSUBS 0.008536f
C72 B.n8 VSUBS 0.008536f
C73 B.n9 VSUBS 0.018834f
C74 B.n10 VSUBS 0.008536f
C75 B.n11 VSUBS 0.008536f
C76 B.n12 VSUBS 0.008536f
C77 B.n13 VSUBS 0.008536f
C78 B.n14 VSUBS 0.008536f
C79 B.n15 VSUBS 0.008536f
C80 B.n16 VSUBS 0.008536f
C81 B.n17 VSUBS 0.008536f
C82 B.n18 VSUBS 0.008536f
C83 B.n19 VSUBS 0.008536f
C84 B.n20 VSUBS 0.008536f
C85 B.n21 VSUBS 0.008536f
C86 B.n22 VSUBS 0.008536f
C87 B.n23 VSUBS 0.008536f
C88 B.n24 VSUBS 0.008536f
C89 B.n25 VSUBS 0.008536f
C90 B.n26 VSUBS 0.008536f
C91 B.n27 VSUBS 0.008536f
C92 B.n28 VSUBS 0.008536f
C93 B.n29 VSUBS 0.008536f
C94 B.n30 VSUBS 0.008536f
C95 B.n31 VSUBS 0.008536f
C96 B.n32 VSUBS 0.008536f
C97 B.n33 VSUBS 0.008536f
C98 B.n34 VSUBS 0.008536f
C99 B.n35 VSUBS 0.008536f
C100 B.n36 VSUBS 0.008536f
C101 B.n37 VSUBS 0.008536f
C102 B.t10 VSUBS 0.390689f
C103 B.t11 VSUBS 0.398211f
C104 B.t9 VSUBS 0.140711f
C105 B.n38 VSUBS 0.405845f
C106 B.n39 VSUBS 0.370035f
C107 B.n40 VSUBS 0.008536f
C108 B.n41 VSUBS 0.008536f
C109 B.n42 VSUBS 0.008536f
C110 B.n43 VSUBS 0.008536f
C111 B.t1 VSUBS 0.390693f
C112 B.t2 VSUBS 0.398215f
C113 B.t0 VSUBS 0.140711f
C114 B.n44 VSUBS 0.405841f
C115 B.n45 VSUBS 0.37003f
C116 B.n46 VSUBS 0.019777f
C117 B.n47 VSUBS 0.008536f
C118 B.n48 VSUBS 0.008536f
C119 B.n49 VSUBS 0.008536f
C120 B.n50 VSUBS 0.008536f
C121 B.n51 VSUBS 0.008536f
C122 B.n52 VSUBS 0.008536f
C123 B.n53 VSUBS 0.008536f
C124 B.n54 VSUBS 0.008536f
C125 B.n55 VSUBS 0.008536f
C126 B.n56 VSUBS 0.008536f
C127 B.n57 VSUBS 0.008536f
C128 B.n58 VSUBS 0.008536f
C129 B.n59 VSUBS 0.008536f
C130 B.n60 VSUBS 0.008536f
C131 B.n61 VSUBS 0.008536f
C132 B.n62 VSUBS 0.008536f
C133 B.n63 VSUBS 0.008536f
C134 B.n64 VSUBS 0.008536f
C135 B.n65 VSUBS 0.008536f
C136 B.n66 VSUBS 0.008536f
C137 B.n67 VSUBS 0.008536f
C138 B.n68 VSUBS 0.008536f
C139 B.n69 VSUBS 0.008536f
C140 B.n70 VSUBS 0.008536f
C141 B.n71 VSUBS 0.008536f
C142 B.n72 VSUBS 0.008536f
C143 B.n73 VSUBS 0.008536f
C144 B.n74 VSUBS 0.02033f
C145 B.n75 VSUBS 0.008536f
C146 B.n76 VSUBS 0.008536f
C147 B.n77 VSUBS 0.008536f
C148 B.n78 VSUBS 0.008536f
C149 B.n79 VSUBS 0.008536f
C150 B.n80 VSUBS 0.008536f
C151 B.n81 VSUBS 0.008536f
C152 B.n82 VSUBS 0.008536f
C153 B.n83 VSUBS 0.008536f
C154 B.n84 VSUBS 0.008536f
C155 B.n85 VSUBS 0.008536f
C156 B.n86 VSUBS 0.008536f
C157 B.n87 VSUBS 0.008536f
C158 B.n88 VSUBS 0.008536f
C159 B.n89 VSUBS 0.008536f
C160 B.n90 VSUBS 0.019874f
C161 B.n91 VSUBS 0.008536f
C162 B.n92 VSUBS 0.008536f
C163 B.n93 VSUBS 0.008536f
C164 B.n94 VSUBS 0.008536f
C165 B.n95 VSUBS 0.008536f
C166 B.n96 VSUBS 0.008536f
C167 B.n97 VSUBS 0.008536f
C168 B.n98 VSUBS 0.008536f
C169 B.n99 VSUBS 0.008536f
C170 B.n100 VSUBS 0.008536f
C171 B.n101 VSUBS 0.008536f
C172 B.n102 VSUBS 0.008536f
C173 B.n103 VSUBS 0.008536f
C174 B.n104 VSUBS 0.008536f
C175 B.n105 VSUBS 0.008536f
C176 B.n106 VSUBS 0.008536f
C177 B.n107 VSUBS 0.008536f
C178 B.n108 VSUBS 0.008536f
C179 B.n109 VSUBS 0.008536f
C180 B.n110 VSUBS 0.008536f
C181 B.n111 VSUBS 0.008536f
C182 B.n112 VSUBS 0.008536f
C183 B.n113 VSUBS 0.008536f
C184 B.n114 VSUBS 0.008536f
C185 B.n115 VSUBS 0.008536f
C186 B.n116 VSUBS 0.008536f
C187 B.n117 VSUBS 0.008536f
C188 B.n118 VSUBS 0.0059f
C189 B.n119 VSUBS 0.008536f
C190 B.n120 VSUBS 0.008536f
C191 B.n121 VSUBS 0.008536f
C192 B.n122 VSUBS 0.008536f
C193 B.n123 VSUBS 0.008536f
C194 B.t8 VSUBS 0.390689f
C195 B.t7 VSUBS 0.398211f
C196 B.t6 VSUBS 0.140711f
C197 B.n124 VSUBS 0.405845f
C198 B.n125 VSUBS 0.370035f
C199 B.n126 VSUBS 0.008536f
C200 B.n127 VSUBS 0.008536f
C201 B.n128 VSUBS 0.008536f
C202 B.n129 VSUBS 0.008536f
C203 B.n130 VSUBS 0.008536f
C204 B.n131 VSUBS 0.008536f
C205 B.n132 VSUBS 0.008536f
C206 B.n133 VSUBS 0.008536f
C207 B.n134 VSUBS 0.008536f
C208 B.n135 VSUBS 0.008536f
C209 B.n136 VSUBS 0.008536f
C210 B.n137 VSUBS 0.008536f
C211 B.n138 VSUBS 0.008536f
C212 B.n139 VSUBS 0.008536f
C213 B.n140 VSUBS 0.008536f
C214 B.n141 VSUBS 0.008536f
C215 B.n142 VSUBS 0.008536f
C216 B.n143 VSUBS 0.008536f
C217 B.n144 VSUBS 0.008536f
C218 B.n145 VSUBS 0.008536f
C219 B.n146 VSUBS 0.008536f
C220 B.n147 VSUBS 0.008536f
C221 B.n148 VSUBS 0.008536f
C222 B.n149 VSUBS 0.008536f
C223 B.n150 VSUBS 0.008536f
C224 B.n151 VSUBS 0.008536f
C225 B.n152 VSUBS 0.008536f
C226 B.n153 VSUBS 0.018834f
C227 B.n154 VSUBS 0.008536f
C228 B.n155 VSUBS 0.008536f
C229 B.n156 VSUBS 0.008536f
C230 B.n157 VSUBS 0.008536f
C231 B.n158 VSUBS 0.008536f
C232 B.n159 VSUBS 0.008536f
C233 B.n160 VSUBS 0.008536f
C234 B.n161 VSUBS 0.008536f
C235 B.n162 VSUBS 0.008536f
C236 B.n163 VSUBS 0.008536f
C237 B.n164 VSUBS 0.008536f
C238 B.n165 VSUBS 0.008536f
C239 B.n166 VSUBS 0.008536f
C240 B.n167 VSUBS 0.008536f
C241 B.n168 VSUBS 0.008536f
C242 B.n169 VSUBS 0.008536f
C243 B.n170 VSUBS 0.008536f
C244 B.n171 VSUBS 0.008536f
C245 B.n172 VSUBS 0.008536f
C246 B.n173 VSUBS 0.008536f
C247 B.n174 VSUBS 0.008536f
C248 B.n175 VSUBS 0.008536f
C249 B.n176 VSUBS 0.008536f
C250 B.n177 VSUBS 0.008536f
C251 B.n178 VSUBS 0.008536f
C252 B.n179 VSUBS 0.008536f
C253 B.n180 VSUBS 0.018834f
C254 B.n181 VSUBS 0.02033f
C255 B.n182 VSUBS 0.02033f
C256 B.n183 VSUBS 0.008536f
C257 B.n184 VSUBS 0.008536f
C258 B.n185 VSUBS 0.008536f
C259 B.n186 VSUBS 0.008536f
C260 B.n187 VSUBS 0.008536f
C261 B.n188 VSUBS 0.008536f
C262 B.n189 VSUBS 0.008536f
C263 B.n190 VSUBS 0.008536f
C264 B.n191 VSUBS 0.008536f
C265 B.n192 VSUBS 0.008536f
C266 B.n193 VSUBS 0.008536f
C267 B.n194 VSUBS 0.008536f
C268 B.n195 VSUBS 0.008536f
C269 B.n196 VSUBS 0.008536f
C270 B.n197 VSUBS 0.008536f
C271 B.n198 VSUBS 0.008536f
C272 B.n199 VSUBS 0.008536f
C273 B.n200 VSUBS 0.008536f
C274 B.n201 VSUBS 0.008536f
C275 B.n202 VSUBS 0.008536f
C276 B.n203 VSUBS 0.008536f
C277 B.n204 VSUBS 0.008536f
C278 B.n205 VSUBS 0.008536f
C279 B.n206 VSUBS 0.008536f
C280 B.n207 VSUBS 0.008536f
C281 B.n208 VSUBS 0.008536f
C282 B.n209 VSUBS 0.008536f
C283 B.n210 VSUBS 0.008536f
C284 B.n211 VSUBS 0.008536f
C285 B.n212 VSUBS 0.008536f
C286 B.n213 VSUBS 0.008536f
C287 B.n214 VSUBS 0.008536f
C288 B.n215 VSUBS 0.008536f
C289 B.n216 VSUBS 0.008536f
C290 B.n217 VSUBS 0.008536f
C291 B.n218 VSUBS 0.008536f
C292 B.n219 VSUBS 0.008536f
C293 B.n220 VSUBS 0.008536f
C294 B.n221 VSUBS 0.008536f
C295 B.n222 VSUBS 0.008536f
C296 B.n223 VSUBS 0.008536f
C297 B.n224 VSUBS 0.008536f
C298 B.n225 VSUBS 0.008536f
C299 B.n226 VSUBS 0.008536f
C300 B.n227 VSUBS 0.008536f
C301 B.n228 VSUBS 0.008536f
C302 B.n229 VSUBS 0.008536f
C303 B.n230 VSUBS 0.008536f
C304 B.n231 VSUBS 0.008536f
C305 B.n232 VSUBS 0.008536f
C306 B.n233 VSUBS 0.008536f
C307 B.n234 VSUBS 0.008536f
C308 B.n235 VSUBS 0.008536f
C309 B.n236 VSUBS 0.008536f
C310 B.n237 VSUBS 0.008536f
C311 B.n238 VSUBS 0.008536f
C312 B.n239 VSUBS 0.008536f
C313 B.n240 VSUBS 0.008536f
C314 B.n241 VSUBS 0.008536f
C315 B.n242 VSUBS 0.008536f
C316 B.n243 VSUBS 0.008536f
C317 B.n244 VSUBS 0.008536f
C318 B.n245 VSUBS 0.008536f
C319 B.n246 VSUBS 0.008536f
C320 B.n247 VSUBS 0.008536f
C321 B.n248 VSUBS 0.008536f
C322 B.n249 VSUBS 0.008536f
C323 B.n250 VSUBS 0.008536f
C324 B.n251 VSUBS 0.008536f
C325 B.n252 VSUBS 0.008536f
C326 B.n253 VSUBS 0.008536f
C327 B.n254 VSUBS 0.008536f
C328 B.n255 VSUBS 0.008536f
C329 B.n256 VSUBS 0.008536f
C330 B.n257 VSUBS 0.008536f
C331 B.n258 VSUBS 0.008536f
C332 B.n259 VSUBS 0.008536f
C333 B.n260 VSUBS 0.008536f
C334 B.n261 VSUBS 0.008536f
C335 B.n262 VSUBS 0.008536f
C336 B.n263 VSUBS 0.008536f
C337 B.n264 VSUBS 0.0059f
C338 B.n265 VSUBS 0.019777f
C339 B.n266 VSUBS 0.006904f
C340 B.n267 VSUBS 0.008536f
C341 B.n268 VSUBS 0.008536f
C342 B.n269 VSUBS 0.008536f
C343 B.n270 VSUBS 0.008536f
C344 B.n271 VSUBS 0.008536f
C345 B.n272 VSUBS 0.008536f
C346 B.n273 VSUBS 0.008536f
C347 B.n274 VSUBS 0.008536f
C348 B.n275 VSUBS 0.008536f
C349 B.n276 VSUBS 0.008536f
C350 B.n277 VSUBS 0.008536f
C351 B.t5 VSUBS 0.390693f
C352 B.t4 VSUBS 0.398215f
C353 B.t3 VSUBS 0.140711f
C354 B.n278 VSUBS 0.405841f
C355 B.n279 VSUBS 0.37003f
C356 B.n280 VSUBS 0.019777f
C357 B.n281 VSUBS 0.006904f
C358 B.n282 VSUBS 0.008536f
C359 B.n283 VSUBS 0.008536f
C360 B.n284 VSUBS 0.008536f
C361 B.n285 VSUBS 0.008536f
C362 B.n286 VSUBS 0.008536f
C363 B.n287 VSUBS 0.008536f
C364 B.n288 VSUBS 0.008536f
C365 B.n289 VSUBS 0.008536f
C366 B.n290 VSUBS 0.008536f
C367 B.n291 VSUBS 0.008536f
C368 B.n292 VSUBS 0.008536f
C369 B.n293 VSUBS 0.008536f
C370 B.n294 VSUBS 0.008536f
C371 B.n295 VSUBS 0.008536f
C372 B.n296 VSUBS 0.008536f
C373 B.n297 VSUBS 0.008536f
C374 B.n298 VSUBS 0.008536f
C375 B.n299 VSUBS 0.008536f
C376 B.n300 VSUBS 0.008536f
C377 B.n301 VSUBS 0.008536f
C378 B.n302 VSUBS 0.008536f
C379 B.n303 VSUBS 0.008536f
C380 B.n304 VSUBS 0.008536f
C381 B.n305 VSUBS 0.008536f
C382 B.n306 VSUBS 0.008536f
C383 B.n307 VSUBS 0.008536f
C384 B.n308 VSUBS 0.008536f
C385 B.n309 VSUBS 0.008536f
C386 B.n310 VSUBS 0.008536f
C387 B.n311 VSUBS 0.008536f
C388 B.n312 VSUBS 0.008536f
C389 B.n313 VSUBS 0.008536f
C390 B.n314 VSUBS 0.008536f
C391 B.n315 VSUBS 0.008536f
C392 B.n316 VSUBS 0.008536f
C393 B.n317 VSUBS 0.008536f
C394 B.n318 VSUBS 0.008536f
C395 B.n319 VSUBS 0.008536f
C396 B.n320 VSUBS 0.008536f
C397 B.n321 VSUBS 0.008536f
C398 B.n322 VSUBS 0.008536f
C399 B.n323 VSUBS 0.008536f
C400 B.n324 VSUBS 0.008536f
C401 B.n325 VSUBS 0.008536f
C402 B.n326 VSUBS 0.008536f
C403 B.n327 VSUBS 0.008536f
C404 B.n328 VSUBS 0.008536f
C405 B.n329 VSUBS 0.008536f
C406 B.n330 VSUBS 0.008536f
C407 B.n331 VSUBS 0.008536f
C408 B.n332 VSUBS 0.008536f
C409 B.n333 VSUBS 0.008536f
C410 B.n334 VSUBS 0.008536f
C411 B.n335 VSUBS 0.008536f
C412 B.n336 VSUBS 0.008536f
C413 B.n337 VSUBS 0.008536f
C414 B.n338 VSUBS 0.008536f
C415 B.n339 VSUBS 0.008536f
C416 B.n340 VSUBS 0.008536f
C417 B.n341 VSUBS 0.008536f
C418 B.n342 VSUBS 0.008536f
C419 B.n343 VSUBS 0.008536f
C420 B.n344 VSUBS 0.008536f
C421 B.n345 VSUBS 0.008536f
C422 B.n346 VSUBS 0.008536f
C423 B.n347 VSUBS 0.008536f
C424 B.n348 VSUBS 0.008536f
C425 B.n349 VSUBS 0.008536f
C426 B.n350 VSUBS 0.008536f
C427 B.n351 VSUBS 0.008536f
C428 B.n352 VSUBS 0.008536f
C429 B.n353 VSUBS 0.008536f
C430 B.n354 VSUBS 0.008536f
C431 B.n355 VSUBS 0.008536f
C432 B.n356 VSUBS 0.008536f
C433 B.n357 VSUBS 0.008536f
C434 B.n358 VSUBS 0.008536f
C435 B.n359 VSUBS 0.008536f
C436 B.n360 VSUBS 0.008536f
C437 B.n361 VSUBS 0.008536f
C438 B.n362 VSUBS 0.008536f
C439 B.n363 VSUBS 0.008536f
C440 B.n364 VSUBS 0.008536f
C441 B.n365 VSUBS 0.019291f
C442 B.n366 VSUBS 0.02033f
C443 B.n367 VSUBS 0.018834f
C444 B.n368 VSUBS 0.008536f
C445 B.n369 VSUBS 0.008536f
C446 B.n370 VSUBS 0.008536f
C447 B.n371 VSUBS 0.008536f
C448 B.n372 VSUBS 0.008536f
C449 B.n373 VSUBS 0.008536f
C450 B.n374 VSUBS 0.008536f
C451 B.n375 VSUBS 0.008536f
C452 B.n376 VSUBS 0.008536f
C453 B.n377 VSUBS 0.008536f
C454 B.n378 VSUBS 0.008536f
C455 B.n379 VSUBS 0.008536f
C456 B.n380 VSUBS 0.008536f
C457 B.n381 VSUBS 0.008536f
C458 B.n382 VSUBS 0.008536f
C459 B.n383 VSUBS 0.008536f
C460 B.n384 VSUBS 0.008536f
C461 B.n385 VSUBS 0.008536f
C462 B.n386 VSUBS 0.008536f
C463 B.n387 VSUBS 0.008536f
C464 B.n388 VSUBS 0.008536f
C465 B.n389 VSUBS 0.008536f
C466 B.n390 VSUBS 0.008536f
C467 B.n391 VSUBS 0.008536f
C468 B.n392 VSUBS 0.008536f
C469 B.n393 VSUBS 0.008536f
C470 B.n394 VSUBS 0.008536f
C471 B.n395 VSUBS 0.008536f
C472 B.n396 VSUBS 0.008536f
C473 B.n397 VSUBS 0.008536f
C474 B.n398 VSUBS 0.008536f
C475 B.n399 VSUBS 0.008536f
C476 B.n400 VSUBS 0.008536f
C477 B.n401 VSUBS 0.008536f
C478 B.n402 VSUBS 0.008536f
C479 B.n403 VSUBS 0.008536f
C480 B.n404 VSUBS 0.008536f
C481 B.n405 VSUBS 0.008536f
C482 B.n406 VSUBS 0.008536f
C483 B.n407 VSUBS 0.008536f
C484 B.n408 VSUBS 0.008536f
C485 B.n409 VSUBS 0.008536f
C486 B.n410 VSUBS 0.008536f
C487 B.n411 VSUBS 0.008536f
C488 B.n412 VSUBS 0.008536f
C489 B.n413 VSUBS 0.018834f
C490 B.n414 VSUBS 0.018834f
C491 B.n415 VSUBS 0.02033f
C492 B.n416 VSUBS 0.008536f
C493 B.n417 VSUBS 0.008536f
C494 B.n418 VSUBS 0.008536f
C495 B.n419 VSUBS 0.008536f
C496 B.n420 VSUBS 0.008536f
C497 B.n421 VSUBS 0.008536f
C498 B.n422 VSUBS 0.008536f
C499 B.n423 VSUBS 0.008536f
C500 B.n424 VSUBS 0.008536f
C501 B.n425 VSUBS 0.008536f
C502 B.n426 VSUBS 0.008536f
C503 B.n427 VSUBS 0.008536f
C504 B.n428 VSUBS 0.008536f
C505 B.n429 VSUBS 0.008536f
C506 B.n430 VSUBS 0.008536f
C507 B.n431 VSUBS 0.008536f
C508 B.n432 VSUBS 0.008536f
C509 B.n433 VSUBS 0.008536f
C510 B.n434 VSUBS 0.008536f
C511 B.n435 VSUBS 0.008536f
C512 B.n436 VSUBS 0.008536f
C513 B.n437 VSUBS 0.008536f
C514 B.n438 VSUBS 0.008536f
C515 B.n439 VSUBS 0.008536f
C516 B.n440 VSUBS 0.008536f
C517 B.n441 VSUBS 0.008536f
C518 B.n442 VSUBS 0.008536f
C519 B.n443 VSUBS 0.008536f
C520 B.n444 VSUBS 0.008536f
C521 B.n445 VSUBS 0.008536f
C522 B.n446 VSUBS 0.008536f
C523 B.n447 VSUBS 0.008536f
C524 B.n448 VSUBS 0.008536f
C525 B.n449 VSUBS 0.008536f
C526 B.n450 VSUBS 0.008536f
C527 B.n451 VSUBS 0.008536f
C528 B.n452 VSUBS 0.008536f
C529 B.n453 VSUBS 0.008536f
C530 B.n454 VSUBS 0.008536f
C531 B.n455 VSUBS 0.008536f
C532 B.n456 VSUBS 0.008536f
C533 B.n457 VSUBS 0.008536f
C534 B.n458 VSUBS 0.008536f
C535 B.n459 VSUBS 0.008536f
C536 B.n460 VSUBS 0.008536f
C537 B.n461 VSUBS 0.008536f
C538 B.n462 VSUBS 0.008536f
C539 B.n463 VSUBS 0.008536f
C540 B.n464 VSUBS 0.008536f
C541 B.n465 VSUBS 0.008536f
C542 B.n466 VSUBS 0.008536f
C543 B.n467 VSUBS 0.008536f
C544 B.n468 VSUBS 0.008536f
C545 B.n469 VSUBS 0.008536f
C546 B.n470 VSUBS 0.008536f
C547 B.n471 VSUBS 0.008536f
C548 B.n472 VSUBS 0.008536f
C549 B.n473 VSUBS 0.008536f
C550 B.n474 VSUBS 0.008536f
C551 B.n475 VSUBS 0.008536f
C552 B.n476 VSUBS 0.008536f
C553 B.n477 VSUBS 0.008536f
C554 B.n478 VSUBS 0.008536f
C555 B.n479 VSUBS 0.008536f
C556 B.n480 VSUBS 0.008536f
C557 B.n481 VSUBS 0.008536f
C558 B.n482 VSUBS 0.008536f
C559 B.n483 VSUBS 0.008536f
C560 B.n484 VSUBS 0.008536f
C561 B.n485 VSUBS 0.008536f
C562 B.n486 VSUBS 0.008536f
C563 B.n487 VSUBS 0.008536f
C564 B.n488 VSUBS 0.008536f
C565 B.n489 VSUBS 0.008536f
C566 B.n490 VSUBS 0.008536f
C567 B.n491 VSUBS 0.008536f
C568 B.n492 VSUBS 0.008536f
C569 B.n493 VSUBS 0.008536f
C570 B.n494 VSUBS 0.008536f
C571 B.n495 VSUBS 0.008536f
C572 B.n496 VSUBS 0.008536f
C573 B.n497 VSUBS 0.0059f
C574 B.n498 VSUBS 0.008536f
C575 B.n499 VSUBS 0.008536f
C576 B.n500 VSUBS 0.006904f
C577 B.n501 VSUBS 0.008536f
C578 B.n502 VSUBS 0.008536f
C579 B.n503 VSUBS 0.008536f
C580 B.n504 VSUBS 0.008536f
C581 B.n505 VSUBS 0.008536f
C582 B.n506 VSUBS 0.008536f
C583 B.n507 VSUBS 0.008536f
C584 B.n508 VSUBS 0.008536f
C585 B.n509 VSUBS 0.008536f
C586 B.n510 VSUBS 0.008536f
C587 B.n511 VSUBS 0.008536f
C588 B.n512 VSUBS 0.006904f
C589 B.n513 VSUBS 0.019777f
C590 B.n514 VSUBS 0.0059f
C591 B.n515 VSUBS 0.008536f
C592 B.n516 VSUBS 0.008536f
C593 B.n517 VSUBS 0.008536f
C594 B.n518 VSUBS 0.008536f
C595 B.n519 VSUBS 0.008536f
C596 B.n520 VSUBS 0.008536f
C597 B.n521 VSUBS 0.008536f
C598 B.n522 VSUBS 0.008536f
C599 B.n523 VSUBS 0.008536f
C600 B.n524 VSUBS 0.008536f
C601 B.n525 VSUBS 0.008536f
C602 B.n526 VSUBS 0.008536f
C603 B.n527 VSUBS 0.008536f
C604 B.n528 VSUBS 0.008536f
C605 B.n529 VSUBS 0.008536f
C606 B.n530 VSUBS 0.008536f
C607 B.n531 VSUBS 0.008536f
C608 B.n532 VSUBS 0.008536f
C609 B.n533 VSUBS 0.008536f
C610 B.n534 VSUBS 0.008536f
C611 B.n535 VSUBS 0.008536f
C612 B.n536 VSUBS 0.008536f
C613 B.n537 VSUBS 0.008536f
C614 B.n538 VSUBS 0.008536f
C615 B.n539 VSUBS 0.008536f
C616 B.n540 VSUBS 0.008536f
C617 B.n541 VSUBS 0.008536f
C618 B.n542 VSUBS 0.008536f
C619 B.n543 VSUBS 0.008536f
C620 B.n544 VSUBS 0.008536f
C621 B.n545 VSUBS 0.008536f
C622 B.n546 VSUBS 0.008536f
C623 B.n547 VSUBS 0.008536f
C624 B.n548 VSUBS 0.008536f
C625 B.n549 VSUBS 0.008536f
C626 B.n550 VSUBS 0.008536f
C627 B.n551 VSUBS 0.008536f
C628 B.n552 VSUBS 0.008536f
C629 B.n553 VSUBS 0.008536f
C630 B.n554 VSUBS 0.008536f
C631 B.n555 VSUBS 0.008536f
C632 B.n556 VSUBS 0.008536f
C633 B.n557 VSUBS 0.008536f
C634 B.n558 VSUBS 0.008536f
C635 B.n559 VSUBS 0.008536f
C636 B.n560 VSUBS 0.008536f
C637 B.n561 VSUBS 0.008536f
C638 B.n562 VSUBS 0.008536f
C639 B.n563 VSUBS 0.008536f
C640 B.n564 VSUBS 0.008536f
C641 B.n565 VSUBS 0.008536f
C642 B.n566 VSUBS 0.008536f
C643 B.n567 VSUBS 0.008536f
C644 B.n568 VSUBS 0.008536f
C645 B.n569 VSUBS 0.008536f
C646 B.n570 VSUBS 0.008536f
C647 B.n571 VSUBS 0.008536f
C648 B.n572 VSUBS 0.008536f
C649 B.n573 VSUBS 0.008536f
C650 B.n574 VSUBS 0.008536f
C651 B.n575 VSUBS 0.008536f
C652 B.n576 VSUBS 0.008536f
C653 B.n577 VSUBS 0.008536f
C654 B.n578 VSUBS 0.008536f
C655 B.n579 VSUBS 0.008536f
C656 B.n580 VSUBS 0.008536f
C657 B.n581 VSUBS 0.008536f
C658 B.n582 VSUBS 0.008536f
C659 B.n583 VSUBS 0.008536f
C660 B.n584 VSUBS 0.008536f
C661 B.n585 VSUBS 0.008536f
C662 B.n586 VSUBS 0.008536f
C663 B.n587 VSUBS 0.008536f
C664 B.n588 VSUBS 0.008536f
C665 B.n589 VSUBS 0.008536f
C666 B.n590 VSUBS 0.008536f
C667 B.n591 VSUBS 0.008536f
C668 B.n592 VSUBS 0.008536f
C669 B.n593 VSUBS 0.008536f
C670 B.n594 VSUBS 0.008536f
C671 B.n595 VSUBS 0.008536f
C672 B.n596 VSUBS 0.02033f
C673 B.n597 VSUBS 0.02033f
C674 B.n598 VSUBS 0.018834f
C675 B.n599 VSUBS 0.008536f
C676 B.n600 VSUBS 0.008536f
C677 B.n601 VSUBS 0.008536f
C678 B.n602 VSUBS 0.008536f
C679 B.n603 VSUBS 0.008536f
C680 B.n604 VSUBS 0.008536f
C681 B.n605 VSUBS 0.008536f
C682 B.n606 VSUBS 0.008536f
C683 B.n607 VSUBS 0.008536f
C684 B.n608 VSUBS 0.008536f
C685 B.n609 VSUBS 0.008536f
C686 B.n610 VSUBS 0.008536f
C687 B.n611 VSUBS 0.008536f
C688 B.n612 VSUBS 0.008536f
C689 B.n613 VSUBS 0.008536f
C690 B.n614 VSUBS 0.008536f
C691 B.n615 VSUBS 0.008536f
C692 B.n616 VSUBS 0.008536f
C693 B.n617 VSUBS 0.008536f
C694 B.n618 VSUBS 0.008536f
C695 B.n619 VSUBS 0.011139f
C696 B.n620 VSUBS 0.011866f
C697 B.n621 VSUBS 0.023596f
C698 VTAIL.t2 VSUBS 0.426295f
C699 VTAIL.t3 VSUBS 0.426295f
C700 VTAIL.n0 VSUBS 3.29534f
C701 VTAIL.n1 VSUBS 0.850873f
C702 VTAIL.n2 VSUBS 0.033245f
C703 VTAIL.n3 VSUBS 0.032245f
C704 VTAIL.n4 VSUBS 0.017327f
C705 VTAIL.n5 VSUBS 0.040955f
C706 VTAIL.n6 VSUBS 0.018346f
C707 VTAIL.n7 VSUBS 0.032245f
C708 VTAIL.n8 VSUBS 0.017327f
C709 VTAIL.n9 VSUBS 0.040955f
C710 VTAIL.n10 VSUBS 0.018346f
C711 VTAIL.n11 VSUBS 0.032245f
C712 VTAIL.n12 VSUBS 0.017327f
C713 VTAIL.n13 VSUBS 0.040955f
C714 VTAIL.n14 VSUBS 0.018346f
C715 VTAIL.n15 VSUBS 0.032245f
C716 VTAIL.n16 VSUBS 0.017327f
C717 VTAIL.n17 VSUBS 0.040955f
C718 VTAIL.n18 VSUBS 0.018346f
C719 VTAIL.n19 VSUBS 0.032245f
C720 VTAIL.n20 VSUBS 0.017327f
C721 VTAIL.n21 VSUBS 0.040955f
C722 VTAIL.n22 VSUBS 0.018346f
C723 VTAIL.n23 VSUBS 0.032245f
C724 VTAIL.n24 VSUBS 0.017327f
C725 VTAIL.n25 VSUBS 0.040955f
C726 VTAIL.n26 VSUBS 0.018346f
C727 VTAIL.n27 VSUBS 0.032245f
C728 VTAIL.n28 VSUBS 0.017327f
C729 VTAIL.n29 VSUBS 0.040955f
C730 VTAIL.n30 VSUBS 0.018346f
C731 VTAIL.n31 VSUBS 0.243752f
C732 VTAIL.t0 VSUBS 0.087814f
C733 VTAIL.n32 VSUBS 0.030716f
C734 VTAIL.n33 VSUBS 0.026053f
C735 VTAIL.n34 VSUBS 0.017327f
C736 VTAIL.n35 VSUBS 2.31214f
C737 VTAIL.n36 VSUBS 0.032245f
C738 VTAIL.n37 VSUBS 0.017327f
C739 VTAIL.n38 VSUBS 0.018346f
C740 VTAIL.n39 VSUBS 0.040955f
C741 VTAIL.n40 VSUBS 0.040955f
C742 VTAIL.n41 VSUBS 0.018346f
C743 VTAIL.n42 VSUBS 0.017327f
C744 VTAIL.n43 VSUBS 0.032245f
C745 VTAIL.n44 VSUBS 0.032245f
C746 VTAIL.n45 VSUBS 0.017327f
C747 VTAIL.n46 VSUBS 0.018346f
C748 VTAIL.n47 VSUBS 0.040955f
C749 VTAIL.n48 VSUBS 0.040955f
C750 VTAIL.n49 VSUBS 0.018346f
C751 VTAIL.n50 VSUBS 0.017327f
C752 VTAIL.n51 VSUBS 0.032245f
C753 VTAIL.n52 VSUBS 0.032245f
C754 VTAIL.n53 VSUBS 0.017327f
C755 VTAIL.n54 VSUBS 0.018346f
C756 VTAIL.n55 VSUBS 0.040955f
C757 VTAIL.n56 VSUBS 0.040955f
C758 VTAIL.n57 VSUBS 0.018346f
C759 VTAIL.n58 VSUBS 0.017327f
C760 VTAIL.n59 VSUBS 0.032245f
C761 VTAIL.n60 VSUBS 0.032245f
C762 VTAIL.n61 VSUBS 0.017327f
C763 VTAIL.n62 VSUBS 0.018346f
C764 VTAIL.n63 VSUBS 0.040955f
C765 VTAIL.n64 VSUBS 0.040955f
C766 VTAIL.n65 VSUBS 0.018346f
C767 VTAIL.n66 VSUBS 0.017327f
C768 VTAIL.n67 VSUBS 0.032245f
C769 VTAIL.n68 VSUBS 0.032245f
C770 VTAIL.n69 VSUBS 0.017327f
C771 VTAIL.n70 VSUBS 0.018346f
C772 VTAIL.n71 VSUBS 0.040955f
C773 VTAIL.n72 VSUBS 0.040955f
C774 VTAIL.n73 VSUBS 0.040955f
C775 VTAIL.n74 VSUBS 0.018346f
C776 VTAIL.n75 VSUBS 0.017327f
C777 VTAIL.n76 VSUBS 0.032245f
C778 VTAIL.n77 VSUBS 0.032245f
C779 VTAIL.n78 VSUBS 0.017327f
C780 VTAIL.n79 VSUBS 0.017837f
C781 VTAIL.n80 VSUBS 0.017837f
C782 VTAIL.n81 VSUBS 0.040955f
C783 VTAIL.n82 VSUBS 0.040955f
C784 VTAIL.n83 VSUBS 0.018346f
C785 VTAIL.n84 VSUBS 0.017327f
C786 VTAIL.n85 VSUBS 0.032245f
C787 VTAIL.n86 VSUBS 0.032245f
C788 VTAIL.n87 VSUBS 0.017327f
C789 VTAIL.n88 VSUBS 0.018346f
C790 VTAIL.n89 VSUBS 0.040955f
C791 VTAIL.n90 VSUBS 0.091704f
C792 VTAIL.n91 VSUBS 0.018346f
C793 VTAIL.n92 VSUBS 0.017327f
C794 VTAIL.n93 VSUBS 0.071449f
C795 VTAIL.n94 VSUBS 0.04569f
C796 VTAIL.n95 VSUBS 0.120296f
C797 VTAIL.n96 VSUBS 0.033245f
C798 VTAIL.n97 VSUBS 0.032245f
C799 VTAIL.n98 VSUBS 0.017327f
C800 VTAIL.n99 VSUBS 0.040955f
C801 VTAIL.n100 VSUBS 0.018346f
C802 VTAIL.n101 VSUBS 0.032245f
C803 VTAIL.n102 VSUBS 0.017327f
C804 VTAIL.n103 VSUBS 0.040955f
C805 VTAIL.n104 VSUBS 0.018346f
C806 VTAIL.n105 VSUBS 0.032245f
C807 VTAIL.n106 VSUBS 0.017327f
C808 VTAIL.n107 VSUBS 0.040955f
C809 VTAIL.n108 VSUBS 0.018346f
C810 VTAIL.n109 VSUBS 0.032245f
C811 VTAIL.n110 VSUBS 0.017327f
C812 VTAIL.n111 VSUBS 0.040955f
C813 VTAIL.n112 VSUBS 0.018346f
C814 VTAIL.n113 VSUBS 0.032245f
C815 VTAIL.n114 VSUBS 0.017327f
C816 VTAIL.n115 VSUBS 0.040955f
C817 VTAIL.n116 VSUBS 0.018346f
C818 VTAIL.n117 VSUBS 0.032245f
C819 VTAIL.n118 VSUBS 0.017327f
C820 VTAIL.n119 VSUBS 0.040955f
C821 VTAIL.n120 VSUBS 0.018346f
C822 VTAIL.n121 VSUBS 0.032245f
C823 VTAIL.n122 VSUBS 0.017327f
C824 VTAIL.n123 VSUBS 0.040955f
C825 VTAIL.n124 VSUBS 0.018346f
C826 VTAIL.n125 VSUBS 0.243752f
C827 VTAIL.t8 VSUBS 0.087814f
C828 VTAIL.n126 VSUBS 0.030716f
C829 VTAIL.n127 VSUBS 0.026053f
C830 VTAIL.n128 VSUBS 0.017327f
C831 VTAIL.n129 VSUBS 2.31214f
C832 VTAIL.n130 VSUBS 0.032245f
C833 VTAIL.n131 VSUBS 0.017327f
C834 VTAIL.n132 VSUBS 0.018346f
C835 VTAIL.n133 VSUBS 0.040955f
C836 VTAIL.n134 VSUBS 0.040955f
C837 VTAIL.n135 VSUBS 0.018346f
C838 VTAIL.n136 VSUBS 0.017327f
C839 VTAIL.n137 VSUBS 0.032245f
C840 VTAIL.n138 VSUBS 0.032245f
C841 VTAIL.n139 VSUBS 0.017327f
C842 VTAIL.n140 VSUBS 0.018346f
C843 VTAIL.n141 VSUBS 0.040955f
C844 VTAIL.n142 VSUBS 0.040955f
C845 VTAIL.n143 VSUBS 0.018346f
C846 VTAIL.n144 VSUBS 0.017327f
C847 VTAIL.n145 VSUBS 0.032245f
C848 VTAIL.n146 VSUBS 0.032245f
C849 VTAIL.n147 VSUBS 0.017327f
C850 VTAIL.n148 VSUBS 0.018346f
C851 VTAIL.n149 VSUBS 0.040955f
C852 VTAIL.n150 VSUBS 0.040955f
C853 VTAIL.n151 VSUBS 0.018346f
C854 VTAIL.n152 VSUBS 0.017327f
C855 VTAIL.n153 VSUBS 0.032245f
C856 VTAIL.n154 VSUBS 0.032245f
C857 VTAIL.n155 VSUBS 0.017327f
C858 VTAIL.n156 VSUBS 0.018346f
C859 VTAIL.n157 VSUBS 0.040955f
C860 VTAIL.n158 VSUBS 0.040955f
C861 VTAIL.n159 VSUBS 0.018346f
C862 VTAIL.n160 VSUBS 0.017327f
C863 VTAIL.n161 VSUBS 0.032245f
C864 VTAIL.n162 VSUBS 0.032245f
C865 VTAIL.n163 VSUBS 0.017327f
C866 VTAIL.n164 VSUBS 0.018346f
C867 VTAIL.n165 VSUBS 0.040955f
C868 VTAIL.n166 VSUBS 0.040955f
C869 VTAIL.n167 VSUBS 0.040955f
C870 VTAIL.n168 VSUBS 0.018346f
C871 VTAIL.n169 VSUBS 0.017327f
C872 VTAIL.n170 VSUBS 0.032245f
C873 VTAIL.n171 VSUBS 0.032245f
C874 VTAIL.n172 VSUBS 0.017327f
C875 VTAIL.n173 VSUBS 0.017837f
C876 VTAIL.n174 VSUBS 0.017837f
C877 VTAIL.n175 VSUBS 0.040955f
C878 VTAIL.n176 VSUBS 0.040955f
C879 VTAIL.n177 VSUBS 0.018346f
C880 VTAIL.n178 VSUBS 0.017327f
C881 VTAIL.n179 VSUBS 0.032245f
C882 VTAIL.n180 VSUBS 0.032245f
C883 VTAIL.n181 VSUBS 0.017327f
C884 VTAIL.n182 VSUBS 0.018346f
C885 VTAIL.n183 VSUBS 0.040955f
C886 VTAIL.n184 VSUBS 0.091704f
C887 VTAIL.n185 VSUBS 0.018346f
C888 VTAIL.n186 VSUBS 0.017327f
C889 VTAIL.n187 VSUBS 0.071449f
C890 VTAIL.n188 VSUBS 0.04569f
C891 VTAIL.n189 VSUBS 0.120296f
C892 VTAIL.t14 VSUBS 0.426295f
C893 VTAIL.t15 VSUBS 0.426295f
C894 VTAIL.n190 VSUBS 3.29534f
C895 VTAIL.n191 VSUBS 0.890507f
C896 VTAIL.n192 VSUBS 0.033245f
C897 VTAIL.n193 VSUBS 0.032245f
C898 VTAIL.n194 VSUBS 0.017327f
C899 VTAIL.n195 VSUBS 0.040955f
C900 VTAIL.n196 VSUBS 0.018346f
C901 VTAIL.n197 VSUBS 0.032245f
C902 VTAIL.n198 VSUBS 0.017327f
C903 VTAIL.n199 VSUBS 0.040955f
C904 VTAIL.n200 VSUBS 0.018346f
C905 VTAIL.n201 VSUBS 0.032245f
C906 VTAIL.n202 VSUBS 0.017327f
C907 VTAIL.n203 VSUBS 0.040955f
C908 VTAIL.n204 VSUBS 0.018346f
C909 VTAIL.n205 VSUBS 0.032245f
C910 VTAIL.n206 VSUBS 0.017327f
C911 VTAIL.n207 VSUBS 0.040955f
C912 VTAIL.n208 VSUBS 0.018346f
C913 VTAIL.n209 VSUBS 0.032245f
C914 VTAIL.n210 VSUBS 0.017327f
C915 VTAIL.n211 VSUBS 0.040955f
C916 VTAIL.n212 VSUBS 0.018346f
C917 VTAIL.n213 VSUBS 0.032245f
C918 VTAIL.n214 VSUBS 0.017327f
C919 VTAIL.n215 VSUBS 0.040955f
C920 VTAIL.n216 VSUBS 0.018346f
C921 VTAIL.n217 VSUBS 0.032245f
C922 VTAIL.n218 VSUBS 0.017327f
C923 VTAIL.n219 VSUBS 0.040955f
C924 VTAIL.n220 VSUBS 0.018346f
C925 VTAIL.n221 VSUBS 0.243752f
C926 VTAIL.t10 VSUBS 0.087814f
C927 VTAIL.n222 VSUBS 0.030716f
C928 VTAIL.n223 VSUBS 0.026053f
C929 VTAIL.n224 VSUBS 0.017327f
C930 VTAIL.n225 VSUBS 2.31214f
C931 VTAIL.n226 VSUBS 0.032245f
C932 VTAIL.n227 VSUBS 0.017327f
C933 VTAIL.n228 VSUBS 0.018346f
C934 VTAIL.n229 VSUBS 0.040955f
C935 VTAIL.n230 VSUBS 0.040955f
C936 VTAIL.n231 VSUBS 0.018346f
C937 VTAIL.n232 VSUBS 0.017327f
C938 VTAIL.n233 VSUBS 0.032245f
C939 VTAIL.n234 VSUBS 0.032245f
C940 VTAIL.n235 VSUBS 0.017327f
C941 VTAIL.n236 VSUBS 0.018346f
C942 VTAIL.n237 VSUBS 0.040955f
C943 VTAIL.n238 VSUBS 0.040955f
C944 VTAIL.n239 VSUBS 0.018346f
C945 VTAIL.n240 VSUBS 0.017327f
C946 VTAIL.n241 VSUBS 0.032245f
C947 VTAIL.n242 VSUBS 0.032245f
C948 VTAIL.n243 VSUBS 0.017327f
C949 VTAIL.n244 VSUBS 0.018346f
C950 VTAIL.n245 VSUBS 0.040955f
C951 VTAIL.n246 VSUBS 0.040955f
C952 VTAIL.n247 VSUBS 0.018346f
C953 VTAIL.n248 VSUBS 0.017327f
C954 VTAIL.n249 VSUBS 0.032245f
C955 VTAIL.n250 VSUBS 0.032245f
C956 VTAIL.n251 VSUBS 0.017327f
C957 VTAIL.n252 VSUBS 0.018346f
C958 VTAIL.n253 VSUBS 0.040955f
C959 VTAIL.n254 VSUBS 0.040955f
C960 VTAIL.n255 VSUBS 0.018346f
C961 VTAIL.n256 VSUBS 0.017327f
C962 VTAIL.n257 VSUBS 0.032245f
C963 VTAIL.n258 VSUBS 0.032245f
C964 VTAIL.n259 VSUBS 0.017327f
C965 VTAIL.n260 VSUBS 0.018346f
C966 VTAIL.n261 VSUBS 0.040955f
C967 VTAIL.n262 VSUBS 0.040955f
C968 VTAIL.n263 VSUBS 0.040955f
C969 VTAIL.n264 VSUBS 0.018346f
C970 VTAIL.n265 VSUBS 0.017327f
C971 VTAIL.n266 VSUBS 0.032245f
C972 VTAIL.n267 VSUBS 0.032245f
C973 VTAIL.n268 VSUBS 0.017327f
C974 VTAIL.n269 VSUBS 0.017837f
C975 VTAIL.n270 VSUBS 0.017837f
C976 VTAIL.n271 VSUBS 0.040955f
C977 VTAIL.n272 VSUBS 0.040955f
C978 VTAIL.n273 VSUBS 0.018346f
C979 VTAIL.n274 VSUBS 0.017327f
C980 VTAIL.n275 VSUBS 0.032245f
C981 VTAIL.n276 VSUBS 0.032245f
C982 VTAIL.n277 VSUBS 0.017327f
C983 VTAIL.n278 VSUBS 0.018346f
C984 VTAIL.n279 VSUBS 0.040955f
C985 VTAIL.n280 VSUBS 0.091704f
C986 VTAIL.n281 VSUBS 0.018346f
C987 VTAIL.n282 VSUBS 0.017327f
C988 VTAIL.n283 VSUBS 0.071449f
C989 VTAIL.n284 VSUBS 0.04569f
C990 VTAIL.n285 VSUBS 2.05366f
C991 VTAIL.n286 VSUBS 0.033245f
C992 VTAIL.n287 VSUBS 0.032245f
C993 VTAIL.n288 VSUBS 0.017327f
C994 VTAIL.n289 VSUBS 0.040955f
C995 VTAIL.n290 VSUBS 0.018346f
C996 VTAIL.n291 VSUBS 0.032245f
C997 VTAIL.n292 VSUBS 0.017327f
C998 VTAIL.n293 VSUBS 0.040955f
C999 VTAIL.n294 VSUBS 0.018346f
C1000 VTAIL.n295 VSUBS 0.032245f
C1001 VTAIL.n296 VSUBS 0.017327f
C1002 VTAIL.n297 VSUBS 0.040955f
C1003 VTAIL.n298 VSUBS 0.040955f
C1004 VTAIL.n299 VSUBS 0.018346f
C1005 VTAIL.n300 VSUBS 0.032245f
C1006 VTAIL.n301 VSUBS 0.017327f
C1007 VTAIL.n302 VSUBS 0.040955f
C1008 VTAIL.n303 VSUBS 0.018346f
C1009 VTAIL.n304 VSUBS 0.032245f
C1010 VTAIL.n305 VSUBS 0.017327f
C1011 VTAIL.n306 VSUBS 0.040955f
C1012 VTAIL.n307 VSUBS 0.018346f
C1013 VTAIL.n308 VSUBS 0.032245f
C1014 VTAIL.n309 VSUBS 0.017327f
C1015 VTAIL.n310 VSUBS 0.040955f
C1016 VTAIL.n311 VSUBS 0.018346f
C1017 VTAIL.n312 VSUBS 0.032245f
C1018 VTAIL.n313 VSUBS 0.017327f
C1019 VTAIL.n314 VSUBS 0.040955f
C1020 VTAIL.n315 VSUBS 0.018346f
C1021 VTAIL.n316 VSUBS 0.243752f
C1022 VTAIL.t7 VSUBS 0.087814f
C1023 VTAIL.n317 VSUBS 0.030716f
C1024 VTAIL.n318 VSUBS 0.026053f
C1025 VTAIL.n319 VSUBS 0.017327f
C1026 VTAIL.n320 VSUBS 2.31214f
C1027 VTAIL.n321 VSUBS 0.032245f
C1028 VTAIL.n322 VSUBS 0.017327f
C1029 VTAIL.n323 VSUBS 0.018346f
C1030 VTAIL.n324 VSUBS 0.040955f
C1031 VTAIL.n325 VSUBS 0.040955f
C1032 VTAIL.n326 VSUBS 0.018346f
C1033 VTAIL.n327 VSUBS 0.017327f
C1034 VTAIL.n328 VSUBS 0.032245f
C1035 VTAIL.n329 VSUBS 0.032245f
C1036 VTAIL.n330 VSUBS 0.017327f
C1037 VTAIL.n331 VSUBS 0.018346f
C1038 VTAIL.n332 VSUBS 0.040955f
C1039 VTAIL.n333 VSUBS 0.040955f
C1040 VTAIL.n334 VSUBS 0.018346f
C1041 VTAIL.n335 VSUBS 0.017327f
C1042 VTAIL.n336 VSUBS 0.032245f
C1043 VTAIL.n337 VSUBS 0.032245f
C1044 VTAIL.n338 VSUBS 0.017327f
C1045 VTAIL.n339 VSUBS 0.018346f
C1046 VTAIL.n340 VSUBS 0.040955f
C1047 VTAIL.n341 VSUBS 0.040955f
C1048 VTAIL.n342 VSUBS 0.018346f
C1049 VTAIL.n343 VSUBS 0.017327f
C1050 VTAIL.n344 VSUBS 0.032245f
C1051 VTAIL.n345 VSUBS 0.032245f
C1052 VTAIL.n346 VSUBS 0.017327f
C1053 VTAIL.n347 VSUBS 0.018346f
C1054 VTAIL.n348 VSUBS 0.040955f
C1055 VTAIL.n349 VSUBS 0.040955f
C1056 VTAIL.n350 VSUBS 0.018346f
C1057 VTAIL.n351 VSUBS 0.017327f
C1058 VTAIL.n352 VSUBS 0.032245f
C1059 VTAIL.n353 VSUBS 0.032245f
C1060 VTAIL.n354 VSUBS 0.017327f
C1061 VTAIL.n355 VSUBS 0.018346f
C1062 VTAIL.n356 VSUBS 0.040955f
C1063 VTAIL.n357 VSUBS 0.040955f
C1064 VTAIL.n358 VSUBS 0.018346f
C1065 VTAIL.n359 VSUBS 0.017327f
C1066 VTAIL.n360 VSUBS 0.032245f
C1067 VTAIL.n361 VSUBS 0.032245f
C1068 VTAIL.n362 VSUBS 0.017327f
C1069 VTAIL.n363 VSUBS 0.017837f
C1070 VTAIL.n364 VSUBS 0.017837f
C1071 VTAIL.n365 VSUBS 0.040955f
C1072 VTAIL.n366 VSUBS 0.040955f
C1073 VTAIL.n367 VSUBS 0.018346f
C1074 VTAIL.n368 VSUBS 0.017327f
C1075 VTAIL.n369 VSUBS 0.032245f
C1076 VTAIL.n370 VSUBS 0.032245f
C1077 VTAIL.n371 VSUBS 0.017327f
C1078 VTAIL.n372 VSUBS 0.018346f
C1079 VTAIL.n373 VSUBS 0.040955f
C1080 VTAIL.n374 VSUBS 0.091704f
C1081 VTAIL.n375 VSUBS 0.018346f
C1082 VTAIL.n376 VSUBS 0.017327f
C1083 VTAIL.n377 VSUBS 0.071449f
C1084 VTAIL.n378 VSUBS 0.04569f
C1085 VTAIL.n379 VSUBS 2.05366f
C1086 VTAIL.t4 VSUBS 0.426295f
C1087 VTAIL.t6 VSUBS 0.426295f
C1088 VTAIL.n380 VSUBS 3.29536f
C1089 VTAIL.n381 VSUBS 0.890486f
C1090 VTAIL.n382 VSUBS 0.033245f
C1091 VTAIL.n383 VSUBS 0.032245f
C1092 VTAIL.n384 VSUBS 0.017327f
C1093 VTAIL.n385 VSUBS 0.040955f
C1094 VTAIL.n386 VSUBS 0.018346f
C1095 VTAIL.n387 VSUBS 0.032245f
C1096 VTAIL.n388 VSUBS 0.017327f
C1097 VTAIL.n389 VSUBS 0.040955f
C1098 VTAIL.n390 VSUBS 0.018346f
C1099 VTAIL.n391 VSUBS 0.032245f
C1100 VTAIL.n392 VSUBS 0.017327f
C1101 VTAIL.n393 VSUBS 0.040955f
C1102 VTAIL.n394 VSUBS 0.040955f
C1103 VTAIL.n395 VSUBS 0.018346f
C1104 VTAIL.n396 VSUBS 0.032245f
C1105 VTAIL.n397 VSUBS 0.017327f
C1106 VTAIL.n398 VSUBS 0.040955f
C1107 VTAIL.n399 VSUBS 0.018346f
C1108 VTAIL.n400 VSUBS 0.032245f
C1109 VTAIL.n401 VSUBS 0.017327f
C1110 VTAIL.n402 VSUBS 0.040955f
C1111 VTAIL.n403 VSUBS 0.018346f
C1112 VTAIL.n404 VSUBS 0.032245f
C1113 VTAIL.n405 VSUBS 0.017327f
C1114 VTAIL.n406 VSUBS 0.040955f
C1115 VTAIL.n407 VSUBS 0.018346f
C1116 VTAIL.n408 VSUBS 0.032245f
C1117 VTAIL.n409 VSUBS 0.017327f
C1118 VTAIL.n410 VSUBS 0.040955f
C1119 VTAIL.n411 VSUBS 0.018346f
C1120 VTAIL.n412 VSUBS 0.243752f
C1121 VTAIL.t1 VSUBS 0.087814f
C1122 VTAIL.n413 VSUBS 0.030716f
C1123 VTAIL.n414 VSUBS 0.026053f
C1124 VTAIL.n415 VSUBS 0.017327f
C1125 VTAIL.n416 VSUBS 2.31214f
C1126 VTAIL.n417 VSUBS 0.032245f
C1127 VTAIL.n418 VSUBS 0.017327f
C1128 VTAIL.n419 VSUBS 0.018346f
C1129 VTAIL.n420 VSUBS 0.040955f
C1130 VTAIL.n421 VSUBS 0.040955f
C1131 VTAIL.n422 VSUBS 0.018346f
C1132 VTAIL.n423 VSUBS 0.017327f
C1133 VTAIL.n424 VSUBS 0.032245f
C1134 VTAIL.n425 VSUBS 0.032245f
C1135 VTAIL.n426 VSUBS 0.017327f
C1136 VTAIL.n427 VSUBS 0.018346f
C1137 VTAIL.n428 VSUBS 0.040955f
C1138 VTAIL.n429 VSUBS 0.040955f
C1139 VTAIL.n430 VSUBS 0.018346f
C1140 VTAIL.n431 VSUBS 0.017327f
C1141 VTAIL.n432 VSUBS 0.032245f
C1142 VTAIL.n433 VSUBS 0.032245f
C1143 VTAIL.n434 VSUBS 0.017327f
C1144 VTAIL.n435 VSUBS 0.018346f
C1145 VTAIL.n436 VSUBS 0.040955f
C1146 VTAIL.n437 VSUBS 0.040955f
C1147 VTAIL.n438 VSUBS 0.018346f
C1148 VTAIL.n439 VSUBS 0.017327f
C1149 VTAIL.n440 VSUBS 0.032245f
C1150 VTAIL.n441 VSUBS 0.032245f
C1151 VTAIL.n442 VSUBS 0.017327f
C1152 VTAIL.n443 VSUBS 0.018346f
C1153 VTAIL.n444 VSUBS 0.040955f
C1154 VTAIL.n445 VSUBS 0.040955f
C1155 VTAIL.n446 VSUBS 0.018346f
C1156 VTAIL.n447 VSUBS 0.017327f
C1157 VTAIL.n448 VSUBS 0.032245f
C1158 VTAIL.n449 VSUBS 0.032245f
C1159 VTAIL.n450 VSUBS 0.017327f
C1160 VTAIL.n451 VSUBS 0.018346f
C1161 VTAIL.n452 VSUBS 0.040955f
C1162 VTAIL.n453 VSUBS 0.040955f
C1163 VTAIL.n454 VSUBS 0.018346f
C1164 VTAIL.n455 VSUBS 0.017327f
C1165 VTAIL.n456 VSUBS 0.032245f
C1166 VTAIL.n457 VSUBS 0.032245f
C1167 VTAIL.n458 VSUBS 0.017327f
C1168 VTAIL.n459 VSUBS 0.017837f
C1169 VTAIL.n460 VSUBS 0.017837f
C1170 VTAIL.n461 VSUBS 0.040955f
C1171 VTAIL.n462 VSUBS 0.040955f
C1172 VTAIL.n463 VSUBS 0.018346f
C1173 VTAIL.n464 VSUBS 0.017327f
C1174 VTAIL.n465 VSUBS 0.032245f
C1175 VTAIL.n466 VSUBS 0.032245f
C1176 VTAIL.n467 VSUBS 0.017327f
C1177 VTAIL.n468 VSUBS 0.018346f
C1178 VTAIL.n469 VSUBS 0.040955f
C1179 VTAIL.n470 VSUBS 0.091704f
C1180 VTAIL.n471 VSUBS 0.018346f
C1181 VTAIL.n472 VSUBS 0.017327f
C1182 VTAIL.n473 VSUBS 0.071449f
C1183 VTAIL.n474 VSUBS 0.04569f
C1184 VTAIL.n475 VSUBS 0.120296f
C1185 VTAIL.n476 VSUBS 0.033245f
C1186 VTAIL.n477 VSUBS 0.032245f
C1187 VTAIL.n478 VSUBS 0.017327f
C1188 VTAIL.n479 VSUBS 0.040955f
C1189 VTAIL.n480 VSUBS 0.018346f
C1190 VTAIL.n481 VSUBS 0.032245f
C1191 VTAIL.n482 VSUBS 0.017327f
C1192 VTAIL.n483 VSUBS 0.040955f
C1193 VTAIL.n484 VSUBS 0.018346f
C1194 VTAIL.n485 VSUBS 0.032245f
C1195 VTAIL.n486 VSUBS 0.017327f
C1196 VTAIL.n487 VSUBS 0.040955f
C1197 VTAIL.n488 VSUBS 0.040955f
C1198 VTAIL.n489 VSUBS 0.018346f
C1199 VTAIL.n490 VSUBS 0.032245f
C1200 VTAIL.n491 VSUBS 0.017327f
C1201 VTAIL.n492 VSUBS 0.040955f
C1202 VTAIL.n493 VSUBS 0.018346f
C1203 VTAIL.n494 VSUBS 0.032245f
C1204 VTAIL.n495 VSUBS 0.017327f
C1205 VTAIL.n496 VSUBS 0.040955f
C1206 VTAIL.n497 VSUBS 0.018346f
C1207 VTAIL.n498 VSUBS 0.032245f
C1208 VTAIL.n499 VSUBS 0.017327f
C1209 VTAIL.n500 VSUBS 0.040955f
C1210 VTAIL.n501 VSUBS 0.018346f
C1211 VTAIL.n502 VSUBS 0.032245f
C1212 VTAIL.n503 VSUBS 0.017327f
C1213 VTAIL.n504 VSUBS 0.040955f
C1214 VTAIL.n505 VSUBS 0.018346f
C1215 VTAIL.n506 VSUBS 0.243752f
C1216 VTAIL.t13 VSUBS 0.087814f
C1217 VTAIL.n507 VSUBS 0.030716f
C1218 VTAIL.n508 VSUBS 0.026053f
C1219 VTAIL.n509 VSUBS 0.017327f
C1220 VTAIL.n510 VSUBS 2.31214f
C1221 VTAIL.n511 VSUBS 0.032245f
C1222 VTAIL.n512 VSUBS 0.017327f
C1223 VTAIL.n513 VSUBS 0.018346f
C1224 VTAIL.n514 VSUBS 0.040955f
C1225 VTAIL.n515 VSUBS 0.040955f
C1226 VTAIL.n516 VSUBS 0.018346f
C1227 VTAIL.n517 VSUBS 0.017327f
C1228 VTAIL.n518 VSUBS 0.032245f
C1229 VTAIL.n519 VSUBS 0.032245f
C1230 VTAIL.n520 VSUBS 0.017327f
C1231 VTAIL.n521 VSUBS 0.018346f
C1232 VTAIL.n522 VSUBS 0.040955f
C1233 VTAIL.n523 VSUBS 0.040955f
C1234 VTAIL.n524 VSUBS 0.018346f
C1235 VTAIL.n525 VSUBS 0.017327f
C1236 VTAIL.n526 VSUBS 0.032245f
C1237 VTAIL.n527 VSUBS 0.032245f
C1238 VTAIL.n528 VSUBS 0.017327f
C1239 VTAIL.n529 VSUBS 0.018346f
C1240 VTAIL.n530 VSUBS 0.040955f
C1241 VTAIL.n531 VSUBS 0.040955f
C1242 VTAIL.n532 VSUBS 0.018346f
C1243 VTAIL.n533 VSUBS 0.017327f
C1244 VTAIL.n534 VSUBS 0.032245f
C1245 VTAIL.n535 VSUBS 0.032245f
C1246 VTAIL.n536 VSUBS 0.017327f
C1247 VTAIL.n537 VSUBS 0.018346f
C1248 VTAIL.n538 VSUBS 0.040955f
C1249 VTAIL.n539 VSUBS 0.040955f
C1250 VTAIL.n540 VSUBS 0.018346f
C1251 VTAIL.n541 VSUBS 0.017327f
C1252 VTAIL.n542 VSUBS 0.032245f
C1253 VTAIL.n543 VSUBS 0.032245f
C1254 VTAIL.n544 VSUBS 0.017327f
C1255 VTAIL.n545 VSUBS 0.018346f
C1256 VTAIL.n546 VSUBS 0.040955f
C1257 VTAIL.n547 VSUBS 0.040955f
C1258 VTAIL.n548 VSUBS 0.018346f
C1259 VTAIL.n549 VSUBS 0.017327f
C1260 VTAIL.n550 VSUBS 0.032245f
C1261 VTAIL.n551 VSUBS 0.032245f
C1262 VTAIL.n552 VSUBS 0.017327f
C1263 VTAIL.n553 VSUBS 0.017837f
C1264 VTAIL.n554 VSUBS 0.017837f
C1265 VTAIL.n555 VSUBS 0.040955f
C1266 VTAIL.n556 VSUBS 0.040955f
C1267 VTAIL.n557 VSUBS 0.018346f
C1268 VTAIL.n558 VSUBS 0.017327f
C1269 VTAIL.n559 VSUBS 0.032245f
C1270 VTAIL.n560 VSUBS 0.032245f
C1271 VTAIL.n561 VSUBS 0.017327f
C1272 VTAIL.n562 VSUBS 0.018346f
C1273 VTAIL.n563 VSUBS 0.040955f
C1274 VTAIL.n564 VSUBS 0.091704f
C1275 VTAIL.n565 VSUBS 0.018346f
C1276 VTAIL.n566 VSUBS 0.017327f
C1277 VTAIL.n567 VSUBS 0.071449f
C1278 VTAIL.n568 VSUBS 0.04569f
C1279 VTAIL.n569 VSUBS 0.120296f
C1280 VTAIL.t12 VSUBS 0.426295f
C1281 VTAIL.t11 VSUBS 0.426295f
C1282 VTAIL.n570 VSUBS 3.29536f
C1283 VTAIL.n571 VSUBS 0.890486f
C1284 VTAIL.n572 VSUBS 0.033245f
C1285 VTAIL.n573 VSUBS 0.032245f
C1286 VTAIL.n574 VSUBS 0.017327f
C1287 VTAIL.n575 VSUBS 0.040955f
C1288 VTAIL.n576 VSUBS 0.018346f
C1289 VTAIL.n577 VSUBS 0.032245f
C1290 VTAIL.n578 VSUBS 0.017327f
C1291 VTAIL.n579 VSUBS 0.040955f
C1292 VTAIL.n580 VSUBS 0.018346f
C1293 VTAIL.n581 VSUBS 0.032245f
C1294 VTAIL.n582 VSUBS 0.017327f
C1295 VTAIL.n583 VSUBS 0.040955f
C1296 VTAIL.n584 VSUBS 0.040955f
C1297 VTAIL.n585 VSUBS 0.018346f
C1298 VTAIL.n586 VSUBS 0.032245f
C1299 VTAIL.n587 VSUBS 0.017327f
C1300 VTAIL.n588 VSUBS 0.040955f
C1301 VTAIL.n589 VSUBS 0.018346f
C1302 VTAIL.n590 VSUBS 0.032245f
C1303 VTAIL.n591 VSUBS 0.017327f
C1304 VTAIL.n592 VSUBS 0.040955f
C1305 VTAIL.n593 VSUBS 0.018346f
C1306 VTAIL.n594 VSUBS 0.032245f
C1307 VTAIL.n595 VSUBS 0.017327f
C1308 VTAIL.n596 VSUBS 0.040955f
C1309 VTAIL.n597 VSUBS 0.018346f
C1310 VTAIL.n598 VSUBS 0.032245f
C1311 VTAIL.n599 VSUBS 0.017327f
C1312 VTAIL.n600 VSUBS 0.040955f
C1313 VTAIL.n601 VSUBS 0.018346f
C1314 VTAIL.n602 VSUBS 0.243752f
C1315 VTAIL.t9 VSUBS 0.087814f
C1316 VTAIL.n603 VSUBS 0.030716f
C1317 VTAIL.n604 VSUBS 0.026053f
C1318 VTAIL.n605 VSUBS 0.017327f
C1319 VTAIL.n606 VSUBS 2.31214f
C1320 VTAIL.n607 VSUBS 0.032245f
C1321 VTAIL.n608 VSUBS 0.017327f
C1322 VTAIL.n609 VSUBS 0.018346f
C1323 VTAIL.n610 VSUBS 0.040955f
C1324 VTAIL.n611 VSUBS 0.040955f
C1325 VTAIL.n612 VSUBS 0.018346f
C1326 VTAIL.n613 VSUBS 0.017327f
C1327 VTAIL.n614 VSUBS 0.032245f
C1328 VTAIL.n615 VSUBS 0.032245f
C1329 VTAIL.n616 VSUBS 0.017327f
C1330 VTAIL.n617 VSUBS 0.018346f
C1331 VTAIL.n618 VSUBS 0.040955f
C1332 VTAIL.n619 VSUBS 0.040955f
C1333 VTAIL.n620 VSUBS 0.018346f
C1334 VTAIL.n621 VSUBS 0.017327f
C1335 VTAIL.n622 VSUBS 0.032245f
C1336 VTAIL.n623 VSUBS 0.032245f
C1337 VTAIL.n624 VSUBS 0.017327f
C1338 VTAIL.n625 VSUBS 0.018346f
C1339 VTAIL.n626 VSUBS 0.040955f
C1340 VTAIL.n627 VSUBS 0.040955f
C1341 VTAIL.n628 VSUBS 0.018346f
C1342 VTAIL.n629 VSUBS 0.017327f
C1343 VTAIL.n630 VSUBS 0.032245f
C1344 VTAIL.n631 VSUBS 0.032245f
C1345 VTAIL.n632 VSUBS 0.017327f
C1346 VTAIL.n633 VSUBS 0.018346f
C1347 VTAIL.n634 VSUBS 0.040955f
C1348 VTAIL.n635 VSUBS 0.040955f
C1349 VTAIL.n636 VSUBS 0.018346f
C1350 VTAIL.n637 VSUBS 0.017327f
C1351 VTAIL.n638 VSUBS 0.032245f
C1352 VTAIL.n639 VSUBS 0.032245f
C1353 VTAIL.n640 VSUBS 0.017327f
C1354 VTAIL.n641 VSUBS 0.018346f
C1355 VTAIL.n642 VSUBS 0.040955f
C1356 VTAIL.n643 VSUBS 0.040955f
C1357 VTAIL.n644 VSUBS 0.018346f
C1358 VTAIL.n645 VSUBS 0.017327f
C1359 VTAIL.n646 VSUBS 0.032245f
C1360 VTAIL.n647 VSUBS 0.032245f
C1361 VTAIL.n648 VSUBS 0.017327f
C1362 VTAIL.n649 VSUBS 0.017837f
C1363 VTAIL.n650 VSUBS 0.017837f
C1364 VTAIL.n651 VSUBS 0.040955f
C1365 VTAIL.n652 VSUBS 0.040955f
C1366 VTAIL.n653 VSUBS 0.018346f
C1367 VTAIL.n654 VSUBS 0.017327f
C1368 VTAIL.n655 VSUBS 0.032245f
C1369 VTAIL.n656 VSUBS 0.032245f
C1370 VTAIL.n657 VSUBS 0.017327f
C1371 VTAIL.n658 VSUBS 0.018346f
C1372 VTAIL.n659 VSUBS 0.040955f
C1373 VTAIL.n660 VSUBS 0.091704f
C1374 VTAIL.n661 VSUBS 0.018346f
C1375 VTAIL.n662 VSUBS 0.017327f
C1376 VTAIL.n663 VSUBS 0.071449f
C1377 VTAIL.n664 VSUBS 0.04569f
C1378 VTAIL.n665 VSUBS 2.05366f
C1379 VTAIL.n666 VSUBS 0.033245f
C1380 VTAIL.n667 VSUBS 0.032245f
C1381 VTAIL.n668 VSUBS 0.017327f
C1382 VTAIL.n669 VSUBS 0.040955f
C1383 VTAIL.n670 VSUBS 0.018346f
C1384 VTAIL.n671 VSUBS 0.032245f
C1385 VTAIL.n672 VSUBS 0.017327f
C1386 VTAIL.n673 VSUBS 0.040955f
C1387 VTAIL.n674 VSUBS 0.018346f
C1388 VTAIL.n675 VSUBS 0.032245f
C1389 VTAIL.n676 VSUBS 0.017327f
C1390 VTAIL.n677 VSUBS 0.040955f
C1391 VTAIL.n678 VSUBS 0.018346f
C1392 VTAIL.n679 VSUBS 0.032245f
C1393 VTAIL.n680 VSUBS 0.017327f
C1394 VTAIL.n681 VSUBS 0.040955f
C1395 VTAIL.n682 VSUBS 0.018346f
C1396 VTAIL.n683 VSUBS 0.032245f
C1397 VTAIL.n684 VSUBS 0.017327f
C1398 VTAIL.n685 VSUBS 0.040955f
C1399 VTAIL.n686 VSUBS 0.018346f
C1400 VTAIL.n687 VSUBS 0.032245f
C1401 VTAIL.n688 VSUBS 0.017327f
C1402 VTAIL.n689 VSUBS 0.040955f
C1403 VTAIL.n690 VSUBS 0.018346f
C1404 VTAIL.n691 VSUBS 0.032245f
C1405 VTAIL.n692 VSUBS 0.017327f
C1406 VTAIL.n693 VSUBS 0.040955f
C1407 VTAIL.n694 VSUBS 0.018346f
C1408 VTAIL.n695 VSUBS 0.243752f
C1409 VTAIL.t5 VSUBS 0.087814f
C1410 VTAIL.n696 VSUBS 0.030716f
C1411 VTAIL.n697 VSUBS 0.026053f
C1412 VTAIL.n698 VSUBS 0.017327f
C1413 VTAIL.n699 VSUBS 2.31214f
C1414 VTAIL.n700 VSUBS 0.032245f
C1415 VTAIL.n701 VSUBS 0.017327f
C1416 VTAIL.n702 VSUBS 0.018346f
C1417 VTAIL.n703 VSUBS 0.040955f
C1418 VTAIL.n704 VSUBS 0.040955f
C1419 VTAIL.n705 VSUBS 0.018346f
C1420 VTAIL.n706 VSUBS 0.017327f
C1421 VTAIL.n707 VSUBS 0.032245f
C1422 VTAIL.n708 VSUBS 0.032245f
C1423 VTAIL.n709 VSUBS 0.017327f
C1424 VTAIL.n710 VSUBS 0.018346f
C1425 VTAIL.n711 VSUBS 0.040955f
C1426 VTAIL.n712 VSUBS 0.040955f
C1427 VTAIL.n713 VSUBS 0.018346f
C1428 VTAIL.n714 VSUBS 0.017327f
C1429 VTAIL.n715 VSUBS 0.032245f
C1430 VTAIL.n716 VSUBS 0.032245f
C1431 VTAIL.n717 VSUBS 0.017327f
C1432 VTAIL.n718 VSUBS 0.018346f
C1433 VTAIL.n719 VSUBS 0.040955f
C1434 VTAIL.n720 VSUBS 0.040955f
C1435 VTAIL.n721 VSUBS 0.018346f
C1436 VTAIL.n722 VSUBS 0.017327f
C1437 VTAIL.n723 VSUBS 0.032245f
C1438 VTAIL.n724 VSUBS 0.032245f
C1439 VTAIL.n725 VSUBS 0.017327f
C1440 VTAIL.n726 VSUBS 0.018346f
C1441 VTAIL.n727 VSUBS 0.040955f
C1442 VTAIL.n728 VSUBS 0.040955f
C1443 VTAIL.n729 VSUBS 0.018346f
C1444 VTAIL.n730 VSUBS 0.017327f
C1445 VTAIL.n731 VSUBS 0.032245f
C1446 VTAIL.n732 VSUBS 0.032245f
C1447 VTAIL.n733 VSUBS 0.017327f
C1448 VTAIL.n734 VSUBS 0.018346f
C1449 VTAIL.n735 VSUBS 0.040955f
C1450 VTAIL.n736 VSUBS 0.040955f
C1451 VTAIL.n737 VSUBS 0.040955f
C1452 VTAIL.n738 VSUBS 0.018346f
C1453 VTAIL.n739 VSUBS 0.017327f
C1454 VTAIL.n740 VSUBS 0.032245f
C1455 VTAIL.n741 VSUBS 0.032245f
C1456 VTAIL.n742 VSUBS 0.017327f
C1457 VTAIL.n743 VSUBS 0.017837f
C1458 VTAIL.n744 VSUBS 0.017837f
C1459 VTAIL.n745 VSUBS 0.040955f
C1460 VTAIL.n746 VSUBS 0.040955f
C1461 VTAIL.n747 VSUBS 0.018346f
C1462 VTAIL.n748 VSUBS 0.017327f
C1463 VTAIL.n749 VSUBS 0.032245f
C1464 VTAIL.n750 VSUBS 0.032245f
C1465 VTAIL.n751 VSUBS 0.017327f
C1466 VTAIL.n752 VSUBS 0.018346f
C1467 VTAIL.n753 VSUBS 0.040955f
C1468 VTAIL.n754 VSUBS 0.091704f
C1469 VTAIL.n755 VSUBS 0.018346f
C1470 VTAIL.n756 VSUBS 0.017327f
C1471 VTAIL.n757 VSUBS 0.071449f
C1472 VTAIL.n758 VSUBS 0.04569f
C1473 VTAIL.n759 VSUBS 2.04762f
C1474 VDD1.t3 VSUBS 0.522234f
C1475 VDD1.t2 VSUBS 0.522234f
C1476 VDD1.n0 VSUBS 4.29192f
C1477 VDD1.t7 VSUBS 0.522234f
C1478 VDD1.t5 VSUBS 0.522234f
C1479 VDD1.n1 VSUBS 4.290411f
C1480 VDD1.t6 VSUBS 0.522234f
C1481 VDD1.t4 VSUBS 0.522234f
C1482 VDD1.n2 VSUBS 4.290411f
C1483 VDD1.n3 VSUBS 4.40626f
C1484 VDD1.t0 VSUBS 0.522234f
C1485 VDD1.t1 VSUBS 0.522234f
C1486 VDD1.n4 VSUBS 4.28828f
C1487 VDD1.n5 VSUBS 4.41391f
C1488 VP.n0 VSUBS 0.075502f
C1489 VP.t0 VSUBS 0.641124f
C1490 VP.t1 VSUBS 0.641124f
C1491 VP.t5 VSUBS 0.645063f
C1492 VP.n1 VSUBS 0.16068f
C1493 VP.t4 VSUBS 0.641124f
C1494 VP.t3 VSUBS 0.641124f
C1495 VP.t2 VSUBS 0.645063f
C1496 VP.n2 VSUBS 0.271415f
C1497 VP.n3 VSUBS 0.252302f
C1498 VP.n4 VSUBS 0.025512f
C1499 VP.n5 VSUBS 0.252302f
C1500 VP.t6 VSUBS 0.645063f
C1501 VP.n6 VSUBS 0.271315f
C1502 VP.n7 VSUBS 3.26267f
C1503 VP.n8 VSUBS 3.32553f
C1504 VP.n9 VSUBS 0.271315f
C1505 VP.n10 VSUBS 0.252302f
C1506 VP.n11 VSUBS 0.025512f
C1507 VP.n12 VSUBS 0.252302f
C1508 VP.t7 VSUBS 0.645063f
C1509 VP.n13 VSUBS 0.271315f
C1510 VP.n14 VSUBS 0.058511f
.ends

