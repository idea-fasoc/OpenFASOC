* NGSPICE file created from diff_pair_sample_1651.ext - technology: sky130A

.subckt diff_pair_sample_1651 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t19 VP.t0 VDD1.t5 w_n5926_n2380# sky130_fd_pr__pfet_01v8 ad=1.1649 pd=7.39 as=1.1649 ps=7.39 w=7.06 l=3.8
X1 VDD1.t7 VP.t1 VTAIL.t18 w_n5926_n2380# sky130_fd_pr__pfet_01v8 ad=2.7534 pd=14.9 as=1.1649 ps=7.39 w=7.06 l=3.8
X2 B.t11 B.t9 B.t10 w_n5926_n2380# sky130_fd_pr__pfet_01v8 ad=2.7534 pd=14.9 as=0 ps=0 w=7.06 l=3.8
X3 VTAIL.t5 VN.t0 VDD2.t9 w_n5926_n2380# sky130_fd_pr__pfet_01v8 ad=1.1649 pd=7.39 as=1.1649 ps=7.39 w=7.06 l=3.8
X4 VDD2.t8 VN.t1 VTAIL.t4 w_n5926_n2380# sky130_fd_pr__pfet_01v8 ad=2.7534 pd=14.9 as=1.1649 ps=7.39 w=7.06 l=3.8
X5 VTAIL.t17 VP.t2 VDD1.t9 w_n5926_n2380# sky130_fd_pr__pfet_01v8 ad=1.1649 pd=7.39 as=1.1649 ps=7.39 w=7.06 l=3.8
X6 VDD1.t2 VP.t3 VTAIL.t16 w_n5926_n2380# sky130_fd_pr__pfet_01v8 ad=1.1649 pd=7.39 as=1.1649 ps=7.39 w=7.06 l=3.8
X7 B.t8 B.t6 B.t7 w_n5926_n2380# sky130_fd_pr__pfet_01v8 ad=2.7534 pd=14.9 as=0 ps=0 w=7.06 l=3.8
X8 VDD2.t7 VN.t2 VTAIL.t8 w_n5926_n2380# sky130_fd_pr__pfet_01v8 ad=1.1649 pd=7.39 as=2.7534 ps=14.9 w=7.06 l=3.8
X9 VTAIL.t9 VN.t3 VDD2.t6 w_n5926_n2380# sky130_fd_pr__pfet_01v8 ad=1.1649 pd=7.39 as=1.1649 ps=7.39 w=7.06 l=3.8
X10 B.t5 B.t3 B.t4 w_n5926_n2380# sky130_fd_pr__pfet_01v8 ad=2.7534 pd=14.9 as=0 ps=0 w=7.06 l=3.8
X11 VDD2.t5 VN.t4 VTAIL.t7 w_n5926_n2380# sky130_fd_pr__pfet_01v8 ad=1.1649 pd=7.39 as=1.1649 ps=7.39 w=7.06 l=3.8
X12 B.t2 B.t0 B.t1 w_n5926_n2380# sky130_fd_pr__pfet_01v8 ad=2.7534 pd=14.9 as=0 ps=0 w=7.06 l=3.8
X13 VTAIL.t15 VP.t4 VDD1.t6 w_n5926_n2380# sky130_fd_pr__pfet_01v8 ad=1.1649 pd=7.39 as=1.1649 ps=7.39 w=7.06 l=3.8
X14 VDD2.t4 VN.t5 VTAIL.t3 w_n5926_n2380# sky130_fd_pr__pfet_01v8 ad=1.1649 pd=7.39 as=2.7534 ps=14.9 w=7.06 l=3.8
X15 VDD1.t3 VP.t5 VTAIL.t14 w_n5926_n2380# sky130_fd_pr__pfet_01v8 ad=1.1649 pd=7.39 as=2.7534 ps=14.9 w=7.06 l=3.8
X16 VTAIL.t13 VP.t6 VDD1.t0 w_n5926_n2380# sky130_fd_pr__pfet_01v8 ad=1.1649 pd=7.39 as=1.1649 ps=7.39 w=7.06 l=3.8
X17 VDD2.t3 VN.t6 VTAIL.t6 w_n5926_n2380# sky130_fd_pr__pfet_01v8 ad=2.7534 pd=14.9 as=1.1649 ps=7.39 w=7.06 l=3.8
X18 VTAIL.t1 VN.t7 VDD2.t2 w_n5926_n2380# sky130_fd_pr__pfet_01v8 ad=1.1649 pd=7.39 as=1.1649 ps=7.39 w=7.06 l=3.8
X19 VDD1.t1 VP.t7 VTAIL.t12 w_n5926_n2380# sky130_fd_pr__pfet_01v8 ad=1.1649 pd=7.39 as=1.1649 ps=7.39 w=7.06 l=3.8
X20 VDD1.t8 VP.t8 VTAIL.t11 w_n5926_n2380# sky130_fd_pr__pfet_01v8 ad=1.1649 pd=7.39 as=2.7534 ps=14.9 w=7.06 l=3.8
X21 VDD1.t4 VP.t9 VTAIL.t10 w_n5926_n2380# sky130_fd_pr__pfet_01v8 ad=2.7534 pd=14.9 as=1.1649 ps=7.39 w=7.06 l=3.8
X22 VTAIL.t0 VN.t8 VDD2.t1 w_n5926_n2380# sky130_fd_pr__pfet_01v8 ad=1.1649 pd=7.39 as=1.1649 ps=7.39 w=7.06 l=3.8
X23 VDD2.t0 VN.t9 VTAIL.t2 w_n5926_n2380# sky130_fd_pr__pfet_01v8 ad=1.1649 pd=7.39 as=1.1649 ps=7.39 w=7.06 l=3.8
R0 VP.n34 VP.n33 161.3
R1 VP.n35 VP.n30 161.3
R2 VP.n37 VP.n36 161.3
R3 VP.n38 VP.n29 161.3
R4 VP.n40 VP.n39 161.3
R5 VP.n41 VP.n28 161.3
R6 VP.n43 VP.n42 161.3
R7 VP.n44 VP.n27 161.3
R8 VP.n47 VP.n46 161.3
R9 VP.n48 VP.n26 161.3
R10 VP.n50 VP.n49 161.3
R11 VP.n51 VP.n25 161.3
R12 VP.n53 VP.n52 161.3
R13 VP.n54 VP.n24 161.3
R14 VP.n56 VP.n55 161.3
R15 VP.n57 VP.n23 161.3
R16 VP.n60 VP.n59 161.3
R17 VP.n61 VP.n22 161.3
R18 VP.n63 VP.n62 161.3
R19 VP.n64 VP.n21 161.3
R20 VP.n66 VP.n65 161.3
R21 VP.n67 VP.n20 161.3
R22 VP.n69 VP.n68 161.3
R23 VP.n70 VP.n19 161.3
R24 VP.n72 VP.n71 161.3
R25 VP.n129 VP.n128 161.3
R26 VP.n127 VP.n1 161.3
R27 VP.n126 VP.n125 161.3
R28 VP.n124 VP.n2 161.3
R29 VP.n123 VP.n122 161.3
R30 VP.n121 VP.n3 161.3
R31 VP.n120 VP.n119 161.3
R32 VP.n118 VP.n4 161.3
R33 VP.n117 VP.n116 161.3
R34 VP.n114 VP.n5 161.3
R35 VP.n113 VP.n112 161.3
R36 VP.n111 VP.n6 161.3
R37 VP.n110 VP.n109 161.3
R38 VP.n108 VP.n7 161.3
R39 VP.n107 VP.n106 161.3
R40 VP.n105 VP.n8 161.3
R41 VP.n104 VP.n103 161.3
R42 VP.n101 VP.n9 161.3
R43 VP.n100 VP.n99 161.3
R44 VP.n98 VP.n10 161.3
R45 VP.n97 VP.n96 161.3
R46 VP.n95 VP.n11 161.3
R47 VP.n94 VP.n93 161.3
R48 VP.n92 VP.n12 161.3
R49 VP.n91 VP.n90 161.3
R50 VP.n88 VP.n13 161.3
R51 VP.n87 VP.n86 161.3
R52 VP.n85 VP.n14 161.3
R53 VP.n84 VP.n83 161.3
R54 VP.n82 VP.n15 161.3
R55 VP.n81 VP.n80 161.3
R56 VP.n79 VP.n16 161.3
R57 VP.n78 VP.n77 161.3
R58 VP.n76 VP.n17 161.3
R59 VP.n75 VP.n74 89.7537
R60 VP.n130 VP.n0 89.7537
R61 VP.n73 VP.n18 89.7537
R62 VP.n31 VP.t9 77.0547
R63 VP.n32 VP.n31 56.597
R64 VP.n96 VP.n95 56.5617
R65 VP.n109 VP.n108 56.5617
R66 VP.n52 VP.n51 56.5617
R67 VP.n39 VP.n38 56.5617
R68 VP.n74 VP.n73 55.9124
R69 VP.n83 VP.n82 45.9053
R70 VP.n122 VP.n121 45.9053
R71 VP.n65 VP.n64 45.9053
R72 VP.n75 VP.t1 44.7758
R73 VP.n89 VP.t2 44.7758
R74 VP.n102 VP.t3 44.7758
R75 VP.n115 VP.t6 44.7758
R76 VP.n0 VP.t5 44.7758
R77 VP.n18 VP.t8 44.7758
R78 VP.n58 VP.t4 44.7758
R79 VP.n45 VP.t7 44.7758
R80 VP.n32 VP.t0 44.7758
R81 VP.n82 VP.n81 35.2488
R82 VP.n122 VP.n2 35.2488
R83 VP.n65 VP.n20 35.2488
R84 VP.n77 VP.n76 24.5923
R85 VP.n77 VP.n16 24.5923
R86 VP.n81 VP.n16 24.5923
R87 VP.n83 VP.n14 24.5923
R88 VP.n87 VP.n14 24.5923
R89 VP.n88 VP.n87 24.5923
R90 VP.n90 VP.n12 24.5923
R91 VP.n94 VP.n12 24.5923
R92 VP.n95 VP.n94 24.5923
R93 VP.n96 VP.n10 24.5923
R94 VP.n100 VP.n10 24.5923
R95 VP.n101 VP.n100 24.5923
R96 VP.n103 VP.n8 24.5923
R97 VP.n107 VP.n8 24.5923
R98 VP.n108 VP.n107 24.5923
R99 VP.n109 VP.n6 24.5923
R100 VP.n113 VP.n6 24.5923
R101 VP.n114 VP.n113 24.5923
R102 VP.n116 VP.n4 24.5923
R103 VP.n120 VP.n4 24.5923
R104 VP.n121 VP.n120 24.5923
R105 VP.n126 VP.n2 24.5923
R106 VP.n127 VP.n126 24.5923
R107 VP.n128 VP.n127 24.5923
R108 VP.n69 VP.n20 24.5923
R109 VP.n70 VP.n69 24.5923
R110 VP.n71 VP.n70 24.5923
R111 VP.n52 VP.n24 24.5923
R112 VP.n56 VP.n24 24.5923
R113 VP.n57 VP.n56 24.5923
R114 VP.n59 VP.n22 24.5923
R115 VP.n63 VP.n22 24.5923
R116 VP.n64 VP.n63 24.5923
R117 VP.n39 VP.n28 24.5923
R118 VP.n43 VP.n28 24.5923
R119 VP.n44 VP.n43 24.5923
R120 VP.n46 VP.n26 24.5923
R121 VP.n50 VP.n26 24.5923
R122 VP.n51 VP.n50 24.5923
R123 VP.n33 VP.n30 24.5923
R124 VP.n37 VP.n30 24.5923
R125 VP.n38 VP.n37 24.5923
R126 VP.n90 VP.n89 18.6903
R127 VP.n115 VP.n114 18.6903
R128 VP.n58 VP.n57 18.6903
R129 VP.n33 VP.n32 18.6903
R130 VP.n102 VP.n101 12.2964
R131 VP.n103 VP.n102 12.2964
R132 VP.n45 VP.n44 12.2964
R133 VP.n46 VP.n45 12.2964
R134 VP.n89 VP.n88 5.90254
R135 VP.n116 VP.n115 5.90254
R136 VP.n59 VP.n58 5.90254
R137 VP.n34 VP.n31 2.50625
R138 VP.n76 VP.n75 0.492337
R139 VP.n128 VP.n0 0.492337
R140 VP.n71 VP.n18 0.492337
R141 VP.n73 VP.n72 0.354861
R142 VP.n74 VP.n17 0.354861
R143 VP.n130 VP.n129 0.354861
R144 VP VP.n130 0.267071
R145 VP.n35 VP.n34 0.189894
R146 VP.n36 VP.n35 0.189894
R147 VP.n36 VP.n29 0.189894
R148 VP.n40 VP.n29 0.189894
R149 VP.n41 VP.n40 0.189894
R150 VP.n42 VP.n41 0.189894
R151 VP.n42 VP.n27 0.189894
R152 VP.n47 VP.n27 0.189894
R153 VP.n48 VP.n47 0.189894
R154 VP.n49 VP.n48 0.189894
R155 VP.n49 VP.n25 0.189894
R156 VP.n53 VP.n25 0.189894
R157 VP.n54 VP.n53 0.189894
R158 VP.n55 VP.n54 0.189894
R159 VP.n55 VP.n23 0.189894
R160 VP.n60 VP.n23 0.189894
R161 VP.n61 VP.n60 0.189894
R162 VP.n62 VP.n61 0.189894
R163 VP.n62 VP.n21 0.189894
R164 VP.n66 VP.n21 0.189894
R165 VP.n67 VP.n66 0.189894
R166 VP.n68 VP.n67 0.189894
R167 VP.n68 VP.n19 0.189894
R168 VP.n72 VP.n19 0.189894
R169 VP.n78 VP.n17 0.189894
R170 VP.n79 VP.n78 0.189894
R171 VP.n80 VP.n79 0.189894
R172 VP.n80 VP.n15 0.189894
R173 VP.n84 VP.n15 0.189894
R174 VP.n85 VP.n84 0.189894
R175 VP.n86 VP.n85 0.189894
R176 VP.n86 VP.n13 0.189894
R177 VP.n91 VP.n13 0.189894
R178 VP.n92 VP.n91 0.189894
R179 VP.n93 VP.n92 0.189894
R180 VP.n93 VP.n11 0.189894
R181 VP.n97 VP.n11 0.189894
R182 VP.n98 VP.n97 0.189894
R183 VP.n99 VP.n98 0.189894
R184 VP.n99 VP.n9 0.189894
R185 VP.n104 VP.n9 0.189894
R186 VP.n105 VP.n104 0.189894
R187 VP.n106 VP.n105 0.189894
R188 VP.n106 VP.n7 0.189894
R189 VP.n110 VP.n7 0.189894
R190 VP.n111 VP.n110 0.189894
R191 VP.n112 VP.n111 0.189894
R192 VP.n112 VP.n5 0.189894
R193 VP.n117 VP.n5 0.189894
R194 VP.n118 VP.n117 0.189894
R195 VP.n119 VP.n118 0.189894
R196 VP.n119 VP.n3 0.189894
R197 VP.n123 VP.n3 0.189894
R198 VP.n124 VP.n123 0.189894
R199 VP.n125 VP.n124 0.189894
R200 VP.n125 VP.n1 0.189894
R201 VP.n129 VP.n1 0.189894
R202 VDD1.n1 VDD1.t4 94.5427
R203 VDD1.n3 VDD1.t7 94.5425
R204 VDD1.n5 VDD1.n4 88.9931
R205 VDD1.n1 VDD1.n0 86.3782
R206 VDD1.n3 VDD1.n2 86.3782
R207 VDD1.n7 VDD1.n6 86.3781
R208 VDD1.n7 VDD1.n5 49.0763
R209 VDD1.n6 VDD1.t6 4.60461
R210 VDD1.n6 VDD1.t8 4.60461
R211 VDD1.n0 VDD1.t5 4.60461
R212 VDD1.n0 VDD1.t1 4.60461
R213 VDD1.n4 VDD1.t0 4.60461
R214 VDD1.n4 VDD1.t3 4.60461
R215 VDD1.n2 VDD1.t9 4.60461
R216 VDD1.n2 VDD1.t2 4.60461
R217 VDD1 VDD1.n7 2.61257
R218 VDD1 VDD1.n1 0.948776
R219 VDD1.n5 VDD1.n3 0.83524
R220 VTAIL.n11 VTAIL.t8 74.3036
R221 VTAIL.n17 VTAIL.t3 74.3033
R222 VTAIL.n2 VTAIL.t14 74.3033
R223 VTAIL.n16 VTAIL.t11 74.3033
R224 VTAIL.n15 VTAIL.n14 69.6995
R225 VTAIL.n13 VTAIL.n12 69.6995
R226 VTAIL.n10 VTAIL.n9 69.6995
R227 VTAIL.n8 VTAIL.n7 69.6995
R228 VTAIL.n19 VTAIL.n18 69.6994
R229 VTAIL.n1 VTAIL.n0 69.6994
R230 VTAIL.n4 VTAIL.n3 69.6994
R231 VTAIL.n6 VTAIL.n5 69.6994
R232 VTAIL.n8 VTAIL.n6 25.5738
R233 VTAIL.n17 VTAIL.n16 22.0134
R234 VTAIL.n18 VTAIL.t2 4.60461
R235 VTAIL.n18 VTAIL.t1 4.60461
R236 VTAIL.n0 VTAIL.t4 4.60461
R237 VTAIL.n0 VTAIL.t5 4.60461
R238 VTAIL.n3 VTAIL.t16 4.60461
R239 VTAIL.n3 VTAIL.t13 4.60461
R240 VTAIL.n5 VTAIL.t18 4.60461
R241 VTAIL.n5 VTAIL.t17 4.60461
R242 VTAIL.n14 VTAIL.t12 4.60461
R243 VTAIL.n14 VTAIL.t15 4.60461
R244 VTAIL.n12 VTAIL.t10 4.60461
R245 VTAIL.n12 VTAIL.t19 4.60461
R246 VTAIL.n9 VTAIL.t7 4.60461
R247 VTAIL.n9 VTAIL.t9 4.60461
R248 VTAIL.n7 VTAIL.t6 4.60461
R249 VTAIL.n7 VTAIL.t0 4.60461
R250 VTAIL.n10 VTAIL.n8 3.56084
R251 VTAIL.n11 VTAIL.n10 3.56084
R252 VTAIL.n15 VTAIL.n13 3.56084
R253 VTAIL.n16 VTAIL.n15 3.56084
R254 VTAIL.n6 VTAIL.n4 3.56084
R255 VTAIL.n4 VTAIL.n2 3.56084
R256 VTAIL.n19 VTAIL.n17 3.56084
R257 VTAIL VTAIL.n1 2.72895
R258 VTAIL.n13 VTAIL.n11 2.2505
R259 VTAIL.n2 VTAIL.n1 2.2505
R260 VTAIL VTAIL.n19 0.832397
R261 B.n700 B.n699 585
R262 B.n701 B.n78 585
R263 B.n703 B.n702 585
R264 B.n704 B.n77 585
R265 B.n706 B.n705 585
R266 B.n707 B.n76 585
R267 B.n709 B.n708 585
R268 B.n710 B.n75 585
R269 B.n712 B.n711 585
R270 B.n713 B.n74 585
R271 B.n715 B.n714 585
R272 B.n716 B.n73 585
R273 B.n718 B.n717 585
R274 B.n719 B.n72 585
R275 B.n721 B.n720 585
R276 B.n722 B.n71 585
R277 B.n724 B.n723 585
R278 B.n725 B.n70 585
R279 B.n727 B.n726 585
R280 B.n728 B.n69 585
R281 B.n730 B.n729 585
R282 B.n731 B.n68 585
R283 B.n733 B.n732 585
R284 B.n734 B.n67 585
R285 B.n736 B.n735 585
R286 B.n737 B.n66 585
R287 B.n739 B.n738 585
R288 B.n741 B.n63 585
R289 B.n743 B.n742 585
R290 B.n744 B.n62 585
R291 B.n746 B.n745 585
R292 B.n747 B.n61 585
R293 B.n749 B.n748 585
R294 B.n750 B.n60 585
R295 B.n752 B.n751 585
R296 B.n753 B.n59 585
R297 B.n755 B.n754 585
R298 B.n757 B.n756 585
R299 B.n758 B.n55 585
R300 B.n760 B.n759 585
R301 B.n761 B.n54 585
R302 B.n763 B.n762 585
R303 B.n764 B.n53 585
R304 B.n766 B.n765 585
R305 B.n767 B.n52 585
R306 B.n769 B.n768 585
R307 B.n770 B.n51 585
R308 B.n772 B.n771 585
R309 B.n773 B.n50 585
R310 B.n775 B.n774 585
R311 B.n776 B.n49 585
R312 B.n778 B.n777 585
R313 B.n779 B.n48 585
R314 B.n781 B.n780 585
R315 B.n782 B.n47 585
R316 B.n784 B.n783 585
R317 B.n785 B.n46 585
R318 B.n787 B.n786 585
R319 B.n788 B.n45 585
R320 B.n790 B.n789 585
R321 B.n791 B.n44 585
R322 B.n793 B.n792 585
R323 B.n794 B.n43 585
R324 B.n796 B.n795 585
R325 B.n698 B.n79 585
R326 B.n697 B.n696 585
R327 B.n695 B.n80 585
R328 B.n694 B.n693 585
R329 B.n692 B.n81 585
R330 B.n691 B.n690 585
R331 B.n689 B.n82 585
R332 B.n688 B.n687 585
R333 B.n686 B.n83 585
R334 B.n685 B.n684 585
R335 B.n683 B.n84 585
R336 B.n682 B.n681 585
R337 B.n680 B.n85 585
R338 B.n679 B.n678 585
R339 B.n677 B.n86 585
R340 B.n676 B.n675 585
R341 B.n674 B.n87 585
R342 B.n673 B.n672 585
R343 B.n671 B.n88 585
R344 B.n670 B.n669 585
R345 B.n668 B.n89 585
R346 B.n667 B.n666 585
R347 B.n665 B.n90 585
R348 B.n664 B.n663 585
R349 B.n662 B.n91 585
R350 B.n661 B.n660 585
R351 B.n659 B.n92 585
R352 B.n658 B.n657 585
R353 B.n656 B.n93 585
R354 B.n655 B.n654 585
R355 B.n653 B.n94 585
R356 B.n652 B.n651 585
R357 B.n650 B.n95 585
R358 B.n649 B.n648 585
R359 B.n647 B.n96 585
R360 B.n646 B.n645 585
R361 B.n644 B.n97 585
R362 B.n643 B.n642 585
R363 B.n641 B.n98 585
R364 B.n640 B.n639 585
R365 B.n638 B.n99 585
R366 B.n637 B.n636 585
R367 B.n635 B.n100 585
R368 B.n634 B.n633 585
R369 B.n632 B.n101 585
R370 B.n631 B.n630 585
R371 B.n629 B.n102 585
R372 B.n628 B.n627 585
R373 B.n626 B.n103 585
R374 B.n625 B.n624 585
R375 B.n623 B.n104 585
R376 B.n622 B.n621 585
R377 B.n620 B.n105 585
R378 B.n619 B.n618 585
R379 B.n617 B.n106 585
R380 B.n616 B.n615 585
R381 B.n614 B.n107 585
R382 B.n613 B.n612 585
R383 B.n611 B.n108 585
R384 B.n610 B.n609 585
R385 B.n608 B.n109 585
R386 B.n607 B.n606 585
R387 B.n605 B.n110 585
R388 B.n604 B.n603 585
R389 B.n602 B.n111 585
R390 B.n601 B.n600 585
R391 B.n599 B.n112 585
R392 B.n598 B.n597 585
R393 B.n596 B.n113 585
R394 B.n595 B.n594 585
R395 B.n593 B.n114 585
R396 B.n592 B.n591 585
R397 B.n590 B.n115 585
R398 B.n589 B.n588 585
R399 B.n587 B.n116 585
R400 B.n586 B.n585 585
R401 B.n584 B.n117 585
R402 B.n583 B.n582 585
R403 B.n581 B.n118 585
R404 B.n580 B.n579 585
R405 B.n578 B.n119 585
R406 B.n577 B.n576 585
R407 B.n575 B.n120 585
R408 B.n574 B.n573 585
R409 B.n572 B.n121 585
R410 B.n571 B.n570 585
R411 B.n569 B.n122 585
R412 B.n568 B.n567 585
R413 B.n566 B.n123 585
R414 B.n565 B.n564 585
R415 B.n563 B.n124 585
R416 B.n562 B.n561 585
R417 B.n560 B.n125 585
R418 B.n559 B.n558 585
R419 B.n557 B.n126 585
R420 B.n556 B.n555 585
R421 B.n554 B.n127 585
R422 B.n553 B.n552 585
R423 B.n551 B.n128 585
R424 B.n550 B.n549 585
R425 B.n548 B.n129 585
R426 B.n547 B.n546 585
R427 B.n545 B.n130 585
R428 B.n544 B.n543 585
R429 B.n542 B.n131 585
R430 B.n541 B.n540 585
R431 B.n539 B.n132 585
R432 B.n538 B.n537 585
R433 B.n536 B.n133 585
R434 B.n535 B.n534 585
R435 B.n533 B.n134 585
R436 B.n532 B.n531 585
R437 B.n530 B.n135 585
R438 B.n529 B.n528 585
R439 B.n527 B.n136 585
R440 B.n526 B.n525 585
R441 B.n524 B.n137 585
R442 B.n523 B.n522 585
R443 B.n521 B.n138 585
R444 B.n520 B.n519 585
R445 B.n518 B.n139 585
R446 B.n517 B.n516 585
R447 B.n515 B.n140 585
R448 B.n514 B.n513 585
R449 B.n512 B.n141 585
R450 B.n511 B.n510 585
R451 B.n509 B.n142 585
R452 B.n508 B.n507 585
R453 B.n506 B.n143 585
R454 B.n505 B.n504 585
R455 B.n503 B.n144 585
R456 B.n502 B.n501 585
R457 B.n500 B.n145 585
R458 B.n499 B.n498 585
R459 B.n497 B.n146 585
R460 B.n496 B.n495 585
R461 B.n494 B.n147 585
R462 B.n493 B.n492 585
R463 B.n491 B.n148 585
R464 B.n490 B.n489 585
R465 B.n488 B.n149 585
R466 B.n487 B.n486 585
R467 B.n485 B.n150 585
R468 B.n484 B.n483 585
R469 B.n482 B.n151 585
R470 B.n481 B.n480 585
R471 B.n479 B.n152 585
R472 B.n478 B.n477 585
R473 B.n476 B.n153 585
R474 B.n475 B.n474 585
R475 B.n473 B.n154 585
R476 B.n472 B.n471 585
R477 B.n470 B.n155 585
R478 B.n469 B.n468 585
R479 B.n467 B.n156 585
R480 B.n466 B.n465 585
R481 B.n464 B.n157 585
R482 B.n463 B.n462 585
R483 B.n461 B.n158 585
R484 B.n460 B.n459 585
R485 B.n458 B.n159 585
R486 B.n457 B.n456 585
R487 B.n455 B.n160 585
R488 B.n358 B.n357 585
R489 B.n359 B.n196 585
R490 B.n361 B.n360 585
R491 B.n362 B.n195 585
R492 B.n364 B.n363 585
R493 B.n365 B.n194 585
R494 B.n367 B.n366 585
R495 B.n368 B.n193 585
R496 B.n370 B.n369 585
R497 B.n371 B.n192 585
R498 B.n373 B.n372 585
R499 B.n374 B.n191 585
R500 B.n376 B.n375 585
R501 B.n377 B.n190 585
R502 B.n379 B.n378 585
R503 B.n380 B.n189 585
R504 B.n382 B.n381 585
R505 B.n383 B.n188 585
R506 B.n385 B.n384 585
R507 B.n386 B.n187 585
R508 B.n388 B.n387 585
R509 B.n389 B.n186 585
R510 B.n391 B.n390 585
R511 B.n392 B.n185 585
R512 B.n394 B.n393 585
R513 B.n395 B.n184 585
R514 B.n397 B.n396 585
R515 B.n399 B.n181 585
R516 B.n401 B.n400 585
R517 B.n402 B.n180 585
R518 B.n404 B.n403 585
R519 B.n405 B.n179 585
R520 B.n407 B.n406 585
R521 B.n408 B.n178 585
R522 B.n410 B.n409 585
R523 B.n411 B.n177 585
R524 B.n413 B.n412 585
R525 B.n415 B.n414 585
R526 B.n416 B.n173 585
R527 B.n418 B.n417 585
R528 B.n419 B.n172 585
R529 B.n421 B.n420 585
R530 B.n422 B.n171 585
R531 B.n424 B.n423 585
R532 B.n425 B.n170 585
R533 B.n427 B.n426 585
R534 B.n428 B.n169 585
R535 B.n430 B.n429 585
R536 B.n431 B.n168 585
R537 B.n433 B.n432 585
R538 B.n434 B.n167 585
R539 B.n436 B.n435 585
R540 B.n437 B.n166 585
R541 B.n439 B.n438 585
R542 B.n440 B.n165 585
R543 B.n442 B.n441 585
R544 B.n443 B.n164 585
R545 B.n445 B.n444 585
R546 B.n446 B.n163 585
R547 B.n448 B.n447 585
R548 B.n449 B.n162 585
R549 B.n451 B.n450 585
R550 B.n452 B.n161 585
R551 B.n454 B.n453 585
R552 B.n356 B.n197 585
R553 B.n355 B.n354 585
R554 B.n353 B.n198 585
R555 B.n352 B.n351 585
R556 B.n350 B.n199 585
R557 B.n349 B.n348 585
R558 B.n347 B.n200 585
R559 B.n346 B.n345 585
R560 B.n344 B.n201 585
R561 B.n343 B.n342 585
R562 B.n341 B.n202 585
R563 B.n340 B.n339 585
R564 B.n338 B.n203 585
R565 B.n337 B.n336 585
R566 B.n335 B.n204 585
R567 B.n334 B.n333 585
R568 B.n332 B.n205 585
R569 B.n331 B.n330 585
R570 B.n329 B.n206 585
R571 B.n328 B.n327 585
R572 B.n326 B.n207 585
R573 B.n325 B.n324 585
R574 B.n323 B.n208 585
R575 B.n322 B.n321 585
R576 B.n320 B.n209 585
R577 B.n319 B.n318 585
R578 B.n317 B.n210 585
R579 B.n316 B.n315 585
R580 B.n314 B.n211 585
R581 B.n313 B.n312 585
R582 B.n311 B.n212 585
R583 B.n310 B.n309 585
R584 B.n308 B.n213 585
R585 B.n307 B.n306 585
R586 B.n305 B.n214 585
R587 B.n304 B.n303 585
R588 B.n302 B.n215 585
R589 B.n301 B.n300 585
R590 B.n299 B.n216 585
R591 B.n298 B.n297 585
R592 B.n296 B.n217 585
R593 B.n295 B.n294 585
R594 B.n293 B.n218 585
R595 B.n292 B.n291 585
R596 B.n290 B.n219 585
R597 B.n289 B.n288 585
R598 B.n287 B.n220 585
R599 B.n286 B.n285 585
R600 B.n284 B.n221 585
R601 B.n283 B.n282 585
R602 B.n281 B.n222 585
R603 B.n280 B.n279 585
R604 B.n278 B.n223 585
R605 B.n277 B.n276 585
R606 B.n275 B.n224 585
R607 B.n274 B.n273 585
R608 B.n272 B.n225 585
R609 B.n271 B.n270 585
R610 B.n269 B.n226 585
R611 B.n268 B.n267 585
R612 B.n266 B.n227 585
R613 B.n265 B.n264 585
R614 B.n263 B.n228 585
R615 B.n262 B.n261 585
R616 B.n260 B.n229 585
R617 B.n259 B.n258 585
R618 B.n257 B.n230 585
R619 B.n256 B.n255 585
R620 B.n254 B.n231 585
R621 B.n253 B.n252 585
R622 B.n251 B.n232 585
R623 B.n250 B.n249 585
R624 B.n248 B.n233 585
R625 B.n247 B.n246 585
R626 B.n245 B.n234 585
R627 B.n244 B.n243 585
R628 B.n242 B.n235 585
R629 B.n241 B.n240 585
R630 B.n239 B.n236 585
R631 B.n238 B.n237 585
R632 B.n2 B.n0 585
R633 B.n917 B.n1 585
R634 B.n916 B.n915 585
R635 B.n914 B.n3 585
R636 B.n913 B.n912 585
R637 B.n911 B.n4 585
R638 B.n910 B.n909 585
R639 B.n908 B.n5 585
R640 B.n907 B.n906 585
R641 B.n905 B.n6 585
R642 B.n904 B.n903 585
R643 B.n902 B.n7 585
R644 B.n901 B.n900 585
R645 B.n899 B.n8 585
R646 B.n898 B.n897 585
R647 B.n896 B.n9 585
R648 B.n895 B.n894 585
R649 B.n893 B.n10 585
R650 B.n892 B.n891 585
R651 B.n890 B.n11 585
R652 B.n889 B.n888 585
R653 B.n887 B.n12 585
R654 B.n886 B.n885 585
R655 B.n884 B.n13 585
R656 B.n883 B.n882 585
R657 B.n881 B.n14 585
R658 B.n880 B.n879 585
R659 B.n878 B.n15 585
R660 B.n877 B.n876 585
R661 B.n875 B.n16 585
R662 B.n874 B.n873 585
R663 B.n872 B.n17 585
R664 B.n871 B.n870 585
R665 B.n869 B.n18 585
R666 B.n868 B.n867 585
R667 B.n866 B.n19 585
R668 B.n865 B.n864 585
R669 B.n863 B.n20 585
R670 B.n862 B.n861 585
R671 B.n860 B.n21 585
R672 B.n859 B.n858 585
R673 B.n857 B.n22 585
R674 B.n856 B.n855 585
R675 B.n854 B.n23 585
R676 B.n853 B.n852 585
R677 B.n851 B.n24 585
R678 B.n850 B.n849 585
R679 B.n848 B.n25 585
R680 B.n847 B.n846 585
R681 B.n845 B.n26 585
R682 B.n844 B.n843 585
R683 B.n842 B.n27 585
R684 B.n841 B.n840 585
R685 B.n839 B.n28 585
R686 B.n838 B.n837 585
R687 B.n836 B.n29 585
R688 B.n835 B.n834 585
R689 B.n833 B.n30 585
R690 B.n832 B.n831 585
R691 B.n830 B.n31 585
R692 B.n829 B.n828 585
R693 B.n827 B.n32 585
R694 B.n826 B.n825 585
R695 B.n824 B.n33 585
R696 B.n823 B.n822 585
R697 B.n821 B.n34 585
R698 B.n820 B.n819 585
R699 B.n818 B.n35 585
R700 B.n817 B.n816 585
R701 B.n815 B.n36 585
R702 B.n814 B.n813 585
R703 B.n812 B.n37 585
R704 B.n811 B.n810 585
R705 B.n809 B.n38 585
R706 B.n808 B.n807 585
R707 B.n806 B.n39 585
R708 B.n805 B.n804 585
R709 B.n803 B.n40 585
R710 B.n802 B.n801 585
R711 B.n800 B.n41 585
R712 B.n799 B.n798 585
R713 B.n797 B.n42 585
R714 B.n919 B.n918 585
R715 B.n358 B.n197 478.086
R716 B.n797 B.n796 478.086
R717 B.n455 B.n454 478.086
R718 B.n700 B.n79 478.086
R719 B.n174 B.t0 254.119
R720 B.n182 B.t9 254.119
R721 B.n56 B.t6 254.119
R722 B.n64 B.t3 254.119
R723 B.n174 B.t2 194.718
R724 B.n64 B.t4 194.718
R725 B.n182 B.t11 194.709
R726 B.n56 B.t7 194.709
R727 B.n354 B.n197 163.367
R728 B.n354 B.n353 163.367
R729 B.n353 B.n352 163.367
R730 B.n352 B.n199 163.367
R731 B.n348 B.n199 163.367
R732 B.n348 B.n347 163.367
R733 B.n347 B.n346 163.367
R734 B.n346 B.n201 163.367
R735 B.n342 B.n201 163.367
R736 B.n342 B.n341 163.367
R737 B.n341 B.n340 163.367
R738 B.n340 B.n203 163.367
R739 B.n336 B.n203 163.367
R740 B.n336 B.n335 163.367
R741 B.n335 B.n334 163.367
R742 B.n334 B.n205 163.367
R743 B.n330 B.n205 163.367
R744 B.n330 B.n329 163.367
R745 B.n329 B.n328 163.367
R746 B.n328 B.n207 163.367
R747 B.n324 B.n207 163.367
R748 B.n324 B.n323 163.367
R749 B.n323 B.n322 163.367
R750 B.n322 B.n209 163.367
R751 B.n318 B.n209 163.367
R752 B.n318 B.n317 163.367
R753 B.n317 B.n316 163.367
R754 B.n316 B.n211 163.367
R755 B.n312 B.n211 163.367
R756 B.n312 B.n311 163.367
R757 B.n311 B.n310 163.367
R758 B.n310 B.n213 163.367
R759 B.n306 B.n213 163.367
R760 B.n306 B.n305 163.367
R761 B.n305 B.n304 163.367
R762 B.n304 B.n215 163.367
R763 B.n300 B.n215 163.367
R764 B.n300 B.n299 163.367
R765 B.n299 B.n298 163.367
R766 B.n298 B.n217 163.367
R767 B.n294 B.n217 163.367
R768 B.n294 B.n293 163.367
R769 B.n293 B.n292 163.367
R770 B.n292 B.n219 163.367
R771 B.n288 B.n219 163.367
R772 B.n288 B.n287 163.367
R773 B.n287 B.n286 163.367
R774 B.n286 B.n221 163.367
R775 B.n282 B.n221 163.367
R776 B.n282 B.n281 163.367
R777 B.n281 B.n280 163.367
R778 B.n280 B.n223 163.367
R779 B.n276 B.n223 163.367
R780 B.n276 B.n275 163.367
R781 B.n275 B.n274 163.367
R782 B.n274 B.n225 163.367
R783 B.n270 B.n225 163.367
R784 B.n270 B.n269 163.367
R785 B.n269 B.n268 163.367
R786 B.n268 B.n227 163.367
R787 B.n264 B.n227 163.367
R788 B.n264 B.n263 163.367
R789 B.n263 B.n262 163.367
R790 B.n262 B.n229 163.367
R791 B.n258 B.n229 163.367
R792 B.n258 B.n257 163.367
R793 B.n257 B.n256 163.367
R794 B.n256 B.n231 163.367
R795 B.n252 B.n231 163.367
R796 B.n252 B.n251 163.367
R797 B.n251 B.n250 163.367
R798 B.n250 B.n233 163.367
R799 B.n246 B.n233 163.367
R800 B.n246 B.n245 163.367
R801 B.n245 B.n244 163.367
R802 B.n244 B.n235 163.367
R803 B.n240 B.n235 163.367
R804 B.n240 B.n239 163.367
R805 B.n239 B.n238 163.367
R806 B.n238 B.n2 163.367
R807 B.n918 B.n2 163.367
R808 B.n918 B.n917 163.367
R809 B.n917 B.n916 163.367
R810 B.n916 B.n3 163.367
R811 B.n912 B.n3 163.367
R812 B.n912 B.n911 163.367
R813 B.n911 B.n910 163.367
R814 B.n910 B.n5 163.367
R815 B.n906 B.n5 163.367
R816 B.n906 B.n905 163.367
R817 B.n905 B.n904 163.367
R818 B.n904 B.n7 163.367
R819 B.n900 B.n7 163.367
R820 B.n900 B.n899 163.367
R821 B.n899 B.n898 163.367
R822 B.n898 B.n9 163.367
R823 B.n894 B.n9 163.367
R824 B.n894 B.n893 163.367
R825 B.n893 B.n892 163.367
R826 B.n892 B.n11 163.367
R827 B.n888 B.n11 163.367
R828 B.n888 B.n887 163.367
R829 B.n887 B.n886 163.367
R830 B.n886 B.n13 163.367
R831 B.n882 B.n13 163.367
R832 B.n882 B.n881 163.367
R833 B.n881 B.n880 163.367
R834 B.n880 B.n15 163.367
R835 B.n876 B.n15 163.367
R836 B.n876 B.n875 163.367
R837 B.n875 B.n874 163.367
R838 B.n874 B.n17 163.367
R839 B.n870 B.n17 163.367
R840 B.n870 B.n869 163.367
R841 B.n869 B.n868 163.367
R842 B.n868 B.n19 163.367
R843 B.n864 B.n19 163.367
R844 B.n864 B.n863 163.367
R845 B.n863 B.n862 163.367
R846 B.n862 B.n21 163.367
R847 B.n858 B.n21 163.367
R848 B.n858 B.n857 163.367
R849 B.n857 B.n856 163.367
R850 B.n856 B.n23 163.367
R851 B.n852 B.n23 163.367
R852 B.n852 B.n851 163.367
R853 B.n851 B.n850 163.367
R854 B.n850 B.n25 163.367
R855 B.n846 B.n25 163.367
R856 B.n846 B.n845 163.367
R857 B.n845 B.n844 163.367
R858 B.n844 B.n27 163.367
R859 B.n840 B.n27 163.367
R860 B.n840 B.n839 163.367
R861 B.n839 B.n838 163.367
R862 B.n838 B.n29 163.367
R863 B.n834 B.n29 163.367
R864 B.n834 B.n833 163.367
R865 B.n833 B.n832 163.367
R866 B.n832 B.n31 163.367
R867 B.n828 B.n31 163.367
R868 B.n828 B.n827 163.367
R869 B.n827 B.n826 163.367
R870 B.n826 B.n33 163.367
R871 B.n822 B.n33 163.367
R872 B.n822 B.n821 163.367
R873 B.n821 B.n820 163.367
R874 B.n820 B.n35 163.367
R875 B.n816 B.n35 163.367
R876 B.n816 B.n815 163.367
R877 B.n815 B.n814 163.367
R878 B.n814 B.n37 163.367
R879 B.n810 B.n37 163.367
R880 B.n810 B.n809 163.367
R881 B.n809 B.n808 163.367
R882 B.n808 B.n39 163.367
R883 B.n804 B.n39 163.367
R884 B.n804 B.n803 163.367
R885 B.n803 B.n802 163.367
R886 B.n802 B.n41 163.367
R887 B.n798 B.n41 163.367
R888 B.n798 B.n797 163.367
R889 B.n359 B.n358 163.367
R890 B.n360 B.n359 163.367
R891 B.n360 B.n195 163.367
R892 B.n364 B.n195 163.367
R893 B.n365 B.n364 163.367
R894 B.n366 B.n365 163.367
R895 B.n366 B.n193 163.367
R896 B.n370 B.n193 163.367
R897 B.n371 B.n370 163.367
R898 B.n372 B.n371 163.367
R899 B.n372 B.n191 163.367
R900 B.n376 B.n191 163.367
R901 B.n377 B.n376 163.367
R902 B.n378 B.n377 163.367
R903 B.n378 B.n189 163.367
R904 B.n382 B.n189 163.367
R905 B.n383 B.n382 163.367
R906 B.n384 B.n383 163.367
R907 B.n384 B.n187 163.367
R908 B.n388 B.n187 163.367
R909 B.n389 B.n388 163.367
R910 B.n390 B.n389 163.367
R911 B.n390 B.n185 163.367
R912 B.n394 B.n185 163.367
R913 B.n395 B.n394 163.367
R914 B.n396 B.n395 163.367
R915 B.n396 B.n181 163.367
R916 B.n401 B.n181 163.367
R917 B.n402 B.n401 163.367
R918 B.n403 B.n402 163.367
R919 B.n403 B.n179 163.367
R920 B.n407 B.n179 163.367
R921 B.n408 B.n407 163.367
R922 B.n409 B.n408 163.367
R923 B.n409 B.n177 163.367
R924 B.n413 B.n177 163.367
R925 B.n414 B.n413 163.367
R926 B.n414 B.n173 163.367
R927 B.n418 B.n173 163.367
R928 B.n419 B.n418 163.367
R929 B.n420 B.n419 163.367
R930 B.n420 B.n171 163.367
R931 B.n424 B.n171 163.367
R932 B.n425 B.n424 163.367
R933 B.n426 B.n425 163.367
R934 B.n426 B.n169 163.367
R935 B.n430 B.n169 163.367
R936 B.n431 B.n430 163.367
R937 B.n432 B.n431 163.367
R938 B.n432 B.n167 163.367
R939 B.n436 B.n167 163.367
R940 B.n437 B.n436 163.367
R941 B.n438 B.n437 163.367
R942 B.n438 B.n165 163.367
R943 B.n442 B.n165 163.367
R944 B.n443 B.n442 163.367
R945 B.n444 B.n443 163.367
R946 B.n444 B.n163 163.367
R947 B.n448 B.n163 163.367
R948 B.n449 B.n448 163.367
R949 B.n450 B.n449 163.367
R950 B.n450 B.n161 163.367
R951 B.n454 B.n161 163.367
R952 B.n456 B.n455 163.367
R953 B.n456 B.n159 163.367
R954 B.n460 B.n159 163.367
R955 B.n461 B.n460 163.367
R956 B.n462 B.n461 163.367
R957 B.n462 B.n157 163.367
R958 B.n466 B.n157 163.367
R959 B.n467 B.n466 163.367
R960 B.n468 B.n467 163.367
R961 B.n468 B.n155 163.367
R962 B.n472 B.n155 163.367
R963 B.n473 B.n472 163.367
R964 B.n474 B.n473 163.367
R965 B.n474 B.n153 163.367
R966 B.n478 B.n153 163.367
R967 B.n479 B.n478 163.367
R968 B.n480 B.n479 163.367
R969 B.n480 B.n151 163.367
R970 B.n484 B.n151 163.367
R971 B.n485 B.n484 163.367
R972 B.n486 B.n485 163.367
R973 B.n486 B.n149 163.367
R974 B.n490 B.n149 163.367
R975 B.n491 B.n490 163.367
R976 B.n492 B.n491 163.367
R977 B.n492 B.n147 163.367
R978 B.n496 B.n147 163.367
R979 B.n497 B.n496 163.367
R980 B.n498 B.n497 163.367
R981 B.n498 B.n145 163.367
R982 B.n502 B.n145 163.367
R983 B.n503 B.n502 163.367
R984 B.n504 B.n503 163.367
R985 B.n504 B.n143 163.367
R986 B.n508 B.n143 163.367
R987 B.n509 B.n508 163.367
R988 B.n510 B.n509 163.367
R989 B.n510 B.n141 163.367
R990 B.n514 B.n141 163.367
R991 B.n515 B.n514 163.367
R992 B.n516 B.n515 163.367
R993 B.n516 B.n139 163.367
R994 B.n520 B.n139 163.367
R995 B.n521 B.n520 163.367
R996 B.n522 B.n521 163.367
R997 B.n522 B.n137 163.367
R998 B.n526 B.n137 163.367
R999 B.n527 B.n526 163.367
R1000 B.n528 B.n527 163.367
R1001 B.n528 B.n135 163.367
R1002 B.n532 B.n135 163.367
R1003 B.n533 B.n532 163.367
R1004 B.n534 B.n533 163.367
R1005 B.n534 B.n133 163.367
R1006 B.n538 B.n133 163.367
R1007 B.n539 B.n538 163.367
R1008 B.n540 B.n539 163.367
R1009 B.n540 B.n131 163.367
R1010 B.n544 B.n131 163.367
R1011 B.n545 B.n544 163.367
R1012 B.n546 B.n545 163.367
R1013 B.n546 B.n129 163.367
R1014 B.n550 B.n129 163.367
R1015 B.n551 B.n550 163.367
R1016 B.n552 B.n551 163.367
R1017 B.n552 B.n127 163.367
R1018 B.n556 B.n127 163.367
R1019 B.n557 B.n556 163.367
R1020 B.n558 B.n557 163.367
R1021 B.n558 B.n125 163.367
R1022 B.n562 B.n125 163.367
R1023 B.n563 B.n562 163.367
R1024 B.n564 B.n563 163.367
R1025 B.n564 B.n123 163.367
R1026 B.n568 B.n123 163.367
R1027 B.n569 B.n568 163.367
R1028 B.n570 B.n569 163.367
R1029 B.n570 B.n121 163.367
R1030 B.n574 B.n121 163.367
R1031 B.n575 B.n574 163.367
R1032 B.n576 B.n575 163.367
R1033 B.n576 B.n119 163.367
R1034 B.n580 B.n119 163.367
R1035 B.n581 B.n580 163.367
R1036 B.n582 B.n581 163.367
R1037 B.n582 B.n117 163.367
R1038 B.n586 B.n117 163.367
R1039 B.n587 B.n586 163.367
R1040 B.n588 B.n587 163.367
R1041 B.n588 B.n115 163.367
R1042 B.n592 B.n115 163.367
R1043 B.n593 B.n592 163.367
R1044 B.n594 B.n593 163.367
R1045 B.n594 B.n113 163.367
R1046 B.n598 B.n113 163.367
R1047 B.n599 B.n598 163.367
R1048 B.n600 B.n599 163.367
R1049 B.n600 B.n111 163.367
R1050 B.n604 B.n111 163.367
R1051 B.n605 B.n604 163.367
R1052 B.n606 B.n605 163.367
R1053 B.n606 B.n109 163.367
R1054 B.n610 B.n109 163.367
R1055 B.n611 B.n610 163.367
R1056 B.n612 B.n611 163.367
R1057 B.n612 B.n107 163.367
R1058 B.n616 B.n107 163.367
R1059 B.n617 B.n616 163.367
R1060 B.n618 B.n617 163.367
R1061 B.n618 B.n105 163.367
R1062 B.n622 B.n105 163.367
R1063 B.n623 B.n622 163.367
R1064 B.n624 B.n623 163.367
R1065 B.n624 B.n103 163.367
R1066 B.n628 B.n103 163.367
R1067 B.n629 B.n628 163.367
R1068 B.n630 B.n629 163.367
R1069 B.n630 B.n101 163.367
R1070 B.n634 B.n101 163.367
R1071 B.n635 B.n634 163.367
R1072 B.n636 B.n635 163.367
R1073 B.n636 B.n99 163.367
R1074 B.n640 B.n99 163.367
R1075 B.n641 B.n640 163.367
R1076 B.n642 B.n641 163.367
R1077 B.n642 B.n97 163.367
R1078 B.n646 B.n97 163.367
R1079 B.n647 B.n646 163.367
R1080 B.n648 B.n647 163.367
R1081 B.n648 B.n95 163.367
R1082 B.n652 B.n95 163.367
R1083 B.n653 B.n652 163.367
R1084 B.n654 B.n653 163.367
R1085 B.n654 B.n93 163.367
R1086 B.n658 B.n93 163.367
R1087 B.n659 B.n658 163.367
R1088 B.n660 B.n659 163.367
R1089 B.n660 B.n91 163.367
R1090 B.n664 B.n91 163.367
R1091 B.n665 B.n664 163.367
R1092 B.n666 B.n665 163.367
R1093 B.n666 B.n89 163.367
R1094 B.n670 B.n89 163.367
R1095 B.n671 B.n670 163.367
R1096 B.n672 B.n671 163.367
R1097 B.n672 B.n87 163.367
R1098 B.n676 B.n87 163.367
R1099 B.n677 B.n676 163.367
R1100 B.n678 B.n677 163.367
R1101 B.n678 B.n85 163.367
R1102 B.n682 B.n85 163.367
R1103 B.n683 B.n682 163.367
R1104 B.n684 B.n683 163.367
R1105 B.n684 B.n83 163.367
R1106 B.n688 B.n83 163.367
R1107 B.n689 B.n688 163.367
R1108 B.n690 B.n689 163.367
R1109 B.n690 B.n81 163.367
R1110 B.n694 B.n81 163.367
R1111 B.n695 B.n694 163.367
R1112 B.n696 B.n695 163.367
R1113 B.n696 B.n79 163.367
R1114 B.n796 B.n43 163.367
R1115 B.n792 B.n43 163.367
R1116 B.n792 B.n791 163.367
R1117 B.n791 B.n790 163.367
R1118 B.n790 B.n45 163.367
R1119 B.n786 B.n45 163.367
R1120 B.n786 B.n785 163.367
R1121 B.n785 B.n784 163.367
R1122 B.n784 B.n47 163.367
R1123 B.n780 B.n47 163.367
R1124 B.n780 B.n779 163.367
R1125 B.n779 B.n778 163.367
R1126 B.n778 B.n49 163.367
R1127 B.n774 B.n49 163.367
R1128 B.n774 B.n773 163.367
R1129 B.n773 B.n772 163.367
R1130 B.n772 B.n51 163.367
R1131 B.n768 B.n51 163.367
R1132 B.n768 B.n767 163.367
R1133 B.n767 B.n766 163.367
R1134 B.n766 B.n53 163.367
R1135 B.n762 B.n53 163.367
R1136 B.n762 B.n761 163.367
R1137 B.n761 B.n760 163.367
R1138 B.n760 B.n55 163.367
R1139 B.n756 B.n55 163.367
R1140 B.n756 B.n755 163.367
R1141 B.n755 B.n59 163.367
R1142 B.n751 B.n59 163.367
R1143 B.n751 B.n750 163.367
R1144 B.n750 B.n749 163.367
R1145 B.n749 B.n61 163.367
R1146 B.n745 B.n61 163.367
R1147 B.n745 B.n744 163.367
R1148 B.n744 B.n743 163.367
R1149 B.n743 B.n63 163.367
R1150 B.n738 B.n63 163.367
R1151 B.n738 B.n737 163.367
R1152 B.n737 B.n736 163.367
R1153 B.n736 B.n67 163.367
R1154 B.n732 B.n67 163.367
R1155 B.n732 B.n731 163.367
R1156 B.n731 B.n730 163.367
R1157 B.n730 B.n69 163.367
R1158 B.n726 B.n69 163.367
R1159 B.n726 B.n725 163.367
R1160 B.n725 B.n724 163.367
R1161 B.n724 B.n71 163.367
R1162 B.n720 B.n71 163.367
R1163 B.n720 B.n719 163.367
R1164 B.n719 B.n718 163.367
R1165 B.n718 B.n73 163.367
R1166 B.n714 B.n73 163.367
R1167 B.n714 B.n713 163.367
R1168 B.n713 B.n712 163.367
R1169 B.n712 B.n75 163.367
R1170 B.n708 B.n75 163.367
R1171 B.n708 B.n707 163.367
R1172 B.n707 B.n706 163.367
R1173 B.n706 B.n77 163.367
R1174 B.n702 B.n77 163.367
R1175 B.n702 B.n701 163.367
R1176 B.n701 B.n700 163.367
R1177 B.n175 B.t1 114.621
R1178 B.n65 B.t5 114.621
R1179 B.n183 B.t10 114.612
R1180 B.n57 B.t8 114.612
R1181 B.n175 B.n174 80.0975
R1182 B.n183 B.n182 80.0975
R1183 B.n57 B.n56 80.0975
R1184 B.n65 B.n64 80.0975
R1185 B.n176 B.n175 59.5399
R1186 B.n398 B.n183 59.5399
R1187 B.n58 B.n57 59.5399
R1188 B.n740 B.n65 59.5399
R1189 B.n795 B.n42 31.0639
R1190 B.n699 B.n698 31.0639
R1191 B.n453 B.n160 31.0639
R1192 B.n357 B.n356 31.0639
R1193 B B.n919 18.0485
R1194 B.n795 B.n794 10.6151
R1195 B.n794 B.n793 10.6151
R1196 B.n793 B.n44 10.6151
R1197 B.n789 B.n44 10.6151
R1198 B.n789 B.n788 10.6151
R1199 B.n788 B.n787 10.6151
R1200 B.n787 B.n46 10.6151
R1201 B.n783 B.n46 10.6151
R1202 B.n783 B.n782 10.6151
R1203 B.n782 B.n781 10.6151
R1204 B.n781 B.n48 10.6151
R1205 B.n777 B.n48 10.6151
R1206 B.n777 B.n776 10.6151
R1207 B.n776 B.n775 10.6151
R1208 B.n775 B.n50 10.6151
R1209 B.n771 B.n50 10.6151
R1210 B.n771 B.n770 10.6151
R1211 B.n770 B.n769 10.6151
R1212 B.n769 B.n52 10.6151
R1213 B.n765 B.n52 10.6151
R1214 B.n765 B.n764 10.6151
R1215 B.n764 B.n763 10.6151
R1216 B.n763 B.n54 10.6151
R1217 B.n759 B.n54 10.6151
R1218 B.n759 B.n758 10.6151
R1219 B.n758 B.n757 10.6151
R1220 B.n754 B.n753 10.6151
R1221 B.n753 B.n752 10.6151
R1222 B.n752 B.n60 10.6151
R1223 B.n748 B.n60 10.6151
R1224 B.n748 B.n747 10.6151
R1225 B.n747 B.n746 10.6151
R1226 B.n746 B.n62 10.6151
R1227 B.n742 B.n62 10.6151
R1228 B.n742 B.n741 10.6151
R1229 B.n739 B.n66 10.6151
R1230 B.n735 B.n66 10.6151
R1231 B.n735 B.n734 10.6151
R1232 B.n734 B.n733 10.6151
R1233 B.n733 B.n68 10.6151
R1234 B.n729 B.n68 10.6151
R1235 B.n729 B.n728 10.6151
R1236 B.n728 B.n727 10.6151
R1237 B.n727 B.n70 10.6151
R1238 B.n723 B.n70 10.6151
R1239 B.n723 B.n722 10.6151
R1240 B.n722 B.n721 10.6151
R1241 B.n721 B.n72 10.6151
R1242 B.n717 B.n72 10.6151
R1243 B.n717 B.n716 10.6151
R1244 B.n716 B.n715 10.6151
R1245 B.n715 B.n74 10.6151
R1246 B.n711 B.n74 10.6151
R1247 B.n711 B.n710 10.6151
R1248 B.n710 B.n709 10.6151
R1249 B.n709 B.n76 10.6151
R1250 B.n705 B.n76 10.6151
R1251 B.n705 B.n704 10.6151
R1252 B.n704 B.n703 10.6151
R1253 B.n703 B.n78 10.6151
R1254 B.n699 B.n78 10.6151
R1255 B.n457 B.n160 10.6151
R1256 B.n458 B.n457 10.6151
R1257 B.n459 B.n458 10.6151
R1258 B.n459 B.n158 10.6151
R1259 B.n463 B.n158 10.6151
R1260 B.n464 B.n463 10.6151
R1261 B.n465 B.n464 10.6151
R1262 B.n465 B.n156 10.6151
R1263 B.n469 B.n156 10.6151
R1264 B.n470 B.n469 10.6151
R1265 B.n471 B.n470 10.6151
R1266 B.n471 B.n154 10.6151
R1267 B.n475 B.n154 10.6151
R1268 B.n476 B.n475 10.6151
R1269 B.n477 B.n476 10.6151
R1270 B.n477 B.n152 10.6151
R1271 B.n481 B.n152 10.6151
R1272 B.n482 B.n481 10.6151
R1273 B.n483 B.n482 10.6151
R1274 B.n483 B.n150 10.6151
R1275 B.n487 B.n150 10.6151
R1276 B.n488 B.n487 10.6151
R1277 B.n489 B.n488 10.6151
R1278 B.n489 B.n148 10.6151
R1279 B.n493 B.n148 10.6151
R1280 B.n494 B.n493 10.6151
R1281 B.n495 B.n494 10.6151
R1282 B.n495 B.n146 10.6151
R1283 B.n499 B.n146 10.6151
R1284 B.n500 B.n499 10.6151
R1285 B.n501 B.n500 10.6151
R1286 B.n501 B.n144 10.6151
R1287 B.n505 B.n144 10.6151
R1288 B.n506 B.n505 10.6151
R1289 B.n507 B.n506 10.6151
R1290 B.n507 B.n142 10.6151
R1291 B.n511 B.n142 10.6151
R1292 B.n512 B.n511 10.6151
R1293 B.n513 B.n512 10.6151
R1294 B.n513 B.n140 10.6151
R1295 B.n517 B.n140 10.6151
R1296 B.n518 B.n517 10.6151
R1297 B.n519 B.n518 10.6151
R1298 B.n519 B.n138 10.6151
R1299 B.n523 B.n138 10.6151
R1300 B.n524 B.n523 10.6151
R1301 B.n525 B.n524 10.6151
R1302 B.n525 B.n136 10.6151
R1303 B.n529 B.n136 10.6151
R1304 B.n530 B.n529 10.6151
R1305 B.n531 B.n530 10.6151
R1306 B.n531 B.n134 10.6151
R1307 B.n535 B.n134 10.6151
R1308 B.n536 B.n535 10.6151
R1309 B.n537 B.n536 10.6151
R1310 B.n537 B.n132 10.6151
R1311 B.n541 B.n132 10.6151
R1312 B.n542 B.n541 10.6151
R1313 B.n543 B.n542 10.6151
R1314 B.n543 B.n130 10.6151
R1315 B.n547 B.n130 10.6151
R1316 B.n548 B.n547 10.6151
R1317 B.n549 B.n548 10.6151
R1318 B.n549 B.n128 10.6151
R1319 B.n553 B.n128 10.6151
R1320 B.n554 B.n553 10.6151
R1321 B.n555 B.n554 10.6151
R1322 B.n555 B.n126 10.6151
R1323 B.n559 B.n126 10.6151
R1324 B.n560 B.n559 10.6151
R1325 B.n561 B.n560 10.6151
R1326 B.n561 B.n124 10.6151
R1327 B.n565 B.n124 10.6151
R1328 B.n566 B.n565 10.6151
R1329 B.n567 B.n566 10.6151
R1330 B.n567 B.n122 10.6151
R1331 B.n571 B.n122 10.6151
R1332 B.n572 B.n571 10.6151
R1333 B.n573 B.n572 10.6151
R1334 B.n573 B.n120 10.6151
R1335 B.n577 B.n120 10.6151
R1336 B.n578 B.n577 10.6151
R1337 B.n579 B.n578 10.6151
R1338 B.n579 B.n118 10.6151
R1339 B.n583 B.n118 10.6151
R1340 B.n584 B.n583 10.6151
R1341 B.n585 B.n584 10.6151
R1342 B.n585 B.n116 10.6151
R1343 B.n589 B.n116 10.6151
R1344 B.n590 B.n589 10.6151
R1345 B.n591 B.n590 10.6151
R1346 B.n591 B.n114 10.6151
R1347 B.n595 B.n114 10.6151
R1348 B.n596 B.n595 10.6151
R1349 B.n597 B.n596 10.6151
R1350 B.n597 B.n112 10.6151
R1351 B.n601 B.n112 10.6151
R1352 B.n602 B.n601 10.6151
R1353 B.n603 B.n602 10.6151
R1354 B.n603 B.n110 10.6151
R1355 B.n607 B.n110 10.6151
R1356 B.n608 B.n607 10.6151
R1357 B.n609 B.n608 10.6151
R1358 B.n609 B.n108 10.6151
R1359 B.n613 B.n108 10.6151
R1360 B.n614 B.n613 10.6151
R1361 B.n615 B.n614 10.6151
R1362 B.n615 B.n106 10.6151
R1363 B.n619 B.n106 10.6151
R1364 B.n620 B.n619 10.6151
R1365 B.n621 B.n620 10.6151
R1366 B.n621 B.n104 10.6151
R1367 B.n625 B.n104 10.6151
R1368 B.n626 B.n625 10.6151
R1369 B.n627 B.n626 10.6151
R1370 B.n627 B.n102 10.6151
R1371 B.n631 B.n102 10.6151
R1372 B.n632 B.n631 10.6151
R1373 B.n633 B.n632 10.6151
R1374 B.n633 B.n100 10.6151
R1375 B.n637 B.n100 10.6151
R1376 B.n638 B.n637 10.6151
R1377 B.n639 B.n638 10.6151
R1378 B.n639 B.n98 10.6151
R1379 B.n643 B.n98 10.6151
R1380 B.n644 B.n643 10.6151
R1381 B.n645 B.n644 10.6151
R1382 B.n645 B.n96 10.6151
R1383 B.n649 B.n96 10.6151
R1384 B.n650 B.n649 10.6151
R1385 B.n651 B.n650 10.6151
R1386 B.n651 B.n94 10.6151
R1387 B.n655 B.n94 10.6151
R1388 B.n656 B.n655 10.6151
R1389 B.n657 B.n656 10.6151
R1390 B.n657 B.n92 10.6151
R1391 B.n661 B.n92 10.6151
R1392 B.n662 B.n661 10.6151
R1393 B.n663 B.n662 10.6151
R1394 B.n663 B.n90 10.6151
R1395 B.n667 B.n90 10.6151
R1396 B.n668 B.n667 10.6151
R1397 B.n669 B.n668 10.6151
R1398 B.n669 B.n88 10.6151
R1399 B.n673 B.n88 10.6151
R1400 B.n674 B.n673 10.6151
R1401 B.n675 B.n674 10.6151
R1402 B.n675 B.n86 10.6151
R1403 B.n679 B.n86 10.6151
R1404 B.n680 B.n679 10.6151
R1405 B.n681 B.n680 10.6151
R1406 B.n681 B.n84 10.6151
R1407 B.n685 B.n84 10.6151
R1408 B.n686 B.n685 10.6151
R1409 B.n687 B.n686 10.6151
R1410 B.n687 B.n82 10.6151
R1411 B.n691 B.n82 10.6151
R1412 B.n692 B.n691 10.6151
R1413 B.n693 B.n692 10.6151
R1414 B.n693 B.n80 10.6151
R1415 B.n697 B.n80 10.6151
R1416 B.n698 B.n697 10.6151
R1417 B.n357 B.n196 10.6151
R1418 B.n361 B.n196 10.6151
R1419 B.n362 B.n361 10.6151
R1420 B.n363 B.n362 10.6151
R1421 B.n363 B.n194 10.6151
R1422 B.n367 B.n194 10.6151
R1423 B.n368 B.n367 10.6151
R1424 B.n369 B.n368 10.6151
R1425 B.n369 B.n192 10.6151
R1426 B.n373 B.n192 10.6151
R1427 B.n374 B.n373 10.6151
R1428 B.n375 B.n374 10.6151
R1429 B.n375 B.n190 10.6151
R1430 B.n379 B.n190 10.6151
R1431 B.n380 B.n379 10.6151
R1432 B.n381 B.n380 10.6151
R1433 B.n381 B.n188 10.6151
R1434 B.n385 B.n188 10.6151
R1435 B.n386 B.n385 10.6151
R1436 B.n387 B.n386 10.6151
R1437 B.n387 B.n186 10.6151
R1438 B.n391 B.n186 10.6151
R1439 B.n392 B.n391 10.6151
R1440 B.n393 B.n392 10.6151
R1441 B.n393 B.n184 10.6151
R1442 B.n397 B.n184 10.6151
R1443 B.n400 B.n399 10.6151
R1444 B.n400 B.n180 10.6151
R1445 B.n404 B.n180 10.6151
R1446 B.n405 B.n404 10.6151
R1447 B.n406 B.n405 10.6151
R1448 B.n406 B.n178 10.6151
R1449 B.n410 B.n178 10.6151
R1450 B.n411 B.n410 10.6151
R1451 B.n412 B.n411 10.6151
R1452 B.n416 B.n415 10.6151
R1453 B.n417 B.n416 10.6151
R1454 B.n417 B.n172 10.6151
R1455 B.n421 B.n172 10.6151
R1456 B.n422 B.n421 10.6151
R1457 B.n423 B.n422 10.6151
R1458 B.n423 B.n170 10.6151
R1459 B.n427 B.n170 10.6151
R1460 B.n428 B.n427 10.6151
R1461 B.n429 B.n428 10.6151
R1462 B.n429 B.n168 10.6151
R1463 B.n433 B.n168 10.6151
R1464 B.n434 B.n433 10.6151
R1465 B.n435 B.n434 10.6151
R1466 B.n435 B.n166 10.6151
R1467 B.n439 B.n166 10.6151
R1468 B.n440 B.n439 10.6151
R1469 B.n441 B.n440 10.6151
R1470 B.n441 B.n164 10.6151
R1471 B.n445 B.n164 10.6151
R1472 B.n446 B.n445 10.6151
R1473 B.n447 B.n446 10.6151
R1474 B.n447 B.n162 10.6151
R1475 B.n451 B.n162 10.6151
R1476 B.n452 B.n451 10.6151
R1477 B.n453 B.n452 10.6151
R1478 B.n356 B.n355 10.6151
R1479 B.n355 B.n198 10.6151
R1480 B.n351 B.n198 10.6151
R1481 B.n351 B.n350 10.6151
R1482 B.n350 B.n349 10.6151
R1483 B.n349 B.n200 10.6151
R1484 B.n345 B.n200 10.6151
R1485 B.n345 B.n344 10.6151
R1486 B.n344 B.n343 10.6151
R1487 B.n343 B.n202 10.6151
R1488 B.n339 B.n202 10.6151
R1489 B.n339 B.n338 10.6151
R1490 B.n338 B.n337 10.6151
R1491 B.n337 B.n204 10.6151
R1492 B.n333 B.n204 10.6151
R1493 B.n333 B.n332 10.6151
R1494 B.n332 B.n331 10.6151
R1495 B.n331 B.n206 10.6151
R1496 B.n327 B.n206 10.6151
R1497 B.n327 B.n326 10.6151
R1498 B.n326 B.n325 10.6151
R1499 B.n325 B.n208 10.6151
R1500 B.n321 B.n208 10.6151
R1501 B.n321 B.n320 10.6151
R1502 B.n320 B.n319 10.6151
R1503 B.n319 B.n210 10.6151
R1504 B.n315 B.n210 10.6151
R1505 B.n315 B.n314 10.6151
R1506 B.n314 B.n313 10.6151
R1507 B.n313 B.n212 10.6151
R1508 B.n309 B.n212 10.6151
R1509 B.n309 B.n308 10.6151
R1510 B.n308 B.n307 10.6151
R1511 B.n307 B.n214 10.6151
R1512 B.n303 B.n214 10.6151
R1513 B.n303 B.n302 10.6151
R1514 B.n302 B.n301 10.6151
R1515 B.n301 B.n216 10.6151
R1516 B.n297 B.n216 10.6151
R1517 B.n297 B.n296 10.6151
R1518 B.n296 B.n295 10.6151
R1519 B.n295 B.n218 10.6151
R1520 B.n291 B.n218 10.6151
R1521 B.n291 B.n290 10.6151
R1522 B.n290 B.n289 10.6151
R1523 B.n289 B.n220 10.6151
R1524 B.n285 B.n220 10.6151
R1525 B.n285 B.n284 10.6151
R1526 B.n284 B.n283 10.6151
R1527 B.n283 B.n222 10.6151
R1528 B.n279 B.n222 10.6151
R1529 B.n279 B.n278 10.6151
R1530 B.n278 B.n277 10.6151
R1531 B.n277 B.n224 10.6151
R1532 B.n273 B.n224 10.6151
R1533 B.n273 B.n272 10.6151
R1534 B.n272 B.n271 10.6151
R1535 B.n271 B.n226 10.6151
R1536 B.n267 B.n226 10.6151
R1537 B.n267 B.n266 10.6151
R1538 B.n266 B.n265 10.6151
R1539 B.n265 B.n228 10.6151
R1540 B.n261 B.n228 10.6151
R1541 B.n261 B.n260 10.6151
R1542 B.n260 B.n259 10.6151
R1543 B.n259 B.n230 10.6151
R1544 B.n255 B.n230 10.6151
R1545 B.n255 B.n254 10.6151
R1546 B.n254 B.n253 10.6151
R1547 B.n253 B.n232 10.6151
R1548 B.n249 B.n232 10.6151
R1549 B.n249 B.n248 10.6151
R1550 B.n248 B.n247 10.6151
R1551 B.n247 B.n234 10.6151
R1552 B.n243 B.n234 10.6151
R1553 B.n243 B.n242 10.6151
R1554 B.n242 B.n241 10.6151
R1555 B.n241 B.n236 10.6151
R1556 B.n237 B.n236 10.6151
R1557 B.n237 B.n0 10.6151
R1558 B.n915 B.n1 10.6151
R1559 B.n915 B.n914 10.6151
R1560 B.n914 B.n913 10.6151
R1561 B.n913 B.n4 10.6151
R1562 B.n909 B.n4 10.6151
R1563 B.n909 B.n908 10.6151
R1564 B.n908 B.n907 10.6151
R1565 B.n907 B.n6 10.6151
R1566 B.n903 B.n6 10.6151
R1567 B.n903 B.n902 10.6151
R1568 B.n902 B.n901 10.6151
R1569 B.n901 B.n8 10.6151
R1570 B.n897 B.n8 10.6151
R1571 B.n897 B.n896 10.6151
R1572 B.n896 B.n895 10.6151
R1573 B.n895 B.n10 10.6151
R1574 B.n891 B.n10 10.6151
R1575 B.n891 B.n890 10.6151
R1576 B.n890 B.n889 10.6151
R1577 B.n889 B.n12 10.6151
R1578 B.n885 B.n12 10.6151
R1579 B.n885 B.n884 10.6151
R1580 B.n884 B.n883 10.6151
R1581 B.n883 B.n14 10.6151
R1582 B.n879 B.n14 10.6151
R1583 B.n879 B.n878 10.6151
R1584 B.n878 B.n877 10.6151
R1585 B.n877 B.n16 10.6151
R1586 B.n873 B.n16 10.6151
R1587 B.n873 B.n872 10.6151
R1588 B.n872 B.n871 10.6151
R1589 B.n871 B.n18 10.6151
R1590 B.n867 B.n18 10.6151
R1591 B.n867 B.n866 10.6151
R1592 B.n866 B.n865 10.6151
R1593 B.n865 B.n20 10.6151
R1594 B.n861 B.n20 10.6151
R1595 B.n861 B.n860 10.6151
R1596 B.n860 B.n859 10.6151
R1597 B.n859 B.n22 10.6151
R1598 B.n855 B.n22 10.6151
R1599 B.n855 B.n854 10.6151
R1600 B.n854 B.n853 10.6151
R1601 B.n853 B.n24 10.6151
R1602 B.n849 B.n24 10.6151
R1603 B.n849 B.n848 10.6151
R1604 B.n848 B.n847 10.6151
R1605 B.n847 B.n26 10.6151
R1606 B.n843 B.n26 10.6151
R1607 B.n843 B.n842 10.6151
R1608 B.n842 B.n841 10.6151
R1609 B.n841 B.n28 10.6151
R1610 B.n837 B.n28 10.6151
R1611 B.n837 B.n836 10.6151
R1612 B.n836 B.n835 10.6151
R1613 B.n835 B.n30 10.6151
R1614 B.n831 B.n30 10.6151
R1615 B.n831 B.n830 10.6151
R1616 B.n830 B.n829 10.6151
R1617 B.n829 B.n32 10.6151
R1618 B.n825 B.n32 10.6151
R1619 B.n825 B.n824 10.6151
R1620 B.n824 B.n823 10.6151
R1621 B.n823 B.n34 10.6151
R1622 B.n819 B.n34 10.6151
R1623 B.n819 B.n818 10.6151
R1624 B.n818 B.n817 10.6151
R1625 B.n817 B.n36 10.6151
R1626 B.n813 B.n36 10.6151
R1627 B.n813 B.n812 10.6151
R1628 B.n812 B.n811 10.6151
R1629 B.n811 B.n38 10.6151
R1630 B.n807 B.n38 10.6151
R1631 B.n807 B.n806 10.6151
R1632 B.n806 B.n805 10.6151
R1633 B.n805 B.n40 10.6151
R1634 B.n801 B.n40 10.6151
R1635 B.n801 B.n800 10.6151
R1636 B.n800 B.n799 10.6151
R1637 B.n799 B.n42 10.6151
R1638 B.n757 B.n58 9.36635
R1639 B.n740 B.n739 9.36635
R1640 B.n398 B.n397 9.36635
R1641 B.n415 B.n176 9.36635
R1642 B.n919 B.n0 2.81026
R1643 B.n919 B.n1 2.81026
R1644 B.n754 B.n58 1.24928
R1645 B.n741 B.n740 1.24928
R1646 B.n399 B.n398 1.24928
R1647 B.n412 B.n176 1.24928
R1648 VN.n110 VN.n109 161.3
R1649 VN.n108 VN.n57 161.3
R1650 VN.n107 VN.n106 161.3
R1651 VN.n105 VN.n58 161.3
R1652 VN.n104 VN.n103 161.3
R1653 VN.n102 VN.n59 161.3
R1654 VN.n101 VN.n100 161.3
R1655 VN.n99 VN.n60 161.3
R1656 VN.n98 VN.n97 161.3
R1657 VN.n95 VN.n61 161.3
R1658 VN.n94 VN.n93 161.3
R1659 VN.n92 VN.n62 161.3
R1660 VN.n91 VN.n90 161.3
R1661 VN.n89 VN.n63 161.3
R1662 VN.n88 VN.n87 161.3
R1663 VN.n86 VN.n64 161.3
R1664 VN.n85 VN.n84 161.3
R1665 VN.n82 VN.n65 161.3
R1666 VN.n81 VN.n80 161.3
R1667 VN.n79 VN.n66 161.3
R1668 VN.n78 VN.n77 161.3
R1669 VN.n76 VN.n67 161.3
R1670 VN.n75 VN.n74 161.3
R1671 VN.n73 VN.n68 161.3
R1672 VN.n72 VN.n71 161.3
R1673 VN.n54 VN.n53 161.3
R1674 VN.n52 VN.n1 161.3
R1675 VN.n51 VN.n50 161.3
R1676 VN.n49 VN.n2 161.3
R1677 VN.n48 VN.n47 161.3
R1678 VN.n46 VN.n3 161.3
R1679 VN.n45 VN.n44 161.3
R1680 VN.n43 VN.n4 161.3
R1681 VN.n42 VN.n41 161.3
R1682 VN.n39 VN.n5 161.3
R1683 VN.n38 VN.n37 161.3
R1684 VN.n36 VN.n6 161.3
R1685 VN.n35 VN.n34 161.3
R1686 VN.n33 VN.n7 161.3
R1687 VN.n32 VN.n31 161.3
R1688 VN.n30 VN.n8 161.3
R1689 VN.n29 VN.n28 161.3
R1690 VN.n26 VN.n9 161.3
R1691 VN.n25 VN.n24 161.3
R1692 VN.n23 VN.n10 161.3
R1693 VN.n22 VN.n21 161.3
R1694 VN.n20 VN.n11 161.3
R1695 VN.n19 VN.n18 161.3
R1696 VN.n17 VN.n12 161.3
R1697 VN.n16 VN.n15 161.3
R1698 VN.n55 VN.n0 89.7537
R1699 VN.n111 VN.n56 89.7537
R1700 VN.n69 VN.t2 77.0548
R1701 VN.n13 VN.t1 77.0548
R1702 VN.n14 VN.n13 56.597
R1703 VN.n70 VN.n69 56.597
R1704 VN.n21 VN.n20 56.5617
R1705 VN.n34 VN.n33 56.5617
R1706 VN.n77 VN.n76 56.5617
R1707 VN.n90 VN.n89 56.5617
R1708 VN VN.n111 56.0777
R1709 VN.n47 VN.n46 45.9053
R1710 VN.n103 VN.n102 45.9053
R1711 VN.n14 VN.t0 44.7758
R1712 VN.n27 VN.t9 44.7758
R1713 VN.n40 VN.t7 44.7758
R1714 VN.n0 VN.t5 44.7758
R1715 VN.n70 VN.t3 44.7758
R1716 VN.n83 VN.t4 44.7758
R1717 VN.n96 VN.t8 44.7758
R1718 VN.n56 VN.t6 44.7758
R1719 VN.n47 VN.n2 35.2488
R1720 VN.n103 VN.n58 35.2488
R1721 VN.n15 VN.n12 24.5923
R1722 VN.n19 VN.n12 24.5923
R1723 VN.n20 VN.n19 24.5923
R1724 VN.n21 VN.n10 24.5923
R1725 VN.n25 VN.n10 24.5923
R1726 VN.n26 VN.n25 24.5923
R1727 VN.n28 VN.n8 24.5923
R1728 VN.n32 VN.n8 24.5923
R1729 VN.n33 VN.n32 24.5923
R1730 VN.n34 VN.n6 24.5923
R1731 VN.n38 VN.n6 24.5923
R1732 VN.n39 VN.n38 24.5923
R1733 VN.n41 VN.n4 24.5923
R1734 VN.n45 VN.n4 24.5923
R1735 VN.n46 VN.n45 24.5923
R1736 VN.n51 VN.n2 24.5923
R1737 VN.n52 VN.n51 24.5923
R1738 VN.n53 VN.n52 24.5923
R1739 VN.n76 VN.n75 24.5923
R1740 VN.n75 VN.n68 24.5923
R1741 VN.n71 VN.n68 24.5923
R1742 VN.n89 VN.n88 24.5923
R1743 VN.n88 VN.n64 24.5923
R1744 VN.n84 VN.n64 24.5923
R1745 VN.n82 VN.n81 24.5923
R1746 VN.n81 VN.n66 24.5923
R1747 VN.n77 VN.n66 24.5923
R1748 VN.n102 VN.n101 24.5923
R1749 VN.n101 VN.n60 24.5923
R1750 VN.n97 VN.n60 24.5923
R1751 VN.n95 VN.n94 24.5923
R1752 VN.n94 VN.n62 24.5923
R1753 VN.n90 VN.n62 24.5923
R1754 VN.n109 VN.n108 24.5923
R1755 VN.n108 VN.n107 24.5923
R1756 VN.n107 VN.n58 24.5923
R1757 VN.n15 VN.n14 18.6903
R1758 VN.n40 VN.n39 18.6903
R1759 VN.n71 VN.n70 18.6903
R1760 VN.n96 VN.n95 18.6903
R1761 VN.n27 VN.n26 12.2964
R1762 VN.n28 VN.n27 12.2964
R1763 VN.n84 VN.n83 12.2964
R1764 VN.n83 VN.n82 12.2964
R1765 VN.n41 VN.n40 5.90254
R1766 VN.n97 VN.n96 5.90254
R1767 VN.n72 VN.n69 2.50626
R1768 VN.n16 VN.n13 2.50626
R1769 VN.n53 VN.n0 0.492337
R1770 VN.n109 VN.n56 0.492337
R1771 VN.n111 VN.n110 0.354861
R1772 VN.n55 VN.n54 0.354861
R1773 VN VN.n55 0.267071
R1774 VN.n110 VN.n57 0.189894
R1775 VN.n106 VN.n57 0.189894
R1776 VN.n106 VN.n105 0.189894
R1777 VN.n105 VN.n104 0.189894
R1778 VN.n104 VN.n59 0.189894
R1779 VN.n100 VN.n59 0.189894
R1780 VN.n100 VN.n99 0.189894
R1781 VN.n99 VN.n98 0.189894
R1782 VN.n98 VN.n61 0.189894
R1783 VN.n93 VN.n61 0.189894
R1784 VN.n93 VN.n92 0.189894
R1785 VN.n92 VN.n91 0.189894
R1786 VN.n91 VN.n63 0.189894
R1787 VN.n87 VN.n63 0.189894
R1788 VN.n87 VN.n86 0.189894
R1789 VN.n86 VN.n85 0.189894
R1790 VN.n85 VN.n65 0.189894
R1791 VN.n80 VN.n65 0.189894
R1792 VN.n80 VN.n79 0.189894
R1793 VN.n79 VN.n78 0.189894
R1794 VN.n78 VN.n67 0.189894
R1795 VN.n74 VN.n67 0.189894
R1796 VN.n74 VN.n73 0.189894
R1797 VN.n73 VN.n72 0.189894
R1798 VN.n17 VN.n16 0.189894
R1799 VN.n18 VN.n17 0.189894
R1800 VN.n18 VN.n11 0.189894
R1801 VN.n22 VN.n11 0.189894
R1802 VN.n23 VN.n22 0.189894
R1803 VN.n24 VN.n23 0.189894
R1804 VN.n24 VN.n9 0.189894
R1805 VN.n29 VN.n9 0.189894
R1806 VN.n30 VN.n29 0.189894
R1807 VN.n31 VN.n30 0.189894
R1808 VN.n31 VN.n7 0.189894
R1809 VN.n35 VN.n7 0.189894
R1810 VN.n36 VN.n35 0.189894
R1811 VN.n37 VN.n36 0.189894
R1812 VN.n37 VN.n5 0.189894
R1813 VN.n42 VN.n5 0.189894
R1814 VN.n43 VN.n42 0.189894
R1815 VN.n44 VN.n43 0.189894
R1816 VN.n44 VN.n3 0.189894
R1817 VN.n48 VN.n3 0.189894
R1818 VN.n49 VN.n48 0.189894
R1819 VN.n50 VN.n49 0.189894
R1820 VN.n50 VN.n1 0.189894
R1821 VN.n54 VN.n1 0.189894
R1822 VDD2.n1 VDD2.t8 94.5425
R1823 VDD2.n4 VDD2.t3 90.9824
R1824 VDD2.n3 VDD2.n2 88.9931
R1825 VDD2 VDD2.n7 88.9901
R1826 VDD2.n6 VDD2.n5 86.3782
R1827 VDD2.n1 VDD2.n0 86.3782
R1828 VDD2.n4 VDD2.n3 46.7131
R1829 VDD2.n7 VDD2.t6 4.60461
R1830 VDD2.n7 VDD2.t7 4.60461
R1831 VDD2.n5 VDD2.t1 4.60461
R1832 VDD2.n5 VDD2.t5 4.60461
R1833 VDD2.n2 VDD2.t2 4.60461
R1834 VDD2.n2 VDD2.t4 4.60461
R1835 VDD2.n0 VDD2.t9 4.60461
R1836 VDD2.n0 VDD2.t0 4.60461
R1837 VDD2.n6 VDD2.n4 3.56084
R1838 VDD2 VDD2.n6 0.948776
R1839 VDD2.n3 VDD2.n1 0.83524
C0 B VDD2 2.71165f
C1 VN VP 9.246429f
C2 VP VDD1 7.49404f
C3 VN VDD2 6.91711f
C4 VDD2 VDD1 2.9557f
C5 B VN 1.53468f
C6 B VDD1 2.54701f
C7 VN VDD1 0.156413f
C8 w_n5926_n2380# VTAIL 2.71816f
C9 VP w_n5926_n2380# 13.7111f
C10 VP VTAIL 8.596901f
C11 VDD2 w_n5926_n2380# 3.11103f
C12 VDD2 VTAIL 9.15909f
C13 B w_n5926_n2380# 11.183f
C14 VDD2 VP 0.736438f
C15 B VTAIL 2.9991f
C16 VN w_n5926_n2380# 12.935901f
C17 w_n5926_n2380# VDD1 2.90511f
C18 VN VTAIL 8.58243f
C19 VTAIL VDD1 9.098371f
C20 B VP 2.84491f
C21 VDD2 VSUBS 2.592846f
C22 VDD1 VSUBS 2.356831f
C23 VTAIL VSUBS 0.833795f
C24 VN VSUBS 9.420589f
C25 VP VSUBS 5.280796f
C26 B VSUBS 6.438031f
C27 w_n5926_n2380# VSUBS 0.175433p
C28 VDD2.t8 VSUBS 1.81462f
C29 VDD2.t9 VSUBS 0.192767f
C30 VDD2.t0 VSUBS 0.192767f
C31 VDD2.n0 VSUBS 1.33233f
C32 VDD2.n1 VSUBS 2.12361f
C33 VDD2.t2 VSUBS 0.192767f
C34 VDD2.t4 VSUBS 0.192767f
C35 VDD2.n2 VSUBS 1.37028f
C36 VDD2.n3 VSUBS 4.76293f
C37 VDD2.t3 VSUBS 1.77379f
C38 VDD2.n4 VSUBS 4.73658f
C39 VDD2.t1 VSUBS 0.192767f
C40 VDD2.t5 VSUBS 0.192767f
C41 VDD2.n5 VSUBS 1.33234f
C42 VDD2.n6 VSUBS 1.09175f
C43 VDD2.t6 VSUBS 0.192767f
C44 VDD2.t7 VSUBS 0.192767f
C45 VDD2.n7 VSUBS 1.37022f
C46 VN.t5 VSUBS 2.04307f
C47 VN.n0 VSUBS 0.843675f
C48 VN.n1 VSUBS 0.028521f
C49 VN.n2 VSUBS 0.057309f
C50 VN.n3 VSUBS 0.028521f
C51 VN.n4 VSUBS 0.052889f
C52 VN.n5 VSUBS 0.028521f
C53 VN.t7 VSUBS 2.04307f
C54 VN.n6 VSUBS 0.052889f
C55 VN.n7 VSUBS 0.028521f
C56 VN.n8 VSUBS 0.052889f
C57 VN.n9 VSUBS 0.028521f
C58 VN.t9 VSUBS 2.04307f
C59 VN.n10 VSUBS 0.052889f
C60 VN.n11 VSUBS 0.028521f
C61 VN.n12 VSUBS 0.052889f
C62 VN.t1 VSUBS 2.44788f
C63 VN.n13 VSUBS 0.818465f
C64 VN.t0 VSUBS 2.04307f
C65 VN.n14 VSUBS 0.849847f
C66 VN.n15 VSUBS 0.046622f
C67 VN.n16 VSUBS 0.367595f
C68 VN.n17 VSUBS 0.028521f
C69 VN.n18 VSUBS 0.028521f
C70 VN.n19 VSUBS 0.052889f
C71 VN.n20 VSUBS 0.03633f
C72 VN.n21 VSUBS 0.046588f
C73 VN.n22 VSUBS 0.028521f
C74 VN.n23 VSUBS 0.028521f
C75 VN.n24 VSUBS 0.028521f
C76 VN.n25 VSUBS 0.052889f
C77 VN.n26 VSUBS 0.039834f
C78 VN.n27 VSUBS 0.74088f
C79 VN.n28 VSUBS 0.039834f
C80 VN.n29 VSUBS 0.028521f
C81 VN.n30 VSUBS 0.028521f
C82 VN.n31 VSUBS 0.028521f
C83 VN.n32 VSUBS 0.052889f
C84 VN.n33 VSUBS 0.046588f
C85 VN.n34 VSUBS 0.03633f
C86 VN.n35 VSUBS 0.028521f
C87 VN.n36 VSUBS 0.028521f
C88 VN.n37 VSUBS 0.028521f
C89 VN.n38 VSUBS 0.052889f
C90 VN.n39 VSUBS 0.046622f
C91 VN.n40 VSUBS 0.74088f
C92 VN.n41 VSUBS 0.033045f
C93 VN.n42 VSUBS 0.028521f
C94 VN.n43 VSUBS 0.028521f
C95 VN.n44 VSUBS 0.028521f
C96 VN.n45 VSUBS 0.052889f
C97 VN.n46 VSUBS 0.054343f
C98 VN.n47 VSUBS 0.024154f
C99 VN.n48 VSUBS 0.028521f
C100 VN.n49 VSUBS 0.028521f
C101 VN.n50 VSUBS 0.028521f
C102 VN.n51 VSUBS 0.052889f
C103 VN.n52 VSUBS 0.052889f
C104 VN.n53 VSUBS 0.027301f
C105 VN.n54 VSUBS 0.046024f
C106 VN.n55 VSUBS 0.089409f
C107 VN.t6 VSUBS 2.04307f
C108 VN.n56 VSUBS 0.843675f
C109 VN.n57 VSUBS 0.028521f
C110 VN.n58 VSUBS 0.057309f
C111 VN.n59 VSUBS 0.028521f
C112 VN.n60 VSUBS 0.052889f
C113 VN.n61 VSUBS 0.028521f
C114 VN.t8 VSUBS 2.04307f
C115 VN.n62 VSUBS 0.052889f
C116 VN.n63 VSUBS 0.028521f
C117 VN.n64 VSUBS 0.052889f
C118 VN.n65 VSUBS 0.028521f
C119 VN.t4 VSUBS 2.04307f
C120 VN.n66 VSUBS 0.052889f
C121 VN.n67 VSUBS 0.028521f
C122 VN.n68 VSUBS 0.052889f
C123 VN.t2 VSUBS 2.44788f
C124 VN.n69 VSUBS 0.818465f
C125 VN.t3 VSUBS 2.04307f
C126 VN.n70 VSUBS 0.849847f
C127 VN.n71 VSUBS 0.046622f
C128 VN.n72 VSUBS 0.367595f
C129 VN.n73 VSUBS 0.028521f
C130 VN.n74 VSUBS 0.028521f
C131 VN.n75 VSUBS 0.052889f
C132 VN.n76 VSUBS 0.03633f
C133 VN.n77 VSUBS 0.046588f
C134 VN.n78 VSUBS 0.028521f
C135 VN.n79 VSUBS 0.028521f
C136 VN.n80 VSUBS 0.028521f
C137 VN.n81 VSUBS 0.052889f
C138 VN.n82 VSUBS 0.039834f
C139 VN.n83 VSUBS 0.74088f
C140 VN.n84 VSUBS 0.039834f
C141 VN.n85 VSUBS 0.028521f
C142 VN.n86 VSUBS 0.028521f
C143 VN.n87 VSUBS 0.028521f
C144 VN.n88 VSUBS 0.052889f
C145 VN.n89 VSUBS 0.046588f
C146 VN.n90 VSUBS 0.03633f
C147 VN.n91 VSUBS 0.028521f
C148 VN.n92 VSUBS 0.028521f
C149 VN.n93 VSUBS 0.028521f
C150 VN.n94 VSUBS 0.052889f
C151 VN.n95 VSUBS 0.046622f
C152 VN.n96 VSUBS 0.74088f
C153 VN.n97 VSUBS 0.033045f
C154 VN.n98 VSUBS 0.028521f
C155 VN.n99 VSUBS 0.028521f
C156 VN.n100 VSUBS 0.028521f
C157 VN.n101 VSUBS 0.052889f
C158 VN.n102 VSUBS 0.054343f
C159 VN.n103 VSUBS 0.024154f
C160 VN.n104 VSUBS 0.028521f
C161 VN.n105 VSUBS 0.028521f
C162 VN.n106 VSUBS 0.028521f
C163 VN.n107 VSUBS 0.052889f
C164 VN.n108 VSUBS 0.052889f
C165 VN.n109 VSUBS 0.027301f
C166 VN.n110 VSUBS 0.046024f
C167 VN.n111 VSUBS 1.92894f
C168 B.n0 VSUBS 0.006832f
C169 B.n1 VSUBS 0.006832f
C170 B.n2 VSUBS 0.010805f
C171 B.n3 VSUBS 0.010805f
C172 B.n4 VSUBS 0.010805f
C173 B.n5 VSUBS 0.010805f
C174 B.n6 VSUBS 0.010805f
C175 B.n7 VSUBS 0.010805f
C176 B.n8 VSUBS 0.010805f
C177 B.n9 VSUBS 0.010805f
C178 B.n10 VSUBS 0.010805f
C179 B.n11 VSUBS 0.010805f
C180 B.n12 VSUBS 0.010805f
C181 B.n13 VSUBS 0.010805f
C182 B.n14 VSUBS 0.010805f
C183 B.n15 VSUBS 0.010805f
C184 B.n16 VSUBS 0.010805f
C185 B.n17 VSUBS 0.010805f
C186 B.n18 VSUBS 0.010805f
C187 B.n19 VSUBS 0.010805f
C188 B.n20 VSUBS 0.010805f
C189 B.n21 VSUBS 0.010805f
C190 B.n22 VSUBS 0.010805f
C191 B.n23 VSUBS 0.010805f
C192 B.n24 VSUBS 0.010805f
C193 B.n25 VSUBS 0.010805f
C194 B.n26 VSUBS 0.010805f
C195 B.n27 VSUBS 0.010805f
C196 B.n28 VSUBS 0.010805f
C197 B.n29 VSUBS 0.010805f
C198 B.n30 VSUBS 0.010805f
C199 B.n31 VSUBS 0.010805f
C200 B.n32 VSUBS 0.010805f
C201 B.n33 VSUBS 0.010805f
C202 B.n34 VSUBS 0.010805f
C203 B.n35 VSUBS 0.010805f
C204 B.n36 VSUBS 0.010805f
C205 B.n37 VSUBS 0.010805f
C206 B.n38 VSUBS 0.010805f
C207 B.n39 VSUBS 0.010805f
C208 B.n40 VSUBS 0.010805f
C209 B.n41 VSUBS 0.010805f
C210 B.n42 VSUBS 0.023701f
C211 B.n43 VSUBS 0.010805f
C212 B.n44 VSUBS 0.010805f
C213 B.n45 VSUBS 0.010805f
C214 B.n46 VSUBS 0.010805f
C215 B.n47 VSUBS 0.010805f
C216 B.n48 VSUBS 0.010805f
C217 B.n49 VSUBS 0.010805f
C218 B.n50 VSUBS 0.010805f
C219 B.n51 VSUBS 0.010805f
C220 B.n52 VSUBS 0.010805f
C221 B.n53 VSUBS 0.010805f
C222 B.n54 VSUBS 0.010805f
C223 B.n55 VSUBS 0.010805f
C224 B.t8 VSUBS 0.32873f
C225 B.t7 VSUBS 0.37081f
C226 B.t6 VSUBS 1.97872f
C227 B.n56 VSUBS 0.222186f
C228 B.n57 VSUBS 0.117704f
C229 B.n58 VSUBS 0.025034f
C230 B.n59 VSUBS 0.010805f
C231 B.n60 VSUBS 0.010805f
C232 B.n61 VSUBS 0.010805f
C233 B.n62 VSUBS 0.010805f
C234 B.n63 VSUBS 0.010805f
C235 B.t5 VSUBS 0.328728f
C236 B.t4 VSUBS 0.370808f
C237 B.t3 VSUBS 1.97872f
C238 B.n64 VSUBS 0.222188f
C239 B.n65 VSUBS 0.117706f
C240 B.n66 VSUBS 0.010805f
C241 B.n67 VSUBS 0.010805f
C242 B.n68 VSUBS 0.010805f
C243 B.n69 VSUBS 0.010805f
C244 B.n70 VSUBS 0.010805f
C245 B.n71 VSUBS 0.010805f
C246 B.n72 VSUBS 0.010805f
C247 B.n73 VSUBS 0.010805f
C248 B.n74 VSUBS 0.010805f
C249 B.n75 VSUBS 0.010805f
C250 B.n76 VSUBS 0.010805f
C251 B.n77 VSUBS 0.010805f
C252 B.n78 VSUBS 0.010805f
C253 B.n79 VSUBS 0.023701f
C254 B.n80 VSUBS 0.010805f
C255 B.n81 VSUBS 0.010805f
C256 B.n82 VSUBS 0.010805f
C257 B.n83 VSUBS 0.010805f
C258 B.n84 VSUBS 0.010805f
C259 B.n85 VSUBS 0.010805f
C260 B.n86 VSUBS 0.010805f
C261 B.n87 VSUBS 0.010805f
C262 B.n88 VSUBS 0.010805f
C263 B.n89 VSUBS 0.010805f
C264 B.n90 VSUBS 0.010805f
C265 B.n91 VSUBS 0.010805f
C266 B.n92 VSUBS 0.010805f
C267 B.n93 VSUBS 0.010805f
C268 B.n94 VSUBS 0.010805f
C269 B.n95 VSUBS 0.010805f
C270 B.n96 VSUBS 0.010805f
C271 B.n97 VSUBS 0.010805f
C272 B.n98 VSUBS 0.010805f
C273 B.n99 VSUBS 0.010805f
C274 B.n100 VSUBS 0.010805f
C275 B.n101 VSUBS 0.010805f
C276 B.n102 VSUBS 0.010805f
C277 B.n103 VSUBS 0.010805f
C278 B.n104 VSUBS 0.010805f
C279 B.n105 VSUBS 0.010805f
C280 B.n106 VSUBS 0.010805f
C281 B.n107 VSUBS 0.010805f
C282 B.n108 VSUBS 0.010805f
C283 B.n109 VSUBS 0.010805f
C284 B.n110 VSUBS 0.010805f
C285 B.n111 VSUBS 0.010805f
C286 B.n112 VSUBS 0.010805f
C287 B.n113 VSUBS 0.010805f
C288 B.n114 VSUBS 0.010805f
C289 B.n115 VSUBS 0.010805f
C290 B.n116 VSUBS 0.010805f
C291 B.n117 VSUBS 0.010805f
C292 B.n118 VSUBS 0.010805f
C293 B.n119 VSUBS 0.010805f
C294 B.n120 VSUBS 0.010805f
C295 B.n121 VSUBS 0.010805f
C296 B.n122 VSUBS 0.010805f
C297 B.n123 VSUBS 0.010805f
C298 B.n124 VSUBS 0.010805f
C299 B.n125 VSUBS 0.010805f
C300 B.n126 VSUBS 0.010805f
C301 B.n127 VSUBS 0.010805f
C302 B.n128 VSUBS 0.010805f
C303 B.n129 VSUBS 0.010805f
C304 B.n130 VSUBS 0.010805f
C305 B.n131 VSUBS 0.010805f
C306 B.n132 VSUBS 0.010805f
C307 B.n133 VSUBS 0.010805f
C308 B.n134 VSUBS 0.010805f
C309 B.n135 VSUBS 0.010805f
C310 B.n136 VSUBS 0.010805f
C311 B.n137 VSUBS 0.010805f
C312 B.n138 VSUBS 0.010805f
C313 B.n139 VSUBS 0.010805f
C314 B.n140 VSUBS 0.010805f
C315 B.n141 VSUBS 0.010805f
C316 B.n142 VSUBS 0.010805f
C317 B.n143 VSUBS 0.010805f
C318 B.n144 VSUBS 0.010805f
C319 B.n145 VSUBS 0.010805f
C320 B.n146 VSUBS 0.010805f
C321 B.n147 VSUBS 0.010805f
C322 B.n148 VSUBS 0.010805f
C323 B.n149 VSUBS 0.010805f
C324 B.n150 VSUBS 0.010805f
C325 B.n151 VSUBS 0.010805f
C326 B.n152 VSUBS 0.010805f
C327 B.n153 VSUBS 0.010805f
C328 B.n154 VSUBS 0.010805f
C329 B.n155 VSUBS 0.010805f
C330 B.n156 VSUBS 0.010805f
C331 B.n157 VSUBS 0.010805f
C332 B.n158 VSUBS 0.010805f
C333 B.n159 VSUBS 0.010805f
C334 B.n160 VSUBS 0.023701f
C335 B.n161 VSUBS 0.010805f
C336 B.n162 VSUBS 0.010805f
C337 B.n163 VSUBS 0.010805f
C338 B.n164 VSUBS 0.010805f
C339 B.n165 VSUBS 0.010805f
C340 B.n166 VSUBS 0.010805f
C341 B.n167 VSUBS 0.010805f
C342 B.n168 VSUBS 0.010805f
C343 B.n169 VSUBS 0.010805f
C344 B.n170 VSUBS 0.010805f
C345 B.n171 VSUBS 0.010805f
C346 B.n172 VSUBS 0.010805f
C347 B.n173 VSUBS 0.010805f
C348 B.t1 VSUBS 0.328728f
C349 B.t2 VSUBS 0.370808f
C350 B.t0 VSUBS 1.97872f
C351 B.n174 VSUBS 0.222188f
C352 B.n175 VSUBS 0.117706f
C353 B.n176 VSUBS 0.025034f
C354 B.n177 VSUBS 0.010805f
C355 B.n178 VSUBS 0.010805f
C356 B.n179 VSUBS 0.010805f
C357 B.n180 VSUBS 0.010805f
C358 B.n181 VSUBS 0.010805f
C359 B.t10 VSUBS 0.32873f
C360 B.t11 VSUBS 0.37081f
C361 B.t9 VSUBS 1.97872f
C362 B.n182 VSUBS 0.222186f
C363 B.n183 VSUBS 0.117704f
C364 B.n184 VSUBS 0.010805f
C365 B.n185 VSUBS 0.010805f
C366 B.n186 VSUBS 0.010805f
C367 B.n187 VSUBS 0.010805f
C368 B.n188 VSUBS 0.010805f
C369 B.n189 VSUBS 0.010805f
C370 B.n190 VSUBS 0.010805f
C371 B.n191 VSUBS 0.010805f
C372 B.n192 VSUBS 0.010805f
C373 B.n193 VSUBS 0.010805f
C374 B.n194 VSUBS 0.010805f
C375 B.n195 VSUBS 0.010805f
C376 B.n196 VSUBS 0.010805f
C377 B.n197 VSUBS 0.023701f
C378 B.n198 VSUBS 0.010805f
C379 B.n199 VSUBS 0.010805f
C380 B.n200 VSUBS 0.010805f
C381 B.n201 VSUBS 0.010805f
C382 B.n202 VSUBS 0.010805f
C383 B.n203 VSUBS 0.010805f
C384 B.n204 VSUBS 0.010805f
C385 B.n205 VSUBS 0.010805f
C386 B.n206 VSUBS 0.010805f
C387 B.n207 VSUBS 0.010805f
C388 B.n208 VSUBS 0.010805f
C389 B.n209 VSUBS 0.010805f
C390 B.n210 VSUBS 0.010805f
C391 B.n211 VSUBS 0.010805f
C392 B.n212 VSUBS 0.010805f
C393 B.n213 VSUBS 0.010805f
C394 B.n214 VSUBS 0.010805f
C395 B.n215 VSUBS 0.010805f
C396 B.n216 VSUBS 0.010805f
C397 B.n217 VSUBS 0.010805f
C398 B.n218 VSUBS 0.010805f
C399 B.n219 VSUBS 0.010805f
C400 B.n220 VSUBS 0.010805f
C401 B.n221 VSUBS 0.010805f
C402 B.n222 VSUBS 0.010805f
C403 B.n223 VSUBS 0.010805f
C404 B.n224 VSUBS 0.010805f
C405 B.n225 VSUBS 0.010805f
C406 B.n226 VSUBS 0.010805f
C407 B.n227 VSUBS 0.010805f
C408 B.n228 VSUBS 0.010805f
C409 B.n229 VSUBS 0.010805f
C410 B.n230 VSUBS 0.010805f
C411 B.n231 VSUBS 0.010805f
C412 B.n232 VSUBS 0.010805f
C413 B.n233 VSUBS 0.010805f
C414 B.n234 VSUBS 0.010805f
C415 B.n235 VSUBS 0.010805f
C416 B.n236 VSUBS 0.010805f
C417 B.n237 VSUBS 0.010805f
C418 B.n238 VSUBS 0.010805f
C419 B.n239 VSUBS 0.010805f
C420 B.n240 VSUBS 0.010805f
C421 B.n241 VSUBS 0.010805f
C422 B.n242 VSUBS 0.010805f
C423 B.n243 VSUBS 0.010805f
C424 B.n244 VSUBS 0.010805f
C425 B.n245 VSUBS 0.010805f
C426 B.n246 VSUBS 0.010805f
C427 B.n247 VSUBS 0.010805f
C428 B.n248 VSUBS 0.010805f
C429 B.n249 VSUBS 0.010805f
C430 B.n250 VSUBS 0.010805f
C431 B.n251 VSUBS 0.010805f
C432 B.n252 VSUBS 0.010805f
C433 B.n253 VSUBS 0.010805f
C434 B.n254 VSUBS 0.010805f
C435 B.n255 VSUBS 0.010805f
C436 B.n256 VSUBS 0.010805f
C437 B.n257 VSUBS 0.010805f
C438 B.n258 VSUBS 0.010805f
C439 B.n259 VSUBS 0.010805f
C440 B.n260 VSUBS 0.010805f
C441 B.n261 VSUBS 0.010805f
C442 B.n262 VSUBS 0.010805f
C443 B.n263 VSUBS 0.010805f
C444 B.n264 VSUBS 0.010805f
C445 B.n265 VSUBS 0.010805f
C446 B.n266 VSUBS 0.010805f
C447 B.n267 VSUBS 0.010805f
C448 B.n268 VSUBS 0.010805f
C449 B.n269 VSUBS 0.010805f
C450 B.n270 VSUBS 0.010805f
C451 B.n271 VSUBS 0.010805f
C452 B.n272 VSUBS 0.010805f
C453 B.n273 VSUBS 0.010805f
C454 B.n274 VSUBS 0.010805f
C455 B.n275 VSUBS 0.010805f
C456 B.n276 VSUBS 0.010805f
C457 B.n277 VSUBS 0.010805f
C458 B.n278 VSUBS 0.010805f
C459 B.n279 VSUBS 0.010805f
C460 B.n280 VSUBS 0.010805f
C461 B.n281 VSUBS 0.010805f
C462 B.n282 VSUBS 0.010805f
C463 B.n283 VSUBS 0.010805f
C464 B.n284 VSUBS 0.010805f
C465 B.n285 VSUBS 0.010805f
C466 B.n286 VSUBS 0.010805f
C467 B.n287 VSUBS 0.010805f
C468 B.n288 VSUBS 0.010805f
C469 B.n289 VSUBS 0.010805f
C470 B.n290 VSUBS 0.010805f
C471 B.n291 VSUBS 0.010805f
C472 B.n292 VSUBS 0.010805f
C473 B.n293 VSUBS 0.010805f
C474 B.n294 VSUBS 0.010805f
C475 B.n295 VSUBS 0.010805f
C476 B.n296 VSUBS 0.010805f
C477 B.n297 VSUBS 0.010805f
C478 B.n298 VSUBS 0.010805f
C479 B.n299 VSUBS 0.010805f
C480 B.n300 VSUBS 0.010805f
C481 B.n301 VSUBS 0.010805f
C482 B.n302 VSUBS 0.010805f
C483 B.n303 VSUBS 0.010805f
C484 B.n304 VSUBS 0.010805f
C485 B.n305 VSUBS 0.010805f
C486 B.n306 VSUBS 0.010805f
C487 B.n307 VSUBS 0.010805f
C488 B.n308 VSUBS 0.010805f
C489 B.n309 VSUBS 0.010805f
C490 B.n310 VSUBS 0.010805f
C491 B.n311 VSUBS 0.010805f
C492 B.n312 VSUBS 0.010805f
C493 B.n313 VSUBS 0.010805f
C494 B.n314 VSUBS 0.010805f
C495 B.n315 VSUBS 0.010805f
C496 B.n316 VSUBS 0.010805f
C497 B.n317 VSUBS 0.010805f
C498 B.n318 VSUBS 0.010805f
C499 B.n319 VSUBS 0.010805f
C500 B.n320 VSUBS 0.010805f
C501 B.n321 VSUBS 0.010805f
C502 B.n322 VSUBS 0.010805f
C503 B.n323 VSUBS 0.010805f
C504 B.n324 VSUBS 0.010805f
C505 B.n325 VSUBS 0.010805f
C506 B.n326 VSUBS 0.010805f
C507 B.n327 VSUBS 0.010805f
C508 B.n328 VSUBS 0.010805f
C509 B.n329 VSUBS 0.010805f
C510 B.n330 VSUBS 0.010805f
C511 B.n331 VSUBS 0.010805f
C512 B.n332 VSUBS 0.010805f
C513 B.n333 VSUBS 0.010805f
C514 B.n334 VSUBS 0.010805f
C515 B.n335 VSUBS 0.010805f
C516 B.n336 VSUBS 0.010805f
C517 B.n337 VSUBS 0.010805f
C518 B.n338 VSUBS 0.010805f
C519 B.n339 VSUBS 0.010805f
C520 B.n340 VSUBS 0.010805f
C521 B.n341 VSUBS 0.010805f
C522 B.n342 VSUBS 0.010805f
C523 B.n343 VSUBS 0.010805f
C524 B.n344 VSUBS 0.010805f
C525 B.n345 VSUBS 0.010805f
C526 B.n346 VSUBS 0.010805f
C527 B.n347 VSUBS 0.010805f
C528 B.n348 VSUBS 0.010805f
C529 B.n349 VSUBS 0.010805f
C530 B.n350 VSUBS 0.010805f
C531 B.n351 VSUBS 0.010805f
C532 B.n352 VSUBS 0.010805f
C533 B.n353 VSUBS 0.010805f
C534 B.n354 VSUBS 0.010805f
C535 B.n355 VSUBS 0.010805f
C536 B.n356 VSUBS 0.023701f
C537 B.n357 VSUBS 0.025239f
C538 B.n358 VSUBS 0.025239f
C539 B.n359 VSUBS 0.010805f
C540 B.n360 VSUBS 0.010805f
C541 B.n361 VSUBS 0.010805f
C542 B.n362 VSUBS 0.010805f
C543 B.n363 VSUBS 0.010805f
C544 B.n364 VSUBS 0.010805f
C545 B.n365 VSUBS 0.010805f
C546 B.n366 VSUBS 0.010805f
C547 B.n367 VSUBS 0.010805f
C548 B.n368 VSUBS 0.010805f
C549 B.n369 VSUBS 0.010805f
C550 B.n370 VSUBS 0.010805f
C551 B.n371 VSUBS 0.010805f
C552 B.n372 VSUBS 0.010805f
C553 B.n373 VSUBS 0.010805f
C554 B.n374 VSUBS 0.010805f
C555 B.n375 VSUBS 0.010805f
C556 B.n376 VSUBS 0.010805f
C557 B.n377 VSUBS 0.010805f
C558 B.n378 VSUBS 0.010805f
C559 B.n379 VSUBS 0.010805f
C560 B.n380 VSUBS 0.010805f
C561 B.n381 VSUBS 0.010805f
C562 B.n382 VSUBS 0.010805f
C563 B.n383 VSUBS 0.010805f
C564 B.n384 VSUBS 0.010805f
C565 B.n385 VSUBS 0.010805f
C566 B.n386 VSUBS 0.010805f
C567 B.n387 VSUBS 0.010805f
C568 B.n388 VSUBS 0.010805f
C569 B.n389 VSUBS 0.010805f
C570 B.n390 VSUBS 0.010805f
C571 B.n391 VSUBS 0.010805f
C572 B.n392 VSUBS 0.010805f
C573 B.n393 VSUBS 0.010805f
C574 B.n394 VSUBS 0.010805f
C575 B.n395 VSUBS 0.010805f
C576 B.n396 VSUBS 0.010805f
C577 B.n397 VSUBS 0.010169f
C578 B.n398 VSUBS 0.025034f
C579 B.n399 VSUBS 0.006038f
C580 B.n400 VSUBS 0.010805f
C581 B.n401 VSUBS 0.010805f
C582 B.n402 VSUBS 0.010805f
C583 B.n403 VSUBS 0.010805f
C584 B.n404 VSUBS 0.010805f
C585 B.n405 VSUBS 0.010805f
C586 B.n406 VSUBS 0.010805f
C587 B.n407 VSUBS 0.010805f
C588 B.n408 VSUBS 0.010805f
C589 B.n409 VSUBS 0.010805f
C590 B.n410 VSUBS 0.010805f
C591 B.n411 VSUBS 0.010805f
C592 B.n412 VSUBS 0.006038f
C593 B.n413 VSUBS 0.010805f
C594 B.n414 VSUBS 0.010805f
C595 B.n415 VSUBS 0.010169f
C596 B.n416 VSUBS 0.010805f
C597 B.n417 VSUBS 0.010805f
C598 B.n418 VSUBS 0.010805f
C599 B.n419 VSUBS 0.010805f
C600 B.n420 VSUBS 0.010805f
C601 B.n421 VSUBS 0.010805f
C602 B.n422 VSUBS 0.010805f
C603 B.n423 VSUBS 0.010805f
C604 B.n424 VSUBS 0.010805f
C605 B.n425 VSUBS 0.010805f
C606 B.n426 VSUBS 0.010805f
C607 B.n427 VSUBS 0.010805f
C608 B.n428 VSUBS 0.010805f
C609 B.n429 VSUBS 0.010805f
C610 B.n430 VSUBS 0.010805f
C611 B.n431 VSUBS 0.010805f
C612 B.n432 VSUBS 0.010805f
C613 B.n433 VSUBS 0.010805f
C614 B.n434 VSUBS 0.010805f
C615 B.n435 VSUBS 0.010805f
C616 B.n436 VSUBS 0.010805f
C617 B.n437 VSUBS 0.010805f
C618 B.n438 VSUBS 0.010805f
C619 B.n439 VSUBS 0.010805f
C620 B.n440 VSUBS 0.010805f
C621 B.n441 VSUBS 0.010805f
C622 B.n442 VSUBS 0.010805f
C623 B.n443 VSUBS 0.010805f
C624 B.n444 VSUBS 0.010805f
C625 B.n445 VSUBS 0.010805f
C626 B.n446 VSUBS 0.010805f
C627 B.n447 VSUBS 0.010805f
C628 B.n448 VSUBS 0.010805f
C629 B.n449 VSUBS 0.010805f
C630 B.n450 VSUBS 0.010805f
C631 B.n451 VSUBS 0.010805f
C632 B.n452 VSUBS 0.010805f
C633 B.n453 VSUBS 0.025239f
C634 B.n454 VSUBS 0.025239f
C635 B.n455 VSUBS 0.023701f
C636 B.n456 VSUBS 0.010805f
C637 B.n457 VSUBS 0.010805f
C638 B.n458 VSUBS 0.010805f
C639 B.n459 VSUBS 0.010805f
C640 B.n460 VSUBS 0.010805f
C641 B.n461 VSUBS 0.010805f
C642 B.n462 VSUBS 0.010805f
C643 B.n463 VSUBS 0.010805f
C644 B.n464 VSUBS 0.010805f
C645 B.n465 VSUBS 0.010805f
C646 B.n466 VSUBS 0.010805f
C647 B.n467 VSUBS 0.010805f
C648 B.n468 VSUBS 0.010805f
C649 B.n469 VSUBS 0.010805f
C650 B.n470 VSUBS 0.010805f
C651 B.n471 VSUBS 0.010805f
C652 B.n472 VSUBS 0.010805f
C653 B.n473 VSUBS 0.010805f
C654 B.n474 VSUBS 0.010805f
C655 B.n475 VSUBS 0.010805f
C656 B.n476 VSUBS 0.010805f
C657 B.n477 VSUBS 0.010805f
C658 B.n478 VSUBS 0.010805f
C659 B.n479 VSUBS 0.010805f
C660 B.n480 VSUBS 0.010805f
C661 B.n481 VSUBS 0.010805f
C662 B.n482 VSUBS 0.010805f
C663 B.n483 VSUBS 0.010805f
C664 B.n484 VSUBS 0.010805f
C665 B.n485 VSUBS 0.010805f
C666 B.n486 VSUBS 0.010805f
C667 B.n487 VSUBS 0.010805f
C668 B.n488 VSUBS 0.010805f
C669 B.n489 VSUBS 0.010805f
C670 B.n490 VSUBS 0.010805f
C671 B.n491 VSUBS 0.010805f
C672 B.n492 VSUBS 0.010805f
C673 B.n493 VSUBS 0.010805f
C674 B.n494 VSUBS 0.010805f
C675 B.n495 VSUBS 0.010805f
C676 B.n496 VSUBS 0.010805f
C677 B.n497 VSUBS 0.010805f
C678 B.n498 VSUBS 0.010805f
C679 B.n499 VSUBS 0.010805f
C680 B.n500 VSUBS 0.010805f
C681 B.n501 VSUBS 0.010805f
C682 B.n502 VSUBS 0.010805f
C683 B.n503 VSUBS 0.010805f
C684 B.n504 VSUBS 0.010805f
C685 B.n505 VSUBS 0.010805f
C686 B.n506 VSUBS 0.010805f
C687 B.n507 VSUBS 0.010805f
C688 B.n508 VSUBS 0.010805f
C689 B.n509 VSUBS 0.010805f
C690 B.n510 VSUBS 0.010805f
C691 B.n511 VSUBS 0.010805f
C692 B.n512 VSUBS 0.010805f
C693 B.n513 VSUBS 0.010805f
C694 B.n514 VSUBS 0.010805f
C695 B.n515 VSUBS 0.010805f
C696 B.n516 VSUBS 0.010805f
C697 B.n517 VSUBS 0.010805f
C698 B.n518 VSUBS 0.010805f
C699 B.n519 VSUBS 0.010805f
C700 B.n520 VSUBS 0.010805f
C701 B.n521 VSUBS 0.010805f
C702 B.n522 VSUBS 0.010805f
C703 B.n523 VSUBS 0.010805f
C704 B.n524 VSUBS 0.010805f
C705 B.n525 VSUBS 0.010805f
C706 B.n526 VSUBS 0.010805f
C707 B.n527 VSUBS 0.010805f
C708 B.n528 VSUBS 0.010805f
C709 B.n529 VSUBS 0.010805f
C710 B.n530 VSUBS 0.010805f
C711 B.n531 VSUBS 0.010805f
C712 B.n532 VSUBS 0.010805f
C713 B.n533 VSUBS 0.010805f
C714 B.n534 VSUBS 0.010805f
C715 B.n535 VSUBS 0.010805f
C716 B.n536 VSUBS 0.010805f
C717 B.n537 VSUBS 0.010805f
C718 B.n538 VSUBS 0.010805f
C719 B.n539 VSUBS 0.010805f
C720 B.n540 VSUBS 0.010805f
C721 B.n541 VSUBS 0.010805f
C722 B.n542 VSUBS 0.010805f
C723 B.n543 VSUBS 0.010805f
C724 B.n544 VSUBS 0.010805f
C725 B.n545 VSUBS 0.010805f
C726 B.n546 VSUBS 0.010805f
C727 B.n547 VSUBS 0.010805f
C728 B.n548 VSUBS 0.010805f
C729 B.n549 VSUBS 0.010805f
C730 B.n550 VSUBS 0.010805f
C731 B.n551 VSUBS 0.010805f
C732 B.n552 VSUBS 0.010805f
C733 B.n553 VSUBS 0.010805f
C734 B.n554 VSUBS 0.010805f
C735 B.n555 VSUBS 0.010805f
C736 B.n556 VSUBS 0.010805f
C737 B.n557 VSUBS 0.010805f
C738 B.n558 VSUBS 0.010805f
C739 B.n559 VSUBS 0.010805f
C740 B.n560 VSUBS 0.010805f
C741 B.n561 VSUBS 0.010805f
C742 B.n562 VSUBS 0.010805f
C743 B.n563 VSUBS 0.010805f
C744 B.n564 VSUBS 0.010805f
C745 B.n565 VSUBS 0.010805f
C746 B.n566 VSUBS 0.010805f
C747 B.n567 VSUBS 0.010805f
C748 B.n568 VSUBS 0.010805f
C749 B.n569 VSUBS 0.010805f
C750 B.n570 VSUBS 0.010805f
C751 B.n571 VSUBS 0.010805f
C752 B.n572 VSUBS 0.010805f
C753 B.n573 VSUBS 0.010805f
C754 B.n574 VSUBS 0.010805f
C755 B.n575 VSUBS 0.010805f
C756 B.n576 VSUBS 0.010805f
C757 B.n577 VSUBS 0.010805f
C758 B.n578 VSUBS 0.010805f
C759 B.n579 VSUBS 0.010805f
C760 B.n580 VSUBS 0.010805f
C761 B.n581 VSUBS 0.010805f
C762 B.n582 VSUBS 0.010805f
C763 B.n583 VSUBS 0.010805f
C764 B.n584 VSUBS 0.010805f
C765 B.n585 VSUBS 0.010805f
C766 B.n586 VSUBS 0.010805f
C767 B.n587 VSUBS 0.010805f
C768 B.n588 VSUBS 0.010805f
C769 B.n589 VSUBS 0.010805f
C770 B.n590 VSUBS 0.010805f
C771 B.n591 VSUBS 0.010805f
C772 B.n592 VSUBS 0.010805f
C773 B.n593 VSUBS 0.010805f
C774 B.n594 VSUBS 0.010805f
C775 B.n595 VSUBS 0.010805f
C776 B.n596 VSUBS 0.010805f
C777 B.n597 VSUBS 0.010805f
C778 B.n598 VSUBS 0.010805f
C779 B.n599 VSUBS 0.010805f
C780 B.n600 VSUBS 0.010805f
C781 B.n601 VSUBS 0.010805f
C782 B.n602 VSUBS 0.010805f
C783 B.n603 VSUBS 0.010805f
C784 B.n604 VSUBS 0.010805f
C785 B.n605 VSUBS 0.010805f
C786 B.n606 VSUBS 0.010805f
C787 B.n607 VSUBS 0.010805f
C788 B.n608 VSUBS 0.010805f
C789 B.n609 VSUBS 0.010805f
C790 B.n610 VSUBS 0.010805f
C791 B.n611 VSUBS 0.010805f
C792 B.n612 VSUBS 0.010805f
C793 B.n613 VSUBS 0.010805f
C794 B.n614 VSUBS 0.010805f
C795 B.n615 VSUBS 0.010805f
C796 B.n616 VSUBS 0.010805f
C797 B.n617 VSUBS 0.010805f
C798 B.n618 VSUBS 0.010805f
C799 B.n619 VSUBS 0.010805f
C800 B.n620 VSUBS 0.010805f
C801 B.n621 VSUBS 0.010805f
C802 B.n622 VSUBS 0.010805f
C803 B.n623 VSUBS 0.010805f
C804 B.n624 VSUBS 0.010805f
C805 B.n625 VSUBS 0.010805f
C806 B.n626 VSUBS 0.010805f
C807 B.n627 VSUBS 0.010805f
C808 B.n628 VSUBS 0.010805f
C809 B.n629 VSUBS 0.010805f
C810 B.n630 VSUBS 0.010805f
C811 B.n631 VSUBS 0.010805f
C812 B.n632 VSUBS 0.010805f
C813 B.n633 VSUBS 0.010805f
C814 B.n634 VSUBS 0.010805f
C815 B.n635 VSUBS 0.010805f
C816 B.n636 VSUBS 0.010805f
C817 B.n637 VSUBS 0.010805f
C818 B.n638 VSUBS 0.010805f
C819 B.n639 VSUBS 0.010805f
C820 B.n640 VSUBS 0.010805f
C821 B.n641 VSUBS 0.010805f
C822 B.n642 VSUBS 0.010805f
C823 B.n643 VSUBS 0.010805f
C824 B.n644 VSUBS 0.010805f
C825 B.n645 VSUBS 0.010805f
C826 B.n646 VSUBS 0.010805f
C827 B.n647 VSUBS 0.010805f
C828 B.n648 VSUBS 0.010805f
C829 B.n649 VSUBS 0.010805f
C830 B.n650 VSUBS 0.010805f
C831 B.n651 VSUBS 0.010805f
C832 B.n652 VSUBS 0.010805f
C833 B.n653 VSUBS 0.010805f
C834 B.n654 VSUBS 0.010805f
C835 B.n655 VSUBS 0.010805f
C836 B.n656 VSUBS 0.010805f
C837 B.n657 VSUBS 0.010805f
C838 B.n658 VSUBS 0.010805f
C839 B.n659 VSUBS 0.010805f
C840 B.n660 VSUBS 0.010805f
C841 B.n661 VSUBS 0.010805f
C842 B.n662 VSUBS 0.010805f
C843 B.n663 VSUBS 0.010805f
C844 B.n664 VSUBS 0.010805f
C845 B.n665 VSUBS 0.010805f
C846 B.n666 VSUBS 0.010805f
C847 B.n667 VSUBS 0.010805f
C848 B.n668 VSUBS 0.010805f
C849 B.n669 VSUBS 0.010805f
C850 B.n670 VSUBS 0.010805f
C851 B.n671 VSUBS 0.010805f
C852 B.n672 VSUBS 0.010805f
C853 B.n673 VSUBS 0.010805f
C854 B.n674 VSUBS 0.010805f
C855 B.n675 VSUBS 0.010805f
C856 B.n676 VSUBS 0.010805f
C857 B.n677 VSUBS 0.010805f
C858 B.n678 VSUBS 0.010805f
C859 B.n679 VSUBS 0.010805f
C860 B.n680 VSUBS 0.010805f
C861 B.n681 VSUBS 0.010805f
C862 B.n682 VSUBS 0.010805f
C863 B.n683 VSUBS 0.010805f
C864 B.n684 VSUBS 0.010805f
C865 B.n685 VSUBS 0.010805f
C866 B.n686 VSUBS 0.010805f
C867 B.n687 VSUBS 0.010805f
C868 B.n688 VSUBS 0.010805f
C869 B.n689 VSUBS 0.010805f
C870 B.n690 VSUBS 0.010805f
C871 B.n691 VSUBS 0.010805f
C872 B.n692 VSUBS 0.010805f
C873 B.n693 VSUBS 0.010805f
C874 B.n694 VSUBS 0.010805f
C875 B.n695 VSUBS 0.010805f
C876 B.n696 VSUBS 0.010805f
C877 B.n697 VSUBS 0.010805f
C878 B.n698 VSUBS 0.025043f
C879 B.n699 VSUBS 0.023897f
C880 B.n700 VSUBS 0.025239f
C881 B.n701 VSUBS 0.010805f
C882 B.n702 VSUBS 0.010805f
C883 B.n703 VSUBS 0.010805f
C884 B.n704 VSUBS 0.010805f
C885 B.n705 VSUBS 0.010805f
C886 B.n706 VSUBS 0.010805f
C887 B.n707 VSUBS 0.010805f
C888 B.n708 VSUBS 0.010805f
C889 B.n709 VSUBS 0.010805f
C890 B.n710 VSUBS 0.010805f
C891 B.n711 VSUBS 0.010805f
C892 B.n712 VSUBS 0.010805f
C893 B.n713 VSUBS 0.010805f
C894 B.n714 VSUBS 0.010805f
C895 B.n715 VSUBS 0.010805f
C896 B.n716 VSUBS 0.010805f
C897 B.n717 VSUBS 0.010805f
C898 B.n718 VSUBS 0.010805f
C899 B.n719 VSUBS 0.010805f
C900 B.n720 VSUBS 0.010805f
C901 B.n721 VSUBS 0.010805f
C902 B.n722 VSUBS 0.010805f
C903 B.n723 VSUBS 0.010805f
C904 B.n724 VSUBS 0.010805f
C905 B.n725 VSUBS 0.010805f
C906 B.n726 VSUBS 0.010805f
C907 B.n727 VSUBS 0.010805f
C908 B.n728 VSUBS 0.010805f
C909 B.n729 VSUBS 0.010805f
C910 B.n730 VSUBS 0.010805f
C911 B.n731 VSUBS 0.010805f
C912 B.n732 VSUBS 0.010805f
C913 B.n733 VSUBS 0.010805f
C914 B.n734 VSUBS 0.010805f
C915 B.n735 VSUBS 0.010805f
C916 B.n736 VSUBS 0.010805f
C917 B.n737 VSUBS 0.010805f
C918 B.n738 VSUBS 0.010805f
C919 B.n739 VSUBS 0.010169f
C920 B.n740 VSUBS 0.025034f
C921 B.n741 VSUBS 0.006038f
C922 B.n742 VSUBS 0.010805f
C923 B.n743 VSUBS 0.010805f
C924 B.n744 VSUBS 0.010805f
C925 B.n745 VSUBS 0.010805f
C926 B.n746 VSUBS 0.010805f
C927 B.n747 VSUBS 0.010805f
C928 B.n748 VSUBS 0.010805f
C929 B.n749 VSUBS 0.010805f
C930 B.n750 VSUBS 0.010805f
C931 B.n751 VSUBS 0.010805f
C932 B.n752 VSUBS 0.010805f
C933 B.n753 VSUBS 0.010805f
C934 B.n754 VSUBS 0.006038f
C935 B.n755 VSUBS 0.010805f
C936 B.n756 VSUBS 0.010805f
C937 B.n757 VSUBS 0.010169f
C938 B.n758 VSUBS 0.010805f
C939 B.n759 VSUBS 0.010805f
C940 B.n760 VSUBS 0.010805f
C941 B.n761 VSUBS 0.010805f
C942 B.n762 VSUBS 0.010805f
C943 B.n763 VSUBS 0.010805f
C944 B.n764 VSUBS 0.010805f
C945 B.n765 VSUBS 0.010805f
C946 B.n766 VSUBS 0.010805f
C947 B.n767 VSUBS 0.010805f
C948 B.n768 VSUBS 0.010805f
C949 B.n769 VSUBS 0.010805f
C950 B.n770 VSUBS 0.010805f
C951 B.n771 VSUBS 0.010805f
C952 B.n772 VSUBS 0.010805f
C953 B.n773 VSUBS 0.010805f
C954 B.n774 VSUBS 0.010805f
C955 B.n775 VSUBS 0.010805f
C956 B.n776 VSUBS 0.010805f
C957 B.n777 VSUBS 0.010805f
C958 B.n778 VSUBS 0.010805f
C959 B.n779 VSUBS 0.010805f
C960 B.n780 VSUBS 0.010805f
C961 B.n781 VSUBS 0.010805f
C962 B.n782 VSUBS 0.010805f
C963 B.n783 VSUBS 0.010805f
C964 B.n784 VSUBS 0.010805f
C965 B.n785 VSUBS 0.010805f
C966 B.n786 VSUBS 0.010805f
C967 B.n787 VSUBS 0.010805f
C968 B.n788 VSUBS 0.010805f
C969 B.n789 VSUBS 0.010805f
C970 B.n790 VSUBS 0.010805f
C971 B.n791 VSUBS 0.010805f
C972 B.n792 VSUBS 0.010805f
C973 B.n793 VSUBS 0.010805f
C974 B.n794 VSUBS 0.010805f
C975 B.n795 VSUBS 0.025239f
C976 B.n796 VSUBS 0.025239f
C977 B.n797 VSUBS 0.023701f
C978 B.n798 VSUBS 0.010805f
C979 B.n799 VSUBS 0.010805f
C980 B.n800 VSUBS 0.010805f
C981 B.n801 VSUBS 0.010805f
C982 B.n802 VSUBS 0.010805f
C983 B.n803 VSUBS 0.010805f
C984 B.n804 VSUBS 0.010805f
C985 B.n805 VSUBS 0.010805f
C986 B.n806 VSUBS 0.010805f
C987 B.n807 VSUBS 0.010805f
C988 B.n808 VSUBS 0.010805f
C989 B.n809 VSUBS 0.010805f
C990 B.n810 VSUBS 0.010805f
C991 B.n811 VSUBS 0.010805f
C992 B.n812 VSUBS 0.010805f
C993 B.n813 VSUBS 0.010805f
C994 B.n814 VSUBS 0.010805f
C995 B.n815 VSUBS 0.010805f
C996 B.n816 VSUBS 0.010805f
C997 B.n817 VSUBS 0.010805f
C998 B.n818 VSUBS 0.010805f
C999 B.n819 VSUBS 0.010805f
C1000 B.n820 VSUBS 0.010805f
C1001 B.n821 VSUBS 0.010805f
C1002 B.n822 VSUBS 0.010805f
C1003 B.n823 VSUBS 0.010805f
C1004 B.n824 VSUBS 0.010805f
C1005 B.n825 VSUBS 0.010805f
C1006 B.n826 VSUBS 0.010805f
C1007 B.n827 VSUBS 0.010805f
C1008 B.n828 VSUBS 0.010805f
C1009 B.n829 VSUBS 0.010805f
C1010 B.n830 VSUBS 0.010805f
C1011 B.n831 VSUBS 0.010805f
C1012 B.n832 VSUBS 0.010805f
C1013 B.n833 VSUBS 0.010805f
C1014 B.n834 VSUBS 0.010805f
C1015 B.n835 VSUBS 0.010805f
C1016 B.n836 VSUBS 0.010805f
C1017 B.n837 VSUBS 0.010805f
C1018 B.n838 VSUBS 0.010805f
C1019 B.n839 VSUBS 0.010805f
C1020 B.n840 VSUBS 0.010805f
C1021 B.n841 VSUBS 0.010805f
C1022 B.n842 VSUBS 0.010805f
C1023 B.n843 VSUBS 0.010805f
C1024 B.n844 VSUBS 0.010805f
C1025 B.n845 VSUBS 0.010805f
C1026 B.n846 VSUBS 0.010805f
C1027 B.n847 VSUBS 0.010805f
C1028 B.n848 VSUBS 0.010805f
C1029 B.n849 VSUBS 0.010805f
C1030 B.n850 VSUBS 0.010805f
C1031 B.n851 VSUBS 0.010805f
C1032 B.n852 VSUBS 0.010805f
C1033 B.n853 VSUBS 0.010805f
C1034 B.n854 VSUBS 0.010805f
C1035 B.n855 VSUBS 0.010805f
C1036 B.n856 VSUBS 0.010805f
C1037 B.n857 VSUBS 0.010805f
C1038 B.n858 VSUBS 0.010805f
C1039 B.n859 VSUBS 0.010805f
C1040 B.n860 VSUBS 0.010805f
C1041 B.n861 VSUBS 0.010805f
C1042 B.n862 VSUBS 0.010805f
C1043 B.n863 VSUBS 0.010805f
C1044 B.n864 VSUBS 0.010805f
C1045 B.n865 VSUBS 0.010805f
C1046 B.n866 VSUBS 0.010805f
C1047 B.n867 VSUBS 0.010805f
C1048 B.n868 VSUBS 0.010805f
C1049 B.n869 VSUBS 0.010805f
C1050 B.n870 VSUBS 0.010805f
C1051 B.n871 VSUBS 0.010805f
C1052 B.n872 VSUBS 0.010805f
C1053 B.n873 VSUBS 0.010805f
C1054 B.n874 VSUBS 0.010805f
C1055 B.n875 VSUBS 0.010805f
C1056 B.n876 VSUBS 0.010805f
C1057 B.n877 VSUBS 0.010805f
C1058 B.n878 VSUBS 0.010805f
C1059 B.n879 VSUBS 0.010805f
C1060 B.n880 VSUBS 0.010805f
C1061 B.n881 VSUBS 0.010805f
C1062 B.n882 VSUBS 0.010805f
C1063 B.n883 VSUBS 0.010805f
C1064 B.n884 VSUBS 0.010805f
C1065 B.n885 VSUBS 0.010805f
C1066 B.n886 VSUBS 0.010805f
C1067 B.n887 VSUBS 0.010805f
C1068 B.n888 VSUBS 0.010805f
C1069 B.n889 VSUBS 0.010805f
C1070 B.n890 VSUBS 0.010805f
C1071 B.n891 VSUBS 0.010805f
C1072 B.n892 VSUBS 0.010805f
C1073 B.n893 VSUBS 0.010805f
C1074 B.n894 VSUBS 0.010805f
C1075 B.n895 VSUBS 0.010805f
C1076 B.n896 VSUBS 0.010805f
C1077 B.n897 VSUBS 0.010805f
C1078 B.n898 VSUBS 0.010805f
C1079 B.n899 VSUBS 0.010805f
C1080 B.n900 VSUBS 0.010805f
C1081 B.n901 VSUBS 0.010805f
C1082 B.n902 VSUBS 0.010805f
C1083 B.n903 VSUBS 0.010805f
C1084 B.n904 VSUBS 0.010805f
C1085 B.n905 VSUBS 0.010805f
C1086 B.n906 VSUBS 0.010805f
C1087 B.n907 VSUBS 0.010805f
C1088 B.n908 VSUBS 0.010805f
C1089 B.n909 VSUBS 0.010805f
C1090 B.n910 VSUBS 0.010805f
C1091 B.n911 VSUBS 0.010805f
C1092 B.n912 VSUBS 0.010805f
C1093 B.n913 VSUBS 0.010805f
C1094 B.n914 VSUBS 0.010805f
C1095 B.n915 VSUBS 0.010805f
C1096 B.n916 VSUBS 0.010805f
C1097 B.n917 VSUBS 0.010805f
C1098 B.n918 VSUBS 0.010805f
C1099 B.n919 VSUBS 0.024466f
C1100 VTAIL.t4 VSUBS 0.189097f
C1101 VTAIL.t5 VSUBS 0.189097f
C1102 VTAIL.n0 VSUBS 1.17007f
C1103 VTAIL.n1 VSUBS 1.21312f
C1104 VTAIL.t14 VSUBS 1.59304f
C1105 VTAIL.n2 VSUBS 1.39672f
C1106 VTAIL.t16 VSUBS 0.189097f
C1107 VTAIL.t13 VSUBS 0.189097f
C1108 VTAIL.n3 VSUBS 1.17007f
C1109 VTAIL.n4 VSUBS 1.44709f
C1110 VTAIL.t18 VSUBS 0.189097f
C1111 VTAIL.t17 VSUBS 0.189097f
C1112 VTAIL.n5 VSUBS 1.17007f
C1113 VTAIL.n6 VSUBS 2.96105f
C1114 VTAIL.t6 VSUBS 0.189097f
C1115 VTAIL.t0 VSUBS 0.189097f
C1116 VTAIL.n7 VSUBS 1.17007f
C1117 VTAIL.n8 VSUBS 2.96105f
C1118 VTAIL.t7 VSUBS 0.189097f
C1119 VTAIL.t9 VSUBS 0.189097f
C1120 VTAIL.n9 VSUBS 1.17007f
C1121 VTAIL.n10 VSUBS 1.44708f
C1122 VTAIL.t8 VSUBS 1.59305f
C1123 VTAIL.n11 VSUBS 1.39671f
C1124 VTAIL.t10 VSUBS 0.189097f
C1125 VTAIL.t19 VSUBS 0.189097f
C1126 VTAIL.n12 VSUBS 1.17007f
C1127 VTAIL.n13 VSUBS 1.30397f
C1128 VTAIL.t12 VSUBS 0.189097f
C1129 VTAIL.t15 VSUBS 0.189097f
C1130 VTAIL.n14 VSUBS 1.17007f
C1131 VTAIL.n15 VSUBS 1.44708f
C1132 VTAIL.t11 VSUBS 1.59304f
C1133 VTAIL.n16 VSUBS 2.66495f
C1134 VTAIL.t3 VSUBS 1.59304f
C1135 VTAIL.n17 VSUBS 2.66495f
C1136 VTAIL.t2 VSUBS 0.189097f
C1137 VTAIL.t1 VSUBS 0.189097f
C1138 VTAIL.n18 VSUBS 1.17007f
C1139 VTAIL.n19 VSUBS 1.1491f
C1140 VDD1.t4 VSUBS 1.81262f
C1141 VDD1.t5 VSUBS 0.192554f
C1142 VDD1.t1 VSUBS 0.192554f
C1143 VDD1.n0 VSUBS 1.33087f
C1144 VDD1.n1 VSUBS 2.13292f
C1145 VDD1.t7 VSUBS 1.81262f
C1146 VDD1.t9 VSUBS 0.192554f
C1147 VDD1.t2 VSUBS 0.192554f
C1148 VDD1.n2 VSUBS 1.33086f
C1149 VDD1.n3 VSUBS 2.12127f
C1150 VDD1.t0 VSUBS 0.192554f
C1151 VDD1.t3 VSUBS 0.192554f
C1152 VDD1.n4 VSUBS 1.36877f
C1153 VDD1.n5 VSUBS 4.9699f
C1154 VDD1.t6 VSUBS 0.192554f
C1155 VDD1.t8 VSUBS 0.192554f
C1156 VDD1.n6 VSUBS 1.33086f
C1157 VDD1.n7 VSUBS 4.85292f
C1158 VP.t5 VSUBS 2.27371f
C1159 VP.n0 VSUBS 0.938917f
C1160 VP.n1 VSUBS 0.03174f
C1161 VP.n2 VSUBS 0.063779f
C1162 VP.n3 VSUBS 0.03174f
C1163 VP.n4 VSUBS 0.058859f
C1164 VP.n5 VSUBS 0.03174f
C1165 VP.t6 VSUBS 2.27371f
C1166 VP.n6 VSUBS 0.058859f
C1167 VP.n7 VSUBS 0.03174f
C1168 VP.n8 VSUBS 0.058859f
C1169 VP.n9 VSUBS 0.03174f
C1170 VP.t3 VSUBS 2.27371f
C1171 VP.n10 VSUBS 0.058859f
C1172 VP.n11 VSUBS 0.03174f
C1173 VP.n12 VSUBS 0.058859f
C1174 VP.n13 VSUBS 0.03174f
C1175 VP.t2 VSUBS 2.27371f
C1176 VP.n14 VSUBS 0.058859f
C1177 VP.n15 VSUBS 0.03174f
C1178 VP.n16 VSUBS 0.058859f
C1179 VP.n17 VSUBS 0.05122f
C1180 VP.t1 VSUBS 2.27371f
C1181 VP.t8 VSUBS 2.27371f
C1182 VP.n18 VSUBS 0.938917f
C1183 VP.n19 VSUBS 0.03174f
C1184 VP.n20 VSUBS 0.063779f
C1185 VP.n21 VSUBS 0.03174f
C1186 VP.n22 VSUBS 0.058859f
C1187 VP.n23 VSUBS 0.03174f
C1188 VP.t4 VSUBS 2.27371f
C1189 VP.n24 VSUBS 0.058859f
C1190 VP.n25 VSUBS 0.03174f
C1191 VP.n26 VSUBS 0.058859f
C1192 VP.n27 VSUBS 0.03174f
C1193 VP.t7 VSUBS 2.27371f
C1194 VP.n28 VSUBS 0.058859f
C1195 VP.n29 VSUBS 0.03174f
C1196 VP.n30 VSUBS 0.058859f
C1197 VP.t9 VSUBS 2.72422f
C1198 VP.n31 VSUBS 0.910861f
C1199 VP.t0 VSUBS 2.27371f
C1200 VP.n32 VSUBS 0.945785f
C1201 VP.n33 VSUBS 0.051886f
C1202 VP.n34 VSUBS 0.409092f
C1203 VP.n35 VSUBS 0.03174f
C1204 VP.n36 VSUBS 0.03174f
C1205 VP.n37 VSUBS 0.058859f
C1206 VP.n38 VSUBS 0.040431f
C1207 VP.n39 VSUBS 0.051847f
C1208 VP.n40 VSUBS 0.03174f
C1209 VP.n41 VSUBS 0.03174f
C1210 VP.n42 VSUBS 0.03174f
C1211 VP.n43 VSUBS 0.058859f
C1212 VP.n44 VSUBS 0.044331f
C1213 VP.n45 VSUBS 0.824517f
C1214 VP.n46 VSUBS 0.044331f
C1215 VP.n47 VSUBS 0.03174f
C1216 VP.n48 VSUBS 0.03174f
C1217 VP.n49 VSUBS 0.03174f
C1218 VP.n50 VSUBS 0.058859f
C1219 VP.n51 VSUBS 0.051847f
C1220 VP.n52 VSUBS 0.040431f
C1221 VP.n53 VSUBS 0.03174f
C1222 VP.n54 VSUBS 0.03174f
C1223 VP.n55 VSUBS 0.03174f
C1224 VP.n56 VSUBS 0.058859f
C1225 VP.n57 VSUBS 0.051886f
C1226 VP.n58 VSUBS 0.824517f
C1227 VP.n59 VSUBS 0.036776f
C1228 VP.n60 VSUBS 0.03174f
C1229 VP.n61 VSUBS 0.03174f
C1230 VP.n62 VSUBS 0.03174f
C1231 VP.n63 VSUBS 0.058859f
C1232 VP.n64 VSUBS 0.060478f
C1233 VP.n65 VSUBS 0.026881f
C1234 VP.n66 VSUBS 0.03174f
C1235 VP.n67 VSUBS 0.03174f
C1236 VP.n68 VSUBS 0.03174f
C1237 VP.n69 VSUBS 0.058859f
C1238 VP.n70 VSUBS 0.058859f
C1239 VP.n71 VSUBS 0.030383f
C1240 VP.n72 VSUBS 0.05122f
C1241 VP.n73 VSUBS 2.13418f
C1242 VP.n74 VSUBS 2.15465f
C1243 VP.n75 VSUBS 0.938917f
C1244 VP.n76 VSUBS 0.030383f
C1245 VP.n77 VSUBS 0.058859f
C1246 VP.n78 VSUBS 0.03174f
C1247 VP.n79 VSUBS 0.03174f
C1248 VP.n80 VSUBS 0.03174f
C1249 VP.n81 VSUBS 0.063779f
C1250 VP.n82 VSUBS 0.026881f
C1251 VP.n83 VSUBS 0.060478f
C1252 VP.n84 VSUBS 0.03174f
C1253 VP.n85 VSUBS 0.03174f
C1254 VP.n86 VSUBS 0.03174f
C1255 VP.n87 VSUBS 0.058859f
C1256 VP.n88 VSUBS 0.036776f
C1257 VP.n89 VSUBS 0.824517f
C1258 VP.n90 VSUBS 0.051886f
C1259 VP.n91 VSUBS 0.03174f
C1260 VP.n92 VSUBS 0.03174f
C1261 VP.n93 VSUBS 0.03174f
C1262 VP.n94 VSUBS 0.058859f
C1263 VP.n95 VSUBS 0.040431f
C1264 VP.n96 VSUBS 0.051847f
C1265 VP.n97 VSUBS 0.03174f
C1266 VP.n98 VSUBS 0.03174f
C1267 VP.n99 VSUBS 0.03174f
C1268 VP.n100 VSUBS 0.058859f
C1269 VP.n101 VSUBS 0.044331f
C1270 VP.n102 VSUBS 0.824517f
C1271 VP.n103 VSUBS 0.044331f
C1272 VP.n104 VSUBS 0.03174f
C1273 VP.n105 VSUBS 0.03174f
C1274 VP.n106 VSUBS 0.03174f
C1275 VP.n107 VSUBS 0.058859f
C1276 VP.n108 VSUBS 0.051847f
C1277 VP.n109 VSUBS 0.040431f
C1278 VP.n110 VSUBS 0.03174f
C1279 VP.n111 VSUBS 0.03174f
C1280 VP.n112 VSUBS 0.03174f
C1281 VP.n113 VSUBS 0.058859f
C1282 VP.n114 VSUBS 0.051886f
C1283 VP.n115 VSUBS 0.824517f
C1284 VP.n116 VSUBS 0.036776f
C1285 VP.n117 VSUBS 0.03174f
C1286 VP.n118 VSUBS 0.03174f
C1287 VP.n119 VSUBS 0.03174f
C1288 VP.n120 VSUBS 0.058859f
C1289 VP.n121 VSUBS 0.060478f
C1290 VP.n122 VSUBS 0.026881f
C1291 VP.n123 VSUBS 0.03174f
C1292 VP.n124 VSUBS 0.03174f
C1293 VP.n125 VSUBS 0.03174f
C1294 VP.n126 VSUBS 0.058859f
C1295 VP.n127 VSUBS 0.058859f
C1296 VP.n128 VSUBS 0.030383f
C1297 VP.n129 VSUBS 0.05122f
C1298 VP.n130 VSUBS 0.099502f
.ends

