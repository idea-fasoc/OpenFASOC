* NGSPICE file created from diff_pair_sample_0430.ext - technology: sky130A

.subckt diff_pair_sample_0430 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t9 VN.t0 VTAIL.t17 w_n2626_n3666# sky130_fd_pr__pfet_01v8 ad=2.22585 pd=13.82 as=2.22585 ps=13.82 w=13.49 l=1.05
X1 VDD2.t8 VN.t1 VTAIL.t14 w_n2626_n3666# sky130_fd_pr__pfet_01v8 ad=2.22585 pd=13.82 as=2.22585 ps=13.82 w=13.49 l=1.05
X2 B.t11 B.t9 B.t10 w_n2626_n3666# sky130_fd_pr__pfet_01v8 ad=5.2611 pd=27.76 as=0 ps=0 w=13.49 l=1.05
X3 VDD1.t9 VP.t0 VTAIL.t9 w_n2626_n3666# sky130_fd_pr__pfet_01v8 ad=2.22585 pd=13.82 as=5.2611 ps=27.76 w=13.49 l=1.05
X4 VTAIL.t1 VP.t1 VDD1.t8 w_n2626_n3666# sky130_fd_pr__pfet_01v8 ad=2.22585 pd=13.82 as=2.22585 ps=13.82 w=13.49 l=1.05
X5 B.t8 B.t6 B.t7 w_n2626_n3666# sky130_fd_pr__pfet_01v8 ad=5.2611 pd=27.76 as=0 ps=0 w=13.49 l=1.05
X6 VDD1.t7 VP.t2 VTAIL.t2 w_n2626_n3666# sky130_fd_pr__pfet_01v8 ad=2.22585 pd=13.82 as=2.22585 ps=13.82 w=13.49 l=1.05
X7 B.t5 B.t3 B.t4 w_n2626_n3666# sky130_fd_pr__pfet_01v8 ad=5.2611 pd=27.76 as=0 ps=0 w=13.49 l=1.05
X8 VTAIL.t10 VN.t2 VDD2.t7 w_n2626_n3666# sky130_fd_pr__pfet_01v8 ad=2.22585 pd=13.82 as=2.22585 ps=13.82 w=13.49 l=1.05
X9 VTAIL.t19 VN.t3 VDD2.t6 w_n2626_n3666# sky130_fd_pr__pfet_01v8 ad=2.22585 pd=13.82 as=2.22585 ps=13.82 w=13.49 l=1.05
X10 B.t2 B.t0 B.t1 w_n2626_n3666# sky130_fd_pr__pfet_01v8 ad=5.2611 pd=27.76 as=0 ps=0 w=13.49 l=1.05
X11 VTAIL.t5 VP.t3 VDD1.t6 w_n2626_n3666# sky130_fd_pr__pfet_01v8 ad=2.22585 pd=13.82 as=2.22585 ps=13.82 w=13.49 l=1.05
X12 VDD2.t5 VN.t4 VTAIL.t11 w_n2626_n3666# sky130_fd_pr__pfet_01v8 ad=2.22585 pd=13.82 as=5.2611 ps=27.76 w=13.49 l=1.05
X13 VDD1.t5 VP.t4 VTAIL.t0 w_n2626_n3666# sky130_fd_pr__pfet_01v8 ad=5.2611 pd=27.76 as=2.22585 ps=13.82 w=13.49 l=1.05
X14 VTAIL.t18 VN.t5 VDD2.t4 w_n2626_n3666# sky130_fd_pr__pfet_01v8 ad=2.22585 pd=13.82 as=2.22585 ps=13.82 w=13.49 l=1.05
X15 VDD1.t4 VP.t5 VTAIL.t4 w_n2626_n3666# sky130_fd_pr__pfet_01v8 ad=5.2611 pd=27.76 as=2.22585 ps=13.82 w=13.49 l=1.05
X16 VDD2.t3 VN.t6 VTAIL.t13 w_n2626_n3666# sky130_fd_pr__pfet_01v8 ad=2.22585 pd=13.82 as=5.2611 ps=27.76 w=13.49 l=1.05
X17 VTAIL.t7 VP.t6 VDD1.t3 w_n2626_n3666# sky130_fd_pr__pfet_01v8 ad=2.22585 pd=13.82 as=2.22585 ps=13.82 w=13.49 l=1.05
X18 VDD1.t2 VP.t7 VTAIL.t6 w_n2626_n3666# sky130_fd_pr__pfet_01v8 ad=2.22585 pd=13.82 as=5.2611 ps=27.76 w=13.49 l=1.05
X19 VDD1.t1 VP.t8 VTAIL.t8 w_n2626_n3666# sky130_fd_pr__pfet_01v8 ad=2.22585 pd=13.82 as=2.22585 ps=13.82 w=13.49 l=1.05
X20 VTAIL.t3 VP.t9 VDD1.t0 w_n2626_n3666# sky130_fd_pr__pfet_01v8 ad=2.22585 pd=13.82 as=2.22585 ps=13.82 w=13.49 l=1.05
X21 VTAIL.t16 VN.t7 VDD2.t2 w_n2626_n3666# sky130_fd_pr__pfet_01v8 ad=2.22585 pd=13.82 as=2.22585 ps=13.82 w=13.49 l=1.05
X22 VDD2.t1 VN.t8 VTAIL.t15 w_n2626_n3666# sky130_fd_pr__pfet_01v8 ad=5.2611 pd=27.76 as=2.22585 ps=13.82 w=13.49 l=1.05
X23 VDD2.t0 VN.t9 VTAIL.t12 w_n2626_n3666# sky130_fd_pr__pfet_01v8 ad=5.2611 pd=27.76 as=2.22585 ps=13.82 w=13.49 l=1.05
R0 VN.n5 VN.t9 362.413
R1 VN.n25 VN.t4 362.413
R2 VN.n18 VN.t6 347.271
R3 VN.n38 VN.t8 347.271
R4 VN.n4 VN.t5 309.628
R5 VN.n10 VN.t1 309.628
R6 VN.n16 VN.t2 309.628
R7 VN.n24 VN.t3 309.628
R8 VN.n30 VN.t0 309.628
R9 VN.n36 VN.t7 309.628
R10 VN.n37 VN.n20 161.3
R11 VN.n35 VN.n34 161.3
R12 VN.n33 VN.n21 161.3
R13 VN.n32 VN.n31 161.3
R14 VN.n29 VN.n22 161.3
R15 VN.n28 VN.n27 161.3
R16 VN.n26 VN.n23 161.3
R17 VN.n17 VN.n0 161.3
R18 VN.n15 VN.n14 161.3
R19 VN.n13 VN.n1 161.3
R20 VN.n12 VN.n11 161.3
R21 VN.n9 VN.n2 161.3
R22 VN.n8 VN.n7 161.3
R23 VN.n6 VN.n3 161.3
R24 VN.n39 VN.n38 80.6037
R25 VN.n19 VN.n18 80.6037
R26 VN.n18 VN.n17 55.7853
R27 VN.n38 VN.n37 55.7853
R28 VN.n5 VN.n4 48.3043
R29 VN.n25 VN.n24 48.3043
R30 VN VN.n39 46.34
R31 VN.n9 VN.n8 46.321
R32 VN.n11 VN.n1 46.321
R33 VN.n29 VN.n28 46.321
R34 VN.n31 VN.n21 46.321
R35 VN.n26 VN.n25 43.9769
R36 VN.n6 VN.n5 43.9769
R37 VN.n8 VN.n3 34.6658
R38 VN.n15 VN.n1 34.6658
R39 VN.n28 VN.n23 34.6658
R40 VN.n35 VN.n21 34.6658
R41 VN.n17 VN.n16 18.1061
R42 VN.n37 VN.n36 18.1061
R43 VN.n10 VN.n9 12.234
R44 VN.n11 VN.n10 12.234
R45 VN.n31 VN.n30 12.234
R46 VN.n30 VN.n29 12.234
R47 VN.n4 VN.n3 6.36192
R48 VN.n16 VN.n15 6.36192
R49 VN.n24 VN.n23 6.36192
R50 VN.n36 VN.n35 6.36192
R51 VN.n39 VN.n20 0.285035
R52 VN.n19 VN.n0 0.285035
R53 VN.n34 VN.n20 0.189894
R54 VN.n34 VN.n33 0.189894
R55 VN.n33 VN.n32 0.189894
R56 VN.n32 VN.n22 0.189894
R57 VN.n27 VN.n22 0.189894
R58 VN.n27 VN.n26 0.189894
R59 VN.n7 VN.n6 0.189894
R60 VN.n7 VN.n2 0.189894
R61 VN.n12 VN.n2 0.189894
R62 VN.n13 VN.n12 0.189894
R63 VN.n14 VN.n13 0.189894
R64 VN.n14 VN.n0 0.189894
R65 VN VN.n19 0.146778
R66 VTAIL.n304 VTAIL.n236 756.745
R67 VTAIL.n70 VTAIL.n2 756.745
R68 VTAIL.n230 VTAIL.n162 756.745
R69 VTAIL.n152 VTAIL.n84 756.745
R70 VTAIL.n261 VTAIL.n260 585
R71 VTAIL.n263 VTAIL.n262 585
R72 VTAIL.n256 VTAIL.n255 585
R73 VTAIL.n269 VTAIL.n268 585
R74 VTAIL.n271 VTAIL.n270 585
R75 VTAIL.n252 VTAIL.n251 585
R76 VTAIL.n278 VTAIL.n277 585
R77 VTAIL.n279 VTAIL.n250 585
R78 VTAIL.n281 VTAIL.n280 585
R79 VTAIL.n248 VTAIL.n247 585
R80 VTAIL.n287 VTAIL.n286 585
R81 VTAIL.n289 VTAIL.n288 585
R82 VTAIL.n244 VTAIL.n243 585
R83 VTAIL.n295 VTAIL.n294 585
R84 VTAIL.n297 VTAIL.n296 585
R85 VTAIL.n240 VTAIL.n239 585
R86 VTAIL.n303 VTAIL.n302 585
R87 VTAIL.n305 VTAIL.n304 585
R88 VTAIL.n27 VTAIL.n26 585
R89 VTAIL.n29 VTAIL.n28 585
R90 VTAIL.n22 VTAIL.n21 585
R91 VTAIL.n35 VTAIL.n34 585
R92 VTAIL.n37 VTAIL.n36 585
R93 VTAIL.n18 VTAIL.n17 585
R94 VTAIL.n44 VTAIL.n43 585
R95 VTAIL.n45 VTAIL.n16 585
R96 VTAIL.n47 VTAIL.n46 585
R97 VTAIL.n14 VTAIL.n13 585
R98 VTAIL.n53 VTAIL.n52 585
R99 VTAIL.n55 VTAIL.n54 585
R100 VTAIL.n10 VTAIL.n9 585
R101 VTAIL.n61 VTAIL.n60 585
R102 VTAIL.n63 VTAIL.n62 585
R103 VTAIL.n6 VTAIL.n5 585
R104 VTAIL.n69 VTAIL.n68 585
R105 VTAIL.n71 VTAIL.n70 585
R106 VTAIL.n231 VTAIL.n230 585
R107 VTAIL.n229 VTAIL.n228 585
R108 VTAIL.n166 VTAIL.n165 585
R109 VTAIL.n223 VTAIL.n222 585
R110 VTAIL.n221 VTAIL.n220 585
R111 VTAIL.n170 VTAIL.n169 585
R112 VTAIL.n215 VTAIL.n214 585
R113 VTAIL.n213 VTAIL.n212 585
R114 VTAIL.n174 VTAIL.n173 585
R115 VTAIL.n178 VTAIL.n176 585
R116 VTAIL.n207 VTAIL.n206 585
R117 VTAIL.n205 VTAIL.n204 585
R118 VTAIL.n180 VTAIL.n179 585
R119 VTAIL.n199 VTAIL.n198 585
R120 VTAIL.n197 VTAIL.n196 585
R121 VTAIL.n184 VTAIL.n183 585
R122 VTAIL.n191 VTAIL.n190 585
R123 VTAIL.n189 VTAIL.n188 585
R124 VTAIL.n153 VTAIL.n152 585
R125 VTAIL.n151 VTAIL.n150 585
R126 VTAIL.n88 VTAIL.n87 585
R127 VTAIL.n145 VTAIL.n144 585
R128 VTAIL.n143 VTAIL.n142 585
R129 VTAIL.n92 VTAIL.n91 585
R130 VTAIL.n137 VTAIL.n136 585
R131 VTAIL.n135 VTAIL.n134 585
R132 VTAIL.n96 VTAIL.n95 585
R133 VTAIL.n100 VTAIL.n98 585
R134 VTAIL.n129 VTAIL.n128 585
R135 VTAIL.n127 VTAIL.n126 585
R136 VTAIL.n102 VTAIL.n101 585
R137 VTAIL.n121 VTAIL.n120 585
R138 VTAIL.n119 VTAIL.n118 585
R139 VTAIL.n106 VTAIL.n105 585
R140 VTAIL.n113 VTAIL.n112 585
R141 VTAIL.n111 VTAIL.n110 585
R142 VTAIL.n259 VTAIL.t13 329.036
R143 VTAIL.n25 VTAIL.t9 329.036
R144 VTAIL.n187 VTAIL.t6 329.036
R145 VTAIL.n109 VTAIL.t11 329.036
R146 VTAIL.n262 VTAIL.n261 171.744
R147 VTAIL.n262 VTAIL.n255 171.744
R148 VTAIL.n269 VTAIL.n255 171.744
R149 VTAIL.n270 VTAIL.n269 171.744
R150 VTAIL.n270 VTAIL.n251 171.744
R151 VTAIL.n278 VTAIL.n251 171.744
R152 VTAIL.n279 VTAIL.n278 171.744
R153 VTAIL.n280 VTAIL.n279 171.744
R154 VTAIL.n280 VTAIL.n247 171.744
R155 VTAIL.n287 VTAIL.n247 171.744
R156 VTAIL.n288 VTAIL.n287 171.744
R157 VTAIL.n288 VTAIL.n243 171.744
R158 VTAIL.n295 VTAIL.n243 171.744
R159 VTAIL.n296 VTAIL.n295 171.744
R160 VTAIL.n296 VTAIL.n239 171.744
R161 VTAIL.n303 VTAIL.n239 171.744
R162 VTAIL.n304 VTAIL.n303 171.744
R163 VTAIL.n28 VTAIL.n27 171.744
R164 VTAIL.n28 VTAIL.n21 171.744
R165 VTAIL.n35 VTAIL.n21 171.744
R166 VTAIL.n36 VTAIL.n35 171.744
R167 VTAIL.n36 VTAIL.n17 171.744
R168 VTAIL.n44 VTAIL.n17 171.744
R169 VTAIL.n45 VTAIL.n44 171.744
R170 VTAIL.n46 VTAIL.n45 171.744
R171 VTAIL.n46 VTAIL.n13 171.744
R172 VTAIL.n53 VTAIL.n13 171.744
R173 VTAIL.n54 VTAIL.n53 171.744
R174 VTAIL.n54 VTAIL.n9 171.744
R175 VTAIL.n61 VTAIL.n9 171.744
R176 VTAIL.n62 VTAIL.n61 171.744
R177 VTAIL.n62 VTAIL.n5 171.744
R178 VTAIL.n69 VTAIL.n5 171.744
R179 VTAIL.n70 VTAIL.n69 171.744
R180 VTAIL.n230 VTAIL.n229 171.744
R181 VTAIL.n229 VTAIL.n165 171.744
R182 VTAIL.n222 VTAIL.n165 171.744
R183 VTAIL.n222 VTAIL.n221 171.744
R184 VTAIL.n221 VTAIL.n169 171.744
R185 VTAIL.n214 VTAIL.n169 171.744
R186 VTAIL.n214 VTAIL.n213 171.744
R187 VTAIL.n213 VTAIL.n173 171.744
R188 VTAIL.n178 VTAIL.n173 171.744
R189 VTAIL.n206 VTAIL.n178 171.744
R190 VTAIL.n206 VTAIL.n205 171.744
R191 VTAIL.n205 VTAIL.n179 171.744
R192 VTAIL.n198 VTAIL.n179 171.744
R193 VTAIL.n198 VTAIL.n197 171.744
R194 VTAIL.n197 VTAIL.n183 171.744
R195 VTAIL.n190 VTAIL.n183 171.744
R196 VTAIL.n190 VTAIL.n189 171.744
R197 VTAIL.n152 VTAIL.n151 171.744
R198 VTAIL.n151 VTAIL.n87 171.744
R199 VTAIL.n144 VTAIL.n87 171.744
R200 VTAIL.n144 VTAIL.n143 171.744
R201 VTAIL.n143 VTAIL.n91 171.744
R202 VTAIL.n136 VTAIL.n91 171.744
R203 VTAIL.n136 VTAIL.n135 171.744
R204 VTAIL.n135 VTAIL.n95 171.744
R205 VTAIL.n100 VTAIL.n95 171.744
R206 VTAIL.n128 VTAIL.n100 171.744
R207 VTAIL.n128 VTAIL.n127 171.744
R208 VTAIL.n127 VTAIL.n101 171.744
R209 VTAIL.n120 VTAIL.n101 171.744
R210 VTAIL.n120 VTAIL.n119 171.744
R211 VTAIL.n119 VTAIL.n105 171.744
R212 VTAIL.n112 VTAIL.n105 171.744
R213 VTAIL.n112 VTAIL.n111 171.744
R214 VTAIL.n261 VTAIL.t13 85.8723
R215 VTAIL.n27 VTAIL.t9 85.8723
R216 VTAIL.n189 VTAIL.t6 85.8723
R217 VTAIL.n111 VTAIL.t11 85.8723
R218 VTAIL.n161 VTAIL.n160 54.2445
R219 VTAIL.n159 VTAIL.n158 54.2445
R220 VTAIL.n83 VTAIL.n82 54.2445
R221 VTAIL.n81 VTAIL.n80 54.2445
R222 VTAIL.n311 VTAIL.n310 54.2443
R223 VTAIL.n1 VTAIL.n0 54.2443
R224 VTAIL.n77 VTAIL.n76 54.2443
R225 VTAIL.n79 VTAIL.n78 54.2443
R226 VTAIL.n309 VTAIL.n308 30.8278
R227 VTAIL.n75 VTAIL.n74 30.8278
R228 VTAIL.n235 VTAIL.n234 30.8278
R229 VTAIL.n157 VTAIL.n156 30.8278
R230 VTAIL.n81 VTAIL.n79 26.3755
R231 VTAIL.n309 VTAIL.n235 25.1858
R232 VTAIL.n281 VTAIL.n248 13.1884
R233 VTAIL.n47 VTAIL.n14 13.1884
R234 VTAIL.n176 VTAIL.n174 13.1884
R235 VTAIL.n98 VTAIL.n96 13.1884
R236 VTAIL.n282 VTAIL.n250 12.8005
R237 VTAIL.n286 VTAIL.n285 12.8005
R238 VTAIL.n48 VTAIL.n16 12.8005
R239 VTAIL.n52 VTAIL.n51 12.8005
R240 VTAIL.n212 VTAIL.n211 12.8005
R241 VTAIL.n208 VTAIL.n207 12.8005
R242 VTAIL.n134 VTAIL.n133 12.8005
R243 VTAIL.n130 VTAIL.n129 12.8005
R244 VTAIL.n277 VTAIL.n276 12.0247
R245 VTAIL.n289 VTAIL.n246 12.0247
R246 VTAIL.n43 VTAIL.n42 12.0247
R247 VTAIL.n55 VTAIL.n12 12.0247
R248 VTAIL.n215 VTAIL.n172 12.0247
R249 VTAIL.n204 VTAIL.n177 12.0247
R250 VTAIL.n137 VTAIL.n94 12.0247
R251 VTAIL.n126 VTAIL.n99 12.0247
R252 VTAIL.n275 VTAIL.n252 11.249
R253 VTAIL.n290 VTAIL.n244 11.249
R254 VTAIL.n41 VTAIL.n18 11.249
R255 VTAIL.n56 VTAIL.n10 11.249
R256 VTAIL.n216 VTAIL.n170 11.249
R257 VTAIL.n203 VTAIL.n180 11.249
R258 VTAIL.n138 VTAIL.n92 11.249
R259 VTAIL.n125 VTAIL.n102 11.249
R260 VTAIL.n260 VTAIL.n259 10.7239
R261 VTAIL.n26 VTAIL.n25 10.7239
R262 VTAIL.n188 VTAIL.n187 10.7239
R263 VTAIL.n110 VTAIL.n109 10.7239
R264 VTAIL.n272 VTAIL.n271 10.4732
R265 VTAIL.n294 VTAIL.n293 10.4732
R266 VTAIL.n38 VTAIL.n37 10.4732
R267 VTAIL.n60 VTAIL.n59 10.4732
R268 VTAIL.n220 VTAIL.n219 10.4732
R269 VTAIL.n200 VTAIL.n199 10.4732
R270 VTAIL.n142 VTAIL.n141 10.4732
R271 VTAIL.n122 VTAIL.n121 10.4732
R272 VTAIL.n268 VTAIL.n254 9.69747
R273 VTAIL.n297 VTAIL.n242 9.69747
R274 VTAIL.n34 VTAIL.n20 9.69747
R275 VTAIL.n63 VTAIL.n8 9.69747
R276 VTAIL.n223 VTAIL.n168 9.69747
R277 VTAIL.n196 VTAIL.n182 9.69747
R278 VTAIL.n145 VTAIL.n90 9.69747
R279 VTAIL.n118 VTAIL.n104 9.69747
R280 VTAIL.n308 VTAIL.n307 9.45567
R281 VTAIL.n74 VTAIL.n73 9.45567
R282 VTAIL.n234 VTAIL.n233 9.45567
R283 VTAIL.n156 VTAIL.n155 9.45567
R284 VTAIL.n307 VTAIL.n306 9.3005
R285 VTAIL.n301 VTAIL.n300 9.3005
R286 VTAIL.n299 VTAIL.n298 9.3005
R287 VTAIL.n242 VTAIL.n241 9.3005
R288 VTAIL.n293 VTAIL.n292 9.3005
R289 VTAIL.n291 VTAIL.n290 9.3005
R290 VTAIL.n246 VTAIL.n245 9.3005
R291 VTAIL.n285 VTAIL.n284 9.3005
R292 VTAIL.n258 VTAIL.n257 9.3005
R293 VTAIL.n265 VTAIL.n264 9.3005
R294 VTAIL.n267 VTAIL.n266 9.3005
R295 VTAIL.n254 VTAIL.n253 9.3005
R296 VTAIL.n273 VTAIL.n272 9.3005
R297 VTAIL.n275 VTAIL.n274 9.3005
R298 VTAIL.n276 VTAIL.n249 9.3005
R299 VTAIL.n283 VTAIL.n282 9.3005
R300 VTAIL.n238 VTAIL.n237 9.3005
R301 VTAIL.n73 VTAIL.n72 9.3005
R302 VTAIL.n67 VTAIL.n66 9.3005
R303 VTAIL.n65 VTAIL.n64 9.3005
R304 VTAIL.n8 VTAIL.n7 9.3005
R305 VTAIL.n59 VTAIL.n58 9.3005
R306 VTAIL.n57 VTAIL.n56 9.3005
R307 VTAIL.n12 VTAIL.n11 9.3005
R308 VTAIL.n51 VTAIL.n50 9.3005
R309 VTAIL.n24 VTAIL.n23 9.3005
R310 VTAIL.n31 VTAIL.n30 9.3005
R311 VTAIL.n33 VTAIL.n32 9.3005
R312 VTAIL.n20 VTAIL.n19 9.3005
R313 VTAIL.n39 VTAIL.n38 9.3005
R314 VTAIL.n41 VTAIL.n40 9.3005
R315 VTAIL.n42 VTAIL.n15 9.3005
R316 VTAIL.n49 VTAIL.n48 9.3005
R317 VTAIL.n4 VTAIL.n3 9.3005
R318 VTAIL.n186 VTAIL.n185 9.3005
R319 VTAIL.n193 VTAIL.n192 9.3005
R320 VTAIL.n195 VTAIL.n194 9.3005
R321 VTAIL.n182 VTAIL.n181 9.3005
R322 VTAIL.n201 VTAIL.n200 9.3005
R323 VTAIL.n203 VTAIL.n202 9.3005
R324 VTAIL.n177 VTAIL.n175 9.3005
R325 VTAIL.n209 VTAIL.n208 9.3005
R326 VTAIL.n233 VTAIL.n232 9.3005
R327 VTAIL.n164 VTAIL.n163 9.3005
R328 VTAIL.n227 VTAIL.n226 9.3005
R329 VTAIL.n225 VTAIL.n224 9.3005
R330 VTAIL.n168 VTAIL.n167 9.3005
R331 VTAIL.n219 VTAIL.n218 9.3005
R332 VTAIL.n217 VTAIL.n216 9.3005
R333 VTAIL.n172 VTAIL.n171 9.3005
R334 VTAIL.n211 VTAIL.n210 9.3005
R335 VTAIL.n108 VTAIL.n107 9.3005
R336 VTAIL.n115 VTAIL.n114 9.3005
R337 VTAIL.n117 VTAIL.n116 9.3005
R338 VTAIL.n104 VTAIL.n103 9.3005
R339 VTAIL.n123 VTAIL.n122 9.3005
R340 VTAIL.n125 VTAIL.n124 9.3005
R341 VTAIL.n99 VTAIL.n97 9.3005
R342 VTAIL.n131 VTAIL.n130 9.3005
R343 VTAIL.n155 VTAIL.n154 9.3005
R344 VTAIL.n86 VTAIL.n85 9.3005
R345 VTAIL.n149 VTAIL.n148 9.3005
R346 VTAIL.n147 VTAIL.n146 9.3005
R347 VTAIL.n90 VTAIL.n89 9.3005
R348 VTAIL.n141 VTAIL.n140 9.3005
R349 VTAIL.n139 VTAIL.n138 9.3005
R350 VTAIL.n94 VTAIL.n93 9.3005
R351 VTAIL.n133 VTAIL.n132 9.3005
R352 VTAIL.n267 VTAIL.n256 8.92171
R353 VTAIL.n298 VTAIL.n240 8.92171
R354 VTAIL.n33 VTAIL.n22 8.92171
R355 VTAIL.n64 VTAIL.n6 8.92171
R356 VTAIL.n224 VTAIL.n166 8.92171
R357 VTAIL.n195 VTAIL.n184 8.92171
R358 VTAIL.n146 VTAIL.n88 8.92171
R359 VTAIL.n117 VTAIL.n106 8.92171
R360 VTAIL.n264 VTAIL.n263 8.14595
R361 VTAIL.n302 VTAIL.n301 8.14595
R362 VTAIL.n30 VTAIL.n29 8.14595
R363 VTAIL.n68 VTAIL.n67 8.14595
R364 VTAIL.n228 VTAIL.n227 8.14595
R365 VTAIL.n192 VTAIL.n191 8.14595
R366 VTAIL.n150 VTAIL.n149 8.14595
R367 VTAIL.n114 VTAIL.n113 8.14595
R368 VTAIL.n260 VTAIL.n258 7.3702
R369 VTAIL.n305 VTAIL.n238 7.3702
R370 VTAIL.n308 VTAIL.n236 7.3702
R371 VTAIL.n26 VTAIL.n24 7.3702
R372 VTAIL.n71 VTAIL.n4 7.3702
R373 VTAIL.n74 VTAIL.n2 7.3702
R374 VTAIL.n234 VTAIL.n162 7.3702
R375 VTAIL.n231 VTAIL.n164 7.3702
R376 VTAIL.n188 VTAIL.n186 7.3702
R377 VTAIL.n156 VTAIL.n84 7.3702
R378 VTAIL.n153 VTAIL.n86 7.3702
R379 VTAIL.n110 VTAIL.n108 7.3702
R380 VTAIL.n306 VTAIL.n305 6.59444
R381 VTAIL.n306 VTAIL.n236 6.59444
R382 VTAIL.n72 VTAIL.n71 6.59444
R383 VTAIL.n72 VTAIL.n2 6.59444
R384 VTAIL.n232 VTAIL.n162 6.59444
R385 VTAIL.n232 VTAIL.n231 6.59444
R386 VTAIL.n154 VTAIL.n84 6.59444
R387 VTAIL.n154 VTAIL.n153 6.59444
R388 VTAIL.n263 VTAIL.n258 5.81868
R389 VTAIL.n302 VTAIL.n238 5.81868
R390 VTAIL.n29 VTAIL.n24 5.81868
R391 VTAIL.n68 VTAIL.n4 5.81868
R392 VTAIL.n228 VTAIL.n164 5.81868
R393 VTAIL.n191 VTAIL.n186 5.81868
R394 VTAIL.n150 VTAIL.n86 5.81868
R395 VTAIL.n113 VTAIL.n108 5.81868
R396 VTAIL.n264 VTAIL.n256 5.04292
R397 VTAIL.n301 VTAIL.n240 5.04292
R398 VTAIL.n30 VTAIL.n22 5.04292
R399 VTAIL.n67 VTAIL.n6 5.04292
R400 VTAIL.n227 VTAIL.n166 5.04292
R401 VTAIL.n192 VTAIL.n184 5.04292
R402 VTAIL.n149 VTAIL.n88 5.04292
R403 VTAIL.n114 VTAIL.n106 5.04292
R404 VTAIL.n268 VTAIL.n267 4.26717
R405 VTAIL.n298 VTAIL.n297 4.26717
R406 VTAIL.n34 VTAIL.n33 4.26717
R407 VTAIL.n64 VTAIL.n63 4.26717
R408 VTAIL.n224 VTAIL.n223 4.26717
R409 VTAIL.n196 VTAIL.n195 4.26717
R410 VTAIL.n146 VTAIL.n145 4.26717
R411 VTAIL.n118 VTAIL.n117 4.26717
R412 VTAIL.n271 VTAIL.n254 3.49141
R413 VTAIL.n294 VTAIL.n242 3.49141
R414 VTAIL.n37 VTAIL.n20 3.49141
R415 VTAIL.n60 VTAIL.n8 3.49141
R416 VTAIL.n220 VTAIL.n168 3.49141
R417 VTAIL.n199 VTAIL.n182 3.49141
R418 VTAIL.n142 VTAIL.n90 3.49141
R419 VTAIL.n121 VTAIL.n104 3.49141
R420 VTAIL.n272 VTAIL.n252 2.71565
R421 VTAIL.n293 VTAIL.n244 2.71565
R422 VTAIL.n38 VTAIL.n18 2.71565
R423 VTAIL.n59 VTAIL.n10 2.71565
R424 VTAIL.n219 VTAIL.n170 2.71565
R425 VTAIL.n200 VTAIL.n180 2.71565
R426 VTAIL.n141 VTAIL.n92 2.71565
R427 VTAIL.n122 VTAIL.n102 2.71565
R428 VTAIL.n259 VTAIL.n257 2.41282
R429 VTAIL.n25 VTAIL.n23 2.41282
R430 VTAIL.n187 VTAIL.n185 2.41282
R431 VTAIL.n109 VTAIL.n107 2.41282
R432 VTAIL.n310 VTAIL.t14 2.41006
R433 VTAIL.n310 VTAIL.t10 2.41006
R434 VTAIL.n0 VTAIL.t12 2.41006
R435 VTAIL.n0 VTAIL.t18 2.41006
R436 VTAIL.n76 VTAIL.t8 2.41006
R437 VTAIL.n76 VTAIL.t7 2.41006
R438 VTAIL.n78 VTAIL.t4 2.41006
R439 VTAIL.n78 VTAIL.t1 2.41006
R440 VTAIL.n160 VTAIL.t2 2.41006
R441 VTAIL.n160 VTAIL.t3 2.41006
R442 VTAIL.n158 VTAIL.t0 2.41006
R443 VTAIL.n158 VTAIL.t5 2.41006
R444 VTAIL.n82 VTAIL.t17 2.41006
R445 VTAIL.n82 VTAIL.t19 2.41006
R446 VTAIL.n80 VTAIL.t15 2.41006
R447 VTAIL.n80 VTAIL.t16 2.41006
R448 VTAIL.n277 VTAIL.n275 1.93989
R449 VTAIL.n290 VTAIL.n289 1.93989
R450 VTAIL.n43 VTAIL.n41 1.93989
R451 VTAIL.n56 VTAIL.n55 1.93989
R452 VTAIL.n216 VTAIL.n215 1.93989
R453 VTAIL.n204 VTAIL.n203 1.93989
R454 VTAIL.n138 VTAIL.n137 1.93989
R455 VTAIL.n126 VTAIL.n125 1.93989
R456 VTAIL.n83 VTAIL.n81 1.19016
R457 VTAIL.n157 VTAIL.n83 1.19016
R458 VTAIL.n161 VTAIL.n159 1.19016
R459 VTAIL.n235 VTAIL.n161 1.19016
R460 VTAIL.n79 VTAIL.n77 1.19016
R461 VTAIL.n77 VTAIL.n75 1.19016
R462 VTAIL.n311 VTAIL.n309 1.19016
R463 VTAIL.n276 VTAIL.n250 1.16414
R464 VTAIL.n286 VTAIL.n246 1.16414
R465 VTAIL.n42 VTAIL.n16 1.16414
R466 VTAIL.n52 VTAIL.n12 1.16414
R467 VTAIL.n212 VTAIL.n172 1.16414
R468 VTAIL.n207 VTAIL.n177 1.16414
R469 VTAIL.n134 VTAIL.n94 1.16414
R470 VTAIL.n129 VTAIL.n99 1.16414
R471 VTAIL.n159 VTAIL.n157 1.06516
R472 VTAIL.n75 VTAIL.n1 1.06516
R473 VTAIL VTAIL.n1 0.950931
R474 VTAIL.n282 VTAIL.n281 0.388379
R475 VTAIL.n285 VTAIL.n248 0.388379
R476 VTAIL.n48 VTAIL.n47 0.388379
R477 VTAIL.n51 VTAIL.n14 0.388379
R478 VTAIL.n211 VTAIL.n174 0.388379
R479 VTAIL.n208 VTAIL.n176 0.388379
R480 VTAIL.n133 VTAIL.n96 0.388379
R481 VTAIL.n130 VTAIL.n98 0.388379
R482 VTAIL VTAIL.n311 0.239724
R483 VTAIL.n265 VTAIL.n257 0.155672
R484 VTAIL.n266 VTAIL.n265 0.155672
R485 VTAIL.n266 VTAIL.n253 0.155672
R486 VTAIL.n273 VTAIL.n253 0.155672
R487 VTAIL.n274 VTAIL.n273 0.155672
R488 VTAIL.n274 VTAIL.n249 0.155672
R489 VTAIL.n283 VTAIL.n249 0.155672
R490 VTAIL.n284 VTAIL.n283 0.155672
R491 VTAIL.n284 VTAIL.n245 0.155672
R492 VTAIL.n291 VTAIL.n245 0.155672
R493 VTAIL.n292 VTAIL.n291 0.155672
R494 VTAIL.n292 VTAIL.n241 0.155672
R495 VTAIL.n299 VTAIL.n241 0.155672
R496 VTAIL.n300 VTAIL.n299 0.155672
R497 VTAIL.n300 VTAIL.n237 0.155672
R498 VTAIL.n307 VTAIL.n237 0.155672
R499 VTAIL.n31 VTAIL.n23 0.155672
R500 VTAIL.n32 VTAIL.n31 0.155672
R501 VTAIL.n32 VTAIL.n19 0.155672
R502 VTAIL.n39 VTAIL.n19 0.155672
R503 VTAIL.n40 VTAIL.n39 0.155672
R504 VTAIL.n40 VTAIL.n15 0.155672
R505 VTAIL.n49 VTAIL.n15 0.155672
R506 VTAIL.n50 VTAIL.n49 0.155672
R507 VTAIL.n50 VTAIL.n11 0.155672
R508 VTAIL.n57 VTAIL.n11 0.155672
R509 VTAIL.n58 VTAIL.n57 0.155672
R510 VTAIL.n58 VTAIL.n7 0.155672
R511 VTAIL.n65 VTAIL.n7 0.155672
R512 VTAIL.n66 VTAIL.n65 0.155672
R513 VTAIL.n66 VTAIL.n3 0.155672
R514 VTAIL.n73 VTAIL.n3 0.155672
R515 VTAIL.n233 VTAIL.n163 0.155672
R516 VTAIL.n226 VTAIL.n163 0.155672
R517 VTAIL.n226 VTAIL.n225 0.155672
R518 VTAIL.n225 VTAIL.n167 0.155672
R519 VTAIL.n218 VTAIL.n167 0.155672
R520 VTAIL.n218 VTAIL.n217 0.155672
R521 VTAIL.n217 VTAIL.n171 0.155672
R522 VTAIL.n210 VTAIL.n171 0.155672
R523 VTAIL.n210 VTAIL.n209 0.155672
R524 VTAIL.n209 VTAIL.n175 0.155672
R525 VTAIL.n202 VTAIL.n175 0.155672
R526 VTAIL.n202 VTAIL.n201 0.155672
R527 VTAIL.n201 VTAIL.n181 0.155672
R528 VTAIL.n194 VTAIL.n181 0.155672
R529 VTAIL.n194 VTAIL.n193 0.155672
R530 VTAIL.n193 VTAIL.n185 0.155672
R531 VTAIL.n155 VTAIL.n85 0.155672
R532 VTAIL.n148 VTAIL.n85 0.155672
R533 VTAIL.n148 VTAIL.n147 0.155672
R534 VTAIL.n147 VTAIL.n89 0.155672
R535 VTAIL.n140 VTAIL.n89 0.155672
R536 VTAIL.n140 VTAIL.n139 0.155672
R537 VTAIL.n139 VTAIL.n93 0.155672
R538 VTAIL.n132 VTAIL.n93 0.155672
R539 VTAIL.n132 VTAIL.n131 0.155672
R540 VTAIL.n131 VTAIL.n97 0.155672
R541 VTAIL.n124 VTAIL.n97 0.155672
R542 VTAIL.n124 VTAIL.n123 0.155672
R543 VTAIL.n123 VTAIL.n103 0.155672
R544 VTAIL.n116 VTAIL.n103 0.155672
R545 VTAIL.n116 VTAIL.n115 0.155672
R546 VTAIL.n115 VTAIL.n107 0.155672
R547 VDD2.n145 VDD2.n77 756.745
R548 VDD2.n68 VDD2.n0 756.745
R549 VDD2.n146 VDD2.n145 585
R550 VDD2.n144 VDD2.n143 585
R551 VDD2.n81 VDD2.n80 585
R552 VDD2.n138 VDD2.n137 585
R553 VDD2.n136 VDD2.n135 585
R554 VDD2.n85 VDD2.n84 585
R555 VDD2.n130 VDD2.n129 585
R556 VDD2.n128 VDD2.n127 585
R557 VDD2.n89 VDD2.n88 585
R558 VDD2.n93 VDD2.n91 585
R559 VDD2.n122 VDD2.n121 585
R560 VDD2.n120 VDD2.n119 585
R561 VDD2.n95 VDD2.n94 585
R562 VDD2.n114 VDD2.n113 585
R563 VDD2.n112 VDD2.n111 585
R564 VDD2.n99 VDD2.n98 585
R565 VDD2.n106 VDD2.n105 585
R566 VDD2.n104 VDD2.n103 585
R567 VDD2.n25 VDD2.n24 585
R568 VDD2.n27 VDD2.n26 585
R569 VDD2.n20 VDD2.n19 585
R570 VDD2.n33 VDD2.n32 585
R571 VDD2.n35 VDD2.n34 585
R572 VDD2.n16 VDD2.n15 585
R573 VDD2.n42 VDD2.n41 585
R574 VDD2.n43 VDD2.n14 585
R575 VDD2.n45 VDD2.n44 585
R576 VDD2.n12 VDD2.n11 585
R577 VDD2.n51 VDD2.n50 585
R578 VDD2.n53 VDD2.n52 585
R579 VDD2.n8 VDD2.n7 585
R580 VDD2.n59 VDD2.n58 585
R581 VDD2.n61 VDD2.n60 585
R582 VDD2.n4 VDD2.n3 585
R583 VDD2.n67 VDD2.n66 585
R584 VDD2.n69 VDD2.n68 585
R585 VDD2.n102 VDD2.t1 329.036
R586 VDD2.n23 VDD2.t0 329.036
R587 VDD2.n145 VDD2.n144 171.744
R588 VDD2.n144 VDD2.n80 171.744
R589 VDD2.n137 VDD2.n80 171.744
R590 VDD2.n137 VDD2.n136 171.744
R591 VDD2.n136 VDD2.n84 171.744
R592 VDD2.n129 VDD2.n84 171.744
R593 VDD2.n129 VDD2.n128 171.744
R594 VDD2.n128 VDD2.n88 171.744
R595 VDD2.n93 VDD2.n88 171.744
R596 VDD2.n121 VDD2.n93 171.744
R597 VDD2.n121 VDD2.n120 171.744
R598 VDD2.n120 VDD2.n94 171.744
R599 VDD2.n113 VDD2.n94 171.744
R600 VDD2.n113 VDD2.n112 171.744
R601 VDD2.n112 VDD2.n98 171.744
R602 VDD2.n105 VDD2.n98 171.744
R603 VDD2.n105 VDD2.n104 171.744
R604 VDD2.n26 VDD2.n25 171.744
R605 VDD2.n26 VDD2.n19 171.744
R606 VDD2.n33 VDD2.n19 171.744
R607 VDD2.n34 VDD2.n33 171.744
R608 VDD2.n34 VDD2.n15 171.744
R609 VDD2.n42 VDD2.n15 171.744
R610 VDD2.n43 VDD2.n42 171.744
R611 VDD2.n44 VDD2.n43 171.744
R612 VDD2.n44 VDD2.n11 171.744
R613 VDD2.n51 VDD2.n11 171.744
R614 VDD2.n52 VDD2.n51 171.744
R615 VDD2.n52 VDD2.n7 171.744
R616 VDD2.n59 VDD2.n7 171.744
R617 VDD2.n60 VDD2.n59 171.744
R618 VDD2.n60 VDD2.n3 171.744
R619 VDD2.n67 VDD2.n3 171.744
R620 VDD2.n68 VDD2.n67 171.744
R621 VDD2.n104 VDD2.t1 85.8723
R622 VDD2.n25 VDD2.t0 85.8723
R623 VDD2.n76 VDD2.n75 71.76
R624 VDD2 VDD2.n153 71.7572
R625 VDD2.n152 VDD2.n151 70.9233
R626 VDD2.n74 VDD2.n73 70.9231
R627 VDD2.n74 VDD2.n72 48.6962
R628 VDD2.n150 VDD2.n149 47.5066
R629 VDD2.n150 VDD2.n76 40.9955
R630 VDD2.n91 VDD2.n89 13.1884
R631 VDD2.n45 VDD2.n12 13.1884
R632 VDD2.n127 VDD2.n126 12.8005
R633 VDD2.n123 VDD2.n122 12.8005
R634 VDD2.n46 VDD2.n14 12.8005
R635 VDD2.n50 VDD2.n49 12.8005
R636 VDD2.n130 VDD2.n87 12.0247
R637 VDD2.n119 VDD2.n92 12.0247
R638 VDD2.n41 VDD2.n40 12.0247
R639 VDD2.n53 VDD2.n10 12.0247
R640 VDD2.n131 VDD2.n85 11.249
R641 VDD2.n118 VDD2.n95 11.249
R642 VDD2.n39 VDD2.n16 11.249
R643 VDD2.n54 VDD2.n8 11.249
R644 VDD2.n103 VDD2.n102 10.7239
R645 VDD2.n24 VDD2.n23 10.7239
R646 VDD2.n135 VDD2.n134 10.4732
R647 VDD2.n115 VDD2.n114 10.4732
R648 VDD2.n36 VDD2.n35 10.4732
R649 VDD2.n58 VDD2.n57 10.4732
R650 VDD2.n138 VDD2.n83 9.69747
R651 VDD2.n111 VDD2.n97 9.69747
R652 VDD2.n32 VDD2.n18 9.69747
R653 VDD2.n61 VDD2.n6 9.69747
R654 VDD2.n149 VDD2.n148 9.45567
R655 VDD2.n72 VDD2.n71 9.45567
R656 VDD2.n101 VDD2.n100 9.3005
R657 VDD2.n108 VDD2.n107 9.3005
R658 VDD2.n110 VDD2.n109 9.3005
R659 VDD2.n97 VDD2.n96 9.3005
R660 VDD2.n116 VDD2.n115 9.3005
R661 VDD2.n118 VDD2.n117 9.3005
R662 VDD2.n92 VDD2.n90 9.3005
R663 VDD2.n124 VDD2.n123 9.3005
R664 VDD2.n148 VDD2.n147 9.3005
R665 VDD2.n79 VDD2.n78 9.3005
R666 VDD2.n142 VDD2.n141 9.3005
R667 VDD2.n140 VDD2.n139 9.3005
R668 VDD2.n83 VDD2.n82 9.3005
R669 VDD2.n134 VDD2.n133 9.3005
R670 VDD2.n132 VDD2.n131 9.3005
R671 VDD2.n87 VDD2.n86 9.3005
R672 VDD2.n126 VDD2.n125 9.3005
R673 VDD2.n71 VDD2.n70 9.3005
R674 VDD2.n65 VDD2.n64 9.3005
R675 VDD2.n63 VDD2.n62 9.3005
R676 VDD2.n6 VDD2.n5 9.3005
R677 VDD2.n57 VDD2.n56 9.3005
R678 VDD2.n55 VDD2.n54 9.3005
R679 VDD2.n10 VDD2.n9 9.3005
R680 VDD2.n49 VDD2.n48 9.3005
R681 VDD2.n22 VDD2.n21 9.3005
R682 VDD2.n29 VDD2.n28 9.3005
R683 VDD2.n31 VDD2.n30 9.3005
R684 VDD2.n18 VDD2.n17 9.3005
R685 VDD2.n37 VDD2.n36 9.3005
R686 VDD2.n39 VDD2.n38 9.3005
R687 VDD2.n40 VDD2.n13 9.3005
R688 VDD2.n47 VDD2.n46 9.3005
R689 VDD2.n2 VDD2.n1 9.3005
R690 VDD2.n139 VDD2.n81 8.92171
R691 VDD2.n110 VDD2.n99 8.92171
R692 VDD2.n31 VDD2.n20 8.92171
R693 VDD2.n62 VDD2.n4 8.92171
R694 VDD2.n143 VDD2.n142 8.14595
R695 VDD2.n107 VDD2.n106 8.14595
R696 VDD2.n28 VDD2.n27 8.14595
R697 VDD2.n66 VDD2.n65 8.14595
R698 VDD2.n149 VDD2.n77 7.3702
R699 VDD2.n146 VDD2.n79 7.3702
R700 VDD2.n103 VDD2.n101 7.3702
R701 VDD2.n24 VDD2.n22 7.3702
R702 VDD2.n69 VDD2.n2 7.3702
R703 VDD2.n72 VDD2.n0 7.3702
R704 VDD2.n147 VDD2.n77 6.59444
R705 VDD2.n147 VDD2.n146 6.59444
R706 VDD2.n70 VDD2.n69 6.59444
R707 VDD2.n70 VDD2.n0 6.59444
R708 VDD2.n143 VDD2.n79 5.81868
R709 VDD2.n106 VDD2.n101 5.81868
R710 VDD2.n27 VDD2.n22 5.81868
R711 VDD2.n66 VDD2.n2 5.81868
R712 VDD2.n142 VDD2.n81 5.04292
R713 VDD2.n107 VDD2.n99 5.04292
R714 VDD2.n28 VDD2.n20 5.04292
R715 VDD2.n65 VDD2.n4 5.04292
R716 VDD2.n139 VDD2.n138 4.26717
R717 VDD2.n111 VDD2.n110 4.26717
R718 VDD2.n32 VDD2.n31 4.26717
R719 VDD2.n62 VDD2.n61 4.26717
R720 VDD2.n135 VDD2.n83 3.49141
R721 VDD2.n114 VDD2.n97 3.49141
R722 VDD2.n35 VDD2.n18 3.49141
R723 VDD2.n58 VDD2.n6 3.49141
R724 VDD2.n134 VDD2.n85 2.71565
R725 VDD2.n115 VDD2.n95 2.71565
R726 VDD2.n36 VDD2.n16 2.71565
R727 VDD2.n57 VDD2.n8 2.71565
R728 VDD2.n102 VDD2.n100 2.41282
R729 VDD2.n23 VDD2.n21 2.41282
R730 VDD2.n153 VDD2.t6 2.41006
R731 VDD2.n153 VDD2.t5 2.41006
R732 VDD2.n151 VDD2.t2 2.41006
R733 VDD2.n151 VDD2.t9 2.41006
R734 VDD2.n75 VDD2.t7 2.41006
R735 VDD2.n75 VDD2.t3 2.41006
R736 VDD2.n73 VDD2.t4 2.41006
R737 VDD2.n73 VDD2.t8 2.41006
R738 VDD2.n131 VDD2.n130 1.93989
R739 VDD2.n119 VDD2.n118 1.93989
R740 VDD2.n41 VDD2.n39 1.93989
R741 VDD2.n54 VDD2.n53 1.93989
R742 VDD2.n152 VDD2.n150 1.19016
R743 VDD2.n127 VDD2.n87 1.16414
R744 VDD2.n122 VDD2.n92 1.16414
R745 VDD2.n40 VDD2.n14 1.16414
R746 VDD2.n50 VDD2.n10 1.16414
R747 VDD2.n126 VDD2.n89 0.388379
R748 VDD2.n123 VDD2.n91 0.388379
R749 VDD2.n46 VDD2.n45 0.388379
R750 VDD2.n49 VDD2.n12 0.388379
R751 VDD2 VDD2.n152 0.356103
R752 VDD2.n76 VDD2.n74 0.242568
R753 VDD2.n148 VDD2.n78 0.155672
R754 VDD2.n141 VDD2.n78 0.155672
R755 VDD2.n141 VDD2.n140 0.155672
R756 VDD2.n140 VDD2.n82 0.155672
R757 VDD2.n133 VDD2.n82 0.155672
R758 VDD2.n133 VDD2.n132 0.155672
R759 VDD2.n132 VDD2.n86 0.155672
R760 VDD2.n125 VDD2.n86 0.155672
R761 VDD2.n125 VDD2.n124 0.155672
R762 VDD2.n124 VDD2.n90 0.155672
R763 VDD2.n117 VDD2.n90 0.155672
R764 VDD2.n117 VDD2.n116 0.155672
R765 VDD2.n116 VDD2.n96 0.155672
R766 VDD2.n109 VDD2.n96 0.155672
R767 VDD2.n109 VDD2.n108 0.155672
R768 VDD2.n108 VDD2.n100 0.155672
R769 VDD2.n29 VDD2.n21 0.155672
R770 VDD2.n30 VDD2.n29 0.155672
R771 VDD2.n30 VDD2.n17 0.155672
R772 VDD2.n37 VDD2.n17 0.155672
R773 VDD2.n38 VDD2.n37 0.155672
R774 VDD2.n38 VDD2.n13 0.155672
R775 VDD2.n47 VDD2.n13 0.155672
R776 VDD2.n48 VDD2.n47 0.155672
R777 VDD2.n48 VDD2.n9 0.155672
R778 VDD2.n55 VDD2.n9 0.155672
R779 VDD2.n56 VDD2.n55 0.155672
R780 VDD2.n56 VDD2.n5 0.155672
R781 VDD2.n63 VDD2.n5 0.155672
R782 VDD2.n64 VDD2.n63 0.155672
R783 VDD2.n64 VDD2.n1 0.155672
R784 VDD2.n71 VDD2.n1 0.155672
R785 B.n378 B.n377 585
R786 B.n376 B.n107 585
R787 B.n375 B.n374 585
R788 B.n373 B.n108 585
R789 B.n372 B.n371 585
R790 B.n370 B.n109 585
R791 B.n369 B.n368 585
R792 B.n367 B.n110 585
R793 B.n366 B.n365 585
R794 B.n364 B.n111 585
R795 B.n363 B.n362 585
R796 B.n361 B.n112 585
R797 B.n360 B.n359 585
R798 B.n358 B.n113 585
R799 B.n357 B.n356 585
R800 B.n355 B.n114 585
R801 B.n354 B.n353 585
R802 B.n352 B.n115 585
R803 B.n351 B.n350 585
R804 B.n349 B.n116 585
R805 B.n348 B.n347 585
R806 B.n346 B.n117 585
R807 B.n345 B.n344 585
R808 B.n343 B.n118 585
R809 B.n342 B.n341 585
R810 B.n340 B.n119 585
R811 B.n339 B.n338 585
R812 B.n337 B.n120 585
R813 B.n336 B.n335 585
R814 B.n334 B.n121 585
R815 B.n333 B.n332 585
R816 B.n331 B.n122 585
R817 B.n330 B.n329 585
R818 B.n328 B.n123 585
R819 B.n327 B.n326 585
R820 B.n325 B.n124 585
R821 B.n324 B.n323 585
R822 B.n322 B.n125 585
R823 B.n321 B.n320 585
R824 B.n319 B.n126 585
R825 B.n318 B.n317 585
R826 B.n316 B.n127 585
R827 B.n315 B.n314 585
R828 B.n313 B.n128 585
R829 B.n312 B.n311 585
R830 B.n310 B.n129 585
R831 B.n308 B.n307 585
R832 B.n306 B.n132 585
R833 B.n305 B.n304 585
R834 B.n303 B.n133 585
R835 B.n302 B.n301 585
R836 B.n300 B.n134 585
R837 B.n299 B.n298 585
R838 B.n297 B.n135 585
R839 B.n296 B.n295 585
R840 B.n294 B.n136 585
R841 B.n293 B.n292 585
R842 B.n288 B.n137 585
R843 B.n287 B.n286 585
R844 B.n285 B.n138 585
R845 B.n284 B.n283 585
R846 B.n282 B.n139 585
R847 B.n281 B.n280 585
R848 B.n279 B.n140 585
R849 B.n278 B.n277 585
R850 B.n276 B.n141 585
R851 B.n275 B.n274 585
R852 B.n273 B.n142 585
R853 B.n272 B.n271 585
R854 B.n270 B.n143 585
R855 B.n269 B.n268 585
R856 B.n267 B.n144 585
R857 B.n266 B.n265 585
R858 B.n264 B.n145 585
R859 B.n263 B.n262 585
R860 B.n261 B.n146 585
R861 B.n260 B.n259 585
R862 B.n258 B.n147 585
R863 B.n257 B.n256 585
R864 B.n255 B.n148 585
R865 B.n254 B.n253 585
R866 B.n252 B.n149 585
R867 B.n251 B.n250 585
R868 B.n249 B.n150 585
R869 B.n248 B.n247 585
R870 B.n246 B.n151 585
R871 B.n245 B.n244 585
R872 B.n243 B.n152 585
R873 B.n242 B.n241 585
R874 B.n240 B.n153 585
R875 B.n239 B.n238 585
R876 B.n237 B.n154 585
R877 B.n236 B.n235 585
R878 B.n234 B.n155 585
R879 B.n233 B.n232 585
R880 B.n231 B.n156 585
R881 B.n230 B.n229 585
R882 B.n228 B.n157 585
R883 B.n227 B.n226 585
R884 B.n225 B.n158 585
R885 B.n224 B.n223 585
R886 B.n222 B.n159 585
R887 B.n379 B.n106 585
R888 B.n381 B.n380 585
R889 B.n382 B.n105 585
R890 B.n384 B.n383 585
R891 B.n385 B.n104 585
R892 B.n387 B.n386 585
R893 B.n388 B.n103 585
R894 B.n390 B.n389 585
R895 B.n391 B.n102 585
R896 B.n393 B.n392 585
R897 B.n394 B.n101 585
R898 B.n396 B.n395 585
R899 B.n397 B.n100 585
R900 B.n399 B.n398 585
R901 B.n400 B.n99 585
R902 B.n402 B.n401 585
R903 B.n403 B.n98 585
R904 B.n405 B.n404 585
R905 B.n406 B.n97 585
R906 B.n408 B.n407 585
R907 B.n409 B.n96 585
R908 B.n411 B.n410 585
R909 B.n412 B.n95 585
R910 B.n414 B.n413 585
R911 B.n415 B.n94 585
R912 B.n417 B.n416 585
R913 B.n418 B.n93 585
R914 B.n420 B.n419 585
R915 B.n421 B.n92 585
R916 B.n423 B.n422 585
R917 B.n424 B.n91 585
R918 B.n426 B.n425 585
R919 B.n427 B.n90 585
R920 B.n429 B.n428 585
R921 B.n430 B.n89 585
R922 B.n432 B.n431 585
R923 B.n433 B.n88 585
R924 B.n435 B.n434 585
R925 B.n436 B.n87 585
R926 B.n438 B.n437 585
R927 B.n439 B.n86 585
R928 B.n441 B.n440 585
R929 B.n442 B.n85 585
R930 B.n444 B.n443 585
R931 B.n445 B.n84 585
R932 B.n447 B.n446 585
R933 B.n448 B.n83 585
R934 B.n450 B.n449 585
R935 B.n451 B.n82 585
R936 B.n453 B.n452 585
R937 B.n454 B.n81 585
R938 B.n456 B.n455 585
R939 B.n457 B.n80 585
R940 B.n459 B.n458 585
R941 B.n460 B.n79 585
R942 B.n462 B.n461 585
R943 B.n463 B.n78 585
R944 B.n465 B.n464 585
R945 B.n466 B.n77 585
R946 B.n468 B.n467 585
R947 B.n469 B.n76 585
R948 B.n471 B.n470 585
R949 B.n472 B.n75 585
R950 B.n474 B.n473 585
R951 B.n475 B.n74 585
R952 B.n477 B.n476 585
R953 B.n631 B.n18 585
R954 B.n630 B.n629 585
R955 B.n628 B.n19 585
R956 B.n627 B.n626 585
R957 B.n625 B.n20 585
R958 B.n624 B.n623 585
R959 B.n622 B.n21 585
R960 B.n621 B.n620 585
R961 B.n619 B.n22 585
R962 B.n618 B.n617 585
R963 B.n616 B.n23 585
R964 B.n615 B.n614 585
R965 B.n613 B.n24 585
R966 B.n612 B.n611 585
R967 B.n610 B.n25 585
R968 B.n609 B.n608 585
R969 B.n607 B.n26 585
R970 B.n606 B.n605 585
R971 B.n604 B.n27 585
R972 B.n603 B.n602 585
R973 B.n601 B.n28 585
R974 B.n600 B.n599 585
R975 B.n598 B.n29 585
R976 B.n597 B.n596 585
R977 B.n595 B.n30 585
R978 B.n594 B.n593 585
R979 B.n592 B.n31 585
R980 B.n591 B.n590 585
R981 B.n589 B.n32 585
R982 B.n588 B.n587 585
R983 B.n586 B.n33 585
R984 B.n585 B.n584 585
R985 B.n583 B.n34 585
R986 B.n582 B.n581 585
R987 B.n580 B.n35 585
R988 B.n579 B.n578 585
R989 B.n577 B.n36 585
R990 B.n576 B.n575 585
R991 B.n574 B.n37 585
R992 B.n573 B.n572 585
R993 B.n571 B.n38 585
R994 B.n570 B.n569 585
R995 B.n568 B.n39 585
R996 B.n567 B.n566 585
R997 B.n565 B.n40 585
R998 B.n564 B.n563 585
R999 B.n561 B.n41 585
R1000 B.n560 B.n559 585
R1001 B.n558 B.n44 585
R1002 B.n557 B.n556 585
R1003 B.n555 B.n45 585
R1004 B.n554 B.n553 585
R1005 B.n552 B.n46 585
R1006 B.n551 B.n550 585
R1007 B.n549 B.n47 585
R1008 B.n548 B.n547 585
R1009 B.n546 B.n545 585
R1010 B.n544 B.n51 585
R1011 B.n543 B.n542 585
R1012 B.n541 B.n52 585
R1013 B.n540 B.n539 585
R1014 B.n538 B.n53 585
R1015 B.n537 B.n536 585
R1016 B.n535 B.n54 585
R1017 B.n534 B.n533 585
R1018 B.n532 B.n55 585
R1019 B.n531 B.n530 585
R1020 B.n529 B.n56 585
R1021 B.n528 B.n527 585
R1022 B.n526 B.n57 585
R1023 B.n525 B.n524 585
R1024 B.n523 B.n58 585
R1025 B.n522 B.n521 585
R1026 B.n520 B.n59 585
R1027 B.n519 B.n518 585
R1028 B.n517 B.n60 585
R1029 B.n516 B.n515 585
R1030 B.n514 B.n61 585
R1031 B.n513 B.n512 585
R1032 B.n511 B.n62 585
R1033 B.n510 B.n509 585
R1034 B.n508 B.n63 585
R1035 B.n507 B.n506 585
R1036 B.n505 B.n64 585
R1037 B.n504 B.n503 585
R1038 B.n502 B.n65 585
R1039 B.n501 B.n500 585
R1040 B.n499 B.n66 585
R1041 B.n498 B.n497 585
R1042 B.n496 B.n67 585
R1043 B.n495 B.n494 585
R1044 B.n493 B.n68 585
R1045 B.n492 B.n491 585
R1046 B.n490 B.n69 585
R1047 B.n489 B.n488 585
R1048 B.n487 B.n70 585
R1049 B.n486 B.n485 585
R1050 B.n484 B.n71 585
R1051 B.n483 B.n482 585
R1052 B.n481 B.n72 585
R1053 B.n480 B.n479 585
R1054 B.n478 B.n73 585
R1055 B.n633 B.n632 585
R1056 B.n634 B.n17 585
R1057 B.n636 B.n635 585
R1058 B.n637 B.n16 585
R1059 B.n639 B.n638 585
R1060 B.n640 B.n15 585
R1061 B.n642 B.n641 585
R1062 B.n643 B.n14 585
R1063 B.n645 B.n644 585
R1064 B.n646 B.n13 585
R1065 B.n648 B.n647 585
R1066 B.n649 B.n12 585
R1067 B.n651 B.n650 585
R1068 B.n652 B.n11 585
R1069 B.n654 B.n653 585
R1070 B.n655 B.n10 585
R1071 B.n657 B.n656 585
R1072 B.n658 B.n9 585
R1073 B.n660 B.n659 585
R1074 B.n661 B.n8 585
R1075 B.n663 B.n662 585
R1076 B.n664 B.n7 585
R1077 B.n666 B.n665 585
R1078 B.n667 B.n6 585
R1079 B.n669 B.n668 585
R1080 B.n670 B.n5 585
R1081 B.n672 B.n671 585
R1082 B.n673 B.n4 585
R1083 B.n675 B.n674 585
R1084 B.n676 B.n3 585
R1085 B.n678 B.n677 585
R1086 B.n679 B.n0 585
R1087 B.n2 B.n1 585
R1088 B.n176 B.n175 585
R1089 B.n177 B.n174 585
R1090 B.n179 B.n178 585
R1091 B.n180 B.n173 585
R1092 B.n182 B.n181 585
R1093 B.n183 B.n172 585
R1094 B.n185 B.n184 585
R1095 B.n186 B.n171 585
R1096 B.n188 B.n187 585
R1097 B.n189 B.n170 585
R1098 B.n191 B.n190 585
R1099 B.n192 B.n169 585
R1100 B.n194 B.n193 585
R1101 B.n195 B.n168 585
R1102 B.n197 B.n196 585
R1103 B.n198 B.n167 585
R1104 B.n200 B.n199 585
R1105 B.n201 B.n166 585
R1106 B.n203 B.n202 585
R1107 B.n204 B.n165 585
R1108 B.n206 B.n205 585
R1109 B.n207 B.n164 585
R1110 B.n209 B.n208 585
R1111 B.n210 B.n163 585
R1112 B.n212 B.n211 585
R1113 B.n213 B.n162 585
R1114 B.n215 B.n214 585
R1115 B.n216 B.n161 585
R1116 B.n218 B.n217 585
R1117 B.n219 B.n160 585
R1118 B.n221 B.n220 585
R1119 B.n289 B.t6 512.883
R1120 B.n130 B.t3 512.883
R1121 B.n48 B.t9 512.883
R1122 B.n42 B.t0 512.883
R1123 B.n220 B.n159 458.866
R1124 B.n379 B.n378 458.866
R1125 B.n476 B.n73 458.866
R1126 B.n632 B.n631 458.866
R1127 B.n130 B.t4 429.31
R1128 B.n48 B.t11 429.31
R1129 B.n289 B.t7 429.31
R1130 B.n42 B.t2 429.31
R1131 B.n131 B.t5 402.546
R1132 B.n49 B.t10 402.546
R1133 B.n290 B.t8 402.546
R1134 B.n43 B.t1 402.546
R1135 B.n681 B.n680 256.663
R1136 B.n680 B.n679 235.042
R1137 B.n680 B.n2 235.042
R1138 B.n224 B.n159 163.367
R1139 B.n225 B.n224 163.367
R1140 B.n226 B.n225 163.367
R1141 B.n226 B.n157 163.367
R1142 B.n230 B.n157 163.367
R1143 B.n231 B.n230 163.367
R1144 B.n232 B.n231 163.367
R1145 B.n232 B.n155 163.367
R1146 B.n236 B.n155 163.367
R1147 B.n237 B.n236 163.367
R1148 B.n238 B.n237 163.367
R1149 B.n238 B.n153 163.367
R1150 B.n242 B.n153 163.367
R1151 B.n243 B.n242 163.367
R1152 B.n244 B.n243 163.367
R1153 B.n244 B.n151 163.367
R1154 B.n248 B.n151 163.367
R1155 B.n249 B.n248 163.367
R1156 B.n250 B.n249 163.367
R1157 B.n250 B.n149 163.367
R1158 B.n254 B.n149 163.367
R1159 B.n255 B.n254 163.367
R1160 B.n256 B.n255 163.367
R1161 B.n256 B.n147 163.367
R1162 B.n260 B.n147 163.367
R1163 B.n261 B.n260 163.367
R1164 B.n262 B.n261 163.367
R1165 B.n262 B.n145 163.367
R1166 B.n266 B.n145 163.367
R1167 B.n267 B.n266 163.367
R1168 B.n268 B.n267 163.367
R1169 B.n268 B.n143 163.367
R1170 B.n272 B.n143 163.367
R1171 B.n273 B.n272 163.367
R1172 B.n274 B.n273 163.367
R1173 B.n274 B.n141 163.367
R1174 B.n278 B.n141 163.367
R1175 B.n279 B.n278 163.367
R1176 B.n280 B.n279 163.367
R1177 B.n280 B.n139 163.367
R1178 B.n284 B.n139 163.367
R1179 B.n285 B.n284 163.367
R1180 B.n286 B.n285 163.367
R1181 B.n286 B.n137 163.367
R1182 B.n293 B.n137 163.367
R1183 B.n294 B.n293 163.367
R1184 B.n295 B.n294 163.367
R1185 B.n295 B.n135 163.367
R1186 B.n299 B.n135 163.367
R1187 B.n300 B.n299 163.367
R1188 B.n301 B.n300 163.367
R1189 B.n301 B.n133 163.367
R1190 B.n305 B.n133 163.367
R1191 B.n306 B.n305 163.367
R1192 B.n307 B.n306 163.367
R1193 B.n307 B.n129 163.367
R1194 B.n312 B.n129 163.367
R1195 B.n313 B.n312 163.367
R1196 B.n314 B.n313 163.367
R1197 B.n314 B.n127 163.367
R1198 B.n318 B.n127 163.367
R1199 B.n319 B.n318 163.367
R1200 B.n320 B.n319 163.367
R1201 B.n320 B.n125 163.367
R1202 B.n324 B.n125 163.367
R1203 B.n325 B.n324 163.367
R1204 B.n326 B.n325 163.367
R1205 B.n326 B.n123 163.367
R1206 B.n330 B.n123 163.367
R1207 B.n331 B.n330 163.367
R1208 B.n332 B.n331 163.367
R1209 B.n332 B.n121 163.367
R1210 B.n336 B.n121 163.367
R1211 B.n337 B.n336 163.367
R1212 B.n338 B.n337 163.367
R1213 B.n338 B.n119 163.367
R1214 B.n342 B.n119 163.367
R1215 B.n343 B.n342 163.367
R1216 B.n344 B.n343 163.367
R1217 B.n344 B.n117 163.367
R1218 B.n348 B.n117 163.367
R1219 B.n349 B.n348 163.367
R1220 B.n350 B.n349 163.367
R1221 B.n350 B.n115 163.367
R1222 B.n354 B.n115 163.367
R1223 B.n355 B.n354 163.367
R1224 B.n356 B.n355 163.367
R1225 B.n356 B.n113 163.367
R1226 B.n360 B.n113 163.367
R1227 B.n361 B.n360 163.367
R1228 B.n362 B.n361 163.367
R1229 B.n362 B.n111 163.367
R1230 B.n366 B.n111 163.367
R1231 B.n367 B.n366 163.367
R1232 B.n368 B.n367 163.367
R1233 B.n368 B.n109 163.367
R1234 B.n372 B.n109 163.367
R1235 B.n373 B.n372 163.367
R1236 B.n374 B.n373 163.367
R1237 B.n374 B.n107 163.367
R1238 B.n378 B.n107 163.367
R1239 B.n476 B.n475 163.367
R1240 B.n475 B.n474 163.367
R1241 B.n474 B.n75 163.367
R1242 B.n470 B.n75 163.367
R1243 B.n470 B.n469 163.367
R1244 B.n469 B.n468 163.367
R1245 B.n468 B.n77 163.367
R1246 B.n464 B.n77 163.367
R1247 B.n464 B.n463 163.367
R1248 B.n463 B.n462 163.367
R1249 B.n462 B.n79 163.367
R1250 B.n458 B.n79 163.367
R1251 B.n458 B.n457 163.367
R1252 B.n457 B.n456 163.367
R1253 B.n456 B.n81 163.367
R1254 B.n452 B.n81 163.367
R1255 B.n452 B.n451 163.367
R1256 B.n451 B.n450 163.367
R1257 B.n450 B.n83 163.367
R1258 B.n446 B.n83 163.367
R1259 B.n446 B.n445 163.367
R1260 B.n445 B.n444 163.367
R1261 B.n444 B.n85 163.367
R1262 B.n440 B.n85 163.367
R1263 B.n440 B.n439 163.367
R1264 B.n439 B.n438 163.367
R1265 B.n438 B.n87 163.367
R1266 B.n434 B.n87 163.367
R1267 B.n434 B.n433 163.367
R1268 B.n433 B.n432 163.367
R1269 B.n432 B.n89 163.367
R1270 B.n428 B.n89 163.367
R1271 B.n428 B.n427 163.367
R1272 B.n427 B.n426 163.367
R1273 B.n426 B.n91 163.367
R1274 B.n422 B.n91 163.367
R1275 B.n422 B.n421 163.367
R1276 B.n421 B.n420 163.367
R1277 B.n420 B.n93 163.367
R1278 B.n416 B.n93 163.367
R1279 B.n416 B.n415 163.367
R1280 B.n415 B.n414 163.367
R1281 B.n414 B.n95 163.367
R1282 B.n410 B.n95 163.367
R1283 B.n410 B.n409 163.367
R1284 B.n409 B.n408 163.367
R1285 B.n408 B.n97 163.367
R1286 B.n404 B.n97 163.367
R1287 B.n404 B.n403 163.367
R1288 B.n403 B.n402 163.367
R1289 B.n402 B.n99 163.367
R1290 B.n398 B.n99 163.367
R1291 B.n398 B.n397 163.367
R1292 B.n397 B.n396 163.367
R1293 B.n396 B.n101 163.367
R1294 B.n392 B.n101 163.367
R1295 B.n392 B.n391 163.367
R1296 B.n391 B.n390 163.367
R1297 B.n390 B.n103 163.367
R1298 B.n386 B.n103 163.367
R1299 B.n386 B.n385 163.367
R1300 B.n385 B.n384 163.367
R1301 B.n384 B.n105 163.367
R1302 B.n380 B.n105 163.367
R1303 B.n380 B.n379 163.367
R1304 B.n631 B.n630 163.367
R1305 B.n630 B.n19 163.367
R1306 B.n626 B.n19 163.367
R1307 B.n626 B.n625 163.367
R1308 B.n625 B.n624 163.367
R1309 B.n624 B.n21 163.367
R1310 B.n620 B.n21 163.367
R1311 B.n620 B.n619 163.367
R1312 B.n619 B.n618 163.367
R1313 B.n618 B.n23 163.367
R1314 B.n614 B.n23 163.367
R1315 B.n614 B.n613 163.367
R1316 B.n613 B.n612 163.367
R1317 B.n612 B.n25 163.367
R1318 B.n608 B.n25 163.367
R1319 B.n608 B.n607 163.367
R1320 B.n607 B.n606 163.367
R1321 B.n606 B.n27 163.367
R1322 B.n602 B.n27 163.367
R1323 B.n602 B.n601 163.367
R1324 B.n601 B.n600 163.367
R1325 B.n600 B.n29 163.367
R1326 B.n596 B.n29 163.367
R1327 B.n596 B.n595 163.367
R1328 B.n595 B.n594 163.367
R1329 B.n594 B.n31 163.367
R1330 B.n590 B.n31 163.367
R1331 B.n590 B.n589 163.367
R1332 B.n589 B.n588 163.367
R1333 B.n588 B.n33 163.367
R1334 B.n584 B.n33 163.367
R1335 B.n584 B.n583 163.367
R1336 B.n583 B.n582 163.367
R1337 B.n582 B.n35 163.367
R1338 B.n578 B.n35 163.367
R1339 B.n578 B.n577 163.367
R1340 B.n577 B.n576 163.367
R1341 B.n576 B.n37 163.367
R1342 B.n572 B.n37 163.367
R1343 B.n572 B.n571 163.367
R1344 B.n571 B.n570 163.367
R1345 B.n570 B.n39 163.367
R1346 B.n566 B.n39 163.367
R1347 B.n566 B.n565 163.367
R1348 B.n565 B.n564 163.367
R1349 B.n564 B.n41 163.367
R1350 B.n559 B.n41 163.367
R1351 B.n559 B.n558 163.367
R1352 B.n558 B.n557 163.367
R1353 B.n557 B.n45 163.367
R1354 B.n553 B.n45 163.367
R1355 B.n553 B.n552 163.367
R1356 B.n552 B.n551 163.367
R1357 B.n551 B.n47 163.367
R1358 B.n547 B.n47 163.367
R1359 B.n547 B.n546 163.367
R1360 B.n546 B.n51 163.367
R1361 B.n542 B.n51 163.367
R1362 B.n542 B.n541 163.367
R1363 B.n541 B.n540 163.367
R1364 B.n540 B.n53 163.367
R1365 B.n536 B.n53 163.367
R1366 B.n536 B.n535 163.367
R1367 B.n535 B.n534 163.367
R1368 B.n534 B.n55 163.367
R1369 B.n530 B.n55 163.367
R1370 B.n530 B.n529 163.367
R1371 B.n529 B.n528 163.367
R1372 B.n528 B.n57 163.367
R1373 B.n524 B.n57 163.367
R1374 B.n524 B.n523 163.367
R1375 B.n523 B.n522 163.367
R1376 B.n522 B.n59 163.367
R1377 B.n518 B.n59 163.367
R1378 B.n518 B.n517 163.367
R1379 B.n517 B.n516 163.367
R1380 B.n516 B.n61 163.367
R1381 B.n512 B.n61 163.367
R1382 B.n512 B.n511 163.367
R1383 B.n511 B.n510 163.367
R1384 B.n510 B.n63 163.367
R1385 B.n506 B.n63 163.367
R1386 B.n506 B.n505 163.367
R1387 B.n505 B.n504 163.367
R1388 B.n504 B.n65 163.367
R1389 B.n500 B.n65 163.367
R1390 B.n500 B.n499 163.367
R1391 B.n499 B.n498 163.367
R1392 B.n498 B.n67 163.367
R1393 B.n494 B.n67 163.367
R1394 B.n494 B.n493 163.367
R1395 B.n493 B.n492 163.367
R1396 B.n492 B.n69 163.367
R1397 B.n488 B.n69 163.367
R1398 B.n488 B.n487 163.367
R1399 B.n487 B.n486 163.367
R1400 B.n486 B.n71 163.367
R1401 B.n482 B.n71 163.367
R1402 B.n482 B.n481 163.367
R1403 B.n481 B.n480 163.367
R1404 B.n480 B.n73 163.367
R1405 B.n632 B.n17 163.367
R1406 B.n636 B.n17 163.367
R1407 B.n637 B.n636 163.367
R1408 B.n638 B.n637 163.367
R1409 B.n638 B.n15 163.367
R1410 B.n642 B.n15 163.367
R1411 B.n643 B.n642 163.367
R1412 B.n644 B.n643 163.367
R1413 B.n644 B.n13 163.367
R1414 B.n648 B.n13 163.367
R1415 B.n649 B.n648 163.367
R1416 B.n650 B.n649 163.367
R1417 B.n650 B.n11 163.367
R1418 B.n654 B.n11 163.367
R1419 B.n655 B.n654 163.367
R1420 B.n656 B.n655 163.367
R1421 B.n656 B.n9 163.367
R1422 B.n660 B.n9 163.367
R1423 B.n661 B.n660 163.367
R1424 B.n662 B.n661 163.367
R1425 B.n662 B.n7 163.367
R1426 B.n666 B.n7 163.367
R1427 B.n667 B.n666 163.367
R1428 B.n668 B.n667 163.367
R1429 B.n668 B.n5 163.367
R1430 B.n672 B.n5 163.367
R1431 B.n673 B.n672 163.367
R1432 B.n674 B.n673 163.367
R1433 B.n674 B.n3 163.367
R1434 B.n678 B.n3 163.367
R1435 B.n679 B.n678 163.367
R1436 B.n176 B.n2 163.367
R1437 B.n177 B.n176 163.367
R1438 B.n178 B.n177 163.367
R1439 B.n178 B.n173 163.367
R1440 B.n182 B.n173 163.367
R1441 B.n183 B.n182 163.367
R1442 B.n184 B.n183 163.367
R1443 B.n184 B.n171 163.367
R1444 B.n188 B.n171 163.367
R1445 B.n189 B.n188 163.367
R1446 B.n190 B.n189 163.367
R1447 B.n190 B.n169 163.367
R1448 B.n194 B.n169 163.367
R1449 B.n195 B.n194 163.367
R1450 B.n196 B.n195 163.367
R1451 B.n196 B.n167 163.367
R1452 B.n200 B.n167 163.367
R1453 B.n201 B.n200 163.367
R1454 B.n202 B.n201 163.367
R1455 B.n202 B.n165 163.367
R1456 B.n206 B.n165 163.367
R1457 B.n207 B.n206 163.367
R1458 B.n208 B.n207 163.367
R1459 B.n208 B.n163 163.367
R1460 B.n212 B.n163 163.367
R1461 B.n213 B.n212 163.367
R1462 B.n214 B.n213 163.367
R1463 B.n214 B.n161 163.367
R1464 B.n218 B.n161 163.367
R1465 B.n219 B.n218 163.367
R1466 B.n220 B.n219 163.367
R1467 B.n291 B.n290 59.5399
R1468 B.n309 B.n131 59.5399
R1469 B.n50 B.n49 59.5399
R1470 B.n562 B.n43 59.5399
R1471 B.n377 B.n106 29.8151
R1472 B.n633 B.n18 29.8151
R1473 B.n478 B.n477 29.8151
R1474 B.n222 B.n221 29.8151
R1475 B.n290 B.n289 26.7641
R1476 B.n131 B.n130 26.7641
R1477 B.n49 B.n48 26.7641
R1478 B.n43 B.n42 26.7641
R1479 B B.n681 18.0485
R1480 B.n634 B.n633 10.6151
R1481 B.n635 B.n634 10.6151
R1482 B.n635 B.n16 10.6151
R1483 B.n639 B.n16 10.6151
R1484 B.n640 B.n639 10.6151
R1485 B.n641 B.n640 10.6151
R1486 B.n641 B.n14 10.6151
R1487 B.n645 B.n14 10.6151
R1488 B.n646 B.n645 10.6151
R1489 B.n647 B.n646 10.6151
R1490 B.n647 B.n12 10.6151
R1491 B.n651 B.n12 10.6151
R1492 B.n652 B.n651 10.6151
R1493 B.n653 B.n652 10.6151
R1494 B.n653 B.n10 10.6151
R1495 B.n657 B.n10 10.6151
R1496 B.n658 B.n657 10.6151
R1497 B.n659 B.n658 10.6151
R1498 B.n659 B.n8 10.6151
R1499 B.n663 B.n8 10.6151
R1500 B.n664 B.n663 10.6151
R1501 B.n665 B.n664 10.6151
R1502 B.n665 B.n6 10.6151
R1503 B.n669 B.n6 10.6151
R1504 B.n670 B.n669 10.6151
R1505 B.n671 B.n670 10.6151
R1506 B.n671 B.n4 10.6151
R1507 B.n675 B.n4 10.6151
R1508 B.n676 B.n675 10.6151
R1509 B.n677 B.n676 10.6151
R1510 B.n677 B.n0 10.6151
R1511 B.n629 B.n18 10.6151
R1512 B.n629 B.n628 10.6151
R1513 B.n628 B.n627 10.6151
R1514 B.n627 B.n20 10.6151
R1515 B.n623 B.n20 10.6151
R1516 B.n623 B.n622 10.6151
R1517 B.n622 B.n621 10.6151
R1518 B.n621 B.n22 10.6151
R1519 B.n617 B.n22 10.6151
R1520 B.n617 B.n616 10.6151
R1521 B.n616 B.n615 10.6151
R1522 B.n615 B.n24 10.6151
R1523 B.n611 B.n24 10.6151
R1524 B.n611 B.n610 10.6151
R1525 B.n610 B.n609 10.6151
R1526 B.n609 B.n26 10.6151
R1527 B.n605 B.n26 10.6151
R1528 B.n605 B.n604 10.6151
R1529 B.n604 B.n603 10.6151
R1530 B.n603 B.n28 10.6151
R1531 B.n599 B.n28 10.6151
R1532 B.n599 B.n598 10.6151
R1533 B.n598 B.n597 10.6151
R1534 B.n597 B.n30 10.6151
R1535 B.n593 B.n30 10.6151
R1536 B.n593 B.n592 10.6151
R1537 B.n592 B.n591 10.6151
R1538 B.n591 B.n32 10.6151
R1539 B.n587 B.n32 10.6151
R1540 B.n587 B.n586 10.6151
R1541 B.n586 B.n585 10.6151
R1542 B.n585 B.n34 10.6151
R1543 B.n581 B.n34 10.6151
R1544 B.n581 B.n580 10.6151
R1545 B.n580 B.n579 10.6151
R1546 B.n579 B.n36 10.6151
R1547 B.n575 B.n36 10.6151
R1548 B.n575 B.n574 10.6151
R1549 B.n574 B.n573 10.6151
R1550 B.n573 B.n38 10.6151
R1551 B.n569 B.n38 10.6151
R1552 B.n569 B.n568 10.6151
R1553 B.n568 B.n567 10.6151
R1554 B.n567 B.n40 10.6151
R1555 B.n563 B.n40 10.6151
R1556 B.n561 B.n560 10.6151
R1557 B.n560 B.n44 10.6151
R1558 B.n556 B.n44 10.6151
R1559 B.n556 B.n555 10.6151
R1560 B.n555 B.n554 10.6151
R1561 B.n554 B.n46 10.6151
R1562 B.n550 B.n46 10.6151
R1563 B.n550 B.n549 10.6151
R1564 B.n549 B.n548 10.6151
R1565 B.n545 B.n544 10.6151
R1566 B.n544 B.n543 10.6151
R1567 B.n543 B.n52 10.6151
R1568 B.n539 B.n52 10.6151
R1569 B.n539 B.n538 10.6151
R1570 B.n538 B.n537 10.6151
R1571 B.n537 B.n54 10.6151
R1572 B.n533 B.n54 10.6151
R1573 B.n533 B.n532 10.6151
R1574 B.n532 B.n531 10.6151
R1575 B.n531 B.n56 10.6151
R1576 B.n527 B.n56 10.6151
R1577 B.n527 B.n526 10.6151
R1578 B.n526 B.n525 10.6151
R1579 B.n525 B.n58 10.6151
R1580 B.n521 B.n58 10.6151
R1581 B.n521 B.n520 10.6151
R1582 B.n520 B.n519 10.6151
R1583 B.n519 B.n60 10.6151
R1584 B.n515 B.n60 10.6151
R1585 B.n515 B.n514 10.6151
R1586 B.n514 B.n513 10.6151
R1587 B.n513 B.n62 10.6151
R1588 B.n509 B.n62 10.6151
R1589 B.n509 B.n508 10.6151
R1590 B.n508 B.n507 10.6151
R1591 B.n507 B.n64 10.6151
R1592 B.n503 B.n64 10.6151
R1593 B.n503 B.n502 10.6151
R1594 B.n502 B.n501 10.6151
R1595 B.n501 B.n66 10.6151
R1596 B.n497 B.n66 10.6151
R1597 B.n497 B.n496 10.6151
R1598 B.n496 B.n495 10.6151
R1599 B.n495 B.n68 10.6151
R1600 B.n491 B.n68 10.6151
R1601 B.n491 B.n490 10.6151
R1602 B.n490 B.n489 10.6151
R1603 B.n489 B.n70 10.6151
R1604 B.n485 B.n70 10.6151
R1605 B.n485 B.n484 10.6151
R1606 B.n484 B.n483 10.6151
R1607 B.n483 B.n72 10.6151
R1608 B.n479 B.n72 10.6151
R1609 B.n479 B.n478 10.6151
R1610 B.n477 B.n74 10.6151
R1611 B.n473 B.n74 10.6151
R1612 B.n473 B.n472 10.6151
R1613 B.n472 B.n471 10.6151
R1614 B.n471 B.n76 10.6151
R1615 B.n467 B.n76 10.6151
R1616 B.n467 B.n466 10.6151
R1617 B.n466 B.n465 10.6151
R1618 B.n465 B.n78 10.6151
R1619 B.n461 B.n78 10.6151
R1620 B.n461 B.n460 10.6151
R1621 B.n460 B.n459 10.6151
R1622 B.n459 B.n80 10.6151
R1623 B.n455 B.n80 10.6151
R1624 B.n455 B.n454 10.6151
R1625 B.n454 B.n453 10.6151
R1626 B.n453 B.n82 10.6151
R1627 B.n449 B.n82 10.6151
R1628 B.n449 B.n448 10.6151
R1629 B.n448 B.n447 10.6151
R1630 B.n447 B.n84 10.6151
R1631 B.n443 B.n84 10.6151
R1632 B.n443 B.n442 10.6151
R1633 B.n442 B.n441 10.6151
R1634 B.n441 B.n86 10.6151
R1635 B.n437 B.n86 10.6151
R1636 B.n437 B.n436 10.6151
R1637 B.n436 B.n435 10.6151
R1638 B.n435 B.n88 10.6151
R1639 B.n431 B.n88 10.6151
R1640 B.n431 B.n430 10.6151
R1641 B.n430 B.n429 10.6151
R1642 B.n429 B.n90 10.6151
R1643 B.n425 B.n90 10.6151
R1644 B.n425 B.n424 10.6151
R1645 B.n424 B.n423 10.6151
R1646 B.n423 B.n92 10.6151
R1647 B.n419 B.n92 10.6151
R1648 B.n419 B.n418 10.6151
R1649 B.n418 B.n417 10.6151
R1650 B.n417 B.n94 10.6151
R1651 B.n413 B.n94 10.6151
R1652 B.n413 B.n412 10.6151
R1653 B.n412 B.n411 10.6151
R1654 B.n411 B.n96 10.6151
R1655 B.n407 B.n96 10.6151
R1656 B.n407 B.n406 10.6151
R1657 B.n406 B.n405 10.6151
R1658 B.n405 B.n98 10.6151
R1659 B.n401 B.n98 10.6151
R1660 B.n401 B.n400 10.6151
R1661 B.n400 B.n399 10.6151
R1662 B.n399 B.n100 10.6151
R1663 B.n395 B.n100 10.6151
R1664 B.n395 B.n394 10.6151
R1665 B.n394 B.n393 10.6151
R1666 B.n393 B.n102 10.6151
R1667 B.n389 B.n102 10.6151
R1668 B.n389 B.n388 10.6151
R1669 B.n388 B.n387 10.6151
R1670 B.n387 B.n104 10.6151
R1671 B.n383 B.n104 10.6151
R1672 B.n383 B.n382 10.6151
R1673 B.n382 B.n381 10.6151
R1674 B.n381 B.n106 10.6151
R1675 B.n175 B.n1 10.6151
R1676 B.n175 B.n174 10.6151
R1677 B.n179 B.n174 10.6151
R1678 B.n180 B.n179 10.6151
R1679 B.n181 B.n180 10.6151
R1680 B.n181 B.n172 10.6151
R1681 B.n185 B.n172 10.6151
R1682 B.n186 B.n185 10.6151
R1683 B.n187 B.n186 10.6151
R1684 B.n187 B.n170 10.6151
R1685 B.n191 B.n170 10.6151
R1686 B.n192 B.n191 10.6151
R1687 B.n193 B.n192 10.6151
R1688 B.n193 B.n168 10.6151
R1689 B.n197 B.n168 10.6151
R1690 B.n198 B.n197 10.6151
R1691 B.n199 B.n198 10.6151
R1692 B.n199 B.n166 10.6151
R1693 B.n203 B.n166 10.6151
R1694 B.n204 B.n203 10.6151
R1695 B.n205 B.n204 10.6151
R1696 B.n205 B.n164 10.6151
R1697 B.n209 B.n164 10.6151
R1698 B.n210 B.n209 10.6151
R1699 B.n211 B.n210 10.6151
R1700 B.n211 B.n162 10.6151
R1701 B.n215 B.n162 10.6151
R1702 B.n216 B.n215 10.6151
R1703 B.n217 B.n216 10.6151
R1704 B.n217 B.n160 10.6151
R1705 B.n221 B.n160 10.6151
R1706 B.n223 B.n222 10.6151
R1707 B.n223 B.n158 10.6151
R1708 B.n227 B.n158 10.6151
R1709 B.n228 B.n227 10.6151
R1710 B.n229 B.n228 10.6151
R1711 B.n229 B.n156 10.6151
R1712 B.n233 B.n156 10.6151
R1713 B.n234 B.n233 10.6151
R1714 B.n235 B.n234 10.6151
R1715 B.n235 B.n154 10.6151
R1716 B.n239 B.n154 10.6151
R1717 B.n240 B.n239 10.6151
R1718 B.n241 B.n240 10.6151
R1719 B.n241 B.n152 10.6151
R1720 B.n245 B.n152 10.6151
R1721 B.n246 B.n245 10.6151
R1722 B.n247 B.n246 10.6151
R1723 B.n247 B.n150 10.6151
R1724 B.n251 B.n150 10.6151
R1725 B.n252 B.n251 10.6151
R1726 B.n253 B.n252 10.6151
R1727 B.n253 B.n148 10.6151
R1728 B.n257 B.n148 10.6151
R1729 B.n258 B.n257 10.6151
R1730 B.n259 B.n258 10.6151
R1731 B.n259 B.n146 10.6151
R1732 B.n263 B.n146 10.6151
R1733 B.n264 B.n263 10.6151
R1734 B.n265 B.n264 10.6151
R1735 B.n265 B.n144 10.6151
R1736 B.n269 B.n144 10.6151
R1737 B.n270 B.n269 10.6151
R1738 B.n271 B.n270 10.6151
R1739 B.n271 B.n142 10.6151
R1740 B.n275 B.n142 10.6151
R1741 B.n276 B.n275 10.6151
R1742 B.n277 B.n276 10.6151
R1743 B.n277 B.n140 10.6151
R1744 B.n281 B.n140 10.6151
R1745 B.n282 B.n281 10.6151
R1746 B.n283 B.n282 10.6151
R1747 B.n283 B.n138 10.6151
R1748 B.n287 B.n138 10.6151
R1749 B.n288 B.n287 10.6151
R1750 B.n292 B.n288 10.6151
R1751 B.n296 B.n136 10.6151
R1752 B.n297 B.n296 10.6151
R1753 B.n298 B.n297 10.6151
R1754 B.n298 B.n134 10.6151
R1755 B.n302 B.n134 10.6151
R1756 B.n303 B.n302 10.6151
R1757 B.n304 B.n303 10.6151
R1758 B.n304 B.n132 10.6151
R1759 B.n308 B.n132 10.6151
R1760 B.n311 B.n310 10.6151
R1761 B.n311 B.n128 10.6151
R1762 B.n315 B.n128 10.6151
R1763 B.n316 B.n315 10.6151
R1764 B.n317 B.n316 10.6151
R1765 B.n317 B.n126 10.6151
R1766 B.n321 B.n126 10.6151
R1767 B.n322 B.n321 10.6151
R1768 B.n323 B.n322 10.6151
R1769 B.n323 B.n124 10.6151
R1770 B.n327 B.n124 10.6151
R1771 B.n328 B.n327 10.6151
R1772 B.n329 B.n328 10.6151
R1773 B.n329 B.n122 10.6151
R1774 B.n333 B.n122 10.6151
R1775 B.n334 B.n333 10.6151
R1776 B.n335 B.n334 10.6151
R1777 B.n335 B.n120 10.6151
R1778 B.n339 B.n120 10.6151
R1779 B.n340 B.n339 10.6151
R1780 B.n341 B.n340 10.6151
R1781 B.n341 B.n118 10.6151
R1782 B.n345 B.n118 10.6151
R1783 B.n346 B.n345 10.6151
R1784 B.n347 B.n346 10.6151
R1785 B.n347 B.n116 10.6151
R1786 B.n351 B.n116 10.6151
R1787 B.n352 B.n351 10.6151
R1788 B.n353 B.n352 10.6151
R1789 B.n353 B.n114 10.6151
R1790 B.n357 B.n114 10.6151
R1791 B.n358 B.n357 10.6151
R1792 B.n359 B.n358 10.6151
R1793 B.n359 B.n112 10.6151
R1794 B.n363 B.n112 10.6151
R1795 B.n364 B.n363 10.6151
R1796 B.n365 B.n364 10.6151
R1797 B.n365 B.n110 10.6151
R1798 B.n369 B.n110 10.6151
R1799 B.n370 B.n369 10.6151
R1800 B.n371 B.n370 10.6151
R1801 B.n371 B.n108 10.6151
R1802 B.n375 B.n108 10.6151
R1803 B.n376 B.n375 10.6151
R1804 B.n377 B.n376 10.6151
R1805 B.n563 B.n562 9.36635
R1806 B.n545 B.n50 9.36635
R1807 B.n292 B.n291 9.36635
R1808 B.n310 B.n309 9.36635
R1809 B.n681 B.n0 8.11757
R1810 B.n681 B.n1 8.11757
R1811 B.n562 B.n561 1.24928
R1812 B.n548 B.n50 1.24928
R1813 B.n291 B.n136 1.24928
R1814 B.n309 B.n308 1.24928
R1815 VP.n9 VP.t4 362.413
R1816 VP.n25 VP.t5 347.271
R1817 VP.n41 VP.t0 347.271
R1818 VP.n22 VP.t7 347.271
R1819 VP.n26 VP.t1 309.628
R1820 VP.n33 VP.t8 309.628
R1821 VP.n39 VP.t6 309.628
R1822 VP.n20 VP.t9 309.628
R1823 VP.n14 VP.t2 309.628
R1824 VP.n8 VP.t3 309.628
R1825 VP.n10 VP.n7 161.3
R1826 VP.n12 VP.n11 161.3
R1827 VP.n13 VP.n6 161.3
R1828 VP.n16 VP.n15 161.3
R1829 VP.n17 VP.n5 161.3
R1830 VP.n19 VP.n18 161.3
R1831 VP.n21 VP.n4 161.3
R1832 VP.n40 VP.n0 161.3
R1833 VP.n38 VP.n37 161.3
R1834 VP.n36 VP.n1 161.3
R1835 VP.n35 VP.n34 161.3
R1836 VP.n32 VP.n2 161.3
R1837 VP.n31 VP.n30 161.3
R1838 VP.n29 VP.n3 161.3
R1839 VP.n28 VP.n27 161.3
R1840 VP.n23 VP.n22 80.6037
R1841 VP.n42 VP.n41 80.6037
R1842 VP.n25 VP.n24 80.6037
R1843 VP.n27 VP.n25 55.7853
R1844 VP.n41 VP.n40 55.7853
R1845 VP.n22 VP.n21 55.7853
R1846 VP.n9 VP.n8 48.3043
R1847 VP.n32 VP.n31 46.321
R1848 VP.n34 VP.n1 46.321
R1849 VP.n15 VP.n5 46.321
R1850 VP.n13 VP.n12 46.321
R1851 VP.n24 VP.n23 46.0544
R1852 VP.n10 VP.n9 43.9769
R1853 VP.n31 VP.n3 34.6658
R1854 VP.n38 VP.n1 34.6658
R1855 VP.n19 VP.n5 34.6658
R1856 VP.n12 VP.n7 34.6658
R1857 VP.n27 VP.n26 18.1061
R1858 VP.n40 VP.n39 18.1061
R1859 VP.n21 VP.n20 18.1061
R1860 VP.n33 VP.n32 12.234
R1861 VP.n34 VP.n33 12.234
R1862 VP.n14 VP.n13 12.234
R1863 VP.n15 VP.n14 12.234
R1864 VP.n26 VP.n3 6.36192
R1865 VP.n39 VP.n38 6.36192
R1866 VP.n20 VP.n19 6.36192
R1867 VP.n8 VP.n7 6.36192
R1868 VP.n23 VP.n4 0.285035
R1869 VP.n28 VP.n24 0.285035
R1870 VP.n42 VP.n0 0.285035
R1871 VP.n11 VP.n10 0.189894
R1872 VP.n11 VP.n6 0.189894
R1873 VP.n16 VP.n6 0.189894
R1874 VP.n17 VP.n16 0.189894
R1875 VP.n18 VP.n17 0.189894
R1876 VP.n18 VP.n4 0.189894
R1877 VP.n29 VP.n28 0.189894
R1878 VP.n30 VP.n29 0.189894
R1879 VP.n30 VP.n2 0.189894
R1880 VP.n35 VP.n2 0.189894
R1881 VP.n36 VP.n35 0.189894
R1882 VP.n37 VP.n36 0.189894
R1883 VP.n37 VP.n0 0.189894
R1884 VP VP.n42 0.146778
R1885 VDD1.n68 VDD1.n0 756.745
R1886 VDD1.n143 VDD1.n75 756.745
R1887 VDD1.n69 VDD1.n68 585
R1888 VDD1.n67 VDD1.n66 585
R1889 VDD1.n4 VDD1.n3 585
R1890 VDD1.n61 VDD1.n60 585
R1891 VDD1.n59 VDD1.n58 585
R1892 VDD1.n8 VDD1.n7 585
R1893 VDD1.n53 VDD1.n52 585
R1894 VDD1.n51 VDD1.n50 585
R1895 VDD1.n12 VDD1.n11 585
R1896 VDD1.n16 VDD1.n14 585
R1897 VDD1.n45 VDD1.n44 585
R1898 VDD1.n43 VDD1.n42 585
R1899 VDD1.n18 VDD1.n17 585
R1900 VDD1.n37 VDD1.n36 585
R1901 VDD1.n35 VDD1.n34 585
R1902 VDD1.n22 VDD1.n21 585
R1903 VDD1.n29 VDD1.n28 585
R1904 VDD1.n27 VDD1.n26 585
R1905 VDD1.n100 VDD1.n99 585
R1906 VDD1.n102 VDD1.n101 585
R1907 VDD1.n95 VDD1.n94 585
R1908 VDD1.n108 VDD1.n107 585
R1909 VDD1.n110 VDD1.n109 585
R1910 VDD1.n91 VDD1.n90 585
R1911 VDD1.n117 VDD1.n116 585
R1912 VDD1.n118 VDD1.n89 585
R1913 VDD1.n120 VDD1.n119 585
R1914 VDD1.n87 VDD1.n86 585
R1915 VDD1.n126 VDD1.n125 585
R1916 VDD1.n128 VDD1.n127 585
R1917 VDD1.n83 VDD1.n82 585
R1918 VDD1.n134 VDD1.n133 585
R1919 VDD1.n136 VDD1.n135 585
R1920 VDD1.n79 VDD1.n78 585
R1921 VDD1.n142 VDD1.n141 585
R1922 VDD1.n144 VDD1.n143 585
R1923 VDD1.n25 VDD1.t5 329.036
R1924 VDD1.n98 VDD1.t4 329.036
R1925 VDD1.n68 VDD1.n67 171.744
R1926 VDD1.n67 VDD1.n3 171.744
R1927 VDD1.n60 VDD1.n3 171.744
R1928 VDD1.n60 VDD1.n59 171.744
R1929 VDD1.n59 VDD1.n7 171.744
R1930 VDD1.n52 VDD1.n7 171.744
R1931 VDD1.n52 VDD1.n51 171.744
R1932 VDD1.n51 VDD1.n11 171.744
R1933 VDD1.n16 VDD1.n11 171.744
R1934 VDD1.n44 VDD1.n16 171.744
R1935 VDD1.n44 VDD1.n43 171.744
R1936 VDD1.n43 VDD1.n17 171.744
R1937 VDD1.n36 VDD1.n17 171.744
R1938 VDD1.n36 VDD1.n35 171.744
R1939 VDD1.n35 VDD1.n21 171.744
R1940 VDD1.n28 VDD1.n21 171.744
R1941 VDD1.n28 VDD1.n27 171.744
R1942 VDD1.n101 VDD1.n100 171.744
R1943 VDD1.n101 VDD1.n94 171.744
R1944 VDD1.n108 VDD1.n94 171.744
R1945 VDD1.n109 VDD1.n108 171.744
R1946 VDD1.n109 VDD1.n90 171.744
R1947 VDD1.n117 VDD1.n90 171.744
R1948 VDD1.n118 VDD1.n117 171.744
R1949 VDD1.n119 VDD1.n118 171.744
R1950 VDD1.n119 VDD1.n86 171.744
R1951 VDD1.n126 VDD1.n86 171.744
R1952 VDD1.n127 VDD1.n126 171.744
R1953 VDD1.n127 VDD1.n82 171.744
R1954 VDD1.n134 VDD1.n82 171.744
R1955 VDD1.n135 VDD1.n134 171.744
R1956 VDD1.n135 VDD1.n78 171.744
R1957 VDD1.n142 VDD1.n78 171.744
R1958 VDD1.n143 VDD1.n142 171.744
R1959 VDD1.n27 VDD1.t5 85.8723
R1960 VDD1.n100 VDD1.t4 85.8723
R1961 VDD1.n151 VDD1.n150 71.76
R1962 VDD1.n74 VDD1.n73 70.9233
R1963 VDD1.n153 VDD1.n152 70.9231
R1964 VDD1.n149 VDD1.n148 70.9231
R1965 VDD1.n74 VDD1.n72 48.6962
R1966 VDD1.n149 VDD1.n147 48.6962
R1967 VDD1.n153 VDD1.n151 42.1733
R1968 VDD1.n14 VDD1.n12 13.1884
R1969 VDD1.n120 VDD1.n87 13.1884
R1970 VDD1.n50 VDD1.n49 12.8005
R1971 VDD1.n46 VDD1.n45 12.8005
R1972 VDD1.n121 VDD1.n89 12.8005
R1973 VDD1.n125 VDD1.n124 12.8005
R1974 VDD1.n53 VDD1.n10 12.0247
R1975 VDD1.n42 VDD1.n15 12.0247
R1976 VDD1.n116 VDD1.n115 12.0247
R1977 VDD1.n128 VDD1.n85 12.0247
R1978 VDD1.n54 VDD1.n8 11.249
R1979 VDD1.n41 VDD1.n18 11.249
R1980 VDD1.n114 VDD1.n91 11.249
R1981 VDD1.n129 VDD1.n83 11.249
R1982 VDD1.n26 VDD1.n25 10.7239
R1983 VDD1.n99 VDD1.n98 10.7239
R1984 VDD1.n58 VDD1.n57 10.4732
R1985 VDD1.n38 VDD1.n37 10.4732
R1986 VDD1.n111 VDD1.n110 10.4732
R1987 VDD1.n133 VDD1.n132 10.4732
R1988 VDD1.n61 VDD1.n6 9.69747
R1989 VDD1.n34 VDD1.n20 9.69747
R1990 VDD1.n107 VDD1.n93 9.69747
R1991 VDD1.n136 VDD1.n81 9.69747
R1992 VDD1.n72 VDD1.n71 9.45567
R1993 VDD1.n147 VDD1.n146 9.45567
R1994 VDD1.n24 VDD1.n23 9.3005
R1995 VDD1.n31 VDD1.n30 9.3005
R1996 VDD1.n33 VDD1.n32 9.3005
R1997 VDD1.n20 VDD1.n19 9.3005
R1998 VDD1.n39 VDD1.n38 9.3005
R1999 VDD1.n41 VDD1.n40 9.3005
R2000 VDD1.n15 VDD1.n13 9.3005
R2001 VDD1.n47 VDD1.n46 9.3005
R2002 VDD1.n71 VDD1.n70 9.3005
R2003 VDD1.n2 VDD1.n1 9.3005
R2004 VDD1.n65 VDD1.n64 9.3005
R2005 VDD1.n63 VDD1.n62 9.3005
R2006 VDD1.n6 VDD1.n5 9.3005
R2007 VDD1.n57 VDD1.n56 9.3005
R2008 VDD1.n55 VDD1.n54 9.3005
R2009 VDD1.n10 VDD1.n9 9.3005
R2010 VDD1.n49 VDD1.n48 9.3005
R2011 VDD1.n146 VDD1.n145 9.3005
R2012 VDD1.n140 VDD1.n139 9.3005
R2013 VDD1.n138 VDD1.n137 9.3005
R2014 VDD1.n81 VDD1.n80 9.3005
R2015 VDD1.n132 VDD1.n131 9.3005
R2016 VDD1.n130 VDD1.n129 9.3005
R2017 VDD1.n85 VDD1.n84 9.3005
R2018 VDD1.n124 VDD1.n123 9.3005
R2019 VDD1.n97 VDD1.n96 9.3005
R2020 VDD1.n104 VDD1.n103 9.3005
R2021 VDD1.n106 VDD1.n105 9.3005
R2022 VDD1.n93 VDD1.n92 9.3005
R2023 VDD1.n112 VDD1.n111 9.3005
R2024 VDD1.n114 VDD1.n113 9.3005
R2025 VDD1.n115 VDD1.n88 9.3005
R2026 VDD1.n122 VDD1.n121 9.3005
R2027 VDD1.n77 VDD1.n76 9.3005
R2028 VDD1.n62 VDD1.n4 8.92171
R2029 VDD1.n33 VDD1.n22 8.92171
R2030 VDD1.n106 VDD1.n95 8.92171
R2031 VDD1.n137 VDD1.n79 8.92171
R2032 VDD1.n66 VDD1.n65 8.14595
R2033 VDD1.n30 VDD1.n29 8.14595
R2034 VDD1.n103 VDD1.n102 8.14595
R2035 VDD1.n141 VDD1.n140 8.14595
R2036 VDD1.n72 VDD1.n0 7.3702
R2037 VDD1.n69 VDD1.n2 7.3702
R2038 VDD1.n26 VDD1.n24 7.3702
R2039 VDD1.n99 VDD1.n97 7.3702
R2040 VDD1.n144 VDD1.n77 7.3702
R2041 VDD1.n147 VDD1.n75 7.3702
R2042 VDD1.n70 VDD1.n0 6.59444
R2043 VDD1.n70 VDD1.n69 6.59444
R2044 VDD1.n145 VDD1.n144 6.59444
R2045 VDD1.n145 VDD1.n75 6.59444
R2046 VDD1.n66 VDD1.n2 5.81868
R2047 VDD1.n29 VDD1.n24 5.81868
R2048 VDD1.n102 VDD1.n97 5.81868
R2049 VDD1.n141 VDD1.n77 5.81868
R2050 VDD1.n65 VDD1.n4 5.04292
R2051 VDD1.n30 VDD1.n22 5.04292
R2052 VDD1.n103 VDD1.n95 5.04292
R2053 VDD1.n140 VDD1.n79 5.04292
R2054 VDD1.n62 VDD1.n61 4.26717
R2055 VDD1.n34 VDD1.n33 4.26717
R2056 VDD1.n107 VDD1.n106 4.26717
R2057 VDD1.n137 VDD1.n136 4.26717
R2058 VDD1.n58 VDD1.n6 3.49141
R2059 VDD1.n37 VDD1.n20 3.49141
R2060 VDD1.n110 VDD1.n93 3.49141
R2061 VDD1.n133 VDD1.n81 3.49141
R2062 VDD1.n57 VDD1.n8 2.71565
R2063 VDD1.n38 VDD1.n18 2.71565
R2064 VDD1.n111 VDD1.n91 2.71565
R2065 VDD1.n132 VDD1.n83 2.71565
R2066 VDD1.n25 VDD1.n23 2.41282
R2067 VDD1.n98 VDD1.n96 2.41282
R2068 VDD1.n152 VDD1.t0 2.41006
R2069 VDD1.n152 VDD1.t2 2.41006
R2070 VDD1.n73 VDD1.t6 2.41006
R2071 VDD1.n73 VDD1.t7 2.41006
R2072 VDD1.n150 VDD1.t3 2.41006
R2073 VDD1.n150 VDD1.t9 2.41006
R2074 VDD1.n148 VDD1.t8 2.41006
R2075 VDD1.n148 VDD1.t1 2.41006
R2076 VDD1.n54 VDD1.n53 1.93989
R2077 VDD1.n42 VDD1.n41 1.93989
R2078 VDD1.n116 VDD1.n114 1.93989
R2079 VDD1.n129 VDD1.n128 1.93989
R2080 VDD1.n50 VDD1.n10 1.16414
R2081 VDD1.n45 VDD1.n15 1.16414
R2082 VDD1.n115 VDD1.n89 1.16414
R2083 VDD1.n125 VDD1.n85 1.16414
R2084 VDD1 VDD1.n153 0.834552
R2085 VDD1.n49 VDD1.n12 0.388379
R2086 VDD1.n46 VDD1.n14 0.388379
R2087 VDD1.n121 VDD1.n120 0.388379
R2088 VDD1.n124 VDD1.n87 0.388379
R2089 VDD1 VDD1.n74 0.356103
R2090 VDD1.n151 VDD1.n149 0.242568
R2091 VDD1.n71 VDD1.n1 0.155672
R2092 VDD1.n64 VDD1.n1 0.155672
R2093 VDD1.n64 VDD1.n63 0.155672
R2094 VDD1.n63 VDD1.n5 0.155672
R2095 VDD1.n56 VDD1.n5 0.155672
R2096 VDD1.n56 VDD1.n55 0.155672
R2097 VDD1.n55 VDD1.n9 0.155672
R2098 VDD1.n48 VDD1.n9 0.155672
R2099 VDD1.n48 VDD1.n47 0.155672
R2100 VDD1.n47 VDD1.n13 0.155672
R2101 VDD1.n40 VDD1.n13 0.155672
R2102 VDD1.n40 VDD1.n39 0.155672
R2103 VDD1.n39 VDD1.n19 0.155672
R2104 VDD1.n32 VDD1.n19 0.155672
R2105 VDD1.n32 VDD1.n31 0.155672
R2106 VDD1.n31 VDD1.n23 0.155672
R2107 VDD1.n104 VDD1.n96 0.155672
R2108 VDD1.n105 VDD1.n104 0.155672
R2109 VDD1.n105 VDD1.n92 0.155672
R2110 VDD1.n112 VDD1.n92 0.155672
R2111 VDD1.n113 VDD1.n112 0.155672
R2112 VDD1.n113 VDD1.n88 0.155672
R2113 VDD1.n122 VDD1.n88 0.155672
R2114 VDD1.n123 VDD1.n122 0.155672
R2115 VDD1.n123 VDD1.n84 0.155672
R2116 VDD1.n130 VDD1.n84 0.155672
R2117 VDD1.n131 VDD1.n130 0.155672
R2118 VDD1.n131 VDD1.n80 0.155672
R2119 VDD1.n138 VDD1.n80 0.155672
R2120 VDD1.n139 VDD1.n138 0.155672
R2121 VDD1.n139 VDD1.n76 0.155672
R2122 VDD1.n146 VDD1.n76 0.155672
C0 VTAIL VN 8.99895f
C1 w_n2626_n3666# VP 5.50169f
C2 B VP 1.46436f
C3 w_n2626_n3666# B 8.358099f
C4 VDD2 VN 9.06157f
C5 VDD1 VP 9.29322f
C6 w_n2626_n3666# VDD1 2.29671f
C7 VTAIL VP 9.01351f
C8 B VDD1 1.96491f
C9 VTAIL w_n2626_n3666# 3.25953f
C10 VTAIL B 3.23971f
C11 VTAIL VDD1 13.2416f
C12 VDD2 VP 0.386222f
C13 VDD2 w_n2626_n3666# 2.35971f
C14 VDD2 B 2.02263f
C15 VDD2 VDD1 1.19293f
C16 VDD2 VTAIL 13.278599f
C17 VN VP 6.38605f
C18 VN w_n2626_n3666# 5.16458f
C19 VN B 0.906046f
C20 VN VDD1 0.149756f
C21 VDD2 VSUBS 1.653965f
C22 VDD1 VSUBS 1.338691f
C23 VTAIL VSUBS 0.945809f
C24 VN VSUBS 5.45849f
C25 VP VSUBS 2.342004f
C26 B VSUBS 3.570511f
C27 w_n2626_n3666# VSUBS 0.118265p
C28 VDD1.n0 VSUBS 0.028107f
C29 VDD1.n1 VSUBS 0.025579f
C30 VDD1.n2 VSUBS 0.013745f
C31 VDD1.n3 VSUBS 0.032488f
C32 VDD1.n4 VSUBS 0.014553f
C33 VDD1.n5 VSUBS 0.025579f
C34 VDD1.n6 VSUBS 0.013745f
C35 VDD1.n7 VSUBS 0.032488f
C36 VDD1.n8 VSUBS 0.014553f
C37 VDD1.n9 VSUBS 0.025579f
C38 VDD1.n10 VSUBS 0.013745f
C39 VDD1.n11 VSUBS 0.032488f
C40 VDD1.n12 VSUBS 0.014149f
C41 VDD1.n13 VSUBS 0.025579f
C42 VDD1.n14 VSUBS 0.014149f
C43 VDD1.n15 VSUBS 0.013745f
C44 VDD1.n16 VSUBS 0.032488f
C45 VDD1.n17 VSUBS 0.032488f
C46 VDD1.n18 VSUBS 0.014553f
C47 VDD1.n19 VSUBS 0.025579f
C48 VDD1.n20 VSUBS 0.013745f
C49 VDD1.n21 VSUBS 0.032488f
C50 VDD1.n22 VSUBS 0.014553f
C51 VDD1.n23 VSUBS 1.42375f
C52 VDD1.n24 VSUBS 0.013745f
C53 VDD1.t5 VSUBS 0.070133f
C54 VDD1.n25 VSUBS 0.218676f
C55 VDD1.n26 VSUBS 0.024439f
C56 VDD1.n27 VSUBS 0.024366f
C57 VDD1.n28 VSUBS 0.032488f
C58 VDD1.n29 VSUBS 0.014553f
C59 VDD1.n30 VSUBS 0.013745f
C60 VDD1.n31 VSUBS 0.025579f
C61 VDD1.n32 VSUBS 0.025579f
C62 VDD1.n33 VSUBS 0.013745f
C63 VDD1.n34 VSUBS 0.014553f
C64 VDD1.n35 VSUBS 0.032488f
C65 VDD1.n36 VSUBS 0.032488f
C66 VDD1.n37 VSUBS 0.014553f
C67 VDD1.n38 VSUBS 0.013745f
C68 VDD1.n39 VSUBS 0.025579f
C69 VDD1.n40 VSUBS 0.025579f
C70 VDD1.n41 VSUBS 0.013745f
C71 VDD1.n42 VSUBS 0.014553f
C72 VDD1.n43 VSUBS 0.032488f
C73 VDD1.n44 VSUBS 0.032488f
C74 VDD1.n45 VSUBS 0.014553f
C75 VDD1.n46 VSUBS 0.013745f
C76 VDD1.n47 VSUBS 0.025579f
C77 VDD1.n48 VSUBS 0.025579f
C78 VDD1.n49 VSUBS 0.013745f
C79 VDD1.n50 VSUBS 0.014553f
C80 VDD1.n51 VSUBS 0.032488f
C81 VDD1.n52 VSUBS 0.032488f
C82 VDD1.n53 VSUBS 0.014553f
C83 VDD1.n54 VSUBS 0.013745f
C84 VDD1.n55 VSUBS 0.025579f
C85 VDD1.n56 VSUBS 0.025579f
C86 VDD1.n57 VSUBS 0.013745f
C87 VDD1.n58 VSUBS 0.014553f
C88 VDD1.n59 VSUBS 0.032488f
C89 VDD1.n60 VSUBS 0.032488f
C90 VDD1.n61 VSUBS 0.014553f
C91 VDD1.n62 VSUBS 0.013745f
C92 VDD1.n63 VSUBS 0.025579f
C93 VDD1.n64 VSUBS 0.025579f
C94 VDD1.n65 VSUBS 0.013745f
C95 VDD1.n66 VSUBS 0.014553f
C96 VDD1.n67 VSUBS 0.032488f
C97 VDD1.n68 VSUBS 0.078654f
C98 VDD1.n69 VSUBS 0.014553f
C99 VDD1.n70 VSUBS 0.013745f
C100 VDD1.n71 VSUBS 0.056678f
C101 VDD1.n72 VSUBS 0.060724f
C102 VDD1.t6 VSUBS 0.272672f
C103 VDD1.t7 VSUBS 0.272672f
C104 VDD1.n73 VSUBS 2.16252f
C105 VDD1.n74 VSUBS 0.766785f
C106 VDD1.n75 VSUBS 0.028107f
C107 VDD1.n76 VSUBS 0.025579f
C108 VDD1.n77 VSUBS 0.013745f
C109 VDD1.n78 VSUBS 0.032488f
C110 VDD1.n79 VSUBS 0.014553f
C111 VDD1.n80 VSUBS 0.025579f
C112 VDD1.n81 VSUBS 0.013745f
C113 VDD1.n82 VSUBS 0.032488f
C114 VDD1.n83 VSUBS 0.014553f
C115 VDD1.n84 VSUBS 0.025579f
C116 VDD1.n85 VSUBS 0.013745f
C117 VDD1.n86 VSUBS 0.032488f
C118 VDD1.n87 VSUBS 0.014149f
C119 VDD1.n88 VSUBS 0.025579f
C120 VDD1.n89 VSUBS 0.014553f
C121 VDD1.n90 VSUBS 0.032488f
C122 VDD1.n91 VSUBS 0.014553f
C123 VDD1.n92 VSUBS 0.025579f
C124 VDD1.n93 VSUBS 0.013745f
C125 VDD1.n94 VSUBS 0.032488f
C126 VDD1.n95 VSUBS 0.014553f
C127 VDD1.n96 VSUBS 1.42375f
C128 VDD1.n97 VSUBS 0.013745f
C129 VDD1.t4 VSUBS 0.070133f
C130 VDD1.n98 VSUBS 0.218676f
C131 VDD1.n99 VSUBS 0.024439f
C132 VDD1.n100 VSUBS 0.024366f
C133 VDD1.n101 VSUBS 0.032488f
C134 VDD1.n102 VSUBS 0.014553f
C135 VDD1.n103 VSUBS 0.013745f
C136 VDD1.n104 VSUBS 0.025579f
C137 VDD1.n105 VSUBS 0.025579f
C138 VDD1.n106 VSUBS 0.013745f
C139 VDD1.n107 VSUBS 0.014553f
C140 VDD1.n108 VSUBS 0.032488f
C141 VDD1.n109 VSUBS 0.032488f
C142 VDD1.n110 VSUBS 0.014553f
C143 VDD1.n111 VSUBS 0.013745f
C144 VDD1.n112 VSUBS 0.025579f
C145 VDD1.n113 VSUBS 0.025579f
C146 VDD1.n114 VSUBS 0.013745f
C147 VDD1.n115 VSUBS 0.013745f
C148 VDD1.n116 VSUBS 0.014553f
C149 VDD1.n117 VSUBS 0.032488f
C150 VDD1.n118 VSUBS 0.032488f
C151 VDD1.n119 VSUBS 0.032488f
C152 VDD1.n120 VSUBS 0.014149f
C153 VDD1.n121 VSUBS 0.013745f
C154 VDD1.n122 VSUBS 0.025579f
C155 VDD1.n123 VSUBS 0.025579f
C156 VDD1.n124 VSUBS 0.013745f
C157 VDD1.n125 VSUBS 0.014553f
C158 VDD1.n126 VSUBS 0.032488f
C159 VDD1.n127 VSUBS 0.032488f
C160 VDD1.n128 VSUBS 0.014553f
C161 VDD1.n129 VSUBS 0.013745f
C162 VDD1.n130 VSUBS 0.025579f
C163 VDD1.n131 VSUBS 0.025579f
C164 VDD1.n132 VSUBS 0.013745f
C165 VDD1.n133 VSUBS 0.014553f
C166 VDD1.n134 VSUBS 0.032488f
C167 VDD1.n135 VSUBS 0.032488f
C168 VDD1.n136 VSUBS 0.014553f
C169 VDD1.n137 VSUBS 0.013745f
C170 VDD1.n138 VSUBS 0.025579f
C171 VDD1.n139 VSUBS 0.025579f
C172 VDD1.n140 VSUBS 0.013745f
C173 VDD1.n141 VSUBS 0.014553f
C174 VDD1.n142 VSUBS 0.032488f
C175 VDD1.n143 VSUBS 0.078654f
C176 VDD1.n144 VSUBS 0.014553f
C177 VDD1.n145 VSUBS 0.013745f
C178 VDD1.n146 VSUBS 0.056678f
C179 VDD1.n147 VSUBS 0.060724f
C180 VDD1.t8 VSUBS 0.272672f
C181 VDD1.t1 VSUBS 0.272672f
C182 VDD1.n148 VSUBS 2.16251f
C183 VDD1.n149 VSUBS 0.759887f
C184 VDD1.t3 VSUBS 0.272672f
C185 VDD1.t9 VSUBS 0.272672f
C186 VDD1.n150 VSUBS 2.17038f
C187 VDD1.n151 VSUBS 2.60331f
C188 VDD1.t0 VSUBS 0.272672f
C189 VDD1.t2 VSUBS 0.272672f
C190 VDD1.n152 VSUBS 2.16251f
C191 VDD1.n153 VSUBS 2.99413f
C192 VP.n0 VSUBS 0.059208f
C193 VP.t6 VSUBS 1.71782f
C194 VP.n1 VSUBS 0.037965f
C195 VP.n2 VSUBS 0.044371f
C196 VP.t8 VSUBS 1.71782f
C197 VP.n3 VSUBS 0.059448f
C198 VP.n4 VSUBS 0.059208f
C199 VP.t7 VSUBS 1.7892f
C200 VP.t9 VSUBS 1.71782f
C201 VP.n5 VSUBS 0.037965f
C202 VP.n6 VSUBS 0.044371f
C203 VP.t2 VSUBS 1.71782f
C204 VP.n7 VSUBS 0.059448f
C205 VP.t3 VSUBS 1.71782f
C206 VP.n8 VSUBS 0.667105f
C207 VP.t4 VSUBS 1.81851f
C208 VP.n9 VSUBS 0.69639f
C209 VP.n10 VSUBS 0.192125f
C210 VP.n11 VSUBS 0.044371f
C211 VP.n12 VSUBS 0.037965f
C212 VP.n13 VSUBS 0.064206f
C213 VP.n14 VSUBS 0.627942f
C214 VP.n15 VSUBS 0.064206f
C215 VP.n16 VSUBS 0.044371f
C216 VP.n17 VSUBS 0.044371f
C217 VP.n18 VSUBS 0.044371f
C218 VP.n19 VSUBS 0.059448f
C219 VP.n20 VSUBS 0.627942f
C220 VP.n21 VSUBS 0.062643f
C221 VP.n22 VSUBS 0.701273f
C222 VP.n23 VSUBS 2.14179f
C223 VP.n24 VSUBS 2.17642f
C224 VP.t5 VSUBS 1.7892f
C225 VP.n25 VSUBS 0.701273f
C226 VP.t1 VSUBS 1.71782f
C227 VP.n26 VSUBS 0.627942f
C228 VP.n27 VSUBS 0.062643f
C229 VP.n28 VSUBS 0.059208f
C230 VP.n29 VSUBS 0.044371f
C231 VP.n30 VSUBS 0.044371f
C232 VP.n31 VSUBS 0.037965f
C233 VP.n32 VSUBS 0.064206f
C234 VP.n33 VSUBS 0.627942f
C235 VP.n34 VSUBS 0.064206f
C236 VP.n35 VSUBS 0.044371f
C237 VP.n36 VSUBS 0.044371f
C238 VP.n37 VSUBS 0.044371f
C239 VP.n38 VSUBS 0.059448f
C240 VP.n39 VSUBS 0.627942f
C241 VP.n40 VSUBS 0.062643f
C242 VP.t0 VSUBS 1.7892f
C243 VP.n41 VSUBS 0.701273f
C244 VP.n42 VSUBS 0.041555f
C245 B.n0 VSUBS 0.007084f
C246 B.n1 VSUBS 0.007084f
C247 B.n2 VSUBS 0.010477f
C248 B.n3 VSUBS 0.008029f
C249 B.n4 VSUBS 0.008029f
C250 B.n5 VSUBS 0.008029f
C251 B.n6 VSUBS 0.008029f
C252 B.n7 VSUBS 0.008029f
C253 B.n8 VSUBS 0.008029f
C254 B.n9 VSUBS 0.008029f
C255 B.n10 VSUBS 0.008029f
C256 B.n11 VSUBS 0.008029f
C257 B.n12 VSUBS 0.008029f
C258 B.n13 VSUBS 0.008029f
C259 B.n14 VSUBS 0.008029f
C260 B.n15 VSUBS 0.008029f
C261 B.n16 VSUBS 0.008029f
C262 B.n17 VSUBS 0.008029f
C263 B.n18 VSUBS 0.018356f
C264 B.n19 VSUBS 0.008029f
C265 B.n20 VSUBS 0.008029f
C266 B.n21 VSUBS 0.008029f
C267 B.n22 VSUBS 0.008029f
C268 B.n23 VSUBS 0.008029f
C269 B.n24 VSUBS 0.008029f
C270 B.n25 VSUBS 0.008029f
C271 B.n26 VSUBS 0.008029f
C272 B.n27 VSUBS 0.008029f
C273 B.n28 VSUBS 0.008029f
C274 B.n29 VSUBS 0.008029f
C275 B.n30 VSUBS 0.008029f
C276 B.n31 VSUBS 0.008029f
C277 B.n32 VSUBS 0.008029f
C278 B.n33 VSUBS 0.008029f
C279 B.n34 VSUBS 0.008029f
C280 B.n35 VSUBS 0.008029f
C281 B.n36 VSUBS 0.008029f
C282 B.n37 VSUBS 0.008029f
C283 B.n38 VSUBS 0.008029f
C284 B.n39 VSUBS 0.008029f
C285 B.n40 VSUBS 0.008029f
C286 B.n41 VSUBS 0.008029f
C287 B.t1 VSUBS 0.280717f
C288 B.t2 VSUBS 0.298991f
C289 B.t0 VSUBS 0.685316f
C290 B.n42 VSUBS 0.424699f
C291 B.n43 VSUBS 0.304572f
C292 B.n44 VSUBS 0.008029f
C293 B.n45 VSUBS 0.008029f
C294 B.n46 VSUBS 0.008029f
C295 B.n47 VSUBS 0.008029f
C296 B.t10 VSUBS 0.280721f
C297 B.t11 VSUBS 0.298994f
C298 B.t9 VSUBS 0.685316f
C299 B.n48 VSUBS 0.424696f
C300 B.n49 VSUBS 0.304568f
C301 B.n50 VSUBS 0.018601f
C302 B.n51 VSUBS 0.008029f
C303 B.n52 VSUBS 0.008029f
C304 B.n53 VSUBS 0.008029f
C305 B.n54 VSUBS 0.008029f
C306 B.n55 VSUBS 0.008029f
C307 B.n56 VSUBS 0.008029f
C308 B.n57 VSUBS 0.008029f
C309 B.n58 VSUBS 0.008029f
C310 B.n59 VSUBS 0.008029f
C311 B.n60 VSUBS 0.008029f
C312 B.n61 VSUBS 0.008029f
C313 B.n62 VSUBS 0.008029f
C314 B.n63 VSUBS 0.008029f
C315 B.n64 VSUBS 0.008029f
C316 B.n65 VSUBS 0.008029f
C317 B.n66 VSUBS 0.008029f
C318 B.n67 VSUBS 0.008029f
C319 B.n68 VSUBS 0.008029f
C320 B.n69 VSUBS 0.008029f
C321 B.n70 VSUBS 0.008029f
C322 B.n71 VSUBS 0.008029f
C323 B.n72 VSUBS 0.008029f
C324 B.n73 VSUBS 0.018356f
C325 B.n74 VSUBS 0.008029f
C326 B.n75 VSUBS 0.008029f
C327 B.n76 VSUBS 0.008029f
C328 B.n77 VSUBS 0.008029f
C329 B.n78 VSUBS 0.008029f
C330 B.n79 VSUBS 0.008029f
C331 B.n80 VSUBS 0.008029f
C332 B.n81 VSUBS 0.008029f
C333 B.n82 VSUBS 0.008029f
C334 B.n83 VSUBS 0.008029f
C335 B.n84 VSUBS 0.008029f
C336 B.n85 VSUBS 0.008029f
C337 B.n86 VSUBS 0.008029f
C338 B.n87 VSUBS 0.008029f
C339 B.n88 VSUBS 0.008029f
C340 B.n89 VSUBS 0.008029f
C341 B.n90 VSUBS 0.008029f
C342 B.n91 VSUBS 0.008029f
C343 B.n92 VSUBS 0.008029f
C344 B.n93 VSUBS 0.008029f
C345 B.n94 VSUBS 0.008029f
C346 B.n95 VSUBS 0.008029f
C347 B.n96 VSUBS 0.008029f
C348 B.n97 VSUBS 0.008029f
C349 B.n98 VSUBS 0.008029f
C350 B.n99 VSUBS 0.008029f
C351 B.n100 VSUBS 0.008029f
C352 B.n101 VSUBS 0.008029f
C353 B.n102 VSUBS 0.008029f
C354 B.n103 VSUBS 0.008029f
C355 B.n104 VSUBS 0.008029f
C356 B.n105 VSUBS 0.008029f
C357 B.n106 VSUBS 0.018103f
C358 B.n107 VSUBS 0.008029f
C359 B.n108 VSUBS 0.008029f
C360 B.n109 VSUBS 0.008029f
C361 B.n110 VSUBS 0.008029f
C362 B.n111 VSUBS 0.008029f
C363 B.n112 VSUBS 0.008029f
C364 B.n113 VSUBS 0.008029f
C365 B.n114 VSUBS 0.008029f
C366 B.n115 VSUBS 0.008029f
C367 B.n116 VSUBS 0.008029f
C368 B.n117 VSUBS 0.008029f
C369 B.n118 VSUBS 0.008029f
C370 B.n119 VSUBS 0.008029f
C371 B.n120 VSUBS 0.008029f
C372 B.n121 VSUBS 0.008029f
C373 B.n122 VSUBS 0.008029f
C374 B.n123 VSUBS 0.008029f
C375 B.n124 VSUBS 0.008029f
C376 B.n125 VSUBS 0.008029f
C377 B.n126 VSUBS 0.008029f
C378 B.n127 VSUBS 0.008029f
C379 B.n128 VSUBS 0.008029f
C380 B.n129 VSUBS 0.008029f
C381 B.t5 VSUBS 0.280721f
C382 B.t4 VSUBS 0.298994f
C383 B.t3 VSUBS 0.685316f
C384 B.n130 VSUBS 0.424696f
C385 B.n131 VSUBS 0.304568f
C386 B.n132 VSUBS 0.008029f
C387 B.n133 VSUBS 0.008029f
C388 B.n134 VSUBS 0.008029f
C389 B.n135 VSUBS 0.008029f
C390 B.n136 VSUBS 0.004487f
C391 B.n137 VSUBS 0.008029f
C392 B.n138 VSUBS 0.008029f
C393 B.n139 VSUBS 0.008029f
C394 B.n140 VSUBS 0.008029f
C395 B.n141 VSUBS 0.008029f
C396 B.n142 VSUBS 0.008029f
C397 B.n143 VSUBS 0.008029f
C398 B.n144 VSUBS 0.008029f
C399 B.n145 VSUBS 0.008029f
C400 B.n146 VSUBS 0.008029f
C401 B.n147 VSUBS 0.008029f
C402 B.n148 VSUBS 0.008029f
C403 B.n149 VSUBS 0.008029f
C404 B.n150 VSUBS 0.008029f
C405 B.n151 VSUBS 0.008029f
C406 B.n152 VSUBS 0.008029f
C407 B.n153 VSUBS 0.008029f
C408 B.n154 VSUBS 0.008029f
C409 B.n155 VSUBS 0.008029f
C410 B.n156 VSUBS 0.008029f
C411 B.n157 VSUBS 0.008029f
C412 B.n158 VSUBS 0.008029f
C413 B.n159 VSUBS 0.018356f
C414 B.n160 VSUBS 0.008029f
C415 B.n161 VSUBS 0.008029f
C416 B.n162 VSUBS 0.008029f
C417 B.n163 VSUBS 0.008029f
C418 B.n164 VSUBS 0.008029f
C419 B.n165 VSUBS 0.008029f
C420 B.n166 VSUBS 0.008029f
C421 B.n167 VSUBS 0.008029f
C422 B.n168 VSUBS 0.008029f
C423 B.n169 VSUBS 0.008029f
C424 B.n170 VSUBS 0.008029f
C425 B.n171 VSUBS 0.008029f
C426 B.n172 VSUBS 0.008029f
C427 B.n173 VSUBS 0.008029f
C428 B.n174 VSUBS 0.008029f
C429 B.n175 VSUBS 0.008029f
C430 B.n176 VSUBS 0.008029f
C431 B.n177 VSUBS 0.008029f
C432 B.n178 VSUBS 0.008029f
C433 B.n179 VSUBS 0.008029f
C434 B.n180 VSUBS 0.008029f
C435 B.n181 VSUBS 0.008029f
C436 B.n182 VSUBS 0.008029f
C437 B.n183 VSUBS 0.008029f
C438 B.n184 VSUBS 0.008029f
C439 B.n185 VSUBS 0.008029f
C440 B.n186 VSUBS 0.008029f
C441 B.n187 VSUBS 0.008029f
C442 B.n188 VSUBS 0.008029f
C443 B.n189 VSUBS 0.008029f
C444 B.n190 VSUBS 0.008029f
C445 B.n191 VSUBS 0.008029f
C446 B.n192 VSUBS 0.008029f
C447 B.n193 VSUBS 0.008029f
C448 B.n194 VSUBS 0.008029f
C449 B.n195 VSUBS 0.008029f
C450 B.n196 VSUBS 0.008029f
C451 B.n197 VSUBS 0.008029f
C452 B.n198 VSUBS 0.008029f
C453 B.n199 VSUBS 0.008029f
C454 B.n200 VSUBS 0.008029f
C455 B.n201 VSUBS 0.008029f
C456 B.n202 VSUBS 0.008029f
C457 B.n203 VSUBS 0.008029f
C458 B.n204 VSUBS 0.008029f
C459 B.n205 VSUBS 0.008029f
C460 B.n206 VSUBS 0.008029f
C461 B.n207 VSUBS 0.008029f
C462 B.n208 VSUBS 0.008029f
C463 B.n209 VSUBS 0.008029f
C464 B.n210 VSUBS 0.008029f
C465 B.n211 VSUBS 0.008029f
C466 B.n212 VSUBS 0.008029f
C467 B.n213 VSUBS 0.008029f
C468 B.n214 VSUBS 0.008029f
C469 B.n215 VSUBS 0.008029f
C470 B.n216 VSUBS 0.008029f
C471 B.n217 VSUBS 0.008029f
C472 B.n218 VSUBS 0.008029f
C473 B.n219 VSUBS 0.008029f
C474 B.n220 VSUBS 0.017064f
C475 B.n221 VSUBS 0.017064f
C476 B.n222 VSUBS 0.018356f
C477 B.n223 VSUBS 0.008029f
C478 B.n224 VSUBS 0.008029f
C479 B.n225 VSUBS 0.008029f
C480 B.n226 VSUBS 0.008029f
C481 B.n227 VSUBS 0.008029f
C482 B.n228 VSUBS 0.008029f
C483 B.n229 VSUBS 0.008029f
C484 B.n230 VSUBS 0.008029f
C485 B.n231 VSUBS 0.008029f
C486 B.n232 VSUBS 0.008029f
C487 B.n233 VSUBS 0.008029f
C488 B.n234 VSUBS 0.008029f
C489 B.n235 VSUBS 0.008029f
C490 B.n236 VSUBS 0.008029f
C491 B.n237 VSUBS 0.008029f
C492 B.n238 VSUBS 0.008029f
C493 B.n239 VSUBS 0.008029f
C494 B.n240 VSUBS 0.008029f
C495 B.n241 VSUBS 0.008029f
C496 B.n242 VSUBS 0.008029f
C497 B.n243 VSUBS 0.008029f
C498 B.n244 VSUBS 0.008029f
C499 B.n245 VSUBS 0.008029f
C500 B.n246 VSUBS 0.008029f
C501 B.n247 VSUBS 0.008029f
C502 B.n248 VSUBS 0.008029f
C503 B.n249 VSUBS 0.008029f
C504 B.n250 VSUBS 0.008029f
C505 B.n251 VSUBS 0.008029f
C506 B.n252 VSUBS 0.008029f
C507 B.n253 VSUBS 0.008029f
C508 B.n254 VSUBS 0.008029f
C509 B.n255 VSUBS 0.008029f
C510 B.n256 VSUBS 0.008029f
C511 B.n257 VSUBS 0.008029f
C512 B.n258 VSUBS 0.008029f
C513 B.n259 VSUBS 0.008029f
C514 B.n260 VSUBS 0.008029f
C515 B.n261 VSUBS 0.008029f
C516 B.n262 VSUBS 0.008029f
C517 B.n263 VSUBS 0.008029f
C518 B.n264 VSUBS 0.008029f
C519 B.n265 VSUBS 0.008029f
C520 B.n266 VSUBS 0.008029f
C521 B.n267 VSUBS 0.008029f
C522 B.n268 VSUBS 0.008029f
C523 B.n269 VSUBS 0.008029f
C524 B.n270 VSUBS 0.008029f
C525 B.n271 VSUBS 0.008029f
C526 B.n272 VSUBS 0.008029f
C527 B.n273 VSUBS 0.008029f
C528 B.n274 VSUBS 0.008029f
C529 B.n275 VSUBS 0.008029f
C530 B.n276 VSUBS 0.008029f
C531 B.n277 VSUBS 0.008029f
C532 B.n278 VSUBS 0.008029f
C533 B.n279 VSUBS 0.008029f
C534 B.n280 VSUBS 0.008029f
C535 B.n281 VSUBS 0.008029f
C536 B.n282 VSUBS 0.008029f
C537 B.n283 VSUBS 0.008029f
C538 B.n284 VSUBS 0.008029f
C539 B.n285 VSUBS 0.008029f
C540 B.n286 VSUBS 0.008029f
C541 B.n287 VSUBS 0.008029f
C542 B.n288 VSUBS 0.008029f
C543 B.t8 VSUBS 0.280717f
C544 B.t7 VSUBS 0.298991f
C545 B.t6 VSUBS 0.685316f
C546 B.n289 VSUBS 0.424699f
C547 B.n290 VSUBS 0.304572f
C548 B.n291 VSUBS 0.018601f
C549 B.n292 VSUBS 0.007556f
C550 B.n293 VSUBS 0.008029f
C551 B.n294 VSUBS 0.008029f
C552 B.n295 VSUBS 0.008029f
C553 B.n296 VSUBS 0.008029f
C554 B.n297 VSUBS 0.008029f
C555 B.n298 VSUBS 0.008029f
C556 B.n299 VSUBS 0.008029f
C557 B.n300 VSUBS 0.008029f
C558 B.n301 VSUBS 0.008029f
C559 B.n302 VSUBS 0.008029f
C560 B.n303 VSUBS 0.008029f
C561 B.n304 VSUBS 0.008029f
C562 B.n305 VSUBS 0.008029f
C563 B.n306 VSUBS 0.008029f
C564 B.n307 VSUBS 0.008029f
C565 B.n308 VSUBS 0.004487f
C566 B.n309 VSUBS 0.018601f
C567 B.n310 VSUBS 0.007556f
C568 B.n311 VSUBS 0.008029f
C569 B.n312 VSUBS 0.008029f
C570 B.n313 VSUBS 0.008029f
C571 B.n314 VSUBS 0.008029f
C572 B.n315 VSUBS 0.008029f
C573 B.n316 VSUBS 0.008029f
C574 B.n317 VSUBS 0.008029f
C575 B.n318 VSUBS 0.008029f
C576 B.n319 VSUBS 0.008029f
C577 B.n320 VSUBS 0.008029f
C578 B.n321 VSUBS 0.008029f
C579 B.n322 VSUBS 0.008029f
C580 B.n323 VSUBS 0.008029f
C581 B.n324 VSUBS 0.008029f
C582 B.n325 VSUBS 0.008029f
C583 B.n326 VSUBS 0.008029f
C584 B.n327 VSUBS 0.008029f
C585 B.n328 VSUBS 0.008029f
C586 B.n329 VSUBS 0.008029f
C587 B.n330 VSUBS 0.008029f
C588 B.n331 VSUBS 0.008029f
C589 B.n332 VSUBS 0.008029f
C590 B.n333 VSUBS 0.008029f
C591 B.n334 VSUBS 0.008029f
C592 B.n335 VSUBS 0.008029f
C593 B.n336 VSUBS 0.008029f
C594 B.n337 VSUBS 0.008029f
C595 B.n338 VSUBS 0.008029f
C596 B.n339 VSUBS 0.008029f
C597 B.n340 VSUBS 0.008029f
C598 B.n341 VSUBS 0.008029f
C599 B.n342 VSUBS 0.008029f
C600 B.n343 VSUBS 0.008029f
C601 B.n344 VSUBS 0.008029f
C602 B.n345 VSUBS 0.008029f
C603 B.n346 VSUBS 0.008029f
C604 B.n347 VSUBS 0.008029f
C605 B.n348 VSUBS 0.008029f
C606 B.n349 VSUBS 0.008029f
C607 B.n350 VSUBS 0.008029f
C608 B.n351 VSUBS 0.008029f
C609 B.n352 VSUBS 0.008029f
C610 B.n353 VSUBS 0.008029f
C611 B.n354 VSUBS 0.008029f
C612 B.n355 VSUBS 0.008029f
C613 B.n356 VSUBS 0.008029f
C614 B.n357 VSUBS 0.008029f
C615 B.n358 VSUBS 0.008029f
C616 B.n359 VSUBS 0.008029f
C617 B.n360 VSUBS 0.008029f
C618 B.n361 VSUBS 0.008029f
C619 B.n362 VSUBS 0.008029f
C620 B.n363 VSUBS 0.008029f
C621 B.n364 VSUBS 0.008029f
C622 B.n365 VSUBS 0.008029f
C623 B.n366 VSUBS 0.008029f
C624 B.n367 VSUBS 0.008029f
C625 B.n368 VSUBS 0.008029f
C626 B.n369 VSUBS 0.008029f
C627 B.n370 VSUBS 0.008029f
C628 B.n371 VSUBS 0.008029f
C629 B.n372 VSUBS 0.008029f
C630 B.n373 VSUBS 0.008029f
C631 B.n374 VSUBS 0.008029f
C632 B.n375 VSUBS 0.008029f
C633 B.n376 VSUBS 0.008029f
C634 B.n377 VSUBS 0.017317f
C635 B.n378 VSUBS 0.018356f
C636 B.n379 VSUBS 0.017064f
C637 B.n380 VSUBS 0.008029f
C638 B.n381 VSUBS 0.008029f
C639 B.n382 VSUBS 0.008029f
C640 B.n383 VSUBS 0.008029f
C641 B.n384 VSUBS 0.008029f
C642 B.n385 VSUBS 0.008029f
C643 B.n386 VSUBS 0.008029f
C644 B.n387 VSUBS 0.008029f
C645 B.n388 VSUBS 0.008029f
C646 B.n389 VSUBS 0.008029f
C647 B.n390 VSUBS 0.008029f
C648 B.n391 VSUBS 0.008029f
C649 B.n392 VSUBS 0.008029f
C650 B.n393 VSUBS 0.008029f
C651 B.n394 VSUBS 0.008029f
C652 B.n395 VSUBS 0.008029f
C653 B.n396 VSUBS 0.008029f
C654 B.n397 VSUBS 0.008029f
C655 B.n398 VSUBS 0.008029f
C656 B.n399 VSUBS 0.008029f
C657 B.n400 VSUBS 0.008029f
C658 B.n401 VSUBS 0.008029f
C659 B.n402 VSUBS 0.008029f
C660 B.n403 VSUBS 0.008029f
C661 B.n404 VSUBS 0.008029f
C662 B.n405 VSUBS 0.008029f
C663 B.n406 VSUBS 0.008029f
C664 B.n407 VSUBS 0.008029f
C665 B.n408 VSUBS 0.008029f
C666 B.n409 VSUBS 0.008029f
C667 B.n410 VSUBS 0.008029f
C668 B.n411 VSUBS 0.008029f
C669 B.n412 VSUBS 0.008029f
C670 B.n413 VSUBS 0.008029f
C671 B.n414 VSUBS 0.008029f
C672 B.n415 VSUBS 0.008029f
C673 B.n416 VSUBS 0.008029f
C674 B.n417 VSUBS 0.008029f
C675 B.n418 VSUBS 0.008029f
C676 B.n419 VSUBS 0.008029f
C677 B.n420 VSUBS 0.008029f
C678 B.n421 VSUBS 0.008029f
C679 B.n422 VSUBS 0.008029f
C680 B.n423 VSUBS 0.008029f
C681 B.n424 VSUBS 0.008029f
C682 B.n425 VSUBS 0.008029f
C683 B.n426 VSUBS 0.008029f
C684 B.n427 VSUBS 0.008029f
C685 B.n428 VSUBS 0.008029f
C686 B.n429 VSUBS 0.008029f
C687 B.n430 VSUBS 0.008029f
C688 B.n431 VSUBS 0.008029f
C689 B.n432 VSUBS 0.008029f
C690 B.n433 VSUBS 0.008029f
C691 B.n434 VSUBS 0.008029f
C692 B.n435 VSUBS 0.008029f
C693 B.n436 VSUBS 0.008029f
C694 B.n437 VSUBS 0.008029f
C695 B.n438 VSUBS 0.008029f
C696 B.n439 VSUBS 0.008029f
C697 B.n440 VSUBS 0.008029f
C698 B.n441 VSUBS 0.008029f
C699 B.n442 VSUBS 0.008029f
C700 B.n443 VSUBS 0.008029f
C701 B.n444 VSUBS 0.008029f
C702 B.n445 VSUBS 0.008029f
C703 B.n446 VSUBS 0.008029f
C704 B.n447 VSUBS 0.008029f
C705 B.n448 VSUBS 0.008029f
C706 B.n449 VSUBS 0.008029f
C707 B.n450 VSUBS 0.008029f
C708 B.n451 VSUBS 0.008029f
C709 B.n452 VSUBS 0.008029f
C710 B.n453 VSUBS 0.008029f
C711 B.n454 VSUBS 0.008029f
C712 B.n455 VSUBS 0.008029f
C713 B.n456 VSUBS 0.008029f
C714 B.n457 VSUBS 0.008029f
C715 B.n458 VSUBS 0.008029f
C716 B.n459 VSUBS 0.008029f
C717 B.n460 VSUBS 0.008029f
C718 B.n461 VSUBS 0.008029f
C719 B.n462 VSUBS 0.008029f
C720 B.n463 VSUBS 0.008029f
C721 B.n464 VSUBS 0.008029f
C722 B.n465 VSUBS 0.008029f
C723 B.n466 VSUBS 0.008029f
C724 B.n467 VSUBS 0.008029f
C725 B.n468 VSUBS 0.008029f
C726 B.n469 VSUBS 0.008029f
C727 B.n470 VSUBS 0.008029f
C728 B.n471 VSUBS 0.008029f
C729 B.n472 VSUBS 0.008029f
C730 B.n473 VSUBS 0.008029f
C731 B.n474 VSUBS 0.008029f
C732 B.n475 VSUBS 0.008029f
C733 B.n476 VSUBS 0.017064f
C734 B.n477 VSUBS 0.017064f
C735 B.n478 VSUBS 0.018356f
C736 B.n479 VSUBS 0.008029f
C737 B.n480 VSUBS 0.008029f
C738 B.n481 VSUBS 0.008029f
C739 B.n482 VSUBS 0.008029f
C740 B.n483 VSUBS 0.008029f
C741 B.n484 VSUBS 0.008029f
C742 B.n485 VSUBS 0.008029f
C743 B.n486 VSUBS 0.008029f
C744 B.n487 VSUBS 0.008029f
C745 B.n488 VSUBS 0.008029f
C746 B.n489 VSUBS 0.008029f
C747 B.n490 VSUBS 0.008029f
C748 B.n491 VSUBS 0.008029f
C749 B.n492 VSUBS 0.008029f
C750 B.n493 VSUBS 0.008029f
C751 B.n494 VSUBS 0.008029f
C752 B.n495 VSUBS 0.008029f
C753 B.n496 VSUBS 0.008029f
C754 B.n497 VSUBS 0.008029f
C755 B.n498 VSUBS 0.008029f
C756 B.n499 VSUBS 0.008029f
C757 B.n500 VSUBS 0.008029f
C758 B.n501 VSUBS 0.008029f
C759 B.n502 VSUBS 0.008029f
C760 B.n503 VSUBS 0.008029f
C761 B.n504 VSUBS 0.008029f
C762 B.n505 VSUBS 0.008029f
C763 B.n506 VSUBS 0.008029f
C764 B.n507 VSUBS 0.008029f
C765 B.n508 VSUBS 0.008029f
C766 B.n509 VSUBS 0.008029f
C767 B.n510 VSUBS 0.008029f
C768 B.n511 VSUBS 0.008029f
C769 B.n512 VSUBS 0.008029f
C770 B.n513 VSUBS 0.008029f
C771 B.n514 VSUBS 0.008029f
C772 B.n515 VSUBS 0.008029f
C773 B.n516 VSUBS 0.008029f
C774 B.n517 VSUBS 0.008029f
C775 B.n518 VSUBS 0.008029f
C776 B.n519 VSUBS 0.008029f
C777 B.n520 VSUBS 0.008029f
C778 B.n521 VSUBS 0.008029f
C779 B.n522 VSUBS 0.008029f
C780 B.n523 VSUBS 0.008029f
C781 B.n524 VSUBS 0.008029f
C782 B.n525 VSUBS 0.008029f
C783 B.n526 VSUBS 0.008029f
C784 B.n527 VSUBS 0.008029f
C785 B.n528 VSUBS 0.008029f
C786 B.n529 VSUBS 0.008029f
C787 B.n530 VSUBS 0.008029f
C788 B.n531 VSUBS 0.008029f
C789 B.n532 VSUBS 0.008029f
C790 B.n533 VSUBS 0.008029f
C791 B.n534 VSUBS 0.008029f
C792 B.n535 VSUBS 0.008029f
C793 B.n536 VSUBS 0.008029f
C794 B.n537 VSUBS 0.008029f
C795 B.n538 VSUBS 0.008029f
C796 B.n539 VSUBS 0.008029f
C797 B.n540 VSUBS 0.008029f
C798 B.n541 VSUBS 0.008029f
C799 B.n542 VSUBS 0.008029f
C800 B.n543 VSUBS 0.008029f
C801 B.n544 VSUBS 0.008029f
C802 B.n545 VSUBS 0.007556f
C803 B.n546 VSUBS 0.008029f
C804 B.n547 VSUBS 0.008029f
C805 B.n548 VSUBS 0.004487f
C806 B.n549 VSUBS 0.008029f
C807 B.n550 VSUBS 0.008029f
C808 B.n551 VSUBS 0.008029f
C809 B.n552 VSUBS 0.008029f
C810 B.n553 VSUBS 0.008029f
C811 B.n554 VSUBS 0.008029f
C812 B.n555 VSUBS 0.008029f
C813 B.n556 VSUBS 0.008029f
C814 B.n557 VSUBS 0.008029f
C815 B.n558 VSUBS 0.008029f
C816 B.n559 VSUBS 0.008029f
C817 B.n560 VSUBS 0.008029f
C818 B.n561 VSUBS 0.004487f
C819 B.n562 VSUBS 0.018601f
C820 B.n563 VSUBS 0.007556f
C821 B.n564 VSUBS 0.008029f
C822 B.n565 VSUBS 0.008029f
C823 B.n566 VSUBS 0.008029f
C824 B.n567 VSUBS 0.008029f
C825 B.n568 VSUBS 0.008029f
C826 B.n569 VSUBS 0.008029f
C827 B.n570 VSUBS 0.008029f
C828 B.n571 VSUBS 0.008029f
C829 B.n572 VSUBS 0.008029f
C830 B.n573 VSUBS 0.008029f
C831 B.n574 VSUBS 0.008029f
C832 B.n575 VSUBS 0.008029f
C833 B.n576 VSUBS 0.008029f
C834 B.n577 VSUBS 0.008029f
C835 B.n578 VSUBS 0.008029f
C836 B.n579 VSUBS 0.008029f
C837 B.n580 VSUBS 0.008029f
C838 B.n581 VSUBS 0.008029f
C839 B.n582 VSUBS 0.008029f
C840 B.n583 VSUBS 0.008029f
C841 B.n584 VSUBS 0.008029f
C842 B.n585 VSUBS 0.008029f
C843 B.n586 VSUBS 0.008029f
C844 B.n587 VSUBS 0.008029f
C845 B.n588 VSUBS 0.008029f
C846 B.n589 VSUBS 0.008029f
C847 B.n590 VSUBS 0.008029f
C848 B.n591 VSUBS 0.008029f
C849 B.n592 VSUBS 0.008029f
C850 B.n593 VSUBS 0.008029f
C851 B.n594 VSUBS 0.008029f
C852 B.n595 VSUBS 0.008029f
C853 B.n596 VSUBS 0.008029f
C854 B.n597 VSUBS 0.008029f
C855 B.n598 VSUBS 0.008029f
C856 B.n599 VSUBS 0.008029f
C857 B.n600 VSUBS 0.008029f
C858 B.n601 VSUBS 0.008029f
C859 B.n602 VSUBS 0.008029f
C860 B.n603 VSUBS 0.008029f
C861 B.n604 VSUBS 0.008029f
C862 B.n605 VSUBS 0.008029f
C863 B.n606 VSUBS 0.008029f
C864 B.n607 VSUBS 0.008029f
C865 B.n608 VSUBS 0.008029f
C866 B.n609 VSUBS 0.008029f
C867 B.n610 VSUBS 0.008029f
C868 B.n611 VSUBS 0.008029f
C869 B.n612 VSUBS 0.008029f
C870 B.n613 VSUBS 0.008029f
C871 B.n614 VSUBS 0.008029f
C872 B.n615 VSUBS 0.008029f
C873 B.n616 VSUBS 0.008029f
C874 B.n617 VSUBS 0.008029f
C875 B.n618 VSUBS 0.008029f
C876 B.n619 VSUBS 0.008029f
C877 B.n620 VSUBS 0.008029f
C878 B.n621 VSUBS 0.008029f
C879 B.n622 VSUBS 0.008029f
C880 B.n623 VSUBS 0.008029f
C881 B.n624 VSUBS 0.008029f
C882 B.n625 VSUBS 0.008029f
C883 B.n626 VSUBS 0.008029f
C884 B.n627 VSUBS 0.008029f
C885 B.n628 VSUBS 0.008029f
C886 B.n629 VSUBS 0.008029f
C887 B.n630 VSUBS 0.008029f
C888 B.n631 VSUBS 0.018356f
C889 B.n632 VSUBS 0.017064f
C890 B.n633 VSUBS 0.017064f
C891 B.n634 VSUBS 0.008029f
C892 B.n635 VSUBS 0.008029f
C893 B.n636 VSUBS 0.008029f
C894 B.n637 VSUBS 0.008029f
C895 B.n638 VSUBS 0.008029f
C896 B.n639 VSUBS 0.008029f
C897 B.n640 VSUBS 0.008029f
C898 B.n641 VSUBS 0.008029f
C899 B.n642 VSUBS 0.008029f
C900 B.n643 VSUBS 0.008029f
C901 B.n644 VSUBS 0.008029f
C902 B.n645 VSUBS 0.008029f
C903 B.n646 VSUBS 0.008029f
C904 B.n647 VSUBS 0.008029f
C905 B.n648 VSUBS 0.008029f
C906 B.n649 VSUBS 0.008029f
C907 B.n650 VSUBS 0.008029f
C908 B.n651 VSUBS 0.008029f
C909 B.n652 VSUBS 0.008029f
C910 B.n653 VSUBS 0.008029f
C911 B.n654 VSUBS 0.008029f
C912 B.n655 VSUBS 0.008029f
C913 B.n656 VSUBS 0.008029f
C914 B.n657 VSUBS 0.008029f
C915 B.n658 VSUBS 0.008029f
C916 B.n659 VSUBS 0.008029f
C917 B.n660 VSUBS 0.008029f
C918 B.n661 VSUBS 0.008029f
C919 B.n662 VSUBS 0.008029f
C920 B.n663 VSUBS 0.008029f
C921 B.n664 VSUBS 0.008029f
C922 B.n665 VSUBS 0.008029f
C923 B.n666 VSUBS 0.008029f
C924 B.n667 VSUBS 0.008029f
C925 B.n668 VSUBS 0.008029f
C926 B.n669 VSUBS 0.008029f
C927 B.n670 VSUBS 0.008029f
C928 B.n671 VSUBS 0.008029f
C929 B.n672 VSUBS 0.008029f
C930 B.n673 VSUBS 0.008029f
C931 B.n674 VSUBS 0.008029f
C932 B.n675 VSUBS 0.008029f
C933 B.n676 VSUBS 0.008029f
C934 B.n677 VSUBS 0.008029f
C935 B.n678 VSUBS 0.008029f
C936 B.n679 VSUBS 0.010477f
C937 B.n680 VSUBS 0.01116f
C938 B.n681 VSUBS 0.022194f
C939 VDD2.n0 VSUBS 0.03049f
C940 VDD2.n1 VSUBS 0.027747f
C941 VDD2.n2 VSUBS 0.01491f
C942 VDD2.n3 VSUBS 0.035242f
C943 VDD2.n4 VSUBS 0.015787f
C944 VDD2.n5 VSUBS 0.027747f
C945 VDD2.n6 VSUBS 0.01491f
C946 VDD2.n7 VSUBS 0.035242f
C947 VDD2.n8 VSUBS 0.015787f
C948 VDD2.n9 VSUBS 0.027747f
C949 VDD2.n10 VSUBS 0.01491f
C950 VDD2.n11 VSUBS 0.035242f
C951 VDD2.n12 VSUBS 0.015349f
C952 VDD2.n13 VSUBS 0.027747f
C953 VDD2.n14 VSUBS 0.015787f
C954 VDD2.n15 VSUBS 0.035242f
C955 VDD2.n16 VSUBS 0.015787f
C956 VDD2.n17 VSUBS 0.027747f
C957 VDD2.n18 VSUBS 0.01491f
C958 VDD2.n19 VSUBS 0.035242f
C959 VDD2.n20 VSUBS 0.015787f
C960 VDD2.n21 VSUBS 1.54445f
C961 VDD2.n22 VSUBS 0.01491f
C962 VDD2.t0 VSUBS 0.076079f
C963 VDD2.n23 VSUBS 0.237215f
C964 VDD2.n24 VSUBS 0.026511f
C965 VDD2.n25 VSUBS 0.026431f
C966 VDD2.n26 VSUBS 0.035242f
C967 VDD2.n27 VSUBS 0.015787f
C968 VDD2.n28 VSUBS 0.01491f
C969 VDD2.n29 VSUBS 0.027747f
C970 VDD2.n30 VSUBS 0.027747f
C971 VDD2.n31 VSUBS 0.01491f
C972 VDD2.n32 VSUBS 0.015787f
C973 VDD2.n33 VSUBS 0.035242f
C974 VDD2.n34 VSUBS 0.035242f
C975 VDD2.n35 VSUBS 0.015787f
C976 VDD2.n36 VSUBS 0.01491f
C977 VDD2.n37 VSUBS 0.027747f
C978 VDD2.n38 VSUBS 0.027747f
C979 VDD2.n39 VSUBS 0.01491f
C980 VDD2.n40 VSUBS 0.01491f
C981 VDD2.n41 VSUBS 0.015787f
C982 VDD2.n42 VSUBS 0.035242f
C983 VDD2.n43 VSUBS 0.035242f
C984 VDD2.n44 VSUBS 0.035242f
C985 VDD2.n45 VSUBS 0.015349f
C986 VDD2.n46 VSUBS 0.01491f
C987 VDD2.n47 VSUBS 0.027747f
C988 VDD2.n48 VSUBS 0.027747f
C989 VDD2.n49 VSUBS 0.01491f
C990 VDD2.n50 VSUBS 0.015787f
C991 VDD2.n51 VSUBS 0.035242f
C992 VDD2.n52 VSUBS 0.035242f
C993 VDD2.n53 VSUBS 0.015787f
C994 VDD2.n54 VSUBS 0.01491f
C995 VDD2.n55 VSUBS 0.027747f
C996 VDD2.n56 VSUBS 0.027747f
C997 VDD2.n57 VSUBS 0.01491f
C998 VDD2.n58 VSUBS 0.015787f
C999 VDD2.n59 VSUBS 0.035242f
C1000 VDD2.n60 VSUBS 0.035242f
C1001 VDD2.n61 VSUBS 0.015787f
C1002 VDD2.n62 VSUBS 0.01491f
C1003 VDD2.n63 VSUBS 0.027747f
C1004 VDD2.n64 VSUBS 0.027747f
C1005 VDD2.n65 VSUBS 0.01491f
C1006 VDD2.n66 VSUBS 0.015787f
C1007 VDD2.n67 VSUBS 0.035242f
C1008 VDD2.n68 VSUBS 0.085322f
C1009 VDD2.n69 VSUBS 0.015787f
C1010 VDD2.n70 VSUBS 0.01491f
C1011 VDD2.n71 VSUBS 0.061482f
C1012 VDD2.n72 VSUBS 0.065872f
C1013 VDD2.t4 VSUBS 0.295789f
C1014 VDD2.t8 VSUBS 0.295789f
C1015 VDD2.n73 VSUBS 2.34584f
C1016 VDD2.n74 VSUBS 0.824309f
C1017 VDD2.t7 VSUBS 0.295789f
C1018 VDD2.t3 VSUBS 0.295789f
C1019 VDD2.n75 VSUBS 2.35438f
C1020 VDD2.n76 VSUBS 2.72865f
C1021 VDD2.n77 VSUBS 0.03049f
C1022 VDD2.n78 VSUBS 0.027747f
C1023 VDD2.n79 VSUBS 0.01491f
C1024 VDD2.n80 VSUBS 0.035242f
C1025 VDD2.n81 VSUBS 0.015787f
C1026 VDD2.n82 VSUBS 0.027747f
C1027 VDD2.n83 VSUBS 0.01491f
C1028 VDD2.n84 VSUBS 0.035242f
C1029 VDD2.n85 VSUBS 0.015787f
C1030 VDD2.n86 VSUBS 0.027747f
C1031 VDD2.n87 VSUBS 0.01491f
C1032 VDD2.n88 VSUBS 0.035242f
C1033 VDD2.n89 VSUBS 0.015349f
C1034 VDD2.n90 VSUBS 0.027747f
C1035 VDD2.n91 VSUBS 0.015349f
C1036 VDD2.n92 VSUBS 0.01491f
C1037 VDD2.n93 VSUBS 0.035242f
C1038 VDD2.n94 VSUBS 0.035242f
C1039 VDD2.n95 VSUBS 0.015787f
C1040 VDD2.n96 VSUBS 0.027747f
C1041 VDD2.n97 VSUBS 0.01491f
C1042 VDD2.n98 VSUBS 0.035242f
C1043 VDD2.n99 VSUBS 0.015787f
C1044 VDD2.n100 VSUBS 1.54445f
C1045 VDD2.n101 VSUBS 0.01491f
C1046 VDD2.t1 VSUBS 0.076079f
C1047 VDD2.n102 VSUBS 0.237215f
C1048 VDD2.n103 VSUBS 0.026511f
C1049 VDD2.n104 VSUBS 0.026431f
C1050 VDD2.n105 VSUBS 0.035242f
C1051 VDD2.n106 VSUBS 0.015787f
C1052 VDD2.n107 VSUBS 0.01491f
C1053 VDD2.n108 VSUBS 0.027747f
C1054 VDD2.n109 VSUBS 0.027747f
C1055 VDD2.n110 VSUBS 0.01491f
C1056 VDD2.n111 VSUBS 0.015787f
C1057 VDD2.n112 VSUBS 0.035242f
C1058 VDD2.n113 VSUBS 0.035242f
C1059 VDD2.n114 VSUBS 0.015787f
C1060 VDD2.n115 VSUBS 0.01491f
C1061 VDD2.n116 VSUBS 0.027747f
C1062 VDD2.n117 VSUBS 0.027747f
C1063 VDD2.n118 VSUBS 0.01491f
C1064 VDD2.n119 VSUBS 0.015787f
C1065 VDD2.n120 VSUBS 0.035242f
C1066 VDD2.n121 VSUBS 0.035242f
C1067 VDD2.n122 VSUBS 0.015787f
C1068 VDD2.n123 VSUBS 0.01491f
C1069 VDD2.n124 VSUBS 0.027747f
C1070 VDD2.n125 VSUBS 0.027747f
C1071 VDD2.n126 VSUBS 0.01491f
C1072 VDD2.n127 VSUBS 0.015787f
C1073 VDD2.n128 VSUBS 0.035242f
C1074 VDD2.n129 VSUBS 0.035242f
C1075 VDD2.n130 VSUBS 0.015787f
C1076 VDD2.n131 VSUBS 0.01491f
C1077 VDD2.n132 VSUBS 0.027747f
C1078 VDD2.n133 VSUBS 0.027747f
C1079 VDD2.n134 VSUBS 0.01491f
C1080 VDD2.n135 VSUBS 0.015787f
C1081 VDD2.n136 VSUBS 0.035242f
C1082 VDD2.n137 VSUBS 0.035242f
C1083 VDD2.n138 VSUBS 0.015787f
C1084 VDD2.n139 VSUBS 0.01491f
C1085 VDD2.n140 VSUBS 0.027747f
C1086 VDD2.n141 VSUBS 0.027747f
C1087 VDD2.n142 VSUBS 0.01491f
C1088 VDD2.n143 VSUBS 0.015787f
C1089 VDD2.n144 VSUBS 0.035242f
C1090 VDD2.n145 VSUBS 0.085322f
C1091 VDD2.n146 VSUBS 0.015787f
C1092 VDD2.n147 VSUBS 0.01491f
C1093 VDD2.n148 VSUBS 0.061482f
C1094 VDD2.n149 VSUBS 0.062006f
C1095 VDD2.n150 VSUBS 2.66777f
C1096 VDD2.t2 VSUBS 0.295789f
C1097 VDD2.t9 VSUBS 0.295789f
C1098 VDD2.n151 VSUBS 2.34585f
C1099 VDD2.n152 VSUBS 0.677384f
C1100 VDD2.t6 VSUBS 0.295789f
C1101 VDD2.t5 VSUBS 0.295789f
C1102 VDD2.n153 VSUBS 2.35434f
C1103 VTAIL.t12 VSUBS 0.298628f
C1104 VTAIL.t18 VSUBS 0.298628f
C1105 VTAIL.n0 VSUBS 2.2026f
C1106 VTAIL.n1 VSUBS 0.853985f
C1107 VTAIL.n2 VSUBS 0.030782f
C1108 VTAIL.n3 VSUBS 0.028013f
C1109 VTAIL.n4 VSUBS 0.015053f
C1110 VTAIL.n5 VSUBS 0.03558f
C1111 VTAIL.n6 VSUBS 0.015939f
C1112 VTAIL.n7 VSUBS 0.028013f
C1113 VTAIL.n8 VSUBS 0.015053f
C1114 VTAIL.n9 VSUBS 0.03558f
C1115 VTAIL.n10 VSUBS 0.015939f
C1116 VTAIL.n11 VSUBS 0.028013f
C1117 VTAIL.n12 VSUBS 0.015053f
C1118 VTAIL.n13 VSUBS 0.03558f
C1119 VTAIL.n14 VSUBS 0.015496f
C1120 VTAIL.n15 VSUBS 0.028013f
C1121 VTAIL.n16 VSUBS 0.015939f
C1122 VTAIL.n17 VSUBS 0.03558f
C1123 VTAIL.n18 VSUBS 0.015939f
C1124 VTAIL.n19 VSUBS 0.028013f
C1125 VTAIL.n20 VSUBS 0.015053f
C1126 VTAIL.n21 VSUBS 0.03558f
C1127 VTAIL.n22 VSUBS 0.015939f
C1128 VTAIL.n23 VSUBS 1.55928f
C1129 VTAIL.n24 VSUBS 0.015053f
C1130 VTAIL.t9 VSUBS 0.076809f
C1131 VTAIL.n25 VSUBS 0.239492f
C1132 VTAIL.n26 VSUBS 0.026765f
C1133 VTAIL.n27 VSUBS 0.026685f
C1134 VTAIL.n28 VSUBS 0.03558f
C1135 VTAIL.n29 VSUBS 0.015939f
C1136 VTAIL.n30 VSUBS 0.015053f
C1137 VTAIL.n31 VSUBS 0.028013f
C1138 VTAIL.n32 VSUBS 0.028013f
C1139 VTAIL.n33 VSUBS 0.015053f
C1140 VTAIL.n34 VSUBS 0.015939f
C1141 VTAIL.n35 VSUBS 0.03558f
C1142 VTAIL.n36 VSUBS 0.03558f
C1143 VTAIL.n37 VSUBS 0.015939f
C1144 VTAIL.n38 VSUBS 0.015053f
C1145 VTAIL.n39 VSUBS 0.028013f
C1146 VTAIL.n40 VSUBS 0.028013f
C1147 VTAIL.n41 VSUBS 0.015053f
C1148 VTAIL.n42 VSUBS 0.015053f
C1149 VTAIL.n43 VSUBS 0.015939f
C1150 VTAIL.n44 VSUBS 0.03558f
C1151 VTAIL.n45 VSUBS 0.03558f
C1152 VTAIL.n46 VSUBS 0.03558f
C1153 VTAIL.n47 VSUBS 0.015496f
C1154 VTAIL.n48 VSUBS 0.015053f
C1155 VTAIL.n49 VSUBS 0.028013f
C1156 VTAIL.n50 VSUBS 0.028013f
C1157 VTAIL.n51 VSUBS 0.015053f
C1158 VTAIL.n52 VSUBS 0.015939f
C1159 VTAIL.n53 VSUBS 0.03558f
C1160 VTAIL.n54 VSUBS 0.03558f
C1161 VTAIL.n55 VSUBS 0.015939f
C1162 VTAIL.n56 VSUBS 0.015053f
C1163 VTAIL.n57 VSUBS 0.028013f
C1164 VTAIL.n58 VSUBS 0.028013f
C1165 VTAIL.n59 VSUBS 0.015053f
C1166 VTAIL.n60 VSUBS 0.015939f
C1167 VTAIL.n61 VSUBS 0.03558f
C1168 VTAIL.n62 VSUBS 0.03558f
C1169 VTAIL.n63 VSUBS 0.015939f
C1170 VTAIL.n64 VSUBS 0.015053f
C1171 VTAIL.n65 VSUBS 0.028013f
C1172 VTAIL.n66 VSUBS 0.028013f
C1173 VTAIL.n67 VSUBS 0.015053f
C1174 VTAIL.n68 VSUBS 0.015939f
C1175 VTAIL.n69 VSUBS 0.03558f
C1176 VTAIL.n70 VSUBS 0.086141f
C1177 VTAIL.n71 VSUBS 0.015939f
C1178 VTAIL.n72 VSUBS 0.015053f
C1179 VTAIL.n73 VSUBS 0.062073f
C1180 VTAIL.n74 VSUBS 0.043236f
C1181 VTAIL.n75 VSUBS 0.225901f
C1182 VTAIL.t8 VSUBS 0.298628f
C1183 VTAIL.t7 VSUBS 0.298628f
C1184 VTAIL.n76 VSUBS 2.2026f
C1185 VTAIL.n77 VSUBS 0.886862f
C1186 VTAIL.t4 VSUBS 0.298628f
C1187 VTAIL.t1 VSUBS 0.298628f
C1188 VTAIL.n78 VSUBS 2.2026f
C1189 VTAIL.n79 VSUBS 2.4245f
C1190 VTAIL.t15 VSUBS 0.298628f
C1191 VTAIL.t16 VSUBS 0.298628f
C1192 VTAIL.n80 VSUBS 2.20262f
C1193 VTAIL.n81 VSUBS 2.42448f
C1194 VTAIL.t17 VSUBS 0.298628f
C1195 VTAIL.t19 VSUBS 0.298628f
C1196 VTAIL.n82 VSUBS 2.20262f
C1197 VTAIL.n83 VSUBS 0.886847f
C1198 VTAIL.n84 VSUBS 0.030782f
C1199 VTAIL.n85 VSUBS 0.028013f
C1200 VTAIL.n86 VSUBS 0.015053f
C1201 VTAIL.n87 VSUBS 0.03558f
C1202 VTAIL.n88 VSUBS 0.015939f
C1203 VTAIL.n89 VSUBS 0.028013f
C1204 VTAIL.n90 VSUBS 0.015053f
C1205 VTAIL.n91 VSUBS 0.03558f
C1206 VTAIL.n92 VSUBS 0.015939f
C1207 VTAIL.n93 VSUBS 0.028013f
C1208 VTAIL.n94 VSUBS 0.015053f
C1209 VTAIL.n95 VSUBS 0.03558f
C1210 VTAIL.n96 VSUBS 0.015496f
C1211 VTAIL.n97 VSUBS 0.028013f
C1212 VTAIL.n98 VSUBS 0.015496f
C1213 VTAIL.n99 VSUBS 0.015053f
C1214 VTAIL.n100 VSUBS 0.03558f
C1215 VTAIL.n101 VSUBS 0.03558f
C1216 VTAIL.n102 VSUBS 0.015939f
C1217 VTAIL.n103 VSUBS 0.028013f
C1218 VTAIL.n104 VSUBS 0.015053f
C1219 VTAIL.n105 VSUBS 0.03558f
C1220 VTAIL.n106 VSUBS 0.015939f
C1221 VTAIL.n107 VSUBS 1.55928f
C1222 VTAIL.n108 VSUBS 0.015053f
C1223 VTAIL.t11 VSUBS 0.076809f
C1224 VTAIL.n109 VSUBS 0.239492f
C1225 VTAIL.n110 VSUBS 0.026765f
C1226 VTAIL.n111 VSUBS 0.026685f
C1227 VTAIL.n112 VSUBS 0.03558f
C1228 VTAIL.n113 VSUBS 0.015939f
C1229 VTAIL.n114 VSUBS 0.015053f
C1230 VTAIL.n115 VSUBS 0.028013f
C1231 VTAIL.n116 VSUBS 0.028013f
C1232 VTAIL.n117 VSUBS 0.015053f
C1233 VTAIL.n118 VSUBS 0.015939f
C1234 VTAIL.n119 VSUBS 0.03558f
C1235 VTAIL.n120 VSUBS 0.03558f
C1236 VTAIL.n121 VSUBS 0.015939f
C1237 VTAIL.n122 VSUBS 0.015053f
C1238 VTAIL.n123 VSUBS 0.028013f
C1239 VTAIL.n124 VSUBS 0.028013f
C1240 VTAIL.n125 VSUBS 0.015053f
C1241 VTAIL.n126 VSUBS 0.015939f
C1242 VTAIL.n127 VSUBS 0.03558f
C1243 VTAIL.n128 VSUBS 0.03558f
C1244 VTAIL.n129 VSUBS 0.015939f
C1245 VTAIL.n130 VSUBS 0.015053f
C1246 VTAIL.n131 VSUBS 0.028013f
C1247 VTAIL.n132 VSUBS 0.028013f
C1248 VTAIL.n133 VSUBS 0.015053f
C1249 VTAIL.n134 VSUBS 0.015939f
C1250 VTAIL.n135 VSUBS 0.03558f
C1251 VTAIL.n136 VSUBS 0.03558f
C1252 VTAIL.n137 VSUBS 0.015939f
C1253 VTAIL.n138 VSUBS 0.015053f
C1254 VTAIL.n139 VSUBS 0.028013f
C1255 VTAIL.n140 VSUBS 0.028013f
C1256 VTAIL.n141 VSUBS 0.015053f
C1257 VTAIL.n142 VSUBS 0.015939f
C1258 VTAIL.n143 VSUBS 0.03558f
C1259 VTAIL.n144 VSUBS 0.03558f
C1260 VTAIL.n145 VSUBS 0.015939f
C1261 VTAIL.n146 VSUBS 0.015053f
C1262 VTAIL.n147 VSUBS 0.028013f
C1263 VTAIL.n148 VSUBS 0.028013f
C1264 VTAIL.n149 VSUBS 0.015053f
C1265 VTAIL.n150 VSUBS 0.015939f
C1266 VTAIL.n151 VSUBS 0.03558f
C1267 VTAIL.n152 VSUBS 0.086141f
C1268 VTAIL.n153 VSUBS 0.015939f
C1269 VTAIL.n154 VSUBS 0.015053f
C1270 VTAIL.n155 VSUBS 0.062073f
C1271 VTAIL.n156 VSUBS 0.043236f
C1272 VTAIL.n157 VSUBS 0.225901f
C1273 VTAIL.t0 VSUBS 0.298628f
C1274 VTAIL.t5 VSUBS 0.298628f
C1275 VTAIL.n158 VSUBS 2.20262f
C1276 VTAIL.n159 VSUBS 0.875564f
C1277 VTAIL.t2 VSUBS 0.298628f
C1278 VTAIL.t3 VSUBS 0.298628f
C1279 VTAIL.n160 VSUBS 2.20262f
C1280 VTAIL.n161 VSUBS 0.886847f
C1281 VTAIL.n162 VSUBS 0.030782f
C1282 VTAIL.n163 VSUBS 0.028013f
C1283 VTAIL.n164 VSUBS 0.015053f
C1284 VTAIL.n165 VSUBS 0.03558f
C1285 VTAIL.n166 VSUBS 0.015939f
C1286 VTAIL.n167 VSUBS 0.028013f
C1287 VTAIL.n168 VSUBS 0.015053f
C1288 VTAIL.n169 VSUBS 0.03558f
C1289 VTAIL.n170 VSUBS 0.015939f
C1290 VTAIL.n171 VSUBS 0.028013f
C1291 VTAIL.n172 VSUBS 0.015053f
C1292 VTAIL.n173 VSUBS 0.03558f
C1293 VTAIL.n174 VSUBS 0.015496f
C1294 VTAIL.n175 VSUBS 0.028013f
C1295 VTAIL.n176 VSUBS 0.015496f
C1296 VTAIL.n177 VSUBS 0.015053f
C1297 VTAIL.n178 VSUBS 0.03558f
C1298 VTAIL.n179 VSUBS 0.03558f
C1299 VTAIL.n180 VSUBS 0.015939f
C1300 VTAIL.n181 VSUBS 0.028013f
C1301 VTAIL.n182 VSUBS 0.015053f
C1302 VTAIL.n183 VSUBS 0.03558f
C1303 VTAIL.n184 VSUBS 0.015939f
C1304 VTAIL.n185 VSUBS 1.55928f
C1305 VTAIL.n186 VSUBS 0.015053f
C1306 VTAIL.t6 VSUBS 0.076809f
C1307 VTAIL.n187 VSUBS 0.239492f
C1308 VTAIL.n188 VSUBS 0.026765f
C1309 VTAIL.n189 VSUBS 0.026685f
C1310 VTAIL.n190 VSUBS 0.03558f
C1311 VTAIL.n191 VSUBS 0.015939f
C1312 VTAIL.n192 VSUBS 0.015053f
C1313 VTAIL.n193 VSUBS 0.028013f
C1314 VTAIL.n194 VSUBS 0.028013f
C1315 VTAIL.n195 VSUBS 0.015053f
C1316 VTAIL.n196 VSUBS 0.015939f
C1317 VTAIL.n197 VSUBS 0.03558f
C1318 VTAIL.n198 VSUBS 0.03558f
C1319 VTAIL.n199 VSUBS 0.015939f
C1320 VTAIL.n200 VSUBS 0.015053f
C1321 VTAIL.n201 VSUBS 0.028013f
C1322 VTAIL.n202 VSUBS 0.028013f
C1323 VTAIL.n203 VSUBS 0.015053f
C1324 VTAIL.n204 VSUBS 0.015939f
C1325 VTAIL.n205 VSUBS 0.03558f
C1326 VTAIL.n206 VSUBS 0.03558f
C1327 VTAIL.n207 VSUBS 0.015939f
C1328 VTAIL.n208 VSUBS 0.015053f
C1329 VTAIL.n209 VSUBS 0.028013f
C1330 VTAIL.n210 VSUBS 0.028013f
C1331 VTAIL.n211 VSUBS 0.015053f
C1332 VTAIL.n212 VSUBS 0.015939f
C1333 VTAIL.n213 VSUBS 0.03558f
C1334 VTAIL.n214 VSUBS 0.03558f
C1335 VTAIL.n215 VSUBS 0.015939f
C1336 VTAIL.n216 VSUBS 0.015053f
C1337 VTAIL.n217 VSUBS 0.028013f
C1338 VTAIL.n218 VSUBS 0.028013f
C1339 VTAIL.n219 VSUBS 0.015053f
C1340 VTAIL.n220 VSUBS 0.015939f
C1341 VTAIL.n221 VSUBS 0.03558f
C1342 VTAIL.n222 VSUBS 0.03558f
C1343 VTAIL.n223 VSUBS 0.015939f
C1344 VTAIL.n224 VSUBS 0.015053f
C1345 VTAIL.n225 VSUBS 0.028013f
C1346 VTAIL.n226 VSUBS 0.028013f
C1347 VTAIL.n227 VSUBS 0.015053f
C1348 VTAIL.n228 VSUBS 0.015939f
C1349 VTAIL.n229 VSUBS 0.03558f
C1350 VTAIL.n230 VSUBS 0.086141f
C1351 VTAIL.n231 VSUBS 0.015939f
C1352 VTAIL.n232 VSUBS 0.015053f
C1353 VTAIL.n233 VSUBS 0.062073f
C1354 VTAIL.n234 VSUBS 0.043236f
C1355 VTAIL.n235 VSUBS 1.66743f
C1356 VTAIL.n236 VSUBS 0.030782f
C1357 VTAIL.n237 VSUBS 0.028013f
C1358 VTAIL.n238 VSUBS 0.015053f
C1359 VTAIL.n239 VSUBS 0.03558f
C1360 VTAIL.n240 VSUBS 0.015939f
C1361 VTAIL.n241 VSUBS 0.028013f
C1362 VTAIL.n242 VSUBS 0.015053f
C1363 VTAIL.n243 VSUBS 0.03558f
C1364 VTAIL.n244 VSUBS 0.015939f
C1365 VTAIL.n245 VSUBS 0.028013f
C1366 VTAIL.n246 VSUBS 0.015053f
C1367 VTAIL.n247 VSUBS 0.03558f
C1368 VTAIL.n248 VSUBS 0.015496f
C1369 VTAIL.n249 VSUBS 0.028013f
C1370 VTAIL.n250 VSUBS 0.015939f
C1371 VTAIL.n251 VSUBS 0.03558f
C1372 VTAIL.n252 VSUBS 0.015939f
C1373 VTAIL.n253 VSUBS 0.028013f
C1374 VTAIL.n254 VSUBS 0.015053f
C1375 VTAIL.n255 VSUBS 0.03558f
C1376 VTAIL.n256 VSUBS 0.015939f
C1377 VTAIL.n257 VSUBS 1.55928f
C1378 VTAIL.n258 VSUBS 0.015053f
C1379 VTAIL.t13 VSUBS 0.076809f
C1380 VTAIL.n259 VSUBS 0.239492f
C1381 VTAIL.n260 VSUBS 0.026765f
C1382 VTAIL.n261 VSUBS 0.026685f
C1383 VTAIL.n262 VSUBS 0.03558f
C1384 VTAIL.n263 VSUBS 0.015939f
C1385 VTAIL.n264 VSUBS 0.015053f
C1386 VTAIL.n265 VSUBS 0.028013f
C1387 VTAIL.n266 VSUBS 0.028013f
C1388 VTAIL.n267 VSUBS 0.015053f
C1389 VTAIL.n268 VSUBS 0.015939f
C1390 VTAIL.n269 VSUBS 0.03558f
C1391 VTAIL.n270 VSUBS 0.03558f
C1392 VTAIL.n271 VSUBS 0.015939f
C1393 VTAIL.n272 VSUBS 0.015053f
C1394 VTAIL.n273 VSUBS 0.028013f
C1395 VTAIL.n274 VSUBS 0.028013f
C1396 VTAIL.n275 VSUBS 0.015053f
C1397 VTAIL.n276 VSUBS 0.015053f
C1398 VTAIL.n277 VSUBS 0.015939f
C1399 VTAIL.n278 VSUBS 0.03558f
C1400 VTAIL.n279 VSUBS 0.03558f
C1401 VTAIL.n280 VSUBS 0.03558f
C1402 VTAIL.n281 VSUBS 0.015496f
C1403 VTAIL.n282 VSUBS 0.015053f
C1404 VTAIL.n283 VSUBS 0.028013f
C1405 VTAIL.n284 VSUBS 0.028013f
C1406 VTAIL.n285 VSUBS 0.015053f
C1407 VTAIL.n286 VSUBS 0.015939f
C1408 VTAIL.n287 VSUBS 0.03558f
C1409 VTAIL.n288 VSUBS 0.03558f
C1410 VTAIL.n289 VSUBS 0.015939f
C1411 VTAIL.n290 VSUBS 0.015053f
C1412 VTAIL.n291 VSUBS 0.028013f
C1413 VTAIL.n292 VSUBS 0.028013f
C1414 VTAIL.n293 VSUBS 0.015053f
C1415 VTAIL.n294 VSUBS 0.015939f
C1416 VTAIL.n295 VSUBS 0.03558f
C1417 VTAIL.n296 VSUBS 0.03558f
C1418 VTAIL.n297 VSUBS 0.015939f
C1419 VTAIL.n298 VSUBS 0.015053f
C1420 VTAIL.n299 VSUBS 0.028013f
C1421 VTAIL.n300 VSUBS 0.028013f
C1422 VTAIL.n301 VSUBS 0.015053f
C1423 VTAIL.n302 VSUBS 0.015939f
C1424 VTAIL.n303 VSUBS 0.03558f
C1425 VTAIL.n304 VSUBS 0.086141f
C1426 VTAIL.n305 VSUBS 0.015939f
C1427 VTAIL.n306 VSUBS 0.015053f
C1428 VTAIL.n307 VSUBS 0.062073f
C1429 VTAIL.n308 VSUBS 0.043236f
C1430 VTAIL.n309 VSUBS 1.66743f
C1431 VTAIL.t14 VSUBS 0.298628f
C1432 VTAIL.t10 VSUBS 0.298628f
C1433 VTAIL.n310 VSUBS 2.2026f
C1434 VTAIL.n311 VSUBS 0.801071f
C1435 VN.n0 VSUBS 0.058108f
C1436 VN.t2 VSUBS 1.6859f
C1437 VN.n1 VSUBS 0.037259f
C1438 VN.n2 VSUBS 0.043547f
C1439 VN.t1 VSUBS 1.6859f
C1440 VN.n3 VSUBS 0.058343f
C1441 VN.t9 VSUBS 1.78472f
C1442 VN.t5 VSUBS 1.6859f
C1443 VN.n4 VSUBS 0.654708f
C1444 VN.n5 VSUBS 0.683449f
C1445 VN.n6 VSUBS 0.188554f
C1446 VN.n7 VSUBS 0.043547f
C1447 VN.n8 VSUBS 0.037259f
C1448 VN.n9 VSUBS 0.063013f
C1449 VN.n10 VSUBS 0.616273f
C1450 VN.n11 VSUBS 0.063013f
C1451 VN.n12 VSUBS 0.043547f
C1452 VN.n13 VSUBS 0.043547f
C1453 VN.n14 VSUBS 0.043547f
C1454 VN.n15 VSUBS 0.058343f
C1455 VN.n16 VSUBS 0.616273f
C1456 VN.n17 VSUBS 0.061478f
C1457 VN.t6 VSUBS 1.75595f
C1458 VN.n18 VSUBS 0.688241f
C1459 VN.n19 VSUBS 0.040783f
C1460 VN.n20 VSUBS 0.058108f
C1461 VN.t7 VSUBS 1.6859f
C1462 VN.n21 VSUBS 0.037259f
C1463 VN.n22 VSUBS 0.043547f
C1464 VN.t0 VSUBS 1.6859f
C1465 VN.n23 VSUBS 0.058343f
C1466 VN.t4 VSUBS 1.78472f
C1467 VN.t3 VSUBS 1.6859f
C1468 VN.n24 VSUBS 0.654708f
C1469 VN.n25 VSUBS 0.683449f
C1470 VN.n26 VSUBS 0.188554f
C1471 VN.n27 VSUBS 0.043547f
C1472 VN.n28 VSUBS 0.037259f
C1473 VN.n29 VSUBS 0.063013f
C1474 VN.n30 VSUBS 0.616273f
C1475 VN.n31 VSUBS 0.063013f
C1476 VN.n32 VSUBS 0.043547f
C1477 VN.n33 VSUBS 0.043547f
C1478 VN.n34 VSUBS 0.043547f
C1479 VN.n35 VSUBS 0.058343f
C1480 VN.n36 VSUBS 0.616273f
C1481 VN.n37 VSUBS 0.061478f
C1482 VN.t8 VSUBS 1.75595f
C1483 VN.n38 VSUBS 0.688241f
C1484 VN.n39 VSUBS 2.12605f
.ends

