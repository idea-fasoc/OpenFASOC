* NGSPICE file created from diff_pair_sample_0198.ext - technology: sky130A

.subckt diff_pair_sample_0198 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t1 VP.t0 VTAIL.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=4.8555 pd=25.68 as=4.8555 ps=25.68 w=12.45 l=3.86
X1 B.t15 B.t13 B.t14 B.t7 sky130_fd_pr__nfet_01v8 ad=4.8555 pd=25.68 as=0 ps=0 w=12.45 l=3.86
X2 VDD2.t1 VN.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=4.8555 pd=25.68 as=4.8555 ps=25.68 w=12.45 l=3.86
X3 B.t12 B.t10 B.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=4.8555 pd=25.68 as=0 ps=0 w=12.45 l=3.86
X4 VDD2.t0 VN.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=4.8555 pd=25.68 as=4.8555 ps=25.68 w=12.45 l=3.86
X5 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=4.8555 pd=25.68 as=0 ps=0 w=12.45 l=3.86
X6 VDD1.t0 VP.t1 VTAIL.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=4.8555 pd=25.68 as=4.8555 ps=25.68 w=12.45 l=3.86
X7 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=4.8555 pd=25.68 as=0 ps=0 w=12.45 l=3.86
R0 VP.n0 VP.t0 161.108
R1 VP.n0 VP.t1 112.769
R2 VP VP.n0 0.621237
R3 VTAIL.n1 VTAIL.t0 46.1172
R4 VTAIL.n3 VTAIL.t1 46.1171
R5 VTAIL.n0 VTAIL.t3 46.1171
R6 VTAIL.n2 VTAIL.t2 46.1171
R7 VTAIL.n1 VTAIL.n0 30.3238
R8 VTAIL.n3 VTAIL.n2 26.7117
R9 VTAIL.n2 VTAIL.n1 2.27636
R10 VTAIL VTAIL.n0 1.43153
R11 VTAIL VTAIL.n3 0.845328
R12 VDD1 VDD1.t0 105.841
R13 VDD1 VDD1.t1 63.7571
R14 B.n747 B.n746 585
R15 B.n748 B.n747 585
R16 B.n301 B.n110 585
R17 B.n300 B.n299 585
R18 B.n298 B.n297 585
R19 B.n296 B.n295 585
R20 B.n294 B.n293 585
R21 B.n292 B.n291 585
R22 B.n290 B.n289 585
R23 B.n288 B.n287 585
R24 B.n286 B.n285 585
R25 B.n284 B.n283 585
R26 B.n282 B.n281 585
R27 B.n280 B.n279 585
R28 B.n278 B.n277 585
R29 B.n276 B.n275 585
R30 B.n274 B.n273 585
R31 B.n272 B.n271 585
R32 B.n270 B.n269 585
R33 B.n268 B.n267 585
R34 B.n266 B.n265 585
R35 B.n264 B.n263 585
R36 B.n262 B.n261 585
R37 B.n260 B.n259 585
R38 B.n258 B.n257 585
R39 B.n256 B.n255 585
R40 B.n254 B.n253 585
R41 B.n252 B.n251 585
R42 B.n250 B.n249 585
R43 B.n248 B.n247 585
R44 B.n246 B.n245 585
R45 B.n244 B.n243 585
R46 B.n242 B.n241 585
R47 B.n240 B.n239 585
R48 B.n238 B.n237 585
R49 B.n236 B.n235 585
R50 B.n234 B.n233 585
R51 B.n232 B.n231 585
R52 B.n230 B.n229 585
R53 B.n228 B.n227 585
R54 B.n226 B.n225 585
R55 B.n224 B.n223 585
R56 B.n222 B.n221 585
R57 B.n220 B.n219 585
R58 B.n218 B.n217 585
R59 B.n216 B.n215 585
R60 B.n214 B.n213 585
R61 B.n212 B.n211 585
R62 B.n210 B.n209 585
R63 B.n208 B.n207 585
R64 B.n206 B.n205 585
R65 B.n204 B.n203 585
R66 B.n202 B.n201 585
R67 B.n199 B.n198 585
R68 B.n197 B.n196 585
R69 B.n195 B.n194 585
R70 B.n193 B.n192 585
R71 B.n191 B.n190 585
R72 B.n189 B.n188 585
R73 B.n187 B.n186 585
R74 B.n185 B.n184 585
R75 B.n183 B.n182 585
R76 B.n181 B.n180 585
R77 B.n179 B.n178 585
R78 B.n177 B.n176 585
R79 B.n175 B.n174 585
R80 B.n173 B.n172 585
R81 B.n171 B.n170 585
R82 B.n169 B.n168 585
R83 B.n167 B.n166 585
R84 B.n165 B.n164 585
R85 B.n163 B.n162 585
R86 B.n161 B.n160 585
R87 B.n159 B.n158 585
R88 B.n157 B.n156 585
R89 B.n155 B.n154 585
R90 B.n153 B.n152 585
R91 B.n151 B.n150 585
R92 B.n149 B.n148 585
R93 B.n147 B.n146 585
R94 B.n145 B.n144 585
R95 B.n143 B.n142 585
R96 B.n141 B.n140 585
R97 B.n139 B.n138 585
R98 B.n137 B.n136 585
R99 B.n135 B.n134 585
R100 B.n133 B.n132 585
R101 B.n131 B.n130 585
R102 B.n129 B.n128 585
R103 B.n127 B.n126 585
R104 B.n125 B.n124 585
R105 B.n123 B.n122 585
R106 B.n121 B.n120 585
R107 B.n119 B.n118 585
R108 B.n117 B.n116 585
R109 B.n61 B.n60 585
R110 B.n745 B.n62 585
R111 B.n749 B.n62 585
R112 B.n744 B.n743 585
R113 B.n743 B.n58 585
R114 B.n742 B.n57 585
R115 B.n755 B.n57 585
R116 B.n741 B.n56 585
R117 B.n756 B.n56 585
R118 B.n740 B.n55 585
R119 B.n757 B.n55 585
R120 B.n739 B.n738 585
R121 B.n738 B.n51 585
R122 B.n737 B.n50 585
R123 B.n763 B.n50 585
R124 B.n736 B.n49 585
R125 B.n764 B.n49 585
R126 B.n735 B.n48 585
R127 B.n765 B.n48 585
R128 B.n734 B.n733 585
R129 B.n733 B.n47 585
R130 B.n732 B.n43 585
R131 B.n771 B.n43 585
R132 B.n731 B.n42 585
R133 B.n772 B.n42 585
R134 B.n730 B.n41 585
R135 B.n773 B.n41 585
R136 B.n729 B.n728 585
R137 B.n728 B.n37 585
R138 B.n727 B.n36 585
R139 B.n779 B.n36 585
R140 B.n726 B.n35 585
R141 B.n780 B.n35 585
R142 B.n725 B.n34 585
R143 B.n781 B.n34 585
R144 B.n724 B.n723 585
R145 B.n723 B.n30 585
R146 B.n722 B.n29 585
R147 B.n787 B.n29 585
R148 B.n721 B.n28 585
R149 B.n788 B.n28 585
R150 B.n720 B.n27 585
R151 B.n789 B.n27 585
R152 B.n719 B.n718 585
R153 B.n718 B.n23 585
R154 B.n717 B.n22 585
R155 B.n795 B.n22 585
R156 B.n716 B.n21 585
R157 B.n796 B.n21 585
R158 B.n715 B.n20 585
R159 B.n797 B.n20 585
R160 B.n714 B.n713 585
R161 B.n713 B.n16 585
R162 B.n712 B.n15 585
R163 B.n803 B.n15 585
R164 B.n711 B.n14 585
R165 B.n804 B.n14 585
R166 B.n710 B.n13 585
R167 B.n805 B.n13 585
R168 B.n709 B.n708 585
R169 B.n708 B.n12 585
R170 B.n707 B.n706 585
R171 B.n707 B.n8 585
R172 B.n705 B.n7 585
R173 B.n812 B.n7 585
R174 B.n704 B.n6 585
R175 B.n813 B.n6 585
R176 B.n703 B.n5 585
R177 B.n814 B.n5 585
R178 B.n702 B.n701 585
R179 B.n701 B.n4 585
R180 B.n700 B.n302 585
R181 B.n700 B.n699 585
R182 B.n690 B.n303 585
R183 B.n304 B.n303 585
R184 B.n692 B.n691 585
R185 B.n693 B.n692 585
R186 B.n689 B.n309 585
R187 B.n309 B.n308 585
R188 B.n688 B.n687 585
R189 B.n687 B.n686 585
R190 B.n311 B.n310 585
R191 B.n312 B.n311 585
R192 B.n679 B.n678 585
R193 B.n680 B.n679 585
R194 B.n677 B.n317 585
R195 B.n317 B.n316 585
R196 B.n676 B.n675 585
R197 B.n675 B.n674 585
R198 B.n319 B.n318 585
R199 B.n320 B.n319 585
R200 B.n667 B.n666 585
R201 B.n668 B.n667 585
R202 B.n665 B.n325 585
R203 B.n325 B.n324 585
R204 B.n664 B.n663 585
R205 B.n663 B.n662 585
R206 B.n327 B.n326 585
R207 B.n328 B.n327 585
R208 B.n655 B.n654 585
R209 B.n656 B.n655 585
R210 B.n653 B.n333 585
R211 B.n333 B.n332 585
R212 B.n652 B.n651 585
R213 B.n651 B.n650 585
R214 B.n335 B.n334 585
R215 B.n336 B.n335 585
R216 B.n643 B.n642 585
R217 B.n644 B.n643 585
R218 B.n641 B.n341 585
R219 B.n341 B.n340 585
R220 B.n640 B.n639 585
R221 B.n639 B.n638 585
R222 B.n343 B.n342 585
R223 B.n631 B.n343 585
R224 B.n630 B.n629 585
R225 B.n632 B.n630 585
R226 B.n628 B.n348 585
R227 B.n348 B.n347 585
R228 B.n627 B.n626 585
R229 B.n626 B.n625 585
R230 B.n350 B.n349 585
R231 B.n351 B.n350 585
R232 B.n618 B.n617 585
R233 B.n619 B.n618 585
R234 B.n616 B.n356 585
R235 B.n356 B.n355 585
R236 B.n615 B.n614 585
R237 B.n614 B.n613 585
R238 B.n358 B.n357 585
R239 B.n359 B.n358 585
R240 B.n606 B.n605 585
R241 B.n607 B.n606 585
R242 B.n362 B.n361 585
R243 B.n415 B.n414 585
R244 B.n416 B.n412 585
R245 B.n412 B.n363 585
R246 B.n418 B.n417 585
R247 B.n420 B.n411 585
R248 B.n423 B.n422 585
R249 B.n424 B.n410 585
R250 B.n426 B.n425 585
R251 B.n428 B.n409 585
R252 B.n431 B.n430 585
R253 B.n432 B.n408 585
R254 B.n434 B.n433 585
R255 B.n436 B.n407 585
R256 B.n439 B.n438 585
R257 B.n440 B.n406 585
R258 B.n442 B.n441 585
R259 B.n444 B.n405 585
R260 B.n447 B.n446 585
R261 B.n448 B.n404 585
R262 B.n450 B.n449 585
R263 B.n452 B.n403 585
R264 B.n455 B.n454 585
R265 B.n456 B.n402 585
R266 B.n458 B.n457 585
R267 B.n460 B.n401 585
R268 B.n463 B.n462 585
R269 B.n464 B.n400 585
R270 B.n466 B.n465 585
R271 B.n468 B.n399 585
R272 B.n471 B.n470 585
R273 B.n472 B.n398 585
R274 B.n474 B.n473 585
R275 B.n476 B.n397 585
R276 B.n479 B.n478 585
R277 B.n480 B.n396 585
R278 B.n482 B.n481 585
R279 B.n484 B.n395 585
R280 B.n487 B.n486 585
R281 B.n488 B.n394 585
R282 B.n490 B.n489 585
R283 B.n492 B.n393 585
R284 B.n495 B.n494 585
R285 B.n496 B.n390 585
R286 B.n499 B.n498 585
R287 B.n501 B.n389 585
R288 B.n504 B.n503 585
R289 B.n505 B.n388 585
R290 B.n507 B.n506 585
R291 B.n509 B.n387 585
R292 B.n512 B.n511 585
R293 B.n513 B.n386 585
R294 B.n518 B.n517 585
R295 B.n520 B.n385 585
R296 B.n523 B.n522 585
R297 B.n524 B.n384 585
R298 B.n526 B.n525 585
R299 B.n528 B.n383 585
R300 B.n531 B.n530 585
R301 B.n532 B.n382 585
R302 B.n534 B.n533 585
R303 B.n536 B.n381 585
R304 B.n539 B.n538 585
R305 B.n540 B.n380 585
R306 B.n542 B.n541 585
R307 B.n544 B.n379 585
R308 B.n547 B.n546 585
R309 B.n548 B.n378 585
R310 B.n550 B.n549 585
R311 B.n552 B.n377 585
R312 B.n555 B.n554 585
R313 B.n556 B.n376 585
R314 B.n558 B.n557 585
R315 B.n560 B.n375 585
R316 B.n563 B.n562 585
R317 B.n564 B.n374 585
R318 B.n566 B.n565 585
R319 B.n568 B.n373 585
R320 B.n571 B.n570 585
R321 B.n572 B.n372 585
R322 B.n574 B.n573 585
R323 B.n576 B.n371 585
R324 B.n579 B.n578 585
R325 B.n580 B.n370 585
R326 B.n582 B.n581 585
R327 B.n584 B.n369 585
R328 B.n587 B.n586 585
R329 B.n588 B.n368 585
R330 B.n590 B.n589 585
R331 B.n592 B.n367 585
R332 B.n595 B.n594 585
R333 B.n596 B.n366 585
R334 B.n598 B.n597 585
R335 B.n600 B.n365 585
R336 B.n603 B.n602 585
R337 B.n604 B.n364 585
R338 B.n609 B.n608 585
R339 B.n608 B.n607 585
R340 B.n610 B.n360 585
R341 B.n360 B.n359 585
R342 B.n612 B.n611 585
R343 B.n613 B.n612 585
R344 B.n354 B.n353 585
R345 B.n355 B.n354 585
R346 B.n621 B.n620 585
R347 B.n620 B.n619 585
R348 B.n622 B.n352 585
R349 B.n352 B.n351 585
R350 B.n624 B.n623 585
R351 B.n625 B.n624 585
R352 B.n346 B.n345 585
R353 B.n347 B.n346 585
R354 B.n634 B.n633 585
R355 B.n633 B.n632 585
R356 B.n635 B.n344 585
R357 B.n631 B.n344 585
R358 B.n637 B.n636 585
R359 B.n638 B.n637 585
R360 B.n339 B.n338 585
R361 B.n340 B.n339 585
R362 B.n646 B.n645 585
R363 B.n645 B.n644 585
R364 B.n647 B.n337 585
R365 B.n337 B.n336 585
R366 B.n649 B.n648 585
R367 B.n650 B.n649 585
R368 B.n331 B.n330 585
R369 B.n332 B.n331 585
R370 B.n658 B.n657 585
R371 B.n657 B.n656 585
R372 B.n659 B.n329 585
R373 B.n329 B.n328 585
R374 B.n661 B.n660 585
R375 B.n662 B.n661 585
R376 B.n323 B.n322 585
R377 B.n324 B.n323 585
R378 B.n670 B.n669 585
R379 B.n669 B.n668 585
R380 B.n671 B.n321 585
R381 B.n321 B.n320 585
R382 B.n673 B.n672 585
R383 B.n674 B.n673 585
R384 B.n315 B.n314 585
R385 B.n316 B.n315 585
R386 B.n682 B.n681 585
R387 B.n681 B.n680 585
R388 B.n683 B.n313 585
R389 B.n313 B.n312 585
R390 B.n685 B.n684 585
R391 B.n686 B.n685 585
R392 B.n307 B.n306 585
R393 B.n308 B.n307 585
R394 B.n695 B.n694 585
R395 B.n694 B.n693 585
R396 B.n696 B.n305 585
R397 B.n305 B.n304 585
R398 B.n698 B.n697 585
R399 B.n699 B.n698 585
R400 B.n3 B.n0 585
R401 B.n4 B.n3 585
R402 B.n811 B.n1 585
R403 B.n812 B.n811 585
R404 B.n810 B.n809 585
R405 B.n810 B.n8 585
R406 B.n808 B.n9 585
R407 B.n12 B.n9 585
R408 B.n807 B.n806 585
R409 B.n806 B.n805 585
R410 B.n11 B.n10 585
R411 B.n804 B.n11 585
R412 B.n802 B.n801 585
R413 B.n803 B.n802 585
R414 B.n800 B.n17 585
R415 B.n17 B.n16 585
R416 B.n799 B.n798 585
R417 B.n798 B.n797 585
R418 B.n19 B.n18 585
R419 B.n796 B.n19 585
R420 B.n794 B.n793 585
R421 B.n795 B.n794 585
R422 B.n792 B.n24 585
R423 B.n24 B.n23 585
R424 B.n791 B.n790 585
R425 B.n790 B.n789 585
R426 B.n26 B.n25 585
R427 B.n788 B.n26 585
R428 B.n786 B.n785 585
R429 B.n787 B.n786 585
R430 B.n784 B.n31 585
R431 B.n31 B.n30 585
R432 B.n783 B.n782 585
R433 B.n782 B.n781 585
R434 B.n33 B.n32 585
R435 B.n780 B.n33 585
R436 B.n778 B.n777 585
R437 B.n779 B.n778 585
R438 B.n776 B.n38 585
R439 B.n38 B.n37 585
R440 B.n775 B.n774 585
R441 B.n774 B.n773 585
R442 B.n40 B.n39 585
R443 B.n772 B.n40 585
R444 B.n770 B.n769 585
R445 B.n771 B.n770 585
R446 B.n768 B.n44 585
R447 B.n47 B.n44 585
R448 B.n767 B.n766 585
R449 B.n766 B.n765 585
R450 B.n46 B.n45 585
R451 B.n764 B.n46 585
R452 B.n762 B.n761 585
R453 B.n763 B.n762 585
R454 B.n760 B.n52 585
R455 B.n52 B.n51 585
R456 B.n759 B.n758 585
R457 B.n758 B.n757 585
R458 B.n54 B.n53 585
R459 B.n756 B.n54 585
R460 B.n754 B.n753 585
R461 B.n755 B.n754 585
R462 B.n752 B.n59 585
R463 B.n59 B.n58 585
R464 B.n751 B.n750 585
R465 B.n750 B.n749 585
R466 B.n815 B.n814 585
R467 B.n813 B.n2 585
R468 B.n750 B.n61 578.989
R469 B.n747 B.n62 578.989
R470 B.n606 B.n364 578.989
R471 B.n608 B.n362 578.989
R472 B.n114 B.t2 287.122
R473 B.n111 B.t10 287.122
R474 B.n514 B.t6 287.122
R475 B.n391 B.t13 287.122
R476 B.n748 B.n109 256.663
R477 B.n748 B.n108 256.663
R478 B.n748 B.n107 256.663
R479 B.n748 B.n106 256.663
R480 B.n748 B.n105 256.663
R481 B.n748 B.n104 256.663
R482 B.n748 B.n103 256.663
R483 B.n748 B.n102 256.663
R484 B.n748 B.n101 256.663
R485 B.n748 B.n100 256.663
R486 B.n748 B.n99 256.663
R487 B.n748 B.n98 256.663
R488 B.n748 B.n97 256.663
R489 B.n748 B.n96 256.663
R490 B.n748 B.n95 256.663
R491 B.n748 B.n94 256.663
R492 B.n748 B.n93 256.663
R493 B.n748 B.n92 256.663
R494 B.n748 B.n91 256.663
R495 B.n748 B.n90 256.663
R496 B.n748 B.n89 256.663
R497 B.n748 B.n88 256.663
R498 B.n748 B.n87 256.663
R499 B.n748 B.n86 256.663
R500 B.n748 B.n85 256.663
R501 B.n748 B.n84 256.663
R502 B.n748 B.n83 256.663
R503 B.n748 B.n82 256.663
R504 B.n748 B.n81 256.663
R505 B.n748 B.n80 256.663
R506 B.n748 B.n79 256.663
R507 B.n748 B.n78 256.663
R508 B.n748 B.n77 256.663
R509 B.n748 B.n76 256.663
R510 B.n748 B.n75 256.663
R511 B.n748 B.n74 256.663
R512 B.n748 B.n73 256.663
R513 B.n748 B.n72 256.663
R514 B.n748 B.n71 256.663
R515 B.n748 B.n70 256.663
R516 B.n748 B.n69 256.663
R517 B.n748 B.n68 256.663
R518 B.n748 B.n67 256.663
R519 B.n748 B.n66 256.663
R520 B.n748 B.n65 256.663
R521 B.n748 B.n64 256.663
R522 B.n748 B.n63 256.663
R523 B.n413 B.n363 256.663
R524 B.n419 B.n363 256.663
R525 B.n421 B.n363 256.663
R526 B.n427 B.n363 256.663
R527 B.n429 B.n363 256.663
R528 B.n435 B.n363 256.663
R529 B.n437 B.n363 256.663
R530 B.n443 B.n363 256.663
R531 B.n445 B.n363 256.663
R532 B.n451 B.n363 256.663
R533 B.n453 B.n363 256.663
R534 B.n459 B.n363 256.663
R535 B.n461 B.n363 256.663
R536 B.n467 B.n363 256.663
R537 B.n469 B.n363 256.663
R538 B.n475 B.n363 256.663
R539 B.n477 B.n363 256.663
R540 B.n483 B.n363 256.663
R541 B.n485 B.n363 256.663
R542 B.n491 B.n363 256.663
R543 B.n493 B.n363 256.663
R544 B.n500 B.n363 256.663
R545 B.n502 B.n363 256.663
R546 B.n508 B.n363 256.663
R547 B.n510 B.n363 256.663
R548 B.n519 B.n363 256.663
R549 B.n521 B.n363 256.663
R550 B.n527 B.n363 256.663
R551 B.n529 B.n363 256.663
R552 B.n535 B.n363 256.663
R553 B.n537 B.n363 256.663
R554 B.n543 B.n363 256.663
R555 B.n545 B.n363 256.663
R556 B.n551 B.n363 256.663
R557 B.n553 B.n363 256.663
R558 B.n559 B.n363 256.663
R559 B.n561 B.n363 256.663
R560 B.n567 B.n363 256.663
R561 B.n569 B.n363 256.663
R562 B.n575 B.n363 256.663
R563 B.n577 B.n363 256.663
R564 B.n583 B.n363 256.663
R565 B.n585 B.n363 256.663
R566 B.n591 B.n363 256.663
R567 B.n593 B.n363 256.663
R568 B.n599 B.n363 256.663
R569 B.n601 B.n363 256.663
R570 B.n817 B.n816 256.663
R571 B.n118 B.n117 163.367
R572 B.n122 B.n121 163.367
R573 B.n126 B.n125 163.367
R574 B.n130 B.n129 163.367
R575 B.n134 B.n133 163.367
R576 B.n138 B.n137 163.367
R577 B.n142 B.n141 163.367
R578 B.n146 B.n145 163.367
R579 B.n150 B.n149 163.367
R580 B.n154 B.n153 163.367
R581 B.n158 B.n157 163.367
R582 B.n162 B.n161 163.367
R583 B.n166 B.n165 163.367
R584 B.n170 B.n169 163.367
R585 B.n174 B.n173 163.367
R586 B.n178 B.n177 163.367
R587 B.n182 B.n181 163.367
R588 B.n186 B.n185 163.367
R589 B.n190 B.n189 163.367
R590 B.n194 B.n193 163.367
R591 B.n198 B.n197 163.367
R592 B.n203 B.n202 163.367
R593 B.n207 B.n206 163.367
R594 B.n211 B.n210 163.367
R595 B.n215 B.n214 163.367
R596 B.n219 B.n218 163.367
R597 B.n223 B.n222 163.367
R598 B.n227 B.n226 163.367
R599 B.n231 B.n230 163.367
R600 B.n235 B.n234 163.367
R601 B.n239 B.n238 163.367
R602 B.n243 B.n242 163.367
R603 B.n247 B.n246 163.367
R604 B.n251 B.n250 163.367
R605 B.n255 B.n254 163.367
R606 B.n259 B.n258 163.367
R607 B.n263 B.n262 163.367
R608 B.n267 B.n266 163.367
R609 B.n271 B.n270 163.367
R610 B.n275 B.n274 163.367
R611 B.n279 B.n278 163.367
R612 B.n283 B.n282 163.367
R613 B.n287 B.n286 163.367
R614 B.n291 B.n290 163.367
R615 B.n295 B.n294 163.367
R616 B.n299 B.n298 163.367
R617 B.n747 B.n110 163.367
R618 B.n606 B.n358 163.367
R619 B.n614 B.n358 163.367
R620 B.n614 B.n356 163.367
R621 B.n618 B.n356 163.367
R622 B.n618 B.n350 163.367
R623 B.n626 B.n350 163.367
R624 B.n626 B.n348 163.367
R625 B.n630 B.n348 163.367
R626 B.n630 B.n343 163.367
R627 B.n639 B.n343 163.367
R628 B.n639 B.n341 163.367
R629 B.n643 B.n341 163.367
R630 B.n643 B.n335 163.367
R631 B.n651 B.n335 163.367
R632 B.n651 B.n333 163.367
R633 B.n655 B.n333 163.367
R634 B.n655 B.n327 163.367
R635 B.n663 B.n327 163.367
R636 B.n663 B.n325 163.367
R637 B.n667 B.n325 163.367
R638 B.n667 B.n319 163.367
R639 B.n675 B.n319 163.367
R640 B.n675 B.n317 163.367
R641 B.n679 B.n317 163.367
R642 B.n679 B.n311 163.367
R643 B.n687 B.n311 163.367
R644 B.n687 B.n309 163.367
R645 B.n692 B.n309 163.367
R646 B.n692 B.n303 163.367
R647 B.n700 B.n303 163.367
R648 B.n701 B.n700 163.367
R649 B.n701 B.n5 163.367
R650 B.n6 B.n5 163.367
R651 B.n7 B.n6 163.367
R652 B.n707 B.n7 163.367
R653 B.n708 B.n707 163.367
R654 B.n708 B.n13 163.367
R655 B.n14 B.n13 163.367
R656 B.n15 B.n14 163.367
R657 B.n713 B.n15 163.367
R658 B.n713 B.n20 163.367
R659 B.n21 B.n20 163.367
R660 B.n22 B.n21 163.367
R661 B.n718 B.n22 163.367
R662 B.n718 B.n27 163.367
R663 B.n28 B.n27 163.367
R664 B.n29 B.n28 163.367
R665 B.n723 B.n29 163.367
R666 B.n723 B.n34 163.367
R667 B.n35 B.n34 163.367
R668 B.n36 B.n35 163.367
R669 B.n728 B.n36 163.367
R670 B.n728 B.n41 163.367
R671 B.n42 B.n41 163.367
R672 B.n43 B.n42 163.367
R673 B.n733 B.n43 163.367
R674 B.n733 B.n48 163.367
R675 B.n49 B.n48 163.367
R676 B.n50 B.n49 163.367
R677 B.n738 B.n50 163.367
R678 B.n738 B.n55 163.367
R679 B.n56 B.n55 163.367
R680 B.n57 B.n56 163.367
R681 B.n743 B.n57 163.367
R682 B.n743 B.n62 163.367
R683 B.n414 B.n412 163.367
R684 B.n418 B.n412 163.367
R685 B.n422 B.n420 163.367
R686 B.n426 B.n410 163.367
R687 B.n430 B.n428 163.367
R688 B.n434 B.n408 163.367
R689 B.n438 B.n436 163.367
R690 B.n442 B.n406 163.367
R691 B.n446 B.n444 163.367
R692 B.n450 B.n404 163.367
R693 B.n454 B.n452 163.367
R694 B.n458 B.n402 163.367
R695 B.n462 B.n460 163.367
R696 B.n466 B.n400 163.367
R697 B.n470 B.n468 163.367
R698 B.n474 B.n398 163.367
R699 B.n478 B.n476 163.367
R700 B.n482 B.n396 163.367
R701 B.n486 B.n484 163.367
R702 B.n490 B.n394 163.367
R703 B.n494 B.n492 163.367
R704 B.n499 B.n390 163.367
R705 B.n503 B.n501 163.367
R706 B.n507 B.n388 163.367
R707 B.n511 B.n509 163.367
R708 B.n518 B.n386 163.367
R709 B.n522 B.n520 163.367
R710 B.n526 B.n384 163.367
R711 B.n530 B.n528 163.367
R712 B.n534 B.n382 163.367
R713 B.n538 B.n536 163.367
R714 B.n542 B.n380 163.367
R715 B.n546 B.n544 163.367
R716 B.n550 B.n378 163.367
R717 B.n554 B.n552 163.367
R718 B.n558 B.n376 163.367
R719 B.n562 B.n560 163.367
R720 B.n566 B.n374 163.367
R721 B.n570 B.n568 163.367
R722 B.n574 B.n372 163.367
R723 B.n578 B.n576 163.367
R724 B.n582 B.n370 163.367
R725 B.n586 B.n584 163.367
R726 B.n590 B.n368 163.367
R727 B.n594 B.n592 163.367
R728 B.n598 B.n366 163.367
R729 B.n602 B.n600 163.367
R730 B.n608 B.n360 163.367
R731 B.n612 B.n360 163.367
R732 B.n612 B.n354 163.367
R733 B.n620 B.n354 163.367
R734 B.n620 B.n352 163.367
R735 B.n624 B.n352 163.367
R736 B.n624 B.n346 163.367
R737 B.n633 B.n346 163.367
R738 B.n633 B.n344 163.367
R739 B.n637 B.n344 163.367
R740 B.n637 B.n339 163.367
R741 B.n645 B.n339 163.367
R742 B.n645 B.n337 163.367
R743 B.n649 B.n337 163.367
R744 B.n649 B.n331 163.367
R745 B.n657 B.n331 163.367
R746 B.n657 B.n329 163.367
R747 B.n661 B.n329 163.367
R748 B.n661 B.n323 163.367
R749 B.n669 B.n323 163.367
R750 B.n669 B.n321 163.367
R751 B.n673 B.n321 163.367
R752 B.n673 B.n315 163.367
R753 B.n681 B.n315 163.367
R754 B.n681 B.n313 163.367
R755 B.n685 B.n313 163.367
R756 B.n685 B.n307 163.367
R757 B.n694 B.n307 163.367
R758 B.n694 B.n305 163.367
R759 B.n698 B.n305 163.367
R760 B.n698 B.n3 163.367
R761 B.n815 B.n3 163.367
R762 B.n811 B.n2 163.367
R763 B.n811 B.n810 163.367
R764 B.n810 B.n9 163.367
R765 B.n806 B.n9 163.367
R766 B.n806 B.n11 163.367
R767 B.n802 B.n11 163.367
R768 B.n802 B.n17 163.367
R769 B.n798 B.n17 163.367
R770 B.n798 B.n19 163.367
R771 B.n794 B.n19 163.367
R772 B.n794 B.n24 163.367
R773 B.n790 B.n24 163.367
R774 B.n790 B.n26 163.367
R775 B.n786 B.n26 163.367
R776 B.n786 B.n31 163.367
R777 B.n782 B.n31 163.367
R778 B.n782 B.n33 163.367
R779 B.n778 B.n33 163.367
R780 B.n778 B.n38 163.367
R781 B.n774 B.n38 163.367
R782 B.n774 B.n40 163.367
R783 B.n770 B.n40 163.367
R784 B.n770 B.n44 163.367
R785 B.n766 B.n44 163.367
R786 B.n766 B.n46 163.367
R787 B.n762 B.n46 163.367
R788 B.n762 B.n52 163.367
R789 B.n758 B.n52 163.367
R790 B.n758 B.n54 163.367
R791 B.n754 B.n54 163.367
R792 B.n754 B.n59 163.367
R793 B.n750 B.n59 163.367
R794 B.n111 B.t11 153.065
R795 B.n514 B.t9 153.065
R796 B.n114 B.t4 153.048
R797 B.n391 B.t15 153.048
R798 B.n607 B.n363 87.504
R799 B.n749 B.n748 87.504
R800 B.n115 B.n114 81.2611
R801 B.n112 B.n111 81.2611
R802 B.n515 B.n514 81.2611
R803 B.n392 B.n391 81.2611
R804 B.n112 B.t12 71.8035
R805 B.n515 B.t8 71.8035
R806 B.n115 B.t5 71.7877
R807 B.n392 B.t14 71.7877
R808 B.n63 B.n61 71.676
R809 B.n118 B.n64 71.676
R810 B.n122 B.n65 71.676
R811 B.n126 B.n66 71.676
R812 B.n130 B.n67 71.676
R813 B.n134 B.n68 71.676
R814 B.n138 B.n69 71.676
R815 B.n142 B.n70 71.676
R816 B.n146 B.n71 71.676
R817 B.n150 B.n72 71.676
R818 B.n154 B.n73 71.676
R819 B.n158 B.n74 71.676
R820 B.n162 B.n75 71.676
R821 B.n166 B.n76 71.676
R822 B.n170 B.n77 71.676
R823 B.n174 B.n78 71.676
R824 B.n178 B.n79 71.676
R825 B.n182 B.n80 71.676
R826 B.n186 B.n81 71.676
R827 B.n190 B.n82 71.676
R828 B.n194 B.n83 71.676
R829 B.n198 B.n84 71.676
R830 B.n203 B.n85 71.676
R831 B.n207 B.n86 71.676
R832 B.n211 B.n87 71.676
R833 B.n215 B.n88 71.676
R834 B.n219 B.n89 71.676
R835 B.n223 B.n90 71.676
R836 B.n227 B.n91 71.676
R837 B.n231 B.n92 71.676
R838 B.n235 B.n93 71.676
R839 B.n239 B.n94 71.676
R840 B.n243 B.n95 71.676
R841 B.n247 B.n96 71.676
R842 B.n251 B.n97 71.676
R843 B.n255 B.n98 71.676
R844 B.n259 B.n99 71.676
R845 B.n263 B.n100 71.676
R846 B.n267 B.n101 71.676
R847 B.n271 B.n102 71.676
R848 B.n275 B.n103 71.676
R849 B.n279 B.n104 71.676
R850 B.n283 B.n105 71.676
R851 B.n287 B.n106 71.676
R852 B.n291 B.n107 71.676
R853 B.n295 B.n108 71.676
R854 B.n299 B.n109 71.676
R855 B.n110 B.n109 71.676
R856 B.n298 B.n108 71.676
R857 B.n294 B.n107 71.676
R858 B.n290 B.n106 71.676
R859 B.n286 B.n105 71.676
R860 B.n282 B.n104 71.676
R861 B.n278 B.n103 71.676
R862 B.n274 B.n102 71.676
R863 B.n270 B.n101 71.676
R864 B.n266 B.n100 71.676
R865 B.n262 B.n99 71.676
R866 B.n258 B.n98 71.676
R867 B.n254 B.n97 71.676
R868 B.n250 B.n96 71.676
R869 B.n246 B.n95 71.676
R870 B.n242 B.n94 71.676
R871 B.n238 B.n93 71.676
R872 B.n234 B.n92 71.676
R873 B.n230 B.n91 71.676
R874 B.n226 B.n90 71.676
R875 B.n222 B.n89 71.676
R876 B.n218 B.n88 71.676
R877 B.n214 B.n87 71.676
R878 B.n210 B.n86 71.676
R879 B.n206 B.n85 71.676
R880 B.n202 B.n84 71.676
R881 B.n197 B.n83 71.676
R882 B.n193 B.n82 71.676
R883 B.n189 B.n81 71.676
R884 B.n185 B.n80 71.676
R885 B.n181 B.n79 71.676
R886 B.n177 B.n78 71.676
R887 B.n173 B.n77 71.676
R888 B.n169 B.n76 71.676
R889 B.n165 B.n75 71.676
R890 B.n161 B.n74 71.676
R891 B.n157 B.n73 71.676
R892 B.n153 B.n72 71.676
R893 B.n149 B.n71 71.676
R894 B.n145 B.n70 71.676
R895 B.n141 B.n69 71.676
R896 B.n137 B.n68 71.676
R897 B.n133 B.n67 71.676
R898 B.n129 B.n66 71.676
R899 B.n125 B.n65 71.676
R900 B.n121 B.n64 71.676
R901 B.n117 B.n63 71.676
R902 B.n413 B.n362 71.676
R903 B.n419 B.n418 71.676
R904 B.n422 B.n421 71.676
R905 B.n427 B.n426 71.676
R906 B.n430 B.n429 71.676
R907 B.n435 B.n434 71.676
R908 B.n438 B.n437 71.676
R909 B.n443 B.n442 71.676
R910 B.n446 B.n445 71.676
R911 B.n451 B.n450 71.676
R912 B.n454 B.n453 71.676
R913 B.n459 B.n458 71.676
R914 B.n462 B.n461 71.676
R915 B.n467 B.n466 71.676
R916 B.n470 B.n469 71.676
R917 B.n475 B.n474 71.676
R918 B.n478 B.n477 71.676
R919 B.n483 B.n482 71.676
R920 B.n486 B.n485 71.676
R921 B.n491 B.n490 71.676
R922 B.n494 B.n493 71.676
R923 B.n500 B.n499 71.676
R924 B.n503 B.n502 71.676
R925 B.n508 B.n507 71.676
R926 B.n511 B.n510 71.676
R927 B.n519 B.n518 71.676
R928 B.n522 B.n521 71.676
R929 B.n527 B.n526 71.676
R930 B.n530 B.n529 71.676
R931 B.n535 B.n534 71.676
R932 B.n538 B.n537 71.676
R933 B.n543 B.n542 71.676
R934 B.n546 B.n545 71.676
R935 B.n551 B.n550 71.676
R936 B.n554 B.n553 71.676
R937 B.n559 B.n558 71.676
R938 B.n562 B.n561 71.676
R939 B.n567 B.n566 71.676
R940 B.n570 B.n569 71.676
R941 B.n575 B.n574 71.676
R942 B.n578 B.n577 71.676
R943 B.n583 B.n582 71.676
R944 B.n586 B.n585 71.676
R945 B.n591 B.n590 71.676
R946 B.n594 B.n593 71.676
R947 B.n599 B.n598 71.676
R948 B.n602 B.n601 71.676
R949 B.n414 B.n413 71.676
R950 B.n420 B.n419 71.676
R951 B.n421 B.n410 71.676
R952 B.n428 B.n427 71.676
R953 B.n429 B.n408 71.676
R954 B.n436 B.n435 71.676
R955 B.n437 B.n406 71.676
R956 B.n444 B.n443 71.676
R957 B.n445 B.n404 71.676
R958 B.n452 B.n451 71.676
R959 B.n453 B.n402 71.676
R960 B.n460 B.n459 71.676
R961 B.n461 B.n400 71.676
R962 B.n468 B.n467 71.676
R963 B.n469 B.n398 71.676
R964 B.n476 B.n475 71.676
R965 B.n477 B.n396 71.676
R966 B.n484 B.n483 71.676
R967 B.n485 B.n394 71.676
R968 B.n492 B.n491 71.676
R969 B.n493 B.n390 71.676
R970 B.n501 B.n500 71.676
R971 B.n502 B.n388 71.676
R972 B.n509 B.n508 71.676
R973 B.n510 B.n386 71.676
R974 B.n520 B.n519 71.676
R975 B.n521 B.n384 71.676
R976 B.n528 B.n527 71.676
R977 B.n529 B.n382 71.676
R978 B.n536 B.n535 71.676
R979 B.n537 B.n380 71.676
R980 B.n544 B.n543 71.676
R981 B.n545 B.n378 71.676
R982 B.n552 B.n551 71.676
R983 B.n553 B.n376 71.676
R984 B.n560 B.n559 71.676
R985 B.n561 B.n374 71.676
R986 B.n568 B.n567 71.676
R987 B.n569 B.n372 71.676
R988 B.n576 B.n575 71.676
R989 B.n577 B.n370 71.676
R990 B.n584 B.n583 71.676
R991 B.n585 B.n368 71.676
R992 B.n592 B.n591 71.676
R993 B.n593 B.n366 71.676
R994 B.n600 B.n599 71.676
R995 B.n601 B.n364 71.676
R996 B.n816 B.n815 71.676
R997 B.n816 B.n2 71.676
R998 B.n200 B.n115 59.5399
R999 B.n113 B.n112 59.5399
R1000 B.n516 B.n515 59.5399
R1001 B.n497 B.n392 59.5399
R1002 B.n607 B.n359 42.2008
R1003 B.n613 B.n359 42.2008
R1004 B.n613 B.n355 42.2008
R1005 B.n619 B.n355 42.2008
R1006 B.n619 B.n351 42.2008
R1007 B.n625 B.n351 42.2008
R1008 B.n625 B.n347 42.2008
R1009 B.n632 B.n347 42.2008
R1010 B.n632 B.n631 42.2008
R1011 B.n638 B.n340 42.2008
R1012 B.n644 B.n340 42.2008
R1013 B.n644 B.n336 42.2008
R1014 B.n650 B.n336 42.2008
R1015 B.n650 B.n332 42.2008
R1016 B.n656 B.n332 42.2008
R1017 B.n656 B.n328 42.2008
R1018 B.n662 B.n328 42.2008
R1019 B.n662 B.n324 42.2008
R1020 B.n668 B.n324 42.2008
R1021 B.n668 B.n320 42.2008
R1022 B.n674 B.n320 42.2008
R1023 B.n674 B.n316 42.2008
R1024 B.n680 B.n316 42.2008
R1025 B.n686 B.n312 42.2008
R1026 B.n686 B.n308 42.2008
R1027 B.n693 B.n308 42.2008
R1028 B.n693 B.n304 42.2008
R1029 B.n699 B.n304 42.2008
R1030 B.n699 B.n4 42.2008
R1031 B.n814 B.n4 42.2008
R1032 B.n814 B.n813 42.2008
R1033 B.n813 B.n812 42.2008
R1034 B.n812 B.n8 42.2008
R1035 B.n12 B.n8 42.2008
R1036 B.n805 B.n12 42.2008
R1037 B.n805 B.n804 42.2008
R1038 B.n804 B.n803 42.2008
R1039 B.n803 B.n16 42.2008
R1040 B.n797 B.n796 42.2008
R1041 B.n796 B.n795 42.2008
R1042 B.n795 B.n23 42.2008
R1043 B.n789 B.n23 42.2008
R1044 B.n789 B.n788 42.2008
R1045 B.n788 B.n787 42.2008
R1046 B.n787 B.n30 42.2008
R1047 B.n781 B.n30 42.2008
R1048 B.n781 B.n780 42.2008
R1049 B.n780 B.n779 42.2008
R1050 B.n779 B.n37 42.2008
R1051 B.n773 B.n37 42.2008
R1052 B.n773 B.n772 42.2008
R1053 B.n772 B.n771 42.2008
R1054 B.n765 B.n47 42.2008
R1055 B.n765 B.n764 42.2008
R1056 B.n764 B.n763 42.2008
R1057 B.n763 B.n51 42.2008
R1058 B.n757 B.n51 42.2008
R1059 B.n757 B.n756 42.2008
R1060 B.n756 B.n755 42.2008
R1061 B.n755 B.n58 42.2008
R1062 B.n749 B.n58 42.2008
R1063 B.n609 B.n361 37.62
R1064 B.n605 B.n604 37.62
R1065 B.n746 B.n745 37.62
R1066 B.n751 B.n60 37.62
R1067 B.n638 B.t7 33.5125
R1068 B.n771 B.t3 33.5125
R1069 B.n680 B.t0 31.0301
R1070 B.n797 B.t1 31.0301
R1071 B B.n817 18.0485
R1072 B.t0 B.n312 11.1712
R1073 B.t1 B.n16 11.1712
R1074 B.n610 B.n609 10.6151
R1075 B.n611 B.n610 10.6151
R1076 B.n611 B.n353 10.6151
R1077 B.n621 B.n353 10.6151
R1078 B.n622 B.n621 10.6151
R1079 B.n623 B.n622 10.6151
R1080 B.n623 B.n345 10.6151
R1081 B.n634 B.n345 10.6151
R1082 B.n635 B.n634 10.6151
R1083 B.n636 B.n635 10.6151
R1084 B.n636 B.n338 10.6151
R1085 B.n646 B.n338 10.6151
R1086 B.n647 B.n646 10.6151
R1087 B.n648 B.n647 10.6151
R1088 B.n648 B.n330 10.6151
R1089 B.n658 B.n330 10.6151
R1090 B.n659 B.n658 10.6151
R1091 B.n660 B.n659 10.6151
R1092 B.n660 B.n322 10.6151
R1093 B.n670 B.n322 10.6151
R1094 B.n671 B.n670 10.6151
R1095 B.n672 B.n671 10.6151
R1096 B.n672 B.n314 10.6151
R1097 B.n682 B.n314 10.6151
R1098 B.n683 B.n682 10.6151
R1099 B.n684 B.n683 10.6151
R1100 B.n684 B.n306 10.6151
R1101 B.n695 B.n306 10.6151
R1102 B.n696 B.n695 10.6151
R1103 B.n697 B.n696 10.6151
R1104 B.n697 B.n0 10.6151
R1105 B.n415 B.n361 10.6151
R1106 B.n416 B.n415 10.6151
R1107 B.n417 B.n416 10.6151
R1108 B.n417 B.n411 10.6151
R1109 B.n423 B.n411 10.6151
R1110 B.n424 B.n423 10.6151
R1111 B.n425 B.n424 10.6151
R1112 B.n425 B.n409 10.6151
R1113 B.n431 B.n409 10.6151
R1114 B.n432 B.n431 10.6151
R1115 B.n433 B.n432 10.6151
R1116 B.n433 B.n407 10.6151
R1117 B.n439 B.n407 10.6151
R1118 B.n440 B.n439 10.6151
R1119 B.n441 B.n440 10.6151
R1120 B.n441 B.n405 10.6151
R1121 B.n447 B.n405 10.6151
R1122 B.n448 B.n447 10.6151
R1123 B.n449 B.n448 10.6151
R1124 B.n449 B.n403 10.6151
R1125 B.n455 B.n403 10.6151
R1126 B.n456 B.n455 10.6151
R1127 B.n457 B.n456 10.6151
R1128 B.n457 B.n401 10.6151
R1129 B.n463 B.n401 10.6151
R1130 B.n464 B.n463 10.6151
R1131 B.n465 B.n464 10.6151
R1132 B.n465 B.n399 10.6151
R1133 B.n471 B.n399 10.6151
R1134 B.n472 B.n471 10.6151
R1135 B.n473 B.n472 10.6151
R1136 B.n473 B.n397 10.6151
R1137 B.n479 B.n397 10.6151
R1138 B.n480 B.n479 10.6151
R1139 B.n481 B.n480 10.6151
R1140 B.n481 B.n395 10.6151
R1141 B.n487 B.n395 10.6151
R1142 B.n488 B.n487 10.6151
R1143 B.n489 B.n488 10.6151
R1144 B.n489 B.n393 10.6151
R1145 B.n495 B.n393 10.6151
R1146 B.n496 B.n495 10.6151
R1147 B.n498 B.n389 10.6151
R1148 B.n504 B.n389 10.6151
R1149 B.n505 B.n504 10.6151
R1150 B.n506 B.n505 10.6151
R1151 B.n506 B.n387 10.6151
R1152 B.n512 B.n387 10.6151
R1153 B.n513 B.n512 10.6151
R1154 B.n517 B.n513 10.6151
R1155 B.n523 B.n385 10.6151
R1156 B.n524 B.n523 10.6151
R1157 B.n525 B.n524 10.6151
R1158 B.n525 B.n383 10.6151
R1159 B.n531 B.n383 10.6151
R1160 B.n532 B.n531 10.6151
R1161 B.n533 B.n532 10.6151
R1162 B.n533 B.n381 10.6151
R1163 B.n539 B.n381 10.6151
R1164 B.n540 B.n539 10.6151
R1165 B.n541 B.n540 10.6151
R1166 B.n541 B.n379 10.6151
R1167 B.n547 B.n379 10.6151
R1168 B.n548 B.n547 10.6151
R1169 B.n549 B.n548 10.6151
R1170 B.n549 B.n377 10.6151
R1171 B.n555 B.n377 10.6151
R1172 B.n556 B.n555 10.6151
R1173 B.n557 B.n556 10.6151
R1174 B.n557 B.n375 10.6151
R1175 B.n563 B.n375 10.6151
R1176 B.n564 B.n563 10.6151
R1177 B.n565 B.n564 10.6151
R1178 B.n565 B.n373 10.6151
R1179 B.n571 B.n373 10.6151
R1180 B.n572 B.n571 10.6151
R1181 B.n573 B.n572 10.6151
R1182 B.n573 B.n371 10.6151
R1183 B.n579 B.n371 10.6151
R1184 B.n580 B.n579 10.6151
R1185 B.n581 B.n580 10.6151
R1186 B.n581 B.n369 10.6151
R1187 B.n587 B.n369 10.6151
R1188 B.n588 B.n587 10.6151
R1189 B.n589 B.n588 10.6151
R1190 B.n589 B.n367 10.6151
R1191 B.n595 B.n367 10.6151
R1192 B.n596 B.n595 10.6151
R1193 B.n597 B.n596 10.6151
R1194 B.n597 B.n365 10.6151
R1195 B.n603 B.n365 10.6151
R1196 B.n604 B.n603 10.6151
R1197 B.n605 B.n357 10.6151
R1198 B.n615 B.n357 10.6151
R1199 B.n616 B.n615 10.6151
R1200 B.n617 B.n616 10.6151
R1201 B.n617 B.n349 10.6151
R1202 B.n627 B.n349 10.6151
R1203 B.n628 B.n627 10.6151
R1204 B.n629 B.n628 10.6151
R1205 B.n629 B.n342 10.6151
R1206 B.n640 B.n342 10.6151
R1207 B.n641 B.n640 10.6151
R1208 B.n642 B.n641 10.6151
R1209 B.n642 B.n334 10.6151
R1210 B.n652 B.n334 10.6151
R1211 B.n653 B.n652 10.6151
R1212 B.n654 B.n653 10.6151
R1213 B.n654 B.n326 10.6151
R1214 B.n664 B.n326 10.6151
R1215 B.n665 B.n664 10.6151
R1216 B.n666 B.n665 10.6151
R1217 B.n666 B.n318 10.6151
R1218 B.n676 B.n318 10.6151
R1219 B.n677 B.n676 10.6151
R1220 B.n678 B.n677 10.6151
R1221 B.n678 B.n310 10.6151
R1222 B.n688 B.n310 10.6151
R1223 B.n689 B.n688 10.6151
R1224 B.n691 B.n689 10.6151
R1225 B.n691 B.n690 10.6151
R1226 B.n690 B.n302 10.6151
R1227 B.n702 B.n302 10.6151
R1228 B.n703 B.n702 10.6151
R1229 B.n704 B.n703 10.6151
R1230 B.n705 B.n704 10.6151
R1231 B.n706 B.n705 10.6151
R1232 B.n709 B.n706 10.6151
R1233 B.n710 B.n709 10.6151
R1234 B.n711 B.n710 10.6151
R1235 B.n712 B.n711 10.6151
R1236 B.n714 B.n712 10.6151
R1237 B.n715 B.n714 10.6151
R1238 B.n716 B.n715 10.6151
R1239 B.n717 B.n716 10.6151
R1240 B.n719 B.n717 10.6151
R1241 B.n720 B.n719 10.6151
R1242 B.n721 B.n720 10.6151
R1243 B.n722 B.n721 10.6151
R1244 B.n724 B.n722 10.6151
R1245 B.n725 B.n724 10.6151
R1246 B.n726 B.n725 10.6151
R1247 B.n727 B.n726 10.6151
R1248 B.n729 B.n727 10.6151
R1249 B.n730 B.n729 10.6151
R1250 B.n731 B.n730 10.6151
R1251 B.n732 B.n731 10.6151
R1252 B.n734 B.n732 10.6151
R1253 B.n735 B.n734 10.6151
R1254 B.n736 B.n735 10.6151
R1255 B.n737 B.n736 10.6151
R1256 B.n739 B.n737 10.6151
R1257 B.n740 B.n739 10.6151
R1258 B.n741 B.n740 10.6151
R1259 B.n742 B.n741 10.6151
R1260 B.n744 B.n742 10.6151
R1261 B.n745 B.n744 10.6151
R1262 B.n809 B.n1 10.6151
R1263 B.n809 B.n808 10.6151
R1264 B.n808 B.n807 10.6151
R1265 B.n807 B.n10 10.6151
R1266 B.n801 B.n10 10.6151
R1267 B.n801 B.n800 10.6151
R1268 B.n800 B.n799 10.6151
R1269 B.n799 B.n18 10.6151
R1270 B.n793 B.n18 10.6151
R1271 B.n793 B.n792 10.6151
R1272 B.n792 B.n791 10.6151
R1273 B.n791 B.n25 10.6151
R1274 B.n785 B.n25 10.6151
R1275 B.n785 B.n784 10.6151
R1276 B.n784 B.n783 10.6151
R1277 B.n783 B.n32 10.6151
R1278 B.n777 B.n32 10.6151
R1279 B.n777 B.n776 10.6151
R1280 B.n776 B.n775 10.6151
R1281 B.n775 B.n39 10.6151
R1282 B.n769 B.n39 10.6151
R1283 B.n769 B.n768 10.6151
R1284 B.n768 B.n767 10.6151
R1285 B.n767 B.n45 10.6151
R1286 B.n761 B.n45 10.6151
R1287 B.n761 B.n760 10.6151
R1288 B.n760 B.n759 10.6151
R1289 B.n759 B.n53 10.6151
R1290 B.n753 B.n53 10.6151
R1291 B.n753 B.n752 10.6151
R1292 B.n752 B.n751 10.6151
R1293 B.n116 B.n60 10.6151
R1294 B.n119 B.n116 10.6151
R1295 B.n120 B.n119 10.6151
R1296 B.n123 B.n120 10.6151
R1297 B.n124 B.n123 10.6151
R1298 B.n127 B.n124 10.6151
R1299 B.n128 B.n127 10.6151
R1300 B.n131 B.n128 10.6151
R1301 B.n132 B.n131 10.6151
R1302 B.n135 B.n132 10.6151
R1303 B.n136 B.n135 10.6151
R1304 B.n139 B.n136 10.6151
R1305 B.n140 B.n139 10.6151
R1306 B.n143 B.n140 10.6151
R1307 B.n144 B.n143 10.6151
R1308 B.n147 B.n144 10.6151
R1309 B.n148 B.n147 10.6151
R1310 B.n151 B.n148 10.6151
R1311 B.n152 B.n151 10.6151
R1312 B.n155 B.n152 10.6151
R1313 B.n156 B.n155 10.6151
R1314 B.n159 B.n156 10.6151
R1315 B.n160 B.n159 10.6151
R1316 B.n163 B.n160 10.6151
R1317 B.n164 B.n163 10.6151
R1318 B.n167 B.n164 10.6151
R1319 B.n168 B.n167 10.6151
R1320 B.n171 B.n168 10.6151
R1321 B.n172 B.n171 10.6151
R1322 B.n175 B.n172 10.6151
R1323 B.n176 B.n175 10.6151
R1324 B.n179 B.n176 10.6151
R1325 B.n180 B.n179 10.6151
R1326 B.n183 B.n180 10.6151
R1327 B.n184 B.n183 10.6151
R1328 B.n187 B.n184 10.6151
R1329 B.n188 B.n187 10.6151
R1330 B.n191 B.n188 10.6151
R1331 B.n192 B.n191 10.6151
R1332 B.n195 B.n192 10.6151
R1333 B.n196 B.n195 10.6151
R1334 B.n199 B.n196 10.6151
R1335 B.n204 B.n201 10.6151
R1336 B.n205 B.n204 10.6151
R1337 B.n208 B.n205 10.6151
R1338 B.n209 B.n208 10.6151
R1339 B.n212 B.n209 10.6151
R1340 B.n213 B.n212 10.6151
R1341 B.n216 B.n213 10.6151
R1342 B.n217 B.n216 10.6151
R1343 B.n221 B.n220 10.6151
R1344 B.n224 B.n221 10.6151
R1345 B.n225 B.n224 10.6151
R1346 B.n228 B.n225 10.6151
R1347 B.n229 B.n228 10.6151
R1348 B.n232 B.n229 10.6151
R1349 B.n233 B.n232 10.6151
R1350 B.n236 B.n233 10.6151
R1351 B.n237 B.n236 10.6151
R1352 B.n240 B.n237 10.6151
R1353 B.n241 B.n240 10.6151
R1354 B.n244 B.n241 10.6151
R1355 B.n245 B.n244 10.6151
R1356 B.n248 B.n245 10.6151
R1357 B.n249 B.n248 10.6151
R1358 B.n252 B.n249 10.6151
R1359 B.n253 B.n252 10.6151
R1360 B.n256 B.n253 10.6151
R1361 B.n257 B.n256 10.6151
R1362 B.n260 B.n257 10.6151
R1363 B.n261 B.n260 10.6151
R1364 B.n264 B.n261 10.6151
R1365 B.n265 B.n264 10.6151
R1366 B.n268 B.n265 10.6151
R1367 B.n269 B.n268 10.6151
R1368 B.n272 B.n269 10.6151
R1369 B.n273 B.n272 10.6151
R1370 B.n276 B.n273 10.6151
R1371 B.n277 B.n276 10.6151
R1372 B.n280 B.n277 10.6151
R1373 B.n281 B.n280 10.6151
R1374 B.n284 B.n281 10.6151
R1375 B.n285 B.n284 10.6151
R1376 B.n288 B.n285 10.6151
R1377 B.n289 B.n288 10.6151
R1378 B.n292 B.n289 10.6151
R1379 B.n293 B.n292 10.6151
R1380 B.n296 B.n293 10.6151
R1381 B.n297 B.n296 10.6151
R1382 B.n300 B.n297 10.6151
R1383 B.n301 B.n300 10.6151
R1384 B.n746 B.n301 10.6151
R1385 B.n631 B.t7 8.68879
R1386 B.n47 B.t3 8.68879
R1387 B.n817 B.n0 8.11757
R1388 B.n817 B.n1 8.11757
R1389 B.n498 B.n497 6.5566
R1390 B.n517 B.n516 6.5566
R1391 B.n201 B.n200 6.5566
R1392 B.n217 B.n113 6.5566
R1393 B.n497 B.n496 4.05904
R1394 B.n516 B.n385 4.05904
R1395 B.n200 B.n199 4.05904
R1396 B.n220 B.n113 4.05904
R1397 VN VN.t1 160.921
R1398 VN VN.t0 113.391
R1399 VDD2.n0 VDD2.t1 104.412
R1400 VDD2.n0 VDD2.t0 62.7959
R1401 VDD2 VDD2.n0 0.961707
C0 VDD2 VN 3.02582f
C1 VDD1 VP 3.26105f
C2 VDD2 VTAIL 5.50042f
C3 VTAIL VN 2.74774f
C4 VDD2 VP 0.38541f
C5 VN VP 6.1316f
C6 VTAIL VP 2.7626f
C7 VDD1 VDD2 0.815613f
C8 VDD1 VN 0.148701f
C9 VDD1 VTAIL 5.44043f
C10 VDD2 B 4.967563f
C11 VDD1 B 8.400661f
C12 VTAIL B 8.139374f
C13 VN B 12.065539f
C14 VP B 7.996813f
C15 VDD2.t1 B 2.91234f
C16 VDD2.t0 B 2.28413f
C17 VDD2.n0 B 3.12112f
C18 VN.t0 B 3.53199f
C19 VN.t1 B 4.22876f
C20 VDD1.t1 B 2.32185f
C21 VDD1.t0 B 3.00129f
C22 VTAIL.t3 B 2.27754f
C23 VTAIL.n0 B 1.88771f
C24 VTAIL.t0 B 2.27756f
C25 VTAIL.n1 B 1.94506f
C26 VTAIL.t2 B 2.27754f
C27 VTAIL.n2 B 1.69984f
C28 VTAIL.t1 B 2.27754f
C29 VTAIL.n3 B 1.60268f
C30 VP.t0 B 4.386509f
C31 VP.t1 B 3.65595f
C32 VP.n0 B 4.0505f
.ends

