* NGSPICE file created from diff_pair_sample_1405.ext - technology: sky130A

.subckt diff_pair_sample_1405 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t9 VN.t0 VTAIL.t10 w_n5674_n2424# sky130_fd_pr__pfet_01v8 ad=1.2012 pd=7.61 as=1.2012 ps=7.61 w=7.28 l=3.59
X1 VDD2.t8 VN.t1 VTAIL.t18 w_n5674_n2424# sky130_fd_pr__pfet_01v8 ad=2.8392 pd=15.34 as=1.2012 ps=7.61 w=7.28 l=3.59
X2 VTAIL.t5 VP.t0 VDD1.t9 w_n5674_n2424# sky130_fd_pr__pfet_01v8 ad=1.2012 pd=7.61 as=1.2012 ps=7.61 w=7.28 l=3.59
X3 VTAIL.t9 VP.t1 VDD1.t8 w_n5674_n2424# sky130_fd_pr__pfet_01v8 ad=1.2012 pd=7.61 as=1.2012 ps=7.61 w=7.28 l=3.59
X4 B.t11 B.t9 B.t10 w_n5674_n2424# sky130_fd_pr__pfet_01v8 ad=2.8392 pd=15.34 as=0 ps=0 w=7.28 l=3.59
X5 VDD2.t7 VN.t2 VTAIL.t14 w_n5674_n2424# sky130_fd_pr__pfet_01v8 ad=1.2012 pd=7.61 as=1.2012 ps=7.61 w=7.28 l=3.59
X6 VTAIL.t4 VP.t2 VDD1.t7 w_n5674_n2424# sky130_fd_pr__pfet_01v8 ad=1.2012 pd=7.61 as=1.2012 ps=7.61 w=7.28 l=3.59
X7 VTAIL.t19 VN.t3 VDD2.t6 w_n5674_n2424# sky130_fd_pr__pfet_01v8 ad=1.2012 pd=7.61 as=1.2012 ps=7.61 w=7.28 l=3.59
X8 VTAIL.t13 VN.t4 VDD2.t5 w_n5674_n2424# sky130_fd_pr__pfet_01v8 ad=1.2012 pd=7.61 as=1.2012 ps=7.61 w=7.28 l=3.59
X9 VDD1.t6 VP.t3 VTAIL.t3 w_n5674_n2424# sky130_fd_pr__pfet_01v8 ad=1.2012 pd=7.61 as=2.8392 ps=15.34 w=7.28 l=3.59
X10 VDD2.t4 VN.t5 VTAIL.t15 w_n5674_n2424# sky130_fd_pr__pfet_01v8 ad=2.8392 pd=15.34 as=1.2012 ps=7.61 w=7.28 l=3.59
X11 VDD1.t5 VP.t4 VTAIL.t7 w_n5674_n2424# sky130_fd_pr__pfet_01v8 ad=2.8392 pd=15.34 as=1.2012 ps=7.61 w=7.28 l=3.59
X12 VDD2.t3 VN.t6 VTAIL.t12 w_n5674_n2424# sky130_fd_pr__pfet_01v8 ad=1.2012 pd=7.61 as=2.8392 ps=15.34 w=7.28 l=3.59
X13 VTAIL.t16 VN.t7 VDD2.t2 w_n5674_n2424# sky130_fd_pr__pfet_01v8 ad=1.2012 pd=7.61 as=1.2012 ps=7.61 w=7.28 l=3.59
X14 VDD2.t1 VN.t8 VTAIL.t11 w_n5674_n2424# sky130_fd_pr__pfet_01v8 ad=1.2012 pd=7.61 as=2.8392 ps=15.34 w=7.28 l=3.59
X15 VDD1.t4 VP.t5 VTAIL.t0 w_n5674_n2424# sky130_fd_pr__pfet_01v8 ad=2.8392 pd=15.34 as=1.2012 ps=7.61 w=7.28 l=3.59
X16 VTAIL.t17 VN.t9 VDD2.t0 w_n5674_n2424# sky130_fd_pr__pfet_01v8 ad=1.2012 pd=7.61 as=1.2012 ps=7.61 w=7.28 l=3.59
X17 B.t8 B.t6 B.t7 w_n5674_n2424# sky130_fd_pr__pfet_01v8 ad=2.8392 pd=15.34 as=0 ps=0 w=7.28 l=3.59
X18 VDD1.t3 VP.t6 VTAIL.t8 w_n5674_n2424# sky130_fd_pr__pfet_01v8 ad=1.2012 pd=7.61 as=1.2012 ps=7.61 w=7.28 l=3.59
X19 VDD1.t2 VP.t7 VTAIL.t6 w_n5674_n2424# sky130_fd_pr__pfet_01v8 ad=1.2012 pd=7.61 as=2.8392 ps=15.34 w=7.28 l=3.59
X20 B.t5 B.t3 B.t4 w_n5674_n2424# sky130_fd_pr__pfet_01v8 ad=2.8392 pd=15.34 as=0 ps=0 w=7.28 l=3.59
X21 VTAIL.t1 VP.t8 VDD1.t1 w_n5674_n2424# sky130_fd_pr__pfet_01v8 ad=1.2012 pd=7.61 as=1.2012 ps=7.61 w=7.28 l=3.59
X22 B.t2 B.t0 B.t1 w_n5674_n2424# sky130_fd_pr__pfet_01v8 ad=2.8392 pd=15.34 as=0 ps=0 w=7.28 l=3.59
X23 VDD1.t0 VP.t9 VTAIL.t2 w_n5674_n2424# sky130_fd_pr__pfet_01v8 ad=1.2012 pd=7.61 as=1.2012 ps=7.61 w=7.28 l=3.59
R0 VN.n106 VN.n105 161.3
R1 VN.n104 VN.n55 161.3
R2 VN.n103 VN.n102 161.3
R3 VN.n101 VN.n56 161.3
R4 VN.n100 VN.n99 161.3
R5 VN.n98 VN.n57 161.3
R6 VN.n97 VN.n96 161.3
R7 VN.n95 VN.n58 161.3
R8 VN.n94 VN.n93 161.3
R9 VN.n92 VN.n59 161.3
R10 VN.n91 VN.n90 161.3
R11 VN.n89 VN.n61 161.3
R12 VN.n88 VN.n87 161.3
R13 VN.n86 VN.n62 161.3
R14 VN.n85 VN.n84 161.3
R15 VN.n83 VN.n63 161.3
R16 VN.n82 VN.n81 161.3
R17 VN.n80 VN.n64 161.3
R18 VN.n79 VN.n78 161.3
R19 VN.n77 VN.n66 161.3
R20 VN.n76 VN.n75 161.3
R21 VN.n74 VN.n67 161.3
R22 VN.n73 VN.n72 161.3
R23 VN.n71 VN.n68 161.3
R24 VN.n52 VN.n51 161.3
R25 VN.n50 VN.n1 161.3
R26 VN.n49 VN.n48 161.3
R27 VN.n47 VN.n2 161.3
R28 VN.n46 VN.n45 161.3
R29 VN.n44 VN.n3 161.3
R30 VN.n43 VN.n42 161.3
R31 VN.n41 VN.n4 161.3
R32 VN.n40 VN.n39 161.3
R33 VN.n37 VN.n5 161.3
R34 VN.n36 VN.n35 161.3
R35 VN.n34 VN.n6 161.3
R36 VN.n33 VN.n32 161.3
R37 VN.n31 VN.n7 161.3
R38 VN.n30 VN.n29 161.3
R39 VN.n28 VN.n8 161.3
R40 VN.n27 VN.n26 161.3
R41 VN.n24 VN.n9 161.3
R42 VN.n23 VN.n22 161.3
R43 VN.n21 VN.n10 161.3
R44 VN.n20 VN.n19 161.3
R45 VN.n18 VN.n11 161.3
R46 VN.n17 VN.n16 161.3
R47 VN.n15 VN.n12 161.3
R48 VN.n53 VN.n0 85.819
R49 VN.n107 VN.n54 85.819
R50 VN.n70 VN.t6 81.2364
R51 VN.n14 VN.t5 81.2364
R52 VN.n14 VN.n13 66.4721
R53 VN.n70 VN.n69 66.4721
R54 VN.n19 VN.n10 56.5617
R55 VN.n32 VN.n6 56.5617
R56 VN.n75 VN.n66 56.5617
R57 VN.n87 VN.n61 56.5617
R58 VN VN.n107 55.1118
R59 VN.n45 VN.n2 53.171
R60 VN.n99 VN.n56 53.171
R61 VN.n13 VN.t9 48.8718
R62 VN.n25 VN.t0 48.8718
R63 VN.n38 VN.t3 48.8718
R64 VN.n0 VN.t8 48.8718
R65 VN.n69 VN.t4 48.8718
R66 VN.n65 VN.t2 48.8718
R67 VN.n60 VN.t7 48.8718
R68 VN.n54 VN.t1 48.8718
R69 VN.n45 VN.n44 27.983
R70 VN.n99 VN.n98 27.983
R71 VN.n17 VN.n12 24.5923
R72 VN.n18 VN.n17 24.5923
R73 VN.n19 VN.n18 24.5923
R74 VN.n23 VN.n10 24.5923
R75 VN.n24 VN.n23 24.5923
R76 VN.n26 VN.n24 24.5923
R77 VN.n30 VN.n8 24.5923
R78 VN.n31 VN.n30 24.5923
R79 VN.n32 VN.n31 24.5923
R80 VN.n36 VN.n6 24.5923
R81 VN.n37 VN.n36 24.5923
R82 VN.n39 VN.n37 24.5923
R83 VN.n43 VN.n4 24.5923
R84 VN.n44 VN.n43 24.5923
R85 VN.n49 VN.n2 24.5923
R86 VN.n50 VN.n49 24.5923
R87 VN.n51 VN.n50 24.5923
R88 VN.n75 VN.n74 24.5923
R89 VN.n74 VN.n73 24.5923
R90 VN.n73 VN.n68 24.5923
R91 VN.n87 VN.n86 24.5923
R92 VN.n86 VN.n85 24.5923
R93 VN.n85 VN.n63 24.5923
R94 VN.n81 VN.n80 24.5923
R95 VN.n80 VN.n79 24.5923
R96 VN.n79 VN.n66 24.5923
R97 VN.n98 VN.n97 24.5923
R98 VN.n97 VN.n58 24.5923
R99 VN.n93 VN.n92 24.5923
R100 VN.n92 VN.n91 24.5923
R101 VN.n91 VN.n61 24.5923
R102 VN.n105 VN.n104 24.5923
R103 VN.n104 VN.n103 24.5923
R104 VN.n103 VN.n56 24.5923
R105 VN.n38 VN.n4 16.2311
R106 VN.n60 VN.n58 16.2311
R107 VN.n26 VN.n25 12.2964
R108 VN.n25 VN.n8 12.2964
R109 VN.n65 VN.n63 12.2964
R110 VN.n81 VN.n65 12.2964
R111 VN.n13 VN.n12 8.36172
R112 VN.n39 VN.n38 8.36172
R113 VN.n69 VN.n68 8.36172
R114 VN.n93 VN.n60 8.36172
R115 VN.n51 VN.n0 4.42703
R116 VN.n105 VN.n54 4.42703
R117 VN.n71 VN.n70 3.32151
R118 VN.n15 VN.n14 3.32151
R119 VN.n107 VN.n106 0.354861
R120 VN.n53 VN.n52 0.354861
R121 VN VN.n53 0.267071
R122 VN.n106 VN.n55 0.189894
R123 VN.n102 VN.n55 0.189894
R124 VN.n102 VN.n101 0.189894
R125 VN.n101 VN.n100 0.189894
R126 VN.n100 VN.n57 0.189894
R127 VN.n96 VN.n57 0.189894
R128 VN.n96 VN.n95 0.189894
R129 VN.n95 VN.n94 0.189894
R130 VN.n94 VN.n59 0.189894
R131 VN.n90 VN.n59 0.189894
R132 VN.n90 VN.n89 0.189894
R133 VN.n89 VN.n88 0.189894
R134 VN.n88 VN.n62 0.189894
R135 VN.n84 VN.n62 0.189894
R136 VN.n84 VN.n83 0.189894
R137 VN.n83 VN.n82 0.189894
R138 VN.n82 VN.n64 0.189894
R139 VN.n78 VN.n64 0.189894
R140 VN.n78 VN.n77 0.189894
R141 VN.n77 VN.n76 0.189894
R142 VN.n76 VN.n67 0.189894
R143 VN.n72 VN.n67 0.189894
R144 VN.n72 VN.n71 0.189894
R145 VN.n16 VN.n15 0.189894
R146 VN.n16 VN.n11 0.189894
R147 VN.n20 VN.n11 0.189894
R148 VN.n21 VN.n20 0.189894
R149 VN.n22 VN.n21 0.189894
R150 VN.n22 VN.n9 0.189894
R151 VN.n27 VN.n9 0.189894
R152 VN.n28 VN.n27 0.189894
R153 VN.n29 VN.n28 0.189894
R154 VN.n29 VN.n7 0.189894
R155 VN.n33 VN.n7 0.189894
R156 VN.n34 VN.n33 0.189894
R157 VN.n35 VN.n34 0.189894
R158 VN.n35 VN.n5 0.189894
R159 VN.n40 VN.n5 0.189894
R160 VN.n41 VN.n40 0.189894
R161 VN.n42 VN.n41 0.189894
R162 VN.n42 VN.n3 0.189894
R163 VN.n46 VN.n3 0.189894
R164 VN.n47 VN.n46 0.189894
R165 VN.n48 VN.n47 0.189894
R166 VN.n48 VN.n1 0.189894
R167 VN.n52 VN.n1 0.189894
R168 VTAIL.n135 VTAIL.n134 585
R169 VTAIL.n137 VTAIL.n136 585
R170 VTAIL.n130 VTAIL.n129 585
R171 VTAIL.n143 VTAIL.n142 585
R172 VTAIL.n145 VTAIL.n144 585
R173 VTAIL.n126 VTAIL.n125 585
R174 VTAIL.n151 VTAIL.n150 585
R175 VTAIL.n153 VTAIL.n152 585
R176 VTAIL.n15 VTAIL.n14 585
R177 VTAIL.n17 VTAIL.n16 585
R178 VTAIL.n10 VTAIL.n9 585
R179 VTAIL.n23 VTAIL.n22 585
R180 VTAIL.n25 VTAIL.n24 585
R181 VTAIL.n6 VTAIL.n5 585
R182 VTAIL.n31 VTAIL.n30 585
R183 VTAIL.n33 VTAIL.n32 585
R184 VTAIL.n117 VTAIL.n116 585
R185 VTAIL.n115 VTAIL.n114 585
R186 VTAIL.n90 VTAIL.n89 585
R187 VTAIL.n109 VTAIL.n108 585
R188 VTAIL.n107 VTAIL.n106 585
R189 VTAIL.n94 VTAIL.n93 585
R190 VTAIL.n101 VTAIL.n100 585
R191 VTAIL.n99 VTAIL.n98 585
R192 VTAIL.n77 VTAIL.n76 585
R193 VTAIL.n75 VTAIL.n74 585
R194 VTAIL.n50 VTAIL.n49 585
R195 VTAIL.n69 VTAIL.n68 585
R196 VTAIL.n67 VTAIL.n66 585
R197 VTAIL.n54 VTAIL.n53 585
R198 VTAIL.n61 VTAIL.n60 585
R199 VTAIL.n59 VTAIL.n58 585
R200 VTAIL.n152 VTAIL.n122 498.474
R201 VTAIL.n32 VTAIL.n2 498.474
R202 VTAIL.n116 VTAIL.n86 498.474
R203 VTAIL.n76 VTAIL.n46 498.474
R204 VTAIL.n133 VTAIL.t11 329.053
R205 VTAIL.n13 VTAIL.t3 329.053
R206 VTAIL.n97 VTAIL.t6 329.053
R207 VTAIL.n57 VTAIL.t12 329.053
R208 VTAIL.n136 VTAIL.n135 171.744
R209 VTAIL.n136 VTAIL.n129 171.744
R210 VTAIL.n143 VTAIL.n129 171.744
R211 VTAIL.n144 VTAIL.n143 171.744
R212 VTAIL.n144 VTAIL.n125 171.744
R213 VTAIL.n151 VTAIL.n125 171.744
R214 VTAIL.n152 VTAIL.n151 171.744
R215 VTAIL.n16 VTAIL.n15 171.744
R216 VTAIL.n16 VTAIL.n9 171.744
R217 VTAIL.n23 VTAIL.n9 171.744
R218 VTAIL.n24 VTAIL.n23 171.744
R219 VTAIL.n24 VTAIL.n5 171.744
R220 VTAIL.n31 VTAIL.n5 171.744
R221 VTAIL.n32 VTAIL.n31 171.744
R222 VTAIL.n116 VTAIL.n115 171.744
R223 VTAIL.n115 VTAIL.n89 171.744
R224 VTAIL.n108 VTAIL.n89 171.744
R225 VTAIL.n108 VTAIL.n107 171.744
R226 VTAIL.n107 VTAIL.n93 171.744
R227 VTAIL.n100 VTAIL.n93 171.744
R228 VTAIL.n100 VTAIL.n99 171.744
R229 VTAIL.n76 VTAIL.n75 171.744
R230 VTAIL.n75 VTAIL.n49 171.744
R231 VTAIL.n68 VTAIL.n49 171.744
R232 VTAIL.n68 VTAIL.n67 171.744
R233 VTAIL.n67 VTAIL.n53 171.744
R234 VTAIL.n60 VTAIL.n53 171.744
R235 VTAIL.n60 VTAIL.n59 171.744
R236 VTAIL.n135 VTAIL.t11 85.8723
R237 VTAIL.n15 VTAIL.t3 85.8723
R238 VTAIL.n99 VTAIL.t6 85.8723
R239 VTAIL.n59 VTAIL.t12 85.8723
R240 VTAIL.n85 VTAIL.n84 72.0388
R241 VTAIL.n83 VTAIL.n82 72.0388
R242 VTAIL.n45 VTAIL.n44 72.0388
R243 VTAIL.n43 VTAIL.n42 72.0388
R244 VTAIL.n159 VTAIL.n158 72.0387
R245 VTAIL.n1 VTAIL.n0 72.0387
R246 VTAIL.n39 VTAIL.n38 72.0387
R247 VTAIL.n41 VTAIL.n40 72.0387
R248 VTAIL.n157 VTAIL.n156 36.0641
R249 VTAIL.n37 VTAIL.n36 36.0641
R250 VTAIL.n121 VTAIL.n120 36.0641
R251 VTAIL.n81 VTAIL.n80 36.0641
R252 VTAIL.n43 VTAIL.n41 25.4014
R253 VTAIL.n157 VTAIL.n121 22.0221
R254 VTAIL.n154 VTAIL.n153 12.8005
R255 VTAIL.n34 VTAIL.n33 12.8005
R256 VTAIL.n118 VTAIL.n117 12.8005
R257 VTAIL.n78 VTAIL.n77 12.8005
R258 VTAIL.n150 VTAIL.n124 12.0247
R259 VTAIL.n30 VTAIL.n4 12.0247
R260 VTAIL.n114 VTAIL.n88 12.0247
R261 VTAIL.n74 VTAIL.n48 12.0247
R262 VTAIL.n149 VTAIL.n126 11.249
R263 VTAIL.n29 VTAIL.n6 11.249
R264 VTAIL.n113 VTAIL.n90 11.249
R265 VTAIL.n73 VTAIL.n50 11.249
R266 VTAIL.n134 VTAIL.n133 10.7237
R267 VTAIL.n14 VTAIL.n13 10.7237
R268 VTAIL.n98 VTAIL.n97 10.7237
R269 VTAIL.n58 VTAIL.n57 10.7237
R270 VTAIL.n146 VTAIL.n145 10.4732
R271 VTAIL.n26 VTAIL.n25 10.4732
R272 VTAIL.n110 VTAIL.n109 10.4732
R273 VTAIL.n70 VTAIL.n69 10.4732
R274 VTAIL.n142 VTAIL.n128 9.69747
R275 VTAIL.n22 VTAIL.n8 9.69747
R276 VTAIL.n106 VTAIL.n92 9.69747
R277 VTAIL.n66 VTAIL.n52 9.69747
R278 VTAIL.n156 VTAIL.n155 9.45567
R279 VTAIL.n36 VTAIL.n35 9.45567
R280 VTAIL.n120 VTAIL.n119 9.45567
R281 VTAIL.n80 VTAIL.n79 9.45567
R282 VTAIL.n132 VTAIL.n131 9.3005
R283 VTAIL.n139 VTAIL.n138 9.3005
R284 VTAIL.n141 VTAIL.n140 9.3005
R285 VTAIL.n128 VTAIL.n127 9.3005
R286 VTAIL.n147 VTAIL.n146 9.3005
R287 VTAIL.n149 VTAIL.n148 9.3005
R288 VTAIL.n124 VTAIL.n123 9.3005
R289 VTAIL.n155 VTAIL.n154 9.3005
R290 VTAIL.n12 VTAIL.n11 9.3005
R291 VTAIL.n19 VTAIL.n18 9.3005
R292 VTAIL.n21 VTAIL.n20 9.3005
R293 VTAIL.n8 VTAIL.n7 9.3005
R294 VTAIL.n27 VTAIL.n26 9.3005
R295 VTAIL.n29 VTAIL.n28 9.3005
R296 VTAIL.n4 VTAIL.n3 9.3005
R297 VTAIL.n35 VTAIL.n34 9.3005
R298 VTAIL.n96 VTAIL.n95 9.3005
R299 VTAIL.n103 VTAIL.n102 9.3005
R300 VTAIL.n105 VTAIL.n104 9.3005
R301 VTAIL.n92 VTAIL.n91 9.3005
R302 VTAIL.n111 VTAIL.n110 9.3005
R303 VTAIL.n113 VTAIL.n112 9.3005
R304 VTAIL.n88 VTAIL.n87 9.3005
R305 VTAIL.n119 VTAIL.n118 9.3005
R306 VTAIL.n56 VTAIL.n55 9.3005
R307 VTAIL.n63 VTAIL.n62 9.3005
R308 VTAIL.n65 VTAIL.n64 9.3005
R309 VTAIL.n52 VTAIL.n51 9.3005
R310 VTAIL.n71 VTAIL.n70 9.3005
R311 VTAIL.n73 VTAIL.n72 9.3005
R312 VTAIL.n48 VTAIL.n47 9.3005
R313 VTAIL.n79 VTAIL.n78 9.3005
R314 VTAIL.n141 VTAIL.n130 8.92171
R315 VTAIL.n21 VTAIL.n10 8.92171
R316 VTAIL.n105 VTAIL.n94 8.92171
R317 VTAIL.n65 VTAIL.n54 8.92171
R318 VTAIL.n138 VTAIL.n137 8.14595
R319 VTAIL.n18 VTAIL.n17 8.14595
R320 VTAIL.n102 VTAIL.n101 8.14595
R321 VTAIL.n62 VTAIL.n61 8.14595
R322 VTAIL.n156 VTAIL.n122 7.75445
R323 VTAIL.n36 VTAIL.n2 7.75445
R324 VTAIL.n120 VTAIL.n86 7.75445
R325 VTAIL.n80 VTAIL.n46 7.75445
R326 VTAIL.n134 VTAIL.n132 7.3702
R327 VTAIL.n14 VTAIL.n12 7.3702
R328 VTAIL.n98 VTAIL.n96 7.3702
R329 VTAIL.n58 VTAIL.n56 7.3702
R330 VTAIL.n154 VTAIL.n122 6.08283
R331 VTAIL.n34 VTAIL.n2 6.08283
R332 VTAIL.n118 VTAIL.n86 6.08283
R333 VTAIL.n78 VTAIL.n46 6.08283
R334 VTAIL.n137 VTAIL.n132 5.81868
R335 VTAIL.n17 VTAIL.n12 5.81868
R336 VTAIL.n101 VTAIL.n96 5.81868
R337 VTAIL.n61 VTAIL.n56 5.81868
R338 VTAIL.n138 VTAIL.n130 5.04292
R339 VTAIL.n18 VTAIL.n10 5.04292
R340 VTAIL.n102 VTAIL.n94 5.04292
R341 VTAIL.n62 VTAIL.n54 5.04292
R342 VTAIL.n158 VTAIL.t10 4.46547
R343 VTAIL.n158 VTAIL.t19 4.46547
R344 VTAIL.n0 VTAIL.t15 4.46547
R345 VTAIL.n0 VTAIL.t17 4.46547
R346 VTAIL.n38 VTAIL.t2 4.46547
R347 VTAIL.n38 VTAIL.t1 4.46547
R348 VTAIL.n40 VTAIL.t0 4.46547
R349 VTAIL.n40 VTAIL.t5 4.46547
R350 VTAIL.n84 VTAIL.t8 4.46547
R351 VTAIL.n84 VTAIL.t4 4.46547
R352 VTAIL.n82 VTAIL.t7 4.46547
R353 VTAIL.n82 VTAIL.t9 4.46547
R354 VTAIL.n44 VTAIL.t14 4.46547
R355 VTAIL.n44 VTAIL.t13 4.46547
R356 VTAIL.n42 VTAIL.t18 4.46547
R357 VTAIL.n42 VTAIL.t16 4.46547
R358 VTAIL.n142 VTAIL.n141 4.26717
R359 VTAIL.n22 VTAIL.n21 4.26717
R360 VTAIL.n106 VTAIL.n105 4.26717
R361 VTAIL.n66 VTAIL.n65 4.26717
R362 VTAIL.n145 VTAIL.n128 3.49141
R363 VTAIL.n25 VTAIL.n8 3.49141
R364 VTAIL.n109 VTAIL.n92 3.49141
R365 VTAIL.n69 VTAIL.n52 3.49141
R366 VTAIL.n45 VTAIL.n43 3.37981
R367 VTAIL.n81 VTAIL.n45 3.37981
R368 VTAIL.n85 VTAIL.n83 3.37981
R369 VTAIL.n121 VTAIL.n85 3.37981
R370 VTAIL.n41 VTAIL.n39 3.37981
R371 VTAIL.n39 VTAIL.n37 3.37981
R372 VTAIL.n159 VTAIL.n157 3.37981
R373 VTAIL.n146 VTAIL.n126 2.71565
R374 VTAIL.n26 VTAIL.n6 2.71565
R375 VTAIL.n110 VTAIL.n90 2.71565
R376 VTAIL.n70 VTAIL.n50 2.71565
R377 VTAIL VTAIL.n1 2.59317
R378 VTAIL.n133 VTAIL.n131 2.41305
R379 VTAIL.n13 VTAIL.n11 2.41305
R380 VTAIL.n97 VTAIL.n95 2.41305
R381 VTAIL.n57 VTAIL.n55 2.41305
R382 VTAIL.n83 VTAIL.n81 2.15998
R383 VTAIL.n37 VTAIL.n1 2.15998
R384 VTAIL.n150 VTAIL.n149 1.93989
R385 VTAIL.n30 VTAIL.n29 1.93989
R386 VTAIL.n114 VTAIL.n113 1.93989
R387 VTAIL.n74 VTAIL.n73 1.93989
R388 VTAIL.n153 VTAIL.n124 1.16414
R389 VTAIL.n33 VTAIL.n4 1.16414
R390 VTAIL.n117 VTAIL.n88 1.16414
R391 VTAIL.n77 VTAIL.n48 1.16414
R392 VTAIL VTAIL.n159 0.787138
R393 VTAIL.n139 VTAIL.n131 0.155672
R394 VTAIL.n140 VTAIL.n139 0.155672
R395 VTAIL.n140 VTAIL.n127 0.155672
R396 VTAIL.n147 VTAIL.n127 0.155672
R397 VTAIL.n148 VTAIL.n147 0.155672
R398 VTAIL.n148 VTAIL.n123 0.155672
R399 VTAIL.n155 VTAIL.n123 0.155672
R400 VTAIL.n19 VTAIL.n11 0.155672
R401 VTAIL.n20 VTAIL.n19 0.155672
R402 VTAIL.n20 VTAIL.n7 0.155672
R403 VTAIL.n27 VTAIL.n7 0.155672
R404 VTAIL.n28 VTAIL.n27 0.155672
R405 VTAIL.n28 VTAIL.n3 0.155672
R406 VTAIL.n35 VTAIL.n3 0.155672
R407 VTAIL.n119 VTAIL.n87 0.155672
R408 VTAIL.n112 VTAIL.n87 0.155672
R409 VTAIL.n112 VTAIL.n111 0.155672
R410 VTAIL.n111 VTAIL.n91 0.155672
R411 VTAIL.n104 VTAIL.n91 0.155672
R412 VTAIL.n104 VTAIL.n103 0.155672
R413 VTAIL.n103 VTAIL.n95 0.155672
R414 VTAIL.n79 VTAIL.n47 0.155672
R415 VTAIL.n72 VTAIL.n47 0.155672
R416 VTAIL.n72 VTAIL.n71 0.155672
R417 VTAIL.n71 VTAIL.n51 0.155672
R418 VTAIL.n64 VTAIL.n51 0.155672
R419 VTAIL.n64 VTAIL.n63 0.155672
R420 VTAIL.n63 VTAIL.n55 0.155672
R421 VDD2.n70 VDD2.n69 585
R422 VDD2.n68 VDD2.n67 585
R423 VDD2.n43 VDD2.n42 585
R424 VDD2.n62 VDD2.n61 585
R425 VDD2.n60 VDD2.n59 585
R426 VDD2.n47 VDD2.n46 585
R427 VDD2.n54 VDD2.n53 585
R428 VDD2.n52 VDD2.n51 585
R429 VDD2.n13 VDD2.n12 585
R430 VDD2.n15 VDD2.n14 585
R431 VDD2.n8 VDD2.n7 585
R432 VDD2.n21 VDD2.n20 585
R433 VDD2.n23 VDD2.n22 585
R434 VDD2.n4 VDD2.n3 585
R435 VDD2.n29 VDD2.n28 585
R436 VDD2.n31 VDD2.n30 585
R437 VDD2.n69 VDD2.n39 498.474
R438 VDD2.n30 VDD2.n0 498.474
R439 VDD2.n50 VDD2.t8 329.053
R440 VDD2.n11 VDD2.t4 329.053
R441 VDD2.n69 VDD2.n68 171.744
R442 VDD2.n68 VDD2.n42 171.744
R443 VDD2.n61 VDD2.n42 171.744
R444 VDD2.n61 VDD2.n60 171.744
R445 VDD2.n60 VDD2.n46 171.744
R446 VDD2.n53 VDD2.n46 171.744
R447 VDD2.n53 VDD2.n52 171.744
R448 VDD2.n14 VDD2.n13 171.744
R449 VDD2.n14 VDD2.n7 171.744
R450 VDD2.n21 VDD2.n7 171.744
R451 VDD2.n22 VDD2.n21 171.744
R452 VDD2.n22 VDD2.n3 171.744
R453 VDD2.n29 VDD2.n3 171.744
R454 VDD2.n30 VDD2.n29 171.744
R455 VDD2.n38 VDD2.n37 91.1966
R456 VDD2 VDD2.n77 91.1938
R457 VDD2.n76 VDD2.n75 88.7176
R458 VDD2.n36 VDD2.n35 88.7175
R459 VDD2.n52 VDD2.t8 85.8723
R460 VDD2.n13 VDD2.t4 85.8723
R461 VDD2.n36 VDD2.n34 56.1222
R462 VDD2.n74 VDD2.n73 52.7429
R463 VDD2.n74 VDD2.n38 46.0429
R464 VDD2.n71 VDD2.n70 12.8005
R465 VDD2.n32 VDD2.n31 12.8005
R466 VDD2.n67 VDD2.n41 12.0247
R467 VDD2.n28 VDD2.n2 12.0247
R468 VDD2.n66 VDD2.n43 11.249
R469 VDD2.n27 VDD2.n4 11.249
R470 VDD2.n51 VDD2.n50 10.7237
R471 VDD2.n12 VDD2.n11 10.7237
R472 VDD2.n63 VDD2.n62 10.4732
R473 VDD2.n24 VDD2.n23 10.4732
R474 VDD2.n59 VDD2.n45 9.69747
R475 VDD2.n20 VDD2.n6 9.69747
R476 VDD2.n73 VDD2.n72 9.45567
R477 VDD2.n34 VDD2.n33 9.45567
R478 VDD2.n49 VDD2.n48 9.3005
R479 VDD2.n56 VDD2.n55 9.3005
R480 VDD2.n58 VDD2.n57 9.3005
R481 VDD2.n45 VDD2.n44 9.3005
R482 VDD2.n64 VDD2.n63 9.3005
R483 VDD2.n66 VDD2.n65 9.3005
R484 VDD2.n41 VDD2.n40 9.3005
R485 VDD2.n72 VDD2.n71 9.3005
R486 VDD2.n10 VDD2.n9 9.3005
R487 VDD2.n17 VDD2.n16 9.3005
R488 VDD2.n19 VDD2.n18 9.3005
R489 VDD2.n6 VDD2.n5 9.3005
R490 VDD2.n25 VDD2.n24 9.3005
R491 VDD2.n27 VDD2.n26 9.3005
R492 VDD2.n2 VDD2.n1 9.3005
R493 VDD2.n33 VDD2.n32 9.3005
R494 VDD2.n58 VDD2.n47 8.92171
R495 VDD2.n19 VDD2.n8 8.92171
R496 VDD2.n55 VDD2.n54 8.14595
R497 VDD2.n16 VDD2.n15 8.14595
R498 VDD2.n73 VDD2.n39 7.75445
R499 VDD2.n34 VDD2.n0 7.75445
R500 VDD2.n51 VDD2.n49 7.3702
R501 VDD2.n12 VDD2.n10 7.3702
R502 VDD2.n71 VDD2.n39 6.08283
R503 VDD2.n32 VDD2.n0 6.08283
R504 VDD2.n54 VDD2.n49 5.81868
R505 VDD2.n15 VDD2.n10 5.81868
R506 VDD2.n55 VDD2.n47 5.04292
R507 VDD2.n16 VDD2.n8 5.04292
R508 VDD2.n77 VDD2.t5 4.46547
R509 VDD2.n77 VDD2.t3 4.46547
R510 VDD2.n75 VDD2.t2 4.46547
R511 VDD2.n75 VDD2.t7 4.46547
R512 VDD2.n37 VDD2.t6 4.46547
R513 VDD2.n37 VDD2.t1 4.46547
R514 VDD2.n35 VDD2.t0 4.46547
R515 VDD2.n35 VDD2.t9 4.46547
R516 VDD2.n59 VDD2.n58 4.26717
R517 VDD2.n20 VDD2.n19 4.26717
R518 VDD2.n62 VDD2.n45 3.49141
R519 VDD2.n23 VDD2.n6 3.49141
R520 VDD2.n76 VDD2.n74 3.37981
R521 VDD2.n63 VDD2.n43 2.71565
R522 VDD2.n24 VDD2.n4 2.71565
R523 VDD2.n50 VDD2.n48 2.41305
R524 VDD2.n11 VDD2.n9 2.41305
R525 VDD2.n67 VDD2.n66 1.93989
R526 VDD2.n28 VDD2.n27 1.93989
R527 VDD2.n70 VDD2.n41 1.16414
R528 VDD2.n31 VDD2.n2 1.16414
R529 VDD2 VDD2.n76 0.903517
R530 VDD2.n38 VDD2.n36 0.789982
R531 VDD2.n72 VDD2.n40 0.155672
R532 VDD2.n65 VDD2.n40 0.155672
R533 VDD2.n65 VDD2.n64 0.155672
R534 VDD2.n64 VDD2.n44 0.155672
R535 VDD2.n57 VDD2.n44 0.155672
R536 VDD2.n57 VDD2.n56 0.155672
R537 VDD2.n56 VDD2.n48 0.155672
R538 VDD2.n17 VDD2.n9 0.155672
R539 VDD2.n18 VDD2.n17 0.155672
R540 VDD2.n18 VDD2.n5 0.155672
R541 VDD2.n25 VDD2.n5 0.155672
R542 VDD2.n26 VDD2.n25 0.155672
R543 VDD2.n26 VDD2.n1 0.155672
R544 VDD2.n33 VDD2.n1 0.155672
R545 VP.n32 VP.n29 161.3
R546 VP.n34 VP.n33 161.3
R547 VP.n35 VP.n28 161.3
R548 VP.n37 VP.n36 161.3
R549 VP.n38 VP.n27 161.3
R550 VP.n40 VP.n39 161.3
R551 VP.n41 VP.n26 161.3
R552 VP.n44 VP.n43 161.3
R553 VP.n45 VP.n25 161.3
R554 VP.n47 VP.n46 161.3
R555 VP.n48 VP.n24 161.3
R556 VP.n50 VP.n49 161.3
R557 VP.n51 VP.n23 161.3
R558 VP.n53 VP.n52 161.3
R559 VP.n54 VP.n22 161.3
R560 VP.n57 VP.n56 161.3
R561 VP.n58 VP.n21 161.3
R562 VP.n60 VP.n59 161.3
R563 VP.n61 VP.n20 161.3
R564 VP.n63 VP.n62 161.3
R565 VP.n64 VP.n19 161.3
R566 VP.n66 VP.n65 161.3
R567 VP.n67 VP.n18 161.3
R568 VP.n69 VP.n68 161.3
R569 VP.n123 VP.n122 161.3
R570 VP.n121 VP.n1 161.3
R571 VP.n120 VP.n119 161.3
R572 VP.n118 VP.n2 161.3
R573 VP.n117 VP.n116 161.3
R574 VP.n115 VP.n3 161.3
R575 VP.n114 VP.n113 161.3
R576 VP.n112 VP.n4 161.3
R577 VP.n111 VP.n110 161.3
R578 VP.n108 VP.n5 161.3
R579 VP.n107 VP.n106 161.3
R580 VP.n105 VP.n6 161.3
R581 VP.n104 VP.n103 161.3
R582 VP.n102 VP.n7 161.3
R583 VP.n101 VP.n100 161.3
R584 VP.n99 VP.n8 161.3
R585 VP.n98 VP.n97 161.3
R586 VP.n95 VP.n9 161.3
R587 VP.n94 VP.n93 161.3
R588 VP.n92 VP.n10 161.3
R589 VP.n91 VP.n90 161.3
R590 VP.n89 VP.n11 161.3
R591 VP.n88 VP.n87 161.3
R592 VP.n86 VP.n12 161.3
R593 VP.n85 VP.n84 161.3
R594 VP.n82 VP.n13 161.3
R595 VP.n81 VP.n80 161.3
R596 VP.n79 VP.n14 161.3
R597 VP.n78 VP.n77 161.3
R598 VP.n76 VP.n15 161.3
R599 VP.n75 VP.n74 161.3
R600 VP.n73 VP.n16 161.3
R601 VP.n72 VP.n71 85.819
R602 VP.n124 VP.n0 85.819
R603 VP.n70 VP.n17 85.819
R604 VP.n31 VP.t4 81.2363
R605 VP.n31 VP.n30 66.4721
R606 VP.n90 VP.n10 56.5617
R607 VP.n103 VP.n6 56.5617
R608 VP.n49 VP.n23 56.5617
R609 VP.n36 VP.n27 56.5617
R610 VP.n72 VP.n70 54.9465
R611 VP.n77 VP.n14 53.171
R612 VP.n116 VP.n2 53.171
R613 VP.n62 VP.n19 53.171
R614 VP.n71 VP.t5 48.8718
R615 VP.n83 VP.t0 48.8718
R616 VP.n96 VP.t9 48.8718
R617 VP.n109 VP.t8 48.8718
R618 VP.n0 VP.t3 48.8718
R619 VP.n17 VP.t7 48.8718
R620 VP.n55 VP.t2 48.8718
R621 VP.n42 VP.t6 48.8718
R622 VP.n30 VP.t1 48.8718
R623 VP.n81 VP.n14 27.983
R624 VP.n116 VP.n115 27.983
R625 VP.n62 VP.n61 27.983
R626 VP.n75 VP.n16 24.5923
R627 VP.n76 VP.n75 24.5923
R628 VP.n77 VP.n76 24.5923
R629 VP.n82 VP.n81 24.5923
R630 VP.n84 VP.n82 24.5923
R631 VP.n88 VP.n12 24.5923
R632 VP.n89 VP.n88 24.5923
R633 VP.n90 VP.n89 24.5923
R634 VP.n94 VP.n10 24.5923
R635 VP.n95 VP.n94 24.5923
R636 VP.n97 VP.n95 24.5923
R637 VP.n101 VP.n8 24.5923
R638 VP.n102 VP.n101 24.5923
R639 VP.n103 VP.n102 24.5923
R640 VP.n107 VP.n6 24.5923
R641 VP.n108 VP.n107 24.5923
R642 VP.n110 VP.n108 24.5923
R643 VP.n114 VP.n4 24.5923
R644 VP.n115 VP.n114 24.5923
R645 VP.n120 VP.n2 24.5923
R646 VP.n121 VP.n120 24.5923
R647 VP.n122 VP.n121 24.5923
R648 VP.n66 VP.n19 24.5923
R649 VP.n67 VP.n66 24.5923
R650 VP.n68 VP.n67 24.5923
R651 VP.n53 VP.n23 24.5923
R652 VP.n54 VP.n53 24.5923
R653 VP.n56 VP.n54 24.5923
R654 VP.n60 VP.n21 24.5923
R655 VP.n61 VP.n60 24.5923
R656 VP.n40 VP.n27 24.5923
R657 VP.n41 VP.n40 24.5923
R658 VP.n43 VP.n41 24.5923
R659 VP.n47 VP.n25 24.5923
R660 VP.n48 VP.n47 24.5923
R661 VP.n49 VP.n48 24.5923
R662 VP.n34 VP.n29 24.5923
R663 VP.n35 VP.n34 24.5923
R664 VP.n36 VP.n35 24.5923
R665 VP.n84 VP.n83 16.2311
R666 VP.n109 VP.n4 16.2311
R667 VP.n55 VP.n21 16.2311
R668 VP.n97 VP.n96 12.2964
R669 VP.n96 VP.n8 12.2964
R670 VP.n43 VP.n42 12.2964
R671 VP.n42 VP.n25 12.2964
R672 VP.n83 VP.n12 8.36172
R673 VP.n110 VP.n109 8.36172
R674 VP.n56 VP.n55 8.36172
R675 VP.n30 VP.n29 8.36172
R676 VP.n71 VP.n16 4.42703
R677 VP.n122 VP.n0 4.42703
R678 VP.n68 VP.n17 4.42703
R679 VP.n32 VP.n31 3.3215
R680 VP.n70 VP.n69 0.354861
R681 VP.n73 VP.n72 0.354861
R682 VP.n124 VP.n123 0.354861
R683 VP VP.n124 0.267071
R684 VP.n33 VP.n32 0.189894
R685 VP.n33 VP.n28 0.189894
R686 VP.n37 VP.n28 0.189894
R687 VP.n38 VP.n37 0.189894
R688 VP.n39 VP.n38 0.189894
R689 VP.n39 VP.n26 0.189894
R690 VP.n44 VP.n26 0.189894
R691 VP.n45 VP.n44 0.189894
R692 VP.n46 VP.n45 0.189894
R693 VP.n46 VP.n24 0.189894
R694 VP.n50 VP.n24 0.189894
R695 VP.n51 VP.n50 0.189894
R696 VP.n52 VP.n51 0.189894
R697 VP.n52 VP.n22 0.189894
R698 VP.n57 VP.n22 0.189894
R699 VP.n58 VP.n57 0.189894
R700 VP.n59 VP.n58 0.189894
R701 VP.n59 VP.n20 0.189894
R702 VP.n63 VP.n20 0.189894
R703 VP.n64 VP.n63 0.189894
R704 VP.n65 VP.n64 0.189894
R705 VP.n65 VP.n18 0.189894
R706 VP.n69 VP.n18 0.189894
R707 VP.n74 VP.n73 0.189894
R708 VP.n74 VP.n15 0.189894
R709 VP.n78 VP.n15 0.189894
R710 VP.n79 VP.n78 0.189894
R711 VP.n80 VP.n79 0.189894
R712 VP.n80 VP.n13 0.189894
R713 VP.n85 VP.n13 0.189894
R714 VP.n86 VP.n85 0.189894
R715 VP.n87 VP.n86 0.189894
R716 VP.n87 VP.n11 0.189894
R717 VP.n91 VP.n11 0.189894
R718 VP.n92 VP.n91 0.189894
R719 VP.n93 VP.n92 0.189894
R720 VP.n93 VP.n9 0.189894
R721 VP.n98 VP.n9 0.189894
R722 VP.n99 VP.n98 0.189894
R723 VP.n100 VP.n99 0.189894
R724 VP.n100 VP.n7 0.189894
R725 VP.n104 VP.n7 0.189894
R726 VP.n105 VP.n104 0.189894
R727 VP.n106 VP.n105 0.189894
R728 VP.n106 VP.n5 0.189894
R729 VP.n111 VP.n5 0.189894
R730 VP.n112 VP.n111 0.189894
R731 VP.n113 VP.n112 0.189894
R732 VP.n113 VP.n3 0.189894
R733 VP.n117 VP.n3 0.189894
R734 VP.n118 VP.n117 0.189894
R735 VP.n119 VP.n118 0.189894
R736 VP.n119 VP.n1 0.189894
R737 VP.n123 VP.n1 0.189894
R738 VDD1.n31 VDD1.n30 585
R739 VDD1.n29 VDD1.n28 585
R740 VDD1.n4 VDD1.n3 585
R741 VDD1.n23 VDD1.n22 585
R742 VDD1.n21 VDD1.n20 585
R743 VDD1.n8 VDD1.n7 585
R744 VDD1.n15 VDD1.n14 585
R745 VDD1.n13 VDD1.n12 585
R746 VDD1.n50 VDD1.n49 585
R747 VDD1.n52 VDD1.n51 585
R748 VDD1.n45 VDD1.n44 585
R749 VDD1.n58 VDD1.n57 585
R750 VDD1.n60 VDD1.n59 585
R751 VDD1.n41 VDD1.n40 585
R752 VDD1.n66 VDD1.n65 585
R753 VDD1.n68 VDD1.n67 585
R754 VDD1.n30 VDD1.n0 498.474
R755 VDD1.n67 VDD1.n37 498.474
R756 VDD1.n11 VDD1.t5 329.053
R757 VDD1.n48 VDD1.t4 329.053
R758 VDD1.n30 VDD1.n29 171.744
R759 VDD1.n29 VDD1.n3 171.744
R760 VDD1.n22 VDD1.n3 171.744
R761 VDD1.n22 VDD1.n21 171.744
R762 VDD1.n21 VDD1.n7 171.744
R763 VDD1.n14 VDD1.n7 171.744
R764 VDD1.n14 VDD1.n13 171.744
R765 VDD1.n51 VDD1.n50 171.744
R766 VDD1.n51 VDD1.n44 171.744
R767 VDD1.n58 VDD1.n44 171.744
R768 VDD1.n59 VDD1.n58 171.744
R769 VDD1.n59 VDD1.n40 171.744
R770 VDD1.n66 VDD1.n40 171.744
R771 VDD1.n67 VDD1.n66 171.744
R772 VDD1.n75 VDD1.n74 91.1966
R773 VDD1.n36 VDD1.n35 88.7176
R774 VDD1.n77 VDD1.n76 88.7175
R775 VDD1.n73 VDD1.n72 88.7175
R776 VDD1.n13 VDD1.t5 85.8723
R777 VDD1.n50 VDD1.t4 85.8723
R778 VDD1.n36 VDD1.n34 56.1222
R779 VDD1.n73 VDD1.n71 56.1222
R780 VDD1.n77 VDD1.n75 48.3155
R781 VDD1.n32 VDD1.n31 12.8005
R782 VDD1.n69 VDD1.n68 12.8005
R783 VDD1.n28 VDD1.n2 12.0247
R784 VDD1.n65 VDD1.n39 12.0247
R785 VDD1.n27 VDD1.n4 11.249
R786 VDD1.n64 VDD1.n41 11.249
R787 VDD1.n12 VDD1.n11 10.7237
R788 VDD1.n49 VDD1.n48 10.7237
R789 VDD1.n24 VDD1.n23 10.4732
R790 VDD1.n61 VDD1.n60 10.4732
R791 VDD1.n20 VDD1.n6 9.69747
R792 VDD1.n57 VDD1.n43 9.69747
R793 VDD1.n34 VDD1.n33 9.45567
R794 VDD1.n71 VDD1.n70 9.45567
R795 VDD1.n10 VDD1.n9 9.3005
R796 VDD1.n17 VDD1.n16 9.3005
R797 VDD1.n19 VDD1.n18 9.3005
R798 VDD1.n6 VDD1.n5 9.3005
R799 VDD1.n25 VDD1.n24 9.3005
R800 VDD1.n27 VDD1.n26 9.3005
R801 VDD1.n2 VDD1.n1 9.3005
R802 VDD1.n33 VDD1.n32 9.3005
R803 VDD1.n47 VDD1.n46 9.3005
R804 VDD1.n54 VDD1.n53 9.3005
R805 VDD1.n56 VDD1.n55 9.3005
R806 VDD1.n43 VDD1.n42 9.3005
R807 VDD1.n62 VDD1.n61 9.3005
R808 VDD1.n64 VDD1.n63 9.3005
R809 VDD1.n39 VDD1.n38 9.3005
R810 VDD1.n70 VDD1.n69 9.3005
R811 VDD1.n19 VDD1.n8 8.92171
R812 VDD1.n56 VDD1.n45 8.92171
R813 VDD1.n16 VDD1.n15 8.14595
R814 VDD1.n53 VDD1.n52 8.14595
R815 VDD1.n34 VDD1.n0 7.75445
R816 VDD1.n71 VDD1.n37 7.75445
R817 VDD1.n12 VDD1.n10 7.3702
R818 VDD1.n49 VDD1.n47 7.3702
R819 VDD1.n32 VDD1.n0 6.08283
R820 VDD1.n69 VDD1.n37 6.08283
R821 VDD1.n15 VDD1.n10 5.81868
R822 VDD1.n52 VDD1.n47 5.81868
R823 VDD1.n16 VDD1.n8 5.04292
R824 VDD1.n53 VDD1.n45 5.04292
R825 VDD1.n76 VDD1.t7 4.46547
R826 VDD1.n76 VDD1.t2 4.46547
R827 VDD1.n35 VDD1.t8 4.46547
R828 VDD1.n35 VDD1.t3 4.46547
R829 VDD1.n74 VDD1.t1 4.46547
R830 VDD1.n74 VDD1.t6 4.46547
R831 VDD1.n72 VDD1.t9 4.46547
R832 VDD1.n72 VDD1.t0 4.46547
R833 VDD1.n20 VDD1.n19 4.26717
R834 VDD1.n57 VDD1.n56 4.26717
R835 VDD1.n23 VDD1.n6 3.49141
R836 VDD1.n60 VDD1.n43 3.49141
R837 VDD1.n24 VDD1.n4 2.71565
R838 VDD1.n61 VDD1.n41 2.71565
R839 VDD1 VDD1.n77 2.47679
R840 VDD1.n11 VDD1.n9 2.41305
R841 VDD1.n48 VDD1.n46 2.41305
R842 VDD1.n28 VDD1.n27 1.93989
R843 VDD1.n65 VDD1.n64 1.93989
R844 VDD1.n31 VDD1.n2 1.16414
R845 VDD1.n68 VDD1.n39 1.16414
R846 VDD1 VDD1.n36 0.903517
R847 VDD1.n75 VDD1.n73 0.789982
R848 VDD1.n33 VDD1.n1 0.155672
R849 VDD1.n26 VDD1.n1 0.155672
R850 VDD1.n26 VDD1.n25 0.155672
R851 VDD1.n25 VDD1.n5 0.155672
R852 VDD1.n18 VDD1.n5 0.155672
R853 VDD1.n18 VDD1.n17 0.155672
R854 VDD1.n17 VDD1.n9 0.155672
R855 VDD1.n54 VDD1.n46 0.155672
R856 VDD1.n55 VDD1.n54 0.155672
R857 VDD1.n55 VDD1.n42 0.155672
R858 VDD1.n62 VDD1.n42 0.155672
R859 VDD1.n63 VDD1.n62 0.155672
R860 VDD1.n63 VDD1.n38 0.155672
R861 VDD1.n70 VDD1.n38 0.155672
R862 B.n443 B.n156 585
R863 B.n442 B.n441 585
R864 B.n440 B.n157 585
R865 B.n439 B.n438 585
R866 B.n437 B.n158 585
R867 B.n436 B.n435 585
R868 B.n434 B.n159 585
R869 B.n433 B.n432 585
R870 B.n431 B.n160 585
R871 B.n430 B.n429 585
R872 B.n428 B.n161 585
R873 B.n427 B.n426 585
R874 B.n425 B.n162 585
R875 B.n424 B.n423 585
R876 B.n422 B.n163 585
R877 B.n421 B.n420 585
R878 B.n419 B.n164 585
R879 B.n418 B.n417 585
R880 B.n416 B.n165 585
R881 B.n415 B.n414 585
R882 B.n413 B.n166 585
R883 B.n412 B.n411 585
R884 B.n410 B.n167 585
R885 B.n409 B.n408 585
R886 B.n407 B.n168 585
R887 B.n406 B.n405 585
R888 B.n404 B.n169 585
R889 B.n403 B.n402 585
R890 B.n400 B.n170 585
R891 B.n399 B.n398 585
R892 B.n397 B.n173 585
R893 B.n396 B.n395 585
R894 B.n394 B.n174 585
R895 B.n393 B.n392 585
R896 B.n391 B.n175 585
R897 B.n390 B.n389 585
R898 B.n388 B.n176 585
R899 B.n386 B.n385 585
R900 B.n384 B.n179 585
R901 B.n383 B.n382 585
R902 B.n381 B.n180 585
R903 B.n380 B.n379 585
R904 B.n378 B.n181 585
R905 B.n377 B.n376 585
R906 B.n375 B.n182 585
R907 B.n374 B.n373 585
R908 B.n372 B.n183 585
R909 B.n371 B.n370 585
R910 B.n369 B.n184 585
R911 B.n368 B.n367 585
R912 B.n366 B.n185 585
R913 B.n365 B.n364 585
R914 B.n363 B.n186 585
R915 B.n362 B.n361 585
R916 B.n360 B.n187 585
R917 B.n359 B.n358 585
R918 B.n357 B.n188 585
R919 B.n356 B.n355 585
R920 B.n354 B.n189 585
R921 B.n353 B.n352 585
R922 B.n351 B.n190 585
R923 B.n350 B.n349 585
R924 B.n348 B.n191 585
R925 B.n347 B.n346 585
R926 B.n345 B.n192 585
R927 B.n445 B.n444 585
R928 B.n446 B.n155 585
R929 B.n448 B.n447 585
R930 B.n449 B.n154 585
R931 B.n451 B.n450 585
R932 B.n452 B.n153 585
R933 B.n454 B.n453 585
R934 B.n455 B.n152 585
R935 B.n457 B.n456 585
R936 B.n458 B.n151 585
R937 B.n460 B.n459 585
R938 B.n461 B.n150 585
R939 B.n463 B.n462 585
R940 B.n464 B.n149 585
R941 B.n466 B.n465 585
R942 B.n467 B.n148 585
R943 B.n469 B.n468 585
R944 B.n470 B.n147 585
R945 B.n472 B.n471 585
R946 B.n473 B.n146 585
R947 B.n475 B.n474 585
R948 B.n476 B.n145 585
R949 B.n478 B.n477 585
R950 B.n479 B.n144 585
R951 B.n481 B.n480 585
R952 B.n482 B.n143 585
R953 B.n484 B.n483 585
R954 B.n485 B.n142 585
R955 B.n487 B.n486 585
R956 B.n488 B.n141 585
R957 B.n490 B.n489 585
R958 B.n491 B.n140 585
R959 B.n493 B.n492 585
R960 B.n494 B.n139 585
R961 B.n496 B.n495 585
R962 B.n497 B.n138 585
R963 B.n499 B.n498 585
R964 B.n500 B.n137 585
R965 B.n502 B.n501 585
R966 B.n503 B.n136 585
R967 B.n505 B.n504 585
R968 B.n506 B.n135 585
R969 B.n508 B.n507 585
R970 B.n509 B.n134 585
R971 B.n511 B.n510 585
R972 B.n512 B.n133 585
R973 B.n514 B.n513 585
R974 B.n515 B.n132 585
R975 B.n517 B.n516 585
R976 B.n518 B.n131 585
R977 B.n520 B.n519 585
R978 B.n521 B.n130 585
R979 B.n523 B.n522 585
R980 B.n524 B.n129 585
R981 B.n526 B.n525 585
R982 B.n527 B.n128 585
R983 B.n529 B.n528 585
R984 B.n530 B.n127 585
R985 B.n532 B.n531 585
R986 B.n533 B.n126 585
R987 B.n535 B.n534 585
R988 B.n536 B.n125 585
R989 B.n538 B.n537 585
R990 B.n539 B.n124 585
R991 B.n541 B.n540 585
R992 B.n542 B.n123 585
R993 B.n544 B.n543 585
R994 B.n545 B.n122 585
R995 B.n547 B.n546 585
R996 B.n548 B.n121 585
R997 B.n550 B.n549 585
R998 B.n551 B.n120 585
R999 B.n553 B.n552 585
R1000 B.n554 B.n119 585
R1001 B.n556 B.n555 585
R1002 B.n557 B.n118 585
R1003 B.n559 B.n558 585
R1004 B.n560 B.n117 585
R1005 B.n562 B.n561 585
R1006 B.n563 B.n116 585
R1007 B.n565 B.n564 585
R1008 B.n566 B.n115 585
R1009 B.n568 B.n567 585
R1010 B.n569 B.n114 585
R1011 B.n571 B.n570 585
R1012 B.n572 B.n113 585
R1013 B.n574 B.n573 585
R1014 B.n575 B.n112 585
R1015 B.n577 B.n576 585
R1016 B.n578 B.n111 585
R1017 B.n580 B.n579 585
R1018 B.n581 B.n110 585
R1019 B.n583 B.n582 585
R1020 B.n584 B.n109 585
R1021 B.n586 B.n585 585
R1022 B.n587 B.n108 585
R1023 B.n589 B.n588 585
R1024 B.n590 B.n107 585
R1025 B.n592 B.n591 585
R1026 B.n593 B.n106 585
R1027 B.n595 B.n594 585
R1028 B.n596 B.n105 585
R1029 B.n598 B.n597 585
R1030 B.n599 B.n104 585
R1031 B.n601 B.n600 585
R1032 B.n602 B.n103 585
R1033 B.n604 B.n603 585
R1034 B.n605 B.n102 585
R1035 B.n607 B.n606 585
R1036 B.n608 B.n101 585
R1037 B.n610 B.n609 585
R1038 B.n611 B.n100 585
R1039 B.n613 B.n612 585
R1040 B.n614 B.n99 585
R1041 B.n616 B.n615 585
R1042 B.n617 B.n98 585
R1043 B.n619 B.n618 585
R1044 B.n620 B.n97 585
R1045 B.n622 B.n621 585
R1046 B.n623 B.n96 585
R1047 B.n625 B.n624 585
R1048 B.n626 B.n95 585
R1049 B.n628 B.n627 585
R1050 B.n629 B.n94 585
R1051 B.n631 B.n630 585
R1052 B.n632 B.n93 585
R1053 B.n634 B.n633 585
R1054 B.n635 B.n92 585
R1055 B.n637 B.n636 585
R1056 B.n638 B.n91 585
R1057 B.n640 B.n639 585
R1058 B.n641 B.n90 585
R1059 B.n643 B.n642 585
R1060 B.n644 B.n89 585
R1061 B.n646 B.n645 585
R1062 B.n647 B.n88 585
R1063 B.n649 B.n648 585
R1064 B.n650 B.n87 585
R1065 B.n652 B.n651 585
R1066 B.n653 B.n86 585
R1067 B.n655 B.n654 585
R1068 B.n656 B.n85 585
R1069 B.n658 B.n657 585
R1070 B.n659 B.n84 585
R1071 B.n661 B.n660 585
R1072 B.n662 B.n83 585
R1073 B.n664 B.n663 585
R1074 B.n665 B.n82 585
R1075 B.n667 B.n666 585
R1076 B.n668 B.n81 585
R1077 B.n670 B.n669 585
R1078 B.n671 B.n80 585
R1079 B.n673 B.n672 585
R1080 B.n674 B.n79 585
R1081 B.n676 B.n675 585
R1082 B.n677 B.n78 585
R1083 B.n776 B.n775 585
R1084 B.n774 B.n41 585
R1085 B.n773 B.n772 585
R1086 B.n771 B.n42 585
R1087 B.n770 B.n769 585
R1088 B.n768 B.n43 585
R1089 B.n767 B.n766 585
R1090 B.n765 B.n44 585
R1091 B.n764 B.n763 585
R1092 B.n762 B.n45 585
R1093 B.n761 B.n760 585
R1094 B.n759 B.n46 585
R1095 B.n758 B.n757 585
R1096 B.n756 B.n47 585
R1097 B.n755 B.n754 585
R1098 B.n753 B.n48 585
R1099 B.n752 B.n751 585
R1100 B.n750 B.n49 585
R1101 B.n749 B.n748 585
R1102 B.n747 B.n50 585
R1103 B.n746 B.n745 585
R1104 B.n744 B.n51 585
R1105 B.n743 B.n742 585
R1106 B.n741 B.n52 585
R1107 B.n740 B.n739 585
R1108 B.n738 B.n53 585
R1109 B.n737 B.n736 585
R1110 B.n735 B.n54 585
R1111 B.n734 B.n733 585
R1112 B.n732 B.n55 585
R1113 B.n731 B.n730 585
R1114 B.n729 B.n59 585
R1115 B.n728 B.n727 585
R1116 B.n726 B.n60 585
R1117 B.n725 B.n724 585
R1118 B.n723 B.n61 585
R1119 B.n722 B.n721 585
R1120 B.n719 B.n62 585
R1121 B.n718 B.n717 585
R1122 B.n716 B.n65 585
R1123 B.n715 B.n714 585
R1124 B.n713 B.n66 585
R1125 B.n712 B.n711 585
R1126 B.n710 B.n67 585
R1127 B.n709 B.n708 585
R1128 B.n707 B.n68 585
R1129 B.n706 B.n705 585
R1130 B.n704 B.n69 585
R1131 B.n703 B.n702 585
R1132 B.n701 B.n70 585
R1133 B.n700 B.n699 585
R1134 B.n698 B.n71 585
R1135 B.n697 B.n696 585
R1136 B.n695 B.n72 585
R1137 B.n694 B.n693 585
R1138 B.n692 B.n73 585
R1139 B.n691 B.n690 585
R1140 B.n689 B.n74 585
R1141 B.n688 B.n687 585
R1142 B.n686 B.n75 585
R1143 B.n685 B.n684 585
R1144 B.n683 B.n76 585
R1145 B.n682 B.n681 585
R1146 B.n680 B.n77 585
R1147 B.n679 B.n678 585
R1148 B.n777 B.n40 585
R1149 B.n779 B.n778 585
R1150 B.n780 B.n39 585
R1151 B.n782 B.n781 585
R1152 B.n783 B.n38 585
R1153 B.n785 B.n784 585
R1154 B.n786 B.n37 585
R1155 B.n788 B.n787 585
R1156 B.n789 B.n36 585
R1157 B.n791 B.n790 585
R1158 B.n792 B.n35 585
R1159 B.n794 B.n793 585
R1160 B.n795 B.n34 585
R1161 B.n797 B.n796 585
R1162 B.n798 B.n33 585
R1163 B.n800 B.n799 585
R1164 B.n801 B.n32 585
R1165 B.n803 B.n802 585
R1166 B.n804 B.n31 585
R1167 B.n806 B.n805 585
R1168 B.n807 B.n30 585
R1169 B.n809 B.n808 585
R1170 B.n810 B.n29 585
R1171 B.n812 B.n811 585
R1172 B.n813 B.n28 585
R1173 B.n815 B.n814 585
R1174 B.n816 B.n27 585
R1175 B.n818 B.n817 585
R1176 B.n819 B.n26 585
R1177 B.n821 B.n820 585
R1178 B.n822 B.n25 585
R1179 B.n824 B.n823 585
R1180 B.n825 B.n24 585
R1181 B.n827 B.n826 585
R1182 B.n828 B.n23 585
R1183 B.n830 B.n829 585
R1184 B.n831 B.n22 585
R1185 B.n833 B.n832 585
R1186 B.n834 B.n21 585
R1187 B.n836 B.n835 585
R1188 B.n837 B.n20 585
R1189 B.n839 B.n838 585
R1190 B.n840 B.n19 585
R1191 B.n842 B.n841 585
R1192 B.n843 B.n18 585
R1193 B.n845 B.n844 585
R1194 B.n846 B.n17 585
R1195 B.n848 B.n847 585
R1196 B.n849 B.n16 585
R1197 B.n851 B.n850 585
R1198 B.n852 B.n15 585
R1199 B.n854 B.n853 585
R1200 B.n855 B.n14 585
R1201 B.n857 B.n856 585
R1202 B.n858 B.n13 585
R1203 B.n860 B.n859 585
R1204 B.n861 B.n12 585
R1205 B.n863 B.n862 585
R1206 B.n864 B.n11 585
R1207 B.n866 B.n865 585
R1208 B.n867 B.n10 585
R1209 B.n869 B.n868 585
R1210 B.n870 B.n9 585
R1211 B.n872 B.n871 585
R1212 B.n873 B.n8 585
R1213 B.n875 B.n874 585
R1214 B.n876 B.n7 585
R1215 B.n878 B.n877 585
R1216 B.n879 B.n6 585
R1217 B.n881 B.n880 585
R1218 B.n882 B.n5 585
R1219 B.n884 B.n883 585
R1220 B.n885 B.n4 585
R1221 B.n887 B.n886 585
R1222 B.n888 B.n3 585
R1223 B.n890 B.n889 585
R1224 B.n891 B.n0 585
R1225 B.n2 B.n1 585
R1226 B.n231 B.n230 585
R1227 B.n233 B.n232 585
R1228 B.n234 B.n229 585
R1229 B.n236 B.n235 585
R1230 B.n237 B.n228 585
R1231 B.n239 B.n238 585
R1232 B.n240 B.n227 585
R1233 B.n242 B.n241 585
R1234 B.n243 B.n226 585
R1235 B.n245 B.n244 585
R1236 B.n246 B.n225 585
R1237 B.n248 B.n247 585
R1238 B.n249 B.n224 585
R1239 B.n251 B.n250 585
R1240 B.n252 B.n223 585
R1241 B.n254 B.n253 585
R1242 B.n255 B.n222 585
R1243 B.n257 B.n256 585
R1244 B.n258 B.n221 585
R1245 B.n260 B.n259 585
R1246 B.n261 B.n220 585
R1247 B.n263 B.n262 585
R1248 B.n264 B.n219 585
R1249 B.n266 B.n265 585
R1250 B.n267 B.n218 585
R1251 B.n269 B.n268 585
R1252 B.n270 B.n217 585
R1253 B.n272 B.n271 585
R1254 B.n273 B.n216 585
R1255 B.n275 B.n274 585
R1256 B.n276 B.n215 585
R1257 B.n278 B.n277 585
R1258 B.n279 B.n214 585
R1259 B.n281 B.n280 585
R1260 B.n282 B.n213 585
R1261 B.n284 B.n283 585
R1262 B.n285 B.n212 585
R1263 B.n287 B.n286 585
R1264 B.n288 B.n211 585
R1265 B.n290 B.n289 585
R1266 B.n291 B.n210 585
R1267 B.n293 B.n292 585
R1268 B.n294 B.n209 585
R1269 B.n296 B.n295 585
R1270 B.n297 B.n208 585
R1271 B.n299 B.n298 585
R1272 B.n300 B.n207 585
R1273 B.n302 B.n301 585
R1274 B.n303 B.n206 585
R1275 B.n305 B.n304 585
R1276 B.n306 B.n205 585
R1277 B.n308 B.n307 585
R1278 B.n309 B.n204 585
R1279 B.n311 B.n310 585
R1280 B.n312 B.n203 585
R1281 B.n314 B.n313 585
R1282 B.n315 B.n202 585
R1283 B.n317 B.n316 585
R1284 B.n318 B.n201 585
R1285 B.n320 B.n319 585
R1286 B.n321 B.n200 585
R1287 B.n323 B.n322 585
R1288 B.n324 B.n199 585
R1289 B.n326 B.n325 585
R1290 B.n327 B.n198 585
R1291 B.n329 B.n328 585
R1292 B.n330 B.n197 585
R1293 B.n332 B.n331 585
R1294 B.n333 B.n196 585
R1295 B.n335 B.n334 585
R1296 B.n336 B.n195 585
R1297 B.n338 B.n337 585
R1298 B.n339 B.n194 585
R1299 B.n341 B.n340 585
R1300 B.n342 B.n193 585
R1301 B.n344 B.n343 585
R1302 B.n343 B.n192 468.476
R1303 B.n445 B.n156 468.476
R1304 B.n679 B.n78 468.476
R1305 B.n777 B.n776 468.476
R1306 B.n171 B.t4 366.769
R1307 B.n63 B.t8 366.769
R1308 B.n177 B.t1 366.769
R1309 B.n56 B.t11 366.769
R1310 B.n172 B.t5 290.743
R1311 B.n64 B.t7 290.743
R1312 B.n178 B.t2 290.743
R1313 B.n57 B.t10 290.743
R1314 B.n177 B.t0 258.045
R1315 B.n171 B.t3 258.045
R1316 B.n63 B.t6 258.045
R1317 B.n56 B.t9 258.045
R1318 B.n893 B.n892 256.663
R1319 B.n892 B.n891 235.042
R1320 B.n892 B.n2 235.042
R1321 B.n347 B.n192 163.367
R1322 B.n348 B.n347 163.367
R1323 B.n349 B.n348 163.367
R1324 B.n349 B.n190 163.367
R1325 B.n353 B.n190 163.367
R1326 B.n354 B.n353 163.367
R1327 B.n355 B.n354 163.367
R1328 B.n355 B.n188 163.367
R1329 B.n359 B.n188 163.367
R1330 B.n360 B.n359 163.367
R1331 B.n361 B.n360 163.367
R1332 B.n361 B.n186 163.367
R1333 B.n365 B.n186 163.367
R1334 B.n366 B.n365 163.367
R1335 B.n367 B.n366 163.367
R1336 B.n367 B.n184 163.367
R1337 B.n371 B.n184 163.367
R1338 B.n372 B.n371 163.367
R1339 B.n373 B.n372 163.367
R1340 B.n373 B.n182 163.367
R1341 B.n377 B.n182 163.367
R1342 B.n378 B.n377 163.367
R1343 B.n379 B.n378 163.367
R1344 B.n379 B.n180 163.367
R1345 B.n383 B.n180 163.367
R1346 B.n384 B.n383 163.367
R1347 B.n385 B.n384 163.367
R1348 B.n385 B.n176 163.367
R1349 B.n390 B.n176 163.367
R1350 B.n391 B.n390 163.367
R1351 B.n392 B.n391 163.367
R1352 B.n392 B.n174 163.367
R1353 B.n396 B.n174 163.367
R1354 B.n397 B.n396 163.367
R1355 B.n398 B.n397 163.367
R1356 B.n398 B.n170 163.367
R1357 B.n403 B.n170 163.367
R1358 B.n404 B.n403 163.367
R1359 B.n405 B.n404 163.367
R1360 B.n405 B.n168 163.367
R1361 B.n409 B.n168 163.367
R1362 B.n410 B.n409 163.367
R1363 B.n411 B.n410 163.367
R1364 B.n411 B.n166 163.367
R1365 B.n415 B.n166 163.367
R1366 B.n416 B.n415 163.367
R1367 B.n417 B.n416 163.367
R1368 B.n417 B.n164 163.367
R1369 B.n421 B.n164 163.367
R1370 B.n422 B.n421 163.367
R1371 B.n423 B.n422 163.367
R1372 B.n423 B.n162 163.367
R1373 B.n427 B.n162 163.367
R1374 B.n428 B.n427 163.367
R1375 B.n429 B.n428 163.367
R1376 B.n429 B.n160 163.367
R1377 B.n433 B.n160 163.367
R1378 B.n434 B.n433 163.367
R1379 B.n435 B.n434 163.367
R1380 B.n435 B.n158 163.367
R1381 B.n439 B.n158 163.367
R1382 B.n440 B.n439 163.367
R1383 B.n441 B.n440 163.367
R1384 B.n441 B.n156 163.367
R1385 B.n675 B.n78 163.367
R1386 B.n675 B.n674 163.367
R1387 B.n674 B.n673 163.367
R1388 B.n673 B.n80 163.367
R1389 B.n669 B.n80 163.367
R1390 B.n669 B.n668 163.367
R1391 B.n668 B.n667 163.367
R1392 B.n667 B.n82 163.367
R1393 B.n663 B.n82 163.367
R1394 B.n663 B.n662 163.367
R1395 B.n662 B.n661 163.367
R1396 B.n661 B.n84 163.367
R1397 B.n657 B.n84 163.367
R1398 B.n657 B.n656 163.367
R1399 B.n656 B.n655 163.367
R1400 B.n655 B.n86 163.367
R1401 B.n651 B.n86 163.367
R1402 B.n651 B.n650 163.367
R1403 B.n650 B.n649 163.367
R1404 B.n649 B.n88 163.367
R1405 B.n645 B.n88 163.367
R1406 B.n645 B.n644 163.367
R1407 B.n644 B.n643 163.367
R1408 B.n643 B.n90 163.367
R1409 B.n639 B.n90 163.367
R1410 B.n639 B.n638 163.367
R1411 B.n638 B.n637 163.367
R1412 B.n637 B.n92 163.367
R1413 B.n633 B.n92 163.367
R1414 B.n633 B.n632 163.367
R1415 B.n632 B.n631 163.367
R1416 B.n631 B.n94 163.367
R1417 B.n627 B.n94 163.367
R1418 B.n627 B.n626 163.367
R1419 B.n626 B.n625 163.367
R1420 B.n625 B.n96 163.367
R1421 B.n621 B.n96 163.367
R1422 B.n621 B.n620 163.367
R1423 B.n620 B.n619 163.367
R1424 B.n619 B.n98 163.367
R1425 B.n615 B.n98 163.367
R1426 B.n615 B.n614 163.367
R1427 B.n614 B.n613 163.367
R1428 B.n613 B.n100 163.367
R1429 B.n609 B.n100 163.367
R1430 B.n609 B.n608 163.367
R1431 B.n608 B.n607 163.367
R1432 B.n607 B.n102 163.367
R1433 B.n603 B.n102 163.367
R1434 B.n603 B.n602 163.367
R1435 B.n602 B.n601 163.367
R1436 B.n601 B.n104 163.367
R1437 B.n597 B.n104 163.367
R1438 B.n597 B.n596 163.367
R1439 B.n596 B.n595 163.367
R1440 B.n595 B.n106 163.367
R1441 B.n591 B.n106 163.367
R1442 B.n591 B.n590 163.367
R1443 B.n590 B.n589 163.367
R1444 B.n589 B.n108 163.367
R1445 B.n585 B.n108 163.367
R1446 B.n585 B.n584 163.367
R1447 B.n584 B.n583 163.367
R1448 B.n583 B.n110 163.367
R1449 B.n579 B.n110 163.367
R1450 B.n579 B.n578 163.367
R1451 B.n578 B.n577 163.367
R1452 B.n577 B.n112 163.367
R1453 B.n573 B.n112 163.367
R1454 B.n573 B.n572 163.367
R1455 B.n572 B.n571 163.367
R1456 B.n571 B.n114 163.367
R1457 B.n567 B.n114 163.367
R1458 B.n567 B.n566 163.367
R1459 B.n566 B.n565 163.367
R1460 B.n565 B.n116 163.367
R1461 B.n561 B.n116 163.367
R1462 B.n561 B.n560 163.367
R1463 B.n560 B.n559 163.367
R1464 B.n559 B.n118 163.367
R1465 B.n555 B.n118 163.367
R1466 B.n555 B.n554 163.367
R1467 B.n554 B.n553 163.367
R1468 B.n553 B.n120 163.367
R1469 B.n549 B.n120 163.367
R1470 B.n549 B.n548 163.367
R1471 B.n548 B.n547 163.367
R1472 B.n547 B.n122 163.367
R1473 B.n543 B.n122 163.367
R1474 B.n543 B.n542 163.367
R1475 B.n542 B.n541 163.367
R1476 B.n541 B.n124 163.367
R1477 B.n537 B.n124 163.367
R1478 B.n537 B.n536 163.367
R1479 B.n536 B.n535 163.367
R1480 B.n535 B.n126 163.367
R1481 B.n531 B.n126 163.367
R1482 B.n531 B.n530 163.367
R1483 B.n530 B.n529 163.367
R1484 B.n529 B.n128 163.367
R1485 B.n525 B.n128 163.367
R1486 B.n525 B.n524 163.367
R1487 B.n524 B.n523 163.367
R1488 B.n523 B.n130 163.367
R1489 B.n519 B.n130 163.367
R1490 B.n519 B.n518 163.367
R1491 B.n518 B.n517 163.367
R1492 B.n517 B.n132 163.367
R1493 B.n513 B.n132 163.367
R1494 B.n513 B.n512 163.367
R1495 B.n512 B.n511 163.367
R1496 B.n511 B.n134 163.367
R1497 B.n507 B.n134 163.367
R1498 B.n507 B.n506 163.367
R1499 B.n506 B.n505 163.367
R1500 B.n505 B.n136 163.367
R1501 B.n501 B.n136 163.367
R1502 B.n501 B.n500 163.367
R1503 B.n500 B.n499 163.367
R1504 B.n499 B.n138 163.367
R1505 B.n495 B.n138 163.367
R1506 B.n495 B.n494 163.367
R1507 B.n494 B.n493 163.367
R1508 B.n493 B.n140 163.367
R1509 B.n489 B.n140 163.367
R1510 B.n489 B.n488 163.367
R1511 B.n488 B.n487 163.367
R1512 B.n487 B.n142 163.367
R1513 B.n483 B.n142 163.367
R1514 B.n483 B.n482 163.367
R1515 B.n482 B.n481 163.367
R1516 B.n481 B.n144 163.367
R1517 B.n477 B.n144 163.367
R1518 B.n477 B.n476 163.367
R1519 B.n476 B.n475 163.367
R1520 B.n475 B.n146 163.367
R1521 B.n471 B.n146 163.367
R1522 B.n471 B.n470 163.367
R1523 B.n470 B.n469 163.367
R1524 B.n469 B.n148 163.367
R1525 B.n465 B.n148 163.367
R1526 B.n465 B.n464 163.367
R1527 B.n464 B.n463 163.367
R1528 B.n463 B.n150 163.367
R1529 B.n459 B.n150 163.367
R1530 B.n459 B.n458 163.367
R1531 B.n458 B.n457 163.367
R1532 B.n457 B.n152 163.367
R1533 B.n453 B.n152 163.367
R1534 B.n453 B.n452 163.367
R1535 B.n452 B.n451 163.367
R1536 B.n451 B.n154 163.367
R1537 B.n447 B.n154 163.367
R1538 B.n447 B.n446 163.367
R1539 B.n446 B.n445 163.367
R1540 B.n776 B.n41 163.367
R1541 B.n772 B.n41 163.367
R1542 B.n772 B.n771 163.367
R1543 B.n771 B.n770 163.367
R1544 B.n770 B.n43 163.367
R1545 B.n766 B.n43 163.367
R1546 B.n766 B.n765 163.367
R1547 B.n765 B.n764 163.367
R1548 B.n764 B.n45 163.367
R1549 B.n760 B.n45 163.367
R1550 B.n760 B.n759 163.367
R1551 B.n759 B.n758 163.367
R1552 B.n758 B.n47 163.367
R1553 B.n754 B.n47 163.367
R1554 B.n754 B.n753 163.367
R1555 B.n753 B.n752 163.367
R1556 B.n752 B.n49 163.367
R1557 B.n748 B.n49 163.367
R1558 B.n748 B.n747 163.367
R1559 B.n747 B.n746 163.367
R1560 B.n746 B.n51 163.367
R1561 B.n742 B.n51 163.367
R1562 B.n742 B.n741 163.367
R1563 B.n741 B.n740 163.367
R1564 B.n740 B.n53 163.367
R1565 B.n736 B.n53 163.367
R1566 B.n736 B.n735 163.367
R1567 B.n735 B.n734 163.367
R1568 B.n734 B.n55 163.367
R1569 B.n730 B.n55 163.367
R1570 B.n730 B.n729 163.367
R1571 B.n729 B.n728 163.367
R1572 B.n728 B.n60 163.367
R1573 B.n724 B.n60 163.367
R1574 B.n724 B.n723 163.367
R1575 B.n723 B.n722 163.367
R1576 B.n722 B.n62 163.367
R1577 B.n717 B.n62 163.367
R1578 B.n717 B.n716 163.367
R1579 B.n716 B.n715 163.367
R1580 B.n715 B.n66 163.367
R1581 B.n711 B.n66 163.367
R1582 B.n711 B.n710 163.367
R1583 B.n710 B.n709 163.367
R1584 B.n709 B.n68 163.367
R1585 B.n705 B.n68 163.367
R1586 B.n705 B.n704 163.367
R1587 B.n704 B.n703 163.367
R1588 B.n703 B.n70 163.367
R1589 B.n699 B.n70 163.367
R1590 B.n699 B.n698 163.367
R1591 B.n698 B.n697 163.367
R1592 B.n697 B.n72 163.367
R1593 B.n693 B.n72 163.367
R1594 B.n693 B.n692 163.367
R1595 B.n692 B.n691 163.367
R1596 B.n691 B.n74 163.367
R1597 B.n687 B.n74 163.367
R1598 B.n687 B.n686 163.367
R1599 B.n686 B.n685 163.367
R1600 B.n685 B.n76 163.367
R1601 B.n681 B.n76 163.367
R1602 B.n681 B.n680 163.367
R1603 B.n680 B.n679 163.367
R1604 B.n778 B.n777 163.367
R1605 B.n778 B.n39 163.367
R1606 B.n782 B.n39 163.367
R1607 B.n783 B.n782 163.367
R1608 B.n784 B.n783 163.367
R1609 B.n784 B.n37 163.367
R1610 B.n788 B.n37 163.367
R1611 B.n789 B.n788 163.367
R1612 B.n790 B.n789 163.367
R1613 B.n790 B.n35 163.367
R1614 B.n794 B.n35 163.367
R1615 B.n795 B.n794 163.367
R1616 B.n796 B.n795 163.367
R1617 B.n796 B.n33 163.367
R1618 B.n800 B.n33 163.367
R1619 B.n801 B.n800 163.367
R1620 B.n802 B.n801 163.367
R1621 B.n802 B.n31 163.367
R1622 B.n806 B.n31 163.367
R1623 B.n807 B.n806 163.367
R1624 B.n808 B.n807 163.367
R1625 B.n808 B.n29 163.367
R1626 B.n812 B.n29 163.367
R1627 B.n813 B.n812 163.367
R1628 B.n814 B.n813 163.367
R1629 B.n814 B.n27 163.367
R1630 B.n818 B.n27 163.367
R1631 B.n819 B.n818 163.367
R1632 B.n820 B.n819 163.367
R1633 B.n820 B.n25 163.367
R1634 B.n824 B.n25 163.367
R1635 B.n825 B.n824 163.367
R1636 B.n826 B.n825 163.367
R1637 B.n826 B.n23 163.367
R1638 B.n830 B.n23 163.367
R1639 B.n831 B.n830 163.367
R1640 B.n832 B.n831 163.367
R1641 B.n832 B.n21 163.367
R1642 B.n836 B.n21 163.367
R1643 B.n837 B.n836 163.367
R1644 B.n838 B.n837 163.367
R1645 B.n838 B.n19 163.367
R1646 B.n842 B.n19 163.367
R1647 B.n843 B.n842 163.367
R1648 B.n844 B.n843 163.367
R1649 B.n844 B.n17 163.367
R1650 B.n848 B.n17 163.367
R1651 B.n849 B.n848 163.367
R1652 B.n850 B.n849 163.367
R1653 B.n850 B.n15 163.367
R1654 B.n854 B.n15 163.367
R1655 B.n855 B.n854 163.367
R1656 B.n856 B.n855 163.367
R1657 B.n856 B.n13 163.367
R1658 B.n860 B.n13 163.367
R1659 B.n861 B.n860 163.367
R1660 B.n862 B.n861 163.367
R1661 B.n862 B.n11 163.367
R1662 B.n866 B.n11 163.367
R1663 B.n867 B.n866 163.367
R1664 B.n868 B.n867 163.367
R1665 B.n868 B.n9 163.367
R1666 B.n872 B.n9 163.367
R1667 B.n873 B.n872 163.367
R1668 B.n874 B.n873 163.367
R1669 B.n874 B.n7 163.367
R1670 B.n878 B.n7 163.367
R1671 B.n879 B.n878 163.367
R1672 B.n880 B.n879 163.367
R1673 B.n880 B.n5 163.367
R1674 B.n884 B.n5 163.367
R1675 B.n885 B.n884 163.367
R1676 B.n886 B.n885 163.367
R1677 B.n886 B.n3 163.367
R1678 B.n890 B.n3 163.367
R1679 B.n891 B.n890 163.367
R1680 B.n230 B.n2 163.367
R1681 B.n233 B.n230 163.367
R1682 B.n234 B.n233 163.367
R1683 B.n235 B.n234 163.367
R1684 B.n235 B.n228 163.367
R1685 B.n239 B.n228 163.367
R1686 B.n240 B.n239 163.367
R1687 B.n241 B.n240 163.367
R1688 B.n241 B.n226 163.367
R1689 B.n245 B.n226 163.367
R1690 B.n246 B.n245 163.367
R1691 B.n247 B.n246 163.367
R1692 B.n247 B.n224 163.367
R1693 B.n251 B.n224 163.367
R1694 B.n252 B.n251 163.367
R1695 B.n253 B.n252 163.367
R1696 B.n253 B.n222 163.367
R1697 B.n257 B.n222 163.367
R1698 B.n258 B.n257 163.367
R1699 B.n259 B.n258 163.367
R1700 B.n259 B.n220 163.367
R1701 B.n263 B.n220 163.367
R1702 B.n264 B.n263 163.367
R1703 B.n265 B.n264 163.367
R1704 B.n265 B.n218 163.367
R1705 B.n269 B.n218 163.367
R1706 B.n270 B.n269 163.367
R1707 B.n271 B.n270 163.367
R1708 B.n271 B.n216 163.367
R1709 B.n275 B.n216 163.367
R1710 B.n276 B.n275 163.367
R1711 B.n277 B.n276 163.367
R1712 B.n277 B.n214 163.367
R1713 B.n281 B.n214 163.367
R1714 B.n282 B.n281 163.367
R1715 B.n283 B.n282 163.367
R1716 B.n283 B.n212 163.367
R1717 B.n287 B.n212 163.367
R1718 B.n288 B.n287 163.367
R1719 B.n289 B.n288 163.367
R1720 B.n289 B.n210 163.367
R1721 B.n293 B.n210 163.367
R1722 B.n294 B.n293 163.367
R1723 B.n295 B.n294 163.367
R1724 B.n295 B.n208 163.367
R1725 B.n299 B.n208 163.367
R1726 B.n300 B.n299 163.367
R1727 B.n301 B.n300 163.367
R1728 B.n301 B.n206 163.367
R1729 B.n305 B.n206 163.367
R1730 B.n306 B.n305 163.367
R1731 B.n307 B.n306 163.367
R1732 B.n307 B.n204 163.367
R1733 B.n311 B.n204 163.367
R1734 B.n312 B.n311 163.367
R1735 B.n313 B.n312 163.367
R1736 B.n313 B.n202 163.367
R1737 B.n317 B.n202 163.367
R1738 B.n318 B.n317 163.367
R1739 B.n319 B.n318 163.367
R1740 B.n319 B.n200 163.367
R1741 B.n323 B.n200 163.367
R1742 B.n324 B.n323 163.367
R1743 B.n325 B.n324 163.367
R1744 B.n325 B.n198 163.367
R1745 B.n329 B.n198 163.367
R1746 B.n330 B.n329 163.367
R1747 B.n331 B.n330 163.367
R1748 B.n331 B.n196 163.367
R1749 B.n335 B.n196 163.367
R1750 B.n336 B.n335 163.367
R1751 B.n337 B.n336 163.367
R1752 B.n337 B.n194 163.367
R1753 B.n341 B.n194 163.367
R1754 B.n342 B.n341 163.367
R1755 B.n343 B.n342 163.367
R1756 B.n178 B.n177 76.0247
R1757 B.n172 B.n171 76.0247
R1758 B.n64 B.n63 76.0247
R1759 B.n57 B.n56 76.0247
R1760 B.n387 B.n178 59.5399
R1761 B.n401 B.n172 59.5399
R1762 B.n720 B.n64 59.5399
R1763 B.n58 B.n57 59.5399
R1764 B.n775 B.n40 30.4395
R1765 B.n678 B.n677 30.4395
R1766 B.n345 B.n344 30.4395
R1767 B.n444 B.n443 30.4395
R1768 B B.n893 18.0485
R1769 B.n779 B.n40 10.6151
R1770 B.n780 B.n779 10.6151
R1771 B.n781 B.n780 10.6151
R1772 B.n781 B.n38 10.6151
R1773 B.n785 B.n38 10.6151
R1774 B.n786 B.n785 10.6151
R1775 B.n787 B.n786 10.6151
R1776 B.n787 B.n36 10.6151
R1777 B.n791 B.n36 10.6151
R1778 B.n792 B.n791 10.6151
R1779 B.n793 B.n792 10.6151
R1780 B.n793 B.n34 10.6151
R1781 B.n797 B.n34 10.6151
R1782 B.n798 B.n797 10.6151
R1783 B.n799 B.n798 10.6151
R1784 B.n799 B.n32 10.6151
R1785 B.n803 B.n32 10.6151
R1786 B.n804 B.n803 10.6151
R1787 B.n805 B.n804 10.6151
R1788 B.n805 B.n30 10.6151
R1789 B.n809 B.n30 10.6151
R1790 B.n810 B.n809 10.6151
R1791 B.n811 B.n810 10.6151
R1792 B.n811 B.n28 10.6151
R1793 B.n815 B.n28 10.6151
R1794 B.n816 B.n815 10.6151
R1795 B.n817 B.n816 10.6151
R1796 B.n817 B.n26 10.6151
R1797 B.n821 B.n26 10.6151
R1798 B.n822 B.n821 10.6151
R1799 B.n823 B.n822 10.6151
R1800 B.n823 B.n24 10.6151
R1801 B.n827 B.n24 10.6151
R1802 B.n828 B.n827 10.6151
R1803 B.n829 B.n828 10.6151
R1804 B.n829 B.n22 10.6151
R1805 B.n833 B.n22 10.6151
R1806 B.n834 B.n833 10.6151
R1807 B.n835 B.n834 10.6151
R1808 B.n835 B.n20 10.6151
R1809 B.n839 B.n20 10.6151
R1810 B.n840 B.n839 10.6151
R1811 B.n841 B.n840 10.6151
R1812 B.n841 B.n18 10.6151
R1813 B.n845 B.n18 10.6151
R1814 B.n846 B.n845 10.6151
R1815 B.n847 B.n846 10.6151
R1816 B.n847 B.n16 10.6151
R1817 B.n851 B.n16 10.6151
R1818 B.n852 B.n851 10.6151
R1819 B.n853 B.n852 10.6151
R1820 B.n853 B.n14 10.6151
R1821 B.n857 B.n14 10.6151
R1822 B.n858 B.n857 10.6151
R1823 B.n859 B.n858 10.6151
R1824 B.n859 B.n12 10.6151
R1825 B.n863 B.n12 10.6151
R1826 B.n864 B.n863 10.6151
R1827 B.n865 B.n864 10.6151
R1828 B.n865 B.n10 10.6151
R1829 B.n869 B.n10 10.6151
R1830 B.n870 B.n869 10.6151
R1831 B.n871 B.n870 10.6151
R1832 B.n871 B.n8 10.6151
R1833 B.n875 B.n8 10.6151
R1834 B.n876 B.n875 10.6151
R1835 B.n877 B.n876 10.6151
R1836 B.n877 B.n6 10.6151
R1837 B.n881 B.n6 10.6151
R1838 B.n882 B.n881 10.6151
R1839 B.n883 B.n882 10.6151
R1840 B.n883 B.n4 10.6151
R1841 B.n887 B.n4 10.6151
R1842 B.n888 B.n887 10.6151
R1843 B.n889 B.n888 10.6151
R1844 B.n889 B.n0 10.6151
R1845 B.n775 B.n774 10.6151
R1846 B.n774 B.n773 10.6151
R1847 B.n773 B.n42 10.6151
R1848 B.n769 B.n42 10.6151
R1849 B.n769 B.n768 10.6151
R1850 B.n768 B.n767 10.6151
R1851 B.n767 B.n44 10.6151
R1852 B.n763 B.n44 10.6151
R1853 B.n763 B.n762 10.6151
R1854 B.n762 B.n761 10.6151
R1855 B.n761 B.n46 10.6151
R1856 B.n757 B.n46 10.6151
R1857 B.n757 B.n756 10.6151
R1858 B.n756 B.n755 10.6151
R1859 B.n755 B.n48 10.6151
R1860 B.n751 B.n48 10.6151
R1861 B.n751 B.n750 10.6151
R1862 B.n750 B.n749 10.6151
R1863 B.n749 B.n50 10.6151
R1864 B.n745 B.n50 10.6151
R1865 B.n745 B.n744 10.6151
R1866 B.n744 B.n743 10.6151
R1867 B.n743 B.n52 10.6151
R1868 B.n739 B.n52 10.6151
R1869 B.n739 B.n738 10.6151
R1870 B.n738 B.n737 10.6151
R1871 B.n737 B.n54 10.6151
R1872 B.n733 B.n732 10.6151
R1873 B.n732 B.n731 10.6151
R1874 B.n731 B.n59 10.6151
R1875 B.n727 B.n59 10.6151
R1876 B.n727 B.n726 10.6151
R1877 B.n726 B.n725 10.6151
R1878 B.n725 B.n61 10.6151
R1879 B.n721 B.n61 10.6151
R1880 B.n719 B.n718 10.6151
R1881 B.n718 B.n65 10.6151
R1882 B.n714 B.n65 10.6151
R1883 B.n714 B.n713 10.6151
R1884 B.n713 B.n712 10.6151
R1885 B.n712 B.n67 10.6151
R1886 B.n708 B.n67 10.6151
R1887 B.n708 B.n707 10.6151
R1888 B.n707 B.n706 10.6151
R1889 B.n706 B.n69 10.6151
R1890 B.n702 B.n69 10.6151
R1891 B.n702 B.n701 10.6151
R1892 B.n701 B.n700 10.6151
R1893 B.n700 B.n71 10.6151
R1894 B.n696 B.n71 10.6151
R1895 B.n696 B.n695 10.6151
R1896 B.n695 B.n694 10.6151
R1897 B.n694 B.n73 10.6151
R1898 B.n690 B.n73 10.6151
R1899 B.n690 B.n689 10.6151
R1900 B.n689 B.n688 10.6151
R1901 B.n688 B.n75 10.6151
R1902 B.n684 B.n75 10.6151
R1903 B.n684 B.n683 10.6151
R1904 B.n683 B.n682 10.6151
R1905 B.n682 B.n77 10.6151
R1906 B.n678 B.n77 10.6151
R1907 B.n677 B.n676 10.6151
R1908 B.n676 B.n79 10.6151
R1909 B.n672 B.n79 10.6151
R1910 B.n672 B.n671 10.6151
R1911 B.n671 B.n670 10.6151
R1912 B.n670 B.n81 10.6151
R1913 B.n666 B.n81 10.6151
R1914 B.n666 B.n665 10.6151
R1915 B.n665 B.n664 10.6151
R1916 B.n664 B.n83 10.6151
R1917 B.n660 B.n83 10.6151
R1918 B.n660 B.n659 10.6151
R1919 B.n659 B.n658 10.6151
R1920 B.n658 B.n85 10.6151
R1921 B.n654 B.n85 10.6151
R1922 B.n654 B.n653 10.6151
R1923 B.n653 B.n652 10.6151
R1924 B.n652 B.n87 10.6151
R1925 B.n648 B.n87 10.6151
R1926 B.n648 B.n647 10.6151
R1927 B.n647 B.n646 10.6151
R1928 B.n646 B.n89 10.6151
R1929 B.n642 B.n89 10.6151
R1930 B.n642 B.n641 10.6151
R1931 B.n641 B.n640 10.6151
R1932 B.n640 B.n91 10.6151
R1933 B.n636 B.n91 10.6151
R1934 B.n636 B.n635 10.6151
R1935 B.n635 B.n634 10.6151
R1936 B.n634 B.n93 10.6151
R1937 B.n630 B.n93 10.6151
R1938 B.n630 B.n629 10.6151
R1939 B.n629 B.n628 10.6151
R1940 B.n628 B.n95 10.6151
R1941 B.n624 B.n95 10.6151
R1942 B.n624 B.n623 10.6151
R1943 B.n623 B.n622 10.6151
R1944 B.n622 B.n97 10.6151
R1945 B.n618 B.n97 10.6151
R1946 B.n618 B.n617 10.6151
R1947 B.n617 B.n616 10.6151
R1948 B.n616 B.n99 10.6151
R1949 B.n612 B.n99 10.6151
R1950 B.n612 B.n611 10.6151
R1951 B.n611 B.n610 10.6151
R1952 B.n610 B.n101 10.6151
R1953 B.n606 B.n101 10.6151
R1954 B.n606 B.n605 10.6151
R1955 B.n605 B.n604 10.6151
R1956 B.n604 B.n103 10.6151
R1957 B.n600 B.n103 10.6151
R1958 B.n600 B.n599 10.6151
R1959 B.n599 B.n598 10.6151
R1960 B.n598 B.n105 10.6151
R1961 B.n594 B.n105 10.6151
R1962 B.n594 B.n593 10.6151
R1963 B.n593 B.n592 10.6151
R1964 B.n592 B.n107 10.6151
R1965 B.n588 B.n107 10.6151
R1966 B.n588 B.n587 10.6151
R1967 B.n587 B.n586 10.6151
R1968 B.n586 B.n109 10.6151
R1969 B.n582 B.n109 10.6151
R1970 B.n582 B.n581 10.6151
R1971 B.n581 B.n580 10.6151
R1972 B.n580 B.n111 10.6151
R1973 B.n576 B.n111 10.6151
R1974 B.n576 B.n575 10.6151
R1975 B.n575 B.n574 10.6151
R1976 B.n574 B.n113 10.6151
R1977 B.n570 B.n113 10.6151
R1978 B.n570 B.n569 10.6151
R1979 B.n569 B.n568 10.6151
R1980 B.n568 B.n115 10.6151
R1981 B.n564 B.n115 10.6151
R1982 B.n564 B.n563 10.6151
R1983 B.n563 B.n562 10.6151
R1984 B.n562 B.n117 10.6151
R1985 B.n558 B.n117 10.6151
R1986 B.n558 B.n557 10.6151
R1987 B.n557 B.n556 10.6151
R1988 B.n556 B.n119 10.6151
R1989 B.n552 B.n119 10.6151
R1990 B.n552 B.n551 10.6151
R1991 B.n551 B.n550 10.6151
R1992 B.n550 B.n121 10.6151
R1993 B.n546 B.n121 10.6151
R1994 B.n546 B.n545 10.6151
R1995 B.n545 B.n544 10.6151
R1996 B.n544 B.n123 10.6151
R1997 B.n540 B.n123 10.6151
R1998 B.n540 B.n539 10.6151
R1999 B.n539 B.n538 10.6151
R2000 B.n538 B.n125 10.6151
R2001 B.n534 B.n125 10.6151
R2002 B.n534 B.n533 10.6151
R2003 B.n533 B.n532 10.6151
R2004 B.n532 B.n127 10.6151
R2005 B.n528 B.n127 10.6151
R2006 B.n528 B.n527 10.6151
R2007 B.n527 B.n526 10.6151
R2008 B.n526 B.n129 10.6151
R2009 B.n522 B.n129 10.6151
R2010 B.n522 B.n521 10.6151
R2011 B.n521 B.n520 10.6151
R2012 B.n520 B.n131 10.6151
R2013 B.n516 B.n131 10.6151
R2014 B.n516 B.n515 10.6151
R2015 B.n515 B.n514 10.6151
R2016 B.n514 B.n133 10.6151
R2017 B.n510 B.n133 10.6151
R2018 B.n510 B.n509 10.6151
R2019 B.n509 B.n508 10.6151
R2020 B.n508 B.n135 10.6151
R2021 B.n504 B.n135 10.6151
R2022 B.n504 B.n503 10.6151
R2023 B.n503 B.n502 10.6151
R2024 B.n502 B.n137 10.6151
R2025 B.n498 B.n137 10.6151
R2026 B.n498 B.n497 10.6151
R2027 B.n497 B.n496 10.6151
R2028 B.n496 B.n139 10.6151
R2029 B.n492 B.n139 10.6151
R2030 B.n492 B.n491 10.6151
R2031 B.n491 B.n490 10.6151
R2032 B.n490 B.n141 10.6151
R2033 B.n486 B.n141 10.6151
R2034 B.n486 B.n485 10.6151
R2035 B.n485 B.n484 10.6151
R2036 B.n484 B.n143 10.6151
R2037 B.n480 B.n143 10.6151
R2038 B.n480 B.n479 10.6151
R2039 B.n479 B.n478 10.6151
R2040 B.n478 B.n145 10.6151
R2041 B.n474 B.n145 10.6151
R2042 B.n474 B.n473 10.6151
R2043 B.n473 B.n472 10.6151
R2044 B.n472 B.n147 10.6151
R2045 B.n468 B.n147 10.6151
R2046 B.n468 B.n467 10.6151
R2047 B.n467 B.n466 10.6151
R2048 B.n466 B.n149 10.6151
R2049 B.n462 B.n149 10.6151
R2050 B.n462 B.n461 10.6151
R2051 B.n461 B.n460 10.6151
R2052 B.n460 B.n151 10.6151
R2053 B.n456 B.n151 10.6151
R2054 B.n456 B.n455 10.6151
R2055 B.n455 B.n454 10.6151
R2056 B.n454 B.n153 10.6151
R2057 B.n450 B.n153 10.6151
R2058 B.n450 B.n449 10.6151
R2059 B.n449 B.n448 10.6151
R2060 B.n448 B.n155 10.6151
R2061 B.n444 B.n155 10.6151
R2062 B.n231 B.n1 10.6151
R2063 B.n232 B.n231 10.6151
R2064 B.n232 B.n229 10.6151
R2065 B.n236 B.n229 10.6151
R2066 B.n237 B.n236 10.6151
R2067 B.n238 B.n237 10.6151
R2068 B.n238 B.n227 10.6151
R2069 B.n242 B.n227 10.6151
R2070 B.n243 B.n242 10.6151
R2071 B.n244 B.n243 10.6151
R2072 B.n244 B.n225 10.6151
R2073 B.n248 B.n225 10.6151
R2074 B.n249 B.n248 10.6151
R2075 B.n250 B.n249 10.6151
R2076 B.n250 B.n223 10.6151
R2077 B.n254 B.n223 10.6151
R2078 B.n255 B.n254 10.6151
R2079 B.n256 B.n255 10.6151
R2080 B.n256 B.n221 10.6151
R2081 B.n260 B.n221 10.6151
R2082 B.n261 B.n260 10.6151
R2083 B.n262 B.n261 10.6151
R2084 B.n262 B.n219 10.6151
R2085 B.n266 B.n219 10.6151
R2086 B.n267 B.n266 10.6151
R2087 B.n268 B.n267 10.6151
R2088 B.n268 B.n217 10.6151
R2089 B.n272 B.n217 10.6151
R2090 B.n273 B.n272 10.6151
R2091 B.n274 B.n273 10.6151
R2092 B.n274 B.n215 10.6151
R2093 B.n278 B.n215 10.6151
R2094 B.n279 B.n278 10.6151
R2095 B.n280 B.n279 10.6151
R2096 B.n280 B.n213 10.6151
R2097 B.n284 B.n213 10.6151
R2098 B.n285 B.n284 10.6151
R2099 B.n286 B.n285 10.6151
R2100 B.n286 B.n211 10.6151
R2101 B.n290 B.n211 10.6151
R2102 B.n291 B.n290 10.6151
R2103 B.n292 B.n291 10.6151
R2104 B.n292 B.n209 10.6151
R2105 B.n296 B.n209 10.6151
R2106 B.n297 B.n296 10.6151
R2107 B.n298 B.n297 10.6151
R2108 B.n298 B.n207 10.6151
R2109 B.n302 B.n207 10.6151
R2110 B.n303 B.n302 10.6151
R2111 B.n304 B.n303 10.6151
R2112 B.n304 B.n205 10.6151
R2113 B.n308 B.n205 10.6151
R2114 B.n309 B.n308 10.6151
R2115 B.n310 B.n309 10.6151
R2116 B.n310 B.n203 10.6151
R2117 B.n314 B.n203 10.6151
R2118 B.n315 B.n314 10.6151
R2119 B.n316 B.n315 10.6151
R2120 B.n316 B.n201 10.6151
R2121 B.n320 B.n201 10.6151
R2122 B.n321 B.n320 10.6151
R2123 B.n322 B.n321 10.6151
R2124 B.n322 B.n199 10.6151
R2125 B.n326 B.n199 10.6151
R2126 B.n327 B.n326 10.6151
R2127 B.n328 B.n327 10.6151
R2128 B.n328 B.n197 10.6151
R2129 B.n332 B.n197 10.6151
R2130 B.n333 B.n332 10.6151
R2131 B.n334 B.n333 10.6151
R2132 B.n334 B.n195 10.6151
R2133 B.n338 B.n195 10.6151
R2134 B.n339 B.n338 10.6151
R2135 B.n340 B.n339 10.6151
R2136 B.n340 B.n193 10.6151
R2137 B.n344 B.n193 10.6151
R2138 B.n346 B.n345 10.6151
R2139 B.n346 B.n191 10.6151
R2140 B.n350 B.n191 10.6151
R2141 B.n351 B.n350 10.6151
R2142 B.n352 B.n351 10.6151
R2143 B.n352 B.n189 10.6151
R2144 B.n356 B.n189 10.6151
R2145 B.n357 B.n356 10.6151
R2146 B.n358 B.n357 10.6151
R2147 B.n358 B.n187 10.6151
R2148 B.n362 B.n187 10.6151
R2149 B.n363 B.n362 10.6151
R2150 B.n364 B.n363 10.6151
R2151 B.n364 B.n185 10.6151
R2152 B.n368 B.n185 10.6151
R2153 B.n369 B.n368 10.6151
R2154 B.n370 B.n369 10.6151
R2155 B.n370 B.n183 10.6151
R2156 B.n374 B.n183 10.6151
R2157 B.n375 B.n374 10.6151
R2158 B.n376 B.n375 10.6151
R2159 B.n376 B.n181 10.6151
R2160 B.n380 B.n181 10.6151
R2161 B.n381 B.n380 10.6151
R2162 B.n382 B.n381 10.6151
R2163 B.n382 B.n179 10.6151
R2164 B.n386 B.n179 10.6151
R2165 B.n389 B.n388 10.6151
R2166 B.n389 B.n175 10.6151
R2167 B.n393 B.n175 10.6151
R2168 B.n394 B.n393 10.6151
R2169 B.n395 B.n394 10.6151
R2170 B.n395 B.n173 10.6151
R2171 B.n399 B.n173 10.6151
R2172 B.n400 B.n399 10.6151
R2173 B.n402 B.n169 10.6151
R2174 B.n406 B.n169 10.6151
R2175 B.n407 B.n406 10.6151
R2176 B.n408 B.n407 10.6151
R2177 B.n408 B.n167 10.6151
R2178 B.n412 B.n167 10.6151
R2179 B.n413 B.n412 10.6151
R2180 B.n414 B.n413 10.6151
R2181 B.n414 B.n165 10.6151
R2182 B.n418 B.n165 10.6151
R2183 B.n419 B.n418 10.6151
R2184 B.n420 B.n419 10.6151
R2185 B.n420 B.n163 10.6151
R2186 B.n424 B.n163 10.6151
R2187 B.n425 B.n424 10.6151
R2188 B.n426 B.n425 10.6151
R2189 B.n426 B.n161 10.6151
R2190 B.n430 B.n161 10.6151
R2191 B.n431 B.n430 10.6151
R2192 B.n432 B.n431 10.6151
R2193 B.n432 B.n159 10.6151
R2194 B.n436 B.n159 10.6151
R2195 B.n437 B.n436 10.6151
R2196 B.n438 B.n437 10.6151
R2197 B.n438 B.n157 10.6151
R2198 B.n442 B.n157 10.6151
R2199 B.n443 B.n442 10.6151
R2200 B.n893 B.n0 8.11757
R2201 B.n893 B.n1 8.11757
R2202 B.n733 B.n58 6.5566
R2203 B.n721 B.n720 6.5566
R2204 B.n388 B.n387 6.5566
R2205 B.n401 B.n400 6.5566
R2206 B.n58 B.n54 4.05904
R2207 B.n720 B.n719 4.05904
R2208 B.n387 B.n386 4.05904
R2209 B.n402 B.n401 4.05904
C0 w_n5674_n2424# VP 13.0781f
C1 VDD2 VTAIL 9.048611f
C2 VDD2 B 2.64152f
C3 VTAIL VDD1 8.989409f
C4 B VDD1 2.48505f
C5 VDD2 VDD1 2.8197f
C6 VN VTAIL 8.348559f
C7 B VN 1.48436f
C8 w_n5674_n2424# VTAIL 2.71821f
C9 VDD2 VN 7.05344f
C10 w_n5674_n2424# B 10.8896f
C11 VN VDD1 0.156062f
C12 VP VTAIL 8.36278f
C13 B VP 2.73717f
C14 VDD2 w_n5674_n2424# 3.03805f
C15 w_n5674_n2424# VDD1 2.84304f
C16 VDD2 VP 0.710014f
C17 VP VDD1 7.6041f
C18 w_n5674_n2424# VN 12.3363f
C19 VP VN 8.978621f
C20 B VTAIL 2.99078f
C21 VDD2 VSUBS 2.471304f
C22 VDD1 VSUBS 2.268249f
C23 VTAIL VSUBS 1.388423f
C24 VN VSUBS 9.336201f
C25 VP VSUBS 5.328822f
C26 B VSUBS 6.19658f
C27 w_n5674_n2424# VSUBS 0.170969p
C28 B.n0 VSUBS 0.009491f
C29 B.n1 VSUBS 0.009491f
C30 B.n2 VSUBS 0.014037f
C31 B.n3 VSUBS 0.010757f
C32 B.n4 VSUBS 0.010757f
C33 B.n5 VSUBS 0.010757f
C34 B.n6 VSUBS 0.010757f
C35 B.n7 VSUBS 0.010757f
C36 B.n8 VSUBS 0.010757f
C37 B.n9 VSUBS 0.010757f
C38 B.n10 VSUBS 0.010757f
C39 B.n11 VSUBS 0.010757f
C40 B.n12 VSUBS 0.010757f
C41 B.n13 VSUBS 0.010757f
C42 B.n14 VSUBS 0.010757f
C43 B.n15 VSUBS 0.010757f
C44 B.n16 VSUBS 0.010757f
C45 B.n17 VSUBS 0.010757f
C46 B.n18 VSUBS 0.010757f
C47 B.n19 VSUBS 0.010757f
C48 B.n20 VSUBS 0.010757f
C49 B.n21 VSUBS 0.010757f
C50 B.n22 VSUBS 0.010757f
C51 B.n23 VSUBS 0.010757f
C52 B.n24 VSUBS 0.010757f
C53 B.n25 VSUBS 0.010757f
C54 B.n26 VSUBS 0.010757f
C55 B.n27 VSUBS 0.010757f
C56 B.n28 VSUBS 0.010757f
C57 B.n29 VSUBS 0.010757f
C58 B.n30 VSUBS 0.010757f
C59 B.n31 VSUBS 0.010757f
C60 B.n32 VSUBS 0.010757f
C61 B.n33 VSUBS 0.010757f
C62 B.n34 VSUBS 0.010757f
C63 B.n35 VSUBS 0.010757f
C64 B.n36 VSUBS 0.010757f
C65 B.n37 VSUBS 0.010757f
C66 B.n38 VSUBS 0.010757f
C67 B.n39 VSUBS 0.010757f
C68 B.n40 VSUBS 0.023662f
C69 B.n41 VSUBS 0.010757f
C70 B.n42 VSUBS 0.010757f
C71 B.n43 VSUBS 0.010757f
C72 B.n44 VSUBS 0.010757f
C73 B.n45 VSUBS 0.010757f
C74 B.n46 VSUBS 0.010757f
C75 B.n47 VSUBS 0.010757f
C76 B.n48 VSUBS 0.010757f
C77 B.n49 VSUBS 0.010757f
C78 B.n50 VSUBS 0.010757f
C79 B.n51 VSUBS 0.010757f
C80 B.n52 VSUBS 0.010757f
C81 B.n53 VSUBS 0.010757f
C82 B.n54 VSUBS 0.007435f
C83 B.n55 VSUBS 0.010757f
C84 B.t10 VSUBS 0.173129f
C85 B.t11 VSUBS 0.228442f
C86 B.t9 VSUBS 1.91193f
C87 B.n56 VSUBS 0.374595f
C88 B.n57 VSUBS 0.282193f
C89 B.n58 VSUBS 0.024922f
C90 B.n59 VSUBS 0.010757f
C91 B.n60 VSUBS 0.010757f
C92 B.n61 VSUBS 0.010757f
C93 B.n62 VSUBS 0.010757f
C94 B.t7 VSUBS 0.173132f
C95 B.t8 VSUBS 0.228445f
C96 B.t6 VSUBS 1.91193f
C97 B.n63 VSUBS 0.374592f
C98 B.n64 VSUBS 0.28219f
C99 B.n65 VSUBS 0.010757f
C100 B.n66 VSUBS 0.010757f
C101 B.n67 VSUBS 0.010757f
C102 B.n68 VSUBS 0.010757f
C103 B.n69 VSUBS 0.010757f
C104 B.n70 VSUBS 0.010757f
C105 B.n71 VSUBS 0.010757f
C106 B.n72 VSUBS 0.010757f
C107 B.n73 VSUBS 0.010757f
C108 B.n74 VSUBS 0.010757f
C109 B.n75 VSUBS 0.010757f
C110 B.n76 VSUBS 0.010757f
C111 B.n77 VSUBS 0.010757f
C112 B.n78 VSUBS 0.023662f
C113 B.n79 VSUBS 0.010757f
C114 B.n80 VSUBS 0.010757f
C115 B.n81 VSUBS 0.010757f
C116 B.n82 VSUBS 0.010757f
C117 B.n83 VSUBS 0.010757f
C118 B.n84 VSUBS 0.010757f
C119 B.n85 VSUBS 0.010757f
C120 B.n86 VSUBS 0.010757f
C121 B.n87 VSUBS 0.010757f
C122 B.n88 VSUBS 0.010757f
C123 B.n89 VSUBS 0.010757f
C124 B.n90 VSUBS 0.010757f
C125 B.n91 VSUBS 0.010757f
C126 B.n92 VSUBS 0.010757f
C127 B.n93 VSUBS 0.010757f
C128 B.n94 VSUBS 0.010757f
C129 B.n95 VSUBS 0.010757f
C130 B.n96 VSUBS 0.010757f
C131 B.n97 VSUBS 0.010757f
C132 B.n98 VSUBS 0.010757f
C133 B.n99 VSUBS 0.010757f
C134 B.n100 VSUBS 0.010757f
C135 B.n101 VSUBS 0.010757f
C136 B.n102 VSUBS 0.010757f
C137 B.n103 VSUBS 0.010757f
C138 B.n104 VSUBS 0.010757f
C139 B.n105 VSUBS 0.010757f
C140 B.n106 VSUBS 0.010757f
C141 B.n107 VSUBS 0.010757f
C142 B.n108 VSUBS 0.010757f
C143 B.n109 VSUBS 0.010757f
C144 B.n110 VSUBS 0.010757f
C145 B.n111 VSUBS 0.010757f
C146 B.n112 VSUBS 0.010757f
C147 B.n113 VSUBS 0.010757f
C148 B.n114 VSUBS 0.010757f
C149 B.n115 VSUBS 0.010757f
C150 B.n116 VSUBS 0.010757f
C151 B.n117 VSUBS 0.010757f
C152 B.n118 VSUBS 0.010757f
C153 B.n119 VSUBS 0.010757f
C154 B.n120 VSUBS 0.010757f
C155 B.n121 VSUBS 0.010757f
C156 B.n122 VSUBS 0.010757f
C157 B.n123 VSUBS 0.010757f
C158 B.n124 VSUBS 0.010757f
C159 B.n125 VSUBS 0.010757f
C160 B.n126 VSUBS 0.010757f
C161 B.n127 VSUBS 0.010757f
C162 B.n128 VSUBS 0.010757f
C163 B.n129 VSUBS 0.010757f
C164 B.n130 VSUBS 0.010757f
C165 B.n131 VSUBS 0.010757f
C166 B.n132 VSUBS 0.010757f
C167 B.n133 VSUBS 0.010757f
C168 B.n134 VSUBS 0.010757f
C169 B.n135 VSUBS 0.010757f
C170 B.n136 VSUBS 0.010757f
C171 B.n137 VSUBS 0.010757f
C172 B.n138 VSUBS 0.010757f
C173 B.n139 VSUBS 0.010757f
C174 B.n140 VSUBS 0.010757f
C175 B.n141 VSUBS 0.010757f
C176 B.n142 VSUBS 0.010757f
C177 B.n143 VSUBS 0.010757f
C178 B.n144 VSUBS 0.010757f
C179 B.n145 VSUBS 0.010757f
C180 B.n146 VSUBS 0.010757f
C181 B.n147 VSUBS 0.010757f
C182 B.n148 VSUBS 0.010757f
C183 B.n149 VSUBS 0.010757f
C184 B.n150 VSUBS 0.010757f
C185 B.n151 VSUBS 0.010757f
C186 B.n152 VSUBS 0.010757f
C187 B.n153 VSUBS 0.010757f
C188 B.n154 VSUBS 0.010757f
C189 B.n155 VSUBS 0.010757f
C190 B.n156 VSUBS 0.024426f
C191 B.n157 VSUBS 0.010757f
C192 B.n158 VSUBS 0.010757f
C193 B.n159 VSUBS 0.010757f
C194 B.n160 VSUBS 0.010757f
C195 B.n161 VSUBS 0.010757f
C196 B.n162 VSUBS 0.010757f
C197 B.n163 VSUBS 0.010757f
C198 B.n164 VSUBS 0.010757f
C199 B.n165 VSUBS 0.010757f
C200 B.n166 VSUBS 0.010757f
C201 B.n167 VSUBS 0.010757f
C202 B.n168 VSUBS 0.010757f
C203 B.n169 VSUBS 0.010757f
C204 B.n170 VSUBS 0.010757f
C205 B.t5 VSUBS 0.173132f
C206 B.t4 VSUBS 0.228445f
C207 B.t3 VSUBS 1.91193f
C208 B.n171 VSUBS 0.374592f
C209 B.n172 VSUBS 0.28219f
C210 B.n173 VSUBS 0.010757f
C211 B.n174 VSUBS 0.010757f
C212 B.n175 VSUBS 0.010757f
C213 B.n176 VSUBS 0.010757f
C214 B.t2 VSUBS 0.173129f
C215 B.t1 VSUBS 0.228442f
C216 B.t0 VSUBS 1.91193f
C217 B.n177 VSUBS 0.374595f
C218 B.n178 VSUBS 0.282193f
C219 B.n179 VSUBS 0.010757f
C220 B.n180 VSUBS 0.010757f
C221 B.n181 VSUBS 0.010757f
C222 B.n182 VSUBS 0.010757f
C223 B.n183 VSUBS 0.010757f
C224 B.n184 VSUBS 0.010757f
C225 B.n185 VSUBS 0.010757f
C226 B.n186 VSUBS 0.010757f
C227 B.n187 VSUBS 0.010757f
C228 B.n188 VSUBS 0.010757f
C229 B.n189 VSUBS 0.010757f
C230 B.n190 VSUBS 0.010757f
C231 B.n191 VSUBS 0.010757f
C232 B.n192 VSUBS 0.024426f
C233 B.n193 VSUBS 0.010757f
C234 B.n194 VSUBS 0.010757f
C235 B.n195 VSUBS 0.010757f
C236 B.n196 VSUBS 0.010757f
C237 B.n197 VSUBS 0.010757f
C238 B.n198 VSUBS 0.010757f
C239 B.n199 VSUBS 0.010757f
C240 B.n200 VSUBS 0.010757f
C241 B.n201 VSUBS 0.010757f
C242 B.n202 VSUBS 0.010757f
C243 B.n203 VSUBS 0.010757f
C244 B.n204 VSUBS 0.010757f
C245 B.n205 VSUBS 0.010757f
C246 B.n206 VSUBS 0.010757f
C247 B.n207 VSUBS 0.010757f
C248 B.n208 VSUBS 0.010757f
C249 B.n209 VSUBS 0.010757f
C250 B.n210 VSUBS 0.010757f
C251 B.n211 VSUBS 0.010757f
C252 B.n212 VSUBS 0.010757f
C253 B.n213 VSUBS 0.010757f
C254 B.n214 VSUBS 0.010757f
C255 B.n215 VSUBS 0.010757f
C256 B.n216 VSUBS 0.010757f
C257 B.n217 VSUBS 0.010757f
C258 B.n218 VSUBS 0.010757f
C259 B.n219 VSUBS 0.010757f
C260 B.n220 VSUBS 0.010757f
C261 B.n221 VSUBS 0.010757f
C262 B.n222 VSUBS 0.010757f
C263 B.n223 VSUBS 0.010757f
C264 B.n224 VSUBS 0.010757f
C265 B.n225 VSUBS 0.010757f
C266 B.n226 VSUBS 0.010757f
C267 B.n227 VSUBS 0.010757f
C268 B.n228 VSUBS 0.010757f
C269 B.n229 VSUBS 0.010757f
C270 B.n230 VSUBS 0.010757f
C271 B.n231 VSUBS 0.010757f
C272 B.n232 VSUBS 0.010757f
C273 B.n233 VSUBS 0.010757f
C274 B.n234 VSUBS 0.010757f
C275 B.n235 VSUBS 0.010757f
C276 B.n236 VSUBS 0.010757f
C277 B.n237 VSUBS 0.010757f
C278 B.n238 VSUBS 0.010757f
C279 B.n239 VSUBS 0.010757f
C280 B.n240 VSUBS 0.010757f
C281 B.n241 VSUBS 0.010757f
C282 B.n242 VSUBS 0.010757f
C283 B.n243 VSUBS 0.010757f
C284 B.n244 VSUBS 0.010757f
C285 B.n245 VSUBS 0.010757f
C286 B.n246 VSUBS 0.010757f
C287 B.n247 VSUBS 0.010757f
C288 B.n248 VSUBS 0.010757f
C289 B.n249 VSUBS 0.010757f
C290 B.n250 VSUBS 0.010757f
C291 B.n251 VSUBS 0.010757f
C292 B.n252 VSUBS 0.010757f
C293 B.n253 VSUBS 0.010757f
C294 B.n254 VSUBS 0.010757f
C295 B.n255 VSUBS 0.010757f
C296 B.n256 VSUBS 0.010757f
C297 B.n257 VSUBS 0.010757f
C298 B.n258 VSUBS 0.010757f
C299 B.n259 VSUBS 0.010757f
C300 B.n260 VSUBS 0.010757f
C301 B.n261 VSUBS 0.010757f
C302 B.n262 VSUBS 0.010757f
C303 B.n263 VSUBS 0.010757f
C304 B.n264 VSUBS 0.010757f
C305 B.n265 VSUBS 0.010757f
C306 B.n266 VSUBS 0.010757f
C307 B.n267 VSUBS 0.010757f
C308 B.n268 VSUBS 0.010757f
C309 B.n269 VSUBS 0.010757f
C310 B.n270 VSUBS 0.010757f
C311 B.n271 VSUBS 0.010757f
C312 B.n272 VSUBS 0.010757f
C313 B.n273 VSUBS 0.010757f
C314 B.n274 VSUBS 0.010757f
C315 B.n275 VSUBS 0.010757f
C316 B.n276 VSUBS 0.010757f
C317 B.n277 VSUBS 0.010757f
C318 B.n278 VSUBS 0.010757f
C319 B.n279 VSUBS 0.010757f
C320 B.n280 VSUBS 0.010757f
C321 B.n281 VSUBS 0.010757f
C322 B.n282 VSUBS 0.010757f
C323 B.n283 VSUBS 0.010757f
C324 B.n284 VSUBS 0.010757f
C325 B.n285 VSUBS 0.010757f
C326 B.n286 VSUBS 0.010757f
C327 B.n287 VSUBS 0.010757f
C328 B.n288 VSUBS 0.010757f
C329 B.n289 VSUBS 0.010757f
C330 B.n290 VSUBS 0.010757f
C331 B.n291 VSUBS 0.010757f
C332 B.n292 VSUBS 0.010757f
C333 B.n293 VSUBS 0.010757f
C334 B.n294 VSUBS 0.010757f
C335 B.n295 VSUBS 0.010757f
C336 B.n296 VSUBS 0.010757f
C337 B.n297 VSUBS 0.010757f
C338 B.n298 VSUBS 0.010757f
C339 B.n299 VSUBS 0.010757f
C340 B.n300 VSUBS 0.010757f
C341 B.n301 VSUBS 0.010757f
C342 B.n302 VSUBS 0.010757f
C343 B.n303 VSUBS 0.010757f
C344 B.n304 VSUBS 0.010757f
C345 B.n305 VSUBS 0.010757f
C346 B.n306 VSUBS 0.010757f
C347 B.n307 VSUBS 0.010757f
C348 B.n308 VSUBS 0.010757f
C349 B.n309 VSUBS 0.010757f
C350 B.n310 VSUBS 0.010757f
C351 B.n311 VSUBS 0.010757f
C352 B.n312 VSUBS 0.010757f
C353 B.n313 VSUBS 0.010757f
C354 B.n314 VSUBS 0.010757f
C355 B.n315 VSUBS 0.010757f
C356 B.n316 VSUBS 0.010757f
C357 B.n317 VSUBS 0.010757f
C358 B.n318 VSUBS 0.010757f
C359 B.n319 VSUBS 0.010757f
C360 B.n320 VSUBS 0.010757f
C361 B.n321 VSUBS 0.010757f
C362 B.n322 VSUBS 0.010757f
C363 B.n323 VSUBS 0.010757f
C364 B.n324 VSUBS 0.010757f
C365 B.n325 VSUBS 0.010757f
C366 B.n326 VSUBS 0.010757f
C367 B.n327 VSUBS 0.010757f
C368 B.n328 VSUBS 0.010757f
C369 B.n329 VSUBS 0.010757f
C370 B.n330 VSUBS 0.010757f
C371 B.n331 VSUBS 0.010757f
C372 B.n332 VSUBS 0.010757f
C373 B.n333 VSUBS 0.010757f
C374 B.n334 VSUBS 0.010757f
C375 B.n335 VSUBS 0.010757f
C376 B.n336 VSUBS 0.010757f
C377 B.n337 VSUBS 0.010757f
C378 B.n338 VSUBS 0.010757f
C379 B.n339 VSUBS 0.010757f
C380 B.n340 VSUBS 0.010757f
C381 B.n341 VSUBS 0.010757f
C382 B.n342 VSUBS 0.010757f
C383 B.n343 VSUBS 0.023662f
C384 B.n344 VSUBS 0.023662f
C385 B.n345 VSUBS 0.024426f
C386 B.n346 VSUBS 0.010757f
C387 B.n347 VSUBS 0.010757f
C388 B.n348 VSUBS 0.010757f
C389 B.n349 VSUBS 0.010757f
C390 B.n350 VSUBS 0.010757f
C391 B.n351 VSUBS 0.010757f
C392 B.n352 VSUBS 0.010757f
C393 B.n353 VSUBS 0.010757f
C394 B.n354 VSUBS 0.010757f
C395 B.n355 VSUBS 0.010757f
C396 B.n356 VSUBS 0.010757f
C397 B.n357 VSUBS 0.010757f
C398 B.n358 VSUBS 0.010757f
C399 B.n359 VSUBS 0.010757f
C400 B.n360 VSUBS 0.010757f
C401 B.n361 VSUBS 0.010757f
C402 B.n362 VSUBS 0.010757f
C403 B.n363 VSUBS 0.010757f
C404 B.n364 VSUBS 0.010757f
C405 B.n365 VSUBS 0.010757f
C406 B.n366 VSUBS 0.010757f
C407 B.n367 VSUBS 0.010757f
C408 B.n368 VSUBS 0.010757f
C409 B.n369 VSUBS 0.010757f
C410 B.n370 VSUBS 0.010757f
C411 B.n371 VSUBS 0.010757f
C412 B.n372 VSUBS 0.010757f
C413 B.n373 VSUBS 0.010757f
C414 B.n374 VSUBS 0.010757f
C415 B.n375 VSUBS 0.010757f
C416 B.n376 VSUBS 0.010757f
C417 B.n377 VSUBS 0.010757f
C418 B.n378 VSUBS 0.010757f
C419 B.n379 VSUBS 0.010757f
C420 B.n380 VSUBS 0.010757f
C421 B.n381 VSUBS 0.010757f
C422 B.n382 VSUBS 0.010757f
C423 B.n383 VSUBS 0.010757f
C424 B.n384 VSUBS 0.010757f
C425 B.n385 VSUBS 0.010757f
C426 B.n386 VSUBS 0.007435f
C427 B.n387 VSUBS 0.024922f
C428 B.n388 VSUBS 0.0087f
C429 B.n389 VSUBS 0.010757f
C430 B.n390 VSUBS 0.010757f
C431 B.n391 VSUBS 0.010757f
C432 B.n392 VSUBS 0.010757f
C433 B.n393 VSUBS 0.010757f
C434 B.n394 VSUBS 0.010757f
C435 B.n395 VSUBS 0.010757f
C436 B.n396 VSUBS 0.010757f
C437 B.n397 VSUBS 0.010757f
C438 B.n398 VSUBS 0.010757f
C439 B.n399 VSUBS 0.010757f
C440 B.n400 VSUBS 0.0087f
C441 B.n401 VSUBS 0.024922f
C442 B.n402 VSUBS 0.007435f
C443 B.n403 VSUBS 0.010757f
C444 B.n404 VSUBS 0.010757f
C445 B.n405 VSUBS 0.010757f
C446 B.n406 VSUBS 0.010757f
C447 B.n407 VSUBS 0.010757f
C448 B.n408 VSUBS 0.010757f
C449 B.n409 VSUBS 0.010757f
C450 B.n410 VSUBS 0.010757f
C451 B.n411 VSUBS 0.010757f
C452 B.n412 VSUBS 0.010757f
C453 B.n413 VSUBS 0.010757f
C454 B.n414 VSUBS 0.010757f
C455 B.n415 VSUBS 0.010757f
C456 B.n416 VSUBS 0.010757f
C457 B.n417 VSUBS 0.010757f
C458 B.n418 VSUBS 0.010757f
C459 B.n419 VSUBS 0.010757f
C460 B.n420 VSUBS 0.010757f
C461 B.n421 VSUBS 0.010757f
C462 B.n422 VSUBS 0.010757f
C463 B.n423 VSUBS 0.010757f
C464 B.n424 VSUBS 0.010757f
C465 B.n425 VSUBS 0.010757f
C466 B.n426 VSUBS 0.010757f
C467 B.n427 VSUBS 0.010757f
C468 B.n428 VSUBS 0.010757f
C469 B.n429 VSUBS 0.010757f
C470 B.n430 VSUBS 0.010757f
C471 B.n431 VSUBS 0.010757f
C472 B.n432 VSUBS 0.010757f
C473 B.n433 VSUBS 0.010757f
C474 B.n434 VSUBS 0.010757f
C475 B.n435 VSUBS 0.010757f
C476 B.n436 VSUBS 0.010757f
C477 B.n437 VSUBS 0.010757f
C478 B.n438 VSUBS 0.010757f
C479 B.n439 VSUBS 0.010757f
C480 B.n440 VSUBS 0.010757f
C481 B.n441 VSUBS 0.010757f
C482 B.n442 VSUBS 0.010757f
C483 B.n443 VSUBS 0.023063f
C484 B.n444 VSUBS 0.025025f
C485 B.n445 VSUBS 0.023662f
C486 B.n446 VSUBS 0.010757f
C487 B.n447 VSUBS 0.010757f
C488 B.n448 VSUBS 0.010757f
C489 B.n449 VSUBS 0.010757f
C490 B.n450 VSUBS 0.010757f
C491 B.n451 VSUBS 0.010757f
C492 B.n452 VSUBS 0.010757f
C493 B.n453 VSUBS 0.010757f
C494 B.n454 VSUBS 0.010757f
C495 B.n455 VSUBS 0.010757f
C496 B.n456 VSUBS 0.010757f
C497 B.n457 VSUBS 0.010757f
C498 B.n458 VSUBS 0.010757f
C499 B.n459 VSUBS 0.010757f
C500 B.n460 VSUBS 0.010757f
C501 B.n461 VSUBS 0.010757f
C502 B.n462 VSUBS 0.010757f
C503 B.n463 VSUBS 0.010757f
C504 B.n464 VSUBS 0.010757f
C505 B.n465 VSUBS 0.010757f
C506 B.n466 VSUBS 0.010757f
C507 B.n467 VSUBS 0.010757f
C508 B.n468 VSUBS 0.010757f
C509 B.n469 VSUBS 0.010757f
C510 B.n470 VSUBS 0.010757f
C511 B.n471 VSUBS 0.010757f
C512 B.n472 VSUBS 0.010757f
C513 B.n473 VSUBS 0.010757f
C514 B.n474 VSUBS 0.010757f
C515 B.n475 VSUBS 0.010757f
C516 B.n476 VSUBS 0.010757f
C517 B.n477 VSUBS 0.010757f
C518 B.n478 VSUBS 0.010757f
C519 B.n479 VSUBS 0.010757f
C520 B.n480 VSUBS 0.010757f
C521 B.n481 VSUBS 0.010757f
C522 B.n482 VSUBS 0.010757f
C523 B.n483 VSUBS 0.010757f
C524 B.n484 VSUBS 0.010757f
C525 B.n485 VSUBS 0.010757f
C526 B.n486 VSUBS 0.010757f
C527 B.n487 VSUBS 0.010757f
C528 B.n488 VSUBS 0.010757f
C529 B.n489 VSUBS 0.010757f
C530 B.n490 VSUBS 0.010757f
C531 B.n491 VSUBS 0.010757f
C532 B.n492 VSUBS 0.010757f
C533 B.n493 VSUBS 0.010757f
C534 B.n494 VSUBS 0.010757f
C535 B.n495 VSUBS 0.010757f
C536 B.n496 VSUBS 0.010757f
C537 B.n497 VSUBS 0.010757f
C538 B.n498 VSUBS 0.010757f
C539 B.n499 VSUBS 0.010757f
C540 B.n500 VSUBS 0.010757f
C541 B.n501 VSUBS 0.010757f
C542 B.n502 VSUBS 0.010757f
C543 B.n503 VSUBS 0.010757f
C544 B.n504 VSUBS 0.010757f
C545 B.n505 VSUBS 0.010757f
C546 B.n506 VSUBS 0.010757f
C547 B.n507 VSUBS 0.010757f
C548 B.n508 VSUBS 0.010757f
C549 B.n509 VSUBS 0.010757f
C550 B.n510 VSUBS 0.010757f
C551 B.n511 VSUBS 0.010757f
C552 B.n512 VSUBS 0.010757f
C553 B.n513 VSUBS 0.010757f
C554 B.n514 VSUBS 0.010757f
C555 B.n515 VSUBS 0.010757f
C556 B.n516 VSUBS 0.010757f
C557 B.n517 VSUBS 0.010757f
C558 B.n518 VSUBS 0.010757f
C559 B.n519 VSUBS 0.010757f
C560 B.n520 VSUBS 0.010757f
C561 B.n521 VSUBS 0.010757f
C562 B.n522 VSUBS 0.010757f
C563 B.n523 VSUBS 0.010757f
C564 B.n524 VSUBS 0.010757f
C565 B.n525 VSUBS 0.010757f
C566 B.n526 VSUBS 0.010757f
C567 B.n527 VSUBS 0.010757f
C568 B.n528 VSUBS 0.010757f
C569 B.n529 VSUBS 0.010757f
C570 B.n530 VSUBS 0.010757f
C571 B.n531 VSUBS 0.010757f
C572 B.n532 VSUBS 0.010757f
C573 B.n533 VSUBS 0.010757f
C574 B.n534 VSUBS 0.010757f
C575 B.n535 VSUBS 0.010757f
C576 B.n536 VSUBS 0.010757f
C577 B.n537 VSUBS 0.010757f
C578 B.n538 VSUBS 0.010757f
C579 B.n539 VSUBS 0.010757f
C580 B.n540 VSUBS 0.010757f
C581 B.n541 VSUBS 0.010757f
C582 B.n542 VSUBS 0.010757f
C583 B.n543 VSUBS 0.010757f
C584 B.n544 VSUBS 0.010757f
C585 B.n545 VSUBS 0.010757f
C586 B.n546 VSUBS 0.010757f
C587 B.n547 VSUBS 0.010757f
C588 B.n548 VSUBS 0.010757f
C589 B.n549 VSUBS 0.010757f
C590 B.n550 VSUBS 0.010757f
C591 B.n551 VSUBS 0.010757f
C592 B.n552 VSUBS 0.010757f
C593 B.n553 VSUBS 0.010757f
C594 B.n554 VSUBS 0.010757f
C595 B.n555 VSUBS 0.010757f
C596 B.n556 VSUBS 0.010757f
C597 B.n557 VSUBS 0.010757f
C598 B.n558 VSUBS 0.010757f
C599 B.n559 VSUBS 0.010757f
C600 B.n560 VSUBS 0.010757f
C601 B.n561 VSUBS 0.010757f
C602 B.n562 VSUBS 0.010757f
C603 B.n563 VSUBS 0.010757f
C604 B.n564 VSUBS 0.010757f
C605 B.n565 VSUBS 0.010757f
C606 B.n566 VSUBS 0.010757f
C607 B.n567 VSUBS 0.010757f
C608 B.n568 VSUBS 0.010757f
C609 B.n569 VSUBS 0.010757f
C610 B.n570 VSUBS 0.010757f
C611 B.n571 VSUBS 0.010757f
C612 B.n572 VSUBS 0.010757f
C613 B.n573 VSUBS 0.010757f
C614 B.n574 VSUBS 0.010757f
C615 B.n575 VSUBS 0.010757f
C616 B.n576 VSUBS 0.010757f
C617 B.n577 VSUBS 0.010757f
C618 B.n578 VSUBS 0.010757f
C619 B.n579 VSUBS 0.010757f
C620 B.n580 VSUBS 0.010757f
C621 B.n581 VSUBS 0.010757f
C622 B.n582 VSUBS 0.010757f
C623 B.n583 VSUBS 0.010757f
C624 B.n584 VSUBS 0.010757f
C625 B.n585 VSUBS 0.010757f
C626 B.n586 VSUBS 0.010757f
C627 B.n587 VSUBS 0.010757f
C628 B.n588 VSUBS 0.010757f
C629 B.n589 VSUBS 0.010757f
C630 B.n590 VSUBS 0.010757f
C631 B.n591 VSUBS 0.010757f
C632 B.n592 VSUBS 0.010757f
C633 B.n593 VSUBS 0.010757f
C634 B.n594 VSUBS 0.010757f
C635 B.n595 VSUBS 0.010757f
C636 B.n596 VSUBS 0.010757f
C637 B.n597 VSUBS 0.010757f
C638 B.n598 VSUBS 0.010757f
C639 B.n599 VSUBS 0.010757f
C640 B.n600 VSUBS 0.010757f
C641 B.n601 VSUBS 0.010757f
C642 B.n602 VSUBS 0.010757f
C643 B.n603 VSUBS 0.010757f
C644 B.n604 VSUBS 0.010757f
C645 B.n605 VSUBS 0.010757f
C646 B.n606 VSUBS 0.010757f
C647 B.n607 VSUBS 0.010757f
C648 B.n608 VSUBS 0.010757f
C649 B.n609 VSUBS 0.010757f
C650 B.n610 VSUBS 0.010757f
C651 B.n611 VSUBS 0.010757f
C652 B.n612 VSUBS 0.010757f
C653 B.n613 VSUBS 0.010757f
C654 B.n614 VSUBS 0.010757f
C655 B.n615 VSUBS 0.010757f
C656 B.n616 VSUBS 0.010757f
C657 B.n617 VSUBS 0.010757f
C658 B.n618 VSUBS 0.010757f
C659 B.n619 VSUBS 0.010757f
C660 B.n620 VSUBS 0.010757f
C661 B.n621 VSUBS 0.010757f
C662 B.n622 VSUBS 0.010757f
C663 B.n623 VSUBS 0.010757f
C664 B.n624 VSUBS 0.010757f
C665 B.n625 VSUBS 0.010757f
C666 B.n626 VSUBS 0.010757f
C667 B.n627 VSUBS 0.010757f
C668 B.n628 VSUBS 0.010757f
C669 B.n629 VSUBS 0.010757f
C670 B.n630 VSUBS 0.010757f
C671 B.n631 VSUBS 0.010757f
C672 B.n632 VSUBS 0.010757f
C673 B.n633 VSUBS 0.010757f
C674 B.n634 VSUBS 0.010757f
C675 B.n635 VSUBS 0.010757f
C676 B.n636 VSUBS 0.010757f
C677 B.n637 VSUBS 0.010757f
C678 B.n638 VSUBS 0.010757f
C679 B.n639 VSUBS 0.010757f
C680 B.n640 VSUBS 0.010757f
C681 B.n641 VSUBS 0.010757f
C682 B.n642 VSUBS 0.010757f
C683 B.n643 VSUBS 0.010757f
C684 B.n644 VSUBS 0.010757f
C685 B.n645 VSUBS 0.010757f
C686 B.n646 VSUBS 0.010757f
C687 B.n647 VSUBS 0.010757f
C688 B.n648 VSUBS 0.010757f
C689 B.n649 VSUBS 0.010757f
C690 B.n650 VSUBS 0.010757f
C691 B.n651 VSUBS 0.010757f
C692 B.n652 VSUBS 0.010757f
C693 B.n653 VSUBS 0.010757f
C694 B.n654 VSUBS 0.010757f
C695 B.n655 VSUBS 0.010757f
C696 B.n656 VSUBS 0.010757f
C697 B.n657 VSUBS 0.010757f
C698 B.n658 VSUBS 0.010757f
C699 B.n659 VSUBS 0.010757f
C700 B.n660 VSUBS 0.010757f
C701 B.n661 VSUBS 0.010757f
C702 B.n662 VSUBS 0.010757f
C703 B.n663 VSUBS 0.010757f
C704 B.n664 VSUBS 0.010757f
C705 B.n665 VSUBS 0.010757f
C706 B.n666 VSUBS 0.010757f
C707 B.n667 VSUBS 0.010757f
C708 B.n668 VSUBS 0.010757f
C709 B.n669 VSUBS 0.010757f
C710 B.n670 VSUBS 0.010757f
C711 B.n671 VSUBS 0.010757f
C712 B.n672 VSUBS 0.010757f
C713 B.n673 VSUBS 0.010757f
C714 B.n674 VSUBS 0.010757f
C715 B.n675 VSUBS 0.010757f
C716 B.n676 VSUBS 0.010757f
C717 B.n677 VSUBS 0.023662f
C718 B.n678 VSUBS 0.024426f
C719 B.n679 VSUBS 0.024426f
C720 B.n680 VSUBS 0.010757f
C721 B.n681 VSUBS 0.010757f
C722 B.n682 VSUBS 0.010757f
C723 B.n683 VSUBS 0.010757f
C724 B.n684 VSUBS 0.010757f
C725 B.n685 VSUBS 0.010757f
C726 B.n686 VSUBS 0.010757f
C727 B.n687 VSUBS 0.010757f
C728 B.n688 VSUBS 0.010757f
C729 B.n689 VSUBS 0.010757f
C730 B.n690 VSUBS 0.010757f
C731 B.n691 VSUBS 0.010757f
C732 B.n692 VSUBS 0.010757f
C733 B.n693 VSUBS 0.010757f
C734 B.n694 VSUBS 0.010757f
C735 B.n695 VSUBS 0.010757f
C736 B.n696 VSUBS 0.010757f
C737 B.n697 VSUBS 0.010757f
C738 B.n698 VSUBS 0.010757f
C739 B.n699 VSUBS 0.010757f
C740 B.n700 VSUBS 0.010757f
C741 B.n701 VSUBS 0.010757f
C742 B.n702 VSUBS 0.010757f
C743 B.n703 VSUBS 0.010757f
C744 B.n704 VSUBS 0.010757f
C745 B.n705 VSUBS 0.010757f
C746 B.n706 VSUBS 0.010757f
C747 B.n707 VSUBS 0.010757f
C748 B.n708 VSUBS 0.010757f
C749 B.n709 VSUBS 0.010757f
C750 B.n710 VSUBS 0.010757f
C751 B.n711 VSUBS 0.010757f
C752 B.n712 VSUBS 0.010757f
C753 B.n713 VSUBS 0.010757f
C754 B.n714 VSUBS 0.010757f
C755 B.n715 VSUBS 0.010757f
C756 B.n716 VSUBS 0.010757f
C757 B.n717 VSUBS 0.010757f
C758 B.n718 VSUBS 0.010757f
C759 B.n719 VSUBS 0.007435f
C760 B.n720 VSUBS 0.024922f
C761 B.n721 VSUBS 0.0087f
C762 B.n722 VSUBS 0.010757f
C763 B.n723 VSUBS 0.010757f
C764 B.n724 VSUBS 0.010757f
C765 B.n725 VSUBS 0.010757f
C766 B.n726 VSUBS 0.010757f
C767 B.n727 VSUBS 0.010757f
C768 B.n728 VSUBS 0.010757f
C769 B.n729 VSUBS 0.010757f
C770 B.n730 VSUBS 0.010757f
C771 B.n731 VSUBS 0.010757f
C772 B.n732 VSUBS 0.010757f
C773 B.n733 VSUBS 0.0087f
C774 B.n734 VSUBS 0.010757f
C775 B.n735 VSUBS 0.010757f
C776 B.n736 VSUBS 0.010757f
C777 B.n737 VSUBS 0.010757f
C778 B.n738 VSUBS 0.010757f
C779 B.n739 VSUBS 0.010757f
C780 B.n740 VSUBS 0.010757f
C781 B.n741 VSUBS 0.010757f
C782 B.n742 VSUBS 0.010757f
C783 B.n743 VSUBS 0.010757f
C784 B.n744 VSUBS 0.010757f
C785 B.n745 VSUBS 0.010757f
C786 B.n746 VSUBS 0.010757f
C787 B.n747 VSUBS 0.010757f
C788 B.n748 VSUBS 0.010757f
C789 B.n749 VSUBS 0.010757f
C790 B.n750 VSUBS 0.010757f
C791 B.n751 VSUBS 0.010757f
C792 B.n752 VSUBS 0.010757f
C793 B.n753 VSUBS 0.010757f
C794 B.n754 VSUBS 0.010757f
C795 B.n755 VSUBS 0.010757f
C796 B.n756 VSUBS 0.010757f
C797 B.n757 VSUBS 0.010757f
C798 B.n758 VSUBS 0.010757f
C799 B.n759 VSUBS 0.010757f
C800 B.n760 VSUBS 0.010757f
C801 B.n761 VSUBS 0.010757f
C802 B.n762 VSUBS 0.010757f
C803 B.n763 VSUBS 0.010757f
C804 B.n764 VSUBS 0.010757f
C805 B.n765 VSUBS 0.010757f
C806 B.n766 VSUBS 0.010757f
C807 B.n767 VSUBS 0.010757f
C808 B.n768 VSUBS 0.010757f
C809 B.n769 VSUBS 0.010757f
C810 B.n770 VSUBS 0.010757f
C811 B.n771 VSUBS 0.010757f
C812 B.n772 VSUBS 0.010757f
C813 B.n773 VSUBS 0.010757f
C814 B.n774 VSUBS 0.010757f
C815 B.n775 VSUBS 0.024426f
C816 B.n776 VSUBS 0.024426f
C817 B.n777 VSUBS 0.023662f
C818 B.n778 VSUBS 0.010757f
C819 B.n779 VSUBS 0.010757f
C820 B.n780 VSUBS 0.010757f
C821 B.n781 VSUBS 0.010757f
C822 B.n782 VSUBS 0.010757f
C823 B.n783 VSUBS 0.010757f
C824 B.n784 VSUBS 0.010757f
C825 B.n785 VSUBS 0.010757f
C826 B.n786 VSUBS 0.010757f
C827 B.n787 VSUBS 0.010757f
C828 B.n788 VSUBS 0.010757f
C829 B.n789 VSUBS 0.010757f
C830 B.n790 VSUBS 0.010757f
C831 B.n791 VSUBS 0.010757f
C832 B.n792 VSUBS 0.010757f
C833 B.n793 VSUBS 0.010757f
C834 B.n794 VSUBS 0.010757f
C835 B.n795 VSUBS 0.010757f
C836 B.n796 VSUBS 0.010757f
C837 B.n797 VSUBS 0.010757f
C838 B.n798 VSUBS 0.010757f
C839 B.n799 VSUBS 0.010757f
C840 B.n800 VSUBS 0.010757f
C841 B.n801 VSUBS 0.010757f
C842 B.n802 VSUBS 0.010757f
C843 B.n803 VSUBS 0.010757f
C844 B.n804 VSUBS 0.010757f
C845 B.n805 VSUBS 0.010757f
C846 B.n806 VSUBS 0.010757f
C847 B.n807 VSUBS 0.010757f
C848 B.n808 VSUBS 0.010757f
C849 B.n809 VSUBS 0.010757f
C850 B.n810 VSUBS 0.010757f
C851 B.n811 VSUBS 0.010757f
C852 B.n812 VSUBS 0.010757f
C853 B.n813 VSUBS 0.010757f
C854 B.n814 VSUBS 0.010757f
C855 B.n815 VSUBS 0.010757f
C856 B.n816 VSUBS 0.010757f
C857 B.n817 VSUBS 0.010757f
C858 B.n818 VSUBS 0.010757f
C859 B.n819 VSUBS 0.010757f
C860 B.n820 VSUBS 0.010757f
C861 B.n821 VSUBS 0.010757f
C862 B.n822 VSUBS 0.010757f
C863 B.n823 VSUBS 0.010757f
C864 B.n824 VSUBS 0.010757f
C865 B.n825 VSUBS 0.010757f
C866 B.n826 VSUBS 0.010757f
C867 B.n827 VSUBS 0.010757f
C868 B.n828 VSUBS 0.010757f
C869 B.n829 VSUBS 0.010757f
C870 B.n830 VSUBS 0.010757f
C871 B.n831 VSUBS 0.010757f
C872 B.n832 VSUBS 0.010757f
C873 B.n833 VSUBS 0.010757f
C874 B.n834 VSUBS 0.010757f
C875 B.n835 VSUBS 0.010757f
C876 B.n836 VSUBS 0.010757f
C877 B.n837 VSUBS 0.010757f
C878 B.n838 VSUBS 0.010757f
C879 B.n839 VSUBS 0.010757f
C880 B.n840 VSUBS 0.010757f
C881 B.n841 VSUBS 0.010757f
C882 B.n842 VSUBS 0.010757f
C883 B.n843 VSUBS 0.010757f
C884 B.n844 VSUBS 0.010757f
C885 B.n845 VSUBS 0.010757f
C886 B.n846 VSUBS 0.010757f
C887 B.n847 VSUBS 0.010757f
C888 B.n848 VSUBS 0.010757f
C889 B.n849 VSUBS 0.010757f
C890 B.n850 VSUBS 0.010757f
C891 B.n851 VSUBS 0.010757f
C892 B.n852 VSUBS 0.010757f
C893 B.n853 VSUBS 0.010757f
C894 B.n854 VSUBS 0.010757f
C895 B.n855 VSUBS 0.010757f
C896 B.n856 VSUBS 0.010757f
C897 B.n857 VSUBS 0.010757f
C898 B.n858 VSUBS 0.010757f
C899 B.n859 VSUBS 0.010757f
C900 B.n860 VSUBS 0.010757f
C901 B.n861 VSUBS 0.010757f
C902 B.n862 VSUBS 0.010757f
C903 B.n863 VSUBS 0.010757f
C904 B.n864 VSUBS 0.010757f
C905 B.n865 VSUBS 0.010757f
C906 B.n866 VSUBS 0.010757f
C907 B.n867 VSUBS 0.010757f
C908 B.n868 VSUBS 0.010757f
C909 B.n869 VSUBS 0.010757f
C910 B.n870 VSUBS 0.010757f
C911 B.n871 VSUBS 0.010757f
C912 B.n872 VSUBS 0.010757f
C913 B.n873 VSUBS 0.010757f
C914 B.n874 VSUBS 0.010757f
C915 B.n875 VSUBS 0.010757f
C916 B.n876 VSUBS 0.010757f
C917 B.n877 VSUBS 0.010757f
C918 B.n878 VSUBS 0.010757f
C919 B.n879 VSUBS 0.010757f
C920 B.n880 VSUBS 0.010757f
C921 B.n881 VSUBS 0.010757f
C922 B.n882 VSUBS 0.010757f
C923 B.n883 VSUBS 0.010757f
C924 B.n884 VSUBS 0.010757f
C925 B.n885 VSUBS 0.010757f
C926 B.n886 VSUBS 0.010757f
C927 B.n887 VSUBS 0.010757f
C928 B.n888 VSUBS 0.010757f
C929 B.n889 VSUBS 0.010757f
C930 B.n890 VSUBS 0.010757f
C931 B.n891 VSUBS 0.014037f
C932 B.n892 VSUBS 0.014953f
C933 B.n893 VSUBS 0.029735f
C934 VDD1.n0 VSUBS 0.037477f
C935 VDD1.n1 VSUBS 0.034001f
C936 VDD1.n2 VSUBS 0.018271f
C937 VDD1.n3 VSUBS 0.043185f
C938 VDD1.n4 VSUBS 0.019345f
C939 VDD1.n5 VSUBS 0.034001f
C940 VDD1.n6 VSUBS 0.018271f
C941 VDD1.n7 VSUBS 0.043185f
C942 VDD1.n8 VSUBS 0.019345f
C943 VDD1.n9 VSUBS 0.966857f
C944 VDD1.n10 VSUBS 0.018271f
C945 VDD1.t5 VSUBS 0.092804f
C946 VDD1.n11 VSUBS 0.19545f
C947 VDD1.n12 VSUBS 0.032484f
C948 VDD1.n13 VSUBS 0.032389f
C949 VDD1.n14 VSUBS 0.043185f
C950 VDD1.n15 VSUBS 0.019345f
C951 VDD1.n16 VSUBS 0.018271f
C952 VDD1.n17 VSUBS 0.034001f
C953 VDD1.n18 VSUBS 0.034001f
C954 VDD1.n19 VSUBS 0.018271f
C955 VDD1.n20 VSUBS 0.019345f
C956 VDD1.n21 VSUBS 0.043185f
C957 VDD1.n22 VSUBS 0.043185f
C958 VDD1.n23 VSUBS 0.019345f
C959 VDD1.n24 VSUBS 0.018271f
C960 VDD1.n25 VSUBS 0.034001f
C961 VDD1.n26 VSUBS 0.034001f
C962 VDD1.n27 VSUBS 0.018271f
C963 VDD1.n28 VSUBS 0.019345f
C964 VDD1.n29 VSUBS 0.043185f
C965 VDD1.n30 VSUBS 0.108818f
C966 VDD1.n31 VSUBS 0.019345f
C967 VDD1.n32 VSUBS 0.035879f
C968 VDD1.n33 VSUBS 0.08788f
C969 VDD1.n34 VSUBS 0.13415f
C970 VDD1.t8 VSUBS 0.195601f
C971 VDD1.t3 VSUBS 0.195601f
C972 VDD1.n35 VSUBS 1.39075f
C973 VDD1.n36 VSUBS 1.44057f
C974 VDD1.n37 VSUBS 0.037477f
C975 VDD1.n38 VSUBS 0.034001f
C976 VDD1.n39 VSUBS 0.018271f
C977 VDD1.n40 VSUBS 0.043185f
C978 VDD1.n41 VSUBS 0.019345f
C979 VDD1.n42 VSUBS 0.034001f
C980 VDD1.n43 VSUBS 0.018271f
C981 VDD1.n44 VSUBS 0.043185f
C982 VDD1.n45 VSUBS 0.019345f
C983 VDD1.n46 VSUBS 0.966857f
C984 VDD1.n47 VSUBS 0.018271f
C985 VDD1.t4 VSUBS 0.092804f
C986 VDD1.n48 VSUBS 0.19545f
C987 VDD1.n49 VSUBS 0.032484f
C988 VDD1.n50 VSUBS 0.032389f
C989 VDD1.n51 VSUBS 0.043185f
C990 VDD1.n52 VSUBS 0.019345f
C991 VDD1.n53 VSUBS 0.018271f
C992 VDD1.n54 VSUBS 0.034001f
C993 VDD1.n55 VSUBS 0.034001f
C994 VDD1.n56 VSUBS 0.018271f
C995 VDD1.n57 VSUBS 0.019345f
C996 VDD1.n58 VSUBS 0.043185f
C997 VDD1.n59 VSUBS 0.043185f
C998 VDD1.n60 VSUBS 0.019345f
C999 VDD1.n61 VSUBS 0.018271f
C1000 VDD1.n62 VSUBS 0.034001f
C1001 VDD1.n63 VSUBS 0.034001f
C1002 VDD1.n64 VSUBS 0.018271f
C1003 VDD1.n65 VSUBS 0.019345f
C1004 VDD1.n66 VSUBS 0.043185f
C1005 VDD1.n67 VSUBS 0.108818f
C1006 VDD1.n68 VSUBS 0.019345f
C1007 VDD1.n69 VSUBS 0.035879f
C1008 VDD1.n70 VSUBS 0.08788f
C1009 VDD1.n71 VSUBS 0.13415f
C1010 VDD1.t9 VSUBS 0.195601f
C1011 VDD1.t0 VSUBS 0.195601f
C1012 VDD1.n72 VSUBS 1.39074f
C1013 VDD1.n73 VSUBS 1.42914f
C1014 VDD1.t1 VSUBS 0.195601f
C1015 VDD1.t6 VSUBS 0.195601f
C1016 VDD1.n74 VSUBS 1.42371f
C1017 VDD1.n75 VSUBS 4.73708f
C1018 VDD1.t7 VSUBS 0.195601f
C1019 VDD1.t2 VSUBS 0.195601f
C1020 VDD1.n76 VSUBS 1.39074f
C1021 VDD1.n77 VSUBS 4.661f
C1022 VP.t3 VSUBS 2.23117f
C1023 VP.n0 VSUBS 0.923888f
C1024 VP.n1 VSUBS 0.031924f
C1025 VP.n2 VSUBS 0.056373f
C1026 VP.n3 VSUBS 0.031924f
C1027 VP.n4 VSUBS 0.049264f
C1028 VP.n5 VSUBS 0.031924f
C1029 VP.n6 VSUBS 0.04994f
C1030 VP.n7 VSUBS 0.031924f
C1031 VP.n8 VSUBS 0.044588f
C1032 VP.n9 VSUBS 0.031924f
C1033 VP.n10 VSUBS 0.042874f
C1034 VP.n11 VSUBS 0.031924f
C1035 VP.n12 VSUBS 0.039912f
C1036 VP.n13 VSUBS 0.031924f
C1037 VP.n14 VSUBS 0.033395f
C1038 VP.n15 VSUBS 0.031924f
C1039 VP.n16 VSUBS 0.035236f
C1040 VP.t7 VSUBS 2.23117f
C1041 VP.n17 VSUBS 0.923888f
C1042 VP.n18 VSUBS 0.031924f
C1043 VP.n19 VSUBS 0.056373f
C1044 VP.n20 VSUBS 0.031924f
C1045 VP.n21 VSUBS 0.049264f
C1046 VP.n22 VSUBS 0.031924f
C1047 VP.n23 VSUBS 0.04994f
C1048 VP.n24 VSUBS 0.031924f
C1049 VP.n25 VSUBS 0.044588f
C1050 VP.n26 VSUBS 0.031924f
C1051 VP.n27 VSUBS 0.042874f
C1052 VP.n28 VSUBS 0.031924f
C1053 VP.n29 VSUBS 0.039912f
C1054 VP.t4 VSUBS 2.64817f
C1055 VP.t1 VSUBS 2.23117f
C1056 VP.n30 VSUBS 0.914396f
C1057 VP.n31 VSUBS 0.87627f
C1058 VP.n32 VSUBS 0.400249f
C1059 VP.n33 VSUBS 0.031924f
C1060 VP.n34 VSUBS 0.059201f
C1061 VP.n35 VSUBS 0.059201f
C1062 VP.n36 VSUBS 0.04994f
C1063 VP.n37 VSUBS 0.031924f
C1064 VP.n38 VSUBS 0.031924f
C1065 VP.n39 VSUBS 0.031924f
C1066 VP.n40 VSUBS 0.059201f
C1067 VP.n41 VSUBS 0.059201f
C1068 VP.t6 VSUBS 2.23117f
C1069 VP.n42 VSUBS 0.808637f
C1070 VP.n43 VSUBS 0.044588f
C1071 VP.n44 VSUBS 0.031924f
C1072 VP.n45 VSUBS 0.031924f
C1073 VP.n46 VSUBS 0.031924f
C1074 VP.n47 VSUBS 0.059201f
C1075 VP.n48 VSUBS 0.059201f
C1076 VP.n49 VSUBS 0.042874f
C1077 VP.n50 VSUBS 0.031924f
C1078 VP.n51 VSUBS 0.031924f
C1079 VP.n52 VSUBS 0.031924f
C1080 VP.n53 VSUBS 0.059201f
C1081 VP.n54 VSUBS 0.059201f
C1082 VP.t2 VSUBS 2.23117f
C1083 VP.n55 VSUBS 0.808637f
C1084 VP.n56 VSUBS 0.039912f
C1085 VP.n57 VSUBS 0.031924f
C1086 VP.n58 VSUBS 0.031924f
C1087 VP.n59 VSUBS 0.031924f
C1088 VP.n60 VSUBS 0.059201f
C1089 VP.n61 VSUBS 0.062246f
C1090 VP.n62 VSUBS 0.033395f
C1091 VP.n63 VSUBS 0.031924f
C1092 VP.n64 VSUBS 0.031924f
C1093 VP.n65 VSUBS 0.031924f
C1094 VP.n66 VSUBS 0.059201f
C1095 VP.n67 VSUBS 0.059201f
C1096 VP.n68 VSUBS 0.035236f
C1097 VP.n69 VSUBS 0.051517f
C1098 VP.n70 VSUBS 2.0884f
C1099 VP.t5 VSUBS 2.23117f
C1100 VP.n71 VSUBS 0.923888f
C1101 VP.n72 VSUBS 2.10934f
C1102 VP.n73 VSUBS 0.051517f
C1103 VP.n74 VSUBS 0.031924f
C1104 VP.n75 VSUBS 0.059201f
C1105 VP.n76 VSUBS 0.059201f
C1106 VP.n77 VSUBS 0.056373f
C1107 VP.n78 VSUBS 0.031924f
C1108 VP.n79 VSUBS 0.031924f
C1109 VP.n80 VSUBS 0.031924f
C1110 VP.n81 VSUBS 0.062246f
C1111 VP.n82 VSUBS 0.059201f
C1112 VP.t0 VSUBS 2.23117f
C1113 VP.n83 VSUBS 0.808637f
C1114 VP.n84 VSUBS 0.049264f
C1115 VP.n85 VSUBS 0.031924f
C1116 VP.n86 VSUBS 0.031924f
C1117 VP.n87 VSUBS 0.031924f
C1118 VP.n88 VSUBS 0.059201f
C1119 VP.n89 VSUBS 0.059201f
C1120 VP.n90 VSUBS 0.04994f
C1121 VP.n91 VSUBS 0.031924f
C1122 VP.n92 VSUBS 0.031924f
C1123 VP.n93 VSUBS 0.031924f
C1124 VP.n94 VSUBS 0.059201f
C1125 VP.n95 VSUBS 0.059201f
C1126 VP.t9 VSUBS 2.23117f
C1127 VP.n96 VSUBS 0.808637f
C1128 VP.n97 VSUBS 0.044588f
C1129 VP.n98 VSUBS 0.031924f
C1130 VP.n99 VSUBS 0.031924f
C1131 VP.n100 VSUBS 0.031924f
C1132 VP.n101 VSUBS 0.059201f
C1133 VP.n102 VSUBS 0.059201f
C1134 VP.n103 VSUBS 0.042874f
C1135 VP.n104 VSUBS 0.031924f
C1136 VP.n105 VSUBS 0.031924f
C1137 VP.n106 VSUBS 0.031924f
C1138 VP.n107 VSUBS 0.059201f
C1139 VP.n108 VSUBS 0.059201f
C1140 VP.t8 VSUBS 2.23117f
C1141 VP.n109 VSUBS 0.808637f
C1142 VP.n110 VSUBS 0.039912f
C1143 VP.n111 VSUBS 0.031924f
C1144 VP.n112 VSUBS 0.031924f
C1145 VP.n113 VSUBS 0.031924f
C1146 VP.n114 VSUBS 0.059201f
C1147 VP.n115 VSUBS 0.062246f
C1148 VP.n116 VSUBS 0.033395f
C1149 VP.n117 VSUBS 0.031924f
C1150 VP.n118 VSUBS 0.031924f
C1151 VP.n119 VSUBS 0.031924f
C1152 VP.n120 VSUBS 0.059201f
C1153 VP.n121 VSUBS 0.059201f
C1154 VP.n122 VSUBS 0.035236f
C1155 VP.n123 VSUBS 0.051517f
C1156 VP.n124 VSUBS 0.092844f
C1157 VDD2.n0 VSUBS 0.037363f
C1158 VDD2.n1 VSUBS 0.033898f
C1159 VDD2.n2 VSUBS 0.018215f
C1160 VDD2.n3 VSUBS 0.043054f
C1161 VDD2.n4 VSUBS 0.019287f
C1162 VDD2.n5 VSUBS 0.033898f
C1163 VDD2.n6 VSUBS 0.018215f
C1164 VDD2.n7 VSUBS 0.043054f
C1165 VDD2.n8 VSUBS 0.019287f
C1166 VDD2.n9 VSUBS 0.963929f
C1167 VDD2.n10 VSUBS 0.018215f
C1168 VDD2.t4 VSUBS 0.092523f
C1169 VDD2.n11 VSUBS 0.194858f
C1170 VDD2.n12 VSUBS 0.032386f
C1171 VDD2.n13 VSUBS 0.03229f
C1172 VDD2.n14 VSUBS 0.043054f
C1173 VDD2.n15 VSUBS 0.019287f
C1174 VDD2.n16 VSUBS 0.018215f
C1175 VDD2.n17 VSUBS 0.033898f
C1176 VDD2.n18 VSUBS 0.033898f
C1177 VDD2.n19 VSUBS 0.018215f
C1178 VDD2.n20 VSUBS 0.019287f
C1179 VDD2.n21 VSUBS 0.043054f
C1180 VDD2.n22 VSUBS 0.043054f
C1181 VDD2.n23 VSUBS 0.019287f
C1182 VDD2.n24 VSUBS 0.018215f
C1183 VDD2.n25 VSUBS 0.033898f
C1184 VDD2.n26 VSUBS 0.033898f
C1185 VDD2.n27 VSUBS 0.018215f
C1186 VDD2.n28 VSUBS 0.019287f
C1187 VDD2.n29 VSUBS 0.043054f
C1188 VDD2.n30 VSUBS 0.108489f
C1189 VDD2.n31 VSUBS 0.019287f
C1190 VDD2.n32 VSUBS 0.03577f
C1191 VDD2.n33 VSUBS 0.087614f
C1192 VDD2.n34 VSUBS 0.133744f
C1193 VDD2.t0 VSUBS 0.195009f
C1194 VDD2.t9 VSUBS 0.195009f
C1195 VDD2.n35 VSUBS 1.38653f
C1196 VDD2.n36 VSUBS 1.42481f
C1197 VDD2.t6 VSUBS 0.195009f
C1198 VDD2.t1 VSUBS 0.195009f
C1199 VDD2.n37 VSUBS 1.4194f
C1200 VDD2.n38 VSUBS 4.52192f
C1201 VDD2.n39 VSUBS 0.037363f
C1202 VDD2.n40 VSUBS 0.033898f
C1203 VDD2.n41 VSUBS 0.018215f
C1204 VDD2.n42 VSUBS 0.043054f
C1205 VDD2.n43 VSUBS 0.019287f
C1206 VDD2.n44 VSUBS 0.033898f
C1207 VDD2.n45 VSUBS 0.018215f
C1208 VDD2.n46 VSUBS 0.043054f
C1209 VDD2.n47 VSUBS 0.019287f
C1210 VDD2.n48 VSUBS 0.963929f
C1211 VDD2.n49 VSUBS 0.018215f
C1212 VDD2.t8 VSUBS 0.092523f
C1213 VDD2.n50 VSUBS 0.194858f
C1214 VDD2.n51 VSUBS 0.032386f
C1215 VDD2.n52 VSUBS 0.03229f
C1216 VDD2.n53 VSUBS 0.043054f
C1217 VDD2.n54 VSUBS 0.019287f
C1218 VDD2.n55 VSUBS 0.018215f
C1219 VDD2.n56 VSUBS 0.033898f
C1220 VDD2.n57 VSUBS 0.033898f
C1221 VDD2.n58 VSUBS 0.018215f
C1222 VDD2.n59 VSUBS 0.019287f
C1223 VDD2.n60 VSUBS 0.043054f
C1224 VDD2.n61 VSUBS 0.043054f
C1225 VDD2.n62 VSUBS 0.019287f
C1226 VDD2.n63 VSUBS 0.018215f
C1227 VDD2.n64 VSUBS 0.033898f
C1228 VDD2.n65 VSUBS 0.033898f
C1229 VDD2.n66 VSUBS 0.018215f
C1230 VDD2.n67 VSUBS 0.019287f
C1231 VDD2.n68 VSUBS 0.043054f
C1232 VDD2.n69 VSUBS 0.108489f
C1233 VDD2.n70 VSUBS 0.019287f
C1234 VDD2.n71 VSUBS 0.03577f
C1235 VDD2.n72 VSUBS 0.087614f
C1236 VDD2.n73 VSUBS 0.107268f
C1237 VDD2.n74 VSUBS 3.95369f
C1238 VDD2.t2 VSUBS 0.195009f
C1239 VDD2.t7 VSUBS 0.195009f
C1240 VDD2.n75 VSUBS 1.38654f
C1241 VDD2.n76 VSUBS 1.023f
C1242 VDD2.t5 VSUBS 0.195009f
C1243 VDD2.t3 VSUBS 0.195009f
C1244 VDD2.n77 VSUBS 1.41935f
C1245 VTAIL.t15 VSUBS 0.189185f
C1246 VTAIL.t17 VSUBS 0.189185f
C1247 VTAIL.n0 VSUBS 1.22185f
C1248 VTAIL.n1 VSUBS 1.1208f
C1249 VTAIL.n2 VSUBS 0.036247f
C1250 VTAIL.n3 VSUBS 0.032885f
C1251 VTAIL.n4 VSUBS 0.017671f
C1252 VTAIL.n5 VSUBS 0.041768f
C1253 VTAIL.n6 VSUBS 0.018711f
C1254 VTAIL.n7 VSUBS 0.032885f
C1255 VTAIL.n8 VSUBS 0.017671f
C1256 VTAIL.n9 VSUBS 0.041768f
C1257 VTAIL.n10 VSUBS 0.018711f
C1258 VTAIL.n11 VSUBS 0.935139f
C1259 VTAIL.n12 VSUBS 0.017671f
C1260 VTAIL.t3 VSUBS 0.089759f
C1261 VTAIL.n13 VSUBS 0.189038f
C1262 VTAIL.n14 VSUBS 0.031418f
C1263 VTAIL.n15 VSUBS 0.031326f
C1264 VTAIL.n16 VSUBS 0.041768f
C1265 VTAIL.n17 VSUBS 0.018711f
C1266 VTAIL.n18 VSUBS 0.017671f
C1267 VTAIL.n19 VSUBS 0.032885f
C1268 VTAIL.n20 VSUBS 0.032885f
C1269 VTAIL.n21 VSUBS 0.017671f
C1270 VTAIL.n22 VSUBS 0.018711f
C1271 VTAIL.n23 VSUBS 0.041768f
C1272 VTAIL.n24 VSUBS 0.041768f
C1273 VTAIL.n25 VSUBS 0.018711f
C1274 VTAIL.n26 VSUBS 0.017671f
C1275 VTAIL.n27 VSUBS 0.032885f
C1276 VTAIL.n28 VSUBS 0.032885f
C1277 VTAIL.n29 VSUBS 0.017671f
C1278 VTAIL.n30 VSUBS 0.018711f
C1279 VTAIL.n31 VSUBS 0.041768f
C1280 VTAIL.n32 VSUBS 0.105249f
C1281 VTAIL.n33 VSUBS 0.018711f
C1282 VTAIL.n34 VSUBS 0.034702f
C1283 VTAIL.n35 VSUBS 0.084997f
C1284 VTAIL.n36 VSUBS 0.08142f
C1285 VTAIL.n37 VSUBS 0.620081f
C1286 VTAIL.t2 VSUBS 0.189185f
C1287 VTAIL.t1 VSUBS 0.189185f
C1288 VTAIL.n38 VSUBS 1.22185f
C1289 VTAIL.n39 VSUBS 1.33342f
C1290 VTAIL.t0 VSUBS 0.189185f
C1291 VTAIL.t5 VSUBS 0.189185f
C1292 VTAIL.n40 VSUBS 1.22185f
C1293 VTAIL.n41 VSUBS 2.80322f
C1294 VTAIL.t18 VSUBS 0.189185f
C1295 VTAIL.t16 VSUBS 0.189185f
C1296 VTAIL.n42 VSUBS 1.22186f
C1297 VTAIL.n43 VSUBS 2.80321f
C1298 VTAIL.t14 VSUBS 0.189185f
C1299 VTAIL.t13 VSUBS 0.189185f
C1300 VTAIL.n44 VSUBS 1.22186f
C1301 VTAIL.n45 VSUBS 1.33341f
C1302 VTAIL.n46 VSUBS 0.036247f
C1303 VTAIL.n47 VSUBS 0.032885f
C1304 VTAIL.n48 VSUBS 0.017671f
C1305 VTAIL.n49 VSUBS 0.041768f
C1306 VTAIL.n50 VSUBS 0.018711f
C1307 VTAIL.n51 VSUBS 0.032885f
C1308 VTAIL.n52 VSUBS 0.017671f
C1309 VTAIL.n53 VSUBS 0.041768f
C1310 VTAIL.n54 VSUBS 0.018711f
C1311 VTAIL.n55 VSUBS 0.935139f
C1312 VTAIL.n56 VSUBS 0.017671f
C1313 VTAIL.t12 VSUBS 0.089759f
C1314 VTAIL.n57 VSUBS 0.189038f
C1315 VTAIL.n58 VSUBS 0.031418f
C1316 VTAIL.n59 VSUBS 0.031326f
C1317 VTAIL.n60 VSUBS 0.041768f
C1318 VTAIL.n61 VSUBS 0.018711f
C1319 VTAIL.n62 VSUBS 0.017671f
C1320 VTAIL.n63 VSUBS 0.032885f
C1321 VTAIL.n64 VSUBS 0.032885f
C1322 VTAIL.n65 VSUBS 0.017671f
C1323 VTAIL.n66 VSUBS 0.018711f
C1324 VTAIL.n67 VSUBS 0.041768f
C1325 VTAIL.n68 VSUBS 0.041768f
C1326 VTAIL.n69 VSUBS 0.018711f
C1327 VTAIL.n70 VSUBS 0.017671f
C1328 VTAIL.n71 VSUBS 0.032885f
C1329 VTAIL.n72 VSUBS 0.032885f
C1330 VTAIL.n73 VSUBS 0.017671f
C1331 VTAIL.n74 VSUBS 0.018711f
C1332 VTAIL.n75 VSUBS 0.041768f
C1333 VTAIL.n76 VSUBS 0.105249f
C1334 VTAIL.n77 VSUBS 0.018711f
C1335 VTAIL.n78 VSUBS 0.034702f
C1336 VTAIL.n79 VSUBS 0.084997f
C1337 VTAIL.n80 VSUBS 0.08142f
C1338 VTAIL.n81 VSUBS 0.620081f
C1339 VTAIL.t7 VSUBS 0.189185f
C1340 VTAIL.t9 VSUBS 0.189185f
C1341 VTAIL.n82 VSUBS 1.22186f
C1342 VTAIL.n83 VSUBS 1.20415f
C1343 VTAIL.t8 VSUBS 0.189185f
C1344 VTAIL.t4 VSUBS 0.189185f
C1345 VTAIL.n84 VSUBS 1.22186f
C1346 VTAIL.n85 VSUBS 1.33341f
C1347 VTAIL.n86 VSUBS 0.036247f
C1348 VTAIL.n87 VSUBS 0.032885f
C1349 VTAIL.n88 VSUBS 0.017671f
C1350 VTAIL.n89 VSUBS 0.041768f
C1351 VTAIL.n90 VSUBS 0.018711f
C1352 VTAIL.n91 VSUBS 0.032885f
C1353 VTAIL.n92 VSUBS 0.017671f
C1354 VTAIL.n93 VSUBS 0.041768f
C1355 VTAIL.n94 VSUBS 0.018711f
C1356 VTAIL.n95 VSUBS 0.935139f
C1357 VTAIL.n96 VSUBS 0.017671f
C1358 VTAIL.t6 VSUBS 0.089759f
C1359 VTAIL.n97 VSUBS 0.189038f
C1360 VTAIL.n98 VSUBS 0.031418f
C1361 VTAIL.n99 VSUBS 0.031326f
C1362 VTAIL.n100 VSUBS 0.041768f
C1363 VTAIL.n101 VSUBS 0.018711f
C1364 VTAIL.n102 VSUBS 0.017671f
C1365 VTAIL.n103 VSUBS 0.032885f
C1366 VTAIL.n104 VSUBS 0.032885f
C1367 VTAIL.n105 VSUBS 0.017671f
C1368 VTAIL.n106 VSUBS 0.018711f
C1369 VTAIL.n107 VSUBS 0.041768f
C1370 VTAIL.n108 VSUBS 0.041768f
C1371 VTAIL.n109 VSUBS 0.018711f
C1372 VTAIL.n110 VSUBS 0.017671f
C1373 VTAIL.n111 VSUBS 0.032885f
C1374 VTAIL.n112 VSUBS 0.032885f
C1375 VTAIL.n113 VSUBS 0.017671f
C1376 VTAIL.n114 VSUBS 0.018711f
C1377 VTAIL.n115 VSUBS 0.041768f
C1378 VTAIL.n116 VSUBS 0.105249f
C1379 VTAIL.n117 VSUBS 0.018711f
C1380 VTAIL.n118 VSUBS 0.034702f
C1381 VTAIL.n119 VSUBS 0.084997f
C1382 VTAIL.n120 VSUBS 0.08142f
C1383 VTAIL.n121 VSUBS 1.86106f
C1384 VTAIL.n122 VSUBS 0.036247f
C1385 VTAIL.n123 VSUBS 0.032885f
C1386 VTAIL.n124 VSUBS 0.017671f
C1387 VTAIL.n125 VSUBS 0.041768f
C1388 VTAIL.n126 VSUBS 0.018711f
C1389 VTAIL.n127 VSUBS 0.032885f
C1390 VTAIL.n128 VSUBS 0.017671f
C1391 VTAIL.n129 VSUBS 0.041768f
C1392 VTAIL.n130 VSUBS 0.018711f
C1393 VTAIL.n131 VSUBS 0.935139f
C1394 VTAIL.n132 VSUBS 0.017671f
C1395 VTAIL.t11 VSUBS 0.089759f
C1396 VTAIL.n133 VSUBS 0.189038f
C1397 VTAIL.n134 VSUBS 0.031418f
C1398 VTAIL.n135 VSUBS 0.031326f
C1399 VTAIL.n136 VSUBS 0.041768f
C1400 VTAIL.n137 VSUBS 0.018711f
C1401 VTAIL.n138 VSUBS 0.017671f
C1402 VTAIL.n139 VSUBS 0.032885f
C1403 VTAIL.n140 VSUBS 0.032885f
C1404 VTAIL.n141 VSUBS 0.017671f
C1405 VTAIL.n142 VSUBS 0.018711f
C1406 VTAIL.n143 VSUBS 0.041768f
C1407 VTAIL.n144 VSUBS 0.041768f
C1408 VTAIL.n145 VSUBS 0.018711f
C1409 VTAIL.n146 VSUBS 0.017671f
C1410 VTAIL.n147 VSUBS 0.032885f
C1411 VTAIL.n148 VSUBS 0.032885f
C1412 VTAIL.n149 VSUBS 0.017671f
C1413 VTAIL.n150 VSUBS 0.018711f
C1414 VTAIL.n151 VSUBS 0.041768f
C1415 VTAIL.n152 VSUBS 0.105249f
C1416 VTAIL.n153 VSUBS 0.018711f
C1417 VTAIL.n154 VSUBS 0.034702f
C1418 VTAIL.n155 VSUBS 0.084997f
C1419 VTAIL.n156 VSUBS 0.08142f
C1420 VTAIL.n157 VSUBS 1.86106f
C1421 VTAIL.t10 VSUBS 0.189185f
C1422 VTAIL.t19 VSUBS 0.189185f
C1423 VTAIL.n158 VSUBS 1.22185f
C1424 VTAIL.n159 VSUBS 1.05869f
C1425 VN.t8 VSUBS 2.00475f
C1426 VN.n0 VSUBS 0.830133f
C1427 VN.n1 VSUBS 0.028685f
C1428 VN.n2 VSUBS 0.050652f
C1429 VN.n3 VSUBS 0.028685f
C1430 VN.n4 VSUBS 0.044265f
C1431 VN.n5 VSUBS 0.028685f
C1432 VN.n6 VSUBS 0.044872f
C1433 VN.n7 VSUBS 0.028685f
C1434 VN.n8 VSUBS 0.040063f
C1435 VN.n9 VSUBS 0.028685f
C1436 VN.n10 VSUBS 0.038523f
C1437 VN.n11 VSUBS 0.028685f
C1438 VN.n12 VSUBS 0.035861f
C1439 VN.t9 VSUBS 2.00475f
C1440 VN.n13 VSUBS 0.821604f
C1441 VN.t5 VSUBS 2.37944f
C1442 VN.n14 VSUBS 0.787346f
C1443 VN.n15 VSUBS 0.359632f
C1444 VN.n16 VSUBS 0.028685f
C1445 VN.n17 VSUBS 0.053193f
C1446 VN.n18 VSUBS 0.053193f
C1447 VN.n19 VSUBS 0.044872f
C1448 VN.n20 VSUBS 0.028685f
C1449 VN.n21 VSUBS 0.028685f
C1450 VN.n22 VSUBS 0.028685f
C1451 VN.n23 VSUBS 0.053193f
C1452 VN.n24 VSUBS 0.053193f
C1453 VN.t0 VSUBS 2.00475f
C1454 VN.n25 VSUBS 0.726577f
C1455 VN.n26 VSUBS 0.040063f
C1456 VN.n27 VSUBS 0.028685f
C1457 VN.n28 VSUBS 0.028685f
C1458 VN.n29 VSUBS 0.028685f
C1459 VN.n30 VSUBS 0.053193f
C1460 VN.n31 VSUBS 0.053193f
C1461 VN.n32 VSUBS 0.038523f
C1462 VN.n33 VSUBS 0.028685f
C1463 VN.n34 VSUBS 0.028685f
C1464 VN.n35 VSUBS 0.028685f
C1465 VN.n36 VSUBS 0.053193f
C1466 VN.n37 VSUBS 0.053193f
C1467 VN.t3 VSUBS 2.00475f
C1468 VN.n38 VSUBS 0.726577f
C1469 VN.n39 VSUBS 0.035861f
C1470 VN.n40 VSUBS 0.028685f
C1471 VN.n41 VSUBS 0.028685f
C1472 VN.n42 VSUBS 0.028685f
C1473 VN.n43 VSUBS 0.053193f
C1474 VN.n44 VSUBS 0.05593f
C1475 VN.n45 VSUBS 0.030006f
C1476 VN.n46 VSUBS 0.028685f
C1477 VN.n47 VSUBS 0.028685f
C1478 VN.n48 VSUBS 0.028685f
C1479 VN.n49 VSUBS 0.053193f
C1480 VN.n50 VSUBS 0.053193f
C1481 VN.n51 VSUBS 0.03166f
C1482 VN.n52 VSUBS 0.046289f
C1483 VN.n53 VSUBS 0.083422f
C1484 VN.t1 VSUBS 2.00475f
C1485 VN.n54 VSUBS 0.830133f
C1486 VN.n55 VSUBS 0.028685f
C1487 VN.n56 VSUBS 0.050652f
C1488 VN.n57 VSUBS 0.028685f
C1489 VN.n58 VSUBS 0.044265f
C1490 VN.n59 VSUBS 0.028685f
C1491 VN.t7 VSUBS 2.00475f
C1492 VN.n60 VSUBS 0.726577f
C1493 VN.n61 VSUBS 0.044872f
C1494 VN.n62 VSUBS 0.028685f
C1495 VN.n63 VSUBS 0.040063f
C1496 VN.n64 VSUBS 0.028685f
C1497 VN.t2 VSUBS 2.00475f
C1498 VN.n65 VSUBS 0.726577f
C1499 VN.n66 VSUBS 0.038523f
C1500 VN.n67 VSUBS 0.028685f
C1501 VN.n68 VSUBS 0.035861f
C1502 VN.t6 VSUBS 2.37944f
C1503 VN.t4 VSUBS 2.00475f
C1504 VN.n69 VSUBS 0.821604f
C1505 VN.n70 VSUBS 0.787346f
C1506 VN.n71 VSUBS 0.359632f
C1507 VN.n72 VSUBS 0.028685f
C1508 VN.n73 VSUBS 0.053193f
C1509 VN.n74 VSUBS 0.053193f
C1510 VN.n75 VSUBS 0.044872f
C1511 VN.n76 VSUBS 0.028685f
C1512 VN.n77 VSUBS 0.028685f
C1513 VN.n78 VSUBS 0.028685f
C1514 VN.n79 VSUBS 0.053193f
C1515 VN.n80 VSUBS 0.053193f
C1516 VN.n81 VSUBS 0.040063f
C1517 VN.n82 VSUBS 0.028685f
C1518 VN.n83 VSUBS 0.028685f
C1519 VN.n84 VSUBS 0.028685f
C1520 VN.n85 VSUBS 0.053193f
C1521 VN.n86 VSUBS 0.053193f
C1522 VN.n87 VSUBS 0.038523f
C1523 VN.n88 VSUBS 0.028685f
C1524 VN.n89 VSUBS 0.028685f
C1525 VN.n90 VSUBS 0.028685f
C1526 VN.n91 VSUBS 0.053193f
C1527 VN.n92 VSUBS 0.053193f
C1528 VN.n93 VSUBS 0.035861f
C1529 VN.n94 VSUBS 0.028685f
C1530 VN.n95 VSUBS 0.028685f
C1531 VN.n96 VSUBS 0.028685f
C1532 VN.n97 VSUBS 0.053193f
C1533 VN.n98 VSUBS 0.05593f
C1534 VN.n99 VSUBS 0.030006f
C1535 VN.n100 VSUBS 0.028685f
C1536 VN.n101 VSUBS 0.028685f
C1537 VN.n102 VSUBS 0.028685f
C1538 VN.n103 VSUBS 0.053193f
C1539 VN.n104 VSUBS 0.053193f
C1540 VN.n105 VSUBS 0.03166f
C1541 VN.n106 VSUBS 0.046289f
C1542 VN.n107 VSUBS 1.88784f
.ends

