* NGSPICE file created from diff_pair_sample_0219.ext - technology: sky130A

.subckt diff_pair_sample_0219 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n2326_n1360# sky130_fd_pr__pfet_01v8 ad=0.7644 pd=4.7 as=0 ps=0 w=1.96 l=1.93
X1 B.t8 B.t6 B.t7 w_n2326_n1360# sky130_fd_pr__pfet_01v8 ad=0.7644 pd=4.7 as=0 ps=0 w=1.96 l=1.93
X2 B.t5 B.t3 B.t4 w_n2326_n1360# sky130_fd_pr__pfet_01v8 ad=0.7644 pd=4.7 as=0 ps=0 w=1.96 l=1.93
X3 VTAIL.t7 VN.t0 VDD2.t3 w_n2326_n1360# sky130_fd_pr__pfet_01v8 ad=0.7644 pd=4.7 as=0.3234 ps=2.29 w=1.96 l=1.93
X4 VDD2.t2 VN.t1 VTAIL.t6 w_n2326_n1360# sky130_fd_pr__pfet_01v8 ad=0.3234 pd=2.29 as=0.7644 ps=4.7 w=1.96 l=1.93
X5 VDD1.t3 VP.t0 VTAIL.t3 w_n2326_n1360# sky130_fd_pr__pfet_01v8 ad=0.3234 pd=2.29 as=0.7644 ps=4.7 w=1.96 l=1.93
X6 VTAIL.t0 VP.t1 VDD1.t2 w_n2326_n1360# sky130_fd_pr__pfet_01v8 ad=0.7644 pd=4.7 as=0.3234 ps=2.29 w=1.96 l=1.93
X7 VDD1.t1 VP.t2 VTAIL.t1 w_n2326_n1360# sky130_fd_pr__pfet_01v8 ad=0.3234 pd=2.29 as=0.7644 ps=4.7 w=1.96 l=1.93
X8 VTAIL.t2 VP.t3 VDD1.t0 w_n2326_n1360# sky130_fd_pr__pfet_01v8 ad=0.7644 pd=4.7 as=0.3234 ps=2.29 w=1.96 l=1.93
X9 B.t2 B.t0 B.t1 w_n2326_n1360# sky130_fd_pr__pfet_01v8 ad=0.7644 pd=4.7 as=0 ps=0 w=1.96 l=1.93
X10 VTAIL.t5 VN.t2 VDD2.t0 w_n2326_n1360# sky130_fd_pr__pfet_01v8 ad=0.7644 pd=4.7 as=0.3234 ps=2.29 w=1.96 l=1.93
X11 VDD2.t1 VN.t3 VTAIL.t4 w_n2326_n1360# sky130_fd_pr__pfet_01v8 ad=0.3234 pd=2.29 as=0.7644 ps=4.7 w=1.96 l=1.93
R0 B.n280 B.n37 585
R1 B.n282 B.n281 585
R2 B.n283 B.n36 585
R3 B.n285 B.n284 585
R4 B.n286 B.n35 585
R5 B.n288 B.n287 585
R6 B.n289 B.n34 585
R7 B.n291 B.n290 585
R8 B.n292 B.n33 585
R9 B.n294 B.n293 585
R10 B.n295 B.n32 585
R11 B.n297 B.n296 585
R12 B.n299 B.n29 585
R13 B.n301 B.n300 585
R14 B.n302 B.n28 585
R15 B.n304 B.n303 585
R16 B.n305 B.n27 585
R17 B.n307 B.n306 585
R18 B.n308 B.n26 585
R19 B.n310 B.n309 585
R20 B.n311 B.n25 585
R21 B.n313 B.n312 585
R22 B.n315 B.n314 585
R23 B.n316 B.n21 585
R24 B.n318 B.n317 585
R25 B.n319 B.n20 585
R26 B.n321 B.n320 585
R27 B.n322 B.n19 585
R28 B.n324 B.n323 585
R29 B.n325 B.n18 585
R30 B.n327 B.n326 585
R31 B.n328 B.n17 585
R32 B.n330 B.n329 585
R33 B.n331 B.n16 585
R34 B.n279 B.n278 585
R35 B.n277 B.n38 585
R36 B.n276 B.n275 585
R37 B.n274 B.n39 585
R38 B.n273 B.n272 585
R39 B.n271 B.n40 585
R40 B.n270 B.n269 585
R41 B.n268 B.n41 585
R42 B.n267 B.n266 585
R43 B.n265 B.n42 585
R44 B.n264 B.n263 585
R45 B.n262 B.n43 585
R46 B.n261 B.n260 585
R47 B.n259 B.n44 585
R48 B.n258 B.n257 585
R49 B.n256 B.n45 585
R50 B.n255 B.n254 585
R51 B.n253 B.n46 585
R52 B.n252 B.n251 585
R53 B.n250 B.n47 585
R54 B.n249 B.n248 585
R55 B.n247 B.n48 585
R56 B.n246 B.n245 585
R57 B.n244 B.n49 585
R58 B.n243 B.n242 585
R59 B.n241 B.n50 585
R60 B.n240 B.n239 585
R61 B.n238 B.n51 585
R62 B.n237 B.n236 585
R63 B.n235 B.n52 585
R64 B.n234 B.n233 585
R65 B.n232 B.n53 585
R66 B.n231 B.n230 585
R67 B.n229 B.n54 585
R68 B.n228 B.n227 585
R69 B.n226 B.n55 585
R70 B.n225 B.n224 585
R71 B.n223 B.n56 585
R72 B.n222 B.n221 585
R73 B.n220 B.n57 585
R74 B.n219 B.n218 585
R75 B.n217 B.n58 585
R76 B.n216 B.n215 585
R77 B.n214 B.n59 585
R78 B.n213 B.n212 585
R79 B.n211 B.n60 585
R80 B.n210 B.n209 585
R81 B.n208 B.n61 585
R82 B.n207 B.n206 585
R83 B.n205 B.n62 585
R84 B.n204 B.n203 585
R85 B.n202 B.n63 585
R86 B.n201 B.n200 585
R87 B.n199 B.n64 585
R88 B.n198 B.n197 585
R89 B.n196 B.n65 585
R90 B.n195 B.n194 585
R91 B.n142 B.n87 585
R92 B.n144 B.n143 585
R93 B.n145 B.n86 585
R94 B.n147 B.n146 585
R95 B.n148 B.n85 585
R96 B.n150 B.n149 585
R97 B.n151 B.n84 585
R98 B.n153 B.n152 585
R99 B.n154 B.n83 585
R100 B.n156 B.n155 585
R101 B.n157 B.n82 585
R102 B.n159 B.n158 585
R103 B.n161 B.n79 585
R104 B.n163 B.n162 585
R105 B.n164 B.n78 585
R106 B.n166 B.n165 585
R107 B.n167 B.n77 585
R108 B.n169 B.n168 585
R109 B.n170 B.n76 585
R110 B.n172 B.n171 585
R111 B.n173 B.n75 585
R112 B.n175 B.n174 585
R113 B.n177 B.n176 585
R114 B.n178 B.n71 585
R115 B.n180 B.n179 585
R116 B.n181 B.n70 585
R117 B.n183 B.n182 585
R118 B.n184 B.n69 585
R119 B.n186 B.n185 585
R120 B.n187 B.n68 585
R121 B.n189 B.n188 585
R122 B.n190 B.n67 585
R123 B.n192 B.n191 585
R124 B.n193 B.n66 585
R125 B.n141 B.n140 585
R126 B.n139 B.n88 585
R127 B.n138 B.n137 585
R128 B.n136 B.n89 585
R129 B.n135 B.n134 585
R130 B.n133 B.n90 585
R131 B.n132 B.n131 585
R132 B.n130 B.n91 585
R133 B.n129 B.n128 585
R134 B.n127 B.n92 585
R135 B.n126 B.n125 585
R136 B.n124 B.n93 585
R137 B.n123 B.n122 585
R138 B.n121 B.n94 585
R139 B.n120 B.n119 585
R140 B.n118 B.n95 585
R141 B.n117 B.n116 585
R142 B.n115 B.n96 585
R143 B.n114 B.n113 585
R144 B.n112 B.n97 585
R145 B.n111 B.n110 585
R146 B.n109 B.n98 585
R147 B.n108 B.n107 585
R148 B.n106 B.n99 585
R149 B.n105 B.n104 585
R150 B.n103 B.n100 585
R151 B.n102 B.n101 585
R152 B.n2 B.n0 585
R153 B.n373 B.n1 585
R154 B.n372 B.n371 585
R155 B.n370 B.n3 585
R156 B.n369 B.n368 585
R157 B.n367 B.n4 585
R158 B.n366 B.n365 585
R159 B.n364 B.n5 585
R160 B.n363 B.n362 585
R161 B.n361 B.n6 585
R162 B.n360 B.n359 585
R163 B.n358 B.n7 585
R164 B.n357 B.n356 585
R165 B.n355 B.n8 585
R166 B.n354 B.n353 585
R167 B.n352 B.n9 585
R168 B.n351 B.n350 585
R169 B.n349 B.n10 585
R170 B.n348 B.n347 585
R171 B.n346 B.n11 585
R172 B.n345 B.n344 585
R173 B.n343 B.n12 585
R174 B.n342 B.n341 585
R175 B.n340 B.n13 585
R176 B.n339 B.n338 585
R177 B.n337 B.n14 585
R178 B.n336 B.n335 585
R179 B.n334 B.n15 585
R180 B.n333 B.n332 585
R181 B.n375 B.n374 585
R182 B.n140 B.n87 487.695
R183 B.n332 B.n331 487.695
R184 B.n194 B.n193 487.695
R185 B.n278 B.n37 487.695
R186 B.n72 B.t2 291.392
R187 B.n30 B.t4 291.392
R188 B.n80 B.t11 291.392
R189 B.n22 B.t7 291.392
R190 B.n73 B.t1 247.561
R191 B.n31 B.t5 247.561
R192 B.n81 B.t10 247.561
R193 B.n23 B.t8 247.561
R194 B.n72 B.t0 231.224
R195 B.n80 B.t9 231.224
R196 B.n22 B.t6 231.224
R197 B.n30 B.t3 231.224
R198 B.n140 B.n139 163.367
R199 B.n139 B.n138 163.367
R200 B.n138 B.n89 163.367
R201 B.n134 B.n89 163.367
R202 B.n134 B.n133 163.367
R203 B.n133 B.n132 163.367
R204 B.n132 B.n91 163.367
R205 B.n128 B.n91 163.367
R206 B.n128 B.n127 163.367
R207 B.n127 B.n126 163.367
R208 B.n126 B.n93 163.367
R209 B.n122 B.n93 163.367
R210 B.n122 B.n121 163.367
R211 B.n121 B.n120 163.367
R212 B.n120 B.n95 163.367
R213 B.n116 B.n95 163.367
R214 B.n116 B.n115 163.367
R215 B.n115 B.n114 163.367
R216 B.n114 B.n97 163.367
R217 B.n110 B.n97 163.367
R218 B.n110 B.n109 163.367
R219 B.n109 B.n108 163.367
R220 B.n108 B.n99 163.367
R221 B.n104 B.n99 163.367
R222 B.n104 B.n103 163.367
R223 B.n103 B.n102 163.367
R224 B.n102 B.n2 163.367
R225 B.n374 B.n2 163.367
R226 B.n374 B.n373 163.367
R227 B.n373 B.n372 163.367
R228 B.n372 B.n3 163.367
R229 B.n368 B.n3 163.367
R230 B.n368 B.n367 163.367
R231 B.n367 B.n366 163.367
R232 B.n366 B.n5 163.367
R233 B.n362 B.n5 163.367
R234 B.n362 B.n361 163.367
R235 B.n361 B.n360 163.367
R236 B.n360 B.n7 163.367
R237 B.n356 B.n7 163.367
R238 B.n356 B.n355 163.367
R239 B.n355 B.n354 163.367
R240 B.n354 B.n9 163.367
R241 B.n350 B.n9 163.367
R242 B.n350 B.n349 163.367
R243 B.n349 B.n348 163.367
R244 B.n348 B.n11 163.367
R245 B.n344 B.n11 163.367
R246 B.n344 B.n343 163.367
R247 B.n343 B.n342 163.367
R248 B.n342 B.n13 163.367
R249 B.n338 B.n13 163.367
R250 B.n338 B.n337 163.367
R251 B.n337 B.n336 163.367
R252 B.n336 B.n15 163.367
R253 B.n332 B.n15 163.367
R254 B.n144 B.n87 163.367
R255 B.n145 B.n144 163.367
R256 B.n146 B.n145 163.367
R257 B.n146 B.n85 163.367
R258 B.n150 B.n85 163.367
R259 B.n151 B.n150 163.367
R260 B.n152 B.n151 163.367
R261 B.n152 B.n83 163.367
R262 B.n156 B.n83 163.367
R263 B.n157 B.n156 163.367
R264 B.n158 B.n157 163.367
R265 B.n158 B.n79 163.367
R266 B.n163 B.n79 163.367
R267 B.n164 B.n163 163.367
R268 B.n165 B.n164 163.367
R269 B.n165 B.n77 163.367
R270 B.n169 B.n77 163.367
R271 B.n170 B.n169 163.367
R272 B.n171 B.n170 163.367
R273 B.n171 B.n75 163.367
R274 B.n175 B.n75 163.367
R275 B.n176 B.n175 163.367
R276 B.n176 B.n71 163.367
R277 B.n180 B.n71 163.367
R278 B.n181 B.n180 163.367
R279 B.n182 B.n181 163.367
R280 B.n182 B.n69 163.367
R281 B.n186 B.n69 163.367
R282 B.n187 B.n186 163.367
R283 B.n188 B.n187 163.367
R284 B.n188 B.n67 163.367
R285 B.n192 B.n67 163.367
R286 B.n193 B.n192 163.367
R287 B.n194 B.n65 163.367
R288 B.n198 B.n65 163.367
R289 B.n199 B.n198 163.367
R290 B.n200 B.n199 163.367
R291 B.n200 B.n63 163.367
R292 B.n204 B.n63 163.367
R293 B.n205 B.n204 163.367
R294 B.n206 B.n205 163.367
R295 B.n206 B.n61 163.367
R296 B.n210 B.n61 163.367
R297 B.n211 B.n210 163.367
R298 B.n212 B.n211 163.367
R299 B.n212 B.n59 163.367
R300 B.n216 B.n59 163.367
R301 B.n217 B.n216 163.367
R302 B.n218 B.n217 163.367
R303 B.n218 B.n57 163.367
R304 B.n222 B.n57 163.367
R305 B.n223 B.n222 163.367
R306 B.n224 B.n223 163.367
R307 B.n224 B.n55 163.367
R308 B.n228 B.n55 163.367
R309 B.n229 B.n228 163.367
R310 B.n230 B.n229 163.367
R311 B.n230 B.n53 163.367
R312 B.n234 B.n53 163.367
R313 B.n235 B.n234 163.367
R314 B.n236 B.n235 163.367
R315 B.n236 B.n51 163.367
R316 B.n240 B.n51 163.367
R317 B.n241 B.n240 163.367
R318 B.n242 B.n241 163.367
R319 B.n242 B.n49 163.367
R320 B.n246 B.n49 163.367
R321 B.n247 B.n246 163.367
R322 B.n248 B.n247 163.367
R323 B.n248 B.n47 163.367
R324 B.n252 B.n47 163.367
R325 B.n253 B.n252 163.367
R326 B.n254 B.n253 163.367
R327 B.n254 B.n45 163.367
R328 B.n258 B.n45 163.367
R329 B.n259 B.n258 163.367
R330 B.n260 B.n259 163.367
R331 B.n260 B.n43 163.367
R332 B.n264 B.n43 163.367
R333 B.n265 B.n264 163.367
R334 B.n266 B.n265 163.367
R335 B.n266 B.n41 163.367
R336 B.n270 B.n41 163.367
R337 B.n271 B.n270 163.367
R338 B.n272 B.n271 163.367
R339 B.n272 B.n39 163.367
R340 B.n276 B.n39 163.367
R341 B.n277 B.n276 163.367
R342 B.n278 B.n277 163.367
R343 B.n331 B.n330 163.367
R344 B.n330 B.n17 163.367
R345 B.n326 B.n17 163.367
R346 B.n326 B.n325 163.367
R347 B.n325 B.n324 163.367
R348 B.n324 B.n19 163.367
R349 B.n320 B.n19 163.367
R350 B.n320 B.n319 163.367
R351 B.n319 B.n318 163.367
R352 B.n318 B.n21 163.367
R353 B.n314 B.n21 163.367
R354 B.n314 B.n313 163.367
R355 B.n313 B.n25 163.367
R356 B.n309 B.n25 163.367
R357 B.n309 B.n308 163.367
R358 B.n308 B.n307 163.367
R359 B.n307 B.n27 163.367
R360 B.n303 B.n27 163.367
R361 B.n303 B.n302 163.367
R362 B.n302 B.n301 163.367
R363 B.n301 B.n29 163.367
R364 B.n296 B.n29 163.367
R365 B.n296 B.n295 163.367
R366 B.n295 B.n294 163.367
R367 B.n294 B.n33 163.367
R368 B.n290 B.n33 163.367
R369 B.n290 B.n289 163.367
R370 B.n289 B.n288 163.367
R371 B.n288 B.n35 163.367
R372 B.n284 B.n35 163.367
R373 B.n284 B.n283 163.367
R374 B.n283 B.n282 163.367
R375 B.n282 B.n37 163.367
R376 B.n74 B.n73 59.5399
R377 B.n160 B.n81 59.5399
R378 B.n24 B.n23 59.5399
R379 B.n298 B.n31 59.5399
R380 B.n73 B.n72 43.8308
R381 B.n81 B.n80 43.8308
R382 B.n23 B.n22 43.8308
R383 B.n31 B.n30 43.8308
R384 B.n333 B.n16 31.6883
R385 B.n280 B.n279 31.6883
R386 B.n195 B.n66 31.6883
R387 B.n142 B.n141 31.6883
R388 B B.n375 18.0485
R389 B.n329 B.n16 10.6151
R390 B.n329 B.n328 10.6151
R391 B.n328 B.n327 10.6151
R392 B.n327 B.n18 10.6151
R393 B.n323 B.n18 10.6151
R394 B.n323 B.n322 10.6151
R395 B.n322 B.n321 10.6151
R396 B.n321 B.n20 10.6151
R397 B.n317 B.n20 10.6151
R398 B.n317 B.n316 10.6151
R399 B.n316 B.n315 10.6151
R400 B.n312 B.n311 10.6151
R401 B.n311 B.n310 10.6151
R402 B.n310 B.n26 10.6151
R403 B.n306 B.n26 10.6151
R404 B.n306 B.n305 10.6151
R405 B.n305 B.n304 10.6151
R406 B.n304 B.n28 10.6151
R407 B.n300 B.n28 10.6151
R408 B.n300 B.n299 10.6151
R409 B.n297 B.n32 10.6151
R410 B.n293 B.n32 10.6151
R411 B.n293 B.n292 10.6151
R412 B.n292 B.n291 10.6151
R413 B.n291 B.n34 10.6151
R414 B.n287 B.n34 10.6151
R415 B.n287 B.n286 10.6151
R416 B.n286 B.n285 10.6151
R417 B.n285 B.n36 10.6151
R418 B.n281 B.n36 10.6151
R419 B.n281 B.n280 10.6151
R420 B.n196 B.n195 10.6151
R421 B.n197 B.n196 10.6151
R422 B.n197 B.n64 10.6151
R423 B.n201 B.n64 10.6151
R424 B.n202 B.n201 10.6151
R425 B.n203 B.n202 10.6151
R426 B.n203 B.n62 10.6151
R427 B.n207 B.n62 10.6151
R428 B.n208 B.n207 10.6151
R429 B.n209 B.n208 10.6151
R430 B.n209 B.n60 10.6151
R431 B.n213 B.n60 10.6151
R432 B.n214 B.n213 10.6151
R433 B.n215 B.n214 10.6151
R434 B.n215 B.n58 10.6151
R435 B.n219 B.n58 10.6151
R436 B.n220 B.n219 10.6151
R437 B.n221 B.n220 10.6151
R438 B.n221 B.n56 10.6151
R439 B.n225 B.n56 10.6151
R440 B.n226 B.n225 10.6151
R441 B.n227 B.n226 10.6151
R442 B.n227 B.n54 10.6151
R443 B.n231 B.n54 10.6151
R444 B.n232 B.n231 10.6151
R445 B.n233 B.n232 10.6151
R446 B.n233 B.n52 10.6151
R447 B.n237 B.n52 10.6151
R448 B.n238 B.n237 10.6151
R449 B.n239 B.n238 10.6151
R450 B.n239 B.n50 10.6151
R451 B.n243 B.n50 10.6151
R452 B.n244 B.n243 10.6151
R453 B.n245 B.n244 10.6151
R454 B.n245 B.n48 10.6151
R455 B.n249 B.n48 10.6151
R456 B.n250 B.n249 10.6151
R457 B.n251 B.n250 10.6151
R458 B.n251 B.n46 10.6151
R459 B.n255 B.n46 10.6151
R460 B.n256 B.n255 10.6151
R461 B.n257 B.n256 10.6151
R462 B.n257 B.n44 10.6151
R463 B.n261 B.n44 10.6151
R464 B.n262 B.n261 10.6151
R465 B.n263 B.n262 10.6151
R466 B.n263 B.n42 10.6151
R467 B.n267 B.n42 10.6151
R468 B.n268 B.n267 10.6151
R469 B.n269 B.n268 10.6151
R470 B.n269 B.n40 10.6151
R471 B.n273 B.n40 10.6151
R472 B.n274 B.n273 10.6151
R473 B.n275 B.n274 10.6151
R474 B.n275 B.n38 10.6151
R475 B.n279 B.n38 10.6151
R476 B.n143 B.n142 10.6151
R477 B.n143 B.n86 10.6151
R478 B.n147 B.n86 10.6151
R479 B.n148 B.n147 10.6151
R480 B.n149 B.n148 10.6151
R481 B.n149 B.n84 10.6151
R482 B.n153 B.n84 10.6151
R483 B.n154 B.n153 10.6151
R484 B.n155 B.n154 10.6151
R485 B.n155 B.n82 10.6151
R486 B.n159 B.n82 10.6151
R487 B.n162 B.n161 10.6151
R488 B.n162 B.n78 10.6151
R489 B.n166 B.n78 10.6151
R490 B.n167 B.n166 10.6151
R491 B.n168 B.n167 10.6151
R492 B.n168 B.n76 10.6151
R493 B.n172 B.n76 10.6151
R494 B.n173 B.n172 10.6151
R495 B.n174 B.n173 10.6151
R496 B.n178 B.n177 10.6151
R497 B.n179 B.n178 10.6151
R498 B.n179 B.n70 10.6151
R499 B.n183 B.n70 10.6151
R500 B.n184 B.n183 10.6151
R501 B.n185 B.n184 10.6151
R502 B.n185 B.n68 10.6151
R503 B.n189 B.n68 10.6151
R504 B.n190 B.n189 10.6151
R505 B.n191 B.n190 10.6151
R506 B.n191 B.n66 10.6151
R507 B.n141 B.n88 10.6151
R508 B.n137 B.n88 10.6151
R509 B.n137 B.n136 10.6151
R510 B.n136 B.n135 10.6151
R511 B.n135 B.n90 10.6151
R512 B.n131 B.n90 10.6151
R513 B.n131 B.n130 10.6151
R514 B.n130 B.n129 10.6151
R515 B.n129 B.n92 10.6151
R516 B.n125 B.n92 10.6151
R517 B.n125 B.n124 10.6151
R518 B.n124 B.n123 10.6151
R519 B.n123 B.n94 10.6151
R520 B.n119 B.n94 10.6151
R521 B.n119 B.n118 10.6151
R522 B.n118 B.n117 10.6151
R523 B.n117 B.n96 10.6151
R524 B.n113 B.n96 10.6151
R525 B.n113 B.n112 10.6151
R526 B.n112 B.n111 10.6151
R527 B.n111 B.n98 10.6151
R528 B.n107 B.n98 10.6151
R529 B.n107 B.n106 10.6151
R530 B.n106 B.n105 10.6151
R531 B.n105 B.n100 10.6151
R532 B.n101 B.n100 10.6151
R533 B.n101 B.n0 10.6151
R534 B.n371 B.n1 10.6151
R535 B.n371 B.n370 10.6151
R536 B.n370 B.n369 10.6151
R537 B.n369 B.n4 10.6151
R538 B.n365 B.n4 10.6151
R539 B.n365 B.n364 10.6151
R540 B.n364 B.n363 10.6151
R541 B.n363 B.n6 10.6151
R542 B.n359 B.n6 10.6151
R543 B.n359 B.n358 10.6151
R544 B.n358 B.n357 10.6151
R545 B.n357 B.n8 10.6151
R546 B.n353 B.n8 10.6151
R547 B.n353 B.n352 10.6151
R548 B.n352 B.n351 10.6151
R549 B.n351 B.n10 10.6151
R550 B.n347 B.n10 10.6151
R551 B.n347 B.n346 10.6151
R552 B.n346 B.n345 10.6151
R553 B.n345 B.n12 10.6151
R554 B.n341 B.n12 10.6151
R555 B.n341 B.n340 10.6151
R556 B.n340 B.n339 10.6151
R557 B.n339 B.n14 10.6151
R558 B.n335 B.n14 10.6151
R559 B.n335 B.n334 10.6151
R560 B.n334 B.n333 10.6151
R561 B.n315 B.n24 9.36635
R562 B.n298 B.n297 9.36635
R563 B.n160 B.n159 9.36635
R564 B.n177 B.n74 9.36635
R565 B.n375 B.n0 2.81026
R566 B.n375 B.n1 2.81026
R567 B.n312 B.n24 1.24928
R568 B.n299 B.n298 1.24928
R569 B.n161 B.n160 1.24928
R570 B.n174 B.n74 1.24928
R571 VN.n0 VN.t2 59.7307
R572 VN.n1 VN.t1 59.7307
R573 VN.n0 VN.t3 59.2093
R574 VN.n1 VN.t0 59.2093
R575 VN VN.n1 44.3718
R576 VN VN.n0 7.52714
R577 VDD2.n2 VDD2.n0 231.304
R578 VDD2.n2 VDD2.n1 200.055
R579 VDD2.n1 VDD2.t3 16.5847
R580 VDD2.n1 VDD2.t2 16.5847
R581 VDD2.n0 VDD2.t0 16.5847
R582 VDD2.n0 VDD2.t1 16.5847
R583 VDD2 VDD2.n2 0.0586897
R584 VTAIL.n58 VTAIL.n56 756.745
R585 VTAIL.n2 VTAIL.n0 756.745
R586 VTAIL.n10 VTAIL.n8 756.745
R587 VTAIL.n18 VTAIL.n16 756.745
R588 VTAIL.n50 VTAIL.n48 756.745
R589 VTAIL.n42 VTAIL.n40 756.745
R590 VTAIL.n34 VTAIL.n32 756.745
R591 VTAIL.n26 VTAIL.n24 756.745
R592 VTAIL.n59 VTAIL.n58 585
R593 VTAIL.n3 VTAIL.n2 585
R594 VTAIL.n11 VTAIL.n10 585
R595 VTAIL.n19 VTAIL.n18 585
R596 VTAIL.n51 VTAIL.n50 585
R597 VTAIL.n43 VTAIL.n42 585
R598 VTAIL.n35 VTAIL.n34 585
R599 VTAIL.n27 VTAIL.n26 585
R600 VTAIL.t4 VTAIL.n57 417.779
R601 VTAIL.t5 VTAIL.n1 417.779
R602 VTAIL.t1 VTAIL.n9 417.779
R603 VTAIL.t2 VTAIL.n17 417.779
R604 VTAIL.t3 VTAIL.n49 417.779
R605 VTAIL.t0 VTAIL.n41 417.779
R606 VTAIL.t6 VTAIL.n33 417.779
R607 VTAIL.t7 VTAIL.n25 417.779
R608 VTAIL.n58 VTAIL.t4 85.8723
R609 VTAIL.n2 VTAIL.t5 85.8723
R610 VTAIL.n10 VTAIL.t1 85.8723
R611 VTAIL.n18 VTAIL.t2 85.8723
R612 VTAIL.n50 VTAIL.t3 85.8723
R613 VTAIL.n42 VTAIL.t0 85.8723
R614 VTAIL.n34 VTAIL.t6 85.8723
R615 VTAIL.n26 VTAIL.t7 85.8723
R616 VTAIL.n63 VTAIL.n62 30.6338
R617 VTAIL.n7 VTAIL.n6 30.6338
R618 VTAIL.n15 VTAIL.n14 30.6338
R619 VTAIL.n23 VTAIL.n22 30.6338
R620 VTAIL.n55 VTAIL.n54 30.6338
R621 VTAIL.n47 VTAIL.n46 30.6338
R622 VTAIL.n39 VTAIL.n38 30.6338
R623 VTAIL.n31 VTAIL.n30 30.6338
R624 VTAIL.n63 VTAIL.n55 16.0048
R625 VTAIL.n31 VTAIL.n23 16.0048
R626 VTAIL.n59 VTAIL.n57 9.84608
R627 VTAIL.n3 VTAIL.n1 9.84608
R628 VTAIL.n11 VTAIL.n9 9.84608
R629 VTAIL.n19 VTAIL.n17 9.84608
R630 VTAIL.n51 VTAIL.n49 9.84608
R631 VTAIL.n43 VTAIL.n41 9.84608
R632 VTAIL.n35 VTAIL.n33 9.84608
R633 VTAIL.n27 VTAIL.n25 9.84608
R634 VTAIL.n62 VTAIL.n61 9.45567
R635 VTAIL.n6 VTAIL.n5 9.45567
R636 VTAIL.n14 VTAIL.n13 9.45567
R637 VTAIL.n22 VTAIL.n21 9.45567
R638 VTAIL.n54 VTAIL.n53 9.45567
R639 VTAIL.n46 VTAIL.n45 9.45567
R640 VTAIL.n38 VTAIL.n37 9.45567
R641 VTAIL.n30 VTAIL.n29 9.45567
R642 VTAIL.n61 VTAIL.n60 9.3005
R643 VTAIL.n5 VTAIL.n4 9.3005
R644 VTAIL.n13 VTAIL.n12 9.3005
R645 VTAIL.n21 VTAIL.n20 9.3005
R646 VTAIL.n53 VTAIL.n52 9.3005
R647 VTAIL.n45 VTAIL.n44 9.3005
R648 VTAIL.n37 VTAIL.n36 9.3005
R649 VTAIL.n29 VTAIL.n28 9.3005
R650 VTAIL.n62 VTAIL.n56 8.14595
R651 VTAIL.n6 VTAIL.n0 8.14595
R652 VTAIL.n14 VTAIL.n8 8.14595
R653 VTAIL.n22 VTAIL.n16 8.14595
R654 VTAIL.n54 VTAIL.n48 8.14595
R655 VTAIL.n46 VTAIL.n40 8.14595
R656 VTAIL.n38 VTAIL.n32 8.14595
R657 VTAIL.n30 VTAIL.n24 8.14595
R658 VTAIL.n60 VTAIL.n59 7.3702
R659 VTAIL.n4 VTAIL.n3 7.3702
R660 VTAIL.n12 VTAIL.n11 7.3702
R661 VTAIL.n20 VTAIL.n19 7.3702
R662 VTAIL.n52 VTAIL.n51 7.3702
R663 VTAIL.n44 VTAIL.n43 7.3702
R664 VTAIL.n36 VTAIL.n35 7.3702
R665 VTAIL.n28 VTAIL.n27 7.3702
R666 VTAIL.n60 VTAIL.n56 5.81868
R667 VTAIL.n4 VTAIL.n0 5.81868
R668 VTAIL.n12 VTAIL.n8 5.81868
R669 VTAIL.n20 VTAIL.n16 5.81868
R670 VTAIL.n52 VTAIL.n48 5.81868
R671 VTAIL.n44 VTAIL.n40 5.81868
R672 VTAIL.n36 VTAIL.n32 5.81868
R673 VTAIL.n28 VTAIL.n24 5.81868
R674 VTAIL.n45 VTAIL.n41 3.32369
R675 VTAIL.n37 VTAIL.n33 3.32369
R676 VTAIL.n29 VTAIL.n25 3.32369
R677 VTAIL.n61 VTAIL.n57 3.32369
R678 VTAIL.n5 VTAIL.n1 3.32369
R679 VTAIL.n13 VTAIL.n9 3.32369
R680 VTAIL.n21 VTAIL.n17 3.32369
R681 VTAIL.n53 VTAIL.n49 3.32369
R682 VTAIL.n39 VTAIL.n31 1.94878
R683 VTAIL.n55 VTAIL.n47 1.94878
R684 VTAIL.n23 VTAIL.n15 1.94878
R685 VTAIL VTAIL.n7 1.03283
R686 VTAIL VTAIL.n63 0.916448
R687 VTAIL.n47 VTAIL.n39 0.470328
R688 VTAIL.n15 VTAIL.n7 0.470328
R689 VP.n10 VP.n0 161.3
R690 VP.n9 VP.n8 161.3
R691 VP.n7 VP.n1 161.3
R692 VP.n6 VP.n5 161.3
R693 VP.n4 VP.n3 92.2184
R694 VP.n12 VP.n11 92.2184
R695 VP.n2 VP.t1 59.7307
R696 VP.n2 VP.t0 59.2093
R697 VP.n9 VP.n1 56.5617
R698 VP.n3 VP.n2 44.093
R699 VP.n5 VP.n1 24.5923
R700 VP.n10 VP.n9 24.5923
R701 VP.n4 VP.t3 24.4751
R702 VP.n11 VP.t2 24.4751
R703 VP.n5 VP.n4 18.6903
R704 VP.n11 VP.n10 18.6903
R705 VP.n6 VP.n3 0.278335
R706 VP.n12 VP.n0 0.278335
R707 VP.n7 VP.n6 0.189894
R708 VP.n8 VP.n7 0.189894
R709 VP.n8 VP.n0 0.189894
R710 VP VP.n12 0.153485
R711 VDD1 VDD1.n1 231.829
R712 VDD1 VDD1.n0 200.113
R713 VDD1.n0 VDD1.t2 16.5847
R714 VDD1.n0 VDD1.t3 16.5847
R715 VDD1.n1 VDD1.t0 16.5847
R716 VDD1.n1 VDD1.t1 16.5847
C0 VTAIL VDD2 2.74152f
C1 VN w_n2326_n1360# 3.61102f
C2 w_n2326_n1360# VP 3.90363f
C3 VN VDD1 0.154653f
C4 w_n2326_n1360# B 5.62268f
C5 VDD1 VP 1.19318f
C6 VDD2 w_n2326_n1360# 1.09028f
C7 VDD1 B 0.87284f
C8 VDD2 VDD1 0.866551f
C9 VN VP 3.85645f
C10 VTAIL w_n2326_n1360# 1.60641f
C11 VN B 0.846584f
C12 VTAIL VDD1 2.6918f
C13 VDD2 VN 0.990572f
C14 B VP 1.33609f
C15 VDD2 VP 0.358784f
C16 VDD2 B 0.914315f
C17 VTAIL VN 1.4029f
C18 VDD1 w_n2326_n1360# 1.04988f
C19 VTAIL VP 1.417f
C20 VTAIL B 1.39419f
C21 VDD2 VSUBS 0.550092f
C22 VDD1 VSUBS 2.950974f
C23 VTAIL VSUBS 0.381941f
C24 VN VSUBS 4.58387f
C25 VP VSUBS 1.423748f
C26 B VSUBS 2.689524f
C27 w_n2326_n1360# VSUBS 40.3887f
C28 VDD1.t2 VSUBS 0.030662f
C29 VDD1.t3 VSUBS 0.030662f
C30 VDD1.n0 VSUBS 0.126916f
C31 VDD1.t0 VSUBS 0.030662f
C32 VDD1.t1 VSUBS 0.030662f
C33 VDD1.n1 VSUBS 0.23885f
C34 VP.n0 VSUBS 0.064845f
C35 VP.t2 VSUBS 0.432763f
C36 VP.n1 VSUBS 0.071501f
C37 VP.t0 VSUBS 0.70435f
C38 VP.t1 VSUBS 0.708413f
C39 VP.n2 VSUBS 2.13287f
C40 VP.n3 VSUBS 2.02416f
C41 VP.t3 VSUBS 0.432763f
C42 VP.n4 VSUBS 0.360166f
C43 VP.n5 VSUBS 0.080406f
C44 VP.n6 VSUBS 0.064845f
C45 VP.n7 VSUBS 0.049187f
C46 VP.n8 VSUBS 0.049187f
C47 VP.n9 VSUBS 0.071501f
C48 VP.n10 VSUBS 0.080406f
C49 VP.n11 VSUBS 0.360166f
C50 VP.n12 VSUBS 0.060724f
C51 VTAIL.n0 VSUBS 0.018835f
C52 VTAIL.n1 VSUBS 0.048649f
C53 VTAIL.t5 VSUBS 0.048788f
C54 VTAIL.n2 VSUBS 0.04746f
C55 VTAIL.n3 VSUBS 0.014037f
C56 VTAIL.n4 VSUBS 0.009105f
C57 VTAIL.n5 VSUBS 0.114542f
C58 VTAIL.n6 VSUBS 0.026547f
C59 VTAIL.n7 VSUBS 0.095447f
C60 VTAIL.n8 VSUBS 0.018835f
C61 VTAIL.n9 VSUBS 0.048649f
C62 VTAIL.t1 VSUBS 0.048788f
C63 VTAIL.n10 VSUBS 0.04746f
C64 VTAIL.n11 VSUBS 0.014037f
C65 VTAIL.n12 VSUBS 0.009105f
C66 VTAIL.n13 VSUBS 0.114542f
C67 VTAIL.n14 VSUBS 0.026547f
C68 VTAIL.n15 VSUBS 0.145458f
C69 VTAIL.n16 VSUBS 0.018835f
C70 VTAIL.n17 VSUBS 0.048649f
C71 VTAIL.t2 VSUBS 0.048788f
C72 VTAIL.n18 VSUBS 0.04746f
C73 VTAIL.n19 VSUBS 0.014037f
C74 VTAIL.n20 VSUBS 0.009105f
C75 VTAIL.n21 VSUBS 0.114542f
C76 VTAIL.n22 VSUBS 0.026547f
C77 VTAIL.n23 VSUBS 0.548616f
C78 VTAIL.n24 VSUBS 0.018835f
C79 VTAIL.n25 VSUBS 0.048649f
C80 VTAIL.t7 VSUBS 0.048788f
C81 VTAIL.n26 VSUBS 0.04746f
C82 VTAIL.n27 VSUBS 0.014037f
C83 VTAIL.n28 VSUBS 0.009105f
C84 VTAIL.n29 VSUBS 0.114542f
C85 VTAIL.n30 VSUBS 0.026547f
C86 VTAIL.n31 VSUBS 0.548616f
C87 VTAIL.n32 VSUBS 0.018835f
C88 VTAIL.n33 VSUBS 0.048649f
C89 VTAIL.t6 VSUBS 0.048788f
C90 VTAIL.n34 VSUBS 0.04746f
C91 VTAIL.n35 VSUBS 0.014037f
C92 VTAIL.n36 VSUBS 0.009105f
C93 VTAIL.n37 VSUBS 0.114542f
C94 VTAIL.n38 VSUBS 0.026547f
C95 VTAIL.n39 VSUBS 0.145458f
C96 VTAIL.n40 VSUBS 0.018835f
C97 VTAIL.n41 VSUBS 0.048649f
C98 VTAIL.t0 VSUBS 0.048788f
C99 VTAIL.n42 VSUBS 0.04746f
C100 VTAIL.n43 VSUBS 0.014037f
C101 VTAIL.n44 VSUBS 0.009105f
C102 VTAIL.n45 VSUBS 0.114542f
C103 VTAIL.n46 VSUBS 0.026547f
C104 VTAIL.n47 VSUBS 0.145458f
C105 VTAIL.n48 VSUBS 0.018835f
C106 VTAIL.n49 VSUBS 0.048649f
C107 VTAIL.t3 VSUBS 0.048788f
C108 VTAIL.n50 VSUBS 0.04746f
C109 VTAIL.n51 VSUBS 0.014037f
C110 VTAIL.n52 VSUBS 0.009105f
C111 VTAIL.n53 VSUBS 0.114542f
C112 VTAIL.n54 VSUBS 0.026547f
C113 VTAIL.n55 VSUBS 0.548616f
C114 VTAIL.n56 VSUBS 0.018835f
C115 VTAIL.n57 VSUBS 0.048649f
C116 VTAIL.t4 VSUBS 0.048788f
C117 VTAIL.n58 VSUBS 0.04746f
C118 VTAIL.n59 VSUBS 0.014037f
C119 VTAIL.n60 VSUBS 0.009105f
C120 VTAIL.n61 VSUBS 0.114542f
C121 VTAIL.n62 VSUBS 0.026547f
C122 VTAIL.n63 VSUBS 0.49225f
C123 VDD2.t0 VSUBS 0.031515f
C124 VDD2.t1 VSUBS 0.031515f
C125 VDD2.n0 VSUBS 0.238241f
C126 VDD2.t3 VSUBS 0.031515f
C127 VDD2.t2 VSUBS 0.031515f
C128 VDD2.n1 VSUBS 0.130344f
C129 VDD2.n2 VSUBS 2.07324f
C130 VN.t2 VSUBS 0.675181f
C131 VN.t3 VSUBS 0.671308f
C132 VN.n0 VSUBS 0.473065f
C133 VN.t1 VSUBS 0.675181f
C134 VN.t0 VSUBS 0.671308f
C135 VN.n1 VSUBS 2.05701f
C136 B.n0 VSUBS 0.005699f
C137 B.n1 VSUBS 0.005699f
C138 B.n2 VSUBS 0.009012f
C139 B.n3 VSUBS 0.009012f
C140 B.n4 VSUBS 0.009012f
C141 B.n5 VSUBS 0.009012f
C142 B.n6 VSUBS 0.009012f
C143 B.n7 VSUBS 0.009012f
C144 B.n8 VSUBS 0.009012f
C145 B.n9 VSUBS 0.009012f
C146 B.n10 VSUBS 0.009012f
C147 B.n11 VSUBS 0.009012f
C148 B.n12 VSUBS 0.009012f
C149 B.n13 VSUBS 0.009012f
C150 B.n14 VSUBS 0.009012f
C151 B.n15 VSUBS 0.009012f
C152 B.n16 VSUBS 0.021357f
C153 B.n17 VSUBS 0.009012f
C154 B.n18 VSUBS 0.009012f
C155 B.n19 VSUBS 0.009012f
C156 B.n20 VSUBS 0.009012f
C157 B.n21 VSUBS 0.009012f
C158 B.t8 VSUBS 0.042946f
C159 B.t7 VSUBS 0.053354f
C160 B.t6 VSUBS 0.238927f
C161 B.n22 VSUBS 0.095562f
C162 B.n23 VSUBS 0.082048f
C163 B.n24 VSUBS 0.02088f
C164 B.n25 VSUBS 0.009012f
C165 B.n26 VSUBS 0.009012f
C166 B.n27 VSUBS 0.009012f
C167 B.n28 VSUBS 0.009012f
C168 B.n29 VSUBS 0.009012f
C169 B.t5 VSUBS 0.042946f
C170 B.t4 VSUBS 0.053354f
C171 B.t3 VSUBS 0.238927f
C172 B.n30 VSUBS 0.095562f
C173 B.n31 VSUBS 0.082048f
C174 B.n32 VSUBS 0.009012f
C175 B.n33 VSUBS 0.009012f
C176 B.n34 VSUBS 0.009012f
C177 B.n35 VSUBS 0.009012f
C178 B.n36 VSUBS 0.009012f
C179 B.n37 VSUBS 0.021357f
C180 B.n38 VSUBS 0.009012f
C181 B.n39 VSUBS 0.009012f
C182 B.n40 VSUBS 0.009012f
C183 B.n41 VSUBS 0.009012f
C184 B.n42 VSUBS 0.009012f
C185 B.n43 VSUBS 0.009012f
C186 B.n44 VSUBS 0.009012f
C187 B.n45 VSUBS 0.009012f
C188 B.n46 VSUBS 0.009012f
C189 B.n47 VSUBS 0.009012f
C190 B.n48 VSUBS 0.009012f
C191 B.n49 VSUBS 0.009012f
C192 B.n50 VSUBS 0.009012f
C193 B.n51 VSUBS 0.009012f
C194 B.n52 VSUBS 0.009012f
C195 B.n53 VSUBS 0.009012f
C196 B.n54 VSUBS 0.009012f
C197 B.n55 VSUBS 0.009012f
C198 B.n56 VSUBS 0.009012f
C199 B.n57 VSUBS 0.009012f
C200 B.n58 VSUBS 0.009012f
C201 B.n59 VSUBS 0.009012f
C202 B.n60 VSUBS 0.009012f
C203 B.n61 VSUBS 0.009012f
C204 B.n62 VSUBS 0.009012f
C205 B.n63 VSUBS 0.009012f
C206 B.n64 VSUBS 0.009012f
C207 B.n65 VSUBS 0.009012f
C208 B.n66 VSUBS 0.021357f
C209 B.n67 VSUBS 0.009012f
C210 B.n68 VSUBS 0.009012f
C211 B.n69 VSUBS 0.009012f
C212 B.n70 VSUBS 0.009012f
C213 B.n71 VSUBS 0.009012f
C214 B.t1 VSUBS 0.042946f
C215 B.t2 VSUBS 0.053354f
C216 B.t0 VSUBS 0.238927f
C217 B.n72 VSUBS 0.095562f
C218 B.n73 VSUBS 0.082048f
C219 B.n74 VSUBS 0.02088f
C220 B.n75 VSUBS 0.009012f
C221 B.n76 VSUBS 0.009012f
C222 B.n77 VSUBS 0.009012f
C223 B.n78 VSUBS 0.009012f
C224 B.n79 VSUBS 0.009012f
C225 B.t10 VSUBS 0.042946f
C226 B.t11 VSUBS 0.053354f
C227 B.t9 VSUBS 0.238927f
C228 B.n80 VSUBS 0.095562f
C229 B.n81 VSUBS 0.082048f
C230 B.n82 VSUBS 0.009012f
C231 B.n83 VSUBS 0.009012f
C232 B.n84 VSUBS 0.009012f
C233 B.n85 VSUBS 0.009012f
C234 B.n86 VSUBS 0.009012f
C235 B.n87 VSUBS 0.021357f
C236 B.n88 VSUBS 0.009012f
C237 B.n89 VSUBS 0.009012f
C238 B.n90 VSUBS 0.009012f
C239 B.n91 VSUBS 0.009012f
C240 B.n92 VSUBS 0.009012f
C241 B.n93 VSUBS 0.009012f
C242 B.n94 VSUBS 0.009012f
C243 B.n95 VSUBS 0.009012f
C244 B.n96 VSUBS 0.009012f
C245 B.n97 VSUBS 0.009012f
C246 B.n98 VSUBS 0.009012f
C247 B.n99 VSUBS 0.009012f
C248 B.n100 VSUBS 0.009012f
C249 B.n101 VSUBS 0.009012f
C250 B.n102 VSUBS 0.009012f
C251 B.n103 VSUBS 0.009012f
C252 B.n104 VSUBS 0.009012f
C253 B.n105 VSUBS 0.009012f
C254 B.n106 VSUBS 0.009012f
C255 B.n107 VSUBS 0.009012f
C256 B.n108 VSUBS 0.009012f
C257 B.n109 VSUBS 0.009012f
C258 B.n110 VSUBS 0.009012f
C259 B.n111 VSUBS 0.009012f
C260 B.n112 VSUBS 0.009012f
C261 B.n113 VSUBS 0.009012f
C262 B.n114 VSUBS 0.009012f
C263 B.n115 VSUBS 0.009012f
C264 B.n116 VSUBS 0.009012f
C265 B.n117 VSUBS 0.009012f
C266 B.n118 VSUBS 0.009012f
C267 B.n119 VSUBS 0.009012f
C268 B.n120 VSUBS 0.009012f
C269 B.n121 VSUBS 0.009012f
C270 B.n122 VSUBS 0.009012f
C271 B.n123 VSUBS 0.009012f
C272 B.n124 VSUBS 0.009012f
C273 B.n125 VSUBS 0.009012f
C274 B.n126 VSUBS 0.009012f
C275 B.n127 VSUBS 0.009012f
C276 B.n128 VSUBS 0.009012f
C277 B.n129 VSUBS 0.009012f
C278 B.n130 VSUBS 0.009012f
C279 B.n131 VSUBS 0.009012f
C280 B.n132 VSUBS 0.009012f
C281 B.n133 VSUBS 0.009012f
C282 B.n134 VSUBS 0.009012f
C283 B.n135 VSUBS 0.009012f
C284 B.n136 VSUBS 0.009012f
C285 B.n137 VSUBS 0.009012f
C286 B.n138 VSUBS 0.009012f
C287 B.n139 VSUBS 0.009012f
C288 B.n140 VSUBS 0.019992f
C289 B.n141 VSUBS 0.019992f
C290 B.n142 VSUBS 0.021357f
C291 B.n143 VSUBS 0.009012f
C292 B.n144 VSUBS 0.009012f
C293 B.n145 VSUBS 0.009012f
C294 B.n146 VSUBS 0.009012f
C295 B.n147 VSUBS 0.009012f
C296 B.n148 VSUBS 0.009012f
C297 B.n149 VSUBS 0.009012f
C298 B.n150 VSUBS 0.009012f
C299 B.n151 VSUBS 0.009012f
C300 B.n152 VSUBS 0.009012f
C301 B.n153 VSUBS 0.009012f
C302 B.n154 VSUBS 0.009012f
C303 B.n155 VSUBS 0.009012f
C304 B.n156 VSUBS 0.009012f
C305 B.n157 VSUBS 0.009012f
C306 B.n158 VSUBS 0.009012f
C307 B.n159 VSUBS 0.008482f
C308 B.n160 VSUBS 0.02088f
C309 B.n161 VSUBS 0.005036f
C310 B.n162 VSUBS 0.009012f
C311 B.n163 VSUBS 0.009012f
C312 B.n164 VSUBS 0.009012f
C313 B.n165 VSUBS 0.009012f
C314 B.n166 VSUBS 0.009012f
C315 B.n167 VSUBS 0.009012f
C316 B.n168 VSUBS 0.009012f
C317 B.n169 VSUBS 0.009012f
C318 B.n170 VSUBS 0.009012f
C319 B.n171 VSUBS 0.009012f
C320 B.n172 VSUBS 0.009012f
C321 B.n173 VSUBS 0.009012f
C322 B.n174 VSUBS 0.005036f
C323 B.n175 VSUBS 0.009012f
C324 B.n176 VSUBS 0.009012f
C325 B.n177 VSUBS 0.008482f
C326 B.n178 VSUBS 0.009012f
C327 B.n179 VSUBS 0.009012f
C328 B.n180 VSUBS 0.009012f
C329 B.n181 VSUBS 0.009012f
C330 B.n182 VSUBS 0.009012f
C331 B.n183 VSUBS 0.009012f
C332 B.n184 VSUBS 0.009012f
C333 B.n185 VSUBS 0.009012f
C334 B.n186 VSUBS 0.009012f
C335 B.n187 VSUBS 0.009012f
C336 B.n188 VSUBS 0.009012f
C337 B.n189 VSUBS 0.009012f
C338 B.n190 VSUBS 0.009012f
C339 B.n191 VSUBS 0.009012f
C340 B.n192 VSUBS 0.009012f
C341 B.n193 VSUBS 0.021357f
C342 B.n194 VSUBS 0.019992f
C343 B.n195 VSUBS 0.019992f
C344 B.n196 VSUBS 0.009012f
C345 B.n197 VSUBS 0.009012f
C346 B.n198 VSUBS 0.009012f
C347 B.n199 VSUBS 0.009012f
C348 B.n200 VSUBS 0.009012f
C349 B.n201 VSUBS 0.009012f
C350 B.n202 VSUBS 0.009012f
C351 B.n203 VSUBS 0.009012f
C352 B.n204 VSUBS 0.009012f
C353 B.n205 VSUBS 0.009012f
C354 B.n206 VSUBS 0.009012f
C355 B.n207 VSUBS 0.009012f
C356 B.n208 VSUBS 0.009012f
C357 B.n209 VSUBS 0.009012f
C358 B.n210 VSUBS 0.009012f
C359 B.n211 VSUBS 0.009012f
C360 B.n212 VSUBS 0.009012f
C361 B.n213 VSUBS 0.009012f
C362 B.n214 VSUBS 0.009012f
C363 B.n215 VSUBS 0.009012f
C364 B.n216 VSUBS 0.009012f
C365 B.n217 VSUBS 0.009012f
C366 B.n218 VSUBS 0.009012f
C367 B.n219 VSUBS 0.009012f
C368 B.n220 VSUBS 0.009012f
C369 B.n221 VSUBS 0.009012f
C370 B.n222 VSUBS 0.009012f
C371 B.n223 VSUBS 0.009012f
C372 B.n224 VSUBS 0.009012f
C373 B.n225 VSUBS 0.009012f
C374 B.n226 VSUBS 0.009012f
C375 B.n227 VSUBS 0.009012f
C376 B.n228 VSUBS 0.009012f
C377 B.n229 VSUBS 0.009012f
C378 B.n230 VSUBS 0.009012f
C379 B.n231 VSUBS 0.009012f
C380 B.n232 VSUBS 0.009012f
C381 B.n233 VSUBS 0.009012f
C382 B.n234 VSUBS 0.009012f
C383 B.n235 VSUBS 0.009012f
C384 B.n236 VSUBS 0.009012f
C385 B.n237 VSUBS 0.009012f
C386 B.n238 VSUBS 0.009012f
C387 B.n239 VSUBS 0.009012f
C388 B.n240 VSUBS 0.009012f
C389 B.n241 VSUBS 0.009012f
C390 B.n242 VSUBS 0.009012f
C391 B.n243 VSUBS 0.009012f
C392 B.n244 VSUBS 0.009012f
C393 B.n245 VSUBS 0.009012f
C394 B.n246 VSUBS 0.009012f
C395 B.n247 VSUBS 0.009012f
C396 B.n248 VSUBS 0.009012f
C397 B.n249 VSUBS 0.009012f
C398 B.n250 VSUBS 0.009012f
C399 B.n251 VSUBS 0.009012f
C400 B.n252 VSUBS 0.009012f
C401 B.n253 VSUBS 0.009012f
C402 B.n254 VSUBS 0.009012f
C403 B.n255 VSUBS 0.009012f
C404 B.n256 VSUBS 0.009012f
C405 B.n257 VSUBS 0.009012f
C406 B.n258 VSUBS 0.009012f
C407 B.n259 VSUBS 0.009012f
C408 B.n260 VSUBS 0.009012f
C409 B.n261 VSUBS 0.009012f
C410 B.n262 VSUBS 0.009012f
C411 B.n263 VSUBS 0.009012f
C412 B.n264 VSUBS 0.009012f
C413 B.n265 VSUBS 0.009012f
C414 B.n266 VSUBS 0.009012f
C415 B.n267 VSUBS 0.009012f
C416 B.n268 VSUBS 0.009012f
C417 B.n269 VSUBS 0.009012f
C418 B.n270 VSUBS 0.009012f
C419 B.n271 VSUBS 0.009012f
C420 B.n272 VSUBS 0.009012f
C421 B.n273 VSUBS 0.009012f
C422 B.n274 VSUBS 0.009012f
C423 B.n275 VSUBS 0.009012f
C424 B.n276 VSUBS 0.009012f
C425 B.n277 VSUBS 0.009012f
C426 B.n278 VSUBS 0.019992f
C427 B.n279 VSUBS 0.02109f
C428 B.n280 VSUBS 0.02026f
C429 B.n281 VSUBS 0.009012f
C430 B.n282 VSUBS 0.009012f
C431 B.n283 VSUBS 0.009012f
C432 B.n284 VSUBS 0.009012f
C433 B.n285 VSUBS 0.009012f
C434 B.n286 VSUBS 0.009012f
C435 B.n287 VSUBS 0.009012f
C436 B.n288 VSUBS 0.009012f
C437 B.n289 VSUBS 0.009012f
C438 B.n290 VSUBS 0.009012f
C439 B.n291 VSUBS 0.009012f
C440 B.n292 VSUBS 0.009012f
C441 B.n293 VSUBS 0.009012f
C442 B.n294 VSUBS 0.009012f
C443 B.n295 VSUBS 0.009012f
C444 B.n296 VSUBS 0.009012f
C445 B.n297 VSUBS 0.008482f
C446 B.n298 VSUBS 0.02088f
C447 B.n299 VSUBS 0.005036f
C448 B.n300 VSUBS 0.009012f
C449 B.n301 VSUBS 0.009012f
C450 B.n302 VSUBS 0.009012f
C451 B.n303 VSUBS 0.009012f
C452 B.n304 VSUBS 0.009012f
C453 B.n305 VSUBS 0.009012f
C454 B.n306 VSUBS 0.009012f
C455 B.n307 VSUBS 0.009012f
C456 B.n308 VSUBS 0.009012f
C457 B.n309 VSUBS 0.009012f
C458 B.n310 VSUBS 0.009012f
C459 B.n311 VSUBS 0.009012f
C460 B.n312 VSUBS 0.005036f
C461 B.n313 VSUBS 0.009012f
C462 B.n314 VSUBS 0.009012f
C463 B.n315 VSUBS 0.008482f
C464 B.n316 VSUBS 0.009012f
C465 B.n317 VSUBS 0.009012f
C466 B.n318 VSUBS 0.009012f
C467 B.n319 VSUBS 0.009012f
C468 B.n320 VSUBS 0.009012f
C469 B.n321 VSUBS 0.009012f
C470 B.n322 VSUBS 0.009012f
C471 B.n323 VSUBS 0.009012f
C472 B.n324 VSUBS 0.009012f
C473 B.n325 VSUBS 0.009012f
C474 B.n326 VSUBS 0.009012f
C475 B.n327 VSUBS 0.009012f
C476 B.n328 VSUBS 0.009012f
C477 B.n329 VSUBS 0.009012f
C478 B.n330 VSUBS 0.009012f
C479 B.n331 VSUBS 0.021357f
C480 B.n332 VSUBS 0.019992f
C481 B.n333 VSUBS 0.019992f
C482 B.n334 VSUBS 0.009012f
C483 B.n335 VSUBS 0.009012f
C484 B.n336 VSUBS 0.009012f
C485 B.n337 VSUBS 0.009012f
C486 B.n338 VSUBS 0.009012f
C487 B.n339 VSUBS 0.009012f
C488 B.n340 VSUBS 0.009012f
C489 B.n341 VSUBS 0.009012f
C490 B.n342 VSUBS 0.009012f
C491 B.n343 VSUBS 0.009012f
C492 B.n344 VSUBS 0.009012f
C493 B.n345 VSUBS 0.009012f
C494 B.n346 VSUBS 0.009012f
C495 B.n347 VSUBS 0.009012f
C496 B.n348 VSUBS 0.009012f
C497 B.n349 VSUBS 0.009012f
C498 B.n350 VSUBS 0.009012f
C499 B.n351 VSUBS 0.009012f
C500 B.n352 VSUBS 0.009012f
C501 B.n353 VSUBS 0.009012f
C502 B.n354 VSUBS 0.009012f
C503 B.n355 VSUBS 0.009012f
C504 B.n356 VSUBS 0.009012f
C505 B.n357 VSUBS 0.009012f
C506 B.n358 VSUBS 0.009012f
C507 B.n359 VSUBS 0.009012f
C508 B.n360 VSUBS 0.009012f
C509 B.n361 VSUBS 0.009012f
C510 B.n362 VSUBS 0.009012f
C511 B.n363 VSUBS 0.009012f
C512 B.n364 VSUBS 0.009012f
C513 B.n365 VSUBS 0.009012f
C514 B.n366 VSUBS 0.009012f
C515 B.n367 VSUBS 0.009012f
C516 B.n368 VSUBS 0.009012f
C517 B.n369 VSUBS 0.009012f
C518 B.n370 VSUBS 0.009012f
C519 B.n371 VSUBS 0.009012f
C520 B.n372 VSUBS 0.009012f
C521 B.n373 VSUBS 0.009012f
C522 B.n374 VSUBS 0.009012f
C523 B.n375 VSUBS 0.020406f
.ends

