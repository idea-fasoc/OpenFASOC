* NGSPICE file created from diff_pair_sample_1246.ext - technology: sky130A

.subckt diff_pair_sample_1246 VTAIL VN VP B VDD2 VDD1
X0 B.t19 B.t17 B.t18 B.t14 sky130_fd_pr__nfet_01v8 ad=4.5279 pd=24 as=0 ps=0 w=11.61 l=3.39
X1 VTAIL.t11 VP.t0 VDD1.t3 B.t4 sky130_fd_pr__nfet_01v8 ad=1.91565 pd=11.94 as=1.91565 ps=11.94 w=11.61 l=3.39
X2 VDD2.t5 VN.t0 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=4.5279 pd=24 as=1.91565 ps=11.94 w=11.61 l=3.39
X3 VTAIL.t10 VP.t1 VDD1.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=1.91565 pd=11.94 as=1.91565 ps=11.94 w=11.61 l=3.39
X4 VTAIL.t3 VN.t1 VDD2.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=1.91565 pd=11.94 as=1.91565 ps=11.94 w=11.61 l=3.39
X5 VDD1.t5 VP.t2 VTAIL.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=4.5279 pd=24 as=1.91565 ps=11.94 w=11.61 l=3.39
X6 B.t16 B.t13 B.t15 B.t14 sky130_fd_pr__nfet_01v8 ad=4.5279 pd=24 as=0 ps=0 w=11.61 l=3.39
X7 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=4.5279 pd=24 as=0 ps=0 w=11.61 l=3.39
X8 VDD2.t3 VN.t2 VTAIL.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=1.91565 pd=11.94 as=4.5279 ps=24 w=11.61 l=3.39
X9 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=4.5279 pd=24 as=0 ps=0 w=11.61 l=3.39
X10 VDD1.t4 VP.t3 VTAIL.t8 B.t0 sky130_fd_pr__nfet_01v8 ad=4.5279 pd=24 as=1.91565 ps=11.94 w=11.61 l=3.39
X11 VDD2.t2 VN.t3 VTAIL.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=1.91565 pd=11.94 as=4.5279 ps=24 w=11.61 l=3.39
X12 VDD1.t1 VP.t4 VTAIL.t7 B.t2 sky130_fd_pr__nfet_01v8 ad=1.91565 pd=11.94 as=4.5279 ps=24 w=11.61 l=3.39
X13 VTAIL.t2 VN.t4 VDD2.t1 B.t4 sky130_fd_pr__nfet_01v8 ad=1.91565 pd=11.94 as=1.91565 ps=11.94 w=11.61 l=3.39
X14 VDD2.t0 VN.t5 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=4.5279 pd=24 as=1.91565 ps=11.94 w=11.61 l=3.39
X15 VDD1.t0 VP.t5 VTAIL.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=1.91565 pd=11.94 as=4.5279 ps=24 w=11.61 l=3.39
R0 B.n884 B.n883 585
R1 B.n885 B.n884 585
R2 B.n325 B.n142 585
R3 B.n324 B.n323 585
R4 B.n322 B.n321 585
R5 B.n320 B.n319 585
R6 B.n318 B.n317 585
R7 B.n316 B.n315 585
R8 B.n314 B.n313 585
R9 B.n312 B.n311 585
R10 B.n310 B.n309 585
R11 B.n308 B.n307 585
R12 B.n306 B.n305 585
R13 B.n304 B.n303 585
R14 B.n302 B.n301 585
R15 B.n300 B.n299 585
R16 B.n298 B.n297 585
R17 B.n296 B.n295 585
R18 B.n294 B.n293 585
R19 B.n292 B.n291 585
R20 B.n290 B.n289 585
R21 B.n288 B.n287 585
R22 B.n286 B.n285 585
R23 B.n284 B.n283 585
R24 B.n282 B.n281 585
R25 B.n280 B.n279 585
R26 B.n278 B.n277 585
R27 B.n276 B.n275 585
R28 B.n274 B.n273 585
R29 B.n272 B.n271 585
R30 B.n270 B.n269 585
R31 B.n268 B.n267 585
R32 B.n266 B.n265 585
R33 B.n264 B.n263 585
R34 B.n262 B.n261 585
R35 B.n260 B.n259 585
R36 B.n258 B.n257 585
R37 B.n256 B.n255 585
R38 B.n254 B.n253 585
R39 B.n252 B.n251 585
R40 B.n250 B.n249 585
R41 B.n248 B.n247 585
R42 B.n246 B.n245 585
R43 B.n244 B.n243 585
R44 B.n242 B.n241 585
R45 B.n240 B.n239 585
R46 B.n238 B.n237 585
R47 B.n236 B.n235 585
R48 B.n234 B.n233 585
R49 B.n232 B.n231 585
R50 B.n230 B.n229 585
R51 B.n227 B.n226 585
R52 B.n225 B.n224 585
R53 B.n223 B.n222 585
R54 B.n221 B.n220 585
R55 B.n219 B.n218 585
R56 B.n217 B.n216 585
R57 B.n215 B.n214 585
R58 B.n213 B.n212 585
R59 B.n211 B.n210 585
R60 B.n209 B.n208 585
R61 B.n207 B.n206 585
R62 B.n205 B.n204 585
R63 B.n203 B.n202 585
R64 B.n201 B.n200 585
R65 B.n199 B.n198 585
R66 B.n197 B.n196 585
R67 B.n195 B.n194 585
R68 B.n193 B.n192 585
R69 B.n191 B.n190 585
R70 B.n189 B.n188 585
R71 B.n187 B.n186 585
R72 B.n185 B.n184 585
R73 B.n183 B.n182 585
R74 B.n181 B.n180 585
R75 B.n179 B.n178 585
R76 B.n177 B.n176 585
R77 B.n175 B.n174 585
R78 B.n173 B.n172 585
R79 B.n171 B.n170 585
R80 B.n169 B.n168 585
R81 B.n167 B.n166 585
R82 B.n165 B.n164 585
R83 B.n163 B.n162 585
R84 B.n161 B.n160 585
R85 B.n159 B.n158 585
R86 B.n157 B.n156 585
R87 B.n155 B.n154 585
R88 B.n153 B.n152 585
R89 B.n151 B.n150 585
R90 B.n149 B.n148 585
R91 B.n95 B.n94 585
R92 B.n882 B.n96 585
R93 B.n886 B.n96 585
R94 B.n881 B.n880 585
R95 B.n880 B.n92 585
R96 B.n879 B.n91 585
R97 B.n892 B.n91 585
R98 B.n878 B.n90 585
R99 B.n893 B.n90 585
R100 B.n877 B.n89 585
R101 B.n894 B.n89 585
R102 B.n876 B.n875 585
R103 B.n875 B.n85 585
R104 B.n874 B.n84 585
R105 B.n900 B.n84 585
R106 B.n873 B.n83 585
R107 B.n901 B.n83 585
R108 B.n872 B.n82 585
R109 B.n902 B.n82 585
R110 B.n871 B.n870 585
R111 B.n870 B.n78 585
R112 B.n869 B.n77 585
R113 B.n908 B.n77 585
R114 B.n868 B.n76 585
R115 B.n909 B.n76 585
R116 B.n867 B.n75 585
R117 B.n910 B.n75 585
R118 B.n866 B.n865 585
R119 B.n865 B.n71 585
R120 B.n864 B.n70 585
R121 B.n916 B.n70 585
R122 B.n863 B.n69 585
R123 B.n917 B.n69 585
R124 B.n862 B.n68 585
R125 B.n918 B.n68 585
R126 B.n861 B.n860 585
R127 B.n860 B.n64 585
R128 B.n859 B.n63 585
R129 B.n924 B.n63 585
R130 B.n858 B.n62 585
R131 B.n925 B.n62 585
R132 B.n857 B.n61 585
R133 B.n926 B.n61 585
R134 B.n856 B.n855 585
R135 B.n855 B.n57 585
R136 B.n854 B.n56 585
R137 B.n932 B.n56 585
R138 B.n853 B.n55 585
R139 B.n933 B.n55 585
R140 B.n852 B.n54 585
R141 B.n934 B.n54 585
R142 B.n851 B.n850 585
R143 B.n850 B.n50 585
R144 B.n849 B.n49 585
R145 B.n940 B.n49 585
R146 B.n848 B.n48 585
R147 B.n941 B.n48 585
R148 B.n847 B.n47 585
R149 B.n942 B.n47 585
R150 B.n846 B.n845 585
R151 B.n845 B.n43 585
R152 B.n844 B.n42 585
R153 B.n948 B.n42 585
R154 B.n843 B.n41 585
R155 B.n949 B.n41 585
R156 B.n842 B.n40 585
R157 B.n950 B.n40 585
R158 B.n841 B.n840 585
R159 B.n840 B.n39 585
R160 B.n839 B.n35 585
R161 B.n956 B.n35 585
R162 B.n838 B.n34 585
R163 B.n957 B.n34 585
R164 B.n837 B.n33 585
R165 B.n958 B.n33 585
R166 B.n836 B.n835 585
R167 B.n835 B.n29 585
R168 B.n834 B.n28 585
R169 B.n964 B.n28 585
R170 B.n833 B.n27 585
R171 B.n965 B.n27 585
R172 B.n832 B.n26 585
R173 B.n966 B.n26 585
R174 B.n831 B.n830 585
R175 B.n830 B.n22 585
R176 B.n829 B.n21 585
R177 B.n972 B.n21 585
R178 B.n828 B.n20 585
R179 B.n973 B.n20 585
R180 B.n827 B.n19 585
R181 B.n974 B.n19 585
R182 B.n826 B.n825 585
R183 B.n825 B.n15 585
R184 B.n824 B.n14 585
R185 B.n980 B.n14 585
R186 B.n823 B.n13 585
R187 B.n981 B.n13 585
R188 B.n822 B.n12 585
R189 B.n982 B.n12 585
R190 B.n821 B.n820 585
R191 B.n820 B.n8 585
R192 B.n819 B.n7 585
R193 B.n988 B.n7 585
R194 B.n818 B.n6 585
R195 B.n989 B.n6 585
R196 B.n817 B.n5 585
R197 B.n990 B.n5 585
R198 B.n816 B.n815 585
R199 B.n815 B.n4 585
R200 B.n814 B.n326 585
R201 B.n814 B.n813 585
R202 B.n804 B.n327 585
R203 B.n328 B.n327 585
R204 B.n806 B.n805 585
R205 B.n807 B.n806 585
R206 B.n803 B.n333 585
R207 B.n333 B.n332 585
R208 B.n802 B.n801 585
R209 B.n801 B.n800 585
R210 B.n335 B.n334 585
R211 B.n336 B.n335 585
R212 B.n793 B.n792 585
R213 B.n794 B.n793 585
R214 B.n791 B.n341 585
R215 B.n341 B.n340 585
R216 B.n790 B.n789 585
R217 B.n789 B.n788 585
R218 B.n343 B.n342 585
R219 B.n344 B.n343 585
R220 B.n781 B.n780 585
R221 B.n782 B.n781 585
R222 B.n779 B.n349 585
R223 B.n349 B.n348 585
R224 B.n778 B.n777 585
R225 B.n777 B.n776 585
R226 B.n351 B.n350 585
R227 B.n352 B.n351 585
R228 B.n769 B.n768 585
R229 B.n770 B.n769 585
R230 B.n767 B.n357 585
R231 B.n357 B.n356 585
R232 B.n766 B.n765 585
R233 B.n765 B.n764 585
R234 B.n359 B.n358 585
R235 B.n757 B.n359 585
R236 B.n756 B.n755 585
R237 B.n758 B.n756 585
R238 B.n754 B.n364 585
R239 B.n364 B.n363 585
R240 B.n753 B.n752 585
R241 B.n752 B.n751 585
R242 B.n366 B.n365 585
R243 B.n367 B.n366 585
R244 B.n744 B.n743 585
R245 B.n745 B.n744 585
R246 B.n742 B.n372 585
R247 B.n372 B.n371 585
R248 B.n741 B.n740 585
R249 B.n740 B.n739 585
R250 B.n374 B.n373 585
R251 B.n375 B.n374 585
R252 B.n732 B.n731 585
R253 B.n733 B.n732 585
R254 B.n730 B.n379 585
R255 B.n383 B.n379 585
R256 B.n729 B.n728 585
R257 B.n728 B.n727 585
R258 B.n381 B.n380 585
R259 B.n382 B.n381 585
R260 B.n720 B.n719 585
R261 B.n721 B.n720 585
R262 B.n718 B.n388 585
R263 B.n388 B.n387 585
R264 B.n717 B.n716 585
R265 B.n716 B.n715 585
R266 B.n390 B.n389 585
R267 B.n391 B.n390 585
R268 B.n708 B.n707 585
R269 B.n709 B.n708 585
R270 B.n706 B.n396 585
R271 B.n396 B.n395 585
R272 B.n705 B.n704 585
R273 B.n704 B.n703 585
R274 B.n398 B.n397 585
R275 B.n399 B.n398 585
R276 B.n696 B.n695 585
R277 B.n697 B.n696 585
R278 B.n694 B.n404 585
R279 B.n404 B.n403 585
R280 B.n693 B.n692 585
R281 B.n692 B.n691 585
R282 B.n406 B.n405 585
R283 B.n407 B.n406 585
R284 B.n684 B.n683 585
R285 B.n685 B.n684 585
R286 B.n682 B.n412 585
R287 B.n412 B.n411 585
R288 B.n681 B.n680 585
R289 B.n680 B.n679 585
R290 B.n414 B.n413 585
R291 B.n415 B.n414 585
R292 B.n672 B.n671 585
R293 B.n673 B.n672 585
R294 B.n670 B.n420 585
R295 B.n420 B.n419 585
R296 B.n669 B.n668 585
R297 B.n668 B.n667 585
R298 B.n422 B.n421 585
R299 B.n423 B.n422 585
R300 B.n660 B.n659 585
R301 B.n661 B.n660 585
R302 B.n426 B.n425 585
R303 B.n480 B.n479 585
R304 B.n481 B.n477 585
R305 B.n477 B.n427 585
R306 B.n483 B.n482 585
R307 B.n485 B.n476 585
R308 B.n488 B.n487 585
R309 B.n489 B.n475 585
R310 B.n491 B.n490 585
R311 B.n493 B.n474 585
R312 B.n496 B.n495 585
R313 B.n497 B.n473 585
R314 B.n499 B.n498 585
R315 B.n501 B.n472 585
R316 B.n504 B.n503 585
R317 B.n505 B.n471 585
R318 B.n507 B.n506 585
R319 B.n509 B.n470 585
R320 B.n512 B.n511 585
R321 B.n513 B.n469 585
R322 B.n515 B.n514 585
R323 B.n517 B.n468 585
R324 B.n520 B.n519 585
R325 B.n521 B.n467 585
R326 B.n523 B.n522 585
R327 B.n525 B.n466 585
R328 B.n528 B.n527 585
R329 B.n529 B.n465 585
R330 B.n531 B.n530 585
R331 B.n533 B.n464 585
R332 B.n536 B.n535 585
R333 B.n537 B.n463 585
R334 B.n539 B.n538 585
R335 B.n541 B.n462 585
R336 B.n544 B.n543 585
R337 B.n545 B.n461 585
R338 B.n547 B.n546 585
R339 B.n549 B.n460 585
R340 B.n552 B.n551 585
R341 B.n553 B.n459 585
R342 B.n555 B.n554 585
R343 B.n557 B.n458 585
R344 B.n560 B.n559 585
R345 B.n561 B.n454 585
R346 B.n563 B.n562 585
R347 B.n565 B.n453 585
R348 B.n568 B.n567 585
R349 B.n569 B.n452 585
R350 B.n571 B.n570 585
R351 B.n573 B.n451 585
R352 B.n576 B.n575 585
R353 B.n578 B.n448 585
R354 B.n580 B.n579 585
R355 B.n582 B.n447 585
R356 B.n585 B.n584 585
R357 B.n586 B.n446 585
R358 B.n588 B.n587 585
R359 B.n590 B.n445 585
R360 B.n593 B.n592 585
R361 B.n594 B.n444 585
R362 B.n596 B.n595 585
R363 B.n598 B.n443 585
R364 B.n601 B.n600 585
R365 B.n602 B.n442 585
R366 B.n604 B.n603 585
R367 B.n606 B.n441 585
R368 B.n609 B.n608 585
R369 B.n610 B.n440 585
R370 B.n612 B.n611 585
R371 B.n614 B.n439 585
R372 B.n617 B.n616 585
R373 B.n618 B.n438 585
R374 B.n620 B.n619 585
R375 B.n622 B.n437 585
R376 B.n625 B.n624 585
R377 B.n626 B.n436 585
R378 B.n628 B.n627 585
R379 B.n630 B.n435 585
R380 B.n633 B.n632 585
R381 B.n634 B.n434 585
R382 B.n636 B.n635 585
R383 B.n638 B.n433 585
R384 B.n641 B.n640 585
R385 B.n642 B.n432 585
R386 B.n644 B.n643 585
R387 B.n646 B.n431 585
R388 B.n649 B.n648 585
R389 B.n650 B.n430 585
R390 B.n652 B.n651 585
R391 B.n654 B.n429 585
R392 B.n657 B.n656 585
R393 B.n658 B.n428 585
R394 B.n663 B.n662 585
R395 B.n662 B.n661 585
R396 B.n664 B.n424 585
R397 B.n424 B.n423 585
R398 B.n666 B.n665 585
R399 B.n667 B.n666 585
R400 B.n418 B.n417 585
R401 B.n419 B.n418 585
R402 B.n675 B.n674 585
R403 B.n674 B.n673 585
R404 B.n676 B.n416 585
R405 B.n416 B.n415 585
R406 B.n678 B.n677 585
R407 B.n679 B.n678 585
R408 B.n410 B.n409 585
R409 B.n411 B.n410 585
R410 B.n687 B.n686 585
R411 B.n686 B.n685 585
R412 B.n688 B.n408 585
R413 B.n408 B.n407 585
R414 B.n690 B.n689 585
R415 B.n691 B.n690 585
R416 B.n402 B.n401 585
R417 B.n403 B.n402 585
R418 B.n699 B.n698 585
R419 B.n698 B.n697 585
R420 B.n700 B.n400 585
R421 B.n400 B.n399 585
R422 B.n702 B.n701 585
R423 B.n703 B.n702 585
R424 B.n394 B.n393 585
R425 B.n395 B.n394 585
R426 B.n711 B.n710 585
R427 B.n710 B.n709 585
R428 B.n712 B.n392 585
R429 B.n392 B.n391 585
R430 B.n714 B.n713 585
R431 B.n715 B.n714 585
R432 B.n386 B.n385 585
R433 B.n387 B.n386 585
R434 B.n723 B.n722 585
R435 B.n722 B.n721 585
R436 B.n724 B.n384 585
R437 B.n384 B.n382 585
R438 B.n726 B.n725 585
R439 B.n727 B.n726 585
R440 B.n378 B.n377 585
R441 B.n383 B.n378 585
R442 B.n735 B.n734 585
R443 B.n734 B.n733 585
R444 B.n736 B.n376 585
R445 B.n376 B.n375 585
R446 B.n738 B.n737 585
R447 B.n739 B.n738 585
R448 B.n370 B.n369 585
R449 B.n371 B.n370 585
R450 B.n747 B.n746 585
R451 B.n746 B.n745 585
R452 B.n748 B.n368 585
R453 B.n368 B.n367 585
R454 B.n750 B.n749 585
R455 B.n751 B.n750 585
R456 B.n362 B.n361 585
R457 B.n363 B.n362 585
R458 B.n760 B.n759 585
R459 B.n759 B.n758 585
R460 B.n761 B.n360 585
R461 B.n757 B.n360 585
R462 B.n763 B.n762 585
R463 B.n764 B.n763 585
R464 B.n355 B.n354 585
R465 B.n356 B.n355 585
R466 B.n772 B.n771 585
R467 B.n771 B.n770 585
R468 B.n773 B.n353 585
R469 B.n353 B.n352 585
R470 B.n775 B.n774 585
R471 B.n776 B.n775 585
R472 B.n347 B.n346 585
R473 B.n348 B.n347 585
R474 B.n784 B.n783 585
R475 B.n783 B.n782 585
R476 B.n785 B.n345 585
R477 B.n345 B.n344 585
R478 B.n787 B.n786 585
R479 B.n788 B.n787 585
R480 B.n339 B.n338 585
R481 B.n340 B.n339 585
R482 B.n796 B.n795 585
R483 B.n795 B.n794 585
R484 B.n797 B.n337 585
R485 B.n337 B.n336 585
R486 B.n799 B.n798 585
R487 B.n800 B.n799 585
R488 B.n331 B.n330 585
R489 B.n332 B.n331 585
R490 B.n809 B.n808 585
R491 B.n808 B.n807 585
R492 B.n810 B.n329 585
R493 B.n329 B.n328 585
R494 B.n812 B.n811 585
R495 B.n813 B.n812 585
R496 B.n2 B.n0 585
R497 B.n4 B.n2 585
R498 B.n3 B.n1 585
R499 B.n989 B.n3 585
R500 B.n987 B.n986 585
R501 B.n988 B.n987 585
R502 B.n985 B.n9 585
R503 B.n9 B.n8 585
R504 B.n984 B.n983 585
R505 B.n983 B.n982 585
R506 B.n11 B.n10 585
R507 B.n981 B.n11 585
R508 B.n979 B.n978 585
R509 B.n980 B.n979 585
R510 B.n977 B.n16 585
R511 B.n16 B.n15 585
R512 B.n976 B.n975 585
R513 B.n975 B.n974 585
R514 B.n18 B.n17 585
R515 B.n973 B.n18 585
R516 B.n971 B.n970 585
R517 B.n972 B.n971 585
R518 B.n969 B.n23 585
R519 B.n23 B.n22 585
R520 B.n968 B.n967 585
R521 B.n967 B.n966 585
R522 B.n25 B.n24 585
R523 B.n965 B.n25 585
R524 B.n963 B.n962 585
R525 B.n964 B.n963 585
R526 B.n961 B.n30 585
R527 B.n30 B.n29 585
R528 B.n960 B.n959 585
R529 B.n959 B.n958 585
R530 B.n32 B.n31 585
R531 B.n957 B.n32 585
R532 B.n955 B.n954 585
R533 B.n956 B.n955 585
R534 B.n953 B.n36 585
R535 B.n39 B.n36 585
R536 B.n952 B.n951 585
R537 B.n951 B.n950 585
R538 B.n38 B.n37 585
R539 B.n949 B.n38 585
R540 B.n947 B.n946 585
R541 B.n948 B.n947 585
R542 B.n945 B.n44 585
R543 B.n44 B.n43 585
R544 B.n944 B.n943 585
R545 B.n943 B.n942 585
R546 B.n46 B.n45 585
R547 B.n941 B.n46 585
R548 B.n939 B.n938 585
R549 B.n940 B.n939 585
R550 B.n937 B.n51 585
R551 B.n51 B.n50 585
R552 B.n936 B.n935 585
R553 B.n935 B.n934 585
R554 B.n53 B.n52 585
R555 B.n933 B.n53 585
R556 B.n931 B.n930 585
R557 B.n932 B.n931 585
R558 B.n929 B.n58 585
R559 B.n58 B.n57 585
R560 B.n928 B.n927 585
R561 B.n927 B.n926 585
R562 B.n60 B.n59 585
R563 B.n925 B.n60 585
R564 B.n923 B.n922 585
R565 B.n924 B.n923 585
R566 B.n921 B.n65 585
R567 B.n65 B.n64 585
R568 B.n920 B.n919 585
R569 B.n919 B.n918 585
R570 B.n67 B.n66 585
R571 B.n917 B.n67 585
R572 B.n915 B.n914 585
R573 B.n916 B.n915 585
R574 B.n913 B.n72 585
R575 B.n72 B.n71 585
R576 B.n912 B.n911 585
R577 B.n911 B.n910 585
R578 B.n74 B.n73 585
R579 B.n909 B.n74 585
R580 B.n907 B.n906 585
R581 B.n908 B.n907 585
R582 B.n905 B.n79 585
R583 B.n79 B.n78 585
R584 B.n904 B.n903 585
R585 B.n903 B.n902 585
R586 B.n81 B.n80 585
R587 B.n901 B.n81 585
R588 B.n899 B.n898 585
R589 B.n900 B.n899 585
R590 B.n897 B.n86 585
R591 B.n86 B.n85 585
R592 B.n896 B.n895 585
R593 B.n895 B.n894 585
R594 B.n88 B.n87 585
R595 B.n893 B.n88 585
R596 B.n891 B.n890 585
R597 B.n892 B.n891 585
R598 B.n889 B.n93 585
R599 B.n93 B.n92 585
R600 B.n888 B.n887 585
R601 B.n887 B.n886 585
R602 B.n992 B.n991 585
R603 B.n991 B.n990 585
R604 B.n662 B.n426 439.647
R605 B.n887 B.n95 439.647
R606 B.n660 B.n428 439.647
R607 B.n884 B.n96 439.647
R608 B.n449 B.t13 291.529
R609 B.n455 B.t17 291.529
R610 B.n146 B.t6 291.529
R611 B.n143 B.t10 291.529
R612 B.n885 B.n141 256.663
R613 B.n885 B.n140 256.663
R614 B.n885 B.n139 256.663
R615 B.n885 B.n138 256.663
R616 B.n885 B.n137 256.663
R617 B.n885 B.n136 256.663
R618 B.n885 B.n135 256.663
R619 B.n885 B.n134 256.663
R620 B.n885 B.n133 256.663
R621 B.n885 B.n132 256.663
R622 B.n885 B.n131 256.663
R623 B.n885 B.n130 256.663
R624 B.n885 B.n129 256.663
R625 B.n885 B.n128 256.663
R626 B.n885 B.n127 256.663
R627 B.n885 B.n126 256.663
R628 B.n885 B.n125 256.663
R629 B.n885 B.n124 256.663
R630 B.n885 B.n123 256.663
R631 B.n885 B.n122 256.663
R632 B.n885 B.n121 256.663
R633 B.n885 B.n120 256.663
R634 B.n885 B.n119 256.663
R635 B.n885 B.n118 256.663
R636 B.n885 B.n117 256.663
R637 B.n885 B.n116 256.663
R638 B.n885 B.n115 256.663
R639 B.n885 B.n114 256.663
R640 B.n885 B.n113 256.663
R641 B.n885 B.n112 256.663
R642 B.n885 B.n111 256.663
R643 B.n885 B.n110 256.663
R644 B.n885 B.n109 256.663
R645 B.n885 B.n108 256.663
R646 B.n885 B.n107 256.663
R647 B.n885 B.n106 256.663
R648 B.n885 B.n105 256.663
R649 B.n885 B.n104 256.663
R650 B.n885 B.n103 256.663
R651 B.n885 B.n102 256.663
R652 B.n885 B.n101 256.663
R653 B.n885 B.n100 256.663
R654 B.n885 B.n99 256.663
R655 B.n885 B.n98 256.663
R656 B.n885 B.n97 256.663
R657 B.n478 B.n427 256.663
R658 B.n484 B.n427 256.663
R659 B.n486 B.n427 256.663
R660 B.n492 B.n427 256.663
R661 B.n494 B.n427 256.663
R662 B.n500 B.n427 256.663
R663 B.n502 B.n427 256.663
R664 B.n508 B.n427 256.663
R665 B.n510 B.n427 256.663
R666 B.n516 B.n427 256.663
R667 B.n518 B.n427 256.663
R668 B.n524 B.n427 256.663
R669 B.n526 B.n427 256.663
R670 B.n532 B.n427 256.663
R671 B.n534 B.n427 256.663
R672 B.n540 B.n427 256.663
R673 B.n542 B.n427 256.663
R674 B.n548 B.n427 256.663
R675 B.n550 B.n427 256.663
R676 B.n556 B.n427 256.663
R677 B.n558 B.n427 256.663
R678 B.n564 B.n427 256.663
R679 B.n566 B.n427 256.663
R680 B.n572 B.n427 256.663
R681 B.n574 B.n427 256.663
R682 B.n581 B.n427 256.663
R683 B.n583 B.n427 256.663
R684 B.n589 B.n427 256.663
R685 B.n591 B.n427 256.663
R686 B.n597 B.n427 256.663
R687 B.n599 B.n427 256.663
R688 B.n605 B.n427 256.663
R689 B.n607 B.n427 256.663
R690 B.n613 B.n427 256.663
R691 B.n615 B.n427 256.663
R692 B.n621 B.n427 256.663
R693 B.n623 B.n427 256.663
R694 B.n629 B.n427 256.663
R695 B.n631 B.n427 256.663
R696 B.n637 B.n427 256.663
R697 B.n639 B.n427 256.663
R698 B.n645 B.n427 256.663
R699 B.n647 B.n427 256.663
R700 B.n653 B.n427 256.663
R701 B.n655 B.n427 256.663
R702 B.n662 B.n424 163.367
R703 B.n666 B.n424 163.367
R704 B.n666 B.n418 163.367
R705 B.n674 B.n418 163.367
R706 B.n674 B.n416 163.367
R707 B.n678 B.n416 163.367
R708 B.n678 B.n410 163.367
R709 B.n686 B.n410 163.367
R710 B.n686 B.n408 163.367
R711 B.n690 B.n408 163.367
R712 B.n690 B.n402 163.367
R713 B.n698 B.n402 163.367
R714 B.n698 B.n400 163.367
R715 B.n702 B.n400 163.367
R716 B.n702 B.n394 163.367
R717 B.n710 B.n394 163.367
R718 B.n710 B.n392 163.367
R719 B.n714 B.n392 163.367
R720 B.n714 B.n386 163.367
R721 B.n722 B.n386 163.367
R722 B.n722 B.n384 163.367
R723 B.n726 B.n384 163.367
R724 B.n726 B.n378 163.367
R725 B.n734 B.n378 163.367
R726 B.n734 B.n376 163.367
R727 B.n738 B.n376 163.367
R728 B.n738 B.n370 163.367
R729 B.n746 B.n370 163.367
R730 B.n746 B.n368 163.367
R731 B.n750 B.n368 163.367
R732 B.n750 B.n362 163.367
R733 B.n759 B.n362 163.367
R734 B.n759 B.n360 163.367
R735 B.n763 B.n360 163.367
R736 B.n763 B.n355 163.367
R737 B.n771 B.n355 163.367
R738 B.n771 B.n353 163.367
R739 B.n775 B.n353 163.367
R740 B.n775 B.n347 163.367
R741 B.n783 B.n347 163.367
R742 B.n783 B.n345 163.367
R743 B.n787 B.n345 163.367
R744 B.n787 B.n339 163.367
R745 B.n795 B.n339 163.367
R746 B.n795 B.n337 163.367
R747 B.n799 B.n337 163.367
R748 B.n799 B.n331 163.367
R749 B.n808 B.n331 163.367
R750 B.n808 B.n329 163.367
R751 B.n812 B.n329 163.367
R752 B.n812 B.n2 163.367
R753 B.n991 B.n2 163.367
R754 B.n991 B.n3 163.367
R755 B.n987 B.n3 163.367
R756 B.n987 B.n9 163.367
R757 B.n983 B.n9 163.367
R758 B.n983 B.n11 163.367
R759 B.n979 B.n11 163.367
R760 B.n979 B.n16 163.367
R761 B.n975 B.n16 163.367
R762 B.n975 B.n18 163.367
R763 B.n971 B.n18 163.367
R764 B.n971 B.n23 163.367
R765 B.n967 B.n23 163.367
R766 B.n967 B.n25 163.367
R767 B.n963 B.n25 163.367
R768 B.n963 B.n30 163.367
R769 B.n959 B.n30 163.367
R770 B.n959 B.n32 163.367
R771 B.n955 B.n32 163.367
R772 B.n955 B.n36 163.367
R773 B.n951 B.n36 163.367
R774 B.n951 B.n38 163.367
R775 B.n947 B.n38 163.367
R776 B.n947 B.n44 163.367
R777 B.n943 B.n44 163.367
R778 B.n943 B.n46 163.367
R779 B.n939 B.n46 163.367
R780 B.n939 B.n51 163.367
R781 B.n935 B.n51 163.367
R782 B.n935 B.n53 163.367
R783 B.n931 B.n53 163.367
R784 B.n931 B.n58 163.367
R785 B.n927 B.n58 163.367
R786 B.n927 B.n60 163.367
R787 B.n923 B.n60 163.367
R788 B.n923 B.n65 163.367
R789 B.n919 B.n65 163.367
R790 B.n919 B.n67 163.367
R791 B.n915 B.n67 163.367
R792 B.n915 B.n72 163.367
R793 B.n911 B.n72 163.367
R794 B.n911 B.n74 163.367
R795 B.n907 B.n74 163.367
R796 B.n907 B.n79 163.367
R797 B.n903 B.n79 163.367
R798 B.n903 B.n81 163.367
R799 B.n899 B.n81 163.367
R800 B.n899 B.n86 163.367
R801 B.n895 B.n86 163.367
R802 B.n895 B.n88 163.367
R803 B.n891 B.n88 163.367
R804 B.n891 B.n93 163.367
R805 B.n887 B.n93 163.367
R806 B.n479 B.n477 163.367
R807 B.n483 B.n477 163.367
R808 B.n487 B.n485 163.367
R809 B.n491 B.n475 163.367
R810 B.n495 B.n493 163.367
R811 B.n499 B.n473 163.367
R812 B.n503 B.n501 163.367
R813 B.n507 B.n471 163.367
R814 B.n511 B.n509 163.367
R815 B.n515 B.n469 163.367
R816 B.n519 B.n517 163.367
R817 B.n523 B.n467 163.367
R818 B.n527 B.n525 163.367
R819 B.n531 B.n465 163.367
R820 B.n535 B.n533 163.367
R821 B.n539 B.n463 163.367
R822 B.n543 B.n541 163.367
R823 B.n547 B.n461 163.367
R824 B.n551 B.n549 163.367
R825 B.n555 B.n459 163.367
R826 B.n559 B.n557 163.367
R827 B.n563 B.n454 163.367
R828 B.n567 B.n565 163.367
R829 B.n571 B.n452 163.367
R830 B.n575 B.n573 163.367
R831 B.n580 B.n448 163.367
R832 B.n584 B.n582 163.367
R833 B.n588 B.n446 163.367
R834 B.n592 B.n590 163.367
R835 B.n596 B.n444 163.367
R836 B.n600 B.n598 163.367
R837 B.n604 B.n442 163.367
R838 B.n608 B.n606 163.367
R839 B.n612 B.n440 163.367
R840 B.n616 B.n614 163.367
R841 B.n620 B.n438 163.367
R842 B.n624 B.n622 163.367
R843 B.n628 B.n436 163.367
R844 B.n632 B.n630 163.367
R845 B.n636 B.n434 163.367
R846 B.n640 B.n638 163.367
R847 B.n644 B.n432 163.367
R848 B.n648 B.n646 163.367
R849 B.n652 B.n430 163.367
R850 B.n656 B.n654 163.367
R851 B.n660 B.n422 163.367
R852 B.n668 B.n422 163.367
R853 B.n668 B.n420 163.367
R854 B.n672 B.n420 163.367
R855 B.n672 B.n414 163.367
R856 B.n680 B.n414 163.367
R857 B.n680 B.n412 163.367
R858 B.n684 B.n412 163.367
R859 B.n684 B.n406 163.367
R860 B.n692 B.n406 163.367
R861 B.n692 B.n404 163.367
R862 B.n696 B.n404 163.367
R863 B.n696 B.n398 163.367
R864 B.n704 B.n398 163.367
R865 B.n704 B.n396 163.367
R866 B.n708 B.n396 163.367
R867 B.n708 B.n390 163.367
R868 B.n716 B.n390 163.367
R869 B.n716 B.n388 163.367
R870 B.n720 B.n388 163.367
R871 B.n720 B.n381 163.367
R872 B.n728 B.n381 163.367
R873 B.n728 B.n379 163.367
R874 B.n732 B.n379 163.367
R875 B.n732 B.n374 163.367
R876 B.n740 B.n374 163.367
R877 B.n740 B.n372 163.367
R878 B.n744 B.n372 163.367
R879 B.n744 B.n366 163.367
R880 B.n752 B.n366 163.367
R881 B.n752 B.n364 163.367
R882 B.n756 B.n364 163.367
R883 B.n756 B.n359 163.367
R884 B.n765 B.n359 163.367
R885 B.n765 B.n357 163.367
R886 B.n769 B.n357 163.367
R887 B.n769 B.n351 163.367
R888 B.n777 B.n351 163.367
R889 B.n777 B.n349 163.367
R890 B.n781 B.n349 163.367
R891 B.n781 B.n343 163.367
R892 B.n789 B.n343 163.367
R893 B.n789 B.n341 163.367
R894 B.n793 B.n341 163.367
R895 B.n793 B.n335 163.367
R896 B.n801 B.n335 163.367
R897 B.n801 B.n333 163.367
R898 B.n806 B.n333 163.367
R899 B.n806 B.n327 163.367
R900 B.n814 B.n327 163.367
R901 B.n815 B.n814 163.367
R902 B.n815 B.n5 163.367
R903 B.n6 B.n5 163.367
R904 B.n7 B.n6 163.367
R905 B.n820 B.n7 163.367
R906 B.n820 B.n12 163.367
R907 B.n13 B.n12 163.367
R908 B.n14 B.n13 163.367
R909 B.n825 B.n14 163.367
R910 B.n825 B.n19 163.367
R911 B.n20 B.n19 163.367
R912 B.n21 B.n20 163.367
R913 B.n830 B.n21 163.367
R914 B.n830 B.n26 163.367
R915 B.n27 B.n26 163.367
R916 B.n28 B.n27 163.367
R917 B.n835 B.n28 163.367
R918 B.n835 B.n33 163.367
R919 B.n34 B.n33 163.367
R920 B.n35 B.n34 163.367
R921 B.n840 B.n35 163.367
R922 B.n840 B.n40 163.367
R923 B.n41 B.n40 163.367
R924 B.n42 B.n41 163.367
R925 B.n845 B.n42 163.367
R926 B.n845 B.n47 163.367
R927 B.n48 B.n47 163.367
R928 B.n49 B.n48 163.367
R929 B.n850 B.n49 163.367
R930 B.n850 B.n54 163.367
R931 B.n55 B.n54 163.367
R932 B.n56 B.n55 163.367
R933 B.n855 B.n56 163.367
R934 B.n855 B.n61 163.367
R935 B.n62 B.n61 163.367
R936 B.n63 B.n62 163.367
R937 B.n860 B.n63 163.367
R938 B.n860 B.n68 163.367
R939 B.n69 B.n68 163.367
R940 B.n70 B.n69 163.367
R941 B.n865 B.n70 163.367
R942 B.n865 B.n75 163.367
R943 B.n76 B.n75 163.367
R944 B.n77 B.n76 163.367
R945 B.n870 B.n77 163.367
R946 B.n870 B.n82 163.367
R947 B.n83 B.n82 163.367
R948 B.n84 B.n83 163.367
R949 B.n875 B.n84 163.367
R950 B.n875 B.n89 163.367
R951 B.n90 B.n89 163.367
R952 B.n91 B.n90 163.367
R953 B.n880 B.n91 163.367
R954 B.n880 B.n96 163.367
R955 B.n150 B.n149 163.367
R956 B.n154 B.n153 163.367
R957 B.n158 B.n157 163.367
R958 B.n162 B.n161 163.367
R959 B.n166 B.n165 163.367
R960 B.n170 B.n169 163.367
R961 B.n174 B.n173 163.367
R962 B.n178 B.n177 163.367
R963 B.n182 B.n181 163.367
R964 B.n186 B.n185 163.367
R965 B.n190 B.n189 163.367
R966 B.n194 B.n193 163.367
R967 B.n198 B.n197 163.367
R968 B.n202 B.n201 163.367
R969 B.n206 B.n205 163.367
R970 B.n210 B.n209 163.367
R971 B.n214 B.n213 163.367
R972 B.n218 B.n217 163.367
R973 B.n222 B.n221 163.367
R974 B.n226 B.n225 163.367
R975 B.n231 B.n230 163.367
R976 B.n235 B.n234 163.367
R977 B.n239 B.n238 163.367
R978 B.n243 B.n242 163.367
R979 B.n247 B.n246 163.367
R980 B.n251 B.n250 163.367
R981 B.n255 B.n254 163.367
R982 B.n259 B.n258 163.367
R983 B.n263 B.n262 163.367
R984 B.n267 B.n266 163.367
R985 B.n271 B.n270 163.367
R986 B.n275 B.n274 163.367
R987 B.n279 B.n278 163.367
R988 B.n283 B.n282 163.367
R989 B.n287 B.n286 163.367
R990 B.n291 B.n290 163.367
R991 B.n295 B.n294 163.367
R992 B.n299 B.n298 163.367
R993 B.n303 B.n302 163.367
R994 B.n307 B.n306 163.367
R995 B.n311 B.n310 163.367
R996 B.n315 B.n314 163.367
R997 B.n319 B.n318 163.367
R998 B.n323 B.n322 163.367
R999 B.n884 B.n142 163.367
R1000 B.n449 B.t16 140.96
R1001 B.n143 B.t11 140.96
R1002 B.n455 B.t19 140.946
R1003 B.n146 B.t8 140.946
R1004 B.n661 B.n427 74.9191
R1005 B.n886 B.n885 74.9191
R1006 B.n450 B.n449 72.146
R1007 B.n456 B.n455 72.146
R1008 B.n147 B.n146 72.146
R1009 B.n144 B.n143 72.146
R1010 B.n478 B.n426 71.676
R1011 B.n484 B.n483 71.676
R1012 B.n487 B.n486 71.676
R1013 B.n492 B.n491 71.676
R1014 B.n495 B.n494 71.676
R1015 B.n500 B.n499 71.676
R1016 B.n503 B.n502 71.676
R1017 B.n508 B.n507 71.676
R1018 B.n511 B.n510 71.676
R1019 B.n516 B.n515 71.676
R1020 B.n519 B.n518 71.676
R1021 B.n524 B.n523 71.676
R1022 B.n527 B.n526 71.676
R1023 B.n532 B.n531 71.676
R1024 B.n535 B.n534 71.676
R1025 B.n540 B.n539 71.676
R1026 B.n543 B.n542 71.676
R1027 B.n548 B.n547 71.676
R1028 B.n551 B.n550 71.676
R1029 B.n556 B.n555 71.676
R1030 B.n559 B.n558 71.676
R1031 B.n564 B.n563 71.676
R1032 B.n567 B.n566 71.676
R1033 B.n572 B.n571 71.676
R1034 B.n575 B.n574 71.676
R1035 B.n581 B.n580 71.676
R1036 B.n584 B.n583 71.676
R1037 B.n589 B.n588 71.676
R1038 B.n592 B.n591 71.676
R1039 B.n597 B.n596 71.676
R1040 B.n600 B.n599 71.676
R1041 B.n605 B.n604 71.676
R1042 B.n608 B.n607 71.676
R1043 B.n613 B.n612 71.676
R1044 B.n616 B.n615 71.676
R1045 B.n621 B.n620 71.676
R1046 B.n624 B.n623 71.676
R1047 B.n629 B.n628 71.676
R1048 B.n632 B.n631 71.676
R1049 B.n637 B.n636 71.676
R1050 B.n640 B.n639 71.676
R1051 B.n645 B.n644 71.676
R1052 B.n648 B.n647 71.676
R1053 B.n653 B.n652 71.676
R1054 B.n656 B.n655 71.676
R1055 B.n97 B.n95 71.676
R1056 B.n150 B.n98 71.676
R1057 B.n154 B.n99 71.676
R1058 B.n158 B.n100 71.676
R1059 B.n162 B.n101 71.676
R1060 B.n166 B.n102 71.676
R1061 B.n170 B.n103 71.676
R1062 B.n174 B.n104 71.676
R1063 B.n178 B.n105 71.676
R1064 B.n182 B.n106 71.676
R1065 B.n186 B.n107 71.676
R1066 B.n190 B.n108 71.676
R1067 B.n194 B.n109 71.676
R1068 B.n198 B.n110 71.676
R1069 B.n202 B.n111 71.676
R1070 B.n206 B.n112 71.676
R1071 B.n210 B.n113 71.676
R1072 B.n214 B.n114 71.676
R1073 B.n218 B.n115 71.676
R1074 B.n222 B.n116 71.676
R1075 B.n226 B.n117 71.676
R1076 B.n231 B.n118 71.676
R1077 B.n235 B.n119 71.676
R1078 B.n239 B.n120 71.676
R1079 B.n243 B.n121 71.676
R1080 B.n247 B.n122 71.676
R1081 B.n251 B.n123 71.676
R1082 B.n255 B.n124 71.676
R1083 B.n259 B.n125 71.676
R1084 B.n263 B.n126 71.676
R1085 B.n267 B.n127 71.676
R1086 B.n271 B.n128 71.676
R1087 B.n275 B.n129 71.676
R1088 B.n279 B.n130 71.676
R1089 B.n283 B.n131 71.676
R1090 B.n287 B.n132 71.676
R1091 B.n291 B.n133 71.676
R1092 B.n295 B.n134 71.676
R1093 B.n299 B.n135 71.676
R1094 B.n303 B.n136 71.676
R1095 B.n307 B.n137 71.676
R1096 B.n311 B.n138 71.676
R1097 B.n315 B.n139 71.676
R1098 B.n319 B.n140 71.676
R1099 B.n323 B.n141 71.676
R1100 B.n142 B.n141 71.676
R1101 B.n322 B.n140 71.676
R1102 B.n318 B.n139 71.676
R1103 B.n314 B.n138 71.676
R1104 B.n310 B.n137 71.676
R1105 B.n306 B.n136 71.676
R1106 B.n302 B.n135 71.676
R1107 B.n298 B.n134 71.676
R1108 B.n294 B.n133 71.676
R1109 B.n290 B.n132 71.676
R1110 B.n286 B.n131 71.676
R1111 B.n282 B.n130 71.676
R1112 B.n278 B.n129 71.676
R1113 B.n274 B.n128 71.676
R1114 B.n270 B.n127 71.676
R1115 B.n266 B.n126 71.676
R1116 B.n262 B.n125 71.676
R1117 B.n258 B.n124 71.676
R1118 B.n254 B.n123 71.676
R1119 B.n250 B.n122 71.676
R1120 B.n246 B.n121 71.676
R1121 B.n242 B.n120 71.676
R1122 B.n238 B.n119 71.676
R1123 B.n234 B.n118 71.676
R1124 B.n230 B.n117 71.676
R1125 B.n225 B.n116 71.676
R1126 B.n221 B.n115 71.676
R1127 B.n217 B.n114 71.676
R1128 B.n213 B.n113 71.676
R1129 B.n209 B.n112 71.676
R1130 B.n205 B.n111 71.676
R1131 B.n201 B.n110 71.676
R1132 B.n197 B.n109 71.676
R1133 B.n193 B.n108 71.676
R1134 B.n189 B.n107 71.676
R1135 B.n185 B.n106 71.676
R1136 B.n181 B.n105 71.676
R1137 B.n177 B.n104 71.676
R1138 B.n173 B.n103 71.676
R1139 B.n169 B.n102 71.676
R1140 B.n165 B.n101 71.676
R1141 B.n161 B.n100 71.676
R1142 B.n157 B.n99 71.676
R1143 B.n153 B.n98 71.676
R1144 B.n149 B.n97 71.676
R1145 B.n479 B.n478 71.676
R1146 B.n485 B.n484 71.676
R1147 B.n486 B.n475 71.676
R1148 B.n493 B.n492 71.676
R1149 B.n494 B.n473 71.676
R1150 B.n501 B.n500 71.676
R1151 B.n502 B.n471 71.676
R1152 B.n509 B.n508 71.676
R1153 B.n510 B.n469 71.676
R1154 B.n517 B.n516 71.676
R1155 B.n518 B.n467 71.676
R1156 B.n525 B.n524 71.676
R1157 B.n526 B.n465 71.676
R1158 B.n533 B.n532 71.676
R1159 B.n534 B.n463 71.676
R1160 B.n541 B.n540 71.676
R1161 B.n542 B.n461 71.676
R1162 B.n549 B.n548 71.676
R1163 B.n550 B.n459 71.676
R1164 B.n557 B.n556 71.676
R1165 B.n558 B.n454 71.676
R1166 B.n565 B.n564 71.676
R1167 B.n566 B.n452 71.676
R1168 B.n573 B.n572 71.676
R1169 B.n574 B.n448 71.676
R1170 B.n582 B.n581 71.676
R1171 B.n583 B.n446 71.676
R1172 B.n590 B.n589 71.676
R1173 B.n591 B.n444 71.676
R1174 B.n598 B.n597 71.676
R1175 B.n599 B.n442 71.676
R1176 B.n606 B.n605 71.676
R1177 B.n607 B.n440 71.676
R1178 B.n614 B.n613 71.676
R1179 B.n615 B.n438 71.676
R1180 B.n622 B.n621 71.676
R1181 B.n623 B.n436 71.676
R1182 B.n630 B.n629 71.676
R1183 B.n631 B.n434 71.676
R1184 B.n638 B.n637 71.676
R1185 B.n639 B.n432 71.676
R1186 B.n646 B.n645 71.676
R1187 B.n647 B.n430 71.676
R1188 B.n654 B.n653 71.676
R1189 B.n655 B.n428 71.676
R1190 B.n450 B.t15 68.8145
R1191 B.n144 B.t12 68.8145
R1192 B.n456 B.t18 68.7998
R1193 B.n147 B.t9 68.7998
R1194 B.n577 B.n450 59.5399
R1195 B.n457 B.n456 59.5399
R1196 B.n228 B.n147 59.5399
R1197 B.n145 B.n144 59.5399
R1198 B.n661 B.n423 44.3002
R1199 B.n667 B.n423 44.3002
R1200 B.n667 B.n419 44.3002
R1201 B.n673 B.n419 44.3002
R1202 B.n673 B.n415 44.3002
R1203 B.n679 B.n415 44.3002
R1204 B.n679 B.n411 44.3002
R1205 B.n685 B.n411 44.3002
R1206 B.n691 B.n407 44.3002
R1207 B.n691 B.n403 44.3002
R1208 B.n697 B.n403 44.3002
R1209 B.n697 B.n399 44.3002
R1210 B.n703 B.n399 44.3002
R1211 B.n703 B.n395 44.3002
R1212 B.n709 B.n395 44.3002
R1213 B.n709 B.n391 44.3002
R1214 B.n715 B.n391 44.3002
R1215 B.n715 B.n387 44.3002
R1216 B.n721 B.n387 44.3002
R1217 B.n721 B.n382 44.3002
R1218 B.n727 B.n382 44.3002
R1219 B.n727 B.n383 44.3002
R1220 B.n733 B.n375 44.3002
R1221 B.n739 B.n375 44.3002
R1222 B.n739 B.n371 44.3002
R1223 B.n745 B.n371 44.3002
R1224 B.n745 B.n367 44.3002
R1225 B.n751 B.n367 44.3002
R1226 B.n751 B.n363 44.3002
R1227 B.n758 B.n363 44.3002
R1228 B.n758 B.n757 44.3002
R1229 B.n764 B.n356 44.3002
R1230 B.n770 B.n356 44.3002
R1231 B.n770 B.n352 44.3002
R1232 B.n776 B.n352 44.3002
R1233 B.n776 B.n348 44.3002
R1234 B.n782 B.n348 44.3002
R1235 B.n782 B.n344 44.3002
R1236 B.n788 B.n344 44.3002
R1237 B.n788 B.n340 44.3002
R1238 B.n794 B.n340 44.3002
R1239 B.n800 B.n336 44.3002
R1240 B.n800 B.n332 44.3002
R1241 B.n807 B.n332 44.3002
R1242 B.n807 B.n328 44.3002
R1243 B.n813 B.n328 44.3002
R1244 B.n813 B.n4 44.3002
R1245 B.n990 B.n4 44.3002
R1246 B.n990 B.n989 44.3002
R1247 B.n989 B.n988 44.3002
R1248 B.n988 B.n8 44.3002
R1249 B.n982 B.n8 44.3002
R1250 B.n982 B.n981 44.3002
R1251 B.n981 B.n980 44.3002
R1252 B.n980 B.n15 44.3002
R1253 B.n974 B.n973 44.3002
R1254 B.n973 B.n972 44.3002
R1255 B.n972 B.n22 44.3002
R1256 B.n966 B.n22 44.3002
R1257 B.n966 B.n965 44.3002
R1258 B.n965 B.n964 44.3002
R1259 B.n964 B.n29 44.3002
R1260 B.n958 B.n29 44.3002
R1261 B.n958 B.n957 44.3002
R1262 B.n957 B.n956 44.3002
R1263 B.n950 B.n39 44.3002
R1264 B.n950 B.n949 44.3002
R1265 B.n949 B.n948 44.3002
R1266 B.n948 B.n43 44.3002
R1267 B.n942 B.n43 44.3002
R1268 B.n942 B.n941 44.3002
R1269 B.n941 B.n940 44.3002
R1270 B.n940 B.n50 44.3002
R1271 B.n934 B.n50 44.3002
R1272 B.n933 B.n932 44.3002
R1273 B.n932 B.n57 44.3002
R1274 B.n926 B.n57 44.3002
R1275 B.n926 B.n925 44.3002
R1276 B.n925 B.n924 44.3002
R1277 B.n924 B.n64 44.3002
R1278 B.n918 B.n64 44.3002
R1279 B.n918 B.n917 44.3002
R1280 B.n917 B.n916 44.3002
R1281 B.n916 B.n71 44.3002
R1282 B.n910 B.n71 44.3002
R1283 B.n910 B.n909 44.3002
R1284 B.n909 B.n908 44.3002
R1285 B.n908 B.n78 44.3002
R1286 B.n902 B.n901 44.3002
R1287 B.n901 B.n900 44.3002
R1288 B.n900 B.n85 44.3002
R1289 B.n894 B.n85 44.3002
R1290 B.n894 B.n893 44.3002
R1291 B.n893 B.n892 44.3002
R1292 B.n892 B.n92 44.3002
R1293 B.n886 B.n92 44.3002
R1294 B.n757 B.t1 43.6487
R1295 B.n39 B.t4 43.6487
R1296 B.n733 B.t5 42.3458
R1297 B.n934 B.t2 42.3458
R1298 B.n794 B.t3 41.0428
R1299 B.n974 B.t0 41.0428
R1300 B.n685 B.t14 39.7399
R1301 B.n902 B.t7 39.7399
R1302 B.n883 B.n882 28.5664
R1303 B.n888 B.n94 28.5664
R1304 B.n659 B.n658 28.5664
R1305 B.n663 B.n425 28.5664
R1306 B B.n992 18.0485
R1307 B.n148 B.n94 10.6151
R1308 B.n151 B.n148 10.6151
R1309 B.n152 B.n151 10.6151
R1310 B.n155 B.n152 10.6151
R1311 B.n156 B.n155 10.6151
R1312 B.n159 B.n156 10.6151
R1313 B.n160 B.n159 10.6151
R1314 B.n163 B.n160 10.6151
R1315 B.n164 B.n163 10.6151
R1316 B.n167 B.n164 10.6151
R1317 B.n168 B.n167 10.6151
R1318 B.n171 B.n168 10.6151
R1319 B.n172 B.n171 10.6151
R1320 B.n175 B.n172 10.6151
R1321 B.n176 B.n175 10.6151
R1322 B.n179 B.n176 10.6151
R1323 B.n180 B.n179 10.6151
R1324 B.n183 B.n180 10.6151
R1325 B.n184 B.n183 10.6151
R1326 B.n187 B.n184 10.6151
R1327 B.n188 B.n187 10.6151
R1328 B.n191 B.n188 10.6151
R1329 B.n192 B.n191 10.6151
R1330 B.n195 B.n192 10.6151
R1331 B.n196 B.n195 10.6151
R1332 B.n199 B.n196 10.6151
R1333 B.n200 B.n199 10.6151
R1334 B.n203 B.n200 10.6151
R1335 B.n204 B.n203 10.6151
R1336 B.n207 B.n204 10.6151
R1337 B.n208 B.n207 10.6151
R1338 B.n211 B.n208 10.6151
R1339 B.n212 B.n211 10.6151
R1340 B.n215 B.n212 10.6151
R1341 B.n216 B.n215 10.6151
R1342 B.n219 B.n216 10.6151
R1343 B.n220 B.n219 10.6151
R1344 B.n223 B.n220 10.6151
R1345 B.n224 B.n223 10.6151
R1346 B.n227 B.n224 10.6151
R1347 B.n232 B.n229 10.6151
R1348 B.n233 B.n232 10.6151
R1349 B.n236 B.n233 10.6151
R1350 B.n237 B.n236 10.6151
R1351 B.n240 B.n237 10.6151
R1352 B.n241 B.n240 10.6151
R1353 B.n244 B.n241 10.6151
R1354 B.n245 B.n244 10.6151
R1355 B.n249 B.n248 10.6151
R1356 B.n252 B.n249 10.6151
R1357 B.n253 B.n252 10.6151
R1358 B.n256 B.n253 10.6151
R1359 B.n257 B.n256 10.6151
R1360 B.n260 B.n257 10.6151
R1361 B.n261 B.n260 10.6151
R1362 B.n264 B.n261 10.6151
R1363 B.n265 B.n264 10.6151
R1364 B.n268 B.n265 10.6151
R1365 B.n269 B.n268 10.6151
R1366 B.n272 B.n269 10.6151
R1367 B.n273 B.n272 10.6151
R1368 B.n276 B.n273 10.6151
R1369 B.n277 B.n276 10.6151
R1370 B.n280 B.n277 10.6151
R1371 B.n281 B.n280 10.6151
R1372 B.n284 B.n281 10.6151
R1373 B.n285 B.n284 10.6151
R1374 B.n288 B.n285 10.6151
R1375 B.n289 B.n288 10.6151
R1376 B.n292 B.n289 10.6151
R1377 B.n293 B.n292 10.6151
R1378 B.n296 B.n293 10.6151
R1379 B.n297 B.n296 10.6151
R1380 B.n300 B.n297 10.6151
R1381 B.n301 B.n300 10.6151
R1382 B.n304 B.n301 10.6151
R1383 B.n305 B.n304 10.6151
R1384 B.n308 B.n305 10.6151
R1385 B.n309 B.n308 10.6151
R1386 B.n312 B.n309 10.6151
R1387 B.n313 B.n312 10.6151
R1388 B.n316 B.n313 10.6151
R1389 B.n317 B.n316 10.6151
R1390 B.n320 B.n317 10.6151
R1391 B.n321 B.n320 10.6151
R1392 B.n324 B.n321 10.6151
R1393 B.n325 B.n324 10.6151
R1394 B.n883 B.n325 10.6151
R1395 B.n659 B.n421 10.6151
R1396 B.n669 B.n421 10.6151
R1397 B.n670 B.n669 10.6151
R1398 B.n671 B.n670 10.6151
R1399 B.n671 B.n413 10.6151
R1400 B.n681 B.n413 10.6151
R1401 B.n682 B.n681 10.6151
R1402 B.n683 B.n682 10.6151
R1403 B.n683 B.n405 10.6151
R1404 B.n693 B.n405 10.6151
R1405 B.n694 B.n693 10.6151
R1406 B.n695 B.n694 10.6151
R1407 B.n695 B.n397 10.6151
R1408 B.n705 B.n397 10.6151
R1409 B.n706 B.n705 10.6151
R1410 B.n707 B.n706 10.6151
R1411 B.n707 B.n389 10.6151
R1412 B.n717 B.n389 10.6151
R1413 B.n718 B.n717 10.6151
R1414 B.n719 B.n718 10.6151
R1415 B.n719 B.n380 10.6151
R1416 B.n729 B.n380 10.6151
R1417 B.n730 B.n729 10.6151
R1418 B.n731 B.n730 10.6151
R1419 B.n731 B.n373 10.6151
R1420 B.n741 B.n373 10.6151
R1421 B.n742 B.n741 10.6151
R1422 B.n743 B.n742 10.6151
R1423 B.n743 B.n365 10.6151
R1424 B.n753 B.n365 10.6151
R1425 B.n754 B.n753 10.6151
R1426 B.n755 B.n754 10.6151
R1427 B.n755 B.n358 10.6151
R1428 B.n766 B.n358 10.6151
R1429 B.n767 B.n766 10.6151
R1430 B.n768 B.n767 10.6151
R1431 B.n768 B.n350 10.6151
R1432 B.n778 B.n350 10.6151
R1433 B.n779 B.n778 10.6151
R1434 B.n780 B.n779 10.6151
R1435 B.n780 B.n342 10.6151
R1436 B.n790 B.n342 10.6151
R1437 B.n791 B.n790 10.6151
R1438 B.n792 B.n791 10.6151
R1439 B.n792 B.n334 10.6151
R1440 B.n802 B.n334 10.6151
R1441 B.n803 B.n802 10.6151
R1442 B.n805 B.n803 10.6151
R1443 B.n805 B.n804 10.6151
R1444 B.n804 B.n326 10.6151
R1445 B.n816 B.n326 10.6151
R1446 B.n817 B.n816 10.6151
R1447 B.n818 B.n817 10.6151
R1448 B.n819 B.n818 10.6151
R1449 B.n821 B.n819 10.6151
R1450 B.n822 B.n821 10.6151
R1451 B.n823 B.n822 10.6151
R1452 B.n824 B.n823 10.6151
R1453 B.n826 B.n824 10.6151
R1454 B.n827 B.n826 10.6151
R1455 B.n828 B.n827 10.6151
R1456 B.n829 B.n828 10.6151
R1457 B.n831 B.n829 10.6151
R1458 B.n832 B.n831 10.6151
R1459 B.n833 B.n832 10.6151
R1460 B.n834 B.n833 10.6151
R1461 B.n836 B.n834 10.6151
R1462 B.n837 B.n836 10.6151
R1463 B.n838 B.n837 10.6151
R1464 B.n839 B.n838 10.6151
R1465 B.n841 B.n839 10.6151
R1466 B.n842 B.n841 10.6151
R1467 B.n843 B.n842 10.6151
R1468 B.n844 B.n843 10.6151
R1469 B.n846 B.n844 10.6151
R1470 B.n847 B.n846 10.6151
R1471 B.n848 B.n847 10.6151
R1472 B.n849 B.n848 10.6151
R1473 B.n851 B.n849 10.6151
R1474 B.n852 B.n851 10.6151
R1475 B.n853 B.n852 10.6151
R1476 B.n854 B.n853 10.6151
R1477 B.n856 B.n854 10.6151
R1478 B.n857 B.n856 10.6151
R1479 B.n858 B.n857 10.6151
R1480 B.n859 B.n858 10.6151
R1481 B.n861 B.n859 10.6151
R1482 B.n862 B.n861 10.6151
R1483 B.n863 B.n862 10.6151
R1484 B.n864 B.n863 10.6151
R1485 B.n866 B.n864 10.6151
R1486 B.n867 B.n866 10.6151
R1487 B.n868 B.n867 10.6151
R1488 B.n869 B.n868 10.6151
R1489 B.n871 B.n869 10.6151
R1490 B.n872 B.n871 10.6151
R1491 B.n873 B.n872 10.6151
R1492 B.n874 B.n873 10.6151
R1493 B.n876 B.n874 10.6151
R1494 B.n877 B.n876 10.6151
R1495 B.n878 B.n877 10.6151
R1496 B.n879 B.n878 10.6151
R1497 B.n881 B.n879 10.6151
R1498 B.n882 B.n881 10.6151
R1499 B.n480 B.n425 10.6151
R1500 B.n481 B.n480 10.6151
R1501 B.n482 B.n481 10.6151
R1502 B.n482 B.n476 10.6151
R1503 B.n488 B.n476 10.6151
R1504 B.n489 B.n488 10.6151
R1505 B.n490 B.n489 10.6151
R1506 B.n490 B.n474 10.6151
R1507 B.n496 B.n474 10.6151
R1508 B.n497 B.n496 10.6151
R1509 B.n498 B.n497 10.6151
R1510 B.n498 B.n472 10.6151
R1511 B.n504 B.n472 10.6151
R1512 B.n505 B.n504 10.6151
R1513 B.n506 B.n505 10.6151
R1514 B.n506 B.n470 10.6151
R1515 B.n512 B.n470 10.6151
R1516 B.n513 B.n512 10.6151
R1517 B.n514 B.n513 10.6151
R1518 B.n514 B.n468 10.6151
R1519 B.n520 B.n468 10.6151
R1520 B.n521 B.n520 10.6151
R1521 B.n522 B.n521 10.6151
R1522 B.n522 B.n466 10.6151
R1523 B.n528 B.n466 10.6151
R1524 B.n529 B.n528 10.6151
R1525 B.n530 B.n529 10.6151
R1526 B.n530 B.n464 10.6151
R1527 B.n536 B.n464 10.6151
R1528 B.n537 B.n536 10.6151
R1529 B.n538 B.n537 10.6151
R1530 B.n538 B.n462 10.6151
R1531 B.n544 B.n462 10.6151
R1532 B.n545 B.n544 10.6151
R1533 B.n546 B.n545 10.6151
R1534 B.n546 B.n460 10.6151
R1535 B.n552 B.n460 10.6151
R1536 B.n553 B.n552 10.6151
R1537 B.n554 B.n553 10.6151
R1538 B.n554 B.n458 10.6151
R1539 B.n561 B.n560 10.6151
R1540 B.n562 B.n561 10.6151
R1541 B.n562 B.n453 10.6151
R1542 B.n568 B.n453 10.6151
R1543 B.n569 B.n568 10.6151
R1544 B.n570 B.n569 10.6151
R1545 B.n570 B.n451 10.6151
R1546 B.n576 B.n451 10.6151
R1547 B.n579 B.n578 10.6151
R1548 B.n579 B.n447 10.6151
R1549 B.n585 B.n447 10.6151
R1550 B.n586 B.n585 10.6151
R1551 B.n587 B.n586 10.6151
R1552 B.n587 B.n445 10.6151
R1553 B.n593 B.n445 10.6151
R1554 B.n594 B.n593 10.6151
R1555 B.n595 B.n594 10.6151
R1556 B.n595 B.n443 10.6151
R1557 B.n601 B.n443 10.6151
R1558 B.n602 B.n601 10.6151
R1559 B.n603 B.n602 10.6151
R1560 B.n603 B.n441 10.6151
R1561 B.n609 B.n441 10.6151
R1562 B.n610 B.n609 10.6151
R1563 B.n611 B.n610 10.6151
R1564 B.n611 B.n439 10.6151
R1565 B.n617 B.n439 10.6151
R1566 B.n618 B.n617 10.6151
R1567 B.n619 B.n618 10.6151
R1568 B.n619 B.n437 10.6151
R1569 B.n625 B.n437 10.6151
R1570 B.n626 B.n625 10.6151
R1571 B.n627 B.n626 10.6151
R1572 B.n627 B.n435 10.6151
R1573 B.n633 B.n435 10.6151
R1574 B.n634 B.n633 10.6151
R1575 B.n635 B.n634 10.6151
R1576 B.n635 B.n433 10.6151
R1577 B.n641 B.n433 10.6151
R1578 B.n642 B.n641 10.6151
R1579 B.n643 B.n642 10.6151
R1580 B.n643 B.n431 10.6151
R1581 B.n649 B.n431 10.6151
R1582 B.n650 B.n649 10.6151
R1583 B.n651 B.n650 10.6151
R1584 B.n651 B.n429 10.6151
R1585 B.n657 B.n429 10.6151
R1586 B.n658 B.n657 10.6151
R1587 B.n664 B.n663 10.6151
R1588 B.n665 B.n664 10.6151
R1589 B.n665 B.n417 10.6151
R1590 B.n675 B.n417 10.6151
R1591 B.n676 B.n675 10.6151
R1592 B.n677 B.n676 10.6151
R1593 B.n677 B.n409 10.6151
R1594 B.n687 B.n409 10.6151
R1595 B.n688 B.n687 10.6151
R1596 B.n689 B.n688 10.6151
R1597 B.n689 B.n401 10.6151
R1598 B.n699 B.n401 10.6151
R1599 B.n700 B.n699 10.6151
R1600 B.n701 B.n700 10.6151
R1601 B.n701 B.n393 10.6151
R1602 B.n711 B.n393 10.6151
R1603 B.n712 B.n711 10.6151
R1604 B.n713 B.n712 10.6151
R1605 B.n713 B.n385 10.6151
R1606 B.n723 B.n385 10.6151
R1607 B.n724 B.n723 10.6151
R1608 B.n725 B.n724 10.6151
R1609 B.n725 B.n377 10.6151
R1610 B.n735 B.n377 10.6151
R1611 B.n736 B.n735 10.6151
R1612 B.n737 B.n736 10.6151
R1613 B.n737 B.n369 10.6151
R1614 B.n747 B.n369 10.6151
R1615 B.n748 B.n747 10.6151
R1616 B.n749 B.n748 10.6151
R1617 B.n749 B.n361 10.6151
R1618 B.n760 B.n361 10.6151
R1619 B.n761 B.n760 10.6151
R1620 B.n762 B.n761 10.6151
R1621 B.n762 B.n354 10.6151
R1622 B.n772 B.n354 10.6151
R1623 B.n773 B.n772 10.6151
R1624 B.n774 B.n773 10.6151
R1625 B.n774 B.n346 10.6151
R1626 B.n784 B.n346 10.6151
R1627 B.n785 B.n784 10.6151
R1628 B.n786 B.n785 10.6151
R1629 B.n786 B.n338 10.6151
R1630 B.n796 B.n338 10.6151
R1631 B.n797 B.n796 10.6151
R1632 B.n798 B.n797 10.6151
R1633 B.n798 B.n330 10.6151
R1634 B.n809 B.n330 10.6151
R1635 B.n810 B.n809 10.6151
R1636 B.n811 B.n810 10.6151
R1637 B.n811 B.n0 10.6151
R1638 B.n986 B.n1 10.6151
R1639 B.n986 B.n985 10.6151
R1640 B.n985 B.n984 10.6151
R1641 B.n984 B.n10 10.6151
R1642 B.n978 B.n10 10.6151
R1643 B.n978 B.n977 10.6151
R1644 B.n977 B.n976 10.6151
R1645 B.n976 B.n17 10.6151
R1646 B.n970 B.n17 10.6151
R1647 B.n970 B.n969 10.6151
R1648 B.n969 B.n968 10.6151
R1649 B.n968 B.n24 10.6151
R1650 B.n962 B.n24 10.6151
R1651 B.n962 B.n961 10.6151
R1652 B.n961 B.n960 10.6151
R1653 B.n960 B.n31 10.6151
R1654 B.n954 B.n31 10.6151
R1655 B.n954 B.n953 10.6151
R1656 B.n953 B.n952 10.6151
R1657 B.n952 B.n37 10.6151
R1658 B.n946 B.n37 10.6151
R1659 B.n946 B.n945 10.6151
R1660 B.n945 B.n944 10.6151
R1661 B.n944 B.n45 10.6151
R1662 B.n938 B.n45 10.6151
R1663 B.n938 B.n937 10.6151
R1664 B.n937 B.n936 10.6151
R1665 B.n936 B.n52 10.6151
R1666 B.n930 B.n52 10.6151
R1667 B.n930 B.n929 10.6151
R1668 B.n929 B.n928 10.6151
R1669 B.n928 B.n59 10.6151
R1670 B.n922 B.n59 10.6151
R1671 B.n922 B.n921 10.6151
R1672 B.n921 B.n920 10.6151
R1673 B.n920 B.n66 10.6151
R1674 B.n914 B.n66 10.6151
R1675 B.n914 B.n913 10.6151
R1676 B.n913 B.n912 10.6151
R1677 B.n912 B.n73 10.6151
R1678 B.n906 B.n73 10.6151
R1679 B.n906 B.n905 10.6151
R1680 B.n905 B.n904 10.6151
R1681 B.n904 B.n80 10.6151
R1682 B.n898 B.n80 10.6151
R1683 B.n898 B.n897 10.6151
R1684 B.n897 B.n896 10.6151
R1685 B.n896 B.n87 10.6151
R1686 B.n890 B.n87 10.6151
R1687 B.n890 B.n889 10.6151
R1688 B.n889 B.n888 10.6151
R1689 B.n229 B.n228 6.5566
R1690 B.n245 B.n145 6.5566
R1691 B.n560 B.n457 6.5566
R1692 B.n577 B.n576 6.5566
R1693 B.t14 B.n407 4.56076
R1694 B.t7 B.n78 4.56076
R1695 B.n228 B.n227 4.05904
R1696 B.n248 B.n145 4.05904
R1697 B.n458 B.n457 4.05904
R1698 B.n578 B.n577 4.05904
R1699 B.t3 B.n336 3.25783
R1700 B.t0 B.n15 3.25783
R1701 B.n992 B.n0 2.81026
R1702 B.n992 B.n1 2.81026
R1703 B.n383 B.t5 1.9549
R1704 B.t2 B.n933 1.9549
R1705 B.n764 B.t1 0.651966
R1706 B.n956 B.t4 0.651966
R1707 VP.n16 VP.n15 161.3
R1708 VP.n17 VP.n12 161.3
R1709 VP.n19 VP.n18 161.3
R1710 VP.n20 VP.n11 161.3
R1711 VP.n22 VP.n21 161.3
R1712 VP.n23 VP.n10 161.3
R1713 VP.n25 VP.n24 161.3
R1714 VP.n50 VP.n49 161.3
R1715 VP.n48 VP.n1 161.3
R1716 VP.n47 VP.n46 161.3
R1717 VP.n45 VP.n2 161.3
R1718 VP.n44 VP.n43 161.3
R1719 VP.n42 VP.n3 161.3
R1720 VP.n41 VP.n40 161.3
R1721 VP.n39 VP.n4 161.3
R1722 VP.n38 VP.n37 161.3
R1723 VP.n36 VP.n5 161.3
R1724 VP.n35 VP.n34 161.3
R1725 VP.n33 VP.n6 161.3
R1726 VP.n32 VP.n31 161.3
R1727 VP.n30 VP.n7 161.3
R1728 VP.n29 VP.n28 161.3
R1729 VP.n14 VP.t3 116.094
R1730 VP.n4 VP.t1 82.5377
R1731 VP.n8 VP.t2 82.5377
R1732 VP.n0 VP.t5 82.5377
R1733 VP.n13 VP.t0 82.5377
R1734 VP.n9 VP.t4 82.5377
R1735 VP.n27 VP.n8 79.3019
R1736 VP.n51 VP.n0 79.3019
R1737 VP.n26 VP.n9 79.3019
R1738 VP.n35 VP.n6 54.0911
R1739 VP.n43 VP.n2 54.0911
R1740 VP.n18 VP.n11 54.0911
R1741 VP.n27 VP.n26 51.5524
R1742 VP.n14 VP.n13 50.1285
R1743 VP.n31 VP.n6 26.8957
R1744 VP.n47 VP.n2 26.8957
R1745 VP.n22 VP.n11 26.8957
R1746 VP.n30 VP.n29 24.4675
R1747 VP.n31 VP.n30 24.4675
R1748 VP.n36 VP.n35 24.4675
R1749 VP.n37 VP.n36 24.4675
R1750 VP.n37 VP.n4 24.4675
R1751 VP.n41 VP.n4 24.4675
R1752 VP.n42 VP.n41 24.4675
R1753 VP.n43 VP.n42 24.4675
R1754 VP.n48 VP.n47 24.4675
R1755 VP.n49 VP.n48 24.4675
R1756 VP.n23 VP.n22 24.4675
R1757 VP.n24 VP.n23 24.4675
R1758 VP.n16 VP.n13 24.4675
R1759 VP.n17 VP.n16 24.4675
R1760 VP.n18 VP.n17 24.4675
R1761 VP.n29 VP.n8 10.766
R1762 VP.n49 VP.n0 10.766
R1763 VP.n24 VP.n9 10.766
R1764 VP.n15 VP.n14 3.1271
R1765 VP.n26 VP.n25 0.354971
R1766 VP.n28 VP.n27 0.354971
R1767 VP.n51 VP.n50 0.354971
R1768 VP VP.n51 0.26696
R1769 VP.n15 VP.n12 0.189894
R1770 VP.n19 VP.n12 0.189894
R1771 VP.n20 VP.n19 0.189894
R1772 VP.n21 VP.n20 0.189894
R1773 VP.n21 VP.n10 0.189894
R1774 VP.n25 VP.n10 0.189894
R1775 VP.n28 VP.n7 0.189894
R1776 VP.n32 VP.n7 0.189894
R1777 VP.n33 VP.n32 0.189894
R1778 VP.n34 VP.n33 0.189894
R1779 VP.n34 VP.n5 0.189894
R1780 VP.n38 VP.n5 0.189894
R1781 VP.n39 VP.n38 0.189894
R1782 VP.n40 VP.n39 0.189894
R1783 VP.n40 VP.n3 0.189894
R1784 VP.n44 VP.n3 0.189894
R1785 VP.n45 VP.n44 0.189894
R1786 VP.n46 VP.n45 0.189894
R1787 VP.n46 VP.n1 0.189894
R1788 VP.n50 VP.n1 0.189894
R1789 VDD1 VDD1.t4 69.5726
R1790 VDD1.n1 VDD1.t5 69.4581
R1791 VDD1.n1 VDD1.n0 66.1492
R1792 VDD1.n3 VDD1.n2 65.4026
R1793 VDD1.n3 VDD1.n1 46.3328
R1794 VDD1.n2 VDD1.t3 1.70593
R1795 VDD1.n2 VDD1.t1 1.70593
R1796 VDD1.n0 VDD1.t2 1.70593
R1797 VDD1.n0 VDD1.t0 1.70593
R1798 VDD1 VDD1.n3 0.744035
R1799 VTAIL.n7 VTAIL.t4 50.4304
R1800 VTAIL.n11 VTAIL.t1 50.4294
R1801 VTAIL.n2 VTAIL.t6 50.4294
R1802 VTAIL.n10 VTAIL.t7 50.4293
R1803 VTAIL.n9 VTAIL.n8 48.725
R1804 VTAIL.n6 VTAIL.n5 48.725
R1805 VTAIL.n1 VTAIL.n0 48.724
R1806 VTAIL.n4 VTAIL.n3 48.724
R1807 VTAIL.n6 VTAIL.n4 28.7893
R1808 VTAIL.n11 VTAIL.n10 25.5824
R1809 VTAIL.n7 VTAIL.n6 3.2074
R1810 VTAIL.n10 VTAIL.n9 3.2074
R1811 VTAIL.n4 VTAIL.n2 3.2074
R1812 VTAIL VTAIL.n11 2.34748
R1813 VTAIL.n9 VTAIL.n7 2.07378
R1814 VTAIL.n2 VTAIL.n1 2.07378
R1815 VTAIL.n0 VTAIL.t0 1.70593
R1816 VTAIL.n0 VTAIL.t2 1.70593
R1817 VTAIL.n3 VTAIL.t9 1.70593
R1818 VTAIL.n3 VTAIL.t10 1.70593
R1819 VTAIL.n8 VTAIL.t8 1.70593
R1820 VTAIL.n8 VTAIL.t11 1.70593
R1821 VTAIL.n5 VTAIL.t5 1.70593
R1822 VTAIL.n5 VTAIL.t3 1.70593
R1823 VTAIL VTAIL.n1 0.860414
R1824 VN.n34 VN.n33 161.3
R1825 VN.n32 VN.n19 161.3
R1826 VN.n31 VN.n30 161.3
R1827 VN.n29 VN.n20 161.3
R1828 VN.n28 VN.n27 161.3
R1829 VN.n26 VN.n21 161.3
R1830 VN.n25 VN.n24 161.3
R1831 VN.n16 VN.n15 161.3
R1832 VN.n14 VN.n1 161.3
R1833 VN.n13 VN.n12 161.3
R1834 VN.n11 VN.n2 161.3
R1835 VN.n10 VN.n9 161.3
R1836 VN.n8 VN.n3 161.3
R1837 VN.n7 VN.n6 161.3
R1838 VN.n23 VN.t3 116.094
R1839 VN.n5 VN.t5 116.094
R1840 VN.n4 VN.t4 82.5377
R1841 VN.n0 VN.t2 82.5377
R1842 VN.n22 VN.t1 82.5377
R1843 VN.n18 VN.t0 82.5377
R1844 VN.n17 VN.n0 79.3019
R1845 VN.n35 VN.n18 79.3019
R1846 VN.n9 VN.n2 54.0911
R1847 VN.n27 VN.n20 54.0911
R1848 VN VN.n35 51.7177
R1849 VN.n23 VN.n22 50.1285
R1850 VN.n5 VN.n4 50.1285
R1851 VN.n13 VN.n2 26.8957
R1852 VN.n31 VN.n20 26.8957
R1853 VN.n7 VN.n4 24.4675
R1854 VN.n8 VN.n7 24.4675
R1855 VN.n9 VN.n8 24.4675
R1856 VN.n14 VN.n13 24.4675
R1857 VN.n15 VN.n14 24.4675
R1858 VN.n27 VN.n26 24.4675
R1859 VN.n26 VN.n25 24.4675
R1860 VN.n25 VN.n22 24.4675
R1861 VN.n33 VN.n32 24.4675
R1862 VN.n32 VN.n31 24.4675
R1863 VN.n15 VN.n0 10.766
R1864 VN.n33 VN.n18 10.766
R1865 VN.n24 VN.n23 3.12711
R1866 VN.n6 VN.n5 3.12711
R1867 VN.n35 VN.n34 0.354971
R1868 VN.n17 VN.n16 0.354971
R1869 VN VN.n17 0.26696
R1870 VN.n34 VN.n19 0.189894
R1871 VN.n30 VN.n19 0.189894
R1872 VN.n30 VN.n29 0.189894
R1873 VN.n29 VN.n28 0.189894
R1874 VN.n28 VN.n21 0.189894
R1875 VN.n24 VN.n21 0.189894
R1876 VN.n6 VN.n3 0.189894
R1877 VN.n10 VN.n3 0.189894
R1878 VN.n11 VN.n10 0.189894
R1879 VN.n12 VN.n11 0.189894
R1880 VN.n12 VN.n1 0.189894
R1881 VN.n16 VN.n1 0.189894
R1882 VDD2.n1 VDD2.t0 69.4581
R1883 VDD2.n2 VDD2.t5 67.1092
R1884 VDD2.n1 VDD2.n0 66.1492
R1885 VDD2 VDD2.n3 66.1462
R1886 VDD2.n2 VDD2.n1 44.1463
R1887 VDD2 VDD2.n2 2.46386
R1888 VDD2.n3 VDD2.t4 1.70593
R1889 VDD2.n3 VDD2.t2 1.70593
R1890 VDD2.n0 VDD2.t1 1.70593
R1891 VDD2.n0 VDD2.t3 1.70593
C0 VP VDD2 0.525324f
C1 VDD1 VTAIL 7.84524f
C2 VP VDD1 7.18572f
C3 VDD2 VN 6.81526f
C4 VP VTAIL 7.19703f
C5 VDD1 VN 0.151859f
C6 VN VTAIL 7.1828f
C7 VDD1 VDD2 1.71541f
C8 VP VN 7.62445f
C9 VDD2 VTAIL 7.90214f
C10 VDD2 B 6.509892f
C11 VDD1 B 6.870287f
C12 VTAIL B 8.166581f
C13 VN B 15.179161f
C14 VP B 13.88411f
C15 VDD2.t0 B 2.24485f
C16 VDD2.t1 B 0.19584f
C17 VDD2.t3 B 0.19584f
C18 VDD2.n0 B 1.75567f
C19 VDD2.n1 B 2.73243f
C20 VDD2.t5 B 2.23163f
C21 VDD2.n2 B 2.53342f
C22 VDD2.t4 B 0.19584f
C23 VDD2.t2 B 0.19584f
C24 VDD2.n3 B 1.75563f
C25 VN.t2 B 2.11178f
C26 VN.n0 B 0.817597f
C27 VN.n1 B 0.019712f
C28 VN.n2 B 0.021528f
C29 VN.n3 B 0.019712f
C30 VN.t4 B 2.11178f
C31 VN.n4 B 0.820635f
C32 VN.t5 B 2.36855f
C33 VN.n5 B 0.77212f
C34 VN.n6 B 0.240663f
C35 VN.n7 B 0.036738f
C36 VN.n8 B 0.036738f
C37 VN.n9 B 0.034551f
C38 VN.n10 B 0.019712f
C39 VN.n11 B 0.019712f
C40 VN.n12 B 0.019712f
C41 VN.n13 B 0.038211f
C42 VN.n14 B 0.036738f
C43 VN.n15 B 0.026581f
C44 VN.n16 B 0.031815f
C45 VN.n17 B 0.051389f
C46 VN.t0 B 2.11178f
C47 VN.n18 B 0.817597f
C48 VN.n19 B 0.019712f
C49 VN.n20 B 0.021528f
C50 VN.n21 B 0.019712f
C51 VN.t1 B 2.11178f
C52 VN.n22 B 0.820635f
C53 VN.t3 B 2.36855f
C54 VN.n23 B 0.77212f
C55 VN.n24 B 0.240663f
C56 VN.n25 B 0.036738f
C57 VN.n26 B 0.036738f
C58 VN.n27 B 0.034551f
C59 VN.n28 B 0.019712f
C60 VN.n29 B 0.019712f
C61 VN.n30 B 0.019712f
C62 VN.n31 B 0.038211f
C63 VN.n32 B 0.036738f
C64 VN.n33 B 0.026581f
C65 VN.n34 B 0.031815f
C66 VN.n35 B 1.18266f
C67 VTAIL.t0 B 0.223414f
C68 VTAIL.t2 B 0.223414f
C69 VTAIL.n0 B 1.9334f
C70 VTAIL.n1 B 0.451434f
C71 VTAIL.t6 B 2.46427f
C72 VTAIL.n2 B 0.714028f
C73 VTAIL.t9 B 0.223414f
C74 VTAIL.t10 B 0.223414f
C75 VTAIL.n3 B 1.9334f
C76 VTAIL.n4 B 2.09229f
C77 VTAIL.t5 B 0.223414f
C78 VTAIL.t3 B 0.223414f
C79 VTAIL.n5 B 1.93339f
C80 VTAIL.n6 B 2.0923f
C81 VTAIL.t4 B 2.46427f
C82 VTAIL.n7 B 0.71403f
C83 VTAIL.t8 B 0.223414f
C84 VTAIL.t11 B 0.223414f
C85 VTAIL.n8 B 1.93339f
C86 VTAIL.n9 B 0.635598f
C87 VTAIL.t7 B 2.46426f
C88 VTAIL.n10 B 1.91911f
C89 VTAIL.t1 B 2.46427f
C90 VTAIL.n11 B 1.85162f
C91 VDD1.t4 B 2.27934f
C92 VDD1.t5 B 2.27844f
C93 VDD1.t2 B 0.198771f
C94 VDD1.t0 B 0.198771f
C95 VDD1.n0 B 1.78194f
C96 VDD1.n1 B 2.89872f
C97 VDD1.t3 B 0.198771f
C98 VDD1.t1 B 0.198771f
C99 VDD1.n2 B 1.7768f
C100 VDD1.n3 B 2.57589f
C101 VP.t5 B 2.15365f
C102 VP.n0 B 0.833807f
C103 VP.n1 B 0.020103f
C104 VP.n2 B 0.021955f
C105 VP.n3 B 0.020103f
C106 VP.t1 B 2.15365f
C107 VP.n4 B 0.776571f
C108 VP.n5 B 0.020103f
C109 VP.n6 B 0.021955f
C110 VP.n7 B 0.020103f
C111 VP.t2 B 2.15365f
C112 VP.n8 B 0.833807f
C113 VP.t4 B 2.15365f
C114 VP.n9 B 0.833807f
C115 VP.n10 B 0.020103f
C116 VP.n11 B 0.021955f
C117 VP.n12 B 0.020103f
C118 VP.t0 B 2.15365f
C119 VP.n13 B 0.836906f
C120 VP.t3 B 2.41551f
C121 VP.n14 B 0.78743f
C122 VP.n15 B 0.245435f
C123 VP.n16 B 0.037466f
C124 VP.n17 B 0.037466f
C125 VP.n18 B 0.035236f
C126 VP.n19 B 0.020103f
C127 VP.n20 B 0.020103f
C128 VP.n21 B 0.020103f
C129 VP.n22 B 0.038968f
C130 VP.n23 B 0.037466f
C131 VP.n24 B 0.027108f
C132 VP.n25 B 0.032445f
C133 VP.n26 B 1.19797f
C134 VP.n27 B 1.21198f
C135 VP.n28 B 0.032445f
C136 VP.n29 B 0.027108f
C137 VP.n30 B 0.037466f
C138 VP.n31 B 0.038968f
C139 VP.n32 B 0.020103f
C140 VP.n33 B 0.020103f
C141 VP.n34 B 0.020103f
C142 VP.n35 B 0.035236f
C143 VP.n36 B 0.037466f
C144 VP.n37 B 0.037466f
C145 VP.n38 B 0.020103f
C146 VP.n39 B 0.020103f
C147 VP.n40 B 0.020103f
C148 VP.n41 B 0.037466f
C149 VP.n42 B 0.037466f
C150 VP.n43 B 0.035236f
C151 VP.n44 B 0.020103f
C152 VP.n45 B 0.020103f
C153 VP.n46 B 0.020103f
C154 VP.n47 B 0.038968f
C155 VP.n48 B 0.037466f
C156 VP.n49 B 0.027108f
C157 VP.n50 B 0.032445f
C158 VP.n51 B 0.052408f
.ends

