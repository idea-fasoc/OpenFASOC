* NGSPICE file created from diff_pair_sample_1203.ext - technology: sky130A

.subckt diff_pair_sample_1203 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t5 VN.t0 VTAIL.t7 w_n1418_n3168# sky130_fd_pr__pfet_01v8 ad=4.29 pd=22.78 as=1.815 ps=11.33 w=11 l=0.23
X1 B.t11 B.t9 B.t10 w_n1418_n3168# sky130_fd_pr__pfet_01v8 ad=4.29 pd=22.78 as=0 ps=0 w=11 l=0.23
X2 VDD2.t4 VN.t1 VTAIL.t8 w_n1418_n3168# sky130_fd_pr__pfet_01v8 ad=1.815 pd=11.33 as=4.29 ps=22.78 w=11 l=0.23
X3 VTAIL.t3 VP.t0 VDD1.t5 w_n1418_n3168# sky130_fd_pr__pfet_01v8 ad=1.815 pd=11.33 as=1.815 ps=11.33 w=11 l=0.23
X4 VDD1.t4 VP.t1 VTAIL.t1 w_n1418_n3168# sky130_fd_pr__pfet_01v8 ad=1.815 pd=11.33 as=4.29 ps=22.78 w=11 l=0.23
X5 VTAIL.t10 VN.t2 VDD2.t3 w_n1418_n3168# sky130_fd_pr__pfet_01v8 ad=1.815 pd=11.33 as=1.815 ps=11.33 w=11 l=0.23
X6 VDD1.t3 VP.t2 VTAIL.t2 w_n1418_n3168# sky130_fd_pr__pfet_01v8 ad=1.815 pd=11.33 as=4.29 ps=22.78 w=11 l=0.23
X7 VDD1.t2 VP.t3 VTAIL.t0 w_n1418_n3168# sky130_fd_pr__pfet_01v8 ad=4.29 pd=22.78 as=1.815 ps=11.33 w=11 l=0.23
X8 B.t8 B.t6 B.t7 w_n1418_n3168# sky130_fd_pr__pfet_01v8 ad=4.29 pd=22.78 as=0 ps=0 w=11 l=0.23
X9 VTAIL.t5 VP.t4 VDD1.t1 w_n1418_n3168# sky130_fd_pr__pfet_01v8 ad=1.815 pd=11.33 as=1.815 ps=11.33 w=11 l=0.23
X10 VDD2.t2 VN.t3 VTAIL.t11 w_n1418_n3168# sky130_fd_pr__pfet_01v8 ad=1.815 pd=11.33 as=4.29 ps=22.78 w=11 l=0.23
X11 VDD1.t0 VP.t5 VTAIL.t4 w_n1418_n3168# sky130_fd_pr__pfet_01v8 ad=4.29 pd=22.78 as=1.815 ps=11.33 w=11 l=0.23
X12 B.t5 B.t3 B.t4 w_n1418_n3168# sky130_fd_pr__pfet_01v8 ad=4.29 pd=22.78 as=0 ps=0 w=11 l=0.23
X13 B.t2 B.t0 B.t1 w_n1418_n3168# sky130_fd_pr__pfet_01v8 ad=4.29 pd=22.78 as=0 ps=0 w=11 l=0.23
X14 VDD2.t1 VN.t4 VTAIL.t6 w_n1418_n3168# sky130_fd_pr__pfet_01v8 ad=4.29 pd=22.78 as=1.815 ps=11.33 w=11 l=0.23
X15 VTAIL.t9 VN.t5 VDD2.t0 w_n1418_n3168# sky130_fd_pr__pfet_01v8 ad=1.815 pd=11.33 as=1.815 ps=11.33 w=11 l=0.23
R0 VN.n2 VN.t1 1334.1
R1 VN.n0 VN.t4 1334.1
R2 VN.n6 VN.t0 1334.1
R3 VN.n4 VN.t3 1334.1
R4 VN.n1 VN.t5 1288.83
R5 VN.n5 VN.t2 1288.83
R6 VN.n7 VN.n4 161.489
R7 VN.n3 VN.n0 161.489
R8 VN.n3 VN.n2 161.3
R9 VN.n7 VN.n6 161.3
R10 VN VN.n7 39.0782
R11 VN.n1 VN.n0 36.5157
R12 VN.n2 VN.n1 36.5157
R13 VN.n6 VN.n5 36.5157
R14 VN.n5 VN.n4 36.5157
R15 VN VN.n3 0.0516364
R16 VTAIL.n7 VTAIL.t11 60.8054
R17 VTAIL.n11 VTAIL.t8 60.8053
R18 VTAIL.n2 VTAIL.t2 60.8053
R19 VTAIL.n10 VTAIL.t1 60.8053
R20 VTAIL.n9 VTAIL.n8 57.8505
R21 VTAIL.n6 VTAIL.n5 57.8505
R22 VTAIL.n1 VTAIL.n0 57.8503
R23 VTAIL.n4 VTAIL.n3 57.8503
R24 VTAIL.n6 VTAIL.n4 22.8152
R25 VTAIL.n11 VTAIL.n10 22.3324
R26 VTAIL.n0 VTAIL.t6 2.9555
R27 VTAIL.n0 VTAIL.t9 2.9555
R28 VTAIL.n3 VTAIL.t4 2.9555
R29 VTAIL.n3 VTAIL.t5 2.9555
R30 VTAIL.n8 VTAIL.t0 2.9555
R31 VTAIL.n8 VTAIL.t3 2.9555
R32 VTAIL.n5 VTAIL.t7 2.9555
R33 VTAIL.n5 VTAIL.t10 2.9555
R34 VTAIL.n9 VTAIL.n7 0.711707
R35 VTAIL.n2 VTAIL.n1 0.711707
R36 VTAIL.n7 VTAIL.n6 0.483259
R37 VTAIL.n10 VTAIL.n9 0.483259
R38 VTAIL.n4 VTAIL.n2 0.483259
R39 VTAIL VTAIL.n11 0.304379
R40 VTAIL VTAIL.n1 0.179379
R41 VDD2.n1 VDD2.t1 77.7908
R42 VDD2.n2 VDD2.t5 77.4842
R43 VDD2.n1 VDD2.n0 74.5944
R44 VDD2 VDD2.n3 74.5916
R45 VDD2.n2 VDD2.n1 34.767
R46 VDD2.n3 VDD2.t3 2.9555
R47 VDD2.n3 VDD2.t2 2.9555
R48 VDD2.n0 VDD2.t0 2.9555
R49 VDD2.n0 VDD2.t4 2.9555
R50 VDD2 VDD2.n2 0.420759
R51 B.n99 B.t0 1381.1
R52 B.n93 B.t9 1381.1
R53 B.n37 B.t3 1381.1
R54 B.n30 B.t6 1381.1
R55 B.n278 B.n277 585
R56 B.n276 B.n73 585
R57 B.n275 B.n274 585
R58 B.n273 B.n74 585
R59 B.n272 B.n271 585
R60 B.n270 B.n75 585
R61 B.n269 B.n268 585
R62 B.n267 B.n76 585
R63 B.n266 B.n265 585
R64 B.n264 B.n77 585
R65 B.n263 B.n262 585
R66 B.n261 B.n78 585
R67 B.n260 B.n259 585
R68 B.n258 B.n79 585
R69 B.n257 B.n256 585
R70 B.n255 B.n80 585
R71 B.n254 B.n253 585
R72 B.n252 B.n81 585
R73 B.n251 B.n250 585
R74 B.n249 B.n82 585
R75 B.n248 B.n247 585
R76 B.n246 B.n83 585
R77 B.n245 B.n244 585
R78 B.n243 B.n84 585
R79 B.n242 B.n241 585
R80 B.n240 B.n85 585
R81 B.n239 B.n238 585
R82 B.n237 B.n86 585
R83 B.n236 B.n235 585
R84 B.n234 B.n87 585
R85 B.n233 B.n232 585
R86 B.n231 B.n88 585
R87 B.n230 B.n229 585
R88 B.n228 B.n89 585
R89 B.n227 B.n226 585
R90 B.n225 B.n90 585
R91 B.n224 B.n223 585
R92 B.n222 B.n91 585
R93 B.n221 B.n220 585
R94 B.n218 B.n92 585
R95 B.n217 B.n216 585
R96 B.n215 B.n95 585
R97 B.n214 B.n213 585
R98 B.n212 B.n96 585
R99 B.n211 B.n210 585
R100 B.n209 B.n97 585
R101 B.n208 B.n207 585
R102 B.n206 B.n98 585
R103 B.n204 B.n203 585
R104 B.n202 B.n101 585
R105 B.n201 B.n200 585
R106 B.n199 B.n102 585
R107 B.n198 B.n197 585
R108 B.n196 B.n103 585
R109 B.n195 B.n194 585
R110 B.n193 B.n104 585
R111 B.n192 B.n191 585
R112 B.n190 B.n105 585
R113 B.n189 B.n188 585
R114 B.n187 B.n106 585
R115 B.n186 B.n185 585
R116 B.n184 B.n107 585
R117 B.n183 B.n182 585
R118 B.n181 B.n108 585
R119 B.n180 B.n179 585
R120 B.n178 B.n109 585
R121 B.n177 B.n176 585
R122 B.n175 B.n110 585
R123 B.n174 B.n173 585
R124 B.n172 B.n111 585
R125 B.n171 B.n170 585
R126 B.n169 B.n112 585
R127 B.n168 B.n167 585
R128 B.n166 B.n113 585
R129 B.n165 B.n164 585
R130 B.n163 B.n114 585
R131 B.n162 B.n161 585
R132 B.n160 B.n115 585
R133 B.n159 B.n158 585
R134 B.n157 B.n116 585
R135 B.n156 B.n155 585
R136 B.n154 B.n117 585
R137 B.n153 B.n152 585
R138 B.n151 B.n118 585
R139 B.n150 B.n149 585
R140 B.n148 B.n119 585
R141 B.n147 B.n146 585
R142 B.n279 B.n72 585
R143 B.n281 B.n280 585
R144 B.n282 B.n71 585
R145 B.n284 B.n283 585
R146 B.n285 B.n70 585
R147 B.n287 B.n286 585
R148 B.n288 B.n69 585
R149 B.n290 B.n289 585
R150 B.n291 B.n68 585
R151 B.n293 B.n292 585
R152 B.n294 B.n67 585
R153 B.n296 B.n295 585
R154 B.n297 B.n66 585
R155 B.n299 B.n298 585
R156 B.n300 B.n65 585
R157 B.n302 B.n301 585
R158 B.n303 B.n64 585
R159 B.n305 B.n304 585
R160 B.n306 B.n63 585
R161 B.n308 B.n307 585
R162 B.n309 B.n62 585
R163 B.n311 B.n310 585
R164 B.n312 B.n61 585
R165 B.n314 B.n313 585
R166 B.n315 B.n60 585
R167 B.n317 B.n316 585
R168 B.n318 B.n59 585
R169 B.n320 B.n319 585
R170 B.n321 B.n58 585
R171 B.n323 B.n322 585
R172 B.n454 B.n9 585
R173 B.n453 B.n452 585
R174 B.n451 B.n10 585
R175 B.n450 B.n449 585
R176 B.n448 B.n11 585
R177 B.n447 B.n446 585
R178 B.n445 B.n12 585
R179 B.n444 B.n443 585
R180 B.n442 B.n13 585
R181 B.n441 B.n440 585
R182 B.n439 B.n14 585
R183 B.n438 B.n437 585
R184 B.n436 B.n15 585
R185 B.n435 B.n434 585
R186 B.n433 B.n16 585
R187 B.n432 B.n431 585
R188 B.n430 B.n17 585
R189 B.n429 B.n428 585
R190 B.n427 B.n18 585
R191 B.n426 B.n425 585
R192 B.n424 B.n19 585
R193 B.n423 B.n422 585
R194 B.n421 B.n20 585
R195 B.n420 B.n419 585
R196 B.n418 B.n21 585
R197 B.n417 B.n416 585
R198 B.n415 B.n22 585
R199 B.n414 B.n413 585
R200 B.n412 B.n23 585
R201 B.n411 B.n410 585
R202 B.n409 B.n24 585
R203 B.n408 B.n407 585
R204 B.n406 B.n25 585
R205 B.n405 B.n404 585
R206 B.n403 B.n26 585
R207 B.n402 B.n401 585
R208 B.n400 B.n27 585
R209 B.n399 B.n398 585
R210 B.n397 B.n28 585
R211 B.n396 B.n395 585
R212 B.n394 B.n29 585
R213 B.n393 B.n392 585
R214 B.n391 B.n33 585
R215 B.n390 B.n389 585
R216 B.n388 B.n34 585
R217 B.n387 B.n386 585
R218 B.n385 B.n35 585
R219 B.n384 B.n383 585
R220 B.n381 B.n36 585
R221 B.n380 B.n379 585
R222 B.n378 B.n39 585
R223 B.n377 B.n376 585
R224 B.n375 B.n40 585
R225 B.n374 B.n373 585
R226 B.n372 B.n41 585
R227 B.n371 B.n370 585
R228 B.n369 B.n42 585
R229 B.n368 B.n367 585
R230 B.n366 B.n43 585
R231 B.n365 B.n364 585
R232 B.n363 B.n44 585
R233 B.n362 B.n361 585
R234 B.n360 B.n45 585
R235 B.n359 B.n358 585
R236 B.n357 B.n46 585
R237 B.n356 B.n355 585
R238 B.n354 B.n47 585
R239 B.n353 B.n352 585
R240 B.n351 B.n48 585
R241 B.n350 B.n349 585
R242 B.n348 B.n49 585
R243 B.n347 B.n346 585
R244 B.n345 B.n50 585
R245 B.n344 B.n343 585
R246 B.n342 B.n51 585
R247 B.n341 B.n340 585
R248 B.n339 B.n52 585
R249 B.n338 B.n337 585
R250 B.n336 B.n53 585
R251 B.n335 B.n334 585
R252 B.n333 B.n54 585
R253 B.n332 B.n331 585
R254 B.n330 B.n55 585
R255 B.n329 B.n328 585
R256 B.n327 B.n56 585
R257 B.n326 B.n325 585
R258 B.n324 B.n57 585
R259 B.n456 B.n455 585
R260 B.n457 B.n8 585
R261 B.n459 B.n458 585
R262 B.n460 B.n7 585
R263 B.n462 B.n461 585
R264 B.n463 B.n6 585
R265 B.n465 B.n464 585
R266 B.n466 B.n5 585
R267 B.n468 B.n467 585
R268 B.n469 B.n4 585
R269 B.n471 B.n470 585
R270 B.n472 B.n3 585
R271 B.n474 B.n473 585
R272 B.n475 B.n0 585
R273 B.n2 B.n1 585
R274 B.n127 B.n126 585
R275 B.n129 B.n128 585
R276 B.n130 B.n125 585
R277 B.n132 B.n131 585
R278 B.n133 B.n124 585
R279 B.n135 B.n134 585
R280 B.n136 B.n123 585
R281 B.n138 B.n137 585
R282 B.n139 B.n122 585
R283 B.n141 B.n140 585
R284 B.n142 B.n121 585
R285 B.n144 B.n143 585
R286 B.n145 B.n120 585
R287 B.n147 B.n120 526.135
R288 B.n277 B.n72 526.135
R289 B.n324 B.n323 526.135
R290 B.n456 B.n9 526.135
R291 B.n477 B.n476 256.663
R292 B.n476 B.n475 235.042
R293 B.n476 B.n2 235.042
R294 B.n148 B.n147 163.367
R295 B.n149 B.n148 163.367
R296 B.n149 B.n118 163.367
R297 B.n153 B.n118 163.367
R298 B.n154 B.n153 163.367
R299 B.n155 B.n154 163.367
R300 B.n155 B.n116 163.367
R301 B.n159 B.n116 163.367
R302 B.n160 B.n159 163.367
R303 B.n161 B.n160 163.367
R304 B.n161 B.n114 163.367
R305 B.n165 B.n114 163.367
R306 B.n166 B.n165 163.367
R307 B.n167 B.n166 163.367
R308 B.n167 B.n112 163.367
R309 B.n171 B.n112 163.367
R310 B.n172 B.n171 163.367
R311 B.n173 B.n172 163.367
R312 B.n173 B.n110 163.367
R313 B.n177 B.n110 163.367
R314 B.n178 B.n177 163.367
R315 B.n179 B.n178 163.367
R316 B.n179 B.n108 163.367
R317 B.n183 B.n108 163.367
R318 B.n184 B.n183 163.367
R319 B.n185 B.n184 163.367
R320 B.n185 B.n106 163.367
R321 B.n189 B.n106 163.367
R322 B.n190 B.n189 163.367
R323 B.n191 B.n190 163.367
R324 B.n191 B.n104 163.367
R325 B.n195 B.n104 163.367
R326 B.n196 B.n195 163.367
R327 B.n197 B.n196 163.367
R328 B.n197 B.n102 163.367
R329 B.n201 B.n102 163.367
R330 B.n202 B.n201 163.367
R331 B.n203 B.n202 163.367
R332 B.n203 B.n98 163.367
R333 B.n208 B.n98 163.367
R334 B.n209 B.n208 163.367
R335 B.n210 B.n209 163.367
R336 B.n210 B.n96 163.367
R337 B.n214 B.n96 163.367
R338 B.n215 B.n214 163.367
R339 B.n216 B.n215 163.367
R340 B.n216 B.n92 163.367
R341 B.n221 B.n92 163.367
R342 B.n222 B.n221 163.367
R343 B.n223 B.n222 163.367
R344 B.n223 B.n90 163.367
R345 B.n227 B.n90 163.367
R346 B.n228 B.n227 163.367
R347 B.n229 B.n228 163.367
R348 B.n229 B.n88 163.367
R349 B.n233 B.n88 163.367
R350 B.n234 B.n233 163.367
R351 B.n235 B.n234 163.367
R352 B.n235 B.n86 163.367
R353 B.n239 B.n86 163.367
R354 B.n240 B.n239 163.367
R355 B.n241 B.n240 163.367
R356 B.n241 B.n84 163.367
R357 B.n245 B.n84 163.367
R358 B.n246 B.n245 163.367
R359 B.n247 B.n246 163.367
R360 B.n247 B.n82 163.367
R361 B.n251 B.n82 163.367
R362 B.n252 B.n251 163.367
R363 B.n253 B.n252 163.367
R364 B.n253 B.n80 163.367
R365 B.n257 B.n80 163.367
R366 B.n258 B.n257 163.367
R367 B.n259 B.n258 163.367
R368 B.n259 B.n78 163.367
R369 B.n263 B.n78 163.367
R370 B.n264 B.n263 163.367
R371 B.n265 B.n264 163.367
R372 B.n265 B.n76 163.367
R373 B.n269 B.n76 163.367
R374 B.n270 B.n269 163.367
R375 B.n271 B.n270 163.367
R376 B.n271 B.n74 163.367
R377 B.n275 B.n74 163.367
R378 B.n276 B.n275 163.367
R379 B.n277 B.n276 163.367
R380 B.n323 B.n58 163.367
R381 B.n319 B.n58 163.367
R382 B.n319 B.n318 163.367
R383 B.n318 B.n317 163.367
R384 B.n317 B.n60 163.367
R385 B.n313 B.n60 163.367
R386 B.n313 B.n312 163.367
R387 B.n312 B.n311 163.367
R388 B.n311 B.n62 163.367
R389 B.n307 B.n62 163.367
R390 B.n307 B.n306 163.367
R391 B.n306 B.n305 163.367
R392 B.n305 B.n64 163.367
R393 B.n301 B.n64 163.367
R394 B.n301 B.n300 163.367
R395 B.n300 B.n299 163.367
R396 B.n299 B.n66 163.367
R397 B.n295 B.n66 163.367
R398 B.n295 B.n294 163.367
R399 B.n294 B.n293 163.367
R400 B.n293 B.n68 163.367
R401 B.n289 B.n68 163.367
R402 B.n289 B.n288 163.367
R403 B.n288 B.n287 163.367
R404 B.n287 B.n70 163.367
R405 B.n283 B.n70 163.367
R406 B.n283 B.n282 163.367
R407 B.n282 B.n281 163.367
R408 B.n281 B.n72 163.367
R409 B.n452 B.n9 163.367
R410 B.n452 B.n451 163.367
R411 B.n451 B.n450 163.367
R412 B.n450 B.n11 163.367
R413 B.n446 B.n11 163.367
R414 B.n446 B.n445 163.367
R415 B.n445 B.n444 163.367
R416 B.n444 B.n13 163.367
R417 B.n440 B.n13 163.367
R418 B.n440 B.n439 163.367
R419 B.n439 B.n438 163.367
R420 B.n438 B.n15 163.367
R421 B.n434 B.n15 163.367
R422 B.n434 B.n433 163.367
R423 B.n433 B.n432 163.367
R424 B.n432 B.n17 163.367
R425 B.n428 B.n17 163.367
R426 B.n428 B.n427 163.367
R427 B.n427 B.n426 163.367
R428 B.n426 B.n19 163.367
R429 B.n422 B.n19 163.367
R430 B.n422 B.n421 163.367
R431 B.n421 B.n420 163.367
R432 B.n420 B.n21 163.367
R433 B.n416 B.n21 163.367
R434 B.n416 B.n415 163.367
R435 B.n415 B.n414 163.367
R436 B.n414 B.n23 163.367
R437 B.n410 B.n23 163.367
R438 B.n410 B.n409 163.367
R439 B.n409 B.n408 163.367
R440 B.n408 B.n25 163.367
R441 B.n404 B.n25 163.367
R442 B.n404 B.n403 163.367
R443 B.n403 B.n402 163.367
R444 B.n402 B.n27 163.367
R445 B.n398 B.n27 163.367
R446 B.n398 B.n397 163.367
R447 B.n397 B.n396 163.367
R448 B.n396 B.n29 163.367
R449 B.n392 B.n29 163.367
R450 B.n392 B.n391 163.367
R451 B.n391 B.n390 163.367
R452 B.n390 B.n34 163.367
R453 B.n386 B.n34 163.367
R454 B.n386 B.n385 163.367
R455 B.n385 B.n384 163.367
R456 B.n384 B.n36 163.367
R457 B.n379 B.n36 163.367
R458 B.n379 B.n378 163.367
R459 B.n378 B.n377 163.367
R460 B.n377 B.n40 163.367
R461 B.n373 B.n40 163.367
R462 B.n373 B.n372 163.367
R463 B.n372 B.n371 163.367
R464 B.n371 B.n42 163.367
R465 B.n367 B.n42 163.367
R466 B.n367 B.n366 163.367
R467 B.n366 B.n365 163.367
R468 B.n365 B.n44 163.367
R469 B.n361 B.n44 163.367
R470 B.n361 B.n360 163.367
R471 B.n360 B.n359 163.367
R472 B.n359 B.n46 163.367
R473 B.n355 B.n46 163.367
R474 B.n355 B.n354 163.367
R475 B.n354 B.n353 163.367
R476 B.n353 B.n48 163.367
R477 B.n349 B.n48 163.367
R478 B.n349 B.n348 163.367
R479 B.n348 B.n347 163.367
R480 B.n347 B.n50 163.367
R481 B.n343 B.n50 163.367
R482 B.n343 B.n342 163.367
R483 B.n342 B.n341 163.367
R484 B.n341 B.n52 163.367
R485 B.n337 B.n52 163.367
R486 B.n337 B.n336 163.367
R487 B.n336 B.n335 163.367
R488 B.n335 B.n54 163.367
R489 B.n331 B.n54 163.367
R490 B.n331 B.n330 163.367
R491 B.n330 B.n329 163.367
R492 B.n329 B.n56 163.367
R493 B.n325 B.n56 163.367
R494 B.n325 B.n324 163.367
R495 B.n457 B.n456 163.367
R496 B.n458 B.n457 163.367
R497 B.n458 B.n7 163.367
R498 B.n462 B.n7 163.367
R499 B.n463 B.n462 163.367
R500 B.n464 B.n463 163.367
R501 B.n464 B.n5 163.367
R502 B.n468 B.n5 163.367
R503 B.n469 B.n468 163.367
R504 B.n470 B.n469 163.367
R505 B.n470 B.n3 163.367
R506 B.n474 B.n3 163.367
R507 B.n475 B.n474 163.367
R508 B.n126 B.n2 163.367
R509 B.n129 B.n126 163.367
R510 B.n130 B.n129 163.367
R511 B.n131 B.n130 163.367
R512 B.n131 B.n124 163.367
R513 B.n135 B.n124 163.367
R514 B.n136 B.n135 163.367
R515 B.n137 B.n136 163.367
R516 B.n137 B.n122 163.367
R517 B.n141 B.n122 163.367
R518 B.n142 B.n141 163.367
R519 B.n143 B.n142 163.367
R520 B.n143 B.n120 163.367
R521 B.n93 B.t10 120.546
R522 B.n37 B.t5 120.546
R523 B.n99 B.t1 120.534
R524 B.n30 B.t8 120.534
R525 B.n94 B.t11 109.686
R526 B.n38 B.t4 109.686
R527 B.n100 B.t2 109.674
R528 B.n31 B.t7 109.674
R529 B.n205 B.n100 59.5399
R530 B.n219 B.n94 59.5399
R531 B.n382 B.n38 59.5399
R532 B.n32 B.n31 59.5399
R533 B.n455 B.n454 34.1859
R534 B.n322 B.n57 34.1859
R535 B.n279 B.n278 34.1859
R536 B.n146 B.n145 34.1859
R537 B B.n477 18.0485
R538 B.n100 B.n99 10.8611
R539 B.n94 B.n93 10.8611
R540 B.n38 B.n37 10.8611
R541 B.n31 B.n30 10.8611
R542 B.n455 B.n8 10.6151
R543 B.n459 B.n8 10.6151
R544 B.n460 B.n459 10.6151
R545 B.n461 B.n460 10.6151
R546 B.n461 B.n6 10.6151
R547 B.n465 B.n6 10.6151
R548 B.n466 B.n465 10.6151
R549 B.n467 B.n466 10.6151
R550 B.n467 B.n4 10.6151
R551 B.n471 B.n4 10.6151
R552 B.n472 B.n471 10.6151
R553 B.n473 B.n472 10.6151
R554 B.n473 B.n0 10.6151
R555 B.n454 B.n453 10.6151
R556 B.n453 B.n10 10.6151
R557 B.n449 B.n10 10.6151
R558 B.n449 B.n448 10.6151
R559 B.n448 B.n447 10.6151
R560 B.n447 B.n12 10.6151
R561 B.n443 B.n12 10.6151
R562 B.n443 B.n442 10.6151
R563 B.n442 B.n441 10.6151
R564 B.n441 B.n14 10.6151
R565 B.n437 B.n14 10.6151
R566 B.n437 B.n436 10.6151
R567 B.n436 B.n435 10.6151
R568 B.n435 B.n16 10.6151
R569 B.n431 B.n16 10.6151
R570 B.n431 B.n430 10.6151
R571 B.n430 B.n429 10.6151
R572 B.n429 B.n18 10.6151
R573 B.n425 B.n18 10.6151
R574 B.n425 B.n424 10.6151
R575 B.n424 B.n423 10.6151
R576 B.n423 B.n20 10.6151
R577 B.n419 B.n20 10.6151
R578 B.n419 B.n418 10.6151
R579 B.n418 B.n417 10.6151
R580 B.n417 B.n22 10.6151
R581 B.n413 B.n22 10.6151
R582 B.n413 B.n412 10.6151
R583 B.n412 B.n411 10.6151
R584 B.n411 B.n24 10.6151
R585 B.n407 B.n24 10.6151
R586 B.n407 B.n406 10.6151
R587 B.n406 B.n405 10.6151
R588 B.n405 B.n26 10.6151
R589 B.n401 B.n26 10.6151
R590 B.n401 B.n400 10.6151
R591 B.n400 B.n399 10.6151
R592 B.n399 B.n28 10.6151
R593 B.n395 B.n394 10.6151
R594 B.n394 B.n393 10.6151
R595 B.n393 B.n33 10.6151
R596 B.n389 B.n33 10.6151
R597 B.n389 B.n388 10.6151
R598 B.n388 B.n387 10.6151
R599 B.n387 B.n35 10.6151
R600 B.n383 B.n35 10.6151
R601 B.n381 B.n380 10.6151
R602 B.n380 B.n39 10.6151
R603 B.n376 B.n39 10.6151
R604 B.n376 B.n375 10.6151
R605 B.n375 B.n374 10.6151
R606 B.n374 B.n41 10.6151
R607 B.n370 B.n41 10.6151
R608 B.n370 B.n369 10.6151
R609 B.n369 B.n368 10.6151
R610 B.n368 B.n43 10.6151
R611 B.n364 B.n43 10.6151
R612 B.n364 B.n363 10.6151
R613 B.n363 B.n362 10.6151
R614 B.n362 B.n45 10.6151
R615 B.n358 B.n45 10.6151
R616 B.n358 B.n357 10.6151
R617 B.n357 B.n356 10.6151
R618 B.n356 B.n47 10.6151
R619 B.n352 B.n47 10.6151
R620 B.n352 B.n351 10.6151
R621 B.n351 B.n350 10.6151
R622 B.n350 B.n49 10.6151
R623 B.n346 B.n49 10.6151
R624 B.n346 B.n345 10.6151
R625 B.n345 B.n344 10.6151
R626 B.n344 B.n51 10.6151
R627 B.n340 B.n51 10.6151
R628 B.n340 B.n339 10.6151
R629 B.n339 B.n338 10.6151
R630 B.n338 B.n53 10.6151
R631 B.n334 B.n53 10.6151
R632 B.n334 B.n333 10.6151
R633 B.n333 B.n332 10.6151
R634 B.n332 B.n55 10.6151
R635 B.n328 B.n55 10.6151
R636 B.n328 B.n327 10.6151
R637 B.n327 B.n326 10.6151
R638 B.n326 B.n57 10.6151
R639 B.n322 B.n321 10.6151
R640 B.n321 B.n320 10.6151
R641 B.n320 B.n59 10.6151
R642 B.n316 B.n59 10.6151
R643 B.n316 B.n315 10.6151
R644 B.n315 B.n314 10.6151
R645 B.n314 B.n61 10.6151
R646 B.n310 B.n61 10.6151
R647 B.n310 B.n309 10.6151
R648 B.n309 B.n308 10.6151
R649 B.n308 B.n63 10.6151
R650 B.n304 B.n63 10.6151
R651 B.n304 B.n303 10.6151
R652 B.n303 B.n302 10.6151
R653 B.n302 B.n65 10.6151
R654 B.n298 B.n65 10.6151
R655 B.n298 B.n297 10.6151
R656 B.n297 B.n296 10.6151
R657 B.n296 B.n67 10.6151
R658 B.n292 B.n67 10.6151
R659 B.n292 B.n291 10.6151
R660 B.n291 B.n290 10.6151
R661 B.n290 B.n69 10.6151
R662 B.n286 B.n69 10.6151
R663 B.n286 B.n285 10.6151
R664 B.n285 B.n284 10.6151
R665 B.n284 B.n71 10.6151
R666 B.n280 B.n71 10.6151
R667 B.n280 B.n279 10.6151
R668 B.n127 B.n1 10.6151
R669 B.n128 B.n127 10.6151
R670 B.n128 B.n125 10.6151
R671 B.n132 B.n125 10.6151
R672 B.n133 B.n132 10.6151
R673 B.n134 B.n133 10.6151
R674 B.n134 B.n123 10.6151
R675 B.n138 B.n123 10.6151
R676 B.n139 B.n138 10.6151
R677 B.n140 B.n139 10.6151
R678 B.n140 B.n121 10.6151
R679 B.n144 B.n121 10.6151
R680 B.n145 B.n144 10.6151
R681 B.n146 B.n119 10.6151
R682 B.n150 B.n119 10.6151
R683 B.n151 B.n150 10.6151
R684 B.n152 B.n151 10.6151
R685 B.n152 B.n117 10.6151
R686 B.n156 B.n117 10.6151
R687 B.n157 B.n156 10.6151
R688 B.n158 B.n157 10.6151
R689 B.n158 B.n115 10.6151
R690 B.n162 B.n115 10.6151
R691 B.n163 B.n162 10.6151
R692 B.n164 B.n163 10.6151
R693 B.n164 B.n113 10.6151
R694 B.n168 B.n113 10.6151
R695 B.n169 B.n168 10.6151
R696 B.n170 B.n169 10.6151
R697 B.n170 B.n111 10.6151
R698 B.n174 B.n111 10.6151
R699 B.n175 B.n174 10.6151
R700 B.n176 B.n175 10.6151
R701 B.n176 B.n109 10.6151
R702 B.n180 B.n109 10.6151
R703 B.n181 B.n180 10.6151
R704 B.n182 B.n181 10.6151
R705 B.n182 B.n107 10.6151
R706 B.n186 B.n107 10.6151
R707 B.n187 B.n186 10.6151
R708 B.n188 B.n187 10.6151
R709 B.n188 B.n105 10.6151
R710 B.n192 B.n105 10.6151
R711 B.n193 B.n192 10.6151
R712 B.n194 B.n193 10.6151
R713 B.n194 B.n103 10.6151
R714 B.n198 B.n103 10.6151
R715 B.n199 B.n198 10.6151
R716 B.n200 B.n199 10.6151
R717 B.n200 B.n101 10.6151
R718 B.n204 B.n101 10.6151
R719 B.n207 B.n206 10.6151
R720 B.n207 B.n97 10.6151
R721 B.n211 B.n97 10.6151
R722 B.n212 B.n211 10.6151
R723 B.n213 B.n212 10.6151
R724 B.n213 B.n95 10.6151
R725 B.n217 B.n95 10.6151
R726 B.n218 B.n217 10.6151
R727 B.n220 B.n91 10.6151
R728 B.n224 B.n91 10.6151
R729 B.n225 B.n224 10.6151
R730 B.n226 B.n225 10.6151
R731 B.n226 B.n89 10.6151
R732 B.n230 B.n89 10.6151
R733 B.n231 B.n230 10.6151
R734 B.n232 B.n231 10.6151
R735 B.n232 B.n87 10.6151
R736 B.n236 B.n87 10.6151
R737 B.n237 B.n236 10.6151
R738 B.n238 B.n237 10.6151
R739 B.n238 B.n85 10.6151
R740 B.n242 B.n85 10.6151
R741 B.n243 B.n242 10.6151
R742 B.n244 B.n243 10.6151
R743 B.n244 B.n83 10.6151
R744 B.n248 B.n83 10.6151
R745 B.n249 B.n248 10.6151
R746 B.n250 B.n249 10.6151
R747 B.n250 B.n81 10.6151
R748 B.n254 B.n81 10.6151
R749 B.n255 B.n254 10.6151
R750 B.n256 B.n255 10.6151
R751 B.n256 B.n79 10.6151
R752 B.n260 B.n79 10.6151
R753 B.n261 B.n260 10.6151
R754 B.n262 B.n261 10.6151
R755 B.n262 B.n77 10.6151
R756 B.n266 B.n77 10.6151
R757 B.n267 B.n266 10.6151
R758 B.n268 B.n267 10.6151
R759 B.n268 B.n75 10.6151
R760 B.n272 B.n75 10.6151
R761 B.n273 B.n272 10.6151
R762 B.n274 B.n273 10.6151
R763 B.n274 B.n73 10.6151
R764 B.n278 B.n73 10.6151
R765 B.n477 B.n0 8.11757
R766 B.n477 B.n1 8.11757
R767 B.n395 B.n32 6.5566
R768 B.n383 B.n382 6.5566
R769 B.n206 B.n205 6.5566
R770 B.n219 B.n218 6.5566
R771 B.n32 B.n28 4.05904
R772 B.n382 B.n381 4.05904
R773 B.n205 B.n204 4.05904
R774 B.n220 B.n219 4.05904
R775 VP.n7 VP.t2 1334.1
R776 VP.n5 VP.t5 1334.1
R777 VP.n0 VP.t3 1334.1
R778 VP.n2 VP.t1 1334.1
R779 VP.n6 VP.t4 1288.83
R780 VP.n1 VP.t0 1288.83
R781 VP.n3 VP.n0 161.489
R782 VP.n8 VP.n7 161.3
R783 VP.n3 VP.n2 161.3
R784 VP.n5 VP.n4 161.3
R785 VP.n4 VP.n3 38.6975
R786 VP.n6 VP.n5 36.5157
R787 VP.n7 VP.n6 36.5157
R788 VP.n1 VP.n0 36.5157
R789 VP.n2 VP.n1 36.5157
R790 VP.n8 VP.n4 0.189894
R791 VP VP.n8 0.0516364
R792 VDD1 VDD1.t2 77.9045
R793 VDD1.n1 VDD1.t0 77.7908
R794 VDD1.n1 VDD1.n0 74.5944
R795 VDD1.n3 VDD1.n2 74.5291
R796 VDD1.n3 VDD1.n1 35.5914
R797 VDD1.n2 VDD1.t5 2.9555
R798 VDD1.n2 VDD1.t4 2.9555
R799 VDD1.n0 VDD1.t1 2.9555
R800 VDD1.n0 VDD1.t3 2.9555
R801 VDD1 VDD1.n3 0.063
C0 VDD1 VTAIL 14.283f
C1 VDD2 w_n1418_n3168# 1.60538f
C2 VTAIL w_n1418_n3168# 2.84938f
C3 VTAIL VDD2 14.312301f
C4 VP VN 4.43611f
C5 B VN 0.651454f
C6 VP B 0.93458f
C7 VDD1 VN 0.147637f
C8 w_n1418_n3168# VN 2.09463f
C9 VDD2 VN 2.16151f
C10 VDD1 VP 2.26708f
C11 VTAIL VN 1.70281f
C12 VDD1 B 1.33905f
C13 VP w_n1418_n3168# 2.27135f
C14 B w_n1418_n3168# 6.16985f
C15 VP VDD2 0.258013f
C16 B VDD2 1.3578f
C17 VTAIL VP 1.71755f
C18 VTAIL B 2.22356f
C19 VDD1 w_n1418_n3168# 1.59517f
C20 VDD1 VDD2 0.54538f
C21 VDD2 VSUBS 1.326684f
C22 VDD1 VSUBS 1.57865f
C23 VTAIL VSUBS 0.535091f
C24 VN VSUBS 3.91109f
C25 VP VSUBS 1.075837f
C26 B VSUBS 2.197097f
C27 w_n1418_n3168# VSUBS 55.3871f
C28 VDD1.t2 VSUBS 2.60808f
C29 VDD1.t0 VSUBS 2.60702f
C30 VDD1.t1 VSUBS 0.25937f
C31 VDD1.t3 VSUBS 0.25937f
C32 VDD1.n0 VSUBS 1.99045f
C33 VDD1.n1 VSUBS 2.87976f
C34 VDD1.t5 VSUBS 0.25937f
C35 VDD1.t4 VSUBS 0.25937f
C36 VDD1.n2 VSUBS 1.9899f
C37 VDD1.n3 VSUBS 2.74531f
C38 VP.t3 VSUBS 0.475616f
C39 VP.n0 VSUBS 0.2127f
C40 VP.t0 VSUBS 0.468996f
C41 VP.n1 VSUBS 0.19344f
C42 VP.t1 VSUBS 0.475616f
C43 VP.n2 VSUBS 0.212607f
C44 VP.n3 VSUBS 2.43049f
C45 VP.n4 VSUBS 2.41195f
C46 VP.t4 VSUBS 0.468996f
C47 VP.t5 VSUBS 0.475616f
C48 VP.n5 VSUBS 0.212607f
C49 VP.n6 VSUBS 0.19344f
C50 VP.t2 VSUBS 0.475616f
C51 VP.n7 VSUBS 0.212607f
C52 VP.n8 VSUBS 0.050799f
C53 B.n0 VSUBS 0.007067f
C54 B.n1 VSUBS 0.007067f
C55 B.n2 VSUBS 0.010452f
C56 B.n3 VSUBS 0.008009f
C57 B.n4 VSUBS 0.008009f
C58 B.n5 VSUBS 0.008009f
C59 B.n6 VSUBS 0.008009f
C60 B.n7 VSUBS 0.008009f
C61 B.n8 VSUBS 0.008009f
C62 B.n9 VSUBS 0.019923f
C63 B.n10 VSUBS 0.008009f
C64 B.n11 VSUBS 0.008009f
C65 B.n12 VSUBS 0.008009f
C66 B.n13 VSUBS 0.008009f
C67 B.n14 VSUBS 0.008009f
C68 B.n15 VSUBS 0.008009f
C69 B.n16 VSUBS 0.008009f
C70 B.n17 VSUBS 0.008009f
C71 B.n18 VSUBS 0.008009f
C72 B.n19 VSUBS 0.008009f
C73 B.n20 VSUBS 0.008009f
C74 B.n21 VSUBS 0.008009f
C75 B.n22 VSUBS 0.008009f
C76 B.n23 VSUBS 0.008009f
C77 B.n24 VSUBS 0.008009f
C78 B.n25 VSUBS 0.008009f
C79 B.n26 VSUBS 0.008009f
C80 B.n27 VSUBS 0.008009f
C81 B.n28 VSUBS 0.005536f
C82 B.n29 VSUBS 0.008009f
C83 B.t7 VSUBS 0.40618f
C84 B.t8 VSUBS 0.411532f
C85 B.t6 VSUBS 0.112933f
C86 B.n30 VSUBS 0.098048f
C87 B.n31 VSUBS 0.070825f
C88 B.n32 VSUBS 0.018557f
C89 B.n33 VSUBS 0.008009f
C90 B.n34 VSUBS 0.008009f
C91 B.n35 VSUBS 0.008009f
C92 B.n36 VSUBS 0.008009f
C93 B.t4 VSUBS 0.406173f
C94 B.t5 VSUBS 0.411526f
C95 B.t3 VSUBS 0.112933f
C96 B.n37 VSUBS 0.098054f
C97 B.n38 VSUBS 0.070831f
C98 B.n39 VSUBS 0.008009f
C99 B.n40 VSUBS 0.008009f
C100 B.n41 VSUBS 0.008009f
C101 B.n42 VSUBS 0.008009f
C102 B.n43 VSUBS 0.008009f
C103 B.n44 VSUBS 0.008009f
C104 B.n45 VSUBS 0.008009f
C105 B.n46 VSUBS 0.008009f
C106 B.n47 VSUBS 0.008009f
C107 B.n48 VSUBS 0.008009f
C108 B.n49 VSUBS 0.008009f
C109 B.n50 VSUBS 0.008009f
C110 B.n51 VSUBS 0.008009f
C111 B.n52 VSUBS 0.008009f
C112 B.n53 VSUBS 0.008009f
C113 B.n54 VSUBS 0.008009f
C114 B.n55 VSUBS 0.008009f
C115 B.n56 VSUBS 0.008009f
C116 B.n57 VSUBS 0.019923f
C117 B.n58 VSUBS 0.008009f
C118 B.n59 VSUBS 0.008009f
C119 B.n60 VSUBS 0.008009f
C120 B.n61 VSUBS 0.008009f
C121 B.n62 VSUBS 0.008009f
C122 B.n63 VSUBS 0.008009f
C123 B.n64 VSUBS 0.008009f
C124 B.n65 VSUBS 0.008009f
C125 B.n66 VSUBS 0.008009f
C126 B.n67 VSUBS 0.008009f
C127 B.n68 VSUBS 0.008009f
C128 B.n69 VSUBS 0.008009f
C129 B.n70 VSUBS 0.008009f
C130 B.n71 VSUBS 0.008009f
C131 B.n72 VSUBS 0.018711f
C132 B.n73 VSUBS 0.008009f
C133 B.n74 VSUBS 0.008009f
C134 B.n75 VSUBS 0.008009f
C135 B.n76 VSUBS 0.008009f
C136 B.n77 VSUBS 0.008009f
C137 B.n78 VSUBS 0.008009f
C138 B.n79 VSUBS 0.008009f
C139 B.n80 VSUBS 0.008009f
C140 B.n81 VSUBS 0.008009f
C141 B.n82 VSUBS 0.008009f
C142 B.n83 VSUBS 0.008009f
C143 B.n84 VSUBS 0.008009f
C144 B.n85 VSUBS 0.008009f
C145 B.n86 VSUBS 0.008009f
C146 B.n87 VSUBS 0.008009f
C147 B.n88 VSUBS 0.008009f
C148 B.n89 VSUBS 0.008009f
C149 B.n90 VSUBS 0.008009f
C150 B.n91 VSUBS 0.008009f
C151 B.n92 VSUBS 0.008009f
C152 B.t11 VSUBS 0.406173f
C153 B.t10 VSUBS 0.411526f
C154 B.t9 VSUBS 0.112933f
C155 B.n93 VSUBS 0.098054f
C156 B.n94 VSUBS 0.070831f
C157 B.n95 VSUBS 0.008009f
C158 B.n96 VSUBS 0.008009f
C159 B.n97 VSUBS 0.008009f
C160 B.n98 VSUBS 0.008009f
C161 B.t2 VSUBS 0.40618f
C162 B.t1 VSUBS 0.411532f
C163 B.t0 VSUBS 0.112933f
C164 B.n99 VSUBS 0.098048f
C165 B.n100 VSUBS 0.070825f
C166 B.n101 VSUBS 0.008009f
C167 B.n102 VSUBS 0.008009f
C168 B.n103 VSUBS 0.008009f
C169 B.n104 VSUBS 0.008009f
C170 B.n105 VSUBS 0.008009f
C171 B.n106 VSUBS 0.008009f
C172 B.n107 VSUBS 0.008009f
C173 B.n108 VSUBS 0.008009f
C174 B.n109 VSUBS 0.008009f
C175 B.n110 VSUBS 0.008009f
C176 B.n111 VSUBS 0.008009f
C177 B.n112 VSUBS 0.008009f
C178 B.n113 VSUBS 0.008009f
C179 B.n114 VSUBS 0.008009f
C180 B.n115 VSUBS 0.008009f
C181 B.n116 VSUBS 0.008009f
C182 B.n117 VSUBS 0.008009f
C183 B.n118 VSUBS 0.008009f
C184 B.n119 VSUBS 0.008009f
C185 B.n120 VSUBS 0.018711f
C186 B.n121 VSUBS 0.008009f
C187 B.n122 VSUBS 0.008009f
C188 B.n123 VSUBS 0.008009f
C189 B.n124 VSUBS 0.008009f
C190 B.n125 VSUBS 0.008009f
C191 B.n126 VSUBS 0.008009f
C192 B.n127 VSUBS 0.008009f
C193 B.n128 VSUBS 0.008009f
C194 B.n129 VSUBS 0.008009f
C195 B.n130 VSUBS 0.008009f
C196 B.n131 VSUBS 0.008009f
C197 B.n132 VSUBS 0.008009f
C198 B.n133 VSUBS 0.008009f
C199 B.n134 VSUBS 0.008009f
C200 B.n135 VSUBS 0.008009f
C201 B.n136 VSUBS 0.008009f
C202 B.n137 VSUBS 0.008009f
C203 B.n138 VSUBS 0.008009f
C204 B.n139 VSUBS 0.008009f
C205 B.n140 VSUBS 0.008009f
C206 B.n141 VSUBS 0.008009f
C207 B.n142 VSUBS 0.008009f
C208 B.n143 VSUBS 0.008009f
C209 B.n144 VSUBS 0.008009f
C210 B.n145 VSUBS 0.018711f
C211 B.n146 VSUBS 0.019923f
C212 B.n147 VSUBS 0.019923f
C213 B.n148 VSUBS 0.008009f
C214 B.n149 VSUBS 0.008009f
C215 B.n150 VSUBS 0.008009f
C216 B.n151 VSUBS 0.008009f
C217 B.n152 VSUBS 0.008009f
C218 B.n153 VSUBS 0.008009f
C219 B.n154 VSUBS 0.008009f
C220 B.n155 VSUBS 0.008009f
C221 B.n156 VSUBS 0.008009f
C222 B.n157 VSUBS 0.008009f
C223 B.n158 VSUBS 0.008009f
C224 B.n159 VSUBS 0.008009f
C225 B.n160 VSUBS 0.008009f
C226 B.n161 VSUBS 0.008009f
C227 B.n162 VSUBS 0.008009f
C228 B.n163 VSUBS 0.008009f
C229 B.n164 VSUBS 0.008009f
C230 B.n165 VSUBS 0.008009f
C231 B.n166 VSUBS 0.008009f
C232 B.n167 VSUBS 0.008009f
C233 B.n168 VSUBS 0.008009f
C234 B.n169 VSUBS 0.008009f
C235 B.n170 VSUBS 0.008009f
C236 B.n171 VSUBS 0.008009f
C237 B.n172 VSUBS 0.008009f
C238 B.n173 VSUBS 0.008009f
C239 B.n174 VSUBS 0.008009f
C240 B.n175 VSUBS 0.008009f
C241 B.n176 VSUBS 0.008009f
C242 B.n177 VSUBS 0.008009f
C243 B.n178 VSUBS 0.008009f
C244 B.n179 VSUBS 0.008009f
C245 B.n180 VSUBS 0.008009f
C246 B.n181 VSUBS 0.008009f
C247 B.n182 VSUBS 0.008009f
C248 B.n183 VSUBS 0.008009f
C249 B.n184 VSUBS 0.008009f
C250 B.n185 VSUBS 0.008009f
C251 B.n186 VSUBS 0.008009f
C252 B.n187 VSUBS 0.008009f
C253 B.n188 VSUBS 0.008009f
C254 B.n189 VSUBS 0.008009f
C255 B.n190 VSUBS 0.008009f
C256 B.n191 VSUBS 0.008009f
C257 B.n192 VSUBS 0.008009f
C258 B.n193 VSUBS 0.008009f
C259 B.n194 VSUBS 0.008009f
C260 B.n195 VSUBS 0.008009f
C261 B.n196 VSUBS 0.008009f
C262 B.n197 VSUBS 0.008009f
C263 B.n198 VSUBS 0.008009f
C264 B.n199 VSUBS 0.008009f
C265 B.n200 VSUBS 0.008009f
C266 B.n201 VSUBS 0.008009f
C267 B.n202 VSUBS 0.008009f
C268 B.n203 VSUBS 0.008009f
C269 B.n204 VSUBS 0.005536f
C270 B.n205 VSUBS 0.018557f
C271 B.n206 VSUBS 0.006478f
C272 B.n207 VSUBS 0.008009f
C273 B.n208 VSUBS 0.008009f
C274 B.n209 VSUBS 0.008009f
C275 B.n210 VSUBS 0.008009f
C276 B.n211 VSUBS 0.008009f
C277 B.n212 VSUBS 0.008009f
C278 B.n213 VSUBS 0.008009f
C279 B.n214 VSUBS 0.008009f
C280 B.n215 VSUBS 0.008009f
C281 B.n216 VSUBS 0.008009f
C282 B.n217 VSUBS 0.008009f
C283 B.n218 VSUBS 0.006478f
C284 B.n219 VSUBS 0.018557f
C285 B.n220 VSUBS 0.005536f
C286 B.n221 VSUBS 0.008009f
C287 B.n222 VSUBS 0.008009f
C288 B.n223 VSUBS 0.008009f
C289 B.n224 VSUBS 0.008009f
C290 B.n225 VSUBS 0.008009f
C291 B.n226 VSUBS 0.008009f
C292 B.n227 VSUBS 0.008009f
C293 B.n228 VSUBS 0.008009f
C294 B.n229 VSUBS 0.008009f
C295 B.n230 VSUBS 0.008009f
C296 B.n231 VSUBS 0.008009f
C297 B.n232 VSUBS 0.008009f
C298 B.n233 VSUBS 0.008009f
C299 B.n234 VSUBS 0.008009f
C300 B.n235 VSUBS 0.008009f
C301 B.n236 VSUBS 0.008009f
C302 B.n237 VSUBS 0.008009f
C303 B.n238 VSUBS 0.008009f
C304 B.n239 VSUBS 0.008009f
C305 B.n240 VSUBS 0.008009f
C306 B.n241 VSUBS 0.008009f
C307 B.n242 VSUBS 0.008009f
C308 B.n243 VSUBS 0.008009f
C309 B.n244 VSUBS 0.008009f
C310 B.n245 VSUBS 0.008009f
C311 B.n246 VSUBS 0.008009f
C312 B.n247 VSUBS 0.008009f
C313 B.n248 VSUBS 0.008009f
C314 B.n249 VSUBS 0.008009f
C315 B.n250 VSUBS 0.008009f
C316 B.n251 VSUBS 0.008009f
C317 B.n252 VSUBS 0.008009f
C318 B.n253 VSUBS 0.008009f
C319 B.n254 VSUBS 0.008009f
C320 B.n255 VSUBS 0.008009f
C321 B.n256 VSUBS 0.008009f
C322 B.n257 VSUBS 0.008009f
C323 B.n258 VSUBS 0.008009f
C324 B.n259 VSUBS 0.008009f
C325 B.n260 VSUBS 0.008009f
C326 B.n261 VSUBS 0.008009f
C327 B.n262 VSUBS 0.008009f
C328 B.n263 VSUBS 0.008009f
C329 B.n264 VSUBS 0.008009f
C330 B.n265 VSUBS 0.008009f
C331 B.n266 VSUBS 0.008009f
C332 B.n267 VSUBS 0.008009f
C333 B.n268 VSUBS 0.008009f
C334 B.n269 VSUBS 0.008009f
C335 B.n270 VSUBS 0.008009f
C336 B.n271 VSUBS 0.008009f
C337 B.n272 VSUBS 0.008009f
C338 B.n273 VSUBS 0.008009f
C339 B.n274 VSUBS 0.008009f
C340 B.n275 VSUBS 0.008009f
C341 B.n276 VSUBS 0.008009f
C342 B.n277 VSUBS 0.019923f
C343 B.n278 VSUBS 0.019019f
C344 B.n279 VSUBS 0.019615f
C345 B.n280 VSUBS 0.008009f
C346 B.n281 VSUBS 0.008009f
C347 B.n282 VSUBS 0.008009f
C348 B.n283 VSUBS 0.008009f
C349 B.n284 VSUBS 0.008009f
C350 B.n285 VSUBS 0.008009f
C351 B.n286 VSUBS 0.008009f
C352 B.n287 VSUBS 0.008009f
C353 B.n288 VSUBS 0.008009f
C354 B.n289 VSUBS 0.008009f
C355 B.n290 VSUBS 0.008009f
C356 B.n291 VSUBS 0.008009f
C357 B.n292 VSUBS 0.008009f
C358 B.n293 VSUBS 0.008009f
C359 B.n294 VSUBS 0.008009f
C360 B.n295 VSUBS 0.008009f
C361 B.n296 VSUBS 0.008009f
C362 B.n297 VSUBS 0.008009f
C363 B.n298 VSUBS 0.008009f
C364 B.n299 VSUBS 0.008009f
C365 B.n300 VSUBS 0.008009f
C366 B.n301 VSUBS 0.008009f
C367 B.n302 VSUBS 0.008009f
C368 B.n303 VSUBS 0.008009f
C369 B.n304 VSUBS 0.008009f
C370 B.n305 VSUBS 0.008009f
C371 B.n306 VSUBS 0.008009f
C372 B.n307 VSUBS 0.008009f
C373 B.n308 VSUBS 0.008009f
C374 B.n309 VSUBS 0.008009f
C375 B.n310 VSUBS 0.008009f
C376 B.n311 VSUBS 0.008009f
C377 B.n312 VSUBS 0.008009f
C378 B.n313 VSUBS 0.008009f
C379 B.n314 VSUBS 0.008009f
C380 B.n315 VSUBS 0.008009f
C381 B.n316 VSUBS 0.008009f
C382 B.n317 VSUBS 0.008009f
C383 B.n318 VSUBS 0.008009f
C384 B.n319 VSUBS 0.008009f
C385 B.n320 VSUBS 0.008009f
C386 B.n321 VSUBS 0.008009f
C387 B.n322 VSUBS 0.018711f
C388 B.n323 VSUBS 0.018711f
C389 B.n324 VSUBS 0.019923f
C390 B.n325 VSUBS 0.008009f
C391 B.n326 VSUBS 0.008009f
C392 B.n327 VSUBS 0.008009f
C393 B.n328 VSUBS 0.008009f
C394 B.n329 VSUBS 0.008009f
C395 B.n330 VSUBS 0.008009f
C396 B.n331 VSUBS 0.008009f
C397 B.n332 VSUBS 0.008009f
C398 B.n333 VSUBS 0.008009f
C399 B.n334 VSUBS 0.008009f
C400 B.n335 VSUBS 0.008009f
C401 B.n336 VSUBS 0.008009f
C402 B.n337 VSUBS 0.008009f
C403 B.n338 VSUBS 0.008009f
C404 B.n339 VSUBS 0.008009f
C405 B.n340 VSUBS 0.008009f
C406 B.n341 VSUBS 0.008009f
C407 B.n342 VSUBS 0.008009f
C408 B.n343 VSUBS 0.008009f
C409 B.n344 VSUBS 0.008009f
C410 B.n345 VSUBS 0.008009f
C411 B.n346 VSUBS 0.008009f
C412 B.n347 VSUBS 0.008009f
C413 B.n348 VSUBS 0.008009f
C414 B.n349 VSUBS 0.008009f
C415 B.n350 VSUBS 0.008009f
C416 B.n351 VSUBS 0.008009f
C417 B.n352 VSUBS 0.008009f
C418 B.n353 VSUBS 0.008009f
C419 B.n354 VSUBS 0.008009f
C420 B.n355 VSUBS 0.008009f
C421 B.n356 VSUBS 0.008009f
C422 B.n357 VSUBS 0.008009f
C423 B.n358 VSUBS 0.008009f
C424 B.n359 VSUBS 0.008009f
C425 B.n360 VSUBS 0.008009f
C426 B.n361 VSUBS 0.008009f
C427 B.n362 VSUBS 0.008009f
C428 B.n363 VSUBS 0.008009f
C429 B.n364 VSUBS 0.008009f
C430 B.n365 VSUBS 0.008009f
C431 B.n366 VSUBS 0.008009f
C432 B.n367 VSUBS 0.008009f
C433 B.n368 VSUBS 0.008009f
C434 B.n369 VSUBS 0.008009f
C435 B.n370 VSUBS 0.008009f
C436 B.n371 VSUBS 0.008009f
C437 B.n372 VSUBS 0.008009f
C438 B.n373 VSUBS 0.008009f
C439 B.n374 VSUBS 0.008009f
C440 B.n375 VSUBS 0.008009f
C441 B.n376 VSUBS 0.008009f
C442 B.n377 VSUBS 0.008009f
C443 B.n378 VSUBS 0.008009f
C444 B.n379 VSUBS 0.008009f
C445 B.n380 VSUBS 0.008009f
C446 B.n381 VSUBS 0.005536f
C447 B.n382 VSUBS 0.018557f
C448 B.n383 VSUBS 0.006478f
C449 B.n384 VSUBS 0.008009f
C450 B.n385 VSUBS 0.008009f
C451 B.n386 VSUBS 0.008009f
C452 B.n387 VSUBS 0.008009f
C453 B.n388 VSUBS 0.008009f
C454 B.n389 VSUBS 0.008009f
C455 B.n390 VSUBS 0.008009f
C456 B.n391 VSUBS 0.008009f
C457 B.n392 VSUBS 0.008009f
C458 B.n393 VSUBS 0.008009f
C459 B.n394 VSUBS 0.008009f
C460 B.n395 VSUBS 0.006478f
C461 B.n396 VSUBS 0.008009f
C462 B.n397 VSUBS 0.008009f
C463 B.n398 VSUBS 0.008009f
C464 B.n399 VSUBS 0.008009f
C465 B.n400 VSUBS 0.008009f
C466 B.n401 VSUBS 0.008009f
C467 B.n402 VSUBS 0.008009f
C468 B.n403 VSUBS 0.008009f
C469 B.n404 VSUBS 0.008009f
C470 B.n405 VSUBS 0.008009f
C471 B.n406 VSUBS 0.008009f
C472 B.n407 VSUBS 0.008009f
C473 B.n408 VSUBS 0.008009f
C474 B.n409 VSUBS 0.008009f
C475 B.n410 VSUBS 0.008009f
C476 B.n411 VSUBS 0.008009f
C477 B.n412 VSUBS 0.008009f
C478 B.n413 VSUBS 0.008009f
C479 B.n414 VSUBS 0.008009f
C480 B.n415 VSUBS 0.008009f
C481 B.n416 VSUBS 0.008009f
C482 B.n417 VSUBS 0.008009f
C483 B.n418 VSUBS 0.008009f
C484 B.n419 VSUBS 0.008009f
C485 B.n420 VSUBS 0.008009f
C486 B.n421 VSUBS 0.008009f
C487 B.n422 VSUBS 0.008009f
C488 B.n423 VSUBS 0.008009f
C489 B.n424 VSUBS 0.008009f
C490 B.n425 VSUBS 0.008009f
C491 B.n426 VSUBS 0.008009f
C492 B.n427 VSUBS 0.008009f
C493 B.n428 VSUBS 0.008009f
C494 B.n429 VSUBS 0.008009f
C495 B.n430 VSUBS 0.008009f
C496 B.n431 VSUBS 0.008009f
C497 B.n432 VSUBS 0.008009f
C498 B.n433 VSUBS 0.008009f
C499 B.n434 VSUBS 0.008009f
C500 B.n435 VSUBS 0.008009f
C501 B.n436 VSUBS 0.008009f
C502 B.n437 VSUBS 0.008009f
C503 B.n438 VSUBS 0.008009f
C504 B.n439 VSUBS 0.008009f
C505 B.n440 VSUBS 0.008009f
C506 B.n441 VSUBS 0.008009f
C507 B.n442 VSUBS 0.008009f
C508 B.n443 VSUBS 0.008009f
C509 B.n444 VSUBS 0.008009f
C510 B.n445 VSUBS 0.008009f
C511 B.n446 VSUBS 0.008009f
C512 B.n447 VSUBS 0.008009f
C513 B.n448 VSUBS 0.008009f
C514 B.n449 VSUBS 0.008009f
C515 B.n450 VSUBS 0.008009f
C516 B.n451 VSUBS 0.008009f
C517 B.n452 VSUBS 0.008009f
C518 B.n453 VSUBS 0.008009f
C519 B.n454 VSUBS 0.019923f
C520 B.n455 VSUBS 0.018711f
C521 B.n456 VSUBS 0.018711f
C522 B.n457 VSUBS 0.008009f
C523 B.n458 VSUBS 0.008009f
C524 B.n459 VSUBS 0.008009f
C525 B.n460 VSUBS 0.008009f
C526 B.n461 VSUBS 0.008009f
C527 B.n462 VSUBS 0.008009f
C528 B.n463 VSUBS 0.008009f
C529 B.n464 VSUBS 0.008009f
C530 B.n465 VSUBS 0.008009f
C531 B.n466 VSUBS 0.008009f
C532 B.n467 VSUBS 0.008009f
C533 B.n468 VSUBS 0.008009f
C534 B.n469 VSUBS 0.008009f
C535 B.n470 VSUBS 0.008009f
C536 B.n471 VSUBS 0.008009f
C537 B.n472 VSUBS 0.008009f
C538 B.n473 VSUBS 0.008009f
C539 B.n474 VSUBS 0.008009f
C540 B.n475 VSUBS 0.010452f
C541 B.n476 VSUBS 0.011134f
C542 B.n477 VSUBS 0.022141f
C543 VDD2.t1 VSUBS 2.60863f
C544 VDD2.t0 VSUBS 0.25953f
C545 VDD2.t4 VSUBS 0.25953f
C546 VDD2.n0 VSUBS 1.99169f
C547 VDD2.n1 VSUBS 2.80243f
C548 VDD2.t5 VSUBS 2.60592f
C549 VDD2.n2 VSUBS 2.79684f
C550 VDD2.t3 VSUBS 0.25953f
C551 VDD2.t2 VSUBS 0.25953f
C552 VDD2.n3 VSUBS 1.99165f
C553 VTAIL.t6 VSUBS 0.280018f
C554 VTAIL.t9 VSUBS 0.280018f
C555 VTAIL.n0 VSUBS 1.97765f
C556 VTAIL.n1 VSUBS 0.817329f
C557 VTAIL.t2 VSUBS 2.62172f
C558 VTAIL.n2 VSUBS 0.968493f
C559 VTAIL.t4 VSUBS 0.280018f
C560 VTAIL.t5 VSUBS 0.280018f
C561 VTAIL.n3 VSUBS 1.97765f
C562 VTAIL.n4 VSUBS 2.29716f
C563 VTAIL.t7 VSUBS 0.280018f
C564 VTAIL.t10 VSUBS 0.280018f
C565 VTAIL.n5 VSUBS 1.97766f
C566 VTAIL.n6 VSUBS 2.29715f
C567 VTAIL.t11 VSUBS 2.62174f
C568 VTAIL.n7 VSUBS 0.968474f
C569 VTAIL.t0 VSUBS 0.280018f
C570 VTAIL.t3 VSUBS 0.280018f
C571 VTAIL.n8 VSUBS 1.97766f
C572 VTAIL.n9 VSUBS 0.848863f
C573 VTAIL.t1 VSUBS 2.62172f
C574 VTAIL.n10 VSUBS 2.36667f
C575 VTAIL.t8 VSUBS 2.62172f
C576 VTAIL.n11 VSUBS 2.3481f
C577 VN.t4 VSUBS 0.455103f
C578 VN.n0 VSUBS 0.203527f
C579 VN.t5 VSUBS 0.448768f
C580 VN.n1 VSUBS 0.185097f
C581 VN.t1 VSUBS 0.455103f
C582 VN.n2 VSUBS 0.203437f
C583 VN.n3 VSUBS 0.124778f
C584 VN.t3 VSUBS 0.455103f
C585 VN.n4 VSUBS 0.203527f
C586 VN.t0 VSUBS 0.455103f
C587 VN.t2 VSUBS 0.448768f
C588 VN.n5 VSUBS 0.185097f
C589 VN.n6 VSUBS 0.203437f
C590 VN.n7 VSUBS 2.36706f
.ends

