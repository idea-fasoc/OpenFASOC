* NGSPICE file created from diff_pair_sample_0957.ext - technology: sky130A

.subckt diff_pair_sample_0957 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VN.t0 VDD2.t1 B.t5 sky130_fd_pr__nfet_01v8 ad=0.15015 pd=1.24 as=0.15015 ps=1.24 w=0.91 l=0.94
X1 VTAIL.t14 VN.t1 VDD2.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=0.3549 pd=2.6 as=0.15015 ps=1.24 w=0.91 l=0.94
X2 B.t21 B.t19 B.t20 B.t9 sky130_fd_pr__nfet_01v8 ad=0.3549 pd=2.6 as=0 ps=0 w=0.91 l=0.94
X3 B.t18 B.t16 B.t17 B.t13 sky130_fd_pr__nfet_01v8 ad=0.3549 pd=2.6 as=0 ps=0 w=0.91 l=0.94
X4 VDD2.t6 VN.t2 VTAIL.t13 B.t4 sky130_fd_pr__nfet_01v8 ad=0.15015 pd=1.24 as=0.15015 ps=1.24 w=0.91 l=0.94
X5 VDD2.t5 VN.t3 VTAIL.t12 B.t3 sky130_fd_pr__nfet_01v8 ad=0.15015 pd=1.24 as=0.3549 ps=2.6 w=0.91 l=0.94
X6 VTAIL.t11 VN.t4 VDD2.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=0.15015 pd=1.24 as=0.15015 ps=1.24 w=0.91 l=0.94
X7 VDD1.t7 VP.t0 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.15015 pd=1.24 as=0.3549 ps=2.6 w=0.91 l=0.94
X8 VDD2.t2 VN.t5 VTAIL.t10 B.t0 sky130_fd_pr__nfet_01v8 ad=0.15015 pd=1.24 as=0.15015 ps=1.24 w=0.91 l=0.94
X9 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=0.3549 pd=2.6 as=0 ps=0 w=0.91 l=0.94
X10 VTAIL.t7 VP.t1 VDD1.t6 B.t7 sky130_fd_pr__nfet_01v8 ad=0.3549 pd=2.6 as=0.15015 ps=1.24 w=0.91 l=0.94
X11 VTAIL.t9 VN.t6 VDD2.t4 B.t7 sky130_fd_pr__nfet_01v8 ad=0.3549 pd=2.6 as=0.15015 ps=1.24 w=0.91 l=0.94
X12 VDD1.t5 VP.t2 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=0.15015 pd=1.24 as=0.15015 ps=1.24 w=0.91 l=0.94
X13 VDD2.t7 VN.t7 VTAIL.t8 B.t6 sky130_fd_pr__nfet_01v8 ad=0.15015 pd=1.24 as=0.3549 ps=2.6 w=0.91 l=0.94
X14 VTAIL.t5 VP.t3 VDD1.t4 B.t5 sky130_fd_pr__nfet_01v8 ad=0.15015 pd=1.24 as=0.15015 ps=1.24 w=0.91 l=0.94
X15 VDD1.t3 VP.t4 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=0.15015 pd=1.24 as=0.3549 ps=2.6 w=0.91 l=0.94
X16 VTAIL.t2 VP.t5 VDD1.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.15015 pd=1.24 as=0.15015 ps=1.24 w=0.91 l=0.94
X17 VDD1.t1 VP.t6 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.15015 pd=1.24 as=0.15015 ps=1.24 w=0.91 l=0.94
X18 VTAIL.t1 VP.t7 VDD1.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=0.3549 pd=2.6 as=0.15015 ps=1.24 w=0.91 l=0.94
X19 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=0.3549 pd=2.6 as=0 ps=0 w=0.91 l=0.94
R0 VN.n23 VN.n13 161.3
R1 VN.n21 VN.n20 161.3
R2 VN.n19 VN.n14 161.3
R3 VN.n18 VN.n17 161.3
R4 VN.n10 VN.n0 161.3
R5 VN.n8 VN.n7 161.3
R6 VN.n6 VN.n1 161.3
R7 VN.n5 VN.n4 161.3
R8 VN.n25 VN.n24 80.6037
R9 VN.n12 VN.n11 80.6037
R10 VN.n2 VN.t1 79.9777
R11 VN.n15 VN.t7 79.9777
R12 VN.n11 VN.t3 65.3782
R13 VN.n24 VN.t6 65.3782
R14 VN.n11 VN.n10 53.3386
R15 VN.n24 VN.n23 53.3386
R16 VN.n3 VN.n2 46.9742
R17 VN.n16 VN.n15 46.9742
R18 VN.n18 VN.n15 44.3395
R19 VN.n5 VN.n2 44.3395
R20 VN.n4 VN.n1 40.4934
R21 VN.n8 VN.n1 40.4934
R22 VN.n17 VN.n14 40.4934
R23 VN.n21 VN.n14 40.4934
R24 VN VN.n25 35.143
R25 VN.n3 VN.t2 23.3314
R26 VN.n9 VN.t0 23.3314
R27 VN.n16 VN.t4 23.3314
R28 VN.n22 VN.t5 23.3314
R29 VN.n10 VN.n9 17.8614
R30 VN.n23 VN.n22 17.8614
R31 VN.n4 VN.n3 6.60659
R32 VN.n9 VN.n8 6.60659
R33 VN.n17 VN.n16 6.60659
R34 VN.n22 VN.n21 6.60659
R35 VN.n25 VN.n13 0.285035
R36 VN.n12 VN.n0 0.285035
R37 VN.n20 VN.n13 0.189894
R38 VN.n20 VN.n19 0.189894
R39 VN.n19 VN.n18 0.189894
R40 VN.n6 VN.n5 0.189894
R41 VN.n7 VN.n6 0.189894
R42 VN.n7 VN.n0 0.189894
R43 VN VN.n12 0.146778
R44 VDD2.n2 VDD2.n1 238.879
R45 VDD2.n2 VDD2.n0 238.879
R46 VDD2 VDD2.n5 238.876
R47 VDD2.n4 VDD2.n3 238.387
R48 VDD2.n4 VDD2.n2 29.4265
R49 VDD2.n5 VDD2.t3 21.7587
R50 VDD2.n5 VDD2.t7 21.7587
R51 VDD2.n3 VDD2.t4 21.7587
R52 VDD2.n3 VDD2.t2 21.7587
R53 VDD2.n1 VDD2.t1 21.7587
R54 VDD2.n1 VDD2.t5 21.7587
R55 VDD2.n0 VDD2.t0 21.7587
R56 VDD2.n0 VDD2.t6 21.7587
R57 VDD2 VDD2.n4 0.606103
R58 VTAIL.n14 VTAIL.t3 243.466
R59 VTAIL.n11 VTAIL.t1 243.466
R60 VTAIL.n10 VTAIL.t8 243.466
R61 VTAIL.n7 VTAIL.t9 243.466
R62 VTAIL.n15 VTAIL.t12 243.465
R63 VTAIL.n2 VTAIL.t14 243.465
R64 VTAIL.n3 VTAIL.t6 243.465
R65 VTAIL.n6 VTAIL.t7 243.465
R66 VTAIL.n13 VTAIL.n12 221.708
R67 VTAIL.n9 VTAIL.n8 221.708
R68 VTAIL.n1 VTAIL.n0 221.708
R69 VTAIL.n5 VTAIL.n4 221.708
R70 VTAIL.n0 VTAIL.t13 21.7587
R71 VTAIL.n0 VTAIL.t15 21.7587
R72 VTAIL.n4 VTAIL.t0 21.7587
R73 VTAIL.n4 VTAIL.t2 21.7587
R74 VTAIL.n12 VTAIL.t4 21.7587
R75 VTAIL.n12 VTAIL.t5 21.7587
R76 VTAIL.n8 VTAIL.t10 21.7587
R77 VTAIL.n8 VTAIL.t11 21.7587
R78 VTAIL.n15 VTAIL.n14 14.2462
R79 VTAIL.n7 VTAIL.n6 14.2462
R80 VTAIL.n9 VTAIL.n7 1.09533
R81 VTAIL.n10 VTAIL.n9 1.09533
R82 VTAIL.n13 VTAIL.n11 1.09533
R83 VTAIL.n14 VTAIL.n13 1.09533
R84 VTAIL.n6 VTAIL.n5 1.09533
R85 VTAIL.n5 VTAIL.n3 1.09533
R86 VTAIL.n2 VTAIL.n1 1.09533
R87 VTAIL VTAIL.n15 1.03714
R88 VTAIL.n11 VTAIL.n10 0.470328
R89 VTAIL.n3 VTAIL.n2 0.470328
R90 VTAIL VTAIL.n1 0.0586897
R91 B.n310 B.n309 585
R92 B.n312 B.n70 585
R93 B.n315 B.n314 585
R94 B.n316 B.n69 585
R95 B.n318 B.n317 585
R96 B.n320 B.n68 585
R97 B.n323 B.n322 585
R98 B.n324 B.n64 585
R99 B.n326 B.n325 585
R100 B.n328 B.n63 585
R101 B.n331 B.n330 585
R102 B.n332 B.n62 585
R103 B.n334 B.n333 585
R104 B.n336 B.n61 585
R105 B.n339 B.n338 585
R106 B.n340 B.n60 585
R107 B.n342 B.n341 585
R108 B.n344 B.n59 585
R109 B.n347 B.n346 585
R110 B.n349 B.n56 585
R111 B.n351 B.n350 585
R112 B.n353 B.n55 585
R113 B.n356 B.n355 585
R114 B.n357 B.n54 585
R115 B.n359 B.n358 585
R116 B.n361 B.n53 585
R117 B.n364 B.n363 585
R118 B.n365 B.n52 585
R119 B.n308 B.n50 585
R120 B.n368 B.n50 585
R121 B.n307 B.n49 585
R122 B.n369 B.n49 585
R123 B.n306 B.n48 585
R124 B.n370 B.n48 585
R125 B.n305 B.n304 585
R126 B.n304 B.n44 585
R127 B.n303 B.n43 585
R128 B.n376 B.n43 585
R129 B.n302 B.n42 585
R130 B.n377 B.n42 585
R131 B.n301 B.n41 585
R132 B.n378 B.n41 585
R133 B.n300 B.n299 585
R134 B.n299 B.n37 585
R135 B.n298 B.n36 585
R136 B.n384 B.n36 585
R137 B.n297 B.n35 585
R138 B.n385 B.n35 585
R139 B.n296 B.n34 585
R140 B.n386 B.n34 585
R141 B.n295 B.n294 585
R142 B.n294 B.n33 585
R143 B.n293 B.n29 585
R144 B.n392 B.n29 585
R145 B.n292 B.n28 585
R146 B.n393 B.n28 585
R147 B.n291 B.n27 585
R148 B.n394 B.n27 585
R149 B.n290 B.n289 585
R150 B.n289 B.n26 585
R151 B.n288 B.n22 585
R152 B.n400 B.n22 585
R153 B.n287 B.n21 585
R154 B.n401 B.n21 585
R155 B.n286 B.n20 585
R156 B.n402 B.n20 585
R157 B.n285 B.n284 585
R158 B.n284 B.n19 585
R159 B.n283 B.n15 585
R160 B.n408 B.n15 585
R161 B.n282 B.n14 585
R162 B.n409 B.n14 585
R163 B.n281 B.n13 585
R164 B.n410 B.n13 585
R165 B.n280 B.n279 585
R166 B.n279 B.n12 585
R167 B.n278 B.n277 585
R168 B.n278 B.n8 585
R169 B.n276 B.n7 585
R170 B.n417 B.n7 585
R171 B.n275 B.n6 585
R172 B.n418 B.n6 585
R173 B.n274 B.n5 585
R174 B.n419 B.n5 585
R175 B.n273 B.n272 585
R176 B.n272 B.n4 585
R177 B.n271 B.n71 585
R178 B.n271 B.n270 585
R179 B.n260 B.n72 585
R180 B.n263 B.n72 585
R181 B.n262 B.n261 585
R182 B.n264 B.n262 585
R183 B.n259 B.n77 585
R184 B.n77 B.n76 585
R185 B.n258 B.n257 585
R186 B.n257 B.n256 585
R187 B.n79 B.n78 585
R188 B.n249 B.n79 585
R189 B.n248 B.n247 585
R190 B.n250 B.n248 585
R191 B.n246 B.n84 585
R192 B.n84 B.n83 585
R193 B.n245 B.n244 585
R194 B.n244 B.n243 585
R195 B.n86 B.n85 585
R196 B.n236 B.n86 585
R197 B.n235 B.n234 585
R198 B.n237 B.n235 585
R199 B.n233 B.n91 585
R200 B.n91 B.n90 585
R201 B.n232 B.n231 585
R202 B.n231 B.n230 585
R203 B.n93 B.n92 585
R204 B.n223 B.n93 585
R205 B.n222 B.n221 585
R206 B.n224 B.n222 585
R207 B.n220 B.n98 585
R208 B.n98 B.n97 585
R209 B.n219 B.n218 585
R210 B.n218 B.n217 585
R211 B.n100 B.n99 585
R212 B.n101 B.n100 585
R213 B.n210 B.n209 585
R214 B.n211 B.n210 585
R215 B.n208 B.n106 585
R216 B.n106 B.n105 585
R217 B.n207 B.n206 585
R218 B.n206 B.n205 585
R219 B.n108 B.n107 585
R220 B.n109 B.n108 585
R221 B.n198 B.n197 585
R222 B.n199 B.n198 585
R223 B.n196 B.n114 585
R224 B.n114 B.n113 585
R225 B.n195 B.n194 585
R226 B.n194 B.n193 585
R227 B.n190 B.n118 585
R228 B.n189 B.n188 585
R229 B.n186 B.n119 585
R230 B.n186 B.n117 585
R231 B.n185 B.n184 585
R232 B.n183 B.n182 585
R233 B.n181 B.n121 585
R234 B.n179 B.n178 585
R235 B.n177 B.n122 585
R236 B.n176 B.n175 585
R237 B.n173 B.n172 585
R238 B.n171 B.n170 585
R239 B.n169 B.n127 585
R240 B.n167 B.n166 585
R241 B.n165 B.n128 585
R242 B.n164 B.n163 585
R243 B.n161 B.n129 585
R244 B.n159 B.n158 585
R245 B.n157 B.n130 585
R246 B.n156 B.n155 585
R247 B.n153 B.n152 585
R248 B.n151 B.n150 585
R249 B.n149 B.n135 585
R250 B.n147 B.n146 585
R251 B.n145 B.n136 585
R252 B.n144 B.n143 585
R253 B.n141 B.n137 585
R254 B.n139 B.n138 585
R255 B.n116 B.n115 585
R256 B.n117 B.n116 585
R257 B.n192 B.n191 585
R258 B.n193 B.n192 585
R259 B.n112 B.n111 585
R260 B.n113 B.n112 585
R261 B.n201 B.n200 585
R262 B.n200 B.n199 585
R263 B.n202 B.n110 585
R264 B.n110 B.n109 585
R265 B.n204 B.n203 585
R266 B.n205 B.n204 585
R267 B.n104 B.n103 585
R268 B.n105 B.n104 585
R269 B.n213 B.n212 585
R270 B.n212 B.n211 585
R271 B.n214 B.n102 585
R272 B.n102 B.n101 585
R273 B.n216 B.n215 585
R274 B.n217 B.n216 585
R275 B.n96 B.n95 585
R276 B.n97 B.n96 585
R277 B.n226 B.n225 585
R278 B.n225 B.n224 585
R279 B.n227 B.n94 585
R280 B.n223 B.n94 585
R281 B.n229 B.n228 585
R282 B.n230 B.n229 585
R283 B.n89 B.n88 585
R284 B.n90 B.n89 585
R285 B.n239 B.n238 585
R286 B.n238 B.n237 585
R287 B.n240 B.n87 585
R288 B.n236 B.n87 585
R289 B.n242 B.n241 585
R290 B.n243 B.n242 585
R291 B.n82 B.n81 585
R292 B.n83 B.n82 585
R293 B.n252 B.n251 585
R294 B.n251 B.n250 585
R295 B.n253 B.n80 585
R296 B.n249 B.n80 585
R297 B.n255 B.n254 585
R298 B.n256 B.n255 585
R299 B.n75 B.n74 585
R300 B.n76 B.n75 585
R301 B.n266 B.n265 585
R302 B.n265 B.n264 585
R303 B.n267 B.n73 585
R304 B.n263 B.n73 585
R305 B.n269 B.n268 585
R306 B.n270 B.n269 585
R307 B.n3 B.n0 585
R308 B.n4 B.n3 585
R309 B.n416 B.n1 585
R310 B.n417 B.n416 585
R311 B.n415 B.n414 585
R312 B.n415 B.n8 585
R313 B.n413 B.n9 585
R314 B.n12 B.n9 585
R315 B.n412 B.n411 585
R316 B.n411 B.n410 585
R317 B.n11 B.n10 585
R318 B.n409 B.n11 585
R319 B.n407 B.n406 585
R320 B.n408 B.n407 585
R321 B.n405 B.n16 585
R322 B.n19 B.n16 585
R323 B.n404 B.n403 585
R324 B.n403 B.n402 585
R325 B.n18 B.n17 585
R326 B.n401 B.n18 585
R327 B.n399 B.n398 585
R328 B.n400 B.n399 585
R329 B.n397 B.n23 585
R330 B.n26 B.n23 585
R331 B.n396 B.n395 585
R332 B.n395 B.n394 585
R333 B.n25 B.n24 585
R334 B.n393 B.n25 585
R335 B.n391 B.n390 585
R336 B.n392 B.n391 585
R337 B.n389 B.n30 585
R338 B.n33 B.n30 585
R339 B.n388 B.n387 585
R340 B.n387 B.n386 585
R341 B.n32 B.n31 585
R342 B.n385 B.n32 585
R343 B.n383 B.n382 585
R344 B.n384 B.n383 585
R345 B.n381 B.n38 585
R346 B.n38 B.n37 585
R347 B.n380 B.n379 585
R348 B.n379 B.n378 585
R349 B.n40 B.n39 585
R350 B.n377 B.n40 585
R351 B.n375 B.n374 585
R352 B.n376 B.n375 585
R353 B.n373 B.n45 585
R354 B.n45 B.n44 585
R355 B.n372 B.n371 585
R356 B.n371 B.n370 585
R357 B.n47 B.n46 585
R358 B.n369 B.n47 585
R359 B.n367 B.n366 585
R360 B.n368 B.n367 585
R361 B.n420 B.n419 585
R362 B.n418 B.n2 585
R363 B.n367 B.n52 511.721
R364 B.n310 B.n50 511.721
R365 B.n194 B.n116 511.721
R366 B.n192 B.n118 511.721
R367 B.n57 B.t17 258.928
R368 B.n65 B.t14 258.928
R369 B.n131 B.t11 258.928
R370 B.n123 B.t21 258.928
R371 B.n311 B.n51 256.663
R372 B.n313 B.n51 256.663
R373 B.n319 B.n51 256.663
R374 B.n321 B.n51 256.663
R375 B.n327 B.n51 256.663
R376 B.n329 B.n51 256.663
R377 B.n335 B.n51 256.663
R378 B.n337 B.n51 256.663
R379 B.n343 B.n51 256.663
R380 B.n345 B.n51 256.663
R381 B.n352 B.n51 256.663
R382 B.n354 B.n51 256.663
R383 B.n360 B.n51 256.663
R384 B.n362 B.n51 256.663
R385 B.n187 B.n117 256.663
R386 B.n120 B.n117 256.663
R387 B.n180 B.n117 256.663
R388 B.n174 B.n117 256.663
R389 B.n126 B.n117 256.663
R390 B.n168 B.n117 256.663
R391 B.n162 B.n117 256.663
R392 B.n160 B.n117 256.663
R393 B.n154 B.n117 256.663
R394 B.n134 B.n117 256.663
R395 B.n148 B.n117 256.663
R396 B.n142 B.n117 256.663
R397 B.n140 B.n117 256.663
R398 B.n422 B.n421 256.663
R399 B.n193 B.n117 254.326
R400 B.n368 B.n51 254.326
R401 B.n58 B.t18 234.298
R402 B.n66 B.t15 234.298
R403 B.n132 B.t10 234.298
R404 B.n124 B.t20 234.298
R405 B.n65 B.t12 226.472
R406 B.n131 B.t8 226.472
R407 B.n57 B.t16 225.881
R408 B.n123 B.t19 225.881
R409 B.n363 B.n361 163.367
R410 B.n359 B.n54 163.367
R411 B.n355 B.n353 163.367
R412 B.n351 B.n56 163.367
R413 B.n346 B.n344 163.367
R414 B.n342 B.n60 163.367
R415 B.n338 B.n336 163.367
R416 B.n334 B.n62 163.367
R417 B.n330 B.n328 163.367
R418 B.n326 B.n64 163.367
R419 B.n322 B.n320 163.367
R420 B.n318 B.n69 163.367
R421 B.n314 B.n312 163.367
R422 B.n194 B.n114 163.367
R423 B.n198 B.n114 163.367
R424 B.n198 B.n108 163.367
R425 B.n206 B.n108 163.367
R426 B.n206 B.n106 163.367
R427 B.n210 B.n106 163.367
R428 B.n210 B.n100 163.367
R429 B.n218 B.n100 163.367
R430 B.n218 B.n98 163.367
R431 B.n222 B.n98 163.367
R432 B.n222 B.n93 163.367
R433 B.n231 B.n93 163.367
R434 B.n231 B.n91 163.367
R435 B.n235 B.n91 163.367
R436 B.n235 B.n86 163.367
R437 B.n244 B.n86 163.367
R438 B.n244 B.n84 163.367
R439 B.n248 B.n84 163.367
R440 B.n248 B.n79 163.367
R441 B.n257 B.n79 163.367
R442 B.n257 B.n77 163.367
R443 B.n262 B.n77 163.367
R444 B.n262 B.n72 163.367
R445 B.n271 B.n72 163.367
R446 B.n272 B.n271 163.367
R447 B.n272 B.n5 163.367
R448 B.n6 B.n5 163.367
R449 B.n7 B.n6 163.367
R450 B.n278 B.n7 163.367
R451 B.n279 B.n278 163.367
R452 B.n279 B.n13 163.367
R453 B.n14 B.n13 163.367
R454 B.n15 B.n14 163.367
R455 B.n284 B.n15 163.367
R456 B.n284 B.n20 163.367
R457 B.n21 B.n20 163.367
R458 B.n22 B.n21 163.367
R459 B.n289 B.n22 163.367
R460 B.n289 B.n27 163.367
R461 B.n28 B.n27 163.367
R462 B.n29 B.n28 163.367
R463 B.n294 B.n29 163.367
R464 B.n294 B.n34 163.367
R465 B.n35 B.n34 163.367
R466 B.n36 B.n35 163.367
R467 B.n299 B.n36 163.367
R468 B.n299 B.n41 163.367
R469 B.n42 B.n41 163.367
R470 B.n43 B.n42 163.367
R471 B.n304 B.n43 163.367
R472 B.n304 B.n48 163.367
R473 B.n49 B.n48 163.367
R474 B.n50 B.n49 163.367
R475 B.n188 B.n186 163.367
R476 B.n186 B.n185 163.367
R477 B.n182 B.n181 163.367
R478 B.n179 B.n122 163.367
R479 B.n175 B.n173 163.367
R480 B.n170 B.n169 163.367
R481 B.n167 B.n128 163.367
R482 B.n163 B.n161 163.367
R483 B.n159 B.n130 163.367
R484 B.n155 B.n153 163.367
R485 B.n150 B.n149 163.367
R486 B.n147 B.n136 163.367
R487 B.n143 B.n141 163.367
R488 B.n139 B.n116 163.367
R489 B.n192 B.n112 163.367
R490 B.n200 B.n112 163.367
R491 B.n200 B.n110 163.367
R492 B.n204 B.n110 163.367
R493 B.n204 B.n104 163.367
R494 B.n212 B.n104 163.367
R495 B.n212 B.n102 163.367
R496 B.n216 B.n102 163.367
R497 B.n216 B.n96 163.367
R498 B.n225 B.n96 163.367
R499 B.n225 B.n94 163.367
R500 B.n229 B.n94 163.367
R501 B.n229 B.n89 163.367
R502 B.n238 B.n89 163.367
R503 B.n238 B.n87 163.367
R504 B.n242 B.n87 163.367
R505 B.n242 B.n82 163.367
R506 B.n251 B.n82 163.367
R507 B.n251 B.n80 163.367
R508 B.n255 B.n80 163.367
R509 B.n255 B.n75 163.367
R510 B.n265 B.n75 163.367
R511 B.n265 B.n73 163.367
R512 B.n269 B.n73 163.367
R513 B.n269 B.n3 163.367
R514 B.n420 B.n3 163.367
R515 B.n416 B.n2 163.367
R516 B.n416 B.n415 163.367
R517 B.n415 B.n9 163.367
R518 B.n411 B.n9 163.367
R519 B.n411 B.n11 163.367
R520 B.n407 B.n11 163.367
R521 B.n407 B.n16 163.367
R522 B.n403 B.n16 163.367
R523 B.n403 B.n18 163.367
R524 B.n399 B.n18 163.367
R525 B.n399 B.n23 163.367
R526 B.n395 B.n23 163.367
R527 B.n395 B.n25 163.367
R528 B.n391 B.n25 163.367
R529 B.n391 B.n30 163.367
R530 B.n387 B.n30 163.367
R531 B.n387 B.n32 163.367
R532 B.n383 B.n32 163.367
R533 B.n383 B.n38 163.367
R534 B.n379 B.n38 163.367
R535 B.n379 B.n40 163.367
R536 B.n375 B.n40 163.367
R537 B.n375 B.n45 163.367
R538 B.n371 B.n45 163.367
R539 B.n371 B.n47 163.367
R540 B.n367 B.n47 163.367
R541 B.n193 B.n113 120.939
R542 B.n199 B.n113 120.939
R543 B.n199 B.n109 120.939
R544 B.n205 B.n109 120.939
R545 B.n211 B.n105 120.939
R546 B.n211 B.n101 120.939
R547 B.n217 B.n101 120.939
R548 B.n217 B.n97 120.939
R549 B.n224 B.n97 120.939
R550 B.n224 B.n223 120.939
R551 B.n230 B.n90 120.939
R552 B.n237 B.n90 120.939
R553 B.n237 B.n236 120.939
R554 B.n243 B.n83 120.939
R555 B.n250 B.n83 120.939
R556 B.n250 B.n249 120.939
R557 B.n256 B.n76 120.939
R558 B.n264 B.n76 120.939
R559 B.n264 B.n263 120.939
R560 B.n270 B.n4 120.939
R561 B.n419 B.n4 120.939
R562 B.n419 B.n418 120.939
R563 B.n418 B.n417 120.939
R564 B.n417 B.n8 120.939
R565 B.n410 B.n12 120.939
R566 B.n410 B.n409 120.939
R567 B.n409 B.n408 120.939
R568 B.n402 B.n19 120.939
R569 B.n402 B.n401 120.939
R570 B.n401 B.n400 120.939
R571 B.n394 B.n26 120.939
R572 B.n394 B.n393 120.939
R573 B.n393 B.n392 120.939
R574 B.n386 B.n33 120.939
R575 B.n386 B.n385 120.939
R576 B.n385 B.n384 120.939
R577 B.n384 B.n37 120.939
R578 B.n378 B.n37 120.939
R579 B.n378 B.n377 120.939
R580 B.n376 B.n44 120.939
R581 B.n370 B.n44 120.939
R582 B.n370 B.n369 120.939
R583 B.n369 B.n368 120.939
R584 B.n270 B.t6 117.382
R585 B.t1 B.n8 117.382
R586 B.n205 B.t9 106.71
R587 B.t13 B.n376 106.71
R588 B.n223 B.t7 99.5963
R589 B.n33 B.t3 99.5963
R590 B.n256 B.t2 85.3683
R591 B.n408 B.t4 85.3683
R592 B.n362 B.n52 71.676
R593 B.n361 B.n360 71.676
R594 B.n354 B.n54 71.676
R595 B.n353 B.n352 71.676
R596 B.n345 B.n56 71.676
R597 B.n344 B.n343 71.676
R598 B.n337 B.n60 71.676
R599 B.n336 B.n335 71.676
R600 B.n329 B.n62 71.676
R601 B.n328 B.n327 71.676
R602 B.n321 B.n64 71.676
R603 B.n320 B.n319 71.676
R604 B.n313 B.n69 71.676
R605 B.n312 B.n311 71.676
R606 B.n311 B.n310 71.676
R607 B.n314 B.n313 71.676
R608 B.n319 B.n318 71.676
R609 B.n322 B.n321 71.676
R610 B.n327 B.n326 71.676
R611 B.n330 B.n329 71.676
R612 B.n335 B.n334 71.676
R613 B.n338 B.n337 71.676
R614 B.n343 B.n342 71.676
R615 B.n346 B.n345 71.676
R616 B.n352 B.n351 71.676
R617 B.n355 B.n354 71.676
R618 B.n360 B.n359 71.676
R619 B.n363 B.n362 71.676
R620 B.n187 B.n118 71.676
R621 B.n185 B.n120 71.676
R622 B.n181 B.n180 71.676
R623 B.n174 B.n122 71.676
R624 B.n173 B.n126 71.676
R625 B.n169 B.n168 71.676
R626 B.n162 B.n128 71.676
R627 B.n161 B.n160 71.676
R628 B.n154 B.n130 71.676
R629 B.n153 B.n134 71.676
R630 B.n149 B.n148 71.676
R631 B.n142 B.n136 71.676
R632 B.n141 B.n140 71.676
R633 B.n188 B.n187 71.676
R634 B.n182 B.n120 71.676
R635 B.n180 B.n179 71.676
R636 B.n175 B.n174 71.676
R637 B.n170 B.n126 71.676
R638 B.n168 B.n167 71.676
R639 B.n163 B.n162 71.676
R640 B.n160 B.n159 71.676
R641 B.n155 B.n154 71.676
R642 B.n150 B.n134 71.676
R643 B.n148 B.n147 71.676
R644 B.n143 B.n142 71.676
R645 B.n140 B.n139 71.676
R646 B.n421 B.n420 71.676
R647 B.n421 B.n2 71.676
R648 B.n236 B.t0 67.5834
R649 B.n26 B.t5 67.5834
R650 B.n348 B.n58 59.5399
R651 B.n67 B.n66 59.5399
R652 B.n133 B.n132 59.5399
R653 B.n125 B.n124 59.5399
R654 B.n243 B.t0 53.3554
R655 B.n400 B.t5 53.3554
R656 B.n249 B.t2 35.5704
R657 B.n19 B.t4 35.5704
R658 B.n191 B.n190 33.2493
R659 B.n195 B.n115 33.2493
R660 B.n309 B.n308 33.2493
R661 B.n366 B.n365 33.2493
R662 B.n58 B.n57 24.6308
R663 B.n66 B.n65 24.6308
R664 B.n132 B.n131 24.6308
R665 B.n124 B.n123 24.6308
R666 B.n230 B.t7 21.3425
R667 B.n392 B.t3 21.3425
R668 B B.n422 18.0485
R669 B.t9 B.n105 14.2285
R670 B.n377 B.t13 14.2285
R671 B.n191 B.n111 10.6151
R672 B.n201 B.n111 10.6151
R673 B.n202 B.n201 10.6151
R674 B.n203 B.n202 10.6151
R675 B.n203 B.n103 10.6151
R676 B.n213 B.n103 10.6151
R677 B.n214 B.n213 10.6151
R678 B.n215 B.n214 10.6151
R679 B.n215 B.n95 10.6151
R680 B.n226 B.n95 10.6151
R681 B.n227 B.n226 10.6151
R682 B.n228 B.n227 10.6151
R683 B.n228 B.n88 10.6151
R684 B.n239 B.n88 10.6151
R685 B.n240 B.n239 10.6151
R686 B.n241 B.n240 10.6151
R687 B.n241 B.n81 10.6151
R688 B.n252 B.n81 10.6151
R689 B.n253 B.n252 10.6151
R690 B.n254 B.n253 10.6151
R691 B.n254 B.n74 10.6151
R692 B.n266 B.n74 10.6151
R693 B.n267 B.n266 10.6151
R694 B.n268 B.n267 10.6151
R695 B.n268 B.n0 10.6151
R696 B.n190 B.n189 10.6151
R697 B.n189 B.n119 10.6151
R698 B.n184 B.n119 10.6151
R699 B.n184 B.n183 10.6151
R700 B.n183 B.n121 10.6151
R701 B.n178 B.n121 10.6151
R702 B.n178 B.n177 10.6151
R703 B.n177 B.n176 10.6151
R704 B.n172 B.n171 10.6151
R705 B.n171 B.n127 10.6151
R706 B.n166 B.n127 10.6151
R707 B.n166 B.n165 10.6151
R708 B.n165 B.n164 10.6151
R709 B.n164 B.n129 10.6151
R710 B.n158 B.n129 10.6151
R711 B.n158 B.n157 10.6151
R712 B.n157 B.n156 10.6151
R713 B.n152 B.n151 10.6151
R714 B.n151 B.n135 10.6151
R715 B.n146 B.n135 10.6151
R716 B.n146 B.n145 10.6151
R717 B.n145 B.n144 10.6151
R718 B.n144 B.n137 10.6151
R719 B.n138 B.n137 10.6151
R720 B.n138 B.n115 10.6151
R721 B.n196 B.n195 10.6151
R722 B.n197 B.n196 10.6151
R723 B.n197 B.n107 10.6151
R724 B.n207 B.n107 10.6151
R725 B.n208 B.n207 10.6151
R726 B.n209 B.n208 10.6151
R727 B.n209 B.n99 10.6151
R728 B.n219 B.n99 10.6151
R729 B.n220 B.n219 10.6151
R730 B.n221 B.n220 10.6151
R731 B.n221 B.n92 10.6151
R732 B.n232 B.n92 10.6151
R733 B.n233 B.n232 10.6151
R734 B.n234 B.n233 10.6151
R735 B.n234 B.n85 10.6151
R736 B.n245 B.n85 10.6151
R737 B.n246 B.n245 10.6151
R738 B.n247 B.n246 10.6151
R739 B.n247 B.n78 10.6151
R740 B.n258 B.n78 10.6151
R741 B.n259 B.n258 10.6151
R742 B.n261 B.n259 10.6151
R743 B.n261 B.n260 10.6151
R744 B.n260 B.n71 10.6151
R745 B.n273 B.n71 10.6151
R746 B.n274 B.n273 10.6151
R747 B.n275 B.n274 10.6151
R748 B.n276 B.n275 10.6151
R749 B.n277 B.n276 10.6151
R750 B.n280 B.n277 10.6151
R751 B.n281 B.n280 10.6151
R752 B.n282 B.n281 10.6151
R753 B.n283 B.n282 10.6151
R754 B.n285 B.n283 10.6151
R755 B.n286 B.n285 10.6151
R756 B.n287 B.n286 10.6151
R757 B.n288 B.n287 10.6151
R758 B.n290 B.n288 10.6151
R759 B.n291 B.n290 10.6151
R760 B.n292 B.n291 10.6151
R761 B.n293 B.n292 10.6151
R762 B.n295 B.n293 10.6151
R763 B.n296 B.n295 10.6151
R764 B.n297 B.n296 10.6151
R765 B.n298 B.n297 10.6151
R766 B.n300 B.n298 10.6151
R767 B.n301 B.n300 10.6151
R768 B.n302 B.n301 10.6151
R769 B.n303 B.n302 10.6151
R770 B.n305 B.n303 10.6151
R771 B.n306 B.n305 10.6151
R772 B.n307 B.n306 10.6151
R773 B.n308 B.n307 10.6151
R774 B.n414 B.n1 10.6151
R775 B.n414 B.n413 10.6151
R776 B.n413 B.n412 10.6151
R777 B.n412 B.n10 10.6151
R778 B.n406 B.n10 10.6151
R779 B.n406 B.n405 10.6151
R780 B.n405 B.n404 10.6151
R781 B.n404 B.n17 10.6151
R782 B.n398 B.n17 10.6151
R783 B.n398 B.n397 10.6151
R784 B.n397 B.n396 10.6151
R785 B.n396 B.n24 10.6151
R786 B.n390 B.n24 10.6151
R787 B.n390 B.n389 10.6151
R788 B.n389 B.n388 10.6151
R789 B.n388 B.n31 10.6151
R790 B.n382 B.n31 10.6151
R791 B.n382 B.n381 10.6151
R792 B.n381 B.n380 10.6151
R793 B.n380 B.n39 10.6151
R794 B.n374 B.n39 10.6151
R795 B.n374 B.n373 10.6151
R796 B.n373 B.n372 10.6151
R797 B.n372 B.n46 10.6151
R798 B.n366 B.n46 10.6151
R799 B.n365 B.n364 10.6151
R800 B.n364 B.n53 10.6151
R801 B.n358 B.n53 10.6151
R802 B.n358 B.n357 10.6151
R803 B.n357 B.n356 10.6151
R804 B.n356 B.n55 10.6151
R805 B.n350 B.n55 10.6151
R806 B.n350 B.n349 10.6151
R807 B.n347 B.n59 10.6151
R808 B.n341 B.n59 10.6151
R809 B.n341 B.n340 10.6151
R810 B.n340 B.n339 10.6151
R811 B.n339 B.n61 10.6151
R812 B.n333 B.n61 10.6151
R813 B.n333 B.n332 10.6151
R814 B.n332 B.n331 10.6151
R815 B.n331 B.n63 10.6151
R816 B.n325 B.n324 10.6151
R817 B.n324 B.n323 10.6151
R818 B.n323 B.n68 10.6151
R819 B.n317 B.n68 10.6151
R820 B.n317 B.n316 10.6151
R821 B.n316 B.n315 10.6151
R822 B.n315 B.n70 10.6151
R823 B.n309 B.n70 10.6151
R824 B.n176 B.n125 9.52245
R825 B.n152 B.n133 9.52245
R826 B.n349 B.n348 9.52245
R827 B.n325 B.n67 9.52245
R828 B.n422 B.n0 8.11757
R829 B.n422 B.n1 8.11757
R830 B.n263 B.t6 3.55749
R831 B.n12 B.t1 3.55749
R832 B.n172 B.n125 1.09318
R833 B.n156 B.n133 1.09318
R834 B.n348 B.n347 1.09318
R835 B.n67 B.n63 1.09318
R836 VP.n8 VP.n7 161.3
R837 VP.n9 VP.n4 161.3
R838 VP.n11 VP.n10 161.3
R839 VP.n13 VP.n3 161.3
R840 VP.n26 VP.n0 161.3
R841 VP.n24 VP.n23 161.3
R842 VP.n22 VP.n1 161.3
R843 VP.n21 VP.n20 161.3
R844 VP.n18 VP.n2 161.3
R845 VP.n15 VP.n14 80.6037
R846 VP.n28 VP.n27 80.6037
R847 VP.n17 VP.n16 80.6037
R848 VP.n5 VP.t7 79.9777
R849 VP.n17 VP.t1 65.3782
R850 VP.n27 VP.t4 65.3782
R851 VP.n14 VP.t0 65.3782
R852 VP.n18 VP.n17 53.3386
R853 VP.n27 VP.n26 53.3386
R854 VP.n14 VP.n13 53.3386
R855 VP.n6 VP.n5 46.9742
R856 VP.n8 VP.n5 44.3395
R857 VP.n20 VP.n1 40.4934
R858 VP.n24 VP.n1 40.4934
R859 VP.n11 VP.n4 40.4934
R860 VP.n7 VP.n4 40.4934
R861 VP.n16 VP.n15 34.8574
R862 VP.n19 VP.t6 23.3314
R863 VP.n25 VP.t5 23.3314
R864 VP.n12 VP.t3 23.3314
R865 VP.n6 VP.t2 23.3314
R866 VP.n19 VP.n18 17.8614
R867 VP.n26 VP.n25 17.8614
R868 VP.n13 VP.n12 17.8614
R869 VP.n20 VP.n19 6.60659
R870 VP.n25 VP.n24 6.60659
R871 VP.n12 VP.n11 6.60659
R872 VP.n7 VP.n6 6.60659
R873 VP.n15 VP.n3 0.285035
R874 VP.n16 VP.n2 0.285035
R875 VP.n28 VP.n0 0.285035
R876 VP.n9 VP.n8 0.189894
R877 VP.n10 VP.n9 0.189894
R878 VP.n10 VP.n3 0.189894
R879 VP.n21 VP.n2 0.189894
R880 VP.n22 VP.n21 0.189894
R881 VP.n23 VP.n22 0.189894
R882 VP.n23 VP.n0 0.189894
R883 VP VP.n28 0.146778
R884 VDD1 VDD1.n0 238.994
R885 VDD1.n3 VDD1.n2 238.879
R886 VDD1.n3 VDD1.n1 238.879
R887 VDD1.n5 VDD1.n4 238.387
R888 VDD1.n5 VDD1.n3 30.0095
R889 VDD1.n4 VDD1.t4 21.7587
R890 VDD1.n4 VDD1.t7 21.7587
R891 VDD1.n0 VDD1.t0 21.7587
R892 VDD1.n0 VDD1.t5 21.7587
R893 VDD1.n2 VDD1.t2 21.7587
R894 VDD1.n2 VDD1.t3 21.7587
R895 VDD1.n1 VDD1.t6 21.7587
R896 VDD1.n1 VDD1.t1 21.7587
R897 VDD1 VDD1.n5 0.489724
C0 VP VDD1 1.04466f
C1 VDD1 VDD2 0.946147f
C2 VP VTAIL 1.36185f
C3 VTAIL VDD2 2.95873f
C4 VN VP 3.59014f
C5 VN VDD2 0.851058f
C6 VTAIL VDD1 2.91544f
C7 VN VDD1 0.156047f
C8 VN VTAIL 1.34774f
C9 VP VDD2 0.351712f
C10 VDD2 B 2.704578f
C11 VDD1 B 2.944176f
C12 VTAIL B 2.492844f
C13 VN B 7.639896f
C14 VP B 6.640119f
C15 VDD1.t0 B 0.013251f
C16 VDD1.t5 B 0.013251f
C17 VDD1.n0 B 0.05201f
C18 VDD1.t6 B 0.013251f
C19 VDD1.t1 B 0.013251f
C20 VDD1.n1 B 0.051889f
C21 VDD1.t2 B 0.013251f
C22 VDD1.t3 B 0.013251f
C23 VDD1.n2 B 0.051889f
C24 VDD1.n3 B 1.20617f
C25 VDD1.t4 B 0.013251f
C26 VDD1.t7 B 0.013251f
C27 VDD1.n4 B 0.051428f
C28 VDD1.n5 B 1.08623f
C29 VP.n0 B 0.038494f
C30 VP.t5 B 0.043317f
C31 VP.n1 B 0.023321f
C32 VP.n2 B 0.038494f
C33 VP.t6 B 0.043317f
C34 VP.n3 B 0.038494f
C35 VP.t0 B 0.084861f
C36 VP.t3 B 0.043317f
C37 VP.n4 B 0.023321f
C38 VP.t7 B 0.101258f
C39 VP.n5 B 0.08749f
C40 VP.t2 B 0.043317f
C41 VP.n6 B 0.071884f
C42 VP.n7 B 0.037956f
C43 VP.n8 B 0.119266f
C44 VP.n9 B 0.028848f
C45 VP.n10 B 0.028848f
C46 VP.n11 B 0.037956f
C47 VP.n12 B 0.049593f
C48 VP.n13 B 0.035966f
C49 VP.n14 B 0.08964f
C50 VP.n15 B 0.863112f
C51 VP.n16 B 0.892861f
C52 VP.t1 B 0.084861f
C53 VP.n17 B 0.08964f
C54 VP.n18 B 0.035966f
C55 VP.n19 B 0.049593f
C56 VP.n20 B 0.037956f
C57 VP.n21 B 0.028848f
C58 VP.n22 B 0.028848f
C59 VP.n23 B 0.028848f
C60 VP.n24 B 0.037956f
C61 VP.n25 B 0.049593f
C62 VP.n26 B 0.035966f
C63 VP.t4 B 0.084861f
C64 VP.n27 B 0.08964f
C65 VP.n28 B 0.027017f
C66 VTAIL.t13 B 0.016392f
C67 VTAIL.t15 B 0.016392f
C68 VTAIL.n0 B 0.052631f
C69 VTAIL.n1 B 0.215048f
C70 VTAIL.t14 B 0.090102f
C71 VTAIL.n2 B 0.252516f
C72 VTAIL.t6 B 0.090102f
C73 VTAIL.n3 B 0.252516f
C74 VTAIL.t0 B 0.016392f
C75 VTAIL.t2 B 0.016392f
C76 VTAIL.n4 B 0.052631f
C77 VTAIL.n5 B 0.291188f
C78 VTAIL.t7 B 0.090102f
C79 VTAIL.n6 B 0.665679f
C80 VTAIL.t9 B 0.090102f
C81 VTAIL.n7 B 0.665679f
C82 VTAIL.t10 B 0.016392f
C83 VTAIL.t11 B 0.016392f
C84 VTAIL.n8 B 0.052631f
C85 VTAIL.n9 B 0.291188f
C86 VTAIL.t8 B 0.090102f
C87 VTAIL.n10 B 0.252516f
C88 VTAIL.t1 B 0.090102f
C89 VTAIL.n11 B 0.252516f
C90 VTAIL.t4 B 0.016392f
C91 VTAIL.t5 B 0.016392f
C92 VTAIL.n12 B 0.052631f
C93 VTAIL.n13 B 0.291188f
C94 VTAIL.t3 B 0.090102f
C95 VTAIL.n14 B 0.665679f
C96 VTAIL.t12 B 0.090102f
C97 VTAIL.n15 B 0.661405f
C98 VDD2.t0 B 0.014038f
C99 VDD2.t6 B 0.014038f
C100 VDD2.n0 B 0.054968f
C101 VDD2.t1 B 0.014038f
C102 VDD2.t5 B 0.014038f
C103 VDD2.n1 B 0.054968f
C104 VDD2.n2 B 1.2361f
C105 VDD2.t4 B 0.014038f
C106 VDD2.t2 B 0.014038f
C107 VDD2.n3 B 0.054479f
C108 VDD2.n4 B 1.12757f
C109 VDD2.t3 B 0.014038f
C110 VDD2.t7 B 0.014038f
C111 VDD2.n5 B 0.054963f
C112 VN.n0 B 0.038065f
C113 VN.t0 B 0.042834f
C114 VN.n1 B 0.023061f
C115 VN.t1 B 0.10013f
C116 VN.n2 B 0.086516f
C117 VN.t2 B 0.042834f
C118 VN.n3 B 0.071083f
C119 VN.n4 B 0.037534f
C120 VN.n5 B 0.117937f
C121 VN.n6 B 0.028527f
C122 VN.n7 B 0.028527f
C123 VN.n8 B 0.037534f
C124 VN.n9 B 0.049041f
C125 VN.n10 B 0.035565f
C126 VN.t3 B 0.083915f
C127 VN.n11 B 0.088641f
C128 VN.n12 B 0.026716f
C129 VN.n13 B 0.038065f
C130 VN.t5 B 0.042834f
C131 VN.n14 B 0.023061f
C132 VN.t7 B 0.10013f
C133 VN.n15 B 0.086516f
C134 VN.t4 B 0.042834f
C135 VN.n16 B 0.071083f
C136 VN.n17 B 0.037534f
C137 VN.n18 B 0.117937f
C138 VN.n19 B 0.028527f
C139 VN.n20 B 0.028527f
C140 VN.n21 B 0.037534f
C141 VN.n22 B 0.049041f
C142 VN.n23 B 0.035565f
C143 VN.t6 B 0.083915f
C144 VN.n24 B 0.088641f
C145 VN.n25 B 0.870081f
.ends

