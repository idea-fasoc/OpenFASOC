* NGSPICE file created from diff_pair_sample_1472.ext - technology: sky130A

.subckt diff_pair_sample_1472 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t1 VN.t0 VTAIL.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=4.9998 pd=26.42 as=4.9998 ps=26.42 w=12.82 l=0.41
X1 B.t15 B.t13 B.t14 B.t10 sky130_fd_pr__nfet_01v8 ad=4.9998 pd=26.42 as=0 ps=0 w=12.82 l=0.41
X2 B.t12 B.t9 B.t11 B.t10 sky130_fd_pr__nfet_01v8 ad=4.9998 pd=26.42 as=0 ps=0 w=12.82 l=0.41
X3 B.t8 B.t6 B.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=4.9998 pd=26.42 as=0 ps=0 w=12.82 l=0.41
X4 VDD1.t1 VP.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=4.9998 pd=26.42 as=4.9998 ps=26.42 w=12.82 l=0.41
X5 VDD1.t0 VP.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=4.9998 pd=26.42 as=4.9998 ps=26.42 w=12.82 l=0.41
X6 VDD2.t0 VN.t1 VTAIL.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=4.9998 pd=26.42 as=4.9998 ps=26.42 w=12.82 l=0.41
X7 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=4.9998 pd=26.42 as=0 ps=0 w=12.82 l=0.41
R0 VN VN.t0 1051.72
R1 VN VN.t1 1011.9
R2 VTAIL.n274 VTAIL.n210 289.615
R3 VTAIL.n64 VTAIL.n0 289.615
R4 VTAIL.n204 VTAIL.n140 289.615
R5 VTAIL.n134 VTAIL.n70 289.615
R6 VTAIL.n233 VTAIL.n232 185
R7 VTAIL.n230 VTAIL.n229 185
R8 VTAIL.n239 VTAIL.n238 185
R9 VTAIL.n241 VTAIL.n240 185
R10 VTAIL.n226 VTAIL.n225 185
R11 VTAIL.n247 VTAIL.n246 185
R12 VTAIL.n250 VTAIL.n249 185
R13 VTAIL.n248 VTAIL.n222 185
R14 VTAIL.n255 VTAIL.n221 185
R15 VTAIL.n257 VTAIL.n256 185
R16 VTAIL.n259 VTAIL.n258 185
R17 VTAIL.n218 VTAIL.n217 185
R18 VTAIL.n265 VTAIL.n264 185
R19 VTAIL.n267 VTAIL.n266 185
R20 VTAIL.n214 VTAIL.n213 185
R21 VTAIL.n273 VTAIL.n272 185
R22 VTAIL.n275 VTAIL.n274 185
R23 VTAIL.n23 VTAIL.n22 185
R24 VTAIL.n20 VTAIL.n19 185
R25 VTAIL.n29 VTAIL.n28 185
R26 VTAIL.n31 VTAIL.n30 185
R27 VTAIL.n16 VTAIL.n15 185
R28 VTAIL.n37 VTAIL.n36 185
R29 VTAIL.n40 VTAIL.n39 185
R30 VTAIL.n38 VTAIL.n12 185
R31 VTAIL.n45 VTAIL.n11 185
R32 VTAIL.n47 VTAIL.n46 185
R33 VTAIL.n49 VTAIL.n48 185
R34 VTAIL.n8 VTAIL.n7 185
R35 VTAIL.n55 VTAIL.n54 185
R36 VTAIL.n57 VTAIL.n56 185
R37 VTAIL.n4 VTAIL.n3 185
R38 VTAIL.n63 VTAIL.n62 185
R39 VTAIL.n65 VTAIL.n64 185
R40 VTAIL.n205 VTAIL.n204 185
R41 VTAIL.n203 VTAIL.n202 185
R42 VTAIL.n144 VTAIL.n143 185
R43 VTAIL.n197 VTAIL.n196 185
R44 VTAIL.n195 VTAIL.n194 185
R45 VTAIL.n148 VTAIL.n147 185
R46 VTAIL.n189 VTAIL.n188 185
R47 VTAIL.n187 VTAIL.n186 185
R48 VTAIL.n185 VTAIL.n151 185
R49 VTAIL.n155 VTAIL.n152 185
R50 VTAIL.n180 VTAIL.n179 185
R51 VTAIL.n178 VTAIL.n177 185
R52 VTAIL.n157 VTAIL.n156 185
R53 VTAIL.n172 VTAIL.n171 185
R54 VTAIL.n170 VTAIL.n169 185
R55 VTAIL.n161 VTAIL.n160 185
R56 VTAIL.n164 VTAIL.n163 185
R57 VTAIL.n135 VTAIL.n134 185
R58 VTAIL.n133 VTAIL.n132 185
R59 VTAIL.n74 VTAIL.n73 185
R60 VTAIL.n127 VTAIL.n126 185
R61 VTAIL.n125 VTAIL.n124 185
R62 VTAIL.n78 VTAIL.n77 185
R63 VTAIL.n119 VTAIL.n118 185
R64 VTAIL.n117 VTAIL.n116 185
R65 VTAIL.n115 VTAIL.n81 185
R66 VTAIL.n85 VTAIL.n82 185
R67 VTAIL.n110 VTAIL.n109 185
R68 VTAIL.n108 VTAIL.n107 185
R69 VTAIL.n87 VTAIL.n86 185
R70 VTAIL.n102 VTAIL.n101 185
R71 VTAIL.n100 VTAIL.n99 185
R72 VTAIL.n91 VTAIL.n90 185
R73 VTAIL.n94 VTAIL.n93 185
R74 VTAIL.t3 VTAIL.n231 149.524
R75 VTAIL.t1 VTAIL.n21 149.524
R76 VTAIL.t0 VTAIL.n162 149.524
R77 VTAIL.t2 VTAIL.n92 149.524
R78 VTAIL.n232 VTAIL.n229 104.615
R79 VTAIL.n239 VTAIL.n229 104.615
R80 VTAIL.n240 VTAIL.n239 104.615
R81 VTAIL.n240 VTAIL.n225 104.615
R82 VTAIL.n247 VTAIL.n225 104.615
R83 VTAIL.n249 VTAIL.n247 104.615
R84 VTAIL.n249 VTAIL.n248 104.615
R85 VTAIL.n248 VTAIL.n221 104.615
R86 VTAIL.n257 VTAIL.n221 104.615
R87 VTAIL.n258 VTAIL.n257 104.615
R88 VTAIL.n258 VTAIL.n217 104.615
R89 VTAIL.n265 VTAIL.n217 104.615
R90 VTAIL.n266 VTAIL.n265 104.615
R91 VTAIL.n266 VTAIL.n213 104.615
R92 VTAIL.n273 VTAIL.n213 104.615
R93 VTAIL.n274 VTAIL.n273 104.615
R94 VTAIL.n22 VTAIL.n19 104.615
R95 VTAIL.n29 VTAIL.n19 104.615
R96 VTAIL.n30 VTAIL.n29 104.615
R97 VTAIL.n30 VTAIL.n15 104.615
R98 VTAIL.n37 VTAIL.n15 104.615
R99 VTAIL.n39 VTAIL.n37 104.615
R100 VTAIL.n39 VTAIL.n38 104.615
R101 VTAIL.n38 VTAIL.n11 104.615
R102 VTAIL.n47 VTAIL.n11 104.615
R103 VTAIL.n48 VTAIL.n47 104.615
R104 VTAIL.n48 VTAIL.n7 104.615
R105 VTAIL.n55 VTAIL.n7 104.615
R106 VTAIL.n56 VTAIL.n55 104.615
R107 VTAIL.n56 VTAIL.n3 104.615
R108 VTAIL.n63 VTAIL.n3 104.615
R109 VTAIL.n64 VTAIL.n63 104.615
R110 VTAIL.n204 VTAIL.n203 104.615
R111 VTAIL.n203 VTAIL.n143 104.615
R112 VTAIL.n196 VTAIL.n143 104.615
R113 VTAIL.n196 VTAIL.n195 104.615
R114 VTAIL.n195 VTAIL.n147 104.615
R115 VTAIL.n188 VTAIL.n147 104.615
R116 VTAIL.n188 VTAIL.n187 104.615
R117 VTAIL.n187 VTAIL.n151 104.615
R118 VTAIL.n155 VTAIL.n151 104.615
R119 VTAIL.n179 VTAIL.n155 104.615
R120 VTAIL.n179 VTAIL.n178 104.615
R121 VTAIL.n178 VTAIL.n156 104.615
R122 VTAIL.n171 VTAIL.n156 104.615
R123 VTAIL.n171 VTAIL.n170 104.615
R124 VTAIL.n170 VTAIL.n160 104.615
R125 VTAIL.n163 VTAIL.n160 104.615
R126 VTAIL.n134 VTAIL.n133 104.615
R127 VTAIL.n133 VTAIL.n73 104.615
R128 VTAIL.n126 VTAIL.n73 104.615
R129 VTAIL.n126 VTAIL.n125 104.615
R130 VTAIL.n125 VTAIL.n77 104.615
R131 VTAIL.n118 VTAIL.n77 104.615
R132 VTAIL.n118 VTAIL.n117 104.615
R133 VTAIL.n117 VTAIL.n81 104.615
R134 VTAIL.n85 VTAIL.n81 104.615
R135 VTAIL.n109 VTAIL.n85 104.615
R136 VTAIL.n109 VTAIL.n108 104.615
R137 VTAIL.n108 VTAIL.n86 104.615
R138 VTAIL.n101 VTAIL.n86 104.615
R139 VTAIL.n101 VTAIL.n100 104.615
R140 VTAIL.n100 VTAIL.n90 104.615
R141 VTAIL.n93 VTAIL.n90 104.615
R142 VTAIL.n232 VTAIL.t3 52.3082
R143 VTAIL.n22 VTAIL.t1 52.3082
R144 VTAIL.n163 VTAIL.t0 52.3082
R145 VTAIL.n93 VTAIL.t2 52.3082
R146 VTAIL.n279 VTAIL.n278 31.7975
R147 VTAIL.n69 VTAIL.n68 31.7975
R148 VTAIL.n209 VTAIL.n208 31.7975
R149 VTAIL.n139 VTAIL.n138 31.7975
R150 VTAIL.n139 VTAIL.n69 24.7117
R151 VTAIL.n279 VTAIL.n209 24.0738
R152 VTAIL.n256 VTAIL.n255 13.1884
R153 VTAIL.n46 VTAIL.n45 13.1884
R154 VTAIL.n186 VTAIL.n185 13.1884
R155 VTAIL.n116 VTAIL.n115 13.1884
R156 VTAIL.n254 VTAIL.n222 12.8005
R157 VTAIL.n259 VTAIL.n220 12.8005
R158 VTAIL.n44 VTAIL.n12 12.8005
R159 VTAIL.n49 VTAIL.n10 12.8005
R160 VTAIL.n189 VTAIL.n150 12.8005
R161 VTAIL.n184 VTAIL.n152 12.8005
R162 VTAIL.n119 VTAIL.n80 12.8005
R163 VTAIL.n114 VTAIL.n82 12.8005
R164 VTAIL.n251 VTAIL.n250 12.0247
R165 VTAIL.n260 VTAIL.n218 12.0247
R166 VTAIL.n41 VTAIL.n40 12.0247
R167 VTAIL.n50 VTAIL.n8 12.0247
R168 VTAIL.n190 VTAIL.n148 12.0247
R169 VTAIL.n181 VTAIL.n180 12.0247
R170 VTAIL.n120 VTAIL.n78 12.0247
R171 VTAIL.n111 VTAIL.n110 12.0247
R172 VTAIL.n246 VTAIL.n224 11.249
R173 VTAIL.n264 VTAIL.n263 11.249
R174 VTAIL.n36 VTAIL.n14 11.249
R175 VTAIL.n54 VTAIL.n53 11.249
R176 VTAIL.n194 VTAIL.n193 11.249
R177 VTAIL.n177 VTAIL.n154 11.249
R178 VTAIL.n124 VTAIL.n123 11.249
R179 VTAIL.n107 VTAIL.n84 11.249
R180 VTAIL.n245 VTAIL.n226 10.4732
R181 VTAIL.n267 VTAIL.n216 10.4732
R182 VTAIL.n35 VTAIL.n16 10.4732
R183 VTAIL.n57 VTAIL.n6 10.4732
R184 VTAIL.n197 VTAIL.n146 10.4732
R185 VTAIL.n176 VTAIL.n157 10.4732
R186 VTAIL.n127 VTAIL.n76 10.4732
R187 VTAIL.n106 VTAIL.n87 10.4732
R188 VTAIL.n233 VTAIL.n231 10.2747
R189 VTAIL.n23 VTAIL.n21 10.2747
R190 VTAIL.n164 VTAIL.n162 10.2747
R191 VTAIL.n94 VTAIL.n92 10.2747
R192 VTAIL.n242 VTAIL.n241 9.69747
R193 VTAIL.n268 VTAIL.n214 9.69747
R194 VTAIL.n32 VTAIL.n31 9.69747
R195 VTAIL.n58 VTAIL.n4 9.69747
R196 VTAIL.n198 VTAIL.n144 9.69747
R197 VTAIL.n173 VTAIL.n172 9.69747
R198 VTAIL.n128 VTAIL.n74 9.69747
R199 VTAIL.n103 VTAIL.n102 9.69747
R200 VTAIL.n278 VTAIL.n277 9.45567
R201 VTAIL.n68 VTAIL.n67 9.45567
R202 VTAIL.n208 VTAIL.n207 9.45567
R203 VTAIL.n138 VTAIL.n137 9.45567
R204 VTAIL.n212 VTAIL.n211 9.3005
R205 VTAIL.n271 VTAIL.n270 9.3005
R206 VTAIL.n269 VTAIL.n268 9.3005
R207 VTAIL.n216 VTAIL.n215 9.3005
R208 VTAIL.n263 VTAIL.n262 9.3005
R209 VTAIL.n261 VTAIL.n260 9.3005
R210 VTAIL.n220 VTAIL.n219 9.3005
R211 VTAIL.n235 VTAIL.n234 9.3005
R212 VTAIL.n237 VTAIL.n236 9.3005
R213 VTAIL.n228 VTAIL.n227 9.3005
R214 VTAIL.n243 VTAIL.n242 9.3005
R215 VTAIL.n245 VTAIL.n244 9.3005
R216 VTAIL.n224 VTAIL.n223 9.3005
R217 VTAIL.n252 VTAIL.n251 9.3005
R218 VTAIL.n254 VTAIL.n253 9.3005
R219 VTAIL.n277 VTAIL.n276 9.3005
R220 VTAIL.n2 VTAIL.n1 9.3005
R221 VTAIL.n61 VTAIL.n60 9.3005
R222 VTAIL.n59 VTAIL.n58 9.3005
R223 VTAIL.n6 VTAIL.n5 9.3005
R224 VTAIL.n53 VTAIL.n52 9.3005
R225 VTAIL.n51 VTAIL.n50 9.3005
R226 VTAIL.n10 VTAIL.n9 9.3005
R227 VTAIL.n25 VTAIL.n24 9.3005
R228 VTAIL.n27 VTAIL.n26 9.3005
R229 VTAIL.n18 VTAIL.n17 9.3005
R230 VTAIL.n33 VTAIL.n32 9.3005
R231 VTAIL.n35 VTAIL.n34 9.3005
R232 VTAIL.n14 VTAIL.n13 9.3005
R233 VTAIL.n42 VTAIL.n41 9.3005
R234 VTAIL.n44 VTAIL.n43 9.3005
R235 VTAIL.n67 VTAIL.n66 9.3005
R236 VTAIL.n166 VTAIL.n165 9.3005
R237 VTAIL.n168 VTAIL.n167 9.3005
R238 VTAIL.n159 VTAIL.n158 9.3005
R239 VTAIL.n174 VTAIL.n173 9.3005
R240 VTAIL.n176 VTAIL.n175 9.3005
R241 VTAIL.n154 VTAIL.n153 9.3005
R242 VTAIL.n182 VTAIL.n181 9.3005
R243 VTAIL.n184 VTAIL.n183 9.3005
R244 VTAIL.n207 VTAIL.n206 9.3005
R245 VTAIL.n142 VTAIL.n141 9.3005
R246 VTAIL.n201 VTAIL.n200 9.3005
R247 VTAIL.n199 VTAIL.n198 9.3005
R248 VTAIL.n146 VTAIL.n145 9.3005
R249 VTAIL.n193 VTAIL.n192 9.3005
R250 VTAIL.n191 VTAIL.n190 9.3005
R251 VTAIL.n150 VTAIL.n149 9.3005
R252 VTAIL.n96 VTAIL.n95 9.3005
R253 VTAIL.n98 VTAIL.n97 9.3005
R254 VTAIL.n89 VTAIL.n88 9.3005
R255 VTAIL.n104 VTAIL.n103 9.3005
R256 VTAIL.n106 VTAIL.n105 9.3005
R257 VTAIL.n84 VTAIL.n83 9.3005
R258 VTAIL.n112 VTAIL.n111 9.3005
R259 VTAIL.n114 VTAIL.n113 9.3005
R260 VTAIL.n137 VTAIL.n136 9.3005
R261 VTAIL.n72 VTAIL.n71 9.3005
R262 VTAIL.n131 VTAIL.n130 9.3005
R263 VTAIL.n129 VTAIL.n128 9.3005
R264 VTAIL.n76 VTAIL.n75 9.3005
R265 VTAIL.n123 VTAIL.n122 9.3005
R266 VTAIL.n121 VTAIL.n120 9.3005
R267 VTAIL.n80 VTAIL.n79 9.3005
R268 VTAIL.n238 VTAIL.n228 8.92171
R269 VTAIL.n272 VTAIL.n271 8.92171
R270 VTAIL.n28 VTAIL.n18 8.92171
R271 VTAIL.n62 VTAIL.n61 8.92171
R272 VTAIL.n202 VTAIL.n201 8.92171
R273 VTAIL.n169 VTAIL.n159 8.92171
R274 VTAIL.n132 VTAIL.n131 8.92171
R275 VTAIL.n99 VTAIL.n89 8.92171
R276 VTAIL.n237 VTAIL.n230 8.14595
R277 VTAIL.n275 VTAIL.n212 8.14595
R278 VTAIL.n27 VTAIL.n20 8.14595
R279 VTAIL.n65 VTAIL.n2 8.14595
R280 VTAIL.n205 VTAIL.n142 8.14595
R281 VTAIL.n168 VTAIL.n161 8.14595
R282 VTAIL.n135 VTAIL.n72 8.14595
R283 VTAIL.n98 VTAIL.n91 8.14595
R284 VTAIL.n234 VTAIL.n233 7.3702
R285 VTAIL.n276 VTAIL.n210 7.3702
R286 VTAIL.n24 VTAIL.n23 7.3702
R287 VTAIL.n66 VTAIL.n0 7.3702
R288 VTAIL.n206 VTAIL.n140 7.3702
R289 VTAIL.n165 VTAIL.n164 7.3702
R290 VTAIL.n136 VTAIL.n70 7.3702
R291 VTAIL.n95 VTAIL.n94 7.3702
R292 VTAIL.n278 VTAIL.n210 6.59444
R293 VTAIL.n68 VTAIL.n0 6.59444
R294 VTAIL.n208 VTAIL.n140 6.59444
R295 VTAIL.n138 VTAIL.n70 6.59444
R296 VTAIL.n234 VTAIL.n230 5.81868
R297 VTAIL.n276 VTAIL.n275 5.81868
R298 VTAIL.n24 VTAIL.n20 5.81868
R299 VTAIL.n66 VTAIL.n65 5.81868
R300 VTAIL.n206 VTAIL.n205 5.81868
R301 VTAIL.n165 VTAIL.n161 5.81868
R302 VTAIL.n136 VTAIL.n135 5.81868
R303 VTAIL.n95 VTAIL.n91 5.81868
R304 VTAIL.n238 VTAIL.n237 5.04292
R305 VTAIL.n272 VTAIL.n212 5.04292
R306 VTAIL.n28 VTAIL.n27 5.04292
R307 VTAIL.n62 VTAIL.n2 5.04292
R308 VTAIL.n202 VTAIL.n142 5.04292
R309 VTAIL.n169 VTAIL.n168 5.04292
R310 VTAIL.n132 VTAIL.n72 5.04292
R311 VTAIL.n99 VTAIL.n98 5.04292
R312 VTAIL.n241 VTAIL.n228 4.26717
R313 VTAIL.n271 VTAIL.n214 4.26717
R314 VTAIL.n31 VTAIL.n18 4.26717
R315 VTAIL.n61 VTAIL.n4 4.26717
R316 VTAIL.n201 VTAIL.n144 4.26717
R317 VTAIL.n172 VTAIL.n159 4.26717
R318 VTAIL.n131 VTAIL.n74 4.26717
R319 VTAIL.n102 VTAIL.n89 4.26717
R320 VTAIL.n242 VTAIL.n226 3.49141
R321 VTAIL.n268 VTAIL.n267 3.49141
R322 VTAIL.n32 VTAIL.n16 3.49141
R323 VTAIL.n58 VTAIL.n57 3.49141
R324 VTAIL.n198 VTAIL.n197 3.49141
R325 VTAIL.n173 VTAIL.n157 3.49141
R326 VTAIL.n128 VTAIL.n127 3.49141
R327 VTAIL.n103 VTAIL.n87 3.49141
R328 VTAIL.n235 VTAIL.n231 2.84303
R329 VTAIL.n25 VTAIL.n21 2.84303
R330 VTAIL.n166 VTAIL.n162 2.84303
R331 VTAIL.n96 VTAIL.n92 2.84303
R332 VTAIL.n246 VTAIL.n245 2.71565
R333 VTAIL.n264 VTAIL.n216 2.71565
R334 VTAIL.n36 VTAIL.n35 2.71565
R335 VTAIL.n54 VTAIL.n6 2.71565
R336 VTAIL.n194 VTAIL.n146 2.71565
R337 VTAIL.n177 VTAIL.n176 2.71565
R338 VTAIL.n124 VTAIL.n76 2.71565
R339 VTAIL.n107 VTAIL.n106 2.71565
R340 VTAIL.n250 VTAIL.n224 1.93989
R341 VTAIL.n263 VTAIL.n218 1.93989
R342 VTAIL.n40 VTAIL.n14 1.93989
R343 VTAIL.n53 VTAIL.n8 1.93989
R344 VTAIL.n193 VTAIL.n148 1.93989
R345 VTAIL.n180 VTAIL.n154 1.93989
R346 VTAIL.n123 VTAIL.n78 1.93989
R347 VTAIL.n110 VTAIL.n84 1.93989
R348 VTAIL.n251 VTAIL.n222 1.16414
R349 VTAIL.n260 VTAIL.n259 1.16414
R350 VTAIL.n41 VTAIL.n12 1.16414
R351 VTAIL.n50 VTAIL.n49 1.16414
R352 VTAIL.n190 VTAIL.n189 1.16414
R353 VTAIL.n181 VTAIL.n152 1.16414
R354 VTAIL.n120 VTAIL.n119 1.16414
R355 VTAIL.n111 VTAIL.n82 1.16414
R356 VTAIL.n209 VTAIL.n139 0.789293
R357 VTAIL VTAIL.n69 0.688
R358 VTAIL.n255 VTAIL.n254 0.388379
R359 VTAIL.n256 VTAIL.n220 0.388379
R360 VTAIL.n45 VTAIL.n44 0.388379
R361 VTAIL.n46 VTAIL.n10 0.388379
R362 VTAIL.n186 VTAIL.n150 0.388379
R363 VTAIL.n185 VTAIL.n184 0.388379
R364 VTAIL.n116 VTAIL.n80 0.388379
R365 VTAIL.n115 VTAIL.n114 0.388379
R366 VTAIL.n236 VTAIL.n235 0.155672
R367 VTAIL.n236 VTAIL.n227 0.155672
R368 VTAIL.n243 VTAIL.n227 0.155672
R369 VTAIL.n244 VTAIL.n243 0.155672
R370 VTAIL.n244 VTAIL.n223 0.155672
R371 VTAIL.n252 VTAIL.n223 0.155672
R372 VTAIL.n253 VTAIL.n252 0.155672
R373 VTAIL.n253 VTAIL.n219 0.155672
R374 VTAIL.n261 VTAIL.n219 0.155672
R375 VTAIL.n262 VTAIL.n261 0.155672
R376 VTAIL.n262 VTAIL.n215 0.155672
R377 VTAIL.n269 VTAIL.n215 0.155672
R378 VTAIL.n270 VTAIL.n269 0.155672
R379 VTAIL.n270 VTAIL.n211 0.155672
R380 VTAIL.n277 VTAIL.n211 0.155672
R381 VTAIL.n26 VTAIL.n25 0.155672
R382 VTAIL.n26 VTAIL.n17 0.155672
R383 VTAIL.n33 VTAIL.n17 0.155672
R384 VTAIL.n34 VTAIL.n33 0.155672
R385 VTAIL.n34 VTAIL.n13 0.155672
R386 VTAIL.n42 VTAIL.n13 0.155672
R387 VTAIL.n43 VTAIL.n42 0.155672
R388 VTAIL.n43 VTAIL.n9 0.155672
R389 VTAIL.n51 VTAIL.n9 0.155672
R390 VTAIL.n52 VTAIL.n51 0.155672
R391 VTAIL.n52 VTAIL.n5 0.155672
R392 VTAIL.n59 VTAIL.n5 0.155672
R393 VTAIL.n60 VTAIL.n59 0.155672
R394 VTAIL.n60 VTAIL.n1 0.155672
R395 VTAIL.n67 VTAIL.n1 0.155672
R396 VTAIL.n207 VTAIL.n141 0.155672
R397 VTAIL.n200 VTAIL.n141 0.155672
R398 VTAIL.n200 VTAIL.n199 0.155672
R399 VTAIL.n199 VTAIL.n145 0.155672
R400 VTAIL.n192 VTAIL.n145 0.155672
R401 VTAIL.n192 VTAIL.n191 0.155672
R402 VTAIL.n191 VTAIL.n149 0.155672
R403 VTAIL.n183 VTAIL.n149 0.155672
R404 VTAIL.n183 VTAIL.n182 0.155672
R405 VTAIL.n182 VTAIL.n153 0.155672
R406 VTAIL.n175 VTAIL.n153 0.155672
R407 VTAIL.n175 VTAIL.n174 0.155672
R408 VTAIL.n174 VTAIL.n158 0.155672
R409 VTAIL.n167 VTAIL.n158 0.155672
R410 VTAIL.n167 VTAIL.n166 0.155672
R411 VTAIL.n137 VTAIL.n71 0.155672
R412 VTAIL.n130 VTAIL.n71 0.155672
R413 VTAIL.n130 VTAIL.n129 0.155672
R414 VTAIL.n129 VTAIL.n75 0.155672
R415 VTAIL.n122 VTAIL.n75 0.155672
R416 VTAIL.n122 VTAIL.n121 0.155672
R417 VTAIL.n121 VTAIL.n79 0.155672
R418 VTAIL.n113 VTAIL.n79 0.155672
R419 VTAIL.n113 VTAIL.n112 0.155672
R420 VTAIL.n112 VTAIL.n83 0.155672
R421 VTAIL.n105 VTAIL.n83 0.155672
R422 VTAIL.n105 VTAIL.n104 0.155672
R423 VTAIL.n104 VTAIL.n88 0.155672
R424 VTAIL.n97 VTAIL.n88 0.155672
R425 VTAIL.n97 VTAIL.n96 0.155672
R426 VTAIL VTAIL.n279 0.101793
R427 VDD2.n133 VDD2.n69 289.615
R428 VDD2.n64 VDD2.n0 289.615
R429 VDD2.n134 VDD2.n133 185
R430 VDD2.n132 VDD2.n131 185
R431 VDD2.n73 VDD2.n72 185
R432 VDD2.n126 VDD2.n125 185
R433 VDD2.n124 VDD2.n123 185
R434 VDD2.n77 VDD2.n76 185
R435 VDD2.n118 VDD2.n117 185
R436 VDD2.n116 VDD2.n115 185
R437 VDD2.n114 VDD2.n80 185
R438 VDD2.n84 VDD2.n81 185
R439 VDD2.n109 VDD2.n108 185
R440 VDD2.n107 VDD2.n106 185
R441 VDD2.n86 VDD2.n85 185
R442 VDD2.n101 VDD2.n100 185
R443 VDD2.n99 VDD2.n98 185
R444 VDD2.n90 VDD2.n89 185
R445 VDD2.n93 VDD2.n92 185
R446 VDD2.n23 VDD2.n22 185
R447 VDD2.n20 VDD2.n19 185
R448 VDD2.n29 VDD2.n28 185
R449 VDD2.n31 VDD2.n30 185
R450 VDD2.n16 VDD2.n15 185
R451 VDD2.n37 VDD2.n36 185
R452 VDD2.n40 VDD2.n39 185
R453 VDD2.n38 VDD2.n12 185
R454 VDD2.n45 VDD2.n11 185
R455 VDD2.n47 VDD2.n46 185
R456 VDD2.n49 VDD2.n48 185
R457 VDD2.n8 VDD2.n7 185
R458 VDD2.n55 VDD2.n54 185
R459 VDD2.n57 VDD2.n56 185
R460 VDD2.n4 VDD2.n3 185
R461 VDD2.n63 VDD2.n62 185
R462 VDD2.n65 VDD2.n64 185
R463 VDD2.t1 VDD2.n91 149.524
R464 VDD2.t0 VDD2.n21 149.524
R465 VDD2.n133 VDD2.n132 104.615
R466 VDD2.n132 VDD2.n72 104.615
R467 VDD2.n125 VDD2.n72 104.615
R468 VDD2.n125 VDD2.n124 104.615
R469 VDD2.n124 VDD2.n76 104.615
R470 VDD2.n117 VDD2.n76 104.615
R471 VDD2.n117 VDD2.n116 104.615
R472 VDD2.n116 VDD2.n80 104.615
R473 VDD2.n84 VDD2.n80 104.615
R474 VDD2.n108 VDD2.n84 104.615
R475 VDD2.n108 VDD2.n107 104.615
R476 VDD2.n107 VDD2.n85 104.615
R477 VDD2.n100 VDD2.n85 104.615
R478 VDD2.n100 VDD2.n99 104.615
R479 VDD2.n99 VDD2.n89 104.615
R480 VDD2.n92 VDD2.n89 104.615
R481 VDD2.n22 VDD2.n19 104.615
R482 VDD2.n29 VDD2.n19 104.615
R483 VDD2.n30 VDD2.n29 104.615
R484 VDD2.n30 VDD2.n15 104.615
R485 VDD2.n37 VDD2.n15 104.615
R486 VDD2.n39 VDD2.n37 104.615
R487 VDD2.n39 VDD2.n38 104.615
R488 VDD2.n38 VDD2.n11 104.615
R489 VDD2.n47 VDD2.n11 104.615
R490 VDD2.n48 VDD2.n47 104.615
R491 VDD2.n48 VDD2.n7 104.615
R492 VDD2.n55 VDD2.n7 104.615
R493 VDD2.n56 VDD2.n55 104.615
R494 VDD2.n56 VDD2.n3 104.615
R495 VDD2.n63 VDD2.n3 104.615
R496 VDD2.n64 VDD2.n63 104.615
R497 VDD2.n138 VDD2.n68 84.4805
R498 VDD2.n92 VDD2.t1 52.3082
R499 VDD2.n22 VDD2.t0 52.3082
R500 VDD2.n138 VDD2.n137 48.4763
R501 VDD2.n115 VDD2.n114 13.1884
R502 VDD2.n46 VDD2.n45 13.1884
R503 VDD2.n118 VDD2.n79 12.8005
R504 VDD2.n113 VDD2.n81 12.8005
R505 VDD2.n44 VDD2.n12 12.8005
R506 VDD2.n49 VDD2.n10 12.8005
R507 VDD2.n119 VDD2.n77 12.0247
R508 VDD2.n110 VDD2.n109 12.0247
R509 VDD2.n41 VDD2.n40 12.0247
R510 VDD2.n50 VDD2.n8 12.0247
R511 VDD2.n123 VDD2.n122 11.249
R512 VDD2.n106 VDD2.n83 11.249
R513 VDD2.n36 VDD2.n14 11.249
R514 VDD2.n54 VDD2.n53 11.249
R515 VDD2.n126 VDD2.n75 10.4732
R516 VDD2.n105 VDD2.n86 10.4732
R517 VDD2.n35 VDD2.n16 10.4732
R518 VDD2.n57 VDD2.n6 10.4732
R519 VDD2.n93 VDD2.n91 10.2747
R520 VDD2.n23 VDD2.n21 10.2747
R521 VDD2.n127 VDD2.n73 9.69747
R522 VDD2.n102 VDD2.n101 9.69747
R523 VDD2.n32 VDD2.n31 9.69747
R524 VDD2.n58 VDD2.n4 9.69747
R525 VDD2.n137 VDD2.n136 9.45567
R526 VDD2.n68 VDD2.n67 9.45567
R527 VDD2.n95 VDD2.n94 9.3005
R528 VDD2.n97 VDD2.n96 9.3005
R529 VDD2.n88 VDD2.n87 9.3005
R530 VDD2.n103 VDD2.n102 9.3005
R531 VDD2.n105 VDD2.n104 9.3005
R532 VDD2.n83 VDD2.n82 9.3005
R533 VDD2.n111 VDD2.n110 9.3005
R534 VDD2.n113 VDD2.n112 9.3005
R535 VDD2.n136 VDD2.n135 9.3005
R536 VDD2.n71 VDD2.n70 9.3005
R537 VDD2.n130 VDD2.n129 9.3005
R538 VDD2.n128 VDD2.n127 9.3005
R539 VDD2.n75 VDD2.n74 9.3005
R540 VDD2.n122 VDD2.n121 9.3005
R541 VDD2.n120 VDD2.n119 9.3005
R542 VDD2.n79 VDD2.n78 9.3005
R543 VDD2.n2 VDD2.n1 9.3005
R544 VDD2.n61 VDD2.n60 9.3005
R545 VDD2.n59 VDD2.n58 9.3005
R546 VDD2.n6 VDD2.n5 9.3005
R547 VDD2.n53 VDD2.n52 9.3005
R548 VDD2.n51 VDD2.n50 9.3005
R549 VDD2.n10 VDD2.n9 9.3005
R550 VDD2.n25 VDD2.n24 9.3005
R551 VDD2.n27 VDD2.n26 9.3005
R552 VDD2.n18 VDD2.n17 9.3005
R553 VDD2.n33 VDD2.n32 9.3005
R554 VDD2.n35 VDD2.n34 9.3005
R555 VDD2.n14 VDD2.n13 9.3005
R556 VDD2.n42 VDD2.n41 9.3005
R557 VDD2.n44 VDD2.n43 9.3005
R558 VDD2.n67 VDD2.n66 9.3005
R559 VDD2.n131 VDD2.n130 8.92171
R560 VDD2.n98 VDD2.n88 8.92171
R561 VDD2.n28 VDD2.n18 8.92171
R562 VDD2.n62 VDD2.n61 8.92171
R563 VDD2.n134 VDD2.n71 8.14595
R564 VDD2.n97 VDD2.n90 8.14595
R565 VDD2.n27 VDD2.n20 8.14595
R566 VDD2.n65 VDD2.n2 8.14595
R567 VDD2.n135 VDD2.n69 7.3702
R568 VDD2.n94 VDD2.n93 7.3702
R569 VDD2.n24 VDD2.n23 7.3702
R570 VDD2.n66 VDD2.n0 7.3702
R571 VDD2.n137 VDD2.n69 6.59444
R572 VDD2.n68 VDD2.n0 6.59444
R573 VDD2.n135 VDD2.n134 5.81868
R574 VDD2.n94 VDD2.n90 5.81868
R575 VDD2.n24 VDD2.n20 5.81868
R576 VDD2.n66 VDD2.n65 5.81868
R577 VDD2.n131 VDD2.n71 5.04292
R578 VDD2.n98 VDD2.n97 5.04292
R579 VDD2.n28 VDD2.n27 5.04292
R580 VDD2.n62 VDD2.n2 5.04292
R581 VDD2.n130 VDD2.n73 4.26717
R582 VDD2.n101 VDD2.n88 4.26717
R583 VDD2.n31 VDD2.n18 4.26717
R584 VDD2.n61 VDD2.n4 4.26717
R585 VDD2.n127 VDD2.n126 3.49141
R586 VDD2.n102 VDD2.n86 3.49141
R587 VDD2.n32 VDD2.n16 3.49141
R588 VDD2.n58 VDD2.n57 3.49141
R589 VDD2.n95 VDD2.n91 2.84303
R590 VDD2.n25 VDD2.n21 2.84303
R591 VDD2.n123 VDD2.n75 2.71565
R592 VDD2.n106 VDD2.n105 2.71565
R593 VDD2.n36 VDD2.n35 2.71565
R594 VDD2.n54 VDD2.n6 2.71565
R595 VDD2.n122 VDD2.n77 1.93989
R596 VDD2.n109 VDD2.n83 1.93989
R597 VDD2.n40 VDD2.n14 1.93989
R598 VDD2.n53 VDD2.n8 1.93989
R599 VDD2.n119 VDD2.n118 1.16414
R600 VDD2.n110 VDD2.n81 1.16414
R601 VDD2.n41 VDD2.n12 1.16414
R602 VDD2.n50 VDD2.n49 1.16414
R603 VDD2.n115 VDD2.n79 0.388379
R604 VDD2.n114 VDD2.n113 0.388379
R605 VDD2.n45 VDD2.n44 0.388379
R606 VDD2.n46 VDD2.n10 0.388379
R607 VDD2 VDD2.n138 0.218172
R608 VDD2.n136 VDD2.n70 0.155672
R609 VDD2.n129 VDD2.n70 0.155672
R610 VDD2.n129 VDD2.n128 0.155672
R611 VDD2.n128 VDD2.n74 0.155672
R612 VDD2.n121 VDD2.n74 0.155672
R613 VDD2.n121 VDD2.n120 0.155672
R614 VDD2.n120 VDD2.n78 0.155672
R615 VDD2.n112 VDD2.n78 0.155672
R616 VDD2.n112 VDD2.n111 0.155672
R617 VDD2.n111 VDD2.n82 0.155672
R618 VDD2.n104 VDD2.n82 0.155672
R619 VDD2.n104 VDD2.n103 0.155672
R620 VDD2.n103 VDD2.n87 0.155672
R621 VDD2.n96 VDD2.n87 0.155672
R622 VDD2.n96 VDD2.n95 0.155672
R623 VDD2.n26 VDD2.n25 0.155672
R624 VDD2.n26 VDD2.n17 0.155672
R625 VDD2.n33 VDD2.n17 0.155672
R626 VDD2.n34 VDD2.n33 0.155672
R627 VDD2.n34 VDD2.n13 0.155672
R628 VDD2.n42 VDD2.n13 0.155672
R629 VDD2.n43 VDD2.n42 0.155672
R630 VDD2.n43 VDD2.n9 0.155672
R631 VDD2.n51 VDD2.n9 0.155672
R632 VDD2.n52 VDD2.n51 0.155672
R633 VDD2.n52 VDD2.n5 0.155672
R634 VDD2.n59 VDD2.n5 0.155672
R635 VDD2.n60 VDD2.n59 0.155672
R636 VDD2.n60 VDD2.n1 0.155672
R637 VDD2.n67 VDD2.n1 0.155672
R638 B.n80 B.t9 962.62
R639 B.n77 B.t13 962.62
R640 B.n452 B.t6 962.62
R641 B.n324 B.t2 962.62
R642 B.n601 B.n600 585
R643 B.n273 B.n76 585
R644 B.n272 B.n271 585
R645 B.n270 B.n269 585
R646 B.n268 B.n267 585
R647 B.n266 B.n265 585
R648 B.n264 B.n263 585
R649 B.n262 B.n261 585
R650 B.n260 B.n259 585
R651 B.n258 B.n257 585
R652 B.n256 B.n255 585
R653 B.n254 B.n253 585
R654 B.n252 B.n251 585
R655 B.n250 B.n249 585
R656 B.n248 B.n247 585
R657 B.n246 B.n245 585
R658 B.n244 B.n243 585
R659 B.n242 B.n241 585
R660 B.n240 B.n239 585
R661 B.n238 B.n237 585
R662 B.n236 B.n235 585
R663 B.n234 B.n233 585
R664 B.n232 B.n231 585
R665 B.n230 B.n229 585
R666 B.n228 B.n227 585
R667 B.n226 B.n225 585
R668 B.n224 B.n223 585
R669 B.n222 B.n221 585
R670 B.n220 B.n219 585
R671 B.n218 B.n217 585
R672 B.n216 B.n215 585
R673 B.n214 B.n213 585
R674 B.n212 B.n211 585
R675 B.n210 B.n209 585
R676 B.n208 B.n207 585
R677 B.n206 B.n205 585
R678 B.n204 B.n203 585
R679 B.n202 B.n201 585
R680 B.n200 B.n199 585
R681 B.n198 B.n197 585
R682 B.n196 B.n195 585
R683 B.n194 B.n193 585
R684 B.n192 B.n191 585
R685 B.n190 B.n189 585
R686 B.n188 B.n187 585
R687 B.n186 B.n185 585
R688 B.n184 B.n183 585
R689 B.n182 B.n181 585
R690 B.n180 B.n179 585
R691 B.n178 B.n177 585
R692 B.n176 B.n175 585
R693 B.n174 B.n173 585
R694 B.n172 B.n171 585
R695 B.n170 B.n169 585
R696 B.n168 B.n167 585
R697 B.n166 B.n165 585
R698 B.n164 B.n163 585
R699 B.n162 B.n161 585
R700 B.n160 B.n159 585
R701 B.n158 B.n157 585
R702 B.n156 B.n155 585
R703 B.n154 B.n153 585
R704 B.n152 B.n151 585
R705 B.n150 B.n149 585
R706 B.n148 B.n147 585
R707 B.n146 B.n145 585
R708 B.n144 B.n143 585
R709 B.n142 B.n141 585
R710 B.n140 B.n139 585
R711 B.n138 B.n137 585
R712 B.n136 B.n135 585
R713 B.n134 B.n133 585
R714 B.n132 B.n131 585
R715 B.n130 B.n129 585
R716 B.n128 B.n127 585
R717 B.n126 B.n125 585
R718 B.n124 B.n123 585
R719 B.n122 B.n121 585
R720 B.n120 B.n119 585
R721 B.n118 B.n117 585
R722 B.n116 B.n115 585
R723 B.n114 B.n113 585
R724 B.n112 B.n111 585
R725 B.n110 B.n109 585
R726 B.n108 B.n107 585
R727 B.n106 B.n105 585
R728 B.n104 B.n103 585
R729 B.n102 B.n101 585
R730 B.n100 B.n99 585
R731 B.n98 B.n97 585
R732 B.n96 B.n95 585
R733 B.n94 B.n93 585
R734 B.n92 B.n91 585
R735 B.n90 B.n89 585
R736 B.n88 B.n87 585
R737 B.n86 B.n85 585
R738 B.n84 B.n83 585
R739 B.n26 B.n25 585
R740 B.n599 B.n27 585
R741 B.n604 B.n27 585
R742 B.n598 B.n597 585
R743 B.n597 B.n23 585
R744 B.n596 B.n22 585
R745 B.n610 B.n22 585
R746 B.n595 B.n21 585
R747 B.n611 B.n21 585
R748 B.n594 B.n20 585
R749 B.n612 B.n20 585
R750 B.n593 B.n592 585
R751 B.n592 B.n16 585
R752 B.n591 B.n15 585
R753 B.n618 B.n15 585
R754 B.n590 B.n14 585
R755 B.n619 B.n14 585
R756 B.n589 B.n13 585
R757 B.n620 B.n13 585
R758 B.n588 B.n587 585
R759 B.n587 B.n12 585
R760 B.n586 B.n585 585
R761 B.n586 B.n8 585
R762 B.n584 B.n7 585
R763 B.n627 B.n7 585
R764 B.n583 B.n6 585
R765 B.n628 B.n6 585
R766 B.n582 B.n5 585
R767 B.n629 B.n5 585
R768 B.n581 B.n580 585
R769 B.n580 B.n4 585
R770 B.n579 B.n274 585
R771 B.n579 B.n578 585
R772 B.n568 B.n275 585
R773 B.n571 B.n275 585
R774 B.n570 B.n569 585
R775 B.n572 B.n570 585
R776 B.n567 B.n280 585
R777 B.n280 B.n279 585
R778 B.n566 B.n565 585
R779 B.n565 B.n564 585
R780 B.n282 B.n281 585
R781 B.n283 B.n282 585
R782 B.n557 B.n556 585
R783 B.n558 B.n557 585
R784 B.n555 B.n288 585
R785 B.n288 B.n287 585
R786 B.n554 B.n553 585
R787 B.n553 B.n552 585
R788 B.n290 B.n289 585
R789 B.n291 B.n290 585
R790 B.n545 B.n544 585
R791 B.n546 B.n545 585
R792 B.n294 B.n293 585
R793 B.n349 B.n347 585
R794 B.n350 B.n346 585
R795 B.n350 B.n295 585
R796 B.n353 B.n352 585
R797 B.n354 B.n345 585
R798 B.n356 B.n355 585
R799 B.n358 B.n344 585
R800 B.n361 B.n360 585
R801 B.n362 B.n343 585
R802 B.n364 B.n363 585
R803 B.n366 B.n342 585
R804 B.n369 B.n368 585
R805 B.n370 B.n341 585
R806 B.n372 B.n371 585
R807 B.n374 B.n340 585
R808 B.n377 B.n376 585
R809 B.n378 B.n339 585
R810 B.n380 B.n379 585
R811 B.n382 B.n338 585
R812 B.n385 B.n384 585
R813 B.n386 B.n337 585
R814 B.n388 B.n387 585
R815 B.n390 B.n336 585
R816 B.n393 B.n392 585
R817 B.n394 B.n335 585
R818 B.n396 B.n395 585
R819 B.n398 B.n334 585
R820 B.n401 B.n400 585
R821 B.n402 B.n333 585
R822 B.n404 B.n403 585
R823 B.n406 B.n332 585
R824 B.n409 B.n408 585
R825 B.n410 B.n331 585
R826 B.n412 B.n411 585
R827 B.n414 B.n330 585
R828 B.n417 B.n416 585
R829 B.n418 B.n329 585
R830 B.n420 B.n419 585
R831 B.n422 B.n328 585
R832 B.n425 B.n424 585
R833 B.n426 B.n327 585
R834 B.n428 B.n427 585
R835 B.n430 B.n326 585
R836 B.n433 B.n432 585
R837 B.n435 B.n323 585
R838 B.n437 B.n436 585
R839 B.n439 B.n322 585
R840 B.n442 B.n441 585
R841 B.n443 B.n321 585
R842 B.n445 B.n444 585
R843 B.n447 B.n320 585
R844 B.n450 B.n449 585
R845 B.n451 B.n319 585
R846 B.n456 B.n455 585
R847 B.n458 B.n318 585
R848 B.n461 B.n460 585
R849 B.n462 B.n317 585
R850 B.n464 B.n463 585
R851 B.n466 B.n316 585
R852 B.n469 B.n468 585
R853 B.n470 B.n315 585
R854 B.n472 B.n471 585
R855 B.n474 B.n314 585
R856 B.n477 B.n476 585
R857 B.n478 B.n313 585
R858 B.n480 B.n479 585
R859 B.n482 B.n312 585
R860 B.n485 B.n484 585
R861 B.n486 B.n311 585
R862 B.n488 B.n487 585
R863 B.n490 B.n310 585
R864 B.n493 B.n492 585
R865 B.n494 B.n309 585
R866 B.n496 B.n495 585
R867 B.n498 B.n308 585
R868 B.n501 B.n500 585
R869 B.n502 B.n307 585
R870 B.n504 B.n503 585
R871 B.n506 B.n306 585
R872 B.n509 B.n508 585
R873 B.n510 B.n305 585
R874 B.n512 B.n511 585
R875 B.n514 B.n304 585
R876 B.n517 B.n516 585
R877 B.n518 B.n303 585
R878 B.n520 B.n519 585
R879 B.n522 B.n302 585
R880 B.n525 B.n524 585
R881 B.n526 B.n301 585
R882 B.n528 B.n527 585
R883 B.n530 B.n300 585
R884 B.n533 B.n532 585
R885 B.n534 B.n299 585
R886 B.n536 B.n535 585
R887 B.n538 B.n298 585
R888 B.n539 B.n297 585
R889 B.n542 B.n541 585
R890 B.n543 B.n296 585
R891 B.n296 B.n295 585
R892 B.n548 B.n547 585
R893 B.n547 B.n546 585
R894 B.n549 B.n292 585
R895 B.n292 B.n291 585
R896 B.n551 B.n550 585
R897 B.n552 B.n551 585
R898 B.n286 B.n285 585
R899 B.n287 B.n286 585
R900 B.n560 B.n559 585
R901 B.n559 B.n558 585
R902 B.n561 B.n284 585
R903 B.n284 B.n283 585
R904 B.n563 B.n562 585
R905 B.n564 B.n563 585
R906 B.n278 B.n277 585
R907 B.n279 B.n278 585
R908 B.n574 B.n573 585
R909 B.n573 B.n572 585
R910 B.n575 B.n276 585
R911 B.n571 B.n276 585
R912 B.n577 B.n576 585
R913 B.n578 B.n577 585
R914 B.n3 B.n0 585
R915 B.n4 B.n3 585
R916 B.n626 B.n1 585
R917 B.n627 B.n626 585
R918 B.n625 B.n624 585
R919 B.n625 B.n8 585
R920 B.n623 B.n9 585
R921 B.n12 B.n9 585
R922 B.n622 B.n621 585
R923 B.n621 B.n620 585
R924 B.n11 B.n10 585
R925 B.n619 B.n11 585
R926 B.n617 B.n616 585
R927 B.n618 B.n617 585
R928 B.n615 B.n17 585
R929 B.n17 B.n16 585
R930 B.n614 B.n613 585
R931 B.n613 B.n612 585
R932 B.n19 B.n18 585
R933 B.n611 B.n19 585
R934 B.n609 B.n608 585
R935 B.n610 B.n609 585
R936 B.n607 B.n24 585
R937 B.n24 B.n23 585
R938 B.n606 B.n605 585
R939 B.n605 B.n604 585
R940 B.n630 B.n629 585
R941 B.n628 B.n2 585
R942 B.n605 B.n26 473.281
R943 B.n601 B.n27 473.281
R944 B.n545 B.n296 473.281
R945 B.n547 B.n294 473.281
R946 B.n77 B.t14 310.788
R947 B.n452 B.t8 310.788
R948 B.n80 B.t11 310.788
R949 B.n324 B.t5 310.788
R950 B.n78 B.t15 296.435
R951 B.n453 B.t7 296.435
R952 B.n81 B.t12 296.435
R953 B.n325 B.t4 296.435
R954 B.n603 B.n602 256.663
R955 B.n603 B.n75 256.663
R956 B.n603 B.n74 256.663
R957 B.n603 B.n73 256.663
R958 B.n603 B.n72 256.663
R959 B.n603 B.n71 256.663
R960 B.n603 B.n70 256.663
R961 B.n603 B.n69 256.663
R962 B.n603 B.n68 256.663
R963 B.n603 B.n67 256.663
R964 B.n603 B.n66 256.663
R965 B.n603 B.n65 256.663
R966 B.n603 B.n64 256.663
R967 B.n603 B.n63 256.663
R968 B.n603 B.n62 256.663
R969 B.n603 B.n61 256.663
R970 B.n603 B.n60 256.663
R971 B.n603 B.n59 256.663
R972 B.n603 B.n58 256.663
R973 B.n603 B.n57 256.663
R974 B.n603 B.n56 256.663
R975 B.n603 B.n55 256.663
R976 B.n603 B.n54 256.663
R977 B.n603 B.n53 256.663
R978 B.n603 B.n52 256.663
R979 B.n603 B.n51 256.663
R980 B.n603 B.n50 256.663
R981 B.n603 B.n49 256.663
R982 B.n603 B.n48 256.663
R983 B.n603 B.n47 256.663
R984 B.n603 B.n46 256.663
R985 B.n603 B.n45 256.663
R986 B.n603 B.n44 256.663
R987 B.n603 B.n43 256.663
R988 B.n603 B.n42 256.663
R989 B.n603 B.n41 256.663
R990 B.n603 B.n40 256.663
R991 B.n603 B.n39 256.663
R992 B.n603 B.n38 256.663
R993 B.n603 B.n37 256.663
R994 B.n603 B.n36 256.663
R995 B.n603 B.n35 256.663
R996 B.n603 B.n34 256.663
R997 B.n603 B.n33 256.663
R998 B.n603 B.n32 256.663
R999 B.n603 B.n31 256.663
R1000 B.n603 B.n30 256.663
R1001 B.n603 B.n29 256.663
R1002 B.n603 B.n28 256.663
R1003 B.n348 B.n295 256.663
R1004 B.n351 B.n295 256.663
R1005 B.n357 B.n295 256.663
R1006 B.n359 B.n295 256.663
R1007 B.n365 B.n295 256.663
R1008 B.n367 B.n295 256.663
R1009 B.n373 B.n295 256.663
R1010 B.n375 B.n295 256.663
R1011 B.n381 B.n295 256.663
R1012 B.n383 B.n295 256.663
R1013 B.n389 B.n295 256.663
R1014 B.n391 B.n295 256.663
R1015 B.n397 B.n295 256.663
R1016 B.n399 B.n295 256.663
R1017 B.n405 B.n295 256.663
R1018 B.n407 B.n295 256.663
R1019 B.n413 B.n295 256.663
R1020 B.n415 B.n295 256.663
R1021 B.n421 B.n295 256.663
R1022 B.n423 B.n295 256.663
R1023 B.n429 B.n295 256.663
R1024 B.n431 B.n295 256.663
R1025 B.n438 B.n295 256.663
R1026 B.n440 B.n295 256.663
R1027 B.n446 B.n295 256.663
R1028 B.n448 B.n295 256.663
R1029 B.n457 B.n295 256.663
R1030 B.n459 B.n295 256.663
R1031 B.n465 B.n295 256.663
R1032 B.n467 B.n295 256.663
R1033 B.n473 B.n295 256.663
R1034 B.n475 B.n295 256.663
R1035 B.n481 B.n295 256.663
R1036 B.n483 B.n295 256.663
R1037 B.n489 B.n295 256.663
R1038 B.n491 B.n295 256.663
R1039 B.n497 B.n295 256.663
R1040 B.n499 B.n295 256.663
R1041 B.n505 B.n295 256.663
R1042 B.n507 B.n295 256.663
R1043 B.n513 B.n295 256.663
R1044 B.n515 B.n295 256.663
R1045 B.n521 B.n295 256.663
R1046 B.n523 B.n295 256.663
R1047 B.n529 B.n295 256.663
R1048 B.n531 B.n295 256.663
R1049 B.n537 B.n295 256.663
R1050 B.n540 B.n295 256.663
R1051 B.n632 B.n631 256.663
R1052 B.n85 B.n84 163.367
R1053 B.n89 B.n88 163.367
R1054 B.n93 B.n92 163.367
R1055 B.n97 B.n96 163.367
R1056 B.n101 B.n100 163.367
R1057 B.n105 B.n104 163.367
R1058 B.n109 B.n108 163.367
R1059 B.n113 B.n112 163.367
R1060 B.n117 B.n116 163.367
R1061 B.n121 B.n120 163.367
R1062 B.n125 B.n124 163.367
R1063 B.n129 B.n128 163.367
R1064 B.n133 B.n132 163.367
R1065 B.n137 B.n136 163.367
R1066 B.n141 B.n140 163.367
R1067 B.n145 B.n144 163.367
R1068 B.n149 B.n148 163.367
R1069 B.n153 B.n152 163.367
R1070 B.n157 B.n156 163.367
R1071 B.n161 B.n160 163.367
R1072 B.n165 B.n164 163.367
R1073 B.n169 B.n168 163.367
R1074 B.n173 B.n172 163.367
R1075 B.n177 B.n176 163.367
R1076 B.n181 B.n180 163.367
R1077 B.n185 B.n184 163.367
R1078 B.n189 B.n188 163.367
R1079 B.n193 B.n192 163.367
R1080 B.n197 B.n196 163.367
R1081 B.n201 B.n200 163.367
R1082 B.n205 B.n204 163.367
R1083 B.n209 B.n208 163.367
R1084 B.n213 B.n212 163.367
R1085 B.n217 B.n216 163.367
R1086 B.n221 B.n220 163.367
R1087 B.n225 B.n224 163.367
R1088 B.n229 B.n228 163.367
R1089 B.n233 B.n232 163.367
R1090 B.n237 B.n236 163.367
R1091 B.n241 B.n240 163.367
R1092 B.n245 B.n244 163.367
R1093 B.n249 B.n248 163.367
R1094 B.n253 B.n252 163.367
R1095 B.n257 B.n256 163.367
R1096 B.n261 B.n260 163.367
R1097 B.n265 B.n264 163.367
R1098 B.n269 B.n268 163.367
R1099 B.n271 B.n76 163.367
R1100 B.n545 B.n290 163.367
R1101 B.n553 B.n290 163.367
R1102 B.n553 B.n288 163.367
R1103 B.n557 B.n288 163.367
R1104 B.n557 B.n282 163.367
R1105 B.n565 B.n282 163.367
R1106 B.n565 B.n280 163.367
R1107 B.n570 B.n280 163.367
R1108 B.n570 B.n275 163.367
R1109 B.n579 B.n275 163.367
R1110 B.n580 B.n579 163.367
R1111 B.n580 B.n5 163.367
R1112 B.n6 B.n5 163.367
R1113 B.n7 B.n6 163.367
R1114 B.n586 B.n7 163.367
R1115 B.n587 B.n586 163.367
R1116 B.n587 B.n13 163.367
R1117 B.n14 B.n13 163.367
R1118 B.n15 B.n14 163.367
R1119 B.n592 B.n15 163.367
R1120 B.n592 B.n20 163.367
R1121 B.n21 B.n20 163.367
R1122 B.n22 B.n21 163.367
R1123 B.n597 B.n22 163.367
R1124 B.n597 B.n27 163.367
R1125 B.n350 B.n349 163.367
R1126 B.n352 B.n350 163.367
R1127 B.n356 B.n345 163.367
R1128 B.n360 B.n358 163.367
R1129 B.n364 B.n343 163.367
R1130 B.n368 B.n366 163.367
R1131 B.n372 B.n341 163.367
R1132 B.n376 B.n374 163.367
R1133 B.n380 B.n339 163.367
R1134 B.n384 B.n382 163.367
R1135 B.n388 B.n337 163.367
R1136 B.n392 B.n390 163.367
R1137 B.n396 B.n335 163.367
R1138 B.n400 B.n398 163.367
R1139 B.n404 B.n333 163.367
R1140 B.n408 B.n406 163.367
R1141 B.n412 B.n331 163.367
R1142 B.n416 B.n414 163.367
R1143 B.n420 B.n329 163.367
R1144 B.n424 B.n422 163.367
R1145 B.n428 B.n327 163.367
R1146 B.n432 B.n430 163.367
R1147 B.n437 B.n323 163.367
R1148 B.n441 B.n439 163.367
R1149 B.n445 B.n321 163.367
R1150 B.n449 B.n447 163.367
R1151 B.n456 B.n319 163.367
R1152 B.n460 B.n458 163.367
R1153 B.n464 B.n317 163.367
R1154 B.n468 B.n466 163.367
R1155 B.n472 B.n315 163.367
R1156 B.n476 B.n474 163.367
R1157 B.n480 B.n313 163.367
R1158 B.n484 B.n482 163.367
R1159 B.n488 B.n311 163.367
R1160 B.n492 B.n490 163.367
R1161 B.n496 B.n309 163.367
R1162 B.n500 B.n498 163.367
R1163 B.n504 B.n307 163.367
R1164 B.n508 B.n506 163.367
R1165 B.n512 B.n305 163.367
R1166 B.n516 B.n514 163.367
R1167 B.n520 B.n303 163.367
R1168 B.n524 B.n522 163.367
R1169 B.n528 B.n301 163.367
R1170 B.n532 B.n530 163.367
R1171 B.n536 B.n299 163.367
R1172 B.n539 B.n538 163.367
R1173 B.n541 B.n296 163.367
R1174 B.n547 B.n292 163.367
R1175 B.n551 B.n292 163.367
R1176 B.n551 B.n286 163.367
R1177 B.n559 B.n286 163.367
R1178 B.n559 B.n284 163.367
R1179 B.n563 B.n284 163.367
R1180 B.n563 B.n278 163.367
R1181 B.n573 B.n278 163.367
R1182 B.n573 B.n276 163.367
R1183 B.n577 B.n276 163.367
R1184 B.n577 B.n3 163.367
R1185 B.n630 B.n3 163.367
R1186 B.n626 B.n2 163.367
R1187 B.n626 B.n625 163.367
R1188 B.n625 B.n9 163.367
R1189 B.n621 B.n9 163.367
R1190 B.n621 B.n11 163.367
R1191 B.n617 B.n11 163.367
R1192 B.n617 B.n17 163.367
R1193 B.n613 B.n17 163.367
R1194 B.n613 B.n19 163.367
R1195 B.n609 B.n19 163.367
R1196 B.n609 B.n24 163.367
R1197 B.n605 B.n24 163.367
R1198 B.n546 B.n295 73.4755
R1199 B.n604 B.n603 73.4755
R1200 B.n28 B.n26 71.676
R1201 B.n85 B.n29 71.676
R1202 B.n89 B.n30 71.676
R1203 B.n93 B.n31 71.676
R1204 B.n97 B.n32 71.676
R1205 B.n101 B.n33 71.676
R1206 B.n105 B.n34 71.676
R1207 B.n109 B.n35 71.676
R1208 B.n113 B.n36 71.676
R1209 B.n117 B.n37 71.676
R1210 B.n121 B.n38 71.676
R1211 B.n125 B.n39 71.676
R1212 B.n129 B.n40 71.676
R1213 B.n133 B.n41 71.676
R1214 B.n137 B.n42 71.676
R1215 B.n141 B.n43 71.676
R1216 B.n145 B.n44 71.676
R1217 B.n149 B.n45 71.676
R1218 B.n153 B.n46 71.676
R1219 B.n157 B.n47 71.676
R1220 B.n161 B.n48 71.676
R1221 B.n165 B.n49 71.676
R1222 B.n169 B.n50 71.676
R1223 B.n173 B.n51 71.676
R1224 B.n177 B.n52 71.676
R1225 B.n181 B.n53 71.676
R1226 B.n185 B.n54 71.676
R1227 B.n189 B.n55 71.676
R1228 B.n193 B.n56 71.676
R1229 B.n197 B.n57 71.676
R1230 B.n201 B.n58 71.676
R1231 B.n205 B.n59 71.676
R1232 B.n209 B.n60 71.676
R1233 B.n213 B.n61 71.676
R1234 B.n217 B.n62 71.676
R1235 B.n221 B.n63 71.676
R1236 B.n225 B.n64 71.676
R1237 B.n229 B.n65 71.676
R1238 B.n233 B.n66 71.676
R1239 B.n237 B.n67 71.676
R1240 B.n241 B.n68 71.676
R1241 B.n245 B.n69 71.676
R1242 B.n249 B.n70 71.676
R1243 B.n253 B.n71 71.676
R1244 B.n257 B.n72 71.676
R1245 B.n261 B.n73 71.676
R1246 B.n265 B.n74 71.676
R1247 B.n269 B.n75 71.676
R1248 B.n602 B.n76 71.676
R1249 B.n602 B.n601 71.676
R1250 B.n271 B.n75 71.676
R1251 B.n268 B.n74 71.676
R1252 B.n264 B.n73 71.676
R1253 B.n260 B.n72 71.676
R1254 B.n256 B.n71 71.676
R1255 B.n252 B.n70 71.676
R1256 B.n248 B.n69 71.676
R1257 B.n244 B.n68 71.676
R1258 B.n240 B.n67 71.676
R1259 B.n236 B.n66 71.676
R1260 B.n232 B.n65 71.676
R1261 B.n228 B.n64 71.676
R1262 B.n224 B.n63 71.676
R1263 B.n220 B.n62 71.676
R1264 B.n216 B.n61 71.676
R1265 B.n212 B.n60 71.676
R1266 B.n208 B.n59 71.676
R1267 B.n204 B.n58 71.676
R1268 B.n200 B.n57 71.676
R1269 B.n196 B.n56 71.676
R1270 B.n192 B.n55 71.676
R1271 B.n188 B.n54 71.676
R1272 B.n184 B.n53 71.676
R1273 B.n180 B.n52 71.676
R1274 B.n176 B.n51 71.676
R1275 B.n172 B.n50 71.676
R1276 B.n168 B.n49 71.676
R1277 B.n164 B.n48 71.676
R1278 B.n160 B.n47 71.676
R1279 B.n156 B.n46 71.676
R1280 B.n152 B.n45 71.676
R1281 B.n148 B.n44 71.676
R1282 B.n144 B.n43 71.676
R1283 B.n140 B.n42 71.676
R1284 B.n136 B.n41 71.676
R1285 B.n132 B.n40 71.676
R1286 B.n128 B.n39 71.676
R1287 B.n124 B.n38 71.676
R1288 B.n120 B.n37 71.676
R1289 B.n116 B.n36 71.676
R1290 B.n112 B.n35 71.676
R1291 B.n108 B.n34 71.676
R1292 B.n104 B.n33 71.676
R1293 B.n100 B.n32 71.676
R1294 B.n96 B.n31 71.676
R1295 B.n92 B.n30 71.676
R1296 B.n88 B.n29 71.676
R1297 B.n84 B.n28 71.676
R1298 B.n348 B.n294 71.676
R1299 B.n352 B.n351 71.676
R1300 B.n357 B.n356 71.676
R1301 B.n360 B.n359 71.676
R1302 B.n365 B.n364 71.676
R1303 B.n368 B.n367 71.676
R1304 B.n373 B.n372 71.676
R1305 B.n376 B.n375 71.676
R1306 B.n381 B.n380 71.676
R1307 B.n384 B.n383 71.676
R1308 B.n389 B.n388 71.676
R1309 B.n392 B.n391 71.676
R1310 B.n397 B.n396 71.676
R1311 B.n400 B.n399 71.676
R1312 B.n405 B.n404 71.676
R1313 B.n408 B.n407 71.676
R1314 B.n413 B.n412 71.676
R1315 B.n416 B.n415 71.676
R1316 B.n421 B.n420 71.676
R1317 B.n424 B.n423 71.676
R1318 B.n429 B.n428 71.676
R1319 B.n432 B.n431 71.676
R1320 B.n438 B.n437 71.676
R1321 B.n441 B.n440 71.676
R1322 B.n446 B.n445 71.676
R1323 B.n449 B.n448 71.676
R1324 B.n457 B.n456 71.676
R1325 B.n460 B.n459 71.676
R1326 B.n465 B.n464 71.676
R1327 B.n468 B.n467 71.676
R1328 B.n473 B.n472 71.676
R1329 B.n476 B.n475 71.676
R1330 B.n481 B.n480 71.676
R1331 B.n484 B.n483 71.676
R1332 B.n489 B.n488 71.676
R1333 B.n492 B.n491 71.676
R1334 B.n497 B.n496 71.676
R1335 B.n500 B.n499 71.676
R1336 B.n505 B.n504 71.676
R1337 B.n508 B.n507 71.676
R1338 B.n513 B.n512 71.676
R1339 B.n516 B.n515 71.676
R1340 B.n521 B.n520 71.676
R1341 B.n524 B.n523 71.676
R1342 B.n529 B.n528 71.676
R1343 B.n532 B.n531 71.676
R1344 B.n537 B.n536 71.676
R1345 B.n540 B.n539 71.676
R1346 B.n349 B.n348 71.676
R1347 B.n351 B.n345 71.676
R1348 B.n358 B.n357 71.676
R1349 B.n359 B.n343 71.676
R1350 B.n366 B.n365 71.676
R1351 B.n367 B.n341 71.676
R1352 B.n374 B.n373 71.676
R1353 B.n375 B.n339 71.676
R1354 B.n382 B.n381 71.676
R1355 B.n383 B.n337 71.676
R1356 B.n390 B.n389 71.676
R1357 B.n391 B.n335 71.676
R1358 B.n398 B.n397 71.676
R1359 B.n399 B.n333 71.676
R1360 B.n406 B.n405 71.676
R1361 B.n407 B.n331 71.676
R1362 B.n414 B.n413 71.676
R1363 B.n415 B.n329 71.676
R1364 B.n422 B.n421 71.676
R1365 B.n423 B.n327 71.676
R1366 B.n430 B.n429 71.676
R1367 B.n431 B.n323 71.676
R1368 B.n439 B.n438 71.676
R1369 B.n440 B.n321 71.676
R1370 B.n447 B.n446 71.676
R1371 B.n448 B.n319 71.676
R1372 B.n458 B.n457 71.676
R1373 B.n459 B.n317 71.676
R1374 B.n466 B.n465 71.676
R1375 B.n467 B.n315 71.676
R1376 B.n474 B.n473 71.676
R1377 B.n475 B.n313 71.676
R1378 B.n482 B.n481 71.676
R1379 B.n483 B.n311 71.676
R1380 B.n490 B.n489 71.676
R1381 B.n491 B.n309 71.676
R1382 B.n498 B.n497 71.676
R1383 B.n499 B.n307 71.676
R1384 B.n506 B.n505 71.676
R1385 B.n507 B.n305 71.676
R1386 B.n514 B.n513 71.676
R1387 B.n515 B.n303 71.676
R1388 B.n522 B.n521 71.676
R1389 B.n523 B.n301 71.676
R1390 B.n530 B.n529 71.676
R1391 B.n531 B.n299 71.676
R1392 B.n538 B.n537 71.676
R1393 B.n541 B.n540 71.676
R1394 B.n631 B.n630 71.676
R1395 B.n631 B.n2 71.676
R1396 B.n82 B.n81 59.5399
R1397 B.n79 B.n78 59.5399
R1398 B.n454 B.n453 59.5399
R1399 B.n434 B.n325 59.5399
R1400 B.n546 B.n291 41.2922
R1401 B.n552 B.n291 41.2922
R1402 B.n552 B.n287 41.2922
R1403 B.n558 B.n287 41.2922
R1404 B.n564 B.n283 41.2922
R1405 B.n564 B.n279 41.2922
R1406 B.n572 B.n279 41.2922
R1407 B.n572 B.n571 41.2922
R1408 B.n578 B.n4 41.2922
R1409 B.n629 B.n4 41.2922
R1410 B.n629 B.n628 41.2922
R1411 B.n628 B.n627 41.2922
R1412 B.n627 B.n8 41.2922
R1413 B.n620 B.n12 41.2922
R1414 B.n620 B.n619 41.2922
R1415 B.n619 B.n618 41.2922
R1416 B.n618 B.n16 41.2922
R1417 B.n612 B.n611 41.2922
R1418 B.n611 B.n610 41.2922
R1419 B.n610 B.n23 41.2922
R1420 B.n604 B.n23 41.2922
R1421 B.n571 B.t1 33.3982
R1422 B.n12 B.t0 33.3982
R1423 B.n548 B.n293 30.7517
R1424 B.n544 B.n543 30.7517
R1425 B.n600 B.n599 30.7517
R1426 B.n606 B.n25 30.7517
R1427 B.t3 B.n283 23.6825
R1428 B.t10 B.n16 23.6825
R1429 B B.n632 18.0485
R1430 B.n558 B.t3 17.6102
R1431 B.n612 B.t10 17.6102
R1432 B.n81 B.n80 14.352
R1433 B.n78 B.n77 14.352
R1434 B.n453 B.n452 14.352
R1435 B.n325 B.n324 14.352
R1436 B.n549 B.n548 10.6151
R1437 B.n550 B.n549 10.6151
R1438 B.n550 B.n285 10.6151
R1439 B.n560 B.n285 10.6151
R1440 B.n561 B.n560 10.6151
R1441 B.n562 B.n561 10.6151
R1442 B.n562 B.n277 10.6151
R1443 B.n574 B.n277 10.6151
R1444 B.n575 B.n574 10.6151
R1445 B.n576 B.n575 10.6151
R1446 B.n576 B.n0 10.6151
R1447 B.n347 B.n293 10.6151
R1448 B.n347 B.n346 10.6151
R1449 B.n353 B.n346 10.6151
R1450 B.n354 B.n353 10.6151
R1451 B.n355 B.n354 10.6151
R1452 B.n355 B.n344 10.6151
R1453 B.n361 B.n344 10.6151
R1454 B.n362 B.n361 10.6151
R1455 B.n363 B.n362 10.6151
R1456 B.n363 B.n342 10.6151
R1457 B.n369 B.n342 10.6151
R1458 B.n370 B.n369 10.6151
R1459 B.n371 B.n370 10.6151
R1460 B.n371 B.n340 10.6151
R1461 B.n377 B.n340 10.6151
R1462 B.n378 B.n377 10.6151
R1463 B.n379 B.n378 10.6151
R1464 B.n379 B.n338 10.6151
R1465 B.n385 B.n338 10.6151
R1466 B.n386 B.n385 10.6151
R1467 B.n387 B.n386 10.6151
R1468 B.n387 B.n336 10.6151
R1469 B.n393 B.n336 10.6151
R1470 B.n394 B.n393 10.6151
R1471 B.n395 B.n394 10.6151
R1472 B.n395 B.n334 10.6151
R1473 B.n401 B.n334 10.6151
R1474 B.n402 B.n401 10.6151
R1475 B.n403 B.n402 10.6151
R1476 B.n403 B.n332 10.6151
R1477 B.n409 B.n332 10.6151
R1478 B.n410 B.n409 10.6151
R1479 B.n411 B.n410 10.6151
R1480 B.n411 B.n330 10.6151
R1481 B.n417 B.n330 10.6151
R1482 B.n418 B.n417 10.6151
R1483 B.n419 B.n418 10.6151
R1484 B.n419 B.n328 10.6151
R1485 B.n425 B.n328 10.6151
R1486 B.n426 B.n425 10.6151
R1487 B.n427 B.n426 10.6151
R1488 B.n427 B.n326 10.6151
R1489 B.n433 B.n326 10.6151
R1490 B.n436 B.n435 10.6151
R1491 B.n436 B.n322 10.6151
R1492 B.n442 B.n322 10.6151
R1493 B.n443 B.n442 10.6151
R1494 B.n444 B.n443 10.6151
R1495 B.n444 B.n320 10.6151
R1496 B.n450 B.n320 10.6151
R1497 B.n451 B.n450 10.6151
R1498 B.n455 B.n451 10.6151
R1499 B.n461 B.n318 10.6151
R1500 B.n462 B.n461 10.6151
R1501 B.n463 B.n462 10.6151
R1502 B.n463 B.n316 10.6151
R1503 B.n469 B.n316 10.6151
R1504 B.n470 B.n469 10.6151
R1505 B.n471 B.n470 10.6151
R1506 B.n471 B.n314 10.6151
R1507 B.n477 B.n314 10.6151
R1508 B.n478 B.n477 10.6151
R1509 B.n479 B.n478 10.6151
R1510 B.n479 B.n312 10.6151
R1511 B.n485 B.n312 10.6151
R1512 B.n486 B.n485 10.6151
R1513 B.n487 B.n486 10.6151
R1514 B.n487 B.n310 10.6151
R1515 B.n493 B.n310 10.6151
R1516 B.n494 B.n493 10.6151
R1517 B.n495 B.n494 10.6151
R1518 B.n495 B.n308 10.6151
R1519 B.n501 B.n308 10.6151
R1520 B.n502 B.n501 10.6151
R1521 B.n503 B.n502 10.6151
R1522 B.n503 B.n306 10.6151
R1523 B.n509 B.n306 10.6151
R1524 B.n510 B.n509 10.6151
R1525 B.n511 B.n510 10.6151
R1526 B.n511 B.n304 10.6151
R1527 B.n517 B.n304 10.6151
R1528 B.n518 B.n517 10.6151
R1529 B.n519 B.n518 10.6151
R1530 B.n519 B.n302 10.6151
R1531 B.n525 B.n302 10.6151
R1532 B.n526 B.n525 10.6151
R1533 B.n527 B.n526 10.6151
R1534 B.n527 B.n300 10.6151
R1535 B.n533 B.n300 10.6151
R1536 B.n534 B.n533 10.6151
R1537 B.n535 B.n534 10.6151
R1538 B.n535 B.n298 10.6151
R1539 B.n298 B.n297 10.6151
R1540 B.n542 B.n297 10.6151
R1541 B.n543 B.n542 10.6151
R1542 B.n544 B.n289 10.6151
R1543 B.n554 B.n289 10.6151
R1544 B.n555 B.n554 10.6151
R1545 B.n556 B.n555 10.6151
R1546 B.n556 B.n281 10.6151
R1547 B.n566 B.n281 10.6151
R1548 B.n567 B.n566 10.6151
R1549 B.n569 B.n567 10.6151
R1550 B.n569 B.n568 10.6151
R1551 B.n568 B.n274 10.6151
R1552 B.n581 B.n274 10.6151
R1553 B.n582 B.n581 10.6151
R1554 B.n583 B.n582 10.6151
R1555 B.n584 B.n583 10.6151
R1556 B.n585 B.n584 10.6151
R1557 B.n588 B.n585 10.6151
R1558 B.n589 B.n588 10.6151
R1559 B.n590 B.n589 10.6151
R1560 B.n591 B.n590 10.6151
R1561 B.n593 B.n591 10.6151
R1562 B.n594 B.n593 10.6151
R1563 B.n595 B.n594 10.6151
R1564 B.n596 B.n595 10.6151
R1565 B.n598 B.n596 10.6151
R1566 B.n599 B.n598 10.6151
R1567 B.n624 B.n1 10.6151
R1568 B.n624 B.n623 10.6151
R1569 B.n623 B.n622 10.6151
R1570 B.n622 B.n10 10.6151
R1571 B.n616 B.n10 10.6151
R1572 B.n616 B.n615 10.6151
R1573 B.n615 B.n614 10.6151
R1574 B.n614 B.n18 10.6151
R1575 B.n608 B.n18 10.6151
R1576 B.n608 B.n607 10.6151
R1577 B.n607 B.n606 10.6151
R1578 B.n83 B.n25 10.6151
R1579 B.n86 B.n83 10.6151
R1580 B.n87 B.n86 10.6151
R1581 B.n90 B.n87 10.6151
R1582 B.n91 B.n90 10.6151
R1583 B.n94 B.n91 10.6151
R1584 B.n95 B.n94 10.6151
R1585 B.n98 B.n95 10.6151
R1586 B.n99 B.n98 10.6151
R1587 B.n102 B.n99 10.6151
R1588 B.n103 B.n102 10.6151
R1589 B.n106 B.n103 10.6151
R1590 B.n107 B.n106 10.6151
R1591 B.n110 B.n107 10.6151
R1592 B.n111 B.n110 10.6151
R1593 B.n114 B.n111 10.6151
R1594 B.n115 B.n114 10.6151
R1595 B.n118 B.n115 10.6151
R1596 B.n119 B.n118 10.6151
R1597 B.n122 B.n119 10.6151
R1598 B.n123 B.n122 10.6151
R1599 B.n126 B.n123 10.6151
R1600 B.n127 B.n126 10.6151
R1601 B.n130 B.n127 10.6151
R1602 B.n131 B.n130 10.6151
R1603 B.n134 B.n131 10.6151
R1604 B.n135 B.n134 10.6151
R1605 B.n138 B.n135 10.6151
R1606 B.n139 B.n138 10.6151
R1607 B.n142 B.n139 10.6151
R1608 B.n143 B.n142 10.6151
R1609 B.n146 B.n143 10.6151
R1610 B.n147 B.n146 10.6151
R1611 B.n150 B.n147 10.6151
R1612 B.n151 B.n150 10.6151
R1613 B.n154 B.n151 10.6151
R1614 B.n155 B.n154 10.6151
R1615 B.n158 B.n155 10.6151
R1616 B.n159 B.n158 10.6151
R1617 B.n162 B.n159 10.6151
R1618 B.n163 B.n162 10.6151
R1619 B.n166 B.n163 10.6151
R1620 B.n167 B.n166 10.6151
R1621 B.n171 B.n170 10.6151
R1622 B.n174 B.n171 10.6151
R1623 B.n175 B.n174 10.6151
R1624 B.n178 B.n175 10.6151
R1625 B.n179 B.n178 10.6151
R1626 B.n182 B.n179 10.6151
R1627 B.n183 B.n182 10.6151
R1628 B.n186 B.n183 10.6151
R1629 B.n187 B.n186 10.6151
R1630 B.n191 B.n190 10.6151
R1631 B.n194 B.n191 10.6151
R1632 B.n195 B.n194 10.6151
R1633 B.n198 B.n195 10.6151
R1634 B.n199 B.n198 10.6151
R1635 B.n202 B.n199 10.6151
R1636 B.n203 B.n202 10.6151
R1637 B.n206 B.n203 10.6151
R1638 B.n207 B.n206 10.6151
R1639 B.n210 B.n207 10.6151
R1640 B.n211 B.n210 10.6151
R1641 B.n214 B.n211 10.6151
R1642 B.n215 B.n214 10.6151
R1643 B.n218 B.n215 10.6151
R1644 B.n219 B.n218 10.6151
R1645 B.n222 B.n219 10.6151
R1646 B.n223 B.n222 10.6151
R1647 B.n226 B.n223 10.6151
R1648 B.n227 B.n226 10.6151
R1649 B.n230 B.n227 10.6151
R1650 B.n231 B.n230 10.6151
R1651 B.n234 B.n231 10.6151
R1652 B.n235 B.n234 10.6151
R1653 B.n238 B.n235 10.6151
R1654 B.n239 B.n238 10.6151
R1655 B.n242 B.n239 10.6151
R1656 B.n243 B.n242 10.6151
R1657 B.n246 B.n243 10.6151
R1658 B.n247 B.n246 10.6151
R1659 B.n250 B.n247 10.6151
R1660 B.n251 B.n250 10.6151
R1661 B.n254 B.n251 10.6151
R1662 B.n255 B.n254 10.6151
R1663 B.n258 B.n255 10.6151
R1664 B.n259 B.n258 10.6151
R1665 B.n262 B.n259 10.6151
R1666 B.n263 B.n262 10.6151
R1667 B.n266 B.n263 10.6151
R1668 B.n267 B.n266 10.6151
R1669 B.n270 B.n267 10.6151
R1670 B.n272 B.n270 10.6151
R1671 B.n273 B.n272 10.6151
R1672 B.n600 B.n273 10.6151
R1673 B.n434 B.n433 8.74196
R1674 B.n454 B.n318 8.74196
R1675 B.n167 B.n82 8.74196
R1676 B.n190 B.n79 8.74196
R1677 B.n632 B.n0 8.11757
R1678 B.n632 B.n1 8.11757
R1679 B.n578 B.t1 7.89451
R1680 B.t0 B.n8 7.89451
R1681 B.n435 B.n434 1.87367
R1682 B.n455 B.n454 1.87367
R1683 B.n170 B.n82 1.87367
R1684 B.n187 B.n79 1.87367
R1685 VP.n0 VP.t1 1051.34
R1686 VP.n0 VP.t0 1011.85
R1687 VP VP.n0 0.0516364
R1688 VDD1.n64 VDD1.n0 289.615
R1689 VDD1.n133 VDD1.n69 289.615
R1690 VDD1.n65 VDD1.n64 185
R1691 VDD1.n63 VDD1.n62 185
R1692 VDD1.n4 VDD1.n3 185
R1693 VDD1.n57 VDD1.n56 185
R1694 VDD1.n55 VDD1.n54 185
R1695 VDD1.n8 VDD1.n7 185
R1696 VDD1.n49 VDD1.n48 185
R1697 VDD1.n47 VDD1.n46 185
R1698 VDD1.n45 VDD1.n11 185
R1699 VDD1.n15 VDD1.n12 185
R1700 VDD1.n40 VDD1.n39 185
R1701 VDD1.n38 VDD1.n37 185
R1702 VDD1.n17 VDD1.n16 185
R1703 VDD1.n32 VDD1.n31 185
R1704 VDD1.n30 VDD1.n29 185
R1705 VDD1.n21 VDD1.n20 185
R1706 VDD1.n24 VDD1.n23 185
R1707 VDD1.n92 VDD1.n91 185
R1708 VDD1.n89 VDD1.n88 185
R1709 VDD1.n98 VDD1.n97 185
R1710 VDD1.n100 VDD1.n99 185
R1711 VDD1.n85 VDD1.n84 185
R1712 VDD1.n106 VDD1.n105 185
R1713 VDD1.n109 VDD1.n108 185
R1714 VDD1.n107 VDD1.n81 185
R1715 VDD1.n114 VDD1.n80 185
R1716 VDD1.n116 VDD1.n115 185
R1717 VDD1.n118 VDD1.n117 185
R1718 VDD1.n77 VDD1.n76 185
R1719 VDD1.n124 VDD1.n123 185
R1720 VDD1.n126 VDD1.n125 185
R1721 VDD1.n73 VDD1.n72 185
R1722 VDD1.n132 VDD1.n131 185
R1723 VDD1.n134 VDD1.n133 185
R1724 VDD1.t0 VDD1.n22 149.524
R1725 VDD1.t1 VDD1.n90 149.524
R1726 VDD1.n64 VDD1.n63 104.615
R1727 VDD1.n63 VDD1.n3 104.615
R1728 VDD1.n56 VDD1.n3 104.615
R1729 VDD1.n56 VDD1.n55 104.615
R1730 VDD1.n55 VDD1.n7 104.615
R1731 VDD1.n48 VDD1.n7 104.615
R1732 VDD1.n48 VDD1.n47 104.615
R1733 VDD1.n47 VDD1.n11 104.615
R1734 VDD1.n15 VDD1.n11 104.615
R1735 VDD1.n39 VDD1.n15 104.615
R1736 VDD1.n39 VDD1.n38 104.615
R1737 VDD1.n38 VDD1.n16 104.615
R1738 VDD1.n31 VDD1.n16 104.615
R1739 VDD1.n31 VDD1.n30 104.615
R1740 VDD1.n30 VDD1.n20 104.615
R1741 VDD1.n23 VDD1.n20 104.615
R1742 VDD1.n91 VDD1.n88 104.615
R1743 VDD1.n98 VDD1.n88 104.615
R1744 VDD1.n99 VDD1.n98 104.615
R1745 VDD1.n99 VDD1.n84 104.615
R1746 VDD1.n106 VDD1.n84 104.615
R1747 VDD1.n108 VDD1.n106 104.615
R1748 VDD1.n108 VDD1.n107 104.615
R1749 VDD1.n107 VDD1.n80 104.615
R1750 VDD1.n116 VDD1.n80 104.615
R1751 VDD1.n117 VDD1.n116 104.615
R1752 VDD1.n117 VDD1.n76 104.615
R1753 VDD1.n124 VDD1.n76 104.615
R1754 VDD1.n125 VDD1.n124 104.615
R1755 VDD1.n125 VDD1.n72 104.615
R1756 VDD1.n132 VDD1.n72 104.615
R1757 VDD1.n133 VDD1.n132 104.615
R1758 VDD1 VDD1.n137 85.1648
R1759 VDD1.n23 VDD1.t0 52.3082
R1760 VDD1.n91 VDD1.t1 52.3082
R1761 VDD1 VDD1.n68 48.6939
R1762 VDD1.n46 VDD1.n45 13.1884
R1763 VDD1.n115 VDD1.n114 13.1884
R1764 VDD1.n49 VDD1.n10 12.8005
R1765 VDD1.n44 VDD1.n12 12.8005
R1766 VDD1.n113 VDD1.n81 12.8005
R1767 VDD1.n118 VDD1.n79 12.8005
R1768 VDD1.n50 VDD1.n8 12.0247
R1769 VDD1.n41 VDD1.n40 12.0247
R1770 VDD1.n110 VDD1.n109 12.0247
R1771 VDD1.n119 VDD1.n77 12.0247
R1772 VDD1.n54 VDD1.n53 11.249
R1773 VDD1.n37 VDD1.n14 11.249
R1774 VDD1.n105 VDD1.n83 11.249
R1775 VDD1.n123 VDD1.n122 11.249
R1776 VDD1.n57 VDD1.n6 10.4732
R1777 VDD1.n36 VDD1.n17 10.4732
R1778 VDD1.n104 VDD1.n85 10.4732
R1779 VDD1.n126 VDD1.n75 10.4732
R1780 VDD1.n24 VDD1.n22 10.2747
R1781 VDD1.n92 VDD1.n90 10.2747
R1782 VDD1.n58 VDD1.n4 9.69747
R1783 VDD1.n33 VDD1.n32 9.69747
R1784 VDD1.n101 VDD1.n100 9.69747
R1785 VDD1.n127 VDD1.n73 9.69747
R1786 VDD1.n68 VDD1.n67 9.45567
R1787 VDD1.n137 VDD1.n136 9.45567
R1788 VDD1.n26 VDD1.n25 9.3005
R1789 VDD1.n28 VDD1.n27 9.3005
R1790 VDD1.n19 VDD1.n18 9.3005
R1791 VDD1.n34 VDD1.n33 9.3005
R1792 VDD1.n36 VDD1.n35 9.3005
R1793 VDD1.n14 VDD1.n13 9.3005
R1794 VDD1.n42 VDD1.n41 9.3005
R1795 VDD1.n44 VDD1.n43 9.3005
R1796 VDD1.n67 VDD1.n66 9.3005
R1797 VDD1.n2 VDD1.n1 9.3005
R1798 VDD1.n61 VDD1.n60 9.3005
R1799 VDD1.n59 VDD1.n58 9.3005
R1800 VDD1.n6 VDD1.n5 9.3005
R1801 VDD1.n53 VDD1.n52 9.3005
R1802 VDD1.n51 VDD1.n50 9.3005
R1803 VDD1.n10 VDD1.n9 9.3005
R1804 VDD1.n71 VDD1.n70 9.3005
R1805 VDD1.n130 VDD1.n129 9.3005
R1806 VDD1.n128 VDD1.n127 9.3005
R1807 VDD1.n75 VDD1.n74 9.3005
R1808 VDD1.n122 VDD1.n121 9.3005
R1809 VDD1.n120 VDD1.n119 9.3005
R1810 VDD1.n79 VDD1.n78 9.3005
R1811 VDD1.n94 VDD1.n93 9.3005
R1812 VDD1.n96 VDD1.n95 9.3005
R1813 VDD1.n87 VDD1.n86 9.3005
R1814 VDD1.n102 VDD1.n101 9.3005
R1815 VDD1.n104 VDD1.n103 9.3005
R1816 VDD1.n83 VDD1.n82 9.3005
R1817 VDD1.n111 VDD1.n110 9.3005
R1818 VDD1.n113 VDD1.n112 9.3005
R1819 VDD1.n136 VDD1.n135 9.3005
R1820 VDD1.n62 VDD1.n61 8.92171
R1821 VDD1.n29 VDD1.n19 8.92171
R1822 VDD1.n97 VDD1.n87 8.92171
R1823 VDD1.n131 VDD1.n130 8.92171
R1824 VDD1.n65 VDD1.n2 8.14595
R1825 VDD1.n28 VDD1.n21 8.14595
R1826 VDD1.n96 VDD1.n89 8.14595
R1827 VDD1.n134 VDD1.n71 8.14595
R1828 VDD1.n66 VDD1.n0 7.3702
R1829 VDD1.n25 VDD1.n24 7.3702
R1830 VDD1.n93 VDD1.n92 7.3702
R1831 VDD1.n135 VDD1.n69 7.3702
R1832 VDD1.n68 VDD1.n0 6.59444
R1833 VDD1.n137 VDD1.n69 6.59444
R1834 VDD1.n66 VDD1.n65 5.81868
R1835 VDD1.n25 VDD1.n21 5.81868
R1836 VDD1.n93 VDD1.n89 5.81868
R1837 VDD1.n135 VDD1.n134 5.81868
R1838 VDD1.n62 VDD1.n2 5.04292
R1839 VDD1.n29 VDD1.n28 5.04292
R1840 VDD1.n97 VDD1.n96 5.04292
R1841 VDD1.n131 VDD1.n71 5.04292
R1842 VDD1.n61 VDD1.n4 4.26717
R1843 VDD1.n32 VDD1.n19 4.26717
R1844 VDD1.n100 VDD1.n87 4.26717
R1845 VDD1.n130 VDD1.n73 4.26717
R1846 VDD1.n58 VDD1.n57 3.49141
R1847 VDD1.n33 VDD1.n17 3.49141
R1848 VDD1.n101 VDD1.n85 3.49141
R1849 VDD1.n127 VDD1.n126 3.49141
R1850 VDD1.n26 VDD1.n22 2.84303
R1851 VDD1.n94 VDD1.n90 2.84303
R1852 VDD1.n54 VDD1.n6 2.71565
R1853 VDD1.n37 VDD1.n36 2.71565
R1854 VDD1.n105 VDD1.n104 2.71565
R1855 VDD1.n123 VDD1.n75 2.71565
R1856 VDD1.n53 VDD1.n8 1.93989
R1857 VDD1.n40 VDD1.n14 1.93989
R1858 VDD1.n109 VDD1.n83 1.93989
R1859 VDD1.n122 VDD1.n77 1.93989
R1860 VDD1.n50 VDD1.n49 1.16414
R1861 VDD1.n41 VDD1.n12 1.16414
R1862 VDD1.n110 VDD1.n81 1.16414
R1863 VDD1.n119 VDD1.n118 1.16414
R1864 VDD1.n46 VDD1.n10 0.388379
R1865 VDD1.n45 VDD1.n44 0.388379
R1866 VDD1.n114 VDD1.n113 0.388379
R1867 VDD1.n115 VDD1.n79 0.388379
R1868 VDD1.n67 VDD1.n1 0.155672
R1869 VDD1.n60 VDD1.n1 0.155672
R1870 VDD1.n60 VDD1.n59 0.155672
R1871 VDD1.n59 VDD1.n5 0.155672
R1872 VDD1.n52 VDD1.n5 0.155672
R1873 VDD1.n52 VDD1.n51 0.155672
R1874 VDD1.n51 VDD1.n9 0.155672
R1875 VDD1.n43 VDD1.n9 0.155672
R1876 VDD1.n43 VDD1.n42 0.155672
R1877 VDD1.n42 VDD1.n13 0.155672
R1878 VDD1.n35 VDD1.n13 0.155672
R1879 VDD1.n35 VDD1.n34 0.155672
R1880 VDD1.n34 VDD1.n18 0.155672
R1881 VDD1.n27 VDD1.n18 0.155672
R1882 VDD1.n27 VDD1.n26 0.155672
R1883 VDD1.n95 VDD1.n94 0.155672
R1884 VDD1.n95 VDD1.n86 0.155672
R1885 VDD1.n102 VDD1.n86 0.155672
R1886 VDD1.n103 VDD1.n102 0.155672
R1887 VDD1.n103 VDD1.n82 0.155672
R1888 VDD1.n111 VDD1.n82 0.155672
R1889 VDD1.n112 VDD1.n111 0.155672
R1890 VDD1.n112 VDD1.n78 0.155672
R1891 VDD1.n120 VDD1.n78 0.155672
R1892 VDD1.n121 VDD1.n120 0.155672
R1893 VDD1.n121 VDD1.n74 0.155672
R1894 VDD1.n128 VDD1.n74 0.155672
R1895 VDD1.n129 VDD1.n128 0.155672
R1896 VDD1.n129 VDD1.n70 0.155672
R1897 VDD1.n136 VDD1.n70 0.155672
C0 VN VTAIL 1.12025f
C1 VDD1 VN 0.148123f
C2 VP VDD2 0.242786f
C3 VP VTAIL 1.135f
C4 VP VDD1 1.80879f
C5 VP VN 4.58435f
C6 VDD2 VTAIL 6.80741f
C7 VDD1 VDD2 0.436168f
C8 VDD1 VTAIL 6.77734f
C9 VDD2 VN 1.71931f
C10 VDD2 B 3.788744f
C11 VDD1 B 5.85711f
C12 VTAIL B 6.032257f
C13 VN B 7.11748f
C14 VP B 3.732842f
C15 VDD1.n0 B 0.024955f
C16 VDD1.n1 B 0.017585f
C17 VDD1.n2 B 0.00945f
C18 VDD1.n3 B 0.022336f
C19 VDD1.n4 B 0.010006f
C20 VDD1.n5 B 0.017585f
C21 VDD1.n6 B 0.00945f
C22 VDD1.n7 B 0.022336f
C23 VDD1.n8 B 0.010006f
C24 VDD1.n9 B 0.017585f
C25 VDD1.n10 B 0.00945f
C26 VDD1.n11 B 0.022336f
C27 VDD1.n12 B 0.010006f
C28 VDD1.n13 B 0.017585f
C29 VDD1.n14 B 0.00945f
C30 VDD1.n15 B 0.022336f
C31 VDD1.n16 B 0.022336f
C32 VDD1.n17 B 0.010006f
C33 VDD1.n18 B 0.017585f
C34 VDD1.n19 B 0.00945f
C35 VDD1.n20 B 0.022336f
C36 VDD1.n21 B 0.010006f
C37 VDD1.n22 B 0.132325f
C38 VDD1.t0 B 0.037801f
C39 VDD1.n23 B 0.016752f
C40 VDD1.n24 B 0.015789f
C41 VDD1.n25 B 0.00945f
C42 VDD1.n26 B 0.951292f
C43 VDD1.n27 B 0.017585f
C44 VDD1.n28 B 0.00945f
C45 VDD1.n29 B 0.010006f
C46 VDD1.n30 B 0.022336f
C47 VDD1.n31 B 0.022336f
C48 VDD1.n32 B 0.010006f
C49 VDD1.n33 B 0.00945f
C50 VDD1.n34 B 0.017585f
C51 VDD1.n35 B 0.017585f
C52 VDD1.n36 B 0.00945f
C53 VDD1.n37 B 0.010006f
C54 VDD1.n38 B 0.022336f
C55 VDD1.n39 B 0.022336f
C56 VDD1.n40 B 0.010006f
C57 VDD1.n41 B 0.00945f
C58 VDD1.n42 B 0.017585f
C59 VDD1.n43 B 0.017585f
C60 VDD1.n44 B 0.00945f
C61 VDD1.n45 B 0.009728f
C62 VDD1.n46 B 0.009728f
C63 VDD1.n47 B 0.022336f
C64 VDD1.n48 B 0.022336f
C65 VDD1.n49 B 0.010006f
C66 VDD1.n50 B 0.00945f
C67 VDD1.n51 B 0.017585f
C68 VDD1.n52 B 0.017585f
C69 VDD1.n53 B 0.00945f
C70 VDD1.n54 B 0.010006f
C71 VDD1.n55 B 0.022336f
C72 VDD1.n56 B 0.022336f
C73 VDD1.n57 B 0.010006f
C74 VDD1.n58 B 0.00945f
C75 VDD1.n59 B 0.017585f
C76 VDD1.n60 B 0.017585f
C77 VDD1.n61 B 0.00945f
C78 VDD1.n62 B 0.010006f
C79 VDD1.n63 B 0.022336f
C80 VDD1.n64 B 0.048772f
C81 VDD1.n65 B 0.010006f
C82 VDD1.n66 B 0.00945f
C83 VDD1.n67 B 0.040167f
C84 VDD1.n68 B 0.03967f
C85 VDD1.n69 B 0.024955f
C86 VDD1.n70 B 0.017585f
C87 VDD1.n71 B 0.00945f
C88 VDD1.n72 B 0.022336f
C89 VDD1.n73 B 0.010006f
C90 VDD1.n74 B 0.017585f
C91 VDD1.n75 B 0.00945f
C92 VDD1.n76 B 0.022336f
C93 VDD1.n77 B 0.010006f
C94 VDD1.n78 B 0.017585f
C95 VDD1.n79 B 0.00945f
C96 VDD1.n80 B 0.022336f
C97 VDD1.n81 B 0.010006f
C98 VDD1.n82 B 0.017585f
C99 VDD1.n83 B 0.00945f
C100 VDD1.n84 B 0.022336f
C101 VDD1.n85 B 0.010006f
C102 VDD1.n86 B 0.017585f
C103 VDD1.n87 B 0.00945f
C104 VDD1.n88 B 0.022336f
C105 VDD1.n89 B 0.010006f
C106 VDD1.n90 B 0.132325f
C107 VDD1.t1 B 0.037801f
C108 VDD1.n91 B 0.016752f
C109 VDD1.n92 B 0.015789f
C110 VDD1.n93 B 0.00945f
C111 VDD1.n94 B 0.951292f
C112 VDD1.n95 B 0.017585f
C113 VDD1.n96 B 0.00945f
C114 VDD1.n97 B 0.010006f
C115 VDD1.n98 B 0.022336f
C116 VDD1.n99 B 0.022336f
C117 VDD1.n100 B 0.010006f
C118 VDD1.n101 B 0.00945f
C119 VDD1.n102 B 0.017585f
C120 VDD1.n103 B 0.017585f
C121 VDD1.n104 B 0.00945f
C122 VDD1.n105 B 0.010006f
C123 VDD1.n106 B 0.022336f
C124 VDD1.n107 B 0.022336f
C125 VDD1.n108 B 0.022336f
C126 VDD1.n109 B 0.010006f
C127 VDD1.n110 B 0.00945f
C128 VDD1.n111 B 0.017585f
C129 VDD1.n112 B 0.017585f
C130 VDD1.n113 B 0.00945f
C131 VDD1.n114 B 0.009728f
C132 VDD1.n115 B 0.009728f
C133 VDD1.n116 B 0.022336f
C134 VDD1.n117 B 0.022336f
C135 VDD1.n118 B 0.010006f
C136 VDD1.n119 B 0.00945f
C137 VDD1.n120 B 0.017585f
C138 VDD1.n121 B 0.017585f
C139 VDD1.n122 B 0.00945f
C140 VDD1.n123 B 0.010006f
C141 VDD1.n124 B 0.022336f
C142 VDD1.n125 B 0.022336f
C143 VDD1.n126 B 0.010006f
C144 VDD1.n127 B 0.00945f
C145 VDD1.n128 B 0.017585f
C146 VDD1.n129 B 0.017585f
C147 VDD1.n130 B 0.00945f
C148 VDD1.n131 B 0.010006f
C149 VDD1.n132 B 0.022336f
C150 VDD1.n133 B 0.048772f
C151 VDD1.n134 B 0.010006f
C152 VDD1.n135 B 0.00945f
C153 VDD1.n136 B 0.040167f
C154 VDD1.n137 B 0.462993f
C155 VP.t1 B 0.689115f
C156 VP.t0 B 0.62696f
C157 VP.n0 B 3.27724f
C158 VDD2.n0 B 0.025196f
C159 VDD2.n1 B 0.017755f
C160 VDD2.n2 B 0.009541f
C161 VDD2.n3 B 0.022551f
C162 VDD2.n4 B 0.010102f
C163 VDD2.n5 B 0.017755f
C164 VDD2.n6 B 0.009541f
C165 VDD2.n7 B 0.022551f
C166 VDD2.n8 B 0.010102f
C167 VDD2.n9 B 0.017755f
C168 VDD2.n10 B 0.009541f
C169 VDD2.n11 B 0.022551f
C170 VDD2.n12 B 0.010102f
C171 VDD2.n13 B 0.017755f
C172 VDD2.n14 B 0.009541f
C173 VDD2.n15 B 0.022551f
C174 VDD2.n16 B 0.010102f
C175 VDD2.n17 B 0.017755f
C176 VDD2.n18 B 0.009541f
C177 VDD2.n19 B 0.022551f
C178 VDD2.n20 B 0.010102f
C179 VDD2.n21 B 0.133601f
C180 VDD2.t0 B 0.038165f
C181 VDD2.n22 B 0.016913f
C182 VDD2.n23 B 0.015942f
C183 VDD2.n24 B 0.009541f
C184 VDD2.n25 B 0.960466f
C185 VDD2.n26 B 0.017755f
C186 VDD2.n27 B 0.009541f
C187 VDD2.n28 B 0.010102f
C188 VDD2.n29 B 0.022551f
C189 VDD2.n30 B 0.022551f
C190 VDD2.n31 B 0.010102f
C191 VDD2.n32 B 0.009541f
C192 VDD2.n33 B 0.017755f
C193 VDD2.n34 B 0.017755f
C194 VDD2.n35 B 0.009541f
C195 VDD2.n36 B 0.010102f
C196 VDD2.n37 B 0.022551f
C197 VDD2.n38 B 0.022551f
C198 VDD2.n39 B 0.022551f
C199 VDD2.n40 B 0.010102f
C200 VDD2.n41 B 0.009541f
C201 VDD2.n42 B 0.017755f
C202 VDD2.n43 B 0.017755f
C203 VDD2.n44 B 0.009541f
C204 VDD2.n45 B 0.009821f
C205 VDD2.n46 B 0.009821f
C206 VDD2.n47 B 0.022551f
C207 VDD2.n48 B 0.022551f
C208 VDD2.n49 B 0.010102f
C209 VDD2.n50 B 0.009541f
C210 VDD2.n51 B 0.017755f
C211 VDD2.n52 B 0.017755f
C212 VDD2.n53 B 0.009541f
C213 VDD2.n54 B 0.010102f
C214 VDD2.n55 B 0.022551f
C215 VDD2.n56 B 0.022551f
C216 VDD2.n57 B 0.010102f
C217 VDD2.n58 B 0.009541f
C218 VDD2.n59 B 0.017755f
C219 VDD2.n60 B 0.017755f
C220 VDD2.n61 B 0.009541f
C221 VDD2.n62 B 0.010102f
C222 VDD2.n63 B 0.022551f
C223 VDD2.n64 B 0.049243f
C224 VDD2.n65 B 0.010102f
C225 VDD2.n66 B 0.009541f
C226 VDD2.n67 B 0.040555f
C227 VDD2.n68 B 0.444958f
C228 VDD2.n69 B 0.025196f
C229 VDD2.n70 B 0.017755f
C230 VDD2.n71 B 0.009541f
C231 VDD2.n72 B 0.022551f
C232 VDD2.n73 B 0.010102f
C233 VDD2.n74 B 0.017755f
C234 VDD2.n75 B 0.009541f
C235 VDD2.n76 B 0.022551f
C236 VDD2.n77 B 0.010102f
C237 VDD2.n78 B 0.017755f
C238 VDD2.n79 B 0.009541f
C239 VDD2.n80 B 0.022551f
C240 VDD2.n81 B 0.010102f
C241 VDD2.n82 B 0.017755f
C242 VDD2.n83 B 0.009541f
C243 VDD2.n84 B 0.022551f
C244 VDD2.n85 B 0.022551f
C245 VDD2.n86 B 0.010102f
C246 VDD2.n87 B 0.017755f
C247 VDD2.n88 B 0.009541f
C248 VDD2.n89 B 0.022551f
C249 VDD2.n90 B 0.010102f
C250 VDD2.n91 B 0.133601f
C251 VDD2.t1 B 0.038165f
C252 VDD2.n92 B 0.016913f
C253 VDD2.n93 B 0.015942f
C254 VDD2.n94 B 0.009541f
C255 VDD2.n95 B 0.960467f
C256 VDD2.n96 B 0.017755f
C257 VDD2.n97 B 0.009541f
C258 VDD2.n98 B 0.010102f
C259 VDD2.n99 B 0.022551f
C260 VDD2.n100 B 0.022551f
C261 VDD2.n101 B 0.010102f
C262 VDD2.n102 B 0.009541f
C263 VDD2.n103 B 0.017755f
C264 VDD2.n104 B 0.017755f
C265 VDD2.n105 B 0.009541f
C266 VDD2.n106 B 0.010102f
C267 VDD2.n107 B 0.022551f
C268 VDD2.n108 B 0.022551f
C269 VDD2.n109 B 0.010102f
C270 VDD2.n110 B 0.009541f
C271 VDD2.n111 B 0.017755f
C272 VDD2.n112 B 0.017755f
C273 VDD2.n113 B 0.009541f
C274 VDD2.n114 B 0.009821f
C275 VDD2.n115 B 0.009821f
C276 VDD2.n116 B 0.022551f
C277 VDD2.n117 B 0.022551f
C278 VDD2.n118 B 0.010102f
C279 VDD2.n119 B 0.009541f
C280 VDD2.n120 B 0.017755f
C281 VDD2.n121 B 0.017755f
C282 VDD2.n122 B 0.009541f
C283 VDD2.n123 B 0.010102f
C284 VDD2.n124 B 0.022551f
C285 VDD2.n125 B 0.022551f
C286 VDD2.n126 B 0.010102f
C287 VDD2.n127 B 0.009541f
C288 VDD2.n128 B 0.017755f
C289 VDD2.n129 B 0.017755f
C290 VDD2.n130 B 0.009541f
C291 VDD2.n131 B 0.010102f
C292 VDD2.n132 B 0.022551f
C293 VDD2.n133 B 0.049243f
C294 VDD2.n134 B 0.010102f
C295 VDD2.n135 B 0.009541f
C296 VDD2.n136 B 0.040555f
C297 VDD2.n137 B 0.039845f
C298 VDD2.n138 B 1.92273f
C299 VTAIL.n0 B 0.026792f
C300 VTAIL.n1 B 0.01888f
C301 VTAIL.n2 B 0.010145f
C302 VTAIL.n3 B 0.02398f
C303 VTAIL.n4 B 0.010742f
C304 VTAIL.n5 B 0.01888f
C305 VTAIL.n6 B 0.010145f
C306 VTAIL.n7 B 0.02398f
C307 VTAIL.n8 B 0.010742f
C308 VTAIL.n9 B 0.01888f
C309 VTAIL.n10 B 0.010145f
C310 VTAIL.n11 B 0.02398f
C311 VTAIL.n12 B 0.010742f
C312 VTAIL.n13 B 0.01888f
C313 VTAIL.n14 B 0.010145f
C314 VTAIL.n15 B 0.02398f
C315 VTAIL.n16 B 0.010742f
C316 VTAIL.n17 B 0.01888f
C317 VTAIL.n18 B 0.010145f
C318 VTAIL.n19 B 0.02398f
C319 VTAIL.n20 B 0.010742f
C320 VTAIL.n21 B 0.142065f
C321 VTAIL.t1 B 0.040583f
C322 VTAIL.n22 B 0.017985f
C323 VTAIL.n23 B 0.016952f
C324 VTAIL.n24 B 0.010145f
C325 VTAIL.n25 B 1.02132f
C326 VTAIL.n26 B 0.01888f
C327 VTAIL.n27 B 0.010145f
C328 VTAIL.n28 B 0.010742f
C329 VTAIL.n29 B 0.02398f
C330 VTAIL.n30 B 0.02398f
C331 VTAIL.n31 B 0.010742f
C332 VTAIL.n32 B 0.010145f
C333 VTAIL.n33 B 0.01888f
C334 VTAIL.n34 B 0.01888f
C335 VTAIL.n35 B 0.010145f
C336 VTAIL.n36 B 0.010742f
C337 VTAIL.n37 B 0.02398f
C338 VTAIL.n38 B 0.02398f
C339 VTAIL.n39 B 0.02398f
C340 VTAIL.n40 B 0.010742f
C341 VTAIL.n41 B 0.010145f
C342 VTAIL.n42 B 0.01888f
C343 VTAIL.n43 B 0.01888f
C344 VTAIL.n44 B 0.010145f
C345 VTAIL.n45 B 0.010444f
C346 VTAIL.n46 B 0.010444f
C347 VTAIL.n47 B 0.02398f
C348 VTAIL.n48 B 0.02398f
C349 VTAIL.n49 B 0.010742f
C350 VTAIL.n50 B 0.010145f
C351 VTAIL.n51 B 0.01888f
C352 VTAIL.n52 B 0.01888f
C353 VTAIL.n53 B 0.010145f
C354 VTAIL.n54 B 0.010742f
C355 VTAIL.n55 B 0.02398f
C356 VTAIL.n56 B 0.02398f
C357 VTAIL.n57 B 0.010742f
C358 VTAIL.n58 B 0.010145f
C359 VTAIL.n59 B 0.01888f
C360 VTAIL.n60 B 0.01888f
C361 VTAIL.n61 B 0.010145f
C362 VTAIL.n62 B 0.010742f
C363 VTAIL.n63 B 0.02398f
C364 VTAIL.n64 B 0.052362f
C365 VTAIL.n65 B 0.010742f
C366 VTAIL.n66 B 0.010145f
C367 VTAIL.n67 B 0.043124f
C368 VTAIL.n68 B 0.029329f
C369 VTAIL.n69 B 1.06512f
C370 VTAIL.n70 B 0.026792f
C371 VTAIL.n71 B 0.01888f
C372 VTAIL.n72 B 0.010145f
C373 VTAIL.n73 B 0.02398f
C374 VTAIL.n74 B 0.010742f
C375 VTAIL.n75 B 0.01888f
C376 VTAIL.n76 B 0.010145f
C377 VTAIL.n77 B 0.02398f
C378 VTAIL.n78 B 0.010742f
C379 VTAIL.n79 B 0.01888f
C380 VTAIL.n80 B 0.010145f
C381 VTAIL.n81 B 0.02398f
C382 VTAIL.n82 B 0.010742f
C383 VTAIL.n83 B 0.01888f
C384 VTAIL.n84 B 0.010145f
C385 VTAIL.n85 B 0.02398f
C386 VTAIL.n86 B 0.02398f
C387 VTAIL.n87 B 0.010742f
C388 VTAIL.n88 B 0.01888f
C389 VTAIL.n89 B 0.010145f
C390 VTAIL.n90 B 0.02398f
C391 VTAIL.n91 B 0.010742f
C392 VTAIL.n92 B 0.142065f
C393 VTAIL.t2 B 0.040583f
C394 VTAIL.n93 B 0.017985f
C395 VTAIL.n94 B 0.016952f
C396 VTAIL.n95 B 0.010145f
C397 VTAIL.n96 B 1.02132f
C398 VTAIL.n97 B 0.01888f
C399 VTAIL.n98 B 0.010145f
C400 VTAIL.n99 B 0.010742f
C401 VTAIL.n100 B 0.02398f
C402 VTAIL.n101 B 0.02398f
C403 VTAIL.n102 B 0.010742f
C404 VTAIL.n103 B 0.010145f
C405 VTAIL.n104 B 0.01888f
C406 VTAIL.n105 B 0.01888f
C407 VTAIL.n106 B 0.010145f
C408 VTAIL.n107 B 0.010742f
C409 VTAIL.n108 B 0.02398f
C410 VTAIL.n109 B 0.02398f
C411 VTAIL.n110 B 0.010742f
C412 VTAIL.n111 B 0.010145f
C413 VTAIL.n112 B 0.01888f
C414 VTAIL.n113 B 0.01888f
C415 VTAIL.n114 B 0.010145f
C416 VTAIL.n115 B 0.010444f
C417 VTAIL.n116 B 0.010444f
C418 VTAIL.n117 B 0.02398f
C419 VTAIL.n118 B 0.02398f
C420 VTAIL.n119 B 0.010742f
C421 VTAIL.n120 B 0.010145f
C422 VTAIL.n121 B 0.01888f
C423 VTAIL.n122 B 0.01888f
C424 VTAIL.n123 B 0.010145f
C425 VTAIL.n124 B 0.010742f
C426 VTAIL.n125 B 0.02398f
C427 VTAIL.n126 B 0.02398f
C428 VTAIL.n127 B 0.010742f
C429 VTAIL.n128 B 0.010145f
C430 VTAIL.n129 B 0.01888f
C431 VTAIL.n130 B 0.01888f
C432 VTAIL.n131 B 0.010145f
C433 VTAIL.n132 B 0.010742f
C434 VTAIL.n133 B 0.02398f
C435 VTAIL.n134 B 0.052362f
C436 VTAIL.n135 B 0.010742f
C437 VTAIL.n136 B 0.010145f
C438 VTAIL.n137 B 0.043124f
C439 VTAIL.n138 B 0.029329f
C440 VTAIL.n139 B 1.07128f
C441 VTAIL.n140 B 0.026792f
C442 VTAIL.n141 B 0.01888f
C443 VTAIL.n142 B 0.010145f
C444 VTAIL.n143 B 0.02398f
C445 VTAIL.n144 B 0.010742f
C446 VTAIL.n145 B 0.01888f
C447 VTAIL.n146 B 0.010145f
C448 VTAIL.n147 B 0.02398f
C449 VTAIL.n148 B 0.010742f
C450 VTAIL.n149 B 0.01888f
C451 VTAIL.n150 B 0.010145f
C452 VTAIL.n151 B 0.02398f
C453 VTAIL.n152 B 0.010742f
C454 VTAIL.n153 B 0.01888f
C455 VTAIL.n154 B 0.010145f
C456 VTAIL.n155 B 0.02398f
C457 VTAIL.n156 B 0.02398f
C458 VTAIL.n157 B 0.010742f
C459 VTAIL.n158 B 0.01888f
C460 VTAIL.n159 B 0.010145f
C461 VTAIL.n160 B 0.02398f
C462 VTAIL.n161 B 0.010742f
C463 VTAIL.n162 B 0.142065f
C464 VTAIL.t0 B 0.040583f
C465 VTAIL.n163 B 0.017985f
C466 VTAIL.n164 B 0.016952f
C467 VTAIL.n165 B 0.010145f
C468 VTAIL.n166 B 1.02132f
C469 VTAIL.n167 B 0.01888f
C470 VTAIL.n168 B 0.010145f
C471 VTAIL.n169 B 0.010742f
C472 VTAIL.n170 B 0.02398f
C473 VTAIL.n171 B 0.02398f
C474 VTAIL.n172 B 0.010742f
C475 VTAIL.n173 B 0.010145f
C476 VTAIL.n174 B 0.01888f
C477 VTAIL.n175 B 0.01888f
C478 VTAIL.n176 B 0.010145f
C479 VTAIL.n177 B 0.010742f
C480 VTAIL.n178 B 0.02398f
C481 VTAIL.n179 B 0.02398f
C482 VTAIL.n180 B 0.010742f
C483 VTAIL.n181 B 0.010145f
C484 VTAIL.n182 B 0.01888f
C485 VTAIL.n183 B 0.01888f
C486 VTAIL.n184 B 0.010145f
C487 VTAIL.n185 B 0.010444f
C488 VTAIL.n186 B 0.010444f
C489 VTAIL.n187 B 0.02398f
C490 VTAIL.n188 B 0.02398f
C491 VTAIL.n189 B 0.010742f
C492 VTAIL.n190 B 0.010145f
C493 VTAIL.n191 B 0.01888f
C494 VTAIL.n192 B 0.01888f
C495 VTAIL.n193 B 0.010145f
C496 VTAIL.n194 B 0.010742f
C497 VTAIL.n195 B 0.02398f
C498 VTAIL.n196 B 0.02398f
C499 VTAIL.n197 B 0.010742f
C500 VTAIL.n198 B 0.010145f
C501 VTAIL.n199 B 0.01888f
C502 VTAIL.n200 B 0.01888f
C503 VTAIL.n201 B 0.010145f
C504 VTAIL.n202 B 0.010742f
C505 VTAIL.n203 B 0.02398f
C506 VTAIL.n204 B 0.052362f
C507 VTAIL.n205 B 0.010742f
C508 VTAIL.n206 B 0.010145f
C509 VTAIL.n207 B 0.043124f
C510 VTAIL.n208 B 0.029329f
C511 VTAIL.n209 B 1.03247f
C512 VTAIL.n210 B 0.026792f
C513 VTAIL.n211 B 0.01888f
C514 VTAIL.n212 B 0.010145f
C515 VTAIL.n213 B 0.02398f
C516 VTAIL.n214 B 0.010742f
C517 VTAIL.n215 B 0.01888f
C518 VTAIL.n216 B 0.010145f
C519 VTAIL.n217 B 0.02398f
C520 VTAIL.n218 B 0.010742f
C521 VTAIL.n219 B 0.01888f
C522 VTAIL.n220 B 0.010145f
C523 VTAIL.n221 B 0.02398f
C524 VTAIL.n222 B 0.010742f
C525 VTAIL.n223 B 0.01888f
C526 VTAIL.n224 B 0.010145f
C527 VTAIL.n225 B 0.02398f
C528 VTAIL.n226 B 0.010742f
C529 VTAIL.n227 B 0.01888f
C530 VTAIL.n228 B 0.010145f
C531 VTAIL.n229 B 0.02398f
C532 VTAIL.n230 B 0.010742f
C533 VTAIL.n231 B 0.142065f
C534 VTAIL.t3 B 0.040583f
C535 VTAIL.n232 B 0.017985f
C536 VTAIL.n233 B 0.016952f
C537 VTAIL.n234 B 0.010145f
C538 VTAIL.n235 B 1.02132f
C539 VTAIL.n236 B 0.01888f
C540 VTAIL.n237 B 0.010145f
C541 VTAIL.n238 B 0.010742f
C542 VTAIL.n239 B 0.02398f
C543 VTAIL.n240 B 0.02398f
C544 VTAIL.n241 B 0.010742f
C545 VTAIL.n242 B 0.010145f
C546 VTAIL.n243 B 0.01888f
C547 VTAIL.n244 B 0.01888f
C548 VTAIL.n245 B 0.010145f
C549 VTAIL.n246 B 0.010742f
C550 VTAIL.n247 B 0.02398f
C551 VTAIL.n248 B 0.02398f
C552 VTAIL.n249 B 0.02398f
C553 VTAIL.n250 B 0.010742f
C554 VTAIL.n251 B 0.010145f
C555 VTAIL.n252 B 0.01888f
C556 VTAIL.n253 B 0.01888f
C557 VTAIL.n254 B 0.010145f
C558 VTAIL.n255 B 0.010444f
C559 VTAIL.n256 B 0.010444f
C560 VTAIL.n257 B 0.02398f
C561 VTAIL.n258 B 0.02398f
C562 VTAIL.n259 B 0.010742f
C563 VTAIL.n260 B 0.010145f
C564 VTAIL.n261 B 0.01888f
C565 VTAIL.n262 B 0.01888f
C566 VTAIL.n263 B 0.010145f
C567 VTAIL.n264 B 0.010742f
C568 VTAIL.n265 B 0.02398f
C569 VTAIL.n266 B 0.02398f
C570 VTAIL.n267 B 0.010742f
C571 VTAIL.n268 B 0.010145f
C572 VTAIL.n269 B 0.01888f
C573 VTAIL.n270 B 0.01888f
C574 VTAIL.n271 B 0.010145f
C575 VTAIL.n272 B 0.010742f
C576 VTAIL.n273 B 0.02398f
C577 VTAIL.n274 B 0.052362f
C578 VTAIL.n275 B 0.010742f
C579 VTAIL.n276 B 0.010145f
C580 VTAIL.n277 B 0.043124f
C581 VTAIL.n278 B 0.029329f
C582 VTAIL.n279 B 0.990649f
C583 VN.t1 B 0.61951f
C584 VN.t0 B 0.682456f
.ends

