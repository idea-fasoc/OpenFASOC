* NGSPICE file created from diff_pair_sample_0215.ext - technology: sky130A

.subckt diff_pair_sample_0215 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t7 VP.t0 VTAIL.t11 B.t1 sky130_fd_pr__nfet_01v8 ad=1.4025 pd=8.83 as=3.315 ps=17.78 w=8.5 l=1.95
X1 VDD2.t7 VN.t0 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.4025 pd=8.83 as=1.4025 ps=8.83 w=8.5 l=1.95
X2 VDD2.t6 VN.t1 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=1.4025 pd=8.83 as=3.315 ps=17.78 w=8.5 l=1.95
X3 VDD1.t6 VP.t1 VTAIL.t13 B.t3 sky130_fd_pr__nfet_01v8 ad=1.4025 pd=8.83 as=1.4025 ps=8.83 w=8.5 l=1.95
X4 VDD1.t5 VP.t2 VTAIL.t9 B.t4 sky130_fd_pr__nfet_01v8 ad=1.4025 pd=8.83 as=1.4025 ps=8.83 w=8.5 l=1.95
X5 VTAIL.t7 VN.t2 VDD2.t5 B.t7 sky130_fd_pr__nfet_01v8 ad=3.315 pd=17.78 as=1.4025 ps=8.83 w=8.5 l=1.95
X6 VTAIL.t2 VN.t3 VDD2.t4 B.t2 sky130_fd_pr__nfet_01v8 ad=1.4025 pd=8.83 as=1.4025 ps=8.83 w=8.5 l=1.95
X7 B.t21 B.t19 B.t20 B.t9 sky130_fd_pr__nfet_01v8 ad=3.315 pd=17.78 as=0 ps=0 w=8.5 l=1.95
X8 VDD1.t4 VP.t3 VTAIL.t10 B.t6 sky130_fd_pr__nfet_01v8 ad=1.4025 pd=8.83 as=3.315 ps=17.78 w=8.5 l=1.95
X9 VTAIL.t0 VN.t4 VDD2.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=1.4025 pd=8.83 as=1.4025 ps=8.83 w=8.5 l=1.95
X10 VTAIL.t12 VP.t4 VDD1.t3 B.t7 sky130_fd_pr__nfet_01v8 ad=3.315 pd=17.78 as=1.4025 ps=8.83 w=8.5 l=1.95
X11 B.t18 B.t16 B.t17 B.t13 sky130_fd_pr__nfet_01v8 ad=3.315 pd=17.78 as=0 ps=0 w=8.5 l=1.95
X12 VDD2.t2 VN.t5 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.4025 pd=8.83 as=3.315 ps=17.78 w=8.5 l=1.95
X13 VTAIL.t14 VP.t5 VDD1.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.4025 pd=8.83 as=1.4025 ps=8.83 w=8.5 l=1.95
X14 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=3.315 pd=17.78 as=0 ps=0 w=8.5 l=1.95
X15 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=3.315 pd=17.78 as=0 ps=0 w=8.5 l=1.95
X16 VDD2.t1 VN.t6 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.4025 pd=8.83 as=1.4025 ps=8.83 w=8.5 l=1.95
X17 VTAIL.t15 VP.t6 VDD1.t1 B.t5 sky130_fd_pr__nfet_01v8 ad=3.315 pd=17.78 as=1.4025 ps=8.83 w=8.5 l=1.95
X18 VTAIL.t8 VP.t7 VDD1.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.4025 pd=8.83 as=1.4025 ps=8.83 w=8.5 l=1.95
X19 VTAIL.t5 VN.t7 VDD2.t0 B.t5 sky130_fd_pr__nfet_01v8 ad=3.315 pd=17.78 as=1.4025 ps=8.83 w=8.5 l=1.95
R0 VP.n14 VP.n11 161.3
R1 VP.n16 VP.n15 161.3
R2 VP.n17 VP.n10 161.3
R3 VP.n19 VP.n18 161.3
R4 VP.n20 VP.n9 161.3
R5 VP.n23 VP.n22 161.3
R6 VP.n24 VP.n8 161.3
R7 VP.n26 VP.n25 161.3
R8 VP.n27 VP.n7 161.3
R9 VP.n52 VP.n0 161.3
R10 VP.n51 VP.n50 161.3
R11 VP.n49 VP.n1 161.3
R12 VP.n48 VP.n47 161.3
R13 VP.n45 VP.n2 161.3
R14 VP.n44 VP.n43 161.3
R15 VP.n42 VP.n3 161.3
R16 VP.n41 VP.n40 161.3
R17 VP.n39 VP.n4 161.3
R18 VP.n37 VP.n36 161.3
R19 VP.n35 VP.n5 161.3
R20 VP.n34 VP.n33 161.3
R21 VP.n32 VP.n6 161.3
R22 VP.n12 VP.t4 135.59
R23 VP.n31 VP.t6 105.052
R24 VP.n38 VP.t2 105.052
R25 VP.n46 VP.t5 105.052
R26 VP.n53 VP.t0 105.052
R27 VP.n28 VP.t3 105.052
R28 VP.n21 VP.t7 105.052
R29 VP.n13 VP.t1 105.052
R30 VP.n31 VP.n30 90.2511
R31 VP.n54 VP.n53 90.2511
R32 VP.n29 VP.n28 90.2511
R33 VP.n13 VP.n12 63.2137
R34 VP.n33 VP.n5 56.5617
R35 VP.n51 VP.n1 56.5617
R36 VP.n26 VP.n8 56.5617
R37 VP.n30 VP.n29 45.2269
R38 VP.n40 VP.n3 40.577
R39 VP.n44 VP.n3 40.577
R40 VP.n19 VP.n10 40.577
R41 VP.n15 VP.n10 40.577
R42 VP.n33 VP.n32 24.5923
R43 VP.n37 VP.n5 24.5923
R44 VP.n40 VP.n39 24.5923
R45 VP.n45 VP.n44 24.5923
R46 VP.n47 VP.n1 24.5923
R47 VP.n52 VP.n51 24.5923
R48 VP.n27 VP.n26 24.5923
R49 VP.n20 VP.n19 24.5923
R50 VP.n22 VP.n8 24.5923
R51 VP.n15 VP.n14 24.5923
R52 VP.n32 VP.n31 20.6576
R53 VP.n53 VP.n52 20.6576
R54 VP.n28 VP.n27 20.6576
R55 VP.n38 VP.n37 17.7066
R56 VP.n47 VP.n46 17.7066
R57 VP.n22 VP.n21 17.7066
R58 VP.n12 VP.n11 13.203
R59 VP.n39 VP.n38 6.88621
R60 VP.n46 VP.n45 6.88621
R61 VP.n21 VP.n20 6.88621
R62 VP.n14 VP.n13 6.88621
R63 VP.n29 VP.n7 0.278335
R64 VP.n30 VP.n6 0.278335
R65 VP.n54 VP.n0 0.278335
R66 VP.n16 VP.n11 0.189894
R67 VP.n17 VP.n16 0.189894
R68 VP.n18 VP.n17 0.189894
R69 VP.n18 VP.n9 0.189894
R70 VP.n23 VP.n9 0.189894
R71 VP.n24 VP.n23 0.189894
R72 VP.n25 VP.n24 0.189894
R73 VP.n25 VP.n7 0.189894
R74 VP.n34 VP.n6 0.189894
R75 VP.n35 VP.n34 0.189894
R76 VP.n36 VP.n35 0.189894
R77 VP.n36 VP.n4 0.189894
R78 VP.n41 VP.n4 0.189894
R79 VP.n42 VP.n41 0.189894
R80 VP.n43 VP.n42 0.189894
R81 VP.n43 VP.n2 0.189894
R82 VP.n48 VP.n2 0.189894
R83 VP.n49 VP.n48 0.189894
R84 VP.n50 VP.n49 0.189894
R85 VP.n50 VP.n0 0.189894
R86 VP VP.n54 0.153485
R87 VTAIL.n11 VTAIL.t12 49.4688
R88 VTAIL.n10 VTAIL.t1 49.4688
R89 VTAIL.n7 VTAIL.t5 49.4688
R90 VTAIL.n14 VTAIL.t10 49.4688
R91 VTAIL.n15 VTAIL.t6 49.4686
R92 VTAIL.n2 VTAIL.t7 49.4686
R93 VTAIL.n3 VTAIL.t11 49.4686
R94 VTAIL.n6 VTAIL.t15 49.4686
R95 VTAIL.n13 VTAIL.n12 47.1394
R96 VTAIL.n9 VTAIL.n8 47.1394
R97 VTAIL.n1 VTAIL.n0 47.1394
R98 VTAIL.n5 VTAIL.n4 47.1394
R99 VTAIL.n15 VTAIL.n14 21.66
R100 VTAIL.n7 VTAIL.n6 21.66
R101 VTAIL.n0 VTAIL.t3 2.32991
R102 VTAIL.n0 VTAIL.t0 2.32991
R103 VTAIL.n4 VTAIL.t9 2.32991
R104 VTAIL.n4 VTAIL.t14 2.32991
R105 VTAIL.n12 VTAIL.t13 2.32991
R106 VTAIL.n12 VTAIL.t8 2.32991
R107 VTAIL.n8 VTAIL.t4 2.32991
R108 VTAIL.n8 VTAIL.t2 2.32991
R109 VTAIL.n9 VTAIL.n7 1.96602
R110 VTAIL.n10 VTAIL.n9 1.96602
R111 VTAIL.n13 VTAIL.n11 1.96602
R112 VTAIL.n14 VTAIL.n13 1.96602
R113 VTAIL.n6 VTAIL.n5 1.96602
R114 VTAIL.n5 VTAIL.n3 1.96602
R115 VTAIL.n2 VTAIL.n1 1.96602
R116 VTAIL VTAIL.n15 1.90783
R117 VTAIL.n11 VTAIL.n10 0.470328
R118 VTAIL.n3 VTAIL.n2 0.470328
R119 VTAIL VTAIL.n1 0.0586897
R120 VDD1 VDD1.n0 64.8591
R121 VDD1.n3 VDD1.n2 64.7456
R122 VDD1.n3 VDD1.n1 64.7456
R123 VDD1.n5 VDD1.n4 63.8182
R124 VDD1.n5 VDD1.n3 40.4707
R125 VDD1.n4 VDD1.t0 2.32991
R126 VDD1.n4 VDD1.t4 2.32991
R127 VDD1.n0 VDD1.t3 2.32991
R128 VDD1.n0 VDD1.t6 2.32991
R129 VDD1.n2 VDD1.t2 2.32991
R130 VDD1.n2 VDD1.t7 2.32991
R131 VDD1.n1 VDD1.t1 2.32991
R132 VDD1.n1 VDD1.t5 2.32991
R133 VDD1 VDD1.n5 0.925069
R134 B.n704 B.n703 585
R135 B.n260 B.n113 585
R136 B.n259 B.n258 585
R137 B.n257 B.n256 585
R138 B.n255 B.n254 585
R139 B.n253 B.n252 585
R140 B.n251 B.n250 585
R141 B.n249 B.n248 585
R142 B.n247 B.n246 585
R143 B.n245 B.n244 585
R144 B.n243 B.n242 585
R145 B.n241 B.n240 585
R146 B.n239 B.n238 585
R147 B.n237 B.n236 585
R148 B.n235 B.n234 585
R149 B.n233 B.n232 585
R150 B.n231 B.n230 585
R151 B.n229 B.n228 585
R152 B.n227 B.n226 585
R153 B.n225 B.n224 585
R154 B.n223 B.n222 585
R155 B.n221 B.n220 585
R156 B.n219 B.n218 585
R157 B.n217 B.n216 585
R158 B.n215 B.n214 585
R159 B.n213 B.n212 585
R160 B.n211 B.n210 585
R161 B.n209 B.n208 585
R162 B.n207 B.n206 585
R163 B.n205 B.n204 585
R164 B.n203 B.n202 585
R165 B.n200 B.n199 585
R166 B.n198 B.n197 585
R167 B.n196 B.n195 585
R168 B.n194 B.n193 585
R169 B.n192 B.n191 585
R170 B.n190 B.n189 585
R171 B.n188 B.n187 585
R172 B.n186 B.n185 585
R173 B.n184 B.n183 585
R174 B.n182 B.n181 585
R175 B.n179 B.n178 585
R176 B.n177 B.n176 585
R177 B.n175 B.n174 585
R178 B.n173 B.n172 585
R179 B.n171 B.n170 585
R180 B.n169 B.n168 585
R181 B.n167 B.n166 585
R182 B.n165 B.n164 585
R183 B.n163 B.n162 585
R184 B.n161 B.n160 585
R185 B.n159 B.n158 585
R186 B.n157 B.n156 585
R187 B.n155 B.n154 585
R188 B.n153 B.n152 585
R189 B.n151 B.n150 585
R190 B.n149 B.n148 585
R191 B.n147 B.n146 585
R192 B.n145 B.n144 585
R193 B.n143 B.n142 585
R194 B.n141 B.n140 585
R195 B.n139 B.n138 585
R196 B.n137 B.n136 585
R197 B.n135 B.n134 585
R198 B.n133 B.n132 585
R199 B.n131 B.n130 585
R200 B.n129 B.n128 585
R201 B.n127 B.n126 585
R202 B.n125 B.n124 585
R203 B.n123 B.n122 585
R204 B.n121 B.n120 585
R205 B.n119 B.n118 585
R206 B.n702 B.n77 585
R207 B.n707 B.n77 585
R208 B.n701 B.n76 585
R209 B.n708 B.n76 585
R210 B.n700 B.n699 585
R211 B.n699 B.n72 585
R212 B.n698 B.n71 585
R213 B.n714 B.n71 585
R214 B.n697 B.n70 585
R215 B.n715 B.n70 585
R216 B.n696 B.n69 585
R217 B.n716 B.n69 585
R218 B.n695 B.n694 585
R219 B.n694 B.n68 585
R220 B.n693 B.n64 585
R221 B.n722 B.n64 585
R222 B.n692 B.n63 585
R223 B.n723 B.n63 585
R224 B.n691 B.n62 585
R225 B.n724 B.n62 585
R226 B.n690 B.n689 585
R227 B.n689 B.n58 585
R228 B.n688 B.n57 585
R229 B.n730 B.n57 585
R230 B.n687 B.n56 585
R231 B.n731 B.n56 585
R232 B.n686 B.n55 585
R233 B.n732 B.n55 585
R234 B.n685 B.n684 585
R235 B.n684 B.n51 585
R236 B.n683 B.n50 585
R237 B.n738 B.n50 585
R238 B.n682 B.n49 585
R239 B.n739 B.n49 585
R240 B.n681 B.n48 585
R241 B.n740 B.n48 585
R242 B.n680 B.n679 585
R243 B.n679 B.n44 585
R244 B.n678 B.n43 585
R245 B.n746 B.n43 585
R246 B.n677 B.n42 585
R247 B.n747 B.n42 585
R248 B.n676 B.n41 585
R249 B.n748 B.n41 585
R250 B.n675 B.n674 585
R251 B.n674 B.n37 585
R252 B.n673 B.n36 585
R253 B.n754 B.n36 585
R254 B.n672 B.n35 585
R255 B.n755 B.n35 585
R256 B.n671 B.n34 585
R257 B.n756 B.n34 585
R258 B.n670 B.n669 585
R259 B.n669 B.n30 585
R260 B.n668 B.n29 585
R261 B.n762 B.n29 585
R262 B.n667 B.n28 585
R263 B.n763 B.n28 585
R264 B.n666 B.n27 585
R265 B.n764 B.n27 585
R266 B.n665 B.n664 585
R267 B.n664 B.n23 585
R268 B.n663 B.n22 585
R269 B.n770 B.n22 585
R270 B.n662 B.n21 585
R271 B.n771 B.n21 585
R272 B.n661 B.n20 585
R273 B.n772 B.n20 585
R274 B.n660 B.n659 585
R275 B.n659 B.n16 585
R276 B.n658 B.n15 585
R277 B.n778 B.n15 585
R278 B.n657 B.n14 585
R279 B.n779 B.n14 585
R280 B.n656 B.n13 585
R281 B.n780 B.n13 585
R282 B.n655 B.n654 585
R283 B.n654 B.n12 585
R284 B.n653 B.n652 585
R285 B.n653 B.n8 585
R286 B.n651 B.n7 585
R287 B.n787 B.n7 585
R288 B.n650 B.n6 585
R289 B.n788 B.n6 585
R290 B.n649 B.n5 585
R291 B.n789 B.n5 585
R292 B.n648 B.n647 585
R293 B.n647 B.n4 585
R294 B.n646 B.n261 585
R295 B.n646 B.n645 585
R296 B.n636 B.n262 585
R297 B.n263 B.n262 585
R298 B.n638 B.n637 585
R299 B.n639 B.n638 585
R300 B.n635 B.n267 585
R301 B.n271 B.n267 585
R302 B.n634 B.n633 585
R303 B.n633 B.n632 585
R304 B.n269 B.n268 585
R305 B.n270 B.n269 585
R306 B.n625 B.n624 585
R307 B.n626 B.n625 585
R308 B.n623 B.n276 585
R309 B.n276 B.n275 585
R310 B.n622 B.n621 585
R311 B.n621 B.n620 585
R312 B.n278 B.n277 585
R313 B.n279 B.n278 585
R314 B.n613 B.n612 585
R315 B.n614 B.n613 585
R316 B.n611 B.n284 585
R317 B.n284 B.n283 585
R318 B.n610 B.n609 585
R319 B.n609 B.n608 585
R320 B.n286 B.n285 585
R321 B.n287 B.n286 585
R322 B.n601 B.n600 585
R323 B.n602 B.n601 585
R324 B.n599 B.n292 585
R325 B.n292 B.n291 585
R326 B.n598 B.n597 585
R327 B.n597 B.n596 585
R328 B.n294 B.n293 585
R329 B.n295 B.n294 585
R330 B.n589 B.n588 585
R331 B.n590 B.n589 585
R332 B.n587 B.n300 585
R333 B.n300 B.n299 585
R334 B.n586 B.n585 585
R335 B.n585 B.n584 585
R336 B.n302 B.n301 585
R337 B.n303 B.n302 585
R338 B.n577 B.n576 585
R339 B.n578 B.n577 585
R340 B.n575 B.n307 585
R341 B.n311 B.n307 585
R342 B.n574 B.n573 585
R343 B.n573 B.n572 585
R344 B.n309 B.n308 585
R345 B.n310 B.n309 585
R346 B.n565 B.n564 585
R347 B.n566 B.n565 585
R348 B.n563 B.n316 585
R349 B.n316 B.n315 585
R350 B.n562 B.n561 585
R351 B.n561 B.n560 585
R352 B.n318 B.n317 585
R353 B.n319 B.n318 585
R354 B.n553 B.n552 585
R355 B.n554 B.n553 585
R356 B.n551 B.n324 585
R357 B.n324 B.n323 585
R358 B.n550 B.n549 585
R359 B.n549 B.n548 585
R360 B.n326 B.n325 585
R361 B.n541 B.n326 585
R362 B.n540 B.n539 585
R363 B.n542 B.n540 585
R364 B.n538 B.n331 585
R365 B.n331 B.n330 585
R366 B.n537 B.n536 585
R367 B.n536 B.n535 585
R368 B.n333 B.n332 585
R369 B.n334 B.n333 585
R370 B.n528 B.n527 585
R371 B.n529 B.n528 585
R372 B.n526 B.n339 585
R373 B.n339 B.n338 585
R374 B.n521 B.n520 585
R375 B.n519 B.n377 585
R376 B.n518 B.n376 585
R377 B.n523 B.n376 585
R378 B.n517 B.n516 585
R379 B.n515 B.n514 585
R380 B.n513 B.n512 585
R381 B.n511 B.n510 585
R382 B.n509 B.n508 585
R383 B.n507 B.n506 585
R384 B.n505 B.n504 585
R385 B.n503 B.n502 585
R386 B.n501 B.n500 585
R387 B.n499 B.n498 585
R388 B.n497 B.n496 585
R389 B.n495 B.n494 585
R390 B.n493 B.n492 585
R391 B.n491 B.n490 585
R392 B.n489 B.n488 585
R393 B.n487 B.n486 585
R394 B.n485 B.n484 585
R395 B.n483 B.n482 585
R396 B.n481 B.n480 585
R397 B.n479 B.n478 585
R398 B.n477 B.n476 585
R399 B.n475 B.n474 585
R400 B.n473 B.n472 585
R401 B.n471 B.n470 585
R402 B.n469 B.n468 585
R403 B.n467 B.n466 585
R404 B.n465 B.n464 585
R405 B.n463 B.n462 585
R406 B.n461 B.n460 585
R407 B.n459 B.n458 585
R408 B.n457 B.n456 585
R409 B.n455 B.n454 585
R410 B.n453 B.n452 585
R411 B.n451 B.n450 585
R412 B.n449 B.n448 585
R413 B.n447 B.n446 585
R414 B.n445 B.n444 585
R415 B.n443 B.n442 585
R416 B.n441 B.n440 585
R417 B.n439 B.n438 585
R418 B.n437 B.n436 585
R419 B.n435 B.n434 585
R420 B.n433 B.n432 585
R421 B.n431 B.n430 585
R422 B.n429 B.n428 585
R423 B.n427 B.n426 585
R424 B.n425 B.n424 585
R425 B.n423 B.n422 585
R426 B.n421 B.n420 585
R427 B.n419 B.n418 585
R428 B.n417 B.n416 585
R429 B.n415 B.n414 585
R430 B.n413 B.n412 585
R431 B.n411 B.n410 585
R432 B.n409 B.n408 585
R433 B.n407 B.n406 585
R434 B.n405 B.n404 585
R435 B.n403 B.n402 585
R436 B.n401 B.n400 585
R437 B.n399 B.n398 585
R438 B.n397 B.n396 585
R439 B.n395 B.n394 585
R440 B.n393 B.n392 585
R441 B.n391 B.n390 585
R442 B.n389 B.n388 585
R443 B.n387 B.n386 585
R444 B.n385 B.n384 585
R445 B.n341 B.n340 585
R446 B.n525 B.n524 585
R447 B.n524 B.n523 585
R448 B.n337 B.n336 585
R449 B.n338 B.n337 585
R450 B.n531 B.n530 585
R451 B.n530 B.n529 585
R452 B.n532 B.n335 585
R453 B.n335 B.n334 585
R454 B.n534 B.n533 585
R455 B.n535 B.n534 585
R456 B.n329 B.n328 585
R457 B.n330 B.n329 585
R458 B.n544 B.n543 585
R459 B.n543 B.n542 585
R460 B.n545 B.n327 585
R461 B.n541 B.n327 585
R462 B.n547 B.n546 585
R463 B.n548 B.n547 585
R464 B.n322 B.n321 585
R465 B.n323 B.n322 585
R466 B.n556 B.n555 585
R467 B.n555 B.n554 585
R468 B.n557 B.n320 585
R469 B.n320 B.n319 585
R470 B.n559 B.n558 585
R471 B.n560 B.n559 585
R472 B.n314 B.n313 585
R473 B.n315 B.n314 585
R474 B.n568 B.n567 585
R475 B.n567 B.n566 585
R476 B.n569 B.n312 585
R477 B.n312 B.n310 585
R478 B.n571 B.n570 585
R479 B.n572 B.n571 585
R480 B.n306 B.n305 585
R481 B.n311 B.n306 585
R482 B.n580 B.n579 585
R483 B.n579 B.n578 585
R484 B.n581 B.n304 585
R485 B.n304 B.n303 585
R486 B.n583 B.n582 585
R487 B.n584 B.n583 585
R488 B.n298 B.n297 585
R489 B.n299 B.n298 585
R490 B.n592 B.n591 585
R491 B.n591 B.n590 585
R492 B.n593 B.n296 585
R493 B.n296 B.n295 585
R494 B.n595 B.n594 585
R495 B.n596 B.n595 585
R496 B.n290 B.n289 585
R497 B.n291 B.n290 585
R498 B.n604 B.n603 585
R499 B.n603 B.n602 585
R500 B.n605 B.n288 585
R501 B.n288 B.n287 585
R502 B.n607 B.n606 585
R503 B.n608 B.n607 585
R504 B.n282 B.n281 585
R505 B.n283 B.n282 585
R506 B.n616 B.n615 585
R507 B.n615 B.n614 585
R508 B.n617 B.n280 585
R509 B.n280 B.n279 585
R510 B.n619 B.n618 585
R511 B.n620 B.n619 585
R512 B.n274 B.n273 585
R513 B.n275 B.n274 585
R514 B.n628 B.n627 585
R515 B.n627 B.n626 585
R516 B.n629 B.n272 585
R517 B.n272 B.n270 585
R518 B.n631 B.n630 585
R519 B.n632 B.n631 585
R520 B.n266 B.n265 585
R521 B.n271 B.n266 585
R522 B.n641 B.n640 585
R523 B.n640 B.n639 585
R524 B.n642 B.n264 585
R525 B.n264 B.n263 585
R526 B.n644 B.n643 585
R527 B.n645 B.n644 585
R528 B.n3 B.n0 585
R529 B.n4 B.n3 585
R530 B.n786 B.n1 585
R531 B.n787 B.n786 585
R532 B.n785 B.n784 585
R533 B.n785 B.n8 585
R534 B.n783 B.n9 585
R535 B.n12 B.n9 585
R536 B.n782 B.n781 585
R537 B.n781 B.n780 585
R538 B.n11 B.n10 585
R539 B.n779 B.n11 585
R540 B.n777 B.n776 585
R541 B.n778 B.n777 585
R542 B.n775 B.n17 585
R543 B.n17 B.n16 585
R544 B.n774 B.n773 585
R545 B.n773 B.n772 585
R546 B.n19 B.n18 585
R547 B.n771 B.n19 585
R548 B.n769 B.n768 585
R549 B.n770 B.n769 585
R550 B.n767 B.n24 585
R551 B.n24 B.n23 585
R552 B.n766 B.n765 585
R553 B.n765 B.n764 585
R554 B.n26 B.n25 585
R555 B.n763 B.n26 585
R556 B.n761 B.n760 585
R557 B.n762 B.n761 585
R558 B.n759 B.n31 585
R559 B.n31 B.n30 585
R560 B.n758 B.n757 585
R561 B.n757 B.n756 585
R562 B.n33 B.n32 585
R563 B.n755 B.n33 585
R564 B.n753 B.n752 585
R565 B.n754 B.n753 585
R566 B.n751 B.n38 585
R567 B.n38 B.n37 585
R568 B.n750 B.n749 585
R569 B.n749 B.n748 585
R570 B.n40 B.n39 585
R571 B.n747 B.n40 585
R572 B.n745 B.n744 585
R573 B.n746 B.n745 585
R574 B.n743 B.n45 585
R575 B.n45 B.n44 585
R576 B.n742 B.n741 585
R577 B.n741 B.n740 585
R578 B.n47 B.n46 585
R579 B.n739 B.n47 585
R580 B.n737 B.n736 585
R581 B.n738 B.n737 585
R582 B.n735 B.n52 585
R583 B.n52 B.n51 585
R584 B.n734 B.n733 585
R585 B.n733 B.n732 585
R586 B.n54 B.n53 585
R587 B.n731 B.n54 585
R588 B.n729 B.n728 585
R589 B.n730 B.n729 585
R590 B.n727 B.n59 585
R591 B.n59 B.n58 585
R592 B.n726 B.n725 585
R593 B.n725 B.n724 585
R594 B.n61 B.n60 585
R595 B.n723 B.n61 585
R596 B.n721 B.n720 585
R597 B.n722 B.n721 585
R598 B.n719 B.n65 585
R599 B.n68 B.n65 585
R600 B.n718 B.n717 585
R601 B.n717 B.n716 585
R602 B.n67 B.n66 585
R603 B.n715 B.n67 585
R604 B.n713 B.n712 585
R605 B.n714 B.n713 585
R606 B.n711 B.n73 585
R607 B.n73 B.n72 585
R608 B.n710 B.n709 585
R609 B.n709 B.n708 585
R610 B.n75 B.n74 585
R611 B.n707 B.n75 585
R612 B.n790 B.n789 585
R613 B.n788 B.n2 585
R614 B.n118 B.n75 540.549
R615 B.n704 B.n77 540.549
R616 B.n524 B.n339 540.549
R617 B.n521 B.n337 540.549
R618 B.n116 B.t16 311.849
R619 B.n114 B.t12 311.849
R620 B.n381 B.t19 311.849
R621 B.n378 B.t8 311.849
R622 B.n706 B.n705 256.663
R623 B.n706 B.n112 256.663
R624 B.n706 B.n111 256.663
R625 B.n706 B.n110 256.663
R626 B.n706 B.n109 256.663
R627 B.n706 B.n108 256.663
R628 B.n706 B.n107 256.663
R629 B.n706 B.n106 256.663
R630 B.n706 B.n105 256.663
R631 B.n706 B.n104 256.663
R632 B.n706 B.n103 256.663
R633 B.n706 B.n102 256.663
R634 B.n706 B.n101 256.663
R635 B.n706 B.n100 256.663
R636 B.n706 B.n99 256.663
R637 B.n706 B.n98 256.663
R638 B.n706 B.n97 256.663
R639 B.n706 B.n96 256.663
R640 B.n706 B.n95 256.663
R641 B.n706 B.n94 256.663
R642 B.n706 B.n93 256.663
R643 B.n706 B.n92 256.663
R644 B.n706 B.n91 256.663
R645 B.n706 B.n90 256.663
R646 B.n706 B.n89 256.663
R647 B.n706 B.n88 256.663
R648 B.n706 B.n87 256.663
R649 B.n706 B.n86 256.663
R650 B.n706 B.n85 256.663
R651 B.n706 B.n84 256.663
R652 B.n706 B.n83 256.663
R653 B.n706 B.n82 256.663
R654 B.n706 B.n81 256.663
R655 B.n706 B.n80 256.663
R656 B.n706 B.n79 256.663
R657 B.n706 B.n78 256.663
R658 B.n523 B.n522 256.663
R659 B.n523 B.n342 256.663
R660 B.n523 B.n343 256.663
R661 B.n523 B.n344 256.663
R662 B.n523 B.n345 256.663
R663 B.n523 B.n346 256.663
R664 B.n523 B.n347 256.663
R665 B.n523 B.n348 256.663
R666 B.n523 B.n349 256.663
R667 B.n523 B.n350 256.663
R668 B.n523 B.n351 256.663
R669 B.n523 B.n352 256.663
R670 B.n523 B.n353 256.663
R671 B.n523 B.n354 256.663
R672 B.n523 B.n355 256.663
R673 B.n523 B.n356 256.663
R674 B.n523 B.n357 256.663
R675 B.n523 B.n358 256.663
R676 B.n523 B.n359 256.663
R677 B.n523 B.n360 256.663
R678 B.n523 B.n361 256.663
R679 B.n523 B.n362 256.663
R680 B.n523 B.n363 256.663
R681 B.n523 B.n364 256.663
R682 B.n523 B.n365 256.663
R683 B.n523 B.n366 256.663
R684 B.n523 B.n367 256.663
R685 B.n523 B.n368 256.663
R686 B.n523 B.n369 256.663
R687 B.n523 B.n370 256.663
R688 B.n523 B.n371 256.663
R689 B.n523 B.n372 256.663
R690 B.n523 B.n373 256.663
R691 B.n523 B.n374 256.663
R692 B.n523 B.n375 256.663
R693 B.n792 B.n791 256.663
R694 B.n122 B.n121 163.367
R695 B.n126 B.n125 163.367
R696 B.n130 B.n129 163.367
R697 B.n134 B.n133 163.367
R698 B.n138 B.n137 163.367
R699 B.n142 B.n141 163.367
R700 B.n146 B.n145 163.367
R701 B.n150 B.n149 163.367
R702 B.n154 B.n153 163.367
R703 B.n158 B.n157 163.367
R704 B.n162 B.n161 163.367
R705 B.n166 B.n165 163.367
R706 B.n170 B.n169 163.367
R707 B.n174 B.n173 163.367
R708 B.n178 B.n177 163.367
R709 B.n183 B.n182 163.367
R710 B.n187 B.n186 163.367
R711 B.n191 B.n190 163.367
R712 B.n195 B.n194 163.367
R713 B.n199 B.n198 163.367
R714 B.n204 B.n203 163.367
R715 B.n208 B.n207 163.367
R716 B.n212 B.n211 163.367
R717 B.n216 B.n215 163.367
R718 B.n220 B.n219 163.367
R719 B.n224 B.n223 163.367
R720 B.n228 B.n227 163.367
R721 B.n232 B.n231 163.367
R722 B.n236 B.n235 163.367
R723 B.n240 B.n239 163.367
R724 B.n244 B.n243 163.367
R725 B.n248 B.n247 163.367
R726 B.n252 B.n251 163.367
R727 B.n256 B.n255 163.367
R728 B.n258 B.n113 163.367
R729 B.n528 B.n339 163.367
R730 B.n528 B.n333 163.367
R731 B.n536 B.n333 163.367
R732 B.n536 B.n331 163.367
R733 B.n540 B.n331 163.367
R734 B.n540 B.n326 163.367
R735 B.n549 B.n326 163.367
R736 B.n549 B.n324 163.367
R737 B.n553 B.n324 163.367
R738 B.n553 B.n318 163.367
R739 B.n561 B.n318 163.367
R740 B.n561 B.n316 163.367
R741 B.n565 B.n316 163.367
R742 B.n565 B.n309 163.367
R743 B.n573 B.n309 163.367
R744 B.n573 B.n307 163.367
R745 B.n577 B.n307 163.367
R746 B.n577 B.n302 163.367
R747 B.n585 B.n302 163.367
R748 B.n585 B.n300 163.367
R749 B.n589 B.n300 163.367
R750 B.n589 B.n294 163.367
R751 B.n597 B.n294 163.367
R752 B.n597 B.n292 163.367
R753 B.n601 B.n292 163.367
R754 B.n601 B.n286 163.367
R755 B.n609 B.n286 163.367
R756 B.n609 B.n284 163.367
R757 B.n613 B.n284 163.367
R758 B.n613 B.n278 163.367
R759 B.n621 B.n278 163.367
R760 B.n621 B.n276 163.367
R761 B.n625 B.n276 163.367
R762 B.n625 B.n269 163.367
R763 B.n633 B.n269 163.367
R764 B.n633 B.n267 163.367
R765 B.n638 B.n267 163.367
R766 B.n638 B.n262 163.367
R767 B.n646 B.n262 163.367
R768 B.n647 B.n646 163.367
R769 B.n647 B.n5 163.367
R770 B.n6 B.n5 163.367
R771 B.n7 B.n6 163.367
R772 B.n653 B.n7 163.367
R773 B.n654 B.n653 163.367
R774 B.n654 B.n13 163.367
R775 B.n14 B.n13 163.367
R776 B.n15 B.n14 163.367
R777 B.n659 B.n15 163.367
R778 B.n659 B.n20 163.367
R779 B.n21 B.n20 163.367
R780 B.n22 B.n21 163.367
R781 B.n664 B.n22 163.367
R782 B.n664 B.n27 163.367
R783 B.n28 B.n27 163.367
R784 B.n29 B.n28 163.367
R785 B.n669 B.n29 163.367
R786 B.n669 B.n34 163.367
R787 B.n35 B.n34 163.367
R788 B.n36 B.n35 163.367
R789 B.n674 B.n36 163.367
R790 B.n674 B.n41 163.367
R791 B.n42 B.n41 163.367
R792 B.n43 B.n42 163.367
R793 B.n679 B.n43 163.367
R794 B.n679 B.n48 163.367
R795 B.n49 B.n48 163.367
R796 B.n50 B.n49 163.367
R797 B.n684 B.n50 163.367
R798 B.n684 B.n55 163.367
R799 B.n56 B.n55 163.367
R800 B.n57 B.n56 163.367
R801 B.n689 B.n57 163.367
R802 B.n689 B.n62 163.367
R803 B.n63 B.n62 163.367
R804 B.n64 B.n63 163.367
R805 B.n694 B.n64 163.367
R806 B.n694 B.n69 163.367
R807 B.n70 B.n69 163.367
R808 B.n71 B.n70 163.367
R809 B.n699 B.n71 163.367
R810 B.n699 B.n76 163.367
R811 B.n77 B.n76 163.367
R812 B.n377 B.n376 163.367
R813 B.n516 B.n376 163.367
R814 B.n514 B.n513 163.367
R815 B.n510 B.n509 163.367
R816 B.n506 B.n505 163.367
R817 B.n502 B.n501 163.367
R818 B.n498 B.n497 163.367
R819 B.n494 B.n493 163.367
R820 B.n490 B.n489 163.367
R821 B.n486 B.n485 163.367
R822 B.n482 B.n481 163.367
R823 B.n478 B.n477 163.367
R824 B.n474 B.n473 163.367
R825 B.n470 B.n469 163.367
R826 B.n466 B.n465 163.367
R827 B.n462 B.n461 163.367
R828 B.n458 B.n457 163.367
R829 B.n454 B.n453 163.367
R830 B.n450 B.n449 163.367
R831 B.n446 B.n445 163.367
R832 B.n442 B.n441 163.367
R833 B.n438 B.n437 163.367
R834 B.n434 B.n433 163.367
R835 B.n430 B.n429 163.367
R836 B.n426 B.n425 163.367
R837 B.n422 B.n421 163.367
R838 B.n418 B.n417 163.367
R839 B.n414 B.n413 163.367
R840 B.n410 B.n409 163.367
R841 B.n406 B.n405 163.367
R842 B.n402 B.n401 163.367
R843 B.n398 B.n397 163.367
R844 B.n394 B.n393 163.367
R845 B.n390 B.n389 163.367
R846 B.n386 B.n385 163.367
R847 B.n524 B.n341 163.367
R848 B.n530 B.n337 163.367
R849 B.n530 B.n335 163.367
R850 B.n534 B.n335 163.367
R851 B.n534 B.n329 163.367
R852 B.n543 B.n329 163.367
R853 B.n543 B.n327 163.367
R854 B.n547 B.n327 163.367
R855 B.n547 B.n322 163.367
R856 B.n555 B.n322 163.367
R857 B.n555 B.n320 163.367
R858 B.n559 B.n320 163.367
R859 B.n559 B.n314 163.367
R860 B.n567 B.n314 163.367
R861 B.n567 B.n312 163.367
R862 B.n571 B.n312 163.367
R863 B.n571 B.n306 163.367
R864 B.n579 B.n306 163.367
R865 B.n579 B.n304 163.367
R866 B.n583 B.n304 163.367
R867 B.n583 B.n298 163.367
R868 B.n591 B.n298 163.367
R869 B.n591 B.n296 163.367
R870 B.n595 B.n296 163.367
R871 B.n595 B.n290 163.367
R872 B.n603 B.n290 163.367
R873 B.n603 B.n288 163.367
R874 B.n607 B.n288 163.367
R875 B.n607 B.n282 163.367
R876 B.n615 B.n282 163.367
R877 B.n615 B.n280 163.367
R878 B.n619 B.n280 163.367
R879 B.n619 B.n274 163.367
R880 B.n627 B.n274 163.367
R881 B.n627 B.n272 163.367
R882 B.n631 B.n272 163.367
R883 B.n631 B.n266 163.367
R884 B.n640 B.n266 163.367
R885 B.n640 B.n264 163.367
R886 B.n644 B.n264 163.367
R887 B.n644 B.n3 163.367
R888 B.n790 B.n3 163.367
R889 B.n786 B.n2 163.367
R890 B.n786 B.n785 163.367
R891 B.n785 B.n9 163.367
R892 B.n781 B.n9 163.367
R893 B.n781 B.n11 163.367
R894 B.n777 B.n11 163.367
R895 B.n777 B.n17 163.367
R896 B.n773 B.n17 163.367
R897 B.n773 B.n19 163.367
R898 B.n769 B.n19 163.367
R899 B.n769 B.n24 163.367
R900 B.n765 B.n24 163.367
R901 B.n765 B.n26 163.367
R902 B.n761 B.n26 163.367
R903 B.n761 B.n31 163.367
R904 B.n757 B.n31 163.367
R905 B.n757 B.n33 163.367
R906 B.n753 B.n33 163.367
R907 B.n753 B.n38 163.367
R908 B.n749 B.n38 163.367
R909 B.n749 B.n40 163.367
R910 B.n745 B.n40 163.367
R911 B.n745 B.n45 163.367
R912 B.n741 B.n45 163.367
R913 B.n741 B.n47 163.367
R914 B.n737 B.n47 163.367
R915 B.n737 B.n52 163.367
R916 B.n733 B.n52 163.367
R917 B.n733 B.n54 163.367
R918 B.n729 B.n54 163.367
R919 B.n729 B.n59 163.367
R920 B.n725 B.n59 163.367
R921 B.n725 B.n61 163.367
R922 B.n721 B.n61 163.367
R923 B.n721 B.n65 163.367
R924 B.n717 B.n65 163.367
R925 B.n717 B.n67 163.367
R926 B.n713 B.n67 163.367
R927 B.n713 B.n73 163.367
R928 B.n709 B.n73 163.367
R929 B.n709 B.n75 163.367
R930 B.n114 B.t14 119.276
R931 B.n381 B.t21 119.276
R932 B.n116 B.t17 119.266
R933 B.n378 B.t11 119.266
R934 B.n523 B.n338 106.207
R935 B.n707 B.n706 106.207
R936 B.n115 B.t15 75.0582
R937 B.n382 B.t20 75.0582
R938 B.n117 B.t18 75.0485
R939 B.n379 B.t10 75.0485
R940 B.n118 B.n78 71.676
R941 B.n122 B.n79 71.676
R942 B.n126 B.n80 71.676
R943 B.n130 B.n81 71.676
R944 B.n134 B.n82 71.676
R945 B.n138 B.n83 71.676
R946 B.n142 B.n84 71.676
R947 B.n146 B.n85 71.676
R948 B.n150 B.n86 71.676
R949 B.n154 B.n87 71.676
R950 B.n158 B.n88 71.676
R951 B.n162 B.n89 71.676
R952 B.n166 B.n90 71.676
R953 B.n170 B.n91 71.676
R954 B.n174 B.n92 71.676
R955 B.n178 B.n93 71.676
R956 B.n183 B.n94 71.676
R957 B.n187 B.n95 71.676
R958 B.n191 B.n96 71.676
R959 B.n195 B.n97 71.676
R960 B.n199 B.n98 71.676
R961 B.n204 B.n99 71.676
R962 B.n208 B.n100 71.676
R963 B.n212 B.n101 71.676
R964 B.n216 B.n102 71.676
R965 B.n220 B.n103 71.676
R966 B.n224 B.n104 71.676
R967 B.n228 B.n105 71.676
R968 B.n232 B.n106 71.676
R969 B.n236 B.n107 71.676
R970 B.n240 B.n108 71.676
R971 B.n244 B.n109 71.676
R972 B.n248 B.n110 71.676
R973 B.n252 B.n111 71.676
R974 B.n256 B.n112 71.676
R975 B.n705 B.n113 71.676
R976 B.n705 B.n704 71.676
R977 B.n258 B.n112 71.676
R978 B.n255 B.n111 71.676
R979 B.n251 B.n110 71.676
R980 B.n247 B.n109 71.676
R981 B.n243 B.n108 71.676
R982 B.n239 B.n107 71.676
R983 B.n235 B.n106 71.676
R984 B.n231 B.n105 71.676
R985 B.n227 B.n104 71.676
R986 B.n223 B.n103 71.676
R987 B.n219 B.n102 71.676
R988 B.n215 B.n101 71.676
R989 B.n211 B.n100 71.676
R990 B.n207 B.n99 71.676
R991 B.n203 B.n98 71.676
R992 B.n198 B.n97 71.676
R993 B.n194 B.n96 71.676
R994 B.n190 B.n95 71.676
R995 B.n186 B.n94 71.676
R996 B.n182 B.n93 71.676
R997 B.n177 B.n92 71.676
R998 B.n173 B.n91 71.676
R999 B.n169 B.n90 71.676
R1000 B.n165 B.n89 71.676
R1001 B.n161 B.n88 71.676
R1002 B.n157 B.n87 71.676
R1003 B.n153 B.n86 71.676
R1004 B.n149 B.n85 71.676
R1005 B.n145 B.n84 71.676
R1006 B.n141 B.n83 71.676
R1007 B.n137 B.n82 71.676
R1008 B.n133 B.n81 71.676
R1009 B.n129 B.n80 71.676
R1010 B.n125 B.n79 71.676
R1011 B.n121 B.n78 71.676
R1012 B.n522 B.n521 71.676
R1013 B.n516 B.n342 71.676
R1014 B.n513 B.n343 71.676
R1015 B.n509 B.n344 71.676
R1016 B.n505 B.n345 71.676
R1017 B.n501 B.n346 71.676
R1018 B.n497 B.n347 71.676
R1019 B.n493 B.n348 71.676
R1020 B.n489 B.n349 71.676
R1021 B.n485 B.n350 71.676
R1022 B.n481 B.n351 71.676
R1023 B.n477 B.n352 71.676
R1024 B.n473 B.n353 71.676
R1025 B.n469 B.n354 71.676
R1026 B.n465 B.n355 71.676
R1027 B.n461 B.n356 71.676
R1028 B.n457 B.n357 71.676
R1029 B.n453 B.n358 71.676
R1030 B.n449 B.n359 71.676
R1031 B.n445 B.n360 71.676
R1032 B.n441 B.n361 71.676
R1033 B.n437 B.n362 71.676
R1034 B.n433 B.n363 71.676
R1035 B.n429 B.n364 71.676
R1036 B.n425 B.n365 71.676
R1037 B.n421 B.n366 71.676
R1038 B.n417 B.n367 71.676
R1039 B.n413 B.n368 71.676
R1040 B.n409 B.n369 71.676
R1041 B.n405 B.n370 71.676
R1042 B.n401 B.n371 71.676
R1043 B.n397 B.n372 71.676
R1044 B.n393 B.n373 71.676
R1045 B.n389 B.n374 71.676
R1046 B.n385 B.n375 71.676
R1047 B.n522 B.n377 71.676
R1048 B.n514 B.n342 71.676
R1049 B.n510 B.n343 71.676
R1050 B.n506 B.n344 71.676
R1051 B.n502 B.n345 71.676
R1052 B.n498 B.n346 71.676
R1053 B.n494 B.n347 71.676
R1054 B.n490 B.n348 71.676
R1055 B.n486 B.n349 71.676
R1056 B.n482 B.n350 71.676
R1057 B.n478 B.n351 71.676
R1058 B.n474 B.n352 71.676
R1059 B.n470 B.n353 71.676
R1060 B.n466 B.n354 71.676
R1061 B.n462 B.n355 71.676
R1062 B.n458 B.n356 71.676
R1063 B.n454 B.n357 71.676
R1064 B.n450 B.n358 71.676
R1065 B.n446 B.n359 71.676
R1066 B.n442 B.n360 71.676
R1067 B.n438 B.n361 71.676
R1068 B.n434 B.n362 71.676
R1069 B.n430 B.n363 71.676
R1070 B.n426 B.n364 71.676
R1071 B.n422 B.n365 71.676
R1072 B.n418 B.n366 71.676
R1073 B.n414 B.n367 71.676
R1074 B.n410 B.n368 71.676
R1075 B.n406 B.n369 71.676
R1076 B.n402 B.n370 71.676
R1077 B.n398 B.n371 71.676
R1078 B.n394 B.n372 71.676
R1079 B.n390 B.n373 71.676
R1080 B.n386 B.n374 71.676
R1081 B.n375 B.n341 71.676
R1082 B.n791 B.n790 71.676
R1083 B.n791 B.n2 71.676
R1084 B.n180 B.n117 59.5399
R1085 B.n201 B.n115 59.5399
R1086 B.n383 B.n382 59.5399
R1087 B.n380 B.n379 59.5399
R1088 B.n529 B.n338 54.3018
R1089 B.n529 B.n334 54.3018
R1090 B.n535 B.n334 54.3018
R1091 B.n535 B.n330 54.3018
R1092 B.n542 B.n330 54.3018
R1093 B.n542 B.n541 54.3018
R1094 B.n548 B.n323 54.3018
R1095 B.n554 B.n323 54.3018
R1096 B.n554 B.n319 54.3018
R1097 B.n560 B.n319 54.3018
R1098 B.n560 B.n315 54.3018
R1099 B.n566 B.n315 54.3018
R1100 B.n566 B.n310 54.3018
R1101 B.n572 B.n310 54.3018
R1102 B.n572 B.n311 54.3018
R1103 B.n578 B.n303 54.3018
R1104 B.n584 B.n303 54.3018
R1105 B.n584 B.n299 54.3018
R1106 B.n590 B.n299 54.3018
R1107 B.n590 B.n295 54.3018
R1108 B.n596 B.n295 54.3018
R1109 B.n602 B.n291 54.3018
R1110 B.n602 B.n287 54.3018
R1111 B.n608 B.n287 54.3018
R1112 B.n608 B.n283 54.3018
R1113 B.n614 B.n283 54.3018
R1114 B.n620 B.n279 54.3018
R1115 B.n620 B.n275 54.3018
R1116 B.n626 B.n275 54.3018
R1117 B.n626 B.n270 54.3018
R1118 B.n632 B.n270 54.3018
R1119 B.n632 B.n271 54.3018
R1120 B.n639 B.n263 54.3018
R1121 B.n645 B.n263 54.3018
R1122 B.n645 B.n4 54.3018
R1123 B.n789 B.n4 54.3018
R1124 B.n789 B.n788 54.3018
R1125 B.n788 B.n787 54.3018
R1126 B.n787 B.n8 54.3018
R1127 B.n12 B.n8 54.3018
R1128 B.n780 B.n12 54.3018
R1129 B.n779 B.n778 54.3018
R1130 B.n778 B.n16 54.3018
R1131 B.n772 B.n16 54.3018
R1132 B.n772 B.n771 54.3018
R1133 B.n771 B.n770 54.3018
R1134 B.n770 B.n23 54.3018
R1135 B.n764 B.n763 54.3018
R1136 B.n763 B.n762 54.3018
R1137 B.n762 B.n30 54.3018
R1138 B.n756 B.n30 54.3018
R1139 B.n756 B.n755 54.3018
R1140 B.n754 B.n37 54.3018
R1141 B.n748 B.n37 54.3018
R1142 B.n748 B.n747 54.3018
R1143 B.n747 B.n746 54.3018
R1144 B.n746 B.n44 54.3018
R1145 B.n740 B.n44 54.3018
R1146 B.n739 B.n738 54.3018
R1147 B.n738 B.n51 54.3018
R1148 B.n732 B.n51 54.3018
R1149 B.n732 B.n731 54.3018
R1150 B.n731 B.n730 54.3018
R1151 B.n730 B.n58 54.3018
R1152 B.n724 B.n58 54.3018
R1153 B.n724 B.n723 54.3018
R1154 B.n723 B.n722 54.3018
R1155 B.n716 B.n68 54.3018
R1156 B.n716 B.n715 54.3018
R1157 B.n715 B.n714 54.3018
R1158 B.n714 B.n72 54.3018
R1159 B.n708 B.n72 54.3018
R1160 B.n708 B.n707 54.3018
R1161 B.t4 B.n291 47.1148
R1162 B.n755 B.t0 47.1148
R1163 B.n614 B.t2 45.5177
R1164 B.n764 B.t3 45.5177
R1165 B.n117 B.n116 44.2187
R1166 B.n115 B.n114 44.2187
R1167 B.n382 B.n381 44.2187
R1168 B.n379 B.n378 44.2187
R1169 B.n520 B.n336 35.1225
R1170 B.n526 B.n525 35.1225
R1171 B.n703 B.n702 35.1225
R1172 B.n119 B.n74 35.1225
R1173 B.n578 B.t5 31.1439
R1174 B.n740 B.t6 31.1439
R1175 B.n271 B.t1 29.5468
R1176 B.t7 B.n779 29.5468
R1177 B.n541 B.t9 27.9497
R1178 B.n68 B.t13 27.9497
R1179 B.n548 B.t9 26.3526
R1180 B.n722 B.t13 26.3526
R1181 B.n639 B.t1 24.7555
R1182 B.n780 B.t7 24.7555
R1183 B.n311 B.t5 23.1584
R1184 B.t6 B.n739 23.1584
R1185 B B.n792 18.0485
R1186 B.n531 B.n336 10.6151
R1187 B.n532 B.n531 10.6151
R1188 B.n533 B.n532 10.6151
R1189 B.n533 B.n328 10.6151
R1190 B.n544 B.n328 10.6151
R1191 B.n545 B.n544 10.6151
R1192 B.n546 B.n545 10.6151
R1193 B.n546 B.n321 10.6151
R1194 B.n556 B.n321 10.6151
R1195 B.n557 B.n556 10.6151
R1196 B.n558 B.n557 10.6151
R1197 B.n558 B.n313 10.6151
R1198 B.n568 B.n313 10.6151
R1199 B.n569 B.n568 10.6151
R1200 B.n570 B.n569 10.6151
R1201 B.n570 B.n305 10.6151
R1202 B.n580 B.n305 10.6151
R1203 B.n581 B.n580 10.6151
R1204 B.n582 B.n581 10.6151
R1205 B.n582 B.n297 10.6151
R1206 B.n592 B.n297 10.6151
R1207 B.n593 B.n592 10.6151
R1208 B.n594 B.n593 10.6151
R1209 B.n594 B.n289 10.6151
R1210 B.n604 B.n289 10.6151
R1211 B.n605 B.n604 10.6151
R1212 B.n606 B.n605 10.6151
R1213 B.n606 B.n281 10.6151
R1214 B.n616 B.n281 10.6151
R1215 B.n617 B.n616 10.6151
R1216 B.n618 B.n617 10.6151
R1217 B.n618 B.n273 10.6151
R1218 B.n628 B.n273 10.6151
R1219 B.n629 B.n628 10.6151
R1220 B.n630 B.n629 10.6151
R1221 B.n630 B.n265 10.6151
R1222 B.n641 B.n265 10.6151
R1223 B.n642 B.n641 10.6151
R1224 B.n643 B.n642 10.6151
R1225 B.n643 B.n0 10.6151
R1226 B.n520 B.n519 10.6151
R1227 B.n519 B.n518 10.6151
R1228 B.n518 B.n517 10.6151
R1229 B.n517 B.n515 10.6151
R1230 B.n515 B.n512 10.6151
R1231 B.n512 B.n511 10.6151
R1232 B.n511 B.n508 10.6151
R1233 B.n508 B.n507 10.6151
R1234 B.n507 B.n504 10.6151
R1235 B.n504 B.n503 10.6151
R1236 B.n503 B.n500 10.6151
R1237 B.n500 B.n499 10.6151
R1238 B.n499 B.n496 10.6151
R1239 B.n496 B.n495 10.6151
R1240 B.n495 B.n492 10.6151
R1241 B.n492 B.n491 10.6151
R1242 B.n491 B.n488 10.6151
R1243 B.n488 B.n487 10.6151
R1244 B.n487 B.n484 10.6151
R1245 B.n484 B.n483 10.6151
R1246 B.n483 B.n480 10.6151
R1247 B.n480 B.n479 10.6151
R1248 B.n479 B.n476 10.6151
R1249 B.n476 B.n475 10.6151
R1250 B.n475 B.n472 10.6151
R1251 B.n472 B.n471 10.6151
R1252 B.n471 B.n468 10.6151
R1253 B.n468 B.n467 10.6151
R1254 B.n467 B.n464 10.6151
R1255 B.n464 B.n463 10.6151
R1256 B.n460 B.n459 10.6151
R1257 B.n459 B.n456 10.6151
R1258 B.n456 B.n455 10.6151
R1259 B.n455 B.n452 10.6151
R1260 B.n452 B.n451 10.6151
R1261 B.n451 B.n448 10.6151
R1262 B.n448 B.n447 10.6151
R1263 B.n447 B.n444 10.6151
R1264 B.n444 B.n443 10.6151
R1265 B.n440 B.n439 10.6151
R1266 B.n439 B.n436 10.6151
R1267 B.n436 B.n435 10.6151
R1268 B.n435 B.n432 10.6151
R1269 B.n432 B.n431 10.6151
R1270 B.n431 B.n428 10.6151
R1271 B.n428 B.n427 10.6151
R1272 B.n427 B.n424 10.6151
R1273 B.n424 B.n423 10.6151
R1274 B.n423 B.n420 10.6151
R1275 B.n420 B.n419 10.6151
R1276 B.n419 B.n416 10.6151
R1277 B.n416 B.n415 10.6151
R1278 B.n415 B.n412 10.6151
R1279 B.n412 B.n411 10.6151
R1280 B.n411 B.n408 10.6151
R1281 B.n408 B.n407 10.6151
R1282 B.n407 B.n404 10.6151
R1283 B.n404 B.n403 10.6151
R1284 B.n403 B.n400 10.6151
R1285 B.n400 B.n399 10.6151
R1286 B.n399 B.n396 10.6151
R1287 B.n396 B.n395 10.6151
R1288 B.n395 B.n392 10.6151
R1289 B.n392 B.n391 10.6151
R1290 B.n391 B.n388 10.6151
R1291 B.n388 B.n387 10.6151
R1292 B.n387 B.n384 10.6151
R1293 B.n384 B.n340 10.6151
R1294 B.n525 B.n340 10.6151
R1295 B.n527 B.n526 10.6151
R1296 B.n527 B.n332 10.6151
R1297 B.n537 B.n332 10.6151
R1298 B.n538 B.n537 10.6151
R1299 B.n539 B.n538 10.6151
R1300 B.n539 B.n325 10.6151
R1301 B.n550 B.n325 10.6151
R1302 B.n551 B.n550 10.6151
R1303 B.n552 B.n551 10.6151
R1304 B.n552 B.n317 10.6151
R1305 B.n562 B.n317 10.6151
R1306 B.n563 B.n562 10.6151
R1307 B.n564 B.n563 10.6151
R1308 B.n564 B.n308 10.6151
R1309 B.n574 B.n308 10.6151
R1310 B.n575 B.n574 10.6151
R1311 B.n576 B.n575 10.6151
R1312 B.n576 B.n301 10.6151
R1313 B.n586 B.n301 10.6151
R1314 B.n587 B.n586 10.6151
R1315 B.n588 B.n587 10.6151
R1316 B.n588 B.n293 10.6151
R1317 B.n598 B.n293 10.6151
R1318 B.n599 B.n598 10.6151
R1319 B.n600 B.n599 10.6151
R1320 B.n600 B.n285 10.6151
R1321 B.n610 B.n285 10.6151
R1322 B.n611 B.n610 10.6151
R1323 B.n612 B.n611 10.6151
R1324 B.n612 B.n277 10.6151
R1325 B.n622 B.n277 10.6151
R1326 B.n623 B.n622 10.6151
R1327 B.n624 B.n623 10.6151
R1328 B.n624 B.n268 10.6151
R1329 B.n634 B.n268 10.6151
R1330 B.n635 B.n634 10.6151
R1331 B.n637 B.n635 10.6151
R1332 B.n637 B.n636 10.6151
R1333 B.n636 B.n261 10.6151
R1334 B.n648 B.n261 10.6151
R1335 B.n649 B.n648 10.6151
R1336 B.n650 B.n649 10.6151
R1337 B.n651 B.n650 10.6151
R1338 B.n652 B.n651 10.6151
R1339 B.n655 B.n652 10.6151
R1340 B.n656 B.n655 10.6151
R1341 B.n657 B.n656 10.6151
R1342 B.n658 B.n657 10.6151
R1343 B.n660 B.n658 10.6151
R1344 B.n661 B.n660 10.6151
R1345 B.n662 B.n661 10.6151
R1346 B.n663 B.n662 10.6151
R1347 B.n665 B.n663 10.6151
R1348 B.n666 B.n665 10.6151
R1349 B.n667 B.n666 10.6151
R1350 B.n668 B.n667 10.6151
R1351 B.n670 B.n668 10.6151
R1352 B.n671 B.n670 10.6151
R1353 B.n672 B.n671 10.6151
R1354 B.n673 B.n672 10.6151
R1355 B.n675 B.n673 10.6151
R1356 B.n676 B.n675 10.6151
R1357 B.n677 B.n676 10.6151
R1358 B.n678 B.n677 10.6151
R1359 B.n680 B.n678 10.6151
R1360 B.n681 B.n680 10.6151
R1361 B.n682 B.n681 10.6151
R1362 B.n683 B.n682 10.6151
R1363 B.n685 B.n683 10.6151
R1364 B.n686 B.n685 10.6151
R1365 B.n687 B.n686 10.6151
R1366 B.n688 B.n687 10.6151
R1367 B.n690 B.n688 10.6151
R1368 B.n691 B.n690 10.6151
R1369 B.n692 B.n691 10.6151
R1370 B.n693 B.n692 10.6151
R1371 B.n695 B.n693 10.6151
R1372 B.n696 B.n695 10.6151
R1373 B.n697 B.n696 10.6151
R1374 B.n698 B.n697 10.6151
R1375 B.n700 B.n698 10.6151
R1376 B.n701 B.n700 10.6151
R1377 B.n702 B.n701 10.6151
R1378 B.n784 B.n1 10.6151
R1379 B.n784 B.n783 10.6151
R1380 B.n783 B.n782 10.6151
R1381 B.n782 B.n10 10.6151
R1382 B.n776 B.n10 10.6151
R1383 B.n776 B.n775 10.6151
R1384 B.n775 B.n774 10.6151
R1385 B.n774 B.n18 10.6151
R1386 B.n768 B.n18 10.6151
R1387 B.n768 B.n767 10.6151
R1388 B.n767 B.n766 10.6151
R1389 B.n766 B.n25 10.6151
R1390 B.n760 B.n25 10.6151
R1391 B.n760 B.n759 10.6151
R1392 B.n759 B.n758 10.6151
R1393 B.n758 B.n32 10.6151
R1394 B.n752 B.n32 10.6151
R1395 B.n752 B.n751 10.6151
R1396 B.n751 B.n750 10.6151
R1397 B.n750 B.n39 10.6151
R1398 B.n744 B.n39 10.6151
R1399 B.n744 B.n743 10.6151
R1400 B.n743 B.n742 10.6151
R1401 B.n742 B.n46 10.6151
R1402 B.n736 B.n46 10.6151
R1403 B.n736 B.n735 10.6151
R1404 B.n735 B.n734 10.6151
R1405 B.n734 B.n53 10.6151
R1406 B.n728 B.n53 10.6151
R1407 B.n728 B.n727 10.6151
R1408 B.n727 B.n726 10.6151
R1409 B.n726 B.n60 10.6151
R1410 B.n720 B.n60 10.6151
R1411 B.n720 B.n719 10.6151
R1412 B.n719 B.n718 10.6151
R1413 B.n718 B.n66 10.6151
R1414 B.n712 B.n66 10.6151
R1415 B.n712 B.n711 10.6151
R1416 B.n711 B.n710 10.6151
R1417 B.n710 B.n74 10.6151
R1418 B.n120 B.n119 10.6151
R1419 B.n123 B.n120 10.6151
R1420 B.n124 B.n123 10.6151
R1421 B.n127 B.n124 10.6151
R1422 B.n128 B.n127 10.6151
R1423 B.n131 B.n128 10.6151
R1424 B.n132 B.n131 10.6151
R1425 B.n135 B.n132 10.6151
R1426 B.n136 B.n135 10.6151
R1427 B.n139 B.n136 10.6151
R1428 B.n140 B.n139 10.6151
R1429 B.n143 B.n140 10.6151
R1430 B.n144 B.n143 10.6151
R1431 B.n147 B.n144 10.6151
R1432 B.n148 B.n147 10.6151
R1433 B.n151 B.n148 10.6151
R1434 B.n152 B.n151 10.6151
R1435 B.n155 B.n152 10.6151
R1436 B.n156 B.n155 10.6151
R1437 B.n159 B.n156 10.6151
R1438 B.n160 B.n159 10.6151
R1439 B.n163 B.n160 10.6151
R1440 B.n164 B.n163 10.6151
R1441 B.n167 B.n164 10.6151
R1442 B.n168 B.n167 10.6151
R1443 B.n171 B.n168 10.6151
R1444 B.n172 B.n171 10.6151
R1445 B.n175 B.n172 10.6151
R1446 B.n176 B.n175 10.6151
R1447 B.n179 B.n176 10.6151
R1448 B.n184 B.n181 10.6151
R1449 B.n185 B.n184 10.6151
R1450 B.n188 B.n185 10.6151
R1451 B.n189 B.n188 10.6151
R1452 B.n192 B.n189 10.6151
R1453 B.n193 B.n192 10.6151
R1454 B.n196 B.n193 10.6151
R1455 B.n197 B.n196 10.6151
R1456 B.n200 B.n197 10.6151
R1457 B.n205 B.n202 10.6151
R1458 B.n206 B.n205 10.6151
R1459 B.n209 B.n206 10.6151
R1460 B.n210 B.n209 10.6151
R1461 B.n213 B.n210 10.6151
R1462 B.n214 B.n213 10.6151
R1463 B.n217 B.n214 10.6151
R1464 B.n218 B.n217 10.6151
R1465 B.n221 B.n218 10.6151
R1466 B.n222 B.n221 10.6151
R1467 B.n225 B.n222 10.6151
R1468 B.n226 B.n225 10.6151
R1469 B.n229 B.n226 10.6151
R1470 B.n230 B.n229 10.6151
R1471 B.n233 B.n230 10.6151
R1472 B.n234 B.n233 10.6151
R1473 B.n237 B.n234 10.6151
R1474 B.n238 B.n237 10.6151
R1475 B.n241 B.n238 10.6151
R1476 B.n242 B.n241 10.6151
R1477 B.n245 B.n242 10.6151
R1478 B.n246 B.n245 10.6151
R1479 B.n249 B.n246 10.6151
R1480 B.n250 B.n249 10.6151
R1481 B.n253 B.n250 10.6151
R1482 B.n254 B.n253 10.6151
R1483 B.n257 B.n254 10.6151
R1484 B.n259 B.n257 10.6151
R1485 B.n260 B.n259 10.6151
R1486 B.n703 B.n260 10.6151
R1487 B.n463 B.n380 9.36635
R1488 B.n440 B.n383 9.36635
R1489 B.n180 B.n179 9.36635
R1490 B.n202 B.n201 9.36635
R1491 B.t2 B.n279 8.78453
R1492 B.t3 B.n23 8.78453
R1493 B.n792 B.n0 8.11757
R1494 B.n792 B.n1 8.11757
R1495 B.n596 B.t4 7.18743
R1496 B.t0 B.n754 7.18743
R1497 B.n460 B.n380 1.24928
R1498 B.n443 B.n383 1.24928
R1499 B.n181 B.n180 1.24928
R1500 B.n201 B.n200 1.24928
R1501 VN.n43 VN.n23 161.3
R1502 VN.n42 VN.n41 161.3
R1503 VN.n40 VN.n24 161.3
R1504 VN.n39 VN.n38 161.3
R1505 VN.n36 VN.n25 161.3
R1506 VN.n35 VN.n34 161.3
R1507 VN.n33 VN.n26 161.3
R1508 VN.n32 VN.n31 161.3
R1509 VN.n30 VN.n27 161.3
R1510 VN.n20 VN.n0 161.3
R1511 VN.n19 VN.n18 161.3
R1512 VN.n17 VN.n1 161.3
R1513 VN.n16 VN.n15 161.3
R1514 VN.n13 VN.n2 161.3
R1515 VN.n12 VN.n11 161.3
R1516 VN.n10 VN.n3 161.3
R1517 VN.n9 VN.n8 161.3
R1518 VN.n7 VN.n4 161.3
R1519 VN.n5 VN.t2 135.59
R1520 VN.n28 VN.t5 135.59
R1521 VN.n6 VN.t6 105.052
R1522 VN.n14 VN.t4 105.052
R1523 VN.n21 VN.t1 105.052
R1524 VN.n29 VN.t3 105.052
R1525 VN.n37 VN.t0 105.052
R1526 VN.n44 VN.t7 105.052
R1527 VN.n22 VN.n21 90.2511
R1528 VN.n45 VN.n44 90.2511
R1529 VN.n6 VN.n5 63.2137
R1530 VN.n29 VN.n28 63.2137
R1531 VN.n19 VN.n1 56.5617
R1532 VN.n42 VN.n24 56.5617
R1533 VN VN.n45 45.5058
R1534 VN.n8 VN.n3 40.577
R1535 VN.n12 VN.n3 40.577
R1536 VN.n31 VN.n26 40.577
R1537 VN.n35 VN.n26 40.577
R1538 VN.n8 VN.n7 24.5923
R1539 VN.n13 VN.n12 24.5923
R1540 VN.n15 VN.n1 24.5923
R1541 VN.n20 VN.n19 24.5923
R1542 VN.n31 VN.n30 24.5923
R1543 VN.n38 VN.n24 24.5923
R1544 VN.n36 VN.n35 24.5923
R1545 VN.n43 VN.n42 24.5923
R1546 VN.n21 VN.n20 20.6576
R1547 VN.n44 VN.n43 20.6576
R1548 VN.n15 VN.n14 17.7066
R1549 VN.n38 VN.n37 17.7066
R1550 VN.n28 VN.n27 13.203
R1551 VN.n5 VN.n4 13.203
R1552 VN.n7 VN.n6 6.88621
R1553 VN.n14 VN.n13 6.88621
R1554 VN.n30 VN.n29 6.88621
R1555 VN.n37 VN.n36 6.88621
R1556 VN.n45 VN.n23 0.278335
R1557 VN.n22 VN.n0 0.278335
R1558 VN.n41 VN.n23 0.189894
R1559 VN.n41 VN.n40 0.189894
R1560 VN.n40 VN.n39 0.189894
R1561 VN.n39 VN.n25 0.189894
R1562 VN.n34 VN.n25 0.189894
R1563 VN.n34 VN.n33 0.189894
R1564 VN.n33 VN.n32 0.189894
R1565 VN.n32 VN.n27 0.189894
R1566 VN.n9 VN.n4 0.189894
R1567 VN.n10 VN.n9 0.189894
R1568 VN.n11 VN.n10 0.189894
R1569 VN.n11 VN.n2 0.189894
R1570 VN.n16 VN.n2 0.189894
R1571 VN.n17 VN.n16 0.189894
R1572 VN.n18 VN.n17 0.189894
R1573 VN.n18 VN.n0 0.189894
R1574 VN VN.n22 0.153485
R1575 VDD2.n2 VDD2.n1 64.7456
R1576 VDD2.n2 VDD2.n0 64.7456
R1577 VDD2 VDD2.n5 64.7428
R1578 VDD2.n4 VDD2.n3 63.8182
R1579 VDD2.n4 VDD2.n2 39.8877
R1580 VDD2.n5 VDD2.t4 2.32991
R1581 VDD2.n5 VDD2.t2 2.32991
R1582 VDD2.n3 VDD2.t0 2.32991
R1583 VDD2.n3 VDD2.t7 2.32991
R1584 VDD2.n1 VDD2.t3 2.32991
R1585 VDD2.n1 VDD2.t6 2.32991
R1586 VDD2.n0 VDD2.t5 2.32991
R1587 VDD2.n0 VDD2.t1 2.32991
R1588 VDD2 VDD2.n4 1.04145
C0 VN VDD1 0.150969f
C1 VN VP 6.21651f
C2 VN VDD2 5.89327f
C3 VTAIL VDD1 6.73786f
C4 VP VTAIL 6.25027f
C5 VTAIL VDD2 6.78792f
C6 VN VTAIL 6.23616f
C7 VP VDD1 6.19216f
C8 VDD1 VDD2 1.43976f
C9 VP VDD2 0.45092f
C10 VDD2 B 4.45974f
C11 VDD1 B 4.826319f
C12 VTAIL B 7.948561f
C13 VN B 12.74309f
C14 VP B 11.308582f
C15 VDD2.t5 B 0.165001f
C16 VDD2.t1 B 0.165001f
C17 VDD2.n0 B 1.43318f
C18 VDD2.t3 B 0.165001f
C19 VDD2.t6 B 0.165001f
C20 VDD2.n1 B 1.43318f
C21 VDD2.n2 B 2.64562f
C22 VDD2.t0 B 0.165001f
C23 VDD2.t7 B 0.165001f
C24 VDD2.n3 B 1.42681f
C25 VDD2.n4 B 2.41446f
C26 VDD2.t4 B 0.165001f
C27 VDD2.t2 B 0.165001f
C28 VDD2.n5 B 1.43315f
C29 VN.n0 B 0.0361f
C30 VN.t1 B 1.22211f
C31 VN.n1 B 0.042079f
C32 VN.n2 B 0.027384f
C33 VN.t4 B 1.22211f
C34 VN.n3 B 0.022117f
C35 VN.n4 B 0.203769f
C36 VN.t6 B 1.22211f
C37 VN.t2 B 1.35278f
C38 VN.n5 B 0.517663f
C39 VN.n6 B 0.507801f
C40 VN.n7 B 0.032731f
C41 VN.n8 B 0.054138f
C42 VN.n9 B 0.027384f
C43 VN.n10 B 0.027384f
C44 VN.n11 B 0.027384f
C45 VN.n12 B 0.054138f
C46 VN.n13 B 0.032731f
C47 VN.n14 B 0.449067f
C48 VN.n15 B 0.043761f
C49 VN.n16 B 0.027384f
C50 VN.n17 B 0.027384f
C51 VN.n18 B 0.027384f
C52 VN.n19 B 0.037533f
C53 VN.n20 B 0.046769f
C54 VN.n21 B 0.531702f
C55 VN.n22 B 0.032415f
C56 VN.n23 B 0.0361f
C57 VN.t7 B 1.22211f
C58 VN.n24 B 0.042079f
C59 VN.n25 B 0.027384f
C60 VN.t0 B 1.22211f
C61 VN.n26 B 0.022117f
C62 VN.n27 B 0.203769f
C63 VN.t3 B 1.22211f
C64 VN.t5 B 1.35278f
C65 VN.n28 B 0.517663f
C66 VN.n29 B 0.507801f
C67 VN.n30 B 0.032731f
C68 VN.n31 B 0.054138f
C69 VN.n32 B 0.027384f
C70 VN.n33 B 0.027384f
C71 VN.n34 B 0.027384f
C72 VN.n35 B 0.054138f
C73 VN.n36 B 0.032731f
C74 VN.n37 B 0.449067f
C75 VN.n38 B 0.043761f
C76 VN.n39 B 0.027384f
C77 VN.n40 B 0.027384f
C78 VN.n41 B 0.027384f
C79 VN.n42 B 0.037533f
C80 VN.n43 B 0.046769f
C81 VN.n44 B 0.531702f
C82 VN.n45 B 1.3119f
C83 VDD1.t3 B 0.16641f
C84 VDD1.t6 B 0.16641f
C85 VDD1.n0 B 1.44634f
C86 VDD1.t1 B 0.16641f
C87 VDD1.t5 B 0.16641f
C88 VDD1.n1 B 1.44543f
C89 VDD1.t2 B 0.16641f
C90 VDD1.t7 B 0.16641f
C91 VDD1.n2 B 1.44543f
C92 VDD1.n3 B 2.72034f
C93 VDD1.t0 B 0.16641f
C94 VDD1.t4 B 0.16641f
C95 VDD1.n4 B 1.439f
C96 VDD1.n5 B 2.46518f
C97 VTAIL.t3 B 0.138278f
C98 VTAIL.t0 B 0.138278f
C99 VTAIL.n0 B 1.13612f
C100 VTAIL.n1 B 0.33826f
C101 VTAIL.t7 B 1.44849f
C102 VTAIL.n2 B 0.430316f
C103 VTAIL.t11 B 1.44849f
C104 VTAIL.n3 B 0.430316f
C105 VTAIL.t9 B 0.138278f
C106 VTAIL.t14 B 0.138278f
C107 VTAIL.n4 B 1.13612f
C108 VTAIL.n5 B 0.464781f
C109 VTAIL.t15 B 1.44849f
C110 VTAIL.n6 B 1.29524f
C111 VTAIL.t5 B 1.4485f
C112 VTAIL.n7 B 1.29524f
C113 VTAIL.t4 B 0.138278f
C114 VTAIL.t2 B 0.138278f
C115 VTAIL.n8 B 1.13612f
C116 VTAIL.n9 B 0.464779f
C117 VTAIL.t1 B 1.4485f
C118 VTAIL.n10 B 0.43031f
C119 VTAIL.t12 B 1.4485f
C120 VTAIL.n11 B 0.43031f
C121 VTAIL.t13 B 0.138278f
C122 VTAIL.t8 B 0.138278f
C123 VTAIL.n12 B 1.13612f
C124 VTAIL.n13 B 0.464779f
C125 VTAIL.t10 B 1.4485f
C126 VTAIL.n14 B 1.29523f
C127 VTAIL.t6 B 1.44849f
C128 VTAIL.n15 B 1.29138f
C129 VP.n0 B 0.036967f
C130 VP.t0 B 1.25146f
C131 VP.n1 B 0.04309f
C132 VP.n2 B 0.028041f
C133 VP.t5 B 1.25146f
C134 VP.n3 B 0.022648f
C135 VP.n4 B 0.028041f
C136 VP.t2 B 1.25146f
C137 VP.n5 B 0.04309f
C138 VP.n6 B 0.036967f
C139 VP.t6 B 1.25146f
C140 VP.n7 B 0.036967f
C141 VP.t3 B 1.25146f
C142 VP.n8 B 0.04309f
C143 VP.n9 B 0.028041f
C144 VP.t7 B 1.25146f
C145 VP.n10 B 0.022648f
C146 VP.n11 B 0.208662f
C147 VP.t1 B 1.25146f
C148 VP.t4 B 1.38526f
C149 VP.n12 B 0.530093f
C150 VP.n13 B 0.519995f
C151 VP.n14 B 0.033517f
C152 VP.n15 B 0.055438f
C153 VP.n16 B 0.028041f
C154 VP.n17 B 0.028041f
C155 VP.n18 B 0.028041f
C156 VP.n19 B 0.055438f
C157 VP.n20 B 0.033517f
C158 VP.n21 B 0.45985f
C159 VP.n22 B 0.044812f
C160 VP.n23 B 0.028041f
C161 VP.n24 B 0.028041f
C162 VP.n25 B 0.028041f
C163 VP.n26 B 0.038435f
C164 VP.n27 B 0.047892f
C165 VP.n28 B 0.544469f
C166 VP.n29 B 1.32808f
C167 VP.n30 B 1.35043f
C168 VP.n31 B 0.544469f
C169 VP.n32 B 0.047892f
C170 VP.n33 B 0.038435f
C171 VP.n34 B 0.028041f
C172 VP.n35 B 0.028041f
C173 VP.n36 B 0.028041f
C174 VP.n37 B 0.044812f
C175 VP.n38 B 0.45985f
C176 VP.n39 B 0.033517f
C177 VP.n40 B 0.055438f
C178 VP.n41 B 0.028041f
C179 VP.n42 B 0.028041f
C180 VP.n43 B 0.028041f
C181 VP.n44 B 0.055438f
C182 VP.n45 B 0.033517f
C183 VP.n46 B 0.45985f
C184 VP.n47 B 0.044812f
C185 VP.n48 B 0.028041f
C186 VP.n49 B 0.028041f
C187 VP.n50 B 0.028041f
C188 VP.n51 B 0.038435f
C189 VP.n52 B 0.047892f
C190 VP.n53 B 0.544469f
C191 VP.n54 B 0.033194f
.ends

