* NGSPICE file created from diff_pair_sample_0016.ext - technology: sky130A

.subckt diff_pair_sample_0016 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VN.t0 VDD2.t1 w_n4260_n3952# sky130_fd_pr__pfet_01v8 ad=2.4618 pd=15.25 as=2.4618 ps=15.25 w=14.92 l=2.96
X1 VTAIL.t4 VP.t0 VDD1.t7 w_n4260_n3952# sky130_fd_pr__pfet_01v8 ad=2.4618 pd=15.25 as=2.4618 ps=15.25 w=14.92 l=2.96
X2 B.t11 B.t9 B.t10 w_n4260_n3952# sky130_fd_pr__pfet_01v8 ad=5.8188 pd=30.62 as=0 ps=0 w=14.92 l=2.96
X3 VDD2.t0 VN.t1 VTAIL.t14 w_n4260_n3952# sky130_fd_pr__pfet_01v8 ad=2.4618 pd=15.25 as=5.8188 ps=30.62 w=14.92 l=2.96
X4 VDD2.t3 VN.t2 VTAIL.t13 w_n4260_n3952# sky130_fd_pr__pfet_01v8 ad=2.4618 pd=15.25 as=2.4618 ps=15.25 w=14.92 l=2.96
X5 VTAIL.t5 VP.t1 VDD1.t6 w_n4260_n3952# sky130_fd_pr__pfet_01v8 ad=5.8188 pd=30.62 as=2.4618 ps=15.25 w=14.92 l=2.96
X6 VDD1.t5 VP.t2 VTAIL.t0 w_n4260_n3952# sky130_fd_pr__pfet_01v8 ad=2.4618 pd=15.25 as=5.8188 ps=30.62 w=14.92 l=2.96
X7 VTAIL.t12 VN.t3 VDD2.t2 w_n4260_n3952# sky130_fd_pr__pfet_01v8 ad=2.4618 pd=15.25 as=2.4618 ps=15.25 w=14.92 l=2.96
X8 VDD1.t4 VP.t3 VTAIL.t7 w_n4260_n3952# sky130_fd_pr__pfet_01v8 ad=2.4618 pd=15.25 as=5.8188 ps=30.62 w=14.92 l=2.96
X9 VDD1.t3 VP.t4 VTAIL.t1 w_n4260_n3952# sky130_fd_pr__pfet_01v8 ad=2.4618 pd=15.25 as=2.4618 ps=15.25 w=14.92 l=2.96
X10 VDD2.t5 VN.t4 VTAIL.t11 w_n4260_n3952# sky130_fd_pr__pfet_01v8 ad=2.4618 pd=15.25 as=5.8188 ps=30.62 w=14.92 l=2.96
X11 VDD2.t4 VN.t5 VTAIL.t10 w_n4260_n3952# sky130_fd_pr__pfet_01v8 ad=2.4618 pd=15.25 as=2.4618 ps=15.25 w=14.92 l=2.96
X12 B.t8 B.t6 B.t7 w_n4260_n3952# sky130_fd_pr__pfet_01v8 ad=5.8188 pd=30.62 as=0 ps=0 w=14.92 l=2.96
X13 VTAIL.t9 VN.t6 VDD2.t7 w_n4260_n3952# sky130_fd_pr__pfet_01v8 ad=5.8188 pd=30.62 as=2.4618 ps=15.25 w=14.92 l=2.96
X14 VTAIL.t3 VP.t5 VDD1.t2 w_n4260_n3952# sky130_fd_pr__pfet_01v8 ad=5.8188 pd=30.62 as=2.4618 ps=15.25 w=14.92 l=2.96
X15 B.t5 B.t3 B.t4 w_n4260_n3952# sky130_fd_pr__pfet_01v8 ad=5.8188 pd=30.62 as=0 ps=0 w=14.92 l=2.96
X16 VTAIL.t2 VP.t6 VDD1.t1 w_n4260_n3952# sky130_fd_pr__pfet_01v8 ad=2.4618 pd=15.25 as=2.4618 ps=15.25 w=14.92 l=2.96
X17 VDD1.t0 VP.t7 VTAIL.t6 w_n4260_n3952# sky130_fd_pr__pfet_01v8 ad=2.4618 pd=15.25 as=2.4618 ps=15.25 w=14.92 l=2.96
X18 VTAIL.t8 VN.t7 VDD2.t6 w_n4260_n3952# sky130_fd_pr__pfet_01v8 ad=5.8188 pd=30.62 as=2.4618 ps=15.25 w=14.92 l=2.96
X19 B.t2 B.t0 B.t1 w_n4260_n3952# sky130_fd_pr__pfet_01v8 ad=5.8188 pd=30.62 as=0 ps=0 w=14.92 l=2.96
R0 VN.n60 VN.n59 161.3
R1 VN.n58 VN.n32 161.3
R2 VN.n57 VN.n56 161.3
R3 VN.n55 VN.n33 161.3
R4 VN.n54 VN.n53 161.3
R5 VN.n52 VN.n34 161.3
R6 VN.n50 VN.n49 161.3
R7 VN.n48 VN.n35 161.3
R8 VN.n47 VN.n46 161.3
R9 VN.n45 VN.n36 161.3
R10 VN.n44 VN.n43 161.3
R11 VN.n42 VN.n37 161.3
R12 VN.n41 VN.n40 161.3
R13 VN.n29 VN.n28 161.3
R14 VN.n27 VN.n1 161.3
R15 VN.n26 VN.n25 161.3
R16 VN.n24 VN.n2 161.3
R17 VN.n23 VN.n22 161.3
R18 VN.n21 VN.n3 161.3
R19 VN.n19 VN.n18 161.3
R20 VN.n17 VN.n4 161.3
R21 VN.n16 VN.n15 161.3
R22 VN.n14 VN.n5 161.3
R23 VN.n13 VN.n12 161.3
R24 VN.n11 VN.n6 161.3
R25 VN.n10 VN.n9 161.3
R26 VN.n38 VN.t4 153.299
R27 VN.n7 VN.t6 153.299
R28 VN.n8 VN.t2 121.478
R29 VN.n20 VN.t3 121.478
R30 VN.n0 VN.t1 121.478
R31 VN.n39 VN.t0 121.478
R32 VN.n51 VN.t5 121.478
R33 VN.n31 VN.t7 121.478
R34 VN.n30 VN.n0 68.8507
R35 VN.n61 VN.n31 68.8507
R36 VN.n8 VN.n7 66.845
R37 VN.n39 VN.n38 66.845
R38 VN.n26 VN.n2 56.5617
R39 VN.n57 VN.n33 56.5617
R40 VN VN.n61 55.089
R41 VN.n14 VN.n13 40.577
R42 VN.n15 VN.n14 40.577
R43 VN.n45 VN.n44 40.577
R44 VN.n46 VN.n45 40.577
R45 VN.n9 VN.n6 24.5923
R46 VN.n13 VN.n6 24.5923
R47 VN.n15 VN.n4 24.5923
R48 VN.n19 VN.n4 24.5923
R49 VN.n22 VN.n21 24.5923
R50 VN.n22 VN.n2 24.5923
R51 VN.n27 VN.n26 24.5923
R52 VN.n28 VN.n27 24.5923
R53 VN.n44 VN.n37 24.5923
R54 VN.n40 VN.n37 24.5923
R55 VN.n53 VN.n33 24.5923
R56 VN.n53 VN.n52 24.5923
R57 VN.n50 VN.n35 24.5923
R58 VN.n46 VN.n35 24.5923
R59 VN.n59 VN.n58 24.5923
R60 VN.n58 VN.n57 24.5923
R61 VN.n28 VN.n0 21.3954
R62 VN.n59 VN.n31 21.3954
R63 VN.n21 VN.n20 17.4607
R64 VN.n52 VN.n51 17.4607
R65 VN.n9 VN.n8 7.13213
R66 VN.n20 VN.n19 7.13213
R67 VN.n40 VN.n39 7.13213
R68 VN.n51 VN.n50 7.13213
R69 VN.n41 VN.n38 5.44405
R70 VN.n10 VN.n7 5.44405
R71 VN.n61 VN.n60 0.354861
R72 VN.n30 VN.n29 0.354861
R73 VN VN.n30 0.267071
R74 VN.n60 VN.n32 0.189894
R75 VN.n56 VN.n32 0.189894
R76 VN.n56 VN.n55 0.189894
R77 VN.n55 VN.n54 0.189894
R78 VN.n54 VN.n34 0.189894
R79 VN.n49 VN.n34 0.189894
R80 VN.n49 VN.n48 0.189894
R81 VN.n48 VN.n47 0.189894
R82 VN.n47 VN.n36 0.189894
R83 VN.n43 VN.n36 0.189894
R84 VN.n43 VN.n42 0.189894
R85 VN.n42 VN.n41 0.189894
R86 VN.n11 VN.n10 0.189894
R87 VN.n12 VN.n11 0.189894
R88 VN.n12 VN.n5 0.189894
R89 VN.n16 VN.n5 0.189894
R90 VN.n17 VN.n16 0.189894
R91 VN.n18 VN.n17 0.189894
R92 VN.n18 VN.n3 0.189894
R93 VN.n23 VN.n3 0.189894
R94 VN.n24 VN.n23 0.189894
R95 VN.n25 VN.n24 0.189894
R96 VN.n25 VN.n1 0.189894
R97 VN.n29 VN.n1 0.189894
R98 VDD2.n2 VDD2.n1 70.8667
R99 VDD2.n2 VDD2.n0 70.8667
R100 VDD2 VDD2.n5 70.864
R101 VDD2.n4 VDD2.n3 69.5041
R102 VDD2.n4 VDD2.n2 49.3403
R103 VDD2.n5 VDD2.t1 2.17912
R104 VDD2.n5 VDD2.t5 2.17912
R105 VDD2.n3 VDD2.t6 2.17912
R106 VDD2.n3 VDD2.t4 2.17912
R107 VDD2.n1 VDD2.t2 2.17912
R108 VDD2.n1 VDD2.t0 2.17912
R109 VDD2.n0 VDD2.t7 2.17912
R110 VDD2.n0 VDD2.t3 2.17912
R111 VDD2 VDD2.n4 1.47679
R112 VTAIL.n658 VTAIL.n582 756.745
R113 VTAIL.n78 VTAIL.n2 756.745
R114 VTAIL.n160 VTAIL.n84 756.745
R115 VTAIL.n244 VTAIL.n168 756.745
R116 VTAIL.n576 VTAIL.n500 756.745
R117 VTAIL.n492 VTAIL.n416 756.745
R118 VTAIL.n410 VTAIL.n334 756.745
R119 VTAIL.n326 VTAIL.n250 756.745
R120 VTAIL.n609 VTAIL.n608 585
R121 VTAIL.n606 VTAIL.n605 585
R122 VTAIL.n615 VTAIL.n614 585
R123 VTAIL.n617 VTAIL.n616 585
R124 VTAIL.n602 VTAIL.n601 585
R125 VTAIL.n623 VTAIL.n622 585
R126 VTAIL.n626 VTAIL.n625 585
R127 VTAIL.n624 VTAIL.n598 585
R128 VTAIL.n631 VTAIL.n597 585
R129 VTAIL.n633 VTAIL.n632 585
R130 VTAIL.n635 VTAIL.n634 585
R131 VTAIL.n594 VTAIL.n593 585
R132 VTAIL.n641 VTAIL.n640 585
R133 VTAIL.n643 VTAIL.n642 585
R134 VTAIL.n590 VTAIL.n589 585
R135 VTAIL.n649 VTAIL.n648 585
R136 VTAIL.n651 VTAIL.n650 585
R137 VTAIL.n586 VTAIL.n585 585
R138 VTAIL.n657 VTAIL.n656 585
R139 VTAIL.n659 VTAIL.n658 585
R140 VTAIL.n29 VTAIL.n28 585
R141 VTAIL.n26 VTAIL.n25 585
R142 VTAIL.n35 VTAIL.n34 585
R143 VTAIL.n37 VTAIL.n36 585
R144 VTAIL.n22 VTAIL.n21 585
R145 VTAIL.n43 VTAIL.n42 585
R146 VTAIL.n46 VTAIL.n45 585
R147 VTAIL.n44 VTAIL.n18 585
R148 VTAIL.n51 VTAIL.n17 585
R149 VTAIL.n53 VTAIL.n52 585
R150 VTAIL.n55 VTAIL.n54 585
R151 VTAIL.n14 VTAIL.n13 585
R152 VTAIL.n61 VTAIL.n60 585
R153 VTAIL.n63 VTAIL.n62 585
R154 VTAIL.n10 VTAIL.n9 585
R155 VTAIL.n69 VTAIL.n68 585
R156 VTAIL.n71 VTAIL.n70 585
R157 VTAIL.n6 VTAIL.n5 585
R158 VTAIL.n77 VTAIL.n76 585
R159 VTAIL.n79 VTAIL.n78 585
R160 VTAIL.n111 VTAIL.n110 585
R161 VTAIL.n108 VTAIL.n107 585
R162 VTAIL.n117 VTAIL.n116 585
R163 VTAIL.n119 VTAIL.n118 585
R164 VTAIL.n104 VTAIL.n103 585
R165 VTAIL.n125 VTAIL.n124 585
R166 VTAIL.n128 VTAIL.n127 585
R167 VTAIL.n126 VTAIL.n100 585
R168 VTAIL.n133 VTAIL.n99 585
R169 VTAIL.n135 VTAIL.n134 585
R170 VTAIL.n137 VTAIL.n136 585
R171 VTAIL.n96 VTAIL.n95 585
R172 VTAIL.n143 VTAIL.n142 585
R173 VTAIL.n145 VTAIL.n144 585
R174 VTAIL.n92 VTAIL.n91 585
R175 VTAIL.n151 VTAIL.n150 585
R176 VTAIL.n153 VTAIL.n152 585
R177 VTAIL.n88 VTAIL.n87 585
R178 VTAIL.n159 VTAIL.n158 585
R179 VTAIL.n161 VTAIL.n160 585
R180 VTAIL.n195 VTAIL.n194 585
R181 VTAIL.n192 VTAIL.n191 585
R182 VTAIL.n201 VTAIL.n200 585
R183 VTAIL.n203 VTAIL.n202 585
R184 VTAIL.n188 VTAIL.n187 585
R185 VTAIL.n209 VTAIL.n208 585
R186 VTAIL.n212 VTAIL.n211 585
R187 VTAIL.n210 VTAIL.n184 585
R188 VTAIL.n217 VTAIL.n183 585
R189 VTAIL.n219 VTAIL.n218 585
R190 VTAIL.n221 VTAIL.n220 585
R191 VTAIL.n180 VTAIL.n179 585
R192 VTAIL.n227 VTAIL.n226 585
R193 VTAIL.n229 VTAIL.n228 585
R194 VTAIL.n176 VTAIL.n175 585
R195 VTAIL.n235 VTAIL.n234 585
R196 VTAIL.n237 VTAIL.n236 585
R197 VTAIL.n172 VTAIL.n171 585
R198 VTAIL.n243 VTAIL.n242 585
R199 VTAIL.n245 VTAIL.n244 585
R200 VTAIL.n577 VTAIL.n576 585
R201 VTAIL.n575 VTAIL.n574 585
R202 VTAIL.n504 VTAIL.n503 585
R203 VTAIL.n569 VTAIL.n568 585
R204 VTAIL.n567 VTAIL.n566 585
R205 VTAIL.n508 VTAIL.n507 585
R206 VTAIL.n561 VTAIL.n560 585
R207 VTAIL.n559 VTAIL.n558 585
R208 VTAIL.n512 VTAIL.n511 585
R209 VTAIL.n553 VTAIL.n552 585
R210 VTAIL.n551 VTAIL.n550 585
R211 VTAIL.n549 VTAIL.n515 585
R212 VTAIL.n519 VTAIL.n516 585
R213 VTAIL.n544 VTAIL.n543 585
R214 VTAIL.n542 VTAIL.n541 585
R215 VTAIL.n521 VTAIL.n520 585
R216 VTAIL.n536 VTAIL.n535 585
R217 VTAIL.n534 VTAIL.n533 585
R218 VTAIL.n525 VTAIL.n524 585
R219 VTAIL.n528 VTAIL.n527 585
R220 VTAIL.n493 VTAIL.n492 585
R221 VTAIL.n491 VTAIL.n490 585
R222 VTAIL.n420 VTAIL.n419 585
R223 VTAIL.n485 VTAIL.n484 585
R224 VTAIL.n483 VTAIL.n482 585
R225 VTAIL.n424 VTAIL.n423 585
R226 VTAIL.n477 VTAIL.n476 585
R227 VTAIL.n475 VTAIL.n474 585
R228 VTAIL.n428 VTAIL.n427 585
R229 VTAIL.n469 VTAIL.n468 585
R230 VTAIL.n467 VTAIL.n466 585
R231 VTAIL.n465 VTAIL.n431 585
R232 VTAIL.n435 VTAIL.n432 585
R233 VTAIL.n460 VTAIL.n459 585
R234 VTAIL.n458 VTAIL.n457 585
R235 VTAIL.n437 VTAIL.n436 585
R236 VTAIL.n452 VTAIL.n451 585
R237 VTAIL.n450 VTAIL.n449 585
R238 VTAIL.n441 VTAIL.n440 585
R239 VTAIL.n444 VTAIL.n443 585
R240 VTAIL.n411 VTAIL.n410 585
R241 VTAIL.n409 VTAIL.n408 585
R242 VTAIL.n338 VTAIL.n337 585
R243 VTAIL.n403 VTAIL.n402 585
R244 VTAIL.n401 VTAIL.n400 585
R245 VTAIL.n342 VTAIL.n341 585
R246 VTAIL.n395 VTAIL.n394 585
R247 VTAIL.n393 VTAIL.n392 585
R248 VTAIL.n346 VTAIL.n345 585
R249 VTAIL.n387 VTAIL.n386 585
R250 VTAIL.n385 VTAIL.n384 585
R251 VTAIL.n383 VTAIL.n349 585
R252 VTAIL.n353 VTAIL.n350 585
R253 VTAIL.n378 VTAIL.n377 585
R254 VTAIL.n376 VTAIL.n375 585
R255 VTAIL.n355 VTAIL.n354 585
R256 VTAIL.n370 VTAIL.n369 585
R257 VTAIL.n368 VTAIL.n367 585
R258 VTAIL.n359 VTAIL.n358 585
R259 VTAIL.n362 VTAIL.n361 585
R260 VTAIL.n327 VTAIL.n326 585
R261 VTAIL.n325 VTAIL.n324 585
R262 VTAIL.n254 VTAIL.n253 585
R263 VTAIL.n319 VTAIL.n318 585
R264 VTAIL.n317 VTAIL.n316 585
R265 VTAIL.n258 VTAIL.n257 585
R266 VTAIL.n311 VTAIL.n310 585
R267 VTAIL.n309 VTAIL.n308 585
R268 VTAIL.n262 VTAIL.n261 585
R269 VTAIL.n303 VTAIL.n302 585
R270 VTAIL.n301 VTAIL.n300 585
R271 VTAIL.n299 VTAIL.n265 585
R272 VTAIL.n269 VTAIL.n266 585
R273 VTAIL.n294 VTAIL.n293 585
R274 VTAIL.n292 VTAIL.n291 585
R275 VTAIL.n271 VTAIL.n270 585
R276 VTAIL.n286 VTAIL.n285 585
R277 VTAIL.n284 VTAIL.n283 585
R278 VTAIL.n275 VTAIL.n274 585
R279 VTAIL.n278 VTAIL.n277 585
R280 VTAIL.t14 VTAIL.n607 329.036
R281 VTAIL.t9 VTAIL.n27 329.036
R282 VTAIL.t0 VTAIL.n109 329.036
R283 VTAIL.t3 VTAIL.n193 329.036
R284 VTAIL.t7 VTAIL.n526 329.036
R285 VTAIL.t5 VTAIL.n442 329.036
R286 VTAIL.t11 VTAIL.n360 329.036
R287 VTAIL.t8 VTAIL.n276 329.036
R288 VTAIL.n608 VTAIL.n605 171.744
R289 VTAIL.n615 VTAIL.n605 171.744
R290 VTAIL.n616 VTAIL.n615 171.744
R291 VTAIL.n616 VTAIL.n601 171.744
R292 VTAIL.n623 VTAIL.n601 171.744
R293 VTAIL.n625 VTAIL.n623 171.744
R294 VTAIL.n625 VTAIL.n624 171.744
R295 VTAIL.n624 VTAIL.n597 171.744
R296 VTAIL.n633 VTAIL.n597 171.744
R297 VTAIL.n634 VTAIL.n633 171.744
R298 VTAIL.n634 VTAIL.n593 171.744
R299 VTAIL.n641 VTAIL.n593 171.744
R300 VTAIL.n642 VTAIL.n641 171.744
R301 VTAIL.n642 VTAIL.n589 171.744
R302 VTAIL.n649 VTAIL.n589 171.744
R303 VTAIL.n650 VTAIL.n649 171.744
R304 VTAIL.n650 VTAIL.n585 171.744
R305 VTAIL.n657 VTAIL.n585 171.744
R306 VTAIL.n658 VTAIL.n657 171.744
R307 VTAIL.n28 VTAIL.n25 171.744
R308 VTAIL.n35 VTAIL.n25 171.744
R309 VTAIL.n36 VTAIL.n35 171.744
R310 VTAIL.n36 VTAIL.n21 171.744
R311 VTAIL.n43 VTAIL.n21 171.744
R312 VTAIL.n45 VTAIL.n43 171.744
R313 VTAIL.n45 VTAIL.n44 171.744
R314 VTAIL.n44 VTAIL.n17 171.744
R315 VTAIL.n53 VTAIL.n17 171.744
R316 VTAIL.n54 VTAIL.n53 171.744
R317 VTAIL.n54 VTAIL.n13 171.744
R318 VTAIL.n61 VTAIL.n13 171.744
R319 VTAIL.n62 VTAIL.n61 171.744
R320 VTAIL.n62 VTAIL.n9 171.744
R321 VTAIL.n69 VTAIL.n9 171.744
R322 VTAIL.n70 VTAIL.n69 171.744
R323 VTAIL.n70 VTAIL.n5 171.744
R324 VTAIL.n77 VTAIL.n5 171.744
R325 VTAIL.n78 VTAIL.n77 171.744
R326 VTAIL.n110 VTAIL.n107 171.744
R327 VTAIL.n117 VTAIL.n107 171.744
R328 VTAIL.n118 VTAIL.n117 171.744
R329 VTAIL.n118 VTAIL.n103 171.744
R330 VTAIL.n125 VTAIL.n103 171.744
R331 VTAIL.n127 VTAIL.n125 171.744
R332 VTAIL.n127 VTAIL.n126 171.744
R333 VTAIL.n126 VTAIL.n99 171.744
R334 VTAIL.n135 VTAIL.n99 171.744
R335 VTAIL.n136 VTAIL.n135 171.744
R336 VTAIL.n136 VTAIL.n95 171.744
R337 VTAIL.n143 VTAIL.n95 171.744
R338 VTAIL.n144 VTAIL.n143 171.744
R339 VTAIL.n144 VTAIL.n91 171.744
R340 VTAIL.n151 VTAIL.n91 171.744
R341 VTAIL.n152 VTAIL.n151 171.744
R342 VTAIL.n152 VTAIL.n87 171.744
R343 VTAIL.n159 VTAIL.n87 171.744
R344 VTAIL.n160 VTAIL.n159 171.744
R345 VTAIL.n194 VTAIL.n191 171.744
R346 VTAIL.n201 VTAIL.n191 171.744
R347 VTAIL.n202 VTAIL.n201 171.744
R348 VTAIL.n202 VTAIL.n187 171.744
R349 VTAIL.n209 VTAIL.n187 171.744
R350 VTAIL.n211 VTAIL.n209 171.744
R351 VTAIL.n211 VTAIL.n210 171.744
R352 VTAIL.n210 VTAIL.n183 171.744
R353 VTAIL.n219 VTAIL.n183 171.744
R354 VTAIL.n220 VTAIL.n219 171.744
R355 VTAIL.n220 VTAIL.n179 171.744
R356 VTAIL.n227 VTAIL.n179 171.744
R357 VTAIL.n228 VTAIL.n227 171.744
R358 VTAIL.n228 VTAIL.n175 171.744
R359 VTAIL.n235 VTAIL.n175 171.744
R360 VTAIL.n236 VTAIL.n235 171.744
R361 VTAIL.n236 VTAIL.n171 171.744
R362 VTAIL.n243 VTAIL.n171 171.744
R363 VTAIL.n244 VTAIL.n243 171.744
R364 VTAIL.n576 VTAIL.n575 171.744
R365 VTAIL.n575 VTAIL.n503 171.744
R366 VTAIL.n568 VTAIL.n503 171.744
R367 VTAIL.n568 VTAIL.n567 171.744
R368 VTAIL.n567 VTAIL.n507 171.744
R369 VTAIL.n560 VTAIL.n507 171.744
R370 VTAIL.n560 VTAIL.n559 171.744
R371 VTAIL.n559 VTAIL.n511 171.744
R372 VTAIL.n552 VTAIL.n511 171.744
R373 VTAIL.n552 VTAIL.n551 171.744
R374 VTAIL.n551 VTAIL.n515 171.744
R375 VTAIL.n519 VTAIL.n515 171.744
R376 VTAIL.n543 VTAIL.n519 171.744
R377 VTAIL.n543 VTAIL.n542 171.744
R378 VTAIL.n542 VTAIL.n520 171.744
R379 VTAIL.n535 VTAIL.n520 171.744
R380 VTAIL.n535 VTAIL.n534 171.744
R381 VTAIL.n534 VTAIL.n524 171.744
R382 VTAIL.n527 VTAIL.n524 171.744
R383 VTAIL.n492 VTAIL.n491 171.744
R384 VTAIL.n491 VTAIL.n419 171.744
R385 VTAIL.n484 VTAIL.n419 171.744
R386 VTAIL.n484 VTAIL.n483 171.744
R387 VTAIL.n483 VTAIL.n423 171.744
R388 VTAIL.n476 VTAIL.n423 171.744
R389 VTAIL.n476 VTAIL.n475 171.744
R390 VTAIL.n475 VTAIL.n427 171.744
R391 VTAIL.n468 VTAIL.n427 171.744
R392 VTAIL.n468 VTAIL.n467 171.744
R393 VTAIL.n467 VTAIL.n431 171.744
R394 VTAIL.n435 VTAIL.n431 171.744
R395 VTAIL.n459 VTAIL.n435 171.744
R396 VTAIL.n459 VTAIL.n458 171.744
R397 VTAIL.n458 VTAIL.n436 171.744
R398 VTAIL.n451 VTAIL.n436 171.744
R399 VTAIL.n451 VTAIL.n450 171.744
R400 VTAIL.n450 VTAIL.n440 171.744
R401 VTAIL.n443 VTAIL.n440 171.744
R402 VTAIL.n410 VTAIL.n409 171.744
R403 VTAIL.n409 VTAIL.n337 171.744
R404 VTAIL.n402 VTAIL.n337 171.744
R405 VTAIL.n402 VTAIL.n401 171.744
R406 VTAIL.n401 VTAIL.n341 171.744
R407 VTAIL.n394 VTAIL.n341 171.744
R408 VTAIL.n394 VTAIL.n393 171.744
R409 VTAIL.n393 VTAIL.n345 171.744
R410 VTAIL.n386 VTAIL.n345 171.744
R411 VTAIL.n386 VTAIL.n385 171.744
R412 VTAIL.n385 VTAIL.n349 171.744
R413 VTAIL.n353 VTAIL.n349 171.744
R414 VTAIL.n377 VTAIL.n353 171.744
R415 VTAIL.n377 VTAIL.n376 171.744
R416 VTAIL.n376 VTAIL.n354 171.744
R417 VTAIL.n369 VTAIL.n354 171.744
R418 VTAIL.n369 VTAIL.n368 171.744
R419 VTAIL.n368 VTAIL.n358 171.744
R420 VTAIL.n361 VTAIL.n358 171.744
R421 VTAIL.n326 VTAIL.n325 171.744
R422 VTAIL.n325 VTAIL.n253 171.744
R423 VTAIL.n318 VTAIL.n253 171.744
R424 VTAIL.n318 VTAIL.n317 171.744
R425 VTAIL.n317 VTAIL.n257 171.744
R426 VTAIL.n310 VTAIL.n257 171.744
R427 VTAIL.n310 VTAIL.n309 171.744
R428 VTAIL.n309 VTAIL.n261 171.744
R429 VTAIL.n302 VTAIL.n261 171.744
R430 VTAIL.n302 VTAIL.n301 171.744
R431 VTAIL.n301 VTAIL.n265 171.744
R432 VTAIL.n269 VTAIL.n265 171.744
R433 VTAIL.n293 VTAIL.n269 171.744
R434 VTAIL.n293 VTAIL.n292 171.744
R435 VTAIL.n292 VTAIL.n270 171.744
R436 VTAIL.n285 VTAIL.n270 171.744
R437 VTAIL.n285 VTAIL.n284 171.744
R438 VTAIL.n284 VTAIL.n274 171.744
R439 VTAIL.n277 VTAIL.n274 171.744
R440 VTAIL.n608 VTAIL.t14 85.8723
R441 VTAIL.n28 VTAIL.t9 85.8723
R442 VTAIL.n110 VTAIL.t0 85.8723
R443 VTAIL.n194 VTAIL.t3 85.8723
R444 VTAIL.n527 VTAIL.t7 85.8723
R445 VTAIL.n443 VTAIL.t5 85.8723
R446 VTAIL.n361 VTAIL.t11 85.8723
R447 VTAIL.n277 VTAIL.t8 85.8723
R448 VTAIL.n499 VTAIL.n498 52.8253
R449 VTAIL.n333 VTAIL.n332 52.8253
R450 VTAIL.n1 VTAIL.n0 52.8251
R451 VTAIL.n167 VTAIL.n166 52.8251
R452 VTAIL.n663 VTAIL.n662 30.6338
R453 VTAIL.n83 VTAIL.n82 30.6338
R454 VTAIL.n165 VTAIL.n164 30.6338
R455 VTAIL.n249 VTAIL.n248 30.6338
R456 VTAIL.n581 VTAIL.n580 30.6338
R457 VTAIL.n497 VTAIL.n496 30.6338
R458 VTAIL.n415 VTAIL.n414 30.6338
R459 VTAIL.n331 VTAIL.n330 30.6338
R460 VTAIL.n663 VTAIL.n581 28.0652
R461 VTAIL.n331 VTAIL.n249 28.0652
R462 VTAIL.n632 VTAIL.n631 13.1884
R463 VTAIL.n52 VTAIL.n51 13.1884
R464 VTAIL.n134 VTAIL.n133 13.1884
R465 VTAIL.n218 VTAIL.n217 13.1884
R466 VTAIL.n550 VTAIL.n549 13.1884
R467 VTAIL.n466 VTAIL.n465 13.1884
R468 VTAIL.n384 VTAIL.n383 13.1884
R469 VTAIL.n300 VTAIL.n299 13.1884
R470 VTAIL.n630 VTAIL.n598 12.8005
R471 VTAIL.n635 VTAIL.n596 12.8005
R472 VTAIL.n50 VTAIL.n18 12.8005
R473 VTAIL.n55 VTAIL.n16 12.8005
R474 VTAIL.n132 VTAIL.n100 12.8005
R475 VTAIL.n137 VTAIL.n98 12.8005
R476 VTAIL.n216 VTAIL.n184 12.8005
R477 VTAIL.n221 VTAIL.n182 12.8005
R478 VTAIL.n553 VTAIL.n514 12.8005
R479 VTAIL.n548 VTAIL.n516 12.8005
R480 VTAIL.n469 VTAIL.n430 12.8005
R481 VTAIL.n464 VTAIL.n432 12.8005
R482 VTAIL.n387 VTAIL.n348 12.8005
R483 VTAIL.n382 VTAIL.n350 12.8005
R484 VTAIL.n303 VTAIL.n264 12.8005
R485 VTAIL.n298 VTAIL.n266 12.8005
R486 VTAIL.n627 VTAIL.n626 12.0247
R487 VTAIL.n636 VTAIL.n594 12.0247
R488 VTAIL.n47 VTAIL.n46 12.0247
R489 VTAIL.n56 VTAIL.n14 12.0247
R490 VTAIL.n129 VTAIL.n128 12.0247
R491 VTAIL.n138 VTAIL.n96 12.0247
R492 VTAIL.n213 VTAIL.n212 12.0247
R493 VTAIL.n222 VTAIL.n180 12.0247
R494 VTAIL.n554 VTAIL.n512 12.0247
R495 VTAIL.n545 VTAIL.n544 12.0247
R496 VTAIL.n470 VTAIL.n428 12.0247
R497 VTAIL.n461 VTAIL.n460 12.0247
R498 VTAIL.n388 VTAIL.n346 12.0247
R499 VTAIL.n379 VTAIL.n378 12.0247
R500 VTAIL.n304 VTAIL.n262 12.0247
R501 VTAIL.n295 VTAIL.n294 12.0247
R502 VTAIL.n622 VTAIL.n600 11.249
R503 VTAIL.n640 VTAIL.n639 11.249
R504 VTAIL.n42 VTAIL.n20 11.249
R505 VTAIL.n60 VTAIL.n59 11.249
R506 VTAIL.n124 VTAIL.n102 11.249
R507 VTAIL.n142 VTAIL.n141 11.249
R508 VTAIL.n208 VTAIL.n186 11.249
R509 VTAIL.n226 VTAIL.n225 11.249
R510 VTAIL.n558 VTAIL.n557 11.249
R511 VTAIL.n541 VTAIL.n518 11.249
R512 VTAIL.n474 VTAIL.n473 11.249
R513 VTAIL.n457 VTAIL.n434 11.249
R514 VTAIL.n392 VTAIL.n391 11.249
R515 VTAIL.n375 VTAIL.n352 11.249
R516 VTAIL.n308 VTAIL.n307 11.249
R517 VTAIL.n291 VTAIL.n268 11.249
R518 VTAIL.n609 VTAIL.n607 10.7239
R519 VTAIL.n29 VTAIL.n27 10.7239
R520 VTAIL.n111 VTAIL.n109 10.7239
R521 VTAIL.n195 VTAIL.n193 10.7239
R522 VTAIL.n528 VTAIL.n526 10.7239
R523 VTAIL.n444 VTAIL.n442 10.7239
R524 VTAIL.n362 VTAIL.n360 10.7239
R525 VTAIL.n278 VTAIL.n276 10.7239
R526 VTAIL.n621 VTAIL.n602 10.4732
R527 VTAIL.n643 VTAIL.n592 10.4732
R528 VTAIL.n41 VTAIL.n22 10.4732
R529 VTAIL.n63 VTAIL.n12 10.4732
R530 VTAIL.n123 VTAIL.n104 10.4732
R531 VTAIL.n145 VTAIL.n94 10.4732
R532 VTAIL.n207 VTAIL.n188 10.4732
R533 VTAIL.n229 VTAIL.n178 10.4732
R534 VTAIL.n561 VTAIL.n510 10.4732
R535 VTAIL.n540 VTAIL.n521 10.4732
R536 VTAIL.n477 VTAIL.n426 10.4732
R537 VTAIL.n456 VTAIL.n437 10.4732
R538 VTAIL.n395 VTAIL.n344 10.4732
R539 VTAIL.n374 VTAIL.n355 10.4732
R540 VTAIL.n311 VTAIL.n260 10.4732
R541 VTAIL.n290 VTAIL.n271 10.4732
R542 VTAIL.n618 VTAIL.n617 9.69747
R543 VTAIL.n644 VTAIL.n590 9.69747
R544 VTAIL.n38 VTAIL.n37 9.69747
R545 VTAIL.n64 VTAIL.n10 9.69747
R546 VTAIL.n120 VTAIL.n119 9.69747
R547 VTAIL.n146 VTAIL.n92 9.69747
R548 VTAIL.n204 VTAIL.n203 9.69747
R549 VTAIL.n230 VTAIL.n176 9.69747
R550 VTAIL.n562 VTAIL.n508 9.69747
R551 VTAIL.n537 VTAIL.n536 9.69747
R552 VTAIL.n478 VTAIL.n424 9.69747
R553 VTAIL.n453 VTAIL.n452 9.69747
R554 VTAIL.n396 VTAIL.n342 9.69747
R555 VTAIL.n371 VTAIL.n370 9.69747
R556 VTAIL.n312 VTAIL.n258 9.69747
R557 VTAIL.n287 VTAIL.n286 9.69747
R558 VTAIL.n662 VTAIL.n661 9.45567
R559 VTAIL.n82 VTAIL.n81 9.45567
R560 VTAIL.n164 VTAIL.n163 9.45567
R561 VTAIL.n248 VTAIL.n247 9.45567
R562 VTAIL.n580 VTAIL.n579 9.45567
R563 VTAIL.n496 VTAIL.n495 9.45567
R564 VTAIL.n414 VTAIL.n413 9.45567
R565 VTAIL.n330 VTAIL.n329 9.45567
R566 VTAIL.n655 VTAIL.n654 9.3005
R567 VTAIL.n584 VTAIL.n583 9.3005
R568 VTAIL.n661 VTAIL.n660 9.3005
R569 VTAIL.n588 VTAIL.n587 9.3005
R570 VTAIL.n647 VTAIL.n646 9.3005
R571 VTAIL.n645 VTAIL.n644 9.3005
R572 VTAIL.n592 VTAIL.n591 9.3005
R573 VTAIL.n639 VTAIL.n638 9.3005
R574 VTAIL.n637 VTAIL.n636 9.3005
R575 VTAIL.n596 VTAIL.n595 9.3005
R576 VTAIL.n611 VTAIL.n610 9.3005
R577 VTAIL.n613 VTAIL.n612 9.3005
R578 VTAIL.n604 VTAIL.n603 9.3005
R579 VTAIL.n619 VTAIL.n618 9.3005
R580 VTAIL.n621 VTAIL.n620 9.3005
R581 VTAIL.n600 VTAIL.n599 9.3005
R582 VTAIL.n628 VTAIL.n627 9.3005
R583 VTAIL.n630 VTAIL.n629 9.3005
R584 VTAIL.n653 VTAIL.n652 9.3005
R585 VTAIL.n75 VTAIL.n74 9.3005
R586 VTAIL.n4 VTAIL.n3 9.3005
R587 VTAIL.n81 VTAIL.n80 9.3005
R588 VTAIL.n8 VTAIL.n7 9.3005
R589 VTAIL.n67 VTAIL.n66 9.3005
R590 VTAIL.n65 VTAIL.n64 9.3005
R591 VTAIL.n12 VTAIL.n11 9.3005
R592 VTAIL.n59 VTAIL.n58 9.3005
R593 VTAIL.n57 VTAIL.n56 9.3005
R594 VTAIL.n16 VTAIL.n15 9.3005
R595 VTAIL.n31 VTAIL.n30 9.3005
R596 VTAIL.n33 VTAIL.n32 9.3005
R597 VTAIL.n24 VTAIL.n23 9.3005
R598 VTAIL.n39 VTAIL.n38 9.3005
R599 VTAIL.n41 VTAIL.n40 9.3005
R600 VTAIL.n20 VTAIL.n19 9.3005
R601 VTAIL.n48 VTAIL.n47 9.3005
R602 VTAIL.n50 VTAIL.n49 9.3005
R603 VTAIL.n73 VTAIL.n72 9.3005
R604 VTAIL.n157 VTAIL.n156 9.3005
R605 VTAIL.n86 VTAIL.n85 9.3005
R606 VTAIL.n163 VTAIL.n162 9.3005
R607 VTAIL.n90 VTAIL.n89 9.3005
R608 VTAIL.n149 VTAIL.n148 9.3005
R609 VTAIL.n147 VTAIL.n146 9.3005
R610 VTAIL.n94 VTAIL.n93 9.3005
R611 VTAIL.n141 VTAIL.n140 9.3005
R612 VTAIL.n139 VTAIL.n138 9.3005
R613 VTAIL.n98 VTAIL.n97 9.3005
R614 VTAIL.n113 VTAIL.n112 9.3005
R615 VTAIL.n115 VTAIL.n114 9.3005
R616 VTAIL.n106 VTAIL.n105 9.3005
R617 VTAIL.n121 VTAIL.n120 9.3005
R618 VTAIL.n123 VTAIL.n122 9.3005
R619 VTAIL.n102 VTAIL.n101 9.3005
R620 VTAIL.n130 VTAIL.n129 9.3005
R621 VTAIL.n132 VTAIL.n131 9.3005
R622 VTAIL.n155 VTAIL.n154 9.3005
R623 VTAIL.n241 VTAIL.n240 9.3005
R624 VTAIL.n170 VTAIL.n169 9.3005
R625 VTAIL.n247 VTAIL.n246 9.3005
R626 VTAIL.n174 VTAIL.n173 9.3005
R627 VTAIL.n233 VTAIL.n232 9.3005
R628 VTAIL.n231 VTAIL.n230 9.3005
R629 VTAIL.n178 VTAIL.n177 9.3005
R630 VTAIL.n225 VTAIL.n224 9.3005
R631 VTAIL.n223 VTAIL.n222 9.3005
R632 VTAIL.n182 VTAIL.n181 9.3005
R633 VTAIL.n197 VTAIL.n196 9.3005
R634 VTAIL.n199 VTAIL.n198 9.3005
R635 VTAIL.n190 VTAIL.n189 9.3005
R636 VTAIL.n205 VTAIL.n204 9.3005
R637 VTAIL.n207 VTAIL.n206 9.3005
R638 VTAIL.n186 VTAIL.n185 9.3005
R639 VTAIL.n214 VTAIL.n213 9.3005
R640 VTAIL.n216 VTAIL.n215 9.3005
R641 VTAIL.n239 VTAIL.n238 9.3005
R642 VTAIL.n502 VTAIL.n501 9.3005
R643 VTAIL.n573 VTAIL.n572 9.3005
R644 VTAIL.n571 VTAIL.n570 9.3005
R645 VTAIL.n506 VTAIL.n505 9.3005
R646 VTAIL.n565 VTAIL.n564 9.3005
R647 VTAIL.n563 VTAIL.n562 9.3005
R648 VTAIL.n510 VTAIL.n509 9.3005
R649 VTAIL.n557 VTAIL.n556 9.3005
R650 VTAIL.n555 VTAIL.n554 9.3005
R651 VTAIL.n514 VTAIL.n513 9.3005
R652 VTAIL.n548 VTAIL.n547 9.3005
R653 VTAIL.n546 VTAIL.n545 9.3005
R654 VTAIL.n518 VTAIL.n517 9.3005
R655 VTAIL.n540 VTAIL.n539 9.3005
R656 VTAIL.n538 VTAIL.n537 9.3005
R657 VTAIL.n523 VTAIL.n522 9.3005
R658 VTAIL.n532 VTAIL.n531 9.3005
R659 VTAIL.n530 VTAIL.n529 9.3005
R660 VTAIL.n579 VTAIL.n578 9.3005
R661 VTAIL.n446 VTAIL.n445 9.3005
R662 VTAIL.n448 VTAIL.n447 9.3005
R663 VTAIL.n439 VTAIL.n438 9.3005
R664 VTAIL.n454 VTAIL.n453 9.3005
R665 VTAIL.n456 VTAIL.n455 9.3005
R666 VTAIL.n434 VTAIL.n433 9.3005
R667 VTAIL.n462 VTAIL.n461 9.3005
R668 VTAIL.n464 VTAIL.n463 9.3005
R669 VTAIL.n418 VTAIL.n417 9.3005
R670 VTAIL.n495 VTAIL.n494 9.3005
R671 VTAIL.n489 VTAIL.n488 9.3005
R672 VTAIL.n487 VTAIL.n486 9.3005
R673 VTAIL.n422 VTAIL.n421 9.3005
R674 VTAIL.n481 VTAIL.n480 9.3005
R675 VTAIL.n479 VTAIL.n478 9.3005
R676 VTAIL.n426 VTAIL.n425 9.3005
R677 VTAIL.n473 VTAIL.n472 9.3005
R678 VTAIL.n471 VTAIL.n470 9.3005
R679 VTAIL.n430 VTAIL.n429 9.3005
R680 VTAIL.n364 VTAIL.n363 9.3005
R681 VTAIL.n366 VTAIL.n365 9.3005
R682 VTAIL.n357 VTAIL.n356 9.3005
R683 VTAIL.n372 VTAIL.n371 9.3005
R684 VTAIL.n374 VTAIL.n373 9.3005
R685 VTAIL.n352 VTAIL.n351 9.3005
R686 VTAIL.n380 VTAIL.n379 9.3005
R687 VTAIL.n382 VTAIL.n381 9.3005
R688 VTAIL.n336 VTAIL.n335 9.3005
R689 VTAIL.n413 VTAIL.n412 9.3005
R690 VTAIL.n407 VTAIL.n406 9.3005
R691 VTAIL.n405 VTAIL.n404 9.3005
R692 VTAIL.n340 VTAIL.n339 9.3005
R693 VTAIL.n399 VTAIL.n398 9.3005
R694 VTAIL.n397 VTAIL.n396 9.3005
R695 VTAIL.n344 VTAIL.n343 9.3005
R696 VTAIL.n391 VTAIL.n390 9.3005
R697 VTAIL.n389 VTAIL.n388 9.3005
R698 VTAIL.n348 VTAIL.n347 9.3005
R699 VTAIL.n280 VTAIL.n279 9.3005
R700 VTAIL.n282 VTAIL.n281 9.3005
R701 VTAIL.n273 VTAIL.n272 9.3005
R702 VTAIL.n288 VTAIL.n287 9.3005
R703 VTAIL.n290 VTAIL.n289 9.3005
R704 VTAIL.n268 VTAIL.n267 9.3005
R705 VTAIL.n296 VTAIL.n295 9.3005
R706 VTAIL.n298 VTAIL.n297 9.3005
R707 VTAIL.n252 VTAIL.n251 9.3005
R708 VTAIL.n329 VTAIL.n328 9.3005
R709 VTAIL.n323 VTAIL.n322 9.3005
R710 VTAIL.n321 VTAIL.n320 9.3005
R711 VTAIL.n256 VTAIL.n255 9.3005
R712 VTAIL.n315 VTAIL.n314 9.3005
R713 VTAIL.n313 VTAIL.n312 9.3005
R714 VTAIL.n260 VTAIL.n259 9.3005
R715 VTAIL.n307 VTAIL.n306 9.3005
R716 VTAIL.n305 VTAIL.n304 9.3005
R717 VTAIL.n264 VTAIL.n263 9.3005
R718 VTAIL.n614 VTAIL.n604 8.92171
R719 VTAIL.n648 VTAIL.n647 8.92171
R720 VTAIL.n662 VTAIL.n582 8.92171
R721 VTAIL.n34 VTAIL.n24 8.92171
R722 VTAIL.n68 VTAIL.n67 8.92171
R723 VTAIL.n82 VTAIL.n2 8.92171
R724 VTAIL.n116 VTAIL.n106 8.92171
R725 VTAIL.n150 VTAIL.n149 8.92171
R726 VTAIL.n164 VTAIL.n84 8.92171
R727 VTAIL.n200 VTAIL.n190 8.92171
R728 VTAIL.n234 VTAIL.n233 8.92171
R729 VTAIL.n248 VTAIL.n168 8.92171
R730 VTAIL.n580 VTAIL.n500 8.92171
R731 VTAIL.n566 VTAIL.n565 8.92171
R732 VTAIL.n533 VTAIL.n523 8.92171
R733 VTAIL.n496 VTAIL.n416 8.92171
R734 VTAIL.n482 VTAIL.n481 8.92171
R735 VTAIL.n449 VTAIL.n439 8.92171
R736 VTAIL.n414 VTAIL.n334 8.92171
R737 VTAIL.n400 VTAIL.n399 8.92171
R738 VTAIL.n367 VTAIL.n357 8.92171
R739 VTAIL.n330 VTAIL.n250 8.92171
R740 VTAIL.n316 VTAIL.n315 8.92171
R741 VTAIL.n283 VTAIL.n273 8.92171
R742 VTAIL.n613 VTAIL.n606 8.14595
R743 VTAIL.n651 VTAIL.n588 8.14595
R744 VTAIL.n660 VTAIL.n659 8.14595
R745 VTAIL.n33 VTAIL.n26 8.14595
R746 VTAIL.n71 VTAIL.n8 8.14595
R747 VTAIL.n80 VTAIL.n79 8.14595
R748 VTAIL.n115 VTAIL.n108 8.14595
R749 VTAIL.n153 VTAIL.n90 8.14595
R750 VTAIL.n162 VTAIL.n161 8.14595
R751 VTAIL.n199 VTAIL.n192 8.14595
R752 VTAIL.n237 VTAIL.n174 8.14595
R753 VTAIL.n246 VTAIL.n245 8.14595
R754 VTAIL.n578 VTAIL.n577 8.14595
R755 VTAIL.n569 VTAIL.n506 8.14595
R756 VTAIL.n532 VTAIL.n525 8.14595
R757 VTAIL.n494 VTAIL.n493 8.14595
R758 VTAIL.n485 VTAIL.n422 8.14595
R759 VTAIL.n448 VTAIL.n441 8.14595
R760 VTAIL.n412 VTAIL.n411 8.14595
R761 VTAIL.n403 VTAIL.n340 8.14595
R762 VTAIL.n366 VTAIL.n359 8.14595
R763 VTAIL.n328 VTAIL.n327 8.14595
R764 VTAIL.n319 VTAIL.n256 8.14595
R765 VTAIL.n282 VTAIL.n275 8.14595
R766 VTAIL.n610 VTAIL.n609 7.3702
R767 VTAIL.n652 VTAIL.n586 7.3702
R768 VTAIL.n656 VTAIL.n584 7.3702
R769 VTAIL.n30 VTAIL.n29 7.3702
R770 VTAIL.n72 VTAIL.n6 7.3702
R771 VTAIL.n76 VTAIL.n4 7.3702
R772 VTAIL.n112 VTAIL.n111 7.3702
R773 VTAIL.n154 VTAIL.n88 7.3702
R774 VTAIL.n158 VTAIL.n86 7.3702
R775 VTAIL.n196 VTAIL.n195 7.3702
R776 VTAIL.n238 VTAIL.n172 7.3702
R777 VTAIL.n242 VTAIL.n170 7.3702
R778 VTAIL.n574 VTAIL.n502 7.3702
R779 VTAIL.n570 VTAIL.n504 7.3702
R780 VTAIL.n529 VTAIL.n528 7.3702
R781 VTAIL.n490 VTAIL.n418 7.3702
R782 VTAIL.n486 VTAIL.n420 7.3702
R783 VTAIL.n445 VTAIL.n444 7.3702
R784 VTAIL.n408 VTAIL.n336 7.3702
R785 VTAIL.n404 VTAIL.n338 7.3702
R786 VTAIL.n363 VTAIL.n362 7.3702
R787 VTAIL.n324 VTAIL.n252 7.3702
R788 VTAIL.n320 VTAIL.n254 7.3702
R789 VTAIL.n279 VTAIL.n278 7.3702
R790 VTAIL.n655 VTAIL.n586 6.59444
R791 VTAIL.n656 VTAIL.n655 6.59444
R792 VTAIL.n75 VTAIL.n6 6.59444
R793 VTAIL.n76 VTAIL.n75 6.59444
R794 VTAIL.n157 VTAIL.n88 6.59444
R795 VTAIL.n158 VTAIL.n157 6.59444
R796 VTAIL.n241 VTAIL.n172 6.59444
R797 VTAIL.n242 VTAIL.n241 6.59444
R798 VTAIL.n574 VTAIL.n573 6.59444
R799 VTAIL.n573 VTAIL.n504 6.59444
R800 VTAIL.n490 VTAIL.n489 6.59444
R801 VTAIL.n489 VTAIL.n420 6.59444
R802 VTAIL.n408 VTAIL.n407 6.59444
R803 VTAIL.n407 VTAIL.n338 6.59444
R804 VTAIL.n324 VTAIL.n323 6.59444
R805 VTAIL.n323 VTAIL.n254 6.59444
R806 VTAIL.n610 VTAIL.n606 5.81868
R807 VTAIL.n652 VTAIL.n651 5.81868
R808 VTAIL.n659 VTAIL.n584 5.81868
R809 VTAIL.n30 VTAIL.n26 5.81868
R810 VTAIL.n72 VTAIL.n71 5.81868
R811 VTAIL.n79 VTAIL.n4 5.81868
R812 VTAIL.n112 VTAIL.n108 5.81868
R813 VTAIL.n154 VTAIL.n153 5.81868
R814 VTAIL.n161 VTAIL.n86 5.81868
R815 VTAIL.n196 VTAIL.n192 5.81868
R816 VTAIL.n238 VTAIL.n237 5.81868
R817 VTAIL.n245 VTAIL.n170 5.81868
R818 VTAIL.n577 VTAIL.n502 5.81868
R819 VTAIL.n570 VTAIL.n569 5.81868
R820 VTAIL.n529 VTAIL.n525 5.81868
R821 VTAIL.n493 VTAIL.n418 5.81868
R822 VTAIL.n486 VTAIL.n485 5.81868
R823 VTAIL.n445 VTAIL.n441 5.81868
R824 VTAIL.n411 VTAIL.n336 5.81868
R825 VTAIL.n404 VTAIL.n403 5.81868
R826 VTAIL.n363 VTAIL.n359 5.81868
R827 VTAIL.n327 VTAIL.n252 5.81868
R828 VTAIL.n320 VTAIL.n319 5.81868
R829 VTAIL.n279 VTAIL.n275 5.81868
R830 VTAIL.n614 VTAIL.n613 5.04292
R831 VTAIL.n648 VTAIL.n588 5.04292
R832 VTAIL.n660 VTAIL.n582 5.04292
R833 VTAIL.n34 VTAIL.n33 5.04292
R834 VTAIL.n68 VTAIL.n8 5.04292
R835 VTAIL.n80 VTAIL.n2 5.04292
R836 VTAIL.n116 VTAIL.n115 5.04292
R837 VTAIL.n150 VTAIL.n90 5.04292
R838 VTAIL.n162 VTAIL.n84 5.04292
R839 VTAIL.n200 VTAIL.n199 5.04292
R840 VTAIL.n234 VTAIL.n174 5.04292
R841 VTAIL.n246 VTAIL.n168 5.04292
R842 VTAIL.n578 VTAIL.n500 5.04292
R843 VTAIL.n566 VTAIL.n506 5.04292
R844 VTAIL.n533 VTAIL.n532 5.04292
R845 VTAIL.n494 VTAIL.n416 5.04292
R846 VTAIL.n482 VTAIL.n422 5.04292
R847 VTAIL.n449 VTAIL.n448 5.04292
R848 VTAIL.n412 VTAIL.n334 5.04292
R849 VTAIL.n400 VTAIL.n340 5.04292
R850 VTAIL.n367 VTAIL.n366 5.04292
R851 VTAIL.n328 VTAIL.n250 5.04292
R852 VTAIL.n316 VTAIL.n256 5.04292
R853 VTAIL.n283 VTAIL.n282 5.04292
R854 VTAIL.n617 VTAIL.n604 4.26717
R855 VTAIL.n647 VTAIL.n590 4.26717
R856 VTAIL.n37 VTAIL.n24 4.26717
R857 VTAIL.n67 VTAIL.n10 4.26717
R858 VTAIL.n119 VTAIL.n106 4.26717
R859 VTAIL.n149 VTAIL.n92 4.26717
R860 VTAIL.n203 VTAIL.n190 4.26717
R861 VTAIL.n233 VTAIL.n176 4.26717
R862 VTAIL.n565 VTAIL.n508 4.26717
R863 VTAIL.n536 VTAIL.n523 4.26717
R864 VTAIL.n481 VTAIL.n424 4.26717
R865 VTAIL.n452 VTAIL.n439 4.26717
R866 VTAIL.n399 VTAIL.n342 4.26717
R867 VTAIL.n370 VTAIL.n357 4.26717
R868 VTAIL.n315 VTAIL.n258 4.26717
R869 VTAIL.n286 VTAIL.n273 4.26717
R870 VTAIL.n618 VTAIL.n602 3.49141
R871 VTAIL.n644 VTAIL.n643 3.49141
R872 VTAIL.n38 VTAIL.n22 3.49141
R873 VTAIL.n64 VTAIL.n63 3.49141
R874 VTAIL.n120 VTAIL.n104 3.49141
R875 VTAIL.n146 VTAIL.n145 3.49141
R876 VTAIL.n204 VTAIL.n188 3.49141
R877 VTAIL.n230 VTAIL.n229 3.49141
R878 VTAIL.n562 VTAIL.n561 3.49141
R879 VTAIL.n537 VTAIL.n521 3.49141
R880 VTAIL.n478 VTAIL.n477 3.49141
R881 VTAIL.n453 VTAIL.n437 3.49141
R882 VTAIL.n396 VTAIL.n395 3.49141
R883 VTAIL.n371 VTAIL.n355 3.49141
R884 VTAIL.n312 VTAIL.n311 3.49141
R885 VTAIL.n287 VTAIL.n271 3.49141
R886 VTAIL.n333 VTAIL.n331 2.83671
R887 VTAIL.n415 VTAIL.n333 2.83671
R888 VTAIL.n499 VTAIL.n497 2.83671
R889 VTAIL.n581 VTAIL.n499 2.83671
R890 VTAIL.n249 VTAIL.n167 2.83671
R891 VTAIL.n167 VTAIL.n165 2.83671
R892 VTAIL.n83 VTAIL.n1 2.83671
R893 VTAIL VTAIL.n663 2.77852
R894 VTAIL.n622 VTAIL.n621 2.71565
R895 VTAIL.n640 VTAIL.n592 2.71565
R896 VTAIL.n42 VTAIL.n41 2.71565
R897 VTAIL.n60 VTAIL.n12 2.71565
R898 VTAIL.n124 VTAIL.n123 2.71565
R899 VTAIL.n142 VTAIL.n94 2.71565
R900 VTAIL.n208 VTAIL.n207 2.71565
R901 VTAIL.n226 VTAIL.n178 2.71565
R902 VTAIL.n558 VTAIL.n510 2.71565
R903 VTAIL.n541 VTAIL.n540 2.71565
R904 VTAIL.n474 VTAIL.n426 2.71565
R905 VTAIL.n457 VTAIL.n456 2.71565
R906 VTAIL.n392 VTAIL.n344 2.71565
R907 VTAIL.n375 VTAIL.n374 2.71565
R908 VTAIL.n308 VTAIL.n260 2.71565
R909 VTAIL.n291 VTAIL.n290 2.71565
R910 VTAIL.n530 VTAIL.n526 2.41282
R911 VTAIL.n446 VTAIL.n442 2.41282
R912 VTAIL.n364 VTAIL.n360 2.41282
R913 VTAIL.n280 VTAIL.n276 2.41282
R914 VTAIL.n611 VTAIL.n607 2.41282
R915 VTAIL.n31 VTAIL.n27 2.41282
R916 VTAIL.n113 VTAIL.n109 2.41282
R917 VTAIL.n197 VTAIL.n193 2.41282
R918 VTAIL.n0 VTAIL.t13 2.17912
R919 VTAIL.n0 VTAIL.t12 2.17912
R920 VTAIL.n166 VTAIL.t6 2.17912
R921 VTAIL.n166 VTAIL.t4 2.17912
R922 VTAIL.n498 VTAIL.t1 2.17912
R923 VTAIL.n498 VTAIL.t2 2.17912
R924 VTAIL.n332 VTAIL.t10 2.17912
R925 VTAIL.n332 VTAIL.t15 2.17912
R926 VTAIL.n626 VTAIL.n600 1.93989
R927 VTAIL.n639 VTAIL.n594 1.93989
R928 VTAIL.n46 VTAIL.n20 1.93989
R929 VTAIL.n59 VTAIL.n14 1.93989
R930 VTAIL.n128 VTAIL.n102 1.93989
R931 VTAIL.n141 VTAIL.n96 1.93989
R932 VTAIL.n212 VTAIL.n186 1.93989
R933 VTAIL.n225 VTAIL.n180 1.93989
R934 VTAIL.n557 VTAIL.n512 1.93989
R935 VTAIL.n544 VTAIL.n518 1.93989
R936 VTAIL.n473 VTAIL.n428 1.93989
R937 VTAIL.n460 VTAIL.n434 1.93989
R938 VTAIL.n391 VTAIL.n346 1.93989
R939 VTAIL.n378 VTAIL.n352 1.93989
R940 VTAIL.n307 VTAIL.n262 1.93989
R941 VTAIL.n294 VTAIL.n268 1.93989
R942 VTAIL.n627 VTAIL.n598 1.16414
R943 VTAIL.n636 VTAIL.n635 1.16414
R944 VTAIL.n47 VTAIL.n18 1.16414
R945 VTAIL.n56 VTAIL.n55 1.16414
R946 VTAIL.n129 VTAIL.n100 1.16414
R947 VTAIL.n138 VTAIL.n137 1.16414
R948 VTAIL.n213 VTAIL.n184 1.16414
R949 VTAIL.n222 VTAIL.n221 1.16414
R950 VTAIL.n554 VTAIL.n553 1.16414
R951 VTAIL.n545 VTAIL.n516 1.16414
R952 VTAIL.n470 VTAIL.n469 1.16414
R953 VTAIL.n461 VTAIL.n432 1.16414
R954 VTAIL.n388 VTAIL.n387 1.16414
R955 VTAIL.n379 VTAIL.n350 1.16414
R956 VTAIL.n304 VTAIL.n303 1.16414
R957 VTAIL.n295 VTAIL.n266 1.16414
R958 VTAIL.n497 VTAIL.n415 0.470328
R959 VTAIL.n165 VTAIL.n83 0.470328
R960 VTAIL.n631 VTAIL.n630 0.388379
R961 VTAIL.n632 VTAIL.n596 0.388379
R962 VTAIL.n51 VTAIL.n50 0.388379
R963 VTAIL.n52 VTAIL.n16 0.388379
R964 VTAIL.n133 VTAIL.n132 0.388379
R965 VTAIL.n134 VTAIL.n98 0.388379
R966 VTAIL.n217 VTAIL.n216 0.388379
R967 VTAIL.n218 VTAIL.n182 0.388379
R968 VTAIL.n550 VTAIL.n514 0.388379
R969 VTAIL.n549 VTAIL.n548 0.388379
R970 VTAIL.n466 VTAIL.n430 0.388379
R971 VTAIL.n465 VTAIL.n464 0.388379
R972 VTAIL.n384 VTAIL.n348 0.388379
R973 VTAIL.n383 VTAIL.n382 0.388379
R974 VTAIL.n300 VTAIL.n264 0.388379
R975 VTAIL.n299 VTAIL.n298 0.388379
R976 VTAIL.n612 VTAIL.n611 0.155672
R977 VTAIL.n612 VTAIL.n603 0.155672
R978 VTAIL.n619 VTAIL.n603 0.155672
R979 VTAIL.n620 VTAIL.n619 0.155672
R980 VTAIL.n620 VTAIL.n599 0.155672
R981 VTAIL.n628 VTAIL.n599 0.155672
R982 VTAIL.n629 VTAIL.n628 0.155672
R983 VTAIL.n629 VTAIL.n595 0.155672
R984 VTAIL.n637 VTAIL.n595 0.155672
R985 VTAIL.n638 VTAIL.n637 0.155672
R986 VTAIL.n638 VTAIL.n591 0.155672
R987 VTAIL.n645 VTAIL.n591 0.155672
R988 VTAIL.n646 VTAIL.n645 0.155672
R989 VTAIL.n646 VTAIL.n587 0.155672
R990 VTAIL.n653 VTAIL.n587 0.155672
R991 VTAIL.n654 VTAIL.n653 0.155672
R992 VTAIL.n654 VTAIL.n583 0.155672
R993 VTAIL.n661 VTAIL.n583 0.155672
R994 VTAIL.n32 VTAIL.n31 0.155672
R995 VTAIL.n32 VTAIL.n23 0.155672
R996 VTAIL.n39 VTAIL.n23 0.155672
R997 VTAIL.n40 VTAIL.n39 0.155672
R998 VTAIL.n40 VTAIL.n19 0.155672
R999 VTAIL.n48 VTAIL.n19 0.155672
R1000 VTAIL.n49 VTAIL.n48 0.155672
R1001 VTAIL.n49 VTAIL.n15 0.155672
R1002 VTAIL.n57 VTAIL.n15 0.155672
R1003 VTAIL.n58 VTAIL.n57 0.155672
R1004 VTAIL.n58 VTAIL.n11 0.155672
R1005 VTAIL.n65 VTAIL.n11 0.155672
R1006 VTAIL.n66 VTAIL.n65 0.155672
R1007 VTAIL.n66 VTAIL.n7 0.155672
R1008 VTAIL.n73 VTAIL.n7 0.155672
R1009 VTAIL.n74 VTAIL.n73 0.155672
R1010 VTAIL.n74 VTAIL.n3 0.155672
R1011 VTAIL.n81 VTAIL.n3 0.155672
R1012 VTAIL.n114 VTAIL.n113 0.155672
R1013 VTAIL.n114 VTAIL.n105 0.155672
R1014 VTAIL.n121 VTAIL.n105 0.155672
R1015 VTAIL.n122 VTAIL.n121 0.155672
R1016 VTAIL.n122 VTAIL.n101 0.155672
R1017 VTAIL.n130 VTAIL.n101 0.155672
R1018 VTAIL.n131 VTAIL.n130 0.155672
R1019 VTAIL.n131 VTAIL.n97 0.155672
R1020 VTAIL.n139 VTAIL.n97 0.155672
R1021 VTAIL.n140 VTAIL.n139 0.155672
R1022 VTAIL.n140 VTAIL.n93 0.155672
R1023 VTAIL.n147 VTAIL.n93 0.155672
R1024 VTAIL.n148 VTAIL.n147 0.155672
R1025 VTAIL.n148 VTAIL.n89 0.155672
R1026 VTAIL.n155 VTAIL.n89 0.155672
R1027 VTAIL.n156 VTAIL.n155 0.155672
R1028 VTAIL.n156 VTAIL.n85 0.155672
R1029 VTAIL.n163 VTAIL.n85 0.155672
R1030 VTAIL.n198 VTAIL.n197 0.155672
R1031 VTAIL.n198 VTAIL.n189 0.155672
R1032 VTAIL.n205 VTAIL.n189 0.155672
R1033 VTAIL.n206 VTAIL.n205 0.155672
R1034 VTAIL.n206 VTAIL.n185 0.155672
R1035 VTAIL.n214 VTAIL.n185 0.155672
R1036 VTAIL.n215 VTAIL.n214 0.155672
R1037 VTAIL.n215 VTAIL.n181 0.155672
R1038 VTAIL.n223 VTAIL.n181 0.155672
R1039 VTAIL.n224 VTAIL.n223 0.155672
R1040 VTAIL.n224 VTAIL.n177 0.155672
R1041 VTAIL.n231 VTAIL.n177 0.155672
R1042 VTAIL.n232 VTAIL.n231 0.155672
R1043 VTAIL.n232 VTAIL.n173 0.155672
R1044 VTAIL.n239 VTAIL.n173 0.155672
R1045 VTAIL.n240 VTAIL.n239 0.155672
R1046 VTAIL.n240 VTAIL.n169 0.155672
R1047 VTAIL.n247 VTAIL.n169 0.155672
R1048 VTAIL.n579 VTAIL.n501 0.155672
R1049 VTAIL.n572 VTAIL.n501 0.155672
R1050 VTAIL.n572 VTAIL.n571 0.155672
R1051 VTAIL.n571 VTAIL.n505 0.155672
R1052 VTAIL.n564 VTAIL.n505 0.155672
R1053 VTAIL.n564 VTAIL.n563 0.155672
R1054 VTAIL.n563 VTAIL.n509 0.155672
R1055 VTAIL.n556 VTAIL.n509 0.155672
R1056 VTAIL.n556 VTAIL.n555 0.155672
R1057 VTAIL.n555 VTAIL.n513 0.155672
R1058 VTAIL.n547 VTAIL.n513 0.155672
R1059 VTAIL.n547 VTAIL.n546 0.155672
R1060 VTAIL.n546 VTAIL.n517 0.155672
R1061 VTAIL.n539 VTAIL.n517 0.155672
R1062 VTAIL.n539 VTAIL.n538 0.155672
R1063 VTAIL.n538 VTAIL.n522 0.155672
R1064 VTAIL.n531 VTAIL.n522 0.155672
R1065 VTAIL.n531 VTAIL.n530 0.155672
R1066 VTAIL.n495 VTAIL.n417 0.155672
R1067 VTAIL.n488 VTAIL.n417 0.155672
R1068 VTAIL.n488 VTAIL.n487 0.155672
R1069 VTAIL.n487 VTAIL.n421 0.155672
R1070 VTAIL.n480 VTAIL.n421 0.155672
R1071 VTAIL.n480 VTAIL.n479 0.155672
R1072 VTAIL.n479 VTAIL.n425 0.155672
R1073 VTAIL.n472 VTAIL.n425 0.155672
R1074 VTAIL.n472 VTAIL.n471 0.155672
R1075 VTAIL.n471 VTAIL.n429 0.155672
R1076 VTAIL.n463 VTAIL.n429 0.155672
R1077 VTAIL.n463 VTAIL.n462 0.155672
R1078 VTAIL.n462 VTAIL.n433 0.155672
R1079 VTAIL.n455 VTAIL.n433 0.155672
R1080 VTAIL.n455 VTAIL.n454 0.155672
R1081 VTAIL.n454 VTAIL.n438 0.155672
R1082 VTAIL.n447 VTAIL.n438 0.155672
R1083 VTAIL.n447 VTAIL.n446 0.155672
R1084 VTAIL.n413 VTAIL.n335 0.155672
R1085 VTAIL.n406 VTAIL.n335 0.155672
R1086 VTAIL.n406 VTAIL.n405 0.155672
R1087 VTAIL.n405 VTAIL.n339 0.155672
R1088 VTAIL.n398 VTAIL.n339 0.155672
R1089 VTAIL.n398 VTAIL.n397 0.155672
R1090 VTAIL.n397 VTAIL.n343 0.155672
R1091 VTAIL.n390 VTAIL.n343 0.155672
R1092 VTAIL.n390 VTAIL.n389 0.155672
R1093 VTAIL.n389 VTAIL.n347 0.155672
R1094 VTAIL.n381 VTAIL.n347 0.155672
R1095 VTAIL.n381 VTAIL.n380 0.155672
R1096 VTAIL.n380 VTAIL.n351 0.155672
R1097 VTAIL.n373 VTAIL.n351 0.155672
R1098 VTAIL.n373 VTAIL.n372 0.155672
R1099 VTAIL.n372 VTAIL.n356 0.155672
R1100 VTAIL.n365 VTAIL.n356 0.155672
R1101 VTAIL.n365 VTAIL.n364 0.155672
R1102 VTAIL.n329 VTAIL.n251 0.155672
R1103 VTAIL.n322 VTAIL.n251 0.155672
R1104 VTAIL.n322 VTAIL.n321 0.155672
R1105 VTAIL.n321 VTAIL.n255 0.155672
R1106 VTAIL.n314 VTAIL.n255 0.155672
R1107 VTAIL.n314 VTAIL.n313 0.155672
R1108 VTAIL.n313 VTAIL.n259 0.155672
R1109 VTAIL.n306 VTAIL.n259 0.155672
R1110 VTAIL.n306 VTAIL.n305 0.155672
R1111 VTAIL.n305 VTAIL.n263 0.155672
R1112 VTAIL.n297 VTAIL.n263 0.155672
R1113 VTAIL.n297 VTAIL.n296 0.155672
R1114 VTAIL.n296 VTAIL.n267 0.155672
R1115 VTAIL.n289 VTAIL.n267 0.155672
R1116 VTAIL.n289 VTAIL.n288 0.155672
R1117 VTAIL.n288 VTAIL.n272 0.155672
R1118 VTAIL.n281 VTAIL.n272 0.155672
R1119 VTAIL.n281 VTAIL.n280 0.155672
R1120 VTAIL VTAIL.n1 0.0586897
R1121 VP.n21 VP.n20 161.3
R1122 VP.n22 VP.n17 161.3
R1123 VP.n24 VP.n23 161.3
R1124 VP.n25 VP.n16 161.3
R1125 VP.n27 VP.n26 161.3
R1126 VP.n28 VP.n15 161.3
R1127 VP.n30 VP.n29 161.3
R1128 VP.n32 VP.n14 161.3
R1129 VP.n34 VP.n33 161.3
R1130 VP.n35 VP.n13 161.3
R1131 VP.n37 VP.n36 161.3
R1132 VP.n38 VP.n12 161.3
R1133 VP.n40 VP.n39 161.3
R1134 VP.n73 VP.n72 161.3
R1135 VP.n71 VP.n1 161.3
R1136 VP.n70 VP.n69 161.3
R1137 VP.n68 VP.n2 161.3
R1138 VP.n67 VP.n66 161.3
R1139 VP.n65 VP.n3 161.3
R1140 VP.n63 VP.n62 161.3
R1141 VP.n61 VP.n4 161.3
R1142 VP.n60 VP.n59 161.3
R1143 VP.n58 VP.n5 161.3
R1144 VP.n57 VP.n56 161.3
R1145 VP.n55 VP.n6 161.3
R1146 VP.n54 VP.n53 161.3
R1147 VP.n51 VP.n7 161.3
R1148 VP.n50 VP.n49 161.3
R1149 VP.n48 VP.n8 161.3
R1150 VP.n47 VP.n46 161.3
R1151 VP.n45 VP.n9 161.3
R1152 VP.n44 VP.n43 161.3
R1153 VP.n18 VP.t1 153.298
R1154 VP.n10 VP.t5 121.478
R1155 VP.n52 VP.t7 121.478
R1156 VP.n64 VP.t0 121.478
R1157 VP.n0 VP.t2 121.478
R1158 VP.n11 VP.t3 121.478
R1159 VP.n31 VP.t6 121.478
R1160 VP.n19 VP.t4 121.478
R1161 VP.n42 VP.n10 68.8507
R1162 VP.n74 VP.n0 68.8507
R1163 VP.n41 VP.n11 68.8507
R1164 VP.n19 VP.n18 66.845
R1165 VP.n46 VP.n8 56.5617
R1166 VP.n70 VP.n2 56.5617
R1167 VP.n37 VP.n13 56.5617
R1168 VP.n42 VP.n41 54.9238
R1169 VP.n58 VP.n57 40.577
R1170 VP.n59 VP.n58 40.577
R1171 VP.n26 VP.n25 40.577
R1172 VP.n25 VP.n24 40.577
R1173 VP.n45 VP.n44 24.5923
R1174 VP.n46 VP.n45 24.5923
R1175 VP.n50 VP.n8 24.5923
R1176 VP.n51 VP.n50 24.5923
R1177 VP.n53 VP.n6 24.5923
R1178 VP.n57 VP.n6 24.5923
R1179 VP.n59 VP.n4 24.5923
R1180 VP.n63 VP.n4 24.5923
R1181 VP.n66 VP.n65 24.5923
R1182 VP.n66 VP.n2 24.5923
R1183 VP.n71 VP.n70 24.5923
R1184 VP.n72 VP.n71 24.5923
R1185 VP.n38 VP.n37 24.5923
R1186 VP.n39 VP.n38 24.5923
R1187 VP.n26 VP.n15 24.5923
R1188 VP.n30 VP.n15 24.5923
R1189 VP.n33 VP.n32 24.5923
R1190 VP.n33 VP.n13 24.5923
R1191 VP.n20 VP.n17 24.5923
R1192 VP.n24 VP.n17 24.5923
R1193 VP.n44 VP.n10 21.3954
R1194 VP.n72 VP.n0 21.3954
R1195 VP.n39 VP.n11 21.3954
R1196 VP.n52 VP.n51 17.4607
R1197 VP.n65 VP.n64 17.4607
R1198 VP.n32 VP.n31 17.4607
R1199 VP.n53 VP.n52 7.13213
R1200 VP.n64 VP.n63 7.13213
R1201 VP.n31 VP.n30 7.13213
R1202 VP.n20 VP.n19 7.13213
R1203 VP.n21 VP.n18 5.44401
R1204 VP.n41 VP.n40 0.354861
R1205 VP.n43 VP.n42 0.354861
R1206 VP.n74 VP.n73 0.354861
R1207 VP VP.n74 0.267071
R1208 VP.n22 VP.n21 0.189894
R1209 VP.n23 VP.n22 0.189894
R1210 VP.n23 VP.n16 0.189894
R1211 VP.n27 VP.n16 0.189894
R1212 VP.n28 VP.n27 0.189894
R1213 VP.n29 VP.n28 0.189894
R1214 VP.n29 VP.n14 0.189894
R1215 VP.n34 VP.n14 0.189894
R1216 VP.n35 VP.n34 0.189894
R1217 VP.n36 VP.n35 0.189894
R1218 VP.n36 VP.n12 0.189894
R1219 VP.n40 VP.n12 0.189894
R1220 VP.n43 VP.n9 0.189894
R1221 VP.n47 VP.n9 0.189894
R1222 VP.n48 VP.n47 0.189894
R1223 VP.n49 VP.n48 0.189894
R1224 VP.n49 VP.n7 0.189894
R1225 VP.n54 VP.n7 0.189894
R1226 VP.n55 VP.n54 0.189894
R1227 VP.n56 VP.n55 0.189894
R1228 VP.n56 VP.n5 0.189894
R1229 VP.n60 VP.n5 0.189894
R1230 VP.n61 VP.n60 0.189894
R1231 VP.n62 VP.n61 0.189894
R1232 VP.n62 VP.n3 0.189894
R1233 VP.n67 VP.n3 0.189894
R1234 VP.n68 VP.n67 0.189894
R1235 VP.n69 VP.n68 0.189894
R1236 VP.n69 VP.n1 0.189894
R1237 VP.n73 VP.n1 0.189894
R1238 VDD1 VDD1.n0 70.9804
R1239 VDD1.n3 VDD1.n2 70.8667
R1240 VDD1.n3 VDD1.n1 70.8667
R1241 VDD1.n5 VDD1.n4 69.5041
R1242 VDD1.n5 VDD1.n3 49.9233
R1243 VDD1.n4 VDD1.t1 2.17912
R1244 VDD1.n4 VDD1.t4 2.17912
R1245 VDD1.n0 VDD1.t6 2.17912
R1246 VDD1.n0 VDD1.t3 2.17912
R1247 VDD1.n2 VDD1.t7 2.17912
R1248 VDD1.n2 VDD1.t5 2.17912
R1249 VDD1.n1 VDD1.t2 2.17912
R1250 VDD1.n1 VDD1.t0 2.17912
R1251 VDD1 VDD1.n5 1.36041
R1252 B.n482 B.n481 585
R1253 B.n480 B.n147 585
R1254 B.n479 B.n478 585
R1255 B.n477 B.n148 585
R1256 B.n476 B.n475 585
R1257 B.n474 B.n149 585
R1258 B.n473 B.n472 585
R1259 B.n471 B.n150 585
R1260 B.n470 B.n469 585
R1261 B.n468 B.n151 585
R1262 B.n467 B.n466 585
R1263 B.n465 B.n152 585
R1264 B.n464 B.n463 585
R1265 B.n462 B.n153 585
R1266 B.n461 B.n460 585
R1267 B.n459 B.n154 585
R1268 B.n458 B.n457 585
R1269 B.n456 B.n155 585
R1270 B.n455 B.n454 585
R1271 B.n453 B.n156 585
R1272 B.n452 B.n451 585
R1273 B.n450 B.n157 585
R1274 B.n449 B.n448 585
R1275 B.n447 B.n158 585
R1276 B.n446 B.n445 585
R1277 B.n444 B.n159 585
R1278 B.n443 B.n442 585
R1279 B.n441 B.n160 585
R1280 B.n440 B.n439 585
R1281 B.n438 B.n161 585
R1282 B.n437 B.n436 585
R1283 B.n435 B.n162 585
R1284 B.n434 B.n433 585
R1285 B.n432 B.n163 585
R1286 B.n431 B.n430 585
R1287 B.n429 B.n164 585
R1288 B.n428 B.n427 585
R1289 B.n426 B.n165 585
R1290 B.n425 B.n424 585
R1291 B.n423 B.n166 585
R1292 B.n422 B.n421 585
R1293 B.n420 B.n167 585
R1294 B.n419 B.n418 585
R1295 B.n417 B.n168 585
R1296 B.n416 B.n415 585
R1297 B.n414 B.n169 585
R1298 B.n413 B.n412 585
R1299 B.n411 B.n170 585
R1300 B.n410 B.n409 585
R1301 B.n408 B.n171 585
R1302 B.n406 B.n405 585
R1303 B.n404 B.n174 585
R1304 B.n403 B.n402 585
R1305 B.n401 B.n175 585
R1306 B.n400 B.n399 585
R1307 B.n398 B.n176 585
R1308 B.n397 B.n396 585
R1309 B.n395 B.n177 585
R1310 B.n394 B.n393 585
R1311 B.n392 B.n178 585
R1312 B.n391 B.n390 585
R1313 B.n386 B.n179 585
R1314 B.n385 B.n384 585
R1315 B.n383 B.n180 585
R1316 B.n382 B.n381 585
R1317 B.n380 B.n181 585
R1318 B.n379 B.n378 585
R1319 B.n377 B.n182 585
R1320 B.n376 B.n375 585
R1321 B.n374 B.n183 585
R1322 B.n373 B.n372 585
R1323 B.n371 B.n184 585
R1324 B.n370 B.n369 585
R1325 B.n368 B.n185 585
R1326 B.n367 B.n366 585
R1327 B.n365 B.n186 585
R1328 B.n364 B.n363 585
R1329 B.n362 B.n187 585
R1330 B.n361 B.n360 585
R1331 B.n359 B.n188 585
R1332 B.n358 B.n357 585
R1333 B.n356 B.n189 585
R1334 B.n355 B.n354 585
R1335 B.n353 B.n190 585
R1336 B.n352 B.n351 585
R1337 B.n350 B.n191 585
R1338 B.n349 B.n348 585
R1339 B.n347 B.n192 585
R1340 B.n346 B.n345 585
R1341 B.n344 B.n193 585
R1342 B.n343 B.n342 585
R1343 B.n341 B.n194 585
R1344 B.n340 B.n339 585
R1345 B.n338 B.n195 585
R1346 B.n337 B.n336 585
R1347 B.n335 B.n196 585
R1348 B.n334 B.n333 585
R1349 B.n332 B.n197 585
R1350 B.n331 B.n330 585
R1351 B.n329 B.n198 585
R1352 B.n328 B.n327 585
R1353 B.n326 B.n199 585
R1354 B.n325 B.n324 585
R1355 B.n323 B.n200 585
R1356 B.n322 B.n321 585
R1357 B.n320 B.n201 585
R1358 B.n319 B.n318 585
R1359 B.n317 B.n202 585
R1360 B.n316 B.n315 585
R1361 B.n314 B.n203 585
R1362 B.n483 B.n146 585
R1363 B.n485 B.n484 585
R1364 B.n486 B.n145 585
R1365 B.n488 B.n487 585
R1366 B.n489 B.n144 585
R1367 B.n491 B.n490 585
R1368 B.n492 B.n143 585
R1369 B.n494 B.n493 585
R1370 B.n495 B.n142 585
R1371 B.n497 B.n496 585
R1372 B.n498 B.n141 585
R1373 B.n500 B.n499 585
R1374 B.n501 B.n140 585
R1375 B.n503 B.n502 585
R1376 B.n504 B.n139 585
R1377 B.n506 B.n505 585
R1378 B.n507 B.n138 585
R1379 B.n509 B.n508 585
R1380 B.n510 B.n137 585
R1381 B.n512 B.n511 585
R1382 B.n513 B.n136 585
R1383 B.n515 B.n514 585
R1384 B.n516 B.n135 585
R1385 B.n518 B.n517 585
R1386 B.n519 B.n134 585
R1387 B.n521 B.n520 585
R1388 B.n522 B.n133 585
R1389 B.n524 B.n523 585
R1390 B.n525 B.n132 585
R1391 B.n527 B.n526 585
R1392 B.n528 B.n131 585
R1393 B.n530 B.n529 585
R1394 B.n531 B.n130 585
R1395 B.n533 B.n532 585
R1396 B.n534 B.n129 585
R1397 B.n536 B.n535 585
R1398 B.n537 B.n128 585
R1399 B.n539 B.n538 585
R1400 B.n540 B.n127 585
R1401 B.n542 B.n541 585
R1402 B.n543 B.n126 585
R1403 B.n545 B.n544 585
R1404 B.n546 B.n125 585
R1405 B.n548 B.n547 585
R1406 B.n549 B.n124 585
R1407 B.n551 B.n550 585
R1408 B.n552 B.n123 585
R1409 B.n554 B.n553 585
R1410 B.n555 B.n122 585
R1411 B.n557 B.n556 585
R1412 B.n558 B.n121 585
R1413 B.n560 B.n559 585
R1414 B.n561 B.n120 585
R1415 B.n563 B.n562 585
R1416 B.n564 B.n119 585
R1417 B.n566 B.n565 585
R1418 B.n567 B.n118 585
R1419 B.n569 B.n568 585
R1420 B.n570 B.n117 585
R1421 B.n572 B.n571 585
R1422 B.n573 B.n116 585
R1423 B.n575 B.n574 585
R1424 B.n576 B.n115 585
R1425 B.n578 B.n577 585
R1426 B.n579 B.n114 585
R1427 B.n581 B.n580 585
R1428 B.n582 B.n113 585
R1429 B.n584 B.n583 585
R1430 B.n585 B.n112 585
R1431 B.n587 B.n586 585
R1432 B.n588 B.n111 585
R1433 B.n590 B.n589 585
R1434 B.n591 B.n110 585
R1435 B.n593 B.n592 585
R1436 B.n594 B.n109 585
R1437 B.n596 B.n595 585
R1438 B.n597 B.n108 585
R1439 B.n599 B.n598 585
R1440 B.n600 B.n107 585
R1441 B.n602 B.n601 585
R1442 B.n603 B.n106 585
R1443 B.n605 B.n604 585
R1444 B.n606 B.n105 585
R1445 B.n608 B.n607 585
R1446 B.n609 B.n104 585
R1447 B.n611 B.n610 585
R1448 B.n612 B.n103 585
R1449 B.n614 B.n613 585
R1450 B.n615 B.n102 585
R1451 B.n617 B.n616 585
R1452 B.n618 B.n101 585
R1453 B.n620 B.n619 585
R1454 B.n621 B.n100 585
R1455 B.n623 B.n622 585
R1456 B.n624 B.n99 585
R1457 B.n626 B.n625 585
R1458 B.n627 B.n98 585
R1459 B.n629 B.n628 585
R1460 B.n630 B.n97 585
R1461 B.n632 B.n631 585
R1462 B.n633 B.n96 585
R1463 B.n635 B.n634 585
R1464 B.n636 B.n95 585
R1465 B.n638 B.n637 585
R1466 B.n639 B.n94 585
R1467 B.n641 B.n640 585
R1468 B.n642 B.n93 585
R1469 B.n644 B.n643 585
R1470 B.n645 B.n92 585
R1471 B.n647 B.n646 585
R1472 B.n648 B.n91 585
R1473 B.n650 B.n649 585
R1474 B.n651 B.n90 585
R1475 B.n653 B.n652 585
R1476 B.n819 B.n30 585
R1477 B.n818 B.n817 585
R1478 B.n816 B.n31 585
R1479 B.n815 B.n814 585
R1480 B.n813 B.n32 585
R1481 B.n812 B.n811 585
R1482 B.n810 B.n33 585
R1483 B.n809 B.n808 585
R1484 B.n807 B.n34 585
R1485 B.n806 B.n805 585
R1486 B.n804 B.n35 585
R1487 B.n803 B.n802 585
R1488 B.n801 B.n36 585
R1489 B.n800 B.n799 585
R1490 B.n798 B.n37 585
R1491 B.n797 B.n796 585
R1492 B.n795 B.n38 585
R1493 B.n794 B.n793 585
R1494 B.n792 B.n39 585
R1495 B.n791 B.n790 585
R1496 B.n789 B.n40 585
R1497 B.n788 B.n787 585
R1498 B.n786 B.n41 585
R1499 B.n785 B.n784 585
R1500 B.n783 B.n42 585
R1501 B.n782 B.n781 585
R1502 B.n780 B.n43 585
R1503 B.n779 B.n778 585
R1504 B.n777 B.n44 585
R1505 B.n776 B.n775 585
R1506 B.n774 B.n45 585
R1507 B.n773 B.n772 585
R1508 B.n771 B.n46 585
R1509 B.n770 B.n769 585
R1510 B.n768 B.n47 585
R1511 B.n767 B.n766 585
R1512 B.n765 B.n48 585
R1513 B.n764 B.n763 585
R1514 B.n762 B.n49 585
R1515 B.n761 B.n760 585
R1516 B.n759 B.n50 585
R1517 B.n758 B.n757 585
R1518 B.n756 B.n51 585
R1519 B.n755 B.n754 585
R1520 B.n753 B.n52 585
R1521 B.n752 B.n751 585
R1522 B.n750 B.n53 585
R1523 B.n749 B.n748 585
R1524 B.n747 B.n54 585
R1525 B.n746 B.n745 585
R1526 B.n743 B.n55 585
R1527 B.n742 B.n741 585
R1528 B.n740 B.n58 585
R1529 B.n739 B.n738 585
R1530 B.n737 B.n59 585
R1531 B.n736 B.n735 585
R1532 B.n734 B.n60 585
R1533 B.n733 B.n732 585
R1534 B.n731 B.n61 585
R1535 B.n730 B.n729 585
R1536 B.n728 B.n727 585
R1537 B.n726 B.n65 585
R1538 B.n725 B.n724 585
R1539 B.n723 B.n66 585
R1540 B.n722 B.n721 585
R1541 B.n720 B.n67 585
R1542 B.n719 B.n718 585
R1543 B.n717 B.n68 585
R1544 B.n716 B.n715 585
R1545 B.n714 B.n69 585
R1546 B.n713 B.n712 585
R1547 B.n711 B.n70 585
R1548 B.n710 B.n709 585
R1549 B.n708 B.n71 585
R1550 B.n707 B.n706 585
R1551 B.n705 B.n72 585
R1552 B.n704 B.n703 585
R1553 B.n702 B.n73 585
R1554 B.n701 B.n700 585
R1555 B.n699 B.n74 585
R1556 B.n698 B.n697 585
R1557 B.n696 B.n75 585
R1558 B.n695 B.n694 585
R1559 B.n693 B.n76 585
R1560 B.n692 B.n691 585
R1561 B.n690 B.n77 585
R1562 B.n689 B.n688 585
R1563 B.n687 B.n78 585
R1564 B.n686 B.n685 585
R1565 B.n684 B.n79 585
R1566 B.n683 B.n682 585
R1567 B.n681 B.n80 585
R1568 B.n680 B.n679 585
R1569 B.n678 B.n81 585
R1570 B.n677 B.n676 585
R1571 B.n675 B.n82 585
R1572 B.n674 B.n673 585
R1573 B.n672 B.n83 585
R1574 B.n671 B.n670 585
R1575 B.n669 B.n84 585
R1576 B.n668 B.n667 585
R1577 B.n666 B.n85 585
R1578 B.n665 B.n664 585
R1579 B.n663 B.n86 585
R1580 B.n662 B.n661 585
R1581 B.n660 B.n87 585
R1582 B.n659 B.n658 585
R1583 B.n657 B.n88 585
R1584 B.n656 B.n655 585
R1585 B.n654 B.n89 585
R1586 B.n821 B.n820 585
R1587 B.n822 B.n29 585
R1588 B.n824 B.n823 585
R1589 B.n825 B.n28 585
R1590 B.n827 B.n826 585
R1591 B.n828 B.n27 585
R1592 B.n830 B.n829 585
R1593 B.n831 B.n26 585
R1594 B.n833 B.n832 585
R1595 B.n834 B.n25 585
R1596 B.n836 B.n835 585
R1597 B.n837 B.n24 585
R1598 B.n839 B.n838 585
R1599 B.n840 B.n23 585
R1600 B.n842 B.n841 585
R1601 B.n843 B.n22 585
R1602 B.n845 B.n844 585
R1603 B.n846 B.n21 585
R1604 B.n848 B.n847 585
R1605 B.n849 B.n20 585
R1606 B.n851 B.n850 585
R1607 B.n852 B.n19 585
R1608 B.n854 B.n853 585
R1609 B.n855 B.n18 585
R1610 B.n857 B.n856 585
R1611 B.n858 B.n17 585
R1612 B.n860 B.n859 585
R1613 B.n861 B.n16 585
R1614 B.n863 B.n862 585
R1615 B.n864 B.n15 585
R1616 B.n866 B.n865 585
R1617 B.n867 B.n14 585
R1618 B.n869 B.n868 585
R1619 B.n870 B.n13 585
R1620 B.n872 B.n871 585
R1621 B.n873 B.n12 585
R1622 B.n875 B.n874 585
R1623 B.n876 B.n11 585
R1624 B.n878 B.n877 585
R1625 B.n879 B.n10 585
R1626 B.n881 B.n880 585
R1627 B.n882 B.n9 585
R1628 B.n884 B.n883 585
R1629 B.n885 B.n8 585
R1630 B.n887 B.n886 585
R1631 B.n888 B.n7 585
R1632 B.n890 B.n889 585
R1633 B.n891 B.n6 585
R1634 B.n893 B.n892 585
R1635 B.n894 B.n5 585
R1636 B.n896 B.n895 585
R1637 B.n897 B.n4 585
R1638 B.n899 B.n898 585
R1639 B.n900 B.n3 585
R1640 B.n902 B.n901 585
R1641 B.n903 B.n0 585
R1642 B.n2 B.n1 585
R1643 B.n232 B.n231 585
R1644 B.n233 B.n230 585
R1645 B.n235 B.n234 585
R1646 B.n236 B.n229 585
R1647 B.n238 B.n237 585
R1648 B.n239 B.n228 585
R1649 B.n241 B.n240 585
R1650 B.n242 B.n227 585
R1651 B.n244 B.n243 585
R1652 B.n245 B.n226 585
R1653 B.n247 B.n246 585
R1654 B.n248 B.n225 585
R1655 B.n250 B.n249 585
R1656 B.n251 B.n224 585
R1657 B.n253 B.n252 585
R1658 B.n254 B.n223 585
R1659 B.n256 B.n255 585
R1660 B.n257 B.n222 585
R1661 B.n259 B.n258 585
R1662 B.n260 B.n221 585
R1663 B.n262 B.n261 585
R1664 B.n263 B.n220 585
R1665 B.n265 B.n264 585
R1666 B.n266 B.n219 585
R1667 B.n268 B.n267 585
R1668 B.n269 B.n218 585
R1669 B.n271 B.n270 585
R1670 B.n272 B.n217 585
R1671 B.n274 B.n273 585
R1672 B.n275 B.n216 585
R1673 B.n277 B.n276 585
R1674 B.n278 B.n215 585
R1675 B.n280 B.n279 585
R1676 B.n281 B.n214 585
R1677 B.n283 B.n282 585
R1678 B.n284 B.n213 585
R1679 B.n286 B.n285 585
R1680 B.n287 B.n212 585
R1681 B.n289 B.n288 585
R1682 B.n290 B.n211 585
R1683 B.n292 B.n291 585
R1684 B.n293 B.n210 585
R1685 B.n295 B.n294 585
R1686 B.n296 B.n209 585
R1687 B.n298 B.n297 585
R1688 B.n299 B.n208 585
R1689 B.n301 B.n300 585
R1690 B.n302 B.n207 585
R1691 B.n304 B.n303 585
R1692 B.n305 B.n206 585
R1693 B.n307 B.n306 585
R1694 B.n308 B.n205 585
R1695 B.n310 B.n309 585
R1696 B.n311 B.n204 585
R1697 B.n313 B.n312 585
R1698 B.n312 B.n203 497.305
R1699 B.n483 B.n482 497.305
R1700 B.n652 B.n89 497.305
R1701 B.n820 B.n819 497.305
R1702 B.n172 B.t7 492.205
R1703 B.n62 B.t11 492.205
R1704 B.n387 B.t1 492.204
R1705 B.n56 B.t5 492.204
R1706 B.n173 B.t8 428.399
R1707 B.n63 B.t10 428.399
R1708 B.n388 B.t2 428.399
R1709 B.n57 B.t4 428.399
R1710 B.n387 B.t0 330.01
R1711 B.n172 B.t6 330.01
R1712 B.n62 B.t9 330.01
R1713 B.n56 B.t3 330.01
R1714 B.n905 B.n904 256.663
R1715 B.n904 B.n903 235.042
R1716 B.n904 B.n2 235.042
R1717 B.n316 B.n203 163.367
R1718 B.n317 B.n316 163.367
R1719 B.n318 B.n317 163.367
R1720 B.n318 B.n201 163.367
R1721 B.n322 B.n201 163.367
R1722 B.n323 B.n322 163.367
R1723 B.n324 B.n323 163.367
R1724 B.n324 B.n199 163.367
R1725 B.n328 B.n199 163.367
R1726 B.n329 B.n328 163.367
R1727 B.n330 B.n329 163.367
R1728 B.n330 B.n197 163.367
R1729 B.n334 B.n197 163.367
R1730 B.n335 B.n334 163.367
R1731 B.n336 B.n335 163.367
R1732 B.n336 B.n195 163.367
R1733 B.n340 B.n195 163.367
R1734 B.n341 B.n340 163.367
R1735 B.n342 B.n341 163.367
R1736 B.n342 B.n193 163.367
R1737 B.n346 B.n193 163.367
R1738 B.n347 B.n346 163.367
R1739 B.n348 B.n347 163.367
R1740 B.n348 B.n191 163.367
R1741 B.n352 B.n191 163.367
R1742 B.n353 B.n352 163.367
R1743 B.n354 B.n353 163.367
R1744 B.n354 B.n189 163.367
R1745 B.n358 B.n189 163.367
R1746 B.n359 B.n358 163.367
R1747 B.n360 B.n359 163.367
R1748 B.n360 B.n187 163.367
R1749 B.n364 B.n187 163.367
R1750 B.n365 B.n364 163.367
R1751 B.n366 B.n365 163.367
R1752 B.n366 B.n185 163.367
R1753 B.n370 B.n185 163.367
R1754 B.n371 B.n370 163.367
R1755 B.n372 B.n371 163.367
R1756 B.n372 B.n183 163.367
R1757 B.n376 B.n183 163.367
R1758 B.n377 B.n376 163.367
R1759 B.n378 B.n377 163.367
R1760 B.n378 B.n181 163.367
R1761 B.n382 B.n181 163.367
R1762 B.n383 B.n382 163.367
R1763 B.n384 B.n383 163.367
R1764 B.n384 B.n179 163.367
R1765 B.n391 B.n179 163.367
R1766 B.n392 B.n391 163.367
R1767 B.n393 B.n392 163.367
R1768 B.n393 B.n177 163.367
R1769 B.n397 B.n177 163.367
R1770 B.n398 B.n397 163.367
R1771 B.n399 B.n398 163.367
R1772 B.n399 B.n175 163.367
R1773 B.n403 B.n175 163.367
R1774 B.n404 B.n403 163.367
R1775 B.n405 B.n404 163.367
R1776 B.n405 B.n171 163.367
R1777 B.n410 B.n171 163.367
R1778 B.n411 B.n410 163.367
R1779 B.n412 B.n411 163.367
R1780 B.n412 B.n169 163.367
R1781 B.n416 B.n169 163.367
R1782 B.n417 B.n416 163.367
R1783 B.n418 B.n417 163.367
R1784 B.n418 B.n167 163.367
R1785 B.n422 B.n167 163.367
R1786 B.n423 B.n422 163.367
R1787 B.n424 B.n423 163.367
R1788 B.n424 B.n165 163.367
R1789 B.n428 B.n165 163.367
R1790 B.n429 B.n428 163.367
R1791 B.n430 B.n429 163.367
R1792 B.n430 B.n163 163.367
R1793 B.n434 B.n163 163.367
R1794 B.n435 B.n434 163.367
R1795 B.n436 B.n435 163.367
R1796 B.n436 B.n161 163.367
R1797 B.n440 B.n161 163.367
R1798 B.n441 B.n440 163.367
R1799 B.n442 B.n441 163.367
R1800 B.n442 B.n159 163.367
R1801 B.n446 B.n159 163.367
R1802 B.n447 B.n446 163.367
R1803 B.n448 B.n447 163.367
R1804 B.n448 B.n157 163.367
R1805 B.n452 B.n157 163.367
R1806 B.n453 B.n452 163.367
R1807 B.n454 B.n453 163.367
R1808 B.n454 B.n155 163.367
R1809 B.n458 B.n155 163.367
R1810 B.n459 B.n458 163.367
R1811 B.n460 B.n459 163.367
R1812 B.n460 B.n153 163.367
R1813 B.n464 B.n153 163.367
R1814 B.n465 B.n464 163.367
R1815 B.n466 B.n465 163.367
R1816 B.n466 B.n151 163.367
R1817 B.n470 B.n151 163.367
R1818 B.n471 B.n470 163.367
R1819 B.n472 B.n471 163.367
R1820 B.n472 B.n149 163.367
R1821 B.n476 B.n149 163.367
R1822 B.n477 B.n476 163.367
R1823 B.n478 B.n477 163.367
R1824 B.n478 B.n147 163.367
R1825 B.n482 B.n147 163.367
R1826 B.n652 B.n651 163.367
R1827 B.n651 B.n650 163.367
R1828 B.n650 B.n91 163.367
R1829 B.n646 B.n91 163.367
R1830 B.n646 B.n645 163.367
R1831 B.n645 B.n644 163.367
R1832 B.n644 B.n93 163.367
R1833 B.n640 B.n93 163.367
R1834 B.n640 B.n639 163.367
R1835 B.n639 B.n638 163.367
R1836 B.n638 B.n95 163.367
R1837 B.n634 B.n95 163.367
R1838 B.n634 B.n633 163.367
R1839 B.n633 B.n632 163.367
R1840 B.n632 B.n97 163.367
R1841 B.n628 B.n97 163.367
R1842 B.n628 B.n627 163.367
R1843 B.n627 B.n626 163.367
R1844 B.n626 B.n99 163.367
R1845 B.n622 B.n99 163.367
R1846 B.n622 B.n621 163.367
R1847 B.n621 B.n620 163.367
R1848 B.n620 B.n101 163.367
R1849 B.n616 B.n101 163.367
R1850 B.n616 B.n615 163.367
R1851 B.n615 B.n614 163.367
R1852 B.n614 B.n103 163.367
R1853 B.n610 B.n103 163.367
R1854 B.n610 B.n609 163.367
R1855 B.n609 B.n608 163.367
R1856 B.n608 B.n105 163.367
R1857 B.n604 B.n105 163.367
R1858 B.n604 B.n603 163.367
R1859 B.n603 B.n602 163.367
R1860 B.n602 B.n107 163.367
R1861 B.n598 B.n107 163.367
R1862 B.n598 B.n597 163.367
R1863 B.n597 B.n596 163.367
R1864 B.n596 B.n109 163.367
R1865 B.n592 B.n109 163.367
R1866 B.n592 B.n591 163.367
R1867 B.n591 B.n590 163.367
R1868 B.n590 B.n111 163.367
R1869 B.n586 B.n111 163.367
R1870 B.n586 B.n585 163.367
R1871 B.n585 B.n584 163.367
R1872 B.n584 B.n113 163.367
R1873 B.n580 B.n113 163.367
R1874 B.n580 B.n579 163.367
R1875 B.n579 B.n578 163.367
R1876 B.n578 B.n115 163.367
R1877 B.n574 B.n115 163.367
R1878 B.n574 B.n573 163.367
R1879 B.n573 B.n572 163.367
R1880 B.n572 B.n117 163.367
R1881 B.n568 B.n117 163.367
R1882 B.n568 B.n567 163.367
R1883 B.n567 B.n566 163.367
R1884 B.n566 B.n119 163.367
R1885 B.n562 B.n119 163.367
R1886 B.n562 B.n561 163.367
R1887 B.n561 B.n560 163.367
R1888 B.n560 B.n121 163.367
R1889 B.n556 B.n121 163.367
R1890 B.n556 B.n555 163.367
R1891 B.n555 B.n554 163.367
R1892 B.n554 B.n123 163.367
R1893 B.n550 B.n123 163.367
R1894 B.n550 B.n549 163.367
R1895 B.n549 B.n548 163.367
R1896 B.n548 B.n125 163.367
R1897 B.n544 B.n125 163.367
R1898 B.n544 B.n543 163.367
R1899 B.n543 B.n542 163.367
R1900 B.n542 B.n127 163.367
R1901 B.n538 B.n127 163.367
R1902 B.n538 B.n537 163.367
R1903 B.n537 B.n536 163.367
R1904 B.n536 B.n129 163.367
R1905 B.n532 B.n129 163.367
R1906 B.n532 B.n531 163.367
R1907 B.n531 B.n530 163.367
R1908 B.n530 B.n131 163.367
R1909 B.n526 B.n131 163.367
R1910 B.n526 B.n525 163.367
R1911 B.n525 B.n524 163.367
R1912 B.n524 B.n133 163.367
R1913 B.n520 B.n133 163.367
R1914 B.n520 B.n519 163.367
R1915 B.n519 B.n518 163.367
R1916 B.n518 B.n135 163.367
R1917 B.n514 B.n135 163.367
R1918 B.n514 B.n513 163.367
R1919 B.n513 B.n512 163.367
R1920 B.n512 B.n137 163.367
R1921 B.n508 B.n137 163.367
R1922 B.n508 B.n507 163.367
R1923 B.n507 B.n506 163.367
R1924 B.n506 B.n139 163.367
R1925 B.n502 B.n139 163.367
R1926 B.n502 B.n501 163.367
R1927 B.n501 B.n500 163.367
R1928 B.n500 B.n141 163.367
R1929 B.n496 B.n141 163.367
R1930 B.n496 B.n495 163.367
R1931 B.n495 B.n494 163.367
R1932 B.n494 B.n143 163.367
R1933 B.n490 B.n143 163.367
R1934 B.n490 B.n489 163.367
R1935 B.n489 B.n488 163.367
R1936 B.n488 B.n145 163.367
R1937 B.n484 B.n145 163.367
R1938 B.n484 B.n483 163.367
R1939 B.n819 B.n818 163.367
R1940 B.n818 B.n31 163.367
R1941 B.n814 B.n31 163.367
R1942 B.n814 B.n813 163.367
R1943 B.n813 B.n812 163.367
R1944 B.n812 B.n33 163.367
R1945 B.n808 B.n33 163.367
R1946 B.n808 B.n807 163.367
R1947 B.n807 B.n806 163.367
R1948 B.n806 B.n35 163.367
R1949 B.n802 B.n35 163.367
R1950 B.n802 B.n801 163.367
R1951 B.n801 B.n800 163.367
R1952 B.n800 B.n37 163.367
R1953 B.n796 B.n37 163.367
R1954 B.n796 B.n795 163.367
R1955 B.n795 B.n794 163.367
R1956 B.n794 B.n39 163.367
R1957 B.n790 B.n39 163.367
R1958 B.n790 B.n789 163.367
R1959 B.n789 B.n788 163.367
R1960 B.n788 B.n41 163.367
R1961 B.n784 B.n41 163.367
R1962 B.n784 B.n783 163.367
R1963 B.n783 B.n782 163.367
R1964 B.n782 B.n43 163.367
R1965 B.n778 B.n43 163.367
R1966 B.n778 B.n777 163.367
R1967 B.n777 B.n776 163.367
R1968 B.n776 B.n45 163.367
R1969 B.n772 B.n45 163.367
R1970 B.n772 B.n771 163.367
R1971 B.n771 B.n770 163.367
R1972 B.n770 B.n47 163.367
R1973 B.n766 B.n47 163.367
R1974 B.n766 B.n765 163.367
R1975 B.n765 B.n764 163.367
R1976 B.n764 B.n49 163.367
R1977 B.n760 B.n49 163.367
R1978 B.n760 B.n759 163.367
R1979 B.n759 B.n758 163.367
R1980 B.n758 B.n51 163.367
R1981 B.n754 B.n51 163.367
R1982 B.n754 B.n753 163.367
R1983 B.n753 B.n752 163.367
R1984 B.n752 B.n53 163.367
R1985 B.n748 B.n53 163.367
R1986 B.n748 B.n747 163.367
R1987 B.n747 B.n746 163.367
R1988 B.n746 B.n55 163.367
R1989 B.n741 B.n55 163.367
R1990 B.n741 B.n740 163.367
R1991 B.n740 B.n739 163.367
R1992 B.n739 B.n59 163.367
R1993 B.n735 B.n59 163.367
R1994 B.n735 B.n734 163.367
R1995 B.n734 B.n733 163.367
R1996 B.n733 B.n61 163.367
R1997 B.n729 B.n61 163.367
R1998 B.n729 B.n728 163.367
R1999 B.n728 B.n65 163.367
R2000 B.n724 B.n65 163.367
R2001 B.n724 B.n723 163.367
R2002 B.n723 B.n722 163.367
R2003 B.n722 B.n67 163.367
R2004 B.n718 B.n67 163.367
R2005 B.n718 B.n717 163.367
R2006 B.n717 B.n716 163.367
R2007 B.n716 B.n69 163.367
R2008 B.n712 B.n69 163.367
R2009 B.n712 B.n711 163.367
R2010 B.n711 B.n710 163.367
R2011 B.n710 B.n71 163.367
R2012 B.n706 B.n71 163.367
R2013 B.n706 B.n705 163.367
R2014 B.n705 B.n704 163.367
R2015 B.n704 B.n73 163.367
R2016 B.n700 B.n73 163.367
R2017 B.n700 B.n699 163.367
R2018 B.n699 B.n698 163.367
R2019 B.n698 B.n75 163.367
R2020 B.n694 B.n75 163.367
R2021 B.n694 B.n693 163.367
R2022 B.n693 B.n692 163.367
R2023 B.n692 B.n77 163.367
R2024 B.n688 B.n77 163.367
R2025 B.n688 B.n687 163.367
R2026 B.n687 B.n686 163.367
R2027 B.n686 B.n79 163.367
R2028 B.n682 B.n79 163.367
R2029 B.n682 B.n681 163.367
R2030 B.n681 B.n680 163.367
R2031 B.n680 B.n81 163.367
R2032 B.n676 B.n81 163.367
R2033 B.n676 B.n675 163.367
R2034 B.n675 B.n674 163.367
R2035 B.n674 B.n83 163.367
R2036 B.n670 B.n83 163.367
R2037 B.n670 B.n669 163.367
R2038 B.n669 B.n668 163.367
R2039 B.n668 B.n85 163.367
R2040 B.n664 B.n85 163.367
R2041 B.n664 B.n663 163.367
R2042 B.n663 B.n662 163.367
R2043 B.n662 B.n87 163.367
R2044 B.n658 B.n87 163.367
R2045 B.n658 B.n657 163.367
R2046 B.n657 B.n656 163.367
R2047 B.n656 B.n89 163.367
R2048 B.n820 B.n29 163.367
R2049 B.n824 B.n29 163.367
R2050 B.n825 B.n824 163.367
R2051 B.n826 B.n825 163.367
R2052 B.n826 B.n27 163.367
R2053 B.n830 B.n27 163.367
R2054 B.n831 B.n830 163.367
R2055 B.n832 B.n831 163.367
R2056 B.n832 B.n25 163.367
R2057 B.n836 B.n25 163.367
R2058 B.n837 B.n836 163.367
R2059 B.n838 B.n837 163.367
R2060 B.n838 B.n23 163.367
R2061 B.n842 B.n23 163.367
R2062 B.n843 B.n842 163.367
R2063 B.n844 B.n843 163.367
R2064 B.n844 B.n21 163.367
R2065 B.n848 B.n21 163.367
R2066 B.n849 B.n848 163.367
R2067 B.n850 B.n849 163.367
R2068 B.n850 B.n19 163.367
R2069 B.n854 B.n19 163.367
R2070 B.n855 B.n854 163.367
R2071 B.n856 B.n855 163.367
R2072 B.n856 B.n17 163.367
R2073 B.n860 B.n17 163.367
R2074 B.n861 B.n860 163.367
R2075 B.n862 B.n861 163.367
R2076 B.n862 B.n15 163.367
R2077 B.n866 B.n15 163.367
R2078 B.n867 B.n866 163.367
R2079 B.n868 B.n867 163.367
R2080 B.n868 B.n13 163.367
R2081 B.n872 B.n13 163.367
R2082 B.n873 B.n872 163.367
R2083 B.n874 B.n873 163.367
R2084 B.n874 B.n11 163.367
R2085 B.n878 B.n11 163.367
R2086 B.n879 B.n878 163.367
R2087 B.n880 B.n879 163.367
R2088 B.n880 B.n9 163.367
R2089 B.n884 B.n9 163.367
R2090 B.n885 B.n884 163.367
R2091 B.n886 B.n885 163.367
R2092 B.n886 B.n7 163.367
R2093 B.n890 B.n7 163.367
R2094 B.n891 B.n890 163.367
R2095 B.n892 B.n891 163.367
R2096 B.n892 B.n5 163.367
R2097 B.n896 B.n5 163.367
R2098 B.n897 B.n896 163.367
R2099 B.n898 B.n897 163.367
R2100 B.n898 B.n3 163.367
R2101 B.n902 B.n3 163.367
R2102 B.n903 B.n902 163.367
R2103 B.n232 B.n2 163.367
R2104 B.n233 B.n232 163.367
R2105 B.n234 B.n233 163.367
R2106 B.n234 B.n229 163.367
R2107 B.n238 B.n229 163.367
R2108 B.n239 B.n238 163.367
R2109 B.n240 B.n239 163.367
R2110 B.n240 B.n227 163.367
R2111 B.n244 B.n227 163.367
R2112 B.n245 B.n244 163.367
R2113 B.n246 B.n245 163.367
R2114 B.n246 B.n225 163.367
R2115 B.n250 B.n225 163.367
R2116 B.n251 B.n250 163.367
R2117 B.n252 B.n251 163.367
R2118 B.n252 B.n223 163.367
R2119 B.n256 B.n223 163.367
R2120 B.n257 B.n256 163.367
R2121 B.n258 B.n257 163.367
R2122 B.n258 B.n221 163.367
R2123 B.n262 B.n221 163.367
R2124 B.n263 B.n262 163.367
R2125 B.n264 B.n263 163.367
R2126 B.n264 B.n219 163.367
R2127 B.n268 B.n219 163.367
R2128 B.n269 B.n268 163.367
R2129 B.n270 B.n269 163.367
R2130 B.n270 B.n217 163.367
R2131 B.n274 B.n217 163.367
R2132 B.n275 B.n274 163.367
R2133 B.n276 B.n275 163.367
R2134 B.n276 B.n215 163.367
R2135 B.n280 B.n215 163.367
R2136 B.n281 B.n280 163.367
R2137 B.n282 B.n281 163.367
R2138 B.n282 B.n213 163.367
R2139 B.n286 B.n213 163.367
R2140 B.n287 B.n286 163.367
R2141 B.n288 B.n287 163.367
R2142 B.n288 B.n211 163.367
R2143 B.n292 B.n211 163.367
R2144 B.n293 B.n292 163.367
R2145 B.n294 B.n293 163.367
R2146 B.n294 B.n209 163.367
R2147 B.n298 B.n209 163.367
R2148 B.n299 B.n298 163.367
R2149 B.n300 B.n299 163.367
R2150 B.n300 B.n207 163.367
R2151 B.n304 B.n207 163.367
R2152 B.n305 B.n304 163.367
R2153 B.n306 B.n305 163.367
R2154 B.n306 B.n205 163.367
R2155 B.n310 B.n205 163.367
R2156 B.n311 B.n310 163.367
R2157 B.n312 B.n311 163.367
R2158 B.n388 B.n387 63.8066
R2159 B.n173 B.n172 63.8066
R2160 B.n63 B.n62 63.8066
R2161 B.n57 B.n56 63.8066
R2162 B.n389 B.n388 59.5399
R2163 B.n407 B.n173 59.5399
R2164 B.n64 B.n63 59.5399
R2165 B.n744 B.n57 59.5399
R2166 B.n821 B.n30 32.3127
R2167 B.n654 B.n653 32.3127
R2168 B.n481 B.n146 32.3127
R2169 B.n314 B.n313 32.3127
R2170 B B.n905 18.0485
R2171 B.n822 B.n821 10.6151
R2172 B.n823 B.n822 10.6151
R2173 B.n823 B.n28 10.6151
R2174 B.n827 B.n28 10.6151
R2175 B.n828 B.n827 10.6151
R2176 B.n829 B.n828 10.6151
R2177 B.n829 B.n26 10.6151
R2178 B.n833 B.n26 10.6151
R2179 B.n834 B.n833 10.6151
R2180 B.n835 B.n834 10.6151
R2181 B.n835 B.n24 10.6151
R2182 B.n839 B.n24 10.6151
R2183 B.n840 B.n839 10.6151
R2184 B.n841 B.n840 10.6151
R2185 B.n841 B.n22 10.6151
R2186 B.n845 B.n22 10.6151
R2187 B.n846 B.n845 10.6151
R2188 B.n847 B.n846 10.6151
R2189 B.n847 B.n20 10.6151
R2190 B.n851 B.n20 10.6151
R2191 B.n852 B.n851 10.6151
R2192 B.n853 B.n852 10.6151
R2193 B.n853 B.n18 10.6151
R2194 B.n857 B.n18 10.6151
R2195 B.n858 B.n857 10.6151
R2196 B.n859 B.n858 10.6151
R2197 B.n859 B.n16 10.6151
R2198 B.n863 B.n16 10.6151
R2199 B.n864 B.n863 10.6151
R2200 B.n865 B.n864 10.6151
R2201 B.n865 B.n14 10.6151
R2202 B.n869 B.n14 10.6151
R2203 B.n870 B.n869 10.6151
R2204 B.n871 B.n870 10.6151
R2205 B.n871 B.n12 10.6151
R2206 B.n875 B.n12 10.6151
R2207 B.n876 B.n875 10.6151
R2208 B.n877 B.n876 10.6151
R2209 B.n877 B.n10 10.6151
R2210 B.n881 B.n10 10.6151
R2211 B.n882 B.n881 10.6151
R2212 B.n883 B.n882 10.6151
R2213 B.n883 B.n8 10.6151
R2214 B.n887 B.n8 10.6151
R2215 B.n888 B.n887 10.6151
R2216 B.n889 B.n888 10.6151
R2217 B.n889 B.n6 10.6151
R2218 B.n893 B.n6 10.6151
R2219 B.n894 B.n893 10.6151
R2220 B.n895 B.n894 10.6151
R2221 B.n895 B.n4 10.6151
R2222 B.n899 B.n4 10.6151
R2223 B.n900 B.n899 10.6151
R2224 B.n901 B.n900 10.6151
R2225 B.n901 B.n0 10.6151
R2226 B.n817 B.n30 10.6151
R2227 B.n817 B.n816 10.6151
R2228 B.n816 B.n815 10.6151
R2229 B.n815 B.n32 10.6151
R2230 B.n811 B.n32 10.6151
R2231 B.n811 B.n810 10.6151
R2232 B.n810 B.n809 10.6151
R2233 B.n809 B.n34 10.6151
R2234 B.n805 B.n34 10.6151
R2235 B.n805 B.n804 10.6151
R2236 B.n804 B.n803 10.6151
R2237 B.n803 B.n36 10.6151
R2238 B.n799 B.n36 10.6151
R2239 B.n799 B.n798 10.6151
R2240 B.n798 B.n797 10.6151
R2241 B.n797 B.n38 10.6151
R2242 B.n793 B.n38 10.6151
R2243 B.n793 B.n792 10.6151
R2244 B.n792 B.n791 10.6151
R2245 B.n791 B.n40 10.6151
R2246 B.n787 B.n40 10.6151
R2247 B.n787 B.n786 10.6151
R2248 B.n786 B.n785 10.6151
R2249 B.n785 B.n42 10.6151
R2250 B.n781 B.n42 10.6151
R2251 B.n781 B.n780 10.6151
R2252 B.n780 B.n779 10.6151
R2253 B.n779 B.n44 10.6151
R2254 B.n775 B.n44 10.6151
R2255 B.n775 B.n774 10.6151
R2256 B.n774 B.n773 10.6151
R2257 B.n773 B.n46 10.6151
R2258 B.n769 B.n46 10.6151
R2259 B.n769 B.n768 10.6151
R2260 B.n768 B.n767 10.6151
R2261 B.n767 B.n48 10.6151
R2262 B.n763 B.n48 10.6151
R2263 B.n763 B.n762 10.6151
R2264 B.n762 B.n761 10.6151
R2265 B.n761 B.n50 10.6151
R2266 B.n757 B.n50 10.6151
R2267 B.n757 B.n756 10.6151
R2268 B.n756 B.n755 10.6151
R2269 B.n755 B.n52 10.6151
R2270 B.n751 B.n52 10.6151
R2271 B.n751 B.n750 10.6151
R2272 B.n750 B.n749 10.6151
R2273 B.n749 B.n54 10.6151
R2274 B.n745 B.n54 10.6151
R2275 B.n743 B.n742 10.6151
R2276 B.n742 B.n58 10.6151
R2277 B.n738 B.n58 10.6151
R2278 B.n738 B.n737 10.6151
R2279 B.n737 B.n736 10.6151
R2280 B.n736 B.n60 10.6151
R2281 B.n732 B.n60 10.6151
R2282 B.n732 B.n731 10.6151
R2283 B.n731 B.n730 10.6151
R2284 B.n727 B.n726 10.6151
R2285 B.n726 B.n725 10.6151
R2286 B.n725 B.n66 10.6151
R2287 B.n721 B.n66 10.6151
R2288 B.n721 B.n720 10.6151
R2289 B.n720 B.n719 10.6151
R2290 B.n719 B.n68 10.6151
R2291 B.n715 B.n68 10.6151
R2292 B.n715 B.n714 10.6151
R2293 B.n714 B.n713 10.6151
R2294 B.n713 B.n70 10.6151
R2295 B.n709 B.n70 10.6151
R2296 B.n709 B.n708 10.6151
R2297 B.n708 B.n707 10.6151
R2298 B.n707 B.n72 10.6151
R2299 B.n703 B.n72 10.6151
R2300 B.n703 B.n702 10.6151
R2301 B.n702 B.n701 10.6151
R2302 B.n701 B.n74 10.6151
R2303 B.n697 B.n74 10.6151
R2304 B.n697 B.n696 10.6151
R2305 B.n696 B.n695 10.6151
R2306 B.n695 B.n76 10.6151
R2307 B.n691 B.n76 10.6151
R2308 B.n691 B.n690 10.6151
R2309 B.n690 B.n689 10.6151
R2310 B.n689 B.n78 10.6151
R2311 B.n685 B.n78 10.6151
R2312 B.n685 B.n684 10.6151
R2313 B.n684 B.n683 10.6151
R2314 B.n683 B.n80 10.6151
R2315 B.n679 B.n80 10.6151
R2316 B.n679 B.n678 10.6151
R2317 B.n678 B.n677 10.6151
R2318 B.n677 B.n82 10.6151
R2319 B.n673 B.n82 10.6151
R2320 B.n673 B.n672 10.6151
R2321 B.n672 B.n671 10.6151
R2322 B.n671 B.n84 10.6151
R2323 B.n667 B.n84 10.6151
R2324 B.n667 B.n666 10.6151
R2325 B.n666 B.n665 10.6151
R2326 B.n665 B.n86 10.6151
R2327 B.n661 B.n86 10.6151
R2328 B.n661 B.n660 10.6151
R2329 B.n660 B.n659 10.6151
R2330 B.n659 B.n88 10.6151
R2331 B.n655 B.n88 10.6151
R2332 B.n655 B.n654 10.6151
R2333 B.n653 B.n90 10.6151
R2334 B.n649 B.n90 10.6151
R2335 B.n649 B.n648 10.6151
R2336 B.n648 B.n647 10.6151
R2337 B.n647 B.n92 10.6151
R2338 B.n643 B.n92 10.6151
R2339 B.n643 B.n642 10.6151
R2340 B.n642 B.n641 10.6151
R2341 B.n641 B.n94 10.6151
R2342 B.n637 B.n94 10.6151
R2343 B.n637 B.n636 10.6151
R2344 B.n636 B.n635 10.6151
R2345 B.n635 B.n96 10.6151
R2346 B.n631 B.n96 10.6151
R2347 B.n631 B.n630 10.6151
R2348 B.n630 B.n629 10.6151
R2349 B.n629 B.n98 10.6151
R2350 B.n625 B.n98 10.6151
R2351 B.n625 B.n624 10.6151
R2352 B.n624 B.n623 10.6151
R2353 B.n623 B.n100 10.6151
R2354 B.n619 B.n100 10.6151
R2355 B.n619 B.n618 10.6151
R2356 B.n618 B.n617 10.6151
R2357 B.n617 B.n102 10.6151
R2358 B.n613 B.n102 10.6151
R2359 B.n613 B.n612 10.6151
R2360 B.n612 B.n611 10.6151
R2361 B.n611 B.n104 10.6151
R2362 B.n607 B.n104 10.6151
R2363 B.n607 B.n606 10.6151
R2364 B.n606 B.n605 10.6151
R2365 B.n605 B.n106 10.6151
R2366 B.n601 B.n106 10.6151
R2367 B.n601 B.n600 10.6151
R2368 B.n600 B.n599 10.6151
R2369 B.n599 B.n108 10.6151
R2370 B.n595 B.n108 10.6151
R2371 B.n595 B.n594 10.6151
R2372 B.n594 B.n593 10.6151
R2373 B.n593 B.n110 10.6151
R2374 B.n589 B.n110 10.6151
R2375 B.n589 B.n588 10.6151
R2376 B.n588 B.n587 10.6151
R2377 B.n587 B.n112 10.6151
R2378 B.n583 B.n112 10.6151
R2379 B.n583 B.n582 10.6151
R2380 B.n582 B.n581 10.6151
R2381 B.n581 B.n114 10.6151
R2382 B.n577 B.n114 10.6151
R2383 B.n577 B.n576 10.6151
R2384 B.n576 B.n575 10.6151
R2385 B.n575 B.n116 10.6151
R2386 B.n571 B.n116 10.6151
R2387 B.n571 B.n570 10.6151
R2388 B.n570 B.n569 10.6151
R2389 B.n569 B.n118 10.6151
R2390 B.n565 B.n118 10.6151
R2391 B.n565 B.n564 10.6151
R2392 B.n564 B.n563 10.6151
R2393 B.n563 B.n120 10.6151
R2394 B.n559 B.n120 10.6151
R2395 B.n559 B.n558 10.6151
R2396 B.n558 B.n557 10.6151
R2397 B.n557 B.n122 10.6151
R2398 B.n553 B.n122 10.6151
R2399 B.n553 B.n552 10.6151
R2400 B.n552 B.n551 10.6151
R2401 B.n551 B.n124 10.6151
R2402 B.n547 B.n124 10.6151
R2403 B.n547 B.n546 10.6151
R2404 B.n546 B.n545 10.6151
R2405 B.n545 B.n126 10.6151
R2406 B.n541 B.n126 10.6151
R2407 B.n541 B.n540 10.6151
R2408 B.n540 B.n539 10.6151
R2409 B.n539 B.n128 10.6151
R2410 B.n535 B.n128 10.6151
R2411 B.n535 B.n534 10.6151
R2412 B.n534 B.n533 10.6151
R2413 B.n533 B.n130 10.6151
R2414 B.n529 B.n130 10.6151
R2415 B.n529 B.n528 10.6151
R2416 B.n528 B.n527 10.6151
R2417 B.n527 B.n132 10.6151
R2418 B.n523 B.n132 10.6151
R2419 B.n523 B.n522 10.6151
R2420 B.n522 B.n521 10.6151
R2421 B.n521 B.n134 10.6151
R2422 B.n517 B.n134 10.6151
R2423 B.n517 B.n516 10.6151
R2424 B.n516 B.n515 10.6151
R2425 B.n515 B.n136 10.6151
R2426 B.n511 B.n136 10.6151
R2427 B.n511 B.n510 10.6151
R2428 B.n510 B.n509 10.6151
R2429 B.n509 B.n138 10.6151
R2430 B.n505 B.n138 10.6151
R2431 B.n505 B.n504 10.6151
R2432 B.n504 B.n503 10.6151
R2433 B.n503 B.n140 10.6151
R2434 B.n499 B.n140 10.6151
R2435 B.n499 B.n498 10.6151
R2436 B.n498 B.n497 10.6151
R2437 B.n497 B.n142 10.6151
R2438 B.n493 B.n142 10.6151
R2439 B.n493 B.n492 10.6151
R2440 B.n492 B.n491 10.6151
R2441 B.n491 B.n144 10.6151
R2442 B.n487 B.n144 10.6151
R2443 B.n487 B.n486 10.6151
R2444 B.n486 B.n485 10.6151
R2445 B.n485 B.n146 10.6151
R2446 B.n231 B.n1 10.6151
R2447 B.n231 B.n230 10.6151
R2448 B.n235 B.n230 10.6151
R2449 B.n236 B.n235 10.6151
R2450 B.n237 B.n236 10.6151
R2451 B.n237 B.n228 10.6151
R2452 B.n241 B.n228 10.6151
R2453 B.n242 B.n241 10.6151
R2454 B.n243 B.n242 10.6151
R2455 B.n243 B.n226 10.6151
R2456 B.n247 B.n226 10.6151
R2457 B.n248 B.n247 10.6151
R2458 B.n249 B.n248 10.6151
R2459 B.n249 B.n224 10.6151
R2460 B.n253 B.n224 10.6151
R2461 B.n254 B.n253 10.6151
R2462 B.n255 B.n254 10.6151
R2463 B.n255 B.n222 10.6151
R2464 B.n259 B.n222 10.6151
R2465 B.n260 B.n259 10.6151
R2466 B.n261 B.n260 10.6151
R2467 B.n261 B.n220 10.6151
R2468 B.n265 B.n220 10.6151
R2469 B.n266 B.n265 10.6151
R2470 B.n267 B.n266 10.6151
R2471 B.n267 B.n218 10.6151
R2472 B.n271 B.n218 10.6151
R2473 B.n272 B.n271 10.6151
R2474 B.n273 B.n272 10.6151
R2475 B.n273 B.n216 10.6151
R2476 B.n277 B.n216 10.6151
R2477 B.n278 B.n277 10.6151
R2478 B.n279 B.n278 10.6151
R2479 B.n279 B.n214 10.6151
R2480 B.n283 B.n214 10.6151
R2481 B.n284 B.n283 10.6151
R2482 B.n285 B.n284 10.6151
R2483 B.n285 B.n212 10.6151
R2484 B.n289 B.n212 10.6151
R2485 B.n290 B.n289 10.6151
R2486 B.n291 B.n290 10.6151
R2487 B.n291 B.n210 10.6151
R2488 B.n295 B.n210 10.6151
R2489 B.n296 B.n295 10.6151
R2490 B.n297 B.n296 10.6151
R2491 B.n297 B.n208 10.6151
R2492 B.n301 B.n208 10.6151
R2493 B.n302 B.n301 10.6151
R2494 B.n303 B.n302 10.6151
R2495 B.n303 B.n206 10.6151
R2496 B.n307 B.n206 10.6151
R2497 B.n308 B.n307 10.6151
R2498 B.n309 B.n308 10.6151
R2499 B.n309 B.n204 10.6151
R2500 B.n313 B.n204 10.6151
R2501 B.n315 B.n314 10.6151
R2502 B.n315 B.n202 10.6151
R2503 B.n319 B.n202 10.6151
R2504 B.n320 B.n319 10.6151
R2505 B.n321 B.n320 10.6151
R2506 B.n321 B.n200 10.6151
R2507 B.n325 B.n200 10.6151
R2508 B.n326 B.n325 10.6151
R2509 B.n327 B.n326 10.6151
R2510 B.n327 B.n198 10.6151
R2511 B.n331 B.n198 10.6151
R2512 B.n332 B.n331 10.6151
R2513 B.n333 B.n332 10.6151
R2514 B.n333 B.n196 10.6151
R2515 B.n337 B.n196 10.6151
R2516 B.n338 B.n337 10.6151
R2517 B.n339 B.n338 10.6151
R2518 B.n339 B.n194 10.6151
R2519 B.n343 B.n194 10.6151
R2520 B.n344 B.n343 10.6151
R2521 B.n345 B.n344 10.6151
R2522 B.n345 B.n192 10.6151
R2523 B.n349 B.n192 10.6151
R2524 B.n350 B.n349 10.6151
R2525 B.n351 B.n350 10.6151
R2526 B.n351 B.n190 10.6151
R2527 B.n355 B.n190 10.6151
R2528 B.n356 B.n355 10.6151
R2529 B.n357 B.n356 10.6151
R2530 B.n357 B.n188 10.6151
R2531 B.n361 B.n188 10.6151
R2532 B.n362 B.n361 10.6151
R2533 B.n363 B.n362 10.6151
R2534 B.n363 B.n186 10.6151
R2535 B.n367 B.n186 10.6151
R2536 B.n368 B.n367 10.6151
R2537 B.n369 B.n368 10.6151
R2538 B.n369 B.n184 10.6151
R2539 B.n373 B.n184 10.6151
R2540 B.n374 B.n373 10.6151
R2541 B.n375 B.n374 10.6151
R2542 B.n375 B.n182 10.6151
R2543 B.n379 B.n182 10.6151
R2544 B.n380 B.n379 10.6151
R2545 B.n381 B.n380 10.6151
R2546 B.n381 B.n180 10.6151
R2547 B.n385 B.n180 10.6151
R2548 B.n386 B.n385 10.6151
R2549 B.n390 B.n386 10.6151
R2550 B.n394 B.n178 10.6151
R2551 B.n395 B.n394 10.6151
R2552 B.n396 B.n395 10.6151
R2553 B.n396 B.n176 10.6151
R2554 B.n400 B.n176 10.6151
R2555 B.n401 B.n400 10.6151
R2556 B.n402 B.n401 10.6151
R2557 B.n402 B.n174 10.6151
R2558 B.n406 B.n174 10.6151
R2559 B.n409 B.n408 10.6151
R2560 B.n409 B.n170 10.6151
R2561 B.n413 B.n170 10.6151
R2562 B.n414 B.n413 10.6151
R2563 B.n415 B.n414 10.6151
R2564 B.n415 B.n168 10.6151
R2565 B.n419 B.n168 10.6151
R2566 B.n420 B.n419 10.6151
R2567 B.n421 B.n420 10.6151
R2568 B.n421 B.n166 10.6151
R2569 B.n425 B.n166 10.6151
R2570 B.n426 B.n425 10.6151
R2571 B.n427 B.n426 10.6151
R2572 B.n427 B.n164 10.6151
R2573 B.n431 B.n164 10.6151
R2574 B.n432 B.n431 10.6151
R2575 B.n433 B.n432 10.6151
R2576 B.n433 B.n162 10.6151
R2577 B.n437 B.n162 10.6151
R2578 B.n438 B.n437 10.6151
R2579 B.n439 B.n438 10.6151
R2580 B.n439 B.n160 10.6151
R2581 B.n443 B.n160 10.6151
R2582 B.n444 B.n443 10.6151
R2583 B.n445 B.n444 10.6151
R2584 B.n445 B.n158 10.6151
R2585 B.n449 B.n158 10.6151
R2586 B.n450 B.n449 10.6151
R2587 B.n451 B.n450 10.6151
R2588 B.n451 B.n156 10.6151
R2589 B.n455 B.n156 10.6151
R2590 B.n456 B.n455 10.6151
R2591 B.n457 B.n456 10.6151
R2592 B.n457 B.n154 10.6151
R2593 B.n461 B.n154 10.6151
R2594 B.n462 B.n461 10.6151
R2595 B.n463 B.n462 10.6151
R2596 B.n463 B.n152 10.6151
R2597 B.n467 B.n152 10.6151
R2598 B.n468 B.n467 10.6151
R2599 B.n469 B.n468 10.6151
R2600 B.n469 B.n150 10.6151
R2601 B.n473 B.n150 10.6151
R2602 B.n474 B.n473 10.6151
R2603 B.n475 B.n474 10.6151
R2604 B.n475 B.n148 10.6151
R2605 B.n479 B.n148 10.6151
R2606 B.n480 B.n479 10.6151
R2607 B.n481 B.n480 10.6151
R2608 B.n745 B.n744 9.36635
R2609 B.n727 B.n64 9.36635
R2610 B.n390 B.n389 9.36635
R2611 B.n408 B.n407 9.36635
R2612 B.n905 B.n0 8.11757
R2613 B.n905 B.n1 8.11757
R2614 B.n744 B.n743 1.24928
R2615 B.n730 B.n64 1.24928
R2616 B.n389 B.n178 1.24928
R2617 B.n407 B.n406 1.24928
C0 VTAIL VDD1 9.094019f
C1 VDD1 VN 0.15283f
C2 VTAIL VP 11.366599f
C3 w_n4260_n3952# VTAIL 4.88181f
C4 VP VN 8.639171f
C5 w_n4260_n3952# VN 8.8173f
C6 VTAIL VDD2 9.150849f
C7 VDD2 VN 10.9563f
C8 VDD1 VP 11.3603f
C9 w_n4260_n3952# VDD1 2.15189f
C10 w_n4260_n3952# VP 9.371401f
C11 B VTAIL 6.11902f
C12 VDD1 VDD2 1.96574f
C13 B VN 1.34735f
C14 VDD2 VP 0.55843f
C15 w_n4260_n3952# VDD2 2.2817f
C16 B VDD1 1.83723f
C17 B VP 2.27813f
C18 w_n4260_n3952# B 11.4856f
C19 B VDD2 1.94459f
C20 VTAIL VN 11.352401f
C21 VDD2 VSUBS 2.086501f
C22 VDD1 VSUBS 2.79446f
C23 VTAIL VSUBS 1.529521f
C24 VN VSUBS 7.32608f
C25 VP VSUBS 4.073168f
C26 B VSUBS 5.652764f
C27 w_n4260_n3952# VSUBS 0.206474p
C28 B.n0 VSUBS 0.006144f
C29 B.n1 VSUBS 0.006144f
C30 B.n2 VSUBS 0.009087f
C31 B.n3 VSUBS 0.006963f
C32 B.n4 VSUBS 0.006963f
C33 B.n5 VSUBS 0.006963f
C34 B.n6 VSUBS 0.006963f
C35 B.n7 VSUBS 0.006963f
C36 B.n8 VSUBS 0.006963f
C37 B.n9 VSUBS 0.006963f
C38 B.n10 VSUBS 0.006963f
C39 B.n11 VSUBS 0.006963f
C40 B.n12 VSUBS 0.006963f
C41 B.n13 VSUBS 0.006963f
C42 B.n14 VSUBS 0.006963f
C43 B.n15 VSUBS 0.006963f
C44 B.n16 VSUBS 0.006963f
C45 B.n17 VSUBS 0.006963f
C46 B.n18 VSUBS 0.006963f
C47 B.n19 VSUBS 0.006963f
C48 B.n20 VSUBS 0.006963f
C49 B.n21 VSUBS 0.006963f
C50 B.n22 VSUBS 0.006963f
C51 B.n23 VSUBS 0.006963f
C52 B.n24 VSUBS 0.006963f
C53 B.n25 VSUBS 0.006963f
C54 B.n26 VSUBS 0.006963f
C55 B.n27 VSUBS 0.006963f
C56 B.n28 VSUBS 0.006963f
C57 B.n29 VSUBS 0.006963f
C58 B.n30 VSUBS 0.016575f
C59 B.n31 VSUBS 0.006963f
C60 B.n32 VSUBS 0.006963f
C61 B.n33 VSUBS 0.006963f
C62 B.n34 VSUBS 0.006963f
C63 B.n35 VSUBS 0.006963f
C64 B.n36 VSUBS 0.006963f
C65 B.n37 VSUBS 0.006963f
C66 B.n38 VSUBS 0.006963f
C67 B.n39 VSUBS 0.006963f
C68 B.n40 VSUBS 0.006963f
C69 B.n41 VSUBS 0.006963f
C70 B.n42 VSUBS 0.006963f
C71 B.n43 VSUBS 0.006963f
C72 B.n44 VSUBS 0.006963f
C73 B.n45 VSUBS 0.006963f
C74 B.n46 VSUBS 0.006963f
C75 B.n47 VSUBS 0.006963f
C76 B.n48 VSUBS 0.006963f
C77 B.n49 VSUBS 0.006963f
C78 B.n50 VSUBS 0.006963f
C79 B.n51 VSUBS 0.006963f
C80 B.n52 VSUBS 0.006963f
C81 B.n53 VSUBS 0.006963f
C82 B.n54 VSUBS 0.006963f
C83 B.n55 VSUBS 0.006963f
C84 B.t4 VSUBS 0.276494f
C85 B.t5 VSUBS 0.312858f
C86 B.t3 VSUBS 1.9915f
C87 B.n56 VSUBS 0.491265f
C88 B.n57 VSUBS 0.290446f
C89 B.n58 VSUBS 0.006963f
C90 B.n59 VSUBS 0.006963f
C91 B.n60 VSUBS 0.006963f
C92 B.n61 VSUBS 0.006963f
C93 B.t10 VSUBS 0.276498f
C94 B.t11 VSUBS 0.312861f
C95 B.t9 VSUBS 1.9915f
C96 B.n62 VSUBS 0.491262f
C97 B.n63 VSUBS 0.290443f
C98 B.n64 VSUBS 0.016133f
C99 B.n65 VSUBS 0.006963f
C100 B.n66 VSUBS 0.006963f
C101 B.n67 VSUBS 0.006963f
C102 B.n68 VSUBS 0.006963f
C103 B.n69 VSUBS 0.006963f
C104 B.n70 VSUBS 0.006963f
C105 B.n71 VSUBS 0.006963f
C106 B.n72 VSUBS 0.006963f
C107 B.n73 VSUBS 0.006963f
C108 B.n74 VSUBS 0.006963f
C109 B.n75 VSUBS 0.006963f
C110 B.n76 VSUBS 0.006963f
C111 B.n77 VSUBS 0.006963f
C112 B.n78 VSUBS 0.006963f
C113 B.n79 VSUBS 0.006963f
C114 B.n80 VSUBS 0.006963f
C115 B.n81 VSUBS 0.006963f
C116 B.n82 VSUBS 0.006963f
C117 B.n83 VSUBS 0.006963f
C118 B.n84 VSUBS 0.006963f
C119 B.n85 VSUBS 0.006963f
C120 B.n86 VSUBS 0.006963f
C121 B.n87 VSUBS 0.006963f
C122 B.n88 VSUBS 0.006963f
C123 B.n89 VSUBS 0.016575f
C124 B.n90 VSUBS 0.006963f
C125 B.n91 VSUBS 0.006963f
C126 B.n92 VSUBS 0.006963f
C127 B.n93 VSUBS 0.006963f
C128 B.n94 VSUBS 0.006963f
C129 B.n95 VSUBS 0.006963f
C130 B.n96 VSUBS 0.006963f
C131 B.n97 VSUBS 0.006963f
C132 B.n98 VSUBS 0.006963f
C133 B.n99 VSUBS 0.006963f
C134 B.n100 VSUBS 0.006963f
C135 B.n101 VSUBS 0.006963f
C136 B.n102 VSUBS 0.006963f
C137 B.n103 VSUBS 0.006963f
C138 B.n104 VSUBS 0.006963f
C139 B.n105 VSUBS 0.006963f
C140 B.n106 VSUBS 0.006963f
C141 B.n107 VSUBS 0.006963f
C142 B.n108 VSUBS 0.006963f
C143 B.n109 VSUBS 0.006963f
C144 B.n110 VSUBS 0.006963f
C145 B.n111 VSUBS 0.006963f
C146 B.n112 VSUBS 0.006963f
C147 B.n113 VSUBS 0.006963f
C148 B.n114 VSUBS 0.006963f
C149 B.n115 VSUBS 0.006963f
C150 B.n116 VSUBS 0.006963f
C151 B.n117 VSUBS 0.006963f
C152 B.n118 VSUBS 0.006963f
C153 B.n119 VSUBS 0.006963f
C154 B.n120 VSUBS 0.006963f
C155 B.n121 VSUBS 0.006963f
C156 B.n122 VSUBS 0.006963f
C157 B.n123 VSUBS 0.006963f
C158 B.n124 VSUBS 0.006963f
C159 B.n125 VSUBS 0.006963f
C160 B.n126 VSUBS 0.006963f
C161 B.n127 VSUBS 0.006963f
C162 B.n128 VSUBS 0.006963f
C163 B.n129 VSUBS 0.006963f
C164 B.n130 VSUBS 0.006963f
C165 B.n131 VSUBS 0.006963f
C166 B.n132 VSUBS 0.006963f
C167 B.n133 VSUBS 0.006963f
C168 B.n134 VSUBS 0.006963f
C169 B.n135 VSUBS 0.006963f
C170 B.n136 VSUBS 0.006963f
C171 B.n137 VSUBS 0.006963f
C172 B.n138 VSUBS 0.006963f
C173 B.n139 VSUBS 0.006963f
C174 B.n140 VSUBS 0.006963f
C175 B.n141 VSUBS 0.006963f
C176 B.n142 VSUBS 0.006963f
C177 B.n143 VSUBS 0.006963f
C178 B.n144 VSUBS 0.006963f
C179 B.n145 VSUBS 0.006963f
C180 B.n146 VSUBS 0.016616f
C181 B.n147 VSUBS 0.006963f
C182 B.n148 VSUBS 0.006963f
C183 B.n149 VSUBS 0.006963f
C184 B.n150 VSUBS 0.006963f
C185 B.n151 VSUBS 0.006963f
C186 B.n152 VSUBS 0.006963f
C187 B.n153 VSUBS 0.006963f
C188 B.n154 VSUBS 0.006963f
C189 B.n155 VSUBS 0.006963f
C190 B.n156 VSUBS 0.006963f
C191 B.n157 VSUBS 0.006963f
C192 B.n158 VSUBS 0.006963f
C193 B.n159 VSUBS 0.006963f
C194 B.n160 VSUBS 0.006963f
C195 B.n161 VSUBS 0.006963f
C196 B.n162 VSUBS 0.006963f
C197 B.n163 VSUBS 0.006963f
C198 B.n164 VSUBS 0.006963f
C199 B.n165 VSUBS 0.006963f
C200 B.n166 VSUBS 0.006963f
C201 B.n167 VSUBS 0.006963f
C202 B.n168 VSUBS 0.006963f
C203 B.n169 VSUBS 0.006963f
C204 B.n170 VSUBS 0.006963f
C205 B.n171 VSUBS 0.006963f
C206 B.t8 VSUBS 0.276498f
C207 B.t7 VSUBS 0.312861f
C208 B.t6 VSUBS 1.9915f
C209 B.n172 VSUBS 0.491262f
C210 B.n173 VSUBS 0.290443f
C211 B.n174 VSUBS 0.006963f
C212 B.n175 VSUBS 0.006963f
C213 B.n176 VSUBS 0.006963f
C214 B.n177 VSUBS 0.006963f
C215 B.n178 VSUBS 0.003891f
C216 B.n179 VSUBS 0.006963f
C217 B.n180 VSUBS 0.006963f
C218 B.n181 VSUBS 0.006963f
C219 B.n182 VSUBS 0.006963f
C220 B.n183 VSUBS 0.006963f
C221 B.n184 VSUBS 0.006963f
C222 B.n185 VSUBS 0.006963f
C223 B.n186 VSUBS 0.006963f
C224 B.n187 VSUBS 0.006963f
C225 B.n188 VSUBS 0.006963f
C226 B.n189 VSUBS 0.006963f
C227 B.n190 VSUBS 0.006963f
C228 B.n191 VSUBS 0.006963f
C229 B.n192 VSUBS 0.006963f
C230 B.n193 VSUBS 0.006963f
C231 B.n194 VSUBS 0.006963f
C232 B.n195 VSUBS 0.006963f
C233 B.n196 VSUBS 0.006963f
C234 B.n197 VSUBS 0.006963f
C235 B.n198 VSUBS 0.006963f
C236 B.n199 VSUBS 0.006963f
C237 B.n200 VSUBS 0.006963f
C238 B.n201 VSUBS 0.006963f
C239 B.n202 VSUBS 0.006963f
C240 B.n203 VSUBS 0.016575f
C241 B.n204 VSUBS 0.006963f
C242 B.n205 VSUBS 0.006963f
C243 B.n206 VSUBS 0.006963f
C244 B.n207 VSUBS 0.006963f
C245 B.n208 VSUBS 0.006963f
C246 B.n209 VSUBS 0.006963f
C247 B.n210 VSUBS 0.006963f
C248 B.n211 VSUBS 0.006963f
C249 B.n212 VSUBS 0.006963f
C250 B.n213 VSUBS 0.006963f
C251 B.n214 VSUBS 0.006963f
C252 B.n215 VSUBS 0.006963f
C253 B.n216 VSUBS 0.006963f
C254 B.n217 VSUBS 0.006963f
C255 B.n218 VSUBS 0.006963f
C256 B.n219 VSUBS 0.006963f
C257 B.n220 VSUBS 0.006963f
C258 B.n221 VSUBS 0.006963f
C259 B.n222 VSUBS 0.006963f
C260 B.n223 VSUBS 0.006963f
C261 B.n224 VSUBS 0.006963f
C262 B.n225 VSUBS 0.006963f
C263 B.n226 VSUBS 0.006963f
C264 B.n227 VSUBS 0.006963f
C265 B.n228 VSUBS 0.006963f
C266 B.n229 VSUBS 0.006963f
C267 B.n230 VSUBS 0.006963f
C268 B.n231 VSUBS 0.006963f
C269 B.n232 VSUBS 0.006963f
C270 B.n233 VSUBS 0.006963f
C271 B.n234 VSUBS 0.006963f
C272 B.n235 VSUBS 0.006963f
C273 B.n236 VSUBS 0.006963f
C274 B.n237 VSUBS 0.006963f
C275 B.n238 VSUBS 0.006963f
C276 B.n239 VSUBS 0.006963f
C277 B.n240 VSUBS 0.006963f
C278 B.n241 VSUBS 0.006963f
C279 B.n242 VSUBS 0.006963f
C280 B.n243 VSUBS 0.006963f
C281 B.n244 VSUBS 0.006963f
C282 B.n245 VSUBS 0.006963f
C283 B.n246 VSUBS 0.006963f
C284 B.n247 VSUBS 0.006963f
C285 B.n248 VSUBS 0.006963f
C286 B.n249 VSUBS 0.006963f
C287 B.n250 VSUBS 0.006963f
C288 B.n251 VSUBS 0.006963f
C289 B.n252 VSUBS 0.006963f
C290 B.n253 VSUBS 0.006963f
C291 B.n254 VSUBS 0.006963f
C292 B.n255 VSUBS 0.006963f
C293 B.n256 VSUBS 0.006963f
C294 B.n257 VSUBS 0.006963f
C295 B.n258 VSUBS 0.006963f
C296 B.n259 VSUBS 0.006963f
C297 B.n260 VSUBS 0.006963f
C298 B.n261 VSUBS 0.006963f
C299 B.n262 VSUBS 0.006963f
C300 B.n263 VSUBS 0.006963f
C301 B.n264 VSUBS 0.006963f
C302 B.n265 VSUBS 0.006963f
C303 B.n266 VSUBS 0.006963f
C304 B.n267 VSUBS 0.006963f
C305 B.n268 VSUBS 0.006963f
C306 B.n269 VSUBS 0.006963f
C307 B.n270 VSUBS 0.006963f
C308 B.n271 VSUBS 0.006963f
C309 B.n272 VSUBS 0.006963f
C310 B.n273 VSUBS 0.006963f
C311 B.n274 VSUBS 0.006963f
C312 B.n275 VSUBS 0.006963f
C313 B.n276 VSUBS 0.006963f
C314 B.n277 VSUBS 0.006963f
C315 B.n278 VSUBS 0.006963f
C316 B.n279 VSUBS 0.006963f
C317 B.n280 VSUBS 0.006963f
C318 B.n281 VSUBS 0.006963f
C319 B.n282 VSUBS 0.006963f
C320 B.n283 VSUBS 0.006963f
C321 B.n284 VSUBS 0.006963f
C322 B.n285 VSUBS 0.006963f
C323 B.n286 VSUBS 0.006963f
C324 B.n287 VSUBS 0.006963f
C325 B.n288 VSUBS 0.006963f
C326 B.n289 VSUBS 0.006963f
C327 B.n290 VSUBS 0.006963f
C328 B.n291 VSUBS 0.006963f
C329 B.n292 VSUBS 0.006963f
C330 B.n293 VSUBS 0.006963f
C331 B.n294 VSUBS 0.006963f
C332 B.n295 VSUBS 0.006963f
C333 B.n296 VSUBS 0.006963f
C334 B.n297 VSUBS 0.006963f
C335 B.n298 VSUBS 0.006963f
C336 B.n299 VSUBS 0.006963f
C337 B.n300 VSUBS 0.006963f
C338 B.n301 VSUBS 0.006963f
C339 B.n302 VSUBS 0.006963f
C340 B.n303 VSUBS 0.006963f
C341 B.n304 VSUBS 0.006963f
C342 B.n305 VSUBS 0.006963f
C343 B.n306 VSUBS 0.006963f
C344 B.n307 VSUBS 0.006963f
C345 B.n308 VSUBS 0.006963f
C346 B.n309 VSUBS 0.006963f
C347 B.n310 VSUBS 0.006963f
C348 B.n311 VSUBS 0.006963f
C349 B.n312 VSUBS 0.015784f
C350 B.n313 VSUBS 0.015784f
C351 B.n314 VSUBS 0.016575f
C352 B.n315 VSUBS 0.006963f
C353 B.n316 VSUBS 0.006963f
C354 B.n317 VSUBS 0.006963f
C355 B.n318 VSUBS 0.006963f
C356 B.n319 VSUBS 0.006963f
C357 B.n320 VSUBS 0.006963f
C358 B.n321 VSUBS 0.006963f
C359 B.n322 VSUBS 0.006963f
C360 B.n323 VSUBS 0.006963f
C361 B.n324 VSUBS 0.006963f
C362 B.n325 VSUBS 0.006963f
C363 B.n326 VSUBS 0.006963f
C364 B.n327 VSUBS 0.006963f
C365 B.n328 VSUBS 0.006963f
C366 B.n329 VSUBS 0.006963f
C367 B.n330 VSUBS 0.006963f
C368 B.n331 VSUBS 0.006963f
C369 B.n332 VSUBS 0.006963f
C370 B.n333 VSUBS 0.006963f
C371 B.n334 VSUBS 0.006963f
C372 B.n335 VSUBS 0.006963f
C373 B.n336 VSUBS 0.006963f
C374 B.n337 VSUBS 0.006963f
C375 B.n338 VSUBS 0.006963f
C376 B.n339 VSUBS 0.006963f
C377 B.n340 VSUBS 0.006963f
C378 B.n341 VSUBS 0.006963f
C379 B.n342 VSUBS 0.006963f
C380 B.n343 VSUBS 0.006963f
C381 B.n344 VSUBS 0.006963f
C382 B.n345 VSUBS 0.006963f
C383 B.n346 VSUBS 0.006963f
C384 B.n347 VSUBS 0.006963f
C385 B.n348 VSUBS 0.006963f
C386 B.n349 VSUBS 0.006963f
C387 B.n350 VSUBS 0.006963f
C388 B.n351 VSUBS 0.006963f
C389 B.n352 VSUBS 0.006963f
C390 B.n353 VSUBS 0.006963f
C391 B.n354 VSUBS 0.006963f
C392 B.n355 VSUBS 0.006963f
C393 B.n356 VSUBS 0.006963f
C394 B.n357 VSUBS 0.006963f
C395 B.n358 VSUBS 0.006963f
C396 B.n359 VSUBS 0.006963f
C397 B.n360 VSUBS 0.006963f
C398 B.n361 VSUBS 0.006963f
C399 B.n362 VSUBS 0.006963f
C400 B.n363 VSUBS 0.006963f
C401 B.n364 VSUBS 0.006963f
C402 B.n365 VSUBS 0.006963f
C403 B.n366 VSUBS 0.006963f
C404 B.n367 VSUBS 0.006963f
C405 B.n368 VSUBS 0.006963f
C406 B.n369 VSUBS 0.006963f
C407 B.n370 VSUBS 0.006963f
C408 B.n371 VSUBS 0.006963f
C409 B.n372 VSUBS 0.006963f
C410 B.n373 VSUBS 0.006963f
C411 B.n374 VSUBS 0.006963f
C412 B.n375 VSUBS 0.006963f
C413 B.n376 VSUBS 0.006963f
C414 B.n377 VSUBS 0.006963f
C415 B.n378 VSUBS 0.006963f
C416 B.n379 VSUBS 0.006963f
C417 B.n380 VSUBS 0.006963f
C418 B.n381 VSUBS 0.006963f
C419 B.n382 VSUBS 0.006963f
C420 B.n383 VSUBS 0.006963f
C421 B.n384 VSUBS 0.006963f
C422 B.n385 VSUBS 0.006963f
C423 B.n386 VSUBS 0.006963f
C424 B.t2 VSUBS 0.276494f
C425 B.t1 VSUBS 0.312858f
C426 B.t0 VSUBS 1.9915f
C427 B.n387 VSUBS 0.491265f
C428 B.n388 VSUBS 0.290446f
C429 B.n389 VSUBS 0.016133f
C430 B.n390 VSUBS 0.006554f
C431 B.n391 VSUBS 0.006963f
C432 B.n392 VSUBS 0.006963f
C433 B.n393 VSUBS 0.006963f
C434 B.n394 VSUBS 0.006963f
C435 B.n395 VSUBS 0.006963f
C436 B.n396 VSUBS 0.006963f
C437 B.n397 VSUBS 0.006963f
C438 B.n398 VSUBS 0.006963f
C439 B.n399 VSUBS 0.006963f
C440 B.n400 VSUBS 0.006963f
C441 B.n401 VSUBS 0.006963f
C442 B.n402 VSUBS 0.006963f
C443 B.n403 VSUBS 0.006963f
C444 B.n404 VSUBS 0.006963f
C445 B.n405 VSUBS 0.006963f
C446 B.n406 VSUBS 0.003891f
C447 B.n407 VSUBS 0.016133f
C448 B.n408 VSUBS 0.006554f
C449 B.n409 VSUBS 0.006963f
C450 B.n410 VSUBS 0.006963f
C451 B.n411 VSUBS 0.006963f
C452 B.n412 VSUBS 0.006963f
C453 B.n413 VSUBS 0.006963f
C454 B.n414 VSUBS 0.006963f
C455 B.n415 VSUBS 0.006963f
C456 B.n416 VSUBS 0.006963f
C457 B.n417 VSUBS 0.006963f
C458 B.n418 VSUBS 0.006963f
C459 B.n419 VSUBS 0.006963f
C460 B.n420 VSUBS 0.006963f
C461 B.n421 VSUBS 0.006963f
C462 B.n422 VSUBS 0.006963f
C463 B.n423 VSUBS 0.006963f
C464 B.n424 VSUBS 0.006963f
C465 B.n425 VSUBS 0.006963f
C466 B.n426 VSUBS 0.006963f
C467 B.n427 VSUBS 0.006963f
C468 B.n428 VSUBS 0.006963f
C469 B.n429 VSUBS 0.006963f
C470 B.n430 VSUBS 0.006963f
C471 B.n431 VSUBS 0.006963f
C472 B.n432 VSUBS 0.006963f
C473 B.n433 VSUBS 0.006963f
C474 B.n434 VSUBS 0.006963f
C475 B.n435 VSUBS 0.006963f
C476 B.n436 VSUBS 0.006963f
C477 B.n437 VSUBS 0.006963f
C478 B.n438 VSUBS 0.006963f
C479 B.n439 VSUBS 0.006963f
C480 B.n440 VSUBS 0.006963f
C481 B.n441 VSUBS 0.006963f
C482 B.n442 VSUBS 0.006963f
C483 B.n443 VSUBS 0.006963f
C484 B.n444 VSUBS 0.006963f
C485 B.n445 VSUBS 0.006963f
C486 B.n446 VSUBS 0.006963f
C487 B.n447 VSUBS 0.006963f
C488 B.n448 VSUBS 0.006963f
C489 B.n449 VSUBS 0.006963f
C490 B.n450 VSUBS 0.006963f
C491 B.n451 VSUBS 0.006963f
C492 B.n452 VSUBS 0.006963f
C493 B.n453 VSUBS 0.006963f
C494 B.n454 VSUBS 0.006963f
C495 B.n455 VSUBS 0.006963f
C496 B.n456 VSUBS 0.006963f
C497 B.n457 VSUBS 0.006963f
C498 B.n458 VSUBS 0.006963f
C499 B.n459 VSUBS 0.006963f
C500 B.n460 VSUBS 0.006963f
C501 B.n461 VSUBS 0.006963f
C502 B.n462 VSUBS 0.006963f
C503 B.n463 VSUBS 0.006963f
C504 B.n464 VSUBS 0.006963f
C505 B.n465 VSUBS 0.006963f
C506 B.n466 VSUBS 0.006963f
C507 B.n467 VSUBS 0.006963f
C508 B.n468 VSUBS 0.006963f
C509 B.n469 VSUBS 0.006963f
C510 B.n470 VSUBS 0.006963f
C511 B.n471 VSUBS 0.006963f
C512 B.n472 VSUBS 0.006963f
C513 B.n473 VSUBS 0.006963f
C514 B.n474 VSUBS 0.006963f
C515 B.n475 VSUBS 0.006963f
C516 B.n476 VSUBS 0.006963f
C517 B.n477 VSUBS 0.006963f
C518 B.n478 VSUBS 0.006963f
C519 B.n479 VSUBS 0.006963f
C520 B.n480 VSUBS 0.006963f
C521 B.n481 VSUBS 0.015743f
C522 B.n482 VSUBS 0.016575f
C523 B.n483 VSUBS 0.015784f
C524 B.n484 VSUBS 0.006963f
C525 B.n485 VSUBS 0.006963f
C526 B.n486 VSUBS 0.006963f
C527 B.n487 VSUBS 0.006963f
C528 B.n488 VSUBS 0.006963f
C529 B.n489 VSUBS 0.006963f
C530 B.n490 VSUBS 0.006963f
C531 B.n491 VSUBS 0.006963f
C532 B.n492 VSUBS 0.006963f
C533 B.n493 VSUBS 0.006963f
C534 B.n494 VSUBS 0.006963f
C535 B.n495 VSUBS 0.006963f
C536 B.n496 VSUBS 0.006963f
C537 B.n497 VSUBS 0.006963f
C538 B.n498 VSUBS 0.006963f
C539 B.n499 VSUBS 0.006963f
C540 B.n500 VSUBS 0.006963f
C541 B.n501 VSUBS 0.006963f
C542 B.n502 VSUBS 0.006963f
C543 B.n503 VSUBS 0.006963f
C544 B.n504 VSUBS 0.006963f
C545 B.n505 VSUBS 0.006963f
C546 B.n506 VSUBS 0.006963f
C547 B.n507 VSUBS 0.006963f
C548 B.n508 VSUBS 0.006963f
C549 B.n509 VSUBS 0.006963f
C550 B.n510 VSUBS 0.006963f
C551 B.n511 VSUBS 0.006963f
C552 B.n512 VSUBS 0.006963f
C553 B.n513 VSUBS 0.006963f
C554 B.n514 VSUBS 0.006963f
C555 B.n515 VSUBS 0.006963f
C556 B.n516 VSUBS 0.006963f
C557 B.n517 VSUBS 0.006963f
C558 B.n518 VSUBS 0.006963f
C559 B.n519 VSUBS 0.006963f
C560 B.n520 VSUBS 0.006963f
C561 B.n521 VSUBS 0.006963f
C562 B.n522 VSUBS 0.006963f
C563 B.n523 VSUBS 0.006963f
C564 B.n524 VSUBS 0.006963f
C565 B.n525 VSUBS 0.006963f
C566 B.n526 VSUBS 0.006963f
C567 B.n527 VSUBS 0.006963f
C568 B.n528 VSUBS 0.006963f
C569 B.n529 VSUBS 0.006963f
C570 B.n530 VSUBS 0.006963f
C571 B.n531 VSUBS 0.006963f
C572 B.n532 VSUBS 0.006963f
C573 B.n533 VSUBS 0.006963f
C574 B.n534 VSUBS 0.006963f
C575 B.n535 VSUBS 0.006963f
C576 B.n536 VSUBS 0.006963f
C577 B.n537 VSUBS 0.006963f
C578 B.n538 VSUBS 0.006963f
C579 B.n539 VSUBS 0.006963f
C580 B.n540 VSUBS 0.006963f
C581 B.n541 VSUBS 0.006963f
C582 B.n542 VSUBS 0.006963f
C583 B.n543 VSUBS 0.006963f
C584 B.n544 VSUBS 0.006963f
C585 B.n545 VSUBS 0.006963f
C586 B.n546 VSUBS 0.006963f
C587 B.n547 VSUBS 0.006963f
C588 B.n548 VSUBS 0.006963f
C589 B.n549 VSUBS 0.006963f
C590 B.n550 VSUBS 0.006963f
C591 B.n551 VSUBS 0.006963f
C592 B.n552 VSUBS 0.006963f
C593 B.n553 VSUBS 0.006963f
C594 B.n554 VSUBS 0.006963f
C595 B.n555 VSUBS 0.006963f
C596 B.n556 VSUBS 0.006963f
C597 B.n557 VSUBS 0.006963f
C598 B.n558 VSUBS 0.006963f
C599 B.n559 VSUBS 0.006963f
C600 B.n560 VSUBS 0.006963f
C601 B.n561 VSUBS 0.006963f
C602 B.n562 VSUBS 0.006963f
C603 B.n563 VSUBS 0.006963f
C604 B.n564 VSUBS 0.006963f
C605 B.n565 VSUBS 0.006963f
C606 B.n566 VSUBS 0.006963f
C607 B.n567 VSUBS 0.006963f
C608 B.n568 VSUBS 0.006963f
C609 B.n569 VSUBS 0.006963f
C610 B.n570 VSUBS 0.006963f
C611 B.n571 VSUBS 0.006963f
C612 B.n572 VSUBS 0.006963f
C613 B.n573 VSUBS 0.006963f
C614 B.n574 VSUBS 0.006963f
C615 B.n575 VSUBS 0.006963f
C616 B.n576 VSUBS 0.006963f
C617 B.n577 VSUBS 0.006963f
C618 B.n578 VSUBS 0.006963f
C619 B.n579 VSUBS 0.006963f
C620 B.n580 VSUBS 0.006963f
C621 B.n581 VSUBS 0.006963f
C622 B.n582 VSUBS 0.006963f
C623 B.n583 VSUBS 0.006963f
C624 B.n584 VSUBS 0.006963f
C625 B.n585 VSUBS 0.006963f
C626 B.n586 VSUBS 0.006963f
C627 B.n587 VSUBS 0.006963f
C628 B.n588 VSUBS 0.006963f
C629 B.n589 VSUBS 0.006963f
C630 B.n590 VSUBS 0.006963f
C631 B.n591 VSUBS 0.006963f
C632 B.n592 VSUBS 0.006963f
C633 B.n593 VSUBS 0.006963f
C634 B.n594 VSUBS 0.006963f
C635 B.n595 VSUBS 0.006963f
C636 B.n596 VSUBS 0.006963f
C637 B.n597 VSUBS 0.006963f
C638 B.n598 VSUBS 0.006963f
C639 B.n599 VSUBS 0.006963f
C640 B.n600 VSUBS 0.006963f
C641 B.n601 VSUBS 0.006963f
C642 B.n602 VSUBS 0.006963f
C643 B.n603 VSUBS 0.006963f
C644 B.n604 VSUBS 0.006963f
C645 B.n605 VSUBS 0.006963f
C646 B.n606 VSUBS 0.006963f
C647 B.n607 VSUBS 0.006963f
C648 B.n608 VSUBS 0.006963f
C649 B.n609 VSUBS 0.006963f
C650 B.n610 VSUBS 0.006963f
C651 B.n611 VSUBS 0.006963f
C652 B.n612 VSUBS 0.006963f
C653 B.n613 VSUBS 0.006963f
C654 B.n614 VSUBS 0.006963f
C655 B.n615 VSUBS 0.006963f
C656 B.n616 VSUBS 0.006963f
C657 B.n617 VSUBS 0.006963f
C658 B.n618 VSUBS 0.006963f
C659 B.n619 VSUBS 0.006963f
C660 B.n620 VSUBS 0.006963f
C661 B.n621 VSUBS 0.006963f
C662 B.n622 VSUBS 0.006963f
C663 B.n623 VSUBS 0.006963f
C664 B.n624 VSUBS 0.006963f
C665 B.n625 VSUBS 0.006963f
C666 B.n626 VSUBS 0.006963f
C667 B.n627 VSUBS 0.006963f
C668 B.n628 VSUBS 0.006963f
C669 B.n629 VSUBS 0.006963f
C670 B.n630 VSUBS 0.006963f
C671 B.n631 VSUBS 0.006963f
C672 B.n632 VSUBS 0.006963f
C673 B.n633 VSUBS 0.006963f
C674 B.n634 VSUBS 0.006963f
C675 B.n635 VSUBS 0.006963f
C676 B.n636 VSUBS 0.006963f
C677 B.n637 VSUBS 0.006963f
C678 B.n638 VSUBS 0.006963f
C679 B.n639 VSUBS 0.006963f
C680 B.n640 VSUBS 0.006963f
C681 B.n641 VSUBS 0.006963f
C682 B.n642 VSUBS 0.006963f
C683 B.n643 VSUBS 0.006963f
C684 B.n644 VSUBS 0.006963f
C685 B.n645 VSUBS 0.006963f
C686 B.n646 VSUBS 0.006963f
C687 B.n647 VSUBS 0.006963f
C688 B.n648 VSUBS 0.006963f
C689 B.n649 VSUBS 0.006963f
C690 B.n650 VSUBS 0.006963f
C691 B.n651 VSUBS 0.006963f
C692 B.n652 VSUBS 0.015784f
C693 B.n653 VSUBS 0.015784f
C694 B.n654 VSUBS 0.016575f
C695 B.n655 VSUBS 0.006963f
C696 B.n656 VSUBS 0.006963f
C697 B.n657 VSUBS 0.006963f
C698 B.n658 VSUBS 0.006963f
C699 B.n659 VSUBS 0.006963f
C700 B.n660 VSUBS 0.006963f
C701 B.n661 VSUBS 0.006963f
C702 B.n662 VSUBS 0.006963f
C703 B.n663 VSUBS 0.006963f
C704 B.n664 VSUBS 0.006963f
C705 B.n665 VSUBS 0.006963f
C706 B.n666 VSUBS 0.006963f
C707 B.n667 VSUBS 0.006963f
C708 B.n668 VSUBS 0.006963f
C709 B.n669 VSUBS 0.006963f
C710 B.n670 VSUBS 0.006963f
C711 B.n671 VSUBS 0.006963f
C712 B.n672 VSUBS 0.006963f
C713 B.n673 VSUBS 0.006963f
C714 B.n674 VSUBS 0.006963f
C715 B.n675 VSUBS 0.006963f
C716 B.n676 VSUBS 0.006963f
C717 B.n677 VSUBS 0.006963f
C718 B.n678 VSUBS 0.006963f
C719 B.n679 VSUBS 0.006963f
C720 B.n680 VSUBS 0.006963f
C721 B.n681 VSUBS 0.006963f
C722 B.n682 VSUBS 0.006963f
C723 B.n683 VSUBS 0.006963f
C724 B.n684 VSUBS 0.006963f
C725 B.n685 VSUBS 0.006963f
C726 B.n686 VSUBS 0.006963f
C727 B.n687 VSUBS 0.006963f
C728 B.n688 VSUBS 0.006963f
C729 B.n689 VSUBS 0.006963f
C730 B.n690 VSUBS 0.006963f
C731 B.n691 VSUBS 0.006963f
C732 B.n692 VSUBS 0.006963f
C733 B.n693 VSUBS 0.006963f
C734 B.n694 VSUBS 0.006963f
C735 B.n695 VSUBS 0.006963f
C736 B.n696 VSUBS 0.006963f
C737 B.n697 VSUBS 0.006963f
C738 B.n698 VSUBS 0.006963f
C739 B.n699 VSUBS 0.006963f
C740 B.n700 VSUBS 0.006963f
C741 B.n701 VSUBS 0.006963f
C742 B.n702 VSUBS 0.006963f
C743 B.n703 VSUBS 0.006963f
C744 B.n704 VSUBS 0.006963f
C745 B.n705 VSUBS 0.006963f
C746 B.n706 VSUBS 0.006963f
C747 B.n707 VSUBS 0.006963f
C748 B.n708 VSUBS 0.006963f
C749 B.n709 VSUBS 0.006963f
C750 B.n710 VSUBS 0.006963f
C751 B.n711 VSUBS 0.006963f
C752 B.n712 VSUBS 0.006963f
C753 B.n713 VSUBS 0.006963f
C754 B.n714 VSUBS 0.006963f
C755 B.n715 VSUBS 0.006963f
C756 B.n716 VSUBS 0.006963f
C757 B.n717 VSUBS 0.006963f
C758 B.n718 VSUBS 0.006963f
C759 B.n719 VSUBS 0.006963f
C760 B.n720 VSUBS 0.006963f
C761 B.n721 VSUBS 0.006963f
C762 B.n722 VSUBS 0.006963f
C763 B.n723 VSUBS 0.006963f
C764 B.n724 VSUBS 0.006963f
C765 B.n725 VSUBS 0.006963f
C766 B.n726 VSUBS 0.006963f
C767 B.n727 VSUBS 0.006554f
C768 B.n728 VSUBS 0.006963f
C769 B.n729 VSUBS 0.006963f
C770 B.n730 VSUBS 0.003891f
C771 B.n731 VSUBS 0.006963f
C772 B.n732 VSUBS 0.006963f
C773 B.n733 VSUBS 0.006963f
C774 B.n734 VSUBS 0.006963f
C775 B.n735 VSUBS 0.006963f
C776 B.n736 VSUBS 0.006963f
C777 B.n737 VSUBS 0.006963f
C778 B.n738 VSUBS 0.006963f
C779 B.n739 VSUBS 0.006963f
C780 B.n740 VSUBS 0.006963f
C781 B.n741 VSUBS 0.006963f
C782 B.n742 VSUBS 0.006963f
C783 B.n743 VSUBS 0.003891f
C784 B.n744 VSUBS 0.016133f
C785 B.n745 VSUBS 0.006554f
C786 B.n746 VSUBS 0.006963f
C787 B.n747 VSUBS 0.006963f
C788 B.n748 VSUBS 0.006963f
C789 B.n749 VSUBS 0.006963f
C790 B.n750 VSUBS 0.006963f
C791 B.n751 VSUBS 0.006963f
C792 B.n752 VSUBS 0.006963f
C793 B.n753 VSUBS 0.006963f
C794 B.n754 VSUBS 0.006963f
C795 B.n755 VSUBS 0.006963f
C796 B.n756 VSUBS 0.006963f
C797 B.n757 VSUBS 0.006963f
C798 B.n758 VSUBS 0.006963f
C799 B.n759 VSUBS 0.006963f
C800 B.n760 VSUBS 0.006963f
C801 B.n761 VSUBS 0.006963f
C802 B.n762 VSUBS 0.006963f
C803 B.n763 VSUBS 0.006963f
C804 B.n764 VSUBS 0.006963f
C805 B.n765 VSUBS 0.006963f
C806 B.n766 VSUBS 0.006963f
C807 B.n767 VSUBS 0.006963f
C808 B.n768 VSUBS 0.006963f
C809 B.n769 VSUBS 0.006963f
C810 B.n770 VSUBS 0.006963f
C811 B.n771 VSUBS 0.006963f
C812 B.n772 VSUBS 0.006963f
C813 B.n773 VSUBS 0.006963f
C814 B.n774 VSUBS 0.006963f
C815 B.n775 VSUBS 0.006963f
C816 B.n776 VSUBS 0.006963f
C817 B.n777 VSUBS 0.006963f
C818 B.n778 VSUBS 0.006963f
C819 B.n779 VSUBS 0.006963f
C820 B.n780 VSUBS 0.006963f
C821 B.n781 VSUBS 0.006963f
C822 B.n782 VSUBS 0.006963f
C823 B.n783 VSUBS 0.006963f
C824 B.n784 VSUBS 0.006963f
C825 B.n785 VSUBS 0.006963f
C826 B.n786 VSUBS 0.006963f
C827 B.n787 VSUBS 0.006963f
C828 B.n788 VSUBS 0.006963f
C829 B.n789 VSUBS 0.006963f
C830 B.n790 VSUBS 0.006963f
C831 B.n791 VSUBS 0.006963f
C832 B.n792 VSUBS 0.006963f
C833 B.n793 VSUBS 0.006963f
C834 B.n794 VSUBS 0.006963f
C835 B.n795 VSUBS 0.006963f
C836 B.n796 VSUBS 0.006963f
C837 B.n797 VSUBS 0.006963f
C838 B.n798 VSUBS 0.006963f
C839 B.n799 VSUBS 0.006963f
C840 B.n800 VSUBS 0.006963f
C841 B.n801 VSUBS 0.006963f
C842 B.n802 VSUBS 0.006963f
C843 B.n803 VSUBS 0.006963f
C844 B.n804 VSUBS 0.006963f
C845 B.n805 VSUBS 0.006963f
C846 B.n806 VSUBS 0.006963f
C847 B.n807 VSUBS 0.006963f
C848 B.n808 VSUBS 0.006963f
C849 B.n809 VSUBS 0.006963f
C850 B.n810 VSUBS 0.006963f
C851 B.n811 VSUBS 0.006963f
C852 B.n812 VSUBS 0.006963f
C853 B.n813 VSUBS 0.006963f
C854 B.n814 VSUBS 0.006963f
C855 B.n815 VSUBS 0.006963f
C856 B.n816 VSUBS 0.006963f
C857 B.n817 VSUBS 0.006963f
C858 B.n818 VSUBS 0.006963f
C859 B.n819 VSUBS 0.016575f
C860 B.n820 VSUBS 0.015784f
C861 B.n821 VSUBS 0.015784f
C862 B.n822 VSUBS 0.006963f
C863 B.n823 VSUBS 0.006963f
C864 B.n824 VSUBS 0.006963f
C865 B.n825 VSUBS 0.006963f
C866 B.n826 VSUBS 0.006963f
C867 B.n827 VSUBS 0.006963f
C868 B.n828 VSUBS 0.006963f
C869 B.n829 VSUBS 0.006963f
C870 B.n830 VSUBS 0.006963f
C871 B.n831 VSUBS 0.006963f
C872 B.n832 VSUBS 0.006963f
C873 B.n833 VSUBS 0.006963f
C874 B.n834 VSUBS 0.006963f
C875 B.n835 VSUBS 0.006963f
C876 B.n836 VSUBS 0.006963f
C877 B.n837 VSUBS 0.006963f
C878 B.n838 VSUBS 0.006963f
C879 B.n839 VSUBS 0.006963f
C880 B.n840 VSUBS 0.006963f
C881 B.n841 VSUBS 0.006963f
C882 B.n842 VSUBS 0.006963f
C883 B.n843 VSUBS 0.006963f
C884 B.n844 VSUBS 0.006963f
C885 B.n845 VSUBS 0.006963f
C886 B.n846 VSUBS 0.006963f
C887 B.n847 VSUBS 0.006963f
C888 B.n848 VSUBS 0.006963f
C889 B.n849 VSUBS 0.006963f
C890 B.n850 VSUBS 0.006963f
C891 B.n851 VSUBS 0.006963f
C892 B.n852 VSUBS 0.006963f
C893 B.n853 VSUBS 0.006963f
C894 B.n854 VSUBS 0.006963f
C895 B.n855 VSUBS 0.006963f
C896 B.n856 VSUBS 0.006963f
C897 B.n857 VSUBS 0.006963f
C898 B.n858 VSUBS 0.006963f
C899 B.n859 VSUBS 0.006963f
C900 B.n860 VSUBS 0.006963f
C901 B.n861 VSUBS 0.006963f
C902 B.n862 VSUBS 0.006963f
C903 B.n863 VSUBS 0.006963f
C904 B.n864 VSUBS 0.006963f
C905 B.n865 VSUBS 0.006963f
C906 B.n866 VSUBS 0.006963f
C907 B.n867 VSUBS 0.006963f
C908 B.n868 VSUBS 0.006963f
C909 B.n869 VSUBS 0.006963f
C910 B.n870 VSUBS 0.006963f
C911 B.n871 VSUBS 0.006963f
C912 B.n872 VSUBS 0.006963f
C913 B.n873 VSUBS 0.006963f
C914 B.n874 VSUBS 0.006963f
C915 B.n875 VSUBS 0.006963f
C916 B.n876 VSUBS 0.006963f
C917 B.n877 VSUBS 0.006963f
C918 B.n878 VSUBS 0.006963f
C919 B.n879 VSUBS 0.006963f
C920 B.n880 VSUBS 0.006963f
C921 B.n881 VSUBS 0.006963f
C922 B.n882 VSUBS 0.006963f
C923 B.n883 VSUBS 0.006963f
C924 B.n884 VSUBS 0.006963f
C925 B.n885 VSUBS 0.006963f
C926 B.n886 VSUBS 0.006963f
C927 B.n887 VSUBS 0.006963f
C928 B.n888 VSUBS 0.006963f
C929 B.n889 VSUBS 0.006963f
C930 B.n890 VSUBS 0.006963f
C931 B.n891 VSUBS 0.006963f
C932 B.n892 VSUBS 0.006963f
C933 B.n893 VSUBS 0.006963f
C934 B.n894 VSUBS 0.006963f
C935 B.n895 VSUBS 0.006963f
C936 B.n896 VSUBS 0.006963f
C937 B.n897 VSUBS 0.006963f
C938 B.n898 VSUBS 0.006963f
C939 B.n899 VSUBS 0.006963f
C940 B.n900 VSUBS 0.006963f
C941 B.n901 VSUBS 0.006963f
C942 B.n902 VSUBS 0.006963f
C943 B.n903 VSUBS 0.009087f
C944 B.n904 VSUBS 0.00968f
C945 B.n905 VSUBS 0.019249f
C946 VDD1.t6 VSUBS 0.320553f
C947 VDD1.t3 VSUBS 0.320553f
C948 VDD1.n0 VSUBS 2.59971f
C949 VDD1.t2 VSUBS 0.320553f
C950 VDD1.t0 VSUBS 0.320553f
C951 VDD1.n1 VSUBS 2.59806f
C952 VDD1.t7 VSUBS 0.320553f
C953 VDD1.t5 VSUBS 0.320553f
C954 VDD1.n2 VSUBS 2.59806f
C955 VDD1.n3 VSUBS 4.6686f
C956 VDD1.t1 VSUBS 0.320553f
C957 VDD1.t4 VSUBS 0.320553f
C958 VDD1.n4 VSUBS 2.58041f
C959 VDD1.n5 VSUBS 3.93394f
C960 VP.t2 VSUBS 3.34119f
C961 VP.n0 VSUBS 1.27403f
C962 VP.n1 VSUBS 0.027613f
C963 VP.n2 VSUBS 0.043196f
C964 VP.n3 VSUBS 0.027613f
C965 VP.t0 VSUBS 3.34119f
C966 VP.n4 VSUBS 0.051206f
C967 VP.n5 VSUBS 0.027613f
C968 VP.n6 VSUBS 0.051206f
C969 VP.n7 VSUBS 0.027613f
C970 VP.t7 VSUBS 3.34119f
C971 VP.n8 VSUBS 0.043196f
C972 VP.n9 VSUBS 0.027613f
C973 VP.t5 VSUBS 3.34119f
C974 VP.n10 VSUBS 1.27403f
C975 VP.t3 VSUBS 3.34119f
C976 VP.n11 VSUBS 1.27403f
C977 VP.n12 VSUBS 0.027613f
C978 VP.n13 VSUBS 0.043196f
C979 VP.n14 VSUBS 0.027613f
C980 VP.t6 VSUBS 3.34119f
C981 VP.n15 VSUBS 0.051206f
C982 VP.n16 VSUBS 0.027613f
C983 VP.n17 VSUBS 0.051206f
C984 VP.t1 VSUBS 3.62098f
C985 VP.n18 VSUBS 1.21105f
C986 VP.t4 VSUBS 3.34119f
C987 VP.n19 VSUBS 1.24596f
C988 VP.n20 VSUBS 0.033258f
C989 VP.n21 VSUBS 0.296651f
C990 VP.n22 VSUBS 0.027613f
C991 VP.n23 VSUBS 0.027613f
C992 VP.n24 VSUBS 0.054591f
C993 VP.n25 VSUBS 0.022302f
C994 VP.n26 VSUBS 0.054591f
C995 VP.n27 VSUBS 0.027613f
C996 VP.n28 VSUBS 0.027613f
C997 VP.n29 VSUBS 0.027613f
C998 VP.n30 VSUBS 0.033258f
C999 VP.n31 VSUBS 1.16446f
C1000 VP.n32 VSUBS 0.043875f
C1001 VP.n33 VSUBS 0.051206f
C1002 VP.n34 VSUBS 0.027613f
C1003 VP.n35 VSUBS 0.027613f
C1004 VP.n36 VSUBS 0.027613f
C1005 VP.n37 VSUBS 0.037084f
C1006 VP.n38 VSUBS 0.051206f
C1007 VP.n39 VSUBS 0.047919f
C1008 VP.n40 VSUBS 0.04456f
C1009 VP.n41 VSUBS 1.78104f
C1010 VP.n42 VSUBS 1.79916f
C1011 VP.n43 VSUBS 0.04456f
C1012 VP.n44 VSUBS 0.047919f
C1013 VP.n45 VSUBS 0.051206f
C1014 VP.n46 VSUBS 0.037084f
C1015 VP.n47 VSUBS 0.027613f
C1016 VP.n48 VSUBS 0.027613f
C1017 VP.n49 VSUBS 0.027613f
C1018 VP.n50 VSUBS 0.051206f
C1019 VP.n51 VSUBS 0.043875f
C1020 VP.n52 VSUBS 1.16446f
C1021 VP.n53 VSUBS 0.033258f
C1022 VP.n54 VSUBS 0.027613f
C1023 VP.n55 VSUBS 0.027613f
C1024 VP.n56 VSUBS 0.027613f
C1025 VP.n57 VSUBS 0.054591f
C1026 VP.n58 VSUBS 0.022302f
C1027 VP.n59 VSUBS 0.054591f
C1028 VP.n60 VSUBS 0.027613f
C1029 VP.n61 VSUBS 0.027613f
C1030 VP.n62 VSUBS 0.027613f
C1031 VP.n63 VSUBS 0.033258f
C1032 VP.n64 VSUBS 1.16446f
C1033 VP.n65 VSUBS 0.043875f
C1034 VP.n66 VSUBS 0.051206f
C1035 VP.n67 VSUBS 0.027613f
C1036 VP.n68 VSUBS 0.027613f
C1037 VP.n69 VSUBS 0.027613f
C1038 VP.n70 VSUBS 0.037084f
C1039 VP.n71 VSUBS 0.051206f
C1040 VP.n72 VSUBS 0.047919f
C1041 VP.n73 VSUBS 0.04456f
C1042 VP.n74 VSUBS 0.055435f
C1043 VTAIL.t13 VSUBS 0.289619f
C1044 VTAIL.t12 VSUBS 0.289619f
C1045 VTAIL.n0 VSUBS 2.17914f
C1046 VTAIL.n1 VSUBS 0.834846f
C1047 VTAIL.n2 VSUBS 0.027721f
C1048 VTAIL.n3 VSUBS 0.024564f
C1049 VTAIL.n4 VSUBS 0.0132f
C1050 VTAIL.n5 VSUBS 0.031199f
C1051 VTAIL.n6 VSUBS 0.013976f
C1052 VTAIL.n7 VSUBS 0.024564f
C1053 VTAIL.n8 VSUBS 0.0132f
C1054 VTAIL.n9 VSUBS 0.031199f
C1055 VTAIL.n10 VSUBS 0.013976f
C1056 VTAIL.n11 VSUBS 0.024564f
C1057 VTAIL.n12 VSUBS 0.0132f
C1058 VTAIL.n13 VSUBS 0.031199f
C1059 VTAIL.n14 VSUBS 0.013976f
C1060 VTAIL.n15 VSUBS 0.024564f
C1061 VTAIL.n16 VSUBS 0.0132f
C1062 VTAIL.n17 VSUBS 0.031199f
C1063 VTAIL.n18 VSUBS 0.013976f
C1064 VTAIL.n19 VSUBS 0.024564f
C1065 VTAIL.n20 VSUBS 0.0132f
C1066 VTAIL.n21 VSUBS 0.031199f
C1067 VTAIL.n22 VSUBS 0.013976f
C1068 VTAIL.n23 VSUBS 0.024564f
C1069 VTAIL.n24 VSUBS 0.0132f
C1070 VTAIL.n25 VSUBS 0.031199f
C1071 VTAIL.n26 VSUBS 0.013976f
C1072 VTAIL.n27 VSUBS 0.225888f
C1073 VTAIL.t9 VSUBS 0.067471f
C1074 VTAIL.n28 VSUBS 0.0234f
C1075 VTAIL.n29 VSUBS 0.02347f
C1076 VTAIL.n30 VSUBS 0.0132f
C1077 VTAIL.n31 VSUBS 1.52121f
C1078 VTAIL.n32 VSUBS 0.024564f
C1079 VTAIL.n33 VSUBS 0.0132f
C1080 VTAIL.n34 VSUBS 0.013976f
C1081 VTAIL.n35 VSUBS 0.031199f
C1082 VTAIL.n36 VSUBS 0.031199f
C1083 VTAIL.n37 VSUBS 0.013976f
C1084 VTAIL.n38 VSUBS 0.0132f
C1085 VTAIL.n39 VSUBS 0.024564f
C1086 VTAIL.n40 VSUBS 0.024564f
C1087 VTAIL.n41 VSUBS 0.0132f
C1088 VTAIL.n42 VSUBS 0.013976f
C1089 VTAIL.n43 VSUBS 0.031199f
C1090 VTAIL.n44 VSUBS 0.031199f
C1091 VTAIL.n45 VSUBS 0.031199f
C1092 VTAIL.n46 VSUBS 0.013976f
C1093 VTAIL.n47 VSUBS 0.0132f
C1094 VTAIL.n48 VSUBS 0.024564f
C1095 VTAIL.n49 VSUBS 0.024564f
C1096 VTAIL.n50 VSUBS 0.0132f
C1097 VTAIL.n51 VSUBS 0.013588f
C1098 VTAIL.n52 VSUBS 0.013588f
C1099 VTAIL.n53 VSUBS 0.031199f
C1100 VTAIL.n54 VSUBS 0.031199f
C1101 VTAIL.n55 VSUBS 0.013976f
C1102 VTAIL.n56 VSUBS 0.0132f
C1103 VTAIL.n57 VSUBS 0.024564f
C1104 VTAIL.n58 VSUBS 0.024564f
C1105 VTAIL.n59 VSUBS 0.0132f
C1106 VTAIL.n60 VSUBS 0.013976f
C1107 VTAIL.n61 VSUBS 0.031199f
C1108 VTAIL.n62 VSUBS 0.031199f
C1109 VTAIL.n63 VSUBS 0.013976f
C1110 VTAIL.n64 VSUBS 0.0132f
C1111 VTAIL.n65 VSUBS 0.024564f
C1112 VTAIL.n66 VSUBS 0.024564f
C1113 VTAIL.n67 VSUBS 0.0132f
C1114 VTAIL.n68 VSUBS 0.013976f
C1115 VTAIL.n69 VSUBS 0.031199f
C1116 VTAIL.n70 VSUBS 0.031199f
C1117 VTAIL.n71 VSUBS 0.013976f
C1118 VTAIL.n72 VSUBS 0.0132f
C1119 VTAIL.n73 VSUBS 0.024564f
C1120 VTAIL.n74 VSUBS 0.024564f
C1121 VTAIL.n75 VSUBS 0.0132f
C1122 VTAIL.n76 VSUBS 0.013976f
C1123 VTAIL.n77 VSUBS 0.031199f
C1124 VTAIL.n78 VSUBS 0.078018f
C1125 VTAIL.n79 VSUBS 0.013976f
C1126 VTAIL.n80 VSUBS 0.0132f
C1127 VTAIL.n81 VSUBS 0.054095f
C1128 VTAIL.n82 VSUBS 0.039261f
C1129 VTAIL.n83 VSUBS 0.281145f
C1130 VTAIL.n84 VSUBS 0.027721f
C1131 VTAIL.n85 VSUBS 0.024564f
C1132 VTAIL.n86 VSUBS 0.0132f
C1133 VTAIL.n87 VSUBS 0.031199f
C1134 VTAIL.n88 VSUBS 0.013976f
C1135 VTAIL.n89 VSUBS 0.024564f
C1136 VTAIL.n90 VSUBS 0.0132f
C1137 VTAIL.n91 VSUBS 0.031199f
C1138 VTAIL.n92 VSUBS 0.013976f
C1139 VTAIL.n93 VSUBS 0.024564f
C1140 VTAIL.n94 VSUBS 0.0132f
C1141 VTAIL.n95 VSUBS 0.031199f
C1142 VTAIL.n96 VSUBS 0.013976f
C1143 VTAIL.n97 VSUBS 0.024564f
C1144 VTAIL.n98 VSUBS 0.0132f
C1145 VTAIL.n99 VSUBS 0.031199f
C1146 VTAIL.n100 VSUBS 0.013976f
C1147 VTAIL.n101 VSUBS 0.024564f
C1148 VTAIL.n102 VSUBS 0.0132f
C1149 VTAIL.n103 VSUBS 0.031199f
C1150 VTAIL.n104 VSUBS 0.013976f
C1151 VTAIL.n105 VSUBS 0.024564f
C1152 VTAIL.n106 VSUBS 0.0132f
C1153 VTAIL.n107 VSUBS 0.031199f
C1154 VTAIL.n108 VSUBS 0.013976f
C1155 VTAIL.n109 VSUBS 0.225888f
C1156 VTAIL.t0 VSUBS 0.067471f
C1157 VTAIL.n110 VSUBS 0.0234f
C1158 VTAIL.n111 VSUBS 0.02347f
C1159 VTAIL.n112 VSUBS 0.0132f
C1160 VTAIL.n113 VSUBS 1.52121f
C1161 VTAIL.n114 VSUBS 0.024564f
C1162 VTAIL.n115 VSUBS 0.0132f
C1163 VTAIL.n116 VSUBS 0.013976f
C1164 VTAIL.n117 VSUBS 0.031199f
C1165 VTAIL.n118 VSUBS 0.031199f
C1166 VTAIL.n119 VSUBS 0.013976f
C1167 VTAIL.n120 VSUBS 0.0132f
C1168 VTAIL.n121 VSUBS 0.024564f
C1169 VTAIL.n122 VSUBS 0.024564f
C1170 VTAIL.n123 VSUBS 0.0132f
C1171 VTAIL.n124 VSUBS 0.013976f
C1172 VTAIL.n125 VSUBS 0.031199f
C1173 VTAIL.n126 VSUBS 0.031199f
C1174 VTAIL.n127 VSUBS 0.031199f
C1175 VTAIL.n128 VSUBS 0.013976f
C1176 VTAIL.n129 VSUBS 0.0132f
C1177 VTAIL.n130 VSUBS 0.024564f
C1178 VTAIL.n131 VSUBS 0.024564f
C1179 VTAIL.n132 VSUBS 0.0132f
C1180 VTAIL.n133 VSUBS 0.013588f
C1181 VTAIL.n134 VSUBS 0.013588f
C1182 VTAIL.n135 VSUBS 0.031199f
C1183 VTAIL.n136 VSUBS 0.031199f
C1184 VTAIL.n137 VSUBS 0.013976f
C1185 VTAIL.n138 VSUBS 0.0132f
C1186 VTAIL.n139 VSUBS 0.024564f
C1187 VTAIL.n140 VSUBS 0.024564f
C1188 VTAIL.n141 VSUBS 0.0132f
C1189 VTAIL.n142 VSUBS 0.013976f
C1190 VTAIL.n143 VSUBS 0.031199f
C1191 VTAIL.n144 VSUBS 0.031199f
C1192 VTAIL.n145 VSUBS 0.013976f
C1193 VTAIL.n146 VSUBS 0.0132f
C1194 VTAIL.n147 VSUBS 0.024564f
C1195 VTAIL.n148 VSUBS 0.024564f
C1196 VTAIL.n149 VSUBS 0.0132f
C1197 VTAIL.n150 VSUBS 0.013976f
C1198 VTAIL.n151 VSUBS 0.031199f
C1199 VTAIL.n152 VSUBS 0.031199f
C1200 VTAIL.n153 VSUBS 0.013976f
C1201 VTAIL.n154 VSUBS 0.0132f
C1202 VTAIL.n155 VSUBS 0.024564f
C1203 VTAIL.n156 VSUBS 0.024564f
C1204 VTAIL.n157 VSUBS 0.0132f
C1205 VTAIL.n158 VSUBS 0.013976f
C1206 VTAIL.n159 VSUBS 0.031199f
C1207 VTAIL.n160 VSUBS 0.078018f
C1208 VTAIL.n161 VSUBS 0.013976f
C1209 VTAIL.n162 VSUBS 0.0132f
C1210 VTAIL.n163 VSUBS 0.054095f
C1211 VTAIL.n164 VSUBS 0.039261f
C1212 VTAIL.n165 VSUBS 0.281145f
C1213 VTAIL.t6 VSUBS 0.289619f
C1214 VTAIL.t4 VSUBS 0.289619f
C1215 VTAIL.n166 VSUBS 2.17914f
C1216 VTAIL.n167 VSUBS 1.05473f
C1217 VTAIL.n168 VSUBS 0.027721f
C1218 VTAIL.n169 VSUBS 0.024564f
C1219 VTAIL.n170 VSUBS 0.0132f
C1220 VTAIL.n171 VSUBS 0.031199f
C1221 VTAIL.n172 VSUBS 0.013976f
C1222 VTAIL.n173 VSUBS 0.024564f
C1223 VTAIL.n174 VSUBS 0.0132f
C1224 VTAIL.n175 VSUBS 0.031199f
C1225 VTAIL.n176 VSUBS 0.013976f
C1226 VTAIL.n177 VSUBS 0.024564f
C1227 VTAIL.n178 VSUBS 0.0132f
C1228 VTAIL.n179 VSUBS 0.031199f
C1229 VTAIL.n180 VSUBS 0.013976f
C1230 VTAIL.n181 VSUBS 0.024564f
C1231 VTAIL.n182 VSUBS 0.0132f
C1232 VTAIL.n183 VSUBS 0.031199f
C1233 VTAIL.n184 VSUBS 0.013976f
C1234 VTAIL.n185 VSUBS 0.024564f
C1235 VTAIL.n186 VSUBS 0.0132f
C1236 VTAIL.n187 VSUBS 0.031199f
C1237 VTAIL.n188 VSUBS 0.013976f
C1238 VTAIL.n189 VSUBS 0.024564f
C1239 VTAIL.n190 VSUBS 0.0132f
C1240 VTAIL.n191 VSUBS 0.031199f
C1241 VTAIL.n192 VSUBS 0.013976f
C1242 VTAIL.n193 VSUBS 0.225888f
C1243 VTAIL.t3 VSUBS 0.067471f
C1244 VTAIL.n194 VSUBS 0.0234f
C1245 VTAIL.n195 VSUBS 0.02347f
C1246 VTAIL.n196 VSUBS 0.0132f
C1247 VTAIL.n197 VSUBS 1.52121f
C1248 VTAIL.n198 VSUBS 0.024564f
C1249 VTAIL.n199 VSUBS 0.0132f
C1250 VTAIL.n200 VSUBS 0.013976f
C1251 VTAIL.n201 VSUBS 0.031199f
C1252 VTAIL.n202 VSUBS 0.031199f
C1253 VTAIL.n203 VSUBS 0.013976f
C1254 VTAIL.n204 VSUBS 0.0132f
C1255 VTAIL.n205 VSUBS 0.024564f
C1256 VTAIL.n206 VSUBS 0.024564f
C1257 VTAIL.n207 VSUBS 0.0132f
C1258 VTAIL.n208 VSUBS 0.013976f
C1259 VTAIL.n209 VSUBS 0.031199f
C1260 VTAIL.n210 VSUBS 0.031199f
C1261 VTAIL.n211 VSUBS 0.031199f
C1262 VTAIL.n212 VSUBS 0.013976f
C1263 VTAIL.n213 VSUBS 0.0132f
C1264 VTAIL.n214 VSUBS 0.024564f
C1265 VTAIL.n215 VSUBS 0.024564f
C1266 VTAIL.n216 VSUBS 0.0132f
C1267 VTAIL.n217 VSUBS 0.013588f
C1268 VTAIL.n218 VSUBS 0.013588f
C1269 VTAIL.n219 VSUBS 0.031199f
C1270 VTAIL.n220 VSUBS 0.031199f
C1271 VTAIL.n221 VSUBS 0.013976f
C1272 VTAIL.n222 VSUBS 0.0132f
C1273 VTAIL.n223 VSUBS 0.024564f
C1274 VTAIL.n224 VSUBS 0.024564f
C1275 VTAIL.n225 VSUBS 0.0132f
C1276 VTAIL.n226 VSUBS 0.013976f
C1277 VTAIL.n227 VSUBS 0.031199f
C1278 VTAIL.n228 VSUBS 0.031199f
C1279 VTAIL.n229 VSUBS 0.013976f
C1280 VTAIL.n230 VSUBS 0.0132f
C1281 VTAIL.n231 VSUBS 0.024564f
C1282 VTAIL.n232 VSUBS 0.024564f
C1283 VTAIL.n233 VSUBS 0.0132f
C1284 VTAIL.n234 VSUBS 0.013976f
C1285 VTAIL.n235 VSUBS 0.031199f
C1286 VTAIL.n236 VSUBS 0.031199f
C1287 VTAIL.n237 VSUBS 0.013976f
C1288 VTAIL.n238 VSUBS 0.0132f
C1289 VTAIL.n239 VSUBS 0.024564f
C1290 VTAIL.n240 VSUBS 0.024564f
C1291 VTAIL.n241 VSUBS 0.0132f
C1292 VTAIL.n242 VSUBS 0.013976f
C1293 VTAIL.n243 VSUBS 0.031199f
C1294 VTAIL.n244 VSUBS 0.078018f
C1295 VTAIL.n245 VSUBS 0.013976f
C1296 VTAIL.n246 VSUBS 0.0132f
C1297 VTAIL.n247 VSUBS 0.054095f
C1298 VTAIL.n248 VSUBS 0.039261f
C1299 VTAIL.n249 VSUBS 1.82018f
C1300 VTAIL.n250 VSUBS 0.027721f
C1301 VTAIL.n251 VSUBS 0.024564f
C1302 VTAIL.n252 VSUBS 0.0132f
C1303 VTAIL.n253 VSUBS 0.031199f
C1304 VTAIL.n254 VSUBS 0.013976f
C1305 VTAIL.n255 VSUBS 0.024564f
C1306 VTAIL.n256 VSUBS 0.0132f
C1307 VTAIL.n257 VSUBS 0.031199f
C1308 VTAIL.n258 VSUBS 0.013976f
C1309 VTAIL.n259 VSUBS 0.024564f
C1310 VTAIL.n260 VSUBS 0.0132f
C1311 VTAIL.n261 VSUBS 0.031199f
C1312 VTAIL.n262 VSUBS 0.013976f
C1313 VTAIL.n263 VSUBS 0.024564f
C1314 VTAIL.n264 VSUBS 0.0132f
C1315 VTAIL.n265 VSUBS 0.031199f
C1316 VTAIL.n266 VSUBS 0.013976f
C1317 VTAIL.n267 VSUBS 0.024564f
C1318 VTAIL.n268 VSUBS 0.0132f
C1319 VTAIL.n269 VSUBS 0.031199f
C1320 VTAIL.n270 VSUBS 0.031199f
C1321 VTAIL.n271 VSUBS 0.013976f
C1322 VTAIL.n272 VSUBS 0.024564f
C1323 VTAIL.n273 VSUBS 0.0132f
C1324 VTAIL.n274 VSUBS 0.031199f
C1325 VTAIL.n275 VSUBS 0.013976f
C1326 VTAIL.n276 VSUBS 0.225888f
C1327 VTAIL.t8 VSUBS 0.067471f
C1328 VTAIL.n277 VSUBS 0.0234f
C1329 VTAIL.n278 VSUBS 0.02347f
C1330 VTAIL.n279 VSUBS 0.0132f
C1331 VTAIL.n280 VSUBS 1.52121f
C1332 VTAIL.n281 VSUBS 0.024564f
C1333 VTAIL.n282 VSUBS 0.0132f
C1334 VTAIL.n283 VSUBS 0.013976f
C1335 VTAIL.n284 VSUBS 0.031199f
C1336 VTAIL.n285 VSUBS 0.031199f
C1337 VTAIL.n286 VSUBS 0.013976f
C1338 VTAIL.n287 VSUBS 0.0132f
C1339 VTAIL.n288 VSUBS 0.024564f
C1340 VTAIL.n289 VSUBS 0.024564f
C1341 VTAIL.n290 VSUBS 0.0132f
C1342 VTAIL.n291 VSUBS 0.013976f
C1343 VTAIL.n292 VSUBS 0.031199f
C1344 VTAIL.n293 VSUBS 0.031199f
C1345 VTAIL.n294 VSUBS 0.013976f
C1346 VTAIL.n295 VSUBS 0.0132f
C1347 VTAIL.n296 VSUBS 0.024564f
C1348 VTAIL.n297 VSUBS 0.024564f
C1349 VTAIL.n298 VSUBS 0.0132f
C1350 VTAIL.n299 VSUBS 0.013588f
C1351 VTAIL.n300 VSUBS 0.013588f
C1352 VTAIL.n301 VSUBS 0.031199f
C1353 VTAIL.n302 VSUBS 0.031199f
C1354 VTAIL.n303 VSUBS 0.013976f
C1355 VTAIL.n304 VSUBS 0.0132f
C1356 VTAIL.n305 VSUBS 0.024564f
C1357 VTAIL.n306 VSUBS 0.024564f
C1358 VTAIL.n307 VSUBS 0.0132f
C1359 VTAIL.n308 VSUBS 0.013976f
C1360 VTAIL.n309 VSUBS 0.031199f
C1361 VTAIL.n310 VSUBS 0.031199f
C1362 VTAIL.n311 VSUBS 0.013976f
C1363 VTAIL.n312 VSUBS 0.0132f
C1364 VTAIL.n313 VSUBS 0.024564f
C1365 VTAIL.n314 VSUBS 0.024564f
C1366 VTAIL.n315 VSUBS 0.0132f
C1367 VTAIL.n316 VSUBS 0.013976f
C1368 VTAIL.n317 VSUBS 0.031199f
C1369 VTAIL.n318 VSUBS 0.031199f
C1370 VTAIL.n319 VSUBS 0.013976f
C1371 VTAIL.n320 VSUBS 0.0132f
C1372 VTAIL.n321 VSUBS 0.024564f
C1373 VTAIL.n322 VSUBS 0.024564f
C1374 VTAIL.n323 VSUBS 0.0132f
C1375 VTAIL.n324 VSUBS 0.013976f
C1376 VTAIL.n325 VSUBS 0.031199f
C1377 VTAIL.n326 VSUBS 0.078018f
C1378 VTAIL.n327 VSUBS 0.013976f
C1379 VTAIL.n328 VSUBS 0.0132f
C1380 VTAIL.n329 VSUBS 0.054095f
C1381 VTAIL.n330 VSUBS 0.039261f
C1382 VTAIL.n331 VSUBS 1.82018f
C1383 VTAIL.t10 VSUBS 0.289619f
C1384 VTAIL.t15 VSUBS 0.289619f
C1385 VTAIL.n332 VSUBS 2.17915f
C1386 VTAIL.n333 VSUBS 1.05472f
C1387 VTAIL.n334 VSUBS 0.027721f
C1388 VTAIL.n335 VSUBS 0.024564f
C1389 VTAIL.n336 VSUBS 0.0132f
C1390 VTAIL.n337 VSUBS 0.031199f
C1391 VTAIL.n338 VSUBS 0.013976f
C1392 VTAIL.n339 VSUBS 0.024564f
C1393 VTAIL.n340 VSUBS 0.0132f
C1394 VTAIL.n341 VSUBS 0.031199f
C1395 VTAIL.n342 VSUBS 0.013976f
C1396 VTAIL.n343 VSUBS 0.024564f
C1397 VTAIL.n344 VSUBS 0.0132f
C1398 VTAIL.n345 VSUBS 0.031199f
C1399 VTAIL.n346 VSUBS 0.013976f
C1400 VTAIL.n347 VSUBS 0.024564f
C1401 VTAIL.n348 VSUBS 0.0132f
C1402 VTAIL.n349 VSUBS 0.031199f
C1403 VTAIL.n350 VSUBS 0.013976f
C1404 VTAIL.n351 VSUBS 0.024564f
C1405 VTAIL.n352 VSUBS 0.0132f
C1406 VTAIL.n353 VSUBS 0.031199f
C1407 VTAIL.n354 VSUBS 0.031199f
C1408 VTAIL.n355 VSUBS 0.013976f
C1409 VTAIL.n356 VSUBS 0.024564f
C1410 VTAIL.n357 VSUBS 0.0132f
C1411 VTAIL.n358 VSUBS 0.031199f
C1412 VTAIL.n359 VSUBS 0.013976f
C1413 VTAIL.n360 VSUBS 0.225888f
C1414 VTAIL.t11 VSUBS 0.067471f
C1415 VTAIL.n361 VSUBS 0.0234f
C1416 VTAIL.n362 VSUBS 0.02347f
C1417 VTAIL.n363 VSUBS 0.0132f
C1418 VTAIL.n364 VSUBS 1.52121f
C1419 VTAIL.n365 VSUBS 0.024564f
C1420 VTAIL.n366 VSUBS 0.0132f
C1421 VTAIL.n367 VSUBS 0.013976f
C1422 VTAIL.n368 VSUBS 0.031199f
C1423 VTAIL.n369 VSUBS 0.031199f
C1424 VTAIL.n370 VSUBS 0.013976f
C1425 VTAIL.n371 VSUBS 0.0132f
C1426 VTAIL.n372 VSUBS 0.024564f
C1427 VTAIL.n373 VSUBS 0.024564f
C1428 VTAIL.n374 VSUBS 0.0132f
C1429 VTAIL.n375 VSUBS 0.013976f
C1430 VTAIL.n376 VSUBS 0.031199f
C1431 VTAIL.n377 VSUBS 0.031199f
C1432 VTAIL.n378 VSUBS 0.013976f
C1433 VTAIL.n379 VSUBS 0.0132f
C1434 VTAIL.n380 VSUBS 0.024564f
C1435 VTAIL.n381 VSUBS 0.024564f
C1436 VTAIL.n382 VSUBS 0.0132f
C1437 VTAIL.n383 VSUBS 0.013588f
C1438 VTAIL.n384 VSUBS 0.013588f
C1439 VTAIL.n385 VSUBS 0.031199f
C1440 VTAIL.n386 VSUBS 0.031199f
C1441 VTAIL.n387 VSUBS 0.013976f
C1442 VTAIL.n388 VSUBS 0.0132f
C1443 VTAIL.n389 VSUBS 0.024564f
C1444 VTAIL.n390 VSUBS 0.024564f
C1445 VTAIL.n391 VSUBS 0.0132f
C1446 VTAIL.n392 VSUBS 0.013976f
C1447 VTAIL.n393 VSUBS 0.031199f
C1448 VTAIL.n394 VSUBS 0.031199f
C1449 VTAIL.n395 VSUBS 0.013976f
C1450 VTAIL.n396 VSUBS 0.0132f
C1451 VTAIL.n397 VSUBS 0.024564f
C1452 VTAIL.n398 VSUBS 0.024564f
C1453 VTAIL.n399 VSUBS 0.0132f
C1454 VTAIL.n400 VSUBS 0.013976f
C1455 VTAIL.n401 VSUBS 0.031199f
C1456 VTAIL.n402 VSUBS 0.031199f
C1457 VTAIL.n403 VSUBS 0.013976f
C1458 VTAIL.n404 VSUBS 0.0132f
C1459 VTAIL.n405 VSUBS 0.024564f
C1460 VTAIL.n406 VSUBS 0.024564f
C1461 VTAIL.n407 VSUBS 0.0132f
C1462 VTAIL.n408 VSUBS 0.013976f
C1463 VTAIL.n409 VSUBS 0.031199f
C1464 VTAIL.n410 VSUBS 0.078018f
C1465 VTAIL.n411 VSUBS 0.013976f
C1466 VTAIL.n412 VSUBS 0.0132f
C1467 VTAIL.n413 VSUBS 0.054095f
C1468 VTAIL.n414 VSUBS 0.039261f
C1469 VTAIL.n415 VSUBS 0.281145f
C1470 VTAIL.n416 VSUBS 0.027721f
C1471 VTAIL.n417 VSUBS 0.024564f
C1472 VTAIL.n418 VSUBS 0.0132f
C1473 VTAIL.n419 VSUBS 0.031199f
C1474 VTAIL.n420 VSUBS 0.013976f
C1475 VTAIL.n421 VSUBS 0.024564f
C1476 VTAIL.n422 VSUBS 0.0132f
C1477 VTAIL.n423 VSUBS 0.031199f
C1478 VTAIL.n424 VSUBS 0.013976f
C1479 VTAIL.n425 VSUBS 0.024564f
C1480 VTAIL.n426 VSUBS 0.0132f
C1481 VTAIL.n427 VSUBS 0.031199f
C1482 VTAIL.n428 VSUBS 0.013976f
C1483 VTAIL.n429 VSUBS 0.024564f
C1484 VTAIL.n430 VSUBS 0.0132f
C1485 VTAIL.n431 VSUBS 0.031199f
C1486 VTAIL.n432 VSUBS 0.013976f
C1487 VTAIL.n433 VSUBS 0.024564f
C1488 VTAIL.n434 VSUBS 0.0132f
C1489 VTAIL.n435 VSUBS 0.031199f
C1490 VTAIL.n436 VSUBS 0.031199f
C1491 VTAIL.n437 VSUBS 0.013976f
C1492 VTAIL.n438 VSUBS 0.024564f
C1493 VTAIL.n439 VSUBS 0.0132f
C1494 VTAIL.n440 VSUBS 0.031199f
C1495 VTAIL.n441 VSUBS 0.013976f
C1496 VTAIL.n442 VSUBS 0.225888f
C1497 VTAIL.t5 VSUBS 0.067471f
C1498 VTAIL.n443 VSUBS 0.0234f
C1499 VTAIL.n444 VSUBS 0.02347f
C1500 VTAIL.n445 VSUBS 0.0132f
C1501 VTAIL.n446 VSUBS 1.52121f
C1502 VTAIL.n447 VSUBS 0.024564f
C1503 VTAIL.n448 VSUBS 0.0132f
C1504 VTAIL.n449 VSUBS 0.013976f
C1505 VTAIL.n450 VSUBS 0.031199f
C1506 VTAIL.n451 VSUBS 0.031199f
C1507 VTAIL.n452 VSUBS 0.013976f
C1508 VTAIL.n453 VSUBS 0.0132f
C1509 VTAIL.n454 VSUBS 0.024564f
C1510 VTAIL.n455 VSUBS 0.024564f
C1511 VTAIL.n456 VSUBS 0.0132f
C1512 VTAIL.n457 VSUBS 0.013976f
C1513 VTAIL.n458 VSUBS 0.031199f
C1514 VTAIL.n459 VSUBS 0.031199f
C1515 VTAIL.n460 VSUBS 0.013976f
C1516 VTAIL.n461 VSUBS 0.0132f
C1517 VTAIL.n462 VSUBS 0.024564f
C1518 VTAIL.n463 VSUBS 0.024564f
C1519 VTAIL.n464 VSUBS 0.0132f
C1520 VTAIL.n465 VSUBS 0.013588f
C1521 VTAIL.n466 VSUBS 0.013588f
C1522 VTAIL.n467 VSUBS 0.031199f
C1523 VTAIL.n468 VSUBS 0.031199f
C1524 VTAIL.n469 VSUBS 0.013976f
C1525 VTAIL.n470 VSUBS 0.0132f
C1526 VTAIL.n471 VSUBS 0.024564f
C1527 VTAIL.n472 VSUBS 0.024564f
C1528 VTAIL.n473 VSUBS 0.0132f
C1529 VTAIL.n474 VSUBS 0.013976f
C1530 VTAIL.n475 VSUBS 0.031199f
C1531 VTAIL.n476 VSUBS 0.031199f
C1532 VTAIL.n477 VSUBS 0.013976f
C1533 VTAIL.n478 VSUBS 0.0132f
C1534 VTAIL.n479 VSUBS 0.024564f
C1535 VTAIL.n480 VSUBS 0.024564f
C1536 VTAIL.n481 VSUBS 0.0132f
C1537 VTAIL.n482 VSUBS 0.013976f
C1538 VTAIL.n483 VSUBS 0.031199f
C1539 VTAIL.n484 VSUBS 0.031199f
C1540 VTAIL.n485 VSUBS 0.013976f
C1541 VTAIL.n486 VSUBS 0.0132f
C1542 VTAIL.n487 VSUBS 0.024564f
C1543 VTAIL.n488 VSUBS 0.024564f
C1544 VTAIL.n489 VSUBS 0.0132f
C1545 VTAIL.n490 VSUBS 0.013976f
C1546 VTAIL.n491 VSUBS 0.031199f
C1547 VTAIL.n492 VSUBS 0.078018f
C1548 VTAIL.n493 VSUBS 0.013976f
C1549 VTAIL.n494 VSUBS 0.0132f
C1550 VTAIL.n495 VSUBS 0.054095f
C1551 VTAIL.n496 VSUBS 0.039261f
C1552 VTAIL.n497 VSUBS 0.281145f
C1553 VTAIL.t1 VSUBS 0.289619f
C1554 VTAIL.t2 VSUBS 0.289619f
C1555 VTAIL.n498 VSUBS 2.17915f
C1556 VTAIL.n499 VSUBS 1.05472f
C1557 VTAIL.n500 VSUBS 0.027721f
C1558 VTAIL.n501 VSUBS 0.024564f
C1559 VTAIL.n502 VSUBS 0.0132f
C1560 VTAIL.n503 VSUBS 0.031199f
C1561 VTAIL.n504 VSUBS 0.013976f
C1562 VTAIL.n505 VSUBS 0.024564f
C1563 VTAIL.n506 VSUBS 0.0132f
C1564 VTAIL.n507 VSUBS 0.031199f
C1565 VTAIL.n508 VSUBS 0.013976f
C1566 VTAIL.n509 VSUBS 0.024564f
C1567 VTAIL.n510 VSUBS 0.0132f
C1568 VTAIL.n511 VSUBS 0.031199f
C1569 VTAIL.n512 VSUBS 0.013976f
C1570 VTAIL.n513 VSUBS 0.024564f
C1571 VTAIL.n514 VSUBS 0.0132f
C1572 VTAIL.n515 VSUBS 0.031199f
C1573 VTAIL.n516 VSUBS 0.013976f
C1574 VTAIL.n517 VSUBS 0.024564f
C1575 VTAIL.n518 VSUBS 0.0132f
C1576 VTAIL.n519 VSUBS 0.031199f
C1577 VTAIL.n520 VSUBS 0.031199f
C1578 VTAIL.n521 VSUBS 0.013976f
C1579 VTAIL.n522 VSUBS 0.024564f
C1580 VTAIL.n523 VSUBS 0.0132f
C1581 VTAIL.n524 VSUBS 0.031199f
C1582 VTAIL.n525 VSUBS 0.013976f
C1583 VTAIL.n526 VSUBS 0.225888f
C1584 VTAIL.t7 VSUBS 0.067471f
C1585 VTAIL.n527 VSUBS 0.0234f
C1586 VTAIL.n528 VSUBS 0.02347f
C1587 VTAIL.n529 VSUBS 0.0132f
C1588 VTAIL.n530 VSUBS 1.52121f
C1589 VTAIL.n531 VSUBS 0.024564f
C1590 VTAIL.n532 VSUBS 0.0132f
C1591 VTAIL.n533 VSUBS 0.013976f
C1592 VTAIL.n534 VSUBS 0.031199f
C1593 VTAIL.n535 VSUBS 0.031199f
C1594 VTAIL.n536 VSUBS 0.013976f
C1595 VTAIL.n537 VSUBS 0.0132f
C1596 VTAIL.n538 VSUBS 0.024564f
C1597 VTAIL.n539 VSUBS 0.024564f
C1598 VTAIL.n540 VSUBS 0.0132f
C1599 VTAIL.n541 VSUBS 0.013976f
C1600 VTAIL.n542 VSUBS 0.031199f
C1601 VTAIL.n543 VSUBS 0.031199f
C1602 VTAIL.n544 VSUBS 0.013976f
C1603 VTAIL.n545 VSUBS 0.0132f
C1604 VTAIL.n546 VSUBS 0.024564f
C1605 VTAIL.n547 VSUBS 0.024564f
C1606 VTAIL.n548 VSUBS 0.0132f
C1607 VTAIL.n549 VSUBS 0.013588f
C1608 VTAIL.n550 VSUBS 0.013588f
C1609 VTAIL.n551 VSUBS 0.031199f
C1610 VTAIL.n552 VSUBS 0.031199f
C1611 VTAIL.n553 VSUBS 0.013976f
C1612 VTAIL.n554 VSUBS 0.0132f
C1613 VTAIL.n555 VSUBS 0.024564f
C1614 VTAIL.n556 VSUBS 0.024564f
C1615 VTAIL.n557 VSUBS 0.0132f
C1616 VTAIL.n558 VSUBS 0.013976f
C1617 VTAIL.n559 VSUBS 0.031199f
C1618 VTAIL.n560 VSUBS 0.031199f
C1619 VTAIL.n561 VSUBS 0.013976f
C1620 VTAIL.n562 VSUBS 0.0132f
C1621 VTAIL.n563 VSUBS 0.024564f
C1622 VTAIL.n564 VSUBS 0.024564f
C1623 VTAIL.n565 VSUBS 0.0132f
C1624 VTAIL.n566 VSUBS 0.013976f
C1625 VTAIL.n567 VSUBS 0.031199f
C1626 VTAIL.n568 VSUBS 0.031199f
C1627 VTAIL.n569 VSUBS 0.013976f
C1628 VTAIL.n570 VSUBS 0.0132f
C1629 VTAIL.n571 VSUBS 0.024564f
C1630 VTAIL.n572 VSUBS 0.024564f
C1631 VTAIL.n573 VSUBS 0.0132f
C1632 VTAIL.n574 VSUBS 0.013976f
C1633 VTAIL.n575 VSUBS 0.031199f
C1634 VTAIL.n576 VSUBS 0.078018f
C1635 VTAIL.n577 VSUBS 0.013976f
C1636 VTAIL.n578 VSUBS 0.0132f
C1637 VTAIL.n579 VSUBS 0.054095f
C1638 VTAIL.n580 VSUBS 0.039261f
C1639 VTAIL.n581 VSUBS 1.82018f
C1640 VTAIL.n582 VSUBS 0.027721f
C1641 VTAIL.n583 VSUBS 0.024564f
C1642 VTAIL.n584 VSUBS 0.0132f
C1643 VTAIL.n585 VSUBS 0.031199f
C1644 VTAIL.n586 VSUBS 0.013976f
C1645 VTAIL.n587 VSUBS 0.024564f
C1646 VTAIL.n588 VSUBS 0.0132f
C1647 VTAIL.n589 VSUBS 0.031199f
C1648 VTAIL.n590 VSUBS 0.013976f
C1649 VTAIL.n591 VSUBS 0.024564f
C1650 VTAIL.n592 VSUBS 0.0132f
C1651 VTAIL.n593 VSUBS 0.031199f
C1652 VTAIL.n594 VSUBS 0.013976f
C1653 VTAIL.n595 VSUBS 0.024564f
C1654 VTAIL.n596 VSUBS 0.0132f
C1655 VTAIL.n597 VSUBS 0.031199f
C1656 VTAIL.n598 VSUBS 0.013976f
C1657 VTAIL.n599 VSUBS 0.024564f
C1658 VTAIL.n600 VSUBS 0.0132f
C1659 VTAIL.n601 VSUBS 0.031199f
C1660 VTAIL.n602 VSUBS 0.013976f
C1661 VTAIL.n603 VSUBS 0.024564f
C1662 VTAIL.n604 VSUBS 0.0132f
C1663 VTAIL.n605 VSUBS 0.031199f
C1664 VTAIL.n606 VSUBS 0.013976f
C1665 VTAIL.n607 VSUBS 0.225888f
C1666 VTAIL.t14 VSUBS 0.067471f
C1667 VTAIL.n608 VSUBS 0.0234f
C1668 VTAIL.n609 VSUBS 0.02347f
C1669 VTAIL.n610 VSUBS 0.0132f
C1670 VTAIL.n611 VSUBS 1.52121f
C1671 VTAIL.n612 VSUBS 0.024564f
C1672 VTAIL.n613 VSUBS 0.0132f
C1673 VTAIL.n614 VSUBS 0.013976f
C1674 VTAIL.n615 VSUBS 0.031199f
C1675 VTAIL.n616 VSUBS 0.031199f
C1676 VTAIL.n617 VSUBS 0.013976f
C1677 VTAIL.n618 VSUBS 0.0132f
C1678 VTAIL.n619 VSUBS 0.024564f
C1679 VTAIL.n620 VSUBS 0.024564f
C1680 VTAIL.n621 VSUBS 0.0132f
C1681 VTAIL.n622 VSUBS 0.013976f
C1682 VTAIL.n623 VSUBS 0.031199f
C1683 VTAIL.n624 VSUBS 0.031199f
C1684 VTAIL.n625 VSUBS 0.031199f
C1685 VTAIL.n626 VSUBS 0.013976f
C1686 VTAIL.n627 VSUBS 0.0132f
C1687 VTAIL.n628 VSUBS 0.024564f
C1688 VTAIL.n629 VSUBS 0.024564f
C1689 VTAIL.n630 VSUBS 0.0132f
C1690 VTAIL.n631 VSUBS 0.013588f
C1691 VTAIL.n632 VSUBS 0.013588f
C1692 VTAIL.n633 VSUBS 0.031199f
C1693 VTAIL.n634 VSUBS 0.031199f
C1694 VTAIL.n635 VSUBS 0.013976f
C1695 VTAIL.n636 VSUBS 0.0132f
C1696 VTAIL.n637 VSUBS 0.024564f
C1697 VTAIL.n638 VSUBS 0.024564f
C1698 VTAIL.n639 VSUBS 0.0132f
C1699 VTAIL.n640 VSUBS 0.013976f
C1700 VTAIL.n641 VSUBS 0.031199f
C1701 VTAIL.n642 VSUBS 0.031199f
C1702 VTAIL.n643 VSUBS 0.013976f
C1703 VTAIL.n644 VSUBS 0.0132f
C1704 VTAIL.n645 VSUBS 0.024564f
C1705 VTAIL.n646 VSUBS 0.024564f
C1706 VTAIL.n647 VSUBS 0.0132f
C1707 VTAIL.n648 VSUBS 0.013976f
C1708 VTAIL.n649 VSUBS 0.031199f
C1709 VTAIL.n650 VSUBS 0.031199f
C1710 VTAIL.n651 VSUBS 0.013976f
C1711 VTAIL.n652 VSUBS 0.0132f
C1712 VTAIL.n653 VSUBS 0.024564f
C1713 VTAIL.n654 VSUBS 0.024564f
C1714 VTAIL.n655 VSUBS 0.0132f
C1715 VTAIL.n656 VSUBS 0.013976f
C1716 VTAIL.n657 VSUBS 0.031199f
C1717 VTAIL.n658 VSUBS 0.078018f
C1718 VTAIL.n659 VSUBS 0.013976f
C1719 VTAIL.n660 VSUBS 0.0132f
C1720 VTAIL.n661 VSUBS 0.054095f
C1721 VTAIL.n662 VSUBS 0.039261f
C1722 VTAIL.n663 VSUBS 1.81557f
C1723 VDD2.t7 VSUBS 0.31914f
C1724 VDD2.t3 VSUBS 0.31914f
C1725 VDD2.n0 VSUBS 2.58661f
C1726 VDD2.t2 VSUBS 0.31914f
C1727 VDD2.t0 VSUBS 0.31914f
C1728 VDD2.n1 VSUBS 2.58661f
C1729 VDD2.n2 VSUBS 4.59198f
C1730 VDD2.t6 VSUBS 0.31914f
C1731 VDD2.t4 VSUBS 0.31914f
C1732 VDD2.n3 VSUBS 2.56904f
C1733 VDD2.n4 VSUBS 3.88283f
C1734 VDD2.t1 VSUBS 0.31914f
C1735 VDD2.t5 VSUBS 0.31914f
C1736 VDD2.n5 VSUBS 2.58657f
C1737 VN.t1 VSUBS 3.08259f
C1738 VN.n0 VSUBS 1.17543f
C1739 VN.n1 VSUBS 0.025476f
C1740 VN.n2 VSUBS 0.039852f
C1741 VN.n3 VSUBS 0.025476f
C1742 VN.t3 VSUBS 3.08259f
C1743 VN.n4 VSUBS 0.047242f
C1744 VN.n5 VSUBS 0.025476f
C1745 VN.n6 VSUBS 0.047242f
C1746 VN.t6 VSUBS 3.34073f
C1747 VN.n7 VSUBS 1.11732f
C1748 VN.t2 VSUBS 3.08259f
C1749 VN.n8 VSUBS 1.14952f
C1750 VN.n9 VSUBS 0.030684f
C1751 VN.n10 VSUBS 0.27369f
C1752 VN.n11 VSUBS 0.025476f
C1753 VN.n12 VSUBS 0.025476f
C1754 VN.n13 VSUBS 0.050366f
C1755 VN.n14 VSUBS 0.020576f
C1756 VN.n15 VSUBS 0.050366f
C1757 VN.n16 VSUBS 0.025476f
C1758 VN.n17 VSUBS 0.025476f
C1759 VN.n18 VSUBS 0.025476f
C1760 VN.n19 VSUBS 0.030684f
C1761 VN.n20 VSUBS 1.07433f
C1762 VN.n21 VSUBS 0.040479f
C1763 VN.n22 VSUBS 0.047242f
C1764 VN.n23 VSUBS 0.025476f
C1765 VN.n24 VSUBS 0.025476f
C1766 VN.n25 VSUBS 0.025476f
C1767 VN.n26 VSUBS 0.034214f
C1768 VN.n27 VSUBS 0.047242f
C1769 VN.n28 VSUBS 0.04421f
C1770 VN.n29 VSUBS 0.041111f
C1771 VN.n30 VSUBS 0.051144f
C1772 VN.t7 VSUBS 3.08259f
C1773 VN.n31 VSUBS 1.17543f
C1774 VN.n32 VSUBS 0.025476f
C1775 VN.n33 VSUBS 0.039852f
C1776 VN.n34 VSUBS 0.025476f
C1777 VN.t5 VSUBS 3.08259f
C1778 VN.n35 VSUBS 0.047242f
C1779 VN.n36 VSUBS 0.025476f
C1780 VN.n37 VSUBS 0.047242f
C1781 VN.t4 VSUBS 3.34073f
C1782 VN.n38 VSUBS 1.11732f
C1783 VN.t0 VSUBS 3.08259f
C1784 VN.n39 VSUBS 1.14952f
C1785 VN.n40 VSUBS 0.030684f
C1786 VN.n41 VSUBS 0.27369f
C1787 VN.n42 VSUBS 0.025476f
C1788 VN.n43 VSUBS 0.025476f
C1789 VN.n44 VSUBS 0.050366f
C1790 VN.n45 VSUBS 0.020576f
C1791 VN.n46 VSUBS 0.050366f
C1792 VN.n47 VSUBS 0.025476f
C1793 VN.n48 VSUBS 0.025476f
C1794 VN.n49 VSUBS 0.025476f
C1795 VN.n50 VSUBS 0.030684f
C1796 VN.n51 VSUBS 1.07433f
C1797 VN.n52 VSUBS 0.040479f
C1798 VN.n53 VSUBS 0.047242f
C1799 VN.n54 VSUBS 0.025476f
C1800 VN.n55 VSUBS 0.025476f
C1801 VN.n56 VSUBS 0.025476f
C1802 VN.n57 VSUBS 0.034214f
C1803 VN.n58 VSUBS 0.047242f
C1804 VN.n59 VSUBS 0.04421f
C1805 VN.n60 VSUBS 0.041111f
C1806 VN.n61 VSUBS 1.65329f
.ends

