* NGSPICE file created from diff_pair_sample_0078.ext - technology: sky130A

.subckt diff_pair_sample_0078 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t7 VP.t0 VTAIL.t13 w_n4360_n1490# sky130_fd_pr__pfet_01v8 ad=0.43065 pd=2.94 as=0.43065 ps=2.94 w=2.61 l=3.06
X1 VTAIL.t7 VN.t0 VDD2.t7 w_n4360_n1490# sky130_fd_pr__pfet_01v8 ad=0.43065 pd=2.94 as=0.43065 ps=2.94 w=2.61 l=3.06
X2 VTAIL.t2 VN.t1 VDD2.t6 w_n4360_n1490# sky130_fd_pr__pfet_01v8 ad=1.0179 pd=6 as=0.43065 ps=2.94 w=2.61 l=3.06
X3 VTAIL.t0 VN.t2 VDD2.t5 w_n4360_n1490# sky130_fd_pr__pfet_01v8 ad=1.0179 pd=6 as=0.43065 ps=2.94 w=2.61 l=3.06
X4 VDD1.t6 VP.t1 VTAIL.t12 w_n4360_n1490# sky130_fd_pr__pfet_01v8 ad=0.43065 pd=2.94 as=1.0179 ps=6 w=2.61 l=3.06
X5 VDD1.t5 VP.t2 VTAIL.t9 w_n4360_n1490# sky130_fd_pr__pfet_01v8 ad=0.43065 pd=2.94 as=1.0179 ps=6 w=2.61 l=3.06
X6 VDD2.t4 VN.t3 VTAIL.t4 w_n4360_n1490# sky130_fd_pr__pfet_01v8 ad=0.43065 pd=2.94 as=1.0179 ps=6 w=2.61 l=3.06
X7 VDD2.t3 VN.t4 VTAIL.t5 w_n4360_n1490# sky130_fd_pr__pfet_01v8 ad=0.43065 pd=2.94 as=0.43065 ps=2.94 w=2.61 l=3.06
X8 VTAIL.t11 VP.t3 VDD1.t4 w_n4360_n1490# sky130_fd_pr__pfet_01v8 ad=0.43065 pd=2.94 as=0.43065 ps=2.94 w=2.61 l=3.06
X9 VTAIL.t6 VN.t5 VDD2.t2 w_n4360_n1490# sky130_fd_pr__pfet_01v8 ad=0.43065 pd=2.94 as=0.43065 ps=2.94 w=2.61 l=3.06
X10 B.t11 B.t9 B.t10 w_n4360_n1490# sky130_fd_pr__pfet_01v8 ad=1.0179 pd=6 as=0 ps=0 w=2.61 l=3.06
X11 B.t8 B.t6 B.t7 w_n4360_n1490# sky130_fd_pr__pfet_01v8 ad=1.0179 pd=6 as=0 ps=0 w=2.61 l=3.06
X12 VDD1.t3 VP.t4 VTAIL.t15 w_n4360_n1490# sky130_fd_pr__pfet_01v8 ad=0.43065 pd=2.94 as=0.43065 ps=2.94 w=2.61 l=3.06
X13 VDD2.t1 VN.t6 VTAIL.t1 w_n4360_n1490# sky130_fd_pr__pfet_01v8 ad=0.43065 pd=2.94 as=0.43065 ps=2.94 w=2.61 l=3.06
X14 VTAIL.t8 VP.t5 VDD1.t2 w_n4360_n1490# sky130_fd_pr__pfet_01v8 ad=1.0179 pd=6 as=0.43065 ps=2.94 w=2.61 l=3.06
X15 VTAIL.t14 VP.t6 VDD1.t1 w_n4360_n1490# sky130_fd_pr__pfet_01v8 ad=0.43065 pd=2.94 as=0.43065 ps=2.94 w=2.61 l=3.06
X16 VDD2.t0 VN.t7 VTAIL.t3 w_n4360_n1490# sky130_fd_pr__pfet_01v8 ad=0.43065 pd=2.94 as=1.0179 ps=6 w=2.61 l=3.06
X17 VTAIL.t10 VP.t7 VDD1.t0 w_n4360_n1490# sky130_fd_pr__pfet_01v8 ad=1.0179 pd=6 as=0.43065 ps=2.94 w=2.61 l=3.06
X18 B.t5 B.t3 B.t4 w_n4360_n1490# sky130_fd_pr__pfet_01v8 ad=1.0179 pd=6 as=0 ps=0 w=2.61 l=3.06
X19 B.t2 B.t0 B.t1 w_n4360_n1490# sky130_fd_pr__pfet_01v8 ad=1.0179 pd=6 as=0 ps=0 w=2.61 l=3.06
R0 VP.n21 VP.n18 161.3
R1 VP.n23 VP.n22 161.3
R2 VP.n24 VP.n17 161.3
R3 VP.n26 VP.n25 161.3
R4 VP.n27 VP.n16 161.3
R5 VP.n29 VP.n28 161.3
R6 VP.n31 VP.n30 161.3
R7 VP.n32 VP.n14 161.3
R8 VP.n34 VP.n33 161.3
R9 VP.n35 VP.n13 161.3
R10 VP.n37 VP.n36 161.3
R11 VP.n38 VP.n12 161.3
R12 VP.n40 VP.n39 161.3
R13 VP.n75 VP.n74 161.3
R14 VP.n73 VP.n1 161.3
R15 VP.n72 VP.n71 161.3
R16 VP.n70 VP.n2 161.3
R17 VP.n69 VP.n68 161.3
R18 VP.n67 VP.n3 161.3
R19 VP.n66 VP.n65 161.3
R20 VP.n64 VP.n63 161.3
R21 VP.n62 VP.n5 161.3
R22 VP.n61 VP.n60 161.3
R23 VP.n59 VP.n6 161.3
R24 VP.n58 VP.n57 161.3
R25 VP.n56 VP.n7 161.3
R26 VP.n54 VP.n53 161.3
R27 VP.n52 VP.n8 161.3
R28 VP.n51 VP.n50 161.3
R29 VP.n49 VP.n9 161.3
R30 VP.n48 VP.n47 161.3
R31 VP.n46 VP.n10 161.3
R32 VP.n45 VP.n44 161.3
R33 VP.n43 VP.n42 73.6745
R34 VP.n76 VP.n0 73.6745
R35 VP.n41 VP.n11 73.6745
R36 VP.n61 VP.n6 56.5193
R37 VP.n26 VP.n17 56.5193
R38 VP.n49 VP.n48 54.0911
R39 VP.n72 VP.n2 54.0911
R40 VP.n37 VP.n13 54.0911
R41 VP.n19 VP.t5 53.7686
R42 VP.n20 VP.n19 52.0468
R43 VP.n42 VP.n41 46.0145
R44 VP.n50 VP.n49 26.8957
R45 VP.n68 VP.n2 26.8957
R46 VP.n33 VP.n13 26.8957
R47 VP.n44 VP.n10 24.4675
R48 VP.n48 VP.n10 24.4675
R49 VP.n50 VP.n8 24.4675
R50 VP.n54 VP.n8 24.4675
R51 VP.n57 VP.n56 24.4675
R52 VP.n57 VP.n6 24.4675
R53 VP.n62 VP.n61 24.4675
R54 VP.n63 VP.n62 24.4675
R55 VP.n67 VP.n66 24.4675
R56 VP.n68 VP.n67 24.4675
R57 VP.n73 VP.n72 24.4675
R58 VP.n74 VP.n73 24.4675
R59 VP.n38 VP.n37 24.4675
R60 VP.n39 VP.n38 24.4675
R61 VP.n27 VP.n26 24.4675
R62 VP.n28 VP.n27 24.4675
R63 VP.n32 VP.n31 24.4675
R64 VP.n33 VP.n32 24.4675
R65 VP.n22 VP.n21 24.4675
R66 VP.n22 VP.n17 24.4675
R67 VP.n56 VP.n55 21.7761
R68 VP.n63 VP.n4 21.7761
R69 VP.n28 VP.n15 21.7761
R70 VP.n21 VP.n20 21.7761
R71 VP.n43 VP.t7 20.5564
R72 VP.n55 VP.t0 20.5564
R73 VP.n4 VP.t6 20.5564
R74 VP.n0 VP.t1 20.5564
R75 VP.n11 VP.t2 20.5564
R76 VP.n15 VP.t3 20.5564
R77 VP.n20 VP.t4 20.5564
R78 VP.n44 VP.n43 16.3934
R79 VP.n74 VP.n0 16.3934
R80 VP.n39 VP.n11 16.3934
R81 VP.n19 VP.n18 4.0838
R82 VP.n55 VP.n54 2.69187
R83 VP.n66 VP.n4 2.69187
R84 VP.n31 VP.n15 2.69187
R85 VP.n41 VP.n40 0.354971
R86 VP.n45 VP.n42 0.354971
R87 VP.n76 VP.n75 0.354971
R88 VP VP.n76 0.26696
R89 VP.n23 VP.n18 0.189894
R90 VP.n24 VP.n23 0.189894
R91 VP.n25 VP.n24 0.189894
R92 VP.n25 VP.n16 0.189894
R93 VP.n29 VP.n16 0.189894
R94 VP.n30 VP.n29 0.189894
R95 VP.n30 VP.n14 0.189894
R96 VP.n34 VP.n14 0.189894
R97 VP.n35 VP.n34 0.189894
R98 VP.n36 VP.n35 0.189894
R99 VP.n36 VP.n12 0.189894
R100 VP.n40 VP.n12 0.189894
R101 VP.n46 VP.n45 0.189894
R102 VP.n47 VP.n46 0.189894
R103 VP.n47 VP.n9 0.189894
R104 VP.n51 VP.n9 0.189894
R105 VP.n52 VP.n51 0.189894
R106 VP.n53 VP.n52 0.189894
R107 VP.n53 VP.n7 0.189894
R108 VP.n58 VP.n7 0.189894
R109 VP.n59 VP.n58 0.189894
R110 VP.n60 VP.n59 0.189894
R111 VP.n60 VP.n5 0.189894
R112 VP.n64 VP.n5 0.189894
R113 VP.n65 VP.n64 0.189894
R114 VP.n65 VP.n3 0.189894
R115 VP.n69 VP.n3 0.189894
R116 VP.n70 VP.n69 0.189894
R117 VP.n71 VP.n70 0.189894
R118 VP.n71 VP.n1 0.189894
R119 VP.n75 VP.n1 0.189894
R120 VTAIL.n98 VTAIL.n92 756.745
R121 VTAIL.n8 VTAIL.n2 756.745
R122 VTAIL.n20 VTAIL.n14 756.745
R123 VTAIL.n34 VTAIL.n28 756.745
R124 VTAIL.n86 VTAIL.n80 756.745
R125 VTAIL.n72 VTAIL.n66 756.745
R126 VTAIL.n60 VTAIL.n54 756.745
R127 VTAIL.n46 VTAIL.n40 756.745
R128 VTAIL.n97 VTAIL.n96 585
R129 VTAIL.n99 VTAIL.n98 585
R130 VTAIL.n7 VTAIL.n6 585
R131 VTAIL.n9 VTAIL.n8 585
R132 VTAIL.n19 VTAIL.n18 585
R133 VTAIL.n21 VTAIL.n20 585
R134 VTAIL.n33 VTAIL.n32 585
R135 VTAIL.n35 VTAIL.n34 585
R136 VTAIL.n87 VTAIL.n86 585
R137 VTAIL.n85 VTAIL.n84 585
R138 VTAIL.n73 VTAIL.n72 585
R139 VTAIL.n71 VTAIL.n70 585
R140 VTAIL.n61 VTAIL.n60 585
R141 VTAIL.n59 VTAIL.n58 585
R142 VTAIL.n47 VTAIL.n46 585
R143 VTAIL.n45 VTAIL.n44 585
R144 VTAIL.n95 VTAIL.t3 355.474
R145 VTAIL.n5 VTAIL.t2 355.474
R146 VTAIL.n17 VTAIL.t12 355.474
R147 VTAIL.n31 VTAIL.t10 355.474
R148 VTAIL.n83 VTAIL.t9 355.474
R149 VTAIL.n69 VTAIL.t8 355.474
R150 VTAIL.n57 VTAIL.t4 355.474
R151 VTAIL.n43 VTAIL.t0 355.474
R152 VTAIL.n98 VTAIL.n97 171.744
R153 VTAIL.n8 VTAIL.n7 171.744
R154 VTAIL.n20 VTAIL.n19 171.744
R155 VTAIL.n34 VTAIL.n33 171.744
R156 VTAIL.n86 VTAIL.n85 171.744
R157 VTAIL.n72 VTAIL.n71 171.744
R158 VTAIL.n60 VTAIL.n59 171.744
R159 VTAIL.n46 VTAIL.n45 171.744
R160 VTAIL.n79 VTAIL.n78 139.114
R161 VTAIL.n53 VTAIL.n52 139.114
R162 VTAIL.n1 VTAIL.n0 139.114
R163 VTAIL.n27 VTAIL.n26 139.114
R164 VTAIL.n97 VTAIL.t3 85.8723
R165 VTAIL.n7 VTAIL.t2 85.8723
R166 VTAIL.n19 VTAIL.t12 85.8723
R167 VTAIL.n33 VTAIL.t10 85.8723
R168 VTAIL.n85 VTAIL.t9 85.8723
R169 VTAIL.n71 VTAIL.t8 85.8723
R170 VTAIL.n59 VTAIL.t4 85.8723
R171 VTAIL.n45 VTAIL.t0 85.8723
R172 VTAIL.n103 VTAIL.n102 36.2581
R173 VTAIL.n13 VTAIL.n12 36.2581
R174 VTAIL.n25 VTAIL.n24 36.2581
R175 VTAIL.n39 VTAIL.n38 36.2581
R176 VTAIL.n91 VTAIL.n90 36.2581
R177 VTAIL.n77 VTAIL.n76 36.2581
R178 VTAIL.n65 VTAIL.n64 36.2581
R179 VTAIL.n51 VTAIL.n50 36.2581
R180 VTAIL.n103 VTAIL.n91 17.5393
R181 VTAIL.n51 VTAIL.n39 17.5393
R182 VTAIL.n96 VTAIL.n95 15.8418
R183 VTAIL.n6 VTAIL.n5 15.8418
R184 VTAIL.n18 VTAIL.n17 15.8418
R185 VTAIL.n32 VTAIL.n31 15.8418
R186 VTAIL.n84 VTAIL.n83 15.8418
R187 VTAIL.n70 VTAIL.n69 15.8418
R188 VTAIL.n58 VTAIL.n57 15.8418
R189 VTAIL.n44 VTAIL.n43 15.8418
R190 VTAIL.n99 VTAIL.n94 12.8005
R191 VTAIL.n9 VTAIL.n4 12.8005
R192 VTAIL.n21 VTAIL.n16 12.8005
R193 VTAIL.n35 VTAIL.n30 12.8005
R194 VTAIL.n87 VTAIL.n82 12.8005
R195 VTAIL.n73 VTAIL.n68 12.8005
R196 VTAIL.n61 VTAIL.n56 12.8005
R197 VTAIL.n47 VTAIL.n42 12.8005
R198 VTAIL.n0 VTAIL.t1 12.4545
R199 VTAIL.n0 VTAIL.t7 12.4545
R200 VTAIL.n26 VTAIL.t13 12.4545
R201 VTAIL.n26 VTAIL.t14 12.4545
R202 VTAIL.n78 VTAIL.t15 12.4545
R203 VTAIL.n78 VTAIL.t11 12.4545
R204 VTAIL.n52 VTAIL.t5 12.4545
R205 VTAIL.n52 VTAIL.t6 12.4545
R206 VTAIL.n100 VTAIL.n92 12.0247
R207 VTAIL.n10 VTAIL.n2 12.0247
R208 VTAIL.n22 VTAIL.n14 12.0247
R209 VTAIL.n36 VTAIL.n28 12.0247
R210 VTAIL.n88 VTAIL.n80 12.0247
R211 VTAIL.n74 VTAIL.n66 12.0247
R212 VTAIL.n62 VTAIL.n54 12.0247
R213 VTAIL.n48 VTAIL.n40 12.0247
R214 VTAIL.n102 VTAIL.n101 9.45567
R215 VTAIL.n12 VTAIL.n11 9.45567
R216 VTAIL.n24 VTAIL.n23 9.45567
R217 VTAIL.n38 VTAIL.n37 9.45567
R218 VTAIL.n90 VTAIL.n89 9.45567
R219 VTAIL.n76 VTAIL.n75 9.45567
R220 VTAIL.n64 VTAIL.n63 9.45567
R221 VTAIL.n50 VTAIL.n49 9.45567
R222 VTAIL.n101 VTAIL.n100 9.3005
R223 VTAIL.n94 VTAIL.n93 9.3005
R224 VTAIL.n11 VTAIL.n10 9.3005
R225 VTAIL.n4 VTAIL.n3 9.3005
R226 VTAIL.n23 VTAIL.n22 9.3005
R227 VTAIL.n16 VTAIL.n15 9.3005
R228 VTAIL.n37 VTAIL.n36 9.3005
R229 VTAIL.n30 VTAIL.n29 9.3005
R230 VTAIL.n89 VTAIL.n88 9.3005
R231 VTAIL.n82 VTAIL.n81 9.3005
R232 VTAIL.n75 VTAIL.n74 9.3005
R233 VTAIL.n68 VTAIL.n67 9.3005
R234 VTAIL.n63 VTAIL.n62 9.3005
R235 VTAIL.n56 VTAIL.n55 9.3005
R236 VTAIL.n49 VTAIL.n48 9.3005
R237 VTAIL.n42 VTAIL.n41 9.3005
R238 VTAIL.n83 VTAIL.n81 4.29255
R239 VTAIL.n69 VTAIL.n67 4.29255
R240 VTAIL.n57 VTAIL.n55 4.29255
R241 VTAIL.n43 VTAIL.n41 4.29255
R242 VTAIL.n95 VTAIL.n93 4.29255
R243 VTAIL.n5 VTAIL.n3 4.29255
R244 VTAIL.n17 VTAIL.n15 4.29255
R245 VTAIL.n31 VTAIL.n29 4.29255
R246 VTAIL.n53 VTAIL.n51 2.92291
R247 VTAIL.n65 VTAIL.n53 2.92291
R248 VTAIL.n79 VTAIL.n77 2.92291
R249 VTAIL.n91 VTAIL.n79 2.92291
R250 VTAIL.n39 VTAIL.n27 2.92291
R251 VTAIL.n27 VTAIL.n25 2.92291
R252 VTAIL.n13 VTAIL.n1 2.92291
R253 VTAIL VTAIL.n103 2.86472
R254 VTAIL.n102 VTAIL.n92 1.93989
R255 VTAIL.n12 VTAIL.n2 1.93989
R256 VTAIL.n24 VTAIL.n14 1.93989
R257 VTAIL.n38 VTAIL.n28 1.93989
R258 VTAIL.n90 VTAIL.n80 1.93989
R259 VTAIL.n76 VTAIL.n66 1.93989
R260 VTAIL.n64 VTAIL.n54 1.93989
R261 VTAIL.n50 VTAIL.n40 1.93989
R262 VTAIL.n100 VTAIL.n99 1.16414
R263 VTAIL.n10 VTAIL.n9 1.16414
R264 VTAIL.n22 VTAIL.n21 1.16414
R265 VTAIL.n36 VTAIL.n35 1.16414
R266 VTAIL.n88 VTAIL.n87 1.16414
R267 VTAIL.n74 VTAIL.n73 1.16414
R268 VTAIL.n62 VTAIL.n61 1.16414
R269 VTAIL.n48 VTAIL.n47 1.16414
R270 VTAIL.n77 VTAIL.n65 0.470328
R271 VTAIL.n25 VTAIL.n13 0.470328
R272 VTAIL.n96 VTAIL.n94 0.388379
R273 VTAIL.n6 VTAIL.n4 0.388379
R274 VTAIL.n18 VTAIL.n16 0.388379
R275 VTAIL.n32 VTAIL.n30 0.388379
R276 VTAIL.n84 VTAIL.n82 0.388379
R277 VTAIL.n70 VTAIL.n68 0.388379
R278 VTAIL.n58 VTAIL.n56 0.388379
R279 VTAIL.n44 VTAIL.n42 0.388379
R280 VTAIL.n101 VTAIL.n93 0.155672
R281 VTAIL.n11 VTAIL.n3 0.155672
R282 VTAIL.n23 VTAIL.n15 0.155672
R283 VTAIL.n37 VTAIL.n29 0.155672
R284 VTAIL.n89 VTAIL.n81 0.155672
R285 VTAIL.n75 VTAIL.n67 0.155672
R286 VTAIL.n63 VTAIL.n55 0.155672
R287 VTAIL.n49 VTAIL.n41 0.155672
R288 VTAIL VTAIL.n1 0.0586897
R289 VDD1 VDD1.n0 157.312
R290 VDD1.n3 VDD1.n2 157.198
R291 VDD1.n3 VDD1.n1 157.198
R292 VDD1.n5 VDD1.n4 155.792
R293 VDD1.n5 VDD1.n3 39.6992
R294 VDD1.n4 VDD1.t4 12.4545
R295 VDD1.n4 VDD1.t5 12.4545
R296 VDD1.n0 VDD1.t2 12.4545
R297 VDD1.n0 VDD1.t3 12.4545
R298 VDD1.n2 VDD1.t1 12.4545
R299 VDD1.n2 VDD1.t6 12.4545
R300 VDD1.n1 VDD1.t0 12.4545
R301 VDD1.n1 VDD1.t7 12.4545
R302 VDD1 VDD1.n5 1.40352
R303 VN.n60 VN.n59 161.3
R304 VN.n58 VN.n32 161.3
R305 VN.n57 VN.n56 161.3
R306 VN.n55 VN.n33 161.3
R307 VN.n54 VN.n53 161.3
R308 VN.n52 VN.n34 161.3
R309 VN.n51 VN.n50 161.3
R310 VN.n49 VN.n48 161.3
R311 VN.n47 VN.n36 161.3
R312 VN.n46 VN.n45 161.3
R313 VN.n44 VN.n37 161.3
R314 VN.n43 VN.n42 161.3
R315 VN.n41 VN.n38 161.3
R316 VN.n29 VN.n28 161.3
R317 VN.n27 VN.n1 161.3
R318 VN.n26 VN.n25 161.3
R319 VN.n24 VN.n2 161.3
R320 VN.n23 VN.n22 161.3
R321 VN.n21 VN.n3 161.3
R322 VN.n20 VN.n19 161.3
R323 VN.n18 VN.n17 161.3
R324 VN.n16 VN.n5 161.3
R325 VN.n15 VN.n14 161.3
R326 VN.n13 VN.n6 161.3
R327 VN.n12 VN.n11 161.3
R328 VN.n10 VN.n7 161.3
R329 VN.n30 VN.n0 73.6745
R330 VN.n61 VN.n31 73.6745
R331 VN.n15 VN.n6 56.5193
R332 VN.n46 VN.n37 56.5193
R333 VN.n26 VN.n2 54.0911
R334 VN.n57 VN.n33 54.0911
R335 VN.n39 VN.t3 53.7689
R336 VN.n8 VN.t1 53.7689
R337 VN.n9 VN.n8 52.0467
R338 VN.n40 VN.n39 52.0467
R339 VN VN.n61 46.1798
R340 VN.n22 VN.n2 26.8957
R341 VN.n53 VN.n33 26.8957
R342 VN.n11 VN.n10 24.4675
R343 VN.n11 VN.n6 24.4675
R344 VN.n16 VN.n15 24.4675
R345 VN.n17 VN.n16 24.4675
R346 VN.n21 VN.n20 24.4675
R347 VN.n22 VN.n21 24.4675
R348 VN.n27 VN.n26 24.4675
R349 VN.n28 VN.n27 24.4675
R350 VN.n42 VN.n37 24.4675
R351 VN.n42 VN.n41 24.4675
R352 VN.n53 VN.n52 24.4675
R353 VN.n52 VN.n51 24.4675
R354 VN.n48 VN.n47 24.4675
R355 VN.n47 VN.n46 24.4675
R356 VN.n59 VN.n58 24.4675
R357 VN.n58 VN.n57 24.4675
R358 VN.n10 VN.n9 21.7761
R359 VN.n17 VN.n4 21.7761
R360 VN.n41 VN.n40 21.7761
R361 VN.n48 VN.n35 21.7761
R362 VN.n9 VN.t6 20.5564
R363 VN.n4 VN.t0 20.5564
R364 VN.n0 VN.t7 20.5564
R365 VN.n40 VN.t5 20.5564
R366 VN.n35 VN.t4 20.5564
R367 VN.n31 VN.t2 20.5564
R368 VN.n28 VN.n0 16.3934
R369 VN.n59 VN.n31 16.3934
R370 VN.n39 VN.n38 4.08382
R371 VN.n8 VN.n7 4.08382
R372 VN.n20 VN.n4 2.69187
R373 VN.n51 VN.n35 2.69187
R374 VN.n61 VN.n60 0.354971
R375 VN.n30 VN.n29 0.354971
R376 VN VN.n30 0.26696
R377 VN.n60 VN.n32 0.189894
R378 VN.n56 VN.n32 0.189894
R379 VN.n56 VN.n55 0.189894
R380 VN.n55 VN.n54 0.189894
R381 VN.n54 VN.n34 0.189894
R382 VN.n50 VN.n34 0.189894
R383 VN.n50 VN.n49 0.189894
R384 VN.n49 VN.n36 0.189894
R385 VN.n45 VN.n36 0.189894
R386 VN.n45 VN.n44 0.189894
R387 VN.n44 VN.n43 0.189894
R388 VN.n43 VN.n38 0.189894
R389 VN.n12 VN.n7 0.189894
R390 VN.n13 VN.n12 0.189894
R391 VN.n14 VN.n13 0.189894
R392 VN.n14 VN.n5 0.189894
R393 VN.n18 VN.n5 0.189894
R394 VN.n19 VN.n18 0.189894
R395 VN.n19 VN.n3 0.189894
R396 VN.n23 VN.n3 0.189894
R397 VN.n24 VN.n23 0.189894
R398 VN.n25 VN.n24 0.189894
R399 VN.n25 VN.n1 0.189894
R400 VN.n29 VN.n1 0.189894
R401 VDD2.n2 VDD2.n1 157.198
R402 VDD2.n2 VDD2.n0 157.198
R403 VDD2 VDD2.n5 157.196
R404 VDD2.n4 VDD2.n3 155.793
R405 VDD2.n4 VDD2.n2 39.1162
R406 VDD2.n5 VDD2.t2 12.4545
R407 VDD2.n5 VDD2.t4 12.4545
R408 VDD2.n3 VDD2.t5 12.4545
R409 VDD2.n3 VDD2.t3 12.4545
R410 VDD2.n1 VDD2.t7 12.4545
R411 VDD2.n1 VDD2.t0 12.4545
R412 VDD2.n0 VDD2.t6 12.4545
R413 VDD2.n0 VDD2.t1 12.4545
R414 VDD2 VDD2.n4 1.5199
R415 B.n485 B.n54 585
R416 B.n487 B.n486 585
R417 B.n488 B.n53 585
R418 B.n490 B.n489 585
R419 B.n491 B.n52 585
R420 B.n493 B.n492 585
R421 B.n494 B.n51 585
R422 B.n496 B.n495 585
R423 B.n497 B.n50 585
R424 B.n499 B.n498 585
R425 B.n500 B.n49 585
R426 B.n502 B.n501 585
R427 B.n503 B.n48 585
R428 B.n505 B.n504 585
R429 B.n507 B.n45 585
R430 B.n509 B.n508 585
R431 B.n510 B.n44 585
R432 B.n512 B.n511 585
R433 B.n513 B.n43 585
R434 B.n515 B.n514 585
R435 B.n516 B.n42 585
R436 B.n518 B.n517 585
R437 B.n519 B.n41 585
R438 B.n521 B.n520 585
R439 B.n523 B.n522 585
R440 B.n524 B.n37 585
R441 B.n526 B.n525 585
R442 B.n527 B.n36 585
R443 B.n529 B.n528 585
R444 B.n530 B.n35 585
R445 B.n532 B.n531 585
R446 B.n533 B.n34 585
R447 B.n535 B.n534 585
R448 B.n536 B.n33 585
R449 B.n538 B.n537 585
R450 B.n539 B.n32 585
R451 B.n541 B.n540 585
R452 B.n542 B.n31 585
R453 B.n484 B.n483 585
R454 B.n482 B.n55 585
R455 B.n481 B.n480 585
R456 B.n479 B.n56 585
R457 B.n478 B.n477 585
R458 B.n476 B.n57 585
R459 B.n475 B.n474 585
R460 B.n473 B.n58 585
R461 B.n472 B.n471 585
R462 B.n470 B.n59 585
R463 B.n469 B.n468 585
R464 B.n467 B.n60 585
R465 B.n466 B.n465 585
R466 B.n464 B.n61 585
R467 B.n463 B.n462 585
R468 B.n461 B.n62 585
R469 B.n460 B.n459 585
R470 B.n458 B.n63 585
R471 B.n457 B.n456 585
R472 B.n455 B.n64 585
R473 B.n454 B.n453 585
R474 B.n452 B.n65 585
R475 B.n451 B.n450 585
R476 B.n449 B.n66 585
R477 B.n448 B.n447 585
R478 B.n446 B.n67 585
R479 B.n445 B.n444 585
R480 B.n443 B.n68 585
R481 B.n442 B.n441 585
R482 B.n440 B.n69 585
R483 B.n439 B.n438 585
R484 B.n437 B.n70 585
R485 B.n436 B.n435 585
R486 B.n434 B.n71 585
R487 B.n433 B.n432 585
R488 B.n431 B.n72 585
R489 B.n430 B.n429 585
R490 B.n428 B.n73 585
R491 B.n427 B.n426 585
R492 B.n425 B.n74 585
R493 B.n424 B.n423 585
R494 B.n422 B.n75 585
R495 B.n421 B.n420 585
R496 B.n419 B.n76 585
R497 B.n418 B.n417 585
R498 B.n416 B.n77 585
R499 B.n415 B.n414 585
R500 B.n413 B.n78 585
R501 B.n412 B.n411 585
R502 B.n410 B.n79 585
R503 B.n409 B.n408 585
R504 B.n407 B.n80 585
R505 B.n406 B.n405 585
R506 B.n404 B.n81 585
R507 B.n403 B.n402 585
R508 B.n401 B.n82 585
R509 B.n400 B.n399 585
R510 B.n398 B.n83 585
R511 B.n397 B.n396 585
R512 B.n395 B.n84 585
R513 B.n394 B.n393 585
R514 B.n392 B.n85 585
R515 B.n391 B.n390 585
R516 B.n389 B.n86 585
R517 B.n388 B.n387 585
R518 B.n386 B.n87 585
R519 B.n385 B.n384 585
R520 B.n383 B.n88 585
R521 B.n382 B.n381 585
R522 B.n380 B.n89 585
R523 B.n379 B.n378 585
R524 B.n377 B.n90 585
R525 B.n376 B.n375 585
R526 B.n374 B.n91 585
R527 B.n373 B.n372 585
R528 B.n371 B.n92 585
R529 B.n370 B.n369 585
R530 B.n368 B.n93 585
R531 B.n367 B.n366 585
R532 B.n365 B.n94 585
R533 B.n364 B.n363 585
R534 B.n362 B.n95 585
R535 B.n361 B.n360 585
R536 B.n359 B.n96 585
R537 B.n358 B.n357 585
R538 B.n356 B.n97 585
R539 B.n355 B.n354 585
R540 B.n353 B.n98 585
R541 B.n352 B.n351 585
R542 B.n350 B.n99 585
R543 B.n349 B.n348 585
R544 B.n347 B.n100 585
R545 B.n346 B.n345 585
R546 B.n344 B.n101 585
R547 B.n343 B.n342 585
R548 B.n341 B.n102 585
R549 B.n340 B.n339 585
R550 B.n338 B.n103 585
R551 B.n337 B.n336 585
R552 B.n335 B.n104 585
R553 B.n334 B.n333 585
R554 B.n332 B.n105 585
R555 B.n331 B.n330 585
R556 B.n329 B.n106 585
R557 B.n328 B.n327 585
R558 B.n326 B.n107 585
R559 B.n325 B.n324 585
R560 B.n323 B.n108 585
R561 B.n322 B.n321 585
R562 B.n320 B.n109 585
R563 B.n319 B.n318 585
R564 B.n317 B.n110 585
R565 B.n316 B.n315 585
R566 B.n314 B.n111 585
R567 B.n313 B.n312 585
R568 B.n311 B.n112 585
R569 B.n310 B.n309 585
R570 B.n251 B.n136 585
R571 B.n253 B.n252 585
R572 B.n254 B.n135 585
R573 B.n256 B.n255 585
R574 B.n257 B.n134 585
R575 B.n259 B.n258 585
R576 B.n260 B.n133 585
R577 B.n262 B.n261 585
R578 B.n263 B.n132 585
R579 B.n265 B.n264 585
R580 B.n266 B.n131 585
R581 B.n268 B.n267 585
R582 B.n269 B.n130 585
R583 B.n271 B.n270 585
R584 B.n273 B.n127 585
R585 B.n275 B.n274 585
R586 B.n276 B.n126 585
R587 B.n278 B.n277 585
R588 B.n279 B.n125 585
R589 B.n281 B.n280 585
R590 B.n282 B.n124 585
R591 B.n284 B.n283 585
R592 B.n285 B.n123 585
R593 B.n287 B.n286 585
R594 B.n289 B.n288 585
R595 B.n290 B.n119 585
R596 B.n292 B.n291 585
R597 B.n293 B.n118 585
R598 B.n295 B.n294 585
R599 B.n296 B.n117 585
R600 B.n298 B.n297 585
R601 B.n299 B.n116 585
R602 B.n301 B.n300 585
R603 B.n302 B.n115 585
R604 B.n304 B.n303 585
R605 B.n305 B.n114 585
R606 B.n307 B.n306 585
R607 B.n308 B.n113 585
R608 B.n250 B.n249 585
R609 B.n248 B.n137 585
R610 B.n247 B.n246 585
R611 B.n245 B.n138 585
R612 B.n244 B.n243 585
R613 B.n242 B.n139 585
R614 B.n241 B.n240 585
R615 B.n239 B.n140 585
R616 B.n238 B.n237 585
R617 B.n236 B.n141 585
R618 B.n235 B.n234 585
R619 B.n233 B.n142 585
R620 B.n232 B.n231 585
R621 B.n230 B.n143 585
R622 B.n229 B.n228 585
R623 B.n227 B.n144 585
R624 B.n226 B.n225 585
R625 B.n224 B.n145 585
R626 B.n223 B.n222 585
R627 B.n221 B.n146 585
R628 B.n220 B.n219 585
R629 B.n218 B.n147 585
R630 B.n217 B.n216 585
R631 B.n215 B.n148 585
R632 B.n214 B.n213 585
R633 B.n212 B.n149 585
R634 B.n211 B.n210 585
R635 B.n209 B.n150 585
R636 B.n208 B.n207 585
R637 B.n206 B.n151 585
R638 B.n205 B.n204 585
R639 B.n203 B.n152 585
R640 B.n202 B.n201 585
R641 B.n200 B.n153 585
R642 B.n199 B.n198 585
R643 B.n197 B.n154 585
R644 B.n196 B.n195 585
R645 B.n194 B.n155 585
R646 B.n193 B.n192 585
R647 B.n191 B.n156 585
R648 B.n190 B.n189 585
R649 B.n188 B.n157 585
R650 B.n187 B.n186 585
R651 B.n185 B.n158 585
R652 B.n184 B.n183 585
R653 B.n182 B.n159 585
R654 B.n181 B.n180 585
R655 B.n179 B.n160 585
R656 B.n178 B.n177 585
R657 B.n176 B.n161 585
R658 B.n175 B.n174 585
R659 B.n173 B.n162 585
R660 B.n172 B.n171 585
R661 B.n170 B.n163 585
R662 B.n169 B.n168 585
R663 B.n167 B.n164 585
R664 B.n166 B.n165 585
R665 B.n2 B.n0 585
R666 B.n629 B.n1 585
R667 B.n628 B.n627 585
R668 B.n626 B.n3 585
R669 B.n625 B.n624 585
R670 B.n623 B.n4 585
R671 B.n622 B.n621 585
R672 B.n620 B.n5 585
R673 B.n619 B.n618 585
R674 B.n617 B.n6 585
R675 B.n616 B.n615 585
R676 B.n614 B.n7 585
R677 B.n613 B.n612 585
R678 B.n611 B.n8 585
R679 B.n610 B.n609 585
R680 B.n608 B.n9 585
R681 B.n607 B.n606 585
R682 B.n605 B.n10 585
R683 B.n604 B.n603 585
R684 B.n602 B.n11 585
R685 B.n601 B.n600 585
R686 B.n599 B.n12 585
R687 B.n598 B.n597 585
R688 B.n596 B.n13 585
R689 B.n595 B.n594 585
R690 B.n593 B.n14 585
R691 B.n592 B.n591 585
R692 B.n590 B.n15 585
R693 B.n589 B.n588 585
R694 B.n587 B.n16 585
R695 B.n586 B.n585 585
R696 B.n584 B.n17 585
R697 B.n583 B.n582 585
R698 B.n581 B.n18 585
R699 B.n580 B.n579 585
R700 B.n578 B.n19 585
R701 B.n577 B.n576 585
R702 B.n575 B.n20 585
R703 B.n574 B.n573 585
R704 B.n572 B.n21 585
R705 B.n571 B.n570 585
R706 B.n569 B.n22 585
R707 B.n568 B.n567 585
R708 B.n566 B.n23 585
R709 B.n565 B.n564 585
R710 B.n563 B.n24 585
R711 B.n562 B.n561 585
R712 B.n560 B.n25 585
R713 B.n559 B.n558 585
R714 B.n557 B.n26 585
R715 B.n556 B.n555 585
R716 B.n554 B.n27 585
R717 B.n553 B.n552 585
R718 B.n551 B.n28 585
R719 B.n550 B.n549 585
R720 B.n548 B.n29 585
R721 B.n547 B.n546 585
R722 B.n545 B.n30 585
R723 B.n544 B.n543 585
R724 B.n631 B.n630 585
R725 B.n251 B.n250 458.866
R726 B.n544 B.n31 458.866
R727 B.n310 B.n113 458.866
R728 B.n485 B.n484 458.866
R729 B.n120 B.t2 292.13
R730 B.n46 B.t4 292.13
R731 B.n128 B.t11 292.13
R732 B.n38 B.t7 292.13
R733 B.n120 B.t0 229.206
R734 B.n128 B.t9 229.206
R735 B.n38 B.t6 229.206
R736 B.n46 B.t3 229.206
R737 B.n121 B.t1 226.385
R738 B.n47 B.t5 226.385
R739 B.n129 B.t10 226.385
R740 B.n39 B.t8 226.385
R741 B.n250 B.n137 163.367
R742 B.n246 B.n137 163.367
R743 B.n246 B.n245 163.367
R744 B.n245 B.n244 163.367
R745 B.n244 B.n139 163.367
R746 B.n240 B.n139 163.367
R747 B.n240 B.n239 163.367
R748 B.n239 B.n238 163.367
R749 B.n238 B.n141 163.367
R750 B.n234 B.n141 163.367
R751 B.n234 B.n233 163.367
R752 B.n233 B.n232 163.367
R753 B.n232 B.n143 163.367
R754 B.n228 B.n143 163.367
R755 B.n228 B.n227 163.367
R756 B.n227 B.n226 163.367
R757 B.n226 B.n145 163.367
R758 B.n222 B.n145 163.367
R759 B.n222 B.n221 163.367
R760 B.n221 B.n220 163.367
R761 B.n220 B.n147 163.367
R762 B.n216 B.n147 163.367
R763 B.n216 B.n215 163.367
R764 B.n215 B.n214 163.367
R765 B.n214 B.n149 163.367
R766 B.n210 B.n149 163.367
R767 B.n210 B.n209 163.367
R768 B.n209 B.n208 163.367
R769 B.n208 B.n151 163.367
R770 B.n204 B.n151 163.367
R771 B.n204 B.n203 163.367
R772 B.n203 B.n202 163.367
R773 B.n202 B.n153 163.367
R774 B.n198 B.n153 163.367
R775 B.n198 B.n197 163.367
R776 B.n197 B.n196 163.367
R777 B.n196 B.n155 163.367
R778 B.n192 B.n155 163.367
R779 B.n192 B.n191 163.367
R780 B.n191 B.n190 163.367
R781 B.n190 B.n157 163.367
R782 B.n186 B.n157 163.367
R783 B.n186 B.n185 163.367
R784 B.n185 B.n184 163.367
R785 B.n184 B.n159 163.367
R786 B.n180 B.n159 163.367
R787 B.n180 B.n179 163.367
R788 B.n179 B.n178 163.367
R789 B.n178 B.n161 163.367
R790 B.n174 B.n161 163.367
R791 B.n174 B.n173 163.367
R792 B.n173 B.n172 163.367
R793 B.n172 B.n163 163.367
R794 B.n168 B.n163 163.367
R795 B.n168 B.n167 163.367
R796 B.n167 B.n166 163.367
R797 B.n166 B.n2 163.367
R798 B.n630 B.n2 163.367
R799 B.n630 B.n629 163.367
R800 B.n629 B.n628 163.367
R801 B.n628 B.n3 163.367
R802 B.n624 B.n3 163.367
R803 B.n624 B.n623 163.367
R804 B.n623 B.n622 163.367
R805 B.n622 B.n5 163.367
R806 B.n618 B.n5 163.367
R807 B.n618 B.n617 163.367
R808 B.n617 B.n616 163.367
R809 B.n616 B.n7 163.367
R810 B.n612 B.n7 163.367
R811 B.n612 B.n611 163.367
R812 B.n611 B.n610 163.367
R813 B.n610 B.n9 163.367
R814 B.n606 B.n9 163.367
R815 B.n606 B.n605 163.367
R816 B.n605 B.n604 163.367
R817 B.n604 B.n11 163.367
R818 B.n600 B.n11 163.367
R819 B.n600 B.n599 163.367
R820 B.n599 B.n598 163.367
R821 B.n598 B.n13 163.367
R822 B.n594 B.n13 163.367
R823 B.n594 B.n593 163.367
R824 B.n593 B.n592 163.367
R825 B.n592 B.n15 163.367
R826 B.n588 B.n15 163.367
R827 B.n588 B.n587 163.367
R828 B.n587 B.n586 163.367
R829 B.n586 B.n17 163.367
R830 B.n582 B.n17 163.367
R831 B.n582 B.n581 163.367
R832 B.n581 B.n580 163.367
R833 B.n580 B.n19 163.367
R834 B.n576 B.n19 163.367
R835 B.n576 B.n575 163.367
R836 B.n575 B.n574 163.367
R837 B.n574 B.n21 163.367
R838 B.n570 B.n21 163.367
R839 B.n570 B.n569 163.367
R840 B.n569 B.n568 163.367
R841 B.n568 B.n23 163.367
R842 B.n564 B.n23 163.367
R843 B.n564 B.n563 163.367
R844 B.n563 B.n562 163.367
R845 B.n562 B.n25 163.367
R846 B.n558 B.n25 163.367
R847 B.n558 B.n557 163.367
R848 B.n557 B.n556 163.367
R849 B.n556 B.n27 163.367
R850 B.n552 B.n27 163.367
R851 B.n552 B.n551 163.367
R852 B.n551 B.n550 163.367
R853 B.n550 B.n29 163.367
R854 B.n546 B.n29 163.367
R855 B.n546 B.n545 163.367
R856 B.n545 B.n544 163.367
R857 B.n252 B.n251 163.367
R858 B.n252 B.n135 163.367
R859 B.n256 B.n135 163.367
R860 B.n257 B.n256 163.367
R861 B.n258 B.n257 163.367
R862 B.n258 B.n133 163.367
R863 B.n262 B.n133 163.367
R864 B.n263 B.n262 163.367
R865 B.n264 B.n263 163.367
R866 B.n264 B.n131 163.367
R867 B.n268 B.n131 163.367
R868 B.n269 B.n268 163.367
R869 B.n270 B.n269 163.367
R870 B.n270 B.n127 163.367
R871 B.n275 B.n127 163.367
R872 B.n276 B.n275 163.367
R873 B.n277 B.n276 163.367
R874 B.n277 B.n125 163.367
R875 B.n281 B.n125 163.367
R876 B.n282 B.n281 163.367
R877 B.n283 B.n282 163.367
R878 B.n283 B.n123 163.367
R879 B.n287 B.n123 163.367
R880 B.n288 B.n287 163.367
R881 B.n288 B.n119 163.367
R882 B.n292 B.n119 163.367
R883 B.n293 B.n292 163.367
R884 B.n294 B.n293 163.367
R885 B.n294 B.n117 163.367
R886 B.n298 B.n117 163.367
R887 B.n299 B.n298 163.367
R888 B.n300 B.n299 163.367
R889 B.n300 B.n115 163.367
R890 B.n304 B.n115 163.367
R891 B.n305 B.n304 163.367
R892 B.n306 B.n305 163.367
R893 B.n306 B.n113 163.367
R894 B.n311 B.n310 163.367
R895 B.n312 B.n311 163.367
R896 B.n312 B.n111 163.367
R897 B.n316 B.n111 163.367
R898 B.n317 B.n316 163.367
R899 B.n318 B.n317 163.367
R900 B.n318 B.n109 163.367
R901 B.n322 B.n109 163.367
R902 B.n323 B.n322 163.367
R903 B.n324 B.n323 163.367
R904 B.n324 B.n107 163.367
R905 B.n328 B.n107 163.367
R906 B.n329 B.n328 163.367
R907 B.n330 B.n329 163.367
R908 B.n330 B.n105 163.367
R909 B.n334 B.n105 163.367
R910 B.n335 B.n334 163.367
R911 B.n336 B.n335 163.367
R912 B.n336 B.n103 163.367
R913 B.n340 B.n103 163.367
R914 B.n341 B.n340 163.367
R915 B.n342 B.n341 163.367
R916 B.n342 B.n101 163.367
R917 B.n346 B.n101 163.367
R918 B.n347 B.n346 163.367
R919 B.n348 B.n347 163.367
R920 B.n348 B.n99 163.367
R921 B.n352 B.n99 163.367
R922 B.n353 B.n352 163.367
R923 B.n354 B.n353 163.367
R924 B.n354 B.n97 163.367
R925 B.n358 B.n97 163.367
R926 B.n359 B.n358 163.367
R927 B.n360 B.n359 163.367
R928 B.n360 B.n95 163.367
R929 B.n364 B.n95 163.367
R930 B.n365 B.n364 163.367
R931 B.n366 B.n365 163.367
R932 B.n366 B.n93 163.367
R933 B.n370 B.n93 163.367
R934 B.n371 B.n370 163.367
R935 B.n372 B.n371 163.367
R936 B.n372 B.n91 163.367
R937 B.n376 B.n91 163.367
R938 B.n377 B.n376 163.367
R939 B.n378 B.n377 163.367
R940 B.n378 B.n89 163.367
R941 B.n382 B.n89 163.367
R942 B.n383 B.n382 163.367
R943 B.n384 B.n383 163.367
R944 B.n384 B.n87 163.367
R945 B.n388 B.n87 163.367
R946 B.n389 B.n388 163.367
R947 B.n390 B.n389 163.367
R948 B.n390 B.n85 163.367
R949 B.n394 B.n85 163.367
R950 B.n395 B.n394 163.367
R951 B.n396 B.n395 163.367
R952 B.n396 B.n83 163.367
R953 B.n400 B.n83 163.367
R954 B.n401 B.n400 163.367
R955 B.n402 B.n401 163.367
R956 B.n402 B.n81 163.367
R957 B.n406 B.n81 163.367
R958 B.n407 B.n406 163.367
R959 B.n408 B.n407 163.367
R960 B.n408 B.n79 163.367
R961 B.n412 B.n79 163.367
R962 B.n413 B.n412 163.367
R963 B.n414 B.n413 163.367
R964 B.n414 B.n77 163.367
R965 B.n418 B.n77 163.367
R966 B.n419 B.n418 163.367
R967 B.n420 B.n419 163.367
R968 B.n420 B.n75 163.367
R969 B.n424 B.n75 163.367
R970 B.n425 B.n424 163.367
R971 B.n426 B.n425 163.367
R972 B.n426 B.n73 163.367
R973 B.n430 B.n73 163.367
R974 B.n431 B.n430 163.367
R975 B.n432 B.n431 163.367
R976 B.n432 B.n71 163.367
R977 B.n436 B.n71 163.367
R978 B.n437 B.n436 163.367
R979 B.n438 B.n437 163.367
R980 B.n438 B.n69 163.367
R981 B.n442 B.n69 163.367
R982 B.n443 B.n442 163.367
R983 B.n444 B.n443 163.367
R984 B.n444 B.n67 163.367
R985 B.n448 B.n67 163.367
R986 B.n449 B.n448 163.367
R987 B.n450 B.n449 163.367
R988 B.n450 B.n65 163.367
R989 B.n454 B.n65 163.367
R990 B.n455 B.n454 163.367
R991 B.n456 B.n455 163.367
R992 B.n456 B.n63 163.367
R993 B.n460 B.n63 163.367
R994 B.n461 B.n460 163.367
R995 B.n462 B.n461 163.367
R996 B.n462 B.n61 163.367
R997 B.n466 B.n61 163.367
R998 B.n467 B.n466 163.367
R999 B.n468 B.n467 163.367
R1000 B.n468 B.n59 163.367
R1001 B.n472 B.n59 163.367
R1002 B.n473 B.n472 163.367
R1003 B.n474 B.n473 163.367
R1004 B.n474 B.n57 163.367
R1005 B.n478 B.n57 163.367
R1006 B.n479 B.n478 163.367
R1007 B.n480 B.n479 163.367
R1008 B.n480 B.n55 163.367
R1009 B.n484 B.n55 163.367
R1010 B.n540 B.n31 163.367
R1011 B.n540 B.n539 163.367
R1012 B.n539 B.n538 163.367
R1013 B.n538 B.n33 163.367
R1014 B.n534 B.n33 163.367
R1015 B.n534 B.n533 163.367
R1016 B.n533 B.n532 163.367
R1017 B.n532 B.n35 163.367
R1018 B.n528 B.n35 163.367
R1019 B.n528 B.n527 163.367
R1020 B.n527 B.n526 163.367
R1021 B.n526 B.n37 163.367
R1022 B.n522 B.n37 163.367
R1023 B.n522 B.n521 163.367
R1024 B.n521 B.n41 163.367
R1025 B.n517 B.n41 163.367
R1026 B.n517 B.n516 163.367
R1027 B.n516 B.n515 163.367
R1028 B.n515 B.n43 163.367
R1029 B.n511 B.n43 163.367
R1030 B.n511 B.n510 163.367
R1031 B.n510 B.n509 163.367
R1032 B.n509 B.n45 163.367
R1033 B.n504 B.n45 163.367
R1034 B.n504 B.n503 163.367
R1035 B.n503 B.n502 163.367
R1036 B.n502 B.n49 163.367
R1037 B.n498 B.n49 163.367
R1038 B.n498 B.n497 163.367
R1039 B.n497 B.n496 163.367
R1040 B.n496 B.n51 163.367
R1041 B.n492 B.n51 163.367
R1042 B.n492 B.n491 163.367
R1043 B.n491 B.n490 163.367
R1044 B.n490 B.n53 163.367
R1045 B.n486 B.n53 163.367
R1046 B.n486 B.n485 163.367
R1047 B.n121 B.n120 65.746
R1048 B.n129 B.n128 65.746
R1049 B.n39 B.n38 65.746
R1050 B.n47 B.n46 65.746
R1051 B.n122 B.n121 59.5399
R1052 B.n272 B.n129 59.5399
R1053 B.n40 B.n39 59.5399
R1054 B.n506 B.n47 59.5399
R1055 B.n483 B.n54 29.8151
R1056 B.n543 B.n542 29.8151
R1057 B.n309 B.n308 29.8151
R1058 B.n249 B.n136 29.8151
R1059 B B.n631 18.0485
R1060 B.n542 B.n541 10.6151
R1061 B.n541 B.n32 10.6151
R1062 B.n537 B.n32 10.6151
R1063 B.n537 B.n536 10.6151
R1064 B.n536 B.n535 10.6151
R1065 B.n535 B.n34 10.6151
R1066 B.n531 B.n34 10.6151
R1067 B.n531 B.n530 10.6151
R1068 B.n530 B.n529 10.6151
R1069 B.n529 B.n36 10.6151
R1070 B.n525 B.n36 10.6151
R1071 B.n525 B.n524 10.6151
R1072 B.n524 B.n523 10.6151
R1073 B.n520 B.n519 10.6151
R1074 B.n519 B.n518 10.6151
R1075 B.n518 B.n42 10.6151
R1076 B.n514 B.n42 10.6151
R1077 B.n514 B.n513 10.6151
R1078 B.n513 B.n512 10.6151
R1079 B.n512 B.n44 10.6151
R1080 B.n508 B.n44 10.6151
R1081 B.n508 B.n507 10.6151
R1082 B.n505 B.n48 10.6151
R1083 B.n501 B.n48 10.6151
R1084 B.n501 B.n500 10.6151
R1085 B.n500 B.n499 10.6151
R1086 B.n499 B.n50 10.6151
R1087 B.n495 B.n50 10.6151
R1088 B.n495 B.n494 10.6151
R1089 B.n494 B.n493 10.6151
R1090 B.n493 B.n52 10.6151
R1091 B.n489 B.n52 10.6151
R1092 B.n489 B.n488 10.6151
R1093 B.n488 B.n487 10.6151
R1094 B.n487 B.n54 10.6151
R1095 B.n309 B.n112 10.6151
R1096 B.n313 B.n112 10.6151
R1097 B.n314 B.n313 10.6151
R1098 B.n315 B.n314 10.6151
R1099 B.n315 B.n110 10.6151
R1100 B.n319 B.n110 10.6151
R1101 B.n320 B.n319 10.6151
R1102 B.n321 B.n320 10.6151
R1103 B.n321 B.n108 10.6151
R1104 B.n325 B.n108 10.6151
R1105 B.n326 B.n325 10.6151
R1106 B.n327 B.n326 10.6151
R1107 B.n327 B.n106 10.6151
R1108 B.n331 B.n106 10.6151
R1109 B.n332 B.n331 10.6151
R1110 B.n333 B.n332 10.6151
R1111 B.n333 B.n104 10.6151
R1112 B.n337 B.n104 10.6151
R1113 B.n338 B.n337 10.6151
R1114 B.n339 B.n338 10.6151
R1115 B.n339 B.n102 10.6151
R1116 B.n343 B.n102 10.6151
R1117 B.n344 B.n343 10.6151
R1118 B.n345 B.n344 10.6151
R1119 B.n345 B.n100 10.6151
R1120 B.n349 B.n100 10.6151
R1121 B.n350 B.n349 10.6151
R1122 B.n351 B.n350 10.6151
R1123 B.n351 B.n98 10.6151
R1124 B.n355 B.n98 10.6151
R1125 B.n356 B.n355 10.6151
R1126 B.n357 B.n356 10.6151
R1127 B.n357 B.n96 10.6151
R1128 B.n361 B.n96 10.6151
R1129 B.n362 B.n361 10.6151
R1130 B.n363 B.n362 10.6151
R1131 B.n363 B.n94 10.6151
R1132 B.n367 B.n94 10.6151
R1133 B.n368 B.n367 10.6151
R1134 B.n369 B.n368 10.6151
R1135 B.n369 B.n92 10.6151
R1136 B.n373 B.n92 10.6151
R1137 B.n374 B.n373 10.6151
R1138 B.n375 B.n374 10.6151
R1139 B.n375 B.n90 10.6151
R1140 B.n379 B.n90 10.6151
R1141 B.n380 B.n379 10.6151
R1142 B.n381 B.n380 10.6151
R1143 B.n381 B.n88 10.6151
R1144 B.n385 B.n88 10.6151
R1145 B.n386 B.n385 10.6151
R1146 B.n387 B.n386 10.6151
R1147 B.n387 B.n86 10.6151
R1148 B.n391 B.n86 10.6151
R1149 B.n392 B.n391 10.6151
R1150 B.n393 B.n392 10.6151
R1151 B.n393 B.n84 10.6151
R1152 B.n397 B.n84 10.6151
R1153 B.n398 B.n397 10.6151
R1154 B.n399 B.n398 10.6151
R1155 B.n399 B.n82 10.6151
R1156 B.n403 B.n82 10.6151
R1157 B.n404 B.n403 10.6151
R1158 B.n405 B.n404 10.6151
R1159 B.n405 B.n80 10.6151
R1160 B.n409 B.n80 10.6151
R1161 B.n410 B.n409 10.6151
R1162 B.n411 B.n410 10.6151
R1163 B.n411 B.n78 10.6151
R1164 B.n415 B.n78 10.6151
R1165 B.n416 B.n415 10.6151
R1166 B.n417 B.n416 10.6151
R1167 B.n417 B.n76 10.6151
R1168 B.n421 B.n76 10.6151
R1169 B.n422 B.n421 10.6151
R1170 B.n423 B.n422 10.6151
R1171 B.n423 B.n74 10.6151
R1172 B.n427 B.n74 10.6151
R1173 B.n428 B.n427 10.6151
R1174 B.n429 B.n428 10.6151
R1175 B.n429 B.n72 10.6151
R1176 B.n433 B.n72 10.6151
R1177 B.n434 B.n433 10.6151
R1178 B.n435 B.n434 10.6151
R1179 B.n435 B.n70 10.6151
R1180 B.n439 B.n70 10.6151
R1181 B.n440 B.n439 10.6151
R1182 B.n441 B.n440 10.6151
R1183 B.n441 B.n68 10.6151
R1184 B.n445 B.n68 10.6151
R1185 B.n446 B.n445 10.6151
R1186 B.n447 B.n446 10.6151
R1187 B.n447 B.n66 10.6151
R1188 B.n451 B.n66 10.6151
R1189 B.n452 B.n451 10.6151
R1190 B.n453 B.n452 10.6151
R1191 B.n453 B.n64 10.6151
R1192 B.n457 B.n64 10.6151
R1193 B.n458 B.n457 10.6151
R1194 B.n459 B.n458 10.6151
R1195 B.n459 B.n62 10.6151
R1196 B.n463 B.n62 10.6151
R1197 B.n464 B.n463 10.6151
R1198 B.n465 B.n464 10.6151
R1199 B.n465 B.n60 10.6151
R1200 B.n469 B.n60 10.6151
R1201 B.n470 B.n469 10.6151
R1202 B.n471 B.n470 10.6151
R1203 B.n471 B.n58 10.6151
R1204 B.n475 B.n58 10.6151
R1205 B.n476 B.n475 10.6151
R1206 B.n477 B.n476 10.6151
R1207 B.n477 B.n56 10.6151
R1208 B.n481 B.n56 10.6151
R1209 B.n482 B.n481 10.6151
R1210 B.n483 B.n482 10.6151
R1211 B.n253 B.n136 10.6151
R1212 B.n254 B.n253 10.6151
R1213 B.n255 B.n254 10.6151
R1214 B.n255 B.n134 10.6151
R1215 B.n259 B.n134 10.6151
R1216 B.n260 B.n259 10.6151
R1217 B.n261 B.n260 10.6151
R1218 B.n261 B.n132 10.6151
R1219 B.n265 B.n132 10.6151
R1220 B.n266 B.n265 10.6151
R1221 B.n267 B.n266 10.6151
R1222 B.n267 B.n130 10.6151
R1223 B.n271 B.n130 10.6151
R1224 B.n274 B.n273 10.6151
R1225 B.n274 B.n126 10.6151
R1226 B.n278 B.n126 10.6151
R1227 B.n279 B.n278 10.6151
R1228 B.n280 B.n279 10.6151
R1229 B.n280 B.n124 10.6151
R1230 B.n284 B.n124 10.6151
R1231 B.n285 B.n284 10.6151
R1232 B.n286 B.n285 10.6151
R1233 B.n290 B.n289 10.6151
R1234 B.n291 B.n290 10.6151
R1235 B.n291 B.n118 10.6151
R1236 B.n295 B.n118 10.6151
R1237 B.n296 B.n295 10.6151
R1238 B.n297 B.n296 10.6151
R1239 B.n297 B.n116 10.6151
R1240 B.n301 B.n116 10.6151
R1241 B.n302 B.n301 10.6151
R1242 B.n303 B.n302 10.6151
R1243 B.n303 B.n114 10.6151
R1244 B.n307 B.n114 10.6151
R1245 B.n308 B.n307 10.6151
R1246 B.n249 B.n248 10.6151
R1247 B.n248 B.n247 10.6151
R1248 B.n247 B.n138 10.6151
R1249 B.n243 B.n138 10.6151
R1250 B.n243 B.n242 10.6151
R1251 B.n242 B.n241 10.6151
R1252 B.n241 B.n140 10.6151
R1253 B.n237 B.n140 10.6151
R1254 B.n237 B.n236 10.6151
R1255 B.n236 B.n235 10.6151
R1256 B.n235 B.n142 10.6151
R1257 B.n231 B.n142 10.6151
R1258 B.n231 B.n230 10.6151
R1259 B.n230 B.n229 10.6151
R1260 B.n229 B.n144 10.6151
R1261 B.n225 B.n144 10.6151
R1262 B.n225 B.n224 10.6151
R1263 B.n224 B.n223 10.6151
R1264 B.n223 B.n146 10.6151
R1265 B.n219 B.n146 10.6151
R1266 B.n219 B.n218 10.6151
R1267 B.n218 B.n217 10.6151
R1268 B.n217 B.n148 10.6151
R1269 B.n213 B.n148 10.6151
R1270 B.n213 B.n212 10.6151
R1271 B.n212 B.n211 10.6151
R1272 B.n211 B.n150 10.6151
R1273 B.n207 B.n150 10.6151
R1274 B.n207 B.n206 10.6151
R1275 B.n206 B.n205 10.6151
R1276 B.n205 B.n152 10.6151
R1277 B.n201 B.n152 10.6151
R1278 B.n201 B.n200 10.6151
R1279 B.n200 B.n199 10.6151
R1280 B.n199 B.n154 10.6151
R1281 B.n195 B.n154 10.6151
R1282 B.n195 B.n194 10.6151
R1283 B.n194 B.n193 10.6151
R1284 B.n193 B.n156 10.6151
R1285 B.n189 B.n156 10.6151
R1286 B.n189 B.n188 10.6151
R1287 B.n188 B.n187 10.6151
R1288 B.n187 B.n158 10.6151
R1289 B.n183 B.n158 10.6151
R1290 B.n183 B.n182 10.6151
R1291 B.n182 B.n181 10.6151
R1292 B.n181 B.n160 10.6151
R1293 B.n177 B.n160 10.6151
R1294 B.n177 B.n176 10.6151
R1295 B.n176 B.n175 10.6151
R1296 B.n175 B.n162 10.6151
R1297 B.n171 B.n162 10.6151
R1298 B.n171 B.n170 10.6151
R1299 B.n170 B.n169 10.6151
R1300 B.n169 B.n164 10.6151
R1301 B.n165 B.n164 10.6151
R1302 B.n165 B.n0 10.6151
R1303 B.n627 B.n1 10.6151
R1304 B.n627 B.n626 10.6151
R1305 B.n626 B.n625 10.6151
R1306 B.n625 B.n4 10.6151
R1307 B.n621 B.n4 10.6151
R1308 B.n621 B.n620 10.6151
R1309 B.n620 B.n619 10.6151
R1310 B.n619 B.n6 10.6151
R1311 B.n615 B.n6 10.6151
R1312 B.n615 B.n614 10.6151
R1313 B.n614 B.n613 10.6151
R1314 B.n613 B.n8 10.6151
R1315 B.n609 B.n8 10.6151
R1316 B.n609 B.n608 10.6151
R1317 B.n608 B.n607 10.6151
R1318 B.n607 B.n10 10.6151
R1319 B.n603 B.n10 10.6151
R1320 B.n603 B.n602 10.6151
R1321 B.n602 B.n601 10.6151
R1322 B.n601 B.n12 10.6151
R1323 B.n597 B.n12 10.6151
R1324 B.n597 B.n596 10.6151
R1325 B.n596 B.n595 10.6151
R1326 B.n595 B.n14 10.6151
R1327 B.n591 B.n14 10.6151
R1328 B.n591 B.n590 10.6151
R1329 B.n590 B.n589 10.6151
R1330 B.n589 B.n16 10.6151
R1331 B.n585 B.n16 10.6151
R1332 B.n585 B.n584 10.6151
R1333 B.n584 B.n583 10.6151
R1334 B.n583 B.n18 10.6151
R1335 B.n579 B.n18 10.6151
R1336 B.n579 B.n578 10.6151
R1337 B.n578 B.n577 10.6151
R1338 B.n577 B.n20 10.6151
R1339 B.n573 B.n20 10.6151
R1340 B.n573 B.n572 10.6151
R1341 B.n572 B.n571 10.6151
R1342 B.n571 B.n22 10.6151
R1343 B.n567 B.n22 10.6151
R1344 B.n567 B.n566 10.6151
R1345 B.n566 B.n565 10.6151
R1346 B.n565 B.n24 10.6151
R1347 B.n561 B.n24 10.6151
R1348 B.n561 B.n560 10.6151
R1349 B.n560 B.n559 10.6151
R1350 B.n559 B.n26 10.6151
R1351 B.n555 B.n26 10.6151
R1352 B.n555 B.n554 10.6151
R1353 B.n554 B.n553 10.6151
R1354 B.n553 B.n28 10.6151
R1355 B.n549 B.n28 10.6151
R1356 B.n549 B.n548 10.6151
R1357 B.n548 B.n547 10.6151
R1358 B.n547 B.n30 10.6151
R1359 B.n543 B.n30 10.6151
R1360 B.n523 B.n40 9.36635
R1361 B.n506 B.n505 9.36635
R1362 B.n272 B.n271 9.36635
R1363 B.n289 B.n122 9.36635
R1364 B.n631 B.n0 2.81026
R1365 B.n631 B.n1 2.81026
R1366 B.n520 B.n40 1.24928
R1367 B.n507 B.n506 1.24928
R1368 B.n273 B.n272 1.24928
R1369 B.n286 B.n122 1.24928
C0 w_n4360_n1490# VTAIL 2.13672f
C1 VN B 1.23587f
C2 w_n4360_n1490# B 8.234019f
C3 VDD1 VN 0.157831f
C4 VP VTAIL 3.59208f
C5 VDD1 w_n4360_n1490# 1.84857f
C6 VDD2 VTAIL 5.37627f
C7 VP B 2.1889f
C8 B VDD2 1.64639f
C9 VP VDD1 2.72565f
C10 VDD1 VDD2 2.01713f
C11 w_n4360_n1490# VN 8.85045f
C12 B VTAIL 1.94215f
C13 VP VN 6.49688f
C14 VN VDD2 2.31149f
C15 VDD1 VTAIL 5.31877f
C16 VP w_n4360_n1490# 9.414809f
C17 w_n4360_n1490# VDD2 1.98197f
C18 VDD1 B 1.5356f
C19 VP VDD2 0.574922f
C20 VN VTAIL 3.57798f
C21 VDD2 VSUBS 1.736618f
C22 VDD1 VSUBS 2.4802f
C23 VTAIL VSUBS 0.630063f
C24 VN VSUBS 7.39285f
C25 VP VSUBS 3.452136f
C26 B VSUBS 4.432795f
C27 w_n4360_n1490# VSUBS 82.5086f
C28 B.n0 VSUBS 0.006359f
C29 B.n1 VSUBS 0.006359f
C30 B.n2 VSUBS 0.010057f
C31 B.n3 VSUBS 0.010057f
C32 B.n4 VSUBS 0.010057f
C33 B.n5 VSUBS 0.010057f
C34 B.n6 VSUBS 0.010057f
C35 B.n7 VSUBS 0.010057f
C36 B.n8 VSUBS 0.010057f
C37 B.n9 VSUBS 0.010057f
C38 B.n10 VSUBS 0.010057f
C39 B.n11 VSUBS 0.010057f
C40 B.n12 VSUBS 0.010057f
C41 B.n13 VSUBS 0.010057f
C42 B.n14 VSUBS 0.010057f
C43 B.n15 VSUBS 0.010057f
C44 B.n16 VSUBS 0.010057f
C45 B.n17 VSUBS 0.010057f
C46 B.n18 VSUBS 0.010057f
C47 B.n19 VSUBS 0.010057f
C48 B.n20 VSUBS 0.010057f
C49 B.n21 VSUBS 0.010057f
C50 B.n22 VSUBS 0.010057f
C51 B.n23 VSUBS 0.010057f
C52 B.n24 VSUBS 0.010057f
C53 B.n25 VSUBS 0.010057f
C54 B.n26 VSUBS 0.010057f
C55 B.n27 VSUBS 0.010057f
C56 B.n28 VSUBS 0.010057f
C57 B.n29 VSUBS 0.010057f
C58 B.n30 VSUBS 0.010057f
C59 B.n31 VSUBS 0.022993f
C60 B.n32 VSUBS 0.010057f
C61 B.n33 VSUBS 0.010057f
C62 B.n34 VSUBS 0.010057f
C63 B.n35 VSUBS 0.010057f
C64 B.n36 VSUBS 0.010057f
C65 B.n37 VSUBS 0.010057f
C66 B.t8 VSUBS 0.058338f
C67 B.t7 VSUBS 0.082483f
C68 B.t6 VSUBS 0.562546f
C69 B.n38 VSUBS 0.144964f
C70 B.n39 VSUBS 0.121629f
C71 B.n40 VSUBS 0.0233f
C72 B.n41 VSUBS 0.010057f
C73 B.n42 VSUBS 0.010057f
C74 B.n43 VSUBS 0.010057f
C75 B.n44 VSUBS 0.010057f
C76 B.n45 VSUBS 0.010057f
C77 B.t5 VSUBS 0.058338f
C78 B.t4 VSUBS 0.082483f
C79 B.t3 VSUBS 0.562546f
C80 B.n46 VSUBS 0.144964f
C81 B.n47 VSUBS 0.121629f
C82 B.n48 VSUBS 0.010057f
C83 B.n49 VSUBS 0.010057f
C84 B.n50 VSUBS 0.010057f
C85 B.n51 VSUBS 0.010057f
C86 B.n52 VSUBS 0.010057f
C87 B.n53 VSUBS 0.010057f
C88 B.n54 VSUBS 0.021691f
C89 B.n55 VSUBS 0.010057f
C90 B.n56 VSUBS 0.010057f
C91 B.n57 VSUBS 0.010057f
C92 B.n58 VSUBS 0.010057f
C93 B.n59 VSUBS 0.010057f
C94 B.n60 VSUBS 0.010057f
C95 B.n61 VSUBS 0.010057f
C96 B.n62 VSUBS 0.010057f
C97 B.n63 VSUBS 0.010057f
C98 B.n64 VSUBS 0.010057f
C99 B.n65 VSUBS 0.010057f
C100 B.n66 VSUBS 0.010057f
C101 B.n67 VSUBS 0.010057f
C102 B.n68 VSUBS 0.010057f
C103 B.n69 VSUBS 0.010057f
C104 B.n70 VSUBS 0.010057f
C105 B.n71 VSUBS 0.010057f
C106 B.n72 VSUBS 0.010057f
C107 B.n73 VSUBS 0.010057f
C108 B.n74 VSUBS 0.010057f
C109 B.n75 VSUBS 0.010057f
C110 B.n76 VSUBS 0.010057f
C111 B.n77 VSUBS 0.010057f
C112 B.n78 VSUBS 0.010057f
C113 B.n79 VSUBS 0.010057f
C114 B.n80 VSUBS 0.010057f
C115 B.n81 VSUBS 0.010057f
C116 B.n82 VSUBS 0.010057f
C117 B.n83 VSUBS 0.010057f
C118 B.n84 VSUBS 0.010057f
C119 B.n85 VSUBS 0.010057f
C120 B.n86 VSUBS 0.010057f
C121 B.n87 VSUBS 0.010057f
C122 B.n88 VSUBS 0.010057f
C123 B.n89 VSUBS 0.010057f
C124 B.n90 VSUBS 0.010057f
C125 B.n91 VSUBS 0.010057f
C126 B.n92 VSUBS 0.010057f
C127 B.n93 VSUBS 0.010057f
C128 B.n94 VSUBS 0.010057f
C129 B.n95 VSUBS 0.010057f
C130 B.n96 VSUBS 0.010057f
C131 B.n97 VSUBS 0.010057f
C132 B.n98 VSUBS 0.010057f
C133 B.n99 VSUBS 0.010057f
C134 B.n100 VSUBS 0.010057f
C135 B.n101 VSUBS 0.010057f
C136 B.n102 VSUBS 0.010057f
C137 B.n103 VSUBS 0.010057f
C138 B.n104 VSUBS 0.010057f
C139 B.n105 VSUBS 0.010057f
C140 B.n106 VSUBS 0.010057f
C141 B.n107 VSUBS 0.010057f
C142 B.n108 VSUBS 0.010057f
C143 B.n109 VSUBS 0.010057f
C144 B.n110 VSUBS 0.010057f
C145 B.n111 VSUBS 0.010057f
C146 B.n112 VSUBS 0.010057f
C147 B.n113 VSUBS 0.022993f
C148 B.n114 VSUBS 0.010057f
C149 B.n115 VSUBS 0.010057f
C150 B.n116 VSUBS 0.010057f
C151 B.n117 VSUBS 0.010057f
C152 B.n118 VSUBS 0.010057f
C153 B.n119 VSUBS 0.010057f
C154 B.t1 VSUBS 0.058338f
C155 B.t2 VSUBS 0.082483f
C156 B.t0 VSUBS 0.562546f
C157 B.n120 VSUBS 0.144964f
C158 B.n121 VSUBS 0.121629f
C159 B.n122 VSUBS 0.0233f
C160 B.n123 VSUBS 0.010057f
C161 B.n124 VSUBS 0.010057f
C162 B.n125 VSUBS 0.010057f
C163 B.n126 VSUBS 0.010057f
C164 B.n127 VSUBS 0.010057f
C165 B.t10 VSUBS 0.058338f
C166 B.t11 VSUBS 0.082483f
C167 B.t9 VSUBS 0.562546f
C168 B.n128 VSUBS 0.144964f
C169 B.n129 VSUBS 0.121629f
C170 B.n130 VSUBS 0.010057f
C171 B.n131 VSUBS 0.010057f
C172 B.n132 VSUBS 0.010057f
C173 B.n133 VSUBS 0.010057f
C174 B.n134 VSUBS 0.010057f
C175 B.n135 VSUBS 0.010057f
C176 B.n136 VSUBS 0.022993f
C177 B.n137 VSUBS 0.010057f
C178 B.n138 VSUBS 0.010057f
C179 B.n139 VSUBS 0.010057f
C180 B.n140 VSUBS 0.010057f
C181 B.n141 VSUBS 0.010057f
C182 B.n142 VSUBS 0.010057f
C183 B.n143 VSUBS 0.010057f
C184 B.n144 VSUBS 0.010057f
C185 B.n145 VSUBS 0.010057f
C186 B.n146 VSUBS 0.010057f
C187 B.n147 VSUBS 0.010057f
C188 B.n148 VSUBS 0.010057f
C189 B.n149 VSUBS 0.010057f
C190 B.n150 VSUBS 0.010057f
C191 B.n151 VSUBS 0.010057f
C192 B.n152 VSUBS 0.010057f
C193 B.n153 VSUBS 0.010057f
C194 B.n154 VSUBS 0.010057f
C195 B.n155 VSUBS 0.010057f
C196 B.n156 VSUBS 0.010057f
C197 B.n157 VSUBS 0.010057f
C198 B.n158 VSUBS 0.010057f
C199 B.n159 VSUBS 0.010057f
C200 B.n160 VSUBS 0.010057f
C201 B.n161 VSUBS 0.010057f
C202 B.n162 VSUBS 0.010057f
C203 B.n163 VSUBS 0.010057f
C204 B.n164 VSUBS 0.010057f
C205 B.n165 VSUBS 0.010057f
C206 B.n166 VSUBS 0.010057f
C207 B.n167 VSUBS 0.010057f
C208 B.n168 VSUBS 0.010057f
C209 B.n169 VSUBS 0.010057f
C210 B.n170 VSUBS 0.010057f
C211 B.n171 VSUBS 0.010057f
C212 B.n172 VSUBS 0.010057f
C213 B.n173 VSUBS 0.010057f
C214 B.n174 VSUBS 0.010057f
C215 B.n175 VSUBS 0.010057f
C216 B.n176 VSUBS 0.010057f
C217 B.n177 VSUBS 0.010057f
C218 B.n178 VSUBS 0.010057f
C219 B.n179 VSUBS 0.010057f
C220 B.n180 VSUBS 0.010057f
C221 B.n181 VSUBS 0.010057f
C222 B.n182 VSUBS 0.010057f
C223 B.n183 VSUBS 0.010057f
C224 B.n184 VSUBS 0.010057f
C225 B.n185 VSUBS 0.010057f
C226 B.n186 VSUBS 0.010057f
C227 B.n187 VSUBS 0.010057f
C228 B.n188 VSUBS 0.010057f
C229 B.n189 VSUBS 0.010057f
C230 B.n190 VSUBS 0.010057f
C231 B.n191 VSUBS 0.010057f
C232 B.n192 VSUBS 0.010057f
C233 B.n193 VSUBS 0.010057f
C234 B.n194 VSUBS 0.010057f
C235 B.n195 VSUBS 0.010057f
C236 B.n196 VSUBS 0.010057f
C237 B.n197 VSUBS 0.010057f
C238 B.n198 VSUBS 0.010057f
C239 B.n199 VSUBS 0.010057f
C240 B.n200 VSUBS 0.010057f
C241 B.n201 VSUBS 0.010057f
C242 B.n202 VSUBS 0.010057f
C243 B.n203 VSUBS 0.010057f
C244 B.n204 VSUBS 0.010057f
C245 B.n205 VSUBS 0.010057f
C246 B.n206 VSUBS 0.010057f
C247 B.n207 VSUBS 0.010057f
C248 B.n208 VSUBS 0.010057f
C249 B.n209 VSUBS 0.010057f
C250 B.n210 VSUBS 0.010057f
C251 B.n211 VSUBS 0.010057f
C252 B.n212 VSUBS 0.010057f
C253 B.n213 VSUBS 0.010057f
C254 B.n214 VSUBS 0.010057f
C255 B.n215 VSUBS 0.010057f
C256 B.n216 VSUBS 0.010057f
C257 B.n217 VSUBS 0.010057f
C258 B.n218 VSUBS 0.010057f
C259 B.n219 VSUBS 0.010057f
C260 B.n220 VSUBS 0.010057f
C261 B.n221 VSUBS 0.010057f
C262 B.n222 VSUBS 0.010057f
C263 B.n223 VSUBS 0.010057f
C264 B.n224 VSUBS 0.010057f
C265 B.n225 VSUBS 0.010057f
C266 B.n226 VSUBS 0.010057f
C267 B.n227 VSUBS 0.010057f
C268 B.n228 VSUBS 0.010057f
C269 B.n229 VSUBS 0.010057f
C270 B.n230 VSUBS 0.010057f
C271 B.n231 VSUBS 0.010057f
C272 B.n232 VSUBS 0.010057f
C273 B.n233 VSUBS 0.010057f
C274 B.n234 VSUBS 0.010057f
C275 B.n235 VSUBS 0.010057f
C276 B.n236 VSUBS 0.010057f
C277 B.n237 VSUBS 0.010057f
C278 B.n238 VSUBS 0.010057f
C279 B.n239 VSUBS 0.010057f
C280 B.n240 VSUBS 0.010057f
C281 B.n241 VSUBS 0.010057f
C282 B.n242 VSUBS 0.010057f
C283 B.n243 VSUBS 0.010057f
C284 B.n244 VSUBS 0.010057f
C285 B.n245 VSUBS 0.010057f
C286 B.n246 VSUBS 0.010057f
C287 B.n247 VSUBS 0.010057f
C288 B.n248 VSUBS 0.010057f
C289 B.n249 VSUBS 0.021374f
C290 B.n250 VSUBS 0.021374f
C291 B.n251 VSUBS 0.022993f
C292 B.n252 VSUBS 0.010057f
C293 B.n253 VSUBS 0.010057f
C294 B.n254 VSUBS 0.010057f
C295 B.n255 VSUBS 0.010057f
C296 B.n256 VSUBS 0.010057f
C297 B.n257 VSUBS 0.010057f
C298 B.n258 VSUBS 0.010057f
C299 B.n259 VSUBS 0.010057f
C300 B.n260 VSUBS 0.010057f
C301 B.n261 VSUBS 0.010057f
C302 B.n262 VSUBS 0.010057f
C303 B.n263 VSUBS 0.010057f
C304 B.n264 VSUBS 0.010057f
C305 B.n265 VSUBS 0.010057f
C306 B.n266 VSUBS 0.010057f
C307 B.n267 VSUBS 0.010057f
C308 B.n268 VSUBS 0.010057f
C309 B.n269 VSUBS 0.010057f
C310 B.n270 VSUBS 0.010057f
C311 B.n271 VSUBS 0.009465f
C312 B.n272 VSUBS 0.0233f
C313 B.n273 VSUBS 0.00562f
C314 B.n274 VSUBS 0.010057f
C315 B.n275 VSUBS 0.010057f
C316 B.n276 VSUBS 0.010057f
C317 B.n277 VSUBS 0.010057f
C318 B.n278 VSUBS 0.010057f
C319 B.n279 VSUBS 0.010057f
C320 B.n280 VSUBS 0.010057f
C321 B.n281 VSUBS 0.010057f
C322 B.n282 VSUBS 0.010057f
C323 B.n283 VSUBS 0.010057f
C324 B.n284 VSUBS 0.010057f
C325 B.n285 VSUBS 0.010057f
C326 B.n286 VSUBS 0.00562f
C327 B.n287 VSUBS 0.010057f
C328 B.n288 VSUBS 0.010057f
C329 B.n289 VSUBS 0.009465f
C330 B.n290 VSUBS 0.010057f
C331 B.n291 VSUBS 0.010057f
C332 B.n292 VSUBS 0.010057f
C333 B.n293 VSUBS 0.010057f
C334 B.n294 VSUBS 0.010057f
C335 B.n295 VSUBS 0.010057f
C336 B.n296 VSUBS 0.010057f
C337 B.n297 VSUBS 0.010057f
C338 B.n298 VSUBS 0.010057f
C339 B.n299 VSUBS 0.010057f
C340 B.n300 VSUBS 0.010057f
C341 B.n301 VSUBS 0.010057f
C342 B.n302 VSUBS 0.010057f
C343 B.n303 VSUBS 0.010057f
C344 B.n304 VSUBS 0.010057f
C345 B.n305 VSUBS 0.010057f
C346 B.n306 VSUBS 0.010057f
C347 B.n307 VSUBS 0.010057f
C348 B.n308 VSUBS 0.022993f
C349 B.n309 VSUBS 0.021374f
C350 B.n310 VSUBS 0.021374f
C351 B.n311 VSUBS 0.010057f
C352 B.n312 VSUBS 0.010057f
C353 B.n313 VSUBS 0.010057f
C354 B.n314 VSUBS 0.010057f
C355 B.n315 VSUBS 0.010057f
C356 B.n316 VSUBS 0.010057f
C357 B.n317 VSUBS 0.010057f
C358 B.n318 VSUBS 0.010057f
C359 B.n319 VSUBS 0.010057f
C360 B.n320 VSUBS 0.010057f
C361 B.n321 VSUBS 0.010057f
C362 B.n322 VSUBS 0.010057f
C363 B.n323 VSUBS 0.010057f
C364 B.n324 VSUBS 0.010057f
C365 B.n325 VSUBS 0.010057f
C366 B.n326 VSUBS 0.010057f
C367 B.n327 VSUBS 0.010057f
C368 B.n328 VSUBS 0.010057f
C369 B.n329 VSUBS 0.010057f
C370 B.n330 VSUBS 0.010057f
C371 B.n331 VSUBS 0.010057f
C372 B.n332 VSUBS 0.010057f
C373 B.n333 VSUBS 0.010057f
C374 B.n334 VSUBS 0.010057f
C375 B.n335 VSUBS 0.010057f
C376 B.n336 VSUBS 0.010057f
C377 B.n337 VSUBS 0.010057f
C378 B.n338 VSUBS 0.010057f
C379 B.n339 VSUBS 0.010057f
C380 B.n340 VSUBS 0.010057f
C381 B.n341 VSUBS 0.010057f
C382 B.n342 VSUBS 0.010057f
C383 B.n343 VSUBS 0.010057f
C384 B.n344 VSUBS 0.010057f
C385 B.n345 VSUBS 0.010057f
C386 B.n346 VSUBS 0.010057f
C387 B.n347 VSUBS 0.010057f
C388 B.n348 VSUBS 0.010057f
C389 B.n349 VSUBS 0.010057f
C390 B.n350 VSUBS 0.010057f
C391 B.n351 VSUBS 0.010057f
C392 B.n352 VSUBS 0.010057f
C393 B.n353 VSUBS 0.010057f
C394 B.n354 VSUBS 0.010057f
C395 B.n355 VSUBS 0.010057f
C396 B.n356 VSUBS 0.010057f
C397 B.n357 VSUBS 0.010057f
C398 B.n358 VSUBS 0.010057f
C399 B.n359 VSUBS 0.010057f
C400 B.n360 VSUBS 0.010057f
C401 B.n361 VSUBS 0.010057f
C402 B.n362 VSUBS 0.010057f
C403 B.n363 VSUBS 0.010057f
C404 B.n364 VSUBS 0.010057f
C405 B.n365 VSUBS 0.010057f
C406 B.n366 VSUBS 0.010057f
C407 B.n367 VSUBS 0.010057f
C408 B.n368 VSUBS 0.010057f
C409 B.n369 VSUBS 0.010057f
C410 B.n370 VSUBS 0.010057f
C411 B.n371 VSUBS 0.010057f
C412 B.n372 VSUBS 0.010057f
C413 B.n373 VSUBS 0.010057f
C414 B.n374 VSUBS 0.010057f
C415 B.n375 VSUBS 0.010057f
C416 B.n376 VSUBS 0.010057f
C417 B.n377 VSUBS 0.010057f
C418 B.n378 VSUBS 0.010057f
C419 B.n379 VSUBS 0.010057f
C420 B.n380 VSUBS 0.010057f
C421 B.n381 VSUBS 0.010057f
C422 B.n382 VSUBS 0.010057f
C423 B.n383 VSUBS 0.010057f
C424 B.n384 VSUBS 0.010057f
C425 B.n385 VSUBS 0.010057f
C426 B.n386 VSUBS 0.010057f
C427 B.n387 VSUBS 0.010057f
C428 B.n388 VSUBS 0.010057f
C429 B.n389 VSUBS 0.010057f
C430 B.n390 VSUBS 0.010057f
C431 B.n391 VSUBS 0.010057f
C432 B.n392 VSUBS 0.010057f
C433 B.n393 VSUBS 0.010057f
C434 B.n394 VSUBS 0.010057f
C435 B.n395 VSUBS 0.010057f
C436 B.n396 VSUBS 0.010057f
C437 B.n397 VSUBS 0.010057f
C438 B.n398 VSUBS 0.010057f
C439 B.n399 VSUBS 0.010057f
C440 B.n400 VSUBS 0.010057f
C441 B.n401 VSUBS 0.010057f
C442 B.n402 VSUBS 0.010057f
C443 B.n403 VSUBS 0.010057f
C444 B.n404 VSUBS 0.010057f
C445 B.n405 VSUBS 0.010057f
C446 B.n406 VSUBS 0.010057f
C447 B.n407 VSUBS 0.010057f
C448 B.n408 VSUBS 0.010057f
C449 B.n409 VSUBS 0.010057f
C450 B.n410 VSUBS 0.010057f
C451 B.n411 VSUBS 0.010057f
C452 B.n412 VSUBS 0.010057f
C453 B.n413 VSUBS 0.010057f
C454 B.n414 VSUBS 0.010057f
C455 B.n415 VSUBS 0.010057f
C456 B.n416 VSUBS 0.010057f
C457 B.n417 VSUBS 0.010057f
C458 B.n418 VSUBS 0.010057f
C459 B.n419 VSUBS 0.010057f
C460 B.n420 VSUBS 0.010057f
C461 B.n421 VSUBS 0.010057f
C462 B.n422 VSUBS 0.010057f
C463 B.n423 VSUBS 0.010057f
C464 B.n424 VSUBS 0.010057f
C465 B.n425 VSUBS 0.010057f
C466 B.n426 VSUBS 0.010057f
C467 B.n427 VSUBS 0.010057f
C468 B.n428 VSUBS 0.010057f
C469 B.n429 VSUBS 0.010057f
C470 B.n430 VSUBS 0.010057f
C471 B.n431 VSUBS 0.010057f
C472 B.n432 VSUBS 0.010057f
C473 B.n433 VSUBS 0.010057f
C474 B.n434 VSUBS 0.010057f
C475 B.n435 VSUBS 0.010057f
C476 B.n436 VSUBS 0.010057f
C477 B.n437 VSUBS 0.010057f
C478 B.n438 VSUBS 0.010057f
C479 B.n439 VSUBS 0.010057f
C480 B.n440 VSUBS 0.010057f
C481 B.n441 VSUBS 0.010057f
C482 B.n442 VSUBS 0.010057f
C483 B.n443 VSUBS 0.010057f
C484 B.n444 VSUBS 0.010057f
C485 B.n445 VSUBS 0.010057f
C486 B.n446 VSUBS 0.010057f
C487 B.n447 VSUBS 0.010057f
C488 B.n448 VSUBS 0.010057f
C489 B.n449 VSUBS 0.010057f
C490 B.n450 VSUBS 0.010057f
C491 B.n451 VSUBS 0.010057f
C492 B.n452 VSUBS 0.010057f
C493 B.n453 VSUBS 0.010057f
C494 B.n454 VSUBS 0.010057f
C495 B.n455 VSUBS 0.010057f
C496 B.n456 VSUBS 0.010057f
C497 B.n457 VSUBS 0.010057f
C498 B.n458 VSUBS 0.010057f
C499 B.n459 VSUBS 0.010057f
C500 B.n460 VSUBS 0.010057f
C501 B.n461 VSUBS 0.010057f
C502 B.n462 VSUBS 0.010057f
C503 B.n463 VSUBS 0.010057f
C504 B.n464 VSUBS 0.010057f
C505 B.n465 VSUBS 0.010057f
C506 B.n466 VSUBS 0.010057f
C507 B.n467 VSUBS 0.010057f
C508 B.n468 VSUBS 0.010057f
C509 B.n469 VSUBS 0.010057f
C510 B.n470 VSUBS 0.010057f
C511 B.n471 VSUBS 0.010057f
C512 B.n472 VSUBS 0.010057f
C513 B.n473 VSUBS 0.010057f
C514 B.n474 VSUBS 0.010057f
C515 B.n475 VSUBS 0.010057f
C516 B.n476 VSUBS 0.010057f
C517 B.n477 VSUBS 0.010057f
C518 B.n478 VSUBS 0.010057f
C519 B.n479 VSUBS 0.010057f
C520 B.n480 VSUBS 0.010057f
C521 B.n481 VSUBS 0.010057f
C522 B.n482 VSUBS 0.010057f
C523 B.n483 VSUBS 0.022675f
C524 B.n484 VSUBS 0.021374f
C525 B.n485 VSUBS 0.022993f
C526 B.n486 VSUBS 0.010057f
C527 B.n487 VSUBS 0.010057f
C528 B.n488 VSUBS 0.010057f
C529 B.n489 VSUBS 0.010057f
C530 B.n490 VSUBS 0.010057f
C531 B.n491 VSUBS 0.010057f
C532 B.n492 VSUBS 0.010057f
C533 B.n493 VSUBS 0.010057f
C534 B.n494 VSUBS 0.010057f
C535 B.n495 VSUBS 0.010057f
C536 B.n496 VSUBS 0.010057f
C537 B.n497 VSUBS 0.010057f
C538 B.n498 VSUBS 0.010057f
C539 B.n499 VSUBS 0.010057f
C540 B.n500 VSUBS 0.010057f
C541 B.n501 VSUBS 0.010057f
C542 B.n502 VSUBS 0.010057f
C543 B.n503 VSUBS 0.010057f
C544 B.n504 VSUBS 0.010057f
C545 B.n505 VSUBS 0.009465f
C546 B.n506 VSUBS 0.0233f
C547 B.n507 VSUBS 0.00562f
C548 B.n508 VSUBS 0.010057f
C549 B.n509 VSUBS 0.010057f
C550 B.n510 VSUBS 0.010057f
C551 B.n511 VSUBS 0.010057f
C552 B.n512 VSUBS 0.010057f
C553 B.n513 VSUBS 0.010057f
C554 B.n514 VSUBS 0.010057f
C555 B.n515 VSUBS 0.010057f
C556 B.n516 VSUBS 0.010057f
C557 B.n517 VSUBS 0.010057f
C558 B.n518 VSUBS 0.010057f
C559 B.n519 VSUBS 0.010057f
C560 B.n520 VSUBS 0.00562f
C561 B.n521 VSUBS 0.010057f
C562 B.n522 VSUBS 0.010057f
C563 B.n523 VSUBS 0.009465f
C564 B.n524 VSUBS 0.010057f
C565 B.n525 VSUBS 0.010057f
C566 B.n526 VSUBS 0.010057f
C567 B.n527 VSUBS 0.010057f
C568 B.n528 VSUBS 0.010057f
C569 B.n529 VSUBS 0.010057f
C570 B.n530 VSUBS 0.010057f
C571 B.n531 VSUBS 0.010057f
C572 B.n532 VSUBS 0.010057f
C573 B.n533 VSUBS 0.010057f
C574 B.n534 VSUBS 0.010057f
C575 B.n535 VSUBS 0.010057f
C576 B.n536 VSUBS 0.010057f
C577 B.n537 VSUBS 0.010057f
C578 B.n538 VSUBS 0.010057f
C579 B.n539 VSUBS 0.010057f
C580 B.n540 VSUBS 0.010057f
C581 B.n541 VSUBS 0.010057f
C582 B.n542 VSUBS 0.022993f
C583 B.n543 VSUBS 0.021374f
C584 B.n544 VSUBS 0.021374f
C585 B.n545 VSUBS 0.010057f
C586 B.n546 VSUBS 0.010057f
C587 B.n547 VSUBS 0.010057f
C588 B.n548 VSUBS 0.010057f
C589 B.n549 VSUBS 0.010057f
C590 B.n550 VSUBS 0.010057f
C591 B.n551 VSUBS 0.010057f
C592 B.n552 VSUBS 0.010057f
C593 B.n553 VSUBS 0.010057f
C594 B.n554 VSUBS 0.010057f
C595 B.n555 VSUBS 0.010057f
C596 B.n556 VSUBS 0.010057f
C597 B.n557 VSUBS 0.010057f
C598 B.n558 VSUBS 0.010057f
C599 B.n559 VSUBS 0.010057f
C600 B.n560 VSUBS 0.010057f
C601 B.n561 VSUBS 0.010057f
C602 B.n562 VSUBS 0.010057f
C603 B.n563 VSUBS 0.010057f
C604 B.n564 VSUBS 0.010057f
C605 B.n565 VSUBS 0.010057f
C606 B.n566 VSUBS 0.010057f
C607 B.n567 VSUBS 0.010057f
C608 B.n568 VSUBS 0.010057f
C609 B.n569 VSUBS 0.010057f
C610 B.n570 VSUBS 0.010057f
C611 B.n571 VSUBS 0.010057f
C612 B.n572 VSUBS 0.010057f
C613 B.n573 VSUBS 0.010057f
C614 B.n574 VSUBS 0.010057f
C615 B.n575 VSUBS 0.010057f
C616 B.n576 VSUBS 0.010057f
C617 B.n577 VSUBS 0.010057f
C618 B.n578 VSUBS 0.010057f
C619 B.n579 VSUBS 0.010057f
C620 B.n580 VSUBS 0.010057f
C621 B.n581 VSUBS 0.010057f
C622 B.n582 VSUBS 0.010057f
C623 B.n583 VSUBS 0.010057f
C624 B.n584 VSUBS 0.010057f
C625 B.n585 VSUBS 0.010057f
C626 B.n586 VSUBS 0.010057f
C627 B.n587 VSUBS 0.010057f
C628 B.n588 VSUBS 0.010057f
C629 B.n589 VSUBS 0.010057f
C630 B.n590 VSUBS 0.010057f
C631 B.n591 VSUBS 0.010057f
C632 B.n592 VSUBS 0.010057f
C633 B.n593 VSUBS 0.010057f
C634 B.n594 VSUBS 0.010057f
C635 B.n595 VSUBS 0.010057f
C636 B.n596 VSUBS 0.010057f
C637 B.n597 VSUBS 0.010057f
C638 B.n598 VSUBS 0.010057f
C639 B.n599 VSUBS 0.010057f
C640 B.n600 VSUBS 0.010057f
C641 B.n601 VSUBS 0.010057f
C642 B.n602 VSUBS 0.010057f
C643 B.n603 VSUBS 0.010057f
C644 B.n604 VSUBS 0.010057f
C645 B.n605 VSUBS 0.010057f
C646 B.n606 VSUBS 0.010057f
C647 B.n607 VSUBS 0.010057f
C648 B.n608 VSUBS 0.010057f
C649 B.n609 VSUBS 0.010057f
C650 B.n610 VSUBS 0.010057f
C651 B.n611 VSUBS 0.010057f
C652 B.n612 VSUBS 0.010057f
C653 B.n613 VSUBS 0.010057f
C654 B.n614 VSUBS 0.010057f
C655 B.n615 VSUBS 0.010057f
C656 B.n616 VSUBS 0.010057f
C657 B.n617 VSUBS 0.010057f
C658 B.n618 VSUBS 0.010057f
C659 B.n619 VSUBS 0.010057f
C660 B.n620 VSUBS 0.010057f
C661 B.n621 VSUBS 0.010057f
C662 B.n622 VSUBS 0.010057f
C663 B.n623 VSUBS 0.010057f
C664 B.n624 VSUBS 0.010057f
C665 B.n625 VSUBS 0.010057f
C666 B.n626 VSUBS 0.010057f
C667 B.n627 VSUBS 0.010057f
C668 B.n628 VSUBS 0.010057f
C669 B.n629 VSUBS 0.010057f
C670 B.n630 VSUBS 0.010057f
C671 B.n631 VSUBS 0.022771f
C672 VDD2.t6 VSUBS 0.062671f
C673 VDD2.t1 VSUBS 0.062671f
C674 VDD2.n0 VSUBS 0.316285f
C675 VDD2.t7 VSUBS 0.062671f
C676 VDD2.t0 VSUBS 0.062671f
C677 VDD2.n1 VSUBS 0.316285f
C678 VDD2.n2 VSUBS 3.85161f
C679 VDD2.t5 VSUBS 0.062671f
C680 VDD2.t3 VSUBS 0.062671f
C681 VDD2.n3 VSUBS 0.309122f
C682 VDD2.n4 VSUBS 3.00979f
C683 VDD2.t2 VSUBS 0.062671f
C684 VDD2.t4 VSUBS 0.062671f
C685 VDD2.n5 VSUBS 0.316263f
C686 VN.t7 VSUBS 0.911161f
C687 VN.n0 VSUBS 0.567584f
C688 VN.n1 VSUBS 0.04667f
C689 VN.n2 VSUBS 0.050969f
C690 VN.n3 VSUBS 0.04667f
C691 VN.t0 VSUBS 0.911161f
C692 VN.n4 VSUBS 0.391127f
C693 VN.n5 VSUBS 0.04667f
C694 VN.n6 VSUBS 0.068129f
C695 VN.n7 VSUBS 0.53345f
C696 VN.t6 VSUBS 0.911161f
C697 VN.t1 VSUBS 1.35193f
C698 VN.n8 VSUBS 0.539516f
C699 VN.n9 VSUBS 0.559191f
C700 VN.n10 VSUBS 0.082254f
C701 VN.n11 VSUBS 0.08698f
C702 VN.n12 VSUBS 0.04667f
C703 VN.n13 VSUBS 0.04667f
C704 VN.n14 VSUBS 0.04667f
C705 VN.n15 VSUBS 0.068129f
C706 VN.n16 VSUBS 0.08698f
C707 VN.n17 VSUBS 0.082254f
C708 VN.n18 VSUBS 0.04667f
C709 VN.n19 VSUBS 0.04667f
C710 VN.n20 VSUBS 0.048759f
C711 VN.n21 VSUBS 0.08698f
C712 VN.n22 VSUBS 0.090467f
C713 VN.n23 VSUBS 0.04667f
C714 VN.n24 VSUBS 0.04667f
C715 VN.n25 VSUBS 0.04667f
C716 VN.n26 VSUBS 0.081802f
C717 VN.n27 VSUBS 0.08698f
C718 VN.n28 VSUBS 0.072807f
C719 VN.n29 VSUBS 0.075324f
C720 VN.n30 VSUBS 0.105273f
C721 VN.t2 VSUBS 0.911161f
C722 VN.n31 VSUBS 0.567584f
C723 VN.n32 VSUBS 0.04667f
C724 VN.n33 VSUBS 0.050969f
C725 VN.n34 VSUBS 0.04667f
C726 VN.t4 VSUBS 0.911161f
C727 VN.n35 VSUBS 0.391127f
C728 VN.n36 VSUBS 0.04667f
C729 VN.n37 VSUBS 0.068129f
C730 VN.n38 VSUBS 0.53345f
C731 VN.t5 VSUBS 0.911161f
C732 VN.t3 VSUBS 1.35193f
C733 VN.n39 VSUBS 0.539516f
C734 VN.n40 VSUBS 0.559191f
C735 VN.n41 VSUBS 0.082254f
C736 VN.n42 VSUBS 0.08698f
C737 VN.n43 VSUBS 0.04667f
C738 VN.n44 VSUBS 0.04667f
C739 VN.n45 VSUBS 0.04667f
C740 VN.n46 VSUBS 0.068129f
C741 VN.n47 VSUBS 0.08698f
C742 VN.n48 VSUBS 0.082254f
C743 VN.n49 VSUBS 0.04667f
C744 VN.n50 VSUBS 0.04667f
C745 VN.n51 VSUBS 0.048759f
C746 VN.n52 VSUBS 0.08698f
C747 VN.n53 VSUBS 0.090467f
C748 VN.n54 VSUBS 0.04667f
C749 VN.n55 VSUBS 0.04667f
C750 VN.n56 VSUBS 0.04667f
C751 VN.n57 VSUBS 0.081802f
C752 VN.n58 VSUBS 0.08698f
C753 VN.n59 VSUBS 0.072807f
C754 VN.n60 VSUBS 0.075324f
C755 VN.n61 VSUBS 2.36018f
C756 VDD1.t2 VSUBS 0.063871f
C757 VDD1.t3 VSUBS 0.063871f
C758 VDD1.n0 VSUBS 0.323027f
C759 VDD1.t0 VSUBS 0.063871f
C760 VDD1.t7 VSUBS 0.063871f
C761 VDD1.n1 VSUBS 0.322337f
C762 VDD1.t1 VSUBS 0.063871f
C763 VDD1.t6 VSUBS 0.063871f
C764 VDD1.n2 VSUBS 0.322337f
C765 VDD1.n3 VSUBS 3.98976f
C766 VDD1.t4 VSUBS 0.063871f
C767 VDD1.t5 VSUBS 0.063871f
C768 VDD1.n4 VSUBS 0.315036f
C769 VDD1.n5 VSUBS 3.10571f
C770 VTAIL.t1 VSUBS 0.07004f
C771 VTAIL.t7 VSUBS 0.07004f
C772 VTAIL.n0 VSUBS 0.297398f
C773 VTAIL.n1 VSUBS 0.735444f
C774 VTAIL.n2 VSUBS 0.037315f
C775 VTAIL.n3 VSUBS 0.251258f
C776 VTAIL.n4 VSUBS 0.018248f
C777 VTAIL.t2 VSUBS 0.098876f
C778 VTAIL.n5 VSUBS 0.116691f
C779 VTAIL.n6 VSUBS 0.025432f
C780 VTAIL.n7 VSUBS 0.032349f
C781 VTAIL.n8 VSUBS 0.104424f
C782 VTAIL.n9 VSUBS 0.019321f
C783 VTAIL.n10 VSUBS 0.018248f
C784 VTAIL.n11 VSUBS 0.088236f
C785 VTAIL.n12 VSUBS 0.052798f
C786 VTAIL.n13 VSUBS 0.405706f
C787 VTAIL.n14 VSUBS 0.037315f
C788 VTAIL.n15 VSUBS 0.251258f
C789 VTAIL.n16 VSUBS 0.018248f
C790 VTAIL.t12 VSUBS 0.098876f
C791 VTAIL.n17 VSUBS 0.116691f
C792 VTAIL.n18 VSUBS 0.025432f
C793 VTAIL.n19 VSUBS 0.032349f
C794 VTAIL.n20 VSUBS 0.104424f
C795 VTAIL.n21 VSUBS 0.019321f
C796 VTAIL.n22 VSUBS 0.018248f
C797 VTAIL.n23 VSUBS 0.088236f
C798 VTAIL.n24 VSUBS 0.052798f
C799 VTAIL.n25 VSUBS 0.405706f
C800 VTAIL.t13 VSUBS 0.07004f
C801 VTAIL.t14 VSUBS 0.07004f
C802 VTAIL.n26 VSUBS 0.297398f
C803 VTAIL.n27 VSUBS 1.04886f
C804 VTAIL.n28 VSUBS 0.037315f
C805 VTAIL.n29 VSUBS 0.251258f
C806 VTAIL.n30 VSUBS 0.018248f
C807 VTAIL.t10 VSUBS 0.098876f
C808 VTAIL.n31 VSUBS 0.116691f
C809 VTAIL.n32 VSUBS 0.025432f
C810 VTAIL.n33 VSUBS 0.032349f
C811 VTAIL.n34 VSUBS 0.104424f
C812 VTAIL.n35 VSUBS 0.019321f
C813 VTAIL.n36 VSUBS 0.018248f
C814 VTAIL.n37 VSUBS 0.088236f
C815 VTAIL.n38 VSUBS 0.052798f
C816 VTAIL.n39 VSUBS 1.38157f
C817 VTAIL.n40 VSUBS 0.037315f
C818 VTAIL.n41 VSUBS 0.251258f
C819 VTAIL.n42 VSUBS 0.018248f
C820 VTAIL.t0 VSUBS 0.098876f
C821 VTAIL.n43 VSUBS 0.116691f
C822 VTAIL.n44 VSUBS 0.025432f
C823 VTAIL.n45 VSUBS 0.032349f
C824 VTAIL.n46 VSUBS 0.104424f
C825 VTAIL.n47 VSUBS 0.019321f
C826 VTAIL.n48 VSUBS 0.018248f
C827 VTAIL.n49 VSUBS 0.088236f
C828 VTAIL.n50 VSUBS 0.052798f
C829 VTAIL.n51 VSUBS 1.38157f
C830 VTAIL.t5 VSUBS 0.07004f
C831 VTAIL.t6 VSUBS 0.07004f
C832 VTAIL.n52 VSUBS 0.297399f
C833 VTAIL.n53 VSUBS 1.04885f
C834 VTAIL.n54 VSUBS 0.037315f
C835 VTAIL.n55 VSUBS 0.251258f
C836 VTAIL.n56 VSUBS 0.018248f
C837 VTAIL.t4 VSUBS 0.098876f
C838 VTAIL.n57 VSUBS 0.116691f
C839 VTAIL.n58 VSUBS 0.025432f
C840 VTAIL.n59 VSUBS 0.032349f
C841 VTAIL.n60 VSUBS 0.104424f
C842 VTAIL.n61 VSUBS 0.019321f
C843 VTAIL.n62 VSUBS 0.018248f
C844 VTAIL.n63 VSUBS 0.088236f
C845 VTAIL.n64 VSUBS 0.052798f
C846 VTAIL.n65 VSUBS 0.405706f
C847 VTAIL.n66 VSUBS 0.037315f
C848 VTAIL.n67 VSUBS 0.251258f
C849 VTAIL.n68 VSUBS 0.018248f
C850 VTAIL.t8 VSUBS 0.098876f
C851 VTAIL.n69 VSUBS 0.116691f
C852 VTAIL.n70 VSUBS 0.025432f
C853 VTAIL.n71 VSUBS 0.032349f
C854 VTAIL.n72 VSUBS 0.104424f
C855 VTAIL.n73 VSUBS 0.019321f
C856 VTAIL.n74 VSUBS 0.018248f
C857 VTAIL.n75 VSUBS 0.088236f
C858 VTAIL.n76 VSUBS 0.052798f
C859 VTAIL.n77 VSUBS 0.405706f
C860 VTAIL.t15 VSUBS 0.07004f
C861 VTAIL.t11 VSUBS 0.07004f
C862 VTAIL.n78 VSUBS 0.297399f
C863 VTAIL.n79 VSUBS 1.04885f
C864 VTAIL.n80 VSUBS 0.037315f
C865 VTAIL.n81 VSUBS 0.251258f
C866 VTAIL.n82 VSUBS 0.018248f
C867 VTAIL.t9 VSUBS 0.098876f
C868 VTAIL.n83 VSUBS 0.116691f
C869 VTAIL.n84 VSUBS 0.025432f
C870 VTAIL.n85 VSUBS 0.032349f
C871 VTAIL.n86 VSUBS 0.104424f
C872 VTAIL.n87 VSUBS 0.019321f
C873 VTAIL.n88 VSUBS 0.018248f
C874 VTAIL.n89 VSUBS 0.088236f
C875 VTAIL.n90 VSUBS 0.052798f
C876 VTAIL.n91 VSUBS 1.38157f
C877 VTAIL.n92 VSUBS 0.037315f
C878 VTAIL.n93 VSUBS 0.251258f
C879 VTAIL.n94 VSUBS 0.018248f
C880 VTAIL.t3 VSUBS 0.098876f
C881 VTAIL.n95 VSUBS 0.116691f
C882 VTAIL.n96 VSUBS 0.025432f
C883 VTAIL.n97 VSUBS 0.032349f
C884 VTAIL.n98 VSUBS 0.104424f
C885 VTAIL.n99 VSUBS 0.019321f
C886 VTAIL.n100 VSUBS 0.018248f
C887 VTAIL.n101 VSUBS 0.088236f
C888 VTAIL.n102 VSUBS 0.052798f
C889 VTAIL.n103 VSUBS 1.3752f
C890 VP.t1 VSUBS 1.047f
C891 VP.n0 VSUBS 0.652199f
C892 VP.n1 VSUBS 0.053627f
C893 VP.n2 VSUBS 0.058568f
C894 VP.n3 VSUBS 0.053627f
C895 VP.t6 VSUBS 1.047f
C896 VP.n4 VSUBS 0.449436f
C897 VP.n5 VSUBS 0.053627f
C898 VP.n6 VSUBS 0.078286f
C899 VP.n7 VSUBS 0.053627f
C900 VP.t0 VSUBS 1.047f
C901 VP.n8 VSUBS 0.099947f
C902 VP.n9 VSUBS 0.053627f
C903 VP.n10 VSUBS 0.099947f
C904 VP.t2 VSUBS 1.047f
C905 VP.n11 VSUBS 0.652199f
C906 VP.n12 VSUBS 0.053627f
C907 VP.n13 VSUBS 0.058568f
C908 VP.n14 VSUBS 0.053627f
C909 VP.t3 VSUBS 1.047f
C910 VP.n15 VSUBS 0.449436f
C911 VP.n16 VSUBS 0.053627f
C912 VP.n17 VSUBS 0.078286f
C913 VP.n18 VSUBS 0.612977f
C914 VP.t4 VSUBS 1.047f
C915 VP.t5 VSUBS 1.55347f
C916 VP.n19 VSUBS 0.619947f
C917 VP.n20 VSUBS 0.642554f
C918 VP.n21 VSUBS 0.094517f
C919 VP.n22 VSUBS 0.099947f
C920 VP.n23 VSUBS 0.053627f
C921 VP.n24 VSUBS 0.053627f
C922 VP.n25 VSUBS 0.053627f
C923 VP.n26 VSUBS 0.078286f
C924 VP.n27 VSUBS 0.099947f
C925 VP.n28 VSUBS 0.094517f
C926 VP.n29 VSUBS 0.053627f
C927 VP.n30 VSUBS 0.053627f
C928 VP.n31 VSUBS 0.056028f
C929 VP.n32 VSUBS 0.099947f
C930 VP.n33 VSUBS 0.103954f
C931 VP.n34 VSUBS 0.053627f
C932 VP.n35 VSUBS 0.053627f
C933 VP.n36 VSUBS 0.053627f
C934 VP.n37 VSUBS 0.093997f
C935 VP.n38 VSUBS 0.099947f
C936 VP.n39 VSUBS 0.083661f
C937 VP.n40 VSUBS 0.086553f
C938 VP.n41 VSUBS 2.68943f
C939 VP.n42 VSUBS 2.73132f
C940 VP.t7 VSUBS 1.047f
C941 VP.n43 VSUBS 0.652199f
C942 VP.n44 VSUBS 0.083661f
C943 VP.n45 VSUBS 0.086553f
C944 VP.n46 VSUBS 0.053627f
C945 VP.n47 VSUBS 0.053627f
C946 VP.n48 VSUBS 0.093997f
C947 VP.n49 VSUBS 0.058568f
C948 VP.n50 VSUBS 0.103954f
C949 VP.n51 VSUBS 0.053627f
C950 VP.n52 VSUBS 0.053627f
C951 VP.n53 VSUBS 0.053627f
C952 VP.n54 VSUBS 0.056028f
C953 VP.n55 VSUBS 0.449436f
C954 VP.n56 VSUBS 0.094517f
C955 VP.n57 VSUBS 0.099947f
C956 VP.n58 VSUBS 0.053627f
C957 VP.n59 VSUBS 0.053627f
C958 VP.n60 VSUBS 0.053627f
C959 VP.n61 VSUBS 0.078286f
C960 VP.n62 VSUBS 0.099947f
C961 VP.n63 VSUBS 0.094517f
C962 VP.n64 VSUBS 0.053627f
C963 VP.n65 VSUBS 0.053627f
C964 VP.n66 VSUBS 0.056028f
C965 VP.n67 VSUBS 0.099947f
C966 VP.n68 VSUBS 0.103954f
C967 VP.n69 VSUBS 0.053627f
C968 VP.n70 VSUBS 0.053627f
C969 VP.n71 VSUBS 0.053627f
C970 VP.n72 VSUBS 0.093997f
C971 VP.n73 VSUBS 0.099947f
C972 VP.n74 VSUBS 0.083661f
C973 VP.n75 VSUBS 0.086553f
C974 VP.n76 VSUBS 0.120967f
.ends

