* NGSPICE file created from diff_pair_sample_0272.ext - technology: sky130A

.subckt diff_pair_sample_0272 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t3 VN.t0 VTAIL.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=0.9075 pd=5.83 as=2.145 ps=11.78 w=5.5 l=3.59
X1 VDD1.t3 VP.t0 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.9075 pd=5.83 as=2.145 ps=11.78 w=5.5 l=3.59
X2 VTAIL.t3 VP.t1 VDD1.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=2.145 pd=11.78 as=0.9075 ps=5.83 w=5.5 l=3.59
X3 B.t17 B.t15 B.t16 B.t12 sky130_fd_pr__nfet_01v8 ad=2.145 pd=11.78 as=0 ps=0 w=5.5 l=3.59
X4 VTAIL.t4 VN.t1 VDD2.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=2.145 pd=11.78 as=0.9075 ps=5.83 w=5.5 l=3.59
X5 B.t14 B.t11 B.t13 B.t12 sky130_fd_pr__nfet_01v8 ad=2.145 pd=11.78 as=0 ps=0 w=5.5 l=3.59
X6 VTAIL.t0 VP.t2 VDD1.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=2.145 pd=11.78 as=0.9075 ps=5.83 w=5.5 l=3.59
X7 VDD2.t1 VN.t2 VTAIL.t5 B.t1 sky130_fd_pr__nfet_01v8 ad=0.9075 pd=5.83 as=2.145 ps=11.78 w=5.5 l=3.59
X8 B.t10 B.t8 B.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=2.145 pd=11.78 as=0 ps=0 w=5.5 l=3.59
X9 VDD1.t0 VP.t3 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.9075 pd=5.83 as=2.145 ps=11.78 w=5.5 l=3.59
X10 VTAIL.t7 VN.t3 VDD2.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.145 pd=11.78 as=0.9075 ps=5.83 w=5.5 l=3.59
X11 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=2.145 pd=11.78 as=0 ps=0 w=5.5 l=3.59
R0 VN.n1 VN.t2 71.8345
R1 VN.n0 VN.t3 71.8345
R2 VN.n0 VN.t0 70.5919
R3 VN.n1 VN.t1 70.5919
R4 VN VN.n1 46.7794
R5 VN VN.n0 2.10136
R6 VTAIL.n5 VTAIL.t0 58.1546
R7 VTAIL.n4 VTAIL.t5 58.1546
R8 VTAIL.n3 VTAIL.t4 58.1546
R9 VTAIL.n6 VTAIL.t2 58.1537
R10 VTAIL.n7 VTAIL.t6 58.1536
R11 VTAIL.n0 VTAIL.t7 58.1536
R12 VTAIL.n1 VTAIL.t1 58.1536
R13 VTAIL.n2 VTAIL.t3 58.1536
R14 VTAIL.n7 VTAIL.n6 20.4876
R15 VTAIL.n3 VTAIL.n2 20.4876
R16 VTAIL.n4 VTAIL.n3 3.37981
R17 VTAIL.n6 VTAIL.n5 3.37981
R18 VTAIL.n2 VTAIL.n1 3.37981
R19 VTAIL VTAIL.n0 1.74834
R20 VTAIL VTAIL.n7 1.63197
R21 VTAIL.n5 VTAIL.n4 0.470328
R22 VTAIL.n1 VTAIL.n0 0.470328
R23 VDD2.n2 VDD2.n0 109.828
R24 VDD2.n2 VDD2.n1 71.2325
R25 VDD2.n1 VDD2.t2 3.6005
R26 VDD2.n1 VDD2.t1 3.6005
R27 VDD2.n0 VDD2.t0 3.6005
R28 VDD2.n0 VDD2.t3 3.6005
R29 VDD2 VDD2.n2 0.0586897
R30 B.n519 B.n518 585
R31 B.n519 B.n79 585
R32 B.n522 B.n521 585
R33 B.n523 B.n111 585
R34 B.n525 B.n524 585
R35 B.n527 B.n110 585
R36 B.n530 B.n529 585
R37 B.n531 B.n109 585
R38 B.n533 B.n532 585
R39 B.n535 B.n108 585
R40 B.n538 B.n537 585
R41 B.n539 B.n107 585
R42 B.n541 B.n540 585
R43 B.n543 B.n106 585
R44 B.n546 B.n545 585
R45 B.n547 B.n105 585
R46 B.n549 B.n548 585
R47 B.n551 B.n104 585
R48 B.n554 B.n553 585
R49 B.n555 B.n103 585
R50 B.n557 B.n556 585
R51 B.n559 B.n102 585
R52 B.n562 B.n561 585
R53 B.n563 B.n99 585
R54 B.n566 B.n565 585
R55 B.n568 B.n98 585
R56 B.n571 B.n570 585
R57 B.n572 B.n97 585
R58 B.n574 B.n573 585
R59 B.n576 B.n96 585
R60 B.n579 B.n578 585
R61 B.n580 B.n92 585
R62 B.n582 B.n581 585
R63 B.n584 B.n91 585
R64 B.n587 B.n586 585
R65 B.n588 B.n90 585
R66 B.n590 B.n589 585
R67 B.n592 B.n89 585
R68 B.n595 B.n594 585
R69 B.n596 B.n88 585
R70 B.n598 B.n597 585
R71 B.n600 B.n87 585
R72 B.n603 B.n602 585
R73 B.n604 B.n86 585
R74 B.n606 B.n605 585
R75 B.n608 B.n85 585
R76 B.n611 B.n610 585
R77 B.n612 B.n84 585
R78 B.n614 B.n613 585
R79 B.n616 B.n83 585
R80 B.n619 B.n618 585
R81 B.n620 B.n82 585
R82 B.n622 B.n621 585
R83 B.n624 B.n81 585
R84 B.n627 B.n626 585
R85 B.n628 B.n80 585
R86 B.n517 B.n78 585
R87 B.n631 B.n78 585
R88 B.n516 B.n77 585
R89 B.n632 B.n77 585
R90 B.n515 B.n76 585
R91 B.n633 B.n76 585
R92 B.n514 B.n513 585
R93 B.n513 B.n72 585
R94 B.n512 B.n71 585
R95 B.n639 B.n71 585
R96 B.n511 B.n70 585
R97 B.n640 B.n70 585
R98 B.n510 B.n69 585
R99 B.n641 B.n69 585
R100 B.n509 B.n508 585
R101 B.n508 B.n65 585
R102 B.n507 B.n64 585
R103 B.n647 B.n64 585
R104 B.n506 B.n63 585
R105 B.n648 B.n63 585
R106 B.n505 B.n62 585
R107 B.n649 B.n62 585
R108 B.n504 B.n503 585
R109 B.n503 B.n58 585
R110 B.n502 B.n57 585
R111 B.n655 B.n57 585
R112 B.n501 B.n56 585
R113 B.n656 B.n56 585
R114 B.n500 B.n55 585
R115 B.n657 B.n55 585
R116 B.n499 B.n498 585
R117 B.n498 B.n51 585
R118 B.n497 B.n50 585
R119 B.n663 B.n50 585
R120 B.n496 B.n49 585
R121 B.n664 B.n49 585
R122 B.n495 B.n48 585
R123 B.n665 B.n48 585
R124 B.n494 B.n493 585
R125 B.n493 B.n44 585
R126 B.n492 B.n43 585
R127 B.n671 B.n43 585
R128 B.n491 B.n42 585
R129 B.n672 B.n42 585
R130 B.n490 B.n41 585
R131 B.n673 B.n41 585
R132 B.n489 B.n488 585
R133 B.n488 B.n40 585
R134 B.n487 B.n36 585
R135 B.n679 B.n36 585
R136 B.n486 B.n35 585
R137 B.n680 B.n35 585
R138 B.n485 B.n34 585
R139 B.n681 B.n34 585
R140 B.n484 B.n483 585
R141 B.n483 B.n30 585
R142 B.n482 B.n29 585
R143 B.n687 B.n29 585
R144 B.n481 B.n28 585
R145 B.n688 B.n28 585
R146 B.n480 B.n27 585
R147 B.n689 B.n27 585
R148 B.n479 B.n478 585
R149 B.n478 B.n23 585
R150 B.n477 B.n22 585
R151 B.n695 B.n22 585
R152 B.n476 B.n21 585
R153 B.n696 B.n21 585
R154 B.n475 B.n20 585
R155 B.n697 B.n20 585
R156 B.n474 B.n473 585
R157 B.n473 B.n19 585
R158 B.n472 B.n15 585
R159 B.n703 B.n15 585
R160 B.n471 B.n14 585
R161 B.n704 B.n14 585
R162 B.n470 B.n13 585
R163 B.n705 B.n13 585
R164 B.n469 B.n468 585
R165 B.n468 B.n12 585
R166 B.n467 B.n466 585
R167 B.n467 B.n8 585
R168 B.n465 B.n7 585
R169 B.n712 B.n7 585
R170 B.n464 B.n6 585
R171 B.n713 B.n6 585
R172 B.n463 B.n5 585
R173 B.n714 B.n5 585
R174 B.n462 B.n461 585
R175 B.n461 B.n4 585
R176 B.n460 B.n112 585
R177 B.n460 B.n459 585
R178 B.n450 B.n113 585
R179 B.n114 B.n113 585
R180 B.n452 B.n451 585
R181 B.n453 B.n452 585
R182 B.n449 B.n119 585
R183 B.n119 B.n118 585
R184 B.n448 B.n447 585
R185 B.n447 B.n446 585
R186 B.n121 B.n120 585
R187 B.n439 B.n121 585
R188 B.n438 B.n437 585
R189 B.n440 B.n438 585
R190 B.n436 B.n126 585
R191 B.n126 B.n125 585
R192 B.n435 B.n434 585
R193 B.n434 B.n433 585
R194 B.n128 B.n127 585
R195 B.n129 B.n128 585
R196 B.n426 B.n425 585
R197 B.n427 B.n426 585
R198 B.n424 B.n134 585
R199 B.n134 B.n133 585
R200 B.n423 B.n422 585
R201 B.n422 B.n421 585
R202 B.n136 B.n135 585
R203 B.n137 B.n136 585
R204 B.n414 B.n413 585
R205 B.n415 B.n414 585
R206 B.n412 B.n142 585
R207 B.n142 B.n141 585
R208 B.n411 B.n410 585
R209 B.n410 B.n409 585
R210 B.n144 B.n143 585
R211 B.n402 B.n144 585
R212 B.n401 B.n400 585
R213 B.n403 B.n401 585
R214 B.n399 B.n149 585
R215 B.n149 B.n148 585
R216 B.n398 B.n397 585
R217 B.n397 B.n396 585
R218 B.n151 B.n150 585
R219 B.n152 B.n151 585
R220 B.n389 B.n388 585
R221 B.n390 B.n389 585
R222 B.n387 B.n157 585
R223 B.n157 B.n156 585
R224 B.n386 B.n385 585
R225 B.n385 B.n384 585
R226 B.n159 B.n158 585
R227 B.n160 B.n159 585
R228 B.n377 B.n376 585
R229 B.n378 B.n377 585
R230 B.n375 B.n165 585
R231 B.n165 B.n164 585
R232 B.n374 B.n373 585
R233 B.n373 B.n372 585
R234 B.n167 B.n166 585
R235 B.n168 B.n167 585
R236 B.n365 B.n364 585
R237 B.n366 B.n365 585
R238 B.n363 B.n173 585
R239 B.n173 B.n172 585
R240 B.n362 B.n361 585
R241 B.n361 B.n360 585
R242 B.n175 B.n174 585
R243 B.n176 B.n175 585
R244 B.n353 B.n352 585
R245 B.n354 B.n353 585
R246 B.n351 B.n181 585
R247 B.n181 B.n180 585
R248 B.n350 B.n349 585
R249 B.n349 B.n348 585
R250 B.n183 B.n182 585
R251 B.n184 B.n183 585
R252 B.n341 B.n340 585
R253 B.n342 B.n341 585
R254 B.n339 B.n189 585
R255 B.n189 B.n188 585
R256 B.n338 B.n337 585
R257 B.n337 B.n336 585
R258 B.n333 B.n193 585
R259 B.n332 B.n331 585
R260 B.n329 B.n194 585
R261 B.n329 B.n192 585
R262 B.n328 B.n327 585
R263 B.n326 B.n325 585
R264 B.n324 B.n196 585
R265 B.n322 B.n321 585
R266 B.n320 B.n197 585
R267 B.n319 B.n318 585
R268 B.n316 B.n198 585
R269 B.n314 B.n313 585
R270 B.n312 B.n199 585
R271 B.n311 B.n310 585
R272 B.n308 B.n200 585
R273 B.n306 B.n305 585
R274 B.n304 B.n201 585
R275 B.n303 B.n302 585
R276 B.n300 B.n202 585
R277 B.n298 B.n297 585
R278 B.n296 B.n203 585
R279 B.n295 B.n294 585
R280 B.n292 B.n204 585
R281 B.n290 B.n289 585
R282 B.n287 B.n205 585
R283 B.n286 B.n285 585
R284 B.n283 B.n208 585
R285 B.n281 B.n280 585
R286 B.n279 B.n209 585
R287 B.n278 B.n277 585
R288 B.n275 B.n210 585
R289 B.n273 B.n272 585
R290 B.n271 B.n211 585
R291 B.n269 B.n268 585
R292 B.n266 B.n214 585
R293 B.n264 B.n263 585
R294 B.n262 B.n215 585
R295 B.n261 B.n260 585
R296 B.n258 B.n216 585
R297 B.n256 B.n255 585
R298 B.n254 B.n217 585
R299 B.n253 B.n252 585
R300 B.n250 B.n218 585
R301 B.n248 B.n247 585
R302 B.n246 B.n219 585
R303 B.n245 B.n244 585
R304 B.n242 B.n220 585
R305 B.n240 B.n239 585
R306 B.n238 B.n221 585
R307 B.n237 B.n236 585
R308 B.n234 B.n222 585
R309 B.n232 B.n231 585
R310 B.n230 B.n223 585
R311 B.n229 B.n228 585
R312 B.n226 B.n224 585
R313 B.n191 B.n190 585
R314 B.n335 B.n334 585
R315 B.n336 B.n335 585
R316 B.n187 B.n186 585
R317 B.n188 B.n187 585
R318 B.n344 B.n343 585
R319 B.n343 B.n342 585
R320 B.n345 B.n185 585
R321 B.n185 B.n184 585
R322 B.n347 B.n346 585
R323 B.n348 B.n347 585
R324 B.n179 B.n178 585
R325 B.n180 B.n179 585
R326 B.n356 B.n355 585
R327 B.n355 B.n354 585
R328 B.n357 B.n177 585
R329 B.n177 B.n176 585
R330 B.n359 B.n358 585
R331 B.n360 B.n359 585
R332 B.n171 B.n170 585
R333 B.n172 B.n171 585
R334 B.n368 B.n367 585
R335 B.n367 B.n366 585
R336 B.n369 B.n169 585
R337 B.n169 B.n168 585
R338 B.n371 B.n370 585
R339 B.n372 B.n371 585
R340 B.n163 B.n162 585
R341 B.n164 B.n163 585
R342 B.n380 B.n379 585
R343 B.n379 B.n378 585
R344 B.n381 B.n161 585
R345 B.n161 B.n160 585
R346 B.n383 B.n382 585
R347 B.n384 B.n383 585
R348 B.n155 B.n154 585
R349 B.n156 B.n155 585
R350 B.n392 B.n391 585
R351 B.n391 B.n390 585
R352 B.n393 B.n153 585
R353 B.n153 B.n152 585
R354 B.n395 B.n394 585
R355 B.n396 B.n395 585
R356 B.n147 B.n146 585
R357 B.n148 B.n147 585
R358 B.n405 B.n404 585
R359 B.n404 B.n403 585
R360 B.n406 B.n145 585
R361 B.n402 B.n145 585
R362 B.n408 B.n407 585
R363 B.n409 B.n408 585
R364 B.n140 B.n139 585
R365 B.n141 B.n140 585
R366 B.n417 B.n416 585
R367 B.n416 B.n415 585
R368 B.n418 B.n138 585
R369 B.n138 B.n137 585
R370 B.n420 B.n419 585
R371 B.n421 B.n420 585
R372 B.n132 B.n131 585
R373 B.n133 B.n132 585
R374 B.n429 B.n428 585
R375 B.n428 B.n427 585
R376 B.n430 B.n130 585
R377 B.n130 B.n129 585
R378 B.n432 B.n431 585
R379 B.n433 B.n432 585
R380 B.n124 B.n123 585
R381 B.n125 B.n124 585
R382 B.n442 B.n441 585
R383 B.n441 B.n440 585
R384 B.n443 B.n122 585
R385 B.n439 B.n122 585
R386 B.n445 B.n444 585
R387 B.n446 B.n445 585
R388 B.n117 B.n116 585
R389 B.n118 B.n117 585
R390 B.n455 B.n454 585
R391 B.n454 B.n453 585
R392 B.n456 B.n115 585
R393 B.n115 B.n114 585
R394 B.n458 B.n457 585
R395 B.n459 B.n458 585
R396 B.n3 B.n0 585
R397 B.n4 B.n3 585
R398 B.n711 B.n1 585
R399 B.n712 B.n711 585
R400 B.n710 B.n709 585
R401 B.n710 B.n8 585
R402 B.n708 B.n9 585
R403 B.n12 B.n9 585
R404 B.n707 B.n706 585
R405 B.n706 B.n705 585
R406 B.n11 B.n10 585
R407 B.n704 B.n11 585
R408 B.n702 B.n701 585
R409 B.n703 B.n702 585
R410 B.n700 B.n16 585
R411 B.n19 B.n16 585
R412 B.n699 B.n698 585
R413 B.n698 B.n697 585
R414 B.n18 B.n17 585
R415 B.n696 B.n18 585
R416 B.n694 B.n693 585
R417 B.n695 B.n694 585
R418 B.n692 B.n24 585
R419 B.n24 B.n23 585
R420 B.n691 B.n690 585
R421 B.n690 B.n689 585
R422 B.n26 B.n25 585
R423 B.n688 B.n26 585
R424 B.n686 B.n685 585
R425 B.n687 B.n686 585
R426 B.n684 B.n31 585
R427 B.n31 B.n30 585
R428 B.n683 B.n682 585
R429 B.n682 B.n681 585
R430 B.n33 B.n32 585
R431 B.n680 B.n33 585
R432 B.n678 B.n677 585
R433 B.n679 B.n678 585
R434 B.n676 B.n37 585
R435 B.n40 B.n37 585
R436 B.n675 B.n674 585
R437 B.n674 B.n673 585
R438 B.n39 B.n38 585
R439 B.n672 B.n39 585
R440 B.n670 B.n669 585
R441 B.n671 B.n670 585
R442 B.n668 B.n45 585
R443 B.n45 B.n44 585
R444 B.n667 B.n666 585
R445 B.n666 B.n665 585
R446 B.n47 B.n46 585
R447 B.n664 B.n47 585
R448 B.n662 B.n661 585
R449 B.n663 B.n662 585
R450 B.n660 B.n52 585
R451 B.n52 B.n51 585
R452 B.n659 B.n658 585
R453 B.n658 B.n657 585
R454 B.n54 B.n53 585
R455 B.n656 B.n54 585
R456 B.n654 B.n653 585
R457 B.n655 B.n654 585
R458 B.n652 B.n59 585
R459 B.n59 B.n58 585
R460 B.n651 B.n650 585
R461 B.n650 B.n649 585
R462 B.n61 B.n60 585
R463 B.n648 B.n61 585
R464 B.n646 B.n645 585
R465 B.n647 B.n646 585
R466 B.n644 B.n66 585
R467 B.n66 B.n65 585
R468 B.n643 B.n642 585
R469 B.n642 B.n641 585
R470 B.n68 B.n67 585
R471 B.n640 B.n68 585
R472 B.n638 B.n637 585
R473 B.n639 B.n638 585
R474 B.n636 B.n73 585
R475 B.n73 B.n72 585
R476 B.n635 B.n634 585
R477 B.n634 B.n633 585
R478 B.n75 B.n74 585
R479 B.n632 B.n75 585
R480 B.n630 B.n629 585
R481 B.n631 B.n630 585
R482 B.n715 B.n714 585
R483 B.n713 B.n2 585
R484 B.n630 B.n80 497.305
R485 B.n519 B.n78 497.305
R486 B.n337 B.n191 497.305
R487 B.n335 B.n193 497.305
R488 B.n520 B.n79 256.663
R489 B.n526 B.n79 256.663
R490 B.n528 B.n79 256.663
R491 B.n534 B.n79 256.663
R492 B.n536 B.n79 256.663
R493 B.n542 B.n79 256.663
R494 B.n544 B.n79 256.663
R495 B.n550 B.n79 256.663
R496 B.n552 B.n79 256.663
R497 B.n558 B.n79 256.663
R498 B.n560 B.n79 256.663
R499 B.n567 B.n79 256.663
R500 B.n569 B.n79 256.663
R501 B.n575 B.n79 256.663
R502 B.n577 B.n79 256.663
R503 B.n583 B.n79 256.663
R504 B.n585 B.n79 256.663
R505 B.n591 B.n79 256.663
R506 B.n593 B.n79 256.663
R507 B.n599 B.n79 256.663
R508 B.n601 B.n79 256.663
R509 B.n607 B.n79 256.663
R510 B.n609 B.n79 256.663
R511 B.n615 B.n79 256.663
R512 B.n617 B.n79 256.663
R513 B.n623 B.n79 256.663
R514 B.n625 B.n79 256.663
R515 B.n330 B.n192 256.663
R516 B.n195 B.n192 256.663
R517 B.n323 B.n192 256.663
R518 B.n317 B.n192 256.663
R519 B.n315 B.n192 256.663
R520 B.n309 B.n192 256.663
R521 B.n307 B.n192 256.663
R522 B.n301 B.n192 256.663
R523 B.n299 B.n192 256.663
R524 B.n293 B.n192 256.663
R525 B.n291 B.n192 256.663
R526 B.n284 B.n192 256.663
R527 B.n282 B.n192 256.663
R528 B.n276 B.n192 256.663
R529 B.n274 B.n192 256.663
R530 B.n267 B.n192 256.663
R531 B.n265 B.n192 256.663
R532 B.n259 B.n192 256.663
R533 B.n257 B.n192 256.663
R534 B.n251 B.n192 256.663
R535 B.n249 B.n192 256.663
R536 B.n243 B.n192 256.663
R537 B.n241 B.n192 256.663
R538 B.n235 B.n192 256.663
R539 B.n233 B.n192 256.663
R540 B.n227 B.n192 256.663
R541 B.n225 B.n192 256.663
R542 B.n717 B.n716 256.663
R543 B.n93 B.t15 246.095
R544 B.n100 B.t11 246.095
R545 B.n212 B.t8 246.095
R546 B.n206 B.t4 246.095
R547 B.n626 B.n624 163.367
R548 B.n622 B.n82 163.367
R549 B.n618 B.n616 163.367
R550 B.n614 B.n84 163.367
R551 B.n610 B.n608 163.367
R552 B.n606 B.n86 163.367
R553 B.n602 B.n600 163.367
R554 B.n598 B.n88 163.367
R555 B.n594 B.n592 163.367
R556 B.n590 B.n90 163.367
R557 B.n586 B.n584 163.367
R558 B.n582 B.n92 163.367
R559 B.n578 B.n576 163.367
R560 B.n574 B.n97 163.367
R561 B.n570 B.n568 163.367
R562 B.n566 B.n99 163.367
R563 B.n561 B.n559 163.367
R564 B.n557 B.n103 163.367
R565 B.n553 B.n551 163.367
R566 B.n549 B.n105 163.367
R567 B.n545 B.n543 163.367
R568 B.n541 B.n107 163.367
R569 B.n537 B.n535 163.367
R570 B.n533 B.n109 163.367
R571 B.n529 B.n527 163.367
R572 B.n525 B.n111 163.367
R573 B.n521 B.n519 163.367
R574 B.n337 B.n189 163.367
R575 B.n341 B.n189 163.367
R576 B.n341 B.n183 163.367
R577 B.n349 B.n183 163.367
R578 B.n349 B.n181 163.367
R579 B.n353 B.n181 163.367
R580 B.n353 B.n175 163.367
R581 B.n361 B.n175 163.367
R582 B.n361 B.n173 163.367
R583 B.n365 B.n173 163.367
R584 B.n365 B.n167 163.367
R585 B.n373 B.n167 163.367
R586 B.n373 B.n165 163.367
R587 B.n377 B.n165 163.367
R588 B.n377 B.n159 163.367
R589 B.n385 B.n159 163.367
R590 B.n385 B.n157 163.367
R591 B.n389 B.n157 163.367
R592 B.n389 B.n151 163.367
R593 B.n397 B.n151 163.367
R594 B.n397 B.n149 163.367
R595 B.n401 B.n149 163.367
R596 B.n401 B.n144 163.367
R597 B.n410 B.n144 163.367
R598 B.n410 B.n142 163.367
R599 B.n414 B.n142 163.367
R600 B.n414 B.n136 163.367
R601 B.n422 B.n136 163.367
R602 B.n422 B.n134 163.367
R603 B.n426 B.n134 163.367
R604 B.n426 B.n128 163.367
R605 B.n434 B.n128 163.367
R606 B.n434 B.n126 163.367
R607 B.n438 B.n126 163.367
R608 B.n438 B.n121 163.367
R609 B.n447 B.n121 163.367
R610 B.n447 B.n119 163.367
R611 B.n452 B.n119 163.367
R612 B.n452 B.n113 163.367
R613 B.n460 B.n113 163.367
R614 B.n461 B.n460 163.367
R615 B.n461 B.n5 163.367
R616 B.n6 B.n5 163.367
R617 B.n7 B.n6 163.367
R618 B.n467 B.n7 163.367
R619 B.n468 B.n467 163.367
R620 B.n468 B.n13 163.367
R621 B.n14 B.n13 163.367
R622 B.n15 B.n14 163.367
R623 B.n473 B.n15 163.367
R624 B.n473 B.n20 163.367
R625 B.n21 B.n20 163.367
R626 B.n22 B.n21 163.367
R627 B.n478 B.n22 163.367
R628 B.n478 B.n27 163.367
R629 B.n28 B.n27 163.367
R630 B.n29 B.n28 163.367
R631 B.n483 B.n29 163.367
R632 B.n483 B.n34 163.367
R633 B.n35 B.n34 163.367
R634 B.n36 B.n35 163.367
R635 B.n488 B.n36 163.367
R636 B.n488 B.n41 163.367
R637 B.n42 B.n41 163.367
R638 B.n43 B.n42 163.367
R639 B.n493 B.n43 163.367
R640 B.n493 B.n48 163.367
R641 B.n49 B.n48 163.367
R642 B.n50 B.n49 163.367
R643 B.n498 B.n50 163.367
R644 B.n498 B.n55 163.367
R645 B.n56 B.n55 163.367
R646 B.n57 B.n56 163.367
R647 B.n503 B.n57 163.367
R648 B.n503 B.n62 163.367
R649 B.n63 B.n62 163.367
R650 B.n64 B.n63 163.367
R651 B.n508 B.n64 163.367
R652 B.n508 B.n69 163.367
R653 B.n70 B.n69 163.367
R654 B.n71 B.n70 163.367
R655 B.n513 B.n71 163.367
R656 B.n513 B.n76 163.367
R657 B.n77 B.n76 163.367
R658 B.n78 B.n77 163.367
R659 B.n331 B.n329 163.367
R660 B.n329 B.n328 163.367
R661 B.n325 B.n324 163.367
R662 B.n322 B.n197 163.367
R663 B.n318 B.n316 163.367
R664 B.n314 B.n199 163.367
R665 B.n310 B.n308 163.367
R666 B.n306 B.n201 163.367
R667 B.n302 B.n300 163.367
R668 B.n298 B.n203 163.367
R669 B.n294 B.n292 163.367
R670 B.n290 B.n205 163.367
R671 B.n285 B.n283 163.367
R672 B.n281 B.n209 163.367
R673 B.n277 B.n275 163.367
R674 B.n273 B.n211 163.367
R675 B.n268 B.n266 163.367
R676 B.n264 B.n215 163.367
R677 B.n260 B.n258 163.367
R678 B.n256 B.n217 163.367
R679 B.n252 B.n250 163.367
R680 B.n248 B.n219 163.367
R681 B.n244 B.n242 163.367
R682 B.n240 B.n221 163.367
R683 B.n236 B.n234 163.367
R684 B.n232 B.n223 163.367
R685 B.n228 B.n226 163.367
R686 B.n335 B.n187 163.367
R687 B.n343 B.n187 163.367
R688 B.n343 B.n185 163.367
R689 B.n347 B.n185 163.367
R690 B.n347 B.n179 163.367
R691 B.n355 B.n179 163.367
R692 B.n355 B.n177 163.367
R693 B.n359 B.n177 163.367
R694 B.n359 B.n171 163.367
R695 B.n367 B.n171 163.367
R696 B.n367 B.n169 163.367
R697 B.n371 B.n169 163.367
R698 B.n371 B.n163 163.367
R699 B.n379 B.n163 163.367
R700 B.n379 B.n161 163.367
R701 B.n383 B.n161 163.367
R702 B.n383 B.n155 163.367
R703 B.n391 B.n155 163.367
R704 B.n391 B.n153 163.367
R705 B.n395 B.n153 163.367
R706 B.n395 B.n147 163.367
R707 B.n404 B.n147 163.367
R708 B.n404 B.n145 163.367
R709 B.n408 B.n145 163.367
R710 B.n408 B.n140 163.367
R711 B.n416 B.n140 163.367
R712 B.n416 B.n138 163.367
R713 B.n420 B.n138 163.367
R714 B.n420 B.n132 163.367
R715 B.n428 B.n132 163.367
R716 B.n428 B.n130 163.367
R717 B.n432 B.n130 163.367
R718 B.n432 B.n124 163.367
R719 B.n441 B.n124 163.367
R720 B.n441 B.n122 163.367
R721 B.n445 B.n122 163.367
R722 B.n445 B.n117 163.367
R723 B.n454 B.n117 163.367
R724 B.n454 B.n115 163.367
R725 B.n458 B.n115 163.367
R726 B.n458 B.n3 163.367
R727 B.n715 B.n3 163.367
R728 B.n711 B.n2 163.367
R729 B.n711 B.n710 163.367
R730 B.n710 B.n9 163.367
R731 B.n706 B.n9 163.367
R732 B.n706 B.n11 163.367
R733 B.n702 B.n11 163.367
R734 B.n702 B.n16 163.367
R735 B.n698 B.n16 163.367
R736 B.n698 B.n18 163.367
R737 B.n694 B.n18 163.367
R738 B.n694 B.n24 163.367
R739 B.n690 B.n24 163.367
R740 B.n690 B.n26 163.367
R741 B.n686 B.n26 163.367
R742 B.n686 B.n31 163.367
R743 B.n682 B.n31 163.367
R744 B.n682 B.n33 163.367
R745 B.n678 B.n33 163.367
R746 B.n678 B.n37 163.367
R747 B.n674 B.n37 163.367
R748 B.n674 B.n39 163.367
R749 B.n670 B.n39 163.367
R750 B.n670 B.n45 163.367
R751 B.n666 B.n45 163.367
R752 B.n666 B.n47 163.367
R753 B.n662 B.n47 163.367
R754 B.n662 B.n52 163.367
R755 B.n658 B.n52 163.367
R756 B.n658 B.n54 163.367
R757 B.n654 B.n54 163.367
R758 B.n654 B.n59 163.367
R759 B.n650 B.n59 163.367
R760 B.n650 B.n61 163.367
R761 B.n646 B.n61 163.367
R762 B.n646 B.n66 163.367
R763 B.n642 B.n66 163.367
R764 B.n642 B.n68 163.367
R765 B.n638 B.n68 163.367
R766 B.n638 B.n73 163.367
R767 B.n634 B.n73 163.367
R768 B.n634 B.n75 163.367
R769 B.n630 B.n75 163.367
R770 B.n100 B.t13 146.952
R771 B.n212 B.t10 146.952
R772 B.n93 B.t16 146.946
R773 B.n206 B.t7 146.946
R774 B.n336 B.n192 139.862
R775 B.n631 B.n79 139.862
R776 B.n94 B.n93 76.0247
R777 B.n101 B.n100 76.0247
R778 B.n213 B.n212 76.0247
R779 B.n207 B.n206 76.0247
R780 B.n625 B.n80 71.676
R781 B.n624 B.n623 71.676
R782 B.n617 B.n82 71.676
R783 B.n616 B.n615 71.676
R784 B.n609 B.n84 71.676
R785 B.n608 B.n607 71.676
R786 B.n601 B.n86 71.676
R787 B.n600 B.n599 71.676
R788 B.n593 B.n88 71.676
R789 B.n592 B.n591 71.676
R790 B.n585 B.n90 71.676
R791 B.n584 B.n583 71.676
R792 B.n577 B.n92 71.676
R793 B.n576 B.n575 71.676
R794 B.n569 B.n97 71.676
R795 B.n568 B.n567 71.676
R796 B.n560 B.n99 71.676
R797 B.n559 B.n558 71.676
R798 B.n552 B.n103 71.676
R799 B.n551 B.n550 71.676
R800 B.n544 B.n105 71.676
R801 B.n543 B.n542 71.676
R802 B.n536 B.n107 71.676
R803 B.n535 B.n534 71.676
R804 B.n528 B.n109 71.676
R805 B.n527 B.n526 71.676
R806 B.n520 B.n111 71.676
R807 B.n521 B.n520 71.676
R808 B.n526 B.n525 71.676
R809 B.n529 B.n528 71.676
R810 B.n534 B.n533 71.676
R811 B.n537 B.n536 71.676
R812 B.n542 B.n541 71.676
R813 B.n545 B.n544 71.676
R814 B.n550 B.n549 71.676
R815 B.n553 B.n552 71.676
R816 B.n558 B.n557 71.676
R817 B.n561 B.n560 71.676
R818 B.n567 B.n566 71.676
R819 B.n570 B.n569 71.676
R820 B.n575 B.n574 71.676
R821 B.n578 B.n577 71.676
R822 B.n583 B.n582 71.676
R823 B.n586 B.n585 71.676
R824 B.n591 B.n590 71.676
R825 B.n594 B.n593 71.676
R826 B.n599 B.n598 71.676
R827 B.n602 B.n601 71.676
R828 B.n607 B.n606 71.676
R829 B.n610 B.n609 71.676
R830 B.n615 B.n614 71.676
R831 B.n618 B.n617 71.676
R832 B.n623 B.n622 71.676
R833 B.n626 B.n625 71.676
R834 B.n330 B.n193 71.676
R835 B.n328 B.n195 71.676
R836 B.n324 B.n323 71.676
R837 B.n317 B.n197 71.676
R838 B.n316 B.n315 71.676
R839 B.n309 B.n199 71.676
R840 B.n308 B.n307 71.676
R841 B.n301 B.n201 71.676
R842 B.n300 B.n299 71.676
R843 B.n293 B.n203 71.676
R844 B.n292 B.n291 71.676
R845 B.n284 B.n205 71.676
R846 B.n283 B.n282 71.676
R847 B.n276 B.n209 71.676
R848 B.n275 B.n274 71.676
R849 B.n267 B.n211 71.676
R850 B.n266 B.n265 71.676
R851 B.n259 B.n215 71.676
R852 B.n258 B.n257 71.676
R853 B.n251 B.n217 71.676
R854 B.n250 B.n249 71.676
R855 B.n243 B.n219 71.676
R856 B.n242 B.n241 71.676
R857 B.n235 B.n221 71.676
R858 B.n234 B.n233 71.676
R859 B.n227 B.n223 71.676
R860 B.n226 B.n225 71.676
R861 B.n331 B.n330 71.676
R862 B.n325 B.n195 71.676
R863 B.n323 B.n322 71.676
R864 B.n318 B.n317 71.676
R865 B.n315 B.n314 71.676
R866 B.n310 B.n309 71.676
R867 B.n307 B.n306 71.676
R868 B.n302 B.n301 71.676
R869 B.n299 B.n298 71.676
R870 B.n294 B.n293 71.676
R871 B.n291 B.n290 71.676
R872 B.n285 B.n284 71.676
R873 B.n282 B.n281 71.676
R874 B.n277 B.n276 71.676
R875 B.n274 B.n273 71.676
R876 B.n268 B.n267 71.676
R877 B.n265 B.n264 71.676
R878 B.n260 B.n259 71.676
R879 B.n257 B.n256 71.676
R880 B.n252 B.n251 71.676
R881 B.n249 B.n248 71.676
R882 B.n244 B.n243 71.676
R883 B.n241 B.n240 71.676
R884 B.n236 B.n235 71.676
R885 B.n233 B.n232 71.676
R886 B.n228 B.n227 71.676
R887 B.n225 B.n191 71.676
R888 B.n716 B.n715 71.676
R889 B.n716 B.n2 71.676
R890 B.n101 B.t14 70.928
R891 B.n213 B.t9 70.928
R892 B.n94 B.t17 70.9222
R893 B.n207 B.t6 70.9222
R894 B.n336 B.n188 69.4205
R895 B.n342 B.n188 69.4205
R896 B.n342 B.n184 69.4205
R897 B.n348 B.n184 69.4205
R898 B.n348 B.n180 69.4205
R899 B.n354 B.n180 69.4205
R900 B.n354 B.n176 69.4205
R901 B.n360 B.n176 69.4205
R902 B.n366 B.n172 69.4205
R903 B.n366 B.n168 69.4205
R904 B.n372 B.n168 69.4205
R905 B.n372 B.n164 69.4205
R906 B.n378 B.n164 69.4205
R907 B.n378 B.n160 69.4205
R908 B.n384 B.n160 69.4205
R909 B.n384 B.n156 69.4205
R910 B.n390 B.n156 69.4205
R911 B.n390 B.n152 69.4205
R912 B.n396 B.n152 69.4205
R913 B.n396 B.n148 69.4205
R914 B.n403 B.n148 69.4205
R915 B.n403 B.n402 69.4205
R916 B.n409 B.n141 69.4205
R917 B.n415 B.n141 69.4205
R918 B.n415 B.n137 69.4205
R919 B.n421 B.n137 69.4205
R920 B.n421 B.n133 69.4205
R921 B.n427 B.n133 69.4205
R922 B.n427 B.n129 69.4205
R923 B.n433 B.n129 69.4205
R924 B.n433 B.n125 69.4205
R925 B.n440 B.n125 69.4205
R926 B.n440 B.n439 69.4205
R927 B.n446 B.n118 69.4205
R928 B.n453 B.n118 69.4205
R929 B.n453 B.n114 69.4205
R930 B.n459 B.n114 69.4205
R931 B.n459 B.n4 69.4205
R932 B.n714 B.n4 69.4205
R933 B.n714 B.n713 69.4205
R934 B.n713 B.n712 69.4205
R935 B.n712 B.n8 69.4205
R936 B.n12 B.n8 69.4205
R937 B.n705 B.n12 69.4205
R938 B.n705 B.n704 69.4205
R939 B.n704 B.n703 69.4205
R940 B.n697 B.n19 69.4205
R941 B.n697 B.n696 69.4205
R942 B.n696 B.n695 69.4205
R943 B.n695 B.n23 69.4205
R944 B.n689 B.n23 69.4205
R945 B.n689 B.n688 69.4205
R946 B.n688 B.n687 69.4205
R947 B.n687 B.n30 69.4205
R948 B.n681 B.n30 69.4205
R949 B.n681 B.n680 69.4205
R950 B.n680 B.n679 69.4205
R951 B.n673 B.n40 69.4205
R952 B.n673 B.n672 69.4205
R953 B.n672 B.n671 69.4205
R954 B.n671 B.n44 69.4205
R955 B.n665 B.n44 69.4205
R956 B.n665 B.n664 69.4205
R957 B.n664 B.n663 69.4205
R958 B.n663 B.n51 69.4205
R959 B.n657 B.n51 69.4205
R960 B.n657 B.n656 69.4205
R961 B.n656 B.n655 69.4205
R962 B.n655 B.n58 69.4205
R963 B.n649 B.n58 69.4205
R964 B.n649 B.n648 69.4205
R965 B.n647 B.n65 69.4205
R966 B.n641 B.n65 69.4205
R967 B.n641 B.n640 69.4205
R968 B.n640 B.n639 69.4205
R969 B.n639 B.n72 69.4205
R970 B.n633 B.n72 69.4205
R971 B.n633 B.n632 69.4205
R972 B.n632 B.n631 69.4205
R973 B.n360 B.t5 60.2325
R974 B.n446 B.t1 60.2325
R975 B.n703 B.t0 60.2325
R976 B.t12 B.n647 60.2325
R977 B.n95 B.n94 59.5399
R978 B.n564 B.n101 59.5399
R979 B.n270 B.n213 59.5399
R980 B.n288 B.n207 59.5399
R981 B.n402 B.t3 41.8566
R982 B.n40 B.t2 41.8566
R983 B.n334 B.n333 32.3127
R984 B.n338 B.n190 32.3127
R985 B.n518 B.n517 32.3127
R986 B.n629 B.n628 32.3127
R987 B.n409 B.t3 27.5643
R988 B.n679 B.t2 27.5643
R989 B B.n717 18.0485
R990 B.n334 B.n186 10.6151
R991 B.n344 B.n186 10.6151
R992 B.n345 B.n344 10.6151
R993 B.n346 B.n345 10.6151
R994 B.n346 B.n178 10.6151
R995 B.n356 B.n178 10.6151
R996 B.n357 B.n356 10.6151
R997 B.n358 B.n357 10.6151
R998 B.n358 B.n170 10.6151
R999 B.n368 B.n170 10.6151
R1000 B.n369 B.n368 10.6151
R1001 B.n370 B.n369 10.6151
R1002 B.n370 B.n162 10.6151
R1003 B.n380 B.n162 10.6151
R1004 B.n381 B.n380 10.6151
R1005 B.n382 B.n381 10.6151
R1006 B.n382 B.n154 10.6151
R1007 B.n392 B.n154 10.6151
R1008 B.n393 B.n392 10.6151
R1009 B.n394 B.n393 10.6151
R1010 B.n394 B.n146 10.6151
R1011 B.n405 B.n146 10.6151
R1012 B.n406 B.n405 10.6151
R1013 B.n407 B.n406 10.6151
R1014 B.n407 B.n139 10.6151
R1015 B.n417 B.n139 10.6151
R1016 B.n418 B.n417 10.6151
R1017 B.n419 B.n418 10.6151
R1018 B.n419 B.n131 10.6151
R1019 B.n429 B.n131 10.6151
R1020 B.n430 B.n429 10.6151
R1021 B.n431 B.n430 10.6151
R1022 B.n431 B.n123 10.6151
R1023 B.n442 B.n123 10.6151
R1024 B.n443 B.n442 10.6151
R1025 B.n444 B.n443 10.6151
R1026 B.n444 B.n116 10.6151
R1027 B.n455 B.n116 10.6151
R1028 B.n456 B.n455 10.6151
R1029 B.n457 B.n456 10.6151
R1030 B.n457 B.n0 10.6151
R1031 B.n333 B.n332 10.6151
R1032 B.n332 B.n194 10.6151
R1033 B.n327 B.n194 10.6151
R1034 B.n327 B.n326 10.6151
R1035 B.n326 B.n196 10.6151
R1036 B.n321 B.n196 10.6151
R1037 B.n321 B.n320 10.6151
R1038 B.n320 B.n319 10.6151
R1039 B.n319 B.n198 10.6151
R1040 B.n313 B.n198 10.6151
R1041 B.n313 B.n312 10.6151
R1042 B.n312 B.n311 10.6151
R1043 B.n311 B.n200 10.6151
R1044 B.n305 B.n200 10.6151
R1045 B.n305 B.n304 10.6151
R1046 B.n304 B.n303 10.6151
R1047 B.n303 B.n202 10.6151
R1048 B.n297 B.n202 10.6151
R1049 B.n297 B.n296 10.6151
R1050 B.n296 B.n295 10.6151
R1051 B.n295 B.n204 10.6151
R1052 B.n289 B.n204 10.6151
R1053 B.n287 B.n286 10.6151
R1054 B.n286 B.n208 10.6151
R1055 B.n280 B.n208 10.6151
R1056 B.n280 B.n279 10.6151
R1057 B.n279 B.n278 10.6151
R1058 B.n278 B.n210 10.6151
R1059 B.n272 B.n210 10.6151
R1060 B.n272 B.n271 10.6151
R1061 B.n269 B.n214 10.6151
R1062 B.n263 B.n214 10.6151
R1063 B.n263 B.n262 10.6151
R1064 B.n262 B.n261 10.6151
R1065 B.n261 B.n216 10.6151
R1066 B.n255 B.n216 10.6151
R1067 B.n255 B.n254 10.6151
R1068 B.n254 B.n253 10.6151
R1069 B.n253 B.n218 10.6151
R1070 B.n247 B.n218 10.6151
R1071 B.n247 B.n246 10.6151
R1072 B.n246 B.n245 10.6151
R1073 B.n245 B.n220 10.6151
R1074 B.n239 B.n220 10.6151
R1075 B.n239 B.n238 10.6151
R1076 B.n238 B.n237 10.6151
R1077 B.n237 B.n222 10.6151
R1078 B.n231 B.n222 10.6151
R1079 B.n231 B.n230 10.6151
R1080 B.n230 B.n229 10.6151
R1081 B.n229 B.n224 10.6151
R1082 B.n224 B.n190 10.6151
R1083 B.n339 B.n338 10.6151
R1084 B.n340 B.n339 10.6151
R1085 B.n340 B.n182 10.6151
R1086 B.n350 B.n182 10.6151
R1087 B.n351 B.n350 10.6151
R1088 B.n352 B.n351 10.6151
R1089 B.n352 B.n174 10.6151
R1090 B.n362 B.n174 10.6151
R1091 B.n363 B.n362 10.6151
R1092 B.n364 B.n363 10.6151
R1093 B.n364 B.n166 10.6151
R1094 B.n374 B.n166 10.6151
R1095 B.n375 B.n374 10.6151
R1096 B.n376 B.n375 10.6151
R1097 B.n376 B.n158 10.6151
R1098 B.n386 B.n158 10.6151
R1099 B.n387 B.n386 10.6151
R1100 B.n388 B.n387 10.6151
R1101 B.n388 B.n150 10.6151
R1102 B.n398 B.n150 10.6151
R1103 B.n399 B.n398 10.6151
R1104 B.n400 B.n399 10.6151
R1105 B.n400 B.n143 10.6151
R1106 B.n411 B.n143 10.6151
R1107 B.n412 B.n411 10.6151
R1108 B.n413 B.n412 10.6151
R1109 B.n413 B.n135 10.6151
R1110 B.n423 B.n135 10.6151
R1111 B.n424 B.n423 10.6151
R1112 B.n425 B.n424 10.6151
R1113 B.n425 B.n127 10.6151
R1114 B.n435 B.n127 10.6151
R1115 B.n436 B.n435 10.6151
R1116 B.n437 B.n436 10.6151
R1117 B.n437 B.n120 10.6151
R1118 B.n448 B.n120 10.6151
R1119 B.n449 B.n448 10.6151
R1120 B.n451 B.n449 10.6151
R1121 B.n451 B.n450 10.6151
R1122 B.n450 B.n112 10.6151
R1123 B.n462 B.n112 10.6151
R1124 B.n463 B.n462 10.6151
R1125 B.n464 B.n463 10.6151
R1126 B.n465 B.n464 10.6151
R1127 B.n466 B.n465 10.6151
R1128 B.n469 B.n466 10.6151
R1129 B.n470 B.n469 10.6151
R1130 B.n471 B.n470 10.6151
R1131 B.n472 B.n471 10.6151
R1132 B.n474 B.n472 10.6151
R1133 B.n475 B.n474 10.6151
R1134 B.n476 B.n475 10.6151
R1135 B.n477 B.n476 10.6151
R1136 B.n479 B.n477 10.6151
R1137 B.n480 B.n479 10.6151
R1138 B.n481 B.n480 10.6151
R1139 B.n482 B.n481 10.6151
R1140 B.n484 B.n482 10.6151
R1141 B.n485 B.n484 10.6151
R1142 B.n486 B.n485 10.6151
R1143 B.n487 B.n486 10.6151
R1144 B.n489 B.n487 10.6151
R1145 B.n490 B.n489 10.6151
R1146 B.n491 B.n490 10.6151
R1147 B.n492 B.n491 10.6151
R1148 B.n494 B.n492 10.6151
R1149 B.n495 B.n494 10.6151
R1150 B.n496 B.n495 10.6151
R1151 B.n497 B.n496 10.6151
R1152 B.n499 B.n497 10.6151
R1153 B.n500 B.n499 10.6151
R1154 B.n501 B.n500 10.6151
R1155 B.n502 B.n501 10.6151
R1156 B.n504 B.n502 10.6151
R1157 B.n505 B.n504 10.6151
R1158 B.n506 B.n505 10.6151
R1159 B.n507 B.n506 10.6151
R1160 B.n509 B.n507 10.6151
R1161 B.n510 B.n509 10.6151
R1162 B.n511 B.n510 10.6151
R1163 B.n512 B.n511 10.6151
R1164 B.n514 B.n512 10.6151
R1165 B.n515 B.n514 10.6151
R1166 B.n516 B.n515 10.6151
R1167 B.n517 B.n516 10.6151
R1168 B.n709 B.n1 10.6151
R1169 B.n709 B.n708 10.6151
R1170 B.n708 B.n707 10.6151
R1171 B.n707 B.n10 10.6151
R1172 B.n701 B.n10 10.6151
R1173 B.n701 B.n700 10.6151
R1174 B.n700 B.n699 10.6151
R1175 B.n699 B.n17 10.6151
R1176 B.n693 B.n17 10.6151
R1177 B.n693 B.n692 10.6151
R1178 B.n692 B.n691 10.6151
R1179 B.n691 B.n25 10.6151
R1180 B.n685 B.n25 10.6151
R1181 B.n685 B.n684 10.6151
R1182 B.n684 B.n683 10.6151
R1183 B.n683 B.n32 10.6151
R1184 B.n677 B.n32 10.6151
R1185 B.n677 B.n676 10.6151
R1186 B.n676 B.n675 10.6151
R1187 B.n675 B.n38 10.6151
R1188 B.n669 B.n38 10.6151
R1189 B.n669 B.n668 10.6151
R1190 B.n668 B.n667 10.6151
R1191 B.n667 B.n46 10.6151
R1192 B.n661 B.n46 10.6151
R1193 B.n661 B.n660 10.6151
R1194 B.n660 B.n659 10.6151
R1195 B.n659 B.n53 10.6151
R1196 B.n653 B.n53 10.6151
R1197 B.n653 B.n652 10.6151
R1198 B.n652 B.n651 10.6151
R1199 B.n651 B.n60 10.6151
R1200 B.n645 B.n60 10.6151
R1201 B.n645 B.n644 10.6151
R1202 B.n644 B.n643 10.6151
R1203 B.n643 B.n67 10.6151
R1204 B.n637 B.n67 10.6151
R1205 B.n637 B.n636 10.6151
R1206 B.n636 B.n635 10.6151
R1207 B.n635 B.n74 10.6151
R1208 B.n629 B.n74 10.6151
R1209 B.n628 B.n627 10.6151
R1210 B.n627 B.n81 10.6151
R1211 B.n621 B.n81 10.6151
R1212 B.n621 B.n620 10.6151
R1213 B.n620 B.n619 10.6151
R1214 B.n619 B.n83 10.6151
R1215 B.n613 B.n83 10.6151
R1216 B.n613 B.n612 10.6151
R1217 B.n612 B.n611 10.6151
R1218 B.n611 B.n85 10.6151
R1219 B.n605 B.n85 10.6151
R1220 B.n605 B.n604 10.6151
R1221 B.n604 B.n603 10.6151
R1222 B.n603 B.n87 10.6151
R1223 B.n597 B.n87 10.6151
R1224 B.n597 B.n596 10.6151
R1225 B.n596 B.n595 10.6151
R1226 B.n595 B.n89 10.6151
R1227 B.n589 B.n89 10.6151
R1228 B.n589 B.n588 10.6151
R1229 B.n588 B.n587 10.6151
R1230 B.n587 B.n91 10.6151
R1231 B.n581 B.n580 10.6151
R1232 B.n580 B.n579 10.6151
R1233 B.n579 B.n96 10.6151
R1234 B.n573 B.n96 10.6151
R1235 B.n573 B.n572 10.6151
R1236 B.n572 B.n571 10.6151
R1237 B.n571 B.n98 10.6151
R1238 B.n565 B.n98 10.6151
R1239 B.n563 B.n562 10.6151
R1240 B.n562 B.n102 10.6151
R1241 B.n556 B.n102 10.6151
R1242 B.n556 B.n555 10.6151
R1243 B.n555 B.n554 10.6151
R1244 B.n554 B.n104 10.6151
R1245 B.n548 B.n104 10.6151
R1246 B.n548 B.n547 10.6151
R1247 B.n547 B.n546 10.6151
R1248 B.n546 B.n106 10.6151
R1249 B.n540 B.n106 10.6151
R1250 B.n540 B.n539 10.6151
R1251 B.n539 B.n538 10.6151
R1252 B.n538 B.n108 10.6151
R1253 B.n532 B.n108 10.6151
R1254 B.n532 B.n531 10.6151
R1255 B.n531 B.n530 10.6151
R1256 B.n530 B.n110 10.6151
R1257 B.n524 B.n110 10.6151
R1258 B.n524 B.n523 10.6151
R1259 B.n523 B.n522 10.6151
R1260 B.n522 B.n518 10.6151
R1261 B.t5 B.n172 9.18843
R1262 B.n439 B.t1 9.18843
R1263 B.n19 B.t0 9.18843
R1264 B.n648 B.t12 9.18843
R1265 B.n717 B.n0 8.11757
R1266 B.n717 B.n1 8.11757
R1267 B.n288 B.n287 6.5566
R1268 B.n271 B.n270 6.5566
R1269 B.n581 B.n95 6.5566
R1270 B.n565 B.n564 6.5566
R1271 B.n289 B.n288 4.05904
R1272 B.n270 B.n269 4.05904
R1273 B.n95 B.n91 4.05904
R1274 B.n564 B.n563 4.05904
R1275 VP.n19 VP.n18 161.3
R1276 VP.n17 VP.n1 161.3
R1277 VP.n16 VP.n15 161.3
R1278 VP.n14 VP.n2 161.3
R1279 VP.n13 VP.n12 161.3
R1280 VP.n11 VP.n3 161.3
R1281 VP.n10 VP.n9 161.3
R1282 VP.n8 VP.n4 161.3
R1283 VP.n7 VP.n6 79.917
R1284 VP.n20 VP.n0 79.917
R1285 VP.n5 VP.t2 71.8343
R1286 VP.n5 VP.t0 70.5919
R1287 VP.n12 VP.n2 56.5617
R1288 VP.n7 VP.n5 46.6141
R1289 VP.n6 VP.t1 36.9225
R1290 VP.n0 VP.t3 36.9225
R1291 VP.n10 VP.n4 24.5923
R1292 VP.n11 VP.n10 24.5923
R1293 VP.n12 VP.n11 24.5923
R1294 VP.n16 VP.n2 24.5923
R1295 VP.n17 VP.n16 24.5923
R1296 VP.n18 VP.n17 24.5923
R1297 VP.n6 VP.n4 10.3291
R1298 VP.n18 VP.n0 10.3291
R1299 VP.n8 VP.n7 0.354861
R1300 VP.n20 VP.n19 0.354861
R1301 VP VP.n20 0.267071
R1302 VP.n9 VP.n8 0.189894
R1303 VP.n9 VP.n3 0.189894
R1304 VP.n13 VP.n3 0.189894
R1305 VP.n14 VP.n13 0.189894
R1306 VP.n15 VP.n14 0.189894
R1307 VP.n15 VP.n1 0.189894
R1308 VP.n19 VP.n1 0.189894
R1309 VDD1 VDD1.n1 110.353
R1310 VDD1 VDD1.n0 71.2907
R1311 VDD1.n0 VDD1.t1 3.6005
R1312 VDD1.n0 VDD1.t3 3.6005
R1313 VDD1.n1 VDD1.t2 3.6005
R1314 VDD1.n1 VDD1.t0 3.6005
C0 VN VDD1 0.15038f
C1 VN VDD2 2.46724f
C2 VTAIL VDD1 4.29406f
C3 VTAIL VDD2 4.3549f
C4 VDD1 VDD2 1.26503f
C5 VP VN 5.694991f
C6 VTAIL VP 3.00448f
C7 VTAIL VN 2.99037f
C8 VP VDD1 2.77365f
C9 VP VDD2 0.457786f
C10 VDD2 B 3.840405f
C11 VDD1 B 7.80785f
C12 VTAIL B 6.350605f
C13 VN B 12.07905f
C14 VP B 10.437232f
C15 VDD1.t1 B 0.12671f
C16 VDD1.t3 B 0.12671f
C17 VDD1.n0 B 1.05831f
C18 VDD1.t2 B 0.12671f
C19 VDD1.t0 B 0.12671f
C20 VDD1.n1 B 1.57525f
C21 VP.t3 B 1.31831f
C22 VP.n0 B 0.590932f
C23 VP.n1 B 0.025361f
C24 VP.n2 B 0.036867f
C25 VP.n3 B 0.025361f
C26 VP.n4 B 0.033564f
C27 VP.t2 B 1.65439f
C28 VP.t0 B 1.6428f
C29 VP.n5 B 2.38261f
C30 VP.t1 B 1.31831f
C31 VP.n6 B 0.590932f
C32 VP.n7 B 1.31511f
C33 VP.n8 B 0.040926f
C34 VP.n9 B 0.025361f
C35 VP.n10 B 0.04703f
C36 VP.n11 B 0.04703f
C37 VP.n12 B 0.036867f
C38 VP.n13 B 0.025361f
C39 VP.n14 B 0.025361f
C40 VP.n15 B 0.025361f
C41 VP.n16 B 0.04703f
C42 VP.n17 B 0.04703f
C43 VP.n18 B 0.033564f
C44 VP.n19 B 0.040926f
C45 VP.n20 B 0.068858f
C46 VDD2.t0 B 0.125037f
C47 VDD2.t3 B 0.125037f
C48 VDD2.n0 B 1.52983f
C49 VDD2.t2 B 0.125037f
C50 VDD2.t1 B 0.125037f
C51 VDD2.n1 B 1.04389f
C52 VDD2.n2 B 3.50667f
C53 VTAIL.t7 B 0.926043f
C54 VTAIL.n0 B 0.390135f
C55 VTAIL.t1 B 0.926043f
C56 VTAIL.n1 B 0.502568f
C57 VTAIL.t3 B 0.926043f
C58 VTAIL.n2 B 1.32035f
C59 VTAIL.t4 B 0.926043f
C60 VTAIL.n3 B 1.32035f
C61 VTAIL.t5 B 0.926043f
C62 VTAIL.n4 B 0.502567f
C63 VTAIL.t0 B 0.926043f
C64 VTAIL.n5 B 0.502567f
C65 VTAIL.t2 B 0.926039f
C66 VTAIL.n6 B 1.32035f
C67 VTAIL.t6 B 0.926043f
C68 VTAIL.n7 B 1.1999f
C69 VN.t0 B 1.595f
C70 VN.t3 B 1.60626f
C71 VN.n0 B 0.935597f
C72 VN.t2 B 1.60626f
C73 VN.t1 B 1.595f
C74 VN.n1 B 2.32355f
.ends

