* NGSPICE file created from diff_pair_sample_1071.ext - technology: sky130A

.subckt diff_pair_sample_1071 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VN.t0 VDD2.t6 w_n4770_n1148# sky130_fd_pr__pfet_01v8 ad=0.1485 pd=1.23 as=0.1485 ps=1.23 w=0.9 l=3.47
X1 VTAIL.t4 VP.t0 VDD1.t7 w_n4770_n1148# sky130_fd_pr__pfet_01v8 ad=0.351 pd=2.58 as=0.1485 ps=1.23 w=0.9 l=3.47
X2 VTAIL.t6 VP.t1 VDD1.t6 w_n4770_n1148# sky130_fd_pr__pfet_01v8 ad=0.1485 pd=1.23 as=0.1485 ps=1.23 w=0.9 l=3.47
X3 VDD1.t5 VP.t2 VTAIL.t5 w_n4770_n1148# sky130_fd_pr__pfet_01v8 ad=0.1485 pd=1.23 as=0.351 ps=2.58 w=0.9 l=3.47
X4 VDD2.t7 VN.t1 VTAIL.t14 w_n4770_n1148# sky130_fd_pr__pfet_01v8 ad=0.1485 pd=1.23 as=0.1485 ps=1.23 w=0.9 l=3.47
X5 VTAIL.t0 VP.t3 VDD1.t4 w_n4770_n1148# sky130_fd_pr__pfet_01v8 ad=0.351 pd=2.58 as=0.1485 ps=1.23 w=0.9 l=3.47
X6 B.t11 B.t9 B.t10 w_n4770_n1148# sky130_fd_pr__pfet_01v8 ad=0.351 pd=2.58 as=0 ps=0 w=0.9 l=3.47
X7 VDD2.t3 VN.t2 VTAIL.t13 w_n4770_n1148# sky130_fd_pr__pfet_01v8 ad=0.1485 pd=1.23 as=0.351 ps=2.58 w=0.9 l=3.47
X8 VDD2.t1 VN.t3 VTAIL.t12 w_n4770_n1148# sky130_fd_pr__pfet_01v8 ad=0.1485 pd=1.23 as=0.351 ps=2.58 w=0.9 l=3.47
X9 VDD1.t3 VP.t4 VTAIL.t2 w_n4770_n1148# sky130_fd_pr__pfet_01v8 ad=0.1485 pd=1.23 as=0.1485 ps=1.23 w=0.9 l=3.47
X10 VDD2.t2 VN.t4 VTAIL.t11 w_n4770_n1148# sky130_fd_pr__pfet_01v8 ad=0.1485 pd=1.23 as=0.1485 ps=1.23 w=0.9 l=3.47
X11 VDD1.t2 VP.t5 VTAIL.t3 w_n4770_n1148# sky130_fd_pr__pfet_01v8 ad=0.1485 pd=1.23 as=0.1485 ps=1.23 w=0.9 l=3.47
X12 B.t8 B.t6 B.t7 w_n4770_n1148# sky130_fd_pr__pfet_01v8 ad=0.351 pd=2.58 as=0 ps=0 w=0.9 l=3.47
X13 VTAIL.t10 VN.t5 VDD2.t4 w_n4770_n1148# sky130_fd_pr__pfet_01v8 ad=0.351 pd=2.58 as=0.1485 ps=1.23 w=0.9 l=3.47
X14 B.t5 B.t3 B.t4 w_n4770_n1148# sky130_fd_pr__pfet_01v8 ad=0.351 pd=2.58 as=0 ps=0 w=0.9 l=3.47
X15 VTAIL.t7 VP.t6 VDD1.t1 w_n4770_n1148# sky130_fd_pr__pfet_01v8 ad=0.1485 pd=1.23 as=0.1485 ps=1.23 w=0.9 l=3.47
X16 VTAIL.t9 VN.t6 VDD2.t5 w_n4770_n1148# sky130_fd_pr__pfet_01v8 ad=0.1485 pd=1.23 as=0.1485 ps=1.23 w=0.9 l=3.47
X17 B.t2 B.t0 B.t1 w_n4770_n1148# sky130_fd_pr__pfet_01v8 ad=0.351 pd=2.58 as=0 ps=0 w=0.9 l=3.47
X18 VTAIL.t8 VN.t7 VDD2.t0 w_n4770_n1148# sky130_fd_pr__pfet_01v8 ad=0.351 pd=2.58 as=0.1485 ps=1.23 w=0.9 l=3.47
X19 VDD1.t0 VP.t7 VTAIL.t1 w_n4770_n1148# sky130_fd_pr__pfet_01v8 ad=0.1485 pd=1.23 as=0.351 ps=2.58 w=0.9 l=3.47
R0 VN.n68 VN.n67 161.3
R1 VN.n66 VN.n36 161.3
R2 VN.n65 VN.n64 161.3
R3 VN.n63 VN.n37 161.3
R4 VN.n62 VN.n61 161.3
R5 VN.n60 VN.n38 161.3
R6 VN.n59 VN.n58 161.3
R7 VN.n57 VN.n39 161.3
R8 VN.n56 VN.n55 161.3
R9 VN.n54 VN.n40 161.3
R10 VN.n53 VN.n52 161.3
R11 VN.n51 VN.n42 161.3
R12 VN.n50 VN.n49 161.3
R13 VN.n48 VN.n43 161.3
R14 VN.n47 VN.n46 161.3
R15 VN.n33 VN.n32 161.3
R16 VN.n31 VN.n1 161.3
R17 VN.n30 VN.n29 161.3
R18 VN.n28 VN.n2 161.3
R19 VN.n27 VN.n26 161.3
R20 VN.n25 VN.n3 161.3
R21 VN.n24 VN.n23 161.3
R22 VN.n22 VN.n4 161.3
R23 VN.n21 VN.n20 161.3
R24 VN.n18 VN.n5 161.3
R25 VN.n17 VN.n16 161.3
R26 VN.n15 VN.n6 161.3
R27 VN.n14 VN.n13 161.3
R28 VN.n12 VN.n7 161.3
R29 VN.n11 VN.n10 161.3
R30 VN.n34 VN.n0 80.4088
R31 VN.n69 VN.n35 80.4088
R32 VN.n26 VN.n2 56.5617
R33 VN.n61 VN.n37 56.5617
R34 VN.n9 VN.n8 55.1568
R35 VN.n45 VN.n44 55.1568
R36 VN VN.n69 46.8012
R37 VN.n13 VN.n6 40.577
R38 VN.n17 VN.n6 40.577
R39 VN.n49 VN.n42 40.577
R40 VN.n53 VN.n42 40.577
R41 VN.n45 VN.t2 39.696
R42 VN.n9 VN.t5 39.696
R43 VN.n12 VN.n11 24.5923
R44 VN.n13 VN.n12 24.5923
R45 VN.n18 VN.n17 24.5923
R46 VN.n20 VN.n18 24.5923
R47 VN.n24 VN.n4 24.5923
R48 VN.n25 VN.n24 24.5923
R49 VN.n26 VN.n25 24.5923
R50 VN.n30 VN.n2 24.5923
R51 VN.n31 VN.n30 24.5923
R52 VN.n32 VN.n31 24.5923
R53 VN.n49 VN.n48 24.5923
R54 VN.n48 VN.n47 24.5923
R55 VN.n61 VN.n60 24.5923
R56 VN.n60 VN.n59 24.5923
R57 VN.n59 VN.n39 24.5923
R58 VN.n55 VN.n54 24.5923
R59 VN.n54 VN.n53 24.5923
R60 VN.n67 VN.n66 24.5923
R61 VN.n66 VN.n65 24.5923
R62 VN.n65 VN.n37 24.5923
R63 VN.n11 VN.n8 19.674
R64 VN.n20 VN.n19 19.674
R65 VN.n47 VN.n44 19.674
R66 VN.n55 VN.n41 19.674
R67 VN.n32 VN.n0 9.83723
R68 VN.n67 VN.n35 9.83723
R69 VN.n8 VN.t1 6.25122
R70 VN.n19 VN.t6 6.25122
R71 VN.n0 VN.t3 6.25122
R72 VN.n44 VN.t0 6.25122
R73 VN.n41 VN.t4 6.25122
R74 VN.n35 VN.t7 6.25122
R75 VN.n19 VN.n4 4.91887
R76 VN.n41 VN.n39 4.91887
R77 VN.n46 VN.n45 3.15112
R78 VN.n10 VN.n9 3.15112
R79 VN.n69 VN.n68 0.354861
R80 VN.n34 VN.n33 0.354861
R81 VN VN.n34 0.267071
R82 VN.n68 VN.n36 0.189894
R83 VN.n64 VN.n36 0.189894
R84 VN.n64 VN.n63 0.189894
R85 VN.n63 VN.n62 0.189894
R86 VN.n62 VN.n38 0.189894
R87 VN.n58 VN.n38 0.189894
R88 VN.n58 VN.n57 0.189894
R89 VN.n57 VN.n56 0.189894
R90 VN.n56 VN.n40 0.189894
R91 VN.n52 VN.n40 0.189894
R92 VN.n52 VN.n51 0.189894
R93 VN.n51 VN.n50 0.189894
R94 VN.n50 VN.n43 0.189894
R95 VN.n46 VN.n43 0.189894
R96 VN.n10 VN.n7 0.189894
R97 VN.n14 VN.n7 0.189894
R98 VN.n15 VN.n14 0.189894
R99 VN.n16 VN.n15 0.189894
R100 VN.n16 VN.n5 0.189894
R101 VN.n21 VN.n5 0.189894
R102 VN.n22 VN.n21 0.189894
R103 VN.n23 VN.n22 0.189894
R104 VN.n23 VN.n3 0.189894
R105 VN.n27 VN.n3 0.189894
R106 VN.n28 VN.n27 0.189894
R107 VN.n29 VN.n28 0.189894
R108 VN.n29 VN.n1 0.189894
R109 VN.n33 VN.n1 0.189894
R110 VDD2.n2 VDD2.n1 639.775
R111 VDD2.n2 VDD2.n0 639.775
R112 VDD2 VDD2.n5 639.774
R113 VDD2.n4 VDD2.n3 638.193
R114 VDD2.n4 VDD2.n2 39.2325
R115 VDD2.n5 VDD2.t6 36.1172
R116 VDD2.n5 VDD2.t3 36.1172
R117 VDD2.n3 VDD2.t0 36.1172
R118 VDD2.n3 VDD2.t2 36.1172
R119 VDD2.n1 VDD2.t5 36.1172
R120 VDD2.n1 VDD2.t1 36.1172
R121 VDD2.n0 VDD2.t4 36.1172
R122 VDD2.n0 VDD2.t7 36.1172
R123 VDD2 VDD2.n4 1.69662
R124 VTAIL.n14 VTAIL.t5 657.631
R125 VTAIL.n11 VTAIL.t4 657.631
R126 VTAIL.n10 VTAIL.t13 657.631
R127 VTAIL.n7 VTAIL.t8 657.631
R128 VTAIL.n15 VTAIL.t12 657.63
R129 VTAIL.n2 VTAIL.t10 657.63
R130 VTAIL.n3 VTAIL.t1 657.63
R131 VTAIL.n6 VTAIL.t0 657.63
R132 VTAIL.n13 VTAIL.n12 621.514
R133 VTAIL.n9 VTAIL.n8 621.514
R134 VTAIL.n1 VTAIL.n0 621.514
R135 VTAIL.n5 VTAIL.n4 621.514
R136 VTAIL.n0 VTAIL.t14 36.1172
R137 VTAIL.n0 VTAIL.t9 36.1172
R138 VTAIL.n4 VTAIL.t3 36.1172
R139 VTAIL.n4 VTAIL.t6 36.1172
R140 VTAIL.n12 VTAIL.t2 36.1172
R141 VTAIL.n12 VTAIL.t7 36.1172
R142 VTAIL.n8 VTAIL.t11 36.1172
R143 VTAIL.n8 VTAIL.t15 36.1172
R144 VTAIL.n15 VTAIL.n14 16.4186
R145 VTAIL.n7 VTAIL.n6 16.4186
R146 VTAIL.n9 VTAIL.n7 3.27636
R147 VTAIL.n10 VTAIL.n9 3.27636
R148 VTAIL.n13 VTAIL.n11 3.27636
R149 VTAIL.n14 VTAIL.n13 3.27636
R150 VTAIL.n6 VTAIL.n5 3.27636
R151 VTAIL.n5 VTAIL.n3 3.27636
R152 VTAIL.n2 VTAIL.n1 3.27636
R153 VTAIL VTAIL.n15 3.21817
R154 VTAIL.n11 VTAIL.n10 0.470328
R155 VTAIL.n3 VTAIL.n2 0.470328
R156 VTAIL VTAIL.n1 0.0586897
R157 VP.n24 VP.n23 161.3
R158 VP.n25 VP.n20 161.3
R159 VP.n27 VP.n26 161.3
R160 VP.n28 VP.n19 161.3
R161 VP.n30 VP.n29 161.3
R162 VP.n31 VP.n18 161.3
R163 VP.n34 VP.n33 161.3
R164 VP.n35 VP.n17 161.3
R165 VP.n37 VP.n36 161.3
R166 VP.n38 VP.n16 161.3
R167 VP.n40 VP.n39 161.3
R168 VP.n41 VP.n15 161.3
R169 VP.n43 VP.n42 161.3
R170 VP.n44 VP.n14 161.3
R171 VP.n46 VP.n45 161.3
R172 VP.n85 VP.n84 161.3
R173 VP.n83 VP.n1 161.3
R174 VP.n82 VP.n81 161.3
R175 VP.n80 VP.n2 161.3
R176 VP.n79 VP.n78 161.3
R177 VP.n77 VP.n3 161.3
R178 VP.n76 VP.n75 161.3
R179 VP.n74 VP.n4 161.3
R180 VP.n73 VP.n72 161.3
R181 VP.n70 VP.n5 161.3
R182 VP.n69 VP.n68 161.3
R183 VP.n67 VP.n6 161.3
R184 VP.n66 VP.n65 161.3
R185 VP.n64 VP.n7 161.3
R186 VP.n63 VP.n62 161.3
R187 VP.n61 VP.n60 161.3
R188 VP.n59 VP.n9 161.3
R189 VP.n58 VP.n57 161.3
R190 VP.n56 VP.n10 161.3
R191 VP.n55 VP.n54 161.3
R192 VP.n53 VP.n11 161.3
R193 VP.n52 VP.n51 161.3
R194 VP.n50 VP.n12 161.3
R195 VP.n49 VP.n48 80.4088
R196 VP.n86 VP.n0 80.4088
R197 VP.n47 VP.n13 80.4088
R198 VP.n54 VP.n10 56.5617
R199 VP.n78 VP.n2 56.5617
R200 VP.n39 VP.n15 56.5617
R201 VP.n22 VP.n21 55.1568
R202 VP.n49 VP.n47 46.6359
R203 VP.n65 VP.n6 40.577
R204 VP.n69 VP.n6 40.577
R205 VP.n30 VP.n19 40.577
R206 VP.n26 VP.n19 40.577
R207 VP.n22 VP.t0 39.6958
R208 VP.n52 VP.n12 24.5923
R209 VP.n53 VP.n52 24.5923
R210 VP.n54 VP.n53 24.5923
R211 VP.n58 VP.n10 24.5923
R212 VP.n59 VP.n58 24.5923
R213 VP.n60 VP.n59 24.5923
R214 VP.n64 VP.n63 24.5923
R215 VP.n65 VP.n64 24.5923
R216 VP.n70 VP.n69 24.5923
R217 VP.n72 VP.n70 24.5923
R218 VP.n76 VP.n4 24.5923
R219 VP.n77 VP.n76 24.5923
R220 VP.n78 VP.n77 24.5923
R221 VP.n82 VP.n2 24.5923
R222 VP.n83 VP.n82 24.5923
R223 VP.n84 VP.n83 24.5923
R224 VP.n43 VP.n15 24.5923
R225 VP.n44 VP.n43 24.5923
R226 VP.n45 VP.n44 24.5923
R227 VP.n31 VP.n30 24.5923
R228 VP.n33 VP.n31 24.5923
R229 VP.n37 VP.n17 24.5923
R230 VP.n38 VP.n37 24.5923
R231 VP.n39 VP.n38 24.5923
R232 VP.n25 VP.n24 24.5923
R233 VP.n26 VP.n25 24.5923
R234 VP.n63 VP.n8 19.674
R235 VP.n72 VP.n71 19.674
R236 VP.n33 VP.n32 19.674
R237 VP.n24 VP.n21 19.674
R238 VP.n48 VP.n12 9.83723
R239 VP.n84 VP.n0 9.83723
R240 VP.n45 VP.n13 9.83723
R241 VP.n48 VP.t3 6.25122
R242 VP.n8 VP.t5 6.25122
R243 VP.n71 VP.t1 6.25122
R244 VP.n0 VP.t7 6.25122
R245 VP.n13 VP.t2 6.25122
R246 VP.n32 VP.t6 6.25122
R247 VP.n21 VP.t4 6.25122
R248 VP.n60 VP.n8 4.91887
R249 VP.n71 VP.n4 4.91887
R250 VP.n32 VP.n17 4.91887
R251 VP.n23 VP.n22 3.1511
R252 VP.n47 VP.n46 0.354861
R253 VP.n50 VP.n49 0.354861
R254 VP.n86 VP.n85 0.354861
R255 VP VP.n86 0.267071
R256 VP.n23 VP.n20 0.189894
R257 VP.n27 VP.n20 0.189894
R258 VP.n28 VP.n27 0.189894
R259 VP.n29 VP.n28 0.189894
R260 VP.n29 VP.n18 0.189894
R261 VP.n34 VP.n18 0.189894
R262 VP.n35 VP.n34 0.189894
R263 VP.n36 VP.n35 0.189894
R264 VP.n36 VP.n16 0.189894
R265 VP.n40 VP.n16 0.189894
R266 VP.n41 VP.n40 0.189894
R267 VP.n42 VP.n41 0.189894
R268 VP.n42 VP.n14 0.189894
R269 VP.n46 VP.n14 0.189894
R270 VP.n51 VP.n50 0.189894
R271 VP.n51 VP.n11 0.189894
R272 VP.n55 VP.n11 0.189894
R273 VP.n56 VP.n55 0.189894
R274 VP.n57 VP.n56 0.189894
R275 VP.n57 VP.n9 0.189894
R276 VP.n61 VP.n9 0.189894
R277 VP.n62 VP.n61 0.189894
R278 VP.n62 VP.n7 0.189894
R279 VP.n66 VP.n7 0.189894
R280 VP.n67 VP.n66 0.189894
R281 VP.n68 VP.n67 0.189894
R282 VP.n68 VP.n5 0.189894
R283 VP.n73 VP.n5 0.189894
R284 VP.n74 VP.n73 0.189894
R285 VP.n75 VP.n74 0.189894
R286 VP.n75 VP.n3 0.189894
R287 VP.n79 VP.n3 0.189894
R288 VP.n80 VP.n79 0.189894
R289 VP.n81 VP.n80 0.189894
R290 VP.n81 VP.n1 0.189894
R291 VP.n85 VP.n1 0.189894
R292 VDD1 VDD1.n0 639.889
R293 VDD1.n3 VDD1.n2 639.775
R294 VDD1.n3 VDD1.n1 639.775
R295 VDD1.n5 VDD1.n4 638.193
R296 VDD1.n5 VDD1.n3 39.8155
R297 VDD1.n4 VDD1.t1 36.1172
R298 VDD1.n4 VDD1.t5 36.1172
R299 VDD1.n0 VDD1.t7 36.1172
R300 VDD1.n0 VDD1.t3 36.1172
R301 VDD1.n2 VDD1.t6 36.1172
R302 VDD1.n2 VDD1.t0 36.1172
R303 VDD1.n1 VDD1.t4 36.1172
R304 VDD1.n1 VDD1.t2 36.1172
R305 VDD1 VDD1.n5 1.58024
R306 B.n285 B.t11 721.966
R307 B.n127 B.t5 721.966
R308 B.n40 B.t1 721.966
R309 B.n47 B.t7 721.966
R310 B.n286 B.t10 648.269
R311 B.n128 B.t4 648.269
R312 B.n41 B.t2 648.269
R313 B.n48 B.t8 648.269
R314 B.n497 B.n52 585
R315 B.n499 B.n498 585
R316 B.n500 B.n51 585
R317 B.n502 B.n501 585
R318 B.n503 B.n50 585
R319 B.n505 B.n504 585
R320 B.n506 B.n49 585
R321 B.n508 B.n507 585
R322 B.n509 B.n46 585
R323 B.n512 B.n511 585
R324 B.n513 B.n45 585
R325 B.n515 B.n514 585
R326 B.n516 B.n44 585
R327 B.n518 B.n517 585
R328 B.n519 B.n43 585
R329 B.n521 B.n520 585
R330 B.n522 B.n39 585
R331 B.n524 B.n523 585
R332 B.n525 B.n38 585
R333 B.n527 B.n526 585
R334 B.n528 B.n37 585
R335 B.n530 B.n529 585
R336 B.n531 B.n36 585
R337 B.n533 B.n532 585
R338 B.n534 B.n35 585
R339 B.n536 B.n535 585
R340 B.n537 B.n34 585
R341 B.n496 B.n495 585
R342 B.n494 B.n53 585
R343 B.n493 B.n492 585
R344 B.n491 B.n54 585
R345 B.n490 B.n489 585
R346 B.n488 B.n55 585
R347 B.n487 B.n486 585
R348 B.n485 B.n56 585
R349 B.n484 B.n483 585
R350 B.n482 B.n57 585
R351 B.n481 B.n480 585
R352 B.n479 B.n58 585
R353 B.n478 B.n477 585
R354 B.n476 B.n59 585
R355 B.n475 B.n474 585
R356 B.n473 B.n60 585
R357 B.n472 B.n471 585
R358 B.n470 B.n61 585
R359 B.n469 B.n468 585
R360 B.n467 B.n62 585
R361 B.n466 B.n465 585
R362 B.n464 B.n63 585
R363 B.n463 B.n462 585
R364 B.n461 B.n64 585
R365 B.n460 B.n459 585
R366 B.n458 B.n65 585
R367 B.n457 B.n456 585
R368 B.n455 B.n66 585
R369 B.n454 B.n453 585
R370 B.n452 B.n67 585
R371 B.n451 B.n450 585
R372 B.n449 B.n68 585
R373 B.n448 B.n447 585
R374 B.n446 B.n69 585
R375 B.n445 B.n444 585
R376 B.n443 B.n70 585
R377 B.n442 B.n441 585
R378 B.n440 B.n71 585
R379 B.n439 B.n438 585
R380 B.n437 B.n72 585
R381 B.n436 B.n435 585
R382 B.n434 B.n73 585
R383 B.n433 B.n432 585
R384 B.n431 B.n74 585
R385 B.n430 B.n429 585
R386 B.n428 B.n75 585
R387 B.n427 B.n426 585
R388 B.n425 B.n76 585
R389 B.n424 B.n423 585
R390 B.n422 B.n77 585
R391 B.n421 B.n420 585
R392 B.n419 B.n78 585
R393 B.n418 B.n417 585
R394 B.n416 B.n79 585
R395 B.n415 B.n414 585
R396 B.n413 B.n80 585
R397 B.n412 B.n411 585
R398 B.n410 B.n81 585
R399 B.n409 B.n408 585
R400 B.n407 B.n82 585
R401 B.n406 B.n405 585
R402 B.n404 B.n83 585
R403 B.n403 B.n402 585
R404 B.n401 B.n84 585
R405 B.n400 B.n399 585
R406 B.n398 B.n85 585
R407 B.n397 B.n396 585
R408 B.n395 B.n86 585
R409 B.n394 B.n393 585
R410 B.n392 B.n87 585
R411 B.n391 B.n390 585
R412 B.n389 B.n88 585
R413 B.n388 B.n387 585
R414 B.n386 B.n89 585
R415 B.n385 B.n384 585
R416 B.n383 B.n90 585
R417 B.n382 B.n381 585
R418 B.n380 B.n91 585
R419 B.n379 B.n378 585
R420 B.n377 B.n92 585
R421 B.n376 B.n375 585
R422 B.n374 B.n93 585
R423 B.n373 B.n372 585
R424 B.n371 B.n94 585
R425 B.n370 B.n369 585
R426 B.n368 B.n95 585
R427 B.n367 B.n366 585
R428 B.n365 B.n96 585
R429 B.n364 B.n363 585
R430 B.n362 B.n97 585
R431 B.n361 B.n360 585
R432 B.n359 B.n98 585
R433 B.n358 B.n357 585
R434 B.n356 B.n99 585
R435 B.n355 B.n354 585
R436 B.n353 B.n100 585
R437 B.n352 B.n351 585
R438 B.n350 B.n101 585
R439 B.n349 B.n348 585
R440 B.n347 B.n102 585
R441 B.n346 B.n345 585
R442 B.n344 B.n103 585
R443 B.n343 B.n342 585
R444 B.n341 B.n104 585
R445 B.n340 B.n339 585
R446 B.n338 B.n105 585
R447 B.n337 B.n336 585
R448 B.n335 B.n106 585
R449 B.n334 B.n333 585
R450 B.n332 B.n107 585
R451 B.n331 B.n330 585
R452 B.n329 B.n108 585
R453 B.n328 B.n327 585
R454 B.n326 B.n109 585
R455 B.n325 B.n324 585
R456 B.n323 B.n110 585
R457 B.n322 B.n321 585
R458 B.n320 B.n111 585
R459 B.n319 B.n318 585
R460 B.n317 B.n112 585
R461 B.n316 B.n315 585
R462 B.n314 B.n113 585
R463 B.n313 B.n312 585
R464 B.n311 B.n114 585
R465 B.n310 B.n309 585
R466 B.n308 B.n115 585
R467 B.n307 B.n306 585
R468 B.n305 B.n116 585
R469 B.n304 B.n303 585
R470 B.n259 B.n132 585
R471 B.n261 B.n260 585
R472 B.n262 B.n131 585
R473 B.n264 B.n263 585
R474 B.n265 B.n130 585
R475 B.n267 B.n266 585
R476 B.n268 B.n129 585
R477 B.n270 B.n269 585
R478 B.n271 B.n126 585
R479 B.n274 B.n273 585
R480 B.n275 B.n125 585
R481 B.n277 B.n276 585
R482 B.n278 B.n124 585
R483 B.n280 B.n279 585
R484 B.n281 B.n123 585
R485 B.n283 B.n282 585
R486 B.n284 B.n122 585
R487 B.n289 B.n288 585
R488 B.n290 B.n121 585
R489 B.n292 B.n291 585
R490 B.n293 B.n120 585
R491 B.n295 B.n294 585
R492 B.n296 B.n119 585
R493 B.n298 B.n297 585
R494 B.n299 B.n118 585
R495 B.n301 B.n300 585
R496 B.n302 B.n117 585
R497 B.n258 B.n257 585
R498 B.n256 B.n133 585
R499 B.n255 B.n254 585
R500 B.n253 B.n134 585
R501 B.n252 B.n251 585
R502 B.n250 B.n135 585
R503 B.n249 B.n248 585
R504 B.n247 B.n136 585
R505 B.n246 B.n245 585
R506 B.n244 B.n137 585
R507 B.n243 B.n242 585
R508 B.n241 B.n138 585
R509 B.n240 B.n239 585
R510 B.n238 B.n139 585
R511 B.n237 B.n236 585
R512 B.n235 B.n140 585
R513 B.n234 B.n233 585
R514 B.n232 B.n141 585
R515 B.n231 B.n230 585
R516 B.n229 B.n142 585
R517 B.n228 B.n227 585
R518 B.n226 B.n143 585
R519 B.n225 B.n224 585
R520 B.n223 B.n144 585
R521 B.n222 B.n221 585
R522 B.n220 B.n145 585
R523 B.n219 B.n218 585
R524 B.n217 B.n146 585
R525 B.n216 B.n215 585
R526 B.n214 B.n147 585
R527 B.n213 B.n212 585
R528 B.n211 B.n148 585
R529 B.n210 B.n209 585
R530 B.n208 B.n149 585
R531 B.n207 B.n206 585
R532 B.n205 B.n150 585
R533 B.n204 B.n203 585
R534 B.n202 B.n151 585
R535 B.n201 B.n200 585
R536 B.n199 B.n152 585
R537 B.n198 B.n197 585
R538 B.n196 B.n153 585
R539 B.n195 B.n194 585
R540 B.n193 B.n154 585
R541 B.n192 B.n191 585
R542 B.n190 B.n155 585
R543 B.n189 B.n188 585
R544 B.n187 B.n156 585
R545 B.n186 B.n185 585
R546 B.n184 B.n157 585
R547 B.n183 B.n182 585
R548 B.n181 B.n158 585
R549 B.n180 B.n179 585
R550 B.n178 B.n159 585
R551 B.n177 B.n176 585
R552 B.n175 B.n160 585
R553 B.n174 B.n173 585
R554 B.n172 B.n161 585
R555 B.n171 B.n170 585
R556 B.n169 B.n162 585
R557 B.n168 B.n167 585
R558 B.n166 B.n163 585
R559 B.n165 B.n164 585
R560 B.n2 B.n0 585
R561 B.n633 B.n1 585
R562 B.n632 B.n631 585
R563 B.n630 B.n3 585
R564 B.n629 B.n628 585
R565 B.n627 B.n4 585
R566 B.n626 B.n625 585
R567 B.n624 B.n5 585
R568 B.n623 B.n622 585
R569 B.n621 B.n6 585
R570 B.n620 B.n619 585
R571 B.n618 B.n7 585
R572 B.n617 B.n616 585
R573 B.n615 B.n8 585
R574 B.n614 B.n613 585
R575 B.n612 B.n9 585
R576 B.n611 B.n610 585
R577 B.n609 B.n10 585
R578 B.n608 B.n607 585
R579 B.n606 B.n11 585
R580 B.n605 B.n604 585
R581 B.n603 B.n12 585
R582 B.n602 B.n601 585
R583 B.n600 B.n13 585
R584 B.n599 B.n598 585
R585 B.n597 B.n14 585
R586 B.n596 B.n595 585
R587 B.n594 B.n15 585
R588 B.n593 B.n592 585
R589 B.n591 B.n16 585
R590 B.n590 B.n589 585
R591 B.n588 B.n17 585
R592 B.n587 B.n586 585
R593 B.n585 B.n18 585
R594 B.n584 B.n583 585
R595 B.n582 B.n19 585
R596 B.n581 B.n580 585
R597 B.n579 B.n20 585
R598 B.n578 B.n577 585
R599 B.n576 B.n21 585
R600 B.n575 B.n574 585
R601 B.n573 B.n22 585
R602 B.n572 B.n571 585
R603 B.n570 B.n23 585
R604 B.n569 B.n568 585
R605 B.n567 B.n24 585
R606 B.n566 B.n565 585
R607 B.n564 B.n25 585
R608 B.n563 B.n562 585
R609 B.n561 B.n26 585
R610 B.n560 B.n559 585
R611 B.n558 B.n27 585
R612 B.n557 B.n556 585
R613 B.n555 B.n28 585
R614 B.n554 B.n553 585
R615 B.n552 B.n29 585
R616 B.n551 B.n550 585
R617 B.n549 B.n30 585
R618 B.n548 B.n547 585
R619 B.n546 B.n31 585
R620 B.n545 B.n544 585
R621 B.n543 B.n32 585
R622 B.n542 B.n541 585
R623 B.n540 B.n33 585
R624 B.n539 B.n538 585
R625 B.n635 B.n634 585
R626 B.n257 B.n132 540.549
R627 B.n538 B.n537 540.549
R628 B.n303 B.n302 540.549
R629 B.n495 B.n52 540.549
R630 B.n285 B.t9 209.823
R631 B.n127 B.t3 209.823
R632 B.n40 B.t0 209.823
R633 B.n47 B.t6 209.823
R634 B.n257 B.n256 163.367
R635 B.n256 B.n255 163.367
R636 B.n255 B.n134 163.367
R637 B.n251 B.n134 163.367
R638 B.n251 B.n250 163.367
R639 B.n250 B.n249 163.367
R640 B.n249 B.n136 163.367
R641 B.n245 B.n136 163.367
R642 B.n245 B.n244 163.367
R643 B.n244 B.n243 163.367
R644 B.n243 B.n138 163.367
R645 B.n239 B.n138 163.367
R646 B.n239 B.n238 163.367
R647 B.n238 B.n237 163.367
R648 B.n237 B.n140 163.367
R649 B.n233 B.n140 163.367
R650 B.n233 B.n232 163.367
R651 B.n232 B.n231 163.367
R652 B.n231 B.n142 163.367
R653 B.n227 B.n142 163.367
R654 B.n227 B.n226 163.367
R655 B.n226 B.n225 163.367
R656 B.n225 B.n144 163.367
R657 B.n221 B.n144 163.367
R658 B.n221 B.n220 163.367
R659 B.n220 B.n219 163.367
R660 B.n219 B.n146 163.367
R661 B.n215 B.n146 163.367
R662 B.n215 B.n214 163.367
R663 B.n214 B.n213 163.367
R664 B.n213 B.n148 163.367
R665 B.n209 B.n148 163.367
R666 B.n209 B.n208 163.367
R667 B.n208 B.n207 163.367
R668 B.n207 B.n150 163.367
R669 B.n203 B.n150 163.367
R670 B.n203 B.n202 163.367
R671 B.n202 B.n201 163.367
R672 B.n201 B.n152 163.367
R673 B.n197 B.n152 163.367
R674 B.n197 B.n196 163.367
R675 B.n196 B.n195 163.367
R676 B.n195 B.n154 163.367
R677 B.n191 B.n154 163.367
R678 B.n191 B.n190 163.367
R679 B.n190 B.n189 163.367
R680 B.n189 B.n156 163.367
R681 B.n185 B.n156 163.367
R682 B.n185 B.n184 163.367
R683 B.n184 B.n183 163.367
R684 B.n183 B.n158 163.367
R685 B.n179 B.n158 163.367
R686 B.n179 B.n178 163.367
R687 B.n178 B.n177 163.367
R688 B.n177 B.n160 163.367
R689 B.n173 B.n160 163.367
R690 B.n173 B.n172 163.367
R691 B.n172 B.n171 163.367
R692 B.n171 B.n162 163.367
R693 B.n167 B.n162 163.367
R694 B.n167 B.n166 163.367
R695 B.n166 B.n165 163.367
R696 B.n165 B.n2 163.367
R697 B.n634 B.n2 163.367
R698 B.n634 B.n633 163.367
R699 B.n633 B.n632 163.367
R700 B.n632 B.n3 163.367
R701 B.n628 B.n3 163.367
R702 B.n628 B.n627 163.367
R703 B.n627 B.n626 163.367
R704 B.n626 B.n5 163.367
R705 B.n622 B.n5 163.367
R706 B.n622 B.n621 163.367
R707 B.n621 B.n620 163.367
R708 B.n620 B.n7 163.367
R709 B.n616 B.n7 163.367
R710 B.n616 B.n615 163.367
R711 B.n615 B.n614 163.367
R712 B.n614 B.n9 163.367
R713 B.n610 B.n9 163.367
R714 B.n610 B.n609 163.367
R715 B.n609 B.n608 163.367
R716 B.n608 B.n11 163.367
R717 B.n604 B.n11 163.367
R718 B.n604 B.n603 163.367
R719 B.n603 B.n602 163.367
R720 B.n602 B.n13 163.367
R721 B.n598 B.n13 163.367
R722 B.n598 B.n597 163.367
R723 B.n597 B.n596 163.367
R724 B.n596 B.n15 163.367
R725 B.n592 B.n15 163.367
R726 B.n592 B.n591 163.367
R727 B.n591 B.n590 163.367
R728 B.n590 B.n17 163.367
R729 B.n586 B.n17 163.367
R730 B.n586 B.n585 163.367
R731 B.n585 B.n584 163.367
R732 B.n584 B.n19 163.367
R733 B.n580 B.n19 163.367
R734 B.n580 B.n579 163.367
R735 B.n579 B.n578 163.367
R736 B.n578 B.n21 163.367
R737 B.n574 B.n21 163.367
R738 B.n574 B.n573 163.367
R739 B.n573 B.n572 163.367
R740 B.n572 B.n23 163.367
R741 B.n568 B.n23 163.367
R742 B.n568 B.n567 163.367
R743 B.n567 B.n566 163.367
R744 B.n566 B.n25 163.367
R745 B.n562 B.n25 163.367
R746 B.n562 B.n561 163.367
R747 B.n561 B.n560 163.367
R748 B.n560 B.n27 163.367
R749 B.n556 B.n27 163.367
R750 B.n556 B.n555 163.367
R751 B.n555 B.n554 163.367
R752 B.n554 B.n29 163.367
R753 B.n550 B.n29 163.367
R754 B.n550 B.n549 163.367
R755 B.n549 B.n548 163.367
R756 B.n548 B.n31 163.367
R757 B.n544 B.n31 163.367
R758 B.n544 B.n543 163.367
R759 B.n543 B.n542 163.367
R760 B.n542 B.n33 163.367
R761 B.n538 B.n33 163.367
R762 B.n261 B.n132 163.367
R763 B.n262 B.n261 163.367
R764 B.n263 B.n262 163.367
R765 B.n263 B.n130 163.367
R766 B.n267 B.n130 163.367
R767 B.n268 B.n267 163.367
R768 B.n269 B.n268 163.367
R769 B.n269 B.n126 163.367
R770 B.n274 B.n126 163.367
R771 B.n275 B.n274 163.367
R772 B.n276 B.n275 163.367
R773 B.n276 B.n124 163.367
R774 B.n280 B.n124 163.367
R775 B.n281 B.n280 163.367
R776 B.n282 B.n281 163.367
R777 B.n282 B.n122 163.367
R778 B.n289 B.n122 163.367
R779 B.n290 B.n289 163.367
R780 B.n291 B.n290 163.367
R781 B.n291 B.n120 163.367
R782 B.n295 B.n120 163.367
R783 B.n296 B.n295 163.367
R784 B.n297 B.n296 163.367
R785 B.n297 B.n118 163.367
R786 B.n301 B.n118 163.367
R787 B.n302 B.n301 163.367
R788 B.n303 B.n116 163.367
R789 B.n307 B.n116 163.367
R790 B.n308 B.n307 163.367
R791 B.n309 B.n308 163.367
R792 B.n309 B.n114 163.367
R793 B.n313 B.n114 163.367
R794 B.n314 B.n313 163.367
R795 B.n315 B.n314 163.367
R796 B.n315 B.n112 163.367
R797 B.n319 B.n112 163.367
R798 B.n320 B.n319 163.367
R799 B.n321 B.n320 163.367
R800 B.n321 B.n110 163.367
R801 B.n325 B.n110 163.367
R802 B.n326 B.n325 163.367
R803 B.n327 B.n326 163.367
R804 B.n327 B.n108 163.367
R805 B.n331 B.n108 163.367
R806 B.n332 B.n331 163.367
R807 B.n333 B.n332 163.367
R808 B.n333 B.n106 163.367
R809 B.n337 B.n106 163.367
R810 B.n338 B.n337 163.367
R811 B.n339 B.n338 163.367
R812 B.n339 B.n104 163.367
R813 B.n343 B.n104 163.367
R814 B.n344 B.n343 163.367
R815 B.n345 B.n344 163.367
R816 B.n345 B.n102 163.367
R817 B.n349 B.n102 163.367
R818 B.n350 B.n349 163.367
R819 B.n351 B.n350 163.367
R820 B.n351 B.n100 163.367
R821 B.n355 B.n100 163.367
R822 B.n356 B.n355 163.367
R823 B.n357 B.n356 163.367
R824 B.n357 B.n98 163.367
R825 B.n361 B.n98 163.367
R826 B.n362 B.n361 163.367
R827 B.n363 B.n362 163.367
R828 B.n363 B.n96 163.367
R829 B.n367 B.n96 163.367
R830 B.n368 B.n367 163.367
R831 B.n369 B.n368 163.367
R832 B.n369 B.n94 163.367
R833 B.n373 B.n94 163.367
R834 B.n374 B.n373 163.367
R835 B.n375 B.n374 163.367
R836 B.n375 B.n92 163.367
R837 B.n379 B.n92 163.367
R838 B.n380 B.n379 163.367
R839 B.n381 B.n380 163.367
R840 B.n381 B.n90 163.367
R841 B.n385 B.n90 163.367
R842 B.n386 B.n385 163.367
R843 B.n387 B.n386 163.367
R844 B.n387 B.n88 163.367
R845 B.n391 B.n88 163.367
R846 B.n392 B.n391 163.367
R847 B.n393 B.n392 163.367
R848 B.n393 B.n86 163.367
R849 B.n397 B.n86 163.367
R850 B.n398 B.n397 163.367
R851 B.n399 B.n398 163.367
R852 B.n399 B.n84 163.367
R853 B.n403 B.n84 163.367
R854 B.n404 B.n403 163.367
R855 B.n405 B.n404 163.367
R856 B.n405 B.n82 163.367
R857 B.n409 B.n82 163.367
R858 B.n410 B.n409 163.367
R859 B.n411 B.n410 163.367
R860 B.n411 B.n80 163.367
R861 B.n415 B.n80 163.367
R862 B.n416 B.n415 163.367
R863 B.n417 B.n416 163.367
R864 B.n417 B.n78 163.367
R865 B.n421 B.n78 163.367
R866 B.n422 B.n421 163.367
R867 B.n423 B.n422 163.367
R868 B.n423 B.n76 163.367
R869 B.n427 B.n76 163.367
R870 B.n428 B.n427 163.367
R871 B.n429 B.n428 163.367
R872 B.n429 B.n74 163.367
R873 B.n433 B.n74 163.367
R874 B.n434 B.n433 163.367
R875 B.n435 B.n434 163.367
R876 B.n435 B.n72 163.367
R877 B.n439 B.n72 163.367
R878 B.n440 B.n439 163.367
R879 B.n441 B.n440 163.367
R880 B.n441 B.n70 163.367
R881 B.n445 B.n70 163.367
R882 B.n446 B.n445 163.367
R883 B.n447 B.n446 163.367
R884 B.n447 B.n68 163.367
R885 B.n451 B.n68 163.367
R886 B.n452 B.n451 163.367
R887 B.n453 B.n452 163.367
R888 B.n453 B.n66 163.367
R889 B.n457 B.n66 163.367
R890 B.n458 B.n457 163.367
R891 B.n459 B.n458 163.367
R892 B.n459 B.n64 163.367
R893 B.n463 B.n64 163.367
R894 B.n464 B.n463 163.367
R895 B.n465 B.n464 163.367
R896 B.n465 B.n62 163.367
R897 B.n469 B.n62 163.367
R898 B.n470 B.n469 163.367
R899 B.n471 B.n470 163.367
R900 B.n471 B.n60 163.367
R901 B.n475 B.n60 163.367
R902 B.n476 B.n475 163.367
R903 B.n477 B.n476 163.367
R904 B.n477 B.n58 163.367
R905 B.n481 B.n58 163.367
R906 B.n482 B.n481 163.367
R907 B.n483 B.n482 163.367
R908 B.n483 B.n56 163.367
R909 B.n487 B.n56 163.367
R910 B.n488 B.n487 163.367
R911 B.n489 B.n488 163.367
R912 B.n489 B.n54 163.367
R913 B.n493 B.n54 163.367
R914 B.n494 B.n493 163.367
R915 B.n495 B.n494 163.367
R916 B.n537 B.n536 163.367
R917 B.n536 B.n35 163.367
R918 B.n532 B.n35 163.367
R919 B.n532 B.n531 163.367
R920 B.n531 B.n530 163.367
R921 B.n530 B.n37 163.367
R922 B.n526 B.n37 163.367
R923 B.n526 B.n525 163.367
R924 B.n525 B.n524 163.367
R925 B.n524 B.n39 163.367
R926 B.n520 B.n39 163.367
R927 B.n520 B.n519 163.367
R928 B.n519 B.n518 163.367
R929 B.n518 B.n44 163.367
R930 B.n514 B.n44 163.367
R931 B.n514 B.n513 163.367
R932 B.n513 B.n512 163.367
R933 B.n512 B.n46 163.367
R934 B.n507 B.n46 163.367
R935 B.n507 B.n506 163.367
R936 B.n506 B.n505 163.367
R937 B.n505 B.n50 163.367
R938 B.n501 B.n50 163.367
R939 B.n501 B.n500 163.367
R940 B.n500 B.n499 163.367
R941 B.n499 B.n52 163.367
R942 B.n286 B.n285 73.6975
R943 B.n128 B.n127 73.6975
R944 B.n41 B.n40 73.6975
R945 B.n48 B.n47 73.6975
R946 B.n287 B.n286 59.5399
R947 B.n272 B.n128 59.5399
R948 B.n42 B.n41 59.5399
R949 B.n510 B.n48 59.5399
R950 B.n539 B.n34 35.1225
R951 B.n497 B.n496 35.1225
R952 B.n304 B.n117 35.1225
R953 B.n259 B.n258 35.1225
R954 B B.n635 18.0485
R955 B.n535 B.n34 10.6151
R956 B.n535 B.n534 10.6151
R957 B.n534 B.n533 10.6151
R958 B.n533 B.n36 10.6151
R959 B.n529 B.n36 10.6151
R960 B.n529 B.n528 10.6151
R961 B.n528 B.n527 10.6151
R962 B.n527 B.n38 10.6151
R963 B.n523 B.n522 10.6151
R964 B.n522 B.n521 10.6151
R965 B.n521 B.n43 10.6151
R966 B.n517 B.n43 10.6151
R967 B.n517 B.n516 10.6151
R968 B.n516 B.n515 10.6151
R969 B.n515 B.n45 10.6151
R970 B.n511 B.n45 10.6151
R971 B.n509 B.n508 10.6151
R972 B.n508 B.n49 10.6151
R973 B.n504 B.n49 10.6151
R974 B.n504 B.n503 10.6151
R975 B.n503 B.n502 10.6151
R976 B.n502 B.n51 10.6151
R977 B.n498 B.n51 10.6151
R978 B.n498 B.n497 10.6151
R979 B.n305 B.n304 10.6151
R980 B.n306 B.n305 10.6151
R981 B.n306 B.n115 10.6151
R982 B.n310 B.n115 10.6151
R983 B.n311 B.n310 10.6151
R984 B.n312 B.n311 10.6151
R985 B.n312 B.n113 10.6151
R986 B.n316 B.n113 10.6151
R987 B.n317 B.n316 10.6151
R988 B.n318 B.n317 10.6151
R989 B.n318 B.n111 10.6151
R990 B.n322 B.n111 10.6151
R991 B.n323 B.n322 10.6151
R992 B.n324 B.n323 10.6151
R993 B.n324 B.n109 10.6151
R994 B.n328 B.n109 10.6151
R995 B.n329 B.n328 10.6151
R996 B.n330 B.n329 10.6151
R997 B.n330 B.n107 10.6151
R998 B.n334 B.n107 10.6151
R999 B.n335 B.n334 10.6151
R1000 B.n336 B.n335 10.6151
R1001 B.n336 B.n105 10.6151
R1002 B.n340 B.n105 10.6151
R1003 B.n341 B.n340 10.6151
R1004 B.n342 B.n341 10.6151
R1005 B.n342 B.n103 10.6151
R1006 B.n346 B.n103 10.6151
R1007 B.n347 B.n346 10.6151
R1008 B.n348 B.n347 10.6151
R1009 B.n348 B.n101 10.6151
R1010 B.n352 B.n101 10.6151
R1011 B.n353 B.n352 10.6151
R1012 B.n354 B.n353 10.6151
R1013 B.n354 B.n99 10.6151
R1014 B.n358 B.n99 10.6151
R1015 B.n359 B.n358 10.6151
R1016 B.n360 B.n359 10.6151
R1017 B.n360 B.n97 10.6151
R1018 B.n364 B.n97 10.6151
R1019 B.n365 B.n364 10.6151
R1020 B.n366 B.n365 10.6151
R1021 B.n366 B.n95 10.6151
R1022 B.n370 B.n95 10.6151
R1023 B.n371 B.n370 10.6151
R1024 B.n372 B.n371 10.6151
R1025 B.n372 B.n93 10.6151
R1026 B.n376 B.n93 10.6151
R1027 B.n377 B.n376 10.6151
R1028 B.n378 B.n377 10.6151
R1029 B.n378 B.n91 10.6151
R1030 B.n382 B.n91 10.6151
R1031 B.n383 B.n382 10.6151
R1032 B.n384 B.n383 10.6151
R1033 B.n384 B.n89 10.6151
R1034 B.n388 B.n89 10.6151
R1035 B.n389 B.n388 10.6151
R1036 B.n390 B.n389 10.6151
R1037 B.n390 B.n87 10.6151
R1038 B.n394 B.n87 10.6151
R1039 B.n395 B.n394 10.6151
R1040 B.n396 B.n395 10.6151
R1041 B.n396 B.n85 10.6151
R1042 B.n400 B.n85 10.6151
R1043 B.n401 B.n400 10.6151
R1044 B.n402 B.n401 10.6151
R1045 B.n402 B.n83 10.6151
R1046 B.n406 B.n83 10.6151
R1047 B.n407 B.n406 10.6151
R1048 B.n408 B.n407 10.6151
R1049 B.n408 B.n81 10.6151
R1050 B.n412 B.n81 10.6151
R1051 B.n413 B.n412 10.6151
R1052 B.n414 B.n413 10.6151
R1053 B.n414 B.n79 10.6151
R1054 B.n418 B.n79 10.6151
R1055 B.n419 B.n418 10.6151
R1056 B.n420 B.n419 10.6151
R1057 B.n420 B.n77 10.6151
R1058 B.n424 B.n77 10.6151
R1059 B.n425 B.n424 10.6151
R1060 B.n426 B.n425 10.6151
R1061 B.n426 B.n75 10.6151
R1062 B.n430 B.n75 10.6151
R1063 B.n431 B.n430 10.6151
R1064 B.n432 B.n431 10.6151
R1065 B.n432 B.n73 10.6151
R1066 B.n436 B.n73 10.6151
R1067 B.n437 B.n436 10.6151
R1068 B.n438 B.n437 10.6151
R1069 B.n438 B.n71 10.6151
R1070 B.n442 B.n71 10.6151
R1071 B.n443 B.n442 10.6151
R1072 B.n444 B.n443 10.6151
R1073 B.n444 B.n69 10.6151
R1074 B.n448 B.n69 10.6151
R1075 B.n449 B.n448 10.6151
R1076 B.n450 B.n449 10.6151
R1077 B.n450 B.n67 10.6151
R1078 B.n454 B.n67 10.6151
R1079 B.n455 B.n454 10.6151
R1080 B.n456 B.n455 10.6151
R1081 B.n456 B.n65 10.6151
R1082 B.n460 B.n65 10.6151
R1083 B.n461 B.n460 10.6151
R1084 B.n462 B.n461 10.6151
R1085 B.n462 B.n63 10.6151
R1086 B.n466 B.n63 10.6151
R1087 B.n467 B.n466 10.6151
R1088 B.n468 B.n467 10.6151
R1089 B.n468 B.n61 10.6151
R1090 B.n472 B.n61 10.6151
R1091 B.n473 B.n472 10.6151
R1092 B.n474 B.n473 10.6151
R1093 B.n474 B.n59 10.6151
R1094 B.n478 B.n59 10.6151
R1095 B.n479 B.n478 10.6151
R1096 B.n480 B.n479 10.6151
R1097 B.n480 B.n57 10.6151
R1098 B.n484 B.n57 10.6151
R1099 B.n485 B.n484 10.6151
R1100 B.n486 B.n485 10.6151
R1101 B.n486 B.n55 10.6151
R1102 B.n490 B.n55 10.6151
R1103 B.n491 B.n490 10.6151
R1104 B.n492 B.n491 10.6151
R1105 B.n492 B.n53 10.6151
R1106 B.n496 B.n53 10.6151
R1107 B.n260 B.n259 10.6151
R1108 B.n260 B.n131 10.6151
R1109 B.n264 B.n131 10.6151
R1110 B.n265 B.n264 10.6151
R1111 B.n266 B.n265 10.6151
R1112 B.n266 B.n129 10.6151
R1113 B.n270 B.n129 10.6151
R1114 B.n271 B.n270 10.6151
R1115 B.n273 B.n125 10.6151
R1116 B.n277 B.n125 10.6151
R1117 B.n278 B.n277 10.6151
R1118 B.n279 B.n278 10.6151
R1119 B.n279 B.n123 10.6151
R1120 B.n283 B.n123 10.6151
R1121 B.n284 B.n283 10.6151
R1122 B.n288 B.n284 10.6151
R1123 B.n292 B.n121 10.6151
R1124 B.n293 B.n292 10.6151
R1125 B.n294 B.n293 10.6151
R1126 B.n294 B.n119 10.6151
R1127 B.n298 B.n119 10.6151
R1128 B.n299 B.n298 10.6151
R1129 B.n300 B.n299 10.6151
R1130 B.n300 B.n117 10.6151
R1131 B.n258 B.n133 10.6151
R1132 B.n254 B.n133 10.6151
R1133 B.n254 B.n253 10.6151
R1134 B.n253 B.n252 10.6151
R1135 B.n252 B.n135 10.6151
R1136 B.n248 B.n135 10.6151
R1137 B.n248 B.n247 10.6151
R1138 B.n247 B.n246 10.6151
R1139 B.n246 B.n137 10.6151
R1140 B.n242 B.n137 10.6151
R1141 B.n242 B.n241 10.6151
R1142 B.n241 B.n240 10.6151
R1143 B.n240 B.n139 10.6151
R1144 B.n236 B.n139 10.6151
R1145 B.n236 B.n235 10.6151
R1146 B.n235 B.n234 10.6151
R1147 B.n234 B.n141 10.6151
R1148 B.n230 B.n141 10.6151
R1149 B.n230 B.n229 10.6151
R1150 B.n229 B.n228 10.6151
R1151 B.n228 B.n143 10.6151
R1152 B.n224 B.n143 10.6151
R1153 B.n224 B.n223 10.6151
R1154 B.n223 B.n222 10.6151
R1155 B.n222 B.n145 10.6151
R1156 B.n218 B.n145 10.6151
R1157 B.n218 B.n217 10.6151
R1158 B.n217 B.n216 10.6151
R1159 B.n216 B.n147 10.6151
R1160 B.n212 B.n147 10.6151
R1161 B.n212 B.n211 10.6151
R1162 B.n211 B.n210 10.6151
R1163 B.n210 B.n149 10.6151
R1164 B.n206 B.n149 10.6151
R1165 B.n206 B.n205 10.6151
R1166 B.n205 B.n204 10.6151
R1167 B.n204 B.n151 10.6151
R1168 B.n200 B.n151 10.6151
R1169 B.n200 B.n199 10.6151
R1170 B.n199 B.n198 10.6151
R1171 B.n198 B.n153 10.6151
R1172 B.n194 B.n153 10.6151
R1173 B.n194 B.n193 10.6151
R1174 B.n193 B.n192 10.6151
R1175 B.n192 B.n155 10.6151
R1176 B.n188 B.n155 10.6151
R1177 B.n188 B.n187 10.6151
R1178 B.n187 B.n186 10.6151
R1179 B.n186 B.n157 10.6151
R1180 B.n182 B.n157 10.6151
R1181 B.n182 B.n181 10.6151
R1182 B.n181 B.n180 10.6151
R1183 B.n180 B.n159 10.6151
R1184 B.n176 B.n159 10.6151
R1185 B.n176 B.n175 10.6151
R1186 B.n175 B.n174 10.6151
R1187 B.n174 B.n161 10.6151
R1188 B.n170 B.n161 10.6151
R1189 B.n170 B.n169 10.6151
R1190 B.n169 B.n168 10.6151
R1191 B.n168 B.n163 10.6151
R1192 B.n164 B.n163 10.6151
R1193 B.n164 B.n0 10.6151
R1194 B.n631 B.n1 10.6151
R1195 B.n631 B.n630 10.6151
R1196 B.n630 B.n629 10.6151
R1197 B.n629 B.n4 10.6151
R1198 B.n625 B.n4 10.6151
R1199 B.n625 B.n624 10.6151
R1200 B.n624 B.n623 10.6151
R1201 B.n623 B.n6 10.6151
R1202 B.n619 B.n6 10.6151
R1203 B.n619 B.n618 10.6151
R1204 B.n618 B.n617 10.6151
R1205 B.n617 B.n8 10.6151
R1206 B.n613 B.n8 10.6151
R1207 B.n613 B.n612 10.6151
R1208 B.n612 B.n611 10.6151
R1209 B.n611 B.n10 10.6151
R1210 B.n607 B.n10 10.6151
R1211 B.n607 B.n606 10.6151
R1212 B.n606 B.n605 10.6151
R1213 B.n605 B.n12 10.6151
R1214 B.n601 B.n12 10.6151
R1215 B.n601 B.n600 10.6151
R1216 B.n600 B.n599 10.6151
R1217 B.n599 B.n14 10.6151
R1218 B.n595 B.n14 10.6151
R1219 B.n595 B.n594 10.6151
R1220 B.n594 B.n593 10.6151
R1221 B.n593 B.n16 10.6151
R1222 B.n589 B.n16 10.6151
R1223 B.n589 B.n588 10.6151
R1224 B.n588 B.n587 10.6151
R1225 B.n587 B.n18 10.6151
R1226 B.n583 B.n18 10.6151
R1227 B.n583 B.n582 10.6151
R1228 B.n582 B.n581 10.6151
R1229 B.n581 B.n20 10.6151
R1230 B.n577 B.n20 10.6151
R1231 B.n577 B.n576 10.6151
R1232 B.n576 B.n575 10.6151
R1233 B.n575 B.n22 10.6151
R1234 B.n571 B.n22 10.6151
R1235 B.n571 B.n570 10.6151
R1236 B.n570 B.n569 10.6151
R1237 B.n569 B.n24 10.6151
R1238 B.n565 B.n24 10.6151
R1239 B.n565 B.n564 10.6151
R1240 B.n564 B.n563 10.6151
R1241 B.n563 B.n26 10.6151
R1242 B.n559 B.n26 10.6151
R1243 B.n559 B.n558 10.6151
R1244 B.n558 B.n557 10.6151
R1245 B.n557 B.n28 10.6151
R1246 B.n553 B.n28 10.6151
R1247 B.n553 B.n552 10.6151
R1248 B.n552 B.n551 10.6151
R1249 B.n551 B.n30 10.6151
R1250 B.n547 B.n30 10.6151
R1251 B.n547 B.n546 10.6151
R1252 B.n546 B.n545 10.6151
R1253 B.n545 B.n32 10.6151
R1254 B.n541 B.n32 10.6151
R1255 B.n541 B.n540 10.6151
R1256 B.n540 B.n539 10.6151
R1257 B.n523 B.n42 6.5566
R1258 B.n511 B.n510 6.5566
R1259 B.n273 B.n272 6.5566
R1260 B.n288 B.n287 6.5566
R1261 B.n42 B.n38 4.05904
R1262 B.n510 B.n509 4.05904
R1263 B.n272 B.n271 4.05904
R1264 B.n287 B.n121 4.05904
R1265 B.n635 B.n0 2.81026
R1266 B.n635 B.n1 2.81026
C0 B VDD1 1.61601f
C1 VDD2 VTAIL 5.25415f
C2 B VN 1.25721f
C3 B w_n4770_n1148# 8.467f
C4 B VTAIL 1.33012f
C5 VP VDD1 1.58677f
C6 VP VN 6.67489f
C7 VP w_n4770_n1148# 10.407f
C8 B VDD2 1.74024f
C9 VP VTAIL 2.87679f
C10 VP VDD2 0.622352f
C11 VN VDD1 0.161059f
C12 w_n4770_n1148# VDD1 1.93043f
C13 VTAIL VDD1 5.1939f
C14 w_n4770_n1148# VN 9.793281f
C15 B VP 2.3029f
C16 VTAIL VN 2.86268f
C17 w_n4770_n1148# VTAIL 1.76773f
C18 VDD2 VDD1 2.22911f
C19 VDD2 VN 1.13029f
C20 w_n4770_n1148# VDD2 2.08051f
C21 VDD2 VSUBS 1.885908f
C22 VDD1 VSUBS 2.386493f
C23 VTAIL VSUBS 0.65284f
C24 VN VSUBS 8.553889f
C25 VP VSUBS 3.805615f
C26 B VSUBS 4.718087f
C27 w_n4770_n1148# VSUBS 70.6914f
C28 B.n0 VSUBS 0.008171f
C29 B.n1 VSUBS 0.008171f
C30 B.n2 VSUBS 0.012921f
C31 B.n3 VSUBS 0.012921f
C32 B.n4 VSUBS 0.012921f
C33 B.n5 VSUBS 0.012921f
C34 B.n6 VSUBS 0.012921f
C35 B.n7 VSUBS 0.012921f
C36 B.n8 VSUBS 0.012921f
C37 B.n9 VSUBS 0.012921f
C38 B.n10 VSUBS 0.012921f
C39 B.n11 VSUBS 0.012921f
C40 B.n12 VSUBS 0.012921f
C41 B.n13 VSUBS 0.012921f
C42 B.n14 VSUBS 0.012921f
C43 B.n15 VSUBS 0.012921f
C44 B.n16 VSUBS 0.012921f
C45 B.n17 VSUBS 0.012921f
C46 B.n18 VSUBS 0.012921f
C47 B.n19 VSUBS 0.012921f
C48 B.n20 VSUBS 0.012921f
C49 B.n21 VSUBS 0.012921f
C50 B.n22 VSUBS 0.012921f
C51 B.n23 VSUBS 0.012921f
C52 B.n24 VSUBS 0.012921f
C53 B.n25 VSUBS 0.012921f
C54 B.n26 VSUBS 0.012921f
C55 B.n27 VSUBS 0.012921f
C56 B.n28 VSUBS 0.012921f
C57 B.n29 VSUBS 0.012921f
C58 B.n30 VSUBS 0.012921f
C59 B.n31 VSUBS 0.012921f
C60 B.n32 VSUBS 0.012921f
C61 B.n33 VSUBS 0.012921f
C62 B.n34 VSUBS 0.032097f
C63 B.n35 VSUBS 0.012921f
C64 B.n36 VSUBS 0.012921f
C65 B.n37 VSUBS 0.012921f
C66 B.n38 VSUBS 0.008931f
C67 B.n39 VSUBS 0.012921f
C68 B.t2 VSUBS 0.032131f
C69 B.t1 VSUBS 0.039244f
C70 B.t0 VSUBS 0.290241f
C71 B.n40 VSUBS 0.130024f
C72 B.n41 VSUBS 0.088117f
C73 B.n42 VSUBS 0.029937f
C74 B.n43 VSUBS 0.012921f
C75 B.n44 VSUBS 0.012921f
C76 B.n45 VSUBS 0.012921f
C77 B.n46 VSUBS 0.012921f
C78 B.t8 VSUBS 0.032131f
C79 B.t7 VSUBS 0.039244f
C80 B.t6 VSUBS 0.290241f
C81 B.n47 VSUBS 0.130024f
C82 B.n48 VSUBS 0.088117f
C83 B.n49 VSUBS 0.012921f
C84 B.n50 VSUBS 0.012921f
C85 B.n51 VSUBS 0.012921f
C86 B.n52 VSUBS 0.032097f
C87 B.n53 VSUBS 0.012921f
C88 B.n54 VSUBS 0.012921f
C89 B.n55 VSUBS 0.012921f
C90 B.n56 VSUBS 0.012921f
C91 B.n57 VSUBS 0.012921f
C92 B.n58 VSUBS 0.012921f
C93 B.n59 VSUBS 0.012921f
C94 B.n60 VSUBS 0.012921f
C95 B.n61 VSUBS 0.012921f
C96 B.n62 VSUBS 0.012921f
C97 B.n63 VSUBS 0.012921f
C98 B.n64 VSUBS 0.012921f
C99 B.n65 VSUBS 0.012921f
C100 B.n66 VSUBS 0.012921f
C101 B.n67 VSUBS 0.012921f
C102 B.n68 VSUBS 0.012921f
C103 B.n69 VSUBS 0.012921f
C104 B.n70 VSUBS 0.012921f
C105 B.n71 VSUBS 0.012921f
C106 B.n72 VSUBS 0.012921f
C107 B.n73 VSUBS 0.012921f
C108 B.n74 VSUBS 0.012921f
C109 B.n75 VSUBS 0.012921f
C110 B.n76 VSUBS 0.012921f
C111 B.n77 VSUBS 0.012921f
C112 B.n78 VSUBS 0.012921f
C113 B.n79 VSUBS 0.012921f
C114 B.n80 VSUBS 0.012921f
C115 B.n81 VSUBS 0.012921f
C116 B.n82 VSUBS 0.012921f
C117 B.n83 VSUBS 0.012921f
C118 B.n84 VSUBS 0.012921f
C119 B.n85 VSUBS 0.012921f
C120 B.n86 VSUBS 0.012921f
C121 B.n87 VSUBS 0.012921f
C122 B.n88 VSUBS 0.012921f
C123 B.n89 VSUBS 0.012921f
C124 B.n90 VSUBS 0.012921f
C125 B.n91 VSUBS 0.012921f
C126 B.n92 VSUBS 0.012921f
C127 B.n93 VSUBS 0.012921f
C128 B.n94 VSUBS 0.012921f
C129 B.n95 VSUBS 0.012921f
C130 B.n96 VSUBS 0.012921f
C131 B.n97 VSUBS 0.012921f
C132 B.n98 VSUBS 0.012921f
C133 B.n99 VSUBS 0.012921f
C134 B.n100 VSUBS 0.012921f
C135 B.n101 VSUBS 0.012921f
C136 B.n102 VSUBS 0.012921f
C137 B.n103 VSUBS 0.012921f
C138 B.n104 VSUBS 0.012921f
C139 B.n105 VSUBS 0.012921f
C140 B.n106 VSUBS 0.012921f
C141 B.n107 VSUBS 0.012921f
C142 B.n108 VSUBS 0.012921f
C143 B.n109 VSUBS 0.012921f
C144 B.n110 VSUBS 0.012921f
C145 B.n111 VSUBS 0.012921f
C146 B.n112 VSUBS 0.012921f
C147 B.n113 VSUBS 0.012921f
C148 B.n114 VSUBS 0.012921f
C149 B.n115 VSUBS 0.012921f
C150 B.n116 VSUBS 0.012921f
C151 B.n117 VSUBS 0.032097f
C152 B.n118 VSUBS 0.012921f
C153 B.n119 VSUBS 0.012921f
C154 B.n120 VSUBS 0.012921f
C155 B.n121 VSUBS 0.008931f
C156 B.n122 VSUBS 0.012921f
C157 B.n123 VSUBS 0.012921f
C158 B.n124 VSUBS 0.012921f
C159 B.n125 VSUBS 0.012921f
C160 B.n126 VSUBS 0.012921f
C161 B.t4 VSUBS 0.032131f
C162 B.t5 VSUBS 0.039244f
C163 B.t3 VSUBS 0.290241f
C164 B.n127 VSUBS 0.130024f
C165 B.n128 VSUBS 0.088117f
C166 B.n129 VSUBS 0.012921f
C167 B.n130 VSUBS 0.012921f
C168 B.n131 VSUBS 0.012921f
C169 B.n132 VSUBS 0.032097f
C170 B.n133 VSUBS 0.012921f
C171 B.n134 VSUBS 0.012921f
C172 B.n135 VSUBS 0.012921f
C173 B.n136 VSUBS 0.012921f
C174 B.n137 VSUBS 0.012921f
C175 B.n138 VSUBS 0.012921f
C176 B.n139 VSUBS 0.012921f
C177 B.n140 VSUBS 0.012921f
C178 B.n141 VSUBS 0.012921f
C179 B.n142 VSUBS 0.012921f
C180 B.n143 VSUBS 0.012921f
C181 B.n144 VSUBS 0.012921f
C182 B.n145 VSUBS 0.012921f
C183 B.n146 VSUBS 0.012921f
C184 B.n147 VSUBS 0.012921f
C185 B.n148 VSUBS 0.012921f
C186 B.n149 VSUBS 0.012921f
C187 B.n150 VSUBS 0.012921f
C188 B.n151 VSUBS 0.012921f
C189 B.n152 VSUBS 0.012921f
C190 B.n153 VSUBS 0.012921f
C191 B.n154 VSUBS 0.012921f
C192 B.n155 VSUBS 0.012921f
C193 B.n156 VSUBS 0.012921f
C194 B.n157 VSUBS 0.012921f
C195 B.n158 VSUBS 0.012921f
C196 B.n159 VSUBS 0.012921f
C197 B.n160 VSUBS 0.012921f
C198 B.n161 VSUBS 0.012921f
C199 B.n162 VSUBS 0.012921f
C200 B.n163 VSUBS 0.012921f
C201 B.n164 VSUBS 0.012921f
C202 B.n165 VSUBS 0.012921f
C203 B.n166 VSUBS 0.012921f
C204 B.n167 VSUBS 0.012921f
C205 B.n168 VSUBS 0.012921f
C206 B.n169 VSUBS 0.012921f
C207 B.n170 VSUBS 0.012921f
C208 B.n171 VSUBS 0.012921f
C209 B.n172 VSUBS 0.012921f
C210 B.n173 VSUBS 0.012921f
C211 B.n174 VSUBS 0.012921f
C212 B.n175 VSUBS 0.012921f
C213 B.n176 VSUBS 0.012921f
C214 B.n177 VSUBS 0.012921f
C215 B.n178 VSUBS 0.012921f
C216 B.n179 VSUBS 0.012921f
C217 B.n180 VSUBS 0.012921f
C218 B.n181 VSUBS 0.012921f
C219 B.n182 VSUBS 0.012921f
C220 B.n183 VSUBS 0.012921f
C221 B.n184 VSUBS 0.012921f
C222 B.n185 VSUBS 0.012921f
C223 B.n186 VSUBS 0.012921f
C224 B.n187 VSUBS 0.012921f
C225 B.n188 VSUBS 0.012921f
C226 B.n189 VSUBS 0.012921f
C227 B.n190 VSUBS 0.012921f
C228 B.n191 VSUBS 0.012921f
C229 B.n192 VSUBS 0.012921f
C230 B.n193 VSUBS 0.012921f
C231 B.n194 VSUBS 0.012921f
C232 B.n195 VSUBS 0.012921f
C233 B.n196 VSUBS 0.012921f
C234 B.n197 VSUBS 0.012921f
C235 B.n198 VSUBS 0.012921f
C236 B.n199 VSUBS 0.012921f
C237 B.n200 VSUBS 0.012921f
C238 B.n201 VSUBS 0.012921f
C239 B.n202 VSUBS 0.012921f
C240 B.n203 VSUBS 0.012921f
C241 B.n204 VSUBS 0.012921f
C242 B.n205 VSUBS 0.012921f
C243 B.n206 VSUBS 0.012921f
C244 B.n207 VSUBS 0.012921f
C245 B.n208 VSUBS 0.012921f
C246 B.n209 VSUBS 0.012921f
C247 B.n210 VSUBS 0.012921f
C248 B.n211 VSUBS 0.012921f
C249 B.n212 VSUBS 0.012921f
C250 B.n213 VSUBS 0.012921f
C251 B.n214 VSUBS 0.012921f
C252 B.n215 VSUBS 0.012921f
C253 B.n216 VSUBS 0.012921f
C254 B.n217 VSUBS 0.012921f
C255 B.n218 VSUBS 0.012921f
C256 B.n219 VSUBS 0.012921f
C257 B.n220 VSUBS 0.012921f
C258 B.n221 VSUBS 0.012921f
C259 B.n222 VSUBS 0.012921f
C260 B.n223 VSUBS 0.012921f
C261 B.n224 VSUBS 0.012921f
C262 B.n225 VSUBS 0.012921f
C263 B.n226 VSUBS 0.012921f
C264 B.n227 VSUBS 0.012921f
C265 B.n228 VSUBS 0.012921f
C266 B.n229 VSUBS 0.012921f
C267 B.n230 VSUBS 0.012921f
C268 B.n231 VSUBS 0.012921f
C269 B.n232 VSUBS 0.012921f
C270 B.n233 VSUBS 0.012921f
C271 B.n234 VSUBS 0.012921f
C272 B.n235 VSUBS 0.012921f
C273 B.n236 VSUBS 0.012921f
C274 B.n237 VSUBS 0.012921f
C275 B.n238 VSUBS 0.012921f
C276 B.n239 VSUBS 0.012921f
C277 B.n240 VSUBS 0.012921f
C278 B.n241 VSUBS 0.012921f
C279 B.n242 VSUBS 0.012921f
C280 B.n243 VSUBS 0.012921f
C281 B.n244 VSUBS 0.012921f
C282 B.n245 VSUBS 0.012921f
C283 B.n246 VSUBS 0.012921f
C284 B.n247 VSUBS 0.012921f
C285 B.n248 VSUBS 0.012921f
C286 B.n249 VSUBS 0.012921f
C287 B.n250 VSUBS 0.012921f
C288 B.n251 VSUBS 0.012921f
C289 B.n252 VSUBS 0.012921f
C290 B.n253 VSUBS 0.012921f
C291 B.n254 VSUBS 0.012921f
C292 B.n255 VSUBS 0.012921f
C293 B.n256 VSUBS 0.012921f
C294 B.n257 VSUBS 0.03137f
C295 B.n258 VSUBS 0.03137f
C296 B.n259 VSUBS 0.032097f
C297 B.n260 VSUBS 0.012921f
C298 B.n261 VSUBS 0.012921f
C299 B.n262 VSUBS 0.012921f
C300 B.n263 VSUBS 0.012921f
C301 B.n264 VSUBS 0.012921f
C302 B.n265 VSUBS 0.012921f
C303 B.n266 VSUBS 0.012921f
C304 B.n267 VSUBS 0.012921f
C305 B.n268 VSUBS 0.012921f
C306 B.n269 VSUBS 0.012921f
C307 B.n270 VSUBS 0.012921f
C308 B.n271 VSUBS 0.008931f
C309 B.n272 VSUBS 0.029937f
C310 B.n273 VSUBS 0.010451f
C311 B.n274 VSUBS 0.012921f
C312 B.n275 VSUBS 0.012921f
C313 B.n276 VSUBS 0.012921f
C314 B.n277 VSUBS 0.012921f
C315 B.n278 VSUBS 0.012921f
C316 B.n279 VSUBS 0.012921f
C317 B.n280 VSUBS 0.012921f
C318 B.n281 VSUBS 0.012921f
C319 B.n282 VSUBS 0.012921f
C320 B.n283 VSUBS 0.012921f
C321 B.n284 VSUBS 0.012921f
C322 B.t10 VSUBS 0.032131f
C323 B.t11 VSUBS 0.039244f
C324 B.t9 VSUBS 0.290241f
C325 B.n285 VSUBS 0.130024f
C326 B.n286 VSUBS 0.088117f
C327 B.n287 VSUBS 0.029937f
C328 B.n288 VSUBS 0.010451f
C329 B.n289 VSUBS 0.012921f
C330 B.n290 VSUBS 0.012921f
C331 B.n291 VSUBS 0.012921f
C332 B.n292 VSUBS 0.012921f
C333 B.n293 VSUBS 0.012921f
C334 B.n294 VSUBS 0.012921f
C335 B.n295 VSUBS 0.012921f
C336 B.n296 VSUBS 0.012921f
C337 B.n297 VSUBS 0.012921f
C338 B.n298 VSUBS 0.012921f
C339 B.n299 VSUBS 0.012921f
C340 B.n300 VSUBS 0.012921f
C341 B.n301 VSUBS 0.012921f
C342 B.n302 VSUBS 0.032097f
C343 B.n303 VSUBS 0.03137f
C344 B.n304 VSUBS 0.03137f
C345 B.n305 VSUBS 0.012921f
C346 B.n306 VSUBS 0.012921f
C347 B.n307 VSUBS 0.012921f
C348 B.n308 VSUBS 0.012921f
C349 B.n309 VSUBS 0.012921f
C350 B.n310 VSUBS 0.012921f
C351 B.n311 VSUBS 0.012921f
C352 B.n312 VSUBS 0.012921f
C353 B.n313 VSUBS 0.012921f
C354 B.n314 VSUBS 0.012921f
C355 B.n315 VSUBS 0.012921f
C356 B.n316 VSUBS 0.012921f
C357 B.n317 VSUBS 0.012921f
C358 B.n318 VSUBS 0.012921f
C359 B.n319 VSUBS 0.012921f
C360 B.n320 VSUBS 0.012921f
C361 B.n321 VSUBS 0.012921f
C362 B.n322 VSUBS 0.012921f
C363 B.n323 VSUBS 0.012921f
C364 B.n324 VSUBS 0.012921f
C365 B.n325 VSUBS 0.012921f
C366 B.n326 VSUBS 0.012921f
C367 B.n327 VSUBS 0.012921f
C368 B.n328 VSUBS 0.012921f
C369 B.n329 VSUBS 0.012921f
C370 B.n330 VSUBS 0.012921f
C371 B.n331 VSUBS 0.012921f
C372 B.n332 VSUBS 0.012921f
C373 B.n333 VSUBS 0.012921f
C374 B.n334 VSUBS 0.012921f
C375 B.n335 VSUBS 0.012921f
C376 B.n336 VSUBS 0.012921f
C377 B.n337 VSUBS 0.012921f
C378 B.n338 VSUBS 0.012921f
C379 B.n339 VSUBS 0.012921f
C380 B.n340 VSUBS 0.012921f
C381 B.n341 VSUBS 0.012921f
C382 B.n342 VSUBS 0.012921f
C383 B.n343 VSUBS 0.012921f
C384 B.n344 VSUBS 0.012921f
C385 B.n345 VSUBS 0.012921f
C386 B.n346 VSUBS 0.012921f
C387 B.n347 VSUBS 0.012921f
C388 B.n348 VSUBS 0.012921f
C389 B.n349 VSUBS 0.012921f
C390 B.n350 VSUBS 0.012921f
C391 B.n351 VSUBS 0.012921f
C392 B.n352 VSUBS 0.012921f
C393 B.n353 VSUBS 0.012921f
C394 B.n354 VSUBS 0.012921f
C395 B.n355 VSUBS 0.012921f
C396 B.n356 VSUBS 0.012921f
C397 B.n357 VSUBS 0.012921f
C398 B.n358 VSUBS 0.012921f
C399 B.n359 VSUBS 0.012921f
C400 B.n360 VSUBS 0.012921f
C401 B.n361 VSUBS 0.012921f
C402 B.n362 VSUBS 0.012921f
C403 B.n363 VSUBS 0.012921f
C404 B.n364 VSUBS 0.012921f
C405 B.n365 VSUBS 0.012921f
C406 B.n366 VSUBS 0.012921f
C407 B.n367 VSUBS 0.012921f
C408 B.n368 VSUBS 0.012921f
C409 B.n369 VSUBS 0.012921f
C410 B.n370 VSUBS 0.012921f
C411 B.n371 VSUBS 0.012921f
C412 B.n372 VSUBS 0.012921f
C413 B.n373 VSUBS 0.012921f
C414 B.n374 VSUBS 0.012921f
C415 B.n375 VSUBS 0.012921f
C416 B.n376 VSUBS 0.012921f
C417 B.n377 VSUBS 0.012921f
C418 B.n378 VSUBS 0.012921f
C419 B.n379 VSUBS 0.012921f
C420 B.n380 VSUBS 0.012921f
C421 B.n381 VSUBS 0.012921f
C422 B.n382 VSUBS 0.012921f
C423 B.n383 VSUBS 0.012921f
C424 B.n384 VSUBS 0.012921f
C425 B.n385 VSUBS 0.012921f
C426 B.n386 VSUBS 0.012921f
C427 B.n387 VSUBS 0.012921f
C428 B.n388 VSUBS 0.012921f
C429 B.n389 VSUBS 0.012921f
C430 B.n390 VSUBS 0.012921f
C431 B.n391 VSUBS 0.012921f
C432 B.n392 VSUBS 0.012921f
C433 B.n393 VSUBS 0.012921f
C434 B.n394 VSUBS 0.012921f
C435 B.n395 VSUBS 0.012921f
C436 B.n396 VSUBS 0.012921f
C437 B.n397 VSUBS 0.012921f
C438 B.n398 VSUBS 0.012921f
C439 B.n399 VSUBS 0.012921f
C440 B.n400 VSUBS 0.012921f
C441 B.n401 VSUBS 0.012921f
C442 B.n402 VSUBS 0.012921f
C443 B.n403 VSUBS 0.012921f
C444 B.n404 VSUBS 0.012921f
C445 B.n405 VSUBS 0.012921f
C446 B.n406 VSUBS 0.012921f
C447 B.n407 VSUBS 0.012921f
C448 B.n408 VSUBS 0.012921f
C449 B.n409 VSUBS 0.012921f
C450 B.n410 VSUBS 0.012921f
C451 B.n411 VSUBS 0.012921f
C452 B.n412 VSUBS 0.012921f
C453 B.n413 VSUBS 0.012921f
C454 B.n414 VSUBS 0.012921f
C455 B.n415 VSUBS 0.012921f
C456 B.n416 VSUBS 0.012921f
C457 B.n417 VSUBS 0.012921f
C458 B.n418 VSUBS 0.012921f
C459 B.n419 VSUBS 0.012921f
C460 B.n420 VSUBS 0.012921f
C461 B.n421 VSUBS 0.012921f
C462 B.n422 VSUBS 0.012921f
C463 B.n423 VSUBS 0.012921f
C464 B.n424 VSUBS 0.012921f
C465 B.n425 VSUBS 0.012921f
C466 B.n426 VSUBS 0.012921f
C467 B.n427 VSUBS 0.012921f
C468 B.n428 VSUBS 0.012921f
C469 B.n429 VSUBS 0.012921f
C470 B.n430 VSUBS 0.012921f
C471 B.n431 VSUBS 0.012921f
C472 B.n432 VSUBS 0.012921f
C473 B.n433 VSUBS 0.012921f
C474 B.n434 VSUBS 0.012921f
C475 B.n435 VSUBS 0.012921f
C476 B.n436 VSUBS 0.012921f
C477 B.n437 VSUBS 0.012921f
C478 B.n438 VSUBS 0.012921f
C479 B.n439 VSUBS 0.012921f
C480 B.n440 VSUBS 0.012921f
C481 B.n441 VSUBS 0.012921f
C482 B.n442 VSUBS 0.012921f
C483 B.n443 VSUBS 0.012921f
C484 B.n444 VSUBS 0.012921f
C485 B.n445 VSUBS 0.012921f
C486 B.n446 VSUBS 0.012921f
C487 B.n447 VSUBS 0.012921f
C488 B.n448 VSUBS 0.012921f
C489 B.n449 VSUBS 0.012921f
C490 B.n450 VSUBS 0.012921f
C491 B.n451 VSUBS 0.012921f
C492 B.n452 VSUBS 0.012921f
C493 B.n453 VSUBS 0.012921f
C494 B.n454 VSUBS 0.012921f
C495 B.n455 VSUBS 0.012921f
C496 B.n456 VSUBS 0.012921f
C497 B.n457 VSUBS 0.012921f
C498 B.n458 VSUBS 0.012921f
C499 B.n459 VSUBS 0.012921f
C500 B.n460 VSUBS 0.012921f
C501 B.n461 VSUBS 0.012921f
C502 B.n462 VSUBS 0.012921f
C503 B.n463 VSUBS 0.012921f
C504 B.n464 VSUBS 0.012921f
C505 B.n465 VSUBS 0.012921f
C506 B.n466 VSUBS 0.012921f
C507 B.n467 VSUBS 0.012921f
C508 B.n468 VSUBS 0.012921f
C509 B.n469 VSUBS 0.012921f
C510 B.n470 VSUBS 0.012921f
C511 B.n471 VSUBS 0.012921f
C512 B.n472 VSUBS 0.012921f
C513 B.n473 VSUBS 0.012921f
C514 B.n474 VSUBS 0.012921f
C515 B.n475 VSUBS 0.012921f
C516 B.n476 VSUBS 0.012921f
C517 B.n477 VSUBS 0.012921f
C518 B.n478 VSUBS 0.012921f
C519 B.n479 VSUBS 0.012921f
C520 B.n480 VSUBS 0.012921f
C521 B.n481 VSUBS 0.012921f
C522 B.n482 VSUBS 0.012921f
C523 B.n483 VSUBS 0.012921f
C524 B.n484 VSUBS 0.012921f
C525 B.n485 VSUBS 0.012921f
C526 B.n486 VSUBS 0.012921f
C527 B.n487 VSUBS 0.012921f
C528 B.n488 VSUBS 0.012921f
C529 B.n489 VSUBS 0.012921f
C530 B.n490 VSUBS 0.012921f
C531 B.n491 VSUBS 0.012921f
C532 B.n492 VSUBS 0.012921f
C533 B.n493 VSUBS 0.012921f
C534 B.n494 VSUBS 0.012921f
C535 B.n495 VSUBS 0.03137f
C536 B.n496 VSUBS 0.032789f
C537 B.n497 VSUBS 0.030677f
C538 B.n498 VSUBS 0.012921f
C539 B.n499 VSUBS 0.012921f
C540 B.n500 VSUBS 0.012921f
C541 B.n501 VSUBS 0.012921f
C542 B.n502 VSUBS 0.012921f
C543 B.n503 VSUBS 0.012921f
C544 B.n504 VSUBS 0.012921f
C545 B.n505 VSUBS 0.012921f
C546 B.n506 VSUBS 0.012921f
C547 B.n507 VSUBS 0.012921f
C548 B.n508 VSUBS 0.012921f
C549 B.n509 VSUBS 0.008931f
C550 B.n510 VSUBS 0.029937f
C551 B.n511 VSUBS 0.010451f
C552 B.n512 VSUBS 0.012921f
C553 B.n513 VSUBS 0.012921f
C554 B.n514 VSUBS 0.012921f
C555 B.n515 VSUBS 0.012921f
C556 B.n516 VSUBS 0.012921f
C557 B.n517 VSUBS 0.012921f
C558 B.n518 VSUBS 0.012921f
C559 B.n519 VSUBS 0.012921f
C560 B.n520 VSUBS 0.012921f
C561 B.n521 VSUBS 0.012921f
C562 B.n522 VSUBS 0.012921f
C563 B.n523 VSUBS 0.010451f
C564 B.n524 VSUBS 0.012921f
C565 B.n525 VSUBS 0.012921f
C566 B.n526 VSUBS 0.012921f
C567 B.n527 VSUBS 0.012921f
C568 B.n528 VSUBS 0.012921f
C569 B.n529 VSUBS 0.012921f
C570 B.n530 VSUBS 0.012921f
C571 B.n531 VSUBS 0.012921f
C572 B.n532 VSUBS 0.012921f
C573 B.n533 VSUBS 0.012921f
C574 B.n534 VSUBS 0.012921f
C575 B.n535 VSUBS 0.012921f
C576 B.n536 VSUBS 0.012921f
C577 B.n537 VSUBS 0.032097f
C578 B.n538 VSUBS 0.03137f
C579 B.n539 VSUBS 0.03137f
C580 B.n540 VSUBS 0.012921f
C581 B.n541 VSUBS 0.012921f
C582 B.n542 VSUBS 0.012921f
C583 B.n543 VSUBS 0.012921f
C584 B.n544 VSUBS 0.012921f
C585 B.n545 VSUBS 0.012921f
C586 B.n546 VSUBS 0.012921f
C587 B.n547 VSUBS 0.012921f
C588 B.n548 VSUBS 0.012921f
C589 B.n549 VSUBS 0.012921f
C590 B.n550 VSUBS 0.012921f
C591 B.n551 VSUBS 0.012921f
C592 B.n552 VSUBS 0.012921f
C593 B.n553 VSUBS 0.012921f
C594 B.n554 VSUBS 0.012921f
C595 B.n555 VSUBS 0.012921f
C596 B.n556 VSUBS 0.012921f
C597 B.n557 VSUBS 0.012921f
C598 B.n558 VSUBS 0.012921f
C599 B.n559 VSUBS 0.012921f
C600 B.n560 VSUBS 0.012921f
C601 B.n561 VSUBS 0.012921f
C602 B.n562 VSUBS 0.012921f
C603 B.n563 VSUBS 0.012921f
C604 B.n564 VSUBS 0.012921f
C605 B.n565 VSUBS 0.012921f
C606 B.n566 VSUBS 0.012921f
C607 B.n567 VSUBS 0.012921f
C608 B.n568 VSUBS 0.012921f
C609 B.n569 VSUBS 0.012921f
C610 B.n570 VSUBS 0.012921f
C611 B.n571 VSUBS 0.012921f
C612 B.n572 VSUBS 0.012921f
C613 B.n573 VSUBS 0.012921f
C614 B.n574 VSUBS 0.012921f
C615 B.n575 VSUBS 0.012921f
C616 B.n576 VSUBS 0.012921f
C617 B.n577 VSUBS 0.012921f
C618 B.n578 VSUBS 0.012921f
C619 B.n579 VSUBS 0.012921f
C620 B.n580 VSUBS 0.012921f
C621 B.n581 VSUBS 0.012921f
C622 B.n582 VSUBS 0.012921f
C623 B.n583 VSUBS 0.012921f
C624 B.n584 VSUBS 0.012921f
C625 B.n585 VSUBS 0.012921f
C626 B.n586 VSUBS 0.012921f
C627 B.n587 VSUBS 0.012921f
C628 B.n588 VSUBS 0.012921f
C629 B.n589 VSUBS 0.012921f
C630 B.n590 VSUBS 0.012921f
C631 B.n591 VSUBS 0.012921f
C632 B.n592 VSUBS 0.012921f
C633 B.n593 VSUBS 0.012921f
C634 B.n594 VSUBS 0.012921f
C635 B.n595 VSUBS 0.012921f
C636 B.n596 VSUBS 0.012921f
C637 B.n597 VSUBS 0.012921f
C638 B.n598 VSUBS 0.012921f
C639 B.n599 VSUBS 0.012921f
C640 B.n600 VSUBS 0.012921f
C641 B.n601 VSUBS 0.012921f
C642 B.n602 VSUBS 0.012921f
C643 B.n603 VSUBS 0.012921f
C644 B.n604 VSUBS 0.012921f
C645 B.n605 VSUBS 0.012921f
C646 B.n606 VSUBS 0.012921f
C647 B.n607 VSUBS 0.012921f
C648 B.n608 VSUBS 0.012921f
C649 B.n609 VSUBS 0.012921f
C650 B.n610 VSUBS 0.012921f
C651 B.n611 VSUBS 0.012921f
C652 B.n612 VSUBS 0.012921f
C653 B.n613 VSUBS 0.012921f
C654 B.n614 VSUBS 0.012921f
C655 B.n615 VSUBS 0.012921f
C656 B.n616 VSUBS 0.012921f
C657 B.n617 VSUBS 0.012921f
C658 B.n618 VSUBS 0.012921f
C659 B.n619 VSUBS 0.012921f
C660 B.n620 VSUBS 0.012921f
C661 B.n621 VSUBS 0.012921f
C662 B.n622 VSUBS 0.012921f
C663 B.n623 VSUBS 0.012921f
C664 B.n624 VSUBS 0.012921f
C665 B.n625 VSUBS 0.012921f
C666 B.n626 VSUBS 0.012921f
C667 B.n627 VSUBS 0.012921f
C668 B.n628 VSUBS 0.012921f
C669 B.n629 VSUBS 0.012921f
C670 B.n630 VSUBS 0.012921f
C671 B.n631 VSUBS 0.012921f
C672 B.n632 VSUBS 0.012921f
C673 B.n633 VSUBS 0.012921f
C674 B.n634 VSUBS 0.012921f
C675 B.n635 VSUBS 0.029258f
C676 VDD1.t7 VSUBS 0.019536f
C677 VDD1.t3 VSUBS 0.019536f
C678 VDD1.n0 VSUBS 0.054519f
C679 VDD1.t4 VSUBS 0.019536f
C680 VDD1.t2 VSUBS 0.019536f
C681 VDD1.n1 VSUBS 0.054379f
C682 VDD1.t6 VSUBS 0.019536f
C683 VDD1.t0 VSUBS 0.019536f
C684 VDD1.n2 VSUBS 0.054379f
C685 VDD1.n3 VSUBS 3.44567f
C686 VDD1.t1 VSUBS 0.019536f
C687 VDD1.t5 VSUBS 0.019536f
C688 VDD1.n4 VSUBS 0.052785f
C689 VDD1.n5 VSUBS 2.63963f
C690 VP.t7 VSUBS 0.376449f
C691 VP.n0 VSUBS 0.520715f
C692 VP.n1 VSUBS 0.068314f
C693 VP.n2 VSUBS 0.089854f
C694 VP.n3 VSUBS 0.068314f
C695 VP.n4 VSUBS 0.07665f
C696 VP.n5 VSUBS 0.068314f
C697 VP.n6 VSUBS 0.055175f
C698 VP.n7 VSUBS 0.068314f
C699 VP.t5 VSUBS 0.376449f
C700 VP.n8 VSUBS 0.261836f
C701 VP.n9 VSUBS 0.068314f
C702 VP.n10 VSUBS 0.108755f
C703 VP.n11 VSUBS 0.068314f
C704 VP.n12 VSUBS 0.089158f
C705 VP.t2 VSUBS 0.376449f
C706 VP.n13 VSUBS 0.520715f
C707 VP.n14 VSUBS 0.068314f
C708 VP.n15 VSUBS 0.089854f
C709 VP.n16 VSUBS 0.068314f
C710 VP.n17 VSUBS 0.07665f
C711 VP.n18 VSUBS 0.068314f
C712 VP.n19 VSUBS 0.055175f
C713 VP.n20 VSUBS 0.068314f
C714 VP.t4 VSUBS 0.376449f
C715 VP.n21 VSUBS 0.51515f
C716 VP.t0 VSUBS 1.02309f
C717 VP.n22 VSUBS 0.628309f
C718 VP.n23 VSUBS 0.841374f
C719 VP.n24 VSUBS 0.114174f
C720 VP.n25 VSUBS 0.126682f
C721 VP.n26 VSUBS 0.135058f
C722 VP.n27 VSUBS 0.068314f
C723 VP.n28 VSUBS 0.068314f
C724 VP.n29 VSUBS 0.068314f
C725 VP.n30 VSUBS 0.135058f
C726 VP.n31 VSUBS 0.126682f
C727 VP.t6 VSUBS 0.376449f
C728 VP.n32 VSUBS 0.261836f
C729 VP.n33 VSUBS 0.114174f
C730 VP.n34 VSUBS 0.068314f
C731 VP.n35 VSUBS 0.068314f
C732 VP.n36 VSUBS 0.068314f
C733 VP.n37 VSUBS 0.126682f
C734 VP.n38 VSUBS 0.126682f
C735 VP.n39 VSUBS 0.108755f
C736 VP.n40 VSUBS 0.068314f
C737 VP.n41 VSUBS 0.068314f
C738 VP.n42 VSUBS 0.068314f
C739 VP.n43 VSUBS 0.126682f
C740 VP.n44 VSUBS 0.126682f
C741 VP.n45 VSUBS 0.089158f
C742 VP.n46 VSUBS 0.11024f
C743 VP.n47 VSUBS 3.52731f
C744 VP.t3 VSUBS 0.376449f
C745 VP.n48 VSUBS 0.520715f
C746 VP.n49 VSUBS 3.58012f
C747 VP.n50 VSUBS 0.11024f
C748 VP.n51 VSUBS 0.068314f
C749 VP.n52 VSUBS 0.126682f
C750 VP.n53 VSUBS 0.126682f
C751 VP.n54 VSUBS 0.089854f
C752 VP.n55 VSUBS 0.068314f
C753 VP.n56 VSUBS 0.068314f
C754 VP.n57 VSUBS 0.068314f
C755 VP.n58 VSUBS 0.126682f
C756 VP.n59 VSUBS 0.126682f
C757 VP.n60 VSUBS 0.07665f
C758 VP.n61 VSUBS 0.068314f
C759 VP.n62 VSUBS 0.068314f
C760 VP.n63 VSUBS 0.114174f
C761 VP.n64 VSUBS 0.126682f
C762 VP.n65 VSUBS 0.135058f
C763 VP.n66 VSUBS 0.068314f
C764 VP.n67 VSUBS 0.068314f
C765 VP.n68 VSUBS 0.068314f
C766 VP.n69 VSUBS 0.135058f
C767 VP.n70 VSUBS 0.126682f
C768 VP.t1 VSUBS 0.376449f
C769 VP.n71 VSUBS 0.261836f
C770 VP.n72 VSUBS 0.114174f
C771 VP.n73 VSUBS 0.068314f
C772 VP.n74 VSUBS 0.068314f
C773 VP.n75 VSUBS 0.068314f
C774 VP.n76 VSUBS 0.126682f
C775 VP.n77 VSUBS 0.126682f
C776 VP.n78 VSUBS 0.108755f
C777 VP.n79 VSUBS 0.068314f
C778 VP.n80 VSUBS 0.068314f
C779 VP.n81 VSUBS 0.068314f
C780 VP.n82 VSUBS 0.126682f
C781 VP.n83 VSUBS 0.126682f
C782 VP.n84 VSUBS 0.089158f
C783 VP.n85 VSUBS 0.11024f
C784 VP.n86 VSUBS 0.182804f
C785 VTAIL.t14 VSUBS 0.029117f
C786 VTAIL.t9 VSUBS 0.029117f
C787 VTAIL.n0 VSUBS 0.070763f
C788 VTAIL.n1 VSUBS 0.694644f
C789 VTAIL.t10 VSUBS 0.143525f
C790 VTAIL.n2 VSUBS 0.755595f
C791 VTAIL.t1 VSUBS 0.143525f
C792 VTAIL.n3 VSUBS 0.755595f
C793 VTAIL.t3 VSUBS 0.029117f
C794 VTAIL.t6 VSUBS 0.029117f
C795 VTAIL.n4 VSUBS 0.070763f
C796 VTAIL.n5 VSUBS 1.11912f
C797 VTAIL.t0 VSUBS 0.143525f
C798 VTAIL.n6 VSUBS 1.78424f
C799 VTAIL.t8 VSUBS 0.143525f
C800 VTAIL.n7 VSUBS 1.78424f
C801 VTAIL.t11 VSUBS 0.029117f
C802 VTAIL.t15 VSUBS 0.029117f
C803 VTAIL.n8 VSUBS 0.070763f
C804 VTAIL.n9 VSUBS 1.11912f
C805 VTAIL.t13 VSUBS 0.143525f
C806 VTAIL.n10 VSUBS 0.755595f
C807 VTAIL.t4 VSUBS 0.143525f
C808 VTAIL.n11 VSUBS 0.755595f
C809 VTAIL.t2 VSUBS 0.029117f
C810 VTAIL.t7 VSUBS 0.029117f
C811 VTAIL.n12 VSUBS 0.070763f
C812 VTAIL.n13 VSUBS 1.11912f
C813 VTAIL.t5 VSUBS 0.143525f
C814 VTAIL.n14 VSUBS 1.78424f
C815 VTAIL.t12 VSUBS 0.143525f
C816 VTAIL.n15 VSUBS 1.77657f
C817 VDD2.t4 VSUBS 0.025696f
C818 VDD2.t7 VSUBS 0.025696f
C819 VDD2.n0 VSUBS 0.071526f
C820 VDD2.t5 VSUBS 0.025696f
C821 VDD2.t1 VSUBS 0.025696f
C822 VDD2.n1 VSUBS 0.071526f
C823 VDD2.n2 VSUBS 4.45732f
C824 VDD2.t0 VSUBS 0.025696f
C825 VDD2.t2 VSUBS 0.025696f
C826 VDD2.n3 VSUBS 0.06943f
C827 VDD2.n4 VSUBS 3.42697f
C828 VDD2.t6 VSUBS 0.025696f
C829 VDD2.t3 VSUBS 0.025696f
C830 VDD2.n5 VSUBS 0.071521f
C831 VN.t3 VSUBS 0.32609f
C832 VN.n0 VSUBS 0.451056f
C833 VN.n1 VSUBS 0.059175f
C834 VN.n2 VSUBS 0.077834f
C835 VN.n3 VSUBS 0.059175f
C836 VN.n4 VSUBS 0.066396f
C837 VN.n5 VSUBS 0.059175f
C838 VN.n6 VSUBS 0.047794f
C839 VN.n7 VSUBS 0.059175f
C840 VN.t1 VSUBS 0.32609f
C841 VN.n8 VSUBS 0.446236f
C842 VN.t5 VSUBS 0.886227f
C843 VN.n9 VSUBS 0.544256f
C844 VN.n10 VSUBS 0.728818f
C845 VN.n11 VSUBS 0.0989f
C846 VN.n12 VSUBS 0.109735f
C847 VN.n13 VSUBS 0.116991f
C848 VN.n14 VSUBS 0.059175f
C849 VN.n15 VSUBS 0.059175f
C850 VN.n16 VSUBS 0.059175f
C851 VN.n17 VSUBS 0.116991f
C852 VN.n18 VSUBS 0.109735f
C853 VN.t6 VSUBS 0.32609f
C854 VN.n19 VSUBS 0.226809f
C855 VN.n20 VSUBS 0.0989f
C856 VN.n21 VSUBS 0.059175f
C857 VN.n22 VSUBS 0.059175f
C858 VN.n23 VSUBS 0.059175f
C859 VN.n24 VSUBS 0.109735f
C860 VN.n25 VSUBS 0.109735f
C861 VN.n26 VSUBS 0.094206f
C862 VN.n27 VSUBS 0.059175f
C863 VN.n28 VSUBS 0.059175f
C864 VN.n29 VSUBS 0.059175f
C865 VN.n30 VSUBS 0.109735f
C866 VN.n31 VSUBS 0.109735f
C867 VN.n32 VSUBS 0.077231f
C868 VN.n33 VSUBS 0.095492f
C869 VN.n34 VSUBS 0.158349f
C870 VN.t7 VSUBS 0.32609f
C871 VN.n35 VSUBS 0.451056f
C872 VN.n36 VSUBS 0.059175f
C873 VN.n37 VSUBS 0.077834f
C874 VN.n38 VSUBS 0.059175f
C875 VN.n39 VSUBS 0.066396f
C876 VN.n40 VSUBS 0.059175f
C877 VN.t4 VSUBS 0.32609f
C878 VN.n41 VSUBS 0.226809f
C879 VN.n42 VSUBS 0.047794f
C880 VN.n43 VSUBS 0.059175f
C881 VN.t0 VSUBS 0.32609f
C882 VN.n44 VSUBS 0.446236f
C883 VN.t2 VSUBS 0.886227f
C884 VN.n45 VSUBS 0.544256f
C885 VN.n46 VSUBS 0.728818f
C886 VN.n47 VSUBS 0.0989f
C887 VN.n48 VSUBS 0.109735f
C888 VN.n49 VSUBS 0.116991f
C889 VN.n50 VSUBS 0.059175f
C890 VN.n51 VSUBS 0.059175f
C891 VN.n52 VSUBS 0.059175f
C892 VN.n53 VSUBS 0.116991f
C893 VN.n54 VSUBS 0.109735f
C894 VN.n55 VSUBS 0.0989f
C895 VN.n56 VSUBS 0.059175f
C896 VN.n57 VSUBS 0.059175f
C897 VN.n58 VSUBS 0.059175f
C898 VN.n59 VSUBS 0.109735f
C899 VN.n60 VSUBS 0.109735f
C900 VN.n61 VSUBS 0.094206f
C901 VN.n62 VSUBS 0.059175f
C902 VN.n63 VSUBS 0.059175f
C903 VN.n64 VSUBS 0.059175f
C904 VN.n65 VSUBS 0.109735f
C905 VN.n66 VSUBS 0.109735f
C906 VN.n67 VSUBS 0.077231f
C907 VN.n68 VSUBS 0.095492f
C908 VN.n69 VSUBS 3.08025f
.ends

