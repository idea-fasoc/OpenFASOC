* NGSPICE file created from diff_pair_sample_1644.ext - technology: sky130A

.subckt diff_pair_sample_1644 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t1 VP.t0 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=2.7573 pd=14.92 as=2.7573 ps=14.92 w=7.07 l=3.6
X1 B.t15 B.t13 B.t14 B.t7 sky130_fd_pr__nfet_01v8 ad=2.7573 pd=14.92 as=0 ps=0 w=7.07 l=3.6
X2 VDD2.t1 VN.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.7573 pd=14.92 as=2.7573 ps=14.92 w=7.07 l=3.6
X3 B.t12 B.t10 B.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=2.7573 pd=14.92 as=0 ps=0 w=7.07 l=3.6
X4 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=2.7573 pd=14.92 as=0 ps=0 w=7.07 l=3.6
X5 VDD2.t0 VN.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.7573 pd=14.92 as=2.7573 ps=14.92 w=7.07 l=3.6
X6 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=2.7573 pd=14.92 as=0 ps=0 w=7.07 l=3.6
X7 VDD1.t0 VP.t1 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=2.7573 pd=14.92 as=2.7573 ps=14.92 w=7.07 l=3.6
R0 VP.n0 VP.t1 129.691
R1 VP.n0 VP.t0 86.118
R2 VP VP.n0 0.52637
R3 VTAIL.n1 VTAIL.t1 51.5391
R4 VTAIL.n3 VTAIL.t0 51.5389
R5 VTAIL.n0 VTAIL.t3 51.5389
R6 VTAIL.n2 VTAIL.t2 51.5389
R7 VTAIL.n1 VTAIL.n0 25.2376
R8 VTAIL.n3 VTAIL.n2 21.8496
R9 VTAIL.n2 VTAIL.n1 2.16429
R10 VTAIL VTAIL.n0 1.3755
R11 VTAIL VTAIL.n3 0.789293
R12 VDD1 VDD1.t1 106.12
R13 VDD1 VDD1.t0 69.1228
R14 B.n578 B.n577 585
R15 B.n219 B.n91 585
R16 B.n218 B.n217 585
R17 B.n216 B.n215 585
R18 B.n214 B.n213 585
R19 B.n212 B.n211 585
R20 B.n210 B.n209 585
R21 B.n208 B.n207 585
R22 B.n206 B.n205 585
R23 B.n204 B.n203 585
R24 B.n202 B.n201 585
R25 B.n200 B.n199 585
R26 B.n198 B.n197 585
R27 B.n196 B.n195 585
R28 B.n194 B.n193 585
R29 B.n192 B.n191 585
R30 B.n190 B.n189 585
R31 B.n188 B.n187 585
R32 B.n186 B.n185 585
R33 B.n184 B.n183 585
R34 B.n182 B.n181 585
R35 B.n180 B.n179 585
R36 B.n178 B.n177 585
R37 B.n176 B.n175 585
R38 B.n174 B.n173 585
R39 B.n172 B.n171 585
R40 B.n170 B.n169 585
R41 B.n167 B.n166 585
R42 B.n165 B.n164 585
R43 B.n163 B.n162 585
R44 B.n161 B.n160 585
R45 B.n159 B.n158 585
R46 B.n157 B.n156 585
R47 B.n155 B.n154 585
R48 B.n153 B.n152 585
R49 B.n151 B.n150 585
R50 B.n149 B.n148 585
R51 B.n146 B.n145 585
R52 B.n144 B.n143 585
R53 B.n142 B.n141 585
R54 B.n140 B.n139 585
R55 B.n138 B.n137 585
R56 B.n136 B.n135 585
R57 B.n134 B.n133 585
R58 B.n132 B.n131 585
R59 B.n130 B.n129 585
R60 B.n128 B.n127 585
R61 B.n126 B.n125 585
R62 B.n124 B.n123 585
R63 B.n122 B.n121 585
R64 B.n120 B.n119 585
R65 B.n118 B.n117 585
R66 B.n116 B.n115 585
R67 B.n114 B.n113 585
R68 B.n112 B.n111 585
R69 B.n110 B.n109 585
R70 B.n108 B.n107 585
R71 B.n106 B.n105 585
R72 B.n104 B.n103 585
R73 B.n102 B.n101 585
R74 B.n100 B.n99 585
R75 B.n98 B.n97 585
R76 B.n60 B.n59 585
R77 B.n583 B.n582 585
R78 B.n576 B.n92 585
R79 B.n92 B.n57 585
R80 B.n575 B.n56 585
R81 B.n587 B.n56 585
R82 B.n574 B.n55 585
R83 B.n588 B.n55 585
R84 B.n573 B.n54 585
R85 B.n589 B.n54 585
R86 B.n572 B.n571 585
R87 B.n571 B.n50 585
R88 B.n570 B.n49 585
R89 B.n595 B.n49 585
R90 B.n569 B.n48 585
R91 B.n596 B.n48 585
R92 B.n568 B.n47 585
R93 B.n597 B.n47 585
R94 B.n567 B.n566 585
R95 B.n566 B.n46 585
R96 B.n565 B.n42 585
R97 B.n603 B.n42 585
R98 B.n564 B.n41 585
R99 B.n604 B.n41 585
R100 B.n563 B.n40 585
R101 B.n605 B.n40 585
R102 B.n562 B.n561 585
R103 B.n561 B.n36 585
R104 B.n560 B.n35 585
R105 B.n611 B.n35 585
R106 B.n559 B.n34 585
R107 B.n612 B.n34 585
R108 B.n558 B.n33 585
R109 B.n613 B.n33 585
R110 B.n557 B.n556 585
R111 B.n556 B.n29 585
R112 B.n555 B.n28 585
R113 B.n619 B.n28 585
R114 B.n554 B.n27 585
R115 B.n620 B.n27 585
R116 B.n553 B.n26 585
R117 B.n621 B.n26 585
R118 B.n552 B.n551 585
R119 B.n551 B.n22 585
R120 B.n550 B.n21 585
R121 B.n627 B.n21 585
R122 B.n549 B.n20 585
R123 B.n628 B.n20 585
R124 B.n548 B.n19 585
R125 B.n629 B.n19 585
R126 B.n547 B.n546 585
R127 B.n546 B.n15 585
R128 B.n545 B.n14 585
R129 B.n635 B.n14 585
R130 B.n544 B.n13 585
R131 B.n636 B.n13 585
R132 B.n543 B.n12 585
R133 B.n637 B.n12 585
R134 B.n542 B.n541 585
R135 B.n541 B.n8 585
R136 B.n540 B.n7 585
R137 B.n643 B.n7 585
R138 B.n539 B.n6 585
R139 B.n644 B.n6 585
R140 B.n538 B.n5 585
R141 B.n645 B.n5 585
R142 B.n537 B.n536 585
R143 B.n536 B.n4 585
R144 B.n535 B.n220 585
R145 B.n535 B.n534 585
R146 B.n525 B.n221 585
R147 B.n222 B.n221 585
R148 B.n527 B.n526 585
R149 B.n528 B.n527 585
R150 B.n524 B.n227 585
R151 B.n227 B.n226 585
R152 B.n523 B.n522 585
R153 B.n522 B.n521 585
R154 B.n229 B.n228 585
R155 B.n230 B.n229 585
R156 B.n514 B.n513 585
R157 B.n515 B.n514 585
R158 B.n512 B.n235 585
R159 B.n235 B.n234 585
R160 B.n511 B.n510 585
R161 B.n510 B.n509 585
R162 B.n237 B.n236 585
R163 B.n238 B.n237 585
R164 B.n502 B.n501 585
R165 B.n503 B.n502 585
R166 B.n500 B.n243 585
R167 B.n243 B.n242 585
R168 B.n499 B.n498 585
R169 B.n498 B.n497 585
R170 B.n245 B.n244 585
R171 B.n246 B.n245 585
R172 B.n490 B.n489 585
R173 B.n491 B.n490 585
R174 B.n488 B.n251 585
R175 B.n251 B.n250 585
R176 B.n487 B.n486 585
R177 B.n486 B.n485 585
R178 B.n253 B.n252 585
R179 B.n254 B.n253 585
R180 B.n478 B.n477 585
R181 B.n479 B.n478 585
R182 B.n476 B.n259 585
R183 B.n259 B.n258 585
R184 B.n475 B.n474 585
R185 B.n474 B.n473 585
R186 B.n261 B.n260 585
R187 B.n466 B.n261 585
R188 B.n465 B.n464 585
R189 B.n467 B.n465 585
R190 B.n463 B.n266 585
R191 B.n266 B.n265 585
R192 B.n462 B.n461 585
R193 B.n461 B.n460 585
R194 B.n268 B.n267 585
R195 B.n269 B.n268 585
R196 B.n453 B.n452 585
R197 B.n454 B.n453 585
R198 B.n451 B.n274 585
R199 B.n274 B.n273 585
R200 B.n450 B.n449 585
R201 B.n449 B.n448 585
R202 B.n276 B.n275 585
R203 B.n277 B.n276 585
R204 B.n444 B.n443 585
R205 B.n280 B.n279 585
R206 B.n440 B.n439 585
R207 B.n441 B.n440 585
R208 B.n438 B.n312 585
R209 B.n437 B.n436 585
R210 B.n435 B.n434 585
R211 B.n433 B.n432 585
R212 B.n431 B.n430 585
R213 B.n429 B.n428 585
R214 B.n427 B.n426 585
R215 B.n425 B.n424 585
R216 B.n423 B.n422 585
R217 B.n421 B.n420 585
R218 B.n419 B.n418 585
R219 B.n417 B.n416 585
R220 B.n415 B.n414 585
R221 B.n413 B.n412 585
R222 B.n411 B.n410 585
R223 B.n409 B.n408 585
R224 B.n407 B.n406 585
R225 B.n405 B.n404 585
R226 B.n403 B.n402 585
R227 B.n401 B.n400 585
R228 B.n399 B.n398 585
R229 B.n397 B.n396 585
R230 B.n395 B.n394 585
R231 B.n393 B.n392 585
R232 B.n391 B.n390 585
R233 B.n389 B.n388 585
R234 B.n387 B.n386 585
R235 B.n385 B.n384 585
R236 B.n383 B.n382 585
R237 B.n381 B.n380 585
R238 B.n379 B.n378 585
R239 B.n377 B.n376 585
R240 B.n375 B.n374 585
R241 B.n373 B.n372 585
R242 B.n371 B.n370 585
R243 B.n369 B.n368 585
R244 B.n367 B.n366 585
R245 B.n365 B.n364 585
R246 B.n363 B.n362 585
R247 B.n361 B.n360 585
R248 B.n359 B.n358 585
R249 B.n357 B.n356 585
R250 B.n355 B.n354 585
R251 B.n353 B.n352 585
R252 B.n351 B.n350 585
R253 B.n349 B.n348 585
R254 B.n347 B.n346 585
R255 B.n345 B.n344 585
R256 B.n343 B.n342 585
R257 B.n341 B.n340 585
R258 B.n339 B.n338 585
R259 B.n337 B.n336 585
R260 B.n335 B.n334 585
R261 B.n333 B.n332 585
R262 B.n331 B.n330 585
R263 B.n329 B.n328 585
R264 B.n327 B.n326 585
R265 B.n325 B.n324 585
R266 B.n323 B.n322 585
R267 B.n321 B.n320 585
R268 B.n319 B.n311 585
R269 B.n441 B.n311 585
R270 B.n445 B.n278 585
R271 B.n278 B.n277 585
R272 B.n447 B.n446 585
R273 B.n448 B.n447 585
R274 B.n272 B.n271 585
R275 B.n273 B.n272 585
R276 B.n456 B.n455 585
R277 B.n455 B.n454 585
R278 B.n457 B.n270 585
R279 B.n270 B.n269 585
R280 B.n459 B.n458 585
R281 B.n460 B.n459 585
R282 B.n264 B.n263 585
R283 B.n265 B.n264 585
R284 B.n469 B.n468 585
R285 B.n468 B.n467 585
R286 B.n470 B.n262 585
R287 B.n466 B.n262 585
R288 B.n472 B.n471 585
R289 B.n473 B.n472 585
R290 B.n257 B.n256 585
R291 B.n258 B.n257 585
R292 B.n481 B.n480 585
R293 B.n480 B.n479 585
R294 B.n482 B.n255 585
R295 B.n255 B.n254 585
R296 B.n484 B.n483 585
R297 B.n485 B.n484 585
R298 B.n249 B.n248 585
R299 B.n250 B.n249 585
R300 B.n493 B.n492 585
R301 B.n492 B.n491 585
R302 B.n494 B.n247 585
R303 B.n247 B.n246 585
R304 B.n496 B.n495 585
R305 B.n497 B.n496 585
R306 B.n241 B.n240 585
R307 B.n242 B.n241 585
R308 B.n505 B.n504 585
R309 B.n504 B.n503 585
R310 B.n506 B.n239 585
R311 B.n239 B.n238 585
R312 B.n508 B.n507 585
R313 B.n509 B.n508 585
R314 B.n233 B.n232 585
R315 B.n234 B.n233 585
R316 B.n517 B.n516 585
R317 B.n516 B.n515 585
R318 B.n518 B.n231 585
R319 B.n231 B.n230 585
R320 B.n520 B.n519 585
R321 B.n521 B.n520 585
R322 B.n225 B.n224 585
R323 B.n226 B.n225 585
R324 B.n530 B.n529 585
R325 B.n529 B.n528 585
R326 B.n531 B.n223 585
R327 B.n223 B.n222 585
R328 B.n533 B.n532 585
R329 B.n534 B.n533 585
R330 B.n2 B.n0 585
R331 B.n4 B.n2 585
R332 B.n3 B.n1 585
R333 B.n644 B.n3 585
R334 B.n642 B.n641 585
R335 B.n643 B.n642 585
R336 B.n640 B.n9 585
R337 B.n9 B.n8 585
R338 B.n639 B.n638 585
R339 B.n638 B.n637 585
R340 B.n11 B.n10 585
R341 B.n636 B.n11 585
R342 B.n634 B.n633 585
R343 B.n635 B.n634 585
R344 B.n632 B.n16 585
R345 B.n16 B.n15 585
R346 B.n631 B.n630 585
R347 B.n630 B.n629 585
R348 B.n18 B.n17 585
R349 B.n628 B.n18 585
R350 B.n626 B.n625 585
R351 B.n627 B.n626 585
R352 B.n624 B.n23 585
R353 B.n23 B.n22 585
R354 B.n623 B.n622 585
R355 B.n622 B.n621 585
R356 B.n25 B.n24 585
R357 B.n620 B.n25 585
R358 B.n618 B.n617 585
R359 B.n619 B.n618 585
R360 B.n616 B.n30 585
R361 B.n30 B.n29 585
R362 B.n615 B.n614 585
R363 B.n614 B.n613 585
R364 B.n32 B.n31 585
R365 B.n612 B.n32 585
R366 B.n610 B.n609 585
R367 B.n611 B.n610 585
R368 B.n608 B.n37 585
R369 B.n37 B.n36 585
R370 B.n607 B.n606 585
R371 B.n606 B.n605 585
R372 B.n39 B.n38 585
R373 B.n604 B.n39 585
R374 B.n602 B.n601 585
R375 B.n603 B.n602 585
R376 B.n600 B.n43 585
R377 B.n46 B.n43 585
R378 B.n599 B.n598 585
R379 B.n598 B.n597 585
R380 B.n45 B.n44 585
R381 B.n596 B.n45 585
R382 B.n594 B.n593 585
R383 B.n595 B.n594 585
R384 B.n592 B.n51 585
R385 B.n51 B.n50 585
R386 B.n591 B.n590 585
R387 B.n590 B.n589 585
R388 B.n53 B.n52 585
R389 B.n588 B.n53 585
R390 B.n586 B.n585 585
R391 B.n587 B.n586 585
R392 B.n584 B.n58 585
R393 B.n58 B.n57 585
R394 B.n647 B.n646 585
R395 B.n646 B.n645 585
R396 B.n443 B.n278 521.33
R397 B.n582 B.n58 521.33
R398 B.n311 B.n276 521.33
R399 B.n578 B.n92 521.33
R400 B.n580 B.n579 256.663
R401 B.n580 B.n90 256.663
R402 B.n580 B.n89 256.663
R403 B.n580 B.n88 256.663
R404 B.n580 B.n87 256.663
R405 B.n580 B.n86 256.663
R406 B.n580 B.n85 256.663
R407 B.n580 B.n84 256.663
R408 B.n580 B.n83 256.663
R409 B.n580 B.n82 256.663
R410 B.n580 B.n81 256.663
R411 B.n580 B.n80 256.663
R412 B.n580 B.n79 256.663
R413 B.n580 B.n78 256.663
R414 B.n580 B.n77 256.663
R415 B.n580 B.n76 256.663
R416 B.n580 B.n75 256.663
R417 B.n580 B.n74 256.663
R418 B.n580 B.n73 256.663
R419 B.n580 B.n72 256.663
R420 B.n580 B.n71 256.663
R421 B.n580 B.n70 256.663
R422 B.n580 B.n69 256.663
R423 B.n580 B.n68 256.663
R424 B.n580 B.n67 256.663
R425 B.n580 B.n66 256.663
R426 B.n580 B.n65 256.663
R427 B.n580 B.n64 256.663
R428 B.n580 B.n63 256.663
R429 B.n580 B.n62 256.663
R430 B.n580 B.n61 256.663
R431 B.n581 B.n580 256.663
R432 B.n442 B.n441 256.663
R433 B.n441 B.n281 256.663
R434 B.n441 B.n282 256.663
R435 B.n441 B.n283 256.663
R436 B.n441 B.n284 256.663
R437 B.n441 B.n285 256.663
R438 B.n441 B.n286 256.663
R439 B.n441 B.n287 256.663
R440 B.n441 B.n288 256.663
R441 B.n441 B.n289 256.663
R442 B.n441 B.n290 256.663
R443 B.n441 B.n291 256.663
R444 B.n441 B.n292 256.663
R445 B.n441 B.n293 256.663
R446 B.n441 B.n294 256.663
R447 B.n441 B.n295 256.663
R448 B.n441 B.n296 256.663
R449 B.n441 B.n297 256.663
R450 B.n441 B.n298 256.663
R451 B.n441 B.n299 256.663
R452 B.n441 B.n300 256.663
R453 B.n441 B.n301 256.663
R454 B.n441 B.n302 256.663
R455 B.n441 B.n303 256.663
R456 B.n441 B.n304 256.663
R457 B.n441 B.n305 256.663
R458 B.n441 B.n306 256.663
R459 B.n441 B.n307 256.663
R460 B.n441 B.n308 256.663
R461 B.n441 B.n309 256.663
R462 B.n441 B.n310 256.663
R463 B.n316 B.t2 256.512
R464 B.n313 B.t10 256.512
R465 B.n95 B.t6 256.512
R466 B.n93 B.t13 256.512
R467 B.n447 B.n278 163.367
R468 B.n447 B.n272 163.367
R469 B.n455 B.n272 163.367
R470 B.n455 B.n270 163.367
R471 B.n459 B.n270 163.367
R472 B.n459 B.n264 163.367
R473 B.n468 B.n264 163.367
R474 B.n468 B.n262 163.367
R475 B.n472 B.n262 163.367
R476 B.n472 B.n257 163.367
R477 B.n480 B.n257 163.367
R478 B.n480 B.n255 163.367
R479 B.n484 B.n255 163.367
R480 B.n484 B.n249 163.367
R481 B.n492 B.n249 163.367
R482 B.n492 B.n247 163.367
R483 B.n496 B.n247 163.367
R484 B.n496 B.n241 163.367
R485 B.n504 B.n241 163.367
R486 B.n504 B.n239 163.367
R487 B.n508 B.n239 163.367
R488 B.n508 B.n233 163.367
R489 B.n516 B.n233 163.367
R490 B.n516 B.n231 163.367
R491 B.n520 B.n231 163.367
R492 B.n520 B.n225 163.367
R493 B.n529 B.n225 163.367
R494 B.n529 B.n223 163.367
R495 B.n533 B.n223 163.367
R496 B.n533 B.n2 163.367
R497 B.n646 B.n2 163.367
R498 B.n646 B.n3 163.367
R499 B.n642 B.n3 163.367
R500 B.n642 B.n9 163.367
R501 B.n638 B.n9 163.367
R502 B.n638 B.n11 163.367
R503 B.n634 B.n11 163.367
R504 B.n634 B.n16 163.367
R505 B.n630 B.n16 163.367
R506 B.n630 B.n18 163.367
R507 B.n626 B.n18 163.367
R508 B.n626 B.n23 163.367
R509 B.n622 B.n23 163.367
R510 B.n622 B.n25 163.367
R511 B.n618 B.n25 163.367
R512 B.n618 B.n30 163.367
R513 B.n614 B.n30 163.367
R514 B.n614 B.n32 163.367
R515 B.n610 B.n32 163.367
R516 B.n610 B.n37 163.367
R517 B.n606 B.n37 163.367
R518 B.n606 B.n39 163.367
R519 B.n602 B.n39 163.367
R520 B.n602 B.n43 163.367
R521 B.n598 B.n43 163.367
R522 B.n598 B.n45 163.367
R523 B.n594 B.n45 163.367
R524 B.n594 B.n51 163.367
R525 B.n590 B.n51 163.367
R526 B.n590 B.n53 163.367
R527 B.n586 B.n53 163.367
R528 B.n586 B.n58 163.367
R529 B.n440 B.n280 163.367
R530 B.n440 B.n312 163.367
R531 B.n436 B.n435 163.367
R532 B.n432 B.n431 163.367
R533 B.n428 B.n427 163.367
R534 B.n424 B.n423 163.367
R535 B.n420 B.n419 163.367
R536 B.n416 B.n415 163.367
R537 B.n412 B.n411 163.367
R538 B.n408 B.n407 163.367
R539 B.n404 B.n403 163.367
R540 B.n400 B.n399 163.367
R541 B.n396 B.n395 163.367
R542 B.n392 B.n391 163.367
R543 B.n388 B.n387 163.367
R544 B.n384 B.n383 163.367
R545 B.n380 B.n379 163.367
R546 B.n376 B.n375 163.367
R547 B.n372 B.n371 163.367
R548 B.n368 B.n367 163.367
R549 B.n364 B.n363 163.367
R550 B.n360 B.n359 163.367
R551 B.n356 B.n355 163.367
R552 B.n352 B.n351 163.367
R553 B.n348 B.n347 163.367
R554 B.n344 B.n343 163.367
R555 B.n340 B.n339 163.367
R556 B.n336 B.n335 163.367
R557 B.n332 B.n331 163.367
R558 B.n328 B.n327 163.367
R559 B.n324 B.n323 163.367
R560 B.n320 B.n311 163.367
R561 B.n449 B.n276 163.367
R562 B.n449 B.n274 163.367
R563 B.n453 B.n274 163.367
R564 B.n453 B.n268 163.367
R565 B.n461 B.n268 163.367
R566 B.n461 B.n266 163.367
R567 B.n465 B.n266 163.367
R568 B.n465 B.n261 163.367
R569 B.n474 B.n261 163.367
R570 B.n474 B.n259 163.367
R571 B.n478 B.n259 163.367
R572 B.n478 B.n253 163.367
R573 B.n486 B.n253 163.367
R574 B.n486 B.n251 163.367
R575 B.n490 B.n251 163.367
R576 B.n490 B.n245 163.367
R577 B.n498 B.n245 163.367
R578 B.n498 B.n243 163.367
R579 B.n502 B.n243 163.367
R580 B.n502 B.n237 163.367
R581 B.n510 B.n237 163.367
R582 B.n510 B.n235 163.367
R583 B.n514 B.n235 163.367
R584 B.n514 B.n229 163.367
R585 B.n522 B.n229 163.367
R586 B.n522 B.n227 163.367
R587 B.n527 B.n227 163.367
R588 B.n527 B.n221 163.367
R589 B.n535 B.n221 163.367
R590 B.n536 B.n535 163.367
R591 B.n536 B.n5 163.367
R592 B.n6 B.n5 163.367
R593 B.n7 B.n6 163.367
R594 B.n541 B.n7 163.367
R595 B.n541 B.n12 163.367
R596 B.n13 B.n12 163.367
R597 B.n14 B.n13 163.367
R598 B.n546 B.n14 163.367
R599 B.n546 B.n19 163.367
R600 B.n20 B.n19 163.367
R601 B.n21 B.n20 163.367
R602 B.n551 B.n21 163.367
R603 B.n551 B.n26 163.367
R604 B.n27 B.n26 163.367
R605 B.n28 B.n27 163.367
R606 B.n556 B.n28 163.367
R607 B.n556 B.n33 163.367
R608 B.n34 B.n33 163.367
R609 B.n35 B.n34 163.367
R610 B.n561 B.n35 163.367
R611 B.n561 B.n40 163.367
R612 B.n41 B.n40 163.367
R613 B.n42 B.n41 163.367
R614 B.n566 B.n42 163.367
R615 B.n566 B.n47 163.367
R616 B.n48 B.n47 163.367
R617 B.n49 B.n48 163.367
R618 B.n571 B.n49 163.367
R619 B.n571 B.n54 163.367
R620 B.n55 B.n54 163.367
R621 B.n56 B.n55 163.367
R622 B.n92 B.n56 163.367
R623 B.n97 B.n60 163.367
R624 B.n101 B.n100 163.367
R625 B.n105 B.n104 163.367
R626 B.n109 B.n108 163.367
R627 B.n113 B.n112 163.367
R628 B.n117 B.n116 163.367
R629 B.n121 B.n120 163.367
R630 B.n125 B.n124 163.367
R631 B.n129 B.n128 163.367
R632 B.n133 B.n132 163.367
R633 B.n137 B.n136 163.367
R634 B.n141 B.n140 163.367
R635 B.n145 B.n144 163.367
R636 B.n150 B.n149 163.367
R637 B.n154 B.n153 163.367
R638 B.n158 B.n157 163.367
R639 B.n162 B.n161 163.367
R640 B.n166 B.n165 163.367
R641 B.n171 B.n170 163.367
R642 B.n175 B.n174 163.367
R643 B.n179 B.n178 163.367
R644 B.n183 B.n182 163.367
R645 B.n187 B.n186 163.367
R646 B.n191 B.n190 163.367
R647 B.n195 B.n194 163.367
R648 B.n199 B.n198 163.367
R649 B.n203 B.n202 163.367
R650 B.n207 B.n206 163.367
R651 B.n211 B.n210 163.367
R652 B.n215 B.n214 163.367
R653 B.n217 B.n91 163.367
R654 B.n316 B.t5 150.392
R655 B.n93 B.t14 150.392
R656 B.n313 B.t12 150.383
R657 B.n95 B.t8 150.383
R658 B.n441 B.n277 123.856
R659 B.n580 B.n57 123.856
R660 B.n317 B.n316 76.2187
R661 B.n314 B.n313 76.2187
R662 B.n96 B.n95 76.2187
R663 B.n94 B.n93 76.2187
R664 B.n317 B.t4 74.1734
R665 B.n94 B.t15 74.1734
R666 B.n314 B.t11 74.1656
R667 B.n96 B.t9 74.1656
R668 B.n443 B.n442 71.676
R669 B.n312 B.n281 71.676
R670 B.n435 B.n282 71.676
R671 B.n431 B.n283 71.676
R672 B.n427 B.n284 71.676
R673 B.n423 B.n285 71.676
R674 B.n419 B.n286 71.676
R675 B.n415 B.n287 71.676
R676 B.n411 B.n288 71.676
R677 B.n407 B.n289 71.676
R678 B.n403 B.n290 71.676
R679 B.n399 B.n291 71.676
R680 B.n395 B.n292 71.676
R681 B.n391 B.n293 71.676
R682 B.n387 B.n294 71.676
R683 B.n383 B.n295 71.676
R684 B.n379 B.n296 71.676
R685 B.n375 B.n297 71.676
R686 B.n371 B.n298 71.676
R687 B.n367 B.n299 71.676
R688 B.n363 B.n300 71.676
R689 B.n359 B.n301 71.676
R690 B.n355 B.n302 71.676
R691 B.n351 B.n303 71.676
R692 B.n347 B.n304 71.676
R693 B.n343 B.n305 71.676
R694 B.n339 B.n306 71.676
R695 B.n335 B.n307 71.676
R696 B.n331 B.n308 71.676
R697 B.n327 B.n309 71.676
R698 B.n323 B.n310 71.676
R699 B.n582 B.n581 71.676
R700 B.n97 B.n61 71.676
R701 B.n101 B.n62 71.676
R702 B.n105 B.n63 71.676
R703 B.n109 B.n64 71.676
R704 B.n113 B.n65 71.676
R705 B.n117 B.n66 71.676
R706 B.n121 B.n67 71.676
R707 B.n125 B.n68 71.676
R708 B.n129 B.n69 71.676
R709 B.n133 B.n70 71.676
R710 B.n137 B.n71 71.676
R711 B.n141 B.n72 71.676
R712 B.n145 B.n73 71.676
R713 B.n150 B.n74 71.676
R714 B.n154 B.n75 71.676
R715 B.n158 B.n76 71.676
R716 B.n162 B.n77 71.676
R717 B.n166 B.n78 71.676
R718 B.n171 B.n79 71.676
R719 B.n175 B.n80 71.676
R720 B.n179 B.n81 71.676
R721 B.n183 B.n82 71.676
R722 B.n187 B.n83 71.676
R723 B.n191 B.n84 71.676
R724 B.n195 B.n85 71.676
R725 B.n199 B.n86 71.676
R726 B.n203 B.n87 71.676
R727 B.n207 B.n88 71.676
R728 B.n211 B.n89 71.676
R729 B.n215 B.n90 71.676
R730 B.n579 B.n91 71.676
R731 B.n579 B.n578 71.676
R732 B.n217 B.n90 71.676
R733 B.n214 B.n89 71.676
R734 B.n210 B.n88 71.676
R735 B.n206 B.n87 71.676
R736 B.n202 B.n86 71.676
R737 B.n198 B.n85 71.676
R738 B.n194 B.n84 71.676
R739 B.n190 B.n83 71.676
R740 B.n186 B.n82 71.676
R741 B.n182 B.n81 71.676
R742 B.n178 B.n80 71.676
R743 B.n174 B.n79 71.676
R744 B.n170 B.n78 71.676
R745 B.n165 B.n77 71.676
R746 B.n161 B.n76 71.676
R747 B.n157 B.n75 71.676
R748 B.n153 B.n74 71.676
R749 B.n149 B.n73 71.676
R750 B.n144 B.n72 71.676
R751 B.n140 B.n71 71.676
R752 B.n136 B.n70 71.676
R753 B.n132 B.n69 71.676
R754 B.n128 B.n68 71.676
R755 B.n124 B.n67 71.676
R756 B.n120 B.n66 71.676
R757 B.n116 B.n65 71.676
R758 B.n112 B.n64 71.676
R759 B.n108 B.n63 71.676
R760 B.n104 B.n62 71.676
R761 B.n100 B.n61 71.676
R762 B.n581 B.n60 71.676
R763 B.n442 B.n280 71.676
R764 B.n436 B.n281 71.676
R765 B.n432 B.n282 71.676
R766 B.n428 B.n283 71.676
R767 B.n424 B.n284 71.676
R768 B.n420 B.n285 71.676
R769 B.n416 B.n286 71.676
R770 B.n412 B.n287 71.676
R771 B.n408 B.n288 71.676
R772 B.n404 B.n289 71.676
R773 B.n400 B.n290 71.676
R774 B.n396 B.n291 71.676
R775 B.n392 B.n292 71.676
R776 B.n388 B.n293 71.676
R777 B.n384 B.n294 71.676
R778 B.n380 B.n295 71.676
R779 B.n376 B.n296 71.676
R780 B.n372 B.n297 71.676
R781 B.n368 B.n298 71.676
R782 B.n364 B.n299 71.676
R783 B.n360 B.n300 71.676
R784 B.n356 B.n301 71.676
R785 B.n352 B.n302 71.676
R786 B.n348 B.n303 71.676
R787 B.n344 B.n304 71.676
R788 B.n340 B.n305 71.676
R789 B.n336 B.n306 71.676
R790 B.n332 B.n307 71.676
R791 B.n328 B.n308 71.676
R792 B.n324 B.n309 71.676
R793 B.n320 B.n310 71.676
R794 B.n448 B.n277 60.5918
R795 B.n448 B.n273 60.5918
R796 B.n454 B.n273 60.5918
R797 B.n454 B.n269 60.5918
R798 B.n460 B.n269 60.5918
R799 B.n460 B.n265 60.5918
R800 B.n467 B.n265 60.5918
R801 B.n467 B.n466 60.5918
R802 B.n473 B.n258 60.5918
R803 B.n479 B.n258 60.5918
R804 B.n479 B.n254 60.5918
R805 B.n485 B.n254 60.5918
R806 B.n485 B.n250 60.5918
R807 B.n491 B.n250 60.5918
R808 B.n491 B.n246 60.5918
R809 B.n497 B.n246 60.5918
R810 B.n497 B.n242 60.5918
R811 B.n503 B.n242 60.5918
R812 B.n503 B.n238 60.5918
R813 B.n509 B.n238 60.5918
R814 B.n509 B.n234 60.5918
R815 B.n515 B.n234 60.5918
R816 B.n521 B.n230 60.5918
R817 B.n521 B.n226 60.5918
R818 B.n528 B.n226 60.5918
R819 B.n528 B.n222 60.5918
R820 B.n534 B.n222 60.5918
R821 B.n534 B.n4 60.5918
R822 B.n645 B.n4 60.5918
R823 B.n645 B.n644 60.5918
R824 B.n644 B.n643 60.5918
R825 B.n643 B.n8 60.5918
R826 B.n637 B.n8 60.5918
R827 B.n637 B.n636 60.5918
R828 B.n636 B.n635 60.5918
R829 B.n635 B.n15 60.5918
R830 B.n629 B.n628 60.5918
R831 B.n628 B.n627 60.5918
R832 B.n627 B.n22 60.5918
R833 B.n621 B.n22 60.5918
R834 B.n621 B.n620 60.5918
R835 B.n620 B.n619 60.5918
R836 B.n619 B.n29 60.5918
R837 B.n613 B.n29 60.5918
R838 B.n613 B.n612 60.5918
R839 B.n612 B.n611 60.5918
R840 B.n611 B.n36 60.5918
R841 B.n605 B.n36 60.5918
R842 B.n605 B.n604 60.5918
R843 B.n604 B.n603 60.5918
R844 B.n597 B.n46 60.5918
R845 B.n597 B.n596 60.5918
R846 B.n596 B.n595 60.5918
R847 B.n595 B.n50 60.5918
R848 B.n589 B.n50 60.5918
R849 B.n589 B.n588 60.5918
R850 B.n588 B.n587 60.5918
R851 B.n587 B.n57 60.5918
R852 B.n318 B.n317 59.5399
R853 B.n315 B.n314 59.5399
R854 B.n147 B.n96 59.5399
R855 B.n168 B.n94 59.5399
R856 B.n466 B.t3 51.6813
R857 B.n46 B.t7 51.6813
R858 B.n515 B.t1 37.4246
R859 B.n629 B.t0 37.4246
R860 B.n584 B.n583 33.8737
R861 B.n577 B.n576 33.8737
R862 B.n319 B.n275 33.8737
R863 B.n445 B.n444 33.8737
R864 B.t1 B.n230 23.1678
R865 B.t0 B.n15 23.1678
R866 B B.n647 18.0485
R867 B.n583 B.n59 10.6151
R868 B.n98 B.n59 10.6151
R869 B.n99 B.n98 10.6151
R870 B.n102 B.n99 10.6151
R871 B.n103 B.n102 10.6151
R872 B.n106 B.n103 10.6151
R873 B.n107 B.n106 10.6151
R874 B.n110 B.n107 10.6151
R875 B.n111 B.n110 10.6151
R876 B.n114 B.n111 10.6151
R877 B.n115 B.n114 10.6151
R878 B.n118 B.n115 10.6151
R879 B.n119 B.n118 10.6151
R880 B.n122 B.n119 10.6151
R881 B.n123 B.n122 10.6151
R882 B.n126 B.n123 10.6151
R883 B.n127 B.n126 10.6151
R884 B.n130 B.n127 10.6151
R885 B.n131 B.n130 10.6151
R886 B.n134 B.n131 10.6151
R887 B.n135 B.n134 10.6151
R888 B.n138 B.n135 10.6151
R889 B.n139 B.n138 10.6151
R890 B.n142 B.n139 10.6151
R891 B.n143 B.n142 10.6151
R892 B.n146 B.n143 10.6151
R893 B.n151 B.n148 10.6151
R894 B.n152 B.n151 10.6151
R895 B.n155 B.n152 10.6151
R896 B.n156 B.n155 10.6151
R897 B.n159 B.n156 10.6151
R898 B.n160 B.n159 10.6151
R899 B.n163 B.n160 10.6151
R900 B.n164 B.n163 10.6151
R901 B.n167 B.n164 10.6151
R902 B.n172 B.n169 10.6151
R903 B.n173 B.n172 10.6151
R904 B.n176 B.n173 10.6151
R905 B.n177 B.n176 10.6151
R906 B.n180 B.n177 10.6151
R907 B.n181 B.n180 10.6151
R908 B.n184 B.n181 10.6151
R909 B.n185 B.n184 10.6151
R910 B.n188 B.n185 10.6151
R911 B.n189 B.n188 10.6151
R912 B.n192 B.n189 10.6151
R913 B.n193 B.n192 10.6151
R914 B.n196 B.n193 10.6151
R915 B.n197 B.n196 10.6151
R916 B.n200 B.n197 10.6151
R917 B.n201 B.n200 10.6151
R918 B.n204 B.n201 10.6151
R919 B.n205 B.n204 10.6151
R920 B.n208 B.n205 10.6151
R921 B.n209 B.n208 10.6151
R922 B.n212 B.n209 10.6151
R923 B.n213 B.n212 10.6151
R924 B.n216 B.n213 10.6151
R925 B.n218 B.n216 10.6151
R926 B.n219 B.n218 10.6151
R927 B.n577 B.n219 10.6151
R928 B.n450 B.n275 10.6151
R929 B.n451 B.n450 10.6151
R930 B.n452 B.n451 10.6151
R931 B.n452 B.n267 10.6151
R932 B.n462 B.n267 10.6151
R933 B.n463 B.n462 10.6151
R934 B.n464 B.n463 10.6151
R935 B.n464 B.n260 10.6151
R936 B.n475 B.n260 10.6151
R937 B.n476 B.n475 10.6151
R938 B.n477 B.n476 10.6151
R939 B.n477 B.n252 10.6151
R940 B.n487 B.n252 10.6151
R941 B.n488 B.n487 10.6151
R942 B.n489 B.n488 10.6151
R943 B.n489 B.n244 10.6151
R944 B.n499 B.n244 10.6151
R945 B.n500 B.n499 10.6151
R946 B.n501 B.n500 10.6151
R947 B.n501 B.n236 10.6151
R948 B.n511 B.n236 10.6151
R949 B.n512 B.n511 10.6151
R950 B.n513 B.n512 10.6151
R951 B.n513 B.n228 10.6151
R952 B.n523 B.n228 10.6151
R953 B.n524 B.n523 10.6151
R954 B.n526 B.n524 10.6151
R955 B.n526 B.n525 10.6151
R956 B.n525 B.n220 10.6151
R957 B.n537 B.n220 10.6151
R958 B.n538 B.n537 10.6151
R959 B.n539 B.n538 10.6151
R960 B.n540 B.n539 10.6151
R961 B.n542 B.n540 10.6151
R962 B.n543 B.n542 10.6151
R963 B.n544 B.n543 10.6151
R964 B.n545 B.n544 10.6151
R965 B.n547 B.n545 10.6151
R966 B.n548 B.n547 10.6151
R967 B.n549 B.n548 10.6151
R968 B.n550 B.n549 10.6151
R969 B.n552 B.n550 10.6151
R970 B.n553 B.n552 10.6151
R971 B.n554 B.n553 10.6151
R972 B.n555 B.n554 10.6151
R973 B.n557 B.n555 10.6151
R974 B.n558 B.n557 10.6151
R975 B.n559 B.n558 10.6151
R976 B.n560 B.n559 10.6151
R977 B.n562 B.n560 10.6151
R978 B.n563 B.n562 10.6151
R979 B.n564 B.n563 10.6151
R980 B.n565 B.n564 10.6151
R981 B.n567 B.n565 10.6151
R982 B.n568 B.n567 10.6151
R983 B.n569 B.n568 10.6151
R984 B.n570 B.n569 10.6151
R985 B.n572 B.n570 10.6151
R986 B.n573 B.n572 10.6151
R987 B.n574 B.n573 10.6151
R988 B.n575 B.n574 10.6151
R989 B.n576 B.n575 10.6151
R990 B.n444 B.n279 10.6151
R991 B.n439 B.n279 10.6151
R992 B.n439 B.n438 10.6151
R993 B.n438 B.n437 10.6151
R994 B.n437 B.n434 10.6151
R995 B.n434 B.n433 10.6151
R996 B.n433 B.n430 10.6151
R997 B.n430 B.n429 10.6151
R998 B.n429 B.n426 10.6151
R999 B.n426 B.n425 10.6151
R1000 B.n425 B.n422 10.6151
R1001 B.n422 B.n421 10.6151
R1002 B.n421 B.n418 10.6151
R1003 B.n418 B.n417 10.6151
R1004 B.n417 B.n414 10.6151
R1005 B.n414 B.n413 10.6151
R1006 B.n413 B.n410 10.6151
R1007 B.n410 B.n409 10.6151
R1008 B.n409 B.n406 10.6151
R1009 B.n406 B.n405 10.6151
R1010 B.n405 B.n402 10.6151
R1011 B.n402 B.n401 10.6151
R1012 B.n401 B.n398 10.6151
R1013 B.n398 B.n397 10.6151
R1014 B.n397 B.n394 10.6151
R1015 B.n394 B.n393 10.6151
R1016 B.n390 B.n389 10.6151
R1017 B.n389 B.n386 10.6151
R1018 B.n386 B.n385 10.6151
R1019 B.n385 B.n382 10.6151
R1020 B.n382 B.n381 10.6151
R1021 B.n381 B.n378 10.6151
R1022 B.n378 B.n377 10.6151
R1023 B.n377 B.n374 10.6151
R1024 B.n374 B.n373 10.6151
R1025 B.n370 B.n369 10.6151
R1026 B.n369 B.n366 10.6151
R1027 B.n366 B.n365 10.6151
R1028 B.n365 B.n362 10.6151
R1029 B.n362 B.n361 10.6151
R1030 B.n361 B.n358 10.6151
R1031 B.n358 B.n357 10.6151
R1032 B.n357 B.n354 10.6151
R1033 B.n354 B.n353 10.6151
R1034 B.n353 B.n350 10.6151
R1035 B.n350 B.n349 10.6151
R1036 B.n349 B.n346 10.6151
R1037 B.n346 B.n345 10.6151
R1038 B.n345 B.n342 10.6151
R1039 B.n342 B.n341 10.6151
R1040 B.n341 B.n338 10.6151
R1041 B.n338 B.n337 10.6151
R1042 B.n337 B.n334 10.6151
R1043 B.n334 B.n333 10.6151
R1044 B.n333 B.n330 10.6151
R1045 B.n330 B.n329 10.6151
R1046 B.n329 B.n326 10.6151
R1047 B.n326 B.n325 10.6151
R1048 B.n325 B.n322 10.6151
R1049 B.n322 B.n321 10.6151
R1050 B.n321 B.n319 10.6151
R1051 B.n446 B.n445 10.6151
R1052 B.n446 B.n271 10.6151
R1053 B.n456 B.n271 10.6151
R1054 B.n457 B.n456 10.6151
R1055 B.n458 B.n457 10.6151
R1056 B.n458 B.n263 10.6151
R1057 B.n469 B.n263 10.6151
R1058 B.n470 B.n469 10.6151
R1059 B.n471 B.n470 10.6151
R1060 B.n471 B.n256 10.6151
R1061 B.n481 B.n256 10.6151
R1062 B.n482 B.n481 10.6151
R1063 B.n483 B.n482 10.6151
R1064 B.n483 B.n248 10.6151
R1065 B.n493 B.n248 10.6151
R1066 B.n494 B.n493 10.6151
R1067 B.n495 B.n494 10.6151
R1068 B.n495 B.n240 10.6151
R1069 B.n505 B.n240 10.6151
R1070 B.n506 B.n505 10.6151
R1071 B.n507 B.n506 10.6151
R1072 B.n507 B.n232 10.6151
R1073 B.n517 B.n232 10.6151
R1074 B.n518 B.n517 10.6151
R1075 B.n519 B.n518 10.6151
R1076 B.n519 B.n224 10.6151
R1077 B.n530 B.n224 10.6151
R1078 B.n531 B.n530 10.6151
R1079 B.n532 B.n531 10.6151
R1080 B.n532 B.n0 10.6151
R1081 B.n641 B.n1 10.6151
R1082 B.n641 B.n640 10.6151
R1083 B.n640 B.n639 10.6151
R1084 B.n639 B.n10 10.6151
R1085 B.n633 B.n10 10.6151
R1086 B.n633 B.n632 10.6151
R1087 B.n632 B.n631 10.6151
R1088 B.n631 B.n17 10.6151
R1089 B.n625 B.n17 10.6151
R1090 B.n625 B.n624 10.6151
R1091 B.n624 B.n623 10.6151
R1092 B.n623 B.n24 10.6151
R1093 B.n617 B.n24 10.6151
R1094 B.n617 B.n616 10.6151
R1095 B.n616 B.n615 10.6151
R1096 B.n615 B.n31 10.6151
R1097 B.n609 B.n31 10.6151
R1098 B.n609 B.n608 10.6151
R1099 B.n608 B.n607 10.6151
R1100 B.n607 B.n38 10.6151
R1101 B.n601 B.n38 10.6151
R1102 B.n601 B.n600 10.6151
R1103 B.n600 B.n599 10.6151
R1104 B.n599 B.n44 10.6151
R1105 B.n593 B.n44 10.6151
R1106 B.n593 B.n592 10.6151
R1107 B.n592 B.n591 10.6151
R1108 B.n591 B.n52 10.6151
R1109 B.n585 B.n52 10.6151
R1110 B.n585 B.n584 10.6151
R1111 B.n147 B.n146 9.36635
R1112 B.n169 B.n168 9.36635
R1113 B.n393 B.n315 9.36635
R1114 B.n370 B.n318 9.36635
R1115 B.n473 B.t3 8.91099
R1116 B.n603 B.t7 8.91099
R1117 B.n647 B.n0 2.81026
R1118 B.n647 B.n1 2.81026
R1119 B.n148 B.n147 1.24928
R1120 B.n168 B.n167 1.24928
R1121 B.n390 B.n315 1.24928
R1122 B.n373 B.n318 1.24928
R1123 VN VN.t1 129.599
R1124 VN VN.t0 86.6438
R1125 VDD2.n0 VDD2.t1 104.748
R1126 VDD2.n0 VDD2.t0 68.2176
R1127 VDD2 VDD2.n0 0.905672
C0 VDD2 VN 1.81463f
C1 VDD2 VDD1 0.78221f
C2 VN VTAIL 1.87969f
C3 VTAIL VDD1 4.02708f
C4 VN VDD1 0.148581f
C5 VDD2 VP 0.374738f
C6 VTAIL VP 1.89392f
C7 VN VP 5.00911f
C8 VP VDD1 2.03935f
C9 VDD2 VTAIL 4.08605f
C10 VDD2 B 3.865546f
C11 VDD1 B 6.90991f
C12 VTAIL B 5.529978f
C13 VN B 9.13908f
C14 VP B 7.167722f
C15 VDD2.t1 B 1.20605f
C16 VDD2.t0 B 0.885173f
C17 VDD2.n0 B 1.88554f
C18 VN.t0 B 1.34697f
C19 VN.t1 B 1.72688f
C20 VDD1.t0 B 1.28234f
C21 VDD1.t1 B 1.7814f
C22 VTAIL.t3 B 0.914804f
C23 VTAIL.n0 B 1.15701f
C24 VTAIL.t1 B 0.914807f
C25 VTAIL.n1 B 1.19781f
C26 VTAIL.t2 B 0.914804f
C27 VTAIL.n2 B 1.02258f
C28 VTAIL.t0 B 0.914804f
C29 VTAIL.n3 B 0.95146f
C30 VP.t1 B 2.42837f
C31 VP.t0 B 1.8909f
C32 VP.n0 B 2.5927f
.ends

