* NGSPICE file created from diff_pair_sample_0089.ext - technology: sky130A

.subckt diff_pair_sample_0089 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t18 VP.t0 VDD1.t2 w_n2950_n4810# sky130_fd_pr__pfet_01v8 ad=3.16965 pd=19.54 as=3.16965 ps=19.54 w=19.21 l=1.32
X1 VDD2.t9 VN.t0 VTAIL.t4 w_n2950_n4810# sky130_fd_pr__pfet_01v8 ad=7.4919 pd=39.2 as=3.16965 ps=19.54 w=19.21 l=1.32
X2 VDD1.t6 VP.t1 VTAIL.t17 w_n2950_n4810# sky130_fd_pr__pfet_01v8 ad=7.4919 pd=39.2 as=3.16965 ps=19.54 w=19.21 l=1.32
X3 B.t11 B.t9 B.t10 w_n2950_n4810# sky130_fd_pr__pfet_01v8 ad=7.4919 pd=39.2 as=0 ps=0 w=19.21 l=1.32
X4 VDD2.t8 VN.t1 VTAIL.t19 w_n2950_n4810# sky130_fd_pr__pfet_01v8 ad=3.16965 pd=19.54 as=3.16965 ps=19.54 w=19.21 l=1.32
X5 VDD2.t7 VN.t2 VTAIL.t0 w_n2950_n4810# sky130_fd_pr__pfet_01v8 ad=3.16965 pd=19.54 as=7.4919 ps=39.2 w=19.21 l=1.32
X6 VTAIL.t7 VN.t3 VDD2.t6 w_n2950_n4810# sky130_fd_pr__pfet_01v8 ad=3.16965 pd=19.54 as=3.16965 ps=19.54 w=19.21 l=1.32
X7 VDD2.t5 VN.t4 VTAIL.t8 w_n2950_n4810# sky130_fd_pr__pfet_01v8 ad=3.16965 pd=19.54 as=3.16965 ps=19.54 w=19.21 l=1.32
X8 VTAIL.t3 VN.t5 VDD2.t4 w_n2950_n4810# sky130_fd_pr__pfet_01v8 ad=3.16965 pd=19.54 as=3.16965 ps=19.54 w=19.21 l=1.32
X9 VDD2.t3 VN.t6 VTAIL.t2 w_n2950_n4810# sky130_fd_pr__pfet_01v8 ad=7.4919 pd=39.2 as=3.16965 ps=19.54 w=19.21 l=1.32
X10 VTAIL.t16 VP.t2 VDD1.t5 w_n2950_n4810# sky130_fd_pr__pfet_01v8 ad=3.16965 pd=19.54 as=3.16965 ps=19.54 w=19.21 l=1.32
X11 B.t8 B.t6 B.t7 w_n2950_n4810# sky130_fd_pr__pfet_01v8 ad=7.4919 pd=39.2 as=0 ps=0 w=19.21 l=1.32
X12 VDD1.t1 VP.t3 VTAIL.t15 w_n2950_n4810# sky130_fd_pr__pfet_01v8 ad=3.16965 pd=19.54 as=7.4919 ps=39.2 w=19.21 l=1.32
X13 VTAIL.t14 VP.t4 VDD1.t0 w_n2950_n4810# sky130_fd_pr__pfet_01v8 ad=3.16965 pd=19.54 as=3.16965 ps=19.54 w=19.21 l=1.32
X14 VDD1.t9 VP.t5 VTAIL.t13 w_n2950_n4810# sky130_fd_pr__pfet_01v8 ad=3.16965 pd=19.54 as=7.4919 ps=39.2 w=19.21 l=1.32
X15 VDD1.t8 VP.t6 VTAIL.t12 w_n2950_n4810# sky130_fd_pr__pfet_01v8 ad=3.16965 pd=19.54 as=3.16965 ps=19.54 w=19.21 l=1.32
X16 VTAIL.t6 VN.t7 VDD2.t2 w_n2950_n4810# sky130_fd_pr__pfet_01v8 ad=3.16965 pd=19.54 as=3.16965 ps=19.54 w=19.21 l=1.32
X17 VDD2.t1 VN.t8 VTAIL.t1 w_n2950_n4810# sky130_fd_pr__pfet_01v8 ad=3.16965 pd=19.54 as=7.4919 ps=39.2 w=19.21 l=1.32
X18 VTAIL.t5 VN.t9 VDD2.t0 w_n2950_n4810# sky130_fd_pr__pfet_01v8 ad=3.16965 pd=19.54 as=3.16965 ps=19.54 w=19.21 l=1.32
X19 VTAIL.t11 VP.t7 VDD1.t4 w_n2950_n4810# sky130_fd_pr__pfet_01v8 ad=3.16965 pd=19.54 as=3.16965 ps=19.54 w=19.21 l=1.32
X20 VDD1.t3 VP.t8 VTAIL.t10 w_n2950_n4810# sky130_fd_pr__pfet_01v8 ad=7.4919 pd=39.2 as=3.16965 ps=19.54 w=19.21 l=1.32
X21 B.t5 B.t3 B.t4 w_n2950_n4810# sky130_fd_pr__pfet_01v8 ad=7.4919 pd=39.2 as=0 ps=0 w=19.21 l=1.32
X22 B.t2 B.t0 B.t1 w_n2950_n4810# sky130_fd_pr__pfet_01v8 ad=7.4919 pd=39.2 as=0 ps=0 w=19.21 l=1.32
X23 VDD1.t7 VP.t9 VTAIL.t9 w_n2950_n4810# sky130_fd_pr__pfet_01v8 ad=3.16965 pd=19.54 as=3.16965 ps=19.54 w=19.21 l=1.32
R0 VP.n14 VP.t1 381.712
R1 VP.n3 VP.t9 350.728
R2 VP.n7 VP.t8 350.728
R3 VP.n5 VP.t7 350.728
R4 VP.n48 VP.t4 350.728
R5 VP.n55 VP.t3 350.728
R6 VP.n11 VP.t6 350.728
R7 VP.n31 VP.t5 350.728
R8 VP.n24 VP.t0 350.728
R9 VP.n13 VP.t2 350.728
R10 VP.n33 VP.n7 171.088
R11 VP.n56 VP.n55 171.088
R12 VP.n32 VP.n31 171.088
R13 VP.n16 VP.n15 161.3
R14 VP.n17 VP.n12 161.3
R15 VP.n19 VP.n18 161.3
R16 VP.n20 VP.n11 161.3
R17 VP.n22 VP.n21 161.3
R18 VP.n23 VP.n10 161.3
R19 VP.n26 VP.n25 161.3
R20 VP.n27 VP.n9 161.3
R21 VP.n29 VP.n28 161.3
R22 VP.n30 VP.n8 161.3
R23 VP.n54 VP.n0 161.3
R24 VP.n53 VP.n52 161.3
R25 VP.n51 VP.n1 161.3
R26 VP.n50 VP.n49 161.3
R27 VP.n47 VP.n2 161.3
R28 VP.n46 VP.n45 161.3
R29 VP.n44 VP.n3 161.3
R30 VP.n43 VP.n42 161.3
R31 VP.n41 VP.n4 161.3
R32 VP.n40 VP.n39 161.3
R33 VP.n38 VP.n37 161.3
R34 VP.n36 VP.n6 161.3
R35 VP.n35 VP.n34 161.3
R36 VP.n14 VP.n13 57.1957
R37 VP.n42 VP.n41 56.5193
R38 VP.n47 VP.n46 56.5193
R39 VP.n23 VP.n22 56.5193
R40 VP.n18 VP.n17 56.5193
R41 VP.n33 VP.n32 51.5725
R42 VP.n37 VP.n36 42.9216
R43 VP.n53 VP.n1 42.9216
R44 VP.n29 VP.n9 42.9216
R45 VP.n36 VP.n35 38.0652
R46 VP.n54 VP.n53 38.0652
R47 VP.n30 VP.n29 38.0652
R48 VP.n15 VP.n14 26.7159
R49 VP.n41 VP.n40 24.4675
R50 VP.n42 VP.n3 24.4675
R51 VP.n46 VP.n3 24.4675
R52 VP.n49 VP.n47 24.4675
R53 VP.n25 VP.n23 24.4675
R54 VP.n18 VP.n11 24.4675
R55 VP.n22 VP.n11 24.4675
R56 VP.n17 VP.n16 24.4675
R57 VP.n37 VP.n5 17.1274
R58 VP.n48 VP.n1 17.1274
R59 VP.n24 VP.n9 17.1274
R60 VP.n35 VP.n7 14.6807
R61 VP.n55 VP.n54 14.6807
R62 VP.n31 VP.n30 14.6807
R63 VP.n40 VP.n5 7.3406
R64 VP.n49 VP.n48 7.3406
R65 VP.n25 VP.n24 7.3406
R66 VP.n16 VP.n13 7.3406
R67 VP.n15 VP.n12 0.189894
R68 VP.n19 VP.n12 0.189894
R69 VP.n20 VP.n19 0.189894
R70 VP.n21 VP.n20 0.189894
R71 VP.n21 VP.n10 0.189894
R72 VP.n26 VP.n10 0.189894
R73 VP.n27 VP.n26 0.189894
R74 VP.n28 VP.n27 0.189894
R75 VP.n28 VP.n8 0.189894
R76 VP.n32 VP.n8 0.189894
R77 VP.n34 VP.n33 0.189894
R78 VP.n34 VP.n6 0.189894
R79 VP.n38 VP.n6 0.189894
R80 VP.n39 VP.n38 0.189894
R81 VP.n39 VP.n4 0.189894
R82 VP.n43 VP.n4 0.189894
R83 VP.n44 VP.n43 0.189894
R84 VP.n45 VP.n44 0.189894
R85 VP.n45 VP.n2 0.189894
R86 VP.n50 VP.n2 0.189894
R87 VP.n51 VP.n50 0.189894
R88 VP.n52 VP.n51 0.189894
R89 VP.n52 VP.n0 0.189894
R90 VP.n56 VP.n0 0.189894
R91 VP VP.n56 0.0516364
R92 VDD1.n1 VDD1.t6 69.2251
R93 VDD1.n3 VDD1.t3 69.2248
R94 VDD1.n5 VDD1.n4 67.122
R95 VDD1.n1 VDD1.n0 66.1106
R96 VDD1.n3 VDD1.n2 66.1105
R97 VDD1.n7 VDD1.n6 66.1104
R98 VDD1.n7 VDD1.n5 48.3263
R99 VDD1.n6 VDD1.t2 1.69259
R100 VDD1.n6 VDD1.t9 1.69259
R101 VDD1.n0 VDD1.t5 1.69259
R102 VDD1.n0 VDD1.t8 1.69259
R103 VDD1.n4 VDD1.t0 1.69259
R104 VDD1.n4 VDD1.t1 1.69259
R105 VDD1.n2 VDD1.t4 1.69259
R106 VDD1.n2 VDD1.t7 1.69259
R107 VDD1 VDD1.n7 1.00912
R108 VDD1 VDD1.n1 0.414293
R109 VDD1.n5 VDD1.n3 0.300757
R110 VTAIL.n11 VTAIL.t0 51.1239
R111 VTAIL.n17 VTAIL.t1 51.1236
R112 VTAIL.n2 VTAIL.t15 51.1236
R113 VTAIL.n16 VTAIL.t13 51.1236
R114 VTAIL.n15 VTAIL.n14 49.4318
R115 VTAIL.n13 VTAIL.n12 49.4318
R116 VTAIL.n10 VTAIL.n9 49.4318
R117 VTAIL.n8 VTAIL.n7 49.4318
R118 VTAIL.n19 VTAIL.n18 49.4317
R119 VTAIL.n1 VTAIL.n0 49.4317
R120 VTAIL.n4 VTAIL.n3 49.4317
R121 VTAIL.n6 VTAIL.n5 49.4317
R122 VTAIL.n8 VTAIL.n6 31.7721
R123 VTAIL.n17 VTAIL.n16 30.3496
R124 VTAIL.n18 VTAIL.t8 1.69259
R125 VTAIL.n18 VTAIL.t7 1.69259
R126 VTAIL.n0 VTAIL.t2 1.69259
R127 VTAIL.n0 VTAIL.t3 1.69259
R128 VTAIL.n3 VTAIL.t9 1.69259
R129 VTAIL.n3 VTAIL.t14 1.69259
R130 VTAIL.n5 VTAIL.t10 1.69259
R131 VTAIL.n5 VTAIL.t11 1.69259
R132 VTAIL.n14 VTAIL.t12 1.69259
R133 VTAIL.n14 VTAIL.t18 1.69259
R134 VTAIL.n12 VTAIL.t17 1.69259
R135 VTAIL.n12 VTAIL.t16 1.69259
R136 VTAIL.n9 VTAIL.t19 1.69259
R137 VTAIL.n9 VTAIL.t6 1.69259
R138 VTAIL.n7 VTAIL.t4 1.69259
R139 VTAIL.n7 VTAIL.t5 1.69259
R140 VTAIL.n10 VTAIL.n8 1.42291
R141 VTAIL.n11 VTAIL.n10 1.42291
R142 VTAIL.n15 VTAIL.n13 1.42291
R143 VTAIL.n16 VTAIL.n15 1.42291
R144 VTAIL.n6 VTAIL.n4 1.42291
R145 VTAIL.n4 VTAIL.n2 1.42291
R146 VTAIL.n19 VTAIL.n17 1.42291
R147 VTAIL.n13 VTAIL.n11 1.18153
R148 VTAIL.n2 VTAIL.n1 1.18153
R149 VTAIL VTAIL.n1 1.1255
R150 VTAIL VTAIL.n19 0.297914
R151 VN.n6 VN.t6 381.712
R152 VN.n32 VN.t2 381.712
R153 VN.n3 VN.t4 350.728
R154 VN.n5 VN.t5 350.728
R155 VN.n16 VN.t3 350.728
R156 VN.n23 VN.t8 350.728
R157 VN.n29 VN.t1 350.728
R158 VN.n31 VN.t7 350.728
R159 VN.n28 VN.t9 350.728
R160 VN.n48 VN.t0 350.728
R161 VN.n24 VN.n23 171.088
R162 VN.n49 VN.n48 171.088
R163 VN.n47 VN.n25 161.3
R164 VN.n46 VN.n45 161.3
R165 VN.n44 VN.n26 161.3
R166 VN.n43 VN.n42 161.3
R167 VN.n41 VN.n27 161.3
R168 VN.n40 VN.n39 161.3
R169 VN.n38 VN.n29 161.3
R170 VN.n37 VN.n36 161.3
R171 VN.n35 VN.n30 161.3
R172 VN.n34 VN.n33 161.3
R173 VN.n22 VN.n0 161.3
R174 VN.n21 VN.n20 161.3
R175 VN.n19 VN.n1 161.3
R176 VN.n18 VN.n17 161.3
R177 VN.n15 VN.n2 161.3
R178 VN.n14 VN.n13 161.3
R179 VN.n12 VN.n3 161.3
R180 VN.n11 VN.n10 161.3
R181 VN.n9 VN.n4 161.3
R182 VN.n8 VN.n7 161.3
R183 VN.n6 VN.n5 57.1957
R184 VN.n32 VN.n31 57.1957
R185 VN.n10 VN.n9 56.5193
R186 VN.n15 VN.n14 56.5193
R187 VN.n36 VN.n35 56.5193
R188 VN.n41 VN.n40 56.5193
R189 VN VN.n49 51.9532
R190 VN.n21 VN.n1 42.9216
R191 VN.n46 VN.n26 42.9216
R192 VN.n22 VN.n21 38.0652
R193 VN.n47 VN.n46 38.0652
R194 VN.n33 VN.n32 26.7159
R195 VN.n7 VN.n6 26.7159
R196 VN.n9 VN.n8 24.4675
R197 VN.n10 VN.n3 24.4675
R198 VN.n14 VN.n3 24.4675
R199 VN.n17 VN.n15 24.4675
R200 VN.n35 VN.n34 24.4675
R201 VN.n40 VN.n29 24.4675
R202 VN.n36 VN.n29 24.4675
R203 VN.n42 VN.n41 24.4675
R204 VN.n16 VN.n1 17.1274
R205 VN.n28 VN.n26 17.1274
R206 VN.n23 VN.n22 14.6807
R207 VN.n48 VN.n47 14.6807
R208 VN.n8 VN.n5 7.3406
R209 VN.n17 VN.n16 7.3406
R210 VN.n34 VN.n31 7.3406
R211 VN.n42 VN.n28 7.3406
R212 VN.n49 VN.n25 0.189894
R213 VN.n45 VN.n25 0.189894
R214 VN.n45 VN.n44 0.189894
R215 VN.n44 VN.n43 0.189894
R216 VN.n43 VN.n27 0.189894
R217 VN.n39 VN.n27 0.189894
R218 VN.n39 VN.n38 0.189894
R219 VN.n38 VN.n37 0.189894
R220 VN.n37 VN.n30 0.189894
R221 VN.n33 VN.n30 0.189894
R222 VN.n7 VN.n4 0.189894
R223 VN.n11 VN.n4 0.189894
R224 VN.n12 VN.n11 0.189894
R225 VN.n13 VN.n12 0.189894
R226 VN.n13 VN.n2 0.189894
R227 VN.n18 VN.n2 0.189894
R228 VN.n19 VN.n18 0.189894
R229 VN.n20 VN.n19 0.189894
R230 VN.n20 VN.n0 0.189894
R231 VN.n24 VN.n0 0.189894
R232 VN VN.n24 0.0516364
R233 VDD2.n1 VDD2.t3 69.2248
R234 VDD2.n4 VDD2.t9 67.8026
R235 VDD2.n3 VDD2.n2 67.122
R236 VDD2 VDD2.n7 67.119
R237 VDD2.n6 VDD2.n5 66.1106
R238 VDD2.n1 VDD2.n0 66.1105
R239 VDD2.n4 VDD2.n3 47.0321
R240 VDD2.n7 VDD2.t2 1.69259
R241 VDD2.n7 VDD2.t7 1.69259
R242 VDD2.n5 VDD2.t0 1.69259
R243 VDD2.n5 VDD2.t8 1.69259
R244 VDD2.n2 VDD2.t6 1.69259
R245 VDD2.n2 VDD2.t1 1.69259
R246 VDD2.n0 VDD2.t4 1.69259
R247 VDD2.n0 VDD2.t5 1.69259
R248 VDD2.n6 VDD2.n4 1.42291
R249 VDD2 VDD2.n6 0.414293
R250 VDD2.n3 VDD2.n1 0.300757
R251 B.n591 B.n92 585
R252 B.n593 B.n592 585
R253 B.n594 B.n91 585
R254 B.n596 B.n595 585
R255 B.n597 B.n90 585
R256 B.n599 B.n598 585
R257 B.n600 B.n89 585
R258 B.n602 B.n601 585
R259 B.n603 B.n88 585
R260 B.n605 B.n604 585
R261 B.n606 B.n87 585
R262 B.n608 B.n607 585
R263 B.n609 B.n86 585
R264 B.n611 B.n610 585
R265 B.n612 B.n85 585
R266 B.n614 B.n613 585
R267 B.n615 B.n84 585
R268 B.n617 B.n616 585
R269 B.n618 B.n83 585
R270 B.n620 B.n619 585
R271 B.n621 B.n82 585
R272 B.n623 B.n622 585
R273 B.n624 B.n81 585
R274 B.n626 B.n625 585
R275 B.n627 B.n80 585
R276 B.n629 B.n628 585
R277 B.n630 B.n79 585
R278 B.n632 B.n631 585
R279 B.n633 B.n78 585
R280 B.n635 B.n634 585
R281 B.n636 B.n77 585
R282 B.n638 B.n637 585
R283 B.n639 B.n76 585
R284 B.n641 B.n640 585
R285 B.n642 B.n75 585
R286 B.n644 B.n643 585
R287 B.n645 B.n74 585
R288 B.n647 B.n646 585
R289 B.n648 B.n73 585
R290 B.n650 B.n649 585
R291 B.n651 B.n72 585
R292 B.n653 B.n652 585
R293 B.n654 B.n71 585
R294 B.n656 B.n655 585
R295 B.n657 B.n70 585
R296 B.n659 B.n658 585
R297 B.n660 B.n69 585
R298 B.n662 B.n661 585
R299 B.n663 B.n68 585
R300 B.n665 B.n664 585
R301 B.n666 B.n67 585
R302 B.n668 B.n667 585
R303 B.n669 B.n66 585
R304 B.n671 B.n670 585
R305 B.n672 B.n65 585
R306 B.n674 B.n673 585
R307 B.n675 B.n64 585
R308 B.n677 B.n676 585
R309 B.n678 B.n63 585
R310 B.n680 B.n679 585
R311 B.n681 B.n62 585
R312 B.n683 B.n682 585
R313 B.n684 B.n59 585
R314 B.n687 B.n686 585
R315 B.n688 B.n58 585
R316 B.n690 B.n689 585
R317 B.n691 B.n57 585
R318 B.n693 B.n692 585
R319 B.n694 B.n56 585
R320 B.n696 B.n695 585
R321 B.n697 B.n55 585
R322 B.n699 B.n698 585
R323 B.n701 B.n700 585
R324 B.n702 B.n51 585
R325 B.n704 B.n703 585
R326 B.n705 B.n50 585
R327 B.n707 B.n706 585
R328 B.n708 B.n49 585
R329 B.n710 B.n709 585
R330 B.n711 B.n48 585
R331 B.n713 B.n712 585
R332 B.n714 B.n47 585
R333 B.n716 B.n715 585
R334 B.n717 B.n46 585
R335 B.n719 B.n718 585
R336 B.n720 B.n45 585
R337 B.n722 B.n721 585
R338 B.n723 B.n44 585
R339 B.n725 B.n724 585
R340 B.n726 B.n43 585
R341 B.n728 B.n727 585
R342 B.n729 B.n42 585
R343 B.n731 B.n730 585
R344 B.n732 B.n41 585
R345 B.n734 B.n733 585
R346 B.n735 B.n40 585
R347 B.n737 B.n736 585
R348 B.n738 B.n39 585
R349 B.n740 B.n739 585
R350 B.n741 B.n38 585
R351 B.n743 B.n742 585
R352 B.n744 B.n37 585
R353 B.n746 B.n745 585
R354 B.n747 B.n36 585
R355 B.n749 B.n748 585
R356 B.n750 B.n35 585
R357 B.n752 B.n751 585
R358 B.n753 B.n34 585
R359 B.n755 B.n754 585
R360 B.n756 B.n33 585
R361 B.n758 B.n757 585
R362 B.n759 B.n32 585
R363 B.n761 B.n760 585
R364 B.n762 B.n31 585
R365 B.n764 B.n763 585
R366 B.n765 B.n30 585
R367 B.n767 B.n766 585
R368 B.n768 B.n29 585
R369 B.n770 B.n769 585
R370 B.n771 B.n28 585
R371 B.n773 B.n772 585
R372 B.n774 B.n27 585
R373 B.n776 B.n775 585
R374 B.n777 B.n26 585
R375 B.n779 B.n778 585
R376 B.n780 B.n25 585
R377 B.n782 B.n781 585
R378 B.n783 B.n24 585
R379 B.n785 B.n784 585
R380 B.n786 B.n23 585
R381 B.n788 B.n787 585
R382 B.n789 B.n22 585
R383 B.n791 B.n790 585
R384 B.n792 B.n21 585
R385 B.n794 B.n793 585
R386 B.n590 B.n589 585
R387 B.n588 B.n93 585
R388 B.n587 B.n586 585
R389 B.n585 B.n94 585
R390 B.n584 B.n583 585
R391 B.n582 B.n95 585
R392 B.n581 B.n580 585
R393 B.n579 B.n96 585
R394 B.n578 B.n577 585
R395 B.n576 B.n97 585
R396 B.n575 B.n574 585
R397 B.n573 B.n98 585
R398 B.n572 B.n571 585
R399 B.n570 B.n99 585
R400 B.n569 B.n568 585
R401 B.n567 B.n100 585
R402 B.n566 B.n565 585
R403 B.n564 B.n101 585
R404 B.n563 B.n562 585
R405 B.n561 B.n102 585
R406 B.n560 B.n559 585
R407 B.n558 B.n103 585
R408 B.n557 B.n556 585
R409 B.n555 B.n104 585
R410 B.n554 B.n553 585
R411 B.n552 B.n105 585
R412 B.n551 B.n550 585
R413 B.n549 B.n106 585
R414 B.n548 B.n547 585
R415 B.n546 B.n107 585
R416 B.n545 B.n544 585
R417 B.n543 B.n108 585
R418 B.n542 B.n541 585
R419 B.n540 B.n109 585
R420 B.n539 B.n538 585
R421 B.n537 B.n110 585
R422 B.n536 B.n535 585
R423 B.n534 B.n111 585
R424 B.n533 B.n532 585
R425 B.n531 B.n112 585
R426 B.n530 B.n529 585
R427 B.n528 B.n113 585
R428 B.n527 B.n526 585
R429 B.n525 B.n114 585
R430 B.n524 B.n523 585
R431 B.n522 B.n115 585
R432 B.n521 B.n520 585
R433 B.n519 B.n116 585
R434 B.n518 B.n517 585
R435 B.n516 B.n117 585
R436 B.n515 B.n514 585
R437 B.n513 B.n118 585
R438 B.n512 B.n511 585
R439 B.n510 B.n119 585
R440 B.n509 B.n508 585
R441 B.n507 B.n120 585
R442 B.n506 B.n505 585
R443 B.n504 B.n121 585
R444 B.n503 B.n502 585
R445 B.n501 B.n122 585
R446 B.n500 B.n499 585
R447 B.n498 B.n123 585
R448 B.n497 B.n496 585
R449 B.n495 B.n124 585
R450 B.n494 B.n493 585
R451 B.n492 B.n125 585
R452 B.n491 B.n490 585
R453 B.n489 B.n126 585
R454 B.n488 B.n487 585
R455 B.n486 B.n127 585
R456 B.n485 B.n484 585
R457 B.n483 B.n128 585
R458 B.n482 B.n481 585
R459 B.n480 B.n129 585
R460 B.n479 B.n478 585
R461 B.n275 B.n274 585
R462 B.n276 B.n201 585
R463 B.n278 B.n277 585
R464 B.n279 B.n200 585
R465 B.n281 B.n280 585
R466 B.n282 B.n199 585
R467 B.n284 B.n283 585
R468 B.n285 B.n198 585
R469 B.n287 B.n286 585
R470 B.n288 B.n197 585
R471 B.n290 B.n289 585
R472 B.n291 B.n196 585
R473 B.n293 B.n292 585
R474 B.n294 B.n195 585
R475 B.n296 B.n295 585
R476 B.n297 B.n194 585
R477 B.n299 B.n298 585
R478 B.n300 B.n193 585
R479 B.n302 B.n301 585
R480 B.n303 B.n192 585
R481 B.n305 B.n304 585
R482 B.n306 B.n191 585
R483 B.n308 B.n307 585
R484 B.n309 B.n190 585
R485 B.n311 B.n310 585
R486 B.n312 B.n189 585
R487 B.n314 B.n313 585
R488 B.n315 B.n188 585
R489 B.n317 B.n316 585
R490 B.n318 B.n187 585
R491 B.n320 B.n319 585
R492 B.n321 B.n186 585
R493 B.n323 B.n322 585
R494 B.n324 B.n185 585
R495 B.n326 B.n325 585
R496 B.n327 B.n184 585
R497 B.n329 B.n328 585
R498 B.n330 B.n183 585
R499 B.n332 B.n331 585
R500 B.n333 B.n182 585
R501 B.n335 B.n334 585
R502 B.n336 B.n181 585
R503 B.n338 B.n337 585
R504 B.n339 B.n180 585
R505 B.n341 B.n340 585
R506 B.n342 B.n179 585
R507 B.n344 B.n343 585
R508 B.n345 B.n178 585
R509 B.n347 B.n346 585
R510 B.n348 B.n177 585
R511 B.n350 B.n349 585
R512 B.n351 B.n176 585
R513 B.n353 B.n352 585
R514 B.n354 B.n175 585
R515 B.n356 B.n355 585
R516 B.n357 B.n174 585
R517 B.n359 B.n358 585
R518 B.n360 B.n173 585
R519 B.n362 B.n361 585
R520 B.n363 B.n172 585
R521 B.n365 B.n364 585
R522 B.n366 B.n171 585
R523 B.n368 B.n367 585
R524 B.n370 B.n369 585
R525 B.n371 B.n167 585
R526 B.n373 B.n372 585
R527 B.n374 B.n166 585
R528 B.n376 B.n375 585
R529 B.n377 B.n165 585
R530 B.n379 B.n378 585
R531 B.n380 B.n164 585
R532 B.n382 B.n381 585
R533 B.n384 B.n161 585
R534 B.n386 B.n385 585
R535 B.n387 B.n160 585
R536 B.n389 B.n388 585
R537 B.n390 B.n159 585
R538 B.n392 B.n391 585
R539 B.n393 B.n158 585
R540 B.n395 B.n394 585
R541 B.n396 B.n157 585
R542 B.n398 B.n397 585
R543 B.n399 B.n156 585
R544 B.n401 B.n400 585
R545 B.n402 B.n155 585
R546 B.n404 B.n403 585
R547 B.n405 B.n154 585
R548 B.n407 B.n406 585
R549 B.n408 B.n153 585
R550 B.n410 B.n409 585
R551 B.n411 B.n152 585
R552 B.n413 B.n412 585
R553 B.n414 B.n151 585
R554 B.n416 B.n415 585
R555 B.n417 B.n150 585
R556 B.n419 B.n418 585
R557 B.n420 B.n149 585
R558 B.n422 B.n421 585
R559 B.n423 B.n148 585
R560 B.n425 B.n424 585
R561 B.n426 B.n147 585
R562 B.n428 B.n427 585
R563 B.n429 B.n146 585
R564 B.n431 B.n430 585
R565 B.n432 B.n145 585
R566 B.n434 B.n433 585
R567 B.n435 B.n144 585
R568 B.n437 B.n436 585
R569 B.n438 B.n143 585
R570 B.n440 B.n439 585
R571 B.n441 B.n142 585
R572 B.n443 B.n442 585
R573 B.n444 B.n141 585
R574 B.n446 B.n445 585
R575 B.n447 B.n140 585
R576 B.n449 B.n448 585
R577 B.n450 B.n139 585
R578 B.n452 B.n451 585
R579 B.n453 B.n138 585
R580 B.n455 B.n454 585
R581 B.n456 B.n137 585
R582 B.n458 B.n457 585
R583 B.n459 B.n136 585
R584 B.n461 B.n460 585
R585 B.n462 B.n135 585
R586 B.n464 B.n463 585
R587 B.n465 B.n134 585
R588 B.n467 B.n466 585
R589 B.n468 B.n133 585
R590 B.n470 B.n469 585
R591 B.n471 B.n132 585
R592 B.n473 B.n472 585
R593 B.n474 B.n131 585
R594 B.n476 B.n475 585
R595 B.n477 B.n130 585
R596 B.n273 B.n202 585
R597 B.n272 B.n271 585
R598 B.n270 B.n203 585
R599 B.n269 B.n268 585
R600 B.n267 B.n204 585
R601 B.n266 B.n265 585
R602 B.n264 B.n205 585
R603 B.n263 B.n262 585
R604 B.n261 B.n206 585
R605 B.n260 B.n259 585
R606 B.n258 B.n207 585
R607 B.n257 B.n256 585
R608 B.n255 B.n208 585
R609 B.n254 B.n253 585
R610 B.n252 B.n209 585
R611 B.n251 B.n250 585
R612 B.n249 B.n210 585
R613 B.n248 B.n247 585
R614 B.n246 B.n211 585
R615 B.n245 B.n244 585
R616 B.n243 B.n212 585
R617 B.n242 B.n241 585
R618 B.n240 B.n213 585
R619 B.n239 B.n238 585
R620 B.n237 B.n214 585
R621 B.n236 B.n235 585
R622 B.n234 B.n215 585
R623 B.n233 B.n232 585
R624 B.n231 B.n216 585
R625 B.n230 B.n229 585
R626 B.n228 B.n217 585
R627 B.n227 B.n226 585
R628 B.n225 B.n218 585
R629 B.n224 B.n223 585
R630 B.n222 B.n219 585
R631 B.n221 B.n220 585
R632 B.n2 B.n0 585
R633 B.n849 B.n1 585
R634 B.n848 B.n847 585
R635 B.n846 B.n3 585
R636 B.n845 B.n844 585
R637 B.n843 B.n4 585
R638 B.n842 B.n841 585
R639 B.n840 B.n5 585
R640 B.n839 B.n838 585
R641 B.n837 B.n6 585
R642 B.n836 B.n835 585
R643 B.n834 B.n7 585
R644 B.n833 B.n832 585
R645 B.n831 B.n8 585
R646 B.n830 B.n829 585
R647 B.n828 B.n9 585
R648 B.n827 B.n826 585
R649 B.n825 B.n10 585
R650 B.n824 B.n823 585
R651 B.n822 B.n11 585
R652 B.n821 B.n820 585
R653 B.n819 B.n12 585
R654 B.n818 B.n817 585
R655 B.n816 B.n13 585
R656 B.n815 B.n814 585
R657 B.n813 B.n14 585
R658 B.n812 B.n811 585
R659 B.n810 B.n15 585
R660 B.n809 B.n808 585
R661 B.n807 B.n16 585
R662 B.n806 B.n805 585
R663 B.n804 B.n17 585
R664 B.n803 B.n802 585
R665 B.n801 B.n18 585
R666 B.n800 B.n799 585
R667 B.n798 B.n19 585
R668 B.n797 B.n796 585
R669 B.n795 B.n20 585
R670 B.n851 B.n850 585
R671 B.n162 B.t3 555.428
R672 B.n168 B.t0 555.428
R673 B.n52 B.t9 555.428
R674 B.n60 B.t6 555.428
R675 B.n274 B.n273 554.963
R676 B.n795 B.n794 554.963
R677 B.n478 B.n477 554.963
R678 B.n591 B.n590 554.963
R679 B.n273 B.n272 163.367
R680 B.n272 B.n203 163.367
R681 B.n268 B.n203 163.367
R682 B.n268 B.n267 163.367
R683 B.n267 B.n266 163.367
R684 B.n266 B.n205 163.367
R685 B.n262 B.n205 163.367
R686 B.n262 B.n261 163.367
R687 B.n261 B.n260 163.367
R688 B.n260 B.n207 163.367
R689 B.n256 B.n207 163.367
R690 B.n256 B.n255 163.367
R691 B.n255 B.n254 163.367
R692 B.n254 B.n209 163.367
R693 B.n250 B.n209 163.367
R694 B.n250 B.n249 163.367
R695 B.n249 B.n248 163.367
R696 B.n248 B.n211 163.367
R697 B.n244 B.n211 163.367
R698 B.n244 B.n243 163.367
R699 B.n243 B.n242 163.367
R700 B.n242 B.n213 163.367
R701 B.n238 B.n213 163.367
R702 B.n238 B.n237 163.367
R703 B.n237 B.n236 163.367
R704 B.n236 B.n215 163.367
R705 B.n232 B.n215 163.367
R706 B.n232 B.n231 163.367
R707 B.n231 B.n230 163.367
R708 B.n230 B.n217 163.367
R709 B.n226 B.n217 163.367
R710 B.n226 B.n225 163.367
R711 B.n225 B.n224 163.367
R712 B.n224 B.n219 163.367
R713 B.n220 B.n219 163.367
R714 B.n220 B.n2 163.367
R715 B.n850 B.n2 163.367
R716 B.n850 B.n849 163.367
R717 B.n849 B.n848 163.367
R718 B.n848 B.n3 163.367
R719 B.n844 B.n3 163.367
R720 B.n844 B.n843 163.367
R721 B.n843 B.n842 163.367
R722 B.n842 B.n5 163.367
R723 B.n838 B.n5 163.367
R724 B.n838 B.n837 163.367
R725 B.n837 B.n836 163.367
R726 B.n836 B.n7 163.367
R727 B.n832 B.n7 163.367
R728 B.n832 B.n831 163.367
R729 B.n831 B.n830 163.367
R730 B.n830 B.n9 163.367
R731 B.n826 B.n9 163.367
R732 B.n826 B.n825 163.367
R733 B.n825 B.n824 163.367
R734 B.n824 B.n11 163.367
R735 B.n820 B.n11 163.367
R736 B.n820 B.n819 163.367
R737 B.n819 B.n818 163.367
R738 B.n818 B.n13 163.367
R739 B.n814 B.n13 163.367
R740 B.n814 B.n813 163.367
R741 B.n813 B.n812 163.367
R742 B.n812 B.n15 163.367
R743 B.n808 B.n15 163.367
R744 B.n808 B.n807 163.367
R745 B.n807 B.n806 163.367
R746 B.n806 B.n17 163.367
R747 B.n802 B.n17 163.367
R748 B.n802 B.n801 163.367
R749 B.n801 B.n800 163.367
R750 B.n800 B.n19 163.367
R751 B.n796 B.n19 163.367
R752 B.n796 B.n795 163.367
R753 B.n274 B.n201 163.367
R754 B.n278 B.n201 163.367
R755 B.n279 B.n278 163.367
R756 B.n280 B.n279 163.367
R757 B.n280 B.n199 163.367
R758 B.n284 B.n199 163.367
R759 B.n285 B.n284 163.367
R760 B.n286 B.n285 163.367
R761 B.n286 B.n197 163.367
R762 B.n290 B.n197 163.367
R763 B.n291 B.n290 163.367
R764 B.n292 B.n291 163.367
R765 B.n292 B.n195 163.367
R766 B.n296 B.n195 163.367
R767 B.n297 B.n296 163.367
R768 B.n298 B.n297 163.367
R769 B.n298 B.n193 163.367
R770 B.n302 B.n193 163.367
R771 B.n303 B.n302 163.367
R772 B.n304 B.n303 163.367
R773 B.n304 B.n191 163.367
R774 B.n308 B.n191 163.367
R775 B.n309 B.n308 163.367
R776 B.n310 B.n309 163.367
R777 B.n310 B.n189 163.367
R778 B.n314 B.n189 163.367
R779 B.n315 B.n314 163.367
R780 B.n316 B.n315 163.367
R781 B.n316 B.n187 163.367
R782 B.n320 B.n187 163.367
R783 B.n321 B.n320 163.367
R784 B.n322 B.n321 163.367
R785 B.n322 B.n185 163.367
R786 B.n326 B.n185 163.367
R787 B.n327 B.n326 163.367
R788 B.n328 B.n327 163.367
R789 B.n328 B.n183 163.367
R790 B.n332 B.n183 163.367
R791 B.n333 B.n332 163.367
R792 B.n334 B.n333 163.367
R793 B.n334 B.n181 163.367
R794 B.n338 B.n181 163.367
R795 B.n339 B.n338 163.367
R796 B.n340 B.n339 163.367
R797 B.n340 B.n179 163.367
R798 B.n344 B.n179 163.367
R799 B.n345 B.n344 163.367
R800 B.n346 B.n345 163.367
R801 B.n346 B.n177 163.367
R802 B.n350 B.n177 163.367
R803 B.n351 B.n350 163.367
R804 B.n352 B.n351 163.367
R805 B.n352 B.n175 163.367
R806 B.n356 B.n175 163.367
R807 B.n357 B.n356 163.367
R808 B.n358 B.n357 163.367
R809 B.n358 B.n173 163.367
R810 B.n362 B.n173 163.367
R811 B.n363 B.n362 163.367
R812 B.n364 B.n363 163.367
R813 B.n364 B.n171 163.367
R814 B.n368 B.n171 163.367
R815 B.n369 B.n368 163.367
R816 B.n369 B.n167 163.367
R817 B.n373 B.n167 163.367
R818 B.n374 B.n373 163.367
R819 B.n375 B.n374 163.367
R820 B.n375 B.n165 163.367
R821 B.n379 B.n165 163.367
R822 B.n380 B.n379 163.367
R823 B.n381 B.n380 163.367
R824 B.n381 B.n161 163.367
R825 B.n386 B.n161 163.367
R826 B.n387 B.n386 163.367
R827 B.n388 B.n387 163.367
R828 B.n388 B.n159 163.367
R829 B.n392 B.n159 163.367
R830 B.n393 B.n392 163.367
R831 B.n394 B.n393 163.367
R832 B.n394 B.n157 163.367
R833 B.n398 B.n157 163.367
R834 B.n399 B.n398 163.367
R835 B.n400 B.n399 163.367
R836 B.n400 B.n155 163.367
R837 B.n404 B.n155 163.367
R838 B.n405 B.n404 163.367
R839 B.n406 B.n405 163.367
R840 B.n406 B.n153 163.367
R841 B.n410 B.n153 163.367
R842 B.n411 B.n410 163.367
R843 B.n412 B.n411 163.367
R844 B.n412 B.n151 163.367
R845 B.n416 B.n151 163.367
R846 B.n417 B.n416 163.367
R847 B.n418 B.n417 163.367
R848 B.n418 B.n149 163.367
R849 B.n422 B.n149 163.367
R850 B.n423 B.n422 163.367
R851 B.n424 B.n423 163.367
R852 B.n424 B.n147 163.367
R853 B.n428 B.n147 163.367
R854 B.n429 B.n428 163.367
R855 B.n430 B.n429 163.367
R856 B.n430 B.n145 163.367
R857 B.n434 B.n145 163.367
R858 B.n435 B.n434 163.367
R859 B.n436 B.n435 163.367
R860 B.n436 B.n143 163.367
R861 B.n440 B.n143 163.367
R862 B.n441 B.n440 163.367
R863 B.n442 B.n441 163.367
R864 B.n442 B.n141 163.367
R865 B.n446 B.n141 163.367
R866 B.n447 B.n446 163.367
R867 B.n448 B.n447 163.367
R868 B.n448 B.n139 163.367
R869 B.n452 B.n139 163.367
R870 B.n453 B.n452 163.367
R871 B.n454 B.n453 163.367
R872 B.n454 B.n137 163.367
R873 B.n458 B.n137 163.367
R874 B.n459 B.n458 163.367
R875 B.n460 B.n459 163.367
R876 B.n460 B.n135 163.367
R877 B.n464 B.n135 163.367
R878 B.n465 B.n464 163.367
R879 B.n466 B.n465 163.367
R880 B.n466 B.n133 163.367
R881 B.n470 B.n133 163.367
R882 B.n471 B.n470 163.367
R883 B.n472 B.n471 163.367
R884 B.n472 B.n131 163.367
R885 B.n476 B.n131 163.367
R886 B.n477 B.n476 163.367
R887 B.n478 B.n129 163.367
R888 B.n482 B.n129 163.367
R889 B.n483 B.n482 163.367
R890 B.n484 B.n483 163.367
R891 B.n484 B.n127 163.367
R892 B.n488 B.n127 163.367
R893 B.n489 B.n488 163.367
R894 B.n490 B.n489 163.367
R895 B.n490 B.n125 163.367
R896 B.n494 B.n125 163.367
R897 B.n495 B.n494 163.367
R898 B.n496 B.n495 163.367
R899 B.n496 B.n123 163.367
R900 B.n500 B.n123 163.367
R901 B.n501 B.n500 163.367
R902 B.n502 B.n501 163.367
R903 B.n502 B.n121 163.367
R904 B.n506 B.n121 163.367
R905 B.n507 B.n506 163.367
R906 B.n508 B.n507 163.367
R907 B.n508 B.n119 163.367
R908 B.n512 B.n119 163.367
R909 B.n513 B.n512 163.367
R910 B.n514 B.n513 163.367
R911 B.n514 B.n117 163.367
R912 B.n518 B.n117 163.367
R913 B.n519 B.n518 163.367
R914 B.n520 B.n519 163.367
R915 B.n520 B.n115 163.367
R916 B.n524 B.n115 163.367
R917 B.n525 B.n524 163.367
R918 B.n526 B.n525 163.367
R919 B.n526 B.n113 163.367
R920 B.n530 B.n113 163.367
R921 B.n531 B.n530 163.367
R922 B.n532 B.n531 163.367
R923 B.n532 B.n111 163.367
R924 B.n536 B.n111 163.367
R925 B.n537 B.n536 163.367
R926 B.n538 B.n537 163.367
R927 B.n538 B.n109 163.367
R928 B.n542 B.n109 163.367
R929 B.n543 B.n542 163.367
R930 B.n544 B.n543 163.367
R931 B.n544 B.n107 163.367
R932 B.n548 B.n107 163.367
R933 B.n549 B.n548 163.367
R934 B.n550 B.n549 163.367
R935 B.n550 B.n105 163.367
R936 B.n554 B.n105 163.367
R937 B.n555 B.n554 163.367
R938 B.n556 B.n555 163.367
R939 B.n556 B.n103 163.367
R940 B.n560 B.n103 163.367
R941 B.n561 B.n560 163.367
R942 B.n562 B.n561 163.367
R943 B.n562 B.n101 163.367
R944 B.n566 B.n101 163.367
R945 B.n567 B.n566 163.367
R946 B.n568 B.n567 163.367
R947 B.n568 B.n99 163.367
R948 B.n572 B.n99 163.367
R949 B.n573 B.n572 163.367
R950 B.n574 B.n573 163.367
R951 B.n574 B.n97 163.367
R952 B.n578 B.n97 163.367
R953 B.n579 B.n578 163.367
R954 B.n580 B.n579 163.367
R955 B.n580 B.n95 163.367
R956 B.n584 B.n95 163.367
R957 B.n585 B.n584 163.367
R958 B.n586 B.n585 163.367
R959 B.n586 B.n93 163.367
R960 B.n590 B.n93 163.367
R961 B.n794 B.n21 163.367
R962 B.n790 B.n21 163.367
R963 B.n790 B.n789 163.367
R964 B.n789 B.n788 163.367
R965 B.n788 B.n23 163.367
R966 B.n784 B.n23 163.367
R967 B.n784 B.n783 163.367
R968 B.n783 B.n782 163.367
R969 B.n782 B.n25 163.367
R970 B.n778 B.n25 163.367
R971 B.n778 B.n777 163.367
R972 B.n777 B.n776 163.367
R973 B.n776 B.n27 163.367
R974 B.n772 B.n27 163.367
R975 B.n772 B.n771 163.367
R976 B.n771 B.n770 163.367
R977 B.n770 B.n29 163.367
R978 B.n766 B.n29 163.367
R979 B.n766 B.n765 163.367
R980 B.n765 B.n764 163.367
R981 B.n764 B.n31 163.367
R982 B.n760 B.n31 163.367
R983 B.n760 B.n759 163.367
R984 B.n759 B.n758 163.367
R985 B.n758 B.n33 163.367
R986 B.n754 B.n33 163.367
R987 B.n754 B.n753 163.367
R988 B.n753 B.n752 163.367
R989 B.n752 B.n35 163.367
R990 B.n748 B.n35 163.367
R991 B.n748 B.n747 163.367
R992 B.n747 B.n746 163.367
R993 B.n746 B.n37 163.367
R994 B.n742 B.n37 163.367
R995 B.n742 B.n741 163.367
R996 B.n741 B.n740 163.367
R997 B.n740 B.n39 163.367
R998 B.n736 B.n39 163.367
R999 B.n736 B.n735 163.367
R1000 B.n735 B.n734 163.367
R1001 B.n734 B.n41 163.367
R1002 B.n730 B.n41 163.367
R1003 B.n730 B.n729 163.367
R1004 B.n729 B.n728 163.367
R1005 B.n728 B.n43 163.367
R1006 B.n724 B.n43 163.367
R1007 B.n724 B.n723 163.367
R1008 B.n723 B.n722 163.367
R1009 B.n722 B.n45 163.367
R1010 B.n718 B.n45 163.367
R1011 B.n718 B.n717 163.367
R1012 B.n717 B.n716 163.367
R1013 B.n716 B.n47 163.367
R1014 B.n712 B.n47 163.367
R1015 B.n712 B.n711 163.367
R1016 B.n711 B.n710 163.367
R1017 B.n710 B.n49 163.367
R1018 B.n706 B.n49 163.367
R1019 B.n706 B.n705 163.367
R1020 B.n705 B.n704 163.367
R1021 B.n704 B.n51 163.367
R1022 B.n700 B.n51 163.367
R1023 B.n700 B.n699 163.367
R1024 B.n699 B.n55 163.367
R1025 B.n695 B.n55 163.367
R1026 B.n695 B.n694 163.367
R1027 B.n694 B.n693 163.367
R1028 B.n693 B.n57 163.367
R1029 B.n689 B.n57 163.367
R1030 B.n689 B.n688 163.367
R1031 B.n688 B.n687 163.367
R1032 B.n687 B.n59 163.367
R1033 B.n682 B.n59 163.367
R1034 B.n682 B.n681 163.367
R1035 B.n681 B.n680 163.367
R1036 B.n680 B.n63 163.367
R1037 B.n676 B.n63 163.367
R1038 B.n676 B.n675 163.367
R1039 B.n675 B.n674 163.367
R1040 B.n674 B.n65 163.367
R1041 B.n670 B.n65 163.367
R1042 B.n670 B.n669 163.367
R1043 B.n669 B.n668 163.367
R1044 B.n668 B.n67 163.367
R1045 B.n664 B.n67 163.367
R1046 B.n664 B.n663 163.367
R1047 B.n663 B.n662 163.367
R1048 B.n662 B.n69 163.367
R1049 B.n658 B.n69 163.367
R1050 B.n658 B.n657 163.367
R1051 B.n657 B.n656 163.367
R1052 B.n656 B.n71 163.367
R1053 B.n652 B.n71 163.367
R1054 B.n652 B.n651 163.367
R1055 B.n651 B.n650 163.367
R1056 B.n650 B.n73 163.367
R1057 B.n646 B.n73 163.367
R1058 B.n646 B.n645 163.367
R1059 B.n645 B.n644 163.367
R1060 B.n644 B.n75 163.367
R1061 B.n640 B.n75 163.367
R1062 B.n640 B.n639 163.367
R1063 B.n639 B.n638 163.367
R1064 B.n638 B.n77 163.367
R1065 B.n634 B.n77 163.367
R1066 B.n634 B.n633 163.367
R1067 B.n633 B.n632 163.367
R1068 B.n632 B.n79 163.367
R1069 B.n628 B.n79 163.367
R1070 B.n628 B.n627 163.367
R1071 B.n627 B.n626 163.367
R1072 B.n626 B.n81 163.367
R1073 B.n622 B.n81 163.367
R1074 B.n622 B.n621 163.367
R1075 B.n621 B.n620 163.367
R1076 B.n620 B.n83 163.367
R1077 B.n616 B.n83 163.367
R1078 B.n616 B.n615 163.367
R1079 B.n615 B.n614 163.367
R1080 B.n614 B.n85 163.367
R1081 B.n610 B.n85 163.367
R1082 B.n610 B.n609 163.367
R1083 B.n609 B.n608 163.367
R1084 B.n608 B.n87 163.367
R1085 B.n604 B.n87 163.367
R1086 B.n604 B.n603 163.367
R1087 B.n603 B.n602 163.367
R1088 B.n602 B.n89 163.367
R1089 B.n598 B.n89 163.367
R1090 B.n598 B.n597 163.367
R1091 B.n597 B.n596 163.367
R1092 B.n596 B.n91 163.367
R1093 B.n592 B.n91 163.367
R1094 B.n592 B.n591 163.367
R1095 B.n162 B.t5 141.388
R1096 B.n60 B.t7 141.388
R1097 B.n168 B.t2 141.363
R1098 B.n52 B.t10 141.363
R1099 B.n163 B.t4 109.388
R1100 B.n61 B.t8 109.388
R1101 B.n169 B.t1 109.365
R1102 B.n53 B.t11 109.365
R1103 B.n383 B.n163 59.5399
R1104 B.n170 B.n169 59.5399
R1105 B.n54 B.n53 59.5399
R1106 B.n685 B.n61 59.5399
R1107 B.n589 B.n92 36.059
R1108 B.n793 B.n20 36.059
R1109 B.n479 B.n130 36.059
R1110 B.n275 B.n202 36.059
R1111 B.n163 B.n162 32.0005
R1112 B.n169 B.n168 32.0005
R1113 B.n53 B.n52 32.0005
R1114 B.n61 B.n60 32.0005
R1115 B B.n851 18.0485
R1116 B.n793 B.n792 10.6151
R1117 B.n792 B.n791 10.6151
R1118 B.n791 B.n22 10.6151
R1119 B.n787 B.n22 10.6151
R1120 B.n787 B.n786 10.6151
R1121 B.n786 B.n785 10.6151
R1122 B.n785 B.n24 10.6151
R1123 B.n781 B.n24 10.6151
R1124 B.n781 B.n780 10.6151
R1125 B.n780 B.n779 10.6151
R1126 B.n779 B.n26 10.6151
R1127 B.n775 B.n26 10.6151
R1128 B.n775 B.n774 10.6151
R1129 B.n774 B.n773 10.6151
R1130 B.n773 B.n28 10.6151
R1131 B.n769 B.n28 10.6151
R1132 B.n769 B.n768 10.6151
R1133 B.n768 B.n767 10.6151
R1134 B.n767 B.n30 10.6151
R1135 B.n763 B.n30 10.6151
R1136 B.n763 B.n762 10.6151
R1137 B.n762 B.n761 10.6151
R1138 B.n761 B.n32 10.6151
R1139 B.n757 B.n32 10.6151
R1140 B.n757 B.n756 10.6151
R1141 B.n756 B.n755 10.6151
R1142 B.n755 B.n34 10.6151
R1143 B.n751 B.n34 10.6151
R1144 B.n751 B.n750 10.6151
R1145 B.n750 B.n749 10.6151
R1146 B.n749 B.n36 10.6151
R1147 B.n745 B.n36 10.6151
R1148 B.n745 B.n744 10.6151
R1149 B.n744 B.n743 10.6151
R1150 B.n743 B.n38 10.6151
R1151 B.n739 B.n38 10.6151
R1152 B.n739 B.n738 10.6151
R1153 B.n738 B.n737 10.6151
R1154 B.n737 B.n40 10.6151
R1155 B.n733 B.n40 10.6151
R1156 B.n733 B.n732 10.6151
R1157 B.n732 B.n731 10.6151
R1158 B.n731 B.n42 10.6151
R1159 B.n727 B.n42 10.6151
R1160 B.n727 B.n726 10.6151
R1161 B.n726 B.n725 10.6151
R1162 B.n725 B.n44 10.6151
R1163 B.n721 B.n44 10.6151
R1164 B.n721 B.n720 10.6151
R1165 B.n720 B.n719 10.6151
R1166 B.n719 B.n46 10.6151
R1167 B.n715 B.n46 10.6151
R1168 B.n715 B.n714 10.6151
R1169 B.n714 B.n713 10.6151
R1170 B.n713 B.n48 10.6151
R1171 B.n709 B.n48 10.6151
R1172 B.n709 B.n708 10.6151
R1173 B.n708 B.n707 10.6151
R1174 B.n707 B.n50 10.6151
R1175 B.n703 B.n50 10.6151
R1176 B.n703 B.n702 10.6151
R1177 B.n702 B.n701 10.6151
R1178 B.n698 B.n697 10.6151
R1179 B.n697 B.n696 10.6151
R1180 B.n696 B.n56 10.6151
R1181 B.n692 B.n56 10.6151
R1182 B.n692 B.n691 10.6151
R1183 B.n691 B.n690 10.6151
R1184 B.n690 B.n58 10.6151
R1185 B.n686 B.n58 10.6151
R1186 B.n684 B.n683 10.6151
R1187 B.n683 B.n62 10.6151
R1188 B.n679 B.n62 10.6151
R1189 B.n679 B.n678 10.6151
R1190 B.n678 B.n677 10.6151
R1191 B.n677 B.n64 10.6151
R1192 B.n673 B.n64 10.6151
R1193 B.n673 B.n672 10.6151
R1194 B.n672 B.n671 10.6151
R1195 B.n671 B.n66 10.6151
R1196 B.n667 B.n66 10.6151
R1197 B.n667 B.n666 10.6151
R1198 B.n666 B.n665 10.6151
R1199 B.n665 B.n68 10.6151
R1200 B.n661 B.n68 10.6151
R1201 B.n661 B.n660 10.6151
R1202 B.n660 B.n659 10.6151
R1203 B.n659 B.n70 10.6151
R1204 B.n655 B.n70 10.6151
R1205 B.n655 B.n654 10.6151
R1206 B.n654 B.n653 10.6151
R1207 B.n653 B.n72 10.6151
R1208 B.n649 B.n72 10.6151
R1209 B.n649 B.n648 10.6151
R1210 B.n648 B.n647 10.6151
R1211 B.n647 B.n74 10.6151
R1212 B.n643 B.n74 10.6151
R1213 B.n643 B.n642 10.6151
R1214 B.n642 B.n641 10.6151
R1215 B.n641 B.n76 10.6151
R1216 B.n637 B.n76 10.6151
R1217 B.n637 B.n636 10.6151
R1218 B.n636 B.n635 10.6151
R1219 B.n635 B.n78 10.6151
R1220 B.n631 B.n78 10.6151
R1221 B.n631 B.n630 10.6151
R1222 B.n630 B.n629 10.6151
R1223 B.n629 B.n80 10.6151
R1224 B.n625 B.n80 10.6151
R1225 B.n625 B.n624 10.6151
R1226 B.n624 B.n623 10.6151
R1227 B.n623 B.n82 10.6151
R1228 B.n619 B.n82 10.6151
R1229 B.n619 B.n618 10.6151
R1230 B.n618 B.n617 10.6151
R1231 B.n617 B.n84 10.6151
R1232 B.n613 B.n84 10.6151
R1233 B.n613 B.n612 10.6151
R1234 B.n612 B.n611 10.6151
R1235 B.n611 B.n86 10.6151
R1236 B.n607 B.n86 10.6151
R1237 B.n607 B.n606 10.6151
R1238 B.n606 B.n605 10.6151
R1239 B.n605 B.n88 10.6151
R1240 B.n601 B.n88 10.6151
R1241 B.n601 B.n600 10.6151
R1242 B.n600 B.n599 10.6151
R1243 B.n599 B.n90 10.6151
R1244 B.n595 B.n90 10.6151
R1245 B.n595 B.n594 10.6151
R1246 B.n594 B.n593 10.6151
R1247 B.n593 B.n92 10.6151
R1248 B.n480 B.n479 10.6151
R1249 B.n481 B.n480 10.6151
R1250 B.n481 B.n128 10.6151
R1251 B.n485 B.n128 10.6151
R1252 B.n486 B.n485 10.6151
R1253 B.n487 B.n486 10.6151
R1254 B.n487 B.n126 10.6151
R1255 B.n491 B.n126 10.6151
R1256 B.n492 B.n491 10.6151
R1257 B.n493 B.n492 10.6151
R1258 B.n493 B.n124 10.6151
R1259 B.n497 B.n124 10.6151
R1260 B.n498 B.n497 10.6151
R1261 B.n499 B.n498 10.6151
R1262 B.n499 B.n122 10.6151
R1263 B.n503 B.n122 10.6151
R1264 B.n504 B.n503 10.6151
R1265 B.n505 B.n504 10.6151
R1266 B.n505 B.n120 10.6151
R1267 B.n509 B.n120 10.6151
R1268 B.n510 B.n509 10.6151
R1269 B.n511 B.n510 10.6151
R1270 B.n511 B.n118 10.6151
R1271 B.n515 B.n118 10.6151
R1272 B.n516 B.n515 10.6151
R1273 B.n517 B.n516 10.6151
R1274 B.n517 B.n116 10.6151
R1275 B.n521 B.n116 10.6151
R1276 B.n522 B.n521 10.6151
R1277 B.n523 B.n522 10.6151
R1278 B.n523 B.n114 10.6151
R1279 B.n527 B.n114 10.6151
R1280 B.n528 B.n527 10.6151
R1281 B.n529 B.n528 10.6151
R1282 B.n529 B.n112 10.6151
R1283 B.n533 B.n112 10.6151
R1284 B.n534 B.n533 10.6151
R1285 B.n535 B.n534 10.6151
R1286 B.n535 B.n110 10.6151
R1287 B.n539 B.n110 10.6151
R1288 B.n540 B.n539 10.6151
R1289 B.n541 B.n540 10.6151
R1290 B.n541 B.n108 10.6151
R1291 B.n545 B.n108 10.6151
R1292 B.n546 B.n545 10.6151
R1293 B.n547 B.n546 10.6151
R1294 B.n547 B.n106 10.6151
R1295 B.n551 B.n106 10.6151
R1296 B.n552 B.n551 10.6151
R1297 B.n553 B.n552 10.6151
R1298 B.n553 B.n104 10.6151
R1299 B.n557 B.n104 10.6151
R1300 B.n558 B.n557 10.6151
R1301 B.n559 B.n558 10.6151
R1302 B.n559 B.n102 10.6151
R1303 B.n563 B.n102 10.6151
R1304 B.n564 B.n563 10.6151
R1305 B.n565 B.n564 10.6151
R1306 B.n565 B.n100 10.6151
R1307 B.n569 B.n100 10.6151
R1308 B.n570 B.n569 10.6151
R1309 B.n571 B.n570 10.6151
R1310 B.n571 B.n98 10.6151
R1311 B.n575 B.n98 10.6151
R1312 B.n576 B.n575 10.6151
R1313 B.n577 B.n576 10.6151
R1314 B.n577 B.n96 10.6151
R1315 B.n581 B.n96 10.6151
R1316 B.n582 B.n581 10.6151
R1317 B.n583 B.n582 10.6151
R1318 B.n583 B.n94 10.6151
R1319 B.n587 B.n94 10.6151
R1320 B.n588 B.n587 10.6151
R1321 B.n589 B.n588 10.6151
R1322 B.n276 B.n275 10.6151
R1323 B.n277 B.n276 10.6151
R1324 B.n277 B.n200 10.6151
R1325 B.n281 B.n200 10.6151
R1326 B.n282 B.n281 10.6151
R1327 B.n283 B.n282 10.6151
R1328 B.n283 B.n198 10.6151
R1329 B.n287 B.n198 10.6151
R1330 B.n288 B.n287 10.6151
R1331 B.n289 B.n288 10.6151
R1332 B.n289 B.n196 10.6151
R1333 B.n293 B.n196 10.6151
R1334 B.n294 B.n293 10.6151
R1335 B.n295 B.n294 10.6151
R1336 B.n295 B.n194 10.6151
R1337 B.n299 B.n194 10.6151
R1338 B.n300 B.n299 10.6151
R1339 B.n301 B.n300 10.6151
R1340 B.n301 B.n192 10.6151
R1341 B.n305 B.n192 10.6151
R1342 B.n306 B.n305 10.6151
R1343 B.n307 B.n306 10.6151
R1344 B.n307 B.n190 10.6151
R1345 B.n311 B.n190 10.6151
R1346 B.n312 B.n311 10.6151
R1347 B.n313 B.n312 10.6151
R1348 B.n313 B.n188 10.6151
R1349 B.n317 B.n188 10.6151
R1350 B.n318 B.n317 10.6151
R1351 B.n319 B.n318 10.6151
R1352 B.n319 B.n186 10.6151
R1353 B.n323 B.n186 10.6151
R1354 B.n324 B.n323 10.6151
R1355 B.n325 B.n324 10.6151
R1356 B.n325 B.n184 10.6151
R1357 B.n329 B.n184 10.6151
R1358 B.n330 B.n329 10.6151
R1359 B.n331 B.n330 10.6151
R1360 B.n331 B.n182 10.6151
R1361 B.n335 B.n182 10.6151
R1362 B.n336 B.n335 10.6151
R1363 B.n337 B.n336 10.6151
R1364 B.n337 B.n180 10.6151
R1365 B.n341 B.n180 10.6151
R1366 B.n342 B.n341 10.6151
R1367 B.n343 B.n342 10.6151
R1368 B.n343 B.n178 10.6151
R1369 B.n347 B.n178 10.6151
R1370 B.n348 B.n347 10.6151
R1371 B.n349 B.n348 10.6151
R1372 B.n349 B.n176 10.6151
R1373 B.n353 B.n176 10.6151
R1374 B.n354 B.n353 10.6151
R1375 B.n355 B.n354 10.6151
R1376 B.n355 B.n174 10.6151
R1377 B.n359 B.n174 10.6151
R1378 B.n360 B.n359 10.6151
R1379 B.n361 B.n360 10.6151
R1380 B.n361 B.n172 10.6151
R1381 B.n365 B.n172 10.6151
R1382 B.n366 B.n365 10.6151
R1383 B.n367 B.n366 10.6151
R1384 B.n371 B.n370 10.6151
R1385 B.n372 B.n371 10.6151
R1386 B.n372 B.n166 10.6151
R1387 B.n376 B.n166 10.6151
R1388 B.n377 B.n376 10.6151
R1389 B.n378 B.n377 10.6151
R1390 B.n378 B.n164 10.6151
R1391 B.n382 B.n164 10.6151
R1392 B.n385 B.n384 10.6151
R1393 B.n385 B.n160 10.6151
R1394 B.n389 B.n160 10.6151
R1395 B.n390 B.n389 10.6151
R1396 B.n391 B.n390 10.6151
R1397 B.n391 B.n158 10.6151
R1398 B.n395 B.n158 10.6151
R1399 B.n396 B.n395 10.6151
R1400 B.n397 B.n396 10.6151
R1401 B.n397 B.n156 10.6151
R1402 B.n401 B.n156 10.6151
R1403 B.n402 B.n401 10.6151
R1404 B.n403 B.n402 10.6151
R1405 B.n403 B.n154 10.6151
R1406 B.n407 B.n154 10.6151
R1407 B.n408 B.n407 10.6151
R1408 B.n409 B.n408 10.6151
R1409 B.n409 B.n152 10.6151
R1410 B.n413 B.n152 10.6151
R1411 B.n414 B.n413 10.6151
R1412 B.n415 B.n414 10.6151
R1413 B.n415 B.n150 10.6151
R1414 B.n419 B.n150 10.6151
R1415 B.n420 B.n419 10.6151
R1416 B.n421 B.n420 10.6151
R1417 B.n421 B.n148 10.6151
R1418 B.n425 B.n148 10.6151
R1419 B.n426 B.n425 10.6151
R1420 B.n427 B.n426 10.6151
R1421 B.n427 B.n146 10.6151
R1422 B.n431 B.n146 10.6151
R1423 B.n432 B.n431 10.6151
R1424 B.n433 B.n432 10.6151
R1425 B.n433 B.n144 10.6151
R1426 B.n437 B.n144 10.6151
R1427 B.n438 B.n437 10.6151
R1428 B.n439 B.n438 10.6151
R1429 B.n439 B.n142 10.6151
R1430 B.n443 B.n142 10.6151
R1431 B.n444 B.n443 10.6151
R1432 B.n445 B.n444 10.6151
R1433 B.n445 B.n140 10.6151
R1434 B.n449 B.n140 10.6151
R1435 B.n450 B.n449 10.6151
R1436 B.n451 B.n450 10.6151
R1437 B.n451 B.n138 10.6151
R1438 B.n455 B.n138 10.6151
R1439 B.n456 B.n455 10.6151
R1440 B.n457 B.n456 10.6151
R1441 B.n457 B.n136 10.6151
R1442 B.n461 B.n136 10.6151
R1443 B.n462 B.n461 10.6151
R1444 B.n463 B.n462 10.6151
R1445 B.n463 B.n134 10.6151
R1446 B.n467 B.n134 10.6151
R1447 B.n468 B.n467 10.6151
R1448 B.n469 B.n468 10.6151
R1449 B.n469 B.n132 10.6151
R1450 B.n473 B.n132 10.6151
R1451 B.n474 B.n473 10.6151
R1452 B.n475 B.n474 10.6151
R1453 B.n475 B.n130 10.6151
R1454 B.n271 B.n202 10.6151
R1455 B.n271 B.n270 10.6151
R1456 B.n270 B.n269 10.6151
R1457 B.n269 B.n204 10.6151
R1458 B.n265 B.n204 10.6151
R1459 B.n265 B.n264 10.6151
R1460 B.n264 B.n263 10.6151
R1461 B.n263 B.n206 10.6151
R1462 B.n259 B.n206 10.6151
R1463 B.n259 B.n258 10.6151
R1464 B.n258 B.n257 10.6151
R1465 B.n257 B.n208 10.6151
R1466 B.n253 B.n208 10.6151
R1467 B.n253 B.n252 10.6151
R1468 B.n252 B.n251 10.6151
R1469 B.n251 B.n210 10.6151
R1470 B.n247 B.n210 10.6151
R1471 B.n247 B.n246 10.6151
R1472 B.n246 B.n245 10.6151
R1473 B.n245 B.n212 10.6151
R1474 B.n241 B.n212 10.6151
R1475 B.n241 B.n240 10.6151
R1476 B.n240 B.n239 10.6151
R1477 B.n239 B.n214 10.6151
R1478 B.n235 B.n214 10.6151
R1479 B.n235 B.n234 10.6151
R1480 B.n234 B.n233 10.6151
R1481 B.n233 B.n216 10.6151
R1482 B.n229 B.n216 10.6151
R1483 B.n229 B.n228 10.6151
R1484 B.n228 B.n227 10.6151
R1485 B.n227 B.n218 10.6151
R1486 B.n223 B.n218 10.6151
R1487 B.n223 B.n222 10.6151
R1488 B.n222 B.n221 10.6151
R1489 B.n221 B.n0 10.6151
R1490 B.n847 B.n1 10.6151
R1491 B.n847 B.n846 10.6151
R1492 B.n846 B.n845 10.6151
R1493 B.n845 B.n4 10.6151
R1494 B.n841 B.n4 10.6151
R1495 B.n841 B.n840 10.6151
R1496 B.n840 B.n839 10.6151
R1497 B.n839 B.n6 10.6151
R1498 B.n835 B.n6 10.6151
R1499 B.n835 B.n834 10.6151
R1500 B.n834 B.n833 10.6151
R1501 B.n833 B.n8 10.6151
R1502 B.n829 B.n8 10.6151
R1503 B.n829 B.n828 10.6151
R1504 B.n828 B.n827 10.6151
R1505 B.n827 B.n10 10.6151
R1506 B.n823 B.n10 10.6151
R1507 B.n823 B.n822 10.6151
R1508 B.n822 B.n821 10.6151
R1509 B.n821 B.n12 10.6151
R1510 B.n817 B.n12 10.6151
R1511 B.n817 B.n816 10.6151
R1512 B.n816 B.n815 10.6151
R1513 B.n815 B.n14 10.6151
R1514 B.n811 B.n14 10.6151
R1515 B.n811 B.n810 10.6151
R1516 B.n810 B.n809 10.6151
R1517 B.n809 B.n16 10.6151
R1518 B.n805 B.n16 10.6151
R1519 B.n805 B.n804 10.6151
R1520 B.n804 B.n803 10.6151
R1521 B.n803 B.n18 10.6151
R1522 B.n799 B.n18 10.6151
R1523 B.n799 B.n798 10.6151
R1524 B.n798 B.n797 10.6151
R1525 B.n797 B.n20 10.6151
R1526 B.n698 B.n54 6.5566
R1527 B.n686 B.n685 6.5566
R1528 B.n370 B.n170 6.5566
R1529 B.n383 B.n382 6.5566
R1530 B.n701 B.n54 4.05904
R1531 B.n685 B.n684 4.05904
R1532 B.n367 B.n170 4.05904
R1533 B.n384 B.n383 4.05904
R1534 B.n851 B.n0 2.81026
R1535 B.n851 B.n1 2.81026
C0 VDD2 VTAIL 16.1192f
C1 VDD2 VDD1 1.34572f
C2 B w_n2950_n4810# 10.4156f
C3 VP w_n2950_n4810# 6.43521f
C4 VP B 1.6743f
C5 VN w_n2950_n4810# 6.05509f
C6 VTAIL w_n2950_n4810# 4.12476f
C7 VN B 1.04216f
C8 VTAIL B 4.53988f
C9 VN VP 7.84604f
C10 VDD1 w_n2950_n4810# 2.81449f
C11 VDD2 w_n2950_n4810# 2.89155f
C12 VTAIL VP 13.7511f
C13 VDD1 B 2.51202f
C14 VDD2 B 2.58009f
C15 VTAIL VN 13.7365f
C16 VDD1 VP 14.175401f
C17 VDD2 VP 0.421198f
C18 VDD1 VN 0.150315f
C19 VDD2 VN 13.9107f
C20 VDD1 VTAIL 16.0818f
C21 VDD2 VSUBS 1.925234f
C22 VDD1 VSUBS 1.648927f
C23 VTAIL VSUBS 1.226311f
C24 VN VSUBS 6.11984f
C25 VP VSUBS 2.866852f
C26 B VSUBS 4.38909f
C27 w_n2950_n4810# VSUBS 0.173354p
C28 B.n0 VSUBS 0.005212f
C29 B.n1 VSUBS 0.005212f
C30 B.n2 VSUBS 0.008242f
C31 B.n3 VSUBS 0.008242f
C32 B.n4 VSUBS 0.008242f
C33 B.n5 VSUBS 0.008242f
C34 B.n6 VSUBS 0.008242f
C35 B.n7 VSUBS 0.008242f
C36 B.n8 VSUBS 0.008242f
C37 B.n9 VSUBS 0.008242f
C38 B.n10 VSUBS 0.008242f
C39 B.n11 VSUBS 0.008242f
C40 B.n12 VSUBS 0.008242f
C41 B.n13 VSUBS 0.008242f
C42 B.n14 VSUBS 0.008242f
C43 B.n15 VSUBS 0.008242f
C44 B.n16 VSUBS 0.008242f
C45 B.n17 VSUBS 0.008242f
C46 B.n18 VSUBS 0.008242f
C47 B.n19 VSUBS 0.008242f
C48 B.n20 VSUBS 0.020098f
C49 B.n21 VSUBS 0.008242f
C50 B.n22 VSUBS 0.008242f
C51 B.n23 VSUBS 0.008242f
C52 B.n24 VSUBS 0.008242f
C53 B.n25 VSUBS 0.008242f
C54 B.n26 VSUBS 0.008242f
C55 B.n27 VSUBS 0.008242f
C56 B.n28 VSUBS 0.008242f
C57 B.n29 VSUBS 0.008242f
C58 B.n30 VSUBS 0.008242f
C59 B.n31 VSUBS 0.008242f
C60 B.n32 VSUBS 0.008242f
C61 B.n33 VSUBS 0.008242f
C62 B.n34 VSUBS 0.008242f
C63 B.n35 VSUBS 0.008242f
C64 B.n36 VSUBS 0.008242f
C65 B.n37 VSUBS 0.008242f
C66 B.n38 VSUBS 0.008242f
C67 B.n39 VSUBS 0.008242f
C68 B.n40 VSUBS 0.008242f
C69 B.n41 VSUBS 0.008242f
C70 B.n42 VSUBS 0.008242f
C71 B.n43 VSUBS 0.008242f
C72 B.n44 VSUBS 0.008242f
C73 B.n45 VSUBS 0.008242f
C74 B.n46 VSUBS 0.008242f
C75 B.n47 VSUBS 0.008242f
C76 B.n48 VSUBS 0.008242f
C77 B.n49 VSUBS 0.008242f
C78 B.n50 VSUBS 0.008242f
C79 B.n51 VSUBS 0.008242f
C80 B.t11 VSUBS 0.766916f
C81 B.t10 VSUBS 0.78207f
C82 B.t9 VSUBS 1.25182f
C83 B.n52 VSUBS 0.321653f
C84 B.n53 VSUBS 0.078702f
C85 B.n54 VSUBS 0.019095f
C86 B.n55 VSUBS 0.008242f
C87 B.n56 VSUBS 0.008242f
C88 B.n57 VSUBS 0.008242f
C89 B.n58 VSUBS 0.008242f
C90 B.n59 VSUBS 0.008242f
C91 B.t8 VSUBS 0.766884f
C92 B.t7 VSUBS 0.782043f
C93 B.t6 VSUBS 1.25182f
C94 B.n60 VSUBS 0.32168f
C95 B.n61 VSUBS 0.078734f
C96 B.n62 VSUBS 0.008242f
C97 B.n63 VSUBS 0.008242f
C98 B.n64 VSUBS 0.008242f
C99 B.n65 VSUBS 0.008242f
C100 B.n66 VSUBS 0.008242f
C101 B.n67 VSUBS 0.008242f
C102 B.n68 VSUBS 0.008242f
C103 B.n69 VSUBS 0.008242f
C104 B.n70 VSUBS 0.008242f
C105 B.n71 VSUBS 0.008242f
C106 B.n72 VSUBS 0.008242f
C107 B.n73 VSUBS 0.008242f
C108 B.n74 VSUBS 0.008242f
C109 B.n75 VSUBS 0.008242f
C110 B.n76 VSUBS 0.008242f
C111 B.n77 VSUBS 0.008242f
C112 B.n78 VSUBS 0.008242f
C113 B.n79 VSUBS 0.008242f
C114 B.n80 VSUBS 0.008242f
C115 B.n81 VSUBS 0.008242f
C116 B.n82 VSUBS 0.008242f
C117 B.n83 VSUBS 0.008242f
C118 B.n84 VSUBS 0.008242f
C119 B.n85 VSUBS 0.008242f
C120 B.n86 VSUBS 0.008242f
C121 B.n87 VSUBS 0.008242f
C122 B.n88 VSUBS 0.008242f
C123 B.n89 VSUBS 0.008242f
C124 B.n90 VSUBS 0.008242f
C125 B.n91 VSUBS 0.008242f
C126 B.n92 VSUBS 0.020227f
C127 B.n93 VSUBS 0.008242f
C128 B.n94 VSUBS 0.008242f
C129 B.n95 VSUBS 0.008242f
C130 B.n96 VSUBS 0.008242f
C131 B.n97 VSUBS 0.008242f
C132 B.n98 VSUBS 0.008242f
C133 B.n99 VSUBS 0.008242f
C134 B.n100 VSUBS 0.008242f
C135 B.n101 VSUBS 0.008242f
C136 B.n102 VSUBS 0.008242f
C137 B.n103 VSUBS 0.008242f
C138 B.n104 VSUBS 0.008242f
C139 B.n105 VSUBS 0.008242f
C140 B.n106 VSUBS 0.008242f
C141 B.n107 VSUBS 0.008242f
C142 B.n108 VSUBS 0.008242f
C143 B.n109 VSUBS 0.008242f
C144 B.n110 VSUBS 0.008242f
C145 B.n111 VSUBS 0.008242f
C146 B.n112 VSUBS 0.008242f
C147 B.n113 VSUBS 0.008242f
C148 B.n114 VSUBS 0.008242f
C149 B.n115 VSUBS 0.008242f
C150 B.n116 VSUBS 0.008242f
C151 B.n117 VSUBS 0.008242f
C152 B.n118 VSUBS 0.008242f
C153 B.n119 VSUBS 0.008242f
C154 B.n120 VSUBS 0.008242f
C155 B.n121 VSUBS 0.008242f
C156 B.n122 VSUBS 0.008242f
C157 B.n123 VSUBS 0.008242f
C158 B.n124 VSUBS 0.008242f
C159 B.n125 VSUBS 0.008242f
C160 B.n126 VSUBS 0.008242f
C161 B.n127 VSUBS 0.008242f
C162 B.n128 VSUBS 0.008242f
C163 B.n129 VSUBS 0.008242f
C164 B.n130 VSUBS 0.021109f
C165 B.n131 VSUBS 0.008242f
C166 B.n132 VSUBS 0.008242f
C167 B.n133 VSUBS 0.008242f
C168 B.n134 VSUBS 0.008242f
C169 B.n135 VSUBS 0.008242f
C170 B.n136 VSUBS 0.008242f
C171 B.n137 VSUBS 0.008242f
C172 B.n138 VSUBS 0.008242f
C173 B.n139 VSUBS 0.008242f
C174 B.n140 VSUBS 0.008242f
C175 B.n141 VSUBS 0.008242f
C176 B.n142 VSUBS 0.008242f
C177 B.n143 VSUBS 0.008242f
C178 B.n144 VSUBS 0.008242f
C179 B.n145 VSUBS 0.008242f
C180 B.n146 VSUBS 0.008242f
C181 B.n147 VSUBS 0.008242f
C182 B.n148 VSUBS 0.008242f
C183 B.n149 VSUBS 0.008242f
C184 B.n150 VSUBS 0.008242f
C185 B.n151 VSUBS 0.008242f
C186 B.n152 VSUBS 0.008242f
C187 B.n153 VSUBS 0.008242f
C188 B.n154 VSUBS 0.008242f
C189 B.n155 VSUBS 0.008242f
C190 B.n156 VSUBS 0.008242f
C191 B.n157 VSUBS 0.008242f
C192 B.n158 VSUBS 0.008242f
C193 B.n159 VSUBS 0.008242f
C194 B.n160 VSUBS 0.008242f
C195 B.n161 VSUBS 0.008242f
C196 B.t4 VSUBS 0.766884f
C197 B.t5 VSUBS 0.782043f
C198 B.t3 VSUBS 1.25182f
C199 B.n162 VSUBS 0.32168f
C200 B.n163 VSUBS 0.078734f
C201 B.n164 VSUBS 0.008242f
C202 B.n165 VSUBS 0.008242f
C203 B.n166 VSUBS 0.008242f
C204 B.n167 VSUBS 0.008242f
C205 B.t1 VSUBS 0.766916f
C206 B.t2 VSUBS 0.78207f
C207 B.t0 VSUBS 1.25182f
C208 B.n168 VSUBS 0.321653f
C209 B.n169 VSUBS 0.078702f
C210 B.n170 VSUBS 0.019095f
C211 B.n171 VSUBS 0.008242f
C212 B.n172 VSUBS 0.008242f
C213 B.n173 VSUBS 0.008242f
C214 B.n174 VSUBS 0.008242f
C215 B.n175 VSUBS 0.008242f
C216 B.n176 VSUBS 0.008242f
C217 B.n177 VSUBS 0.008242f
C218 B.n178 VSUBS 0.008242f
C219 B.n179 VSUBS 0.008242f
C220 B.n180 VSUBS 0.008242f
C221 B.n181 VSUBS 0.008242f
C222 B.n182 VSUBS 0.008242f
C223 B.n183 VSUBS 0.008242f
C224 B.n184 VSUBS 0.008242f
C225 B.n185 VSUBS 0.008242f
C226 B.n186 VSUBS 0.008242f
C227 B.n187 VSUBS 0.008242f
C228 B.n188 VSUBS 0.008242f
C229 B.n189 VSUBS 0.008242f
C230 B.n190 VSUBS 0.008242f
C231 B.n191 VSUBS 0.008242f
C232 B.n192 VSUBS 0.008242f
C233 B.n193 VSUBS 0.008242f
C234 B.n194 VSUBS 0.008242f
C235 B.n195 VSUBS 0.008242f
C236 B.n196 VSUBS 0.008242f
C237 B.n197 VSUBS 0.008242f
C238 B.n198 VSUBS 0.008242f
C239 B.n199 VSUBS 0.008242f
C240 B.n200 VSUBS 0.008242f
C241 B.n201 VSUBS 0.008242f
C242 B.n202 VSUBS 0.020098f
C243 B.n203 VSUBS 0.008242f
C244 B.n204 VSUBS 0.008242f
C245 B.n205 VSUBS 0.008242f
C246 B.n206 VSUBS 0.008242f
C247 B.n207 VSUBS 0.008242f
C248 B.n208 VSUBS 0.008242f
C249 B.n209 VSUBS 0.008242f
C250 B.n210 VSUBS 0.008242f
C251 B.n211 VSUBS 0.008242f
C252 B.n212 VSUBS 0.008242f
C253 B.n213 VSUBS 0.008242f
C254 B.n214 VSUBS 0.008242f
C255 B.n215 VSUBS 0.008242f
C256 B.n216 VSUBS 0.008242f
C257 B.n217 VSUBS 0.008242f
C258 B.n218 VSUBS 0.008242f
C259 B.n219 VSUBS 0.008242f
C260 B.n220 VSUBS 0.008242f
C261 B.n221 VSUBS 0.008242f
C262 B.n222 VSUBS 0.008242f
C263 B.n223 VSUBS 0.008242f
C264 B.n224 VSUBS 0.008242f
C265 B.n225 VSUBS 0.008242f
C266 B.n226 VSUBS 0.008242f
C267 B.n227 VSUBS 0.008242f
C268 B.n228 VSUBS 0.008242f
C269 B.n229 VSUBS 0.008242f
C270 B.n230 VSUBS 0.008242f
C271 B.n231 VSUBS 0.008242f
C272 B.n232 VSUBS 0.008242f
C273 B.n233 VSUBS 0.008242f
C274 B.n234 VSUBS 0.008242f
C275 B.n235 VSUBS 0.008242f
C276 B.n236 VSUBS 0.008242f
C277 B.n237 VSUBS 0.008242f
C278 B.n238 VSUBS 0.008242f
C279 B.n239 VSUBS 0.008242f
C280 B.n240 VSUBS 0.008242f
C281 B.n241 VSUBS 0.008242f
C282 B.n242 VSUBS 0.008242f
C283 B.n243 VSUBS 0.008242f
C284 B.n244 VSUBS 0.008242f
C285 B.n245 VSUBS 0.008242f
C286 B.n246 VSUBS 0.008242f
C287 B.n247 VSUBS 0.008242f
C288 B.n248 VSUBS 0.008242f
C289 B.n249 VSUBS 0.008242f
C290 B.n250 VSUBS 0.008242f
C291 B.n251 VSUBS 0.008242f
C292 B.n252 VSUBS 0.008242f
C293 B.n253 VSUBS 0.008242f
C294 B.n254 VSUBS 0.008242f
C295 B.n255 VSUBS 0.008242f
C296 B.n256 VSUBS 0.008242f
C297 B.n257 VSUBS 0.008242f
C298 B.n258 VSUBS 0.008242f
C299 B.n259 VSUBS 0.008242f
C300 B.n260 VSUBS 0.008242f
C301 B.n261 VSUBS 0.008242f
C302 B.n262 VSUBS 0.008242f
C303 B.n263 VSUBS 0.008242f
C304 B.n264 VSUBS 0.008242f
C305 B.n265 VSUBS 0.008242f
C306 B.n266 VSUBS 0.008242f
C307 B.n267 VSUBS 0.008242f
C308 B.n268 VSUBS 0.008242f
C309 B.n269 VSUBS 0.008242f
C310 B.n270 VSUBS 0.008242f
C311 B.n271 VSUBS 0.008242f
C312 B.n272 VSUBS 0.008242f
C313 B.n273 VSUBS 0.020098f
C314 B.n274 VSUBS 0.021109f
C315 B.n275 VSUBS 0.021109f
C316 B.n276 VSUBS 0.008242f
C317 B.n277 VSUBS 0.008242f
C318 B.n278 VSUBS 0.008242f
C319 B.n279 VSUBS 0.008242f
C320 B.n280 VSUBS 0.008242f
C321 B.n281 VSUBS 0.008242f
C322 B.n282 VSUBS 0.008242f
C323 B.n283 VSUBS 0.008242f
C324 B.n284 VSUBS 0.008242f
C325 B.n285 VSUBS 0.008242f
C326 B.n286 VSUBS 0.008242f
C327 B.n287 VSUBS 0.008242f
C328 B.n288 VSUBS 0.008242f
C329 B.n289 VSUBS 0.008242f
C330 B.n290 VSUBS 0.008242f
C331 B.n291 VSUBS 0.008242f
C332 B.n292 VSUBS 0.008242f
C333 B.n293 VSUBS 0.008242f
C334 B.n294 VSUBS 0.008242f
C335 B.n295 VSUBS 0.008242f
C336 B.n296 VSUBS 0.008242f
C337 B.n297 VSUBS 0.008242f
C338 B.n298 VSUBS 0.008242f
C339 B.n299 VSUBS 0.008242f
C340 B.n300 VSUBS 0.008242f
C341 B.n301 VSUBS 0.008242f
C342 B.n302 VSUBS 0.008242f
C343 B.n303 VSUBS 0.008242f
C344 B.n304 VSUBS 0.008242f
C345 B.n305 VSUBS 0.008242f
C346 B.n306 VSUBS 0.008242f
C347 B.n307 VSUBS 0.008242f
C348 B.n308 VSUBS 0.008242f
C349 B.n309 VSUBS 0.008242f
C350 B.n310 VSUBS 0.008242f
C351 B.n311 VSUBS 0.008242f
C352 B.n312 VSUBS 0.008242f
C353 B.n313 VSUBS 0.008242f
C354 B.n314 VSUBS 0.008242f
C355 B.n315 VSUBS 0.008242f
C356 B.n316 VSUBS 0.008242f
C357 B.n317 VSUBS 0.008242f
C358 B.n318 VSUBS 0.008242f
C359 B.n319 VSUBS 0.008242f
C360 B.n320 VSUBS 0.008242f
C361 B.n321 VSUBS 0.008242f
C362 B.n322 VSUBS 0.008242f
C363 B.n323 VSUBS 0.008242f
C364 B.n324 VSUBS 0.008242f
C365 B.n325 VSUBS 0.008242f
C366 B.n326 VSUBS 0.008242f
C367 B.n327 VSUBS 0.008242f
C368 B.n328 VSUBS 0.008242f
C369 B.n329 VSUBS 0.008242f
C370 B.n330 VSUBS 0.008242f
C371 B.n331 VSUBS 0.008242f
C372 B.n332 VSUBS 0.008242f
C373 B.n333 VSUBS 0.008242f
C374 B.n334 VSUBS 0.008242f
C375 B.n335 VSUBS 0.008242f
C376 B.n336 VSUBS 0.008242f
C377 B.n337 VSUBS 0.008242f
C378 B.n338 VSUBS 0.008242f
C379 B.n339 VSUBS 0.008242f
C380 B.n340 VSUBS 0.008242f
C381 B.n341 VSUBS 0.008242f
C382 B.n342 VSUBS 0.008242f
C383 B.n343 VSUBS 0.008242f
C384 B.n344 VSUBS 0.008242f
C385 B.n345 VSUBS 0.008242f
C386 B.n346 VSUBS 0.008242f
C387 B.n347 VSUBS 0.008242f
C388 B.n348 VSUBS 0.008242f
C389 B.n349 VSUBS 0.008242f
C390 B.n350 VSUBS 0.008242f
C391 B.n351 VSUBS 0.008242f
C392 B.n352 VSUBS 0.008242f
C393 B.n353 VSUBS 0.008242f
C394 B.n354 VSUBS 0.008242f
C395 B.n355 VSUBS 0.008242f
C396 B.n356 VSUBS 0.008242f
C397 B.n357 VSUBS 0.008242f
C398 B.n358 VSUBS 0.008242f
C399 B.n359 VSUBS 0.008242f
C400 B.n360 VSUBS 0.008242f
C401 B.n361 VSUBS 0.008242f
C402 B.n362 VSUBS 0.008242f
C403 B.n363 VSUBS 0.008242f
C404 B.n364 VSUBS 0.008242f
C405 B.n365 VSUBS 0.008242f
C406 B.n366 VSUBS 0.008242f
C407 B.n367 VSUBS 0.005696f
C408 B.n368 VSUBS 0.008242f
C409 B.n369 VSUBS 0.008242f
C410 B.n370 VSUBS 0.006666f
C411 B.n371 VSUBS 0.008242f
C412 B.n372 VSUBS 0.008242f
C413 B.n373 VSUBS 0.008242f
C414 B.n374 VSUBS 0.008242f
C415 B.n375 VSUBS 0.008242f
C416 B.n376 VSUBS 0.008242f
C417 B.n377 VSUBS 0.008242f
C418 B.n378 VSUBS 0.008242f
C419 B.n379 VSUBS 0.008242f
C420 B.n380 VSUBS 0.008242f
C421 B.n381 VSUBS 0.008242f
C422 B.n382 VSUBS 0.006666f
C423 B.n383 VSUBS 0.019095f
C424 B.n384 VSUBS 0.005696f
C425 B.n385 VSUBS 0.008242f
C426 B.n386 VSUBS 0.008242f
C427 B.n387 VSUBS 0.008242f
C428 B.n388 VSUBS 0.008242f
C429 B.n389 VSUBS 0.008242f
C430 B.n390 VSUBS 0.008242f
C431 B.n391 VSUBS 0.008242f
C432 B.n392 VSUBS 0.008242f
C433 B.n393 VSUBS 0.008242f
C434 B.n394 VSUBS 0.008242f
C435 B.n395 VSUBS 0.008242f
C436 B.n396 VSUBS 0.008242f
C437 B.n397 VSUBS 0.008242f
C438 B.n398 VSUBS 0.008242f
C439 B.n399 VSUBS 0.008242f
C440 B.n400 VSUBS 0.008242f
C441 B.n401 VSUBS 0.008242f
C442 B.n402 VSUBS 0.008242f
C443 B.n403 VSUBS 0.008242f
C444 B.n404 VSUBS 0.008242f
C445 B.n405 VSUBS 0.008242f
C446 B.n406 VSUBS 0.008242f
C447 B.n407 VSUBS 0.008242f
C448 B.n408 VSUBS 0.008242f
C449 B.n409 VSUBS 0.008242f
C450 B.n410 VSUBS 0.008242f
C451 B.n411 VSUBS 0.008242f
C452 B.n412 VSUBS 0.008242f
C453 B.n413 VSUBS 0.008242f
C454 B.n414 VSUBS 0.008242f
C455 B.n415 VSUBS 0.008242f
C456 B.n416 VSUBS 0.008242f
C457 B.n417 VSUBS 0.008242f
C458 B.n418 VSUBS 0.008242f
C459 B.n419 VSUBS 0.008242f
C460 B.n420 VSUBS 0.008242f
C461 B.n421 VSUBS 0.008242f
C462 B.n422 VSUBS 0.008242f
C463 B.n423 VSUBS 0.008242f
C464 B.n424 VSUBS 0.008242f
C465 B.n425 VSUBS 0.008242f
C466 B.n426 VSUBS 0.008242f
C467 B.n427 VSUBS 0.008242f
C468 B.n428 VSUBS 0.008242f
C469 B.n429 VSUBS 0.008242f
C470 B.n430 VSUBS 0.008242f
C471 B.n431 VSUBS 0.008242f
C472 B.n432 VSUBS 0.008242f
C473 B.n433 VSUBS 0.008242f
C474 B.n434 VSUBS 0.008242f
C475 B.n435 VSUBS 0.008242f
C476 B.n436 VSUBS 0.008242f
C477 B.n437 VSUBS 0.008242f
C478 B.n438 VSUBS 0.008242f
C479 B.n439 VSUBS 0.008242f
C480 B.n440 VSUBS 0.008242f
C481 B.n441 VSUBS 0.008242f
C482 B.n442 VSUBS 0.008242f
C483 B.n443 VSUBS 0.008242f
C484 B.n444 VSUBS 0.008242f
C485 B.n445 VSUBS 0.008242f
C486 B.n446 VSUBS 0.008242f
C487 B.n447 VSUBS 0.008242f
C488 B.n448 VSUBS 0.008242f
C489 B.n449 VSUBS 0.008242f
C490 B.n450 VSUBS 0.008242f
C491 B.n451 VSUBS 0.008242f
C492 B.n452 VSUBS 0.008242f
C493 B.n453 VSUBS 0.008242f
C494 B.n454 VSUBS 0.008242f
C495 B.n455 VSUBS 0.008242f
C496 B.n456 VSUBS 0.008242f
C497 B.n457 VSUBS 0.008242f
C498 B.n458 VSUBS 0.008242f
C499 B.n459 VSUBS 0.008242f
C500 B.n460 VSUBS 0.008242f
C501 B.n461 VSUBS 0.008242f
C502 B.n462 VSUBS 0.008242f
C503 B.n463 VSUBS 0.008242f
C504 B.n464 VSUBS 0.008242f
C505 B.n465 VSUBS 0.008242f
C506 B.n466 VSUBS 0.008242f
C507 B.n467 VSUBS 0.008242f
C508 B.n468 VSUBS 0.008242f
C509 B.n469 VSUBS 0.008242f
C510 B.n470 VSUBS 0.008242f
C511 B.n471 VSUBS 0.008242f
C512 B.n472 VSUBS 0.008242f
C513 B.n473 VSUBS 0.008242f
C514 B.n474 VSUBS 0.008242f
C515 B.n475 VSUBS 0.008242f
C516 B.n476 VSUBS 0.008242f
C517 B.n477 VSUBS 0.021109f
C518 B.n478 VSUBS 0.020098f
C519 B.n479 VSUBS 0.020098f
C520 B.n480 VSUBS 0.008242f
C521 B.n481 VSUBS 0.008242f
C522 B.n482 VSUBS 0.008242f
C523 B.n483 VSUBS 0.008242f
C524 B.n484 VSUBS 0.008242f
C525 B.n485 VSUBS 0.008242f
C526 B.n486 VSUBS 0.008242f
C527 B.n487 VSUBS 0.008242f
C528 B.n488 VSUBS 0.008242f
C529 B.n489 VSUBS 0.008242f
C530 B.n490 VSUBS 0.008242f
C531 B.n491 VSUBS 0.008242f
C532 B.n492 VSUBS 0.008242f
C533 B.n493 VSUBS 0.008242f
C534 B.n494 VSUBS 0.008242f
C535 B.n495 VSUBS 0.008242f
C536 B.n496 VSUBS 0.008242f
C537 B.n497 VSUBS 0.008242f
C538 B.n498 VSUBS 0.008242f
C539 B.n499 VSUBS 0.008242f
C540 B.n500 VSUBS 0.008242f
C541 B.n501 VSUBS 0.008242f
C542 B.n502 VSUBS 0.008242f
C543 B.n503 VSUBS 0.008242f
C544 B.n504 VSUBS 0.008242f
C545 B.n505 VSUBS 0.008242f
C546 B.n506 VSUBS 0.008242f
C547 B.n507 VSUBS 0.008242f
C548 B.n508 VSUBS 0.008242f
C549 B.n509 VSUBS 0.008242f
C550 B.n510 VSUBS 0.008242f
C551 B.n511 VSUBS 0.008242f
C552 B.n512 VSUBS 0.008242f
C553 B.n513 VSUBS 0.008242f
C554 B.n514 VSUBS 0.008242f
C555 B.n515 VSUBS 0.008242f
C556 B.n516 VSUBS 0.008242f
C557 B.n517 VSUBS 0.008242f
C558 B.n518 VSUBS 0.008242f
C559 B.n519 VSUBS 0.008242f
C560 B.n520 VSUBS 0.008242f
C561 B.n521 VSUBS 0.008242f
C562 B.n522 VSUBS 0.008242f
C563 B.n523 VSUBS 0.008242f
C564 B.n524 VSUBS 0.008242f
C565 B.n525 VSUBS 0.008242f
C566 B.n526 VSUBS 0.008242f
C567 B.n527 VSUBS 0.008242f
C568 B.n528 VSUBS 0.008242f
C569 B.n529 VSUBS 0.008242f
C570 B.n530 VSUBS 0.008242f
C571 B.n531 VSUBS 0.008242f
C572 B.n532 VSUBS 0.008242f
C573 B.n533 VSUBS 0.008242f
C574 B.n534 VSUBS 0.008242f
C575 B.n535 VSUBS 0.008242f
C576 B.n536 VSUBS 0.008242f
C577 B.n537 VSUBS 0.008242f
C578 B.n538 VSUBS 0.008242f
C579 B.n539 VSUBS 0.008242f
C580 B.n540 VSUBS 0.008242f
C581 B.n541 VSUBS 0.008242f
C582 B.n542 VSUBS 0.008242f
C583 B.n543 VSUBS 0.008242f
C584 B.n544 VSUBS 0.008242f
C585 B.n545 VSUBS 0.008242f
C586 B.n546 VSUBS 0.008242f
C587 B.n547 VSUBS 0.008242f
C588 B.n548 VSUBS 0.008242f
C589 B.n549 VSUBS 0.008242f
C590 B.n550 VSUBS 0.008242f
C591 B.n551 VSUBS 0.008242f
C592 B.n552 VSUBS 0.008242f
C593 B.n553 VSUBS 0.008242f
C594 B.n554 VSUBS 0.008242f
C595 B.n555 VSUBS 0.008242f
C596 B.n556 VSUBS 0.008242f
C597 B.n557 VSUBS 0.008242f
C598 B.n558 VSUBS 0.008242f
C599 B.n559 VSUBS 0.008242f
C600 B.n560 VSUBS 0.008242f
C601 B.n561 VSUBS 0.008242f
C602 B.n562 VSUBS 0.008242f
C603 B.n563 VSUBS 0.008242f
C604 B.n564 VSUBS 0.008242f
C605 B.n565 VSUBS 0.008242f
C606 B.n566 VSUBS 0.008242f
C607 B.n567 VSUBS 0.008242f
C608 B.n568 VSUBS 0.008242f
C609 B.n569 VSUBS 0.008242f
C610 B.n570 VSUBS 0.008242f
C611 B.n571 VSUBS 0.008242f
C612 B.n572 VSUBS 0.008242f
C613 B.n573 VSUBS 0.008242f
C614 B.n574 VSUBS 0.008242f
C615 B.n575 VSUBS 0.008242f
C616 B.n576 VSUBS 0.008242f
C617 B.n577 VSUBS 0.008242f
C618 B.n578 VSUBS 0.008242f
C619 B.n579 VSUBS 0.008242f
C620 B.n580 VSUBS 0.008242f
C621 B.n581 VSUBS 0.008242f
C622 B.n582 VSUBS 0.008242f
C623 B.n583 VSUBS 0.008242f
C624 B.n584 VSUBS 0.008242f
C625 B.n585 VSUBS 0.008242f
C626 B.n586 VSUBS 0.008242f
C627 B.n587 VSUBS 0.008242f
C628 B.n588 VSUBS 0.008242f
C629 B.n589 VSUBS 0.02098f
C630 B.n590 VSUBS 0.020098f
C631 B.n591 VSUBS 0.021109f
C632 B.n592 VSUBS 0.008242f
C633 B.n593 VSUBS 0.008242f
C634 B.n594 VSUBS 0.008242f
C635 B.n595 VSUBS 0.008242f
C636 B.n596 VSUBS 0.008242f
C637 B.n597 VSUBS 0.008242f
C638 B.n598 VSUBS 0.008242f
C639 B.n599 VSUBS 0.008242f
C640 B.n600 VSUBS 0.008242f
C641 B.n601 VSUBS 0.008242f
C642 B.n602 VSUBS 0.008242f
C643 B.n603 VSUBS 0.008242f
C644 B.n604 VSUBS 0.008242f
C645 B.n605 VSUBS 0.008242f
C646 B.n606 VSUBS 0.008242f
C647 B.n607 VSUBS 0.008242f
C648 B.n608 VSUBS 0.008242f
C649 B.n609 VSUBS 0.008242f
C650 B.n610 VSUBS 0.008242f
C651 B.n611 VSUBS 0.008242f
C652 B.n612 VSUBS 0.008242f
C653 B.n613 VSUBS 0.008242f
C654 B.n614 VSUBS 0.008242f
C655 B.n615 VSUBS 0.008242f
C656 B.n616 VSUBS 0.008242f
C657 B.n617 VSUBS 0.008242f
C658 B.n618 VSUBS 0.008242f
C659 B.n619 VSUBS 0.008242f
C660 B.n620 VSUBS 0.008242f
C661 B.n621 VSUBS 0.008242f
C662 B.n622 VSUBS 0.008242f
C663 B.n623 VSUBS 0.008242f
C664 B.n624 VSUBS 0.008242f
C665 B.n625 VSUBS 0.008242f
C666 B.n626 VSUBS 0.008242f
C667 B.n627 VSUBS 0.008242f
C668 B.n628 VSUBS 0.008242f
C669 B.n629 VSUBS 0.008242f
C670 B.n630 VSUBS 0.008242f
C671 B.n631 VSUBS 0.008242f
C672 B.n632 VSUBS 0.008242f
C673 B.n633 VSUBS 0.008242f
C674 B.n634 VSUBS 0.008242f
C675 B.n635 VSUBS 0.008242f
C676 B.n636 VSUBS 0.008242f
C677 B.n637 VSUBS 0.008242f
C678 B.n638 VSUBS 0.008242f
C679 B.n639 VSUBS 0.008242f
C680 B.n640 VSUBS 0.008242f
C681 B.n641 VSUBS 0.008242f
C682 B.n642 VSUBS 0.008242f
C683 B.n643 VSUBS 0.008242f
C684 B.n644 VSUBS 0.008242f
C685 B.n645 VSUBS 0.008242f
C686 B.n646 VSUBS 0.008242f
C687 B.n647 VSUBS 0.008242f
C688 B.n648 VSUBS 0.008242f
C689 B.n649 VSUBS 0.008242f
C690 B.n650 VSUBS 0.008242f
C691 B.n651 VSUBS 0.008242f
C692 B.n652 VSUBS 0.008242f
C693 B.n653 VSUBS 0.008242f
C694 B.n654 VSUBS 0.008242f
C695 B.n655 VSUBS 0.008242f
C696 B.n656 VSUBS 0.008242f
C697 B.n657 VSUBS 0.008242f
C698 B.n658 VSUBS 0.008242f
C699 B.n659 VSUBS 0.008242f
C700 B.n660 VSUBS 0.008242f
C701 B.n661 VSUBS 0.008242f
C702 B.n662 VSUBS 0.008242f
C703 B.n663 VSUBS 0.008242f
C704 B.n664 VSUBS 0.008242f
C705 B.n665 VSUBS 0.008242f
C706 B.n666 VSUBS 0.008242f
C707 B.n667 VSUBS 0.008242f
C708 B.n668 VSUBS 0.008242f
C709 B.n669 VSUBS 0.008242f
C710 B.n670 VSUBS 0.008242f
C711 B.n671 VSUBS 0.008242f
C712 B.n672 VSUBS 0.008242f
C713 B.n673 VSUBS 0.008242f
C714 B.n674 VSUBS 0.008242f
C715 B.n675 VSUBS 0.008242f
C716 B.n676 VSUBS 0.008242f
C717 B.n677 VSUBS 0.008242f
C718 B.n678 VSUBS 0.008242f
C719 B.n679 VSUBS 0.008242f
C720 B.n680 VSUBS 0.008242f
C721 B.n681 VSUBS 0.008242f
C722 B.n682 VSUBS 0.008242f
C723 B.n683 VSUBS 0.008242f
C724 B.n684 VSUBS 0.005696f
C725 B.n685 VSUBS 0.019095f
C726 B.n686 VSUBS 0.006666f
C727 B.n687 VSUBS 0.008242f
C728 B.n688 VSUBS 0.008242f
C729 B.n689 VSUBS 0.008242f
C730 B.n690 VSUBS 0.008242f
C731 B.n691 VSUBS 0.008242f
C732 B.n692 VSUBS 0.008242f
C733 B.n693 VSUBS 0.008242f
C734 B.n694 VSUBS 0.008242f
C735 B.n695 VSUBS 0.008242f
C736 B.n696 VSUBS 0.008242f
C737 B.n697 VSUBS 0.008242f
C738 B.n698 VSUBS 0.006666f
C739 B.n699 VSUBS 0.008242f
C740 B.n700 VSUBS 0.008242f
C741 B.n701 VSUBS 0.005696f
C742 B.n702 VSUBS 0.008242f
C743 B.n703 VSUBS 0.008242f
C744 B.n704 VSUBS 0.008242f
C745 B.n705 VSUBS 0.008242f
C746 B.n706 VSUBS 0.008242f
C747 B.n707 VSUBS 0.008242f
C748 B.n708 VSUBS 0.008242f
C749 B.n709 VSUBS 0.008242f
C750 B.n710 VSUBS 0.008242f
C751 B.n711 VSUBS 0.008242f
C752 B.n712 VSUBS 0.008242f
C753 B.n713 VSUBS 0.008242f
C754 B.n714 VSUBS 0.008242f
C755 B.n715 VSUBS 0.008242f
C756 B.n716 VSUBS 0.008242f
C757 B.n717 VSUBS 0.008242f
C758 B.n718 VSUBS 0.008242f
C759 B.n719 VSUBS 0.008242f
C760 B.n720 VSUBS 0.008242f
C761 B.n721 VSUBS 0.008242f
C762 B.n722 VSUBS 0.008242f
C763 B.n723 VSUBS 0.008242f
C764 B.n724 VSUBS 0.008242f
C765 B.n725 VSUBS 0.008242f
C766 B.n726 VSUBS 0.008242f
C767 B.n727 VSUBS 0.008242f
C768 B.n728 VSUBS 0.008242f
C769 B.n729 VSUBS 0.008242f
C770 B.n730 VSUBS 0.008242f
C771 B.n731 VSUBS 0.008242f
C772 B.n732 VSUBS 0.008242f
C773 B.n733 VSUBS 0.008242f
C774 B.n734 VSUBS 0.008242f
C775 B.n735 VSUBS 0.008242f
C776 B.n736 VSUBS 0.008242f
C777 B.n737 VSUBS 0.008242f
C778 B.n738 VSUBS 0.008242f
C779 B.n739 VSUBS 0.008242f
C780 B.n740 VSUBS 0.008242f
C781 B.n741 VSUBS 0.008242f
C782 B.n742 VSUBS 0.008242f
C783 B.n743 VSUBS 0.008242f
C784 B.n744 VSUBS 0.008242f
C785 B.n745 VSUBS 0.008242f
C786 B.n746 VSUBS 0.008242f
C787 B.n747 VSUBS 0.008242f
C788 B.n748 VSUBS 0.008242f
C789 B.n749 VSUBS 0.008242f
C790 B.n750 VSUBS 0.008242f
C791 B.n751 VSUBS 0.008242f
C792 B.n752 VSUBS 0.008242f
C793 B.n753 VSUBS 0.008242f
C794 B.n754 VSUBS 0.008242f
C795 B.n755 VSUBS 0.008242f
C796 B.n756 VSUBS 0.008242f
C797 B.n757 VSUBS 0.008242f
C798 B.n758 VSUBS 0.008242f
C799 B.n759 VSUBS 0.008242f
C800 B.n760 VSUBS 0.008242f
C801 B.n761 VSUBS 0.008242f
C802 B.n762 VSUBS 0.008242f
C803 B.n763 VSUBS 0.008242f
C804 B.n764 VSUBS 0.008242f
C805 B.n765 VSUBS 0.008242f
C806 B.n766 VSUBS 0.008242f
C807 B.n767 VSUBS 0.008242f
C808 B.n768 VSUBS 0.008242f
C809 B.n769 VSUBS 0.008242f
C810 B.n770 VSUBS 0.008242f
C811 B.n771 VSUBS 0.008242f
C812 B.n772 VSUBS 0.008242f
C813 B.n773 VSUBS 0.008242f
C814 B.n774 VSUBS 0.008242f
C815 B.n775 VSUBS 0.008242f
C816 B.n776 VSUBS 0.008242f
C817 B.n777 VSUBS 0.008242f
C818 B.n778 VSUBS 0.008242f
C819 B.n779 VSUBS 0.008242f
C820 B.n780 VSUBS 0.008242f
C821 B.n781 VSUBS 0.008242f
C822 B.n782 VSUBS 0.008242f
C823 B.n783 VSUBS 0.008242f
C824 B.n784 VSUBS 0.008242f
C825 B.n785 VSUBS 0.008242f
C826 B.n786 VSUBS 0.008242f
C827 B.n787 VSUBS 0.008242f
C828 B.n788 VSUBS 0.008242f
C829 B.n789 VSUBS 0.008242f
C830 B.n790 VSUBS 0.008242f
C831 B.n791 VSUBS 0.008242f
C832 B.n792 VSUBS 0.008242f
C833 B.n793 VSUBS 0.021109f
C834 B.n794 VSUBS 0.021109f
C835 B.n795 VSUBS 0.020098f
C836 B.n796 VSUBS 0.008242f
C837 B.n797 VSUBS 0.008242f
C838 B.n798 VSUBS 0.008242f
C839 B.n799 VSUBS 0.008242f
C840 B.n800 VSUBS 0.008242f
C841 B.n801 VSUBS 0.008242f
C842 B.n802 VSUBS 0.008242f
C843 B.n803 VSUBS 0.008242f
C844 B.n804 VSUBS 0.008242f
C845 B.n805 VSUBS 0.008242f
C846 B.n806 VSUBS 0.008242f
C847 B.n807 VSUBS 0.008242f
C848 B.n808 VSUBS 0.008242f
C849 B.n809 VSUBS 0.008242f
C850 B.n810 VSUBS 0.008242f
C851 B.n811 VSUBS 0.008242f
C852 B.n812 VSUBS 0.008242f
C853 B.n813 VSUBS 0.008242f
C854 B.n814 VSUBS 0.008242f
C855 B.n815 VSUBS 0.008242f
C856 B.n816 VSUBS 0.008242f
C857 B.n817 VSUBS 0.008242f
C858 B.n818 VSUBS 0.008242f
C859 B.n819 VSUBS 0.008242f
C860 B.n820 VSUBS 0.008242f
C861 B.n821 VSUBS 0.008242f
C862 B.n822 VSUBS 0.008242f
C863 B.n823 VSUBS 0.008242f
C864 B.n824 VSUBS 0.008242f
C865 B.n825 VSUBS 0.008242f
C866 B.n826 VSUBS 0.008242f
C867 B.n827 VSUBS 0.008242f
C868 B.n828 VSUBS 0.008242f
C869 B.n829 VSUBS 0.008242f
C870 B.n830 VSUBS 0.008242f
C871 B.n831 VSUBS 0.008242f
C872 B.n832 VSUBS 0.008242f
C873 B.n833 VSUBS 0.008242f
C874 B.n834 VSUBS 0.008242f
C875 B.n835 VSUBS 0.008242f
C876 B.n836 VSUBS 0.008242f
C877 B.n837 VSUBS 0.008242f
C878 B.n838 VSUBS 0.008242f
C879 B.n839 VSUBS 0.008242f
C880 B.n840 VSUBS 0.008242f
C881 B.n841 VSUBS 0.008242f
C882 B.n842 VSUBS 0.008242f
C883 B.n843 VSUBS 0.008242f
C884 B.n844 VSUBS 0.008242f
C885 B.n845 VSUBS 0.008242f
C886 B.n846 VSUBS 0.008242f
C887 B.n847 VSUBS 0.008242f
C888 B.n848 VSUBS 0.008242f
C889 B.n849 VSUBS 0.008242f
C890 B.n850 VSUBS 0.008242f
C891 B.n851 VSUBS 0.018662f
C892 VDD2.t3 VSUBS 4.39522f
C893 VDD2.t4 VSUBS 0.40484f
C894 VDD2.t5 VSUBS 0.40484f
C895 VDD2.n0 VSUBS 3.37686f
C896 VDD2.n1 VSUBS 1.45504f
C897 VDD2.t6 VSUBS 0.40484f
C898 VDD2.t1 VSUBS 0.40484f
C899 VDD2.n2 VSUBS 3.38837f
C900 VDD2.n3 VSUBS 3.18009f
C901 VDD2.t9 VSUBS 4.37925f
C902 VDD2.n4 VSUBS 3.74683f
C903 VDD2.t0 VSUBS 0.40484f
C904 VDD2.t8 VSUBS 0.40484f
C905 VDD2.n5 VSUBS 3.37686f
C906 VDD2.n6 VSUBS 0.700904f
C907 VDD2.t2 VSUBS 0.40484f
C908 VDD2.t7 VSUBS 0.40484f
C909 VDD2.n7 VSUBS 3.38831f
C910 VN.n0 VSUBS 0.036654f
C911 VN.t8 VSUBS 2.55953f
C912 VN.n1 VSUBS 0.061676f
C913 VN.n2 VSUBS 0.036654f
C914 VN.t4 VSUBS 2.55953f
C915 VN.n3 VSUBS 0.936557f
C916 VN.n4 VSUBS 0.036654f
C917 VN.t5 VSUBS 2.55953f
C918 VN.n5 VSUBS 0.955332f
C919 VN.t6 VSUBS 2.64252f
C920 VN.n6 VSUBS 0.991303f
C921 VN.n7 VSUBS 0.195219f
C922 VN.n8 VSUBS 0.044705f
C923 VN.n9 VSUBS 0.045851f
C924 VN.n10 VSUBS 0.061172f
C925 VN.n11 VSUBS 0.036654f
C926 VN.n12 VSUBS 0.036654f
C927 VN.n13 VSUBS 0.036654f
C928 VN.n14 VSUBS 0.061172f
C929 VN.n15 VSUBS 0.045851f
C930 VN.t3 VSUBS 2.55953f
C931 VN.n16 VSUBS 0.901971f
C932 VN.n17 VSUBS 0.044705f
C933 VN.n18 VSUBS 0.036654f
C934 VN.n19 VSUBS 0.036654f
C935 VN.n20 VSUBS 0.036654f
C936 VN.n21 VSUBS 0.029928f
C937 VN.n22 VSUBS 0.060124f
C938 VN.n23 VSUBS 0.974008f
C939 VN.n24 VSUBS 0.032776f
C940 VN.n25 VSUBS 0.036654f
C941 VN.t0 VSUBS 2.55953f
C942 VN.n26 VSUBS 0.061676f
C943 VN.n27 VSUBS 0.036654f
C944 VN.t9 VSUBS 2.55953f
C945 VN.n28 VSUBS 0.901971f
C946 VN.t1 VSUBS 2.55953f
C947 VN.n29 VSUBS 0.936557f
C948 VN.n30 VSUBS 0.036654f
C949 VN.t7 VSUBS 2.55953f
C950 VN.n31 VSUBS 0.955332f
C951 VN.t2 VSUBS 2.64252f
C952 VN.n32 VSUBS 0.991303f
C953 VN.n33 VSUBS 0.195219f
C954 VN.n34 VSUBS 0.044705f
C955 VN.n35 VSUBS 0.045851f
C956 VN.n36 VSUBS 0.061172f
C957 VN.n37 VSUBS 0.036654f
C958 VN.n38 VSUBS 0.036654f
C959 VN.n39 VSUBS 0.036654f
C960 VN.n40 VSUBS 0.061172f
C961 VN.n41 VSUBS 0.045851f
C962 VN.n42 VSUBS 0.044705f
C963 VN.n43 VSUBS 0.036654f
C964 VN.n44 VSUBS 0.036654f
C965 VN.n45 VSUBS 0.036654f
C966 VN.n46 VSUBS 0.029928f
C967 VN.n47 VSUBS 0.060124f
C968 VN.n48 VSUBS 0.974008f
C969 VN.n49 VSUBS 2.11514f
C970 VTAIL.t2 VSUBS 0.408217f
C971 VTAIL.t3 VSUBS 0.408217f
C972 VTAIL.n0 VSUBS 3.22197f
C973 VTAIL.n1 VSUBS 0.893965f
C974 VTAIL.t15 VSUBS 4.20531f
C975 VTAIL.n2 VSUBS 1.04972f
C976 VTAIL.t9 VSUBS 0.408217f
C977 VTAIL.t14 VSUBS 0.408217f
C978 VTAIL.n3 VSUBS 3.22197f
C979 VTAIL.n4 VSUBS 0.940651f
C980 VTAIL.t10 VSUBS 0.408217f
C981 VTAIL.t11 VSUBS 0.408217f
C982 VTAIL.n5 VSUBS 3.22197f
C983 VTAIL.n6 VSUBS 2.86413f
C984 VTAIL.t4 VSUBS 0.408217f
C985 VTAIL.t5 VSUBS 0.408217f
C986 VTAIL.n7 VSUBS 3.22197f
C987 VTAIL.n8 VSUBS 2.86413f
C988 VTAIL.t19 VSUBS 0.408217f
C989 VTAIL.t6 VSUBS 0.408217f
C990 VTAIL.n9 VSUBS 3.22197f
C991 VTAIL.n10 VSUBS 0.940651f
C992 VTAIL.t0 VSUBS 4.20531f
C993 VTAIL.n11 VSUBS 1.04971f
C994 VTAIL.t17 VSUBS 0.408217f
C995 VTAIL.t16 VSUBS 0.408217f
C996 VTAIL.n12 VSUBS 3.22197f
C997 VTAIL.n13 VSUBS 0.919736f
C998 VTAIL.t12 VSUBS 0.408217f
C999 VTAIL.t18 VSUBS 0.408217f
C1000 VTAIL.n14 VSUBS 3.22197f
C1001 VTAIL.n15 VSUBS 0.940651f
C1002 VTAIL.t13 VSUBS 4.20531f
C1003 VTAIL.n16 VSUBS 2.87087f
C1004 VTAIL.t1 VSUBS 4.20531f
C1005 VTAIL.n17 VSUBS 2.87087f
C1006 VTAIL.t8 VSUBS 0.408217f
C1007 VTAIL.t7 VSUBS 0.408217f
C1008 VTAIL.n18 VSUBS 3.22197f
C1009 VTAIL.n19 VSUBS 0.84317f
C1010 VDD1.t6 VSUBS 4.39541f
C1011 VDD1.t5 VSUBS 0.404857f
C1012 VDD1.t8 VSUBS 0.404857f
C1013 VDD1.n0 VSUBS 3.377f
C1014 VDD1.n1 VSUBS 1.46279f
C1015 VDD1.t3 VSUBS 4.39541f
C1016 VDD1.t4 VSUBS 0.404857f
C1017 VDD1.t7 VSUBS 0.404857f
C1018 VDD1.n2 VSUBS 3.377f
C1019 VDD1.n3 VSUBS 1.4551f
C1020 VDD1.t0 VSUBS 0.404857f
C1021 VDD1.t1 VSUBS 0.404857f
C1022 VDD1.n4 VSUBS 3.38851f
C1023 VDD1.n5 VSUBS 3.28126f
C1024 VDD1.t2 VSUBS 0.404857f
C1025 VDD1.t9 VSUBS 0.404857f
C1026 VDD1.n6 VSUBS 3.37699f
C1027 VDD1.n7 VSUBS 3.72942f
C1028 VP.n0 VSUBS 0.037319f
C1029 VP.t3 VSUBS 2.60594f
C1030 VP.n1 VSUBS 0.062794f
C1031 VP.n2 VSUBS 0.037319f
C1032 VP.t9 VSUBS 2.60594f
C1033 VP.n3 VSUBS 0.953539f
C1034 VP.n4 VSUBS 0.037319f
C1035 VP.t7 VSUBS 2.60594f
C1036 VP.n5 VSUBS 0.918325f
C1037 VP.n6 VSUBS 0.037319f
C1038 VP.t8 VSUBS 2.60594f
C1039 VP.n7 VSUBS 0.991669f
C1040 VP.n8 VSUBS 0.037319f
C1041 VP.t5 VSUBS 2.60594f
C1042 VP.n9 VSUBS 0.062794f
C1043 VP.n10 VSUBS 0.037319f
C1044 VP.t6 VSUBS 2.60594f
C1045 VP.n11 VSUBS 0.953539f
C1046 VP.n12 VSUBS 0.037319f
C1047 VP.t2 VSUBS 2.60594f
C1048 VP.n13 VSUBS 0.972654f
C1049 VP.t1 VSUBS 2.69043f
C1050 VP.n14 VSUBS 1.00928f
C1051 VP.n15 VSUBS 0.198759f
C1052 VP.n16 VSUBS 0.045516f
C1053 VP.n17 VSUBS 0.046683f
C1054 VP.n18 VSUBS 0.062281f
C1055 VP.n19 VSUBS 0.037319f
C1056 VP.n20 VSUBS 0.037319f
C1057 VP.n21 VSUBS 0.037319f
C1058 VP.n22 VSUBS 0.062281f
C1059 VP.n23 VSUBS 0.046683f
C1060 VP.t0 VSUBS 2.60594f
C1061 VP.n24 VSUBS 0.918325f
C1062 VP.n25 VSUBS 0.045516f
C1063 VP.n26 VSUBS 0.037319f
C1064 VP.n27 VSUBS 0.037319f
C1065 VP.n28 VSUBS 0.037319f
C1066 VP.n29 VSUBS 0.030471f
C1067 VP.n30 VSUBS 0.061214f
C1068 VP.n31 VSUBS 0.991669f
C1069 VP.n32 VSUBS 2.12926f
C1070 VP.n33 VSUBS 2.15528f
C1071 VP.n34 VSUBS 0.037319f
C1072 VP.n35 VSUBS 0.061214f
C1073 VP.n36 VSUBS 0.030471f
C1074 VP.n37 VSUBS 0.062794f
C1075 VP.n38 VSUBS 0.037319f
C1076 VP.n39 VSUBS 0.037319f
C1077 VP.n40 VSUBS 0.045516f
C1078 VP.n41 VSUBS 0.046683f
C1079 VP.n42 VSUBS 0.062281f
C1080 VP.n43 VSUBS 0.037319f
C1081 VP.n44 VSUBS 0.037319f
C1082 VP.n45 VSUBS 0.037319f
C1083 VP.n46 VSUBS 0.062281f
C1084 VP.n47 VSUBS 0.046683f
C1085 VP.t4 VSUBS 2.60594f
C1086 VP.n48 VSUBS 0.918325f
C1087 VP.n49 VSUBS 0.045516f
C1088 VP.n50 VSUBS 0.037319f
C1089 VP.n51 VSUBS 0.037319f
C1090 VP.n52 VSUBS 0.037319f
C1091 VP.n53 VSUBS 0.030471f
C1092 VP.n54 VSUBS 0.061214f
C1093 VP.n55 VSUBS 0.991669f
C1094 VP.n56 VSUBS 0.03337f
.ends

