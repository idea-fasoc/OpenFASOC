* NGSPICE file created from diff_pair_sample_0216.ext - technology: sky130A

.subckt diff_pair_sample_0216 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t5 VN.t0 VTAIL.t5 w_n3538_n1970# sky130_fd_pr__pfet_01v8 ad=0.82665 pd=5.34 as=1.9539 ps=10.8 w=5.01 l=2.88
X1 VTAIL.t8 VN.t1 VDD2.t4 w_n3538_n1970# sky130_fd_pr__pfet_01v8 ad=0.82665 pd=5.34 as=0.82665 ps=5.34 w=5.01 l=2.88
X2 B.t11 B.t9 B.t10 w_n3538_n1970# sky130_fd_pr__pfet_01v8 ad=1.9539 pd=10.8 as=0 ps=0 w=5.01 l=2.88
X3 VDD2.t3 VN.t2 VTAIL.t3 w_n3538_n1970# sky130_fd_pr__pfet_01v8 ad=1.9539 pd=10.8 as=0.82665 ps=5.34 w=5.01 l=2.88
X4 VDD1.t5 VP.t0 VTAIL.t9 w_n3538_n1970# sky130_fd_pr__pfet_01v8 ad=0.82665 pd=5.34 as=1.9539 ps=10.8 w=5.01 l=2.88
X5 VDD1.t4 VP.t1 VTAIL.t11 w_n3538_n1970# sky130_fd_pr__pfet_01v8 ad=1.9539 pd=10.8 as=0.82665 ps=5.34 w=5.01 l=2.88
X6 B.t8 B.t6 B.t7 w_n3538_n1970# sky130_fd_pr__pfet_01v8 ad=1.9539 pd=10.8 as=0 ps=0 w=5.01 l=2.88
X7 VDD2.t2 VN.t3 VTAIL.t4 w_n3538_n1970# sky130_fd_pr__pfet_01v8 ad=0.82665 pd=5.34 as=1.9539 ps=10.8 w=5.01 l=2.88
X8 VTAIL.t10 VP.t2 VDD1.t3 w_n3538_n1970# sky130_fd_pr__pfet_01v8 ad=0.82665 pd=5.34 as=0.82665 ps=5.34 w=5.01 l=2.88
X9 VDD1.t2 VP.t3 VTAIL.t2 w_n3538_n1970# sky130_fd_pr__pfet_01v8 ad=1.9539 pd=10.8 as=0.82665 ps=5.34 w=5.01 l=2.88
X10 VDD1.t1 VP.t4 VTAIL.t1 w_n3538_n1970# sky130_fd_pr__pfet_01v8 ad=0.82665 pd=5.34 as=1.9539 ps=10.8 w=5.01 l=2.88
X11 B.t5 B.t3 B.t4 w_n3538_n1970# sky130_fd_pr__pfet_01v8 ad=1.9539 pd=10.8 as=0 ps=0 w=5.01 l=2.88
X12 VTAIL.t0 VP.t5 VDD1.t0 w_n3538_n1970# sky130_fd_pr__pfet_01v8 ad=0.82665 pd=5.34 as=0.82665 ps=5.34 w=5.01 l=2.88
X13 B.t2 B.t0 B.t1 w_n3538_n1970# sky130_fd_pr__pfet_01v8 ad=1.9539 pd=10.8 as=0 ps=0 w=5.01 l=2.88
X14 VDD2.t1 VN.t4 VTAIL.t7 w_n3538_n1970# sky130_fd_pr__pfet_01v8 ad=1.9539 pd=10.8 as=0.82665 ps=5.34 w=5.01 l=2.88
X15 VTAIL.t6 VN.t5 VDD2.t0 w_n3538_n1970# sky130_fd_pr__pfet_01v8 ad=0.82665 pd=5.34 as=0.82665 ps=5.34 w=5.01 l=2.88
R0 VN.n30 VN.n29 161.3
R1 VN.n28 VN.n17 161.3
R2 VN.n27 VN.n26 161.3
R3 VN.n25 VN.n18 161.3
R4 VN.n24 VN.n23 161.3
R5 VN.n22 VN.n19 161.3
R6 VN.n14 VN.n13 161.3
R7 VN.n12 VN.n1 161.3
R8 VN.n11 VN.n10 161.3
R9 VN.n9 VN.n2 161.3
R10 VN.n8 VN.n7 161.3
R11 VN.n6 VN.n3 161.3
R12 VN.n20 VN.t3 73.7447
R13 VN.n4 VN.t2 73.7447
R14 VN.n15 VN.n0 67.5578
R15 VN.n31 VN.n16 67.5578
R16 VN.n5 VN.n4 61.5425
R17 VN.n21 VN.n20 61.5425
R18 VN.n11 VN.n2 54.5767
R19 VN.n27 VN.n18 54.5767
R20 VN VN.n31 44.7745
R21 VN.n5 VN.t1 41.9245
R22 VN.n0 VN.t0 41.9245
R23 VN.n21 VN.t5 41.9245
R24 VN.n16 VN.t4 41.9245
R25 VN.n12 VN.n11 26.41
R26 VN.n28 VN.n27 26.41
R27 VN.n7 VN.n6 24.4675
R28 VN.n7 VN.n2 24.4675
R29 VN.n13 VN.n12 24.4675
R30 VN.n23 VN.n18 24.4675
R31 VN.n23 VN.n22 24.4675
R32 VN.n29 VN.n28 24.4675
R33 VN.n13 VN.n0 22.5101
R34 VN.n29 VN.n16 22.5101
R35 VN.n6 VN.n5 12.234
R36 VN.n22 VN.n21 12.234
R37 VN.n20 VN.n19 5.36474
R38 VN.n4 VN.n3 5.36474
R39 VN.n31 VN.n30 0.354971
R40 VN.n15 VN.n14 0.354971
R41 VN VN.n15 0.26696
R42 VN.n30 VN.n17 0.189894
R43 VN.n26 VN.n17 0.189894
R44 VN.n26 VN.n25 0.189894
R45 VN.n25 VN.n24 0.189894
R46 VN.n24 VN.n19 0.189894
R47 VN.n8 VN.n3 0.189894
R48 VN.n9 VN.n8 0.189894
R49 VN.n10 VN.n9 0.189894
R50 VN.n10 VN.n1 0.189894
R51 VN.n14 VN.n1 0.189894
R52 VTAIL.n7 VTAIL.t4 91.9954
R53 VTAIL.n11 VTAIL.t5 91.9953
R54 VTAIL.n2 VTAIL.t1 91.9953
R55 VTAIL.n10 VTAIL.t9 91.9953
R56 VTAIL.n9 VTAIL.n8 85.5075
R57 VTAIL.n6 VTAIL.n5 85.5075
R58 VTAIL.n1 VTAIL.n0 85.5072
R59 VTAIL.n4 VTAIL.n3 85.5072
R60 VTAIL.n6 VTAIL.n4 22.2203
R61 VTAIL.n11 VTAIL.n10 19.4531
R62 VTAIL.n0 VTAIL.t3 6.48852
R63 VTAIL.n0 VTAIL.t8 6.48852
R64 VTAIL.n3 VTAIL.t2 6.48852
R65 VTAIL.n3 VTAIL.t10 6.48852
R66 VTAIL.n8 VTAIL.t11 6.48852
R67 VTAIL.n8 VTAIL.t0 6.48852
R68 VTAIL.n5 VTAIL.t7 6.48852
R69 VTAIL.n5 VTAIL.t6 6.48852
R70 VTAIL.n7 VTAIL.n6 2.76774
R71 VTAIL.n10 VTAIL.n9 2.76774
R72 VTAIL.n4 VTAIL.n2 2.76774
R73 VTAIL VTAIL.n11 2.01774
R74 VTAIL.n9 VTAIL.n7 1.85395
R75 VTAIL.n2 VTAIL.n1 1.85395
R76 VTAIL VTAIL.n1 0.7505
R77 VDD2.n1 VDD2.t3 110.695
R78 VDD2.n2 VDD2.t1 108.674
R79 VDD2.n1 VDD2.n0 102.823
R80 VDD2 VDD2.n3 102.82
R81 VDD2.n2 VDD2.n1 37.0278
R82 VDD2.n3 VDD2.t0 6.48852
R83 VDD2.n3 VDD2.t2 6.48852
R84 VDD2.n0 VDD2.t4 6.48852
R85 VDD2.n0 VDD2.t5 6.48852
R86 VDD2 VDD2.n2 2.13412
R87 B.n443 B.n442 585
R88 B.n444 B.n55 585
R89 B.n446 B.n445 585
R90 B.n447 B.n54 585
R91 B.n449 B.n448 585
R92 B.n450 B.n53 585
R93 B.n452 B.n451 585
R94 B.n453 B.n52 585
R95 B.n455 B.n454 585
R96 B.n456 B.n51 585
R97 B.n458 B.n457 585
R98 B.n459 B.n50 585
R99 B.n461 B.n460 585
R100 B.n462 B.n49 585
R101 B.n464 B.n463 585
R102 B.n465 B.n48 585
R103 B.n467 B.n466 585
R104 B.n468 B.n47 585
R105 B.n470 B.n469 585
R106 B.n471 B.n43 585
R107 B.n473 B.n472 585
R108 B.n474 B.n42 585
R109 B.n476 B.n475 585
R110 B.n477 B.n41 585
R111 B.n479 B.n478 585
R112 B.n480 B.n40 585
R113 B.n482 B.n481 585
R114 B.n483 B.n39 585
R115 B.n485 B.n484 585
R116 B.n486 B.n38 585
R117 B.n488 B.n487 585
R118 B.n490 B.n35 585
R119 B.n492 B.n491 585
R120 B.n493 B.n34 585
R121 B.n495 B.n494 585
R122 B.n496 B.n33 585
R123 B.n498 B.n497 585
R124 B.n499 B.n32 585
R125 B.n501 B.n500 585
R126 B.n502 B.n31 585
R127 B.n504 B.n503 585
R128 B.n505 B.n30 585
R129 B.n507 B.n506 585
R130 B.n508 B.n29 585
R131 B.n510 B.n509 585
R132 B.n511 B.n28 585
R133 B.n513 B.n512 585
R134 B.n514 B.n27 585
R135 B.n516 B.n515 585
R136 B.n517 B.n26 585
R137 B.n519 B.n518 585
R138 B.n520 B.n25 585
R139 B.n441 B.n56 585
R140 B.n440 B.n439 585
R141 B.n438 B.n57 585
R142 B.n437 B.n436 585
R143 B.n435 B.n58 585
R144 B.n434 B.n433 585
R145 B.n432 B.n59 585
R146 B.n431 B.n430 585
R147 B.n429 B.n60 585
R148 B.n428 B.n427 585
R149 B.n426 B.n61 585
R150 B.n425 B.n424 585
R151 B.n423 B.n62 585
R152 B.n422 B.n421 585
R153 B.n420 B.n63 585
R154 B.n419 B.n418 585
R155 B.n417 B.n64 585
R156 B.n416 B.n415 585
R157 B.n414 B.n65 585
R158 B.n413 B.n412 585
R159 B.n411 B.n66 585
R160 B.n410 B.n409 585
R161 B.n408 B.n67 585
R162 B.n407 B.n406 585
R163 B.n405 B.n68 585
R164 B.n404 B.n403 585
R165 B.n402 B.n69 585
R166 B.n401 B.n400 585
R167 B.n399 B.n70 585
R168 B.n398 B.n397 585
R169 B.n396 B.n71 585
R170 B.n395 B.n394 585
R171 B.n393 B.n72 585
R172 B.n392 B.n391 585
R173 B.n390 B.n73 585
R174 B.n389 B.n388 585
R175 B.n387 B.n74 585
R176 B.n386 B.n385 585
R177 B.n384 B.n75 585
R178 B.n383 B.n382 585
R179 B.n381 B.n76 585
R180 B.n380 B.n379 585
R181 B.n378 B.n77 585
R182 B.n377 B.n376 585
R183 B.n375 B.n78 585
R184 B.n374 B.n373 585
R185 B.n372 B.n79 585
R186 B.n371 B.n370 585
R187 B.n369 B.n80 585
R188 B.n368 B.n367 585
R189 B.n366 B.n81 585
R190 B.n365 B.n364 585
R191 B.n363 B.n82 585
R192 B.n362 B.n361 585
R193 B.n360 B.n83 585
R194 B.n359 B.n358 585
R195 B.n357 B.n84 585
R196 B.n356 B.n355 585
R197 B.n354 B.n85 585
R198 B.n353 B.n352 585
R199 B.n351 B.n86 585
R200 B.n350 B.n349 585
R201 B.n348 B.n87 585
R202 B.n347 B.n346 585
R203 B.n345 B.n88 585
R204 B.n344 B.n343 585
R205 B.n342 B.n89 585
R206 B.n341 B.n340 585
R207 B.n339 B.n90 585
R208 B.n338 B.n337 585
R209 B.n336 B.n91 585
R210 B.n335 B.n334 585
R211 B.n333 B.n92 585
R212 B.n332 B.n331 585
R213 B.n330 B.n93 585
R214 B.n329 B.n328 585
R215 B.n327 B.n94 585
R216 B.n326 B.n325 585
R217 B.n324 B.n95 585
R218 B.n323 B.n322 585
R219 B.n321 B.n96 585
R220 B.n320 B.n319 585
R221 B.n318 B.n97 585
R222 B.n317 B.n316 585
R223 B.n315 B.n98 585
R224 B.n314 B.n313 585
R225 B.n312 B.n99 585
R226 B.n311 B.n310 585
R227 B.n309 B.n100 585
R228 B.n308 B.n307 585
R229 B.n306 B.n101 585
R230 B.n305 B.n304 585
R231 B.n303 B.n102 585
R232 B.n224 B.n223 585
R233 B.n225 B.n132 585
R234 B.n227 B.n226 585
R235 B.n228 B.n131 585
R236 B.n230 B.n229 585
R237 B.n231 B.n130 585
R238 B.n233 B.n232 585
R239 B.n234 B.n129 585
R240 B.n236 B.n235 585
R241 B.n237 B.n128 585
R242 B.n239 B.n238 585
R243 B.n240 B.n127 585
R244 B.n242 B.n241 585
R245 B.n243 B.n126 585
R246 B.n245 B.n244 585
R247 B.n246 B.n125 585
R248 B.n248 B.n247 585
R249 B.n249 B.n124 585
R250 B.n251 B.n250 585
R251 B.n252 B.n123 585
R252 B.n254 B.n253 585
R253 B.n256 B.n120 585
R254 B.n258 B.n257 585
R255 B.n259 B.n119 585
R256 B.n261 B.n260 585
R257 B.n262 B.n118 585
R258 B.n264 B.n263 585
R259 B.n265 B.n117 585
R260 B.n267 B.n266 585
R261 B.n268 B.n116 585
R262 B.n270 B.n269 585
R263 B.n272 B.n271 585
R264 B.n273 B.n112 585
R265 B.n275 B.n274 585
R266 B.n276 B.n111 585
R267 B.n278 B.n277 585
R268 B.n279 B.n110 585
R269 B.n281 B.n280 585
R270 B.n282 B.n109 585
R271 B.n284 B.n283 585
R272 B.n285 B.n108 585
R273 B.n287 B.n286 585
R274 B.n288 B.n107 585
R275 B.n290 B.n289 585
R276 B.n291 B.n106 585
R277 B.n293 B.n292 585
R278 B.n294 B.n105 585
R279 B.n296 B.n295 585
R280 B.n297 B.n104 585
R281 B.n299 B.n298 585
R282 B.n300 B.n103 585
R283 B.n302 B.n301 585
R284 B.n222 B.n133 585
R285 B.n221 B.n220 585
R286 B.n219 B.n134 585
R287 B.n218 B.n217 585
R288 B.n216 B.n135 585
R289 B.n215 B.n214 585
R290 B.n213 B.n136 585
R291 B.n212 B.n211 585
R292 B.n210 B.n137 585
R293 B.n209 B.n208 585
R294 B.n207 B.n138 585
R295 B.n206 B.n205 585
R296 B.n204 B.n139 585
R297 B.n203 B.n202 585
R298 B.n201 B.n140 585
R299 B.n200 B.n199 585
R300 B.n198 B.n141 585
R301 B.n197 B.n196 585
R302 B.n195 B.n142 585
R303 B.n194 B.n193 585
R304 B.n192 B.n143 585
R305 B.n191 B.n190 585
R306 B.n189 B.n144 585
R307 B.n188 B.n187 585
R308 B.n186 B.n145 585
R309 B.n185 B.n184 585
R310 B.n183 B.n146 585
R311 B.n182 B.n181 585
R312 B.n180 B.n147 585
R313 B.n179 B.n178 585
R314 B.n177 B.n148 585
R315 B.n176 B.n175 585
R316 B.n174 B.n149 585
R317 B.n173 B.n172 585
R318 B.n171 B.n150 585
R319 B.n170 B.n169 585
R320 B.n168 B.n151 585
R321 B.n167 B.n166 585
R322 B.n165 B.n152 585
R323 B.n164 B.n163 585
R324 B.n162 B.n153 585
R325 B.n161 B.n160 585
R326 B.n159 B.n154 585
R327 B.n158 B.n157 585
R328 B.n156 B.n155 585
R329 B.n2 B.n0 585
R330 B.n589 B.n1 585
R331 B.n588 B.n587 585
R332 B.n586 B.n3 585
R333 B.n585 B.n584 585
R334 B.n583 B.n4 585
R335 B.n582 B.n581 585
R336 B.n580 B.n5 585
R337 B.n579 B.n578 585
R338 B.n577 B.n6 585
R339 B.n576 B.n575 585
R340 B.n574 B.n7 585
R341 B.n573 B.n572 585
R342 B.n571 B.n8 585
R343 B.n570 B.n569 585
R344 B.n568 B.n9 585
R345 B.n567 B.n566 585
R346 B.n565 B.n10 585
R347 B.n564 B.n563 585
R348 B.n562 B.n11 585
R349 B.n561 B.n560 585
R350 B.n559 B.n12 585
R351 B.n558 B.n557 585
R352 B.n556 B.n13 585
R353 B.n555 B.n554 585
R354 B.n553 B.n14 585
R355 B.n552 B.n551 585
R356 B.n550 B.n15 585
R357 B.n549 B.n548 585
R358 B.n547 B.n16 585
R359 B.n546 B.n545 585
R360 B.n544 B.n17 585
R361 B.n543 B.n542 585
R362 B.n541 B.n18 585
R363 B.n540 B.n539 585
R364 B.n538 B.n19 585
R365 B.n537 B.n536 585
R366 B.n535 B.n20 585
R367 B.n534 B.n533 585
R368 B.n532 B.n21 585
R369 B.n531 B.n530 585
R370 B.n529 B.n22 585
R371 B.n528 B.n527 585
R372 B.n526 B.n23 585
R373 B.n525 B.n524 585
R374 B.n523 B.n24 585
R375 B.n522 B.n521 585
R376 B.n591 B.n590 585
R377 B.n223 B.n222 454.062
R378 B.n522 B.n25 454.062
R379 B.n301 B.n102 454.062
R380 B.n443 B.n56 454.062
R381 B.n113 B.t9 250.357
R382 B.n121 B.t3 250.357
R383 B.n36 B.t6 250.357
R384 B.n44 B.t0 250.357
R385 B.n113 B.t11 181.609
R386 B.n44 B.t1 181.609
R387 B.n121 B.t5 181.606
R388 B.n36 B.t7 181.606
R389 B.n222 B.n221 163.367
R390 B.n221 B.n134 163.367
R391 B.n217 B.n134 163.367
R392 B.n217 B.n216 163.367
R393 B.n216 B.n215 163.367
R394 B.n215 B.n136 163.367
R395 B.n211 B.n136 163.367
R396 B.n211 B.n210 163.367
R397 B.n210 B.n209 163.367
R398 B.n209 B.n138 163.367
R399 B.n205 B.n138 163.367
R400 B.n205 B.n204 163.367
R401 B.n204 B.n203 163.367
R402 B.n203 B.n140 163.367
R403 B.n199 B.n140 163.367
R404 B.n199 B.n198 163.367
R405 B.n198 B.n197 163.367
R406 B.n197 B.n142 163.367
R407 B.n193 B.n142 163.367
R408 B.n193 B.n192 163.367
R409 B.n192 B.n191 163.367
R410 B.n191 B.n144 163.367
R411 B.n187 B.n144 163.367
R412 B.n187 B.n186 163.367
R413 B.n186 B.n185 163.367
R414 B.n185 B.n146 163.367
R415 B.n181 B.n146 163.367
R416 B.n181 B.n180 163.367
R417 B.n180 B.n179 163.367
R418 B.n179 B.n148 163.367
R419 B.n175 B.n148 163.367
R420 B.n175 B.n174 163.367
R421 B.n174 B.n173 163.367
R422 B.n173 B.n150 163.367
R423 B.n169 B.n150 163.367
R424 B.n169 B.n168 163.367
R425 B.n168 B.n167 163.367
R426 B.n167 B.n152 163.367
R427 B.n163 B.n152 163.367
R428 B.n163 B.n162 163.367
R429 B.n162 B.n161 163.367
R430 B.n161 B.n154 163.367
R431 B.n157 B.n154 163.367
R432 B.n157 B.n156 163.367
R433 B.n156 B.n2 163.367
R434 B.n590 B.n2 163.367
R435 B.n590 B.n589 163.367
R436 B.n589 B.n588 163.367
R437 B.n588 B.n3 163.367
R438 B.n584 B.n3 163.367
R439 B.n584 B.n583 163.367
R440 B.n583 B.n582 163.367
R441 B.n582 B.n5 163.367
R442 B.n578 B.n5 163.367
R443 B.n578 B.n577 163.367
R444 B.n577 B.n576 163.367
R445 B.n576 B.n7 163.367
R446 B.n572 B.n7 163.367
R447 B.n572 B.n571 163.367
R448 B.n571 B.n570 163.367
R449 B.n570 B.n9 163.367
R450 B.n566 B.n9 163.367
R451 B.n566 B.n565 163.367
R452 B.n565 B.n564 163.367
R453 B.n564 B.n11 163.367
R454 B.n560 B.n11 163.367
R455 B.n560 B.n559 163.367
R456 B.n559 B.n558 163.367
R457 B.n558 B.n13 163.367
R458 B.n554 B.n13 163.367
R459 B.n554 B.n553 163.367
R460 B.n553 B.n552 163.367
R461 B.n552 B.n15 163.367
R462 B.n548 B.n15 163.367
R463 B.n548 B.n547 163.367
R464 B.n547 B.n546 163.367
R465 B.n546 B.n17 163.367
R466 B.n542 B.n17 163.367
R467 B.n542 B.n541 163.367
R468 B.n541 B.n540 163.367
R469 B.n540 B.n19 163.367
R470 B.n536 B.n19 163.367
R471 B.n536 B.n535 163.367
R472 B.n535 B.n534 163.367
R473 B.n534 B.n21 163.367
R474 B.n530 B.n21 163.367
R475 B.n530 B.n529 163.367
R476 B.n529 B.n528 163.367
R477 B.n528 B.n23 163.367
R478 B.n524 B.n23 163.367
R479 B.n524 B.n523 163.367
R480 B.n523 B.n522 163.367
R481 B.n223 B.n132 163.367
R482 B.n227 B.n132 163.367
R483 B.n228 B.n227 163.367
R484 B.n229 B.n228 163.367
R485 B.n229 B.n130 163.367
R486 B.n233 B.n130 163.367
R487 B.n234 B.n233 163.367
R488 B.n235 B.n234 163.367
R489 B.n235 B.n128 163.367
R490 B.n239 B.n128 163.367
R491 B.n240 B.n239 163.367
R492 B.n241 B.n240 163.367
R493 B.n241 B.n126 163.367
R494 B.n245 B.n126 163.367
R495 B.n246 B.n245 163.367
R496 B.n247 B.n246 163.367
R497 B.n247 B.n124 163.367
R498 B.n251 B.n124 163.367
R499 B.n252 B.n251 163.367
R500 B.n253 B.n252 163.367
R501 B.n253 B.n120 163.367
R502 B.n258 B.n120 163.367
R503 B.n259 B.n258 163.367
R504 B.n260 B.n259 163.367
R505 B.n260 B.n118 163.367
R506 B.n264 B.n118 163.367
R507 B.n265 B.n264 163.367
R508 B.n266 B.n265 163.367
R509 B.n266 B.n116 163.367
R510 B.n270 B.n116 163.367
R511 B.n271 B.n270 163.367
R512 B.n271 B.n112 163.367
R513 B.n275 B.n112 163.367
R514 B.n276 B.n275 163.367
R515 B.n277 B.n276 163.367
R516 B.n277 B.n110 163.367
R517 B.n281 B.n110 163.367
R518 B.n282 B.n281 163.367
R519 B.n283 B.n282 163.367
R520 B.n283 B.n108 163.367
R521 B.n287 B.n108 163.367
R522 B.n288 B.n287 163.367
R523 B.n289 B.n288 163.367
R524 B.n289 B.n106 163.367
R525 B.n293 B.n106 163.367
R526 B.n294 B.n293 163.367
R527 B.n295 B.n294 163.367
R528 B.n295 B.n104 163.367
R529 B.n299 B.n104 163.367
R530 B.n300 B.n299 163.367
R531 B.n301 B.n300 163.367
R532 B.n305 B.n102 163.367
R533 B.n306 B.n305 163.367
R534 B.n307 B.n306 163.367
R535 B.n307 B.n100 163.367
R536 B.n311 B.n100 163.367
R537 B.n312 B.n311 163.367
R538 B.n313 B.n312 163.367
R539 B.n313 B.n98 163.367
R540 B.n317 B.n98 163.367
R541 B.n318 B.n317 163.367
R542 B.n319 B.n318 163.367
R543 B.n319 B.n96 163.367
R544 B.n323 B.n96 163.367
R545 B.n324 B.n323 163.367
R546 B.n325 B.n324 163.367
R547 B.n325 B.n94 163.367
R548 B.n329 B.n94 163.367
R549 B.n330 B.n329 163.367
R550 B.n331 B.n330 163.367
R551 B.n331 B.n92 163.367
R552 B.n335 B.n92 163.367
R553 B.n336 B.n335 163.367
R554 B.n337 B.n336 163.367
R555 B.n337 B.n90 163.367
R556 B.n341 B.n90 163.367
R557 B.n342 B.n341 163.367
R558 B.n343 B.n342 163.367
R559 B.n343 B.n88 163.367
R560 B.n347 B.n88 163.367
R561 B.n348 B.n347 163.367
R562 B.n349 B.n348 163.367
R563 B.n349 B.n86 163.367
R564 B.n353 B.n86 163.367
R565 B.n354 B.n353 163.367
R566 B.n355 B.n354 163.367
R567 B.n355 B.n84 163.367
R568 B.n359 B.n84 163.367
R569 B.n360 B.n359 163.367
R570 B.n361 B.n360 163.367
R571 B.n361 B.n82 163.367
R572 B.n365 B.n82 163.367
R573 B.n366 B.n365 163.367
R574 B.n367 B.n366 163.367
R575 B.n367 B.n80 163.367
R576 B.n371 B.n80 163.367
R577 B.n372 B.n371 163.367
R578 B.n373 B.n372 163.367
R579 B.n373 B.n78 163.367
R580 B.n377 B.n78 163.367
R581 B.n378 B.n377 163.367
R582 B.n379 B.n378 163.367
R583 B.n379 B.n76 163.367
R584 B.n383 B.n76 163.367
R585 B.n384 B.n383 163.367
R586 B.n385 B.n384 163.367
R587 B.n385 B.n74 163.367
R588 B.n389 B.n74 163.367
R589 B.n390 B.n389 163.367
R590 B.n391 B.n390 163.367
R591 B.n391 B.n72 163.367
R592 B.n395 B.n72 163.367
R593 B.n396 B.n395 163.367
R594 B.n397 B.n396 163.367
R595 B.n397 B.n70 163.367
R596 B.n401 B.n70 163.367
R597 B.n402 B.n401 163.367
R598 B.n403 B.n402 163.367
R599 B.n403 B.n68 163.367
R600 B.n407 B.n68 163.367
R601 B.n408 B.n407 163.367
R602 B.n409 B.n408 163.367
R603 B.n409 B.n66 163.367
R604 B.n413 B.n66 163.367
R605 B.n414 B.n413 163.367
R606 B.n415 B.n414 163.367
R607 B.n415 B.n64 163.367
R608 B.n419 B.n64 163.367
R609 B.n420 B.n419 163.367
R610 B.n421 B.n420 163.367
R611 B.n421 B.n62 163.367
R612 B.n425 B.n62 163.367
R613 B.n426 B.n425 163.367
R614 B.n427 B.n426 163.367
R615 B.n427 B.n60 163.367
R616 B.n431 B.n60 163.367
R617 B.n432 B.n431 163.367
R618 B.n433 B.n432 163.367
R619 B.n433 B.n58 163.367
R620 B.n437 B.n58 163.367
R621 B.n438 B.n437 163.367
R622 B.n439 B.n438 163.367
R623 B.n439 B.n56 163.367
R624 B.n518 B.n25 163.367
R625 B.n518 B.n517 163.367
R626 B.n517 B.n516 163.367
R627 B.n516 B.n27 163.367
R628 B.n512 B.n27 163.367
R629 B.n512 B.n511 163.367
R630 B.n511 B.n510 163.367
R631 B.n510 B.n29 163.367
R632 B.n506 B.n29 163.367
R633 B.n506 B.n505 163.367
R634 B.n505 B.n504 163.367
R635 B.n504 B.n31 163.367
R636 B.n500 B.n31 163.367
R637 B.n500 B.n499 163.367
R638 B.n499 B.n498 163.367
R639 B.n498 B.n33 163.367
R640 B.n494 B.n33 163.367
R641 B.n494 B.n493 163.367
R642 B.n493 B.n492 163.367
R643 B.n492 B.n35 163.367
R644 B.n487 B.n35 163.367
R645 B.n487 B.n486 163.367
R646 B.n486 B.n485 163.367
R647 B.n485 B.n39 163.367
R648 B.n481 B.n39 163.367
R649 B.n481 B.n480 163.367
R650 B.n480 B.n479 163.367
R651 B.n479 B.n41 163.367
R652 B.n475 B.n41 163.367
R653 B.n475 B.n474 163.367
R654 B.n474 B.n473 163.367
R655 B.n473 B.n43 163.367
R656 B.n469 B.n43 163.367
R657 B.n469 B.n468 163.367
R658 B.n468 B.n467 163.367
R659 B.n467 B.n48 163.367
R660 B.n463 B.n48 163.367
R661 B.n463 B.n462 163.367
R662 B.n462 B.n461 163.367
R663 B.n461 B.n50 163.367
R664 B.n457 B.n50 163.367
R665 B.n457 B.n456 163.367
R666 B.n456 B.n455 163.367
R667 B.n455 B.n52 163.367
R668 B.n451 B.n52 163.367
R669 B.n451 B.n450 163.367
R670 B.n450 B.n449 163.367
R671 B.n449 B.n54 163.367
R672 B.n445 B.n54 163.367
R673 B.n445 B.n444 163.367
R674 B.n444 B.n443 163.367
R675 B.n114 B.t10 119.356
R676 B.n45 B.t2 119.356
R677 B.n122 B.t4 119.35
R678 B.n37 B.t8 119.35
R679 B.n114 B.n113 62.255
R680 B.n122 B.n121 62.255
R681 B.n37 B.n36 62.255
R682 B.n45 B.n44 62.255
R683 B.n115 B.n114 59.5399
R684 B.n255 B.n122 59.5399
R685 B.n489 B.n37 59.5399
R686 B.n46 B.n45 59.5399
R687 B.n521 B.n520 29.5029
R688 B.n442 B.n441 29.5029
R689 B.n303 B.n302 29.5029
R690 B.n224 B.n133 29.5029
R691 B B.n591 18.0485
R692 B.n520 B.n519 10.6151
R693 B.n519 B.n26 10.6151
R694 B.n515 B.n26 10.6151
R695 B.n515 B.n514 10.6151
R696 B.n514 B.n513 10.6151
R697 B.n513 B.n28 10.6151
R698 B.n509 B.n28 10.6151
R699 B.n509 B.n508 10.6151
R700 B.n508 B.n507 10.6151
R701 B.n507 B.n30 10.6151
R702 B.n503 B.n30 10.6151
R703 B.n503 B.n502 10.6151
R704 B.n502 B.n501 10.6151
R705 B.n501 B.n32 10.6151
R706 B.n497 B.n32 10.6151
R707 B.n497 B.n496 10.6151
R708 B.n496 B.n495 10.6151
R709 B.n495 B.n34 10.6151
R710 B.n491 B.n34 10.6151
R711 B.n491 B.n490 10.6151
R712 B.n488 B.n38 10.6151
R713 B.n484 B.n38 10.6151
R714 B.n484 B.n483 10.6151
R715 B.n483 B.n482 10.6151
R716 B.n482 B.n40 10.6151
R717 B.n478 B.n40 10.6151
R718 B.n478 B.n477 10.6151
R719 B.n477 B.n476 10.6151
R720 B.n476 B.n42 10.6151
R721 B.n472 B.n471 10.6151
R722 B.n471 B.n470 10.6151
R723 B.n470 B.n47 10.6151
R724 B.n466 B.n47 10.6151
R725 B.n466 B.n465 10.6151
R726 B.n465 B.n464 10.6151
R727 B.n464 B.n49 10.6151
R728 B.n460 B.n49 10.6151
R729 B.n460 B.n459 10.6151
R730 B.n459 B.n458 10.6151
R731 B.n458 B.n51 10.6151
R732 B.n454 B.n51 10.6151
R733 B.n454 B.n453 10.6151
R734 B.n453 B.n452 10.6151
R735 B.n452 B.n53 10.6151
R736 B.n448 B.n53 10.6151
R737 B.n448 B.n447 10.6151
R738 B.n447 B.n446 10.6151
R739 B.n446 B.n55 10.6151
R740 B.n442 B.n55 10.6151
R741 B.n304 B.n303 10.6151
R742 B.n304 B.n101 10.6151
R743 B.n308 B.n101 10.6151
R744 B.n309 B.n308 10.6151
R745 B.n310 B.n309 10.6151
R746 B.n310 B.n99 10.6151
R747 B.n314 B.n99 10.6151
R748 B.n315 B.n314 10.6151
R749 B.n316 B.n315 10.6151
R750 B.n316 B.n97 10.6151
R751 B.n320 B.n97 10.6151
R752 B.n321 B.n320 10.6151
R753 B.n322 B.n321 10.6151
R754 B.n322 B.n95 10.6151
R755 B.n326 B.n95 10.6151
R756 B.n327 B.n326 10.6151
R757 B.n328 B.n327 10.6151
R758 B.n328 B.n93 10.6151
R759 B.n332 B.n93 10.6151
R760 B.n333 B.n332 10.6151
R761 B.n334 B.n333 10.6151
R762 B.n334 B.n91 10.6151
R763 B.n338 B.n91 10.6151
R764 B.n339 B.n338 10.6151
R765 B.n340 B.n339 10.6151
R766 B.n340 B.n89 10.6151
R767 B.n344 B.n89 10.6151
R768 B.n345 B.n344 10.6151
R769 B.n346 B.n345 10.6151
R770 B.n346 B.n87 10.6151
R771 B.n350 B.n87 10.6151
R772 B.n351 B.n350 10.6151
R773 B.n352 B.n351 10.6151
R774 B.n352 B.n85 10.6151
R775 B.n356 B.n85 10.6151
R776 B.n357 B.n356 10.6151
R777 B.n358 B.n357 10.6151
R778 B.n358 B.n83 10.6151
R779 B.n362 B.n83 10.6151
R780 B.n363 B.n362 10.6151
R781 B.n364 B.n363 10.6151
R782 B.n364 B.n81 10.6151
R783 B.n368 B.n81 10.6151
R784 B.n369 B.n368 10.6151
R785 B.n370 B.n369 10.6151
R786 B.n370 B.n79 10.6151
R787 B.n374 B.n79 10.6151
R788 B.n375 B.n374 10.6151
R789 B.n376 B.n375 10.6151
R790 B.n376 B.n77 10.6151
R791 B.n380 B.n77 10.6151
R792 B.n381 B.n380 10.6151
R793 B.n382 B.n381 10.6151
R794 B.n382 B.n75 10.6151
R795 B.n386 B.n75 10.6151
R796 B.n387 B.n386 10.6151
R797 B.n388 B.n387 10.6151
R798 B.n388 B.n73 10.6151
R799 B.n392 B.n73 10.6151
R800 B.n393 B.n392 10.6151
R801 B.n394 B.n393 10.6151
R802 B.n394 B.n71 10.6151
R803 B.n398 B.n71 10.6151
R804 B.n399 B.n398 10.6151
R805 B.n400 B.n399 10.6151
R806 B.n400 B.n69 10.6151
R807 B.n404 B.n69 10.6151
R808 B.n405 B.n404 10.6151
R809 B.n406 B.n405 10.6151
R810 B.n406 B.n67 10.6151
R811 B.n410 B.n67 10.6151
R812 B.n411 B.n410 10.6151
R813 B.n412 B.n411 10.6151
R814 B.n412 B.n65 10.6151
R815 B.n416 B.n65 10.6151
R816 B.n417 B.n416 10.6151
R817 B.n418 B.n417 10.6151
R818 B.n418 B.n63 10.6151
R819 B.n422 B.n63 10.6151
R820 B.n423 B.n422 10.6151
R821 B.n424 B.n423 10.6151
R822 B.n424 B.n61 10.6151
R823 B.n428 B.n61 10.6151
R824 B.n429 B.n428 10.6151
R825 B.n430 B.n429 10.6151
R826 B.n430 B.n59 10.6151
R827 B.n434 B.n59 10.6151
R828 B.n435 B.n434 10.6151
R829 B.n436 B.n435 10.6151
R830 B.n436 B.n57 10.6151
R831 B.n440 B.n57 10.6151
R832 B.n441 B.n440 10.6151
R833 B.n225 B.n224 10.6151
R834 B.n226 B.n225 10.6151
R835 B.n226 B.n131 10.6151
R836 B.n230 B.n131 10.6151
R837 B.n231 B.n230 10.6151
R838 B.n232 B.n231 10.6151
R839 B.n232 B.n129 10.6151
R840 B.n236 B.n129 10.6151
R841 B.n237 B.n236 10.6151
R842 B.n238 B.n237 10.6151
R843 B.n238 B.n127 10.6151
R844 B.n242 B.n127 10.6151
R845 B.n243 B.n242 10.6151
R846 B.n244 B.n243 10.6151
R847 B.n244 B.n125 10.6151
R848 B.n248 B.n125 10.6151
R849 B.n249 B.n248 10.6151
R850 B.n250 B.n249 10.6151
R851 B.n250 B.n123 10.6151
R852 B.n254 B.n123 10.6151
R853 B.n257 B.n256 10.6151
R854 B.n257 B.n119 10.6151
R855 B.n261 B.n119 10.6151
R856 B.n262 B.n261 10.6151
R857 B.n263 B.n262 10.6151
R858 B.n263 B.n117 10.6151
R859 B.n267 B.n117 10.6151
R860 B.n268 B.n267 10.6151
R861 B.n269 B.n268 10.6151
R862 B.n273 B.n272 10.6151
R863 B.n274 B.n273 10.6151
R864 B.n274 B.n111 10.6151
R865 B.n278 B.n111 10.6151
R866 B.n279 B.n278 10.6151
R867 B.n280 B.n279 10.6151
R868 B.n280 B.n109 10.6151
R869 B.n284 B.n109 10.6151
R870 B.n285 B.n284 10.6151
R871 B.n286 B.n285 10.6151
R872 B.n286 B.n107 10.6151
R873 B.n290 B.n107 10.6151
R874 B.n291 B.n290 10.6151
R875 B.n292 B.n291 10.6151
R876 B.n292 B.n105 10.6151
R877 B.n296 B.n105 10.6151
R878 B.n297 B.n296 10.6151
R879 B.n298 B.n297 10.6151
R880 B.n298 B.n103 10.6151
R881 B.n302 B.n103 10.6151
R882 B.n220 B.n133 10.6151
R883 B.n220 B.n219 10.6151
R884 B.n219 B.n218 10.6151
R885 B.n218 B.n135 10.6151
R886 B.n214 B.n135 10.6151
R887 B.n214 B.n213 10.6151
R888 B.n213 B.n212 10.6151
R889 B.n212 B.n137 10.6151
R890 B.n208 B.n137 10.6151
R891 B.n208 B.n207 10.6151
R892 B.n207 B.n206 10.6151
R893 B.n206 B.n139 10.6151
R894 B.n202 B.n139 10.6151
R895 B.n202 B.n201 10.6151
R896 B.n201 B.n200 10.6151
R897 B.n200 B.n141 10.6151
R898 B.n196 B.n141 10.6151
R899 B.n196 B.n195 10.6151
R900 B.n195 B.n194 10.6151
R901 B.n194 B.n143 10.6151
R902 B.n190 B.n143 10.6151
R903 B.n190 B.n189 10.6151
R904 B.n189 B.n188 10.6151
R905 B.n188 B.n145 10.6151
R906 B.n184 B.n145 10.6151
R907 B.n184 B.n183 10.6151
R908 B.n183 B.n182 10.6151
R909 B.n182 B.n147 10.6151
R910 B.n178 B.n147 10.6151
R911 B.n178 B.n177 10.6151
R912 B.n177 B.n176 10.6151
R913 B.n176 B.n149 10.6151
R914 B.n172 B.n149 10.6151
R915 B.n172 B.n171 10.6151
R916 B.n171 B.n170 10.6151
R917 B.n170 B.n151 10.6151
R918 B.n166 B.n151 10.6151
R919 B.n166 B.n165 10.6151
R920 B.n165 B.n164 10.6151
R921 B.n164 B.n153 10.6151
R922 B.n160 B.n153 10.6151
R923 B.n160 B.n159 10.6151
R924 B.n159 B.n158 10.6151
R925 B.n158 B.n155 10.6151
R926 B.n155 B.n0 10.6151
R927 B.n587 B.n1 10.6151
R928 B.n587 B.n586 10.6151
R929 B.n586 B.n585 10.6151
R930 B.n585 B.n4 10.6151
R931 B.n581 B.n4 10.6151
R932 B.n581 B.n580 10.6151
R933 B.n580 B.n579 10.6151
R934 B.n579 B.n6 10.6151
R935 B.n575 B.n6 10.6151
R936 B.n575 B.n574 10.6151
R937 B.n574 B.n573 10.6151
R938 B.n573 B.n8 10.6151
R939 B.n569 B.n8 10.6151
R940 B.n569 B.n568 10.6151
R941 B.n568 B.n567 10.6151
R942 B.n567 B.n10 10.6151
R943 B.n563 B.n10 10.6151
R944 B.n563 B.n562 10.6151
R945 B.n562 B.n561 10.6151
R946 B.n561 B.n12 10.6151
R947 B.n557 B.n12 10.6151
R948 B.n557 B.n556 10.6151
R949 B.n556 B.n555 10.6151
R950 B.n555 B.n14 10.6151
R951 B.n551 B.n14 10.6151
R952 B.n551 B.n550 10.6151
R953 B.n550 B.n549 10.6151
R954 B.n549 B.n16 10.6151
R955 B.n545 B.n16 10.6151
R956 B.n545 B.n544 10.6151
R957 B.n544 B.n543 10.6151
R958 B.n543 B.n18 10.6151
R959 B.n539 B.n18 10.6151
R960 B.n539 B.n538 10.6151
R961 B.n538 B.n537 10.6151
R962 B.n537 B.n20 10.6151
R963 B.n533 B.n20 10.6151
R964 B.n533 B.n532 10.6151
R965 B.n532 B.n531 10.6151
R966 B.n531 B.n22 10.6151
R967 B.n527 B.n22 10.6151
R968 B.n527 B.n526 10.6151
R969 B.n526 B.n525 10.6151
R970 B.n525 B.n24 10.6151
R971 B.n521 B.n24 10.6151
R972 B.n490 B.n489 9.36635
R973 B.n472 B.n46 9.36635
R974 B.n255 B.n254 9.36635
R975 B.n272 B.n115 9.36635
R976 B.n591 B.n0 2.81026
R977 B.n591 B.n1 2.81026
R978 B.n489 B.n488 1.24928
R979 B.n46 B.n42 1.24928
R980 B.n256 B.n255 1.24928
R981 B.n269 B.n115 1.24928
R982 VP.n13 VP.n10 161.3
R983 VP.n15 VP.n14 161.3
R984 VP.n16 VP.n9 161.3
R985 VP.n18 VP.n17 161.3
R986 VP.n19 VP.n8 161.3
R987 VP.n21 VP.n20 161.3
R988 VP.n43 VP.n42 161.3
R989 VP.n41 VP.n1 161.3
R990 VP.n40 VP.n39 161.3
R991 VP.n38 VP.n2 161.3
R992 VP.n37 VP.n36 161.3
R993 VP.n35 VP.n3 161.3
R994 VP.n33 VP.n32 161.3
R995 VP.n31 VP.n4 161.3
R996 VP.n30 VP.n29 161.3
R997 VP.n28 VP.n5 161.3
R998 VP.n27 VP.n26 161.3
R999 VP.n25 VP.n6 161.3
R1000 VP.n11 VP.t1 73.7445
R1001 VP.n24 VP.n23 67.5578
R1002 VP.n44 VP.n0 67.5578
R1003 VP.n22 VP.n7 67.5578
R1004 VP.n12 VP.n11 61.5426
R1005 VP.n29 VP.n28 54.5767
R1006 VP.n40 VP.n2 54.5767
R1007 VP.n18 VP.n9 54.5767
R1008 VP.n24 VP.n22 44.6092
R1009 VP.n23 VP.t3 41.9245
R1010 VP.n34 VP.t2 41.9245
R1011 VP.n0 VP.t4 41.9245
R1012 VP.n7 VP.t0 41.9245
R1013 VP.n12 VP.t5 41.9245
R1014 VP.n28 VP.n27 26.41
R1015 VP.n41 VP.n40 26.41
R1016 VP.n19 VP.n18 26.41
R1017 VP.n27 VP.n6 24.4675
R1018 VP.n29 VP.n4 24.4675
R1019 VP.n33 VP.n4 24.4675
R1020 VP.n36 VP.n35 24.4675
R1021 VP.n36 VP.n2 24.4675
R1022 VP.n42 VP.n41 24.4675
R1023 VP.n20 VP.n19 24.4675
R1024 VP.n14 VP.n13 24.4675
R1025 VP.n14 VP.n9 24.4675
R1026 VP.n23 VP.n6 22.5101
R1027 VP.n42 VP.n0 22.5101
R1028 VP.n20 VP.n7 22.5101
R1029 VP.n34 VP.n33 12.234
R1030 VP.n35 VP.n34 12.234
R1031 VP.n13 VP.n12 12.234
R1032 VP.n11 VP.n10 5.36471
R1033 VP.n22 VP.n21 0.354971
R1034 VP.n25 VP.n24 0.354971
R1035 VP.n44 VP.n43 0.354971
R1036 VP VP.n44 0.26696
R1037 VP.n15 VP.n10 0.189894
R1038 VP.n16 VP.n15 0.189894
R1039 VP.n17 VP.n16 0.189894
R1040 VP.n17 VP.n8 0.189894
R1041 VP.n21 VP.n8 0.189894
R1042 VP.n26 VP.n25 0.189894
R1043 VP.n26 VP.n5 0.189894
R1044 VP.n30 VP.n5 0.189894
R1045 VP.n31 VP.n30 0.189894
R1046 VP.n32 VP.n31 0.189894
R1047 VP.n32 VP.n3 0.189894
R1048 VP.n37 VP.n3 0.189894
R1049 VP.n38 VP.n37 0.189894
R1050 VP.n39 VP.n38 0.189894
R1051 VP.n39 VP.n1 0.189894
R1052 VP.n43 VP.n1 0.189894
R1053 VDD1 VDD1.t4 110.808
R1054 VDD1.n1 VDD1.t2 110.695
R1055 VDD1.n1 VDD1.n0 102.823
R1056 VDD1.n3 VDD1.n2 102.186
R1057 VDD1.n3 VDD1.n1 38.9944
R1058 VDD1.n2 VDD1.t0 6.48852
R1059 VDD1.n2 VDD1.t5 6.48852
R1060 VDD1.n0 VDD1.t3 6.48852
R1061 VDD1.n0 VDD1.t1 6.48852
R1062 VDD1 VDD1.n3 0.634121
C0 VN VTAIL 3.8016f
C1 w_n3538_n1970# VP 7.10957f
C2 VP B 1.93574f
C3 VDD2 VTAIL 5.40627f
C4 VDD2 VN 3.08788f
C5 VTAIL VDD1 5.35181f
C6 w_n3538_n1970# VTAIL 2.02289f
C7 VTAIL B 2.1877f
C8 VN VDD1 0.151163f
C9 VN w_n3538_n1970# 6.65147f
C10 VN B 1.16939f
C11 VDD2 VDD1 1.51571f
C12 VDD2 w_n3538_n1970# 1.96975f
C13 VDD2 B 1.69161f
C14 VP VTAIL 3.81577f
C15 w_n3538_n1970# VDD1 1.87603f
C16 VDD1 B 1.61069f
C17 VN VP 5.9068f
C18 w_n3538_n1970# B 8.11712f
C19 VDD2 VP 0.48579f
C20 VP VDD1 3.41619f
C21 VDD2 VSUBS 1.455622f
C22 VDD1 VSUBS 1.968177f
C23 VTAIL VSUBS 0.687125f
C24 VN VSUBS 5.86245f
C25 VP VSUBS 2.697573f
C26 B VSUBS 4.079394f
C27 w_n3538_n1970# VSUBS 87.332f
C28 VDD1.t4 VSUBS 0.773655f
C29 VDD1.t2 VSUBS 0.772951f
C30 VDD1.t3 VSUBS 0.089296f
C31 VDD1.t1 VSUBS 0.089296f
C32 VDD1.n0 VSUBS 0.565997f
C33 VDD1.n1 VSUBS 2.76651f
C34 VDD1.t0 VSUBS 0.089296f
C35 VDD1.t5 VSUBS 0.089296f
C36 VDD1.n2 VSUBS 0.56227f
C37 VDD1.n3 VSUBS 2.25922f
C38 VP.t4 VSUBS 1.53016f
C39 VP.n0 VSUBS 0.745239f
C40 VP.n1 VSUBS 0.040539f
C41 VP.n2 VSUBS 0.070615f
C42 VP.n3 VSUBS 0.040539f
C43 VP.t2 VSUBS 1.53016f
C44 VP.n4 VSUBS 0.075553f
C45 VP.n5 VSUBS 0.040539f
C46 VP.n6 VSUBS 0.07257f
C47 VP.t0 VSUBS 1.53016f
C48 VP.n7 VSUBS 0.745239f
C49 VP.n8 VSUBS 0.040539f
C50 VP.n9 VSUBS 0.070615f
C51 VP.n10 VSUBS 0.430946f
C52 VP.t5 VSUBS 1.53016f
C53 VP.t1 VSUBS 1.89804f
C54 VP.n11 VSUBS 0.685271f
C55 VP.n12 VSUBS 0.709877f
C56 VP.n13 VSUBS 0.056903f
C57 VP.n14 VSUBS 0.075553f
C58 VP.n15 VSUBS 0.040539f
C59 VP.n16 VSUBS 0.040539f
C60 VP.n17 VSUBS 0.040539f
C61 VP.n18 VSUBS 0.045226f
C62 VP.n19 VSUBS 0.078078f
C63 VP.n20 VSUBS 0.07257f
C64 VP.n21 VSUBS 0.065428f
C65 VP.n22 VSUBS 1.92745f
C66 VP.t3 VSUBS 1.53016f
C67 VP.n23 VSUBS 0.745239f
C68 VP.n24 VSUBS 1.96011f
C69 VP.n25 VSUBS 0.065428f
C70 VP.n26 VSUBS 0.040539f
C71 VP.n27 VSUBS 0.078078f
C72 VP.n28 VSUBS 0.045226f
C73 VP.n29 VSUBS 0.070615f
C74 VP.n30 VSUBS 0.040539f
C75 VP.n31 VSUBS 0.040539f
C76 VP.n32 VSUBS 0.040539f
C77 VP.n33 VSUBS 0.056903f
C78 VP.n34 VSUBS 0.583709f
C79 VP.n35 VSUBS 0.056903f
C80 VP.n36 VSUBS 0.075553f
C81 VP.n37 VSUBS 0.040539f
C82 VP.n38 VSUBS 0.040539f
C83 VP.n39 VSUBS 0.040539f
C84 VP.n40 VSUBS 0.045226f
C85 VP.n41 VSUBS 0.078078f
C86 VP.n42 VSUBS 0.07257f
C87 VP.n43 VSUBS 0.065428f
C88 VP.n44 VSUBS 0.078105f
C89 B.n0 VSUBS 0.005103f
C90 B.n1 VSUBS 0.005103f
C91 B.n2 VSUBS 0.008071f
C92 B.n3 VSUBS 0.008071f
C93 B.n4 VSUBS 0.008071f
C94 B.n5 VSUBS 0.008071f
C95 B.n6 VSUBS 0.008071f
C96 B.n7 VSUBS 0.008071f
C97 B.n8 VSUBS 0.008071f
C98 B.n9 VSUBS 0.008071f
C99 B.n10 VSUBS 0.008071f
C100 B.n11 VSUBS 0.008071f
C101 B.n12 VSUBS 0.008071f
C102 B.n13 VSUBS 0.008071f
C103 B.n14 VSUBS 0.008071f
C104 B.n15 VSUBS 0.008071f
C105 B.n16 VSUBS 0.008071f
C106 B.n17 VSUBS 0.008071f
C107 B.n18 VSUBS 0.008071f
C108 B.n19 VSUBS 0.008071f
C109 B.n20 VSUBS 0.008071f
C110 B.n21 VSUBS 0.008071f
C111 B.n22 VSUBS 0.008071f
C112 B.n23 VSUBS 0.008071f
C113 B.n24 VSUBS 0.008071f
C114 B.n25 VSUBS 0.018212f
C115 B.n26 VSUBS 0.008071f
C116 B.n27 VSUBS 0.008071f
C117 B.n28 VSUBS 0.008071f
C118 B.n29 VSUBS 0.008071f
C119 B.n30 VSUBS 0.008071f
C120 B.n31 VSUBS 0.008071f
C121 B.n32 VSUBS 0.008071f
C122 B.n33 VSUBS 0.008071f
C123 B.n34 VSUBS 0.008071f
C124 B.n35 VSUBS 0.008071f
C125 B.t8 VSUBS 0.161242f
C126 B.t7 VSUBS 0.185532f
C127 B.t6 VSUBS 0.796575f
C128 B.n36 VSUBS 0.122316f
C129 B.n37 VSUBS 0.082369f
C130 B.n38 VSUBS 0.008071f
C131 B.n39 VSUBS 0.008071f
C132 B.n40 VSUBS 0.008071f
C133 B.n41 VSUBS 0.008071f
C134 B.n42 VSUBS 0.00451f
C135 B.n43 VSUBS 0.008071f
C136 B.t2 VSUBS 0.161242f
C137 B.t1 VSUBS 0.185531f
C138 B.t0 VSUBS 0.796575f
C139 B.n44 VSUBS 0.122316f
C140 B.n45 VSUBS 0.082369f
C141 B.n46 VSUBS 0.018699f
C142 B.n47 VSUBS 0.008071f
C143 B.n48 VSUBS 0.008071f
C144 B.n49 VSUBS 0.008071f
C145 B.n50 VSUBS 0.008071f
C146 B.n51 VSUBS 0.008071f
C147 B.n52 VSUBS 0.008071f
C148 B.n53 VSUBS 0.008071f
C149 B.n54 VSUBS 0.008071f
C150 B.n55 VSUBS 0.008071f
C151 B.n56 VSUBS 0.017156f
C152 B.n57 VSUBS 0.008071f
C153 B.n58 VSUBS 0.008071f
C154 B.n59 VSUBS 0.008071f
C155 B.n60 VSUBS 0.008071f
C156 B.n61 VSUBS 0.008071f
C157 B.n62 VSUBS 0.008071f
C158 B.n63 VSUBS 0.008071f
C159 B.n64 VSUBS 0.008071f
C160 B.n65 VSUBS 0.008071f
C161 B.n66 VSUBS 0.008071f
C162 B.n67 VSUBS 0.008071f
C163 B.n68 VSUBS 0.008071f
C164 B.n69 VSUBS 0.008071f
C165 B.n70 VSUBS 0.008071f
C166 B.n71 VSUBS 0.008071f
C167 B.n72 VSUBS 0.008071f
C168 B.n73 VSUBS 0.008071f
C169 B.n74 VSUBS 0.008071f
C170 B.n75 VSUBS 0.008071f
C171 B.n76 VSUBS 0.008071f
C172 B.n77 VSUBS 0.008071f
C173 B.n78 VSUBS 0.008071f
C174 B.n79 VSUBS 0.008071f
C175 B.n80 VSUBS 0.008071f
C176 B.n81 VSUBS 0.008071f
C177 B.n82 VSUBS 0.008071f
C178 B.n83 VSUBS 0.008071f
C179 B.n84 VSUBS 0.008071f
C180 B.n85 VSUBS 0.008071f
C181 B.n86 VSUBS 0.008071f
C182 B.n87 VSUBS 0.008071f
C183 B.n88 VSUBS 0.008071f
C184 B.n89 VSUBS 0.008071f
C185 B.n90 VSUBS 0.008071f
C186 B.n91 VSUBS 0.008071f
C187 B.n92 VSUBS 0.008071f
C188 B.n93 VSUBS 0.008071f
C189 B.n94 VSUBS 0.008071f
C190 B.n95 VSUBS 0.008071f
C191 B.n96 VSUBS 0.008071f
C192 B.n97 VSUBS 0.008071f
C193 B.n98 VSUBS 0.008071f
C194 B.n99 VSUBS 0.008071f
C195 B.n100 VSUBS 0.008071f
C196 B.n101 VSUBS 0.008071f
C197 B.n102 VSUBS 0.017156f
C198 B.n103 VSUBS 0.008071f
C199 B.n104 VSUBS 0.008071f
C200 B.n105 VSUBS 0.008071f
C201 B.n106 VSUBS 0.008071f
C202 B.n107 VSUBS 0.008071f
C203 B.n108 VSUBS 0.008071f
C204 B.n109 VSUBS 0.008071f
C205 B.n110 VSUBS 0.008071f
C206 B.n111 VSUBS 0.008071f
C207 B.n112 VSUBS 0.008071f
C208 B.t10 VSUBS 0.161242f
C209 B.t11 VSUBS 0.185531f
C210 B.t9 VSUBS 0.796575f
C211 B.n113 VSUBS 0.122316f
C212 B.n114 VSUBS 0.082369f
C213 B.n115 VSUBS 0.018699f
C214 B.n116 VSUBS 0.008071f
C215 B.n117 VSUBS 0.008071f
C216 B.n118 VSUBS 0.008071f
C217 B.n119 VSUBS 0.008071f
C218 B.n120 VSUBS 0.008071f
C219 B.t4 VSUBS 0.161242f
C220 B.t5 VSUBS 0.185532f
C221 B.t3 VSUBS 0.796575f
C222 B.n121 VSUBS 0.122316f
C223 B.n122 VSUBS 0.082369f
C224 B.n123 VSUBS 0.008071f
C225 B.n124 VSUBS 0.008071f
C226 B.n125 VSUBS 0.008071f
C227 B.n126 VSUBS 0.008071f
C228 B.n127 VSUBS 0.008071f
C229 B.n128 VSUBS 0.008071f
C230 B.n129 VSUBS 0.008071f
C231 B.n130 VSUBS 0.008071f
C232 B.n131 VSUBS 0.008071f
C233 B.n132 VSUBS 0.008071f
C234 B.n133 VSUBS 0.017156f
C235 B.n134 VSUBS 0.008071f
C236 B.n135 VSUBS 0.008071f
C237 B.n136 VSUBS 0.008071f
C238 B.n137 VSUBS 0.008071f
C239 B.n138 VSUBS 0.008071f
C240 B.n139 VSUBS 0.008071f
C241 B.n140 VSUBS 0.008071f
C242 B.n141 VSUBS 0.008071f
C243 B.n142 VSUBS 0.008071f
C244 B.n143 VSUBS 0.008071f
C245 B.n144 VSUBS 0.008071f
C246 B.n145 VSUBS 0.008071f
C247 B.n146 VSUBS 0.008071f
C248 B.n147 VSUBS 0.008071f
C249 B.n148 VSUBS 0.008071f
C250 B.n149 VSUBS 0.008071f
C251 B.n150 VSUBS 0.008071f
C252 B.n151 VSUBS 0.008071f
C253 B.n152 VSUBS 0.008071f
C254 B.n153 VSUBS 0.008071f
C255 B.n154 VSUBS 0.008071f
C256 B.n155 VSUBS 0.008071f
C257 B.n156 VSUBS 0.008071f
C258 B.n157 VSUBS 0.008071f
C259 B.n158 VSUBS 0.008071f
C260 B.n159 VSUBS 0.008071f
C261 B.n160 VSUBS 0.008071f
C262 B.n161 VSUBS 0.008071f
C263 B.n162 VSUBS 0.008071f
C264 B.n163 VSUBS 0.008071f
C265 B.n164 VSUBS 0.008071f
C266 B.n165 VSUBS 0.008071f
C267 B.n166 VSUBS 0.008071f
C268 B.n167 VSUBS 0.008071f
C269 B.n168 VSUBS 0.008071f
C270 B.n169 VSUBS 0.008071f
C271 B.n170 VSUBS 0.008071f
C272 B.n171 VSUBS 0.008071f
C273 B.n172 VSUBS 0.008071f
C274 B.n173 VSUBS 0.008071f
C275 B.n174 VSUBS 0.008071f
C276 B.n175 VSUBS 0.008071f
C277 B.n176 VSUBS 0.008071f
C278 B.n177 VSUBS 0.008071f
C279 B.n178 VSUBS 0.008071f
C280 B.n179 VSUBS 0.008071f
C281 B.n180 VSUBS 0.008071f
C282 B.n181 VSUBS 0.008071f
C283 B.n182 VSUBS 0.008071f
C284 B.n183 VSUBS 0.008071f
C285 B.n184 VSUBS 0.008071f
C286 B.n185 VSUBS 0.008071f
C287 B.n186 VSUBS 0.008071f
C288 B.n187 VSUBS 0.008071f
C289 B.n188 VSUBS 0.008071f
C290 B.n189 VSUBS 0.008071f
C291 B.n190 VSUBS 0.008071f
C292 B.n191 VSUBS 0.008071f
C293 B.n192 VSUBS 0.008071f
C294 B.n193 VSUBS 0.008071f
C295 B.n194 VSUBS 0.008071f
C296 B.n195 VSUBS 0.008071f
C297 B.n196 VSUBS 0.008071f
C298 B.n197 VSUBS 0.008071f
C299 B.n198 VSUBS 0.008071f
C300 B.n199 VSUBS 0.008071f
C301 B.n200 VSUBS 0.008071f
C302 B.n201 VSUBS 0.008071f
C303 B.n202 VSUBS 0.008071f
C304 B.n203 VSUBS 0.008071f
C305 B.n204 VSUBS 0.008071f
C306 B.n205 VSUBS 0.008071f
C307 B.n206 VSUBS 0.008071f
C308 B.n207 VSUBS 0.008071f
C309 B.n208 VSUBS 0.008071f
C310 B.n209 VSUBS 0.008071f
C311 B.n210 VSUBS 0.008071f
C312 B.n211 VSUBS 0.008071f
C313 B.n212 VSUBS 0.008071f
C314 B.n213 VSUBS 0.008071f
C315 B.n214 VSUBS 0.008071f
C316 B.n215 VSUBS 0.008071f
C317 B.n216 VSUBS 0.008071f
C318 B.n217 VSUBS 0.008071f
C319 B.n218 VSUBS 0.008071f
C320 B.n219 VSUBS 0.008071f
C321 B.n220 VSUBS 0.008071f
C322 B.n221 VSUBS 0.008071f
C323 B.n222 VSUBS 0.017156f
C324 B.n223 VSUBS 0.018212f
C325 B.n224 VSUBS 0.018212f
C326 B.n225 VSUBS 0.008071f
C327 B.n226 VSUBS 0.008071f
C328 B.n227 VSUBS 0.008071f
C329 B.n228 VSUBS 0.008071f
C330 B.n229 VSUBS 0.008071f
C331 B.n230 VSUBS 0.008071f
C332 B.n231 VSUBS 0.008071f
C333 B.n232 VSUBS 0.008071f
C334 B.n233 VSUBS 0.008071f
C335 B.n234 VSUBS 0.008071f
C336 B.n235 VSUBS 0.008071f
C337 B.n236 VSUBS 0.008071f
C338 B.n237 VSUBS 0.008071f
C339 B.n238 VSUBS 0.008071f
C340 B.n239 VSUBS 0.008071f
C341 B.n240 VSUBS 0.008071f
C342 B.n241 VSUBS 0.008071f
C343 B.n242 VSUBS 0.008071f
C344 B.n243 VSUBS 0.008071f
C345 B.n244 VSUBS 0.008071f
C346 B.n245 VSUBS 0.008071f
C347 B.n246 VSUBS 0.008071f
C348 B.n247 VSUBS 0.008071f
C349 B.n248 VSUBS 0.008071f
C350 B.n249 VSUBS 0.008071f
C351 B.n250 VSUBS 0.008071f
C352 B.n251 VSUBS 0.008071f
C353 B.n252 VSUBS 0.008071f
C354 B.n253 VSUBS 0.008071f
C355 B.n254 VSUBS 0.007596f
C356 B.n255 VSUBS 0.018699f
C357 B.n256 VSUBS 0.00451f
C358 B.n257 VSUBS 0.008071f
C359 B.n258 VSUBS 0.008071f
C360 B.n259 VSUBS 0.008071f
C361 B.n260 VSUBS 0.008071f
C362 B.n261 VSUBS 0.008071f
C363 B.n262 VSUBS 0.008071f
C364 B.n263 VSUBS 0.008071f
C365 B.n264 VSUBS 0.008071f
C366 B.n265 VSUBS 0.008071f
C367 B.n266 VSUBS 0.008071f
C368 B.n267 VSUBS 0.008071f
C369 B.n268 VSUBS 0.008071f
C370 B.n269 VSUBS 0.00451f
C371 B.n270 VSUBS 0.008071f
C372 B.n271 VSUBS 0.008071f
C373 B.n272 VSUBS 0.007596f
C374 B.n273 VSUBS 0.008071f
C375 B.n274 VSUBS 0.008071f
C376 B.n275 VSUBS 0.008071f
C377 B.n276 VSUBS 0.008071f
C378 B.n277 VSUBS 0.008071f
C379 B.n278 VSUBS 0.008071f
C380 B.n279 VSUBS 0.008071f
C381 B.n280 VSUBS 0.008071f
C382 B.n281 VSUBS 0.008071f
C383 B.n282 VSUBS 0.008071f
C384 B.n283 VSUBS 0.008071f
C385 B.n284 VSUBS 0.008071f
C386 B.n285 VSUBS 0.008071f
C387 B.n286 VSUBS 0.008071f
C388 B.n287 VSUBS 0.008071f
C389 B.n288 VSUBS 0.008071f
C390 B.n289 VSUBS 0.008071f
C391 B.n290 VSUBS 0.008071f
C392 B.n291 VSUBS 0.008071f
C393 B.n292 VSUBS 0.008071f
C394 B.n293 VSUBS 0.008071f
C395 B.n294 VSUBS 0.008071f
C396 B.n295 VSUBS 0.008071f
C397 B.n296 VSUBS 0.008071f
C398 B.n297 VSUBS 0.008071f
C399 B.n298 VSUBS 0.008071f
C400 B.n299 VSUBS 0.008071f
C401 B.n300 VSUBS 0.008071f
C402 B.n301 VSUBS 0.018212f
C403 B.n302 VSUBS 0.018212f
C404 B.n303 VSUBS 0.017156f
C405 B.n304 VSUBS 0.008071f
C406 B.n305 VSUBS 0.008071f
C407 B.n306 VSUBS 0.008071f
C408 B.n307 VSUBS 0.008071f
C409 B.n308 VSUBS 0.008071f
C410 B.n309 VSUBS 0.008071f
C411 B.n310 VSUBS 0.008071f
C412 B.n311 VSUBS 0.008071f
C413 B.n312 VSUBS 0.008071f
C414 B.n313 VSUBS 0.008071f
C415 B.n314 VSUBS 0.008071f
C416 B.n315 VSUBS 0.008071f
C417 B.n316 VSUBS 0.008071f
C418 B.n317 VSUBS 0.008071f
C419 B.n318 VSUBS 0.008071f
C420 B.n319 VSUBS 0.008071f
C421 B.n320 VSUBS 0.008071f
C422 B.n321 VSUBS 0.008071f
C423 B.n322 VSUBS 0.008071f
C424 B.n323 VSUBS 0.008071f
C425 B.n324 VSUBS 0.008071f
C426 B.n325 VSUBS 0.008071f
C427 B.n326 VSUBS 0.008071f
C428 B.n327 VSUBS 0.008071f
C429 B.n328 VSUBS 0.008071f
C430 B.n329 VSUBS 0.008071f
C431 B.n330 VSUBS 0.008071f
C432 B.n331 VSUBS 0.008071f
C433 B.n332 VSUBS 0.008071f
C434 B.n333 VSUBS 0.008071f
C435 B.n334 VSUBS 0.008071f
C436 B.n335 VSUBS 0.008071f
C437 B.n336 VSUBS 0.008071f
C438 B.n337 VSUBS 0.008071f
C439 B.n338 VSUBS 0.008071f
C440 B.n339 VSUBS 0.008071f
C441 B.n340 VSUBS 0.008071f
C442 B.n341 VSUBS 0.008071f
C443 B.n342 VSUBS 0.008071f
C444 B.n343 VSUBS 0.008071f
C445 B.n344 VSUBS 0.008071f
C446 B.n345 VSUBS 0.008071f
C447 B.n346 VSUBS 0.008071f
C448 B.n347 VSUBS 0.008071f
C449 B.n348 VSUBS 0.008071f
C450 B.n349 VSUBS 0.008071f
C451 B.n350 VSUBS 0.008071f
C452 B.n351 VSUBS 0.008071f
C453 B.n352 VSUBS 0.008071f
C454 B.n353 VSUBS 0.008071f
C455 B.n354 VSUBS 0.008071f
C456 B.n355 VSUBS 0.008071f
C457 B.n356 VSUBS 0.008071f
C458 B.n357 VSUBS 0.008071f
C459 B.n358 VSUBS 0.008071f
C460 B.n359 VSUBS 0.008071f
C461 B.n360 VSUBS 0.008071f
C462 B.n361 VSUBS 0.008071f
C463 B.n362 VSUBS 0.008071f
C464 B.n363 VSUBS 0.008071f
C465 B.n364 VSUBS 0.008071f
C466 B.n365 VSUBS 0.008071f
C467 B.n366 VSUBS 0.008071f
C468 B.n367 VSUBS 0.008071f
C469 B.n368 VSUBS 0.008071f
C470 B.n369 VSUBS 0.008071f
C471 B.n370 VSUBS 0.008071f
C472 B.n371 VSUBS 0.008071f
C473 B.n372 VSUBS 0.008071f
C474 B.n373 VSUBS 0.008071f
C475 B.n374 VSUBS 0.008071f
C476 B.n375 VSUBS 0.008071f
C477 B.n376 VSUBS 0.008071f
C478 B.n377 VSUBS 0.008071f
C479 B.n378 VSUBS 0.008071f
C480 B.n379 VSUBS 0.008071f
C481 B.n380 VSUBS 0.008071f
C482 B.n381 VSUBS 0.008071f
C483 B.n382 VSUBS 0.008071f
C484 B.n383 VSUBS 0.008071f
C485 B.n384 VSUBS 0.008071f
C486 B.n385 VSUBS 0.008071f
C487 B.n386 VSUBS 0.008071f
C488 B.n387 VSUBS 0.008071f
C489 B.n388 VSUBS 0.008071f
C490 B.n389 VSUBS 0.008071f
C491 B.n390 VSUBS 0.008071f
C492 B.n391 VSUBS 0.008071f
C493 B.n392 VSUBS 0.008071f
C494 B.n393 VSUBS 0.008071f
C495 B.n394 VSUBS 0.008071f
C496 B.n395 VSUBS 0.008071f
C497 B.n396 VSUBS 0.008071f
C498 B.n397 VSUBS 0.008071f
C499 B.n398 VSUBS 0.008071f
C500 B.n399 VSUBS 0.008071f
C501 B.n400 VSUBS 0.008071f
C502 B.n401 VSUBS 0.008071f
C503 B.n402 VSUBS 0.008071f
C504 B.n403 VSUBS 0.008071f
C505 B.n404 VSUBS 0.008071f
C506 B.n405 VSUBS 0.008071f
C507 B.n406 VSUBS 0.008071f
C508 B.n407 VSUBS 0.008071f
C509 B.n408 VSUBS 0.008071f
C510 B.n409 VSUBS 0.008071f
C511 B.n410 VSUBS 0.008071f
C512 B.n411 VSUBS 0.008071f
C513 B.n412 VSUBS 0.008071f
C514 B.n413 VSUBS 0.008071f
C515 B.n414 VSUBS 0.008071f
C516 B.n415 VSUBS 0.008071f
C517 B.n416 VSUBS 0.008071f
C518 B.n417 VSUBS 0.008071f
C519 B.n418 VSUBS 0.008071f
C520 B.n419 VSUBS 0.008071f
C521 B.n420 VSUBS 0.008071f
C522 B.n421 VSUBS 0.008071f
C523 B.n422 VSUBS 0.008071f
C524 B.n423 VSUBS 0.008071f
C525 B.n424 VSUBS 0.008071f
C526 B.n425 VSUBS 0.008071f
C527 B.n426 VSUBS 0.008071f
C528 B.n427 VSUBS 0.008071f
C529 B.n428 VSUBS 0.008071f
C530 B.n429 VSUBS 0.008071f
C531 B.n430 VSUBS 0.008071f
C532 B.n431 VSUBS 0.008071f
C533 B.n432 VSUBS 0.008071f
C534 B.n433 VSUBS 0.008071f
C535 B.n434 VSUBS 0.008071f
C536 B.n435 VSUBS 0.008071f
C537 B.n436 VSUBS 0.008071f
C538 B.n437 VSUBS 0.008071f
C539 B.n438 VSUBS 0.008071f
C540 B.n439 VSUBS 0.008071f
C541 B.n440 VSUBS 0.008071f
C542 B.n441 VSUBS 0.018212f
C543 B.n442 VSUBS 0.017156f
C544 B.n443 VSUBS 0.018212f
C545 B.n444 VSUBS 0.008071f
C546 B.n445 VSUBS 0.008071f
C547 B.n446 VSUBS 0.008071f
C548 B.n447 VSUBS 0.008071f
C549 B.n448 VSUBS 0.008071f
C550 B.n449 VSUBS 0.008071f
C551 B.n450 VSUBS 0.008071f
C552 B.n451 VSUBS 0.008071f
C553 B.n452 VSUBS 0.008071f
C554 B.n453 VSUBS 0.008071f
C555 B.n454 VSUBS 0.008071f
C556 B.n455 VSUBS 0.008071f
C557 B.n456 VSUBS 0.008071f
C558 B.n457 VSUBS 0.008071f
C559 B.n458 VSUBS 0.008071f
C560 B.n459 VSUBS 0.008071f
C561 B.n460 VSUBS 0.008071f
C562 B.n461 VSUBS 0.008071f
C563 B.n462 VSUBS 0.008071f
C564 B.n463 VSUBS 0.008071f
C565 B.n464 VSUBS 0.008071f
C566 B.n465 VSUBS 0.008071f
C567 B.n466 VSUBS 0.008071f
C568 B.n467 VSUBS 0.008071f
C569 B.n468 VSUBS 0.008071f
C570 B.n469 VSUBS 0.008071f
C571 B.n470 VSUBS 0.008071f
C572 B.n471 VSUBS 0.008071f
C573 B.n472 VSUBS 0.007596f
C574 B.n473 VSUBS 0.008071f
C575 B.n474 VSUBS 0.008071f
C576 B.n475 VSUBS 0.008071f
C577 B.n476 VSUBS 0.008071f
C578 B.n477 VSUBS 0.008071f
C579 B.n478 VSUBS 0.008071f
C580 B.n479 VSUBS 0.008071f
C581 B.n480 VSUBS 0.008071f
C582 B.n481 VSUBS 0.008071f
C583 B.n482 VSUBS 0.008071f
C584 B.n483 VSUBS 0.008071f
C585 B.n484 VSUBS 0.008071f
C586 B.n485 VSUBS 0.008071f
C587 B.n486 VSUBS 0.008071f
C588 B.n487 VSUBS 0.008071f
C589 B.n488 VSUBS 0.00451f
C590 B.n489 VSUBS 0.018699f
C591 B.n490 VSUBS 0.007596f
C592 B.n491 VSUBS 0.008071f
C593 B.n492 VSUBS 0.008071f
C594 B.n493 VSUBS 0.008071f
C595 B.n494 VSUBS 0.008071f
C596 B.n495 VSUBS 0.008071f
C597 B.n496 VSUBS 0.008071f
C598 B.n497 VSUBS 0.008071f
C599 B.n498 VSUBS 0.008071f
C600 B.n499 VSUBS 0.008071f
C601 B.n500 VSUBS 0.008071f
C602 B.n501 VSUBS 0.008071f
C603 B.n502 VSUBS 0.008071f
C604 B.n503 VSUBS 0.008071f
C605 B.n504 VSUBS 0.008071f
C606 B.n505 VSUBS 0.008071f
C607 B.n506 VSUBS 0.008071f
C608 B.n507 VSUBS 0.008071f
C609 B.n508 VSUBS 0.008071f
C610 B.n509 VSUBS 0.008071f
C611 B.n510 VSUBS 0.008071f
C612 B.n511 VSUBS 0.008071f
C613 B.n512 VSUBS 0.008071f
C614 B.n513 VSUBS 0.008071f
C615 B.n514 VSUBS 0.008071f
C616 B.n515 VSUBS 0.008071f
C617 B.n516 VSUBS 0.008071f
C618 B.n517 VSUBS 0.008071f
C619 B.n518 VSUBS 0.008071f
C620 B.n519 VSUBS 0.008071f
C621 B.n520 VSUBS 0.018212f
C622 B.n521 VSUBS 0.017156f
C623 B.n522 VSUBS 0.017156f
C624 B.n523 VSUBS 0.008071f
C625 B.n524 VSUBS 0.008071f
C626 B.n525 VSUBS 0.008071f
C627 B.n526 VSUBS 0.008071f
C628 B.n527 VSUBS 0.008071f
C629 B.n528 VSUBS 0.008071f
C630 B.n529 VSUBS 0.008071f
C631 B.n530 VSUBS 0.008071f
C632 B.n531 VSUBS 0.008071f
C633 B.n532 VSUBS 0.008071f
C634 B.n533 VSUBS 0.008071f
C635 B.n534 VSUBS 0.008071f
C636 B.n535 VSUBS 0.008071f
C637 B.n536 VSUBS 0.008071f
C638 B.n537 VSUBS 0.008071f
C639 B.n538 VSUBS 0.008071f
C640 B.n539 VSUBS 0.008071f
C641 B.n540 VSUBS 0.008071f
C642 B.n541 VSUBS 0.008071f
C643 B.n542 VSUBS 0.008071f
C644 B.n543 VSUBS 0.008071f
C645 B.n544 VSUBS 0.008071f
C646 B.n545 VSUBS 0.008071f
C647 B.n546 VSUBS 0.008071f
C648 B.n547 VSUBS 0.008071f
C649 B.n548 VSUBS 0.008071f
C650 B.n549 VSUBS 0.008071f
C651 B.n550 VSUBS 0.008071f
C652 B.n551 VSUBS 0.008071f
C653 B.n552 VSUBS 0.008071f
C654 B.n553 VSUBS 0.008071f
C655 B.n554 VSUBS 0.008071f
C656 B.n555 VSUBS 0.008071f
C657 B.n556 VSUBS 0.008071f
C658 B.n557 VSUBS 0.008071f
C659 B.n558 VSUBS 0.008071f
C660 B.n559 VSUBS 0.008071f
C661 B.n560 VSUBS 0.008071f
C662 B.n561 VSUBS 0.008071f
C663 B.n562 VSUBS 0.008071f
C664 B.n563 VSUBS 0.008071f
C665 B.n564 VSUBS 0.008071f
C666 B.n565 VSUBS 0.008071f
C667 B.n566 VSUBS 0.008071f
C668 B.n567 VSUBS 0.008071f
C669 B.n568 VSUBS 0.008071f
C670 B.n569 VSUBS 0.008071f
C671 B.n570 VSUBS 0.008071f
C672 B.n571 VSUBS 0.008071f
C673 B.n572 VSUBS 0.008071f
C674 B.n573 VSUBS 0.008071f
C675 B.n574 VSUBS 0.008071f
C676 B.n575 VSUBS 0.008071f
C677 B.n576 VSUBS 0.008071f
C678 B.n577 VSUBS 0.008071f
C679 B.n578 VSUBS 0.008071f
C680 B.n579 VSUBS 0.008071f
C681 B.n580 VSUBS 0.008071f
C682 B.n581 VSUBS 0.008071f
C683 B.n582 VSUBS 0.008071f
C684 B.n583 VSUBS 0.008071f
C685 B.n584 VSUBS 0.008071f
C686 B.n585 VSUBS 0.008071f
C687 B.n586 VSUBS 0.008071f
C688 B.n587 VSUBS 0.008071f
C689 B.n588 VSUBS 0.008071f
C690 B.n589 VSUBS 0.008071f
C691 B.n590 VSUBS 0.008071f
C692 B.n591 VSUBS 0.018274f
C693 VDD2.t3 VSUBS 0.753736f
C694 VDD2.t4 VSUBS 0.087077f
C695 VDD2.t5 VSUBS 0.087077f
C696 VDD2.n0 VSUBS 0.551927f
C697 VDD2.n1 VSUBS 2.5883f
C698 VDD2.t1 VSUBS 0.744063f
C699 VDD2.n2 VSUBS 2.18316f
C700 VDD2.t0 VSUBS 0.087077f
C701 VDD2.t2 VSUBS 0.087077f
C702 VDD2.n3 VSUBS 0.551904f
C703 VTAIL.t3 VSUBS 0.138841f
C704 VTAIL.t8 VSUBS 0.138841f
C705 VTAIL.n0 VSUBS 0.770973f
C706 VTAIL.n1 VSUBS 0.885888f
C707 VTAIL.t1 VSUBS 1.07834f
C708 VTAIL.n2 VSUBS 1.18513f
C709 VTAIL.t2 VSUBS 0.138841f
C710 VTAIL.t10 VSUBS 0.138841f
C711 VTAIL.n3 VSUBS 0.770973f
C712 VTAIL.n4 VSUBS 2.49423f
C713 VTAIL.t7 VSUBS 0.138841f
C714 VTAIL.t6 VSUBS 0.138841f
C715 VTAIL.n5 VSUBS 0.770977f
C716 VTAIL.n6 VSUBS 2.49422f
C717 VTAIL.t4 VSUBS 1.07835f
C718 VTAIL.n7 VSUBS 1.18512f
C719 VTAIL.t11 VSUBS 0.138841f
C720 VTAIL.t0 VSUBS 0.138841f
C721 VTAIL.n8 VSUBS 0.770977f
C722 VTAIL.n9 VSUBS 1.11383f
C723 VTAIL.t9 VSUBS 1.07834f
C724 VTAIL.n10 VSUBS 2.25281f
C725 VTAIL.t5 VSUBS 1.07834f
C726 VTAIL.n11 VSUBS 2.16806f
C727 VN.t0 VSUBS 1.47298f
C728 VN.n0 VSUBS 0.717391f
C729 VN.n1 VSUBS 0.039024f
C730 VN.n2 VSUBS 0.067976f
C731 VN.n3 VSUBS 0.414841f
C732 VN.t1 VSUBS 1.47298f
C733 VN.t2 VSUBS 1.82711f
C734 VN.n4 VSUBS 0.659662f
C735 VN.n5 VSUBS 0.683349f
C736 VN.n6 VSUBS 0.054777f
C737 VN.n7 VSUBS 0.07273f
C738 VN.n8 VSUBS 0.039024f
C739 VN.n9 VSUBS 0.039024f
C740 VN.n10 VSUBS 0.039024f
C741 VN.n11 VSUBS 0.043536f
C742 VN.n12 VSUBS 0.07516f
C743 VN.n13 VSUBS 0.069858f
C744 VN.n14 VSUBS 0.062983f
C745 VN.n15 VSUBS 0.075186f
C746 VN.t4 VSUBS 1.47298f
C747 VN.n16 VSUBS 0.717391f
C748 VN.n17 VSUBS 0.039024f
C749 VN.n18 VSUBS 0.067976f
C750 VN.n19 VSUBS 0.414841f
C751 VN.t5 VSUBS 1.47298f
C752 VN.t3 VSUBS 1.82711f
C753 VN.n20 VSUBS 0.659662f
C754 VN.n21 VSUBS 0.683349f
C755 VN.n22 VSUBS 0.054777f
C756 VN.n23 VSUBS 0.07273f
C757 VN.n24 VSUBS 0.039024f
C758 VN.n25 VSUBS 0.039024f
C759 VN.n26 VSUBS 0.039024f
C760 VN.n27 VSUBS 0.043536f
C761 VN.n28 VSUBS 0.07516f
C762 VN.n29 VSUBS 0.069858f
C763 VN.n30 VSUBS 0.062983f
C764 VN.n31 VSUBS 1.87205f
.ends

