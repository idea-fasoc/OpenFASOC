* NGSPICE file created from diff_pair_sample_1198.ext - technology: sky130A

.subckt diff_pair_sample_1198 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t3 VP.t0 VTAIL.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=1.79355 pd=11.2 as=4.2393 ps=22.52 w=10.87 l=3.37
X1 B.t17 B.t15 B.t16 B.t12 sky130_fd_pr__nfet_01v8 ad=4.2393 pd=22.52 as=0 ps=0 w=10.87 l=3.37
X2 B.t14 B.t11 B.t13 B.t12 sky130_fd_pr__nfet_01v8 ad=4.2393 pd=22.52 as=0 ps=0 w=10.87 l=3.37
X3 VTAIL.t4 VN.t0 VDD2.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=4.2393 pd=22.52 as=1.79355 ps=11.2 w=10.87 l=3.37
X4 B.t10 B.t8 B.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=4.2393 pd=22.52 as=0 ps=0 w=10.87 l=3.37
X5 VTAIL.t3 VP.t1 VDD1.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=4.2393 pd=22.52 as=1.79355 ps=11.2 w=10.87 l=3.37
X6 VTAIL.t7 VN.t1 VDD2.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=4.2393 pd=22.52 as=1.79355 ps=11.2 w=10.87 l=3.37
X7 VDD2.t1 VN.t2 VTAIL.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=1.79355 pd=11.2 as=4.2393 ps=22.52 w=10.87 l=3.37
X8 VDD2.t0 VN.t3 VTAIL.t5 B.t3 sky130_fd_pr__nfet_01v8 ad=1.79355 pd=11.2 as=4.2393 ps=22.52 w=10.87 l=3.37
X9 VDD1.t1 VP.t2 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.79355 pd=11.2 as=4.2393 ps=22.52 w=10.87 l=3.37
X10 VTAIL.t0 VP.t3 VDD1.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=4.2393 pd=22.52 as=1.79355 ps=11.2 w=10.87 l=3.37
X11 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=4.2393 pd=22.52 as=0 ps=0 w=10.87 l=3.37
R0 VP.n17 VP.n16 161.3
R1 VP.n15 VP.n1 161.3
R2 VP.n14 VP.n13 161.3
R3 VP.n12 VP.n2 161.3
R4 VP.n11 VP.n10 161.3
R5 VP.n9 VP.n3 161.3
R6 VP.n8 VP.n7 161.3
R7 VP.n5 VP.t3 112.817
R8 VP.n5 VP.t2 111.683
R9 VP.n4 VP.t1 77.7355
R10 VP.n0 VP.t0 77.7355
R11 VP.n6 VP.n4 72.9405
R12 VP.n18 VP.n0 72.9405
R13 VP.n6 VP.n5 50.3307
R14 VP.n10 VP.n2 40.4934
R15 VP.n14 VP.n2 40.4934
R16 VP.n9 VP.n8 24.4675
R17 VP.n10 VP.n9 24.4675
R18 VP.n15 VP.n14 24.4675
R19 VP.n16 VP.n15 24.4675
R20 VP.n8 VP.n4 17.1274
R21 VP.n16 VP.n0 17.1274
R22 VP.n7 VP.n6 0.354971
R23 VP.n18 VP.n17 0.354971
R24 VP VP.n18 0.26696
R25 VP.n7 VP.n3 0.189894
R26 VP.n11 VP.n3 0.189894
R27 VP.n12 VP.n11 0.189894
R28 VP.n13 VP.n12 0.189894
R29 VP.n13 VP.n1 0.189894
R30 VP.n17 VP.n1 0.189894
R31 VTAIL.n458 VTAIL.n406 289.615
R32 VTAIL.n52 VTAIL.n0 289.615
R33 VTAIL.n110 VTAIL.n58 289.615
R34 VTAIL.n168 VTAIL.n116 289.615
R35 VTAIL.n400 VTAIL.n348 289.615
R36 VTAIL.n342 VTAIL.n290 289.615
R37 VTAIL.n284 VTAIL.n232 289.615
R38 VTAIL.n226 VTAIL.n174 289.615
R39 VTAIL.n425 VTAIL.n424 185
R40 VTAIL.n422 VTAIL.n421 185
R41 VTAIL.n431 VTAIL.n430 185
R42 VTAIL.n433 VTAIL.n432 185
R43 VTAIL.n418 VTAIL.n417 185
R44 VTAIL.n439 VTAIL.n438 185
R45 VTAIL.n442 VTAIL.n441 185
R46 VTAIL.n440 VTAIL.n414 185
R47 VTAIL.n447 VTAIL.n413 185
R48 VTAIL.n449 VTAIL.n448 185
R49 VTAIL.n451 VTAIL.n450 185
R50 VTAIL.n410 VTAIL.n409 185
R51 VTAIL.n457 VTAIL.n456 185
R52 VTAIL.n459 VTAIL.n458 185
R53 VTAIL.n19 VTAIL.n18 185
R54 VTAIL.n16 VTAIL.n15 185
R55 VTAIL.n25 VTAIL.n24 185
R56 VTAIL.n27 VTAIL.n26 185
R57 VTAIL.n12 VTAIL.n11 185
R58 VTAIL.n33 VTAIL.n32 185
R59 VTAIL.n36 VTAIL.n35 185
R60 VTAIL.n34 VTAIL.n8 185
R61 VTAIL.n41 VTAIL.n7 185
R62 VTAIL.n43 VTAIL.n42 185
R63 VTAIL.n45 VTAIL.n44 185
R64 VTAIL.n4 VTAIL.n3 185
R65 VTAIL.n51 VTAIL.n50 185
R66 VTAIL.n53 VTAIL.n52 185
R67 VTAIL.n77 VTAIL.n76 185
R68 VTAIL.n74 VTAIL.n73 185
R69 VTAIL.n83 VTAIL.n82 185
R70 VTAIL.n85 VTAIL.n84 185
R71 VTAIL.n70 VTAIL.n69 185
R72 VTAIL.n91 VTAIL.n90 185
R73 VTAIL.n94 VTAIL.n93 185
R74 VTAIL.n92 VTAIL.n66 185
R75 VTAIL.n99 VTAIL.n65 185
R76 VTAIL.n101 VTAIL.n100 185
R77 VTAIL.n103 VTAIL.n102 185
R78 VTAIL.n62 VTAIL.n61 185
R79 VTAIL.n109 VTAIL.n108 185
R80 VTAIL.n111 VTAIL.n110 185
R81 VTAIL.n135 VTAIL.n134 185
R82 VTAIL.n132 VTAIL.n131 185
R83 VTAIL.n141 VTAIL.n140 185
R84 VTAIL.n143 VTAIL.n142 185
R85 VTAIL.n128 VTAIL.n127 185
R86 VTAIL.n149 VTAIL.n148 185
R87 VTAIL.n152 VTAIL.n151 185
R88 VTAIL.n150 VTAIL.n124 185
R89 VTAIL.n157 VTAIL.n123 185
R90 VTAIL.n159 VTAIL.n158 185
R91 VTAIL.n161 VTAIL.n160 185
R92 VTAIL.n120 VTAIL.n119 185
R93 VTAIL.n167 VTAIL.n166 185
R94 VTAIL.n169 VTAIL.n168 185
R95 VTAIL.n401 VTAIL.n400 185
R96 VTAIL.n399 VTAIL.n398 185
R97 VTAIL.n352 VTAIL.n351 185
R98 VTAIL.n393 VTAIL.n392 185
R99 VTAIL.n391 VTAIL.n390 185
R100 VTAIL.n389 VTAIL.n355 185
R101 VTAIL.n359 VTAIL.n356 185
R102 VTAIL.n384 VTAIL.n383 185
R103 VTAIL.n382 VTAIL.n381 185
R104 VTAIL.n361 VTAIL.n360 185
R105 VTAIL.n376 VTAIL.n375 185
R106 VTAIL.n374 VTAIL.n373 185
R107 VTAIL.n365 VTAIL.n364 185
R108 VTAIL.n368 VTAIL.n367 185
R109 VTAIL.n343 VTAIL.n342 185
R110 VTAIL.n341 VTAIL.n340 185
R111 VTAIL.n294 VTAIL.n293 185
R112 VTAIL.n335 VTAIL.n334 185
R113 VTAIL.n333 VTAIL.n332 185
R114 VTAIL.n331 VTAIL.n297 185
R115 VTAIL.n301 VTAIL.n298 185
R116 VTAIL.n326 VTAIL.n325 185
R117 VTAIL.n324 VTAIL.n323 185
R118 VTAIL.n303 VTAIL.n302 185
R119 VTAIL.n318 VTAIL.n317 185
R120 VTAIL.n316 VTAIL.n315 185
R121 VTAIL.n307 VTAIL.n306 185
R122 VTAIL.n310 VTAIL.n309 185
R123 VTAIL.n285 VTAIL.n284 185
R124 VTAIL.n283 VTAIL.n282 185
R125 VTAIL.n236 VTAIL.n235 185
R126 VTAIL.n277 VTAIL.n276 185
R127 VTAIL.n275 VTAIL.n274 185
R128 VTAIL.n273 VTAIL.n239 185
R129 VTAIL.n243 VTAIL.n240 185
R130 VTAIL.n268 VTAIL.n267 185
R131 VTAIL.n266 VTAIL.n265 185
R132 VTAIL.n245 VTAIL.n244 185
R133 VTAIL.n260 VTAIL.n259 185
R134 VTAIL.n258 VTAIL.n257 185
R135 VTAIL.n249 VTAIL.n248 185
R136 VTAIL.n252 VTAIL.n251 185
R137 VTAIL.n227 VTAIL.n226 185
R138 VTAIL.n225 VTAIL.n224 185
R139 VTAIL.n178 VTAIL.n177 185
R140 VTAIL.n219 VTAIL.n218 185
R141 VTAIL.n217 VTAIL.n216 185
R142 VTAIL.n215 VTAIL.n181 185
R143 VTAIL.n185 VTAIL.n182 185
R144 VTAIL.n210 VTAIL.n209 185
R145 VTAIL.n208 VTAIL.n207 185
R146 VTAIL.n187 VTAIL.n186 185
R147 VTAIL.n202 VTAIL.n201 185
R148 VTAIL.n200 VTAIL.n199 185
R149 VTAIL.n191 VTAIL.n190 185
R150 VTAIL.n194 VTAIL.n193 185
R151 VTAIL.t6 VTAIL.n423 149.524
R152 VTAIL.t4 VTAIL.n17 149.524
R153 VTAIL.t2 VTAIL.n75 149.524
R154 VTAIL.t3 VTAIL.n133 149.524
R155 VTAIL.t1 VTAIL.n366 149.524
R156 VTAIL.t0 VTAIL.n308 149.524
R157 VTAIL.t5 VTAIL.n250 149.524
R158 VTAIL.t7 VTAIL.n192 149.524
R159 VTAIL.n424 VTAIL.n421 104.615
R160 VTAIL.n431 VTAIL.n421 104.615
R161 VTAIL.n432 VTAIL.n431 104.615
R162 VTAIL.n432 VTAIL.n417 104.615
R163 VTAIL.n439 VTAIL.n417 104.615
R164 VTAIL.n441 VTAIL.n439 104.615
R165 VTAIL.n441 VTAIL.n440 104.615
R166 VTAIL.n440 VTAIL.n413 104.615
R167 VTAIL.n449 VTAIL.n413 104.615
R168 VTAIL.n450 VTAIL.n449 104.615
R169 VTAIL.n450 VTAIL.n409 104.615
R170 VTAIL.n457 VTAIL.n409 104.615
R171 VTAIL.n458 VTAIL.n457 104.615
R172 VTAIL.n18 VTAIL.n15 104.615
R173 VTAIL.n25 VTAIL.n15 104.615
R174 VTAIL.n26 VTAIL.n25 104.615
R175 VTAIL.n26 VTAIL.n11 104.615
R176 VTAIL.n33 VTAIL.n11 104.615
R177 VTAIL.n35 VTAIL.n33 104.615
R178 VTAIL.n35 VTAIL.n34 104.615
R179 VTAIL.n34 VTAIL.n7 104.615
R180 VTAIL.n43 VTAIL.n7 104.615
R181 VTAIL.n44 VTAIL.n43 104.615
R182 VTAIL.n44 VTAIL.n3 104.615
R183 VTAIL.n51 VTAIL.n3 104.615
R184 VTAIL.n52 VTAIL.n51 104.615
R185 VTAIL.n76 VTAIL.n73 104.615
R186 VTAIL.n83 VTAIL.n73 104.615
R187 VTAIL.n84 VTAIL.n83 104.615
R188 VTAIL.n84 VTAIL.n69 104.615
R189 VTAIL.n91 VTAIL.n69 104.615
R190 VTAIL.n93 VTAIL.n91 104.615
R191 VTAIL.n93 VTAIL.n92 104.615
R192 VTAIL.n92 VTAIL.n65 104.615
R193 VTAIL.n101 VTAIL.n65 104.615
R194 VTAIL.n102 VTAIL.n101 104.615
R195 VTAIL.n102 VTAIL.n61 104.615
R196 VTAIL.n109 VTAIL.n61 104.615
R197 VTAIL.n110 VTAIL.n109 104.615
R198 VTAIL.n134 VTAIL.n131 104.615
R199 VTAIL.n141 VTAIL.n131 104.615
R200 VTAIL.n142 VTAIL.n141 104.615
R201 VTAIL.n142 VTAIL.n127 104.615
R202 VTAIL.n149 VTAIL.n127 104.615
R203 VTAIL.n151 VTAIL.n149 104.615
R204 VTAIL.n151 VTAIL.n150 104.615
R205 VTAIL.n150 VTAIL.n123 104.615
R206 VTAIL.n159 VTAIL.n123 104.615
R207 VTAIL.n160 VTAIL.n159 104.615
R208 VTAIL.n160 VTAIL.n119 104.615
R209 VTAIL.n167 VTAIL.n119 104.615
R210 VTAIL.n168 VTAIL.n167 104.615
R211 VTAIL.n400 VTAIL.n399 104.615
R212 VTAIL.n399 VTAIL.n351 104.615
R213 VTAIL.n392 VTAIL.n351 104.615
R214 VTAIL.n392 VTAIL.n391 104.615
R215 VTAIL.n391 VTAIL.n355 104.615
R216 VTAIL.n359 VTAIL.n355 104.615
R217 VTAIL.n383 VTAIL.n359 104.615
R218 VTAIL.n383 VTAIL.n382 104.615
R219 VTAIL.n382 VTAIL.n360 104.615
R220 VTAIL.n375 VTAIL.n360 104.615
R221 VTAIL.n375 VTAIL.n374 104.615
R222 VTAIL.n374 VTAIL.n364 104.615
R223 VTAIL.n367 VTAIL.n364 104.615
R224 VTAIL.n342 VTAIL.n341 104.615
R225 VTAIL.n341 VTAIL.n293 104.615
R226 VTAIL.n334 VTAIL.n293 104.615
R227 VTAIL.n334 VTAIL.n333 104.615
R228 VTAIL.n333 VTAIL.n297 104.615
R229 VTAIL.n301 VTAIL.n297 104.615
R230 VTAIL.n325 VTAIL.n301 104.615
R231 VTAIL.n325 VTAIL.n324 104.615
R232 VTAIL.n324 VTAIL.n302 104.615
R233 VTAIL.n317 VTAIL.n302 104.615
R234 VTAIL.n317 VTAIL.n316 104.615
R235 VTAIL.n316 VTAIL.n306 104.615
R236 VTAIL.n309 VTAIL.n306 104.615
R237 VTAIL.n284 VTAIL.n283 104.615
R238 VTAIL.n283 VTAIL.n235 104.615
R239 VTAIL.n276 VTAIL.n235 104.615
R240 VTAIL.n276 VTAIL.n275 104.615
R241 VTAIL.n275 VTAIL.n239 104.615
R242 VTAIL.n243 VTAIL.n239 104.615
R243 VTAIL.n267 VTAIL.n243 104.615
R244 VTAIL.n267 VTAIL.n266 104.615
R245 VTAIL.n266 VTAIL.n244 104.615
R246 VTAIL.n259 VTAIL.n244 104.615
R247 VTAIL.n259 VTAIL.n258 104.615
R248 VTAIL.n258 VTAIL.n248 104.615
R249 VTAIL.n251 VTAIL.n248 104.615
R250 VTAIL.n226 VTAIL.n225 104.615
R251 VTAIL.n225 VTAIL.n177 104.615
R252 VTAIL.n218 VTAIL.n177 104.615
R253 VTAIL.n218 VTAIL.n217 104.615
R254 VTAIL.n217 VTAIL.n181 104.615
R255 VTAIL.n185 VTAIL.n181 104.615
R256 VTAIL.n209 VTAIL.n185 104.615
R257 VTAIL.n209 VTAIL.n208 104.615
R258 VTAIL.n208 VTAIL.n186 104.615
R259 VTAIL.n201 VTAIL.n186 104.615
R260 VTAIL.n201 VTAIL.n200 104.615
R261 VTAIL.n200 VTAIL.n190 104.615
R262 VTAIL.n193 VTAIL.n190 104.615
R263 VTAIL.n424 VTAIL.t6 52.3082
R264 VTAIL.n18 VTAIL.t4 52.3082
R265 VTAIL.n76 VTAIL.t2 52.3082
R266 VTAIL.n134 VTAIL.t3 52.3082
R267 VTAIL.n367 VTAIL.t1 52.3082
R268 VTAIL.n309 VTAIL.t0 52.3082
R269 VTAIL.n251 VTAIL.t5 52.3082
R270 VTAIL.n193 VTAIL.t7 52.3082
R271 VTAIL.n463 VTAIL.n462 35.8702
R272 VTAIL.n57 VTAIL.n56 35.8702
R273 VTAIL.n115 VTAIL.n114 35.8702
R274 VTAIL.n173 VTAIL.n172 35.8702
R275 VTAIL.n405 VTAIL.n404 35.8702
R276 VTAIL.n347 VTAIL.n346 35.8702
R277 VTAIL.n289 VTAIL.n288 35.8702
R278 VTAIL.n231 VTAIL.n230 35.8702
R279 VTAIL.n463 VTAIL.n405 24.9272
R280 VTAIL.n231 VTAIL.n173 24.9272
R281 VTAIL.n448 VTAIL.n447 13.1884
R282 VTAIL.n42 VTAIL.n41 13.1884
R283 VTAIL.n100 VTAIL.n99 13.1884
R284 VTAIL.n158 VTAIL.n157 13.1884
R285 VTAIL.n390 VTAIL.n389 13.1884
R286 VTAIL.n332 VTAIL.n331 13.1884
R287 VTAIL.n274 VTAIL.n273 13.1884
R288 VTAIL.n216 VTAIL.n215 13.1884
R289 VTAIL.n446 VTAIL.n414 12.8005
R290 VTAIL.n451 VTAIL.n412 12.8005
R291 VTAIL.n40 VTAIL.n8 12.8005
R292 VTAIL.n45 VTAIL.n6 12.8005
R293 VTAIL.n98 VTAIL.n66 12.8005
R294 VTAIL.n103 VTAIL.n64 12.8005
R295 VTAIL.n156 VTAIL.n124 12.8005
R296 VTAIL.n161 VTAIL.n122 12.8005
R297 VTAIL.n393 VTAIL.n354 12.8005
R298 VTAIL.n388 VTAIL.n356 12.8005
R299 VTAIL.n335 VTAIL.n296 12.8005
R300 VTAIL.n330 VTAIL.n298 12.8005
R301 VTAIL.n277 VTAIL.n238 12.8005
R302 VTAIL.n272 VTAIL.n240 12.8005
R303 VTAIL.n219 VTAIL.n180 12.8005
R304 VTAIL.n214 VTAIL.n182 12.8005
R305 VTAIL.n443 VTAIL.n442 12.0247
R306 VTAIL.n452 VTAIL.n410 12.0247
R307 VTAIL.n37 VTAIL.n36 12.0247
R308 VTAIL.n46 VTAIL.n4 12.0247
R309 VTAIL.n95 VTAIL.n94 12.0247
R310 VTAIL.n104 VTAIL.n62 12.0247
R311 VTAIL.n153 VTAIL.n152 12.0247
R312 VTAIL.n162 VTAIL.n120 12.0247
R313 VTAIL.n394 VTAIL.n352 12.0247
R314 VTAIL.n385 VTAIL.n384 12.0247
R315 VTAIL.n336 VTAIL.n294 12.0247
R316 VTAIL.n327 VTAIL.n326 12.0247
R317 VTAIL.n278 VTAIL.n236 12.0247
R318 VTAIL.n269 VTAIL.n268 12.0247
R319 VTAIL.n220 VTAIL.n178 12.0247
R320 VTAIL.n211 VTAIL.n210 12.0247
R321 VTAIL.n438 VTAIL.n416 11.249
R322 VTAIL.n456 VTAIL.n455 11.249
R323 VTAIL.n32 VTAIL.n10 11.249
R324 VTAIL.n50 VTAIL.n49 11.249
R325 VTAIL.n90 VTAIL.n68 11.249
R326 VTAIL.n108 VTAIL.n107 11.249
R327 VTAIL.n148 VTAIL.n126 11.249
R328 VTAIL.n166 VTAIL.n165 11.249
R329 VTAIL.n398 VTAIL.n397 11.249
R330 VTAIL.n381 VTAIL.n358 11.249
R331 VTAIL.n340 VTAIL.n339 11.249
R332 VTAIL.n323 VTAIL.n300 11.249
R333 VTAIL.n282 VTAIL.n281 11.249
R334 VTAIL.n265 VTAIL.n242 11.249
R335 VTAIL.n224 VTAIL.n223 11.249
R336 VTAIL.n207 VTAIL.n184 11.249
R337 VTAIL.n437 VTAIL.n418 10.4732
R338 VTAIL.n459 VTAIL.n408 10.4732
R339 VTAIL.n31 VTAIL.n12 10.4732
R340 VTAIL.n53 VTAIL.n2 10.4732
R341 VTAIL.n89 VTAIL.n70 10.4732
R342 VTAIL.n111 VTAIL.n60 10.4732
R343 VTAIL.n147 VTAIL.n128 10.4732
R344 VTAIL.n169 VTAIL.n118 10.4732
R345 VTAIL.n401 VTAIL.n350 10.4732
R346 VTAIL.n380 VTAIL.n361 10.4732
R347 VTAIL.n343 VTAIL.n292 10.4732
R348 VTAIL.n322 VTAIL.n303 10.4732
R349 VTAIL.n285 VTAIL.n234 10.4732
R350 VTAIL.n264 VTAIL.n245 10.4732
R351 VTAIL.n227 VTAIL.n176 10.4732
R352 VTAIL.n206 VTAIL.n187 10.4732
R353 VTAIL.n425 VTAIL.n423 10.2747
R354 VTAIL.n19 VTAIL.n17 10.2747
R355 VTAIL.n77 VTAIL.n75 10.2747
R356 VTAIL.n135 VTAIL.n133 10.2747
R357 VTAIL.n368 VTAIL.n366 10.2747
R358 VTAIL.n310 VTAIL.n308 10.2747
R359 VTAIL.n252 VTAIL.n250 10.2747
R360 VTAIL.n194 VTAIL.n192 10.2747
R361 VTAIL.n434 VTAIL.n433 9.69747
R362 VTAIL.n460 VTAIL.n406 9.69747
R363 VTAIL.n28 VTAIL.n27 9.69747
R364 VTAIL.n54 VTAIL.n0 9.69747
R365 VTAIL.n86 VTAIL.n85 9.69747
R366 VTAIL.n112 VTAIL.n58 9.69747
R367 VTAIL.n144 VTAIL.n143 9.69747
R368 VTAIL.n170 VTAIL.n116 9.69747
R369 VTAIL.n402 VTAIL.n348 9.69747
R370 VTAIL.n377 VTAIL.n376 9.69747
R371 VTAIL.n344 VTAIL.n290 9.69747
R372 VTAIL.n319 VTAIL.n318 9.69747
R373 VTAIL.n286 VTAIL.n232 9.69747
R374 VTAIL.n261 VTAIL.n260 9.69747
R375 VTAIL.n228 VTAIL.n174 9.69747
R376 VTAIL.n203 VTAIL.n202 9.69747
R377 VTAIL.n462 VTAIL.n461 9.45567
R378 VTAIL.n56 VTAIL.n55 9.45567
R379 VTAIL.n114 VTAIL.n113 9.45567
R380 VTAIL.n172 VTAIL.n171 9.45567
R381 VTAIL.n404 VTAIL.n403 9.45567
R382 VTAIL.n346 VTAIL.n345 9.45567
R383 VTAIL.n288 VTAIL.n287 9.45567
R384 VTAIL.n230 VTAIL.n229 9.45567
R385 VTAIL.n461 VTAIL.n460 9.3005
R386 VTAIL.n408 VTAIL.n407 9.3005
R387 VTAIL.n455 VTAIL.n454 9.3005
R388 VTAIL.n453 VTAIL.n452 9.3005
R389 VTAIL.n412 VTAIL.n411 9.3005
R390 VTAIL.n427 VTAIL.n426 9.3005
R391 VTAIL.n429 VTAIL.n428 9.3005
R392 VTAIL.n420 VTAIL.n419 9.3005
R393 VTAIL.n435 VTAIL.n434 9.3005
R394 VTAIL.n437 VTAIL.n436 9.3005
R395 VTAIL.n416 VTAIL.n415 9.3005
R396 VTAIL.n444 VTAIL.n443 9.3005
R397 VTAIL.n446 VTAIL.n445 9.3005
R398 VTAIL.n55 VTAIL.n54 9.3005
R399 VTAIL.n2 VTAIL.n1 9.3005
R400 VTAIL.n49 VTAIL.n48 9.3005
R401 VTAIL.n47 VTAIL.n46 9.3005
R402 VTAIL.n6 VTAIL.n5 9.3005
R403 VTAIL.n21 VTAIL.n20 9.3005
R404 VTAIL.n23 VTAIL.n22 9.3005
R405 VTAIL.n14 VTAIL.n13 9.3005
R406 VTAIL.n29 VTAIL.n28 9.3005
R407 VTAIL.n31 VTAIL.n30 9.3005
R408 VTAIL.n10 VTAIL.n9 9.3005
R409 VTAIL.n38 VTAIL.n37 9.3005
R410 VTAIL.n40 VTAIL.n39 9.3005
R411 VTAIL.n113 VTAIL.n112 9.3005
R412 VTAIL.n60 VTAIL.n59 9.3005
R413 VTAIL.n107 VTAIL.n106 9.3005
R414 VTAIL.n105 VTAIL.n104 9.3005
R415 VTAIL.n64 VTAIL.n63 9.3005
R416 VTAIL.n79 VTAIL.n78 9.3005
R417 VTAIL.n81 VTAIL.n80 9.3005
R418 VTAIL.n72 VTAIL.n71 9.3005
R419 VTAIL.n87 VTAIL.n86 9.3005
R420 VTAIL.n89 VTAIL.n88 9.3005
R421 VTAIL.n68 VTAIL.n67 9.3005
R422 VTAIL.n96 VTAIL.n95 9.3005
R423 VTAIL.n98 VTAIL.n97 9.3005
R424 VTAIL.n171 VTAIL.n170 9.3005
R425 VTAIL.n118 VTAIL.n117 9.3005
R426 VTAIL.n165 VTAIL.n164 9.3005
R427 VTAIL.n163 VTAIL.n162 9.3005
R428 VTAIL.n122 VTAIL.n121 9.3005
R429 VTAIL.n137 VTAIL.n136 9.3005
R430 VTAIL.n139 VTAIL.n138 9.3005
R431 VTAIL.n130 VTAIL.n129 9.3005
R432 VTAIL.n145 VTAIL.n144 9.3005
R433 VTAIL.n147 VTAIL.n146 9.3005
R434 VTAIL.n126 VTAIL.n125 9.3005
R435 VTAIL.n154 VTAIL.n153 9.3005
R436 VTAIL.n156 VTAIL.n155 9.3005
R437 VTAIL.n370 VTAIL.n369 9.3005
R438 VTAIL.n372 VTAIL.n371 9.3005
R439 VTAIL.n363 VTAIL.n362 9.3005
R440 VTAIL.n378 VTAIL.n377 9.3005
R441 VTAIL.n380 VTAIL.n379 9.3005
R442 VTAIL.n358 VTAIL.n357 9.3005
R443 VTAIL.n386 VTAIL.n385 9.3005
R444 VTAIL.n388 VTAIL.n387 9.3005
R445 VTAIL.n403 VTAIL.n402 9.3005
R446 VTAIL.n350 VTAIL.n349 9.3005
R447 VTAIL.n397 VTAIL.n396 9.3005
R448 VTAIL.n395 VTAIL.n394 9.3005
R449 VTAIL.n354 VTAIL.n353 9.3005
R450 VTAIL.n312 VTAIL.n311 9.3005
R451 VTAIL.n314 VTAIL.n313 9.3005
R452 VTAIL.n305 VTAIL.n304 9.3005
R453 VTAIL.n320 VTAIL.n319 9.3005
R454 VTAIL.n322 VTAIL.n321 9.3005
R455 VTAIL.n300 VTAIL.n299 9.3005
R456 VTAIL.n328 VTAIL.n327 9.3005
R457 VTAIL.n330 VTAIL.n329 9.3005
R458 VTAIL.n345 VTAIL.n344 9.3005
R459 VTAIL.n292 VTAIL.n291 9.3005
R460 VTAIL.n339 VTAIL.n338 9.3005
R461 VTAIL.n337 VTAIL.n336 9.3005
R462 VTAIL.n296 VTAIL.n295 9.3005
R463 VTAIL.n254 VTAIL.n253 9.3005
R464 VTAIL.n256 VTAIL.n255 9.3005
R465 VTAIL.n247 VTAIL.n246 9.3005
R466 VTAIL.n262 VTAIL.n261 9.3005
R467 VTAIL.n264 VTAIL.n263 9.3005
R468 VTAIL.n242 VTAIL.n241 9.3005
R469 VTAIL.n270 VTAIL.n269 9.3005
R470 VTAIL.n272 VTAIL.n271 9.3005
R471 VTAIL.n287 VTAIL.n286 9.3005
R472 VTAIL.n234 VTAIL.n233 9.3005
R473 VTAIL.n281 VTAIL.n280 9.3005
R474 VTAIL.n279 VTAIL.n278 9.3005
R475 VTAIL.n238 VTAIL.n237 9.3005
R476 VTAIL.n196 VTAIL.n195 9.3005
R477 VTAIL.n198 VTAIL.n197 9.3005
R478 VTAIL.n189 VTAIL.n188 9.3005
R479 VTAIL.n204 VTAIL.n203 9.3005
R480 VTAIL.n206 VTAIL.n205 9.3005
R481 VTAIL.n184 VTAIL.n183 9.3005
R482 VTAIL.n212 VTAIL.n211 9.3005
R483 VTAIL.n214 VTAIL.n213 9.3005
R484 VTAIL.n229 VTAIL.n228 9.3005
R485 VTAIL.n176 VTAIL.n175 9.3005
R486 VTAIL.n223 VTAIL.n222 9.3005
R487 VTAIL.n221 VTAIL.n220 9.3005
R488 VTAIL.n180 VTAIL.n179 9.3005
R489 VTAIL.n430 VTAIL.n420 8.92171
R490 VTAIL.n24 VTAIL.n14 8.92171
R491 VTAIL.n82 VTAIL.n72 8.92171
R492 VTAIL.n140 VTAIL.n130 8.92171
R493 VTAIL.n373 VTAIL.n363 8.92171
R494 VTAIL.n315 VTAIL.n305 8.92171
R495 VTAIL.n257 VTAIL.n247 8.92171
R496 VTAIL.n199 VTAIL.n189 8.92171
R497 VTAIL.n429 VTAIL.n422 8.14595
R498 VTAIL.n23 VTAIL.n16 8.14595
R499 VTAIL.n81 VTAIL.n74 8.14595
R500 VTAIL.n139 VTAIL.n132 8.14595
R501 VTAIL.n372 VTAIL.n365 8.14595
R502 VTAIL.n314 VTAIL.n307 8.14595
R503 VTAIL.n256 VTAIL.n249 8.14595
R504 VTAIL.n198 VTAIL.n191 8.14595
R505 VTAIL.n426 VTAIL.n425 7.3702
R506 VTAIL.n20 VTAIL.n19 7.3702
R507 VTAIL.n78 VTAIL.n77 7.3702
R508 VTAIL.n136 VTAIL.n135 7.3702
R509 VTAIL.n369 VTAIL.n368 7.3702
R510 VTAIL.n311 VTAIL.n310 7.3702
R511 VTAIL.n253 VTAIL.n252 7.3702
R512 VTAIL.n195 VTAIL.n194 7.3702
R513 VTAIL.n426 VTAIL.n422 5.81868
R514 VTAIL.n20 VTAIL.n16 5.81868
R515 VTAIL.n78 VTAIL.n74 5.81868
R516 VTAIL.n136 VTAIL.n132 5.81868
R517 VTAIL.n369 VTAIL.n365 5.81868
R518 VTAIL.n311 VTAIL.n307 5.81868
R519 VTAIL.n253 VTAIL.n249 5.81868
R520 VTAIL.n195 VTAIL.n191 5.81868
R521 VTAIL.n430 VTAIL.n429 5.04292
R522 VTAIL.n24 VTAIL.n23 5.04292
R523 VTAIL.n82 VTAIL.n81 5.04292
R524 VTAIL.n140 VTAIL.n139 5.04292
R525 VTAIL.n373 VTAIL.n372 5.04292
R526 VTAIL.n315 VTAIL.n314 5.04292
R527 VTAIL.n257 VTAIL.n256 5.04292
R528 VTAIL.n199 VTAIL.n198 5.04292
R529 VTAIL.n433 VTAIL.n420 4.26717
R530 VTAIL.n462 VTAIL.n406 4.26717
R531 VTAIL.n27 VTAIL.n14 4.26717
R532 VTAIL.n56 VTAIL.n0 4.26717
R533 VTAIL.n85 VTAIL.n72 4.26717
R534 VTAIL.n114 VTAIL.n58 4.26717
R535 VTAIL.n143 VTAIL.n130 4.26717
R536 VTAIL.n172 VTAIL.n116 4.26717
R537 VTAIL.n404 VTAIL.n348 4.26717
R538 VTAIL.n376 VTAIL.n363 4.26717
R539 VTAIL.n346 VTAIL.n290 4.26717
R540 VTAIL.n318 VTAIL.n305 4.26717
R541 VTAIL.n288 VTAIL.n232 4.26717
R542 VTAIL.n260 VTAIL.n247 4.26717
R543 VTAIL.n230 VTAIL.n174 4.26717
R544 VTAIL.n202 VTAIL.n189 4.26717
R545 VTAIL.n434 VTAIL.n418 3.49141
R546 VTAIL.n460 VTAIL.n459 3.49141
R547 VTAIL.n28 VTAIL.n12 3.49141
R548 VTAIL.n54 VTAIL.n53 3.49141
R549 VTAIL.n86 VTAIL.n70 3.49141
R550 VTAIL.n112 VTAIL.n111 3.49141
R551 VTAIL.n144 VTAIL.n128 3.49141
R552 VTAIL.n170 VTAIL.n169 3.49141
R553 VTAIL.n402 VTAIL.n401 3.49141
R554 VTAIL.n377 VTAIL.n361 3.49141
R555 VTAIL.n344 VTAIL.n343 3.49141
R556 VTAIL.n319 VTAIL.n303 3.49141
R557 VTAIL.n286 VTAIL.n285 3.49141
R558 VTAIL.n261 VTAIL.n245 3.49141
R559 VTAIL.n228 VTAIL.n227 3.49141
R560 VTAIL.n203 VTAIL.n187 3.49141
R561 VTAIL.n289 VTAIL.n231 3.19016
R562 VTAIL.n405 VTAIL.n347 3.19016
R563 VTAIL.n173 VTAIL.n115 3.19016
R564 VTAIL.n427 VTAIL.n423 2.84303
R565 VTAIL.n21 VTAIL.n17 2.84303
R566 VTAIL.n79 VTAIL.n75 2.84303
R567 VTAIL.n137 VTAIL.n133 2.84303
R568 VTAIL.n370 VTAIL.n366 2.84303
R569 VTAIL.n312 VTAIL.n308 2.84303
R570 VTAIL.n254 VTAIL.n250 2.84303
R571 VTAIL.n196 VTAIL.n192 2.84303
R572 VTAIL.n438 VTAIL.n437 2.71565
R573 VTAIL.n456 VTAIL.n408 2.71565
R574 VTAIL.n32 VTAIL.n31 2.71565
R575 VTAIL.n50 VTAIL.n2 2.71565
R576 VTAIL.n90 VTAIL.n89 2.71565
R577 VTAIL.n108 VTAIL.n60 2.71565
R578 VTAIL.n148 VTAIL.n147 2.71565
R579 VTAIL.n166 VTAIL.n118 2.71565
R580 VTAIL.n398 VTAIL.n350 2.71565
R581 VTAIL.n381 VTAIL.n380 2.71565
R582 VTAIL.n340 VTAIL.n292 2.71565
R583 VTAIL.n323 VTAIL.n322 2.71565
R584 VTAIL.n282 VTAIL.n234 2.71565
R585 VTAIL.n265 VTAIL.n264 2.71565
R586 VTAIL.n224 VTAIL.n176 2.71565
R587 VTAIL.n207 VTAIL.n206 2.71565
R588 VTAIL.n442 VTAIL.n416 1.93989
R589 VTAIL.n455 VTAIL.n410 1.93989
R590 VTAIL.n36 VTAIL.n10 1.93989
R591 VTAIL.n49 VTAIL.n4 1.93989
R592 VTAIL.n94 VTAIL.n68 1.93989
R593 VTAIL.n107 VTAIL.n62 1.93989
R594 VTAIL.n152 VTAIL.n126 1.93989
R595 VTAIL.n165 VTAIL.n120 1.93989
R596 VTAIL.n397 VTAIL.n352 1.93989
R597 VTAIL.n384 VTAIL.n358 1.93989
R598 VTAIL.n339 VTAIL.n294 1.93989
R599 VTAIL.n326 VTAIL.n300 1.93989
R600 VTAIL.n281 VTAIL.n236 1.93989
R601 VTAIL.n268 VTAIL.n242 1.93989
R602 VTAIL.n223 VTAIL.n178 1.93989
R603 VTAIL.n210 VTAIL.n184 1.93989
R604 VTAIL VTAIL.n57 1.65352
R605 VTAIL VTAIL.n463 1.53714
R606 VTAIL.n443 VTAIL.n414 1.16414
R607 VTAIL.n452 VTAIL.n451 1.16414
R608 VTAIL.n37 VTAIL.n8 1.16414
R609 VTAIL.n46 VTAIL.n45 1.16414
R610 VTAIL.n95 VTAIL.n66 1.16414
R611 VTAIL.n104 VTAIL.n103 1.16414
R612 VTAIL.n153 VTAIL.n124 1.16414
R613 VTAIL.n162 VTAIL.n161 1.16414
R614 VTAIL.n394 VTAIL.n393 1.16414
R615 VTAIL.n385 VTAIL.n356 1.16414
R616 VTAIL.n336 VTAIL.n335 1.16414
R617 VTAIL.n327 VTAIL.n298 1.16414
R618 VTAIL.n278 VTAIL.n277 1.16414
R619 VTAIL.n269 VTAIL.n240 1.16414
R620 VTAIL.n220 VTAIL.n219 1.16414
R621 VTAIL.n211 VTAIL.n182 1.16414
R622 VTAIL.n347 VTAIL.n289 0.470328
R623 VTAIL.n115 VTAIL.n57 0.470328
R624 VTAIL.n447 VTAIL.n446 0.388379
R625 VTAIL.n448 VTAIL.n412 0.388379
R626 VTAIL.n41 VTAIL.n40 0.388379
R627 VTAIL.n42 VTAIL.n6 0.388379
R628 VTAIL.n99 VTAIL.n98 0.388379
R629 VTAIL.n100 VTAIL.n64 0.388379
R630 VTAIL.n157 VTAIL.n156 0.388379
R631 VTAIL.n158 VTAIL.n122 0.388379
R632 VTAIL.n390 VTAIL.n354 0.388379
R633 VTAIL.n389 VTAIL.n388 0.388379
R634 VTAIL.n332 VTAIL.n296 0.388379
R635 VTAIL.n331 VTAIL.n330 0.388379
R636 VTAIL.n274 VTAIL.n238 0.388379
R637 VTAIL.n273 VTAIL.n272 0.388379
R638 VTAIL.n216 VTAIL.n180 0.388379
R639 VTAIL.n215 VTAIL.n214 0.388379
R640 VTAIL.n428 VTAIL.n427 0.155672
R641 VTAIL.n428 VTAIL.n419 0.155672
R642 VTAIL.n435 VTAIL.n419 0.155672
R643 VTAIL.n436 VTAIL.n435 0.155672
R644 VTAIL.n436 VTAIL.n415 0.155672
R645 VTAIL.n444 VTAIL.n415 0.155672
R646 VTAIL.n445 VTAIL.n444 0.155672
R647 VTAIL.n445 VTAIL.n411 0.155672
R648 VTAIL.n453 VTAIL.n411 0.155672
R649 VTAIL.n454 VTAIL.n453 0.155672
R650 VTAIL.n454 VTAIL.n407 0.155672
R651 VTAIL.n461 VTAIL.n407 0.155672
R652 VTAIL.n22 VTAIL.n21 0.155672
R653 VTAIL.n22 VTAIL.n13 0.155672
R654 VTAIL.n29 VTAIL.n13 0.155672
R655 VTAIL.n30 VTAIL.n29 0.155672
R656 VTAIL.n30 VTAIL.n9 0.155672
R657 VTAIL.n38 VTAIL.n9 0.155672
R658 VTAIL.n39 VTAIL.n38 0.155672
R659 VTAIL.n39 VTAIL.n5 0.155672
R660 VTAIL.n47 VTAIL.n5 0.155672
R661 VTAIL.n48 VTAIL.n47 0.155672
R662 VTAIL.n48 VTAIL.n1 0.155672
R663 VTAIL.n55 VTAIL.n1 0.155672
R664 VTAIL.n80 VTAIL.n79 0.155672
R665 VTAIL.n80 VTAIL.n71 0.155672
R666 VTAIL.n87 VTAIL.n71 0.155672
R667 VTAIL.n88 VTAIL.n87 0.155672
R668 VTAIL.n88 VTAIL.n67 0.155672
R669 VTAIL.n96 VTAIL.n67 0.155672
R670 VTAIL.n97 VTAIL.n96 0.155672
R671 VTAIL.n97 VTAIL.n63 0.155672
R672 VTAIL.n105 VTAIL.n63 0.155672
R673 VTAIL.n106 VTAIL.n105 0.155672
R674 VTAIL.n106 VTAIL.n59 0.155672
R675 VTAIL.n113 VTAIL.n59 0.155672
R676 VTAIL.n138 VTAIL.n137 0.155672
R677 VTAIL.n138 VTAIL.n129 0.155672
R678 VTAIL.n145 VTAIL.n129 0.155672
R679 VTAIL.n146 VTAIL.n145 0.155672
R680 VTAIL.n146 VTAIL.n125 0.155672
R681 VTAIL.n154 VTAIL.n125 0.155672
R682 VTAIL.n155 VTAIL.n154 0.155672
R683 VTAIL.n155 VTAIL.n121 0.155672
R684 VTAIL.n163 VTAIL.n121 0.155672
R685 VTAIL.n164 VTAIL.n163 0.155672
R686 VTAIL.n164 VTAIL.n117 0.155672
R687 VTAIL.n171 VTAIL.n117 0.155672
R688 VTAIL.n403 VTAIL.n349 0.155672
R689 VTAIL.n396 VTAIL.n349 0.155672
R690 VTAIL.n396 VTAIL.n395 0.155672
R691 VTAIL.n395 VTAIL.n353 0.155672
R692 VTAIL.n387 VTAIL.n353 0.155672
R693 VTAIL.n387 VTAIL.n386 0.155672
R694 VTAIL.n386 VTAIL.n357 0.155672
R695 VTAIL.n379 VTAIL.n357 0.155672
R696 VTAIL.n379 VTAIL.n378 0.155672
R697 VTAIL.n378 VTAIL.n362 0.155672
R698 VTAIL.n371 VTAIL.n362 0.155672
R699 VTAIL.n371 VTAIL.n370 0.155672
R700 VTAIL.n345 VTAIL.n291 0.155672
R701 VTAIL.n338 VTAIL.n291 0.155672
R702 VTAIL.n338 VTAIL.n337 0.155672
R703 VTAIL.n337 VTAIL.n295 0.155672
R704 VTAIL.n329 VTAIL.n295 0.155672
R705 VTAIL.n329 VTAIL.n328 0.155672
R706 VTAIL.n328 VTAIL.n299 0.155672
R707 VTAIL.n321 VTAIL.n299 0.155672
R708 VTAIL.n321 VTAIL.n320 0.155672
R709 VTAIL.n320 VTAIL.n304 0.155672
R710 VTAIL.n313 VTAIL.n304 0.155672
R711 VTAIL.n313 VTAIL.n312 0.155672
R712 VTAIL.n287 VTAIL.n233 0.155672
R713 VTAIL.n280 VTAIL.n233 0.155672
R714 VTAIL.n280 VTAIL.n279 0.155672
R715 VTAIL.n279 VTAIL.n237 0.155672
R716 VTAIL.n271 VTAIL.n237 0.155672
R717 VTAIL.n271 VTAIL.n270 0.155672
R718 VTAIL.n270 VTAIL.n241 0.155672
R719 VTAIL.n263 VTAIL.n241 0.155672
R720 VTAIL.n263 VTAIL.n262 0.155672
R721 VTAIL.n262 VTAIL.n246 0.155672
R722 VTAIL.n255 VTAIL.n246 0.155672
R723 VTAIL.n255 VTAIL.n254 0.155672
R724 VTAIL.n229 VTAIL.n175 0.155672
R725 VTAIL.n222 VTAIL.n175 0.155672
R726 VTAIL.n222 VTAIL.n221 0.155672
R727 VTAIL.n221 VTAIL.n179 0.155672
R728 VTAIL.n213 VTAIL.n179 0.155672
R729 VTAIL.n213 VTAIL.n212 0.155672
R730 VTAIL.n212 VTAIL.n183 0.155672
R731 VTAIL.n205 VTAIL.n183 0.155672
R732 VTAIL.n205 VTAIL.n204 0.155672
R733 VTAIL.n204 VTAIL.n188 0.155672
R734 VTAIL.n197 VTAIL.n188 0.155672
R735 VTAIL.n197 VTAIL.n196 0.155672
R736 VDD1 VDD1.n1 109.204
R737 VDD1 VDD1.n0 66.0832
R738 VDD1.n0 VDD1.t0 1.82203
R739 VDD1.n0 VDD1.t1 1.82203
R740 VDD1.n1 VDD1.t2 1.82203
R741 VDD1.n1 VDD1.t3 1.82203
R742 B.n765 B.n764 585
R743 B.n292 B.n119 585
R744 B.n291 B.n290 585
R745 B.n289 B.n288 585
R746 B.n287 B.n286 585
R747 B.n285 B.n284 585
R748 B.n283 B.n282 585
R749 B.n281 B.n280 585
R750 B.n279 B.n278 585
R751 B.n277 B.n276 585
R752 B.n275 B.n274 585
R753 B.n273 B.n272 585
R754 B.n271 B.n270 585
R755 B.n269 B.n268 585
R756 B.n267 B.n266 585
R757 B.n265 B.n264 585
R758 B.n263 B.n262 585
R759 B.n261 B.n260 585
R760 B.n259 B.n258 585
R761 B.n257 B.n256 585
R762 B.n255 B.n254 585
R763 B.n253 B.n252 585
R764 B.n251 B.n250 585
R765 B.n249 B.n248 585
R766 B.n247 B.n246 585
R767 B.n245 B.n244 585
R768 B.n243 B.n242 585
R769 B.n241 B.n240 585
R770 B.n239 B.n238 585
R771 B.n237 B.n236 585
R772 B.n235 B.n234 585
R773 B.n233 B.n232 585
R774 B.n231 B.n230 585
R775 B.n229 B.n228 585
R776 B.n227 B.n226 585
R777 B.n225 B.n224 585
R778 B.n223 B.n222 585
R779 B.n221 B.n220 585
R780 B.n219 B.n218 585
R781 B.n217 B.n216 585
R782 B.n215 B.n214 585
R783 B.n213 B.n212 585
R784 B.n211 B.n210 585
R785 B.n209 B.n208 585
R786 B.n207 B.n206 585
R787 B.n205 B.n204 585
R788 B.n203 B.n202 585
R789 B.n201 B.n200 585
R790 B.n199 B.n198 585
R791 B.n197 B.n196 585
R792 B.n195 B.n194 585
R793 B.n193 B.n192 585
R794 B.n191 B.n190 585
R795 B.n189 B.n188 585
R796 B.n187 B.n186 585
R797 B.n185 B.n184 585
R798 B.n183 B.n182 585
R799 B.n181 B.n180 585
R800 B.n179 B.n178 585
R801 B.n177 B.n176 585
R802 B.n175 B.n174 585
R803 B.n173 B.n172 585
R804 B.n171 B.n170 585
R805 B.n169 B.n168 585
R806 B.n167 B.n166 585
R807 B.n165 B.n164 585
R808 B.n163 B.n162 585
R809 B.n161 B.n160 585
R810 B.n159 B.n158 585
R811 B.n157 B.n156 585
R812 B.n155 B.n154 585
R813 B.n153 B.n152 585
R814 B.n151 B.n150 585
R815 B.n149 B.n148 585
R816 B.n147 B.n146 585
R817 B.n145 B.n144 585
R818 B.n143 B.n142 585
R819 B.n141 B.n140 585
R820 B.n139 B.n138 585
R821 B.n137 B.n136 585
R822 B.n135 B.n134 585
R823 B.n133 B.n132 585
R824 B.n131 B.n130 585
R825 B.n129 B.n128 585
R826 B.n127 B.n126 585
R827 B.n75 B.n74 585
R828 B.n763 B.n76 585
R829 B.n768 B.n76 585
R830 B.n762 B.n761 585
R831 B.n761 B.n72 585
R832 B.n760 B.n71 585
R833 B.n774 B.n71 585
R834 B.n759 B.n70 585
R835 B.n775 B.n70 585
R836 B.n758 B.n69 585
R837 B.n776 B.n69 585
R838 B.n757 B.n756 585
R839 B.n756 B.n65 585
R840 B.n755 B.n64 585
R841 B.n782 B.n64 585
R842 B.n754 B.n63 585
R843 B.n783 B.n63 585
R844 B.n753 B.n62 585
R845 B.n784 B.n62 585
R846 B.n752 B.n751 585
R847 B.n751 B.n58 585
R848 B.n750 B.n57 585
R849 B.n790 B.n57 585
R850 B.n749 B.n56 585
R851 B.n791 B.n56 585
R852 B.n748 B.n55 585
R853 B.n792 B.n55 585
R854 B.n747 B.n746 585
R855 B.n746 B.n51 585
R856 B.n745 B.n50 585
R857 B.n798 B.n50 585
R858 B.n744 B.n49 585
R859 B.n799 B.n49 585
R860 B.n743 B.n48 585
R861 B.n800 B.n48 585
R862 B.n742 B.n741 585
R863 B.n741 B.n44 585
R864 B.n740 B.n43 585
R865 B.n806 B.n43 585
R866 B.n739 B.n42 585
R867 B.n807 B.n42 585
R868 B.n738 B.n41 585
R869 B.n808 B.n41 585
R870 B.n737 B.n736 585
R871 B.n736 B.n37 585
R872 B.n735 B.n36 585
R873 B.n814 B.n36 585
R874 B.n734 B.n35 585
R875 B.n815 B.n35 585
R876 B.n733 B.n34 585
R877 B.n816 B.n34 585
R878 B.n732 B.n731 585
R879 B.n731 B.n30 585
R880 B.n730 B.n29 585
R881 B.n822 B.n29 585
R882 B.n729 B.n28 585
R883 B.n823 B.n28 585
R884 B.n728 B.n27 585
R885 B.n824 B.n27 585
R886 B.n727 B.n726 585
R887 B.n726 B.n23 585
R888 B.n725 B.n22 585
R889 B.n830 B.n22 585
R890 B.n724 B.n21 585
R891 B.n831 B.n21 585
R892 B.n723 B.n20 585
R893 B.n832 B.n20 585
R894 B.n722 B.n721 585
R895 B.n721 B.n19 585
R896 B.n720 B.n15 585
R897 B.n838 B.n15 585
R898 B.n719 B.n14 585
R899 B.n839 B.n14 585
R900 B.n718 B.n13 585
R901 B.n840 B.n13 585
R902 B.n717 B.n716 585
R903 B.n716 B.n12 585
R904 B.n715 B.n714 585
R905 B.n715 B.n8 585
R906 B.n713 B.n7 585
R907 B.n847 B.n7 585
R908 B.n712 B.n6 585
R909 B.n848 B.n6 585
R910 B.n711 B.n5 585
R911 B.n849 B.n5 585
R912 B.n710 B.n709 585
R913 B.n709 B.n4 585
R914 B.n708 B.n293 585
R915 B.n708 B.n707 585
R916 B.n698 B.n294 585
R917 B.n295 B.n294 585
R918 B.n700 B.n699 585
R919 B.n701 B.n700 585
R920 B.n697 B.n300 585
R921 B.n300 B.n299 585
R922 B.n696 B.n695 585
R923 B.n695 B.n694 585
R924 B.n302 B.n301 585
R925 B.n687 B.n302 585
R926 B.n686 B.n685 585
R927 B.n688 B.n686 585
R928 B.n684 B.n307 585
R929 B.n307 B.n306 585
R930 B.n683 B.n682 585
R931 B.n682 B.n681 585
R932 B.n309 B.n308 585
R933 B.n310 B.n309 585
R934 B.n674 B.n673 585
R935 B.n675 B.n674 585
R936 B.n672 B.n315 585
R937 B.n315 B.n314 585
R938 B.n671 B.n670 585
R939 B.n670 B.n669 585
R940 B.n317 B.n316 585
R941 B.n318 B.n317 585
R942 B.n662 B.n661 585
R943 B.n663 B.n662 585
R944 B.n660 B.n323 585
R945 B.n323 B.n322 585
R946 B.n659 B.n658 585
R947 B.n658 B.n657 585
R948 B.n325 B.n324 585
R949 B.n326 B.n325 585
R950 B.n650 B.n649 585
R951 B.n651 B.n650 585
R952 B.n648 B.n331 585
R953 B.n331 B.n330 585
R954 B.n647 B.n646 585
R955 B.n646 B.n645 585
R956 B.n333 B.n332 585
R957 B.n334 B.n333 585
R958 B.n638 B.n637 585
R959 B.n639 B.n638 585
R960 B.n636 B.n339 585
R961 B.n339 B.n338 585
R962 B.n635 B.n634 585
R963 B.n634 B.n633 585
R964 B.n341 B.n340 585
R965 B.n342 B.n341 585
R966 B.n626 B.n625 585
R967 B.n627 B.n626 585
R968 B.n624 B.n347 585
R969 B.n347 B.n346 585
R970 B.n623 B.n622 585
R971 B.n622 B.n621 585
R972 B.n349 B.n348 585
R973 B.n350 B.n349 585
R974 B.n614 B.n613 585
R975 B.n615 B.n614 585
R976 B.n612 B.n355 585
R977 B.n355 B.n354 585
R978 B.n611 B.n610 585
R979 B.n610 B.n609 585
R980 B.n357 B.n356 585
R981 B.n358 B.n357 585
R982 B.n602 B.n601 585
R983 B.n603 B.n602 585
R984 B.n600 B.n363 585
R985 B.n363 B.n362 585
R986 B.n599 B.n598 585
R987 B.n598 B.n597 585
R988 B.n365 B.n364 585
R989 B.n366 B.n365 585
R990 B.n590 B.n589 585
R991 B.n591 B.n590 585
R992 B.n369 B.n368 585
R993 B.n418 B.n416 585
R994 B.n419 B.n415 585
R995 B.n419 B.n370 585
R996 B.n422 B.n421 585
R997 B.n423 B.n414 585
R998 B.n425 B.n424 585
R999 B.n427 B.n413 585
R1000 B.n430 B.n429 585
R1001 B.n431 B.n412 585
R1002 B.n433 B.n432 585
R1003 B.n435 B.n411 585
R1004 B.n438 B.n437 585
R1005 B.n439 B.n410 585
R1006 B.n441 B.n440 585
R1007 B.n443 B.n409 585
R1008 B.n446 B.n445 585
R1009 B.n447 B.n408 585
R1010 B.n449 B.n448 585
R1011 B.n451 B.n407 585
R1012 B.n454 B.n453 585
R1013 B.n455 B.n406 585
R1014 B.n457 B.n456 585
R1015 B.n459 B.n405 585
R1016 B.n462 B.n461 585
R1017 B.n463 B.n404 585
R1018 B.n465 B.n464 585
R1019 B.n467 B.n403 585
R1020 B.n470 B.n469 585
R1021 B.n471 B.n402 585
R1022 B.n473 B.n472 585
R1023 B.n475 B.n401 585
R1024 B.n478 B.n477 585
R1025 B.n479 B.n400 585
R1026 B.n481 B.n480 585
R1027 B.n483 B.n399 585
R1028 B.n486 B.n485 585
R1029 B.n487 B.n398 585
R1030 B.n492 B.n491 585
R1031 B.n494 B.n397 585
R1032 B.n497 B.n496 585
R1033 B.n498 B.n396 585
R1034 B.n500 B.n499 585
R1035 B.n502 B.n395 585
R1036 B.n505 B.n504 585
R1037 B.n506 B.n394 585
R1038 B.n508 B.n507 585
R1039 B.n510 B.n393 585
R1040 B.n513 B.n512 585
R1041 B.n515 B.n390 585
R1042 B.n517 B.n516 585
R1043 B.n519 B.n389 585
R1044 B.n522 B.n521 585
R1045 B.n523 B.n388 585
R1046 B.n525 B.n524 585
R1047 B.n527 B.n387 585
R1048 B.n530 B.n529 585
R1049 B.n531 B.n386 585
R1050 B.n533 B.n532 585
R1051 B.n535 B.n385 585
R1052 B.n538 B.n537 585
R1053 B.n539 B.n384 585
R1054 B.n541 B.n540 585
R1055 B.n543 B.n383 585
R1056 B.n546 B.n545 585
R1057 B.n547 B.n382 585
R1058 B.n549 B.n548 585
R1059 B.n551 B.n381 585
R1060 B.n554 B.n553 585
R1061 B.n555 B.n380 585
R1062 B.n557 B.n556 585
R1063 B.n559 B.n379 585
R1064 B.n562 B.n561 585
R1065 B.n563 B.n378 585
R1066 B.n565 B.n564 585
R1067 B.n567 B.n377 585
R1068 B.n570 B.n569 585
R1069 B.n571 B.n376 585
R1070 B.n573 B.n572 585
R1071 B.n575 B.n375 585
R1072 B.n578 B.n577 585
R1073 B.n579 B.n374 585
R1074 B.n581 B.n580 585
R1075 B.n583 B.n373 585
R1076 B.n584 B.n372 585
R1077 B.n587 B.n586 585
R1078 B.n588 B.n371 585
R1079 B.n371 B.n370 585
R1080 B.n593 B.n592 585
R1081 B.n592 B.n591 585
R1082 B.n594 B.n367 585
R1083 B.n367 B.n366 585
R1084 B.n596 B.n595 585
R1085 B.n597 B.n596 585
R1086 B.n361 B.n360 585
R1087 B.n362 B.n361 585
R1088 B.n605 B.n604 585
R1089 B.n604 B.n603 585
R1090 B.n606 B.n359 585
R1091 B.n359 B.n358 585
R1092 B.n608 B.n607 585
R1093 B.n609 B.n608 585
R1094 B.n353 B.n352 585
R1095 B.n354 B.n353 585
R1096 B.n617 B.n616 585
R1097 B.n616 B.n615 585
R1098 B.n618 B.n351 585
R1099 B.n351 B.n350 585
R1100 B.n620 B.n619 585
R1101 B.n621 B.n620 585
R1102 B.n345 B.n344 585
R1103 B.n346 B.n345 585
R1104 B.n629 B.n628 585
R1105 B.n628 B.n627 585
R1106 B.n630 B.n343 585
R1107 B.n343 B.n342 585
R1108 B.n632 B.n631 585
R1109 B.n633 B.n632 585
R1110 B.n337 B.n336 585
R1111 B.n338 B.n337 585
R1112 B.n641 B.n640 585
R1113 B.n640 B.n639 585
R1114 B.n642 B.n335 585
R1115 B.n335 B.n334 585
R1116 B.n644 B.n643 585
R1117 B.n645 B.n644 585
R1118 B.n329 B.n328 585
R1119 B.n330 B.n329 585
R1120 B.n653 B.n652 585
R1121 B.n652 B.n651 585
R1122 B.n654 B.n327 585
R1123 B.n327 B.n326 585
R1124 B.n656 B.n655 585
R1125 B.n657 B.n656 585
R1126 B.n321 B.n320 585
R1127 B.n322 B.n321 585
R1128 B.n665 B.n664 585
R1129 B.n664 B.n663 585
R1130 B.n666 B.n319 585
R1131 B.n319 B.n318 585
R1132 B.n668 B.n667 585
R1133 B.n669 B.n668 585
R1134 B.n313 B.n312 585
R1135 B.n314 B.n313 585
R1136 B.n677 B.n676 585
R1137 B.n676 B.n675 585
R1138 B.n678 B.n311 585
R1139 B.n311 B.n310 585
R1140 B.n680 B.n679 585
R1141 B.n681 B.n680 585
R1142 B.n305 B.n304 585
R1143 B.n306 B.n305 585
R1144 B.n690 B.n689 585
R1145 B.n689 B.n688 585
R1146 B.n691 B.n303 585
R1147 B.n687 B.n303 585
R1148 B.n693 B.n692 585
R1149 B.n694 B.n693 585
R1150 B.n298 B.n297 585
R1151 B.n299 B.n298 585
R1152 B.n703 B.n702 585
R1153 B.n702 B.n701 585
R1154 B.n704 B.n296 585
R1155 B.n296 B.n295 585
R1156 B.n706 B.n705 585
R1157 B.n707 B.n706 585
R1158 B.n3 B.n0 585
R1159 B.n4 B.n3 585
R1160 B.n846 B.n1 585
R1161 B.n847 B.n846 585
R1162 B.n845 B.n844 585
R1163 B.n845 B.n8 585
R1164 B.n843 B.n9 585
R1165 B.n12 B.n9 585
R1166 B.n842 B.n841 585
R1167 B.n841 B.n840 585
R1168 B.n11 B.n10 585
R1169 B.n839 B.n11 585
R1170 B.n837 B.n836 585
R1171 B.n838 B.n837 585
R1172 B.n835 B.n16 585
R1173 B.n19 B.n16 585
R1174 B.n834 B.n833 585
R1175 B.n833 B.n832 585
R1176 B.n18 B.n17 585
R1177 B.n831 B.n18 585
R1178 B.n829 B.n828 585
R1179 B.n830 B.n829 585
R1180 B.n827 B.n24 585
R1181 B.n24 B.n23 585
R1182 B.n826 B.n825 585
R1183 B.n825 B.n824 585
R1184 B.n26 B.n25 585
R1185 B.n823 B.n26 585
R1186 B.n821 B.n820 585
R1187 B.n822 B.n821 585
R1188 B.n819 B.n31 585
R1189 B.n31 B.n30 585
R1190 B.n818 B.n817 585
R1191 B.n817 B.n816 585
R1192 B.n33 B.n32 585
R1193 B.n815 B.n33 585
R1194 B.n813 B.n812 585
R1195 B.n814 B.n813 585
R1196 B.n811 B.n38 585
R1197 B.n38 B.n37 585
R1198 B.n810 B.n809 585
R1199 B.n809 B.n808 585
R1200 B.n40 B.n39 585
R1201 B.n807 B.n40 585
R1202 B.n805 B.n804 585
R1203 B.n806 B.n805 585
R1204 B.n803 B.n45 585
R1205 B.n45 B.n44 585
R1206 B.n802 B.n801 585
R1207 B.n801 B.n800 585
R1208 B.n47 B.n46 585
R1209 B.n799 B.n47 585
R1210 B.n797 B.n796 585
R1211 B.n798 B.n797 585
R1212 B.n795 B.n52 585
R1213 B.n52 B.n51 585
R1214 B.n794 B.n793 585
R1215 B.n793 B.n792 585
R1216 B.n54 B.n53 585
R1217 B.n791 B.n54 585
R1218 B.n789 B.n788 585
R1219 B.n790 B.n789 585
R1220 B.n787 B.n59 585
R1221 B.n59 B.n58 585
R1222 B.n786 B.n785 585
R1223 B.n785 B.n784 585
R1224 B.n61 B.n60 585
R1225 B.n783 B.n61 585
R1226 B.n781 B.n780 585
R1227 B.n782 B.n781 585
R1228 B.n779 B.n66 585
R1229 B.n66 B.n65 585
R1230 B.n778 B.n777 585
R1231 B.n777 B.n776 585
R1232 B.n68 B.n67 585
R1233 B.n775 B.n68 585
R1234 B.n773 B.n772 585
R1235 B.n774 B.n773 585
R1236 B.n771 B.n73 585
R1237 B.n73 B.n72 585
R1238 B.n770 B.n769 585
R1239 B.n769 B.n768 585
R1240 B.n850 B.n849 585
R1241 B.n848 B.n2 585
R1242 B.n769 B.n75 554.963
R1243 B.n765 B.n76 554.963
R1244 B.n590 B.n371 554.963
R1245 B.n592 B.n369 554.963
R1246 B.n120 B.t13 334.801
R1247 B.n391 B.t7 334.801
R1248 B.n123 B.t16 334.801
R1249 B.n488 B.t10 334.801
R1250 B.n123 B.t15 286.709
R1251 B.n120 B.t11 286.709
R1252 B.n391 B.t4 286.709
R1253 B.n488 B.t8 286.709
R1254 B.n121 B.t14 263.045
R1255 B.n392 B.t6 263.045
R1256 B.n124 B.t17 263.045
R1257 B.n489 B.t9 263.045
R1258 B.n767 B.n766 256.663
R1259 B.n767 B.n118 256.663
R1260 B.n767 B.n117 256.663
R1261 B.n767 B.n116 256.663
R1262 B.n767 B.n115 256.663
R1263 B.n767 B.n114 256.663
R1264 B.n767 B.n113 256.663
R1265 B.n767 B.n112 256.663
R1266 B.n767 B.n111 256.663
R1267 B.n767 B.n110 256.663
R1268 B.n767 B.n109 256.663
R1269 B.n767 B.n108 256.663
R1270 B.n767 B.n107 256.663
R1271 B.n767 B.n106 256.663
R1272 B.n767 B.n105 256.663
R1273 B.n767 B.n104 256.663
R1274 B.n767 B.n103 256.663
R1275 B.n767 B.n102 256.663
R1276 B.n767 B.n101 256.663
R1277 B.n767 B.n100 256.663
R1278 B.n767 B.n99 256.663
R1279 B.n767 B.n98 256.663
R1280 B.n767 B.n97 256.663
R1281 B.n767 B.n96 256.663
R1282 B.n767 B.n95 256.663
R1283 B.n767 B.n94 256.663
R1284 B.n767 B.n93 256.663
R1285 B.n767 B.n92 256.663
R1286 B.n767 B.n91 256.663
R1287 B.n767 B.n90 256.663
R1288 B.n767 B.n89 256.663
R1289 B.n767 B.n88 256.663
R1290 B.n767 B.n87 256.663
R1291 B.n767 B.n86 256.663
R1292 B.n767 B.n85 256.663
R1293 B.n767 B.n84 256.663
R1294 B.n767 B.n83 256.663
R1295 B.n767 B.n82 256.663
R1296 B.n767 B.n81 256.663
R1297 B.n767 B.n80 256.663
R1298 B.n767 B.n79 256.663
R1299 B.n767 B.n78 256.663
R1300 B.n767 B.n77 256.663
R1301 B.n417 B.n370 256.663
R1302 B.n420 B.n370 256.663
R1303 B.n426 B.n370 256.663
R1304 B.n428 B.n370 256.663
R1305 B.n434 B.n370 256.663
R1306 B.n436 B.n370 256.663
R1307 B.n442 B.n370 256.663
R1308 B.n444 B.n370 256.663
R1309 B.n450 B.n370 256.663
R1310 B.n452 B.n370 256.663
R1311 B.n458 B.n370 256.663
R1312 B.n460 B.n370 256.663
R1313 B.n466 B.n370 256.663
R1314 B.n468 B.n370 256.663
R1315 B.n474 B.n370 256.663
R1316 B.n476 B.n370 256.663
R1317 B.n482 B.n370 256.663
R1318 B.n484 B.n370 256.663
R1319 B.n493 B.n370 256.663
R1320 B.n495 B.n370 256.663
R1321 B.n501 B.n370 256.663
R1322 B.n503 B.n370 256.663
R1323 B.n509 B.n370 256.663
R1324 B.n511 B.n370 256.663
R1325 B.n518 B.n370 256.663
R1326 B.n520 B.n370 256.663
R1327 B.n526 B.n370 256.663
R1328 B.n528 B.n370 256.663
R1329 B.n534 B.n370 256.663
R1330 B.n536 B.n370 256.663
R1331 B.n542 B.n370 256.663
R1332 B.n544 B.n370 256.663
R1333 B.n550 B.n370 256.663
R1334 B.n552 B.n370 256.663
R1335 B.n558 B.n370 256.663
R1336 B.n560 B.n370 256.663
R1337 B.n566 B.n370 256.663
R1338 B.n568 B.n370 256.663
R1339 B.n574 B.n370 256.663
R1340 B.n576 B.n370 256.663
R1341 B.n582 B.n370 256.663
R1342 B.n585 B.n370 256.663
R1343 B.n852 B.n851 256.663
R1344 B.n128 B.n127 163.367
R1345 B.n132 B.n131 163.367
R1346 B.n136 B.n135 163.367
R1347 B.n140 B.n139 163.367
R1348 B.n144 B.n143 163.367
R1349 B.n148 B.n147 163.367
R1350 B.n152 B.n151 163.367
R1351 B.n156 B.n155 163.367
R1352 B.n160 B.n159 163.367
R1353 B.n164 B.n163 163.367
R1354 B.n168 B.n167 163.367
R1355 B.n172 B.n171 163.367
R1356 B.n176 B.n175 163.367
R1357 B.n180 B.n179 163.367
R1358 B.n184 B.n183 163.367
R1359 B.n188 B.n187 163.367
R1360 B.n192 B.n191 163.367
R1361 B.n196 B.n195 163.367
R1362 B.n200 B.n199 163.367
R1363 B.n204 B.n203 163.367
R1364 B.n208 B.n207 163.367
R1365 B.n212 B.n211 163.367
R1366 B.n216 B.n215 163.367
R1367 B.n220 B.n219 163.367
R1368 B.n224 B.n223 163.367
R1369 B.n228 B.n227 163.367
R1370 B.n232 B.n231 163.367
R1371 B.n236 B.n235 163.367
R1372 B.n240 B.n239 163.367
R1373 B.n244 B.n243 163.367
R1374 B.n248 B.n247 163.367
R1375 B.n252 B.n251 163.367
R1376 B.n256 B.n255 163.367
R1377 B.n260 B.n259 163.367
R1378 B.n264 B.n263 163.367
R1379 B.n268 B.n267 163.367
R1380 B.n272 B.n271 163.367
R1381 B.n276 B.n275 163.367
R1382 B.n280 B.n279 163.367
R1383 B.n284 B.n283 163.367
R1384 B.n288 B.n287 163.367
R1385 B.n290 B.n119 163.367
R1386 B.n590 B.n365 163.367
R1387 B.n598 B.n365 163.367
R1388 B.n598 B.n363 163.367
R1389 B.n602 B.n363 163.367
R1390 B.n602 B.n357 163.367
R1391 B.n610 B.n357 163.367
R1392 B.n610 B.n355 163.367
R1393 B.n614 B.n355 163.367
R1394 B.n614 B.n349 163.367
R1395 B.n622 B.n349 163.367
R1396 B.n622 B.n347 163.367
R1397 B.n626 B.n347 163.367
R1398 B.n626 B.n341 163.367
R1399 B.n634 B.n341 163.367
R1400 B.n634 B.n339 163.367
R1401 B.n638 B.n339 163.367
R1402 B.n638 B.n333 163.367
R1403 B.n646 B.n333 163.367
R1404 B.n646 B.n331 163.367
R1405 B.n650 B.n331 163.367
R1406 B.n650 B.n325 163.367
R1407 B.n658 B.n325 163.367
R1408 B.n658 B.n323 163.367
R1409 B.n662 B.n323 163.367
R1410 B.n662 B.n317 163.367
R1411 B.n670 B.n317 163.367
R1412 B.n670 B.n315 163.367
R1413 B.n674 B.n315 163.367
R1414 B.n674 B.n309 163.367
R1415 B.n682 B.n309 163.367
R1416 B.n682 B.n307 163.367
R1417 B.n686 B.n307 163.367
R1418 B.n686 B.n302 163.367
R1419 B.n695 B.n302 163.367
R1420 B.n695 B.n300 163.367
R1421 B.n700 B.n300 163.367
R1422 B.n700 B.n294 163.367
R1423 B.n708 B.n294 163.367
R1424 B.n709 B.n708 163.367
R1425 B.n709 B.n5 163.367
R1426 B.n6 B.n5 163.367
R1427 B.n7 B.n6 163.367
R1428 B.n715 B.n7 163.367
R1429 B.n716 B.n715 163.367
R1430 B.n716 B.n13 163.367
R1431 B.n14 B.n13 163.367
R1432 B.n15 B.n14 163.367
R1433 B.n721 B.n15 163.367
R1434 B.n721 B.n20 163.367
R1435 B.n21 B.n20 163.367
R1436 B.n22 B.n21 163.367
R1437 B.n726 B.n22 163.367
R1438 B.n726 B.n27 163.367
R1439 B.n28 B.n27 163.367
R1440 B.n29 B.n28 163.367
R1441 B.n731 B.n29 163.367
R1442 B.n731 B.n34 163.367
R1443 B.n35 B.n34 163.367
R1444 B.n36 B.n35 163.367
R1445 B.n736 B.n36 163.367
R1446 B.n736 B.n41 163.367
R1447 B.n42 B.n41 163.367
R1448 B.n43 B.n42 163.367
R1449 B.n741 B.n43 163.367
R1450 B.n741 B.n48 163.367
R1451 B.n49 B.n48 163.367
R1452 B.n50 B.n49 163.367
R1453 B.n746 B.n50 163.367
R1454 B.n746 B.n55 163.367
R1455 B.n56 B.n55 163.367
R1456 B.n57 B.n56 163.367
R1457 B.n751 B.n57 163.367
R1458 B.n751 B.n62 163.367
R1459 B.n63 B.n62 163.367
R1460 B.n64 B.n63 163.367
R1461 B.n756 B.n64 163.367
R1462 B.n756 B.n69 163.367
R1463 B.n70 B.n69 163.367
R1464 B.n71 B.n70 163.367
R1465 B.n761 B.n71 163.367
R1466 B.n761 B.n76 163.367
R1467 B.n419 B.n418 163.367
R1468 B.n421 B.n419 163.367
R1469 B.n425 B.n414 163.367
R1470 B.n429 B.n427 163.367
R1471 B.n433 B.n412 163.367
R1472 B.n437 B.n435 163.367
R1473 B.n441 B.n410 163.367
R1474 B.n445 B.n443 163.367
R1475 B.n449 B.n408 163.367
R1476 B.n453 B.n451 163.367
R1477 B.n457 B.n406 163.367
R1478 B.n461 B.n459 163.367
R1479 B.n465 B.n404 163.367
R1480 B.n469 B.n467 163.367
R1481 B.n473 B.n402 163.367
R1482 B.n477 B.n475 163.367
R1483 B.n481 B.n400 163.367
R1484 B.n485 B.n483 163.367
R1485 B.n492 B.n398 163.367
R1486 B.n496 B.n494 163.367
R1487 B.n500 B.n396 163.367
R1488 B.n504 B.n502 163.367
R1489 B.n508 B.n394 163.367
R1490 B.n512 B.n510 163.367
R1491 B.n517 B.n390 163.367
R1492 B.n521 B.n519 163.367
R1493 B.n525 B.n388 163.367
R1494 B.n529 B.n527 163.367
R1495 B.n533 B.n386 163.367
R1496 B.n537 B.n535 163.367
R1497 B.n541 B.n384 163.367
R1498 B.n545 B.n543 163.367
R1499 B.n549 B.n382 163.367
R1500 B.n553 B.n551 163.367
R1501 B.n557 B.n380 163.367
R1502 B.n561 B.n559 163.367
R1503 B.n565 B.n378 163.367
R1504 B.n569 B.n567 163.367
R1505 B.n573 B.n376 163.367
R1506 B.n577 B.n575 163.367
R1507 B.n581 B.n374 163.367
R1508 B.n584 B.n583 163.367
R1509 B.n586 B.n371 163.367
R1510 B.n592 B.n367 163.367
R1511 B.n596 B.n367 163.367
R1512 B.n596 B.n361 163.367
R1513 B.n604 B.n361 163.367
R1514 B.n604 B.n359 163.367
R1515 B.n608 B.n359 163.367
R1516 B.n608 B.n353 163.367
R1517 B.n616 B.n353 163.367
R1518 B.n616 B.n351 163.367
R1519 B.n620 B.n351 163.367
R1520 B.n620 B.n345 163.367
R1521 B.n628 B.n345 163.367
R1522 B.n628 B.n343 163.367
R1523 B.n632 B.n343 163.367
R1524 B.n632 B.n337 163.367
R1525 B.n640 B.n337 163.367
R1526 B.n640 B.n335 163.367
R1527 B.n644 B.n335 163.367
R1528 B.n644 B.n329 163.367
R1529 B.n652 B.n329 163.367
R1530 B.n652 B.n327 163.367
R1531 B.n656 B.n327 163.367
R1532 B.n656 B.n321 163.367
R1533 B.n664 B.n321 163.367
R1534 B.n664 B.n319 163.367
R1535 B.n668 B.n319 163.367
R1536 B.n668 B.n313 163.367
R1537 B.n676 B.n313 163.367
R1538 B.n676 B.n311 163.367
R1539 B.n680 B.n311 163.367
R1540 B.n680 B.n305 163.367
R1541 B.n689 B.n305 163.367
R1542 B.n689 B.n303 163.367
R1543 B.n693 B.n303 163.367
R1544 B.n693 B.n298 163.367
R1545 B.n702 B.n298 163.367
R1546 B.n702 B.n296 163.367
R1547 B.n706 B.n296 163.367
R1548 B.n706 B.n3 163.367
R1549 B.n850 B.n3 163.367
R1550 B.n846 B.n2 163.367
R1551 B.n846 B.n845 163.367
R1552 B.n845 B.n9 163.367
R1553 B.n841 B.n9 163.367
R1554 B.n841 B.n11 163.367
R1555 B.n837 B.n11 163.367
R1556 B.n837 B.n16 163.367
R1557 B.n833 B.n16 163.367
R1558 B.n833 B.n18 163.367
R1559 B.n829 B.n18 163.367
R1560 B.n829 B.n24 163.367
R1561 B.n825 B.n24 163.367
R1562 B.n825 B.n26 163.367
R1563 B.n821 B.n26 163.367
R1564 B.n821 B.n31 163.367
R1565 B.n817 B.n31 163.367
R1566 B.n817 B.n33 163.367
R1567 B.n813 B.n33 163.367
R1568 B.n813 B.n38 163.367
R1569 B.n809 B.n38 163.367
R1570 B.n809 B.n40 163.367
R1571 B.n805 B.n40 163.367
R1572 B.n805 B.n45 163.367
R1573 B.n801 B.n45 163.367
R1574 B.n801 B.n47 163.367
R1575 B.n797 B.n47 163.367
R1576 B.n797 B.n52 163.367
R1577 B.n793 B.n52 163.367
R1578 B.n793 B.n54 163.367
R1579 B.n789 B.n54 163.367
R1580 B.n789 B.n59 163.367
R1581 B.n785 B.n59 163.367
R1582 B.n785 B.n61 163.367
R1583 B.n781 B.n61 163.367
R1584 B.n781 B.n66 163.367
R1585 B.n777 B.n66 163.367
R1586 B.n777 B.n68 163.367
R1587 B.n773 B.n68 163.367
R1588 B.n773 B.n73 163.367
R1589 B.n769 B.n73 163.367
R1590 B.n591 B.n370 96.0674
R1591 B.n768 B.n767 96.0674
R1592 B.n124 B.n123 71.7581
R1593 B.n121 B.n120 71.7581
R1594 B.n392 B.n391 71.7581
R1595 B.n489 B.n488 71.7581
R1596 B.n77 B.n75 71.676
R1597 B.n128 B.n78 71.676
R1598 B.n132 B.n79 71.676
R1599 B.n136 B.n80 71.676
R1600 B.n140 B.n81 71.676
R1601 B.n144 B.n82 71.676
R1602 B.n148 B.n83 71.676
R1603 B.n152 B.n84 71.676
R1604 B.n156 B.n85 71.676
R1605 B.n160 B.n86 71.676
R1606 B.n164 B.n87 71.676
R1607 B.n168 B.n88 71.676
R1608 B.n172 B.n89 71.676
R1609 B.n176 B.n90 71.676
R1610 B.n180 B.n91 71.676
R1611 B.n184 B.n92 71.676
R1612 B.n188 B.n93 71.676
R1613 B.n192 B.n94 71.676
R1614 B.n196 B.n95 71.676
R1615 B.n200 B.n96 71.676
R1616 B.n204 B.n97 71.676
R1617 B.n208 B.n98 71.676
R1618 B.n212 B.n99 71.676
R1619 B.n216 B.n100 71.676
R1620 B.n220 B.n101 71.676
R1621 B.n224 B.n102 71.676
R1622 B.n228 B.n103 71.676
R1623 B.n232 B.n104 71.676
R1624 B.n236 B.n105 71.676
R1625 B.n240 B.n106 71.676
R1626 B.n244 B.n107 71.676
R1627 B.n248 B.n108 71.676
R1628 B.n252 B.n109 71.676
R1629 B.n256 B.n110 71.676
R1630 B.n260 B.n111 71.676
R1631 B.n264 B.n112 71.676
R1632 B.n268 B.n113 71.676
R1633 B.n272 B.n114 71.676
R1634 B.n276 B.n115 71.676
R1635 B.n280 B.n116 71.676
R1636 B.n284 B.n117 71.676
R1637 B.n288 B.n118 71.676
R1638 B.n766 B.n119 71.676
R1639 B.n766 B.n765 71.676
R1640 B.n290 B.n118 71.676
R1641 B.n287 B.n117 71.676
R1642 B.n283 B.n116 71.676
R1643 B.n279 B.n115 71.676
R1644 B.n275 B.n114 71.676
R1645 B.n271 B.n113 71.676
R1646 B.n267 B.n112 71.676
R1647 B.n263 B.n111 71.676
R1648 B.n259 B.n110 71.676
R1649 B.n255 B.n109 71.676
R1650 B.n251 B.n108 71.676
R1651 B.n247 B.n107 71.676
R1652 B.n243 B.n106 71.676
R1653 B.n239 B.n105 71.676
R1654 B.n235 B.n104 71.676
R1655 B.n231 B.n103 71.676
R1656 B.n227 B.n102 71.676
R1657 B.n223 B.n101 71.676
R1658 B.n219 B.n100 71.676
R1659 B.n215 B.n99 71.676
R1660 B.n211 B.n98 71.676
R1661 B.n207 B.n97 71.676
R1662 B.n203 B.n96 71.676
R1663 B.n199 B.n95 71.676
R1664 B.n195 B.n94 71.676
R1665 B.n191 B.n93 71.676
R1666 B.n187 B.n92 71.676
R1667 B.n183 B.n91 71.676
R1668 B.n179 B.n90 71.676
R1669 B.n175 B.n89 71.676
R1670 B.n171 B.n88 71.676
R1671 B.n167 B.n87 71.676
R1672 B.n163 B.n86 71.676
R1673 B.n159 B.n85 71.676
R1674 B.n155 B.n84 71.676
R1675 B.n151 B.n83 71.676
R1676 B.n147 B.n82 71.676
R1677 B.n143 B.n81 71.676
R1678 B.n139 B.n80 71.676
R1679 B.n135 B.n79 71.676
R1680 B.n131 B.n78 71.676
R1681 B.n127 B.n77 71.676
R1682 B.n417 B.n369 71.676
R1683 B.n421 B.n420 71.676
R1684 B.n426 B.n425 71.676
R1685 B.n429 B.n428 71.676
R1686 B.n434 B.n433 71.676
R1687 B.n437 B.n436 71.676
R1688 B.n442 B.n441 71.676
R1689 B.n445 B.n444 71.676
R1690 B.n450 B.n449 71.676
R1691 B.n453 B.n452 71.676
R1692 B.n458 B.n457 71.676
R1693 B.n461 B.n460 71.676
R1694 B.n466 B.n465 71.676
R1695 B.n469 B.n468 71.676
R1696 B.n474 B.n473 71.676
R1697 B.n477 B.n476 71.676
R1698 B.n482 B.n481 71.676
R1699 B.n485 B.n484 71.676
R1700 B.n493 B.n492 71.676
R1701 B.n496 B.n495 71.676
R1702 B.n501 B.n500 71.676
R1703 B.n504 B.n503 71.676
R1704 B.n509 B.n508 71.676
R1705 B.n512 B.n511 71.676
R1706 B.n518 B.n517 71.676
R1707 B.n521 B.n520 71.676
R1708 B.n526 B.n525 71.676
R1709 B.n529 B.n528 71.676
R1710 B.n534 B.n533 71.676
R1711 B.n537 B.n536 71.676
R1712 B.n542 B.n541 71.676
R1713 B.n545 B.n544 71.676
R1714 B.n550 B.n549 71.676
R1715 B.n553 B.n552 71.676
R1716 B.n558 B.n557 71.676
R1717 B.n561 B.n560 71.676
R1718 B.n566 B.n565 71.676
R1719 B.n569 B.n568 71.676
R1720 B.n574 B.n573 71.676
R1721 B.n577 B.n576 71.676
R1722 B.n582 B.n581 71.676
R1723 B.n585 B.n584 71.676
R1724 B.n418 B.n417 71.676
R1725 B.n420 B.n414 71.676
R1726 B.n427 B.n426 71.676
R1727 B.n428 B.n412 71.676
R1728 B.n435 B.n434 71.676
R1729 B.n436 B.n410 71.676
R1730 B.n443 B.n442 71.676
R1731 B.n444 B.n408 71.676
R1732 B.n451 B.n450 71.676
R1733 B.n452 B.n406 71.676
R1734 B.n459 B.n458 71.676
R1735 B.n460 B.n404 71.676
R1736 B.n467 B.n466 71.676
R1737 B.n468 B.n402 71.676
R1738 B.n475 B.n474 71.676
R1739 B.n476 B.n400 71.676
R1740 B.n483 B.n482 71.676
R1741 B.n484 B.n398 71.676
R1742 B.n494 B.n493 71.676
R1743 B.n495 B.n396 71.676
R1744 B.n502 B.n501 71.676
R1745 B.n503 B.n394 71.676
R1746 B.n510 B.n509 71.676
R1747 B.n511 B.n390 71.676
R1748 B.n519 B.n518 71.676
R1749 B.n520 B.n388 71.676
R1750 B.n527 B.n526 71.676
R1751 B.n528 B.n386 71.676
R1752 B.n535 B.n534 71.676
R1753 B.n536 B.n384 71.676
R1754 B.n543 B.n542 71.676
R1755 B.n544 B.n382 71.676
R1756 B.n551 B.n550 71.676
R1757 B.n552 B.n380 71.676
R1758 B.n559 B.n558 71.676
R1759 B.n560 B.n378 71.676
R1760 B.n567 B.n566 71.676
R1761 B.n568 B.n376 71.676
R1762 B.n575 B.n574 71.676
R1763 B.n576 B.n374 71.676
R1764 B.n583 B.n582 71.676
R1765 B.n586 B.n585 71.676
R1766 B.n851 B.n850 71.676
R1767 B.n851 B.n2 71.676
R1768 B.n125 B.n124 59.5399
R1769 B.n122 B.n121 59.5399
R1770 B.n514 B.n392 59.5399
R1771 B.n490 B.n489 59.5399
R1772 B.n591 B.n366 46.3306
R1773 B.n597 B.n366 46.3306
R1774 B.n597 B.n362 46.3306
R1775 B.n603 B.n362 46.3306
R1776 B.n603 B.n358 46.3306
R1777 B.n609 B.n358 46.3306
R1778 B.n609 B.n354 46.3306
R1779 B.n615 B.n354 46.3306
R1780 B.n621 B.n350 46.3306
R1781 B.n621 B.n346 46.3306
R1782 B.n627 B.n346 46.3306
R1783 B.n627 B.n342 46.3306
R1784 B.n633 B.n342 46.3306
R1785 B.n633 B.n338 46.3306
R1786 B.n639 B.n338 46.3306
R1787 B.n639 B.n334 46.3306
R1788 B.n645 B.n334 46.3306
R1789 B.n645 B.n330 46.3306
R1790 B.n651 B.n330 46.3306
R1791 B.n651 B.n326 46.3306
R1792 B.n657 B.n326 46.3306
R1793 B.n663 B.n322 46.3306
R1794 B.n663 B.n318 46.3306
R1795 B.n669 B.n318 46.3306
R1796 B.n669 B.n314 46.3306
R1797 B.n675 B.n314 46.3306
R1798 B.n675 B.n310 46.3306
R1799 B.n681 B.n310 46.3306
R1800 B.n681 B.n306 46.3306
R1801 B.n688 B.n306 46.3306
R1802 B.n688 B.n687 46.3306
R1803 B.n694 B.n299 46.3306
R1804 B.n701 B.n299 46.3306
R1805 B.n701 B.n295 46.3306
R1806 B.n707 B.n295 46.3306
R1807 B.n707 B.n4 46.3306
R1808 B.n849 B.n4 46.3306
R1809 B.n849 B.n848 46.3306
R1810 B.n848 B.n847 46.3306
R1811 B.n847 B.n8 46.3306
R1812 B.n12 B.n8 46.3306
R1813 B.n840 B.n12 46.3306
R1814 B.n840 B.n839 46.3306
R1815 B.n839 B.n838 46.3306
R1816 B.n832 B.n19 46.3306
R1817 B.n832 B.n831 46.3306
R1818 B.n831 B.n830 46.3306
R1819 B.n830 B.n23 46.3306
R1820 B.n824 B.n23 46.3306
R1821 B.n824 B.n823 46.3306
R1822 B.n823 B.n822 46.3306
R1823 B.n822 B.n30 46.3306
R1824 B.n816 B.n30 46.3306
R1825 B.n816 B.n815 46.3306
R1826 B.n814 B.n37 46.3306
R1827 B.n808 B.n37 46.3306
R1828 B.n808 B.n807 46.3306
R1829 B.n807 B.n806 46.3306
R1830 B.n806 B.n44 46.3306
R1831 B.n800 B.n44 46.3306
R1832 B.n800 B.n799 46.3306
R1833 B.n799 B.n798 46.3306
R1834 B.n798 B.n51 46.3306
R1835 B.n792 B.n51 46.3306
R1836 B.n792 B.n791 46.3306
R1837 B.n791 B.n790 46.3306
R1838 B.n790 B.n58 46.3306
R1839 B.n784 B.n783 46.3306
R1840 B.n783 B.n782 46.3306
R1841 B.n782 B.n65 46.3306
R1842 B.n776 B.n65 46.3306
R1843 B.n776 B.n775 46.3306
R1844 B.n775 B.n774 46.3306
R1845 B.n774 B.n72 46.3306
R1846 B.n768 B.n72 46.3306
R1847 B.n764 B.n763 36.059
R1848 B.n593 B.n368 36.059
R1849 B.n589 B.n588 36.059
R1850 B.n770 B.n74 36.059
R1851 B.n657 B.t2 26.5722
R1852 B.t1 B.n814 26.5722
R1853 B.n694 B.t3 25.2095
R1854 B.n838 B.t0 25.2095
R1855 B.t5 B.n350 23.8469
R1856 B.t12 B.n58 23.8469
R1857 B.n615 B.t5 22.4842
R1858 B.n784 B.t12 22.4842
R1859 B.n687 B.t3 21.1216
R1860 B.n19 B.t0 21.1216
R1861 B.t2 B.n322 19.7589
R1862 B.n815 B.t1 19.7589
R1863 B B.n852 18.0485
R1864 B.n594 B.n593 10.6151
R1865 B.n595 B.n594 10.6151
R1866 B.n595 B.n360 10.6151
R1867 B.n605 B.n360 10.6151
R1868 B.n606 B.n605 10.6151
R1869 B.n607 B.n606 10.6151
R1870 B.n607 B.n352 10.6151
R1871 B.n617 B.n352 10.6151
R1872 B.n618 B.n617 10.6151
R1873 B.n619 B.n618 10.6151
R1874 B.n619 B.n344 10.6151
R1875 B.n629 B.n344 10.6151
R1876 B.n630 B.n629 10.6151
R1877 B.n631 B.n630 10.6151
R1878 B.n631 B.n336 10.6151
R1879 B.n641 B.n336 10.6151
R1880 B.n642 B.n641 10.6151
R1881 B.n643 B.n642 10.6151
R1882 B.n643 B.n328 10.6151
R1883 B.n653 B.n328 10.6151
R1884 B.n654 B.n653 10.6151
R1885 B.n655 B.n654 10.6151
R1886 B.n655 B.n320 10.6151
R1887 B.n665 B.n320 10.6151
R1888 B.n666 B.n665 10.6151
R1889 B.n667 B.n666 10.6151
R1890 B.n667 B.n312 10.6151
R1891 B.n677 B.n312 10.6151
R1892 B.n678 B.n677 10.6151
R1893 B.n679 B.n678 10.6151
R1894 B.n679 B.n304 10.6151
R1895 B.n690 B.n304 10.6151
R1896 B.n691 B.n690 10.6151
R1897 B.n692 B.n691 10.6151
R1898 B.n692 B.n297 10.6151
R1899 B.n703 B.n297 10.6151
R1900 B.n704 B.n703 10.6151
R1901 B.n705 B.n704 10.6151
R1902 B.n705 B.n0 10.6151
R1903 B.n416 B.n368 10.6151
R1904 B.n416 B.n415 10.6151
R1905 B.n422 B.n415 10.6151
R1906 B.n423 B.n422 10.6151
R1907 B.n424 B.n423 10.6151
R1908 B.n424 B.n413 10.6151
R1909 B.n430 B.n413 10.6151
R1910 B.n431 B.n430 10.6151
R1911 B.n432 B.n431 10.6151
R1912 B.n432 B.n411 10.6151
R1913 B.n438 B.n411 10.6151
R1914 B.n439 B.n438 10.6151
R1915 B.n440 B.n439 10.6151
R1916 B.n440 B.n409 10.6151
R1917 B.n446 B.n409 10.6151
R1918 B.n447 B.n446 10.6151
R1919 B.n448 B.n447 10.6151
R1920 B.n448 B.n407 10.6151
R1921 B.n454 B.n407 10.6151
R1922 B.n455 B.n454 10.6151
R1923 B.n456 B.n455 10.6151
R1924 B.n456 B.n405 10.6151
R1925 B.n462 B.n405 10.6151
R1926 B.n463 B.n462 10.6151
R1927 B.n464 B.n463 10.6151
R1928 B.n464 B.n403 10.6151
R1929 B.n470 B.n403 10.6151
R1930 B.n471 B.n470 10.6151
R1931 B.n472 B.n471 10.6151
R1932 B.n472 B.n401 10.6151
R1933 B.n478 B.n401 10.6151
R1934 B.n479 B.n478 10.6151
R1935 B.n480 B.n479 10.6151
R1936 B.n480 B.n399 10.6151
R1937 B.n486 B.n399 10.6151
R1938 B.n487 B.n486 10.6151
R1939 B.n491 B.n487 10.6151
R1940 B.n497 B.n397 10.6151
R1941 B.n498 B.n497 10.6151
R1942 B.n499 B.n498 10.6151
R1943 B.n499 B.n395 10.6151
R1944 B.n505 B.n395 10.6151
R1945 B.n506 B.n505 10.6151
R1946 B.n507 B.n506 10.6151
R1947 B.n507 B.n393 10.6151
R1948 B.n513 B.n393 10.6151
R1949 B.n516 B.n515 10.6151
R1950 B.n516 B.n389 10.6151
R1951 B.n522 B.n389 10.6151
R1952 B.n523 B.n522 10.6151
R1953 B.n524 B.n523 10.6151
R1954 B.n524 B.n387 10.6151
R1955 B.n530 B.n387 10.6151
R1956 B.n531 B.n530 10.6151
R1957 B.n532 B.n531 10.6151
R1958 B.n532 B.n385 10.6151
R1959 B.n538 B.n385 10.6151
R1960 B.n539 B.n538 10.6151
R1961 B.n540 B.n539 10.6151
R1962 B.n540 B.n383 10.6151
R1963 B.n546 B.n383 10.6151
R1964 B.n547 B.n546 10.6151
R1965 B.n548 B.n547 10.6151
R1966 B.n548 B.n381 10.6151
R1967 B.n554 B.n381 10.6151
R1968 B.n555 B.n554 10.6151
R1969 B.n556 B.n555 10.6151
R1970 B.n556 B.n379 10.6151
R1971 B.n562 B.n379 10.6151
R1972 B.n563 B.n562 10.6151
R1973 B.n564 B.n563 10.6151
R1974 B.n564 B.n377 10.6151
R1975 B.n570 B.n377 10.6151
R1976 B.n571 B.n570 10.6151
R1977 B.n572 B.n571 10.6151
R1978 B.n572 B.n375 10.6151
R1979 B.n578 B.n375 10.6151
R1980 B.n579 B.n578 10.6151
R1981 B.n580 B.n579 10.6151
R1982 B.n580 B.n373 10.6151
R1983 B.n373 B.n372 10.6151
R1984 B.n587 B.n372 10.6151
R1985 B.n588 B.n587 10.6151
R1986 B.n589 B.n364 10.6151
R1987 B.n599 B.n364 10.6151
R1988 B.n600 B.n599 10.6151
R1989 B.n601 B.n600 10.6151
R1990 B.n601 B.n356 10.6151
R1991 B.n611 B.n356 10.6151
R1992 B.n612 B.n611 10.6151
R1993 B.n613 B.n612 10.6151
R1994 B.n613 B.n348 10.6151
R1995 B.n623 B.n348 10.6151
R1996 B.n624 B.n623 10.6151
R1997 B.n625 B.n624 10.6151
R1998 B.n625 B.n340 10.6151
R1999 B.n635 B.n340 10.6151
R2000 B.n636 B.n635 10.6151
R2001 B.n637 B.n636 10.6151
R2002 B.n637 B.n332 10.6151
R2003 B.n647 B.n332 10.6151
R2004 B.n648 B.n647 10.6151
R2005 B.n649 B.n648 10.6151
R2006 B.n649 B.n324 10.6151
R2007 B.n659 B.n324 10.6151
R2008 B.n660 B.n659 10.6151
R2009 B.n661 B.n660 10.6151
R2010 B.n661 B.n316 10.6151
R2011 B.n671 B.n316 10.6151
R2012 B.n672 B.n671 10.6151
R2013 B.n673 B.n672 10.6151
R2014 B.n673 B.n308 10.6151
R2015 B.n683 B.n308 10.6151
R2016 B.n684 B.n683 10.6151
R2017 B.n685 B.n684 10.6151
R2018 B.n685 B.n301 10.6151
R2019 B.n696 B.n301 10.6151
R2020 B.n697 B.n696 10.6151
R2021 B.n699 B.n697 10.6151
R2022 B.n699 B.n698 10.6151
R2023 B.n698 B.n293 10.6151
R2024 B.n710 B.n293 10.6151
R2025 B.n711 B.n710 10.6151
R2026 B.n712 B.n711 10.6151
R2027 B.n713 B.n712 10.6151
R2028 B.n714 B.n713 10.6151
R2029 B.n717 B.n714 10.6151
R2030 B.n718 B.n717 10.6151
R2031 B.n719 B.n718 10.6151
R2032 B.n720 B.n719 10.6151
R2033 B.n722 B.n720 10.6151
R2034 B.n723 B.n722 10.6151
R2035 B.n724 B.n723 10.6151
R2036 B.n725 B.n724 10.6151
R2037 B.n727 B.n725 10.6151
R2038 B.n728 B.n727 10.6151
R2039 B.n729 B.n728 10.6151
R2040 B.n730 B.n729 10.6151
R2041 B.n732 B.n730 10.6151
R2042 B.n733 B.n732 10.6151
R2043 B.n734 B.n733 10.6151
R2044 B.n735 B.n734 10.6151
R2045 B.n737 B.n735 10.6151
R2046 B.n738 B.n737 10.6151
R2047 B.n739 B.n738 10.6151
R2048 B.n740 B.n739 10.6151
R2049 B.n742 B.n740 10.6151
R2050 B.n743 B.n742 10.6151
R2051 B.n744 B.n743 10.6151
R2052 B.n745 B.n744 10.6151
R2053 B.n747 B.n745 10.6151
R2054 B.n748 B.n747 10.6151
R2055 B.n749 B.n748 10.6151
R2056 B.n750 B.n749 10.6151
R2057 B.n752 B.n750 10.6151
R2058 B.n753 B.n752 10.6151
R2059 B.n754 B.n753 10.6151
R2060 B.n755 B.n754 10.6151
R2061 B.n757 B.n755 10.6151
R2062 B.n758 B.n757 10.6151
R2063 B.n759 B.n758 10.6151
R2064 B.n760 B.n759 10.6151
R2065 B.n762 B.n760 10.6151
R2066 B.n763 B.n762 10.6151
R2067 B.n844 B.n1 10.6151
R2068 B.n844 B.n843 10.6151
R2069 B.n843 B.n842 10.6151
R2070 B.n842 B.n10 10.6151
R2071 B.n836 B.n10 10.6151
R2072 B.n836 B.n835 10.6151
R2073 B.n835 B.n834 10.6151
R2074 B.n834 B.n17 10.6151
R2075 B.n828 B.n17 10.6151
R2076 B.n828 B.n827 10.6151
R2077 B.n827 B.n826 10.6151
R2078 B.n826 B.n25 10.6151
R2079 B.n820 B.n25 10.6151
R2080 B.n820 B.n819 10.6151
R2081 B.n819 B.n818 10.6151
R2082 B.n818 B.n32 10.6151
R2083 B.n812 B.n32 10.6151
R2084 B.n812 B.n811 10.6151
R2085 B.n811 B.n810 10.6151
R2086 B.n810 B.n39 10.6151
R2087 B.n804 B.n39 10.6151
R2088 B.n804 B.n803 10.6151
R2089 B.n803 B.n802 10.6151
R2090 B.n802 B.n46 10.6151
R2091 B.n796 B.n46 10.6151
R2092 B.n796 B.n795 10.6151
R2093 B.n795 B.n794 10.6151
R2094 B.n794 B.n53 10.6151
R2095 B.n788 B.n53 10.6151
R2096 B.n788 B.n787 10.6151
R2097 B.n787 B.n786 10.6151
R2098 B.n786 B.n60 10.6151
R2099 B.n780 B.n60 10.6151
R2100 B.n780 B.n779 10.6151
R2101 B.n779 B.n778 10.6151
R2102 B.n778 B.n67 10.6151
R2103 B.n772 B.n67 10.6151
R2104 B.n772 B.n771 10.6151
R2105 B.n771 B.n770 10.6151
R2106 B.n126 B.n74 10.6151
R2107 B.n129 B.n126 10.6151
R2108 B.n130 B.n129 10.6151
R2109 B.n133 B.n130 10.6151
R2110 B.n134 B.n133 10.6151
R2111 B.n137 B.n134 10.6151
R2112 B.n138 B.n137 10.6151
R2113 B.n141 B.n138 10.6151
R2114 B.n142 B.n141 10.6151
R2115 B.n145 B.n142 10.6151
R2116 B.n146 B.n145 10.6151
R2117 B.n149 B.n146 10.6151
R2118 B.n150 B.n149 10.6151
R2119 B.n153 B.n150 10.6151
R2120 B.n154 B.n153 10.6151
R2121 B.n157 B.n154 10.6151
R2122 B.n158 B.n157 10.6151
R2123 B.n161 B.n158 10.6151
R2124 B.n162 B.n161 10.6151
R2125 B.n165 B.n162 10.6151
R2126 B.n166 B.n165 10.6151
R2127 B.n169 B.n166 10.6151
R2128 B.n170 B.n169 10.6151
R2129 B.n173 B.n170 10.6151
R2130 B.n174 B.n173 10.6151
R2131 B.n177 B.n174 10.6151
R2132 B.n178 B.n177 10.6151
R2133 B.n181 B.n178 10.6151
R2134 B.n182 B.n181 10.6151
R2135 B.n185 B.n182 10.6151
R2136 B.n186 B.n185 10.6151
R2137 B.n189 B.n186 10.6151
R2138 B.n190 B.n189 10.6151
R2139 B.n193 B.n190 10.6151
R2140 B.n194 B.n193 10.6151
R2141 B.n197 B.n194 10.6151
R2142 B.n198 B.n197 10.6151
R2143 B.n202 B.n201 10.6151
R2144 B.n205 B.n202 10.6151
R2145 B.n206 B.n205 10.6151
R2146 B.n209 B.n206 10.6151
R2147 B.n210 B.n209 10.6151
R2148 B.n213 B.n210 10.6151
R2149 B.n214 B.n213 10.6151
R2150 B.n217 B.n214 10.6151
R2151 B.n218 B.n217 10.6151
R2152 B.n222 B.n221 10.6151
R2153 B.n225 B.n222 10.6151
R2154 B.n226 B.n225 10.6151
R2155 B.n229 B.n226 10.6151
R2156 B.n230 B.n229 10.6151
R2157 B.n233 B.n230 10.6151
R2158 B.n234 B.n233 10.6151
R2159 B.n237 B.n234 10.6151
R2160 B.n238 B.n237 10.6151
R2161 B.n241 B.n238 10.6151
R2162 B.n242 B.n241 10.6151
R2163 B.n245 B.n242 10.6151
R2164 B.n246 B.n245 10.6151
R2165 B.n249 B.n246 10.6151
R2166 B.n250 B.n249 10.6151
R2167 B.n253 B.n250 10.6151
R2168 B.n254 B.n253 10.6151
R2169 B.n257 B.n254 10.6151
R2170 B.n258 B.n257 10.6151
R2171 B.n261 B.n258 10.6151
R2172 B.n262 B.n261 10.6151
R2173 B.n265 B.n262 10.6151
R2174 B.n266 B.n265 10.6151
R2175 B.n269 B.n266 10.6151
R2176 B.n270 B.n269 10.6151
R2177 B.n273 B.n270 10.6151
R2178 B.n274 B.n273 10.6151
R2179 B.n277 B.n274 10.6151
R2180 B.n278 B.n277 10.6151
R2181 B.n281 B.n278 10.6151
R2182 B.n282 B.n281 10.6151
R2183 B.n285 B.n282 10.6151
R2184 B.n286 B.n285 10.6151
R2185 B.n289 B.n286 10.6151
R2186 B.n291 B.n289 10.6151
R2187 B.n292 B.n291 10.6151
R2188 B.n764 B.n292 10.6151
R2189 B.n491 B.n490 9.36635
R2190 B.n515 B.n514 9.36635
R2191 B.n198 B.n125 9.36635
R2192 B.n221 B.n122 9.36635
R2193 B.n852 B.n0 8.11757
R2194 B.n852 B.n1 8.11757
R2195 B.n490 B.n397 1.24928
R2196 B.n514 B.n513 1.24928
R2197 B.n201 B.n125 1.24928
R2198 B.n218 B.n122 1.24928
R2199 VN.n1 VN.t3 112.817
R2200 VN.n0 VN.t0 112.817
R2201 VN.n0 VN.t2 111.683
R2202 VN.n1 VN.t1 111.683
R2203 VN VN.n1 50.4961
R2204 VN VN.n0 2.39381
R2205 VDD2.n2 VDD2.n0 108.68
R2206 VDD2.n2 VDD2.n1 66.025
R2207 VDD2.n1 VDD2.t2 1.82203
R2208 VDD2.n1 VDD2.t0 1.82203
R2209 VDD2.n0 VDD2.t3 1.82203
R2210 VDD2.n0 VDD2.t1 1.82203
R2211 VDD2 VDD2.n2 0.0586897
C0 VN VDD1 0.149543f
C1 VDD1 VP 4.81271f
C2 VDD1 VTAIL 5.35311f
C3 VDD2 VN 4.52004f
C4 VDD2 VP 0.443149f
C5 VDD2 VTAIL 5.41248f
C6 VN VP 6.53462f
C7 VN VTAIL 4.5932f
C8 VTAIL VP 4.6073f
C9 VDD2 VDD1 1.20559f
C10 VDD2 B 4.122184f
C11 VDD1 B 8.48366f
C12 VTAIL B 9.817608f
C13 VN B 12.087449f
C14 VP B 10.500535f
C15 VDD2.t3 B 0.233399f
C16 VDD2.t1 B 0.233399f
C17 VDD2.n0 B 2.72376f
C18 VDD2.t2 B 0.233399f
C19 VDD2.t0 B 0.233399f
C20 VDD2.n1 B 2.0702f
C21 VDD2.n2 B 3.88733f
C22 VN.t2 B 2.45564f
C23 VN.t0 B 2.46462f
C24 VN.n0 B 1.47188f
C25 VN.t1 B 2.45564f
C26 VN.t3 B 2.46462f
C27 VN.n1 B 2.80524f
C28 VDD1.t0 B 0.238059f
C29 VDD1.t1 B 0.238059f
C30 VDD1.n0 B 2.11199f
C31 VDD1.t2 B 0.238059f
C32 VDD1.t3 B 0.238059f
C33 VDD1.n1 B 2.80479f
C34 VTAIL.n0 B 0.025618f
C35 VTAIL.n1 B 0.017312f
C36 VTAIL.n2 B 0.009303f
C37 VTAIL.n3 B 0.021988f
C38 VTAIL.n4 B 0.00985f
C39 VTAIL.n5 B 0.017312f
C40 VTAIL.n6 B 0.009303f
C41 VTAIL.n7 B 0.021988f
C42 VTAIL.n8 B 0.00985f
C43 VTAIL.n9 B 0.017312f
C44 VTAIL.n10 B 0.009303f
C45 VTAIL.n11 B 0.021988f
C46 VTAIL.n12 B 0.00985f
C47 VTAIL.n13 B 0.017312f
C48 VTAIL.n14 B 0.009303f
C49 VTAIL.n15 B 0.021988f
C50 VTAIL.n16 B 0.00985f
C51 VTAIL.n17 B 0.117309f
C52 VTAIL.t4 B 0.037032f
C53 VTAIL.n18 B 0.016491f
C54 VTAIL.n19 B 0.015544f
C55 VTAIL.n20 B 0.009303f
C56 VTAIL.n21 B 0.786349f
C57 VTAIL.n22 B 0.017312f
C58 VTAIL.n23 B 0.009303f
C59 VTAIL.n24 B 0.00985f
C60 VTAIL.n25 B 0.021988f
C61 VTAIL.n26 B 0.021988f
C62 VTAIL.n27 B 0.00985f
C63 VTAIL.n28 B 0.009303f
C64 VTAIL.n29 B 0.017312f
C65 VTAIL.n30 B 0.017312f
C66 VTAIL.n31 B 0.009303f
C67 VTAIL.n32 B 0.00985f
C68 VTAIL.n33 B 0.021988f
C69 VTAIL.n34 B 0.021988f
C70 VTAIL.n35 B 0.021988f
C71 VTAIL.n36 B 0.00985f
C72 VTAIL.n37 B 0.009303f
C73 VTAIL.n38 B 0.017312f
C74 VTAIL.n39 B 0.017312f
C75 VTAIL.n40 B 0.009303f
C76 VTAIL.n41 B 0.009576f
C77 VTAIL.n42 B 0.009576f
C78 VTAIL.n43 B 0.021988f
C79 VTAIL.n44 B 0.021988f
C80 VTAIL.n45 B 0.00985f
C81 VTAIL.n46 B 0.009303f
C82 VTAIL.n47 B 0.017312f
C83 VTAIL.n48 B 0.017312f
C84 VTAIL.n49 B 0.009303f
C85 VTAIL.n50 B 0.00985f
C86 VTAIL.n51 B 0.021988f
C87 VTAIL.n52 B 0.049873f
C88 VTAIL.n53 B 0.00985f
C89 VTAIL.n54 B 0.009303f
C90 VTAIL.n55 B 0.044509f
C91 VTAIL.n56 B 0.028271f
C92 VTAIL.n57 B 0.135748f
C93 VTAIL.n58 B 0.025618f
C94 VTAIL.n59 B 0.017312f
C95 VTAIL.n60 B 0.009303f
C96 VTAIL.n61 B 0.021988f
C97 VTAIL.n62 B 0.00985f
C98 VTAIL.n63 B 0.017312f
C99 VTAIL.n64 B 0.009303f
C100 VTAIL.n65 B 0.021988f
C101 VTAIL.n66 B 0.00985f
C102 VTAIL.n67 B 0.017312f
C103 VTAIL.n68 B 0.009303f
C104 VTAIL.n69 B 0.021988f
C105 VTAIL.n70 B 0.00985f
C106 VTAIL.n71 B 0.017312f
C107 VTAIL.n72 B 0.009303f
C108 VTAIL.n73 B 0.021988f
C109 VTAIL.n74 B 0.00985f
C110 VTAIL.n75 B 0.117309f
C111 VTAIL.t2 B 0.037032f
C112 VTAIL.n76 B 0.016491f
C113 VTAIL.n77 B 0.015544f
C114 VTAIL.n78 B 0.009303f
C115 VTAIL.n79 B 0.786349f
C116 VTAIL.n80 B 0.017312f
C117 VTAIL.n81 B 0.009303f
C118 VTAIL.n82 B 0.00985f
C119 VTAIL.n83 B 0.021988f
C120 VTAIL.n84 B 0.021988f
C121 VTAIL.n85 B 0.00985f
C122 VTAIL.n86 B 0.009303f
C123 VTAIL.n87 B 0.017312f
C124 VTAIL.n88 B 0.017312f
C125 VTAIL.n89 B 0.009303f
C126 VTAIL.n90 B 0.00985f
C127 VTAIL.n91 B 0.021988f
C128 VTAIL.n92 B 0.021988f
C129 VTAIL.n93 B 0.021988f
C130 VTAIL.n94 B 0.00985f
C131 VTAIL.n95 B 0.009303f
C132 VTAIL.n96 B 0.017312f
C133 VTAIL.n97 B 0.017312f
C134 VTAIL.n98 B 0.009303f
C135 VTAIL.n99 B 0.009576f
C136 VTAIL.n100 B 0.009576f
C137 VTAIL.n101 B 0.021988f
C138 VTAIL.n102 B 0.021988f
C139 VTAIL.n103 B 0.00985f
C140 VTAIL.n104 B 0.009303f
C141 VTAIL.n105 B 0.017312f
C142 VTAIL.n106 B 0.017312f
C143 VTAIL.n107 B 0.009303f
C144 VTAIL.n108 B 0.00985f
C145 VTAIL.n109 B 0.021988f
C146 VTAIL.n110 B 0.049873f
C147 VTAIL.n111 B 0.00985f
C148 VTAIL.n112 B 0.009303f
C149 VTAIL.n113 B 0.044509f
C150 VTAIL.n114 B 0.028271f
C151 VTAIL.n115 B 0.221466f
C152 VTAIL.n116 B 0.025618f
C153 VTAIL.n117 B 0.017312f
C154 VTAIL.n118 B 0.009303f
C155 VTAIL.n119 B 0.021988f
C156 VTAIL.n120 B 0.00985f
C157 VTAIL.n121 B 0.017312f
C158 VTAIL.n122 B 0.009303f
C159 VTAIL.n123 B 0.021988f
C160 VTAIL.n124 B 0.00985f
C161 VTAIL.n125 B 0.017312f
C162 VTAIL.n126 B 0.009303f
C163 VTAIL.n127 B 0.021988f
C164 VTAIL.n128 B 0.00985f
C165 VTAIL.n129 B 0.017312f
C166 VTAIL.n130 B 0.009303f
C167 VTAIL.n131 B 0.021988f
C168 VTAIL.n132 B 0.00985f
C169 VTAIL.n133 B 0.117309f
C170 VTAIL.t3 B 0.037032f
C171 VTAIL.n134 B 0.016491f
C172 VTAIL.n135 B 0.015544f
C173 VTAIL.n136 B 0.009303f
C174 VTAIL.n137 B 0.786349f
C175 VTAIL.n138 B 0.017312f
C176 VTAIL.n139 B 0.009303f
C177 VTAIL.n140 B 0.00985f
C178 VTAIL.n141 B 0.021988f
C179 VTAIL.n142 B 0.021988f
C180 VTAIL.n143 B 0.00985f
C181 VTAIL.n144 B 0.009303f
C182 VTAIL.n145 B 0.017312f
C183 VTAIL.n146 B 0.017312f
C184 VTAIL.n147 B 0.009303f
C185 VTAIL.n148 B 0.00985f
C186 VTAIL.n149 B 0.021988f
C187 VTAIL.n150 B 0.021988f
C188 VTAIL.n151 B 0.021988f
C189 VTAIL.n152 B 0.00985f
C190 VTAIL.n153 B 0.009303f
C191 VTAIL.n154 B 0.017312f
C192 VTAIL.n155 B 0.017312f
C193 VTAIL.n156 B 0.009303f
C194 VTAIL.n157 B 0.009576f
C195 VTAIL.n158 B 0.009576f
C196 VTAIL.n159 B 0.021988f
C197 VTAIL.n160 B 0.021988f
C198 VTAIL.n161 B 0.00985f
C199 VTAIL.n162 B 0.009303f
C200 VTAIL.n163 B 0.017312f
C201 VTAIL.n164 B 0.017312f
C202 VTAIL.n165 B 0.009303f
C203 VTAIL.n166 B 0.00985f
C204 VTAIL.n167 B 0.021988f
C205 VTAIL.n168 B 0.049873f
C206 VTAIL.n169 B 0.00985f
C207 VTAIL.n170 B 0.009303f
C208 VTAIL.n171 B 0.044509f
C209 VTAIL.n172 B 0.028271f
C210 VTAIL.n173 B 1.13108f
C211 VTAIL.n174 B 0.025618f
C212 VTAIL.n175 B 0.017312f
C213 VTAIL.n176 B 0.009303f
C214 VTAIL.n177 B 0.021988f
C215 VTAIL.n178 B 0.00985f
C216 VTAIL.n179 B 0.017312f
C217 VTAIL.n180 B 0.009303f
C218 VTAIL.n181 B 0.021988f
C219 VTAIL.n182 B 0.00985f
C220 VTAIL.n183 B 0.017312f
C221 VTAIL.n184 B 0.009303f
C222 VTAIL.n185 B 0.021988f
C223 VTAIL.n186 B 0.021988f
C224 VTAIL.n187 B 0.00985f
C225 VTAIL.n188 B 0.017312f
C226 VTAIL.n189 B 0.009303f
C227 VTAIL.n190 B 0.021988f
C228 VTAIL.n191 B 0.00985f
C229 VTAIL.n192 B 0.117309f
C230 VTAIL.t7 B 0.037032f
C231 VTAIL.n193 B 0.016491f
C232 VTAIL.n194 B 0.015544f
C233 VTAIL.n195 B 0.009303f
C234 VTAIL.n196 B 0.786349f
C235 VTAIL.n197 B 0.017312f
C236 VTAIL.n198 B 0.009303f
C237 VTAIL.n199 B 0.00985f
C238 VTAIL.n200 B 0.021988f
C239 VTAIL.n201 B 0.021988f
C240 VTAIL.n202 B 0.00985f
C241 VTAIL.n203 B 0.009303f
C242 VTAIL.n204 B 0.017312f
C243 VTAIL.n205 B 0.017312f
C244 VTAIL.n206 B 0.009303f
C245 VTAIL.n207 B 0.00985f
C246 VTAIL.n208 B 0.021988f
C247 VTAIL.n209 B 0.021988f
C248 VTAIL.n210 B 0.00985f
C249 VTAIL.n211 B 0.009303f
C250 VTAIL.n212 B 0.017312f
C251 VTAIL.n213 B 0.017312f
C252 VTAIL.n214 B 0.009303f
C253 VTAIL.n215 B 0.009576f
C254 VTAIL.n216 B 0.009576f
C255 VTAIL.n217 B 0.021988f
C256 VTAIL.n218 B 0.021988f
C257 VTAIL.n219 B 0.00985f
C258 VTAIL.n220 B 0.009303f
C259 VTAIL.n221 B 0.017312f
C260 VTAIL.n222 B 0.017312f
C261 VTAIL.n223 B 0.009303f
C262 VTAIL.n224 B 0.00985f
C263 VTAIL.n225 B 0.021988f
C264 VTAIL.n226 B 0.049873f
C265 VTAIL.n227 B 0.00985f
C266 VTAIL.n228 B 0.009303f
C267 VTAIL.n229 B 0.044509f
C268 VTAIL.n230 B 0.028271f
C269 VTAIL.n231 B 1.13108f
C270 VTAIL.n232 B 0.025618f
C271 VTAIL.n233 B 0.017312f
C272 VTAIL.n234 B 0.009303f
C273 VTAIL.n235 B 0.021988f
C274 VTAIL.n236 B 0.00985f
C275 VTAIL.n237 B 0.017312f
C276 VTAIL.n238 B 0.009303f
C277 VTAIL.n239 B 0.021988f
C278 VTAIL.n240 B 0.00985f
C279 VTAIL.n241 B 0.017312f
C280 VTAIL.n242 B 0.009303f
C281 VTAIL.n243 B 0.021988f
C282 VTAIL.n244 B 0.021988f
C283 VTAIL.n245 B 0.00985f
C284 VTAIL.n246 B 0.017312f
C285 VTAIL.n247 B 0.009303f
C286 VTAIL.n248 B 0.021988f
C287 VTAIL.n249 B 0.00985f
C288 VTAIL.n250 B 0.117309f
C289 VTAIL.t5 B 0.037032f
C290 VTAIL.n251 B 0.016491f
C291 VTAIL.n252 B 0.015544f
C292 VTAIL.n253 B 0.009303f
C293 VTAIL.n254 B 0.786349f
C294 VTAIL.n255 B 0.017312f
C295 VTAIL.n256 B 0.009303f
C296 VTAIL.n257 B 0.00985f
C297 VTAIL.n258 B 0.021988f
C298 VTAIL.n259 B 0.021988f
C299 VTAIL.n260 B 0.00985f
C300 VTAIL.n261 B 0.009303f
C301 VTAIL.n262 B 0.017312f
C302 VTAIL.n263 B 0.017312f
C303 VTAIL.n264 B 0.009303f
C304 VTAIL.n265 B 0.00985f
C305 VTAIL.n266 B 0.021988f
C306 VTAIL.n267 B 0.021988f
C307 VTAIL.n268 B 0.00985f
C308 VTAIL.n269 B 0.009303f
C309 VTAIL.n270 B 0.017312f
C310 VTAIL.n271 B 0.017312f
C311 VTAIL.n272 B 0.009303f
C312 VTAIL.n273 B 0.009576f
C313 VTAIL.n274 B 0.009576f
C314 VTAIL.n275 B 0.021988f
C315 VTAIL.n276 B 0.021988f
C316 VTAIL.n277 B 0.00985f
C317 VTAIL.n278 B 0.009303f
C318 VTAIL.n279 B 0.017312f
C319 VTAIL.n280 B 0.017312f
C320 VTAIL.n281 B 0.009303f
C321 VTAIL.n282 B 0.00985f
C322 VTAIL.n283 B 0.021988f
C323 VTAIL.n284 B 0.049873f
C324 VTAIL.n285 B 0.00985f
C325 VTAIL.n286 B 0.009303f
C326 VTAIL.n287 B 0.044509f
C327 VTAIL.n288 B 0.028271f
C328 VTAIL.n289 B 0.221466f
C329 VTAIL.n290 B 0.025618f
C330 VTAIL.n291 B 0.017312f
C331 VTAIL.n292 B 0.009303f
C332 VTAIL.n293 B 0.021988f
C333 VTAIL.n294 B 0.00985f
C334 VTAIL.n295 B 0.017312f
C335 VTAIL.n296 B 0.009303f
C336 VTAIL.n297 B 0.021988f
C337 VTAIL.n298 B 0.00985f
C338 VTAIL.n299 B 0.017312f
C339 VTAIL.n300 B 0.009303f
C340 VTAIL.n301 B 0.021988f
C341 VTAIL.n302 B 0.021988f
C342 VTAIL.n303 B 0.00985f
C343 VTAIL.n304 B 0.017312f
C344 VTAIL.n305 B 0.009303f
C345 VTAIL.n306 B 0.021988f
C346 VTAIL.n307 B 0.00985f
C347 VTAIL.n308 B 0.117309f
C348 VTAIL.t0 B 0.037032f
C349 VTAIL.n309 B 0.016491f
C350 VTAIL.n310 B 0.015544f
C351 VTAIL.n311 B 0.009303f
C352 VTAIL.n312 B 0.786349f
C353 VTAIL.n313 B 0.017312f
C354 VTAIL.n314 B 0.009303f
C355 VTAIL.n315 B 0.00985f
C356 VTAIL.n316 B 0.021988f
C357 VTAIL.n317 B 0.021988f
C358 VTAIL.n318 B 0.00985f
C359 VTAIL.n319 B 0.009303f
C360 VTAIL.n320 B 0.017312f
C361 VTAIL.n321 B 0.017312f
C362 VTAIL.n322 B 0.009303f
C363 VTAIL.n323 B 0.00985f
C364 VTAIL.n324 B 0.021988f
C365 VTAIL.n325 B 0.021988f
C366 VTAIL.n326 B 0.00985f
C367 VTAIL.n327 B 0.009303f
C368 VTAIL.n328 B 0.017312f
C369 VTAIL.n329 B 0.017312f
C370 VTAIL.n330 B 0.009303f
C371 VTAIL.n331 B 0.009576f
C372 VTAIL.n332 B 0.009576f
C373 VTAIL.n333 B 0.021988f
C374 VTAIL.n334 B 0.021988f
C375 VTAIL.n335 B 0.00985f
C376 VTAIL.n336 B 0.009303f
C377 VTAIL.n337 B 0.017312f
C378 VTAIL.n338 B 0.017312f
C379 VTAIL.n339 B 0.009303f
C380 VTAIL.n340 B 0.00985f
C381 VTAIL.n341 B 0.021988f
C382 VTAIL.n342 B 0.049873f
C383 VTAIL.n343 B 0.00985f
C384 VTAIL.n344 B 0.009303f
C385 VTAIL.n345 B 0.044509f
C386 VTAIL.n346 B 0.028271f
C387 VTAIL.n347 B 0.221466f
C388 VTAIL.n348 B 0.025618f
C389 VTAIL.n349 B 0.017312f
C390 VTAIL.n350 B 0.009303f
C391 VTAIL.n351 B 0.021988f
C392 VTAIL.n352 B 0.00985f
C393 VTAIL.n353 B 0.017312f
C394 VTAIL.n354 B 0.009303f
C395 VTAIL.n355 B 0.021988f
C396 VTAIL.n356 B 0.00985f
C397 VTAIL.n357 B 0.017312f
C398 VTAIL.n358 B 0.009303f
C399 VTAIL.n359 B 0.021988f
C400 VTAIL.n360 B 0.021988f
C401 VTAIL.n361 B 0.00985f
C402 VTAIL.n362 B 0.017312f
C403 VTAIL.n363 B 0.009303f
C404 VTAIL.n364 B 0.021988f
C405 VTAIL.n365 B 0.00985f
C406 VTAIL.n366 B 0.117309f
C407 VTAIL.t1 B 0.037032f
C408 VTAIL.n367 B 0.016491f
C409 VTAIL.n368 B 0.015544f
C410 VTAIL.n369 B 0.009303f
C411 VTAIL.n370 B 0.786349f
C412 VTAIL.n371 B 0.017312f
C413 VTAIL.n372 B 0.009303f
C414 VTAIL.n373 B 0.00985f
C415 VTAIL.n374 B 0.021988f
C416 VTAIL.n375 B 0.021988f
C417 VTAIL.n376 B 0.00985f
C418 VTAIL.n377 B 0.009303f
C419 VTAIL.n378 B 0.017312f
C420 VTAIL.n379 B 0.017312f
C421 VTAIL.n380 B 0.009303f
C422 VTAIL.n381 B 0.00985f
C423 VTAIL.n382 B 0.021988f
C424 VTAIL.n383 B 0.021988f
C425 VTAIL.n384 B 0.00985f
C426 VTAIL.n385 B 0.009303f
C427 VTAIL.n386 B 0.017312f
C428 VTAIL.n387 B 0.017312f
C429 VTAIL.n388 B 0.009303f
C430 VTAIL.n389 B 0.009576f
C431 VTAIL.n390 B 0.009576f
C432 VTAIL.n391 B 0.021988f
C433 VTAIL.n392 B 0.021988f
C434 VTAIL.n393 B 0.00985f
C435 VTAIL.n394 B 0.009303f
C436 VTAIL.n395 B 0.017312f
C437 VTAIL.n396 B 0.017312f
C438 VTAIL.n397 B 0.009303f
C439 VTAIL.n398 B 0.00985f
C440 VTAIL.n399 B 0.021988f
C441 VTAIL.n400 B 0.049873f
C442 VTAIL.n401 B 0.00985f
C443 VTAIL.n402 B 0.009303f
C444 VTAIL.n403 B 0.044509f
C445 VTAIL.n404 B 0.028271f
C446 VTAIL.n405 B 1.13108f
C447 VTAIL.n406 B 0.025618f
C448 VTAIL.n407 B 0.017312f
C449 VTAIL.n408 B 0.009303f
C450 VTAIL.n409 B 0.021988f
C451 VTAIL.n410 B 0.00985f
C452 VTAIL.n411 B 0.017312f
C453 VTAIL.n412 B 0.009303f
C454 VTAIL.n413 B 0.021988f
C455 VTAIL.n414 B 0.00985f
C456 VTAIL.n415 B 0.017312f
C457 VTAIL.n416 B 0.009303f
C458 VTAIL.n417 B 0.021988f
C459 VTAIL.n418 B 0.00985f
C460 VTAIL.n419 B 0.017312f
C461 VTAIL.n420 B 0.009303f
C462 VTAIL.n421 B 0.021988f
C463 VTAIL.n422 B 0.00985f
C464 VTAIL.n423 B 0.117309f
C465 VTAIL.t6 B 0.037032f
C466 VTAIL.n424 B 0.016491f
C467 VTAIL.n425 B 0.015544f
C468 VTAIL.n426 B 0.009303f
C469 VTAIL.n427 B 0.786349f
C470 VTAIL.n428 B 0.017312f
C471 VTAIL.n429 B 0.009303f
C472 VTAIL.n430 B 0.00985f
C473 VTAIL.n431 B 0.021988f
C474 VTAIL.n432 B 0.021988f
C475 VTAIL.n433 B 0.00985f
C476 VTAIL.n434 B 0.009303f
C477 VTAIL.n435 B 0.017312f
C478 VTAIL.n436 B 0.017312f
C479 VTAIL.n437 B 0.009303f
C480 VTAIL.n438 B 0.00985f
C481 VTAIL.n439 B 0.021988f
C482 VTAIL.n440 B 0.021988f
C483 VTAIL.n441 B 0.021988f
C484 VTAIL.n442 B 0.00985f
C485 VTAIL.n443 B 0.009303f
C486 VTAIL.n444 B 0.017312f
C487 VTAIL.n445 B 0.017312f
C488 VTAIL.n446 B 0.009303f
C489 VTAIL.n447 B 0.009576f
C490 VTAIL.n448 B 0.009576f
C491 VTAIL.n449 B 0.021988f
C492 VTAIL.n450 B 0.021988f
C493 VTAIL.n451 B 0.00985f
C494 VTAIL.n452 B 0.009303f
C495 VTAIL.n453 B 0.017312f
C496 VTAIL.n454 B 0.017312f
C497 VTAIL.n455 B 0.009303f
C498 VTAIL.n456 B 0.00985f
C499 VTAIL.n457 B 0.021988f
C500 VTAIL.n458 B 0.049873f
C501 VTAIL.n459 B 0.00985f
C502 VTAIL.n460 B 0.009303f
C503 VTAIL.n461 B 0.044509f
C504 VTAIL.n462 B 0.028271f
C505 VTAIL.n463 B 1.03887f
C506 VP.t0 B 2.21953f
C507 VP.n0 B 0.876889f
C508 VP.n1 B 0.022304f
C509 VP.n2 B 0.018031f
C510 VP.n3 B 0.022304f
C511 VP.t1 B 2.21953f
C512 VP.n4 B 0.876889f
C513 VP.t3 B 2.51697f
C514 VP.t2 B 2.5078f
C515 VP.n5 B 2.85578f
C516 VP.n6 B 1.28077f
C517 VP.n7 B 0.035999f
C518 VP.n8 B 0.035412f
C519 VP.n9 B 0.041569f
C520 VP.n10 B 0.044329f
C521 VP.n11 B 0.022304f
C522 VP.n12 B 0.022304f
C523 VP.n13 B 0.022304f
C524 VP.n14 B 0.044329f
C525 VP.n15 B 0.041569f
C526 VP.n16 B 0.035412f
C527 VP.n17 B 0.035999f
C528 VP.n18 B 0.052241f
.ends

