# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_9T_clkbuf_16
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_9T_clkbuf_16 0 0 ;
  SIZE 15.8 BY 6.15 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.05 2.2 1.55 2.5 ;
      LAYER MET2 ;
        RECT 1.05 2.2 1.55 2.5 ;
        RECT 1.1 2.15 1.5 2.55 ;
      LAYER VIA12 ;
        RECT 1.17 2.22 1.43 2.48 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 5.55 15.8 6.15 ;
        RECT 15 3.5 15.25 6.15 ;
        RECT 13.3 3.5 13.55 6.15 ;
        RECT 11.6 3.5 11.85 6.15 ;
        RECT 9.9 3.5 10.15 6.15 ;
        RECT 8.2 3.5 8.45 6.15 ;
        RECT 6.5 3.5 6.75 6.15 ;
        RECT 4.8 3.5 5.05 6.15 ;
        RECT 3.1 3.5 3.35 6.15 ;
        RECT 1.4 3.5 1.65 6.15 ;
      LAYER MET2 ;
        RECT 13.65 5.6 14.15 5.9 ;
        RECT 13.7 5.55 14.1 5.95 ;
        RECT 12.45 5.6 12.95 5.9 ;
        RECT 12.5 5.55 12.9 5.95 ;
        RECT 11.25 5.6 11.75 5.9 ;
        RECT 11.3 5.55 11.7 5.95 ;
        RECT 10.05 5.6 10.55 5.9 ;
        RECT 10.1 5.55 10.5 5.95 ;
        RECT 8.85 5.6 9.35 5.9 ;
        RECT 8.9 5.55 9.3 5.95 ;
        RECT 7.65 5.6 8.15 5.9 ;
        RECT 7.7 5.55 8.1 5.95 ;
        RECT 6.45 5.6 6.95 5.9 ;
        RECT 6.5 5.55 6.9 5.95 ;
        RECT 5.25 5.6 5.75 5.9 ;
        RECT 5.3 5.55 5.7 5.95 ;
        RECT 4.05 5.6 4.55 5.9 ;
        RECT 4.1 5.55 4.5 5.95 ;
        RECT 2.85 5.6 3.35 5.9 ;
        RECT 2.9 5.55 3.3 5.95 ;
        RECT 1.65 5.6 2.15 5.9 ;
        RECT 1.7 5.55 2.1 5.95 ;
        RECT 0.45 5.6 0.95 5.9 ;
        RECT 0.5 5.55 0.9 5.95 ;
      LAYER VIA12 ;
        RECT 0.57 5.62 0.83 5.88 ;
        RECT 1.77 5.62 2.03 5.88 ;
        RECT 2.97 5.62 3.23 5.88 ;
        RECT 4.17 5.62 4.43 5.88 ;
        RECT 5.37 5.62 5.63 5.88 ;
        RECT 6.57 5.62 6.83 5.88 ;
        RECT 7.77 5.62 8.03 5.88 ;
        RECT 8.97 5.62 9.23 5.88 ;
        RECT 10.17 5.62 10.43 5.88 ;
        RECT 11.37 5.62 11.63 5.88 ;
        RECT 12.57 5.62 12.83 5.88 ;
        RECT 13.77 5.62 14.03 5.88 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 15.8 0.6 ;
        RECT 15 0 15.25 1.8 ;
        RECT 13.3 0 13.55 1.8 ;
        RECT 11.6 0 11.85 1.8 ;
        RECT 9.9 0 10.15 1.8 ;
        RECT 8.2 0 8.45 1.8 ;
        RECT 6.5 0 6.75 1.8 ;
        RECT 4.8 0 5.05 1.8 ;
        RECT 3.1 0 3.35 1.8 ;
        RECT 1.4 0 1.65 1.8 ;
      LAYER MET2 ;
        RECT 13.65 0.25 14.15 0.55 ;
        RECT 13.7 0.2 14.1 0.6 ;
        RECT 12.45 0.25 12.95 0.55 ;
        RECT 12.5 0.2 12.9 0.6 ;
        RECT 11.25 0.25 11.75 0.55 ;
        RECT 11.3 0.2 11.7 0.6 ;
        RECT 10.05 0.25 10.55 0.55 ;
        RECT 10.1 0.2 10.5 0.6 ;
        RECT 8.85 0.25 9.35 0.55 ;
        RECT 8.9 0.2 9.3 0.6 ;
        RECT 7.65 0.25 8.15 0.55 ;
        RECT 7.7 0.2 8.1 0.6 ;
        RECT 6.45 0.25 6.95 0.55 ;
        RECT 6.5 0.2 6.9 0.6 ;
        RECT 5.25 0.25 5.75 0.55 ;
        RECT 5.3 0.2 5.7 0.6 ;
        RECT 4.05 0.25 4.55 0.55 ;
        RECT 4.1 0.2 4.5 0.6 ;
        RECT 2.85 0.25 3.35 0.55 ;
        RECT 2.9 0.2 3.3 0.6 ;
        RECT 1.65 0.25 2.15 0.55 ;
        RECT 1.7 0.2 2.1 0.6 ;
        RECT 0.45 0.25 0.95 0.55 ;
        RECT 0.5 0.2 0.9 0.6 ;
      LAYER VIA12 ;
        RECT 0.57 0.27 0.83 0.53 ;
        RECT 1.77 0.27 2.03 0.53 ;
        RECT 2.97 0.27 3.23 0.53 ;
        RECT 4.17 0.27 4.43 0.53 ;
        RECT 5.37 0.27 5.63 0.53 ;
        RECT 6.57 0.27 6.83 0.53 ;
        RECT 7.77 0.27 8.03 0.53 ;
        RECT 8.97 0.27 9.23 0.53 ;
        RECT 10.17 0.27 10.43 0.53 ;
        RECT 11.37 0.27 11.63 0.53 ;
        RECT 12.57 0.27 12.83 0.53 ;
        RECT 13.77 0.27 14.03 0.53 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 14.05 3.5 14.55 3.8 ;
        RECT 14.15 0.95 14.4 5.2 ;
        RECT 2.25 2.95 14.4 3.25 ;
        RECT 2.25 2.05 14.4 2.35 ;
        RECT 12.45 0.95 12.7 5.2 ;
        RECT 10.75 0.95 11 5.2 ;
        RECT 9.05 0.95 9.3 5.2 ;
        RECT 7.35 0.95 7.6 5.2 ;
        RECT 5.65 0.95 5.9 5.2 ;
        RECT 3.95 0.95 4.2 5.2 ;
        RECT 2.25 0.95 2.5 5.2 ;
      LAYER MET2 ;
        RECT 14.05 3.45 14.55 3.85 ;
      LAYER VIA12 ;
        RECT 14.17 3.52 14.43 3.78 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.55 0.95 0.8 5.2 ;
      RECT 0.55 2.95 2 3.25 ;
  END
END gf180mcu_osu_sc_9T_clkbuf_16
