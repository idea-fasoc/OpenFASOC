* NGSPICE file created from diff_pair_sample_1758.ext - technology: sky130A

.subckt diff_pair_sample_1758 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t7 VN.t0 VTAIL.t9 B.t1 sky130_fd_pr__nfet_01v8 ad=3.14985 pd=19.42 as=7.4451 ps=38.96 w=19.09 l=2.39
X1 VTAIL.t12 VN.t1 VDD2.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=3.14985 pd=19.42 as=3.14985 ps=19.42 w=19.09 l=2.39
X2 VDD1.t7 VP.t0 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=3.14985 pd=19.42 as=7.4451 ps=38.96 w=19.09 l=2.39
X3 VTAIL.t5 VP.t1 VDD1.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=7.4451 pd=38.96 as=3.14985 ps=19.42 w=19.09 l=2.39
X4 VTAIL.t7 VP.t2 VDD1.t5 B.t7 sky130_fd_pr__nfet_01v8 ad=7.4451 pd=38.96 as=3.14985 ps=19.42 w=19.09 l=2.39
X5 B.t21 B.t19 B.t20 B.t9 sky130_fd_pr__nfet_01v8 ad=7.4451 pd=38.96 as=0 ps=0 w=19.09 l=2.39
X6 VDD1.t4 VP.t3 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=3.14985 pd=19.42 as=3.14985 ps=19.42 w=19.09 l=2.39
X7 VTAIL.t8 VN.t2 VDD2.t5 B.t7 sky130_fd_pr__nfet_01v8 ad=7.4451 pd=38.96 as=3.14985 ps=19.42 w=19.09 l=2.39
X8 VDD2.t4 VN.t3 VTAIL.t14 B.t0 sky130_fd_pr__nfet_01v8 ad=3.14985 pd=19.42 as=3.14985 ps=19.42 w=19.09 l=2.39
X9 B.t18 B.t16 B.t17 B.t13 sky130_fd_pr__nfet_01v8 ad=7.4451 pd=38.96 as=0 ps=0 w=19.09 l=2.39
X10 VDD2.t3 VN.t4 VTAIL.t15 B.t6 sky130_fd_pr__nfet_01v8 ad=3.14985 pd=19.42 as=3.14985 ps=19.42 w=19.09 l=2.39
X11 VTAIL.t4 VP.t4 VDD1.t3 B.t4 sky130_fd_pr__nfet_01v8 ad=3.14985 pd=19.42 as=3.14985 ps=19.42 w=19.09 l=2.39
X12 VTAIL.t10 VN.t5 VDD2.t2 B.t5 sky130_fd_pr__nfet_01v8 ad=7.4451 pd=38.96 as=3.14985 ps=19.42 w=19.09 l=2.39
X13 VDD1.t2 VP.t5 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=3.14985 pd=19.42 as=7.4451 ps=38.96 w=19.09 l=2.39
X14 VDD2.t1 VN.t6 VTAIL.t11 B.t2 sky130_fd_pr__nfet_01v8 ad=3.14985 pd=19.42 as=7.4451 ps=38.96 w=19.09 l=2.39
X15 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=7.4451 pd=38.96 as=0 ps=0 w=19.09 l=2.39
X16 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=7.4451 pd=38.96 as=0 ps=0 w=19.09 l=2.39
X17 VTAIL.t3 VP.t6 VDD1.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=3.14985 pd=19.42 as=3.14985 ps=19.42 w=19.09 l=2.39
X18 VDD1.t0 VP.t7 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=3.14985 pd=19.42 as=3.14985 ps=19.42 w=19.09 l=2.39
X19 VTAIL.t13 VN.t7 VDD2.t0 B.t4 sky130_fd_pr__nfet_01v8 ad=3.14985 pd=19.42 as=3.14985 ps=19.42 w=19.09 l=2.39
R0 VN.n7 VN.t2 225.333
R1 VN.n34 VN.t6 225.333
R2 VN.n6 VN.t4 192.498
R3 VN.n17 VN.t1 192.498
R4 VN.n25 VN.t0 192.498
R5 VN.n33 VN.t7 192.498
R6 VN.n44 VN.t3 192.498
R7 VN.n52 VN.t5 192.498
R8 VN.n51 VN.n27 161.3
R9 VN.n50 VN.n49 161.3
R10 VN.n48 VN.n28 161.3
R11 VN.n47 VN.n46 161.3
R12 VN.n45 VN.n29 161.3
R13 VN.n43 VN.n42 161.3
R14 VN.n41 VN.n30 161.3
R15 VN.n40 VN.n39 161.3
R16 VN.n38 VN.n31 161.3
R17 VN.n37 VN.n36 161.3
R18 VN.n35 VN.n32 161.3
R19 VN.n24 VN.n0 161.3
R20 VN.n23 VN.n22 161.3
R21 VN.n21 VN.n1 161.3
R22 VN.n20 VN.n19 161.3
R23 VN.n18 VN.n2 161.3
R24 VN.n16 VN.n15 161.3
R25 VN.n14 VN.n3 161.3
R26 VN.n13 VN.n12 161.3
R27 VN.n11 VN.n4 161.3
R28 VN.n10 VN.n9 161.3
R29 VN.n8 VN.n5 161.3
R30 VN.n26 VN.n25 94.6082
R31 VN.n53 VN.n52 94.6082
R32 VN.n7 VN.n6 66.7382
R33 VN.n34 VN.n33 66.7382
R34 VN.n12 VN.n11 56.5193
R35 VN.n39 VN.n38 56.5193
R36 VN VN.n53 55.6269
R37 VN.n19 VN.n1 43.4072
R38 VN.n46 VN.n28 43.4072
R39 VN.n23 VN.n1 37.5796
R40 VN.n50 VN.n28 37.5796
R41 VN.n10 VN.n5 24.4675
R42 VN.n11 VN.n10 24.4675
R43 VN.n12 VN.n3 24.4675
R44 VN.n16 VN.n3 24.4675
R45 VN.n19 VN.n18 24.4675
R46 VN.n24 VN.n23 24.4675
R47 VN.n38 VN.n37 24.4675
R48 VN.n37 VN.n32 24.4675
R49 VN.n46 VN.n45 24.4675
R50 VN.n43 VN.n30 24.4675
R51 VN.n39 VN.n30 24.4675
R52 VN.n51 VN.n50 24.4675
R53 VN.n18 VN.n17 19.0848
R54 VN.n45 VN.n44 19.0848
R55 VN.n25 VN.n24 16.1487
R56 VN.n52 VN.n51 16.1487
R57 VN.n35 VN.n34 9.37577
R58 VN.n8 VN.n7 9.37577
R59 VN.n6 VN.n5 5.38324
R60 VN.n17 VN.n16 5.38324
R61 VN.n33 VN.n32 5.38324
R62 VN.n44 VN.n43 5.38324
R63 VN.n53 VN.n27 0.278367
R64 VN.n26 VN.n0 0.278367
R65 VN.n49 VN.n27 0.189894
R66 VN.n49 VN.n48 0.189894
R67 VN.n48 VN.n47 0.189894
R68 VN.n47 VN.n29 0.189894
R69 VN.n42 VN.n29 0.189894
R70 VN.n42 VN.n41 0.189894
R71 VN.n41 VN.n40 0.189894
R72 VN.n40 VN.n31 0.189894
R73 VN.n36 VN.n31 0.189894
R74 VN.n36 VN.n35 0.189894
R75 VN.n9 VN.n8 0.189894
R76 VN.n9 VN.n4 0.189894
R77 VN.n13 VN.n4 0.189894
R78 VN.n14 VN.n13 0.189894
R79 VN.n15 VN.n14 0.189894
R80 VN.n15 VN.n2 0.189894
R81 VN.n20 VN.n2 0.189894
R82 VN.n21 VN.n20 0.189894
R83 VN.n22 VN.n21 0.189894
R84 VN.n22 VN.n0 0.189894
R85 VN VN.n26 0.153454
R86 VTAIL.n11 VTAIL.t7 47.0791
R87 VTAIL.n10 VTAIL.t11 47.0791
R88 VTAIL.n7 VTAIL.t10 47.0791
R89 VTAIL.n15 VTAIL.t9 47.079
R90 VTAIL.n2 VTAIL.t8 47.079
R91 VTAIL.n3 VTAIL.t2 47.079
R92 VTAIL.n6 VTAIL.t5 47.079
R93 VTAIL.n14 VTAIL.t1 47.079
R94 VTAIL.n13 VTAIL.n12 46.042
R95 VTAIL.n9 VTAIL.n8 46.042
R96 VTAIL.n1 VTAIL.n0 46.0408
R97 VTAIL.n5 VTAIL.n4 46.0408
R98 VTAIL.n15 VTAIL.n14 31.1686
R99 VTAIL.n7 VTAIL.n6 31.1686
R100 VTAIL.n9 VTAIL.n7 2.34533
R101 VTAIL.n10 VTAIL.n9 2.34533
R102 VTAIL.n13 VTAIL.n11 2.34533
R103 VTAIL.n14 VTAIL.n13 2.34533
R104 VTAIL.n6 VTAIL.n5 2.34533
R105 VTAIL.n5 VTAIL.n3 2.34533
R106 VTAIL.n2 VTAIL.n1 2.34533
R107 VTAIL VTAIL.n15 2.28714
R108 VTAIL.n0 VTAIL.t15 1.03769
R109 VTAIL.n0 VTAIL.t12 1.03769
R110 VTAIL.n4 VTAIL.t0 1.03769
R111 VTAIL.n4 VTAIL.t4 1.03769
R112 VTAIL.n12 VTAIL.t6 1.03769
R113 VTAIL.n12 VTAIL.t3 1.03769
R114 VTAIL.n8 VTAIL.t14 1.03769
R115 VTAIL.n8 VTAIL.t13 1.03769
R116 VTAIL.n11 VTAIL.n10 0.470328
R117 VTAIL.n3 VTAIL.n2 0.470328
R118 VTAIL VTAIL.n1 0.0586897
R119 VDD2.n2 VDD2.n1 63.8366
R120 VDD2.n2 VDD2.n0 63.8366
R121 VDD2 VDD2.n5 63.8348
R122 VDD2.n4 VDD2.n3 62.7207
R123 VDD2.n4 VDD2.n2 50.7239
R124 VDD2 VDD2.n4 1.2311
R125 VDD2.n5 VDD2.t0 1.03769
R126 VDD2.n5 VDD2.t1 1.03769
R127 VDD2.n3 VDD2.t2 1.03769
R128 VDD2.n3 VDD2.t4 1.03769
R129 VDD2.n1 VDD2.t6 1.03769
R130 VDD2.n1 VDD2.t7 1.03769
R131 VDD2.n0 VDD2.t5 1.03769
R132 VDD2.n0 VDD2.t3 1.03769
R133 B.n1072 B.n1071 585
R134 B.n1073 B.n1072 585
R135 B.n428 B.n157 585
R136 B.n427 B.n426 585
R137 B.n425 B.n424 585
R138 B.n423 B.n422 585
R139 B.n421 B.n420 585
R140 B.n419 B.n418 585
R141 B.n417 B.n416 585
R142 B.n415 B.n414 585
R143 B.n413 B.n412 585
R144 B.n411 B.n410 585
R145 B.n409 B.n408 585
R146 B.n407 B.n406 585
R147 B.n405 B.n404 585
R148 B.n403 B.n402 585
R149 B.n401 B.n400 585
R150 B.n399 B.n398 585
R151 B.n397 B.n396 585
R152 B.n395 B.n394 585
R153 B.n393 B.n392 585
R154 B.n391 B.n390 585
R155 B.n389 B.n388 585
R156 B.n387 B.n386 585
R157 B.n385 B.n384 585
R158 B.n383 B.n382 585
R159 B.n381 B.n380 585
R160 B.n379 B.n378 585
R161 B.n377 B.n376 585
R162 B.n375 B.n374 585
R163 B.n373 B.n372 585
R164 B.n371 B.n370 585
R165 B.n369 B.n368 585
R166 B.n367 B.n366 585
R167 B.n365 B.n364 585
R168 B.n363 B.n362 585
R169 B.n361 B.n360 585
R170 B.n359 B.n358 585
R171 B.n357 B.n356 585
R172 B.n355 B.n354 585
R173 B.n353 B.n352 585
R174 B.n351 B.n350 585
R175 B.n349 B.n348 585
R176 B.n347 B.n346 585
R177 B.n345 B.n344 585
R178 B.n343 B.n342 585
R179 B.n341 B.n340 585
R180 B.n339 B.n338 585
R181 B.n337 B.n336 585
R182 B.n335 B.n334 585
R183 B.n333 B.n332 585
R184 B.n331 B.n330 585
R185 B.n329 B.n328 585
R186 B.n327 B.n326 585
R187 B.n325 B.n324 585
R188 B.n323 B.n322 585
R189 B.n321 B.n320 585
R190 B.n319 B.n318 585
R191 B.n317 B.n316 585
R192 B.n315 B.n314 585
R193 B.n313 B.n312 585
R194 B.n311 B.n310 585
R195 B.n309 B.n308 585
R196 B.n307 B.n306 585
R197 B.n305 B.n304 585
R198 B.n303 B.n302 585
R199 B.n301 B.n300 585
R200 B.n299 B.n298 585
R201 B.n297 B.n296 585
R202 B.n295 B.n294 585
R203 B.n293 B.n292 585
R204 B.n291 B.n290 585
R205 B.n289 B.n288 585
R206 B.n286 B.n285 585
R207 B.n284 B.n283 585
R208 B.n282 B.n281 585
R209 B.n280 B.n279 585
R210 B.n278 B.n277 585
R211 B.n276 B.n275 585
R212 B.n274 B.n273 585
R213 B.n272 B.n271 585
R214 B.n270 B.n269 585
R215 B.n268 B.n267 585
R216 B.n266 B.n265 585
R217 B.n264 B.n263 585
R218 B.n262 B.n261 585
R219 B.n260 B.n259 585
R220 B.n258 B.n257 585
R221 B.n256 B.n255 585
R222 B.n254 B.n253 585
R223 B.n252 B.n251 585
R224 B.n250 B.n249 585
R225 B.n248 B.n247 585
R226 B.n246 B.n245 585
R227 B.n244 B.n243 585
R228 B.n242 B.n241 585
R229 B.n240 B.n239 585
R230 B.n238 B.n237 585
R231 B.n236 B.n235 585
R232 B.n234 B.n233 585
R233 B.n232 B.n231 585
R234 B.n230 B.n229 585
R235 B.n228 B.n227 585
R236 B.n226 B.n225 585
R237 B.n224 B.n223 585
R238 B.n222 B.n221 585
R239 B.n220 B.n219 585
R240 B.n218 B.n217 585
R241 B.n216 B.n215 585
R242 B.n214 B.n213 585
R243 B.n212 B.n211 585
R244 B.n210 B.n209 585
R245 B.n208 B.n207 585
R246 B.n206 B.n205 585
R247 B.n204 B.n203 585
R248 B.n202 B.n201 585
R249 B.n200 B.n199 585
R250 B.n198 B.n197 585
R251 B.n196 B.n195 585
R252 B.n194 B.n193 585
R253 B.n192 B.n191 585
R254 B.n190 B.n189 585
R255 B.n188 B.n187 585
R256 B.n186 B.n185 585
R257 B.n184 B.n183 585
R258 B.n182 B.n181 585
R259 B.n180 B.n179 585
R260 B.n178 B.n177 585
R261 B.n176 B.n175 585
R262 B.n174 B.n173 585
R263 B.n172 B.n171 585
R264 B.n170 B.n169 585
R265 B.n168 B.n167 585
R266 B.n166 B.n165 585
R267 B.n164 B.n163 585
R268 B.n88 B.n87 585
R269 B.n1070 B.n89 585
R270 B.n1074 B.n89 585
R271 B.n1069 B.n1068 585
R272 B.n1068 B.n85 585
R273 B.n1067 B.n84 585
R274 B.n1080 B.n84 585
R275 B.n1066 B.n83 585
R276 B.n1081 B.n83 585
R277 B.n1065 B.n82 585
R278 B.n1082 B.n82 585
R279 B.n1064 B.n1063 585
R280 B.n1063 B.n78 585
R281 B.n1062 B.n77 585
R282 B.n1088 B.n77 585
R283 B.n1061 B.n76 585
R284 B.n1089 B.n76 585
R285 B.n1060 B.n75 585
R286 B.n1090 B.n75 585
R287 B.n1059 B.n1058 585
R288 B.n1058 B.n71 585
R289 B.n1057 B.n70 585
R290 B.n1096 B.n70 585
R291 B.n1056 B.n69 585
R292 B.n1097 B.n69 585
R293 B.n1055 B.n68 585
R294 B.n1098 B.n68 585
R295 B.n1054 B.n1053 585
R296 B.n1053 B.n64 585
R297 B.n1052 B.n63 585
R298 B.n1104 B.n63 585
R299 B.n1051 B.n62 585
R300 B.n1105 B.n62 585
R301 B.n1050 B.n61 585
R302 B.n1106 B.n61 585
R303 B.n1049 B.n1048 585
R304 B.n1048 B.n57 585
R305 B.n1047 B.n56 585
R306 B.n1112 B.n56 585
R307 B.n1046 B.n55 585
R308 B.n1113 B.n55 585
R309 B.n1045 B.n54 585
R310 B.n1114 B.n54 585
R311 B.n1044 B.n1043 585
R312 B.n1043 B.n50 585
R313 B.n1042 B.n49 585
R314 B.n1120 B.n49 585
R315 B.n1041 B.n48 585
R316 B.n1121 B.n48 585
R317 B.n1040 B.n47 585
R318 B.n1122 B.n47 585
R319 B.n1039 B.n1038 585
R320 B.n1038 B.n43 585
R321 B.n1037 B.n42 585
R322 B.n1128 B.n42 585
R323 B.n1036 B.n41 585
R324 B.n1129 B.n41 585
R325 B.n1035 B.n40 585
R326 B.n1130 B.n40 585
R327 B.n1034 B.n1033 585
R328 B.n1033 B.n36 585
R329 B.n1032 B.n35 585
R330 B.n1136 B.n35 585
R331 B.n1031 B.n34 585
R332 B.n1137 B.n34 585
R333 B.n1030 B.n33 585
R334 B.n1138 B.n33 585
R335 B.n1029 B.n1028 585
R336 B.n1028 B.n29 585
R337 B.n1027 B.n28 585
R338 B.n1144 B.n28 585
R339 B.n1026 B.n27 585
R340 B.n1145 B.n27 585
R341 B.n1025 B.n26 585
R342 B.n1146 B.n26 585
R343 B.n1024 B.n1023 585
R344 B.n1023 B.n22 585
R345 B.n1022 B.n21 585
R346 B.n1152 B.n21 585
R347 B.n1021 B.n20 585
R348 B.n1153 B.n20 585
R349 B.n1020 B.n19 585
R350 B.n1154 B.n19 585
R351 B.n1019 B.n1018 585
R352 B.n1018 B.n15 585
R353 B.n1017 B.n14 585
R354 B.n1160 B.n14 585
R355 B.n1016 B.n13 585
R356 B.n1161 B.n13 585
R357 B.n1015 B.n12 585
R358 B.n1162 B.n12 585
R359 B.n1014 B.n1013 585
R360 B.n1013 B.n8 585
R361 B.n1012 B.n7 585
R362 B.n1168 B.n7 585
R363 B.n1011 B.n6 585
R364 B.n1169 B.n6 585
R365 B.n1010 B.n5 585
R366 B.n1170 B.n5 585
R367 B.n1009 B.n1008 585
R368 B.n1008 B.n4 585
R369 B.n1007 B.n429 585
R370 B.n1007 B.n1006 585
R371 B.n997 B.n430 585
R372 B.n431 B.n430 585
R373 B.n999 B.n998 585
R374 B.n1000 B.n999 585
R375 B.n996 B.n436 585
R376 B.n436 B.n435 585
R377 B.n995 B.n994 585
R378 B.n994 B.n993 585
R379 B.n438 B.n437 585
R380 B.n439 B.n438 585
R381 B.n986 B.n985 585
R382 B.n987 B.n986 585
R383 B.n984 B.n444 585
R384 B.n444 B.n443 585
R385 B.n983 B.n982 585
R386 B.n982 B.n981 585
R387 B.n446 B.n445 585
R388 B.n447 B.n446 585
R389 B.n974 B.n973 585
R390 B.n975 B.n974 585
R391 B.n972 B.n452 585
R392 B.n452 B.n451 585
R393 B.n971 B.n970 585
R394 B.n970 B.n969 585
R395 B.n454 B.n453 585
R396 B.n455 B.n454 585
R397 B.n962 B.n961 585
R398 B.n963 B.n962 585
R399 B.n960 B.n460 585
R400 B.n460 B.n459 585
R401 B.n959 B.n958 585
R402 B.n958 B.n957 585
R403 B.n462 B.n461 585
R404 B.n463 B.n462 585
R405 B.n950 B.n949 585
R406 B.n951 B.n950 585
R407 B.n948 B.n468 585
R408 B.n468 B.n467 585
R409 B.n947 B.n946 585
R410 B.n946 B.n945 585
R411 B.n470 B.n469 585
R412 B.n471 B.n470 585
R413 B.n938 B.n937 585
R414 B.n939 B.n938 585
R415 B.n936 B.n476 585
R416 B.n476 B.n475 585
R417 B.n935 B.n934 585
R418 B.n934 B.n933 585
R419 B.n478 B.n477 585
R420 B.n479 B.n478 585
R421 B.n926 B.n925 585
R422 B.n927 B.n926 585
R423 B.n924 B.n484 585
R424 B.n484 B.n483 585
R425 B.n923 B.n922 585
R426 B.n922 B.n921 585
R427 B.n486 B.n485 585
R428 B.n487 B.n486 585
R429 B.n914 B.n913 585
R430 B.n915 B.n914 585
R431 B.n912 B.n492 585
R432 B.n492 B.n491 585
R433 B.n911 B.n910 585
R434 B.n910 B.n909 585
R435 B.n494 B.n493 585
R436 B.n495 B.n494 585
R437 B.n902 B.n901 585
R438 B.n903 B.n902 585
R439 B.n900 B.n500 585
R440 B.n500 B.n499 585
R441 B.n899 B.n898 585
R442 B.n898 B.n897 585
R443 B.n502 B.n501 585
R444 B.n503 B.n502 585
R445 B.n890 B.n889 585
R446 B.n891 B.n890 585
R447 B.n888 B.n507 585
R448 B.n511 B.n507 585
R449 B.n887 B.n886 585
R450 B.n886 B.n885 585
R451 B.n509 B.n508 585
R452 B.n510 B.n509 585
R453 B.n878 B.n877 585
R454 B.n879 B.n878 585
R455 B.n876 B.n516 585
R456 B.n516 B.n515 585
R457 B.n875 B.n874 585
R458 B.n874 B.n873 585
R459 B.n518 B.n517 585
R460 B.n519 B.n518 585
R461 B.n866 B.n865 585
R462 B.n867 B.n866 585
R463 B.n522 B.n521 585
R464 B.n595 B.n594 585
R465 B.n596 B.n592 585
R466 B.n592 B.n523 585
R467 B.n598 B.n597 585
R468 B.n600 B.n591 585
R469 B.n603 B.n602 585
R470 B.n604 B.n590 585
R471 B.n606 B.n605 585
R472 B.n608 B.n589 585
R473 B.n611 B.n610 585
R474 B.n612 B.n588 585
R475 B.n614 B.n613 585
R476 B.n616 B.n587 585
R477 B.n619 B.n618 585
R478 B.n620 B.n586 585
R479 B.n622 B.n621 585
R480 B.n624 B.n585 585
R481 B.n627 B.n626 585
R482 B.n628 B.n584 585
R483 B.n630 B.n629 585
R484 B.n632 B.n583 585
R485 B.n635 B.n634 585
R486 B.n636 B.n582 585
R487 B.n638 B.n637 585
R488 B.n640 B.n581 585
R489 B.n643 B.n642 585
R490 B.n644 B.n580 585
R491 B.n646 B.n645 585
R492 B.n648 B.n579 585
R493 B.n651 B.n650 585
R494 B.n652 B.n578 585
R495 B.n654 B.n653 585
R496 B.n656 B.n577 585
R497 B.n659 B.n658 585
R498 B.n660 B.n576 585
R499 B.n662 B.n661 585
R500 B.n664 B.n575 585
R501 B.n667 B.n666 585
R502 B.n668 B.n574 585
R503 B.n670 B.n669 585
R504 B.n672 B.n573 585
R505 B.n675 B.n674 585
R506 B.n676 B.n572 585
R507 B.n678 B.n677 585
R508 B.n680 B.n571 585
R509 B.n683 B.n682 585
R510 B.n684 B.n570 585
R511 B.n686 B.n685 585
R512 B.n688 B.n569 585
R513 B.n691 B.n690 585
R514 B.n692 B.n568 585
R515 B.n694 B.n693 585
R516 B.n696 B.n567 585
R517 B.n699 B.n698 585
R518 B.n700 B.n566 585
R519 B.n702 B.n701 585
R520 B.n704 B.n565 585
R521 B.n707 B.n706 585
R522 B.n708 B.n564 585
R523 B.n710 B.n709 585
R524 B.n712 B.n563 585
R525 B.n715 B.n714 585
R526 B.n716 B.n560 585
R527 B.n719 B.n718 585
R528 B.n721 B.n559 585
R529 B.n724 B.n723 585
R530 B.n725 B.n558 585
R531 B.n727 B.n726 585
R532 B.n729 B.n557 585
R533 B.n732 B.n731 585
R534 B.n733 B.n556 585
R535 B.n738 B.n737 585
R536 B.n740 B.n555 585
R537 B.n743 B.n742 585
R538 B.n744 B.n554 585
R539 B.n746 B.n745 585
R540 B.n748 B.n553 585
R541 B.n751 B.n750 585
R542 B.n752 B.n552 585
R543 B.n754 B.n753 585
R544 B.n756 B.n551 585
R545 B.n759 B.n758 585
R546 B.n760 B.n550 585
R547 B.n762 B.n761 585
R548 B.n764 B.n549 585
R549 B.n767 B.n766 585
R550 B.n768 B.n548 585
R551 B.n770 B.n769 585
R552 B.n772 B.n547 585
R553 B.n775 B.n774 585
R554 B.n776 B.n546 585
R555 B.n778 B.n777 585
R556 B.n780 B.n545 585
R557 B.n783 B.n782 585
R558 B.n784 B.n544 585
R559 B.n786 B.n785 585
R560 B.n788 B.n543 585
R561 B.n791 B.n790 585
R562 B.n792 B.n542 585
R563 B.n794 B.n793 585
R564 B.n796 B.n541 585
R565 B.n799 B.n798 585
R566 B.n800 B.n540 585
R567 B.n802 B.n801 585
R568 B.n804 B.n539 585
R569 B.n807 B.n806 585
R570 B.n808 B.n538 585
R571 B.n810 B.n809 585
R572 B.n812 B.n537 585
R573 B.n815 B.n814 585
R574 B.n816 B.n536 585
R575 B.n818 B.n817 585
R576 B.n820 B.n535 585
R577 B.n823 B.n822 585
R578 B.n824 B.n534 585
R579 B.n826 B.n825 585
R580 B.n828 B.n533 585
R581 B.n831 B.n830 585
R582 B.n832 B.n532 585
R583 B.n834 B.n833 585
R584 B.n836 B.n531 585
R585 B.n839 B.n838 585
R586 B.n840 B.n530 585
R587 B.n842 B.n841 585
R588 B.n844 B.n529 585
R589 B.n847 B.n846 585
R590 B.n848 B.n528 585
R591 B.n850 B.n849 585
R592 B.n852 B.n527 585
R593 B.n855 B.n854 585
R594 B.n856 B.n526 585
R595 B.n858 B.n857 585
R596 B.n860 B.n525 585
R597 B.n863 B.n862 585
R598 B.n864 B.n524 585
R599 B.n869 B.n868 585
R600 B.n868 B.n867 585
R601 B.n870 B.n520 585
R602 B.n520 B.n519 585
R603 B.n872 B.n871 585
R604 B.n873 B.n872 585
R605 B.n514 B.n513 585
R606 B.n515 B.n514 585
R607 B.n881 B.n880 585
R608 B.n880 B.n879 585
R609 B.n882 B.n512 585
R610 B.n512 B.n510 585
R611 B.n884 B.n883 585
R612 B.n885 B.n884 585
R613 B.n506 B.n505 585
R614 B.n511 B.n506 585
R615 B.n893 B.n892 585
R616 B.n892 B.n891 585
R617 B.n894 B.n504 585
R618 B.n504 B.n503 585
R619 B.n896 B.n895 585
R620 B.n897 B.n896 585
R621 B.n498 B.n497 585
R622 B.n499 B.n498 585
R623 B.n905 B.n904 585
R624 B.n904 B.n903 585
R625 B.n906 B.n496 585
R626 B.n496 B.n495 585
R627 B.n908 B.n907 585
R628 B.n909 B.n908 585
R629 B.n490 B.n489 585
R630 B.n491 B.n490 585
R631 B.n917 B.n916 585
R632 B.n916 B.n915 585
R633 B.n918 B.n488 585
R634 B.n488 B.n487 585
R635 B.n920 B.n919 585
R636 B.n921 B.n920 585
R637 B.n482 B.n481 585
R638 B.n483 B.n482 585
R639 B.n929 B.n928 585
R640 B.n928 B.n927 585
R641 B.n930 B.n480 585
R642 B.n480 B.n479 585
R643 B.n932 B.n931 585
R644 B.n933 B.n932 585
R645 B.n474 B.n473 585
R646 B.n475 B.n474 585
R647 B.n941 B.n940 585
R648 B.n940 B.n939 585
R649 B.n942 B.n472 585
R650 B.n472 B.n471 585
R651 B.n944 B.n943 585
R652 B.n945 B.n944 585
R653 B.n466 B.n465 585
R654 B.n467 B.n466 585
R655 B.n953 B.n952 585
R656 B.n952 B.n951 585
R657 B.n954 B.n464 585
R658 B.n464 B.n463 585
R659 B.n956 B.n955 585
R660 B.n957 B.n956 585
R661 B.n458 B.n457 585
R662 B.n459 B.n458 585
R663 B.n965 B.n964 585
R664 B.n964 B.n963 585
R665 B.n966 B.n456 585
R666 B.n456 B.n455 585
R667 B.n968 B.n967 585
R668 B.n969 B.n968 585
R669 B.n450 B.n449 585
R670 B.n451 B.n450 585
R671 B.n977 B.n976 585
R672 B.n976 B.n975 585
R673 B.n978 B.n448 585
R674 B.n448 B.n447 585
R675 B.n980 B.n979 585
R676 B.n981 B.n980 585
R677 B.n442 B.n441 585
R678 B.n443 B.n442 585
R679 B.n989 B.n988 585
R680 B.n988 B.n987 585
R681 B.n990 B.n440 585
R682 B.n440 B.n439 585
R683 B.n992 B.n991 585
R684 B.n993 B.n992 585
R685 B.n434 B.n433 585
R686 B.n435 B.n434 585
R687 B.n1002 B.n1001 585
R688 B.n1001 B.n1000 585
R689 B.n1003 B.n432 585
R690 B.n432 B.n431 585
R691 B.n1005 B.n1004 585
R692 B.n1006 B.n1005 585
R693 B.n2 B.n0 585
R694 B.n4 B.n2 585
R695 B.n3 B.n1 585
R696 B.n1169 B.n3 585
R697 B.n1167 B.n1166 585
R698 B.n1168 B.n1167 585
R699 B.n1165 B.n9 585
R700 B.n9 B.n8 585
R701 B.n1164 B.n1163 585
R702 B.n1163 B.n1162 585
R703 B.n11 B.n10 585
R704 B.n1161 B.n11 585
R705 B.n1159 B.n1158 585
R706 B.n1160 B.n1159 585
R707 B.n1157 B.n16 585
R708 B.n16 B.n15 585
R709 B.n1156 B.n1155 585
R710 B.n1155 B.n1154 585
R711 B.n18 B.n17 585
R712 B.n1153 B.n18 585
R713 B.n1151 B.n1150 585
R714 B.n1152 B.n1151 585
R715 B.n1149 B.n23 585
R716 B.n23 B.n22 585
R717 B.n1148 B.n1147 585
R718 B.n1147 B.n1146 585
R719 B.n25 B.n24 585
R720 B.n1145 B.n25 585
R721 B.n1143 B.n1142 585
R722 B.n1144 B.n1143 585
R723 B.n1141 B.n30 585
R724 B.n30 B.n29 585
R725 B.n1140 B.n1139 585
R726 B.n1139 B.n1138 585
R727 B.n32 B.n31 585
R728 B.n1137 B.n32 585
R729 B.n1135 B.n1134 585
R730 B.n1136 B.n1135 585
R731 B.n1133 B.n37 585
R732 B.n37 B.n36 585
R733 B.n1132 B.n1131 585
R734 B.n1131 B.n1130 585
R735 B.n39 B.n38 585
R736 B.n1129 B.n39 585
R737 B.n1127 B.n1126 585
R738 B.n1128 B.n1127 585
R739 B.n1125 B.n44 585
R740 B.n44 B.n43 585
R741 B.n1124 B.n1123 585
R742 B.n1123 B.n1122 585
R743 B.n46 B.n45 585
R744 B.n1121 B.n46 585
R745 B.n1119 B.n1118 585
R746 B.n1120 B.n1119 585
R747 B.n1117 B.n51 585
R748 B.n51 B.n50 585
R749 B.n1116 B.n1115 585
R750 B.n1115 B.n1114 585
R751 B.n53 B.n52 585
R752 B.n1113 B.n53 585
R753 B.n1111 B.n1110 585
R754 B.n1112 B.n1111 585
R755 B.n1109 B.n58 585
R756 B.n58 B.n57 585
R757 B.n1108 B.n1107 585
R758 B.n1107 B.n1106 585
R759 B.n60 B.n59 585
R760 B.n1105 B.n60 585
R761 B.n1103 B.n1102 585
R762 B.n1104 B.n1103 585
R763 B.n1101 B.n65 585
R764 B.n65 B.n64 585
R765 B.n1100 B.n1099 585
R766 B.n1099 B.n1098 585
R767 B.n67 B.n66 585
R768 B.n1097 B.n67 585
R769 B.n1095 B.n1094 585
R770 B.n1096 B.n1095 585
R771 B.n1093 B.n72 585
R772 B.n72 B.n71 585
R773 B.n1092 B.n1091 585
R774 B.n1091 B.n1090 585
R775 B.n74 B.n73 585
R776 B.n1089 B.n74 585
R777 B.n1087 B.n1086 585
R778 B.n1088 B.n1087 585
R779 B.n1085 B.n79 585
R780 B.n79 B.n78 585
R781 B.n1084 B.n1083 585
R782 B.n1083 B.n1082 585
R783 B.n81 B.n80 585
R784 B.n1081 B.n81 585
R785 B.n1079 B.n1078 585
R786 B.n1080 B.n1079 585
R787 B.n1077 B.n86 585
R788 B.n86 B.n85 585
R789 B.n1076 B.n1075 585
R790 B.n1075 B.n1074 585
R791 B.n1172 B.n1171 585
R792 B.n1171 B.n1170 585
R793 B.n868 B.n522 478.086
R794 B.n1075 B.n88 478.086
R795 B.n866 B.n524 478.086
R796 B.n1072 B.n89 478.086
R797 B.n734 B.t8 400.204
R798 B.n561 B.t19 400.204
R799 B.n161 B.t16 400.204
R800 B.n158 B.t12 400.204
R801 B.n1073 B.n156 256.663
R802 B.n1073 B.n155 256.663
R803 B.n1073 B.n154 256.663
R804 B.n1073 B.n153 256.663
R805 B.n1073 B.n152 256.663
R806 B.n1073 B.n151 256.663
R807 B.n1073 B.n150 256.663
R808 B.n1073 B.n149 256.663
R809 B.n1073 B.n148 256.663
R810 B.n1073 B.n147 256.663
R811 B.n1073 B.n146 256.663
R812 B.n1073 B.n145 256.663
R813 B.n1073 B.n144 256.663
R814 B.n1073 B.n143 256.663
R815 B.n1073 B.n142 256.663
R816 B.n1073 B.n141 256.663
R817 B.n1073 B.n140 256.663
R818 B.n1073 B.n139 256.663
R819 B.n1073 B.n138 256.663
R820 B.n1073 B.n137 256.663
R821 B.n1073 B.n136 256.663
R822 B.n1073 B.n135 256.663
R823 B.n1073 B.n134 256.663
R824 B.n1073 B.n133 256.663
R825 B.n1073 B.n132 256.663
R826 B.n1073 B.n131 256.663
R827 B.n1073 B.n130 256.663
R828 B.n1073 B.n129 256.663
R829 B.n1073 B.n128 256.663
R830 B.n1073 B.n127 256.663
R831 B.n1073 B.n126 256.663
R832 B.n1073 B.n125 256.663
R833 B.n1073 B.n124 256.663
R834 B.n1073 B.n123 256.663
R835 B.n1073 B.n122 256.663
R836 B.n1073 B.n121 256.663
R837 B.n1073 B.n120 256.663
R838 B.n1073 B.n119 256.663
R839 B.n1073 B.n118 256.663
R840 B.n1073 B.n117 256.663
R841 B.n1073 B.n116 256.663
R842 B.n1073 B.n115 256.663
R843 B.n1073 B.n114 256.663
R844 B.n1073 B.n113 256.663
R845 B.n1073 B.n112 256.663
R846 B.n1073 B.n111 256.663
R847 B.n1073 B.n110 256.663
R848 B.n1073 B.n109 256.663
R849 B.n1073 B.n108 256.663
R850 B.n1073 B.n107 256.663
R851 B.n1073 B.n106 256.663
R852 B.n1073 B.n105 256.663
R853 B.n1073 B.n104 256.663
R854 B.n1073 B.n103 256.663
R855 B.n1073 B.n102 256.663
R856 B.n1073 B.n101 256.663
R857 B.n1073 B.n100 256.663
R858 B.n1073 B.n99 256.663
R859 B.n1073 B.n98 256.663
R860 B.n1073 B.n97 256.663
R861 B.n1073 B.n96 256.663
R862 B.n1073 B.n95 256.663
R863 B.n1073 B.n94 256.663
R864 B.n1073 B.n93 256.663
R865 B.n1073 B.n92 256.663
R866 B.n1073 B.n91 256.663
R867 B.n1073 B.n90 256.663
R868 B.n593 B.n523 256.663
R869 B.n599 B.n523 256.663
R870 B.n601 B.n523 256.663
R871 B.n607 B.n523 256.663
R872 B.n609 B.n523 256.663
R873 B.n615 B.n523 256.663
R874 B.n617 B.n523 256.663
R875 B.n623 B.n523 256.663
R876 B.n625 B.n523 256.663
R877 B.n631 B.n523 256.663
R878 B.n633 B.n523 256.663
R879 B.n639 B.n523 256.663
R880 B.n641 B.n523 256.663
R881 B.n647 B.n523 256.663
R882 B.n649 B.n523 256.663
R883 B.n655 B.n523 256.663
R884 B.n657 B.n523 256.663
R885 B.n663 B.n523 256.663
R886 B.n665 B.n523 256.663
R887 B.n671 B.n523 256.663
R888 B.n673 B.n523 256.663
R889 B.n679 B.n523 256.663
R890 B.n681 B.n523 256.663
R891 B.n687 B.n523 256.663
R892 B.n689 B.n523 256.663
R893 B.n695 B.n523 256.663
R894 B.n697 B.n523 256.663
R895 B.n703 B.n523 256.663
R896 B.n705 B.n523 256.663
R897 B.n711 B.n523 256.663
R898 B.n713 B.n523 256.663
R899 B.n720 B.n523 256.663
R900 B.n722 B.n523 256.663
R901 B.n728 B.n523 256.663
R902 B.n730 B.n523 256.663
R903 B.n739 B.n523 256.663
R904 B.n741 B.n523 256.663
R905 B.n747 B.n523 256.663
R906 B.n749 B.n523 256.663
R907 B.n755 B.n523 256.663
R908 B.n757 B.n523 256.663
R909 B.n763 B.n523 256.663
R910 B.n765 B.n523 256.663
R911 B.n771 B.n523 256.663
R912 B.n773 B.n523 256.663
R913 B.n779 B.n523 256.663
R914 B.n781 B.n523 256.663
R915 B.n787 B.n523 256.663
R916 B.n789 B.n523 256.663
R917 B.n795 B.n523 256.663
R918 B.n797 B.n523 256.663
R919 B.n803 B.n523 256.663
R920 B.n805 B.n523 256.663
R921 B.n811 B.n523 256.663
R922 B.n813 B.n523 256.663
R923 B.n819 B.n523 256.663
R924 B.n821 B.n523 256.663
R925 B.n827 B.n523 256.663
R926 B.n829 B.n523 256.663
R927 B.n835 B.n523 256.663
R928 B.n837 B.n523 256.663
R929 B.n843 B.n523 256.663
R930 B.n845 B.n523 256.663
R931 B.n851 B.n523 256.663
R932 B.n853 B.n523 256.663
R933 B.n859 B.n523 256.663
R934 B.n861 B.n523 256.663
R935 B.n868 B.n520 163.367
R936 B.n872 B.n520 163.367
R937 B.n872 B.n514 163.367
R938 B.n880 B.n514 163.367
R939 B.n880 B.n512 163.367
R940 B.n884 B.n512 163.367
R941 B.n884 B.n506 163.367
R942 B.n892 B.n506 163.367
R943 B.n892 B.n504 163.367
R944 B.n896 B.n504 163.367
R945 B.n896 B.n498 163.367
R946 B.n904 B.n498 163.367
R947 B.n904 B.n496 163.367
R948 B.n908 B.n496 163.367
R949 B.n908 B.n490 163.367
R950 B.n916 B.n490 163.367
R951 B.n916 B.n488 163.367
R952 B.n920 B.n488 163.367
R953 B.n920 B.n482 163.367
R954 B.n928 B.n482 163.367
R955 B.n928 B.n480 163.367
R956 B.n932 B.n480 163.367
R957 B.n932 B.n474 163.367
R958 B.n940 B.n474 163.367
R959 B.n940 B.n472 163.367
R960 B.n944 B.n472 163.367
R961 B.n944 B.n466 163.367
R962 B.n952 B.n466 163.367
R963 B.n952 B.n464 163.367
R964 B.n956 B.n464 163.367
R965 B.n956 B.n458 163.367
R966 B.n964 B.n458 163.367
R967 B.n964 B.n456 163.367
R968 B.n968 B.n456 163.367
R969 B.n968 B.n450 163.367
R970 B.n976 B.n450 163.367
R971 B.n976 B.n448 163.367
R972 B.n980 B.n448 163.367
R973 B.n980 B.n442 163.367
R974 B.n988 B.n442 163.367
R975 B.n988 B.n440 163.367
R976 B.n992 B.n440 163.367
R977 B.n992 B.n434 163.367
R978 B.n1001 B.n434 163.367
R979 B.n1001 B.n432 163.367
R980 B.n1005 B.n432 163.367
R981 B.n1005 B.n2 163.367
R982 B.n1171 B.n2 163.367
R983 B.n1171 B.n3 163.367
R984 B.n1167 B.n3 163.367
R985 B.n1167 B.n9 163.367
R986 B.n1163 B.n9 163.367
R987 B.n1163 B.n11 163.367
R988 B.n1159 B.n11 163.367
R989 B.n1159 B.n16 163.367
R990 B.n1155 B.n16 163.367
R991 B.n1155 B.n18 163.367
R992 B.n1151 B.n18 163.367
R993 B.n1151 B.n23 163.367
R994 B.n1147 B.n23 163.367
R995 B.n1147 B.n25 163.367
R996 B.n1143 B.n25 163.367
R997 B.n1143 B.n30 163.367
R998 B.n1139 B.n30 163.367
R999 B.n1139 B.n32 163.367
R1000 B.n1135 B.n32 163.367
R1001 B.n1135 B.n37 163.367
R1002 B.n1131 B.n37 163.367
R1003 B.n1131 B.n39 163.367
R1004 B.n1127 B.n39 163.367
R1005 B.n1127 B.n44 163.367
R1006 B.n1123 B.n44 163.367
R1007 B.n1123 B.n46 163.367
R1008 B.n1119 B.n46 163.367
R1009 B.n1119 B.n51 163.367
R1010 B.n1115 B.n51 163.367
R1011 B.n1115 B.n53 163.367
R1012 B.n1111 B.n53 163.367
R1013 B.n1111 B.n58 163.367
R1014 B.n1107 B.n58 163.367
R1015 B.n1107 B.n60 163.367
R1016 B.n1103 B.n60 163.367
R1017 B.n1103 B.n65 163.367
R1018 B.n1099 B.n65 163.367
R1019 B.n1099 B.n67 163.367
R1020 B.n1095 B.n67 163.367
R1021 B.n1095 B.n72 163.367
R1022 B.n1091 B.n72 163.367
R1023 B.n1091 B.n74 163.367
R1024 B.n1087 B.n74 163.367
R1025 B.n1087 B.n79 163.367
R1026 B.n1083 B.n79 163.367
R1027 B.n1083 B.n81 163.367
R1028 B.n1079 B.n81 163.367
R1029 B.n1079 B.n86 163.367
R1030 B.n1075 B.n86 163.367
R1031 B.n594 B.n592 163.367
R1032 B.n598 B.n592 163.367
R1033 B.n602 B.n600 163.367
R1034 B.n606 B.n590 163.367
R1035 B.n610 B.n608 163.367
R1036 B.n614 B.n588 163.367
R1037 B.n618 B.n616 163.367
R1038 B.n622 B.n586 163.367
R1039 B.n626 B.n624 163.367
R1040 B.n630 B.n584 163.367
R1041 B.n634 B.n632 163.367
R1042 B.n638 B.n582 163.367
R1043 B.n642 B.n640 163.367
R1044 B.n646 B.n580 163.367
R1045 B.n650 B.n648 163.367
R1046 B.n654 B.n578 163.367
R1047 B.n658 B.n656 163.367
R1048 B.n662 B.n576 163.367
R1049 B.n666 B.n664 163.367
R1050 B.n670 B.n574 163.367
R1051 B.n674 B.n672 163.367
R1052 B.n678 B.n572 163.367
R1053 B.n682 B.n680 163.367
R1054 B.n686 B.n570 163.367
R1055 B.n690 B.n688 163.367
R1056 B.n694 B.n568 163.367
R1057 B.n698 B.n696 163.367
R1058 B.n702 B.n566 163.367
R1059 B.n706 B.n704 163.367
R1060 B.n710 B.n564 163.367
R1061 B.n714 B.n712 163.367
R1062 B.n719 B.n560 163.367
R1063 B.n723 B.n721 163.367
R1064 B.n727 B.n558 163.367
R1065 B.n731 B.n729 163.367
R1066 B.n738 B.n556 163.367
R1067 B.n742 B.n740 163.367
R1068 B.n746 B.n554 163.367
R1069 B.n750 B.n748 163.367
R1070 B.n754 B.n552 163.367
R1071 B.n758 B.n756 163.367
R1072 B.n762 B.n550 163.367
R1073 B.n766 B.n764 163.367
R1074 B.n770 B.n548 163.367
R1075 B.n774 B.n772 163.367
R1076 B.n778 B.n546 163.367
R1077 B.n782 B.n780 163.367
R1078 B.n786 B.n544 163.367
R1079 B.n790 B.n788 163.367
R1080 B.n794 B.n542 163.367
R1081 B.n798 B.n796 163.367
R1082 B.n802 B.n540 163.367
R1083 B.n806 B.n804 163.367
R1084 B.n810 B.n538 163.367
R1085 B.n814 B.n812 163.367
R1086 B.n818 B.n536 163.367
R1087 B.n822 B.n820 163.367
R1088 B.n826 B.n534 163.367
R1089 B.n830 B.n828 163.367
R1090 B.n834 B.n532 163.367
R1091 B.n838 B.n836 163.367
R1092 B.n842 B.n530 163.367
R1093 B.n846 B.n844 163.367
R1094 B.n850 B.n528 163.367
R1095 B.n854 B.n852 163.367
R1096 B.n858 B.n526 163.367
R1097 B.n862 B.n860 163.367
R1098 B.n866 B.n518 163.367
R1099 B.n874 B.n518 163.367
R1100 B.n874 B.n516 163.367
R1101 B.n878 B.n516 163.367
R1102 B.n878 B.n509 163.367
R1103 B.n886 B.n509 163.367
R1104 B.n886 B.n507 163.367
R1105 B.n890 B.n507 163.367
R1106 B.n890 B.n502 163.367
R1107 B.n898 B.n502 163.367
R1108 B.n898 B.n500 163.367
R1109 B.n902 B.n500 163.367
R1110 B.n902 B.n494 163.367
R1111 B.n910 B.n494 163.367
R1112 B.n910 B.n492 163.367
R1113 B.n914 B.n492 163.367
R1114 B.n914 B.n486 163.367
R1115 B.n922 B.n486 163.367
R1116 B.n922 B.n484 163.367
R1117 B.n926 B.n484 163.367
R1118 B.n926 B.n478 163.367
R1119 B.n934 B.n478 163.367
R1120 B.n934 B.n476 163.367
R1121 B.n938 B.n476 163.367
R1122 B.n938 B.n470 163.367
R1123 B.n946 B.n470 163.367
R1124 B.n946 B.n468 163.367
R1125 B.n950 B.n468 163.367
R1126 B.n950 B.n462 163.367
R1127 B.n958 B.n462 163.367
R1128 B.n958 B.n460 163.367
R1129 B.n962 B.n460 163.367
R1130 B.n962 B.n454 163.367
R1131 B.n970 B.n454 163.367
R1132 B.n970 B.n452 163.367
R1133 B.n974 B.n452 163.367
R1134 B.n974 B.n446 163.367
R1135 B.n982 B.n446 163.367
R1136 B.n982 B.n444 163.367
R1137 B.n986 B.n444 163.367
R1138 B.n986 B.n438 163.367
R1139 B.n994 B.n438 163.367
R1140 B.n994 B.n436 163.367
R1141 B.n999 B.n436 163.367
R1142 B.n999 B.n430 163.367
R1143 B.n1007 B.n430 163.367
R1144 B.n1008 B.n1007 163.367
R1145 B.n1008 B.n5 163.367
R1146 B.n6 B.n5 163.367
R1147 B.n7 B.n6 163.367
R1148 B.n1013 B.n7 163.367
R1149 B.n1013 B.n12 163.367
R1150 B.n13 B.n12 163.367
R1151 B.n14 B.n13 163.367
R1152 B.n1018 B.n14 163.367
R1153 B.n1018 B.n19 163.367
R1154 B.n20 B.n19 163.367
R1155 B.n21 B.n20 163.367
R1156 B.n1023 B.n21 163.367
R1157 B.n1023 B.n26 163.367
R1158 B.n27 B.n26 163.367
R1159 B.n28 B.n27 163.367
R1160 B.n1028 B.n28 163.367
R1161 B.n1028 B.n33 163.367
R1162 B.n34 B.n33 163.367
R1163 B.n35 B.n34 163.367
R1164 B.n1033 B.n35 163.367
R1165 B.n1033 B.n40 163.367
R1166 B.n41 B.n40 163.367
R1167 B.n42 B.n41 163.367
R1168 B.n1038 B.n42 163.367
R1169 B.n1038 B.n47 163.367
R1170 B.n48 B.n47 163.367
R1171 B.n49 B.n48 163.367
R1172 B.n1043 B.n49 163.367
R1173 B.n1043 B.n54 163.367
R1174 B.n55 B.n54 163.367
R1175 B.n56 B.n55 163.367
R1176 B.n1048 B.n56 163.367
R1177 B.n1048 B.n61 163.367
R1178 B.n62 B.n61 163.367
R1179 B.n63 B.n62 163.367
R1180 B.n1053 B.n63 163.367
R1181 B.n1053 B.n68 163.367
R1182 B.n69 B.n68 163.367
R1183 B.n70 B.n69 163.367
R1184 B.n1058 B.n70 163.367
R1185 B.n1058 B.n75 163.367
R1186 B.n76 B.n75 163.367
R1187 B.n77 B.n76 163.367
R1188 B.n1063 B.n77 163.367
R1189 B.n1063 B.n82 163.367
R1190 B.n83 B.n82 163.367
R1191 B.n84 B.n83 163.367
R1192 B.n1068 B.n84 163.367
R1193 B.n1068 B.n89 163.367
R1194 B.n165 B.n164 163.367
R1195 B.n169 B.n168 163.367
R1196 B.n173 B.n172 163.367
R1197 B.n177 B.n176 163.367
R1198 B.n181 B.n180 163.367
R1199 B.n185 B.n184 163.367
R1200 B.n189 B.n188 163.367
R1201 B.n193 B.n192 163.367
R1202 B.n197 B.n196 163.367
R1203 B.n201 B.n200 163.367
R1204 B.n205 B.n204 163.367
R1205 B.n209 B.n208 163.367
R1206 B.n213 B.n212 163.367
R1207 B.n217 B.n216 163.367
R1208 B.n221 B.n220 163.367
R1209 B.n225 B.n224 163.367
R1210 B.n229 B.n228 163.367
R1211 B.n233 B.n232 163.367
R1212 B.n237 B.n236 163.367
R1213 B.n241 B.n240 163.367
R1214 B.n245 B.n244 163.367
R1215 B.n249 B.n248 163.367
R1216 B.n253 B.n252 163.367
R1217 B.n257 B.n256 163.367
R1218 B.n261 B.n260 163.367
R1219 B.n265 B.n264 163.367
R1220 B.n269 B.n268 163.367
R1221 B.n273 B.n272 163.367
R1222 B.n277 B.n276 163.367
R1223 B.n281 B.n280 163.367
R1224 B.n285 B.n284 163.367
R1225 B.n290 B.n289 163.367
R1226 B.n294 B.n293 163.367
R1227 B.n298 B.n297 163.367
R1228 B.n302 B.n301 163.367
R1229 B.n306 B.n305 163.367
R1230 B.n310 B.n309 163.367
R1231 B.n314 B.n313 163.367
R1232 B.n318 B.n317 163.367
R1233 B.n322 B.n321 163.367
R1234 B.n326 B.n325 163.367
R1235 B.n330 B.n329 163.367
R1236 B.n334 B.n333 163.367
R1237 B.n338 B.n337 163.367
R1238 B.n342 B.n341 163.367
R1239 B.n346 B.n345 163.367
R1240 B.n350 B.n349 163.367
R1241 B.n354 B.n353 163.367
R1242 B.n358 B.n357 163.367
R1243 B.n362 B.n361 163.367
R1244 B.n366 B.n365 163.367
R1245 B.n370 B.n369 163.367
R1246 B.n374 B.n373 163.367
R1247 B.n378 B.n377 163.367
R1248 B.n382 B.n381 163.367
R1249 B.n386 B.n385 163.367
R1250 B.n390 B.n389 163.367
R1251 B.n394 B.n393 163.367
R1252 B.n398 B.n397 163.367
R1253 B.n402 B.n401 163.367
R1254 B.n406 B.n405 163.367
R1255 B.n410 B.n409 163.367
R1256 B.n414 B.n413 163.367
R1257 B.n418 B.n417 163.367
R1258 B.n422 B.n421 163.367
R1259 B.n426 B.n425 163.367
R1260 B.n1072 B.n157 163.367
R1261 B.n734 B.t11 120.909
R1262 B.n158 B.t14 120.909
R1263 B.n561 B.t21 120.883
R1264 B.n161 B.t17 120.883
R1265 B.n593 B.n522 71.676
R1266 B.n599 B.n598 71.676
R1267 B.n602 B.n601 71.676
R1268 B.n607 B.n606 71.676
R1269 B.n610 B.n609 71.676
R1270 B.n615 B.n614 71.676
R1271 B.n618 B.n617 71.676
R1272 B.n623 B.n622 71.676
R1273 B.n626 B.n625 71.676
R1274 B.n631 B.n630 71.676
R1275 B.n634 B.n633 71.676
R1276 B.n639 B.n638 71.676
R1277 B.n642 B.n641 71.676
R1278 B.n647 B.n646 71.676
R1279 B.n650 B.n649 71.676
R1280 B.n655 B.n654 71.676
R1281 B.n658 B.n657 71.676
R1282 B.n663 B.n662 71.676
R1283 B.n666 B.n665 71.676
R1284 B.n671 B.n670 71.676
R1285 B.n674 B.n673 71.676
R1286 B.n679 B.n678 71.676
R1287 B.n682 B.n681 71.676
R1288 B.n687 B.n686 71.676
R1289 B.n690 B.n689 71.676
R1290 B.n695 B.n694 71.676
R1291 B.n698 B.n697 71.676
R1292 B.n703 B.n702 71.676
R1293 B.n706 B.n705 71.676
R1294 B.n711 B.n710 71.676
R1295 B.n714 B.n713 71.676
R1296 B.n720 B.n719 71.676
R1297 B.n723 B.n722 71.676
R1298 B.n728 B.n727 71.676
R1299 B.n731 B.n730 71.676
R1300 B.n739 B.n738 71.676
R1301 B.n742 B.n741 71.676
R1302 B.n747 B.n746 71.676
R1303 B.n750 B.n749 71.676
R1304 B.n755 B.n754 71.676
R1305 B.n758 B.n757 71.676
R1306 B.n763 B.n762 71.676
R1307 B.n766 B.n765 71.676
R1308 B.n771 B.n770 71.676
R1309 B.n774 B.n773 71.676
R1310 B.n779 B.n778 71.676
R1311 B.n782 B.n781 71.676
R1312 B.n787 B.n786 71.676
R1313 B.n790 B.n789 71.676
R1314 B.n795 B.n794 71.676
R1315 B.n798 B.n797 71.676
R1316 B.n803 B.n802 71.676
R1317 B.n806 B.n805 71.676
R1318 B.n811 B.n810 71.676
R1319 B.n814 B.n813 71.676
R1320 B.n819 B.n818 71.676
R1321 B.n822 B.n821 71.676
R1322 B.n827 B.n826 71.676
R1323 B.n830 B.n829 71.676
R1324 B.n835 B.n834 71.676
R1325 B.n838 B.n837 71.676
R1326 B.n843 B.n842 71.676
R1327 B.n846 B.n845 71.676
R1328 B.n851 B.n850 71.676
R1329 B.n854 B.n853 71.676
R1330 B.n859 B.n858 71.676
R1331 B.n862 B.n861 71.676
R1332 B.n90 B.n88 71.676
R1333 B.n165 B.n91 71.676
R1334 B.n169 B.n92 71.676
R1335 B.n173 B.n93 71.676
R1336 B.n177 B.n94 71.676
R1337 B.n181 B.n95 71.676
R1338 B.n185 B.n96 71.676
R1339 B.n189 B.n97 71.676
R1340 B.n193 B.n98 71.676
R1341 B.n197 B.n99 71.676
R1342 B.n201 B.n100 71.676
R1343 B.n205 B.n101 71.676
R1344 B.n209 B.n102 71.676
R1345 B.n213 B.n103 71.676
R1346 B.n217 B.n104 71.676
R1347 B.n221 B.n105 71.676
R1348 B.n225 B.n106 71.676
R1349 B.n229 B.n107 71.676
R1350 B.n233 B.n108 71.676
R1351 B.n237 B.n109 71.676
R1352 B.n241 B.n110 71.676
R1353 B.n245 B.n111 71.676
R1354 B.n249 B.n112 71.676
R1355 B.n253 B.n113 71.676
R1356 B.n257 B.n114 71.676
R1357 B.n261 B.n115 71.676
R1358 B.n265 B.n116 71.676
R1359 B.n269 B.n117 71.676
R1360 B.n273 B.n118 71.676
R1361 B.n277 B.n119 71.676
R1362 B.n281 B.n120 71.676
R1363 B.n285 B.n121 71.676
R1364 B.n290 B.n122 71.676
R1365 B.n294 B.n123 71.676
R1366 B.n298 B.n124 71.676
R1367 B.n302 B.n125 71.676
R1368 B.n306 B.n126 71.676
R1369 B.n310 B.n127 71.676
R1370 B.n314 B.n128 71.676
R1371 B.n318 B.n129 71.676
R1372 B.n322 B.n130 71.676
R1373 B.n326 B.n131 71.676
R1374 B.n330 B.n132 71.676
R1375 B.n334 B.n133 71.676
R1376 B.n338 B.n134 71.676
R1377 B.n342 B.n135 71.676
R1378 B.n346 B.n136 71.676
R1379 B.n350 B.n137 71.676
R1380 B.n354 B.n138 71.676
R1381 B.n358 B.n139 71.676
R1382 B.n362 B.n140 71.676
R1383 B.n366 B.n141 71.676
R1384 B.n370 B.n142 71.676
R1385 B.n374 B.n143 71.676
R1386 B.n378 B.n144 71.676
R1387 B.n382 B.n145 71.676
R1388 B.n386 B.n146 71.676
R1389 B.n390 B.n147 71.676
R1390 B.n394 B.n148 71.676
R1391 B.n398 B.n149 71.676
R1392 B.n402 B.n150 71.676
R1393 B.n406 B.n151 71.676
R1394 B.n410 B.n152 71.676
R1395 B.n414 B.n153 71.676
R1396 B.n418 B.n154 71.676
R1397 B.n422 B.n155 71.676
R1398 B.n426 B.n156 71.676
R1399 B.n157 B.n156 71.676
R1400 B.n425 B.n155 71.676
R1401 B.n421 B.n154 71.676
R1402 B.n417 B.n153 71.676
R1403 B.n413 B.n152 71.676
R1404 B.n409 B.n151 71.676
R1405 B.n405 B.n150 71.676
R1406 B.n401 B.n149 71.676
R1407 B.n397 B.n148 71.676
R1408 B.n393 B.n147 71.676
R1409 B.n389 B.n146 71.676
R1410 B.n385 B.n145 71.676
R1411 B.n381 B.n144 71.676
R1412 B.n377 B.n143 71.676
R1413 B.n373 B.n142 71.676
R1414 B.n369 B.n141 71.676
R1415 B.n365 B.n140 71.676
R1416 B.n361 B.n139 71.676
R1417 B.n357 B.n138 71.676
R1418 B.n353 B.n137 71.676
R1419 B.n349 B.n136 71.676
R1420 B.n345 B.n135 71.676
R1421 B.n341 B.n134 71.676
R1422 B.n337 B.n133 71.676
R1423 B.n333 B.n132 71.676
R1424 B.n329 B.n131 71.676
R1425 B.n325 B.n130 71.676
R1426 B.n321 B.n129 71.676
R1427 B.n317 B.n128 71.676
R1428 B.n313 B.n127 71.676
R1429 B.n309 B.n126 71.676
R1430 B.n305 B.n125 71.676
R1431 B.n301 B.n124 71.676
R1432 B.n297 B.n123 71.676
R1433 B.n293 B.n122 71.676
R1434 B.n289 B.n121 71.676
R1435 B.n284 B.n120 71.676
R1436 B.n280 B.n119 71.676
R1437 B.n276 B.n118 71.676
R1438 B.n272 B.n117 71.676
R1439 B.n268 B.n116 71.676
R1440 B.n264 B.n115 71.676
R1441 B.n260 B.n114 71.676
R1442 B.n256 B.n113 71.676
R1443 B.n252 B.n112 71.676
R1444 B.n248 B.n111 71.676
R1445 B.n244 B.n110 71.676
R1446 B.n240 B.n109 71.676
R1447 B.n236 B.n108 71.676
R1448 B.n232 B.n107 71.676
R1449 B.n228 B.n106 71.676
R1450 B.n224 B.n105 71.676
R1451 B.n220 B.n104 71.676
R1452 B.n216 B.n103 71.676
R1453 B.n212 B.n102 71.676
R1454 B.n208 B.n101 71.676
R1455 B.n204 B.n100 71.676
R1456 B.n200 B.n99 71.676
R1457 B.n196 B.n98 71.676
R1458 B.n192 B.n97 71.676
R1459 B.n188 B.n96 71.676
R1460 B.n184 B.n95 71.676
R1461 B.n180 B.n94 71.676
R1462 B.n176 B.n93 71.676
R1463 B.n172 B.n92 71.676
R1464 B.n168 B.n91 71.676
R1465 B.n164 B.n90 71.676
R1466 B.n594 B.n593 71.676
R1467 B.n600 B.n599 71.676
R1468 B.n601 B.n590 71.676
R1469 B.n608 B.n607 71.676
R1470 B.n609 B.n588 71.676
R1471 B.n616 B.n615 71.676
R1472 B.n617 B.n586 71.676
R1473 B.n624 B.n623 71.676
R1474 B.n625 B.n584 71.676
R1475 B.n632 B.n631 71.676
R1476 B.n633 B.n582 71.676
R1477 B.n640 B.n639 71.676
R1478 B.n641 B.n580 71.676
R1479 B.n648 B.n647 71.676
R1480 B.n649 B.n578 71.676
R1481 B.n656 B.n655 71.676
R1482 B.n657 B.n576 71.676
R1483 B.n664 B.n663 71.676
R1484 B.n665 B.n574 71.676
R1485 B.n672 B.n671 71.676
R1486 B.n673 B.n572 71.676
R1487 B.n680 B.n679 71.676
R1488 B.n681 B.n570 71.676
R1489 B.n688 B.n687 71.676
R1490 B.n689 B.n568 71.676
R1491 B.n696 B.n695 71.676
R1492 B.n697 B.n566 71.676
R1493 B.n704 B.n703 71.676
R1494 B.n705 B.n564 71.676
R1495 B.n712 B.n711 71.676
R1496 B.n713 B.n560 71.676
R1497 B.n721 B.n720 71.676
R1498 B.n722 B.n558 71.676
R1499 B.n729 B.n728 71.676
R1500 B.n730 B.n556 71.676
R1501 B.n740 B.n739 71.676
R1502 B.n741 B.n554 71.676
R1503 B.n748 B.n747 71.676
R1504 B.n749 B.n552 71.676
R1505 B.n756 B.n755 71.676
R1506 B.n757 B.n550 71.676
R1507 B.n764 B.n763 71.676
R1508 B.n765 B.n548 71.676
R1509 B.n772 B.n771 71.676
R1510 B.n773 B.n546 71.676
R1511 B.n780 B.n779 71.676
R1512 B.n781 B.n544 71.676
R1513 B.n788 B.n787 71.676
R1514 B.n789 B.n542 71.676
R1515 B.n796 B.n795 71.676
R1516 B.n797 B.n540 71.676
R1517 B.n804 B.n803 71.676
R1518 B.n805 B.n538 71.676
R1519 B.n812 B.n811 71.676
R1520 B.n813 B.n536 71.676
R1521 B.n820 B.n819 71.676
R1522 B.n821 B.n534 71.676
R1523 B.n828 B.n827 71.676
R1524 B.n829 B.n532 71.676
R1525 B.n836 B.n835 71.676
R1526 B.n837 B.n530 71.676
R1527 B.n844 B.n843 71.676
R1528 B.n845 B.n528 71.676
R1529 B.n852 B.n851 71.676
R1530 B.n853 B.n526 71.676
R1531 B.n860 B.n859 71.676
R1532 B.n861 B.n524 71.676
R1533 B.n735 B.t10 68.1573
R1534 B.n159 B.t15 68.1573
R1535 B.n562 B.t20 68.1316
R1536 B.n162 B.t18 68.1316
R1537 B.n736 B.n735 59.5399
R1538 B.n717 B.n562 59.5399
R1539 B.n287 B.n162 59.5399
R1540 B.n160 B.n159 59.5399
R1541 B.n867 B.n523 59.1427
R1542 B.n1074 B.n1073 59.1427
R1543 B.n735 B.n734 52.752
R1544 B.n562 B.n561 52.752
R1545 B.n162 B.n161 52.752
R1546 B.n159 B.n158 52.752
R1547 B.n1076 B.n87 31.0639
R1548 B.n1071 B.n1070 31.0639
R1549 B.n865 B.n864 31.0639
R1550 B.n869 B.n521 31.0639
R1551 B.n867 B.n519 30.7003
R1552 B.n873 B.n519 30.7003
R1553 B.n873 B.n515 30.7003
R1554 B.n879 B.n515 30.7003
R1555 B.n879 B.n510 30.7003
R1556 B.n885 B.n510 30.7003
R1557 B.n885 B.n511 30.7003
R1558 B.n891 B.n503 30.7003
R1559 B.n897 B.n503 30.7003
R1560 B.n897 B.n499 30.7003
R1561 B.n903 B.n499 30.7003
R1562 B.n903 B.n495 30.7003
R1563 B.n909 B.n495 30.7003
R1564 B.n909 B.n491 30.7003
R1565 B.n915 B.n491 30.7003
R1566 B.n915 B.n487 30.7003
R1567 B.n921 B.n487 30.7003
R1568 B.n927 B.n483 30.7003
R1569 B.n927 B.n479 30.7003
R1570 B.n933 B.n479 30.7003
R1571 B.n933 B.n475 30.7003
R1572 B.n939 B.n475 30.7003
R1573 B.n939 B.n471 30.7003
R1574 B.n945 B.n471 30.7003
R1575 B.n951 B.n467 30.7003
R1576 B.n951 B.n463 30.7003
R1577 B.n957 B.n463 30.7003
R1578 B.n957 B.n459 30.7003
R1579 B.n963 B.n459 30.7003
R1580 B.n963 B.n455 30.7003
R1581 B.n969 B.n455 30.7003
R1582 B.n975 B.n451 30.7003
R1583 B.n975 B.n447 30.7003
R1584 B.n981 B.n447 30.7003
R1585 B.n981 B.n443 30.7003
R1586 B.n987 B.n443 30.7003
R1587 B.n987 B.n439 30.7003
R1588 B.n993 B.n439 30.7003
R1589 B.n1000 B.n435 30.7003
R1590 B.n1000 B.n431 30.7003
R1591 B.n1006 B.n431 30.7003
R1592 B.n1006 B.n4 30.7003
R1593 B.n1170 B.n4 30.7003
R1594 B.n1170 B.n1169 30.7003
R1595 B.n1169 B.n1168 30.7003
R1596 B.n1168 B.n8 30.7003
R1597 B.n1162 B.n8 30.7003
R1598 B.n1162 B.n1161 30.7003
R1599 B.n1160 B.n15 30.7003
R1600 B.n1154 B.n15 30.7003
R1601 B.n1154 B.n1153 30.7003
R1602 B.n1153 B.n1152 30.7003
R1603 B.n1152 B.n22 30.7003
R1604 B.n1146 B.n22 30.7003
R1605 B.n1146 B.n1145 30.7003
R1606 B.n1144 B.n29 30.7003
R1607 B.n1138 B.n29 30.7003
R1608 B.n1138 B.n1137 30.7003
R1609 B.n1137 B.n1136 30.7003
R1610 B.n1136 B.n36 30.7003
R1611 B.n1130 B.n36 30.7003
R1612 B.n1130 B.n1129 30.7003
R1613 B.n1128 B.n43 30.7003
R1614 B.n1122 B.n43 30.7003
R1615 B.n1122 B.n1121 30.7003
R1616 B.n1121 B.n1120 30.7003
R1617 B.n1120 B.n50 30.7003
R1618 B.n1114 B.n50 30.7003
R1619 B.n1114 B.n1113 30.7003
R1620 B.n1112 B.n57 30.7003
R1621 B.n1106 B.n57 30.7003
R1622 B.n1106 B.n1105 30.7003
R1623 B.n1105 B.n1104 30.7003
R1624 B.n1104 B.n64 30.7003
R1625 B.n1098 B.n64 30.7003
R1626 B.n1098 B.n1097 30.7003
R1627 B.n1097 B.n1096 30.7003
R1628 B.n1096 B.n71 30.7003
R1629 B.n1090 B.n71 30.7003
R1630 B.n1089 B.n1088 30.7003
R1631 B.n1088 B.n78 30.7003
R1632 B.n1082 B.n78 30.7003
R1633 B.n1082 B.n1081 30.7003
R1634 B.n1081 B.n1080 30.7003
R1635 B.n1080 B.n85 30.7003
R1636 B.n1074 B.n85 30.7003
R1637 B.n891 B.t9 24.8312
R1638 B.n1090 B.t13 24.8312
R1639 B.t5 B.n483 18.5107
R1640 B.t0 B.n467 18.5107
R1641 B.t4 B.n451 18.5107
R1642 B.t2 B.n435 18.5107
R1643 B.n1161 B.t7 18.5107
R1644 B.n1145 B.t6 18.5107
R1645 B.n1129 B.t3 18.5107
R1646 B.n1113 B.t1 18.5107
R1647 B B.n1172 18.0485
R1648 B.n921 B.t5 12.1901
R1649 B.n945 B.t0 12.1901
R1650 B.n969 B.t4 12.1901
R1651 B.n993 B.t2 12.1901
R1652 B.t7 B.n1160 12.1901
R1653 B.t6 B.n1144 12.1901
R1654 B.t3 B.n1128 12.1901
R1655 B.t1 B.n1112 12.1901
R1656 B.n163 B.n87 10.6151
R1657 B.n166 B.n163 10.6151
R1658 B.n167 B.n166 10.6151
R1659 B.n170 B.n167 10.6151
R1660 B.n171 B.n170 10.6151
R1661 B.n174 B.n171 10.6151
R1662 B.n175 B.n174 10.6151
R1663 B.n178 B.n175 10.6151
R1664 B.n179 B.n178 10.6151
R1665 B.n182 B.n179 10.6151
R1666 B.n183 B.n182 10.6151
R1667 B.n186 B.n183 10.6151
R1668 B.n187 B.n186 10.6151
R1669 B.n190 B.n187 10.6151
R1670 B.n191 B.n190 10.6151
R1671 B.n194 B.n191 10.6151
R1672 B.n195 B.n194 10.6151
R1673 B.n198 B.n195 10.6151
R1674 B.n199 B.n198 10.6151
R1675 B.n202 B.n199 10.6151
R1676 B.n203 B.n202 10.6151
R1677 B.n206 B.n203 10.6151
R1678 B.n207 B.n206 10.6151
R1679 B.n210 B.n207 10.6151
R1680 B.n211 B.n210 10.6151
R1681 B.n214 B.n211 10.6151
R1682 B.n215 B.n214 10.6151
R1683 B.n218 B.n215 10.6151
R1684 B.n219 B.n218 10.6151
R1685 B.n222 B.n219 10.6151
R1686 B.n223 B.n222 10.6151
R1687 B.n226 B.n223 10.6151
R1688 B.n227 B.n226 10.6151
R1689 B.n230 B.n227 10.6151
R1690 B.n231 B.n230 10.6151
R1691 B.n234 B.n231 10.6151
R1692 B.n235 B.n234 10.6151
R1693 B.n238 B.n235 10.6151
R1694 B.n239 B.n238 10.6151
R1695 B.n242 B.n239 10.6151
R1696 B.n243 B.n242 10.6151
R1697 B.n246 B.n243 10.6151
R1698 B.n247 B.n246 10.6151
R1699 B.n250 B.n247 10.6151
R1700 B.n251 B.n250 10.6151
R1701 B.n254 B.n251 10.6151
R1702 B.n255 B.n254 10.6151
R1703 B.n258 B.n255 10.6151
R1704 B.n259 B.n258 10.6151
R1705 B.n262 B.n259 10.6151
R1706 B.n263 B.n262 10.6151
R1707 B.n266 B.n263 10.6151
R1708 B.n267 B.n266 10.6151
R1709 B.n270 B.n267 10.6151
R1710 B.n271 B.n270 10.6151
R1711 B.n274 B.n271 10.6151
R1712 B.n275 B.n274 10.6151
R1713 B.n278 B.n275 10.6151
R1714 B.n279 B.n278 10.6151
R1715 B.n282 B.n279 10.6151
R1716 B.n283 B.n282 10.6151
R1717 B.n286 B.n283 10.6151
R1718 B.n291 B.n288 10.6151
R1719 B.n292 B.n291 10.6151
R1720 B.n295 B.n292 10.6151
R1721 B.n296 B.n295 10.6151
R1722 B.n299 B.n296 10.6151
R1723 B.n300 B.n299 10.6151
R1724 B.n303 B.n300 10.6151
R1725 B.n304 B.n303 10.6151
R1726 B.n308 B.n307 10.6151
R1727 B.n311 B.n308 10.6151
R1728 B.n312 B.n311 10.6151
R1729 B.n315 B.n312 10.6151
R1730 B.n316 B.n315 10.6151
R1731 B.n319 B.n316 10.6151
R1732 B.n320 B.n319 10.6151
R1733 B.n323 B.n320 10.6151
R1734 B.n324 B.n323 10.6151
R1735 B.n327 B.n324 10.6151
R1736 B.n328 B.n327 10.6151
R1737 B.n331 B.n328 10.6151
R1738 B.n332 B.n331 10.6151
R1739 B.n335 B.n332 10.6151
R1740 B.n336 B.n335 10.6151
R1741 B.n339 B.n336 10.6151
R1742 B.n340 B.n339 10.6151
R1743 B.n343 B.n340 10.6151
R1744 B.n344 B.n343 10.6151
R1745 B.n347 B.n344 10.6151
R1746 B.n348 B.n347 10.6151
R1747 B.n351 B.n348 10.6151
R1748 B.n352 B.n351 10.6151
R1749 B.n355 B.n352 10.6151
R1750 B.n356 B.n355 10.6151
R1751 B.n359 B.n356 10.6151
R1752 B.n360 B.n359 10.6151
R1753 B.n363 B.n360 10.6151
R1754 B.n364 B.n363 10.6151
R1755 B.n367 B.n364 10.6151
R1756 B.n368 B.n367 10.6151
R1757 B.n371 B.n368 10.6151
R1758 B.n372 B.n371 10.6151
R1759 B.n375 B.n372 10.6151
R1760 B.n376 B.n375 10.6151
R1761 B.n379 B.n376 10.6151
R1762 B.n380 B.n379 10.6151
R1763 B.n383 B.n380 10.6151
R1764 B.n384 B.n383 10.6151
R1765 B.n387 B.n384 10.6151
R1766 B.n388 B.n387 10.6151
R1767 B.n391 B.n388 10.6151
R1768 B.n392 B.n391 10.6151
R1769 B.n395 B.n392 10.6151
R1770 B.n396 B.n395 10.6151
R1771 B.n399 B.n396 10.6151
R1772 B.n400 B.n399 10.6151
R1773 B.n403 B.n400 10.6151
R1774 B.n404 B.n403 10.6151
R1775 B.n407 B.n404 10.6151
R1776 B.n408 B.n407 10.6151
R1777 B.n411 B.n408 10.6151
R1778 B.n412 B.n411 10.6151
R1779 B.n415 B.n412 10.6151
R1780 B.n416 B.n415 10.6151
R1781 B.n419 B.n416 10.6151
R1782 B.n420 B.n419 10.6151
R1783 B.n423 B.n420 10.6151
R1784 B.n424 B.n423 10.6151
R1785 B.n427 B.n424 10.6151
R1786 B.n428 B.n427 10.6151
R1787 B.n1071 B.n428 10.6151
R1788 B.n865 B.n517 10.6151
R1789 B.n875 B.n517 10.6151
R1790 B.n876 B.n875 10.6151
R1791 B.n877 B.n876 10.6151
R1792 B.n877 B.n508 10.6151
R1793 B.n887 B.n508 10.6151
R1794 B.n888 B.n887 10.6151
R1795 B.n889 B.n888 10.6151
R1796 B.n889 B.n501 10.6151
R1797 B.n899 B.n501 10.6151
R1798 B.n900 B.n899 10.6151
R1799 B.n901 B.n900 10.6151
R1800 B.n901 B.n493 10.6151
R1801 B.n911 B.n493 10.6151
R1802 B.n912 B.n911 10.6151
R1803 B.n913 B.n912 10.6151
R1804 B.n913 B.n485 10.6151
R1805 B.n923 B.n485 10.6151
R1806 B.n924 B.n923 10.6151
R1807 B.n925 B.n924 10.6151
R1808 B.n925 B.n477 10.6151
R1809 B.n935 B.n477 10.6151
R1810 B.n936 B.n935 10.6151
R1811 B.n937 B.n936 10.6151
R1812 B.n937 B.n469 10.6151
R1813 B.n947 B.n469 10.6151
R1814 B.n948 B.n947 10.6151
R1815 B.n949 B.n948 10.6151
R1816 B.n949 B.n461 10.6151
R1817 B.n959 B.n461 10.6151
R1818 B.n960 B.n959 10.6151
R1819 B.n961 B.n960 10.6151
R1820 B.n961 B.n453 10.6151
R1821 B.n971 B.n453 10.6151
R1822 B.n972 B.n971 10.6151
R1823 B.n973 B.n972 10.6151
R1824 B.n973 B.n445 10.6151
R1825 B.n983 B.n445 10.6151
R1826 B.n984 B.n983 10.6151
R1827 B.n985 B.n984 10.6151
R1828 B.n985 B.n437 10.6151
R1829 B.n995 B.n437 10.6151
R1830 B.n996 B.n995 10.6151
R1831 B.n998 B.n996 10.6151
R1832 B.n998 B.n997 10.6151
R1833 B.n997 B.n429 10.6151
R1834 B.n1009 B.n429 10.6151
R1835 B.n1010 B.n1009 10.6151
R1836 B.n1011 B.n1010 10.6151
R1837 B.n1012 B.n1011 10.6151
R1838 B.n1014 B.n1012 10.6151
R1839 B.n1015 B.n1014 10.6151
R1840 B.n1016 B.n1015 10.6151
R1841 B.n1017 B.n1016 10.6151
R1842 B.n1019 B.n1017 10.6151
R1843 B.n1020 B.n1019 10.6151
R1844 B.n1021 B.n1020 10.6151
R1845 B.n1022 B.n1021 10.6151
R1846 B.n1024 B.n1022 10.6151
R1847 B.n1025 B.n1024 10.6151
R1848 B.n1026 B.n1025 10.6151
R1849 B.n1027 B.n1026 10.6151
R1850 B.n1029 B.n1027 10.6151
R1851 B.n1030 B.n1029 10.6151
R1852 B.n1031 B.n1030 10.6151
R1853 B.n1032 B.n1031 10.6151
R1854 B.n1034 B.n1032 10.6151
R1855 B.n1035 B.n1034 10.6151
R1856 B.n1036 B.n1035 10.6151
R1857 B.n1037 B.n1036 10.6151
R1858 B.n1039 B.n1037 10.6151
R1859 B.n1040 B.n1039 10.6151
R1860 B.n1041 B.n1040 10.6151
R1861 B.n1042 B.n1041 10.6151
R1862 B.n1044 B.n1042 10.6151
R1863 B.n1045 B.n1044 10.6151
R1864 B.n1046 B.n1045 10.6151
R1865 B.n1047 B.n1046 10.6151
R1866 B.n1049 B.n1047 10.6151
R1867 B.n1050 B.n1049 10.6151
R1868 B.n1051 B.n1050 10.6151
R1869 B.n1052 B.n1051 10.6151
R1870 B.n1054 B.n1052 10.6151
R1871 B.n1055 B.n1054 10.6151
R1872 B.n1056 B.n1055 10.6151
R1873 B.n1057 B.n1056 10.6151
R1874 B.n1059 B.n1057 10.6151
R1875 B.n1060 B.n1059 10.6151
R1876 B.n1061 B.n1060 10.6151
R1877 B.n1062 B.n1061 10.6151
R1878 B.n1064 B.n1062 10.6151
R1879 B.n1065 B.n1064 10.6151
R1880 B.n1066 B.n1065 10.6151
R1881 B.n1067 B.n1066 10.6151
R1882 B.n1069 B.n1067 10.6151
R1883 B.n1070 B.n1069 10.6151
R1884 B.n595 B.n521 10.6151
R1885 B.n596 B.n595 10.6151
R1886 B.n597 B.n596 10.6151
R1887 B.n597 B.n591 10.6151
R1888 B.n603 B.n591 10.6151
R1889 B.n604 B.n603 10.6151
R1890 B.n605 B.n604 10.6151
R1891 B.n605 B.n589 10.6151
R1892 B.n611 B.n589 10.6151
R1893 B.n612 B.n611 10.6151
R1894 B.n613 B.n612 10.6151
R1895 B.n613 B.n587 10.6151
R1896 B.n619 B.n587 10.6151
R1897 B.n620 B.n619 10.6151
R1898 B.n621 B.n620 10.6151
R1899 B.n621 B.n585 10.6151
R1900 B.n627 B.n585 10.6151
R1901 B.n628 B.n627 10.6151
R1902 B.n629 B.n628 10.6151
R1903 B.n629 B.n583 10.6151
R1904 B.n635 B.n583 10.6151
R1905 B.n636 B.n635 10.6151
R1906 B.n637 B.n636 10.6151
R1907 B.n637 B.n581 10.6151
R1908 B.n643 B.n581 10.6151
R1909 B.n644 B.n643 10.6151
R1910 B.n645 B.n644 10.6151
R1911 B.n645 B.n579 10.6151
R1912 B.n651 B.n579 10.6151
R1913 B.n652 B.n651 10.6151
R1914 B.n653 B.n652 10.6151
R1915 B.n653 B.n577 10.6151
R1916 B.n659 B.n577 10.6151
R1917 B.n660 B.n659 10.6151
R1918 B.n661 B.n660 10.6151
R1919 B.n661 B.n575 10.6151
R1920 B.n667 B.n575 10.6151
R1921 B.n668 B.n667 10.6151
R1922 B.n669 B.n668 10.6151
R1923 B.n669 B.n573 10.6151
R1924 B.n675 B.n573 10.6151
R1925 B.n676 B.n675 10.6151
R1926 B.n677 B.n676 10.6151
R1927 B.n677 B.n571 10.6151
R1928 B.n683 B.n571 10.6151
R1929 B.n684 B.n683 10.6151
R1930 B.n685 B.n684 10.6151
R1931 B.n685 B.n569 10.6151
R1932 B.n691 B.n569 10.6151
R1933 B.n692 B.n691 10.6151
R1934 B.n693 B.n692 10.6151
R1935 B.n693 B.n567 10.6151
R1936 B.n699 B.n567 10.6151
R1937 B.n700 B.n699 10.6151
R1938 B.n701 B.n700 10.6151
R1939 B.n701 B.n565 10.6151
R1940 B.n707 B.n565 10.6151
R1941 B.n708 B.n707 10.6151
R1942 B.n709 B.n708 10.6151
R1943 B.n709 B.n563 10.6151
R1944 B.n715 B.n563 10.6151
R1945 B.n716 B.n715 10.6151
R1946 B.n718 B.n559 10.6151
R1947 B.n724 B.n559 10.6151
R1948 B.n725 B.n724 10.6151
R1949 B.n726 B.n725 10.6151
R1950 B.n726 B.n557 10.6151
R1951 B.n732 B.n557 10.6151
R1952 B.n733 B.n732 10.6151
R1953 B.n737 B.n733 10.6151
R1954 B.n743 B.n555 10.6151
R1955 B.n744 B.n743 10.6151
R1956 B.n745 B.n744 10.6151
R1957 B.n745 B.n553 10.6151
R1958 B.n751 B.n553 10.6151
R1959 B.n752 B.n751 10.6151
R1960 B.n753 B.n752 10.6151
R1961 B.n753 B.n551 10.6151
R1962 B.n759 B.n551 10.6151
R1963 B.n760 B.n759 10.6151
R1964 B.n761 B.n760 10.6151
R1965 B.n761 B.n549 10.6151
R1966 B.n767 B.n549 10.6151
R1967 B.n768 B.n767 10.6151
R1968 B.n769 B.n768 10.6151
R1969 B.n769 B.n547 10.6151
R1970 B.n775 B.n547 10.6151
R1971 B.n776 B.n775 10.6151
R1972 B.n777 B.n776 10.6151
R1973 B.n777 B.n545 10.6151
R1974 B.n783 B.n545 10.6151
R1975 B.n784 B.n783 10.6151
R1976 B.n785 B.n784 10.6151
R1977 B.n785 B.n543 10.6151
R1978 B.n791 B.n543 10.6151
R1979 B.n792 B.n791 10.6151
R1980 B.n793 B.n792 10.6151
R1981 B.n793 B.n541 10.6151
R1982 B.n799 B.n541 10.6151
R1983 B.n800 B.n799 10.6151
R1984 B.n801 B.n800 10.6151
R1985 B.n801 B.n539 10.6151
R1986 B.n807 B.n539 10.6151
R1987 B.n808 B.n807 10.6151
R1988 B.n809 B.n808 10.6151
R1989 B.n809 B.n537 10.6151
R1990 B.n815 B.n537 10.6151
R1991 B.n816 B.n815 10.6151
R1992 B.n817 B.n816 10.6151
R1993 B.n817 B.n535 10.6151
R1994 B.n823 B.n535 10.6151
R1995 B.n824 B.n823 10.6151
R1996 B.n825 B.n824 10.6151
R1997 B.n825 B.n533 10.6151
R1998 B.n831 B.n533 10.6151
R1999 B.n832 B.n831 10.6151
R2000 B.n833 B.n832 10.6151
R2001 B.n833 B.n531 10.6151
R2002 B.n839 B.n531 10.6151
R2003 B.n840 B.n839 10.6151
R2004 B.n841 B.n840 10.6151
R2005 B.n841 B.n529 10.6151
R2006 B.n847 B.n529 10.6151
R2007 B.n848 B.n847 10.6151
R2008 B.n849 B.n848 10.6151
R2009 B.n849 B.n527 10.6151
R2010 B.n855 B.n527 10.6151
R2011 B.n856 B.n855 10.6151
R2012 B.n857 B.n856 10.6151
R2013 B.n857 B.n525 10.6151
R2014 B.n863 B.n525 10.6151
R2015 B.n864 B.n863 10.6151
R2016 B.n870 B.n869 10.6151
R2017 B.n871 B.n870 10.6151
R2018 B.n871 B.n513 10.6151
R2019 B.n881 B.n513 10.6151
R2020 B.n882 B.n881 10.6151
R2021 B.n883 B.n882 10.6151
R2022 B.n883 B.n505 10.6151
R2023 B.n893 B.n505 10.6151
R2024 B.n894 B.n893 10.6151
R2025 B.n895 B.n894 10.6151
R2026 B.n895 B.n497 10.6151
R2027 B.n905 B.n497 10.6151
R2028 B.n906 B.n905 10.6151
R2029 B.n907 B.n906 10.6151
R2030 B.n907 B.n489 10.6151
R2031 B.n917 B.n489 10.6151
R2032 B.n918 B.n917 10.6151
R2033 B.n919 B.n918 10.6151
R2034 B.n919 B.n481 10.6151
R2035 B.n929 B.n481 10.6151
R2036 B.n930 B.n929 10.6151
R2037 B.n931 B.n930 10.6151
R2038 B.n931 B.n473 10.6151
R2039 B.n941 B.n473 10.6151
R2040 B.n942 B.n941 10.6151
R2041 B.n943 B.n942 10.6151
R2042 B.n943 B.n465 10.6151
R2043 B.n953 B.n465 10.6151
R2044 B.n954 B.n953 10.6151
R2045 B.n955 B.n954 10.6151
R2046 B.n955 B.n457 10.6151
R2047 B.n965 B.n457 10.6151
R2048 B.n966 B.n965 10.6151
R2049 B.n967 B.n966 10.6151
R2050 B.n967 B.n449 10.6151
R2051 B.n977 B.n449 10.6151
R2052 B.n978 B.n977 10.6151
R2053 B.n979 B.n978 10.6151
R2054 B.n979 B.n441 10.6151
R2055 B.n989 B.n441 10.6151
R2056 B.n990 B.n989 10.6151
R2057 B.n991 B.n990 10.6151
R2058 B.n991 B.n433 10.6151
R2059 B.n1002 B.n433 10.6151
R2060 B.n1003 B.n1002 10.6151
R2061 B.n1004 B.n1003 10.6151
R2062 B.n1004 B.n0 10.6151
R2063 B.n1166 B.n1 10.6151
R2064 B.n1166 B.n1165 10.6151
R2065 B.n1165 B.n1164 10.6151
R2066 B.n1164 B.n10 10.6151
R2067 B.n1158 B.n10 10.6151
R2068 B.n1158 B.n1157 10.6151
R2069 B.n1157 B.n1156 10.6151
R2070 B.n1156 B.n17 10.6151
R2071 B.n1150 B.n17 10.6151
R2072 B.n1150 B.n1149 10.6151
R2073 B.n1149 B.n1148 10.6151
R2074 B.n1148 B.n24 10.6151
R2075 B.n1142 B.n24 10.6151
R2076 B.n1142 B.n1141 10.6151
R2077 B.n1141 B.n1140 10.6151
R2078 B.n1140 B.n31 10.6151
R2079 B.n1134 B.n31 10.6151
R2080 B.n1134 B.n1133 10.6151
R2081 B.n1133 B.n1132 10.6151
R2082 B.n1132 B.n38 10.6151
R2083 B.n1126 B.n38 10.6151
R2084 B.n1126 B.n1125 10.6151
R2085 B.n1125 B.n1124 10.6151
R2086 B.n1124 B.n45 10.6151
R2087 B.n1118 B.n45 10.6151
R2088 B.n1118 B.n1117 10.6151
R2089 B.n1117 B.n1116 10.6151
R2090 B.n1116 B.n52 10.6151
R2091 B.n1110 B.n52 10.6151
R2092 B.n1110 B.n1109 10.6151
R2093 B.n1109 B.n1108 10.6151
R2094 B.n1108 B.n59 10.6151
R2095 B.n1102 B.n59 10.6151
R2096 B.n1102 B.n1101 10.6151
R2097 B.n1101 B.n1100 10.6151
R2098 B.n1100 B.n66 10.6151
R2099 B.n1094 B.n66 10.6151
R2100 B.n1094 B.n1093 10.6151
R2101 B.n1093 B.n1092 10.6151
R2102 B.n1092 B.n73 10.6151
R2103 B.n1086 B.n73 10.6151
R2104 B.n1086 B.n1085 10.6151
R2105 B.n1085 B.n1084 10.6151
R2106 B.n1084 B.n80 10.6151
R2107 B.n1078 B.n80 10.6151
R2108 B.n1078 B.n1077 10.6151
R2109 B.n1077 B.n1076 10.6151
R2110 B.n288 B.n287 6.5566
R2111 B.n304 B.n160 6.5566
R2112 B.n718 B.n717 6.5566
R2113 B.n737 B.n736 6.5566
R2114 B.n511 B.t9 5.86957
R2115 B.t13 B.n1089 5.86957
R2116 B.n287 B.n286 4.05904
R2117 B.n307 B.n160 4.05904
R2118 B.n717 B.n716 4.05904
R2119 B.n736 B.n555 4.05904
R2120 B.n1172 B.n0 2.81026
R2121 B.n1172 B.n1 2.81026
R2122 VP.n15 VP.t2 225.333
R2123 VP.n36 VP.t1 192.498
R2124 VP.n43 VP.t7 192.498
R2125 VP.n55 VP.t4 192.498
R2126 VP.n63 VP.t0 192.498
R2127 VP.n33 VP.t5 192.498
R2128 VP.n25 VP.t6 192.498
R2129 VP.n14 VP.t3 192.498
R2130 VP.n16 VP.n13 161.3
R2131 VP.n18 VP.n17 161.3
R2132 VP.n19 VP.n12 161.3
R2133 VP.n21 VP.n20 161.3
R2134 VP.n22 VP.n11 161.3
R2135 VP.n24 VP.n23 161.3
R2136 VP.n26 VP.n10 161.3
R2137 VP.n28 VP.n27 161.3
R2138 VP.n29 VP.n9 161.3
R2139 VP.n31 VP.n30 161.3
R2140 VP.n32 VP.n8 161.3
R2141 VP.n62 VP.n0 161.3
R2142 VP.n61 VP.n60 161.3
R2143 VP.n59 VP.n1 161.3
R2144 VP.n58 VP.n57 161.3
R2145 VP.n56 VP.n2 161.3
R2146 VP.n54 VP.n53 161.3
R2147 VP.n52 VP.n3 161.3
R2148 VP.n51 VP.n50 161.3
R2149 VP.n49 VP.n4 161.3
R2150 VP.n48 VP.n47 161.3
R2151 VP.n46 VP.n5 161.3
R2152 VP.n45 VP.n44 161.3
R2153 VP.n42 VP.n6 161.3
R2154 VP.n41 VP.n40 161.3
R2155 VP.n39 VP.n7 161.3
R2156 VP.n38 VP.n37 161.3
R2157 VP.n36 VP.n35 94.6082
R2158 VP.n64 VP.n63 94.6082
R2159 VP.n34 VP.n33 94.6082
R2160 VP.n15 VP.n14 66.7382
R2161 VP.n50 VP.n49 56.5193
R2162 VP.n20 VP.n19 56.5193
R2163 VP.n35 VP.n34 55.3481
R2164 VP.n42 VP.n41 43.4072
R2165 VP.n57 VP.n1 43.4072
R2166 VP.n27 VP.n9 43.4072
R2167 VP.n41 VP.n7 37.5796
R2168 VP.n61 VP.n1 37.5796
R2169 VP.n31 VP.n9 37.5796
R2170 VP.n37 VP.n7 24.4675
R2171 VP.n44 VP.n42 24.4675
R2172 VP.n48 VP.n5 24.4675
R2173 VP.n49 VP.n48 24.4675
R2174 VP.n50 VP.n3 24.4675
R2175 VP.n54 VP.n3 24.4675
R2176 VP.n57 VP.n56 24.4675
R2177 VP.n62 VP.n61 24.4675
R2178 VP.n32 VP.n31 24.4675
R2179 VP.n20 VP.n11 24.4675
R2180 VP.n24 VP.n11 24.4675
R2181 VP.n27 VP.n26 24.4675
R2182 VP.n18 VP.n13 24.4675
R2183 VP.n19 VP.n18 24.4675
R2184 VP.n44 VP.n43 19.0848
R2185 VP.n56 VP.n55 19.0848
R2186 VP.n26 VP.n25 19.0848
R2187 VP.n37 VP.n36 16.1487
R2188 VP.n63 VP.n62 16.1487
R2189 VP.n33 VP.n32 16.1487
R2190 VP.n16 VP.n15 9.37577
R2191 VP.n43 VP.n5 5.38324
R2192 VP.n55 VP.n54 5.38324
R2193 VP.n25 VP.n24 5.38324
R2194 VP.n14 VP.n13 5.38324
R2195 VP.n34 VP.n8 0.278367
R2196 VP.n38 VP.n35 0.278367
R2197 VP.n64 VP.n0 0.278367
R2198 VP.n17 VP.n16 0.189894
R2199 VP.n17 VP.n12 0.189894
R2200 VP.n21 VP.n12 0.189894
R2201 VP.n22 VP.n21 0.189894
R2202 VP.n23 VP.n22 0.189894
R2203 VP.n23 VP.n10 0.189894
R2204 VP.n28 VP.n10 0.189894
R2205 VP.n29 VP.n28 0.189894
R2206 VP.n30 VP.n29 0.189894
R2207 VP.n30 VP.n8 0.189894
R2208 VP.n39 VP.n38 0.189894
R2209 VP.n40 VP.n39 0.189894
R2210 VP.n40 VP.n6 0.189894
R2211 VP.n45 VP.n6 0.189894
R2212 VP.n46 VP.n45 0.189894
R2213 VP.n47 VP.n46 0.189894
R2214 VP.n47 VP.n4 0.189894
R2215 VP.n51 VP.n4 0.189894
R2216 VP.n52 VP.n51 0.189894
R2217 VP.n53 VP.n52 0.189894
R2218 VP.n53 VP.n2 0.189894
R2219 VP.n58 VP.n2 0.189894
R2220 VP.n59 VP.n58 0.189894
R2221 VP.n60 VP.n59 0.189894
R2222 VP.n60 VP.n0 0.189894
R2223 VP VP.n64 0.153454
R2224 VDD1 VDD1.n0 63.9513
R2225 VDD1.n3 VDD1.n2 63.8366
R2226 VDD1.n3 VDD1.n1 63.8366
R2227 VDD1.n5 VDD1.n4 62.7206
R2228 VDD1.n5 VDD1.n3 51.3069
R2229 VDD1 VDD1.n5 1.11472
R2230 VDD1.n4 VDD1.t1 1.03769
R2231 VDD1.n4 VDD1.t2 1.03769
R2232 VDD1.n0 VDD1.t5 1.03769
R2233 VDD1.n0 VDD1.t4 1.03769
R2234 VDD1.n2 VDD1.t3 1.03769
R2235 VDD1.n2 VDD1.t7 1.03769
R2236 VDD1.n1 VDD1.t6 1.03769
R2237 VDD1.n1 VDD1.t0 1.03769
C0 VN VTAIL 13.348599f
C1 VDD2 VDD1 1.66534f
C2 VP VTAIL 13.3627f
C3 VN VP 8.716691f
C4 VDD1 VTAIL 10.5507f
C5 VN VDD1 0.150952f
C6 VDD2 VTAIL 10.603701f
C7 VDD1 VP 13.6862f
C8 VDD2 VN 13.3415f
C9 VDD2 VP 0.496928f
C10 VDD2 B 5.679608f
C11 VDD1 B 6.094728f
C12 VTAIL B 14.575555f
C13 VN B 15.314769f
C14 VP B 13.743596f
C15 VDD1.t5 B 0.372333f
C16 VDD1.t4 B 0.372333f
C17 VDD1.n0 B 3.41698f
C18 VDD1.t6 B 0.372333f
C19 VDD1.t0 B 0.372333f
C20 VDD1.n1 B 3.41597f
C21 VDD1.t3 B 0.372333f
C22 VDD1.t7 B 0.372333f
C23 VDD1.n2 B 3.41597f
C24 VDD1.n3 B 3.59992f
C25 VDD1.t1 B 0.372333f
C26 VDD1.t2 B 0.372333f
C27 VDD1.n4 B 3.40749f
C28 VDD1.n5 B 3.3956f
C29 VP.n0 B 0.029785f
C30 VP.t0 B 2.83823f
C31 VP.n1 B 0.018526f
C32 VP.n2 B 0.022592f
C33 VP.t4 B 2.83823f
C34 VP.n3 B 0.042106f
C35 VP.n4 B 0.022592f
C36 VP.n5 B 0.025891f
C37 VP.n6 B 0.022592f
C38 VP.n7 B 0.04544f
C39 VP.n8 B 0.029785f
C40 VP.t5 B 2.83823f
C41 VP.n9 B 0.018526f
C42 VP.n10 B 0.022592f
C43 VP.t6 B 2.83823f
C44 VP.n11 B 0.042106f
C45 VP.n12 B 0.022592f
C46 VP.n13 B 0.025891f
C47 VP.t2 B 3.00055f
C48 VP.t3 B 2.83823f
C49 VP.n14 B 1.04004f
C50 VP.n15 B 1.03085f
C51 VP.n16 B 0.196531f
C52 VP.n17 B 0.022592f
C53 VP.n18 B 0.042106f
C54 VP.n19 B 0.03298f
C55 VP.n20 B 0.03298f
C56 VP.n21 B 0.022592f
C57 VP.n22 B 0.022592f
C58 VP.n23 B 0.022592f
C59 VP.n24 B 0.025891f
C60 VP.n25 B 0.983676f
C61 VP.n26 B 0.037532f
C62 VP.n27 B 0.044099f
C63 VP.n28 B 0.022592f
C64 VP.n29 B 0.022592f
C65 VP.n30 B 0.022592f
C66 VP.n31 B 0.04544f
C67 VP.n32 B 0.035038f
C68 VP.n33 B 1.06102f
C69 VP.n34 B 1.44962f
C70 VP.n35 B 1.46429f
C71 VP.t1 B 2.83823f
C72 VP.n36 B 1.06102f
C73 VP.n37 B 0.035038f
C74 VP.n38 B 0.029785f
C75 VP.n39 B 0.022592f
C76 VP.n40 B 0.022592f
C77 VP.n41 B 0.018526f
C78 VP.n42 B 0.044099f
C79 VP.t7 B 2.83823f
C80 VP.n43 B 0.983676f
C81 VP.n44 B 0.037532f
C82 VP.n45 B 0.022592f
C83 VP.n46 B 0.022592f
C84 VP.n47 B 0.022592f
C85 VP.n48 B 0.042106f
C86 VP.n49 B 0.03298f
C87 VP.n50 B 0.03298f
C88 VP.n51 B 0.022592f
C89 VP.n52 B 0.022592f
C90 VP.n53 B 0.022592f
C91 VP.n54 B 0.025891f
C92 VP.n55 B 0.983676f
C93 VP.n56 B 0.037532f
C94 VP.n57 B 0.044099f
C95 VP.n58 B 0.022592f
C96 VP.n59 B 0.022592f
C97 VP.n60 B 0.022592f
C98 VP.n61 B 0.04544f
C99 VP.n62 B 0.035038f
C100 VP.n63 B 1.06102f
C101 VP.n64 B 0.031569f
C102 VDD2.t5 B 0.367583f
C103 VDD2.t3 B 0.367583f
C104 VDD2.n0 B 3.37239f
C105 VDD2.t6 B 0.367583f
C106 VDD2.t7 B 0.367583f
C107 VDD2.n1 B 3.37239f
C108 VDD2.n2 B 3.50343f
C109 VDD2.t2 B 0.367583f
C110 VDD2.t4 B 0.367583f
C111 VDD2.n3 B 3.36404f
C112 VDD2.n4 B 3.32197f
C113 VDD2.t0 B 0.367583f
C114 VDD2.t1 B 0.367583f
C115 VDD2.n5 B 3.37235f
C116 VTAIL.t15 B 0.276841f
C117 VTAIL.t12 B 0.276841f
C118 VTAIL.n0 B 2.48149f
C119 VTAIL.n1 B 0.316544f
C120 VTAIL.t8 B 3.17129f
C121 VTAIL.n2 B 0.406101f
C122 VTAIL.t2 B 3.17129f
C123 VTAIL.n3 B 0.406101f
C124 VTAIL.t0 B 0.276841f
C125 VTAIL.t4 B 0.276841f
C126 VTAIL.n4 B 2.48149f
C127 VTAIL.n5 B 0.451758f
C128 VTAIL.t5 B 3.17129f
C129 VTAIL.n6 B 1.73939f
C130 VTAIL.t10 B 3.17131f
C131 VTAIL.n7 B 1.73937f
C132 VTAIL.t14 B 0.276841f
C133 VTAIL.t13 B 0.276841f
C134 VTAIL.n8 B 2.48149f
C135 VTAIL.n9 B 0.451751f
C136 VTAIL.t11 B 3.17131f
C137 VTAIL.n10 B 0.406078f
C138 VTAIL.t7 B 3.17131f
C139 VTAIL.n11 B 0.406078f
C140 VTAIL.t6 B 0.276841f
C141 VTAIL.t3 B 0.276841f
C142 VTAIL.n12 B 2.48149f
C143 VTAIL.n13 B 0.451751f
C144 VTAIL.t1 B 3.17129f
C145 VTAIL.n14 B 1.73939f
C146 VTAIL.t9 B 3.17129f
C147 VTAIL.n15 B 1.73595f
C148 VN.n0 B 0.029343f
C149 VN.t0 B 2.79611f
C150 VN.n1 B 0.018251f
C151 VN.n2 B 0.022257f
C152 VN.t1 B 2.79611f
C153 VN.n3 B 0.041481f
C154 VN.n4 B 0.022257f
C155 VN.n5 B 0.025507f
C156 VN.t2 B 2.95602f
C157 VN.t4 B 2.79611f
C158 VN.n6 B 1.02461f
C159 VN.n7 B 1.01555f
C160 VN.n8 B 0.193614f
C161 VN.n9 B 0.022257f
C162 VN.n10 B 0.041481f
C163 VN.n11 B 0.032491f
C164 VN.n12 B 0.032491f
C165 VN.n13 B 0.022257f
C166 VN.n14 B 0.022257f
C167 VN.n15 B 0.022257f
C168 VN.n16 B 0.025507f
C169 VN.n17 B 0.969078f
C170 VN.n18 B 0.036975f
C171 VN.n19 B 0.043445f
C172 VN.n20 B 0.022257f
C173 VN.n21 B 0.022257f
C174 VN.n22 B 0.022257f
C175 VN.n23 B 0.044766f
C176 VN.n24 B 0.034518f
C177 VN.n25 B 1.04527f
C178 VN.n26 B 0.031101f
C179 VN.n27 B 0.029343f
C180 VN.t5 B 2.79611f
C181 VN.n28 B 0.018251f
C182 VN.n29 B 0.022257f
C183 VN.t3 B 2.79611f
C184 VN.n30 B 0.041481f
C185 VN.n31 B 0.022257f
C186 VN.n32 B 0.025507f
C187 VN.t6 B 2.95602f
C188 VN.t7 B 2.79611f
C189 VN.n33 B 1.02461f
C190 VN.n34 B 1.01555f
C191 VN.n35 B 0.193614f
C192 VN.n36 B 0.022257f
C193 VN.n37 B 0.041481f
C194 VN.n38 B 0.032491f
C195 VN.n39 B 0.032491f
C196 VN.n40 B 0.022257f
C197 VN.n41 B 0.022257f
C198 VN.n42 B 0.022257f
C199 VN.n43 B 0.025507f
C200 VN.n44 B 0.969078f
C201 VN.n45 B 0.036975f
C202 VN.n46 B 0.043445f
C203 VN.n47 B 0.022257f
C204 VN.n48 B 0.022257f
C205 VN.n49 B 0.022257f
C206 VN.n50 B 0.044766f
C207 VN.n51 B 0.034518f
C208 VN.n52 B 1.04527f
C209 VN.n53 B 1.43988f
.ends

