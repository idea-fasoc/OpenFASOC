* NGSPICE file created from diff_pair_sample_1784.ext - technology: sky130A

.subckt diff_pair_sample_1784 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t7 VN.t0 VTAIL.t14 B.t5 sky130_fd_pr__nfet_01v8 ad=1.78695 pd=11.16 as=1.78695 ps=11.16 w=10.83 l=2.16
X1 VDD1.t7 VP.t0 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.78695 pd=11.16 as=4.2237 ps=22.44 w=10.83 l=2.16
X2 VDD1.t6 VP.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.78695 pd=11.16 as=4.2237 ps=22.44 w=10.83 l=2.16
X3 VTAIL.t7 VP.t2 VDD1.t5 B.t7 sky130_fd_pr__nfet_01v8 ad=1.78695 pd=11.16 as=1.78695 ps=11.16 w=10.83 l=2.16
X4 VTAIL.t12 VN.t1 VDD2.t6 B.t7 sky130_fd_pr__nfet_01v8 ad=1.78695 pd=11.16 as=1.78695 ps=11.16 w=10.83 l=2.16
X5 VTAIL.t8 VN.t2 VDD2.t5 B.t0 sky130_fd_pr__nfet_01v8 ad=4.2237 pd=22.44 as=1.78695 ps=11.16 w=10.83 l=2.16
X6 VDD2.t4 VN.t3 VTAIL.t11 B.t1 sky130_fd_pr__nfet_01v8 ad=1.78695 pd=11.16 as=4.2237 ps=22.44 w=10.83 l=2.16
X7 VTAIL.t6 VP.t3 VDD1.t4 B.t6 sky130_fd_pr__nfet_01v8 ad=1.78695 pd=11.16 as=1.78695 ps=11.16 w=10.83 l=2.16
X8 B.t21 B.t19 B.t20 B.t9 sky130_fd_pr__nfet_01v8 ad=4.2237 pd=22.44 as=0 ps=0 w=10.83 l=2.16
X9 VDD1.t3 VP.t4 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=1.78695 pd=11.16 as=1.78695 ps=11.16 w=10.83 l=2.16
X10 B.t18 B.t16 B.t17 B.t13 sky130_fd_pr__nfet_01v8 ad=4.2237 pd=22.44 as=0 ps=0 w=10.83 l=2.16
X11 VTAIL.t0 VP.t5 VDD1.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=4.2237 pd=22.44 as=1.78695 ps=11.16 w=10.83 l=2.16
X12 VDD2.t3 VN.t4 VTAIL.t10 B.t2 sky130_fd_pr__nfet_01v8 ad=1.78695 pd=11.16 as=4.2237 ps=22.44 w=10.83 l=2.16
X13 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=4.2237 pd=22.44 as=0 ps=0 w=10.83 l=2.16
X14 VTAIL.t15 VN.t5 VDD2.t2 B.t4 sky130_fd_pr__nfet_01v8 ad=4.2237 pd=22.44 as=1.78695 ps=11.16 w=10.83 l=2.16
X15 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=4.2237 pd=22.44 as=0 ps=0 w=10.83 l=2.16
X16 VTAIL.t13 VN.t6 VDD2.t1 B.t6 sky130_fd_pr__nfet_01v8 ad=1.78695 pd=11.16 as=1.78695 ps=11.16 w=10.83 l=2.16
X17 VDD2.t0 VN.t7 VTAIL.t9 B.t3 sky130_fd_pr__nfet_01v8 ad=1.78695 pd=11.16 as=1.78695 ps=11.16 w=10.83 l=2.16
X18 VTAIL.t4 VP.t6 VDD1.t1 B.t4 sky130_fd_pr__nfet_01v8 ad=4.2237 pd=22.44 as=1.78695 ps=11.16 w=10.83 l=2.16
X19 VDD1.t0 VP.t7 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.78695 pd=11.16 as=1.78695 ps=11.16 w=10.83 l=2.16
R0 VN.n47 VN.n25 161.3
R1 VN.n46 VN.n45 161.3
R2 VN.n44 VN.n26 161.3
R3 VN.n43 VN.n42 161.3
R4 VN.n41 VN.n27 161.3
R5 VN.n39 VN.n38 161.3
R6 VN.n37 VN.n28 161.3
R7 VN.n36 VN.n35 161.3
R8 VN.n34 VN.n29 161.3
R9 VN.n33 VN.n32 161.3
R10 VN.n22 VN.n0 161.3
R11 VN.n21 VN.n20 161.3
R12 VN.n19 VN.n1 161.3
R13 VN.n18 VN.n17 161.3
R14 VN.n16 VN.n2 161.3
R15 VN.n14 VN.n13 161.3
R16 VN.n12 VN.n3 161.3
R17 VN.n11 VN.n10 161.3
R18 VN.n9 VN.n4 161.3
R19 VN.n8 VN.n7 161.3
R20 VN.n6 VN.t5 152.594
R21 VN.n31 VN.t4 152.594
R22 VN.n5 VN.t7 120.835
R23 VN.n15 VN.t1 120.835
R24 VN.n23 VN.t3 120.835
R25 VN.n30 VN.t6 120.835
R26 VN.n40 VN.t0 120.835
R27 VN.n48 VN.t2 120.835
R28 VN.n24 VN.n23 99.257
R29 VN.n49 VN.n48 99.257
R30 VN.n6 VN.n5 59.5219
R31 VN.n31 VN.n30 59.5219
R32 VN VN.n49 48.1648
R33 VN.n17 VN.n1 41.4647
R34 VN.n42 VN.n26 41.4647
R35 VN.n10 VN.n9 40.4934
R36 VN.n10 VN.n3 40.4934
R37 VN.n35 VN.n34 40.4934
R38 VN.n35 VN.n28 40.4934
R39 VN.n21 VN.n1 39.5221
R40 VN.n46 VN.n26 39.5221
R41 VN.n9 VN.n8 24.4675
R42 VN.n14 VN.n3 24.4675
R43 VN.n17 VN.n16 24.4675
R44 VN.n22 VN.n21 24.4675
R45 VN.n34 VN.n33 24.4675
R46 VN.n42 VN.n41 24.4675
R47 VN.n39 VN.n28 24.4675
R48 VN.n47 VN.n46 24.4675
R49 VN.n16 VN.n15 12.4787
R50 VN.n41 VN.n40 12.4787
R51 VN.n8 VN.n5 11.9893
R52 VN.n15 VN.n14 11.9893
R53 VN.n33 VN.n30 11.9893
R54 VN.n40 VN.n39 11.9893
R55 VN.n23 VN.n22 11.5
R56 VN.n48 VN.n47 11.5
R57 VN.n32 VN.n31 9.80091
R58 VN.n7 VN.n6 9.80091
R59 VN.n49 VN.n25 0.278367
R60 VN.n24 VN.n0 0.278367
R61 VN.n45 VN.n25 0.189894
R62 VN.n45 VN.n44 0.189894
R63 VN.n44 VN.n43 0.189894
R64 VN.n43 VN.n27 0.189894
R65 VN.n38 VN.n27 0.189894
R66 VN.n38 VN.n37 0.189894
R67 VN.n37 VN.n36 0.189894
R68 VN.n36 VN.n29 0.189894
R69 VN.n32 VN.n29 0.189894
R70 VN.n7 VN.n4 0.189894
R71 VN.n11 VN.n4 0.189894
R72 VN.n12 VN.n11 0.189894
R73 VN.n13 VN.n12 0.189894
R74 VN.n13 VN.n2 0.189894
R75 VN.n18 VN.n2 0.189894
R76 VN.n19 VN.n18 0.189894
R77 VN.n20 VN.n19 0.189894
R78 VN.n20 VN.n0 0.189894
R79 VN VN.n24 0.153454
R80 VTAIL.n466 VTAIL.n414 289.615
R81 VTAIL.n54 VTAIL.n2 289.615
R82 VTAIL.n112 VTAIL.n60 289.615
R83 VTAIL.n172 VTAIL.n120 289.615
R84 VTAIL.n408 VTAIL.n356 289.615
R85 VTAIL.n348 VTAIL.n296 289.615
R86 VTAIL.n290 VTAIL.n238 289.615
R87 VTAIL.n230 VTAIL.n178 289.615
R88 VTAIL.n433 VTAIL.n432 185
R89 VTAIL.n430 VTAIL.n429 185
R90 VTAIL.n439 VTAIL.n438 185
R91 VTAIL.n441 VTAIL.n440 185
R92 VTAIL.n426 VTAIL.n425 185
R93 VTAIL.n447 VTAIL.n446 185
R94 VTAIL.n450 VTAIL.n449 185
R95 VTAIL.n448 VTAIL.n422 185
R96 VTAIL.n455 VTAIL.n421 185
R97 VTAIL.n457 VTAIL.n456 185
R98 VTAIL.n459 VTAIL.n458 185
R99 VTAIL.n418 VTAIL.n417 185
R100 VTAIL.n465 VTAIL.n464 185
R101 VTAIL.n467 VTAIL.n466 185
R102 VTAIL.n21 VTAIL.n20 185
R103 VTAIL.n18 VTAIL.n17 185
R104 VTAIL.n27 VTAIL.n26 185
R105 VTAIL.n29 VTAIL.n28 185
R106 VTAIL.n14 VTAIL.n13 185
R107 VTAIL.n35 VTAIL.n34 185
R108 VTAIL.n38 VTAIL.n37 185
R109 VTAIL.n36 VTAIL.n10 185
R110 VTAIL.n43 VTAIL.n9 185
R111 VTAIL.n45 VTAIL.n44 185
R112 VTAIL.n47 VTAIL.n46 185
R113 VTAIL.n6 VTAIL.n5 185
R114 VTAIL.n53 VTAIL.n52 185
R115 VTAIL.n55 VTAIL.n54 185
R116 VTAIL.n79 VTAIL.n78 185
R117 VTAIL.n76 VTAIL.n75 185
R118 VTAIL.n85 VTAIL.n84 185
R119 VTAIL.n87 VTAIL.n86 185
R120 VTAIL.n72 VTAIL.n71 185
R121 VTAIL.n93 VTAIL.n92 185
R122 VTAIL.n96 VTAIL.n95 185
R123 VTAIL.n94 VTAIL.n68 185
R124 VTAIL.n101 VTAIL.n67 185
R125 VTAIL.n103 VTAIL.n102 185
R126 VTAIL.n105 VTAIL.n104 185
R127 VTAIL.n64 VTAIL.n63 185
R128 VTAIL.n111 VTAIL.n110 185
R129 VTAIL.n113 VTAIL.n112 185
R130 VTAIL.n139 VTAIL.n138 185
R131 VTAIL.n136 VTAIL.n135 185
R132 VTAIL.n145 VTAIL.n144 185
R133 VTAIL.n147 VTAIL.n146 185
R134 VTAIL.n132 VTAIL.n131 185
R135 VTAIL.n153 VTAIL.n152 185
R136 VTAIL.n156 VTAIL.n155 185
R137 VTAIL.n154 VTAIL.n128 185
R138 VTAIL.n161 VTAIL.n127 185
R139 VTAIL.n163 VTAIL.n162 185
R140 VTAIL.n165 VTAIL.n164 185
R141 VTAIL.n124 VTAIL.n123 185
R142 VTAIL.n171 VTAIL.n170 185
R143 VTAIL.n173 VTAIL.n172 185
R144 VTAIL.n409 VTAIL.n408 185
R145 VTAIL.n407 VTAIL.n406 185
R146 VTAIL.n360 VTAIL.n359 185
R147 VTAIL.n401 VTAIL.n400 185
R148 VTAIL.n399 VTAIL.n398 185
R149 VTAIL.n397 VTAIL.n363 185
R150 VTAIL.n367 VTAIL.n364 185
R151 VTAIL.n392 VTAIL.n391 185
R152 VTAIL.n390 VTAIL.n389 185
R153 VTAIL.n369 VTAIL.n368 185
R154 VTAIL.n384 VTAIL.n383 185
R155 VTAIL.n382 VTAIL.n381 185
R156 VTAIL.n373 VTAIL.n372 185
R157 VTAIL.n376 VTAIL.n375 185
R158 VTAIL.n349 VTAIL.n348 185
R159 VTAIL.n347 VTAIL.n346 185
R160 VTAIL.n300 VTAIL.n299 185
R161 VTAIL.n341 VTAIL.n340 185
R162 VTAIL.n339 VTAIL.n338 185
R163 VTAIL.n337 VTAIL.n303 185
R164 VTAIL.n307 VTAIL.n304 185
R165 VTAIL.n332 VTAIL.n331 185
R166 VTAIL.n330 VTAIL.n329 185
R167 VTAIL.n309 VTAIL.n308 185
R168 VTAIL.n324 VTAIL.n323 185
R169 VTAIL.n322 VTAIL.n321 185
R170 VTAIL.n313 VTAIL.n312 185
R171 VTAIL.n316 VTAIL.n315 185
R172 VTAIL.n291 VTAIL.n290 185
R173 VTAIL.n289 VTAIL.n288 185
R174 VTAIL.n242 VTAIL.n241 185
R175 VTAIL.n283 VTAIL.n282 185
R176 VTAIL.n281 VTAIL.n280 185
R177 VTAIL.n279 VTAIL.n245 185
R178 VTAIL.n249 VTAIL.n246 185
R179 VTAIL.n274 VTAIL.n273 185
R180 VTAIL.n272 VTAIL.n271 185
R181 VTAIL.n251 VTAIL.n250 185
R182 VTAIL.n266 VTAIL.n265 185
R183 VTAIL.n264 VTAIL.n263 185
R184 VTAIL.n255 VTAIL.n254 185
R185 VTAIL.n258 VTAIL.n257 185
R186 VTAIL.n231 VTAIL.n230 185
R187 VTAIL.n229 VTAIL.n228 185
R188 VTAIL.n182 VTAIL.n181 185
R189 VTAIL.n223 VTAIL.n222 185
R190 VTAIL.n221 VTAIL.n220 185
R191 VTAIL.n219 VTAIL.n185 185
R192 VTAIL.n189 VTAIL.n186 185
R193 VTAIL.n214 VTAIL.n213 185
R194 VTAIL.n212 VTAIL.n211 185
R195 VTAIL.n191 VTAIL.n190 185
R196 VTAIL.n206 VTAIL.n205 185
R197 VTAIL.n204 VTAIL.n203 185
R198 VTAIL.n195 VTAIL.n194 185
R199 VTAIL.n198 VTAIL.n197 185
R200 VTAIL.t11 VTAIL.n431 149.524
R201 VTAIL.t15 VTAIL.n19 149.524
R202 VTAIL.t2 VTAIL.n77 149.524
R203 VTAIL.t0 VTAIL.n137 149.524
R204 VTAIL.t1 VTAIL.n374 149.524
R205 VTAIL.t4 VTAIL.n314 149.524
R206 VTAIL.t10 VTAIL.n256 149.524
R207 VTAIL.t8 VTAIL.n196 149.524
R208 VTAIL.n432 VTAIL.n429 104.615
R209 VTAIL.n439 VTAIL.n429 104.615
R210 VTAIL.n440 VTAIL.n439 104.615
R211 VTAIL.n440 VTAIL.n425 104.615
R212 VTAIL.n447 VTAIL.n425 104.615
R213 VTAIL.n449 VTAIL.n447 104.615
R214 VTAIL.n449 VTAIL.n448 104.615
R215 VTAIL.n448 VTAIL.n421 104.615
R216 VTAIL.n457 VTAIL.n421 104.615
R217 VTAIL.n458 VTAIL.n457 104.615
R218 VTAIL.n458 VTAIL.n417 104.615
R219 VTAIL.n465 VTAIL.n417 104.615
R220 VTAIL.n466 VTAIL.n465 104.615
R221 VTAIL.n20 VTAIL.n17 104.615
R222 VTAIL.n27 VTAIL.n17 104.615
R223 VTAIL.n28 VTAIL.n27 104.615
R224 VTAIL.n28 VTAIL.n13 104.615
R225 VTAIL.n35 VTAIL.n13 104.615
R226 VTAIL.n37 VTAIL.n35 104.615
R227 VTAIL.n37 VTAIL.n36 104.615
R228 VTAIL.n36 VTAIL.n9 104.615
R229 VTAIL.n45 VTAIL.n9 104.615
R230 VTAIL.n46 VTAIL.n45 104.615
R231 VTAIL.n46 VTAIL.n5 104.615
R232 VTAIL.n53 VTAIL.n5 104.615
R233 VTAIL.n54 VTAIL.n53 104.615
R234 VTAIL.n78 VTAIL.n75 104.615
R235 VTAIL.n85 VTAIL.n75 104.615
R236 VTAIL.n86 VTAIL.n85 104.615
R237 VTAIL.n86 VTAIL.n71 104.615
R238 VTAIL.n93 VTAIL.n71 104.615
R239 VTAIL.n95 VTAIL.n93 104.615
R240 VTAIL.n95 VTAIL.n94 104.615
R241 VTAIL.n94 VTAIL.n67 104.615
R242 VTAIL.n103 VTAIL.n67 104.615
R243 VTAIL.n104 VTAIL.n103 104.615
R244 VTAIL.n104 VTAIL.n63 104.615
R245 VTAIL.n111 VTAIL.n63 104.615
R246 VTAIL.n112 VTAIL.n111 104.615
R247 VTAIL.n138 VTAIL.n135 104.615
R248 VTAIL.n145 VTAIL.n135 104.615
R249 VTAIL.n146 VTAIL.n145 104.615
R250 VTAIL.n146 VTAIL.n131 104.615
R251 VTAIL.n153 VTAIL.n131 104.615
R252 VTAIL.n155 VTAIL.n153 104.615
R253 VTAIL.n155 VTAIL.n154 104.615
R254 VTAIL.n154 VTAIL.n127 104.615
R255 VTAIL.n163 VTAIL.n127 104.615
R256 VTAIL.n164 VTAIL.n163 104.615
R257 VTAIL.n164 VTAIL.n123 104.615
R258 VTAIL.n171 VTAIL.n123 104.615
R259 VTAIL.n172 VTAIL.n171 104.615
R260 VTAIL.n408 VTAIL.n407 104.615
R261 VTAIL.n407 VTAIL.n359 104.615
R262 VTAIL.n400 VTAIL.n359 104.615
R263 VTAIL.n400 VTAIL.n399 104.615
R264 VTAIL.n399 VTAIL.n363 104.615
R265 VTAIL.n367 VTAIL.n363 104.615
R266 VTAIL.n391 VTAIL.n367 104.615
R267 VTAIL.n391 VTAIL.n390 104.615
R268 VTAIL.n390 VTAIL.n368 104.615
R269 VTAIL.n383 VTAIL.n368 104.615
R270 VTAIL.n383 VTAIL.n382 104.615
R271 VTAIL.n382 VTAIL.n372 104.615
R272 VTAIL.n375 VTAIL.n372 104.615
R273 VTAIL.n348 VTAIL.n347 104.615
R274 VTAIL.n347 VTAIL.n299 104.615
R275 VTAIL.n340 VTAIL.n299 104.615
R276 VTAIL.n340 VTAIL.n339 104.615
R277 VTAIL.n339 VTAIL.n303 104.615
R278 VTAIL.n307 VTAIL.n303 104.615
R279 VTAIL.n331 VTAIL.n307 104.615
R280 VTAIL.n331 VTAIL.n330 104.615
R281 VTAIL.n330 VTAIL.n308 104.615
R282 VTAIL.n323 VTAIL.n308 104.615
R283 VTAIL.n323 VTAIL.n322 104.615
R284 VTAIL.n322 VTAIL.n312 104.615
R285 VTAIL.n315 VTAIL.n312 104.615
R286 VTAIL.n290 VTAIL.n289 104.615
R287 VTAIL.n289 VTAIL.n241 104.615
R288 VTAIL.n282 VTAIL.n241 104.615
R289 VTAIL.n282 VTAIL.n281 104.615
R290 VTAIL.n281 VTAIL.n245 104.615
R291 VTAIL.n249 VTAIL.n245 104.615
R292 VTAIL.n273 VTAIL.n249 104.615
R293 VTAIL.n273 VTAIL.n272 104.615
R294 VTAIL.n272 VTAIL.n250 104.615
R295 VTAIL.n265 VTAIL.n250 104.615
R296 VTAIL.n265 VTAIL.n264 104.615
R297 VTAIL.n264 VTAIL.n254 104.615
R298 VTAIL.n257 VTAIL.n254 104.615
R299 VTAIL.n230 VTAIL.n229 104.615
R300 VTAIL.n229 VTAIL.n181 104.615
R301 VTAIL.n222 VTAIL.n181 104.615
R302 VTAIL.n222 VTAIL.n221 104.615
R303 VTAIL.n221 VTAIL.n185 104.615
R304 VTAIL.n189 VTAIL.n185 104.615
R305 VTAIL.n213 VTAIL.n189 104.615
R306 VTAIL.n213 VTAIL.n212 104.615
R307 VTAIL.n212 VTAIL.n190 104.615
R308 VTAIL.n205 VTAIL.n190 104.615
R309 VTAIL.n205 VTAIL.n204 104.615
R310 VTAIL.n204 VTAIL.n194 104.615
R311 VTAIL.n197 VTAIL.n194 104.615
R312 VTAIL.n432 VTAIL.t11 52.3082
R313 VTAIL.n20 VTAIL.t15 52.3082
R314 VTAIL.n78 VTAIL.t2 52.3082
R315 VTAIL.n138 VTAIL.t0 52.3082
R316 VTAIL.n375 VTAIL.t1 52.3082
R317 VTAIL.n315 VTAIL.t4 52.3082
R318 VTAIL.n257 VTAIL.t10 52.3082
R319 VTAIL.n197 VTAIL.t8 52.3082
R320 VTAIL.n355 VTAIL.n354 48.5706
R321 VTAIL.n237 VTAIL.n236 48.5706
R322 VTAIL.n1 VTAIL.n0 48.5704
R323 VTAIL.n119 VTAIL.n118 48.5704
R324 VTAIL.n471 VTAIL.n470 35.0944
R325 VTAIL.n59 VTAIL.n58 35.0944
R326 VTAIL.n117 VTAIL.n116 35.0944
R327 VTAIL.n177 VTAIL.n176 35.0944
R328 VTAIL.n413 VTAIL.n412 35.0944
R329 VTAIL.n353 VTAIL.n352 35.0944
R330 VTAIL.n295 VTAIL.n294 35.0944
R331 VTAIL.n235 VTAIL.n234 35.0944
R332 VTAIL.n471 VTAIL.n413 23.8496
R333 VTAIL.n235 VTAIL.n177 23.8496
R334 VTAIL.n456 VTAIL.n455 13.1884
R335 VTAIL.n44 VTAIL.n43 13.1884
R336 VTAIL.n102 VTAIL.n101 13.1884
R337 VTAIL.n162 VTAIL.n161 13.1884
R338 VTAIL.n398 VTAIL.n397 13.1884
R339 VTAIL.n338 VTAIL.n337 13.1884
R340 VTAIL.n280 VTAIL.n279 13.1884
R341 VTAIL.n220 VTAIL.n219 13.1884
R342 VTAIL.n454 VTAIL.n422 12.8005
R343 VTAIL.n459 VTAIL.n420 12.8005
R344 VTAIL.n42 VTAIL.n10 12.8005
R345 VTAIL.n47 VTAIL.n8 12.8005
R346 VTAIL.n100 VTAIL.n68 12.8005
R347 VTAIL.n105 VTAIL.n66 12.8005
R348 VTAIL.n160 VTAIL.n128 12.8005
R349 VTAIL.n165 VTAIL.n126 12.8005
R350 VTAIL.n401 VTAIL.n362 12.8005
R351 VTAIL.n396 VTAIL.n364 12.8005
R352 VTAIL.n341 VTAIL.n302 12.8005
R353 VTAIL.n336 VTAIL.n304 12.8005
R354 VTAIL.n283 VTAIL.n244 12.8005
R355 VTAIL.n278 VTAIL.n246 12.8005
R356 VTAIL.n223 VTAIL.n184 12.8005
R357 VTAIL.n218 VTAIL.n186 12.8005
R358 VTAIL.n451 VTAIL.n450 12.0247
R359 VTAIL.n460 VTAIL.n418 12.0247
R360 VTAIL.n39 VTAIL.n38 12.0247
R361 VTAIL.n48 VTAIL.n6 12.0247
R362 VTAIL.n97 VTAIL.n96 12.0247
R363 VTAIL.n106 VTAIL.n64 12.0247
R364 VTAIL.n157 VTAIL.n156 12.0247
R365 VTAIL.n166 VTAIL.n124 12.0247
R366 VTAIL.n402 VTAIL.n360 12.0247
R367 VTAIL.n393 VTAIL.n392 12.0247
R368 VTAIL.n342 VTAIL.n300 12.0247
R369 VTAIL.n333 VTAIL.n332 12.0247
R370 VTAIL.n284 VTAIL.n242 12.0247
R371 VTAIL.n275 VTAIL.n274 12.0247
R372 VTAIL.n224 VTAIL.n182 12.0247
R373 VTAIL.n215 VTAIL.n214 12.0247
R374 VTAIL.n446 VTAIL.n424 11.249
R375 VTAIL.n464 VTAIL.n463 11.249
R376 VTAIL.n34 VTAIL.n12 11.249
R377 VTAIL.n52 VTAIL.n51 11.249
R378 VTAIL.n92 VTAIL.n70 11.249
R379 VTAIL.n110 VTAIL.n109 11.249
R380 VTAIL.n152 VTAIL.n130 11.249
R381 VTAIL.n170 VTAIL.n169 11.249
R382 VTAIL.n406 VTAIL.n405 11.249
R383 VTAIL.n389 VTAIL.n366 11.249
R384 VTAIL.n346 VTAIL.n345 11.249
R385 VTAIL.n329 VTAIL.n306 11.249
R386 VTAIL.n288 VTAIL.n287 11.249
R387 VTAIL.n271 VTAIL.n248 11.249
R388 VTAIL.n228 VTAIL.n227 11.249
R389 VTAIL.n211 VTAIL.n188 11.249
R390 VTAIL.n445 VTAIL.n426 10.4732
R391 VTAIL.n467 VTAIL.n416 10.4732
R392 VTAIL.n33 VTAIL.n14 10.4732
R393 VTAIL.n55 VTAIL.n4 10.4732
R394 VTAIL.n91 VTAIL.n72 10.4732
R395 VTAIL.n113 VTAIL.n62 10.4732
R396 VTAIL.n151 VTAIL.n132 10.4732
R397 VTAIL.n173 VTAIL.n122 10.4732
R398 VTAIL.n409 VTAIL.n358 10.4732
R399 VTAIL.n388 VTAIL.n369 10.4732
R400 VTAIL.n349 VTAIL.n298 10.4732
R401 VTAIL.n328 VTAIL.n309 10.4732
R402 VTAIL.n291 VTAIL.n240 10.4732
R403 VTAIL.n270 VTAIL.n251 10.4732
R404 VTAIL.n231 VTAIL.n180 10.4732
R405 VTAIL.n210 VTAIL.n191 10.4732
R406 VTAIL.n433 VTAIL.n431 10.2747
R407 VTAIL.n21 VTAIL.n19 10.2747
R408 VTAIL.n79 VTAIL.n77 10.2747
R409 VTAIL.n139 VTAIL.n137 10.2747
R410 VTAIL.n376 VTAIL.n374 10.2747
R411 VTAIL.n316 VTAIL.n314 10.2747
R412 VTAIL.n258 VTAIL.n256 10.2747
R413 VTAIL.n198 VTAIL.n196 10.2747
R414 VTAIL.n442 VTAIL.n441 9.69747
R415 VTAIL.n468 VTAIL.n414 9.69747
R416 VTAIL.n30 VTAIL.n29 9.69747
R417 VTAIL.n56 VTAIL.n2 9.69747
R418 VTAIL.n88 VTAIL.n87 9.69747
R419 VTAIL.n114 VTAIL.n60 9.69747
R420 VTAIL.n148 VTAIL.n147 9.69747
R421 VTAIL.n174 VTAIL.n120 9.69747
R422 VTAIL.n410 VTAIL.n356 9.69747
R423 VTAIL.n385 VTAIL.n384 9.69747
R424 VTAIL.n350 VTAIL.n296 9.69747
R425 VTAIL.n325 VTAIL.n324 9.69747
R426 VTAIL.n292 VTAIL.n238 9.69747
R427 VTAIL.n267 VTAIL.n266 9.69747
R428 VTAIL.n232 VTAIL.n178 9.69747
R429 VTAIL.n207 VTAIL.n206 9.69747
R430 VTAIL.n470 VTAIL.n469 9.45567
R431 VTAIL.n58 VTAIL.n57 9.45567
R432 VTAIL.n116 VTAIL.n115 9.45567
R433 VTAIL.n176 VTAIL.n175 9.45567
R434 VTAIL.n412 VTAIL.n411 9.45567
R435 VTAIL.n352 VTAIL.n351 9.45567
R436 VTAIL.n294 VTAIL.n293 9.45567
R437 VTAIL.n234 VTAIL.n233 9.45567
R438 VTAIL.n469 VTAIL.n468 9.3005
R439 VTAIL.n416 VTAIL.n415 9.3005
R440 VTAIL.n463 VTAIL.n462 9.3005
R441 VTAIL.n461 VTAIL.n460 9.3005
R442 VTAIL.n420 VTAIL.n419 9.3005
R443 VTAIL.n435 VTAIL.n434 9.3005
R444 VTAIL.n437 VTAIL.n436 9.3005
R445 VTAIL.n428 VTAIL.n427 9.3005
R446 VTAIL.n443 VTAIL.n442 9.3005
R447 VTAIL.n445 VTAIL.n444 9.3005
R448 VTAIL.n424 VTAIL.n423 9.3005
R449 VTAIL.n452 VTAIL.n451 9.3005
R450 VTAIL.n454 VTAIL.n453 9.3005
R451 VTAIL.n57 VTAIL.n56 9.3005
R452 VTAIL.n4 VTAIL.n3 9.3005
R453 VTAIL.n51 VTAIL.n50 9.3005
R454 VTAIL.n49 VTAIL.n48 9.3005
R455 VTAIL.n8 VTAIL.n7 9.3005
R456 VTAIL.n23 VTAIL.n22 9.3005
R457 VTAIL.n25 VTAIL.n24 9.3005
R458 VTAIL.n16 VTAIL.n15 9.3005
R459 VTAIL.n31 VTAIL.n30 9.3005
R460 VTAIL.n33 VTAIL.n32 9.3005
R461 VTAIL.n12 VTAIL.n11 9.3005
R462 VTAIL.n40 VTAIL.n39 9.3005
R463 VTAIL.n42 VTAIL.n41 9.3005
R464 VTAIL.n115 VTAIL.n114 9.3005
R465 VTAIL.n62 VTAIL.n61 9.3005
R466 VTAIL.n109 VTAIL.n108 9.3005
R467 VTAIL.n107 VTAIL.n106 9.3005
R468 VTAIL.n66 VTAIL.n65 9.3005
R469 VTAIL.n81 VTAIL.n80 9.3005
R470 VTAIL.n83 VTAIL.n82 9.3005
R471 VTAIL.n74 VTAIL.n73 9.3005
R472 VTAIL.n89 VTAIL.n88 9.3005
R473 VTAIL.n91 VTAIL.n90 9.3005
R474 VTAIL.n70 VTAIL.n69 9.3005
R475 VTAIL.n98 VTAIL.n97 9.3005
R476 VTAIL.n100 VTAIL.n99 9.3005
R477 VTAIL.n175 VTAIL.n174 9.3005
R478 VTAIL.n122 VTAIL.n121 9.3005
R479 VTAIL.n169 VTAIL.n168 9.3005
R480 VTAIL.n167 VTAIL.n166 9.3005
R481 VTAIL.n126 VTAIL.n125 9.3005
R482 VTAIL.n141 VTAIL.n140 9.3005
R483 VTAIL.n143 VTAIL.n142 9.3005
R484 VTAIL.n134 VTAIL.n133 9.3005
R485 VTAIL.n149 VTAIL.n148 9.3005
R486 VTAIL.n151 VTAIL.n150 9.3005
R487 VTAIL.n130 VTAIL.n129 9.3005
R488 VTAIL.n158 VTAIL.n157 9.3005
R489 VTAIL.n160 VTAIL.n159 9.3005
R490 VTAIL.n378 VTAIL.n377 9.3005
R491 VTAIL.n380 VTAIL.n379 9.3005
R492 VTAIL.n371 VTAIL.n370 9.3005
R493 VTAIL.n386 VTAIL.n385 9.3005
R494 VTAIL.n388 VTAIL.n387 9.3005
R495 VTAIL.n366 VTAIL.n365 9.3005
R496 VTAIL.n394 VTAIL.n393 9.3005
R497 VTAIL.n396 VTAIL.n395 9.3005
R498 VTAIL.n411 VTAIL.n410 9.3005
R499 VTAIL.n358 VTAIL.n357 9.3005
R500 VTAIL.n405 VTAIL.n404 9.3005
R501 VTAIL.n403 VTAIL.n402 9.3005
R502 VTAIL.n362 VTAIL.n361 9.3005
R503 VTAIL.n318 VTAIL.n317 9.3005
R504 VTAIL.n320 VTAIL.n319 9.3005
R505 VTAIL.n311 VTAIL.n310 9.3005
R506 VTAIL.n326 VTAIL.n325 9.3005
R507 VTAIL.n328 VTAIL.n327 9.3005
R508 VTAIL.n306 VTAIL.n305 9.3005
R509 VTAIL.n334 VTAIL.n333 9.3005
R510 VTAIL.n336 VTAIL.n335 9.3005
R511 VTAIL.n351 VTAIL.n350 9.3005
R512 VTAIL.n298 VTAIL.n297 9.3005
R513 VTAIL.n345 VTAIL.n344 9.3005
R514 VTAIL.n343 VTAIL.n342 9.3005
R515 VTAIL.n302 VTAIL.n301 9.3005
R516 VTAIL.n260 VTAIL.n259 9.3005
R517 VTAIL.n262 VTAIL.n261 9.3005
R518 VTAIL.n253 VTAIL.n252 9.3005
R519 VTAIL.n268 VTAIL.n267 9.3005
R520 VTAIL.n270 VTAIL.n269 9.3005
R521 VTAIL.n248 VTAIL.n247 9.3005
R522 VTAIL.n276 VTAIL.n275 9.3005
R523 VTAIL.n278 VTAIL.n277 9.3005
R524 VTAIL.n293 VTAIL.n292 9.3005
R525 VTAIL.n240 VTAIL.n239 9.3005
R526 VTAIL.n287 VTAIL.n286 9.3005
R527 VTAIL.n285 VTAIL.n284 9.3005
R528 VTAIL.n244 VTAIL.n243 9.3005
R529 VTAIL.n200 VTAIL.n199 9.3005
R530 VTAIL.n202 VTAIL.n201 9.3005
R531 VTAIL.n193 VTAIL.n192 9.3005
R532 VTAIL.n208 VTAIL.n207 9.3005
R533 VTAIL.n210 VTAIL.n209 9.3005
R534 VTAIL.n188 VTAIL.n187 9.3005
R535 VTAIL.n216 VTAIL.n215 9.3005
R536 VTAIL.n218 VTAIL.n217 9.3005
R537 VTAIL.n233 VTAIL.n232 9.3005
R538 VTAIL.n180 VTAIL.n179 9.3005
R539 VTAIL.n227 VTAIL.n226 9.3005
R540 VTAIL.n225 VTAIL.n224 9.3005
R541 VTAIL.n184 VTAIL.n183 9.3005
R542 VTAIL.n438 VTAIL.n428 8.92171
R543 VTAIL.n26 VTAIL.n16 8.92171
R544 VTAIL.n84 VTAIL.n74 8.92171
R545 VTAIL.n144 VTAIL.n134 8.92171
R546 VTAIL.n381 VTAIL.n371 8.92171
R547 VTAIL.n321 VTAIL.n311 8.92171
R548 VTAIL.n263 VTAIL.n253 8.92171
R549 VTAIL.n203 VTAIL.n193 8.92171
R550 VTAIL.n437 VTAIL.n430 8.14595
R551 VTAIL.n25 VTAIL.n18 8.14595
R552 VTAIL.n83 VTAIL.n76 8.14595
R553 VTAIL.n143 VTAIL.n136 8.14595
R554 VTAIL.n380 VTAIL.n373 8.14595
R555 VTAIL.n320 VTAIL.n313 8.14595
R556 VTAIL.n262 VTAIL.n255 8.14595
R557 VTAIL.n202 VTAIL.n195 8.14595
R558 VTAIL.n434 VTAIL.n433 7.3702
R559 VTAIL.n22 VTAIL.n21 7.3702
R560 VTAIL.n80 VTAIL.n79 7.3702
R561 VTAIL.n140 VTAIL.n139 7.3702
R562 VTAIL.n377 VTAIL.n376 7.3702
R563 VTAIL.n317 VTAIL.n316 7.3702
R564 VTAIL.n259 VTAIL.n258 7.3702
R565 VTAIL.n199 VTAIL.n198 7.3702
R566 VTAIL.n434 VTAIL.n430 5.81868
R567 VTAIL.n22 VTAIL.n18 5.81868
R568 VTAIL.n80 VTAIL.n76 5.81868
R569 VTAIL.n140 VTAIL.n136 5.81868
R570 VTAIL.n377 VTAIL.n373 5.81868
R571 VTAIL.n317 VTAIL.n313 5.81868
R572 VTAIL.n259 VTAIL.n255 5.81868
R573 VTAIL.n199 VTAIL.n195 5.81868
R574 VTAIL.n438 VTAIL.n437 5.04292
R575 VTAIL.n26 VTAIL.n25 5.04292
R576 VTAIL.n84 VTAIL.n83 5.04292
R577 VTAIL.n144 VTAIL.n143 5.04292
R578 VTAIL.n381 VTAIL.n380 5.04292
R579 VTAIL.n321 VTAIL.n320 5.04292
R580 VTAIL.n263 VTAIL.n262 5.04292
R581 VTAIL.n203 VTAIL.n202 5.04292
R582 VTAIL.n441 VTAIL.n428 4.26717
R583 VTAIL.n470 VTAIL.n414 4.26717
R584 VTAIL.n29 VTAIL.n16 4.26717
R585 VTAIL.n58 VTAIL.n2 4.26717
R586 VTAIL.n87 VTAIL.n74 4.26717
R587 VTAIL.n116 VTAIL.n60 4.26717
R588 VTAIL.n147 VTAIL.n134 4.26717
R589 VTAIL.n176 VTAIL.n120 4.26717
R590 VTAIL.n412 VTAIL.n356 4.26717
R591 VTAIL.n384 VTAIL.n371 4.26717
R592 VTAIL.n352 VTAIL.n296 4.26717
R593 VTAIL.n324 VTAIL.n311 4.26717
R594 VTAIL.n294 VTAIL.n238 4.26717
R595 VTAIL.n266 VTAIL.n253 4.26717
R596 VTAIL.n234 VTAIL.n178 4.26717
R597 VTAIL.n206 VTAIL.n193 4.26717
R598 VTAIL.n442 VTAIL.n426 3.49141
R599 VTAIL.n468 VTAIL.n467 3.49141
R600 VTAIL.n30 VTAIL.n14 3.49141
R601 VTAIL.n56 VTAIL.n55 3.49141
R602 VTAIL.n88 VTAIL.n72 3.49141
R603 VTAIL.n114 VTAIL.n113 3.49141
R604 VTAIL.n148 VTAIL.n132 3.49141
R605 VTAIL.n174 VTAIL.n173 3.49141
R606 VTAIL.n410 VTAIL.n409 3.49141
R607 VTAIL.n385 VTAIL.n369 3.49141
R608 VTAIL.n350 VTAIL.n349 3.49141
R609 VTAIL.n325 VTAIL.n309 3.49141
R610 VTAIL.n292 VTAIL.n291 3.49141
R611 VTAIL.n267 VTAIL.n251 3.49141
R612 VTAIL.n232 VTAIL.n231 3.49141
R613 VTAIL.n207 VTAIL.n191 3.49141
R614 VTAIL.n435 VTAIL.n431 2.84303
R615 VTAIL.n23 VTAIL.n19 2.84303
R616 VTAIL.n81 VTAIL.n77 2.84303
R617 VTAIL.n141 VTAIL.n137 2.84303
R618 VTAIL.n378 VTAIL.n374 2.84303
R619 VTAIL.n318 VTAIL.n314 2.84303
R620 VTAIL.n260 VTAIL.n256 2.84303
R621 VTAIL.n200 VTAIL.n196 2.84303
R622 VTAIL.n446 VTAIL.n445 2.71565
R623 VTAIL.n464 VTAIL.n416 2.71565
R624 VTAIL.n34 VTAIL.n33 2.71565
R625 VTAIL.n52 VTAIL.n4 2.71565
R626 VTAIL.n92 VTAIL.n91 2.71565
R627 VTAIL.n110 VTAIL.n62 2.71565
R628 VTAIL.n152 VTAIL.n151 2.71565
R629 VTAIL.n170 VTAIL.n122 2.71565
R630 VTAIL.n406 VTAIL.n358 2.71565
R631 VTAIL.n389 VTAIL.n388 2.71565
R632 VTAIL.n346 VTAIL.n298 2.71565
R633 VTAIL.n329 VTAIL.n328 2.71565
R634 VTAIL.n288 VTAIL.n240 2.71565
R635 VTAIL.n271 VTAIL.n270 2.71565
R636 VTAIL.n228 VTAIL.n180 2.71565
R637 VTAIL.n211 VTAIL.n210 2.71565
R638 VTAIL.n237 VTAIL.n235 2.14705
R639 VTAIL.n295 VTAIL.n237 2.14705
R640 VTAIL.n355 VTAIL.n353 2.14705
R641 VTAIL.n413 VTAIL.n355 2.14705
R642 VTAIL.n177 VTAIL.n119 2.14705
R643 VTAIL.n119 VTAIL.n117 2.14705
R644 VTAIL.n59 VTAIL.n1 2.14705
R645 VTAIL VTAIL.n471 2.08886
R646 VTAIL.n450 VTAIL.n424 1.93989
R647 VTAIL.n463 VTAIL.n418 1.93989
R648 VTAIL.n38 VTAIL.n12 1.93989
R649 VTAIL.n51 VTAIL.n6 1.93989
R650 VTAIL.n96 VTAIL.n70 1.93989
R651 VTAIL.n109 VTAIL.n64 1.93989
R652 VTAIL.n156 VTAIL.n130 1.93989
R653 VTAIL.n169 VTAIL.n124 1.93989
R654 VTAIL.n405 VTAIL.n360 1.93989
R655 VTAIL.n392 VTAIL.n366 1.93989
R656 VTAIL.n345 VTAIL.n300 1.93989
R657 VTAIL.n332 VTAIL.n306 1.93989
R658 VTAIL.n287 VTAIL.n242 1.93989
R659 VTAIL.n274 VTAIL.n248 1.93989
R660 VTAIL.n227 VTAIL.n182 1.93989
R661 VTAIL.n214 VTAIL.n188 1.93989
R662 VTAIL.n0 VTAIL.t9 1.82875
R663 VTAIL.n0 VTAIL.t12 1.82875
R664 VTAIL.n118 VTAIL.t5 1.82875
R665 VTAIL.n118 VTAIL.t6 1.82875
R666 VTAIL.n354 VTAIL.t3 1.82875
R667 VTAIL.n354 VTAIL.t7 1.82875
R668 VTAIL.n236 VTAIL.t14 1.82875
R669 VTAIL.n236 VTAIL.t13 1.82875
R670 VTAIL.n451 VTAIL.n422 1.16414
R671 VTAIL.n460 VTAIL.n459 1.16414
R672 VTAIL.n39 VTAIL.n10 1.16414
R673 VTAIL.n48 VTAIL.n47 1.16414
R674 VTAIL.n97 VTAIL.n68 1.16414
R675 VTAIL.n106 VTAIL.n105 1.16414
R676 VTAIL.n157 VTAIL.n128 1.16414
R677 VTAIL.n166 VTAIL.n165 1.16414
R678 VTAIL.n402 VTAIL.n401 1.16414
R679 VTAIL.n393 VTAIL.n364 1.16414
R680 VTAIL.n342 VTAIL.n341 1.16414
R681 VTAIL.n333 VTAIL.n304 1.16414
R682 VTAIL.n284 VTAIL.n283 1.16414
R683 VTAIL.n275 VTAIL.n246 1.16414
R684 VTAIL.n224 VTAIL.n223 1.16414
R685 VTAIL.n215 VTAIL.n186 1.16414
R686 VTAIL.n353 VTAIL.n295 0.470328
R687 VTAIL.n117 VTAIL.n59 0.470328
R688 VTAIL.n455 VTAIL.n454 0.388379
R689 VTAIL.n456 VTAIL.n420 0.388379
R690 VTAIL.n43 VTAIL.n42 0.388379
R691 VTAIL.n44 VTAIL.n8 0.388379
R692 VTAIL.n101 VTAIL.n100 0.388379
R693 VTAIL.n102 VTAIL.n66 0.388379
R694 VTAIL.n161 VTAIL.n160 0.388379
R695 VTAIL.n162 VTAIL.n126 0.388379
R696 VTAIL.n398 VTAIL.n362 0.388379
R697 VTAIL.n397 VTAIL.n396 0.388379
R698 VTAIL.n338 VTAIL.n302 0.388379
R699 VTAIL.n337 VTAIL.n336 0.388379
R700 VTAIL.n280 VTAIL.n244 0.388379
R701 VTAIL.n279 VTAIL.n278 0.388379
R702 VTAIL.n220 VTAIL.n184 0.388379
R703 VTAIL.n219 VTAIL.n218 0.388379
R704 VTAIL.n436 VTAIL.n435 0.155672
R705 VTAIL.n436 VTAIL.n427 0.155672
R706 VTAIL.n443 VTAIL.n427 0.155672
R707 VTAIL.n444 VTAIL.n443 0.155672
R708 VTAIL.n444 VTAIL.n423 0.155672
R709 VTAIL.n452 VTAIL.n423 0.155672
R710 VTAIL.n453 VTAIL.n452 0.155672
R711 VTAIL.n453 VTAIL.n419 0.155672
R712 VTAIL.n461 VTAIL.n419 0.155672
R713 VTAIL.n462 VTAIL.n461 0.155672
R714 VTAIL.n462 VTAIL.n415 0.155672
R715 VTAIL.n469 VTAIL.n415 0.155672
R716 VTAIL.n24 VTAIL.n23 0.155672
R717 VTAIL.n24 VTAIL.n15 0.155672
R718 VTAIL.n31 VTAIL.n15 0.155672
R719 VTAIL.n32 VTAIL.n31 0.155672
R720 VTAIL.n32 VTAIL.n11 0.155672
R721 VTAIL.n40 VTAIL.n11 0.155672
R722 VTAIL.n41 VTAIL.n40 0.155672
R723 VTAIL.n41 VTAIL.n7 0.155672
R724 VTAIL.n49 VTAIL.n7 0.155672
R725 VTAIL.n50 VTAIL.n49 0.155672
R726 VTAIL.n50 VTAIL.n3 0.155672
R727 VTAIL.n57 VTAIL.n3 0.155672
R728 VTAIL.n82 VTAIL.n81 0.155672
R729 VTAIL.n82 VTAIL.n73 0.155672
R730 VTAIL.n89 VTAIL.n73 0.155672
R731 VTAIL.n90 VTAIL.n89 0.155672
R732 VTAIL.n90 VTAIL.n69 0.155672
R733 VTAIL.n98 VTAIL.n69 0.155672
R734 VTAIL.n99 VTAIL.n98 0.155672
R735 VTAIL.n99 VTAIL.n65 0.155672
R736 VTAIL.n107 VTAIL.n65 0.155672
R737 VTAIL.n108 VTAIL.n107 0.155672
R738 VTAIL.n108 VTAIL.n61 0.155672
R739 VTAIL.n115 VTAIL.n61 0.155672
R740 VTAIL.n142 VTAIL.n141 0.155672
R741 VTAIL.n142 VTAIL.n133 0.155672
R742 VTAIL.n149 VTAIL.n133 0.155672
R743 VTAIL.n150 VTAIL.n149 0.155672
R744 VTAIL.n150 VTAIL.n129 0.155672
R745 VTAIL.n158 VTAIL.n129 0.155672
R746 VTAIL.n159 VTAIL.n158 0.155672
R747 VTAIL.n159 VTAIL.n125 0.155672
R748 VTAIL.n167 VTAIL.n125 0.155672
R749 VTAIL.n168 VTAIL.n167 0.155672
R750 VTAIL.n168 VTAIL.n121 0.155672
R751 VTAIL.n175 VTAIL.n121 0.155672
R752 VTAIL.n411 VTAIL.n357 0.155672
R753 VTAIL.n404 VTAIL.n357 0.155672
R754 VTAIL.n404 VTAIL.n403 0.155672
R755 VTAIL.n403 VTAIL.n361 0.155672
R756 VTAIL.n395 VTAIL.n361 0.155672
R757 VTAIL.n395 VTAIL.n394 0.155672
R758 VTAIL.n394 VTAIL.n365 0.155672
R759 VTAIL.n387 VTAIL.n365 0.155672
R760 VTAIL.n387 VTAIL.n386 0.155672
R761 VTAIL.n386 VTAIL.n370 0.155672
R762 VTAIL.n379 VTAIL.n370 0.155672
R763 VTAIL.n379 VTAIL.n378 0.155672
R764 VTAIL.n351 VTAIL.n297 0.155672
R765 VTAIL.n344 VTAIL.n297 0.155672
R766 VTAIL.n344 VTAIL.n343 0.155672
R767 VTAIL.n343 VTAIL.n301 0.155672
R768 VTAIL.n335 VTAIL.n301 0.155672
R769 VTAIL.n335 VTAIL.n334 0.155672
R770 VTAIL.n334 VTAIL.n305 0.155672
R771 VTAIL.n327 VTAIL.n305 0.155672
R772 VTAIL.n327 VTAIL.n326 0.155672
R773 VTAIL.n326 VTAIL.n310 0.155672
R774 VTAIL.n319 VTAIL.n310 0.155672
R775 VTAIL.n319 VTAIL.n318 0.155672
R776 VTAIL.n293 VTAIL.n239 0.155672
R777 VTAIL.n286 VTAIL.n239 0.155672
R778 VTAIL.n286 VTAIL.n285 0.155672
R779 VTAIL.n285 VTAIL.n243 0.155672
R780 VTAIL.n277 VTAIL.n243 0.155672
R781 VTAIL.n277 VTAIL.n276 0.155672
R782 VTAIL.n276 VTAIL.n247 0.155672
R783 VTAIL.n269 VTAIL.n247 0.155672
R784 VTAIL.n269 VTAIL.n268 0.155672
R785 VTAIL.n268 VTAIL.n252 0.155672
R786 VTAIL.n261 VTAIL.n252 0.155672
R787 VTAIL.n261 VTAIL.n260 0.155672
R788 VTAIL.n233 VTAIL.n179 0.155672
R789 VTAIL.n226 VTAIL.n179 0.155672
R790 VTAIL.n226 VTAIL.n225 0.155672
R791 VTAIL.n225 VTAIL.n183 0.155672
R792 VTAIL.n217 VTAIL.n183 0.155672
R793 VTAIL.n217 VTAIL.n216 0.155672
R794 VTAIL.n216 VTAIL.n187 0.155672
R795 VTAIL.n209 VTAIL.n187 0.155672
R796 VTAIL.n209 VTAIL.n208 0.155672
R797 VTAIL.n208 VTAIL.n192 0.155672
R798 VTAIL.n201 VTAIL.n192 0.155672
R799 VTAIL.n201 VTAIL.n200 0.155672
R800 VTAIL VTAIL.n1 0.0586897
R801 VDD2.n2 VDD2.n1 66.2671
R802 VDD2.n2 VDD2.n0 66.2671
R803 VDD2 VDD2.n5 66.2643
R804 VDD2.n4 VDD2.n3 65.2494
R805 VDD2.n4 VDD2.n2 42.711
R806 VDD2.n5 VDD2.t1 1.82875
R807 VDD2.n5 VDD2.t3 1.82875
R808 VDD2.n3 VDD2.t5 1.82875
R809 VDD2.n3 VDD2.t7 1.82875
R810 VDD2.n1 VDD2.t6 1.82875
R811 VDD2.n1 VDD2.t4 1.82875
R812 VDD2.n0 VDD2.t2 1.82875
R813 VDD2.n0 VDD2.t0 1.82875
R814 VDD2 VDD2.n4 1.13197
R815 B.n797 B.n796 585
R816 B.n299 B.n126 585
R817 B.n298 B.n297 585
R818 B.n296 B.n295 585
R819 B.n294 B.n293 585
R820 B.n292 B.n291 585
R821 B.n290 B.n289 585
R822 B.n288 B.n287 585
R823 B.n286 B.n285 585
R824 B.n284 B.n283 585
R825 B.n282 B.n281 585
R826 B.n280 B.n279 585
R827 B.n278 B.n277 585
R828 B.n276 B.n275 585
R829 B.n274 B.n273 585
R830 B.n272 B.n271 585
R831 B.n270 B.n269 585
R832 B.n268 B.n267 585
R833 B.n266 B.n265 585
R834 B.n264 B.n263 585
R835 B.n262 B.n261 585
R836 B.n260 B.n259 585
R837 B.n258 B.n257 585
R838 B.n256 B.n255 585
R839 B.n254 B.n253 585
R840 B.n252 B.n251 585
R841 B.n250 B.n249 585
R842 B.n248 B.n247 585
R843 B.n246 B.n245 585
R844 B.n244 B.n243 585
R845 B.n242 B.n241 585
R846 B.n240 B.n239 585
R847 B.n238 B.n237 585
R848 B.n236 B.n235 585
R849 B.n234 B.n233 585
R850 B.n232 B.n231 585
R851 B.n230 B.n229 585
R852 B.n228 B.n227 585
R853 B.n226 B.n225 585
R854 B.n224 B.n223 585
R855 B.n222 B.n221 585
R856 B.n220 B.n219 585
R857 B.n218 B.n217 585
R858 B.n216 B.n215 585
R859 B.n214 B.n213 585
R860 B.n212 B.n211 585
R861 B.n210 B.n209 585
R862 B.n208 B.n207 585
R863 B.n206 B.n205 585
R864 B.n204 B.n203 585
R865 B.n202 B.n201 585
R866 B.n200 B.n199 585
R867 B.n198 B.n197 585
R868 B.n196 B.n195 585
R869 B.n194 B.n193 585
R870 B.n192 B.n191 585
R871 B.n190 B.n189 585
R872 B.n188 B.n187 585
R873 B.n186 B.n185 585
R874 B.n184 B.n183 585
R875 B.n182 B.n181 585
R876 B.n180 B.n179 585
R877 B.n178 B.n177 585
R878 B.n176 B.n175 585
R879 B.n174 B.n173 585
R880 B.n172 B.n171 585
R881 B.n170 B.n169 585
R882 B.n168 B.n167 585
R883 B.n166 B.n165 585
R884 B.n164 B.n163 585
R885 B.n162 B.n161 585
R886 B.n160 B.n159 585
R887 B.n158 B.n157 585
R888 B.n156 B.n155 585
R889 B.n154 B.n153 585
R890 B.n152 B.n151 585
R891 B.n150 B.n149 585
R892 B.n148 B.n147 585
R893 B.n146 B.n145 585
R894 B.n144 B.n143 585
R895 B.n142 B.n141 585
R896 B.n140 B.n139 585
R897 B.n138 B.n137 585
R898 B.n136 B.n135 585
R899 B.n134 B.n133 585
R900 B.n82 B.n81 585
R901 B.n795 B.n83 585
R902 B.n800 B.n83 585
R903 B.n794 B.n793 585
R904 B.n793 B.n79 585
R905 B.n792 B.n78 585
R906 B.n806 B.n78 585
R907 B.n791 B.n77 585
R908 B.n807 B.n77 585
R909 B.n790 B.n76 585
R910 B.n808 B.n76 585
R911 B.n789 B.n788 585
R912 B.n788 B.n72 585
R913 B.n787 B.n71 585
R914 B.n814 B.n71 585
R915 B.n786 B.n70 585
R916 B.n815 B.n70 585
R917 B.n785 B.n69 585
R918 B.n816 B.n69 585
R919 B.n784 B.n783 585
R920 B.n783 B.n65 585
R921 B.n782 B.n64 585
R922 B.n822 B.n64 585
R923 B.n781 B.n63 585
R924 B.n823 B.n63 585
R925 B.n780 B.n62 585
R926 B.n824 B.n62 585
R927 B.n779 B.n778 585
R928 B.n778 B.n58 585
R929 B.n777 B.n57 585
R930 B.n830 B.n57 585
R931 B.n776 B.n56 585
R932 B.n831 B.n56 585
R933 B.n775 B.n55 585
R934 B.n832 B.n55 585
R935 B.n774 B.n773 585
R936 B.n773 B.n54 585
R937 B.n772 B.n50 585
R938 B.n838 B.n50 585
R939 B.n771 B.n49 585
R940 B.n839 B.n49 585
R941 B.n770 B.n48 585
R942 B.n840 B.n48 585
R943 B.n769 B.n768 585
R944 B.n768 B.n44 585
R945 B.n767 B.n43 585
R946 B.n846 B.n43 585
R947 B.n766 B.n42 585
R948 B.n847 B.n42 585
R949 B.n765 B.n41 585
R950 B.n848 B.n41 585
R951 B.n764 B.n763 585
R952 B.n763 B.n37 585
R953 B.n762 B.n36 585
R954 B.n854 B.n36 585
R955 B.n761 B.n35 585
R956 B.n855 B.n35 585
R957 B.n760 B.n34 585
R958 B.n856 B.n34 585
R959 B.n759 B.n758 585
R960 B.n758 B.n30 585
R961 B.n757 B.n29 585
R962 B.n862 B.n29 585
R963 B.n756 B.n28 585
R964 B.n863 B.n28 585
R965 B.n755 B.n27 585
R966 B.n864 B.n27 585
R967 B.n754 B.n753 585
R968 B.n753 B.n23 585
R969 B.n752 B.n22 585
R970 B.n870 B.n22 585
R971 B.n751 B.n21 585
R972 B.n871 B.n21 585
R973 B.n750 B.n20 585
R974 B.n872 B.n20 585
R975 B.n749 B.n748 585
R976 B.n748 B.n16 585
R977 B.n747 B.n15 585
R978 B.n878 B.n15 585
R979 B.n746 B.n14 585
R980 B.n879 B.n14 585
R981 B.n745 B.n13 585
R982 B.n880 B.n13 585
R983 B.n744 B.n743 585
R984 B.n743 B.n12 585
R985 B.n742 B.n741 585
R986 B.n742 B.n8 585
R987 B.n740 B.n7 585
R988 B.n887 B.n7 585
R989 B.n739 B.n6 585
R990 B.n888 B.n6 585
R991 B.n738 B.n5 585
R992 B.n889 B.n5 585
R993 B.n737 B.n736 585
R994 B.n736 B.n4 585
R995 B.n735 B.n300 585
R996 B.n735 B.n734 585
R997 B.n725 B.n301 585
R998 B.n302 B.n301 585
R999 B.n727 B.n726 585
R1000 B.n728 B.n727 585
R1001 B.n724 B.n306 585
R1002 B.n310 B.n306 585
R1003 B.n723 B.n722 585
R1004 B.n722 B.n721 585
R1005 B.n308 B.n307 585
R1006 B.n309 B.n308 585
R1007 B.n714 B.n713 585
R1008 B.n715 B.n714 585
R1009 B.n712 B.n315 585
R1010 B.n315 B.n314 585
R1011 B.n711 B.n710 585
R1012 B.n710 B.n709 585
R1013 B.n317 B.n316 585
R1014 B.n318 B.n317 585
R1015 B.n702 B.n701 585
R1016 B.n703 B.n702 585
R1017 B.n700 B.n322 585
R1018 B.n326 B.n322 585
R1019 B.n699 B.n698 585
R1020 B.n698 B.n697 585
R1021 B.n324 B.n323 585
R1022 B.n325 B.n324 585
R1023 B.n690 B.n689 585
R1024 B.n691 B.n690 585
R1025 B.n688 B.n331 585
R1026 B.n331 B.n330 585
R1027 B.n687 B.n686 585
R1028 B.n686 B.n685 585
R1029 B.n333 B.n332 585
R1030 B.n334 B.n333 585
R1031 B.n678 B.n677 585
R1032 B.n679 B.n678 585
R1033 B.n676 B.n339 585
R1034 B.n339 B.n338 585
R1035 B.n675 B.n674 585
R1036 B.n674 B.n673 585
R1037 B.n341 B.n340 585
R1038 B.n342 B.n341 585
R1039 B.n666 B.n665 585
R1040 B.n667 B.n666 585
R1041 B.n664 B.n347 585
R1042 B.n347 B.n346 585
R1043 B.n663 B.n662 585
R1044 B.n662 B.n661 585
R1045 B.n349 B.n348 585
R1046 B.n654 B.n349 585
R1047 B.n653 B.n652 585
R1048 B.n655 B.n653 585
R1049 B.n651 B.n354 585
R1050 B.n354 B.n353 585
R1051 B.n650 B.n649 585
R1052 B.n649 B.n648 585
R1053 B.n356 B.n355 585
R1054 B.n357 B.n356 585
R1055 B.n641 B.n640 585
R1056 B.n642 B.n641 585
R1057 B.n639 B.n362 585
R1058 B.n362 B.n361 585
R1059 B.n638 B.n637 585
R1060 B.n637 B.n636 585
R1061 B.n364 B.n363 585
R1062 B.n365 B.n364 585
R1063 B.n629 B.n628 585
R1064 B.n630 B.n629 585
R1065 B.n627 B.n370 585
R1066 B.n370 B.n369 585
R1067 B.n626 B.n625 585
R1068 B.n625 B.n624 585
R1069 B.n372 B.n371 585
R1070 B.n373 B.n372 585
R1071 B.n617 B.n616 585
R1072 B.n618 B.n617 585
R1073 B.n615 B.n378 585
R1074 B.n378 B.n377 585
R1075 B.n614 B.n613 585
R1076 B.n613 B.n612 585
R1077 B.n380 B.n379 585
R1078 B.n381 B.n380 585
R1079 B.n605 B.n604 585
R1080 B.n606 B.n605 585
R1081 B.n384 B.n383 585
R1082 B.n433 B.n431 585
R1083 B.n434 B.n430 585
R1084 B.n434 B.n385 585
R1085 B.n437 B.n436 585
R1086 B.n438 B.n429 585
R1087 B.n440 B.n439 585
R1088 B.n442 B.n428 585
R1089 B.n445 B.n444 585
R1090 B.n446 B.n427 585
R1091 B.n448 B.n447 585
R1092 B.n450 B.n426 585
R1093 B.n453 B.n452 585
R1094 B.n454 B.n425 585
R1095 B.n456 B.n455 585
R1096 B.n458 B.n424 585
R1097 B.n461 B.n460 585
R1098 B.n462 B.n423 585
R1099 B.n464 B.n463 585
R1100 B.n466 B.n422 585
R1101 B.n469 B.n468 585
R1102 B.n470 B.n421 585
R1103 B.n472 B.n471 585
R1104 B.n474 B.n420 585
R1105 B.n477 B.n476 585
R1106 B.n478 B.n419 585
R1107 B.n480 B.n479 585
R1108 B.n482 B.n418 585
R1109 B.n485 B.n484 585
R1110 B.n486 B.n417 585
R1111 B.n488 B.n487 585
R1112 B.n490 B.n416 585
R1113 B.n493 B.n492 585
R1114 B.n494 B.n415 585
R1115 B.n496 B.n495 585
R1116 B.n498 B.n414 585
R1117 B.n501 B.n500 585
R1118 B.n502 B.n413 585
R1119 B.n507 B.n506 585
R1120 B.n509 B.n412 585
R1121 B.n512 B.n511 585
R1122 B.n513 B.n411 585
R1123 B.n515 B.n514 585
R1124 B.n517 B.n410 585
R1125 B.n520 B.n519 585
R1126 B.n521 B.n409 585
R1127 B.n523 B.n522 585
R1128 B.n525 B.n408 585
R1129 B.n528 B.n527 585
R1130 B.n530 B.n405 585
R1131 B.n532 B.n531 585
R1132 B.n534 B.n404 585
R1133 B.n537 B.n536 585
R1134 B.n538 B.n403 585
R1135 B.n540 B.n539 585
R1136 B.n542 B.n402 585
R1137 B.n545 B.n544 585
R1138 B.n546 B.n401 585
R1139 B.n548 B.n547 585
R1140 B.n550 B.n400 585
R1141 B.n553 B.n552 585
R1142 B.n554 B.n399 585
R1143 B.n556 B.n555 585
R1144 B.n558 B.n398 585
R1145 B.n561 B.n560 585
R1146 B.n562 B.n397 585
R1147 B.n564 B.n563 585
R1148 B.n566 B.n396 585
R1149 B.n569 B.n568 585
R1150 B.n570 B.n395 585
R1151 B.n572 B.n571 585
R1152 B.n574 B.n394 585
R1153 B.n577 B.n576 585
R1154 B.n578 B.n393 585
R1155 B.n580 B.n579 585
R1156 B.n582 B.n392 585
R1157 B.n585 B.n584 585
R1158 B.n586 B.n391 585
R1159 B.n588 B.n587 585
R1160 B.n590 B.n390 585
R1161 B.n593 B.n592 585
R1162 B.n594 B.n389 585
R1163 B.n596 B.n595 585
R1164 B.n598 B.n388 585
R1165 B.n599 B.n387 585
R1166 B.n602 B.n601 585
R1167 B.n603 B.n386 585
R1168 B.n386 B.n385 585
R1169 B.n608 B.n607 585
R1170 B.n607 B.n606 585
R1171 B.n609 B.n382 585
R1172 B.n382 B.n381 585
R1173 B.n611 B.n610 585
R1174 B.n612 B.n611 585
R1175 B.n376 B.n375 585
R1176 B.n377 B.n376 585
R1177 B.n620 B.n619 585
R1178 B.n619 B.n618 585
R1179 B.n621 B.n374 585
R1180 B.n374 B.n373 585
R1181 B.n623 B.n622 585
R1182 B.n624 B.n623 585
R1183 B.n368 B.n367 585
R1184 B.n369 B.n368 585
R1185 B.n632 B.n631 585
R1186 B.n631 B.n630 585
R1187 B.n633 B.n366 585
R1188 B.n366 B.n365 585
R1189 B.n635 B.n634 585
R1190 B.n636 B.n635 585
R1191 B.n360 B.n359 585
R1192 B.n361 B.n360 585
R1193 B.n644 B.n643 585
R1194 B.n643 B.n642 585
R1195 B.n645 B.n358 585
R1196 B.n358 B.n357 585
R1197 B.n647 B.n646 585
R1198 B.n648 B.n647 585
R1199 B.n352 B.n351 585
R1200 B.n353 B.n352 585
R1201 B.n657 B.n656 585
R1202 B.n656 B.n655 585
R1203 B.n658 B.n350 585
R1204 B.n654 B.n350 585
R1205 B.n660 B.n659 585
R1206 B.n661 B.n660 585
R1207 B.n345 B.n344 585
R1208 B.n346 B.n345 585
R1209 B.n669 B.n668 585
R1210 B.n668 B.n667 585
R1211 B.n670 B.n343 585
R1212 B.n343 B.n342 585
R1213 B.n672 B.n671 585
R1214 B.n673 B.n672 585
R1215 B.n337 B.n336 585
R1216 B.n338 B.n337 585
R1217 B.n681 B.n680 585
R1218 B.n680 B.n679 585
R1219 B.n682 B.n335 585
R1220 B.n335 B.n334 585
R1221 B.n684 B.n683 585
R1222 B.n685 B.n684 585
R1223 B.n329 B.n328 585
R1224 B.n330 B.n329 585
R1225 B.n693 B.n692 585
R1226 B.n692 B.n691 585
R1227 B.n694 B.n327 585
R1228 B.n327 B.n325 585
R1229 B.n696 B.n695 585
R1230 B.n697 B.n696 585
R1231 B.n321 B.n320 585
R1232 B.n326 B.n321 585
R1233 B.n705 B.n704 585
R1234 B.n704 B.n703 585
R1235 B.n706 B.n319 585
R1236 B.n319 B.n318 585
R1237 B.n708 B.n707 585
R1238 B.n709 B.n708 585
R1239 B.n313 B.n312 585
R1240 B.n314 B.n313 585
R1241 B.n717 B.n716 585
R1242 B.n716 B.n715 585
R1243 B.n718 B.n311 585
R1244 B.n311 B.n309 585
R1245 B.n720 B.n719 585
R1246 B.n721 B.n720 585
R1247 B.n305 B.n304 585
R1248 B.n310 B.n305 585
R1249 B.n730 B.n729 585
R1250 B.n729 B.n728 585
R1251 B.n731 B.n303 585
R1252 B.n303 B.n302 585
R1253 B.n733 B.n732 585
R1254 B.n734 B.n733 585
R1255 B.n3 B.n0 585
R1256 B.n4 B.n3 585
R1257 B.n886 B.n1 585
R1258 B.n887 B.n886 585
R1259 B.n885 B.n884 585
R1260 B.n885 B.n8 585
R1261 B.n883 B.n9 585
R1262 B.n12 B.n9 585
R1263 B.n882 B.n881 585
R1264 B.n881 B.n880 585
R1265 B.n11 B.n10 585
R1266 B.n879 B.n11 585
R1267 B.n877 B.n876 585
R1268 B.n878 B.n877 585
R1269 B.n875 B.n17 585
R1270 B.n17 B.n16 585
R1271 B.n874 B.n873 585
R1272 B.n873 B.n872 585
R1273 B.n19 B.n18 585
R1274 B.n871 B.n19 585
R1275 B.n869 B.n868 585
R1276 B.n870 B.n869 585
R1277 B.n867 B.n24 585
R1278 B.n24 B.n23 585
R1279 B.n866 B.n865 585
R1280 B.n865 B.n864 585
R1281 B.n26 B.n25 585
R1282 B.n863 B.n26 585
R1283 B.n861 B.n860 585
R1284 B.n862 B.n861 585
R1285 B.n859 B.n31 585
R1286 B.n31 B.n30 585
R1287 B.n858 B.n857 585
R1288 B.n857 B.n856 585
R1289 B.n33 B.n32 585
R1290 B.n855 B.n33 585
R1291 B.n853 B.n852 585
R1292 B.n854 B.n853 585
R1293 B.n851 B.n38 585
R1294 B.n38 B.n37 585
R1295 B.n850 B.n849 585
R1296 B.n849 B.n848 585
R1297 B.n40 B.n39 585
R1298 B.n847 B.n40 585
R1299 B.n845 B.n844 585
R1300 B.n846 B.n845 585
R1301 B.n843 B.n45 585
R1302 B.n45 B.n44 585
R1303 B.n842 B.n841 585
R1304 B.n841 B.n840 585
R1305 B.n47 B.n46 585
R1306 B.n839 B.n47 585
R1307 B.n837 B.n836 585
R1308 B.n838 B.n837 585
R1309 B.n835 B.n51 585
R1310 B.n54 B.n51 585
R1311 B.n834 B.n833 585
R1312 B.n833 B.n832 585
R1313 B.n53 B.n52 585
R1314 B.n831 B.n53 585
R1315 B.n829 B.n828 585
R1316 B.n830 B.n829 585
R1317 B.n827 B.n59 585
R1318 B.n59 B.n58 585
R1319 B.n826 B.n825 585
R1320 B.n825 B.n824 585
R1321 B.n61 B.n60 585
R1322 B.n823 B.n61 585
R1323 B.n821 B.n820 585
R1324 B.n822 B.n821 585
R1325 B.n819 B.n66 585
R1326 B.n66 B.n65 585
R1327 B.n818 B.n817 585
R1328 B.n817 B.n816 585
R1329 B.n68 B.n67 585
R1330 B.n815 B.n68 585
R1331 B.n813 B.n812 585
R1332 B.n814 B.n813 585
R1333 B.n811 B.n73 585
R1334 B.n73 B.n72 585
R1335 B.n810 B.n809 585
R1336 B.n809 B.n808 585
R1337 B.n75 B.n74 585
R1338 B.n807 B.n75 585
R1339 B.n805 B.n804 585
R1340 B.n806 B.n805 585
R1341 B.n803 B.n80 585
R1342 B.n80 B.n79 585
R1343 B.n802 B.n801 585
R1344 B.n801 B.n800 585
R1345 B.n890 B.n889 585
R1346 B.n888 B.n2 585
R1347 B.n801 B.n82 530.939
R1348 B.n797 B.n83 530.939
R1349 B.n605 B.n386 530.939
R1350 B.n607 B.n384 530.939
R1351 B.n130 B.t8 328.104
R1352 B.n127 B.t19 328.104
R1353 B.n406 B.t16 328.104
R1354 B.n503 B.t12 328.104
R1355 B.n127 B.t20 310.56
R1356 B.n406 B.t18 310.56
R1357 B.n130 B.t10 310.56
R1358 B.n503 B.t15 310.56
R1359 B.n128 B.t21 262.269
R1360 B.n407 B.t17 262.269
R1361 B.n131 B.t11 262.269
R1362 B.n504 B.t14 262.269
R1363 B.n799 B.n798 256.663
R1364 B.n799 B.n125 256.663
R1365 B.n799 B.n124 256.663
R1366 B.n799 B.n123 256.663
R1367 B.n799 B.n122 256.663
R1368 B.n799 B.n121 256.663
R1369 B.n799 B.n120 256.663
R1370 B.n799 B.n119 256.663
R1371 B.n799 B.n118 256.663
R1372 B.n799 B.n117 256.663
R1373 B.n799 B.n116 256.663
R1374 B.n799 B.n115 256.663
R1375 B.n799 B.n114 256.663
R1376 B.n799 B.n113 256.663
R1377 B.n799 B.n112 256.663
R1378 B.n799 B.n111 256.663
R1379 B.n799 B.n110 256.663
R1380 B.n799 B.n109 256.663
R1381 B.n799 B.n108 256.663
R1382 B.n799 B.n107 256.663
R1383 B.n799 B.n106 256.663
R1384 B.n799 B.n105 256.663
R1385 B.n799 B.n104 256.663
R1386 B.n799 B.n103 256.663
R1387 B.n799 B.n102 256.663
R1388 B.n799 B.n101 256.663
R1389 B.n799 B.n100 256.663
R1390 B.n799 B.n99 256.663
R1391 B.n799 B.n98 256.663
R1392 B.n799 B.n97 256.663
R1393 B.n799 B.n96 256.663
R1394 B.n799 B.n95 256.663
R1395 B.n799 B.n94 256.663
R1396 B.n799 B.n93 256.663
R1397 B.n799 B.n92 256.663
R1398 B.n799 B.n91 256.663
R1399 B.n799 B.n90 256.663
R1400 B.n799 B.n89 256.663
R1401 B.n799 B.n88 256.663
R1402 B.n799 B.n87 256.663
R1403 B.n799 B.n86 256.663
R1404 B.n799 B.n85 256.663
R1405 B.n799 B.n84 256.663
R1406 B.n432 B.n385 256.663
R1407 B.n435 B.n385 256.663
R1408 B.n441 B.n385 256.663
R1409 B.n443 B.n385 256.663
R1410 B.n449 B.n385 256.663
R1411 B.n451 B.n385 256.663
R1412 B.n457 B.n385 256.663
R1413 B.n459 B.n385 256.663
R1414 B.n465 B.n385 256.663
R1415 B.n467 B.n385 256.663
R1416 B.n473 B.n385 256.663
R1417 B.n475 B.n385 256.663
R1418 B.n481 B.n385 256.663
R1419 B.n483 B.n385 256.663
R1420 B.n489 B.n385 256.663
R1421 B.n491 B.n385 256.663
R1422 B.n497 B.n385 256.663
R1423 B.n499 B.n385 256.663
R1424 B.n508 B.n385 256.663
R1425 B.n510 B.n385 256.663
R1426 B.n516 B.n385 256.663
R1427 B.n518 B.n385 256.663
R1428 B.n524 B.n385 256.663
R1429 B.n526 B.n385 256.663
R1430 B.n533 B.n385 256.663
R1431 B.n535 B.n385 256.663
R1432 B.n541 B.n385 256.663
R1433 B.n543 B.n385 256.663
R1434 B.n549 B.n385 256.663
R1435 B.n551 B.n385 256.663
R1436 B.n557 B.n385 256.663
R1437 B.n559 B.n385 256.663
R1438 B.n565 B.n385 256.663
R1439 B.n567 B.n385 256.663
R1440 B.n573 B.n385 256.663
R1441 B.n575 B.n385 256.663
R1442 B.n581 B.n385 256.663
R1443 B.n583 B.n385 256.663
R1444 B.n589 B.n385 256.663
R1445 B.n591 B.n385 256.663
R1446 B.n597 B.n385 256.663
R1447 B.n600 B.n385 256.663
R1448 B.n892 B.n891 256.663
R1449 B.n135 B.n134 163.367
R1450 B.n139 B.n138 163.367
R1451 B.n143 B.n142 163.367
R1452 B.n147 B.n146 163.367
R1453 B.n151 B.n150 163.367
R1454 B.n155 B.n154 163.367
R1455 B.n159 B.n158 163.367
R1456 B.n163 B.n162 163.367
R1457 B.n167 B.n166 163.367
R1458 B.n171 B.n170 163.367
R1459 B.n175 B.n174 163.367
R1460 B.n179 B.n178 163.367
R1461 B.n183 B.n182 163.367
R1462 B.n187 B.n186 163.367
R1463 B.n191 B.n190 163.367
R1464 B.n195 B.n194 163.367
R1465 B.n199 B.n198 163.367
R1466 B.n203 B.n202 163.367
R1467 B.n207 B.n206 163.367
R1468 B.n211 B.n210 163.367
R1469 B.n215 B.n214 163.367
R1470 B.n219 B.n218 163.367
R1471 B.n223 B.n222 163.367
R1472 B.n227 B.n226 163.367
R1473 B.n231 B.n230 163.367
R1474 B.n235 B.n234 163.367
R1475 B.n239 B.n238 163.367
R1476 B.n243 B.n242 163.367
R1477 B.n247 B.n246 163.367
R1478 B.n251 B.n250 163.367
R1479 B.n255 B.n254 163.367
R1480 B.n259 B.n258 163.367
R1481 B.n263 B.n262 163.367
R1482 B.n267 B.n266 163.367
R1483 B.n271 B.n270 163.367
R1484 B.n275 B.n274 163.367
R1485 B.n279 B.n278 163.367
R1486 B.n283 B.n282 163.367
R1487 B.n287 B.n286 163.367
R1488 B.n291 B.n290 163.367
R1489 B.n295 B.n294 163.367
R1490 B.n297 B.n126 163.367
R1491 B.n605 B.n380 163.367
R1492 B.n613 B.n380 163.367
R1493 B.n613 B.n378 163.367
R1494 B.n617 B.n378 163.367
R1495 B.n617 B.n372 163.367
R1496 B.n625 B.n372 163.367
R1497 B.n625 B.n370 163.367
R1498 B.n629 B.n370 163.367
R1499 B.n629 B.n364 163.367
R1500 B.n637 B.n364 163.367
R1501 B.n637 B.n362 163.367
R1502 B.n641 B.n362 163.367
R1503 B.n641 B.n356 163.367
R1504 B.n649 B.n356 163.367
R1505 B.n649 B.n354 163.367
R1506 B.n653 B.n354 163.367
R1507 B.n653 B.n349 163.367
R1508 B.n662 B.n349 163.367
R1509 B.n662 B.n347 163.367
R1510 B.n666 B.n347 163.367
R1511 B.n666 B.n341 163.367
R1512 B.n674 B.n341 163.367
R1513 B.n674 B.n339 163.367
R1514 B.n678 B.n339 163.367
R1515 B.n678 B.n333 163.367
R1516 B.n686 B.n333 163.367
R1517 B.n686 B.n331 163.367
R1518 B.n690 B.n331 163.367
R1519 B.n690 B.n324 163.367
R1520 B.n698 B.n324 163.367
R1521 B.n698 B.n322 163.367
R1522 B.n702 B.n322 163.367
R1523 B.n702 B.n317 163.367
R1524 B.n710 B.n317 163.367
R1525 B.n710 B.n315 163.367
R1526 B.n714 B.n315 163.367
R1527 B.n714 B.n308 163.367
R1528 B.n722 B.n308 163.367
R1529 B.n722 B.n306 163.367
R1530 B.n727 B.n306 163.367
R1531 B.n727 B.n301 163.367
R1532 B.n735 B.n301 163.367
R1533 B.n736 B.n735 163.367
R1534 B.n736 B.n5 163.367
R1535 B.n6 B.n5 163.367
R1536 B.n7 B.n6 163.367
R1537 B.n742 B.n7 163.367
R1538 B.n743 B.n742 163.367
R1539 B.n743 B.n13 163.367
R1540 B.n14 B.n13 163.367
R1541 B.n15 B.n14 163.367
R1542 B.n748 B.n15 163.367
R1543 B.n748 B.n20 163.367
R1544 B.n21 B.n20 163.367
R1545 B.n22 B.n21 163.367
R1546 B.n753 B.n22 163.367
R1547 B.n753 B.n27 163.367
R1548 B.n28 B.n27 163.367
R1549 B.n29 B.n28 163.367
R1550 B.n758 B.n29 163.367
R1551 B.n758 B.n34 163.367
R1552 B.n35 B.n34 163.367
R1553 B.n36 B.n35 163.367
R1554 B.n763 B.n36 163.367
R1555 B.n763 B.n41 163.367
R1556 B.n42 B.n41 163.367
R1557 B.n43 B.n42 163.367
R1558 B.n768 B.n43 163.367
R1559 B.n768 B.n48 163.367
R1560 B.n49 B.n48 163.367
R1561 B.n50 B.n49 163.367
R1562 B.n773 B.n50 163.367
R1563 B.n773 B.n55 163.367
R1564 B.n56 B.n55 163.367
R1565 B.n57 B.n56 163.367
R1566 B.n778 B.n57 163.367
R1567 B.n778 B.n62 163.367
R1568 B.n63 B.n62 163.367
R1569 B.n64 B.n63 163.367
R1570 B.n783 B.n64 163.367
R1571 B.n783 B.n69 163.367
R1572 B.n70 B.n69 163.367
R1573 B.n71 B.n70 163.367
R1574 B.n788 B.n71 163.367
R1575 B.n788 B.n76 163.367
R1576 B.n77 B.n76 163.367
R1577 B.n78 B.n77 163.367
R1578 B.n793 B.n78 163.367
R1579 B.n793 B.n83 163.367
R1580 B.n434 B.n433 163.367
R1581 B.n436 B.n434 163.367
R1582 B.n440 B.n429 163.367
R1583 B.n444 B.n442 163.367
R1584 B.n448 B.n427 163.367
R1585 B.n452 B.n450 163.367
R1586 B.n456 B.n425 163.367
R1587 B.n460 B.n458 163.367
R1588 B.n464 B.n423 163.367
R1589 B.n468 B.n466 163.367
R1590 B.n472 B.n421 163.367
R1591 B.n476 B.n474 163.367
R1592 B.n480 B.n419 163.367
R1593 B.n484 B.n482 163.367
R1594 B.n488 B.n417 163.367
R1595 B.n492 B.n490 163.367
R1596 B.n496 B.n415 163.367
R1597 B.n500 B.n498 163.367
R1598 B.n507 B.n413 163.367
R1599 B.n511 B.n509 163.367
R1600 B.n515 B.n411 163.367
R1601 B.n519 B.n517 163.367
R1602 B.n523 B.n409 163.367
R1603 B.n527 B.n525 163.367
R1604 B.n532 B.n405 163.367
R1605 B.n536 B.n534 163.367
R1606 B.n540 B.n403 163.367
R1607 B.n544 B.n542 163.367
R1608 B.n548 B.n401 163.367
R1609 B.n552 B.n550 163.367
R1610 B.n556 B.n399 163.367
R1611 B.n560 B.n558 163.367
R1612 B.n564 B.n397 163.367
R1613 B.n568 B.n566 163.367
R1614 B.n572 B.n395 163.367
R1615 B.n576 B.n574 163.367
R1616 B.n580 B.n393 163.367
R1617 B.n584 B.n582 163.367
R1618 B.n588 B.n391 163.367
R1619 B.n592 B.n590 163.367
R1620 B.n596 B.n389 163.367
R1621 B.n599 B.n598 163.367
R1622 B.n601 B.n386 163.367
R1623 B.n607 B.n382 163.367
R1624 B.n611 B.n382 163.367
R1625 B.n611 B.n376 163.367
R1626 B.n619 B.n376 163.367
R1627 B.n619 B.n374 163.367
R1628 B.n623 B.n374 163.367
R1629 B.n623 B.n368 163.367
R1630 B.n631 B.n368 163.367
R1631 B.n631 B.n366 163.367
R1632 B.n635 B.n366 163.367
R1633 B.n635 B.n360 163.367
R1634 B.n643 B.n360 163.367
R1635 B.n643 B.n358 163.367
R1636 B.n647 B.n358 163.367
R1637 B.n647 B.n352 163.367
R1638 B.n656 B.n352 163.367
R1639 B.n656 B.n350 163.367
R1640 B.n660 B.n350 163.367
R1641 B.n660 B.n345 163.367
R1642 B.n668 B.n345 163.367
R1643 B.n668 B.n343 163.367
R1644 B.n672 B.n343 163.367
R1645 B.n672 B.n337 163.367
R1646 B.n680 B.n337 163.367
R1647 B.n680 B.n335 163.367
R1648 B.n684 B.n335 163.367
R1649 B.n684 B.n329 163.367
R1650 B.n692 B.n329 163.367
R1651 B.n692 B.n327 163.367
R1652 B.n696 B.n327 163.367
R1653 B.n696 B.n321 163.367
R1654 B.n704 B.n321 163.367
R1655 B.n704 B.n319 163.367
R1656 B.n708 B.n319 163.367
R1657 B.n708 B.n313 163.367
R1658 B.n716 B.n313 163.367
R1659 B.n716 B.n311 163.367
R1660 B.n720 B.n311 163.367
R1661 B.n720 B.n305 163.367
R1662 B.n729 B.n305 163.367
R1663 B.n729 B.n303 163.367
R1664 B.n733 B.n303 163.367
R1665 B.n733 B.n3 163.367
R1666 B.n890 B.n3 163.367
R1667 B.n886 B.n2 163.367
R1668 B.n886 B.n885 163.367
R1669 B.n885 B.n9 163.367
R1670 B.n881 B.n9 163.367
R1671 B.n881 B.n11 163.367
R1672 B.n877 B.n11 163.367
R1673 B.n877 B.n17 163.367
R1674 B.n873 B.n17 163.367
R1675 B.n873 B.n19 163.367
R1676 B.n869 B.n19 163.367
R1677 B.n869 B.n24 163.367
R1678 B.n865 B.n24 163.367
R1679 B.n865 B.n26 163.367
R1680 B.n861 B.n26 163.367
R1681 B.n861 B.n31 163.367
R1682 B.n857 B.n31 163.367
R1683 B.n857 B.n33 163.367
R1684 B.n853 B.n33 163.367
R1685 B.n853 B.n38 163.367
R1686 B.n849 B.n38 163.367
R1687 B.n849 B.n40 163.367
R1688 B.n845 B.n40 163.367
R1689 B.n845 B.n45 163.367
R1690 B.n841 B.n45 163.367
R1691 B.n841 B.n47 163.367
R1692 B.n837 B.n47 163.367
R1693 B.n837 B.n51 163.367
R1694 B.n833 B.n51 163.367
R1695 B.n833 B.n53 163.367
R1696 B.n829 B.n53 163.367
R1697 B.n829 B.n59 163.367
R1698 B.n825 B.n59 163.367
R1699 B.n825 B.n61 163.367
R1700 B.n821 B.n61 163.367
R1701 B.n821 B.n66 163.367
R1702 B.n817 B.n66 163.367
R1703 B.n817 B.n68 163.367
R1704 B.n813 B.n68 163.367
R1705 B.n813 B.n73 163.367
R1706 B.n809 B.n73 163.367
R1707 B.n809 B.n75 163.367
R1708 B.n805 B.n75 163.367
R1709 B.n805 B.n80 163.367
R1710 B.n801 B.n80 163.367
R1711 B.n606 B.n385 94.94
R1712 B.n800 B.n799 94.94
R1713 B.n84 B.n82 71.676
R1714 B.n135 B.n85 71.676
R1715 B.n139 B.n86 71.676
R1716 B.n143 B.n87 71.676
R1717 B.n147 B.n88 71.676
R1718 B.n151 B.n89 71.676
R1719 B.n155 B.n90 71.676
R1720 B.n159 B.n91 71.676
R1721 B.n163 B.n92 71.676
R1722 B.n167 B.n93 71.676
R1723 B.n171 B.n94 71.676
R1724 B.n175 B.n95 71.676
R1725 B.n179 B.n96 71.676
R1726 B.n183 B.n97 71.676
R1727 B.n187 B.n98 71.676
R1728 B.n191 B.n99 71.676
R1729 B.n195 B.n100 71.676
R1730 B.n199 B.n101 71.676
R1731 B.n203 B.n102 71.676
R1732 B.n207 B.n103 71.676
R1733 B.n211 B.n104 71.676
R1734 B.n215 B.n105 71.676
R1735 B.n219 B.n106 71.676
R1736 B.n223 B.n107 71.676
R1737 B.n227 B.n108 71.676
R1738 B.n231 B.n109 71.676
R1739 B.n235 B.n110 71.676
R1740 B.n239 B.n111 71.676
R1741 B.n243 B.n112 71.676
R1742 B.n247 B.n113 71.676
R1743 B.n251 B.n114 71.676
R1744 B.n255 B.n115 71.676
R1745 B.n259 B.n116 71.676
R1746 B.n263 B.n117 71.676
R1747 B.n267 B.n118 71.676
R1748 B.n271 B.n119 71.676
R1749 B.n275 B.n120 71.676
R1750 B.n279 B.n121 71.676
R1751 B.n283 B.n122 71.676
R1752 B.n287 B.n123 71.676
R1753 B.n291 B.n124 71.676
R1754 B.n295 B.n125 71.676
R1755 B.n798 B.n126 71.676
R1756 B.n798 B.n797 71.676
R1757 B.n297 B.n125 71.676
R1758 B.n294 B.n124 71.676
R1759 B.n290 B.n123 71.676
R1760 B.n286 B.n122 71.676
R1761 B.n282 B.n121 71.676
R1762 B.n278 B.n120 71.676
R1763 B.n274 B.n119 71.676
R1764 B.n270 B.n118 71.676
R1765 B.n266 B.n117 71.676
R1766 B.n262 B.n116 71.676
R1767 B.n258 B.n115 71.676
R1768 B.n254 B.n114 71.676
R1769 B.n250 B.n113 71.676
R1770 B.n246 B.n112 71.676
R1771 B.n242 B.n111 71.676
R1772 B.n238 B.n110 71.676
R1773 B.n234 B.n109 71.676
R1774 B.n230 B.n108 71.676
R1775 B.n226 B.n107 71.676
R1776 B.n222 B.n106 71.676
R1777 B.n218 B.n105 71.676
R1778 B.n214 B.n104 71.676
R1779 B.n210 B.n103 71.676
R1780 B.n206 B.n102 71.676
R1781 B.n202 B.n101 71.676
R1782 B.n198 B.n100 71.676
R1783 B.n194 B.n99 71.676
R1784 B.n190 B.n98 71.676
R1785 B.n186 B.n97 71.676
R1786 B.n182 B.n96 71.676
R1787 B.n178 B.n95 71.676
R1788 B.n174 B.n94 71.676
R1789 B.n170 B.n93 71.676
R1790 B.n166 B.n92 71.676
R1791 B.n162 B.n91 71.676
R1792 B.n158 B.n90 71.676
R1793 B.n154 B.n89 71.676
R1794 B.n150 B.n88 71.676
R1795 B.n146 B.n87 71.676
R1796 B.n142 B.n86 71.676
R1797 B.n138 B.n85 71.676
R1798 B.n134 B.n84 71.676
R1799 B.n432 B.n384 71.676
R1800 B.n436 B.n435 71.676
R1801 B.n441 B.n440 71.676
R1802 B.n444 B.n443 71.676
R1803 B.n449 B.n448 71.676
R1804 B.n452 B.n451 71.676
R1805 B.n457 B.n456 71.676
R1806 B.n460 B.n459 71.676
R1807 B.n465 B.n464 71.676
R1808 B.n468 B.n467 71.676
R1809 B.n473 B.n472 71.676
R1810 B.n476 B.n475 71.676
R1811 B.n481 B.n480 71.676
R1812 B.n484 B.n483 71.676
R1813 B.n489 B.n488 71.676
R1814 B.n492 B.n491 71.676
R1815 B.n497 B.n496 71.676
R1816 B.n500 B.n499 71.676
R1817 B.n508 B.n507 71.676
R1818 B.n511 B.n510 71.676
R1819 B.n516 B.n515 71.676
R1820 B.n519 B.n518 71.676
R1821 B.n524 B.n523 71.676
R1822 B.n527 B.n526 71.676
R1823 B.n533 B.n532 71.676
R1824 B.n536 B.n535 71.676
R1825 B.n541 B.n540 71.676
R1826 B.n544 B.n543 71.676
R1827 B.n549 B.n548 71.676
R1828 B.n552 B.n551 71.676
R1829 B.n557 B.n556 71.676
R1830 B.n560 B.n559 71.676
R1831 B.n565 B.n564 71.676
R1832 B.n568 B.n567 71.676
R1833 B.n573 B.n572 71.676
R1834 B.n576 B.n575 71.676
R1835 B.n581 B.n580 71.676
R1836 B.n584 B.n583 71.676
R1837 B.n589 B.n588 71.676
R1838 B.n592 B.n591 71.676
R1839 B.n597 B.n596 71.676
R1840 B.n600 B.n599 71.676
R1841 B.n433 B.n432 71.676
R1842 B.n435 B.n429 71.676
R1843 B.n442 B.n441 71.676
R1844 B.n443 B.n427 71.676
R1845 B.n450 B.n449 71.676
R1846 B.n451 B.n425 71.676
R1847 B.n458 B.n457 71.676
R1848 B.n459 B.n423 71.676
R1849 B.n466 B.n465 71.676
R1850 B.n467 B.n421 71.676
R1851 B.n474 B.n473 71.676
R1852 B.n475 B.n419 71.676
R1853 B.n482 B.n481 71.676
R1854 B.n483 B.n417 71.676
R1855 B.n490 B.n489 71.676
R1856 B.n491 B.n415 71.676
R1857 B.n498 B.n497 71.676
R1858 B.n499 B.n413 71.676
R1859 B.n509 B.n508 71.676
R1860 B.n510 B.n411 71.676
R1861 B.n517 B.n516 71.676
R1862 B.n518 B.n409 71.676
R1863 B.n525 B.n524 71.676
R1864 B.n526 B.n405 71.676
R1865 B.n534 B.n533 71.676
R1866 B.n535 B.n403 71.676
R1867 B.n542 B.n541 71.676
R1868 B.n543 B.n401 71.676
R1869 B.n550 B.n549 71.676
R1870 B.n551 B.n399 71.676
R1871 B.n558 B.n557 71.676
R1872 B.n559 B.n397 71.676
R1873 B.n566 B.n565 71.676
R1874 B.n567 B.n395 71.676
R1875 B.n574 B.n573 71.676
R1876 B.n575 B.n393 71.676
R1877 B.n582 B.n581 71.676
R1878 B.n583 B.n391 71.676
R1879 B.n590 B.n589 71.676
R1880 B.n591 B.n389 71.676
R1881 B.n598 B.n597 71.676
R1882 B.n601 B.n600 71.676
R1883 B.n891 B.n890 71.676
R1884 B.n891 B.n2 71.676
R1885 B.n132 B.n131 59.5399
R1886 B.n129 B.n128 59.5399
R1887 B.n529 B.n407 59.5399
R1888 B.n505 B.n504 59.5399
R1889 B.n131 B.n130 48.2914
R1890 B.n128 B.n127 48.2914
R1891 B.n407 B.n406 48.2914
R1892 B.n504 B.n503 48.2914
R1893 B.n606 B.n381 46.4457
R1894 B.n612 B.n381 46.4457
R1895 B.n612 B.n377 46.4457
R1896 B.n618 B.n377 46.4457
R1897 B.n618 B.n373 46.4457
R1898 B.n624 B.n373 46.4457
R1899 B.n630 B.n369 46.4457
R1900 B.n630 B.n365 46.4457
R1901 B.n636 B.n365 46.4457
R1902 B.n636 B.n361 46.4457
R1903 B.n642 B.n361 46.4457
R1904 B.n642 B.n357 46.4457
R1905 B.n648 B.n357 46.4457
R1906 B.n648 B.n353 46.4457
R1907 B.n655 B.n353 46.4457
R1908 B.n655 B.n654 46.4457
R1909 B.n661 B.n346 46.4457
R1910 B.n667 B.n346 46.4457
R1911 B.n667 B.n342 46.4457
R1912 B.n673 B.n342 46.4457
R1913 B.n673 B.n338 46.4457
R1914 B.n679 B.n338 46.4457
R1915 B.n685 B.n334 46.4457
R1916 B.n685 B.n330 46.4457
R1917 B.n691 B.n330 46.4457
R1918 B.n691 B.n325 46.4457
R1919 B.n697 B.n325 46.4457
R1920 B.n697 B.n326 46.4457
R1921 B.n703 B.n318 46.4457
R1922 B.n709 B.n318 46.4457
R1923 B.n709 B.n314 46.4457
R1924 B.n715 B.n314 46.4457
R1925 B.n715 B.n309 46.4457
R1926 B.n721 B.n309 46.4457
R1927 B.n721 B.n310 46.4457
R1928 B.n728 B.n302 46.4457
R1929 B.n734 B.n302 46.4457
R1930 B.n734 B.n4 46.4457
R1931 B.n889 B.n4 46.4457
R1932 B.n889 B.n888 46.4457
R1933 B.n888 B.n887 46.4457
R1934 B.n887 B.n8 46.4457
R1935 B.n12 B.n8 46.4457
R1936 B.n880 B.n12 46.4457
R1937 B.n879 B.n878 46.4457
R1938 B.n878 B.n16 46.4457
R1939 B.n872 B.n16 46.4457
R1940 B.n872 B.n871 46.4457
R1941 B.n871 B.n870 46.4457
R1942 B.n870 B.n23 46.4457
R1943 B.n864 B.n23 46.4457
R1944 B.n863 B.n862 46.4457
R1945 B.n862 B.n30 46.4457
R1946 B.n856 B.n30 46.4457
R1947 B.n856 B.n855 46.4457
R1948 B.n855 B.n854 46.4457
R1949 B.n854 B.n37 46.4457
R1950 B.n848 B.n847 46.4457
R1951 B.n847 B.n846 46.4457
R1952 B.n846 B.n44 46.4457
R1953 B.n840 B.n44 46.4457
R1954 B.n840 B.n839 46.4457
R1955 B.n839 B.n838 46.4457
R1956 B.n832 B.n54 46.4457
R1957 B.n832 B.n831 46.4457
R1958 B.n831 B.n830 46.4457
R1959 B.n830 B.n58 46.4457
R1960 B.n824 B.n58 46.4457
R1961 B.n824 B.n823 46.4457
R1962 B.n823 B.n822 46.4457
R1963 B.n822 B.n65 46.4457
R1964 B.n816 B.n65 46.4457
R1965 B.n816 B.n815 46.4457
R1966 B.n814 B.n72 46.4457
R1967 B.n808 B.n72 46.4457
R1968 B.n808 B.n807 46.4457
R1969 B.n807 B.n806 46.4457
R1970 B.n806 B.n79 46.4457
R1971 B.n800 B.n79 46.4457
R1972 B.n326 B.t6 42.3476
R1973 B.t3 B.n863 42.3476
R1974 B.n728 B.t2 35.5174
R1975 B.n880 B.t4 35.5174
R1976 B.n608 B.n383 34.4981
R1977 B.n604 B.n603 34.4981
R1978 B.n796 B.n795 34.4981
R1979 B.n802 B.n81 34.4981
R1980 B.n624 B.t13 34.1514
R1981 B.n661 B.t0 34.1514
R1982 B.n838 B.t1 34.1514
R1983 B.t9 B.n814 34.1514
R1984 B.n679 B.t5 27.3212
R1985 B.n848 B.t7 27.3212
R1986 B.t5 B.n334 19.125
R1987 B.t7 B.n37 19.125
R1988 B B.n892 18.0485
R1989 B.t13 B.n369 12.2948
R1990 B.n654 B.t0 12.2948
R1991 B.n54 B.t1 12.2948
R1992 B.n815 B.t9 12.2948
R1993 B.n310 B.t2 10.9288
R1994 B.t4 B.n879 10.9288
R1995 B.n609 B.n608 10.6151
R1996 B.n610 B.n609 10.6151
R1997 B.n610 B.n375 10.6151
R1998 B.n620 B.n375 10.6151
R1999 B.n621 B.n620 10.6151
R2000 B.n622 B.n621 10.6151
R2001 B.n622 B.n367 10.6151
R2002 B.n632 B.n367 10.6151
R2003 B.n633 B.n632 10.6151
R2004 B.n634 B.n633 10.6151
R2005 B.n634 B.n359 10.6151
R2006 B.n644 B.n359 10.6151
R2007 B.n645 B.n644 10.6151
R2008 B.n646 B.n645 10.6151
R2009 B.n646 B.n351 10.6151
R2010 B.n657 B.n351 10.6151
R2011 B.n658 B.n657 10.6151
R2012 B.n659 B.n658 10.6151
R2013 B.n659 B.n344 10.6151
R2014 B.n669 B.n344 10.6151
R2015 B.n670 B.n669 10.6151
R2016 B.n671 B.n670 10.6151
R2017 B.n671 B.n336 10.6151
R2018 B.n681 B.n336 10.6151
R2019 B.n682 B.n681 10.6151
R2020 B.n683 B.n682 10.6151
R2021 B.n683 B.n328 10.6151
R2022 B.n693 B.n328 10.6151
R2023 B.n694 B.n693 10.6151
R2024 B.n695 B.n694 10.6151
R2025 B.n695 B.n320 10.6151
R2026 B.n705 B.n320 10.6151
R2027 B.n706 B.n705 10.6151
R2028 B.n707 B.n706 10.6151
R2029 B.n707 B.n312 10.6151
R2030 B.n717 B.n312 10.6151
R2031 B.n718 B.n717 10.6151
R2032 B.n719 B.n718 10.6151
R2033 B.n719 B.n304 10.6151
R2034 B.n730 B.n304 10.6151
R2035 B.n731 B.n730 10.6151
R2036 B.n732 B.n731 10.6151
R2037 B.n732 B.n0 10.6151
R2038 B.n431 B.n383 10.6151
R2039 B.n431 B.n430 10.6151
R2040 B.n437 B.n430 10.6151
R2041 B.n438 B.n437 10.6151
R2042 B.n439 B.n438 10.6151
R2043 B.n439 B.n428 10.6151
R2044 B.n445 B.n428 10.6151
R2045 B.n446 B.n445 10.6151
R2046 B.n447 B.n446 10.6151
R2047 B.n447 B.n426 10.6151
R2048 B.n453 B.n426 10.6151
R2049 B.n454 B.n453 10.6151
R2050 B.n455 B.n454 10.6151
R2051 B.n455 B.n424 10.6151
R2052 B.n461 B.n424 10.6151
R2053 B.n462 B.n461 10.6151
R2054 B.n463 B.n462 10.6151
R2055 B.n463 B.n422 10.6151
R2056 B.n469 B.n422 10.6151
R2057 B.n470 B.n469 10.6151
R2058 B.n471 B.n470 10.6151
R2059 B.n471 B.n420 10.6151
R2060 B.n477 B.n420 10.6151
R2061 B.n478 B.n477 10.6151
R2062 B.n479 B.n478 10.6151
R2063 B.n479 B.n418 10.6151
R2064 B.n485 B.n418 10.6151
R2065 B.n486 B.n485 10.6151
R2066 B.n487 B.n486 10.6151
R2067 B.n487 B.n416 10.6151
R2068 B.n493 B.n416 10.6151
R2069 B.n494 B.n493 10.6151
R2070 B.n495 B.n494 10.6151
R2071 B.n495 B.n414 10.6151
R2072 B.n501 B.n414 10.6151
R2073 B.n502 B.n501 10.6151
R2074 B.n506 B.n502 10.6151
R2075 B.n512 B.n412 10.6151
R2076 B.n513 B.n512 10.6151
R2077 B.n514 B.n513 10.6151
R2078 B.n514 B.n410 10.6151
R2079 B.n520 B.n410 10.6151
R2080 B.n521 B.n520 10.6151
R2081 B.n522 B.n521 10.6151
R2082 B.n522 B.n408 10.6151
R2083 B.n528 B.n408 10.6151
R2084 B.n531 B.n530 10.6151
R2085 B.n531 B.n404 10.6151
R2086 B.n537 B.n404 10.6151
R2087 B.n538 B.n537 10.6151
R2088 B.n539 B.n538 10.6151
R2089 B.n539 B.n402 10.6151
R2090 B.n545 B.n402 10.6151
R2091 B.n546 B.n545 10.6151
R2092 B.n547 B.n546 10.6151
R2093 B.n547 B.n400 10.6151
R2094 B.n553 B.n400 10.6151
R2095 B.n554 B.n553 10.6151
R2096 B.n555 B.n554 10.6151
R2097 B.n555 B.n398 10.6151
R2098 B.n561 B.n398 10.6151
R2099 B.n562 B.n561 10.6151
R2100 B.n563 B.n562 10.6151
R2101 B.n563 B.n396 10.6151
R2102 B.n569 B.n396 10.6151
R2103 B.n570 B.n569 10.6151
R2104 B.n571 B.n570 10.6151
R2105 B.n571 B.n394 10.6151
R2106 B.n577 B.n394 10.6151
R2107 B.n578 B.n577 10.6151
R2108 B.n579 B.n578 10.6151
R2109 B.n579 B.n392 10.6151
R2110 B.n585 B.n392 10.6151
R2111 B.n586 B.n585 10.6151
R2112 B.n587 B.n586 10.6151
R2113 B.n587 B.n390 10.6151
R2114 B.n593 B.n390 10.6151
R2115 B.n594 B.n593 10.6151
R2116 B.n595 B.n594 10.6151
R2117 B.n595 B.n388 10.6151
R2118 B.n388 B.n387 10.6151
R2119 B.n602 B.n387 10.6151
R2120 B.n603 B.n602 10.6151
R2121 B.n604 B.n379 10.6151
R2122 B.n614 B.n379 10.6151
R2123 B.n615 B.n614 10.6151
R2124 B.n616 B.n615 10.6151
R2125 B.n616 B.n371 10.6151
R2126 B.n626 B.n371 10.6151
R2127 B.n627 B.n626 10.6151
R2128 B.n628 B.n627 10.6151
R2129 B.n628 B.n363 10.6151
R2130 B.n638 B.n363 10.6151
R2131 B.n639 B.n638 10.6151
R2132 B.n640 B.n639 10.6151
R2133 B.n640 B.n355 10.6151
R2134 B.n650 B.n355 10.6151
R2135 B.n651 B.n650 10.6151
R2136 B.n652 B.n651 10.6151
R2137 B.n652 B.n348 10.6151
R2138 B.n663 B.n348 10.6151
R2139 B.n664 B.n663 10.6151
R2140 B.n665 B.n664 10.6151
R2141 B.n665 B.n340 10.6151
R2142 B.n675 B.n340 10.6151
R2143 B.n676 B.n675 10.6151
R2144 B.n677 B.n676 10.6151
R2145 B.n677 B.n332 10.6151
R2146 B.n687 B.n332 10.6151
R2147 B.n688 B.n687 10.6151
R2148 B.n689 B.n688 10.6151
R2149 B.n689 B.n323 10.6151
R2150 B.n699 B.n323 10.6151
R2151 B.n700 B.n699 10.6151
R2152 B.n701 B.n700 10.6151
R2153 B.n701 B.n316 10.6151
R2154 B.n711 B.n316 10.6151
R2155 B.n712 B.n711 10.6151
R2156 B.n713 B.n712 10.6151
R2157 B.n713 B.n307 10.6151
R2158 B.n723 B.n307 10.6151
R2159 B.n724 B.n723 10.6151
R2160 B.n726 B.n724 10.6151
R2161 B.n726 B.n725 10.6151
R2162 B.n725 B.n300 10.6151
R2163 B.n737 B.n300 10.6151
R2164 B.n738 B.n737 10.6151
R2165 B.n739 B.n738 10.6151
R2166 B.n740 B.n739 10.6151
R2167 B.n741 B.n740 10.6151
R2168 B.n744 B.n741 10.6151
R2169 B.n745 B.n744 10.6151
R2170 B.n746 B.n745 10.6151
R2171 B.n747 B.n746 10.6151
R2172 B.n749 B.n747 10.6151
R2173 B.n750 B.n749 10.6151
R2174 B.n751 B.n750 10.6151
R2175 B.n752 B.n751 10.6151
R2176 B.n754 B.n752 10.6151
R2177 B.n755 B.n754 10.6151
R2178 B.n756 B.n755 10.6151
R2179 B.n757 B.n756 10.6151
R2180 B.n759 B.n757 10.6151
R2181 B.n760 B.n759 10.6151
R2182 B.n761 B.n760 10.6151
R2183 B.n762 B.n761 10.6151
R2184 B.n764 B.n762 10.6151
R2185 B.n765 B.n764 10.6151
R2186 B.n766 B.n765 10.6151
R2187 B.n767 B.n766 10.6151
R2188 B.n769 B.n767 10.6151
R2189 B.n770 B.n769 10.6151
R2190 B.n771 B.n770 10.6151
R2191 B.n772 B.n771 10.6151
R2192 B.n774 B.n772 10.6151
R2193 B.n775 B.n774 10.6151
R2194 B.n776 B.n775 10.6151
R2195 B.n777 B.n776 10.6151
R2196 B.n779 B.n777 10.6151
R2197 B.n780 B.n779 10.6151
R2198 B.n781 B.n780 10.6151
R2199 B.n782 B.n781 10.6151
R2200 B.n784 B.n782 10.6151
R2201 B.n785 B.n784 10.6151
R2202 B.n786 B.n785 10.6151
R2203 B.n787 B.n786 10.6151
R2204 B.n789 B.n787 10.6151
R2205 B.n790 B.n789 10.6151
R2206 B.n791 B.n790 10.6151
R2207 B.n792 B.n791 10.6151
R2208 B.n794 B.n792 10.6151
R2209 B.n795 B.n794 10.6151
R2210 B.n884 B.n1 10.6151
R2211 B.n884 B.n883 10.6151
R2212 B.n883 B.n882 10.6151
R2213 B.n882 B.n10 10.6151
R2214 B.n876 B.n10 10.6151
R2215 B.n876 B.n875 10.6151
R2216 B.n875 B.n874 10.6151
R2217 B.n874 B.n18 10.6151
R2218 B.n868 B.n18 10.6151
R2219 B.n868 B.n867 10.6151
R2220 B.n867 B.n866 10.6151
R2221 B.n866 B.n25 10.6151
R2222 B.n860 B.n25 10.6151
R2223 B.n860 B.n859 10.6151
R2224 B.n859 B.n858 10.6151
R2225 B.n858 B.n32 10.6151
R2226 B.n852 B.n32 10.6151
R2227 B.n852 B.n851 10.6151
R2228 B.n851 B.n850 10.6151
R2229 B.n850 B.n39 10.6151
R2230 B.n844 B.n39 10.6151
R2231 B.n844 B.n843 10.6151
R2232 B.n843 B.n842 10.6151
R2233 B.n842 B.n46 10.6151
R2234 B.n836 B.n46 10.6151
R2235 B.n836 B.n835 10.6151
R2236 B.n835 B.n834 10.6151
R2237 B.n834 B.n52 10.6151
R2238 B.n828 B.n52 10.6151
R2239 B.n828 B.n827 10.6151
R2240 B.n827 B.n826 10.6151
R2241 B.n826 B.n60 10.6151
R2242 B.n820 B.n60 10.6151
R2243 B.n820 B.n819 10.6151
R2244 B.n819 B.n818 10.6151
R2245 B.n818 B.n67 10.6151
R2246 B.n812 B.n67 10.6151
R2247 B.n812 B.n811 10.6151
R2248 B.n811 B.n810 10.6151
R2249 B.n810 B.n74 10.6151
R2250 B.n804 B.n74 10.6151
R2251 B.n804 B.n803 10.6151
R2252 B.n803 B.n802 10.6151
R2253 B.n133 B.n81 10.6151
R2254 B.n136 B.n133 10.6151
R2255 B.n137 B.n136 10.6151
R2256 B.n140 B.n137 10.6151
R2257 B.n141 B.n140 10.6151
R2258 B.n144 B.n141 10.6151
R2259 B.n145 B.n144 10.6151
R2260 B.n148 B.n145 10.6151
R2261 B.n149 B.n148 10.6151
R2262 B.n152 B.n149 10.6151
R2263 B.n153 B.n152 10.6151
R2264 B.n156 B.n153 10.6151
R2265 B.n157 B.n156 10.6151
R2266 B.n160 B.n157 10.6151
R2267 B.n161 B.n160 10.6151
R2268 B.n164 B.n161 10.6151
R2269 B.n165 B.n164 10.6151
R2270 B.n168 B.n165 10.6151
R2271 B.n169 B.n168 10.6151
R2272 B.n172 B.n169 10.6151
R2273 B.n173 B.n172 10.6151
R2274 B.n176 B.n173 10.6151
R2275 B.n177 B.n176 10.6151
R2276 B.n180 B.n177 10.6151
R2277 B.n181 B.n180 10.6151
R2278 B.n184 B.n181 10.6151
R2279 B.n185 B.n184 10.6151
R2280 B.n188 B.n185 10.6151
R2281 B.n189 B.n188 10.6151
R2282 B.n192 B.n189 10.6151
R2283 B.n193 B.n192 10.6151
R2284 B.n196 B.n193 10.6151
R2285 B.n197 B.n196 10.6151
R2286 B.n200 B.n197 10.6151
R2287 B.n201 B.n200 10.6151
R2288 B.n204 B.n201 10.6151
R2289 B.n205 B.n204 10.6151
R2290 B.n209 B.n208 10.6151
R2291 B.n212 B.n209 10.6151
R2292 B.n213 B.n212 10.6151
R2293 B.n216 B.n213 10.6151
R2294 B.n217 B.n216 10.6151
R2295 B.n220 B.n217 10.6151
R2296 B.n221 B.n220 10.6151
R2297 B.n224 B.n221 10.6151
R2298 B.n225 B.n224 10.6151
R2299 B.n229 B.n228 10.6151
R2300 B.n232 B.n229 10.6151
R2301 B.n233 B.n232 10.6151
R2302 B.n236 B.n233 10.6151
R2303 B.n237 B.n236 10.6151
R2304 B.n240 B.n237 10.6151
R2305 B.n241 B.n240 10.6151
R2306 B.n244 B.n241 10.6151
R2307 B.n245 B.n244 10.6151
R2308 B.n248 B.n245 10.6151
R2309 B.n249 B.n248 10.6151
R2310 B.n252 B.n249 10.6151
R2311 B.n253 B.n252 10.6151
R2312 B.n256 B.n253 10.6151
R2313 B.n257 B.n256 10.6151
R2314 B.n260 B.n257 10.6151
R2315 B.n261 B.n260 10.6151
R2316 B.n264 B.n261 10.6151
R2317 B.n265 B.n264 10.6151
R2318 B.n268 B.n265 10.6151
R2319 B.n269 B.n268 10.6151
R2320 B.n272 B.n269 10.6151
R2321 B.n273 B.n272 10.6151
R2322 B.n276 B.n273 10.6151
R2323 B.n277 B.n276 10.6151
R2324 B.n280 B.n277 10.6151
R2325 B.n281 B.n280 10.6151
R2326 B.n284 B.n281 10.6151
R2327 B.n285 B.n284 10.6151
R2328 B.n288 B.n285 10.6151
R2329 B.n289 B.n288 10.6151
R2330 B.n292 B.n289 10.6151
R2331 B.n293 B.n292 10.6151
R2332 B.n296 B.n293 10.6151
R2333 B.n298 B.n296 10.6151
R2334 B.n299 B.n298 10.6151
R2335 B.n796 B.n299 10.6151
R2336 B.n506 B.n505 9.36635
R2337 B.n530 B.n529 9.36635
R2338 B.n205 B.n132 9.36635
R2339 B.n228 B.n129 9.36635
R2340 B.n892 B.n0 8.11757
R2341 B.n892 B.n1 8.11757
R2342 B.n703 B.t6 4.09861
R2343 B.n864 B.t3 4.09861
R2344 B.n505 B.n412 1.24928
R2345 B.n529 B.n528 1.24928
R2346 B.n208 B.n132 1.24928
R2347 B.n225 B.n129 1.24928
R2348 VP.n16 VP.n15 161.3
R2349 VP.n17 VP.n12 161.3
R2350 VP.n19 VP.n18 161.3
R2351 VP.n20 VP.n11 161.3
R2352 VP.n22 VP.n21 161.3
R2353 VP.n24 VP.n10 161.3
R2354 VP.n26 VP.n25 161.3
R2355 VP.n27 VP.n9 161.3
R2356 VP.n29 VP.n28 161.3
R2357 VP.n30 VP.n8 161.3
R2358 VP.n58 VP.n0 161.3
R2359 VP.n57 VP.n56 161.3
R2360 VP.n55 VP.n1 161.3
R2361 VP.n54 VP.n53 161.3
R2362 VP.n52 VP.n2 161.3
R2363 VP.n50 VP.n49 161.3
R2364 VP.n48 VP.n3 161.3
R2365 VP.n47 VP.n46 161.3
R2366 VP.n45 VP.n4 161.3
R2367 VP.n44 VP.n43 161.3
R2368 VP.n42 VP.n41 161.3
R2369 VP.n40 VP.n6 161.3
R2370 VP.n39 VP.n38 161.3
R2371 VP.n37 VP.n7 161.3
R2372 VP.n36 VP.n35 161.3
R2373 VP.n14 VP.t6 152.594
R2374 VP.n34 VP.t5 120.835
R2375 VP.n5 VP.t4 120.835
R2376 VP.n51 VP.t3 120.835
R2377 VP.n59 VP.t0 120.835
R2378 VP.n31 VP.t1 120.835
R2379 VP.n23 VP.t2 120.835
R2380 VP.n13 VP.t7 120.835
R2381 VP.n34 VP.n33 99.257
R2382 VP.n60 VP.n59 99.257
R2383 VP.n32 VP.n31 99.257
R2384 VP.n14 VP.n13 59.5219
R2385 VP.n33 VP.n32 47.886
R2386 VP.n40 VP.n39 41.4647
R2387 VP.n53 VP.n1 41.4647
R2388 VP.n25 VP.n9 41.4647
R2389 VP.n46 VP.n45 40.4934
R2390 VP.n46 VP.n3 40.4934
R2391 VP.n18 VP.n11 40.4934
R2392 VP.n18 VP.n17 40.4934
R2393 VP.n39 VP.n7 39.5221
R2394 VP.n57 VP.n1 39.5221
R2395 VP.n29 VP.n9 39.5221
R2396 VP.n35 VP.n7 24.4675
R2397 VP.n41 VP.n40 24.4675
R2398 VP.n45 VP.n44 24.4675
R2399 VP.n50 VP.n3 24.4675
R2400 VP.n53 VP.n52 24.4675
R2401 VP.n58 VP.n57 24.4675
R2402 VP.n30 VP.n29 24.4675
R2403 VP.n22 VP.n11 24.4675
R2404 VP.n25 VP.n24 24.4675
R2405 VP.n17 VP.n16 24.4675
R2406 VP.n41 VP.n5 12.4787
R2407 VP.n52 VP.n51 12.4787
R2408 VP.n24 VP.n23 12.4787
R2409 VP.n44 VP.n5 11.9893
R2410 VP.n51 VP.n50 11.9893
R2411 VP.n23 VP.n22 11.9893
R2412 VP.n16 VP.n13 11.9893
R2413 VP.n35 VP.n34 11.5
R2414 VP.n59 VP.n58 11.5
R2415 VP.n31 VP.n30 11.5
R2416 VP.n15 VP.n14 9.80091
R2417 VP.n32 VP.n8 0.278367
R2418 VP.n36 VP.n33 0.278367
R2419 VP.n60 VP.n0 0.278367
R2420 VP.n15 VP.n12 0.189894
R2421 VP.n19 VP.n12 0.189894
R2422 VP.n20 VP.n19 0.189894
R2423 VP.n21 VP.n20 0.189894
R2424 VP.n21 VP.n10 0.189894
R2425 VP.n26 VP.n10 0.189894
R2426 VP.n27 VP.n26 0.189894
R2427 VP.n28 VP.n27 0.189894
R2428 VP.n28 VP.n8 0.189894
R2429 VP.n37 VP.n36 0.189894
R2430 VP.n38 VP.n37 0.189894
R2431 VP.n38 VP.n6 0.189894
R2432 VP.n42 VP.n6 0.189894
R2433 VP.n43 VP.n42 0.189894
R2434 VP.n43 VP.n4 0.189894
R2435 VP.n47 VP.n4 0.189894
R2436 VP.n48 VP.n47 0.189894
R2437 VP.n49 VP.n48 0.189894
R2438 VP.n49 VP.n2 0.189894
R2439 VP.n54 VP.n2 0.189894
R2440 VP.n55 VP.n54 0.189894
R2441 VP.n56 VP.n55 0.189894
R2442 VP.n56 VP.n0 0.189894
R2443 VP VP.n60 0.153454
R2444 VDD1 VDD1.n0 66.3808
R2445 VDD1.n3 VDD1.n2 66.2671
R2446 VDD1.n3 VDD1.n1 66.2671
R2447 VDD1.n5 VDD1.n4 65.2492
R2448 VDD1.n5 VDD1.n3 43.294
R2449 VDD1.n4 VDD1.t5 1.82875
R2450 VDD1.n4 VDD1.t6 1.82875
R2451 VDD1.n0 VDD1.t1 1.82875
R2452 VDD1.n0 VDD1.t0 1.82875
R2453 VDD1.n2 VDD1.t4 1.82875
R2454 VDD1.n2 VDD1.t7 1.82875
R2455 VDD1.n1 VDD1.t2 1.82875
R2456 VDD1.n1 VDD1.t3 1.82875
R2457 VDD1 VDD1.n5 1.01559
C0 VDD1 VP 7.91293f
C1 VDD1 VN 0.150457f
C2 VDD2 VP 0.472375f
C3 VDD2 VN 7.59219f
C4 VDD1 VTAIL 7.62886f
C5 VDD2 VTAIL 7.68033f
C6 VP VN 6.912529f
C7 VDD1 VDD2 1.54508f
C8 VP VTAIL 7.90482f
C9 VN VTAIL 7.89071f
C10 VDD2 B 4.825999f
C11 VDD1 B 5.213513f
C12 VTAIL B 9.47539f
C13 VN B 13.750831f
C14 VP B 12.301099f
C15 VDD1.t1 B 0.211303f
C16 VDD1.t0 B 0.211303f
C17 VDD1.n0 B 1.8812f
C18 VDD1.t2 B 0.211303f
C19 VDD1.t3 B 0.211303f
C20 VDD1.n1 B 1.88027f
C21 VDD1.t4 B 0.211303f
C22 VDD1.t7 B 0.211303f
C23 VDD1.n2 B 1.88027f
C24 VDD1.n3 B 2.9599f
C25 VDD1.t5 B 0.211303f
C26 VDD1.t6 B 0.211303f
C27 VDD1.n4 B 1.87317f
C28 VDD1.n5 B 2.70104f
C29 VP.n0 B 0.033697f
C30 VP.t0 B 1.62402f
C31 VP.n1 B 0.020695f
C32 VP.n2 B 0.025559f
C33 VP.t3 B 1.62402f
C34 VP.n3 B 0.050799f
C35 VP.n4 B 0.025559f
C36 VP.t4 B 1.62402f
C37 VP.n5 B 0.582047f
C38 VP.n6 B 0.025559f
C39 VP.n7 B 0.051038f
C40 VP.n8 B 0.033697f
C41 VP.t1 B 1.62402f
C42 VP.n9 B 0.020695f
C43 VP.n10 B 0.025559f
C44 VP.t2 B 1.62402f
C45 VP.n11 B 0.050799f
C46 VP.n12 B 0.025559f
C47 VP.t7 B 1.62402f
C48 VP.n13 B 0.647049f
C49 VP.t6 B 1.77294f
C50 VP.n14 B 0.642243f
C51 VP.n15 B 0.216279f
C52 VP.n16 B 0.03564f
C53 VP.n17 B 0.050799f
C54 VP.n18 B 0.020662f
C55 VP.n19 B 0.025559f
C56 VP.n20 B 0.025559f
C57 VP.n21 B 0.025559f
C58 VP.n22 B 0.03564f
C59 VP.n23 B 0.582047f
C60 VP.n24 B 0.036111f
C61 VP.n25 B 0.050526f
C62 VP.n26 B 0.025559f
C63 VP.n27 B 0.025559f
C64 VP.n28 B 0.025559f
C65 VP.n29 B 0.051038f
C66 VP.n30 B 0.03517f
C67 VP.n31 B 0.654422f
C68 VP.n32 B 1.32812f
C69 VP.n33 B 1.3473f
C70 VP.t5 B 1.62402f
C71 VP.n34 B 0.654422f
C72 VP.n35 B 0.03517f
C73 VP.n36 B 0.033697f
C74 VP.n37 B 0.025559f
C75 VP.n38 B 0.025559f
C76 VP.n39 B 0.020695f
C77 VP.n40 B 0.050526f
C78 VP.n41 B 0.036111f
C79 VP.n42 B 0.025559f
C80 VP.n43 B 0.025559f
C81 VP.n44 B 0.03564f
C82 VP.n45 B 0.050799f
C83 VP.n46 B 0.020662f
C84 VP.n47 B 0.025559f
C85 VP.n48 B 0.025559f
C86 VP.n49 B 0.025559f
C87 VP.n50 B 0.03564f
C88 VP.n51 B 0.582047f
C89 VP.n52 B 0.036111f
C90 VP.n53 B 0.050526f
C91 VP.n54 B 0.025559f
C92 VP.n55 B 0.025559f
C93 VP.n56 B 0.025559f
C94 VP.n57 B 0.051038f
C95 VP.n58 B 0.03517f
C96 VP.n59 B 0.654422f
C97 VP.n60 B 0.037287f
C98 VDD2.t2 B 0.209811f
C99 VDD2.t0 B 0.209811f
C100 VDD2.n0 B 1.867f
C101 VDD2.t6 B 0.209811f
C102 VDD2.t4 B 0.209811f
C103 VDD2.n1 B 1.867f
C104 VDD2.n2 B 2.88764f
C105 VDD2.t5 B 0.209811f
C106 VDD2.t7 B 0.209811f
C107 VDD2.n3 B 1.85995f
C108 VDD2.n4 B 2.65197f
C109 VDD2.t1 B 0.209811f
C110 VDD2.t3 B 0.209811f
C111 VDD2.n5 B 1.86697f
C112 VTAIL.t9 B 0.169998f
C113 VTAIL.t12 B 0.169998f
C114 VTAIL.n0 B 1.45299f
C115 VTAIL.n1 B 0.329235f
C116 VTAIL.n2 B 0.028858f
C117 VTAIL.n3 B 0.019864f
C118 VTAIL.n4 B 0.010674f
C119 VTAIL.n5 B 0.025229f
C120 VTAIL.n6 B 0.011302f
C121 VTAIL.n7 B 0.019864f
C122 VTAIL.n8 B 0.010674f
C123 VTAIL.n9 B 0.025229f
C124 VTAIL.n10 B 0.011302f
C125 VTAIL.n11 B 0.019864f
C126 VTAIL.n12 B 0.010674f
C127 VTAIL.n13 B 0.025229f
C128 VTAIL.n14 B 0.011302f
C129 VTAIL.n15 B 0.019864f
C130 VTAIL.n16 B 0.010674f
C131 VTAIL.n17 B 0.025229f
C132 VTAIL.n18 B 0.011302f
C133 VTAIL.n19 B 0.134295f
C134 VTAIL.t15 B 0.042486f
C135 VTAIL.n20 B 0.018922f
C136 VTAIL.n21 B 0.017835f
C137 VTAIL.n22 B 0.010674f
C138 VTAIL.n23 B 0.898721f
C139 VTAIL.n24 B 0.019864f
C140 VTAIL.n25 B 0.010674f
C141 VTAIL.n26 B 0.011302f
C142 VTAIL.n27 B 0.025229f
C143 VTAIL.n28 B 0.025229f
C144 VTAIL.n29 B 0.011302f
C145 VTAIL.n30 B 0.010674f
C146 VTAIL.n31 B 0.019864f
C147 VTAIL.n32 B 0.019864f
C148 VTAIL.n33 B 0.010674f
C149 VTAIL.n34 B 0.011302f
C150 VTAIL.n35 B 0.025229f
C151 VTAIL.n36 B 0.025229f
C152 VTAIL.n37 B 0.025229f
C153 VTAIL.n38 B 0.011302f
C154 VTAIL.n39 B 0.010674f
C155 VTAIL.n40 B 0.019864f
C156 VTAIL.n41 B 0.019864f
C157 VTAIL.n42 B 0.010674f
C158 VTAIL.n43 B 0.010988f
C159 VTAIL.n44 B 0.010988f
C160 VTAIL.n45 B 0.025229f
C161 VTAIL.n46 B 0.025229f
C162 VTAIL.n47 B 0.011302f
C163 VTAIL.n48 B 0.010674f
C164 VTAIL.n49 B 0.019864f
C165 VTAIL.n50 B 0.019864f
C166 VTAIL.n51 B 0.010674f
C167 VTAIL.n52 B 0.011302f
C168 VTAIL.n53 B 0.025229f
C169 VTAIL.n54 B 0.056276f
C170 VTAIL.n55 B 0.011302f
C171 VTAIL.n56 B 0.010674f
C172 VTAIL.n57 B 0.049985f
C173 VTAIL.n58 B 0.03178f
C174 VTAIL.n59 B 0.18673f
C175 VTAIL.n60 B 0.028858f
C176 VTAIL.n61 B 0.019864f
C177 VTAIL.n62 B 0.010674f
C178 VTAIL.n63 B 0.025229f
C179 VTAIL.n64 B 0.011302f
C180 VTAIL.n65 B 0.019864f
C181 VTAIL.n66 B 0.010674f
C182 VTAIL.n67 B 0.025229f
C183 VTAIL.n68 B 0.011302f
C184 VTAIL.n69 B 0.019864f
C185 VTAIL.n70 B 0.010674f
C186 VTAIL.n71 B 0.025229f
C187 VTAIL.n72 B 0.011302f
C188 VTAIL.n73 B 0.019864f
C189 VTAIL.n74 B 0.010674f
C190 VTAIL.n75 B 0.025229f
C191 VTAIL.n76 B 0.011302f
C192 VTAIL.n77 B 0.134295f
C193 VTAIL.t2 B 0.042486f
C194 VTAIL.n78 B 0.018922f
C195 VTAIL.n79 B 0.017835f
C196 VTAIL.n80 B 0.010674f
C197 VTAIL.n81 B 0.898721f
C198 VTAIL.n82 B 0.019864f
C199 VTAIL.n83 B 0.010674f
C200 VTAIL.n84 B 0.011302f
C201 VTAIL.n85 B 0.025229f
C202 VTAIL.n86 B 0.025229f
C203 VTAIL.n87 B 0.011302f
C204 VTAIL.n88 B 0.010674f
C205 VTAIL.n89 B 0.019864f
C206 VTAIL.n90 B 0.019864f
C207 VTAIL.n91 B 0.010674f
C208 VTAIL.n92 B 0.011302f
C209 VTAIL.n93 B 0.025229f
C210 VTAIL.n94 B 0.025229f
C211 VTAIL.n95 B 0.025229f
C212 VTAIL.n96 B 0.011302f
C213 VTAIL.n97 B 0.010674f
C214 VTAIL.n98 B 0.019864f
C215 VTAIL.n99 B 0.019864f
C216 VTAIL.n100 B 0.010674f
C217 VTAIL.n101 B 0.010988f
C218 VTAIL.n102 B 0.010988f
C219 VTAIL.n103 B 0.025229f
C220 VTAIL.n104 B 0.025229f
C221 VTAIL.n105 B 0.011302f
C222 VTAIL.n106 B 0.010674f
C223 VTAIL.n107 B 0.019864f
C224 VTAIL.n108 B 0.019864f
C225 VTAIL.n109 B 0.010674f
C226 VTAIL.n110 B 0.011302f
C227 VTAIL.n111 B 0.025229f
C228 VTAIL.n112 B 0.056276f
C229 VTAIL.n113 B 0.011302f
C230 VTAIL.n114 B 0.010674f
C231 VTAIL.n115 B 0.049985f
C232 VTAIL.n116 B 0.03178f
C233 VTAIL.n117 B 0.18673f
C234 VTAIL.t5 B 0.169998f
C235 VTAIL.t6 B 0.169998f
C236 VTAIL.n118 B 1.45299f
C237 VTAIL.n119 B 0.462902f
C238 VTAIL.n120 B 0.028858f
C239 VTAIL.n121 B 0.019864f
C240 VTAIL.n122 B 0.010674f
C241 VTAIL.n123 B 0.025229f
C242 VTAIL.n124 B 0.011302f
C243 VTAIL.n125 B 0.019864f
C244 VTAIL.n126 B 0.010674f
C245 VTAIL.n127 B 0.025229f
C246 VTAIL.n128 B 0.011302f
C247 VTAIL.n129 B 0.019864f
C248 VTAIL.n130 B 0.010674f
C249 VTAIL.n131 B 0.025229f
C250 VTAIL.n132 B 0.011302f
C251 VTAIL.n133 B 0.019864f
C252 VTAIL.n134 B 0.010674f
C253 VTAIL.n135 B 0.025229f
C254 VTAIL.n136 B 0.011302f
C255 VTAIL.n137 B 0.134295f
C256 VTAIL.t0 B 0.042486f
C257 VTAIL.n138 B 0.018922f
C258 VTAIL.n139 B 0.017835f
C259 VTAIL.n140 B 0.010674f
C260 VTAIL.n141 B 0.898721f
C261 VTAIL.n142 B 0.019864f
C262 VTAIL.n143 B 0.010674f
C263 VTAIL.n144 B 0.011302f
C264 VTAIL.n145 B 0.025229f
C265 VTAIL.n146 B 0.025229f
C266 VTAIL.n147 B 0.011302f
C267 VTAIL.n148 B 0.010674f
C268 VTAIL.n149 B 0.019864f
C269 VTAIL.n150 B 0.019864f
C270 VTAIL.n151 B 0.010674f
C271 VTAIL.n152 B 0.011302f
C272 VTAIL.n153 B 0.025229f
C273 VTAIL.n154 B 0.025229f
C274 VTAIL.n155 B 0.025229f
C275 VTAIL.n156 B 0.011302f
C276 VTAIL.n157 B 0.010674f
C277 VTAIL.n158 B 0.019864f
C278 VTAIL.n159 B 0.019864f
C279 VTAIL.n160 B 0.010674f
C280 VTAIL.n161 B 0.010988f
C281 VTAIL.n162 B 0.010988f
C282 VTAIL.n163 B 0.025229f
C283 VTAIL.n164 B 0.025229f
C284 VTAIL.n165 B 0.011302f
C285 VTAIL.n166 B 0.010674f
C286 VTAIL.n167 B 0.019864f
C287 VTAIL.n168 B 0.019864f
C288 VTAIL.n169 B 0.010674f
C289 VTAIL.n170 B 0.011302f
C290 VTAIL.n171 B 0.025229f
C291 VTAIL.n172 B 0.056276f
C292 VTAIL.n173 B 0.011302f
C293 VTAIL.n174 B 0.010674f
C294 VTAIL.n175 B 0.049985f
C295 VTAIL.n176 B 0.03178f
C296 VTAIL.n177 B 1.16145f
C297 VTAIL.n178 B 0.028858f
C298 VTAIL.n179 B 0.019864f
C299 VTAIL.n180 B 0.010674f
C300 VTAIL.n181 B 0.025229f
C301 VTAIL.n182 B 0.011302f
C302 VTAIL.n183 B 0.019864f
C303 VTAIL.n184 B 0.010674f
C304 VTAIL.n185 B 0.025229f
C305 VTAIL.n186 B 0.011302f
C306 VTAIL.n187 B 0.019864f
C307 VTAIL.n188 B 0.010674f
C308 VTAIL.n189 B 0.025229f
C309 VTAIL.n190 B 0.025229f
C310 VTAIL.n191 B 0.011302f
C311 VTAIL.n192 B 0.019864f
C312 VTAIL.n193 B 0.010674f
C313 VTAIL.n194 B 0.025229f
C314 VTAIL.n195 B 0.011302f
C315 VTAIL.n196 B 0.134295f
C316 VTAIL.t8 B 0.042486f
C317 VTAIL.n197 B 0.018922f
C318 VTAIL.n198 B 0.017835f
C319 VTAIL.n199 B 0.010674f
C320 VTAIL.n200 B 0.898721f
C321 VTAIL.n201 B 0.019864f
C322 VTAIL.n202 B 0.010674f
C323 VTAIL.n203 B 0.011302f
C324 VTAIL.n204 B 0.025229f
C325 VTAIL.n205 B 0.025229f
C326 VTAIL.n206 B 0.011302f
C327 VTAIL.n207 B 0.010674f
C328 VTAIL.n208 B 0.019864f
C329 VTAIL.n209 B 0.019864f
C330 VTAIL.n210 B 0.010674f
C331 VTAIL.n211 B 0.011302f
C332 VTAIL.n212 B 0.025229f
C333 VTAIL.n213 B 0.025229f
C334 VTAIL.n214 B 0.011302f
C335 VTAIL.n215 B 0.010674f
C336 VTAIL.n216 B 0.019864f
C337 VTAIL.n217 B 0.019864f
C338 VTAIL.n218 B 0.010674f
C339 VTAIL.n219 B 0.010988f
C340 VTAIL.n220 B 0.010988f
C341 VTAIL.n221 B 0.025229f
C342 VTAIL.n222 B 0.025229f
C343 VTAIL.n223 B 0.011302f
C344 VTAIL.n224 B 0.010674f
C345 VTAIL.n225 B 0.019864f
C346 VTAIL.n226 B 0.019864f
C347 VTAIL.n227 B 0.010674f
C348 VTAIL.n228 B 0.011302f
C349 VTAIL.n229 B 0.025229f
C350 VTAIL.n230 B 0.056276f
C351 VTAIL.n231 B 0.011302f
C352 VTAIL.n232 B 0.010674f
C353 VTAIL.n233 B 0.049985f
C354 VTAIL.n234 B 0.03178f
C355 VTAIL.n235 B 1.16145f
C356 VTAIL.t14 B 0.169998f
C357 VTAIL.t13 B 0.169998f
C358 VTAIL.n236 B 1.45299f
C359 VTAIL.n237 B 0.462894f
C360 VTAIL.n238 B 0.028858f
C361 VTAIL.n239 B 0.019864f
C362 VTAIL.n240 B 0.010674f
C363 VTAIL.n241 B 0.025229f
C364 VTAIL.n242 B 0.011302f
C365 VTAIL.n243 B 0.019864f
C366 VTAIL.n244 B 0.010674f
C367 VTAIL.n245 B 0.025229f
C368 VTAIL.n246 B 0.011302f
C369 VTAIL.n247 B 0.019864f
C370 VTAIL.n248 B 0.010674f
C371 VTAIL.n249 B 0.025229f
C372 VTAIL.n250 B 0.025229f
C373 VTAIL.n251 B 0.011302f
C374 VTAIL.n252 B 0.019864f
C375 VTAIL.n253 B 0.010674f
C376 VTAIL.n254 B 0.025229f
C377 VTAIL.n255 B 0.011302f
C378 VTAIL.n256 B 0.134295f
C379 VTAIL.t10 B 0.042486f
C380 VTAIL.n257 B 0.018922f
C381 VTAIL.n258 B 0.017835f
C382 VTAIL.n259 B 0.010674f
C383 VTAIL.n260 B 0.898721f
C384 VTAIL.n261 B 0.019864f
C385 VTAIL.n262 B 0.010674f
C386 VTAIL.n263 B 0.011302f
C387 VTAIL.n264 B 0.025229f
C388 VTAIL.n265 B 0.025229f
C389 VTAIL.n266 B 0.011302f
C390 VTAIL.n267 B 0.010674f
C391 VTAIL.n268 B 0.019864f
C392 VTAIL.n269 B 0.019864f
C393 VTAIL.n270 B 0.010674f
C394 VTAIL.n271 B 0.011302f
C395 VTAIL.n272 B 0.025229f
C396 VTAIL.n273 B 0.025229f
C397 VTAIL.n274 B 0.011302f
C398 VTAIL.n275 B 0.010674f
C399 VTAIL.n276 B 0.019864f
C400 VTAIL.n277 B 0.019864f
C401 VTAIL.n278 B 0.010674f
C402 VTAIL.n279 B 0.010988f
C403 VTAIL.n280 B 0.010988f
C404 VTAIL.n281 B 0.025229f
C405 VTAIL.n282 B 0.025229f
C406 VTAIL.n283 B 0.011302f
C407 VTAIL.n284 B 0.010674f
C408 VTAIL.n285 B 0.019864f
C409 VTAIL.n286 B 0.019864f
C410 VTAIL.n287 B 0.010674f
C411 VTAIL.n288 B 0.011302f
C412 VTAIL.n289 B 0.025229f
C413 VTAIL.n290 B 0.056276f
C414 VTAIL.n291 B 0.011302f
C415 VTAIL.n292 B 0.010674f
C416 VTAIL.n293 B 0.049985f
C417 VTAIL.n294 B 0.03178f
C418 VTAIL.n295 B 0.18673f
C419 VTAIL.n296 B 0.028858f
C420 VTAIL.n297 B 0.019864f
C421 VTAIL.n298 B 0.010674f
C422 VTAIL.n299 B 0.025229f
C423 VTAIL.n300 B 0.011302f
C424 VTAIL.n301 B 0.019864f
C425 VTAIL.n302 B 0.010674f
C426 VTAIL.n303 B 0.025229f
C427 VTAIL.n304 B 0.011302f
C428 VTAIL.n305 B 0.019864f
C429 VTAIL.n306 B 0.010674f
C430 VTAIL.n307 B 0.025229f
C431 VTAIL.n308 B 0.025229f
C432 VTAIL.n309 B 0.011302f
C433 VTAIL.n310 B 0.019864f
C434 VTAIL.n311 B 0.010674f
C435 VTAIL.n312 B 0.025229f
C436 VTAIL.n313 B 0.011302f
C437 VTAIL.n314 B 0.134295f
C438 VTAIL.t4 B 0.042486f
C439 VTAIL.n315 B 0.018922f
C440 VTAIL.n316 B 0.017835f
C441 VTAIL.n317 B 0.010674f
C442 VTAIL.n318 B 0.898721f
C443 VTAIL.n319 B 0.019864f
C444 VTAIL.n320 B 0.010674f
C445 VTAIL.n321 B 0.011302f
C446 VTAIL.n322 B 0.025229f
C447 VTAIL.n323 B 0.025229f
C448 VTAIL.n324 B 0.011302f
C449 VTAIL.n325 B 0.010674f
C450 VTAIL.n326 B 0.019864f
C451 VTAIL.n327 B 0.019864f
C452 VTAIL.n328 B 0.010674f
C453 VTAIL.n329 B 0.011302f
C454 VTAIL.n330 B 0.025229f
C455 VTAIL.n331 B 0.025229f
C456 VTAIL.n332 B 0.011302f
C457 VTAIL.n333 B 0.010674f
C458 VTAIL.n334 B 0.019864f
C459 VTAIL.n335 B 0.019864f
C460 VTAIL.n336 B 0.010674f
C461 VTAIL.n337 B 0.010988f
C462 VTAIL.n338 B 0.010988f
C463 VTAIL.n339 B 0.025229f
C464 VTAIL.n340 B 0.025229f
C465 VTAIL.n341 B 0.011302f
C466 VTAIL.n342 B 0.010674f
C467 VTAIL.n343 B 0.019864f
C468 VTAIL.n344 B 0.019864f
C469 VTAIL.n345 B 0.010674f
C470 VTAIL.n346 B 0.011302f
C471 VTAIL.n347 B 0.025229f
C472 VTAIL.n348 B 0.056276f
C473 VTAIL.n349 B 0.011302f
C474 VTAIL.n350 B 0.010674f
C475 VTAIL.n351 B 0.049985f
C476 VTAIL.n352 B 0.03178f
C477 VTAIL.n353 B 0.18673f
C478 VTAIL.t3 B 0.169998f
C479 VTAIL.t7 B 0.169998f
C480 VTAIL.n354 B 1.45299f
C481 VTAIL.n355 B 0.462894f
C482 VTAIL.n356 B 0.028858f
C483 VTAIL.n357 B 0.019864f
C484 VTAIL.n358 B 0.010674f
C485 VTAIL.n359 B 0.025229f
C486 VTAIL.n360 B 0.011302f
C487 VTAIL.n361 B 0.019864f
C488 VTAIL.n362 B 0.010674f
C489 VTAIL.n363 B 0.025229f
C490 VTAIL.n364 B 0.011302f
C491 VTAIL.n365 B 0.019864f
C492 VTAIL.n366 B 0.010674f
C493 VTAIL.n367 B 0.025229f
C494 VTAIL.n368 B 0.025229f
C495 VTAIL.n369 B 0.011302f
C496 VTAIL.n370 B 0.019864f
C497 VTAIL.n371 B 0.010674f
C498 VTAIL.n372 B 0.025229f
C499 VTAIL.n373 B 0.011302f
C500 VTAIL.n374 B 0.134295f
C501 VTAIL.t1 B 0.042486f
C502 VTAIL.n375 B 0.018922f
C503 VTAIL.n376 B 0.017835f
C504 VTAIL.n377 B 0.010674f
C505 VTAIL.n378 B 0.898721f
C506 VTAIL.n379 B 0.019864f
C507 VTAIL.n380 B 0.010674f
C508 VTAIL.n381 B 0.011302f
C509 VTAIL.n382 B 0.025229f
C510 VTAIL.n383 B 0.025229f
C511 VTAIL.n384 B 0.011302f
C512 VTAIL.n385 B 0.010674f
C513 VTAIL.n386 B 0.019864f
C514 VTAIL.n387 B 0.019864f
C515 VTAIL.n388 B 0.010674f
C516 VTAIL.n389 B 0.011302f
C517 VTAIL.n390 B 0.025229f
C518 VTAIL.n391 B 0.025229f
C519 VTAIL.n392 B 0.011302f
C520 VTAIL.n393 B 0.010674f
C521 VTAIL.n394 B 0.019864f
C522 VTAIL.n395 B 0.019864f
C523 VTAIL.n396 B 0.010674f
C524 VTAIL.n397 B 0.010988f
C525 VTAIL.n398 B 0.010988f
C526 VTAIL.n399 B 0.025229f
C527 VTAIL.n400 B 0.025229f
C528 VTAIL.n401 B 0.011302f
C529 VTAIL.n402 B 0.010674f
C530 VTAIL.n403 B 0.019864f
C531 VTAIL.n404 B 0.019864f
C532 VTAIL.n405 B 0.010674f
C533 VTAIL.n406 B 0.011302f
C534 VTAIL.n407 B 0.025229f
C535 VTAIL.n408 B 0.056276f
C536 VTAIL.n409 B 0.011302f
C537 VTAIL.n410 B 0.010674f
C538 VTAIL.n411 B 0.049985f
C539 VTAIL.n412 B 0.03178f
C540 VTAIL.n413 B 1.16145f
C541 VTAIL.n414 B 0.028858f
C542 VTAIL.n415 B 0.019864f
C543 VTAIL.n416 B 0.010674f
C544 VTAIL.n417 B 0.025229f
C545 VTAIL.n418 B 0.011302f
C546 VTAIL.n419 B 0.019864f
C547 VTAIL.n420 B 0.010674f
C548 VTAIL.n421 B 0.025229f
C549 VTAIL.n422 B 0.011302f
C550 VTAIL.n423 B 0.019864f
C551 VTAIL.n424 B 0.010674f
C552 VTAIL.n425 B 0.025229f
C553 VTAIL.n426 B 0.011302f
C554 VTAIL.n427 B 0.019864f
C555 VTAIL.n428 B 0.010674f
C556 VTAIL.n429 B 0.025229f
C557 VTAIL.n430 B 0.011302f
C558 VTAIL.n431 B 0.134295f
C559 VTAIL.t11 B 0.042486f
C560 VTAIL.n432 B 0.018922f
C561 VTAIL.n433 B 0.017835f
C562 VTAIL.n434 B 0.010674f
C563 VTAIL.n435 B 0.898721f
C564 VTAIL.n436 B 0.019864f
C565 VTAIL.n437 B 0.010674f
C566 VTAIL.n438 B 0.011302f
C567 VTAIL.n439 B 0.025229f
C568 VTAIL.n440 B 0.025229f
C569 VTAIL.n441 B 0.011302f
C570 VTAIL.n442 B 0.010674f
C571 VTAIL.n443 B 0.019864f
C572 VTAIL.n444 B 0.019864f
C573 VTAIL.n445 B 0.010674f
C574 VTAIL.n446 B 0.011302f
C575 VTAIL.n447 B 0.025229f
C576 VTAIL.n448 B 0.025229f
C577 VTAIL.n449 B 0.025229f
C578 VTAIL.n450 B 0.011302f
C579 VTAIL.n451 B 0.010674f
C580 VTAIL.n452 B 0.019864f
C581 VTAIL.n453 B 0.019864f
C582 VTAIL.n454 B 0.010674f
C583 VTAIL.n455 B 0.010988f
C584 VTAIL.n456 B 0.010988f
C585 VTAIL.n457 B 0.025229f
C586 VTAIL.n458 B 0.025229f
C587 VTAIL.n459 B 0.011302f
C588 VTAIL.n460 B 0.010674f
C589 VTAIL.n461 B 0.019864f
C590 VTAIL.n462 B 0.019864f
C591 VTAIL.n463 B 0.010674f
C592 VTAIL.n464 B 0.011302f
C593 VTAIL.n465 B 0.025229f
C594 VTAIL.n466 B 0.056276f
C595 VTAIL.n467 B 0.011302f
C596 VTAIL.n468 B 0.010674f
C597 VTAIL.n469 B 0.049985f
C598 VTAIL.n470 B 0.03178f
C599 VTAIL.n471 B 1.15772f
C600 VN.n0 B 0.033199f
C601 VN.t3 B 1.60003f
C602 VN.n1 B 0.020389f
C603 VN.n2 B 0.025181f
C604 VN.t1 B 1.60003f
C605 VN.n3 B 0.050048f
C606 VN.n4 B 0.025181f
C607 VN.t7 B 1.60003f
C608 VN.n5 B 0.637488f
C609 VN.t5 B 1.74674f
C610 VN.n6 B 0.632754f
C611 VN.n7 B 0.213084f
C612 VN.n8 B 0.035114f
C613 VN.n9 B 0.050048f
C614 VN.n10 B 0.020357f
C615 VN.n11 B 0.025181f
C616 VN.n12 B 0.025181f
C617 VN.n13 B 0.025181f
C618 VN.n14 B 0.035114f
C619 VN.n15 B 0.573447f
C620 VN.n16 B 0.035577f
C621 VN.n17 B 0.049779f
C622 VN.n18 B 0.025181f
C623 VN.n19 B 0.025181f
C624 VN.n20 B 0.025181f
C625 VN.n21 B 0.050284f
C626 VN.n22 B 0.03465f
C627 VN.n23 B 0.644753f
C628 VN.n24 B 0.036736f
C629 VN.n25 B 0.033199f
C630 VN.t2 B 1.60003f
C631 VN.n26 B 0.020389f
C632 VN.n27 B 0.025181f
C633 VN.t0 B 1.60003f
C634 VN.n28 B 0.050048f
C635 VN.n29 B 0.025181f
C636 VN.t6 B 1.60003f
C637 VN.n30 B 0.637488f
C638 VN.t4 B 1.74674f
C639 VN.n31 B 0.632754f
C640 VN.n32 B 0.213084f
C641 VN.n33 B 0.035114f
C642 VN.n34 B 0.050048f
C643 VN.n35 B 0.020357f
C644 VN.n36 B 0.025181f
C645 VN.n37 B 0.025181f
C646 VN.n38 B 0.025181f
C647 VN.n39 B 0.035114f
C648 VN.n40 B 0.573447f
C649 VN.n41 B 0.035577f
C650 VN.n42 B 0.049779f
C651 VN.n43 B 0.025181f
C652 VN.n44 B 0.025181f
C653 VN.n45 B 0.025181f
C654 VN.n46 B 0.050284f
C655 VN.n47 B 0.03465f
C656 VN.n48 B 0.644753f
C657 VN.n49 B 1.32212f
.ends

