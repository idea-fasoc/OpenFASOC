* NGSPICE file created from diff_pair_sample_0669.ext - technology: sky130A

.subckt diff_pair_sample_0669 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t3 VP.t0 VTAIL.t5 w_n1594_n3298# sky130_fd_pr__pfet_01v8 ad=1.92225 pd=11.98 as=4.5435 ps=24.08 w=11.65 l=0.71
X1 VTAIL.t1 VN.t0 VDD2.t3 w_n1594_n3298# sky130_fd_pr__pfet_01v8 ad=4.5435 pd=24.08 as=1.92225 ps=11.98 w=11.65 l=0.71
X2 B.t11 B.t9 B.t10 w_n1594_n3298# sky130_fd_pr__pfet_01v8 ad=4.5435 pd=24.08 as=0 ps=0 w=11.65 l=0.71
X3 VTAIL.t4 VP.t1 VDD1.t2 w_n1594_n3298# sky130_fd_pr__pfet_01v8 ad=4.5435 pd=24.08 as=1.92225 ps=11.98 w=11.65 l=0.71
X4 B.t8 B.t6 B.t7 w_n1594_n3298# sky130_fd_pr__pfet_01v8 ad=4.5435 pd=24.08 as=0 ps=0 w=11.65 l=0.71
X5 VDD2.t2 VN.t1 VTAIL.t0 w_n1594_n3298# sky130_fd_pr__pfet_01v8 ad=1.92225 pd=11.98 as=4.5435 ps=24.08 w=11.65 l=0.71
X6 VTAIL.t3 VN.t2 VDD2.t1 w_n1594_n3298# sky130_fd_pr__pfet_01v8 ad=4.5435 pd=24.08 as=1.92225 ps=11.98 w=11.65 l=0.71
X7 B.t5 B.t3 B.t4 w_n1594_n3298# sky130_fd_pr__pfet_01v8 ad=4.5435 pd=24.08 as=0 ps=0 w=11.65 l=0.71
X8 VDD2.t0 VN.t3 VTAIL.t2 w_n1594_n3298# sky130_fd_pr__pfet_01v8 ad=1.92225 pd=11.98 as=4.5435 ps=24.08 w=11.65 l=0.71
X9 B.t2 B.t0 B.t1 w_n1594_n3298# sky130_fd_pr__pfet_01v8 ad=4.5435 pd=24.08 as=0 ps=0 w=11.65 l=0.71
X10 VDD1.t1 VP.t2 VTAIL.t6 w_n1594_n3298# sky130_fd_pr__pfet_01v8 ad=1.92225 pd=11.98 as=4.5435 ps=24.08 w=11.65 l=0.71
X11 VTAIL.t7 VP.t3 VDD1.t0 w_n1594_n3298# sky130_fd_pr__pfet_01v8 ad=4.5435 pd=24.08 as=1.92225 ps=11.98 w=11.65 l=0.71
R0 VP.n1 VP.t1 472.108
R1 VP.n1 VP.t0 472.058
R2 VP.n3 VP.t3 451.111
R3 VP.n5 VP.t2 451.111
R4 VP.n6 VP.n5 161.3
R5 VP.n4 VP.n0 161.3
R6 VP.n3 VP.n2 161.3
R7 VP.n2 VP.n1 84.8439
R8 VP.n4 VP.n3 24.1005
R9 VP.n5 VP.n4 24.1005
R10 VP.n2 VP.n0 0.189894
R11 VP.n6 VP.n0 0.189894
R12 VP VP.n6 0.0516364
R13 VTAIL.n5 VTAIL.t4 58.2729
R14 VTAIL.n4 VTAIL.t0 58.2729
R15 VTAIL.n3 VTAIL.t1 58.2729
R16 VTAIL.n7 VTAIL.t2 58.2727
R17 VTAIL.n0 VTAIL.t3 58.2727
R18 VTAIL.n1 VTAIL.t6 58.2727
R19 VTAIL.n2 VTAIL.t7 58.2727
R20 VTAIL.n6 VTAIL.t5 58.2727
R21 VTAIL.n7 VTAIL.n6 23.3065
R22 VTAIL.n3 VTAIL.n2 23.3065
R23 VTAIL.n4 VTAIL.n3 0.897052
R24 VTAIL.n6 VTAIL.n5 0.897052
R25 VTAIL.n2 VTAIL.n1 0.897052
R26 VTAIL VTAIL.n0 0.506965
R27 VTAIL.n5 VTAIL.n4 0.470328
R28 VTAIL.n1 VTAIL.n0 0.470328
R29 VTAIL VTAIL.n7 0.390586
R30 VDD1 VDD1.n1 109.133
R31 VDD1 VDD1.n0 72.2196
R32 VDD1.n0 VDD1.t2 2.79063
R33 VDD1.n0 VDD1.t3 2.79063
R34 VDD1.n1 VDD1.t0 2.79063
R35 VDD1.n1 VDD1.t1 2.79063
R36 VN.n0 VN.t2 472.108
R37 VN.n1 VN.t1 472.108
R38 VN.n0 VN.t3 472.058
R39 VN.n1 VN.t0 472.058
R40 VN VN.n1 85.2246
R41 VN VN.n0 44.7132
R42 VDD2.n2 VDD2.n0 108.609
R43 VDD2.n2 VDD2.n1 72.1614
R44 VDD2.n1 VDD2.t3 2.79063
R45 VDD2.n1 VDD2.t2 2.79063
R46 VDD2.n0 VDD2.t1 2.79063
R47 VDD2.n0 VDD2.t0 2.79063
R48 VDD2 VDD2.n2 0.0586897
R49 B.n104 B.t0 598.288
R50 B.n232 B.t9 598.288
R51 B.n38 B.t6 598.288
R52 B.n32 B.t3 598.288
R53 B.n297 B.n78 585
R54 B.n296 B.n295 585
R55 B.n294 B.n79 585
R56 B.n293 B.n292 585
R57 B.n291 B.n80 585
R58 B.n290 B.n289 585
R59 B.n288 B.n81 585
R60 B.n287 B.n286 585
R61 B.n285 B.n82 585
R62 B.n284 B.n283 585
R63 B.n282 B.n83 585
R64 B.n281 B.n280 585
R65 B.n279 B.n84 585
R66 B.n278 B.n277 585
R67 B.n276 B.n85 585
R68 B.n275 B.n274 585
R69 B.n273 B.n86 585
R70 B.n272 B.n271 585
R71 B.n270 B.n87 585
R72 B.n269 B.n268 585
R73 B.n267 B.n88 585
R74 B.n266 B.n265 585
R75 B.n264 B.n89 585
R76 B.n263 B.n262 585
R77 B.n261 B.n90 585
R78 B.n260 B.n259 585
R79 B.n258 B.n91 585
R80 B.n257 B.n256 585
R81 B.n255 B.n92 585
R82 B.n254 B.n253 585
R83 B.n252 B.n93 585
R84 B.n251 B.n250 585
R85 B.n249 B.n94 585
R86 B.n248 B.n247 585
R87 B.n246 B.n95 585
R88 B.n245 B.n244 585
R89 B.n243 B.n96 585
R90 B.n242 B.n241 585
R91 B.n240 B.n97 585
R92 B.n239 B.n238 585
R93 B.n237 B.n98 585
R94 B.n236 B.n235 585
R95 B.n231 B.n99 585
R96 B.n230 B.n229 585
R97 B.n228 B.n100 585
R98 B.n227 B.n226 585
R99 B.n225 B.n101 585
R100 B.n224 B.n223 585
R101 B.n222 B.n102 585
R102 B.n221 B.n220 585
R103 B.n218 B.n103 585
R104 B.n217 B.n216 585
R105 B.n215 B.n106 585
R106 B.n214 B.n213 585
R107 B.n212 B.n107 585
R108 B.n211 B.n210 585
R109 B.n209 B.n108 585
R110 B.n208 B.n207 585
R111 B.n206 B.n109 585
R112 B.n205 B.n204 585
R113 B.n203 B.n110 585
R114 B.n202 B.n201 585
R115 B.n200 B.n111 585
R116 B.n199 B.n198 585
R117 B.n197 B.n112 585
R118 B.n196 B.n195 585
R119 B.n194 B.n113 585
R120 B.n193 B.n192 585
R121 B.n191 B.n114 585
R122 B.n190 B.n189 585
R123 B.n188 B.n115 585
R124 B.n187 B.n186 585
R125 B.n185 B.n116 585
R126 B.n184 B.n183 585
R127 B.n182 B.n117 585
R128 B.n181 B.n180 585
R129 B.n179 B.n118 585
R130 B.n178 B.n177 585
R131 B.n176 B.n119 585
R132 B.n175 B.n174 585
R133 B.n173 B.n120 585
R134 B.n172 B.n171 585
R135 B.n170 B.n121 585
R136 B.n169 B.n168 585
R137 B.n167 B.n122 585
R138 B.n166 B.n165 585
R139 B.n164 B.n123 585
R140 B.n163 B.n162 585
R141 B.n161 B.n124 585
R142 B.n160 B.n159 585
R143 B.n158 B.n125 585
R144 B.n299 B.n298 585
R145 B.n300 B.n77 585
R146 B.n302 B.n301 585
R147 B.n303 B.n76 585
R148 B.n305 B.n304 585
R149 B.n306 B.n75 585
R150 B.n308 B.n307 585
R151 B.n309 B.n74 585
R152 B.n311 B.n310 585
R153 B.n312 B.n73 585
R154 B.n314 B.n313 585
R155 B.n315 B.n72 585
R156 B.n317 B.n316 585
R157 B.n318 B.n71 585
R158 B.n320 B.n319 585
R159 B.n321 B.n70 585
R160 B.n323 B.n322 585
R161 B.n324 B.n69 585
R162 B.n326 B.n325 585
R163 B.n327 B.n68 585
R164 B.n329 B.n328 585
R165 B.n330 B.n67 585
R166 B.n332 B.n331 585
R167 B.n333 B.n66 585
R168 B.n335 B.n334 585
R169 B.n336 B.n65 585
R170 B.n338 B.n337 585
R171 B.n339 B.n64 585
R172 B.n341 B.n340 585
R173 B.n342 B.n63 585
R174 B.n344 B.n343 585
R175 B.n345 B.n62 585
R176 B.n347 B.n346 585
R177 B.n348 B.n61 585
R178 B.n350 B.n349 585
R179 B.n351 B.n60 585
R180 B.n490 B.n489 585
R181 B.n488 B.n11 585
R182 B.n487 B.n486 585
R183 B.n485 B.n12 585
R184 B.n484 B.n483 585
R185 B.n482 B.n13 585
R186 B.n481 B.n480 585
R187 B.n479 B.n14 585
R188 B.n478 B.n477 585
R189 B.n476 B.n15 585
R190 B.n475 B.n474 585
R191 B.n473 B.n16 585
R192 B.n472 B.n471 585
R193 B.n470 B.n17 585
R194 B.n469 B.n468 585
R195 B.n467 B.n18 585
R196 B.n466 B.n465 585
R197 B.n464 B.n19 585
R198 B.n463 B.n462 585
R199 B.n461 B.n20 585
R200 B.n460 B.n459 585
R201 B.n458 B.n21 585
R202 B.n457 B.n456 585
R203 B.n455 B.n22 585
R204 B.n454 B.n453 585
R205 B.n452 B.n23 585
R206 B.n451 B.n450 585
R207 B.n449 B.n24 585
R208 B.n448 B.n447 585
R209 B.n446 B.n25 585
R210 B.n445 B.n444 585
R211 B.n443 B.n26 585
R212 B.n442 B.n441 585
R213 B.n440 B.n27 585
R214 B.n439 B.n438 585
R215 B.n437 B.n28 585
R216 B.n436 B.n435 585
R217 B.n434 B.n29 585
R218 B.n433 B.n432 585
R219 B.n431 B.n30 585
R220 B.n430 B.n429 585
R221 B.n427 B.n31 585
R222 B.n426 B.n425 585
R223 B.n424 B.n34 585
R224 B.n423 B.n422 585
R225 B.n421 B.n35 585
R226 B.n420 B.n419 585
R227 B.n418 B.n36 585
R228 B.n417 B.n416 585
R229 B.n415 B.n37 585
R230 B.n413 B.n412 585
R231 B.n411 B.n40 585
R232 B.n410 B.n409 585
R233 B.n408 B.n41 585
R234 B.n407 B.n406 585
R235 B.n405 B.n42 585
R236 B.n404 B.n403 585
R237 B.n402 B.n43 585
R238 B.n401 B.n400 585
R239 B.n399 B.n44 585
R240 B.n398 B.n397 585
R241 B.n396 B.n45 585
R242 B.n395 B.n394 585
R243 B.n393 B.n46 585
R244 B.n392 B.n391 585
R245 B.n390 B.n47 585
R246 B.n389 B.n388 585
R247 B.n387 B.n48 585
R248 B.n386 B.n385 585
R249 B.n384 B.n49 585
R250 B.n383 B.n382 585
R251 B.n381 B.n50 585
R252 B.n380 B.n379 585
R253 B.n378 B.n51 585
R254 B.n377 B.n376 585
R255 B.n375 B.n52 585
R256 B.n374 B.n373 585
R257 B.n372 B.n53 585
R258 B.n371 B.n370 585
R259 B.n369 B.n54 585
R260 B.n368 B.n367 585
R261 B.n366 B.n55 585
R262 B.n365 B.n364 585
R263 B.n363 B.n56 585
R264 B.n362 B.n361 585
R265 B.n360 B.n57 585
R266 B.n359 B.n358 585
R267 B.n357 B.n58 585
R268 B.n356 B.n355 585
R269 B.n354 B.n59 585
R270 B.n353 B.n352 585
R271 B.n491 B.n10 585
R272 B.n493 B.n492 585
R273 B.n494 B.n9 585
R274 B.n496 B.n495 585
R275 B.n497 B.n8 585
R276 B.n499 B.n498 585
R277 B.n500 B.n7 585
R278 B.n502 B.n501 585
R279 B.n503 B.n6 585
R280 B.n505 B.n504 585
R281 B.n506 B.n5 585
R282 B.n508 B.n507 585
R283 B.n509 B.n4 585
R284 B.n511 B.n510 585
R285 B.n512 B.n3 585
R286 B.n514 B.n513 585
R287 B.n515 B.n0 585
R288 B.n2 B.n1 585
R289 B.n134 B.n133 585
R290 B.n136 B.n135 585
R291 B.n137 B.n132 585
R292 B.n139 B.n138 585
R293 B.n140 B.n131 585
R294 B.n142 B.n141 585
R295 B.n143 B.n130 585
R296 B.n145 B.n144 585
R297 B.n146 B.n129 585
R298 B.n148 B.n147 585
R299 B.n149 B.n128 585
R300 B.n151 B.n150 585
R301 B.n152 B.n127 585
R302 B.n154 B.n153 585
R303 B.n155 B.n126 585
R304 B.n157 B.n156 585
R305 B.n156 B.n125 444.452
R306 B.n298 B.n297 444.452
R307 B.n352 B.n351 444.452
R308 B.n491 B.n490 444.452
R309 B.n517 B.n516 256.663
R310 B.n516 B.n515 235.042
R311 B.n516 B.n2 235.042
R312 B.n160 B.n125 163.367
R313 B.n161 B.n160 163.367
R314 B.n162 B.n161 163.367
R315 B.n162 B.n123 163.367
R316 B.n166 B.n123 163.367
R317 B.n167 B.n166 163.367
R318 B.n168 B.n167 163.367
R319 B.n168 B.n121 163.367
R320 B.n172 B.n121 163.367
R321 B.n173 B.n172 163.367
R322 B.n174 B.n173 163.367
R323 B.n174 B.n119 163.367
R324 B.n178 B.n119 163.367
R325 B.n179 B.n178 163.367
R326 B.n180 B.n179 163.367
R327 B.n180 B.n117 163.367
R328 B.n184 B.n117 163.367
R329 B.n185 B.n184 163.367
R330 B.n186 B.n185 163.367
R331 B.n186 B.n115 163.367
R332 B.n190 B.n115 163.367
R333 B.n191 B.n190 163.367
R334 B.n192 B.n191 163.367
R335 B.n192 B.n113 163.367
R336 B.n196 B.n113 163.367
R337 B.n197 B.n196 163.367
R338 B.n198 B.n197 163.367
R339 B.n198 B.n111 163.367
R340 B.n202 B.n111 163.367
R341 B.n203 B.n202 163.367
R342 B.n204 B.n203 163.367
R343 B.n204 B.n109 163.367
R344 B.n208 B.n109 163.367
R345 B.n209 B.n208 163.367
R346 B.n210 B.n209 163.367
R347 B.n210 B.n107 163.367
R348 B.n214 B.n107 163.367
R349 B.n215 B.n214 163.367
R350 B.n216 B.n215 163.367
R351 B.n216 B.n103 163.367
R352 B.n221 B.n103 163.367
R353 B.n222 B.n221 163.367
R354 B.n223 B.n222 163.367
R355 B.n223 B.n101 163.367
R356 B.n227 B.n101 163.367
R357 B.n228 B.n227 163.367
R358 B.n229 B.n228 163.367
R359 B.n229 B.n99 163.367
R360 B.n236 B.n99 163.367
R361 B.n237 B.n236 163.367
R362 B.n238 B.n237 163.367
R363 B.n238 B.n97 163.367
R364 B.n242 B.n97 163.367
R365 B.n243 B.n242 163.367
R366 B.n244 B.n243 163.367
R367 B.n244 B.n95 163.367
R368 B.n248 B.n95 163.367
R369 B.n249 B.n248 163.367
R370 B.n250 B.n249 163.367
R371 B.n250 B.n93 163.367
R372 B.n254 B.n93 163.367
R373 B.n255 B.n254 163.367
R374 B.n256 B.n255 163.367
R375 B.n256 B.n91 163.367
R376 B.n260 B.n91 163.367
R377 B.n261 B.n260 163.367
R378 B.n262 B.n261 163.367
R379 B.n262 B.n89 163.367
R380 B.n266 B.n89 163.367
R381 B.n267 B.n266 163.367
R382 B.n268 B.n267 163.367
R383 B.n268 B.n87 163.367
R384 B.n272 B.n87 163.367
R385 B.n273 B.n272 163.367
R386 B.n274 B.n273 163.367
R387 B.n274 B.n85 163.367
R388 B.n278 B.n85 163.367
R389 B.n279 B.n278 163.367
R390 B.n280 B.n279 163.367
R391 B.n280 B.n83 163.367
R392 B.n284 B.n83 163.367
R393 B.n285 B.n284 163.367
R394 B.n286 B.n285 163.367
R395 B.n286 B.n81 163.367
R396 B.n290 B.n81 163.367
R397 B.n291 B.n290 163.367
R398 B.n292 B.n291 163.367
R399 B.n292 B.n79 163.367
R400 B.n296 B.n79 163.367
R401 B.n297 B.n296 163.367
R402 B.n351 B.n350 163.367
R403 B.n350 B.n61 163.367
R404 B.n346 B.n61 163.367
R405 B.n346 B.n345 163.367
R406 B.n345 B.n344 163.367
R407 B.n344 B.n63 163.367
R408 B.n340 B.n63 163.367
R409 B.n340 B.n339 163.367
R410 B.n339 B.n338 163.367
R411 B.n338 B.n65 163.367
R412 B.n334 B.n65 163.367
R413 B.n334 B.n333 163.367
R414 B.n333 B.n332 163.367
R415 B.n332 B.n67 163.367
R416 B.n328 B.n67 163.367
R417 B.n328 B.n327 163.367
R418 B.n327 B.n326 163.367
R419 B.n326 B.n69 163.367
R420 B.n322 B.n69 163.367
R421 B.n322 B.n321 163.367
R422 B.n321 B.n320 163.367
R423 B.n320 B.n71 163.367
R424 B.n316 B.n71 163.367
R425 B.n316 B.n315 163.367
R426 B.n315 B.n314 163.367
R427 B.n314 B.n73 163.367
R428 B.n310 B.n73 163.367
R429 B.n310 B.n309 163.367
R430 B.n309 B.n308 163.367
R431 B.n308 B.n75 163.367
R432 B.n304 B.n75 163.367
R433 B.n304 B.n303 163.367
R434 B.n303 B.n302 163.367
R435 B.n302 B.n77 163.367
R436 B.n298 B.n77 163.367
R437 B.n490 B.n11 163.367
R438 B.n486 B.n11 163.367
R439 B.n486 B.n485 163.367
R440 B.n485 B.n484 163.367
R441 B.n484 B.n13 163.367
R442 B.n480 B.n13 163.367
R443 B.n480 B.n479 163.367
R444 B.n479 B.n478 163.367
R445 B.n478 B.n15 163.367
R446 B.n474 B.n15 163.367
R447 B.n474 B.n473 163.367
R448 B.n473 B.n472 163.367
R449 B.n472 B.n17 163.367
R450 B.n468 B.n17 163.367
R451 B.n468 B.n467 163.367
R452 B.n467 B.n466 163.367
R453 B.n466 B.n19 163.367
R454 B.n462 B.n19 163.367
R455 B.n462 B.n461 163.367
R456 B.n461 B.n460 163.367
R457 B.n460 B.n21 163.367
R458 B.n456 B.n21 163.367
R459 B.n456 B.n455 163.367
R460 B.n455 B.n454 163.367
R461 B.n454 B.n23 163.367
R462 B.n450 B.n23 163.367
R463 B.n450 B.n449 163.367
R464 B.n449 B.n448 163.367
R465 B.n448 B.n25 163.367
R466 B.n444 B.n25 163.367
R467 B.n444 B.n443 163.367
R468 B.n443 B.n442 163.367
R469 B.n442 B.n27 163.367
R470 B.n438 B.n27 163.367
R471 B.n438 B.n437 163.367
R472 B.n437 B.n436 163.367
R473 B.n436 B.n29 163.367
R474 B.n432 B.n29 163.367
R475 B.n432 B.n431 163.367
R476 B.n431 B.n430 163.367
R477 B.n430 B.n31 163.367
R478 B.n425 B.n31 163.367
R479 B.n425 B.n424 163.367
R480 B.n424 B.n423 163.367
R481 B.n423 B.n35 163.367
R482 B.n419 B.n35 163.367
R483 B.n419 B.n418 163.367
R484 B.n418 B.n417 163.367
R485 B.n417 B.n37 163.367
R486 B.n412 B.n37 163.367
R487 B.n412 B.n411 163.367
R488 B.n411 B.n410 163.367
R489 B.n410 B.n41 163.367
R490 B.n406 B.n41 163.367
R491 B.n406 B.n405 163.367
R492 B.n405 B.n404 163.367
R493 B.n404 B.n43 163.367
R494 B.n400 B.n43 163.367
R495 B.n400 B.n399 163.367
R496 B.n399 B.n398 163.367
R497 B.n398 B.n45 163.367
R498 B.n394 B.n45 163.367
R499 B.n394 B.n393 163.367
R500 B.n393 B.n392 163.367
R501 B.n392 B.n47 163.367
R502 B.n388 B.n47 163.367
R503 B.n388 B.n387 163.367
R504 B.n387 B.n386 163.367
R505 B.n386 B.n49 163.367
R506 B.n382 B.n49 163.367
R507 B.n382 B.n381 163.367
R508 B.n381 B.n380 163.367
R509 B.n380 B.n51 163.367
R510 B.n376 B.n51 163.367
R511 B.n376 B.n375 163.367
R512 B.n375 B.n374 163.367
R513 B.n374 B.n53 163.367
R514 B.n370 B.n53 163.367
R515 B.n370 B.n369 163.367
R516 B.n369 B.n368 163.367
R517 B.n368 B.n55 163.367
R518 B.n364 B.n55 163.367
R519 B.n364 B.n363 163.367
R520 B.n363 B.n362 163.367
R521 B.n362 B.n57 163.367
R522 B.n358 B.n57 163.367
R523 B.n358 B.n357 163.367
R524 B.n357 B.n356 163.367
R525 B.n356 B.n59 163.367
R526 B.n352 B.n59 163.367
R527 B.n492 B.n491 163.367
R528 B.n492 B.n9 163.367
R529 B.n496 B.n9 163.367
R530 B.n497 B.n496 163.367
R531 B.n498 B.n497 163.367
R532 B.n498 B.n7 163.367
R533 B.n502 B.n7 163.367
R534 B.n503 B.n502 163.367
R535 B.n504 B.n503 163.367
R536 B.n504 B.n5 163.367
R537 B.n508 B.n5 163.367
R538 B.n509 B.n508 163.367
R539 B.n510 B.n509 163.367
R540 B.n510 B.n3 163.367
R541 B.n514 B.n3 163.367
R542 B.n515 B.n514 163.367
R543 B.n133 B.n2 163.367
R544 B.n136 B.n133 163.367
R545 B.n137 B.n136 163.367
R546 B.n138 B.n137 163.367
R547 B.n138 B.n131 163.367
R548 B.n142 B.n131 163.367
R549 B.n143 B.n142 163.367
R550 B.n144 B.n143 163.367
R551 B.n144 B.n129 163.367
R552 B.n148 B.n129 163.367
R553 B.n149 B.n148 163.367
R554 B.n150 B.n149 163.367
R555 B.n150 B.n127 163.367
R556 B.n154 B.n127 163.367
R557 B.n155 B.n154 163.367
R558 B.n156 B.n155 163.367
R559 B.n232 B.t10 129.103
R560 B.n38 B.t8 129.103
R561 B.n104 B.t1 129.089
R562 B.n32 B.t5 129.089
R563 B.n233 B.t11 108.933
R564 B.n39 B.t7 108.933
R565 B.n105 B.t2 108.919
R566 B.n33 B.t4 108.919
R567 B.n219 B.n105 59.5399
R568 B.n234 B.n233 59.5399
R569 B.n414 B.n39 59.5399
R570 B.n428 B.n33 59.5399
R571 B.n489 B.n10 28.8785
R572 B.n353 B.n60 28.8785
R573 B.n158 B.n157 28.8785
R574 B.n299 B.n78 28.8785
R575 B.n105 B.n104 20.1702
R576 B.n233 B.n232 20.1702
R577 B.n39 B.n38 20.1702
R578 B.n33 B.n32 20.1702
R579 B B.n517 18.0485
R580 B.n493 B.n10 10.6151
R581 B.n494 B.n493 10.6151
R582 B.n495 B.n494 10.6151
R583 B.n495 B.n8 10.6151
R584 B.n499 B.n8 10.6151
R585 B.n500 B.n499 10.6151
R586 B.n501 B.n500 10.6151
R587 B.n501 B.n6 10.6151
R588 B.n505 B.n6 10.6151
R589 B.n506 B.n505 10.6151
R590 B.n507 B.n506 10.6151
R591 B.n507 B.n4 10.6151
R592 B.n511 B.n4 10.6151
R593 B.n512 B.n511 10.6151
R594 B.n513 B.n512 10.6151
R595 B.n513 B.n0 10.6151
R596 B.n489 B.n488 10.6151
R597 B.n488 B.n487 10.6151
R598 B.n487 B.n12 10.6151
R599 B.n483 B.n12 10.6151
R600 B.n483 B.n482 10.6151
R601 B.n482 B.n481 10.6151
R602 B.n481 B.n14 10.6151
R603 B.n477 B.n14 10.6151
R604 B.n477 B.n476 10.6151
R605 B.n476 B.n475 10.6151
R606 B.n475 B.n16 10.6151
R607 B.n471 B.n16 10.6151
R608 B.n471 B.n470 10.6151
R609 B.n470 B.n469 10.6151
R610 B.n469 B.n18 10.6151
R611 B.n465 B.n18 10.6151
R612 B.n465 B.n464 10.6151
R613 B.n464 B.n463 10.6151
R614 B.n463 B.n20 10.6151
R615 B.n459 B.n20 10.6151
R616 B.n459 B.n458 10.6151
R617 B.n458 B.n457 10.6151
R618 B.n457 B.n22 10.6151
R619 B.n453 B.n22 10.6151
R620 B.n453 B.n452 10.6151
R621 B.n452 B.n451 10.6151
R622 B.n451 B.n24 10.6151
R623 B.n447 B.n24 10.6151
R624 B.n447 B.n446 10.6151
R625 B.n446 B.n445 10.6151
R626 B.n445 B.n26 10.6151
R627 B.n441 B.n26 10.6151
R628 B.n441 B.n440 10.6151
R629 B.n440 B.n439 10.6151
R630 B.n439 B.n28 10.6151
R631 B.n435 B.n28 10.6151
R632 B.n435 B.n434 10.6151
R633 B.n434 B.n433 10.6151
R634 B.n433 B.n30 10.6151
R635 B.n429 B.n30 10.6151
R636 B.n427 B.n426 10.6151
R637 B.n426 B.n34 10.6151
R638 B.n422 B.n34 10.6151
R639 B.n422 B.n421 10.6151
R640 B.n421 B.n420 10.6151
R641 B.n420 B.n36 10.6151
R642 B.n416 B.n36 10.6151
R643 B.n416 B.n415 10.6151
R644 B.n413 B.n40 10.6151
R645 B.n409 B.n40 10.6151
R646 B.n409 B.n408 10.6151
R647 B.n408 B.n407 10.6151
R648 B.n407 B.n42 10.6151
R649 B.n403 B.n42 10.6151
R650 B.n403 B.n402 10.6151
R651 B.n402 B.n401 10.6151
R652 B.n401 B.n44 10.6151
R653 B.n397 B.n44 10.6151
R654 B.n397 B.n396 10.6151
R655 B.n396 B.n395 10.6151
R656 B.n395 B.n46 10.6151
R657 B.n391 B.n46 10.6151
R658 B.n391 B.n390 10.6151
R659 B.n390 B.n389 10.6151
R660 B.n389 B.n48 10.6151
R661 B.n385 B.n48 10.6151
R662 B.n385 B.n384 10.6151
R663 B.n384 B.n383 10.6151
R664 B.n383 B.n50 10.6151
R665 B.n379 B.n50 10.6151
R666 B.n379 B.n378 10.6151
R667 B.n378 B.n377 10.6151
R668 B.n377 B.n52 10.6151
R669 B.n373 B.n52 10.6151
R670 B.n373 B.n372 10.6151
R671 B.n372 B.n371 10.6151
R672 B.n371 B.n54 10.6151
R673 B.n367 B.n54 10.6151
R674 B.n367 B.n366 10.6151
R675 B.n366 B.n365 10.6151
R676 B.n365 B.n56 10.6151
R677 B.n361 B.n56 10.6151
R678 B.n361 B.n360 10.6151
R679 B.n360 B.n359 10.6151
R680 B.n359 B.n58 10.6151
R681 B.n355 B.n58 10.6151
R682 B.n355 B.n354 10.6151
R683 B.n354 B.n353 10.6151
R684 B.n349 B.n60 10.6151
R685 B.n349 B.n348 10.6151
R686 B.n348 B.n347 10.6151
R687 B.n347 B.n62 10.6151
R688 B.n343 B.n62 10.6151
R689 B.n343 B.n342 10.6151
R690 B.n342 B.n341 10.6151
R691 B.n341 B.n64 10.6151
R692 B.n337 B.n64 10.6151
R693 B.n337 B.n336 10.6151
R694 B.n336 B.n335 10.6151
R695 B.n335 B.n66 10.6151
R696 B.n331 B.n66 10.6151
R697 B.n331 B.n330 10.6151
R698 B.n330 B.n329 10.6151
R699 B.n329 B.n68 10.6151
R700 B.n325 B.n68 10.6151
R701 B.n325 B.n324 10.6151
R702 B.n324 B.n323 10.6151
R703 B.n323 B.n70 10.6151
R704 B.n319 B.n70 10.6151
R705 B.n319 B.n318 10.6151
R706 B.n318 B.n317 10.6151
R707 B.n317 B.n72 10.6151
R708 B.n313 B.n72 10.6151
R709 B.n313 B.n312 10.6151
R710 B.n312 B.n311 10.6151
R711 B.n311 B.n74 10.6151
R712 B.n307 B.n74 10.6151
R713 B.n307 B.n306 10.6151
R714 B.n306 B.n305 10.6151
R715 B.n305 B.n76 10.6151
R716 B.n301 B.n76 10.6151
R717 B.n301 B.n300 10.6151
R718 B.n300 B.n299 10.6151
R719 B.n134 B.n1 10.6151
R720 B.n135 B.n134 10.6151
R721 B.n135 B.n132 10.6151
R722 B.n139 B.n132 10.6151
R723 B.n140 B.n139 10.6151
R724 B.n141 B.n140 10.6151
R725 B.n141 B.n130 10.6151
R726 B.n145 B.n130 10.6151
R727 B.n146 B.n145 10.6151
R728 B.n147 B.n146 10.6151
R729 B.n147 B.n128 10.6151
R730 B.n151 B.n128 10.6151
R731 B.n152 B.n151 10.6151
R732 B.n153 B.n152 10.6151
R733 B.n153 B.n126 10.6151
R734 B.n157 B.n126 10.6151
R735 B.n159 B.n158 10.6151
R736 B.n159 B.n124 10.6151
R737 B.n163 B.n124 10.6151
R738 B.n164 B.n163 10.6151
R739 B.n165 B.n164 10.6151
R740 B.n165 B.n122 10.6151
R741 B.n169 B.n122 10.6151
R742 B.n170 B.n169 10.6151
R743 B.n171 B.n170 10.6151
R744 B.n171 B.n120 10.6151
R745 B.n175 B.n120 10.6151
R746 B.n176 B.n175 10.6151
R747 B.n177 B.n176 10.6151
R748 B.n177 B.n118 10.6151
R749 B.n181 B.n118 10.6151
R750 B.n182 B.n181 10.6151
R751 B.n183 B.n182 10.6151
R752 B.n183 B.n116 10.6151
R753 B.n187 B.n116 10.6151
R754 B.n188 B.n187 10.6151
R755 B.n189 B.n188 10.6151
R756 B.n189 B.n114 10.6151
R757 B.n193 B.n114 10.6151
R758 B.n194 B.n193 10.6151
R759 B.n195 B.n194 10.6151
R760 B.n195 B.n112 10.6151
R761 B.n199 B.n112 10.6151
R762 B.n200 B.n199 10.6151
R763 B.n201 B.n200 10.6151
R764 B.n201 B.n110 10.6151
R765 B.n205 B.n110 10.6151
R766 B.n206 B.n205 10.6151
R767 B.n207 B.n206 10.6151
R768 B.n207 B.n108 10.6151
R769 B.n211 B.n108 10.6151
R770 B.n212 B.n211 10.6151
R771 B.n213 B.n212 10.6151
R772 B.n213 B.n106 10.6151
R773 B.n217 B.n106 10.6151
R774 B.n218 B.n217 10.6151
R775 B.n220 B.n102 10.6151
R776 B.n224 B.n102 10.6151
R777 B.n225 B.n224 10.6151
R778 B.n226 B.n225 10.6151
R779 B.n226 B.n100 10.6151
R780 B.n230 B.n100 10.6151
R781 B.n231 B.n230 10.6151
R782 B.n235 B.n231 10.6151
R783 B.n239 B.n98 10.6151
R784 B.n240 B.n239 10.6151
R785 B.n241 B.n240 10.6151
R786 B.n241 B.n96 10.6151
R787 B.n245 B.n96 10.6151
R788 B.n246 B.n245 10.6151
R789 B.n247 B.n246 10.6151
R790 B.n247 B.n94 10.6151
R791 B.n251 B.n94 10.6151
R792 B.n252 B.n251 10.6151
R793 B.n253 B.n252 10.6151
R794 B.n253 B.n92 10.6151
R795 B.n257 B.n92 10.6151
R796 B.n258 B.n257 10.6151
R797 B.n259 B.n258 10.6151
R798 B.n259 B.n90 10.6151
R799 B.n263 B.n90 10.6151
R800 B.n264 B.n263 10.6151
R801 B.n265 B.n264 10.6151
R802 B.n265 B.n88 10.6151
R803 B.n269 B.n88 10.6151
R804 B.n270 B.n269 10.6151
R805 B.n271 B.n270 10.6151
R806 B.n271 B.n86 10.6151
R807 B.n275 B.n86 10.6151
R808 B.n276 B.n275 10.6151
R809 B.n277 B.n276 10.6151
R810 B.n277 B.n84 10.6151
R811 B.n281 B.n84 10.6151
R812 B.n282 B.n281 10.6151
R813 B.n283 B.n282 10.6151
R814 B.n283 B.n82 10.6151
R815 B.n287 B.n82 10.6151
R816 B.n288 B.n287 10.6151
R817 B.n289 B.n288 10.6151
R818 B.n289 B.n80 10.6151
R819 B.n293 B.n80 10.6151
R820 B.n294 B.n293 10.6151
R821 B.n295 B.n294 10.6151
R822 B.n295 B.n78 10.6151
R823 B.n517 B.n0 8.11757
R824 B.n517 B.n1 8.11757
R825 B.n428 B.n427 6.5566
R826 B.n415 B.n414 6.5566
R827 B.n220 B.n219 6.5566
R828 B.n235 B.n234 6.5566
R829 B.n429 B.n428 4.05904
R830 B.n414 B.n413 4.05904
R831 B.n219 B.n218 4.05904
R832 B.n234 B.n98 4.05904
C0 VDD2 B 0.940107f
C1 w_n1594_n3298# VN 2.35062f
C2 VN VP 4.76606f
C3 VDD2 w_n1594_n3298# 1.06857f
C4 VTAIL VDD1 6.60083f
C5 VDD2 VP 0.273848f
C6 B w_n1594_n3298# 6.82176f
C7 B VP 1.06751f
C8 VDD1 VN 0.147098f
C9 w_n1594_n3298# VP 2.55076f
C10 VTAIL VN 2.71827f
C11 VDD2 VDD1 0.568716f
C12 VDD2 VTAIL 6.64236f
C13 B VDD1 0.91843f
C14 B VTAIL 3.72971f
C15 w_n1594_n3298# VDD1 1.05386f
C16 VDD2 VN 3.09778f
C17 VDD1 VP 3.22427f
C18 VTAIL w_n1594_n3298# 4.03037f
C19 VTAIL VP 2.73237f
C20 B VN 0.744189f
C21 VDD2 VSUBS 0.668517f
C22 VDD1 VSUBS 4.893106f
C23 VTAIL VSUBS 0.852293f
C24 VN VSUBS 5.7222f
C25 VP VSUBS 1.282035f
C26 B VSUBS 2.598994f
C27 w_n1594_n3298# VSUBS 64.74831f
C28 B.n0 VSUBS 0.007233f
C29 B.n1 VSUBS 0.007233f
C30 B.n2 VSUBS 0.010697f
C31 B.n3 VSUBS 0.008197f
C32 B.n4 VSUBS 0.008197f
C33 B.n5 VSUBS 0.008197f
C34 B.n6 VSUBS 0.008197f
C35 B.n7 VSUBS 0.008197f
C36 B.n8 VSUBS 0.008197f
C37 B.n9 VSUBS 0.008197f
C38 B.n10 VSUBS 0.01728f
C39 B.n11 VSUBS 0.008197f
C40 B.n12 VSUBS 0.008197f
C41 B.n13 VSUBS 0.008197f
C42 B.n14 VSUBS 0.008197f
C43 B.n15 VSUBS 0.008197f
C44 B.n16 VSUBS 0.008197f
C45 B.n17 VSUBS 0.008197f
C46 B.n18 VSUBS 0.008197f
C47 B.n19 VSUBS 0.008197f
C48 B.n20 VSUBS 0.008197f
C49 B.n21 VSUBS 0.008197f
C50 B.n22 VSUBS 0.008197f
C51 B.n23 VSUBS 0.008197f
C52 B.n24 VSUBS 0.008197f
C53 B.n25 VSUBS 0.008197f
C54 B.n26 VSUBS 0.008197f
C55 B.n27 VSUBS 0.008197f
C56 B.n28 VSUBS 0.008197f
C57 B.n29 VSUBS 0.008197f
C58 B.n30 VSUBS 0.008197f
C59 B.n31 VSUBS 0.008197f
C60 B.t4 VSUBS 0.443159f
C61 B.t5 VSUBS 0.453032f
C62 B.t3 VSUBS 0.400671f
C63 B.n32 VSUBS 0.155538f
C64 B.n33 VSUBS 0.074881f
C65 B.n34 VSUBS 0.008197f
C66 B.n35 VSUBS 0.008197f
C67 B.n36 VSUBS 0.008197f
C68 B.n37 VSUBS 0.008197f
C69 B.t7 VSUBS 0.443151f
C70 B.t8 VSUBS 0.453024f
C71 B.t6 VSUBS 0.400671f
C72 B.n38 VSUBS 0.155546f
C73 B.n39 VSUBS 0.074889f
C74 B.n40 VSUBS 0.008197f
C75 B.n41 VSUBS 0.008197f
C76 B.n42 VSUBS 0.008197f
C77 B.n43 VSUBS 0.008197f
C78 B.n44 VSUBS 0.008197f
C79 B.n45 VSUBS 0.008197f
C80 B.n46 VSUBS 0.008197f
C81 B.n47 VSUBS 0.008197f
C82 B.n48 VSUBS 0.008197f
C83 B.n49 VSUBS 0.008197f
C84 B.n50 VSUBS 0.008197f
C85 B.n51 VSUBS 0.008197f
C86 B.n52 VSUBS 0.008197f
C87 B.n53 VSUBS 0.008197f
C88 B.n54 VSUBS 0.008197f
C89 B.n55 VSUBS 0.008197f
C90 B.n56 VSUBS 0.008197f
C91 B.n57 VSUBS 0.008197f
C92 B.n58 VSUBS 0.008197f
C93 B.n59 VSUBS 0.008197f
C94 B.n60 VSUBS 0.01728f
C95 B.n61 VSUBS 0.008197f
C96 B.n62 VSUBS 0.008197f
C97 B.n63 VSUBS 0.008197f
C98 B.n64 VSUBS 0.008197f
C99 B.n65 VSUBS 0.008197f
C100 B.n66 VSUBS 0.008197f
C101 B.n67 VSUBS 0.008197f
C102 B.n68 VSUBS 0.008197f
C103 B.n69 VSUBS 0.008197f
C104 B.n70 VSUBS 0.008197f
C105 B.n71 VSUBS 0.008197f
C106 B.n72 VSUBS 0.008197f
C107 B.n73 VSUBS 0.008197f
C108 B.n74 VSUBS 0.008197f
C109 B.n75 VSUBS 0.008197f
C110 B.n76 VSUBS 0.008197f
C111 B.n77 VSUBS 0.008197f
C112 B.n78 VSUBS 0.017066f
C113 B.n79 VSUBS 0.008197f
C114 B.n80 VSUBS 0.008197f
C115 B.n81 VSUBS 0.008197f
C116 B.n82 VSUBS 0.008197f
C117 B.n83 VSUBS 0.008197f
C118 B.n84 VSUBS 0.008197f
C119 B.n85 VSUBS 0.008197f
C120 B.n86 VSUBS 0.008197f
C121 B.n87 VSUBS 0.008197f
C122 B.n88 VSUBS 0.008197f
C123 B.n89 VSUBS 0.008197f
C124 B.n90 VSUBS 0.008197f
C125 B.n91 VSUBS 0.008197f
C126 B.n92 VSUBS 0.008197f
C127 B.n93 VSUBS 0.008197f
C128 B.n94 VSUBS 0.008197f
C129 B.n95 VSUBS 0.008197f
C130 B.n96 VSUBS 0.008197f
C131 B.n97 VSUBS 0.008197f
C132 B.n98 VSUBS 0.005666f
C133 B.n99 VSUBS 0.008197f
C134 B.n100 VSUBS 0.008197f
C135 B.n101 VSUBS 0.008197f
C136 B.n102 VSUBS 0.008197f
C137 B.n103 VSUBS 0.008197f
C138 B.t2 VSUBS 0.443159f
C139 B.t1 VSUBS 0.453032f
C140 B.t0 VSUBS 0.400671f
C141 B.n104 VSUBS 0.155538f
C142 B.n105 VSUBS 0.074881f
C143 B.n106 VSUBS 0.008197f
C144 B.n107 VSUBS 0.008197f
C145 B.n108 VSUBS 0.008197f
C146 B.n109 VSUBS 0.008197f
C147 B.n110 VSUBS 0.008197f
C148 B.n111 VSUBS 0.008197f
C149 B.n112 VSUBS 0.008197f
C150 B.n113 VSUBS 0.008197f
C151 B.n114 VSUBS 0.008197f
C152 B.n115 VSUBS 0.008197f
C153 B.n116 VSUBS 0.008197f
C154 B.n117 VSUBS 0.008197f
C155 B.n118 VSUBS 0.008197f
C156 B.n119 VSUBS 0.008197f
C157 B.n120 VSUBS 0.008197f
C158 B.n121 VSUBS 0.008197f
C159 B.n122 VSUBS 0.008197f
C160 B.n123 VSUBS 0.008197f
C161 B.n124 VSUBS 0.008197f
C162 B.n125 VSUBS 0.018161f
C163 B.n126 VSUBS 0.008197f
C164 B.n127 VSUBS 0.008197f
C165 B.n128 VSUBS 0.008197f
C166 B.n129 VSUBS 0.008197f
C167 B.n130 VSUBS 0.008197f
C168 B.n131 VSUBS 0.008197f
C169 B.n132 VSUBS 0.008197f
C170 B.n133 VSUBS 0.008197f
C171 B.n134 VSUBS 0.008197f
C172 B.n135 VSUBS 0.008197f
C173 B.n136 VSUBS 0.008197f
C174 B.n137 VSUBS 0.008197f
C175 B.n138 VSUBS 0.008197f
C176 B.n139 VSUBS 0.008197f
C177 B.n140 VSUBS 0.008197f
C178 B.n141 VSUBS 0.008197f
C179 B.n142 VSUBS 0.008197f
C180 B.n143 VSUBS 0.008197f
C181 B.n144 VSUBS 0.008197f
C182 B.n145 VSUBS 0.008197f
C183 B.n146 VSUBS 0.008197f
C184 B.n147 VSUBS 0.008197f
C185 B.n148 VSUBS 0.008197f
C186 B.n149 VSUBS 0.008197f
C187 B.n150 VSUBS 0.008197f
C188 B.n151 VSUBS 0.008197f
C189 B.n152 VSUBS 0.008197f
C190 B.n153 VSUBS 0.008197f
C191 B.n154 VSUBS 0.008197f
C192 B.n155 VSUBS 0.008197f
C193 B.n156 VSUBS 0.01728f
C194 B.n157 VSUBS 0.01728f
C195 B.n158 VSUBS 0.018161f
C196 B.n159 VSUBS 0.008197f
C197 B.n160 VSUBS 0.008197f
C198 B.n161 VSUBS 0.008197f
C199 B.n162 VSUBS 0.008197f
C200 B.n163 VSUBS 0.008197f
C201 B.n164 VSUBS 0.008197f
C202 B.n165 VSUBS 0.008197f
C203 B.n166 VSUBS 0.008197f
C204 B.n167 VSUBS 0.008197f
C205 B.n168 VSUBS 0.008197f
C206 B.n169 VSUBS 0.008197f
C207 B.n170 VSUBS 0.008197f
C208 B.n171 VSUBS 0.008197f
C209 B.n172 VSUBS 0.008197f
C210 B.n173 VSUBS 0.008197f
C211 B.n174 VSUBS 0.008197f
C212 B.n175 VSUBS 0.008197f
C213 B.n176 VSUBS 0.008197f
C214 B.n177 VSUBS 0.008197f
C215 B.n178 VSUBS 0.008197f
C216 B.n179 VSUBS 0.008197f
C217 B.n180 VSUBS 0.008197f
C218 B.n181 VSUBS 0.008197f
C219 B.n182 VSUBS 0.008197f
C220 B.n183 VSUBS 0.008197f
C221 B.n184 VSUBS 0.008197f
C222 B.n185 VSUBS 0.008197f
C223 B.n186 VSUBS 0.008197f
C224 B.n187 VSUBS 0.008197f
C225 B.n188 VSUBS 0.008197f
C226 B.n189 VSUBS 0.008197f
C227 B.n190 VSUBS 0.008197f
C228 B.n191 VSUBS 0.008197f
C229 B.n192 VSUBS 0.008197f
C230 B.n193 VSUBS 0.008197f
C231 B.n194 VSUBS 0.008197f
C232 B.n195 VSUBS 0.008197f
C233 B.n196 VSUBS 0.008197f
C234 B.n197 VSUBS 0.008197f
C235 B.n198 VSUBS 0.008197f
C236 B.n199 VSUBS 0.008197f
C237 B.n200 VSUBS 0.008197f
C238 B.n201 VSUBS 0.008197f
C239 B.n202 VSUBS 0.008197f
C240 B.n203 VSUBS 0.008197f
C241 B.n204 VSUBS 0.008197f
C242 B.n205 VSUBS 0.008197f
C243 B.n206 VSUBS 0.008197f
C244 B.n207 VSUBS 0.008197f
C245 B.n208 VSUBS 0.008197f
C246 B.n209 VSUBS 0.008197f
C247 B.n210 VSUBS 0.008197f
C248 B.n211 VSUBS 0.008197f
C249 B.n212 VSUBS 0.008197f
C250 B.n213 VSUBS 0.008197f
C251 B.n214 VSUBS 0.008197f
C252 B.n215 VSUBS 0.008197f
C253 B.n216 VSUBS 0.008197f
C254 B.n217 VSUBS 0.008197f
C255 B.n218 VSUBS 0.005666f
C256 B.n219 VSUBS 0.018992f
C257 B.n220 VSUBS 0.00663f
C258 B.n221 VSUBS 0.008197f
C259 B.n222 VSUBS 0.008197f
C260 B.n223 VSUBS 0.008197f
C261 B.n224 VSUBS 0.008197f
C262 B.n225 VSUBS 0.008197f
C263 B.n226 VSUBS 0.008197f
C264 B.n227 VSUBS 0.008197f
C265 B.n228 VSUBS 0.008197f
C266 B.n229 VSUBS 0.008197f
C267 B.n230 VSUBS 0.008197f
C268 B.n231 VSUBS 0.008197f
C269 B.t11 VSUBS 0.443151f
C270 B.t10 VSUBS 0.453024f
C271 B.t9 VSUBS 0.400671f
C272 B.n232 VSUBS 0.155546f
C273 B.n233 VSUBS 0.074889f
C274 B.n234 VSUBS 0.018992f
C275 B.n235 VSUBS 0.00663f
C276 B.n236 VSUBS 0.008197f
C277 B.n237 VSUBS 0.008197f
C278 B.n238 VSUBS 0.008197f
C279 B.n239 VSUBS 0.008197f
C280 B.n240 VSUBS 0.008197f
C281 B.n241 VSUBS 0.008197f
C282 B.n242 VSUBS 0.008197f
C283 B.n243 VSUBS 0.008197f
C284 B.n244 VSUBS 0.008197f
C285 B.n245 VSUBS 0.008197f
C286 B.n246 VSUBS 0.008197f
C287 B.n247 VSUBS 0.008197f
C288 B.n248 VSUBS 0.008197f
C289 B.n249 VSUBS 0.008197f
C290 B.n250 VSUBS 0.008197f
C291 B.n251 VSUBS 0.008197f
C292 B.n252 VSUBS 0.008197f
C293 B.n253 VSUBS 0.008197f
C294 B.n254 VSUBS 0.008197f
C295 B.n255 VSUBS 0.008197f
C296 B.n256 VSUBS 0.008197f
C297 B.n257 VSUBS 0.008197f
C298 B.n258 VSUBS 0.008197f
C299 B.n259 VSUBS 0.008197f
C300 B.n260 VSUBS 0.008197f
C301 B.n261 VSUBS 0.008197f
C302 B.n262 VSUBS 0.008197f
C303 B.n263 VSUBS 0.008197f
C304 B.n264 VSUBS 0.008197f
C305 B.n265 VSUBS 0.008197f
C306 B.n266 VSUBS 0.008197f
C307 B.n267 VSUBS 0.008197f
C308 B.n268 VSUBS 0.008197f
C309 B.n269 VSUBS 0.008197f
C310 B.n270 VSUBS 0.008197f
C311 B.n271 VSUBS 0.008197f
C312 B.n272 VSUBS 0.008197f
C313 B.n273 VSUBS 0.008197f
C314 B.n274 VSUBS 0.008197f
C315 B.n275 VSUBS 0.008197f
C316 B.n276 VSUBS 0.008197f
C317 B.n277 VSUBS 0.008197f
C318 B.n278 VSUBS 0.008197f
C319 B.n279 VSUBS 0.008197f
C320 B.n280 VSUBS 0.008197f
C321 B.n281 VSUBS 0.008197f
C322 B.n282 VSUBS 0.008197f
C323 B.n283 VSUBS 0.008197f
C324 B.n284 VSUBS 0.008197f
C325 B.n285 VSUBS 0.008197f
C326 B.n286 VSUBS 0.008197f
C327 B.n287 VSUBS 0.008197f
C328 B.n288 VSUBS 0.008197f
C329 B.n289 VSUBS 0.008197f
C330 B.n290 VSUBS 0.008197f
C331 B.n291 VSUBS 0.008197f
C332 B.n292 VSUBS 0.008197f
C333 B.n293 VSUBS 0.008197f
C334 B.n294 VSUBS 0.008197f
C335 B.n295 VSUBS 0.008197f
C336 B.n296 VSUBS 0.008197f
C337 B.n297 VSUBS 0.018161f
C338 B.n298 VSUBS 0.01728f
C339 B.n299 VSUBS 0.018375f
C340 B.n300 VSUBS 0.008197f
C341 B.n301 VSUBS 0.008197f
C342 B.n302 VSUBS 0.008197f
C343 B.n303 VSUBS 0.008197f
C344 B.n304 VSUBS 0.008197f
C345 B.n305 VSUBS 0.008197f
C346 B.n306 VSUBS 0.008197f
C347 B.n307 VSUBS 0.008197f
C348 B.n308 VSUBS 0.008197f
C349 B.n309 VSUBS 0.008197f
C350 B.n310 VSUBS 0.008197f
C351 B.n311 VSUBS 0.008197f
C352 B.n312 VSUBS 0.008197f
C353 B.n313 VSUBS 0.008197f
C354 B.n314 VSUBS 0.008197f
C355 B.n315 VSUBS 0.008197f
C356 B.n316 VSUBS 0.008197f
C357 B.n317 VSUBS 0.008197f
C358 B.n318 VSUBS 0.008197f
C359 B.n319 VSUBS 0.008197f
C360 B.n320 VSUBS 0.008197f
C361 B.n321 VSUBS 0.008197f
C362 B.n322 VSUBS 0.008197f
C363 B.n323 VSUBS 0.008197f
C364 B.n324 VSUBS 0.008197f
C365 B.n325 VSUBS 0.008197f
C366 B.n326 VSUBS 0.008197f
C367 B.n327 VSUBS 0.008197f
C368 B.n328 VSUBS 0.008197f
C369 B.n329 VSUBS 0.008197f
C370 B.n330 VSUBS 0.008197f
C371 B.n331 VSUBS 0.008197f
C372 B.n332 VSUBS 0.008197f
C373 B.n333 VSUBS 0.008197f
C374 B.n334 VSUBS 0.008197f
C375 B.n335 VSUBS 0.008197f
C376 B.n336 VSUBS 0.008197f
C377 B.n337 VSUBS 0.008197f
C378 B.n338 VSUBS 0.008197f
C379 B.n339 VSUBS 0.008197f
C380 B.n340 VSUBS 0.008197f
C381 B.n341 VSUBS 0.008197f
C382 B.n342 VSUBS 0.008197f
C383 B.n343 VSUBS 0.008197f
C384 B.n344 VSUBS 0.008197f
C385 B.n345 VSUBS 0.008197f
C386 B.n346 VSUBS 0.008197f
C387 B.n347 VSUBS 0.008197f
C388 B.n348 VSUBS 0.008197f
C389 B.n349 VSUBS 0.008197f
C390 B.n350 VSUBS 0.008197f
C391 B.n351 VSUBS 0.01728f
C392 B.n352 VSUBS 0.018161f
C393 B.n353 VSUBS 0.018161f
C394 B.n354 VSUBS 0.008197f
C395 B.n355 VSUBS 0.008197f
C396 B.n356 VSUBS 0.008197f
C397 B.n357 VSUBS 0.008197f
C398 B.n358 VSUBS 0.008197f
C399 B.n359 VSUBS 0.008197f
C400 B.n360 VSUBS 0.008197f
C401 B.n361 VSUBS 0.008197f
C402 B.n362 VSUBS 0.008197f
C403 B.n363 VSUBS 0.008197f
C404 B.n364 VSUBS 0.008197f
C405 B.n365 VSUBS 0.008197f
C406 B.n366 VSUBS 0.008197f
C407 B.n367 VSUBS 0.008197f
C408 B.n368 VSUBS 0.008197f
C409 B.n369 VSUBS 0.008197f
C410 B.n370 VSUBS 0.008197f
C411 B.n371 VSUBS 0.008197f
C412 B.n372 VSUBS 0.008197f
C413 B.n373 VSUBS 0.008197f
C414 B.n374 VSUBS 0.008197f
C415 B.n375 VSUBS 0.008197f
C416 B.n376 VSUBS 0.008197f
C417 B.n377 VSUBS 0.008197f
C418 B.n378 VSUBS 0.008197f
C419 B.n379 VSUBS 0.008197f
C420 B.n380 VSUBS 0.008197f
C421 B.n381 VSUBS 0.008197f
C422 B.n382 VSUBS 0.008197f
C423 B.n383 VSUBS 0.008197f
C424 B.n384 VSUBS 0.008197f
C425 B.n385 VSUBS 0.008197f
C426 B.n386 VSUBS 0.008197f
C427 B.n387 VSUBS 0.008197f
C428 B.n388 VSUBS 0.008197f
C429 B.n389 VSUBS 0.008197f
C430 B.n390 VSUBS 0.008197f
C431 B.n391 VSUBS 0.008197f
C432 B.n392 VSUBS 0.008197f
C433 B.n393 VSUBS 0.008197f
C434 B.n394 VSUBS 0.008197f
C435 B.n395 VSUBS 0.008197f
C436 B.n396 VSUBS 0.008197f
C437 B.n397 VSUBS 0.008197f
C438 B.n398 VSUBS 0.008197f
C439 B.n399 VSUBS 0.008197f
C440 B.n400 VSUBS 0.008197f
C441 B.n401 VSUBS 0.008197f
C442 B.n402 VSUBS 0.008197f
C443 B.n403 VSUBS 0.008197f
C444 B.n404 VSUBS 0.008197f
C445 B.n405 VSUBS 0.008197f
C446 B.n406 VSUBS 0.008197f
C447 B.n407 VSUBS 0.008197f
C448 B.n408 VSUBS 0.008197f
C449 B.n409 VSUBS 0.008197f
C450 B.n410 VSUBS 0.008197f
C451 B.n411 VSUBS 0.008197f
C452 B.n412 VSUBS 0.008197f
C453 B.n413 VSUBS 0.005666f
C454 B.n414 VSUBS 0.018992f
C455 B.n415 VSUBS 0.00663f
C456 B.n416 VSUBS 0.008197f
C457 B.n417 VSUBS 0.008197f
C458 B.n418 VSUBS 0.008197f
C459 B.n419 VSUBS 0.008197f
C460 B.n420 VSUBS 0.008197f
C461 B.n421 VSUBS 0.008197f
C462 B.n422 VSUBS 0.008197f
C463 B.n423 VSUBS 0.008197f
C464 B.n424 VSUBS 0.008197f
C465 B.n425 VSUBS 0.008197f
C466 B.n426 VSUBS 0.008197f
C467 B.n427 VSUBS 0.00663f
C468 B.n428 VSUBS 0.018992f
C469 B.n429 VSUBS 0.005666f
C470 B.n430 VSUBS 0.008197f
C471 B.n431 VSUBS 0.008197f
C472 B.n432 VSUBS 0.008197f
C473 B.n433 VSUBS 0.008197f
C474 B.n434 VSUBS 0.008197f
C475 B.n435 VSUBS 0.008197f
C476 B.n436 VSUBS 0.008197f
C477 B.n437 VSUBS 0.008197f
C478 B.n438 VSUBS 0.008197f
C479 B.n439 VSUBS 0.008197f
C480 B.n440 VSUBS 0.008197f
C481 B.n441 VSUBS 0.008197f
C482 B.n442 VSUBS 0.008197f
C483 B.n443 VSUBS 0.008197f
C484 B.n444 VSUBS 0.008197f
C485 B.n445 VSUBS 0.008197f
C486 B.n446 VSUBS 0.008197f
C487 B.n447 VSUBS 0.008197f
C488 B.n448 VSUBS 0.008197f
C489 B.n449 VSUBS 0.008197f
C490 B.n450 VSUBS 0.008197f
C491 B.n451 VSUBS 0.008197f
C492 B.n452 VSUBS 0.008197f
C493 B.n453 VSUBS 0.008197f
C494 B.n454 VSUBS 0.008197f
C495 B.n455 VSUBS 0.008197f
C496 B.n456 VSUBS 0.008197f
C497 B.n457 VSUBS 0.008197f
C498 B.n458 VSUBS 0.008197f
C499 B.n459 VSUBS 0.008197f
C500 B.n460 VSUBS 0.008197f
C501 B.n461 VSUBS 0.008197f
C502 B.n462 VSUBS 0.008197f
C503 B.n463 VSUBS 0.008197f
C504 B.n464 VSUBS 0.008197f
C505 B.n465 VSUBS 0.008197f
C506 B.n466 VSUBS 0.008197f
C507 B.n467 VSUBS 0.008197f
C508 B.n468 VSUBS 0.008197f
C509 B.n469 VSUBS 0.008197f
C510 B.n470 VSUBS 0.008197f
C511 B.n471 VSUBS 0.008197f
C512 B.n472 VSUBS 0.008197f
C513 B.n473 VSUBS 0.008197f
C514 B.n474 VSUBS 0.008197f
C515 B.n475 VSUBS 0.008197f
C516 B.n476 VSUBS 0.008197f
C517 B.n477 VSUBS 0.008197f
C518 B.n478 VSUBS 0.008197f
C519 B.n479 VSUBS 0.008197f
C520 B.n480 VSUBS 0.008197f
C521 B.n481 VSUBS 0.008197f
C522 B.n482 VSUBS 0.008197f
C523 B.n483 VSUBS 0.008197f
C524 B.n484 VSUBS 0.008197f
C525 B.n485 VSUBS 0.008197f
C526 B.n486 VSUBS 0.008197f
C527 B.n487 VSUBS 0.008197f
C528 B.n488 VSUBS 0.008197f
C529 B.n489 VSUBS 0.018161f
C530 B.n490 VSUBS 0.018161f
C531 B.n491 VSUBS 0.01728f
C532 B.n492 VSUBS 0.008197f
C533 B.n493 VSUBS 0.008197f
C534 B.n494 VSUBS 0.008197f
C535 B.n495 VSUBS 0.008197f
C536 B.n496 VSUBS 0.008197f
C537 B.n497 VSUBS 0.008197f
C538 B.n498 VSUBS 0.008197f
C539 B.n499 VSUBS 0.008197f
C540 B.n500 VSUBS 0.008197f
C541 B.n501 VSUBS 0.008197f
C542 B.n502 VSUBS 0.008197f
C543 B.n503 VSUBS 0.008197f
C544 B.n504 VSUBS 0.008197f
C545 B.n505 VSUBS 0.008197f
C546 B.n506 VSUBS 0.008197f
C547 B.n507 VSUBS 0.008197f
C548 B.n508 VSUBS 0.008197f
C549 B.n509 VSUBS 0.008197f
C550 B.n510 VSUBS 0.008197f
C551 B.n511 VSUBS 0.008197f
C552 B.n512 VSUBS 0.008197f
C553 B.n513 VSUBS 0.008197f
C554 B.n514 VSUBS 0.008197f
C555 B.n515 VSUBS 0.010697f
C556 B.n516 VSUBS 0.011395f
C557 B.n517 VSUBS 0.02266f
C558 VDD2.t1 VSUBS 0.258142f
C559 VDD2.t0 VSUBS 0.258142f
C560 VDD2.n0 VSUBS 2.63148f
C561 VDD2.t3 VSUBS 0.258142f
C562 VDD2.t2 VSUBS 0.258142f
C563 VDD2.n1 VSUBS 1.99505f
C564 VDD2.n2 VSUBS 3.95387f
C565 VN.t2 VSUBS 1.44872f
C566 VN.t3 VSUBS 1.44866f
C567 VN.n0 VSUBS 1.09458f
C568 VN.t1 VSUBS 1.44872f
C569 VN.t0 VSUBS 1.44866f
C570 VN.n1 VSUBS 2.27406f
C571 VDD1.t2 VSUBS 0.258048f
C572 VDD1.t3 VSUBS 0.258048f
C573 VDD1.n0 VSUBS 1.99483f
C574 VDD1.t0 VSUBS 0.258048f
C575 VDD1.t1 VSUBS 0.258048f
C576 VDD1.n1 VSUBS 2.65585f
C577 VTAIL.t3 VSUBS 2.00806f
C578 VTAIL.n0 VSUBS 0.702387f
C579 VTAIL.t6 VSUBS 2.00806f
C580 VTAIL.n1 VSUBS 0.731497f
C581 VTAIL.t7 VSUBS 2.00806f
C582 VTAIL.n2 VSUBS 1.82737f
C583 VTAIL.t1 VSUBS 2.00807f
C584 VTAIL.n3 VSUBS 1.82737f
C585 VTAIL.t0 VSUBS 2.00807f
C586 VTAIL.n4 VSUBS 0.73149f
C587 VTAIL.t4 VSUBS 2.00807f
C588 VTAIL.n5 VSUBS 0.73149f
C589 VTAIL.t5 VSUBS 2.00806f
C590 VTAIL.n6 VSUBS 1.82737f
C591 VTAIL.t2 VSUBS 2.00806f
C592 VTAIL.n7 VSUBS 1.78958f
C593 VP.n0 VSUBS 0.062096f
C594 VP.t0 VSUBS 1.49181f
C595 VP.t1 VSUBS 1.49188f
C596 VP.n1 VSUBS 2.31645f
C597 VP.n2 VSUBS 3.75583f
C598 VP.t3 VSUBS 1.46578f
C599 VP.n3 VSUBS 0.582306f
C600 VP.n4 VSUBS 0.014091f
C601 VP.t2 VSUBS 1.46578f
C602 VP.n5 VSUBS 0.582306f
C603 VP.n6 VSUBS 0.048122f
.ends

