* NGSPICE file created from diff_pair_sample_1199.ext - technology: sky130A

.subckt diff_pair_sample_1199 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t9 VN.t0 VTAIL.t6 B.t9 sky130_fd_pr__nfet_01v8 ad=0.4875 pd=3.28 as=0.20625 ps=1.58 w=1.25 l=2.38
X1 VDD1.t9 VP.t0 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.20625 pd=1.58 as=0.4875 ps=3.28 w=1.25 l=2.38
X2 VDD1.t8 VP.t1 VTAIL.t14 B.t8 sky130_fd_pr__nfet_01v8 ad=0.4875 pd=3.28 as=0.20625 ps=1.58 w=1.25 l=2.38
X3 VTAIL.t7 VN.t1 VDD2.t8 B.t1 sky130_fd_pr__nfet_01v8 ad=0.20625 pd=1.58 as=0.20625 ps=1.58 w=1.25 l=2.38
X4 VTAIL.t2 VP.t2 VDD1.t7 B.t2 sky130_fd_pr__nfet_01v8 ad=0.20625 pd=1.58 as=0.20625 ps=1.58 w=1.25 l=2.38
X5 VDD2.t7 VN.t2 VTAIL.t8 B.t8 sky130_fd_pr__nfet_01v8 ad=0.4875 pd=3.28 as=0.20625 ps=1.58 w=1.25 l=2.38
X6 VDD2.t6 VN.t3 VTAIL.t12 B.t7 sky130_fd_pr__nfet_01v8 ad=0.20625 pd=1.58 as=0.20625 ps=1.58 w=1.25 l=2.38
X7 B.t23 B.t21 B.t22 B.t15 sky130_fd_pr__nfet_01v8 ad=0.4875 pd=3.28 as=0 ps=0 w=1.25 l=2.38
X8 B.t20 B.t18 B.t19 B.t11 sky130_fd_pr__nfet_01v8 ad=0.4875 pd=3.28 as=0 ps=0 w=1.25 l=2.38
X9 VTAIL.t9 VN.t4 VDD2.t5 B.t6 sky130_fd_pr__nfet_01v8 ad=0.20625 pd=1.58 as=0.20625 ps=1.58 w=1.25 l=2.38
X10 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=0.4875 pd=3.28 as=0 ps=0 w=1.25 l=2.38
X11 VTAIL.t13 VN.t5 VDD2.t4 B.t5 sky130_fd_pr__nfet_01v8 ad=0.20625 pd=1.58 as=0.20625 ps=1.58 w=1.25 l=2.38
X12 VTAIL.t1 VP.t3 VDD1.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=0.20625 pd=1.58 as=0.20625 ps=1.58 w=1.25 l=2.38
X13 VDD2.t3 VN.t6 VTAIL.t10 B.t4 sky130_fd_pr__nfet_01v8 ad=0.20625 pd=1.58 as=0.4875 ps=3.28 w=1.25 l=2.38
X14 VDD2.t2 VN.t7 VTAIL.t4 B.t0 sky130_fd_pr__nfet_01v8 ad=0.20625 pd=1.58 as=0.20625 ps=1.58 w=1.25 l=2.38
X15 VDD1.t5 VP.t4 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.20625 pd=1.58 as=0.20625 ps=1.58 w=1.25 l=2.38
X16 VDD1.t4 VP.t5 VTAIL.t17 B.t7 sky130_fd_pr__nfet_01v8 ad=0.20625 pd=1.58 as=0.20625 ps=1.58 w=1.25 l=2.38
X17 VTAIL.t5 VN.t8 VDD2.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=0.20625 pd=1.58 as=0.20625 ps=1.58 w=1.25 l=2.38
X18 VTAIL.t19 VP.t6 VDD1.t3 B.t5 sky130_fd_pr__nfet_01v8 ad=0.20625 pd=1.58 as=0.20625 ps=1.58 w=1.25 l=2.38
X19 VDD1.t2 VP.t7 VTAIL.t18 B.t4 sky130_fd_pr__nfet_01v8 ad=0.20625 pd=1.58 as=0.4875 ps=3.28 w=1.25 l=2.38
X20 VDD2.t0 VN.t9 VTAIL.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=0.20625 pd=1.58 as=0.4875 ps=3.28 w=1.25 l=2.38
X21 VTAIL.t16 VP.t8 VDD1.t1 B.t6 sky130_fd_pr__nfet_01v8 ad=0.20625 pd=1.58 as=0.20625 ps=1.58 w=1.25 l=2.38
X22 VDD1.t0 VP.t9 VTAIL.t15 B.t9 sky130_fd_pr__nfet_01v8 ad=0.4875 pd=3.28 as=0.20625 ps=1.58 w=1.25 l=2.38
X23 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=0.4875 pd=3.28 as=0 ps=0 w=1.25 l=2.38
R0 VN.n73 VN.n38 161.3
R1 VN.n72 VN.n71 161.3
R2 VN.n70 VN.n39 161.3
R3 VN.n69 VN.n68 161.3
R4 VN.n67 VN.n40 161.3
R5 VN.n66 VN.n65 161.3
R6 VN.n64 VN.n63 161.3
R7 VN.n62 VN.n42 161.3
R8 VN.n61 VN.n60 161.3
R9 VN.n59 VN.n43 161.3
R10 VN.n58 VN.n57 161.3
R11 VN.n55 VN.n44 161.3
R12 VN.n54 VN.n53 161.3
R13 VN.n52 VN.n45 161.3
R14 VN.n51 VN.n50 161.3
R15 VN.n49 VN.n46 161.3
R16 VN.n35 VN.n0 161.3
R17 VN.n34 VN.n33 161.3
R18 VN.n32 VN.n1 161.3
R19 VN.n31 VN.n30 161.3
R20 VN.n29 VN.n2 161.3
R21 VN.n28 VN.n27 161.3
R22 VN.n26 VN.n25 161.3
R23 VN.n24 VN.n4 161.3
R24 VN.n23 VN.n22 161.3
R25 VN.n21 VN.n5 161.3
R26 VN.n20 VN.n19 161.3
R27 VN.n17 VN.n6 161.3
R28 VN.n16 VN.n15 161.3
R29 VN.n14 VN.n7 161.3
R30 VN.n13 VN.n12 161.3
R31 VN.n11 VN.n8 161.3
R32 VN.n37 VN.n36 102.438
R33 VN.n75 VN.n74 102.438
R34 VN.n30 VN.n1 56.5193
R35 VN.n68 VN.n39 56.5193
R36 VN.n12 VN.n7 50.6917
R37 VN.n24 VN.n23 50.6917
R38 VN.n50 VN.n45 50.6917
R39 VN.n62 VN.n61 50.6917
R40 VN.n10 VN.n9 49.8376
R41 VN.n48 VN.n47 49.8376
R42 VN.n9 VN.t0 45.7749
R43 VN.n47 VN.t6 45.7749
R44 VN VN.n75 43.9944
R45 VN.n16 VN.n7 30.2951
R46 VN.n23 VN.n5 30.2951
R47 VN.n54 VN.n45 30.2951
R48 VN.n61 VN.n43 30.2951
R49 VN.n12 VN.n11 24.4675
R50 VN.n17 VN.n16 24.4675
R51 VN.n19 VN.n5 24.4675
R52 VN.n25 VN.n24 24.4675
R53 VN.n29 VN.n28 24.4675
R54 VN.n30 VN.n29 24.4675
R55 VN.n34 VN.n1 24.4675
R56 VN.n35 VN.n34 24.4675
R57 VN.n50 VN.n49 24.4675
R58 VN.n57 VN.n43 24.4675
R59 VN.n55 VN.n54 24.4675
R60 VN.n68 VN.n67 24.4675
R61 VN.n67 VN.n66 24.4675
R62 VN.n63 VN.n62 24.4675
R63 VN.n73 VN.n72 24.4675
R64 VN.n72 VN.n39 24.4675
R65 VN.n11 VN.n10 22.5101
R66 VN.n25 VN.n3 22.5101
R67 VN.n49 VN.n48 22.5101
R68 VN.n63 VN.n41 22.5101
R69 VN.n10 VN.t1 12.6581
R70 VN.n18 VN.t3 12.6581
R71 VN.n3 VN.t8 12.6581
R72 VN.n36 VN.t9 12.6581
R73 VN.n48 VN.t4 12.6581
R74 VN.n56 VN.t7 12.6581
R75 VN.n41 VN.t5 12.6581
R76 VN.n74 VN.t2 12.6581
R77 VN.n18 VN.n17 12.234
R78 VN.n19 VN.n18 12.234
R79 VN.n57 VN.n56 12.234
R80 VN.n56 VN.n55 12.234
R81 VN.n36 VN.n35 8.31928
R82 VN.n74 VN.n73 8.31928
R83 VN.n47 VN.n46 6.95571
R84 VN.n9 VN.n8 6.95571
R85 VN.n28 VN.n3 1.95786
R86 VN.n66 VN.n41 1.95786
R87 VN.n75 VN.n38 0.278367
R88 VN.n37 VN.n0 0.278367
R89 VN.n71 VN.n38 0.189894
R90 VN.n71 VN.n70 0.189894
R91 VN.n70 VN.n69 0.189894
R92 VN.n69 VN.n40 0.189894
R93 VN.n65 VN.n40 0.189894
R94 VN.n65 VN.n64 0.189894
R95 VN.n64 VN.n42 0.189894
R96 VN.n60 VN.n42 0.189894
R97 VN.n60 VN.n59 0.189894
R98 VN.n59 VN.n58 0.189894
R99 VN.n58 VN.n44 0.189894
R100 VN.n53 VN.n44 0.189894
R101 VN.n53 VN.n52 0.189894
R102 VN.n52 VN.n51 0.189894
R103 VN.n51 VN.n46 0.189894
R104 VN.n13 VN.n8 0.189894
R105 VN.n14 VN.n13 0.189894
R106 VN.n15 VN.n14 0.189894
R107 VN.n15 VN.n6 0.189894
R108 VN.n20 VN.n6 0.189894
R109 VN.n21 VN.n20 0.189894
R110 VN.n22 VN.n21 0.189894
R111 VN.n22 VN.n4 0.189894
R112 VN.n26 VN.n4 0.189894
R113 VN.n27 VN.n26 0.189894
R114 VN.n27 VN.n2 0.189894
R115 VN.n31 VN.n2 0.189894
R116 VN.n32 VN.n31 0.189894
R117 VN.n33 VN.n32 0.189894
R118 VN.n33 VN.n0 0.189894
R119 VN VN.n37 0.153454
R120 VTAIL.n17 VTAIL.t11 155.327
R121 VTAIL.n2 VTAIL.t18 155.327
R122 VTAIL.n16 VTAIL.t3 155.327
R123 VTAIL.n11 VTAIL.t10 155.327
R124 VTAIL.n19 VTAIL.n18 129.168
R125 VTAIL.n1 VTAIL.n0 129.168
R126 VTAIL.n4 VTAIL.n3 129.168
R127 VTAIL.n6 VTAIL.n5 129.168
R128 VTAIL.n15 VTAIL.n14 129.167
R129 VTAIL.n13 VTAIL.n12 129.167
R130 VTAIL.n10 VTAIL.n9 129.167
R131 VTAIL.n8 VTAIL.n7 129.167
R132 VTAIL.n8 VTAIL.n6 18.1169
R133 VTAIL.n18 VTAIL.t12 15.8405
R134 VTAIL.n18 VTAIL.t5 15.8405
R135 VTAIL.n0 VTAIL.t6 15.8405
R136 VTAIL.n0 VTAIL.t7 15.8405
R137 VTAIL.n3 VTAIL.t0 15.8405
R138 VTAIL.n3 VTAIL.t16 15.8405
R139 VTAIL.n5 VTAIL.t14 15.8405
R140 VTAIL.n5 VTAIL.t19 15.8405
R141 VTAIL.n14 VTAIL.t17 15.8405
R142 VTAIL.n14 VTAIL.t2 15.8405
R143 VTAIL.n12 VTAIL.t15 15.8405
R144 VTAIL.n12 VTAIL.t1 15.8405
R145 VTAIL.n9 VTAIL.t4 15.8405
R146 VTAIL.n9 VTAIL.t9 15.8405
R147 VTAIL.n7 VTAIL.t8 15.8405
R148 VTAIL.n7 VTAIL.t13 15.8405
R149 VTAIL.n17 VTAIL.n16 15.7807
R150 VTAIL.n10 VTAIL.n8 2.33671
R151 VTAIL.n11 VTAIL.n10 2.33671
R152 VTAIL.n15 VTAIL.n13 2.33671
R153 VTAIL.n16 VTAIL.n15 2.33671
R154 VTAIL.n6 VTAIL.n4 2.33671
R155 VTAIL.n4 VTAIL.n2 2.33671
R156 VTAIL.n19 VTAIL.n17 2.33671
R157 VTAIL VTAIL.n1 1.81084
R158 VTAIL.n13 VTAIL.n11 1.63843
R159 VTAIL.n2 VTAIL.n1 1.63843
R160 VTAIL VTAIL.n19 0.526362
R161 VDD2.n1 VDD2.t9 174.341
R162 VDD2.n4 VDD2.t7 172.006
R163 VDD2.n3 VDD2.n2 147.544
R164 VDD2 VDD2.n7 147.542
R165 VDD2.n1 VDD2.n0 145.847
R166 VDD2.n6 VDD2.n5 145.846
R167 VDD2.n4 VDD2.n3 35.8899
R168 VDD2.n7 VDD2.t5 15.8405
R169 VDD2.n7 VDD2.t3 15.8405
R170 VDD2.n5 VDD2.t4 15.8405
R171 VDD2.n5 VDD2.t2 15.8405
R172 VDD2.n2 VDD2.t1 15.8405
R173 VDD2.n2 VDD2.t0 15.8405
R174 VDD2.n0 VDD2.t8 15.8405
R175 VDD2.n0 VDD2.t6 15.8405
R176 VDD2.n6 VDD2.n4 2.33671
R177 VDD2 VDD2.n6 0.642741
R178 VDD2.n3 VDD2.n1 0.529206
R179 B.n610 B.n609 585
R180 B.n179 B.n118 585
R181 B.n178 B.n177 585
R182 B.n176 B.n175 585
R183 B.n174 B.n173 585
R184 B.n172 B.n171 585
R185 B.n170 B.n169 585
R186 B.n168 B.n167 585
R187 B.n166 B.n165 585
R188 B.n164 B.n163 585
R189 B.n162 B.n161 585
R190 B.n160 B.n159 585
R191 B.n158 B.n157 585
R192 B.n156 B.n155 585
R193 B.n154 B.n153 585
R194 B.n152 B.n151 585
R195 B.n150 B.n149 585
R196 B.n148 B.n147 585
R197 B.n146 B.n145 585
R198 B.n144 B.n143 585
R199 B.n142 B.n141 585
R200 B.n140 B.n139 585
R201 B.n138 B.n137 585
R202 B.n136 B.n135 585
R203 B.n134 B.n133 585
R204 B.n132 B.n131 585
R205 B.n130 B.n129 585
R206 B.n128 B.n127 585
R207 B.n126 B.n125 585
R208 B.n102 B.n101 585
R209 B.n608 B.n103 585
R210 B.n613 B.n103 585
R211 B.n607 B.n606 585
R212 B.n606 B.n99 585
R213 B.n605 B.n98 585
R214 B.n619 B.n98 585
R215 B.n604 B.n97 585
R216 B.n620 B.n97 585
R217 B.n603 B.n96 585
R218 B.n621 B.n96 585
R219 B.n602 B.n601 585
R220 B.n601 B.n92 585
R221 B.n600 B.n91 585
R222 B.n627 B.n91 585
R223 B.n599 B.n90 585
R224 B.n628 B.n90 585
R225 B.n598 B.n89 585
R226 B.n629 B.n89 585
R227 B.n597 B.n596 585
R228 B.n596 B.n85 585
R229 B.n595 B.n84 585
R230 B.n635 B.n84 585
R231 B.n594 B.n83 585
R232 B.n636 B.n83 585
R233 B.n593 B.n82 585
R234 B.n637 B.n82 585
R235 B.n592 B.n591 585
R236 B.n591 B.n78 585
R237 B.n590 B.n77 585
R238 B.n643 B.n77 585
R239 B.n589 B.n76 585
R240 B.n644 B.n76 585
R241 B.n588 B.n75 585
R242 B.n645 B.n75 585
R243 B.n587 B.n586 585
R244 B.n586 B.n71 585
R245 B.n585 B.n70 585
R246 B.n651 B.n70 585
R247 B.n584 B.n69 585
R248 B.n652 B.n69 585
R249 B.n583 B.n68 585
R250 B.n653 B.n68 585
R251 B.n582 B.n581 585
R252 B.n581 B.n64 585
R253 B.n580 B.n63 585
R254 B.n659 B.n63 585
R255 B.n579 B.n62 585
R256 B.n660 B.n62 585
R257 B.n578 B.n61 585
R258 B.n661 B.n61 585
R259 B.n577 B.n576 585
R260 B.n576 B.n57 585
R261 B.n575 B.n56 585
R262 B.n667 B.n56 585
R263 B.n574 B.n55 585
R264 B.n668 B.n55 585
R265 B.n573 B.n54 585
R266 B.n669 B.n54 585
R267 B.n572 B.n571 585
R268 B.n571 B.n50 585
R269 B.n570 B.n49 585
R270 B.n675 B.n49 585
R271 B.n569 B.n48 585
R272 B.n676 B.n48 585
R273 B.n568 B.n47 585
R274 B.n677 B.n47 585
R275 B.n567 B.n566 585
R276 B.n566 B.n43 585
R277 B.n565 B.n42 585
R278 B.n683 B.n42 585
R279 B.n564 B.n41 585
R280 B.n684 B.n41 585
R281 B.n563 B.n40 585
R282 B.n685 B.n40 585
R283 B.n562 B.n561 585
R284 B.n561 B.n36 585
R285 B.n560 B.n35 585
R286 B.n691 B.n35 585
R287 B.n559 B.n34 585
R288 B.n692 B.n34 585
R289 B.n558 B.n33 585
R290 B.n693 B.n33 585
R291 B.n557 B.n556 585
R292 B.n556 B.n29 585
R293 B.n555 B.n28 585
R294 B.n699 B.n28 585
R295 B.n554 B.n27 585
R296 B.n700 B.n27 585
R297 B.n553 B.n26 585
R298 B.n701 B.n26 585
R299 B.n552 B.n551 585
R300 B.n551 B.n22 585
R301 B.n550 B.n21 585
R302 B.n707 B.n21 585
R303 B.n549 B.n20 585
R304 B.n708 B.n20 585
R305 B.n548 B.n19 585
R306 B.n709 B.n19 585
R307 B.n547 B.n546 585
R308 B.n546 B.n15 585
R309 B.n545 B.n14 585
R310 B.n715 B.n14 585
R311 B.n544 B.n13 585
R312 B.n716 B.n13 585
R313 B.n543 B.n12 585
R314 B.n717 B.n12 585
R315 B.n542 B.n541 585
R316 B.n541 B.n8 585
R317 B.n540 B.n7 585
R318 B.n723 B.n7 585
R319 B.n539 B.n6 585
R320 B.n724 B.n6 585
R321 B.n538 B.n5 585
R322 B.n725 B.n5 585
R323 B.n537 B.n536 585
R324 B.n536 B.n4 585
R325 B.n535 B.n180 585
R326 B.n535 B.n534 585
R327 B.n525 B.n181 585
R328 B.n182 B.n181 585
R329 B.n527 B.n526 585
R330 B.n528 B.n527 585
R331 B.n524 B.n187 585
R332 B.n187 B.n186 585
R333 B.n523 B.n522 585
R334 B.n522 B.n521 585
R335 B.n189 B.n188 585
R336 B.n190 B.n189 585
R337 B.n514 B.n513 585
R338 B.n515 B.n514 585
R339 B.n512 B.n195 585
R340 B.n195 B.n194 585
R341 B.n511 B.n510 585
R342 B.n510 B.n509 585
R343 B.n197 B.n196 585
R344 B.n198 B.n197 585
R345 B.n502 B.n501 585
R346 B.n503 B.n502 585
R347 B.n500 B.n203 585
R348 B.n203 B.n202 585
R349 B.n499 B.n498 585
R350 B.n498 B.n497 585
R351 B.n205 B.n204 585
R352 B.n206 B.n205 585
R353 B.n490 B.n489 585
R354 B.n491 B.n490 585
R355 B.n488 B.n211 585
R356 B.n211 B.n210 585
R357 B.n487 B.n486 585
R358 B.n486 B.n485 585
R359 B.n213 B.n212 585
R360 B.n214 B.n213 585
R361 B.n478 B.n477 585
R362 B.n479 B.n478 585
R363 B.n476 B.n219 585
R364 B.n219 B.n218 585
R365 B.n475 B.n474 585
R366 B.n474 B.n473 585
R367 B.n221 B.n220 585
R368 B.n222 B.n221 585
R369 B.n466 B.n465 585
R370 B.n467 B.n466 585
R371 B.n464 B.n227 585
R372 B.n227 B.n226 585
R373 B.n463 B.n462 585
R374 B.n462 B.n461 585
R375 B.n229 B.n228 585
R376 B.n230 B.n229 585
R377 B.n454 B.n453 585
R378 B.n455 B.n454 585
R379 B.n452 B.n235 585
R380 B.n235 B.n234 585
R381 B.n451 B.n450 585
R382 B.n450 B.n449 585
R383 B.n237 B.n236 585
R384 B.n238 B.n237 585
R385 B.n442 B.n441 585
R386 B.n443 B.n442 585
R387 B.n440 B.n243 585
R388 B.n243 B.n242 585
R389 B.n439 B.n438 585
R390 B.n438 B.n437 585
R391 B.n245 B.n244 585
R392 B.n246 B.n245 585
R393 B.n430 B.n429 585
R394 B.n431 B.n430 585
R395 B.n428 B.n251 585
R396 B.n251 B.n250 585
R397 B.n427 B.n426 585
R398 B.n426 B.n425 585
R399 B.n253 B.n252 585
R400 B.n254 B.n253 585
R401 B.n418 B.n417 585
R402 B.n419 B.n418 585
R403 B.n416 B.n259 585
R404 B.n259 B.n258 585
R405 B.n415 B.n414 585
R406 B.n414 B.n413 585
R407 B.n261 B.n260 585
R408 B.n262 B.n261 585
R409 B.n406 B.n405 585
R410 B.n407 B.n406 585
R411 B.n404 B.n267 585
R412 B.n267 B.n266 585
R413 B.n403 B.n402 585
R414 B.n402 B.n401 585
R415 B.n269 B.n268 585
R416 B.n270 B.n269 585
R417 B.n394 B.n393 585
R418 B.n395 B.n394 585
R419 B.n392 B.n274 585
R420 B.n278 B.n274 585
R421 B.n391 B.n390 585
R422 B.n390 B.n389 585
R423 B.n276 B.n275 585
R424 B.n277 B.n276 585
R425 B.n382 B.n381 585
R426 B.n383 B.n382 585
R427 B.n380 B.n283 585
R428 B.n283 B.n282 585
R429 B.n379 B.n378 585
R430 B.n378 B.n377 585
R431 B.n285 B.n284 585
R432 B.n286 B.n285 585
R433 B.n370 B.n369 585
R434 B.n371 B.n370 585
R435 B.n289 B.n288 585
R436 B.n310 B.n308 585
R437 B.n311 B.n307 585
R438 B.n311 B.n290 585
R439 B.n314 B.n313 585
R440 B.n315 B.n306 585
R441 B.n317 B.n316 585
R442 B.n319 B.n305 585
R443 B.n322 B.n321 585
R444 B.n323 B.n304 585
R445 B.n328 B.n327 585
R446 B.n330 B.n303 585
R447 B.n333 B.n332 585
R448 B.n334 B.n302 585
R449 B.n336 B.n335 585
R450 B.n338 B.n301 585
R451 B.n341 B.n340 585
R452 B.n342 B.n300 585
R453 B.n344 B.n343 585
R454 B.n346 B.n299 585
R455 B.n349 B.n348 585
R456 B.n351 B.n296 585
R457 B.n353 B.n352 585
R458 B.n355 B.n295 585
R459 B.n358 B.n357 585
R460 B.n359 B.n294 585
R461 B.n361 B.n360 585
R462 B.n363 B.n293 585
R463 B.n364 B.n292 585
R464 B.n367 B.n366 585
R465 B.n368 B.n291 585
R466 B.n291 B.n290 585
R467 B.n373 B.n372 585
R468 B.n372 B.n371 585
R469 B.n374 B.n287 585
R470 B.n287 B.n286 585
R471 B.n376 B.n375 585
R472 B.n377 B.n376 585
R473 B.n281 B.n280 585
R474 B.n282 B.n281 585
R475 B.n385 B.n384 585
R476 B.n384 B.n383 585
R477 B.n386 B.n279 585
R478 B.n279 B.n277 585
R479 B.n388 B.n387 585
R480 B.n389 B.n388 585
R481 B.n273 B.n272 585
R482 B.n278 B.n273 585
R483 B.n397 B.n396 585
R484 B.n396 B.n395 585
R485 B.n398 B.n271 585
R486 B.n271 B.n270 585
R487 B.n400 B.n399 585
R488 B.n401 B.n400 585
R489 B.n265 B.n264 585
R490 B.n266 B.n265 585
R491 B.n409 B.n408 585
R492 B.n408 B.n407 585
R493 B.n410 B.n263 585
R494 B.n263 B.n262 585
R495 B.n412 B.n411 585
R496 B.n413 B.n412 585
R497 B.n257 B.n256 585
R498 B.n258 B.n257 585
R499 B.n421 B.n420 585
R500 B.n420 B.n419 585
R501 B.n422 B.n255 585
R502 B.n255 B.n254 585
R503 B.n424 B.n423 585
R504 B.n425 B.n424 585
R505 B.n249 B.n248 585
R506 B.n250 B.n249 585
R507 B.n433 B.n432 585
R508 B.n432 B.n431 585
R509 B.n434 B.n247 585
R510 B.n247 B.n246 585
R511 B.n436 B.n435 585
R512 B.n437 B.n436 585
R513 B.n241 B.n240 585
R514 B.n242 B.n241 585
R515 B.n445 B.n444 585
R516 B.n444 B.n443 585
R517 B.n446 B.n239 585
R518 B.n239 B.n238 585
R519 B.n448 B.n447 585
R520 B.n449 B.n448 585
R521 B.n233 B.n232 585
R522 B.n234 B.n233 585
R523 B.n457 B.n456 585
R524 B.n456 B.n455 585
R525 B.n458 B.n231 585
R526 B.n231 B.n230 585
R527 B.n460 B.n459 585
R528 B.n461 B.n460 585
R529 B.n225 B.n224 585
R530 B.n226 B.n225 585
R531 B.n469 B.n468 585
R532 B.n468 B.n467 585
R533 B.n470 B.n223 585
R534 B.n223 B.n222 585
R535 B.n472 B.n471 585
R536 B.n473 B.n472 585
R537 B.n217 B.n216 585
R538 B.n218 B.n217 585
R539 B.n481 B.n480 585
R540 B.n480 B.n479 585
R541 B.n482 B.n215 585
R542 B.n215 B.n214 585
R543 B.n484 B.n483 585
R544 B.n485 B.n484 585
R545 B.n209 B.n208 585
R546 B.n210 B.n209 585
R547 B.n493 B.n492 585
R548 B.n492 B.n491 585
R549 B.n494 B.n207 585
R550 B.n207 B.n206 585
R551 B.n496 B.n495 585
R552 B.n497 B.n496 585
R553 B.n201 B.n200 585
R554 B.n202 B.n201 585
R555 B.n505 B.n504 585
R556 B.n504 B.n503 585
R557 B.n506 B.n199 585
R558 B.n199 B.n198 585
R559 B.n508 B.n507 585
R560 B.n509 B.n508 585
R561 B.n193 B.n192 585
R562 B.n194 B.n193 585
R563 B.n517 B.n516 585
R564 B.n516 B.n515 585
R565 B.n518 B.n191 585
R566 B.n191 B.n190 585
R567 B.n520 B.n519 585
R568 B.n521 B.n520 585
R569 B.n185 B.n184 585
R570 B.n186 B.n185 585
R571 B.n530 B.n529 585
R572 B.n529 B.n528 585
R573 B.n531 B.n183 585
R574 B.n183 B.n182 585
R575 B.n533 B.n532 585
R576 B.n534 B.n533 585
R577 B.n2 B.n0 585
R578 B.n4 B.n2 585
R579 B.n3 B.n1 585
R580 B.n724 B.n3 585
R581 B.n722 B.n721 585
R582 B.n723 B.n722 585
R583 B.n720 B.n9 585
R584 B.n9 B.n8 585
R585 B.n719 B.n718 585
R586 B.n718 B.n717 585
R587 B.n11 B.n10 585
R588 B.n716 B.n11 585
R589 B.n714 B.n713 585
R590 B.n715 B.n714 585
R591 B.n712 B.n16 585
R592 B.n16 B.n15 585
R593 B.n711 B.n710 585
R594 B.n710 B.n709 585
R595 B.n18 B.n17 585
R596 B.n708 B.n18 585
R597 B.n706 B.n705 585
R598 B.n707 B.n706 585
R599 B.n704 B.n23 585
R600 B.n23 B.n22 585
R601 B.n703 B.n702 585
R602 B.n702 B.n701 585
R603 B.n25 B.n24 585
R604 B.n700 B.n25 585
R605 B.n698 B.n697 585
R606 B.n699 B.n698 585
R607 B.n696 B.n30 585
R608 B.n30 B.n29 585
R609 B.n695 B.n694 585
R610 B.n694 B.n693 585
R611 B.n32 B.n31 585
R612 B.n692 B.n32 585
R613 B.n690 B.n689 585
R614 B.n691 B.n690 585
R615 B.n688 B.n37 585
R616 B.n37 B.n36 585
R617 B.n687 B.n686 585
R618 B.n686 B.n685 585
R619 B.n39 B.n38 585
R620 B.n684 B.n39 585
R621 B.n682 B.n681 585
R622 B.n683 B.n682 585
R623 B.n680 B.n44 585
R624 B.n44 B.n43 585
R625 B.n679 B.n678 585
R626 B.n678 B.n677 585
R627 B.n46 B.n45 585
R628 B.n676 B.n46 585
R629 B.n674 B.n673 585
R630 B.n675 B.n674 585
R631 B.n672 B.n51 585
R632 B.n51 B.n50 585
R633 B.n671 B.n670 585
R634 B.n670 B.n669 585
R635 B.n53 B.n52 585
R636 B.n668 B.n53 585
R637 B.n666 B.n665 585
R638 B.n667 B.n666 585
R639 B.n664 B.n58 585
R640 B.n58 B.n57 585
R641 B.n663 B.n662 585
R642 B.n662 B.n661 585
R643 B.n60 B.n59 585
R644 B.n660 B.n60 585
R645 B.n658 B.n657 585
R646 B.n659 B.n658 585
R647 B.n656 B.n65 585
R648 B.n65 B.n64 585
R649 B.n655 B.n654 585
R650 B.n654 B.n653 585
R651 B.n67 B.n66 585
R652 B.n652 B.n67 585
R653 B.n650 B.n649 585
R654 B.n651 B.n650 585
R655 B.n648 B.n72 585
R656 B.n72 B.n71 585
R657 B.n647 B.n646 585
R658 B.n646 B.n645 585
R659 B.n74 B.n73 585
R660 B.n644 B.n74 585
R661 B.n642 B.n641 585
R662 B.n643 B.n642 585
R663 B.n640 B.n79 585
R664 B.n79 B.n78 585
R665 B.n639 B.n638 585
R666 B.n638 B.n637 585
R667 B.n81 B.n80 585
R668 B.n636 B.n81 585
R669 B.n634 B.n633 585
R670 B.n635 B.n634 585
R671 B.n632 B.n86 585
R672 B.n86 B.n85 585
R673 B.n631 B.n630 585
R674 B.n630 B.n629 585
R675 B.n88 B.n87 585
R676 B.n628 B.n88 585
R677 B.n626 B.n625 585
R678 B.n627 B.n626 585
R679 B.n624 B.n93 585
R680 B.n93 B.n92 585
R681 B.n623 B.n622 585
R682 B.n622 B.n621 585
R683 B.n95 B.n94 585
R684 B.n620 B.n95 585
R685 B.n618 B.n617 585
R686 B.n619 B.n618 585
R687 B.n616 B.n100 585
R688 B.n100 B.n99 585
R689 B.n615 B.n614 585
R690 B.n614 B.n613 585
R691 B.n727 B.n726 585
R692 B.n726 B.n725 585
R693 B.n372 B.n289 454.062
R694 B.n614 B.n102 454.062
R695 B.n370 B.n291 454.062
R696 B.n610 B.n103 454.062
R697 B.n612 B.n611 256.663
R698 B.n612 B.n117 256.663
R699 B.n612 B.n116 256.663
R700 B.n612 B.n115 256.663
R701 B.n612 B.n114 256.663
R702 B.n612 B.n113 256.663
R703 B.n612 B.n112 256.663
R704 B.n612 B.n111 256.663
R705 B.n612 B.n110 256.663
R706 B.n612 B.n109 256.663
R707 B.n612 B.n108 256.663
R708 B.n612 B.n107 256.663
R709 B.n612 B.n106 256.663
R710 B.n612 B.n105 256.663
R711 B.n612 B.n104 256.663
R712 B.n309 B.n290 256.663
R713 B.n312 B.n290 256.663
R714 B.n318 B.n290 256.663
R715 B.n320 B.n290 256.663
R716 B.n329 B.n290 256.663
R717 B.n331 B.n290 256.663
R718 B.n337 B.n290 256.663
R719 B.n339 B.n290 256.663
R720 B.n345 B.n290 256.663
R721 B.n347 B.n290 256.663
R722 B.n354 B.n290 256.663
R723 B.n356 B.n290 256.663
R724 B.n362 B.n290 256.663
R725 B.n365 B.n290 256.663
R726 B.n297 B.t10 208.487
R727 B.n324 B.t18 208.487
R728 B.n122 B.t14 208.487
R729 B.n119 B.t21 208.487
R730 B.n297 B.t13 201.767
R731 B.n324 B.t20 201.767
R732 B.n122 B.t16 201.767
R733 B.n119 B.t22 201.767
R734 B.n371 B.n290 200.613
R735 B.n613 B.n612 200.613
R736 B.n372 B.n287 163.367
R737 B.n376 B.n287 163.367
R738 B.n376 B.n281 163.367
R739 B.n384 B.n281 163.367
R740 B.n384 B.n279 163.367
R741 B.n388 B.n279 163.367
R742 B.n388 B.n273 163.367
R743 B.n396 B.n273 163.367
R744 B.n396 B.n271 163.367
R745 B.n400 B.n271 163.367
R746 B.n400 B.n265 163.367
R747 B.n408 B.n265 163.367
R748 B.n408 B.n263 163.367
R749 B.n412 B.n263 163.367
R750 B.n412 B.n257 163.367
R751 B.n420 B.n257 163.367
R752 B.n420 B.n255 163.367
R753 B.n424 B.n255 163.367
R754 B.n424 B.n249 163.367
R755 B.n432 B.n249 163.367
R756 B.n432 B.n247 163.367
R757 B.n436 B.n247 163.367
R758 B.n436 B.n241 163.367
R759 B.n444 B.n241 163.367
R760 B.n444 B.n239 163.367
R761 B.n448 B.n239 163.367
R762 B.n448 B.n233 163.367
R763 B.n456 B.n233 163.367
R764 B.n456 B.n231 163.367
R765 B.n460 B.n231 163.367
R766 B.n460 B.n225 163.367
R767 B.n468 B.n225 163.367
R768 B.n468 B.n223 163.367
R769 B.n472 B.n223 163.367
R770 B.n472 B.n217 163.367
R771 B.n480 B.n217 163.367
R772 B.n480 B.n215 163.367
R773 B.n484 B.n215 163.367
R774 B.n484 B.n209 163.367
R775 B.n492 B.n209 163.367
R776 B.n492 B.n207 163.367
R777 B.n496 B.n207 163.367
R778 B.n496 B.n201 163.367
R779 B.n504 B.n201 163.367
R780 B.n504 B.n199 163.367
R781 B.n508 B.n199 163.367
R782 B.n508 B.n193 163.367
R783 B.n516 B.n193 163.367
R784 B.n516 B.n191 163.367
R785 B.n520 B.n191 163.367
R786 B.n520 B.n185 163.367
R787 B.n529 B.n185 163.367
R788 B.n529 B.n183 163.367
R789 B.n533 B.n183 163.367
R790 B.n533 B.n2 163.367
R791 B.n726 B.n2 163.367
R792 B.n726 B.n3 163.367
R793 B.n722 B.n3 163.367
R794 B.n722 B.n9 163.367
R795 B.n718 B.n9 163.367
R796 B.n718 B.n11 163.367
R797 B.n714 B.n11 163.367
R798 B.n714 B.n16 163.367
R799 B.n710 B.n16 163.367
R800 B.n710 B.n18 163.367
R801 B.n706 B.n18 163.367
R802 B.n706 B.n23 163.367
R803 B.n702 B.n23 163.367
R804 B.n702 B.n25 163.367
R805 B.n698 B.n25 163.367
R806 B.n698 B.n30 163.367
R807 B.n694 B.n30 163.367
R808 B.n694 B.n32 163.367
R809 B.n690 B.n32 163.367
R810 B.n690 B.n37 163.367
R811 B.n686 B.n37 163.367
R812 B.n686 B.n39 163.367
R813 B.n682 B.n39 163.367
R814 B.n682 B.n44 163.367
R815 B.n678 B.n44 163.367
R816 B.n678 B.n46 163.367
R817 B.n674 B.n46 163.367
R818 B.n674 B.n51 163.367
R819 B.n670 B.n51 163.367
R820 B.n670 B.n53 163.367
R821 B.n666 B.n53 163.367
R822 B.n666 B.n58 163.367
R823 B.n662 B.n58 163.367
R824 B.n662 B.n60 163.367
R825 B.n658 B.n60 163.367
R826 B.n658 B.n65 163.367
R827 B.n654 B.n65 163.367
R828 B.n654 B.n67 163.367
R829 B.n650 B.n67 163.367
R830 B.n650 B.n72 163.367
R831 B.n646 B.n72 163.367
R832 B.n646 B.n74 163.367
R833 B.n642 B.n74 163.367
R834 B.n642 B.n79 163.367
R835 B.n638 B.n79 163.367
R836 B.n638 B.n81 163.367
R837 B.n634 B.n81 163.367
R838 B.n634 B.n86 163.367
R839 B.n630 B.n86 163.367
R840 B.n630 B.n88 163.367
R841 B.n626 B.n88 163.367
R842 B.n626 B.n93 163.367
R843 B.n622 B.n93 163.367
R844 B.n622 B.n95 163.367
R845 B.n618 B.n95 163.367
R846 B.n618 B.n100 163.367
R847 B.n614 B.n100 163.367
R848 B.n311 B.n310 163.367
R849 B.n313 B.n311 163.367
R850 B.n317 B.n306 163.367
R851 B.n321 B.n319 163.367
R852 B.n328 B.n304 163.367
R853 B.n332 B.n330 163.367
R854 B.n336 B.n302 163.367
R855 B.n340 B.n338 163.367
R856 B.n344 B.n300 163.367
R857 B.n348 B.n346 163.367
R858 B.n353 B.n296 163.367
R859 B.n357 B.n355 163.367
R860 B.n361 B.n294 163.367
R861 B.n364 B.n363 163.367
R862 B.n366 B.n291 163.367
R863 B.n370 B.n285 163.367
R864 B.n378 B.n285 163.367
R865 B.n378 B.n283 163.367
R866 B.n382 B.n283 163.367
R867 B.n382 B.n276 163.367
R868 B.n390 B.n276 163.367
R869 B.n390 B.n274 163.367
R870 B.n394 B.n274 163.367
R871 B.n394 B.n269 163.367
R872 B.n402 B.n269 163.367
R873 B.n402 B.n267 163.367
R874 B.n406 B.n267 163.367
R875 B.n406 B.n261 163.367
R876 B.n414 B.n261 163.367
R877 B.n414 B.n259 163.367
R878 B.n418 B.n259 163.367
R879 B.n418 B.n253 163.367
R880 B.n426 B.n253 163.367
R881 B.n426 B.n251 163.367
R882 B.n430 B.n251 163.367
R883 B.n430 B.n245 163.367
R884 B.n438 B.n245 163.367
R885 B.n438 B.n243 163.367
R886 B.n442 B.n243 163.367
R887 B.n442 B.n237 163.367
R888 B.n450 B.n237 163.367
R889 B.n450 B.n235 163.367
R890 B.n454 B.n235 163.367
R891 B.n454 B.n229 163.367
R892 B.n462 B.n229 163.367
R893 B.n462 B.n227 163.367
R894 B.n466 B.n227 163.367
R895 B.n466 B.n221 163.367
R896 B.n474 B.n221 163.367
R897 B.n474 B.n219 163.367
R898 B.n478 B.n219 163.367
R899 B.n478 B.n213 163.367
R900 B.n486 B.n213 163.367
R901 B.n486 B.n211 163.367
R902 B.n490 B.n211 163.367
R903 B.n490 B.n205 163.367
R904 B.n498 B.n205 163.367
R905 B.n498 B.n203 163.367
R906 B.n502 B.n203 163.367
R907 B.n502 B.n197 163.367
R908 B.n510 B.n197 163.367
R909 B.n510 B.n195 163.367
R910 B.n514 B.n195 163.367
R911 B.n514 B.n189 163.367
R912 B.n522 B.n189 163.367
R913 B.n522 B.n187 163.367
R914 B.n527 B.n187 163.367
R915 B.n527 B.n181 163.367
R916 B.n535 B.n181 163.367
R917 B.n536 B.n535 163.367
R918 B.n536 B.n5 163.367
R919 B.n6 B.n5 163.367
R920 B.n7 B.n6 163.367
R921 B.n541 B.n7 163.367
R922 B.n541 B.n12 163.367
R923 B.n13 B.n12 163.367
R924 B.n14 B.n13 163.367
R925 B.n546 B.n14 163.367
R926 B.n546 B.n19 163.367
R927 B.n20 B.n19 163.367
R928 B.n21 B.n20 163.367
R929 B.n551 B.n21 163.367
R930 B.n551 B.n26 163.367
R931 B.n27 B.n26 163.367
R932 B.n28 B.n27 163.367
R933 B.n556 B.n28 163.367
R934 B.n556 B.n33 163.367
R935 B.n34 B.n33 163.367
R936 B.n35 B.n34 163.367
R937 B.n561 B.n35 163.367
R938 B.n561 B.n40 163.367
R939 B.n41 B.n40 163.367
R940 B.n42 B.n41 163.367
R941 B.n566 B.n42 163.367
R942 B.n566 B.n47 163.367
R943 B.n48 B.n47 163.367
R944 B.n49 B.n48 163.367
R945 B.n571 B.n49 163.367
R946 B.n571 B.n54 163.367
R947 B.n55 B.n54 163.367
R948 B.n56 B.n55 163.367
R949 B.n576 B.n56 163.367
R950 B.n576 B.n61 163.367
R951 B.n62 B.n61 163.367
R952 B.n63 B.n62 163.367
R953 B.n581 B.n63 163.367
R954 B.n581 B.n68 163.367
R955 B.n69 B.n68 163.367
R956 B.n70 B.n69 163.367
R957 B.n586 B.n70 163.367
R958 B.n586 B.n75 163.367
R959 B.n76 B.n75 163.367
R960 B.n77 B.n76 163.367
R961 B.n591 B.n77 163.367
R962 B.n591 B.n82 163.367
R963 B.n83 B.n82 163.367
R964 B.n84 B.n83 163.367
R965 B.n596 B.n84 163.367
R966 B.n596 B.n89 163.367
R967 B.n90 B.n89 163.367
R968 B.n91 B.n90 163.367
R969 B.n601 B.n91 163.367
R970 B.n601 B.n96 163.367
R971 B.n97 B.n96 163.367
R972 B.n98 B.n97 163.367
R973 B.n606 B.n98 163.367
R974 B.n606 B.n103 163.367
R975 B.n127 B.n126 163.367
R976 B.n131 B.n130 163.367
R977 B.n135 B.n134 163.367
R978 B.n139 B.n138 163.367
R979 B.n143 B.n142 163.367
R980 B.n147 B.n146 163.367
R981 B.n151 B.n150 163.367
R982 B.n155 B.n154 163.367
R983 B.n159 B.n158 163.367
R984 B.n163 B.n162 163.367
R985 B.n167 B.n166 163.367
R986 B.n171 B.n170 163.367
R987 B.n175 B.n174 163.367
R988 B.n177 B.n118 163.367
R989 B.n298 B.t12 149.208
R990 B.n325 B.t19 149.208
R991 B.n123 B.t17 149.208
R992 B.n120 B.t23 149.208
R993 B.n371 B.n286 114.636
R994 B.n377 B.n286 114.636
R995 B.n377 B.n282 114.636
R996 B.n383 B.n282 114.636
R997 B.n383 B.n277 114.636
R998 B.n389 B.n277 114.636
R999 B.n389 B.n278 114.636
R1000 B.n395 B.n270 114.636
R1001 B.n401 B.n270 114.636
R1002 B.n401 B.n266 114.636
R1003 B.n407 B.n266 114.636
R1004 B.n407 B.n262 114.636
R1005 B.n413 B.n262 114.636
R1006 B.n413 B.n258 114.636
R1007 B.n419 B.n258 114.636
R1008 B.n419 B.n254 114.636
R1009 B.n425 B.n254 114.636
R1010 B.n431 B.n250 114.636
R1011 B.n431 B.n246 114.636
R1012 B.n437 B.n246 114.636
R1013 B.n437 B.n242 114.636
R1014 B.n443 B.n242 114.636
R1015 B.n443 B.n238 114.636
R1016 B.n449 B.n238 114.636
R1017 B.n455 B.n234 114.636
R1018 B.n455 B.n230 114.636
R1019 B.n461 B.n230 114.636
R1020 B.n461 B.n226 114.636
R1021 B.n467 B.n226 114.636
R1022 B.n467 B.n222 114.636
R1023 B.n473 B.n222 114.636
R1024 B.n479 B.n218 114.636
R1025 B.n479 B.n214 114.636
R1026 B.n485 B.n214 114.636
R1027 B.n485 B.n210 114.636
R1028 B.n491 B.n210 114.636
R1029 B.n491 B.n206 114.636
R1030 B.n497 B.n206 114.636
R1031 B.n503 B.n202 114.636
R1032 B.n503 B.n198 114.636
R1033 B.n509 B.n198 114.636
R1034 B.n509 B.n194 114.636
R1035 B.n515 B.n194 114.636
R1036 B.n515 B.n190 114.636
R1037 B.n521 B.n190 114.636
R1038 B.n528 B.n186 114.636
R1039 B.n528 B.n182 114.636
R1040 B.n534 B.n182 114.636
R1041 B.n534 B.n4 114.636
R1042 B.n725 B.n4 114.636
R1043 B.n725 B.n724 114.636
R1044 B.n724 B.n723 114.636
R1045 B.n723 B.n8 114.636
R1046 B.n717 B.n8 114.636
R1047 B.n717 B.n716 114.636
R1048 B.n715 B.n15 114.636
R1049 B.n709 B.n15 114.636
R1050 B.n709 B.n708 114.636
R1051 B.n708 B.n707 114.636
R1052 B.n707 B.n22 114.636
R1053 B.n701 B.n22 114.636
R1054 B.n701 B.n700 114.636
R1055 B.n699 B.n29 114.636
R1056 B.n693 B.n29 114.636
R1057 B.n693 B.n692 114.636
R1058 B.n692 B.n691 114.636
R1059 B.n691 B.n36 114.636
R1060 B.n685 B.n36 114.636
R1061 B.n685 B.n684 114.636
R1062 B.n683 B.n43 114.636
R1063 B.n677 B.n43 114.636
R1064 B.n677 B.n676 114.636
R1065 B.n676 B.n675 114.636
R1066 B.n675 B.n50 114.636
R1067 B.n669 B.n50 114.636
R1068 B.n669 B.n668 114.636
R1069 B.n667 B.n57 114.636
R1070 B.n661 B.n57 114.636
R1071 B.n661 B.n660 114.636
R1072 B.n660 B.n659 114.636
R1073 B.n659 B.n64 114.636
R1074 B.n653 B.n64 114.636
R1075 B.n653 B.n652 114.636
R1076 B.n651 B.n71 114.636
R1077 B.n645 B.n71 114.636
R1078 B.n645 B.n644 114.636
R1079 B.n644 B.n643 114.636
R1080 B.n643 B.n78 114.636
R1081 B.n637 B.n78 114.636
R1082 B.n637 B.n636 114.636
R1083 B.n636 B.n635 114.636
R1084 B.n635 B.n85 114.636
R1085 B.n629 B.n85 114.636
R1086 B.n628 B.n627 114.636
R1087 B.n627 B.n92 114.636
R1088 B.n621 B.n92 114.636
R1089 B.n621 B.n620 114.636
R1090 B.n620 B.n619 114.636
R1091 B.n619 B.n99 114.636
R1092 B.n613 B.n99 114.636
R1093 B.n395 B.t11 74.1767
R1094 B.n629 B.t15 74.1767
R1095 B.n309 B.n289 71.676
R1096 B.n313 B.n312 71.676
R1097 B.n318 B.n317 71.676
R1098 B.n321 B.n320 71.676
R1099 B.n329 B.n328 71.676
R1100 B.n332 B.n331 71.676
R1101 B.n337 B.n336 71.676
R1102 B.n340 B.n339 71.676
R1103 B.n345 B.n344 71.676
R1104 B.n348 B.n347 71.676
R1105 B.n354 B.n353 71.676
R1106 B.n357 B.n356 71.676
R1107 B.n362 B.n361 71.676
R1108 B.n365 B.n364 71.676
R1109 B.n104 B.n102 71.676
R1110 B.n127 B.n105 71.676
R1111 B.n131 B.n106 71.676
R1112 B.n135 B.n107 71.676
R1113 B.n139 B.n108 71.676
R1114 B.n143 B.n109 71.676
R1115 B.n147 B.n110 71.676
R1116 B.n151 B.n111 71.676
R1117 B.n155 B.n112 71.676
R1118 B.n159 B.n113 71.676
R1119 B.n163 B.n114 71.676
R1120 B.n167 B.n115 71.676
R1121 B.n171 B.n116 71.676
R1122 B.n175 B.n117 71.676
R1123 B.n611 B.n118 71.676
R1124 B.n611 B.n610 71.676
R1125 B.n177 B.n117 71.676
R1126 B.n174 B.n116 71.676
R1127 B.n170 B.n115 71.676
R1128 B.n166 B.n114 71.676
R1129 B.n162 B.n113 71.676
R1130 B.n158 B.n112 71.676
R1131 B.n154 B.n111 71.676
R1132 B.n150 B.n110 71.676
R1133 B.n146 B.n109 71.676
R1134 B.n142 B.n108 71.676
R1135 B.n138 B.n107 71.676
R1136 B.n134 B.n106 71.676
R1137 B.n130 B.n105 71.676
R1138 B.n126 B.n104 71.676
R1139 B.n310 B.n309 71.676
R1140 B.n312 B.n306 71.676
R1141 B.n319 B.n318 71.676
R1142 B.n320 B.n304 71.676
R1143 B.n330 B.n329 71.676
R1144 B.n331 B.n302 71.676
R1145 B.n338 B.n337 71.676
R1146 B.n339 B.n300 71.676
R1147 B.n346 B.n345 71.676
R1148 B.n347 B.n296 71.676
R1149 B.n355 B.n354 71.676
R1150 B.n356 B.n294 71.676
R1151 B.n363 B.n362 71.676
R1152 B.n366 B.n365 71.676
R1153 B.t4 B.n186 67.4335
R1154 B.n716 B.t9 67.4335
R1155 B.t6 B.n202 64.0618
R1156 B.n700 B.t1 64.0618
R1157 B.n425 B.t8 60.6902
R1158 B.t0 B.n218 60.6902
R1159 B.n684 B.t7 60.6902
R1160 B.t3 B.n651 60.6902
R1161 B.n350 B.n298 59.5399
R1162 B.n326 B.n325 59.5399
R1163 B.n124 B.n123 59.5399
R1164 B.n121 B.n120 59.5399
R1165 B.n449 B.t5 57.3185
R1166 B.t5 B.n234 57.3185
R1167 B.n668 B.t2 57.3185
R1168 B.t2 B.n667 57.3185
R1169 B.t8 B.n250 53.9469
R1170 B.n473 B.t0 53.9469
R1171 B.t7 B.n683 53.9469
R1172 B.n652 B.t3 53.9469
R1173 B.n298 B.n297 52.5581
R1174 B.n325 B.n324 52.5581
R1175 B.n123 B.n122 52.5581
R1176 B.n120 B.n119 52.5581
R1177 B.n497 B.t6 50.5752
R1178 B.t1 B.n699 50.5752
R1179 B.n521 B.t4 47.2036
R1180 B.t9 B.n715 47.2036
R1181 B.n278 B.t11 40.4603
R1182 B.t15 B.n628 40.4603
R1183 B.n609 B.n608 29.5029
R1184 B.n615 B.n101 29.5029
R1185 B.n369 B.n368 29.5029
R1186 B.n373 B.n288 29.5029
R1187 B B.n727 18.0485
R1188 B.n125 B.n101 10.6151
R1189 B.n128 B.n125 10.6151
R1190 B.n129 B.n128 10.6151
R1191 B.n132 B.n129 10.6151
R1192 B.n133 B.n132 10.6151
R1193 B.n136 B.n133 10.6151
R1194 B.n137 B.n136 10.6151
R1195 B.n140 B.n137 10.6151
R1196 B.n141 B.n140 10.6151
R1197 B.n145 B.n144 10.6151
R1198 B.n148 B.n145 10.6151
R1199 B.n149 B.n148 10.6151
R1200 B.n152 B.n149 10.6151
R1201 B.n153 B.n152 10.6151
R1202 B.n156 B.n153 10.6151
R1203 B.n157 B.n156 10.6151
R1204 B.n160 B.n157 10.6151
R1205 B.n161 B.n160 10.6151
R1206 B.n165 B.n164 10.6151
R1207 B.n168 B.n165 10.6151
R1208 B.n169 B.n168 10.6151
R1209 B.n172 B.n169 10.6151
R1210 B.n173 B.n172 10.6151
R1211 B.n176 B.n173 10.6151
R1212 B.n178 B.n176 10.6151
R1213 B.n179 B.n178 10.6151
R1214 B.n609 B.n179 10.6151
R1215 B.n369 B.n284 10.6151
R1216 B.n379 B.n284 10.6151
R1217 B.n380 B.n379 10.6151
R1218 B.n381 B.n380 10.6151
R1219 B.n381 B.n275 10.6151
R1220 B.n391 B.n275 10.6151
R1221 B.n392 B.n391 10.6151
R1222 B.n393 B.n392 10.6151
R1223 B.n393 B.n268 10.6151
R1224 B.n403 B.n268 10.6151
R1225 B.n404 B.n403 10.6151
R1226 B.n405 B.n404 10.6151
R1227 B.n405 B.n260 10.6151
R1228 B.n415 B.n260 10.6151
R1229 B.n416 B.n415 10.6151
R1230 B.n417 B.n416 10.6151
R1231 B.n417 B.n252 10.6151
R1232 B.n427 B.n252 10.6151
R1233 B.n428 B.n427 10.6151
R1234 B.n429 B.n428 10.6151
R1235 B.n429 B.n244 10.6151
R1236 B.n439 B.n244 10.6151
R1237 B.n440 B.n439 10.6151
R1238 B.n441 B.n440 10.6151
R1239 B.n441 B.n236 10.6151
R1240 B.n451 B.n236 10.6151
R1241 B.n452 B.n451 10.6151
R1242 B.n453 B.n452 10.6151
R1243 B.n453 B.n228 10.6151
R1244 B.n463 B.n228 10.6151
R1245 B.n464 B.n463 10.6151
R1246 B.n465 B.n464 10.6151
R1247 B.n465 B.n220 10.6151
R1248 B.n475 B.n220 10.6151
R1249 B.n476 B.n475 10.6151
R1250 B.n477 B.n476 10.6151
R1251 B.n477 B.n212 10.6151
R1252 B.n487 B.n212 10.6151
R1253 B.n488 B.n487 10.6151
R1254 B.n489 B.n488 10.6151
R1255 B.n489 B.n204 10.6151
R1256 B.n499 B.n204 10.6151
R1257 B.n500 B.n499 10.6151
R1258 B.n501 B.n500 10.6151
R1259 B.n501 B.n196 10.6151
R1260 B.n511 B.n196 10.6151
R1261 B.n512 B.n511 10.6151
R1262 B.n513 B.n512 10.6151
R1263 B.n513 B.n188 10.6151
R1264 B.n523 B.n188 10.6151
R1265 B.n524 B.n523 10.6151
R1266 B.n526 B.n524 10.6151
R1267 B.n526 B.n525 10.6151
R1268 B.n525 B.n180 10.6151
R1269 B.n537 B.n180 10.6151
R1270 B.n538 B.n537 10.6151
R1271 B.n539 B.n538 10.6151
R1272 B.n540 B.n539 10.6151
R1273 B.n542 B.n540 10.6151
R1274 B.n543 B.n542 10.6151
R1275 B.n544 B.n543 10.6151
R1276 B.n545 B.n544 10.6151
R1277 B.n547 B.n545 10.6151
R1278 B.n548 B.n547 10.6151
R1279 B.n549 B.n548 10.6151
R1280 B.n550 B.n549 10.6151
R1281 B.n552 B.n550 10.6151
R1282 B.n553 B.n552 10.6151
R1283 B.n554 B.n553 10.6151
R1284 B.n555 B.n554 10.6151
R1285 B.n557 B.n555 10.6151
R1286 B.n558 B.n557 10.6151
R1287 B.n559 B.n558 10.6151
R1288 B.n560 B.n559 10.6151
R1289 B.n562 B.n560 10.6151
R1290 B.n563 B.n562 10.6151
R1291 B.n564 B.n563 10.6151
R1292 B.n565 B.n564 10.6151
R1293 B.n567 B.n565 10.6151
R1294 B.n568 B.n567 10.6151
R1295 B.n569 B.n568 10.6151
R1296 B.n570 B.n569 10.6151
R1297 B.n572 B.n570 10.6151
R1298 B.n573 B.n572 10.6151
R1299 B.n574 B.n573 10.6151
R1300 B.n575 B.n574 10.6151
R1301 B.n577 B.n575 10.6151
R1302 B.n578 B.n577 10.6151
R1303 B.n579 B.n578 10.6151
R1304 B.n580 B.n579 10.6151
R1305 B.n582 B.n580 10.6151
R1306 B.n583 B.n582 10.6151
R1307 B.n584 B.n583 10.6151
R1308 B.n585 B.n584 10.6151
R1309 B.n587 B.n585 10.6151
R1310 B.n588 B.n587 10.6151
R1311 B.n589 B.n588 10.6151
R1312 B.n590 B.n589 10.6151
R1313 B.n592 B.n590 10.6151
R1314 B.n593 B.n592 10.6151
R1315 B.n594 B.n593 10.6151
R1316 B.n595 B.n594 10.6151
R1317 B.n597 B.n595 10.6151
R1318 B.n598 B.n597 10.6151
R1319 B.n599 B.n598 10.6151
R1320 B.n600 B.n599 10.6151
R1321 B.n602 B.n600 10.6151
R1322 B.n603 B.n602 10.6151
R1323 B.n604 B.n603 10.6151
R1324 B.n605 B.n604 10.6151
R1325 B.n607 B.n605 10.6151
R1326 B.n608 B.n607 10.6151
R1327 B.n308 B.n288 10.6151
R1328 B.n308 B.n307 10.6151
R1329 B.n314 B.n307 10.6151
R1330 B.n315 B.n314 10.6151
R1331 B.n316 B.n315 10.6151
R1332 B.n316 B.n305 10.6151
R1333 B.n322 B.n305 10.6151
R1334 B.n323 B.n322 10.6151
R1335 B.n327 B.n323 10.6151
R1336 B.n333 B.n303 10.6151
R1337 B.n334 B.n333 10.6151
R1338 B.n335 B.n334 10.6151
R1339 B.n335 B.n301 10.6151
R1340 B.n341 B.n301 10.6151
R1341 B.n342 B.n341 10.6151
R1342 B.n343 B.n342 10.6151
R1343 B.n343 B.n299 10.6151
R1344 B.n349 B.n299 10.6151
R1345 B.n352 B.n351 10.6151
R1346 B.n352 B.n295 10.6151
R1347 B.n358 B.n295 10.6151
R1348 B.n359 B.n358 10.6151
R1349 B.n360 B.n359 10.6151
R1350 B.n360 B.n293 10.6151
R1351 B.n293 B.n292 10.6151
R1352 B.n367 B.n292 10.6151
R1353 B.n368 B.n367 10.6151
R1354 B.n374 B.n373 10.6151
R1355 B.n375 B.n374 10.6151
R1356 B.n375 B.n280 10.6151
R1357 B.n385 B.n280 10.6151
R1358 B.n386 B.n385 10.6151
R1359 B.n387 B.n386 10.6151
R1360 B.n387 B.n272 10.6151
R1361 B.n397 B.n272 10.6151
R1362 B.n398 B.n397 10.6151
R1363 B.n399 B.n398 10.6151
R1364 B.n399 B.n264 10.6151
R1365 B.n409 B.n264 10.6151
R1366 B.n410 B.n409 10.6151
R1367 B.n411 B.n410 10.6151
R1368 B.n411 B.n256 10.6151
R1369 B.n421 B.n256 10.6151
R1370 B.n422 B.n421 10.6151
R1371 B.n423 B.n422 10.6151
R1372 B.n423 B.n248 10.6151
R1373 B.n433 B.n248 10.6151
R1374 B.n434 B.n433 10.6151
R1375 B.n435 B.n434 10.6151
R1376 B.n435 B.n240 10.6151
R1377 B.n445 B.n240 10.6151
R1378 B.n446 B.n445 10.6151
R1379 B.n447 B.n446 10.6151
R1380 B.n447 B.n232 10.6151
R1381 B.n457 B.n232 10.6151
R1382 B.n458 B.n457 10.6151
R1383 B.n459 B.n458 10.6151
R1384 B.n459 B.n224 10.6151
R1385 B.n469 B.n224 10.6151
R1386 B.n470 B.n469 10.6151
R1387 B.n471 B.n470 10.6151
R1388 B.n471 B.n216 10.6151
R1389 B.n481 B.n216 10.6151
R1390 B.n482 B.n481 10.6151
R1391 B.n483 B.n482 10.6151
R1392 B.n483 B.n208 10.6151
R1393 B.n493 B.n208 10.6151
R1394 B.n494 B.n493 10.6151
R1395 B.n495 B.n494 10.6151
R1396 B.n495 B.n200 10.6151
R1397 B.n505 B.n200 10.6151
R1398 B.n506 B.n505 10.6151
R1399 B.n507 B.n506 10.6151
R1400 B.n507 B.n192 10.6151
R1401 B.n517 B.n192 10.6151
R1402 B.n518 B.n517 10.6151
R1403 B.n519 B.n518 10.6151
R1404 B.n519 B.n184 10.6151
R1405 B.n530 B.n184 10.6151
R1406 B.n531 B.n530 10.6151
R1407 B.n532 B.n531 10.6151
R1408 B.n532 B.n0 10.6151
R1409 B.n721 B.n1 10.6151
R1410 B.n721 B.n720 10.6151
R1411 B.n720 B.n719 10.6151
R1412 B.n719 B.n10 10.6151
R1413 B.n713 B.n10 10.6151
R1414 B.n713 B.n712 10.6151
R1415 B.n712 B.n711 10.6151
R1416 B.n711 B.n17 10.6151
R1417 B.n705 B.n17 10.6151
R1418 B.n705 B.n704 10.6151
R1419 B.n704 B.n703 10.6151
R1420 B.n703 B.n24 10.6151
R1421 B.n697 B.n24 10.6151
R1422 B.n697 B.n696 10.6151
R1423 B.n696 B.n695 10.6151
R1424 B.n695 B.n31 10.6151
R1425 B.n689 B.n31 10.6151
R1426 B.n689 B.n688 10.6151
R1427 B.n688 B.n687 10.6151
R1428 B.n687 B.n38 10.6151
R1429 B.n681 B.n38 10.6151
R1430 B.n681 B.n680 10.6151
R1431 B.n680 B.n679 10.6151
R1432 B.n679 B.n45 10.6151
R1433 B.n673 B.n45 10.6151
R1434 B.n673 B.n672 10.6151
R1435 B.n672 B.n671 10.6151
R1436 B.n671 B.n52 10.6151
R1437 B.n665 B.n52 10.6151
R1438 B.n665 B.n664 10.6151
R1439 B.n664 B.n663 10.6151
R1440 B.n663 B.n59 10.6151
R1441 B.n657 B.n59 10.6151
R1442 B.n657 B.n656 10.6151
R1443 B.n656 B.n655 10.6151
R1444 B.n655 B.n66 10.6151
R1445 B.n649 B.n66 10.6151
R1446 B.n649 B.n648 10.6151
R1447 B.n648 B.n647 10.6151
R1448 B.n647 B.n73 10.6151
R1449 B.n641 B.n73 10.6151
R1450 B.n641 B.n640 10.6151
R1451 B.n640 B.n639 10.6151
R1452 B.n639 B.n80 10.6151
R1453 B.n633 B.n80 10.6151
R1454 B.n633 B.n632 10.6151
R1455 B.n632 B.n631 10.6151
R1456 B.n631 B.n87 10.6151
R1457 B.n625 B.n87 10.6151
R1458 B.n625 B.n624 10.6151
R1459 B.n624 B.n623 10.6151
R1460 B.n623 B.n94 10.6151
R1461 B.n617 B.n94 10.6151
R1462 B.n617 B.n616 10.6151
R1463 B.n616 B.n615 10.6151
R1464 B.n141 B.n124 9.36635
R1465 B.n164 B.n121 9.36635
R1466 B.n327 B.n326 9.36635
R1467 B.n351 B.n350 9.36635
R1468 B.n727 B.n0 2.81026
R1469 B.n727 B.n1 2.81026
R1470 B.n144 B.n124 1.24928
R1471 B.n161 B.n121 1.24928
R1472 B.n326 B.n303 1.24928
R1473 B.n350 B.n349 1.24928
R1474 VP.n23 VP.n20 161.3
R1475 VP.n25 VP.n24 161.3
R1476 VP.n26 VP.n19 161.3
R1477 VP.n28 VP.n27 161.3
R1478 VP.n29 VP.n18 161.3
R1479 VP.n32 VP.n31 161.3
R1480 VP.n33 VP.n17 161.3
R1481 VP.n35 VP.n34 161.3
R1482 VP.n36 VP.n16 161.3
R1483 VP.n38 VP.n37 161.3
R1484 VP.n40 VP.n39 161.3
R1485 VP.n41 VP.n14 161.3
R1486 VP.n43 VP.n42 161.3
R1487 VP.n44 VP.n13 161.3
R1488 VP.n46 VP.n45 161.3
R1489 VP.n47 VP.n12 161.3
R1490 VP.n86 VP.n0 161.3
R1491 VP.n85 VP.n84 161.3
R1492 VP.n83 VP.n1 161.3
R1493 VP.n82 VP.n81 161.3
R1494 VP.n80 VP.n2 161.3
R1495 VP.n79 VP.n78 161.3
R1496 VP.n77 VP.n76 161.3
R1497 VP.n75 VP.n4 161.3
R1498 VP.n74 VP.n73 161.3
R1499 VP.n72 VP.n5 161.3
R1500 VP.n71 VP.n70 161.3
R1501 VP.n68 VP.n6 161.3
R1502 VP.n67 VP.n66 161.3
R1503 VP.n65 VP.n7 161.3
R1504 VP.n64 VP.n63 161.3
R1505 VP.n62 VP.n8 161.3
R1506 VP.n60 VP.n59 161.3
R1507 VP.n58 VP.n9 161.3
R1508 VP.n57 VP.n56 161.3
R1509 VP.n55 VP.n10 161.3
R1510 VP.n54 VP.n53 161.3
R1511 VP.n52 VP.n11 161.3
R1512 VP.n51 VP.n50 102.438
R1513 VP.n88 VP.n87 102.438
R1514 VP.n49 VP.n48 102.438
R1515 VP.n56 VP.n55 56.5193
R1516 VP.n81 VP.n1 56.5193
R1517 VP.n42 VP.n13 56.5193
R1518 VP.n63 VP.n7 50.6917
R1519 VP.n75 VP.n74 50.6917
R1520 VP.n36 VP.n35 50.6917
R1521 VP.n24 VP.n19 50.6917
R1522 VP.n22 VP.n21 49.8376
R1523 VP.n21 VP.t9 45.7749
R1524 VP.n51 VP.n49 43.7155
R1525 VP.n67 VP.n7 30.2951
R1526 VP.n74 VP.n5 30.2951
R1527 VP.n35 VP.n17 30.2951
R1528 VP.n28 VP.n19 30.2951
R1529 VP.n54 VP.n11 24.4675
R1530 VP.n55 VP.n54 24.4675
R1531 VP.n56 VP.n9 24.4675
R1532 VP.n60 VP.n9 24.4675
R1533 VP.n63 VP.n62 24.4675
R1534 VP.n68 VP.n67 24.4675
R1535 VP.n70 VP.n5 24.4675
R1536 VP.n76 VP.n75 24.4675
R1537 VP.n80 VP.n79 24.4675
R1538 VP.n81 VP.n80 24.4675
R1539 VP.n85 VP.n1 24.4675
R1540 VP.n86 VP.n85 24.4675
R1541 VP.n46 VP.n13 24.4675
R1542 VP.n47 VP.n46 24.4675
R1543 VP.n37 VP.n36 24.4675
R1544 VP.n41 VP.n40 24.4675
R1545 VP.n42 VP.n41 24.4675
R1546 VP.n29 VP.n28 24.4675
R1547 VP.n31 VP.n17 24.4675
R1548 VP.n24 VP.n23 24.4675
R1549 VP.n62 VP.n61 22.5101
R1550 VP.n76 VP.n3 22.5101
R1551 VP.n37 VP.n15 22.5101
R1552 VP.n23 VP.n22 22.5101
R1553 VP.n50 VP.t1 12.6581
R1554 VP.n61 VP.t6 12.6581
R1555 VP.n69 VP.t4 12.6581
R1556 VP.n3 VP.t8 12.6581
R1557 VP.n87 VP.t7 12.6581
R1558 VP.n48 VP.t0 12.6581
R1559 VP.n15 VP.t2 12.6581
R1560 VP.n30 VP.t5 12.6581
R1561 VP.n22 VP.t3 12.6581
R1562 VP.n69 VP.n68 12.234
R1563 VP.n70 VP.n69 12.234
R1564 VP.n30 VP.n29 12.234
R1565 VP.n31 VP.n30 12.234
R1566 VP.n50 VP.n11 8.31928
R1567 VP.n87 VP.n86 8.31928
R1568 VP.n48 VP.n47 8.31928
R1569 VP.n21 VP.n20 6.95571
R1570 VP.n61 VP.n60 1.95786
R1571 VP.n79 VP.n3 1.95786
R1572 VP.n40 VP.n15 1.95786
R1573 VP.n49 VP.n12 0.278367
R1574 VP.n52 VP.n51 0.278367
R1575 VP.n88 VP.n0 0.278367
R1576 VP.n25 VP.n20 0.189894
R1577 VP.n26 VP.n25 0.189894
R1578 VP.n27 VP.n26 0.189894
R1579 VP.n27 VP.n18 0.189894
R1580 VP.n32 VP.n18 0.189894
R1581 VP.n33 VP.n32 0.189894
R1582 VP.n34 VP.n33 0.189894
R1583 VP.n34 VP.n16 0.189894
R1584 VP.n38 VP.n16 0.189894
R1585 VP.n39 VP.n38 0.189894
R1586 VP.n39 VP.n14 0.189894
R1587 VP.n43 VP.n14 0.189894
R1588 VP.n44 VP.n43 0.189894
R1589 VP.n45 VP.n44 0.189894
R1590 VP.n45 VP.n12 0.189894
R1591 VP.n53 VP.n52 0.189894
R1592 VP.n53 VP.n10 0.189894
R1593 VP.n57 VP.n10 0.189894
R1594 VP.n58 VP.n57 0.189894
R1595 VP.n59 VP.n58 0.189894
R1596 VP.n59 VP.n8 0.189894
R1597 VP.n64 VP.n8 0.189894
R1598 VP.n65 VP.n64 0.189894
R1599 VP.n66 VP.n65 0.189894
R1600 VP.n66 VP.n6 0.189894
R1601 VP.n71 VP.n6 0.189894
R1602 VP.n72 VP.n71 0.189894
R1603 VP.n73 VP.n72 0.189894
R1604 VP.n73 VP.n4 0.189894
R1605 VP.n77 VP.n4 0.189894
R1606 VP.n78 VP.n77 0.189894
R1607 VP.n78 VP.n2 0.189894
R1608 VP.n82 VP.n2 0.189894
R1609 VP.n83 VP.n82 0.189894
R1610 VP.n84 VP.n83 0.189894
R1611 VP.n84 VP.n0 0.189894
R1612 VP VP.n88 0.153454
R1613 VDD1.n3 VDD1.t8 174.341
R1614 VDD1.n1 VDD1.t0 174.341
R1615 VDD1.n5 VDD1.n4 147.544
R1616 VDD1.n7 VDD1.n6 145.847
R1617 VDD1.n3 VDD1.n2 145.847
R1618 VDD1.n1 VDD1.n0 145.846
R1619 VDD1.n7 VDD1.n5 37.641
R1620 VDD1.n6 VDD1.t7 15.8405
R1621 VDD1.n6 VDD1.t9 15.8405
R1622 VDD1.n0 VDD1.t6 15.8405
R1623 VDD1.n0 VDD1.t4 15.8405
R1624 VDD1.n4 VDD1.t1 15.8405
R1625 VDD1.n4 VDD1.t2 15.8405
R1626 VDD1.n2 VDD1.t3 15.8405
R1627 VDD1.n2 VDD1.t5 15.8405
R1628 VDD1 VDD1.n7 1.69447
R1629 VDD1 VDD1.n1 0.642741
R1630 VDD1.n5 VDD1.n3 0.529206
C0 VN VTAIL 2.94863f
C1 VDD2 VP 0.564044f
C2 VDD1 VP 1.95184f
C3 VDD2 VDD1 2.03018f
C4 VP VTAIL 2.96276f
C5 VP VN 6.09564f
C6 VDD2 VTAIL 5.23454f
C7 VDD1 VTAIL 5.18261f
C8 VDD2 VN 1.55243f
C9 VDD1 VN 0.16048f
C10 VDD2 B 5.043318f
C11 VDD1 B 5.001898f
C12 VTAIL B 3.261116f
C13 VN B 16.05728f
C14 VP B 14.608521f
C15 VDD1.t0 B 0.167687f
C16 VDD1.t6 B 0.024418f
C17 VDD1.t4 B 0.024418f
C18 VDD1.n0 B 0.122093f
C19 VDD1.n1 B 0.800595f
C20 VDD1.t8 B 0.167687f
C21 VDD1.t3 B 0.024418f
C22 VDD1.t5 B 0.024418f
C23 VDD1.n2 B 0.122094f
C24 VDD1.n3 B 0.792635f
C25 VDD1.t1 B 0.024418f
C26 VDD1.t2 B 0.024418f
C27 VDD1.n4 B 0.127898f
C28 VDD1.n5 B 2.20991f
C29 VDD1.t7 B 0.024418f
C30 VDD1.t9 B 0.024418f
C31 VDD1.n6 B 0.122094f
C32 VDD1.n7 B 2.18587f
C33 VP.n0 B 0.037538f
C34 VP.t7 B 0.174082f
C35 VP.n1 B 0.03641f
C36 VP.n2 B 0.028472f
C37 VP.t8 B 0.174082f
C38 VP.n3 B 0.105327f
C39 VP.n4 B 0.028472f
C40 VP.n5 B 0.056896f
C41 VP.n6 B 0.028472f
C42 VP.t4 B 0.174082f
C43 VP.n7 B 0.027323f
C44 VP.n8 B 0.028472f
C45 VP.t6 B 0.174082f
C46 VP.n9 B 0.053065f
C47 VP.n10 B 0.028472f
C48 VP.n11 B 0.035774f
C49 VP.n12 B 0.037538f
C50 VP.t0 B 0.174082f
C51 VP.n13 B 0.03641f
C52 VP.n14 B 0.028472f
C53 VP.t2 B 0.174082f
C54 VP.n15 B 0.105327f
C55 VP.n16 B 0.028472f
C56 VP.n17 B 0.056896f
C57 VP.n18 B 0.028472f
C58 VP.t5 B 0.174082f
C59 VP.n19 B 0.027323f
C60 VP.n20 B 0.268738f
C61 VP.t3 B 0.174082f
C62 VP.t9 B 0.369575f
C63 VP.n21 B 0.173434f
C64 VP.n22 B 0.195855f
C65 VP.n23 B 0.05097f
C66 VP.n24 B 0.051981f
C67 VP.n25 B 0.028472f
C68 VP.n26 B 0.028472f
C69 VP.n27 B 0.028472f
C70 VP.n28 B 0.056896f
C71 VP.n29 B 0.039966f
C72 VP.n30 B 0.105327f
C73 VP.n31 B 0.039966f
C74 VP.n32 B 0.028472f
C75 VP.n33 B 0.028472f
C76 VP.n34 B 0.028472f
C77 VP.n35 B 0.027323f
C78 VP.n36 B 0.051981f
C79 VP.n37 B 0.05097f
C80 VP.n38 B 0.028472f
C81 VP.n39 B 0.028472f
C82 VP.n40 B 0.028963f
C83 VP.n41 B 0.053065f
C84 VP.n42 B 0.046724f
C85 VP.n43 B 0.028472f
C86 VP.n44 B 0.028472f
C87 VP.n45 B 0.028472f
C88 VP.n46 B 0.053065f
C89 VP.n47 B 0.035774f
C90 VP.n48 B 0.189768f
C91 VP.n49 B 1.28951f
C92 VP.t1 B 0.174082f
C93 VP.n50 B 0.189768f
C94 VP.n51 B 1.31293f
C95 VP.n52 B 0.037538f
C96 VP.n53 B 0.028472f
C97 VP.n54 B 0.053065f
C98 VP.n55 B 0.03641f
C99 VP.n56 B 0.046724f
C100 VP.n57 B 0.028472f
C101 VP.n58 B 0.028472f
C102 VP.n59 B 0.028472f
C103 VP.n60 B 0.028963f
C104 VP.n61 B 0.105327f
C105 VP.n62 B 0.05097f
C106 VP.n63 B 0.051981f
C107 VP.n64 B 0.028472f
C108 VP.n65 B 0.028472f
C109 VP.n66 B 0.028472f
C110 VP.n67 B 0.056896f
C111 VP.n68 B 0.039966f
C112 VP.n69 B 0.105327f
C113 VP.n70 B 0.039966f
C114 VP.n71 B 0.028472f
C115 VP.n72 B 0.028472f
C116 VP.n73 B 0.028472f
C117 VP.n74 B 0.027323f
C118 VP.n75 B 0.051981f
C119 VP.n76 B 0.05097f
C120 VP.n77 B 0.028472f
C121 VP.n78 B 0.028472f
C122 VP.n79 B 0.028963f
C123 VP.n80 B 0.053065f
C124 VP.n81 B 0.046724f
C125 VP.n82 B 0.028472f
C126 VP.n83 B 0.028472f
C127 VP.n84 B 0.028472f
C128 VP.n85 B 0.053065f
C129 VP.n86 B 0.035774f
C130 VP.n87 B 0.189768f
C131 VP.n88 B 0.04543f
C132 VDD2.t9 B 0.169841f
C133 VDD2.t8 B 0.024732f
C134 VDD2.t6 B 0.024732f
C135 VDD2.n0 B 0.123662f
C136 VDD2.n1 B 0.802815f
C137 VDD2.t1 B 0.024732f
C138 VDD2.t0 B 0.024732f
C139 VDD2.n2 B 0.129541f
C140 VDD2.n3 B 2.12877f
C141 VDD2.t7 B 0.164473f
C142 VDD2.n4 B 2.12097f
C143 VDD2.t4 B 0.024732f
C144 VDD2.t2 B 0.024732f
C145 VDD2.n5 B 0.123662f
C146 VDD2.n6 B 0.415668f
C147 VDD2.t5 B 0.024732f
C148 VDD2.t3 B 0.024732f
C149 VDD2.n7 B 0.129524f
C150 VTAIL.t6 B 0.039411f
C151 VTAIL.t7 B 0.039411f
C152 VTAIL.n0 B 0.161954f
C153 VTAIL.n1 B 0.703657f
C154 VTAIL.t18 B 0.228342f
C155 VTAIL.n2 B 0.812359f
C156 VTAIL.t0 B 0.039411f
C157 VTAIL.t16 B 0.039411f
C158 VTAIL.n3 B 0.161954f
C159 VTAIL.n4 B 0.861033f
C160 VTAIL.t14 B 0.039411f
C161 VTAIL.t19 B 0.039411f
C162 VTAIL.n5 B 0.161954f
C163 VTAIL.n6 B 1.84189f
C164 VTAIL.t8 B 0.039411f
C165 VTAIL.t13 B 0.039411f
C166 VTAIL.n7 B 0.161953f
C167 VTAIL.n8 B 1.84189f
C168 VTAIL.t4 B 0.039411f
C169 VTAIL.t9 B 0.039411f
C170 VTAIL.n9 B 0.161953f
C171 VTAIL.n10 B 0.861034f
C172 VTAIL.t10 B 0.228342f
C173 VTAIL.n11 B 0.812359f
C174 VTAIL.t15 B 0.039411f
C175 VTAIL.t1 B 0.039411f
C176 VTAIL.n12 B 0.161953f
C177 VTAIL.n13 B 0.771263f
C178 VTAIL.t17 B 0.039411f
C179 VTAIL.t2 B 0.039411f
C180 VTAIL.n14 B 0.161953f
C181 VTAIL.n15 B 0.861034f
C182 VTAIL.t3 B 0.228342f
C183 VTAIL.n16 B 1.58264f
C184 VTAIL.t11 B 0.228342f
C185 VTAIL.n17 B 1.58264f
C186 VTAIL.t12 B 0.039411f
C187 VTAIL.t5 B 0.039411f
C188 VTAIL.n18 B 0.161954f
C189 VTAIL.n19 B 0.628293f
C190 VN.n0 B 0.036963f
C191 VN.t9 B 0.171415f
C192 VN.n1 B 0.035852f
C193 VN.n2 B 0.028036f
C194 VN.t8 B 0.171415f
C195 VN.n3 B 0.103713f
C196 VN.n4 B 0.028036f
C197 VN.n5 B 0.056024f
C198 VN.n6 B 0.028036f
C199 VN.t3 B 0.171415f
C200 VN.n7 B 0.026905f
C201 VN.n8 B 0.264621f
C202 VN.t1 B 0.171415f
C203 VN.t0 B 0.363913f
C204 VN.n9 B 0.170777f
C205 VN.n10 B 0.192855f
C206 VN.n11 B 0.050189f
C207 VN.n12 B 0.051185f
C208 VN.n13 B 0.028036f
C209 VN.n14 B 0.028036f
C210 VN.n15 B 0.028036f
C211 VN.n16 B 0.056024f
C212 VN.n17 B 0.039354f
C213 VN.n18 B 0.103713f
C214 VN.n19 B 0.039354f
C215 VN.n20 B 0.028036f
C216 VN.n21 B 0.028036f
C217 VN.n22 B 0.028036f
C218 VN.n23 B 0.026905f
C219 VN.n24 B 0.051185f
C220 VN.n25 B 0.050189f
C221 VN.n26 B 0.028036f
C222 VN.n27 B 0.028036f
C223 VN.n28 B 0.028519f
C224 VN.n29 B 0.052253f
C225 VN.n30 B 0.046009f
C226 VN.n31 B 0.028036f
C227 VN.n32 B 0.028036f
C228 VN.n33 B 0.028036f
C229 VN.n34 B 0.052253f
C230 VN.n35 B 0.035226f
C231 VN.n36 B 0.186861f
C232 VN.n37 B 0.044734f
C233 VN.n38 B 0.036963f
C234 VN.t2 B 0.171415f
C235 VN.n39 B 0.035852f
C236 VN.n40 B 0.028036f
C237 VN.t5 B 0.171415f
C238 VN.n41 B 0.103713f
C239 VN.n42 B 0.028036f
C240 VN.n43 B 0.056024f
C241 VN.n44 B 0.028036f
C242 VN.t7 B 0.171415f
C243 VN.n45 B 0.026905f
C244 VN.n46 B 0.264621f
C245 VN.t4 B 0.171415f
C246 VN.t6 B 0.363913f
C247 VN.n47 B 0.170777f
C248 VN.n48 B 0.192855f
C249 VN.n49 B 0.050189f
C250 VN.n50 B 0.051185f
C251 VN.n51 B 0.028036f
C252 VN.n52 B 0.028036f
C253 VN.n53 B 0.028036f
C254 VN.n54 B 0.056024f
C255 VN.n55 B 0.039354f
C256 VN.n56 B 0.103713f
C257 VN.n57 B 0.039354f
C258 VN.n58 B 0.028036f
C259 VN.n59 B 0.028036f
C260 VN.n60 B 0.028036f
C261 VN.n61 B 0.026905f
C262 VN.n62 B 0.051185f
C263 VN.n63 B 0.050189f
C264 VN.n64 B 0.028036f
C265 VN.n65 B 0.028036f
C266 VN.n66 B 0.028519f
C267 VN.n67 B 0.052253f
C268 VN.n68 B 0.046009f
C269 VN.n69 B 0.028036f
C270 VN.n70 B 0.028036f
C271 VN.n71 B 0.028036f
C272 VN.n72 B 0.052253f
C273 VN.n73 B 0.035226f
C274 VN.n74 B 0.186861f
C275 VN.n75 B 1.28517f
.ends

