* NGSPICE file created from diff_pair_sample_0451.ext - technology: sky130A

.subckt diff_pair_sample_0451 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t9 VN.t0 VTAIL.t18 w_n5866_n2130# sky130_fd_pr__pfet_01v8 ad=0.95865 pd=6.14 as=2.2659 ps=12.4 w=5.81 l=3.75
X1 VDD2.t8 VN.t1 VTAIL.t17 w_n5866_n2130# sky130_fd_pr__pfet_01v8 ad=0.95865 pd=6.14 as=0.95865 ps=6.14 w=5.81 l=3.75
X2 B.t11 B.t9 B.t10 w_n5866_n2130# sky130_fd_pr__pfet_01v8 ad=2.2659 pd=12.4 as=0 ps=0 w=5.81 l=3.75
X3 VTAIL.t6 VP.t0 VDD1.t9 w_n5866_n2130# sky130_fd_pr__pfet_01v8 ad=0.95865 pd=6.14 as=0.95865 ps=6.14 w=5.81 l=3.75
X4 VTAIL.t16 VN.t2 VDD2.t7 w_n5866_n2130# sky130_fd_pr__pfet_01v8 ad=0.95865 pd=6.14 as=0.95865 ps=6.14 w=5.81 l=3.75
X5 VTAIL.t11 VN.t3 VDD2.t6 w_n5866_n2130# sky130_fd_pr__pfet_01v8 ad=0.95865 pd=6.14 as=0.95865 ps=6.14 w=5.81 l=3.75
X6 VDD1.t8 VP.t1 VTAIL.t4 w_n5866_n2130# sky130_fd_pr__pfet_01v8 ad=0.95865 pd=6.14 as=2.2659 ps=12.4 w=5.81 l=3.75
X7 VDD1.t7 VP.t2 VTAIL.t7 w_n5866_n2130# sky130_fd_pr__pfet_01v8 ad=0.95865 pd=6.14 as=0.95865 ps=6.14 w=5.81 l=3.75
X8 VDD2.t5 VN.t4 VTAIL.t19 w_n5866_n2130# sky130_fd_pr__pfet_01v8 ad=0.95865 pd=6.14 as=0.95865 ps=6.14 w=5.81 l=3.75
X9 B.t8 B.t6 B.t7 w_n5866_n2130# sky130_fd_pr__pfet_01v8 ad=2.2659 pd=12.4 as=0 ps=0 w=5.81 l=3.75
X10 VDD2.t4 VN.t5 VTAIL.t13 w_n5866_n2130# sky130_fd_pr__pfet_01v8 ad=0.95865 pd=6.14 as=2.2659 ps=12.4 w=5.81 l=3.75
X11 VTAIL.t14 VN.t6 VDD2.t3 w_n5866_n2130# sky130_fd_pr__pfet_01v8 ad=0.95865 pd=6.14 as=0.95865 ps=6.14 w=5.81 l=3.75
X12 VTAIL.t9 VP.t3 VDD1.t6 w_n5866_n2130# sky130_fd_pr__pfet_01v8 ad=0.95865 pd=6.14 as=0.95865 ps=6.14 w=5.81 l=3.75
X13 VTAIL.t5 VP.t4 VDD1.t5 w_n5866_n2130# sky130_fd_pr__pfet_01v8 ad=0.95865 pd=6.14 as=0.95865 ps=6.14 w=5.81 l=3.75
X14 B.t5 B.t3 B.t4 w_n5866_n2130# sky130_fd_pr__pfet_01v8 ad=2.2659 pd=12.4 as=0 ps=0 w=5.81 l=3.75
X15 VDD1.t4 VP.t5 VTAIL.t1 w_n5866_n2130# sky130_fd_pr__pfet_01v8 ad=2.2659 pd=12.4 as=0.95865 ps=6.14 w=5.81 l=3.75
X16 VDD1.t3 VP.t6 VTAIL.t3 w_n5866_n2130# sky130_fd_pr__pfet_01v8 ad=0.95865 pd=6.14 as=0.95865 ps=6.14 w=5.81 l=3.75
X17 VDD2.t2 VN.t7 VTAIL.t10 w_n5866_n2130# sky130_fd_pr__pfet_01v8 ad=2.2659 pd=12.4 as=0.95865 ps=6.14 w=5.81 l=3.75
X18 B.t2 B.t0 B.t1 w_n5866_n2130# sky130_fd_pr__pfet_01v8 ad=2.2659 pd=12.4 as=0 ps=0 w=5.81 l=3.75
X19 VTAIL.t8 VP.t7 VDD1.t2 w_n5866_n2130# sky130_fd_pr__pfet_01v8 ad=0.95865 pd=6.14 as=0.95865 ps=6.14 w=5.81 l=3.75
X20 VTAIL.t15 VN.t8 VDD2.t1 w_n5866_n2130# sky130_fd_pr__pfet_01v8 ad=0.95865 pd=6.14 as=0.95865 ps=6.14 w=5.81 l=3.75
X21 VDD2.t0 VN.t9 VTAIL.t12 w_n5866_n2130# sky130_fd_pr__pfet_01v8 ad=2.2659 pd=12.4 as=0.95865 ps=6.14 w=5.81 l=3.75
X22 VDD1.t1 VP.t8 VTAIL.t0 w_n5866_n2130# sky130_fd_pr__pfet_01v8 ad=2.2659 pd=12.4 as=0.95865 ps=6.14 w=5.81 l=3.75
X23 VDD1.t0 VP.t9 VTAIL.t2 w_n5866_n2130# sky130_fd_pr__pfet_01v8 ad=0.95865 pd=6.14 as=2.2659 ps=12.4 w=5.81 l=3.75
R0 VN.n108 VN.n107 161.3
R1 VN.n106 VN.n56 161.3
R2 VN.n105 VN.n104 161.3
R3 VN.n103 VN.n57 161.3
R4 VN.n102 VN.n101 161.3
R5 VN.n100 VN.n58 161.3
R6 VN.n99 VN.n98 161.3
R7 VN.n97 VN.n59 161.3
R8 VN.n96 VN.n95 161.3
R9 VN.n94 VN.n60 161.3
R10 VN.n93 VN.n92 161.3
R11 VN.n91 VN.n62 161.3
R12 VN.n90 VN.n89 161.3
R13 VN.n88 VN.n63 161.3
R14 VN.n87 VN.n86 161.3
R15 VN.n85 VN.n64 161.3
R16 VN.n84 VN.n83 161.3
R17 VN.n82 VN.n65 161.3
R18 VN.n81 VN.n80 161.3
R19 VN.n79 VN.n66 161.3
R20 VN.n78 VN.n77 161.3
R21 VN.n76 VN.n67 161.3
R22 VN.n75 VN.n74 161.3
R23 VN.n73 VN.n68 161.3
R24 VN.n72 VN.n71 161.3
R25 VN.n53 VN.n52 161.3
R26 VN.n51 VN.n1 161.3
R27 VN.n50 VN.n49 161.3
R28 VN.n48 VN.n2 161.3
R29 VN.n47 VN.n46 161.3
R30 VN.n45 VN.n3 161.3
R31 VN.n44 VN.n43 161.3
R32 VN.n42 VN.n4 161.3
R33 VN.n41 VN.n40 161.3
R34 VN.n38 VN.n5 161.3
R35 VN.n37 VN.n36 161.3
R36 VN.n35 VN.n6 161.3
R37 VN.n34 VN.n33 161.3
R38 VN.n32 VN.n7 161.3
R39 VN.n31 VN.n30 161.3
R40 VN.n29 VN.n8 161.3
R41 VN.n28 VN.n27 161.3
R42 VN.n26 VN.n9 161.3
R43 VN.n25 VN.n24 161.3
R44 VN.n23 VN.n10 161.3
R45 VN.n22 VN.n21 161.3
R46 VN.n20 VN.n11 161.3
R47 VN.n19 VN.n18 161.3
R48 VN.n17 VN.n12 161.3
R49 VN.n16 VN.n15 161.3
R50 VN.n54 VN.n0 82.238
R51 VN.n109 VN.n55 82.238
R52 VN.n14 VN.n13 70.8482
R53 VN.n70 VN.n69 70.8482
R54 VN.n69 VN.t5 70.3424
R55 VN.n13 VN.t7 70.3424
R56 VN VN.n109 54.9601
R57 VN.n46 VN.n2 52.1486
R58 VN.n101 VN.n57 52.1486
R59 VN.n21 VN.n20 44.3785
R60 VN.n33 VN.n6 44.3785
R61 VN.n77 VN.n76 44.3785
R62 VN.n89 VN.n62 44.3785
R63 VN.n27 VN.t1 37.3394
R64 VN.n14 VN.t3 37.3394
R65 VN.n39 VN.t2 37.3394
R66 VN.n0 VN.t0 37.3394
R67 VN.n83 VN.t4 37.3394
R68 VN.n70 VN.t8 37.3394
R69 VN.n61 VN.t6 37.3394
R70 VN.n55 VN.t9 37.3394
R71 VN.n21 VN.n10 36.6083
R72 VN.n33 VN.n32 36.6083
R73 VN.n77 VN.n66 36.6083
R74 VN.n89 VN.n88 36.6083
R75 VN.n46 VN.n45 28.8382
R76 VN.n101 VN.n100 28.8382
R77 VN.n15 VN.n12 24.4675
R78 VN.n19 VN.n12 24.4675
R79 VN.n20 VN.n19 24.4675
R80 VN.n25 VN.n10 24.4675
R81 VN.n26 VN.n25 24.4675
R82 VN.n27 VN.n26 24.4675
R83 VN.n27 VN.n8 24.4675
R84 VN.n31 VN.n8 24.4675
R85 VN.n32 VN.n31 24.4675
R86 VN.n37 VN.n6 24.4675
R87 VN.n38 VN.n37 24.4675
R88 VN.n40 VN.n38 24.4675
R89 VN.n44 VN.n4 24.4675
R90 VN.n45 VN.n44 24.4675
R91 VN.n50 VN.n2 24.4675
R92 VN.n51 VN.n50 24.4675
R93 VN.n52 VN.n51 24.4675
R94 VN.n76 VN.n75 24.4675
R95 VN.n75 VN.n68 24.4675
R96 VN.n71 VN.n68 24.4675
R97 VN.n88 VN.n87 24.4675
R98 VN.n87 VN.n64 24.4675
R99 VN.n83 VN.n64 24.4675
R100 VN.n83 VN.n82 24.4675
R101 VN.n82 VN.n81 24.4675
R102 VN.n81 VN.n66 24.4675
R103 VN.n100 VN.n99 24.4675
R104 VN.n99 VN.n59 24.4675
R105 VN.n95 VN.n94 24.4675
R106 VN.n94 VN.n93 24.4675
R107 VN.n93 VN.n62 24.4675
R108 VN.n107 VN.n106 24.4675
R109 VN.n106 VN.n105 24.4675
R110 VN.n105 VN.n57 24.4675
R111 VN.n39 VN.n4 20.5528
R112 VN.n61 VN.n59 20.5528
R113 VN.n52 VN.n0 7.82994
R114 VN.n107 VN.n55 7.82994
R115 VN.n15 VN.n14 3.91522
R116 VN.n40 VN.n39 3.91522
R117 VN.n71 VN.n70 3.91522
R118 VN.n95 VN.n61 3.91522
R119 VN.n72 VN.n69 3.22187
R120 VN.n16 VN.n13 3.22187
R121 VN.n109 VN.n108 0.354971
R122 VN.n54 VN.n53 0.354971
R123 VN VN.n54 0.26696
R124 VN.n108 VN.n56 0.189894
R125 VN.n104 VN.n56 0.189894
R126 VN.n104 VN.n103 0.189894
R127 VN.n103 VN.n102 0.189894
R128 VN.n102 VN.n58 0.189894
R129 VN.n98 VN.n58 0.189894
R130 VN.n98 VN.n97 0.189894
R131 VN.n97 VN.n96 0.189894
R132 VN.n96 VN.n60 0.189894
R133 VN.n92 VN.n60 0.189894
R134 VN.n92 VN.n91 0.189894
R135 VN.n91 VN.n90 0.189894
R136 VN.n90 VN.n63 0.189894
R137 VN.n86 VN.n63 0.189894
R138 VN.n86 VN.n85 0.189894
R139 VN.n85 VN.n84 0.189894
R140 VN.n84 VN.n65 0.189894
R141 VN.n80 VN.n65 0.189894
R142 VN.n80 VN.n79 0.189894
R143 VN.n79 VN.n78 0.189894
R144 VN.n78 VN.n67 0.189894
R145 VN.n74 VN.n67 0.189894
R146 VN.n74 VN.n73 0.189894
R147 VN.n73 VN.n72 0.189894
R148 VN.n17 VN.n16 0.189894
R149 VN.n18 VN.n17 0.189894
R150 VN.n18 VN.n11 0.189894
R151 VN.n22 VN.n11 0.189894
R152 VN.n23 VN.n22 0.189894
R153 VN.n24 VN.n23 0.189894
R154 VN.n24 VN.n9 0.189894
R155 VN.n28 VN.n9 0.189894
R156 VN.n29 VN.n28 0.189894
R157 VN.n30 VN.n29 0.189894
R158 VN.n30 VN.n7 0.189894
R159 VN.n34 VN.n7 0.189894
R160 VN.n35 VN.n34 0.189894
R161 VN.n36 VN.n35 0.189894
R162 VN.n36 VN.n5 0.189894
R163 VN.n41 VN.n5 0.189894
R164 VN.n42 VN.n41 0.189894
R165 VN.n43 VN.n42 0.189894
R166 VN.n43 VN.n3 0.189894
R167 VN.n47 VN.n3 0.189894
R168 VN.n48 VN.n47 0.189894
R169 VN.n49 VN.n48 0.189894
R170 VN.n49 VN.n1 0.189894
R171 VN.n53 VN.n1 0.189894
R172 VTAIL.n132 VTAIL.n131 756.745
R173 VTAIL.n30 VTAIL.n29 756.745
R174 VTAIL.n102 VTAIL.n101 756.745
R175 VTAIL.n68 VTAIL.n67 756.745
R176 VTAIL.n115 VTAIL.n114 585
R177 VTAIL.n117 VTAIL.n116 585
R178 VTAIL.n110 VTAIL.n109 585
R179 VTAIL.n123 VTAIL.n122 585
R180 VTAIL.n125 VTAIL.n124 585
R181 VTAIL.n106 VTAIL.n105 585
R182 VTAIL.n131 VTAIL.n130 585
R183 VTAIL.n13 VTAIL.n12 585
R184 VTAIL.n15 VTAIL.n14 585
R185 VTAIL.n8 VTAIL.n7 585
R186 VTAIL.n21 VTAIL.n20 585
R187 VTAIL.n23 VTAIL.n22 585
R188 VTAIL.n4 VTAIL.n3 585
R189 VTAIL.n29 VTAIL.n28 585
R190 VTAIL.n101 VTAIL.n100 585
R191 VTAIL.n76 VTAIL.n75 585
R192 VTAIL.n95 VTAIL.n94 585
R193 VTAIL.n93 VTAIL.n92 585
R194 VTAIL.n80 VTAIL.n79 585
R195 VTAIL.n87 VTAIL.n86 585
R196 VTAIL.n85 VTAIL.n84 585
R197 VTAIL.n67 VTAIL.n66 585
R198 VTAIL.n42 VTAIL.n41 585
R199 VTAIL.n61 VTAIL.n60 585
R200 VTAIL.n59 VTAIL.n58 585
R201 VTAIL.n46 VTAIL.n45 585
R202 VTAIL.n53 VTAIL.n52 585
R203 VTAIL.n51 VTAIL.n50 585
R204 VTAIL.n113 VTAIL.t18 329.175
R205 VTAIL.n11 VTAIL.t4 329.175
R206 VTAIL.n83 VTAIL.t2 329.175
R207 VTAIL.n49 VTAIL.t13 329.175
R208 VTAIL.n116 VTAIL.n115 171.744
R209 VTAIL.n116 VTAIL.n109 171.744
R210 VTAIL.n123 VTAIL.n109 171.744
R211 VTAIL.n124 VTAIL.n123 171.744
R212 VTAIL.n124 VTAIL.n105 171.744
R213 VTAIL.n131 VTAIL.n105 171.744
R214 VTAIL.n14 VTAIL.n13 171.744
R215 VTAIL.n14 VTAIL.n7 171.744
R216 VTAIL.n21 VTAIL.n7 171.744
R217 VTAIL.n22 VTAIL.n21 171.744
R218 VTAIL.n22 VTAIL.n3 171.744
R219 VTAIL.n29 VTAIL.n3 171.744
R220 VTAIL.n101 VTAIL.n75 171.744
R221 VTAIL.n94 VTAIL.n75 171.744
R222 VTAIL.n94 VTAIL.n93 171.744
R223 VTAIL.n93 VTAIL.n79 171.744
R224 VTAIL.n86 VTAIL.n79 171.744
R225 VTAIL.n86 VTAIL.n85 171.744
R226 VTAIL.n67 VTAIL.n41 171.744
R227 VTAIL.n60 VTAIL.n41 171.744
R228 VTAIL.n60 VTAIL.n59 171.744
R229 VTAIL.n59 VTAIL.n45 171.744
R230 VTAIL.n52 VTAIL.n45 171.744
R231 VTAIL.n52 VTAIL.n51 171.744
R232 VTAIL.n115 VTAIL.t18 85.8723
R233 VTAIL.n13 VTAIL.t4 85.8723
R234 VTAIL.n85 VTAIL.t2 85.8723
R235 VTAIL.n51 VTAIL.t13 85.8723
R236 VTAIL.n73 VTAIL.n72 78.2402
R237 VTAIL.n71 VTAIL.n70 78.2402
R238 VTAIL.n39 VTAIL.n38 78.2402
R239 VTAIL.n37 VTAIL.n36 78.2402
R240 VTAIL.n135 VTAIL.n134 78.2392
R241 VTAIL.n1 VTAIL.n0 78.2392
R242 VTAIL.n33 VTAIL.n32 78.2392
R243 VTAIL.n35 VTAIL.n34 78.2392
R244 VTAIL.n133 VTAIL.n132 34.3187
R245 VTAIL.n31 VTAIL.n30 34.3187
R246 VTAIL.n103 VTAIL.n102 34.3187
R247 VTAIL.n69 VTAIL.n68 34.3187
R248 VTAIL.n37 VTAIL.n35 24.41
R249 VTAIL.n133 VTAIL.n103 20.8927
R250 VTAIL.n130 VTAIL.n104 12.0247
R251 VTAIL.n28 VTAIL.n2 12.0247
R252 VTAIL.n100 VTAIL.n74 12.0247
R253 VTAIL.n66 VTAIL.n40 12.0247
R254 VTAIL.n129 VTAIL.n106 11.249
R255 VTAIL.n27 VTAIL.n4 11.249
R256 VTAIL.n99 VTAIL.n76 11.249
R257 VTAIL.n65 VTAIL.n42 11.249
R258 VTAIL.n114 VTAIL.n113 10.722
R259 VTAIL.n12 VTAIL.n11 10.722
R260 VTAIL.n84 VTAIL.n83 10.722
R261 VTAIL.n50 VTAIL.n49 10.722
R262 VTAIL.n126 VTAIL.n125 10.4732
R263 VTAIL.n24 VTAIL.n23 10.4732
R264 VTAIL.n96 VTAIL.n95 10.4732
R265 VTAIL.n62 VTAIL.n61 10.4732
R266 VTAIL.n122 VTAIL.n108 9.69747
R267 VTAIL.n20 VTAIL.n6 9.69747
R268 VTAIL.n92 VTAIL.n78 9.69747
R269 VTAIL.n58 VTAIL.n44 9.69747
R270 VTAIL.n128 VTAIL.n104 9.45567
R271 VTAIL.n26 VTAIL.n2 9.45567
R272 VTAIL.n98 VTAIL.n74 9.45567
R273 VTAIL.n64 VTAIL.n40 9.45567
R274 VTAIL.n112 VTAIL.n111 9.3005
R275 VTAIL.n119 VTAIL.n118 9.3005
R276 VTAIL.n121 VTAIL.n120 9.3005
R277 VTAIL.n108 VTAIL.n107 9.3005
R278 VTAIL.n127 VTAIL.n126 9.3005
R279 VTAIL.n129 VTAIL.n128 9.3005
R280 VTAIL.n10 VTAIL.n9 9.3005
R281 VTAIL.n17 VTAIL.n16 9.3005
R282 VTAIL.n19 VTAIL.n18 9.3005
R283 VTAIL.n6 VTAIL.n5 9.3005
R284 VTAIL.n25 VTAIL.n24 9.3005
R285 VTAIL.n27 VTAIL.n26 9.3005
R286 VTAIL.n99 VTAIL.n98 9.3005
R287 VTAIL.n97 VTAIL.n96 9.3005
R288 VTAIL.n78 VTAIL.n77 9.3005
R289 VTAIL.n91 VTAIL.n90 9.3005
R290 VTAIL.n89 VTAIL.n88 9.3005
R291 VTAIL.n82 VTAIL.n81 9.3005
R292 VTAIL.n55 VTAIL.n54 9.3005
R293 VTAIL.n57 VTAIL.n56 9.3005
R294 VTAIL.n44 VTAIL.n43 9.3005
R295 VTAIL.n63 VTAIL.n62 9.3005
R296 VTAIL.n65 VTAIL.n64 9.3005
R297 VTAIL.n48 VTAIL.n47 9.3005
R298 VTAIL.n121 VTAIL.n110 8.92171
R299 VTAIL.n19 VTAIL.n8 8.92171
R300 VTAIL.n91 VTAIL.n80 8.92171
R301 VTAIL.n57 VTAIL.n46 8.92171
R302 VTAIL.n118 VTAIL.n117 8.14595
R303 VTAIL.n16 VTAIL.n15 8.14595
R304 VTAIL.n88 VTAIL.n87 8.14595
R305 VTAIL.n54 VTAIL.n53 8.14595
R306 VTAIL.n114 VTAIL.n112 7.3702
R307 VTAIL.n12 VTAIL.n10 7.3702
R308 VTAIL.n84 VTAIL.n82 7.3702
R309 VTAIL.n50 VTAIL.n48 7.3702
R310 VTAIL.n117 VTAIL.n112 5.81868
R311 VTAIL.n15 VTAIL.n10 5.81868
R312 VTAIL.n87 VTAIL.n82 5.81868
R313 VTAIL.n53 VTAIL.n48 5.81868
R314 VTAIL.n134 VTAIL.t17 5.59516
R315 VTAIL.n134 VTAIL.t16 5.59516
R316 VTAIL.n0 VTAIL.t10 5.59516
R317 VTAIL.n0 VTAIL.t11 5.59516
R318 VTAIL.n32 VTAIL.t7 5.59516
R319 VTAIL.n32 VTAIL.t9 5.59516
R320 VTAIL.n34 VTAIL.t1 5.59516
R321 VTAIL.n34 VTAIL.t6 5.59516
R322 VTAIL.n72 VTAIL.t3 5.59516
R323 VTAIL.n72 VTAIL.t8 5.59516
R324 VTAIL.n70 VTAIL.t0 5.59516
R325 VTAIL.n70 VTAIL.t5 5.59516
R326 VTAIL.n38 VTAIL.t19 5.59516
R327 VTAIL.n38 VTAIL.t15 5.59516
R328 VTAIL.n36 VTAIL.t12 5.59516
R329 VTAIL.n36 VTAIL.t14 5.59516
R330 VTAIL.n118 VTAIL.n110 5.04292
R331 VTAIL.n16 VTAIL.n8 5.04292
R332 VTAIL.n88 VTAIL.n80 5.04292
R333 VTAIL.n54 VTAIL.n46 5.04292
R334 VTAIL.n122 VTAIL.n121 4.26717
R335 VTAIL.n20 VTAIL.n19 4.26717
R336 VTAIL.n92 VTAIL.n91 4.26717
R337 VTAIL.n58 VTAIL.n57 4.26717
R338 VTAIL.n39 VTAIL.n37 3.51774
R339 VTAIL.n69 VTAIL.n39 3.51774
R340 VTAIL.n73 VTAIL.n71 3.51774
R341 VTAIL.n103 VTAIL.n73 3.51774
R342 VTAIL.n35 VTAIL.n33 3.51774
R343 VTAIL.n33 VTAIL.n31 3.51774
R344 VTAIL.n135 VTAIL.n133 3.51774
R345 VTAIL.n125 VTAIL.n108 3.49141
R346 VTAIL.n23 VTAIL.n6 3.49141
R347 VTAIL.n95 VTAIL.n78 3.49141
R348 VTAIL.n61 VTAIL.n44 3.49141
R349 VTAIL.n126 VTAIL.n106 2.71565
R350 VTAIL.n24 VTAIL.n4 2.71565
R351 VTAIL.n96 VTAIL.n76 2.71565
R352 VTAIL.n62 VTAIL.n42 2.71565
R353 VTAIL VTAIL.n1 2.69662
R354 VTAIL.n113 VTAIL.n111 2.4147
R355 VTAIL.n11 VTAIL.n9 2.4147
R356 VTAIL.n83 VTAIL.n81 2.4147
R357 VTAIL.n49 VTAIL.n47 2.4147
R358 VTAIL.n71 VTAIL.n69 2.22895
R359 VTAIL.n31 VTAIL.n1 2.22895
R360 VTAIL.n130 VTAIL.n129 1.93989
R361 VTAIL.n28 VTAIL.n27 1.93989
R362 VTAIL.n100 VTAIL.n99 1.93989
R363 VTAIL.n66 VTAIL.n65 1.93989
R364 VTAIL.n132 VTAIL.n104 1.16414
R365 VTAIL.n30 VTAIL.n2 1.16414
R366 VTAIL.n102 VTAIL.n74 1.16414
R367 VTAIL.n68 VTAIL.n40 1.16414
R368 VTAIL VTAIL.n135 0.821621
R369 VTAIL.n119 VTAIL.n111 0.155672
R370 VTAIL.n120 VTAIL.n119 0.155672
R371 VTAIL.n120 VTAIL.n107 0.155672
R372 VTAIL.n127 VTAIL.n107 0.155672
R373 VTAIL.n128 VTAIL.n127 0.155672
R374 VTAIL.n17 VTAIL.n9 0.155672
R375 VTAIL.n18 VTAIL.n17 0.155672
R376 VTAIL.n18 VTAIL.n5 0.155672
R377 VTAIL.n25 VTAIL.n5 0.155672
R378 VTAIL.n26 VTAIL.n25 0.155672
R379 VTAIL.n98 VTAIL.n97 0.155672
R380 VTAIL.n97 VTAIL.n77 0.155672
R381 VTAIL.n90 VTAIL.n77 0.155672
R382 VTAIL.n90 VTAIL.n89 0.155672
R383 VTAIL.n89 VTAIL.n81 0.155672
R384 VTAIL.n64 VTAIL.n63 0.155672
R385 VTAIL.n63 VTAIL.n43 0.155672
R386 VTAIL.n56 VTAIL.n43 0.155672
R387 VTAIL.n56 VTAIL.n55 0.155672
R388 VTAIL.n55 VTAIL.n47 0.155672
R389 VDD2.n61 VDD2.n60 756.745
R390 VDD2.n28 VDD2.n27 756.745
R391 VDD2.n60 VDD2.n59 585
R392 VDD2.n35 VDD2.n34 585
R393 VDD2.n54 VDD2.n53 585
R394 VDD2.n52 VDD2.n51 585
R395 VDD2.n39 VDD2.n38 585
R396 VDD2.n46 VDD2.n45 585
R397 VDD2.n44 VDD2.n43 585
R398 VDD2.n11 VDD2.n10 585
R399 VDD2.n13 VDD2.n12 585
R400 VDD2.n6 VDD2.n5 585
R401 VDD2.n19 VDD2.n18 585
R402 VDD2.n21 VDD2.n20 585
R403 VDD2.n2 VDD2.n1 585
R404 VDD2.n27 VDD2.n26 585
R405 VDD2.n9 VDD2.t2 329.175
R406 VDD2.n42 VDD2.t0 329.175
R407 VDD2.n60 VDD2.n34 171.744
R408 VDD2.n53 VDD2.n34 171.744
R409 VDD2.n53 VDD2.n52 171.744
R410 VDD2.n52 VDD2.n38 171.744
R411 VDD2.n45 VDD2.n38 171.744
R412 VDD2.n45 VDD2.n44 171.744
R413 VDD2.n12 VDD2.n11 171.744
R414 VDD2.n12 VDD2.n5 171.744
R415 VDD2.n19 VDD2.n5 171.744
R416 VDD2.n20 VDD2.n19 171.744
R417 VDD2.n20 VDD2.n1 171.744
R418 VDD2.n27 VDD2.n1 171.744
R419 VDD2.n32 VDD2.n31 97.5006
R420 VDD2 VDD2.n65 97.4976
R421 VDD2.n64 VDD2.n63 94.919
R422 VDD2.n30 VDD2.n29 94.918
R423 VDD2.n44 VDD2.t0 85.8723
R424 VDD2.n11 VDD2.t2 85.8723
R425 VDD2.n30 VDD2.n28 54.5147
R426 VDD2.n62 VDD2.n61 50.9975
R427 VDD2.n62 VDD2.n32 45.4308
R428 VDD2.n59 VDD2.n33 12.0247
R429 VDD2.n26 VDD2.n0 12.0247
R430 VDD2.n58 VDD2.n35 11.249
R431 VDD2.n25 VDD2.n2 11.249
R432 VDD2.n10 VDD2.n9 10.722
R433 VDD2.n43 VDD2.n42 10.722
R434 VDD2.n55 VDD2.n54 10.4732
R435 VDD2.n22 VDD2.n21 10.4732
R436 VDD2.n51 VDD2.n37 9.69747
R437 VDD2.n18 VDD2.n4 9.69747
R438 VDD2.n57 VDD2.n33 9.45567
R439 VDD2.n24 VDD2.n0 9.45567
R440 VDD2.n48 VDD2.n47 9.3005
R441 VDD2.n50 VDD2.n49 9.3005
R442 VDD2.n37 VDD2.n36 9.3005
R443 VDD2.n56 VDD2.n55 9.3005
R444 VDD2.n58 VDD2.n57 9.3005
R445 VDD2.n41 VDD2.n40 9.3005
R446 VDD2.n8 VDD2.n7 9.3005
R447 VDD2.n15 VDD2.n14 9.3005
R448 VDD2.n17 VDD2.n16 9.3005
R449 VDD2.n4 VDD2.n3 9.3005
R450 VDD2.n23 VDD2.n22 9.3005
R451 VDD2.n25 VDD2.n24 9.3005
R452 VDD2.n50 VDD2.n39 8.92171
R453 VDD2.n17 VDD2.n6 8.92171
R454 VDD2.n47 VDD2.n46 8.14595
R455 VDD2.n14 VDD2.n13 8.14595
R456 VDD2.n43 VDD2.n41 7.3702
R457 VDD2.n10 VDD2.n8 7.3702
R458 VDD2.n46 VDD2.n41 5.81868
R459 VDD2.n13 VDD2.n8 5.81868
R460 VDD2.n65 VDD2.t1 5.59516
R461 VDD2.n65 VDD2.t4 5.59516
R462 VDD2.n63 VDD2.t3 5.59516
R463 VDD2.n63 VDD2.t5 5.59516
R464 VDD2.n31 VDD2.t7 5.59516
R465 VDD2.n31 VDD2.t9 5.59516
R466 VDD2.n29 VDD2.t6 5.59516
R467 VDD2.n29 VDD2.t8 5.59516
R468 VDD2.n47 VDD2.n39 5.04292
R469 VDD2.n14 VDD2.n6 5.04292
R470 VDD2.n51 VDD2.n50 4.26717
R471 VDD2.n18 VDD2.n17 4.26717
R472 VDD2.n64 VDD2.n62 3.51774
R473 VDD2.n54 VDD2.n37 3.49141
R474 VDD2.n21 VDD2.n4 3.49141
R475 VDD2.n55 VDD2.n35 2.71565
R476 VDD2.n22 VDD2.n2 2.71565
R477 VDD2.n9 VDD2.n7 2.4147
R478 VDD2.n42 VDD2.n40 2.4147
R479 VDD2.n59 VDD2.n58 1.93989
R480 VDD2.n26 VDD2.n25 1.93989
R481 VDD2.n61 VDD2.n33 1.16414
R482 VDD2.n28 VDD2.n0 1.16414
R483 VDD2 VDD2.n64 0.938
R484 VDD2.n32 VDD2.n30 0.824464
R485 VDD2.n57 VDD2.n56 0.155672
R486 VDD2.n56 VDD2.n36 0.155672
R487 VDD2.n49 VDD2.n36 0.155672
R488 VDD2.n49 VDD2.n48 0.155672
R489 VDD2.n48 VDD2.n40 0.155672
R490 VDD2.n15 VDD2.n7 0.155672
R491 VDD2.n16 VDD2.n15 0.155672
R492 VDD2.n16 VDD2.n3 0.155672
R493 VDD2.n23 VDD2.n3 0.155672
R494 VDD2.n24 VDD2.n23 0.155672
R495 B.n674 B.n673 585
R496 B.n675 B.n74 585
R497 B.n677 B.n676 585
R498 B.n678 B.n73 585
R499 B.n680 B.n679 585
R500 B.n681 B.n72 585
R501 B.n683 B.n682 585
R502 B.n684 B.n71 585
R503 B.n686 B.n685 585
R504 B.n687 B.n70 585
R505 B.n689 B.n688 585
R506 B.n690 B.n69 585
R507 B.n692 B.n691 585
R508 B.n693 B.n68 585
R509 B.n695 B.n694 585
R510 B.n696 B.n67 585
R511 B.n698 B.n697 585
R512 B.n699 B.n66 585
R513 B.n701 B.n700 585
R514 B.n702 B.n65 585
R515 B.n704 B.n703 585
R516 B.n705 B.n61 585
R517 B.n707 B.n706 585
R518 B.n708 B.n60 585
R519 B.n710 B.n709 585
R520 B.n711 B.n59 585
R521 B.n713 B.n712 585
R522 B.n714 B.n58 585
R523 B.n716 B.n715 585
R524 B.n717 B.n57 585
R525 B.n719 B.n718 585
R526 B.n720 B.n56 585
R527 B.n722 B.n721 585
R528 B.n724 B.n53 585
R529 B.n726 B.n725 585
R530 B.n727 B.n52 585
R531 B.n729 B.n728 585
R532 B.n730 B.n51 585
R533 B.n732 B.n731 585
R534 B.n733 B.n50 585
R535 B.n735 B.n734 585
R536 B.n736 B.n49 585
R537 B.n738 B.n737 585
R538 B.n739 B.n48 585
R539 B.n741 B.n740 585
R540 B.n742 B.n47 585
R541 B.n744 B.n743 585
R542 B.n745 B.n46 585
R543 B.n747 B.n746 585
R544 B.n748 B.n45 585
R545 B.n750 B.n749 585
R546 B.n751 B.n44 585
R547 B.n753 B.n752 585
R548 B.n754 B.n43 585
R549 B.n756 B.n755 585
R550 B.n757 B.n42 585
R551 B.n672 B.n75 585
R552 B.n671 B.n670 585
R553 B.n669 B.n76 585
R554 B.n668 B.n667 585
R555 B.n666 B.n77 585
R556 B.n665 B.n664 585
R557 B.n663 B.n78 585
R558 B.n662 B.n661 585
R559 B.n660 B.n79 585
R560 B.n659 B.n658 585
R561 B.n657 B.n80 585
R562 B.n656 B.n655 585
R563 B.n654 B.n81 585
R564 B.n653 B.n652 585
R565 B.n651 B.n82 585
R566 B.n650 B.n649 585
R567 B.n648 B.n83 585
R568 B.n647 B.n646 585
R569 B.n645 B.n84 585
R570 B.n644 B.n643 585
R571 B.n642 B.n85 585
R572 B.n641 B.n640 585
R573 B.n639 B.n86 585
R574 B.n638 B.n637 585
R575 B.n636 B.n87 585
R576 B.n635 B.n634 585
R577 B.n633 B.n88 585
R578 B.n632 B.n631 585
R579 B.n630 B.n89 585
R580 B.n629 B.n628 585
R581 B.n627 B.n90 585
R582 B.n626 B.n625 585
R583 B.n624 B.n91 585
R584 B.n623 B.n622 585
R585 B.n621 B.n92 585
R586 B.n620 B.n619 585
R587 B.n618 B.n93 585
R588 B.n617 B.n616 585
R589 B.n615 B.n94 585
R590 B.n614 B.n613 585
R591 B.n612 B.n95 585
R592 B.n611 B.n610 585
R593 B.n609 B.n96 585
R594 B.n608 B.n607 585
R595 B.n606 B.n97 585
R596 B.n605 B.n604 585
R597 B.n603 B.n98 585
R598 B.n602 B.n601 585
R599 B.n600 B.n99 585
R600 B.n599 B.n598 585
R601 B.n597 B.n100 585
R602 B.n596 B.n595 585
R603 B.n594 B.n101 585
R604 B.n593 B.n592 585
R605 B.n591 B.n102 585
R606 B.n590 B.n589 585
R607 B.n588 B.n103 585
R608 B.n587 B.n586 585
R609 B.n585 B.n104 585
R610 B.n584 B.n583 585
R611 B.n582 B.n105 585
R612 B.n581 B.n580 585
R613 B.n579 B.n106 585
R614 B.n578 B.n577 585
R615 B.n576 B.n107 585
R616 B.n575 B.n574 585
R617 B.n573 B.n108 585
R618 B.n572 B.n571 585
R619 B.n570 B.n109 585
R620 B.n569 B.n568 585
R621 B.n567 B.n110 585
R622 B.n566 B.n565 585
R623 B.n564 B.n111 585
R624 B.n563 B.n562 585
R625 B.n561 B.n112 585
R626 B.n560 B.n559 585
R627 B.n558 B.n113 585
R628 B.n557 B.n556 585
R629 B.n555 B.n114 585
R630 B.n554 B.n553 585
R631 B.n552 B.n115 585
R632 B.n551 B.n550 585
R633 B.n549 B.n116 585
R634 B.n548 B.n547 585
R635 B.n546 B.n117 585
R636 B.n545 B.n544 585
R637 B.n543 B.n118 585
R638 B.n542 B.n541 585
R639 B.n540 B.n119 585
R640 B.n539 B.n538 585
R641 B.n537 B.n120 585
R642 B.n536 B.n535 585
R643 B.n534 B.n121 585
R644 B.n533 B.n532 585
R645 B.n531 B.n122 585
R646 B.n530 B.n529 585
R647 B.n528 B.n123 585
R648 B.n527 B.n526 585
R649 B.n525 B.n124 585
R650 B.n524 B.n523 585
R651 B.n522 B.n125 585
R652 B.n521 B.n520 585
R653 B.n519 B.n126 585
R654 B.n518 B.n517 585
R655 B.n516 B.n127 585
R656 B.n515 B.n514 585
R657 B.n513 B.n128 585
R658 B.n512 B.n511 585
R659 B.n510 B.n129 585
R660 B.n509 B.n508 585
R661 B.n507 B.n130 585
R662 B.n506 B.n505 585
R663 B.n504 B.n131 585
R664 B.n503 B.n502 585
R665 B.n501 B.n132 585
R666 B.n500 B.n499 585
R667 B.n498 B.n133 585
R668 B.n497 B.n496 585
R669 B.n495 B.n134 585
R670 B.n494 B.n493 585
R671 B.n492 B.n135 585
R672 B.n491 B.n490 585
R673 B.n489 B.n136 585
R674 B.n488 B.n487 585
R675 B.n486 B.n137 585
R676 B.n485 B.n484 585
R677 B.n483 B.n138 585
R678 B.n482 B.n481 585
R679 B.n480 B.n139 585
R680 B.n479 B.n478 585
R681 B.n477 B.n140 585
R682 B.n476 B.n475 585
R683 B.n474 B.n141 585
R684 B.n473 B.n472 585
R685 B.n471 B.n142 585
R686 B.n470 B.n469 585
R687 B.n468 B.n143 585
R688 B.n467 B.n466 585
R689 B.n465 B.n144 585
R690 B.n464 B.n463 585
R691 B.n462 B.n145 585
R692 B.n461 B.n460 585
R693 B.n459 B.n146 585
R694 B.n458 B.n457 585
R695 B.n456 B.n147 585
R696 B.n455 B.n454 585
R697 B.n453 B.n148 585
R698 B.n452 B.n451 585
R699 B.n450 B.n149 585
R700 B.n449 B.n448 585
R701 B.n447 B.n150 585
R702 B.n446 B.n445 585
R703 B.n444 B.n151 585
R704 B.n443 B.n442 585
R705 B.n441 B.n152 585
R706 B.n440 B.n439 585
R707 B.n438 B.n153 585
R708 B.n437 B.n436 585
R709 B.n435 B.n154 585
R710 B.n434 B.n433 585
R711 B.n432 B.n155 585
R712 B.n347 B.n346 585
R713 B.n348 B.n187 585
R714 B.n350 B.n349 585
R715 B.n351 B.n186 585
R716 B.n353 B.n352 585
R717 B.n354 B.n185 585
R718 B.n356 B.n355 585
R719 B.n357 B.n184 585
R720 B.n359 B.n358 585
R721 B.n360 B.n183 585
R722 B.n362 B.n361 585
R723 B.n363 B.n182 585
R724 B.n365 B.n364 585
R725 B.n366 B.n181 585
R726 B.n368 B.n367 585
R727 B.n369 B.n180 585
R728 B.n371 B.n370 585
R729 B.n372 B.n179 585
R730 B.n374 B.n373 585
R731 B.n375 B.n178 585
R732 B.n377 B.n376 585
R733 B.n378 B.n177 585
R734 B.n380 B.n379 585
R735 B.n382 B.n174 585
R736 B.n384 B.n383 585
R737 B.n385 B.n173 585
R738 B.n387 B.n386 585
R739 B.n388 B.n172 585
R740 B.n390 B.n389 585
R741 B.n391 B.n171 585
R742 B.n393 B.n392 585
R743 B.n394 B.n170 585
R744 B.n396 B.n395 585
R745 B.n398 B.n397 585
R746 B.n399 B.n166 585
R747 B.n401 B.n400 585
R748 B.n402 B.n165 585
R749 B.n404 B.n403 585
R750 B.n405 B.n164 585
R751 B.n407 B.n406 585
R752 B.n408 B.n163 585
R753 B.n410 B.n409 585
R754 B.n411 B.n162 585
R755 B.n413 B.n412 585
R756 B.n414 B.n161 585
R757 B.n416 B.n415 585
R758 B.n417 B.n160 585
R759 B.n419 B.n418 585
R760 B.n420 B.n159 585
R761 B.n422 B.n421 585
R762 B.n423 B.n158 585
R763 B.n425 B.n424 585
R764 B.n426 B.n157 585
R765 B.n428 B.n427 585
R766 B.n429 B.n156 585
R767 B.n431 B.n430 585
R768 B.n345 B.n188 585
R769 B.n344 B.n343 585
R770 B.n342 B.n189 585
R771 B.n341 B.n340 585
R772 B.n339 B.n190 585
R773 B.n338 B.n337 585
R774 B.n336 B.n191 585
R775 B.n335 B.n334 585
R776 B.n333 B.n192 585
R777 B.n332 B.n331 585
R778 B.n330 B.n193 585
R779 B.n329 B.n328 585
R780 B.n327 B.n194 585
R781 B.n326 B.n325 585
R782 B.n324 B.n195 585
R783 B.n323 B.n322 585
R784 B.n321 B.n196 585
R785 B.n320 B.n319 585
R786 B.n318 B.n197 585
R787 B.n317 B.n316 585
R788 B.n315 B.n198 585
R789 B.n314 B.n313 585
R790 B.n312 B.n199 585
R791 B.n311 B.n310 585
R792 B.n309 B.n200 585
R793 B.n308 B.n307 585
R794 B.n306 B.n201 585
R795 B.n305 B.n304 585
R796 B.n303 B.n202 585
R797 B.n302 B.n301 585
R798 B.n300 B.n203 585
R799 B.n299 B.n298 585
R800 B.n297 B.n204 585
R801 B.n296 B.n295 585
R802 B.n294 B.n205 585
R803 B.n293 B.n292 585
R804 B.n291 B.n206 585
R805 B.n290 B.n289 585
R806 B.n288 B.n207 585
R807 B.n287 B.n286 585
R808 B.n285 B.n208 585
R809 B.n284 B.n283 585
R810 B.n282 B.n209 585
R811 B.n281 B.n280 585
R812 B.n279 B.n210 585
R813 B.n278 B.n277 585
R814 B.n276 B.n211 585
R815 B.n275 B.n274 585
R816 B.n273 B.n212 585
R817 B.n272 B.n271 585
R818 B.n270 B.n213 585
R819 B.n269 B.n268 585
R820 B.n267 B.n214 585
R821 B.n266 B.n265 585
R822 B.n264 B.n215 585
R823 B.n263 B.n262 585
R824 B.n261 B.n216 585
R825 B.n260 B.n259 585
R826 B.n258 B.n217 585
R827 B.n257 B.n256 585
R828 B.n255 B.n218 585
R829 B.n254 B.n253 585
R830 B.n252 B.n219 585
R831 B.n251 B.n250 585
R832 B.n249 B.n220 585
R833 B.n248 B.n247 585
R834 B.n246 B.n221 585
R835 B.n245 B.n244 585
R836 B.n243 B.n222 585
R837 B.n242 B.n241 585
R838 B.n240 B.n223 585
R839 B.n239 B.n238 585
R840 B.n237 B.n224 585
R841 B.n236 B.n235 585
R842 B.n234 B.n225 585
R843 B.n233 B.n232 585
R844 B.n231 B.n226 585
R845 B.n230 B.n229 585
R846 B.n228 B.n227 585
R847 B.n2 B.n0 585
R848 B.n877 B.n1 585
R849 B.n876 B.n875 585
R850 B.n874 B.n3 585
R851 B.n873 B.n872 585
R852 B.n871 B.n4 585
R853 B.n870 B.n869 585
R854 B.n868 B.n5 585
R855 B.n867 B.n866 585
R856 B.n865 B.n6 585
R857 B.n864 B.n863 585
R858 B.n862 B.n7 585
R859 B.n861 B.n860 585
R860 B.n859 B.n8 585
R861 B.n858 B.n857 585
R862 B.n856 B.n9 585
R863 B.n855 B.n854 585
R864 B.n853 B.n10 585
R865 B.n852 B.n851 585
R866 B.n850 B.n11 585
R867 B.n849 B.n848 585
R868 B.n847 B.n12 585
R869 B.n846 B.n845 585
R870 B.n844 B.n13 585
R871 B.n843 B.n842 585
R872 B.n841 B.n14 585
R873 B.n840 B.n839 585
R874 B.n838 B.n15 585
R875 B.n837 B.n836 585
R876 B.n835 B.n16 585
R877 B.n834 B.n833 585
R878 B.n832 B.n17 585
R879 B.n831 B.n830 585
R880 B.n829 B.n18 585
R881 B.n828 B.n827 585
R882 B.n826 B.n19 585
R883 B.n825 B.n824 585
R884 B.n823 B.n20 585
R885 B.n822 B.n821 585
R886 B.n820 B.n21 585
R887 B.n819 B.n818 585
R888 B.n817 B.n22 585
R889 B.n816 B.n815 585
R890 B.n814 B.n23 585
R891 B.n813 B.n812 585
R892 B.n811 B.n24 585
R893 B.n810 B.n809 585
R894 B.n808 B.n25 585
R895 B.n807 B.n806 585
R896 B.n805 B.n26 585
R897 B.n804 B.n803 585
R898 B.n802 B.n27 585
R899 B.n801 B.n800 585
R900 B.n799 B.n28 585
R901 B.n798 B.n797 585
R902 B.n796 B.n29 585
R903 B.n795 B.n794 585
R904 B.n793 B.n30 585
R905 B.n792 B.n791 585
R906 B.n790 B.n31 585
R907 B.n789 B.n788 585
R908 B.n787 B.n32 585
R909 B.n786 B.n785 585
R910 B.n784 B.n33 585
R911 B.n783 B.n782 585
R912 B.n781 B.n34 585
R913 B.n780 B.n779 585
R914 B.n778 B.n35 585
R915 B.n777 B.n776 585
R916 B.n775 B.n36 585
R917 B.n774 B.n773 585
R918 B.n772 B.n37 585
R919 B.n771 B.n770 585
R920 B.n769 B.n38 585
R921 B.n768 B.n767 585
R922 B.n766 B.n39 585
R923 B.n765 B.n764 585
R924 B.n763 B.n40 585
R925 B.n762 B.n761 585
R926 B.n760 B.n41 585
R927 B.n759 B.n758 585
R928 B.n879 B.n878 585
R929 B.n347 B.n188 550.159
R930 B.n758 B.n757 550.159
R931 B.n432 B.n431 550.159
R932 B.n673 B.n672 550.159
R933 B.n167 B.t8 343.635
R934 B.n62 B.t10 343.635
R935 B.n175 B.t5 343.635
R936 B.n54 B.t1 343.635
R937 B.n168 B.t7 264.509
R938 B.n63 B.t11 264.509
R939 B.n176 B.t4 264.509
R940 B.n55 B.t2 264.509
R941 B.n167 B.t6 246.643
R942 B.n175 B.t3 246.643
R943 B.n54 B.t0 246.643
R944 B.n62 B.t9 246.643
R945 B.n343 B.n188 163.367
R946 B.n343 B.n342 163.367
R947 B.n342 B.n341 163.367
R948 B.n341 B.n190 163.367
R949 B.n337 B.n190 163.367
R950 B.n337 B.n336 163.367
R951 B.n336 B.n335 163.367
R952 B.n335 B.n192 163.367
R953 B.n331 B.n192 163.367
R954 B.n331 B.n330 163.367
R955 B.n330 B.n329 163.367
R956 B.n329 B.n194 163.367
R957 B.n325 B.n194 163.367
R958 B.n325 B.n324 163.367
R959 B.n324 B.n323 163.367
R960 B.n323 B.n196 163.367
R961 B.n319 B.n196 163.367
R962 B.n319 B.n318 163.367
R963 B.n318 B.n317 163.367
R964 B.n317 B.n198 163.367
R965 B.n313 B.n198 163.367
R966 B.n313 B.n312 163.367
R967 B.n312 B.n311 163.367
R968 B.n311 B.n200 163.367
R969 B.n307 B.n200 163.367
R970 B.n307 B.n306 163.367
R971 B.n306 B.n305 163.367
R972 B.n305 B.n202 163.367
R973 B.n301 B.n202 163.367
R974 B.n301 B.n300 163.367
R975 B.n300 B.n299 163.367
R976 B.n299 B.n204 163.367
R977 B.n295 B.n204 163.367
R978 B.n295 B.n294 163.367
R979 B.n294 B.n293 163.367
R980 B.n293 B.n206 163.367
R981 B.n289 B.n206 163.367
R982 B.n289 B.n288 163.367
R983 B.n288 B.n287 163.367
R984 B.n287 B.n208 163.367
R985 B.n283 B.n208 163.367
R986 B.n283 B.n282 163.367
R987 B.n282 B.n281 163.367
R988 B.n281 B.n210 163.367
R989 B.n277 B.n210 163.367
R990 B.n277 B.n276 163.367
R991 B.n276 B.n275 163.367
R992 B.n275 B.n212 163.367
R993 B.n271 B.n212 163.367
R994 B.n271 B.n270 163.367
R995 B.n270 B.n269 163.367
R996 B.n269 B.n214 163.367
R997 B.n265 B.n214 163.367
R998 B.n265 B.n264 163.367
R999 B.n264 B.n263 163.367
R1000 B.n263 B.n216 163.367
R1001 B.n259 B.n216 163.367
R1002 B.n259 B.n258 163.367
R1003 B.n258 B.n257 163.367
R1004 B.n257 B.n218 163.367
R1005 B.n253 B.n218 163.367
R1006 B.n253 B.n252 163.367
R1007 B.n252 B.n251 163.367
R1008 B.n251 B.n220 163.367
R1009 B.n247 B.n220 163.367
R1010 B.n247 B.n246 163.367
R1011 B.n246 B.n245 163.367
R1012 B.n245 B.n222 163.367
R1013 B.n241 B.n222 163.367
R1014 B.n241 B.n240 163.367
R1015 B.n240 B.n239 163.367
R1016 B.n239 B.n224 163.367
R1017 B.n235 B.n224 163.367
R1018 B.n235 B.n234 163.367
R1019 B.n234 B.n233 163.367
R1020 B.n233 B.n226 163.367
R1021 B.n229 B.n226 163.367
R1022 B.n229 B.n228 163.367
R1023 B.n228 B.n2 163.367
R1024 B.n878 B.n2 163.367
R1025 B.n878 B.n877 163.367
R1026 B.n877 B.n876 163.367
R1027 B.n876 B.n3 163.367
R1028 B.n872 B.n3 163.367
R1029 B.n872 B.n871 163.367
R1030 B.n871 B.n870 163.367
R1031 B.n870 B.n5 163.367
R1032 B.n866 B.n5 163.367
R1033 B.n866 B.n865 163.367
R1034 B.n865 B.n864 163.367
R1035 B.n864 B.n7 163.367
R1036 B.n860 B.n7 163.367
R1037 B.n860 B.n859 163.367
R1038 B.n859 B.n858 163.367
R1039 B.n858 B.n9 163.367
R1040 B.n854 B.n9 163.367
R1041 B.n854 B.n853 163.367
R1042 B.n853 B.n852 163.367
R1043 B.n852 B.n11 163.367
R1044 B.n848 B.n11 163.367
R1045 B.n848 B.n847 163.367
R1046 B.n847 B.n846 163.367
R1047 B.n846 B.n13 163.367
R1048 B.n842 B.n13 163.367
R1049 B.n842 B.n841 163.367
R1050 B.n841 B.n840 163.367
R1051 B.n840 B.n15 163.367
R1052 B.n836 B.n15 163.367
R1053 B.n836 B.n835 163.367
R1054 B.n835 B.n834 163.367
R1055 B.n834 B.n17 163.367
R1056 B.n830 B.n17 163.367
R1057 B.n830 B.n829 163.367
R1058 B.n829 B.n828 163.367
R1059 B.n828 B.n19 163.367
R1060 B.n824 B.n19 163.367
R1061 B.n824 B.n823 163.367
R1062 B.n823 B.n822 163.367
R1063 B.n822 B.n21 163.367
R1064 B.n818 B.n21 163.367
R1065 B.n818 B.n817 163.367
R1066 B.n817 B.n816 163.367
R1067 B.n816 B.n23 163.367
R1068 B.n812 B.n23 163.367
R1069 B.n812 B.n811 163.367
R1070 B.n811 B.n810 163.367
R1071 B.n810 B.n25 163.367
R1072 B.n806 B.n25 163.367
R1073 B.n806 B.n805 163.367
R1074 B.n805 B.n804 163.367
R1075 B.n804 B.n27 163.367
R1076 B.n800 B.n27 163.367
R1077 B.n800 B.n799 163.367
R1078 B.n799 B.n798 163.367
R1079 B.n798 B.n29 163.367
R1080 B.n794 B.n29 163.367
R1081 B.n794 B.n793 163.367
R1082 B.n793 B.n792 163.367
R1083 B.n792 B.n31 163.367
R1084 B.n788 B.n31 163.367
R1085 B.n788 B.n787 163.367
R1086 B.n787 B.n786 163.367
R1087 B.n786 B.n33 163.367
R1088 B.n782 B.n33 163.367
R1089 B.n782 B.n781 163.367
R1090 B.n781 B.n780 163.367
R1091 B.n780 B.n35 163.367
R1092 B.n776 B.n35 163.367
R1093 B.n776 B.n775 163.367
R1094 B.n775 B.n774 163.367
R1095 B.n774 B.n37 163.367
R1096 B.n770 B.n37 163.367
R1097 B.n770 B.n769 163.367
R1098 B.n769 B.n768 163.367
R1099 B.n768 B.n39 163.367
R1100 B.n764 B.n39 163.367
R1101 B.n764 B.n763 163.367
R1102 B.n763 B.n762 163.367
R1103 B.n762 B.n41 163.367
R1104 B.n758 B.n41 163.367
R1105 B.n348 B.n347 163.367
R1106 B.n349 B.n348 163.367
R1107 B.n349 B.n186 163.367
R1108 B.n353 B.n186 163.367
R1109 B.n354 B.n353 163.367
R1110 B.n355 B.n354 163.367
R1111 B.n355 B.n184 163.367
R1112 B.n359 B.n184 163.367
R1113 B.n360 B.n359 163.367
R1114 B.n361 B.n360 163.367
R1115 B.n361 B.n182 163.367
R1116 B.n365 B.n182 163.367
R1117 B.n366 B.n365 163.367
R1118 B.n367 B.n366 163.367
R1119 B.n367 B.n180 163.367
R1120 B.n371 B.n180 163.367
R1121 B.n372 B.n371 163.367
R1122 B.n373 B.n372 163.367
R1123 B.n373 B.n178 163.367
R1124 B.n377 B.n178 163.367
R1125 B.n378 B.n377 163.367
R1126 B.n379 B.n378 163.367
R1127 B.n379 B.n174 163.367
R1128 B.n384 B.n174 163.367
R1129 B.n385 B.n384 163.367
R1130 B.n386 B.n385 163.367
R1131 B.n386 B.n172 163.367
R1132 B.n390 B.n172 163.367
R1133 B.n391 B.n390 163.367
R1134 B.n392 B.n391 163.367
R1135 B.n392 B.n170 163.367
R1136 B.n396 B.n170 163.367
R1137 B.n397 B.n396 163.367
R1138 B.n397 B.n166 163.367
R1139 B.n401 B.n166 163.367
R1140 B.n402 B.n401 163.367
R1141 B.n403 B.n402 163.367
R1142 B.n403 B.n164 163.367
R1143 B.n407 B.n164 163.367
R1144 B.n408 B.n407 163.367
R1145 B.n409 B.n408 163.367
R1146 B.n409 B.n162 163.367
R1147 B.n413 B.n162 163.367
R1148 B.n414 B.n413 163.367
R1149 B.n415 B.n414 163.367
R1150 B.n415 B.n160 163.367
R1151 B.n419 B.n160 163.367
R1152 B.n420 B.n419 163.367
R1153 B.n421 B.n420 163.367
R1154 B.n421 B.n158 163.367
R1155 B.n425 B.n158 163.367
R1156 B.n426 B.n425 163.367
R1157 B.n427 B.n426 163.367
R1158 B.n427 B.n156 163.367
R1159 B.n431 B.n156 163.367
R1160 B.n433 B.n432 163.367
R1161 B.n433 B.n154 163.367
R1162 B.n437 B.n154 163.367
R1163 B.n438 B.n437 163.367
R1164 B.n439 B.n438 163.367
R1165 B.n439 B.n152 163.367
R1166 B.n443 B.n152 163.367
R1167 B.n444 B.n443 163.367
R1168 B.n445 B.n444 163.367
R1169 B.n445 B.n150 163.367
R1170 B.n449 B.n150 163.367
R1171 B.n450 B.n449 163.367
R1172 B.n451 B.n450 163.367
R1173 B.n451 B.n148 163.367
R1174 B.n455 B.n148 163.367
R1175 B.n456 B.n455 163.367
R1176 B.n457 B.n456 163.367
R1177 B.n457 B.n146 163.367
R1178 B.n461 B.n146 163.367
R1179 B.n462 B.n461 163.367
R1180 B.n463 B.n462 163.367
R1181 B.n463 B.n144 163.367
R1182 B.n467 B.n144 163.367
R1183 B.n468 B.n467 163.367
R1184 B.n469 B.n468 163.367
R1185 B.n469 B.n142 163.367
R1186 B.n473 B.n142 163.367
R1187 B.n474 B.n473 163.367
R1188 B.n475 B.n474 163.367
R1189 B.n475 B.n140 163.367
R1190 B.n479 B.n140 163.367
R1191 B.n480 B.n479 163.367
R1192 B.n481 B.n480 163.367
R1193 B.n481 B.n138 163.367
R1194 B.n485 B.n138 163.367
R1195 B.n486 B.n485 163.367
R1196 B.n487 B.n486 163.367
R1197 B.n487 B.n136 163.367
R1198 B.n491 B.n136 163.367
R1199 B.n492 B.n491 163.367
R1200 B.n493 B.n492 163.367
R1201 B.n493 B.n134 163.367
R1202 B.n497 B.n134 163.367
R1203 B.n498 B.n497 163.367
R1204 B.n499 B.n498 163.367
R1205 B.n499 B.n132 163.367
R1206 B.n503 B.n132 163.367
R1207 B.n504 B.n503 163.367
R1208 B.n505 B.n504 163.367
R1209 B.n505 B.n130 163.367
R1210 B.n509 B.n130 163.367
R1211 B.n510 B.n509 163.367
R1212 B.n511 B.n510 163.367
R1213 B.n511 B.n128 163.367
R1214 B.n515 B.n128 163.367
R1215 B.n516 B.n515 163.367
R1216 B.n517 B.n516 163.367
R1217 B.n517 B.n126 163.367
R1218 B.n521 B.n126 163.367
R1219 B.n522 B.n521 163.367
R1220 B.n523 B.n522 163.367
R1221 B.n523 B.n124 163.367
R1222 B.n527 B.n124 163.367
R1223 B.n528 B.n527 163.367
R1224 B.n529 B.n528 163.367
R1225 B.n529 B.n122 163.367
R1226 B.n533 B.n122 163.367
R1227 B.n534 B.n533 163.367
R1228 B.n535 B.n534 163.367
R1229 B.n535 B.n120 163.367
R1230 B.n539 B.n120 163.367
R1231 B.n540 B.n539 163.367
R1232 B.n541 B.n540 163.367
R1233 B.n541 B.n118 163.367
R1234 B.n545 B.n118 163.367
R1235 B.n546 B.n545 163.367
R1236 B.n547 B.n546 163.367
R1237 B.n547 B.n116 163.367
R1238 B.n551 B.n116 163.367
R1239 B.n552 B.n551 163.367
R1240 B.n553 B.n552 163.367
R1241 B.n553 B.n114 163.367
R1242 B.n557 B.n114 163.367
R1243 B.n558 B.n557 163.367
R1244 B.n559 B.n558 163.367
R1245 B.n559 B.n112 163.367
R1246 B.n563 B.n112 163.367
R1247 B.n564 B.n563 163.367
R1248 B.n565 B.n564 163.367
R1249 B.n565 B.n110 163.367
R1250 B.n569 B.n110 163.367
R1251 B.n570 B.n569 163.367
R1252 B.n571 B.n570 163.367
R1253 B.n571 B.n108 163.367
R1254 B.n575 B.n108 163.367
R1255 B.n576 B.n575 163.367
R1256 B.n577 B.n576 163.367
R1257 B.n577 B.n106 163.367
R1258 B.n581 B.n106 163.367
R1259 B.n582 B.n581 163.367
R1260 B.n583 B.n582 163.367
R1261 B.n583 B.n104 163.367
R1262 B.n587 B.n104 163.367
R1263 B.n588 B.n587 163.367
R1264 B.n589 B.n588 163.367
R1265 B.n589 B.n102 163.367
R1266 B.n593 B.n102 163.367
R1267 B.n594 B.n593 163.367
R1268 B.n595 B.n594 163.367
R1269 B.n595 B.n100 163.367
R1270 B.n599 B.n100 163.367
R1271 B.n600 B.n599 163.367
R1272 B.n601 B.n600 163.367
R1273 B.n601 B.n98 163.367
R1274 B.n605 B.n98 163.367
R1275 B.n606 B.n605 163.367
R1276 B.n607 B.n606 163.367
R1277 B.n607 B.n96 163.367
R1278 B.n611 B.n96 163.367
R1279 B.n612 B.n611 163.367
R1280 B.n613 B.n612 163.367
R1281 B.n613 B.n94 163.367
R1282 B.n617 B.n94 163.367
R1283 B.n618 B.n617 163.367
R1284 B.n619 B.n618 163.367
R1285 B.n619 B.n92 163.367
R1286 B.n623 B.n92 163.367
R1287 B.n624 B.n623 163.367
R1288 B.n625 B.n624 163.367
R1289 B.n625 B.n90 163.367
R1290 B.n629 B.n90 163.367
R1291 B.n630 B.n629 163.367
R1292 B.n631 B.n630 163.367
R1293 B.n631 B.n88 163.367
R1294 B.n635 B.n88 163.367
R1295 B.n636 B.n635 163.367
R1296 B.n637 B.n636 163.367
R1297 B.n637 B.n86 163.367
R1298 B.n641 B.n86 163.367
R1299 B.n642 B.n641 163.367
R1300 B.n643 B.n642 163.367
R1301 B.n643 B.n84 163.367
R1302 B.n647 B.n84 163.367
R1303 B.n648 B.n647 163.367
R1304 B.n649 B.n648 163.367
R1305 B.n649 B.n82 163.367
R1306 B.n653 B.n82 163.367
R1307 B.n654 B.n653 163.367
R1308 B.n655 B.n654 163.367
R1309 B.n655 B.n80 163.367
R1310 B.n659 B.n80 163.367
R1311 B.n660 B.n659 163.367
R1312 B.n661 B.n660 163.367
R1313 B.n661 B.n78 163.367
R1314 B.n665 B.n78 163.367
R1315 B.n666 B.n665 163.367
R1316 B.n667 B.n666 163.367
R1317 B.n667 B.n76 163.367
R1318 B.n671 B.n76 163.367
R1319 B.n672 B.n671 163.367
R1320 B.n757 B.n756 163.367
R1321 B.n756 B.n43 163.367
R1322 B.n752 B.n43 163.367
R1323 B.n752 B.n751 163.367
R1324 B.n751 B.n750 163.367
R1325 B.n750 B.n45 163.367
R1326 B.n746 B.n45 163.367
R1327 B.n746 B.n745 163.367
R1328 B.n745 B.n744 163.367
R1329 B.n744 B.n47 163.367
R1330 B.n740 B.n47 163.367
R1331 B.n740 B.n739 163.367
R1332 B.n739 B.n738 163.367
R1333 B.n738 B.n49 163.367
R1334 B.n734 B.n49 163.367
R1335 B.n734 B.n733 163.367
R1336 B.n733 B.n732 163.367
R1337 B.n732 B.n51 163.367
R1338 B.n728 B.n51 163.367
R1339 B.n728 B.n727 163.367
R1340 B.n727 B.n726 163.367
R1341 B.n726 B.n53 163.367
R1342 B.n721 B.n53 163.367
R1343 B.n721 B.n720 163.367
R1344 B.n720 B.n719 163.367
R1345 B.n719 B.n57 163.367
R1346 B.n715 B.n57 163.367
R1347 B.n715 B.n714 163.367
R1348 B.n714 B.n713 163.367
R1349 B.n713 B.n59 163.367
R1350 B.n709 B.n59 163.367
R1351 B.n709 B.n708 163.367
R1352 B.n708 B.n707 163.367
R1353 B.n707 B.n61 163.367
R1354 B.n703 B.n61 163.367
R1355 B.n703 B.n702 163.367
R1356 B.n702 B.n701 163.367
R1357 B.n701 B.n66 163.367
R1358 B.n697 B.n66 163.367
R1359 B.n697 B.n696 163.367
R1360 B.n696 B.n695 163.367
R1361 B.n695 B.n68 163.367
R1362 B.n691 B.n68 163.367
R1363 B.n691 B.n690 163.367
R1364 B.n690 B.n689 163.367
R1365 B.n689 B.n70 163.367
R1366 B.n685 B.n70 163.367
R1367 B.n685 B.n684 163.367
R1368 B.n684 B.n683 163.367
R1369 B.n683 B.n72 163.367
R1370 B.n679 B.n72 163.367
R1371 B.n679 B.n678 163.367
R1372 B.n678 B.n677 163.367
R1373 B.n677 B.n74 163.367
R1374 B.n673 B.n74 163.367
R1375 B.n168 B.n167 79.1278
R1376 B.n176 B.n175 79.1278
R1377 B.n55 B.n54 79.1278
R1378 B.n63 B.n62 79.1278
R1379 B.n169 B.n168 59.5399
R1380 B.n381 B.n176 59.5399
R1381 B.n723 B.n55 59.5399
R1382 B.n64 B.n63 59.5399
R1383 B.n759 B.n42 35.7468
R1384 B.n430 B.n155 35.7468
R1385 B.n346 B.n345 35.7468
R1386 B.n674 B.n75 35.7468
R1387 B B.n879 18.0485
R1388 B.n755 B.n42 10.6151
R1389 B.n755 B.n754 10.6151
R1390 B.n754 B.n753 10.6151
R1391 B.n753 B.n44 10.6151
R1392 B.n749 B.n44 10.6151
R1393 B.n749 B.n748 10.6151
R1394 B.n748 B.n747 10.6151
R1395 B.n747 B.n46 10.6151
R1396 B.n743 B.n46 10.6151
R1397 B.n743 B.n742 10.6151
R1398 B.n742 B.n741 10.6151
R1399 B.n741 B.n48 10.6151
R1400 B.n737 B.n48 10.6151
R1401 B.n737 B.n736 10.6151
R1402 B.n736 B.n735 10.6151
R1403 B.n735 B.n50 10.6151
R1404 B.n731 B.n50 10.6151
R1405 B.n731 B.n730 10.6151
R1406 B.n730 B.n729 10.6151
R1407 B.n729 B.n52 10.6151
R1408 B.n725 B.n52 10.6151
R1409 B.n725 B.n724 10.6151
R1410 B.n722 B.n56 10.6151
R1411 B.n718 B.n56 10.6151
R1412 B.n718 B.n717 10.6151
R1413 B.n717 B.n716 10.6151
R1414 B.n716 B.n58 10.6151
R1415 B.n712 B.n58 10.6151
R1416 B.n712 B.n711 10.6151
R1417 B.n711 B.n710 10.6151
R1418 B.n710 B.n60 10.6151
R1419 B.n706 B.n705 10.6151
R1420 B.n705 B.n704 10.6151
R1421 B.n704 B.n65 10.6151
R1422 B.n700 B.n65 10.6151
R1423 B.n700 B.n699 10.6151
R1424 B.n699 B.n698 10.6151
R1425 B.n698 B.n67 10.6151
R1426 B.n694 B.n67 10.6151
R1427 B.n694 B.n693 10.6151
R1428 B.n693 B.n692 10.6151
R1429 B.n692 B.n69 10.6151
R1430 B.n688 B.n69 10.6151
R1431 B.n688 B.n687 10.6151
R1432 B.n687 B.n686 10.6151
R1433 B.n686 B.n71 10.6151
R1434 B.n682 B.n71 10.6151
R1435 B.n682 B.n681 10.6151
R1436 B.n681 B.n680 10.6151
R1437 B.n680 B.n73 10.6151
R1438 B.n676 B.n73 10.6151
R1439 B.n676 B.n675 10.6151
R1440 B.n675 B.n674 10.6151
R1441 B.n434 B.n155 10.6151
R1442 B.n435 B.n434 10.6151
R1443 B.n436 B.n435 10.6151
R1444 B.n436 B.n153 10.6151
R1445 B.n440 B.n153 10.6151
R1446 B.n441 B.n440 10.6151
R1447 B.n442 B.n441 10.6151
R1448 B.n442 B.n151 10.6151
R1449 B.n446 B.n151 10.6151
R1450 B.n447 B.n446 10.6151
R1451 B.n448 B.n447 10.6151
R1452 B.n448 B.n149 10.6151
R1453 B.n452 B.n149 10.6151
R1454 B.n453 B.n452 10.6151
R1455 B.n454 B.n453 10.6151
R1456 B.n454 B.n147 10.6151
R1457 B.n458 B.n147 10.6151
R1458 B.n459 B.n458 10.6151
R1459 B.n460 B.n459 10.6151
R1460 B.n460 B.n145 10.6151
R1461 B.n464 B.n145 10.6151
R1462 B.n465 B.n464 10.6151
R1463 B.n466 B.n465 10.6151
R1464 B.n466 B.n143 10.6151
R1465 B.n470 B.n143 10.6151
R1466 B.n471 B.n470 10.6151
R1467 B.n472 B.n471 10.6151
R1468 B.n472 B.n141 10.6151
R1469 B.n476 B.n141 10.6151
R1470 B.n477 B.n476 10.6151
R1471 B.n478 B.n477 10.6151
R1472 B.n478 B.n139 10.6151
R1473 B.n482 B.n139 10.6151
R1474 B.n483 B.n482 10.6151
R1475 B.n484 B.n483 10.6151
R1476 B.n484 B.n137 10.6151
R1477 B.n488 B.n137 10.6151
R1478 B.n489 B.n488 10.6151
R1479 B.n490 B.n489 10.6151
R1480 B.n490 B.n135 10.6151
R1481 B.n494 B.n135 10.6151
R1482 B.n495 B.n494 10.6151
R1483 B.n496 B.n495 10.6151
R1484 B.n496 B.n133 10.6151
R1485 B.n500 B.n133 10.6151
R1486 B.n501 B.n500 10.6151
R1487 B.n502 B.n501 10.6151
R1488 B.n502 B.n131 10.6151
R1489 B.n506 B.n131 10.6151
R1490 B.n507 B.n506 10.6151
R1491 B.n508 B.n507 10.6151
R1492 B.n508 B.n129 10.6151
R1493 B.n512 B.n129 10.6151
R1494 B.n513 B.n512 10.6151
R1495 B.n514 B.n513 10.6151
R1496 B.n514 B.n127 10.6151
R1497 B.n518 B.n127 10.6151
R1498 B.n519 B.n518 10.6151
R1499 B.n520 B.n519 10.6151
R1500 B.n520 B.n125 10.6151
R1501 B.n524 B.n125 10.6151
R1502 B.n525 B.n524 10.6151
R1503 B.n526 B.n525 10.6151
R1504 B.n526 B.n123 10.6151
R1505 B.n530 B.n123 10.6151
R1506 B.n531 B.n530 10.6151
R1507 B.n532 B.n531 10.6151
R1508 B.n532 B.n121 10.6151
R1509 B.n536 B.n121 10.6151
R1510 B.n537 B.n536 10.6151
R1511 B.n538 B.n537 10.6151
R1512 B.n538 B.n119 10.6151
R1513 B.n542 B.n119 10.6151
R1514 B.n543 B.n542 10.6151
R1515 B.n544 B.n543 10.6151
R1516 B.n544 B.n117 10.6151
R1517 B.n548 B.n117 10.6151
R1518 B.n549 B.n548 10.6151
R1519 B.n550 B.n549 10.6151
R1520 B.n550 B.n115 10.6151
R1521 B.n554 B.n115 10.6151
R1522 B.n555 B.n554 10.6151
R1523 B.n556 B.n555 10.6151
R1524 B.n556 B.n113 10.6151
R1525 B.n560 B.n113 10.6151
R1526 B.n561 B.n560 10.6151
R1527 B.n562 B.n561 10.6151
R1528 B.n562 B.n111 10.6151
R1529 B.n566 B.n111 10.6151
R1530 B.n567 B.n566 10.6151
R1531 B.n568 B.n567 10.6151
R1532 B.n568 B.n109 10.6151
R1533 B.n572 B.n109 10.6151
R1534 B.n573 B.n572 10.6151
R1535 B.n574 B.n573 10.6151
R1536 B.n574 B.n107 10.6151
R1537 B.n578 B.n107 10.6151
R1538 B.n579 B.n578 10.6151
R1539 B.n580 B.n579 10.6151
R1540 B.n580 B.n105 10.6151
R1541 B.n584 B.n105 10.6151
R1542 B.n585 B.n584 10.6151
R1543 B.n586 B.n585 10.6151
R1544 B.n586 B.n103 10.6151
R1545 B.n590 B.n103 10.6151
R1546 B.n591 B.n590 10.6151
R1547 B.n592 B.n591 10.6151
R1548 B.n592 B.n101 10.6151
R1549 B.n596 B.n101 10.6151
R1550 B.n597 B.n596 10.6151
R1551 B.n598 B.n597 10.6151
R1552 B.n598 B.n99 10.6151
R1553 B.n602 B.n99 10.6151
R1554 B.n603 B.n602 10.6151
R1555 B.n604 B.n603 10.6151
R1556 B.n604 B.n97 10.6151
R1557 B.n608 B.n97 10.6151
R1558 B.n609 B.n608 10.6151
R1559 B.n610 B.n609 10.6151
R1560 B.n610 B.n95 10.6151
R1561 B.n614 B.n95 10.6151
R1562 B.n615 B.n614 10.6151
R1563 B.n616 B.n615 10.6151
R1564 B.n616 B.n93 10.6151
R1565 B.n620 B.n93 10.6151
R1566 B.n621 B.n620 10.6151
R1567 B.n622 B.n621 10.6151
R1568 B.n622 B.n91 10.6151
R1569 B.n626 B.n91 10.6151
R1570 B.n627 B.n626 10.6151
R1571 B.n628 B.n627 10.6151
R1572 B.n628 B.n89 10.6151
R1573 B.n632 B.n89 10.6151
R1574 B.n633 B.n632 10.6151
R1575 B.n634 B.n633 10.6151
R1576 B.n634 B.n87 10.6151
R1577 B.n638 B.n87 10.6151
R1578 B.n639 B.n638 10.6151
R1579 B.n640 B.n639 10.6151
R1580 B.n640 B.n85 10.6151
R1581 B.n644 B.n85 10.6151
R1582 B.n645 B.n644 10.6151
R1583 B.n646 B.n645 10.6151
R1584 B.n646 B.n83 10.6151
R1585 B.n650 B.n83 10.6151
R1586 B.n651 B.n650 10.6151
R1587 B.n652 B.n651 10.6151
R1588 B.n652 B.n81 10.6151
R1589 B.n656 B.n81 10.6151
R1590 B.n657 B.n656 10.6151
R1591 B.n658 B.n657 10.6151
R1592 B.n658 B.n79 10.6151
R1593 B.n662 B.n79 10.6151
R1594 B.n663 B.n662 10.6151
R1595 B.n664 B.n663 10.6151
R1596 B.n664 B.n77 10.6151
R1597 B.n668 B.n77 10.6151
R1598 B.n669 B.n668 10.6151
R1599 B.n670 B.n669 10.6151
R1600 B.n670 B.n75 10.6151
R1601 B.n346 B.n187 10.6151
R1602 B.n350 B.n187 10.6151
R1603 B.n351 B.n350 10.6151
R1604 B.n352 B.n351 10.6151
R1605 B.n352 B.n185 10.6151
R1606 B.n356 B.n185 10.6151
R1607 B.n357 B.n356 10.6151
R1608 B.n358 B.n357 10.6151
R1609 B.n358 B.n183 10.6151
R1610 B.n362 B.n183 10.6151
R1611 B.n363 B.n362 10.6151
R1612 B.n364 B.n363 10.6151
R1613 B.n364 B.n181 10.6151
R1614 B.n368 B.n181 10.6151
R1615 B.n369 B.n368 10.6151
R1616 B.n370 B.n369 10.6151
R1617 B.n370 B.n179 10.6151
R1618 B.n374 B.n179 10.6151
R1619 B.n375 B.n374 10.6151
R1620 B.n376 B.n375 10.6151
R1621 B.n376 B.n177 10.6151
R1622 B.n380 B.n177 10.6151
R1623 B.n383 B.n382 10.6151
R1624 B.n383 B.n173 10.6151
R1625 B.n387 B.n173 10.6151
R1626 B.n388 B.n387 10.6151
R1627 B.n389 B.n388 10.6151
R1628 B.n389 B.n171 10.6151
R1629 B.n393 B.n171 10.6151
R1630 B.n394 B.n393 10.6151
R1631 B.n395 B.n394 10.6151
R1632 B.n399 B.n398 10.6151
R1633 B.n400 B.n399 10.6151
R1634 B.n400 B.n165 10.6151
R1635 B.n404 B.n165 10.6151
R1636 B.n405 B.n404 10.6151
R1637 B.n406 B.n405 10.6151
R1638 B.n406 B.n163 10.6151
R1639 B.n410 B.n163 10.6151
R1640 B.n411 B.n410 10.6151
R1641 B.n412 B.n411 10.6151
R1642 B.n412 B.n161 10.6151
R1643 B.n416 B.n161 10.6151
R1644 B.n417 B.n416 10.6151
R1645 B.n418 B.n417 10.6151
R1646 B.n418 B.n159 10.6151
R1647 B.n422 B.n159 10.6151
R1648 B.n423 B.n422 10.6151
R1649 B.n424 B.n423 10.6151
R1650 B.n424 B.n157 10.6151
R1651 B.n428 B.n157 10.6151
R1652 B.n429 B.n428 10.6151
R1653 B.n430 B.n429 10.6151
R1654 B.n345 B.n344 10.6151
R1655 B.n344 B.n189 10.6151
R1656 B.n340 B.n189 10.6151
R1657 B.n340 B.n339 10.6151
R1658 B.n339 B.n338 10.6151
R1659 B.n338 B.n191 10.6151
R1660 B.n334 B.n191 10.6151
R1661 B.n334 B.n333 10.6151
R1662 B.n333 B.n332 10.6151
R1663 B.n332 B.n193 10.6151
R1664 B.n328 B.n193 10.6151
R1665 B.n328 B.n327 10.6151
R1666 B.n327 B.n326 10.6151
R1667 B.n326 B.n195 10.6151
R1668 B.n322 B.n195 10.6151
R1669 B.n322 B.n321 10.6151
R1670 B.n321 B.n320 10.6151
R1671 B.n320 B.n197 10.6151
R1672 B.n316 B.n197 10.6151
R1673 B.n316 B.n315 10.6151
R1674 B.n315 B.n314 10.6151
R1675 B.n314 B.n199 10.6151
R1676 B.n310 B.n199 10.6151
R1677 B.n310 B.n309 10.6151
R1678 B.n309 B.n308 10.6151
R1679 B.n308 B.n201 10.6151
R1680 B.n304 B.n201 10.6151
R1681 B.n304 B.n303 10.6151
R1682 B.n303 B.n302 10.6151
R1683 B.n302 B.n203 10.6151
R1684 B.n298 B.n203 10.6151
R1685 B.n298 B.n297 10.6151
R1686 B.n297 B.n296 10.6151
R1687 B.n296 B.n205 10.6151
R1688 B.n292 B.n205 10.6151
R1689 B.n292 B.n291 10.6151
R1690 B.n291 B.n290 10.6151
R1691 B.n290 B.n207 10.6151
R1692 B.n286 B.n207 10.6151
R1693 B.n286 B.n285 10.6151
R1694 B.n285 B.n284 10.6151
R1695 B.n284 B.n209 10.6151
R1696 B.n280 B.n209 10.6151
R1697 B.n280 B.n279 10.6151
R1698 B.n279 B.n278 10.6151
R1699 B.n278 B.n211 10.6151
R1700 B.n274 B.n211 10.6151
R1701 B.n274 B.n273 10.6151
R1702 B.n273 B.n272 10.6151
R1703 B.n272 B.n213 10.6151
R1704 B.n268 B.n213 10.6151
R1705 B.n268 B.n267 10.6151
R1706 B.n267 B.n266 10.6151
R1707 B.n266 B.n215 10.6151
R1708 B.n262 B.n215 10.6151
R1709 B.n262 B.n261 10.6151
R1710 B.n261 B.n260 10.6151
R1711 B.n260 B.n217 10.6151
R1712 B.n256 B.n217 10.6151
R1713 B.n256 B.n255 10.6151
R1714 B.n255 B.n254 10.6151
R1715 B.n254 B.n219 10.6151
R1716 B.n250 B.n219 10.6151
R1717 B.n250 B.n249 10.6151
R1718 B.n249 B.n248 10.6151
R1719 B.n248 B.n221 10.6151
R1720 B.n244 B.n221 10.6151
R1721 B.n244 B.n243 10.6151
R1722 B.n243 B.n242 10.6151
R1723 B.n242 B.n223 10.6151
R1724 B.n238 B.n223 10.6151
R1725 B.n238 B.n237 10.6151
R1726 B.n237 B.n236 10.6151
R1727 B.n236 B.n225 10.6151
R1728 B.n232 B.n225 10.6151
R1729 B.n232 B.n231 10.6151
R1730 B.n231 B.n230 10.6151
R1731 B.n230 B.n227 10.6151
R1732 B.n227 B.n0 10.6151
R1733 B.n875 B.n1 10.6151
R1734 B.n875 B.n874 10.6151
R1735 B.n874 B.n873 10.6151
R1736 B.n873 B.n4 10.6151
R1737 B.n869 B.n4 10.6151
R1738 B.n869 B.n868 10.6151
R1739 B.n868 B.n867 10.6151
R1740 B.n867 B.n6 10.6151
R1741 B.n863 B.n6 10.6151
R1742 B.n863 B.n862 10.6151
R1743 B.n862 B.n861 10.6151
R1744 B.n861 B.n8 10.6151
R1745 B.n857 B.n8 10.6151
R1746 B.n857 B.n856 10.6151
R1747 B.n856 B.n855 10.6151
R1748 B.n855 B.n10 10.6151
R1749 B.n851 B.n10 10.6151
R1750 B.n851 B.n850 10.6151
R1751 B.n850 B.n849 10.6151
R1752 B.n849 B.n12 10.6151
R1753 B.n845 B.n12 10.6151
R1754 B.n845 B.n844 10.6151
R1755 B.n844 B.n843 10.6151
R1756 B.n843 B.n14 10.6151
R1757 B.n839 B.n14 10.6151
R1758 B.n839 B.n838 10.6151
R1759 B.n838 B.n837 10.6151
R1760 B.n837 B.n16 10.6151
R1761 B.n833 B.n16 10.6151
R1762 B.n833 B.n832 10.6151
R1763 B.n832 B.n831 10.6151
R1764 B.n831 B.n18 10.6151
R1765 B.n827 B.n18 10.6151
R1766 B.n827 B.n826 10.6151
R1767 B.n826 B.n825 10.6151
R1768 B.n825 B.n20 10.6151
R1769 B.n821 B.n20 10.6151
R1770 B.n821 B.n820 10.6151
R1771 B.n820 B.n819 10.6151
R1772 B.n819 B.n22 10.6151
R1773 B.n815 B.n22 10.6151
R1774 B.n815 B.n814 10.6151
R1775 B.n814 B.n813 10.6151
R1776 B.n813 B.n24 10.6151
R1777 B.n809 B.n24 10.6151
R1778 B.n809 B.n808 10.6151
R1779 B.n808 B.n807 10.6151
R1780 B.n807 B.n26 10.6151
R1781 B.n803 B.n26 10.6151
R1782 B.n803 B.n802 10.6151
R1783 B.n802 B.n801 10.6151
R1784 B.n801 B.n28 10.6151
R1785 B.n797 B.n28 10.6151
R1786 B.n797 B.n796 10.6151
R1787 B.n796 B.n795 10.6151
R1788 B.n795 B.n30 10.6151
R1789 B.n791 B.n30 10.6151
R1790 B.n791 B.n790 10.6151
R1791 B.n790 B.n789 10.6151
R1792 B.n789 B.n32 10.6151
R1793 B.n785 B.n32 10.6151
R1794 B.n785 B.n784 10.6151
R1795 B.n784 B.n783 10.6151
R1796 B.n783 B.n34 10.6151
R1797 B.n779 B.n34 10.6151
R1798 B.n779 B.n778 10.6151
R1799 B.n778 B.n777 10.6151
R1800 B.n777 B.n36 10.6151
R1801 B.n773 B.n36 10.6151
R1802 B.n773 B.n772 10.6151
R1803 B.n772 B.n771 10.6151
R1804 B.n771 B.n38 10.6151
R1805 B.n767 B.n38 10.6151
R1806 B.n767 B.n766 10.6151
R1807 B.n766 B.n765 10.6151
R1808 B.n765 B.n40 10.6151
R1809 B.n761 B.n40 10.6151
R1810 B.n761 B.n760 10.6151
R1811 B.n760 B.n759 10.6151
R1812 B.n724 B.n723 9.36635
R1813 B.n706 B.n64 9.36635
R1814 B.n381 B.n380 9.36635
R1815 B.n398 B.n169 9.36635
R1816 B.n879 B.n0 2.81026
R1817 B.n879 B.n1 2.81026
R1818 B.n723 B.n722 1.24928
R1819 B.n64 B.n60 1.24928
R1820 B.n382 B.n381 1.24928
R1821 B.n395 B.n169 1.24928
R1822 VP.n33 VP.n32 161.3
R1823 VP.n34 VP.n29 161.3
R1824 VP.n36 VP.n35 161.3
R1825 VP.n37 VP.n28 161.3
R1826 VP.n39 VP.n38 161.3
R1827 VP.n40 VP.n27 161.3
R1828 VP.n42 VP.n41 161.3
R1829 VP.n43 VP.n26 161.3
R1830 VP.n45 VP.n44 161.3
R1831 VP.n46 VP.n25 161.3
R1832 VP.n48 VP.n47 161.3
R1833 VP.n49 VP.n24 161.3
R1834 VP.n51 VP.n50 161.3
R1835 VP.n52 VP.n23 161.3
R1836 VP.n54 VP.n53 161.3
R1837 VP.n55 VP.n22 161.3
R1838 VP.n58 VP.n57 161.3
R1839 VP.n59 VP.n21 161.3
R1840 VP.n61 VP.n60 161.3
R1841 VP.n62 VP.n20 161.3
R1842 VP.n64 VP.n63 161.3
R1843 VP.n65 VP.n19 161.3
R1844 VP.n67 VP.n66 161.3
R1845 VP.n68 VP.n18 161.3
R1846 VP.n70 VP.n69 161.3
R1847 VP.n125 VP.n124 161.3
R1848 VP.n123 VP.n1 161.3
R1849 VP.n122 VP.n121 161.3
R1850 VP.n120 VP.n2 161.3
R1851 VP.n119 VP.n118 161.3
R1852 VP.n117 VP.n3 161.3
R1853 VP.n116 VP.n115 161.3
R1854 VP.n114 VP.n4 161.3
R1855 VP.n113 VP.n112 161.3
R1856 VP.n110 VP.n5 161.3
R1857 VP.n109 VP.n108 161.3
R1858 VP.n107 VP.n6 161.3
R1859 VP.n106 VP.n105 161.3
R1860 VP.n104 VP.n7 161.3
R1861 VP.n103 VP.n102 161.3
R1862 VP.n101 VP.n8 161.3
R1863 VP.n100 VP.n99 161.3
R1864 VP.n98 VP.n9 161.3
R1865 VP.n97 VP.n96 161.3
R1866 VP.n95 VP.n10 161.3
R1867 VP.n94 VP.n93 161.3
R1868 VP.n92 VP.n11 161.3
R1869 VP.n91 VP.n90 161.3
R1870 VP.n89 VP.n12 161.3
R1871 VP.n88 VP.n87 161.3
R1872 VP.n85 VP.n13 161.3
R1873 VP.n84 VP.n83 161.3
R1874 VP.n82 VP.n14 161.3
R1875 VP.n81 VP.n80 161.3
R1876 VP.n79 VP.n15 161.3
R1877 VP.n78 VP.n77 161.3
R1878 VP.n76 VP.n16 161.3
R1879 VP.n75 VP.n74 161.3
R1880 VP.n73 VP.n72 82.238
R1881 VP.n126 VP.n0 82.238
R1882 VP.n71 VP.n17 82.238
R1883 VP.n31 VP.n30 70.8482
R1884 VP.n30 VP.t8 70.3423
R1885 VP.n72 VP.n71 54.7948
R1886 VP.n80 VP.n79 52.1486
R1887 VP.n118 VP.n2 52.1486
R1888 VP.n63 VP.n19 52.1486
R1889 VP.n93 VP.n92 44.3785
R1890 VP.n105 VP.n6 44.3785
R1891 VP.n50 VP.n23 44.3785
R1892 VP.n38 VP.n37 44.3785
R1893 VP.n99 VP.t2 37.3394
R1894 VP.n73 VP.t5 37.3394
R1895 VP.n86 VP.t0 37.3394
R1896 VP.n111 VP.t3 37.3394
R1897 VP.n0 VP.t1 37.3394
R1898 VP.n44 VP.t6 37.3394
R1899 VP.n17 VP.t9 37.3394
R1900 VP.n56 VP.t7 37.3394
R1901 VP.n31 VP.t4 37.3394
R1902 VP.n93 VP.n10 36.6083
R1903 VP.n105 VP.n104 36.6083
R1904 VP.n50 VP.n49 36.6083
R1905 VP.n38 VP.n27 36.6083
R1906 VP.n80 VP.n14 28.8382
R1907 VP.n118 VP.n117 28.8382
R1908 VP.n63 VP.n62 28.8382
R1909 VP.n74 VP.n16 24.4675
R1910 VP.n78 VP.n16 24.4675
R1911 VP.n79 VP.n78 24.4675
R1912 VP.n84 VP.n14 24.4675
R1913 VP.n85 VP.n84 24.4675
R1914 VP.n87 VP.n12 24.4675
R1915 VP.n91 VP.n12 24.4675
R1916 VP.n92 VP.n91 24.4675
R1917 VP.n97 VP.n10 24.4675
R1918 VP.n98 VP.n97 24.4675
R1919 VP.n99 VP.n98 24.4675
R1920 VP.n99 VP.n8 24.4675
R1921 VP.n103 VP.n8 24.4675
R1922 VP.n104 VP.n103 24.4675
R1923 VP.n109 VP.n6 24.4675
R1924 VP.n110 VP.n109 24.4675
R1925 VP.n112 VP.n110 24.4675
R1926 VP.n116 VP.n4 24.4675
R1927 VP.n117 VP.n116 24.4675
R1928 VP.n122 VP.n2 24.4675
R1929 VP.n123 VP.n122 24.4675
R1930 VP.n124 VP.n123 24.4675
R1931 VP.n67 VP.n19 24.4675
R1932 VP.n68 VP.n67 24.4675
R1933 VP.n69 VP.n68 24.4675
R1934 VP.n54 VP.n23 24.4675
R1935 VP.n55 VP.n54 24.4675
R1936 VP.n57 VP.n55 24.4675
R1937 VP.n61 VP.n21 24.4675
R1938 VP.n62 VP.n61 24.4675
R1939 VP.n42 VP.n27 24.4675
R1940 VP.n43 VP.n42 24.4675
R1941 VP.n44 VP.n43 24.4675
R1942 VP.n44 VP.n25 24.4675
R1943 VP.n48 VP.n25 24.4675
R1944 VP.n49 VP.n48 24.4675
R1945 VP.n32 VP.n29 24.4675
R1946 VP.n36 VP.n29 24.4675
R1947 VP.n37 VP.n36 24.4675
R1948 VP.n86 VP.n85 20.5528
R1949 VP.n111 VP.n4 20.5528
R1950 VP.n56 VP.n21 20.5528
R1951 VP.n74 VP.n73 7.82994
R1952 VP.n124 VP.n0 7.82994
R1953 VP.n69 VP.n17 7.82994
R1954 VP.n87 VP.n86 3.91522
R1955 VP.n112 VP.n111 3.91522
R1956 VP.n57 VP.n56 3.91522
R1957 VP.n32 VP.n31 3.91522
R1958 VP.n33 VP.n30 3.22185
R1959 VP.n71 VP.n70 0.354971
R1960 VP.n75 VP.n72 0.354971
R1961 VP.n126 VP.n125 0.354971
R1962 VP VP.n126 0.26696
R1963 VP.n34 VP.n33 0.189894
R1964 VP.n35 VP.n34 0.189894
R1965 VP.n35 VP.n28 0.189894
R1966 VP.n39 VP.n28 0.189894
R1967 VP.n40 VP.n39 0.189894
R1968 VP.n41 VP.n40 0.189894
R1969 VP.n41 VP.n26 0.189894
R1970 VP.n45 VP.n26 0.189894
R1971 VP.n46 VP.n45 0.189894
R1972 VP.n47 VP.n46 0.189894
R1973 VP.n47 VP.n24 0.189894
R1974 VP.n51 VP.n24 0.189894
R1975 VP.n52 VP.n51 0.189894
R1976 VP.n53 VP.n52 0.189894
R1977 VP.n53 VP.n22 0.189894
R1978 VP.n58 VP.n22 0.189894
R1979 VP.n59 VP.n58 0.189894
R1980 VP.n60 VP.n59 0.189894
R1981 VP.n60 VP.n20 0.189894
R1982 VP.n64 VP.n20 0.189894
R1983 VP.n65 VP.n64 0.189894
R1984 VP.n66 VP.n65 0.189894
R1985 VP.n66 VP.n18 0.189894
R1986 VP.n70 VP.n18 0.189894
R1987 VP.n76 VP.n75 0.189894
R1988 VP.n77 VP.n76 0.189894
R1989 VP.n77 VP.n15 0.189894
R1990 VP.n81 VP.n15 0.189894
R1991 VP.n82 VP.n81 0.189894
R1992 VP.n83 VP.n82 0.189894
R1993 VP.n83 VP.n13 0.189894
R1994 VP.n88 VP.n13 0.189894
R1995 VP.n89 VP.n88 0.189894
R1996 VP.n90 VP.n89 0.189894
R1997 VP.n90 VP.n11 0.189894
R1998 VP.n94 VP.n11 0.189894
R1999 VP.n95 VP.n94 0.189894
R2000 VP.n96 VP.n95 0.189894
R2001 VP.n96 VP.n9 0.189894
R2002 VP.n100 VP.n9 0.189894
R2003 VP.n101 VP.n100 0.189894
R2004 VP.n102 VP.n101 0.189894
R2005 VP.n102 VP.n7 0.189894
R2006 VP.n106 VP.n7 0.189894
R2007 VP.n107 VP.n106 0.189894
R2008 VP.n108 VP.n107 0.189894
R2009 VP.n108 VP.n5 0.189894
R2010 VP.n113 VP.n5 0.189894
R2011 VP.n114 VP.n113 0.189894
R2012 VP.n115 VP.n114 0.189894
R2013 VP.n115 VP.n3 0.189894
R2014 VP.n119 VP.n3 0.189894
R2015 VP.n120 VP.n119 0.189894
R2016 VP.n121 VP.n120 0.189894
R2017 VP.n121 VP.n1 0.189894
R2018 VP.n125 VP.n1 0.189894
R2019 VDD1.n28 VDD1.n27 756.745
R2020 VDD1.n59 VDD1.n58 756.745
R2021 VDD1.n27 VDD1.n26 585
R2022 VDD1.n2 VDD1.n1 585
R2023 VDD1.n21 VDD1.n20 585
R2024 VDD1.n19 VDD1.n18 585
R2025 VDD1.n6 VDD1.n5 585
R2026 VDD1.n13 VDD1.n12 585
R2027 VDD1.n11 VDD1.n10 585
R2028 VDD1.n42 VDD1.n41 585
R2029 VDD1.n44 VDD1.n43 585
R2030 VDD1.n37 VDD1.n36 585
R2031 VDD1.n50 VDD1.n49 585
R2032 VDD1.n52 VDD1.n51 585
R2033 VDD1.n33 VDD1.n32 585
R2034 VDD1.n58 VDD1.n57 585
R2035 VDD1.n40 VDD1.t4 329.175
R2036 VDD1.n9 VDD1.t1 329.175
R2037 VDD1.n27 VDD1.n1 171.744
R2038 VDD1.n20 VDD1.n1 171.744
R2039 VDD1.n20 VDD1.n19 171.744
R2040 VDD1.n19 VDD1.n5 171.744
R2041 VDD1.n12 VDD1.n5 171.744
R2042 VDD1.n12 VDD1.n11 171.744
R2043 VDD1.n43 VDD1.n42 171.744
R2044 VDD1.n43 VDD1.n36 171.744
R2045 VDD1.n50 VDD1.n36 171.744
R2046 VDD1.n51 VDD1.n50 171.744
R2047 VDD1.n51 VDD1.n32 171.744
R2048 VDD1.n58 VDD1.n32 171.744
R2049 VDD1.n63 VDD1.n62 97.5006
R2050 VDD1.n30 VDD1.n29 94.919
R2051 VDD1.n61 VDD1.n60 94.918
R2052 VDD1.n65 VDD1.n64 94.9178
R2053 VDD1.n11 VDD1.t1 85.8723
R2054 VDD1.n42 VDD1.t4 85.8723
R2055 VDD1.n30 VDD1.n28 54.5147
R2056 VDD1.n61 VDD1.n59 54.5147
R2057 VDD1.n65 VDD1.n63 47.7724
R2058 VDD1.n26 VDD1.n0 12.0247
R2059 VDD1.n57 VDD1.n31 12.0247
R2060 VDD1.n25 VDD1.n2 11.249
R2061 VDD1.n56 VDD1.n33 11.249
R2062 VDD1.n41 VDD1.n40 10.722
R2063 VDD1.n10 VDD1.n9 10.722
R2064 VDD1.n22 VDD1.n21 10.4732
R2065 VDD1.n53 VDD1.n52 10.4732
R2066 VDD1.n18 VDD1.n4 9.69747
R2067 VDD1.n49 VDD1.n35 9.69747
R2068 VDD1.n24 VDD1.n0 9.45567
R2069 VDD1.n55 VDD1.n31 9.45567
R2070 VDD1.n15 VDD1.n14 9.3005
R2071 VDD1.n17 VDD1.n16 9.3005
R2072 VDD1.n4 VDD1.n3 9.3005
R2073 VDD1.n23 VDD1.n22 9.3005
R2074 VDD1.n25 VDD1.n24 9.3005
R2075 VDD1.n8 VDD1.n7 9.3005
R2076 VDD1.n39 VDD1.n38 9.3005
R2077 VDD1.n46 VDD1.n45 9.3005
R2078 VDD1.n48 VDD1.n47 9.3005
R2079 VDD1.n35 VDD1.n34 9.3005
R2080 VDD1.n54 VDD1.n53 9.3005
R2081 VDD1.n56 VDD1.n55 9.3005
R2082 VDD1.n17 VDD1.n6 8.92171
R2083 VDD1.n48 VDD1.n37 8.92171
R2084 VDD1.n14 VDD1.n13 8.14595
R2085 VDD1.n45 VDD1.n44 8.14595
R2086 VDD1.n10 VDD1.n8 7.3702
R2087 VDD1.n41 VDD1.n39 7.3702
R2088 VDD1.n13 VDD1.n8 5.81868
R2089 VDD1.n44 VDD1.n39 5.81868
R2090 VDD1.n64 VDD1.t2 5.59516
R2091 VDD1.n64 VDD1.t0 5.59516
R2092 VDD1.n29 VDD1.t5 5.59516
R2093 VDD1.n29 VDD1.t3 5.59516
R2094 VDD1.n62 VDD1.t6 5.59516
R2095 VDD1.n62 VDD1.t8 5.59516
R2096 VDD1.n60 VDD1.t9 5.59516
R2097 VDD1.n60 VDD1.t7 5.59516
R2098 VDD1.n14 VDD1.n6 5.04292
R2099 VDD1.n45 VDD1.n37 5.04292
R2100 VDD1.n18 VDD1.n17 4.26717
R2101 VDD1.n49 VDD1.n48 4.26717
R2102 VDD1.n21 VDD1.n4 3.49141
R2103 VDD1.n52 VDD1.n35 3.49141
R2104 VDD1.n22 VDD1.n2 2.71565
R2105 VDD1.n53 VDD1.n33 2.71565
R2106 VDD1 VDD1.n65 2.58024
R2107 VDD1.n40 VDD1.n38 2.4147
R2108 VDD1.n9 VDD1.n7 2.4147
R2109 VDD1.n26 VDD1.n25 1.93989
R2110 VDD1.n57 VDD1.n56 1.93989
R2111 VDD1.n28 VDD1.n0 1.16414
R2112 VDD1.n59 VDD1.n31 1.16414
R2113 VDD1 VDD1.n30 0.938
R2114 VDD1.n63 VDD1.n61 0.824464
R2115 VDD1.n24 VDD1.n23 0.155672
R2116 VDD1.n23 VDD1.n3 0.155672
R2117 VDD1.n16 VDD1.n3 0.155672
R2118 VDD1.n16 VDD1.n15 0.155672
R2119 VDD1.n15 VDD1.n7 0.155672
R2120 VDD1.n46 VDD1.n38 0.155672
R2121 VDD1.n47 VDD1.n46 0.155672
R2122 VDD1.n47 VDD1.n34 0.155672
R2123 VDD1.n54 VDD1.n34 0.155672
R2124 VDD1.n55 VDD1.n54 0.155672
C0 VN B 1.49586f
C1 VN VDD1 0.15585f
C2 VTAIL VN 7.50061f
C3 w_n5866_n2130# VP 13.5609f
C4 B VP 2.79241f
C5 w_n5866_n2130# B 10.762f
C6 VDD2 VN 5.78605f
C7 VDD1 VP 6.35681f
C8 w_n5866_n2130# VDD1 2.79876f
C9 VTAIL VP 7.51496f
C10 B VDD1 2.42729f
C11 VTAIL w_n5866_n2130# 2.5328f
C12 VTAIL B 2.67223f
C13 VTAIL VDD1 8.56394f
C14 VDD2 VP 0.729631f
C15 VDD2 w_n5866_n2130# 3.00204f
C16 VDD2 B 2.59007f
C17 VDD2 VDD1 2.92219f
C18 VDD2 VTAIL 8.624499f
C19 VN VP 8.94608f
C20 VN w_n5866_n2130# 12.793599f
C21 VDD2 VSUBS 2.534949f
C22 VDD1 VSUBS 2.310606f
C23 VTAIL VSUBS 0.799623f
C24 VN VSUBS 9.40225f
C25 VP VSUBS 5.182269f
C26 B VSUBS 6.271456f
C27 w_n5866_n2130# VSUBS 0.156059p
C28 VDD1.n0 VSUBS 0.020167f
C29 VDD1.n1 VSUBS 0.045487f
C30 VDD1.n2 VSUBS 0.020377f
C31 VDD1.n3 VSUBS 0.035813f
C32 VDD1.n4 VSUBS 0.019245f
C33 VDD1.n5 VSUBS 0.045487f
C34 VDD1.n6 VSUBS 0.020377f
C35 VDD1.n7 VSUBS 0.787087f
C36 VDD1.n8 VSUBS 0.019245f
C37 VDD1.t1 VSUBS 0.097948f
C38 VDD1.n9 VSUBS 0.182352f
C39 VDD1.n10 VSUBS 0.034203f
C40 VDD1.n11 VSUBS 0.034115f
C41 VDD1.n12 VSUBS 0.045487f
C42 VDD1.n13 VSUBS 0.020377f
C43 VDD1.n14 VSUBS 0.019245f
C44 VDD1.n15 VSUBS 0.035813f
C45 VDD1.n16 VSUBS 0.035813f
C46 VDD1.n17 VSUBS 0.019245f
C47 VDD1.n18 VSUBS 0.020377f
C48 VDD1.n19 VSUBS 0.045487f
C49 VDD1.n20 VSUBS 0.045487f
C50 VDD1.n21 VSUBS 0.020377f
C51 VDD1.n22 VSUBS 0.019245f
C52 VDD1.n23 VSUBS 0.035813f
C53 VDD1.n24 VSUBS 0.091098f
C54 VDD1.n25 VSUBS 0.019245f
C55 VDD1.n26 VSUBS 0.020377f
C56 VDD1.n27 VSUBS 0.099784f
C57 VDD1.n28 VSUBS 0.122172f
C58 VDD1.t5 VSUBS 0.164428f
C59 VDD1.t3 VSUBS 0.164428f
C60 VDD1.n29 VSUBS 1.10443f
C61 VDD1.n30 VSUBS 1.51242f
C62 VDD1.n31 VSUBS 0.020167f
C63 VDD1.n32 VSUBS 0.045487f
C64 VDD1.n33 VSUBS 0.020377f
C65 VDD1.n34 VSUBS 0.035813f
C66 VDD1.n35 VSUBS 0.019245f
C67 VDD1.n36 VSUBS 0.045487f
C68 VDD1.n37 VSUBS 0.020377f
C69 VDD1.n38 VSUBS 0.787087f
C70 VDD1.n39 VSUBS 0.019245f
C71 VDD1.t4 VSUBS 0.097948f
C72 VDD1.n40 VSUBS 0.182352f
C73 VDD1.n41 VSUBS 0.034203f
C74 VDD1.n42 VSUBS 0.034115f
C75 VDD1.n43 VSUBS 0.045487f
C76 VDD1.n44 VSUBS 0.020377f
C77 VDD1.n45 VSUBS 0.019245f
C78 VDD1.n46 VSUBS 0.035813f
C79 VDD1.n47 VSUBS 0.035813f
C80 VDD1.n48 VSUBS 0.019245f
C81 VDD1.n49 VSUBS 0.020377f
C82 VDD1.n50 VSUBS 0.045487f
C83 VDD1.n51 VSUBS 0.045487f
C84 VDD1.n52 VSUBS 0.020377f
C85 VDD1.n53 VSUBS 0.019245f
C86 VDD1.n54 VSUBS 0.035813f
C87 VDD1.n55 VSUBS 0.091098f
C88 VDD1.n56 VSUBS 0.019245f
C89 VDD1.n57 VSUBS 0.020377f
C90 VDD1.n58 VSUBS 0.099784f
C91 VDD1.n59 VSUBS 0.122172f
C92 VDD1.t9 VSUBS 0.164428f
C93 VDD1.t7 VSUBS 0.164428f
C94 VDD1.n60 VSUBS 1.10443f
C95 VDD1.n61 VSUBS 1.50033f
C96 VDD1.t6 VSUBS 0.164428f
C97 VDD1.t8 VSUBS 0.164428f
C98 VDD1.n62 VSUBS 1.13807f
C99 VDD1.n63 VSUBS 4.95212f
C100 VDD1.t2 VSUBS 0.164428f
C101 VDD1.t0 VSUBS 0.164428f
C102 VDD1.n64 VSUBS 1.10442f
C103 VDD1.n65 VSUBS 4.80778f
C104 VP.t1 VSUBS 2.00987f
C105 VP.n0 VSUBS 0.881911f
C106 VP.n1 VSUBS 0.03492f
C107 VP.n2 VSUBS 0.062692f
C108 VP.n3 VSUBS 0.03492f
C109 VP.n4 VSUBS 0.059942f
C110 VP.n5 VSUBS 0.03492f
C111 VP.n6 VSUBS 0.067675f
C112 VP.n7 VSUBS 0.03492f
C113 VP.n8 VSUBS 0.065083f
C114 VP.n9 VSUBS 0.03492f
C115 VP.t2 VSUBS 2.00987f
C116 VP.n10 VSUBS 0.070409f
C117 VP.n11 VSUBS 0.03492f
C118 VP.n12 VSUBS 0.065083f
C119 VP.n13 VSUBS 0.03492f
C120 VP.t0 VSUBS 2.00987f
C121 VP.n14 VSUBS 0.069074f
C122 VP.n15 VSUBS 0.03492f
C123 VP.n16 VSUBS 0.065083f
C124 VP.t9 VSUBS 2.00987f
C125 VP.n17 VSUBS 0.881911f
C126 VP.n18 VSUBS 0.03492f
C127 VP.n19 VSUBS 0.062692f
C128 VP.n20 VSUBS 0.03492f
C129 VP.n21 VSUBS 0.059942f
C130 VP.n22 VSUBS 0.03492f
C131 VP.n23 VSUBS 0.067675f
C132 VP.n24 VSUBS 0.03492f
C133 VP.n25 VSUBS 0.065083f
C134 VP.n26 VSUBS 0.03492f
C135 VP.t6 VSUBS 2.00987f
C136 VP.n27 VSUBS 0.070409f
C137 VP.n28 VSUBS 0.03492f
C138 VP.n29 VSUBS 0.065083f
C139 VP.t8 VSUBS 2.48547f
C140 VP.n30 VSUBS 0.828335f
C141 VP.t4 VSUBS 2.00987f
C142 VP.n31 VSUBS 0.856713f
C143 VP.n32 VSUBS 0.038092f
C144 VP.n33 VSUBS 0.443451f
C145 VP.n34 VSUBS 0.03492f
C146 VP.n35 VSUBS 0.03492f
C147 VP.n36 VSUBS 0.065083f
C148 VP.n37 VSUBS 0.067675f
C149 VP.n38 VSUBS 0.028954f
C150 VP.n39 VSUBS 0.03492f
C151 VP.n40 VSUBS 0.03492f
C152 VP.n41 VSUBS 0.03492f
C153 VP.n42 VSUBS 0.065083f
C154 VP.n43 VSUBS 0.065083f
C155 VP.n44 VSUBS 0.775814f
C156 VP.n45 VSUBS 0.03492f
C157 VP.n46 VSUBS 0.03492f
C158 VP.n47 VSUBS 0.03492f
C159 VP.n48 VSUBS 0.065083f
C160 VP.n49 VSUBS 0.070409f
C161 VP.n50 VSUBS 0.028954f
C162 VP.n51 VSUBS 0.03492f
C163 VP.n52 VSUBS 0.03492f
C164 VP.n53 VSUBS 0.03492f
C165 VP.n54 VSUBS 0.065083f
C166 VP.n55 VSUBS 0.065083f
C167 VP.t7 VSUBS 2.00987f
C168 VP.n56 VSUBS 0.742863f
C169 VP.n57 VSUBS 0.038092f
C170 VP.n58 VSUBS 0.03492f
C171 VP.n59 VSUBS 0.03492f
C172 VP.n60 VSUBS 0.03492f
C173 VP.n61 VSUBS 0.065083f
C174 VP.n62 VSUBS 0.069074f
C175 VP.n63 VSUBS 0.035271f
C176 VP.n64 VSUBS 0.03492f
C177 VP.n65 VSUBS 0.03492f
C178 VP.n66 VSUBS 0.03492f
C179 VP.n67 VSUBS 0.065083f
C180 VP.n68 VSUBS 0.065083f
C181 VP.n69 VSUBS 0.043233f
C182 VP.n70 VSUBS 0.056361f
C183 VP.n71 VSUBS 2.27861f
C184 VP.n72 VSUBS 2.30152f
C185 VP.t5 VSUBS 2.00987f
C186 VP.n73 VSUBS 0.881911f
C187 VP.n74 VSUBS 0.043233f
C188 VP.n75 VSUBS 0.056361f
C189 VP.n76 VSUBS 0.03492f
C190 VP.n77 VSUBS 0.03492f
C191 VP.n78 VSUBS 0.065083f
C192 VP.n79 VSUBS 0.062692f
C193 VP.n80 VSUBS 0.035271f
C194 VP.n81 VSUBS 0.03492f
C195 VP.n82 VSUBS 0.03492f
C196 VP.n83 VSUBS 0.03492f
C197 VP.n84 VSUBS 0.065083f
C198 VP.n85 VSUBS 0.059942f
C199 VP.n86 VSUBS 0.742863f
C200 VP.n87 VSUBS 0.038092f
C201 VP.n88 VSUBS 0.03492f
C202 VP.n89 VSUBS 0.03492f
C203 VP.n90 VSUBS 0.03492f
C204 VP.n91 VSUBS 0.065083f
C205 VP.n92 VSUBS 0.067675f
C206 VP.n93 VSUBS 0.028954f
C207 VP.n94 VSUBS 0.03492f
C208 VP.n95 VSUBS 0.03492f
C209 VP.n96 VSUBS 0.03492f
C210 VP.n97 VSUBS 0.065083f
C211 VP.n98 VSUBS 0.065083f
C212 VP.n99 VSUBS 0.775814f
C213 VP.n100 VSUBS 0.03492f
C214 VP.n101 VSUBS 0.03492f
C215 VP.n102 VSUBS 0.03492f
C216 VP.n103 VSUBS 0.065083f
C217 VP.n104 VSUBS 0.070409f
C218 VP.n105 VSUBS 0.028954f
C219 VP.n106 VSUBS 0.03492f
C220 VP.n107 VSUBS 0.03492f
C221 VP.n108 VSUBS 0.03492f
C222 VP.n109 VSUBS 0.065083f
C223 VP.n110 VSUBS 0.065083f
C224 VP.t3 VSUBS 2.00987f
C225 VP.n111 VSUBS 0.742863f
C226 VP.n112 VSUBS 0.038092f
C227 VP.n113 VSUBS 0.03492f
C228 VP.n114 VSUBS 0.03492f
C229 VP.n115 VSUBS 0.03492f
C230 VP.n116 VSUBS 0.065083f
C231 VP.n117 VSUBS 0.069074f
C232 VP.n118 VSUBS 0.035271f
C233 VP.n119 VSUBS 0.03492f
C234 VP.n120 VSUBS 0.03492f
C235 VP.n121 VSUBS 0.03492f
C236 VP.n122 VSUBS 0.065083f
C237 VP.n123 VSUBS 0.065083f
C238 VP.n124 VSUBS 0.043233f
C239 VP.n125 VSUBS 0.056361f
C240 VP.n126 VSUBS 0.100743f
C241 B.n0 VSUBS 0.007395f
C242 B.n1 VSUBS 0.007395f
C243 B.n2 VSUBS 0.011694f
C244 B.n3 VSUBS 0.011694f
C245 B.n4 VSUBS 0.011694f
C246 B.n5 VSUBS 0.011694f
C247 B.n6 VSUBS 0.011694f
C248 B.n7 VSUBS 0.011694f
C249 B.n8 VSUBS 0.011694f
C250 B.n9 VSUBS 0.011694f
C251 B.n10 VSUBS 0.011694f
C252 B.n11 VSUBS 0.011694f
C253 B.n12 VSUBS 0.011694f
C254 B.n13 VSUBS 0.011694f
C255 B.n14 VSUBS 0.011694f
C256 B.n15 VSUBS 0.011694f
C257 B.n16 VSUBS 0.011694f
C258 B.n17 VSUBS 0.011694f
C259 B.n18 VSUBS 0.011694f
C260 B.n19 VSUBS 0.011694f
C261 B.n20 VSUBS 0.011694f
C262 B.n21 VSUBS 0.011694f
C263 B.n22 VSUBS 0.011694f
C264 B.n23 VSUBS 0.011694f
C265 B.n24 VSUBS 0.011694f
C266 B.n25 VSUBS 0.011694f
C267 B.n26 VSUBS 0.011694f
C268 B.n27 VSUBS 0.011694f
C269 B.n28 VSUBS 0.011694f
C270 B.n29 VSUBS 0.011694f
C271 B.n30 VSUBS 0.011694f
C272 B.n31 VSUBS 0.011694f
C273 B.n32 VSUBS 0.011694f
C274 B.n33 VSUBS 0.011694f
C275 B.n34 VSUBS 0.011694f
C276 B.n35 VSUBS 0.011694f
C277 B.n36 VSUBS 0.011694f
C278 B.n37 VSUBS 0.011694f
C279 B.n38 VSUBS 0.011694f
C280 B.n39 VSUBS 0.011694f
C281 B.n40 VSUBS 0.011694f
C282 B.n41 VSUBS 0.011694f
C283 B.n42 VSUBS 0.029572f
C284 B.n43 VSUBS 0.011694f
C285 B.n44 VSUBS 0.011694f
C286 B.n45 VSUBS 0.011694f
C287 B.n46 VSUBS 0.011694f
C288 B.n47 VSUBS 0.011694f
C289 B.n48 VSUBS 0.011694f
C290 B.n49 VSUBS 0.011694f
C291 B.n50 VSUBS 0.011694f
C292 B.n51 VSUBS 0.011694f
C293 B.n52 VSUBS 0.011694f
C294 B.n53 VSUBS 0.011694f
C295 B.t2 VSUBS 0.143371f
C296 B.t1 VSUBS 0.200312f
C297 B.t0 VSUBS 1.751f
C298 B.n54 VSUBS 0.332713f
C299 B.n55 VSUBS 0.263965f
C300 B.n56 VSUBS 0.011694f
C301 B.n57 VSUBS 0.011694f
C302 B.n58 VSUBS 0.011694f
C303 B.n59 VSUBS 0.011694f
C304 B.n60 VSUBS 0.006535f
C305 B.n61 VSUBS 0.011694f
C306 B.t11 VSUBS 0.143374f
C307 B.t10 VSUBS 0.200315f
C308 B.t9 VSUBS 1.751f
C309 B.n62 VSUBS 0.33271f
C310 B.n63 VSUBS 0.263962f
C311 B.n64 VSUBS 0.027095f
C312 B.n65 VSUBS 0.011694f
C313 B.n66 VSUBS 0.011694f
C314 B.n67 VSUBS 0.011694f
C315 B.n68 VSUBS 0.011694f
C316 B.n69 VSUBS 0.011694f
C317 B.n70 VSUBS 0.011694f
C318 B.n71 VSUBS 0.011694f
C319 B.n72 VSUBS 0.011694f
C320 B.n73 VSUBS 0.011694f
C321 B.n74 VSUBS 0.011694f
C322 B.n75 VSUBS 0.029818f
C323 B.n76 VSUBS 0.011694f
C324 B.n77 VSUBS 0.011694f
C325 B.n78 VSUBS 0.011694f
C326 B.n79 VSUBS 0.011694f
C327 B.n80 VSUBS 0.011694f
C328 B.n81 VSUBS 0.011694f
C329 B.n82 VSUBS 0.011694f
C330 B.n83 VSUBS 0.011694f
C331 B.n84 VSUBS 0.011694f
C332 B.n85 VSUBS 0.011694f
C333 B.n86 VSUBS 0.011694f
C334 B.n87 VSUBS 0.011694f
C335 B.n88 VSUBS 0.011694f
C336 B.n89 VSUBS 0.011694f
C337 B.n90 VSUBS 0.011694f
C338 B.n91 VSUBS 0.011694f
C339 B.n92 VSUBS 0.011694f
C340 B.n93 VSUBS 0.011694f
C341 B.n94 VSUBS 0.011694f
C342 B.n95 VSUBS 0.011694f
C343 B.n96 VSUBS 0.011694f
C344 B.n97 VSUBS 0.011694f
C345 B.n98 VSUBS 0.011694f
C346 B.n99 VSUBS 0.011694f
C347 B.n100 VSUBS 0.011694f
C348 B.n101 VSUBS 0.011694f
C349 B.n102 VSUBS 0.011694f
C350 B.n103 VSUBS 0.011694f
C351 B.n104 VSUBS 0.011694f
C352 B.n105 VSUBS 0.011694f
C353 B.n106 VSUBS 0.011694f
C354 B.n107 VSUBS 0.011694f
C355 B.n108 VSUBS 0.011694f
C356 B.n109 VSUBS 0.011694f
C357 B.n110 VSUBS 0.011694f
C358 B.n111 VSUBS 0.011694f
C359 B.n112 VSUBS 0.011694f
C360 B.n113 VSUBS 0.011694f
C361 B.n114 VSUBS 0.011694f
C362 B.n115 VSUBS 0.011694f
C363 B.n116 VSUBS 0.011694f
C364 B.n117 VSUBS 0.011694f
C365 B.n118 VSUBS 0.011694f
C366 B.n119 VSUBS 0.011694f
C367 B.n120 VSUBS 0.011694f
C368 B.n121 VSUBS 0.011694f
C369 B.n122 VSUBS 0.011694f
C370 B.n123 VSUBS 0.011694f
C371 B.n124 VSUBS 0.011694f
C372 B.n125 VSUBS 0.011694f
C373 B.n126 VSUBS 0.011694f
C374 B.n127 VSUBS 0.011694f
C375 B.n128 VSUBS 0.011694f
C376 B.n129 VSUBS 0.011694f
C377 B.n130 VSUBS 0.011694f
C378 B.n131 VSUBS 0.011694f
C379 B.n132 VSUBS 0.011694f
C380 B.n133 VSUBS 0.011694f
C381 B.n134 VSUBS 0.011694f
C382 B.n135 VSUBS 0.011694f
C383 B.n136 VSUBS 0.011694f
C384 B.n137 VSUBS 0.011694f
C385 B.n138 VSUBS 0.011694f
C386 B.n139 VSUBS 0.011694f
C387 B.n140 VSUBS 0.011694f
C388 B.n141 VSUBS 0.011694f
C389 B.n142 VSUBS 0.011694f
C390 B.n143 VSUBS 0.011694f
C391 B.n144 VSUBS 0.011694f
C392 B.n145 VSUBS 0.011694f
C393 B.n146 VSUBS 0.011694f
C394 B.n147 VSUBS 0.011694f
C395 B.n148 VSUBS 0.011694f
C396 B.n149 VSUBS 0.011694f
C397 B.n150 VSUBS 0.011694f
C398 B.n151 VSUBS 0.011694f
C399 B.n152 VSUBS 0.011694f
C400 B.n153 VSUBS 0.011694f
C401 B.n154 VSUBS 0.011694f
C402 B.n155 VSUBS 0.028556f
C403 B.n156 VSUBS 0.011694f
C404 B.n157 VSUBS 0.011694f
C405 B.n158 VSUBS 0.011694f
C406 B.n159 VSUBS 0.011694f
C407 B.n160 VSUBS 0.011694f
C408 B.n161 VSUBS 0.011694f
C409 B.n162 VSUBS 0.011694f
C410 B.n163 VSUBS 0.011694f
C411 B.n164 VSUBS 0.011694f
C412 B.n165 VSUBS 0.011694f
C413 B.n166 VSUBS 0.011694f
C414 B.t7 VSUBS 0.143374f
C415 B.t8 VSUBS 0.200315f
C416 B.t6 VSUBS 1.751f
C417 B.n167 VSUBS 0.33271f
C418 B.n168 VSUBS 0.263962f
C419 B.n169 VSUBS 0.027095f
C420 B.n170 VSUBS 0.011694f
C421 B.n171 VSUBS 0.011694f
C422 B.n172 VSUBS 0.011694f
C423 B.n173 VSUBS 0.011694f
C424 B.n174 VSUBS 0.011694f
C425 B.t4 VSUBS 0.143371f
C426 B.t5 VSUBS 0.200312f
C427 B.t3 VSUBS 1.751f
C428 B.n175 VSUBS 0.332713f
C429 B.n176 VSUBS 0.263965f
C430 B.n177 VSUBS 0.011694f
C431 B.n178 VSUBS 0.011694f
C432 B.n179 VSUBS 0.011694f
C433 B.n180 VSUBS 0.011694f
C434 B.n181 VSUBS 0.011694f
C435 B.n182 VSUBS 0.011694f
C436 B.n183 VSUBS 0.011694f
C437 B.n184 VSUBS 0.011694f
C438 B.n185 VSUBS 0.011694f
C439 B.n186 VSUBS 0.011694f
C440 B.n187 VSUBS 0.011694f
C441 B.n188 VSUBS 0.028556f
C442 B.n189 VSUBS 0.011694f
C443 B.n190 VSUBS 0.011694f
C444 B.n191 VSUBS 0.011694f
C445 B.n192 VSUBS 0.011694f
C446 B.n193 VSUBS 0.011694f
C447 B.n194 VSUBS 0.011694f
C448 B.n195 VSUBS 0.011694f
C449 B.n196 VSUBS 0.011694f
C450 B.n197 VSUBS 0.011694f
C451 B.n198 VSUBS 0.011694f
C452 B.n199 VSUBS 0.011694f
C453 B.n200 VSUBS 0.011694f
C454 B.n201 VSUBS 0.011694f
C455 B.n202 VSUBS 0.011694f
C456 B.n203 VSUBS 0.011694f
C457 B.n204 VSUBS 0.011694f
C458 B.n205 VSUBS 0.011694f
C459 B.n206 VSUBS 0.011694f
C460 B.n207 VSUBS 0.011694f
C461 B.n208 VSUBS 0.011694f
C462 B.n209 VSUBS 0.011694f
C463 B.n210 VSUBS 0.011694f
C464 B.n211 VSUBS 0.011694f
C465 B.n212 VSUBS 0.011694f
C466 B.n213 VSUBS 0.011694f
C467 B.n214 VSUBS 0.011694f
C468 B.n215 VSUBS 0.011694f
C469 B.n216 VSUBS 0.011694f
C470 B.n217 VSUBS 0.011694f
C471 B.n218 VSUBS 0.011694f
C472 B.n219 VSUBS 0.011694f
C473 B.n220 VSUBS 0.011694f
C474 B.n221 VSUBS 0.011694f
C475 B.n222 VSUBS 0.011694f
C476 B.n223 VSUBS 0.011694f
C477 B.n224 VSUBS 0.011694f
C478 B.n225 VSUBS 0.011694f
C479 B.n226 VSUBS 0.011694f
C480 B.n227 VSUBS 0.011694f
C481 B.n228 VSUBS 0.011694f
C482 B.n229 VSUBS 0.011694f
C483 B.n230 VSUBS 0.011694f
C484 B.n231 VSUBS 0.011694f
C485 B.n232 VSUBS 0.011694f
C486 B.n233 VSUBS 0.011694f
C487 B.n234 VSUBS 0.011694f
C488 B.n235 VSUBS 0.011694f
C489 B.n236 VSUBS 0.011694f
C490 B.n237 VSUBS 0.011694f
C491 B.n238 VSUBS 0.011694f
C492 B.n239 VSUBS 0.011694f
C493 B.n240 VSUBS 0.011694f
C494 B.n241 VSUBS 0.011694f
C495 B.n242 VSUBS 0.011694f
C496 B.n243 VSUBS 0.011694f
C497 B.n244 VSUBS 0.011694f
C498 B.n245 VSUBS 0.011694f
C499 B.n246 VSUBS 0.011694f
C500 B.n247 VSUBS 0.011694f
C501 B.n248 VSUBS 0.011694f
C502 B.n249 VSUBS 0.011694f
C503 B.n250 VSUBS 0.011694f
C504 B.n251 VSUBS 0.011694f
C505 B.n252 VSUBS 0.011694f
C506 B.n253 VSUBS 0.011694f
C507 B.n254 VSUBS 0.011694f
C508 B.n255 VSUBS 0.011694f
C509 B.n256 VSUBS 0.011694f
C510 B.n257 VSUBS 0.011694f
C511 B.n258 VSUBS 0.011694f
C512 B.n259 VSUBS 0.011694f
C513 B.n260 VSUBS 0.011694f
C514 B.n261 VSUBS 0.011694f
C515 B.n262 VSUBS 0.011694f
C516 B.n263 VSUBS 0.011694f
C517 B.n264 VSUBS 0.011694f
C518 B.n265 VSUBS 0.011694f
C519 B.n266 VSUBS 0.011694f
C520 B.n267 VSUBS 0.011694f
C521 B.n268 VSUBS 0.011694f
C522 B.n269 VSUBS 0.011694f
C523 B.n270 VSUBS 0.011694f
C524 B.n271 VSUBS 0.011694f
C525 B.n272 VSUBS 0.011694f
C526 B.n273 VSUBS 0.011694f
C527 B.n274 VSUBS 0.011694f
C528 B.n275 VSUBS 0.011694f
C529 B.n276 VSUBS 0.011694f
C530 B.n277 VSUBS 0.011694f
C531 B.n278 VSUBS 0.011694f
C532 B.n279 VSUBS 0.011694f
C533 B.n280 VSUBS 0.011694f
C534 B.n281 VSUBS 0.011694f
C535 B.n282 VSUBS 0.011694f
C536 B.n283 VSUBS 0.011694f
C537 B.n284 VSUBS 0.011694f
C538 B.n285 VSUBS 0.011694f
C539 B.n286 VSUBS 0.011694f
C540 B.n287 VSUBS 0.011694f
C541 B.n288 VSUBS 0.011694f
C542 B.n289 VSUBS 0.011694f
C543 B.n290 VSUBS 0.011694f
C544 B.n291 VSUBS 0.011694f
C545 B.n292 VSUBS 0.011694f
C546 B.n293 VSUBS 0.011694f
C547 B.n294 VSUBS 0.011694f
C548 B.n295 VSUBS 0.011694f
C549 B.n296 VSUBS 0.011694f
C550 B.n297 VSUBS 0.011694f
C551 B.n298 VSUBS 0.011694f
C552 B.n299 VSUBS 0.011694f
C553 B.n300 VSUBS 0.011694f
C554 B.n301 VSUBS 0.011694f
C555 B.n302 VSUBS 0.011694f
C556 B.n303 VSUBS 0.011694f
C557 B.n304 VSUBS 0.011694f
C558 B.n305 VSUBS 0.011694f
C559 B.n306 VSUBS 0.011694f
C560 B.n307 VSUBS 0.011694f
C561 B.n308 VSUBS 0.011694f
C562 B.n309 VSUBS 0.011694f
C563 B.n310 VSUBS 0.011694f
C564 B.n311 VSUBS 0.011694f
C565 B.n312 VSUBS 0.011694f
C566 B.n313 VSUBS 0.011694f
C567 B.n314 VSUBS 0.011694f
C568 B.n315 VSUBS 0.011694f
C569 B.n316 VSUBS 0.011694f
C570 B.n317 VSUBS 0.011694f
C571 B.n318 VSUBS 0.011694f
C572 B.n319 VSUBS 0.011694f
C573 B.n320 VSUBS 0.011694f
C574 B.n321 VSUBS 0.011694f
C575 B.n322 VSUBS 0.011694f
C576 B.n323 VSUBS 0.011694f
C577 B.n324 VSUBS 0.011694f
C578 B.n325 VSUBS 0.011694f
C579 B.n326 VSUBS 0.011694f
C580 B.n327 VSUBS 0.011694f
C581 B.n328 VSUBS 0.011694f
C582 B.n329 VSUBS 0.011694f
C583 B.n330 VSUBS 0.011694f
C584 B.n331 VSUBS 0.011694f
C585 B.n332 VSUBS 0.011694f
C586 B.n333 VSUBS 0.011694f
C587 B.n334 VSUBS 0.011694f
C588 B.n335 VSUBS 0.011694f
C589 B.n336 VSUBS 0.011694f
C590 B.n337 VSUBS 0.011694f
C591 B.n338 VSUBS 0.011694f
C592 B.n339 VSUBS 0.011694f
C593 B.n340 VSUBS 0.011694f
C594 B.n341 VSUBS 0.011694f
C595 B.n342 VSUBS 0.011694f
C596 B.n343 VSUBS 0.011694f
C597 B.n344 VSUBS 0.011694f
C598 B.n345 VSUBS 0.028556f
C599 B.n346 VSUBS 0.029572f
C600 B.n347 VSUBS 0.029572f
C601 B.n348 VSUBS 0.011694f
C602 B.n349 VSUBS 0.011694f
C603 B.n350 VSUBS 0.011694f
C604 B.n351 VSUBS 0.011694f
C605 B.n352 VSUBS 0.011694f
C606 B.n353 VSUBS 0.011694f
C607 B.n354 VSUBS 0.011694f
C608 B.n355 VSUBS 0.011694f
C609 B.n356 VSUBS 0.011694f
C610 B.n357 VSUBS 0.011694f
C611 B.n358 VSUBS 0.011694f
C612 B.n359 VSUBS 0.011694f
C613 B.n360 VSUBS 0.011694f
C614 B.n361 VSUBS 0.011694f
C615 B.n362 VSUBS 0.011694f
C616 B.n363 VSUBS 0.011694f
C617 B.n364 VSUBS 0.011694f
C618 B.n365 VSUBS 0.011694f
C619 B.n366 VSUBS 0.011694f
C620 B.n367 VSUBS 0.011694f
C621 B.n368 VSUBS 0.011694f
C622 B.n369 VSUBS 0.011694f
C623 B.n370 VSUBS 0.011694f
C624 B.n371 VSUBS 0.011694f
C625 B.n372 VSUBS 0.011694f
C626 B.n373 VSUBS 0.011694f
C627 B.n374 VSUBS 0.011694f
C628 B.n375 VSUBS 0.011694f
C629 B.n376 VSUBS 0.011694f
C630 B.n377 VSUBS 0.011694f
C631 B.n378 VSUBS 0.011694f
C632 B.n379 VSUBS 0.011694f
C633 B.n380 VSUBS 0.011006f
C634 B.n381 VSUBS 0.027095f
C635 B.n382 VSUBS 0.006535f
C636 B.n383 VSUBS 0.011694f
C637 B.n384 VSUBS 0.011694f
C638 B.n385 VSUBS 0.011694f
C639 B.n386 VSUBS 0.011694f
C640 B.n387 VSUBS 0.011694f
C641 B.n388 VSUBS 0.011694f
C642 B.n389 VSUBS 0.011694f
C643 B.n390 VSUBS 0.011694f
C644 B.n391 VSUBS 0.011694f
C645 B.n392 VSUBS 0.011694f
C646 B.n393 VSUBS 0.011694f
C647 B.n394 VSUBS 0.011694f
C648 B.n395 VSUBS 0.006535f
C649 B.n396 VSUBS 0.011694f
C650 B.n397 VSUBS 0.011694f
C651 B.n398 VSUBS 0.011006f
C652 B.n399 VSUBS 0.011694f
C653 B.n400 VSUBS 0.011694f
C654 B.n401 VSUBS 0.011694f
C655 B.n402 VSUBS 0.011694f
C656 B.n403 VSUBS 0.011694f
C657 B.n404 VSUBS 0.011694f
C658 B.n405 VSUBS 0.011694f
C659 B.n406 VSUBS 0.011694f
C660 B.n407 VSUBS 0.011694f
C661 B.n408 VSUBS 0.011694f
C662 B.n409 VSUBS 0.011694f
C663 B.n410 VSUBS 0.011694f
C664 B.n411 VSUBS 0.011694f
C665 B.n412 VSUBS 0.011694f
C666 B.n413 VSUBS 0.011694f
C667 B.n414 VSUBS 0.011694f
C668 B.n415 VSUBS 0.011694f
C669 B.n416 VSUBS 0.011694f
C670 B.n417 VSUBS 0.011694f
C671 B.n418 VSUBS 0.011694f
C672 B.n419 VSUBS 0.011694f
C673 B.n420 VSUBS 0.011694f
C674 B.n421 VSUBS 0.011694f
C675 B.n422 VSUBS 0.011694f
C676 B.n423 VSUBS 0.011694f
C677 B.n424 VSUBS 0.011694f
C678 B.n425 VSUBS 0.011694f
C679 B.n426 VSUBS 0.011694f
C680 B.n427 VSUBS 0.011694f
C681 B.n428 VSUBS 0.011694f
C682 B.n429 VSUBS 0.011694f
C683 B.n430 VSUBS 0.029572f
C684 B.n431 VSUBS 0.029572f
C685 B.n432 VSUBS 0.028556f
C686 B.n433 VSUBS 0.011694f
C687 B.n434 VSUBS 0.011694f
C688 B.n435 VSUBS 0.011694f
C689 B.n436 VSUBS 0.011694f
C690 B.n437 VSUBS 0.011694f
C691 B.n438 VSUBS 0.011694f
C692 B.n439 VSUBS 0.011694f
C693 B.n440 VSUBS 0.011694f
C694 B.n441 VSUBS 0.011694f
C695 B.n442 VSUBS 0.011694f
C696 B.n443 VSUBS 0.011694f
C697 B.n444 VSUBS 0.011694f
C698 B.n445 VSUBS 0.011694f
C699 B.n446 VSUBS 0.011694f
C700 B.n447 VSUBS 0.011694f
C701 B.n448 VSUBS 0.011694f
C702 B.n449 VSUBS 0.011694f
C703 B.n450 VSUBS 0.011694f
C704 B.n451 VSUBS 0.011694f
C705 B.n452 VSUBS 0.011694f
C706 B.n453 VSUBS 0.011694f
C707 B.n454 VSUBS 0.011694f
C708 B.n455 VSUBS 0.011694f
C709 B.n456 VSUBS 0.011694f
C710 B.n457 VSUBS 0.011694f
C711 B.n458 VSUBS 0.011694f
C712 B.n459 VSUBS 0.011694f
C713 B.n460 VSUBS 0.011694f
C714 B.n461 VSUBS 0.011694f
C715 B.n462 VSUBS 0.011694f
C716 B.n463 VSUBS 0.011694f
C717 B.n464 VSUBS 0.011694f
C718 B.n465 VSUBS 0.011694f
C719 B.n466 VSUBS 0.011694f
C720 B.n467 VSUBS 0.011694f
C721 B.n468 VSUBS 0.011694f
C722 B.n469 VSUBS 0.011694f
C723 B.n470 VSUBS 0.011694f
C724 B.n471 VSUBS 0.011694f
C725 B.n472 VSUBS 0.011694f
C726 B.n473 VSUBS 0.011694f
C727 B.n474 VSUBS 0.011694f
C728 B.n475 VSUBS 0.011694f
C729 B.n476 VSUBS 0.011694f
C730 B.n477 VSUBS 0.011694f
C731 B.n478 VSUBS 0.011694f
C732 B.n479 VSUBS 0.011694f
C733 B.n480 VSUBS 0.011694f
C734 B.n481 VSUBS 0.011694f
C735 B.n482 VSUBS 0.011694f
C736 B.n483 VSUBS 0.011694f
C737 B.n484 VSUBS 0.011694f
C738 B.n485 VSUBS 0.011694f
C739 B.n486 VSUBS 0.011694f
C740 B.n487 VSUBS 0.011694f
C741 B.n488 VSUBS 0.011694f
C742 B.n489 VSUBS 0.011694f
C743 B.n490 VSUBS 0.011694f
C744 B.n491 VSUBS 0.011694f
C745 B.n492 VSUBS 0.011694f
C746 B.n493 VSUBS 0.011694f
C747 B.n494 VSUBS 0.011694f
C748 B.n495 VSUBS 0.011694f
C749 B.n496 VSUBS 0.011694f
C750 B.n497 VSUBS 0.011694f
C751 B.n498 VSUBS 0.011694f
C752 B.n499 VSUBS 0.011694f
C753 B.n500 VSUBS 0.011694f
C754 B.n501 VSUBS 0.011694f
C755 B.n502 VSUBS 0.011694f
C756 B.n503 VSUBS 0.011694f
C757 B.n504 VSUBS 0.011694f
C758 B.n505 VSUBS 0.011694f
C759 B.n506 VSUBS 0.011694f
C760 B.n507 VSUBS 0.011694f
C761 B.n508 VSUBS 0.011694f
C762 B.n509 VSUBS 0.011694f
C763 B.n510 VSUBS 0.011694f
C764 B.n511 VSUBS 0.011694f
C765 B.n512 VSUBS 0.011694f
C766 B.n513 VSUBS 0.011694f
C767 B.n514 VSUBS 0.011694f
C768 B.n515 VSUBS 0.011694f
C769 B.n516 VSUBS 0.011694f
C770 B.n517 VSUBS 0.011694f
C771 B.n518 VSUBS 0.011694f
C772 B.n519 VSUBS 0.011694f
C773 B.n520 VSUBS 0.011694f
C774 B.n521 VSUBS 0.011694f
C775 B.n522 VSUBS 0.011694f
C776 B.n523 VSUBS 0.011694f
C777 B.n524 VSUBS 0.011694f
C778 B.n525 VSUBS 0.011694f
C779 B.n526 VSUBS 0.011694f
C780 B.n527 VSUBS 0.011694f
C781 B.n528 VSUBS 0.011694f
C782 B.n529 VSUBS 0.011694f
C783 B.n530 VSUBS 0.011694f
C784 B.n531 VSUBS 0.011694f
C785 B.n532 VSUBS 0.011694f
C786 B.n533 VSUBS 0.011694f
C787 B.n534 VSUBS 0.011694f
C788 B.n535 VSUBS 0.011694f
C789 B.n536 VSUBS 0.011694f
C790 B.n537 VSUBS 0.011694f
C791 B.n538 VSUBS 0.011694f
C792 B.n539 VSUBS 0.011694f
C793 B.n540 VSUBS 0.011694f
C794 B.n541 VSUBS 0.011694f
C795 B.n542 VSUBS 0.011694f
C796 B.n543 VSUBS 0.011694f
C797 B.n544 VSUBS 0.011694f
C798 B.n545 VSUBS 0.011694f
C799 B.n546 VSUBS 0.011694f
C800 B.n547 VSUBS 0.011694f
C801 B.n548 VSUBS 0.011694f
C802 B.n549 VSUBS 0.011694f
C803 B.n550 VSUBS 0.011694f
C804 B.n551 VSUBS 0.011694f
C805 B.n552 VSUBS 0.011694f
C806 B.n553 VSUBS 0.011694f
C807 B.n554 VSUBS 0.011694f
C808 B.n555 VSUBS 0.011694f
C809 B.n556 VSUBS 0.011694f
C810 B.n557 VSUBS 0.011694f
C811 B.n558 VSUBS 0.011694f
C812 B.n559 VSUBS 0.011694f
C813 B.n560 VSUBS 0.011694f
C814 B.n561 VSUBS 0.011694f
C815 B.n562 VSUBS 0.011694f
C816 B.n563 VSUBS 0.011694f
C817 B.n564 VSUBS 0.011694f
C818 B.n565 VSUBS 0.011694f
C819 B.n566 VSUBS 0.011694f
C820 B.n567 VSUBS 0.011694f
C821 B.n568 VSUBS 0.011694f
C822 B.n569 VSUBS 0.011694f
C823 B.n570 VSUBS 0.011694f
C824 B.n571 VSUBS 0.011694f
C825 B.n572 VSUBS 0.011694f
C826 B.n573 VSUBS 0.011694f
C827 B.n574 VSUBS 0.011694f
C828 B.n575 VSUBS 0.011694f
C829 B.n576 VSUBS 0.011694f
C830 B.n577 VSUBS 0.011694f
C831 B.n578 VSUBS 0.011694f
C832 B.n579 VSUBS 0.011694f
C833 B.n580 VSUBS 0.011694f
C834 B.n581 VSUBS 0.011694f
C835 B.n582 VSUBS 0.011694f
C836 B.n583 VSUBS 0.011694f
C837 B.n584 VSUBS 0.011694f
C838 B.n585 VSUBS 0.011694f
C839 B.n586 VSUBS 0.011694f
C840 B.n587 VSUBS 0.011694f
C841 B.n588 VSUBS 0.011694f
C842 B.n589 VSUBS 0.011694f
C843 B.n590 VSUBS 0.011694f
C844 B.n591 VSUBS 0.011694f
C845 B.n592 VSUBS 0.011694f
C846 B.n593 VSUBS 0.011694f
C847 B.n594 VSUBS 0.011694f
C848 B.n595 VSUBS 0.011694f
C849 B.n596 VSUBS 0.011694f
C850 B.n597 VSUBS 0.011694f
C851 B.n598 VSUBS 0.011694f
C852 B.n599 VSUBS 0.011694f
C853 B.n600 VSUBS 0.011694f
C854 B.n601 VSUBS 0.011694f
C855 B.n602 VSUBS 0.011694f
C856 B.n603 VSUBS 0.011694f
C857 B.n604 VSUBS 0.011694f
C858 B.n605 VSUBS 0.011694f
C859 B.n606 VSUBS 0.011694f
C860 B.n607 VSUBS 0.011694f
C861 B.n608 VSUBS 0.011694f
C862 B.n609 VSUBS 0.011694f
C863 B.n610 VSUBS 0.011694f
C864 B.n611 VSUBS 0.011694f
C865 B.n612 VSUBS 0.011694f
C866 B.n613 VSUBS 0.011694f
C867 B.n614 VSUBS 0.011694f
C868 B.n615 VSUBS 0.011694f
C869 B.n616 VSUBS 0.011694f
C870 B.n617 VSUBS 0.011694f
C871 B.n618 VSUBS 0.011694f
C872 B.n619 VSUBS 0.011694f
C873 B.n620 VSUBS 0.011694f
C874 B.n621 VSUBS 0.011694f
C875 B.n622 VSUBS 0.011694f
C876 B.n623 VSUBS 0.011694f
C877 B.n624 VSUBS 0.011694f
C878 B.n625 VSUBS 0.011694f
C879 B.n626 VSUBS 0.011694f
C880 B.n627 VSUBS 0.011694f
C881 B.n628 VSUBS 0.011694f
C882 B.n629 VSUBS 0.011694f
C883 B.n630 VSUBS 0.011694f
C884 B.n631 VSUBS 0.011694f
C885 B.n632 VSUBS 0.011694f
C886 B.n633 VSUBS 0.011694f
C887 B.n634 VSUBS 0.011694f
C888 B.n635 VSUBS 0.011694f
C889 B.n636 VSUBS 0.011694f
C890 B.n637 VSUBS 0.011694f
C891 B.n638 VSUBS 0.011694f
C892 B.n639 VSUBS 0.011694f
C893 B.n640 VSUBS 0.011694f
C894 B.n641 VSUBS 0.011694f
C895 B.n642 VSUBS 0.011694f
C896 B.n643 VSUBS 0.011694f
C897 B.n644 VSUBS 0.011694f
C898 B.n645 VSUBS 0.011694f
C899 B.n646 VSUBS 0.011694f
C900 B.n647 VSUBS 0.011694f
C901 B.n648 VSUBS 0.011694f
C902 B.n649 VSUBS 0.011694f
C903 B.n650 VSUBS 0.011694f
C904 B.n651 VSUBS 0.011694f
C905 B.n652 VSUBS 0.011694f
C906 B.n653 VSUBS 0.011694f
C907 B.n654 VSUBS 0.011694f
C908 B.n655 VSUBS 0.011694f
C909 B.n656 VSUBS 0.011694f
C910 B.n657 VSUBS 0.011694f
C911 B.n658 VSUBS 0.011694f
C912 B.n659 VSUBS 0.011694f
C913 B.n660 VSUBS 0.011694f
C914 B.n661 VSUBS 0.011694f
C915 B.n662 VSUBS 0.011694f
C916 B.n663 VSUBS 0.011694f
C917 B.n664 VSUBS 0.011694f
C918 B.n665 VSUBS 0.011694f
C919 B.n666 VSUBS 0.011694f
C920 B.n667 VSUBS 0.011694f
C921 B.n668 VSUBS 0.011694f
C922 B.n669 VSUBS 0.011694f
C923 B.n670 VSUBS 0.011694f
C924 B.n671 VSUBS 0.011694f
C925 B.n672 VSUBS 0.028556f
C926 B.n673 VSUBS 0.029572f
C927 B.n674 VSUBS 0.028309f
C928 B.n675 VSUBS 0.011694f
C929 B.n676 VSUBS 0.011694f
C930 B.n677 VSUBS 0.011694f
C931 B.n678 VSUBS 0.011694f
C932 B.n679 VSUBS 0.011694f
C933 B.n680 VSUBS 0.011694f
C934 B.n681 VSUBS 0.011694f
C935 B.n682 VSUBS 0.011694f
C936 B.n683 VSUBS 0.011694f
C937 B.n684 VSUBS 0.011694f
C938 B.n685 VSUBS 0.011694f
C939 B.n686 VSUBS 0.011694f
C940 B.n687 VSUBS 0.011694f
C941 B.n688 VSUBS 0.011694f
C942 B.n689 VSUBS 0.011694f
C943 B.n690 VSUBS 0.011694f
C944 B.n691 VSUBS 0.011694f
C945 B.n692 VSUBS 0.011694f
C946 B.n693 VSUBS 0.011694f
C947 B.n694 VSUBS 0.011694f
C948 B.n695 VSUBS 0.011694f
C949 B.n696 VSUBS 0.011694f
C950 B.n697 VSUBS 0.011694f
C951 B.n698 VSUBS 0.011694f
C952 B.n699 VSUBS 0.011694f
C953 B.n700 VSUBS 0.011694f
C954 B.n701 VSUBS 0.011694f
C955 B.n702 VSUBS 0.011694f
C956 B.n703 VSUBS 0.011694f
C957 B.n704 VSUBS 0.011694f
C958 B.n705 VSUBS 0.011694f
C959 B.n706 VSUBS 0.011006f
C960 B.n707 VSUBS 0.011694f
C961 B.n708 VSUBS 0.011694f
C962 B.n709 VSUBS 0.011694f
C963 B.n710 VSUBS 0.011694f
C964 B.n711 VSUBS 0.011694f
C965 B.n712 VSUBS 0.011694f
C966 B.n713 VSUBS 0.011694f
C967 B.n714 VSUBS 0.011694f
C968 B.n715 VSUBS 0.011694f
C969 B.n716 VSUBS 0.011694f
C970 B.n717 VSUBS 0.011694f
C971 B.n718 VSUBS 0.011694f
C972 B.n719 VSUBS 0.011694f
C973 B.n720 VSUBS 0.011694f
C974 B.n721 VSUBS 0.011694f
C975 B.n722 VSUBS 0.006535f
C976 B.n723 VSUBS 0.027095f
C977 B.n724 VSUBS 0.011006f
C978 B.n725 VSUBS 0.011694f
C979 B.n726 VSUBS 0.011694f
C980 B.n727 VSUBS 0.011694f
C981 B.n728 VSUBS 0.011694f
C982 B.n729 VSUBS 0.011694f
C983 B.n730 VSUBS 0.011694f
C984 B.n731 VSUBS 0.011694f
C985 B.n732 VSUBS 0.011694f
C986 B.n733 VSUBS 0.011694f
C987 B.n734 VSUBS 0.011694f
C988 B.n735 VSUBS 0.011694f
C989 B.n736 VSUBS 0.011694f
C990 B.n737 VSUBS 0.011694f
C991 B.n738 VSUBS 0.011694f
C992 B.n739 VSUBS 0.011694f
C993 B.n740 VSUBS 0.011694f
C994 B.n741 VSUBS 0.011694f
C995 B.n742 VSUBS 0.011694f
C996 B.n743 VSUBS 0.011694f
C997 B.n744 VSUBS 0.011694f
C998 B.n745 VSUBS 0.011694f
C999 B.n746 VSUBS 0.011694f
C1000 B.n747 VSUBS 0.011694f
C1001 B.n748 VSUBS 0.011694f
C1002 B.n749 VSUBS 0.011694f
C1003 B.n750 VSUBS 0.011694f
C1004 B.n751 VSUBS 0.011694f
C1005 B.n752 VSUBS 0.011694f
C1006 B.n753 VSUBS 0.011694f
C1007 B.n754 VSUBS 0.011694f
C1008 B.n755 VSUBS 0.011694f
C1009 B.n756 VSUBS 0.011694f
C1010 B.n757 VSUBS 0.029572f
C1011 B.n758 VSUBS 0.028556f
C1012 B.n759 VSUBS 0.028556f
C1013 B.n760 VSUBS 0.011694f
C1014 B.n761 VSUBS 0.011694f
C1015 B.n762 VSUBS 0.011694f
C1016 B.n763 VSUBS 0.011694f
C1017 B.n764 VSUBS 0.011694f
C1018 B.n765 VSUBS 0.011694f
C1019 B.n766 VSUBS 0.011694f
C1020 B.n767 VSUBS 0.011694f
C1021 B.n768 VSUBS 0.011694f
C1022 B.n769 VSUBS 0.011694f
C1023 B.n770 VSUBS 0.011694f
C1024 B.n771 VSUBS 0.011694f
C1025 B.n772 VSUBS 0.011694f
C1026 B.n773 VSUBS 0.011694f
C1027 B.n774 VSUBS 0.011694f
C1028 B.n775 VSUBS 0.011694f
C1029 B.n776 VSUBS 0.011694f
C1030 B.n777 VSUBS 0.011694f
C1031 B.n778 VSUBS 0.011694f
C1032 B.n779 VSUBS 0.011694f
C1033 B.n780 VSUBS 0.011694f
C1034 B.n781 VSUBS 0.011694f
C1035 B.n782 VSUBS 0.011694f
C1036 B.n783 VSUBS 0.011694f
C1037 B.n784 VSUBS 0.011694f
C1038 B.n785 VSUBS 0.011694f
C1039 B.n786 VSUBS 0.011694f
C1040 B.n787 VSUBS 0.011694f
C1041 B.n788 VSUBS 0.011694f
C1042 B.n789 VSUBS 0.011694f
C1043 B.n790 VSUBS 0.011694f
C1044 B.n791 VSUBS 0.011694f
C1045 B.n792 VSUBS 0.011694f
C1046 B.n793 VSUBS 0.011694f
C1047 B.n794 VSUBS 0.011694f
C1048 B.n795 VSUBS 0.011694f
C1049 B.n796 VSUBS 0.011694f
C1050 B.n797 VSUBS 0.011694f
C1051 B.n798 VSUBS 0.011694f
C1052 B.n799 VSUBS 0.011694f
C1053 B.n800 VSUBS 0.011694f
C1054 B.n801 VSUBS 0.011694f
C1055 B.n802 VSUBS 0.011694f
C1056 B.n803 VSUBS 0.011694f
C1057 B.n804 VSUBS 0.011694f
C1058 B.n805 VSUBS 0.011694f
C1059 B.n806 VSUBS 0.011694f
C1060 B.n807 VSUBS 0.011694f
C1061 B.n808 VSUBS 0.011694f
C1062 B.n809 VSUBS 0.011694f
C1063 B.n810 VSUBS 0.011694f
C1064 B.n811 VSUBS 0.011694f
C1065 B.n812 VSUBS 0.011694f
C1066 B.n813 VSUBS 0.011694f
C1067 B.n814 VSUBS 0.011694f
C1068 B.n815 VSUBS 0.011694f
C1069 B.n816 VSUBS 0.011694f
C1070 B.n817 VSUBS 0.011694f
C1071 B.n818 VSUBS 0.011694f
C1072 B.n819 VSUBS 0.011694f
C1073 B.n820 VSUBS 0.011694f
C1074 B.n821 VSUBS 0.011694f
C1075 B.n822 VSUBS 0.011694f
C1076 B.n823 VSUBS 0.011694f
C1077 B.n824 VSUBS 0.011694f
C1078 B.n825 VSUBS 0.011694f
C1079 B.n826 VSUBS 0.011694f
C1080 B.n827 VSUBS 0.011694f
C1081 B.n828 VSUBS 0.011694f
C1082 B.n829 VSUBS 0.011694f
C1083 B.n830 VSUBS 0.011694f
C1084 B.n831 VSUBS 0.011694f
C1085 B.n832 VSUBS 0.011694f
C1086 B.n833 VSUBS 0.011694f
C1087 B.n834 VSUBS 0.011694f
C1088 B.n835 VSUBS 0.011694f
C1089 B.n836 VSUBS 0.011694f
C1090 B.n837 VSUBS 0.011694f
C1091 B.n838 VSUBS 0.011694f
C1092 B.n839 VSUBS 0.011694f
C1093 B.n840 VSUBS 0.011694f
C1094 B.n841 VSUBS 0.011694f
C1095 B.n842 VSUBS 0.011694f
C1096 B.n843 VSUBS 0.011694f
C1097 B.n844 VSUBS 0.011694f
C1098 B.n845 VSUBS 0.011694f
C1099 B.n846 VSUBS 0.011694f
C1100 B.n847 VSUBS 0.011694f
C1101 B.n848 VSUBS 0.011694f
C1102 B.n849 VSUBS 0.011694f
C1103 B.n850 VSUBS 0.011694f
C1104 B.n851 VSUBS 0.011694f
C1105 B.n852 VSUBS 0.011694f
C1106 B.n853 VSUBS 0.011694f
C1107 B.n854 VSUBS 0.011694f
C1108 B.n855 VSUBS 0.011694f
C1109 B.n856 VSUBS 0.011694f
C1110 B.n857 VSUBS 0.011694f
C1111 B.n858 VSUBS 0.011694f
C1112 B.n859 VSUBS 0.011694f
C1113 B.n860 VSUBS 0.011694f
C1114 B.n861 VSUBS 0.011694f
C1115 B.n862 VSUBS 0.011694f
C1116 B.n863 VSUBS 0.011694f
C1117 B.n864 VSUBS 0.011694f
C1118 B.n865 VSUBS 0.011694f
C1119 B.n866 VSUBS 0.011694f
C1120 B.n867 VSUBS 0.011694f
C1121 B.n868 VSUBS 0.011694f
C1122 B.n869 VSUBS 0.011694f
C1123 B.n870 VSUBS 0.011694f
C1124 B.n871 VSUBS 0.011694f
C1125 B.n872 VSUBS 0.011694f
C1126 B.n873 VSUBS 0.011694f
C1127 B.n874 VSUBS 0.011694f
C1128 B.n875 VSUBS 0.011694f
C1129 B.n876 VSUBS 0.011694f
C1130 B.n877 VSUBS 0.011694f
C1131 B.n878 VSUBS 0.011694f
C1132 B.n879 VSUBS 0.02648f
C1133 VDD2.n0 VSUBS 0.020108f
C1134 VDD2.n1 VSUBS 0.045353f
C1135 VDD2.n2 VSUBS 0.020317f
C1136 VDD2.n3 VSUBS 0.035708f
C1137 VDD2.n4 VSUBS 0.019188f
C1138 VDD2.n5 VSUBS 0.045353f
C1139 VDD2.n6 VSUBS 0.020317f
C1140 VDD2.n7 VSUBS 0.784766f
C1141 VDD2.n8 VSUBS 0.019188f
C1142 VDD2.t2 VSUBS 0.097659f
C1143 VDD2.n9 VSUBS 0.181814f
C1144 VDD2.n10 VSUBS 0.034102f
C1145 VDD2.n11 VSUBS 0.034015f
C1146 VDD2.n12 VSUBS 0.045353f
C1147 VDD2.n13 VSUBS 0.020317f
C1148 VDD2.n14 VSUBS 0.019188f
C1149 VDD2.n15 VSUBS 0.035708f
C1150 VDD2.n16 VSUBS 0.035708f
C1151 VDD2.n17 VSUBS 0.019188f
C1152 VDD2.n18 VSUBS 0.020317f
C1153 VDD2.n19 VSUBS 0.045353f
C1154 VDD2.n20 VSUBS 0.045353f
C1155 VDD2.n21 VSUBS 0.020317f
C1156 VDD2.n22 VSUBS 0.019188f
C1157 VDD2.n23 VSUBS 0.035708f
C1158 VDD2.n24 VSUBS 0.09083f
C1159 VDD2.n25 VSUBS 0.019188f
C1160 VDD2.n26 VSUBS 0.020317f
C1161 VDD2.n27 VSUBS 0.09949f
C1162 VDD2.n28 VSUBS 0.121812f
C1163 VDD2.t6 VSUBS 0.163943f
C1164 VDD2.t8 VSUBS 0.163943f
C1165 VDD2.n29 VSUBS 1.10117f
C1166 VDD2.n30 VSUBS 1.49591f
C1167 VDD2.t7 VSUBS 0.163943f
C1168 VDD2.t9 VSUBS 0.163943f
C1169 VDD2.n31 VSUBS 1.13471f
C1170 VDD2.n32 VSUBS 4.72182f
C1171 VDD2.n33 VSUBS 0.020108f
C1172 VDD2.n34 VSUBS 0.045353f
C1173 VDD2.n35 VSUBS 0.020317f
C1174 VDD2.n36 VSUBS 0.035708f
C1175 VDD2.n37 VSUBS 0.019188f
C1176 VDD2.n38 VSUBS 0.045353f
C1177 VDD2.n39 VSUBS 0.020317f
C1178 VDD2.n40 VSUBS 0.784766f
C1179 VDD2.n41 VSUBS 0.019188f
C1180 VDD2.t0 VSUBS 0.097659f
C1181 VDD2.n42 VSUBS 0.181814f
C1182 VDD2.n43 VSUBS 0.034102f
C1183 VDD2.n44 VSUBS 0.034015f
C1184 VDD2.n45 VSUBS 0.045353f
C1185 VDD2.n46 VSUBS 0.020317f
C1186 VDD2.n47 VSUBS 0.019188f
C1187 VDD2.n48 VSUBS 0.035708f
C1188 VDD2.n49 VSUBS 0.035708f
C1189 VDD2.n50 VSUBS 0.019188f
C1190 VDD2.n51 VSUBS 0.020317f
C1191 VDD2.n52 VSUBS 0.045353f
C1192 VDD2.n53 VSUBS 0.045353f
C1193 VDD2.n54 VSUBS 0.020317f
C1194 VDD2.n55 VSUBS 0.019188f
C1195 VDD2.n56 VSUBS 0.035708f
C1196 VDD2.n57 VSUBS 0.09083f
C1197 VDD2.n58 VSUBS 0.019188f
C1198 VDD2.n59 VSUBS 0.020317f
C1199 VDD2.n60 VSUBS 0.09949f
C1200 VDD2.n61 VSUBS 0.091067f
C1201 VDD2.n62 VSUBS 4.08841f
C1202 VDD2.t3 VSUBS 0.163943f
C1203 VDD2.t5 VSUBS 0.163943f
C1204 VDD2.n63 VSUBS 1.10117f
C1205 VDD2.n64 VSUBS 1.06219f
C1206 VDD2.t1 VSUBS 0.163943f
C1207 VDD2.t4 VSUBS 0.163943f
C1208 VDD2.n65 VSUBS 1.13465f
C1209 VTAIL.t10 VSUBS 0.162153f
C1210 VTAIL.t11 VSUBS 0.162153f
C1211 VTAIL.n0 VSUBS 0.97469f
C1212 VTAIL.n1 VSUBS 1.17051f
C1213 VTAIL.n2 VSUBS 0.019888f
C1214 VTAIL.n3 VSUBS 0.044858f
C1215 VTAIL.n4 VSUBS 0.020095f
C1216 VTAIL.n5 VSUBS 0.035318f
C1217 VTAIL.n6 VSUBS 0.018978f
C1218 VTAIL.n7 VSUBS 0.044858f
C1219 VTAIL.n8 VSUBS 0.020095f
C1220 VTAIL.n9 VSUBS 0.776196f
C1221 VTAIL.n10 VSUBS 0.018978f
C1222 VTAIL.t4 VSUBS 0.096593f
C1223 VTAIL.n11 VSUBS 0.179829f
C1224 VTAIL.n12 VSUBS 0.03373f
C1225 VTAIL.n13 VSUBS 0.033643f
C1226 VTAIL.n14 VSUBS 0.044858f
C1227 VTAIL.n15 VSUBS 0.020095f
C1228 VTAIL.n16 VSUBS 0.018978f
C1229 VTAIL.n17 VSUBS 0.035318f
C1230 VTAIL.n18 VSUBS 0.035318f
C1231 VTAIL.n19 VSUBS 0.018978f
C1232 VTAIL.n20 VSUBS 0.020095f
C1233 VTAIL.n21 VSUBS 0.044858f
C1234 VTAIL.n22 VSUBS 0.044858f
C1235 VTAIL.n23 VSUBS 0.020095f
C1236 VTAIL.n24 VSUBS 0.018978f
C1237 VTAIL.n25 VSUBS 0.035318f
C1238 VTAIL.n26 VSUBS 0.089838f
C1239 VTAIL.n27 VSUBS 0.018978f
C1240 VTAIL.n28 VSUBS 0.020095f
C1241 VTAIL.n29 VSUBS 0.098404f
C1242 VTAIL.n30 VSUBS 0.065726f
C1243 VTAIL.n31 VSUBS 0.687036f
C1244 VTAIL.t7 VSUBS 0.162153f
C1245 VTAIL.t9 VSUBS 0.162153f
C1246 VTAIL.n32 VSUBS 0.97469f
C1247 VTAIL.n33 VSUBS 1.41062f
C1248 VTAIL.t1 VSUBS 0.162153f
C1249 VTAIL.t6 VSUBS 0.162153f
C1250 VTAIL.n34 VSUBS 0.97469f
C1251 VTAIL.n35 VSUBS 2.86064f
C1252 VTAIL.t12 VSUBS 0.162153f
C1253 VTAIL.t14 VSUBS 0.162153f
C1254 VTAIL.n36 VSUBS 0.974694f
C1255 VTAIL.n37 VSUBS 2.86063f
C1256 VTAIL.t19 VSUBS 0.162153f
C1257 VTAIL.t15 VSUBS 0.162153f
C1258 VTAIL.n38 VSUBS 0.974694f
C1259 VTAIL.n39 VSUBS 1.41062f
C1260 VTAIL.n40 VSUBS 0.019888f
C1261 VTAIL.n41 VSUBS 0.044858f
C1262 VTAIL.n42 VSUBS 0.020095f
C1263 VTAIL.n43 VSUBS 0.035318f
C1264 VTAIL.n44 VSUBS 0.018978f
C1265 VTAIL.n45 VSUBS 0.044858f
C1266 VTAIL.n46 VSUBS 0.020095f
C1267 VTAIL.n47 VSUBS 0.776196f
C1268 VTAIL.n48 VSUBS 0.018978f
C1269 VTAIL.t13 VSUBS 0.096593f
C1270 VTAIL.n49 VSUBS 0.179829f
C1271 VTAIL.n50 VSUBS 0.03373f
C1272 VTAIL.n51 VSUBS 0.033643f
C1273 VTAIL.n52 VSUBS 0.044858f
C1274 VTAIL.n53 VSUBS 0.020095f
C1275 VTAIL.n54 VSUBS 0.018978f
C1276 VTAIL.n55 VSUBS 0.035318f
C1277 VTAIL.n56 VSUBS 0.035318f
C1278 VTAIL.n57 VSUBS 0.018978f
C1279 VTAIL.n58 VSUBS 0.020095f
C1280 VTAIL.n59 VSUBS 0.044858f
C1281 VTAIL.n60 VSUBS 0.044858f
C1282 VTAIL.n61 VSUBS 0.020095f
C1283 VTAIL.n62 VSUBS 0.018978f
C1284 VTAIL.n63 VSUBS 0.035318f
C1285 VTAIL.n64 VSUBS 0.089838f
C1286 VTAIL.n65 VSUBS 0.018978f
C1287 VTAIL.n66 VSUBS 0.020095f
C1288 VTAIL.n67 VSUBS 0.098404f
C1289 VTAIL.n68 VSUBS 0.065726f
C1290 VTAIL.n69 VSUBS 0.687036f
C1291 VTAIL.t0 VSUBS 0.162153f
C1292 VTAIL.t5 VSUBS 0.162153f
C1293 VTAIL.n70 VSUBS 0.974694f
C1294 VTAIL.n71 VSUBS 1.26395f
C1295 VTAIL.t3 VSUBS 0.162153f
C1296 VTAIL.t8 VSUBS 0.162153f
C1297 VTAIL.n72 VSUBS 0.974694f
C1298 VTAIL.n73 VSUBS 1.41062f
C1299 VTAIL.n74 VSUBS 0.019888f
C1300 VTAIL.n75 VSUBS 0.044858f
C1301 VTAIL.n76 VSUBS 0.020095f
C1302 VTAIL.n77 VSUBS 0.035318f
C1303 VTAIL.n78 VSUBS 0.018978f
C1304 VTAIL.n79 VSUBS 0.044858f
C1305 VTAIL.n80 VSUBS 0.020095f
C1306 VTAIL.n81 VSUBS 0.776196f
C1307 VTAIL.n82 VSUBS 0.018978f
C1308 VTAIL.t2 VSUBS 0.096593f
C1309 VTAIL.n83 VSUBS 0.179829f
C1310 VTAIL.n84 VSUBS 0.03373f
C1311 VTAIL.n85 VSUBS 0.033643f
C1312 VTAIL.n86 VSUBS 0.044858f
C1313 VTAIL.n87 VSUBS 0.020095f
C1314 VTAIL.n88 VSUBS 0.018978f
C1315 VTAIL.n89 VSUBS 0.035318f
C1316 VTAIL.n90 VSUBS 0.035318f
C1317 VTAIL.n91 VSUBS 0.018978f
C1318 VTAIL.n92 VSUBS 0.020095f
C1319 VTAIL.n93 VSUBS 0.044858f
C1320 VTAIL.n94 VSUBS 0.044858f
C1321 VTAIL.n95 VSUBS 0.020095f
C1322 VTAIL.n96 VSUBS 0.018978f
C1323 VTAIL.n97 VSUBS 0.035318f
C1324 VTAIL.n98 VSUBS 0.089838f
C1325 VTAIL.n99 VSUBS 0.018978f
C1326 VTAIL.n100 VSUBS 0.020095f
C1327 VTAIL.n101 VSUBS 0.098404f
C1328 VTAIL.n102 VSUBS 0.065726f
C1329 VTAIL.n103 VSUBS 1.88345f
C1330 VTAIL.n104 VSUBS 0.019888f
C1331 VTAIL.n105 VSUBS 0.044858f
C1332 VTAIL.n106 VSUBS 0.020095f
C1333 VTAIL.n107 VSUBS 0.035318f
C1334 VTAIL.n108 VSUBS 0.018978f
C1335 VTAIL.n109 VSUBS 0.044858f
C1336 VTAIL.n110 VSUBS 0.020095f
C1337 VTAIL.n111 VSUBS 0.776196f
C1338 VTAIL.n112 VSUBS 0.018978f
C1339 VTAIL.t18 VSUBS 0.096593f
C1340 VTAIL.n113 VSUBS 0.179829f
C1341 VTAIL.n114 VSUBS 0.03373f
C1342 VTAIL.n115 VSUBS 0.033643f
C1343 VTAIL.n116 VSUBS 0.044858f
C1344 VTAIL.n117 VSUBS 0.020095f
C1345 VTAIL.n118 VSUBS 0.018978f
C1346 VTAIL.n119 VSUBS 0.035318f
C1347 VTAIL.n120 VSUBS 0.035318f
C1348 VTAIL.n121 VSUBS 0.018978f
C1349 VTAIL.n122 VSUBS 0.020095f
C1350 VTAIL.n123 VSUBS 0.044858f
C1351 VTAIL.n124 VSUBS 0.044858f
C1352 VTAIL.n125 VSUBS 0.020095f
C1353 VTAIL.n126 VSUBS 0.018978f
C1354 VTAIL.n127 VSUBS 0.035318f
C1355 VTAIL.n128 VSUBS 0.089838f
C1356 VTAIL.n129 VSUBS 0.018978f
C1357 VTAIL.n130 VSUBS 0.020095f
C1358 VTAIL.n131 VSUBS 0.098404f
C1359 VTAIL.n132 VSUBS 0.065726f
C1360 VTAIL.n133 VSUBS 1.88345f
C1361 VTAIL.t17 VSUBS 0.162153f
C1362 VTAIL.t16 VSUBS 0.162153f
C1363 VTAIL.n134 VSUBS 0.97469f
C1364 VTAIL.n135 VSUBS 1.1038f
C1365 VN.t0 VSUBS 1.79228f
C1366 VN.n0 VSUBS 0.786435f
C1367 VN.n1 VSUBS 0.03114f
C1368 VN.n2 VSUBS 0.055905f
C1369 VN.n3 VSUBS 0.03114f
C1370 VN.n4 VSUBS 0.053452f
C1371 VN.n5 VSUBS 0.03114f
C1372 VN.n6 VSUBS 0.060349f
C1373 VN.n7 VSUBS 0.03114f
C1374 VN.n8 VSUBS 0.058037f
C1375 VN.n9 VSUBS 0.03114f
C1376 VN.t1 VSUBS 1.79228f
C1377 VN.n10 VSUBS 0.062786f
C1378 VN.n11 VSUBS 0.03114f
C1379 VN.n12 VSUBS 0.058037f
C1380 VN.t7 VSUBS 2.21639f
C1381 VN.n13 VSUBS 0.738659f
C1382 VN.t3 VSUBS 1.79228f
C1383 VN.n14 VSUBS 0.763966f
C1384 VN.n15 VSUBS 0.033968f
C1385 VN.n16 VSUBS 0.395442f
C1386 VN.n17 VSUBS 0.03114f
C1387 VN.n18 VSUBS 0.03114f
C1388 VN.n19 VSUBS 0.058037f
C1389 VN.n20 VSUBS 0.060349f
C1390 VN.n21 VSUBS 0.02582f
C1391 VN.n22 VSUBS 0.03114f
C1392 VN.n23 VSUBS 0.03114f
C1393 VN.n24 VSUBS 0.03114f
C1394 VN.n25 VSUBS 0.058037f
C1395 VN.n26 VSUBS 0.058037f
C1396 VN.n27 VSUBS 0.691825f
C1397 VN.n28 VSUBS 0.03114f
C1398 VN.n29 VSUBS 0.03114f
C1399 VN.n30 VSUBS 0.03114f
C1400 VN.n31 VSUBS 0.058037f
C1401 VN.n32 VSUBS 0.062786f
C1402 VN.n33 VSUBS 0.02582f
C1403 VN.n34 VSUBS 0.03114f
C1404 VN.n35 VSUBS 0.03114f
C1405 VN.n36 VSUBS 0.03114f
C1406 VN.n37 VSUBS 0.058037f
C1407 VN.n38 VSUBS 0.058037f
C1408 VN.t2 VSUBS 1.79228f
C1409 VN.n39 VSUBS 0.662441f
C1410 VN.n40 VSUBS 0.033968f
C1411 VN.n41 VSUBS 0.03114f
C1412 VN.n42 VSUBS 0.03114f
C1413 VN.n43 VSUBS 0.03114f
C1414 VN.n44 VSUBS 0.058037f
C1415 VN.n45 VSUBS 0.061596f
C1416 VN.n46 VSUBS 0.031453f
C1417 VN.n47 VSUBS 0.03114f
C1418 VN.n48 VSUBS 0.03114f
C1419 VN.n49 VSUBS 0.03114f
C1420 VN.n50 VSUBS 0.058037f
C1421 VN.n51 VSUBS 0.058037f
C1422 VN.n52 VSUBS 0.038553f
C1423 VN.n53 VSUBS 0.050259f
C1424 VN.n54 VSUBS 0.089837f
C1425 VN.t9 VSUBS 1.79228f
C1426 VN.n55 VSUBS 0.786435f
C1427 VN.n56 VSUBS 0.03114f
C1428 VN.n57 VSUBS 0.055905f
C1429 VN.n58 VSUBS 0.03114f
C1430 VN.n59 VSUBS 0.053452f
C1431 VN.n60 VSUBS 0.03114f
C1432 VN.t6 VSUBS 1.79228f
C1433 VN.n61 VSUBS 0.662441f
C1434 VN.n62 VSUBS 0.060349f
C1435 VN.n63 VSUBS 0.03114f
C1436 VN.n64 VSUBS 0.058037f
C1437 VN.n65 VSUBS 0.03114f
C1438 VN.t4 VSUBS 1.79228f
C1439 VN.n66 VSUBS 0.062786f
C1440 VN.n67 VSUBS 0.03114f
C1441 VN.n68 VSUBS 0.058037f
C1442 VN.t5 VSUBS 2.21639f
C1443 VN.n69 VSUBS 0.738659f
C1444 VN.t8 VSUBS 1.79228f
C1445 VN.n70 VSUBS 0.763966f
C1446 VN.n71 VSUBS 0.033968f
C1447 VN.n72 VSUBS 0.395442f
C1448 VN.n73 VSUBS 0.03114f
C1449 VN.n74 VSUBS 0.03114f
C1450 VN.n75 VSUBS 0.058037f
C1451 VN.n76 VSUBS 0.060349f
C1452 VN.n77 VSUBS 0.02582f
C1453 VN.n78 VSUBS 0.03114f
C1454 VN.n79 VSUBS 0.03114f
C1455 VN.n80 VSUBS 0.03114f
C1456 VN.n81 VSUBS 0.058037f
C1457 VN.n82 VSUBS 0.058037f
C1458 VN.n83 VSUBS 0.691825f
C1459 VN.n84 VSUBS 0.03114f
C1460 VN.n85 VSUBS 0.03114f
C1461 VN.n86 VSUBS 0.03114f
C1462 VN.n87 VSUBS 0.058037f
C1463 VN.n88 VSUBS 0.062786f
C1464 VN.n89 VSUBS 0.02582f
C1465 VN.n90 VSUBS 0.03114f
C1466 VN.n91 VSUBS 0.03114f
C1467 VN.n92 VSUBS 0.03114f
C1468 VN.n93 VSUBS 0.058037f
C1469 VN.n94 VSUBS 0.058037f
C1470 VN.n95 VSUBS 0.033968f
C1471 VN.n96 VSUBS 0.03114f
C1472 VN.n97 VSUBS 0.03114f
C1473 VN.n98 VSUBS 0.03114f
C1474 VN.n99 VSUBS 0.058037f
C1475 VN.n100 VSUBS 0.061596f
C1476 VN.n101 VSUBS 0.031453f
C1477 VN.n102 VSUBS 0.03114f
C1478 VN.n103 VSUBS 0.03114f
C1479 VN.n104 VSUBS 0.03114f
C1480 VN.n105 VSUBS 0.058037f
C1481 VN.n106 VSUBS 0.058037f
C1482 VN.n107 VSUBS 0.038553f
C1483 VN.n108 VSUBS 0.050259f
C1484 VN.n109 VSUBS 2.04427f
.ends

