* NGSPICE file created from diff_pair_sample_1223.ext - technology: sky130A

.subckt diff_pair_sample_1223 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t15 w_n3334_n3172# sky130_fd_pr__pfet_01v8 ad=1.8183 pd=11.35 as=4.2978 ps=22.82 w=11.02 l=1.64
X1 VTAIL.t19 VP.t1 VDD1.t8 w_n3334_n3172# sky130_fd_pr__pfet_01v8 ad=1.8183 pd=11.35 as=1.8183 ps=11.35 w=11.02 l=1.64
X2 VTAIL.t4 VN.t0 VDD2.t9 w_n3334_n3172# sky130_fd_pr__pfet_01v8 ad=1.8183 pd=11.35 as=1.8183 ps=11.35 w=11.02 l=1.64
X3 B.t11 B.t9 B.t10 w_n3334_n3172# sky130_fd_pr__pfet_01v8 ad=4.2978 pd=22.82 as=0 ps=0 w=11.02 l=1.64
X4 VTAIL.t5 VN.t1 VDD2.t8 w_n3334_n3172# sky130_fd_pr__pfet_01v8 ad=1.8183 pd=11.35 as=1.8183 ps=11.35 w=11.02 l=1.64
X5 VTAIL.t12 VP.t2 VDD1.t7 w_n3334_n3172# sky130_fd_pr__pfet_01v8 ad=1.8183 pd=11.35 as=1.8183 ps=11.35 w=11.02 l=1.64
X6 B.t8 B.t6 B.t7 w_n3334_n3172# sky130_fd_pr__pfet_01v8 ad=4.2978 pd=22.82 as=0 ps=0 w=11.02 l=1.64
X7 VDD1.t6 VP.t3 VTAIL.t18 w_n3334_n3172# sky130_fd_pr__pfet_01v8 ad=4.2978 pd=22.82 as=1.8183 ps=11.35 w=11.02 l=1.64
X8 VTAIL.t6 VN.t2 VDD2.t7 w_n3334_n3172# sky130_fd_pr__pfet_01v8 ad=1.8183 pd=11.35 as=1.8183 ps=11.35 w=11.02 l=1.64
X9 VTAIL.t13 VP.t4 VDD1.t5 w_n3334_n3172# sky130_fd_pr__pfet_01v8 ad=1.8183 pd=11.35 as=1.8183 ps=11.35 w=11.02 l=1.64
X10 VDD2.t6 VN.t3 VTAIL.t7 w_n3334_n3172# sky130_fd_pr__pfet_01v8 ad=1.8183 pd=11.35 as=4.2978 ps=22.82 w=11.02 l=1.64
X11 VTAIL.t14 VP.t5 VDD1.t4 w_n3334_n3172# sky130_fd_pr__pfet_01v8 ad=1.8183 pd=11.35 as=1.8183 ps=11.35 w=11.02 l=1.64
X12 B.t5 B.t3 B.t4 w_n3334_n3172# sky130_fd_pr__pfet_01v8 ad=4.2978 pd=22.82 as=0 ps=0 w=11.02 l=1.64
X13 VDD2.t5 VN.t4 VTAIL.t9 w_n3334_n3172# sky130_fd_pr__pfet_01v8 ad=4.2978 pd=22.82 as=1.8183 ps=11.35 w=11.02 l=1.64
X14 B.t2 B.t0 B.t1 w_n3334_n3172# sky130_fd_pr__pfet_01v8 ad=4.2978 pd=22.82 as=0 ps=0 w=11.02 l=1.64
X15 VDD1.t3 VP.t6 VTAIL.t11 w_n3334_n3172# sky130_fd_pr__pfet_01v8 ad=1.8183 pd=11.35 as=4.2978 ps=22.82 w=11.02 l=1.64
X16 VDD1.t2 VP.t7 VTAIL.t16 w_n3334_n3172# sky130_fd_pr__pfet_01v8 ad=1.8183 pd=11.35 as=1.8183 ps=11.35 w=11.02 l=1.64
X17 VTAIL.t2 VN.t5 VDD2.t4 w_n3334_n3172# sky130_fd_pr__pfet_01v8 ad=1.8183 pd=11.35 as=1.8183 ps=11.35 w=11.02 l=1.64
X18 VDD2.t3 VN.t6 VTAIL.t0 w_n3334_n3172# sky130_fd_pr__pfet_01v8 ad=4.2978 pd=22.82 as=1.8183 ps=11.35 w=11.02 l=1.64
X19 VDD1.t1 VP.t8 VTAIL.t17 w_n3334_n3172# sky130_fd_pr__pfet_01v8 ad=1.8183 pd=11.35 as=1.8183 ps=11.35 w=11.02 l=1.64
X20 VDD2.t2 VN.t7 VTAIL.t8 w_n3334_n3172# sky130_fd_pr__pfet_01v8 ad=1.8183 pd=11.35 as=4.2978 ps=22.82 w=11.02 l=1.64
X21 VDD2.t1 VN.t8 VTAIL.t1 w_n3334_n3172# sky130_fd_pr__pfet_01v8 ad=1.8183 pd=11.35 as=1.8183 ps=11.35 w=11.02 l=1.64
X22 VDD2.t0 VN.t9 VTAIL.t3 w_n3334_n3172# sky130_fd_pr__pfet_01v8 ad=1.8183 pd=11.35 as=1.8183 ps=11.35 w=11.02 l=1.64
X23 VDD1.t0 VP.t9 VTAIL.t10 w_n3334_n3172# sky130_fd_pr__pfet_01v8 ad=4.2978 pd=22.82 as=1.8183 ps=11.35 w=11.02 l=1.64
R0 VP.n14 VP.t3 195.387
R1 VP.n39 VP.n38 176.548
R2 VP.n68 VP.n67 176.548
R3 VP.n37 VP.n36 176.548
R4 VP.n39 VP.t9 161.94
R5 VP.n46 VP.t2 161.94
R6 VP.n53 VP.t8 161.94
R7 VP.n60 VP.t4 161.94
R8 VP.n67 VP.t6 161.94
R9 VP.n36 VP.t0 161.94
R10 VP.n29 VP.t5 161.94
R11 VP.n22 VP.t7 161.94
R12 VP.n15 VP.t1 161.94
R13 VP.n17 VP.n16 161.3
R14 VP.n18 VP.n13 161.3
R15 VP.n20 VP.n19 161.3
R16 VP.n21 VP.n12 161.3
R17 VP.n24 VP.n23 161.3
R18 VP.n25 VP.n11 161.3
R19 VP.n27 VP.n26 161.3
R20 VP.n28 VP.n10 161.3
R21 VP.n31 VP.n30 161.3
R22 VP.n32 VP.n9 161.3
R23 VP.n34 VP.n33 161.3
R24 VP.n35 VP.n8 161.3
R25 VP.n66 VP.n0 161.3
R26 VP.n65 VP.n64 161.3
R27 VP.n63 VP.n1 161.3
R28 VP.n62 VP.n61 161.3
R29 VP.n59 VP.n2 161.3
R30 VP.n58 VP.n57 161.3
R31 VP.n56 VP.n3 161.3
R32 VP.n55 VP.n54 161.3
R33 VP.n52 VP.n4 161.3
R34 VP.n51 VP.n50 161.3
R35 VP.n49 VP.n5 161.3
R36 VP.n48 VP.n47 161.3
R37 VP.n45 VP.n6 161.3
R38 VP.n44 VP.n43 161.3
R39 VP.n42 VP.n7 161.3
R40 VP.n41 VP.n40 161.3
R41 VP.n44 VP.n7 56.5617
R42 VP.n65 VP.n1 56.5617
R43 VP.n34 VP.n9 56.5617
R44 VP.n51 VP.n5 56.5617
R45 VP.n58 VP.n3 56.5617
R46 VP.n27 VP.n11 56.5617
R47 VP.n20 VP.n13 56.5617
R48 VP.n15 VP.n14 55.694
R49 VP.n38 VP.n37 47.1028
R50 VP.n40 VP.n7 24.5923
R51 VP.n45 VP.n44 24.5923
R52 VP.n47 VP.n5 24.5923
R53 VP.n52 VP.n51 24.5923
R54 VP.n54 VP.n3 24.5923
R55 VP.n59 VP.n58 24.5923
R56 VP.n61 VP.n1 24.5923
R57 VP.n66 VP.n65 24.5923
R58 VP.n35 VP.n34 24.5923
R59 VP.n28 VP.n27 24.5923
R60 VP.n30 VP.n9 24.5923
R61 VP.n21 VP.n20 24.5923
R62 VP.n23 VP.n11 24.5923
R63 VP.n16 VP.n13 24.5923
R64 VP.n17 VP.n14 17.8292
R65 VP.n46 VP.n45 13.7719
R66 VP.n61 VP.n60 13.7719
R67 VP.n30 VP.n29 13.7719
R68 VP.n53 VP.n52 12.2964
R69 VP.n54 VP.n53 12.2964
R70 VP.n22 VP.n21 12.2964
R71 VP.n23 VP.n22 12.2964
R72 VP.n47 VP.n46 10.8209
R73 VP.n60 VP.n59 10.8209
R74 VP.n29 VP.n28 10.8209
R75 VP.n16 VP.n15 10.8209
R76 VP.n40 VP.n39 9.3454
R77 VP.n67 VP.n66 9.3454
R78 VP.n36 VP.n35 9.3454
R79 VP.n18 VP.n17 0.189894
R80 VP.n19 VP.n18 0.189894
R81 VP.n19 VP.n12 0.189894
R82 VP.n24 VP.n12 0.189894
R83 VP.n25 VP.n24 0.189894
R84 VP.n26 VP.n25 0.189894
R85 VP.n26 VP.n10 0.189894
R86 VP.n31 VP.n10 0.189894
R87 VP.n32 VP.n31 0.189894
R88 VP.n33 VP.n32 0.189894
R89 VP.n33 VP.n8 0.189894
R90 VP.n37 VP.n8 0.189894
R91 VP.n41 VP.n38 0.189894
R92 VP.n42 VP.n41 0.189894
R93 VP.n43 VP.n42 0.189894
R94 VP.n43 VP.n6 0.189894
R95 VP.n48 VP.n6 0.189894
R96 VP.n49 VP.n48 0.189894
R97 VP.n50 VP.n49 0.189894
R98 VP.n50 VP.n4 0.189894
R99 VP.n55 VP.n4 0.189894
R100 VP.n56 VP.n55 0.189894
R101 VP.n57 VP.n56 0.189894
R102 VP.n57 VP.n2 0.189894
R103 VP.n62 VP.n2 0.189894
R104 VP.n63 VP.n62 0.189894
R105 VP.n64 VP.n63 0.189894
R106 VP.n64 VP.n0 0.189894
R107 VP.n68 VP.n0 0.189894
R108 VP VP.n68 0.0516364
R109 VTAIL.n11 VTAIL.t7 61.188
R110 VTAIL.n17 VTAIL.t8 61.1878
R111 VTAIL.n2 VTAIL.t11 61.1878
R112 VTAIL.n16 VTAIL.t15 61.1878
R113 VTAIL.n15 VTAIL.n14 58.2384
R114 VTAIL.n13 VTAIL.n12 58.2384
R115 VTAIL.n10 VTAIL.n9 58.2384
R116 VTAIL.n8 VTAIL.n7 58.2384
R117 VTAIL.n19 VTAIL.n18 58.2381
R118 VTAIL.n1 VTAIL.n0 58.2381
R119 VTAIL.n4 VTAIL.n3 58.2381
R120 VTAIL.n6 VTAIL.n5 58.2381
R121 VTAIL.n8 VTAIL.n6 25.2634
R122 VTAIL.n17 VTAIL.n16 23.5652
R123 VTAIL.n18 VTAIL.t1 2.95014
R124 VTAIL.n18 VTAIL.t6 2.95014
R125 VTAIL.n0 VTAIL.t0 2.95014
R126 VTAIL.n0 VTAIL.t5 2.95014
R127 VTAIL.n3 VTAIL.t17 2.95014
R128 VTAIL.n3 VTAIL.t13 2.95014
R129 VTAIL.n5 VTAIL.t10 2.95014
R130 VTAIL.n5 VTAIL.t12 2.95014
R131 VTAIL.n14 VTAIL.t16 2.95014
R132 VTAIL.n14 VTAIL.t14 2.95014
R133 VTAIL.n12 VTAIL.t18 2.95014
R134 VTAIL.n12 VTAIL.t19 2.95014
R135 VTAIL.n9 VTAIL.t3 2.95014
R136 VTAIL.n9 VTAIL.t4 2.95014
R137 VTAIL.n7 VTAIL.t9 2.95014
R138 VTAIL.n7 VTAIL.t2 2.95014
R139 VTAIL.n10 VTAIL.n8 1.69878
R140 VTAIL.n11 VTAIL.n10 1.69878
R141 VTAIL.n15 VTAIL.n13 1.69878
R142 VTAIL.n16 VTAIL.n15 1.69878
R143 VTAIL.n6 VTAIL.n4 1.69878
R144 VTAIL.n4 VTAIL.n2 1.69878
R145 VTAIL.n19 VTAIL.n17 1.69878
R146 VTAIL VTAIL.n1 1.3324
R147 VTAIL.n13 VTAIL.n11 1.31947
R148 VTAIL.n2 VTAIL.n1 1.31947
R149 VTAIL VTAIL.n19 0.366879
R150 VDD1.n1 VDD1.t6 79.565
R151 VDD1.n3 VDD1.t0 79.5649
R152 VDD1.n5 VDD1.n4 76.1353
R153 VDD1.n1 VDD1.n0 74.9172
R154 VDD1.n7 VDD1.n6 74.917
R155 VDD1.n3 VDD1.n2 74.9169
R156 VDD1.n7 VDD1.n5 42.7143
R157 VDD1.n6 VDD1.t4 2.95014
R158 VDD1.n6 VDD1.t9 2.95014
R159 VDD1.n0 VDD1.t8 2.95014
R160 VDD1.n0 VDD1.t2 2.95014
R161 VDD1.n4 VDD1.t5 2.95014
R162 VDD1.n4 VDD1.t3 2.95014
R163 VDD1.n2 VDD1.t7 2.95014
R164 VDD1.n2 VDD1.t1 2.95014
R165 VDD1 VDD1.n7 1.21602
R166 VDD1 VDD1.n1 0.483259
R167 VDD1.n5 VDD1.n3 0.369723
R168 VN.n6 VN.t6 195.387
R169 VN.n36 VN.t3 195.387
R170 VN.n29 VN.n28 176.548
R171 VN.n59 VN.n58 176.548
R172 VN.n7 VN.t1 161.94
R173 VN.n14 VN.t8 161.94
R174 VN.n21 VN.t2 161.94
R175 VN.n28 VN.t7 161.94
R176 VN.n37 VN.t0 161.94
R177 VN.n44 VN.t9 161.94
R178 VN.n51 VN.t5 161.94
R179 VN.n58 VN.t4 161.94
R180 VN.n57 VN.n30 161.3
R181 VN.n56 VN.n55 161.3
R182 VN.n54 VN.n31 161.3
R183 VN.n53 VN.n52 161.3
R184 VN.n50 VN.n32 161.3
R185 VN.n49 VN.n48 161.3
R186 VN.n47 VN.n33 161.3
R187 VN.n46 VN.n45 161.3
R188 VN.n43 VN.n34 161.3
R189 VN.n42 VN.n41 161.3
R190 VN.n40 VN.n35 161.3
R191 VN.n39 VN.n38 161.3
R192 VN.n27 VN.n0 161.3
R193 VN.n26 VN.n25 161.3
R194 VN.n24 VN.n1 161.3
R195 VN.n23 VN.n22 161.3
R196 VN.n20 VN.n2 161.3
R197 VN.n19 VN.n18 161.3
R198 VN.n17 VN.n3 161.3
R199 VN.n16 VN.n15 161.3
R200 VN.n13 VN.n4 161.3
R201 VN.n12 VN.n11 161.3
R202 VN.n10 VN.n5 161.3
R203 VN.n9 VN.n8 161.3
R204 VN.n26 VN.n1 56.5617
R205 VN.n56 VN.n31 56.5617
R206 VN.n12 VN.n5 56.5617
R207 VN.n19 VN.n3 56.5617
R208 VN.n42 VN.n35 56.5617
R209 VN.n49 VN.n33 56.5617
R210 VN.n7 VN.n6 55.694
R211 VN.n37 VN.n36 55.694
R212 VN VN.n59 47.4835
R213 VN.n8 VN.n5 24.5923
R214 VN.n13 VN.n12 24.5923
R215 VN.n15 VN.n3 24.5923
R216 VN.n20 VN.n19 24.5923
R217 VN.n22 VN.n1 24.5923
R218 VN.n27 VN.n26 24.5923
R219 VN.n38 VN.n35 24.5923
R220 VN.n45 VN.n33 24.5923
R221 VN.n43 VN.n42 24.5923
R222 VN.n52 VN.n31 24.5923
R223 VN.n50 VN.n49 24.5923
R224 VN.n57 VN.n56 24.5923
R225 VN.n39 VN.n36 17.8292
R226 VN.n9 VN.n6 17.8292
R227 VN.n22 VN.n21 13.7719
R228 VN.n52 VN.n51 13.7719
R229 VN.n14 VN.n13 12.2964
R230 VN.n15 VN.n14 12.2964
R231 VN.n45 VN.n44 12.2964
R232 VN.n44 VN.n43 12.2964
R233 VN.n8 VN.n7 10.8209
R234 VN.n21 VN.n20 10.8209
R235 VN.n38 VN.n37 10.8209
R236 VN.n51 VN.n50 10.8209
R237 VN.n28 VN.n27 9.3454
R238 VN.n58 VN.n57 9.3454
R239 VN.n59 VN.n30 0.189894
R240 VN.n55 VN.n30 0.189894
R241 VN.n55 VN.n54 0.189894
R242 VN.n54 VN.n53 0.189894
R243 VN.n53 VN.n32 0.189894
R244 VN.n48 VN.n32 0.189894
R245 VN.n48 VN.n47 0.189894
R246 VN.n47 VN.n46 0.189894
R247 VN.n46 VN.n34 0.189894
R248 VN.n41 VN.n34 0.189894
R249 VN.n41 VN.n40 0.189894
R250 VN.n40 VN.n39 0.189894
R251 VN.n10 VN.n9 0.189894
R252 VN.n11 VN.n10 0.189894
R253 VN.n11 VN.n4 0.189894
R254 VN.n16 VN.n4 0.189894
R255 VN.n17 VN.n16 0.189894
R256 VN.n18 VN.n17 0.189894
R257 VN.n18 VN.n2 0.189894
R258 VN.n23 VN.n2 0.189894
R259 VN.n24 VN.n23 0.189894
R260 VN.n25 VN.n24 0.189894
R261 VN.n25 VN.n0 0.189894
R262 VN.n29 VN.n0 0.189894
R263 VN VN.n29 0.0516364
R264 VDD2.n1 VDD2.t3 79.5649
R265 VDD2.n4 VDD2.t5 77.8667
R266 VDD2.n3 VDD2.n2 76.1353
R267 VDD2 VDD2.n7 76.1325
R268 VDD2.n6 VDD2.n5 74.9172
R269 VDD2.n1 VDD2.n0 74.9169
R270 VDD2.n4 VDD2.n3 41.2821
R271 VDD2.n7 VDD2.t9 2.95014
R272 VDD2.n7 VDD2.t6 2.95014
R273 VDD2.n5 VDD2.t4 2.95014
R274 VDD2.n5 VDD2.t0 2.95014
R275 VDD2.n2 VDD2.t7 2.95014
R276 VDD2.n2 VDD2.t2 2.95014
R277 VDD2.n0 VDD2.t8 2.95014
R278 VDD2.n0 VDD2.t1 2.95014
R279 VDD2.n6 VDD2.n4 1.69878
R280 VDD2 VDD2.n6 0.483259
R281 VDD2.n3 VDD2.n1 0.369723
R282 B.n510 B.n509 585
R283 B.n511 B.n70 585
R284 B.n513 B.n512 585
R285 B.n514 B.n69 585
R286 B.n516 B.n515 585
R287 B.n517 B.n68 585
R288 B.n519 B.n518 585
R289 B.n520 B.n67 585
R290 B.n522 B.n521 585
R291 B.n523 B.n66 585
R292 B.n525 B.n524 585
R293 B.n526 B.n65 585
R294 B.n528 B.n527 585
R295 B.n529 B.n64 585
R296 B.n531 B.n530 585
R297 B.n532 B.n63 585
R298 B.n534 B.n533 585
R299 B.n535 B.n62 585
R300 B.n537 B.n536 585
R301 B.n538 B.n61 585
R302 B.n540 B.n539 585
R303 B.n541 B.n60 585
R304 B.n543 B.n542 585
R305 B.n544 B.n59 585
R306 B.n546 B.n545 585
R307 B.n547 B.n58 585
R308 B.n549 B.n548 585
R309 B.n550 B.n57 585
R310 B.n552 B.n551 585
R311 B.n553 B.n56 585
R312 B.n555 B.n554 585
R313 B.n556 B.n55 585
R314 B.n558 B.n557 585
R315 B.n559 B.n54 585
R316 B.n561 B.n560 585
R317 B.n562 B.n53 585
R318 B.n564 B.n563 585
R319 B.n565 B.n52 585
R320 B.n567 B.n566 585
R321 B.n569 B.n49 585
R322 B.n571 B.n570 585
R323 B.n572 B.n48 585
R324 B.n574 B.n573 585
R325 B.n575 B.n47 585
R326 B.n577 B.n576 585
R327 B.n578 B.n46 585
R328 B.n580 B.n579 585
R329 B.n581 B.n43 585
R330 B.n584 B.n583 585
R331 B.n585 B.n42 585
R332 B.n587 B.n586 585
R333 B.n588 B.n41 585
R334 B.n590 B.n589 585
R335 B.n591 B.n40 585
R336 B.n593 B.n592 585
R337 B.n594 B.n39 585
R338 B.n596 B.n595 585
R339 B.n597 B.n38 585
R340 B.n599 B.n598 585
R341 B.n600 B.n37 585
R342 B.n602 B.n601 585
R343 B.n603 B.n36 585
R344 B.n605 B.n604 585
R345 B.n606 B.n35 585
R346 B.n608 B.n607 585
R347 B.n609 B.n34 585
R348 B.n611 B.n610 585
R349 B.n612 B.n33 585
R350 B.n614 B.n613 585
R351 B.n615 B.n32 585
R352 B.n617 B.n616 585
R353 B.n618 B.n31 585
R354 B.n620 B.n619 585
R355 B.n621 B.n30 585
R356 B.n623 B.n622 585
R357 B.n624 B.n29 585
R358 B.n626 B.n625 585
R359 B.n627 B.n28 585
R360 B.n629 B.n628 585
R361 B.n630 B.n27 585
R362 B.n632 B.n631 585
R363 B.n633 B.n26 585
R364 B.n635 B.n634 585
R365 B.n636 B.n25 585
R366 B.n638 B.n637 585
R367 B.n639 B.n24 585
R368 B.n641 B.n640 585
R369 B.n508 B.n71 585
R370 B.n507 B.n506 585
R371 B.n505 B.n72 585
R372 B.n504 B.n503 585
R373 B.n502 B.n73 585
R374 B.n501 B.n500 585
R375 B.n499 B.n74 585
R376 B.n498 B.n497 585
R377 B.n496 B.n75 585
R378 B.n495 B.n494 585
R379 B.n493 B.n76 585
R380 B.n492 B.n491 585
R381 B.n490 B.n77 585
R382 B.n489 B.n488 585
R383 B.n487 B.n78 585
R384 B.n486 B.n485 585
R385 B.n484 B.n79 585
R386 B.n483 B.n482 585
R387 B.n481 B.n80 585
R388 B.n480 B.n479 585
R389 B.n478 B.n81 585
R390 B.n477 B.n476 585
R391 B.n475 B.n82 585
R392 B.n474 B.n473 585
R393 B.n472 B.n83 585
R394 B.n471 B.n470 585
R395 B.n469 B.n84 585
R396 B.n468 B.n467 585
R397 B.n466 B.n85 585
R398 B.n465 B.n464 585
R399 B.n463 B.n86 585
R400 B.n462 B.n461 585
R401 B.n460 B.n87 585
R402 B.n459 B.n458 585
R403 B.n457 B.n88 585
R404 B.n456 B.n455 585
R405 B.n454 B.n89 585
R406 B.n453 B.n452 585
R407 B.n451 B.n90 585
R408 B.n450 B.n449 585
R409 B.n448 B.n91 585
R410 B.n447 B.n446 585
R411 B.n445 B.n92 585
R412 B.n444 B.n443 585
R413 B.n442 B.n93 585
R414 B.n441 B.n440 585
R415 B.n439 B.n94 585
R416 B.n438 B.n437 585
R417 B.n436 B.n95 585
R418 B.n435 B.n434 585
R419 B.n433 B.n96 585
R420 B.n432 B.n431 585
R421 B.n430 B.n97 585
R422 B.n429 B.n428 585
R423 B.n427 B.n98 585
R424 B.n426 B.n425 585
R425 B.n424 B.n99 585
R426 B.n423 B.n422 585
R427 B.n421 B.n100 585
R428 B.n420 B.n419 585
R429 B.n418 B.n101 585
R430 B.n417 B.n416 585
R431 B.n415 B.n102 585
R432 B.n414 B.n413 585
R433 B.n412 B.n103 585
R434 B.n411 B.n410 585
R435 B.n409 B.n104 585
R436 B.n408 B.n407 585
R437 B.n406 B.n105 585
R438 B.n405 B.n404 585
R439 B.n403 B.n106 585
R440 B.n402 B.n401 585
R441 B.n400 B.n107 585
R442 B.n399 B.n398 585
R443 B.n397 B.n108 585
R444 B.n396 B.n395 585
R445 B.n394 B.n109 585
R446 B.n393 B.n392 585
R447 B.n391 B.n110 585
R448 B.n390 B.n389 585
R449 B.n388 B.n111 585
R450 B.n387 B.n386 585
R451 B.n385 B.n112 585
R452 B.n384 B.n383 585
R453 B.n382 B.n113 585
R454 B.n381 B.n380 585
R455 B.n379 B.n114 585
R456 B.n247 B.n162 585
R457 B.n249 B.n248 585
R458 B.n250 B.n161 585
R459 B.n252 B.n251 585
R460 B.n253 B.n160 585
R461 B.n255 B.n254 585
R462 B.n256 B.n159 585
R463 B.n258 B.n257 585
R464 B.n259 B.n158 585
R465 B.n261 B.n260 585
R466 B.n262 B.n157 585
R467 B.n264 B.n263 585
R468 B.n265 B.n156 585
R469 B.n267 B.n266 585
R470 B.n268 B.n155 585
R471 B.n270 B.n269 585
R472 B.n271 B.n154 585
R473 B.n273 B.n272 585
R474 B.n274 B.n153 585
R475 B.n276 B.n275 585
R476 B.n277 B.n152 585
R477 B.n279 B.n278 585
R478 B.n280 B.n151 585
R479 B.n282 B.n281 585
R480 B.n283 B.n150 585
R481 B.n285 B.n284 585
R482 B.n286 B.n149 585
R483 B.n288 B.n287 585
R484 B.n289 B.n148 585
R485 B.n291 B.n290 585
R486 B.n292 B.n147 585
R487 B.n294 B.n293 585
R488 B.n295 B.n146 585
R489 B.n297 B.n296 585
R490 B.n298 B.n145 585
R491 B.n300 B.n299 585
R492 B.n301 B.n144 585
R493 B.n303 B.n302 585
R494 B.n304 B.n141 585
R495 B.n307 B.n306 585
R496 B.n308 B.n140 585
R497 B.n310 B.n309 585
R498 B.n311 B.n139 585
R499 B.n313 B.n312 585
R500 B.n314 B.n138 585
R501 B.n316 B.n315 585
R502 B.n317 B.n137 585
R503 B.n319 B.n318 585
R504 B.n321 B.n320 585
R505 B.n322 B.n133 585
R506 B.n324 B.n323 585
R507 B.n325 B.n132 585
R508 B.n327 B.n326 585
R509 B.n328 B.n131 585
R510 B.n330 B.n329 585
R511 B.n331 B.n130 585
R512 B.n333 B.n332 585
R513 B.n334 B.n129 585
R514 B.n336 B.n335 585
R515 B.n337 B.n128 585
R516 B.n339 B.n338 585
R517 B.n340 B.n127 585
R518 B.n342 B.n341 585
R519 B.n343 B.n126 585
R520 B.n345 B.n344 585
R521 B.n346 B.n125 585
R522 B.n348 B.n347 585
R523 B.n349 B.n124 585
R524 B.n351 B.n350 585
R525 B.n352 B.n123 585
R526 B.n354 B.n353 585
R527 B.n355 B.n122 585
R528 B.n357 B.n356 585
R529 B.n358 B.n121 585
R530 B.n360 B.n359 585
R531 B.n361 B.n120 585
R532 B.n363 B.n362 585
R533 B.n364 B.n119 585
R534 B.n366 B.n365 585
R535 B.n367 B.n118 585
R536 B.n369 B.n368 585
R537 B.n370 B.n117 585
R538 B.n372 B.n371 585
R539 B.n373 B.n116 585
R540 B.n375 B.n374 585
R541 B.n376 B.n115 585
R542 B.n378 B.n377 585
R543 B.n246 B.n245 585
R544 B.n244 B.n163 585
R545 B.n243 B.n242 585
R546 B.n241 B.n164 585
R547 B.n240 B.n239 585
R548 B.n238 B.n165 585
R549 B.n237 B.n236 585
R550 B.n235 B.n166 585
R551 B.n234 B.n233 585
R552 B.n232 B.n167 585
R553 B.n231 B.n230 585
R554 B.n229 B.n168 585
R555 B.n228 B.n227 585
R556 B.n226 B.n169 585
R557 B.n225 B.n224 585
R558 B.n223 B.n170 585
R559 B.n222 B.n221 585
R560 B.n220 B.n171 585
R561 B.n219 B.n218 585
R562 B.n217 B.n172 585
R563 B.n216 B.n215 585
R564 B.n214 B.n173 585
R565 B.n213 B.n212 585
R566 B.n211 B.n174 585
R567 B.n210 B.n209 585
R568 B.n208 B.n175 585
R569 B.n207 B.n206 585
R570 B.n205 B.n176 585
R571 B.n204 B.n203 585
R572 B.n202 B.n177 585
R573 B.n201 B.n200 585
R574 B.n199 B.n178 585
R575 B.n198 B.n197 585
R576 B.n196 B.n179 585
R577 B.n195 B.n194 585
R578 B.n193 B.n180 585
R579 B.n192 B.n191 585
R580 B.n190 B.n181 585
R581 B.n189 B.n188 585
R582 B.n187 B.n182 585
R583 B.n186 B.n185 585
R584 B.n184 B.n183 585
R585 B.n2 B.n0 585
R586 B.n705 B.n1 585
R587 B.n704 B.n703 585
R588 B.n702 B.n3 585
R589 B.n701 B.n700 585
R590 B.n699 B.n4 585
R591 B.n698 B.n697 585
R592 B.n696 B.n5 585
R593 B.n695 B.n694 585
R594 B.n693 B.n6 585
R595 B.n692 B.n691 585
R596 B.n690 B.n7 585
R597 B.n689 B.n688 585
R598 B.n687 B.n8 585
R599 B.n686 B.n685 585
R600 B.n684 B.n9 585
R601 B.n683 B.n682 585
R602 B.n681 B.n10 585
R603 B.n680 B.n679 585
R604 B.n678 B.n11 585
R605 B.n677 B.n676 585
R606 B.n675 B.n12 585
R607 B.n674 B.n673 585
R608 B.n672 B.n13 585
R609 B.n671 B.n670 585
R610 B.n669 B.n14 585
R611 B.n668 B.n667 585
R612 B.n666 B.n15 585
R613 B.n665 B.n664 585
R614 B.n663 B.n16 585
R615 B.n662 B.n661 585
R616 B.n660 B.n17 585
R617 B.n659 B.n658 585
R618 B.n657 B.n18 585
R619 B.n656 B.n655 585
R620 B.n654 B.n19 585
R621 B.n653 B.n652 585
R622 B.n651 B.n20 585
R623 B.n650 B.n649 585
R624 B.n648 B.n21 585
R625 B.n647 B.n646 585
R626 B.n645 B.n22 585
R627 B.n644 B.n643 585
R628 B.n642 B.n23 585
R629 B.n707 B.n706 585
R630 B.n247 B.n246 482.89
R631 B.n640 B.n23 482.89
R632 B.n379 B.n378 482.89
R633 B.n510 B.n71 482.89
R634 B.n134 B.t9 367.865
R635 B.n142 B.t0 367.865
R636 B.n44 B.t6 367.865
R637 B.n50 B.t3 367.865
R638 B.n246 B.n163 163.367
R639 B.n242 B.n163 163.367
R640 B.n242 B.n241 163.367
R641 B.n241 B.n240 163.367
R642 B.n240 B.n165 163.367
R643 B.n236 B.n165 163.367
R644 B.n236 B.n235 163.367
R645 B.n235 B.n234 163.367
R646 B.n234 B.n167 163.367
R647 B.n230 B.n167 163.367
R648 B.n230 B.n229 163.367
R649 B.n229 B.n228 163.367
R650 B.n228 B.n169 163.367
R651 B.n224 B.n169 163.367
R652 B.n224 B.n223 163.367
R653 B.n223 B.n222 163.367
R654 B.n222 B.n171 163.367
R655 B.n218 B.n171 163.367
R656 B.n218 B.n217 163.367
R657 B.n217 B.n216 163.367
R658 B.n216 B.n173 163.367
R659 B.n212 B.n173 163.367
R660 B.n212 B.n211 163.367
R661 B.n211 B.n210 163.367
R662 B.n210 B.n175 163.367
R663 B.n206 B.n175 163.367
R664 B.n206 B.n205 163.367
R665 B.n205 B.n204 163.367
R666 B.n204 B.n177 163.367
R667 B.n200 B.n177 163.367
R668 B.n200 B.n199 163.367
R669 B.n199 B.n198 163.367
R670 B.n198 B.n179 163.367
R671 B.n194 B.n179 163.367
R672 B.n194 B.n193 163.367
R673 B.n193 B.n192 163.367
R674 B.n192 B.n181 163.367
R675 B.n188 B.n181 163.367
R676 B.n188 B.n187 163.367
R677 B.n187 B.n186 163.367
R678 B.n186 B.n183 163.367
R679 B.n183 B.n2 163.367
R680 B.n706 B.n2 163.367
R681 B.n706 B.n705 163.367
R682 B.n705 B.n704 163.367
R683 B.n704 B.n3 163.367
R684 B.n700 B.n3 163.367
R685 B.n700 B.n699 163.367
R686 B.n699 B.n698 163.367
R687 B.n698 B.n5 163.367
R688 B.n694 B.n5 163.367
R689 B.n694 B.n693 163.367
R690 B.n693 B.n692 163.367
R691 B.n692 B.n7 163.367
R692 B.n688 B.n7 163.367
R693 B.n688 B.n687 163.367
R694 B.n687 B.n686 163.367
R695 B.n686 B.n9 163.367
R696 B.n682 B.n9 163.367
R697 B.n682 B.n681 163.367
R698 B.n681 B.n680 163.367
R699 B.n680 B.n11 163.367
R700 B.n676 B.n11 163.367
R701 B.n676 B.n675 163.367
R702 B.n675 B.n674 163.367
R703 B.n674 B.n13 163.367
R704 B.n670 B.n13 163.367
R705 B.n670 B.n669 163.367
R706 B.n669 B.n668 163.367
R707 B.n668 B.n15 163.367
R708 B.n664 B.n15 163.367
R709 B.n664 B.n663 163.367
R710 B.n663 B.n662 163.367
R711 B.n662 B.n17 163.367
R712 B.n658 B.n17 163.367
R713 B.n658 B.n657 163.367
R714 B.n657 B.n656 163.367
R715 B.n656 B.n19 163.367
R716 B.n652 B.n19 163.367
R717 B.n652 B.n651 163.367
R718 B.n651 B.n650 163.367
R719 B.n650 B.n21 163.367
R720 B.n646 B.n21 163.367
R721 B.n646 B.n645 163.367
R722 B.n645 B.n644 163.367
R723 B.n644 B.n23 163.367
R724 B.n248 B.n247 163.367
R725 B.n248 B.n161 163.367
R726 B.n252 B.n161 163.367
R727 B.n253 B.n252 163.367
R728 B.n254 B.n253 163.367
R729 B.n254 B.n159 163.367
R730 B.n258 B.n159 163.367
R731 B.n259 B.n258 163.367
R732 B.n260 B.n259 163.367
R733 B.n260 B.n157 163.367
R734 B.n264 B.n157 163.367
R735 B.n265 B.n264 163.367
R736 B.n266 B.n265 163.367
R737 B.n266 B.n155 163.367
R738 B.n270 B.n155 163.367
R739 B.n271 B.n270 163.367
R740 B.n272 B.n271 163.367
R741 B.n272 B.n153 163.367
R742 B.n276 B.n153 163.367
R743 B.n277 B.n276 163.367
R744 B.n278 B.n277 163.367
R745 B.n278 B.n151 163.367
R746 B.n282 B.n151 163.367
R747 B.n283 B.n282 163.367
R748 B.n284 B.n283 163.367
R749 B.n284 B.n149 163.367
R750 B.n288 B.n149 163.367
R751 B.n289 B.n288 163.367
R752 B.n290 B.n289 163.367
R753 B.n290 B.n147 163.367
R754 B.n294 B.n147 163.367
R755 B.n295 B.n294 163.367
R756 B.n296 B.n295 163.367
R757 B.n296 B.n145 163.367
R758 B.n300 B.n145 163.367
R759 B.n301 B.n300 163.367
R760 B.n302 B.n301 163.367
R761 B.n302 B.n141 163.367
R762 B.n307 B.n141 163.367
R763 B.n308 B.n307 163.367
R764 B.n309 B.n308 163.367
R765 B.n309 B.n139 163.367
R766 B.n313 B.n139 163.367
R767 B.n314 B.n313 163.367
R768 B.n315 B.n314 163.367
R769 B.n315 B.n137 163.367
R770 B.n319 B.n137 163.367
R771 B.n320 B.n319 163.367
R772 B.n320 B.n133 163.367
R773 B.n324 B.n133 163.367
R774 B.n325 B.n324 163.367
R775 B.n326 B.n325 163.367
R776 B.n326 B.n131 163.367
R777 B.n330 B.n131 163.367
R778 B.n331 B.n330 163.367
R779 B.n332 B.n331 163.367
R780 B.n332 B.n129 163.367
R781 B.n336 B.n129 163.367
R782 B.n337 B.n336 163.367
R783 B.n338 B.n337 163.367
R784 B.n338 B.n127 163.367
R785 B.n342 B.n127 163.367
R786 B.n343 B.n342 163.367
R787 B.n344 B.n343 163.367
R788 B.n344 B.n125 163.367
R789 B.n348 B.n125 163.367
R790 B.n349 B.n348 163.367
R791 B.n350 B.n349 163.367
R792 B.n350 B.n123 163.367
R793 B.n354 B.n123 163.367
R794 B.n355 B.n354 163.367
R795 B.n356 B.n355 163.367
R796 B.n356 B.n121 163.367
R797 B.n360 B.n121 163.367
R798 B.n361 B.n360 163.367
R799 B.n362 B.n361 163.367
R800 B.n362 B.n119 163.367
R801 B.n366 B.n119 163.367
R802 B.n367 B.n366 163.367
R803 B.n368 B.n367 163.367
R804 B.n368 B.n117 163.367
R805 B.n372 B.n117 163.367
R806 B.n373 B.n372 163.367
R807 B.n374 B.n373 163.367
R808 B.n374 B.n115 163.367
R809 B.n378 B.n115 163.367
R810 B.n380 B.n379 163.367
R811 B.n380 B.n113 163.367
R812 B.n384 B.n113 163.367
R813 B.n385 B.n384 163.367
R814 B.n386 B.n385 163.367
R815 B.n386 B.n111 163.367
R816 B.n390 B.n111 163.367
R817 B.n391 B.n390 163.367
R818 B.n392 B.n391 163.367
R819 B.n392 B.n109 163.367
R820 B.n396 B.n109 163.367
R821 B.n397 B.n396 163.367
R822 B.n398 B.n397 163.367
R823 B.n398 B.n107 163.367
R824 B.n402 B.n107 163.367
R825 B.n403 B.n402 163.367
R826 B.n404 B.n403 163.367
R827 B.n404 B.n105 163.367
R828 B.n408 B.n105 163.367
R829 B.n409 B.n408 163.367
R830 B.n410 B.n409 163.367
R831 B.n410 B.n103 163.367
R832 B.n414 B.n103 163.367
R833 B.n415 B.n414 163.367
R834 B.n416 B.n415 163.367
R835 B.n416 B.n101 163.367
R836 B.n420 B.n101 163.367
R837 B.n421 B.n420 163.367
R838 B.n422 B.n421 163.367
R839 B.n422 B.n99 163.367
R840 B.n426 B.n99 163.367
R841 B.n427 B.n426 163.367
R842 B.n428 B.n427 163.367
R843 B.n428 B.n97 163.367
R844 B.n432 B.n97 163.367
R845 B.n433 B.n432 163.367
R846 B.n434 B.n433 163.367
R847 B.n434 B.n95 163.367
R848 B.n438 B.n95 163.367
R849 B.n439 B.n438 163.367
R850 B.n440 B.n439 163.367
R851 B.n440 B.n93 163.367
R852 B.n444 B.n93 163.367
R853 B.n445 B.n444 163.367
R854 B.n446 B.n445 163.367
R855 B.n446 B.n91 163.367
R856 B.n450 B.n91 163.367
R857 B.n451 B.n450 163.367
R858 B.n452 B.n451 163.367
R859 B.n452 B.n89 163.367
R860 B.n456 B.n89 163.367
R861 B.n457 B.n456 163.367
R862 B.n458 B.n457 163.367
R863 B.n458 B.n87 163.367
R864 B.n462 B.n87 163.367
R865 B.n463 B.n462 163.367
R866 B.n464 B.n463 163.367
R867 B.n464 B.n85 163.367
R868 B.n468 B.n85 163.367
R869 B.n469 B.n468 163.367
R870 B.n470 B.n469 163.367
R871 B.n470 B.n83 163.367
R872 B.n474 B.n83 163.367
R873 B.n475 B.n474 163.367
R874 B.n476 B.n475 163.367
R875 B.n476 B.n81 163.367
R876 B.n480 B.n81 163.367
R877 B.n481 B.n480 163.367
R878 B.n482 B.n481 163.367
R879 B.n482 B.n79 163.367
R880 B.n486 B.n79 163.367
R881 B.n487 B.n486 163.367
R882 B.n488 B.n487 163.367
R883 B.n488 B.n77 163.367
R884 B.n492 B.n77 163.367
R885 B.n493 B.n492 163.367
R886 B.n494 B.n493 163.367
R887 B.n494 B.n75 163.367
R888 B.n498 B.n75 163.367
R889 B.n499 B.n498 163.367
R890 B.n500 B.n499 163.367
R891 B.n500 B.n73 163.367
R892 B.n504 B.n73 163.367
R893 B.n505 B.n504 163.367
R894 B.n506 B.n505 163.367
R895 B.n506 B.n71 163.367
R896 B.n640 B.n639 163.367
R897 B.n639 B.n638 163.367
R898 B.n638 B.n25 163.367
R899 B.n634 B.n25 163.367
R900 B.n634 B.n633 163.367
R901 B.n633 B.n632 163.367
R902 B.n632 B.n27 163.367
R903 B.n628 B.n27 163.367
R904 B.n628 B.n627 163.367
R905 B.n627 B.n626 163.367
R906 B.n626 B.n29 163.367
R907 B.n622 B.n29 163.367
R908 B.n622 B.n621 163.367
R909 B.n621 B.n620 163.367
R910 B.n620 B.n31 163.367
R911 B.n616 B.n31 163.367
R912 B.n616 B.n615 163.367
R913 B.n615 B.n614 163.367
R914 B.n614 B.n33 163.367
R915 B.n610 B.n33 163.367
R916 B.n610 B.n609 163.367
R917 B.n609 B.n608 163.367
R918 B.n608 B.n35 163.367
R919 B.n604 B.n35 163.367
R920 B.n604 B.n603 163.367
R921 B.n603 B.n602 163.367
R922 B.n602 B.n37 163.367
R923 B.n598 B.n37 163.367
R924 B.n598 B.n597 163.367
R925 B.n597 B.n596 163.367
R926 B.n596 B.n39 163.367
R927 B.n592 B.n39 163.367
R928 B.n592 B.n591 163.367
R929 B.n591 B.n590 163.367
R930 B.n590 B.n41 163.367
R931 B.n586 B.n41 163.367
R932 B.n586 B.n585 163.367
R933 B.n585 B.n584 163.367
R934 B.n584 B.n43 163.367
R935 B.n579 B.n43 163.367
R936 B.n579 B.n578 163.367
R937 B.n578 B.n577 163.367
R938 B.n577 B.n47 163.367
R939 B.n573 B.n47 163.367
R940 B.n573 B.n572 163.367
R941 B.n572 B.n571 163.367
R942 B.n571 B.n49 163.367
R943 B.n566 B.n49 163.367
R944 B.n566 B.n565 163.367
R945 B.n565 B.n564 163.367
R946 B.n564 B.n53 163.367
R947 B.n560 B.n53 163.367
R948 B.n560 B.n559 163.367
R949 B.n559 B.n558 163.367
R950 B.n558 B.n55 163.367
R951 B.n554 B.n55 163.367
R952 B.n554 B.n553 163.367
R953 B.n553 B.n552 163.367
R954 B.n552 B.n57 163.367
R955 B.n548 B.n57 163.367
R956 B.n548 B.n547 163.367
R957 B.n547 B.n546 163.367
R958 B.n546 B.n59 163.367
R959 B.n542 B.n59 163.367
R960 B.n542 B.n541 163.367
R961 B.n541 B.n540 163.367
R962 B.n540 B.n61 163.367
R963 B.n536 B.n61 163.367
R964 B.n536 B.n535 163.367
R965 B.n535 B.n534 163.367
R966 B.n534 B.n63 163.367
R967 B.n530 B.n63 163.367
R968 B.n530 B.n529 163.367
R969 B.n529 B.n528 163.367
R970 B.n528 B.n65 163.367
R971 B.n524 B.n65 163.367
R972 B.n524 B.n523 163.367
R973 B.n523 B.n522 163.367
R974 B.n522 B.n67 163.367
R975 B.n518 B.n67 163.367
R976 B.n518 B.n517 163.367
R977 B.n517 B.n516 163.367
R978 B.n516 B.n69 163.367
R979 B.n512 B.n69 163.367
R980 B.n512 B.n511 163.367
R981 B.n511 B.n510 163.367
R982 B.n134 B.t11 148.274
R983 B.n50 B.t4 148.274
R984 B.n142 B.t2 148.262
R985 B.n44 B.t7 148.262
R986 B.n135 B.t10 110.069
R987 B.n51 B.t5 110.069
R988 B.n143 B.t1 110.055
R989 B.n45 B.t8 110.055
R990 B.n136 B.n135 59.5399
R991 B.n305 B.n143 59.5399
R992 B.n582 B.n45 59.5399
R993 B.n568 B.n51 59.5399
R994 B.n135 B.n134 38.2066
R995 B.n143 B.n142 38.2066
R996 B.n45 B.n44 38.2066
R997 B.n51 B.n50 38.2066
R998 B.n642 B.n641 31.3761
R999 B.n509 B.n508 31.3761
R1000 B.n377 B.n114 31.3761
R1001 B.n245 B.n162 31.3761
R1002 B B.n707 18.0485
R1003 B.n641 B.n24 10.6151
R1004 B.n637 B.n24 10.6151
R1005 B.n637 B.n636 10.6151
R1006 B.n636 B.n635 10.6151
R1007 B.n635 B.n26 10.6151
R1008 B.n631 B.n26 10.6151
R1009 B.n631 B.n630 10.6151
R1010 B.n630 B.n629 10.6151
R1011 B.n629 B.n28 10.6151
R1012 B.n625 B.n28 10.6151
R1013 B.n625 B.n624 10.6151
R1014 B.n624 B.n623 10.6151
R1015 B.n623 B.n30 10.6151
R1016 B.n619 B.n30 10.6151
R1017 B.n619 B.n618 10.6151
R1018 B.n618 B.n617 10.6151
R1019 B.n617 B.n32 10.6151
R1020 B.n613 B.n32 10.6151
R1021 B.n613 B.n612 10.6151
R1022 B.n612 B.n611 10.6151
R1023 B.n611 B.n34 10.6151
R1024 B.n607 B.n34 10.6151
R1025 B.n607 B.n606 10.6151
R1026 B.n606 B.n605 10.6151
R1027 B.n605 B.n36 10.6151
R1028 B.n601 B.n36 10.6151
R1029 B.n601 B.n600 10.6151
R1030 B.n600 B.n599 10.6151
R1031 B.n599 B.n38 10.6151
R1032 B.n595 B.n38 10.6151
R1033 B.n595 B.n594 10.6151
R1034 B.n594 B.n593 10.6151
R1035 B.n593 B.n40 10.6151
R1036 B.n589 B.n40 10.6151
R1037 B.n589 B.n588 10.6151
R1038 B.n588 B.n587 10.6151
R1039 B.n587 B.n42 10.6151
R1040 B.n583 B.n42 10.6151
R1041 B.n581 B.n580 10.6151
R1042 B.n580 B.n46 10.6151
R1043 B.n576 B.n46 10.6151
R1044 B.n576 B.n575 10.6151
R1045 B.n575 B.n574 10.6151
R1046 B.n574 B.n48 10.6151
R1047 B.n570 B.n48 10.6151
R1048 B.n570 B.n569 10.6151
R1049 B.n567 B.n52 10.6151
R1050 B.n563 B.n52 10.6151
R1051 B.n563 B.n562 10.6151
R1052 B.n562 B.n561 10.6151
R1053 B.n561 B.n54 10.6151
R1054 B.n557 B.n54 10.6151
R1055 B.n557 B.n556 10.6151
R1056 B.n556 B.n555 10.6151
R1057 B.n555 B.n56 10.6151
R1058 B.n551 B.n56 10.6151
R1059 B.n551 B.n550 10.6151
R1060 B.n550 B.n549 10.6151
R1061 B.n549 B.n58 10.6151
R1062 B.n545 B.n58 10.6151
R1063 B.n545 B.n544 10.6151
R1064 B.n544 B.n543 10.6151
R1065 B.n543 B.n60 10.6151
R1066 B.n539 B.n60 10.6151
R1067 B.n539 B.n538 10.6151
R1068 B.n538 B.n537 10.6151
R1069 B.n537 B.n62 10.6151
R1070 B.n533 B.n62 10.6151
R1071 B.n533 B.n532 10.6151
R1072 B.n532 B.n531 10.6151
R1073 B.n531 B.n64 10.6151
R1074 B.n527 B.n64 10.6151
R1075 B.n527 B.n526 10.6151
R1076 B.n526 B.n525 10.6151
R1077 B.n525 B.n66 10.6151
R1078 B.n521 B.n66 10.6151
R1079 B.n521 B.n520 10.6151
R1080 B.n520 B.n519 10.6151
R1081 B.n519 B.n68 10.6151
R1082 B.n515 B.n68 10.6151
R1083 B.n515 B.n514 10.6151
R1084 B.n514 B.n513 10.6151
R1085 B.n513 B.n70 10.6151
R1086 B.n509 B.n70 10.6151
R1087 B.n381 B.n114 10.6151
R1088 B.n382 B.n381 10.6151
R1089 B.n383 B.n382 10.6151
R1090 B.n383 B.n112 10.6151
R1091 B.n387 B.n112 10.6151
R1092 B.n388 B.n387 10.6151
R1093 B.n389 B.n388 10.6151
R1094 B.n389 B.n110 10.6151
R1095 B.n393 B.n110 10.6151
R1096 B.n394 B.n393 10.6151
R1097 B.n395 B.n394 10.6151
R1098 B.n395 B.n108 10.6151
R1099 B.n399 B.n108 10.6151
R1100 B.n400 B.n399 10.6151
R1101 B.n401 B.n400 10.6151
R1102 B.n401 B.n106 10.6151
R1103 B.n405 B.n106 10.6151
R1104 B.n406 B.n405 10.6151
R1105 B.n407 B.n406 10.6151
R1106 B.n407 B.n104 10.6151
R1107 B.n411 B.n104 10.6151
R1108 B.n412 B.n411 10.6151
R1109 B.n413 B.n412 10.6151
R1110 B.n413 B.n102 10.6151
R1111 B.n417 B.n102 10.6151
R1112 B.n418 B.n417 10.6151
R1113 B.n419 B.n418 10.6151
R1114 B.n419 B.n100 10.6151
R1115 B.n423 B.n100 10.6151
R1116 B.n424 B.n423 10.6151
R1117 B.n425 B.n424 10.6151
R1118 B.n425 B.n98 10.6151
R1119 B.n429 B.n98 10.6151
R1120 B.n430 B.n429 10.6151
R1121 B.n431 B.n430 10.6151
R1122 B.n431 B.n96 10.6151
R1123 B.n435 B.n96 10.6151
R1124 B.n436 B.n435 10.6151
R1125 B.n437 B.n436 10.6151
R1126 B.n437 B.n94 10.6151
R1127 B.n441 B.n94 10.6151
R1128 B.n442 B.n441 10.6151
R1129 B.n443 B.n442 10.6151
R1130 B.n443 B.n92 10.6151
R1131 B.n447 B.n92 10.6151
R1132 B.n448 B.n447 10.6151
R1133 B.n449 B.n448 10.6151
R1134 B.n449 B.n90 10.6151
R1135 B.n453 B.n90 10.6151
R1136 B.n454 B.n453 10.6151
R1137 B.n455 B.n454 10.6151
R1138 B.n455 B.n88 10.6151
R1139 B.n459 B.n88 10.6151
R1140 B.n460 B.n459 10.6151
R1141 B.n461 B.n460 10.6151
R1142 B.n461 B.n86 10.6151
R1143 B.n465 B.n86 10.6151
R1144 B.n466 B.n465 10.6151
R1145 B.n467 B.n466 10.6151
R1146 B.n467 B.n84 10.6151
R1147 B.n471 B.n84 10.6151
R1148 B.n472 B.n471 10.6151
R1149 B.n473 B.n472 10.6151
R1150 B.n473 B.n82 10.6151
R1151 B.n477 B.n82 10.6151
R1152 B.n478 B.n477 10.6151
R1153 B.n479 B.n478 10.6151
R1154 B.n479 B.n80 10.6151
R1155 B.n483 B.n80 10.6151
R1156 B.n484 B.n483 10.6151
R1157 B.n485 B.n484 10.6151
R1158 B.n485 B.n78 10.6151
R1159 B.n489 B.n78 10.6151
R1160 B.n490 B.n489 10.6151
R1161 B.n491 B.n490 10.6151
R1162 B.n491 B.n76 10.6151
R1163 B.n495 B.n76 10.6151
R1164 B.n496 B.n495 10.6151
R1165 B.n497 B.n496 10.6151
R1166 B.n497 B.n74 10.6151
R1167 B.n501 B.n74 10.6151
R1168 B.n502 B.n501 10.6151
R1169 B.n503 B.n502 10.6151
R1170 B.n503 B.n72 10.6151
R1171 B.n507 B.n72 10.6151
R1172 B.n508 B.n507 10.6151
R1173 B.n249 B.n162 10.6151
R1174 B.n250 B.n249 10.6151
R1175 B.n251 B.n250 10.6151
R1176 B.n251 B.n160 10.6151
R1177 B.n255 B.n160 10.6151
R1178 B.n256 B.n255 10.6151
R1179 B.n257 B.n256 10.6151
R1180 B.n257 B.n158 10.6151
R1181 B.n261 B.n158 10.6151
R1182 B.n262 B.n261 10.6151
R1183 B.n263 B.n262 10.6151
R1184 B.n263 B.n156 10.6151
R1185 B.n267 B.n156 10.6151
R1186 B.n268 B.n267 10.6151
R1187 B.n269 B.n268 10.6151
R1188 B.n269 B.n154 10.6151
R1189 B.n273 B.n154 10.6151
R1190 B.n274 B.n273 10.6151
R1191 B.n275 B.n274 10.6151
R1192 B.n275 B.n152 10.6151
R1193 B.n279 B.n152 10.6151
R1194 B.n280 B.n279 10.6151
R1195 B.n281 B.n280 10.6151
R1196 B.n281 B.n150 10.6151
R1197 B.n285 B.n150 10.6151
R1198 B.n286 B.n285 10.6151
R1199 B.n287 B.n286 10.6151
R1200 B.n287 B.n148 10.6151
R1201 B.n291 B.n148 10.6151
R1202 B.n292 B.n291 10.6151
R1203 B.n293 B.n292 10.6151
R1204 B.n293 B.n146 10.6151
R1205 B.n297 B.n146 10.6151
R1206 B.n298 B.n297 10.6151
R1207 B.n299 B.n298 10.6151
R1208 B.n299 B.n144 10.6151
R1209 B.n303 B.n144 10.6151
R1210 B.n304 B.n303 10.6151
R1211 B.n306 B.n140 10.6151
R1212 B.n310 B.n140 10.6151
R1213 B.n311 B.n310 10.6151
R1214 B.n312 B.n311 10.6151
R1215 B.n312 B.n138 10.6151
R1216 B.n316 B.n138 10.6151
R1217 B.n317 B.n316 10.6151
R1218 B.n318 B.n317 10.6151
R1219 B.n322 B.n321 10.6151
R1220 B.n323 B.n322 10.6151
R1221 B.n323 B.n132 10.6151
R1222 B.n327 B.n132 10.6151
R1223 B.n328 B.n327 10.6151
R1224 B.n329 B.n328 10.6151
R1225 B.n329 B.n130 10.6151
R1226 B.n333 B.n130 10.6151
R1227 B.n334 B.n333 10.6151
R1228 B.n335 B.n334 10.6151
R1229 B.n335 B.n128 10.6151
R1230 B.n339 B.n128 10.6151
R1231 B.n340 B.n339 10.6151
R1232 B.n341 B.n340 10.6151
R1233 B.n341 B.n126 10.6151
R1234 B.n345 B.n126 10.6151
R1235 B.n346 B.n345 10.6151
R1236 B.n347 B.n346 10.6151
R1237 B.n347 B.n124 10.6151
R1238 B.n351 B.n124 10.6151
R1239 B.n352 B.n351 10.6151
R1240 B.n353 B.n352 10.6151
R1241 B.n353 B.n122 10.6151
R1242 B.n357 B.n122 10.6151
R1243 B.n358 B.n357 10.6151
R1244 B.n359 B.n358 10.6151
R1245 B.n359 B.n120 10.6151
R1246 B.n363 B.n120 10.6151
R1247 B.n364 B.n363 10.6151
R1248 B.n365 B.n364 10.6151
R1249 B.n365 B.n118 10.6151
R1250 B.n369 B.n118 10.6151
R1251 B.n370 B.n369 10.6151
R1252 B.n371 B.n370 10.6151
R1253 B.n371 B.n116 10.6151
R1254 B.n375 B.n116 10.6151
R1255 B.n376 B.n375 10.6151
R1256 B.n377 B.n376 10.6151
R1257 B.n245 B.n244 10.6151
R1258 B.n244 B.n243 10.6151
R1259 B.n243 B.n164 10.6151
R1260 B.n239 B.n164 10.6151
R1261 B.n239 B.n238 10.6151
R1262 B.n238 B.n237 10.6151
R1263 B.n237 B.n166 10.6151
R1264 B.n233 B.n166 10.6151
R1265 B.n233 B.n232 10.6151
R1266 B.n232 B.n231 10.6151
R1267 B.n231 B.n168 10.6151
R1268 B.n227 B.n168 10.6151
R1269 B.n227 B.n226 10.6151
R1270 B.n226 B.n225 10.6151
R1271 B.n225 B.n170 10.6151
R1272 B.n221 B.n170 10.6151
R1273 B.n221 B.n220 10.6151
R1274 B.n220 B.n219 10.6151
R1275 B.n219 B.n172 10.6151
R1276 B.n215 B.n172 10.6151
R1277 B.n215 B.n214 10.6151
R1278 B.n214 B.n213 10.6151
R1279 B.n213 B.n174 10.6151
R1280 B.n209 B.n174 10.6151
R1281 B.n209 B.n208 10.6151
R1282 B.n208 B.n207 10.6151
R1283 B.n207 B.n176 10.6151
R1284 B.n203 B.n176 10.6151
R1285 B.n203 B.n202 10.6151
R1286 B.n202 B.n201 10.6151
R1287 B.n201 B.n178 10.6151
R1288 B.n197 B.n178 10.6151
R1289 B.n197 B.n196 10.6151
R1290 B.n196 B.n195 10.6151
R1291 B.n195 B.n180 10.6151
R1292 B.n191 B.n180 10.6151
R1293 B.n191 B.n190 10.6151
R1294 B.n190 B.n189 10.6151
R1295 B.n189 B.n182 10.6151
R1296 B.n185 B.n182 10.6151
R1297 B.n185 B.n184 10.6151
R1298 B.n184 B.n0 10.6151
R1299 B.n703 B.n1 10.6151
R1300 B.n703 B.n702 10.6151
R1301 B.n702 B.n701 10.6151
R1302 B.n701 B.n4 10.6151
R1303 B.n697 B.n4 10.6151
R1304 B.n697 B.n696 10.6151
R1305 B.n696 B.n695 10.6151
R1306 B.n695 B.n6 10.6151
R1307 B.n691 B.n6 10.6151
R1308 B.n691 B.n690 10.6151
R1309 B.n690 B.n689 10.6151
R1310 B.n689 B.n8 10.6151
R1311 B.n685 B.n8 10.6151
R1312 B.n685 B.n684 10.6151
R1313 B.n684 B.n683 10.6151
R1314 B.n683 B.n10 10.6151
R1315 B.n679 B.n10 10.6151
R1316 B.n679 B.n678 10.6151
R1317 B.n678 B.n677 10.6151
R1318 B.n677 B.n12 10.6151
R1319 B.n673 B.n12 10.6151
R1320 B.n673 B.n672 10.6151
R1321 B.n672 B.n671 10.6151
R1322 B.n671 B.n14 10.6151
R1323 B.n667 B.n14 10.6151
R1324 B.n667 B.n666 10.6151
R1325 B.n666 B.n665 10.6151
R1326 B.n665 B.n16 10.6151
R1327 B.n661 B.n16 10.6151
R1328 B.n661 B.n660 10.6151
R1329 B.n660 B.n659 10.6151
R1330 B.n659 B.n18 10.6151
R1331 B.n655 B.n18 10.6151
R1332 B.n655 B.n654 10.6151
R1333 B.n654 B.n653 10.6151
R1334 B.n653 B.n20 10.6151
R1335 B.n649 B.n20 10.6151
R1336 B.n649 B.n648 10.6151
R1337 B.n648 B.n647 10.6151
R1338 B.n647 B.n22 10.6151
R1339 B.n643 B.n22 10.6151
R1340 B.n643 B.n642 10.6151
R1341 B.n582 B.n581 6.5566
R1342 B.n569 B.n568 6.5566
R1343 B.n306 B.n305 6.5566
R1344 B.n318 B.n136 6.5566
R1345 B.n583 B.n582 4.05904
R1346 B.n568 B.n567 4.05904
R1347 B.n305 B.n304 4.05904
R1348 B.n321 B.n136 4.05904
R1349 B.n707 B.n0 2.81026
R1350 B.n707 B.n1 2.81026
C0 VN B 1.03054f
C1 B VDD2 2.10378f
C2 VN VP 6.79455f
C3 VN VDD1 0.15164f
C4 VDD2 VP 0.461571f
C5 VDD1 VDD2 1.55096f
C6 VTAIL B 3.08639f
C7 B w_n3334_n3172# 8.65751f
C8 VTAIL VP 9.069969f
C9 VTAIL VDD1 10.153099f
C10 w_n3334_n3172# VP 7.23269f
C11 VN VDD2 8.77509f
C12 VDD1 w_n3334_n3172# 2.3552f
C13 VTAIL VN 9.055599f
C14 B VP 1.75018f
C15 VN w_n3334_n3172# 6.80158f
C16 VTAIL VDD2 10.1966f
C17 VDD1 B 2.02325f
C18 w_n3334_n3172# VDD2 2.44896f
C19 VDD1 VP 9.081231f
C20 VTAIL w_n3334_n3172# 2.95612f
C21 VDD2 VSUBS 1.76113f
C22 VDD1 VSUBS 1.53316f
C23 VTAIL VSUBS 1.028453f
C24 VN VSUBS 6.10356f
C25 VP VSUBS 2.969588f
C26 B VSUBS 4.093238f
C27 w_n3334_n3172# VSUBS 0.130386p
C28 B.n0 VSUBS 0.005796f
C29 B.n1 VSUBS 0.005796f
C30 B.n2 VSUBS 0.009165f
C31 B.n3 VSUBS 0.009165f
C32 B.n4 VSUBS 0.009165f
C33 B.n5 VSUBS 0.009165f
C34 B.n6 VSUBS 0.009165f
C35 B.n7 VSUBS 0.009165f
C36 B.n8 VSUBS 0.009165f
C37 B.n9 VSUBS 0.009165f
C38 B.n10 VSUBS 0.009165f
C39 B.n11 VSUBS 0.009165f
C40 B.n12 VSUBS 0.009165f
C41 B.n13 VSUBS 0.009165f
C42 B.n14 VSUBS 0.009165f
C43 B.n15 VSUBS 0.009165f
C44 B.n16 VSUBS 0.009165f
C45 B.n17 VSUBS 0.009165f
C46 B.n18 VSUBS 0.009165f
C47 B.n19 VSUBS 0.009165f
C48 B.n20 VSUBS 0.009165f
C49 B.n21 VSUBS 0.009165f
C50 B.n22 VSUBS 0.009165f
C51 B.n23 VSUBS 0.020493f
C52 B.n24 VSUBS 0.009165f
C53 B.n25 VSUBS 0.009165f
C54 B.n26 VSUBS 0.009165f
C55 B.n27 VSUBS 0.009165f
C56 B.n28 VSUBS 0.009165f
C57 B.n29 VSUBS 0.009165f
C58 B.n30 VSUBS 0.009165f
C59 B.n31 VSUBS 0.009165f
C60 B.n32 VSUBS 0.009165f
C61 B.n33 VSUBS 0.009165f
C62 B.n34 VSUBS 0.009165f
C63 B.n35 VSUBS 0.009165f
C64 B.n36 VSUBS 0.009165f
C65 B.n37 VSUBS 0.009165f
C66 B.n38 VSUBS 0.009165f
C67 B.n39 VSUBS 0.009165f
C68 B.n40 VSUBS 0.009165f
C69 B.n41 VSUBS 0.009165f
C70 B.n42 VSUBS 0.009165f
C71 B.n43 VSUBS 0.009165f
C72 B.t8 VSUBS 0.465739f
C73 B.t7 VSUBS 0.485227f
C74 B.t6 VSUBS 1.04832f
C75 B.n44 VSUBS 0.224593f
C76 B.n45 VSUBS 0.088694f
C77 B.n46 VSUBS 0.009165f
C78 B.n47 VSUBS 0.009165f
C79 B.n48 VSUBS 0.009165f
C80 B.n49 VSUBS 0.009165f
C81 B.t5 VSUBS 0.465732f
C82 B.t4 VSUBS 0.485219f
C83 B.t3 VSUBS 1.04832f
C84 B.n50 VSUBS 0.2246f
C85 B.n51 VSUBS 0.088702f
C86 B.n52 VSUBS 0.009165f
C87 B.n53 VSUBS 0.009165f
C88 B.n54 VSUBS 0.009165f
C89 B.n55 VSUBS 0.009165f
C90 B.n56 VSUBS 0.009165f
C91 B.n57 VSUBS 0.009165f
C92 B.n58 VSUBS 0.009165f
C93 B.n59 VSUBS 0.009165f
C94 B.n60 VSUBS 0.009165f
C95 B.n61 VSUBS 0.009165f
C96 B.n62 VSUBS 0.009165f
C97 B.n63 VSUBS 0.009165f
C98 B.n64 VSUBS 0.009165f
C99 B.n65 VSUBS 0.009165f
C100 B.n66 VSUBS 0.009165f
C101 B.n67 VSUBS 0.009165f
C102 B.n68 VSUBS 0.009165f
C103 B.n69 VSUBS 0.009165f
C104 B.n70 VSUBS 0.009165f
C105 B.n71 VSUBS 0.020493f
C106 B.n72 VSUBS 0.009165f
C107 B.n73 VSUBS 0.009165f
C108 B.n74 VSUBS 0.009165f
C109 B.n75 VSUBS 0.009165f
C110 B.n76 VSUBS 0.009165f
C111 B.n77 VSUBS 0.009165f
C112 B.n78 VSUBS 0.009165f
C113 B.n79 VSUBS 0.009165f
C114 B.n80 VSUBS 0.009165f
C115 B.n81 VSUBS 0.009165f
C116 B.n82 VSUBS 0.009165f
C117 B.n83 VSUBS 0.009165f
C118 B.n84 VSUBS 0.009165f
C119 B.n85 VSUBS 0.009165f
C120 B.n86 VSUBS 0.009165f
C121 B.n87 VSUBS 0.009165f
C122 B.n88 VSUBS 0.009165f
C123 B.n89 VSUBS 0.009165f
C124 B.n90 VSUBS 0.009165f
C125 B.n91 VSUBS 0.009165f
C126 B.n92 VSUBS 0.009165f
C127 B.n93 VSUBS 0.009165f
C128 B.n94 VSUBS 0.009165f
C129 B.n95 VSUBS 0.009165f
C130 B.n96 VSUBS 0.009165f
C131 B.n97 VSUBS 0.009165f
C132 B.n98 VSUBS 0.009165f
C133 B.n99 VSUBS 0.009165f
C134 B.n100 VSUBS 0.009165f
C135 B.n101 VSUBS 0.009165f
C136 B.n102 VSUBS 0.009165f
C137 B.n103 VSUBS 0.009165f
C138 B.n104 VSUBS 0.009165f
C139 B.n105 VSUBS 0.009165f
C140 B.n106 VSUBS 0.009165f
C141 B.n107 VSUBS 0.009165f
C142 B.n108 VSUBS 0.009165f
C143 B.n109 VSUBS 0.009165f
C144 B.n110 VSUBS 0.009165f
C145 B.n111 VSUBS 0.009165f
C146 B.n112 VSUBS 0.009165f
C147 B.n113 VSUBS 0.009165f
C148 B.n114 VSUBS 0.020493f
C149 B.n115 VSUBS 0.009165f
C150 B.n116 VSUBS 0.009165f
C151 B.n117 VSUBS 0.009165f
C152 B.n118 VSUBS 0.009165f
C153 B.n119 VSUBS 0.009165f
C154 B.n120 VSUBS 0.009165f
C155 B.n121 VSUBS 0.009165f
C156 B.n122 VSUBS 0.009165f
C157 B.n123 VSUBS 0.009165f
C158 B.n124 VSUBS 0.009165f
C159 B.n125 VSUBS 0.009165f
C160 B.n126 VSUBS 0.009165f
C161 B.n127 VSUBS 0.009165f
C162 B.n128 VSUBS 0.009165f
C163 B.n129 VSUBS 0.009165f
C164 B.n130 VSUBS 0.009165f
C165 B.n131 VSUBS 0.009165f
C166 B.n132 VSUBS 0.009165f
C167 B.n133 VSUBS 0.009165f
C168 B.t10 VSUBS 0.465732f
C169 B.t11 VSUBS 0.485219f
C170 B.t9 VSUBS 1.04832f
C171 B.n134 VSUBS 0.2246f
C172 B.n135 VSUBS 0.088702f
C173 B.n136 VSUBS 0.021235f
C174 B.n137 VSUBS 0.009165f
C175 B.n138 VSUBS 0.009165f
C176 B.n139 VSUBS 0.009165f
C177 B.n140 VSUBS 0.009165f
C178 B.n141 VSUBS 0.009165f
C179 B.t1 VSUBS 0.465739f
C180 B.t2 VSUBS 0.485227f
C181 B.t0 VSUBS 1.04832f
C182 B.n142 VSUBS 0.224593f
C183 B.n143 VSUBS 0.088694f
C184 B.n144 VSUBS 0.009165f
C185 B.n145 VSUBS 0.009165f
C186 B.n146 VSUBS 0.009165f
C187 B.n147 VSUBS 0.009165f
C188 B.n148 VSUBS 0.009165f
C189 B.n149 VSUBS 0.009165f
C190 B.n150 VSUBS 0.009165f
C191 B.n151 VSUBS 0.009165f
C192 B.n152 VSUBS 0.009165f
C193 B.n153 VSUBS 0.009165f
C194 B.n154 VSUBS 0.009165f
C195 B.n155 VSUBS 0.009165f
C196 B.n156 VSUBS 0.009165f
C197 B.n157 VSUBS 0.009165f
C198 B.n158 VSUBS 0.009165f
C199 B.n159 VSUBS 0.009165f
C200 B.n160 VSUBS 0.009165f
C201 B.n161 VSUBS 0.009165f
C202 B.n162 VSUBS 0.02129f
C203 B.n163 VSUBS 0.009165f
C204 B.n164 VSUBS 0.009165f
C205 B.n165 VSUBS 0.009165f
C206 B.n166 VSUBS 0.009165f
C207 B.n167 VSUBS 0.009165f
C208 B.n168 VSUBS 0.009165f
C209 B.n169 VSUBS 0.009165f
C210 B.n170 VSUBS 0.009165f
C211 B.n171 VSUBS 0.009165f
C212 B.n172 VSUBS 0.009165f
C213 B.n173 VSUBS 0.009165f
C214 B.n174 VSUBS 0.009165f
C215 B.n175 VSUBS 0.009165f
C216 B.n176 VSUBS 0.009165f
C217 B.n177 VSUBS 0.009165f
C218 B.n178 VSUBS 0.009165f
C219 B.n179 VSUBS 0.009165f
C220 B.n180 VSUBS 0.009165f
C221 B.n181 VSUBS 0.009165f
C222 B.n182 VSUBS 0.009165f
C223 B.n183 VSUBS 0.009165f
C224 B.n184 VSUBS 0.009165f
C225 B.n185 VSUBS 0.009165f
C226 B.n186 VSUBS 0.009165f
C227 B.n187 VSUBS 0.009165f
C228 B.n188 VSUBS 0.009165f
C229 B.n189 VSUBS 0.009165f
C230 B.n190 VSUBS 0.009165f
C231 B.n191 VSUBS 0.009165f
C232 B.n192 VSUBS 0.009165f
C233 B.n193 VSUBS 0.009165f
C234 B.n194 VSUBS 0.009165f
C235 B.n195 VSUBS 0.009165f
C236 B.n196 VSUBS 0.009165f
C237 B.n197 VSUBS 0.009165f
C238 B.n198 VSUBS 0.009165f
C239 B.n199 VSUBS 0.009165f
C240 B.n200 VSUBS 0.009165f
C241 B.n201 VSUBS 0.009165f
C242 B.n202 VSUBS 0.009165f
C243 B.n203 VSUBS 0.009165f
C244 B.n204 VSUBS 0.009165f
C245 B.n205 VSUBS 0.009165f
C246 B.n206 VSUBS 0.009165f
C247 B.n207 VSUBS 0.009165f
C248 B.n208 VSUBS 0.009165f
C249 B.n209 VSUBS 0.009165f
C250 B.n210 VSUBS 0.009165f
C251 B.n211 VSUBS 0.009165f
C252 B.n212 VSUBS 0.009165f
C253 B.n213 VSUBS 0.009165f
C254 B.n214 VSUBS 0.009165f
C255 B.n215 VSUBS 0.009165f
C256 B.n216 VSUBS 0.009165f
C257 B.n217 VSUBS 0.009165f
C258 B.n218 VSUBS 0.009165f
C259 B.n219 VSUBS 0.009165f
C260 B.n220 VSUBS 0.009165f
C261 B.n221 VSUBS 0.009165f
C262 B.n222 VSUBS 0.009165f
C263 B.n223 VSUBS 0.009165f
C264 B.n224 VSUBS 0.009165f
C265 B.n225 VSUBS 0.009165f
C266 B.n226 VSUBS 0.009165f
C267 B.n227 VSUBS 0.009165f
C268 B.n228 VSUBS 0.009165f
C269 B.n229 VSUBS 0.009165f
C270 B.n230 VSUBS 0.009165f
C271 B.n231 VSUBS 0.009165f
C272 B.n232 VSUBS 0.009165f
C273 B.n233 VSUBS 0.009165f
C274 B.n234 VSUBS 0.009165f
C275 B.n235 VSUBS 0.009165f
C276 B.n236 VSUBS 0.009165f
C277 B.n237 VSUBS 0.009165f
C278 B.n238 VSUBS 0.009165f
C279 B.n239 VSUBS 0.009165f
C280 B.n240 VSUBS 0.009165f
C281 B.n241 VSUBS 0.009165f
C282 B.n242 VSUBS 0.009165f
C283 B.n243 VSUBS 0.009165f
C284 B.n244 VSUBS 0.009165f
C285 B.n245 VSUBS 0.020493f
C286 B.n246 VSUBS 0.020493f
C287 B.n247 VSUBS 0.02129f
C288 B.n248 VSUBS 0.009165f
C289 B.n249 VSUBS 0.009165f
C290 B.n250 VSUBS 0.009165f
C291 B.n251 VSUBS 0.009165f
C292 B.n252 VSUBS 0.009165f
C293 B.n253 VSUBS 0.009165f
C294 B.n254 VSUBS 0.009165f
C295 B.n255 VSUBS 0.009165f
C296 B.n256 VSUBS 0.009165f
C297 B.n257 VSUBS 0.009165f
C298 B.n258 VSUBS 0.009165f
C299 B.n259 VSUBS 0.009165f
C300 B.n260 VSUBS 0.009165f
C301 B.n261 VSUBS 0.009165f
C302 B.n262 VSUBS 0.009165f
C303 B.n263 VSUBS 0.009165f
C304 B.n264 VSUBS 0.009165f
C305 B.n265 VSUBS 0.009165f
C306 B.n266 VSUBS 0.009165f
C307 B.n267 VSUBS 0.009165f
C308 B.n268 VSUBS 0.009165f
C309 B.n269 VSUBS 0.009165f
C310 B.n270 VSUBS 0.009165f
C311 B.n271 VSUBS 0.009165f
C312 B.n272 VSUBS 0.009165f
C313 B.n273 VSUBS 0.009165f
C314 B.n274 VSUBS 0.009165f
C315 B.n275 VSUBS 0.009165f
C316 B.n276 VSUBS 0.009165f
C317 B.n277 VSUBS 0.009165f
C318 B.n278 VSUBS 0.009165f
C319 B.n279 VSUBS 0.009165f
C320 B.n280 VSUBS 0.009165f
C321 B.n281 VSUBS 0.009165f
C322 B.n282 VSUBS 0.009165f
C323 B.n283 VSUBS 0.009165f
C324 B.n284 VSUBS 0.009165f
C325 B.n285 VSUBS 0.009165f
C326 B.n286 VSUBS 0.009165f
C327 B.n287 VSUBS 0.009165f
C328 B.n288 VSUBS 0.009165f
C329 B.n289 VSUBS 0.009165f
C330 B.n290 VSUBS 0.009165f
C331 B.n291 VSUBS 0.009165f
C332 B.n292 VSUBS 0.009165f
C333 B.n293 VSUBS 0.009165f
C334 B.n294 VSUBS 0.009165f
C335 B.n295 VSUBS 0.009165f
C336 B.n296 VSUBS 0.009165f
C337 B.n297 VSUBS 0.009165f
C338 B.n298 VSUBS 0.009165f
C339 B.n299 VSUBS 0.009165f
C340 B.n300 VSUBS 0.009165f
C341 B.n301 VSUBS 0.009165f
C342 B.n302 VSUBS 0.009165f
C343 B.n303 VSUBS 0.009165f
C344 B.n304 VSUBS 0.006335f
C345 B.n305 VSUBS 0.021235f
C346 B.n306 VSUBS 0.007413f
C347 B.n307 VSUBS 0.009165f
C348 B.n308 VSUBS 0.009165f
C349 B.n309 VSUBS 0.009165f
C350 B.n310 VSUBS 0.009165f
C351 B.n311 VSUBS 0.009165f
C352 B.n312 VSUBS 0.009165f
C353 B.n313 VSUBS 0.009165f
C354 B.n314 VSUBS 0.009165f
C355 B.n315 VSUBS 0.009165f
C356 B.n316 VSUBS 0.009165f
C357 B.n317 VSUBS 0.009165f
C358 B.n318 VSUBS 0.007413f
C359 B.n319 VSUBS 0.009165f
C360 B.n320 VSUBS 0.009165f
C361 B.n321 VSUBS 0.006335f
C362 B.n322 VSUBS 0.009165f
C363 B.n323 VSUBS 0.009165f
C364 B.n324 VSUBS 0.009165f
C365 B.n325 VSUBS 0.009165f
C366 B.n326 VSUBS 0.009165f
C367 B.n327 VSUBS 0.009165f
C368 B.n328 VSUBS 0.009165f
C369 B.n329 VSUBS 0.009165f
C370 B.n330 VSUBS 0.009165f
C371 B.n331 VSUBS 0.009165f
C372 B.n332 VSUBS 0.009165f
C373 B.n333 VSUBS 0.009165f
C374 B.n334 VSUBS 0.009165f
C375 B.n335 VSUBS 0.009165f
C376 B.n336 VSUBS 0.009165f
C377 B.n337 VSUBS 0.009165f
C378 B.n338 VSUBS 0.009165f
C379 B.n339 VSUBS 0.009165f
C380 B.n340 VSUBS 0.009165f
C381 B.n341 VSUBS 0.009165f
C382 B.n342 VSUBS 0.009165f
C383 B.n343 VSUBS 0.009165f
C384 B.n344 VSUBS 0.009165f
C385 B.n345 VSUBS 0.009165f
C386 B.n346 VSUBS 0.009165f
C387 B.n347 VSUBS 0.009165f
C388 B.n348 VSUBS 0.009165f
C389 B.n349 VSUBS 0.009165f
C390 B.n350 VSUBS 0.009165f
C391 B.n351 VSUBS 0.009165f
C392 B.n352 VSUBS 0.009165f
C393 B.n353 VSUBS 0.009165f
C394 B.n354 VSUBS 0.009165f
C395 B.n355 VSUBS 0.009165f
C396 B.n356 VSUBS 0.009165f
C397 B.n357 VSUBS 0.009165f
C398 B.n358 VSUBS 0.009165f
C399 B.n359 VSUBS 0.009165f
C400 B.n360 VSUBS 0.009165f
C401 B.n361 VSUBS 0.009165f
C402 B.n362 VSUBS 0.009165f
C403 B.n363 VSUBS 0.009165f
C404 B.n364 VSUBS 0.009165f
C405 B.n365 VSUBS 0.009165f
C406 B.n366 VSUBS 0.009165f
C407 B.n367 VSUBS 0.009165f
C408 B.n368 VSUBS 0.009165f
C409 B.n369 VSUBS 0.009165f
C410 B.n370 VSUBS 0.009165f
C411 B.n371 VSUBS 0.009165f
C412 B.n372 VSUBS 0.009165f
C413 B.n373 VSUBS 0.009165f
C414 B.n374 VSUBS 0.009165f
C415 B.n375 VSUBS 0.009165f
C416 B.n376 VSUBS 0.009165f
C417 B.n377 VSUBS 0.02129f
C418 B.n378 VSUBS 0.02129f
C419 B.n379 VSUBS 0.020493f
C420 B.n380 VSUBS 0.009165f
C421 B.n381 VSUBS 0.009165f
C422 B.n382 VSUBS 0.009165f
C423 B.n383 VSUBS 0.009165f
C424 B.n384 VSUBS 0.009165f
C425 B.n385 VSUBS 0.009165f
C426 B.n386 VSUBS 0.009165f
C427 B.n387 VSUBS 0.009165f
C428 B.n388 VSUBS 0.009165f
C429 B.n389 VSUBS 0.009165f
C430 B.n390 VSUBS 0.009165f
C431 B.n391 VSUBS 0.009165f
C432 B.n392 VSUBS 0.009165f
C433 B.n393 VSUBS 0.009165f
C434 B.n394 VSUBS 0.009165f
C435 B.n395 VSUBS 0.009165f
C436 B.n396 VSUBS 0.009165f
C437 B.n397 VSUBS 0.009165f
C438 B.n398 VSUBS 0.009165f
C439 B.n399 VSUBS 0.009165f
C440 B.n400 VSUBS 0.009165f
C441 B.n401 VSUBS 0.009165f
C442 B.n402 VSUBS 0.009165f
C443 B.n403 VSUBS 0.009165f
C444 B.n404 VSUBS 0.009165f
C445 B.n405 VSUBS 0.009165f
C446 B.n406 VSUBS 0.009165f
C447 B.n407 VSUBS 0.009165f
C448 B.n408 VSUBS 0.009165f
C449 B.n409 VSUBS 0.009165f
C450 B.n410 VSUBS 0.009165f
C451 B.n411 VSUBS 0.009165f
C452 B.n412 VSUBS 0.009165f
C453 B.n413 VSUBS 0.009165f
C454 B.n414 VSUBS 0.009165f
C455 B.n415 VSUBS 0.009165f
C456 B.n416 VSUBS 0.009165f
C457 B.n417 VSUBS 0.009165f
C458 B.n418 VSUBS 0.009165f
C459 B.n419 VSUBS 0.009165f
C460 B.n420 VSUBS 0.009165f
C461 B.n421 VSUBS 0.009165f
C462 B.n422 VSUBS 0.009165f
C463 B.n423 VSUBS 0.009165f
C464 B.n424 VSUBS 0.009165f
C465 B.n425 VSUBS 0.009165f
C466 B.n426 VSUBS 0.009165f
C467 B.n427 VSUBS 0.009165f
C468 B.n428 VSUBS 0.009165f
C469 B.n429 VSUBS 0.009165f
C470 B.n430 VSUBS 0.009165f
C471 B.n431 VSUBS 0.009165f
C472 B.n432 VSUBS 0.009165f
C473 B.n433 VSUBS 0.009165f
C474 B.n434 VSUBS 0.009165f
C475 B.n435 VSUBS 0.009165f
C476 B.n436 VSUBS 0.009165f
C477 B.n437 VSUBS 0.009165f
C478 B.n438 VSUBS 0.009165f
C479 B.n439 VSUBS 0.009165f
C480 B.n440 VSUBS 0.009165f
C481 B.n441 VSUBS 0.009165f
C482 B.n442 VSUBS 0.009165f
C483 B.n443 VSUBS 0.009165f
C484 B.n444 VSUBS 0.009165f
C485 B.n445 VSUBS 0.009165f
C486 B.n446 VSUBS 0.009165f
C487 B.n447 VSUBS 0.009165f
C488 B.n448 VSUBS 0.009165f
C489 B.n449 VSUBS 0.009165f
C490 B.n450 VSUBS 0.009165f
C491 B.n451 VSUBS 0.009165f
C492 B.n452 VSUBS 0.009165f
C493 B.n453 VSUBS 0.009165f
C494 B.n454 VSUBS 0.009165f
C495 B.n455 VSUBS 0.009165f
C496 B.n456 VSUBS 0.009165f
C497 B.n457 VSUBS 0.009165f
C498 B.n458 VSUBS 0.009165f
C499 B.n459 VSUBS 0.009165f
C500 B.n460 VSUBS 0.009165f
C501 B.n461 VSUBS 0.009165f
C502 B.n462 VSUBS 0.009165f
C503 B.n463 VSUBS 0.009165f
C504 B.n464 VSUBS 0.009165f
C505 B.n465 VSUBS 0.009165f
C506 B.n466 VSUBS 0.009165f
C507 B.n467 VSUBS 0.009165f
C508 B.n468 VSUBS 0.009165f
C509 B.n469 VSUBS 0.009165f
C510 B.n470 VSUBS 0.009165f
C511 B.n471 VSUBS 0.009165f
C512 B.n472 VSUBS 0.009165f
C513 B.n473 VSUBS 0.009165f
C514 B.n474 VSUBS 0.009165f
C515 B.n475 VSUBS 0.009165f
C516 B.n476 VSUBS 0.009165f
C517 B.n477 VSUBS 0.009165f
C518 B.n478 VSUBS 0.009165f
C519 B.n479 VSUBS 0.009165f
C520 B.n480 VSUBS 0.009165f
C521 B.n481 VSUBS 0.009165f
C522 B.n482 VSUBS 0.009165f
C523 B.n483 VSUBS 0.009165f
C524 B.n484 VSUBS 0.009165f
C525 B.n485 VSUBS 0.009165f
C526 B.n486 VSUBS 0.009165f
C527 B.n487 VSUBS 0.009165f
C528 B.n488 VSUBS 0.009165f
C529 B.n489 VSUBS 0.009165f
C530 B.n490 VSUBS 0.009165f
C531 B.n491 VSUBS 0.009165f
C532 B.n492 VSUBS 0.009165f
C533 B.n493 VSUBS 0.009165f
C534 B.n494 VSUBS 0.009165f
C535 B.n495 VSUBS 0.009165f
C536 B.n496 VSUBS 0.009165f
C537 B.n497 VSUBS 0.009165f
C538 B.n498 VSUBS 0.009165f
C539 B.n499 VSUBS 0.009165f
C540 B.n500 VSUBS 0.009165f
C541 B.n501 VSUBS 0.009165f
C542 B.n502 VSUBS 0.009165f
C543 B.n503 VSUBS 0.009165f
C544 B.n504 VSUBS 0.009165f
C545 B.n505 VSUBS 0.009165f
C546 B.n506 VSUBS 0.009165f
C547 B.n507 VSUBS 0.009165f
C548 B.n508 VSUBS 0.02162f
C549 B.n509 VSUBS 0.020163f
C550 B.n510 VSUBS 0.02129f
C551 B.n511 VSUBS 0.009165f
C552 B.n512 VSUBS 0.009165f
C553 B.n513 VSUBS 0.009165f
C554 B.n514 VSUBS 0.009165f
C555 B.n515 VSUBS 0.009165f
C556 B.n516 VSUBS 0.009165f
C557 B.n517 VSUBS 0.009165f
C558 B.n518 VSUBS 0.009165f
C559 B.n519 VSUBS 0.009165f
C560 B.n520 VSUBS 0.009165f
C561 B.n521 VSUBS 0.009165f
C562 B.n522 VSUBS 0.009165f
C563 B.n523 VSUBS 0.009165f
C564 B.n524 VSUBS 0.009165f
C565 B.n525 VSUBS 0.009165f
C566 B.n526 VSUBS 0.009165f
C567 B.n527 VSUBS 0.009165f
C568 B.n528 VSUBS 0.009165f
C569 B.n529 VSUBS 0.009165f
C570 B.n530 VSUBS 0.009165f
C571 B.n531 VSUBS 0.009165f
C572 B.n532 VSUBS 0.009165f
C573 B.n533 VSUBS 0.009165f
C574 B.n534 VSUBS 0.009165f
C575 B.n535 VSUBS 0.009165f
C576 B.n536 VSUBS 0.009165f
C577 B.n537 VSUBS 0.009165f
C578 B.n538 VSUBS 0.009165f
C579 B.n539 VSUBS 0.009165f
C580 B.n540 VSUBS 0.009165f
C581 B.n541 VSUBS 0.009165f
C582 B.n542 VSUBS 0.009165f
C583 B.n543 VSUBS 0.009165f
C584 B.n544 VSUBS 0.009165f
C585 B.n545 VSUBS 0.009165f
C586 B.n546 VSUBS 0.009165f
C587 B.n547 VSUBS 0.009165f
C588 B.n548 VSUBS 0.009165f
C589 B.n549 VSUBS 0.009165f
C590 B.n550 VSUBS 0.009165f
C591 B.n551 VSUBS 0.009165f
C592 B.n552 VSUBS 0.009165f
C593 B.n553 VSUBS 0.009165f
C594 B.n554 VSUBS 0.009165f
C595 B.n555 VSUBS 0.009165f
C596 B.n556 VSUBS 0.009165f
C597 B.n557 VSUBS 0.009165f
C598 B.n558 VSUBS 0.009165f
C599 B.n559 VSUBS 0.009165f
C600 B.n560 VSUBS 0.009165f
C601 B.n561 VSUBS 0.009165f
C602 B.n562 VSUBS 0.009165f
C603 B.n563 VSUBS 0.009165f
C604 B.n564 VSUBS 0.009165f
C605 B.n565 VSUBS 0.009165f
C606 B.n566 VSUBS 0.009165f
C607 B.n567 VSUBS 0.006335f
C608 B.n568 VSUBS 0.021235f
C609 B.n569 VSUBS 0.007413f
C610 B.n570 VSUBS 0.009165f
C611 B.n571 VSUBS 0.009165f
C612 B.n572 VSUBS 0.009165f
C613 B.n573 VSUBS 0.009165f
C614 B.n574 VSUBS 0.009165f
C615 B.n575 VSUBS 0.009165f
C616 B.n576 VSUBS 0.009165f
C617 B.n577 VSUBS 0.009165f
C618 B.n578 VSUBS 0.009165f
C619 B.n579 VSUBS 0.009165f
C620 B.n580 VSUBS 0.009165f
C621 B.n581 VSUBS 0.007413f
C622 B.n582 VSUBS 0.021235f
C623 B.n583 VSUBS 0.006335f
C624 B.n584 VSUBS 0.009165f
C625 B.n585 VSUBS 0.009165f
C626 B.n586 VSUBS 0.009165f
C627 B.n587 VSUBS 0.009165f
C628 B.n588 VSUBS 0.009165f
C629 B.n589 VSUBS 0.009165f
C630 B.n590 VSUBS 0.009165f
C631 B.n591 VSUBS 0.009165f
C632 B.n592 VSUBS 0.009165f
C633 B.n593 VSUBS 0.009165f
C634 B.n594 VSUBS 0.009165f
C635 B.n595 VSUBS 0.009165f
C636 B.n596 VSUBS 0.009165f
C637 B.n597 VSUBS 0.009165f
C638 B.n598 VSUBS 0.009165f
C639 B.n599 VSUBS 0.009165f
C640 B.n600 VSUBS 0.009165f
C641 B.n601 VSUBS 0.009165f
C642 B.n602 VSUBS 0.009165f
C643 B.n603 VSUBS 0.009165f
C644 B.n604 VSUBS 0.009165f
C645 B.n605 VSUBS 0.009165f
C646 B.n606 VSUBS 0.009165f
C647 B.n607 VSUBS 0.009165f
C648 B.n608 VSUBS 0.009165f
C649 B.n609 VSUBS 0.009165f
C650 B.n610 VSUBS 0.009165f
C651 B.n611 VSUBS 0.009165f
C652 B.n612 VSUBS 0.009165f
C653 B.n613 VSUBS 0.009165f
C654 B.n614 VSUBS 0.009165f
C655 B.n615 VSUBS 0.009165f
C656 B.n616 VSUBS 0.009165f
C657 B.n617 VSUBS 0.009165f
C658 B.n618 VSUBS 0.009165f
C659 B.n619 VSUBS 0.009165f
C660 B.n620 VSUBS 0.009165f
C661 B.n621 VSUBS 0.009165f
C662 B.n622 VSUBS 0.009165f
C663 B.n623 VSUBS 0.009165f
C664 B.n624 VSUBS 0.009165f
C665 B.n625 VSUBS 0.009165f
C666 B.n626 VSUBS 0.009165f
C667 B.n627 VSUBS 0.009165f
C668 B.n628 VSUBS 0.009165f
C669 B.n629 VSUBS 0.009165f
C670 B.n630 VSUBS 0.009165f
C671 B.n631 VSUBS 0.009165f
C672 B.n632 VSUBS 0.009165f
C673 B.n633 VSUBS 0.009165f
C674 B.n634 VSUBS 0.009165f
C675 B.n635 VSUBS 0.009165f
C676 B.n636 VSUBS 0.009165f
C677 B.n637 VSUBS 0.009165f
C678 B.n638 VSUBS 0.009165f
C679 B.n639 VSUBS 0.009165f
C680 B.n640 VSUBS 0.02129f
C681 B.n641 VSUBS 0.02129f
C682 B.n642 VSUBS 0.020493f
C683 B.n643 VSUBS 0.009165f
C684 B.n644 VSUBS 0.009165f
C685 B.n645 VSUBS 0.009165f
C686 B.n646 VSUBS 0.009165f
C687 B.n647 VSUBS 0.009165f
C688 B.n648 VSUBS 0.009165f
C689 B.n649 VSUBS 0.009165f
C690 B.n650 VSUBS 0.009165f
C691 B.n651 VSUBS 0.009165f
C692 B.n652 VSUBS 0.009165f
C693 B.n653 VSUBS 0.009165f
C694 B.n654 VSUBS 0.009165f
C695 B.n655 VSUBS 0.009165f
C696 B.n656 VSUBS 0.009165f
C697 B.n657 VSUBS 0.009165f
C698 B.n658 VSUBS 0.009165f
C699 B.n659 VSUBS 0.009165f
C700 B.n660 VSUBS 0.009165f
C701 B.n661 VSUBS 0.009165f
C702 B.n662 VSUBS 0.009165f
C703 B.n663 VSUBS 0.009165f
C704 B.n664 VSUBS 0.009165f
C705 B.n665 VSUBS 0.009165f
C706 B.n666 VSUBS 0.009165f
C707 B.n667 VSUBS 0.009165f
C708 B.n668 VSUBS 0.009165f
C709 B.n669 VSUBS 0.009165f
C710 B.n670 VSUBS 0.009165f
C711 B.n671 VSUBS 0.009165f
C712 B.n672 VSUBS 0.009165f
C713 B.n673 VSUBS 0.009165f
C714 B.n674 VSUBS 0.009165f
C715 B.n675 VSUBS 0.009165f
C716 B.n676 VSUBS 0.009165f
C717 B.n677 VSUBS 0.009165f
C718 B.n678 VSUBS 0.009165f
C719 B.n679 VSUBS 0.009165f
C720 B.n680 VSUBS 0.009165f
C721 B.n681 VSUBS 0.009165f
C722 B.n682 VSUBS 0.009165f
C723 B.n683 VSUBS 0.009165f
C724 B.n684 VSUBS 0.009165f
C725 B.n685 VSUBS 0.009165f
C726 B.n686 VSUBS 0.009165f
C727 B.n687 VSUBS 0.009165f
C728 B.n688 VSUBS 0.009165f
C729 B.n689 VSUBS 0.009165f
C730 B.n690 VSUBS 0.009165f
C731 B.n691 VSUBS 0.009165f
C732 B.n692 VSUBS 0.009165f
C733 B.n693 VSUBS 0.009165f
C734 B.n694 VSUBS 0.009165f
C735 B.n695 VSUBS 0.009165f
C736 B.n696 VSUBS 0.009165f
C737 B.n697 VSUBS 0.009165f
C738 B.n698 VSUBS 0.009165f
C739 B.n699 VSUBS 0.009165f
C740 B.n700 VSUBS 0.009165f
C741 B.n701 VSUBS 0.009165f
C742 B.n702 VSUBS 0.009165f
C743 B.n703 VSUBS 0.009165f
C744 B.n704 VSUBS 0.009165f
C745 B.n705 VSUBS 0.009165f
C746 B.n706 VSUBS 0.009165f
C747 B.n707 VSUBS 0.020753f
C748 VDD2.t3 VSUBS 2.44655f
C749 VDD2.t8 VSUBS 0.241781f
C750 VDD2.t1 VSUBS 0.241781f
C751 VDD2.n0 VSUBS 1.85702f
C752 VDD2.n1 VSUBS 1.44811f
C753 VDD2.t7 VSUBS 0.241781f
C754 VDD2.t2 VSUBS 0.241781f
C755 VDD2.n2 VSUBS 1.86961f
C756 VDD2.n3 VSUBS 2.88344f
C757 VDD2.t5 VSUBS 2.43027f
C758 VDD2.n4 VSUBS 3.26938f
C759 VDD2.t4 VSUBS 0.241781f
C760 VDD2.t0 VSUBS 0.241781f
C761 VDD2.n5 VSUBS 1.85703f
C762 VDD2.n6 VSUBS 0.709323f
C763 VDD2.t9 VSUBS 0.241781f
C764 VDD2.t6 VSUBS 0.241781f
C765 VDD2.n7 VSUBS 1.86957f
C766 VN.n0 VSUBS 0.036619f
C767 VN.t7 VSUBS 1.79858f
C768 VN.n1 VSUBS 0.048672f
C769 VN.n2 VSUBS 0.036619f
C770 VN.t2 VSUBS 1.79858f
C771 VN.n3 VSUBS 0.051711f
C772 VN.n4 VSUBS 0.036619f
C773 VN.t8 VSUBS 1.79858f
C774 VN.n5 VSUBS 0.054751f
C775 VN.t6 VSUBS 1.93621f
C776 VN.n6 VSUBS 0.736903f
C777 VN.t1 VSUBS 1.79858f
C778 VN.n7 VSUBS 0.721992f
C779 VN.n8 VSUBS 0.049133f
C780 VN.n9 VSUBS 0.235203f
C781 VN.n10 VSUBS 0.036619f
C782 VN.n11 VSUBS 0.036619f
C783 VN.n12 VSUBS 0.051711f
C784 VN.n13 VSUBS 0.051144f
C785 VN.n14 VSUBS 0.651751f
C786 VN.n15 VSUBS 0.051144f
C787 VN.n16 VSUBS 0.036619f
C788 VN.n17 VSUBS 0.036619f
C789 VN.n18 VSUBS 0.036619f
C790 VN.n19 VSUBS 0.054751f
C791 VN.n20 VSUBS 0.049133f
C792 VN.n21 VSUBS 0.651751f
C793 VN.n22 VSUBS 0.053156f
C794 VN.n23 VSUBS 0.036619f
C795 VN.n24 VSUBS 0.036619f
C796 VN.n25 VSUBS 0.036619f
C797 VN.n26 VSUBS 0.05779f
C798 VN.n27 VSUBS 0.047121f
C799 VN.n28 VSUBS 0.734007f
C800 VN.n29 VSUBS 0.036153f
C801 VN.n30 VSUBS 0.036619f
C802 VN.t4 VSUBS 1.79858f
C803 VN.n31 VSUBS 0.048672f
C804 VN.n32 VSUBS 0.036619f
C805 VN.t5 VSUBS 1.79858f
C806 VN.n33 VSUBS 0.051711f
C807 VN.n34 VSUBS 0.036619f
C808 VN.t9 VSUBS 1.79858f
C809 VN.n35 VSUBS 0.054751f
C810 VN.t3 VSUBS 1.93621f
C811 VN.n36 VSUBS 0.736903f
C812 VN.t0 VSUBS 1.79858f
C813 VN.n37 VSUBS 0.721992f
C814 VN.n38 VSUBS 0.049133f
C815 VN.n39 VSUBS 0.235203f
C816 VN.n40 VSUBS 0.036619f
C817 VN.n41 VSUBS 0.036619f
C818 VN.n42 VSUBS 0.051711f
C819 VN.n43 VSUBS 0.051144f
C820 VN.n44 VSUBS 0.651751f
C821 VN.n45 VSUBS 0.051144f
C822 VN.n46 VSUBS 0.036619f
C823 VN.n47 VSUBS 0.036619f
C824 VN.n48 VSUBS 0.036619f
C825 VN.n49 VSUBS 0.054751f
C826 VN.n50 VSUBS 0.049133f
C827 VN.n51 VSUBS 0.651751f
C828 VN.n52 VSUBS 0.053156f
C829 VN.n53 VSUBS 0.036619f
C830 VN.n54 VSUBS 0.036619f
C831 VN.n55 VSUBS 0.036619f
C832 VN.n56 VSUBS 0.05779f
C833 VN.n57 VSUBS 0.047121f
C834 VN.n58 VSUBS 0.734007f
C835 VN.n59 VSUBS 1.84896f
C836 VDD1.t6 VSUBS 2.45667f
C837 VDD1.t8 VSUBS 0.242779f
C838 VDD1.t2 VSUBS 0.242779f
C839 VDD1.n0 VSUBS 1.8647f
C840 VDD1.n1 VSUBS 1.46252f
C841 VDD1.t0 VSUBS 2.45665f
C842 VDD1.t7 VSUBS 0.242779f
C843 VDD1.t1 VSUBS 0.242779f
C844 VDD1.n2 VSUBS 1.86469f
C845 VDD1.n3 VSUBS 1.45409f
C846 VDD1.t5 VSUBS 0.242779f
C847 VDD1.t3 VSUBS 0.242779f
C848 VDD1.n4 VSUBS 1.87733f
C849 VDD1.n5 VSUBS 3.00622f
C850 VDD1.t4 VSUBS 0.242779f
C851 VDD1.t9 VSUBS 0.242779f
C852 VDD1.n6 VSUBS 1.86469f
C853 VDD1.n7 VSUBS 3.29766f
C854 VTAIL.t0 VSUBS 0.249998f
C855 VTAIL.t5 VSUBS 0.249998f
C856 VTAIL.n0 VSUBS 1.76943f
C857 VTAIL.n1 VSUBS 0.888582f
C858 VTAIL.t11 VSUBS 2.34513f
C859 VTAIL.n2 VSUBS 1.02859f
C860 VTAIL.t17 VSUBS 0.249998f
C861 VTAIL.t13 VSUBS 0.249998f
C862 VTAIL.n3 VSUBS 1.76943f
C863 VTAIL.n4 VSUBS 0.957561f
C864 VTAIL.t10 VSUBS 0.249998f
C865 VTAIL.t12 VSUBS 0.249998f
C866 VTAIL.n5 VSUBS 1.76943f
C867 VTAIL.n6 VSUBS 2.3834f
C868 VTAIL.t9 VSUBS 0.249998f
C869 VTAIL.t2 VSUBS 0.249998f
C870 VTAIL.n7 VSUBS 1.76944f
C871 VTAIL.n8 VSUBS 2.3834f
C872 VTAIL.t3 VSUBS 0.249998f
C873 VTAIL.t4 VSUBS 0.249998f
C874 VTAIL.n9 VSUBS 1.76944f
C875 VTAIL.n10 VSUBS 0.957553f
C876 VTAIL.t7 VSUBS 2.34514f
C877 VTAIL.n11 VSUBS 1.02858f
C878 VTAIL.t18 VSUBS 0.249998f
C879 VTAIL.t19 VSUBS 0.249998f
C880 VTAIL.n12 VSUBS 1.76944f
C881 VTAIL.n13 VSUBS 0.922466f
C882 VTAIL.t16 VSUBS 0.249998f
C883 VTAIL.t14 VSUBS 0.249998f
C884 VTAIL.n14 VSUBS 1.76944f
C885 VTAIL.n15 VSUBS 0.957553f
C886 VTAIL.t15 VSUBS 2.34513f
C887 VTAIL.n16 VSUBS 2.33243f
C888 VTAIL.t8 VSUBS 2.34513f
C889 VTAIL.n17 VSUBS 2.33243f
C890 VTAIL.t1 VSUBS 0.249998f
C891 VTAIL.t6 VSUBS 0.249998f
C892 VTAIL.n18 VSUBS 1.76943f
C893 VTAIL.n19 VSUBS 0.834356f
C894 VP.n0 VSUBS 0.037494f
C895 VP.t6 VSUBS 1.84156f
C896 VP.n1 VSUBS 0.049835f
C897 VP.n2 VSUBS 0.037494f
C898 VP.t4 VSUBS 1.84156f
C899 VP.n3 VSUBS 0.052947f
C900 VP.n4 VSUBS 0.037494f
C901 VP.t8 VSUBS 1.84156f
C902 VP.n5 VSUBS 0.056059f
C903 VP.n6 VSUBS 0.037494f
C904 VP.t2 VSUBS 1.84156f
C905 VP.n7 VSUBS 0.059171f
C906 VP.n8 VSUBS 0.037494f
C907 VP.t0 VSUBS 1.84156f
C908 VP.n9 VSUBS 0.049835f
C909 VP.n10 VSUBS 0.037494f
C910 VP.t5 VSUBS 1.84156f
C911 VP.n11 VSUBS 0.052947f
C912 VP.n12 VSUBS 0.037494f
C913 VP.t7 VSUBS 1.84156f
C914 VP.n13 VSUBS 0.056059f
C915 VP.t3 VSUBS 1.98247f
C916 VP.n14 VSUBS 0.754511f
C917 VP.t1 VSUBS 1.84156f
C918 VP.n15 VSUBS 0.739244f
C919 VP.n16 VSUBS 0.050307f
C920 VP.n17 VSUBS 0.240823f
C921 VP.n18 VSUBS 0.037494f
C922 VP.n19 VSUBS 0.037494f
C923 VP.n20 VSUBS 0.052947f
C924 VP.n21 VSUBS 0.052366f
C925 VP.n22 VSUBS 0.667325f
C926 VP.n23 VSUBS 0.052366f
C927 VP.n24 VSUBS 0.037494f
C928 VP.n25 VSUBS 0.037494f
C929 VP.n26 VSUBS 0.037494f
C930 VP.n27 VSUBS 0.056059f
C931 VP.n28 VSUBS 0.050307f
C932 VP.n29 VSUBS 0.667325f
C933 VP.n30 VSUBS 0.054426f
C934 VP.n31 VSUBS 0.037494f
C935 VP.n32 VSUBS 0.037494f
C936 VP.n33 VSUBS 0.037494f
C937 VP.n34 VSUBS 0.059171f
C938 VP.n35 VSUBS 0.048248f
C939 VP.n36 VSUBS 0.751546f
C940 VP.n37 VSUBS 1.86869f
C941 VP.n38 VSUBS 1.89739f
C942 VP.t9 VSUBS 1.84156f
C943 VP.n39 VSUBS 0.751546f
C944 VP.n40 VSUBS 0.048248f
C945 VP.n41 VSUBS 0.037494f
C946 VP.n42 VSUBS 0.037494f
C947 VP.n43 VSUBS 0.037494f
C948 VP.n44 VSUBS 0.049835f
C949 VP.n45 VSUBS 0.054426f
C950 VP.n46 VSUBS 0.667325f
C951 VP.n47 VSUBS 0.050307f
C952 VP.n48 VSUBS 0.037494f
C953 VP.n49 VSUBS 0.037494f
C954 VP.n50 VSUBS 0.037494f
C955 VP.n51 VSUBS 0.052947f
C956 VP.n52 VSUBS 0.052366f
C957 VP.n53 VSUBS 0.667325f
C958 VP.n54 VSUBS 0.052366f
C959 VP.n55 VSUBS 0.037494f
C960 VP.n56 VSUBS 0.037494f
C961 VP.n57 VSUBS 0.037494f
C962 VP.n58 VSUBS 0.056059f
C963 VP.n59 VSUBS 0.050307f
C964 VP.n60 VSUBS 0.667325f
C965 VP.n61 VSUBS 0.054426f
C966 VP.n62 VSUBS 0.037494f
C967 VP.n63 VSUBS 0.037494f
C968 VP.n64 VSUBS 0.037494f
C969 VP.n65 VSUBS 0.059171f
C970 VP.n66 VSUBS 0.048248f
C971 VP.n67 VSUBS 0.751546f
C972 VP.n68 VSUBS 0.037017f
.ends

