* NGSPICE file created from diff_pair_sample_0392.ext - technology: sky130A

.subckt diff_pair_sample_0392 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t6 VN.t0 VDD2.t0 w_n2656_n2314# sky130_fd_pr__pfet_01v8 ad=2.6247 pd=14.24 as=1.11045 ps=7.06 w=6.73 l=2.48
X1 VTAIL.t2 VP.t0 VDD1.t3 w_n2656_n2314# sky130_fd_pr__pfet_01v8 ad=2.6247 pd=14.24 as=1.11045 ps=7.06 w=6.73 l=2.48
X2 VTAIL.t5 VN.t1 VDD2.t2 w_n2656_n2314# sky130_fd_pr__pfet_01v8 ad=2.6247 pd=14.24 as=1.11045 ps=7.06 w=6.73 l=2.48
X3 VDD1.t2 VP.t1 VTAIL.t7 w_n2656_n2314# sky130_fd_pr__pfet_01v8 ad=1.11045 pd=7.06 as=2.6247 ps=14.24 w=6.73 l=2.48
X4 B.t11 B.t9 B.t10 w_n2656_n2314# sky130_fd_pr__pfet_01v8 ad=2.6247 pd=14.24 as=0 ps=0 w=6.73 l=2.48
X5 VDD2.t1 VN.t2 VTAIL.t4 w_n2656_n2314# sky130_fd_pr__pfet_01v8 ad=1.11045 pd=7.06 as=2.6247 ps=14.24 w=6.73 l=2.48
X6 B.t8 B.t6 B.t7 w_n2656_n2314# sky130_fd_pr__pfet_01v8 ad=2.6247 pd=14.24 as=0 ps=0 w=6.73 l=2.48
X7 VDD2.t3 VN.t3 VTAIL.t3 w_n2656_n2314# sky130_fd_pr__pfet_01v8 ad=1.11045 pd=7.06 as=2.6247 ps=14.24 w=6.73 l=2.48
X8 VTAIL.t0 VP.t2 VDD1.t1 w_n2656_n2314# sky130_fd_pr__pfet_01v8 ad=2.6247 pd=14.24 as=1.11045 ps=7.06 w=6.73 l=2.48
X9 VDD1.t0 VP.t3 VTAIL.t1 w_n2656_n2314# sky130_fd_pr__pfet_01v8 ad=1.11045 pd=7.06 as=2.6247 ps=14.24 w=6.73 l=2.48
X10 B.t5 B.t3 B.t4 w_n2656_n2314# sky130_fd_pr__pfet_01v8 ad=2.6247 pd=14.24 as=0 ps=0 w=6.73 l=2.48
X11 B.t2 B.t0 B.t1 w_n2656_n2314# sky130_fd_pr__pfet_01v8 ad=2.6247 pd=14.24 as=0 ps=0 w=6.73 l=2.48
R0 VN.n0 VN.t1 100.665
R1 VN.n1 VN.t2 100.665
R2 VN.n0 VN.t3 99.9113
R3 VN.n1 VN.t0 99.9113
R4 VN VN.n1 46.7318
R5 VN VN.n0 4.56892
R6 VDD2.n2 VDD2.n0 125.376
R7 VDD2.n2 VDD2.n1 88.5927
R8 VDD2.n1 VDD2.t0 4.83037
R9 VDD2.n1 VDD2.t1 4.83037
R10 VDD2.n0 VDD2.t2 4.83037
R11 VDD2.n0 VDD2.t3 4.83037
R12 VDD2 VDD2.n2 0.0586897
R13 VTAIL.n282 VTAIL.n252 756.745
R14 VTAIL.n30 VTAIL.n0 756.745
R15 VTAIL.n66 VTAIL.n36 756.745
R16 VTAIL.n102 VTAIL.n72 756.745
R17 VTAIL.n246 VTAIL.n216 756.745
R18 VTAIL.n210 VTAIL.n180 756.745
R19 VTAIL.n174 VTAIL.n144 756.745
R20 VTAIL.n138 VTAIL.n108 756.745
R21 VTAIL.n265 VTAIL.n264 585
R22 VTAIL.n267 VTAIL.n266 585
R23 VTAIL.n260 VTAIL.n259 585
R24 VTAIL.n273 VTAIL.n272 585
R25 VTAIL.n275 VTAIL.n274 585
R26 VTAIL.n256 VTAIL.n255 585
R27 VTAIL.n281 VTAIL.n280 585
R28 VTAIL.n283 VTAIL.n282 585
R29 VTAIL.n13 VTAIL.n12 585
R30 VTAIL.n15 VTAIL.n14 585
R31 VTAIL.n8 VTAIL.n7 585
R32 VTAIL.n21 VTAIL.n20 585
R33 VTAIL.n23 VTAIL.n22 585
R34 VTAIL.n4 VTAIL.n3 585
R35 VTAIL.n29 VTAIL.n28 585
R36 VTAIL.n31 VTAIL.n30 585
R37 VTAIL.n49 VTAIL.n48 585
R38 VTAIL.n51 VTAIL.n50 585
R39 VTAIL.n44 VTAIL.n43 585
R40 VTAIL.n57 VTAIL.n56 585
R41 VTAIL.n59 VTAIL.n58 585
R42 VTAIL.n40 VTAIL.n39 585
R43 VTAIL.n65 VTAIL.n64 585
R44 VTAIL.n67 VTAIL.n66 585
R45 VTAIL.n85 VTAIL.n84 585
R46 VTAIL.n87 VTAIL.n86 585
R47 VTAIL.n80 VTAIL.n79 585
R48 VTAIL.n93 VTAIL.n92 585
R49 VTAIL.n95 VTAIL.n94 585
R50 VTAIL.n76 VTAIL.n75 585
R51 VTAIL.n101 VTAIL.n100 585
R52 VTAIL.n103 VTAIL.n102 585
R53 VTAIL.n247 VTAIL.n246 585
R54 VTAIL.n245 VTAIL.n244 585
R55 VTAIL.n220 VTAIL.n219 585
R56 VTAIL.n239 VTAIL.n238 585
R57 VTAIL.n237 VTAIL.n236 585
R58 VTAIL.n224 VTAIL.n223 585
R59 VTAIL.n231 VTAIL.n230 585
R60 VTAIL.n229 VTAIL.n228 585
R61 VTAIL.n211 VTAIL.n210 585
R62 VTAIL.n209 VTAIL.n208 585
R63 VTAIL.n184 VTAIL.n183 585
R64 VTAIL.n203 VTAIL.n202 585
R65 VTAIL.n201 VTAIL.n200 585
R66 VTAIL.n188 VTAIL.n187 585
R67 VTAIL.n195 VTAIL.n194 585
R68 VTAIL.n193 VTAIL.n192 585
R69 VTAIL.n175 VTAIL.n174 585
R70 VTAIL.n173 VTAIL.n172 585
R71 VTAIL.n148 VTAIL.n147 585
R72 VTAIL.n167 VTAIL.n166 585
R73 VTAIL.n165 VTAIL.n164 585
R74 VTAIL.n152 VTAIL.n151 585
R75 VTAIL.n159 VTAIL.n158 585
R76 VTAIL.n157 VTAIL.n156 585
R77 VTAIL.n139 VTAIL.n138 585
R78 VTAIL.n137 VTAIL.n136 585
R79 VTAIL.n112 VTAIL.n111 585
R80 VTAIL.n131 VTAIL.n130 585
R81 VTAIL.n129 VTAIL.n128 585
R82 VTAIL.n116 VTAIL.n115 585
R83 VTAIL.n123 VTAIL.n122 585
R84 VTAIL.n121 VTAIL.n120 585
R85 VTAIL.n263 VTAIL.t3 327.514
R86 VTAIL.n11 VTAIL.t5 327.514
R87 VTAIL.n47 VTAIL.t1 327.514
R88 VTAIL.n83 VTAIL.t0 327.514
R89 VTAIL.n227 VTAIL.t7 327.514
R90 VTAIL.n191 VTAIL.t2 327.514
R91 VTAIL.n155 VTAIL.t4 327.514
R92 VTAIL.n119 VTAIL.t6 327.514
R93 VTAIL.n266 VTAIL.n265 171.744
R94 VTAIL.n266 VTAIL.n259 171.744
R95 VTAIL.n273 VTAIL.n259 171.744
R96 VTAIL.n274 VTAIL.n273 171.744
R97 VTAIL.n274 VTAIL.n255 171.744
R98 VTAIL.n281 VTAIL.n255 171.744
R99 VTAIL.n282 VTAIL.n281 171.744
R100 VTAIL.n14 VTAIL.n13 171.744
R101 VTAIL.n14 VTAIL.n7 171.744
R102 VTAIL.n21 VTAIL.n7 171.744
R103 VTAIL.n22 VTAIL.n21 171.744
R104 VTAIL.n22 VTAIL.n3 171.744
R105 VTAIL.n29 VTAIL.n3 171.744
R106 VTAIL.n30 VTAIL.n29 171.744
R107 VTAIL.n50 VTAIL.n49 171.744
R108 VTAIL.n50 VTAIL.n43 171.744
R109 VTAIL.n57 VTAIL.n43 171.744
R110 VTAIL.n58 VTAIL.n57 171.744
R111 VTAIL.n58 VTAIL.n39 171.744
R112 VTAIL.n65 VTAIL.n39 171.744
R113 VTAIL.n66 VTAIL.n65 171.744
R114 VTAIL.n86 VTAIL.n85 171.744
R115 VTAIL.n86 VTAIL.n79 171.744
R116 VTAIL.n93 VTAIL.n79 171.744
R117 VTAIL.n94 VTAIL.n93 171.744
R118 VTAIL.n94 VTAIL.n75 171.744
R119 VTAIL.n101 VTAIL.n75 171.744
R120 VTAIL.n102 VTAIL.n101 171.744
R121 VTAIL.n246 VTAIL.n245 171.744
R122 VTAIL.n245 VTAIL.n219 171.744
R123 VTAIL.n238 VTAIL.n219 171.744
R124 VTAIL.n238 VTAIL.n237 171.744
R125 VTAIL.n237 VTAIL.n223 171.744
R126 VTAIL.n230 VTAIL.n223 171.744
R127 VTAIL.n230 VTAIL.n229 171.744
R128 VTAIL.n210 VTAIL.n209 171.744
R129 VTAIL.n209 VTAIL.n183 171.744
R130 VTAIL.n202 VTAIL.n183 171.744
R131 VTAIL.n202 VTAIL.n201 171.744
R132 VTAIL.n201 VTAIL.n187 171.744
R133 VTAIL.n194 VTAIL.n187 171.744
R134 VTAIL.n194 VTAIL.n193 171.744
R135 VTAIL.n174 VTAIL.n173 171.744
R136 VTAIL.n173 VTAIL.n147 171.744
R137 VTAIL.n166 VTAIL.n147 171.744
R138 VTAIL.n166 VTAIL.n165 171.744
R139 VTAIL.n165 VTAIL.n151 171.744
R140 VTAIL.n158 VTAIL.n151 171.744
R141 VTAIL.n158 VTAIL.n157 171.744
R142 VTAIL.n138 VTAIL.n137 171.744
R143 VTAIL.n137 VTAIL.n111 171.744
R144 VTAIL.n130 VTAIL.n111 171.744
R145 VTAIL.n130 VTAIL.n129 171.744
R146 VTAIL.n129 VTAIL.n115 171.744
R147 VTAIL.n122 VTAIL.n115 171.744
R148 VTAIL.n122 VTAIL.n121 171.744
R149 VTAIL.n265 VTAIL.t3 85.8723
R150 VTAIL.n13 VTAIL.t5 85.8723
R151 VTAIL.n49 VTAIL.t1 85.8723
R152 VTAIL.n85 VTAIL.t0 85.8723
R153 VTAIL.n229 VTAIL.t7 85.8723
R154 VTAIL.n193 VTAIL.t2 85.8723
R155 VTAIL.n157 VTAIL.t4 85.8723
R156 VTAIL.n121 VTAIL.t6 85.8723
R157 VTAIL.n287 VTAIL.n286 32.3793
R158 VTAIL.n35 VTAIL.n34 32.3793
R159 VTAIL.n71 VTAIL.n70 32.3793
R160 VTAIL.n107 VTAIL.n106 32.3793
R161 VTAIL.n251 VTAIL.n250 32.3793
R162 VTAIL.n215 VTAIL.n214 32.3793
R163 VTAIL.n179 VTAIL.n178 32.3793
R164 VTAIL.n143 VTAIL.n142 32.3793
R165 VTAIL.n287 VTAIL.n251 20.591
R166 VTAIL.n143 VTAIL.n107 20.591
R167 VTAIL.n264 VTAIL.n263 16.3884
R168 VTAIL.n12 VTAIL.n11 16.3884
R169 VTAIL.n48 VTAIL.n47 16.3884
R170 VTAIL.n84 VTAIL.n83 16.3884
R171 VTAIL.n228 VTAIL.n227 16.3884
R172 VTAIL.n192 VTAIL.n191 16.3884
R173 VTAIL.n156 VTAIL.n155 16.3884
R174 VTAIL.n120 VTAIL.n119 16.3884
R175 VTAIL.n267 VTAIL.n262 12.8005
R176 VTAIL.n15 VTAIL.n10 12.8005
R177 VTAIL.n51 VTAIL.n46 12.8005
R178 VTAIL.n87 VTAIL.n82 12.8005
R179 VTAIL.n231 VTAIL.n226 12.8005
R180 VTAIL.n195 VTAIL.n190 12.8005
R181 VTAIL.n159 VTAIL.n154 12.8005
R182 VTAIL.n123 VTAIL.n118 12.8005
R183 VTAIL.n268 VTAIL.n260 12.0247
R184 VTAIL.n16 VTAIL.n8 12.0247
R185 VTAIL.n52 VTAIL.n44 12.0247
R186 VTAIL.n88 VTAIL.n80 12.0247
R187 VTAIL.n232 VTAIL.n224 12.0247
R188 VTAIL.n196 VTAIL.n188 12.0247
R189 VTAIL.n160 VTAIL.n152 12.0247
R190 VTAIL.n124 VTAIL.n116 12.0247
R191 VTAIL.n272 VTAIL.n271 11.249
R192 VTAIL.n20 VTAIL.n19 11.249
R193 VTAIL.n56 VTAIL.n55 11.249
R194 VTAIL.n92 VTAIL.n91 11.249
R195 VTAIL.n236 VTAIL.n235 11.249
R196 VTAIL.n200 VTAIL.n199 11.249
R197 VTAIL.n164 VTAIL.n163 11.249
R198 VTAIL.n128 VTAIL.n127 11.249
R199 VTAIL.n275 VTAIL.n258 10.4732
R200 VTAIL.n23 VTAIL.n6 10.4732
R201 VTAIL.n59 VTAIL.n42 10.4732
R202 VTAIL.n95 VTAIL.n78 10.4732
R203 VTAIL.n239 VTAIL.n222 10.4732
R204 VTAIL.n203 VTAIL.n186 10.4732
R205 VTAIL.n167 VTAIL.n150 10.4732
R206 VTAIL.n131 VTAIL.n114 10.4732
R207 VTAIL.n276 VTAIL.n256 9.69747
R208 VTAIL.n24 VTAIL.n4 9.69747
R209 VTAIL.n60 VTAIL.n40 9.69747
R210 VTAIL.n96 VTAIL.n76 9.69747
R211 VTAIL.n240 VTAIL.n220 9.69747
R212 VTAIL.n204 VTAIL.n184 9.69747
R213 VTAIL.n168 VTAIL.n148 9.69747
R214 VTAIL.n132 VTAIL.n112 9.69747
R215 VTAIL.n286 VTAIL.n285 9.45567
R216 VTAIL.n34 VTAIL.n33 9.45567
R217 VTAIL.n70 VTAIL.n69 9.45567
R218 VTAIL.n106 VTAIL.n105 9.45567
R219 VTAIL.n250 VTAIL.n249 9.45567
R220 VTAIL.n214 VTAIL.n213 9.45567
R221 VTAIL.n178 VTAIL.n177 9.45567
R222 VTAIL.n142 VTAIL.n141 9.45567
R223 VTAIL.n254 VTAIL.n253 9.3005
R224 VTAIL.n279 VTAIL.n278 9.3005
R225 VTAIL.n277 VTAIL.n276 9.3005
R226 VTAIL.n258 VTAIL.n257 9.3005
R227 VTAIL.n271 VTAIL.n270 9.3005
R228 VTAIL.n269 VTAIL.n268 9.3005
R229 VTAIL.n262 VTAIL.n261 9.3005
R230 VTAIL.n285 VTAIL.n284 9.3005
R231 VTAIL.n2 VTAIL.n1 9.3005
R232 VTAIL.n27 VTAIL.n26 9.3005
R233 VTAIL.n25 VTAIL.n24 9.3005
R234 VTAIL.n6 VTAIL.n5 9.3005
R235 VTAIL.n19 VTAIL.n18 9.3005
R236 VTAIL.n17 VTAIL.n16 9.3005
R237 VTAIL.n10 VTAIL.n9 9.3005
R238 VTAIL.n33 VTAIL.n32 9.3005
R239 VTAIL.n38 VTAIL.n37 9.3005
R240 VTAIL.n63 VTAIL.n62 9.3005
R241 VTAIL.n61 VTAIL.n60 9.3005
R242 VTAIL.n42 VTAIL.n41 9.3005
R243 VTAIL.n55 VTAIL.n54 9.3005
R244 VTAIL.n53 VTAIL.n52 9.3005
R245 VTAIL.n46 VTAIL.n45 9.3005
R246 VTAIL.n69 VTAIL.n68 9.3005
R247 VTAIL.n74 VTAIL.n73 9.3005
R248 VTAIL.n99 VTAIL.n98 9.3005
R249 VTAIL.n97 VTAIL.n96 9.3005
R250 VTAIL.n78 VTAIL.n77 9.3005
R251 VTAIL.n91 VTAIL.n90 9.3005
R252 VTAIL.n89 VTAIL.n88 9.3005
R253 VTAIL.n82 VTAIL.n81 9.3005
R254 VTAIL.n105 VTAIL.n104 9.3005
R255 VTAIL.n249 VTAIL.n248 9.3005
R256 VTAIL.n218 VTAIL.n217 9.3005
R257 VTAIL.n243 VTAIL.n242 9.3005
R258 VTAIL.n241 VTAIL.n240 9.3005
R259 VTAIL.n222 VTAIL.n221 9.3005
R260 VTAIL.n235 VTAIL.n234 9.3005
R261 VTAIL.n233 VTAIL.n232 9.3005
R262 VTAIL.n226 VTAIL.n225 9.3005
R263 VTAIL.n213 VTAIL.n212 9.3005
R264 VTAIL.n182 VTAIL.n181 9.3005
R265 VTAIL.n207 VTAIL.n206 9.3005
R266 VTAIL.n205 VTAIL.n204 9.3005
R267 VTAIL.n186 VTAIL.n185 9.3005
R268 VTAIL.n199 VTAIL.n198 9.3005
R269 VTAIL.n197 VTAIL.n196 9.3005
R270 VTAIL.n190 VTAIL.n189 9.3005
R271 VTAIL.n177 VTAIL.n176 9.3005
R272 VTAIL.n146 VTAIL.n145 9.3005
R273 VTAIL.n171 VTAIL.n170 9.3005
R274 VTAIL.n169 VTAIL.n168 9.3005
R275 VTAIL.n150 VTAIL.n149 9.3005
R276 VTAIL.n163 VTAIL.n162 9.3005
R277 VTAIL.n161 VTAIL.n160 9.3005
R278 VTAIL.n154 VTAIL.n153 9.3005
R279 VTAIL.n141 VTAIL.n140 9.3005
R280 VTAIL.n110 VTAIL.n109 9.3005
R281 VTAIL.n135 VTAIL.n134 9.3005
R282 VTAIL.n133 VTAIL.n132 9.3005
R283 VTAIL.n114 VTAIL.n113 9.3005
R284 VTAIL.n127 VTAIL.n126 9.3005
R285 VTAIL.n125 VTAIL.n124 9.3005
R286 VTAIL.n118 VTAIL.n117 9.3005
R287 VTAIL.n280 VTAIL.n279 8.92171
R288 VTAIL.n28 VTAIL.n27 8.92171
R289 VTAIL.n64 VTAIL.n63 8.92171
R290 VTAIL.n100 VTAIL.n99 8.92171
R291 VTAIL.n244 VTAIL.n243 8.92171
R292 VTAIL.n208 VTAIL.n207 8.92171
R293 VTAIL.n172 VTAIL.n171 8.92171
R294 VTAIL.n136 VTAIL.n135 8.92171
R295 VTAIL.n283 VTAIL.n254 8.14595
R296 VTAIL.n31 VTAIL.n2 8.14595
R297 VTAIL.n67 VTAIL.n38 8.14595
R298 VTAIL.n103 VTAIL.n74 8.14595
R299 VTAIL.n247 VTAIL.n218 8.14595
R300 VTAIL.n211 VTAIL.n182 8.14595
R301 VTAIL.n175 VTAIL.n146 8.14595
R302 VTAIL.n139 VTAIL.n110 8.14595
R303 VTAIL.n284 VTAIL.n252 7.3702
R304 VTAIL.n32 VTAIL.n0 7.3702
R305 VTAIL.n68 VTAIL.n36 7.3702
R306 VTAIL.n104 VTAIL.n72 7.3702
R307 VTAIL.n248 VTAIL.n216 7.3702
R308 VTAIL.n212 VTAIL.n180 7.3702
R309 VTAIL.n176 VTAIL.n144 7.3702
R310 VTAIL.n140 VTAIL.n108 7.3702
R311 VTAIL.n286 VTAIL.n252 6.59444
R312 VTAIL.n34 VTAIL.n0 6.59444
R313 VTAIL.n70 VTAIL.n36 6.59444
R314 VTAIL.n106 VTAIL.n72 6.59444
R315 VTAIL.n250 VTAIL.n216 6.59444
R316 VTAIL.n214 VTAIL.n180 6.59444
R317 VTAIL.n178 VTAIL.n144 6.59444
R318 VTAIL.n142 VTAIL.n108 6.59444
R319 VTAIL.n284 VTAIL.n283 5.81868
R320 VTAIL.n32 VTAIL.n31 5.81868
R321 VTAIL.n68 VTAIL.n67 5.81868
R322 VTAIL.n104 VTAIL.n103 5.81868
R323 VTAIL.n248 VTAIL.n247 5.81868
R324 VTAIL.n212 VTAIL.n211 5.81868
R325 VTAIL.n176 VTAIL.n175 5.81868
R326 VTAIL.n140 VTAIL.n139 5.81868
R327 VTAIL.n280 VTAIL.n254 5.04292
R328 VTAIL.n28 VTAIL.n2 5.04292
R329 VTAIL.n64 VTAIL.n38 5.04292
R330 VTAIL.n100 VTAIL.n74 5.04292
R331 VTAIL.n244 VTAIL.n218 5.04292
R332 VTAIL.n208 VTAIL.n182 5.04292
R333 VTAIL.n172 VTAIL.n146 5.04292
R334 VTAIL.n136 VTAIL.n110 5.04292
R335 VTAIL.n279 VTAIL.n256 4.26717
R336 VTAIL.n27 VTAIL.n4 4.26717
R337 VTAIL.n63 VTAIL.n40 4.26717
R338 VTAIL.n99 VTAIL.n76 4.26717
R339 VTAIL.n243 VTAIL.n220 4.26717
R340 VTAIL.n207 VTAIL.n184 4.26717
R341 VTAIL.n171 VTAIL.n148 4.26717
R342 VTAIL.n135 VTAIL.n112 4.26717
R343 VTAIL.n263 VTAIL.n261 3.71088
R344 VTAIL.n11 VTAIL.n9 3.71088
R345 VTAIL.n47 VTAIL.n45 3.71088
R346 VTAIL.n83 VTAIL.n81 3.71088
R347 VTAIL.n227 VTAIL.n225 3.71088
R348 VTAIL.n191 VTAIL.n189 3.71088
R349 VTAIL.n155 VTAIL.n153 3.71088
R350 VTAIL.n119 VTAIL.n117 3.71088
R351 VTAIL.n276 VTAIL.n275 3.49141
R352 VTAIL.n24 VTAIL.n23 3.49141
R353 VTAIL.n60 VTAIL.n59 3.49141
R354 VTAIL.n96 VTAIL.n95 3.49141
R355 VTAIL.n240 VTAIL.n239 3.49141
R356 VTAIL.n204 VTAIL.n203 3.49141
R357 VTAIL.n168 VTAIL.n167 3.49141
R358 VTAIL.n132 VTAIL.n131 3.49141
R359 VTAIL.n272 VTAIL.n258 2.71565
R360 VTAIL.n20 VTAIL.n6 2.71565
R361 VTAIL.n56 VTAIL.n42 2.71565
R362 VTAIL.n92 VTAIL.n78 2.71565
R363 VTAIL.n236 VTAIL.n222 2.71565
R364 VTAIL.n200 VTAIL.n186 2.71565
R365 VTAIL.n164 VTAIL.n150 2.71565
R366 VTAIL.n128 VTAIL.n114 2.71565
R367 VTAIL.n179 VTAIL.n143 2.42291
R368 VTAIL.n251 VTAIL.n215 2.42291
R369 VTAIL.n107 VTAIL.n71 2.42291
R370 VTAIL.n271 VTAIL.n260 1.93989
R371 VTAIL.n19 VTAIL.n8 1.93989
R372 VTAIL.n55 VTAIL.n44 1.93989
R373 VTAIL.n91 VTAIL.n80 1.93989
R374 VTAIL.n235 VTAIL.n224 1.93989
R375 VTAIL.n199 VTAIL.n188 1.93989
R376 VTAIL.n163 VTAIL.n152 1.93989
R377 VTAIL.n127 VTAIL.n116 1.93989
R378 VTAIL VTAIL.n35 1.2699
R379 VTAIL.n268 VTAIL.n267 1.16414
R380 VTAIL.n16 VTAIL.n15 1.16414
R381 VTAIL.n52 VTAIL.n51 1.16414
R382 VTAIL.n88 VTAIL.n87 1.16414
R383 VTAIL.n232 VTAIL.n231 1.16414
R384 VTAIL.n196 VTAIL.n195 1.16414
R385 VTAIL.n160 VTAIL.n159 1.16414
R386 VTAIL.n124 VTAIL.n123 1.16414
R387 VTAIL VTAIL.n287 1.15352
R388 VTAIL.n215 VTAIL.n179 0.470328
R389 VTAIL.n71 VTAIL.n35 0.470328
R390 VTAIL.n264 VTAIL.n262 0.388379
R391 VTAIL.n12 VTAIL.n10 0.388379
R392 VTAIL.n48 VTAIL.n46 0.388379
R393 VTAIL.n84 VTAIL.n82 0.388379
R394 VTAIL.n228 VTAIL.n226 0.388379
R395 VTAIL.n192 VTAIL.n190 0.388379
R396 VTAIL.n156 VTAIL.n154 0.388379
R397 VTAIL.n120 VTAIL.n118 0.388379
R398 VTAIL.n269 VTAIL.n261 0.155672
R399 VTAIL.n270 VTAIL.n269 0.155672
R400 VTAIL.n270 VTAIL.n257 0.155672
R401 VTAIL.n277 VTAIL.n257 0.155672
R402 VTAIL.n278 VTAIL.n277 0.155672
R403 VTAIL.n278 VTAIL.n253 0.155672
R404 VTAIL.n285 VTAIL.n253 0.155672
R405 VTAIL.n17 VTAIL.n9 0.155672
R406 VTAIL.n18 VTAIL.n17 0.155672
R407 VTAIL.n18 VTAIL.n5 0.155672
R408 VTAIL.n25 VTAIL.n5 0.155672
R409 VTAIL.n26 VTAIL.n25 0.155672
R410 VTAIL.n26 VTAIL.n1 0.155672
R411 VTAIL.n33 VTAIL.n1 0.155672
R412 VTAIL.n53 VTAIL.n45 0.155672
R413 VTAIL.n54 VTAIL.n53 0.155672
R414 VTAIL.n54 VTAIL.n41 0.155672
R415 VTAIL.n61 VTAIL.n41 0.155672
R416 VTAIL.n62 VTAIL.n61 0.155672
R417 VTAIL.n62 VTAIL.n37 0.155672
R418 VTAIL.n69 VTAIL.n37 0.155672
R419 VTAIL.n89 VTAIL.n81 0.155672
R420 VTAIL.n90 VTAIL.n89 0.155672
R421 VTAIL.n90 VTAIL.n77 0.155672
R422 VTAIL.n97 VTAIL.n77 0.155672
R423 VTAIL.n98 VTAIL.n97 0.155672
R424 VTAIL.n98 VTAIL.n73 0.155672
R425 VTAIL.n105 VTAIL.n73 0.155672
R426 VTAIL.n249 VTAIL.n217 0.155672
R427 VTAIL.n242 VTAIL.n217 0.155672
R428 VTAIL.n242 VTAIL.n241 0.155672
R429 VTAIL.n241 VTAIL.n221 0.155672
R430 VTAIL.n234 VTAIL.n221 0.155672
R431 VTAIL.n234 VTAIL.n233 0.155672
R432 VTAIL.n233 VTAIL.n225 0.155672
R433 VTAIL.n213 VTAIL.n181 0.155672
R434 VTAIL.n206 VTAIL.n181 0.155672
R435 VTAIL.n206 VTAIL.n205 0.155672
R436 VTAIL.n205 VTAIL.n185 0.155672
R437 VTAIL.n198 VTAIL.n185 0.155672
R438 VTAIL.n198 VTAIL.n197 0.155672
R439 VTAIL.n197 VTAIL.n189 0.155672
R440 VTAIL.n177 VTAIL.n145 0.155672
R441 VTAIL.n170 VTAIL.n145 0.155672
R442 VTAIL.n170 VTAIL.n169 0.155672
R443 VTAIL.n169 VTAIL.n149 0.155672
R444 VTAIL.n162 VTAIL.n149 0.155672
R445 VTAIL.n162 VTAIL.n161 0.155672
R446 VTAIL.n161 VTAIL.n153 0.155672
R447 VTAIL.n141 VTAIL.n109 0.155672
R448 VTAIL.n134 VTAIL.n109 0.155672
R449 VTAIL.n134 VTAIL.n133 0.155672
R450 VTAIL.n133 VTAIL.n113 0.155672
R451 VTAIL.n126 VTAIL.n113 0.155672
R452 VTAIL.n126 VTAIL.n125 0.155672
R453 VTAIL.n125 VTAIL.n117 0.155672
R454 VP.n14 VP.n0 161.3
R455 VP.n13 VP.n12 161.3
R456 VP.n11 VP.n1 161.3
R457 VP.n10 VP.n9 161.3
R458 VP.n8 VP.n2 161.3
R459 VP.n7 VP.n6 161.3
R460 VP.n5 VP.n3 103.171
R461 VP.n16 VP.n15 103.171
R462 VP.n4 VP.t0 100.665
R463 VP.n4 VP.t1 99.9113
R464 VP.n3 VP.t2 65.4009
R465 VP.n15 VP.t3 65.4009
R466 VP.n9 VP.n1 56.5193
R467 VP.n5 VP.n4 46.4529
R468 VP.n8 VP.n7 24.4675
R469 VP.n9 VP.n8 24.4675
R470 VP.n13 VP.n1 24.4675
R471 VP.n14 VP.n13 24.4675
R472 VP.n7 VP.n3 7.58527
R473 VP.n15 VP.n14 7.58527
R474 VP.n6 VP.n5 0.278367
R475 VP.n16 VP.n0 0.278367
R476 VP.n6 VP.n2 0.189894
R477 VP.n10 VP.n2 0.189894
R478 VP.n11 VP.n10 0.189894
R479 VP.n12 VP.n11 0.189894
R480 VP.n12 VP.n0 0.189894
R481 VP VP.n16 0.153454
R482 VDD1 VDD1.n1 125.901
R483 VDD1 VDD1.n0 88.6509
R484 VDD1.n0 VDD1.t3 4.83037
R485 VDD1.n0 VDD1.t2 4.83037
R486 VDD1.n1 VDD1.t1 4.83037
R487 VDD1.n1 VDD1.t0 4.83037
R488 B.n383 B.n54 585
R489 B.n385 B.n384 585
R490 B.n386 B.n53 585
R491 B.n388 B.n387 585
R492 B.n389 B.n52 585
R493 B.n391 B.n390 585
R494 B.n392 B.n51 585
R495 B.n394 B.n393 585
R496 B.n395 B.n50 585
R497 B.n397 B.n396 585
R498 B.n398 B.n49 585
R499 B.n400 B.n399 585
R500 B.n401 B.n48 585
R501 B.n403 B.n402 585
R502 B.n404 B.n47 585
R503 B.n406 B.n405 585
R504 B.n407 B.n46 585
R505 B.n409 B.n408 585
R506 B.n410 B.n45 585
R507 B.n412 B.n411 585
R508 B.n413 B.n44 585
R509 B.n415 B.n414 585
R510 B.n416 B.n43 585
R511 B.n418 B.n417 585
R512 B.n419 B.n39 585
R513 B.n421 B.n420 585
R514 B.n422 B.n38 585
R515 B.n424 B.n423 585
R516 B.n425 B.n37 585
R517 B.n427 B.n426 585
R518 B.n428 B.n36 585
R519 B.n430 B.n429 585
R520 B.n431 B.n35 585
R521 B.n433 B.n432 585
R522 B.n434 B.n34 585
R523 B.n436 B.n435 585
R524 B.n438 B.n31 585
R525 B.n440 B.n439 585
R526 B.n441 B.n30 585
R527 B.n443 B.n442 585
R528 B.n444 B.n29 585
R529 B.n446 B.n445 585
R530 B.n447 B.n28 585
R531 B.n449 B.n448 585
R532 B.n450 B.n27 585
R533 B.n452 B.n451 585
R534 B.n453 B.n26 585
R535 B.n455 B.n454 585
R536 B.n456 B.n25 585
R537 B.n458 B.n457 585
R538 B.n459 B.n24 585
R539 B.n461 B.n460 585
R540 B.n462 B.n23 585
R541 B.n464 B.n463 585
R542 B.n465 B.n22 585
R543 B.n467 B.n466 585
R544 B.n468 B.n21 585
R545 B.n470 B.n469 585
R546 B.n471 B.n20 585
R547 B.n473 B.n472 585
R548 B.n474 B.n19 585
R549 B.n476 B.n475 585
R550 B.n382 B.n381 585
R551 B.n380 B.n55 585
R552 B.n379 B.n378 585
R553 B.n377 B.n56 585
R554 B.n376 B.n375 585
R555 B.n374 B.n57 585
R556 B.n373 B.n372 585
R557 B.n371 B.n58 585
R558 B.n370 B.n369 585
R559 B.n368 B.n59 585
R560 B.n367 B.n366 585
R561 B.n365 B.n60 585
R562 B.n364 B.n363 585
R563 B.n362 B.n61 585
R564 B.n361 B.n360 585
R565 B.n359 B.n62 585
R566 B.n358 B.n357 585
R567 B.n356 B.n63 585
R568 B.n355 B.n354 585
R569 B.n353 B.n64 585
R570 B.n352 B.n351 585
R571 B.n350 B.n65 585
R572 B.n349 B.n348 585
R573 B.n347 B.n66 585
R574 B.n346 B.n345 585
R575 B.n344 B.n67 585
R576 B.n343 B.n342 585
R577 B.n341 B.n68 585
R578 B.n340 B.n339 585
R579 B.n338 B.n69 585
R580 B.n337 B.n336 585
R581 B.n335 B.n70 585
R582 B.n334 B.n333 585
R583 B.n332 B.n71 585
R584 B.n331 B.n330 585
R585 B.n329 B.n72 585
R586 B.n328 B.n327 585
R587 B.n326 B.n73 585
R588 B.n325 B.n324 585
R589 B.n323 B.n74 585
R590 B.n322 B.n321 585
R591 B.n320 B.n75 585
R592 B.n319 B.n318 585
R593 B.n317 B.n76 585
R594 B.n316 B.n315 585
R595 B.n314 B.n77 585
R596 B.n313 B.n312 585
R597 B.n311 B.n78 585
R598 B.n310 B.n309 585
R599 B.n308 B.n79 585
R600 B.n307 B.n306 585
R601 B.n305 B.n80 585
R602 B.n304 B.n303 585
R603 B.n302 B.n81 585
R604 B.n301 B.n300 585
R605 B.n299 B.n82 585
R606 B.n298 B.n297 585
R607 B.n296 B.n83 585
R608 B.n295 B.n294 585
R609 B.n293 B.n84 585
R610 B.n292 B.n291 585
R611 B.n290 B.n85 585
R612 B.n289 B.n288 585
R613 B.n287 B.n86 585
R614 B.n286 B.n285 585
R615 B.n284 B.n87 585
R616 B.n283 B.n282 585
R617 B.n188 B.n123 585
R618 B.n190 B.n189 585
R619 B.n191 B.n122 585
R620 B.n193 B.n192 585
R621 B.n194 B.n121 585
R622 B.n196 B.n195 585
R623 B.n197 B.n120 585
R624 B.n199 B.n198 585
R625 B.n200 B.n119 585
R626 B.n202 B.n201 585
R627 B.n203 B.n118 585
R628 B.n205 B.n204 585
R629 B.n206 B.n117 585
R630 B.n208 B.n207 585
R631 B.n209 B.n116 585
R632 B.n211 B.n210 585
R633 B.n212 B.n115 585
R634 B.n214 B.n213 585
R635 B.n215 B.n114 585
R636 B.n217 B.n216 585
R637 B.n218 B.n113 585
R638 B.n220 B.n219 585
R639 B.n221 B.n112 585
R640 B.n223 B.n222 585
R641 B.n224 B.n111 585
R642 B.n226 B.n225 585
R643 B.n228 B.n108 585
R644 B.n230 B.n229 585
R645 B.n231 B.n107 585
R646 B.n233 B.n232 585
R647 B.n234 B.n106 585
R648 B.n236 B.n235 585
R649 B.n237 B.n105 585
R650 B.n239 B.n238 585
R651 B.n240 B.n104 585
R652 B.n242 B.n241 585
R653 B.n244 B.n243 585
R654 B.n245 B.n100 585
R655 B.n247 B.n246 585
R656 B.n248 B.n99 585
R657 B.n250 B.n249 585
R658 B.n251 B.n98 585
R659 B.n253 B.n252 585
R660 B.n254 B.n97 585
R661 B.n256 B.n255 585
R662 B.n257 B.n96 585
R663 B.n259 B.n258 585
R664 B.n260 B.n95 585
R665 B.n262 B.n261 585
R666 B.n263 B.n94 585
R667 B.n265 B.n264 585
R668 B.n266 B.n93 585
R669 B.n268 B.n267 585
R670 B.n269 B.n92 585
R671 B.n271 B.n270 585
R672 B.n272 B.n91 585
R673 B.n274 B.n273 585
R674 B.n275 B.n90 585
R675 B.n277 B.n276 585
R676 B.n278 B.n89 585
R677 B.n280 B.n279 585
R678 B.n281 B.n88 585
R679 B.n187 B.n186 585
R680 B.n185 B.n124 585
R681 B.n184 B.n183 585
R682 B.n182 B.n125 585
R683 B.n181 B.n180 585
R684 B.n179 B.n126 585
R685 B.n178 B.n177 585
R686 B.n176 B.n127 585
R687 B.n175 B.n174 585
R688 B.n173 B.n128 585
R689 B.n172 B.n171 585
R690 B.n170 B.n129 585
R691 B.n169 B.n168 585
R692 B.n167 B.n130 585
R693 B.n166 B.n165 585
R694 B.n164 B.n131 585
R695 B.n163 B.n162 585
R696 B.n161 B.n132 585
R697 B.n160 B.n159 585
R698 B.n158 B.n133 585
R699 B.n157 B.n156 585
R700 B.n155 B.n134 585
R701 B.n154 B.n153 585
R702 B.n152 B.n135 585
R703 B.n151 B.n150 585
R704 B.n149 B.n136 585
R705 B.n148 B.n147 585
R706 B.n146 B.n137 585
R707 B.n145 B.n144 585
R708 B.n143 B.n138 585
R709 B.n142 B.n141 585
R710 B.n140 B.n139 585
R711 B.n2 B.n0 585
R712 B.n525 B.n1 585
R713 B.n524 B.n523 585
R714 B.n522 B.n3 585
R715 B.n521 B.n520 585
R716 B.n519 B.n4 585
R717 B.n518 B.n517 585
R718 B.n516 B.n5 585
R719 B.n515 B.n514 585
R720 B.n513 B.n6 585
R721 B.n512 B.n511 585
R722 B.n510 B.n7 585
R723 B.n509 B.n508 585
R724 B.n507 B.n8 585
R725 B.n506 B.n505 585
R726 B.n504 B.n9 585
R727 B.n503 B.n502 585
R728 B.n501 B.n10 585
R729 B.n500 B.n499 585
R730 B.n498 B.n11 585
R731 B.n497 B.n496 585
R732 B.n495 B.n12 585
R733 B.n494 B.n493 585
R734 B.n492 B.n13 585
R735 B.n491 B.n490 585
R736 B.n489 B.n14 585
R737 B.n488 B.n487 585
R738 B.n486 B.n15 585
R739 B.n485 B.n484 585
R740 B.n483 B.n16 585
R741 B.n482 B.n481 585
R742 B.n480 B.n17 585
R743 B.n479 B.n478 585
R744 B.n477 B.n18 585
R745 B.n527 B.n526 585
R746 B.n188 B.n187 468.476
R747 B.n477 B.n476 468.476
R748 B.n283 B.n88 468.476
R749 B.n381 B.n54 468.476
R750 B.n101 B.t2 335.654
R751 B.n40 B.t10 335.654
R752 B.n109 B.t5 335.654
R753 B.n32 B.t7 335.654
R754 B.n102 B.t1 281.156
R755 B.n41 B.t11 281.156
R756 B.n110 B.t4 281.156
R757 B.n33 B.t8 281.156
R758 B.n101 B.t0 273.259
R759 B.n109 B.t3 273.259
R760 B.n32 B.t6 273.259
R761 B.n40 B.t9 273.259
R762 B.n187 B.n124 163.367
R763 B.n183 B.n124 163.367
R764 B.n183 B.n182 163.367
R765 B.n182 B.n181 163.367
R766 B.n181 B.n126 163.367
R767 B.n177 B.n126 163.367
R768 B.n177 B.n176 163.367
R769 B.n176 B.n175 163.367
R770 B.n175 B.n128 163.367
R771 B.n171 B.n128 163.367
R772 B.n171 B.n170 163.367
R773 B.n170 B.n169 163.367
R774 B.n169 B.n130 163.367
R775 B.n165 B.n130 163.367
R776 B.n165 B.n164 163.367
R777 B.n164 B.n163 163.367
R778 B.n163 B.n132 163.367
R779 B.n159 B.n132 163.367
R780 B.n159 B.n158 163.367
R781 B.n158 B.n157 163.367
R782 B.n157 B.n134 163.367
R783 B.n153 B.n134 163.367
R784 B.n153 B.n152 163.367
R785 B.n152 B.n151 163.367
R786 B.n151 B.n136 163.367
R787 B.n147 B.n136 163.367
R788 B.n147 B.n146 163.367
R789 B.n146 B.n145 163.367
R790 B.n145 B.n138 163.367
R791 B.n141 B.n138 163.367
R792 B.n141 B.n140 163.367
R793 B.n140 B.n2 163.367
R794 B.n526 B.n2 163.367
R795 B.n526 B.n525 163.367
R796 B.n525 B.n524 163.367
R797 B.n524 B.n3 163.367
R798 B.n520 B.n3 163.367
R799 B.n520 B.n519 163.367
R800 B.n519 B.n518 163.367
R801 B.n518 B.n5 163.367
R802 B.n514 B.n5 163.367
R803 B.n514 B.n513 163.367
R804 B.n513 B.n512 163.367
R805 B.n512 B.n7 163.367
R806 B.n508 B.n7 163.367
R807 B.n508 B.n507 163.367
R808 B.n507 B.n506 163.367
R809 B.n506 B.n9 163.367
R810 B.n502 B.n9 163.367
R811 B.n502 B.n501 163.367
R812 B.n501 B.n500 163.367
R813 B.n500 B.n11 163.367
R814 B.n496 B.n11 163.367
R815 B.n496 B.n495 163.367
R816 B.n495 B.n494 163.367
R817 B.n494 B.n13 163.367
R818 B.n490 B.n13 163.367
R819 B.n490 B.n489 163.367
R820 B.n489 B.n488 163.367
R821 B.n488 B.n15 163.367
R822 B.n484 B.n15 163.367
R823 B.n484 B.n483 163.367
R824 B.n483 B.n482 163.367
R825 B.n482 B.n17 163.367
R826 B.n478 B.n17 163.367
R827 B.n478 B.n477 163.367
R828 B.n189 B.n188 163.367
R829 B.n189 B.n122 163.367
R830 B.n193 B.n122 163.367
R831 B.n194 B.n193 163.367
R832 B.n195 B.n194 163.367
R833 B.n195 B.n120 163.367
R834 B.n199 B.n120 163.367
R835 B.n200 B.n199 163.367
R836 B.n201 B.n200 163.367
R837 B.n201 B.n118 163.367
R838 B.n205 B.n118 163.367
R839 B.n206 B.n205 163.367
R840 B.n207 B.n206 163.367
R841 B.n207 B.n116 163.367
R842 B.n211 B.n116 163.367
R843 B.n212 B.n211 163.367
R844 B.n213 B.n212 163.367
R845 B.n213 B.n114 163.367
R846 B.n217 B.n114 163.367
R847 B.n218 B.n217 163.367
R848 B.n219 B.n218 163.367
R849 B.n219 B.n112 163.367
R850 B.n223 B.n112 163.367
R851 B.n224 B.n223 163.367
R852 B.n225 B.n224 163.367
R853 B.n225 B.n108 163.367
R854 B.n230 B.n108 163.367
R855 B.n231 B.n230 163.367
R856 B.n232 B.n231 163.367
R857 B.n232 B.n106 163.367
R858 B.n236 B.n106 163.367
R859 B.n237 B.n236 163.367
R860 B.n238 B.n237 163.367
R861 B.n238 B.n104 163.367
R862 B.n242 B.n104 163.367
R863 B.n243 B.n242 163.367
R864 B.n243 B.n100 163.367
R865 B.n247 B.n100 163.367
R866 B.n248 B.n247 163.367
R867 B.n249 B.n248 163.367
R868 B.n249 B.n98 163.367
R869 B.n253 B.n98 163.367
R870 B.n254 B.n253 163.367
R871 B.n255 B.n254 163.367
R872 B.n255 B.n96 163.367
R873 B.n259 B.n96 163.367
R874 B.n260 B.n259 163.367
R875 B.n261 B.n260 163.367
R876 B.n261 B.n94 163.367
R877 B.n265 B.n94 163.367
R878 B.n266 B.n265 163.367
R879 B.n267 B.n266 163.367
R880 B.n267 B.n92 163.367
R881 B.n271 B.n92 163.367
R882 B.n272 B.n271 163.367
R883 B.n273 B.n272 163.367
R884 B.n273 B.n90 163.367
R885 B.n277 B.n90 163.367
R886 B.n278 B.n277 163.367
R887 B.n279 B.n278 163.367
R888 B.n279 B.n88 163.367
R889 B.n284 B.n283 163.367
R890 B.n285 B.n284 163.367
R891 B.n285 B.n86 163.367
R892 B.n289 B.n86 163.367
R893 B.n290 B.n289 163.367
R894 B.n291 B.n290 163.367
R895 B.n291 B.n84 163.367
R896 B.n295 B.n84 163.367
R897 B.n296 B.n295 163.367
R898 B.n297 B.n296 163.367
R899 B.n297 B.n82 163.367
R900 B.n301 B.n82 163.367
R901 B.n302 B.n301 163.367
R902 B.n303 B.n302 163.367
R903 B.n303 B.n80 163.367
R904 B.n307 B.n80 163.367
R905 B.n308 B.n307 163.367
R906 B.n309 B.n308 163.367
R907 B.n309 B.n78 163.367
R908 B.n313 B.n78 163.367
R909 B.n314 B.n313 163.367
R910 B.n315 B.n314 163.367
R911 B.n315 B.n76 163.367
R912 B.n319 B.n76 163.367
R913 B.n320 B.n319 163.367
R914 B.n321 B.n320 163.367
R915 B.n321 B.n74 163.367
R916 B.n325 B.n74 163.367
R917 B.n326 B.n325 163.367
R918 B.n327 B.n326 163.367
R919 B.n327 B.n72 163.367
R920 B.n331 B.n72 163.367
R921 B.n332 B.n331 163.367
R922 B.n333 B.n332 163.367
R923 B.n333 B.n70 163.367
R924 B.n337 B.n70 163.367
R925 B.n338 B.n337 163.367
R926 B.n339 B.n338 163.367
R927 B.n339 B.n68 163.367
R928 B.n343 B.n68 163.367
R929 B.n344 B.n343 163.367
R930 B.n345 B.n344 163.367
R931 B.n345 B.n66 163.367
R932 B.n349 B.n66 163.367
R933 B.n350 B.n349 163.367
R934 B.n351 B.n350 163.367
R935 B.n351 B.n64 163.367
R936 B.n355 B.n64 163.367
R937 B.n356 B.n355 163.367
R938 B.n357 B.n356 163.367
R939 B.n357 B.n62 163.367
R940 B.n361 B.n62 163.367
R941 B.n362 B.n361 163.367
R942 B.n363 B.n362 163.367
R943 B.n363 B.n60 163.367
R944 B.n367 B.n60 163.367
R945 B.n368 B.n367 163.367
R946 B.n369 B.n368 163.367
R947 B.n369 B.n58 163.367
R948 B.n373 B.n58 163.367
R949 B.n374 B.n373 163.367
R950 B.n375 B.n374 163.367
R951 B.n375 B.n56 163.367
R952 B.n379 B.n56 163.367
R953 B.n380 B.n379 163.367
R954 B.n381 B.n380 163.367
R955 B.n476 B.n19 163.367
R956 B.n472 B.n19 163.367
R957 B.n472 B.n471 163.367
R958 B.n471 B.n470 163.367
R959 B.n470 B.n21 163.367
R960 B.n466 B.n21 163.367
R961 B.n466 B.n465 163.367
R962 B.n465 B.n464 163.367
R963 B.n464 B.n23 163.367
R964 B.n460 B.n23 163.367
R965 B.n460 B.n459 163.367
R966 B.n459 B.n458 163.367
R967 B.n458 B.n25 163.367
R968 B.n454 B.n25 163.367
R969 B.n454 B.n453 163.367
R970 B.n453 B.n452 163.367
R971 B.n452 B.n27 163.367
R972 B.n448 B.n27 163.367
R973 B.n448 B.n447 163.367
R974 B.n447 B.n446 163.367
R975 B.n446 B.n29 163.367
R976 B.n442 B.n29 163.367
R977 B.n442 B.n441 163.367
R978 B.n441 B.n440 163.367
R979 B.n440 B.n31 163.367
R980 B.n435 B.n31 163.367
R981 B.n435 B.n434 163.367
R982 B.n434 B.n433 163.367
R983 B.n433 B.n35 163.367
R984 B.n429 B.n35 163.367
R985 B.n429 B.n428 163.367
R986 B.n428 B.n427 163.367
R987 B.n427 B.n37 163.367
R988 B.n423 B.n37 163.367
R989 B.n423 B.n422 163.367
R990 B.n422 B.n421 163.367
R991 B.n421 B.n39 163.367
R992 B.n417 B.n39 163.367
R993 B.n417 B.n416 163.367
R994 B.n416 B.n415 163.367
R995 B.n415 B.n44 163.367
R996 B.n411 B.n44 163.367
R997 B.n411 B.n410 163.367
R998 B.n410 B.n409 163.367
R999 B.n409 B.n46 163.367
R1000 B.n405 B.n46 163.367
R1001 B.n405 B.n404 163.367
R1002 B.n404 B.n403 163.367
R1003 B.n403 B.n48 163.367
R1004 B.n399 B.n48 163.367
R1005 B.n399 B.n398 163.367
R1006 B.n398 B.n397 163.367
R1007 B.n397 B.n50 163.367
R1008 B.n393 B.n50 163.367
R1009 B.n393 B.n392 163.367
R1010 B.n392 B.n391 163.367
R1011 B.n391 B.n52 163.367
R1012 B.n387 B.n52 163.367
R1013 B.n387 B.n386 163.367
R1014 B.n386 B.n385 163.367
R1015 B.n385 B.n54 163.367
R1016 B.n103 B.n102 59.5399
R1017 B.n227 B.n110 59.5399
R1018 B.n437 B.n33 59.5399
R1019 B.n42 B.n41 59.5399
R1020 B.n102 B.n101 54.4975
R1021 B.n110 B.n109 54.4975
R1022 B.n33 B.n32 54.4975
R1023 B.n41 B.n40 54.4975
R1024 B.n475 B.n18 30.4395
R1025 B.n383 B.n382 30.4395
R1026 B.n282 B.n281 30.4395
R1027 B.n186 B.n123 30.4395
R1028 B B.n527 18.0485
R1029 B.n475 B.n474 10.6151
R1030 B.n474 B.n473 10.6151
R1031 B.n473 B.n20 10.6151
R1032 B.n469 B.n20 10.6151
R1033 B.n469 B.n468 10.6151
R1034 B.n468 B.n467 10.6151
R1035 B.n467 B.n22 10.6151
R1036 B.n463 B.n22 10.6151
R1037 B.n463 B.n462 10.6151
R1038 B.n462 B.n461 10.6151
R1039 B.n461 B.n24 10.6151
R1040 B.n457 B.n24 10.6151
R1041 B.n457 B.n456 10.6151
R1042 B.n456 B.n455 10.6151
R1043 B.n455 B.n26 10.6151
R1044 B.n451 B.n26 10.6151
R1045 B.n451 B.n450 10.6151
R1046 B.n450 B.n449 10.6151
R1047 B.n449 B.n28 10.6151
R1048 B.n445 B.n28 10.6151
R1049 B.n445 B.n444 10.6151
R1050 B.n444 B.n443 10.6151
R1051 B.n443 B.n30 10.6151
R1052 B.n439 B.n30 10.6151
R1053 B.n439 B.n438 10.6151
R1054 B.n436 B.n34 10.6151
R1055 B.n432 B.n34 10.6151
R1056 B.n432 B.n431 10.6151
R1057 B.n431 B.n430 10.6151
R1058 B.n430 B.n36 10.6151
R1059 B.n426 B.n36 10.6151
R1060 B.n426 B.n425 10.6151
R1061 B.n425 B.n424 10.6151
R1062 B.n424 B.n38 10.6151
R1063 B.n420 B.n419 10.6151
R1064 B.n419 B.n418 10.6151
R1065 B.n418 B.n43 10.6151
R1066 B.n414 B.n43 10.6151
R1067 B.n414 B.n413 10.6151
R1068 B.n413 B.n412 10.6151
R1069 B.n412 B.n45 10.6151
R1070 B.n408 B.n45 10.6151
R1071 B.n408 B.n407 10.6151
R1072 B.n407 B.n406 10.6151
R1073 B.n406 B.n47 10.6151
R1074 B.n402 B.n47 10.6151
R1075 B.n402 B.n401 10.6151
R1076 B.n401 B.n400 10.6151
R1077 B.n400 B.n49 10.6151
R1078 B.n396 B.n49 10.6151
R1079 B.n396 B.n395 10.6151
R1080 B.n395 B.n394 10.6151
R1081 B.n394 B.n51 10.6151
R1082 B.n390 B.n51 10.6151
R1083 B.n390 B.n389 10.6151
R1084 B.n389 B.n388 10.6151
R1085 B.n388 B.n53 10.6151
R1086 B.n384 B.n53 10.6151
R1087 B.n384 B.n383 10.6151
R1088 B.n282 B.n87 10.6151
R1089 B.n286 B.n87 10.6151
R1090 B.n287 B.n286 10.6151
R1091 B.n288 B.n287 10.6151
R1092 B.n288 B.n85 10.6151
R1093 B.n292 B.n85 10.6151
R1094 B.n293 B.n292 10.6151
R1095 B.n294 B.n293 10.6151
R1096 B.n294 B.n83 10.6151
R1097 B.n298 B.n83 10.6151
R1098 B.n299 B.n298 10.6151
R1099 B.n300 B.n299 10.6151
R1100 B.n300 B.n81 10.6151
R1101 B.n304 B.n81 10.6151
R1102 B.n305 B.n304 10.6151
R1103 B.n306 B.n305 10.6151
R1104 B.n306 B.n79 10.6151
R1105 B.n310 B.n79 10.6151
R1106 B.n311 B.n310 10.6151
R1107 B.n312 B.n311 10.6151
R1108 B.n312 B.n77 10.6151
R1109 B.n316 B.n77 10.6151
R1110 B.n317 B.n316 10.6151
R1111 B.n318 B.n317 10.6151
R1112 B.n318 B.n75 10.6151
R1113 B.n322 B.n75 10.6151
R1114 B.n323 B.n322 10.6151
R1115 B.n324 B.n323 10.6151
R1116 B.n324 B.n73 10.6151
R1117 B.n328 B.n73 10.6151
R1118 B.n329 B.n328 10.6151
R1119 B.n330 B.n329 10.6151
R1120 B.n330 B.n71 10.6151
R1121 B.n334 B.n71 10.6151
R1122 B.n335 B.n334 10.6151
R1123 B.n336 B.n335 10.6151
R1124 B.n336 B.n69 10.6151
R1125 B.n340 B.n69 10.6151
R1126 B.n341 B.n340 10.6151
R1127 B.n342 B.n341 10.6151
R1128 B.n342 B.n67 10.6151
R1129 B.n346 B.n67 10.6151
R1130 B.n347 B.n346 10.6151
R1131 B.n348 B.n347 10.6151
R1132 B.n348 B.n65 10.6151
R1133 B.n352 B.n65 10.6151
R1134 B.n353 B.n352 10.6151
R1135 B.n354 B.n353 10.6151
R1136 B.n354 B.n63 10.6151
R1137 B.n358 B.n63 10.6151
R1138 B.n359 B.n358 10.6151
R1139 B.n360 B.n359 10.6151
R1140 B.n360 B.n61 10.6151
R1141 B.n364 B.n61 10.6151
R1142 B.n365 B.n364 10.6151
R1143 B.n366 B.n365 10.6151
R1144 B.n366 B.n59 10.6151
R1145 B.n370 B.n59 10.6151
R1146 B.n371 B.n370 10.6151
R1147 B.n372 B.n371 10.6151
R1148 B.n372 B.n57 10.6151
R1149 B.n376 B.n57 10.6151
R1150 B.n377 B.n376 10.6151
R1151 B.n378 B.n377 10.6151
R1152 B.n378 B.n55 10.6151
R1153 B.n382 B.n55 10.6151
R1154 B.n190 B.n123 10.6151
R1155 B.n191 B.n190 10.6151
R1156 B.n192 B.n191 10.6151
R1157 B.n192 B.n121 10.6151
R1158 B.n196 B.n121 10.6151
R1159 B.n197 B.n196 10.6151
R1160 B.n198 B.n197 10.6151
R1161 B.n198 B.n119 10.6151
R1162 B.n202 B.n119 10.6151
R1163 B.n203 B.n202 10.6151
R1164 B.n204 B.n203 10.6151
R1165 B.n204 B.n117 10.6151
R1166 B.n208 B.n117 10.6151
R1167 B.n209 B.n208 10.6151
R1168 B.n210 B.n209 10.6151
R1169 B.n210 B.n115 10.6151
R1170 B.n214 B.n115 10.6151
R1171 B.n215 B.n214 10.6151
R1172 B.n216 B.n215 10.6151
R1173 B.n216 B.n113 10.6151
R1174 B.n220 B.n113 10.6151
R1175 B.n221 B.n220 10.6151
R1176 B.n222 B.n221 10.6151
R1177 B.n222 B.n111 10.6151
R1178 B.n226 B.n111 10.6151
R1179 B.n229 B.n228 10.6151
R1180 B.n229 B.n107 10.6151
R1181 B.n233 B.n107 10.6151
R1182 B.n234 B.n233 10.6151
R1183 B.n235 B.n234 10.6151
R1184 B.n235 B.n105 10.6151
R1185 B.n239 B.n105 10.6151
R1186 B.n240 B.n239 10.6151
R1187 B.n241 B.n240 10.6151
R1188 B.n245 B.n244 10.6151
R1189 B.n246 B.n245 10.6151
R1190 B.n246 B.n99 10.6151
R1191 B.n250 B.n99 10.6151
R1192 B.n251 B.n250 10.6151
R1193 B.n252 B.n251 10.6151
R1194 B.n252 B.n97 10.6151
R1195 B.n256 B.n97 10.6151
R1196 B.n257 B.n256 10.6151
R1197 B.n258 B.n257 10.6151
R1198 B.n258 B.n95 10.6151
R1199 B.n262 B.n95 10.6151
R1200 B.n263 B.n262 10.6151
R1201 B.n264 B.n263 10.6151
R1202 B.n264 B.n93 10.6151
R1203 B.n268 B.n93 10.6151
R1204 B.n269 B.n268 10.6151
R1205 B.n270 B.n269 10.6151
R1206 B.n270 B.n91 10.6151
R1207 B.n274 B.n91 10.6151
R1208 B.n275 B.n274 10.6151
R1209 B.n276 B.n275 10.6151
R1210 B.n276 B.n89 10.6151
R1211 B.n280 B.n89 10.6151
R1212 B.n281 B.n280 10.6151
R1213 B.n186 B.n185 10.6151
R1214 B.n185 B.n184 10.6151
R1215 B.n184 B.n125 10.6151
R1216 B.n180 B.n125 10.6151
R1217 B.n180 B.n179 10.6151
R1218 B.n179 B.n178 10.6151
R1219 B.n178 B.n127 10.6151
R1220 B.n174 B.n127 10.6151
R1221 B.n174 B.n173 10.6151
R1222 B.n173 B.n172 10.6151
R1223 B.n172 B.n129 10.6151
R1224 B.n168 B.n129 10.6151
R1225 B.n168 B.n167 10.6151
R1226 B.n167 B.n166 10.6151
R1227 B.n166 B.n131 10.6151
R1228 B.n162 B.n131 10.6151
R1229 B.n162 B.n161 10.6151
R1230 B.n161 B.n160 10.6151
R1231 B.n160 B.n133 10.6151
R1232 B.n156 B.n133 10.6151
R1233 B.n156 B.n155 10.6151
R1234 B.n155 B.n154 10.6151
R1235 B.n154 B.n135 10.6151
R1236 B.n150 B.n135 10.6151
R1237 B.n150 B.n149 10.6151
R1238 B.n149 B.n148 10.6151
R1239 B.n148 B.n137 10.6151
R1240 B.n144 B.n137 10.6151
R1241 B.n144 B.n143 10.6151
R1242 B.n143 B.n142 10.6151
R1243 B.n142 B.n139 10.6151
R1244 B.n139 B.n0 10.6151
R1245 B.n523 B.n1 10.6151
R1246 B.n523 B.n522 10.6151
R1247 B.n522 B.n521 10.6151
R1248 B.n521 B.n4 10.6151
R1249 B.n517 B.n4 10.6151
R1250 B.n517 B.n516 10.6151
R1251 B.n516 B.n515 10.6151
R1252 B.n515 B.n6 10.6151
R1253 B.n511 B.n6 10.6151
R1254 B.n511 B.n510 10.6151
R1255 B.n510 B.n509 10.6151
R1256 B.n509 B.n8 10.6151
R1257 B.n505 B.n8 10.6151
R1258 B.n505 B.n504 10.6151
R1259 B.n504 B.n503 10.6151
R1260 B.n503 B.n10 10.6151
R1261 B.n499 B.n10 10.6151
R1262 B.n499 B.n498 10.6151
R1263 B.n498 B.n497 10.6151
R1264 B.n497 B.n12 10.6151
R1265 B.n493 B.n12 10.6151
R1266 B.n493 B.n492 10.6151
R1267 B.n492 B.n491 10.6151
R1268 B.n491 B.n14 10.6151
R1269 B.n487 B.n14 10.6151
R1270 B.n487 B.n486 10.6151
R1271 B.n486 B.n485 10.6151
R1272 B.n485 B.n16 10.6151
R1273 B.n481 B.n16 10.6151
R1274 B.n481 B.n480 10.6151
R1275 B.n480 B.n479 10.6151
R1276 B.n479 B.n18 10.6151
R1277 B.n438 B.n437 9.36635
R1278 B.n420 B.n42 9.36635
R1279 B.n227 B.n226 9.36635
R1280 B.n244 B.n103 9.36635
R1281 B.n527 B.n0 2.81026
R1282 B.n527 B.n1 2.81026
R1283 B.n437 B.n436 1.24928
R1284 B.n42 B.n38 1.24928
R1285 B.n228 B.n227 1.24928
R1286 B.n241 B.n103 1.24928
C0 VN B 1.02242f
C1 VDD2 w_n2656_n2314# 1.34503f
C2 VDD1 VP 3.0157f
C3 VP VTAIL 3.02433f
C4 VDD1 VTAIL 4.11398f
C5 VDD2 B 1.14779f
C6 VP VN 5.13077f
C7 VDD1 VN 0.149025f
C8 VTAIL VN 3.01023f
C9 w_n2656_n2314# B 7.62602f
C10 VDD2 VP 0.386803f
C11 VDD1 VDD2 1.00451f
C12 VDD2 VTAIL 4.16738f
C13 VP w_n2656_n2314# 4.72292f
C14 VDD1 w_n2656_n2314# 1.29154f
C15 w_n2656_n2314# VTAIL 2.7828f
C16 VDD2 VN 2.77863f
C17 VP B 1.58796f
C18 w_n2656_n2314# VN 4.38178f
C19 VDD1 B 1.09765f
C20 VTAIL B 3.17092f
C21 VDD2 VSUBS 0.79196f
C22 VDD1 VSUBS 4.961635f
C23 VTAIL VSUBS 0.721164f
C24 VN VSUBS 5.21798f
C25 VP VSUBS 1.905687f
C26 B VSUBS 3.729722f
C27 w_n2656_n2314# VSUBS 76.524704f
C28 B.n0 VSUBS 0.005077f
C29 B.n1 VSUBS 0.005077f
C30 B.n2 VSUBS 0.008029f
C31 B.n3 VSUBS 0.008029f
C32 B.n4 VSUBS 0.008029f
C33 B.n5 VSUBS 0.008029f
C34 B.n6 VSUBS 0.008029f
C35 B.n7 VSUBS 0.008029f
C36 B.n8 VSUBS 0.008029f
C37 B.n9 VSUBS 0.008029f
C38 B.n10 VSUBS 0.008029f
C39 B.n11 VSUBS 0.008029f
C40 B.n12 VSUBS 0.008029f
C41 B.n13 VSUBS 0.008029f
C42 B.n14 VSUBS 0.008029f
C43 B.n15 VSUBS 0.008029f
C44 B.n16 VSUBS 0.008029f
C45 B.n17 VSUBS 0.008029f
C46 B.n18 VSUBS 0.017463f
C47 B.n19 VSUBS 0.008029f
C48 B.n20 VSUBS 0.008029f
C49 B.n21 VSUBS 0.008029f
C50 B.n22 VSUBS 0.008029f
C51 B.n23 VSUBS 0.008029f
C52 B.n24 VSUBS 0.008029f
C53 B.n25 VSUBS 0.008029f
C54 B.n26 VSUBS 0.008029f
C55 B.n27 VSUBS 0.008029f
C56 B.n28 VSUBS 0.008029f
C57 B.n29 VSUBS 0.008029f
C58 B.n30 VSUBS 0.008029f
C59 B.n31 VSUBS 0.008029f
C60 B.t8 VSUBS 0.117743f
C61 B.t7 VSUBS 0.147389f
C62 B.t6 VSUBS 0.898235f
C63 B.n32 VSUBS 0.248995f
C64 B.n33 VSUBS 0.194039f
C65 B.n34 VSUBS 0.008029f
C66 B.n35 VSUBS 0.008029f
C67 B.n36 VSUBS 0.008029f
C68 B.n37 VSUBS 0.008029f
C69 B.n38 VSUBS 0.004487f
C70 B.n39 VSUBS 0.008029f
C71 B.t11 VSUBS 0.117746f
C72 B.t10 VSUBS 0.14739f
C73 B.t9 VSUBS 0.898235f
C74 B.n40 VSUBS 0.248993f
C75 B.n41 VSUBS 0.194037f
C76 B.n42 VSUBS 0.018602f
C77 B.n43 VSUBS 0.008029f
C78 B.n44 VSUBS 0.008029f
C79 B.n45 VSUBS 0.008029f
C80 B.n46 VSUBS 0.008029f
C81 B.n47 VSUBS 0.008029f
C82 B.n48 VSUBS 0.008029f
C83 B.n49 VSUBS 0.008029f
C84 B.n50 VSUBS 0.008029f
C85 B.n51 VSUBS 0.008029f
C86 B.n52 VSUBS 0.008029f
C87 B.n53 VSUBS 0.008029f
C88 B.n54 VSUBS 0.018431f
C89 B.n55 VSUBS 0.008029f
C90 B.n56 VSUBS 0.008029f
C91 B.n57 VSUBS 0.008029f
C92 B.n58 VSUBS 0.008029f
C93 B.n59 VSUBS 0.008029f
C94 B.n60 VSUBS 0.008029f
C95 B.n61 VSUBS 0.008029f
C96 B.n62 VSUBS 0.008029f
C97 B.n63 VSUBS 0.008029f
C98 B.n64 VSUBS 0.008029f
C99 B.n65 VSUBS 0.008029f
C100 B.n66 VSUBS 0.008029f
C101 B.n67 VSUBS 0.008029f
C102 B.n68 VSUBS 0.008029f
C103 B.n69 VSUBS 0.008029f
C104 B.n70 VSUBS 0.008029f
C105 B.n71 VSUBS 0.008029f
C106 B.n72 VSUBS 0.008029f
C107 B.n73 VSUBS 0.008029f
C108 B.n74 VSUBS 0.008029f
C109 B.n75 VSUBS 0.008029f
C110 B.n76 VSUBS 0.008029f
C111 B.n77 VSUBS 0.008029f
C112 B.n78 VSUBS 0.008029f
C113 B.n79 VSUBS 0.008029f
C114 B.n80 VSUBS 0.008029f
C115 B.n81 VSUBS 0.008029f
C116 B.n82 VSUBS 0.008029f
C117 B.n83 VSUBS 0.008029f
C118 B.n84 VSUBS 0.008029f
C119 B.n85 VSUBS 0.008029f
C120 B.n86 VSUBS 0.008029f
C121 B.n87 VSUBS 0.008029f
C122 B.n88 VSUBS 0.018431f
C123 B.n89 VSUBS 0.008029f
C124 B.n90 VSUBS 0.008029f
C125 B.n91 VSUBS 0.008029f
C126 B.n92 VSUBS 0.008029f
C127 B.n93 VSUBS 0.008029f
C128 B.n94 VSUBS 0.008029f
C129 B.n95 VSUBS 0.008029f
C130 B.n96 VSUBS 0.008029f
C131 B.n97 VSUBS 0.008029f
C132 B.n98 VSUBS 0.008029f
C133 B.n99 VSUBS 0.008029f
C134 B.n100 VSUBS 0.008029f
C135 B.t1 VSUBS 0.117746f
C136 B.t2 VSUBS 0.14739f
C137 B.t0 VSUBS 0.898235f
C138 B.n101 VSUBS 0.248993f
C139 B.n102 VSUBS 0.194037f
C140 B.n103 VSUBS 0.018602f
C141 B.n104 VSUBS 0.008029f
C142 B.n105 VSUBS 0.008029f
C143 B.n106 VSUBS 0.008029f
C144 B.n107 VSUBS 0.008029f
C145 B.n108 VSUBS 0.008029f
C146 B.t4 VSUBS 0.117743f
C147 B.t5 VSUBS 0.147389f
C148 B.t3 VSUBS 0.898235f
C149 B.n109 VSUBS 0.248995f
C150 B.n110 VSUBS 0.194039f
C151 B.n111 VSUBS 0.008029f
C152 B.n112 VSUBS 0.008029f
C153 B.n113 VSUBS 0.008029f
C154 B.n114 VSUBS 0.008029f
C155 B.n115 VSUBS 0.008029f
C156 B.n116 VSUBS 0.008029f
C157 B.n117 VSUBS 0.008029f
C158 B.n118 VSUBS 0.008029f
C159 B.n119 VSUBS 0.008029f
C160 B.n120 VSUBS 0.008029f
C161 B.n121 VSUBS 0.008029f
C162 B.n122 VSUBS 0.008029f
C163 B.n123 VSUBS 0.018431f
C164 B.n124 VSUBS 0.008029f
C165 B.n125 VSUBS 0.008029f
C166 B.n126 VSUBS 0.008029f
C167 B.n127 VSUBS 0.008029f
C168 B.n128 VSUBS 0.008029f
C169 B.n129 VSUBS 0.008029f
C170 B.n130 VSUBS 0.008029f
C171 B.n131 VSUBS 0.008029f
C172 B.n132 VSUBS 0.008029f
C173 B.n133 VSUBS 0.008029f
C174 B.n134 VSUBS 0.008029f
C175 B.n135 VSUBS 0.008029f
C176 B.n136 VSUBS 0.008029f
C177 B.n137 VSUBS 0.008029f
C178 B.n138 VSUBS 0.008029f
C179 B.n139 VSUBS 0.008029f
C180 B.n140 VSUBS 0.008029f
C181 B.n141 VSUBS 0.008029f
C182 B.n142 VSUBS 0.008029f
C183 B.n143 VSUBS 0.008029f
C184 B.n144 VSUBS 0.008029f
C185 B.n145 VSUBS 0.008029f
C186 B.n146 VSUBS 0.008029f
C187 B.n147 VSUBS 0.008029f
C188 B.n148 VSUBS 0.008029f
C189 B.n149 VSUBS 0.008029f
C190 B.n150 VSUBS 0.008029f
C191 B.n151 VSUBS 0.008029f
C192 B.n152 VSUBS 0.008029f
C193 B.n153 VSUBS 0.008029f
C194 B.n154 VSUBS 0.008029f
C195 B.n155 VSUBS 0.008029f
C196 B.n156 VSUBS 0.008029f
C197 B.n157 VSUBS 0.008029f
C198 B.n158 VSUBS 0.008029f
C199 B.n159 VSUBS 0.008029f
C200 B.n160 VSUBS 0.008029f
C201 B.n161 VSUBS 0.008029f
C202 B.n162 VSUBS 0.008029f
C203 B.n163 VSUBS 0.008029f
C204 B.n164 VSUBS 0.008029f
C205 B.n165 VSUBS 0.008029f
C206 B.n166 VSUBS 0.008029f
C207 B.n167 VSUBS 0.008029f
C208 B.n168 VSUBS 0.008029f
C209 B.n169 VSUBS 0.008029f
C210 B.n170 VSUBS 0.008029f
C211 B.n171 VSUBS 0.008029f
C212 B.n172 VSUBS 0.008029f
C213 B.n173 VSUBS 0.008029f
C214 B.n174 VSUBS 0.008029f
C215 B.n175 VSUBS 0.008029f
C216 B.n176 VSUBS 0.008029f
C217 B.n177 VSUBS 0.008029f
C218 B.n178 VSUBS 0.008029f
C219 B.n179 VSUBS 0.008029f
C220 B.n180 VSUBS 0.008029f
C221 B.n181 VSUBS 0.008029f
C222 B.n182 VSUBS 0.008029f
C223 B.n183 VSUBS 0.008029f
C224 B.n184 VSUBS 0.008029f
C225 B.n185 VSUBS 0.008029f
C226 B.n186 VSUBS 0.017463f
C227 B.n187 VSUBS 0.017463f
C228 B.n188 VSUBS 0.018431f
C229 B.n189 VSUBS 0.008029f
C230 B.n190 VSUBS 0.008029f
C231 B.n191 VSUBS 0.008029f
C232 B.n192 VSUBS 0.008029f
C233 B.n193 VSUBS 0.008029f
C234 B.n194 VSUBS 0.008029f
C235 B.n195 VSUBS 0.008029f
C236 B.n196 VSUBS 0.008029f
C237 B.n197 VSUBS 0.008029f
C238 B.n198 VSUBS 0.008029f
C239 B.n199 VSUBS 0.008029f
C240 B.n200 VSUBS 0.008029f
C241 B.n201 VSUBS 0.008029f
C242 B.n202 VSUBS 0.008029f
C243 B.n203 VSUBS 0.008029f
C244 B.n204 VSUBS 0.008029f
C245 B.n205 VSUBS 0.008029f
C246 B.n206 VSUBS 0.008029f
C247 B.n207 VSUBS 0.008029f
C248 B.n208 VSUBS 0.008029f
C249 B.n209 VSUBS 0.008029f
C250 B.n210 VSUBS 0.008029f
C251 B.n211 VSUBS 0.008029f
C252 B.n212 VSUBS 0.008029f
C253 B.n213 VSUBS 0.008029f
C254 B.n214 VSUBS 0.008029f
C255 B.n215 VSUBS 0.008029f
C256 B.n216 VSUBS 0.008029f
C257 B.n217 VSUBS 0.008029f
C258 B.n218 VSUBS 0.008029f
C259 B.n219 VSUBS 0.008029f
C260 B.n220 VSUBS 0.008029f
C261 B.n221 VSUBS 0.008029f
C262 B.n222 VSUBS 0.008029f
C263 B.n223 VSUBS 0.008029f
C264 B.n224 VSUBS 0.008029f
C265 B.n225 VSUBS 0.008029f
C266 B.n226 VSUBS 0.007557f
C267 B.n227 VSUBS 0.018602f
C268 B.n228 VSUBS 0.004487f
C269 B.n229 VSUBS 0.008029f
C270 B.n230 VSUBS 0.008029f
C271 B.n231 VSUBS 0.008029f
C272 B.n232 VSUBS 0.008029f
C273 B.n233 VSUBS 0.008029f
C274 B.n234 VSUBS 0.008029f
C275 B.n235 VSUBS 0.008029f
C276 B.n236 VSUBS 0.008029f
C277 B.n237 VSUBS 0.008029f
C278 B.n238 VSUBS 0.008029f
C279 B.n239 VSUBS 0.008029f
C280 B.n240 VSUBS 0.008029f
C281 B.n241 VSUBS 0.004487f
C282 B.n242 VSUBS 0.008029f
C283 B.n243 VSUBS 0.008029f
C284 B.n244 VSUBS 0.007557f
C285 B.n245 VSUBS 0.008029f
C286 B.n246 VSUBS 0.008029f
C287 B.n247 VSUBS 0.008029f
C288 B.n248 VSUBS 0.008029f
C289 B.n249 VSUBS 0.008029f
C290 B.n250 VSUBS 0.008029f
C291 B.n251 VSUBS 0.008029f
C292 B.n252 VSUBS 0.008029f
C293 B.n253 VSUBS 0.008029f
C294 B.n254 VSUBS 0.008029f
C295 B.n255 VSUBS 0.008029f
C296 B.n256 VSUBS 0.008029f
C297 B.n257 VSUBS 0.008029f
C298 B.n258 VSUBS 0.008029f
C299 B.n259 VSUBS 0.008029f
C300 B.n260 VSUBS 0.008029f
C301 B.n261 VSUBS 0.008029f
C302 B.n262 VSUBS 0.008029f
C303 B.n263 VSUBS 0.008029f
C304 B.n264 VSUBS 0.008029f
C305 B.n265 VSUBS 0.008029f
C306 B.n266 VSUBS 0.008029f
C307 B.n267 VSUBS 0.008029f
C308 B.n268 VSUBS 0.008029f
C309 B.n269 VSUBS 0.008029f
C310 B.n270 VSUBS 0.008029f
C311 B.n271 VSUBS 0.008029f
C312 B.n272 VSUBS 0.008029f
C313 B.n273 VSUBS 0.008029f
C314 B.n274 VSUBS 0.008029f
C315 B.n275 VSUBS 0.008029f
C316 B.n276 VSUBS 0.008029f
C317 B.n277 VSUBS 0.008029f
C318 B.n278 VSUBS 0.008029f
C319 B.n279 VSUBS 0.008029f
C320 B.n280 VSUBS 0.008029f
C321 B.n281 VSUBS 0.018431f
C322 B.n282 VSUBS 0.017463f
C323 B.n283 VSUBS 0.017463f
C324 B.n284 VSUBS 0.008029f
C325 B.n285 VSUBS 0.008029f
C326 B.n286 VSUBS 0.008029f
C327 B.n287 VSUBS 0.008029f
C328 B.n288 VSUBS 0.008029f
C329 B.n289 VSUBS 0.008029f
C330 B.n290 VSUBS 0.008029f
C331 B.n291 VSUBS 0.008029f
C332 B.n292 VSUBS 0.008029f
C333 B.n293 VSUBS 0.008029f
C334 B.n294 VSUBS 0.008029f
C335 B.n295 VSUBS 0.008029f
C336 B.n296 VSUBS 0.008029f
C337 B.n297 VSUBS 0.008029f
C338 B.n298 VSUBS 0.008029f
C339 B.n299 VSUBS 0.008029f
C340 B.n300 VSUBS 0.008029f
C341 B.n301 VSUBS 0.008029f
C342 B.n302 VSUBS 0.008029f
C343 B.n303 VSUBS 0.008029f
C344 B.n304 VSUBS 0.008029f
C345 B.n305 VSUBS 0.008029f
C346 B.n306 VSUBS 0.008029f
C347 B.n307 VSUBS 0.008029f
C348 B.n308 VSUBS 0.008029f
C349 B.n309 VSUBS 0.008029f
C350 B.n310 VSUBS 0.008029f
C351 B.n311 VSUBS 0.008029f
C352 B.n312 VSUBS 0.008029f
C353 B.n313 VSUBS 0.008029f
C354 B.n314 VSUBS 0.008029f
C355 B.n315 VSUBS 0.008029f
C356 B.n316 VSUBS 0.008029f
C357 B.n317 VSUBS 0.008029f
C358 B.n318 VSUBS 0.008029f
C359 B.n319 VSUBS 0.008029f
C360 B.n320 VSUBS 0.008029f
C361 B.n321 VSUBS 0.008029f
C362 B.n322 VSUBS 0.008029f
C363 B.n323 VSUBS 0.008029f
C364 B.n324 VSUBS 0.008029f
C365 B.n325 VSUBS 0.008029f
C366 B.n326 VSUBS 0.008029f
C367 B.n327 VSUBS 0.008029f
C368 B.n328 VSUBS 0.008029f
C369 B.n329 VSUBS 0.008029f
C370 B.n330 VSUBS 0.008029f
C371 B.n331 VSUBS 0.008029f
C372 B.n332 VSUBS 0.008029f
C373 B.n333 VSUBS 0.008029f
C374 B.n334 VSUBS 0.008029f
C375 B.n335 VSUBS 0.008029f
C376 B.n336 VSUBS 0.008029f
C377 B.n337 VSUBS 0.008029f
C378 B.n338 VSUBS 0.008029f
C379 B.n339 VSUBS 0.008029f
C380 B.n340 VSUBS 0.008029f
C381 B.n341 VSUBS 0.008029f
C382 B.n342 VSUBS 0.008029f
C383 B.n343 VSUBS 0.008029f
C384 B.n344 VSUBS 0.008029f
C385 B.n345 VSUBS 0.008029f
C386 B.n346 VSUBS 0.008029f
C387 B.n347 VSUBS 0.008029f
C388 B.n348 VSUBS 0.008029f
C389 B.n349 VSUBS 0.008029f
C390 B.n350 VSUBS 0.008029f
C391 B.n351 VSUBS 0.008029f
C392 B.n352 VSUBS 0.008029f
C393 B.n353 VSUBS 0.008029f
C394 B.n354 VSUBS 0.008029f
C395 B.n355 VSUBS 0.008029f
C396 B.n356 VSUBS 0.008029f
C397 B.n357 VSUBS 0.008029f
C398 B.n358 VSUBS 0.008029f
C399 B.n359 VSUBS 0.008029f
C400 B.n360 VSUBS 0.008029f
C401 B.n361 VSUBS 0.008029f
C402 B.n362 VSUBS 0.008029f
C403 B.n363 VSUBS 0.008029f
C404 B.n364 VSUBS 0.008029f
C405 B.n365 VSUBS 0.008029f
C406 B.n366 VSUBS 0.008029f
C407 B.n367 VSUBS 0.008029f
C408 B.n368 VSUBS 0.008029f
C409 B.n369 VSUBS 0.008029f
C410 B.n370 VSUBS 0.008029f
C411 B.n371 VSUBS 0.008029f
C412 B.n372 VSUBS 0.008029f
C413 B.n373 VSUBS 0.008029f
C414 B.n374 VSUBS 0.008029f
C415 B.n375 VSUBS 0.008029f
C416 B.n376 VSUBS 0.008029f
C417 B.n377 VSUBS 0.008029f
C418 B.n378 VSUBS 0.008029f
C419 B.n379 VSUBS 0.008029f
C420 B.n380 VSUBS 0.008029f
C421 B.n381 VSUBS 0.017463f
C422 B.n382 VSUBS 0.018481f
C423 B.n383 VSUBS 0.017413f
C424 B.n384 VSUBS 0.008029f
C425 B.n385 VSUBS 0.008029f
C426 B.n386 VSUBS 0.008029f
C427 B.n387 VSUBS 0.008029f
C428 B.n388 VSUBS 0.008029f
C429 B.n389 VSUBS 0.008029f
C430 B.n390 VSUBS 0.008029f
C431 B.n391 VSUBS 0.008029f
C432 B.n392 VSUBS 0.008029f
C433 B.n393 VSUBS 0.008029f
C434 B.n394 VSUBS 0.008029f
C435 B.n395 VSUBS 0.008029f
C436 B.n396 VSUBS 0.008029f
C437 B.n397 VSUBS 0.008029f
C438 B.n398 VSUBS 0.008029f
C439 B.n399 VSUBS 0.008029f
C440 B.n400 VSUBS 0.008029f
C441 B.n401 VSUBS 0.008029f
C442 B.n402 VSUBS 0.008029f
C443 B.n403 VSUBS 0.008029f
C444 B.n404 VSUBS 0.008029f
C445 B.n405 VSUBS 0.008029f
C446 B.n406 VSUBS 0.008029f
C447 B.n407 VSUBS 0.008029f
C448 B.n408 VSUBS 0.008029f
C449 B.n409 VSUBS 0.008029f
C450 B.n410 VSUBS 0.008029f
C451 B.n411 VSUBS 0.008029f
C452 B.n412 VSUBS 0.008029f
C453 B.n413 VSUBS 0.008029f
C454 B.n414 VSUBS 0.008029f
C455 B.n415 VSUBS 0.008029f
C456 B.n416 VSUBS 0.008029f
C457 B.n417 VSUBS 0.008029f
C458 B.n418 VSUBS 0.008029f
C459 B.n419 VSUBS 0.008029f
C460 B.n420 VSUBS 0.007557f
C461 B.n421 VSUBS 0.008029f
C462 B.n422 VSUBS 0.008029f
C463 B.n423 VSUBS 0.008029f
C464 B.n424 VSUBS 0.008029f
C465 B.n425 VSUBS 0.008029f
C466 B.n426 VSUBS 0.008029f
C467 B.n427 VSUBS 0.008029f
C468 B.n428 VSUBS 0.008029f
C469 B.n429 VSUBS 0.008029f
C470 B.n430 VSUBS 0.008029f
C471 B.n431 VSUBS 0.008029f
C472 B.n432 VSUBS 0.008029f
C473 B.n433 VSUBS 0.008029f
C474 B.n434 VSUBS 0.008029f
C475 B.n435 VSUBS 0.008029f
C476 B.n436 VSUBS 0.004487f
C477 B.n437 VSUBS 0.018602f
C478 B.n438 VSUBS 0.007557f
C479 B.n439 VSUBS 0.008029f
C480 B.n440 VSUBS 0.008029f
C481 B.n441 VSUBS 0.008029f
C482 B.n442 VSUBS 0.008029f
C483 B.n443 VSUBS 0.008029f
C484 B.n444 VSUBS 0.008029f
C485 B.n445 VSUBS 0.008029f
C486 B.n446 VSUBS 0.008029f
C487 B.n447 VSUBS 0.008029f
C488 B.n448 VSUBS 0.008029f
C489 B.n449 VSUBS 0.008029f
C490 B.n450 VSUBS 0.008029f
C491 B.n451 VSUBS 0.008029f
C492 B.n452 VSUBS 0.008029f
C493 B.n453 VSUBS 0.008029f
C494 B.n454 VSUBS 0.008029f
C495 B.n455 VSUBS 0.008029f
C496 B.n456 VSUBS 0.008029f
C497 B.n457 VSUBS 0.008029f
C498 B.n458 VSUBS 0.008029f
C499 B.n459 VSUBS 0.008029f
C500 B.n460 VSUBS 0.008029f
C501 B.n461 VSUBS 0.008029f
C502 B.n462 VSUBS 0.008029f
C503 B.n463 VSUBS 0.008029f
C504 B.n464 VSUBS 0.008029f
C505 B.n465 VSUBS 0.008029f
C506 B.n466 VSUBS 0.008029f
C507 B.n467 VSUBS 0.008029f
C508 B.n468 VSUBS 0.008029f
C509 B.n469 VSUBS 0.008029f
C510 B.n470 VSUBS 0.008029f
C511 B.n471 VSUBS 0.008029f
C512 B.n472 VSUBS 0.008029f
C513 B.n473 VSUBS 0.008029f
C514 B.n474 VSUBS 0.008029f
C515 B.n475 VSUBS 0.018431f
C516 B.n476 VSUBS 0.018431f
C517 B.n477 VSUBS 0.017463f
C518 B.n478 VSUBS 0.008029f
C519 B.n479 VSUBS 0.008029f
C520 B.n480 VSUBS 0.008029f
C521 B.n481 VSUBS 0.008029f
C522 B.n482 VSUBS 0.008029f
C523 B.n483 VSUBS 0.008029f
C524 B.n484 VSUBS 0.008029f
C525 B.n485 VSUBS 0.008029f
C526 B.n486 VSUBS 0.008029f
C527 B.n487 VSUBS 0.008029f
C528 B.n488 VSUBS 0.008029f
C529 B.n489 VSUBS 0.008029f
C530 B.n490 VSUBS 0.008029f
C531 B.n491 VSUBS 0.008029f
C532 B.n492 VSUBS 0.008029f
C533 B.n493 VSUBS 0.008029f
C534 B.n494 VSUBS 0.008029f
C535 B.n495 VSUBS 0.008029f
C536 B.n496 VSUBS 0.008029f
C537 B.n497 VSUBS 0.008029f
C538 B.n498 VSUBS 0.008029f
C539 B.n499 VSUBS 0.008029f
C540 B.n500 VSUBS 0.008029f
C541 B.n501 VSUBS 0.008029f
C542 B.n502 VSUBS 0.008029f
C543 B.n503 VSUBS 0.008029f
C544 B.n504 VSUBS 0.008029f
C545 B.n505 VSUBS 0.008029f
C546 B.n506 VSUBS 0.008029f
C547 B.n507 VSUBS 0.008029f
C548 B.n508 VSUBS 0.008029f
C549 B.n509 VSUBS 0.008029f
C550 B.n510 VSUBS 0.008029f
C551 B.n511 VSUBS 0.008029f
C552 B.n512 VSUBS 0.008029f
C553 B.n513 VSUBS 0.008029f
C554 B.n514 VSUBS 0.008029f
C555 B.n515 VSUBS 0.008029f
C556 B.n516 VSUBS 0.008029f
C557 B.n517 VSUBS 0.008029f
C558 B.n518 VSUBS 0.008029f
C559 B.n519 VSUBS 0.008029f
C560 B.n520 VSUBS 0.008029f
C561 B.n521 VSUBS 0.008029f
C562 B.n522 VSUBS 0.008029f
C563 B.n523 VSUBS 0.008029f
C564 B.n524 VSUBS 0.008029f
C565 B.n525 VSUBS 0.008029f
C566 B.n526 VSUBS 0.008029f
C567 B.n527 VSUBS 0.01818f
C568 VDD1.t3 VSUBS 0.146732f
C569 VDD1.t2 VSUBS 0.146732f
C570 VDD1.n0 VSUBS 1.00331f
C571 VDD1.t1 VSUBS 0.146732f
C572 VDD1.t0 VSUBS 0.146732f
C573 VDD1.n1 VSUBS 1.49065f
C574 VP.n0 VSUBS 0.054931f
C575 VP.t3 VSUBS 1.85232f
C576 VP.n1 VSUBS 0.060823f
C577 VP.n2 VSUBS 0.041665f
C578 VP.t2 VSUBS 1.85232f
C579 VP.n3 VSUBS 0.815495f
C580 VP.t1 VSUBS 2.17701f
C581 VP.t0 VSUBS 2.18399f
C582 VP.n4 VSUBS 3.31786f
C583 VP.n5 VSUBS 2.01402f
C584 VP.n6 VSUBS 0.054931f
C585 VP.n7 VSUBS 0.051198f
C586 VP.n8 VSUBS 0.077653f
C587 VP.n9 VSUBS 0.060823f
C588 VP.n10 VSUBS 0.041665f
C589 VP.n11 VSUBS 0.041665f
C590 VP.n12 VSUBS 0.041665f
C591 VP.n13 VSUBS 0.077653f
C592 VP.n14 VSUBS 0.051198f
C593 VP.n15 VSUBS 0.815495f
C594 VP.n16 VSUBS 0.068546f
C595 VTAIL.n0 VSUBS 0.029836f
C596 VTAIL.n1 VSUBS 0.026739f
C597 VTAIL.n2 VSUBS 0.014368f
C598 VTAIL.n3 VSUBS 0.033962f
C599 VTAIL.n4 VSUBS 0.015214f
C600 VTAIL.n5 VSUBS 0.026739f
C601 VTAIL.n6 VSUBS 0.014368f
C602 VTAIL.n7 VSUBS 0.033962f
C603 VTAIL.n8 VSUBS 0.015214f
C604 VTAIL.n9 VSUBS 0.70249f
C605 VTAIL.n10 VSUBS 0.014368f
C606 VTAIL.t5 VSUBS 0.072655f
C607 VTAIL.n11 VSUBS 0.123747f
C608 VTAIL.n12 VSUBS 0.021601f
C609 VTAIL.n13 VSUBS 0.025471f
C610 VTAIL.n14 VSUBS 0.033962f
C611 VTAIL.n15 VSUBS 0.015214f
C612 VTAIL.n16 VSUBS 0.014368f
C613 VTAIL.n17 VSUBS 0.026739f
C614 VTAIL.n18 VSUBS 0.026739f
C615 VTAIL.n19 VSUBS 0.014368f
C616 VTAIL.n20 VSUBS 0.015214f
C617 VTAIL.n21 VSUBS 0.033962f
C618 VTAIL.n22 VSUBS 0.033962f
C619 VTAIL.n23 VSUBS 0.015214f
C620 VTAIL.n24 VSUBS 0.014368f
C621 VTAIL.n25 VSUBS 0.026739f
C622 VTAIL.n26 VSUBS 0.026739f
C623 VTAIL.n27 VSUBS 0.014368f
C624 VTAIL.n28 VSUBS 0.015214f
C625 VTAIL.n29 VSUBS 0.033962f
C626 VTAIL.n30 VSUBS 0.083768f
C627 VTAIL.n31 VSUBS 0.015214f
C628 VTAIL.n32 VSUBS 0.014368f
C629 VTAIL.n33 VSUBS 0.062172f
C630 VTAIL.n34 VSUBS 0.042206f
C631 VTAIL.n35 VSUBS 0.172895f
C632 VTAIL.n36 VSUBS 0.029836f
C633 VTAIL.n37 VSUBS 0.026739f
C634 VTAIL.n38 VSUBS 0.014368f
C635 VTAIL.n39 VSUBS 0.033962f
C636 VTAIL.n40 VSUBS 0.015214f
C637 VTAIL.n41 VSUBS 0.026739f
C638 VTAIL.n42 VSUBS 0.014368f
C639 VTAIL.n43 VSUBS 0.033962f
C640 VTAIL.n44 VSUBS 0.015214f
C641 VTAIL.n45 VSUBS 0.70249f
C642 VTAIL.n46 VSUBS 0.014368f
C643 VTAIL.t1 VSUBS 0.072655f
C644 VTAIL.n47 VSUBS 0.123747f
C645 VTAIL.n48 VSUBS 0.021601f
C646 VTAIL.n49 VSUBS 0.025471f
C647 VTAIL.n50 VSUBS 0.033962f
C648 VTAIL.n51 VSUBS 0.015214f
C649 VTAIL.n52 VSUBS 0.014368f
C650 VTAIL.n53 VSUBS 0.026739f
C651 VTAIL.n54 VSUBS 0.026739f
C652 VTAIL.n55 VSUBS 0.014368f
C653 VTAIL.n56 VSUBS 0.015214f
C654 VTAIL.n57 VSUBS 0.033962f
C655 VTAIL.n58 VSUBS 0.033962f
C656 VTAIL.n59 VSUBS 0.015214f
C657 VTAIL.n60 VSUBS 0.014368f
C658 VTAIL.n61 VSUBS 0.026739f
C659 VTAIL.n62 VSUBS 0.026739f
C660 VTAIL.n63 VSUBS 0.014368f
C661 VTAIL.n64 VSUBS 0.015214f
C662 VTAIL.n65 VSUBS 0.033962f
C663 VTAIL.n66 VSUBS 0.083768f
C664 VTAIL.n67 VSUBS 0.015214f
C665 VTAIL.n68 VSUBS 0.014368f
C666 VTAIL.n69 VSUBS 0.062172f
C667 VTAIL.n70 VSUBS 0.042206f
C668 VTAIL.n71 VSUBS 0.272238f
C669 VTAIL.n72 VSUBS 0.029836f
C670 VTAIL.n73 VSUBS 0.026739f
C671 VTAIL.n74 VSUBS 0.014368f
C672 VTAIL.n75 VSUBS 0.033962f
C673 VTAIL.n76 VSUBS 0.015214f
C674 VTAIL.n77 VSUBS 0.026739f
C675 VTAIL.n78 VSUBS 0.014368f
C676 VTAIL.n79 VSUBS 0.033962f
C677 VTAIL.n80 VSUBS 0.015214f
C678 VTAIL.n81 VSUBS 0.70249f
C679 VTAIL.n82 VSUBS 0.014368f
C680 VTAIL.t0 VSUBS 0.072655f
C681 VTAIL.n83 VSUBS 0.123747f
C682 VTAIL.n84 VSUBS 0.021601f
C683 VTAIL.n85 VSUBS 0.025471f
C684 VTAIL.n86 VSUBS 0.033962f
C685 VTAIL.n87 VSUBS 0.015214f
C686 VTAIL.n88 VSUBS 0.014368f
C687 VTAIL.n89 VSUBS 0.026739f
C688 VTAIL.n90 VSUBS 0.026739f
C689 VTAIL.n91 VSUBS 0.014368f
C690 VTAIL.n92 VSUBS 0.015214f
C691 VTAIL.n93 VSUBS 0.033962f
C692 VTAIL.n94 VSUBS 0.033962f
C693 VTAIL.n95 VSUBS 0.015214f
C694 VTAIL.n96 VSUBS 0.014368f
C695 VTAIL.n97 VSUBS 0.026739f
C696 VTAIL.n98 VSUBS 0.026739f
C697 VTAIL.n99 VSUBS 0.014368f
C698 VTAIL.n100 VSUBS 0.015214f
C699 VTAIL.n101 VSUBS 0.033962f
C700 VTAIL.n102 VSUBS 0.083768f
C701 VTAIL.n103 VSUBS 0.015214f
C702 VTAIL.n104 VSUBS 0.014368f
C703 VTAIL.n105 VSUBS 0.062172f
C704 VTAIL.n106 VSUBS 0.042206f
C705 VTAIL.n107 VSUBS 1.30357f
C706 VTAIL.n108 VSUBS 0.029836f
C707 VTAIL.n109 VSUBS 0.026739f
C708 VTAIL.n110 VSUBS 0.014368f
C709 VTAIL.n111 VSUBS 0.033962f
C710 VTAIL.n112 VSUBS 0.015214f
C711 VTAIL.n113 VSUBS 0.026739f
C712 VTAIL.n114 VSUBS 0.014368f
C713 VTAIL.n115 VSUBS 0.033962f
C714 VTAIL.n116 VSUBS 0.015214f
C715 VTAIL.n117 VSUBS 0.70249f
C716 VTAIL.n118 VSUBS 0.014368f
C717 VTAIL.t6 VSUBS 0.072655f
C718 VTAIL.n119 VSUBS 0.123747f
C719 VTAIL.n120 VSUBS 0.021601f
C720 VTAIL.n121 VSUBS 0.025471f
C721 VTAIL.n122 VSUBS 0.033962f
C722 VTAIL.n123 VSUBS 0.015214f
C723 VTAIL.n124 VSUBS 0.014368f
C724 VTAIL.n125 VSUBS 0.026739f
C725 VTAIL.n126 VSUBS 0.026739f
C726 VTAIL.n127 VSUBS 0.014368f
C727 VTAIL.n128 VSUBS 0.015214f
C728 VTAIL.n129 VSUBS 0.033962f
C729 VTAIL.n130 VSUBS 0.033962f
C730 VTAIL.n131 VSUBS 0.015214f
C731 VTAIL.n132 VSUBS 0.014368f
C732 VTAIL.n133 VSUBS 0.026739f
C733 VTAIL.n134 VSUBS 0.026739f
C734 VTAIL.n135 VSUBS 0.014368f
C735 VTAIL.n136 VSUBS 0.015214f
C736 VTAIL.n137 VSUBS 0.033962f
C737 VTAIL.n138 VSUBS 0.083768f
C738 VTAIL.n139 VSUBS 0.015214f
C739 VTAIL.n140 VSUBS 0.014368f
C740 VTAIL.n141 VSUBS 0.062172f
C741 VTAIL.n142 VSUBS 0.042206f
C742 VTAIL.n143 VSUBS 1.30357f
C743 VTAIL.n144 VSUBS 0.029836f
C744 VTAIL.n145 VSUBS 0.026739f
C745 VTAIL.n146 VSUBS 0.014368f
C746 VTAIL.n147 VSUBS 0.033962f
C747 VTAIL.n148 VSUBS 0.015214f
C748 VTAIL.n149 VSUBS 0.026739f
C749 VTAIL.n150 VSUBS 0.014368f
C750 VTAIL.n151 VSUBS 0.033962f
C751 VTAIL.n152 VSUBS 0.015214f
C752 VTAIL.n153 VSUBS 0.70249f
C753 VTAIL.n154 VSUBS 0.014368f
C754 VTAIL.t4 VSUBS 0.072655f
C755 VTAIL.n155 VSUBS 0.123747f
C756 VTAIL.n156 VSUBS 0.021601f
C757 VTAIL.n157 VSUBS 0.025471f
C758 VTAIL.n158 VSUBS 0.033962f
C759 VTAIL.n159 VSUBS 0.015214f
C760 VTAIL.n160 VSUBS 0.014368f
C761 VTAIL.n161 VSUBS 0.026739f
C762 VTAIL.n162 VSUBS 0.026739f
C763 VTAIL.n163 VSUBS 0.014368f
C764 VTAIL.n164 VSUBS 0.015214f
C765 VTAIL.n165 VSUBS 0.033962f
C766 VTAIL.n166 VSUBS 0.033962f
C767 VTAIL.n167 VSUBS 0.015214f
C768 VTAIL.n168 VSUBS 0.014368f
C769 VTAIL.n169 VSUBS 0.026739f
C770 VTAIL.n170 VSUBS 0.026739f
C771 VTAIL.n171 VSUBS 0.014368f
C772 VTAIL.n172 VSUBS 0.015214f
C773 VTAIL.n173 VSUBS 0.033962f
C774 VTAIL.n174 VSUBS 0.083768f
C775 VTAIL.n175 VSUBS 0.015214f
C776 VTAIL.n176 VSUBS 0.014368f
C777 VTAIL.n177 VSUBS 0.062172f
C778 VTAIL.n178 VSUBS 0.042206f
C779 VTAIL.n179 VSUBS 0.272238f
C780 VTAIL.n180 VSUBS 0.029836f
C781 VTAIL.n181 VSUBS 0.026739f
C782 VTAIL.n182 VSUBS 0.014368f
C783 VTAIL.n183 VSUBS 0.033962f
C784 VTAIL.n184 VSUBS 0.015214f
C785 VTAIL.n185 VSUBS 0.026739f
C786 VTAIL.n186 VSUBS 0.014368f
C787 VTAIL.n187 VSUBS 0.033962f
C788 VTAIL.n188 VSUBS 0.015214f
C789 VTAIL.n189 VSUBS 0.70249f
C790 VTAIL.n190 VSUBS 0.014368f
C791 VTAIL.t2 VSUBS 0.072655f
C792 VTAIL.n191 VSUBS 0.123747f
C793 VTAIL.n192 VSUBS 0.021601f
C794 VTAIL.n193 VSUBS 0.025471f
C795 VTAIL.n194 VSUBS 0.033962f
C796 VTAIL.n195 VSUBS 0.015214f
C797 VTAIL.n196 VSUBS 0.014368f
C798 VTAIL.n197 VSUBS 0.026739f
C799 VTAIL.n198 VSUBS 0.026739f
C800 VTAIL.n199 VSUBS 0.014368f
C801 VTAIL.n200 VSUBS 0.015214f
C802 VTAIL.n201 VSUBS 0.033962f
C803 VTAIL.n202 VSUBS 0.033962f
C804 VTAIL.n203 VSUBS 0.015214f
C805 VTAIL.n204 VSUBS 0.014368f
C806 VTAIL.n205 VSUBS 0.026739f
C807 VTAIL.n206 VSUBS 0.026739f
C808 VTAIL.n207 VSUBS 0.014368f
C809 VTAIL.n208 VSUBS 0.015214f
C810 VTAIL.n209 VSUBS 0.033962f
C811 VTAIL.n210 VSUBS 0.083768f
C812 VTAIL.n211 VSUBS 0.015214f
C813 VTAIL.n212 VSUBS 0.014368f
C814 VTAIL.n213 VSUBS 0.062172f
C815 VTAIL.n214 VSUBS 0.042206f
C816 VTAIL.n215 VSUBS 0.272238f
C817 VTAIL.n216 VSUBS 0.029836f
C818 VTAIL.n217 VSUBS 0.026739f
C819 VTAIL.n218 VSUBS 0.014368f
C820 VTAIL.n219 VSUBS 0.033962f
C821 VTAIL.n220 VSUBS 0.015214f
C822 VTAIL.n221 VSUBS 0.026739f
C823 VTAIL.n222 VSUBS 0.014368f
C824 VTAIL.n223 VSUBS 0.033962f
C825 VTAIL.n224 VSUBS 0.015214f
C826 VTAIL.n225 VSUBS 0.70249f
C827 VTAIL.n226 VSUBS 0.014368f
C828 VTAIL.t7 VSUBS 0.072655f
C829 VTAIL.n227 VSUBS 0.123747f
C830 VTAIL.n228 VSUBS 0.021601f
C831 VTAIL.n229 VSUBS 0.025471f
C832 VTAIL.n230 VSUBS 0.033962f
C833 VTAIL.n231 VSUBS 0.015214f
C834 VTAIL.n232 VSUBS 0.014368f
C835 VTAIL.n233 VSUBS 0.026739f
C836 VTAIL.n234 VSUBS 0.026739f
C837 VTAIL.n235 VSUBS 0.014368f
C838 VTAIL.n236 VSUBS 0.015214f
C839 VTAIL.n237 VSUBS 0.033962f
C840 VTAIL.n238 VSUBS 0.033962f
C841 VTAIL.n239 VSUBS 0.015214f
C842 VTAIL.n240 VSUBS 0.014368f
C843 VTAIL.n241 VSUBS 0.026739f
C844 VTAIL.n242 VSUBS 0.026739f
C845 VTAIL.n243 VSUBS 0.014368f
C846 VTAIL.n244 VSUBS 0.015214f
C847 VTAIL.n245 VSUBS 0.033962f
C848 VTAIL.n246 VSUBS 0.083768f
C849 VTAIL.n247 VSUBS 0.015214f
C850 VTAIL.n248 VSUBS 0.014368f
C851 VTAIL.n249 VSUBS 0.062172f
C852 VTAIL.n250 VSUBS 0.042206f
C853 VTAIL.n251 VSUBS 1.30357f
C854 VTAIL.n252 VSUBS 0.029836f
C855 VTAIL.n253 VSUBS 0.026739f
C856 VTAIL.n254 VSUBS 0.014368f
C857 VTAIL.n255 VSUBS 0.033962f
C858 VTAIL.n256 VSUBS 0.015214f
C859 VTAIL.n257 VSUBS 0.026739f
C860 VTAIL.n258 VSUBS 0.014368f
C861 VTAIL.n259 VSUBS 0.033962f
C862 VTAIL.n260 VSUBS 0.015214f
C863 VTAIL.n261 VSUBS 0.70249f
C864 VTAIL.n262 VSUBS 0.014368f
C865 VTAIL.t3 VSUBS 0.072655f
C866 VTAIL.n263 VSUBS 0.123747f
C867 VTAIL.n264 VSUBS 0.021601f
C868 VTAIL.n265 VSUBS 0.025471f
C869 VTAIL.n266 VSUBS 0.033962f
C870 VTAIL.n267 VSUBS 0.015214f
C871 VTAIL.n268 VSUBS 0.014368f
C872 VTAIL.n269 VSUBS 0.026739f
C873 VTAIL.n270 VSUBS 0.026739f
C874 VTAIL.n271 VSUBS 0.014368f
C875 VTAIL.n272 VSUBS 0.015214f
C876 VTAIL.n273 VSUBS 0.033962f
C877 VTAIL.n274 VSUBS 0.033962f
C878 VTAIL.n275 VSUBS 0.015214f
C879 VTAIL.n276 VSUBS 0.014368f
C880 VTAIL.n277 VSUBS 0.026739f
C881 VTAIL.n278 VSUBS 0.026739f
C882 VTAIL.n279 VSUBS 0.014368f
C883 VTAIL.n280 VSUBS 0.015214f
C884 VTAIL.n281 VSUBS 0.033962f
C885 VTAIL.n282 VSUBS 0.083768f
C886 VTAIL.n283 VSUBS 0.015214f
C887 VTAIL.n284 VSUBS 0.014368f
C888 VTAIL.n285 VSUBS 0.062172f
C889 VTAIL.n286 VSUBS 0.042206f
C890 VTAIL.n287 VSUBS 1.1942f
C891 VDD2.t2 VSUBS 0.146772f
C892 VDD2.t3 VSUBS 0.146772f
C893 VDD2.n0 VSUBS 1.46991f
C894 VDD2.t0 VSUBS 0.146772f
C895 VDD2.t1 VSUBS 0.146772f
C896 VDD2.n1 VSUBS 1.00312f
C897 VDD2.n2 VSUBS 3.71852f
C898 VN.t1 VSUBS 2.10707f
C899 VN.t3 VSUBS 2.10033f
C900 VN.n0 VSUBS 1.34736f
C901 VN.t2 VSUBS 2.10707f
C902 VN.t0 VSUBS 2.10033f
C903 VN.n1 VSUBS 3.22232f
.ends

