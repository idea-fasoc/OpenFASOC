* NGSPICE file created from diff_pair_sample_0400.ext - technology: sky130A

.subckt diff_pair_sample_0400 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t5 VN.t0 VTAIL.t10 B.t0 sky130_fd_pr__nfet_01v8 ad=3.2331 pd=17.36 as=1.36785 ps=8.62 w=8.29 l=1.23
X1 VTAIL.t2 VP.t0 VDD1.t5 B.t2 sky130_fd_pr__nfet_01v8 ad=1.36785 pd=8.62 as=1.36785 ps=8.62 w=8.29 l=1.23
X2 B.t18 B.t16 B.t17 B.t13 sky130_fd_pr__nfet_01v8 ad=3.2331 pd=17.36 as=0 ps=0 w=8.29 l=1.23
X3 VDD1.t4 VP.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=3.2331 pd=17.36 as=1.36785 ps=8.62 w=8.29 l=1.23
X4 VTAIL.t11 VP.t2 VDD1.t3 B.t19 sky130_fd_pr__nfet_01v8 ad=1.36785 pd=8.62 as=1.36785 ps=8.62 w=8.29 l=1.23
X5 VDD1.t2 VP.t3 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.36785 pd=8.62 as=3.2331 ps=17.36 w=8.29 l=1.23
X6 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=3.2331 pd=17.36 as=0 ps=0 w=8.29 l=1.23
X7 VDD1.t1 VP.t4 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.36785 pd=8.62 as=3.2331 ps=17.36 w=8.29 l=1.23
X8 VDD2.t4 VN.t1 VTAIL.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=1.36785 pd=8.62 as=3.2331 ps=17.36 w=8.29 l=1.23
X9 VDD2.t3 VN.t2 VTAIL.t9 B.t4 sky130_fd_pr__nfet_01v8 ad=1.36785 pd=8.62 as=3.2331 ps=17.36 w=8.29 l=1.23
X10 VTAIL.t8 VN.t3 VDD2.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.36785 pd=8.62 as=1.36785 ps=8.62 w=8.29 l=1.23
X11 VTAIL.t5 VN.t4 VDD2.t1 B.t19 sky130_fd_pr__nfet_01v8 ad=1.36785 pd=8.62 as=1.36785 ps=8.62 w=8.29 l=1.23
X12 B.t11 B.t9 B.t10 B.t6 sky130_fd_pr__nfet_01v8 ad=3.2331 pd=17.36 as=0 ps=0 w=8.29 l=1.23
X13 VDD2.t0 VN.t5 VTAIL.t7 B.t1 sky130_fd_pr__nfet_01v8 ad=3.2331 pd=17.36 as=1.36785 ps=8.62 w=8.29 l=1.23
X14 VDD1.t0 VP.t5 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=3.2331 pd=17.36 as=1.36785 ps=8.62 w=8.29 l=1.23
X15 B.t8 B.t5 B.t7 B.t6 sky130_fd_pr__nfet_01v8 ad=3.2331 pd=17.36 as=0 ps=0 w=8.29 l=1.23
R0 VN.n2 VN.t5 213.067
R1 VN.n10 VN.t1 213.067
R2 VN.n6 VN.t2 194.564
R3 VN.n14 VN.t0 194.564
R4 VN.n1 VN.t3 162.43
R5 VN.n9 VN.t4 162.43
R6 VN.n13 VN.n8 161.3
R7 VN.n12 VN.n11 161.3
R8 VN.n5 VN.n0 161.3
R9 VN.n4 VN.n3 161.3
R10 VN.n15 VN.n14 80.6037
R11 VN.n7 VN.n6 80.6037
R12 VN.n2 VN.n1 45.5344
R13 VN.n10 VN.n9 45.5344
R14 VN VN.n15 40.9081
R15 VN.n5 VN.n4 37.5796
R16 VN.n13 VN.n12 37.5796
R17 VN.n11 VN.n10 29.7304
R18 VN.n3 VN.n2 29.7304
R19 VN.n6 VN.n5 28.4823
R20 VN.n14 VN.n13 28.4823
R21 VN.n4 VN.n1 12.234
R22 VN.n12 VN.n9 12.234
R23 VN.n15 VN.n8 0.285035
R24 VN.n7 VN.n0 0.285035
R25 VN.n11 VN.n8 0.189894
R26 VN.n3 VN.n0 0.189894
R27 VN VN.n7 0.146778
R28 VTAIL.n7 VTAIL.t6 51.9265
R29 VTAIL.n10 VTAIL.t4 51.9264
R30 VTAIL.n11 VTAIL.t9 51.9264
R31 VTAIL.n2 VTAIL.t3 51.9264
R32 VTAIL.n9 VTAIL.n8 49.5381
R33 VTAIL.n6 VTAIL.n5 49.5381
R34 VTAIL.n1 VTAIL.n0 49.5379
R35 VTAIL.n4 VTAIL.n3 49.5379
R36 VTAIL.n6 VTAIL.n4 22.2031
R37 VTAIL.n11 VTAIL.n10 20.8583
R38 VTAIL.n0 VTAIL.t7 2.38892
R39 VTAIL.n0 VTAIL.t8 2.38892
R40 VTAIL.n3 VTAIL.t0 2.38892
R41 VTAIL.n3 VTAIL.t11 2.38892
R42 VTAIL.n8 VTAIL.t1 2.38892
R43 VTAIL.n8 VTAIL.t2 2.38892
R44 VTAIL.n5 VTAIL.t10 2.38892
R45 VTAIL.n5 VTAIL.t5 2.38892
R46 VTAIL.n7 VTAIL.n6 1.34533
R47 VTAIL.n10 VTAIL.n9 1.34533
R48 VTAIL.n4 VTAIL.n2 1.34533
R49 VTAIL.n9 VTAIL.n7 1.14274
R50 VTAIL.n2 VTAIL.n1 1.14274
R51 VTAIL VTAIL.n11 0.950931
R52 VTAIL VTAIL.n1 0.394897
R53 VDD2.n1 VDD2.t0 69.5585
R54 VDD2.n2 VDD2.t5 68.6053
R55 VDD2.n1 VDD2.n0 66.4975
R56 VDD2 VDD2.n3 66.4948
R57 VDD2.n2 VDD2.n1 35.2325
R58 VDD2.n3 VDD2.t1 2.38892
R59 VDD2.n3 VDD2.t4 2.38892
R60 VDD2.n0 VDD2.t2 2.38892
R61 VDD2.n0 VDD2.t3 2.38892
R62 VDD2 VDD2.n2 1.06731
R63 B.n439 B.n438 585
R64 B.n439 B.n50 585
R65 B.n442 B.n441 585
R66 B.n443 B.n90 585
R67 B.n445 B.n444 585
R68 B.n447 B.n89 585
R69 B.n450 B.n449 585
R70 B.n451 B.n88 585
R71 B.n453 B.n452 585
R72 B.n455 B.n87 585
R73 B.n458 B.n457 585
R74 B.n459 B.n86 585
R75 B.n461 B.n460 585
R76 B.n463 B.n85 585
R77 B.n466 B.n465 585
R78 B.n467 B.n84 585
R79 B.n469 B.n468 585
R80 B.n471 B.n83 585
R81 B.n474 B.n473 585
R82 B.n475 B.n82 585
R83 B.n477 B.n476 585
R84 B.n479 B.n81 585
R85 B.n482 B.n481 585
R86 B.n483 B.n80 585
R87 B.n485 B.n484 585
R88 B.n487 B.n79 585
R89 B.n490 B.n489 585
R90 B.n491 B.n78 585
R91 B.n493 B.n492 585
R92 B.n495 B.n77 585
R93 B.n498 B.n497 585
R94 B.n499 B.n74 585
R95 B.n502 B.n501 585
R96 B.n504 B.n73 585
R97 B.n507 B.n506 585
R98 B.n508 B.n72 585
R99 B.n510 B.n509 585
R100 B.n512 B.n71 585
R101 B.n515 B.n514 585
R102 B.n516 B.n67 585
R103 B.n518 B.n517 585
R104 B.n520 B.n66 585
R105 B.n523 B.n522 585
R106 B.n524 B.n65 585
R107 B.n526 B.n525 585
R108 B.n528 B.n64 585
R109 B.n531 B.n530 585
R110 B.n532 B.n63 585
R111 B.n534 B.n533 585
R112 B.n536 B.n62 585
R113 B.n539 B.n538 585
R114 B.n540 B.n61 585
R115 B.n542 B.n541 585
R116 B.n544 B.n60 585
R117 B.n547 B.n546 585
R118 B.n548 B.n59 585
R119 B.n550 B.n549 585
R120 B.n552 B.n58 585
R121 B.n555 B.n554 585
R122 B.n556 B.n57 585
R123 B.n558 B.n557 585
R124 B.n560 B.n56 585
R125 B.n563 B.n562 585
R126 B.n564 B.n55 585
R127 B.n566 B.n565 585
R128 B.n568 B.n54 585
R129 B.n571 B.n570 585
R130 B.n572 B.n53 585
R131 B.n574 B.n573 585
R132 B.n576 B.n52 585
R133 B.n579 B.n578 585
R134 B.n580 B.n51 585
R135 B.n437 B.n49 585
R136 B.n583 B.n49 585
R137 B.n436 B.n48 585
R138 B.n584 B.n48 585
R139 B.n435 B.n47 585
R140 B.n585 B.n47 585
R141 B.n434 B.n433 585
R142 B.n433 B.n43 585
R143 B.n432 B.n42 585
R144 B.n591 B.n42 585
R145 B.n431 B.n41 585
R146 B.n592 B.n41 585
R147 B.n430 B.n40 585
R148 B.n593 B.n40 585
R149 B.n429 B.n428 585
R150 B.n428 B.n36 585
R151 B.n427 B.n35 585
R152 B.n599 B.n35 585
R153 B.n426 B.n34 585
R154 B.n600 B.n34 585
R155 B.n425 B.n33 585
R156 B.n601 B.n33 585
R157 B.n424 B.n423 585
R158 B.n423 B.n29 585
R159 B.n422 B.n28 585
R160 B.n607 B.n28 585
R161 B.n421 B.n27 585
R162 B.n608 B.n27 585
R163 B.n420 B.n26 585
R164 B.n609 B.n26 585
R165 B.n419 B.n418 585
R166 B.n418 B.n22 585
R167 B.n417 B.n21 585
R168 B.n615 B.n21 585
R169 B.n416 B.n20 585
R170 B.n616 B.n20 585
R171 B.n415 B.n19 585
R172 B.n617 B.n19 585
R173 B.n414 B.n413 585
R174 B.n413 B.n15 585
R175 B.n412 B.n14 585
R176 B.n623 B.n14 585
R177 B.n411 B.n13 585
R178 B.n624 B.n13 585
R179 B.n410 B.n12 585
R180 B.n625 B.n12 585
R181 B.n409 B.n408 585
R182 B.n408 B.n407 585
R183 B.n406 B.n405 585
R184 B.n406 B.n8 585
R185 B.n404 B.n7 585
R186 B.n632 B.n7 585
R187 B.n403 B.n6 585
R188 B.n633 B.n6 585
R189 B.n402 B.n5 585
R190 B.n634 B.n5 585
R191 B.n401 B.n400 585
R192 B.n400 B.n4 585
R193 B.n399 B.n91 585
R194 B.n399 B.n398 585
R195 B.n389 B.n92 585
R196 B.n93 B.n92 585
R197 B.n391 B.n390 585
R198 B.n392 B.n391 585
R199 B.n388 B.n98 585
R200 B.n98 B.n97 585
R201 B.n387 B.n386 585
R202 B.n386 B.n385 585
R203 B.n100 B.n99 585
R204 B.n101 B.n100 585
R205 B.n378 B.n377 585
R206 B.n379 B.n378 585
R207 B.n376 B.n106 585
R208 B.n106 B.n105 585
R209 B.n375 B.n374 585
R210 B.n374 B.n373 585
R211 B.n108 B.n107 585
R212 B.n109 B.n108 585
R213 B.n366 B.n365 585
R214 B.n367 B.n366 585
R215 B.n364 B.n113 585
R216 B.n117 B.n113 585
R217 B.n363 B.n362 585
R218 B.n362 B.n361 585
R219 B.n115 B.n114 585
R220 B.n116 B.n115 585
R221 B.n354 B.n353 585
R222 B.n355 B.n354 585
R223 B.n352 B.n122 585
R224 B.n122 B.n121 585
R225 B.n351 B.n350 585
R226 B.n350 B.n349 585
R227 B.n124 B.n123 585
R228 B.n125 B.n124 585
R229 B.n342 B.n341 585
R230 B.n343 B.n342 585
R231 B.n340 B.n129 585
R232 B.n133 B.n129 585
R233 B.n339 B.n338 585
R234 B.n338 B.n337 585
R235 B.n131 B.n130 585
R236 B.n132 B.n131 585
R237 B.n330 B.n329 585
R238 B.n331 B.n330 585
R239 B.n328 B.n138 585
R240 B.n138 B.n137 585
R241 B.n327 B.n326 585
R242 B.n326 B.n325 585
R243 B.n322 B.n142 585
R244 B.n321 B.n320 585
R245 B.n318 B.n143 585
R246 B.n318 B.n141 585
R247 B.n317 B.n316 585
R248 B.n315 B.n314 585
R249 B.n313 B.n145 585
R250 B.n311 B.n310 585
R251 B.n309 B.n146 585
R252 B.n308 B.n307 585
R253 B.n305 B.n147 585
R254 B.n303 B.n302 585
R255 B.n301 B.n148 585
R256 B.n300 B.n299 585
R257 B.n297 B.n149 585
R258 B.n295 B.n294 585
R259 B.n293 B.n150 585
R260 B.n292 B.n291 585
R261 B.n289 B.n151 585
R262 B.n287 B.n286 585
R263 B.n285 B.n152 585
R264 B.n284 B.n283 585
R265 B.n281 B.n153 585
R266 B.n279 B.n278 585
R267 B.n277 B.n154 585
R268 B.n276 B.n275 585
R269 B.n273 B.n155 585
R270 B.n271 B.n270 585
R271 B.n269 B.n156 585
R272 B.n268 B.n267 585
R273 B.n265 B.n157 585
R274 B.n263 B.n262 585
R275 B.n260 B.n158 585
R276 B.n259 B.n258 585
R277 B.n256 B.n161 585
R278 B.n254 B.n253 585
R279 B.n252 B.n162 585
R280 B.n251 B.n250 585
R281 B.n248 B.n163 585
R282 B.n246 B.n245 585
R283 B.n244 B.n164 585
R284 B.n242 B.n241 585
R285 B.n239 B.n167 585
R286 B.n237 B.n236 585
R287 B.n235 B.n168 585
R288 B.n234 B.n233 585
R289 B.n231 B.n169 585
R290 B.n229 B.n228 585
R291 B.n227 B.n170 585
R292 B.n226 B.n225 585
R293 B.n223 B.n171 585
R294 B.n221 B.n220 585
R295 B.n219 B.n172 585
R296 B.n218 B.n217 585
R297 B.n215 B.n173 585
R298 B.n213 B.n212 585
R299 B.n211 B.n174 585
R300 B.n210 B.n209 585
R301 B.n207 B.n175 585
R302 B.n205 B.n204 585
R303 B.n203 B.n176 585
R304 B.n202 B.n201 585
R305 B.n199 B.n177 585
R306 B.n197 B.n196 585
R307 B.n195 B.n178 585
R308 B.n194 B.n193 585
R309 B.n191 B.n179 585
R310 B.n189 B.n188 585
R311 B.n187 B.n180 585
R312 B.n186 B.n185 585
R313 B.n183 B.n181 585
R314 B.n140 B.n139 585
R315 B.n324 B.n323 585
R316 B.n325 B.n324 585
R317 B.n136 B.n135 585
R318 B.n137 B.n136 585
R319 B.n333 B.n332 585
R320 B.n332 B.n331 585
R321 B.n334 B.n134 585
R322 B.n134 B.n132 585
R323 B.n336 B.n335 585
R324 B.n337 B.n336 585
R325 B.n128 B.n127 585
R326 B.n133 B.n128 585
R327 B.n345 B.n344 585
R328 B.n344 B.n343 585
R329 B.n346 B.n126 585
R330 B.n126 B.n125 585
R331 B.n348 B.n347 585
R332 B.n349 B.n348 585
R333 B.n120 B.n119 585
R334 B.n121 B.n120 585
R335 B.n357 B.n356 585
R336 B.n356 B.n355 585
R337 B.n358 B.n118 585
R338 B.n118 B.n116 585
R339 B.n360 B.n359 585
R340 B.n361 B.n360 585
R341 B.n112 B.n111 585
R342 B.n117 B.n112 585
R343 B.n369 B.n368 585
R344 B.n368 B.n367 585
R345 B.n370 B.n110 585
R346 B.n110 B.n109 585
R347 B.n372 B.n371 585
R348 B.n373 B.n372 585
R349 B.n104 B.n103 585
R350 B.n105 B.n104 585
R351 B.n381 B.n380 585
R352 B.n380 B.n379 585
R353 B.n382 B.n102 585
R354 B.n102 B.n101 585
R355 B.n384 B.n383 585
R356 B.n385 B.n384 585
R357 B.n96 B.n95 585
R358 B.n97 B.n96 585
R359 B.n394 B.n393 585
R360 B.n393 B.n392 585
R361 B.n395 B.n94 585
R362 B.n94 B.n93 585
R363 B.n397 B.n396 585
R364 B.n398 B.n397 585
R365 B.n3 B.n0 585
R366 B.n4 B.n3 585
R367 B.n631 B.n1 585
R368 B.n632 B.n631 585
R369 B.n630 B.n629 585
R370 B.n630 B.n8 585
R371 B.n628 B.n9 585
R372 B.n407 B.n9 585
R373 B.n627 B.n626 585
R374 B.n626 B.n625 585
R375 B.n11 B.n10 585
R376 B.n624 B.n11 585
R377 B.n622 B.n621 585
R378 B.n623 B.n622 585
R379 B.n620 B.n16 585
R380 B.n16 B.n15 585
R381 B.n619 B.n618 585
R382 B.n618 B.n617 585
R383 B.n18 B.n17 585
R384 B.n616 B.n18 585
R385 B.n614 B.n613 585
R386 B.n615 B.n614 585
R387 B.n612 B.n23 585
R388 B.n23 B.n22 585
R389 B.n611 B.n610 585
R390 B.n610 B.n609 585
R391 B.n25 B.n24 585
R392 B.n608 B.n25 585
R393 B.n606 B.n605 585
R394 B.n607 B.n606 585
R395 B.n604 B.n30 585
R396 B.n30 B.n29 585
R397 B.n603 B.n602 585
R398 B.n602 B.n601 585
R399 B.n32 B.n31 585
R400 B.n600 B.n32 585
R401 B.n598 B.n597 585
R402 B.n599 B.n598 585
R403 B.n596 B.n37 585
R404 B.n37 B.n36 585
R405 B.n595 B.n594 585
R406 B.n594 B.n593 585
R407 B.n39 B.n38 585
R408 B.n592 B.n39 585
R409 B.n590 B.n589 585
R410 B.n591 B.n590 585
R411 B.n588 B.n44 585
R412 B.n44 B.n43 585
R413 B.n587 B.n586 585
R414 B.n586 B.n585 585
R415 B.n46 B.n45 585
R416 B.n584 B.n46 585
R417 B.n582 B.n581 585
R418 B.n583 B.n582 585
R419 B.n635 B.n634 585
R420 B.n633 B.n2 585
R421 B.n582 B.n51 492.5
R422 B.n439 B.n49 492.5
R423 B.n326 B.n140 492.5
R424 B.n324 B.n142 492.5
R425 B.n68 B.t16 366.702
R426 B.n75 B.t12 366.702
R427 B.n165 B.t5 366.702
R428 B.n159 B.t9 366.702
R429 B.n440 B.n50 256.663
R430 B.n446 B.n50 256.663
R431 B.n448 B.n50 256.663
R432 B.n454 B.n50 256.663
R433 B.n456 B.n50 256.663
R434 B.n462 B.n50 256.663
R435 B.n464 B.n50 256.663
R436 B.n470 B.n50 256.663
R437 B.n472 B.n50 256.663
R438 B.n478 B.n50 256.663
R439 B.n480 B.n50 256.663
R440 B.n486 B.n50 256.663
R441 B.n488 B.n50 256.663
R442 B.n494 B.n50 256.663
R443 B.n496 B.n50 256.663
R444 B.n503 B.n50 256.663
R445 B.n505 B.n50 256.663
R446 B.n511 B.n50 256.663
R447 B.n513 B.n50 256.663
R448 B.n519 B.n50 256.663
R449 B.n521 B.n50 256.663
R450 B.n527 B.n50 256.663
R451 B.n529 B.n50 256.663
R452 B.n535 B.n50 256.663
R453 B.n537 B.n50 256.663
R454 B.n543 B.n50 256.663
R455 B.n545 B.n50 256.663
R456 B.n551 B.n50 256.663
R457 B.n553 B.n50 256.663
R458 B.n559 B.n50 256.663
R459 B.n561 B.n50 256.663
R460 B.n567 B.n50 256.663
R461 B.n569 B.n50 256.663
R462 B.n575 B.n50 256.663
R463 B.n577 B.n50 256.663
R464 B.n319 B.n141 256.663
R465 B.n144 B.n141 256.663
R466 B.n312 B.n141 256.663
R467 B.n306 B.n141 256.663
R468 B.n304 B.n141 256.663
R469 B.n298 B.n141 256.663
R470 B.n296 B.n141 256.663
R471 B.n290 B.n141 256.663
R472 B.n288 B.n141 256.663
R473 B.n282 B.n141 256.663
R474 B.n280 B.n141 256.663
R475 B.n274 B.n141 256.663
R476 B.n272 B.n141 256.663
R477 B.n266 B.n141 256.663
R478 B.n264 B.n141 256.663
R479 B.n257 B.n141 256.663
R480 B.n255 B.n141 256.663
R481 B.n249 B.n141 256.663
R482 B.n247 B.n141 256.663
R483 B.n240 B.n141 256.663
R484 B.n238 B.n141 256.663
R485 B.n232 B.n141 256.663
R486 B.n230 B.n141 256.663
R487 B.n224 B.n141 256.663
R488 B.n222 B.n141 256.663
R489 B.n216 B.n141 256.663
R490 B.n214 B.n141 256.663
R491 B.n208 B.n141 256.663
R492 B.n206 B.n141 256.663
R493 B.n200 B.n141 256.663
R494 B.n198 B.n141 256.663
R495 B.n192 B.n141 256.663
R496 B.n190 B.n141 256.663
R497 B.n184 B.n141 256.663
R498 B.n182 B.n141 256.663
R499 B.n637 B.n636 256.663
R500 B.n578 B.n576 163.367
R501 B.n574 B.n53 163.367
R502 B.n570 B.n568 163.367
R503 B.n566 B.n55 163.367
R504 B.n562 B.n560 163.367
R505 B.n558 B.n57 163.367
R506 B.n554 B.n552 163.367
R507 B.n550 B.n59 163.367
R508 B.n546 B.n544 163.367
R509 B.n542 B.n61 163.367
R510 B.n538 B.n536 163.367
R511 B.n534 B.n63 163.367
R512 B.n530 B.n528 163.367
R513 B.n526 B.n65 163.367
R514 B.n522 B.n520 163.367
R515 B.n518 B.n67 163.367
R516 B.n514 B.n512 163.367
R517 B.n510 B.n72 163.367
R518 B.n506 B.n504 163.367
R519 B.n502 B.n74 163.367
R520 B.n497 B.n495 163.367
R521 B.n493 B.n78 163.367
R522 B.n489 B.n487 163.367
R523 B.n485 B.n80 163.367
R524 B.n481 B.n479 163.367
R525 B.n477 B.n82 163.367
R526 B.n473 B.n471 163.367
R527 B.n469 B.n84 163.367
R528 B.n465 B.n463 163.367
R529 B.n461 B.n86 163.367
R530 B.n457 B.n455 163.367
R531 B.n453 B.n88 163.367
R532 B.n449 B.n447 163.367
R533 B.n445 B.n90 163.367
R534 B.n441 B.n439 163.367
R535 B.n326 B.n138 163.367
R536 B.n330 B.n138 163.367
R537 B.n330 B.n131 163.367
R538 B.n338 B.n131 163.367
R539 B.n338 B.n129 163.367
R540 B.n342 B.n129 163.367
R541 B.n342 B.n124 163.367
R542 B.n350 B.n124 163.367
R543 B.n350 B.n122 163.367
R544 B.n354 B.n122 163.367
R545 B.n354 B.n115 163.367
R546 B.n362 B.n115 163.367
R547 B.n362 B.n113 163.367
R548 B.n366 B.n113 163.367
R549 B.n366 B.n108 163.367
R550 B.n374 B.n108 163.367
R551 B.n374 B.n106 163.367
R552 B.n378 B.n106 163.367
R553 B.n378 B.n100 163.367
R554 B.n386 B.n100 163.367
R555 B.n386 B.n98 163.367
R556 B.n391 B.n98 163.367
R557 B.n391 B.n92 163.367
R558 B.n399 B.n92 163.367
R559 B.n400 B.n399 163.367
R560 B.n400 B.n5 163.367
R561 B.n6 B.n5 163.367
R562 B.n7 B.n6 163.367
R563 B.n406 B.n7 163.367
R564 B.n408 B.n406 163.367
R565 B.n408 B.n12 163.367
R566 B.n13 B.n12 163.367
R567 B.n14 B.n13 163.367
R568 B.n413 B.n14 163.367
R569 B.n413 B.n19 163.367
R570 B.n20 B.n19 163.367
R571 B.n21 B.n20 163.367
R572 B.n418 B.n21 163.367
R573 B.n418 B.n26 163.367
R574 B.n27 B.n26 163.367
R575 B.n28 B.n27 163.367
R576 B.n423 B.n28 163.367
R577 B.n423 B.n33 163.367
R578 B.n34 B.n33 163.367
R579 B.n35 B.n34 163.367
R580 B.n428 B.n35 163.367
R581 B.n428 B.n40 163.367
R582 B.n41 B.n40 163.367
R583 B.n42 B.n41 163.367
R584 B.n433 B.n42 163.367
R585 B.n433 B.n47 163.367
R586 B.n48 B.n47 163.367
R587 B.n49 B.n48 163.367
R588 B.n320 B.n318 163.367
R589 B.n318 B.n317 163.367
R590 B.n314 B.n313 163.367
R591 B.n311 B.n146 163.367
R592 B.n307 B.n305 163.367
R593 B.n303 B.n148 163.367
R594 B.n299 B.n297 163.367
R595 B.n295 B.n150 163.367
R596 B.n291 B.n289 163.367
R597 B.n287 B.n152 163.367
R598 B.n283 B.n281 163.367
R599 B.n279 B.n154 163.367
R600 B.n275 B.n273 163.367
R601 B.n271 B.n156 163.367
R602 B.n267 B.n265 163.367
R603 B.n263 B.n158 163.367
R604 B.n258 B.n256 163.367
R605 B.n254 B.n162 163.367
R606 B.n250 B.n248 163.367
R607 B.n246 B.n164 163.367
R608 B.n241 B.n239 163.367
R609 B.n237 B.n168 163.367
R610 B.n233 B.n231 163.367
R611 B.n229 B.n170 163.367
R612 B.n225 B.n223 163.367
R613 B.n221 B.n172 163.367
R614 B.n217 B.n215 163.367
R615 B.n213 B.n174 163.367
R616 B.n209 B.n207 163.367
R617 B.n205 B.n176 163.367
R618 B.n201 B.n199 163.367
R619 B.n197 B.n178 163.367
R620 B.n193 B.n191 163.367
R621 B.n189 B.n180 163.367
R622 B.n185 B.n183 163.367
R623 B.n324 B.n136 163.367
R624 B.n332 B.n136 163.367
R625 B.n332 B.n134 163.367
R626 B.n336 B.n134 163.367
R627 B.n336 B.n128 163.367
R628 B.n344 B.n128 163.367
R629 B.n344 B.n126 163.367
R630 B.n348 B.n126 163.367
R631 B.n348 B.n120 163.367
R632 B.n356 B.n120 163.367
R633 B.n356 B.n118 163.367
R634 B.n360 B.n118 163.367
R635 B.n360 B.n112 163.367
R636 B.n368 B.n112 163.367
R637 B.n368 B.n110 163.367
R638 B.n372 B.n110 163.367
R639 B.n372 B.n104 163.367
R640 B.n380 B.n104 163.367
R641 B.n380 B.n102 163.367
R642 B.n384 B.n102 163.367
R643 B.n384 B.n96 163.367
R644 B.n393 B.n96 163.367
R645 B.n393 B.n94 163.367
R646 B.n397 B.n94 163.367
R647 B.n397 B.n3 163.367
R648 B.n635 B.n3 163.367
R649 B.n631 B.n2 163.367
R650 B.n631 B.n630 163.367
R651 B.n630 B.n9 163.367
R652 B.n626 B.n9 163.367
R653 B.n626 B.n11 163.367
R654 B.n622 B.n11 163.367
R655 B.n622 B.n16 163.367
R656 B.n618 B.n16 163.367
R657 B.n618 B.n18 163.367
R658 B.n614 B.n18 163.367
R659 B.n614 B.n23 163.367
R660 B.n610 B.n23 163.367
R661 B.n610 B.n25 163.367
R662 B.n606 B.n25 163.367
R663 B.n606 B.n30 163.367
R664 B.n602 B.n30 163.367
R665 B.n602 B.n32 163.367
R666 B.n598 B.n32 163.367
R667 B.n598 B.n37 163.367
R668 B.n594 B.n37 163.367
R669 B.n594 B.n39 163.367
R670 B.n590 B.n39 163.367
R671 B.n590 B.n44 163.367
R672 B.n586 B.n44 163.367
R673 B.n586 B.n46 163.367
R674 B.n582 B.n46 163.367
R675 B.n75 B.t14 101.299
R676 B.n165 B.t8 101.299
R677 B.n68 B.t17 101.29
R678 B.n159 B.t11 101.29
R679 B.n325 B.n141 98.1207
R680 B.n583 B.n50 98.1207
R681 B.n577 B.n51 71.676
R682 B.n576 B.n575 71.676
R683 B.n569 B.n53 71.676
R684 B.n568 B.n567 71.676
R685 B.n561 B.n55 71.676
R686 B.n560 B.n559 71.676
R687 B.n553 B.n57 71.676
R688 B.n552 B.n551 71.676
R689 B.n545 B.n59 71.676
R690 B.n544 B.n543 71.676
R691 B.n537 B.n61 71.676
R692 B.n536 B.n535 71.676
R693 B.n529 B.n63 71.676
R694 B.n528 B.n527 71.676
R695 B.n521 B.n65 71.676
R696 B.n520 B.n519 71.676
R697 B.n513 B.n67 71.676
R698 B.n512 B.n511 71.676
R699 B.n505 B.n72 71.676
R700 B.n504 B.n503 71.676
R701 B.n496 B.n74 71.676
R702 B.n495 B.n494 71.676
R703 B.n488 B.n78 71.676
R704 B.n487 B.n486 71.676
R705 B.n480 B.n80 71.676
R706 B.n479 B.n478 71.676
R707 B.n472 B.n82 71.676
R708 B.n471 B.n470 71.676
R709 B.n464 B.n84 71.676
R710 B.n463 B.n462 71.676
R711 B.n456 B.n86 71.676
R712 B.n455 B.n454 71.676
R713 B.n448 B.n88 71.676
R714 B.n447 B.n446 71.676
R715 B.n440 B.n90 71.676
R716 B.n441 B.n440 71.676
R717 B.n446 B.n445 71.676
R718 B.n449 B.n448 71.676
R719 B.n454 B.n453 71.676
R720 B.n457 B.n456 71.676
R721 B.n462 B.n461 71.676
R722 B.n465 B.n464 71.676
R723 B.n470 B.n469 71.676
R724 B.n473 B.n472 71.676
R725 B.n478 B.n477 71.676
R726 B.n481 B.n480 71.676
R727 B.n486 B.n485 71.676
R728 B.n489 B.n488 71.676
R729 B.n494 B.n493 71.676
R730 B.n497 B.n496 71.676
R731 B.n503 B.n502 71.676
R732 B.n506 B.n505 71.676
R733 B.n511 B.n510 71.676
R734 B.n514 B.n513 71.676
R735 B.n519 B.n518 71.676
R736 B.n522 B.n521 71.676
R737 B.n527 B.n526 71.676
R738 B.n530 B.n529 71.676
R739 B.n535 B.n534 71.676
R740 B.n538 B.n537 71.676
R741 B.n543 B.n542 71.676
R742 B.n546 B.n545 71.676
R743 B.n551 B.n550 71.676
R744 B.n554 B.n553 71.676
R745 B.n559 B.n558 71.676
R746 B.n562 B.n561 71.676
R747 B.n567 B.n566 71.676
R748 B.n570 B.n569 71.676
R749 B.n575 B.n574 71.676
R750 B.n578 B.n577 71.676
R751 B.n319 B.n142 71.676
R752 B.n317 B.n144 71.676
R753 B.n313 B.n312 71.676
R754 B.n306 B.n146 71.676
R755 B.n305 B.n304 71.676
R756 B.n298 B.n148 71.676
R757 B.n297 B.n296 71.676
R758 B.n290 B.n150 71.676
R759 B.n289 B.n288 71.676
R760 B.n282 B.n152 71.676
R761 B.n281 B.n280 71.676
R762 B.n274 B.n154 71.676
R763 B.n273 B.n272 71.676
R764 B.n266 B.n156 71.676
R765 B.n265 B.n264 71.676
R766 B.n257 B.n158 71.676
R767 B.n256 B.n255 71.676
R768 B.n249 B.n162 71.676
R769 B.n248 B.n247 71.676
R770 B.n240 B.n164 71.676
R771 B.n239 B.n238 71.676
R772 B.n232 B.n168 71.676
R773 B.n231 B.n230 71.676
R774 B.n224 B.n170 71.676
R775 B.n223 B.n222 71.676
R776 B.n216 B.n172 71.676
R777 B.n215 B.n214 71.676
R778 B.n208 B.n174 71.676
R779 B.n207 B.n206 71.676
R780 B.n200 B.n176 71.676
R781 B.n199 B.n198 71.676
R782 B.n192 B.n178 71.676
R783 B.n191 B.n190 71.676
R784 B.n184 B.n180 71.676
R785 B.n183 B.n182 71.676
R786 B.n320 B.n319 71.676
R787 B.n314 B.n144 71.676
R788 B.n312 B.n311 71.676
R789 B.n307 B.n306 71.676
R790 B.n304 B.n303 71.676
R791 B.n299 B.n298 71.676
R792 B.n296 B.n295 71.676
R793 B.n291 B.n290 71.676
R794 B.n288 B.n287 71.676
R795 B.n283 B.n282 71.676
R796 B.n280 B.n279 71.676
R797 B.n275 B.n274 71.676
R798 B.n272 B.n271 71.676
R799 B.n267 B.n266 71.676
R800 B.n264 B.n263 71.676
R801 B.n258 B.n257 71.676
R802 B.n255 B.n254 71.676
R803 B.n250 B.n249 71.676
R804 B.n247 B.n246 71.676
R805 B.n241 B.n240 71.676
R806 B.n238 B.n237 71.676
R807 B.n233 B.n232 71.676
R808 B.n230 B.n229 71.676
R809 B.n225 B.n224 71.676
R810 B.n222 B.n221 71.676
R811 B.n217 B.n216 71.676
R812 B.n214 B.n213 71.676
R813 B.n209 B.n208 71.676
R814 B.n206 B.n205 71.676
R815 B.n201 B.n200 71.676
R816 B.n198 B.n197 71.676
R817 B.n193 B.n192 71.676
R818 B.n190 B.n189 71.676
R819 B.n185 B.n184 71.676
R820 B.n182 B.n140 71.676
R821 B.n636 B.n635 71.676
R822 B.n636 B.n2 71.676
R823 B.n76 B.t15 71.0445
R824 B.n166 B.t7 71.0445
R825 B.n69 B.t18 71.0348
R826 B.n160 B.t10 71.0348
R827 B.n70 B.n69 59.5399
R828 B.n500 B.n76 59.5399
R829 B.n243 B.n166 59.5399
R830 B.n261 B.n160 59.5399
R831 B.n325 B.n137 55.1424
R832 B.n331 B.n137 55.1424
R833 B.n331 B.n132 55.1424
R834 B.n337 B.n132 55.1424
R835 B.n337 B.n133 55.1424
R836 B.n343 B.n125 55.1424
R837 B.n349 B.n125 55.1424
R838 B.n349 B.n121 55.1424
R839 B.n355 B.n121 55.1424
R840 B.n355 B.n116 55.1424
R841 B.n361 B.n116 55.1424
R842 B.n361 B.n117 55.1424
R843 B.n367 B.n109 55.1424
R844 B.n373 B.n109 55.1424
R845 B.n373 B.n105 55.1424
R846 B.n379 B.n105 55.1424
R847 B.n385 B.n101 55.1424
R848 B.n385 B.n97 55.1424
R849 B.n392 B.n97 55.1424
R850 B.n398 B.n93 55.1424
R851 B.n398 B.n4 55.1424
R852 B.n634 B.n4 55.1424
R853 B.n634 B.n633 55.1424
R854 B.n633 B.n632 55.1424
R855 B.n632 B.n8 55.1424
R856 B.n407 B.n8 55.1424
R857 B.n625 B.n624 55.1424
R858 B.n624 B.n623 55.1424
R859 B.n623 B.n15 55.1424
R860 B.n617 B.n616 55.1424
R861 B.n616 B.n615 55.1424
R862 B.n615 B.n22 55.1424
R863 B.n609 B.n22 55.1424
R864 B.n608 B.n607 55.1424
R865 B.n607 B.n29 55.1424
R866 B.n601 B.n29 55.1424
R867 B.n601 B.n600 55.1424
R868 B.n600 B.n599 55.1424
R869 B.n599 B.n36 55.1424
R870 B.n593 B.n36 55.1424
R871 B.n592 B.n591 55.1424
R872 B.n591 B.n43 55.1424
R873 B.n585 B.n43 55.1424
R874 B.n585 B.n584 55.1424
R875 B.n584 B.n583 55.1424
R876 B.t19 B.n101 54.3315
R877 B.t2 B.n15 54.3315
R878 B.n133 B.t6 34.8696
R879 B.t13 B.n592 34.8696
R880 B.n392 B.t3 33.2478
R881 B.n625 B.t1 33.2478
R882 B.n323 B.n322 32.0005
R883 B.n327 B.n139 32.0005
R884 B.n438 B.n437 32.0005
R885 B.n581 B.n580 32.0005
R886 B.n367 B.t0 31.626
R887 B.n609 B.t4 31.626
R888 B.n69 B.n68 30.255
R889 B.n76 B.n75 30.255
R890 B.n166 B.n165 30.255
R891 B.n160 B.n159 30.255
R892 B.n117 B.t0 23.5169
R893 B.t4 B.n608 23.5169
R894 B.t3 B.n93 21.8951
R895 B.n407 B.t1 21.8951
R896 B.n343 B.t6 20.2733
R897 B.n593 B.t13 20.2733
R898 B B.n637 18.0485
R899 B.n323 B.n135 10.6151
R900 B.n333 B.n135 10.6151
R901 B.n334 B.n333 10.6151
R902 B.n335 B.n334 10.6151
R903 B.n335 B.n127 10.6151
R904 B.n345 B.n127 10.6151
R905 B.n346 B.n345 10.6151
R906 B.n347 B.n346 10.6151
R907 B.n347 B.n119 10.6151
R908 B.n357 B.n119 10.6151
R909 B.n358 B.n357 10.6151
R910 B.n359 B.n358 10.6151
R911 B.n359 B.n111 10.6151
R912 B.n369 B.n111 10.6151
R913 B.n370 B.n369 10.6151
R914 B.n371 B.n370 10.6151
R915 B.n371 B.n103 10.6151
R916 B.n381 B.n103 10.6151
R917 B.n382 B.n381 10.6151
R918 B.n383 B.n382 10.6151
R919 B.n383 B.n95 10.6151
R920 B.n394 B.n95 10.6151
R921 B.n395 B.n394 10.6151
R922 B.n396 B.n395 10.6151
R923 B.n396 B.n0 10.6151
R924 B.n322 B.n321 10.6151
R925 B.n321 B.n143 10.6151
R926 B.n316 B.n143 10.6151
R927 B.n316 B.n315 10.6151
R928 B.n315 B.n145 10.6151
R929 B.n310 B.n145 10.6151
R930 B.n310 B.n309 10.6151
R931 B.n309 B.n308 10.6151
R932 B.n308 B.n147 10.6151
R933 B.n302 B.n147 10.6151
R934 B.n302 B.n301 10.6151
R935 B.n301 B.n300 10.6151
R936 B.n300 B.n149 10.6151
R937 B.n294 B.n149 10.6151
R938 B.n294 B.n293 10.6151
R939 B.n293 B.n292 10.6151
R940 B.n292 B.n151 10.6151
R941 B.n286 B.n151 10.6151
R942 B.n286 B.n285 10.6151
R943 B.n285 B.n284 10.6151
R944 B.n284 B.n153 10.6151
R945 B.n278 B.n153 10.6151
R946 B.n278 B.n277 10.6151
R947 B.n277 B.n276 10.6151
R948 B.n276 B.n155 10.6151
R949 B.n270 B.n155 10.6151
R950 B.n270 B.n269 10.6151
R951 B.n269 B.n268 10.6151
R952 B.n268 B.n157 10.6151
R953 B.n262 B.n157 10.6151
R954 B.n260 B.n259 10.6151
R955 B.n259 B.n161 10.6151
R956 B.n253 B.n161 10.6151
R957 B.n253 B.n252 10.6151
R958 B.n252 B.n251 10.6151
R959 B.n251 B.n163 10.6151
R960 B.n245 B.n163 10.6151
R961 B.n245 B.n244 10.6151
R962 B.n242 B.n167 10.6151
R963 B.n236 B.n167 10.6151
R964 B.n236 B.n235 10.6151
R965 B.n235 B.n234 10.6151
R966 B.n234 B.n169 10.6151
R967 B.n228 B.n169 10.6151
R968 B.n228 B.n227 10.6151
R969 B.n227 B.n226 10.6151
R970 B.n226 B.n171 10.6151
R971 B.n220 B.n171 10.6151
R972 B.n220 B.n219 10.6151
R973 B.n219 B.n218 10.6151
R974 B.n218 B.n173 10.6151
R975 B.n212 B.n173 10.6151
R976 B.n212 B.n211 10.6151
R977 B.n211 B.n210 10.6151
R978 B.n210 B.n175 10.6151
R979 B.n204 B.n175 10.6151
R980 B.n204 B.n203 10.6151
R981 B.n203 B.n202 10.6151
R982 B.n202 B.n177 10.6151
R983 B.n196 B.n177 10.6151
R984 B.n196 B.n195 10.6151
R985 B.n195 B.n194 10.6151
R986 B.n194 B.n179 10.6151
R987 B.n188 B.n179 10.6151
R988 B.n188 B.n187 10.6151
R989 B.n187 B.n186 10.6151
R990 B.n186 B.n181 10.6151
R991 B.n181 B.n139 10.6151
R992 B.n328 B.n327 10.6151
R993 B.n329 B.n328 10.6151
R994 B.n329 B.n130 10.6151
R995 B.n339 B.n130 10.6151
R996 B.n340 B.n339 10.6151
R997 B.n341 B.n340 10.6151
R998 B.n341 B.n123 10.6151
R999 B.n351 B.n123 10.6151
R1000 B.n352 B.n351 10.6151
R1001 B.n353 B.n352 10.6151
R1002 B.n353 B.n114 10.6151
R1003 B.n363 B.n114 10.6151
R1004 B.n364 B.n363 10.6151
R1005 B.n365 B.n364 10.6151
R1006 B.n365 B.n107 10.6151
R1007 B.n375 B.n107 10.6151
R1008 B.n376 B.n375 10.6151
R1009 B.n377 B.n376 10.6151
R1010 B.n377 B.n99 10.6151
R1011 B.n387 B.n99 10.6151
R1012 B.n388 B.n387 10.6151
R1013 B.n390 B.n388 10.6151
R1014 B.n390 B.n389 10.6151
R1015 B.n389 B.n91 10.6151
R1016 B.n401 B.n91 10.6151
R1017 B.n402 B.n401 10.6151
R1018 B.n403 B.n402 10.6151
R1019 B.n404 B.n403 10.6151
R1020 B.n405 B.n404 10.6151
R1021 B.n409 B.n405 10.6151
R1022 B.n410 B.n409 10.6151
R1023 B.n411 B.n410 10.6151
R1024 B.n412 B.n411 10.6151
R1025 B.n414 B.n412 10.6151
R1026 B.n415 B.n414 10.6151
R1027 B.n416 B.n415 10.6151
R1028 B.n417 B.n416 10.6151
R1029 B.n419 B.n417 10.6151
R1030 B.n420 B.n419 10.6151
R1031 B.n421 B.n420 10.6151
R1032 B.n422 B.n421 10.6151
R1033 B.n424 B.n422 10.6151
R1034 B.n425 B.n424 10.6151
R1035 B.n426 B.n425 10.6151
R1036 B.n427 B.n426 10.6151
R1037 B.n429 B.n427 10.6151
R1038 B.n430 B.n429 10.6151
R1039 B.n431 B.n430 10.6151
R1040 B.n432 B.n431 10.6151
R1041 B.n434 B.n432 10.6151
R1042 B.n435 B.n434 10.6151
R1043 B.n436 B.n435 10.6151
R1044 B.n437 B.n436 10.6151
R1045 B.n629 B.n1 10.6151
R1046 B.n629 B.n628 10.6151
R1047 B.n628 B.n627 10.6151
R1048 B.n627 B.n10 10.6151
R1049 B.n621 B.n10 10.6151
R1050 B.n621 B.n620 10.6151
R1051 B.n620 B.n619 10.6151
R1052 B.n619 B.n17 10.6151
R1053 B.n613 B.n17 10.6151
R1054 B.n613 B.n612 10.6151
R1055 B.n612 B.n611 10.6151
R1056 B.n611 B.n24 10.6151
R1057 B.n605 B.n24 10.6151
R1058 B.n605 B.n604 10.6151
R1059 B.n604 B.n603 10.6151
R1060 B.n603 B.n31 10.6151
R1061 B.n597 B.n31 10.6151
R1062 B.n597 B.n596 10.6151
R1063 B.n596 B.n595 10.6151
R1064 B.n595 B.n38 10.6151
R1065 B.n589 B.n38 10.6151
R1066 B.n589 B.n588 10.6151
R1067 B.n588 B.n587 10.6151
R1068 B.n587 B.n45 10.6151
R1069 B.n581 B.n45 10.6151
R1070 B.n580 B.n579 10.6151
R1071 B.n579 B.n52 10.6151
R1072 B.n573 B.n52 10.6151
R1073 B.n573 B.n572 10.6151
R1074 B.n572 B.n571 10.6151
R1075 B.n571 B.n54 10.6151
R1076 B.n565 B.n54 10.6151
R1077 B.n565 B.n564 10.6151
R1078 B.n564 B.n563 10.6151
R1079 B.n563 B.n56 10.6151
R1080 B.n557 B.n56 10.6151
R1081 B.n557 B.n556 10.6151
R1082 B.n556 B.n555 10.6151
R1083 B.n555 B.n58 10.6151
R1084 B.n549 B.n58 10.6151
R1085 B.n549 B.n548 10.6151
R1086 B.n548 B.n547 10.6151
R1087 B.n547 B.n60 10.6151
R1088 B.n541 B.n60 10.6151
R1089 B.n541 B.n540 10.6151
R1090 B.n540 B.n539 10.6151
R1091 B.n539 B.n62 10.6151
R1092 B.n533 B.n62 10.6151
R1093 B.n533 B.n532 10.6151
R1094 B.n532 B.n531 10.6151
R1095 B.n531 B.n64 10.6151
R1096 B.n525 B.n64 10.6151
R1097 B.n525 B.n524 10.6151
R1098 B.n524 B.n523 10.6151
R1099 B.n523 B.n66 10.6151
R1100 B.n517 B.n516 10.6151
R1101 B.n516 B.n515 10.6151
R1102 B.n515 B.n71 10.6151
R1103 B.n509 B.n71 10.6151
R1104 B.n509 B.n508 10.6151
R1105 B.n508 B.n507 10.6151
R1106 B.n507 B.n73 10.6151
R1107 B.n501 B.n73 10.6151
R1108 B.n499 B.n498 10.6151
R1109 B.n498 B.n77 10.6151
R1110 B.n492 B.n77 10.6151
R1111 B.n492 B.n491 10.6151
R1112 B.n491 B.n490 10.6151
R1113 B.n490 B.n79 10.6151
R1114 B.n484 B.n79 10.6151
R1115 B.n484 B.n483 10.6151
R1116 B.n483 B.n482 10.6151
R1117 B.n482 B.n81 10.6151
R1118 B.n476 B.n81 10.6151
R1119 B.n476 B.n475 10.6151
R1120 B.n475 B.n474 10.6151
R1121 B.n474 B.n83 10.6151
R1122 B.n468 B.n83 10.6151
R1123 B.n468 B.n467 10.6151
R1124 B.n467 B.n466 10.6151
R1125 B.n466 B.n85 10.6151
R1126 B.n460 B.n85 10.6151
R1127 B.n460 B.n459 10.6151
R1128 B.n459 B.n458 10.6151
R1129 B.n458 B.n87 10.6151
R1130 B.n452 B.n87 10.6151
R1131 B.n452 B.n451 10.6151
R1132 B.n451 B.n450 10.6151
R1133 B.n450 B.n89 10.6151
R1134 B.n444 B.n89 10.6151
R1135 B.n444 B.n443 10.6151
R1136 B.n443 B.n442 10.6151
R1137 B.n442 B.n438 10.6151
R1138 B.n637 B.n0 8.11757
R1139 B.n637 B.n1 8.11757
R1140 B.n261 B.n260 6.5566
R1141 B.n244 B.n243 6.5566
R1142 B.n517 B.n70 6.5566
R1143 B.n501 B.n500 6.5566
R1144 B.n262 B.n261 4.05904
R1145 B.n243 B.n242 4.05904
R1146 B.n70 B.n66 4.05904
R1147 B.n500 B.n499 4.05904
R1148 B.n379 B.t19 0.81141
R1149 B.n617 B.t2 0.81141
R1150 VP.n5 VP.t5 213.067
R1151 VP.n12 VP.t1 194.564
R1152 VP.n19 VP.t4 194.564
R1153 VP.n9 VP.t3 194.564
R1154 VP.n1 VP.t2 162.43
R1155 VP.n4 VP.t0 162.43
R1156 VP.n7 VP.n6 161.3
R1157 VP.n8 VP.n3 161.3
R1158 VP.n18 VP.n0 161.3
R1159 VP.n17 VP.n16 161.3
R1160 VP.n15 VP.n14 161.3
R1161 VP.n13 VP.n2 161.3
R1162 VP.n10 VP.n9 80.6037
R1163 VP.n20 VP.n19 80.6037
R1164 VP.n12 VP.n11 80.6037
R1165 VP.n5 VP.n4 45.5344
R1166 VP.n11 VP.n10 40.6226
R1167 VP.n14 VP.n13 37.5796
R1168 VP.n18 VP.n17 37.5796
R1169 VP.n8 VP.n7 37.5796
R1170 VP.n6 VP.n5 29.7304
R1171 VP.n13 VP.n12 28.4823
R1172 VP.n19 VP.n18 28.4823
R1173 VP.n9 VP.n8 28.4823
R1174 VP.n14 VP.n1 12.234
R1175 VP.n17 VP.n1 12.234
R1176 VP.n7 VP.n4 12.234
R1177 VP.n10 VP.n3 0.285035
R1178 VP.n11 VP.n2 0.285035
R1179 VP.n20 VP.n0 0.285035
R1180 VP.n6 VP.n3 0.189894
R1181 VP.n15 VP.n2 0.189894
R1182 VP.n16 VP.n15 0.189894
R1183 VP.n16 VP.n0 0.189894
R1184 VP VP.n20 0.146778
R1185 VDD1 VDD1.t0 69.6721
R1186 VDD1.n1 VDD1.t4 69.5585
R1187 VDD1.n1 VDD1.n0 66.4975
R1188 VDD1.n3 VDD1.n2 66.2168
R1189 VDD1.n3 VDD1.n1 36.488
R1190 VDD1.n2 VDD1.t5 2.38892
R1191 VDD1.n2 VDD1.t2 2.38892
R1192 VDD1.n0 VDD1.t3 2.38892
R1193 VDD1.n0 VDD1.t1 2.38892
R1194 VDD1 VDD1.n3 0.278517
C0 VDD1 VN 0.148682f
C1 VDD1 VTAIL 6.45892f
C2 VDD2 VDD1 0.903748f
C3 VDD1 VP 4.10562f
C4 VN VTAIL 3.90232f
C5 VDD2 VN 3.91548f
C6 VP VN 4.90888f
C7 VDD2 VTAIL 6.4998f
C8 VP VTAIL 3.91668f
C9 VDD2 VP 0.341715f
C10 VDD2 B 4.233115f
C11 VDD1 B 4.488052f
C12 VTAIL B 5.40869f
C13 VN B 8.698421f
C14 VP B 7.131883f
C15 VDD1.t0 B 1.6235f
C16 VDD1.t4 B 1.62288f
C17 VDD1.t3 B 0.146424f
C18 VDD1.t1 B 0.146424f
C19 VDD1.n0 B 1.27371f
C20 VDD1.n1 B 1.92981f
C21 VDD1.t5 B 0.146424f
C22 VDD1.t2 B 0.146424f
C23 VDD1.n2 B 1.27241f
C24 VDD1.n3 B 1.88336f
C25 VP.n0 B 0.050095f
C26 VP.t2 B 1.02966f
C27 VP.n1 B 0.392142f
C28 VP.n2 B 0.050095f
C29 VP.n3 B 0.050095f
C30 VP.t3 B 1.1004f
C31 VP.t0 B 1.02966f
C32 VP.n4 B 0.439737f
C33 VP.t5 B 1.14137f
C34 VP.n5 B 0.456472f
C35 VP.n6 B 0.194087f
C36 VP.n7 B 0.058238f
C37 VP.n8 B 0.021989f
C38 VP.n9 B 0.463086f
C39 VP.n10 B 1.47826f
C40 VP.n11 B 1.51148f
C41 VP.t1 B 1.1004f
C42 VP.n12 B 0.463086f
C43 VP.n13 B 0.021989f
C44 VP.n14 B 0.058238f
C45 VP.n15 B 0.037542f
C46 VP.n16 B 0.037542f
C47 VP.n17 B 0.058238f
C48 VP.n18 B 0.021989f
C49 VP.t4 B 1.1004f
C50 VP.n19 B 0.463086f
C51 VP.n20 B 0.035159f
C52 VDD2.t0 B 1.60476f
C53 VDD2.t2 B 0.144788f
C54 VDD2.t3 B 0.144788f
C55 VDD2.n0 B 1.25948f
C56 VDD2.n1 B 1.83078f
C57 VDD2.t5 B 1.60058f
C58 VDD2.n2 B 1.87108f
C59 VDD2.t1 B 0.144788f
C60 VDD2.t4 B 0.144788f
C61 VDD2.n3 B 1.25946f
C62 VTAIL.t7 B 0.159582f
C63 VTAIL.t8 B 0.159582f
C64 VTAIL.n0 B 1.32311f
C65 VTAIL.n1 B 0.344822f
C66 VTAIL.t3 B 1.6848f
C67 VTAIL.n2 B 0.492965f
C68 VTAIL.t0 B 0.159582f
C69 VTAIL.t11 B 0.159582f
C70 VTAIL.n3 B 1.32311f
C71 VTAIL.n4 B 1.43274f
C72 VTAIL.t10 B 0.159582f
C73 VTAIL.t5 B 0.159582f
C74 VTAIL.n5 B 1.32312f
C75 VTAIL.n6 B 1.43274f
C76 VTAIL.t6 B 1.68481f
C77 VTAIL.n7 B 0.492953f
C78 VTAIL.t1 B 0.159582f
C79 VTAIL.t2 B 0.159582f
C80 VTAIL.n8 B 1.32312f
C81 VTAIL.n9 B 0.41942f
C82 VTAIL.t4 B 1.6848f
C83 VTAIL.n10 B 1.40072f
C84 VTAIL.t9 B 1.6848f
C85 VTAIL.n11 B 1.36976f
C86 VN.n0 B 0.049117f
C87 VN.t3 B 1.00956f
C88 VN.n1 B 0.431155f
C89 VN.t5 B 1.1191f
C90 VN.n2 B 0.447564f
C91 VN.n3 B 0.190299f
C92 VN.n4 B 0.057102f
C93 VN.n5 B 0.02156f
C94 VN.t2 B 1.07893f
C95 VN.n6 B 0.454049f
C96 VN.n7 B 0.034473f
C97 VN.n8 B 0.049117f
C98 VN.t4 B 1.00956f
C99 VN.n9 B 0.431155f
C100 VN.t1 B 1.1191f
C101 VN.n10 B 0.447564f
C102 VN.n11 B 0.190299f
C103 VN.n12 B 0.057102f
C104 VN.n13 B 0.02156f
C105 VN.t0 B 1.07893f
C106 VN.n14 B 0.454049f
C107 VN.n15 B 1.47019f
.ends

