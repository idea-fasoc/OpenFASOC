* NGSPICE file created from diff_pair_sample_0979.ext - technology: sky130A

.subckt diff_pair_sample_0979 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t19 VN.t0 VDD2.t5 w_n3802_n1648# sky130_fd_pr__pfet_01v8 ad=0.561 pd=3.73 as=0.561 ps=3.73 w=3.4 l=2.03
X1 VDD1.t9 VP.t0 VTAIL.t1 w_n3802_n1648# sky130_fd_pr__pfet_01v8 ad=0.561 pd=3.73 as=1.326 ps=7.58 w=3.4 l=2.03
X2 VDD1.t8 VP.t1 VTAIL.t6 w_n3802_n1648# sky130_fd_pr__pfet_01v8 ad=0.561 pd=3.73 as=0.561 ps=3.73 w=3.4 l=2.03
X3 VTAIL.t18 VN.t1 VDD2.t8 w_n3802_n1648# sky130_fd_pr__pfet_01v8 ad=0.561 pd=3.73 as=0.561 ps=3.73 w=3.4 l=2.03
X4 B.t11 B.t9 B.t10 w_n3802_n1648# sky130_fd_pr__pfet_01v8 ad=1.326 pd=7.58 as=0 ps=0 w=3.4 l=2.03
X5 VTAIL.t17 VN.t2 VDD2.t0 w_n3802_n1648# sky130_fd_pr__pfet_01v8 ad=0.561 pd=3.73 as=0.561 ps=3.73 w=3.4 l=2.03
X6 VTAIL.t7 VP.t2 VDD1.t7 w_n3802_n1648# sky130_fd_pr__pfet_01v8 ad=0.561 pd=3.73 as=0.561 ps=3.73 w=3.4 l=2.03
X7 VDD1.t6 VP.t3 VTAIL.t0 w_n3802_n1648# sky130_fd_pr__pfet_01v8 ad=1.326 pd=7.58 as=0.561 ps=3.73 w=3.4 l=2.03
X8 VTAIL.t16 VN.t3 VDD2.t2 w_n3802_n1648# sky130_fd_pr__pfet_01v8 ad=0.561 pd=3.73 as=0.561 ps=3.73 w=3.4 l=2.03
X9 VDD1.t5 VP.t4 VTAIL.t2 w_n3802_n1648# sky130_fd_pr__pfet_01v8 ad=0.561 pd=3.73 as=0.561 ps=3.73 w=3.4 l=2.03
X10 VDD1.t4 VP.t5 VTAIL.t5 w_n3802_n1648# sky130_fd_pr__pfet_01v8 ad=1.326 pd=7.58 as=0.561 ps=3.73 w=3.4 l=2.03
X11 VDD2.t7 VN.t4 VTAIL.t15 w_n3802_n1648# sky130_fd_pr__pfet_01v8 ad=0.561 pd=3.73 as=0.561 ps=3.73 w=3.4 l=2.03
X12 VDD2.t9 VN.t5 VTAIL.t14 w_n3802_n1648# sky130_fd_pr__pfet_01v8 ad=0.561 pd=3.73 as=1.326 ps=7.58 w=3.4 l=2.03
X13 VDD2.t6 VN.t6 VTAIL.t13 w_n3802_n1648# sky130_fd_pr__pfet_01v8 ad=1.326 pd=7.58 as=0.561 ps=3.73 w=3.4 l=2.03
X14 VDD1.t3 VP.t6 VTAIL.t3 w_n3802_n1648# sky130_fd_pr__pfet_01v8 ad=0.561 pd=3.73 as=1.326 ps=7.58 w=3.4 l=2.03
X15 VDD2.t4 VN.t7 VTAIL.t12 w_n3802_n1648# sky130_fd_pr__pfet_01v8 ad=0.561 pd=3.73 as=0.561 ps=3.73 w=3.4 l=2.03
X16 VDD2.t3 VN.t8 VTAIL.t11 w_n3802_n1648# sky130_fd_pr__pfet_01v8 ad=0.561 pd=3.73 as=1.326 ps=7.58 w=3.4 l=2.03
X17 VDD2.t1 VN.t9 VTAIL.t10 w_n3802_n1648# sky130_fd_pr__pfet_01v8 ad=1.326 pd=7.58 as=0.561 ps=3.73 w=3.4 l=2.03
X18 B.t8 B.t6 B.t7 w_n3802_n1648# sky130_fd_pr__pfet_01v8 ad=1.326 pd=7.58 as=0 ps=0 w=3.4 l=2.03
X19 VTAIL.t9 VP.t7 VDD1.t2 w_n3802_n1648# sky130_fd_pr__pfet_01v8 ad=0.561 pd=3.73 as=0.561 ps=3.73 w=3.4 l=2.03
X20 VTAIL.t8 VP.t8 VDD1.t1 w_n3802_n1648# sky130_fd_pr__pfet_01v8 ad=0.561 pd=3.73 as=0.561 ps=3.73 w=3.4 l=2.03
X21 B.t5 B.t3 B.t4 w_n3802_n1648# sky130_fd_pr__pfet_01v8 ad=1.326 pd=7.58 as=0 ps=0 w=3.4 l=2.03
X22 B.t2 B.t0 B.t1 w_n3802_n1648# sky130_fd_pr__pfet_01v8 ad=1.326 pd=7.58 as=0 ps=0 w=3.4 l=2.03
X23 VTAIL.t4 VP.t9 VDD1.t0 w_n3802_n1648# sky130_fd_pr__pfet_01v8 ad=0.561 pd=3.73 as=0.561 ps=3.73 w=3.4 l=2.03
R0 VN.n65 VN.n34 161.3
R1 VN.n64 VN.n63 161.3
R2 VN.n62 VN.n35 161.3
R3 VN.n61 VN.n60 161.3
R4 VN.n58 VN.n36 161.3
R5 VN.n57 VN.n56 161.3
R6 VN.n55 VN.n37 161.3
R7 VN.n54 VN.n53 161.3
R8 VN.n52 VN.n38 161.3
R9 VN.n50 VN.n49 161.3
R10 VN.n48 VN.n39 161.3
R11 VN.n47 VN.n46 161.3
R12 VN.n45 VN.n40 161.3
R13 VN.n44 VN.n43 161.3
R14 VN.n31 VN.n0 161.3
R15 VN.n30 VN.n29 161.3
R16 VN.n28 VN.n1 161.3
R17 VN.n27 VN.n26 161.3
R18 VN.n24 VN.n2 161.3
R19 VN.n23 VN.n22 161.3
R20 VN.n21 VN.n3 161.3
R21 VN.n20 VN.n19 161.3
R22 VN.n18 VN.n4 161.3
R23 VN.n16 VN.n15 161.3
R24 VN.n14 VN.n5 161.3
R25 VN.n13 VN.n12 161.3
R26 VN.n11 VN.n6 161.3
R27 VN.n10 VN.n9 161.3
R28 VN.n33 VN.n32 87.7919
R29 VN.n67 VN.n66 87.7919
R30 VN.n8 VN.t9 71.3343
R31 VN.n42 VN.t5 71.3343
R32 VN.n8 VN.n7 65.0363
R33 VN.n42 VN.n41 65.0363
R34 VN.n30 VN.n1 56.5617
R35 VN.n64 VN.n35 56.5617
R36 VN.n12 VN.n5 47.3584
R37 VN.n19 VN.n3 47.3584
R38 VN.n46 VN.n39 47.3584
R39 VN.n53 VN.n37 47.3584
R40 VN VN.n67 43.8618
R41 VN.n7 VN.t3 40.365
R42 VN.n17 VN.t4 40.365
R43 VN.n25 VN.t0 40.365
R44 VN.n32 VN.t8 40.365
R45 VN.n41 VN.t1 40.365
R46 VN.n51 VN.t7 40.365
R47 VN.n59 VN.t2 40.365
R48 VN.n66 VN.t6 40.365
R49 VN.n12 VN.n11 33.7956
R50 VN.n23 VN.n3 33.7956
R51 VN.n46 VN.n45 33.7956
R52 VN.n57 VN.n37 33.7956
R53 VN.n11 VN.n10 24.5923
R54 VN.n16 VN.n5 24.5923
R55 VN.n19 VN.n18 24.5923
R56 VN.n24 VN.n23 24.5923
R57 VN.n26 VN.n1 24.5923
R58 VN.n31 VN.n30 24.5923
R59 VN.n45 VN.n44 24.5923
R60 VN.n53 VN.n52 24.5923
R61 VN.n50 VN.n39 24.5923
R62 VN.n60 VN.n35 24.5923
R63 VN.n58 VN.n57 24.5923
R64 VN.n65 VN.n64 24.5923
R65 VN.n32 VN.n31 23.1168
R66 VN.n66 VN.n65 23.1168
R67 VN.n26 VN.n25 19.1821
R68 VN.n60 VN.n59 19.1821
R69 VN.n43 VN.n42 12.856
R70 VN.n9 VN.n8 12.856
R71 VN.n17 VN.n16 12.2964
R72 VN.n18 VN.n17 12.2964
R73 VN.n52 VN.n51 12.2964
R74 VN.n51 VN.n50 12.2964
R75 VN.n10 VN.n7 5.4107
R76 VN.n25 VN.n24 5.4107
R77 VN.n44 VN.n41 5.4107
R78 VN.n59 VN.n58 5.4107
R79 VN.n67 VN.n34 0.278335
R80 VN.n33 VN.n0 0.278335
R81 VN.n63 VN.n34 0.189894
R82 VN.n63 VN.n62 0.189894
R83 VN.n62 VN.n61 0.189894
R84 VN.n61 VN.n36 0.189894
R85 VN.n56 VN.n36 0.189894
R86 VN.n56 VN.n55 0.189894
R87 VN.n55 VN.n54 0.189894
R88 VN.n54 VN.n38 0.189894
R89 VN.n49 VN.n38 0.189894
R90 VN.n49 VN.n48 0.189894
R91 VN.n48 VN.n47 0.189894
R92 VN.n47 VN.n40 0.189894
R93 VN.n43 VN.n40 0.189894
R94 VN.n9 VN.n6 0.189894
R95 VN.n13 VN.n6 0.189894
R96 VN.n14 VN.n13 0.189894
R97 VN.n15 VN.n14 0.189894
R98 VN.n15 VN.n4 0.189894
R99 VN.n20 VN.n4 0.189894
R100 VN.n21 VN.n20 0.189894
R101 VN.n22 VN.n21 0.189894
R102 VN.n22 VN.n2 0.189894
R103 VN.n27 VN.n2 0.189894
R104 VN.n28 VN.n27 0.189894
R105 VN.n29 VN.n28 0.189894
R106 VN.n29 VN.n0 0.189894
R107 VN VN.n33 0.153485
R108 VDD2.n29 VDD2.n19 756.745
R109 VDD2.n10 VDD2.n0 756.745
R110 VDD2.n30 VDD2.n29 585
R111 VDD2.n28 VDD2.n27 585
R112 VDD2.n23 VDD2.n22 585
R113 VDD2.n4 VDD2.n3 585
R114 VDD2.n9 VDD2.n8 585
R115 VDD2.n11 VDD2.n10 585
R116 VDD2.n24 VDD2.t6 338.558
R117 VDD2.n5 VDD2.t1 338.558
R118 VDD2.n29 VDD2.n28 171.744
R119 VDD2.n28 VDD2.n22 171.744
R120 VDD2.n9 VDD2.n3 171.744
R121 VDD2.n10 VDD2.n9 171.744
R122 VDD2.n18 VDD2.n17 128.837
R123 VDD2 VDD2.n37 128.833
R124 VDD2.n36 VDD2.n35 127.367
R125 VDD2.n16 VDD2.n15 127.367
R126 VDD2.t6 VDD2.n22 85.8723
R127 VDD2.t1 VDD2.n3 85.8723
R128 VDD2.n16 VDD2.n14 49.3471
R129 VDD2.n34 VDD2.n33 47.3126
R130 VDD2.n34 VDD2.n18 36.3101
R131 VDD2.n24 VDD2.n23 10.6058
R132 VDD2.n5 VDD2.n4 10.6058
R133 VDD2.n33 VDD2.n19 9.69747
R134 VDD2.n14 VDD2.n0 9.69747
R135 VDD2.n37 VDD2.t8 9.56079
R136 VDD2.n37 VDD2.t9 9.56079
R137 VDD2.n35 VDD2.t0 9.56079
R138 VDD2.n35 VDD2.t4 9.56079
R139 VDD2.n17 VDD2.t5 9.56079
R140 VDD2.n17 VDD2.t3 9.56079
R141 VDD2.n15 VDD2.t2 9.56079
R142 VDD2.n15 VDD2.t7 9.56079
R143 VDD2.n33 VDD2.n32 9.45567
R144 VDD2.n14 VDD2.n13 9.45567
R145 VDD2.n21 VDD2.n20 9.3005
R146 VDD2.n32 VDD2.n31 9.3005
R147 VDD2.n26 VDD2.n25 9.3005
R148 VDD2.n7 VDD2.n6 9.3005
R149 VDD2.n2 VDD2.n1 9.3005
R150 VDD2.n13 VDD2.n12 9.3005
R151 VDD2.n31 VDD2.n30 8.92171
R152 VDD2.n12 VDD2.n11 8.92171
R153 VDD2.n27 VDD2.n21 8.14595
R154 VDD2.n8 VDD2.n2 8.14595
R155 VDD2.n26 VDD2.n23 7.3702
R156 VDD2.n7 VDD2.n4 7.3702
R157 VDD2.n27 VDD2.n26 5.81868
R158 VDD2.n8 VDD2.n7 5.81868
R159 VDD2.n30 VDD2.n21 5.04292
R160 VDD2.n11 VDD2.n2 5.04292
R161 VDD2.n31 VDD2.n19 4.26717
R162 VDD2.n12 VDD2.n0 4.26717
R163 VDD2.n25 VDD2.n24 2.5326
R164 VDD2.n6 VDD2.n5 2.5326
R165 VDD2.n36 VDD2.n34 2.03498
R166 VDD2 VDD2.n36 0.56731
R167 VDD2.n18 VDD2.n16 0.453775
R168 VDD2.n32 VDD2.n20 0.155672
R169 VDD2.n25 VDD2.n20 0.155672
R170 VDD2.n6 VDD2.n1 0.155672
R171 VDD2.n13 VDD2.n1 0.155672
R172 VTAIL.n72 VTAIL.n62 756.745
R173 VTAIL.n12 VTAIL.n2 756.745
R174 VTAIL.n56 VTAIL.n46 756.745
R175 VTAIL.n36 VTAIL.n26 756.745
R176 VTAIL.n66 VTAIL.n65 585
R177 VTAIL.n71 VTAIL.n70 585
R178 VTAIL.n73 VTAIL.n72 585
R179 VTAIL.n6 VTAIL.n5 585
R180 VTAIL.n11 VTAIL.n10 585
R181 VTAIL.n13 VTAIL.n12 585
R182 VTAIL.n57 VTAIL.n56 585
R183 VTAIL.n55 VTAIL.n54 585
R184 VTAIL.n50 VTAIL.n49 585
R185 VTAIL.n37 VTAIL.n36 585
R186 VTAIL.n35 VTAIL.n34 585
R187 VTAIL.n30 VTAIL.n29 585
R188 VTAIL.n67 VTAIL.t11 338.558
R189 VTAIL.n7 VTAIL.t3 338.558
R190 VTAIL.n31 VTAIL.t14 338.558
R191 VTAIL.n51 VTAIL.t1 338.558
R192 VTAIL.n71 VTAIL.n65 171.744
R193 VTAIL.n72 VTAIL.n71 171.744
R194 VTAIL.n11 VTAIL.n5 171.744
R195 VTAIL.n12 VTAIL.n11 171.744
R196 VTAIL.n56 VTAIL.n55 171.744
R197 VTAIL.n55 VTAIL.n49 171.744
R198 VTAIL.n36 VTAIL.n35 171.744
R199 VTAIL.n35 VTAIL.n29 171.744
R200 VTAIL.n79 VTAIL.n78 110.688
R201 VTAIL.n1 VTAIL.n0 110.688
R202 VTAIL.n19 VTAIL.n18 110.688
R203 VTAIL.n21 VTAIL.n20 110.688
R204 VTAIL.n45 VTAIL.n44 110.688
R205 VTAIL.n43 VTAIL.n42 110.688
R206 VTAIL.n25 VTAIL.n24 110.688
R207 VTAIL.n23 VTAIL.n22 110.688
R208 VTAIL.t11 VTAIL.n65 85.8723
R209 VTAIL.t3 VTAIL.n5 85.8723
R210 VTAIL.t1 VTAIL.n49 85.8723
R211 VTAIL.t14 VTAIL.n29 85.8723
R212 VTAIL.n77 VTAIL.n76 30.6338
R213 VTAIL.n17 VTAIL.n16 30.6338
R214 VTAIL.n61 VTAIL.n60 30.6338
R215 VTAIL.n41 VTAIL.n40 30.6338
R216 VTAIL.n23 VTAIL.n21 19.3669
R217 VTAIL.n77 VTAIL.n61 17.3324
R218 VTAIL.n67 VTAIL.n66 10.6058
R219 VTAIL.n7 VTAIL.n6 10.6058
R220 VTAIL.n51 VTAIL.n50 10.6058
R221 VTAIL.n31 VTAIL.n30 10.6058
R222 VTAIL.n76 VTAIL.n62 9.69747
R223 VTAIL.n16 VTAIL.n2 9.69747
R224 VTAIL.n60 VTAIL.n46 9.69747
R225 VTAIL.n40 VTAIL.n26 9.69747
R226 VTAIL.n78 VTAIL.t15 9.56079
R227 VTAIL.n78 VTAIL.t19 9.56079
R228 VTAIL.n0 VTAIL.t10 9.56079
R229 VTAIL.n0 VTAIL.t16 9.56079
R230 VTAIL.n18 VTAIL.t2 9.56079
R231 VTAIL.n18 VTAIL.t7 9.56079
R232 VTAIL.n20 VTAIL.t5 9.56079
R233 VTAIL.n20 VTAIL.t4 9.56079
R234 VTAIL.n44 VTAIL.t6 9.56079
R235 VTAIL.n44 VTAIL.t9 9.56079
R236 VTAIL.n42 VTAIL.t0 9.56079
R237 VTAIL.n42 VTAIL.t8 9.56079
R238 VTAIL.n24 VTAIL.t12 9.56079
R239 VTAIL.n24 VTAIL.t18 9.56079
R240 VTAIL.n22 VTAIL.t13 9.56079
R241 VTAIL.n22 VTAIL.t17 9.56079
R242 VTAIL.n76 VTAIL.n75 9.45567
R243 VTAIL.n16 VTAIL.n15 9.45567
R244 VTAIL.n60 VTAIL.n59 9.45567
R245 VTAIL.n40 VTAIL.n39 9.45567
R246 VTAIL.n69 VTAIL.n68 9.3005
R247 VTAIL.n64 VTAIL.n63 9.3005
R248 VTAIL.n75 VTAIL.n74 9.3005
R249 VTAIL.n9 VTAIL.n8 9.3005
R250 VTAIL.n4 VTAIL.n3 9.3005
R251 VTAIL.n15 VTAIL.n14 9.3005
R252 VTAIL.n48 VTAIL.n47 9.3005
R253 VTAIL.n53 VTAIL.n52 9.3005
R254 VTAIL.n59 VTAIL.n58 9.3005
R255 VTAIL.n28 VTAIL.n27 9.3005
R256 VTAIL.n39 VTAIL.n38 9.3005
R257 VTAIL.n33 VTAIL.n32 9.3005
R258 VTAIL.n74 VTAIL.n73 8.92171
R259 VTAIL.n14 VTAIL.n13 8.92171
R260 VTAIL.n58 VTAIL.n57 8.92171
R261 VTAIL.n38 VTAIL.n37 8.92171
R262 VTAIL.n70 VTAIL.n64 8.14595
R263 VTAIL.n10 VTAIL.n4 8.14595
R264 VTAIL.n54 VTAIL.n48 8.14595
R265 VTAIL.n34 VTAIL.n28 8.14595
R266 VTAIL.n69 VTAIL.n66 7.3702
R267 VTAIL.n9 VTAIL.n6 7.3702
R268 VTAIL.n53 VTAIL.n50 7.3702
R269 VTAIL.n33 VTAIL.n30 7.3702
R270 VTAIL.n70 VTAIL.n69 5.81868
R271 VTAIL.n10 VTAIL.n9 5.81868
R272 VTAIL.n54 VTAIL.n53 5.81868
R273 VTAIL.n34 VTAIL.n33 5.81868
R274 VTAIL.n73 VTAIL.n64 5.04292
R275 VTAIL.n13 VTAIL.n4 5.04292
R276 VTAIL.n57 VTAIL.n48 5.04292
R277 VTAIL.n37 VTAIL.n28 5.04292
R278 VTAIL.n74 VTAIL.n62 4.26717
R279 VTAIL.n14 VTAIL.n2 4.26717
R280 VTAIL.n58 VTAIL.n46 4.26717
R281 VTAIL.n38 VTAIL.n26 4.26717
R282 VTAIL.n68 VTAIL.n67 2.5326
R283 VTAIL.n8 VTAIL.n7 2.5326
R284 VTAIL.n52 VTAIL.n51 2.5326
R285 VTAIL.n32 VTAIL.n31 2.5326
R286 VTAIL.n25 VTAIL.n23 2.03498
R287 VTAIL.n41 VTAIL.n25 2.03498
R288 VTAIL.n45 VTAIL.n43 2.03498
R289 VTAIL.n61 VTAIL.n45 2.03498
R290 VTAIL.n21 VTAIL.n19 2.03498
R291 VTAIL.n19 VTAIL.n17 2.03498
R292 VTAIL.n79 VTAIL.n77 2.03498
R293 VTAIL VTAIL.n1 1.58455
R294 VTAIL.n43 VTAIL.n41 1.48757
R295 VTAIL.n17 VTAIL.n1 1.48757
R296 VTAIL VTAIL.n79 0.450931
R297 VTAIL.n68 VTAIL.n63 0.155672
R298 VTAIL.n75 VTAIL.n63 0.155672
R299 VTAIL.n8 VTAIL.n3 0.155672
R300 VTAIL.n15 VTAIL.n3 0.155672
R301 VTAIL.n59 VTAIL.n47 0.155672
R302 VTAIL.n52 VTAIL.n47 0.155672
R303 VTAIL.n39 VTAIL.n27 0.155672
R304 VTAIL.n32 VTAIL.n27 0.155672
R305 VP.n20 VP.n19 161.3
R306 VP.n21 VP.n16 161.3
R307 VP.n23 VP.n22 161.3
R308 VP.n24 VP.n15 161.3
R309 VP.n26 VP.n25 161.3
R310 VP.n28 VP.n14 161.3
R311 VP.n30 VP.n29 161.3
R312 VP.n31 VP.n13 161.3
R313 VP.n33 VP.n32 161.3
R314 VP.n34 VP.n12 161.3
R315 VP.n37 VP.n36 161.3
R316 VP.n38 VP.n11 161.3
R317 VP.n40 VP.n39 161.3
R318 VP.n41 VP.n10 161.3
R319 VP.n74 VP.n0 161.3
R320 VP.n73 VP.n72 161.3
R321 VP.n71 VP.n1 161.3
R322 VP.n70 VP.n69 161.3
R323 VP.n67 VP.n2 161.3
R324 VP.n66 VP.n65 161.3
R325 VP.n64 VP.n3 161.3
R326 VP.n63 VP.n62 161.3
R327 VP.n61 VP.n4 161.3
R328 VP.n59 VP.n58 161.3
R329 VP.n57 VP.n5 161.3
R330 VP.n56 VP.n55 161.3
R331 VP.n54 VP.n6 161.3
R332 VP.n53 VP.n52 161.3
R333 VP.n51 VP.n50 161.3
R334 VP.n49 VP.n8 161.3
R335 VP.n48 VP.n47 161.3
R336 VP.n46 VP.n9 161.3
R337 VP.n45 VP.n44 87.7919
R338 VP.n76 VP.n75 87.7919
R339 VP.n43 VP.n42 87.7919
R340 VP.n18 VP.t3 71.3343
R341 VP.n18 VP.n17 65.0363
R342 VP.n49 VP.n48 56.5617
R343 VP.n73 VP.n1 56.5617
R344 VP.n40 VP.n11 56.5617
R345 VP.n55 VP.n5 47.3584
R346 VP.n62 VP.n3 47.3584
R347 VP.n29 VP.n13 47.3584
R348 VP.n22 VP.n15 47.3584
R349 VP.n45 VP.n43 43.583
R350 VP.n44 VP.t5 40.365
R351 VP.n7 VP.t9 40.365
R352 VP.n60 VP.t4 40.365
R353 VP.n68 VP.t2 40.365
R354 VP.n75 VP.t6 40.365
R355 VP.n42 VP.t0 40.365
R356 VP.n35 VP.t7 40.365
R357 VP.n27 VP.t1 40.365
R358 VP.n17 VP.t8 40.365
R359 VP.n55 VP.n54 33.7956
R360 VP.n66 VP.n3 33.7956
R361 VP.n33 VP.n13 33.7956
R362 VP.n22 VP.n21 33.7956
R363 VP.n48 VP.n9 24.5923
R364 VP.n50 VP.n49 24.5923
R365 VP.n54 VP.n53 24.5923
R366 VP.n59 VP.n5 24.5923
R367 VP.n62 VP.n61 24.5923
R368 VP.n67 VP.n66 24.5923
R369 VP.n69 VP.n1 24.5923
R370 VP.n74 VP.n73 24.5923
R371 VP.n41 VP.n40 24.5923
R372 VP.n34 VP.n33 24.5923
R373 VP.n36 VP.n11 24.5923
R374 VP.n26 VP.n15 24.5923
R375 VP.n29 VP.n28 24.5923
R376 VP.n21 VP.n20 24.5923
R377 VP.n44 VP.n9 23.1168
R378 VP.n75 VP.n74 23.1168
R379 VP.n42 VP.n41 23.1168
R380 VP.n50 VP.n7 19.1821
R381 VP.n69 VP.n68 19.1821
R382 VP.n36 VP.n35 19.1821
R383 VP.n19 VP.n18 12.856
R384 VP.n60 VP.n59 12.2964
R385 VP.n61 VP.n60 12.2964
R386 VP.n27 VP.n26 12.2964
R387 VP.n28 VP.n27 12.2964
R388 VP.n53 VP.n7 5.4107
R389 VP.n68 VP.n67 5.4107
R390 VP.n35 VP.n34 5.4107
R391 VP.n20 VP.n17 5.4107
R392 VP.n43 VP.n10 0.278335
R393 VP.n46 VP.n45 0.278335
R394 VP.n76 VP.n0 0.278335
R395 VP.n19 VP.n16 0.189894
R396 VP.n23 VP.n16 0.189894
R397 VP.n24 VP.n23 0.189894
R398 VP.n25 VP.n24 0.189894
R399 VP.n25 VP.n14 0.189894
R400 VP.n30 VP.n14 0.189894
R401 VP.n31 VP.n30 0.189894
R402 VP.n32 VP.n31 0.189894
R403 VP.n32 VP.n12 0.189894
R404 VP.n37 VP.n12 0.189894
R405 VP.n38 VP.n37 0.189894
R406 VP.n39 VP.n38 0.189894
R407 VP.n39 VP.n10 0.189894
R408 VP.n47 VP.n46 0.189894
R409 VP.n47 VP.n8 0.189894
R410 VP.n51 VP.n8 0.189894
R411 VP.n52 VP.n51 0.189894
R412 VP.n52 VP.n6 0.189894
R413 VP.n56 VP.n6 0.189894
R414 VP.n57 VP.n56 0.189894
R415 VP.n58 VP.n57 0.189894
R416 VP.n58 VP.n4 0.189894
R417 VP.n63 VP.n4 0.189894
R418 VP.n64 VP.n63 0.189894
R419 VP.n65 VP.n64 0.189894
R420 VP.n65 VP.n2 0.189894
R421 VP.n70 VP.n2 0.189894
R422 VP.n71 VP.n70 0.189894
R423 VP.n72 VP.n71 0.189894
R424 VP.n72 VP.n0 0.189894
R425 VP VP.n76 0.153485
R426 VDD1.n10 VDD1.n0 756.745
R427 VDD1.n27 VDD1.n17 756.745
R428 VDD1.n11 VDD1.n10 585
R429 VDD1.n9 VDD1.n8 585
R430 VDD1.n4 VDD1.n3 585
R431 VDD1.n21 VDD1.n20 585
R432 VDD1.n26 VDD1.n25 585
R433 VDD1.n28 VDD1.n27 585
R434 VDD1.n5 VDD1.t6 338.558
R435 VDD1.n22 VDD1.t4 338.558
R436 VDD1.n10 VDD1.n9 171.744
R437 VDD1.n9 VDD1.n3 171.744
R438 VDD1.n26 VDD1.n20 171.744
R439 VDD1.n27 VDD1.n26 171.744
R440 VDD1.n35 VDD1.n34 128.837
R441 VDD1.n37 VDD1.n36 127.367
R442 VDD1.n16 VDD1.n15 127.367
R443 VDD1.n33 VDD1.n32 127.367
R444 VDD1.t6 VDD1.n3 85.8723
R445 VDD1.t4 VDD1.n20 85.8723
R446 VDD1.n16 VDD1.n14 49.3471
R447 VDD1.n33 VDD1.n31 49.3471
R448 VDD1.n37 VDD1.n35 37.9104
R449 VDD1.n5 VDD1.n4 10.6058
R450 VDD1.n22 VDD1.n21 10.6058
R451 VDD1.n14 VDD1.n0 9.69747
R452 VDD1.n31 VDD1.n17 9.69747
R453 VDD1.n36 VDD1.t2 9.56079
R454 VDD1.n36 VDD1.t9 9.56079
R455 VDD1.n15 VDD1.t1 9.56079
R456 VDD1.n15 VDD1.t8 9.56079
R457 VDD1.n34 VDD1.t7 9.56079
R458 VDD1.n34 VDD1.t3 9.56079
R459 VDD1.n32 VDD1.t0 9.56079
R460 VDD1.n32 VDD1.t5 9.56079
R461 VDD1.n14 VDD1.n13 9.45567
R462 VDD1.n31 VDD1.n30 9.45567
R463 VDD1.n2 VDD1.n1 9.3005
R464 VDD1.n13 VDD1.n12 9.3005
R465 VDD1.n7 VDD1.n6 9.3005
R466 VDD1.n24 VDD1.n23 9.3005
R467 VDD1.n19 VDD1.n18 9.3005
R468 VDD1.n30 VDD1.n29 9.3005
R469 VDD1.n12 VDD1.n11 8.92171
R470 VDD1.n29 VDD1.n28 8.92171
R471 VDD1.n8 VDD1.n2 8.14595
R472 VDD1.n25 VDD1.n19 8.14595
R473 VDD1.n7 VDD1.n4 7.3702
R474 VDD1.n24 VDD1.n21 7.3702
R475 VDD1.n8 VDD1.n7 5.81868
R476 VDD1.n25 VDD1.n24 5.81868
R477 VDD1.n11 VDD1.n2 5.04292
R478 VDD1.n28 VDD1.n19 5.04292
R479 VDD1.n12 VDD1.n0 4.26717
R480 VDD1.n29 VDD1.n17 4.26717
R481 VDD1.n6 VDD1.n5 2.5326
R482 VDD1.n23 VDD1.n22 2.5326
R483 VDD1 VDD1.n37 1.46817
R484 VDD1 VDD1.n16 0.56731
R485 VDD1.n35 VDD1.n33 0.453775
R486 VDD1.n13 VDD1.n1 0.155672
R487 VDD1.n6 VDD1.n1 0.155672
R488 VDD1.n23 VDD1.n18 0.155672
R489 VDD1.n30 VDD1.n18 0.155672
R490 B.n288 B.n287 585
R491 B.n286 B.n103 585
R492 B.n285 B.n284 585
R493 B.n283 B.n104 585
R494 B.n282 B.n281 585
R495 B.n280 B.n105 585
R496 B.n279 B.n278 585
R497 B.n277 B.n106 585
R498 B.n276 B.n275 585
R499 B.n274 B.n107 585
R500 B.n273 B.n272 585
R501 B.n271 B.n108 585
R502 B.n270 B.n269 585
R503 B.n268 B.n109 585
R504 B.n267 B.n266 585
R505 B.n265 B.n110 585
R506 B.n263 B.n262 585
R507 B.n261 B.n113 585
R508 B.n260 B.n259 585
R509 B.n258 B.n114 585
R510 B.n257 B.n256 585
R511 B.n255 B.n115 585
R512 B.n254 B.n253 585
R513 B.n252 B.n116 585
R514 B.n251 B.n250 585
R515 B.n249 B.n117 585
R516 B.n248 B.n247 585
R517 B.n243 B.n118 585
R518 B.n242 B.n241 585
R519 B.n240 B.n119 585
R520 B.n239 B.n238 585
R521 B.n237 B.n120 585
R522 B.n236 B.n235 585
R523 B.n234 B.n121 585
R524 B.n233 B.n232 585
R525 B.n231 B.n122 585
R526 B.n230 B.n229 585
R527 B.n228 B.n123 585
R528 B.n227 B.n226 585
R529 B.n225 B.n124 585
R530 B.n224 B.n223 585
R531 B.n222 B.n125 585
R532 B.n289 B.n102 585
R533 B.n291 B.n290 585
R534 B.n292 B.n101 585
R535 B.n294 B.n293 585
R536 B.n295 B.n100 585
R537 B.n297 B.n296 585
R538 B.n298 B.n99 585
R539 B.n300 B.n299 585
R540 B.n301 B.n98 585
R541 B.n303 B.n302 585
R542 B.n304 B.n97 585
R543 B.n306 B.n305 585
R544 B.n307 B.n96 585
R545 B.n309 B.n308 585
R546 B.n310 B.n95 585
R547 B.n312 B.n311 585
R548 B.n313 B.n94 585
R549 B.n315 B.n314 585
R550 B.n316 B.n93 585
R551 B.n318 B.n317 585
R552 B.n319 B.n92 585
R553 B.n321 B.n320 585
R554 B.n322 B.n91 585
R555 B.n324 B.n323 585
R556 B.n325 B.n90 585
R557 B.n327 B.n326 585
R558 B.n328 B.n89 585
R559 B.n330 B.n329 585
R560 B.n331 B.n88 585
R561 B.n333 B.n332 585
R562 B.n334 B.n87 585
R563 B.n336 B.n335 585
R564 B.n337 B.n86 585
R565 B.n339 B.n338 585
R566 B.n340 B.n85 585
R567 B.n342 B.n341 585
R568 B.n343 B.n84 585
R569 B.n345 B.n344 585
R570 B.n346 B.n83 585
R571 B.n348 B.n347 585
R572 B.n349 B.n82 585
R573 B.n351 B.n350 585
R574 B.n352 B.n81 585
R575 B.n354 B.n353 585
R576 B.n355 B.n80 585
R577 B.n357 B.n356 585
R578 B.n358 B.n79 585
R579 B.n360 B.n359 585
R580 B.n361 B.n78 585
R581 B.n363 B.n362 585
R582 B.n364 B.n77 585
R583 B.n366 B.n365 585
R584 B.n367 B.n76 585
R585 B.n369 B.n368 585
R586 B.n370 B.n75 585
R587 B.n372 B.n371 585
R588 B.n373 B.n74 585
R589 B.n375 B.n374 585
R590 B.n376 B.n73 585
R591 B.n378 B.n377 585
R592 B.n379 B.n72 585
R593 B.n381 B.n380 585
R594 B.n382 B.n71 585
R595 B.n384 B.n383 585
R596 B.n385 B.n70 585
R597 B.n387 B.n386 585
R598 B.n388 B.n69 585
R599 B.n390 B.n389 585
R600 B.n391 B.n68 585
R601 B.n393 B.n392 585
R602 B.n394 B.n67 585
R603 B.n396 B.n395 585
R604 B.n397 B.n66 585
R605 B.n399 B.n398 585
R606 B.n400 B.n65 585
R607 B.n402 B.n401 585
R608 B.n403 B.n64 585
R609 B.n405 B.n404 585
R610 B.n406 B.n63 585
R611 B.n408 B.n407 585
R612 B.n409 B.n62 585
R613 B.n411 B.n410 585
R614 B.n412 B.n61 585
R615 B.n414 B.n413 585
R616 B.n415 B.n60 585
R617 B.n417 B.n416 585
R618 B.n418 B.n59 585
R619 B.n420 B.n419 585
R620 B.n421 B.n58 585
R621 B.n423 B.n422 585
R622 B.n424 B.n57 585
R623 B.n426 B.n425 585
R624 B.n427 B.n56 585
R625 B.n429 B.n428 585
R626 B.n430 B.n55 585
R627 B.n432 B.n431 585
R628 B.n433 B.n54 585
R629 B.n435 B.n434 585
R630 B.n436 B.n53 585
R631 B.n438 B.n437 585
R632 B.n502 B.n501 585
R633 B.n500 B.n27 585
R634 B.n499 B.n498 585
R635 B.n497 B.n28 585
R636 B.n496 B.n495 585
R637 B.n494 B.n29 585
R638 B.n493 B.n492 585
R639 B.n491 B.n30 585
R640 B.n490 B.n489 585
R641 B.n488 B.n31 585
R642 B.n487 B.n486 585
R643 B.n485 B.n32 585
R644 B.n484 B.n483 585
R645 B.n482 B.n33 585
R646 B.n481 B.n480 585
R647 B.n479 B.n34 585
R648 B.n478 B.n477 585
R649 B.n476 B.n35 585
R650 B.n475 B.n474 585
R651 B.n473 B.n39 585
R652 B.n472 B.n471 585
R653 B.n470 B.n40 585
R654 B.n469 B.n468 585
R655 B.n467 B.n41 585
R656 B.n466 B.n465 585
R657 B.n464 B.n42 585
R658 B.n462 B.n461 585
R659 B.n460 B.n45 585
R660 B.n459 B.n458 585
R661 B.n457 B.n46 585
R662 B.n456 B.n455 585
R663 B.n454 B.n47 585
R664 B.n453 B.n452 585
R665 B.n451 B.n48 585
R666 B.n450 B.n449 585
R667 B.n448 B.n49 585
R668 B.n447 B.n446 585
R669 B.n445 B.n50 585
R670 B.n444 B.n443 585
R671 B.n442 B.n51 585
R672 B.n441 B.n440 585
R673 B.n439 B.n52 585
R674 B.n503 B.n26 585
R675 B.n505 B.n504 585
R676 B.n506 B.n25 585
R677 B.n508 B.n507 585
R678 B.n509 B.n24 585
R679 B.n511 B.n510 585
R680 B.n512 B.n23 585
R681 B.n514 B.n513 585
R682 B.n515 B.n22 585
R683 B.n517 B.n516 585
R684 B.n518 B.n21 585
R685 B.n520 B.n519 585
R686 B.n521 B.n20 585
R687 B.n523 B.n522 585
R688 B.n524 B.n19 585
R689 B.n526 B.n525 585
R690 B.n527 B.n18 585
R691 B.n529 B.n528 585
R692 B.n530 B.n17 585
R693 B.n532 B.n531 585
R694 B.n533 B.n16 585
R695 B.n535 B.n534 585
R696 B.n536 B.n15 585
R697 B.n538 B.n537 585
R698 B.n539 B.n14 585
R699 B.n541 B.n540 585
R700 B.n542 B.n13 585
R701 B.n544 B.n543 585
R702 B.n545 B.n12 585
R703 B.n547 B.n546 585
R704 B.n548 B.n11 585
R705 B.n550 B.n549 585
R706 B.n551 B.n10 585
R707 B.n553 B.n552 585
R708 B.n554 B.n9 585
R709 B.n556 B.n555 585
R710 B.n557 B.n8 585
R711 B.n559 B.n558 585
R712 B.n560 B.n7 585
R713 B.n562 B.n561 585
R714 B.n563 B.n6 585
R715 B.n565 B.n564 585
R716 B.n566 B.n5 585
R717 B.n568 B.n567 585
R718 B.n569 B.n4 585
R719 B.n571 B.n570 585
R720 B.n572 B.n3 585
R721 B.n574 B.n573 585
R722 B.n575 B.n0 585
R723 B.n2 B.n1 585
R724 B.n150 B.n149 585
R725 B.n152 B.n151 585
R726 B.n153 B.n148 585
R727 B.n155 B.n154 585
R728 B.n156 B.n147 585
R729 B.n158 B.n157 585
R730 B.n159 B.n146 585
R731 B.n161 B.n160 585
R732 B.n162 B.n145 585
R733 B.n164 B.n163 585
R734 B.n165 B.n144 585
R735 B.n167 B.n166 585
R736 B.n168 B.n143 585
R737 B.n170 B.n169 585
R738 B.n171 B.n142 585
R739 B.n173 B.n172 585
R740 B.n174 B.n141 585
R741 B.n176 B.n175 585
R742 B.n177 B.n140 585
R743 B.n179 B.n178 585
R744 B.n180 B.n139 585
R745 B.n182 B.n181 585
R746 B.n183 B.n138 585
R747 B.n185 B.n184 585
R748 B.n186 B.n137 585
R749 B.n188 B.n187 585
R750 B.n189 B.n136 585
R751 B.n191 B.n190 585
R752 B.n192 B.n135 585
R753 B.n194 B.n193 585
R754 B.n195 B.n134 585
R755 B.n197 B.n196 585
R756 B.n198 B.n133 585
R757 B.n200 B.n199 585
R758 B.n201 B.n132 585
R759 B.n203 B.n202 585
R760 B.n204 B.n131 585
R761 B.n206 B.n205 585
R762 B.n207 B.n130 585
R763 B.n209 B.n208 585
R764 B.n210 B.n129 585
R765 B.n212 B.n211 585
R766 B.n213 B.n128 585
R767 B.n215 B.n214 585
R768 B.n216 B.n127 585
R769 B.n218 B.n217 585
R770 B.n219 B.n126 585
R771 B.n221 B.n220 585
R772 B.n222 B.n221 559.769
R773 B.n287 B.n102 559.769
R774 B.n437 B.n52 559.769
R775 B.n503 B.n502 559.769
R776 B.n111 B.t10 275.209
R777 B.n43 B.t5 275.209
R778 B.n244 B.t1 275.209
R779 B.n36 B.t8 275.209
R780 B.n577 B.n576 256.663
R781 B.n244 B.t0 247.352
R782 B.n111 B.t9 247.352
R783 B.n43 B.t3 247.352
R784 B.n36 B.t6 247.352
R785 B.n576 B.n575 235.042
R786 B.n576 B.n2 235.042
R787 B.n112 B.t11 229.44
R788 B.n44 B.t4 229.44
R789 B.n245 B.t2 229.44
R790 B.n37 B.t7 229.44
R791 B.n223 B.n222 163.367
R792 B.n223 B.n124 163.367
R793 B.n227 B.n124 163.367
R794 B.n228 B.n227 163.367
R795 B.n229 B.n228 163.367
R796 B.n229 B.n122 163.367
R797 B.n233 B.n122 163.367
R798 B.n234 B.n233 163.367
R799 B.n235 B.n234 163.367
R800 B.n235 B.n120 163.367
R801 B.n239 B.n120 163.367
R802 B.n240 B.n239 163.367
R803 B.n241 B.n240 163.367
R804 B.n241 B.n118 163.367
R805 B.n248 B.n118 163.367
R806 B.n249 B.n248 163.367
R807 B.n250 B.n249 163.367
R808 B.n250 B.n116 163.367
R809 B.n254 B.n116 163.367
R810 B.n255 B.n254 163.367
R811 B.n256 B.n255 163.367
R812 B.n256 B.n114 163.367
R813 B.n260 B.n114 163.367
R814 B.n261 B.n260 163.367
R815 B.n262 B.n261 163.367
R816 B.n262 B.n110 163.367
R817 B.n267 B.n110 163.367
R818 B.n268 B.n267 163.367
R819 B.n269 B.n268 163.367
R820 B.n269 B.n108 163.367
R821 B.n273 B.n108 163.367
R822 B.n274 B.n273 163.367
R823 B.n275 B.n274 163.367
R824 B.n275 B.n106 163.367
R825 B.n279 B.n106 163.367
R826 B.n280 B.n279 163.367
R827 B.n281 B.n280 163.367
R828 B.n281 B.n104 163.367
R829 B.n285 B.n104 163.367
R830 B.n286 B.n285 163.367
R831 B.n287 B.n286 163.367
R832 B.n437 B.n436 163.367
R833 B.n436 B.n435 163.367
R834 B.n435 B.n54 163.367
R835 B.n431 B.n54 163.367
R836 B.n431 B.n430 163.367
R837 B.n430 B.n429 163.367
R838 B.n429 B.n56 163.367
R839 B.n425 B.n56 163.367
R840 B.n425 B.n424 163.367
R841 B.n424 B.n423 163.367
R842 B.n423 B.n58 163.367
R843 B.n419 B.n58 163.367
R844 B.n419 B.n418 163.367
R845 B.n418 B.n417 163.367
R846 B.n417 B.n60 163.367
R847 B.n413 B.n60 163.367
R848 B.n413 B.n412 163.367
R849 B.n412 B.n411 163.367
R850 B.n411 B.n62 163.367
R851 B.n407 B.n62 163.367
R852 B.n407 B.n406 163.367
R853 B.n406 B.n405 163.367
R854 B.n405 B.n64 163.367
R855 B.n401 B.n64 163.367
R856 B.n401 B.n400 163.367
R857 B.n400 B.n399 163.367
R858 B.n399 B.n66 163.367
R859 B.n395 B.n66 163.367
R860 B.n395 B.n394 163.367
R861 B.n394 B.n393 163.367
R862 B.n393 B.n68 163.367
R863 B.n389 B.n68 163.367
R864 B.n389 B.n388 163.367
R865 B.n388 B.n387 163.367
R866 B.n387 B.n70 163.367
R867 B.n383 B.n70 163.367
R868 B.n383 B.n382 163.367
R869 B.n382 B.n381 163.367
R870 B.n381 B.n72 163.367
R871 B.n377 B.n72 163.367
R872 B.n377 B.n376 163.367
R873 B.n376 B.n375 163.367
R874 B.n375 B.n74 163.367
R875 B.n371 B.n74 163.367
R876 B.n371 B.n370 163.367
R877 B.n370 B.n369 163.367
R878 B.n369 B.n76 163.367
R879 B.n365 B.n76 163.367
R880 B.n365 B.n364 163.367
R881 B.n364 B.n363 163.367
R882 B.n363 B.n78 163.367
R883 B.n359 B.n78 163.367
R884 B.n359 B.n358 163.367
R885 B.n358 B.n357 163.367
R886 B.n357 B.n80 163.367
R887 B.n353 B.n80 163.367
R888 B.n353 B.n352 163.367
R889 B.n352 B.n351 163.367
R890 B.n351 B.n82 163.367
R891 B.n347 B.n82 163.367
R892 B.n347 B.n346 163.367
R893 B.n346 B.n345 163.367
R894 B.n345 B.n84 163.367
R895 B.n341 B.n84 163.367
R896 B.n341 B.n340 163.367
R897 B.n340 B.n339 163.367
R898 B.n339 B.n86 163.367
R899 B.n335 B.n86 163.367
R900 B.n335 B.n334 163.367
R901 B.n334 B.n333 163.367
R902 B.n333 B.n88 163.367
R903 B.n329 B.n88 163.367
R904 B.n329 B.n328 163.367
R905 B.n328 B.n327 163.367
R906 B.n327 B.n90 163.367
R907 B.n323 B.n90 163.367
R908 B.n323 B.n322 163.367
R909 B.n322 B.n321 163.367
R910 B.n321 B.n92 163.367
R911 B.n317 B.n92 163.367
R912 B.n317 B.n316 163.367
R913 B.n316 B.n315 163.367
R914 B.n315 B.n94 163.367
R915 B.n311 B.n94 163.367
R916 B.n311 B.n310 163.367
R917 B.n310 B.n309 163.367
R918 B.n309 B.n96 163.367
R919 B.n305 B.n96 163.367
R920 B.n305 B.n304 163.367
R921 B.n304 B.n303 163.367
R922 B.n303 B.n98 163.367
R923 B.n299 B.n98 163.367
R924 B.n299 B.n298 163.367
R925 B.n298 B.n297 163.367
R926 B.n297 B.n100 163.367
R927 B.n293 B.n100 163.367
R928 B.n293 B.n292 163.367
R929 B.n292 B.n291 163.367
R930 B.n291 B.n102 163.367
R931 B.n502 B.n27 163.367
R932 B.n498 B.n27 163.367
R933 B.n498 B.n497 163.367
R934 B.n497 B.n496 163.367
R935 B.n496 B.n29 163.367
R936 B.n492 B.n29 163.367
R937 B.n492 B.n491 163.367
R938 B.n491 B.n490 163.367
R939 B.n490 B.n31 163.367
R940 B.n486 B.n31 163.367
R941 B.n486 B.n485 163.367
R942 B.n485 B.n484 163.367
R943 B.n484 B.n33 163.367
R944 B.n480 B.n33 163.367
R945 B.n480 B.n479 163.367
R946 B.n479 B.n478 163.367
R947 B.n478 B.n35 163.367
R948 B.n474 B.n35 163.367
R949 B.n474 B.n473 163.367
R950 B.n473 B.n472 163.367
R951 B.n472 B.n40 163.367
R952 B.n468 B.n40 163.367
R953 B.n468 B.n467 163.367
R954 B.n467 B.n466 163.367
R955 B.n466 B.n42 163.367
R956 B.n461 B.n42 163.367
R957 B.n461 B.n460 163.367
R958 B.n460 B.n459 163.367
R959 B.n459 B.n46 163.367
R960 B.n455 B.n46 163.367
R961 B.n455 B.n454 163.367
R962 B.n454 B.n453 163.367
R963 B.n453 B.n48 163.367
R964 B.n449 B.n48 163.367
R965 B.n449 B.n448 163.367
R966 B.n448 B.n447 163.367
R967 B.n447 B.n50 163.367
R968 B.n443 B.n50 163.367
R969 B.n443 B.n442 163.367
R970 B.n442 B.n441 163.367
R971 B.n441 B.n52 163.367
R972 B.n504 B.n503 163.367
R973 B.n504 B.n25 163.367
R974 B.n508 B.n25 163.367
R975 B.n509 B.n508 163.367
R976 B.n510 B.n509 163.367
R977 B.n510 B.n23 163.367
R978 B.n514 B.n23 163.367
R979 B.n515 B.n514 163.367
R980 B.n516 B.n515 163.367
R981 B.n516 B.n21 163.367
R982 B.n520 B.n21 163.367
R983 B.n521 B.n520 163.367
R984 B.n522 B.n521 163.367
R985 B.n522 B.n19 163.367
R986 B.n526 B.n19 163.367
R987 B.n527 B.n526 163.367
R988 B.n528 B.n527 163.367
R989 B.n528 B.n17 163.367
R990 B.n532 B.n17 163.367
R991 B.n533 B.n532 163.367
R992 B.n534 B.n533 163.367
R993 B.n534 B.n15 163.367
R994 B.n538 B.n15 163.367
R995 B.n539 B.n538 163.367
R996 B.n540 B.n539 163.367
R997 B.n540 B.n13 163.367
R998 B.n544 B.n13 163.367
R999 B.n545 B.n544 163.367
R1000 B.n546 B.n545 163.367
R1001 B.n546 B.n11 163.367
R1002 B.n550 B.n11 163.367
R1003 B.n551 B.n550 163.367
R1004 B.n552 B.n551 163.367
R1005 B.n552 B.n9 163.367
R1006 B.n556 B.n9 163.367
R1007 B.n557 B.n556 163.367
R1008 B.n558 B.n557 163.367
R1009 B.n558 B.n7 163.367
R1010 B.n562 B.n7 163.367
R1011 B.n563 B.n562 163.367
R1012 B.n564 B.n563 163.367
R1013 B.n564 B.n5 163.367
R1014 B.n568 B.n5 163.367
R1015 B.n569 B.n568 163.367
R1016 B.n570 B.n569 163.367
R1017 B.n570 B.n3 163.367
R1018 B.n574 B.n3 163.367
R1019 B.n575 B.n574 163.367
R1020 B.n150 B.n2 163.367
R1021 B.n151 B.n150 163.367
R1022 B.n151 B.n148 163.367
R1023 B.n155 B.n148 163.367
R1024 B.n156 B.n155 163.367
R1025 B.n157 B.n156 163.367
R1026 B.n157 B.n146 163.367
R1027 B.n161 B.n146 163.367
R1028 B.n162 B.n161 163.367
R1029 B.n163 B.n162 163.367
R1030 B.n163 B.n144 163.367
R1031 B.n167 B.n144 163.367
R1032 B.n168 B.n167 163.367
R1033 B.n169 B.n168 163.367
R1034 B.n169 B.n142 163.367
R1035 B.n173 B.n142 163.367
R1036 B.n174 B.n173 163.367
R1037 B.n175 B.n174 163.367
R1038 B.n175 B.n140 163.367
R1039 B.n179 B.n140 163.367
R1040 B.n180 B.n179 163.367
R1041 B.n181 B.n180 163.367
R1042 B.n181 B.n138 163.367
R1043 B.n185 B.n138 163.367
R1044 B.n186 B.n185 163.367
R1045 B.n187 B.n186 163.367
R1046 B.n187 B.n136 163.367
R1047 B.n191 B.n136 163.367
R1048 B.n192 B.n191 163.367
R1049 B.n193 B.n192 163.367
R1050 B.n193 B.n134 163.367
R1051 B.n197 B.n134 163.367
R1052 B.n198 B.n197 163.367
R1053 B.n199 B.n198 163.367
R1054 B.n199 B.n132 163.367
R1055 B.n203 B.n132 163.367
R1056 B.n204 B.n203 163.367
R1057 B.n205 B.n204 163.367
R1058 B.n205 B.n130 163.367
R1059 B.n209 B.n130 163.367
R1060 B.n210 B.n209 163.367
R1061 B.n211 B.n210 163.367
R1062 B.n211 B.n128 163.367
R1063 B.n215 B.n128 163.367
R1064 B.n216 B.n215 163.367
R1065 B.n217 B.n216 163.367
R1066 B.n217 B.n126 163.367
R1067 B.n221 B.n126 163.367
R1068 B.n246 B.n245 59.5399
R1069 B.n264 B.n112 59.5399
R1070 B.n463 B.n44 59.5399
R1071 B.n38 B.n37 59.5399
R1072 B.n245 B.n244 45.7702
R1073 B.n112 B.n111 45.7702
R1074 B.n44 B.n43 45.7702
R1075 B.n37 B.n36 45.7702
R1076 B.n289 B.n288 36.3712
R1077 B.n501 B.n26 36.3712
R1078 B.n439 B.n438 36.3712
R1079 B.n220 B.n125 36.3712
R1080 B B.n577 18.0485
R1081 B.n505 B.n26 10.6151
R1082 B.n506 B.n505 10.6151
R1083 B.n507 B.n506 10.6151
R1084 B.n507 B.n24 10.6151
R1085 B.n511 B.n24 10.6151
R1086 B.n512 B.n511 10.6151
R1087 B.n513 B.n512 10.6151
R1088 B.n513 B.n22 10.6151
R1089 B.n517 B.n22 10.6151
R1090 B.n518 B.n517 10.6151
R1091 B.n519 B.n518 10.6151
R1092 B.n519 B.n20 10.6151
R1093 B.n523 B.n20 10.6151
R1094 B.n524 B.n523 10.6151
R1095 B.n525 B.n524 10.6151
R1096 B.n525 B.n18 10.6151
R1097 B.n529 B.n18 10.6151
R1098 B.n530 B.n529 10.6151
R1099 B.n531 B.n530 10.6151
R1100 B.n531 B.n16 10.6151
R1101 B.n535 B.n16 10.6151
R1102 B.n536 B.n535 10.6151
R1103 B.n537 B.n536 10.6151
R1104 B.n537 B.n14 10.6151
R1105 B.n541 B.n14 10.6151
R1106 B.n542 B.n541 10.6151
R1107 B.n543 B.n542 10.6151
R1108 B.n543 B.n12 10.6151
R1109 B.n547 B.n12 10.6151
R1110 B.n548 B.n547 10.6151
R1111 B.n549 B.n548 10.6151
R1112 B.n549 B.n10 10.6151
R1113 B.n553 B.n10 10.6151
R1114 B.n554 B.n553 10.6151
R1115 B.n555 B.n554 10.6151
R1116 B.n555 B.n8 10.6151
R1117 B.n559 B.n8 10.6151
R1118 B.n560 B.n559 10.6151
R1119 B.n561 B.n560 10.6151
R1120 B.n561 B.n6 10.6151
R1121 B.n565 B.n6 10.6151
R1122 B.n566 B.n565 10.6151
R1123 B.n567 B.n566 10.6151
R1124 B.n567 B.n4 10.6151
R1125 B.n571 B.n4 10.6151
R1126 B.n572 B.n571 10.6151
R1127 B.n573 B.n572 10.6151
R1128 B.n573 B.n0 10.6151
R1129 B.n501 B.n500 10.6151
R1130 B.n500 B.n499 10.6151
R1131 B.n499 B.n28 10.6151
R1132 B.n495 B.n28 10.6151
R1133 B.n495 B.n494 10.6151
R1134 B.n494 B.n493 10.6151
R1135 B.n493 B.n30 10.6151
R1136 B.n489 B.n30 10.6151
R1137 B.n489 B.n488 10.6151
R1138 B.n488 B.n487 10.6151
R1139 B.n487 B.n32 10.6151
R1140 B.n483 B.n32 10.6151
R1141 B.n483 B.n482 10.6151
R1142 B.n482 B.n481 10.6151
R1143 B.n481 B.n34 10.6151
R1144 B.n477 B.n476 10.6151
R1145 B.n476 B.n475 10.6151
R1146 B.n475 B.n39 10.6151
R1147 B.n471 B.n39 10.6151
R1148 B.n471 B.n470 10.6151
R1149 B.n470 B.n469 10.6151
R1150 B.n469 B.n41 10.6151
R1151 B.n465 B.n41 10.6151
R1152 B.n465 B.n464 10.6151
R1153 B.n462 B.n45 10.6151
R1154 B.n458 B.n45 10.6151
R1155 B.n458 B.n457 10.6151
R1156 B.n457 B.n456 10.6151
R1157 B.n456 B.n47 10.6151
R1158 B.n452 B.n47 10.6151
R1159 B.n452 B.n451 10.6151
R1160 B.n451 B.n450 10.6151
R1161 B.n450 B.n49 10.6151
R1162 B.n446 B.n49 10.6151
R1163 B.n446 B.n445 10.6151
R1164 B.n445 B.n444 10.6151
R1165 B.n444 B.n51 10.6151
R1166 B.n440 B.n51 10.6151
R1167 B.n440 B.n439 10.6151
R1168 B.n438 B.n53 10.6151
R1169 B.n434 B.n53 10.6151
R1170 B.n434 B.n433 10.6151
R1171 B.n433 B.n432 10.6151
R1172 B.n432 B.n55 10.6151
R1173 B.n428 B.n55 10.6151
R1174 B.n428 B.n427 10.6151
R1175 B.n427 B.n426 10.6151
R1176 B.n426 B.n57 10.6151
R1177 B.n422 B.n57 10.6151
R1178 B.n422 B.n421 10.6151
R1179 B.n421 B.n420 10.6151
R1180 B.n420 B.n59 10.6151
R1181 B.n416 B.n59 10.6151
R1182 B.n416 B.n415 10.6151
R1183 B.n415 B.n414 10.6151
R1184 B.n414 B.n61 10.6151
R1185 B.n410 B.n61 10.6151
R1186 B.n410 B.n409 10.6151
R1187 B.n409 B.n408 10.6151
R1188 B.n408 B.n63 10.6151
R1189 B.n404 B.n63 10.6151
R1190 B.n404 B.n403 10.6151
R1191 B.n403 B.n402 10.6151
R1192 B.n402 B.n65 10.6151
R1193 B.n398 B.n65 10.6151
R1194 B.n398 B.n397 10.6151
R1195 B.n397 B.n396 10.6151
R1196 B.n396 B.n67 10.6151
R1197 B.n392 B.n67 10.6151
R1198 B.n392 B.n391 10.6151
R1199 B.n391 B.n390 10.6151
R1200 B.n390 B.n69 10.6151
R1201 B.n386 B.n69 10.6151
R1202 B.n386 B.n385 10.6151
R1203 B.n385 B.n384 10.6151
R1204 B.n384 B.n71 10.6151
R1205 B.n380 B.n71 10.6151
R1206 B.n380 B.n379 10.6151
R1207 B.n379 B.n378 10.6151
R1208 B.n378 B.n73 10.6151
R1209 B.n374 B.n73 10.6151
R1210 B.n374 B.n373 10.6151
R1211 B.n373 B.n372 10.6151
R1212 B.n372 B.n75 10.6151
R1213 B.n368 B.n75 10.6151
R1214 B.n368 B.n367 10.6151
R1215 B.n367 B.n366 10.6151
R1216 B.n366 B.n77 10.6151
R1217 B.n362 B.n77 10.6151
R1218 B.n362 B.n361 10.6151
R1219 B.n361 B.n360 10.6151
R1220 B.n360 B.n79 10.6151
R1221 B.n356 B.n79 10.6151
R1222 B.n356 B.n355 10.6151
R1223 B.n355 B.n354 10.6151
R1224 B.n354 B.n81 10.6151
R1225 B.n350 B.n81 10.6151
R1226 B.n350 B.n349 10.6151
R1227 B.n349 B.n348 10.6151
R1228 B.n348 B.n83 10.6151
R1229 B.n344 B.n83 10.6151
R1230 B.n344 B.n343 10.6151
R1231 B.n343 B.n342 10.6151
R1232 B.n342 B.n85 10.6151
R1233 B.n338 B.n85 10.6151
R1234 B.n338 B.n337 10.6151
R1235 B.n337 B.n336 10.6151
R1236 B.n336 B.n87 10.6151
R1237 B.n332 B.n87 10.6151
R1238 B.n332 B.n331 10.6151
R1239 B.n331 B.n330 10.6151
R1240 B.n330 B.n89 10.6151
R1241 B.n326 B.n89 10.6151
R1242 B.n326 B.n325 10.6151
R1243 B.n325 B.n324 10.6151
R1244 B.n324 B.n91 10.6151
R1245 B.n320 B.n91 10.6151
R1246 B.n320 B.n319 10.6151
R1247 B.n319 B.n318 10.6151
R1248 B.n318 B.n93 10.6151
R1249 B.n314 B.n93 10.6151
R1250 B.n314 B.n313 10.6151
R1251 B.n313 B.n312 10.6151
R1252 B.n312 B.n95 10.6151
R1253 B.n308 B.n95 10.6151
R1254 B.n308 B.n307 10.6151
R1255 B.n307 B.n306 10.6151
R1256 B.n306 B.n97 10.6151
R1257 B.n302 B.n97 10.6151
R1258 B.n302 B.n301 10.6151
R1259 B.n301 B.n300 10.6151
R1260 B.n300 B.n99 10.6151
R1261 B.n296 B.n99 10.6151
R1262 B.n296 B.n295 10.6151
R1263 B.n295 B.n294 10.6151
R1264 B.n294 B.n101 10.6151
R1265 B.n290 B.n101 10.6151
R1266 B.n290 B.n289 10.6151
R1267 B.n149 B.n1 10.6151
R1268 B.n152 B.n149 10.6151
R1269 B.n153 B.n152 10.6151
R1270 B.n154 B.n153 10.6151
R1271 B.n154 B.n147 10.6151
R1272 B.n158 B.n147 10.6151
R1273 B.n159 B.n158 10.6151
R1274 B.n160 B.n159 10.6151
R1275 B.n160 B.n145 10.6151
R1276 B.n164 B.n145 10.6151
R1277 B.n165 B.n164 10.6151
R1278 B.n166 B.n165 10.6151
R1279 B.n166 B.n143 10.6151
R1280 B.n170 B.n143 10.6151
R1281 B.n171 B.n170 10.6151
R1282 B.n172 B.n171 10.6151
R1283 B.n172 B.n141 10.6151
R1284 B.n176 B.n141 10.6151
R1285 B.n177 B.n176 10.6151
R1286 B.n178 B.n177 10.6151
R1287 B.n178 B.n139 10.6151
R1288 B.n182 B.n139 10.6151
R1289 B.n183 B.n182 10.6151
R1290 B.n184 B.n183 10.6151
R1291 B.n184 B.n137 10.6151
R1292 B.n188 B.n137 10.6151
R1293 B.n189 B.n188 10.6151
R1294 B.n190 B.n189 10.6151
R1295 B.n190 B.n135 10.6151
R1296 B.n194 B.n135 10.6151
R1297 B.n195 B.n194 10.6151
R1298 B.n196 B.n195 10.6151
R1299 B.n196 B.n133 10.6151
R1300 B.n200 B.n133 10.6151
R1301 B.n201 B.n200 10.6151
R1302 B.n202 B.n201 10.6151
R1303 B.n202 B.n131 10.6151
R1304 B.n206 B.n131 10.6151
R1305 B.n207 B.n206 10.6151
R1306 B.n208 B.n207 10.6151
R1307 B.n208 B.n129 10.6151
R1308 B.n212 B.n129 10.6151
R1309 B.n213 B.n212 10.6151
R1310 B.n214 B.n213 10.6151
R1311 B.n214 B.n127 10.6151
R1312 B.n218 B.n127 10.6151
R1313 B.n219 B.n218 10.6151
R1314 B.n220 B.n219 10.6151
R1315 B.n224 B.n125 10.6151
R1316 B.n225 B.n224 10.6151
R1317 B.n226 B.n225 10.6151
R1318 B.n226 B.n123 10.6151
R1319 B.n230 B.n123 10.6151
R1320 B.n231 B.n230 10.6151
R1321 B.n232 B.n231 10.6151
R1322 B.n232 B.n121 10.6151
R1323 B.n236 B.n121 10.6151
R1324 B.n237 B.n236 10.6151
R1325 B.n238 B.n237 10.6151
R1326 B.n238 B.n119 10.6151
R1327 B.n242 B.n119 10.6151
R1328 B.n243 B.n242 10.6151
R1329 B.n247 B.n243 10.6151
R1330 B.n251 B.n117 10.6151
R1331 B.n252 B.n251 10.6151
R1332 B.n253 B.n252 10.6151
R1333 B.n253 B.n115 10.6151
R1334 B.n257 B.n115 10.6151
R1335 B.n258 B.n257 10.6151
R1336 B.n259 B.n258 10.6151
R1337 B.n259 B.n113 10.6151
R1338 B.n263 B.n113 10.6151
R1339 B.n266 B.n265 10.6151
R1340 B.n266 B.n109 10.6151
R1341 B.n270 B.n109 10.6151
R1342 B.n271 B.n270 10.6151
R1343 B.n272 B.n271 10.6151
R1344 B.n272 B.n107 10.6151
R1345 B.n276 B.n107 10.6151
R1346 B.n277 B.n276 10.6151
R1347 B.n278 B.n277 10.6151
R1348 B.n278 B.n105 10.6151
R1349 B.n282 B.n105 10.6151
R1350 B.n283 B.n282 10.6151
R1351 B.n284 B.n283 10.6151
R1352 B.n284 B.n103 10.6151
R1353 B.n288 B.n103 10.6151
R1354 B.n38 B.n34 9.36635
R1355 B.n463 B.n462 9.36635
R1356 B.n247 B.n246 9.36635
R1357 B.n265 B.n264 9.36635
R1358 B.n577 B.n0 8.11757
R1359 B.n577 B.n1 8.11757
R1360 B.n477 B.n38 1.24928
R1361 B.n464 B.n463 1.24928
R1362 B.n246 B.n117 1.24928
R1363 B.n264 B.n263 1.24928
C0 VDD2 VDD1 1.80213f
C1 VDD1 w_n3802_n1648# 1.96382f
C2 VN VTAIL 4.1983f
C3 VDD1 VP 3.57462f
C4 VN B 1.06254f
C5 B VTAIL 1.59782f
C6 VDD2 w_n3802_n1648# 2.0774f
C7 VDD2 VP 0.515887f
C8 VDD1 VN 0.157161f
C9 VP w_n3802_n1648# 8.28483f
C10 VDD1 VTAIL 5.92706f
C11 VDD1 B 1.58614f
C12 VDD2 VN 3.21886f
C13 VN w_n3802_n1648# 7.793299f
C14 VN VP 5.96498f
C15 VDD2 VTAIL 5.97596f
C16 VTAIL w_n3802_n1648# 1.88447f
C17 VDD2 B 1.68202f
C18 VP VTAIL 4.21248f
C19 B w_n3802_n1648# 7.19829f
C20 VP B 1.88849f
C21 VDD2 VSUBS 1.536774f
C22 VDD1 VSUBS 1.422974f
C23 VTAIL VSUBS 0.515918f
C24 VN VSUBS 6.53222f
C25 VP VSUBS 2.957406f
C26 B VSUBS 3.69944f
C27 w_n3802_n1648# VSUBS 79.1576f
C28 B.n0 VSUBS 0.00649f
C29 B.n1 VSUBS 0.00649f
C30 B.n2 VSUBS 0.009598f
C31 B.n3 VSUBS 0.007355f
C32 B.n4 VSUBS 0.007355f
C33 B.n5 VSUBS 0.007355f
C34 B.n6 VSUBS 0.007355f
C35 B.n7 VSUBS 0.007355f
C36 B.n8 VSUBS 0.007355f
C37 B.n9 VSUBS 0.007355f
C38 B.n10 VSUBS 0.007355f
C39 B.n11 VSUBS 0.007355f
C40 B.n12 VSUBS 0.007355f
C41 B.n13 VSUBS 0.007355f
C42 B.n14 VSUBS 0.007355f
C43 B.n15 VSUBS 0.007355f
C44 B.n16 VSUBS 0.007355f
C45 B.n17 VSUBS 0.007355f
C46 B.n18 VSUBS 0.007355f
C47 B.n19 VSUBS 0.007355f
C48 B.n20 VSUBS 0.007355f
C49 B.n21 VSUBS 0.007355f
C50 B.n22 VSUBS 0.007355f
C51 B.n23 VSUBS 0.007355f
C52 B.n24 VSUBS 0.007355f
C53 B.n25 VSUBS 0.007355f
C54 B.n26 VSUBS 0.01803f
C55 B.n27 VSUBS 0.007355f
C56 B.n28 VSUBS 0.007355f
C57 B.n29 VSUBS 0.007355f
C58 B.n30 VSUBS 0.007355f
C59 B.n31 VSUBS 0.007355f
C60 B.n32 VSUBS 0.007355f
C61 B.n33 VSUBS 0.007355f
C62 B.n34 VSUBS 0.006923f
C63 B.n35 VSUBS 0.007355f
C64 B.t7 VSUBS 0.053099f
C65 B.t8 VSUBS 0.068661f
C66 B.t6 VSUBS 0.348094f
C67 B.n36 VSUBS 0.120389f
C68 B.n37 VSUBS 0.104059f
C69 B.n38 VSUBS 0.017042f
C70 B.n39 VSUBS 0.007355f
C71 B.n40 VSUBS 0.007355f
C72 B.n41 VSUBS 0.007355f
C73 B.n42 VSUBS 0.007355f
C74 B.t4 VSUBS 0.0531f
C75 B.t5 VSUBS 0.068661f
C76 B.t3 VSUBS 0.348094f
C77 B.n43 VSUBS 0.120389f
C78 B.n44 VSUBS 0.104059f
C79 B.n45 VSUBS 0.007355f
C80 B.n46 VSUBS 0.007355f
C81 B.n47 VSUBS 0.007355f
C82 B.n48 VSUBS 0.007355f
C83 B.n49 VSUBS 0.007355f
C84 B.n50 VSUBS 0.007355f
C85 B.n51 VSUBS 0.007355f
C86 B.n52 VSUBS 0.018963f
C87 B.n53 VSUBS 0.007355f
C88 B.n54 VSUBS 0.007355f
C89 B.n55 VSUBS 0.007355f
C90 B.n56 VSUBS 0.007355f
C91 B.n57 VSUBS 0.007355f
C92 B.n58 VSUBS 0.007355f
C93 B.n59 VSUBS 0.007355f
C94 B.n60 VSUBS 0.007355f
C95 B.n61 VSUBS 0.007355f
C96 B.n62 VSUBS 0.007355f
C97 B.n63 VSUBS 0.007355f
C98 B.n64 VSUBS 0.007355f
C99 B.n65 VSUBS 0.007355f
C100 B.n66 VSUBS 0.007355f
C101 B.n67 VSUBS 0.007355f
C102 B.n68 VSUBS 0.007355f
C103 B.n69 VSUBS 0.007355f
C104 B.n70 VSUBS 0.007355f
C105 B.n71 VSUBS 0.007355f
C106 B.n72 VSUBS 0.007355f
C107 B.n73 VSUBS 0.007355f
C108 B.n74 VSUBS 0.007355f
C109 B.n75 VSUBS 0.007355f
C110 B.n76 VSUBS 0.007355f
C111 B.n77 VSUBS 0.007355f
C112 B.n78 VSUBS 0.007355f
C113 B.n79 VSUBS 0.007355f
C114 B.n80 VSUBS 0.007355f
C115 B.n81 VSUBS 0.007355f
C116 B.n82 VSUBS 0.007355f
C117 B.n83 VSUBS 0.007355f
C118 B.n84 VSUBS 0.007355f
C119 B.n85 VSUBS 0.007355f
C120 B.n86 VSUBS 0.007355f
C121 B.n87 VSUBS 0.007355f
C122 B.n88 VSUBS 0.007355f
C123 B.n89 VSUBS 0.007355f
C124 B.n90 VSUBS 0.007355f
C125 B.n91 VSUBS 0.007355f
C126 B.n92 VSUBS 0.007355f
C127 B.n93 VSUBS 0.007355f
C128 B.n94 VSUBS 0.007355f
C129 B.n95 VSUBS 0.007355f
C130 B.n96 VSUBS 0.007355f
C131 B.n97 VSUBS 0.007355f
C132 B.n98 VSUBS 0.007355f
C133 B.n99 VSUBS 0.007355f
C134 B.n100 VSUBS 0.007355f
C135 B.n101 VSUBS 0.007355f
C136 B.n102 VSUBS 0.01803f
C137 B.n103 VSUBS 0.007355f
C138 B.n104 VSUBS 0.007355f
C139 B.n105 VSUBS 0.007355f
C140 B.n106 VSUBS 0.007355f
C141 B.n107 VSUBS 0.007355f
C142 B.n108 VSUBS 0.007355f
C143 B.n109 VSUBS 0.007355f
C144 B.n110 VSUBS 0.007355f
C145 B.t11 VSUBS 0.0531f
C146 B.t10 VSUBS 0.068661f
C147 B.t9 VSUBS 0.348094f
C148 B.n111 VSUBS 0.120389f
C149 B.n112 VSUBS 0.104059f
C150 B.n113 VSUBS 0.007355f
C151 B.n114 VSUBS 0.007355f
C152 B.n115 VSUBS 0.007355f
C153 B.n116 VSUBS 0.007355f
C154 B.n117 VSUBS 0.00411f
C155 B.n118 VSUBS 0.007355f
C156 B.n119 VSUBS 0.007355f
C157 B.n120 VSUBS 0.007355f
C158 B.n121 VSUBS 0.007355f
C159 B.n122 VSUBS 0.007355f
C160 B.n123 VSUBS 0.007355f
C161 B.n124 VSUBS 0.007355f
C162 B.n125 VSUBS 0.018963f
C163 B.n126 VSUBS 0.007355f
C164 B.n127 VSUBS 0.007355f
C165 B.n128 VSUBS 0.007355f
C166 B.n129 VSUBS 0.007355f
C167 B.n130 VSUBS 0.007355f
C168 B.n131 VSUBS 0.007355f
C169 B.n132 VSUBS 0.007355f
C170 B.n133 VSUBS 0.007355f
C171 B.n134 VSUBS 0.007355f
C172 B.n135 VSUBS 0.007355f
C173 B.n136 VSUBS 0.007355f
C174 B.n137 VSUBS 0.007355f
C175 B.n138 VSUBS 0.007355f
C176 B.n139 VSUBS 0.007355f
C177 B.n140 VSUBS 0.007355f
C178 B.n141 VSUBS 0.007355f
C179 B.n142 VSUBS 0.007355f
C180 B.n143 VSUBS 0.007355f
C181 B.n144 VSUBS 0.007355f
C182 B.n145 VSUBS 0.007355f
C183 B.n146 VSUBS 0.007355f
C184 B.n147 VSUBS 0.007355f
C185 B.n148 VSUBS 0.007355f
C186 B.n149 VSUBS 0.007355f
C187 B.n150 VSUBS 0.007355f
C188 B.n151 VSUBS 0.007355f
C189 B.n152 VSUBS 0.007355f
C190 B.n153 VSUBS 0.007355f
C191 B.n154 VSUBS 0.007355f
C192 B.n155 VSUBS 0.007355f
C193 B.n156 VSUBS 0.007355f
C194 B.n157 VSUBS 0.007355f
C195 B.n158 VSUBS 0.007355f
C196 B.n159 VSUBS 0.007355f
C197 B.n160 VSUBS 0.007355f
C198 B.n161 VSUBS 0.007355f
C199 B.n162 VSUBS 0.007355f
C200 B.n163 VSUBS 0.007355f
C201 B.n164 VSUBS 0.007355f
C202 B.n165 VSUBS 0.007355f
C203 B.n166 VSUBS 0.007355f
C204 B.n167 VSUBS 0.007355f
C205 B.n168 VSUBS 0.007355f
C206 B.n169 VSUBS 0.007355f
C207 B.n170 VSUBS 0.007355f
C208 B.n171 VSUBS 0.007355f
C209 B.n172 VSUBS 0.007355f
C210 B.n173 VSUBS 0.007355f
C211 B.n174 VSUBS 0.007355f
C212 B.n175 VSUBS 0.007355f
C213 B.n176 VSUBS 0.007355f
C214 B.n177 VSUBS 0.007355f
C215 B.n178 VSUBS 0.007355f
C216 B.n179 VSUBS 0.007355f
C217 B.n180 VSUBS 0.007355f
C218 B.n181 VSUBS 0.007355f
C219 B.n182 VSUBS 0.007355f
C220 B.n183 VSUBS 0.007355f
C221 B.n184 VSUBS 0.007355f
C222 B.n185 VSUBS 0.007355f
C223 B.n186 VSUBS 0.007355f
C224 B.n187 VSUBS 0.007355f
C225 B.n188 VSUBS 0.007355f
C226 B.n189 VSUBS 0.007355f
C227 B.n190 VSUBS 0.007355f
C228 B.n191 VSUBS 0.007355f
C229 B.n192 VSUBS 0.007355f
C230 B.n193 VSUBS 0.007355f
C231 B.n194 VSUBS 0.007355f
C232 B.n195 VSUBS 0.007355f
C233 B.n196 VSUBS 0.007355f
C234 B.n197 VSUBS 0.007355f
C235 B.n198 VSUBS 0.007355f
C236 B.n199 VSUBS 0.007355f
C237 B.n200 VSUBS 0.007355f
C238 B.n201 VSUBS 0.007355f
C239 B.n202 VSUBS 0.007355f
C240 B.n203 VSUBS 0.007355f
C241 B.n204 VSUBS 0.007355f
C242 B.n205 VSUBS 0.007355f
C243 B.n206 VSUBS 0.007355f
C244 B.n207 VSUBS 0.007355f
C245 B.n208 VSUBS 0.007355f
C246 B.n209 VSUBS 0.007355f
C247 B.n210 VSUBS 0.007355f
C248 B.n211 VSUBS 0.007355f
C249 B.n212 VSUBS 0.007355f
C250 B.n213 VSUBS 0.007355f
C251 B.n214 VSUBS 0.007355f
C252 B.n215 VSUBS 0.007355f
C253 B.n216 VSUBS 0.007355f
C254 B.n217 VSUBS 0.007355f
C255 B.n218 VSUBS 0.007355f
C256 B.n219 VSUBS 0.007355f
C257 B.n220 VSUBS 0.01803f
C258 B.n221 VSUBS 0.01803f
C259 B.n222 VSUBS 0.018963f
C260 B.n223 VSUBS 0.007355f
C261 B.n224 VSUBS 0.007355f
C262 B.n225 VSUBS 0.007355f
C263 B.n226 VSUBS 0.007355f
C264 B.n227 VSUBS 0.007355f
C265 B.n228 VSUBS 0.007355f
C266 B.n229 VSUBS 0.007355f
C267 B.n230 VSUBS 0.007355f
C268 B.n231 VSUBS 0.007355f
C269 B.n232 VSUBS 0.007355f
C270 B.n233 VSUBS 0.007355f
C271 B.n234 VSUBS 0.007355f
C272 B.n235 VSUBS 0.007355f
C273 B.n236 VSUBS 0.007355f
C274 B.n237 VSUBS 0.007355f
C275 B.n238 VSUBS 0.007355f
C276 B.n239 VSUBS 0.007355f
C277 B.n240 VSUBS 0.007355f
C278 B.n241 VSUBS 0.007355f
C279 B.n242 VSUBS 0.007355f
C280 B.n243 VSUBS 0.007355f
C281 B.t2 VSUBS 0.053099f
C282 B.t1 VSUBS 0.068661f
C283 B.t0 VSUBS 0.348094f
C284 B.n244 VSUBS 0.120389f
C285 B.n245 VSUBS 0.104059f
C286 B.n246 VSUBS 0.017042f
C287 B.n247 VSUBS 0.006923f
C288 B.n248 VSUBS 0.007355f
C289 B.n249 VSUBS 0.007355f
C290 B.n250 VSUBS 0.007355f
C291 B.n251 VSUBS 0.007355f
C292 B.n252 VSUBS 0.007355f
C293 B.n253 VSUBS 0.007355f
C294 B.n254 VSUBS 0.007355f
C295 B.n255 VSUBS 0.007355f
C296 B.n256 VSUBS 0.007355f
C297 B.n257 VSUBS 0.007355f
C298 B.n258 VSUBS 0.007355f
C299 B.n259 VSUBS 0.007355f
C300 B.n260 VSUBS 0.007355f
C301 B.n261 VSUBS 0.007355f
C302 B.n262 VSUBS 0.007355f
C303 B.n263 VSUBS 0.00411f
C304 B.n264 VSUBS 0.017042f
C305 B.n265 VSUBS 0.006923f
C306 B.n266 VSUBS 0.007355f
C307 B.n267 VSUBS 0.007355f
C308 B.n268 VSUBS 0.007355f
C309 B.n269 VSUBS 0.007355f
C310 B.n270 VSUBS 0.007355f
C311 B.n271 VSUBS 0.007355f
C312 B.n272 VSUBS 0.007355f
C313 B.n273 VSUBS 0.007355f
C314 B.n274 VSUBS 0.007355f
C315 B.n275 VSUBS 0.007355f
C316 B.n276 VSUBS 0.007355f
C317 B.n277 VSUBS 0.007355f
C318 B.n278 VSUBS 0.007355f
C319 B.n279 VSUBS 0.007355f
C320 B.n280 VSUBS 0.007355f
C321 B.n281 VSUBS 0.007355f
C322 B.n282 VSUBS 0.007355f
C323 B.n283 VSUBS 0.007355f
C324 B.n284 VSUBS 0.007355f
C325 B.n285 VSUBS 0.007355f
C326 B.n286 VSUBS 0.007355f
C327 B.n287 VSUBS 0.018963f
C328 B.n288 VSUBS 0.018183f
C329 B.n289 VSUBS 0.018811f
C330 B.n290 VSUBS 0.007355f
C331 B.n291 VSUBS 0.007355f
C332 B.n292 VSUBS 0.007355f
C333 B.n293 VSUBS 0.007355f
C334 B.n294 VSUBS 0.007355f
C335 B.n295 VSUBS 0.007355f
C336 B.n296 VSUBS 0.007355f
C337 B.n297 VSUBS 0.007355f
C338 B.n298 VSUBS 0.007355f
C339 B.n299 VSUBS 0.007355f
C340 B.n300 VSUBS 0.007355f
C341 B.n301 VSUBS 0.007355f
C342 B.n302 VSUBS 0.007355f
C343 B.n303 VSUBS 0.007355f
C344 B.n304 VSUBS 0.007355f
C345 B.n305 VSUBS 0.007355f
C346 B.n306 VSUBS 0.007355f
C347 B.n307 VSUBS 0.007355f
C348 B.n308 VSUBS 0.007355f
C349 B.n309 VSUBS 0.007355f
C350 B.n310 VSUBS 0.007355f
C351 B.n311 VSUBS 0.007355f
C352 B.n312 VSUBS 0.007355f
C353 B.n313 VSUBS 0.007355f
C354 B.n314 VSUBS 0.007355f
C355 B.n315 VSUBS 0.007355f
C356 B.n316 VSUBS 0.007355f
C357 B.n317 VSUBS 0.007355f
C358 B.n318 VSUBS 0.007355f
C359 B.n319 VSUBS 0.007355f
C360 B.n320 VSUBS 0.007355f
C361 B.n321 VSUBS 0.007355f
C362 B.n322 VSUBS 0.007355f
C363 B.n323 VSUBS 0.007355f
C364 B.n324 VSUBS 0.007355f
C365 B.n325 VSUBS 0.007355f
C366 B.n326 VSUBS 0.007355f
C367 B.n327 VSUBS 0.007355f
C368 B.n328 VSUBS 0.007355f
C369 B.n329 VSUBS 0.007355f
C370 B.n330 VSUBS 0.007355f
C371 B.n331 VSUBS 0.007355f
C372 B.n332 VSUBS 0.007355f
C373 B.n333 VSUBS 0.007355f
C374 B.n334 VSUBS 0.007355f
C375 B.n335 VSUBS 0.007355f
C376 B.n336 VSUBS 0.007355f
C377 B.n337 VSUBS 0.007355f
C378 B.n338 VSUBS 0.007355f
C379 B.n339 VSUBS 0.007355f
C380 B.n340 VSUBS 0.007355f
C381 B.n341 VSUBS 0.007355f
C382 B.n342 VSUBS 0.007355f
C383 B.n343 VSUBS 0.007355f
C384 B.n344 VSUBS 0.007355f
C385 B.n345 VSUBS 0.007355f
C386 B.n346 VSUBS 0.007355f
C387 B.n347 VSUBS 0.007355f
C388 B.n348 VSUBS 0.007355f
C389 B.n349 VSUBS 0.007355f
C390 B.n350 VSUBS 0.007355f
C391 B.n351 VSUBS 0.007355f
C392 B.n352 VSUBS 0.007355f
C393 B.n353 VSUBS 0.007355f
C394 B.n354 VSUBS 0.007355f
C395 B.n355 VSUBS 0.007355f
C396 B.n356 VSUBS 0.007355f
C397 B.n357 VSUBS 0.007355f
C398 B.n358 VSUBS 0.007355f
C399 B.n359 VSUBS 0.007355f
C400 B.n360 VSUBS 0.007355f
C401 B.n361 VSUBS 0.007355f
C402 B.n362 VSUBS 0.007355f
C403 B.n363 VSUBS 0.007355f
C404 B.n364 VSUBS 0.007355f
C405 B.n365 VSUBS 0.007355f
C406 B.n366 VSUBS 0.007355f
C407 B.n367 VSUBS 0.007355f
C408 B.n368 VSUBS 0.007355f
C409 B.n369 VSUBS 0.007355f
C410 B.n370 VSUBS 0.007355f
C411 B.n371 VSUBS 0.007355f
C412 B.n372 VSUBS 0.007355f
C413 B.n373 VSUBS 0.007355f
C414 B.n374 VSUBS 0.007355f
C415 B.n375 VSUBS 0.007355f
C416 B.n376 VSUBS 0.007355f
C417 B.n377 VSUBS 0.007355f
C418 B.n378 VSUBS 0.007355f
C419 B.n379 VSUBS 0.007355f
C420 B.n380 VSUBS 0.007355f
C421 B.n381 VSUBS 0.007355f
C422 B.n382 VSUBS 0.007355f
C423 B.n383 VSUBS 0.007355f
C424 B.n384 VSUBS 0.007355f
C425 B.n385 VSUBS 0.007355f
C426 B.n386 VSUBS 0.007355f
C427 B.n387 VSUBS 0.007355f
C428 B.n388 VSUBS 0.007355f
C429 B.n389 VSUBS 0.007355f
C430 B.n390 VSUBS 0.007355f
C431 B.n391 VSUBS 0.007355f
C432 B.n392 VSUBS 0.007355f
C433 B.n393 VSUBS 0.007355f
C434 B.n394 VSUBS 0.007355f
C435 B.n395 VSUBS 0.007355f
C436 B.n396 VSUBS 0.007355f
C437 B.n397 VSUBS 0.007355f
C438 B.n398 VSUBS 0.007355f
C439 B.n399 VSUBS 0.007355f
C440 B.n400 VSUBS 0.007355f
C441 B.n401 VSUBS 0.007355f
C442 B.n402 VSUBS 0.007355f
C443 B.n403 VSUBS 0.007355f
C444 B.n404 VSUBS 0.007355f
C445 B.n405 VSUBS 0.007355f
C446 B.n406 VSUBS 0.007355f
C447 B.n407 VSUBS 0.007355f
C448 B.n408 VSUBS 0.007355f
C449 B.n409 VSUBS 0.007355f
C450 B.n410 VSUBS 0.007355f
C451 B.n411 VSUBS 0.007355f
C452 B.n412 VSUBS 0.007355f
C453 B.n413 VSUBS 0.007355f
C454 B.n414 VSUBS 0.007355f
C455 B.n415 VSUBS 0.007355f
C456 B.n416 VSUBS 0.007355f
C457 B.n417 VSUBS 0.007355f
C458 B.n418 VSUBS 0.007355f
C459 B.n419 VSUBS 0.007355f
C460 B.n420 VSUBS 0.007355f
C461 B.n421 VSUBS 0.007355f
C462 B.n422 VSUBS 0.007355f
C463 B.n423 VSUBS 0.007355f
C464 B.n424 VSUBS 0.007355f
C465 B.n425 VSUBS 0.007355f
C466 B.n426 VSUBS 0.007355f
C467 B.n427 VSUBS 0.007355f
C468 B.n428 VSUBS 0.007355f
C469 B.n429 VSUBS 0.007355f
C470 B.n430 VSUBS 0.007355f
C471 B.n431 VSUBS 0.007355f
C472 B.n432 VSUBS 0.007355f
C473 B.n433 VSUBS 0.007355f
C474 B.n434 VSUBS 0.007355f
C475 B.n435 VSUBS 0.007355f
C476 B.n436 VSUBS 0.007355f
C477 B.n437 VSUBS 0.01803f
C478 B.n438 VSUBS 0.01803f
C479 B.n439 VSUBS 0.018963f
C480 B.n440 VSUBS 0.007355f
C481 B.n441 VSUBS 0.007355f
C482 B.n442 VSUBS 0.007355f
C483 B.n443 VSUBS 0.007355f
C484 B.n444 VSUBS 0.007355f
C485 B.n445 VSUBS 0.007355f
C486 B.n446 VSUBS 0.007355f
C487 B.n447 VSUBS 0.007355f
C488 B.n448 VSUBS 0.007355f
C489 B.n449 VSUBS 0.007355f
C490 B.n450 VSUBS 0.007355f
C491 B.n451 VSUBS 0.007355f
C492 B.n452 VSUBS 0.007355f
C493 B.n453 VSUBS 0.007355f
C494 B.n454 VSUBS 0.007355f
C495 B.n455 VSUBS 0.007355f
C496 B.n456 VSUBS 0.007355f
C497 B.n457 VSUBS 0.007355f
C498 B.n458 VSUBS 0.007355f
C499 B.n459 VSUBS 0.007355f
C500 B.n460 VSUBS 0.007355f
C501 B.n461 VSUBS 0.007355f
C502 B.n462 VSUBS 0.006923f
C503 B.n463 VSUBS 0.017042f
C504 B.n464 VSUBS 0.00411f
C505 B.n465 VSUBS 0.007355f
C506 B.n466 VSUBS 0.007355f
C507 B.n467 VSUBS 0.007355f
C508 B.n468 VSUBS 0.007355f
C509 B.n469 VSUBS 0.007355f
C510 B.n470 VSUBS 0.007355f
C511 B.n471 VSUBS 0.007355f
C512 B.n472 VSUBS 0.007355f
C513 B.n473 VSUBS 0.007355f
C514 B.n474 VSUBS 0.007355f
C515 B.n475 VSUBS 0.007355f
C516 B.n476 VSUBS 0.007355f
C517 B.n477 VSUBS 0.00411f
C518 B.n478 VSUBS 0.007355f
C519 B.n479 VSUBS 0.007355f
C520 B.n480 VSUBS 0.007355f
C521 B.n481 VSUBS 0.007355f
C522 B.n482 VSUBS 0.007355f
C523 B.n483 VSUBS 0.007355f
C524 B.n484 VSUBS 0.007355f
C525 B.n485 VSUBS 0.007355f
C526 B.n486 VSUBS 0.007355f
C527 B.n487 VSUBS 0.007355f
C528 B.n488 VSUBS 0.007355f
C529 B.n489 VSUBS 0.007355f
C530 B.n490 VSUBS 0.007355f
C531 B.n491 VSUBS 0.007355f
C532 B.n492 VSUBS 0.007355f
C533 B.n493 VSUBS 0.007355f
C534 B.n494 VSUBS 0.007355f
C535 B.n495 VSUBS 0.007355f
C536 B.n496 VSUBS 0.007355f
C537 B.n497 VSUBS 0.007355f
C538 B.n498 VSUBS 0.007355f
C539 B.n499 VSUBS 0.007355f
C540 B.n500 VSUBS 0.007355f
C541 B.n501 VSUBS 0.018963f
C542 B.n502 VSUBS 0.018963f
C543 B.n503 VSUBS 0.01803f
C544 B.n504 VSUBS 0.007355f
C545 B.n505 VSUBS 0.007355f
C546 B.n506 VSUBS 0.007355f
C547 B.n507 VSUBS 0.007355f
C548 B.n508 VSUBS 0.007355f
C549 B.n509 VSUBS 0.007355f
C550 B.n510 VSUBS 0.007355f
C551 B.n511 VSUBS 0.007355f
C552 B.n512 VSUBS 0.007355f
C553 B.n513 VSUBS 0.007355f
C554 B.n514 VSUBS 0.007355f
C555 B.n515 VSUBS 0.007355f
C556 B.n516 VSUBS 0.007355f
C557 B.n517 VSUBS 0.007355f
C558 B.n518 VSUBS 0.007355f
C559 B.n519 VSUBS 0.007355f
C560 B.n520 VSUBS 0.007355f
C561 B.n521 VSUBS 0.007355f
C562 B.n522 VSUBS 0.007355f
C563 B.n523 VSUBS 0.007355f
C564 B.n524 VSUBS 0.007355f
C565 B.n525 VSUBS 0.007355f
C566 B.n526 VSUBS 0.007355f
C567 B.n527 VSUBS 0.007355f
C568 B.n528 VSUBS 0.007355f
C569 B.n529 VSUBS 0.007355f
C570 B.n530 VSUBS 0.007355f
C571 B.n531 VSUBS 0.007355f
C572 B.n532 VSUBS 0.007355f
C573 B.n533 VSUBS 0.007355f
C574 B.n534 VSUBS 0.007355f
C575 B.n535 VSUBS 0.007355f
C576 B.n536 VSUBS 0.007355f
C577 B.n537 VSUBS 0.007355f
C578 B.n538 VSUBS 0.007355f
C579 B.n539 VSUBS 0.007355f
C580 B.n540 VSUBS 0.007355f
C581 B.n541 VSUBS 0.007355f
C582 B.n542 VSUBS 0.007355f
C583 B.n543 VSUBS 0.007355f
C584 B.n544 VSUBS 0.007355f
C585 B.n545 VSUBS 0.007355f
C586 B.n546 VSUBS 0.007355f
C587 B.n547 VSUBS 0.007355f
C588 B.n548 VSUBS 0.007355f
C589 B.n549 VSUBS 0.007355f
C590 B.n550 VSUBS 0.007355f
C591 B.n551 VSUBS 0.007355f
C592 B.n552 VSUBS 0.007355f
C593 B.n553 VSUBS 0.007355f
C594 B.n554 VSUBS 0.007355f
C595 B.n555 VSUBS 0.007355f
C596 B.n556 VSUBS 0.007355f
C597 B.n557 VSUBS 0.007355f
C598 B.n558 VSUBS 0.007355f
C599 B.n559 VSUBS 0.007355f
C600 B.n560 VSUBS 0.007355f
C601 B.n561 VSUBS 0.007355f
C602 B.n562 VSUBS 0.007355f
C603 B.n563 VSUBS 0.007355f
C604 B.n564 VSUBS 0.007355f
C605 B.n565 VSUBS 0.007355f
C606 B.n566 VSUBS 0.007355f
C607 B.n567 VSUBS 0.007355f
C608 B.n568 VSUBS 0.007355f
C609 B.n569 VSUBS 0.007355f
C610 B.n570 VSUBS 0.007355f
C611 B.n571 VSUBS 0.007355f
C612 B.n572 VSUBS 0.007355f
C613 B.n573 VSUBS 0.007355f
C614 B.n574 VSUBS 0.007355f
C615 B.n575 VSUBS 0.009598f
C616 B.n576 VSUBS 0.010225f
C617 B.n577 VSUBS 0.020333f
C618 VDD1.n0 VSUBS 0.026929f
C619 VDD1.n1 VSUBS 0.023509f
C620 VDD1.n2 VSUBS 0.012633f
C621 VDD1.n3 VSUBS 0.022394f
C622 VDD1.n4 VSUBS 0.021946f
C623 VDD1.t6 VSUBS 0.069036f
C624 VDD1.n5 VSUBS 0.095297f
C625 VDD1.n6 VSUBS 0.262777f
C626 VDD1.n7 VSUBS 0.012633f
C627 VDD1.n8 VSUBS 0.013376f
C628 VDD1.n9 VSUBS 0.029859f
C629 VDD1.n10 VSUBS 0.076024f
C630 VDD1.n11 VSUBS 0.013376f
C631 VDD1.n12 VSUBS 0.012633f
C632 VDD1.n13 VSUBS 0.05177f
C633 VDD1.n14 VSUBS 0.06273f
C634 VDD1.t1 VSUBS 0.063163f
C635 VDD1.t8 VSUBS 0.063163f
C636 VDD1.n15 VSUBS 0.334684f
C637 VDD1.n16 VSUBS 0.712946f
C638 VDD1.n17 VSUBS 0.026929f
C639 VDD1.n18 VSUBS 0.023509f
C640 VDD1.n19 VSUBS 0.012633f
C641 VDD1.n20 VSUBS 0.022394f
C642 VDD1.n21 VSUBS 0.021946f
C643 VDD1.t4 VSUBS 0.069036f
C644 VDD1.n22 VSUBS 0.095297f
C645 VDD1.n23 VSUBS 0.262777f
C646 VDD1.n24 VSUBS 0.012633f
C647 VDD1.n25 VSUBS 0.013376f
C648 VDD1.n26 VSUBS 0.029859f
C649 VDD1.n27 VSUBS 0.076024f
C650 VDD1.n28 VSUBS 0.013376f
C651 VDD1.n29 VSUBS 0.012633f
C652 VDD1.n30 VSUBS 0.05177f
C653 VDD1.n31 VSUBS 0.06273f
C654 VDD1.t0 VSUBS 0.063163f
C655 VDD1.t5 VSUBS 0.063163f
C656 VDD1.n32 VSUBS 0.334683f
C657 VDD1.n33 VSUBS 0.705549f
C658 VDD1.t7 VSUBS 0.063163f
C659 VDD1.t3 VSUBS 0.063163f
C660 VDD1.n34 VSUBS 0.341548f
C661 VDD1.n35 VSUBS 2.19999f
C662 VDD1.t2 VSUBS 0.063163f
C663 VDD1.t9 VSUBS 0.063163f
C664 VDD1.n36 VSUBS 0.334684f
C665 VDD1.n37 VSUBS 2.26266f
C666 VP.n0 VSUBS 0.065027f
C667 VP.t6 VSUBS 0.860552f
C668 VP.n1 VSUBS 0.077161f
C669 VP.n2 VSUBS 0.049326f
C670 VP.t2 VSUBS 0.860552f
C671 VP.n3 VSUBS 0.043008f
C672 VP.n4 VSUBS 0.049326f
C673 VP.t4 VSUBS 0.860552f
C674 VP.n5 VSUBS 0.092772f
C675 VP.n6 VSUBS 0.049326f
C676 VP.t9 VSUBS 0.860552f
C677 VP.n7 VSUBS 0.363186f
C678 VP.n8 VSUBS 0.049326f
C679 VP.n9 VSUBS 0.088761f
C680 VP.n10 VSUBS 0.065027f
C681 VP.t0 VSUBS 0.860552f
C682 VP.n11 VSUBS 0.077161f
C683 VP.n12 VSUBS 0.049326f
C684 VP.t7 VSUBS 0.860552f
C685 VP.n13 VSUBS 0.043008f
C686 VP.n14 VSUBS 0.049326f
C687 VP.t1 VSUBS 0.860552f
C688 VP.n15 VSUBS 0.092772f
C689 VP.n16 VSUBS 0.049326f
C690 VP.t8 VSUBS 0.860552f
C691 VP.n17 VSUBS 0.470233f
C692 VP.t3 VSUBS 1.1262f
C693 VP.n18 VSUBS 0.47643f
C694 VP.n19 VSUBS 0.370278f
C695 VP.n20 VSUBS 0.056248f
C696 VP.n21 VSUBS 0.099094f
C697 VP.n22 VSUBS 0.043008f
C698 VP.n23 VSUBS 0.049326f
C699 VP.n24 VSUBS 0.049326f
C700 VP.n25 VSUBS 0.049326f
C701 VP.n26 VSUBS 0.068892f
C702 VP.n27 VSUBS 0.363186f
C703 VP.n28 VSUBS 0.068892f
C704 VP.n29 VSUBS 0.092772f
C705 VP.n30 VSUBS 0.049326f
C706 VP.n31 VSUBS 0.049326f
C707 VP.n32 VSUBS 0.049326f
C708 VP.n33 VSUBS 0.099094f
C709 VP.n34 VSUBS 0.056248f
C710 VP.n35 VSUBS 0.363186f
C711 VP.n36 VSUBS 0.081536f
C712 VP.n37 VSUBS 0.049326f
C713 VP.n38 VSUBS 0.049326f
C714 VP.n39 VSUBS 0.049326f
C715 VP.n40 VSUBS 0.066244f
C716 VP.n41 VSUBS 0.088761f
C717 VP.n42 VSUBS 0.525634f
C718 VP.n43 VSUBS 2.20158f
C719 VP.t5 VSUBS 0.860552f
C720 VP.n44 VSUBS 0.525634f
C721 VP.n45 VSUBS 2.24238f
C722 VP.n46 VSUBS 0.065027f
C723 VP.n47 VSUBS 0.049326f
C724 VP.n48 VSUBS 0.066244f
C725 VP.n49 VSUBS 0.077161f
C726 VP.n50 VSUBS 0.081536f
C727 VP.n51 VSUBS 0.049326f
C728 VP.n52 VSUBS 0.049326f
C729 VP.n53 VSUBS 0.056248f
C730 VP.n54 VSUBS 0.099094f
C731 VP.n55 VSUBS 0.043008f
C732 VP.n56 VSUBS 0.049326f
C733 VP.n57 VSUBS 0.049326f
C734 VP.n58 VSUBS 0.049326f
C735 VP.n59 VSUBS 0.068892f
C736 VP.n60 VSUBS 0.363186f
C737 VP.n61 VSUBS 0.068892f
C738 VP.n62 VSUBS 0.092772f
C739 VP.n63 VSUBS 0.049326f
C740 VP.n64 VSUBS 0.049326f
C741 VP.n65 VSUBS 0.049326f
C742 VP.n66 VSUBS 0.099094f
C743 VP.n67 VSUBS 0.056248f
C744 VP.n68 VSUBS 0.363186f
C745 VP.n69 VSUBS 0.081536f
C746 VP.n70 VSUBS 0.049326f
C747 VP.n71 VSUBS 0.049326f
C748 VP.n72 VSUBS 0.049326f
C749 VP.n73 VSUBS 0.066244f
C750 VP.n74 VSUBS 0.088761f
C751 VP.n75 VSUBS 0.525634f
C752 VP.n76 VSUBS 0.0551f
C753 VTAIL.t10 VSUBS 0.084065f
C754 VTAIL.t16 VSUBS 0.084065f
C755 VTAIL.n0 VSUBS 0.380923f
C756 VTAIL.n1 VSUBS 0.765675f
C757 VTAIL.n2 VSUBS 0.03584f
C758 VTAIL.n3 VSUBS 0.031288f
C759 VTAIL.n4 VSUBS 0.016813f
C760 VTAIL.n5 VSUBS 0.029805f
C761 VTAIL.n6 VSUBS 0.029208f
C762 VTAIL.t3 VSUBS 0.091881f
C763 VTAIL.n7 VSUBS 0.126831f
C764 VTAIL.n8 VSUBS 0.349732f
C765 VTAIL.n9 VSUBS 0.016813f
C766 VTAIL.n10 VSUBS 0.017802f
C767 VTAIL.n11 VSUBS 0.03974f
C768 VTAIL.n12 VSUBS 0.101181f
C769 VTAIL.n13 VSUBS 0.017802f
C770 VTAIL.n14 VSUBS 0.016813f
C771 VTAIL.n15 VSUBS 0.068902f
C772 VTAIL.n16 VSUBS 0.050996f
C773 VTAIL.n17 VSUBS 0.379829f
C774 VTAIL.t2 VSUBS 0.084065f
C775 VTAIL.t7 VSUBS 0.084065f
C776 VTAIL.n18 VSUBS 0.380923f
C777 VTAIL.n19 VSUBS 0.866275f
C778 VTAIL.t5 VSUBS 0.084065f
C779 VTAIL.t4 VSUBS 0.084065f
C780 VTAIL.n20 VSUBS 0.380923f
C781 VTAIL.n21 VSUBS 1.7919f
C782 VTAIL.t13 VSUBS 0.084065f
C783 VTAIL.t17 VSUBS 0.084065f
C784 VTAIL.n22 VSUBS 0.380925f
C785 VTAIL.n23 VSUBS 1.7919f
C786 VTAIL.t12 VSUBS 0.084065f
C787 VTAIL.t18 VSUBS 0.084065f
C788 VTAIL.n24 VSUBS 0.380925f
C789 VTAIL.n25 VSUBS 0.866273f
C790 VTAIL.n26 VSUBS 0.03584f
C791 VTAIL.n27 VSUBS 0.031288f
C792 VTAIL.n28 VSUBS 0.016813f
C793 VTAIL.n29 VSUBS 0.029805f
C794 VTAIL.n30 VSUBS 0.029208f
C795 VTAIL.t14 VSUBS 0.091881f
C796 VTAIL.n31 VSUBS 0.126831f
C797 VTAIL.n32 VSUBS 0.349732f
C798 VTAIL.n33 VSUBS 0.016813f
C799 VTAIL.n34 VSUBS 0.017802f
C800 VTAIL.n35 VSUBS 0.03974f
C801 VTAIL.n36 VSUBS 0.101181f
C802 VTAIL.n37 VSUBS 0.017802f
C803 VTAIL.n38 VSUBS 0.016813f
C804 VTAIL.n39 VSUBS 0.068902f
C805 VTAIL.n40 VSUBS 0.050996f
C806 VTAIL.n41 VSUBS 0.379829f
C807 VTAIL.t0 VSUBS 0.084065f
C808 VTAIL.t8 VSUBS 0.084065f
C809 VTAIL.n42 VSUBS 0.380925f
C810 VTAIL.n43 VSUBS 0.811084f
C811 VTAIL.t6 VSUBS 0.084065f
C812 VTAIL.t9 VSUBS 0.084065f
C813 VTAIL.n44 VSUBS 0.380925f
C814 VTAIL.n45 VSUBS 0.866273f
C815 VTAIL.n46 VSUBS 0.03584f
C816 VTAIL.n47 VSUBS 0.031288f
C817 VTAIL.n48 VSUBS 0.016813f
C818 VTAIL.n49 VSUBS 0.029805f
C819 VTAIL.n50 VSUBS 0.029208f
C820 VTAIL.t1 VSUBS 0.091881f
C821 VTAIL.n51 VSUBS 0.126831f
C822 VTAIL.n52 VSUBS 0.349732f
C823 VTAIL.n53 VSUBS 0.016813f
C824 VTAIL.n54 VSUBS 0.017802f
C825 VTAIL.n55 VSUBS 0.03974f
C826 VTAIL.n56 VSUBS 0.101181f
C827 VTAIL.n57 VSUBS 0.017802f
C828 VTAIL.n58 VSUBS 0.016813f
C829 VTAIL.n59 VSUBS 0.068902f
C830 VTAIL.n60 VSUBS 0.050996f
C831 VTAIL.n61 VSUBS 1.15553f
C832 VTAIL.n62 VSUBS 0.03584f
C833 VTAIL.n63 VSUBS 0.031288f
C834 VTAIL.n64 VSUBS 0.016813f
C835 VTAIL.n65 VSUBS 0.029805f
C836 VTAIL.n66 VSUBS 0.029208f
C837 VTAIL.t11 VSUBS 0.091881f
C838 VTAIL.n67 VSUBS 0.126831f
C839 VTAIL.n68 VSUBS 0.349732f
C840 VTAIL.n69 VSUBS 0.016813f
C841 VTAIL.n70 VSUBS 0.017802f
C842 VTAIL.n71 VSUBS 0.03974f
C843 VTAIL.n72 VSUBS 0.101181f
C844 VTAIL.n73 VSUBS 0.017802f
C845 VTAIL.n74 VSUBS 0.016813f
C846 VTAIL.n75 VSUBS 0.068902f
C847 VTAIL.n76 VSUBS 0.050996f
C848 VTAIL.n77 VSUBS 1.15553f
C849 VTAIL.t15 VSUBS 0.084065f
C850 VTAIL.t19 VSUBS 0.084065f
C851 VTAIL.n78 VSUBS 0.380923f
C852 VTAIL.n79 VSUBS 0.706575f
C853 VDD2.n0 VSUBS 0.032327f
C854 VDD2.n1 VSUBS 0.028221f
C855 VDD2.n2 VSUBS 0.015165f
C856 VDD2.n3 VSUBS 0.026883f
C857 VDD2.n4 VSUBS 0.026345f
C858 VDD2.t1 VSUBS 0.082875f
C859 VDD2.n5 VSUBS 0.114398f
C860 VDD2.n6 VSUBS 0.315449f
C861 VDD2.n7 VSUBS 0.015165f
C862 VDD2.n8 VSUBS 0.016057f
C863 VDD2.n9 VSUBS 0.035844f
C864 VDD2.n10 VSUBS 0.091263f
C865 VDD2.n11 VSUBS 0.016057f
C866 VDD2.n12 VSUBS 0.015165f
C867 VDD2.n13 VSUBS 0.062148f
C868 VDD2.n14 VSUBS 0.075305f
C869 VDD2.t2 VSUBS 0.075824f
C870 VDD2.t7 VSUBS 0.075824f
C871 VDD2.n15 VSUBS 0.401768f
C872 VDD2.n16 VSUBS 0.846973f
C873 VDD2.t5 VSUBS 0.075824f
C874 VDD2.t3 VSUBS 0.075824f
C875 VDD2.n17 VSUBS 0.41001f
C876 VDD2.n18 VSUBS 2.5245f
C877 VDD2.n19 VSUBS 0.032327f
C878 VDD2.n20 VSUBS 0.028221f
C879 VDD2.n21 VSUBS 0.015165f
C880 VDD2.n22 VSUBS 0.026883f
C881 VDD2.n23 VSUBS 0.026345f
C882 VDD2.t6 VSUBS 0.082875f
C883 VDD2.n24 VSUBS 0.114398f
C884 VDD2.n25 VSUBS 0.315449f
C885 VDD2.n26 VSUBS 0.015165f
C886 VDD2.n27 VSUBS 0.016057f
C887 VDD2.n28 VSUBS 0.035844f
C888 VDD2.n29 VSUBS 0.091263f
C889 VDD2.n30 VSUBS 0.016057f
C890 VDD2.n31 VSUBS 0.015165f
C891 VDD2.n32 VSUBS 0.062148f
C892 VDD2.n33 VSUBS 0.065509f
C893 VDD2.n34 VSUBS 2.24466f
C894 VDD2.t0 VSUBS 0.075824f
C895 VDD2.t4 VSUBS 0.075824f
C896 VDD2.n35 VSUBS 0.40177f
C897 VDD2.n36 VSUBS 0.628065f
C898 VDD2.t8 VSUBS 0.075824f
C899 VDD2.t9 VSUBS 0.075824f
C900 VDD2.n37 VSUBS 0.409988f
C901 VN.n0 VSUBS 0.062184f
C902 VN.t8 VSUBS 0.822925f
C903 VN.n1 VSUBS 0.073788f
C904 VN.n2 VSUBS 0.047169f
C905 VN.t0 VSUBS 0.822925f
C906 VN.n3 VSUBS 0.041128f
C907 VN.n4 VSUBS 0.047169f
C908 VN.t4 VSUBS 0.822925f
C909 VN.n5 VSUBS 0.088716f
C910 VN.n6 VSUBS 0.047169f
C911 VN.t3 VSUBS 0.822925f
C912 VN.n7 VSUBS 0.449673f
C913 VN.t9 VSUBS 1.07696f
C914 VN.n8 VSUBS 0.455599f
C915 VN.n9 VSUBS 0.354088f
C916 VN.n10 VSUBS 0.053789f
C917 VN.n11 VSUBS 0.094761f
C918 VN.n12 VSUBS 0.041128f
C919 VN.n13 VSUBS 0.047169f
C920 VN.n14 VSUBS 0.047169f
C921 VN.n15 VSUBS 0.047169f
C922 VN.n16 VSUBS 0.06588f
C923 VN.n17 VSUBS 0.347306f
C924 VN.n18 VSUBS 0.06588f
C925 VN.n19 VSUBS 0.088716f
C926 VN.n20 VSUBS 0.047169f
C927 VN.n21 VSUBS 0.047169f
C928 VN.n22 VSUBS 0.047169f
C929 VN.n23 VSUBS 0.094761f
C930 VN.n24 VSUBS 0.053789f
C931 VN.n25 VSUBS 0.347306f
C932 VN.n26 VSUBS 0.077971f
C933 VN.n27 VSUBS 0.047169f
C934 VN.n28 VSUBS 0.047169f
C935 VN.n29 VSUBS 0.047169f
C936 VN.n30 VSUBS 0.063347f
C937 VN.n31 VSUBS 0.08488f
C938 VN.n32 VSUBS 0.502651f
C939 VN.n33 VSUBS 0.052691f
C940 VN.n34 VSUBS 0.062184f
C941 VN.t6 VSUBS 0.822925f
C942 VN.n35 VSUBS 0.073788f
C943 VN.n36 VSUBS 0.047169f
C944 VN.t2 VSUBS 0.822925f
C945 VN.n37 VSUBS 0.041128f
C946 VN.n38 VSUBS 0.047169f
C947 VN.t7 VSUBS 0.822925f
C948 VN.n39 VSUBS 0.088716f
C949 VN.n40 VSUBS 0.047169f
C950 VN.t1 VSUBS 0.822925f
C951 VN.n41 VSUBS 0.449673f
C952 VN.t5 VSUBS 1.07696f
C953 VN.n42 VSUBS 0.455599f
C954 VN.n43 VSUBS 0.354088f
C955 VN.n44 VSUBS 0.053789f
C956 VN.n45 VSUBS 0.094761f
C957 VN.n46 VSUBS 0.041128f
C958 VN.n47 VSUBS 0.047169f
C959 VN.n48 VSUBS 0.047169f
C960 VN.n49 VSUBS 0.047169f
C961 VN.n50 VSUBS 0.06588f
C962 VN.n51 VSUBS 0.347306f
C963 VN.n52 VSUBS 0.06588f
C964 VN.n53 VSUBS 0.088716f
C965 VN.n54 VSUBS 0.047169f
C966 VN.n55 VSUBS 0.047169f
C967 VN.n56 VSUBS 0.047169f
C968 VN.n57 VSUBS 0.094761f
C969 VN.n58 VSUBS 0.053789f
C970 VN.n59 VSUBS 0.347306f
C971 VN.n60 VSUBS 0.077971f
C972 VN.n61 VSUBS 0.047169f
C973 VN.n62 VSUBS 0.047169f
C974 VN.n63 VSUBS 0.047169f
C975 VN.n64 VSUBS 0.063347f
C976 VN.n65 VSUBS 0.08488f
C977 VN.n66 VSUBS 0.502651f
C978 VN.n67 VSUBS 2.13125f
.ends

