* NGSPICE file created from diff_pair_sample_0860.ext - technology: sky130A

.subckt diff_pair_sample_0860 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VP.t0 VDD1.t5 w_n2860_n2596# sky130_fd_pr__pfet_01v8 ad=1.3431 pd=8.47 as=1.3431 ps=8.47 w=8.14 l=1.56
X1 B.t11 B.t9 B.t10 w_n2860_n2596# sky130_fd_pr__pfet_01v8 ad=3.1746 pd=17.06 as=0 ps=0 w=8.14 l=1.56
X2 VDD1.t7 VP.t1 VTAIL.t14 w_n2860_n2596# sky130_fd_pr__pfet_01v8 ad=1.3431 pd=8.47 as=3.1746 ps=17.06 w=8.14 l=1.56
X3 VDD2.t7 VN.t0 VTAIL.t6 w_n2860_n2596# sky130_fd_pr__pfet_01v8 ad=1.3431 pd=8.47 as=1.3431 ps=8.47 w=8.14 l=1.56
X4 VTAIL.t0 VN.t1 VDD2.t6 w_n2860_n2596# sky130_fd_pr__pfet_01v8 ad=1.3431 pd=8.47 as=1.3431 ps=8.47 w=8.14 l=1.56
X5 VTAIL.t7 VN.t2 VDD2.t5 w_n2860_n2596# sky130_fd_pr__pfet_01v8 ad=3.1746 pd=17.06 as=1.3431 ps=8.47 w=8.14 l=1.56
X6 VTAIL.t13 VP.t2 VDD1.t6 w_n2860_n2596# sky130_fd_pr__pfet_01v8 ad=3.1746 pd=17.06 as=1.3431 ps=8.47 w=8.14 l=1.56
X7 VDD2.t4 VN.t3 VTAIL.t1 w_n2860_n2596# sky130_fd_pr__pfet_01v8 ad=1.3431 pd=8.47 as=1.3431 ps=8.47 w=8.14 l=1.56
X8 VDD1.t4 VP.t3 VTAIL.t12 w_n2860_n2596# sky130_fd_pr__pfet_01v8 ad=1.3431 pd=8.47 as=3.1746 ps=17.06 w=8.14 l=1.56
X9 B.t8 B.t6 B.t7 w_n2860_n2596# sky130_fd_pr__pfet_01v8 ad=3.1746 pd=17.06 as=0 ps=0 w=8.14 l=1.56
X10 VTAIL.t4 VN.t4 VDD2.t3 w_n2860_n2596# sky130_fd_pr__pfet_01v8 ad=1.3431 pd=8.47 as=1.3431 ps=8.47 w=8.14 l=1.56
X11 VTAIL.t11 VP.t4 VDD1.t3 w_n2860_n2596# sky130_fd_pr__pfet_01v8 ad=1.3431 pd=8.47 as=1.3431 ps=8.47 w=8.14 l=1.56
X12 VDD2.t2 VN.t5 VTAIL.t5 w_n2860_n2596# sky130_fd_pr__pfet_01v8 ad=1.3431 pd=8.47 as=3.1746 ps=17.06 w=8.14 l=1.56
X13 VDD1.t1 VP.t5 VTAIL.t10 w_n2860_n2596# sky130_fd_pr__pfet_01v8 ad=1.3431 pd=8.47 as=1.3431 ps=8.47 w=8.14 l=1.56
X14 VTAIL.t2 VN.t6 VDD2.t1 w_n2860_n2596# sky130_fd_pr__pfet_01v8 ad=3.1746 pd=17.06 as=1.3431 ps=8.47 w=8.14 l=1.56
X15 VTAIL.t9 VP.t6 VDD1.t0 w_n2860_n2596# sky130_fd_pr__pfet_01v8 ad=3.1746 pd=17.06 as=1.3431 ps=8.47 w=8.14 l=1.56
X16 VDD2.t0 VN.t7 VTAIL.t3 w_n2860_n2596# sky130_fd_pr__pfet_01v8 ad=1.3431 pd=8.47 as=3.1746 ps=17.06 w=8.14 l=1.56
X17 VDD1.t2 VP.t7 VTAIL.t8 w_n2860_n2596# sky130_fd_pr__pfet_01v8 ad=1.3431 pd=8.47 as=1.3431 ps=8.47 w=8.14 l=1.56
X18 B.t5 B.t3 B.t4 w_n2860_n2596# sky130_fd_pr__pfet_01v8 ad=3.1746 pd=17.06 as=0 ps=0 w=8.14 l=1.56
X19 B.t2 B.t0 B.t1 w_n2860_n2596# sky130_fd_pr__pfet_01v8 ad=3.1746 pd=17.06 as=0 ps=0 w=8.14 l=1.56
R0 VP.n28 VP.n27 181.506
R1 VP.n50 VP.n49 181.506
R2 VP.n26 VP.n25 181.506
R3 VP.n13 VP.n12 161.3
R4 VP.n14 VP.n9 161.3
R5 VP.n16 VP.n15 161.3
R6 VP.n17 VP.n8 161.3
R7 VP.n20 VP.n19 161.3
R8 VP.n21 VP.n7 161.3
R9 VP.n23 VP.n22 161.3
R10 VP.n24 VP.n6 161.3
R11 VP.n48 VP.n0 161.3
R12 VP.n47 VP.n46 161.3
R13 VP.n45 VP.n1 161.3
R14 VP.n44 VP.n43 161.3
R15 VP.n41 VP.n2 161.3
R16 VP.n40 VP.n39 161.3
R17 VP.n38 VP.n3 161.3
R18 VP.n37 VP.n36 161.3
R19 VP.n34 VP.n4 161.3
R20 VP.n33 VP.n32 161.3
R21 VP.n31 VP.n5 161.3
R22 VP.n30 VP.n29 161.3
R23 VP.n10 VP.t6 156.085
R24 VP.n28 VP.t2 125.754
R25 VP.n35 VP.t7 125.754
R26 VP.n42 VP.t0 125.754
R27 VP.n49 VP.t3 125.754
R28 VP.n25 VP.t1 125.754
R29 VP.n18 VP.t4 125.754
R30 VP.n11 VP.t5 125.754
R31 VP.n11 VP.n10 56.704
R32 VP.n40 VP.n3 56.4773
R33 VP.n16 VP.n9 56.4773
R34 VP.n33 VP.n5 54.0429
R35 VP.n47 VP.n1 54.0429
R36 VP.n23 VP.n7 54.0429
R37 VP.n27 VP.n26 42.955
R38 VP.n34 VP.n33 26.7783
R39 VP.n43 VP.n1 26.7783
R40 VP.n19 VP.n7 26.7783
R41 VP.n29 VP.n5 24.3439
R42 VP.n36 VP.n3 24.3439
R43 VP.n41 VP.n40 24.3439
R44 VP.n48 VP.n47 24.3439
R45 VP.n24 VP.n23 24.3439
R46 VP.n17 VP.n16 24.3439
R47 VP.n12 VP.n9 24.3439
R48 VP.n13 VP.n10 18.4239
R49 VP.n35 VP.n34 14.85
R50 VP.n43 VP.n42 14.85
R51 VP.n19 VP.n18 14.85
R52 VP.n36 VP.n35 9.49444
R53 VP.n42 VP.n41 9.49444
R54 VP.n18 VP.n17 9.49444
R55 VP.n12 VP.n11 9.49444
R56 VP.n29 VP.n28 4.13888
R57 VP.n49 VP.n48 4.13888
R58 VP.n25 VP.n24 4.13888
R59 VP.n14 VP.n13 0.189894
R60 VP.n15 VP.n14 0.189894
R61 VP.n15 VP.n8 0.189894
R62 VP.n20 VP.n8 0.189894
R63 VP.n21 VP.n20 0.189894
R64 VP.n22 VP.n21 0.189894
R65 VP.n22 VP.n6 0.189894
R66 VP.n26 VP.n6 0.189894
R67 VP.n30 VP.n27 0.189894
R68 VP.n31 VP.n30 0.189894
R69 VP.n32 VP.n31 0.189894
R70 VP.n32 VP.n4 0.189894
R71 VP.n37 VP.n4 0.189894
R72 VP.n38 VP.n37 0.189894
R73 VP.n39 VP.n38 0.189894
R74 VP.n39 VP.n2 0.189894
R75 VP.n44 VP.n2 0.189894
R76 VP.n45 VP.n44 0.189894
R77 VP.n46 VP.n45 0.189894
R78 VP.n46 VP.n0 0.189894
R79 VP.n50 VP.n0 0.189894
R80 VP VP.n50 0.0516364
R81 VDD1 VDD1.n0 83.2719
R82 VDD1.n3 VDD1.n2 83.1582
R83 VDD1.n3 VDD1.n1 83.1582
R84 VDD1.n5 VDD1.n4 82.3991
R85 VDD1.n5 VDD1.n3 38.6474
R86 VDD1.n4 VDD1.t3 3.99374
R87 VDD1.n4 VDD1.t7 3.99374
R88 VDD1.n0 VDD1.t0 3.99374
R89 VDD1.n0 VDD1.t1 3.99374
R90 VDD1.n2 VDD1.t5 3.99374
R91 VDD1.n2 VDD1.t4 3.99374
R92 VDD1.n1 VDD1.t6 3.99374
R93 VDD1.n1 VDD1.t2 3.99374
R94 VDD1 VDD1.n5 0.756965
R95 VTAIL.n354 VTAIL.n316 756.745
R96 VTAIL.n40 VTAIL.n2 756.745
R97 VTAIL.n84 VTAIL.n46 756.745
R98 VTAIL.n130 VTAIL.n92 756.745
R99 VTAIL.n310 VTAIL.n272 756.745
R100 VTAIL.n264 VTAIL.n226 756.745
R101 VTAIL.n220 VTAIL.n182 756.745
R102 VTAIL.n174 VTAIL.n136 756.745
R103 VTAIL.n331 VTAIL.n330 585
R104 VTAIL.n328 VTAIL.n327 585
R105 VTAIL.n337 VTAIL.n336 585
R106 VTAIL.n339 VTAIL.n338 585
R107 VTAIL.n324 VTAIL.n323 585
R108 VTAIL.n345 VTAIL.n344 585
R109 VTAIL.n347 VTAIL.n346 585
R110 VTAIL.n320 VTAIL.n319 585
R111 VTAIL.n353 VTAIL.n352 585
R112 VTAIL.n355 VTAIL.n354 585
R113 VTAIL.n17 VTAIL.n16 585
R114 VTAIL.n14 VTAIL.n13 585
R115 VTAIL.n23 VTAIL.n22 585
R116 VTAIL.n25 VTAIL.n24 585
R117 VTAIL.n10 VTAIL.n9 585
R118 VTAIL.n31 VTAIL.n30 585
R119 VTAIL.n33 VTAIL.n32 585
R120 VTAIL.n6 VTAIL.n5 585
R121 VTAIL.n39 VTAIL.n38 585
R122 VTAIL.n41 VTAIL.n40 585
R123 VTAIL.n61 VTAIL.n60 585
R124 VTAIL.n58 VTAIL.n57 585
R125 VTAIL.n67 VTAIL.n66 585
R126 VTAIL.n69 VTAIL.n68 585
R127 VTAIL.n54 VTAIL.n53 585
R128 VTAIL.n75 VTAIL.n74 585
R129 VTAIL.n77 VTAIL.n76 585
R130 VTAIL.n50 VTAIL.n49 585
R131 VTAIL.n83 VTAIL.n82 585
R132 VTAIL.n85 VTAIL.n84 585
R133 VTAIL.n107 VTAIL.n106 585
R134 VTAIL.n104 VTAIL.n103 585
R135 VTAIL.n113 VTAIL.n112 585
R136 VTAIL.n115 VTAIL.n114 585
R137 VTAIL.n100 VTAIL.n99 585
R138 VTAIL.n121 VTAIL.n120 585
R139 VTAIL.n123 VTAIL.n122 585
R140 VTAIL.n96 VTAIL.n95 585
R141 VTAIL.n129 VTAIL.n128 585
R142 VTAIL.n131 VTAIL.n130 585
R143 VTAIL.n311 VTAIL.n310 585
R144 VTAIL.n309 VTAIL.n308 585
R145 VTAIL.n276 VTAIL.n275 585
R146 VTAIL.n303 VTAIL.n302 585
R147 VTAIL.n301 VTAIL.n300 585
R148 VTAIL.n280 VTAIL.n279 585
R149 VTAIL.n295 VTAIL.n294 585
R150 VTAIL.n293 VTAIL.n292 585
R151 VTAIL.n284 VTAIL.n283 585
R152 VTAIL.n287 VTAIL.n286 585
R153 VTAIL.n265 VTAIL.n264 585
R154 VTAIL.n263 VTAIL.n262 585
R155 VTAIL.n230 VTAIL.n229 585
R156 VTAIL.n257 VTAIL.n256 585
R157 VTAIL.n255 VTAIL.n254 585
R158 VTAIL.n234 VTAIL.n233 585
R159 VTAIL.n249 VTAIL.n248 585
R160 VTAIL.n247 VTAIL.n246 585
R161 VTAIL.n238 VTAIL.n237 585
R162 VTAIL.n241 VTAIL.n240 585
R163 VTAIL.n221 VTAIL.n220 585
R164 VTAIL.n219 VTAIL.n218 585
R165 VTAIL.n186 VTAIL.n185 585
R166 VTAIL.n213 VTAIL.n212 585
R167 VTAIL.n211 VTAIL.n210 585
R168 VTAIL.n190 VTAIL.n189 585
R169 VTAIL.n205 VTAIL.n204 585
R170 VTAIL.n203 VTAIL.n202 585
R171 VTAIL.n194 VTAIL.n193 585
R172 VTAIL.n197 VTAIL.n196 585
R173 VTAIL.n175 VTAIL.n174 585
R174 VTAIL.n173 VTAIL.n172 585
R175 VTAIL.n140 VTAIL.n139 585
R176 VTAIL.n167 VTAIL.n166 585
R177 VTAIL.n165 VTAIL.n164 585
R178 VTAIL.n144 VTAIL.n143 585
R179 VTAIL.n159 VTAIL.n158 585
R180 VTAIL.n157 VTAIL.n156 585
R181 VTAIL.n148 VTAIL.n147 585
R182 VTAIL.n151 VTAIL.n150 585
R183 VTAIL.t3 VTAIL.n329 327.473
R184 VTAIL.t2 VTAIL.n15 327.473
R185 VTAIL.t12 VTAIL.n59 327.473
R186 VTAIL.t13 VTAIL.n105 327.473
R187 VTAIL.t14 VTAIL.n285 327.473
R188 VTAIL.t9 VTAIL.n239 327.473
R189 VTAIL.t5 VTAIL.n195 327.473
R190 VTAIL.t7 VTAIL.n149 327.473
R191 VTAIL.n330 VTAIL.n327 171.744
R192 VTAIL.n337 VTAIL.n327 171.744
R193 VTAIL.n338 VTAIL.n337 171.744
R194 VTAIL.n338 VTAIL.n323 171.744
R195 VTAIL.n345 VTAIL.n323 171.744
R196 VTAIL.n346 VTAIL.n345 171.744
R197 VTAIL.n346 VTAIL.n319 171.744
R198 VTAIL.n353 VTAIL.n319 171.744
R199 VTAIL.n354 VTAIL.n353 171.744
R200 VTAIL.n16 VTAIL.n13 171.744
R201 VTAIL.n23 VTAIL.n13 171.744
R202 VTAIL.n24 VTAIL.n23 171.744
R203 VTAIL.n24 VTAIL.n9 171.744
R204 VTAIL.n31 VTAIL.n9 171.744
R205 VTAIL.n32 VTAIL.n31 171.744
R206 VTAIL.n32 VTAIL.n5 171.744
R207 VTAIL.n39 VTAIL.n5 171.744
R208 VTAIL.n40 VTAIL.n39 171.744
R209 VTAIL.n60 VTAIL.n57 171.744
R210 VTAIL.n67 VTAIL.n57 171.744
R211 VTAIL.n68 VTAIL.n67 171.744
R212 VTAIL.n68 VTAIL.n53 171.744
R213 VTAIL.n75 VTAIL.n53 171.744
R214 VTAIL.n76 VTAIL.n75 171.744
R215 VTAIL.n76 VTAIL.n49 171.744
R216 VTAIL.n83 VTAIL.n49 171.744
R217 VTAIL.n84 VTAIL.n83 171.744
R218 VTAIL.n106 VTAIL.n103 171.744
R219 VTAIL.n113 VTAIL.n103 171.744
R220 VTAIL.n114 VTAIL.n113 171.744
R221 VTAIL.n114 VTAIL.n99 171.744
R222 VTAIL.n121 VTAIL.n99 171.744
R223 VTAIL.n122 VTAIL.n121 171.744
R224 VTAIL.n122 VTAIL.n95 171.744
R225 VTAIL.n129 VTAIL.n95 171.744
R226 VTAIL.n130 VTAIL.n129 171.744
R227 VTAIL.n310 VTAIL.n309 171.744
R228 VTAIL.n309 VTAIL.n275 171.744
R229 VTAIL.n302 VTAIL.n275 171.744
R230 VTAIL.n302 VTAIL.n301 171.744
R231 VTAIL.n301 VTAIL.n279 171.744
R232 VTAIL.n294 VTAIL.n279 171.744
R233 VTAIL.n294 VTAIL.n293 171.744
R234 VTAIL.n293 VTAIL.n283 171.744
R235 VTAIL.n286 VTAIL.n283 171.744
R236 VTAIL.n264 VTAIL.n263 171.744
R237 VTAIL.n263 VTAIL.n229 171.744
R238 VTAIL.n256 VTAIL.n229 171.744
R239 VTAIL.n256 VTAIL.n255 171.744
R240 VTAIL.n255 VTAIL.n233 171.744
R241 VTAIL.n248 VTAIL.n233 171.744
R242 VTAIL.n248 VTAIL.n247 171.744
R243 VTAIL.n247 VTAIL.n237 171.744
R244 VTAIL.n240 VTAIL.n237 171.744
R245 VTAIL.n220 VTAIL.n219 171.744
R246 VTAIL.n219 VTAIL.n185 171.744
R247 VTAIL.n212 VTAIL.n185 171.744
R248 VTAIL.n212 VTAIL.n211 171.744
R249 VTAIL.n211 VTAIL.n189 171.744
R250 VTAIL.n204 VTAIL.n189 171.744
R251 VTAIL.n204 VTAIL.n203 171.744
R252 VTAIL.n203 VTAIL.n193 171.744
R253 VTAIL.n196 VTAIL.n193 171.744
R254 VTAIL.n174 VTAIL.n173 171.744
R255 VTAIL.n173 VTAIL.n139 171.744
R256 VTAIL.n166 VTAIL.n139 171.744
R257 VTAIL.n166 VTAIL.n165 171.744
R258 VTAIL.n165 VTAIL.n143 171.744
R259 VTAIL.n158 VTAIL.n143 171.744
R260 VTAIL.n158 VTAIL.n157 171.744
R261 VTAIL.n157 VTAIL.n147 171.744
R262 VTAIL.n150 VTAIL.n147 171.744
R263 VTAIL.n330 VTAIL.t3 85.8723
R264 VTAIL.n16 VTAIL.t2 85.8723
R265 VTAIL.n60 VTAIL.t12 85.8723
R266 VTAIL.n106 VTAIL.t13 85.8723
R267 VTAIL.n286 VTAIL.t14 85.8723
R268 VTAIL.n240 VTAIL.t9 85.8723
R269 VTAIL.n196 VTAIL.t5 85.8723
R270 VTAIL.n150 VTAIL.t7 85.8723
R271 VTAIL.n271 VTAIL.n270 65.7203
R272 VTAIL.n181 VTAIL.n180 65.7203
R273 VTAIL.n1 VTAIL.n0 65.7201
R274 VTAIL.n91 VTAIL.n90 65.7201
R275 VTAIL.n359 VTAIL.n358 31.7975
R276 VTAIL.n45 VTAIL.n44 31.7975
R277 VTAIL.n89 VTAIL.n88 31.7975
R278 VTAIL.n135 VTAIL.n134 31.7975
R279 VTAIL.n315 VTAIL.n314 31.7975
R280 VTAIL.n269 VTAIL.n268 31.7975
R281 VTAIL.n225 VTAIL.n224 31.7975
R282 VTAIL.n179 VTAIL.n178 31.7975
R283 VTAIL.n359 VTAIL.n315 21.0134
R284 VTAIL.n179 VTAIL.n135 21.0134
R285 VTAIL.n331 VTAIL.n329 16.3894
R286 VTAIL.n17 VTAIL.n15 16.3894
R287 VTAIL.n61 VTAIL.n59 16.3894
R288 VTAIL.n107 VTAIL.n105 16.3894
R289 VTAIL.n287 VTAIL.n285 16.3894
R290 VTAIL.n241 VTAIL.n239 16.3894
R291 VTAIL.n197 VTAIL.n195 16.3894
R292 VTAIL.n151 VTAIL.n149 16.3894
R293 VTAIL.n332 VTAIL.n328 12.8005
R294 VTAIL.n18 VTAIL.n14 12.8005
R295 VTAIL.n62 VTAIL.n58 12.8005
R296 VTAIL.n108 VTAIL.n104 12.8005
R297 VTAIL.n288 VTAIL.n284 12.8005
R298 VTAIL.n242 VTAIL.n238 12.8005
R299 VTAIL.n198 VTAIL.n194 12.8005
R300 VTAIL.n152 VTAIL.n148 12.8005
R301 VTAIL.n336 VTAIL.n335 12.0247
R302 VTAIL.n22 VTAIL.n21 12.0247
R303 VTAIL.n66 VTAIL.n65 12.0247
R304 VTAIL.n112 VTAIL.n111 12.0247
R305 VTAIL.n292 VTAIL.n291 12.0247
R306 VTAIL.n246 VTAIL.n245 12.0247
R307 VTAIL.n202 VTAIL.n201 12.0247
R308 VTAIL.n156 VTAIL.n155 12.0247
R309 VTAIL.n339 VTAIL.n326 11.249
R310 VTAIL.n25 VTAIL.n12 11.249
R311 VTAIL.n69 VTAIL.n56 11.249
R312 VTAIL.n115 VTAIL.n102 11.249
R313 VTAIL.n295 VTAIL.n282 11.249
R314 VTAIL.n249 VTAIL.n236 11.249
R315 VTAIL.n205 VTAIL.n192 11.249
R316 VTAIL.n159 VTAIL.n146 11.249
R317 VTAIL.n340 VTAIL.n324 10.4732
R318 VTAIL.n26 VTAIL.n10 10.4732
R319 VTAIL.n70 VTAIL.n54 10.4732
R320 VTAIL.n116 VTAIL.n100 10.4732
R321 VTAIL.n296 VTAIL.n280 10.4732
R322 VTAIL.n250 VTAIL.n234 10.4732
R323 VTAIL.n206 VTAIL.n190 10.4732
R324 VTAIL.n160 VTAIL.n144 10.4732
R325 VTAIL.n344 VTAIL.n343 9.69747
R326 VTAIL.n30 VTAIL.n29 9.69747
R327 VTAIL.n74 VTAIL.n73 9.69747
R328 VTAIL.n120 VTAIL.n119 9.69747
R329 VTAIL.n300 VTAIL.n299 9.69747
R330 VTAIL.n254 VTAIL.n253 9.69747
R331 VTAIL.n210 VTAIL.n209 9.69747
R332 VTAIL.n164 VTAIL.n163 9.69747
R333 VTAIL.n358 VTAIL.n357 9.45567
R334 VTAIL.n44 VTAIL.n43 9.45567
R335 VTAIL.n88 VTAIL.n87 9.45567
R336 VTAIL.n134 VTAIL.n133 9.45567
R337 VTAIL.n314 VTAIL.n313 9.45567
R338 VTAIL.n268 VTAIL.n267 9.45567
R339 VTAIL.n224 VTAIL.n223 9.45567
R340 VTAIL.n178 VTAIL.n177 9.45567
R341 VTAIL.n318 VTAIL.n317 9.3005
R342 VTAIL.n357 VTAIL.n356 9.3005
R343 VTAIL.n349 VTAIL.n348 9.3005
R344 VTAIL.n322 VTAIL.n321 9.3005
R345 VTAIL.n343 VTAIL.n342 9.3005
R346 VTAIL.n341 VTAIL.n340 9.3005
R347 VTAIL.n326 VTAIL.n325 9.3005
R348 VTAIL.n335 VTAIL.n334 9.3005
R349 VTAIL.n333 VTAIL.n332 9.3005
R350 VTAIL.n351 VTAIL.n350 9.3005
R351 VTAIL.n4 VTAIL.n3 9.3005
R352 VTAIL.n43 VTAIL.n42 9.3005
R353 VTAIL.n35 VTAIL.n34 9.3005
R354 VTAIL.n8 VTAIL.n7 9.3005
R355 VTAIL.n29 VTAIL.n28 9.3005
R356 VTAIL.n27 VTAIL.n26 9.3005
R357 VTAIL.n12 VTAIL.n11 9.3005
R358 VTAIL.n21 VTAIL.n20 9.3005
R359 VTAIL.n19 VTAIL.n18 9.3005
R360 VTAIL.n37 VTAIL.n36 9.3005
R361 VTAIL.n48 VTAIL.n47 9.3005
R362 VTAIL.n87 VTAIL.n86 9.3005
R363 VTAIL.n79 VTAIL.n78 9.3005
R364 VTAIL.n52 VTAIL.n51 9.3005
R365 VTAIL.n73 VTAIL.n72 9.3005
R366 VTAIL.n71 VTAIL.n70 9.3005
R367 VTAIL.n56 VTAIL.n55 9.3005
R368 VTAIL.n65 VTAIL.n64 9.3005
R369 VTAIL.n63 VTAIL.n62 9.3005
R370 VTAIL.n81 VTAIL.n80 9.3005
R371 VTAIL.n94 VTAIL.n93 9.3005
R372 VTAIL.n133 VTAIL.n132 9.3005
R373 VTAIL.n125 VTAIL.n124 9.3005
R374 VTAIL.n98 VTAIL.n97 9.3005
R375 VTAIL.n119 VTAIL.n118 9.3005
R376 VTAIL.n117 VTAIL.n116 9.3005
R377 VTAIL.n102 VTAIL.n101 9.3005
R378 VTAIL.n111 VTAIL.n110 9.3005
R379 VTAIL.n109 VTAIL.n108 9.3005
R380 VTAIL.n127 VTAIL.n126 9.3005
R381 VTAIL.n274 VTAIL.n273 9.3005
R382 VTAIL.n307 VTAIL.n306 9.3005
R383 VTAIL.n305 VTAIL.n304 9.3005
R384 VTAIL.n278 VTAIL.n277 9.3005
R385 VTAIL.n299 VTAIL.n298 9.3005
R386 VTAIL.n297 VTAIL.n296 9.3005
R387 VTAIL.n282 VTAIL.n281 9.3005
R388 VTAIL.n291 VTAIL.n290 9.3005
R389 VTAIL.n289 VTAIL.n288 9.3005
R390 VTAIL.n313 VTAIL.n312 9.3005
R391 VTAIL.n267 VTAIL.n266 9.3005
R392 VTAIL.n228 VTAIL.n227 9.3005
R393 VTAIL.n261 VTAIL.n260 9.3005
R394 VTAIL.n259 VTAIL.n258 9.3005
R395 VTAIL.n232 VTAIL.n231 9.3005
R396 VTAIL.n253 VTAIL.n252 9.3005
R397 VTAIL.n251 VTAIL.n250 9.3005
R398 VTAIL.n236 VTAIL.n235 9.3005
R399 VTAIL.n245 VTAIL.n244 9.3005
R400 VTAIL.n243 VTAIL.n242 9.3005
R401 VTAIL.n223 VTAIL.n222 9.3005
R402 VTAIL.n184 VTAIL.n183 9.3005
R403 VTAIL.n217 VTAIL.n216 9.3005
R404 VTAIL.n215 VTAIL.n214 9.3005
R405 VTAIL.n188 VTAIL.n187 9.3005
R406 VTAIL.n209 VTAIL.n208 9.3005
R407 VTAIL.n207 VTAIL.n206 9.3005
R408 VTAIL.n192 VTAIL.n191 9.3005
R409 VTAIL.n201 VTAIL.n200 9.3005
R410 VTAIL.n199 VTAIL.n198 9.3005
R411 VTAIL.n177 VTAIL.n176 9.3005
R412 VTAIL.n138 VTAIL.n137 9.3005
R413 VTAIL.n171 VTAIL.n170 9.3005
R414 VTAIL.n169 VTAIL.n168 9.3005
R415 VTAIL.n142 VTAIL.n141 9.3005
R416 VTAIL.n163 VTAIL.n162 9.3005
R417 VTAIL.n161 VTAIL.n160 9.3005
R418 VTAIL.n146 VTAIL.n145 9.3005
R419 VTAIL.n155 VTAIL.n154 9.3005
R420 VTAIL.n153 VTAIL.n152 9.3005
R421 VTAIL.n347 VTAIL.n322 8.92171
R422 VTAIL.n33 VTAIL.n8 8.92171
R423 VTAIL.n77 VTAIL.n52 8.92171
R424 VTAIL.n123 VTAIL.n98 8.92171
R425 VTAIL.n303 VTAIL.n278 8.92171
R426 VTAIL.n257 VTAIL.n232 8.92171
R427 VTAIL.n213 VTAIL.n188 8.92171
R428 VTAIL.n167 VTAIL.n142 8.92171
R429 VTAIL.n348 VTAIL.n320 8.14595
R430 VTAIL.n358 VTAIL.n316 8.14595
R431 VTAIL.n34 VTAIL.n6 8.14595
R432 VTAIL.n44 VTAIL.n2 8.14595
R433 VTAIL.n78 VTAIL.n50 8.14595
R434 VTAIL.n88 VTAIL.n46 8.14595
R435 VTAIL.n124 VTAIL.n96 8.14595
R436 VTAIL.n134 VTAIL.n92 8.14595
R437 VTAIL.n314 VTAIL.n272 8.14595
R438 VTAIL.n304 VTAIL.n276 8.14595
R439 VTAIL.n268 VTAIL.n226 8.14595
R440 VTAIL.n258 VTAIL.n230 8.14595
R441 VTAIL.n224 VTAIL.n182 8.14595
R442 VTAIL.n214 VTAIL.n186 8.14595
R443 VTAIL.n178 VTAIL.n136 8.14595
R444 VTAIL.n168 VTAIL.n140 8.14595
R445 VTAIL.n352 VTAIL.n351 7.3702
R446 VTAIL.n356 VTAIL.n355 7.3702
R447 VTAIL.n38 VTAIL.n37 7.3702
R448 VTAIL.n42 VTAIL.n41 7.3702
R449 VTAIL.n82 VTAIL.n81 7.3702
R450 VTAIL.n86 VTAIL.n85 7.3702
R451 VTAIL.n128 VTAIL.n127 7.3702
R452 VTAIL.n132 VTAIL.n131 7.3702
R453 VTAIL.n312 VTAIL.n311 7.3702
R454 VTAIL.n308 VTAIL.n307 7.3702
R455 VTAIL.n266 VTAIL.n265 7.3702
R456 VTAIL.n262 VTAIL.n261 7.3702
R457 VTAIL.n222 VTAIL.n221 7.3702
R458 VTAIL.n218 VTAIL.n217 7.3702
R459 VTAIL.n176 VTAIL.n175 7.3702
R460 VTAIL.n172 VTAIL.n171 7.3702
R461 VTAIL.n352 VTAIL.n318 6.59444
R462 VTAIL.n355 VTAIL.n318 6.59444
R463 VTAIL.n38 VTAIL.n4 6.59444
R464 VTAIL.n41 VTAIL.n4 6.59444
R465 VTAIL.n82 VTAIL.n48 6.59444
R466 VTAIL.n85 VTAIL.n48 6.59444
R467 VTAIL.n128 VTAIL.n94 6.59444
R468 VTAIL.n131 VTAIL.n94 6.59444
R469 VTAIL.n311 VTAIL.n274 6.59444
R470 VTAIL.n308 VTAIL.n274 6.59444
R471 VTAIL.n265 VTAIL.n228 6.59444
R472 VTAIL.n262 VTAIL.n228 6.59444
R473 VTAIL.n221 VTAIL.n184 6.59444
R474 VTAIL.n218 VTAIL.n184 6.59444
R475 VTAIL.n175 VTAIL.n138 6.59444
R476 VTAIL.n172 VTAIL.n138 6.59444
R477 VTAIL.n351 VTAIL.n320 5.81868
R478 VTAIL.n356 VTAIL.n316 5.81868
R479 VTAIL.n37 VTAIL.n6 5.81868
R480 VTAIL.n42 VTAIL.n2 5.81868
R481 VTAIL.n81 VTAIL.n50 5.81868
R482 VTAIL.n86 VTAIL.n46 5.81868
R483 VTAIL.n127 VTAIL.n96 5.81868
R484 VTAIL.n132 VTAIL.n92 5.81868
R485 VTAIL.n312 VTAIL.n272 5.81868
R486 VTAIL.n307 VTAIL.n276 5.81868
R487 VTAIL.n266 VTAIL.n226 5.81868
R488 VTAIL.n261 VTAIL.n230 5.81868
R489 VTAIL.n222 VTAIL.n182 5.81868
R490 VTAIL.n217 VTAIL.n186 5.81868
R491 VTAIL.n176 VTAIL.n136 5.81868
R492 VTAIL.n171 VTAIL.n140 5.81868
R493 VTAIL.n348 VTAIL.n347 5.04292
R494 VTAIL.n34 VTAIL.n33 5.04292
R495 VTAIL.n78 VTAIL.n77 5.04292
R496 VTAIL.n124 VTAIL.n123 5.04292
R497 VTAIL.n304 VTAIL.n303 5.04292
R498 VTAIL.n258 VTAIL.n257 5.04292
R499 VTAIL.n214 VTAIL.n213 5.04292
R500 VTAIL.n168 VTAIL.n167 5.04292
R501 VTAIL.n344 VTAIL.n322 4.26717
R502 VTAIL.n30 VTAIL.n8 4.26717
R503 VTAIL.n74 VTAIL.n52 4.26717
R504 VTAIL.n120 VTAIL.n98 4.26717
R505 VTAIL.n300 VTAIL.n278 4.26717
R506 VTAIL.n254 VTAIL.n232 4.26717
R507 VTAIL.n210 VTAIL.n188 4.26717
R508 VTAIL.n164 VTAIL.n142 4.26717
R509 VTAIL.n0 VTAIL.t1 3.99374
R510 VTAIL.n0 VTAIL.t0 3.99374
R511 VTAIL.n90 VTAIL.t8 3.99374
R512 VTAIL.n90 VTAIL.t15 3.99374
R513 VTAIL.n270 VTAIL.t10 3.99374
R514 VTAIL.n270 VTAIL.t11 3.99374
R515 VTAIL.n180 VTAIL.t6 3.99374
R516 VTAIL.n180 VTAIL.t4 3.99374
R517 VTAIL.n333 VTAIL.n329 3.70995
R518 VTAIL.n19 VTAIL.n15 3.70995
R519 VTAIL.n63 VTAIL.n59 3.70995
R520 VTAIL.n109 VTAIL.n105 3.70995
R521 VTAIL.n243 VTAIL.n239 3.70995
R522 VTAIL.n199 VTAIL.n195 3.70995
R523 VTAIL.n153 VTAIL.n149 3.70995
R524 VTAIL.n289 VTAIL.n285 3.70995
R525 VTAIL.n343 VTAIL.n324 3.49141
R526 VTAIL.n29 VTAIL.n10 3.49141
R527 VTAIL.n73 VTAIL.n54 3.49141
R528 VTAIL.n119 VTAIL.n100 3.49141
R529 VTAIL.n299 VTAIL.n280 3.49141
R530 VTAIL.n253 VTAIL.n234 3.49141
R531 VTAIL.n209 VTAIL.n190 3.49141
R532 VTAIL.n163 VTAIL.n144 3.49141
R533 VTAIL.n340 VTAIL.n339 2.71565
R534 VTAIL.n26 VTAIL.n25 2.71565
R535 VTAIL.n70 VTAIL.n69 2.71565
R536 VTAIL.n116 VTAIL.n115 2.71565
R537 VTAIL.n296 VTAIL.n295 2.71565
R538 VTAIL.n250 VTAIL.n249 2.71565
R539 VTAIL.n206 VTAIL.n205 2.71565
R540 VTAIL.n160 VTAIL.n159 2.71565
R541 VTAIL.n336 VTAIL.n326 1.93989
R542 VTAIL.n22 VTAIL.n12 1.93989
R543 VTAIL.n66 VTAIL.n56 1.93989
R544 VTAIL.n112 VTAIL.n102 1.93989
R545 VTAIL.n292 VTAIL.n282 1.93989
R546 VTAIL.n246 VTAIL.n236 1.93989
R547 VTAIL.n202 VTAIL.n192 1.93989
R548 VTAIL.n156 VTAIL.n146 1.93989
R549 VTAIL.n181 VTAIL.n179 1.62981
R550 VTAIL.n225 VTAIL.n181 1.62981
R551 VTAIL.n271 VTAIL.n269 1.62981
R552 VTAIL.n315 VTAIL.n271 1.62981
R553 VTAIL.n135 VTAIL.n91 1.62981
R554 VTAIL.n91 VTAIL.n89 1.62981
R555 VTAIL.n45 VTAIL.n1 1.62981
R556 VTAIL VTAIL.n359 1.57162
R557 VTAIL.n335 VTAIL.n328 1.16414
R558 VTAIL.n21 VTAIL.n14 1.16414
R559 VTAIL.n65 VTAIL.n58 1.16414
R560 VTAIL.n111 VTAIL.n104 1.16414
R561 VTAIL.n291 VTAIL.n284 1.16414
R562 VTAIL.n245 VTAIL.n238 1.16414
R563 VTAIL.n201 VTAIL.n194 1.16414
R564 VTAIL.n155 VTAIL.n148 1.16414
R565 VTAIL.n269 VTAIL.n225 0.470328
R566 VTAIL.n89 VTAIL.n45 0.470328
R567 VTAIL.n332 VTAIL.n331 0.388379
R568 VTAIL.n18 VTAIL.n17 0.388379
R569 VTAIL.n62 VTAIL.n61 0.388379
R570 VTAIL.n108 VTAIL.n107 0.388379
R571 VTAIL.n288 VTAIL.n287 0.388379
R572 VTAIL.n242 VTAIL.n241 0.388379
R573 VTAIL.n198 VTAIL.n197 0.388379
R574 VTAIL.n152 VTAIL.n151 0.388379
R575 VTAIL.n334 VTAIL.n333 0.155672
R576 VTAIL.n334 VTAIL.n325 0.155672
R577 VTAIL.n341 VTAIL.n325 0.155672
R578 VTAIL.n342 VTAIL.n341 0.155672
R579 VTAIL.n342 VTAIL.n321 0.155672
R580 VTAIL.n349 VTAIL.n321 0.155672
R581 VTAIL.n350 VTAIL.n349 0.155672
R582 VTAIL.n350 VTAIL.n317 0.155672
R583 VTAIL.n357 VTAIL.n317 0.155672
R584 VTAIL.n20 VTAIL.n19 0.155672
R585 VTAIL.n20 VTAIL.n11 0.155672
R586 VTAIL.n27 VTAIL.n11 0.155672
R587 VTAIL.n28 VTAIL.n27 0.155672
R588 VTAIL.n28 VTAIL.n7 0.155672
R589 VTAIL.n35 VTAIL.n7 0.155672
R590 VTAIL.n36 VTAIL.n35 0.155672
R591 VTAIL.n36 VTAIL.n3 0.155672
R592 VTAIL.n43 VTAIL.n3 0.155672
R593 VTAIL.n64 VTAIL.n63 0.155672
R594 VTAIL.n64 VTAIL.n55 0.155672
R595 VTAIL.n71 VTAIL.n55 0.155672
R596 VTAIL.n72 VTAIL.n71 0.155672
R597 VTAIL.n72 VTAIL.n51 0.155672
R598 VTAIL.n79 VTAIL.n51 0.155672
R599 VTAIL.n80 VTAIL.n79 0.155672
R600 VTAIL.n80 VTAIL.n47 0.155672
R601 VTAIL.n87 VTAIL.n47 0.155672
R602 VTAIL.n110 VTAIL.n109 0.155672
R603 VTAIL.n110 VTAIL.n101 0.155672
R604 VTAIL.n117 VTAIL.n101 0.155672
R605 VTAIL.n118 VTAIL.n117 0.155672
R606 VTAIL.n118 VTAIL.n97 0.155672
R607 VTAIL.n125 VTAIL.n97 0.155672
R608 VTAIL.n126 VTAIL.n125 0.155672
R609 VTAIL.n126 VTAIL.n93 0.155672
R610 VTAIL.n133 VTAIL.n93 0.155672
R611 VTAIL.n313 VTAIL.n273 0.155672
R612 VTAIL.n306 VTAIL.n273 0.155672
R613 VTAIL.n306 VTAIL.n305 0.155672
R614 VTAIL.n305 VTAIL.n277 0.155672
R615 VTAIL.n298 VTAIL.n277 0.155672
R616 VTAIL.n298 VTAIL.n297 0.155672
R617 VTAIL.n297 VTAIL.n281 0.155672
R618 VTAIL.n290 VTAIL.n281 0.155672
R619 VTAIL.n290 VTAIL.n289 0.155672
R620 VTAIL.n267 VTAIL.n227 0.155672
R621 VTAIL.n260 VTAIL.n227 0.155672
R622 VTAIL.n260 VTAIL.n259 0.155672
R623 VTAIL.n259 VTAIL.n231 0.155672
R624 VTAIL.n252 VTAIL.n231 0.155672
R625 VTAIL.n252 VTAIL.n251 0.155672
R626 VTAIL.n251 VTAIL.n235 0.155672
R627 VTAIL.n244 VTAIL.n235 0.155672
R628 VTAIL.n244 VTAIL.n243 0.155672
R629 VTAIL.n223 VTAIL.n183 0.155672
R630 VTAIL.n216 VTAIL.n183 0.155672
R631 VTAIL.n216 VTAIL.n215 0.155672
R632 VTAIL.n215 VTAIL.n187 0.155672
R633 VTAIL.n208 VTAIL.n187 0.155672
R634 VTAIL.n208 VTAIL.n207 0.155672
R635 VTAIL.n207 VTAIL.n191 0.155672
R636 VTAIL.n200 VTAIL.n191 0.155672
R637 VTAIL.n200 VTAIL.n199 0.155672
R638 VTAIL.n177 VTAIL.n137 0.155672
R639 VTAIL.n170 VTAIL.n137 0.155672
R640 VTAIL.n170 VTAIL.n169 0.155672
R641 VTAIL.n169 VTAIL.n141 0.155672
R642 VTAIL.n162 VTAIL.n141 0.155672
R643 VTAIL.n162 VTAIL.n161 0.155672
R644 VTAIL.n161 VTAIL.n145 0.155672
R645 VTAIL.n154 VTAIL.n145 0.155672
R646 VTAIL.n154 VTAIL.n153 0.155672
R647 VTAIL VTAIL.n1 0.0586897
R648 B.n422 B.n59 585
R649 B.n424 B.n423 585
R650 B.n425 B.n58 585
R651 B.n427 B.n426 585
R652 B.n428 B.n57 585
R653 B.n430 B.n429 585
R654 B.n431 B.n56 585
R655 B.n433 B.n432 585
R656 B.n434 B.n55 585
R657 B.n436 B.n435 585
R658 B.n437 B.n54 585
R659 B.n439 B.n438 585
R660 B.n440 B.n53 585
R661 B.n442 B.n441 585
R662 B.n443 B.n52 585
R663 B.n445 B.n444 585
R664 B.n446 B.n51 585
R665 B.n448 B.n447 585
R666 B.n449 B.n50 585
R667 B.n451 B.n450 585
R668 B.n452 B.n49 585
R669 B.n454 B.n453 585
R670 B.n455 B.n48 585
R671 B.n457 B.n456 585
R672 B.n458 B.n47 585
R673 B.n460 B.n459 585
R674 B.n461 B.n46 585
R675 B.n463 B.n462 585
R676 B.n464 B.n45 585
R677 B.n466 B.n465 585
R678 B.n468 B.n467 585
R679 B.n469 B.n41 585
R680 B.n471 B.n470 585
R681 B.n472 B.n40 585
R682 B.n474 B.n473 585
R683 B.n475 B.n39 585
R684 B.n477 B.n476 585
R685 B.n478 B.n38 585
R686 B.n480 B.n479 585
R687 B.n481 B.n35 585
R688 B.n484 B.n483 585
R689 B.n485 B.n34 585
R690 B.n487 B.n486 585
R691 B.n488 B.n33 585
R692 B.n490 B.n489 585
R693 B.n491 B.n32 585
R694 B.n493 B.n492 585
R695 B.n494 B.n31 585
R696 B.n496 B.n495 585
R697 B.n497 B.n30 585
R698 B.n499 B.n498 585
R699 B.n500 B.n29 585
R700 B.n502 B.n501 585
R701 B.n503 B.n28 585
R702 B.n505 B.n504 585
R703 B.n506 B.n27 585
R704 B.n508 B.n507 585
R705 B.n509 B.n26 585
R706 B.n511 B.n510 585
R707 B.n512 B.n25 585
R708 B.n514 B.n513 585
R709 B.n515 B.n24 585
R710 B.n517 B.n516 585
R711 B.n518 B.n23 585
R712 B.n520 B.n519 585
R713 B.n521 B.n22 585
R714 B.n523 B.n522 585
R715 B.n524 B.n21 585
R716 B.n526 B.n525 585
R717 B.n527 B.n20 585
R718 B.n421 B.n420 585
R719 B.n419 B.n60 585
R720 B.n418 B.n417 585
R721 B.n416 B.n61 585
R722 B.n415 B.n414 585
R723 B.n413 B.n62 585
R724 B.n412 B.n411 585
R725 B.n410 B.n63 585
R726 B.n409 B.n408 585
R727 B.n407 B.n64 585
R728 B.n406 B.n405 585
R729 B.n404 B.n65 585
R730 B.n403 B.n402 585
R731 B.n401 B.n66 585
R732 B.n400 B.n399 585
R733 B.n398 B.n67 585
R734 B.n397 B.n396 585
R735 B.n395 B.n68 585
R736 B.n394 B.n393 585
R737 B.n392 B.n69 585
R738 B.n391 B.n390 585
R739 B.n389 B.n70 585
R740 B.n388 B.n387 585
R741 B.n386 B.n71 585
R742 B.n385 B.n384 585
R743 B.n383 B.n72 585
R744 B.n382 B.n381 585
R745 B.n380 B.n73 585
R746 B.n379 B.n378 585
R747 B.n377 B.n74 585
R748 B.n376 B.n375 585
R749 B.n374 B.n75 585
R750 B.n373 B.n372 585
R751 B.n371 B.n76 585
R752 B.n370 B.n369 585
R753 B.n368 B.n77 585
R754 B.n367 B.n366 585
R755 B.n365 B.n78 585
R756 B.n364 B.n363 585
R757 B.n362 B.n79 585
R758 B.n361 B.n360 585
R759 B.n359 B.n80 585
R760 B.n358 B.n357 585
R761 B.n356 B.n81 585
R762 B.n355 B.n354 585
R763 B.n353 B.n82 585
R764 B.n352 B.n351 585
R765 B.n350 B.n83 585
R766 B.n349 B.n348 585
R767 B.n347 B.n84 585
R768 B.n346 B.n345 585
R769 B.n344 B.n85 585
R770 B.n343 B.n342 585
R771 B.n341 B.n86 585
R772 B.n340 B.n339 585
R773 B.n338 B.n87 585
R774 B.n337 B.n336 585
R775 B.n335 B.n88 585
R776 B.n334 B.n333 585
R777 B.n332 B.n89 585
R778 B.n331 B.n330 585
R779 B.n329 B.n90 585
R780 B.n328 B.n327 585
R781 B.n326 B.n91 585
R782 B.n325 B.n324 585
R783 B.n323 B.n92 585
R784 B.n322 B.n321 585
R785 B.n320 B.n93 585
R786 B.n319 B.n318 585
R787 B.n317 B.n94 585
R788 B.n316 B.n315 585
R789 B.n314 B.n95 585
R790 B.n313 B.n312 585
R791 B.n206 B.n135 585
R792 B.n208 B.n207 585
R793 B.n209 B.n134 585
R794 B.n211 B.n210 585
R795 B.n212 B.n133 585
R796 B.n214 B.n213 585
R797 B.n215 B.n132 585
R798 B.n217 B.n216 585
R799 B.n218 B.n131 585
R800 B.n220 B.n219 585
R801 B.n221 B.n130 585
R802 B.n223 B.n222 585
R803 B.n224 B.n129 585
R804 B.n226 B.n225 585
R805 B.n227 B.n128 585
R806 B.n229 B.n228 585
R807 B.n230 B.n127 585
R808 B.n232 B.n231 585
R809 B.n233 B.n126 585
R810 B.n235 B.n234 585
R811 B.n236 B.n125 585
R812 B.n238 B.n237 585
R813 B.n239 B.n124 585
R814 B.n241 B.n240 585
R815 B.n242 B.n123 585
R816 B.n244 B.n243 585
R817 B.n245 B.n122 585
R818 B.n247 B.n246 585
R819 B.n248 B.n121 585
R820 B.n250 B.n249 585
R821 B.n252 B.n251 585
R822 B.n253 B.n117 585
R823 B.n255 B.n254 585
R824 B.n256 B.n116 585
R825 B.n258 B.n257 585
R826 B.n259 B.n115 585
R827 B.n261 B.n260 585
R828 B.n262 B.n114 585
R829 B.n264 B.n263 585
R830 B.n265 B.n111 585
R831 B.n268 B.n267 585
R832 B.n269 B.n110 585
R833 B.n271 B.n270 585
R834 B.n272 B.n109 585
R835 B.n274 B.n273 585
R836 B.n275 B.n108 585
R837 B.n277 B.n276 585
R838 B.n278 B.n107 585
R839 B.n280 B.n279 585
R840 B.n281 B.n106 585
R841 B.n283 B.n282 585
R842 B.n284 B.n105 585
R843 B.n286 B.n285 585
R844 B.n287 B.n104 585
R845 B.n289 B.n288 585
R846 B.n290 B.n103 585
R847 B.n292 B.n291 585
R848 B.n293 B.n102 585
R849 B.n295 B.n294 585
R850 B.n296 B.n101 585
R851 B.n298 B.n297 585
R852 B.n299 B.n100 585
R853 B.n301 B.n300 585
R854 B.n302 B.n99 585
R855 B.n304 B.n303 585
R856 B.n305 B.n98 585
R857 B.n307 B.n306 585
R858 B.n308 B.n97 585
R859 B.n310 B.n309 585
R860 B.n311 B.n96 585
R861 B.n205 B.n204 585
R862 B.n203 B.n136 585
R863 B.n202 B.n201 585
R864 B.n200 B.n137 585
R865 B.n199 B.n198 585
R866 B.n197 B.n138 585
R867 B.n196 B.n195 585
R868 B.n194 B.n139 585
R869 B.n193 B.n192 585
R870 B.n191 B.n140 585
R871 B.n190 B.n189 585
R872 B.n188 B.n141 585
R873 B.n187 B.n186 585
R874 B.n185 B.n142 585
R875 B.n184 B.n183 585
R876 B.n182 B.n143 585
R877 B.n181 B.n180 585
R878 B.n179 B.n144 585
R879 B.n178 B.n177 585
R880 B.n176 B.n145 585
R881 B.n175 B.n174 585
R882 B.n173 B.n146 585
R883 B.n172 B.n171 585
R884 B.n170 B.n147 585
R885 B.n169 B.n168 585
R886 B.n167 B.n148 585
R887 B.n166 B.n165 585
R888 B.n164 B.n149 585
R889 B.n163 B.n162 585
R890 B.n161 B.n150 585
R891 B.n160 B.n159 585
R892 B.n158 B.n151 585
R893 B.n157 B.n156 585
R894 B.n155 B.n152 585
R895 B.n154 B.n153 585
R896 B.n2 B.n0 585
R897 B.n581 B.n1 585
R898 B.n580 B.n579 585
R899 B.n578 B.n3 585
R900 B.n577 B.n576 585
R901 B.n575 B.n4 585
R902 B.n574 B.n573 585
R903 B.n572 B.n5 585
R904 B.n571 B.n570 585
R905 B.n569 B.n6 585
R906 B.n568 B.n567 585
R907 B.n566 B.n7 585
R908 B.n565 B.n564 585
R909 B.n563 B.n8 585
R910 B.n562 B.n561 585
R911 B.n560 B.n9 585
R912 B.n559 B.n558 585
R913 B.n557 B.n10 585
R914 B.n556 B.n555 585
R915 B.n554 B.n11 585
R916 B.n553 B.n552 585
R917 B.n551 B.n12 585
R918 B.n550 B.n549 585
R919 B.n548 B.n13 585
R920 B.n547 B.n546 585
R921 B.n545 B.n14 585
R922 B.n544 B.n543 585
R923 B.n542 B.n15 585
R924 B.n541 B.n540 585
R925 B.n539 B.n16 585
R926 B.n538 B.n537 585
R927 B.n536 B.n17 585
R928 B.n535 B.n534 585
R929 B.n533 B.n18 585
R930 B.n532 B.n531 585
R931 B.n530 B.n19 585
R932 B.n529 B.n528 585
R933 B.n583 B.n582 585
R934 B.n204 B.n135 492.5
R935 B.n528 B.n527 492.5
R936 B.n312 B.n311 492.5
R937 B.n420 B.n59 492.5
R938 B.n112 B.t2 343.06
R939 B.n42 B.t10 343.06
R940 B.n118 B.t5 343.06
R941 B.n36 B.t7 343.06
R942 B.n112 B.t0 331.409
R943 B.n118 B.t3 331.409
R944 B.n36 B.t6 331.409
R945 B.n42 B.t9 331.409
R946 B.n113 B.t1 306.406
R947 B.n43 B.t11 306.406
R948 B.n119 B.t4 306.406
R949 B.n37 B.t8 306.406
R950 B.n204 B.n203 163.367
R951 B.n203 B.n202 163.367
R952 B.n202 B.n137 163.367
R953 B.n198 B.n137 163.367
R954 B.n198 B.n197 163.367
R955 B.n197 B.n196 163.367
R956 B.n196 B.n139 163.367
R957 B.n192 B.n139 163.367
R958 B.n192 B.n191 163.367
R959 B.n191 B.n190 163.367
R960 B.n190 B.n141 163.367
R961 B.n186 B.n141 163.367
R962 B.n186 B.n185 163.367
R963 B.n185 B.n184 163.367
R964 B.n184 B.n143 163.367
R965 B.n180 B.n143 163.367
R966 B.n180 B.n179 163.367
R967 B.n179 B.n178 163.367
R968 B.n178 B.n145 163.367
R969 B.n174 B.n145 163.367
R970 B.n174 B.n173 163.367
R971 B.n173 B.n172 163.367
R972 B.n172 B.n147 163.367
R973 B.n168 B.n147 163.367
R974 B.n168 B.n167 163.367
R975 B.n167 B.n166 163.367
R976 B.n166 B.n149 163.367
R977 B.n162 B.n149 163.367
R978 B.n162 B.n161 163.367
R979 B.n161 B.n160 163.367
R980 B.n160 B.n151 163.367
R981 B.n156 B.n151 163.367
R982 B.n156 B.n155 163.367
R983 B.n155 B.n154 163.367
R984 B.n154 B.n2 163.367
R985 B.n582 B.n2 163.367
R986 B.n582 B.n581 163.367
R987 B.n581 B.n580 163.367
R988 B.n580 B.n3 163.367
R989 B.n576 B.n3 163.367
R990 B.n576 B.n575 163.367
R991 B.n575 B.n574 163.367
R992 B.n574 B.n5 163.367
R993 B.n570 B.n5 163.367
R994 B.n570 B.n569 163.367
R995 B.n569 B.n568 163.367
R996 B.n568 B.n7 163.367
R997 B.n564 B.n7 163.367
R998 B.n564 B.n563 163.367
R999 B.n563 B.n562 163.367
R1000 B.n562 B.n9 163.367
R1001 B.n558 B.n9 163.367
R1002 B.n558 B.n557 163.367
R1003 B.n557 B.n556 163.367
R1004 B.n556 B.n11 163.367
R1005 B.n552 B.n11 163.367
R1006 B.n552 B.n551 163.367
R1007 B.n551 B.n550 163.367
R1008 B.n550 B.n13 163.367
R1009 B.n546 B.n13 163.367
R1010 B.n546 B.n545 163.367
R1011 B.n545 B.n544 163.367
R1012 B.n544 B.n15 163.367
R1013 B.n540 B.n15 163.367
R1014 B.n540 B.n539 163.367
R1015 B.n539 B.n538 163.367
R1016 B.n538 B.n17 163.367
R1017 B.n534 B.n17 163.367
R1018 B.n534 B.n533 163.367
R1019 B.n533 B.n532 163.367
R1020 B.n532 B.n19 163.367
R1021 B.n528 B.n19 163.367
R1022 B.n208 B.n135 163.367
R1023 B.n209 B.n208 163.367
R1024 B.n210 B.n209 163.367
R1025 B.n210 B.n133 163.367
R1026 B.n214 B.n133 163.367
R1027 B.n215 B.n214 163.367
R1028 B.n216 B.n215 163.367
R1029 B.n216 B.n131 163.367
R1030 B.n220 B.n131 163.367
R1031 B.n221 B.n220 163.367
R1032 B.n222 B.n221 163.367
R1033 B.n222 B.n129 163.367
R1034 B.n226 B.n129 163.367
R1035 B.n227 B.n226 163.367
R1036 B.n228 B.n227 163.367
R1037 B.n228 B.n127 163.367
R1038 B.n232 B.n127 163.367
R1039 B.n233 B.n232 163.367
R1040 B.n234 B.n233 163.367
R1041 B.n234 B.n125 163.367
R1042 B.n238 B.n125 163.367
R1043 B.n239 B.n238 163.367
R1044 B.n240 B.n239 163.367
R1045 B.n240 B.n123 163.367
R1046 B.n244 B.n123 163.367
R1047 B.n245 B.n244 163.367
R1048 B.n246 B.n245 163.367
R1049 B.n246 B.n121 163.367
R1050 B.n250 B.n121 163.367
R1051 B.n251 B.n250 163.367
R1052 B.n251 B.n117 163.367
R1053 B.n255 B.n117 163.367
R1054 B.n256 B.n255 163.367
R1055 B.n257 B.n256 163.367
R1056 B.n257 B.n115 163.367
R1057 B.n261 B.n115 163.367
R1058 B.n262 B.n261 163.367
R1059 B.n263 B.n262 163.367
R1060 B.n263 B.n111 163.367
R1061 B.n268 B.n111 163.367
R1062 B.n269 B.n268 163.367
R1063 B.n270 B.n269 163.367
R1064 B.n270 B.n109 163.367
R1065 B.n274 B.n109 163.367
R1066 B.n275 B.n274 163.367
R1067 B.n276 B.n275 163.367
R1068 B.n276 B.n107 163.367
R1069 B.n280 B.n107 163.367
R1070 B.n281 B.n280 163.367
R1071 B.n282 B.n281 163.367
R1072 B.n282 B.n105 163.367
R1073 B.n286 B.n105 163.367
R1074 B.n287 B.n286 163.367
R1075 B.n288 B.n287 163.367
R1076 B.n288 B.n103 163.367
R1077 B.n292 B.n103 163.367
R1078 B.n293 B.n292 163.367
R1079 B.n294 B.n293 163.367
R1080 B.n294 B.n101 163.367
R1081 B.n298 B.n101 163.367
R1082 B.n299 B.n298 163.367
R1083 B.n300 B.n299 163.367
R1084 B.n300 B.n99 163.367
R1085 B.n304 B.n99 163.367
R1086 B.n305 B.n304 163.367
R1087 B.n306 B.n305 163.367
R1088 B.n306 B.n97 163.367
R1089 B.n310 B.n97 163.367
R1090 B.n311 B.n310 163.367
R1091 B.n312 B.n95 163.367
R1092 B.n316 B.n95 163.367
R1093 B.n317 B.n316 163.367
R1094 B.n318 B.n317 163.367
R1095 B.n318 B.n93 163.367
R1096 B.n322 B.n93 163.367
R1097 B.n323 B.n322 163.367
R1098 B.n324 B.n323 163.367
R1099 B.n324 B.n91 163.367
R1100 B.n328 B.n91 163.367
R1101 B.n329 B.n328 163.367
R1102 B.n330 B.n329 163.367
R1103 B.n330 B.n89 163.367
R1104 B.n334 B.n89 163.367
R1105 B.n335 B.n334 163.367
R1106 B.n336 B.n335 163.367
R1107 B.n336 B.n87 163.367
R1108 B.n340 B.n87 163.367
R1109 B.n341 B.n340 163.367
R1110 B.n342 B.n341 163.367
R1111 B.n342 B.n85 163.367
R1112 B.n346 B.n85 163.367
R1113 B.n347 B.n346 163.367
R1114 B.n348 B.n347 163.367
R1115 B.n348 B.n83 163.367
R1116 B.n352 B.n83 163.367
R1117 B.n353 B.n352 163.367
R1118 B.n354 B.n353 163.367
R1119 B.n354 B.n81 163.367
R1120 B.n358 B.n81 163.367
R1121 B.n359 B.n358 163.367
R1122 B.n360 B.n359 163.367
R1123 B.n360 B.n79 163.367
R1124 B.n364 B.n79 163.367
R1125 B.n365 B.n364 163.367
R1126 B.n366 B.n365 163.367
R1127 B.n366 B.n77 163.367
R1128 B.n370 B.n77 163.367
R1129 B.n371 B.n370 163.367
R1130 B.n372 B.n371 163.367
R1131 B.n372 B.n75 163.367
R1132 B.n376 B.n75 163.367
R1133 B.n377 B.n376 163.367
R1134 B.n378 B.n377 163.367
R1135 B.n378 B.n73 163.367
R1136 B.n382 B.n73 163.367
R1137 B.n383 B.n382 163.367
R1138 B.n384 B.n383 163.367
R1139 B.n384 B.n71 163.367
R1140 B.n388 B.n71 163.367
R1141 B.n389 B.n388 163.367
R1142 B.n390 B.n389 163.367
R1143 B.n390 B.n69 163.367
R1144 B.n394 B.n69 163.367
R1145 B.n395 B.n394 163.367
R1146 B.n396 B.n395 163.367
R1147 B.n396 B.n67 163.367
R1148 B.n400 B.n67 163.367
R1149 B.n401 B.n400 163.367
R1150 B.n402 B.n401 163.367
R1151 B.n402 B.n65 163.367
R1152 B.n406 B.n65 163.367
R1153 B.n407 B.n406 163.367
R1154 B.n408 B.n407 163.367
R1155 B.n408 B.n63 163.367
R1156 B.n412 B.n63 163.367
R1157 B.n413 B.n412 163.367
R1158 B.n414 B.n413 163.367
R1159 B.n414 B.n61 163.367
R1160 B.n418 B.n61 163.367
R1161 B.n419 B.n418 163.367
R1162 B.n420 B.n419 163.367
R1163 B.n527 B.n526 163.367
R1164 B.n526 B.n21 163.367
R1165 B.n522 B.n21 163.367
R1166 B.n522 B.n521 163.367
R1167 B.n521 B.n520 163.367
R1168 B.n520 B.n23 163.367
R1169 B.n516 B.n23 163.367
R1170 B.n516 B.n515 163.367
R1171 B.n515 B.n514 163.367
R1172 B.n514 B.n25 163.367
R1173 B.n510 B.n25 163.367
R1174 B.n510 B.n509 163.367
R1175 B.n509 B.n508 163.367
R1176 B.n508 B.n27 163.367
R1177 B.n504 B.n27 163.367
R1178 B.n504 B.n503 163.367
R1179 B.n503 B.n502 163.367
R1180 B.n502 B.n29 163.367
R1181 B.n498 B.n29 163.367
R1182 B.n498 B.n497 163.367
R1183 B.n497 B.n496 163.367
R1184 B.n496 B.n31 163.367
R1185 B.n492 B.n31 163.367
R1186 B.n492 B.n491 163.367
R1187 B.n491 B.n490 163.367
R1188 B.n490 B.n33 163.367
R1189 B.n486 B.n33 163.367
R1190 B.n486 B.n485 163.367
R1191 B.n485 B.n484 163.367
R1192 B.n484 B.n35 163.367
R1193 B.n479 B.n35 163.367
R1194 B.n479 B.n478 163.367
R1195 B.n478 B.n477 163.367
R1196 B.n477 B.n39 163.367
R1197 B.n473 B.n39 163.367
R1198 B.n473 B.n472 163.367
R1199 B.n472 B.n471 163.367
R1200 B.n471 B.n41 163.367
R1201 B.n467 B.n41 163.367
R1202 B.n467 B.n466 163.367
R1203 B.n466 B.n45 163.367
R1204 B.n462 B.n45 163.367
R1205 B.n462 B.n461 163.367
R1206 B.n461 B.n460 163.367
R1207 B.n460 B.n47 163.367
R1208 B.n456 B.n47 163.367
R1209 B.n456 B.n455 163.367
R1210 B.n455 B.n454 163.367
R1211 B.n454 B.n49 163.367
R1212 B.n450 B.n49 163.367
R1213 B.n450 B.n449 163.367
R1214 B.n449 B.n448 163.367
R1215 B.n448 B.n51 163.367
R1216 B.n444 B.n51 163.367
R1217 B.n444 B.n443 163.367
R1218 B.n443 B.n442 163.367
R1219 B.n442 B.n53 163.367
R1220 B.n438 B.n53 163.367
R1221 B.n438 B.n437 163.367
R1222 B.n437 B.n436 163.367
R1223 B.n436 B.n55 163.367
R1224 B.n432 B.n55 163.367
R1225 B.n432 B.n431 163.367
R1226 B.n431 B.n430 163.367
R1227 B.n430 B.n57 163.367
R1228 B.n426 B.n57 163.367
R1229 B.n426 B.n425 163.367
R1230 B.n425 B.n424 163.367
R1231 B.n424 B.n59 163.367
R1232 B.n266 B.n113 59.5399
R1233 B.n120 B.n119 59.5399
R1234 B.n482 B.n37 59.5399
R1235 B.n44 B.n43 59.5399
R1236 B.n113 B.n112 36.655
R1237 B.n119 B.n118 36.655
R1238 B.n37 B.n36 36.655
R1239 B.n43 B.n42 36.655
R1240 B.n529 B.n20 32.0005
R1241 B.n422 B.n421 32.0005
R1242 B.n313 B.n96 32.0005
R1243 B.n206 B.n205 32.0005
R1244 B B.n583 18.0485
R1245 B.n525 B.n20 10.6151
R1246 B.n525 B.n524 10.6151
R1247 B.n524 B.n523 10.6151
R1248 B.n523 B.n22 10.6151
R1249 B.n519 B.n22 10.6151
R1250 B.n519 B.n518 10.6151
R1251 B.n518 B.n517 10.6151
R1252 B.n517 B.n24 10.6151
R1253 B.n513 B.n24 10.6151
R1254 B.n513 B.n512 10.6151
R1255 B.n512 B.n511 10.6151
R1256 B.n511 B.n26 10.6151
R1257 B.n507 B.n26 10.6151
R1258 B.n507 B.n506 10.6151
R1259 B.n506 B.n505 10.6151
R1260 B.n505 B.n28 10.6151
R1261 B.n501 B.n28 10.6151
R1262 B.n501 B.n500 10.6151
R1263 B.n500 B.n499 10.6151
R1264 B.n499 B.n30 10.6151
R1265 B.n495 B.n30 10.6151
R1266 B.n495 B.n494 10.6151
R1267 B.n494 B.n493 10.6151
R1268 B.n493 B.n32 10.6151
R1269 B.n489 B.n32 10.6151
R1270 B.n489 B.n488 10.6151
R1271 B.n488 B.n487 10.6151
R1272 B.n487 B.n34 10.6151
R1273 B.n483 B.n34 10.6151
R1274 B.n481 B.n480 10.6151
R1275 B.n480 B.n38 10.6151
R1276 B.n476 B.n38 10.6151
R1277 B.n476 B.n475 10.6151
R1278 B.n475 B.n474 10.6151
R1279 B.n474 B.n40 10.6151
R1280 B.n470 B.n40 10.6151
R1281 B.n470 B.n469 10.6151
R1282 B.n469 B.n468 10.6151
R1283 B.n465 B.n464 10.6151
R1284 B.n464 B.n463 10.6151
R1285 B.n463 B.n46 10.6151
R1286 B.n459 B.n46 10.6151
R1287 B.n459 B.n458 10.6151
R1288 B.n458 B.n457 10.6151
R1289 B.n457 B.n48 10.6151
R1290 B.n453 B.n48 10.6151
R1291 B.n453 B.n452 10.6151
R1292 B.n452 B.n451 10.6151
R1293 B.n451 B.n50 10.6151
R1294 B.n447 B.n50 10.6151
R1295 B.n447 B.n446 10.6151
R1296 B.n446 B.n445 10.6151
R1297 B.n445 B.n52 10.6151
R1298 B.n441 B.n52 10.6151
R1299 B.n441 B.n440 10.6151
R1300 B.n440 B.n439 10.6151
R1301 B.n439 B.n54 10.6151
R1302 B.n435 B.n54 10.6151
R1303 B.n435 B.n434 10.6151
R1304 B.n434 B.n433 10.6151
R1305 B.n433 B.n56 10.6151
R1306 B.n429 B.n56 10.6151
R1307 B.n429 B.n428 10.6151
R1308 B.n428 B.n427 10.6151
R1309 B.n427 B.n58 10.6151
R1310 B.n423 B.n58 10.6151
R1311 B.n423 B.n422 10.6151
R1312 B.n314 B.n313 10.6151
R1313 B.n315 B.n314 10.6151
R1314 B.n315 B.n94 10.6151
R1315 B.n319 B.n94 10.6151
R1316 B.n320 B.n319 10.6151
R1317 B.n321 B.n320 10.6151
R1318 B.n321 B.n92 10.6151
R1319 B.n325 B.n92 10.6151
R1320 B.n326 B.n325 10.6151
R1321 B.n327 B.n326 10.6151
R1322 B.n327 B.n90 10.6151
R1323 B.n331 B.n90 10.6151
R1324 B.n332 B.n331 10.6151
R1325 B.n333 B.n332 10.6151
R1326 B.n333 B.n88 10.6151
R1327 B.n337 B.n88 10.6151
R1328 B.n338 B.n337 10.6151
R1329 B.n339 B.n338 10.6151
R1330 B.n339 B.n86 10.6151
R1331 B.n343 B.n86 10.6151
R1332 B.n344 B.n343 10.6151
R1333 B.n345 B.n344 10.6151
R1334 B.n345 B.n84 10.6151
R1335 B.n349 B.n84 10.6151
R1336 B.n350 B.n349 10.6151
R1337 B.n351 B.n350 10.6151
R1338 B.n351 B.n82 10.6151
R1339 B.n355 B.n82 10.6151
R1340 B.n356 B.n355 10.6151
R1341 B.n357 B.n356 10.6151
R1342 B.n357 B.n80 10.6151
R1343 B.n361 B.n80 10.6151
R1344 B.n362 B.n361 10.6151
R1345 B.n363 B.n362 10.6151
R1346 B.n363 B.n78 10.6151
R1347 B.n367 B.n78 10.6151
R1348 B.n368 B.n367 10.6151
R1349 B.n369 B.n368 10.6151
R1350 B.n369 B.n76 10.6151
R1351 B.n373 B.n76 10.6151
R1352 B.n374 B.n373 10.6151
R1353 B.n375 B.n374 10.6151
R1354 B.n375 B.n74 10.6151
R1355 B.n379 B.n74 10.6151
R1356 B.n380 B.n379 10.6151
R1357 B.n381 B.n380 10.6151
R1358 B.n381 B.n72 10.6151
R1359 B.n385 B.n72 10.6151
R1360 B.n386 B.n385 10.6151
R1361 B.n387 B.n386 10.6151
R1362 B.n387 B.n70 10.6151
R1363 B.n391 B.n70 10.6151
R1364 B.n392 B.n391 10.6151
R1365 B.n393 B.n392 10.6151
R1366 B.n393 B.n68 10.6151
R1367 B.n397 B.n68 10.6151
R1368 B.n398 B.n397 10.6151
R1369 B.n399 B.n398 10.6151
R1370 B.n399 B.n66 10.6151
R1371 B.n403 B.n66 10.6151
R1372 B.n404 B.n403 10.6151
R1373 B.n405 B.n404 10.6151
R1374 B.n405 B.n64 10.6151
R1375 B.n409 B.n64 10.6151
R1376 B.n410 B.n409 10.6151
R1377 B.n411 B.n410 10.6151
R1378 B.n411 B.n62 10.6151
R1379 B.n415 B.n62 10.6151
R1380 B.n416 B.n415 10.6151
R1381 B.n417 B.n416 10.6151
R1382 B.n417 B.n60 10.6151
R1383 B.n421 B.n60 10.6151
R1384 B.n207 B.n206 10.6151
R1385 B.n207 B.n134 10.6151
R1386 B.n211 B.n134 10.6151
R1387 B.n212 B.n211 10.6151
R1388 B.n213 B.n212 10.6151
R1389 B.n213 B.n132 10.6151
R1390 B.n217 B.n132 10.6151
R1391 B.n218 B.n217 10.6151
R1392 B.n219 B.n218 10.6151
R1393 B.n219 B.n130 10.6151
R1394 B.n223 B.n130 10.6151
R1395 B.n224 B.n223 10.6151
R1396 B.n225 B.n224 10.6151
R1397 B.n225 B.n128 10.6151
R1398 B.n229 B.n128 10.6151
R1399 B.n230 B.n229 10.6151
R1400 B.n231 B.n230 10.6151
R1401 B.n231 B.n126 10.6151
R1402 B.n235 B.n126 10.6151
R1403 B.n236 B.n235 10.6151
R1404 B.n237 B.n236 10.6151
R1405 B.n237 B.n124 10.6151
R1406 B.n241 B.n124 10.6151
R1407 B.n242 B.n241 10.6151
R1408 B.n243 B.n242 10.6151
R1409 B.n243 B.n122 10.6151
R1410 B.n247 B.n122 10.6151
R1411 B.n248 B.n247 10.6151
R1412 B.n249 B.n248 10.6151
R1413 B.n253 B.n252 10.6151
R1414 B.n254 B.n253 10.6151
R1415 B.n254 B.n116 10.6151
R1416 B.n258 B.n116 10.6151
R1417 B.n259 B.n258 10.6151
R1418 B.n260 B.n259 10.6151
R1419 B.n260 B.n114 10.6151
R1420 B.n264 B.n114 10.6151
R1421 B.n265 B.n264 10.6151
R1422 B.n267 B.n110 10.6151
R1423 B.n271 B.n110 10.6151
R1424 B.n272 B.n271 10.6151
R1425 B.n273 B.n272 10.6151
R1426 B.n273 B.n108 10.6151
R1427 B.n277 B.n108 10.6151
R1428 B.n278 B.n277 10.6151
R1429 B.n279 B.n278 10.6151
R1430 B.n279 B.n106 10.6151
R1431 B.n283 B.n106 10.6151
R1432 B.n284 B.n283 10.6151
R1433 B.n285 B.n284 10.6151
R1434 B.n285 B.n104 10.6151
R1435 B.n289 B.n104 10.6151
R1436 B.n290 B.n289 10.6151
R1437 B.n291 B.n290 10.6151
R1438 B.n291 B.n102 10.6151
R1439 B.n295 B.n102 10.6151
R1440 B.n296 B.n295 10.6151
R1441 B.n297 B.n296 10.6151
R1442 B.n297 B.n100 10.6151
R1443 B.n301 B.n100 10.6151
R1444 B.n302 B.n301 10.6151
R1445 B.n303 B.n302 10.6151
R1446 B.n303 B.n98 10.6151
R1447 B.n307 B.n98 10.6151
R1448 B.n308 B.n307 10.6151
R1449 B.n309 B.n308 10.6151
R1450 B.n309 B.n96 10.6151
R1451 B.n205 B.n136 10.6151
R1452 B.n201 B.n136 10.6151
R1453 B.n201 B.n200 10.6151
R1454 B.n200 B.n199 10.6151
R1455 B.n199 B.n138 10.6151
R1456 B.n195 B.n138 10.6151
R1457 B.n195 B.n194 10.6151
R1458 B.n194 B.n193 10.6151
R1459 B.n193 B.n140 10.6151
R1460 B.n189 B.n140 10.6151
R1461 B.n189 B.n188 10.6151
R1462 B.n188 B.n187 10.6151
R1463 B.n187 B.n142 10.6151
R1464 B.n183 B.n142 10.6151
R1465 B.n183 B.n182 10.6151
R1466 B.n182 B.n181 10.6151
R1467 B.n181 B.n144 10.6151
R1468 B.n177 B.n144 10.6151
R1469 B.n177 B.n176 10.6151
R1470 B.n176 B.n175 10.6151
R1471 B.n175 B.n146 10.6151
R1472 B.n171 B.n146 10.6151
R1473 B.n171 B.n170 10.6151
R1474 B.n170 B.n169 10.6151
R1475 B.n169 B.n148 10.6151
R1476 B.n165 B.n148 10.6151
R1477 B.n165 B.n164 10.6151
R1478 B.n164 B.n163 10.6151
R1479 B.n163 B.n150 10.6151
R1480 B.n159 B.n150 10.6151
R1481 B.n159 B.n158 10.6151
R1482 B.n158 B.n157 10.6151
R1483 B.n157 B.n152 10.6151
R1484 B.n153 B.n152 10.6151
R1485 B.n153 B.n0 10.6151
R1486 B.n579 B.n1 10.6151
R1487 B.n579 B.n578 10.6151
R1488 B.n578 B.n577 10.6151
R1489 B.n577 B.n4 10.6151
R1490 B.n573 B.n4 10.6151
R1491 B.n573 B.n572 10.6151
R1492 B.n572 B.n571 10.6151
R1493 B.n571 B.n6 10.6151
R1494 B.n567 B.n6 10.6151
R1495 B.n567 B.n566 10.6151
R1496 B.n566 B.n565 10.6151
R1497 B.n565 B.n8 10.6151
R1498 B.n561 B.n8 10.6151
R1499 B.n561 B.n560 10.6151
R1500 B.n560 B.n559 10.6151
R1501 B.n559 B.n10 10.6151
R1502 B.n555 B.n10 10.6151
R1503 B.n555 B.n554 10.6151
R1504 B.n554 B.n553 10.6151
R1505 B.n553 B.n12 10.6151
R1506 B.n549 B.n12 10.6151
R1507 B.n549 B.n548 10.6151
R1508 B.n548 B.n547 10.6151
R1509 B.n547 B.n14 10.6151
R1510 B.n543 B.n14 10.6151
R1511 B.n543 B.n542 10.6151
R1512 B.n542 B.n541 10.6151
R1513 B.n541 B.n16 10.6151
R1514 B.n537 B.n16 10.6151
R1515 B.n537 B.n536 10.6151
R1516 B.n536 B.n535 10.6151
R1517 B.n535 B.n18 10.6151
R1518 B.n531 B.n18 10.6151
R1519 B.n531 B.n530 10.6151
R1520 B.n530 B.n529 10.6151
R1521 B.n483 B.n482 9.36635
R1522 B.n465 B.n44 9.36635
R1523 B.n249 B.n120 9.36635
R1524 B.n267 B.n266 9.36635
R1525 B.n583 B.n0 2.81026
R1526 B.n583 B.n1 2.81026
R1527 B.n482 B.n481 1.24928
R1528 B.n468 B.n44 1.24928
R1529 B.n252 B.n120 1.24928
R1530 B.n266 B.n265 1.24928
R1531 VN.n20 VN.n19 181.506
R1532 VN.n41 VN.n40 181.506
R1533 VN.n39 VN.n21 161.3
R1534 VN.n38 VN.n37 161.3
R1535 VN.n36 VN.n22 161.3
R1536 VN.n35 VN.n34 161.3
R1537 VN.n32 VN.n23 161.3
R1538 VN.n31 VN.n30 161.3
R1539 VN.n29 VN.n24 161.3
R1540 VN.n28 VN.n27 161.3
R1541 VN.n18 VN.n0 161.3
R1542 VN.n17 VN.n16 161.3
R1543 VN.n15 VN.n1 161.3
R1544 VN.n14 VN.n13 161.3
R1545 VN.n11 VN.n2 161.3
R1546 VN.n10 VN.n9 161.3
R1547 VN.n8 VN.n3 161.3
R1548 VN.n7 VN.n6 161.3
R1549 VN.n4 VN.t6 156.085
R1550 VN.n25 VN.t5 156.085
R1551 VN.n5 VN.t3 125.754
R1552 VN.n12 VN.t1 125.754
R1553 VN.n19 VN.t7 125.754
R1554 VN.n26 VN.t4 125.754
R1555 VN.n33 VN.t0 125.754
R1556 VN.n40 VN.t2 125.754
R1557 VN.n5 VN.n4 56.704
R1558 VN.n26 VN.n25 56.704
R1559 VN.n10 VN.n3 56.4773
R1560 VN.n31 VN.n24 56.4773
R1561 VN.n17 VN.n1 54.0429
R1562 VN.n38 VN.n22 54.0429
R1563 VN VN.n41 43.3357
R1564 VN.n13 VN.n1 26.7783
R1565 VN.n34 VN.n22 26.7783
R1566 VN.n6 VN.n3 24.3439
R1567 VN.n11 VN.n10 24.3439
R1568 VN.n18 VN.n17 24.3439
R1569 VN.n27 VN.n24 24.3439
R1570 VN.n32 VN.n31 24.3439
R1571 VN.n39 VN.n38 24.3439
R1572 VN.n28 VN.n25 18.4239
R1573 VN.n7 VN.n4 18.4239
R1574 VN.n13 VN.n12 14.85
R1575 VN.n34 VN.n33 14.85
R1576 VN.n6 VN.n5 9.49444
R1577 VN.n12 VN.n11 9.49444
R1578 VN.n27 VN.n26 9.49444
R1579 VN.n33 VN.n32 9.49444
R1580 VN.n19 VN.n18 4.13888
R1581 VN.n40 VN.n39 4.13888
R1582 VN.n41 VN.n21 0.189894
R1583 VN.n37 VN.n21 0.189894
R1584 VN.n37 VN.n36 0.189894
R1585 VN.n36 VN.n35 0.189894
R1586 VN.n35 VN.n23 0.189894
R1587 VN.n30 VN.n23 0.189894
R1588 VN.n30 VN.n29 0.189894
R1589 VN.n29 VN.n28 0.189894
R1590 VN.n8 VN.n7 0.189894
R1591 VN.n9 VN.n8 0.189894
R1592 VN.n9 VN.n2 0.189894
R1593 VN.n14 VN.n2 0.189894
R1594 VN.n15 VN.n14 0.189894
R1595 VN.n16 VN.n15 0.189894
R1596 VN.n16 VN.n0 0.189894
R1597 VN.n20 VN.n0 0.189894
R1598 VN VN.n20 0.0516364
R1599 VDD2.n2 VDD2.n1 83.1582
R1600 VDD2.n2 VDD2.n0 83.1582
R1601 VDD2 VDD2.n5 83.1555
R1602 VDD2.n4 VDD2.n3 82.3991
R1603 VDD2.n4 VDD2.n2 38.0644
R1604 VDD2.n5 VDD2.t3 3.99374
R1605 VDD2.n5 VDD2.t2 3.99374
R1606 VDD2.n3 VDD2.t5 3.99374
R1607 VDD2.n3 VDD2.t7 3.99374
R1608 VDD2.n1 VDD2.t6 3.99374
R1609 VDD2.n1 VDD2.t0 3.99374
R1610 VDD2.n0 VDD2.t1 3.99374
R1611 VDD2.n0 VDD2.t4 3.99374
R1612 VDD2 VDD2.n4 0.873345
C0 B VDD1 1.22883f
C1 VTAIL VP 5.55379f
C2 w_n2860_n2596# VN 5.469f
C3 VDD2 VN 5.32519f
C4 B VP 1.54663f
C5 VN VDD1 0.14948f
C6 w_n2860_n2596# VDD2 1.58036f
C7 w_n2860_n2596# VDD1 1.50925f
C8 VDD2 VDD1 1.25099f
C9 B VTAIL 3.27138f
C10 VN VP 5.68299f
C11 w_n2860_n2596# VP 5.83722f
C12 VDD2 VP 0.408636f
C13 VDD1 VP 5.58348f
C14 VN VTAIL 5.53968f
C15 w_n2860_n2596# VTAIL 3.25561f
C16 B VN 0.934904f
C17 VDD2 VTAIL 6.70391f
C18 w_n2860_n2596# B 7.44024f
C19 VTAIL VDD1 6.65647f
C20 B VDD2 1.29215f
C21 VDD2 VSUBS 1.393499f
C22 VDD1 VSUBS 1.862478f
C23 VTAIL VSUBS 0.951708f
C24 VN VSUBS 5.27987f
C25 VP VSUBS 2.364542f
C26 B VSUBS 3.516276f
C27 w_n2860_n2596# VSUBS 92.0806f
C28 VDD2.t1 VSUBS 0.159297f
C29 VDD2.t4 VSUBS 0.159297f
C30 VDD2.n0 VSUBS 1.1456f
C31 VDD2.t6 VSUBS 0.159297f
C32 VDD2.t0 VSUBS 0.159297f
C33 VDD2.n1 VSUBS 1.1456f
C34 VDD2.n2 VSUBS 2.883f
C35 VDD2.t5 VSUBS 0.159297f
C36 VDD2.t7 VSUBS 0.159297f
C37 VDD2.n3 VSUBS 1.13976f
C38 VDD2.n4 VSUBS 2.50254f
C39 VDD2.t3 VSUBS 0.159297f
C40 VDD2.t2 VSUBS 0.159297f
C41 VDD2.n5 VSUBS 1.14558f
C42 VN.n0 VSUBS 0.041399f
C43 VN.t7 VSUBS 1.41295f
C44 VN.n1 VSUBS 0.045349f
C45 VN.n2 VSUBS 0.041399f
C46 VN.t1 VSUBS 1.41295f
C47 VN.n3 VSUBS 0.060699f
C48 VN.t6 VSUBS 1.54776f
C49 VN.n4 VSUBS 0.631279f
C50 VN.t3 VSUBS 1.41295f
C51 VN.n5 VSUBS 0.605477f
C52 VN.n6 VSUBS 0.05419f
C53 VN.n7 VSUBS 0.259884f
C54 VN.n8 VSUBS 0.041399f
C55 VN.n9 VSUBS 0.041399f
C56 VN.n10 VSUBS 0.060699f
C57 VN.n11 VSUBS 0.05419f
C58 VN.n12 VSUBS 0.529379f
C59 VN.n13 VSUBS 0.065746f
C60 VN.n14 VSUBS 0.041399f
C61 VN.n15 VSUBS 0.041399f
C62 VN.n16 VSUBS 0.041399f
C63 VN.n17 VSUBS 0.072916f
C64 VN.n18 VSUBS 0.045767f
C65 VN.n19 VSUBS 0.608159f
C66 VN.n20 VSUBS 0.041951f
C67 VN.n21 VSUBS 0.041399f
C68 VN.t2 VSUBS 1.41295f
C69 VN.n22 VSUBS 0.045349f
C70 VN.n23 VSUBS 0.041399f
C71 VN.t0 VSUBS 1.41295f
C72 VN.n24 VSUBS 0.060699f
C73 VN.t5 VSUBS 1.54776f
C74 VN.n25 VSUBS 0.631279f
C75 VN.t4 VSUBS 1.41295f
C76 VN.n26 VSUBS 0.605477f
C77 VN.n27 VSUBS 0.05419f
C78 VN.n28 VSUBS 0.259884f
C79 VN.n29 VSUBS 0.041399f
C80 VN.n30 VSUBS 0.041399f
C81 VN.n31 VSUBS 0.060699f
C82 VN.n32 VSUBS 0.05419f
C83 VN.n33 VSUBS 0.529379f
C84 VN.n34 VSUBS 0.065746f
C85 VN.n35 VSUBS 0.041399f
C86 VN.n36 VSUBS 0.041399f
C87 VN.n37 VSUBS 0.041399f
C88 VN.n38 VSUBS 0.072916f
C89 VN.n39 VSUBS 0.045767f
C90 VN.n40 VSUBS 0.608159f
C91 VN.n41 VSUBS 1.81065f
C92 B.n0 VSUBS 0.00506f
C93 B.n1 VSUBS 0.00506f
C94 B.n2 VSUBS 0.008001f
C95 B.n3 VSUBS 0.008001f
C96 B.n4 VSUBS 0.008001f
C97 B.n5 VSUBS 0.008001f
C98 B.n6 VSUBS 0.008001f
C99 B.n7 VSUBS 0.008001f
C100 B.n8 VSUBS 0.008001f
C101 B.n9 VSUBS 0.008001f
C102 B.n10 VSUBS 0.008001f
C103 B.n11 VSUBS 0.008001f
C104 B.n12 VSUBS 0.008001f
C105 B.n13 VSUBS 0.008001f
C106 B.n14 VSUBS 0.008001f
C107 B.n15 VSUBS 0.008001f
C108 B.n16 VSUBS 0.008001f
C109 B.n17 VSUBS 0.008001f
C110 B.n18 VSUBS 0.008001f
C111 B.n19 VSUBS 0.008001f
C112 B.n20 VSUBS 0.018815f
C113 B.n21 VSUBS 0.008001f
C114 B.n22 VSUBS 0.008001f
C115 B.n23 VSUBS 0.008001f
C116 B.n24 VSUBS 0.008001f
C117 B.n25 VSUBS 0.008001f
C118 B.n26 VSUBS 0.008001f
C119 B.n27 VSUBS 0.008001f
C120 B.n28 VSUBS 0.008001f
C121 B.n29 VSUBS 0.008001f
C122 B.n30 VSUBS 0.008001f
C123 B.n31 VSUBS 0.008001f
C124 B.n32 VSUBS 0.008001f
C125 B.n33 VSUBS 0.008001f
C126 B.n34 VSUBS 0.008001f
C127 B.n35 VSUBS 0.008001f
C128 B.t8 VSUBS 0.1482f
C129 B.t7 VSUBS 0.170104f
C130 B.t6 VSUBS 0.653861f
C131 B.n36 VSUBS 0.28224f
C132 B.n37 VSUBS 0.216415f
C133 B.n38 VSUBS 0.008001f
C134 B.n39 VSUBS 0.008001f
C135 B.n40 VSUBS 0.008001f
C136 B.n41 VSUBS 0.008001f
C137 B.t11 VSUBS 0.148203f
C138 B.t10 VSUBS 0.170106f
C139 B.t9 VSUBS 0.653861f
C140 B.n42 VSUBS 0.282238f
C141 B.n43 VSUBS 0.216413f
C142 B.n44 VSUBS 0.018538f
C143 B.n45 VSUBS 0.008001f
C144 B.n46 VSUBS 0.008001f
C145 B.n47 VSUBS 0.008001f
C146 B.n48 VSUBS 0.008001f
C147 B.n49 VSUBS 0.008001f
C148 B.n50 VSUBS 0.008001f
C149 B.n51 VSUBS 0.008001f
C150 B.n52 VSUBS 0.008001f
C151 B.n53 VSUBS 0.008001f
C152 B.n54 VSUBS 0.008001f
C153 B.n55 VSUBS 0.008001f
C154 B.n56 VSUBS 0.008001f
C155 B.n57 VSUBS 0.008001f
C156 B.n58 VSUBS 0.008001f
C157 B.n59 VSUBS 0.018815f
C158 B.n60 VSUBS 0.008001f
C159 B.n61 VSUBS 0.008001f
C160 B.n62 VSUBS 0.008001f
C161 B.n63 VSUBS 0.008001f
C162 B.n64 VSUBS 0.008001f
C163 B.n65 VSUBS 0.008001f
C164 B.n66 VSUBS 0.008001f
C165 B.n67 VSUBS 0.008001f
C166 B.n68 VSUBS 0.008001f
C167 B.n69 VSUBS 0.008001f
C168 B.n70 VSUBS 0.008001f
C169 B.n71 VSUBS 0.008001f
C170 B.n72 VSUBS 0.008001f
C171 B.n73 VSUBS 0.008001f
C172 B.n74 VSUBS 0.008001f
C173 B.n75 VSUBS 0.008001f
C174 B.n76 VSUBS 0.008001f
C175 B.n77 VSUBS 0.008001f
C176 B.n78 VSUBS 0.008001f
C177 B.n79 VSUBS 0.008001f
C178 B.n80 VSUBS 0.008001f
C179 B.n81 VSUBS 0.008001f
C180 B.n82 VSUBS 0.008001f
C181 B.n83 VSUBS 0.008001f
C182 B.n84 VSUBS 0.008001f
C183 B.n85 VSUBS 0.008001f
C184 B.n86 VSUBS 0.008001f
C185 B.n87 VSUBS 0.008001f
C186 B.n88 VSUBS 0.008001f
C187 B.n89 VSUBS 0.008001f
C188 B.n90 VSUBS 0.008001f
C189 B.n91 VSUBS 0.008001f
C190 B.n92 VSUBS 0.008001f
C191 B.n93 VSUBS 0.008001f
C192 B.n94 VSUBS 0.008001f
C193 B.n95 VSUBS 0.008001f
C194 B.n96 VSUBS 0.018815f
C195 B.n97 VSUBS 0.008001f
C196 B.n98 VSUBS 0.008001f
C197 B.n99 VSUBS 0.008001f
C198 B.n100 VSUBS 0.008001f
C199 B.n101 VSUBS 0.008001f
C200 B.n102 VSUBS 0.008001f
C201 B.n103 VSUBS 0.008001f
C202 B.n104 VSUBS 0.008001f
C203 B.n105 VSUBS 0.008001f
C204 B.n106 VSUBS 0.008001f
C205 B.n107 VSUBS 0.008001f
C206 B.n108 VSUBS 0.008001f
C207 B.n109 VSUBS 0.008001f
C208 B.n110 VSUBS 0.008001f
C209 B.n111 VSUBS 0.008001f
C210 B.t1 VSUBS 0.148203f
C211 B.t2 VSUBS 0.170106f
C212 B.t0 VSUBS 0.653861f
C213 B.n112 VSUBS 0.282238f
C214 B.n113 VSUBS 0.216413f
C215 B.n114 VSUBS 0.008001f
C216 B.n115 VSUBS 0.008001f
C217 B.n116 VSUBS 0.008001f
C218 B.n117 VSUBS 0.008001f
C219 B.t4 VSUBS 0.1482f
C220 B.t5 VSUBS 0.170104f
C221 B.t3 VSUBS 0.653861f
C222 B.n118 VSUBS 0.28224f
C223 B.n119 VSUBS 0.216415f
C224 B.n120 VSUBS 0.018538f
C225 B.n121 VSUBS 0.008001f
C226 B.n122 VSUBS 0.008001f
C227 B.n123 VSUBS 0.008001f
C228 B.n124 VSUBS 0.008001f
C229 B.n125 VSUBS 0.008001f
C230 B.n126 VSUBS 0.008001f
C231 B.n127 VSUBS 0.008001f
C232 B.n128 VSUBS 0.008001f
C233 B.n129 VSUBS 0.008001f
C234 B.n130 VSUBS 0.008001f
C235 B.n131 VSUBS 0.008001f
C236 B.n132 VSUBS 0.008001f
C237 B.n133 VSUBS 0.008001f
C238 B.n134 VSUBS 0.008001f
C239 B.n135 VSUBS 0.018815f
C240 B.n136 VSUBS 0.008001f
C241 B.n137 VSUBS 0.008001f
C242 B.n138 VSUBS 0.008001f
C243 B.n139 VSUBS 0.008001f
C244 B.n140 VSUBS 0.008001f
C245 B.n141 VSUBS 0.008001f
C246 B.n142 VSUBS 0.008001f
C247 B.n143 VSUBS 0.008001f
C248 B.n144 VSUBS 0.008001f
C249 B.n145 VSUBS 0.008001f
C250 B.n146 VSUBS 0.008001f
C251 B.n147 VSUBS 0.008001f
C252 B.n148 VSUBS 0.008001f
C253 B.n149 VSUBS 0.008001f
C254 B.n150 VSUBS 0.008001f
C255 B.n151 VSUBS 0.008001f
C256 B.n152 VSUBS 0.008001f
C257 B.n153 VSUBS 0.008001f
C258 B.n154 VSUBS 0.008001f
C259 B.n155 VSUBS 0.008001f
C260 B.n156 VSUBS 0.008001f
C261 B.n157 VSUBS 0.008001f
C262 B.n158 VSUBS 0.008001f
C263 B.n159 VSUBS 0.008001f
C264 B.n160 VSUBS 0.008001f
C265 B.n161 VSUBS 0.008001f
C266 B.n162 VSUBS 0.008001f
C267 B.n163 VSUBS 0.008001f
C268 B.n164 VSUBS 0.008001f
C269 B.n165 VSUBS 0.008001f
C270 B.n166 VSUBS 0.008001f
C271 B.n167 VSUBS 0.008001f
C272 B.n168 VSUBS 0.008001f
C273 B.n169 VSUBS 0.008001f
C274 B.n170 VSUBS 0.008001f
C275 B.n171 VSUBS 0.008001f
C276 B.n172 VSUBS 0.008001f
C277 B.n173 VSUBS 0.008001f
C278 B.n174 VSUBS 0.008001f
C279 B.n175 VSUBS 0.008001f
C280 B.n176 VSUBS 0.008001f
C281 B.n177 VSUBS 0.008001f
C282 B.n178 VSUBS 0.008001f
C283 B.n179 VSUBS 0.008001f
C284 B.n180 VSUBS 0.008001f
C285 B.n181 VSUBS 0.008001f
C286 B.n182 VSUBS 0.008001f
C287 B.n183 VSUBS 0.008001f
C288 B.n184 VSUBS 0.008001f
C289 B.n185 VSUBS 0.008001f
C290 B.n186 VSUBS 0.008001f
C291 B.n187 VSUBS 0.008001f
C292 B.n188 VSUBS 0.008001f
C293 B.n189 VSUBS 0.008001f
C294 B.n190 VSUBS 0.008001f
C295 B.n191 VSUBS 0.008001f
C296 B.n192 VSUBS 0.008001f
C297 B.n193 VSUBS 0.008001f
C298 B.n194 VSUBS 0.008001f
C299 B.n195 VSUBS 0.008001f
C300 B.n196 VSUBS 0.008001f
C301 B.n197 VSUBS 0.008001f
C302 B.n198 VSUBS 0.008001f
C303 B.n199 VSUBS 0.008001f
C304 B.n200 VSUBS 0.008001f
C305 B.n201 VSUBS 0.008001f
C306 B.n202 VSUBS 0.008001f
C307 B.n203 VSUBS 0.008001f
C308 B.n204 VSUBS 0.018132f
C309 B.n205 VSUBS 0.018132f
C310 B.n206 VSUBS 0.018815f
C311 B.n207 VSUBS 0.008001f
C312 B.n208 VSUBS 0.008001f
C313 B.n209 VSUBS 0.008001f
C314 B.n210 VSUBS 0.008001f
C315 B.n211 VSUBS 0.008001f
C316 B.n212 VSUBS 0.008001f
C317 B.n213 VSUBS 0.008001f
C318 B.n214 VSUBS 0.008001f
C319 B.n215 VSUBS 0.008001f
C320 B.n216 VSUBS 0.008001f
C321 B.n217 VSUBS 0.008001f
C322 B.n218 VSUBS 0.008001f
C323 B.n219 VSUBS 0.008001f
C324 B.n220 VSUBS 0.008001f
C325 B.n221 VSUBS 0.008001f
C326 B.n222 VSUBS 0.008001f
C327 B.n223 VSUBS 0.008001f
C328 B.n224 VSUBS 0.008001f
C329 B.n225 VSUBS 0.008001f
C330 B.n226 VSUBS 0.008001f
C331 B.n227 VSUBS 0.008001f
C332 B.n228 VSUBS 0.008001f
C333 B.n229 VSUBS 0.008001f
C334 B.n230 VSUBS 0.008001f
C335 B.n231 VSUBS 0.008001f
C336 B.n232 VSUBS 0.008001f
C337 B.n233 VSUBS 0.008001f
C338 B.n234 VSUBS 0.008001f
C339 B.n235 VSUBS 0.008001f
C340 B.n236 VSUBS 0.008001f
C341 B.n237 VSUBS 0.008001f
C342 B.n238 VSUBS 0.008001f
C343 B.n239 VSUBS 0.008001f
C344 B.n240 VSUBS 0.008001f
C345 B.n241 VSUBS 0.008001f
C346 B.n242 VSUBS 0.008001f
C347 B.n243 VSUBS 0.008001f
C348 B.n244 VSUBS 0.008001f
C349 B.n245 VSUBS 0.008001f
C350 B.n246 VSUBS 0.008001f
C351 B.n247 VSUBS 0.008001f
C352 B.n248 VSUBS 0.008001f
C353 B.n249 VSUBS 0.007531f
C354 B.n250 VSUBS 0.008001f
C355 B.n251 VSUBS 0.008001f
C356 B.n252 VSUBS 0.004471f
C357 B.n253 VSUBS 0.008001f
C358 B.n254 VSUBS 0.008001f
C359 B.n255 VSUBS 0.008001f
C360 B.n256 VSUBS 0.008001f
C361 B.n257 VSUBS 0.008001f
C362 B.n258 VSUBS 0.008001f
C363 B.n259 VSUBS 0.008001f
C364 B.n260 VSUBS 0.008001f
C365 B.n261 VSUBS 0.008001f
C366 B.n262 VSUBS 0.008001f
C367 B.n263 VSUBS 0.008001f
C368 B.n264 VSUBS 0.008001f
C369 B.n265 VSUBS 0.004471f
C370 B.n266 VSUBS 0.018538f
C371 B.n267 VSUBS 0.007531f
C372 B.n268 VSUBS 0.008001f
C373 B.n269 VSUBS 0.008001f
C374 B.n270 VSUBS 0.008001f
C375 B.n271 VSUBS 0.008001f
C376 B.n272 VSUBS 0.008001f
C377 B.n273 VSUBS 0.008001f
C378 B.n274 VSUBS 0.008001f
C379 B.n275 VSUBS 0.008001f
C380 B.n276 VSUBS 0.008001f
C381 B.n277 VSUBS 0.008001f
C382 B.n278 VSUBS 0.008001f
C383 B.n279 VSUBS 0.008001f
C384 B.n280 VSUBS 0.008001f
C385 B.n281 VSUBS 0.008001f
C386 B.n282 VSUBS 0.008001f
C387 B.n283 VSUBS 0.008001f
C388 B.n284 VSUBS 0.008001f
C389 B.n285 VSUBS 0.008001f
C390 B.n286 VSUBS 0.008001f
C391 B.n287 VSUBS 0.008001f
C392 B.n288 VSUBS 0.008001f
C393 B.n289 VSUBS 0.008001f
C394 B.n290 VSUBS 0.008001f
C395 B.n291 VSUBS 0.008001f
C396 B.n292 VSUBS 0.008001f
C397 B.n293 VSUBS 0.008001f
C398 B.n294 VSUBS 0.008001f
C399 B.n295 VSUBS 0.008001f
C400 B.n296 VSUBS 0.008001f
C401 B.n297 VSUBS 0.008001f
C402 B.n298 VSUBS 0.008001f
C403 B.n299 VSUBS 0.008001f
C404 B.n300 VSUBS 0.008001f
C405 B.n301 VSUBS 0.008001f
C406 B.n302 VSUBS 0.008001f
C407 B.n303 VSUBS 0.008001f
C408 B.n304 VSUBS 0.008001f
C409 B.n305 VSUBS 0.008001f
C410 B.n306 VSUBS 0.008001f
C411 B.n307 VSUBS 0.008001f
C412 B.n308 VSUBS 0.008001f
C413 B.n309 VSUBS 0.008001f
C414 B.n310 VSUBS 0.008001f
C415 B.n311 VSUBS 0.018815f
C416 B.n312 VSUBS 0.018132f
C417 B.n313 VSUBS 0.018132f
C418 B.n314 VSUBS 0.008001f
C419 B.n315 VSUBS 0.008001f
C420 B.n316 VSUBS 0.008001f
C421 B.n317 VSUBS 0.008001f
C422 B.n318 VSUBS 0.008001f
C423 B.n319 VSUBS 0.008001f
C424 B.n320 VSUBS 0.008001f
C425 B.n321 VSUBS 0.008001f
C426 B.n322 VSUBS 0.008001f
C427 B.n323 VSUBS 0.008001f
C428 B.n324 VSUBS 0.008001f
C429 B.n325 VSUBS 0.008001f
C430 B.n326 VSUBS 0.008001f
C431 B.n327 VSUBS 0.008001f
C432 B.n328 VSUBS 0.008001f
C433 B.n329 VSUBS 0.008001f
C434 B.n330 VSUBS 0.008001f
C435 B.n331 VSUBS 0.008001f
C436 B.n332 VSUBS 0.008001f
C437 B.n333 VSUBS 0.008001f
C438 B.n334 VSUBS 0.008001f
C439 B.n335 VSUBS 0.008001f
C440 B.n336 VSUBS 0.008001f
C441 B.n337 VSUBS 0.008001f
C442 B.n338 VSUBS 0.008001f
C443 B.n339 VSUBS 0.008001f
C444 B.n340 VSUBS 0.008001f
C445 B.n341 VSUBS 0.008001f
C446 B.n342 VSUBS 0.008001f
C447 B.n343 VSUBS 0.008001f
C448 B.n344 VSUBS 0.008001f
C449 B.n345 VSUBS 0.008001f
C450 B.n346 VSUBS 0.008001f
C451 B.n347 VSUBS 0.008001f
C452 B.n348 VSUBS 0.008001f
C453 B.n349 VSUBS 0.008001f
C454 B.n350 VSUBS 0.008001f
C455 B.n351 VSUBS 0.008001f
C456 B.n352 VSUBS 0.008001f
C457 B.n353 VSUBS 0.008001f
C458 B.n354 VSUBS 0.008001f
C459 B.n355 VSUBS 0.008001f
C460 B.n356 VSUBS 0.008001f
C461 B.n357 VSUBS 0.008001f
C462 B.n358 VSUBS 0.008001f
C463 B.n359 VSUBS 0.008001f
C464 B.n360 VSUBS 0.008001f
C465 B.n361 VSUBS 0.008001f
C466 B.n362 VSUBS 0.008001f
C467 B.n363 VSUBS 0.008001f
C468 B.n364 VSUBS 0.008001f
C469 B.n365 VSUBS 0.008001f
C470 B.n366 VSUBS 0.008001f
C471 B.n367 VSUBS 0.008001f
C472 B.n368 VSUBS 0.008001f
C473 B.n369 VSUBS 0.008001f
C474 B.n370 VSUBS 0.008001f
C475 B.n371 VSUBS 0.008001f
C476 B.n372 VSUBS 0.008001f
C477 B.n373 VSUBS 0.008001f
C478 B.n374 VSUBS 0.008001f
C479 B.n375 VSUBS 0.008001f
C480 B.n376 VSUBS 0.008001f
C481 B.n377 VSUBS 0.008001f
C482 B.n378 VSUBS 0.008001f
C483 B.n379 VSUBS 0.008001f
C484 B.n380 VSUBS 0.008001f
C485 B.n381 VSUBS 0.008001f
C486 B.n382 VSUBS 0.008001f
C487 B.n383 VSUBS 0.008001f
C488 B.n384 VSUBS 0.008001f
C489 B.n385 VSUBS 0.008001f
C490 B.n386 VSUBS 0.008001f
C491 B.n387 VSUBS 0.008001f
C492 B.n388 VSUBS 0.008001f
C493 B.n389 VSUBS 0.008001f
C494 B.n390 VSUBS 0.008001f
C495 B.n391 VSUBS 0.008001f
C496 B.n392 VSUBS 0.008001f
C497 B.n393 VSUBS 0.008001f
C498 B.n394 VSUBS 0.008001f
C499 B.n395 VSUBS 0.008001f
C500 B.n396 VSUBS 0.008001f
C501 B.n397 VSUBS 0.008001f
C502 B.n398 VSUBS 0.008001f
C503 B.n399 VSUBS 0.008001f
C504 B.n400 VSUBS 0.008001f
C505 B.n401 VSUBS 0.008001f
C506 B.n402 VSUBS 0.008001f
C507 B.n403 VSUBS 0.008001f
C508 B.n404 VSUBS 0.008001f
C509 B.n405 VSUBS 0.008001f
C510 B.n406 VSUBS 0.008001f
C511 B.n407 VSUBS 0.008001f
C512 B.n408 VSUBS 0.008001f
C513 B.n409 VSUBS 0.008001f
C514 B.n410 VSUBS 0.008001f
C515 B.n411 VSUBS 0.008001f
C516 B.n412 VSUBS 0.008001f
C517 B.n413 VSUBS 0.008001f
C518 B.n414 VSUBS 0.008001f
C519 B.n415 VSUBS 0.008001f
C520 B.n416 VSUBS 0.008001f
C521 B.n417 VSUBS 0.008001f
C522 B.n418 VSUBS 0.008001f
C523 B.n419 VSUBS 0.008001f
C524 B.n420 VSUBS 0.018132f
C525 B.n421 VSUBS 0.019097f
C526 B.n422 VSUBS 0.01785f
C527 B.n423 VSUBS 0.008001f
C528 B.n424 VSUBS 0.008001f
C529 B.n425 VSUBS 0.008001f
C530 B.n426 VSUBS 0.008001f
C531 B.n427 VSUBS 0.008001f
C532 B.n428 VSUBS 0.008001f
C533 B.n429 VSUBS 0.008001f
C534 B.n430 VSUBS 0.008001f
C535 B.n431 VSUBS 0.008001f
C536 B.n432 VSUBS 0.008001f
C537 B.n433 VSUBS 0.008001f
C538 B.n434 VSUBS 0.008001f
C539 B.n435 VSUBS 0.008001f
C540 B.n436 VSUBS 0.008001f
C541 B.n437 VSUBS 0.008001f
C542 B.n438 VSUBS 0.008001f
C543 B.n439 VSUBS 0.008001f
C544 B.n440 VSUBS 0.008001f
C545 B.n441 VSUBS 0.008001f
C546 B.n442 VSUBS 0.008001f
C547 B.n443 VSUBS 0.008001f
C548 B.n444 VSUBS 0.008001f
C549 B.n445 VSUBS 0.008001f
C550 B.n446 VSUBS 0.008001f
C551 B.n447 VSUBS 0.008001f
C552 B.n448 VSUBS 0.008001f
C553 B.n449 VSUBS 0.008001f
C554 B.n450 VSUBS 0.008001f
C555 B.n451 VSUBS 0.008001f
C556 B.n452 VSUBS 0.008001f
C557 B.n453 VSUBS 0.008001f
C558 B.n454 VSUBS 0.008001f
C559 B.n455 VSUBS 0.008001f
C560 B.n456 VSUBS 0.008001f
C561 B.n457 VSUBS 0.008001f
C562 B.n458 VSUBS 0.008001f
C563 B.n459 VSUBS 0.008001f
C564 B.n460 VSUBS 0.008001f
C565 B.n461 VSUBS 0.008001f
C566 B.n462 VSUBS 0.008001f
C567 B.n463 VSUBS 0.008001f
C568 B.n464 VSUBS 0.008001f
C569 B.n465 VSUBS 0.007531f
C570 B.n466 VSUBS 0.008001f
C571 B.n467 VSUBS 0.008001f
C572 B.n468 VSUBS 0.004471f
C573 B.n469 VSUBS 0.008001f
C574 B.n470 VSUBS 0.008001f
C575 B.n471 VSUBS 0.008001f
C576 B.n472 VSUBS 0.008001f
C577 B.n473 VSUBS 0.008001f
C578 B.n474 VSUBS 0.008001f
C579 B.n475 VSUBS 0.008001f
C580 B.n476 VSUBS 0.008001f
C581 B.n477 VSUBS 0.008001f
C582 B.n478 VSUBS 0.008001f
C583 B.n479 VSUBS 0.008001f
C584 B.n480 VSUBS 0.008001f
C585 B.n481 VSUBS 0.004471f
C586 B.n482 VSUBS 0.018538f
C587 B.n483 VSUBS 0.007531f
C588 B.n484 VSUBS 0.008001f
C589 B.n485 VSUBS 0.008001f
C590 B.n486 VSUBS 0.008001f
C591 B.n487 VSUBS 0.008001f
C592 B.n488 VSUBS 0.008001f
C593 B.n489 VSUBS 0.008001f
C594 B.n490 VSUBS 0.008001f
C595 B.n491 VSUBS 0.008001f
C596 B.n492 VSUBS 0.008001f
C597 B.n493 VSUBS 0.008001f
C598 B.n494 VSUBS 0.008001f
C599 B.n495 VSUBS 0.008001f
C600 B.n496 VSUBS 0.008001f
C601 B.n497 VSUBS 0.008001f
C602 B.n498 VSUBS 0.008001f
C603 B.n499 VSUBS 0.008001f
C604 B.n500 VSUBS 0.008001f
C605 B.n501 VSUBS 0.008001f
C606 B.n502 VSUBS 0.008001f
C607 B.n503 VSUBS 0.008001f
C608 B.n504 VSUBS 0.008001f
C609 B.n505 VSUBS 0.008001f
C610 B.n506 VSUBS 0.008001f
C611 B.n507 VSUBS 0.008001f
C612 B.n508 VSUBS 0.008001f
C613 B.n509 VSUBS 0.008001f
C614 B.n510 VSUBS 0.008001f
C615 B.n511 VSUBS 0.008001f
C616 B.n512 VSUBS 0.008001f
C617 B.n513 VSUBS 0.008001f
C618 B.n514 VSUBS 0.008001f
C619 B.n515 VSUBS 0.008001f
C620 B.n516 VSUBS 0.008001f
C621 B.n517 VSUBS 0.008001f
C622 B.n518 VSUBS 0.008001f
C623 B.n519 VSUBS 0.008001f
C624 B.n520 VSUBS 0.008001f
C625 B.n521 VSUBS 0.008001f
C626 B.n522 VSUBS 0.008001f
C627 B.n523 VSUBS 0.008001f
C628 B.n524 VSUBS 0.008001f
C629 B.n525 VSUBS 0.008001f
C630 B.n526 VSUBS 0.008001f
C631 B.n527 VSUBS 0.018815f
C632 B.n528 VSUBS 0.018132f
C633 B.n529 VSUBS 0.018132f
C634 B.n530 VSUBS 0.008001f
C635 B.n531 VSUBS 0.008001f
C636 B.n532 VSUBS 0.008001f
C637 B.n533 VSUBS 0.008001f
C638 B.n534 VSUBS 0.008001f
C639 B.n535 VSUBS 0.008001f
C640 B.n536 VSUBS 0.008001f
C641 B.n537 VSUBS 0.008001f
C642 B.n538 VSUBS 0.008001f
C643 B.n539 VSUBS 0.008001f
C644 B.n540 VSUBS 0.008001f
C645 B.n541 VSUBS 0.008001f
C646 B.n542 VSUBS 0.008001f
C647 B.n543 VSUBS 0.008001f
C648 B.n544 VSUBS 0.008001f
C649 B.n545 VSUBS 0.008001f
C650 B.n546 VSUBS 0.008001f
C651 B.n547 VSUBS 0.008001f
C652 B.n548 VSUBS 0.008001f
C653 B.n549 VSUBS 0.008001f
C654 B.n550 VSUBS 0.008001f
C655 B.n551 VSUBS 0.008001f
C656 B.n552 VSUBS 0.008001f
C657 B.n553 VSUBS 0.008001f
C658 B.n554 VSUBS 0.008001f
C659 B.n555 VSUBS 0.008001f
C660 B.n556 VSUBS 0.008001f
C661 B.n557 VSUBS 0.008001f
C662 B.n558 VSUBS 0.008001f
C663 B.n559 VSUBS 0.008001f
C664 B.n560 VSUBS 0.008001f
C665 B.n561 VSUBS 0.008001f
C666 B.n562 VSUBS 0.008001f
C667 B.n563 VSUBS 0.008001f
C668 B.n564 VSUBS 0.008001f
C669 B.n565 VSUBS 0.008001f
C670 B.n566 VSUBS 0.008001f
C671 B.n567 VSUBS 0.008001f
C672 B.n568 VSUBS 0.008001f
C673 B.n569 VSUBS 0.008001f
C674 B.n570 VSUBS 0.008001f
C675 B.n571 VSUBS 0.008001f
C676 B.n572 VSUBS 0.008001f
C677 B.n573 VSUBS 0.008001f
C678 B.n574 VSUBS 0.008001f
C679 B.n575 VSUBS 0.008001f
C680 B.n576 VSUBS 0.008001f
C681 B.n577 VSUBS 0.008001f
C682 B.n578 VSUBS 0.008001f
C683 B.n579 VSUBS 0.008001f
C684 B.n580 VSUBS 0.008001f
C685 B.n581 VSUBS 0.008001f
C686 B.n582 VSUBS 0.008001f
C687 B.n583 VSUBS 0.018117f
C688 VTAIL.t1 VSUBS 0.167219f
C689 VTAIL.t0 VSUBS 0.167219f
C690 VTAIL.n0 VSUBS 1.08074f
C691 VTAIL.n1 VSUBS 0.682544f
C692 VTAIL.n2 VSUBS 0.029557f
C693 VTAIL.n3 VSUBS 0.025996f
C694 VTAIL.n4 VSUBS 0.013969f
C695 VTAIL.n5 VSUBS 0.033018f
C696 VTAIL.n6 VSUBS 0.014791f
C697 VTAIL.n7 VSUBS 0.025996f
C698 VTAIL.n8 VSUBS 0.013969f
C699 VTAIL.n9 VSUBS 0.033018f
C700 VTAIL.n10 VSUBS 0.014791f
C701 VTAIL.n11 VSUBS 0.025996f
C702 VTAIL.n12 VSUBS 0.013969f
C703 VTAIL.n13 VSUBS 0.033018f
C704 VTAIL.n14 VSUBS 0.014791f
C705 VTAIL.n15 VSUBS 0.130831f
C706 VTAIL.t2 VSUBS 0.070426f
C707 VTAIL.n16 VSUBS 0.024764f
C708 VTAIL.n17 VSUBS 0.021004f
C709 VTAIL.n18 VSUBS 0.013969f
C710 VTAIL.n19 VSUBS 0.849952f
C711 VTAIL.n20 VSUBS 0.025996f
C712 VTAIL.n21 VSUBS 0.013969f
C713 VTAIL.n22 VSUBS 0.014791f
C714 VTAIL.n23 VSUBS 0.033018f
C715 VTAIL.n24 VSUBS 0.033018f
C716 VTAIL.n25 VSUBS 0.014791f
C717 VTAIL.n26 VSUBS 0.013969f
C718 VTAIL.n27 VSUBS 0.025996f
C719 VTAIL.n28 VSUBS 0.025996f
C720 VTAIL.n29 VSUBS 0.013969f
C721 VTAIL.n30 VSUBS 0.014791f
C722 VTAIL.n31 VSUBS 0.033018f
C723 VTAIL.n32 VSUBS 0.033018f
C724 VTAIL.n33 VSUBS 0.014791f
C725 VTAIL.n34 VSUBS 0.013969f
C726 VTAIL.n35 VSUBS 0.025996f
C727 VTAIL.n36 VSUBS 0.025996f
C728 VTAIL.n37 VSUBS 0.013969f
C729 VTAIL.n38 VSUBS 0.014791f
C730 VTAIL.n39 VSUBS 0.033018f
C731 VTAIL.n40 VSUBS 0.083316f
C732 VTAIL.n41 VSUBS 0.014791f
C733 VTAIL.n42 VSUBS 0.013969f
C734 VTAIL.n43 VSUBS 0.059378f
C735 VTAIL.n44 VSUBS 0.042027f
C736 VTAIL.n45 VSUBS 0.197636f
C737 VTAIL.n46 VSUBS 0.029557f
C738 VTAIL.n47 VSUBS 0.025996f
C739 VTAIL.n48 VSUBS 0.013969f
C740 VTAIL.n49 VSUBS 0.033018f
C741 VTAIL.n50 VSUBS 0.014791f
C742 VTAIL.n51 VSUBS 0.025996f
C743 VTAIL.n52 VSUBS 0.013969f
C744 VTAIL.n53 VSUBS 0.033018f
C745 VTAIL.n54 VSUBS 0.014791f
C746 VTAIL.n55 VSUBS 0.025996f
C747 VTAIL.n56 VSUBS 0.013969f
C748 VTAIL.n57 VSUBS 0.033018f
C749 VTAIL.n58 VSUBS 0.014791f
C750 VTAIL.n59 VSUBS 0.130831f
C751 VTAIL.t12 VSUBS 0.070426f
C752 VTAIL.n60 VSUBS 0.024764f
C753 VTAIL.n61 VSUBS 0.021004f
C754 VTAIL.n62 VSUBS 0.013969f
C755 VTAIL.n63 VSUBS 0.849952f
C756 VTAIL.n64 VSUBS 0.025996f
C757 VTAIL.n65 VSUBS 0.013969f
C758 VTAIL.n66 VSUBS 0.014791f
C759 VTAIL.n67 VSUBS 0.033018f
C760 VTAIL.n68 VSUBS 0.033018f
C761 VTAIL.n69 VSUBS 0.014791f
C762 VTAIL.n70 VSUBS 0.013969f
C763 VTAIL.n71 VSUBS 0.025996f
C764 VTAIL.n72 VSUBS 0.025996f
C765 VTAIL.n73 VSUBS 0.013969f
C766 VTAIL.n74 VSUBS 0.014791f
C767 VTAIL.n75 VSUBS 0.033018f
C768 VTAIL.n76 VSUBS 0.033018f
C769 VTAIL.n77 VSUBS 0.014791f
C770 VTAIL.n78 VSUBS 0.013969f
C771 VTAIL.n79 VSUBS 0.025996f
C772 VTAIL.n80 VSUBS 0.025996f
C773 VTAIL.n81 VSUBS 0.013969f
C774 VTAIL.n82 VSUBS 0.014791f
C775 VTAIL.n83 VSUBS 0.033018f
C776 VTAIL.n84 VSUBS 0.083316f
C777 VTAIL.n85 VSUBS 0.014791f
C778 VTAIL.n86 VSUBS 0.013969f
C779 VTAIL.n87 VSUBS 0.059378f
C780 VTAIL.n88 VSUBS 0.042027f
C781 VTAIL.n89 VSUBS 0.197636f
C782 VTAIL.t8 VSUBS 0.167219f
C783 VTAIL.t15 VSUBS 0.167219f
C784 VTAIL.n90 VSUBS 1.08074f
C785 VTAIL.n91 VSUBS 0.814149f
C786 VTAIL.n92 VSUBS 0.029557f
C787 VTAIL.n93 VSUBS 0.025996f
C788 VTAIL.n94 VSUBS 0.013969f
C789 VTAIL.n95 VSUBS 0.033018f
C790 VTAIL.n96 VSUBS 0.014791f
C791 VTAIL.n97 VSUBS 0.025996f
C792 VTAIL.n98 VSUBS 0.013969f
C793 VTAIL.n99 VSUBS 0.033018f
C794 VTAIL.n100 VSUBS 0.014791f
C795 VTAIL.n101 VSUBS 0.025996f
C796 VTAIL.n102 VSUBS 0.013969f
C797 VTAIL.n103 VSUBS 0.033018f
C798 VTAIL.n104 VSUBS 0.014791f
C799 VTAIL.n105 VSUBS 0.130831f
C800 VTAIL.t13 VSUBS 0.070426f
C801 VTAIL.n106 VSUBS 0.024764f
C802 VTAIL.n107 VSUBS 0.021004f
C803 VTAIL.n108 VSUBS 0.013969f
C804 VTAIL.n109 VSUBS 0.849952f
C805 VTAIL.n110 VSUBS 0.025996f
C806 VTAIL.n111 VSUBS 0.013969f
C807 VTAIL.n112 VSUBS 0.014791f
C808 VTAIL.n113 VSUBS 0.033018f
C809 VTAIL.n114 VSUBS 0.033018f
C810 VTAIL.n115 VSUBS 0.014791f
C811 VTAIL.n116 VSUBS 0.013969f
C812 VTAIL.n117 VSUBS 0.025996f
C813 VTAIL.n118 VSUBS 0.025996f
C814 VTAIL.n119 VSUBS 0.013969f
C815 VTAIL.n120 VSUBS 0.014791f
C816 VTAIL.n121 VSUBS 0.033018f
C817 VTAIL.n122 VSUBS 0.033018f
C818 VTAIL.n123 VSUBS 0.014791f
C819 VTAIL.n124 VSUBS 0.013969f
C820 VTAIL.n125 VSUBS 0.025996f
C821 VTAIL.n126 VSUBS 0.025996f
C822 VTAIL.n127 VSUBS 0.013969f
C823 VTAIL.n128 VSUBS 0.014791f
C824 VTAIL.n129 VSUBS 0.033018f
C825 VTAIL.n130 VSUBS 0.083316f
C826 VTAIL.n131 VSUBS 0.014791f
C827 VTAIL.n132 VSUBS 0.013969f
C828 VTAIL.n133 VSUBS 0.059378f
C829 VTAIL.n134 VSUBS 0.042027f
C830 VTAIL.n135 VSUBS 1.23569f
C831 VTAIL.n136 VSUBS 0.029557f
C832 VTAIL.n137 VSUBS 0.025996f
C833 VTAIL.n138 VSUBS 0.013969f
C834 VTAIL.n139 VSUBS 0.033018f
C835 VTAIL.n140 VSUBS 0.014791f
C836 VTAIL.n141 VSUBS 0.025996f
C837 VTAIL.n142 VSUBS 0.013969f
C838 VTAIL.n143 VSUBS 0.033018f
C839 VTAIL.n144 VSUBS 0.014791f
C840 VTAIL.n145 VSUBS 0.025996f
C841 VTAIL.n146 VSUBS 0.013969f
C842 VTAIL.n147 VSUBS 0.033018f
C843 VTAIL.n148 VSUBS 0.014791f
C844 VTAIL.n149 VSUBS 0.130831f
C845 VTAIL.t7 VSUBS 0.070426f
C846 VTAIL.n150 VSUBS 0.024764f
C847 VTAIL.n151 VSUBS 0.021004f
C848 VTAIL.n152 VSUBS 0.013969f
C849 VTAIL.n153 VSUBS 0.849952f
C850 VTAIL.n154 VSUBS 0.025996f
C851 VTAIL.n155 VSUBS 0.013969f
C852 VTAIL.n156 VSUBS 0.014791f
C853 VTAIL.n157 VSUBS 0.033018f
C854 VTAIL.n158 VSUBS 0.033018f
C855 VTAIL.n159 VSUBS 0.014791f
C856 VTAIL.n160 VSUBS 0.013969f
C857 VTAIL.n161 VSUBS 0.025996f
C858 VTAIL.n162 VSUBS 0.025996f
C859 VTAIL.n163 VSUBS 0.013969f
C860 VTAIL.n164 VSUBS 0.014791f
C861 VTAIL.n165 VSUBS 0.033018f
C862 VTAIL.n166 VSUBS 0.033018f
C863 VTAIL.n167 VSUBS 0.014791f
C864 VTAIL.n168 VSUBS 0.013969f
C865 VTAIL.n169 VSUBS 0.025996f
C866 VTAIL.n170 VSUBS 0.025996f
C867 VTAIL.n171 VSUBS 0.013969f
C868 VTAIL.n172 VSUBS 0.014791f
C869 VTAIL.n173 VSUBS 0.033018f
C870 VTAIL.n174 VSUBS 0.083316f
C871 VTAIL.n175 VSUBS 0.014791f
C872 VTAIL.n176 VSUBS 0.013969f
C873 VTAIL.n177 VSUBS 0.059378f
C874 VTAIL.n178 VSUBS 0.042027f
C875 VTAIL.n179 VSUBS 1.23569f
C876 VTAIL.t6 VSUBS 0.167219f
C877 VTAIL.t4 VSUBS 0.167219f
C878 VTAIL.n180 VSUBS 1.08074f
C879 VTAIL.n181 VSUBS 0.814141f
C880 VTAIL.n182 VSUBS 0.029557f
C881 VTAIL.n183 VSUBS 0.025996f
C882 VTAIL.n184 VSUBS 0.013969f
C883 VTAIL.n185 VSUBS 0.033018f
C884 VTAIL.n186 VSUBS 0.014791f
C885 VTAIL.n187 VSUBS 0.025996f
C886 VTAIL.n188 VSUBS 0.013969f
C887 VTAIL.n189 VSUBS 0.033018f
C888 VTAIL.n190 VSUBS 0.014791f
C889 VTAIL.n191 VSUBS 0.025996f
C890 VTAIL.n192 VSUBS 0.013969f
C891 VTAIL.n193 VSUBS 0.033018f
C892 VTAIL.n194 VSUBS 0.014791f
C893 VTAIL.n195 VSUBS 0.130831f
C894 VTAIL.t5 VSUBS 0.070426f
C895 VTAIL.n196 VSUBS 0.024764f
C896 VTAIL.n197 VSUBS 0.021004f
C897 VTAIL.n198 VSUBS 0.013969f
C898 VTAIL.n199 VSUBS 0.849952f
C899 VTAIL.n200 VSUBS 0.025996f
C900 VTAIL.n201 VSUBS 0.013969f
C901 VTAIL.n202 VSUBS 0.014791f
C902 VTAIL.n203 VSUBS 0.033018f
C903 VTAIL.n204 VSUBS 0.033018f
C904 VTAIL.n205 VSUBS 0.014791f
C905 VTAIL.n206 VSUBS 0.013969f
C906 VTAIL.n207 VSUBS 0.025996f
C907 VTAIL.n208 VSUBS 0.025996f
C908 VTAIL.n209 VSUBS 0.013969f
C909 VTAIL.n210 VSUBS 0.014791f
C910 VTAIL.n211 VSUBS 0.033018f
C911 VTAIL.n212 VSUBS 0.033018f
C912 VTAIL.n213 VSUBS 0.014791f
C913 VTAIL.n214 VSUBS 0.013969f
C914 VTAIL.n215 VSUBS 0.025996f
C915 VTAIL.n216 VSUBS 0.025996f
C916 VTAIL.n217 VSUBS 0.013969f
C917 VTAIL.n218 VSUBS 0.014791f
C918 VTAIL.n219 VSUBS 0.033018f
C919 VTAIL.n220 VSUBS 0.083316f
C920 VTAIL.n221 VSUBS 0.014791f
C921 VTAIL.n222 VSUBS 0.013969f
C922 VTAIL.n223 VSUBS 0.059378f
C923 VTAIL.n224 VSUBS 0.042027f
C924 VTAIL.n225 VSUBS 0.197636f
C925 VTAIL.n226 VSUBS 0.029557f
C926 VTAIL.n227 VSUBS 0.025996f
C927 VTAIL.n228 VSUBS 0.013969f
C928 VTAIL.n229 VSUBS 0.033018f
C929 VTAIL.n230 VSUBS 0.014791f
C930 VTAIL.n231 VSUBS 0.025996f
C931 VTAIL.n232 VSUBS 0.013969f
C932 VTAIL.n233 VSUBS 0.033018f
C933 VTAIL.n234 VSUBS 0.014791f
C934 VTAIL.n235 VSUBS 0.025996f
C935 VTAIL.n236 VSUBS 0.013969f
C936 VTAIL.n237 VSUBS 0.033018f
C937 VTAIL.n238 VSUBS 0.014791f
C938 VTAIL.n239 VSUBS 0.130831f
C939 VTAIL.t9 VSUBS 0.070426f
C940 VTAIL.n240 VSUBS 0.024764f
C941 VTAIL.n241 VSUBS 0.021004f
C942 VTAIL.n242 VSUBS 0.013969f
C943 VTAIL.n243 VSUBS 0.849952f
C944 VTAIL.n244 VSUBS 0.025996f
C945 VTAIL.n245 VSUBS 0.013969f
C946 VTAIL.n246 VSUBS 0.014791f
C947 VTAIL.n247 VSUBS 0.033018f
C948 VTAIL.n248 VSUBS 0.033018f
C949 VTAIL.n249 VSUBS 0.014791f
C950 VTAIL.n250 VSUBS 0.013969f
C951 VTAIL.n251 VSUBS 0.025996f
C952 VTAIL.n252 VSUBS 0.025996f
C953 VTAIL.n253 VSUBS 0.013969f
C954 VTAIL.n254 VSUBS 0.014791f
C955 VTAIL.n255 VSUBS 0.033018f
C956 VTAIL.n256 VSUBS 0.033018f
C957 VTAIL.n257 VSUBS 0.014791f
C958 VTAIL.n258 VSUBS 0.013969f
C959 VTAIL.n259 VSUBS 0.025996f
C960 VTAIL.n260 VSUBS 0.025996f
C961 VTAIL.n261 VSUBS 0.013969f
C962 VTAIL.n262 VSUBS 0.014791f
C963 VTAIL.n263 VSUBS 0.033018f
C964 VTAIL.n264 VSUBS 0.083316f
C965 VTAIL.n265 VSUBS 0.014791f
C966 VTAIL.n266 VSUBS 0.013969f
C967 VTAIL.n267 VSUBS 0.059378f
C968 VTAIL.n268 VSUBS 0.042027f
C969 VTAIL.n269 VSUBS 0.197636f
C970 VTAIL.t10 VSUBS 0.167219f
C971 VTAIL.t11 VSUBS 0.167219f
C972 VTAIL.n270 VSUBS 1.08074f
C973 VTAIL.n271 VSUBS 0.814141f
C974 VTAIL.n272 VSUBS 0.029557f
C975 VTAIL.n273 VSUBS 0.025996f
C976 VTAIL.n274 VSUBS 0.013969f
C977 VTAIL.n275 VSUBS 0.033018f
C978 VTAIL.n276 VSUBS 0.014791f
C979 VTAIL.n277 VSUBS 0.025996f
C980 VTAIL.n278 VSUBS 0.013969f
C981 VTAIL.n279 VSUBS 0.033018f
C982 VTAIL.n280 VSUBS 0.014791f
C983 VTAIL.n281 VSUBS 0.025996f
C984 VTAIL.n282 VSUBS 0.013969f
C985 VTAIL.n283 VSUBS 0.033018f
C986 VTAIL.n284 VSUBS 0.014791f
C987 VTAIL.n285 VSUBS 0.130831f
C988 VTAIL.t14 VSUBS 0.070426f
C989 VTAIL.n286 VSUBS 0.024764f
C990 VTAIL.n287 VSUBS 0.021004f
C991 VTAIL.n288 VSUBS 0.013969f
C992 VTAIL.n289 VSUBS 0.849952f
C993 VTAIL.n290 VSUBS 0.025996f
C994 VTAIL.n291 VSUBS 0.013969f
C995 VTAIL.n292 VSUBS 0.014791f
C996 VTAIL.n293 VSUBS 0.033018f
C997 VTAIL.n294 VSUBS 0.033018f
C998 VTAIL.n295 VSUBS 0.014791f
C999 VTAIL.n296 VSUBS 0.013969f
C1000 VTAIL.n297 VSUBS 0.025996f
C1001 VTAIL.n298 VSUBS 0.025996f
C1002 VTAIL.n299 VSUBS 0.013969f
C1003 VTAIL.n300 VSUBS 0.014791f
C1004 VTAIL.n301 VSUBS 0.033018f
C1005 VTAIL.n302 VSUBS 0.033018f
C1006 VTAIL.n303 VSUBS 0.014791f
C1007 VTAIL.n304 VSUBS 0.013969f
C1008 VTAIL.n305 VSUBS 0.025996f
C1009 VTAIL.n306 VSUBS 0.025996f
C1010 VTAIL.n307 VSUBS 0.013969f
C1011 VTAIL.n308 VSUBS 0.014791f
C1012 VTAIL.n309 VSUBS 0.033018f
C1013 VTAIL.n310 VSUBS 0.083316f
C1014 VTAIL.n311 VSUBS 0.014791f
C1015 VTAIL.n312 VSUBS 0.013969f
C1016 VTAIL.n313 VSUBS 0.059378f
C1017 VTAIL.n314 VSUBS 0.042027f
C1018 VTAIL.n315 VSUBS 1.23569f
C1019 VTAIL.n316 VSUBS 0.029557f
C1020 VTAIL.n317 VSUBS 0.025996f
C1021 VTAIL.n318 VSUBS 0.013969f
C1022 VTAIL.n319 VSUBS 0.033018f
C1023 VTAIL.n320 VSUBS 0.014791f
C1024 VTAIL.n321 VSUBS 0.025996f
C1025 VTAIL.n322 VSUBS 0.013969f
C1026 VTAIL.n323 VSUBS 0.033018f
C1027 VTAIL.n324 VSUBS 0.014791f
C1028 VTAIL.n325 VSUBS 0.025996f
C1029 VTAIL.n326 VSUBS 0.013969f
C1030 VTAIL.n327 VSUBS 0.033018f
C1031 VTAIL.n328 VSUBS 0.014791f
C1032 VTAIL.n329 VSUBS 0.130831f
C1033 VTAIL.t3 VSUBS 0.070426f
C1034 VTAIL.n330 VSUBS 0.024764f
C1035 VTAIL.n331 VSUBS 0.021004f
C1036 VTAIL.n332 VSUBS 0.013969f
C1037 VTAIL.n333 VSUBS 0.849952f
C1038 VTAIL.n334 VSUBS 0.025996f
C1039 VTAIL.n335 VSUBS 0.013969f
C1040 VTAIL.n336 VSUBS 0.014791f
C1041 VTAIL.n337 VSUBS 0.033018f
C1042 VTAIL.n338 VSUBS 0.033018f
C1043 VTAIL.n339 VSUBS 0.014791f
C1044 VTAIL.n340 VSUBS 0.013969f
C1045 VTAIL.n341 VSUBS 0.025996f
C1046 VTAIL.n342 VSUBS 0.025996f
C1047 VTAIL.n343 VSUBS 0.013969f
C1048 VTAIL.n344 VSUBS 0.014791f
C1049 VTAIL.n345 VSUBS 0.033018f
C1050 VTAIL.n346 VSUBS 0.033018f
C1051 VTAIL.n347 VSUBS 0.014791f
C1052 VTAIL.n348 VSUBS 0.013969f
C1053 VTAIL.n349 VSUBS 0.025996f
C1054 VTAIL.n350 VSUBS 0.025996f
C1055 VTAIL.n351 VSUBS 0.013969f
C1056 VTAIL.n352 VSUBS 0.014791f
C1057 VTAIL.n353 VSUBS 0.033018f
C1058 VTAIL.n354 VSUBS 0.083316f
C1059 VTAIL.n355 VSUBS 0.014791f
C1060 VTAIL.n356 VSUBS 0.013969f
C1061 VTAIL.n357 VSUBS 0.059378f
C1062 VTAIL.n358 VSUBS 0.042027f
C1063 VTAIL.n359 VSUBS 1.23081f
C1064 VDD1.t0 VSUBS 0.162045f
C1065 VDD1.t1 VSUBS 0.162045f
C1066 VDD1.n0 VSUBS 1.16633f
C1067 VDD1.t6 VSUBS 0.162045f
C1068 VDD1.t2 VSUBS 0.162045f
C1069 VDD1.n1 VSUBS 1.16536f
C1070 VDD1.t5 VSUBS 0.162045f
C1071 VDD1.t4 VSUBS 0.162045f
C1072 VDD1.n2 VSUBS 1.16536f
C1073 VDD1.n3 VSUBS 2.98599f
C1074 VDD1.t3 VSUBS 0.162045f
C1075 VDD1.t7 VSUBS 0.162045f
C1076 VDD1.n4 VSUBS 1.15942f
C1077 VDD1.n5 VSUBS 2.57602f
C1078 VP.n0 VSUBS 0.04283f
C1079 VP.t3 VSUBS 1.46177f
C1080 VP.n1 VSUBS 0.046916f
C1081 VP.n2 VSUBS 0.04283f
C1082 VP.t0 VSUBS 1.46177f
C1083 VP.n3 VSUBS 0.062796f
C1084 VP.n4 VSUBS 0.04283f
C1085 VP.t7 VSUBS 1.46177f
C1086 VP.n5 VSUBS 0.075436f
C1087 VP.n6 VSUBS 0.04283f
C1088 VP.t1 VSUBS 1.46177f
C1089 VP.n7 VSUBS 0.046916f
C1090 VP.n8 VSUBS 0.04283f
C1091 VP.t4 VSUBS 1.46177f
C1092 VP.n9 VSUBS 0.062796f
C1093 VP.t6 VSUBS 1.60124f
C1094 VP.n10 VSUBS 0.653093f
C1095 VP.t5 VSUBS 1.46177f
C1096 VP.n11 VSUBS 0.626399f
C1097 VP.n12 VSUBS 0.056062f
C1098 VP.n13 VSUBS 0.268864f
C1099 VP.n14 VSUBS 0.04283f
C1100 VP.n15 VSUBS 0.04283f
C1101 VP.n16 VSUBS 0.062796f
C1102 VP.n17 VSUBS 0.056062f
C1103 VP.n18 VSUBS 0.547671f
C1104 VP.n19 VSUBS 0.068017f
C1105 VP.n20 VSUBS 0.04283f
C1106 VP.n21 VSUBS 0.04283f
C1107 VP.n22 VSUBS 0.04283f
C1108 VP.n23 VSUBS 0.075436f
C1109 VP.n24 VSUBS 0.047348f
C1110 VP.n25 VSUBS 0.629174f
C1111 VP.n26 VSUBS 1.84514f
C1112 VP.n27 VSUBS 1.88088f
C1113 VP.t2 VSUBS 1.46177f
C1114 VP.n28 VSUBS 0.629174f
C1115 VP.n29 VSUBS 0.047348f
C1116 VP.n30 VSUBS 0.04283f
C1117 VP.n31 VSUBS 0.04283f
C1118 VP.n32 VSUBS 0.04283f
C1119 VP.n33 VSUBS 0.046916f
C1120 VP.n34 VSUBS 0.068017f
C1121 VP.n35 VSUBS 0.547671f
C1122 VP.n36 VSUBS 0.056062f
C1123 VP.n37 VSUBS 0.04283f
C1124 VP.n38 VSUBS 0.04283f
C1125 VP.n39 VSUBS 0.04283f
C1126 VP.n40 VSUBS 0.062796f
C1127 VP.n41 VSUBS 0.056062f
C1128 VP.n42 VSUBS 0.547671f
C1129 VP.n43 VSUBS 0.068017f
C1130 VP.n44 VSUBS 0.04283f
C1131 VP.n45 VSUBS 0.04283f
C1132 VP.n46 VSUBS 0.04283f
C1133 VP.n47 VSUBS 0.075436f
C1134 VP.n48 VSUBS 0.047348f
C1135 VP.n49 VSUBS 0.629174f
C1136 VP.n50 VSUBS 0.043401f
.ends

