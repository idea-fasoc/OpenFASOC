* NGSPICE file created from diff_pair_sample_1556.ext - technology: sky130A

.subckt diff_pair_sample_1556 VTAIL VN VP B VDD2 VDD1
X0 B.t17 B.t15 B.t16 B.t12 sky130_fd_pr__nfet_01v8 ad=0.6708 pd=4.22 as=0 ps=0 w=1.72 l=1.23
X1 VDD1.t3 VP.t0 VTAIL.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=0.2838 pd=2.05 as=0.6708 ps=4.22 w=1.72 l=1.23
X2 VTAIL.t7 VN.t0 VDD2.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=0.6708 pd=4.22 as=0.2838 ps=2.05 w=1.72 l=1.23
X3 VDD1.t2 VP.t1 VTAIL.t5 B.t0 sky130_fd_pr__nfet_01v8 ad=0.2838 pd=2.05 as=0.6708 ps=4.22 w=1.72 l=1.23
X4 B.t14 B.t11 B.t13 B.t12 sky130_fd_pr__nfet_01v8 ad=0.6708 pd=4.22 as=0 ps=0 w=1.72 l=1.23
X5 B.t10 B.t8 B.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=0.6708 pd=4.22 as=0 ps=0 w=1.72 l=1.23
X6 VDD2.t2 VN.t1 VTAIL.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=0.2838 pd=2.05 as=0.6708 ps=4.22 w=1.72 l=1.23
X7 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=0.6708 pd=4.22 as=0 ps=0 w=1.72 l=1.23
X8 VTAIL.t0 VN.t2 VDD2.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.6708 pd=4.22 as=0.2838 ps=2.05 w=1.72 l=1.23
X9 VDD2.t0 VN.t3 VTAIL.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=0.2838 pd=2.05 as=0.6708 ps=4.22 w=1.72 l=1.23
X10 VTAIL.t4 VP.t2 VDD1.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.6708 pd=4.22 as=0.2838 ps=2.05 w=1.72 l=1.23
X11 VTAIL.t3 VP.t3 VDD1.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=0.6708 pd=4.22 as=0.2838 ps=2.05 w=1.72 l=1.23
R0 B.n287 B.n286 585
R1 B.n289 B.n64 585
R2 B.n292 B.n291 585
R3 B.n293 B.n63 585
R4 B.n295 B.n294 585
R5 B.n297 B.n62 585
R6 B.n300 B.n299 585
R7 B.n301 B.n61 585
R8 B.n303 B.n302 585
R9 B.n305 B.n60 585
R10 B.n308 B.n307 585
R11 B.n310 B.n57 585
R12 B.n312 B.n311 585
R13 B.n314 B.n56 585
R14 B.n317 B.n316 585
R15 B.n318 B.n55 585
R16 B.n320 B.n319 585
R17 B.n322 B.n54 585
R18 B.n325 B.n324 585
R19 B.n326 B.n50 585
R20 B.n328 B.n327 585
R21 B.n330 B.n49 585
R22 B.n333 B.n332 585
R23 B.n334 B.n48 585
R24 B.n336 B.n335 585
R25 B.n338 B.n47 585
R26 B.n341 B.n340 585
R27 B.n342 B.n46 585
R28 B.n344 B.n343 585
R29 B.n346 B.n45 585
R30 B.n349 B.n348 585
R31 B.n350 B.n44 585
R32 B.n285 B.n42 585
R33 B.n353 B.n42 585
R34 B.n284 B.n41 585
R35 B.n354 B.n41 585
R36 B.n283 B.n40 585
R37 B.n355 B.n40 585
R38 B.n282 B.n281 585
R39 B.n281 B.n36 585
R40 B.n280 B.n35 585
R41 B.n361 B.n35 585
R42 B.n279 B.n34 585
R43 B.n362 B.n34 585
R44 B.n278 B.n33 585
R45 B.n363 B.n33 585
R46 B.n277 B.n276 585
R47 B.n276 B.n29 585
R48 B.n275 B.n28 585
R49 B.n369 B.n28 585
R50 B.n274 B.n27 585
R51 B.n370 B.n27 585
R52 B.n273 B.n26 585
R53 B.n371 B.n26 585
R54 B.n272 B.n271 585
R55 B.n271 B.n22 585
R56 B.n270 B.n21 585
R57 B.n377 B.n21 585
R58 B.n269 B.n20 585
R59 B.n378 B.n20 585
R60 B.n268 B.n19 585
R61 B.n379 B.n19 585
R62 B.n267 B.n266 585
R63 B.n266 B.n15 585
R64 B.n265 B.n14 585
R65 B.n385 B.n14 585
R66 B.n264 B.n13 585
R67 B.n386 B.n13 585
R68 B.n263 B.n12 585
R69 B.n387 B.n12 585
R70 B.n262 B.n261 585
R71 B.n261 B.n8 585
R72 B.n260 B.n7 585
R73 B.n393 B.n7 585
R74 B.n259 B.n6 585
R75 B.n394 B.n6 585
R76 B.n258 B.n5 585
R77 B.n395 B.n5 585
R78 B.n257 B.n256 585
R79 B.n256 B.n4 585
R80 B.n255 B.n65 585
R81 B.n255 B.n254 585
R82 B.n245 B.n66 585
R83 B.n67 B.n66 585
R84 B.n247 B.n246 585
R85 B.n248 B.n247 585
R86 B.n244 B.n72 585
R87 B.n72 B.n71 585
R88 B.n243 B.n242 585
R89 B.n242 B.n241 585
R90 B.n74 B.n73 585
R91 B.n75 B.n74 585
R92 B.n234 B.n233 585
R93 B.n235 B.n234 585
R94 B.n232 B.n79 585
R95 B.n83 B.n79 585
R96 B.n231 B.n230 585
R97 B.n230 B.n229 585
R98 B.n81 B.n80 585
R99 B.n82 B.n81 585
R100 B.n222 B.n221 585
R101 B.n223 B.n222 585
R102 B.n220 B.n88 585
R103 B.n88 B.n87 585
R104 B.n219 B.n218 585
R105 B.n218 B.n217 585
R106 B.n90 B.n89 585
R107 B.n91 B.n90 585
R108 B.n210 B.n209 585
R109 B.n211 B.n210 585
R110 B.n208 B.n95 585
R111 B.n99 B.n95 585
R112 B.n207 B.n206 585
R113 B.n206 B.n205 585
R114 B.n97 B.n96 585
R115 B.n98 B.n97 585
R116 B.n198 B.n197 585
R117 B.n199 B.n198 585
R118 B.n196 B.n104 585
R119 B.n104 B.n103 585
R120 B.n195 B.n194 585
R121 B.n194 B.n193 585
R122 B.n190 B.n108 585
R123 B.n189 B.n188 585
R124 B.n186 B.n109 585
R125 B.n186 B.n107 585
R126 B.n185 B.n184 585
R127 B.n183 B.n182 585
R128 B.n181 B.n111 585
R129 B.n179 B.n178 585
R130 B.n177 B.n112 585
R131 B.n176 B.n175 585
R132 B.n173 B.n113 585
R133 B.n171 B.n170 585
R134 B.n168 B.n114 585
R135 B.n167 B.n166 585
R136 B.n164 B.n117 585
R137 B.n162 B.n161 585
R138 B.n160 B.n118 585
R139 B.n159 B.n158 585
R140 B.n156 B.n119 585
R141 B.n154 B.n153 585
R142 B.n152 B.n120 585
R143 B.n151 B.n150 585
R144 B.n148 B.n147 585
R145 B.n146 B.n145 585
R146 B.n144 B.n125 585
R147 B.n142 B.n141 585
R148 B.n140 B.n126 585
R149 B.n139 B.n138 585
R150 B.n136 B.n127 585
R151 B.n134 B.n133 585
R152 B.n132 B.n128 585
R153 B.n131 B.n130 585
R154 B.n106 B.n105 585
R155 B.n107 B.n106 585
R156 B.n192 B.n191 585
R157 B.n193 B.n192 585
R158 B.n102 B.n101 585
R159 B.n103 B.n102 585
R160 B.n201 B.n200 585
R161 B.n200 B.n199 585
R162 B.n202 B.n100 585
R163 B.n100 B.n98 585
R164 B.n204 B.n203 585
R165 B.n205 B.n204 585
R166 B.n94 B.n93 585
R167 B.n99 B.n94 585
R168 B.n213 B.n212 585
R169 B.n212 B.n211 585
R170 B.n214 B.n92 585
R171 B.n92 B.n91 585
R172 B.n216 B.n215 585
R173 B.n217 B.n216 585
R174 B.n86 B.n85 585
R175 B.n87 B.n86 585
R176 B.n225 B.n224 585
R177 B.n224 B.n223 585
R178 B.n226 B.n84 585
R179 B.n84 B.n82 585
R180 B.n228 B.n227 585
R181 B.n229 B.n228 585
R182 B.n78 B.n77 585
R183 B.n83 B.n78 585
R184 B.n237 B.n236 585
R185 B.n236 B.n235 585
R186 B.n238 B.n76 585
R187 B.n76 B.n75 585
R188 B.n240 B.n239 585
R189 B.n241 B.n240 585
R190 B.n70 B.n69 585
R191 B.n71 B.n70 585
R192 B.n250 B.n249 585
R193 B.n249 B.n248 585
R194 B.n251 B.n68 585
R195 B.n68 B.n67 585
R196 B.n253 B.n252 585
R197 B.n254 B.n253 585
R198 B.n2 B.n0 585
R199 B.n4 B.n2 585
R200 B.n3 B.n1 585
R201 B.n394 B.n3 585
R202 B.n392 B.n391 585
R203 B.n393 B.n392 585
R204 B.n390 B.n9 585
R205 B.n9 B.n8 585
R206 B.n389 B.n388 585
R207 B.n388 B.n387 585
R208 B.n11 B.n10 585
R209 B.n386 B.n11 585
R210 B.n384 B.n383 585
R211 B.n385 B.n384 585
R212 B.n382 B.n16 585
R213 B.n16 B.n15 585
R214 B.n381 B.n380 585
R215 B.n380 B.n379 585
R216 B.n18 B.n17 585
R217 B.n378 B.n18 585
R218 B.n376 B.n375 585
R219 B.n377 B.n376 585
R220 B.n374 B.n23 585
R221 B.n23 B.n22 585
R222 B.n373 B.n372 585
R223 B.n372 B.n371 585
R224 B.n25 B.n24 585
R225 B.n370 B.n25 585
R226 B.n368 B.n367 585
R227 B.n369 B.n368 585
R228 B.n366 B.n30 585
R229 B.n30 B.n29 585
R230 B.n365 B.n364 585
R231 B.n364 B.n363 585
R232 B.n32 B.n31 585
R233 B.n362 B.n32 585
R234 B.n360 B.n359 585
R235 B.n361 B.n360 585
R236 B.n358 B.n37 585
R237 B.n37 B.n36 585
R238 B.n357 B.n356 585
R239 B.n356 B.n355 585
R240 B.n39 B.n38 585
R241 B.n354 B.n39 585
R242 B.n352 B.n351 585
R243 B.n353 B.n352 585
R244 B.n397 B.n396 585
R245 B.n396 B.n395 585
R246 B.n192 B.n108 506.916
R247 B.n352 B.n44 506.916
R248 B.n194 B.n106 506.916
R249 B.n287 B.n42 506.916
R250 B.n288 B.n43 256.663
R251 B.n290 B.n43 256.663
R252 B.n296 B.n43 256.663
R253 B.n298 B.n43 256.663
R254 B.n304 B.n43 256.663
R255 B.n306 B.n43 256.663
R256 B.n313 B.n43 256.663
R257 B.n315 B.n43 256.663
R258 B.n321 B.n43 256.663
R259 B.n323 B.n43 256.663
R260 B.n329 B.n43 256.663
R261 B.n331 B.n43 256.663
R262 B.n337 B.n43 256.663
R263 B.n339 B.n43 256.663
R264 B.n345 B.n43 256.663
R265 B.n347 B.n43 256.663
R266 B.n187 B.n107 256.663
R267 B.n110 B.n107 256.663
R268 B.n180 B.n107 256.663
R269 B.n174 B.n107 256.663
R270 B.n172 B.n107 256.663
R271 B.n165 B.n107 256.663
R272 B.n163 B.n107 256.663
R273 B.n157 B.n107 256.663
R274 B.n155 B.n107 256.663
R275 B.n149 B.n107 256.663
R276 B.n124 B.n107 256.663
R277 B.n143 B.n107 256.663
R278 B.n137 B.n107 256.663
R279 B.n135 B.n107 256.663
R280 B.n129 B.n107 256.663
R281 B.n121 B.t4 237.972
R282 B.n115 B.t8 237.972
R283 B.n51 B.t15 237.972
R284 B.n58 B.t11 237.972
R285 B.n193 B.n107 180.844
R286 B.n353 B.n43 180.844
R287 B.n192 B.n102 163.367
R288 B.n200 B.n102 163.367
R289 B.n200 B.n100 163.367
R290 B.n204 B.n100 163.367
R291 B.n204 B.n94 163.367
R292 B.n212 B.n94 163.367
R293 B.n212 B.n92 163.367
R294 B.n216 B.n92 163.367
R295 B.n216 B.n86 163.367
R296 B.n224 B.n86 163.367
R297 B.n224 B.n84 163.367
R298 B.n228 B.n84 163.367
R299 B.n228 B.n78 163.367
R300 B.n236 B.n78 163.367
R301 B.n236 B.n76 163.367
R302 B.n240 B.n76 163.367
R303 B.n240 B.n70 163.367
R304 B.n249 B.n70 163.367
R305 B.n249 B.n68 163.367
R306 B.n253 B.n68 163.367
R307 B.n253 B.n2 163.367
R308 B.n396 B.n2 163.367
R309 B.n396 B.n3 163.367
R310 B.n392 B.n3 163.367
R311 B.n392 B.n9 163.367
R312 B.n388 B.n9 163.367
R313 B.n388 B.n11 163.367
R314 B.n384 B.n11 163.367
R315 B.n384 B.n16 163.367
R316 B.n380 B.n16 163.367
R317 B.n380 B.n18 163.367
R318 B.n376 B.n18 163.367
R319 B.n376 B.n23 163.367
R320 B.n372 B.n23 163.367
R321 B.n372 B.n25 163.367
R322 B.n368 B.n25 163.367
R323 B.n368 B.n30 163.367
R324 B.n364 B.n30 163.367
R325 B.n364 B.n32 163.367
R326 B.n360 B.n32 163.367
R327 B.n360 B.n37 163.367
R328 B.n356 B.n37 163.367
R329 B.n356 B.n39 163.367
R330 B.n352 B.n39 163.367
R331 B.n188 B.n186 163.367
R332 B.n186 B.n185 163.367
R333 B.n182 B.n181 163.367
R334 B.n179 B.n112 163.367
R335 B.n175 B.n173 163.367
R336 B.n171 B.n114 163.367
R337 B.n166 B.n164 163.367
R338 B.n162 B.n118 163.367
R339 B.n158 B.n156 163.367
R340 B.n154 B.n120 163.367
R341 B.n150 B.n148 163.367
R342 B.n145 B.n144 163.367
R343 B.n142 B.n126 163.367
R344 B.n138 B.n136 163.367
R345 B.n134 B.n128 163.367
R346 B.n130 B.n106 163.367
R347 B.n194 B.n104 163.367
R348 B.n198 B.n104 163.367
R349 B.n198 B.n97 163.367
R350 B.n206 B.n97 163.367
R351 B.n206 B.n95 163.367
R352 B.n210 B.n95 163.367
R353 B.n210 B.n90 163.367
R354 B.n218 B.n90 163.367
R355 B.n218 B.n88 163.367
R356 B.n222 B.n88 163.367
R357 B.n222 B.n81 163.367
R358 B.n230 B.n81 163.367
R359 B.n230 B.n79 163.367
R360 B.n234 B.n79 163.367
R361 B.n234 B.n74 163.367
R362 B.n242 B.n74 163.367
R363 B.n242 B.n72 163.367
R364 B.n247 B.n72 163.367
R365 B.n247 B.n66 163.367
R366 B.n255 B.n66 163.367
R367 B.n256 B.n255 163.367
R368 B.n256 B.n5 163.367
R369 B.n6 B.n5 163.367
R370 B.n7 B.n6 163.367
R371 B.n261 B.n7 163.367
R372 B.n261 B.n12 163.367
R373 B.n13 B.n12 163.367
R374 B.n14 B.n13 163.367
R375 B.n266 B.n14 163.367
R376 B.n266 B.n19 163.367
R377 B.n20 B.n19 163.367
R378 B.n21 B.n20 163.367
R379 B.n271 B.n21 163.367
R380 B.n271 B.n26 163.367
R381 B.n27 B.n26 163.367
R382 B.n28 B.n27 163.367
R383 B.n276 B.n28 163.367
R384 B.n276 B.n33 163.367
R385 B.n34 B.n33 163.367
R386 B.n35 B.n34 163.367
R387 B.n281 B.n35 163.367
R388 B.n281 B.n40 163.367
R389 B.n41 B.n40 163.367
R390 B.n42 B.n41 163.367
R391 B.n348 B.n346 163.367
R392 B.n344 B.n46 163.367
R393 B.n340 B.n338 163.367
R394 B.n336 B.n48 163.367
R395 B.n332 B.n330 163.367
R396 B.n328 B.n50 163.367
R397 B.n324 B.n322 163.367
R398 B.n320 B.n55 163.367
R399 B.n316 B.n314 163.367
R400 B.n312 B.n57 163.367
R401 B.n307 B.n305 163.367
R402 B.n303 B.n61 163.367
R403 B.n299 B.n297 163.367
R404 B.n295 B.n63 163.367
R405 B.n291 B.n289 163.367
R406 B.n121 B.t7 147.843
R407 B.n58 B.t13 147.843
R408 B.n115 B.t10 147.843
R409 B.n51 B.t16 147.843
R410 B.n122 B.t6 117.588
R411 B.n59 B.t14 117.588
R412 B.n116 B.t9 117.588
R413 B.n52 B.t17 117.588
R414 B.n193 B.n103 106.934
R415 B.n199 B.n103 106.934
R416 B.n199 B.n98 106.934
R417 B.n205 B.n98 106.934
R418 B.n205 B.n99 106.934
R419 B.n211 B.n91 106.934
R420 B.n217 B.n91 106.934
R421 B.n217 B.n87 106.934
R422 B.n223 B.n87 106.934
R423 B.n223 B.n82 106.934
R424 B.n229 B.n82 106.934
R425 B.n229 B.n83 106.934
R426 B.n235 B.n75 106.934
R427 B.n241 B.n75 106.934
R428 B.n241 B.n71 106.934
R429 B.n248 B.n71 106.934
R430 B.n254 B.n67 106.934
R431 B.n254 B.n4 106.934
R432 B.n395 B.n4 106.934
R433 B.n395 B.n394 106.934
R434 B.n394 B.n393 106.934
R435 B.n393 B.n8 106.934
R436 B.n387 B.n386 106.934
R437 B.n386 B.n385 106.934
R438 B.n385 B.n15 106.934
R439 B.n379 B.n15 106.934
R440 B.n378 B.n377 106.934
R441 B.n377 B.n22 106.934
R442 B.n371 B.n22 106.934
R443 B.n371 B.n370 106.934
R444 B.n370 B.n369 106.934
R445 B.n369 B.n29 106.934
R446 B.n363 B.n29 106.934
R447 B.n362 B.n361 106.934
R448 B.n361 B.n36 106.934
R449 B.n355 B.n36 106.934
R450 B.n355 B.n354 106.934
R451 B.n354 B.n353 106.934
R452 B.t0 B.n67 95.9262
R453 B.t2 B.n8 95.9262
R454 B.n99 B.t5 77.0555
R455 B.t12 B.n362 77.0555
R456 B.n187 B.n108 71.676
R457 B.n185 B.n110 71.676
R458 B.n181 B.n180 71.676
R459 B.n174 B.n112 71.676
R460 B.n173 B.n172 71.676
R461 B.n165 B.n114 71.676
R462 B.n164 B.n163 71.676
R463 B.n157 B.n118 71.676
R464 B.n156 B.n155 71.676
R465 B.n149 B.n120 71.676
R466 B.n148 B.n124 71.676
R467 B.n144 B.n143 71.676
R468 B.n137 B.n126 71.676
R469 B.n136 B.n135 71.676
R470 B.n129 B.n128 71.676
R471 B.n347 B.n44 71.676
R472 B.n346 B.n345 71.676
R473 B.n339 B.n46 71.676
R474 B.n338 B.n337 71.676
R475 B.n331 B.n48 71.676
R476 B.n330 B.n329 71.676
R477 B.n323 B.n50 71.676
R478 B.n322 B.n321 71.676
R479 B.n315 B.n55 71.676
R480 B.n314 B.n313 71.676
R481 B.n306 B.n57 71.676
R482 B.n305 B.n304 71.676
R483 B.n298 B.n61 71.676
R484 B.n297 B.n296 71.676
R485 B.n290 B.n63 71.676
R486 B.n289 B.n288 71.676
R487 B.n288 B.n287 71.676
R488 B.n291 B.n290 71.676
R489 B.n296 B.n295 71.676
R490 B.n299 B.n298 71.676
R491 B.n304 B.n303 71.676
R492 B.n307 B.n306 71.676
R493 B.n313 B.n312 71.676
R494 B.n316 B.n315 71.676
R495 B.n321 B.n320 71.676
R496 B.n324 B.n323 71.676
R497 B.n329 B.n328 71.676
R498 B.n332 B.n331 71.676
R499 B.n337 B.n336 71.676
R500 B.n340 B.n339 71.676
R501 B.n345 B.n344 71.676
R502 B.n348 B.n347 71.676
R503 B.n188 B.n187 71.676
R504 B.n182 B.n110 71.676
R505 B.n180 B.n179 71.676
R506 B.n175 B.n174 71.676
R507 B.n172 B.n171 71.676
R508 B.n166 B.n165 71.676
R509 B.n163 B.n162 71.676
R510 B.n158 B.n157 71.676
R511 B.n155 B.n154 71.676
R512 B.n150 B.n149 71.676
R513 B.n145 B.n124 71.676
R514 B.n143 B.n142 71.676
R515 B.n138 B.n137 71.676
R516 B.n135 B.n134 71.676
R517 B.n130 B.n129 71.676
R518 B.n123 B.n122 59.5399
R519 B.n169 B.n116 59.5399
R520 B.n53 B.n52 59.5399
R521 B.n309 B.n59 59.5399
R522 B.n83 B.t1 55.0398
R523 B.t3 B.n378 55.0398
R524 B.n235 B.t1 51.8947
R525 B.n379 B.t3 51.8947
R526 B.n351 B.n350 32.9371
R527 B.n286 B.n285 32.9371
R528 B.n195 B.n105 32.9371
R529 B.n191 B.n190 32.9371
R530 B.n122 B.n121 30.255
R531 B.n116 B.n115 30.255
R532 B.n52 B.n51 30.255
R533 B.n59 B.n58 30.255
R534 B.n211 B.t5 29.879
R535 B.n363 B.t12 29.879
R536 B B.n397 18.0485
R537 B.n248 B.t0 11.0084
R538 B.n387 B.t2 11.0084
R539 B.n350 B.n349 10.6151
R540 B.n349 B.n45 10.6151
R541 B.n343 B.n45 10.6151
R542 B.n343 B.n342 10.6151
R543 B.n342 B.n341 10.6151
R544 B.n341 B.n47 10.6151
R545 B.n335 B.n47 10.6151
R546 B.n335 B.n334 10.6151
R547 B.n334 B.n333 10.6151
R548 B.n333 B.n49 10.6151
R549 B.n327 B.n326 10.6151
R550 B.n326 B.n325 10.6151
R551 B.n325 B.n54 10.6151
R552 B.n319 B.n54 10.6151
R553 B.n319 B.n318 10.6151
R554 B.n318 B.n317 10.6151
R555 B.n317 B.n56 10.6151
R556 B.n311 B.n56 10.6151
R557 B.n311 B.n310 10.6151
R558 B.n308 B.n60 10.6151
R559 B.n302 B.n60 10.6151
R560 B.n302 B.n301 10.6151
R561 B.n301 B.n300 10.6151
R562 B.n300 B.n62 10.6151
R563 B.n294 B.n62 10.6151
R564 B.n294 B.n293 10.6151
R565 B.n293 B.n292 10.6151
R566 B.n292 B.n64 10.6151
R567 B.n286 B.n64 10.6151
R568 B.n196 B.n195 10.6151
R569 B.n197 B.n196 10.6151
R570 B.n197 B.n96 10.6151
R571 B.n207 B.n96 10.6151
R572 B.n208 B.n207 10.6151
R573 B.n209 B.n208 10.6151
R574 B.n209 B.n89 10.6151
R575 B.n219 B.n89 10.6151
R576 B.n220 B.n219 10.6151
R577 B.n221 B.n220 10.6151
R578 B.n221 B.n80 10.6151
R579 B.n231 B.n80 10.6151
R580 B.n232 B.n231 10.6151
R581 B.n233 B.n232 10.6151
R582 B.n233 B.n73 10.6151
R583 B.n243 B.n73 10.6151
R584 B.n244 B.n243 10.6151
R585 B.n246 B.n244 10.6151
R586 B.n246 B.n245 10.6151
R587 B.n245 B.n65 10.6151
R588 B.n257 B.n65 10.6151
R589 B.n258 B.n257 10.6151
R590 B.n259 B.n258 10.6151
R591 B.n260 B.n259 10.6151
R592 B.n262 B.n260 10.6151
R593 B.n263 B.n262 10.6151
R594 B.n264 B.n263 10.6151
R595 B.n265 B.n264 10.6151
R596 B.n267 B.n265 10.6151
R597 B.n268 B.n267 10.6151
R598 B.n269 B.n268 10.6151
R599 B.n270 B.n269 10.6151
R600 B.n272 B.n270 10.6151
R601 B.n273 B.n272 10.6151
R602 B.n274 B.n273 10.6151
R603 B.n275 B.n274 10.6151
R604 B.n277 B.n275 10.6151
R605 B.n278 B.n277 10.6151
R606 B.n279 B.n278 10.6151
R607 B.n280 B.n279 10.6151
R608 B.n282 B.n280 10.6151
R609 B.n283 B.n282 10.6151
R610 B.n284 B.n283 10.6151
R611 B.n285 B.n284 10.6151
R612 B.n190 B.n189 10.6151
R613 B.n189 B.n109 10.6151
R614 B.n184 B.n109 10.6151
R615 B.n184 B.n183 10.6151
R616 B.n183 B.n111 10.6151
R617 B.n178 B.n111 10.6151
R618 B.n178 B.n177 10.6151
R619 B.n177 B.n176 10.6151
R620 B.n176 B.n113 10.6151
R621 B.n170 B.n113 10.6151
R622 B.n168 B.n167 10.6151
R623 B.n167 B.n117 10.6151
R624 B.n161 B.n117 10.6151
R625 B.n161 B.n160 10.6151
R626 B.n160 B.n159 10.6151
R627 B.n159 B.n119 10.6151
R628 B.n153 B.n119 10.6151
R629 B.n153 B.n152 10.6151
R630 B.n152 B.n151 10.6151
R631 B.n147 B.n146 10.6151
R632 B.n146 B.n125 10.6151
R633 B.n141 B.n125 10.6151
R634 B.n141 B.n140 10.6151
R635 B.n140 B.n139 10.6151
R636 B.n139 B.n127 10.6151
R637 B.n133 B.n127 10.6151
R638 B.n133 B.n132 10.6151
R639 B.n132 B.n131 10.6151
R640 B.n131 B.n105 10.6151
R641 B.n191 B.n101 10.6151
R642 B.n201 B.n101 10.6151
R643 B.n202 B.n201 10.6151
R644 B.n203 B.n202 10.6151
R645 B.n203 B.n93 10.6151
R646 B.n213 B.n93 10.6151
R647 B.n214 B.n213 10.6151
R648 B.n215 B.n214 10.6151
R649 B.n215 B.n85 10.6151
R650 B.n225 B.n85 10.6151
R651 B.n226 B.n225 10.6151
R652 B.n227 B.n226 10.6151
R653 B.n227 B.n77 10.6151
R654 B.n237 B.n77 10.6151
R655 B.n238 B.n237 10.6151
R656 B.n239 B.n238 10.6151
R657 B.n239 B.n69 10.6151
R658 B.n250 B.n69 10.6151
R659 B.n251 B.n250 10.6151
R660 B.n252 B.n251 10.6151
R661 B.n252 B.n0 10.6151
R662 B.n391 B.n1 10.6151
R663 B.n391 B.n390 10.6151
R664 B.n390 B.n389 10.6151
R665 B.n389 B.n10 10.6151
R666 B.n383 B.n10 10.6151
R667 B.n383 B.n382 10.6151
R668 B.n382 B.n381 10.6151
R669 B.n381 B.n17 10.6151
R670 B.n375 B.n17 10.6151
R671 B.n375 B.n374 10.6151
R672 B.n374 B.n373 10.6151
R673 B.n373 B.n24 10.6151
R674 B.n367 B.n24 10.6151
R675 B.n367 B.n366 10.6151
R676 B.n366 B.n365 10.6151
R677 B.n365 B.n31 10.6151
R678 B.n359 B.n31 10.6151
R679 B.n359 B.n358 10.6151
R680 B.n358 B.n357 10.6151
R681 B.n357 B.n38 10.6151
R682 B.n351 B.n38 10.6151
R683 B.n53 B.n49 9.36635
R684 B.n309 B.n308 9.36635
R685 B.n170 B.n169 9.36635
R686 B.n147 B.n123 9.36635
R687 B.n397 B.n0 2.81026
R688 B.n397 B.n1 2.81026
R689 B.n327 B.n53 1.24928
R690 B.n310 B.n309 1.24928
R691 B.n169 B.n168 1.24928
R692 B.n151 B.n123 1.24928
R693 VP.n4 VP.n3 172.012
R694 VP.n10 VP.n9 172.012
R695 VP.n8 VP.n0 161.3
R696 VP.n7 VP.n6 161.3
R697 VP.n5 VP.n1 161.3
R698 VP.n2 VP.t3 70.1085
R699 VP.n2 VP.t0 69.8876
R700 VP.n4 VP.n2 52.5757
R701 VP.n7 VP.n1 40.4106
R702 VP.n8 VP.n7 40.4106
R703 VP.n3 VP.t2 33.7013
R704 VP.n9 VP.t1 33.7013
R705 VP.n3 VP.n1 13.6328
R706 VP.n9 VP.n8 13.6328
R707 VP.n5 VP.n4 0.189894
R708 VP.n6 VP.n5 0.189894
R709 VP.n6 VP.n0 0.189894
R710 VP.n10 VP.n0 0.189894
R711 VP VP.n10 0.0516364
R712 VTAIL.n58 VTAIL.n56 289.615
R713 VTAIL.n2 VTAIL.n0 289.615
R714 VTAIL.n10 VTAIL.n8 289.615
R715 VTAIL.n18 VTAIL.n16 289.615
R716 VTAIL.n50 VTAIL.n48 289.615
R717 VTAIL.n42 VTAIL.n40 289.615
R718 VTAIL.n34 VTAIL.n32 289.615
R719 VTAIL.n26 VTAIL.n24 289.615
R720 VTAIL.n59 VTAIL.n58 185
R721 VTAIL.n3 VTAIL.n2 185
R722 VTAIL.n11 VTAIL.n10 185
R723 VTAIL.n19 VTAIL.n18 185
R724 VTAIL.n51 VTAIL.n50 185
R725 VTAIL.n43 VTAIL.n42 185
R726 VTAIL.n35 VTAIL.n34 185
R727 VTAIL.n27 VTAIL.n26 185
R728 VTAIL.t6 VTAIL.n57 164.876
R729 VTAIL.t7 VTAIL.n1 164.876
R730 VTAIL.t5 VTAIL.n9 164.876
R731 VTAIL.t4 VTAIL.n17 164.876
R732 VTAIL.t2 VTAIL.n49 164.876
R733 VTAIL.t3 VTAIL.n41 164.876
R734 VTAIL.t1 VTAIL.n33 164.876
R735 VTAIL.t0 VTAIL.n25 164.876
R736 VTAIL.n58 VTAIL.t6 52.3082
R737 VTAIL.n2 VTAIL.t7 52.3082
R738 VTAIL.n10 VTAIL.t5 52.3082
R739 VTAIL.n18 VTAIL.t4 52.3082
R740 VTAIL.n50 VTAIL.t2 52.3082
R741 VTAIL.n42 VTAIL.t3 52.3082
R742 VTAIL.n34 VTAIL.t1 52.3082
R743 VTAIL.n26 VTAIL.t0 52.3082
R744 VTAIL.n63 VTAIL.n62 32.9611
R745 VTAIL.n7 VTAIL.n6 32.9611
R746 VTAIL.n15 VTAIL.n14 32.9611
R747 VTAIL.n23 VTAIL.n22 32.9611
R748 VTAIL.n55 VTAIL.n54 32.9611
R749 VTAIL.n47 VTAIL.n46 32.9611
R750 VTAIL.n39 VTAIL.n38 32.9611
R751 VTAIL.n31 VTAIL.n30 32.9611
R752 VTAIL.n63 VTAIL.n55 15.1945
R753 VTAIL.n31 VTAIL.n23 15.1945
R754 VTAIL.n59 VTAIL.n57 14.7318
R755 VTAIL.n3 VTAIL.n1 14.7318
R756 VTAIL.n11 VTAIL.n9 14.7318
R757 VTAIL.n19 VTAIL.n17 14.7318
R758 VTAIL.n51 VTAIL.n49 14.7318
R759 VTAIL.n43 VTAIL.n41 14.7318
R760 VTAIL.n35 VTAIL.n33 14.7318
R761 VTAIL.n27 VTAIL.n25 14.7318
R762 VTAIL.n60 VTAIL.n56 12.8005
R763 VTAIL.n4 VTAIL.n0 12.8005
R764 VTAIL.n12 VTAIL.n8 12.8005
R765 VTAIL.n20 VTAIL.n16 12.8005
R766 VTAIL.n52 VTAIL.n48 12.8005
R767 VTAIL.n44 VTAIL.n40 12.8005
R768 VTAIL.n36 VTAIL.n32 12.8005
R769 VTAIL.n28 VTAIL.n24 12.8005
R770 VTAIL.n62 VTAIL.n61 9.45567
R771 VTAIL.n6 VTAIL.n5 9.45567
R772 VTAIL.n14 VTAIL.n13 9.45567
R773 VTAIL.n22 VTAIL.n21 9.45567
R774 VTAIL.n54 VTAIL.n53 9.45567
R775 VTAIL.n46 VTAIL.n45 9.45567
R776 VTAIL.n38 VTAIL.n37 9.45567
R777 VTAIL.n30 VTAIL.n29 9.45567
R778 VTAIL.n61 VTAIL.n60 9.3005
R779 VTAIL.n5 VTAIL.n4 9.3005
R780 VTAIL.n13 VTAIL.n12 9.3005
R781 VTAIL.n21 VTAIL.n20 9.3005
R782 VTAIL.n53 VTAIL.n52 9.3005
R783 VTAIL.n45 VTAIL.n44 9.3005
R784 VTAIL.n37 VTAIL.n36 9.3005
R785 VTAIL.n29 VTAIL.n28 9.3005
R786 VTAIL.n61 VTAIL.n57 5.62509
R787 VTAIL.n5 VTAIL.n1 5.62509
R788 VTAIL.n13 VTAIL.n9 5.62509
R789 VTAIL.n21 VTAIL.n17 5.62509
R790 VTAIL.n53 VTAIL.n49 5.62509
R791 VTAIL.n45 VTAIL.n41 5.62509
R792 VTAIL.n37 VTAIL.n33 5.62509
R793 VTAIL.n29 VTAIL.n25 5.62509
R794 VTAIL.n39 VTAIL.n31 1.34533
R795 VTAIL.n55 VTAIL.n47 1.34533
R796 VTAIL.n23 VTAIL.n15 1.34533
R797 VTAIL.n62 VTAIL.n56 1.16414
R798 VTAIL.n6 VTAIL.n0 1.16414
R799 VTAIL.n14 VTAIL.n8 1.16414
R800 VTAIL.n22 VTAIL.n16 1.16414
R801 VTAIL.n54 VTAIL.n48 1.16414
R802 VTAIL.n46 VTAIL.n40 1.16414
R803 VTAIL.n38 VTAIL.n32 1.16414
R804 VTAIL.n30 VTAIL.n24 1.16414
R805 VTAIL VTAIL.n7 0.731103
R806 VTAIL VTAIL.n63 0.614724
R807 VTAIL.n47 VTAIL.n39 0.470328
R808 VTAIL.n15 VTAIL.n7 0.470328
R809 VTAIL.n60 VTAIL.n59 0.388379
R810 VTAIL.n4 VTAIL.n3 0.388379
R811 VTAIL.n12 VTAIL.n11 0.388379
R812 VTAIL.n20 VTAIL.n19 0.388379
R813 VTAIL.n52 VTAIL.n51 0.388379
R814 VTAIL.n44 VTAIL.n43 0.388379
R815 VTAIL.n36 VTAIL.n35 0.388379
R816 VTAIL.n28 VTAIL.n27 0.388379
R817 VDD1 VDD1.n1 130.017
R818 VDD1 VDD1.n0 100.317
R819 VDD1.n0 VDD1.t0 11.5121
R820 VDD1.n0 VDD1.t3 11.5121
R821 VDD1.n1 VDD1.t1 11.5121
R822 VDD1.n1 VDD1.t2 11.5121
R823 VN.n0 VN.t0 70.1085
R824 VN.n1 VN.t1 70.1085
R825 VN.n0 VN.t3 69.8876
R826 VN.n1 VN.t2 69.8876
R827 VN VN.n1 52.9564
R828 VN VN.n0 18.3769
R829 VDD2.n2 VDD2.n0 129.492
R830 VDD2.n2 VDD2.n1 100.26
R831 VDD2.n1 VDD2.t1 11.5121
R832 VDD2.n1 VDD2.t2 11.5121
R833 VDD2.n0 VDD2.t3 11.5121
R834 VDD2.n0 VDD2.t0 11.5121
R835 VDD2 VDD2.n2 0.0586897
C0 VN VP 3.31223f
C1 VDD1 VN 0.153291f
C2 VTAIL VN 1.08278f
C3 VDD1 VP 0.98767f
C4 VDD2 VN 0.828735f
C5 VTAIL VP 1.09689f
C6 VDD1 VTAIL 2.33373f
C7 VDD2 VP 0.313487f
C8 VDD1 VDD2 0.691975f
C9 VTAIL VDD2 2.37875f
C10 VDD2 B 2.154549f
C11 VDD1 B 3.97683f
C12 VTAIL B 2.951793f
C13 VN B 6.60092f
C14 VP B 5.142353f
C15 VDD2.t3 B 0.027816f
C16 VDD2.t0 B 0.027816f
C17 VDD2.n0 B 0.331127f
C18 VDD2.t1 B 0.027816f
C19 VDD2.t2 B 0.027816f
C20 VDD2.n1 B 0.177599f
C21 VDD2.n2 B 1.68692f
C22 VN.t0 B 0.230756f
C23 VN.t3 B 0.230187f
C24 VN.n0 B 0.202597f
C25 VN.t1 B 0.230756f
C26 VN.t2 B 0.230187f
C27 VN.n1 B 0.836966f
C28 VDD1.t0 B 0.025843f
C29 VDD1.t3 B 0.025843f
C30 VDD1.n0 B 0.165132f
C31 VDD1.t1 B 0.025843f
C32 VDD1.t2 B 0.025843f
C33 VDD1.n1 B 0.31857f
C34 VTAIL.n0 B 0.021788f
C35 VTAIL.n1 B 0.051034f
C36 VTAIL.t7 B 0.036937f
C37 VTAIL.n2 B 0.03761f
C38 VTAIL.n3 B 0.011351f
C39 VTAIL.n4 B 0.009214f
C40 VTAIL.n5 B 0.098838f
C41 VTAIL.n6 B 0.023699f
C42 VTAIL.n7 B 0.081498f
C43 VTAIL.n8 B 0.021788f
C44 VTAIL.n9 B 0.051034f
C45 VTAIL.t5 B 0.036937f
C46 VTAIL.n10 B 0.03761f
C47 VTAIL.n11 B 0.011351f
C48 VTAIL.n12 B 0.009214f
C49 VTAIL.n13 B 0.098838f
C50 VTAIL.n14 B 0.023699f
C51 VTAIL.n15 B 0.115435f
C52 VTAIL.n16 B 0.021788f
C53 VTAIL.n17 B 0.051034f
C54 VTAIL.t4 B 0.036937f
C55 VTAIL.n18 B 0.03761f
C56 VTAIL.n19 B 0.011351f
C57 VTAIL.n20 B 0.009214f
C58 VTAIL.n21 B 0.098838f
C59 VTAIL.n22 B 0.023699f
C60 VTAIL.n23 B 0.478622f
C61 VTAIL.n24 B 0.021788f
C62 VTAIL.n25 B 0.051034f
C63 VTAIL.t0 B 0.036937f
C64 VTAIL.n26 B 0.03761f
C65 VTAIL.n27 B 0.011351f
C66 VTAIL.n28 B 0.009214f
C67 VTAIL.n29 B 0.098838f
C68 VTAIL.n30 B 0.023699f
C69 VTAIL.n31 B 0.478622f
C70 VTAIL.n32 B 0.021788f
C71 VTAIL.n33 B 0.051034f
C72 VTAIL.t1 B 0.036937f
C73 VTAIL.n34 B 0.03761f
C74 VTAIL.n35 B 0.011351f
C75 VTAIL.n36 B 0.009214f
C76 VTAIL.n37 B 0.098838f
C77 VTAIL.n38 B 0.023699f
C78 VTAIL.n39 B 0.115435f
C79 VTAIL.n40 B 0.021788f
C80 VTAIL.n41 B 0.051034f
C81 VTAIL.t3 B 0.036937f
C82 VTAIL.n42 B 0.03761f
C83 VTAIL.n43 B 0.011351f
C84 VTAIL.n44 B 0.009214f
C85 VTAIL.n45 B 0.098838f
C86 VTAIL.n46 B 0.023699f
C87 VTAIL.n47 B 0.115435f
C88 VTAIL.n48 B 0.021788f
C89 VTAIL.n49 B 0.051034f
C90 VTAIL.t2 B 0.036937f
C91 VTAIL.n50 B 0.03761f
C92 VTAIL.n51 B 0.011351f
C93 VTAIL.n52 B 0.009214f
C94 VTAIL.n53 B 0.098838f
C95 VTAIL.n54 B 0.023699f
C96 VTAIL.n55 B 0.478622f
C97 VTAIL.n56 B 0.021788f
C98 VTAIL.n57 B 0.051034f
C99 VTAIL.t6 B 0.036937f
C100 VTAIL.n58 B 0.03761f
C101 VTAIL.n59 B 0.011351f
C102 VTAIL.n60 B 0.009214f
C103 VTAIL.n61 B 0.098838f
C104 VTAIL.n62 B 0.023699f
C105 VTAIL.n63 B 0.438256f
C106 VP.n0 B 0.029252f
C107 VP.t1 B 0.13982f
C108 VP.n1 B 0.046545f
C109 VP.t3 B 0.233631f
C110 VP.t0 B 0.233055f
C111 VP.n2 B 0.832246f
C112 VP.t2 B 0.13982f
C113 VP.n3 B 0.13675f
C114 VP.n4 B 1.20548f
C115 VP.n5 B 0.029252f
C116 VP.n6 B 0.029252f
C117 VP.n7 B 0.023671f
C118 VP.n8 B 0.046545f
C119 VP.n9 B 0.13675f
C120 VP.n10 B 0.026115f
.ends

