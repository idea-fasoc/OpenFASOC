* NGSPICE file created from diff_pair_sample_0736.ext - technology: sky130A

.subckt diff_pair_sample_0736 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VN.t0 VDD2.t3 w_n5050_n4556# sky130_fd_pr__pfet_01v8 ad=6.9966 pd=36.66 as=2.9601 ps=18.27 w=17.94 l=3.75
X1 VDD2.t2 VN.t1 VTAIL.t14 w_n5050_n4556# sky130_fd_pr__pfet_01v8 ad=2.9601 pd=18.27 as=2.9601 ps=18.27 w=17.94 l=3.75
X2 VDD2.t5 VN.t2 VTAIL.t13 w_n5050_n4556# sky130_fd_pr__pfet_01v8 ad=2.9601 pd=18.27 as=6.9966 ps=36.66 w=17.94 l=3.75
X3 B.t11 B.t9 B.t10 w_n5050_n4556# sky130_fd_pr__pfet_01v8 ad=6.9966 pd=36.66 as=0 ps=0 w=17.94 l=3.75
X4 B.t8 B.t6 B.t7 w_n5050_n4556# sky130_fd_pr__pfet_01v8 ad=6.9966 pd=36.66 as=0 ps=0 w=17.94 l=3.75
X5 VTAIL.t12 VN.t3 VDD2.t4 w_n5050_n4556# sky130_fd_pr__pfet_01v8 ad=6.9966 pd=36.66 as=2.9601 ps=18.27 w=17.94 l=3.75
X6 B.t5 B.t3 B.t4 w_n5050_n4556# sky130_fd_pr__pfet_01v8 ad=6.9966 pd=36.66 as=0 ps=0 w=17.94 l=3.75
X7 VTAIL.t11 VN.t4 VDD2.t1 w_n5050_n4556# sky130_fd_pr__pfet_01v8 ad=2.9601 pd=18.27 as=2.9601 ps=18.27 w=17.94 l=3.75
X8 VDD1.t7 VP.t0 VTAIL.t5 w_n5050_n4556# sky130_fd_pr__pfet_01v8 ad=2.9601 pd=18.27 as=2.9601 ps=18.27 w=17.94 l=3.75
X9 VTAIL.t7 VP.t1 VDD1.t6 w_n5050_n4556# sky130_fd_pr__pfet_01v8 ad=6.9966 pd=36.66 as=2.9601 ps=18.27 w=17.94 l=3.75
X10 VDD2.t0 VN.t5 VTAIL.t10 w_n5050_n4556# sky130_fd_pr__pfet_01v8 ad=2.9601 pd=18.27 as=6.9966 ps=36.66 w=17.94 l=3.75
X11 VDD2.t7 VN.t6 VTAIL.t9 w_n5050_n4556# sky130_fd_pr__pfet_01v8 ad=2.9601 pd=18.27 as=2.9601 ps=18.27 w=17.94 l=3.75
X12 VDD1.t5 VP.t2 VTAIL.t6 w_n5050_n4556# sky130_fd_pr__pfet_01v8 ad=2.9601 pd=18.27 as=6.9966 ps=36.66 w=17.94 l=3.75
X13 VTAIL.t3 VP.t3 VDD1.t4 w_n5050_n4556# sky130_fd_pr__pfet_01v8 ad=2.9601 pd=18.27 as=2.9601 ps=18.27 w=17.94 l=3.75
X14 VDD1.t3 VP.t4 VTAIL.t4 w_n5050_n4556# sky130_fd_pr__pfet_01v8 ad=2.9601 pd=18.27 as=2.9601 ps=18.27 w=17.94 l=3.75
X15 VDD1.t2 VP.t5 VTAIL.t2 w_n5050_n4556# sky130_fd_pr__pfet_01v8 ad=2.9601 pd=18.27 as=6.9966 ps=36.66 w=17.94 l=3.75
X16 VTAIL.t8 VN.t7 VDD2.t6 w_n5050_n4556# sky130_fd_pr__pfet_01v8 ad=2.9601 pd=18.27 as=2.9601 ps=18.27 w=17.94 l=3.75
X17 VTAIL.t1 VP.t6 VDD1.t1 w_n5050_n4556# sky130_fd_pr__pfet_01v8 ad=2.9601 pd=18.27 as=2.9601 ps=18.27 w=17.94 l=3.75
X18 B.t2 B.t0 B.t1 w_n5050_n4556# sky130_fd_pr__pfet_01v8 ad=6.9966 pd=36.66 as=0 ps=0 w=17.94 l=3.75
X19 VTAIL.t0 VP.t7 VDD1.t0 w_n5050_n4556# sky130_fd_pr__pfet_01v8 ad=6.9966 pd=36.66 as=2.9601 ps=18.27 w=17.94 l=3.75
R0 VN.n76 VN.n75 161.3
R1 VN.n74 VN.n40 161.3
R2 VN.n73 VN.n72 161.3
R3 VN.n71 VN.n41 161.3
R4 VN.n70 VN.n69 161.3
R5 VN.n68 VN.n42 161.3
R6 VN.n67 VN.n66 161.3
R7 VN.n65 VN.n43 161.3
R8 VN.n64 VN.n63 161.3
R9 VN.n62 VN.n44 161.3
R10 VN.n61 VN.n60 161.3
R11 VN.n59 VN.n46 161.3
R12 VN.n58 VN.n57 161.3
R13 VN.n56 VN.n47 161.3
R14 VN.n55 VN.n54 161.3
R15 VN.n53 VN.n48 161.3
R16 VN.n52 VN.n51 161.3
R17 VN.n37 VN.n36 161.3
R18 VN.n35 VN.n1 161.3
R19 VN.n34 VN.n33 161.3
R20 VN.n32 VN.n2 161.3
R21 VN.n31 VN.n30 161.3
R22 VN.n29 VN.n3 161.3
R23 VN.n28 VN.n27 161.3
R24 VN.n26 VN.n4 161.3
R25 VN.n25 VN.n24 161.3
R26 VN.n22 VN.n5 161.3
R27 VN.n21 VN.n20 161.3
R28 VN.n19 VN.n6 161.3
R29 VN.n18 VN.n17 161.3
R30 VN.n16 VN.n7 161.3
R31 VN.n15 VN.n14 161.3
R32 VN.n13 VN.n8 161.3
R33 VN.n12 VN.n11 161.3
R34 VN.n49 VN.t2 147.802
R35 VN.n9 VN.t0 147.802
R36 VN.n10 VN.t6 115.294
R37 VN.n23 VN.t4 115.294
R38 VN.n0 VN.t5 115.294
R39 VN.n50 VN.t7 115.294
R40 VN.n45 VN.t1 115.294
R41 VN.n39 VN.t3 115.294
R42 VN.n38 VN.n0 84.0486
R43 VN.n77 VN.n39 84.0486
R44 VN.n10 VN.n9 72.7154
R45 VN.n50 VN.n49 72.7153
R46 VN VN.n77 61.0282
R47 VN.n30 VN.n2 48.2005
R48 VN.n69 VN.n41 48.2005
R49 VN.n17 VN.n16 40.4106
R50 VN.n17 VN.n6 40.4106
R51 VN.n57 VN.n56 40.4106
R52 VN.n57 VN.n46 40.4106
R53 VN.n30 VN.n29 32.6207
R54 VN.n69 VN.n68 32.6207
R55 VN.n11 VN.n8 24.3439
R56 VN.n15 VN.n8 24.3439
R57 VN.n16 VN.n15 24.3439
R58 VN.n21 VN.n6 24.3439
R59 VN.n22 VN.n21 24.3439
R60 VN.n24 VN.n22 24.3439
R61 VN.n28 VN.n4 24.3439
R62 VN.n29 VN.n28 24.3439
R63 VN.n34 VN.n2 24.3439
R64 VN.n35 VN.n34 24.3439
R65 VN.n36 VN.n35 24.3439
R66 VN.n56 VN.n55 24.3439
R67 VN.n55 VN.n48 24.3439
R68 VN.n51 VN.n48 24.3439
R69 VN.n68 VN.n67 24.3439
R70 VN.n67 VN.n43 24.3439
R71 VN.n63 VN.n62 24.3439
R72 VN.n62 VN.n61 24.3439
R73 VN.n61 VN.n46 24.3439
R74 VN.n75 VN.n74 24.3439
R75 VN.n74 VN.n73 24.3439
R76 VN.n73 VN.n41 24.3439
R77 VN.n23 VN.n4 22.3965
R78 VN.n45 VN.n43 22.3965
R79 VN.n36 VN.n0 5.84292
R80 VN.n75 VN.n39 5.84292
R81 VN.n12 VN.n9 3.29535
R82 VN.n52 VN.n49 3.29535
R83 VN.n11 VN.n10 1.94797
R84 VN.n24 VN.n23 1.94797
R85 VN.n51 VN.n50 1.94797
R86 VN.n63 VN.n45 1.94797
R87 VN.n77 VN.n76 0.355081
R88 VN.n38 VN.n37 0.355081
R89 VN VN.n38 0.26685
R90 VN.n76 VN.n40 0.189894
R91 VN.n72 VN.n40 0.189894
R92 VN.n72 VN.n71 0.189894
R93 VN.n71 VN.n70 0.189894
R94 VN.n70 VN.n42 0.189894
R95 VN.n66 VN.n42 0.189894
R96 VN.n66 VN.n65 0.189894
R97 VN.n65 VN.n64 0.189894
R98 VN.n64 VN.n44 0.189894
R99 VN.n60 VN.n44 0.189894
R100 VN.n60 VN.n59 0.189894
R101 VN.n59 VN.n58 0.189894
R102 VN.n58 VN.n47 0.189894
R103 VN.n54 VN.n47 0.189894
R104 VN.n54 VN.n53 0.189894
R105 VN.n53 VN.n52 0.189894
R106 VN.n13 VN.n12 0.189894
R107 VN.n14 VN.n13 0.189894
R108 VN.n14 VN.n7 0.189894
R109 VN.n18 VN.n7 0.189894
R110 VN.n19 VN.n18 0.189894
R111 VN.n20 VN.n19 0.189894
R112 VN.n20 VN.n5 0.189894
R113 VN.n25 VN.n5 0.189894
R114 VN.n26 VN.n25 0.189894
R115 VN.n27 VN.n26 0.189894
R116 VN.n27 VN.n3 0.189894
R117 VN.n31 VN.n3 0.189894
R118 VN.n32 VN.n31 0.189894
R119 VN.n33 VN.n32 0.189894
R120 VN.n33 VN.n1 0.189894
R121 VN.n37 VN.n1 0.189894
R122 VDD2.n2 VDD2.n1 71.7174
R123 VDD2.n2 VDD2.n0 71.7174
R124 VDD2 VDD2.n5 71.7146
R125 VDD2.n4 VDD2.n3 70.0143
R126 VDD2.n4 VDD2.n2 55.0084
R127 VDD2 VDD2.n4 1.81731
R128 VDD2.n5 VDD2.t6 1.81237
R129 VDD2.n5 VDD2.t5 1.81237
R130 VDD2.n3 VDD2.t4 1.81237
R131 VDD2.n3 VDD2.t2 1.81237
R132 VDD2.n1 VDD2.t1 1.81237
R133 VDD2.n1 VDD2.t0 1.81237
R134 VDD2.n0 VDD2.t3 1.81237
R135 VDD2.n0 VDD2.t7 1.81237
R136 VTAIL.n11 VTAIL.t0 55.1474
R137 VTAIL.n10 VTAIL.t13 55.1474
R138 VTAIL.n7 VTAIL.t12 55.1474
R139 VTAIL.n15 VTAIL.t10 55.1472
R140 VTAIL.n2 VTAIL.t15 55.1472
R141 VTAIL.n3 VTAIL.t6 55.1472
R142 VTAIL.n6 VTAIL.t7 55.1472
R143 VTAIL.n14 VTAIL.t2 55.1472
R144 VTAIL.n13 VTAIL.n12 53.3355
R145 VTAIL.n9 VTAIL.n8 53.3355
R146 VTAIL.n1 VTAIL.n0 53.3353
R147 VTAIL.n5 VTAIL.n4 53.3353
R148 VTAIL.n15 VTAIL.n14 31.3496
R149 VTAIL.n7 VTAIL.n6 31.3496
R150 VTAIL.n9 VTAIL.n7 3.51774
R151 VTAIL.n10 VTAIL.n9 3.51774
R152 VTAIL.n13 VTAIL.n11 3.51774
R153 VTAIL.n14 VTAIL.n13 3.51774
R154 VTAIL.n6 VTAIL.n5 3.51774
R155 VTAIL.n5 VTAIL.n3 3.51774
R156 VTAIL.n2 VTAIL.n1 3.51774
R157 VTAIL VTAIL.n15 3.45955
R158 VTAIL.n0 VTAIL.t9 1.81237
R159 VTAIL.n0 VTAIL.t11 1.81237
R160 VTAIL.n4 VTAIL.t4 1.81237
R161 VTAIL.n4 VTAIL.t1 1.81237
R162 VTAIL.n12 VTAIL.t5 1.81237
R163 VTAIL.n12 VTAIL.t3 1.81237
R164 VTAIL.n8 VTAIL.t14 1.81237
R165 VTAIL.n8 VTAIL.t8 1.81237
R166 VTAIL.n11 VTAIL.n10 0.470328
R167 VTAIL.n3 VTAIL.n2 0.470328
R168 VTAIL VTAIL.n1 0.0586897
R169 B.n776 B.n775 585
R170 B.n777 B.n104 585
R171 B.n779 B.n778 585
R172 B.n780 B.n103 585
R173 B.n782 B.n781 585
R174 B.n783 B.n102 585
R175 B.n785 B.n784 585
R176 B.n786 B.n101 585
R177 B.n788 B.n787 585
R178 B.n789 B.n100 585
R179 B.n791 B.n790 585
R180 B.n792 B.n99 585
R181 B.n794 B.n793 585
R182 B.n795 B.n98 585
R183 B.n797 B.n796 585
R184 B.n798 B.n97 585
R185 B.n800 B.n799 585
R186 B.n801 B.n96 585
R187 B.n803 B.n802 585
R188 B.n804 B.n95 585
R189 B.n806 B.n805 585
R190 B.n807 B.n94 585
R191 B.n809 B.n808 585
R192 B.n810 B.n93 585
R193 B.n812 B.n811 585
R194 B.n813 B.n92 585
R195 B.n815 B.n814 585
R196 B.n816 B.n91 585
R197 B.n818 B.n817 585
R198 B.n819 B.n90 585
R199 B.n821 B.n820 585
R200 B.n822 B.n89 585
R201 B.n824 B.n823 585
R202 B.n825 B.n88 585
R203 B.n827 B.n826 585
R204 B.n828 B.n87 585
R205 B.n830 B.n829 585
R206 B.n831 B.n86 585
R207 B.n833 B.n832 585
R208 B.n834 B.n85 585
R209 B.n836 B.n835 585
R210 B.n837 B.n84 585
R211 B.n839 B.n838 585
R212 B.n840 B.n83 585
R213 B.n842 B.n841 585
R214 B.n843 B.n82 585
R215 B.n845 B.n844 585
R216 B.n846 B.n81 585
R217 B.n848 B.n847 585
R218 B.n849 B.n80 585
R219 B.n851 B.n850 585
R220 B.n852 B.n79 585
R221 B.n854 B.n853 585
R222 B.n855 B.n78 585
R223 B.n857 B.n856 585
R224 B.n858 B.n77 585
R225 B.n860 B.n859 585
R226 B.n861 B.n73 585
R227 B.n863 B.n862 585
R228 B.n864 B.n72 585
R229 B.n866 B.n865 585
R230 B.n867 B.n71 585
R231 B.n869 B.n868 585
R232 B.n870 B.n70 585
R233 B.n872 B.n871 585
R234 B.n873 B.n69 585
R235 B.n875 B.n874 585
R236 B.n876 B.n68 585
R237 B.n878 B.n877 585
R238 B.n880 B.n65 585
R239 B.n882 B.n881 585
R240 B.n883 B.n64 585
R241 B.n885 B.n884 585
R242 B.n886 B.n63 585
R243 B.n888 B.n887 585
R244 B.n889 B.n62 585
R245 B.n891 B.n890 585
R246 B.n892 B.n61 585
R247 B.n894 B.n893 585
R248 B.n895 B.n60 585
R249 B.n897 B.n896 585
R250 B.n898 B.n59 585
R251 B.n900 B.n899 585
R252 B.n901 B.n58 585
R253 B.n903 B.n902 585
R254 B.n904 B.n57 585
R255 B.n906 B.n905 585
R256 B.n907 B.n56 585
R257 B.n909 B.n908 585
R258 B.n910 B.n55 585
R259 B.n912 B.n911 585
R260 B.n913 B.n54 585
R261 B.n915 B.n914 585
R262 B.n916 B.n53 585
R263 B.n918 B.n917 585
R264 B.n919 B.n52 585
R265 B.n921 B.n920 585
R266 B.n922 B.n51 585
R267 B.n924 B.n923 585
R268 B.n925 B.n50 585
R269 B.n927 B.n926 585
R270 B.n928 B.n49 585
R271 B.n930 B.n929 585
R272 B.n931 B.n48 585
R273 B.n933 B.n932 585
R274 B.n934 B.n47 585
R275 B.n936 B.n935 585
R276 B.n937 B.n46 585
R277 B.n939 B.n938 585
R278 B.n940 B.n45 585
R279 B.n942 B.n941 585
R280 B.n943 B.n44 585
R281 B.n945 B.n944 585
R282 B.n946 B.n43 585
R283 B.n948 B.n947 585
R284 B.n949 B.n42 585
R285 B.n951 B.n950 585
R286 B.n952 B.n41 585
R287 B.n954 B.n953 585
R288 B.n955 B.n40 585
R289 B.n957 B.n956 585
R290 B.n958 B.n39 585
R291 B.n960 B.n959 585
R292 B.n961 B.n38 585
R293 B.n963 B.n962 585
R294 B.n964 B.n37 585
R295 B.n966 B.n965 585
R296 B.n967 B.n36 585
R297 B.n774 B.n105 585
R298 B.n773 B.n772 585
R299 B.n771 B.n106 585
R300 B.n770 B.n769 585
R301 B.n768 B.n107 585
R302 B.n767 B.n766 585
R303 B.n765 B.n108 585
R304 B.n764 B.n763 585
R305 B.n762 B.n109 585
R306 B.n761 B.n760 585
R307 B.n759 B.n110 585
R308 B.n758 B.n757 585
R309 B.n756 B.n111 585
R310 B.n755 B.n754 585
R311 B.n753 B.n112 585
R312 B.n752 B.n751 585
R313 B.n750 B.n113 585
R314 B.n749 B.n748 585
R315 B.n747 B.n114 585
R316 B.n746 B.n745 585
R317 B.n744 B.n115 585
R318 B.n743 B.n742 585
R319 B.n741 B.n116 585
R320 B.n740 B.n739 585
R321 B.n738 B.n117 585
R322 B.n737 B.n736 585
R323 B.n735 B.n118 585
R324 B.n734 B.n733 585
R325 B.n732 B.n119 585
R326 B.n731 B.n730 585
R327 B.n729 B.n120 585
R328 B.n728 B.n727 585
R329 B.n726 B.n121 585
R330 B.n725 B.n724 585
R331 B.n723 B.n122 585
R332 B.n722 B.n721 585
R333 B.n720 B.n123 585
R334 B.n719 B.n718 585
R335 B.n717 B.n124 585
R336 B.n716 B.n715 585
R337 B.n714 B.n125 585
R338 B.n713 B.n712 585
R339 B.n711 B.n126 585
R340 B.n710 B.n709 585
R341 B.n708 B.n127 585
R342 B.n707 B.n706 585
R343 B.n705 B.n128 585
R344 B.n704 B.n703 585
R345 B.n702 B.n129 585
R346 B.n701 B.n700 585
R347 B.n699 B.n130 585
R348 B.n698 B.n697 585
R349 B.n696 B.n131 585
R350 B.n695 B.n694 585
R351 B.n693 B.n132 585
R352 B.n692 B.n691 585
R353 B.n690 B.n133 585
R354 B.n689 B.n688 585
R355 B.n687 B.n134 585
R356 B.n686 B.n685 585
R357 B.n684 B.n135 585
R358 B.n683 B.n682 585
R359 B.n681 B.n136 585
R360 B.n680 B.n679 585
R361 B.n678 B.n137 585
R362 B.n677 B.n676 585
R363 B.n675 B.n138 585
R364 B.n674 B.n673 585
R365 B.n672 B.n139 585
R366 B.n671 B.n670 585
R367 B.n669 B.n140 585
R368 B.n668 B.n667 585
R369 B.n666 B.n141 585
R370 B.n665 B.n664 585
R371 B.n663 B.n142 585
R372 B.n662 B.n661 585
R373 B.n660 B.n143 585
R374 B.n659 B.n658 585
R375 B.n657 B.n144 585
R376 B.n656 B.n655 585
R377 B.n654 B.n145 585
R378 B.n653 B.n652 585
R379 B.n651 B.n146 585
R380 B.n650 B.n649 585
R381 B.n648 B.n147 585
R382 B.n647 B.n646 585
R383 B.n645 B.n148 585
R384 B.n644 B.n643 585
R385 B.n642 B.n149 585
R386 B.n641 B.n640 585
R387 B.n639 B.n150 585
R388 B.n638 B.n637 585
R389 B.n636 B.n151 585
R390 B.n635 B.n634 585
R391 B.n633 B.n152 585
R392 B.n632 B.n631 585
R393 B.n630 B.n153 585
R394 B.n629 B.n628 585
R395 B.n627 B.n154 585
R396 B.n626 B.n625 585
R397 B.n624 B.n155 585
R398 B.n623 B.n622 585
R399 B.n621 B.n156 585
R400 B.n620 B.n619 585
R401 B.n618 B.n157 585
R402 B.n617 B.n616 585
R403 B.n615 B.n158 585
R404 B.n614 B.n613 585
R405 B.n612 B.n159 585
R406 B.n611 B.n610 585
R407 B.n609 B.n160 585
R408 B.n608 B.n607 585
R409 B.n606 B.n161 585
R410 B.n605 B.n604 585
R411 B.n603 B.n162 585
R412 B.n602 B.n601 585
R413 B.n600 B.n163 585
R414 B.n599 B.n598 585
R415 B.n597 B.n164 585
R416 B.n596 B.n595 585
R417 B.n594 B.n165 585
R418 B.n593 B.n592 585
R419 B.n591 B.n166 585
R420 B.n590 B.n589 585
R421 B.n588 B.n167 585
R422 B.n587 B.n586 585
R423 B.n585 B.n168 585
R424 B.n584 B.n583 585
R425 B.n582 B.n169 585
R426 B.n581 B.n580 585
R427 B.n579 B.n170 585
R428 B.n578 B.n577 585
R429 B.n576 B.n171 585
R430 B.n575 B.n574 585
R431 B.n573 B.n172 585
R432 B.n572 B.n571 585
R433 B.n570 B.n173 585
R434 B.n377 B.n376 585
R435 B.n378 B.n241 585
R436 B.n380 B.n379 585
R437 B.n381 B.n240 585
R438 B.n383 B.n382 585
R439 B.n384 B.n239 585
R440 B.n386 B.n385 585
R441 B.n387 B.n238 585
R442 B.n389 B.n388 585
R443 B.n390 B.n237 585
R444 B.n392 B.n391 585
R445 B.n393 B.n236 585
R446 B.n395 B.n394 585
R447 B.n396 B.n235 585
R448 B.n398 B.n397 585
R449 B.n399 B.n234 585
R450 B.n401 B.n400 585
R451 B.n402 B.n233 585
R452 B.n404 B.n403 585
R453 B.n405 B.n232 585
R454 B.n407 B.n406 585
R455 B.n408 B.n231 585
R456 B.n410 B.n409 585
R457 B.n411 B.n230 585
R458 B.n413 B.n412 585
R459 B.n414 B.n229 585
R460 B.n416 B.n415 585
R461 B.n417 B.n228 585
R462 B.n419 B.n418 585
R463 B.n420 B.n227 585
R464 B.n422 B.n421 585
R465 B.n423 B.n226 585
R466 B.n425 B.n424 585
R467 B.n426 B.n225 585
R468 B.n428 B.n427 585
R469 B.n429 B.n224 585
R470 B.n431 B.n430 585
R471 B.n432 B.n223 585
R472 B.n434 B.n433 585
R473 B.n435 B.n222 585
R474 B.n437 B.n436 585
R475 B.n438 B.n221 585
R476 B.n440 B.n439 585
R477 B.n441 B.n220 585
R478 B.n443 B.n442 585
R479 B.n444 B.n219 585
R480 B.n446 B.n445 585
R481 B.n447 B.n218 585
R482 B.n449 B.n448 585
R483 B.n450 B.n217 585
R484 B.n452 B.n451 585
R485 B.n453 B.n216 585
R486 B.n455 B.n454 585
R487 B.n456 B.n215 585
R488 B.n458 B.n457 585
R489 B.n459 B.n214 585
R490 B.n461 B.n460 585
R491 B.n462 B.n213 585
R492 B.n464 B.n463 585
R493 B.n466 B.n210 585
R494 B.n468 B.n467 585
R495 B.n469 B.n209 585
R496 B.n471 B.n470 585
R497 B.n472 B.n208 585
R498 B.n474 B.n473 585
R499 B.n475 B.n207 585
R500 B.n477 B.n476 585
R501 B.n478 B.n206 585
R502 B.n480 B.n479 585
R503 B.n482 B.n481 585
R504 B.n483 B.n202 585
R505 B.n485 B.n484 585
R506 B.n486 B.n201 585
R507 B.n488 B.n487 585
R508 B.n489 B.n200 585
R509 B.n491 B.n490 585
R510 B.n492 B.n199 585
R511 B.n494 B.n493 585
R512 B.n495 B.n198 585
R513 B.n497 B.n496 585
R514 B.n498 B.n197 585
R515 B.n500 B.n499 585
R516 B.n501 B.n196 585
R517 B.n503 B.n502 585
R518 B.n504 B.n195 585
R519 B.n506 B.n505 585
R520 B.n507 B.n194 585
R521 B.n509 B.n508 585
R522 B.n510 B.n193 585
R523 B.n512 B.n511 585
R524 B.n513 B.n192 585
R525 B.n515 B.n514 585
R526 B.n516 B.n191 585
R527 B.n518 B.n517 585
R528 B.n519 B.n190 585
R529 B.n521 B.n520 585
R530 B.n522 B.n189 585
R531 B.n524 B.n523 585
R532 B.n525 B.n188 585
R533 B.n527 B.n526 585
R534 B.n528 B.n187 585
R535 B.n530 B.n529 585
R536 B.n531 B.n186 585
R537 B.n533 B.n532 585
R538 B.n534 B.n185 585
R539 B.n536 B.n535 585
R540 B.n537 B.n184 585
R541 B.n539 B.n538 585
R542 B.n540 B.n183 585
R543 B.n542 B.n541 585
R544 B.n543 B.n182 585
R545 B.n545 B.n544 585
R546 B.n546 B.n181 585
R547 B.n548 B.n547 585
R548 B.n549 B.n180 585
R549 B.n551 B.n550 585
R550 B.n552 B.n179 585
R551 B.n554 B.n553 585
R552 B.n555 B.n178 585
R553 B.n557 B.n556 585
R554 B.n558 B.n177 585
R555 B.n560 B.n559 585
R556 B.n561 B.n176 585
R557 B.n563 B.n562 585
R558 B.n564 B.n175 585
R559 B.n566 B.n565 585
R560 B.n567 B.n174 585
R561 B.n569 B.n568 585
R562 B.n375 B.n242 585
R563 B.n374 B.n373 585
R564 B.n372 B.n243 585
R565 B.n371 B.n370 585
R566 B.n369 B.n244 585
R567 B.n368 B.n367 585
R568 B.n366 B.n245 585
R569 B.n365 B.n364 585
R570 B.n363 B.n246 585
R571 B.n362 B.n361 585
R572 B.n360 B.n247 585
R573 B.n359 B.n358 585
R574 B.n357 B.n248 585
R575 B.n356 B.n355 585
R576 B.n354 B.n249 585
R577 B.n353 B.n352 585
R578 B.n351 B.n250 585
R579 B.n350 B.n349 585
R580 B.n348 B.n251 585
R581 B.n347 B.n346 585
R582 B.n345 B.n252 585
R583 B.n344 B.n343 585
R584 B.n342 B.n253 585
R585 B.n341 B.n340 585
R586 B.n339 B.n254 585
R587 B.n338 B.n337 585
R588 B.n336 B.n255 585
R589 B.n335 B.n334 585
R590 B.n333 B.n256 585
R591 B.n332 B.n331 585
R592 B.n330 B.n257 585
R593 B.n329 B.n328 585
R594 B.n327 B.n258 585
R595 B.n326 B.n325 585
R596 B.n324 B.n259 585
R597 B.n323 B.n322 585
R598 B.n321 B.n260 585
R599 B.n320 B.n319 585
R600 B.n318 B.n261 585
R601 B.n317 B.n316 585
R602 B.n315 B.n262 585
R603 B.n314 B.n313 585
R604 B.n312 B.n263 585
R605 B.n311 B.n310 585
R606 B.n309 B.n264 585
R607 B.n308 B.n307 585
R608 B.n306 B.n265 585
R609 B.n305 B.n304 585
R610 B.n303 B.n266 585
R611 B.n302 B.n301 585
R612 B.n300 B.n267 585
R613 B.n299 B.n298 585
R614 B.n297 B.n268 585
R615 B.n296 B.n295 585
R616 B.n294 B.n269 585
R617 B.n293 B.n292 585
R618 B.n291 B.n270 585
R619 B.n290 B.n289 585
R620 B.n288 B.n271 585
R621 B.n287 B.n286 585
R622 B.n285 B.n272 585
R623 B.n284 B.n283 585
R624 B.n282 B.n273 585
R625 B.n281 B.n280 585
R626 B.n279 B.n274 585
R627 B.n278 B.n277 585
R628 B.n276 B.n275 585
R629 B.n2 B.n0 585
R630 B.n1069 B.n1 585
R631 B.n1068 B.n1067 585
R632 B.n1066 B.n3 585
R633 B.n1065 B.n1064 585
R634 B.n1063 B.n4 585
R635 B.n1062 B.n1061 585
R636 B.n1060 B.n5 585
R637 B.n1059 B.n1058 585
R638 B.n1057 B.n6 585
R639 B.n1056 B.n1055 585
R640 B.n1054 B.n7 585
R641 B.n1053 B.n1052 585
R642 B.n1051 B.n8 585
R643 B.n1050 B.n1049 585
R644 B.n1048 B.n9 585
R645 B.n1047 B.n1046 585
R646 B.n1045 B.n10 585
R647 B.n1044 B.n1043 585
R648 B.n1042 B.n11 585
R649 B.n1041 B.n1040 585
R650 B.n1039 B.n12 585
R651 B.n1038 B.n1037 585
R652 B.n1036 B.n13 585
R653 B.n1035 B.n1034 585
R654 B.n1033 B.n14 585
R655 B.n1032 B.n1031 585
R656 B.n1030 B.n15 585
R657 B.n1029 B.n1028 585
R658 B.n1027 B.n16 585
R659 B.n1026 B.n1025 585
R660 B.n1024 B.n17 585
R661 B.n1023 B.n1022 585
R662 B.n1021 B.n18 585
R663 B.n1020 B.n1019 585
R664 B.n1018 B.n19 585
R665 B.n1017 B.n1016 585
R666 B.n1015 B.n20 585
R667 B.n1014 B.n1013 585
R668 B.n1012 B.n21 585
R669 B.n1011 B.n1010 585
R670 B.n1009 B.n22 585
R671 B.n1008 B.n1007 585
R672 B.n1006 B.n23 585
R673 B.n1005 B.n1004 585
R674 B.n1003 B.n24 585
R675 B.n1002 B.n1001 585
R676 B.n1000 B.n25 585
R677 B.n999 B.n998 585
R678 B.n997 B.n26 585
R679 B.n996 B.n995 585
R680 B.n994 B.n27 585
R681 B.n993 B.n992 585
R682 B.n991 B.n28 585
R683 B.n990 B.n989 585
R684 B.n988 B.n29 585
R685 B.n987 B.n986 585
R686 B.n985 B.n30 585
R687 B.n984 B.n983 585
R688 B.n982 B.n31 585
R689 B.n981 B.n980 585
R690 B.n979 B.n32 585
R691 B.n978 B.n977 585
R692 B.n976 B.n33 585
R693 B.n975 B.n974 585
R694 B.n973 B.n34 585
R695 B.n972 B.n971 585
R696 B.n970 B.n35 585
R697 B.n969 B.n968 585
R698 B.n1071 B.n1070 585
R699 B.n377 B.n242 497.305
R700 B.n968 B.n967 497.305
R701 B.n570 B.n569 497.305
R702 B.n775 B.n774 497.305
R703 B.n203 B.t0 324.599
R704 B.n211 B.t9 324.599
R705 B.n66 B.t3 324.599
R706 B.n74 B.t6 324.599
R707 B.n203 B.t2 190.38
R708 B.n74 B.t7 190.38
R709 B.n211 B.t11 190.357
R710 B.n66 B.t4 190.357
R711 B.n373 B.n242 163.367
R712 B.n373 B.n372 163.367
R713 B.n372 B.n371 163.367
R714 B.n371 B.n244 163.367
R715 B.n367 B.n244 163.367
R716 B.n367 B.n366 163.367
R717 B.n366 B.n365 163.367
R718 B.n365 B.n246 163.367
R719 B.n361 B.n246 163.367
R720 B.n361 B.n360 163.367
R721 B.n360 B.n359 163.367
R722 B.n359 B.n248 163.367
R723 B.n355 B.n248 163.367
R724 B.n355 B.n354 163.367
R725 B.n354 B.n353 163.367
R726 B.n353 B.n250 163.367
R727 B.n349 B.n250 163.367
R728 B.n349 B.n348 163.367
R729 B.n348 B.n347 163.367
R730 B.n347 B.n252 163.367
R731 B.n343 B.n252 163.367
R732 B.n343 B.n342 163.367
R733 B.n342 B.n341 163.367
R734 B.n341 B.n254 163.367
R735 B.n337 B.n254 163.367
R736 B.n337 B.n336 163.367
R737 B.n336 B.n335 163.367
R738 B.n335 B.n256 163.367
R739 B.n331 B.n256 163.367
R740 B.n331 B.n330 163.367
R741 B.n330 B.n329 163.367
R742 B.n329 B.n258 163.367
R743 B.n325 B.n258 163.367
R744 B.n325 B.n324 163.367
R745 B.n324 B.n323 163.367
R746 B.n323 B.n260 163.367
R747 B.n319 B.n260 163.367
R748 B.n319 B.n318 163.367
R749 B.n318 B.n317 163.367
R750 B.n317 B.n262 163.367
R751 B.n313 B.n262 163.367
R752 B.n313 B.n312 163.367
R753 B.n312 B.n311 163.367
R754 B.n311 B.n264 163.367
R755 B.n307 B.n264 163.367
R756 B.n307 B.n306 163.367
R757 B.n306 B.n305 163.367
R758 B.n305 B.n266 163.367
R759 B.n301 B.n266 163.367
R760 B.n301 B.n300 163.367
R761 B.n300 B.n299 163.367
R762 B.n299 B.n268 163.367
R763 B.n295 B.n268 163.367
R764 B.n295 B.n294 163.367
R765 B.n294 B.n293 163.367
R766 B.n293 B.n270 163.367
R767 B.n289 B.n270 163.367
R768 B.n289 B.n288 163.367
R769 B.n288 B.n287 163.367
R770 B.n287 B.n272 163.367
R771 B.n283 B.n272 163.367
R772 B.n283 B.n282 163.367
R773 B.n282 B.n281 163.367
R774 B.n281 B.n274 163.367
R775 B.n277 B.n274 163.367
R776 B.n277 B.n276 163.367
R777 B.n276 B.n2 163.367
R778 B.n1070 B.n2 163.367
R779 B.n1070 B.n1069 163.367
R780 B.n1069 B.n1068 163.367
R781 B.n1068 B.n3 163.367
R782 B.n1064 B.n3 163.367
R783 B.n1064 B.n1063 163.367
R784 B.n1063 B.n1062 163.367
R785 B.n1062 B.n5 163.367
R786 B.n1058 B.n5 163.367
R787 B.n1058 B.n1057 163.367
R788 B.n1057 B.n1056 163.367
R789 B.n1056 B.n7 163.367
R790 B.n1052 B.n7 163.367
R791 B.n1052 B.n1051 163.367
R792 B.n1051 B.n1050 163.367
R793 B.n1050 B.n9 163.367
R794 B.n1046 B.n9 163.367
R795 B.n1046 B.n1045 163.367
R796 B.n1045 B.n1044 163.367
R797 B.n1044 B.n11 163.367
R798 B.n1040 B.n11 163.367
R799 B.n1040 B.n1039 163.367
R800 B.n1039 B.n1038 163.367
R801 B.n1038 B.n13 163.367
R802 B.n1034 B.n13 163.367
R803 B.n1034 B.n1033 163.367
R804 B.n1033 B.n1032 163.367
R805 B.n1032 B.n15 163.367
R806 B.n1028 B.n15 163.367
R807 B.n1028 B.n1027 163.367
R808 B.n1027 B.n1026 163.367
R809 B.n1026 B.n17 163.367
R810 B.n1022 B.n17 163.367
R811 B.n1022 B.n1021 163.367
R812 B.n1021 B.n1020 163.367
R813 B.n1020 B.n19 163.367
R814 B.n1016 B.n19 163.367
R815 B.n1016 B.n1015 163.367
R816 B.n1015 B.n1014 163.367
R817 B.n1014 B.n21 163.367
R818 B.n1010 B.n21 163.367
R819 B.n1010 B.n1009 163.367
R820 B.n1009 B.n1008 163.367
R821 B.n1008 B.n23 163.367
R822 B.n1004 B.n23 163.367
R823 B.n1004 B.n1003 163.367
R824 B.n1003 B.n1002 163.367
R825 B.n1002 B.n25 163.367
R826 B.n998 B.n25 163.367
R827 B.n998 B.n997 163.367
R828 B.n997 B.n996 163.367
R829 B.n996 B.n27 163.367
R830 B.n992 B.n27 163.367
R831 B.n992 B.n991 163.367
R832 B.n991 B.n990 163.367
R833 B.n990 B.n29 163.367
R834 B.n986 B.n29 163.367
R835 B.n986 B.n985 163.367
R836 B.n985 B.n984 163.367
R837 B.n984 B.n31 163.367
R838 B.n980 B.n31 163.367
R839 B.n980 B.n979 163.367
R840 B.n979 B.n978 163.367
R841 B.n978 B.n33 163.367
R842 B.n974 B.n33 163.367
R843 B.n974 B.n973 163.367
R844 B.n973 B.n972 163.367
R845 B.n972 B.n35 163.367
R846 B.n968 B.n35 163.367
R847 B.n378 B.n377 163.367
R848 B.n379 B.n378 163.367
R849 B.n379 B.n240 163.367
R850 B.n383 B.n240 163.367
R851 B.n384 B.n383 163.367
R852 B.n385 B.n384 163.367
R853 B.n385 B.n238 163.367
R854 B.n389 B.n238 163.367
R855 B.n390 B.n389 163.367
R856 B.n391 B.n390 163.367
R857 B.n391 B.n236 163.367
R858 B.n395 B.n236 163.367
R859 B.n396 B.n395 163.367
R860 B.n397 B.n396 163.367
R861 B.n397 B.n234 163.367
R862 B.n401 B.n234 163.367
R863 B.n402 B.n401 163.367
R864 B.n403 B.n402 163.367
R865 B.n403 B.n232 163.367
R866 B.n407 B.n232 163.367
R867 B.n408 B.n407 163.367
R868 B.n409 B.n408 163.367
R869 B.n409 B.n230 163.367
R870 B.n413 B.n230 163.367
R871 B.n414 B.n413 163.367
R872 B.n415 B.n414 163.367
R873 B.n415 B.n228 163.367
R874 B.n419 B.n228 163.367
R875 B.n420 B.n419 163.367
R876 B.n421 B.n420 163.367
R877 B.n421 B.n226 163.367
R878 B.n425 B.n226 163.367
R879 B.n426 B.n425 163.367
R880 B.n427 B.n426 163.367
R881 B.n427 B.n224 163.367
R882 B.n431 B.n224 163.367
R883 B.n432 B.n431 163.367
R884 B.n433 B.n432 163.367
R885 B.n433 B.n222 163.367
R886 B.n437 B.n222 163.367
R887 B.n438 B.n437 163.367
R888 B.n439 B.n438 163.367
R889 B.n439 B.n220 163.367
R890 B.n443 B.n220 163.367
R891 B.n444 B.n443 163.367
R892 B.n445 B.n444 163.367
R893 B.n445 B.n218 163.367
R894 B.n449 B.n218 163.367
R895 B.n450 B.n449 163.367
R896 B.n451 B.n450 163.367
R897 B.n451 B.n216 163.367
R898 B.n455 B.n216 163.367
R899 B.n456 B.n455 163.367
R900 B.n457 B.n456 163.367
R901 B.n457 B.n214 163.367
R902 B.n461 B.n214 163.367
R903 B.n462 B.n461 163.367
R904 B.n463 B.n462 163.367
R905 B.n463 B.n210 163.367
R906 B.n468 B.n210 163.367
R907 B.n469 B.n468 163.367
R908 B.n470 B.n469 163.367
R909 B.n470 B.n208 163.367
R910 B.n474 B.n208 163.367
R911 B.n475 B.n474 163.367
R912 B.n476 B.n475 163.367
R913 B.n476 B.n206 163.367
R914 B.n480 B.n206 163.367
R915 B.n481 B.n480 163.367
R916 B.n481 B.n202 163.367
R917 B.n485 B.n202 163.367
R918 B.n486 B.n485 163.367
R919 B.n487 B.n486 163.367
R920 B.n487 B.n200 163.367
R921 B.n491 B.n200 163.367
R922 B.n492 B.n491 163.367
R923 B.n493 B.n492 163.367
R924 B.n493 B.n198 163.367
R925 B.n497 B.n198 163.367
R926 B.n498 B.n497 163.367
R927 B.n499 B.n498 163.367
R928 B.n499 B.n196 163.367
R929 B.n503 B.n196 163.367
R930 B.n504 B.n503 163.367
R931 B.n505 B.n504 163.367
R932 B.n505 B.n194 163.367
R933 B.n509 B.n194 163.367
R934 B.n510 B.n509 163.367
R935 B.n511 B.n510 163.367
R936 B.n511 B.n192 163.367
R937 B.n515 B.n192 163.367
R938 B.n516 B.n515 163.367
R939 B.n517 B.n516 163.367
R940 B.n517 B.n190 163.367
R941 B.n521 B.n190 163.367
R942 B.n522 B.n521 163.367
R943 B.n523 B.n522 163.367
R944 B.n523 B.n188 163.367
R945 B.n527 B.n188 163.367
R946 B.n528 B.n527 163.367
R947 B.n529 B.n528 163.367
R948 B.n529 B.n186 163.367
R949 B.n533 B.n186 163.367
R950 B.n534 B.n533 163.367
R951 B.n535 B.n534 163.367
R952 B.n535 B.n184 163.367
R953 B.n539 B.n184 163.367
R954 B.n540 B.n539 163.367
R955 B.n541 B.n540 163.367
R956 B.n541 B.n182 163.367
R957 B.n545 B.n182 163.367
R958 B.n546 B.n545 163.367
R959 B.n547 B.n546 163.367
R960 B.n547 B.n180 163.367
R961 B.n551 B.n180 163.367
R962 B.n552 B.n551 163.367
R963 B.n553 B.n552 163.367
R964 B.n553 B.n178 163.367
R965 B.n557 B.n178 163.367
R966 B.n558 B.n557 163.367
R967 B.n559 B.n558 163.367
R968 B.n559 B.n176 163.367
R969 B.n563 B.n176 163.367
R970 B.n564 B.n563 163.367
R971 B.n565 B.n564 163.367
R972 B.n565 B.n174 163.367
R973 B.n569 B.n174 163.367
R974 B.n571 B.n570 163.367
R975 B.n571 B.n172 163.367
R976 B.n575 B.n172 163.367
R977 B.n576 B.n575 163.367
R978 B.n577 B.n576 163.367
R979 B.n577 B.n170 163.367
R980 B.n581 B.n170 163.367
R981 B.n582 B.n581 163.367
R982 B.n583 B.n582 163.367
R983 B.n583 B.n168 163.367
R984 B.n587 B.n168 163.367
R985 B.n588 B.n587 163.367
R986 B.n589 B.n588 163.367
R987 B.n589 B.n166 163.367
R988 B.n593 B.n166 163.367
R989 B.n594 B.n593 163.367
R990 B.n595 B.n594 163.367
R991 B.n595 B.n164 163.367
R992 B.n599 B.n164 163.367
R993 B.n600 B.n599 163.367
R994 B.n601 B.n600 163.367
R995 B.n601 B.n162 163.367
R996 B.n605 B.n162 163.367
R997 B.n606 B.n605 163.367
R998 B.n607 B.n606 163.367
R999 B.n607 B.n160 163.367
R1000 B.n611 B.n160 163.367
R1001 B.n612 B.n611 163.367
R1002 B.n613 B.n612 163.367
R1003 B.n613 B.n158 163.367
R1004 B.n617 B.n158 163.367
R1005 B.n618 B.n617 163.367
R1006 B.n619 B.n618 163.367
R1007 B.n619 B.n156 163.367
R1008 B.n623 B.n156 163.367
R1009 B.n624 B.n623 163.367
R1010 B.n625 B.n624 163.367
R1011 B.n625 B.n154 163.367
R1012 B.n629 B.n154 163.367
R1013 B.n630 B.n629 163.367
R1014 B.n631 B.n630 163.367
R1015 B.n631 B.n152 163.367
R1016 B.n635 B.n152 163.367
R1017 B.n636 B.n635 163.367
R1018 B.n637 B.n636 163.367
R1019 B.n637 B.n150 163.367
R1020 B.n641 B.n150 163.367
R1021 B.n642 B.n641 163.367
R1022 B.n643 B.n642 163.367
R1023 B.n643 B.n148 163.367
R1024 B.n647 B.n148 163.367
R1025 B.n648 B.n647 163.367
R1026 B.n649 B.n648 163.367
R1027 B.n649 B.n146 163.367
R1028 B.n653 B.n146 163.367
R1029 B.n654 B.n653 163.367
R1030 B.n655 B.n654 163.367
R1031 B.n655 B.n144 163.367
R1032 B.n659 B.n144 163.367
R1033 B.n660 B.n659 163.367
R1034 B.n661 B.n660 163.367
R1035 B.n661 B.n142 163.367
R1036 B.n665 B.n142 163.367
R1037 B.n666 B.n665 163.367
R1038 B.n667 B.n666 163.367
R1039 B.n667 B.n140 163.367
R1040 B.n671 B.n140 163.367
R1041 B.n672 B.n671 163.367
R1042 B.n673 B.n672 163.367
R1043 B.n673 B.n138 163.367
R1044 B.n677 B.n138 163.367
R1045 B.n678 B.n677 163.367
R1046 B.n679 B.n678 163.367
R1047 B.n679 B.n136 163.367
R1048 B.n683 B.n136 163.367
R1049 B.n684 B.n683 163.367
R1050 B.n685 B.n684 163.367
R1051 B.n685 B.n134 163.367
R1052 B.n689 B.n134 163.367
R1053 B.n690 B.n689 163.367
R1054 B.n691 B.n690 163.367
R1055 B.n691 B.n132 163.367
R1056 B.n695 B.n132 163.367
R1057 B.n696 B.n695 163.367
R1058 B.n697 B.n696 163.367
R1059 B.n697 B.n130 163.367
R1060 B.n701 B.n130 163.367
R1061 B.n702 B.n701 163.367
R1062 B.n703 B.n702 163.367
R1063 B.n703 B.n128 163.367
R1064 B.n707 B.n128 163.367
R1065 B.n708 B.n707 163.367
R1066 B.n709 B.n708 163.367
R1067 B.n709 B.n126 163.367
R1068 B.n713 B.n126 163.367
R1069 B.n714 B.n713 163.367
R1070 B.n715 B.n714 163.367
R1071 B.n715 B.n124 163.367
R1072 B.n719 B.n124 163.367
R1073 B.n720 B.n719 163.367
R1074 B.n721 B.n720 163.367
R1075 B.n721 B.n122 163.367
R1076 B.n725 B.n122 163.367
R1077 B.n726 B.n725 163.367
R1078 B.n727 B.n726 163.367
R1079 B.n727 B.n120 163.367
R1080 B.n731 B.n120 163.367
R1081 B.n732 B.n731 163.367
R1082 B.n733 B.n732 163.367
R1083 B.n733 B.n118 163.367
R1084 B.n737 B.n118 163.367
R1085 B.n738 B.n737 163.367
R1086 B.n739 B.n738 163.367
R1087 B.n739 B.n116 163.367
R1088 B.n743 B.n116 163.367
R1089 B.n744 B.n743 163.367
R1090 B.n745 B.n744 163.367
R1091 B.n745 B.n114 163.367
R1092 B.n749 B.n114 163.367
R1093 B.n750 B.n749 163.367
R1094 B.n751 B.n750 163.367
R1095 B.n751 B.n112 163.367
R1096 B.n755 B.n112 163.367
R1097 B.n756 B.n755 163.367
R1098 B.n757 B.n756 163.367
R1099 B.n757 B.n110 163.367
R1100 B.n761 B.n110 163.367
R1101 B.n762 B.n761 163.367
R1102 B.n763 B.n762 163.367
R1103 B.n763 B.n108 163.367
R1104 B.n767 B.n108 163.367
R1105 B.n768 B.n767 163.367
R1106 B.n769 B.n768 163.367
R1107 B.n769 B.n106 163.367
R1108 B.n773 B.n106 163.367
R1109 B.n774 B.n773 163.367
R1110 B.n967 B.n966 163.367
R1111 B.n966 B.n37 163.367
R1112 B.n962 B.n37 163.367
R1113 B.n962 B.n961 163.367
R1114 B.n961 B.n960 163.367
R1115 B.n960 B.n39 163.367
R1116 B.n956 B.n39 163.367
R1117 B.n956 B.n955 163.367
R1118 B.n955 B.n954 163.367
R1119 B.n954 B.n41 163.367
R1120 B.n950 B.n41 163.367
R1121 B.n950 B.n949 163.367
R1122 B.n949 B.n948 163.367
R1123 B.n948 B.n43 163.367
R1124 B.n944 B.n43 163.367
R1125 B.n944 B.n943 163.367
R1126 B.n943 B.n942 163.367
R1127 B.n942 B.n45 163.367
R1128 B.n938 B.n45 163.367
R1129 B.n938 B.n937 163.367
R1130 B.n937 B.n936 163.367
R1131 B.n936 B.n47 163.367
R1132 B.n932 B.n47 163.367
R1133 B.n932 B.n931 163.367
R1134 B.n931 B.n930 163.367
R1135 B.n930 B.n49 163.367
R1136 B.n926 B.n49 163.367
R1137 B.n926 B.n925 163.367
R1138 B.n925 B.n924 163.367
R1139 B.n924 B.n51 163.367
R1140 B.n920 B.n51 163.367
R1141 B.n920 B.n919 163.367
R1142 B.n919 B.n918 163.367
R1143 B.n918 B.n53 163.367
R1144 B.n914 B.n53 163.367
R1145 B.n914 B.n913 163.367
R1146 B.n913 B.n912 163.367
R1147 B.n912 B.n55 163.367
R1148 B.n908 B.n55 163.367
R1149 B.n908 B.n907 163.367
R1150 B.n907 B.n906 163.367
R1151 B.n906 B.n57 163.367
R1152 B.n902 B.n57 163.367
R1153 B.n902 B.n901 163.367
R1154 B.n901 B.n900 163.367
R1155 B.n900 B.n59 163.367
R1156 B.n896 B.n59 163.367
R1157 B.n896 B.n895 163.367
R1158 B.n895 B.n894 163.367
R1159 B.n894 B.n61 163.367
R1160 B.n890 B.n61 163.367
R1161 B.n890 B.n889 163.367
R1162 B.n889 B.n888 163.367
R1163 B.n888 B.n63 163.367
R1164 B.n884 B.n63 163.367
R1165 B.n884 B.n883 163.367
R1166 B.n883 B.n882 163.367
R1167 B.n882 B.n65 163.367
R1168 B.n877 B.n65 163.367
R1169 B.n877 B.n876 163.367
R1170 B.n876 B.n875 163.367
R1171 B.n875 B.n69 163.367
R1172 B.n871 B.n69 163.367
R1173 B.n871 B.n870 163.367
R1174 B.n870 B.n869 163.367
R1175 B.n869 B.n71 163.367
R1176 B.n865 B.n71 163.367
R1177 B.n865 B.n864 163.367
R1178 B.n864 B.n863 163.367
R1179 B.n863 B.n73 163.367
R1180 B.n859 B.n73 163.367
R1181 B.n859 B.n858 163.367
R1182 B.n858 B.n857 163.367
R1183 B.n857 B.n78 163.367
R1184 B.n853 B.n78 163.367
R1185 B.n853 B.n852 163.367
R1186 B.n852 B.n851 163.367
R1187 B.n851 B.n80 163.367
R1188 B.n847 B.n80 163.367
R1189 B.n847 B.n846 163.367
R1190 B.n846 B.n845 163.367
R1191 B.n845 B.n82 163.367
R1192 B.n841 B.n82 163.367
R1193 B.n841 B.n840 163.367
R1194 B.n840 B.n839 163.367
R1195 B.n839 B.n84 163.367
R1196 B.n835 B.n84 163.367
R1197 B.n835 B.n834 163.367
R1198 B.n834 B.n833 163.367
R1199 B.n833 B.n86 163.367
R1200 B.n829 B.n86 163.367
R1201 B.n829 B.n828 163.367
R1202 B.n828 B.n827 163.367
R1203 B.n827 B.n88 163.367
R1204 B.n823 B.n88 163.367
R1205 B.n823 B.n822 163.367
R1206 B.n822 B.n821 163.367
R1207 B.n821 B.n90 163.367
R1208 B.n817 B.n90 163.367
R1209 B.n817 B.n816 163.367
R1210 B.n816 B.n815 163.367
R1211 B.n815 B.n92 163.367
R1212 B.n811 B.n92 163.367
R1213 B.n811 B.n810 163.367
R1214 B.n810 B.n809 163.367
R1215 B.n809 B.n94 163.367
R1216 B.n805 B.n94 163.367
R1217 B.n805 B.n804 163.367
R1218 B.n804 B.n803 163.367
R1219 B.n803 B.n96 163.367
R1220 B.n799 B.n96 163.367
R1221 B.n799 B.n798 163.367
R1222 B.n798 B.n797 163.367
R1223 B.n797 B.n98 163.367
R1224 B.n793 B.n98 163.367
R1225 B.n793 B.n792 163.367
R1226 B.n792 B.n791 163.367
R1227 B.n791 B.n100 163.367
R1228 B.n787 B.n100 163.367
R1229 B.n787 B.n786 163.367
R1230 B.n786 B.n785 163.367
R1231 B.n785 B.n102 163.367
R1232 B.n781 B.n102 163.367
R1233 B.n781 B.n780 163.367
R1234 B.n780 B.n779 163.367
R1235 B.n779 B.n104 163.367
R1236 B.n775 B.n104 163.367
R1237 B.n204 B.t1 111.252
R1238 B.n75 B.t8 111.252
R1239 B.n212 B.t10 111.23
R1240 B.n67 B.t5 111.23
R1241 B.n204 B.n203 79.1278
R1242 B.n212 B.n211 79.1278
R1243 B.n67 B.n66 79.1278
R1244 B.n75 B.n74 79.1278
R1245 B.n205 B.n204 59.5399
R1246 B.n465 B.n212 59.5399
R1247 B.n879 B.n67 59.5399
R1248 B.n76 B.n75 59.5399
R1249 B.n969 B.n36 32.3127
R1250 B.n776 B.n105 32.3127
R1251 B.n568 B.n173 32.3127
R1252 B.n376 B.n375 32.3127
R1253 B B.n1071 18.0485
R1254 B.n965 B.n36 10.6151
R1255 B.n965 B.n964 10.6151
R1256 B.n964 B.n963 10.6151
R1257 B.n963 B.n38 10.6151
R1258 B.n959 B.n38 10.6151
R1259 B.n959 B.n958 10.6151
R1260 B.n958 B.n957 10.6151
R1261 B.n957 B.n40 10.6151
R1262 B.n953 B.n40 10.6151
R1263 B.n953 B.n952 10.6151
R1264 B.n952 B.n951 10.6151
R1265 B.n951 B.n42 10.6151
R1266 B.n947 B.n42 10.6151
R1267 B.n947 B.n946 10.6151
R1268 B.n946 B.n945 10.6151
R1269 B.n945 B.n44 10.6151
R1270 B.n941 B.n44 10.6151
R1271 B.n941 B.n940 10.6151
R1272 B.n940 B.n939 10.6151
R1273 B.n939 B.n46 10.6151
R1274 B.n935 B.n46 10.6151
R1275 B.n935 B.n934 10.6151
R1276 B.n934 B.n933 10.6151
R1277 B.n933 B.n48 10.6151
R1278 B.n929 B.n48 10.6151
R1279 B.n929 B.n928 10.6151
R1280 B.n928 B.n927 10.6151
R1281 B.n927 B.n50 10.6151
R1282 B.n923 B.n50 10.6151
R1283 B.n923 B.n922 10.6151
R1284 B.n922 B.n921 10.6151
R1285 B.n921 B.n52 10.6151
R1286 B.n917 B.n52 10.6151
R1287 B.n917 B.n916 10.6151
R1288 B.n916 B.n915 10.6151
R1289 B.n915 B.n54 10.6151
R1290 B.n911 B.n54 10.6151
R1291 B.n911 B.n910 10.6151
R1292 B.n910 B.n909 10.6151
R1293 B.n909 B.n56 10.6151
R1294 B.n905 B.n56 10.6151
R1295 B.n905 B.n904 10.6151
R1296 B.n904 B.n903 10.6151
R1297 B.n903 B.n58 10.6151
R1298 B.n899 B.n58 10.6151
R1299 B.n899 B.n898 10.6151
R1300 B.n898 B.n897 10.6151
R1301 B.n897 B.n60 10.6151
R1302 B.n893 B.n60 10.6151
R1303 B.n893 B.n892 10.6151
R1304 B.n892 B.n891 10.6151
R1305 B.n891 B.n62 10.6151
R1306 B.n887 B.n62 10.6151
R1307 B.n887 B.n886 10.6151
R1308 B.n886 B.n885 10.6151
R1309 B.n885 B.n64 10.6151
R1310 B.n881 B.n64 10.6151
R1311 B.n881 B.n880 10.6151
R1312 B.n878 B.n68 10.6151
R1313 B.n874 B.n68 10.6151
R1314 B.n874 B.n873 10.6151
R1315 B.n873 B.n872 10.6151
R1316 B.n872 B.n70 10.6151
R1317 B.n868 B.n70 10.6151
R1318 B.n868 B.n867 10.6151
R1319 B.n867 B.n866 10.6151
R1320 B.n866 B.n72 10.6151
R1321 B.n862 B.n861 10.6151
R1322 B.n861 B.n860 10.6151
R1323 B.n860 B.n77 10.6151
R1324 B.n856 B.n77 10.6151
R1325 B.n856 B.n855 10.6151
R1326 B.n855 B.n854 10.6151
R1327 B.n854 B.n79 10.6151
R1328 B.n850 B.n79 10.6151
R1329 B.n850 B.n849 10.6151
R1330 B.n849 B.n848 10.6151
R1331 B.n848 B.n81 10.6151
R1332 B.n844 B.n81 10.6151
R1333 B.n844 B.n843 10.6151
R1334 B.n843 B.n842 10.6151
R1335 B.n842 B.n83 10.6151
R1336 B.n838 B.n83 10.6151
R1337 B.n838 B.n837 10.6151
R1338 B.n837 B.n836 10.6151
R1339 B.n836 B.n85 10.6151
R1340 B.n832 B.n85 10.6151
R1341 B.n832 B.n831 10.6151
R1342 B.n831 B.n830 10.6151
R1343 B.n830 B.n87 10.6151
R1344 B.n826 B.n87 10.6151
R1345 B.n826 B.n825 10.6151
R1346 B.n825 B.n824 10.6151
R1347 B.n824 B.n89 10.6151
R1348 B.n820 B.n89 10.6151
R1349 B.n820 B.n819 10.6151
R1350 B.n819 B.n818 10.6151
R1351 B.n818 B.n91 10.6151
R1352 B.n814 B.n91 10.6151
R1353 B.n814 B.n813 10.6151
R1354 B.n813 B.n812 10.6151
R1355 B.n812 B.n93 10.6151
R1356 B.n808 B.n93 10.6151
R1357 B.n808 B.n807 10.6151
R1358 B.n807 B.n806 10.6151
R1359 B.n806 B.n95 10.6151
R1360 B.n802 B.n95 10.6151
R1361 B.n802 B.n801 10.6151
R1362 B.n801 B.n800 10.6151
R1363 B.n800 B.n97 10.6151
R1364 B.n796 B.n97 10.6151
R1365 B.n796 B.n795 10.6151
R1366 B.n795 B.n794 10.6151
R1367 B.n794 B.n99 10.6151
R1368 B.n790 B.n99 10.6151
R1369 B.n790 B.n789 10.6151
R1370 B.n789 B.n788 10.6151
R1371 B.n788 B.n101 10.6151
R1372 B.n784 B.n101 10.6151
R1373 B.n784 B.n783 10.6151
R1374 B.n783 B.n782 10.6151
R1375 B.n782 B.n103 10.6151
R1376 B.n778 B.n103 10.6151
R1377 B.n778 B.n777 10.6151
R1378 B.n777 B.n776 10.6151
R1379 B.n572 B.n173 10.6151
R1380 B.n573 B.n572 10.6151
R1381 B.n574 B.n573 10.6151
R1382 B.n574 B.n171 10.6151
R1383 B.n578 B.n171 10.6151
R1384 B.n579 B.n578 10.6151
R1385 B.n580 B.n579 10.6151
R1386 B.n580 B.n169 10.6151
R1387 B.n584 B.n169 10.6151
R1388 B.n585 B.n584 10.6151
R1389 B.n586 B.n585 10.6151
R1390 B.n586 B.n167 10.6151
R1391 B.n590 B.n167 10.6151
R1392 B.n591 B.n590 10.6151
R1393 B.n592 B.n591 10.6151
R1394 B.n592 B.n165 10.6151
R1395 B.n596 B.n165 10.6151
R1396 B.n597 B.n596 10.6151
R1397 B.n598 B.n597 10.6151
R1398 B.n598 B.n163 10.6151
R1399 B.n602 B.n163 10.6151
R1400 B.n603 B.n602 10.6151
R1401 B.n604 B.n603 10.6151
R1402 B.n604 B.n161 10.6151
R1403 B.n608 B.n161 10.6151
R1404 B.n609 B.n608 10.6151
R1405 B.n610 B.n609 10.6151
R1406 B.n610 B.n159 10.6151
R1407 B.n614 B.n159 10.6151
R1408 B.n615 B.n614 10.6151
R1409 B.n616 B.n615 10.6151
R1410 B.n616 B.n157 10.6151
R1411 B.n620 B.n157 10.6151
R1412 B.n621 B.n620 10.6151
R1413 B.n622 B.n621 10.6151
R1414 B.n622 B.n155 10.6151
R1415 B.n626 B.n155 10.6151
R1416 B.n627 B.n626 10.6151
R1417 B.n628 B.n627 10.6151
R1418 B.n628 B.n153 10.6151
R1419 B.n632 B.n153 10.6151
R1420 B.n633 B.n632 10.6151
R1421 B.n634 B.n633 10.6151
R1422 B.n634 B.n151 10.6151
R1423 B.n638 B.n151 10.6151
R1424 B.n639 B.n638 10.6151
R1425 B.n640 B.n639 10.6151
R1426 B.n640 B.n149 10.6151
R1427 B.n644 B.n149 10.6151
R1428 B.n645 B.n644 10.6151
R1429 B.n646 B.n645 10.6151
R1430 B.n646 B.n147 10.6151
R1431 B.n650 B.n147 10.6151
R1432 B.n651 B.n650 10.6151
R1433 B.n652 B.n651 10.6151
R1434 B.n652 B.n145 10.6151
R1435 B.n656 B.n145 10.6151
R1436 B.n657 B.n656 10.6151
R1437 B.n658 B.n657 10.6151
R1438 B.n658 B.n143 10.6151
R1439 B.n662 B.n143 10.6151
R1440 B.n663 B.n662 10.6151
R1441 B.n664 B.n663 10.6151
R1442 B.n664 B.n141 10.6151
R1443 B.n668 B.n141 10.6151
R1444 B.n669 B.n668 10.6151
R1445 B.n670 B.n669 10.6151
R1446 B.n670 B.n139 10.6151
R1447 B.n674 B.n139 10.6151
R1448 B.n675 B.n674 10.6151
R1449 B.n676 B.n675 10.6151
R1450 B.n676 B.n137 10.6151
R1451 B.n680 B.n137 10.6151
R1452 B.n681 B.n680 10.6151
R1453 B.n682 B.n681 10.6151
R1454 B.n682 B.n135 10.6151
R1455 B.n686 B.n135 10.6151
R1456 B.n687 B.n686 10.6151
R1457 B.n688 B.n687 10.6151
R1458 B.n688 B.n133 10.6151
R1459 B.n692 B.n133 10.6151
R1460 B.n693 B.n692 10.6151
R1461 B.n694 B.n693 10.6151
R1462 B.n694 B.n131 10.6151
R1463 B.n698 B.n131 10.6151
R1464 B.n699 B.n698 10.6151
R1465 B.n700 B.n699 10.6151
R1466 B.n700 B.n129 10.6151
R1467 B.n704 B.n129 10.6151
R1468 B.n705 B.n704 10.6151
R1469 B.n706 B.n705 10.6151
R1470 B.n706 B.n127 10.6151
R1471 B.n710 B.n127 10.6151
R1472 B.n711 B.n710 10.6151
R1473 B.n712 B.n711 10.6151
R1474 B.n712 B.n125 10.6151
R1475 B.n716 B.n125 10.6151
R1476 B.n717 B.n716 10.6151
R1477 B.n718 B.n717 10.6151
R1478 B.n718 B.n123 10.6151
R1479 B.n722 B.n123 10.6151
R1480 B.n723 B.n722 10.6151
R1481 B.n724 B.n723 10.6151
R1482 B.n724 B.n121 10.6151
R1483 B.n728 B.n121 10.6151
R1484 B.n729 B.n728 10.6151
R1485 B.n730 B.n729 10.6151
R1486 B.n730 B.n119 10.6151
R1487 B.n734 B.n119 10.6151
R1488 B.n735 B.n734 10.6151
R1489 B.n736 B.n735 10.6151
R1490 B.n736 B.n117 10.6151
R1491 B.n740 B.n117 10.6151
R1492 B.n741 B.n740 10.6151
R1493 B.n742 B.n741 10.6151
R1494 B.n742 B.n115 10.6151
R1495 B.n746 B.n115 10.6151
R1496 B.n747 B.n746 10.6151
R1497 B.n748 B.n747 10.6151
R1498 B.n748 B.n113 10.6151
R1499 B.n752 B.n113 10.6151
R1500 B.n753 B.n752 10.6151
R1501 B.n754 B.n753 10.6151
R1502 B.n754 B.n111 10.6151
R1503 B.n758 B.n111 10.6151
R1504 B.n759 B.n758 10.6151
R1505 B.n760 B.n759 10.6151
R1506 B.n760 B.n109 10.6151
R1507 B.n764 B.n109 10.6151
R1508 B.n765 B.n764 10.6151
R1509 B.n766 B.n765 10.6151
R1510 B.n766 B.n107 10.6151
R1511 B.n770 B.n107 10.6151
R1512 B.n771 B.n770 10.6151
R1513 B.n772 B.n771 10.6151
R1514 B.n772 B.n105 10.6151
R1515 B.n376 B.n241 10.6151
R1516 B.n380 B.n241 10.6151
R1517 B.n381 B.n380 10.6151
R1518 B.n382 B.n381 10.6151
R1519 B.n382 B.n239 10.6151
R1520 B.n386 B.n239 10.6151
R1521 B.n387 B.n386 10.6151
R1522 B.n388 B.n387 10.6151
R1523 B.n388 B.n237 10.6151
R1524 B.n392 B.n237 10.6151
R1525 B.n393 B.n392 10.6151
R1526 B.n394 B.n393 10.6151
R1527 B.n394 B.n235 10.6151
R1528 B.n398 B.n235 10.6151
R1529 B.n399 B.n398 10.6151
R1530 B.n400 B.n399 10.6151
R1531 B.n400 B.n233 10.6151
R1532 B.n404 B.n233 10.6151
R1533 B.n405 B.n404 10.6151
R1534 B.n406 B.n405 10.6151
R1535 B.n406 B.n231 10.6151
R1536 B.n410 B.n231 10.6151
R1537 B.n411 B.n410 10.6151
R1538 B.n412 B.n411 10.6151
R1539 B.n412 B.n229 10.6151
R1540 B.n416 B.n229 10.6151
R1541 B.n417 B.n416 10.6151
R1542 B.n418 B.n417 10.6151
R1543 B.n418 B.n227 10.6151
R1544 B.n422 B.n227 10.6151
R1545 B.n423 B.n422 10.6151
R1546 B.n424 B.n423 10.6151
R1547 B.n424 B.n225 10.6151
R1548 B.n428 B.n225 10.6151
R1549 B.n429 B.n428 10.6151
R1550 B.n430 B.n429 10.6151
R1551 B.n430 B.n223 10.6151
R1552 B.n434 B.n223 10.6151
R1553 B.n435 B.n434 10.6151
R1554 B.n436 B.n435 10.6151
R1555 B.n436 B.n221 10.6151
R1556 B.n440 B.n221 10.6151
R1557 B.n441 B.n440 10.6151
R1558 B.n442 B.n441 10.6151
R1559 B.n442 B.n219 10.6151
R1560 B.n446 B.n219 10.6151
R1561 B.n447 B.n446 10.6151
R1562 B.n448 B.n447 10.6151
R1563 B.n448 B.n217 10.6151
R1564 B.n452 B.n217 10.6151
R1565 B.n453 B.n452 10.6151
R1566 B.n454 B.n453 10.6151
R1567 B.n454 B.n215 10.6151
R1568 B.n458 B.n215 10.6151
R1569 B.n459 B.n458 10.6151
R1570 B.n460 B.n459 10.6151
R1571 B.n460 B.n213 10.6151
R1572 B.n464 B.n213 10.6151
R1573 B.n467 B.n466 10.6151
R1574 B.n467 B.n209 10.6151
R1575 B.n471 B.n209 10.6151
R1576 B.n472 B.n471 10.6151
R1577 B.n473 B.n472 10.6151
R1578 B.n473 B.n207 10.6151
R1579 B.n477 B.n207 10.6151
R1580 B.n478 B.n477 10.6151
R1581 B.n479 B.n478 10.6151
R1582 B.n483 B.n482 10.6151
R1583 B.n484 B.n483 10.6151
R1584 B.n484 B.n201 10.6151
R1585 B.n488 B.n201 10.6151
R1586 B.n489 B.n488 10.6151
R1587 B.n490 B.n489 10.6151
R1588 B.n490 B.n199 10.6151
R1589 B.n494 B.n199 10.6151
R1590 B.n495 B.n494 10.6151
R1591 B.n496 B.n495 10.6151
R1592 B.n496 B.n197 10.6151
R1593 B.n500 B.n197 10.6151
R1594 B.n501 B.n500 10.6151
R1595 B.n502 B.n501 10.6151
R1596 B.n502 B.n195 10.6151
R1597 B.n506 B.n195 10.6151
R1598 B.n507 B.n506 10.6151
R1599 B.n508 B.n507 10.6151
R1600 B.n508 B.n193 10.6151
R1601 B.n512 B.n193 10.6151
R1602 B.n513 B.n512 10.6151
R1603 B.n514 B.n513 10.6151
R1604 B.n514 B.n191 10.6151
R1605 B.n518 B.n191 10.6151
R1606 B.n519 B.n518 10.6151
R1607 B.n520 B.n519 10.6151
R1608 B.n520 B.n189 10.6151
R1609 B.n524 B.n189 10.6151
R1610 B.n525 B.n524 10.6151
R1611 B.n526 B.n525 10.6151
R1612 B.n526 B.n187 10.6151
R1613 B.n530 B.n187 10.6151
R1614 B.n531 B.n530 10.6151
R1615 B.n532 B.n531 10.6151
R1616 B.n532 B.n185 10.6151
R1617 B.n536 B.n185 10.6151
R1618 B.n537 B.n536 10.6151
R1619 B.n538 B.n537 10.6151
R1620 B.n538 B.n183 10.6151
R1621 B.n542 B.n183 10.6151
R1622 B.n543 B.n542 10.6151
R1623 B.n544 B.n543 10.6151
R1624 B.n544 B.n181 10.6151
R1625 B.n548 B.n181 10.6151
R1626 B.n549 B.n548 10.6151
R1627 B.n550 B.n549 10.6151
R1628 B.n550 B.n179 10.6151
R1629 B.n554 B.n179 10.6151
R1630 B.n555 B.n554 10.6151
R1631 B.n556 B.n555 10.6151
R1632 B.n556 B.n177 10.6151
R1633 B.n560 B.n177 10.6151
R1634 B.n561 B.n560 10.6151
R1635 B.n562 B.n561 10.6151
R1636 B.n562 B.n175 10.6151
R1637 B.n566 B.n175 10.6151
R1638 B.n567 B.n566 10.6151
R1639 B.n568 B.n567 10.6151
R1640 B.n375 B.n374 10.6151
R1641 B.n374 B.n243 10.6151
R1642 B.n370 B.n243 10.6151
R1643 B.n370 B.n369 10.6151
R1644 B.n369 B.n368 10.6151
R1645 B.n368 B.n245 10.6151
R1646 B.n364 B.n245 10.6151
R1647 B.n364 B.n363 10.6151
R1648 B.n363 B.n362 10.6151
R1649 B.n362 B.n247 10.6151
R1650 B.n358 B.n247 10.6151
R1651 B.n358 B.n357 10.6151
R1652 B.n357 B.n356 10.6151
R1653 B.n356 B.n249 10.6151
R1654 B.n352 B.n249 10.6151
R1655 B.n352 B.n351 10.6151
R1656 B.n351 B.n350 10.6151
R1657 B.n350 B.n251 10.6151
R1658 B.n346 B.n251 10.6151
R1659 B.n346 B.n345 10.6151
R1660 B.n345 B.n344 10.6151
R1661 B.n344 B.n253 10.6151
R1662 B.n340 B.n253 10.6151
R1663 B.n340 B.n339 10.6151
R1664 B.n339 B.n338 10.6151
R1665 B.n338 B.n255 10.6151
R1666 B.n334 B.n255 10.6151
R1667 B.n334 B.n333 10.6151
R1668 B.n333 B.n332 10.6151
R1669 B.n332 B.n257 10.6151
R1670 B.n328 B.n257 10.6151
R1671 B.n328 B.n327 10.6151
R1672 B.n327 B.n326 10.6151
R1673 B.n326 B.n259 10.6151
R1674 B.n322 B.n259 10.6151
R1675 B.n322 B.n321 10.6151
R1676 B.n321 B.n320 10.6151
R1677 B.n320 B.n261 10.6151
R1678 B.n316 B.n261 10.6151
R1679 B.n316 B.n315 10.6151
R1680 B.n315 B.n314 10.6151
R1681 B.n314 B.n263 10.6151
R1682 B.n310 B.n263 10.6151
R1683 B.n310 B.n309 10.6151
R1684 B.n309 B.n308 10.6151
R1685 B.n308 B.n265 10.6151
R1686 B.n304 B.n265 10.6151
R1687 B.n304 B.n303 10.6151
R1688 B.n303 B.n302 10.6151
R1689 B.n302 B.n267 10.6151
R1690 B.n298 B.n267 10.6151
R1691 B.n298 B.n297 10.6151
R1692 B.n297 B.n296 10.6151
R1693 B.n296 B.n269 10.6151
R1694 B.n292 B.n269 10.6151
R1695 B.n292 B.n291 10.6151
R1696 B.n291 B.n290 10.6151
R1697 B.n290 B.n271 10.6151
R1698 B.n286 B.n271 10.6151
R1699 B.n286 B.n285 10.6151
R1700 B.n285 B.n284 10.6151
R1701 B.n284 B.n273 10.6151
R1702 B.n280 B.n273 10.6151
R1703 B.n280 B.n279 10.6151
R1704 B.n279 B.n278 10.6151
R1705 B.n278 B.n275 10.6151
R1706 B.n275 B.n0 10.6151
R1707 B.n1067 B.n1 10.6151
R1708 B.n1067 B.n1066 10.6151
R1709 B.n1066 B.n1065 10.6151
R1710 B.n1065 B.n4 10.6151
R1711 B.n1061 B.n4 10.6151
R1712 B.n1061 B.n1060 10.6151
R1713 B.n1060 B.n1059 10.6151
R1714 B.n1059 B.n6 10.6151
R1715 B.n1055 B.n6 10.6151
R1716 B.n1055 B.n1054 10.6151
R1717 B.n1054 B.n1053 10.6151
R1718 B.n1053 B.n8 10.6151
R1719 B.n1049 B.n8 10.6151
R1720 B.n1049 B.n1048 10.6151
R1721 B.n1048 B.n1047 10.6151
R1722 B.n1047 B.n10 10.6151
R1723 B.n1043 B.n10 10.6151
R1724 B.n1043 B.n1042 10.6151
R1725 B.n1042 B.n1041 10.6151
R1726 B.n1041 B.n12 10.6151
R1727 B.n1037 B.n12 10.6151
R1728 B.n1037 B.n1036 10.6151
R1729 B.n1036 B.n1035 10.6151
R1730 B.n1035 B.n14 10.6151
R1731 B.n1031 B.n14 10.6151
R1732 B.n1031 B.n1030 10.6151
R1733 B.n1030 B.n1029 10.6151
R1734 B.n1029 B.n16 10.6151
R1735 B.n1025 B.n16 10.6151
R1736 B.n1025 B.n1024 10.6151
R1737 B.n1024 B.n1023 10.6151
R1738 B.n1023 B.n18 10.6151
R1739 B.n1019 B.n18 10.6151
R1740 B.n1019 B.n1018 10.6151
R1741 B.n1018 B.n1017 10.6151
R1742 B.n1017 B.n20 10.6151
R1743 B.n1013 B.n20 10.6151
R1744 B.n1013 B.n1012 10.6151
R1745 B.n1012 B.n1011 10.6151
R1746 B.n1011 B.n22 10.6151
R1747 B.n1007 B.n22 10.6151
R1748 B.n1007 B.n1006 10.6151
R1749 B.n1006 B.n1005 10.6151
R1750 B.n1005 B.n24 10.6151
R1751 B.n1001 B.n24 10.6151
R1752 B.n1001 B.n1000 10.6151
R1753 B.n1000 B.n999 10.6151
R1754 B.n999 B.n26 10.6151
R1755 B.n995 B.n26 10.6151
R1756 B.n995 B.n994 10.6151
R1757 B.n994 B.n993 10.6151
R1758 B.n993 B.n28 10.6151
R1759 B.n989 B.n28 10.6151
R1760 B.n989 B.n988 10.6151
R1761 B.n988 B.n987 10.6151
R1762 B.n987 B.n30 10.6151
R1763 B.n983 B.n30 10.6151
R1764 B.n983 B.n982 10.6151
R1765 B.n982 B.n981 10.6151
R1766 B.n981 B.n32 10.6151
R1767 B.n977 B.n32 10.6151
R1768 B.n977 B.n976 10.6151
R1769 B.n976 B.n975 10.6151
R1770 B.n975 B.n34 10.6151
R1771 B.n971 B.n34 10.6151
R1772 B.n971 B.n970 10.6151
R1773 B.n970 B.n969 10.6151
R1774 B.n880 B.n879 9.36635
R1775 B.n862 B.n76 9.36635
R1776 B.n465 B.n464 9.36635
R1777 B.n482 B.n205 9.36635
R1778 B.n1071 B.n0 2.81026
R1779 B.n1071 B.n1 2.81026
R1780 B.n879 B.n878 1.24928
R1781 B.n76 B.n72 1.24928
R1782 B.n466 B.n465 1.24928
R1783 B.n479 B.n205 1.24928
R1784 VP.n25 VP.n24 161.3
R1785 VP.n26 VP.n21 161.3
R1786 VP.n28 VP.n27 161.3
R1787 VP.n29 VP.n20 161.3
R1788 VP.n31 VP.n30 161.3
R1789 VP.n32 VP.n19 161.3
R1790 VP.n34 VP.n33 161.3
R1791 VP.n35 VP.n18 161.3
R1792 VP.n38 VP.n37 161.3
R1793 VP.n39 VP.n17 161.3
R1794 VP.n41 VP.n40 161.3
R1795 VP.n42 VP.n16 161.3
R1796 VP.n44 VP.n43 161.3
R1797 VP.n45 VP.n15 161.3
R1798 VP.n47 VP.n46 161.3
R1799 VP.n48 VP.n14 161.3
R1800 VP.n50 VP.n49 161.3
R1801 VP.n93 VP.n92 161.3
R1802 VP.n91 VP.n1 161.3
R1803 VP.n90 VP.n89 161.3
R1804 VP.n88 VP.n2 161.3
R1805 VP.n87 VP.n86 161.3
R1806 VP.n85 VP.n3 161.3
R1807 VP.n84 VP.n83 161.3
R1808 VP.n82 VP.n4 161.3
R1809 VP.n81 VP.n80 161.3
R1810 VP.n78 VP.n5 161.3
R1811 VP.n77 VP.n76 161.3
R1812 VP.n75 VP.n6 161.3
R1813 VP.n74 VP.n73 161.3
R1814 VP.n72 VP.n7 161.3
R1815 VP.n71 VP.n70 161.3
R1816 VP.n69 VP.n8 161.3
R1817 VP.n68 VP.n67 161.3
R1818 VP.n65 VP.n9 161.3
R1819 VP.n64 VP.n63 161.3
R1820 VP.n62 VP.n10 161.3
R1821 VP.n61 VP.n60 161.3
R1822 VP.n59 VP.n11 161.3
R1823 VP.n58 VP.n57 161.3
R1824 VP.n56 VP.n12 161.3
R1825 VP.n55 VP.n54 161.3
R1826 VP.n22 VP.t7 147.802
R1827 VP.n53 VP.t1 115.294
R1828 VP.n66 VP.t4 115.294
R1829 VP.n79 VP.t6 115.294
R1830 VP.n0 VP.t2 115.294
R1831 VP.n13 VP.t5 115.294
R1832 VP.n36 VP.t3 115.294
R1833 VP.n23 VP.t0 115.294
R1834 VP.n53 VP.n52 84.0486
R1835 VP.n94 VP.n0 84.0486
R1836 VP.n51 VP.n13 84.0486
R1837 VP.n23 VP.n22 72.7154
R1838 VP.n52 VP.n51 60.8628
R1839 VP.n60 VP.n59 48.2005
R1840 VP.n86 VP.n2 48.2005
R1841 VP.n43 VP.n15 48.2005
R1842 VP.n73 VP.n72 40.4106
R1843 VP.n73 VP.n6 40.4106
R1844 VP.n30 VP.n19 40.4106
R1845 VP.n30 VP.n29 40.4106
R1846 VP.n60 VP.n10 32.6207
R1847 VP.n86 VP.n85 32.6207
R1848 VP.n43 VP.n42 32.6207
R1849 VP.n54 VP.n12 24.3439
R1850 VP.n58 VP.n12 24.3439
R1851 VP.n59 VP.n58 24.3439
R1852 VP.n64 VP.n10 24.3439
R1853 VP.n65 VP.n64 24.3439
R1854 VP.n67 VP.n8 24.3439
R1855 VP.n71 VP.n8 24.3439
R1856 VP.n72 VP.n71 24.3439
R1857 VP.n77 VP.n6 24.3439
R1858 VP.n78 VP.n77 24.3439
R1859 VP.n80 VP.n78 24.3439
R1860 VP.n84 VP.n4 24.3439
R1861 VP.n85 VP.n84 24.3439
R1862 VP.n90 VP.n2 24.3439
R1863 VP.n91 VP.n90 24.3439
R1864 VP.n92 VP.n91 24.3439
R1865 VP.n47 VP.n15 24.3439
R1866 VP.n48 VP.n47 24.3439
R1867 VP.n49 VP.n48 24.3439
R1868 VP.n34 VP.n19 24.3439
R1869 VP.n35 VP.n34 24.3439
R1870 VP.n37 VP.n35 24.3439
R1871 VP.n41 VP.n17 24.3439
R1872 VP.n42 VP.n41 24.3439
R1873 VP.n24 VP.n21 24.3439
R1874 VP.n28 VP.n21 24.3439
R1875 VP.n29 VP.n28 24.3439
R1876 VP.n66 VP.n65 22.3965
R1877 VP.n79 VP.n4 22.3965
R1878 VP.n36 VP.n17 22.3965
R1879 VP.n54 VP.n53 5.84292
R1880 VP.n92 VP.n0 5.84292
R1881 VP.n49 VP.n13 5.84292
R1882 VP.n25 VP.n22 3.29533
R1883 VP.n67 VP.n66 1.94797
R1884 VP.n80 VP.n79 1.94797
R1885 VP.n37 VP.n36 1.94797
R1886 VP.n24 VP.n23 1.94797
R1887 VP.n51 VP.n50 0.355081
R1888 VP.n55 VP.n52 0.355081
R1889 VP.n94 VP.n93 0.355081
R1890 VP VP.n94 0.26685
R1891 VP.n26 VP.n25 0.189894
R1892 VP.n27 VP.n26 0.189894
R1893 VP.n27 VP.n20 0.189894
R1894 VP.n31 VP.n20 0.189894
R1895 VP.n32 VP.n31 0.189894
R1896 VP.n33 VP.n32 0.189894
R1897 VP.n33 VP.n18 0.189894
R1898 VP.n38 VP.n18 0.189894
R1899 VP.n39 VP.n38 0.189894
R1900 VP.n40 VP.n39 0.189894
R1901 VP.n40 VP.n16 0.189894
R1902 VP.n44 VP.n16 0.189894
R1903 VP.n45 VP.n44 0.189894
R1904 VP.n46 VP.n45 0.189894
R1905 VP.n46 VP.n14 0.189894
R1906 VP.n50 VP.n14 0.189894
R1907 VP.n56 VP.n55 0.189894
R1908 VP.n57 VP.n56 0.189894
R1909 VP.n57 VP.n11 0.189894
R1910 VP.n61 VP.n11 0.189894
R1911 VP.n62 VP.n61 0.189894
R1912 VP.n63 VP.n62 0.189894
R1913 VP.n63 VP.n9 0.189894
R1914 VP.n68 VP.n9 0.189894
R1915 VP.n69 VP.n68 0.189894
R1916 VP.n70 VP.n69 0.189894
R1917 VP.n70 VP.n7 0.189894
R1918 VP.n74 VP.n7 0.189894
R1919 VP.n75 VP.n74 0.189894
R1920 VP.n76 VP.n75 0.189894
R1921 VP.n76 VP.n5 0.189894
R1922 VP.n81 VP.n5 0.189894
R1923 VP.n82 VP.n81 0.189894
R1924 VP.n83 VP.n82 0.189894
R1925 VP.n83 VP.n3 0.189894
R1926 VP.n87 VP.n3 0.189894
R1927 VP.n88 VP.n87 0.189894
R1928 VP.n89 VP.n88 0.189894
R1929 VP.n89 VP.n1 0.189894
R1930 VP.n93 VP.n1 0.189894
R1931 VDD1 VDD1.n0 71.8311
R1932 VDD1.n3 VDD1.n2 71.7174
R1933 VDD1.n3 VDD1.n1 71.7174
R1934 VDD1.n5 VDD1.n4 70.0141
R1935 VDD1.n5 VDD1.n3 55.5914
R1936 VDD1.n4 VDD1.t4 1.81237
R1937 VDD1.n4 VDD1.t2 1.81237
R1938 VDD1.n0 VDD1.t0 1.81237
R1939 VDD1.n0 VDD1.t7 1.81237
R1940 VDD1.n2 VDD1.t1 1.81237
R1941 VDD1.n2 VDD1.t5 1.81237
R1942 VDD1.n1 VDD1.t6 1.81237
R1943 VDD1.n1 VDD1.t3 1.81237
R1944 VDD1 VDD1.n5 1.70093
C0 VTAIL VDD1 10.2312f
C1 w_n5050_n4556# VP 11.3831f
C2 VDD2 w_n5050_n4556# 2.64362f
C3 VDD2 VP 0.641537f
C4 VTAIL B 7.509359f
C5 B VDD1 2.16071f
C6 VN w_n5050_n4556# 10.7242f
C7 VN VP 10.1766f
C8 VN VDD2 13.5839f
C9 VTAIL w_n5050_n4556# 5.59429f
C10 VTAIL VP 14.0966f
C11 w_n5050_n4556# VDD1 2.48067f
C12 VDD1 VP 14.0702f
C13 VTAIL VDD2 10.2934f
C14 VDD2 VDD1 2.37298f
C15 VTAIL VN 14.0825f
C16 VN VDD1 0.153301f
C17 w_n5050_n4556# B 13.540901f
C18 B VP 2.66869f
C19 VDD2 B 2.29292f
C20 VN B 1.55787f
C21 VDD2 VSUBS 2.57555f
C22 VDD1 VSUBS 3.42298f
C23 VTAIL VSUBS 1.806974f
C24 VN VSUBS 8.47009f
C25 VP VSUBS 4.977206f
C26 B VSUBS 6.78732f
C27 w_n5050_n4556# VSUBS 0.281366p
C28 VDD1.t0 VSUBS 0.446605f
C29 VDD1.t7 VSUBS 0.446605f
C30 VDD1.n0 VSUBS 3.7438f
C31 VDD1.t6 VSUBS 0.446605f
C32 VDD1.t3 VSUBS 0.446605f
C33 VDD1.n1 VSUBS 3.74173f
C34 VDD1.t1 VSUBS 0.446605f
C35 VDD1.t5 VSUBS 0.446605f
C36 VDD1.n2 VSUBS 3.74173f
C37 VDD1.n3 VSUBS 6.20941f
C38 VDD1.t4 VSUBS 0.446605f
C39 VDD1.t2 VSUBS 0.446605f
C40 VDD1.n4 VSUBS 3.7142f
C41 VDD1.n5 VSUBS 5.17924f
C42 VP.t2 VSUBS 4.22006f
C43 VP.n0 VSUBS 1.54326f
C44 VP.n1 VSUBS 0.022807f
C45 VP.n2 VSUBS 0.042928f
C46 VP.n3 VSUBS 0.022807f
C47 VP.n4 VSUBS 0.041032f
C48 VP.n5 VSUBS 0.022807f
C49 VP.n6 VSUBS 0.045571f
C50 VP.n7 VSUBS 0.022807f
C51 VP.n8 VSUBS 0.04272f
C52 VP.n9 VSUBS 0.022807f
C53 VP.t4 VSUBS 4.22006f
C54 VP.n10 VSUBS 0.046252f
C55 VP.n11 VSUBS 0.022807f
C56 VP.n12 VSUBS 0.04272f
C57 VP.t5 VSUBS 4.22006f
C58 VP.n13 VSUBS 1.54326f
C59 VP.n14 VSUBS 0.022807f
C60 VP.n15 VSUBS 0.042928f
C61 VP.n16 VSUBS 0.022807f
C62 VP.n17 VSUBS 0.041032f
C63 VP.n18 VSUBS 0.022807f
C64 VP.n19 VSUBS 0.045571f
C65 VP.n20 VSUBS 0.022807f
C66 VP.n21 VSUBS 0.04272f
C67 VP.t7 VSUBS 4.57887f
C68 VP.n22 VSUBS 1.46108f
C69 VP.t0 VSUBS 4.22006f
C70 VP.n23 VSUBS 1.52814f
C71 VP.n24 VSUBS 0.023315f
C72 VP.n25 VSUBS 0.290619f
C73 VP.n26 VSUBS 0.022807f
C74 VP.n27 VSUBS 0.022807f
C75 VP.n28 VSUBS 0.04272f
C76 VP.n29 VSUBS 0.045571f
C77 VP.n30 VSUBS 0.018456f
C78 VP.n31 VSUBS 0.022807f
C79 VP.n32 VSUBS 0.022807f
C80 VP.n33 VSUBS 0.022807f
C81 VP.n34 VSUBS 0.04272f
C82 VP.n35 VSUBS 0.04272f
C83 VP.t3 VSUBS 4.22006f
C84 VP.n36 VSUBS 1.45441f
C85 VP.n37 VSUBS 0.023315f
C86 VP.n38 VSUBS 0.022807f
C87 VP.n39 VSUBS 0.022807f
C88 VP.n40 VSUBS 0.022807f
C89 VP.n41 VSUBS 0.04272f
C90 VP.n42 VSUBS 0.046252f
C91 VP.n43 VSUBS 0.020417f
C92 VP.n44 VSUBS 0.022807f
C93 VP.n45 VSUBS 0.022807f
C94 VP.n46 VSUBS 0.022807f
C95 VP.n47 VSUBS 0.04272f
C96 VP.n48 VSUBS 0.04272f
C97 VP.n49 VSUBS 0.02669f
C98 VP.n50 VSUBS 0.036816f
C99 VP.n51 VSUBS 1.71522f
C100 VP.n52 VSUBS 1.72866f
C101 VP.t1 VSUBS 4.22006f
C102 VP.n53 VSUBS 1.54326f
C103 VP.n54 VSUBS 0.02669f
C104 VP.n55 VSUBS 0.036816f
C105 VP.n56 VSUBS 0.022807f
C106 VP.n57 VSUBS 0.022807f
C107 VP.n58 VSUBS 0.04272f
C108 VP.n59 VSUBS 0.042928f
C109 VP.n60 VSUBS 0.020417f
C110 VP.n61 VSUBS 0.022807f
C111 VP.n62 VSUBS 0.022807f
C112 VP.n63 VSUBS 0.022807f
C113 VP.n64 VSUBS 0.04272f
C114 VP.n65 VSUBS 0.041032f
C115 VP.n66 VSUBS 1.45441f
C116 VP.n67 VSUBS 0.023315f
C117 VP.n68 VSUBS 0.022807f
C118 VP.n69 VSUBS 0.022807f
C119 VP.n70 VSUBS 0.022807f
C120 VP.n71 VSUBS 0.04272f
C121 VP.n72 VSUBS 0.045571f
C122 VP.n73 VSUBS 0.018456f
C123 VP.n74 VSUBS 0.022807f
C124 VP.n75 VSUBS 0.022807f
C125 VP.n76 VSUBS 0.022807f
C126 VP.n77 VSUBS 0.04272f
C127 VP.n78 VSUBS 0.04272f
C128 VP.t6 VSUBS 4.22006f
C129 VP.n79 VSUBS 1.45441f
C130 VP.n80 VSUBS 0.023315f
C131 VP.n81 VSUBS 0.022807f
C132 VP.n82 VSUBS 0.022807f
C133 VP.n83 VSUBS 0.022807f
C134 VP.n84 VSUBS 0.04272f
C135 VP.n85 VSUBS 0.046252f
C136 VP.n86 VSUBS 0.020417f
C137 VP.n87 VSUBS 0.022807f
C138 VP.n88 VSUBS 0.022807f
C139 VP.n89 VSUBS 0.022807f
C140 VP.n90 VSUBS 0.04272f
C141 VP.n91 VSUBS 0.04272f
C142 VP.n92 VSUBS 0.02669f
C143 VP.n93 VSUBS 0.036816f
C144 VP.n94 VSUBS 0.067412f
C145 B.n0 VSUBS 0.004672f
C146 B.n1 VSUBS 0.004672f
C147 B.n2 VSUBS 0.007387f
C148 B.n3 VSUBS 0.007387f
C149 B.n4 VSUBS 0.007387f
C150 B.n5 VSUBS 0.007387f
C151 B.n6 VSUBS 0.007387f
C152 B.n7 VSUBS 0.007387f
C153 B.n8 VSUBS 0.007387f
C154 B.n9 VSUBS 0.007387f
C155 B.n10 VSUBS 0.007387f
C156 B.n11 VSUBS 0.007387f
C157 B.n12 VSUBS 0.007387f
C158 B.n13 VSUBS 0.007387f
C159 B.n14 VSUBS 0.007387f
C160 B.n15 VSUBS 0.007387f
C161 B.n16 VSUBS 0.007387f
C162 B.n17 VSUBS 0.007387f
C163 B.n18 VSUBS 0.007387f
C164 B.n19 VSUBS 0.007387f
C165 B.n20 VSUBS 0.007387f
C166 B.n21 VSUBS 0.007387f
C167 B.n22 VSUBS 0.007387f
C168 B.n23 VSUBS 0.007387f
C169 B.n24 VSUBS 0.007387f
C170 B.n25 VSUBS 0.007387f
C171 B.n26 VSUBS 0.007387f
C172 B.n27 VSUBS 0.007387f
C173 B.n28 VSUBS 0.007387f
C174 B.n29 VSUBS 0.007387f
C175 B.n30 VSUBS 0.007387f
C176 B.n31 VSUBS 0.007387f
C177 B.n32 VSUBS 0.007387f
C178 B.n33 VSUBS 0.007387f
C179 B.n34 VSUBS 0.007387f
C180 B.n35 VSUBS 0.007387f
C181 B.n36 VSUBS 0.017757f
C182 B.n37 VSUBS 0.007387f
C183 B.n38 VSUBS 0.007387f
C184 B.n39 VSUBS 0.007387f
C185 B.n40 VSUBS 0.007387f
C186 B.n41 VSUBS 0.007387f
C187 B.n42 VSUBS 0.007387f
C188 B.n43 VSUBS 0.007387f
C189 B.n44 VSUBS 0.007387f
C190 B.n45 VSUBS 0.007387f
C191 B.n46 VSUBS 0.007387f
C192 B.n47 VSUBS 0.007387f
C193 B.n48 VSUBS 0.007387f
C194 B.n49 VSUBS 0.007387f
C195 B.n50 VSUBS 0.007387f
C196 B.n51 VSUBS 0.007387f
C197 B.n52 VSUBS 0.007387f
C198 B.n53 VSUBS 0.007387f
C199 B.n54 VSUBS 0.007387f
C200 B.n55 VSUBS 0.007387f
C201 B.n56 VSUBS 0.007387f
C202 B.n57 VSUBS 0.007387f
C203 B.n58 VSUBS 0.007387f
C204 B.n59 VSUBS 0.007387f
C205 B.n60 VSUBS 0.007387f
C206 B.n61 VSUBS 0.007387f
C207 B.n62 VSUBS 0.007387f
C208 B.n63 VSUBS 0.007387f
C209 B.n64 VSUBS 0.007387f
C210 B.n65 VSUBS 0.007387f
C211 B.t5 VSUBS 0.639049f
C212 B.t4 VSUBS 0.668385f
C213 B.t3 VSUBS 3.23308f
C214 B.n66 VSUBS 0.41484f
C215 B.n67 VSUBS 0.081109f
C216 B.n68 VSUBS 0.007387f
C217 B.n69 VSUBS 0.007387f
C218 B.n70 VSUBS 0.007387f
C219 B.n71 VSUBS 0.007387f
C220 B.n72 VSUBS 0.004128f
C221 B.n73 VSUBS 0.007387f
C222 B.t8 VSUBS 0.639026f
C223 B.t7 VSUBS 0.668368f
C224 B.t6 VSUBS 3.23308f
C225 B.n74 VSUBS 0.414857f
C226 B.n75 VSUBS 0.081132f
C227 B.n76 VSUBS 0.017116f
C228 B.n77 VSUBS 0.007387f
C229 B.n78 VSUBS 0.007387f
C230 B.n79 VSUBS 0.007387f
C231 B.n80 VSUBS 0.007387f
C232 B.n81 VSUBS 0.007387f
C233 B.n82 VSUBS 0.007387f
C234 B.n83 VSUBS 0.007387f
C235 B.n84 VSUBS 0.007387f
C236 B.n85 VSUBS 0.007387f
C237 B.n86 VSUBS 0.007387f
C238 B.n87 VSUBS 0.007387f
C239 B.n88 VSUBS 0.007387f
C240 B.n89 VSUBS 0.007387f
C241 B.n90 VSUBS 0.007387f
C242 B.n91 VSUBS 0.007387f
C243 B.n92 VSUBS 0.007387f
C244 B.n93 VSUBS 0.007387f
C245 B.n94 VSUBS 0.007387f
C246 B.n95 VSUBS 0.007387f
C247 B.n96 VSUBS 0.007387f
C248 B.n97 VSUBS 0.007387f
C249 B.n98 VSUBS 0.007387f
C250 B.n99 VSUBS 0.007387f
C251 B.n100 VSUBS 0.007387f
C252 B.n101 VSUBS 0.007387f
C253 B.n102 VSUBS 0.007387f
C254 B.n103 VSUBS 0.007387f
C255 B.n104 VSUBS 0.007387f
C256 B.n105 VSUBS 0.017456f
C257 B.n106 VSUBS 0.007387f
C258 B.n107 VSUBS 0.007387f
C259 B.n108 VSUBS 0.007387f
C260 B.n109 VSUBS 0.007387f
C261 B.n110 VSUBS 0.007387f
C262 B.n111 VSUBS 0.007387f
C263 B.n112 VSUBS 0.007387f
C264 B.n113 VSUBS 0.007387f
C265 B.n114 VSUBS 0.007387f
C266 B.n115 VSUBS 0.007387f
C267 B.n116 VSUBS 0.007387f
C268 B.n117 VSUBS 0.007387f
C269 B.n118 VSUBS 0.007387f
C270 B.n119 VSUBS 0.007387f
C271 B.n120 VSUBS 0.007387f
C272 B.n121 VSUBS 0.007387f
C273 B.n122 VSUBS 0.007387f
C274 B.n123 VSUBS 0.007387f
C275 B.n124 VSUBS 0.007387f
C276 B.n125 VSUBS 0.007387f
C277 B.n126 VSUBS 0.007387f
C278 B.n127 VSUBS 0.007387f
C279 B.n128 VSUBS 0.007387f
C280 B.n129 VSUBS 0.007387f
C281 B.n130 VSUBS 0.007387f
C282 B.n131 VSUBS 0.007387f
C283 B.n132 VSUBS 0.007387f
C284 B.n133 VSUBS 0.007387f
C285 B.n134 VSUBS 0.007387f
C286 B.n135 VSUBS 0.007387f
C287 B.n136 VSUBS 0.007387f
C288 B.n137 VSUBS 0.007387f
C289 B.n138 VSUBS 0.007387f
C290 B.n139 VSUBS 0.007387f
C291 B.n140 VSUBS 0.007387f
C292 B.n141 VSUBS 0.007387f
C293 B.n142 VSUBS 0.007387f
C294 B.n143 VSUBS 0.007387f
C295 B.n144 VSUBS 0.007387f
C296 B.n145 VSUBS 0.007387f
C297 B.n146 VSUBS 0.007387f
C298 B.n147 VSUBS 0.007387f
C299 B.n148 VSUBS 0.007387f
C300 B.n149 VSUBS 0.007387f
C301 B.n150 VSUBS 0.007387f
C302 B.n151 VSUBS 0.007387f
C303 B.n152 VSUBS 0.007387f
C304 B.n153 VSUBS 0.007387f
C305 B.n154 VSUBS 0.007387f
C306 B.n155 VSUBS 0.007387f
C307 B.n156 VSUBS 0.007387f
C308 B.n157 VSUBS 0.007387f
C309 B.n158 VSUBS 0.007387f
C310 B.n159 VSUBS 0.007387f
C311 B.n160 VSUBS 0.007387f
C312 B.n161 VSUBS 0.007387f
C313 B.n162 VSUBS 0.007387f
C314 B.n163 VSUBS 0.007387f
C315 B.n164 VSUBS 0.007387f
C316 B.n165 VSUBS 0.007387f
C317 B.n166 VSUBS 0.007387f
C318 B.n167 VSUBS 0.007387f
C319 B.n168 VSUBS 0.007387f
C320 B.n169 VSUBS 0.007387f
C321 B.n170 VSUBS 0.007387f
C322 B.n171 VSUBS 0.007387f
C323 B.n172 VSUBS 0.007387f
C324 B.n173 VSUBS 0.016573f
C325 B.n174 VSUBS 0.007387f
C326 B.n175 VSUBS 0.007387f
C327 B.n176 VSUBS 0.007387f
C328 B.n177 VSUBS 0.007387f
C329 B.n178 VSUBS 0.007387f
C330 B.n179 VSUBS 0.007387f
C331 B.n180 VSUBS 0.007387f
C332 B.n181 VSUBS 0.007387f
C333 B.n182 VSUBS 0.007387f
C334 B.n183 VSUBS 0.007387f
C335 B.n184 VSUBS 0.007387f
C336 B.n185 VSUBS 0.007387f
C337 B.n186 VSUBS 0.007387f
C338 B.n187 VSUBS 0.007387f
C339 B.n188 VSUBS 0.007387f
C340 B.n189 VSUBS 0.007387f
C341 B.n190 VSUBS 0.007387f
C342 B.n191 VSUBS 0.007387f
C343 B.n192 VSUBS 0.007387f
C344 B.n193 VSUBS 0.007387f
C345 B.n194 VSUBS 0.007387f
C346 B.n195 VSUBS 0.007387f
C347 B.n196 VSUBS 0.007387f
C348 B.n197 VSUBS 0.007387f
C349 B.n198 VSUBS 0.007387f
C350 B.n199 VSUBS 0.007387f
C351 B.n200 VSUBS 0.007387f
C352 B.n201 VSUBS 0.007387f
C353 B.n202 VSUBS 0.007387f
C354 B.t1 VSUBS 0.639026f
C355 B.t2 VSUBS 0.668368f
C356 B.t0 VSUBS 3.23308f
C357 B.n203 VSUBS 0.414857f
C358 B.n204 VSUBS 0.081132f
C359 B.n205 VSUBS 0.017116f
C360 B.n206 VSUBS 0.007387f
C361 B.n207 VSUBS 0.007387f
C362 B.n208 VSUBS 0.007387f
C363 B.n209 VSUBS 0.007387f
C364 B.n210 VSUBS 0.007387f
C365 B.t10 VSUBS 0.639049f
C366 B.t11 VSUBS 0.668385f
C367 B.t9 VSUBS 3.23308f
C368 B.n211 VSUBS 0.41484f
C369 B.n212 VSUBS 0.081109f
C370 B.n213 VSUBS 0.007387f
C371 B.n214 VSUBS 0.007387f
C372 B.n215 VSUBS 0.007387f
C373 B.n216 VSUBS 0.007387f
C374 B.n217 VSUBS 0.007387f
C375 B.n218 VSUBS 0.007387f
C376 B.n219 VSUBS 0.007387f
C377 B.n220 VSUBS 0.007387f
C378 B.n221 VSUBS 0.007387f
C379 B.n222 VSUBS 0.007387f
C380 B.n223 VSUBS 0.007387f
C381 B.n224 VSUBS 0.007387f
C382 B.n225 VSUBS 0.007387f
C383 B.n226 VSUBS 0.007387f
C384 B.n227 VSUBS 0.007387f
C385 B.n228 VSUBS 0.007387f
C386 B.n229 VSUBS 0.007387f
C387 B.n230 VSUBS 0.007387f
C388 B.n231 VSUBS 0.007387f
C389 B.n232 VSUBS 0.007387f
C390 B.n233 VSUBS 0.007387f
C391 B.n234 VSUBS 0.007387f
C392 B.n235 VSUBS 0.007387f
C393 B.n236 VSUBS 0.007387f
C394 B.n237 VSUBS 0.007387f
C395 B.n238 VSUBS 0.007387f
C396 B.n239 VSUBS 0.007387f
C397 B.n240 VSUBS 0.007387f
C398 B.n241 VSUBS 0.007387f
C399 B.n242 VSUBS 0.016573f
C400 B.n243 VSUBS 0.007387f
C401 B.n244 VSUBS 0.007387f
C402 B.n245 VSUBS 0.007387f
C403 B.n246 VSUBS 0.007387f
C404 B.n247 VSUBS 0.007387f
C405 B.n248 VSUBS 0.007387f
C406 B.n249 VSUBS 0.007387f
C407 B.n250 VSUBS 0.007387f
C408 B.n251 VSUBS 0.007387f
C409 B.n252 VSUBS 0.007387f
C410 B.n253 VSUBS 0.007387f
C411 B.n254 VSUBS 0.007387f
C412 B.n255 VSUBS 0.007387f
C413 B.n256 VSUBS 0.007387f
C414 B.n257 VSUBS 0.007387f
C415 B.n258 VSUBS 0.007387f
C416 B.n259 VSUBS 0.007387f
C417 B.n260 VSUBS 0.007387f
C418 B.n261 VSUBS 0.007387f
C419 B.n262 VSUBS 0.007387f
C420 B.n263 VSUBS 0.007387f
C421 B.n264 VSUBS 0.007387f
C422 B.n265 VSUBS 0.007387f
C423 B.n266 VSUBS 0.007387f
C424 B.n267 VSUBS 0.007387f
C425 B.n268 VSUBS 0.007387f
C426 B.n269 VSUBS 0.007387f
C427 B.n270 VSUBS 0.007387f
C428 B.n271 VSUBS 0.007387f
C429 B.n272 VSUBS 0.007387f
C430 B.n273 VSUBS 0.007387f
C431 B.n274 VSUBS 0.007387f
C432 B.n275 VSUBS 0.007387f
C433 B.n276 VSUBS 0.007387f
C434 B.n277 VSUBS 0.007387f
C435 B.n278 VSUBS 0.007387f
C436 B.n279 VSUBS 0.007387f
C437 B.n280 VSUBS 0.007387f
C438 B.n281 VSUBS 0.007387f
C439 B.n282 VSUBS 0.007387f
C440 B.n283 VSUBS 0.007387f
C441 B.n284 VSUBS 0.007387f
C442 B.n285 VSUBS 0.007387f
C443 B.n286 VSUBS 0.007387f
C444 B.n287 VSUBS 0.007387f
C445 B.n288 VSUBS 0.007387f
C446 B.n289 VSUBS 0.007387f
C447 B.n290 VSUBS 0.007387f
C448 B.n291 VSUBS 0.007387f
C449 B.n292 VSUBS 0.007387f
C450 B.n293 VSUBS 0.007387f
C451 B.n294 VSUBS 0.007387f
C452 B.n295 VSUBS 0.007387f
C453 B.n296 VSUBS 0.007387f
C454 B.n297 VSUBS 0.007387f
C455 B.n298 VSUBS 0.007387f
C456 B.n299 VSUBS 0.007387f
C457 B.n300 VSUBS 0.007387f
C458 B.n301 VSUBS 0.007387f
C459 B.n302 VSUBS 0.007387f
C460 B.n303 VSUBS 0.007387f
C461 B.n304 VSUBS 0.007387f
C462 B.n305 VSUBS 0.007387f
C463 B.n306 VSUBS 0.007387f
C464 B.n307 VSUBS 0.007387f
C465 B.n308 VSUBS 0.007387f
C466 B.n309 VSUBS 0.007387f
C467 B.n310 VSUBS 0.007387f
C468 B.n311 VSUBS 0.007387f
C469 B.n312 VSUBS 0.007387f
C470 B.n313 VSUBS 0.007387f
C471 B.n314 VSUBS 0.007387f
C472 B.n315 VSUBS 0.007387f
C473 B.n316 VSUBS 0.007387f
C474 B.n317 VSUBS 0.007387f
C475 B.n318 VSUBS 0.007387f
C476 B.n319 VSUBS 0.007387f
C477 B.n320 VSUBS 0.007387f
C478 B.n321 VSUBS 0.007387f
C479 B.n322 VSUBS 0.007387f
C480 B.n323 VSUBS 0.007387f
C481 B.n324 VSUBS 0.007387f
C482 B.n325 VSUBS 0.007387f
C483 B.n326 VSUBS 0.007387f
C484 B.n327 VSUBS 0.007387f
C485 B.n328 VSUBS 0.007387f
C486 B.n329 VSUBS 0.007387f
C487 B.n330 VSUBS 0.007387f
C488 B.n331 VSUBS 0.007387f
C489 B.n332 VSUBS 0.007387f
C490 B.n333 VSUBS 0.007387f
C491 B.n334 VSUBS 0.007387f
C492 B.n335 VSUBS 0.007387f
C493 B.n336 VSUBS 0.007387f
C494 B.n337 VSUBS 0.007387f
C495 B.n338 VSUBS 0.007387f
C496 B.n339 VSUBS 0.007387f
C497 B.n340 VSUBS 0.007387f
C498 B.n341 VSUBS 0.007387f
C499 B.n342 VSUBS 0.007387f
C500 B.n343 VSUBS 0.007387f
C501 B.n344 VSUBS 0.007387f
C502 B.n345 VSUBS 0.007387f
C503 B.n346 VSUBS 0.007387f
C504 B.n347 VSUBS 0.007387f
C505 B.n348 VSUBS 0.007387f
C506 B.n349 VSUBS 0.007387f
C507 B.n350 VSUBS 0.007387f
C508 B.n351 VSUBS 0.007387f
C509 B.n352 VSUBS 0.007387f
C510 B.n353 VSUBS 0.007387f
C511 B.n354 VSUBS 0.007387f
C512 B.n355 VSUBS 0.007387f
C513 B.n356 VSUBS 0.007387f
C514 B.n357 VSUBS 0.007387f
C515 B.n358 VSUBS 0.007387f
C516 B.n359 VSUBS 0.007387f
C517 B.n360 VSUBS 0.007387f
C518 B.n361 VSUBS 0.007387f
C519 B.n362 VSUBS 0.007387f
C520 B.n363 VSUBS 0.007387f
C521 B.n364 VSUBS 0.007387f
C522 B.n365 VSUBS 0.007387f
C523 B.n366 VSUBS 0.007387f
C524 B.n367 VSUBS 0.007387f
C525 B.n368 VSUBS 0.007387f
C526 B.n369 VSUBS 0.007387f
C527 B.n370 VSUBS 0.007387f
C528 B.n371 VSUBS 0.007387f
C529 B.n372 VSUBS 0.007387f
C530 B.n373 VSUBS 0.007387f
C531 B.n374 VSUBS 0.007387f
C532 B.n375 VSUBS 0.016573f
C533 B.n376 VSUBS 0.017757f
C534 B.n377 VSUBS 0.017757f
C535 B.n378 VSUBS 0.007387f
C536 B.n379 VSUBS 0.007387f
C537 B.n380 VSUBS 0.007387f
C538 B.n381 VSUBS 0.007387f
C539 B.n382 VSUBS 0.007387f
C540 B.n383 VSUBS 0.007387f
C541 B.n384 VSUBS 0.007387f
C542 B.n385 VSUBS 0.007387f
C543 B.n386 VSUBS 0.007387f
C544 B.n387 VSUBS 0.007387f
C545 B.n388 VSUBS 0.007387f
C546 B.n389 VSUBS 0.007387f
C547 B.n390 VSUBS 0.007387f
C548 B.n391 VSUBS 0.007387f
C549 B.n392 VSUBS 0.007387f
C550 B.n393 VSUBS 0.007387f
C551 B.n394 VSUBS 0.007387f
C552 B.n395 VSUBS 0.007387f
C553 B.n396 VSUBS 0.007387f
C554 B.n397 VSUBS 0.007387f
C555 B.n398 VSUBS 0.007387f
C556 B.n399 VSUBS 0.007387f
C557 B.n400 VSUBS 0.007387f
C558 B.n401 VSUBS 0.007387f
C559 B.n402 VSUBS 0.007387f
C560 B.n403 VSUBS 0.007387f
C561 B.n404 VSUBS 0.007387f
C562 B.n405 VSUBS 0.007387f
C563 B.n406 VSUBS 0.007387f
C564 B.n407 VSUBS 0.007387f
C565 B.n408 VSUBS 0.007387f
C566 B.n409 VSUBS 0.007387f
C567 B.n410 VSUBS 0.007387f
C568 B.n411 VSUBS 0.007387f
C569 B.n412 VSUBS 0.007387f
C570 B.n413 VSUBS 0.007387f
C571 B.n414 VSUBS 0.007387f
C572 B.n415 VSUBS 0.007387f
C573 B.n416 VSUBS 0.007387f
C574 B.n417 VSUBS 0.007387f
C575 B.n418 VSUBS 0.007387f
C576 B.n419 VSUBS 0.007387f
C577 B.n420 VSUBS 0.007387f
C578 B.n421 VSUBS 0.007387f
C579 B.n422 VSUBS 0.007387f
C580 B.n423 VSUBS 0.007387f
C581 B.n424 VSUBS 0.007387f
C582 B.n425 VSUBS 0.007387f
C583 B.n426 VSUBS 0.007387f
C584 B.n427 VSUBS 0.007387f
C585 B.n428 VSUBS 0.007387f
C586 B.n429 VSUBS 0.007387f
C587 B.n430 VSUBS 0.007387f
C588 B.n431 VSUBS 0.007387f
C589 B.n432 VSUBS 0.007387f
C590 B.n433 VSUBS 0.007387f
C591 B.n434 VSUBS 0.007387f
C592 B.n435 VSUBS 0.007387f
C593 B.n436 VSUBS 0.007387f
C594 B.n437 VSUBS 0.007387f
C595 B.n438 VSUBS 0.007387f
C596 B.n439 VSUBS 0.007387f
C597 B.n440 VSUBS 0.007387f
C598 B.n441 VSUBS 0.007387f
C599 B.n442 VSUBS 0.007387f
C600 B.n443 VSUBS 0.007387f
C601 B.n444 VSUBS 0.007387f
C602 B.n445 VSUBS 0.007387f
C603 B.n446 VSUBS 0.007387f
C604 B.n447 VSUBS 0.007387f
C605 B.n448 VSUBS 0.007387f
C606 B.n449 VSUBS 0.007387f
C607 B.n450 VSUBS 0.007387f
C608 B.n451 VSUBS 0.007387f
C609 B.n452 VSUBS 0.007387f
C610 B.n453 VSUBS 0.007387f
C611 B.n454 VSUBS 0.007387f
C612 B.n455 VSUBS 0.007387f
C613 B.n456 VSUBS 0.007387f
C614 B.n457 VSUBS 0.007387f
C615 B.n458 VSUBS 0.007387f
C616 B.n459 VSUBS 0.007387f
C617 B.n460 VSUBS 0.007387f
C618 B.n461 VSUBS 0.007387f
C619 B.n462 VSUBS 0.007387f
C620 B.n463 VSUBS 0.007387f
C621 B.n464 VSUBS 0.006953f
C622 B.n465 VSUBS 0.017116f
C623 B.n466 VSUBS 0.004128f
C624 B.n467 VSUBS 0.007387f
C625 B.n468 VSUBS 0.007387f
C626 B.n469 VSUBS 0.007387f
C627 B.n470 VSUBS 0.007387f
C628 B.n471 VSUBS 0.007387f
C629 B.n472 VSUBS 0.007387f
C630 B.n473 VSUBS 0.007387f
C631 B.n474 VSUBS 0.007387f
C632 B.n475 VSUBS 0.007387f
C633 B.n476 VSUBS 0.007387f
C634 B.n477 VSUBS 0.007387f
C635 B.n478 VSUBS 0.007387f
C636 B.n479 VSUBS 0.004128f
C637 B.n480 VSUBS 0.007387f
C638 B.n481 VSUBS 0.007387f
C639 B.n482 VSUBS 0.006953f
C640 B.n483 VSUBS 0.007387f
C641 B.n484 VSUBS 0.007387f
C642 B.n485 VSUBS 0.007387f
C643 B.n486 VSUBS 0.007387f
C644 B.n487 VSUBS 0.007387f
C645 B.n488 VSUBS 0.007387f
C646 B.n489 VSUBS 0.007387f
C647 B.n490 VSUBS 0.007387f
C648 B.n491 VSUBS 0.007387f
C649 B.n492 VSUBS 0.007387f
C650 B.n493 VSUBS 0.007387f
C651 B.n494 VSUBS 0.007387f
C652 B.n495 VSUBS 0.007387f
C653 B.n496 VSUBS 0.007387f
C654 B.n497 VSUBS 0.007387f
C655 B.n498 VSUBS 0.007387f
C656 B.n499 VSUBS 0.007387f
C657 B.n500 VSUBS 0.007387f
C658 B.n501 VSUBS 0.007387f
C659 B.n502 VSUBS 0.007387f
C660 B.n503 VSUBS 0.007387f
C661 B.n504 VSUBS 0.007387f
C662 B.n505 VSUBS 0.007387f
C663 B.n506 VSUBS 0.007387f
C664 B.n507 VSUBS 0.007387f
C665 B.n508 VSUBS 0.007387f
C666 B.n509 VSUBS 0.007387f
C667 B.n510 VSUBS 0.007387f
C668 B.n511 VSUBS 0.007387f
C669 B.n512 VSUBS 0.007387f
C670 B.n513 VSUBS 0.007387f
C671 B.n514 VSUBS 0.007387f
C672 B.n515 VSUBS 0.007387f
C673 B.n516 VSUBS 0.007387f
C674 B.n517 VSUBS 0.007387f
C675 B.n518 VSUBS 0.007387f
C676 B.n519 VSUBS 0.007387f
C677 B.n520 VSUBS 0.007387f
C678 B.n521 VSUBS 0.007387f
C679 B.n522 VSUBS 0.007387f
C680 B.n523 VSUBS 0.007387f
C681 B.n524 VSUBS 0.007387f
C682 B.n525 VSUBS 0.007387f
C683 B.n526 VSUBS 0.007387f
C684 B.n527 VSUBS 0.007387f
C685 B.n528 VSUBS 0.007387f
C686 B.n529 VSUBS 0.007387f
C687 B.n530 VSUBS 0.007387f
C688 B.n531 VSUBS 0.007387f
C689 B.n532 VSUBS 0.007387f
C690 B.n533 VSUBS 0.007387f
C691 B.n534 VSUBS 0.007387f
C692 B.n535 VSUBS 0.007387f
C693 B.n536 VSUBS 0.007387f
C694 B.n537 VSUBS 0.007387f
C695 B.n538 VSUBS 0.007387f
C696 B.n539 VSUBS 0.007387f
C697 B.n540 VSUBS 0.007387f
C698 B.n541 VSUBS 0.007387f
C699 B.n542 VSUBS 0.007387f
C700 B.n543 VSUBS 0.007387f
C701 B.n544 VSUBS 0.007387f
C702 B.n545 VSUBS 0.007387f
C703 B.n546 VSUBS 0.007387f
C704 B.n547 VSUBS 0.007387f
C705 B.n548 VSUBS 0.007387f
C706 B.n549 VSUBS 0.007387f
C707 B.n550 VSUBS 0.007387f
C708 B.n551 VSUBS 0.007387f
C709 B.n552 VSUBS 0.007387f
C710 B.n553 VSUBS 0.007387f
C711 B.n554 VSUBS 0.007387f
C712 B.n555 VSUBS 0.007387f
C713 B.n556 VSUBS 0.007387f
C714 B.n557 VSUBS 0.007387f
C715 B.n558 VSUBS 0.007387f
C716 B.n559 VSUBS 0.007387f
C717 B.n560 VSUBS 0.007387f
C718 B.n561 VSUBS 0.007387f
C719 B.n562 VSUBS 0.007387f
C720 B.n563 VSUBS 0.007387f
C721 B.n564 VSUBS 0.007387f
C722 B.n565 VSUBS 0.007387f
C723 B.n566 VSUBS 0.007387f
C724 B.n567 VSUBS 0.007387f
C725 B.n568 VSUBS 0.017757f
C726 B.n569 VSUBS 0.017757f
C727 B.n570 VSUBS 0.016573f
C728 B.n571 VSUBS 0.007387f
C729 B.n572 VSUBS 0.007387f
C730 B.n573 VSUBS 0.007387f
C731 B.n574 VSUBS 0.007387f
C732 B.n575 VSUBS 0.007387f
C733 B.n576 VSUBS 0.007387f
C734 B.n577 VSUBS 0.007387f
C735 B.n578 VSUBS 0.007387f
C736 B.n579 VSUBS 0.007387f
C737 B.n580 VSUBS 0.007387f
C738 B.n581 VSUBS 0.007387f
C739 B.n582 VSUBS 0.007387f
C740 B.n583 VSUBS 0.007387f
C741 B.n584 VSUBS 0.007387f
C742 B.n585 VSUBS 0.007387f
C743 B.n586 VSUBS 0.007387f
C744 B.n587 VSUBS 0.007387f
C745 B.n588 VSUBS 0.007387f
C746 B.n589 VSUBS 0.007387f
C747 B.n590 VSUBS 0.007387f
C748 B.n591 VSUBS 0.007387f
C749 B.n592 VSUBS 0.007387f
C750 B.n593 VSUBS 0.007387f
C751 B.n594 VSUBS 0.007387f
C752 B.n595 VSUBS 0.007387f
C753 B.n596 VSUBS 0.007387f
C754 B.n597 VSUBS 0.007387f
C755 B.n598 VSUBS 0.007387f
C756 B.n599 VSUBS 0.007387f
C757 B.n600 VSUBS 0.007387f
C758 B.n601 VSUBS 0.007387f
C759 B.n602 VSUBS 0.007387f
C760 B.n603 VSUBS 0.007387f
C761 B.n604 VSUBS 0.007387f
C762 B.n605 VSUBS 0.007387f
C763 B.n606 VSUBS 0.007387f
C764 B.n607 VSUBS 0.007387f
C765 B.n608 VSUBS 0.007387f
C766 B.n609 VSUBS 0.007387f
C767 B.n610 VSUBS 0.007387f
C768 B.n611 VSUBS 0.007387f
C769 B.n612 VSUBS 0.007387f
C770 B.n613 VSUBS 0.007387f
C771 B.n614 VSUBS 0.007387f
C772 B.n615 VSUBS 0.007387f
C773 B.n616 VSUBS 0.007387f
C774 B.n617 VSUBS 0.007387f
C775 B.n618 VSUBS 0.007387f
C776 B.n619 VSUBS 0.007387f
C777 B.n620 VSUBS 0.007387f
C778 B.n621 VSUBS 0.007387f
C779 B.n622 VSUBS 0.007387f
C780 B.n623 VSUBS 0.007387f
C781 B.n624 VSUBS 0.007387f
C782 B.n625 VSUBS 0.007387f
C783 B.n626 VSUBS 0.007387f
C784 B.n627 VSUBS 0.007387f
C785 B.n628 VSUBS 0.007387f
C786 B.n629 VSUBS 0.007387f
C787 B.n630 VSUBS 0.007387f
C788 B.n631 VSUBS 0.007387f
C789 B.n632 VSUBS 0.007387f
C790 B.n633 VSUBS 0.007387f
C791 B.n634 VSUBS 0.007387f
C792 B.n635 VSUBS 0.007387f
C793 B.n636 VSUBS 0.007387f
C794 B.n637 VSUBS 0.007387f
C795 B.n638 VSUBS 0.007387f
C796 B.n639 VSUBS 0.007387f
C797 B.n640 VSUBS 0.007387f
C798 B.n641 VSUBS 0.007387f
C799 B.n642 VSUBS 0.007387f
C800 B.n643 VSUBS 0.007387f
C801 B.n644 VSUBS 0.007387f
C802 B.n645 VSUBS 0.007387f
C803 B.n646 VSUBS 0.007387f
C804 B.n647 VSUBS 0.007387f
C805 B.n648 VSUBS 0.007387f
C806 B.n649 VSUBS 0.007387f
C807 B.n650 VSUBS 0.007387f
C808 B.n651 VSUBS 0.007387f
C809 B.n652 VSUBS 0.007387f
C810 B.n653 VSUBS 0.007387f
C811 B.n654 VSUBS 0.007387f
C812 B.n655 VSUBS 0.007387f
C813 B.n656 VSUBS 0.007387f
C814 B.n657 VSUBS 0.007387f
C815 B.n658 VSUBS 0.007387f
C816 B.n659 VSUBS 0.007387f
C817 B.n660 VSUBS 0.007387f
C818 B.n661 VSUBS 0.007387f
C819 B.n662 VSUBS 0.007387f
C820 B.n663 VSUBS 0.007387f
C821 B.n664 VSUBS 0.007387f
C822 B.n665 VSUBS 0.007387f
C823 B.n666 VSUBS 0.007387f
C824 B.n667 VSUBS 0.007387f
C825 B.n668 VSUBS 0.007387f
C826 B.n669 VSUBS 0.007387f
C827 B.n670 VSUBS 0.007387f
C828 B.n671 VSUBS 0.007387f
C829 B.n672 VSUBS 0.007387f
C830 B.n673 VSUBS 0.007387f
C831 B.n674 VSUBS 0.007387f
C832 B.n675 VSUBS 0.007387f
C833 B.n676 VSUBS 0.007387f
C834 B.n677 VSUBS 0.007387f
C835 B.n678 VSUBS 0.007387f
C836 B.n679 VSUBS 0.007387f
C837 B.n680 VSUBS 0.007387f
C838 B.n681 VSUBS 0.007387f
C839 B.n682 VSUBS 0.007387f
C840 B.n683 VSUBS 0.007387f
C841 B.n684 VSUBS 0.007387f
C842 B.n685 VSUBS 0.007387f
C843 B.n686 VSUBS 0.007387f
C844 B.n687 VSUBS 0.007387f
C845 B.n688 VSUBS 0.007387f
C846 B.n689 VSUBS 0.007387f
C847 B.n690 VSUBS 0.007387f
C848 B.n691 VSUBS 0.007387f
C849 B.n692 VSUBS 0.007387f
C850 B.n693 VSUBS 0.007387f
C851 B.n694 VSUBS 0.007387f
C852 B.n695 VSUBS 0.007387f
C853 B.n696 VSUBS 0.007387f
C854 B.n697 VSUBS 0.007387f
C855 B.n698 VSUBS 0.007387f
C856 B.n699 VSUBS 0.007387f
C857 B.n700 VSUBS 0.007387f
C858 B.n701 VSUBS 0.007387f
C859 B.n702 VSUBS 0.007387f
C860 B.n703 VSUBS 0.007387f
C861 B.n704 VSUBS 0.007387f
C862 B.n705 VSUBS 0.007387f
C863 B.n706 VSUBS 0.007387f
C864 B.n707 VSUBS 0.007387f
C865 B.n708 VSUBS 0.007387f
C866 B.n709 VSUBS 0.007387f
C867 B.n710 VSUBS 0.007387f
C868 B.n711 VSUBS 0.007387f
C869 B.n712 VSUBS 0.007387f
C870 B.n713 VSUBS 0.007387f
C871 B.n714 VSUBS 0.007387f
C872 B.n715 VSUBS 0.007387f
C873 B.n716 VSUBS 0.007387f
C874 B.n717 VSUBS 0.007387f
C875 B.n718 VSUBS 0.007387f
C876 B.n719 VSUBS 0.007387f
C877 B.n720 VSUBS 0.007387f
C878 B.n721 VSUBS 0.007387f
C879 B.n722 VSUBS 0.007387f
C880 B.n723 VSUBS 0.007387f
C881 B.n724 VSUBS 0.007387f
C882 B.n725 VSUBS 0.007387f
C883 B.n726 VSUBS 0.007387f
C884 B.n727 VSUBS 0.007387f
C885 B.n728 VSUBS 0.007387f
C886 B.n729 VSUBS 0.007387f
C887 B.n730 VSUBS 0.007387f
C888 B.n731 VSUBS 0.007387f
C889 B.n732 VSUBS 0.007387f
C890 B.n733 VSUBS 0.007387f
C891 B.n734 VSUBS 0.007387f
C892 B.n735 VSUBS 0.007387f
C893 B.n736 VSUBS 0.007387f
C894 B.n737 VSUBS 0.007387f
C895 B.n738 VSUBS 0.007387f
C896 B.n739 VSUBS 0.007387f
C897 B.n740 VSUBS 0.007387f
C898 B.n741 VSUBS 0.007387f
C899 B.n742 VSUBS 0.007387f
C900 B.n743 VSUBS 0.007387f
C901 B.n744 VSUBS 0.007387f
C902 B.n745 VSUBS 0.007387f
C903 B.n746 VSUBS 0.007387f
C904 B.n747 VSUBS 0.007387f
C905 B.n748 VSUBS 0.007387f
C906 B.n749 VSUBS 0.007387f
C907 B.n750 VSUBS 0.007387f
C908 B.n751 VSUBS 0.007387f
C909 B.n752 VSUBS 0.007387f
C910 B.n753 VSUBS 0.007387f
C911 B.n754 VSUBS 0.007387f
C912 B.n755 VSUBS 0.007387f
C913 B.n756 VSUBS 0.007387f
C914 B.n757 VSUBS 0.007387f
C915 B.n758 VSUBS 0.007387f
C916 B.n759 VSUBS 0.007387f
C917 B.n760 VSUBS 0.007387f
C918 B.n761 VSUBS 0.007387f
C919 B.n762 VSUBS 0.007387f
C920 B.n763 VSUBS 0.007387f
C921 B.n764 VSUBS 0.007387f
C922 B.n765 VSUBS 0.007387f
C923 B.n766 VSUBS 0.007387f
C924 B.n767 VSUBS 0.007387f
C925 B.n768 VSUBS 0.007387f
C926 B.n769 VSUBS 0.007387f
C927 B.n770 VSUBS 0.007387f
C928 B.n771 VSUBS 0.007387f
C929 B.n772 VSUBS 0.007387f
C930 B.n773 VSUBS 0.007387f
C931 B.n774 VSUBS 0.016573f
C932 B.n775 VSUBS 0.017757f
C933 B.n776 VSUBS 0.016875f
C934 B.n777 VSUBS 0.007387f
C935 B.n778 VSUBS 0.007387f
C936 B.n779 VSUBS 0.007387f
C937 B.n780 VSUBS 0.007387f
C938 B.n781 VSUBS 0.007387f
C939 B.n782 VSUBS 0.007387f
C940 B.n783 VSUBS 0.007387f
C941 B.n784 VSUBS 0.007387f
C942 B.n785 VSUBS 0.007387f
C943 B.n786 VSUBS 0.007387f
C944 B.n787 VSUBS 0.007387f
C945 B.n788 VSUBS 0.007387f
C946 B.n789 VSUBS 0.007387f
C947 B.n790 VSUBS 0.007387f
C948 B.n791 VSUBS 0.007387f
C949 B.n792 VSUBS 0.007387f
C950 B.n793 VSUBS 0.007387f
C951 B.n794 VSUBS 0.007387f
C952 B.n795 VSUBS 0.007387f
C953 B.n796 VSUBS 0.007387f
C954 B.n797 VSUBS 0.007387f
C955 B.n798 VSUBS 0.007387f
C956 B.n799 VSUBS 0.007387f
C957 B.n800 VSUBS 0.007387f
C958 B.n801 VSUBS 0.007387f
C959 B.n802 VSUBS 0.007387f
C960 B.n803 VSUBS 0.007387f
C961 B.n804 VSUBS 0.007387f
C962 B.n805 VSUBS 0.007387f
C963 B.n806 VSUBS 0.007387f
C964 B.n807 VSUBS 0.007387f
C965 B.n808 VSUBS 0.007387f
C966 B.n809 VSUBS 0.007387f
C967 B.n810 VSUBS 0.007387f
C968 B.n811 VSUBS 0.007387f
C969 B.n812 VSUBS 0.007387f
C970 B.n813 VSUBS 0.007387f
C971 B.n814 VSUBS 0.007387f
C972 B.n815 VSUBS 0.007387f
C973 B.n816 VSUBS 0.007387f
C974 B.n817 VSUBS 0.007387f
C975 B.n818 VSUBS 0.007387f
C976 B.n819 VSUBS 0.007387f
C977 B.n820 VSUBS 0.007387f
C978 B.n821 VSUBS 0.007387f
C979 B.n822 VSUBS 0.007387f
C980 B.n823 VSUBS 0.007387f
C981 B.n824 VSUBS 0.007387f
C982 B.n825 VSUBS 0.007387f
C983 B.n826 VSUBS 0.007387f
C984 B.n827 VSUBS 0.007387f
C985 B.n828 VSUBS 0.007387f
C986 B.n829 VSUBS 0.007387f
C987 B.n830 VSUBS 0.007387f
C988 B.n831 VSUBS 0.007387f
C989 B.n832 VSUBS 0.007387f
C990 B.n833 VSUBS 0.007387f
C991 B.n834 VSUBS 0.007387f
C992 B.n835 VSUBS 0.007387f
C993 B.n836 VSUBS 0.007387f
C994 B.n837 VSUBS 0.007387f
C995 B.n838 VSUBS 0.007387f
C996 B.n839 VSUBS 0.007387f
C997 B.n840 VSUBS 0.007387f
C998 B.n841 VSUBS 0.007387f
C999 B.n842 VSUBS 0.007387f
C1000 B.n843 VSUBS 0.007387f
C1001 B.n844 VSUBS 0.007387f
C1002 B.n845 VSUBS 0.007387f
C1003 B.n846 VSUBS 0.007387f
C1004 B.n847 VSUBS 0.007387f
C1005 B.n848 VSUBS 0.007387f
C1006 B.n849 VSUBS 0.007387f
C1007 B.n850 VSUBS 0.007387f
C1008 B.n851 VSUBS 0.007387f
C1009 B.n852 VSUBS 0.007387f
C1010 B.n853 VSUBS 0.007387f
C1011 B.n854 VSUBS 0.007387f
C1012 B.n855 VSUBS 0.007387f
C1013 B.n856 VSUBS 0.007387f
C1014 B.n857 VSUBS 0.007387f
C1015 B.n858 VSUBS 0.007387f
C1016 B.n859 VSUBS 0.007387f
C1017 B.n860 VSUBS 0.007387f
C1018 B.n861 VSUBS 0.007387f
C1019 B.n862 VSUBS 0.006953f
C1020 B.n863 VSUBS 0.007387f
C1021 B.n864 VSUBS 0.007387f
C1022 B.n865 VSUBS 0.007387f
C1023 B.n866 VSUBS 0.007387f
C1024 B.n867 VSUBS 0.007387f
C1025 B.n868 VSUBS 0.007387f
C1026 B.n869 VSUBS 0.007387f
C1027 B.n870 VSUBS 0.007387f
C1028 B.n871 VSUBS 0.007387f
C1029 B.n872 VSUBS 0.007387f
C1030 B.n873 VSUBS 0.007387f
C1031 B.n874 VSUBS 0.007387f
C1032 B.n875 VSUBS 0.007387f
C1033 B.n876 VSUBS 0.007387f
C1034 B.n877 VSUBS 0.007387f
C1035 B.n878 VSUBS 0.004128f
C1036 B.n879 VSUBS 0.017116f
C1037 B.n880 VSUBS 0.006953f
C1038 B.n881 VSUBS 0.007387f
C1039 B.n882 VSUBS 0.007387f
C1040 B.n883 VSUBS 0.007387f
C1041 B.n884 VSUBS 0.007387f
C1042 B.n885 VSUBS 0.007387f
C1043 B.n886 VSUBS 0.007387f
C1044 B.n887 VSUBS 0.007387f
C1045 B.n888 VSUBS 0.007387f
C1046 B.n889 VSUBS 0.007387f
C1047 B.n890 VSUBS 0.007387f
C1048 B.n891 VSUBS 0.007387f
C1049 B.n892 VSUBS 0.007387f
C1050 B.n893 VSUBS 0.007387f
C1051 B.n894 VSUBS 0.007387f
C1052 B.n895 VSUBS 0.007387f
C1053 B.n896 VSUBS 0.007387f
C1054 B.n897 VSUBS 0.007387f
C1055 B.n898 VSUBS 0.007387f
C1056 B.n899 VSUBS 0.007387f
C1057 B.n900 VSUBS 0.007387f
C1058 B.n901 VSUBS 0.007387f
C1059 B.n902 VSUBS 0.007387f
C1060 B.n903 VSUBS 0.007387f
C1061 B.n904 VSUBS 0.007387f
C1062 B.n905 VSUBS 0.007387f
C1063 B.n906 VSUBS 0.007387f
C1064 B.n907 VSUBS 0.007387f
C1065 B.n908 VSUBS 0.007387f
C1066 B.n909 VSUBS 0.007387f
C1067 B.n910 VSUBS 0.007387f
C1068 B.n911 VSUBS 0.007387f
C1069 B.n912 VSUBS 0.007387f
C1070 B.n913 VSUBS 0.007387f
C1071 B.n914 VSUBS 0.007387f
C1072 B.n915 VSUBS 0.007387f
C1073 B.n916 VSUBS 0.007387f
C1074 B.n917 VSUBS 0.007387f
C1075 B.n918 VSUBS 0.007387f
C1076 B.n919 VSUBS 0.007387f
C1077 B.n920 VSUBS 0.007387f
C1078 B.n921 VSUBS 0.007387f
C1079 B.n922 VSUBS 0.007387f
C1080 B.n923 VSUBS 0.007387f
C1081 B.n924 VSUBS 0.007387f
C1082 B.n925 VSUBS 0.007387f
C1083 B.n926 VSUBS 0.007387f
C1084 B.n927 VSUBS 0.007387f
C1085 B.n928 VSUBS 0.007387f
C1086 B.n929 VSUBS 0.007387f
C1087 B.n930 VSUBS 0.007387f
C1088 B.n931 VSUBS 0.007387f
C1089 B.n932 VSUBS 0.007387f
C1090 B.n933 VSUBS 0.007387f
C1091 B.n934 VSUBS 0.007387f
C1092 B.n935 VSUBS 0.007387f
C1093 B.n936 VSUBS 0.007387f
C1094 B.n937 VSUBS 0.007387f
C1095 B.n938 VSUBS 0.007387f
C1096 B.n939 VSUBS 0.007387f
C1097 B.n940 VSUBS 0.007387f
C1098 B.n941 VSUBS 0.007387f
C1099 B.n942 VSUBS 0.007387f
C1100 B.n943 VSUBS 0.007387f
C1101 B.n944 VSUBS 0.007387f
C1102 B.n945 VSUBS 0.007387f
C1103 B.n946 VSUBS 0.007387f
C1104 B.n947 VSUBS 0.007387f
C1105 B.n948 VSUBS 0.007387f
C1106 B.n949 VSUBS 0.007387f
C1107 B.n950 VSUBS 0.007387f
C1108 B.n951 VSUBS 0.007387f
C1109 B.n952 VSUBS 0.007387f
C1110 B.n953 VSUBS 0.007387f
C1111 B.n954 VSUBS 0.007387f
C1112 B.n955 VSUBS 0.007387f
C1113 B.n956 VSUBS 0.007387f
C1114 B.n957 VSUBS 0.007387f
C1115 B.n958 VSUBS 0.007387f
C1116 B.n959 VSUBS 0.007387f
C1117 B.n960 VSUBS 0.007387f
C1118 B.n961 VSUBS 0.007387f
C1119 B.n962 VSUBS 0.007387f
C1120 B.n963 VSUBS 0.007387f
C1121 B.n964 VSUBS 0.007387f
C1122 B.n965 VSUBS 0.007387f
C1123 B.n966 VSUBS 0.007387f
C1124 B.n967 VSUBS 0.017757f
C1125 B.n968 VSUBS 0.016573f
C1126 B.n969 VSUBS 0.016573f
C1127 B.n970 VSUBS 0.007387f
C1128 B.n971 VSUBS 0.007387f
C1129 B.n972 VSUBS 0.007387f
C1130 B.n973 VSUBS 0.007387f
C1131 B.n974 VSUBS 0.007387f
C1132 B.n975 VSUBS 0.007387f
C1133 B.n976 VSUBS 0.007387f
C1134 B.n977 VSUBS 0.007387f
C1135 B.n978 VSUBS 0.007387f
C1136 B.n979 VSUBS 0.007387f
C1137 B.n980 VSUBS 0.007387f
C1138 B.n981 VSUBS 0.007387f
C1139 B.n982 VSUBS 0.007387f
C1140 B.n983 VSUBS 0.007387f
C1141 B.n984 VSUBS 0.007387f
C1142 B.n985 VSUBS 0.007387f
C1143 B.n986 VSUBS 0.007387f
C1144 B.n987 VSUBS 0.007387f
C1145 B.n988 VSUBS 0.007387f
C1146 B.n989 VSUBS 0.007387f
C1147 B.n990 VSUBS 0.007387f
C1148 B.n991 VSUBS 0.007387f
C1149 B.n992 VSUBS 0.007387f
C1150 B.n993 VSUBS 0.007387f
C1151 B.n994 VSUBS 0.007387f
C1152 B.n995 VSUBS 0.007387f
C1153 B.n996 VSUBS 0.007387f
C1154 B.n997 VSUBS 0.007387f
C1155 B.n998 VSUBS 0.007387f
C1156 B.n999 VSUBS 0.007387f
C1157 B.n1000 VSUBS 0.007387f
C1158 B.n1001 VSUBS 0.007387f
C1159 B.n1002 VSUBS 0.007387f
C1160 B.n1003 VSUBS 0.007387f
C1161 B.n1004 VSUBS 0.007387f
C1162 B.n1005 VSUBS 0.007387f
C1163 B.n1006 VSUBS 0.007387f
C1164 B.n1007 VSUBS 0.007387f
C1165 B.n1008 VSUBS 0.007387f
C1166 B.n1009 VSUBS 0.007387f
C1167 B.n1010 VSUBS 0.007387f
C1168 B.n1011 VSUBS 0.007387f
C1169 B.n1012 VSUBS 0.007387f
C1170 B.n1013 VSUBS 0.007387f
C1171 B.n1014 VSUBS 0.007387f
C1172 B.n1015 VSUBS 0.007387f
C1173 B.n1016 VSUBS 0.007387f
C1174 B.n1017 VSUBS 0.007387f
C1175 B.n1018 VSUBS 0.007387f
C1176 B.n1019 VSUBS 0.007387f
C1177 B.n1020 VSUBS 0.007387f
C1178 B.n1021 VSUBS 0.007387f
C1179 B.n1022 VSUBS 0.007387f
C1180 B.n1023 VSUBS 0.007387f
C1181 B.n1024 VSUBS 0.007387f
C1182 B.n1025 VSUBS 0.007387f
C1183 B.n1026 VSUBS 0.007387f
C1184 B.n1027 VSUBS 0.007387f
C1185 B.n1028 VSUBS 0.007387f
C1186 B.n1029 VSUBS 0.007387f
C1187 B.n1030 VSUBS 0.007387f
C1188 B.n1031 VSUBS 0.007387f
C1189 B.n1032 VSUBS 0.007387f
C1190 B.n1033 VSUBS 0.007387f
C1191 B.n1034 VSUBS 0.007387f
C1192 B.n1035 VSUBS 0.007387f
C1193 B.n1036 VSUBS 0.007387f
C1194 B.n1037 VSUBS 0.007387f
C1195 B.n1038 VSUBS 0.007387f
C1196 B.n1039 VSUBS 0.007387f
C1197 B.n1040 VSUBS 0.007387f
C1198 B.n1041 VSUBS 0.007387f
C1199 B.n1042 VSUBS 0.007387f
C1200 B.n1043 VSUBS 0.007387f
C1201 B.n1044 VSUBS 0.007387f
C1202 B.n1045 VSUBS 0.007387f
C1203 B.n1046 VSUBS 0.007387f
C1204 B.n1047 VSUBS 0.007387f
C1205 B.n1048 VSUBS 0.007387f
C1206 B.n1049 VSUBS 0.007387f
C1207 B.n1050 VSUBS 0.007387f
C1208 B.n1051 VSUBS 0.007387f
C1209 B.n1052 VSUBS 0.007387f
C1210 B.n1053 VSUBS 0.007387f
C1211 B.n1054 VSUBS 0.007387f
C1212 B.n1055 VSUBS 0.007387f
C1213 B.n1056 VSUBS 0.007387f
C1214 B.n1057 VSUBS 0.007387f
C1215 B.n1058 VSUBS 0.007387f
C1216 B.n1059 VSUBS 0.007387f
C1217 B.n1060 VSUBS 0.007387f
C1218 B.n1061 VSUBS 0.007387f
C1219 B.n1062 VSUBS 0.007387f
C1220 B.n1063 VSUBS 0.007387f
C1221 B.n1064 VSUBS 0.007387f
C1222 B.n1065 VSUBS 0.007387f
C1223 B.n1066 VSUBS 0.007387f
C1224 B.n1067 VSUBS 0.007387f
C1225 B.n1068 VSUBS 0.007387f
C1226 B.n1069 VSUBS 0.007387f
C1227 B.n1070 VSUBS 0.007387f
C1228 B.n1071 VSUBS 0.016728f
C1229 VTAIL.t9 VSUBS 0.34465f
C1230 VTAIL.t11 VSUBS 0.34465f
C1231 VTAIL.n0 VSUBS 2.71921f
C1232 VTAIL.n1 VSUBS 0.869079f
C1233 VTAIL.t15 VSUBS 3.55027f
C1234 VTAIL.n2 VSUBS 1.01022f
C1235 VTAIL.t6 VSUBS 3.55027f
C1236 VTAIL.n3 VSUBS 1.01022f
C1237 VTAIL.t4 VSUBS 0.34465f
C1238 VTAIL.t1 VSUBS 0.34465f
C1239 VTAIL.n4 VSUBS 2.71921f
C1240 VTAIL.n5 VSUBS 1.14004f
C1241 VTAIL.t7 VSUBS 3.55027f
C1242 VTAIL.n6 VSUBS 2.79068f
C1243 VTAIL.t12 VSUBS 3.55027f
C1244 VTAIL.n7 VSUBS 2.79067f
C1245 VTAIL.t14 VSUBS 0.34465f
C1246 VTAIL.t8 VSUBS 0.34465f
C1247 VTAIL.n8 VSUBS 2.71922f
C1248 VTAIL.n9 VSUBS 1.14004f
C1249 VTAIL.t13 VSUBS 3.55027f
C1250 VTAIL.n10 VSUBS 1.01022f
C1251 VTAIL.t0 VSUBS 3.55027f
C1252 VTAIL.n11 VSUBS 1.01022f
C1253 VTAIL.t5 VSUBS 0.34465f
C1254 VTAIL.t3 VSUBS 0.34465f
C1255 VTAIL.n12 VSUBS 2.71922f
C1256 VTAIL.n13 VSUBS 1.14004f
C1257 VTAIL.t2 VSUBS 3.55027f
C1258 VTAIL.n14 VSUBS 2.79068f
C1259 VTAIL.t10 VSUBS 3.55027f
C1260 VTAIL.n15 VSUBS 2.78612f
C1261 VDD2.t3 VSUBS 0.445411f
C1262 VDD2.t7 VSUBS 0.445411f
C1263 VDD2.n0 VSUBS 3.73172f
C1264 VDD2.t1 VSUBS 0.445411f
C1265 VDD2.t0 VSUBS 0.445411f
C1266 VDD2.n1 VSUBS 3.73172f
C1267 VDD2.n2 VSUBS 6.12837f
C1268 VDD2.t4 VSUBS 0.445411f
C1269 VDD2.t2 VSUBS 0.445411f
C1270 VDD2.n3 VSUBS 3.70429f
C1271 VDD2.n4 VSUBS 5.12555f
C1272 VDD2.t6 VSUBS 0.445411f
C1273 VDD2.t5 VSUBS 0.445411f
C1274 VDD2.n5 VSUBS 3.73165f
C1275 VN.t5 VSUBS 3.90419f
C1276 VN.n0 VSUBS 1.42775f
C1277 VN.n1 VSUBS 0.0211f
C1278 VN.n2 VSUBS 0.039715f
C1279 VN.n3 VSUBS 0.0211f
C1280 VN.n4 VSUBS 0.037961f
C1281 VN.n5 VSUBS 0.0211f
C1282 VN.n6 VSUBS 0.04216f
C1283 VN.n7 VSUBS 0.0211f
C1284 VN.n8 VSUBS 0.039522f
C1285 VN.t0 VSUBS 4.23614f
C1286 VN.n9 VSUBS 1.35171f
C1287 VN.t6 VSUBS 3.90419f
C1288 VN.n10 VSUBS 1.41376f
C1289 VN.n11 VSUBS 0.02157f
C1290 VN.n12 VSUBS 0.268866f
C1291 VN.n13 VSUBS 0.0211f
C1292 VN.n14 VSUBS 0.0211f
C1293 VN.n15 VSUBS 0.039522f
C1294 VN.n16 VSUBS 0.04216f
C1295 VN.n17 VSUBS 0.017074f
C1296 VN.n18 VSUBS 0.0211f
C1297 VN.n19 VSUBS 0.0211f
C1298 VN.n20 VSUBS 0.0211f
C1299 VN.n21 VSUBS 0.039522f
C1300 VN.n22 VSUBS 0.039522f
C1301 VN.t4 VSUBS 3.90419f
C1302 VN.n23 VSUBS 1.34555f
C1303 VN.n24 VSUBS 0.02157f
C1304 VN.n25 VSUBS 0.0211f
C1305 VN.n26 VSUBS 0.0211f
C1306 VN.n27 VSUBS 0.0211f
C1307 VN.n28 VSUBS 0.039522f
C1308 VN.n29 VSUBS 0.04279f
C1309 VN.n30 VSUBS 0.018889f
C1310 VN.n31 VSUBS 0.0211f
C1311 VN.n32 VSUBS 0.0211f
C1312 VN.n33 VSUBS 0.0211f
C1313 VN.n34 VSUBS 0.039522f
C1314 VN.n35 VSUBS 0.039522f
C1315 VN.n36 VSUBS 0.024692f
C1316 VN.n37 VSUBS 0.03406f
C1317 VN.n38 VSUBS 0.062366f
C1318 VN.t3 VSUBS 3.90419f
C1319 VN.n39 VSUBS 1.42775f
C1320 VN.n40 VSUBS 0.0211f
C1321 VN.n41 VSUBS 0.039715f
C1322 VN.n42 VSUBS 0.0211f
C1323 VN.n43 VSUBS 0.037961f
C1324 VN.n44 VSUBS 0.0211f
C1325 VN.t1 VSUBS 3.90419f
C1326 VN.n45 VSUBS 1.34555f
C1327 VN.n46 VSUBS 0.04216f
C1328 VN.n47 VSUBS 0.0211f
C1329 VN.n48 VSUBS 0.039522f
C1330 VN.t2 VSUBS 4.23614f
C1331 VN.n49 VSUBS 1.35171f
C1332 VN.t7 VSUBS 3.90419f
C1333 VN.n50 VSUBS 1.41376f
C1334 VN.n51 VSUBS 0.02157f
C1335 VN.n52 VSUBS 0.268866f
C1336 VN.n53 VSUBS 0.0211f
C1337 VN.n54 VSUBS 0.0211f
C1338 VN.n55 VSUBS 0.039522f
C1339 VN.n56 VSUBS 0.04216f
C1340 VN.n57 VSUBS 0.017074f
C1341 VN.n58 VSUBS 0.0211f
C1342 VN.n59 VSUBS 0.0211f
C1343 VN.n60 VSUBS 0.0211f
C1344 VN.n61 VSUBS 0.039522f
C1345 VN.n62 VSUBS 0.039522f
C1346 VN.n63 VSUBS 0.02157f
C1347 VN.n64 VSUBS 0.0211f
C1348 VN.n65 VSUBS 0.0211f
C1349 VN.n66 VSUBS 0.0211f
C1350 VN.n67 VSUBS 0.039522f
C1351 VN.n68 VSUBS 0.04279f
C1352 VN.n69 VSUBS 0.018889f
C1353 VN.n70 VSUBS 0.0211f
C1354 VN.n71 VSUBS 0.0211f
C1355 VN.n72 VSUBS 0.0211f
C1356 VN.n73 VSUBS 0.039522f
C1357 VN.n74 VSUBS 0.039522f
C1358 VN.n75 VSUBS 0.024692f
C1359 VN.n76 VSUBS 0.03406f
C1360 VN.n77 VSUBS 1.59494f
.ends

