* NGSPICE file created from diff_pair_sample_0236.ext - technology: sky130A

.subckt diff_pair_sample_0236 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t11 VN.t0 VDD2.t3 w_n1730_n2028# sky130_fd_pr__pfet_01v8 ad=0.8745 pd=5.63 as=0.8745 ps=5.63 w=5.3 l=0.62
X1 VDD1.t5 VP.t0 VTAIL.t5 w_n1730_n2028# sky130_fd_pr__pfet_01v8 ad=2.067 pd=11.38 as=0.8745 ps=5.63 w=5.3 l=0.62
X2 VDD2.t0 VN.t1 VTAIL.t10 w_n1730_n2028# sky130_fd_pr__pfet_01v8 ad=2.067 pd=11.38 as=0.8745 ps=5.63 w=5.3 l=0.62
X3 VDD2.t2 VN.t2 VTAIL.t9 w_n1730_n2028# sky130_fd_pr__pfet_01v8 ad=0.8745 pd=5.63 as=2.067 ps=11.38 w=5.3 l=0.62
X4 B.t11 B.t9 B.t10 w_n1730_n2028# sky130_fd_pr__pfet_01v8 ad=2.067 pd=11.38 as=0 ps=0 w=5.3 l=0.62
X5 VTAIL.t8 VN.t3 VDD2.t1 w_n1730_n2028# sky130_fd_pr__pfet_01v8 ad=0.8745 pd=5.63 as=0.8745 ps=5.63 w=5.3 l=0.62
X6 VDD2.t4 VN.t4 VTAIL.t7 w_n1730_n2028# sky130_fd_pr__pfet_01v8 ad=0.8745 pd=5.63 as=2.067 ps=11.38 w=5.3 l=0.62
X7 VDD1.t4 VP.t1 VTAIL.t2 w_n1730_n2028# sky130_fd_pr__pfet_01v8 ad=0.8745 pd=5.63 as=2.067 ps=11.38 w=5.3 l=0.62
X8 B.t8 B.t6 B.t7 w_n1730_n2028# sky130_fd_pr__pfet_01v8 ad=2.067 pd=11.38 as=0 ps=0 w=5.3 l=0.62
X9 VDD2.t5 VN.t5 VTAIL.t6 w_n1730_n2028# sky130_fd_pr__pfet_01v8 ad=2.067 pd=11.38 as=0.8745 ps=5.63 w=5.3 l=0.62
X10 VDD1.t3 VP.t2 VTAIL.t4 w_n1730_n2028# sky130_fd_pr__pfet_01v8 ad=0.8745 pd=5.63 as=2.067 ps=11.38 w=5.3 l=0.62
X11 VTAIL.t3 VP.t3 VDD1.t2 w_n1730_n2028# sky130_fd_pr__pfet_01v8 ad=0.8745 pd=5.63 as=0.8745 ps=5.63 w=5.3 l=0.62
X12 VTAIL.t0 VP.t4 VDD1.t1 w_n1730_n2028# sky130_fd_pr__pfet_01v8 ad=0.8745 pd=5.63 as=0.8745 ps=5.63 w=5.3 l=0.62
X13 B.t5 B.t3 B.t4 w_n1730_n2028# sky130_fd_pr__pfet_01v8 ad=2.067 pd=11.38 as=0 ps=0 w=5.3 l=0.62
X14 VDD1.t0 VP.t5 VTAIL.t1 w_n1730_n2028# sky130_fd_pr__pfet_01v8 ad=2.067 pd=11.38 as=0.8745 ps=5.63 w=5.3 l=0.62
X15 B.t2 B.t0 B.t1 w_n1730_n2028# sky130_fd_pr__pfet_01v8 ad=2.067 pd=11.38 as=0 ps=0 w=5.3 l=0.62
R0 VN.n0 VN.t1 296.197
R1 VN.n4 VN.t2 296.197
R2 VN.n1 VN.t3 269.377
R3 VN.n2 VN.t4 269.377
R4 VN.n5 VN.t0 269.377
R5 VN.n6 VN.t5 269.377
R6 VN.n3 VN.n2 161.3
R7 VN.n7 VN.n6 161.3
R8 VN.n2 VN.n1 48.2005
R9 VN.n6 VN.n5 48.2005
R10 VN.n7 VN.n4 45.1367
R11 VN.n3 VN.n0 45.1367
R12 VN VN.n7 36.3016
R13 VN.n5 VN.n4 13.3799
R14 VN.n1 VN.n0 13.3799
R15 VN VN.n3 0.0516364
R16 VDD2.n51 VDD2.n29 756.745
R17 VDD2.n22 VDD2.n0 756.745
R18 VDD2.n52 VDD2.n51 585
R19 VDD2.n50 VDD2.n49 585
R20 VDD2.n33 VDD2.n32 585
R21 VDD2.n44 VDD2.n43 585
R22 VDD2.n42 VDD2.n41 585
R23 VDD2.n37 VDD2.n36 585
R24 VDD2.n8 VDD2.n7 585
R25 VDD2.n13 VDD2.n12 585
R26 VDD2.n15 VDD2.n14 585
R27 VDD2.n4 VDD2.n3 585
R28 VDD2.n21 VDD2.n20 585
R29 VDD2.n23 VDD2.n22 585
R30 VDD2.n38 VDD2.t5 327.856
R31 VDD2.n9 VDD2.t0 327.856
R32 VDD2.n51 VDD2.n50 171.744
R33 VDD2.n50 VDD2.n32 171.744
R34 VDD2.n43 VDD2.n32 171.744
R35 VDD2.n43 VDD2.n42 171.744
R36 VDD2.n42 VDD2.n36 171.744
R37 VDD2.n13 VDD2.n7 171.744
R38 VDD2.n14 VDD2.n13 171.744
R39 VDD2.n14 VDD2.n3 171.744
R40 VDD2.n21 VDD2.n3 171.744
R41 VDD2.n22 VDD2.n21 171.744
R42 VDD2.n28 VDD2.n27 97.868
R43 VDD2 VDD2.n57 97.8652
R44 VDD2.t5 VDD2.n36 85.8723
R45 VDD2.t0 VDD2.n7 85.8723
R46 VDD2.n28 VDD2.n26 49.8109
R47 VDD2.n56 VDD2.n55 49.252
R48 VDD2.n56 VDD2.n28 30.9459
R49 VDD2.n38 VDD2.n37 16.381
R50 VDD2.n9 VDD2.n8 16.381
R51 VDD2.n41 VDD2.n40 12.8005
R52 VDD2.n12 VDD2.n11 12.8005
R53 VDD2.n44 VDD2.n35 12.0247
R54 VDD2.n15 VDD2.n6 12.0247
R55 VDD2.n45 VDD2.n33 11.249
R56 VDD2.n16 VDD2.n4 11.249
R57 VDD2.n49 VDD2.n48 10.4732
R58 VDD2.n20 VDD2.n19 10.4732
R59 VDD2.n52 VDD2.n31 9.69747
R60 VDD2.n23 VDD2.n2 9.69747
R61 VDD2.n55 VDD2.n54 9.45567
R62 VDD2.n26 VDD2.n25 9.45567
R63 VDD2.n54 VDD2.n53 9.3005
R64 VDD2.n31 VDD2.n30 9.3005
R65 VDD2.n48 VDD2.n47 9.3005
R66 VDD2.n46 VDD2.n45 9.3005
R67 VDD2.n35 VDD2.n34 9.3005
R68 VDD2.n40 VDD2.n39 9.3005
R69 VDD2.n25 VDD2.n24 9.3005
R70 VDD2.n2 VDD2.n1 9.3005
R71 VDD2.n19 VDD2.n18 9.3005
R72 VDD2.n17 VDD2.n16 9.3005
R73 VDD2.n6 VDD2.n5 9.3005
R74 VDD2.n11 VDD2.n10 9.3005
R75 VDD2.n53 VDD2.n29 8.92171
R76 VDD2.n24 VDD2.n0 8.92171
R77 VDD2.n57 VDD2.t3 6.13352
R78 VDD2.n57 VDD2.t2 6.13352
R79 VDD2.n27 VDD2.t1 6.13352
R80 VDD2.n27 VDD2.t4 6.13352
R81 VDD2.n55 VDD2.n29 5.04292
R82 VDD2.n26 VDD2.n0 5.04292
R83 VDD2.n53 VDD2.n52 4.26717
R84 VDD2.n24 VDD2.n23 4.26717
R85 VDD2.n39 VDD2.n38 3.71853
R86 VDD2.n10 VDD2.n9 3.71853
R87 VDD2.n49 VDD2.n31 3.49141
R88 VDD2.n20 VDD2.n2 3.49141
R89 VDD2.n48 VDD2.n33 2.71565
R90 VDD2.n19 VDD2.n4 2.71565
R91 VDD2.n45 VDD2.n44 1.93989
R92 VDD2.n16 VDD2.n15 1.93989
R93 VDD2.n41 VDD2.n35 1.16414
R94 VDD2.n12 VDD2.n6 1.16414
R95 VDD2 VDD2.n56 0.672914
R96 VDD2.n40 VDD2.n37 0.388379
R97 VDD2.n11 VDD2.n8 0.388379
R98 VDD2.n54 VDD2.n30 0.155672
R99 VDD2.n47 VDD2.n30 0.155672
R100 VDD2.n47 VDD2.n46 0.155672
R101 VDD2.n46 VDD2.n34 0.155672
R102 VDD2.n39 VDD2.n34 0.155672
R103 VDD2.n10 VDD2.n5 0.155672
R104 VDD2.n17 VDD2.n5 0.155672
R105 VDD2.n18 VDD2.n17 0.155672
R106 VDD2.n18 VDD2.n1 0.155672
R107 VDD2.n25 VDD2.n1 0.155672
R108 VTAIL.n114 VTAIL.n92 756.745
R109 VTAIL.n24 VTAIL.n2 756.745
R110 VTAIL.n86 VTAIL.n64 756.745
R111 VTAIL.n56 VTAIL.n34 756.745
R112 VTAIL.n100 VTAIL.n99 585
R113 VTAIL.n105 VTAIL.n104 585
R114 VTAIL.n107 VTAIL.n106 585
R115 VTAIL.n96 VTAIL.n95 585
R116 VTAIL.n113 VTAIL.n112 585
R117 VTAIL.n115 VTAIL.n114 585
R118 VTAIL.n10 VTAIL.n9 585
R119 VTAIL.n15 VTAIL.n14 585
R120 VTAIL.n17 VTAIL.n16 585
R121 VTAIL.n6 VTAIL.n5 585
R122 VTAIL.n23 VTAIL.n22 585
R123 VTAIL.n25 VTAIL.n24 585
R124 VTAIL.n87 VTAIL.n86 585
R125 VTAIL.n85 VTAIL.n84 585
R126 VTAIL.n68 VTAIL.n67 585
R127 VTAIL.n79 VTAIL.n78 585
R128 VTAIL.n77 VTAIL.n76 585
R129 VTAIL.n72 VTAIL.n71 585
R130 VTAIL.n57 VTAIL.n56 585
R131 VTAIL.n55 VTAIL.n54 585
R132 VTAIL.n38 VTAIL.n37 585
R133 VTAIL.n49 VTAIL.n48 585
R134 VTAIL.n47 VTAIL.n46 585
R135 VTAIL.n42 VTAIL.n41 585
R136 VTAIL.n101 VTAIL.t7 327.856
R137 VTAIL.n11 VTAIL.t4 327.856
R138 VTAIL.n73 VTAIL.t2 327.856
R139 VTAIL.n43 VTAIL.t9 327.856
R140 VTAIL.n105 VTAIL.n99 171.744
R141 VTAIL.n106 VTAIL.n105 171.744
R142 VTAIL.n106 VTAIL.n95 171.744
R143 VTAIL.n113 VTAIL.n95 171.744
R144 VTAIL.n114 VTAIL.n113 171.744
R145 VTAIL.n15 VTAIL.n9 171.744
R146 VTAIL.n16 VTAIL.n15 171.744
R147 VTAIL.n16 VTAIL.n5 171.744
R148 VTAIL.n23 VTAIL.n5 171.744
R149 VTAIL.n24 VTAIL.n23 171.744
R150 VTAIL.n86 VTAIL.n85 171.744
R151 VTAIL.n85 VTAIL.n67 171.744
R152 VTAIL.n78 VTAIL.n67 171.744
R153 VTAIL.n78 VTAIL.n77 171.744
R154 VTAIL.n77 VTAIL.n71 171.744
R155 VTAIL.n56 VTAIL.n55 171.744
R156 VTAIL.n55 VTAIL.n37 171.744
R157 VTAIL.n48 VTAIL.n37 171.744
R158 VTAIL.n48 VTAIL.n47 171.744
R159 VTAIL.n47 VTAIL.n41 171.744
R160 VTAIL.t7 VTAIL.n99 85.8723
R161 VTAIL.t4 VTAIL.n9 85.8723
R162 VTAIL.t2 VTAIL.n71 85.8723
R163 VTAIL.t9 VTAIL.n41 85.8723
R164 VTAIL.n63 VTAIL.n62 81.04
R165 VTAIL.n33 VTAIL.n32 81.04
R166 VTAIL.n1 VTAIL.n0 81.0399
R167 VTAIL.n31 VTAIL.n30 81.0399
R168 VTAIL.n119 VTAIL.n118 32.5732
R169 VTAIL.n29 VTAIL.n28 32.5732
R170 VTAIL.n91 VTAIL.n90 32.5732
R171 VTAIL.n61 VTAIL.n60 32.5732
R172 VTAIL.n33 VTAIL.n31 18.5738
R173 VTAIL.n119 VTAIL.n91 17.7548
R174 VTAIL.n101 VTAIL.n100 16.381
R175 VTAIL.n11 VTAIL.n10 16.381
R176 VTAIL.n73 VTAIL.n72 16.381
R177 VTAIL.n43 VTAIL.n42 16.381
R178 VTAIL.n104 VTAIL.n103 12.8005
R179 VTAIL.n14 VTAIL.n13 12.8005
R180 VTAIL.n76 VTAIL.n75 12.8005
R181 VTAIL.n46 VTAIL.n45 12.8005
R182 VTAIL.n107 VTAIL.n98 12.0247
R183 VTAIL.n17 VTAIL.n8 12.0247
R184 VTAIL.n79 VTAIL.n70 12.0247
R185 VTAIL.n49 VTAIL.n40 12.0247
R186 VTAIL.n108 VTAIL.n96 11.249
R187 VTAIL.n18 VTAIL.n6 11.249
R188 VTAIL.n80 VTAIL.n68 11.249
R189 VTAIL.n50 VTAIL.n38 11.249
R190 VTAIL.n112 VTAIL.n111 10.4732
R191 VTAIL.n22 VTAIL.n21 10.4732
R192 VTAIL.n84 VTAIL.n83 10.4732
R193 VTAIL.n54 VTAIL.n53 10.4732
R194 VTAIL.n115 VTAIL.n94 9.69747
R195 VTAIL.n25 VTAIL.n4 9.69747
R196 VTAIL.n87 VTAIL.n66 9.69747
R197 VTAIL.n57 VTAIL.n36 9.69747
R198 VTAIL.n118 VTAIL.n117 9.45567
R199 VTAIL.n28 VTAIL.n27 9.45567
R200 VTAIL.n90 VTAIL.n89 9.45567
R201 VTAIL.n60 VTAIL.n59 9.45567
R202 VTAIL.n117 VTAIL.n116 9.3005
R203 VTAIL.n94 VTAIL.n93 9.3005
R204 VTAIL.n111 VTAIL.n110 9.3005
R205 VTAIL.n109 VTAIL.n108 9.3005
R206 VTAIL.n98 VTAIL.n97 9.3005
R207 VTAIL.n103 VTAIL.n102 9.3005
R208 VTAIL.n27 VTAIL.n26 9.3005
R209 VTAIL.n4 VTAIL.n3 9.3005
R210 VTAIL.n21 VTAIL.n20 9.3005
R211 VTAIL.n19 VTAIL.n18 9.3005
R212 VTAIL.n8 VTAIL.n7 9.3005
R213 VTAIL.n13 VTAIL.n12 9.3005
R214 VTAIL.n89 VTAIL.n88 9.3005
R215 VTAIL.n66 VTAIL.n65 9.3005
R216 VTAIL.n83 VTAIL.n82 9.3005
R217 VTAIL.n81 VTAIL.n80 9.3005
R218 VTAIL.n70 VTAIL.n69 9.3005
R219 VTAIL.n75 VTAIL.n74 9.3005
R220 VTAIL.n59 VTAIL.n58 9.3005
R221 VTAIL.n36 VTAIL.n35 9.3005
R222 VTAIL.n53 VTAIL.n52 9.3005
R223 VTAIL.n51 VTAIL.n50 9.3005
R224 VTAIL.n40 VTAIL.n39 9.3005
R225 VTAIL.n45 VTAIL.n44 9.3005
R226 VTAIL.n116 VTAIL.n92 8.92171
R227 VTAIL.n26 VTAIL.n2 8.92171
R228 VTAIL.n88 VTAIL.n64 8.92171
R229 VTAIL.n58 VTAIL.n34 8.92171
R230 VTAIL.n0 VTAIL.t10 6.13352
R231 VTAIL.n0 VTAIL.t8 6.13352
R232 VTAIL.n30 VTAIL.t1 6.13352
R233 VTAIL.n30 VTAIL.t0 6.13352
R234 VTAIL.n62 VTAIL.t5 6.13352
R235 VTAIL.n62 VTAIL.t3 6.13352
R236 VTAIL.n32 VTAIL.t6 6.13352
R237 VTAIL.n32 VTAIL.t11 6.13352
R238 VTAIL.n118 VTAIL.n92 5.04292
R239 VTAIL.n28 VTAIL.n2 5.04292
R240 VTAIL.n90 VTAIL.n64 5.04292
R241 VTAIL.n60 VTAIL.n34 5.04292
R242 VTAIL.n116 VTAIL.n115 4.26717
R243 VTAIL.n26 VTAIL.n25 4.26717
R244 VTAIL.n88 VTAIL.n87 4.26717
R245 VTAIL.n58 VTAIL.n57 4.26717
R246 VTAIL.n74 VTAIL.n73 3.71853
R247 VTAIL.n44 VTAIL.n43 3.71853
R248 VTAIL.n102 VTAIL.n101 3.71853
R249 VTAIL.n12 VTAIL.n11 3.71853
R250 VTAIL.n112 VTAIL.n94 3.49141
R251 VTAIL.n22 VTAIL.n4 3.49141
R252 VTAIL.n84 VTAIL.n66 3.49141
R253 VTAIL.n54 VTAIL.n36 3.49141
R254 VTAIL.n111 VTAIL.n96 2.71565
R255 VTAIL.n21 VTAIL.n6 2.71565
R256 VTAIL.n83 VTAIL.n68 2.71565
R257 VTAIL.n53 VTAIL.n38 2.71565
R258 VTAIL.n108 VTAIL.n107 1.93989
R259 VTAIL.n18 VTAIL.n17 1.93989
R260 VTAIL.n80 VTAIL.n79 1.93989
R261 VTAIL.n50 VTAIL.n49 1.93989
R262 VTAIL.n104 VTAIL.n98 1.16414
R263 VTAIL.n14 VTAIL.n8 1.16414
R264 VTAIL.n76 VTAIL.n70 1.16414
R265 VTAIL.n46 VTAIL.n40 1.16414
R266 VTAIL.n63 VTAIL.n61 0.87981
R267 VTAIL.n29 VTAIL.n1 0.87981
R268 VTAIL.n61 VTAIL.n33 0.819465
R269 VTAIL.n91 VTAIL.n63 0.819465
R270 VTAIL.n31 VTAIL.n29 0.819465
R271 VTAIL VTAIL.n119 0.556535
R272 VTAIL.n103 VTAIL.n100 0.388379
R273 VTAIL.n13 VTAIL.n10 0.388379
R274 VTAIL.n75 VTAIL.n72 0.388379
R275 VTAIL.n45 VTAIL.n42 0.388379
R276 VTAIL VTAIL.n1 0.263431
R277 VTAIL.n102 VTAIL.n97 0.155672
R278 VTAIL.n109 VTAIL.n97 0.155672
R279 VTAIL.n110 VTAIL.n109 0.155672
R280 VTAIL.n110 VTAIL.n93 0.155672
R281 VTAIL.n117 VTAIL.n93 0.155672
R282 VTAIL.n12 VTAIL.n7 0.155672
R283 VTAIL.n19 VTAIL.n7 0.155672
R284 VTAIL.n20 VTAIL.n19 0.155672
R285 VTAIL.n20 VTAIL.n3 0.155672
R286 VTAIL.n27 VTAIL.n3 0.155672
R287 VTAIL.n89 VTAIL.n65 0.155672
R288 VTAIL.n82 VTAIL.n65 0.155672
R289 VTAIL.n82 VTAIL.n81 0.155672
R290 VTAIL.n81 VTAIL.n69 0.155672
R291 VTAIL.n74 VTAIL.n69 0.155672
R292 VTAIL.n59 VTAIL.n35 0.155672
R293 VTAIL.n52 VTAIL.n35 0.155672
R294 VTAIL.n52 VTAIL.n51 0.155672
R295 VTAIL.n51 VTAIL.n39 0.155672
R296 VTAIL.n44 VTAIL.n39 0.155672
R297 VP.n1 VP.t0 296.197
R298 VP.n6 VP.t5 269.377
R299 VP.n7 VP.t4 269.377
R300 VP.n8 VP.t2 269.377
R301 VP.n3 VP.t1 269.377
R302 VP.n2 VP.t3 269.377
R303 VP.n9 VP.n8 161.3
R304 VP.n4 VP.n3 161.3
R305 VP.n6 VP.n5 161.3
R306 VP.n7 VP.n0 80.6037
R307 VP.n7 VP.n6 48.2005
R308 VP.n8 VP.n7 48.2005
R309 VP.n3 VP.n2 48.2005
R310 VP.n4 VP.n1 45.1367
R311 VP.n5 VP.n4 35.921
R312 VP.n2 VP.n1 13.3799
R313 VP.n5 VP.n0 0.285035
R314 VP.n9 VP.n0 0.285035
R315 VP VP.n9 0.0516364
R316 VDD1.n22 VDD1.n0 756.745
R317 VDD1.n49 VDD1.n27 756.745
R318 VDD1.n23 VDD1.n22 585
R319 VDD1.n21 VDD1.n20 585
R320 VDD1.n4 VDD1.n3 585
R321 VDD1.n15 VDD1.n14 585
R322 VDD1.n13 VDD1.n12 585
R323 VDD1.n8 VDD1.n7 585
R324 VDD1.n35 VDD1.n34 585
R325 VDD1.n40 VDD1.n39 585
R326 VDD1.n42 VDD1.n41 585
R327 VDD1.n31 VDD1.n30 585
R328 VDD1.n48 VDD1.n47 585
R329 VDD1.n50 VDD1.n49 585
R330 VDD1.n9 VDD1.t5 327.856
R331 VDD1.n36 VDD1.t0 327.856
R332 VDD1.n22 VDD1.n21 171.744
R333 VDD1.n21 VDD1.n3 171.744
R334 VDD1.n14 VDD1.n3 171.744
R335 VDD1.n14 VDD1.n13 171.744
R336 VDD1.n13 VDD1.n7 171.744
R337 VDD1.n40 VDD1.n34 171.744
R338 VDD1.n41 VDD1.n40 171.744
R339 VDD1.n41 VDD1.n30 171.744
R340 VDD1.n48 VDD1.n30 171.744
R341 VDD1.n49 VDD1.n48 171.744
R342 VDD1.n55 VDD1.n54 97.868
R343 VDD1.n57 VDD1.n56 97.7186
R344 VDD1.t5 VDD1.n7 85.8723
R345 VDD1.t0 VDD1.n34 85.8723
R346 VDD1 VDD1.n26 49.9244
R347 VDD1.n55 VDD1.n53 49.8109
R348 VDD1.n57 VDD1.n55 31.9384
R349 VDD1.n9 VDD1.n8 16.381
R350 VDD1.n36 VDD1.n35 16.381
R351 VDD1.n12 VDD1.n11 12.8005
R352 VDD1.n39 VDD1.n38 12.8005
R353 VDD1.n15 VDD1.n6 12.0247
R354 VDD1.n42 VDD1.n33 12.0247
R355 VDD1.n16 VDD1.n4 11.249
R356 VDD1.n43 VDD1.n31 11.249
R357 VDD1.n20 VDD1.n19 10.4732
R358 VDD1.n47 VDD1.n46 10.4732
R359 VDD1.n23 VDD1.n2 9.69747
R360 VDD1.n50 VDD1.n29 9.69747
R361 VDD1.n26 VDD1.n25 9.45567
R362 VDD1.n53 VDD1.n52 9.45567
R363 VDD1.n25 VDD1.n24 9.3005
R364 VDD1.n2 VDD1.n1 9.3005
R365 VDD1.n19 VDD1.n18 9.3005
R366 VDD1.n17 VDD1.n16 9.3005
R367 VDD1.n6 VDD1.n5 9.3005
R368 VDD1.n11 VDD1.n10 9.3005
R369 VDD1.n52 VDD1.n51 9.3005
R370 VDD1.n29 VDD1.n28 9.3005
R371 VDD1.n46 VDD1.n45 9.3005
R372 VDD1.n44 VDD1.n43 9.3005
R373 VDD1.n33 VDD1.n32 9.3005
R374 VDD1.n38 VDD1.n37 9.3005
R375 VDD1.n24 VDD1.n0 8.92171
R376 VDD1.n51 VDD1.n27 8.92171
R377 VDD1.n56 VDD1.t2 6.13352
R378 VDD1.n56 VDD1.t4 6.13352
R379 VDD1.n54 VDD1.t1 6.13352
R380 VDD1.n54 VDD1.t3 6.13352
R381 VDD1.n26 VDD1.n0 5.04292
R382 VDD1.n53 VDD1.n27 5.04292
R383 VDD1.n24 VDD1.n23 4.26717
R384 VDD1.n51 VDD1.n50 4.26717
R385 VDD1.n10 VDD1.n9 3.71853
R386 VDD1.n37 VDD1.n36 3.71853
R387 VDD1.n20 VDD1.n2 3.49141
R388 VDD1.n47 VDD1.n29 3.49141
R389 VDD1.n19 VDD1.n4 2.71565
R390 VDD1.n46 VDD1.n31 2.71565
R391 VDD1.n16 VDD1.n15 1.93989
R392 VDD1.n43 VDD1.n42 1.93989
R393 VDD1.n12 VDD1.n6 1.16414
R394 VDD1.n39 VDD1.n33 1.16414
R395 VDD1.n11 VDD1.n8 0.388379
R396 VDD1.n38 VDD1.n35 0.388379
R397 VDD1.n25 VDD1.n1 0.155672
R398 VDD1.n18 VDD1.n1 0.155672
R399 VDD1.n18 VDD1.n17 0.155672
R400 VDD1.n17 VDD1.n5 0.155672
R401 VDD1.n10 VDD1.n5 0.155672
R402 VDD1.n37 VDD1.n32 0.155672
R403 VDD1.n44 VDD1.n32 0.155672
R404 VDD1.n45 VDD1.n44 0.155672
R405 VDD1.n45 VDD1.n28 0.155672
R406 VDD1.n52 VDD1.n28 0.155672
R407 VDD1 VDD1.n57 0.147052
R408 B.n270 B.n269 585
R409 B.n271 B.n42 585
R410 B.n273 B.n272 585
R411 B.n274 B.n41 585
R412 B.n276 B.n275 585
R413 B.n277 B.n40 585
R414 B.n279 B.n278 585
R415 B.n280 B.n39 585
R416 B.n282 B.n281 585
R417 B.n283 B.n38 585
R418 B.n285 B.n284 585
R419 B.n286 B.n37 585
R420 B.n288 B.n287 585
R421 B.n289 B.n36 585
R422 B.n291 B.n290 585
R423 B.n292 B.n35 585
R424 B.n294 B.n293 585
R425 B.n295 B.n34 585
R426 B.n297 B.n296 585
R427 B.n298 B.n33 585
R428 B.n300 B.n299 585
R429 B.n301 B.n30 585
R430 B.n304 B.n303 585
R431 B.n305 B.n29 585
R432 B.n307 B.n306 585
R433 B.n308 B.n28 585
R434 B.n310 B.n309 585
R435 B.n311 B.n27 585
R436 B.n313 B.n312 585
R437 B.n314 B.n23 585
R438 B.n316 B.n315 585
R439 B.n317 B.n22 585
R440 B.n319 B.n318 585
R441 B.n320 B.n21 585
R442 B.n322 B.n321 585
R443 B.n323 B.n20 585
R444 B.n325 B.n324 585
R445 B.n326 B.n19 585
R446 B.n328 B.n327 585
R447 B.n329 B.n18 585
R448 B.n331 B.n330 585
R449 B.n332 B.n17 585
R450 B.n334 B.n333 585
R451 B.n335 B.n16 585
R452 B.n337 B.n336 585
R453 B.n338 B.n15 585
R454 B.n340 B.n339 585
R455 B.n341 B.n14 585
R456 B.n343 B.n342 585
R457 B.n344 B.n13 585
R458 B.n346 B.n345 585
R459 B.n347 B.n12 585
R460 B.n349 B.n348 585
R461 B.n268 B.n43 585
R462 B.n267 B.n266 585
R463 B.n265 B.n44 585
R464 B.n264 B.n263 585
R465 B.n262 B.n45 585
R466 B.n261 B.n260 585
R467 B.n259 B.n46 585
R468 B.n258 B.n257 585
R469 B.n256 B.n47 585
R470 B.n255 B.n254 585
R471 B.n253 B.n48 585
R472 B.n252 B.n251 585
R473 B.n250 B.n49 585
R474 B.n249 B.n248 585
R475 B.n247 B.n50 585
R476 B.n246 B.n245 585
R477 B.n244 B.n51 585
R478 B.n243 B.n242 585
R479 B.n241 B.n52 585
R480 B.n240 B.n239 585
R481 B.n238 B.n53 585
R482 B.n237 B.n236 585
R483 B.n235 B.n54 585
R484 B.n234 B.n233 585
R485 B.n232 B.n55 585
R486 B.n231 B.n230 585
R487 B.n229 B.n56 585
R488 B.n228 B.n227 585
R489 B.n226 B.n57 585
R490 B.n225 B.n224 585
R491 B.n223 B.n58 585
R492 B.n222 B.n221 585
R493 B.n220 B.n59 585
R494 B.n219 B.n218 585
R495 B.n217 B.n60 585
R496 B.n216 B.n215 585
R497 B.n214 B.n61 585
R498 B.n213 B.n212 585
R499 B.n211 B.n62 585
R500 B.n128 B.n127 585
R501 B.n129 B.n90 585
R502 B.n131 B.n130 585
R503 B.n132 B.n89 585
R504 B.n134 B.n133 585
R505 B.n135 B.n88 585
R506 B.n137 B.n136 585
R507 B.n138 B.n87 585
R508 B.n140 B.n139 585
R509 B.n141 B.n86 585
R510 B.n143 B.n142 585
R511 B.n144 B.n85 585
R512 B.n146 B.n145 585
R513 B.n147 B.n84 585
R514 B.n149 B.n148 585
R515 B.n150 B.n83 585
R516 B.n152 B.n151 585
R517 B.n153 B.n82 585
R518 B.n155 B.n154 585
R519 B.n156 B.n81 585
R520 B.n158 B.n157 585
R521 B.n159 B.n78 585
R522 B.n162 B.n161 585
R523 B.n163 B.n77 585
R524 B.n165 B.n164 585
R525 B.n166 B.n76 585
R526 B.n168 B.n167 585
R527 B.n169 B.n75 585
R528 B.n171 B.n170 585
R529 B.n172 B.n74 585
R530 B.n177 B.n176 585
R531 B.n178 B.n73 585
R532 B.n180 B.n179 585
R533 B.n181 B.n72 585
R534 B.n183 B.n182 585
R535 B.n184 B.n71 585
R536 B.n186 B.n185 585
R537 B.n187 B.n70 585
R538 B.n189 B.n188 585
R539 B.n190 B.n69 585
R540 B.n192 B.n191 585
R541 B.n193 B.n68 585
R542 B.n195 B.n194 585
R543 B.n196 B.n67 585
R544 B.n198 B.n197 585
R545 B.n199 B.n66 585
R546 B.n201 B.n200 585
R547 B.n202 B.n65 585
R548 B.n204 B.n203 585
R549 B.n205 B.n64 585
R550 B.n207 B.n206 585
R551 B.n208 B.n63 585
R552 B.n210 B.n209 585
R553 B.n126 B.n91 585
R554 B.n125 B.n124 585
R555 B.n123 B.n92 585
R556 B.n122 B.n121 585
R557 B.n120 B.n93 585
R558 B.n119 B.n118 585
R559 B.n117 B.n94 585
R560 B.n116 B.n115 585
R561 B.n114 B.n95 585
R562 B.n113 B.n112 585
R563 B.n111 B.n96 585
R564 B.n110 B.n109 585
R565 B.n108 B.n97 585
R566 B.n107 B.n106 585
R567 B.n105 B.n98 585
R568 B.n104 B.n103 585
R569 B.n102 B.n99 585
R570 B.n101 B.n100 585
R571 B.n2 B.n0 585
R572 B.n377 B.n1 585
R573 B.n376 B.n375 585
R574 B.n374 B.n3 585
R575 B.n373 B.n372 585
R576 B.n371 B.n4 585
R577 B.n370 B.n369 585
R578 B.n368 B.n5 585
R579 B.n367 B.n366 585
R580 B.n365 B.n6 585
R581 B.n364 B.n363 585
R582 B.n362 B.n7 585
R583 B.n361 B.n360 585
R584 B.n359 B.n8 585
R585 B.n358 B.n357 585
R586 B.n356 B.n9 585
R587 B.n355 B.n354 585
R588 B.n353 B.n10 585
R589 B.n352 B.n351 585
R590 B.n350 B.n11 585
R591 B.n379 B.n378 585
R592 B.n127 B.n126 578.989
R593 B.n348 B.n11 578.989
R594 B.n209 B.n62 578.989
R595 B.n269 B.n268 578.989
R596 B.n173 B.t0 410.091
R597 B.n79 B.t3 410.091
R598 B.n24 B.t6 410.091
R599 B.n31 B.t9 410.091
R600 B.n173 B.t2 274.461
R601 B.n31 B.t10 274.461
R602 B.n79 B.t5 274.461
R603 B.n24 B.t7 274.461
R604 B.n174 B.t1 256.036
R605 B.n32 B.t11 256.036
R606 B.n80 B.t4 256.036
R607 B.n25 B.t8 256.036
R608 B.n126 B.n125 163.367
R609 B.n125 B.n92 163.367
R610 B.n121 B.n92 163.367
R611 B.n121 B.n120 163.367
R612 B.n120 B.n119 163.367
R613 B.n119 B.n94 163.367
R614 B.n115 B.n94 163.367
R615 B.n115 B.n114 163.367
R616 B.n114 B.n113 163.367
R617 B.n113 B.n96 163.367
R618 B.n109 B.n96 163.367
R619 B.n109 B.n108 163.367
R620 B.n108 B.n107 163.367
R621 B.n107 B.n98 163.367
R622 B.n103 B.n98 163.367
R623 B.n103 B.n102 163.367
R624 B.n102 B.n101 163.367
R625 B.n101 B.n2 163.367
R626 B.n378 B.n2 163.367
R627 B.n378 B.n377 163.367
R628 B.n377 B.n376 163.367
R629 B.n376 B.n3 163.367
R630 B.n372 B.n3 163.367
R631 B.n372 B.n371 163.367
R632 B.n371 B.n370 163.367
R633 B.n370 B.n5 163.367
R634 B.n366 B.n5 163.367
R635 B.n366 B.n365 163.367
R636 B.n365 B.n364 163.367
R637 B.n364 B.n7 163.367
R638 B.n360 B.n7 163.367
R639 B.n360 B.n359 163.367
R640 B.n359 B.n358 163.367
R641 B.n358 B.n9 163.367
R642 B.n354 B.n9 163.367
R643 B.n354 B.n353 163.367
R644 B.n353 B.n352 163.367
R645 B.n352 B.n11 163.367
R646 B.n127 B.n90 163.367
R647 B.n131 B.n90 163.367
R648 B.n132 B.n131 163.367
R649 B.n133 B.n132 163.367
R650 B.n133 B.n88 163.367
R651 B.n137 B.n88 163.367
R652 B.n138 B.n137 163.367
R653 B.n139 B.n138 163.367
R654 B.n139 B.n86 163.367
R655 B.n143 B.n86 163.367
R656 B.n144 B.n143 163.367
R657 B.n145 B.n144 163.367
R658 B.n145 B.n84 163.367
R659 B.n149 B.n84 163.367
R660 B.n150 B.n149 163.367
R661 B.n151 B.n150 163.367
R662 B.n151 B.n82 163.367
R663 B.n155 B.n82 163.367
R664 B.n156 B.n155 163.367
R665 B.n157 B.n156 163.367
R666 B.n157 B.n78 163.367
R667 B.n162 B.n78 163.367
R668 B.n163 B.n162 163.367
R669 B.n164 B.n163 163.367
R670 B.n164 B.n76 163.367
R671 B.n168 B.n76 163.367
R672 B.n169 B.n168 163.367
R673 B.n170 B.n169 163.367
R674 B.n170 B.n74 163.367
R675 B.n177 B.n74 163.367
R676 B.n178 B.n177 163.367
R677 B.n179 B.n178 163.367
R678 B.n179 B.n72 163.367
R679 B.n183 B.n72 163.367
R680 B.n184 B.n183 163.367
R681 B.n185 B.n184 163.367
R682 B.n185 B.n70 163.367
R683 B.n189 B.n70 163.367
R684 B.n190 B.n189 163.367
R685 B.n191 B.n190 163.367
R686 B.n191 B.n68 163.367
R687 B.n195 B.n68 163.367
R688 B.n196 B.n195 163.367
R689 B.n197 B.n196 163.367
R690 B.n197 B.n66 163.367
R691 B.n201 B.n66 163.367
R692 B.n202 B.n201 163.367
R693 B.n203 B.n202 163.367
R694 B.n203 B.n64 163.367
R695 B.n207 B.n64 163.367
R696 B.n208 B.n207 163.367
R697 B.n209 B.n208 163.367
R698 B.n213 B.n62 163.367
R699 B.n214 B.n213 163.367
R700 B.n215 B.n214 163.367
R701 B.n215 B.n60 163.367
R702 B.n219 B.n60 163.367
R703 B.n220 B.n219 163.367
R704 B.n221 B.n220 163.367
R705 B.n221 B.n58 163.367
R706 B.n225 B.n58 163.367
R707 B.n226 B.n225 163.367
R708 B.n227 B.n226 163.367
R709 B.n227 B.n56 163.367
R710 B.n231 B.n56 163.367
R711 B.n232 B.n231 163.367
R712 B.n233 B.n232 163.367
R713 B.n233 B.n54 163.367
R714 B.n237 B.n54 163.367
R715 B.n238 B.n237 163.367
R716 B.n239 B.n238 163.367
R717 B.n239 B.n52 163.367
R718 B.n243 B.n52 163.367
R719 B.n244 B.n243 163.367
R720 B.n245 B.n244 163.367
R721 B.n245 B.n50 163.367
R722 B.n249 B.n50 163.367
R723 B.n250 B.n249 163.367
R724 B.n251 B.n250 163.367
R725 B.n251 B.n48 163.367
R726 B.n255 B.n48 163.367
R727 B.n256 B.n255 163.367
R728 B.n257 B.n256 163.367
R729 B.n257 B.n46 163.367
R730 B.n261 B.n46 163.367
R731 B.n262 B.n261 163.367
R732 B.n263 B.n262 163.367
R733 B.n263 B.n44 163.367
R734 B.n267 B.n44 163.367
R735 B.n268 B.n267 163.367
R736 B.n348 B.n347 163.367
R737 B.n347 B.n346 163.367
R738 B.n346 B.n13 163.367
R739 B.n342 B.n13 163.367
R740 B.n342 B.n341 163.367
R741 B.n341 B.n340 163.367
R742 B.n340 B.n15 163.367
R743 B.n336 B.n15 163.367
R744 B.n336 B.n335 163.367
R745 B.n335 B.n334 163.367
R746 B.n334 B.n17 163.367
R747 B.n330 B.n17 163.367
R748 B.n330 B.n329 163.367
R749 B.n329 B.n328 163.367
R750 B.n328 B.n19 163.367
R751 B.n324 B.n19 163.367
R752 B.n324 B.n323 163.367
R753 B.n323 B.n322 163.367
R754 B.n322 B.n21 163.367
R755 B.n318 B.n21 163.367
R756 B.n318 B.n317 163.367
R757 B.n317 B.n316 163.367
R758 B.n316 B.n23 163.367
R759 B.n312 B.n23 163.367
R760 B.n312 B.n311 163.367
R761 B.n311 B.n310 163.367
R762 B.n310 B.n28 163.367
R763 B.n306 B.n28 163.367
R764 B.n306 B.n305 163.367
R765 B.n305 B.n304 163.367
R766 B.n304 B.n30 163.367
R767 B.n299 B.n30 163.367
R768 B.n299 B.n298 163.367
R769 B.n298 B.n297 163.367
R770 B.n297 B.n34 163.367
R771 B.n293 B.n34 163.367
R772 B.n293 B.n292 163.367
R773 B.n292 B.n291 163.367
R774 B.n291 B.n36 163.367
R775 B.n287 B.n36 163.367
R776 B.n287 B.n286 163.367
R777 B.n286 B.n285 163.367
R778 B.n285 B.n38 163.367
R779 B.n281 B.n38 163.367
R780 B.n281 B.n280 163.367
R781 B.n280 B.n279 163.367
R782 B.n279 B.n40 163.367
R783 B.n275 B.n40 163.367
R784 B.n275 B.n274 163.367
R785 B.n274 B.n273 163.367
R786 B.n273 B.n42 163.367
R787 B.n269 B.n42 163.367
R788 B.n175 B.n174 59.5399
R789 B.n160 B.n80 59.5399
R790 B.n26 B.n25 59.5399
R791 B.n302 B.n32 59.5399
R792 B.n350 B.n349 37.62
R793 B.n270 B.n43 37.62
R794 B.n211 B.n210 37.62
R795 B.n128 B.n91 37.62
R796 B.n174 B.n173 18.4247
R797 B.n80 B.n79 18.4247
R798 B.n25 B.n24 18.4247
R799 B.n32 B.n31 18.4247
R800 B B.n379 18.0485
R801 B.n349 B.n12 10.6151
R802 B.n345 B.n12 10.6151
R803 B.n345 B.n344 10.6151
R804 B.n344 B.n343 10.6151
R805 B.n343 B.n14 10.6151
R806 B.n339 B.n14 10.6151
R807 B.n339 B.n338 10.6151
R808 B.n338 B.n337 10.6151
R809 B.n337 B.n16 10.6151
R810 B.n333 B.n16 10.6151
R811 B.n333 B.n332 10.6151
R812 B.n332 B.n331 10.6151
R813 B.n331 B.n18 10.6151
R814 B.n327 B.n18 10.6151
R815 B.n327 B.n326 10.6151
R816 B.n326 B.n325 10.6151
R817 B.n325 B.n20 10.6151
R818 B.n321 B.n20 10.6151
R819 B.n321 B.n320 10.6151
R820 B.n320 B.n319 10.6151
R821 B.n319 B.n22 10.6151
R822 B.n315 B.n314 10.6151
R823 B.n314 B.n313 10.6151
R824 B.n313 B.n27 10.6151
R825 B.n309 B.n27 10.6151
R826 B.n309 B.n308 10.6151
R827 B.n308 B.n307 10.6151
R828 B.n307 B.n29 10.6151
R829 B.n303 B.n29 10.6151
R830 B.n301 B.n300 10.6151
R831 B.n300 B.n33 10.6151
R832 B.n296 B.n33 10.6151
R833 B.n296 B.n295 10.6151
R834 B.n295 B.n294 10.6151
R835 B.n294 B.n35 10.6151
R836 B.n290 B.n35 10.6151
R837 B.n290 B.n289 10.6151
R838 B.n289 B.n288 10.6151
R839 B.n288 B.n37 10.6151
R840 B.n284 B.n37 10.6151
R841 B.n284 B.n283 10.6151
R842 B.n283 B.n282 10.6151
R843 B.n282 B.n39 10.6151
R844 B.n278 B.n39 10.6151
R845 B.n278 B.n277 10.6151
R846 B.n277 B.n276 10.6151
R847 B.n276 B.n41 10.6151
R848 B.n272 B.n41 10.6151
R849 B.n272 B.n271 10.6151
R850 B.n271 B.n270 10.6151
R851 B.n212 B.n211 10.6151
R852 B.n212 B.n61 10.6151
R853 B.n216 B.n61 10.6151
R854 B.n217 B.n216 10.6151
R855 B.n218 B.n217 10.6151
R856 B.n218 B.n59 10.6151
R857 B.n222 B.n59 10.6151
R858 B.n223 B.n222 10.6151
R859 B.n224 B.n223 10.6151
R860 B.n224 B.n57 10.6151
R861 B.n228 B.n57 10.6151
R862 B.n229 B.n228 10.6151
R863 B.n230 B.n229 10.6151
R864 B.n230 B.n55 10.6151
R865 B.n234 B.n55 10.6151
R866 B.n235 B.n234 10.6151
R867 B.n236 B.n235 10.6151
R868 B.n236 B.n53 10.6151
R869 B.n240 B.n53 10.6151
R870 B.n241 B.n240 10.6151
R871 B.n242 B.n241 10.6151
R872 B.n242 B.n51 10.6151
R873 B.n246 B.n51 10.6151
R874 B.n247 B.n246 10.6151
R875 B.n248 B.n247 10.6151
R876 B.n248 B.n49 10.6151
R877 B.n252 B.n49 10.6151
R878 B.n253 B.n252 10.6151
R879 B.n254 B.n253 10.6151
R880 B.n254 B.n47 10.6151
R881 B.n258 B.n47 10.6151
R882 B.n259 B.n258 10.6151
R883 B.n260 B.n259 10.6151
R884 B.n260 B.n45 10.6151
R885 B.n264 B.n45 10.6151
R886 B.n265 B.n264 10.6151
R887 B.n266 B.n265 10.6151
R888 B.n266 B.n43 10.6151
R889 B.n129 B.n128 10.6151
R890 B.n130 B.n129 10.6151
R891 B.n130 B.n89 10.6151
R892 B.n134 B.n89 10.6151
R893 B.n135 B.n134 10.6151
R894 B.n136 B.n135 10.6151
R895 B.n136 B.n87 10.6151
R896 B.n140 B.n87 10.6151
R897 B.n141 B.n140 10.6151
R898 B.n142 B.n141 10.6151
R899 B.n142 B.n85 10.6151
R900 B.n146 B.n85 10.6151
R901 B.n147 B.n146 10.6151
R902 B.n148 B.n147 10.6151
R903 B.n148 B.n83 10.6151
R904 B.n152 B.n83 10.6151
R905 B.n153 B.n152 10.6151
R906 B.n154 B.n153 10.6151
R907 B.n154 B.n81 10.6151
R908 B.n158 B.n81 10.6151
R909 B.n159 B.n158 10.6151
R910 B.n161 B.n77 10.6151
R911 B.n165 B.n77 10.6151
R912 B.n166 B.n165 10.6151
R913 B.n167 B.n166 10.6151
R914 B.n167 B.n75 10.6151
R915 B.n171 B.n75 10.6151
R916 B.n172 B.n171 10.6151
R917 B.n176 B.n172 10.6151
R918 B.n180 B.n73 10.6151
R919 B.n181 B.n180 10.6151
R920 B.n182 B.n181 10.6151
R921 B.n182 B.n71 10.6151
R922 B.n186 B.n71 10.6151
R923 B.n187 B.n186 10.6151
R924 B.n188 B.n187 10.6151
R925 B.n188 B.n69 10.6151
R926 B.n192 B.n69 10.6151
R927 B.n193 B.n192 10.6151
R928 B.n194 B.n193 10.6151
R929 B.n194 B.n67 10.6151
R930 B.n198 B.n67 10.6151
R931 B.n199 B.n198 10.6151
R932 B.n200 B.n199 10.6151
R933 B.n200 B.n65 10.6151
R934 B.n204 B.n65 10.6151
R935 B.n205 B.n204 10.6151
R936 B.n206 B.n205 10.6151
R937 B.n206 B.n63 10.6151
R938 B.n210 B.n63 10.6151
R939 B.n124 B.n91 10.6151
R940 B.n124 B.n123 10.6151
R941 B.n123 B.n122 10.6151
R942 B.n122 B.n93 10.6151
R943 B.n118 B.n93 10.6151
R944 B.n118 B.n117 10.6151
R945 B.n117 B.n116 10.6151
R946 B.n116 B.n95 10.6151
R947 B.n112 B.n95 10.6151
R948 B.n112 B.n111 10.6151
R949 B.n111 B.n110 10.6151
R950 B.n110 B.n97 10.6151
R951 B.n106 B.n97 10.6151
R952 B.n106 B.n105 10.6151
R953 B.n105 B.n104 10.6151
R954 B.n104 B.n99 10.6151
R955 B.n100 B.n99 10.6151
R956 B.n100 B.n0 10.6151
R957 B.n375 B.n1 10.6151
R958 B.n375 B.n374 10.6151
R959 B.n374 B.n373 10.6151
R960 B.n373 B.n4 10.6151
R961 B.n369 B.n4 10.6151
R962 B.n369 B.n368 10.6151
R963 B.n368 B.n367 10.6151
R964 B.n367 B.n6 10.6151
R965 B.n363 B.n6 10.6151
R966 B.n363 B.n362 10.6151
R967 B.n362 B.n361 10.6151
R968 B.n361 B.n8 10.6151
R969 B.n357 B.n8 10.6151
R970 B.n357 B.n356 10.6151
R971 B.n356 B.n355 10.6151
R972 B.n355 B.n10 10.6151
R973 B.n351 B.n10 10.6151
R974 B.n351 B.n350 10.6151
R975 B.n315 B.n26 6.5566
R976 B.n303 B.n302 6.5566
R977 B.n161 B.n160 6.5566
R978 B.n176 B.n175 6.5566
R979 B.n26 B.n22 4.05904
R980 B.n302 B.n301 4.05904
R981 B.n160 B.n159 4.05904
R982 B.n175 B.n73 4.05904
R983 B.n379 B.n0 2.81026
R984 B.n379 B.n1 2.81026
C0 VP VTAIL 1.98789f
C1 VDD2 VN 1.98566f
C2 VP B 1.02797f
C3 VDD2 w_n1730_n2028# 1.31428f
C4 w_n1730_n2028# VN 2.65702f
C5 VTAIL VDD1 5.60676f
C6 VP VDD2 0.294148f
C7 B VDD1 1.05026f
C8 VP VN 3.7565f
C9 VP w_n1730_n2028# 2.87509f
C10 VTAIL B 1.47278f
C11 VDD2 VDD1 0.680573f
C12 VN VDD1 0.148421f
C13 VDD2 VTAIL 5.64388f
C14 w_n1730_n2028# VDD1 1.29298f
C15 VDD2 B 1.07746f
C16 VTAIL VN 1.97355f
C17 VN B 0.673722f
C18 VTAIL w_n1730_n2028# 1.86978f
C19 w_n1730_n2028# B 5.06662f
C20 VP VDD1 2.12519f
C21 VDD2 VSUBS 0.87064f
C22 VDD1 VSUBS 0.896332f
C23 VTAIL VSUBS 0.385076f
C24 VN VSUBS 3.07488f
C25 VP VSUBS 1.08699f
C26 B VSUBS 2.02036f
C27 w_n1730_n2028# VSUBS 43.9074f
C28 B.n0 VSUBS 0.004351f
C29 B.n1 VSUBS 0.004351f
C30 B.n2 VSUBS 0.006881f
C31 B.n3 VSUBS 0.006881f
C32 B.n4 VSUBS 0.006881f
C33 B.n5 VSUBS 0.006881f
C34 B.n6 VSUBS 0.006881f
C35 B.n7 VSUBS 0.006881f
C36 B.n8 VSUBS 0.006881f
C37 B.n9 VSUBS 0.006881f
C38 B.n10 VSUBS 0.006881f
C39 B.n11 VSUBS 0.01732f
C40 B.n12 VSUBS 0.006881f
C41 B.n13 VSUBS 0.006881f
C42 B.n14 VSUBS 0.006881f
C43 B.n15 VSUBS 0.006881f
C44 B.n16 VSUBS 0.006881f
C45 B.n17 VSUBS 0.006881f
C46 B.n18 VSUBS 0.006881f
C47 B.n19 VSUBS 0.006881f
C48 B.n20 VSUBS 0.006881f
C49 B.n21 VSUBS 0.006881f
C50 B.n22 VSUBS 0.004756f
C51 B.n23 VSUBS 0.006881f
C52 B.t8 VSUBS 0.076301f
C53 B.t7 VSUBS 0.084537f
C54 B.t6 VSUBS 0.139869f
C55 B.n24 VSUBS 0.149881f
C56 B.n25 VSUBS 0.132496f
C57 B.n26 VSUBS 0.015942f
C58 B.n27 VSUBS 0.006881f
C59 B.n28 VSUBS 0.006881f
C60 B.n29 VSUBS 0.006881f
C61 B.n30 VSUBS 0.006881f
C62 B.t11 VSUBS 0.076302f
C63 B.t10 VSUBS 0.084538f
C64 B.t9 VSUBS 0.139869f
C65 B.n31 VSUBS 0.14988f
C66 B.n32 VSUBS 0.132494f
C67 B.n33 VSUBS 0.006881f
C68 B.n34 VSUBS 0.006881f
C69 B.n35 VSUBS 0.006881f
C70 B.n36 VSUBS 0.006881f
C71 B.n37 VSUBS 0.006881f
C72 B.n38 VSUBS 0.006881f
C73 B.n39 VSUBS 0.006881f
C74 B.n40 VSUBS 0.006881f
C75 B.n41 VSUBS 0.006881f
C76 B.n42 VSUBS 0.006881f
C77 B.n43 VSUBS 0.018026f
C78 B.n44 VSUBS 0.006881f
C79 B.n45 VSUBS 0.006881f
C80 B.n46 VSUBS 0.006881f
C81 B.n47 VSUBS 0.006881f
C82 B.n48 VSUBS 0.006881f
C83 B.n49 VSUBS 0.006881f
C84 B.n50 VSUBS 0.006881f
C85 B.n51 VSUBS 0.006881f
C86 B.n52 VSUBS 0.006881f
C87 B.n53 VSUBS 0.006881f
C88 B.n54 VSUBS 0.006881f
C89 B.n55 VSUBS 0.006881f
C90 B.n56 VSUBS 0.006881f
C91 B.n57 VSUBS 0.006881f
C92 B.n58 VSUBS 0.006881f
C93 B.n59 VSUBS 0.006881f
C94 B.n60 VSUBS 0.006881f
C95 B.n61 VSUBS 0.006881f
C96 B.n62 VSUBS 0.01732f
C97 B.n63 VSUBS 0.006881f
C98 B.n64 VSUBS 0.006881f
C99 B.n65 VSUBS 0.006881f
C100 B.n66 VSUBS 0.006881f
C101 B.n67 VSUBS 0.006881f
C102 B.n68 VSUBS 0.006881f
C103 B.n69 VSUBS 0.006881f
C104 B.n70 VSUBS 0.006881f
C105 B.n71 VSUBS 0.006881f
C106 B.n72 VSUBS 0.006881f
C107 B.n73 VSUBS 0.004756f
C108 B.n74 VSUBS 0.006881f
C109 B.n75 VSUBS 0.006881f
C110 B.n76 VSUBS 0.006881f
C111 B.n77 VSUBS 0.006881f
C112 B.n78 VSUBS 0.006881f
C113 B.t4 VSUBS 0.076301f
C114 B.t5 VSUBS 0.084537f
C115 B.t3 VSUBS 0.139869f
C116 B.n79 VSUBS 0.149881f
C117 B.n80 VSUBS 0.132496f
C118 B.n81 VSUBS 0.006881f
C119 B.n82 VSUBS 0.006881f
C120 B.n83 VSUBS 0.006881f
C121 B.n84 VSUBS 0.006881f
C122 B.n85 VSUBS 0.006881f
C123 B.n86 VSUBS 0.006881f
C124 B.n87 VSUBS 0.006881f
C125 B.n88 VSUBS 0.006881f
C126 B.n89 VSUBS 0.006881f
C127 B.n90 VSUBS 0.006881f
C128 B.n91 VSUBS 0.01732f
C129 B.n92 VSUBS 0.006881f
C130 B.n93 VSUBS 0.006881f
C131 B.n94 VSUBS 0.006881f
C132 B.n95 VSUBS 0.006881f
C133 B.n96 VSUBS 0.006881f
C134 B.n97 VSUBS 0.006881f
C135 B.n98 VSUBS 0.006881f
C136 B.n99 VSUBS 0.006881f
C137 B.n100 VSUBS 0.006881f
C138 B.n101 VSUBS 0.006881f
C139 B.n102 VSUBS 0.006881f
C140 B.n103 VSUBS 0.006881f
C141 B.n104 VSUBS 0.006881f
C142 B.n105 VSUBS 0.006881f
C143 B.n106 VSUBS 0.006881f
C144 B.n107 VSUBS 0.006881f
C145 B.n108 VSUBS 0.006881f
C146 B.n109 VSUBS 0.006881f
C147 B.n110 VSUBS 0.006881f
C148 B.n111 VSUBS 0.006881f
C149 B.n112 VSUBS 0.006881f
C150 B.n113 VSUBS 0.006881f
C151 B.n114 VSUBS 0.006881f
C152 B.n115 VSUBS 0.006881f
C153 B.n116 VSUBS 0.006881f
C154 B.n117 VSUBS 0.006881f
C155 B.n118 VSUBS 0.006881f
C156 B.n119 VSUBS 0.006881f
C157 B.n120 VSUBS 0.006881f
C158 B.n121 VSUBS 0.006881f
C159 B.n122 VSUBS 0.006881f
C160 B.n123 VSUBS 0.006881f
C161 B.n124 VSUBS 0.006881f
C162 B.n125 VSUBS 0.006881f
C163 B.n126 VSUBS 0.01732f
C164 B.n127 VSUBS 0.018095f
C165 B.n128 VSUBS 0.018095f
C166 B.n129 VSUBS 0.006881f
C167 B.n130 VSUBS 0.006881f
C168 B.n131 VSUBS 0.006881f
C169 B.n132 VSUBS 0.006881f
C170 B.n133 VSUBS 0.006881f
C171 B.n134 VSUBS 0.006881f
C172 B.n135 VSUBS 0.006881f
C173 B.n136 VSUBS 0.006881f
C174 B.n137 VSUBS 0.006881f
C175 B.n138 VSUBS 0.006881f
C176 B.n139 VSUBS 0.006881f
C177 B.n140 VSUBS 0.006881f
C178 B.n141 VSUBS 0.006881f
C179 B.n142 VSUBS 0.006881f
C180 B.n143 VSUBS 0.006881f
C181 B.n144 VSUBS 0.006881f
C182 B.n145 VSUBS 0.006881f
C183 B.n146 VSUBS 0.006881f
C184 B.n147 VSUBS 0.006881f
C185 B.n148 VSUBS 0.006881f
C186 B.n149 VSUBS 0.006881f
C187 B.n150 VSUBS 0.006881f
C188 B.n151 VSUBS 0.006881f
C189 B.n152 VSUBS 0.006881f
C190 B.n153 VSUBS 0.006881f
C191 B.n154 VSUBS 0.006881f
C192 B.n155 VSUBS 0.006881f
C193 B.n156 VSUBS 0.006881f
C194 B.n157 VSUBS 0.006881f
C195 B.n158 VSUBS 0.006881f
C196 B.n159 VSUBS 0.004756f
C197 B.n160 VSUBS 0.015942f
C198 B.n161 VSUBS 0.005565f
C199 B.n162 VSUBS 0.006881f
C200 B.n163 VSUBS 0.006881f
C201 B.n164 VSUBS 0.006881f
C202 B.n165 VSUBS 0.006881f
C203 B.n166 VSUBS 0.006881f
C204 B.n167 VSUBS 0.006881f
C205 B.n168 VSUBS 0.006881f
C206 B.n169 VSUBS 0.006881f
C207 B.n170 VSUBS 0.006881f
C208 B.n171 VSUBS 0.006881f
C209 B.n172 VSUBS 0.006881f
C210 B.t1 VSUBS 0.076302f
C211 B.t2 VSUBS 0.084538f
C212 B.t0 VSUBS 0.139869f
C213 B.n173 VSUBS 0.14988f
C214 B.n174 VSUBS 0.132494f
C215 B.n175 VSUBS 0.015942f
C216 B.n176 VSUBS 0.005565f
C217 B.n177 VSUBS 0.006881f
C218 B.n178 VSUBS 0.006881f
C219 B.n179 VSUBS 0.006881f
C220 B.n180 VSUBS 0.006881f
C221 B.n181 VSUBS 0.006881f
C222 B.n182 VSUBS 0.006881f
C223 B.n183 VSUBS 0.006881f
C224 B.n184 VSUBS 0.006881f
C225 B.n185 VSUBS 0.006881f
C226 B.n186 VSUBS 0.006881f
C227 B.n187 VSUBS 0.006881f
C228 B.n188 VSUBS 0.006881f
C229 B.n189 VSUBS 0.006881f
C230 B.n190 VSUBS 0.006881f
C231 B.n191 VSUBS 0.006881f
C232 B.n192 VSUBS 0.006881f
C233 B.n193 VSUBS 0.006881f
C234 B.n194 VSUBS 0.006881f
C235 B.n195 VSUBS 0.006881f
C236 B.n196 VSUBS 0.006881f
C237 B.n197 VSUBS 0.006881f
C238 B.n198 VSUBS 0.006881f
C239 B.n199 VSUBS 0.006881f
C240 B.n200 VSUBS 0.006881f
C241 B.n201 VSUBS 0.006881f
C242 B.n202 VSUBS 0.006881f
C243 B.n203 VSUBS 0.006881f
C244 B.n204 VSUBS 0.006881f
C245 B.n205 VSUBS 0.006881f
C246 B.n206 VSUBS 0.006881f
C247 B.n207 VSUBS 0.006881f
C248 B.n208 VSUBS 0.006881f
C249 B.n209 VSUBS 0.018095f
C250 B.n210 VSUBS 0.018095f
C251 B.n211 VSUBS 0.01732f
C252 B.n212 VSUBS 0.006881f
C253 B.n213 VSUBS 0.006881f
C254 B.n214 VSUBS 0.006881f
C255 B.n215 VSUBS 0.006881f
C256 B.n216 VSUBS 0.006881f
C257 B.n217 VSUBS 0.006881f
C258 B.n218 VSUBS 0.006881f
C259 B.n219 VSUBS 0.006881f
C260 B.n220 VSUBS 0.006881f
C261 B.n221 VSUBS 0.006881f
C262 B.n222 VSUBS 0.006881f
C263 B.n223 VSUBS 0.006881f
C264 B.n224 VSUBS 0.006881f
C265 B.n225 VSUBS 0.006881f
C266 B.n226 VSUBS 0.006881f
C267 B.n227 VSUBS 0.006881f
C268 B.n228 VSUBS 0.006881f
C269 B.n229 VSUBS 0.006881f
C270 B.n230 VSUBS 0.006881f
C271 B.n231 VSUBS 0.006881f
C272 B.n232 VSUBS 0.006881f
C273 B.n233 VSUBS 0.006881f
C274 B.n234 VSUBS 0.006881f
C275 B.n235 VSUBS 0.006881f
C276 B.n236 VSUBS 0.006881f
C277 B.n237 VSUBS 0.006881f
C278 B.n238 VSUBS 0.006881f
C279 B.n239 VSUBS 0.006881f
C280 B.n240 VSUBS 0.006881f
C281 B.n241 VSUBS 0.006881f
C282 B.n242 VSUBS 0.006881f
C283 B.n243 VSUBS 0.006881f
C284 B.n244 VSUBS 0.006881f
C285 B.n245 VSUBS 0.006881f
C286 B.n246 VSUBS 0.006881f
C287 B.n247 VSUBS 0.006881f
C288 B.n248 VSUBS 0.006881f
C289 B.n249 VSUBS 0.006881f
C290 B.n250 VSUBS 0.006881f
C291 B.n251 VSUBS 0.006881f
C292 B.n252 VSUBS 0.006881f
C293 B.n253 VSUBS 0.006881f
C294 B.n254 VSUBS 0.006881f
C295 B.n255 VSUBS 0.006881f
C296 B.n256 VSUBS 0.006881f
C297 B.n257 VSUBS 0.006881f
C298 B.n258 VSUBS 0.006881f
C299 B.n259 VSUBS 0.006881f
C300 B.n260 VSUBS 0.006881f
C301 B.n261 VSUBS 0.006881f
C302 B.n262 VSUBS 0.006881f
C303 B.n263 VSUBS 0.006881f
C304 B.n264 VSUBS 0.006881f
C305 B.n265 VSUBS 0.006881f
C306 B.n266 VSUBS 0.006881f
C307 B.n267 VSUBS 0.006881f
C308 B.n268 VSUBS 0.01732f
C309 B.n269 VSUBS 0.018095f
C310 B.n270 VSUBS 0.017389f
C311 B.n271 VSUBS 0.006881f
C312 B.n272 VSUBS 0.006881f
C313 B.n273 VSUBS 0.006881f
C314 B.n274 VSUBS 0.006881f
C315 B.n275 VSUBS 0.006881f
C316 B.n276 VSUBS 0.006881f
C317 B.n277 VSUBS 0.006881f
C318 B.n278 VSUBS 0.006881f
C319 B.n279 VSUBS 0.006881f
C320 B.n280 VSUBS 0.006881f
C321 B.n281 VSUBS 0.006881f
C322 B.n282 VSUBS 0.006881f
C323 B.n283 VSUBS 0.006881f
C324 B.n284 VSUBS 0.006881f
C325 B.n285 VSUBS 0.006881f
C326 B.n286 VSUBS 0.006881f
C327 B.n287 VSUBS 0.006881f
C328 B.n288 VSUBS 0.006881f
C329 B.n289 VSUBS 0.006881f
C330 B.n290 VSUBS 0.006881f
C331 B.n291 VSUBS 0.006881f
C332 B.n292 VSUBS 0.006881f
C333 B.n293 VSUBS 0.006881f
C334 B.n294 VSUBS 0.006881f
C335 B.n295 VSUBS 0.006881f
C336 B.n296 VSUBS 0.006881f
C337 B.n297 VSUBS 0.006881f
C338 B.n298 VSUBS 0.006881f
C339 B.n299 VSUBS 0.006881f
C340 B.n300 VSUBS 0.006881f
C341 B.n301 VSUBS 0.004756f
C342 B.n302 VSUBS 0.015942f
C343 B.n303 VSUBS 0.005565f
C344 B.n304 VSUBS 0.006881f
C345 B.n305 VSUBS 0.006881f
C346 B.n306 VSUBS 0.006881f
C347 B.n307 VSUBS 0.006881f
C348 B.n308 VSUBS 0.006881f
C349 B.n309 VSUBS 0.006881f
C350 B.n310 VSUBS 0.006881f
C351 B.n311 VSUBS 0.006881f
C352 B.n312 VSUBS 0.006881f
C353 B.n313 VSUBS 0.006881f
C354 B.n314 VSUBS 0.006881f
C355 B.n315 VSUBS 0.005565f
C356 B.n316 VSUBS 0.006881f
C357 B.n317 VSUBS 0.006881f
C358 B.n318 VSUBS 0.006881f
C359 B.n319 VSUBS 0.006881f
C360 B.n320 VSUBS 0.006881f
C361 B.n321 VSUBS 0.006881f
C362 B.n322 VSUBS 0.006881f
C363 B.n323 VSUBS 0.006881f
C364 B.n324 VSUBS 0.006881f
C365 B.n325 VSUBS 0.006881f
C366 B.n326 VSUBS 0.006881f
C367 B.n327 VSUBS 0.006881f
C368 B.n328 VSUBS 0.006881f
C369 B.n329 VSUBS 0.006881f
C370 B.n330 VSUBS 0.006881f
C371 B.n331 VSUBS 0.006881f
C372 B.n332 VSUBS 0.006881f
C373 B.n333 VSUBS 0.006881f
C374 B.n334 VSUBS 0.006881f
C375 B.n335 VSUBS 0.006881f
C376 B.n336 VSUBS 0.006881f
C377 B.n337 VSUBS 0.006881f
C378 B.n338 VSUBS 0.006881f
C379 B.n339 VSUBS 0.006881f
C380 B.n340 VSUBS 0.006881f
C381 B.n341 VSUBS 0.006881f
C382 B.n342 VSUBS 0.006881f
C383 B.n343 VSUBS 0.006881f
C384 B.n344 VSUBS 0.006881f
C385 B.n345 VSUBS 0.006881f
C386 B.n346 VSUBS 0.006881f
C387 B.n347 VSUBS 0.006881f
C388 B.n348 VSUBS 0.018095f
C389 B.n349 VSUBS 0.018095f
C390 B.n350 VSUBS 0.01732f
C391 B.n351 VSUBS 0.006881f
C392 B.n352 VSUBS 0.006881f
C393 B.n353 VSUBS 0.006881f
C394 B.n354 VSUBS 0.006881f
C395 B.n355 VSUBS 0.006881f
C396 B.n356 VSUBS 0.006881f
C397 B.n357 VSUBS 0.006881f
C398 B.n358 VSUBS 0.006881f
C399 B.n359 VSUBS 0.006881f
C400 B.n360 VSUBS 0.006881f
C401 B.n361 VSUBS 0.006881f
C402 B.n362 VSUBS 0.006881f
C403 B.n363 VSUBS 0.006881f
C404 B.n364 VSUBS 0.006881f
C405 B.n365 VSUBS 0.006881f
C406 B.n366 VSUBS 0.006881f
C407 B.n367 VSUBS 0.006881f
C408 B.n368 VSUBS 0.006881f
C409 B.n369 VSUBS 0.006881f
C410 B.n370 VSUBS 0.006881f
C411 B.n371 VSUBS 0.006881f
C412 B.n372 VSUBS 0.006881f
C413 B.n373 VSUBS 0.006881f
C414 B.n374 VSUBS 0.006881f
C415 B.n375 VSUBS 0.006881f
C416 B.n376 VSUBS 0.006881f
C417 B.n377 VSUBS 0.006881f
C418 B.n378 VSUBS 0.006881f
C419 B.n379 VSUBS 0.01558f
C420 VDD1.n0 VSUBS 0.025797f
C421 VDD1.n1 VSUBS 0.023752f
C422 VDD1.n2 VSUBS 0.012763f
C423 VDD1.n3 VSUBS 0.030168f
C424 VDD1.n4 VSUBS 0.013514f
C425 VDD1.n5 VSUBS 0.023752f
C426 VDD1.n6 VSUBS 0.012763f
C427 VDD1.n7 VSUBS 0.022626f
C428 VDD1.n8 VSUBS 0.019163f
C429 VDD1.t5 VSUBS 0.065095f
C430 VDD1.n9 VSUBS 0.100452f
C431 VDD1.n10 VSUBS 0.468648f
C432 VDD1.n11 VSUBS 0.012763f
C433 VDD1.n12 VSUBS 0.013514f
C434 VDD1.n13 VSUBS 0.030168f
C435 VDD1.n14 VSUBS 0.030168f
C436 VDD1.n15 VSUBS 0.013514f
C437 VDD1.n16 VSUBS 0.012763f
C438 VDD1.n17 VSUBS 0.023752f
C439 VDD1.n18 VSUBS 0.023752f
C440 VDD1.n19 VSUBS 0.012763f
C441 VDD1.n20 VSUBS 0.013514f
C442 VDD1.n21 VSUBS 0.030168f
C443 VDD1.n22 VSUBS 0.072008f
C444 VDD1.n23 VSUBS 0.013514f
C445 VDD1.n24 VSUBS 0.012763f
C446 VDD1.n25 VSUBS 0.05555f
C447 VDD1.n26 VSUBS 0.053896f
C448 VDD1.n27 VSUBS 0.025797f
C449 VDD1.n28 VSUBS 0.023752f
C450 VDD1.n29 VSUBS 0.012763f
C451 VDD1.n30 VSUBS 0.030168f
C452 VDD1.n31 VSUBS 0.013514f
C453 VDD1.n32 VSUBS 0.023752f
C454 VDD1.n33 VSUBS 0.012763f
C455 VDD1.n34 VSUBS 0.022626f
C456 VDD1.n35 VSUBS 0.019163f
C457 VDD1.t0 VSUBS 0.065095f
C458 VDD1.n36 VSUBS 0.100452f
C459 VDD1.n37 VSUBS 0.468648f
C460 VDD1.n38 VSUBS 0.012763f
C461 VDD1.n39 VSUBS 0.013514f
C462 VDD1.n40 VSUBS 0.030168f
C463 VDD1.n41 VSUBS 0.030168f
C464 VDD1.n42 VSUBS 0.013514f
C465 VDD1.n43 VSUBS 0.012763f
C466 VDD1.n44 VSUBS 0.023752f
C467 VDD1.n45 VSUBS 0.023752f
C468 VDD1.n46 VSUBS 0.012763f
C469 VDD1.n47 VSUBS 0.013514f
C470 VDD1.n48 VSUBS 0.030168f
C471 VDD1.n49 VSUBS 0.072008f
C472 VDD1.n50 VSUBS 0.013514f
C473 VDD1.n51 VSUBS 0.012763f
C474 VDD1.n52 VSUBS 0.05555f
C475 VDD1.n53 VSUBS 0.05359f
C476 VDD1.t1 VSUBS 0.099478f
C477 VDD1.t3 VSUBS 0.099478f
C478 VDD1.n54 VSUBS 0.636868f
C479 VDD1.n55 VSUBS 1.59501f
C480 VDD1.t2 VSUBS 0.099478f
C481 VDD1.t4 VSUBS 0.099478f
C482 VDD1.n56 VSUBS 0.636168f
C483 VDD1.n57 VSUBS 1.7893f
C484 VP.n0 VSUBS 0.075147f
C485 VP.t0 VSUBS 0.564067f
C486 VP.n1 VSUBS 0.238534f
C487 VP.t1 VSUBS 0.540423f
C488 VP.t3 VSUBS 0.540423f
C489 VP.n2 VSUBS 0.273762f
C490 VP.n3 VSUBS 0.260952f
C491 VP.n4 VSUBS 1.95351f
C492 VP.n5 VSUBS 1.84282f
C493 VP.t5 VSUBS 0.540423f
C494 VP.n6 VSUBS 0.260952f
C495 VP.t4 VSUBS 0.540423f
C496 VP.n7 VSUBS 0.273762f
C497 VP.t2 VSUBS 0.540423f
C498 VP.n8 VSUBS 0.260952f
C499 VP.n9 VSUBS 0.06262f
C500 VTAIL.t10 VSUBS 0.08244f
C501 VTAIL.t8 VSUBS 0.08244f
C502 VTAIL.n0 VSUBS 0.464737f
C503 VTAIL.n1 VSUBS 0.415477f
C504 VTAIL.n2 VSUBS 0.021379f
C505 VTAIL.n3 VSUBS 0.019684f
C506 VTAIL.n4 VSUBS 0.010577f
C507 VTAIL.n5 VSUBS 0.025001f
C508 VTAIL.n6 VSUBS 0.0112f
C509 VTAIL.n7 VSUBS 0.019684f
C510 VTAIL.n8 VSUBS 0.010577f
C511 VTAIL.n9 VSUBS 0.018751f
C512 VTAIL.n10 VSUBS 0.015881f
C513 VTAIL.t4 VSUBS 0.053946f
C514 VTAIL.n11 VSUBS 0.083248f
C515 VTAIL.n12 VSUBS 0.388384f
C516 VTAIL.n13 VSUBS 0.010577f
C517 VTAIL.n14 VSUBS 0.0112f
C518 VTAIL.n15 VSUBS 0.025001f
C519 VTAIL.n16 VSUBS 0.025001f
C520 VTAIL.n17 VSUBS 0.0112f
C521 VTAIL.n18 VSUBS 0.010577f
C522 VTAIL.n19 VSUBS 0.019684f
C523 VTAIL.n20 VSUBS 0.019684f
C524 VTAIL.n21 VSUBS 0.010577f
C525 VTAIL.n22 VSUBS 0.0112f
C526 VTAIL.n23 VSUBS 0.025001f
C527 VTAIL.n24 VSUBS 0.059675f
C528 VTAIL.n25 VSUBS 0.0112f
C529 VTAIL.n26 VSUBS 0.010577f
C530 VTAIL.n27 VSUBS 0.046036f
C531 VTAIL.n28 VSUBS 0.029989f
C532 VTAIL.n29 VSUBS 0.12483f
C533 VTAIL.t1 VSUBS 0.08244f
C534 VTAIL.t0 VSUBS 0.08244f
C535 VTAIL.n30 VSUBS 0.464737f
C536 VTAIL.n31 VSUBS 1.05603f
C537 VTAIL.t6 VSUBS 0.08244f
C538 VTAIL.t11 VSUBS 0.08244f
C539 VTAIL.n32 VSUBS 0.46474f
C540 VTAIL.n33 VSUBS 1.05603f
C541 VTAIL.n34 VSUBS 0.021379f
C542 VTAIL.n35 VSUBS 0.019684f
C543 VTAIL.n36 VSUBS 0.010577f
C544 VTAIL.n37 VSUBS 0.025001f
C545 VTAIL.n38 VSUBS 0.0112f
C546 VTAIL.n39 VSUBS 0.019684f
C547 VTAIL.n40 VSUBS 0.010577f
C548 VTAIL.n41 VSUBS 0.018751f
C549 VTAIL.n42 VSUBS 0.015881f
C550 VTAIL.t9 VSUBS 0.053946f
C551 VTAIL.n43 VSUBS 0.083248f
C552 VTAIL.n44 VSUBS 0.388384f
C553 VTAIL.n45 VSUBS 0.010577f
C554 VTAIL.n46 VSUBS 0.0112f
C555 VTAIL.n47 VSUBS 0.025001f
C556 VTAIL.n48 VSUBS 0.025001f
C557 VTAIL.n49 VSUBS 0.0112f
C558 VTAIL.n50 VSUBS 0.010577f
C559 VTAIL.n51 VSUBS 0.019684f
C560 VTAIL.n52 VSUBS 0.019684f
C561 VTAIL.n53 VSUBS 0.010577f
C562 VTAIL.n54 VSUBS 0.0112f
C563 VTAIL.n55 VSUBS 0.025001f
C564 VTAIL.n56 VSUBS 0.059675f
C565 VTAIL.n57 VSUBS 0.0112f
C566 VTAIL.n58 VSUBS 0.010577f
C567 VTAIL.n59 VSUBS 0.046036f
C568 VTAIL.n60 VSUBS 0.029989f
C569 VTAIL.n61 VSUBS 0.12483f
C570 VTAIL.t5 VSUBS 0.08244f
C571 VTAIL.t3 VSUBS 0.08244f
C572 VTAIL.n62 VSUBS 0.46474f
C573 VTAIL.n63 VSUBS 0.450741f
C574 VTAIL.n64 VSUBS 0.021379f
C575 VTAIL.n65 VSUBS 0.019684f
C576 VTAIL.n66 VSUBS 0.010577f
C577 VTAIL.n67 VSUBS 0.025001f
C578 VTAIL.n68 VSUBS 0.0112f
C579 VTAIL.n69 VSUBS 0.019684f
C580 VTAIL.n70 VSUBS 0.010577f
C581 VTAIL.n71 VSUBS 0.018751f
C582 VTAIL.n72 VSUBS 0.015881f
C583 VTAIL.t2 VSUBS 0.053946f
C584 VTAIL.n73 VSUBS 0.083248f
C585 VTAIL.n74 VSUBS 0.388384f
C586 VTAIL.n75 VSUBS 0.010577f
C587 VTAIL.n76 VSUBS 0.0112f
C588 VTAIL.n77 VSUBS 0.025001f
C589 VTAIL.n78 VSUBS 0.025001f
C590 VTAIL.n79 VSUBS 0.0112f
C591 VTAIL.n80 VSUBS 0.010577f
C592 VTAIL.n81 VSUBS 0.019684f
C593 VTAIL.n82 VSUBS 0.019684f
C594 VTAIL.n83 VSUBS 0.010577f
C595 VTAIL.n84 VSUBS 0.0112f
C596 VTAIL.n85 VSUBS 0.025001f
C597 VTAIL.n86 VSUBS 0.059675f
C598 VTAIL.n87 VSUBS 0.0112f
C599 VTAIL.n88 VSUBS 0.010577f
C600 VTAIL.n89 VSUBS 0.046036f
C601 VTAIL.n90 VSUBS 0.029989f
C602 VTAIL.n91 VSUBS 0.678176f
C603 VTAIL.n92 VSUBS 0.021379f
C604 VTAIL.n93 VSUBS 0.019684f
C605 VTAIL.n94 VSUBS 0.010577f
C606 VTAIL.n95 VSUBS 0.025001f
C607 VTAIL.n96 VSUBS 0.0112f
C608 VTAIL.n97 VSUBS 0.019684f
C609 VTAIL.n98 VSUBS 0.010577f
C610 VTAIL.n99 VSUBS 0.018751f
C611 VTAIL.n100 VSUBS 0.015881f
C612 VTAIL.t7 VSUBS 0.053946f
C613 VTAIL.n101 VSUBS 0.083248f
C614 VTAIL.n102 VSUBS 0.388384f
C615 VTAIL.n103 VSUBS 0.010577f
C616 VTAIL.n104 VSUBS 0.0112f
C617 VTAIL.n105 VSUBS 0.025001f
C618 VTAIL.n106 VSUBS 0.025001f
C619 VTAIL.n107 VSUBS 0.0112f
C620 VTAIL.n108 VSUBS 0.010577f
C621 VTAIL.n109 VSUBS 0.019684f
C622 VTAIL.n110 VSUBS 0.019684f
C623 VTAIL.n111 VSUBS 0.010577f
C624 VTAIL.n112 VSUBS 0.0112f
C625 VTAIL.n113 VSUBS 0.025001f
C626 VTAIL.n114 VSUBS 0.059675f
C627 VTAIL.n115 VSUBS 0.0112f
C628 VTAIL.n116 VSUBS 0.010577f
C629 VTAIL.n117 VSUBS 0.046036f
C630 VTAIL.n118 VSUBS 0.029989f
C631 VTAIL.n119 VSUBS 0.661499f
C632 VDD2.n0 VSUBS 0.018978f
C633 VDD2.n1 VSUBS 0.017473f
C634 VDD2.n2 VSUBS 0.009389f
C635 VDD2.n3 VSUBS 0.022193f
C636 VDD2.n4 VSUBS 0.009942f
C637 VDD2.n5 VSUBS 0.017473f
C638 VDD2.n6 VSUBS 0.009389f
C639 VDD2.n7 VSUBS 0.016645f
C640 VDD2.n8 VSUBS 0.014097f
C641 VDD2.t0 VSUBS 0.047888f
C642 VDD2.n9 VSUBS 0.073898f
C643 VDD2.n10 VSUBS 0.344763f
C644 VDD2.n11 VSUBS 0.009389f
C645 VDD2.n12 VSUBS 0.009942f
C646 VDD2.n13 VSUBS 0.022193f
C647 VDD2.n14 VSUBS 0.022193f
C648 VDD2.n15 VSUBS 0.009942f
C649 VDD2.n16 VSUBS 0.009389f
C650 VDD2.n17 VSUBS 0.017473f
C651 VDD2.n18 VSUBS 0.017473f
C652 VDD2.n19 VSUBS 0.009389f
C653 VDD2.n20 VSUBS 0.009942f
C654 VDD2.n21 VSUBS 0.022193f
C655 VDD2.n22 VSUBS 0.052973f
C656 VDD2.n23 VSUBS 0.009942f
C657 VDD2.n24 VSUBS 0.009389f
C658 VDD2.n25 VSUBS 0.040866f
C659 VDD2.n26 VSUBS 0.039424f
C660 VDD2.t1 VSUBS 0.073181f
C661 VDD2.t4 VSUBS 0.073181f
C662 VDD2.n27 VSUBS 0.468514f
C663 VDD2.n28 VSUBS 1.12266f
C664 VDD2.n29 VSUBS 0.018978f
C665 VDD2.n30 VSUBS 0.017473f
C666 VDD2.n31 VSUBS 0.009389f
C667 VDD2.n32 VSUBS 0.022193f
C668 VDD2.n33 VSUBS 0.009942f
C669 VDD2.n34 VSUBS 0.017473f
C670 VDD2.n35 VSUBS 0.009389f
C671 VDD2.n36 VSUBS 0.016645f
C672 VDD2.n37 VSUBS 0.014097f
C673 VDD2.t5 VSUBS 0.047888f
C674 VDD2.n38 VSUBS 0.073898f
C675 VDD2.n39 VSUBS 0.344763f
C676 VDD2.n40 VSUBS 0.009389f
C677 VDD2.n41 VSUBS 0.009942f
C678 VDD2.n42 VSUBS 0.022193f
C679 VDD2.n43 VSUBS 0.022193f
C680 VDD2.n44 VSUBS 0.009942f
C681 VDD2.n45 VSUBS 0.009389f
C682 VDD2.n46 VSUBS 0.017473f
C683 VDD2.n47 VSUBS 0.017473f
C684 VDD2.n48 VSUBS 0.009389f
C685 VDD2.n49 VSUBS 0.009942f
C686 VDD2.n50 VSUBS 0.022193f
C687 VDD2.n51 VSUBS 0.052973f
C688 VDD2.n52 VSUBS 0.009942f
C689 VDD2.n53 VSUBS 0.009389f
C690 VDD2.n54 VSUBS 0.040866f
C691 VDD2.n55 VSUBS 0.038682f
C692 VDD2.n56 VSUBS 1.04006f
C693 VDD2.t3 VSUBS 0.073181f
C694 VDD2.t2 VSUBS 0.073181f
C695 VDD2.n57 VSUBS 0.4685f
C696 VN.t1 VSUBS 0.412917f
C697 VN.n0 VSUBS 0.174615f
C698 VN.t3 VSUBS 0.395609f
C699 VN.n1 VSUBS 0.200403f
C700 VN.t4 VSUBS 0.395609f
C701 VN.n2 VSUBS 0.191027f
C702 VN.n3 VSUBS 0.16834f
C703 VN.t2 VSUBS 0.412917f
C704 VN.n4 VSUBS 0.174615f
C705 VN.t0 VSUBS 0.395609f
C706 VN.n5 VSUBS 0.200403f
C707 VN.t5 VSUBS 0.395609f
C708 VN.n6 VSUBS 0.191027f
C709 VN.n7 VSUBS 1.45745f
.ends

