* NGSPICE file created from diff_pair_sample_1107.ext - technology: sky130A

.subckt diff_pair_sample_1107 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t3 VP.t0 VTAIL.t4 B.t0 sky130_fd_pr__nfet_01v8 ad=0.4719 pd=3.19 as=1.1154 ps=6.5 w=2.86 l=1.1
X1 B.t17 B.t15 B.t16 B.t9 sky130_fd_pr__nfet_01v8 ad=1.1154 pd=6.5 as=0 ps=0 w=2.86 l=1.1
X2 VTAIL.t6 VP.t1 VDD1.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.1154 pd=6.5 as=0.4719 ps=3.19 w=2.86 l=1.1
X3 B.t14 B.t12 B.t13 B.t5 sky130_fd_pr__nfet_01v8 ad=1.1154 pd=6.5 as=0 ps=0 w=2.86 l=1.1
X4 VTAIL.t2 VN.t0 VDD2.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=1.1154 pd=6.5 as=0.4719 ps=3.19 w=2.86 l=1.1
X5 VDD2.t2 VN.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.4719 pd=3.19 as=1.1154 ps=6.5 w=2.86 l=1.1
X6 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=1.1154 pd=6.5 as=0 ps=0 w=2.86 l=1.1
X7 VTAIL.t5 VP.t2 VDD1.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=1.1154 pd=6.5 as=0.4719 ps=3.19 w=2.86 l=1.1
X8 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=1.1154 pd=6.5 as=0 ps=0 w=2.86 l=1.1
X9 VDD2.t1 VN.t2 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.4719 pd=3.19 as=1.1154 ps=6.5 w=2.86 l=1.1
X10 VDD1.t0 VP.t3 VTAIL.t7 B.t1 sky130_fd_pr__nfet_01v8 ad=0.4719 pd=3.19 as=1.1154 ps=6.5 w=2.86 l=1.1
X11 VTAIL.t3 VN.t3 VDD2.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=1.1154 pd=6.5 as=0.4719 ps=3.19 w=2.86 l=1.1
R0 VP.n0 VP.t2 116.98
R1 VP.n0 VP.t0 116.892
R2 VP.n2 VP.t1 98.3723
R3 VP.n3 VP.t3 98.3723
R4 VP.n4 VP.n3 80.6037
R5 VP.n2 VP.n1 80.6037
R6 VP.n1 VP.n0 66.1168
R7 VP.n3 VP.n2 48.2005
R8 VP.n4 VP.n1 0.380177
R9 VP VP.n4 0.146778
R10 VTAIL.n5 VTAIL.t5 73.0123
R11 VTAIL.n4 VTAIL.t1 73.0123
R12 VTAIL.n3 VTAIL.t2 73.0123
R13 VTAIL.n7 VTAIL.t0 73.012
R14 VTAIL.n0 VTAIL.t3 73.012
R15 VTAIL.n1 VTAIL.t7 73.012
R16 VTAIL.n2 VTAIL.t6 73.012
R17 VTAIL.n6 VTAIL.t4 73.012
R18 VTAIL.n7 VTAIL.n6 16.0652
R19 VTAIL.n3 VTAIL.n2 16.0652
R20 VTAIL.n4 VTAIL.n3 1.23326
R21 VTAIL.n6 VTAIL.n5 1.23326
R22 VTAIL.n2 VTAIL.n1 1.23326
R23 VTAIL VTAIL.n0 0.675069
R24 VTAIL VTAIL.n7 0.55869
R25 VTAIL.n5 VTAIL.n4 0.470328
R26 VTAIL.n1 VTAIL.n0 0.470328
R27 VDD1 VDD1.n1 113.171
R28 VDD1 VDD1.n0 82.8261
R29 VDD1.n0 VDD1.t1 6.92358
R30 VDD1.n0 VDD1.t3 6.92358
R31 VDD1.n1 VDD1.t2 6.92358
R32 VDD1.n1 VDD1.t0 6.92358
R33 B.n371 B.n370 585
R34 B.n372 B.n371 585
R35 B.n139 B.n60 585
R36 B.n138 B.n137 585
R37 B.n136 B.n135 585
R38 B.n134 B.n133 585
R39 B.n132 B.n131 585
R40 B.n130 B.n129 585
R41 B.n128 B.n127 585
R42 B.n126 B.n125 585
R43 B.n124 B.n123 585
R44 B.n122 B.n121 585
R45 B.n120 B.n119 585
R46 B.n118 B.n117 585
R47 B.n116 B.n115 585
R48 B.n114 B.n113 585
R49 B.n112 B.n111 585
R50 B.n110 B.n109 585
R51 B.n108 B.n107 585
R52 B.n106 B.n105 585
R53 B.n104 B.n103 585
R54 B.n102 B.n101 585
R55 B.n100 B.n99 585
R56 B.n98 B.n97 585
R57 B.n96 B.n95 585
R58 B.n93 B.n92 585
R59 B.n91 B.n90 585
R60 B.n89 B.n88 585
R61 B.n87 B.n86 585
R62 B.n85 B.n84 585
R63 B.n83 B.n82 585
R64 B.n81 B.n80 585
R65 B.n79 B.n78 585
R66 B.n77 B.n76 585
R67 B.n75 B.n74 585
R68 B.n73 B.n72 585
R69 B.n71 B.n70 585
R70 B.n69 B.n68 585
R71 B.n67 B.n66 585
R72 B.n39 B.n38 585
R73 B.n369 B.n40 585
R74 B.n373 B.n40 585
R75 B.n368 B.n367 585
R76 B.n367 B.n36 585
R77 B.n366 B.n35 585
R78 B.n379 B.n35 585
R79 B.n365 B.n34 585
R80 B.n380 B.n34 585
R81 B.n364 B.n33 585
R82 B.n381 B.n33 585
R83 B.n363 B.n362 585
R84 B.n362 B.n32 585
R85 B.n361 B.n28 585
R86 B.n387 B.n28 585
R87 B.n360 B.n27 585
R88 B.n388 B.n27 585
R89 B.n359 B.n26 585
R90 B.n389 B.n26 585
R91 B.n358 B.n357 585
R92 B.n357 B.n22 585
R93 B.n356 B.n21 585
R94 B.n395 B.n21 585
R95 B.n355 B.n20 585
R96 B.n396 B.n20 585
R97 B.n354 B.n19 585
R98 B.n397 B.n19 585
R99 B.n353 B.n352 585
R100 B.n352 B.n15 585
R101 B.n351 B.n14 585
R102 B.n403 B.n14 585
R103 B.n350 B.n13 585
R104 B.n404 B.n13 585
R105 B.n349 B.n12 585
R106 B.n405 B.n12 585
R107 B.n348 B.n347 585
R108 B.n347 B.n346 585
R109 B.n345 B.n344 585
R110 B.n345 B.n8 585
R111 B.n343 B.n7 585
R112 B.n412 B.n7 585
R113 B.n342 B.n6 585
R114 B.n413 B.n6 585
R115 B.n341 B.n5 585
R116 B.n414 B.n5 585
R117 B.n340 B.n339 585
R118 B.n339 B.n4 585
R119 B.n338 B.n140 585
R120 B.n338 B.n337 585
R121 B.n328 B.n141 585
R122 B.n142 B.n141 585
R123 B.n330 B.n329 585
R124 B.n331 B.n330 585
R125 B.n327 B.n147 585
R126 B.n147 B.n146 585
R127 B.n326 B.n325 585
R128 B.n325 B.n324 585
R129 B.n149 B.n148 585
R130 B.n150 B.n149 585
R131 B.n317 B.n316 585
R132 B.n318 B.n317 585
R133 B.n315 B.n155 585
R134 B.n155 B.n154 585
R135 B.n314 B.n313 585
R136 B.n313 B.n312 585
R137 B.n157 B.n156 585
R138 B.n158 B.n157 585
R139 B.n305 B.n304 585
R140 B.n306 B.n305 585
R141 B.n303 B.n163 585
R142 B.n163 B.n162 585
R143 B.n302 B.n301 585
R144 B.n301 B.n300 585
R145 B.n165 B.n164 585
R146 B.n293 B.n165 585
R147 B.n292 B.n291 585
R148 B.n294 B.n292 585
R149 B.n290 B.n170 585
R150 B.n170 B.n169 585
R151 B.n289 B.n288 585
R152 B.n288 B.n287 585
R153 B.n172 B.n171 585
R154 B.n173 B.n172 585
R155 B.n280 B.n279 585
R156 B.n281 B.n280 585
R157 B.n176 B.n175 585
R158 B.n201 B.n200 585
R159 B.n202 B.n198 585
R160 B.n198 B.n177 585
R161 B.n204 B.n203 585
R162 B.n206 B.n197 585
R163 B.n209 B.n208 585
R164 B.n210 B.n196 585
R165 B.n212 B.n211 585
R166 B.n214 B.n195 585
R167 B.n217 B.n216 585
R168 B.n218 B.n194 585
R169 B.n220 B.n219 585
R170 B.n222 B.n193 585
R171 B.n225 B.n224 585
R172 B.n226 B.n190 585
R173 B.n229 B.n228 585
R174 B.n231 B.n189 585
R175 B.n234 B.n233 585
R176 B.n235 B.n188 585
R177 B.n237 B.n236 585
R178 B.n239 B.n187 585
R179 B.n242 B.n241 585
R180 B.n243 B.n186 585
R181 B.n248 B.n247 585
R182 B.n250 B.n185 585
R183 B.n253 B.n252 585
R184 B.n254 B.n184 585
R185 B.n256 B.n255 585
R186 B.n258 B.n183 585
R187 B.n261 B.n260 585
R188 B.n262 B.n182 585
R189 B.n264 B.n263 585
R190 B.n266 B.n181 585
R191 B.n269 B.n268 585
R192 B.n270 B.n180 585
R193 B.n272 B.n271 585
R194 B.n274 B.n179 585
R195 B.n277 B.n276 585
R196 B.n278 B.n178 585
R197 B.n283 B.n282 585
R198 B.n282 B.n281 585
R199 B.n284 B.n174 585
R200 B.n174 B.n173 585
R201 B.n286 B.n285 585
R202 B.n287 B.n286 585
R203 B.n168 B.n167 585
R204 B.n169 B.n168 585
R205 B.n296 B.n295 585
R206 B.n295 B.n294 585
R207 B.n297 B.n166 585
R208 B.n293 B.n166 585
R209 B.n299 B.n298 585
R210 B.n300 B.n299 585
R211 B.n161 B.n160 585
R212 B.n162 B.n161 585
R213 B.n308 B.n307 585
R214 B.n307 B.n306 585
R215 B.n309 B.n159 585
R216 B.n159 B.n158 585
R217 B.n311 B.n310 585
R218 B.n312 B.n311 585
R219 B.n153 B.n152 585
R220 B.n154 B.n153 585
R221 B.n320 B.n319 585
R222 B.n319 B.n318 585
R223 B.n321 B.n151 585
R224 B.n151 B.n150 585
R225 B.n323 B.n322 585
R226 B.n324 B.n323 585
R227 B.n145 B.n144 585
R228 B.n146 B.n145 585
R229 B.n333 B.n332 585
R230 B.n332 B.n331 585
R231 B.n334 B.n143 585
R232 B.n143 B.n142 585
R233 B.n336 B.n335 585
R234 B.n337 B.n336 585
R235 B.n3 B.n0 585
R236 B.n4 B.n3 585
R237 B.n411 B.n1 585
R238 B.n412 B.n411 585
R239 B.n410 B.n409 585
R240 B.n410 B.n8 585
R241 B.n408 B.n9 585
R242 B.n346 B.n9 585
R243 B.n407 B.n406 585
R244 B.n406 B.n405 585
R245 B.n11 B.n10 585
R246 B.n404 B.n11 585
R247 B.n402 B.n401 585
R248 B.n403 B.n402 585
R249 B.n400 B.n16 585
R250 B.n16 B.n15 585
R251 B.n399 B.n398 585
R252 B.n398 B.n397 585
R253 B.n18 B.n17 585
R254 B.n396 B.n18 585
R255 B.n394 B.n393 585
R256 B.n395 B.n394 585
R257 B.n392 B.n23 585
R258 B.n23 B.n22 585
R259 B.n391 B.n390 585
R260 B.n390 B.n389 585
R261 B.n25 B.n24 585
R262 B.n388 B.n25 585
R263 B.n386 B.n385 585
R264 B.n387 B.n386 585
R265 B.n384 B.n29 585
R266 B.n32 B.n29 585
R267 B.n383 B.n382 585
R268 B.n382 B.n381 585
R269 B.n31 B.n30 585
R270 B.n380 B.n31 585
R271 B.n378 B.n377 585
R272 B.n379 B.n378 585
R273 B.n376 B.n37 585
R274 B.n37 B.n36 585
R275 B.n375 B.n374 585
R276 B.n374 B.n373 585
R277 B.n415 B.n414 585
R278 B.n413 B.n2 585
R279 B.n374 B.n39 540.549
R280 B.n371 B.n40 540.549
R281 B.n280 B.n178 540.549
R282 B.n282 B.n176 540.549
R283 B.n64 B.t15 266.221
R284 B.n61 B.t8 266.221
R285 B.n244 B.t12 266.221
R286 B.n191 B.t4 266.221
R287 B.n372 B.n59 256.663
R288 B.n372 B.n58 256.663
R289 B.n372 B.n57 256.663
R290 B.n372 B.n56 256.663
R291 B.n372 B.n55 256.663
R292 B.n372 B.n54 256.663
R293 B.n372 B.n53 256.663
R294 B.n372 B.n52 256.663
R295 B.n372 B.n51 256.663
R296 B.n372 B.n50 256.663
R297 B.n372 B.n49 256.663
R298 B.n372 B.n48 256.663
R299 B.n372 B.n47 256.663
R300 B.n372 B.n46 256.663
R301 B.n372 B.n45 256.663
R302 B.n372 B.n44 256.663
R303 B.n372 B.n43 256.663
R304 B.n372 B.n42 256.663
R305 B.n372 B.n41 256.663
R306 B.n199 B.n177 256.663
R307 B.n205 B.n177 256.663
R308 B.n207 B.n177 256.663
R309 B.n213 B.n177 256.663
R310 B.n215 B.n177 256.663
R311 B.n221 B.n177 256.663
R312 B.n223 B.n177 256.663
R313 B.n230 B.n177 256.663
R314 B.n232 B.n177 256.663
R315 B.n238 B.n177 256.663
R316 B.n240 B.n177 256.663
R317 B.n249 B.n177 256.663
R318 B.n251 B.n177 256.663
R319 B.n257 B.n177 256.663
R320 B.n259 B.n177 256.663
R321 B.n265 B.n177 256.663
R322 B.n267 B.n177 256.663
R323 B.n273 B.n177 256.663
R324 B.n275 B.n177 256.663
R325 B.n417 B.n416 256.663
R326 B.n281 B.n177 187.953
R327 B.n373 B.n372 187.953
R328 B.n68 B.n67 163.367
R329 B.n72 B.n71 163.367
R330 B.n76 B.n75 163.367
R331 B.n80 B.n79 163.367
R332 B.n84 B.n83 163.367
R333 B.n88 B.n87 163.367
R334 B.n92 B.n91 163.367
R335 B.n97 B.n96 163.367
R336 B.n101 B.n100 163.367
R337 B.n105 B.n104 163.367
R338 B.n109 B.n108 163.367
R339 B.n113 B.n112 163.367
R340 B.n117 B.n116 163.367
R341 B.n121 B.n120 163.367
R342 B.n125 B.n124 163.367
R343 B.n129 B.n128 163.367
R344 B.n133 B.n132 163.367
R345 B.n137 B.n136 163.367
R346 B.n371 B.n60 163.367
R347 B.n280 B.n172 163.367
R348 B.n288 B.n172 163.367
R349 B.n288 B.n170 163.367
R350 B.n292 B.n170 163.367
R351 B.n292 B.n165 163.367
R352 B.n301 B.n165 163.367
R353 B.n301 B.n163 163.367
R354 B.n305 B.n163 163.367
R355 B.n305 B.n157 163.367
R356 B.n313 B.n157 163.367
R357 B.n313 B.n155 163.367
R358 B.n317 B.n155 163.367
R359 B.n317 B.n149 163.367
R360 B.n325 B.n149 163.367
R361 B.n325 B.n147 163.367
R362 B.n330 B.n147 163.367
R363 B.n330 B.n141 163.367
R364 B.n338 B.n141 163.367
R365 B.n339 B.n338 163.367
R366 B.n339 B.n5 163.367
R367 B.n6 B.n5 163.367
R368 B.n7 B.n6 163.367
R369 B.n345 B.n7 163.367
R370 B.n347 B.n345 163.367
R371 B.n347 B.n12 163.367
R372 B.n13 B.n12 163.367
R373 B.n14 B.n13 163.367
R374 B.n352 B.n14 163.367
R375 B.n352 B.n19 163.367
R376 B.n20 B.n19 163.367
R377 B.n21 B.n20 163.367
R378 B.n357 B.n21 163.367
R379 B.n357 B.n26 163.367
R380 B.n27 B.n26 163.367
R381 B.n28 B.n27 163.367
R382 B.n362 B.n28 163.367
R383 B.n362 B.n33 163.367
R384 B.n34 B.n33 163.367
R385 B.n35 B.n34 163.367
R386 B.n367 B.n35 163.367
R387 B.n367 B.n40 163.367
R388 B.n200 B.n198 163.367
R389 B.n204 B.n198 163.367
R390 B.n208 B.n206 163.367
R391 B.n212 B.n196 163.367
R392 B.n216 B.n214 163.367
R393 B.n220 B.n194 163.367
R394 B.n224 B.n222 163.367
R395 B.n229 B.n190 163.367
R396 B.n233 B.n231 163.367
R397 B.n237 B.n188 163.367
R398 B.n241 B.n239 163.367
R399 B.n248 B.n186 163.367
R400 B.n252 B.n250 163.367
R401 B.n256 B.n184 163.367
R402 B.n260 B.n258 163.367
R403 B.n264 B.n182 163.367
R404 B.n268 B.n266 163.367
R405 B.n272 B.n180 163.367
R406 B.n276 B.n274 163.367
R407 B.n282 B.n174 163.367
R408 B.n286 B.n174 163.367
R409 B.n286 B.n168 163.367
R410 B.n295 B.n168 163.367
R411 B.n295 B.n166 163.367
R412 B.n299 B.n166 163.367
R413 B.n299 B.n161 163.367
R414 B.n307 B.n161 163.367
R415 B.n307 B.n159 163.367
R416 B.n311 B.n159 163.367
R417 B.n311 B.n153 163.367
R418 B.n319 B.n153 163.367
R419 B.n319 B.n151 163.367
R420 B.n323 B.n151 163.367
R421 B.n323 B.n145 163.367
R422 B.n332 B.n145 163.367
R423 B.n332 B.n143 163.367
R424 B.n336 B.n143 163.367
R425 B.n336 B.n3 163.367
R426 B.n415 B.n3 163.367
R427 B.n411 B.n2 163.367
R428 B.n411 B.n410 163.367
R429 B.n410 B.n9 163.367
R430 B.n406 B.n9 163.367
R431 B.n406 B.n11 163.367
R432 B.n402 B.n11 163.367
R433 B.n402 B.n16 163.367
R434 B.n398 B.n16 163.367
R435 B.n398 B.n18 163.367
R436 B.n394 B.n18 163.367
R437 B.n394 B.n23 163.367
R438 B.n390 B.n23 163.367
R439 B.n390 B.n25 163.367
R440 B.n386 B.n25 163.367
R441 B.n386 B.n29 163.367
R442 B.n382 B.n29 163.367
R443 B.n382 B.n31 163.367
R444 B.n378 B.n31 163.367
R445 B.n378 B.n37 163.367
R446 B.n374 B.n37 163.367
R447 B.n61 B.t10 105.957
R448 B.n244 B.t14 105.957
R449 B.n64 B.t16 105.954
R450 B.n191 B.t7 105.954
R451 B.n281 B.n173 91.9489
R452 B.n287 B.n173 91.9489
R453 B.n287 B.n169 91.9489
R454 B.n294 B.n169 91.9489
R455 B.n294 B.n293 91.9489
R456 B.n300 B.n162 91.9489
R457 B.n306 B.n162 91.9489
R458 B.n306 B.n158 91.9489
R459 B.n312 B.n158 91.9489
R460 B.n312 B.n154 91.9489
R461 B.n318 B.n154 91.9489
R462 B.n324 B.n150 91.9489
R463 B.n324 B.n146 91.9489
R464 B.n331 B.n146 91.9489
R465 B.n337 B.n142 91.9489
R466 B.n337 B.n4 91.9489
R467 B.n414 B.n4 91.9489
R468 B.n414 B.n413 91.9489
R469 B.n413 B.n412 91.9489
R470 B.n412 B.n8 91.9489
R471 B.n346 B.n8 91.9489
R472 B.n405 B.n404 91.9489
R473 B.n404 B.n403 91.9489
R474 B.n403 B.n15 91.9489
R475 B.n397 B.n396 91.9489
R476 B.n396 B.n395 91.9489
R477 B.n395 B.n22 91.9489
R478 B.n389 B.n22 91.9489
R479 B.n389 B.n388 91.9489
R480 B.n388 B.n387 91.9489
R481 B.n381 B.n32 91.9489
R482 B.n381 B.n380 91.9489
R483 B.n380 B.n379 91.9489
R484 B.n379 B.n36 91.9489
R485 B.n373 B.n36 91.9489
R486 B.n62 B.t11 78.2227
R487 B.n245 B.t13 78.2227
R488 B.n65 B.t17 78.2209
R489 B.n192 B.t6 78.2209
R490 B.n300 B.t5 75.7227
R491 B.n387 B.t9 75.7227
R492 B.n331 B.t1 73.0183
R493 B.n405 B.t3 73.0183
R494 B.n41 B.n39 71.676
R495 B.n68 B.n42 71.676
R496 B.n72 B.n43 71.676
R497 B.n76 B.n44 71.676
R498 B.n80 B.n45 71.676
R499 B.n84 B.n46 71.676
R500 B.n88 B.n47 71.676
R501 B.n92 B.n48 71.676
R502 B.n97 B.n49 71.676
R503 B.n101 B.n50 71.676
R504 B.n105 B.n51 71.676
R505 B.n109 B.n52 71.676
R506 B.n113 B.n53 71.676
R507 B.n117 B.n54 71.676
R508 B.n121 B.n55 71.676
R509 B.n125 B.n56 71.676
R510 B.n129 B.n57 71.676
R511 B.n133 B.n58 71.676
R512 B.n137 B.n59 71.676
R513 B.n60 B.n59 71.676
R514 B.n136 B.n58 71.676
R515 B.n132 B.n57 71.676
R516 B.n128 B.n56 71.676
R517 B.n124 B.n55 71.676
R518 B.n120 B.n54 71.676
R519 B.n116 B.n53 71.676
R520 B.n112 B.n52 71.676
R521 B.n108 B.n51 71.676
R522 B.n104 B.n50 71.676
R523 B.n100 B.n49 71.676
R524 B.n96 B.n48 71.676
R525 B.n91 B.n47 71.676
R526 B.n87 B.n46 71.676
R527 B.n83 B.n45 71.676
R528 B.n79 B.n44 71.676
R529 B.n75 B.n43 71.676
R530 B.n71 B.n42 71.676
R531 B.n67 B.n41 71.676
R532 B.n199 B.n176 71.676
R533 B.n205 B.n204 71.676
R534 B.n208 B.n207 71.676
R535 B.n213 B.n212 71.676
R536 B.n216 B.n215 71.676
R537 B.n221 B.n220 71.676
R538 B.n224 B.n223 71.676
R539 B.n230 B.n229 71.676
R540 B.n233 B.n232 71.676
R541 B.n238 B.n237 71.676
R542 B.n241 B.n240 71.676
R543 B.n249 B.n248 71.676
R544 B.n252 B.n251 71.676
R545 B.n257 B.n256 71.676
R546 B.n260 B.n259 71.676
R547 B.n265 B.n264 71.676
R548 B.n268 B.n267 71.676
R549 B.n273 B.n272 71.676
R550 B.n276 B.n275 71.676
R551 B.n200 B.n199 71.676
R552 B.n206 B.n205 71.676
R553 B.n207 B.n196 71.676
R554 B.n214 B.n213 71.676
R555 B.n215 B.n194 71.676
R556 B.n222 B.n221 71.676
R557 B.n223 B.n190 71.676
R558 B.n231 B.n230 71.676
R559 B.n232 B.n188 71.676
R560 B.n239 B.n238 71.676
R561 B.n240 B.n186 71.676
R562 B.n250 B.n249 71.676
R563 B.n251 B.n184 71.676
R564 B.n258 B.n257 71.676
R565 B.n259 B.n182 71.676
R566 B.n266 B.n265 71.676
R567 B.n267 B.n180 71.676
R568 B.n274 B.n273 71.676
R569 B.n275 B.n178 71.676
R570 B.n416 B.n415 71.676
R571 B.n416 B.n2 71.676
R572 B.n94 B.n65 59.5399
R573 B.n63 B.n62 59.5399
R574 B.n246 B.n245 59.5399
R575 B.n227 B.n192 59.5399
R576 B.n318 B.t2 54.0878
R577 B.n397 B.t0 54.0878
R578 B.t2 B.n150 37.8616
R579 B.t0 B.n15 37.8616
R580 B.n283 B.n175 35.1225
R581 B.n279 B.n278 35.1225
R582 B.n370 B.n369 35.1225
R583 B.n375 B.n38 35.1225
R584 B.n65 B.n64 27.7338
R585 B.n62 B.n61 27.7338
R586 B.n245 B.n244 27.7338
R587 B.n192 B.n191 27.7338
R588 B.t1 B.n142 18.931
R589 B.n346 B.t3 18.931
R590 B B.n417 18.0485
R591 B.n293 B.t5 16.2267
R592 B.n32 B.t9 16.2267
R593 B.n284 B.n283 10.6151
R594 B.n285 B.n284 10.6151
R595 B.n285 B.n167 10.6151
R596 B.n296 B.n167 10.6151
R597 B.n297 B.n296 10.6151
R598 B.n298 B.n297 10.6151
R599 B.n298 B.n160 10.6151
R600 B.n308 B.n160 10.6151
R601 B.n309 B.n308 10.6151
R602 B.n310 B.n309 10.6151
R603 B.n310 B.n152 10.6151
R604 B.n320 B.n152 10.6151
R605 B.n321 B.n320 10.6151
R606 B.n322 B.n321 10.6151
R607 B.n322 B.n144 10.6151
R608 B.n333 B.n144 10.6151
R609 B.n334 B.n333 10.6151
R610 B.n335 B.n334 10.6151
R611 B.n335 B.n0 10.6151
R612 B.n201 B.n175 10.6151
R613 B.n202 B.n201 10.6151
R614 B.n203 B.n202 10.6151
R615 B.n203 B.n197 10.6151
R616 B.n209 B.n197 10.6151
R617 B.n210 B.n209 10.6151
R618 B.n211 B.n210 10.6151
R619 B.n211 B.n195 10.6151
R620 B.n217 B.n195 10.6151
R621 B.n218 B.n217 10.6151
R622 B.n219 B.n218 10.6151
R623 B.n219 B.n193 10.6151
R624 B.n225 B.n193 10.6151
R625 B.n226 B.n225 10.6151
R626 B.n228 B.n189 10.6151
R627 B.n234 B.n189 10.6151
R628 B.n235 B.n234 10.6151
R629 B.n236 B.n235 10.6151
R630 B.n236 B.n187 10.6151
R631 B.n242 B.n187 10.6151
R632 B.n243 B.n242 10.6151
R633 B.n247 B.n243 10.6151
R634 B.n253 B.n185 10.6151
R635 B.n254 B.n253 10.6151
R636 B.n255 B.n254 10.6151
R637 B.n255 B.n183 10.6151
R638 B.n261 B.n183 10.6151
R639 B.n262 B.n261 10.6151
R640 B.n263 B.n262 10.6151
R641 B.n263 B.n181 10.6151
R642 B.n269 B.n181 10.6151
R643 B.n270 B.n269 10.6151
R644 B.n271 B.n270 10.6151
R645 B.n271 B.n179 10.6151
R646 B.n277 B.n179 10.6151
R647 B.n278 B.n277 10.6151
R648 B.n279 B.n171 10.6151
R649 B.n289 B.n171 10.6151
R650 B.n290 B.n289 10.6151
R651 B.n291 B.n290 10.6151
R652 B.n291 B.n164 10.6151
R653 B.n302 B.n164 10.6151
R654 B.n303 B.n302 10.6151
R655 B.n304 B.n303 10.6151
R656 B.n304 B.n156 10.6151
R657 B.n314 B.n156 10.6151
R658 B.n315 B.n314 10.6151
R659 B.n316 B.n315 10.6151
R660 B.n316 B.n148 10.6151
R661 B.n326 B.n148 10.6151
R662 B.n327 B.n326 10.6151
R663 B.n329 B.n327 10.6151
R664 B.n329 B.n328 10.6151
R665 B.n328 B.n140 10.6151
R666 B.n340 B.n140 10.6151
R667 B.n341 B.n340 10.6151
R668 B.n342 B.n341 10.6151
R669 B.n343 B.n342 10.6151
R670 B.n344 B.n343 10.6151
R671 B.n348 B.n344 10.6151
R672 B.n349 B.n348 10.6151
R673 B.n350 B.n349 10.6151
R674 B.n351 B.n350 10.6151
R675 B.n353 B.n351 10.6151
R676 B.n354 B.n353 10.6151
R677 B.n355 B.n354 10.6151
R678 B.n356 B.n355 10.6151
R679 B.n358 B.n356 10.6151
R680 B.n359 B.n358 10.6151
R681 B.n360 B.n359 10.6151
R682 B.n361 B.n360 10.6151
R683 B.n363 B.n361 10.6151
R684 B.n364 B.n363 10.6151
R685 B.n365 B.n364 10.6151
R686 B.n366 B.n365 10.6151
R687 B.n368 B.n366 10.6151
R688 B.n369 B.n368 10.6151
R689 B.n409 B.n1 10.6151
R690 B.n409 B.n408 10.6151
R691 B.n408 B.n407 10.6151
R692 B.n407 B.n10 10.6151
R693 B.n401 B.n10 10.6151
R694 B.n401 B.n400 10.6151
R695 B.n400 B.n399 10.6151
R696 B.n399 B.n17 10.6151
R697 B.n393 B.n17 10.6151
R698 B.n393 B.n392 10.6151
R699 B.n392 B.n391 10.6151
R700 B.n391 B.n24 10.6151
R701 B.n385 B.n24 10.6151
R702 B.n385 B.n384 10.6151
R703 B.n384 B.n383 10.6151
R704 B.n383 B.n30 10.6151
R705 B.n377 B.n30 10.6151
R706 B.n377 B.n376 10.6151
R707 B.n376 B.n375 10.6151
R708 B.n66 B.n38 10.6151
R709 B.n69 B.n66 10.6151
R710 B.n70 B.n69 10.6151
R711 B.n73 B.n70 10.6151
R712 B.n74 B.n73 10.6151
R713 B.n77 B.n74 10.6151
R714 B.n78 B.n77 10.6151
R715 B.n81 B.n78 10.6151
R716 B.n82 B.n81 10.6151
R717 B.n85 B.n82 10.6151
R718 B.n86 B.n85 10.6151
R719 B.n89 B.n86 10.6151
R720 B.n90 B.n89 10.6151
R721 B.n93 B.n90 10.6151
R722 B.n98 B.n95 10.6151
R723 B.n99 B.n98 10.6151
R724 B.n102 B.n99 10.6151
R725 B.n103 B.n102 10.6151
R726 B.n106 B.n103 10.6151
R727 B.n107 B.n106 10.6151
R728 B.n110 B.n107 10.6151
R729 B.n111 B.n110 10.6151
R730 B.n115 B.n114 10.6151
R731 B.n118 B.n115 10.6151
R732 B.n119 B.n118 10.6151
R733 B.n122 B.n119 10.6151
R734 B.n123 B.n122 10.6151
R735 B.n126 B.n123 10.6151
R736 B.n127 B.n126 10.6151
R737 B.n130 B.n127 10.6151
R738 B.n131 B.n130 10.6151
R739 B.n134 B.n131 10.6151
R740 B.n135 B.n134 10.6151
R741 B.n138 B.n135 10.6151
R742 B.n139 B.n138 10.6151
R743 B.n370 B.n139 10.6151
R744 B.n417 B.n0 8.11757
R745 B.n417 B.n1 8.11757
R746 B.n228 B.n227 6.5566
R747 B.n247 B.n246 6.5566
R748 B.n95 B.n94 6.5566
R749 B.n111 B.n63 6.5566
R750 B.n227 B.n226 4.05904
R751 B.n246 B.n185 4.05904
R752 B.n94 B.n93 4.05904
R753 B.n114 B.n63 4.05904
R754 VN.n0 VN.t3 116.98
R755 VN.n1 VN.t2 116.98
R756 VN.n1 VN.t0 116.892
R757 VN.n0 VN.t1 116.892
R758 VN VN.n1 66.4023
R759 VN VN.n0 31.2622
R760 VDD2.n2 VDD2.n0 112.647
R761 VDD2.n2 VDD2.n1 82.7679
R762 VDD2.n1 VDD2.t3 6.92358
R763 VDD2.n1 VDD2.t1 6.92358
R764 VDD2.n0 VDD2.t0 6.92358
R765 VDD2.n0 VDD2.t2 6.92358
R766 VDD2 VDD2.n2 0.0586897
C0 VDD1 VP 1.27889f
C1 VP VTAIL 1.29371f
C2 VP VN 3.41865f
C3 VP VDD2 0.304835f
C4 VDD1 VTAIL 2.69272f
C5 VDD1 VN 0.153096f
C6 VN VTAIL 1.2796f
C7 VDD1 VDD2 0.662501f
C8 VDD2 VTAIL 2.73687f
C9 VN VDD2 1.12807f
C10 VDD2 B 2.171837f
C11 VDD1 B 4.01883f
C12 VTAIL B 3.612058f
C13 VN B 6.41926f
C14 VP B 4.986817f
C15 VDD2.t0 B 0.042808f
C16 VDD2.t2 B 0.042808f
C17 VDD2.n0 B 0.49598f
C18 VDD2.t3 B 0.042808f
C19 VDD2.t1 B 0.042808f
C20 VDD2.n1 B 0.314037f
C21 VDD2.n2 B 1.63943f
C22 VN.t3 B 0.274652f
C23 VN.t1 B 0.274513f
C24 VN.n0 B 0.248208f
C25 VN.t2 B 0.274652f
C26 VN.t0 B 0.274513f
C27 VN.n1 B 0.718677f
C28 VDD1.t1 B 0.041727f
C29 VDD1.t3 B 0.041727f
C30 VDD1.n0 B 0.306261f
C31 VDD1.t2 B 0.041727f
C32 VDD1.t0 B 0.041727f
C33 VDD1.n1 B 0.495935f
C34 VTAIL.t3 B 0.278811f
C35 VTAIL.n0 B 0.195263f
C36 VTAIL.t7 B 0.278811f
C37 VTAIL.n1 B 0.221466f
C38 VTAIL.t6 B 0.278811f
C39 VTAIL.n2 B 0.570911f
C40 VTAIL.t2 B 0.278812f
C41 VTAIL.n3 B 0.57091f
C42 VTAIL.t1 B 0.278812f
C43 VTAIL.n4 B 0.221465f
C44 VTAIL.t5 B 0.278812f
C45 VTAIL.n5 B 0.221465f
C46 VTAIL.t4 B 0.278811f
C47 VTAIL.n6 B 0.570911f
C48 VTAIL.t0 B 0.278811f
C49 VTAIL.n7 B 0.539245f
C50 VP.t0 B 0.27756f
C51 VP.t2 B 0.277699f
C52 VP.n0 B 0.716585f
C53 VP.n1 B 1.26023f
C54 VP.t1 B 0.253993f
C55 VP.n2 B 0.148746f
C56 VP.t3 B 0.253993f
C57 VP.n3 B 0.148746f
C58 VP.n4 B 0.034109f
.ends

