* NGSPICE file created from diff_pair_sample_1211.ext - technology: sky130A

.subckt diff_pair_sample_1211 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n2818_n2870# sky130_fd_pr__pfet_01v8 ad=3.7089 pd=19.8 as=0 ps=0 w=9.51 l=2.75
X1 B.t8 B.t6 B.t7 w_n2818_n2870# sky130_fd_pr__pfet_01v8 ad=3.7089 pd=19.8 as=0 ps=0 w=9.51 l=2.75
X2 B.t5 B.t3 B.t4 w_n2818_n2870# sky130_fd_pr__pfet_01v8 ad=3.7089 pd=19.8 as=0 ps=0 w=9.51 l=2.75
X3 B.t2 B.t0 B.t1 w_n2818_n2870# sky130_fd_pr__pfet_01v8 ad=3.7089 pd=19.8 as=0 ps=0 w=9.51 l=2.75
X4 VDD2.t3 VN.t0 VTAIL.t5 w_n2818_n2870# sky130_fd_pr__pfet_01v8 ad=1.56915 pd=9.84 as=3.7089 ps=19.8 w=9.51 l=2.75
X5 VTAIL.t0 VP.t0 VDD1.t3 w_n2818_n2870# sky130_fd_pr__pfet_01v8 ad=3.7089 pd=19.8 as=1.56915 ps=9.84 w=9.51 l=2.75
X6 VDD2.t2 VN.t1 VTAIL.t7 w_n2818_n2870# sky130_fd_pr__pfet_01v8 ad=1.56915 pd=9.84 as=3.7089 ps=19.8 w=9.51 l=2.75
X7 VTAIL.t6 VN.t2 VDD2.t1 w_n2818_n2870# sky130_fd_pr__pfet_01v8 ad=3.7089 pd=19.8 as=1.56915 ps=9.84 w=9.51 l=2.75
X8 VTAIL.t4 VN.t3 VDD2.t0 w_n2818_n2870# sky130_fd_pr__pfet_01v8 ad=3.7089 pd=19.8 as=1.56915 ps=9.84 w=9.51 l=2.75
X9 VTAIL.t2 VP.t1 VDD1.t2 w_n2818_n2870# sky130_fd_pr__pfet_01v8 ad=3.7089 pd=19.8 as=1.56915 ps=9.84 w=9.51 l=2.75
X10 VDD1.t1 VP.t2 VTAIL.t1 w_n2818_n2870# sky130_fd_pr__pfet_01v8 ad=1.56915 pd=9.84 as=3.7089 ps=19.8 w=9.51 l=2.75
X11 VDD1.t0 VP.t3 VTAIL.t3 w_n2818_n2870# sky130_fd_pr__pfet_01v8 ad=1.56915 pd=9.84 as=3.7089 ps=19.8 w=9.51 l=2.75
R0 B.n329 B.n328 585
R1 B.n327 B.n100 585
R2 B.n326 B.n325 585
R3 B.n324 B.n101 585
R4 B.n323 B.n322 585
R5 B.n321 B.n102 585
R6 B.n320 B.n319 585
R7 B.n318 B.n103 585
R8 B.n317 B.n316 585
R9 B.n315 B.n104 585
R10 B.n314 B.n313 585
R11 B.n312 B.n105 585
R12 B.n311 B.n310 585
R13 B.n309 B.n106 585
R14 B.n308 B.n307 585
R15 B.n306 B.n107 585
R16 B.n305 B.n304 585
R17 B.n303 B.n108 585
R18 B.n302 B.n301 585
R19 B.n300 B.n109 585
R20 B.n299 B.n298 585
R21 B.n297 B.n110 585
R22 B.n296 B.n295 585
R23 B.n294 B.n111 585
R24 B.n293 B.n292 585
R25 B.n291 B.n112 585
R26 B.n290 B.n289 585
R27 B.n288 B.n113 585
R28 B.n287 B.n286 585
R29 B.n285 B.n114 585
R30 B.n284 B.n283 585
R31 B.n282 B.n115 585
R32 B.n281 B.n280 585
R33 B.n279 B.n116 585
R34 B.n277 B.n276 585
R35 B.n275 B.n119 585
R36 B.n274 B.n273 585
R37 B.n272 B.n120 585
R38 B.n271 B.n270 585
R39 B.n269 B.n121 585
R40 B.n268 B.n267 585
R41 B.n266 B.n122 585
R42 B.n265 B.n264 585
R43 B.n263 B.n123 585
R44 B.n262 B.n261 585
R45 B.n257 B.n124 585
R46 B.n256 B.n255 585
R47 B.n254 B.n125 585
R48 B.n253 B.n252 585
R49 B.n251 B.n126 585
R50 B.n250 B.n249 585
R51 B.n248 B.n127 585
R52 B.n247 B.n246 585
R53 B.n245 B.n128 585
R54 B.n244 B.n243 585
R55 B.n242 B.n129 585
R56 B.n241 B.n240 585
R57 B.n239 B.n130 585
R58 B.n238 B.n237 585
R59 B.n236 B.n131 585
R60 B.n235 B.n234 585
R61 B.n233 B.n132 585
R62 B.n232 B.n231 585
R63 B.n230 B.n133 585
R64 B.n229 B.n228 585
R65 B.n227 B.n134 585
R66 B.n226 B.n225 585
R67 B.n224 B.n135 585
R68 B.n223 B.n222 585
R69 B.n221 B.n136 585
R70 B.n220 B.n219 585
R71 B.n218 B.n137 585
R72 B.n217 B.n216 585
R73 B.n215 B.n138 585
R74 B.n214 B.n213 585
R75 B.n212 B.n139 585
R76 B.n211 B.n210 585
R77 B.n209 B.n140 585
R78 B.n330 B.n99 585
R79 B.n332 B.n331 585
R80 B.n333 B.n98 585
R81 B.n335 B.n334 585
R82 B.n336 B.n97 585
R83 B.n338 B.n337 585
R84 B.n339 B.n96 585
R85 B.n341 B.n340 585
R86 B.n342 B.n95 585
R87 B.n344 B.n343 585
R88 B.n345 B.n94 585
R89 B.n347 B.n346 585
R90 B.n348 B.n93 585
R91 B.n350 B.n349 585
R92 B.n351 B.n92 585
R93 B.n353 B.n352 585
R94 B.n354 B.n91 585
R95 B.n356 B.n355 585
R96 B.n357 B.n90 585
R97 B.n359 B.n358 585
R98 B.n360 B.n89 585
R99 B.n362 B.n361 585
R100 B.n363 B.n88 585
R101 B.n365 B.n364 585
R102 B.n366 B.n87 585
R103 B.n368 B.n367 585
R104 B.n369 B.n86 585
R105 B.n371 B.n370 585
R106 B.n372 B.n85 585
R107 B.n374 B.n373 585
R108 B.n375 B.n84 585
R109 B.n377 B.n376 585
R110 B.n378 B.n83 585
R111 B.n380 B.n379 585
R112 B.n381 B.n82 585
R113 B.n383 B.n382 585
R114 B.n384 B.n81 585
R115 B.n386 B.n385 585
R116 B.n387 B.n80 585
R117 B.n389 B.n388 585
R118 B.n390 B.n79 585
R119 B.n392 B.n391 585
R120 B.n393 B.n78 585
R121 B.n395 B.n394 585
R122 B.n396 B.n77 585
R123 B.n398 B.n397 585
R124 B.n399 B.n76 585
R125 B.n401 B.n400 585
R126 B.n402 B.n75 585
R127 B.n404 B.n403 585
R128 B.n405 B.n74 585
R129 B.n407 B.n406 585
R130 B.n408 B.n73 585
R131 B.n410 B.n409 585
R132 B.n411 B.n72 585
R133 B.n413 B.n412 585
R134 B.n414 B.n71 585
R135 B.n416 B.n415 585
R136 B.n417 B.n70 585
R137 B.n419 B.n418 585
R138 B.n420 B.n69 585
R139 B.n422 B.n421 585
R140 B.n423 B.n68 585
R141 B.n425 B.n424 585
R142 B.n426 B.n67 585
R143 B.n428 B.n427 585
R144 B.n429 B.n66 585
R145 B.n431 B.n430 585
R146 B.n432 B.n65 585
R147 B.n434 B.n433 585
R148 B.n435 B.n64 585
R149 B.n437 B.n436 585
R150 B.n555 B.n554 585
R151 B.n553 B.n20 585
R152 B.n552 B.n551 585
R153 B.n550 B.n21 585
R154 B.n549 B.n548 585
R155 B.n547 B.n22 585
R156 B.n546 B.n545 585
R157 B.n544 B.n23 585
R158 B.n543 B.n542 585
R159 B.n541 B.n24 585
R160 B.n540 B.n539 585
R161 B.n538 B.n25 585
R162 B.n537 B.n536 585
R163 B.n535 B.n26 585
R164 B.n534 B.n533 585
R165 B.n532 B.n27 585
R166 B.n531 B.n530 585
R167 B.n529 B.n28 585
R168 B.n528 B.n527 585
R169 B.n526 B.n29 585
R170 B.n525 B.n524 585
R171 B.n523 B.n30 585
R172 B.n522 B.n521 585
R173 B.n520 B.n31 585
R174 B.n519 B.n518 585
R175 B.n517 B.n32 585
R176 B.n516 B.n515 585
R177 B.n514 B.n33 585
R178 B.n513 B.n512 585
R179 B.n511 B.n34 585
R180 B.n510 B.n509 585
R181 B.n508 B.n35 585
R182 B.n507 B.n506 585
R183 B.n505 B.n36 585
R184 B.n504 B.n503 585
R185 B.n502 B.n37 585
R186 B.n501 B.n500 585
R187 B.n499 B.n41 585
R188 B.n498 B.n497 585
R189 B.n496 B.n42 585
R190 B.n495 B.n494 585
R191 B.n493 B.n43 585
R192 B.n492 B.n491 585
R193 B.n490 B.n44 585
R194 B.n488 B.n487 585
R195 B.n486 B.n47 585
R196 B.n485 B.n484 585
R197 B.n483 B.n48 585
R198 B.n482 B.n481 585
R199 B.n480 B.n49 585
R200 B.n479 B.n478 585
R201 B.n477 B.n50 585
R202 B.n476 B.n475 585
R203 B.n474 B.n51 585
R204 B.n473 B.n472 585
R205 B.n471 B.n52 585
R206 B.n470 B.n469 585
R207 B.n468 B.n53 585
R208 B.n467 B.n466 585
R209 B.n465 B.n54 585
R210 B.n464 B.n463 585
R211 B.n462 B.n55 585
R212 B.n461 B.n460 585
R213 B.n459 B.n56 585
R214 B.n458 B.n457 585
R215 B.n456 B.n57 585
R216 B.n455 B.n454 585
R217 B.n453 B.n58 585
R218 B.n452 B.n451 585
R219 B.n450 B.n59 585
R220 B.n449 B.n448 585
R221 B.n447 B.n60 585
R222 B.n446 B.n445 585
R223 B.n444 B.n61 585
R224 B.n443 B.n442 585
R225 B.n441 B.n62 585
R226 B.n440 B.n439 585
R227 B.n438 B.n63 585
R228 B.n556 B.n19 585
R229 B.n558 B.n557 585
R230 B.n559 B.n18 585
R231 B.n561 B.n560 585
R232 B.n562 B.n17 585
R233 B.n564 B.n563 585
R234 B.n565 B.n16 585
R235 B.n567 B.n566 585
R236 B.n568 B.n15 585
R237 B.n570 B.n569 585
R238 B.n571 B.n14 585
R239 B.n573 B.n572 585
R240 B.n574 B.n13 585
R241 B.n576 B.n575 585
R242 B.n577 B.n12 585
R243 B.n579 B.n578 585
R244 B.n580 B.n11 585
R245 B.n582 B.n581 585
R246 B.n583 B.n10 585
R247 B.n585 B.n584 585
R248 B.n586 B.n9 585
R249 B.n588 B.n587 585
R250 B.n589 B.n8 585
R251 B.n591 B.n590 585
R252 B.n592 B.n7 585
R253 B.n594 B.n593 585
R254 B.n595 B.n6 585
R255 B.n597 B.n596 585
R256 B.n598 B.n5 585
R257 B.n600 B.n599 585
R258 B.n601 B.n4 585
R259 B.n603 B.n602 585
R260 B.n604 B.n3 585
R261 B.n606 B.n605 585
R262 B.n607 B.n0 585
R263 B.n2 B.n1 585
R264 B.n158 B.n157 585
R265 B.n160 B.n159 585
R266 B.n161 B.n156 585
R267 B.n163 B.n162 585
R268 B.n164 B.n155 585
R269 B.n166 B.n165 585
R270 B.n167 B.n154 585
R271 B.n169 B.n168 585
R272 B.n170 B.n153 585
R273 B.n172 B.n171 585
R274 B.n173 B.n152 585
R275 B.n175 B.n174 585
R276 B.n176 B.n151 585
R277 B.n178 B.n177 585
R278 B.n179 B.n150 585
R279 B.n181 B.n180 585
R280 B.n182 B.n149 585
R281 B.n184 B.n183 585
R282 B.n185 B.n148 585
R283 B.n187 B.n186 585
R284 B.n188 B.n147 585
R285 B.n190 B.n189 585
R286 B.n191 B.n146 585
R287 B.n193 B.n192 585
R288 B.n194 B.n145 585
R289 B.n196 B.n195 585
R290 B.n197 B.n144 585
R291 B.n199 B.n198 585
R292 B.n200 B.n143 585
R293 B.n202 B.n201 585
R294 B.n203 B.n142 585
R295 B.n205 B.n204 585
R296 B.n206 B.n141 585
R297 B.n208 B.n207 585
R298 B.n207 B.n140 478.086
R299 B.n330 B.n329 478.086
R300 B.n438 B.n437 478.086
R301 B.n554 B.n19 478.086
R302 B.n117 B.t1 390.76
R303 B.n45 B.t5 390.76
R304 B.n258 B.t10 390.76
R305 B.n38 B.t8 390.76
R306 B.n118 B.t2 331.027
R307 B.n46 B.t4 331.027
R308 B.n259 B.t11 331.026
R309 B.n39 B.t7 331.026
R310 B.n258 B.t9 291.604
R311 B.n117 B.t0 291.604
R312 B.n45 B.t3 291.604
R313 B.n38 B.t6 291.604
R314 B.n609 B.n608 256.663
R315 B.n608 B.n607 235.042
R316 B.n608 B.n2 235.042
R317 B.n211 B.n140 163.367
R318 B.n212 B.n211 163.367
R319 B.n213 B.n212 163.367
R320 B.n213 B.n138 163.367
R321 B.n217 B.n138 163.367
R322 B.n218 B.n217 163.367
R323 B.n219 B.n218 163.367
R324 B.n219 B.n136 163.367
R325 B.n223 B.n136 163.367
R326 B.n224 B.n223 163.367
R327 B.n225 B.n224 163.367
R328 B.n225 B.n134 163.367
R329 B.n229 B.n134 163.367
R330 B.n230 B.n229 163.367
R331 B.n231 B.n230 163.367
R332 B.n231 B.n132 163.367
R333 B.n235 B.n132 163.367
R334 B.n236 B.n235 163.367
R335 B.n237 B.n236 163.367
R336 B.n237 B.n130 163.367
R337 B.n241 B.n130 163.367
R338 B.n242 B.n241 163.367
R339 B.n243 B.n242 163.367
R340 B.n243 B.n128 163.367
R341 B.n247 B.n128 163.367
R342 B.n248 B.n247 163.367
R343 B.n249 B.n248 163.367
R344 B.n249 B.n126 163.367
R345 B.n253 B.n126 163.367
R346 B.n254 B.n253 163.367
R347 B.n255 B.n254 163.367
R348 B.n255 B.n124 163.367
R349 B.n262 B.n124 163.367
R350 B.n263 B.n262 163.367
R351 B.n264 B.n263 163.367
R352 B.n264 B.n122 163.367
R353 B.n268 B.n122 163.367
R354 B.n269 B.n268 163.367
R355 B.n270 B.n269 163.367
R356 B.n270 B.n120 163.367
R357 B.n274 B.n120 163.367
R358 B.n275 B.n274 163.367
R359 B.n276 B.n275 163.367
R360 B.n276 B.n116 163.367
R361 B.n281 B.n116 163.367
R362 B.n282 B.n281 163.367
R363 B.n283 B.n282 163.367
R364 B.n283 B.n114 163.367
R365 B.n287 B.n114 163.367
R366 B.n288 B.n287 163.367
R367 B.n289 B.n288 163.367
R368 B.n289 B.n112 163.367
R369 B.n293 B.n112 163.367
R370 B.n294 B.n293 163.367
R371 B.n295 B.n294 163.367
R372 B.n295 B.n110 163.367
R373 B.n299 B.n110 163.367
R374 B.n300 B.n299 163.367
R375 B.n301 B.n300 163.367
R376 B.n301 B.n108 163.367
R377 B.n305 B.n108 163.367
R378 B.n306 B.n305 163.367
R379 B.n307 B.n306 163.367
R380 B.n307 B.n106 163.367
R381 B.n311 B.n106 163.367
R382 B.n312 B.n311 163.367
R383 B.n313 B.n312 163.367
R384 B.n313 B.n104 163.367
R385 B.n317 B.n104 163.367
R386 B.n318 B.n317 163.367
R387 B.n319 B.n318 163.367
R388 B.n319 B.n102 163.367
R389 B.n323 B.n102 163.367
R390 B.n324 B.n323 163.367
R391 B.n325 B.n324 163.367
R392 B.n325 B.n100 163.367
R393 B.n329 B.n100 163.367
R394 B.n437 B.n64 163.367
R395 B.n433 B.n64 163.367
R396 B.n433 B.n432 163.367
R397 B.n432 B.n431 163.367
R398 B.n431 B.n66 163.367
R399 B.n427 B.n66 163.367
R400 B.n427 B.n426 163.367
R401 B.n426 B.n425 163.367
R402 B.n425 B.n68 163.367
R403 B.n421 B.n68 163.367
R404 B.n421 B.n420 163.367
R405 B.n420 B.n419 163.367
R406 B.n419 B.n70 163.367
R407 B.n415 B.n70 163.367
R408 B.n415 B.n414 163.367
R409 B.n414 B.n413 163.367
R410 B.n413 B.n72 163.367
R411 B.n409 B.n72 163.367
R412 B.n409 B.n408 163.367
R413 B.n408 B.n407 163.367
R414 B.n407 B.n74 163.367
R415 B.n403 B.n74 163.367
R416 B.n403 B.n402 163.367
R417 B.n402 B.n401 163.367
R418 B.n401 B.n76 163.367
R419 B.n397 B.n76 163.367
R420 B.n397 B.n396 163.367
R421 B.n396 B.n395 163.367
R422 B.n395 B.n78 163.367
R423 B.n391 B.n78 163.367
R424 B.n391 B.n390 163.367
R425 B.n390 B.n389 163.367
R426 B.n389 B.n80 163.367
R427 B.n385 B.n80 163.367
R428 B.n385 B.n384 163.367
R429 B.n384 B.n383 163.367
R430 B.n383 B.n82 163.367
R431 B.n379 B.n82 163.367
R432 B.n379 B.n378 163.367
R433 B.n378 B.n377 163.367
R434 B.n377 B.n84 163.367
R435 B.n373 B.n84 163.367
R436 B.n373 B.n372 163.367
R437 B.n372 B.n371 163.367
R438 B.n371 B.n86 163.367
R439 B.n367 B.n86 163.367
R440 B.n367 B.n366 163.367
R441 B.n366 B.n365 163.367
R442 B.n365 B.n88 163.367
R443 B.n361 B.n88 163.367
R444 B.n361 B.n360 163.367
R445 B.n360 B.n359 163.367
R446 B.n359 B.n90 163.367
R447 B.n355 B.n90 163.367
R448 B.n355 B.n354 163.367
R449 B.n354 B.n353 163.367
R450 B.n353 B.n92 163.367
R451 B.n349 B.n92 163.367
R452 B.n349 B.n348 163.367
R453 B.n348 B.n347 163.367
R454 B.n347 B.n94 163.367
R455 B.n343 B.n94 163.367
R456 B.n343 B.n342 163.367
R457 B.n342 B.n341 163.367
R458 B.n341 B.n96 163.367
R459 B.n337 B.n96 163.367
R460 B.n337 B.n336 163.367
R461 B.n336 B.n335 163.367
R462 B.n335 B.n98 163.367
R463 B.n331 B.n98 163.367
R464 B.n331 B.n330 163.367
R465 B.n554 B.n553 163.367
R466 B.n553 B.n552 163.367
R467 B.n552 B.n21 163.367
R468 B.n548 B.n21 163.367
R469 B.n548 B.n547 163.367
R470 B.n547 B.n546 163.367
R471 B.n546 B.n23 163.367
R472 B.n542 B.n23 163.367
R473 B.n542 B.n541 163.367
R474 B.n541 B.n540 163.367
R475 B.n540 B.n25 163.367
R476 B.n536 B.n25 163.367
R477 B.n536 B.n535 163.367
R478 B.n535 B.n534 163.367
R479 B.n534 B.n27 163.367
R480 B.n530 B.n27 163.367
R481 B.n530 B.n529 163.367
R482 B.n529 B.n528 163.367
R483 B.n528 B.n29 163.367
R484 B.n524 B.n29 163.367
R485 B.n524 B.n523 163.367
R486 B.n523 B.n522 163.367
R487 B.n522 B.n31 163.367
R488 B.n518 B.n31 163.367
R489 B.n518 B.n517 163.367
R490 B.n517 B.n516 163.367
R491 B.n516 B.n33 163.367
R492 B.n512 B.n33 163.367
R493 B.n512 B.n511 163.367
R494 B.n511 B.n510 163.367
R495 B.n510 B.n35 163.367
R496 B.n506 B.n35 163.367
R497 B.n506 B.n505 163.367
R498 B.n505 B.n504 163.367
R499 B.n504 B.n37 163.367
R500 B.n500 B.n37 163.367
R501 B.n500 B.n499 163.367
R502 B.n499 B.n498 163.367
R503 B.n498 B.n42 163.367
R504 B.n494 B.n42 163.367
R505 B.n494 B.n493 163.367
R506 B.n493 B.n492 163.367
R507 B.n492 B.n44 163.367
R508 B.n487 B.n44 163.367
R509 B.n487 B.n486 163.367
R510 B.n486 B.n485 163.367
R511 B.n485 B.n48 163.367
R512 B.n481 B.n48 163.367
R513 B.n481 B.n480 163.367
R514 B.n480 B.n479 163.367
R515 B.n479 B.n50 163.367
R516 B.n475 B.n50 163.367
R517 B.n475 B.n474 163.367
R518 B.n474 B.n473 163.367
R519 B.n473 B.n52 163.367
R520 B.n469 B.n52 163.367
R521 B.n469 B.n468 163.367
R522 B.n468 B.n467 163.367
R523 B.n467 B.n54 163.367
R524 B.n463 B.n54 163.367
R525 B.n463 B.n462 163.367
R526 B.n462 B.n461 163.367
R527 B.n461 B.n56 163.367
R528 B.n457 B.n56 163.367
R529 B.n457 B.n456 163.367
R530 B.n456 B.n455 163.367
R531 B.n455 B.n58 163.367
R532 B.n451 B.n58 163.367
R533 B.n451 B.n450 163.367
R534 B.n450 B.n449 163.367
R535 B.n449 B.n60 163.367
R536 B.n445 B.n60 163.367
R537 B.n445 B.n444 163.367
R538 B.n444 B.n443 163.367
R539 B.n443 B.n62 163.367
R540 B.n439 B.n62 163.367
R541 B.n439 B.n438 163.367
R542 B.n558 B.n19 163.367
R543 B.n559 B.n558 163.367
R544 B.n560 B.n559 163.367
R545 B.n560 B.n17 163.367
R546 B.n564 B.n17 163.367
R547 B.n565 B.n564 163.367
R548 B.n566 B.n565 163.367
R549 B.n566 B.n15 163.367
R550 B.n570 B.n15 163.367
R551 B.n571 B.n570 163.367
R552 B.n572 B.n571 163.367
R553 B.n572 B.n13 163.367
R554 B.n576 B.n13 163.367
R555 B.n577 B.n576 163.367
R556 B.n578 B.n577 163.367
R557 B.n578 B.n11 163.367
R558 B.n582 B.n11 163.367
R559 B.n583 B.n582 163.367
R560 B.n584 B.n583 163.367
R561 B.n584 B.n9 163.367
R562 B.n588 B.n9 163.367
R563 B.n589 B.n588 163.367
R564 B.n590 B.n589 163.367
R565 B.n590 B.n7 163.367
R566 B.n594 B.n7 163.367
R567 B.n595 B.n594 163.367
R568 B.n596 B.n595 163.367
R569 B.n596 B.n5 163.367
R570 B.n600 B.n5 163.367
R571 B.n601 B.n600 163.367
R572 B.n602 B.n601 163.367
R573 B.n602 B.n3 163.367
R574 B.n606 B.n3 163.367
R575 B.n607 B.n606 163.367
R576 B.n158 B.n2 163.367
R577 B.n159 B.n158 163.367
R578 B.n159 B.n156 163.367
R579 B.n163 B.n156 163.367
R580 B.n164 B.n163 163.367
R581 B.n165 B.n164 163.367
R582 B.n165 B.n154 163.367
R583 B.n169 B.n154 163.367
R584 B.n170 B.n169 163.367
R585 B.n171 B.n170 163.367
R586 B.n171 B.n152 163.367
R587 B.n175 B.n152 163.367
R588 B.n176 B.n175 163.367
R589 B.n177 B.n176 163.367
R590 B.n177 B.n150 163.367
R591 B.n181 B.n150 163.367
R592 B.n182 B.n181 163.367
R593 B.n183 B.n182 163.367
R594 B.n183 B.n148 163.367
R595 B.n187 B.n148 163.367
R596 B.n188 B.n187 163.367
R597 B.n189 B.n188 163.367
R598 B.n189 B.n146 163.367
R599 B.n193 B.n146 163.367
R600 B.n194 B.n193 163.367
R601 B.n195 B.n194 163.367
R602 B.n195 B.n144 163.367
R603 B.n199 B.n144 163.367
R604 B.n200 B.n199 163.367
R605 B.n201 B.n200 163.367
R606 B.n201 B.n142 163.367
R607 B.n205 B.n142 163.367
R608 B.n206 B.n205 163.367
R609 B.n207 B.n206 163.367
R610 B.n259 B.n258 59.7338
R611 B.n118 B.n117 59.7338
R612 B.n46 B.n45 59.7338
R613 B.n39 B.n38 59.7338
R614 B.n260 B.n259 59.5399
R615 B.n278 B.n118 59.5399
R616 B.n489 B.n46 59.5399
R617 B.n40 B.n39 59.5399
R618 B.n556 B.n555 31.0639
R619 B.n436 B.n63 31.0639
R620 B.n328 B.n99 31.0639
R621 B.n209 B.n208 31.0639
R622 B B.n609 18.0485
R623 B.n557 B.n556 10.6151
R624 B.n557 B.n18 10.6151
R625 B.n561 B.n18 10.6151
R626 B.n562 B.n561 10.6151
R627 B.n563 B.n562 10.6151
R628 B.n563 B.n16 10.6151
R629 B.n567 B.n16 10.6151
R630 B.n568 B.n567 10.6151
R631 B.n569 B.n568 10.6151
R632 B.n569 B.n14 10.6151
R633 B.n573 B.n14 10.6151
R634 B.n574 B.n573 10.6151
R635 B.n575 B.n574 10.6151
R636 B.n575 B.n12 10.6151
R637 B.n579 B.n12 10.6151
R638 B.n580 B.n579 10.6151
R639 B.n581 B.n580 10.6151
R640 B.n581 B.n10 10.6151
R641 B.n585 B.n10 10.6151
R642 B.n586 B.n585 10.6151
R643 B.n587 B.n586 10.6151
R644 B.n587 B.n8 10.6151
R645 B.n591 B.n8 10.6151
R646 B.n592 B.n591 10.6151
R647 B.n593 B.n592 10.6151
R648 B.n593 B.n6 10.6151
R649 B.n597 B.n6 10.6151
R650 B.n598 B.n597 10.6151
R651 B.n599 B.n598 10.6151
R652 B.n599 B.n4 10.6151
R653 B.n603 B.n4 10.6151
R654 B.n604 B.n603 10.6151
R655 B.n605 B.n604 10.6151
R656 B.n605 B.n0 10.6151
R657 B.n555 B.n20 10.6151
R658 B.n551 B.n20 10.6151
R659 B.n551 B.n550 10.6151
R660 B.n550 B.n549 10.6151
R661 B.n549 B.n22 10.6151
R662 B.n545 B.n22 10.6151
R663 B.n545 B.n544 10.6151
R664 B.n544 B.n543 10.6151
R665 B.n543 B.n24 10.6151
R666 B.n539 B.n24 10.6151
R667 B.n539 B.n538 10.6151
R668 B.n538 B.n537 10.6151
R669 B.n537 B.n26 10.6151
R670 B.n533 B.n26 10.6151
R671 B.n533 B.n532 10.6151
R672 B.n532 B.n531 10.6151
R673 B.n531 B.n28 10.6151
R674 B.n527 B.n28 10.6151
R675 B.n527 B.n526 10.6151
R676 B.n526 B.n525 10.6151
R677 B.n525 B.n30 10.6151
R678 B.n521 B.n30 10.6151
R679 B.n521 B.n520 10.6151
R680 B.n520 B.n519 10.6151
R681 B.n519 B.n32 10.6151
R682 B.n515 B.n32 10.6151
R683 B.n515 B.n514 10.6151
R684 B.n514 B.n513 10.6151
R685 B.n513 B.n34 10.6151
R686 B.n509 B.n34 10.6151
R687 B.n509 B.n508 10.6151
R688 B.n508 B.n507 10.6151
R689 B.n507 B.n36 10.6151
R690 B.n503 B.n502 10.6151
R691 B.n502 B.n501 10.6151
R692 B.n501 B.n41 10.6151
R693 B.n497 B.n41 10.6151
R694 B.n497 B.n496 10.6151
R695 B.n496 B.n495 10.6151
R696 B.n495 B.n43 10.6151
R697 B.n491 B.n43 10.6151
R698 B.n491 B.n490 10.6151
R699 B.n488 B.n47 10.6151
R700 B.n484 B.n47 10.6151
R701 B.n484 B.n483 10.6151
R702 B.n483 B.n482 10.6151
R703 B.n482 B.n49 10.6151
R704 B.n478 B.n49 10.6151
R705 B.n478 B.n477 10.6151
R706 B.n477 B.n476 10.6151
R707 B.n476 B.n51 10.6151
R708 B.n472 B.n51 10.6151
R709 B.n472 B.n471 10.6151
R710 B.n471 B.n470 10.6151
R711 B.n470 B.n53 10.6151
R712 B.n466 B.n53 10.6151
R713 B.n466 B.n465 10.6151
R714 B.n465 B.n464 10.6151
R715 B.n464 B.n55 10.6151
R716 B.n460 B.n55 10.6151
R717 B.n460 B.n459 10.6151
R718 B.n459 B.n458 10.6151
R719 B.n458 B.n57 10.6151
R720 B.n454 B.n57 10.6151
R721 B.n454 B.n453 10.6151
R722 B.n453 B.n452 10.6151
R723 B.n452 B.n59 10.6151
R724 B.n448 B.n59 10.6151
R725 B.n448 B.n447 10.6151
R726 B.n447 B.n446 10.6151
R727 B.n446 B.n61 10.6151
R728 B.n442 B.n61 10.6151
R729 B.n442 B.n441 10.6151
R730 B.n441 B.n440 10.6151
R731 B.n440 B.n63 10.6151
R732 B.n436 B.n435 10.6151
R733 B.n435 B.n434 10.6151
R734 B.n434 B.n65 10.6151
R735 B.n430 B.n65 10.6151
R736 B.n430 B.n429 10.6151
R737 B.n429 B.n428 10.6151
R738 B.n428 B.n67 10.6151
R739 B.n424 B.n67 10.6151
R740 B.n424 B.n423 10.6151
R741 B.n423 B.n422 10.6151
R742 B.n422 B.n69 10.6151
R743 B.n418 B.n69 10.6151
R744 B.n418 B.n417 10.6151
R745 B.n417 B.n416 10.6151
R746 B.n416 B.n71 10.6151
R747 B.n412 B.n71 10.6151
R748 B.n412 B.n411 10.6151
R749 B.n411 B.n410 10.6151
R750 B.n410 B.n73 10.6151
R751 B.n406 B.n73 10.6151
R752 B.n406 B.n405 10.6151
R753 B.n405 B.n404 10.6151
R754 B.n404 B.n75 10.6151
R755 B.n400 B.n75 10.6151
R756 B.n400 B.n399 10.6151
R757 B.n399 B.n398 10.6151
R758 B.n398 B.n77 10.6151
R759 B.n394 B.n77 10.6151
R760 B.n394 B.n393 10.6151
R761 B.n393 B.n392 10.6151
R762 B.n392 B.n79 10.6151
R763 B.n388 B.n79 10.6151
R764 B.n388 B.n387 10.6151
R765 B.n387 B.n386 10.6151
R766 B.n386 B.n81 10.6151
R767 B.n382 B.n81 10.6151
R768 B.n382 B.n381 10.6151
R769 B.n381 B.n380 10.6151
R770 B.n380 B.n83 10.6151
R771 B.n376 B.n83 10.6151
R772 B.n376 B.n375 10.6151
R773 B.n375 B.n374 10.6151
R774 B.n374 B.n85 10.6151
R775 B.n370 B.n85 10.6151
R776 B.n370 B.n369 10.6151
R777 B.n369 B.n368 10.6151
R778 B.n368 B.n87 10.6151
R779 B.n364 B.n87 10.6151
R780 B.n364 B.n363 10.6151
R781 B.n363 B.n362 10.6151
R782 B.n362 B.n89 10.6151
R783 B.n358 B.n89 10.6151
R784 B.n358 B.n357 10.6151
R785 B.n357 B.n356 10.6151
R786 B.n356 B.n91 10.6151
R787 B.n352 B.n91 10.6151
R788 B.n352 B.n351 10.6151
R789 B.n351 B.n350 10.6151
R790 B.n350 B.n93 10.6151
R791 B.n346 B.n93 10.6151
R792 B.n346 B.n345 10.6151
R793 B.n345 B.n344 10.6151
R794 B.n344 B.n95 10.6151
R795 B.n340 B.n95 10.6151
R796 B.n340 B.n339 10.6151
R797 B.n339 B.n338 10.6151
R798 B.n338 B.n97 10.6151
R799 B.n334 B.n97 10.6151
R800 B.n334 B.n333 10.6151
R801 B.n333 B.n332 10.6151
R802 B.n332 B.n99 10.6151
R803 B.n157 B.n1 10.6151
R804 B.n160 B.n157 10.6151
R805 B.n161 B.n160 10.6151
R806 B.n162 B.n161 10.6151
R807 B.n162 B.n155 10.6151
R808 B.n166 B.n155 10.6151
R809 B.n167 B.n166 10.6151
R810 B.n168 B.n167 10.6151
R811 B.n168 B.n153 10.6151
R812 B.n172 B.n153 10.6151
R813 B.n173 B.n172 10.6151
R814 B.n174 B.n173 10.6151
R815 B.n174 B.n151 10.6151
R816 B.n178 B.n151 10.6151
R817 B.n179 B.n178 10.6151
R818 B.n180 B.n179 10.6151
R819 B.n180 B.n149 10.6151
R820 B.n184 B.n149 10.6151
R821 B.n185 B.n184 10.6151
R822 B.n186 B.n185 10.6151
R823 B.n186 B.n147 10.6151
R824 B.n190 B.n147 10.6151
R825 B.n191 B.n190 10.6151
R826 B.n192 B.n191 10.6151
R827 B.n192 B.n145 10.6151
R828 B.n196 B.n145 10.6151
R829 B.n197 B.n196 10.6151
R830 B.n198 B.n197 10.6151
R831 B.n198 B.n143 10.6151
R832 B.n202 B.n143 10.6151
R833 B.n203 B.n202 10.6151
R834 B.n204 B.n203 10.6151
R835 B.n204 B.n141 10.6151
R836 B.n208 B.n141 10.6151
R837 B.n210 B.n209 10.6151
R838 B.n210 B.n139 10.6151
R839 B.n214 B.n139 10.6151
R840 B.n215 B.n214 10.6151
R841 B.n216 B.n215 10.6151
R842 B.n216 B.n137 10.6151
R843 B.n220 B.n137 10.6151
R844 B.n221 B.n220 10.6151
R845 B.n222 B.n221 10.6151
R846 B.n222 B.n135 10.6151
R847 B.n226 B.n135 10.6151
R848 B.n227 B.n226 10.6151
R849 B.n228 B.n227 10.6151
R850 B.n228 B.n133 10.6151
R851 B.n232 B.n133 10.6151
R852 B.n233 B.n232 10.6151
R853 B.n234 B.n233 10.6151
R854 B.n234 B.n131 10.6151
R855 B.n238 B.n131 10.6151
R856 B.n239 B.n238 10.6151
R857 B.n240 B.n239 10.6151
R858 B.n240 B.n129 10.6151
R859 B.n244 B.n129 10.6151
R860 B.n245 B.n244 10.6151
R861 B.n246 B.n245 10.6151
R862 B.n246 B.n127 10.6151
R863 B.n250 B.n127 10.6151
R864 B.n251 B.n250 10.6151
R865 B.n252 B.n251 10.6151
R866 B.n252 B.n125 10.6151
R867 B.n256 B.n125 10.6151
R868 B.n257 B.n256 10.6151
R869 B.n261 B.n257 10.6151
R870 B.n265 B.n123 10.6151
R871 B.n266 B.n265 10.6151
R872 B.n267 B.n266 10.6151
R873 B.n267 B.n121 10.6151
R874 B.n271 B.n121 10.6151
R875 B.n272 B.n271 10.6151
R876 B.n273 B.n272 10.6151
R877 B.n273 B.n119 10.6151
R878 B.n277 B.n119 10.6151
R879 B.n280 B.n279 10.6151
R880 B.n280 B.n115 10.6151
R881 B.n284 B.n115 10.6151
R882 B.n285 B.n284 10.6151
R883 B.n286 B.n285 10.6151
R884 B.n286 B.n113 10.6151
R885 B.n290 B.n113 10.6151
R886 B.n291 B.n290 10.6151
R887 B.n292 B.n291 10.6151
R888 B.n292 B.n111 10.6151
R889 B.n296 B.n111 10.6151
R890 B.n297 B.n296 10.6151
R891 B.n298 B.n297 10.6151
R892 B.n298 B.n109 10.6151
R893 B.n302 B.n109 10.6151
R894 B.n303 B.n302 10.6151
R895 B.n304 B.n303 10.6151
R896 B.n304 B.n107 10.6151
R897 B.n308 B.n107 10.6151
R898 B.n309 B.n308 10.6151
R899 B.n310 B.n309 10.6151
R900 B.n310 B.n105 10.6151
R901 B.n314 B.n105 10.6151
R902 B.n315 B.n314 10.6151
R903 B.n316 B.n315 10.6151
R904 B.n316 B.n103 10.6151
R905 B.n320 B.n103 10.6151
R906 B.n321 B.n320 10.6151
R907 B.n322 B.n321 10.6151
R908 B.n322 B.n101 10.6151
R909 B.n326 B.n101 10.6151
R910 B.n327 B.n326 10.6151
R911 B.n328 B.n327 10.6151
R912 B.n40 B.n36 9.36635
R913 B.n489 B.n488 9.36635
R914 B.n261 B.n260 9.36635
R915 B.n279 B.n278 9.36635
R916 B.n609 B.n0 8.11757
R917 B.n609 B.n1 8.11757
R918 B.n503 B.n40 1.24928
R919 B.n490 B.n489 1.24928
R920 B.n260 B.n123 1.24928
R921 B.n278 B.n277 1.24928
R922 VN.n0 VN.t3 117.838
R923 VN.n1 VN.t1 117.838
R924 VN.n0 VN.t0 116.959
R925 VN.n1 VN.t2 116.959
R926 VN VN.n1 48.6824
R927 VN VN.n0 3.58008
R928 VTAIL.n410 VTAIL.n364 756.745
R929 VTAIL.n46 VTAIL.n0 756.745
R930 VTAIL.n98 VTAIL.n52 756.745
R931 VTAIL.n150 VTAIL.n104 756.745
R932 VTAIL.n358 VTAIL.n312 756.745
R933 VTAIL.n306 VTAIL.n260 756.745
R934 VTAIL.n254 VTAIL.n208 756.745
R935 VTAIL.n202 VTAIL.n156 756.745
R936 VTAIL.n380 VTAIL.n379 585
R937 VTAIL.n385 VTAIL.n384 585
R938 VTAIL.n387 VTAIL.n386 585
R939 VTAIL.n376 VTAIL.n375 585
R940 VTAIL.n393 VTAIL.n392 585
R941 VTAIL.n395 VTAIL.n394 585
R942 VTAIL.n372 VTAIL.n371 585
R943 VTAIL.n401 VTAIL.n400 585
R944 VTAIL.n403 VTAIL.n402 585
R945 VTAIL.n368 VTAIL.n367 585
R946 VTAIL.n409 VTAIL.n408 585
R947 VTAIL.n411 VTAIL.n410 585
R948 VTAIL.n16 VTAIL.n15 585
R949 VTAIL.n21 VTAIL.n20 585
R950 VTAIL.n23 VTAIL.n22 585
R951 VTAIL.n12 VTAIL.n11 585
R952 VTAIL.n29 VTAIL.n28 585
R953 VTAIL.n31 VTAIL.n30 585
R954 VTAIL.n8 VTAIL.n7 585
R955 VTAIL.n37 VTAIL.n36 585
R956 VTAIL.n39 VTAIL.n38 585
R957 VTAIL.n4 VTAIL.n3 585
R958 VTAIL.n45 VTAIL.n44 585
R959 VTAIL.n47 VTAIL.n46 585
R960 VTAIL.n68 VTAIL.n67 585
R961 VTAIL.n73 VTAIL.n72 585
R962 VTAIL.n75 VTAIL.n74 585
R963 VTAIL.n64 VTAIL.n63 585
R964 VTAIL.n81 VTAIL.n80 585
R965 VTAIL.n83 VTAIL.n82 585
R966 VTAIL.n60 VTAIL.n59 585
R967 VTAIL.n89 VTAIL.n88 585
R968 VTAIL.n91 VTAIL.n90 585
R969 VTAIL.n56 VTAIL.n55 585
R970 VTAIL.n97 VTAIL.n96 585
R971 VTAIL.n99 VTAIL.n98 585
R972 VTAIL.n120 VTAIL.n119 585
R973 VTAIL.n125 VTAIL.n124 585
R974 VTAIL.n127 VTAIL.n126 585
R975 VTAIL.n116 VTAIL.n115 585
R976 VTAIL.n133 VTAIL.n132 585
R977 VTAIL.n135 VTAIL.n134 585
R978 VTAIL.n112 VTAIL.n111 585
R979 VTAIL.n141 VTAIL.n140 585
R980 VTAIL.n143 VTAIL.n142 585
R981 VTAIL.n108 VTAIL.n107 585
R982 VTAIL.n149 VTAIL.n148 585
R983 VTAIL.n151 VTAIL.n150 585
R984 VTAIL.n359 VTAIL.n358 585
R985 VTAIL.n357 VTAIL.n356 585
R986 VTAIL.n316 VTAIL.n315 585
R987 VTAIL.n351 VTAIL.n350 585
R988 VTAIL.n349 VTAIL.n348 585
R989 VTAIL.n320 VTAIL.n319 585
R990 VTAIL.n343 VTAIL.n342 585
R991 VTAIL.n341 VTAIL.n340 585
R992 VTAIL.n324 VTAIL.n323 585
R993 VTAIL.n335 VTAIL.n334 585
R994 VTAIL.n333 VTAIL.n332 585
R995 VTAIL.n328 VTAIL.n327 585
R996 VTAIL.n307 VTAIL.n306 585
R997 VTAIL.n305 VTAIL.n304 585
R998 VTAIL.n264 VTAIL.n263 585
R999 VTAIL.n299 VTAIL.n298 585
R1000 VTAIL.n297 VTAIL.n296 585
R1001 VTAIL.n268 VTAIL.n267 585
R1002 VTAIL.n291 VTAIL.n290 585
R1003 VTAIL.n289 VTAIL.n288 585
R1004 VTAIL.n272 VTAIL.n271 585
R1005 VTAIL.n283 VTAIL.n282 585
R1006 VTAIL.n281 VTAIL.n280 585
R1007 VTAIL.n276 VTAIL.n275 585
R1008 VTAIL.n255 VTAIL.n254 585
R1009 VTAIL.n253 VTAIL.n252 585
R1010 VTAIL.n212 VTAIL.n211 585
R1011 VTAIL.n247 VTAIL.n246 585
R1012 VTAIL.n245 VTAIL.n244 585
R1013 VTAIL.n216 VTAIL.n215 585
R1014 VTAIL.n239 VTAIL.n238 585
R1015 VTAIL.n237 VTAIL.n236 585
R1016 VTAIL.n220 VTAIL.n219 585
R1017 VTAIL.n231 VTAIL.n230 585
R1018 VTAIL.n229 VTAIL.n228 585
R1019 VTAIL.n224 VTAIL.n223 585
R1020 VTAIL.n203 VTAIL.n202 585
R1021 VTAIL.n201 VTAIL.n200 585
R1022 VTAIL.n160 VTAIL.n159 585
R1023 VTAIL.n195 VTAIL.n194 585
R1024 VTAIL.n193 VTAIL.n192 585
R1025 VTAIL.n164 VTAIL.n163 585
R1026 VTAIL.n187 VTAIL.n186 585
R1027 VTAIL.n185 VTAIL.n184 585
R1028 VTAIL.n168 VTAIL.n167 585
R1029 VTAIL.n179 VTAIL.n178 585
R1030 VTAIL.n177 VTAIL.n176 585
R1031 VTAIL.n172 VTAIL.n171 585
R1032 VTAIL.n381 VTAIL.t5 327.467
R1033 VTAIL.n17 VTAIL.t4 327.467
R1034 VTAIL.n69 VTAIL.t3 327.467
R1035 VTAIL.n121 VTAIL.t0 327.467
R1036 VTAIL.n277 VTAIL.t2 327.467
R1037 VTAIL.n225 VTAIL.t7 327.467
R1038 VTAIL.n173 VTAIL.t6 327.467
R1039 VTAIL.n329 VTAIL.t1 327.467
R1040 VTAIL.n385 VTAIL.n379 171.744
R1041 VTAIL.n386 VTAIL.n385 171.744
R1042 VTAIL.n386 VTAIL.n375 171.744
R1043 VTAIL.n393 VTAIL.n375 171.744
R1044 VTAIL.n394 VTAIL.n393 171.744
R1045 VTAIL.n394 VTAIL.n371 171.744
R1046 VTAIL.n401 VTAIL.n371 171.744
R1047 VTAIL.n402 VTAIL.n401 171.744
R1048 VTAIL.n402 VTAIL.n367 171.744
R1049 VTAIL.n409 VTAIL.n367 171.744
R1050 VTAIL.n410 VTAIL.n409 171.744
R1051 VTAIL.n21 VTAIL.n15 171.744
R1052 VTAIL.n22 VTAIL.n21 171.744
R1053 VTAIL.n22 VTAIL.n11 171.744
R1054 VTAIL.n29 VTAIL.n11 171.744
R1055 VTAIL.n30 VTAIL.n29 171.744
R1056 VTAIL.n30 VTAIL.n7 171.744
R1057 VTAIL.n37 VTAIL.n7 171.744
R1058 VTAIL.n38 VTAIL.n37 171.744
R1059 VTAIL.n38 VTAIL.n3 171.744
R1060 VTAIL.n45 VTAIL.n3 171.744
R1061 VTAIL.n46 VTAIL.n45 171.744
R1062 VTAIL.n73 VTAIL.n67 171.744
R1063 VTAIL.n74 VTAIL.n73 171.744
R1064 VTAIL.n74 VTAIL.n63 171.744
R1065 VTAIL.n81 VTAIL.n63 171.744
R1066 VTAIL.n82 VTAIL.n81 171.744
R1067 VTAIL.n82 VTAIL.n59 171.744
R1068 VTAIL.n89 VTAIL.n59 171.744
R1069 VTAIL.n90 VTAIL.n89 171.744
R1070 VTAIL.n90 VTAIL.n55 171.744
R1071 VTAIL.n97 VTAIL.n55 171.744
R1072 VTAIL.n98 VTAIL.n97 171.744
R1073 VTAIL.n125 VTAIL.n119 171.744
R1074 VTAIL.n126 VTAIL.n125 171.744
R1075 VTAIL.n126 VTAIL.n115 171.744
R1076 VTAIL.n133 VTAIL.n115 171.744
R1077 VTAIL.n134 VTAIL.n133 171.744
R1078 VTAIL.n134 VTAIL.n111 171.744
R1079 VTAIL.n141 VTAIL.n111 171.744
R1080 VTAIL.n142 VTAIL.n141 171.744
R1081 VTAIL.n142 VTAIL.n107 171.744
R1082 VTAIL.n149 VTAIL.n107 171.744
R1083 VTAIL.n150 VTAIL.n149 171.744
R1084 VTAIL.n358 VTAIL.n357 171.744
R1085 VTAIL.n357 VTAIL.n315 171.744
R1086 VTAIL.n350 VTAIL.n315 171.744
R1087 VTAIL.n350 VTAIL.n349 171.744
R1088 VTAIL.n349 VTAIL.n319 171.744
R1089 VTAIL.n342 VTAIL.n319 171.744
R1090 VTAIL.n342 VTAIL.n341 171.744
R1091 VTAIL.n341 VTAIL.n323 171.744
R1092 VTAIL.n334 VTAIL.n323 171.744
R1093 VTAIL.n334 VTAIL.n333 171.744
R1094 VTAIL.n333 VTAIL.n327 171.744
R1095 VTAIL.n306 VTAIL.n305 171.744
R1096 VTAIL.n305 VTAIL.n263 171.744
R1097 VTAIL.n298 VTAIL.n263 171.744
R1098 VTAIL.n298 VTAIL.n297 171.744
R1099 VTAIL.n297 VTAIL.n267 171.744
R1100 VTAIL.n290 VTAIL.n267 171.744
R1101 VTAIL.n290 VTAIL.n289 171.744
R1102 VTAIL.n289 VTAIL.n271 171.744
R1103 VTAIL.n282 VTAIL.n271 171.744
R1104 VTAIL.n282 VTAIL.n281 171.744
R1105 VTAIL.n281 VTAIL.n275 171.744
R1106 VTAIL.n254 VTAIL.n253 171.744
R1107 VTAIL.n253 VTAIL.n211 171.744
R1108 VTAIL.n246 VTAIL.n211 171.744
R1109 VTAIL.n246 VTAIL.n245 171.744
R1110 VTAIL.n245 VTAIL.n215 171.744
R1111 VTAIL.n238 VTAIL.n215 171.744
R1112 VTAIL.n238 VTAIL.n237 171.744
R1113 VTAIL.n237 VTAIL.n219 171.744
R1114 VTAIL.n230 VTAIL.n219 171.744
R1115 VTAIL.n230 VTAIL.n229 171.744
R1116 VTAIL.n229 VTAIL.n223 171.744
R1117 VTAIL.n202 VTAIL.n201 171.744
R1118 VTAIL.n201 VTAIL.n159 171.744
R1119 VTAIL.n194 VTAIL.n159 171.744
R1120 VTAIL.n194 VTAIL.n193 171.744
R1121 VTAIL.n193 VTAIL.n163 171.744
R1122 VTAIL.n186 VTAIL.n163 171.744
R1123 VTAIL.n186 VTAIL.n185 171.744
R1124 VTAIL.n185 VTAIL.n167 171.744
R1125 VTAIL.n178 VTAIL.n167 171.744
R1126 VTAIL.n178 VTAIL.n177 171.744
R1127 VTAIL.n177 VTAIL.n171 171.744
R1128 VTAIL.t5 VTAIL.n379 85.8723
R1129 VTAIL.t4 VTAIL.n15 85.8723
R1130 VTAIL.t3 VTAIL.n67 85.8723
R1131 VTAIL.t0 VTAIL.n119 85.8723
R1132 VTAIL.t1 VTAIL.n327 85.8723
R1133 VTAIL.t2 VTAIL.n275 85.8723
R1134 VTAIL.t7 VTAIL.n223 85.8723
R1135 VTAIL.t6 VTAIL.n171 85.8723
R1136 VTAIL.n415 VTAIL.n414 30.4399
R1137 VTAIL.n51 VTAIL.n50 30.4399
R1138 VTAIL.n103 VTAIL.n102 30.4399
R1139 VTAIL.n155 VTAIL.n154 30.4399
R1140 VTAIL.n363 VTAIL.n362 30.4399
R1141 VTAIL.n311 VTAIL.n310 30.4399
R1142 VTAIL.n259 VTAIL.n258 30.4399
R1143 VTAIL.n207 VTAIL.n206 30.4399
R1144 VTAIL.n415 VTAIL.n363 23.2203
R1145 VTAIL.n207 VTAIL.n155 23.2203
R1146 VTAIL.n381 VTAIL.n380 16.3895
R1147 VTAIL.n17 VTAIL.n16 16.3895
R1148 VTAIL.n69 VTAIL.n68 16.3895
R1149 VTAIL.n121 VTAIL.n120 16.3895
R1150 VTAIL.n329 VTAIL.n328 16.3895
R1151 VTAIL.n277 VTAIL.n276 16.3895
R1152 VTAIL.n225 VTAIL.n224 16.3895
R1153 VTAIL.n173 VTAIL.n172 16.3895
R1154 VTAIL.n384 VTAIL.n383 12.8005
R1155 VTAIL.n20 VTAIL.n19 12.8005
R1156 VTAIL.n72 VTAIL.n71 12.8005
R1157 VTAIL.n124 VTAIL.n123 12.8005
R1158 VTAIL.n332 VTAIL.n331 12.8005
R1159 VTAIL.n280 VTAIL.n279 12.8005
R1160 VTAIL.n228 VTAIL.n227 12.8005
R1161 VTAIL.n176 VTAIL.n175 12.8005
R1162 VTAIL.n387 VTAIL.n378 12.0247
R1163 VTAIL.n23 VTAIL.n14 12.0247
R1164 VTAIL.n75 VTAIL.n66 12.0247
R1165 VTAIL.n127 VTAIL.n118 12.0247
R1166 VTAIL.n335 VTAIL.n326 12.0247
R1167 VTAIL.n283 VTAIL.n274 12.0247
R1168 VTAIL.n231 VTAIL.n222 12.0247
R1169 VTAIL.n179 VTAIL.n170 12.0247
R1170 VTAIL.n388 VTAIL.n376 11.249
R1171 VTAIL.n24 VTAIL.n12 11.249
R1172 VTAIL.n76 VTAIL.n64 11.249
R1173 VTAIL.n128 VTAIL.n116 11.249
R1174 VTAIL.n336 VTAIL.n324 11.249
R1175 VTAIL.n284 VTAIL.n272 11.249
R1176 VTAIL.n232 VTAIL.n220 11.249
R1177 VTAIL.n180 VTAIL.n168 11.249
R1178 VTAIL.n392 VTAIL.n391 10.4732
R1179 VTAIL.n28 VTAIL.n27 10.4732
R1180 VTAIL.n80 VTAIL.n79 10.4732
R1181 VTAIL.n132 VTAIL.n131 10.4732
R1182 VTAIL.n340 VTAIL.n339 10.4732
R1183 VTAIL.n288 VTAIL.n287 10.4732
R1184 VTAIL.n236 VTAIL.n235 10.4732
R1185 VTAIL.n184 VTAIL.n183 10.4732
R1186 VTAIL.n395 VTAIL.n374 9.69747
R1187 VTAIL.n414 VTAIL.n364 9.69747
R1188 VTAIL.n31 VTAIL.n10 9.69747
R1189 VTAIL.n50 VTAIL.n0 9.69747
R1190 VTAIL.n83 VTAIL.n62 9.69747
R1191 VTAIL.n102 VTAIL.n52 9.69747
R1192 VTAIL.n135 VTAIL.n114 9.69747
R1193 VTAIL.n154 VTAIL.n104 9.69747
R1194 VTAIL.n362 VTAIL.n312 9.69747
R1195 VTAIL.n343 VTAIL.n322 9.69747
R1196 VTAIL.n310 VTAIL.n260 9.69747
R1197 VTAIL.n291 VTAIL.n270 9.69747
R1198 VTAIL.n258 VTAIL.n208 9.69747
R1199 VTAIL.n239 VTAIL.n218 9.69747
R1200 VTAIL.n206 VTAIL.n156 9.69747
R1201 VTAIL.n187 VTAIL.n166 9.69747
R1202 VTAIL.n414 VTAIL.n413 9.45567
R1203 VTAIL.n50 VTAIL.n49 9.45567
R1204 VTAIL.n102 VTAIL.n101 9.45567
R1205 VTAIL.n154 VTAIL.n153 9.45567
R1206 VTAIL.n362 VTAIL.n361 9.45567
R1207 VTAIL.n310 VTAIL.n309 9.45567
R1208 VTAIL.n258 VTAIL.n257 9.45567
R1209 VTAIL.n206 VTAIL.n205 9.45567
R1210 VTAIL.n405 VTAIL.n404 9.3005
R1211 VTAIL.n407 VTAIL.n406 9.3005
R1212 VTAIL.n366 VTAIL.n365 9.3005
R1213 VTAIL.n413 VTAIL.n412 9.3005
R1214 VTAIL.n399 VTAIL.n398 9.3005
R1215 VTAIL.n397 VTAIL.n396 9.3005
R1216 VTAIL.n374 VTAIL.n373 9.3005
R1217 VTAIL.n391 VTAIL.n390 9.3005
R1218 VTAIL.n389 VTAIL.n388 9.3005
R1219 VTAIL.n378 VTAIL.n377 9.3005
R1220 VTAIL.n383 VTAIL.n382 9.3005
R1221 VTAIL.n370 VTAIL.n369 9.3005
R1222 VTAIL.n41 VTAIL.n40 9.3005
R1223 VTAIL.n43 VTAIL.n42 9.3005
R1224 VTAIL.n2 VTAIL.n1 9.3005
R1225 VTAIL.n49 VTAIL.n48 9.3005
R1226 VTAIL.n35 VTAIL.n34 9.3005
R1227 VTAIL.n33 VTAIL.n32 9.3005
R1228 VTAIL.n10 VTAIL.n9 9.3005
R1229 VTAIL.n27 VTAIL.n26 9.3005
R1230 VTAIL.n25 VTAIL.n24 9.3005
R1231 VTAIL.n14 VTAIL.n13 9.3005
R1232 VTAIL.n19 VTAIL.n18 9.3005
R1233 VTAIL.n6 VTAIL.n5 9.3005
R1234 VTAIL.n93 VTAIL.n92 9.3005
R1235 VTAIL.n95 VTAIL.n94 9.3005
R1236 VTAIL.n54 VTAIL.n53 9.3005
R1237 VTAIL.n101 VTAIL.n100 9.3005
R1238 VTAIL.n87 VTAIL.n86 9.3005
R1239 VTAIL.n85 VTAIL.n84 9.3005
R1240 VTAIL.n62 VTAIL.n61 9.3005
R1241 VTAIL.n79 VTAIL.n78 9.3005
R1242 VTAIL.n77 VTAIL.n76 9.3005
R1243 VTAIL.n66 VTAIL.n65 9.3005
R1244 VTAIL.n71 VTAIL.n70 9.3005
R1245 VTAIL.n58 VTAIL.n57 9.3005
R1246 VTAIL.n145 VTAIL.n144 9.3005
R1247 VTAIL.n147 VTAIL.n146 9.3005
R1248 VTAIL.n106 VTAIL.n105 9.3005
R1249 VTAIL.n153 VTAIL.n152 9.3005
R1250 VTAIL.n139 VTAIL.n138 9.3005
R1251 VTAIL.n137 VTAIL.n136 9.3005
R1252 VTAIL.n114 VTAIL.n113 9.3005
R1253 VTAIL.n131 VTAIL.n130 9.3005
R1254 VTAIL.n129 VTAIL.n128 9.3005
R1255 VTAIL.n118 VTAIL.n117 9.3005
R1256 VTAIL.n123 VTAIL.n122 9.3005
R1257 VTAIL.n110 VTAIL.n109 9.3005
R1258 VTAIL.n314 VTAIL.n313 9.3005
R1259 VTAIL.n355 VTAIL.n354 9.3005
R1260 VTAIL.n353 VTAIL.n352 9.3005
R1261 VTAIL.n318 VTAIL.n317 9.3005
R1262 VTAIL.n347 VTAIL.n346 9.3005
R1263 VTAIL.n345 VTAIL.n344 9.3005
R1264 VTAIL.n322 VTAIL.n321 9.3005
R1265 VTAIL.n339 VTAIL.n338 9.3005
R1266 VTAIL.n337 VTAIL.n336 9.3005
R1267 VTAIL.n326 VTAIL.n325 9.3005
R1268 VTAIL.n331 VTAIL.n330 9.3005
R1269 VTAIL.n361 VTAIL.n360 9.3005
R1270 VTAIL.n303 VTAIL.n302 9.3005
R1271 VTAIL.n262 VTAIL.n261 9.3005
R1272 VTAIL.n309 VTAIL.n308 9.3005
R1273 VTAIL.n301 VTAIL.n300 9.3005
R1274 VTAIL.n266 VTAIL.n265 9.3005
R1275 VTAIL.n295 VTAIL.n294 9.3005
R1276 VTAIL.n293 VTAIL.n292 9.3005
R1277 VTAIL.n270 VTAIL.n269 9.3005
R1278 VTAIL.n287 VTAIL.n286 9.3005
R1279 VTAIL.n285 VTAIL.n284 9.3005
R1280 VTAIL.n274 VTAIL.n273 9.3005
R1281 VTAIL.n279 VTAIL.n278 9.3005
R1282 VTAIL.n251 VTAIL.n250 9.3005
R1283 VTAIL.n210 VTAIL.n209 9.3005
R1284 VTAIL.n257 VTAIL.n256 9.3005
R1285 VTAIL.n249 VTAIL.n248 9.3005
R1286 VTAIL.n214 VTAIL.n213 9.3005
R1287 VTAIL.n243 VTAIL.n242 9.3005
R1288 VTAIL.n241 VTAIL.n240 9.3005
R1289 VTAIL.n218 VTAIL.n217 9.3005
R1290 VTAIL.n235 VTAIL.n234 9.3005
R1291 VTAIL.n233 VTAIL.n232 9.3005
R1292 VTAIL.n222 VTAIL.n221 9.3005
R1293 VTAIL.n227 VTAIL.n226 9.3005
R1294 VTAIL.n199 VTAIL.n198 9.3005
R1295 VTAIL.n158 VTAIL.n157 9.3005
R1296 VTAIL.n205 VTAIL.n204 9.3005
R1297 VTAIL.n197 VTAIL.n196 9.3005
R1298 VTAIL.n162 VTAIL.n161 9.3005
R1299 VTAIL.n191 VTAIL.n190 9.3005
R1300 VTAIL.n189 VTAIL.n188 9.3005
R1301 VTAIL.n166 VTAIL.n165 9.3005
R1302 VTAIL.n183 VTAIL.n182 9.3005
R1303 VTAIL.n181 VTAIL.n180 9.3005
R1304 VTAIL.n170 VTAIL.n169 9.3005
R1305 VTAIL.n175 VTAIL.n174 9.3005
R1306 VTAIL.n396 VTAIL.n372 8.92171
R1307 VTAIL.n412 VTAIL.n411 8.92171
R1308 VTAIL.n32 VTAIL.n8 8.92171
R1309 VTAIL.n48 VTAIL.n47 8.92171
R1310 VTAIL.n84 VTAIL.n60 8.92171
R1311 VTAIL.n100 VTAIL.n99 8.92171
R1312 VTAIL.n136 VTAIL.n112 8.92171
R1313 VTAIL.n152 VTAIL.n151 8.92171
R1314 VTAIL.n360 VTAIL.n359 8.92171
R1315 VTAIL.n344 VTAIL.n320 8.92171
R1316 VTAIL.n308 VTAIL.n307 8.92171
R1317 VTAIL.n292 VTAIL.n268 8.92171
R1318 VTAIL.n256 VTAIL.n255 8.92171
R1319 VTAIL.n240 VTAIL.n216 8.92171
R1320 VTAIL.n204 VTAIL.n203 8.92171
R1321 VTAIL.n188 VTAIL.n164 8.92171
R1322 VTAIL.n400 VTAIL.n399 8.14595
R1323 VTAIL.n408 VTAIL.n366 8.14595
R1324 VTAIL.n36 VTAIL.n35 8.14595
R1325 VTAIL.n44 VTAIL.n2 8.14595
R1326 VTAIL.n88 VTAIL.n87 8.14595
R1327 VTAIL.n96 VTAIL.n54 8.14595
R1328 VTAIL.n140 VTAIL.n139 8.14595
R1329 VTAIL.n148 VTAIL.n106 8.14595
R1330 VTAIL.n356 VTAIL.n314 8.14595
R1331 VTAIL.n348 VTAIL.n347 8.14595
R1332 VTAIL.n304 VTAIL.n262 8.14595
R1333 VTAIL.n296 VTAIL.n295 8.14595
R1334 VTAIL.n252 VTAIL.n210 8.14595
R1335 VTAIL.n244 VTAIL.n243 8.14595
R1336 VTAIL.n200 VTAIL.n158 8.14595
R1337 VTAIL.n192 VTAIL.n191 8.14595
R1338 VTAIL.n403 VTAIL.n370 7.3702
R1339 VTAIL.n407 VTAIL.n368 7.3702
R1340 VTAIL.n39 VTAIL.n6 7.3702
R1341 VTAIL.n43 VTAIL.n4 7.3702
R1342 VTAIL.n91 VTAIL.n58 7.3702
R1343 VTAIL.n95 VTAIL.n56 7.3702
R1344 VTAIL.n143 VTAIL.n110 7.3702
R1345 VTAIL.n147 VTAIL.n108 7.3702
R1346 VTAIL.n355 VTAIL.n316 7.3702
R1347 VTAIL.n351 VTAIL.n318 7.3702
R1348 VTAIL.n303 VTAIL.n264 7.3702
R1349 VTAIL.n299 VTAIL.n266 7.3702
R1350 VTAIL.n251 VTAIL.n212 7.3702
R1351 VTAIL.n247 VTAIL.n214 7.3702
R1352 VTAIL.n199 VTAIL.n160 7.3702
R1353 VTAIL.n195 VTAIL.n162 7.3702
R1354 VTAIL.n404 VTAIL.n403 6.59444
R1355 VTAIL.n404 VTAIL.n368 6.59444
R1356 VTAIL.n40 VTAIL.n39 6.59444
R1357 VTAIL.n40 VTAIL.n4 6.59444
R1358 VTAIL.n92 VTAIL.n91 6.59444
R1359 VTAIL.n92 VTAIL.n56 6.59444
R1360 VTAIL.n144 VTAIL.n143 6.59444
R1361 VTAIL.n144 VTAIL.n108 6.59444
R1362 VTAIL.n352 VTAIL.n316 6.59444
R1363 VTAIL.n352 VTAIL.n351 6.59444
R1364 VTAIL.n300 VTAIL.n264 6.59444
R1365 VTAIL.n300 VTAIL.n299 6.59444
R1366 VTAIL.n248 VTAIL.n212 6.59444
R1367 VTAIL.n248 VTAIL.n247 6.59444
R1368 VTAIL.n196 VTAIL.n160 6.59444
R1369 VTAIL.n196 VTAIL.n195 6.59444
R1370 VTAIL.n400 VTAIL.n370 5.81868
R1371 VTAIL.n408 VTAIL.n407 5.81868
R1372 VTAIL.n36 VTAIL.n6 5.81868
R1373 VTAIL.n44 VTAIL.n43 5.81868
R1374 VTAIL.n88 VTAIL.n58 5.81868
R1375 VTAIL.n96 VTAIL.n95 5.81868
R1376 VTAIL.n140 VTAIL.n110 5.81868
R1377 VTAIL.n148 VTAIL.n147 5.81868
R1378 VTAIL.n356 VTAIL.n355 5.81868
R1379 VTAIL.n348 VTAIL.n318 5.81868
R1380 VTAIL.n304 VTAIL.n303 5.81868
R1381 VTAIL.n296 VTAIL.n266 5.81868
R1382 VTAIL.n252 VTAIL.n251 5.81868
R1383 VTAIL.n244 VTAIL.n214 5.81868
R1384 VTAIL.n200 VTAIL.n199 5.81868
R1385 VTAIL.n192 VTAIL.n162 5.81868
R1386 VTAIL.n399 VTAIL.n372 5.04292
R1387 VTAIL.n411 VTAIL.n366 5.04292
R1388 VTAIL.n35 VTAIL.n8 5.04292
R1389 VTAIL.n47 VTAIL.n2 5.04292
R1390 VTAIL.n87 VTAIL.n60 5.04292
R1391 VTAIL.n99 VTAIL.n54 5.04292
R1392 VTAIL.n139 VTAIL.n112 5.04292
R1393 VTAIL.n151 VTAIL.n106 5.04292
R1394 VTAIL.n359 VTAIL.n314 5.04292
R1395 VTAIL.n347 VTAIL.n320 5.04292
R1396 VTAIL.n307 VTAIL.n262 5.04292
R1397 VTAIL.n295 VTAIL.n268 5.04292
R1398 VTAIL.n255 VTAIL.n210 5.04292
R1399 VTAIL.n243 VTAIL.n216 5.04292
R1400 VTAIL.n203 VTAIL.n158 5.04292
R1401 VTAIL.n191 VTAIL.n164 5.04292
R1402 VTAIL.n396 VTAIL.n395 4.26717
R1403 VTAIL.n412 VTAIL.n364 4.26717
R1404 VTAIL.n32 VTAIL.n31 4.26717
R1405 VTAIL.n48 VTAIL.n0 4.26717
R1406 VTAIL.n84 VTAIL.n83 4.26717
R1407 VTAIL.n100 VTAIL.n52 4.26717
R1408 VTAIL.n136 VTAIL.n135 4.26717
R1409 VTAIL.n152 VTAIL.n104 4.26717
R1410 VTAIL.n360 VTAIL.n312 4.26717
R1411 VTAIL.n344 VTAIL.n343 4.26717
R1412 VTAIL.n308 VTAIL.n260 4.26717
R1413 VTAIL.n292 VTAIL.n291 4.26717
R1414 VTAIL.n256 VTAIL.n208 4.26717
R1415 VTAIL.n240 VTAIL.n239 4.26717
R1416 VTAIL.n204 VTAIL.n156 4.26717
R1417 VTAIL.n188 VTAIL.n187 4.26717
R1418 VTAIL.n382 VTAIL.n381 3.70984
R1419 VTAIL.n18 VTAIL.n17 3.70984
R1420 VTAIL.n70 VTAIL.n69 3.70984
R1421 VTAIL.n122 VTAIL.n121 3.70984
R1422 VTAIL.n278 VTAIL.n277 3.70984
R1423 VTAIL.n226 VTAIL.n225 3.70984
R1424 VTAIL.n174 VTAIL.n173 3.70984
R1425 VTAIL.n330 VTAIL.n329 3.70984
R1426 VTAIL.n392 VTAIL.n374 3.49141
R1427 VTAIL.n28 VTAIL.n10 3.49141
R1428 VTAIL.n80 VTAIL.n62 3.49141
R1429 VTAIL.n132 VTAIL.n114 3.49141
R1430 VTAIL.n340 VTAIL.n322 3.49141
R1431 VTAIL.n288 VTAIL.n270 3.49141
R1432 VTAIL.n236 VTAIL.n218 3.49141
R1433 VTAIL.n184 VTAIL.n166 3.49141
R1434 VTAIL.n391 VTAIL.n376 2.71565
R1435 VTAIL.n27 VTAIL.n12 2.71565
R1436 VTAIL.n79 VTAIL.n64 2.71565
R1437 VTAIL.n131 VTAIL.n116 2.71565
R1438 VTAIL.n339 VTAIL.n324 2.71565
R1439 VTAIL.n287 VTAIL.n272 2.71565
R1440 VTAIL.n235 VTAIL.n220 2.71565
R1441 VTAIL.n183 VTAIL.n168 2.71565
R1442 VTAIL.n259 VTAIL.n207 2.65567
R1443 VTAIL.n363 VTAIL.n311 2.65567
R1444 VTAIL.n155 VTAIL.n103 2.65567
R1445 VTAIL.n388 VTAIL.n387 1.93989
R1446 VTAIL.n24 VTAIL.n23 1.93989
R1447 VTAIL.n76 VTAIL.n75 1.93989
R1448 VTAIL.n128 VTAIL.n127 1.93989
R1449 VTAIL.n336 VTAIL.n335 1.93989
R1450 VTAIL.n284 VTAIL.n283 1.93989
R1451 VTAIL.n232 VTAIL.n231 1.93989
R1452 VTAIL.n180 VTAIL.n179 1.93989
R1453 VTAIL VTAIL.n51 1.38628
R1454 VTAIL VTAIL.n415 1.2699
R1455 VTAIL.n384 VTAIL.n378 1.16414
R1456 VTAIL.n20 VTAIL.n14 1.16414
R1457 VTAIL.n72 VTAIL.n66 1.16414
R1458 VTAIL.n124 VTAIL.n118 1.16414
R1459 VTAIL.n332 VTAIL.n326 1.16414
R1460 VTAIL.n280 VTAIL.n274 1.16414
R1461 VTAIL.n228 VTAIL.n222 1.16414
R1462 VTAIL.n176 VTAIL.n170 1.16414
R1463 VTAIL.n311 VTAIL.n259 0.470328
R1464 VTAIL.n103 VTAIL.n51 0.470328
R1465 VTAIL.n383 VTAIL.n380 0.388379
R1466 VTAIL.n19 VTAIL.n16 0.388379
R1467 VTAIL.n71 VTAIL.n68 0.388379
R1468 VTAIL.n123 VTAIL.n120 0.388379
R1469 VTAIL.n331 VTAIL.n328 0.388379
R1470 VTAIL.n279 VTAIL.n276 0.388379
R1471 VTAIL.n227 VTAIL.n224 0.388379
R1472 VTAIL.n175 VTAIL.n172 0.388379
R1473 VTAIL.n382 VTAIL.n377 0.155672
R1474 VTAIL.n389 VTAIL.n377 0.155672
R1475 VTAIL.n390 VTAIL.n389 0.155672
R1476 VTAIL.n390 VTAIL.n373 0.155672
R1477 VTAIL.n397 VTAIL.n373 0.155672
R1478 VTAIL.n398 VTAIL.n397 0.155672
R1479 VTAIL.n398 VTAIL.n369 0.155672
R1480 VTAIL.n405 VTAIL.n369 0.155672
R1481 VTAIL.n406 VTAIL.n405 0.155672
R1482 VTAIL.n406 VTAIL.n365 0.155672
R1483 VTAIL.n413 VTAIL.n365 0.155672
R1484 VTAIL.n18 VTAIL.n13 0.155672
R1485 VTAIL.n25 VTAIL.n13 0.155672
R1486 VTAIL.n26 VTAIL.n25 0.155672
R1487 VTAIL.n26 VTAIL.n9 0.155672
R1488 VTAIL.n33 VTAIL.n9 0.155672
R1489 VTAIL.n34 VTAIL.n33 0.155672
R1490 VTAIL.n34 VTAIL.n5 0.155672
R1491 VTAIL.n41 VTAIL.n5 0.155672
R1492 VTAIL.n42 VTAIL.n41 0.155672
R1493 VTAIL.n42 VTAIL.n1 0.155672
R1494 VTAIL.n49 VTAIL.n1 0.155672
R1495 VTAIL.n70 VTAIL.n65 0.155672
R1496 VTAIL.n77 VTAIL.n65 0.155672
R1497 VTAIL.n78 VTAIL.n77 0.155672
R1498 VTAIL.n78 VTAIL.n61 0.155672
R1499 VTAIL.n85 VTAIL.n61 0.155672
R1500 VTAIL.n86 VTAIL.n85 0.155672
R1501 VTAIL.n86 VTAIL.n57 0.155672
R1502 VTAIL.n93 VTAIL.n57 0.155672
R1503 VTAIL.n94 VTAIL.n93 0.155672
R1504 VTAIL.n94 VTAIL.n53 0.155672
R1505 VTAIL.n101 VTAIL.n53 0.155672
R1506 VTAIL.n122 VTAIL.n117 0.155672
R1507 VTAIL.n129 VTAIL.n117 0.155672
R1508 VTAIL.n130 VTAIL.n129 0.155672
R1509 VTAIL.n130 VTAIL.n113 0.155672
R1510 VTAIL.n137 VTAIL.n113 0.155672
R1511 VTAIL.n138 VTAIL.n137 0.155672
R1512 VTAIL.n138 VTAIL.n109 0.155672
R1513 VTAIL.n145 VTAIL.n109 0.155672
R1514 VTAIL.n146 VTAIL.n145 0.155672
R1515 VTAIL.n146 VTAIL.n105 0.155672
R1516 VTAIL.n153 VTAIL.n105 0.155672
R1517 VTAIL.n361 VTAIL.n313 0.155672
R1518 VTAIL.n354 VTAIL.n313 0.155672
R1519 VTAIL.n354 VTAIL.n353 0.155672
R1520 VTAIL.n353 VTAIL.n317 0.155672
R1521 VTAIL.n346 VTAIL.n317 0.155672
R1522 VTAIL.n346 VTAIL.n345 0.155672
R1523 VTAIL.n345 VTAIL.n321 0.155672
R1524 VTAIL.n338 VTAIL.n321 0.155672
R1525 VTAIL.n338 VTAIL.n337 0.155672
R1526 VTAIL.n337 VTAIL.n325 0.155672
R1527 VTAIL.n330 VTAIL.n325 0.155672
R1528 VTAIL.n309 VTAIL.n261 0.155672
R1529 VTAIL.n302 VTAIL.n261 0.155672
R1530 VTAIL.n302 VTAIL.n301 0.155672
R1531 VTAIL.n301 VTAIL.n265 0.155672
R1532 VTAIL.n294 VTAIL.n265 0.155672
R1533 VTAIL.n294 VTAIL.n293 0.155672
R1534 VTAIL.n293 VTAIL.n269 0.155672
R1535 VTAIL.n286 VTAIL.n269 0.155672
R1536 VTAIL.n286 VTAIL.n285 0.155672
R1537 VTAIL.n285 VTAIL.n273 0.155672
R1538 VTAIL.n278 VTAIL.n273 0.155672
R1539 VTAIL.n257 VTAIL.n209 0.155672
R1540 VTAIL.n250 VTAIL.n209 0.155672
R1541 VTAIL.n250 VTAIL.n249 0.155672
R1542 VTAIL.n249 VTAIL.n213 0.155672
R1543 VTAIL.n242 VTAIL.n213 0.155672
R1544 VTAIL.n242 VTAIL.n241 0.155672
R1545 VTAIL.n241 VTAIL.n217 0.155672
R1546 VTAIL.n234 VTAIL.n217 0.155672
R1547 VTAIL.n234 VTAIL.n233 0.155672
R1548 VTAIL.n233 VTAIL.n221 0.155672
R1549 VTAIL.n226 VTAIL.n221 0.155672
R1550 VTAIL.n205 VTAIL.n157 0.155672
R1551 VTAIL.n198 VTAIL.n157 0.155672
R1552 VTAIL.n198 VTAIL.n197 0.155672
R1553 VTAIL.n197 VTAIL.n161 0.155672
R1554 VTAIL.n190 VTAIL.n161 0.155672
R1555 VTAIL.n190 VTAIL.n189 0.155672
R1556 VTAIL.n189 VTAIL.n165 0.155672
R1557 VTAIL.n182 VTAIL.n165 0.155672
R1558 VTAIL.n182 VTAIL.n181 0.155672
R1559 VTAIL.n181 VTAIL.n169 0.155672
R1560 VTAIL.n174 VTAIL.n169 0.155672
R1561 VDD2.n2 VDD2.n0 117.094
R1562 VDD2.n2 VDD2.n1 77.2163
R1563 VDD2.n1 VDD2.t1 3.41848
R1564 VDD2.n1 VDD2.t2 3.41848
R1565 VDD2.n0 VDD2.t0 3.41848
R1566 VDD2.n0 VDD2.t3 3.41848
R1567 VDD2 VDD2.n2 0.0586897
R1568 VP.n16 VP.n0 161.3
R1569 VP.n15 VP.n14 161.3
R1570 VP.n13 VP.n1 161.3
R1571 VP.n12 VP.n11 161.3
R1572 VP.n10 VP.n2 161.3
R1573 VP.n9 VP.n8 161.3
R1574 VP.n7 VP.n3 161.3
R1575 VP.n4 VP.t1 117.838
R1576 VP.n4 VP.t2 116.959
R1577 VP.n6 VP.n5 108.799
R1578 VP.n18 VP.n17 108.799
R1579 VP.n5 VP.t0 83.3427
R1580 VP.n17 VP.t3 83.3427
R1581 VP.n6 VP.n4 48.4035
R1582 VP.n11 VP.n10 40.4934
R1583 VP.n11 VP.n1 40.4934
R1584 VP.n9 VP.n3 24.4675
R1585 VP.n10 VP.n9 24.4675
R1586 VP.n15 VP.n1 24.4675
R1587 VP.n16 VP.n15 24.4675
R1588 VP.n5 VP.n3 1.95786
R1589 VP.n17 VP.n16 1.95786
R1590 VP.n7 VP.n6 0.278367
R1591 VP.n18 VP.n0 0.278367
R1592 VP.n8 VP.n7 0.189894
R1593 VP.n8 VP.n2 0.189894
R1594 VP.n12 VP.n2 0.189894
R1595 VP.n13 VP.n12 0.189894
R1596 VP.n14 VP.n13 0.189894
R1597 VP.n14 VP.n0 0.189894
R1598 VP VP.n18 0.153454
R1599 VDD1 VDD1.n1 117.62
R1600 VDD1 VDD1.n0 77.2745
R1601 VDD1.n0 VDD1.t2 3.41848
R1602 VDD1.n0 VDD1.t1 3.41848
R1603 VDD1.n1 VDD1.t3 3.41848
R1604 VDD1.n1 VDD1.t0 3.41848
C0 w_n2818_n2870# VDD1 1.41256f
C1 B VDD1 1.2204f
C2 VP w_n2818_n2870# 5.12268f
C3 VP B 1.71041f
C4 VDD2 VDD1 1.05686f
C5 VP VDD2 0.403687f
C6 VP VDD1 4.12531f
C7 VN VTAIL 3.90924f
C8 VTAIL w_n2818_n2870# 3.42204f
C9 VTAIL B 4.18887f
C10 VN w_n2818_n2870# 4.76004f
C11 VN B 1.10792f
C12 w_n2818_n2870# B 8.732519f
C13 VTAIL VDD2 4.90954f
C14 VTAIL VDD1 4.85433f
C15 VP VTAIL 3.92334f
C16 VN VDD2 3.87137f
C17 VN VDD1 0.148973f
C18 w_n2818_n2870# VDD2 1.472f
C19 VDD2 B 1.27503f
C20 VP VN 5.83965f
C21 VDD2 VSUBS 0.917969f
C22 VDD1 VSUBS 5.544271f
C23 VTAIL VSUBS 1.11781f
C24 VN VSUBS 5.47188f
C25 VP VSUBS 2.264085f
C26 B VSUBS 4.195889f
C27 w_n2818_n2870# VSUBS 0.099994p
C28 VDD1.t2 VSUBS 0.206758f
C29 VDD1.t1 VSUBS 0.206758f
C30 VDD1.n0 VSUBS 1.52732f
C31 VDD1.t3 VSUBS 0.206758f
C32 VDD1.t0 VSUBS 0.206758f
C33 VDD1.n1 VSUBS 2.17741f
C34 VP.n0 VSUBS 0.046551f
C35 VP.t3 VSUBS 2.49715f
C36 VP.n1 VSUBS 0.070177f
C37 VP.n2 VSUBS 0.035309f
C38 VP.n3 VSUBS 0.035917f
C39 VP.t2 VSUBS 2.82124f
C40 VP.t1 VSUBS 2.8295f
C41 VP.n4 VSUBS 3.64211f
C42 VP.t0 VSUBS 2.49715f
C43 VP.n5 VSUBS 1.00532f
C44 VP.n6 VSUBS 1.8534f
C45 VP.n7 VSUBS 0.046551f
C46 VP.n8 VSUBS 0.035309f
C47 VP.n9 VSUBS 0.065807f
C48 VP.n10 VSUBS 0.070177f
C49 VP.n11 VSUBS 0.028544f
C50 VP.n12 VSUBS 0.035309f
C51 VP.n13 VSUBS 0.035309f
C52 VP.n14 VSUBS 0.035309f
C53 VP.n15 VSUBS 0.065807f
C54 VP.n16 VSUBS 0.035917f
C55 VP.n17 VSUBS 1.00532f
C56 VP.n18 VSUBS 0.065808f
C57 VDD2.t0 VSUBS 0.204472f
C58 VDD2.t3 VSUBS 0.204472f
C59 VDD2.n0 VSUBS 2.12932f
C60 VDD2.t1 VSUBS 0.204472f
C61 VDD2.t2 VSUBS 0.204472f
C62 VDD2.n1 VSUBS 1.50987f
C63 VDD2.n2 VSUBS 4.10428f
C64 VTAIL.n0 VSUBS 0.028356f
C65 VTAIL.n1 VSUBS 0.024846f
C66 VTAIL.n2 VSUBS 0.013351f
C67 VTAIL.n3 VSUBS 0.031558f
C68 VTAIL.n4 VSUBS 0.014137f
C69 VTAIL.n5 VSUBS 0.024846f
C70 VTAIL.n6 VSUBS 0.013351f
C71 VTAIL.n7 VSUBS 0.031558f
C72 VTAIL.n8 VSUBS 0.014137f
C73 VTAIL.n9 VSUBS 0.024846f
C74 VTAIL.n10 VSUBS 0.013351f
C75 VTAIL.n11 VSUBS 0.031558f
C76 VTAIL.n12 VSUBS 0.014137f
C77 VTAIL.n13 VSUBS 0.024846f
C78 VTAIL.n14 VSUBS 0.013351f
C79 VTAIL.n15 VSUBS 0.023668f
C80 VTAIL.n16 VSUBS 0.020076f
C81 VTAIL.t4 VSUBS 0.067281f
C82 VTAIL.n17 VSUBS 0.134973f
C83 VTAIL.n18 VSUBS 0.967122f
C84 VTAIL.n19 VSUBS 0.013351f
C85 VTAIL.n20 VSUBS 0.014137f
C86 VTAIL.n21 VSUBS 0.031558f
C87 VTAIL.n22 VSUBS 0.031558f
C88 VTAIL.n23 VSUBS 0.014137f
C89 VTAIL.n24 VSUBS 0.013351f
C90 VTAIL.n25 VSUBS 0.024846f
C91 VTAIL.n26 VSUBS 0.024846f
C92 VTAIL.n27 VSUBS 0.013351f
C93 VTAIL.n28 VSUBS 0.014137f
C94 VTAIL.n29 VSUBS 0.031558f
C95 VTAIL.n30 VSUBS 0.031558f
C96 VTAIL.n31 VSUBS 0.014137f
C97 VTAIL.n32 VSUBS 0.013351f
C98 VTAIL.n33 VSUBS 0.024846f
C99 VTAIL.n34 VSUBS 0.024846f
C100 VTAIL.n35 VSUBS 0.013351f
C101 VTAIL.n36 VSUBS 0.014137f
C102 VTAIL.n37 VSUBS 0.031558f
C103 VTAIL.n38 VSUBS 0.031558f
C104 VTAIL.n39 VSUBS 0.014137f
C105 VTAIL.n40 VSUBS 0.013351f
C106 VTAIL.n41 VSUBS 0.024846f
C107 VTAIL.n42 VSUBS 0.024846f
C108 VTAIL.n43 VSUBS 0.013351f
C109 VTAIL.n44 VSUBS 0.014137f
C110 VTAIL.n45 VSUBS 0.031558f
C111 VTAIL.n46 VSUBS 0.079991f
C112 VTAIL.n47 VSUBS 0.014137f
C113 VTAIL.n48 VSUBS 0.013351f
C114 VTAIL.n49 VSUBS 0.054376f
C115 VTAIL.n50 VSUBS 0.04029f
C116 VTAIL.n51 VSUBS 0.16806f
C117 VTAIL.n52 VSUBS 0.028356f
C118 VTAIL.n53 VSUBS 0.024846f
C119 VTAIL.n54 VSUBS 0.013351f
C120 VTAIL.n55 VSUBS 0.031558f
C121 VTAIL.n56 VSUBS 0.014137f
C122 VTAIL.n57 VSUBS 0.024846f
C123 VTAIL.n58 VSUBS 0.013351f
C124 VTAIL.n59 VSUBS 0.031558f
C125 VTAIL.n60 VSUBS 0.014137f
C126 VTAIL.n61 VSUBS 0.024846f
C127 VTAIL.n62 VSUBS 0.013351f
C128 VTAIL.n63 VSUBS 0.031558f
C129 VTAIL.n64 VSUBS 0.014137f
C130 VTAIL.n65 VSUBS 0.024846f
C131 VTAIL.n66 VSUBS 0.013351f
C132 VTAIL.n67 VSUBS 0.023668f
C133 VTAIL.n68 VSUBS 0.020076f
C134 VTAIL.t3 VSUBS 0.067281f
C135 VTAIL.n69 VSUBS 0.134973f
C136 VTAIL.n70 VSUBS 0.967122f
C137 VTAIL.n71 VSUBS 0.013351f
C138 VTAIL.n72 VSUBS 0.014137f
C139 VTAIL.n73 VSUBS 0.031558f
C140 VTAIL.n74 VSUBS 0.031558f
C141 VTAIL.n75 VSUBS 0.014137f
C142 VTAIL.n76 VSUBS 0.013351f
C143 VTAIL.n77 VSUBS 0.024846f
C144 VTAIL.n78 VSUBS 0.024846f
C145 VTAIL.n79 VSUBS 0.013351f
C146 VTAIL.n80 VSUBS 0.014137f
C147 VTAIL.n81 VSUBS 0.031558f
C148 VTAIL.n82 VSUBS 0.031558f
C149 VTAIL.n83 VSUBS 0.014137f
C150 VTAIL.n84 VSUBS 0.013351f
C151 VTAIL.n85 VSUBS 0.024846f
C152 VTAIL.n86 VSUBS 0.024846f
C153 VTAIL.n87 VSUBS 0.013351f
C154 VTAIL.n88 VSUBS 0.014137f
C155 VTAIL.n89 VSUBS 0.031558f
C156 VTAIL.n90 VSUBS 0.031558f
C157 VTAIL.n91 VSUBS 0.014137f
C158 VTAIL.n92 VSUBS 0.013351f
C159 VTAIL.n93 VSUBS 0.024846f
C160 VTAIL.n94 VSUBS 0.024846f
C161 VTAIL.n95 VSUBS 0.013351f
C162 VTAIL.n96 VSUBS 0.014137f
C163 VTAIL.n97 VSUBS 0.031558f
C164 VTAIL.n98 VSUBS 0.079991f
C165 VTAIL.n99 VSUBS 0.014137f
C166 VTAIL.n100 VSUBS 0.013351f
C167 VTAIL.n101 VSUBS 0.054376f
C168 VTAIL.n102 VSUBS 0.04029f
C169 VTAIL.n103 VSUBS 0.269689f
C170 VTAIL.n104 VSUBS 0.028356f
C171 VTAIL.n105 VSUBS 0.024846f
C172 VTAIL.n106 VSUBS 0.013351f
C173 VTAIL.n107 VSUBS 0.031558f
C174 VTAIL.n108 VSUBS 0.014137f
C175 VTAIL.n109 VSUBS 0.024846f
C176 VTAIL.n110 VSUBS 0.013351f
C177 VTAIL.n111 VSUBS 0.031558f
C178 VTAIL.n112 VSUBS 0.014137f
C179 VTAIL.n113 VSUBS 0.024846f
C180 VTAIL.n114 VSUBS 0.013351f
C181 VTAIL.n115 VSUBS 0.031558f
C182 VTAIL.n116 VSUBS 0.014137f
C183 VTAIL.n117 VSUBS 0.024846f
C184 VTAIL.n118 VSUBS 0.013351f
C185 VTAIL.n119 VSUBS 0.023668f
C186 VTAIL.n120 VSUBS 0.020076f
C187 VTAIL.t0 VSUBS 0.067281f
C188 VTAIL.n121 VSUBS 0.134973f
C189 VTAIL.n122 VSUBS 0.967122f
C190 VTAIL.n123 VSUBS 0.013351f
C191 VTAIL.n124 VSUBS 0.014137f
C192 VTAIL.n125 VSUBS 0.031558f
C193 VTAIL.n126 VSUBS 0.031558f
C194 VTAIL.n127 VSUBS 0.014137f
C195 VTAIL.n128 VSUBS 0.013351f
C196 VTAIL.n129 VSUBS 0.024846f
C197 VTAIL.n130 VSUBS 0.024846f
C198 VTAIL.n131 VSUBS 0.013351f
C199 VTAIL.n132 VSUBS 0.014137f
C200 VTAIL.n133 VSUBS 0.031558f
C201 VTAIL.n134 VSUBS 0.031558f
C202 VTAIL.n135 VSUBS 0.014137f
C203 VTAIL.n136 VSUBS 0.013351f
C204 VTAIL.n137 VSUBS 0.024846f
C205 VTAIL.n138 VSUBS 0.024846f
C206 VTAIL.n139 VSUBS 0.013351f
C207 VTAIL.n140 VSUBS 0.014137f
C208 VTAIL.n141 VSUBS 0.031558f
C209 VTAIL.n142 VSUBS 0.031558f
C210 VTAIL.n143 VSUBS 0.014137f
C211 VTAIL.n144 VSUBS 0.013351f
C212 VTAIL.n145 VSUBS 0.024846f
C213 VTAIL.n146 VSUBS 0.024846f
C214 VTAIL.n147 VSUBS 0.013351f
C215 VTAIL.n148 VSUBS 0.014137f
C216 VTAIL.n149 VSUBS 0.031558f
C217 VTAIL.n150 VSUBS 0.079991f
C218 VTAIL.n151 VSUBS 0.014137f
C219 VTAIL.n152 VSUBS 0.013351f
C220 VTAIL.n153 VSUBS 0.054376f
C221 VTAIL.n154 VSUBS 0.04029f
C222 VTAIL.n155 VSUBS 1.43852f
C223 VTAIL.n156 VSUBS 0.028356f
C224 VTAIL.n157 VSUBS 0.024846f
C225 VTAIL.n158 VSUBS 0.013351f
C226 VTAIL.n159 VSUBS 0.031558f
C227 VTAIL.n160 VSUBS 0.014137f
C228 VTAIL.n161 VSUBS 0.024846f
C229 VTAIL.n162 VSUBS 0.013351f
C230 VTAIL.n163 VSUBS 0.031558f
C231 VTAIL.n164 VSUBS 0.014137f
C232 VTAIL.n165 VSUBS 0.024846f
C233 VTAIL.n166 VSUBS 0.013351f
C234 VTAIL.n167 VSUBS 0.031558f
C235 VTAIL.n168 VSUBS 0.014137f
C236 VTAIL.n169 VSUBS 0.024846f
C237 VTAIL.n170 VSUBS 0.013351f
C238 VTAIL.n171 VSUBS 0.023668f
C239 VTAIL.n172 VSUBS 0.020076f
C240 VTAIL.t6 VSUBS 0.067281f
C241 VTAIL.n173 VSUBS 0.134973f
C242 VTAIL.n174 VSUBS 0.967121f
C243 VTAIL.n175 VSUBS 0.013351f
C244 VTAIL.n176 VSUBS 0.014137f
C245 VTAIL.n177 VSUBS 0.031558f
C246 VTAIL.n178 VSUBS 0.031558f
C247 VTAIL.n179 VSUBS 0.014137f
C248 VTAIL.n180 VSUBS 0.013351f
C249 VTAIL.n181 VSUBS 0.024846f
C250 VTAIL.n182 VSUBS 0.024846f
C251 VTAIL.n183 VSUBS 0.013351f
C252 VTAIL.n184 VSUBS 0.014137f
C253 VTAIL.n185 VSUBS 0.031558f
C254 VTAIL.n186 VSUBS 0.031558f
C255 VTAIL.n187 VSUBS 0.014137f
C256 VTAIL.n188 VSUBS 0.013351f
C257 VTAIL.n189 VSUBS 0.024846f
C258 VTAIL.n190 VSUBS 0.024846f
C259 VTAIL.n191 VSUBS 0.013351f
C260 VTAIL.n192 VSUBS 0.014137f
C261 VTAIL.n193 VSUBS 0.031558f
C262 VTAIL.n194 VSUBS 0.031558f
C263 VTAIL.n195 VSUBS 0.014137f
C264 VTAIL.n196 VSUBS 0.013351f
C265 VTAIL.n197 VSUBS 0.024846f
C266 VTAIL.n198 VSUBS 0.024846f
C267 VTAIL.n199 VSUBS 0.013351f
C268 VTAIL.n200 VSUBS 0.014137f
C269 VTAIL.n201 VSUBS 0.031558f
C270 VTAIL.n202 VSUBS 0.079991f
C271 VTAIL.n203 VSUBS 0.014137f
C272 VTAIL.n204 VSUBS 0.013351f
C273 VTAIL.n205 VSUBS 0.054376f
C274 VTAIL.n206 VSUBS 0.04029f
C275 VTAIL.n207 VSUBS 1.43852f
C276 VTAIL.n208 VSUBS 0.028356f
C277 VTAIL.n209 VSUBS 0.024846f
C278 VTAIL.n210 VSUBS 0.013351f
C279 VTAIL.n211 VSUBS 0.031558f
C280 VTAIL.n212 VSUBS 0.014137f
C281 VTAIL.n213 VSUBS 0.024846f
C282 VTAIL.n214 VSUBS 0.013351f
C283 VTAIL.n215 VSUBS 0.031558f
C284 VTAIL.n216 VSUBS 0.014137f
C285 VTAIL.n217 VSUBS 0.024846f
C286 VTAIL.n218 VSUBS 0.013351f
C287 VTAIL.n219 VSUBS 0.031558f
C288 VTAIL.n220 VSUBS 0.014137f
C289 VTAIL.n221 VSUBS 0.024846f
C290 VTAIL.n222 VSUBS 0.013351f
C291 VTAIL.n223 VSUBS 0.023668f
C292 VTAIL.n224 VSUBS 0.020076f
C293 VTAIL.t7 VSUBS 0.067281f
C294 VTAIL.n225 VSUBS 0.134973f
C295 VTAIL.n226 VSUBS 0.967121f
C296 VTAIL.n227 VSUBS 0.013351f
C297 VTAIL.n228 VSUBS 0.014137f
C298 VTAIL.n229 VSUBS 0.031558f
C299 VTAIL.n230 VSUBS 0.031558f
C300 VTAIL.n231 VSUBS 0.014137f
C301 VTAIL.n232 VSUBS 0.013351f
C302 VTAIL.n233 VSUBS 0.024846f
C303 VTAIL.n234 VSUBS 0.024846f
C304 VTAIL.n235 VSUBS 0.013351f
C305 VTAIL.n236 VSUBS 0.014137f
C306 VTAIL.n237 VSUBS 0.031558f
C307 VTAIL.n238 VSUBS 0.031558f
C308 VTAIL.n239 VSUBS 0.014137f
C309 VTAIL.n240 VSUBS 0.013351f
C310 VTAIL.n241 VSUBS 0.024846f
C311 VTAIL.n242 VSUBS 0.024846f
C312 VTAIL.n243 VSUBS 0.013351f
C313 VTAIL.n244 VSUBS 0.014137f
C314 VTAIL.n245 VSUBS 0.031558f
C315 VTAIL.n246 VSUBS 0.031558f
C316 VTAIL.n247 VSUBS 0.014137f
C317 VTAIL.n248 VSUBS 0.013351f
C318 VTAIL.n249 VSUBS 0.024846f
C319 VTAIL.n250 VSUBS 0.024846f
C320 VTAIL.n251 VSUBS 0.013351f
C321 VTAIL.n252 VSUBS 0.014137f
C322 VTAIL.n253 VSUBS 0.031558f
C323 VTAIL.n254 VSUBS 0.079991f
C324 VTAIL.n255 VSUBS 0.014137f
C325 VTAIL.n256 VSUBS 0.013351f
C326 VTAIL.n257 VSUBS 0.054376f
C327 VTAIL.n258 VSUBS 0.04029f
C328 VTAIL.n259 VSUBS 0.269689f
C329 VTAIL.n260 VSUBS 0.028356f
C330 VTAIL.n261 VSUBS 0.024846f
C331 VTAIL.n262 VSUBS 0.013351f
C332 VTAIL.n263 VSUBS 0.031558f
C333 VTAIL.n264 VSUBS 0.014137f
C334 VTAIL.n265 VSUBS 0.024846f
C335 VTAIL.n266 VSUBS 0.013351f
C336 VTAIL.n267 VSUBS 0.031558f
C337 VTAIL.n268 VSUBS 0.014137f
C338 VTAIL.n269 VSUBS 0.024846f
C339 VTAIL.n270 VSUBS 0.013351f
C340 VTAIL.n271 VSUBS 0.031558f
C341 VTAIL.n272 VSUBS 0.014137f
C342 VTAIL.n273 VSUBS 0.024846f
C343 VTAIL.n274 VSUBS 0.013351f
C344 VTAIL.n275 VSUBS 0.023668f
C345 VTAIL.n276 VSUBS 0.020076f
C346 VTAIL.t2 VSUBS 0.067281f
C347 VTAIL.n277 VSUBS 0.134973f
C348 VTAIL.n278 VSUBS 0.967121f
C349 VTAIL.n279 VSUBS 0.013351f
C350 VTAIL.n280 VSUBS 0.014137f
C351 VTAIL.n281 VSUBS 0.031558f
C352 VTAIL.n282 VSUBS 0.031558f
C353 VTAIL.n283 VSUBS 0.014137f
C354 VTAIL.n284 VSUBS 0.013351f
C355 VTAIL.n285 VSUBS 0.024846f
C356 VTAIL.n286 VSUBS 0.024846f
C357 VTAIL.n287 VSUBS 0.013351f
C358 VTAIL.n288 VSUBS 0.014137f
C359 VTAIL.n289 VSUBS 0.031558f
C360 VTAIL.n290 VSUBS 0.031558f
C361 VTAIL.n291 VSUBS 0.014137f
C362 VTAIL.n292 VSUBS 0.013351f
C363 VTAIL.n293 VSUBS 0.024846f
C364 VTAIL.n294 VSUBS 0.024846f
C365 VTAIL.n295 VSUBS 0.013351f
C366 VTAIL.n296 VSUBS 0.014137f
C367 VTAIL.n297 VSUBS 0.031558f
C368 VTAIL.n298 VSUBS 0.031558f
C369 VTAIL.n299 VSUBS 0.014137f
C370 VTAIL.n300 VSUBS 0.013351f
C371 VTAIL.n301 VSUBS 0.024846f
C372 VTAIL.n302 VSUBS 0.024846f
C373 VTAIL.n303 VSUBS 0.013351f
C374 VTAIL.n304 VSUBS 0.014137f
C375 VTAIL.n305 VSUBS 0.031558f
C376 VTAIL.n306 VSUBS 0.079991f
C377 VTAIL.n307 VSUBS 0.014137f
C378 VTAIL.n308 VSUBS 0.013351f
C379 VTAIL.n309 VSUBS 0.054376f
C380 VTAIL.n310 VSUBS 0.04029f
C381 VTAIL.n311 VSUBS 0.269689f
C382 VTAIL.n312 VSUBS 0.028356f
C383 VTAIL.n313 VSUBS 0.024846f
C384 VTAIL.n314 VSUBS 0.013351f
C385 VTAIL.n315 VSUBS 0.031558f
C386 VTAIL.n316 VSUBS 0.014137f
C387 VTAIL.n317 VSUBS 0.024846f
C388 VTAIL.n318 VSUBS 0.013351f
C389 VTAIL.n319 VSUBS 0.031558f
C390 VTAIL.n320 VSUBS 0.014137f
C391 VTAIL.n321 VSUBS 0.024846f
C392 VTAIL.n322 VSUBS 0.013351f
C393 VTAIL.n323 VSUBS 0.031558f
C394 VTAIL.n324 VSUBS 0.014137f
C395 VTAIL.n325 VSUBS 0.024846f
C396 VTAIL.n326 VSUBS 0.013351f
C397 VTAIL.n327 VSUBS 0.023668f
C398 VTAIL.n328 VSUBS 0.020076f
C399 VTAIL.t1 VSUBS 0.067281f
C400 VTAIL.n329 VSUBS 0.134973f
C401 VTAIL.n330 VSUBS 0.967122f
C402 VTAIL.n331 VSUBS 0.013351f
C403 VTAIL.n332 VSUBS 0.014137f
C404 VTAIL.n333 VSUBS 0.031558f
C405 VTAIL.n334 VSUBS 0.031558f
C406 VTAIL.n335 VSUBS 0.014137f
C407 VTAIL.n336 VSUBS 0.013351f
C408 VTAIL.n337 VSUBS 0.024846f
C409 VTAIL.n338 VSUBS 0.024846f
C410 VTAIL.n339 VSUBS 0.013351f
C411 VTAIL.n340 VSUBS 0.014137f
C412 VTAIL.n341 VSUBS 0.031558f
C413 VTAIL.n342 VSUBS 0.031558f
C414 VTAIL.n343 VSUBS 0.014137f
C415 VTAIL.n344 VSUBS 0.013351f
C416 VTAIL.n345 VSUBS 0.024846f
C417 VTAIL.n346 VSUBS 0.024846f
C418 VTAIL.n347 VSUBS 0.013351f
C419 VTAIL.n348 VSUBS 0.014137f
C420 VTAIL.n349 VSUBS 0.031558f
C421 VTAIL.n350 VSUBS 0.031558f
C422 VTAIL.n351 VSUBS 0.014137f
C423 VTAIL.n352 VSUBS 0.013351f
C424 VTAIL.n353 VSUBS 0.024846f
C425 VTAIL.n354 VSUBS 0.024846f
C426 VTAIL.n355 VSUBS 0.013351f
C427 VTAIL.n356 VSUBS 0.014137f
C428 VTAIL.n357 VSUBS 0.031558f
C429 VTAIL.n358 VSUBS 0.079991f
C430 VTAIL.n359 VSUBS 0.014137f
C431 VTAIL.n360 VSUBS 0.013351f
C432 VTAIL.n361 VSUBS 0.054376f
C433 VTAIL.n362 VSUBS 0.04029f
C434 VTAIL.n363 VSUBS 1.43852f
C435 VTAIL.n364 VSUBS 0.028356f
C436 VTAIL.n365 VSUBS 0.024846f
C437 VTAIL.n366 VSUBS 0.013351f
C438 VTAIL.n367 VSUBS 0.031558f
C439 VTAIL.n368 VSUBS 0.014137f
C440 VTAIL.n369 VSUBS 0.024846f
C441 VTAIL.n370 VSUBS 0.013351f
C442 VTAIL.n371 VSUBS 0.031558f
C443 VTAIL.n372 VSUBS 0.014137f
C444 VTAIL.n373 VSUBS 0.024846f
C445 VTAIL.n374 VSUBS 0.013351f
C446 VTAIL.n375 VSUBS 0.031558f
C447 VTAIL.n376 VSUBS 0.014137f
C448 VTAIL.n377 VSUBS 0.024846f
C449 VTAIL.n378 VSUBS 0.013351f
C450 VTAIL.n379 VSUBS 0.023668f
C451 VTAIL.n380 VSUBS 0.020076f
C452 VTAIL.t5 VSUBS 0.067281f
C453 VTAIL.n381 VSUBS 0.134973f
C454 VTAIL.n382 VSUBS 0.967122f
C455 VTAIL.n383 VSUBS 0.013351f
C456 VTAIL.n384 VSUBS 0.014137f
C457 VTAIL.n385 VSUBS 0.031558f
C458 VTAIL.n386 VSUBS 0.031558f
C459 VTAIL.n387 VSUBS 0.014137f
C460 VTAIL.n388 VSUBS 0.013351f
C461 VTAIL.n389 VSUBS 0.024846f
C462 VTAIL.n390 VSUBS 0.024846f
C463 VTAIL.n391 VSUBS 0.013351f
C464 VTAIL.n392 VSUBS 0.014137f
C465 VTAIL.n393 VSUBS 0.031558f
C466 VTAIL.n394 VSUBS 0.031558f
C467 VTAIL.n395 VSUBS 0.014137f
C468 VTAIL.n396 VSUBS 0.013351f
C469 VTAIL.n397 VSUBS 0.024846f
C470 VTAIL.n398 VSUBS 0.024846f
C471 VTAIL.n399 VSUBS 0.013351f
C472 VTAIL.n400 VSUBS 0.014137f
C473 VTAIL.n401 VSUBS 0.031558f
C474 VTAIL.n402 VSUBS 0.031558f
C475 VTAIL.n403 VSUBS 0.014137f
C476 VTAIL.n404 VSUBS 0.013351f
C477 VTAIL.n405 VSUBS 0.024846f
C478 VTAIL.n406 VSUBS 0.024846f
C479 VTAIL.n407 VSUBS 0.013351f
C480 VTAIL.n408 VSUBS 0.014137f
C481 VTAIL.n409 VSUBS 0.031558f
C482 VTAIL.n410 VSUBS 0.079991f
C483 VTAIL.n411 VSUBS 0.014137f
C484 VTAIL.n412 VSUBS 0.013351f
C485 VTAIL.n413 VSUBS 0.054376f
C486 VTAIL.n414 VSUBS 0.04029f
C487 VTAIL.n415 VSUBS 1.32757f
C488 VN.t3 VSUBS 2.74743f
C489 VN.t0 VSUBS 2.73941f
C490 VN.n0 VSUBS 1.73023f
C491 VN.t1 VSUBS 2.74743f
C492 VN.t2 VSUBS 2.73941f
C493 VN.n1 VSUBS 3.5547f
C494 B.n0 VSUBS 0.006259f
C495 B.n1 VSUBS 0.006259f
C496 B.n2 VSUBS 0.009257f
C497 B.n3 VSUBS 0.007094f
C498 B.n4 VSUBS 0.007094f
C499 B.n5 VSUBS 0.007094f
C500 B.n6 VSUBS 0.007094f
C501 B.n7 VSUBS 0.007094f
C502 B.n8 VSUBS 0.007094f
C503 B.n9 VSUBS 0.007094f
C504 B.n10 VSUBS 0.007094f
C505 B.n11 VSUBS 0.007094f
C506 B.n12 VSUBS 0.007094f
C507 B.n13 VSUBS 0.007094f
C508 B.n14 VSUBS 0.007094f
C509 B.n15 VSUBS 0.007094f
C510 B.n16 VSUBS 0.007094f
C511 B.n17 VSUBS 0.007094f
C512 B.n18 VSUBS 0.007094f
C513 B.n19 VSUBS 0.015861f
C514 B.n20 VSUBS 0.007094f
C515 B.n21 VSUBS 0.007094f
C516 B.n22 VSUBS 0.007094f
C517 B.n23 VSUBS 0.007094f
C518 B.n24 VSUBS 0.007094f
C519 B.n25 VSUBS 0.007094f
C520 B.n26 VSUBS 0.007094f
C521 B.n27 VSUBS 0.007094f
C522 B.n28 VSUBS 0.007094f
C523 B.n29 VSUBS 0.007094f
C524 B.n30 VSUBS 0.007094f
C525 B.n31 VSUBS 0.007094f
C526 B.n32 VSUBS 0.007094f
C527 B.n33 VSUBS 0.007094f
C528 B.n34 VSUBS 0.007094f
C529 B.n35 VSUBS 0.007094f
C530 B.n36 VSUBS 0.006676f
C531 B.n37 VSUBS 0.007094f
C532 B.t7 VSUBS 0.159624f
C533 B.t8 VSUBS 0.191528f
C534 B.t6 VSUBS 1.22815f
C535 B.n38 VSUBS 0.310873f
C536 B.n39 VSUBS 0.218825f
C537 B.n40 VSUBS 0.016435f
C538 B.n41 VSUBS 0.007094f
C539 B.n42 VSUBS 0.007094f
C540 B.n43 VSUBS 0.007094f
C541 B.n44 VSUBS 0.007094f
C542 B.t4 VSUBS 0.159627f
C543 B.t5 VSUBS 0.191531f
C544 B.t3 VSUBS 1.22815f
C545 B.n45 VSUBS 0.310871f
C546 B.n46 VSUBS 0.218822f
C547 B.n47 VSUBS 0.007094f
C548 B.n48 VSUBS 0.007094f
C549 B.n49 VSUBS 0.007094f
C550 B.n50 VSUBS 0.007094f
C551 B.n51 VSUBS 0.007094f
C552 B.n52 VSUBS 0.007094f
C553 B.n53 VSUBS 0.007094f
C554 B.n54 VSUBS 0.007094f
C555 B.n55 VSUBS 0.007094f
C556 B.n56 VSUBS 0.007094f
C557 B.n57 VSUBS 0.007094f
C558 B.n58 VSUBS 0.007094f
C559 B.n59 VSUBS 0.007094f
C560 B.n60 VSUBS 0.007094f
C561 B.n61 VSUBS 0.007094f
C562 B.n62 VSUBS 0.007094f
C563 B.n63 VSUBS 0.016269f
C564 B.n64 VSUBS 0.007094f
C565 B.n65 VSUBS 0.007094f
C566 B.n66 VSUBS 0.007094f
C567 B.n67 VSUBS 0.007094f
C568 B.n68 VSUBS 0.007094f
C569 B.n69 VSUBS 0.007094f
C570 B.n70 VSUBS 0.007094f
C571 B.n71 VSUBS 0.007094f
C572 B.n72 VSUBS 0.007094f
C573 B.n73 VSUBS 0.007094f
C574 B.n74 VSUBS 0.007094f
C575 B.n75 VSUBS 0.007094f
C576 B.n76 VSUBS 0.007094f
C577 B.n77 VSUBS 0.007094f
C578 B.n78 VSUBS 0.007094f
C579 B.n79 VSUBS 0.007094f
C580 B.n80 VSUBS 0.007094f
C581 B.n81 VSUBS 0.007094f
C582 B.n82 VSUBS 0.007094f
C583 B.n83 VSUBS 0.007094f
C584 B.n84 VSUBS 0.007094f
C585 B.n85 VSUBS 0.007094f
C586 B.n86 VSUBS 0.007094f
C587 B.n87 VSUBS 0.007094f
C588 B.n88 VSUBS 0.007094f
C589 B.n89 VSUBS 0.007094f
C590 B.n90 VSUBS 0.007094f
C591 B.n91 VSUBS 0.007094f
C592 B.n92 VSUBS 0.007094f
C593 B.n93 VSUBS 0.007094f
C594 B.n94 VSUBS 0.007094f
C595 B.n95 VSUBS 0.007094f
C596 B.n96 VSUBS 0.007094f
C597 B.n97 VSUBS 0.007094f
C598 B.n98 VSUBS 0.007094f
C599 B.n99 VSUBS 0.016742f
C600 B.n100 VSUBS 0.007094f
C601 B.n101 VSUBS 0.007094f
C602 B.n102 VSUBS 0.007094f
C603 B.n103 VSUBS 0.007094f
C604 B.n104 VSUBS 0.007094f
C605 B.n105 VSUBS 0.007094f
C606 B.n106 VSUBS 0.007094f
C607 B.n107 VSUBS 0.007094f
C608 B.n108 VSUBS 0.007094f
C609 B.n109 VSUBS 0.007094f
C610 B.n110 VSUBS 0.007094f
C611 B.n111 VSUBS 0.007094f
C612 B.n112 VSUBS 0.007094f
C613 B.n113 VSUBS 0.007094f
C614 B.n114 VSUBS 0.007094f
C615 B.n115 VSUBS 0.007094f
C616 B.n116 VSUBS 0.007094f
C617 B.t2 VSUBS 0.159627f
C618 B.t1 VSUBS 0.191531f
C619 B.t0 VSUBS 1.22815f
C620 B.n117 VSUBS 0.310871f
C621 B.n118 VSUBS 0.218822f
C622 B.n119 VSUBS 0.007094f
C623 B.n120 VSUBS 0.007094f
C624 B.n121 VSUBS 0.007094f
C625 B.n122 VSUBS 0.007094f
C626 B.n123 VSUBS 0.003964f
C627 B.n124 VSUBS 0.007094f
C628 B.n125 VSUBS 0.007094f
C629 B.n126 VSUBS 0.007094f
C630 B.n127 VSUBS 0.007094f
C631 B.n128 VSUBS 0.007094f
C632 B.n129 VSUBS 0.007094f
C633 B.n130 VSUBS 0.007094f
C634 B.n131 VSUBS 0.007094f
C635 B.n132 VSUBS 0.007094f
C636 B.n133 VSUBS 0.007094f
C637 B.n134 VSUBS 0.007094f
C638 B.n135 VSUBS 0.007094f
C639 B.n136 VSUBS 0.007094f
C640 B.n137 VSUBS 0.007094f
C641 B.n138 VSUBS 0.007094f
C642 B.n139 VSUBS 0.007094f
C643 B.n140 VSUBS 0.016269f
C644 B.n141 VSUBS 0.007094f
C645 B.n142 VSUBS 0.007094f
C646 B.n143 VSUBS 0.007094f
C647 B.n144 VSUBS 0.007094f
C648 B.n145 VSUBS 0.007094f
C649 B.n146 VSUBS 0.007094f
C650 B.n147 VSUBS 0.007094f
C651 B.n148 VSUBS 0.007094f
C652 B.n149 VSUBS 0.007094f
C653 B.n150 VSUBS 0.007094f
C654 B.n151 VSUBS 0.007094f
C655 B.n152 VSUBS 0.007094f
C656 B.n153 VSUBS 0.007094f
C657 B.n154 VSUBS 0.007094f
C658 B.n155 VSUBS 0.007094f
C659 B.n156 VSUBS 0.007094f
C660 B.n157 VSUBS 0.007094f
C661 B.n158 VSUBS 0.007094f
C662 B.n159 VSUBS 0.007094f
C663 B.n160 VSUBS 0.007094f
C664 B.n161 VSUBS 0.007094f
C665 B.n162 VSUBS 0.007094f
C666 B.n163 VSUBS 0.007094f
C667 B.n164 VSUBS 0.007094f
C668 B.n165 VSUBS 0.007094f
C669 B.n166 VSUBS 0.007094f
C670 B.n167 VSUBS 0.007094f
C671 B.n168 VSUBS 0.007094f
C672 B.n169 VSUBS 0.007094f
C673 B.n170 VSUBS 0.007094f
C674 B.n171 VSUBS 0.007094f
C675 B.n172 VSUBS 0.007094f
C676 B.n173 VSUBS 0.007094f
C677 B.n174 VSUBS 0.007094f
C678 B.n175 VSUBS 0.007094f
C679 B.n176 VSUBS 0.007094f
C680 B.n177 VSUBS 0.007094f
C681 B.n178 VSUBS 0.007094f
C682 B.n179 VSUBS 0.007094f
C683 B.n180 VSUBS 0.007094f
C684 B.n181 VSUBS 0.007094f
C685 B.n182 VSUBS 0.007094f
C686 B.n183 VSUBS 0.007094f
C687 B.n184 VSUBS 0.007094f
C688 B.n185 VSUBS 0.007094f
C689 B.n186 VSUBS 0.007094f
C690 B.n187 VSUBS 0.007094f
C691 B.n188 VSUBS 0.007094f
C692 B.n189 VSUBS 0.007094f
C693 B.n190 VSUBS 0.007094f
C694 B.n191 VSUBS 0.007094f
C695 B.n192 VSUBS 0.007094f
C696 B.n193 VSUBS 0.007094f
C697 B.n194 VSUBS 0.007094f
C698 B.n195 VSUBS 0.007094f
C699 B.n196 VSUBS 0.007094f
C700 B.n197 VSUBS 0.007094f
C701 B.n198 VSUBS 0.007094f
C702 B.n199 VSUBS 0.007094f
C703 B.n200 VSUBS 0.007094f
C704 B.n201 VSUBS 0.007094f
C705 B.n202 VSUBS 0.007094f
C706 B.n203 VSUBS 0.007094f
C707 B.n204 VSUBS 0.007094f
C708 B.n205 VSUBS 0.007094f
C709 B.n206 VSUBS 0.007094f
C710 B.n207 VSUBS 0.015861f
C711 B.n208 VSUBS 0.015861f
C712 B.n209 VSUBS 0.016269f
C713 B.n210 VSUBS 0.007094f
C714 B.n211 VSUBS 0.007094f
C715 B.n212 VSUBS 0.007094f
C716 B.n213 VSUBS 0.007094f
C717 B.n214 VSUBS 0.007094f
C718 B.n215 VSUBS 0.007094f
C719 B.n216 VSUBS 0.007094f
C720 B.n217 VSUBS 0.007094f
C721 B.n218 VSUBS 0.007094f
C722 B.n219 VSUBS 0.007094f
C723 B.n220 VSUBS 0.007094f
C724 B.n221 VSUBS 0.007094f
C725 B.n222 VSUBS 0.007094f
C726 B.n223 VSUBS 0.007094f
C727 B.n224 VSUBS 0.007094f
C728 B.n225 VSUBS 0.007094f
C729 B.n226 VSUBS 0.007094f
C730 B.n227 VSUBS 0.007094f
C731 B.n228 VSUBS 0.007094f
C732 B.n229 VSUBS 0.007094f
C733 B.n230 VSUBS 0.007094f
C734 B.n231 VSUBS 0.007094f
C735 B.n232 VSUBS 0.007094f
C736 B.n233 VSUBS 0.007094f
C737 B.n234 VSUBS 0.007094f
C738 B.n235 VSUBS 0.007094f
C739 B.n236 VSUBS 0.007094f
C740 B.n237 VSUBS 0.007094f
C741 B.n238 VSUBS 0.007094f
C742 B.n239 VSUBS 0.007094f
C743 B.n240 VSUBS 0.007094f
C744 B.n241 VSUBS 0.007094f
C745 B.n242 VSUBS 0.007094f
C746 B.n243 VSUBS 0.007094f
C747 B.n244 VSUBS 0.007094f
C748 B.n245 VSUBS 0.007094f
C749 B.n246 VSUBS 0.007094f
C750 B.n247 VSUBS 0.007094f
C751 B.n248 VSUBS 0.007094f
C752 B.n249 VSUBS 0.007094f
C753 B.n250 VSUBS 0.007094f
C754 B.n251 VSUBS 0.007094f
C755 B.n252 VSUBS 0.007094f
C756 B.n253 VSUBS 0.007094f
C757 B.n254 VSUBS 0.007094f
C758 B.n255 VSUBS 0.007094f
C759 B.n256 VSUBS 0.007094f
C760 B.n257 VSUBS 0.007094f
C761 B.t11 VSUBS 0.159624f
C762 B.t10 VSUBS 0.191528f
C763 B.t9 VSUBS 1.22815f
C764 B.n258 VSUBS 0.310873f
C765 B.n259 VSUBS 0.218825f
C766 B.n260 VSUBS 0.016435f
C767 B.n261 VSUBS 0.006676f
C768 B.n262 VSUBS 0.007094f
C769 B.n263 VSUBS 0.007094f
C770 B.n264 VSUBS 0.007094f
C771 B.n265 VSUBS 0.007094f
C772 B.n266 VSUBS 0.007094f
C773 B.n267 VSUBS 0.007094f
C774 B.n268 VSUBS 0.007094f
C775 B.n269 VSUBS 0.007094f
C776 B.n270 VSUBS 0.007094f
C777 B.n271 VSUBS 0.007094f
C778 B.n272 VSUBS 0.007094f
C779 B.n273 VSUBS 0.007094f
C780 B.n274 VSUBS 0.007094f
C781 B.n275 VSUBS 0.007094f
C782 B.n276 VSUBS 0.007094f
C783 B.n277 VSUBS 0.003964f
C784 B.n278 VSUBS 0.016435f
C785 B.n279 VSUBS 0.006676f
C786 B.n280 VSUBS 0.007094f
C787 B.n281 VSUBS 0.007094f
C788 B.n282 VSUBS 0.007094f
C789 B.n283 VSUBS 0.007094f
C790 B.n284 VSUBS 0.007094f
C791 B.n285 VSUBS 0.007094f
C792 B.n286 VSUBS 0.007094f
C793 B.n287 VSUBS 0.007094f
C794 B.n288 VSUBS 0.007094f
C795 B.n289 VSUBS 0.007094f
C796 B.n290 VSUBS 0.007094f
C797 B.n291 VSUBS 0.007094f
C798 B.n292 VSUBS 0.007094f
C799 B.n293 VSUBS 0.007094f
C800 B.n294 VSUBS 0.007094f
C801 B.n295 VSUBS 0.007094f
C802 B.n296 VSUBS 0.007094f
C803 B.n297 VSUBS 0.007094f
C804 B.n298 VSUBS 0.007094f
C805 B.n299 VSUBS 0.007094f
C806 B.n300 VSUBS 0.007094f
C807 B.n301 VSUBS 0.007094f
C808 B.n302 VSUBS 0.007094f
C809 B.n303 VSUBS 0.007094f
C810 B.n304 VSUBS 0.007094f
C811 B.n305 VSUBS 0.007094f
C812 B.n306 VSUBS 0.007094f
C813 B.n307 VSUBS 0.007094f
C814 B.n308 VSUBS 0.007094f
C815 B.n309 VSUBS 0.007094f
C816 B.n310 VSUBS 0.007094f
C817 B.n311 VSUBS 0.007094f
C818 B.n312 VSUBS 0.007094f
C819 B.n313 VSUBS 0.007094f
C820 B.n314 VSUBS 0.007094f
C821 B.n315 VSUBS 0.007094f
C822 B.n316 VSUBS 0.007094f
C823 B.n317 VSUBS 0.007094f
C824 B.n318 VSUBS 0.007094f
C825 B.n319 VSUBS 0.007094f
C826 B.n320 VSUBS 0.007094f
C827 B.n321 VSUBS 0.007094f
C828 B.n322 VSUBS 0.007094f
C829 B.n323 VSUBS 0.007094f
C830 B.n324 VSUBS 0.007094f
C831 B.n325 VSUBS 0.007094f
C832 B.n326 VSUBS 0.007094f
C833 B.n327 VSUBS 0.007094f
C834 B.n328 VSUBS 0.015388f
C835 B.n329 VSUBS 0.016269f
C836 B.n330 VSUBS 0.015861f
C837 B.n331 VSUBS 0.007094f
C838 B.n332 VSUBS 0.007094f
C839 B.n333 VSUBS 0.007094f
C840 B.n334 VSUBS 0.007094f
C841 B.n335 VSUBS 0.007094f
C842 B.n336 VSUBS 0.007094f
C843 B.n337 VSUBS 0.007094f
C844 B.n338 VSUBS 0.007094f
C845 B.n339 VSUBS 0.007094f
C846 B.n340 VSUBS 0.007094f
C847 B.n341 VSUBS 0.007094f
C848 B.n342 VSUBS 0.007094f
C849 B.n343 VSUBS 0.007094f
C850 B.n344 VSUBS 0.007094f
C851 B.n345 VSUBS 0.007094f
C852 B.n346 VSUBS 0.007094f
C853 B.n347 VSUBS 0.007094f
C854 B.n348 VSUBS 0.007094f
C855 B.n349 VSUBS 0.007094f
C856 B.n350 VSUBS 0.007094f
C857 B.n351 VSUBS 0.007094f
C858 B.n352 VSUBS 0.007094f
C859 B.n353 VSUBS 0.007094f
C860 B.n354 VSUBS 0.007094f
C861 B.n355 VSUBS 0.007094f
C862 B.n356 VSUBS 0.007094f
C863 B.n357 VSUBS 0.007094f
C864 B.n358 VSUBS 0.007094f
C865 B.n359 VSUBS 0.007094f
C866 B.n360 VSUBS 0.007094f
C867 B.n361 VSUBS 0.007094f
C868 B.n362 VSUBS 0.007094f
C869 B.n363 VSUBS 0.007094f
C870 B.n364 VSUBS 0.007094f
C871 B.n365 VSUBS 0.007094f
C872 B.n366 VSUBS 0.007094f
C873 B.n367 VSUBS 0.007094f
C874 B.n368 VSUBS 0.007094f
C875 B.n369 VSUBS 0.007094f
C876 B.n370 VSUBS 0.007094f
C877 B.n371 VSUBS 0.007094f
C878 B.n372 VSUBS 0.007094f
C879 B.n373 VSUBS 0.007094f
C880 B.n374 VSUBS 0.007094f
C881 B.n375 VSUBS 0.007094f
C882 B.n376 VSUBS 0.007094f
C883 B.n377 VSUBS 0.007094f
C884 B.n378 VSUBS 0.007094f
C885 B.n379 VSUBS 0.007094f
C886 B.n380 VSUBS 0.007094f
C887 B.n381 VSUBS 0.007094f
C888 B.n382 VSUBS 0.007094f
C889 B.n383 VSUBS 0.007094f
C890 B.n384 VSUBS 0.007094f
C891 B.n385 VSUBS 0.007094f
C892 B.n386 VSUBS 0.007094f
C893 B.n387 VSUBS 0.007094f
C894 B.n388 VSUBS 0.007094f
C895 B.n389 VSUBS 0.007094f
C896 B.n390 VSUBS 0.007094f
C897 B.n391 VSUBS 0.007094f
C898 B.n392 VSUBS 0.007094f
C899 B.n393 VSUBS 0.007094f
C900 B.n394 VSUBS 0.007094f
C901 B.n395 VSUBS 0.007094f
C902 B.n396 VSUBS 0.007094f
C903 B.n397 VSUBS 0.007094f
C904 B.n398 VSUBS 0.007094f
C905 B.n399 VSUBS 0.007094f
C906 B.n400 VSUBS 0.007094f
C907 B.n401 VSUBS 0.007094f
C908 B.n402 VSUBS 0.007094f
C909 B.n403 VSUBS 0.007094f
C910 B.n404 VSUBS 0.007094f
C911 B.n405 VSUBS 0.007094f
C912 B.n406 VSUBS 0.007094f
C913 B.n407 VSUBS 0.007094f
C914 B.n408 VSUBS 0.007094f
C915 B.n409 VSUBS 0.007094f
C916 B.n410 VSUBS 0.007094f
C917 B.n411 VSUBS 0.007094f
C918 B.n412 VSUBS 0.007094f
C919 B.n413 VSUBS 0.007094f
C920 B.n414 VSUBS 0.007094f
C921 B.n415 VSUBS 0.007094f
C922 B.n416 VSUBS 0.007094f
C923 B.n417 VSUBS 0.007094f
C924 B.n418 VSUBS 0.007094f
C925 B.n419 VSUBS 0.007094f
C926 B.n420 VSUBS 0.007094f
C927 B.n421 VSUBS 0.007094f
C928 B.n422 VSUBS 0.007094f
C929 B.n423 VSUBS 0.007094f
C930 B.n424 VSUBS 0.007094f
C931 B.n425 VSUBS 0.007094f
C932 B.n426 VSUBS 0.007094f
C933 B.n427 VSUBS 0.007094f
C934 B.n428 VSUBS 0.007094f
C935 B.n429 VSUBS 0.007094f
C936 B.n430 VSUBS 0.007094f
C937 B.n431 VSUBS 0.007094f
C938 B.n432 VSUBS 0.007094f
C939 B.n433 VSUBS 0.007094f
C940 B.n434 VSUBS 0.007094f
C941 B.n435 VSUBS 0.007094f
C942 B.n436 VSUBS 0.015861f
C943 B.n437 VSUBS 0.015861f
C944 B.n438 VSUBS 0.016269f
C945 B.n439 VSUBS 0.007094f
C946 B.n440 VSUBS 0.007094f
C947 B.n441 VSUBS 0.007094f
C948 B.n442 VSUBS 0.007094f
C949 B.n443 VSUBS 0.007094f
C950 B.n444 VSUBS 0.007094f
C951 B.n445 VSUBS 0.007094f
C952 B.n446 VSUBS 0.007094f
C953 B.n447 VSUBS 0.007094f
C954 B.n448 VSUBS 0.007094f
C955 B.n449 VSUBS 0.007094f
C956 B.n450 VSUBS 0.007094f
C957 B.n451 VSUBS 0.007094f
C958 B.n452 VSUBS 0.007094f
C959 B.n453 VSUBS 0.007094f
C960 B.n454 VSUBS 0.007094f
C961 B.n455 VSUBS 0.007094f
C962 B.n456 VSUBS 0.007094f
C963 B.n457 VSUBS 0.007094f
C964 B.n458 VSUBS 0.007094f
C965 B.n459 VSUBS 0.007094f
C966 B.n460 VSUBS 0.007094f
C967 B.n461 VSUBS 0.007094f
C968 B.n462 VSUBS 0.007094f
C969 B.n463 VSUBS 0.007094f
C970 B.n464 VSUBS 0.007094f
C971 B.n465 VSUBS 0.007094f
C972 B.n466 VSUBS 0.007094f
C973 B.n467 VSUBS 0.007094f
C974 B.n468 VSUBS 0.007094f
C975 B.n469 VSUBS 0.007094f
C976 B.n470 VSUBS 0.007094f
C977 B.n471 VSUBS 0.007094f
C978 B.n472 VSUBS 0.007094f
C979 B.n473 VSUBS 0.007094f
C980 B.n474 VSUBS 0.007094f
C981 B.n475 VSUBS 0.007094f
C982 B.n476 VSUBS 0.007094f
C983 B.n477 VSUBS 0.007094f
C984 B.n478 VSUBS 0.007094f
C985 B.n479 VSUBS 0.007094f
C986 B.n480 VSUBS 0.007094f
C987 B.n481 VSUBS 0.007094f
C988 B.n482 VSUBS 0.007094f
C989 B.n483 VSUBS 0.007094f
C990 B.n484 VSUBS 0.007094f
C991 B.n485 VSUBS 0.007094f
C992 B.n486 VSUBS 0.007094f
C993 B.n487 VSUBS 0.007094f
C994 B.n488 VSUBS 0.006676f
C995 B.n489 VSUBS 0.016435f
C996 B.n490 VSUBS 0.003964f
C997 B.n491 VSUBS 0.007094f
C998 B.n492 VSUBS 0.007094f
C999 B.n493 VSUBS 0.007094f
C1000 B.n494 VSUBS 0.007094f
C1001 B.n495 VSUBS 0.007094f
C1002 B.n496 VSUBS 0.007094f
C1003 B.n497 VSUBS 0.007094f
C1004 B.n498 VSUBS 0.007094f
C1005 B.n499 VSUBS 0.007094f
C1006 B.n500 VSUBS 0.007094f
C1007 B.n501 VSUBS 0.007094f
C1008 B.n502 VSUBS 0.007094f
C1009 B.n503 VSUBS 0.003964f
C1010 B.n504 VSUBS 0.007094f
C1011 B.n505 VSUBS 0.007094f
C1012 B.n506 VSUBS 0.007094f
C1013 B.n507 VSUBS 0.007094f
C1014 B.n508 VSUBS 0.007094f
C1015 B.n509 VSUBS 0.007094f
C1016 B.n510 VSUBS 0.007094f
C1017 B.n511 VSUBS 0.007094f
C1018 B.n512 VSUBS 0.007094f
C1019 B.n513 VSUBS 0.007094f
C1020 B.n514 VSUBS 0.007094f
C1021 B.n515 VSUBS 0.007094f
C1022 B.n516 VSUBS 0.007094f
C1023 B.n517 VSUBS 0.007094f
C1024 B.n518 VSUBS 0.007094f
C1025 B.n519 VSUBS 0.007094f
C1026 B.n520 VSUBS 0.007094f
C1027 B.n521 VSUBS 0.007094f
C1028 B.n522 VSUBS 0.007094f
C1029 B.n523 VSUBS 0.007094f
C1030 B.n524 VSUBS 0.007094f
C1031 B.n525 VSUBS 0.007094f
C1032 B.n526 VSUBS 0.007094f
C1033 B.n527 VSUBS 0.007094f
C1034 B.n528 VSUBS 0.007094f
C1035 B.n529 VSUBS 0.007094f
C1036 B.n530 VSUBS 0.007094f
C1037 B.n531 VSUBS 0.007094f
C1038 B.n532 VSUBS 0.007094f
C1039 B.n533 VSUBS 0.007094f
C1040 B.n534 VSUBS 0.007094f
C1041 B.n535 VSUBS 0.007094f
C1042 B.n536 VSUBS 0.007094f
C1043 B.n537 VSUBS 0.007094f
C1044 B.n538 VSUBS 0.007094f
C1045 B.n539 VSUBS 0.007094f
C1046 B.n540 VSUBS 0.007094f
C1047 B.n541 VSUBS 0.007094f
C1048 B.n542 VSUBS 0.007094f
C1049 B.n543 VSUBS 0.007094f
C1050 B.n544 VSUBS 0.007094f
C1051 B.n545 VSUBS 0.007094f
C1052 B.n546 VSUBS 0.007094f
C1053 B.n547 VSUBS 0.007094f
C1054 B.n548 VSUBS 0.007094f
C1055 B.n549 VSUBS 0.007094f
C1056 B.n550 VSUBS 0.007094f
C1057 B.n551 VSUBS 0.007094f
C1058 B.n552 VSUBS 0.007094f
C1059 B.n553 VSUBS 0.007094f
C1060 B.n554 VSUBS 0.016269f
C1061 B.n555 VSUBS 0.016269f
C1062 B.n556 VSUBS 0.015861f
C1063 B.n557 VSUBS 0.007094f
C1064 B.n558 VSUBS 0.007094f
C1065 B.n559 VSUBS 0.007094f
C1066 B.n560 VSUBS 0.007094f
C1067 B.n561 VSUBS 0.007094f
C1068 B.n562 VSUBS 0.007094f
C1069 B.n563 VSUBS 0.007094f
C1070 B.n564 VSUBS 0.007094f
C1071 B.n565 VSUBS 0.007094f
C1072 B.n566 VSUBS 0.007094f
C1073 B.n567 VSUBS 0.007094f
C1074 B.n568 VSUBS 0.007094f
C1075 B.n569 VSUBS 0.007094f
C1076 B.n570 VSUBS 0.007094f
C1077 B.n571 VSUBS 0.007094f
C1078 B.n572 VSUBS 0.007094f
C1079 B.n573 VSUBS 0.007094f
C1080 B.n574 VSUBS 0.007094f
C1081 B.n575 VSUBS 0.007094f
C1082 B.n576 VSUBS 0.007094f
C1083 B.n577 VSUBS 0.007094f
C1084 B.n578 VSUBS 0.007094f
C1085 B.n579 VSUBS 0.007094f
C1086 B.n580 VSUBS 0.007094f
C1087 B.n581 VSUBS 0.007094f
C1088 B.n582 VSUBS 0.007094f
C1089 B.n583 VSUBS 0.007094f
C1090 B.n584 VSUBS 0.007094f
C1091 B.n585 VSUBS 0.007094f
C1092 B.n586 VSUBS 0.007094f
C1093 B.n587 VSUBS 0.007094f
C1094 B.n588 VSUBS 0.007094f
C1095 B.n589 VSUBS 0.007094f
C1096 B.n590 VSUBS 0.007094f
C1097 B.n591 VSUBS 0.007094f
C1098 B.n592 VSUBS 0.007094f
C1099 B.n593 VSUBS 0.007094f
C1100 B.n594 VSUBS 0.007094f
C1101 B.n595 VSUBS 0.007094f
C1102 B.n596 VSUBS 0.007094f
C1103 B.n597 VSUBS 0.007094f
C1104 B.n598 VSUBS 0.007094f
C1105 B.n599 VSUBS 0.007094f
C1106 B.n600 VSUBS 0.007094f
C1107 B.n601 VSUBS 0.007094f
C1108 B.n602 VSUBS 0.007094f
C1109 B.n603 VSUBS 0.007094f
C1110 B.n604 VSUBS 0.007094f
C1111 B.n605 VSUBS 0.007094f
C1112 B.n606 VSUBS 0.007094f
C1113 B.n607 VSUBS 0.009257f
C1114 B.n608 VSUBS 0.009861f
C1115 B.n609 VSUBS 0.019609f
.ends

