* NGSPICE file created from diff_pair_sample_0281.ext - technology: sky130A

.subckt diff_pair_sample_0281 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t7 VP.t0 VTAIL.t14 w_n3410_n2636# sky130_fd_pr__pfet_01v8 ad=1.3761 pd=8.67 as=3.2526 ps=17.46 w=8.34 l=2.11
X1 VDD2.t7 VN.t0 VTAIL.t2 w_n3410_n2636# sky130_fd_pr__pfet_01v8 ad=1.3761 pd=8.67 as=3.2526 ps=17.46 w=8.34 l=2.11
X2 VDD2.t6 VN.t1 VTAIL.t7 w_n3410_n2636# sky130_fd_pr__pfet_01v8 ad=1.3761 pd=8.67 as=1.3761 ps=8.67 w=8.34 l=2.11
X3 VDD1.t6 VP.t1 VTAIL.t12 w_n3410_n2636# sky130_fd_pr__pfet_01v8 ad=1.3761 pd=8.67 as=1.3761 ps=8.67 w=8.34 l=2.11
X4 VTAIL.t13 VP.t2 VDD1.t5 w_n3410_n2636# sky130_fd_pr__pfet_01v8 ad=3.2526 pd=17.46 as=1.3761 ps=8.67 w=8.34 l=2.11
X5 VDD2.t5 VN.t2 VTAIL.t6 w_n3410_n2636# sky130_fd_pr__pfet_01v8 ad=1.3761 pd=8.67 as=1.3761 ps=8.67 w=8.34 l=2.11
X6 VDD2.t4 VN.t3 VTAIL.t0 w_n3410_n2636# sky130_fd_pr__pfet_01v8 ad=1.3761 pd=8.67 as=3.2526 ps=17.46 w=8.34 l=2.11
X7 B.t11 B.t9 B.t10 w_n3410_n2636# sky130_fd_pr__pfet_01v8 ad=3.2526 pd=17.46 as=0 ps=0 w=8.34 l=2.11
X8 VTAIL.t10 VP.t3 VDD1.t4 w_n3410_n2636# sky130_fd_pr__pfet_01v8 ad=1.3761 pd=8.67 as=1.3761 ps=8.67 w=8.34 l=2.11
X9 B.t8 B.t6 B.t7 w_n3410_n2636# sky130_fd_pr__pfet_01v8 ad=3.2526 pd=17.46 as=0 ps=0 w=8.34 l=2.11
X10 B.t5 B.t3 B.t4 w_n3410_n2636# sky130_fd_pr__pfet_01v8 ad=3.2526 pd=17.46 as=0 ps=0 w=8.34 l=2.11
X11 VTAIL.t11 VP.t4 VDD1.t3 w_n3410_n2636# sky130_fd_pr__pfet_01v8 ad=1.3761 pd=8.67 as=1.3761 ps=8.67 w=8.34 l=2.11
X12 VTAIL.t4 VN.t4 VDD2.t3 w_n3410_n2636# sky130_fd_pr__pfet_01v8 ad=3.2526 pd=17.46 as=1.3761 ps=8.67 w=8.34 l=2.11
X13 B.t2 B.t0 B.t1 w_n3410_n2636# sky130_fd_pr__pfet_01v8 ad=3.2526 pd=17.46 as=0 ps=0 w=8.34 l=2.11
X14 VTAIL.t5 VN.t5 VDD2.t2 w_n3410_n2636# sky130_fd_pr__pfet_01v8 ad=1.3761 pd=8.67 as=1.3761 ps=8.67 w=8.34 l=2.11
X15 VDD1.t2 VP.t5 VTAIL.t8 w_n3410_n2636# sky130_fd_pr__pfet_01v8 ad=1.3761 pd=8.67 as=3.2526 ps=17.46 w=8.34 l=2.11
X16 VTAIL.t1 VN.t6 VDD2.t1 w_n3410_n2636# sky130_fd_pr__pfet_01v8 ad=1.3761 pd=8.67 as=1.3761 ps=8.67 w=8.34 l=2.11
X17 VTAIL.t3 VN.t7 VDD2.t0 w_n3410_n2636# sky130_fd_pr__pfet_01v8 ad=3.2526 pd=17.46 as=1.3761 ps=8.67 w=8.34 l=2.11
X18 VDD1.t1 VP.t6 VTAIL.t15 w_n3410_n2636# sky130_fd_pr__pfet_01v8 ad=1.3761 pd=8.67 as=1.3761 ps=8.67 w=8.34 l=2.11
X19 VTAIL.t9 VP.t7 VDD1.t0 w_n3410_n2636# sky130_fd_pr__pfet_01v8 ad=3.2526 pd=17.46 as=1.3761 ps=8.67 w=8.34 l=2.11
R0 VP.n15 VP.n12 161.3
R1 VP.n17 VP.n16 161.3
R2 VP.n18 VP.n11 161.3
R3 VP.n20 VP.n19 161.3
R4 VP.n22 VP.n10 161.3
R5 VP.n24 VP.n23 161.3
R6 VP.n25 VP.n9 161.3
R7 VP.n27 VP.n26 161.3
R8 VP.n28 VP.n8 161.3
R9 VP.n54 VP.n0 161.3
R10 VP.n53 VP.n52 161.3
R11 VP.n51 VP.n1 161.3
R12 VP.n50 VP.n49 161.3
R13 VP.n48 VP.n2 161.3
R14 VP.n46 VP.n45 161.3
R15 VP.n44 VP.n3 161.3
R16 VP.n43 VP.n42 161.3
R17 VP.n41 VP.n4 161.3
R18 VP.n39 VP.n38 161.3
R19 VP.n37 VP.n5 161.3
R20 VP.n36 VP.n35 161.3
R21 VP.n34 VP.n6 161.3
R22 VP.n33 VP.n32 161.3
R23 VP.n13 VP.t7 129.504
R24 VP.n7 VP.t2 95.2583
R25 VP.n40 VP.t6 95.2583
R26 VP.n47 VP.t3 95.2583
R27 VP.n55 VP.t0 95.2583
R28 VP.n29 VP.t5 95.2583
R29 VP.n21 VP.t4 95.2583
R30 VP.n14 VP.t1 95.2583
R31 VP.n31 VP.n7 90.7429
R32 VP.n56 VP.n55 90.7429
R33 VP.n30 VP.n29 90.7429
R34 VP.n35 VP.n34 56.5617
R35 VP.n42 VP.n3 56.5617
R36 VP.n53 VP.n1 56.5617
R37 VP.n27 VP.n9 56.5617
R38 VP.n16 VP.n11 56.5617
R39 VP.n14 VP.n13 47.6568
R40 VP.n31 VP.n30 45.886
R41 VP.n34 VP.n33 24.5923
R42 VP.n35 VP.n5 24.5923
R43 VP.n39 VP.n5 24.5923
R44 VP.n42 VP.n41 24.5923
R45 VP.n46 VP.n3 24.5923
R46 VP.n49 VP.n48 24.5923
R47 VP.n49 VP.n1 24.5923
R48 VP.n54 VP.n53 24.5923
R49 VP.n28 VP.n27 24.5923
R50 VP.n20 VP.n11 24.5923
R51 VP.n23 VP.n22 24.5923
R52 VP.n23 VP.n9 24.5923
R53 VP.n16 VP.n15 24.5923
R54 VP.n41 VP.n40 23.1168
R55 VP.n47 VP.n46 23.1168
R56 VP.n21 VP.n20 23.1168
R57 VP.n15 VP.n14 23.1168
R58 VP.n33 VP.n7 20.1658
R59 VP.n55 VP.n54 20.1658
R60 VP.n29 VP.n28 20.1658
R61 VP.n13 VP.n12 8.94243
R62 VP.n40 VP.n39 1.47601
R63 VP.n48 VP.n47 1.47601
R64 VP.n22 VP.n21 1.47601
R65 VP.n30 VP.n8 0.278335
R66 VP.n32 VP.n31 0.278335
R67 VP.n56 VP.n0 0.278335
R68 VP.n17 VP.n12 0.189894
R69 VP.n18 VP.n17 0.189894
R70 VP.n19 VP.n18 0.189894
R71 VP.n19 VP.n10 0.189894
R72 VP.n24 VP.n10 0.189894
R73 VP.n25 VP.n24 0.189894
R74 VP.n26 VP.n25 0.189894
R75 VP.n26 VP.n8 0.189894
R76 VP.n32 VP.n6 0.189894
R77 VP.n36 VP.n6 0.189894
R78 VP.n37 VP.n36 0.189894
R79 VP.n38 VP.n37 0.189894
R80 VP.n38 VP.n4 0.189894
R81 VP.n43 VP.n4 0.189894
R82 VP.n44 VP.n43 0.189894
R83 VP.n45 VP.n44 0.189894
R84 VP.n45 VP.n2 0.189894
R85 VP.n50 VP.n2 0.189894
R86 VP.n51 VP.n50 0.189894
R87 VP.n52 VP.n51 0.189894
R88 VP.n52 VP.n0 0.189894
R89 VP VP.n56 0.153485
R90 VTAIL.n11 VTAIL.t9 71.9944
R91 VTAIL.n10 VTAIL.t0 71.9944
R92 VTAIL.n7 VTAIL.t4 71.9944
R93 VTAIL.n15 VTAIL.t2 71.9943
R94 VTAIL.n2 VTAIL.t3 71.9943
R95 VTAIL.n3 VTAIL.t14 71.9943
R96 VTAIL.n6 VTAIL.t13 71.9943
R97 VTAIL.n14 VTAIL.t8 71.9943
R98 VTAIL.n13 VTAIL.n12 68.097
R99 VTAIL.n9 VTAIL.n8 68.097
R100 VTAIL.n1 VTAIL.n0 68.0967
R101 VTAIL.n5 VTAIL.n4 68.0967
R102 VTAIL.n15 VTAIL.n14 21.66
R103 VTAIL.n7 VTAIL.n6 21.66
R104 VTAIL.n0 VTAIL.t7 3.89798
R105 VTAIL.n0 VTAIL.t1 3.89798
R106 VTAIL.n4 VTAIL.t15 3.89798
R107 VTAIL.n4 VTAIL.t10 3.89798
R108 VTAIL.n12 VTAIL.t12 3.89798
R109 VTAIL.n12 VTAIL.t11 3.89798
R110 VTAIL.n8 VTAIL.t6 3.89798
R111 VTAIL.n8 VTAIL.t5 3.89798
R112 VTAIL.n9 VTAIL.n7 2.10395
R113 VTAIL.n10 VTAIL.n9 2.10395
R114 VTAIL.n13 VTAIL.n11 2.10395
R115 VTAIL.n14 VTAIL.n13 2.10395
R116 VTAIL.n6 VTAIL.n5 2.10395
R117 VTAIL.n5 VTAIL.n3 2.10395
R118 VTAIL.n2 VTAIL.n1 2.10395
R119 VTAIL VTAIL.n15 2.04576
R120 VTAIL.n11 VTAIL.n10 0.470328
R121 VTAIL.n3 VTAIL.n2 0.470328
R122 VTAIL VTAIL.n1 0.0586897
R123 VDD1 VDD1.n0 85.8857
R124 VDD1.n3 VDD1.n2 85.7719
R125 VDD1.n3 VDD1.n1 85.7719
R126 VDD1.n5 VDD1.n4 84.7756
R127 VDD1.n5 VDD1.n3 40.9535
R128 VDD1.n4 VDD1.t3 3.89798
R129 VDD1.n4 VDD1.t2 3.89798
R130 VDD1.n0 VDD1.t0 3.89798
R131 VDD1.n0 VDD1.t6 3.89798
R132 VDD1.n2 VDD1.t4 3.89798
R133 VDD1.n2 VDD1.t7 3.89798
R134 VDD1.n1 VDD1.t5 3.89798
R135 VDD1.n1 VDD1.t1 3.89798
R136 VDD1 VDD1.n5 0.994035
R137 VN.n43 VN.n23 161.3
R138 VN.n42 VN.n41 161.3
R139 VN.n40 VN.n24 161.3
R140 VN.n39 VN.n38 161.3
R141 VN.n37 VN.n25 161.3
R142 VN.n35 VN.n34 161.3
R143 VN.n33 VN.n26 161.3
R144 VN.n32 VN.n31 161.3
R145 VN.n30 VN.n27 161.3
R146 VN.n20 VN.n0 161.3
R147 VN.n19 VN.n18 161.3
R148 VN.n17 VN.n1 161.3
R149 VN.n16 VN.n15 161.3
R150 VN.n14 VN.n2 161.3
R151 VN.n12 VN.n11 161.3
R152 VN.n10 VN.n3 161.3
R153 VN.n9 VN.n8 161.3
R154 VN.n7 VN.n4 161.3
R155 VN.n5 VN.t7 129.504
R156 VN.n28 VN.t3 129.504
R157 VN.n6 VN.t1 95.2583
R158 VN.n13 VN.t6 95.2583
R159 VN.n21 VN.t0 95.2583
R160 VN.n29 VN.t5 95.2583
R161 VN.n36 VN.t2 95.2583
R162 VN.n44 VN.t4 95.2583
R163 VN.n22 VN.n21 90.7429
R164 VN.n45 VN.n44 90.7429
R165 VN.n8 VN.n3 56.5617
R166 VN.n19 VN.n1 56.5617
R167 VN.n31 VN.n26 56.5617
R168 VN.n42 VN.n24 56.5617
R169 VN.n6 VN.n5 47.6568
R170 VN.n29 VN.n28 47.6568
R171 VN VN.n45 46.1649
R172 VN.n8 VN.n7 24.5923
R173 VN.n12 VN.n3 24.5923
R174 VN.n15 VN.n14 24.5923
R175 VN.n15 VN.n1 24.5923
R176 VN.n20 VN.n19 24.5923
R177 VN.n31 VN.n30 24.5923
R178 VN.n38 VN.n24 24.5923
R179 VN.n38 VN.n37 24.5923
R180 VN.n35 VN.n26 24.5923
R181 VN.n43 VN.n42 24.5923
R182 VN.n7 VN.n6 23.1168
R183 VN.n13 VN.n12 23.1168
R184 VN.n30 VN.n29 23.1168
R185 VN.n36 VN.n35 23.1168
R186 VN.n21 VN.n20 20.1658
R187 VN.n44 VN.n43 20.1658
R188 VN.n28 VN.n27 8.94243
R189 VN.n5 VN.n4 8.94243
R190 VN.n14 VN.n13 1.47601
R191 VN.n37 VN.n36 1.47601
R192 VN.n45 VN.n23 0.278335
R193 VN.n22 VN.n0 0.278335
R194 VN.n41 VN.n23 0.189894
R195 VN.n41 VN.n40 0.189894
R196 VN.n40 VN.n39 0.189894
R197 VN.n39 VN.n25 0.189894
R198 VN.n34 VN.n25 0.189894
R199 VN.n34 VN.n33 0.189894
R200 VN.n33 VN.n32 0.189894
R201 VN.n32 VN.n27 0.189894
R202 VN.n9 VN.n4 0.189894
R203 VN.n10 VN.n9 0.189894
R204 VN.n11 VN.n10 0.189894
R205 VN.n11 VN.n2 0.189894
R206 VN.n16 VN.n2 0.189894
R207 VN.n17 VN.n16 0.189894
R208 VN.n18 VN.n17 0.189894
R209 VN.n18 VN.n0 0.189894
R210 VN VN.n22 0.153485
R211 VDD2.n2 VDD2.n1 85.7719
R212 VDD2.n2 VDD2.n0 85.7719
R213 VDD2 VDD2.n5 85.7691
R214 VDD2.n4 VDD2.n3 84.7758
R215 VDD2.n4 VDD2.n2 40.3705
R216 VDD2.n5 VDD2.t2 3.89798
R217 VDD2.n5 VDD2.t4 3.89798
R218 VDD2.n3 VDD2.t3 3.89798
R219 VDD2.n3 VDD2.t5 3.89798
R220 VDD2.n1 VDD2.t1 3.89798
R221 VDD2.n1 VDD2.t7 3.89798
R222 VDD2.n0 VDD2.t0 3.89798
R223 VDD2.n0 VDD2.t6 3.89798
R224 VDD2 VDD2.n4 1.11041
R225 B.n477 B.n476 585
R226 B.n478 B.n63 585
R227 B.n480 B.n479 585
R228 B.n481 B.n62 585
R229 B.n483 B.n482 585
R230 B.n484 B.n61 585
R231 B.n486 B.n485 585
R232 B.n487 B.n60 585
R233 B.n489 B.n488 585
R234 B.n490 B.n59 585
R235 B.n492 B.n491 585
R236 B.n493 B.n58 585
R237 B.n495 B.n494 585
R238 B.n496 B.n57 585
R239 B.n498 B.n497 585
R240 B.n499 B.n56 585
R241 B.n501 B.n500 585
R242 B.n502 B.n55 585
R243 B.n504 B.n503 585
R244 B.n505 B.n54 585
R245 B.n507 B.n506 585
R246 B.n508 B.n53 585
R247 B.n510 B.n509 585
R248 B.n511 B.n52 585
R249 B.n513 B.n512 585
R250 B.n514 B.n51 585
R251 B.n516 B.n515 585
R252 B.n517 B.n50 585
R253 B.n519 B.n518 585
R254 B.n520 B.n49 585
R255 B.n522 B.n521 585
R256 B.n524 B.n523 585
R257 B.n525 B.n45 585
R258 B.n527 B.n526 585
R259 B.n528 B.n44 585
R260 B.n530 B.n529 585
R261 B.n531 B.n43 585
R262 B.n533 B.n532 585
R263 B.n534 B.n42 585
R264 B.n536 B.n535 585
R265 B.n538 B.n39 585
R266 B.n540 B.n539 585
R267 B.n541 B.n38 585
R268 B.n543 B.n542 585
R269 B.n544 B.n37 585
R270 B.n546 B.n545 585
R271 B.n547 B.n36 585
R272 B.n549 B.n548 585
R273 B.n550 B.n35 585
R274 B.n552 B.n551 585
R275 B.n553 B.n34 585
R276 B.n555 B.n554 585
R277 B.n556 B.n33 585
R278 B.n558 B.n557 585
R279 B.n559 B.n32 585
R280 B.n561 B.n560 585
R281 B.n562 B.n31 585
R282 B.n564 B.n563 585
R283 B.n565 B.n30 585
R284 B.n567 B.n566 585
R285 B.n568 B.n29 585
R286 B.n570 B.n569 585
R287 B.n571 B.n28 585
R288 B.n573 B.n572 585
R289 B.n574 B.n27 585
R290 B.n576 B.n575 585
R291 B.n577 B.n26 585
R292 B.n579 B.n578 585
R293 B.n580 B.n25 585
R294 B.n582 B.n581 585
R295 B.n583 B.n24 585
R296 B.n475 B.n64 585
R297 B.n474 B.n473 585
R298 B.n472 B.n65 585
R299 B.n471 B.n470 585
R300 B.n469 B.n66 585
R301 B.n468 B.n467 585
R302 B.n466 B.n67 585
R303 B.n465 B.n464 585
R304 B.n463 B.n68 585
R305 B.n462 B.n461 585
R306 B.n460 B.n69 585
R307 B.n459 B.n458 585
R308 B.n457 B.n70 585
R309 B.n456 B.n455 585
R310 B.n454 B.n71 585
R311 B.n453 B.n452 585
R312 B.n451 B.n72 585
R313 B.n450 B.n449 585
R314 B.n448 B.n73 585
R315 B.n447 B.n446 585
R316 B.n445 B.n74 585
R317 B.n444 B.n443 585
R318 B.n442 B.n75 585
R319 B.n441 B.n440 585
R320 B.n439 B.n76 585
R321 B.n438 B.n437 585
R322 B.n436 B.n77 585
R323 B.n435 B.n434 585
R324 B.n433 B.n78 585
R325 B.n432 B.n431 585
R326 B.n430 B.n79 585
R327 B.n429 B.n428 585
R328 B.n427 B.n80 585
R329 B.n426 B.n425 585
R330 B.n424 B.n81 585
R331 B.n423 B.n422 585
R332 B.n421 B.n82 585
R333 B.n420 B.n419 585
R334 B.n418 B.n83 585
R335 B.n417 B.n416 585
R336 B.n415 B.n84 585
R337 B.n414 B.n413 585
R338 B.n412 B.n85 585
R339 B.n411 B.n410 585
R340 B.n409 B.n86 585
R341 B.n408 B.n407 585
R342 B.n406 B.n87 585
R343 B.n405 B.n404 585
R344 B.n403 B.n88 585
R345 B.n402 B.n401 585
R346 B.n400 B.n89 585
R347 B.n399 B.n398 585
R348 B.n397 B.n90 585
R349 B.n396 B.n395 585
R350 B.n394 B.n91 585
R351 B.n393 B.n392 585
R352 B.n391 B.n92 585
R353 B.n390 B.n389 585
R354 B.n388 B.n93 585
R355 B.n387 B.n386 585
R356 B.n385 B.n94 585
R357 B.n384 B.n383 585
R358 B.n382 B.n95 585
R359 B.n381 B.n380 585
R360 B.n379 B.n96 585
R361 B.n378 B.n377 585
R362 B.n376 B.n97 585
R363 B.n375 B.n374 585
R364 B.n373 B.n98 585
R365 B.n372 B.n371 585
R366 B.n370 B.n99 585
R367 B.n369 B.n368 585
R368 B.n367 B.n100 585
R369 B.n366 B.n365 585
R370 B.n364 B.n101 585
R371 B.n363 B.n362 585
R372 B.n361 B.n102 585
R373 B.n360 B.n359 585
R374 B.n358 B.n103 585
R375 B.n357 B.n356 585
R376 B.n355 B.n104 585
R377 B.n354 B.n353 585
R378 B.n352 B.n105 585
R379 B.n351 B.n350 585
R380 B.n349 B.n106 585
R381 B.n348 B.n347 585
R382 B.n346 B.n107 585
R383 B.n345 B.n344 585
R384 B.n343 B.n108 585
R385 B.n235 B.n148 585
R386 B.n237 B.n236 585
R387 B.n238 B.n147 585
R388 B.n240 B.n239 585
R389 B.n241 B.n146 585
R390 B.n243 B.n242 585
R391 B.n244 B.n145 585
R392 B.n246 B.n245 585
R393 B.n247 B.n144 585
R394 B.n249 B.n248 585
R395 B.n250 B.n143 585
R396 B.n252 B.n251 585
R397 B.n253 B.n142 585
R398 B.n255 B.n254 585
R399 B.n256 B.n141 585
R400 B.n258 B.n257 585
R401 B.n259 B.n140 585
R402 B.n261 B.n260 585
R403 B.n262 B.n139 585
R404 B.n264 B.n263 585
R405 B.n265 B.n138 585
R406 B.n267 B.n266 585
R407 B.n268 B.n137 585
R408 B.n270 B.n269 585
R409 B.n271 B.n136 585
R410 B.n273 B.n272 585
R411 B.n274 B.n135 585
R412 B.n276 B.n275 585
R413 B.n277 B.n134 585
R414 B.n279 B.n278 585
R415 B.n280 B.n131 585
R416 B.n283 B.n282 585
R417 B.n284 B.n130 585
R418 B.n286 B.n285 585
R419 B.n287 B.n129 585
R420 B.n289 B.n288 585
R421 B.n290 B.n128 585
R422 B.n292 B.n291 585
R423 B.n293 B.n127 585
R424 B.n295 B.n294 585
R425 B.n297 B.n296 585
R426 B.n298 B.n123 585
R427 B.n300 B.n299 585
R428 B.n301 B.n122 585
R429 B.n303 B.n302 585
R430 B.n304 B.n121 585
R431 B.n306 B.n305 585
R432 B.n307 B.n120 585
R433 B.n309 B.n308 585
R434 B.n310 B.n119 585
R435 B.n312 B.n311 585
R436 B.n313 B.n118 585
R437 B.n315 B.n314 585
R438 B.n316 B.n117 585
R439 B.n318 B.n317 585
R440 B.n319 B.n116 585
R441 B.n321 B.n320 585
R442 B.n322 B.n115 585
R443 B.n324 B.n323 585
R444 B.n325 B.n114 585
R445 B.n327 B.n326 585
R446 B.n328 B.n113 585
R447 B.n330 B.n329 585
R448 B.n331 B.n112 585
R449 B.n333 B.n332 585
R450 B.n334 B.n111 585
R451 B.n336 B.n335 585
R452 B.n337 B.n110 585
R453 B.n339 B.n338 585
R454 B.n340 B.n109 585
R455 B.n342 B.n341 585
R456 B.n234 B.n233 585
R457 B.n232 B.n149 585
R458 B.n231 B.n230 585
R459 B.n229 B.n150 585
R460 B.n228 B.n227 585
R461 B.n226 B.n151 585
R462 B.n225 B.n224 585
R463 B.n223 B.n152 585
R464 B.n222 B.n221 585
R465 B.n220 B.n153 585
R466 B.n219 B.n218 585
R467 B.n217 B.n154 585
R468 B.n216 B.n215 585
R469 B.n214 B.n155 585
R470 B.n213 B.n212 585
R471 B.n211 B.n156 585
R472 B.n210 B.n209 585
R473 B.n208 B.n157 585
R474 B.n207 B.n206 585
R475 B.n205 B.n158 585
R476 B.n204 B.n203 585
R477 B.n202 B.n159 585
R478 B.n201 B.n200 585
R479 B.n199 B.n160 585
R480 B.n198 B.n197 585
R481 B.n196 B.n161 585
R482 B.n195 B.n194 585
R483 B.n193 B.n162 585
R484 B.n192 B.n191 585
R485 B.n190 B.n163 585
R486 B.n189 B.n188 585
R487 B.n187 B.n164 585
R488 B.n186 B.n185 585
R489 B.n184 B.n165 585
R490 B.n183 B.n182 585
R491 B.n181 B.n166 585
R492 B.n180 B.n179 585
R493 B.n178 B.n167 585
R494 B.n177 B.n176 585
R495 B.n175 B.n168 585
R496 B.n174 B.n173 585
R497 B.n172 B.n169 585
R498 B.n171 B.n170 585
R499 B.n2 B.n0 585
R500 B.n649 B.n1 585
R501 B.n648 B.n647 585
R502 B.n646 B.n3 585
R503 B.n645 B.n644 585
R504 B.n643 B.n4 585
R505 B.n642 B.n641 585
R506 B.n640 B.n5 585
R507 B.n639 B.n638 585
R508 B.n637 B.n6 585
R509 B.n636 B.n635 585
R510 B.n634 B.n7 585
R511 B.n633 B.n632 585
R512 B.n631 B.n8 585
R513 B.n630 B.n629 585
R514 B.n628 B.n9 585
R515 B.n627 B.n626 585
R516 B.n625 B.n10 585
R517 B.n624 B.n623 585
R518 B.n622 B.n11 585
R519 B.n621 B.n620 585
R520 B.n619 B.n12 585
R521 B.n618 B.n617 585
R522 B.n616 B.n13 585
R523 B.n615 B.n614 585
R524 B.n613 B.n14 585
R525 B.n612 B.n611 585
R526 B.n610 B.n15 585
R527 B.n609 B.n608 585
R528 B.n607 B.n16 585
R529 B.n606 B.n605 585
R530 B.n604 B.n17 585
R531 B.n603 B.n602 585
R532 B.n601 B.n18 585
R533 B.n600 B.n599 585
R534 B.n598 B.n19 585
R535 B.n597 B.n596 585
R536 B.n595 B.n20 585
R537 B.n594 B.n593 585
R538 B.n592 B.n21 585
R539 B.n591 B.n590 585
R540 B.n589 B.n22 585
R541 B.n588 B.n587 585
R542 B.n586 B.n23 585
R543 B.n585 B.n584 585
R544 B.n651 B.n650 585
R545 B.n235 B.n234 521.33
R546 B.n584 B.n583 521.33
R547 B.n343 B.n342 521.33
R548 B.n476 B.n475 521.33
R549 B.n124 B.t6 302.423
R550 B.n132 B.t9 302.423
R551 B.n40 B.t0 302.423
R552 B.n46 B.t3 302.423
R553 B.n234 B.n149 163.367
R554 B.n230 B.n149 163.367
R555 B.n230 B.n229 163.367
R556 B.n229 B.n228 163.367
R557 B.n228 B.n151 163.367
R558 B.n224 B.n151 163.367
R559 B.n224 B.n223 163.367
R560 B.n223 B.n222 163.367
R561 B.n222 B.n153 163.367
R562 B.n218 B.n153 163.367
R563 B.n218 B.n217 163.367
R564 B.n217 B.n216 163.367
R565 B.n216 B.n155 163.367
R566 B.n212 B.n155 163.367
R567 B.n212 B.n211 163.367
R568 B.n211 B.n210 163.367
R569 B.n210 B.n157 163.367
R570 B.n206 B.n157 163.367
R571 B.n206 B.n205 163.367
R572 B.n205 B.n204 163.367
R573 B.n204 B.n159 163.367
R574 B.n200 B.n159 163.367
R575 B.n200 B.n199 163.367
R576 B.n199 B.n198 163.367
R577 B.n198 B.n161 163.367
R578 B.n194 B.n161 163.367
R579 B.n194 B.n193 163.367
R580 B.n193 B.n192 163.367
R581 B.n192 B.n163 163.367
R582 B.n188 B.n163 163.367
R583 B.n188 B.n187 163.367
R584 B.n187 B.n186 163.367
R585 B.n186 B.n165 163.367
R586 B.n182 B.n165 163.367
R587 B.n182 B.n181 163.367
R588 B.n181 B.n180 163.367
R589 B.n180 B.n167 163.367
R590 B.n176 B.n167 163.367
R591 B.n176 B.n175 163.367
R592 B.n175 B.n174 163.367
R593 B.n174 B.n169 163.367
R594 B.n170 B.n169 163.367
R595 B.n170 B.n2 163.367
R596 B.n650 B.n2 163.367
R597 B.n650 B.n649 163.367
R598 B.n649 B.n648 163.367
R599 B.n648 B.n3 163.367
R600 B.n644 B.n3 163.367
R601 B.n644 B.n643 163.367
R602 B.n643 B.n642 163.367
R603 B.n642 B.n5 163.367
R604 B.n638 B.n5 163.367
R605 B.n638 B.n637 163.367
R606 B.n637 B.n636 163.367
R607 B.n636 B.n7 163.367
R608 B.n632 B.n7 163.367
R609 B.n632 B.n631 163.367
R610 B.n631 B.n630 163.367
R611 B.n630 B.n9 163.367
R612 B.n626 B.n9 163.367
R613 B.n626 B.n625 163.367
R614 B.n625 B.n624 163.367
R615 B.n624 B.n11 163.367
R616 B.n620 B.n11 163.367
R617 B.n620 B.n619 163.367
R618 B.n619 B.n618 163.367
R619 B.n618 B.n13 163.367
R620 B.n614 B.n13 163.367
R621 B.n614 B.n613 163.367
R622 B.n613 B.n612 163.367
R623 B.n612 B.n15 163.367
R624 B.n608 B.n15 163.367
R625 B.n608 B.n607 163.367
R626 B.n607 B.n606 163.367
R627 B.n606 B.n17 163.367
R628 B.n602 B.n17 163.367
R629 B.n602 B.n601 163.367
R630 B.n601 B.n600 163.367
R631 B.n600 B.n19 163.367
R632 B.n596 B.n19 163.367
R633 B.n596 B.n595 163.367
R634 B.n595 B.n594 163.367
R635 B.n594 B.n21 163.367
R636 B.n590 B.n21 163.367
R637 B.n590 B.n589 163.367
R638 B.n589 B.n588 163.367
R639 B.n588 B.n23 163.367
R640 B.n584 B.n23 163.367
R641 B.n236 B.n235 163.367
R642 B.n236 B.n147 163.367
R643 B.n240 B.n147 163.367
R644 B.n241 B.n240 163.367
R645 B.n242 B.n241 163.367
R646 B.n242 B.n145 163.367
R647 B.n246 B.n145 163.367
R648 B.n247 B.n246 163.367
R649 B.n248 B.n247 163.367
R650 B.n248 B.n143 163.367
R651 B.n252 B.n143 163.367
R652 B.n253 B.n252 163.367
R653 B.n254 B.n253 163.367
R654 B.n254 B.n141 163.367
R655 B.n258 B.n141 163.367
R656 B.n259 B.n258 163.367
R657 B.n260 B.n259 163.367
R658 B.n260 B.n139 163.367
R659 B.n264 B.n139 163.367
R660 B.n265 B.n264 163.367
R661 B.n266 B.n265 163.367
R662 B.n266 B.n137 163.367
R663 B.n270 B.n137 163.367
R664 B.n271 B.n270 163.367
R665 B.n272 B.n271 163.367
R666 B.n272 B.n135 163.367
R667 B.n276 B.n135 163.367
R668 B.n277 B.n276 163.367
R669 B.n278 B.n277 163.367
R670 B.n278 B.n131 163.367
R671 B.n283 B.n131 163.367
R672 B.n284 B.n283 163.367
R673 B.n285 B.n284 163.367
R674 B.n285 B.n129 163.367
R675 B.n289 B.n129 163.367
R676 B.n290 B.n289 163.367
R677 B.n291 B.n290 163.367
R678 B.n291 B.n127 163.367
R679 B.n295 B.n127 163.367
R680 B.n296 B.n295 163.367
R681 B.n296 B.n123 163.367
R682 B.n300 B.n123 163.367
R683 B.n301 B.n300 163.367
R684 B.n302 B.n301 163.367
R685 B.n302 B.n121 163.367
R686 B.n306 B.n121 163.367
R687 B.n307 B.n306 163.367
R688 B.n308 B.n307 163.367
R689 B.n308 B.n119 163.367
R690 B.n312 B.n119 163.367
R691 B.n313 B.n312 163.367
R692 B.n314 B.n313 163.367
R693 B.n314 B.n117 163.367
R694 B.n318 B.n117 163.367
R695 B.n319 B.n318 163.367
R696 B.n320 B.n319 163.367
R697 B.n320 B.n115 163.367
R698 B.n324 B.n115 163.367
R699 B.n325 B.n324 163.367
R700 B.n326 B.n325 163.367
R701 B.n326 B.n113 163.367
R702 B.n330 B.n113 163.367
R703 B.n331 B.n330 163.367
R704 B.n332 B.n331 163.367
R705 B.n332 B.n111 163.367
R706 B.n336 B.n111 163.367
R707 B.n337 B.n336 163.367
R708 B.n338 B.n337 163.367
R709 B.n338 B.n109 163.367
R710 B.n342 B.n109 163.367
R711 B.n344 B.n343 163.367
R712 B.n344 B.n107 163.367
R713 B.n348 B.n107 163.367
R714 B.n349 B.n348 163.367
R715 B.n350 B.n349 163.367
R716 B.n350 B.n105 163.367
R717 B.n354 B.n105 163.367
R718 B.n355 B.n354 163.367
R719 B.n356 B.n355 163.367
R720 B.n356 B.n103 163.367
R721 B.n360 B.n103 163.367
R722 B.n361 B.n360 163.367
R723 B.n362 B.n361 163.367
R724 B.n362 B.n101 163.367
R725 B.n366 B.n101 163.367
R726 B.n367 B.n366 163.367
R727 B.n368 B.n367 163.367
R728 B.n368 B.n99 163.367
R729 B.n372 B.n99 163.367
R730 B.n373 B.n372 163.367
R731 B.n374 B.n373 163.367
R732 B.n374 B.n97 163.367
R733 B.n378 B.n97 163.367
R734 B.n379 B.n378 163.367
R735 B.n380 B.n379 163.367
R736 B.n380 B.n95 163.367
R737 B.n384 B.n95 163.367
R738 B.n385 B.n384 163.367
R739 B.n386 B.n385 163.367
R740 B.n386 B.n93 163.367
R741 B.n390 B.n93 163.367
R742 B.n391 B.n390 163.367
R743 B.n392 B.n391 163.367
R744 B.n392 B.n91 163.367
R745 B.n396 B.n91 163.367
R746 B.n397 B.n396 163.367
R747 B.n398 B.n397 163.367
R748 B.n398 B.n89 163.367
R749 B.n402 B.n89 163.367
R750 B.n403 B.n402 163.367
R751 B.n404 B.n403 163.367
R752 B.n404 B.n87 163.367
R753 B.n408 B.n87 163.367
R754 B.n409 B.n408 163.367
R755 B.n410 B.n409 163.367
R756 B.n410 B.n85 163.367
R757 B.n414 B.n85 163.367
R758 B.n415 B.n414 163.367
R759 B.n416 B.n415 163.367
R760 B.n416 B.n83 163.367
R761 B.n420 B.n83 163.367
R762 B.n421 B.n420 163.367
R763 B.n422 B.n421 163.367
R764 B.n422 B.n81 163.367
R765 B.n426 B.n81 163.367
R766 B.n427 B.n426 163.367
R767 B.n428 B.n427 163.367
R768 B.n428 B.n79 163.367
R769 B.n432 B.n79 163.367
R770 B.n433 B.n432 163.367
R771 B.n434 B.n433 163.367
R772 B.n434 B.n77 163.367
R773 B.n438 B.n77 163.367
R774 B.n439 B.n438 163.367
R775 B.n440 B.n439 163.367
R776 B.n440 B.n75 163.367
R777 B.n444 B.n75 163.367
R778 B.n445 B.n444 163.367
R779 B.n446 B.n445 163.367
R780 B.n446 B.n73 163.367
R781 B.n450 B.n73 163.367
R782 B.n451 B.n450 163.367
R783 B.n452 B.n451 163.367
R784 B.n452 B.n71 163.367
R785 B.n456 B.n71 163.367
R786 B.n457 B.n456 163.367
R787 B.n458 B.n457 163.367
R788 B.n458 B.n69 163.367
R789 B.n462 B.n69 163.367
R790 B.n463 B.n462 163.367
R791 B.n464 B.n463 163.367
R792 B.n464 B.n67 163.367
R793 B.n468 B.n67 163.367
R794 B.n469 B.n468 163.367
R795 B.n470 B.n469 163.367
R796 B.n470 B.n65 163.367
R797 B.n474 B.n65 163.367
R798 B.n475 B.n474 163.367
R799 B.n583 B.n582 163.367
R800 B.n582 B.n25 163.367
R801 B.n578 B.n25 163.367
R802 B.n578 B.n577 163.367
R803 B.n577 B.n576 163.367
R804 B.n576 B.n27 163.367
R805 B.n572 B.n27 163.367
R806 B.n572 B.n571 163.367
R807 B.n571 B.n570 163.367
R808 B.n570 B.n29 163.367
R809 B.n566 B.n29 163.367
R810 B.n566 B.n565 163.367
R811 B.n565 B.n564 163.367
R812 B.n564 B.n31 163.367
R813 B.n560 B.n31 163.367
R814 B.n560 B.n559 163.367
R815 B.n559 B.n558 163.367
R816 B.n558 B.n33 163.367
R817 B.n554 B.n33 163.367
R818 B.n554 B.n553 163.367
R819 B.n553 B.n552 163.367
R820 B.n552 B.n35 163.367
R821 B.n548 B.n35 163.367
R822 B.n548 B.n547 163.367
R823 B.n547 B.n546 163.367
R824 B.n546 B.n37 163.367
R825 B.n542 B.n37 163.367
R826 B.n542 B.n541 163.367
R827 B.n541 B.n540 163.367
R828 B.n540 B.n39 163.367
R829 B.n535 B.n39 163.367
R830 B.n535 B.n534 163.367
R831 B.n534 B.n533 163.367
R832 B.n533 B.n43 163.367
R833 B.n529 B.n43 163.367
R834 B.n529 B.n528 163.367
R835 B.n528 B.n527 163.367
R836 B.n527 B.n45 163.367
R837 B.n523 B.n45 163.367
R838 B.n523 B.n522 163.367
R839 B.n522 B.n49 163.367
R840 B.n518 B.n49 163.367
R841 B.n518 B.n517 163.367
R842 B.n517 B.n516 163.367
R843 B.n516 B.n51 163.367
R844 B.n512 B.n51 163.367
R845 B.n512 B.n511 163.367
R846 B.n511 B.n510 163.367
R847 B.n510 B.n53 163.367
R848 B.n506 B.n53 163.367
R849 B.n506 B.n505 163.367
R850 B.n505 B.n504 163.367
R851 B.n504 B.n55 163.367
R852 B.n500 B.n55 163.367
R853 B.n500 B.n499 163.367
R854 B.n499 B.n498 163.367
R855 B.n498 B.n57 163.367
R856 B.n494 B.n57 163.367
R857 B.n494 B.n493 163.367
R858 B.n493 B.n492 163.367
R859 B.n492 B.n59 163.367
R860 B.n488 B.n59 163.367
R861 B.n488 B.n487 163.367
R862 B.n487 B.n486 163.367
R863 B.n486 B.n61 163.367
R864 B.n482 B.n61 163.367
R865 B.n482 B.n481 163.367
R866 B.n481 B.n480 163.367
R867 B.n480 B.n63 163.367
R868 B.n476 B.n63 163.367
R869 B.n124 B.t8 159.272
R870 B.n46 B.t4 159.272
R871 B.n132 B.t11 159.262
R872 B.n40 B.t1 159.262
R873 B.n125 B.t7 111.951
R874 B.n47 B.t5 111.951
R875 B.n133 B.t10 111.941
R876 B.n41 B.t2 111.941
R877 B.n126 B.n125 59.5399
R878 B.n281 B.n133 59.5399
R879 B.n537 B.n41 59.5399
R880 B.n48 B.n47 59.5399
R881 B.n125 B.n124 47.3217
R882 B.n133 B.n132 47.3217
R883 B.n41 B.n40 47.3217
R884 B.n47 B.n46 47.3217
R885 B.n585 B.n24 33.8737
R886 B.n477 B.n64 33.8737
R887 B.n341 B.n108 33.8737
R888 B.n233 B.n148 33.8737
R889 B B.n651 18.0485
R890 B.n581 B.n24 10.6151
R891 B.n581 B.n580 10.6151
R892 B.n580 B.n579 10.6151
R893 B.n579 B.n26 10.6151
R894 B.n575 B.n26 10.6151
R895 B.n575 B.n574 10.6151
R896 B.n574 B.n573 10.6151
R897 B.n573 B.n28 10.6151
R898 B.n569 B.n28 10.6151
R899 B.n569 B.n568 10.6151
R900 B.n568 B.n567 10.6151
R901 B.n567 B.n30 10.6151
R902 B.n563 B.n30 10.6151
R903 B.n563 B.n562 10.6151
R904 B.n562 B.n561 10.6151
R905 B.n561 B.n32 10.6151
R906 B.n557 B.n32 10.6151
R907 B.n557 B.n556 10.6151
R908 B.n556 B.n555 10.6151
R909 B.n555 B.n34 10.6151
R910 B.n551 B.n34 10.6151
R911 B.n551 B.n550 10.6151
R912 B.n550 B.n549 10.6151
R913 B.n549 B.n36 10.6151
R914 B.n545 B.n36 10.6151
R915 B.n545 B.n544 10.6151
R916 B.n544 B.n543 10.6151
R917 B.n543 B.n38 10.6151
R918 B.n539 B.n38 10.6151
R919 B.n539 B.n538 10.6151
R920 B.n536 B.n42 10.6151
R921 B.n532 B.n42 10.6151
R922 B.n532 B.n531 10.6151
R923 B.n531 B.n530 10.6151
R924 B.n530 B.n44 10.6151
R925 B.n526 B.n44 10.6151
R926 B.n526 B.n525 10.6151
R927 B.n525 B.n524 10.6151
R928 B.n521 B.n520 10.6151
R929 B.n520 B.n519 10.6151
R930 B.n519 B.n50 10.6151
R931 B.n515 B.n50 10.6151
R932 B.n515 B.n514 10.6151
R933 B.n514 B.n513 10.6151
R934 B.n513 B.n52 10.6151
R935 B.n509 B.n52 10.6151
R936 B.n509 B.n508 10.6151
R937 B.n508 B.n507 10.6151
R938 B.n507 B.n54 10.6151
R939 B.n503 B.n54 10.6151
R940 B.n503 B.n502 10.6151
R941 B.n502 B.n501 10.6151
R942 B.n501 B.n56 10.6151
R943 B.n497 B.n56 10.6151
R944 B.n497 B.n496 10.6151
R945 B.n496 B.n495 10.6151
R946 B.n495 B.n58 10.6151
R947 B.n491 B.n58 10.6151
R948 B.n491 B.n490 10.6151
R949 B.n490 B.n489 10.6151
R950 B.n489 B.n60 10.6151
R951 B.n485 B.n60 10.6151
R952 B.n485 B.n484 10.6151
R953 B.n484 B.n483 10.6151
R954 B.n483 B.n62 10.6151
R955 B.n479 B.n62 10.6151
R956 B.n479 B.n478 10.6151
R957 B.n478 B.n477 10.6151
R958 B.n345 B.n108 10.6151
R959 B.n346 B.n345 10.6151
R960 B.n347 B.n346 10.6151
R961 B.n347 B.n106 10.6151
R962 B.n351 B.n106 10.6151
R963 B.n352 B.n351 10.6151
R964 B.n353 B.n352 10.6151
R965 B.n353 B.n104 10.6151
R966 B.n357 B.n104 10.6151
R967 B.n358 B.n357 10.6151
R968 B.n359 B.n358 10.6151
R969 B.n359 B.n102 10.6151
R970 B.n363 B.n102 10.6151
R971 B.n364 B.n363 10.6151
R972 B.n365 B.n364 10.6151
R973 B.n365 B.n100 10.6151
R974 B.n369 B.n100 10.6151
R975 B.n370 B.n369 10.6151
R976 B.n371 B.n370 10.6151
R977 B.n371 B.n98 10.6151
R978 B.n375 B.n98 10.6151
R979 B.n376 B.n375 10.6151
R980 B.n377 B.n376 10.6151
R981 B.n377 B.n96 10.6151
R982 B.n381 B.n96 10.6151
R983 B.n382 B.n381 10.6151
R984 B.n383 B.n382 10.6151
R985 B.n383 B.n94 10.6151
R986 B.n387 B.n94 10.6151
R987 B.n388 B.n387 10.6151
R988 B.n389 B.n388 10.6151
R989 B.n389 B.n92 10.6151
R990 B.n393 B.n92 10.6151
R991 B.n394 B.n393 10.6151
R992 B.n395 B.n394 10.6151
R993 B.n395 B.n90 10.6151
R994 B.n399 B.n90 10.6151
R995 B.n400 B.n399 10.6151
R996 B.n401 B.n400 10.6151
R997 B.n401 B.n88 10.6151
R998 B.n405 B.n88 10.6151
R999 B.n406 B.n405 10.6151
R1000 B.n407 B.n406 10.6151
R1001 B.n407 B.n86 10.6151
R1002 B.n411 B.n86 10.6151
R1003 B.n412 B.n411 10.6151
R1004 B.n413 B.n412 10.6151
R1005 B.n413 B.n84 10.6151
R1006 B.n417 B.n84 10.6151
R1007 B.n418 B.n417 10.6151
R1008 B.n419 B.n418 10.6151
R1009 B.n419 B.n82 10.6151
R1010 B.n423 B.n82 10.6151
R1011 B.n424 B.n423 10.6151
R1012 B.n425 B.n424 10.6151
R1013 B.n425 B.n80 10.6151
R1014 B.n429 B.n80 10.6151
R1015 B.n430 B.n429 10.6151
R1016 B.n431 B.n430 10.6151
R1017 B.n431 B.n78 10.6151
R1018 B.n435 B.n78 10.6151
R1019 B.n436 B.n435 10.6151
R1020 B.n437 B.n436 10.6151
R1021 B.n437 B.n76 10.6151
R1022 B.n441 B.n76 10.6151
R1023 B.n442 B.n441 10.6151
R1024 B.n443 B.n442 10.6151
R1025 B.n443 B.n74 10.6151
R1026 B.n447 B.n74 10.6151
R1027 B.n448 B.n447 10.6151
R1028 B.n449 B.n448 10.6151
R1029 B.n449 B.n72 10.6151
R1030 B.n453 B.n72 10.6151
R1031 B.n454 B.n453 10.6151
R1032 B.n455 B.n454 10.6151
R1033 B.n455 B.n70 10.6151
R1034 B.n459 B.n70 10.6151
R1035 B.n460 B.n459 10.6151
R1036 B.n461 B.n460 10.6151
R1037 B.n461 B.n68 10.6151
R1038 B.n465 B.n68 10.6151
R1039 B.n466 B.n465 10.6151
R1040 B.n467 B.n466 10.6151
R1041 B.n467 B.n66 10.6151
R1042 B.n471 B.n66 10.6151
R1043 B.n472 B.n471 10.6151
R1044 B.n473 B.n472 10.6151
R1045 B.n473 B.n64 10.6151
R1046 B.n237 B.n148 10.6151
R1047 B.n238 B.n237 10.6151
R1048 B.n239 B.n238 10.6151
R1049 B.n239 B.n146 10.6151
R1050 B.n243 B.n146 10.6151
R1051 B.n244 B.n243 10.6151
R1052 B.n245 B.n244 10.6151
R1053 B.n245 B.n144 10.6151
R1054 B.n249 B.n144 10.6151
R1055 B.n250 B.n249 10.6151
R1056 B.n251 B.n250 10.6151
R1057 B.n251 B.n142 10.6151
R1058 B.n255 B.n142 10.6151
R1059 B.n256 B.n255 10.6151
R1060 B.n257 B.n256 10.6151
R1061 B.n257 B.n140 10.6151
R1062 B.n261 B.n140 10.6151
R1063 B.n262 B.n261 10.6151
R1064 B.n263 B.n262 10.6151
R1065 B.n263 B.n138 10.6151
R1066 B.n267 B.n138 10.6151
R1067 B.n268 B.n267 10.6151
R1068 B.n269 B.n268 10.6151
R1069 B.n269 B.n136 10.6151
R1070 B.n273 B.n136 10.6151
R1071 B.n274 B.n273 10.6151
R1072 B.n275 B.n274 10.6151
R1073 B.n275 B.n134 10.6151
R1074 B.n279 B.n134 10.6151
R1075 B.n280 B.n279 10.6151
R1076 B.n282 B.n130 10.6151
R1077 B.n286 B.n130 10.6151
R1078 B.n287 B.n286 10.6151
R1079 B.n288 B.n287 10.6151
R1080 B.n288 B.n128 10.6151
R1081 B.n292 B.n128 10.6151
R1082 B.n293 B.n292 10.6151
R1083 B.n294 B.n293 10.6151
R1084 B.n298 B.n297 10.6151
R1085 B.n299 B.n298 10.6151
R1086 B.n299 B.n122 10.6151
R1087 B.n303 B.n122 10.6151
R1088 B.n304 B.n303 10.6151
R1089 B.n305 B.n304 10.6151
R1090 B.n305 B.n120 10.6151
R1091 B.n309 B.n120 10.6151
R1092 B.n310 B.n309 10.6151
R1093 B.n311 B.n310 10.6151
R1094 B.n311 B.n118 10.6151
R1095 B.n315 B.n118 10.6151
R1096 B.n316 B.n315 10.6151
R1097 B.n317 B.n316 10.6151
R1098 B.n317 B.n116 10.6151
R1099 B.n321 B.n116 10.6151
R1100 B.n322 B.n321 10.6151
R1101 B.n323 B.n322 10.6151
R1102 B.n323 B.n114 10.6151
R1103 B.n327 B.n114 10.6151
R1104 B.n328 B.n327 10.6151
R1105 B.n329 B.n328 10.6151
R1106 B.n329 B.n112 10.6151
R1107 B.n333 B.n112 10.6151
R1108 B.n334 B.n333 10.6151
R1109 B.n335 B.n334 10.6151
R1110 B.n335 B.n110 10.6151
R1111 B.n339 B.n110 10.6151
R1112 B.n340 B.n339 10.6151
R1113 B.n341 B.n340 10.6151
R1114 B.n233 B.n232 10.6151
R1115 B.n232 B.n231 10.6151
R1116 B.n231 B.n150 10.6151
R1117 B.n227 B.n150 10.6151
R1118 B.n227 B.n226 10.6151
R1119 B.n226 B.n225 10.6151
R1120 B.n225 B.n152 10.6151
R1121 B.n221 B.n152 10.6151
R1122 B.n221 B.n220 10.6151
R1123 B.n220 B.n219 10.6151
R1124 B.n219 B.n154 10.6151
R1125 B.n215 B.n154 10.6151
R1126 B.n215 B.n214 10.6151
R1127 B.n214 B.n213 10.6151
R1128 B.n213 B.n156 10.6151
R1129 B.n209 B.n156 10.6151
R1130 B.n209 B.n208 10.6151
R1131 B.n208 B.n207 10.6151
R1132 B.n207 B.n158 10.6151
R1133 B.n203 B.n158 10.6151
R1134 B.n203 B.n202 10.6151
R1135 B.n202 B.n201 10.6151
R1136 B.n201 B.n160 10.6151
R1137 B.n197 B.n160 10.6151
R1138 B.n197 B.n196 10.6151
R1139 B.n196 B.n195 10.6151
R1140 B.n195 B.n162 10.6151
R1141 B.n191 B.n162 10.6151
R1142 B.n191 B.n190 10.6151
R1143 B.n190 B.n189 10.6151
R1144 B.n189 B.n164 10.6151
R1145 B.n185 B.n164 10.6151
R1146 B.n185 B.n184 10.6151
R1147 B.n184 B.n183 10.6151
R1148 B.n183 B.n166 10.6151
R1149 B.n179 B.n166 10.6151
R1150 B.n179 B.n178 10.6151
R1151 B.n178 B.n177 10.6151
R1152 B.n177 B.n168 10.6151
R1153 B.n173 B.n168 10.6151
R1154 B.n173 B.n172 10.6151
R1155 B.n172 B.n171 10.6151
R1156 B.n171 B.n0 10.6151
R1157 B.n647 B.n1 10.6151
R1158 B.n647 B.n646 10.6151
R1159 B.n646 B.n645 10.6151
R1160 B.n645 B.n4 10.6151
R1161 B.n641 B.n4 10.6151
R1162 B.n641 B.n640 10.6151
R1163 B.n640 B.n639 10.6151
R1164 B.n639 B.n6 10.6151
R1165 B.n635 B.n6 10.6151
R1166 B.n635 B.n634 10.6151
R1167 B.n634 B.n633 10.6151
R1168 B.n633 B.n8 10.6151
R1169 B.n629 B.n8 10.6151
R1170 B.n629 B.n628 10.6151
R1171 B.n628 B.n627 10.6151
R1172 B.n627 B.n10 10.6151
R1173 B.n623 B.n10 10.6151
R1174 B.n623 B.n622 10.6151
R1175 B.n622 B.n621 10.6151
R1176 B.n621 B.n12 10.6151
R1177 B.n617 B.n12 10.6151
R1178 B.n617 B.n616 10.6151
R1179 B.n616 B.n615 10.6151
R1180 B.n615 B.n14 10.6151
R1181 B.n611 B.n14 10.6151
R1182 B.n611 B.n610 10.6151
R1183 B.n610 B.n609 10.6151
R1184 B.n609 B.n16 10.6151
R1185 B.n605 B.n16 10.6151
R1186 B.n605 B.n604 10.6151
R1187 B.n604 B.n603 10.6151
R1188 B.n603 B.n18 10.6151
R1189 B.n599 B.n18 10.6151
R1190 B.n599 B.n598 10.6151
R1191 B.n598 B.n597 10.6151
R1192 B.n597 B.n20 10.6151
R1193 B.n593 B.n20 10.6151
R1194 B.n593 B.n592 10.6151
R1195 B.n592 B.n591 10.6151
R1196 B.n591 B.n22 10.6151
R1197 B.n587 B.n22 10.6151
R1198 B.n587 B.n586 10.6151
R1199 B.n586 B.n585 10.6151
R1200 B.n537 B.n536 6.5566
R1201 B.n524 B.n48 6.5566
R1202 B.n282 B.n281 6.5566
R1203 B.n294 B.n126 6.5566
R1204 B.n538 B.n537 4.05904
R1205 B.n521 B.n48 4.05904
R1206 B.n281 B.n280 4.05904
R1207 B.n297 B.n126 4.05904
R1208 B.n651 B.n0 2.81026
R1209 B.n651 B.n1 2.81026
C0 VN B 1.07163f
C1 w_n3410_n2636# VDD1 1.69913f
C2 VDD1 VTAIL 6.69112f
C3 VN VDD2 5.9024f
C4 B VDD1 1.40236f
C5 VP w_n3410_n2636# 7.16234f
C6 VP VTAIL 6.31177f
C7 VDD1 VDD2 1.52302f
C8 VN VDD1 0.151264f
C9 w_n3410_n2636# VTAIL 3.3448f
C10 VP B 1.8087f
C11 VP VDD2 0.467951f
C12 B w_n3410_n2636# 8.339139f
C13 B VTAIL 3.58329f
C14 VP VN 6.38013f
C15 w_n3410_n2636# VDD2 1.79329f
C16 VDD2 VTAIL 6.74225f
C17 VN w_n3410_n2636# 6.72109f
C18 VN VTAIL 6.29766f
C19 B VDD2 1.48297f
C20 VP VDD1 6.21794f
C21 VDD2 VSUBS 1.529712f
C22 VDD1 VSUBS 2.096008f
C23 VTAIL VSUBS 1.083936f
C24 VN VSUBS 6.00413f
C25 VP VSUBS 2.95872f
C26 B VSUBS 4.14419f
C27 w_n3410_n2636# VSUBS 0.111425p
C28 B.n0 VSUBS 0.004821f
C29 B.n1 VSUBS 0.004821f
C30 B.n2 VSUBS 0.007624f
C31 B.n3 VSUBS 0.007624f
C32 B.n4 VSUBS 0.007624f
C33 B.n5 VSUBS 0.007624f
C34 B.n6 VSUBS 0.007624f
C35 B.n7 VSUBS 0.007624f
C36 B.n8 VSUBS 0.007624f
C37 B.n9 VSUBS 0.007624f
C38 B.n10 VSUBS 0.007624f
C39 B.n11 VSUBS 0.007624f
C40 B.n12 VSUBS 0.007624f
C41 B.n13 VSUBS 0.007624f
C42 B.n14 VSUBS 0.007624f
C43 B.n15 VSUBS 0.007624f
C44 B.n16 VSUBS 0.007624f
C45 B.n17 VSUBS 0.007624f
C46 B.n18 VSUBS 0.007624f
C47 B.n19 VSUBS 0.007624f
C48 B.n20 VSUBS 0.007624f
C49 B.n21 VSUBS 0.007624f
C50 B.n22 VSUBS 0.007624f
C51 B.n23 VSUBS 0.007624f
C52 B.n24 VSUBS 0.018583f
C53 B.n25 VSUBS 0.007624f
C54 B.n26 VSUBS 0.007624f
C55 B.n27 VSUBS 0.007624f
C56 B.n28 VSUBS 0.007624f
C57 B.n29 VSUBS 0.007624f
C58 B.n30 VSUBS 0.007624f
C59 B.n31 VSUBS 0.007624f
C60 B.n32 VSUBS 0.007624f
C61 B.n33 VSUBS 0.007624f
C62 B.n34 VSUBS 0.007624f
C63 B.n35 VSUBS 0.007624f
C64 B.n36 VSUBS 0.007624f
C65 B.n37 VSUBS 0.007624f
C66 B.n38 VSUBS 0.007624f
C67 B.n39 VSUBS 0.007624f
C68 B.t2 VSUBS 0.282195f
C69 B.t1 VSUBS 0.301431f
C70 B.t0 VSUBS 0.880252f
C71 B.n40 VSUBS 0.155715f
C72 B.n41 VSUBS 0.075612f
C73 B.n42 VSUBS 0.007624f
C74 B.n43 VSUBS 0.007624f
C75 B.n44 VSUBS 0.007624f
C76 B.n45 VSUBS 0.007624f
C77 B.t5 VSUBS 0.282193f
C78 B.t4 VSUBS 0.301428f
C79 B.t3 VSUBS 0.880252f
C80 B.n46 VSUBS 0.155718f
C81 B.n47 VSUBS 0.075615f
C82 B.n48 VSUBS 0.017665f
C83 B.n49 VSUBS 0.007624f
C84 B.n50 VSUBS 0.007624f
C85 B.n51 VSUBS 0.007624f
C86 B.n52 VSUBS 0.007624f
C87 B.n53 VSUBS 0.007624f
C88 B.n54 VSUBS 0.007624f
C89 B.n55 VSUBS 0.007624f
C90 B.n56 VSUBS 0.007624f
C91 B.n57 VSUBS 0.007624f
C92 B.n58 VSUBS 0.007624f
C93 B.n59 VSUBS 0.007624f
C94 B.n60 VSUBS 0.007624f
C95 B.n61 VSUBS 0.007624f
C96 B.n62 VSUBS 0.007624f
C97 B.n63 VSUBS 0.007624f
C98 B.n64 VSUBS 0.018838f
C99 B.n65 VSUBS 0.007624f
C100 B.n66 VSUBS 0.007624f
C101 B.n67 VSUBS 0.007624f
C102 B.n68 VSUBS 0.007624f
C103 B.n69 VSUBS 0.007624f
C104 B.n70 VSUBS 0.007624f
C105 B.n71 VSUBS 0.007624f
C106 B.n72 VSUBS 0.007624f
C107 B.n73 VSUBS 0.007624f
C108 B.n74 VSUBS 0.007624f
C109 B.n75 VSUBS 0.007624f
C110 B.n76 VSUBS 0.007624f
C111 B.n77 VSUBS 0.007624f
C112 B.n78 VSUBS 0.007624f
C113 B.n79 VSUBS 0.007624f
C114 B.n80 VSUBS 0.007624f
C115 B.n81 VSUBS 0.007624f
C116 B.n82 VSUBS 0.007624f
C117 B.n83 VSUBS 0.007624f
C118 B.n84 VSUBS 0.007624f
C119 B.n85 VSUBS 0.007624f
C120 B.n86 VSUBS 0.007624f
C121 B.n87 VSUBS 0.007624f
C122 B.n88 VSUBS 0.007624f
C123 B.n89 VSUBS 0.007624f
C124 B.n90 VSUBS 0.007624f
C125 B.n91 VSUBS 0.007624f
C126 B.n92 VSUBS 0.007624f
C127 B.n93 VSUBS 0.007624f
C128 B.n94 VSUBS 0.007624f
C129 B.n95 VSUBS 0.007624f
C130 B.n96 VSUBS 0.007624f
C131 B.n97 VSUBS 0.007624f
C132 B.n98 VSUBS 0.007624f
C133 B.n99 VSUBS 0.007624f
C134 B.n100 VSUBS 0.007624f
C135 B.n101 VSUBS 0.007624f
C136 B.n102 VSUBS 0.007624f
C137 B.n103 VSUBS 0.007624f
C138 B.n104 VSUBS 0.007624f
C139 B.n105 VSUBS 0.007624f
C140 B.n106 VSUBS 0.007624f
C141 B.n107 VSUBS 0.007624f
C142 B.n108 VSUBS 0.017969f
C143 B.n109 VSUBS 0.007624f
C144 B.n110 VSUBS 0.007624f
C145 B.n111 VSUBS 0.007624f
C146 B.n112 VSUBS 0.007624f
C147 B.n113 VSUBS 0.007624f
C148 B.n114 VSUBS 0.007624f
C149 B.n115 VSUBS 0.007624f
C150 B.n116 VSUBS 0.007624f
C151 B.n117 VSUBS 0.007624f
C152 B.n118 VSUBS 0.007624f
C153 B.n119 VSUBS 0.007624f
C154 B.n120 VSUBS 0.007624f
C155 B.n121 VSUBS 0.007624f
C156 B.n122 VSUBS 0.007624f
C157 B.n123 VSUBS 0.007624f
C158 B.t7 VSUBS 0.282193f
C159 B.t8 VSUBS 0.301428f
C160 B.t6 VSUBS 0.880252f
C161 B.n124 VSUBS 0.155718f
C162 B.n125 VSUBS 0.075615f
C163 B.n126 VSUBS 0.017665f
C164 B.n127 VSUBS 0.007624f
C165 B.n128 VSUBS 0.007624f
C166 B.n129 VSUBS 0.007624f
C167 B.n130 VSUBS 0.007624f
C168 B.n131 VSUBS 0.007624f
C169 B.t10 VSUBS 0.282195f
C170 B.t11 VSUBS 0.301431f
C171 B.t9 VSUBS 0.880252f
C172 B.n132 VSUBS 0.155715f
C173 B.n133 VSUBS 0.075612f
C174 B.n134 VSUBS 0.007624f
C175 B.n135 VSUBS 0.007624f
C176 B.n136 VSUBS 0.007624f
C177 B.n137 VSUBS 0.007624f
C178 B.n138 VSUBS 0.007624f
C179 B.n139 VSUBS 0.007624f
C180 B.n140 VSUBS 0.007624f
C181 B.n141 VSUBS 0.007624f
C182 B.n142 VSUBS 0.007624f
C183 B.n143 VSUBS 0.007624f
C184 B.n144 VSUBS 0.007624f
C185 B.n145 VSUBS 0.007624f
C186 B.n146 VSUBS 0.007624f
C187 B.n147 VSUBS 0.007624f
C188 B.n148 VSUBS 0.018583f
C189 B.n149 VSUBS 0.007624f
C190 B.n150 VSUBS 0.007624f
C191 B.n151 VSUBS 0.007624f
C192 B.n152 VSUBS 0.007624f
C193 B.n153 VSUBS 0.007624f
C194 B.n154 VSUBS 0.007624f
C195 B.n155 VSUBS 0.007624f
C196 B.n156 VSUBS 0.007624f
C197 B.n157 VSUBS 0.007624f
C198 B.n158 VSUBS 0.007624f
C199 B.n159 VSUBS 0.007624f
C200 B.n160 VSUBS 0.007624f
C201 B.n161 VSUBS 0.007624f
C202 B.n162 VSUBS 0.007624f
C203 B.n163 VSUBS 0.007624f
C204 B.n164 VSUBS 0.007624f
C205 B.n165 VSUBS 0.007624f
C206 B.n166 VSUBS 0.007624f
C207 B.n167 VSUBS 0.007624f
C208 B.n168 VSUBS 0.007624f
C209 B.n169 VSUBS 0.007624f
C210 B.n170 VSUBS 0.007624f
C211 B.n171 VSUBS 0.007624f
C212 B.n172 VSUBS 0.007624f
C213 B.n173 VSUBS 0.007624f
C214 B.n174 VSUBS 0.007624f
C215 B.n175 VSUBS 0.007624f
C216 B.n176 VSUBS 0.007624f
C217 B.n177 VSUBS 0.007624f
C218 B.n178 VSUBS 0.007624f
C219 B.n179 VSUBS 0.007624f
C220 B.n180 VSUBS 0.007624f
C221 B.n181 VSUBS 0.007624f
C222 B.n182 VSUBS 0.007624f
C223 B.n183 VSUBS 0.007624f
C224 B.n184 VSUBS 0.007624f
C225 B.n185 VSUBS 0.007624f
C226 B.n186 VSUBS 0.007624f
C227 B.n187 VSUBS 0.007624f
C228 B.n188 VSUBS 0.007624f
C229 B.n189 VSUBS 0.007624f
C230 B.n190 VSUBS 0.007624f
C231 B.n191 VSUBS 0.007624f
C232 B.n192 VSUBS 0.007624f
C233 B.n193 VSUBS 0.007624f
C234 B.n194 VSUBS 0.007624f
C235 B.n195 VSUBS 0.007624f
C236 B.n196 VSUBS 0.007624f
C237 B.n197 VSUBS 0.007624f
C238 B.n198 VSUBS 0.007624f
C239 B.n199 VSUBS 0.007624f
C240 B.n200 VSUBS 0.007624f
C241 B.n201 VSUBS 0.007624f
C242 B.n202 VSUBS 0.007624f
C243 B.n203 VSUBS 0.007624f
C244 B.n204 VSUBS 0.007624f
C245 B.n205 VSUBS 0.007624f
C246 B.n206 VSUBS 0.007624f
C247 B.n207 VSUBS 0.007624f
C248 B.n208 VSUBS 0.007624f
C249 B.n209 VSUBS 0.007624f
C250 B.n210 VSUBS 0.007624f
C251 B.n211 VSUBS 0.007624f
C252 B.n212 VSUBS 0.007624f
C253 B.n213 VSUBS 0.007624f
C254 B.n214 VSUBS 0.007624f
C255 B.n215 VSUBS 0.007624f
C256 B.n216 VSUBS 0.007624f
C257 B.n217 VSUBS 0.007624f
C258 B.n218 VSUBS 0.007624f
C259 B.n219 VSUBS 0.007624f
C260 B.n220 VSUBS 0.007624f
C261 B.n221 VSUBS 0.007624f
C262 B.n222 VSUBS 0.007624f
C263 B.n223 VSUBS 0.007624f
C264 B.n224 VSUBS 0.007624f
C265 B.n225 VSUBS 0.007624f
C266 B.n226 VSUBS 0.007624f
C267 B.n227 VSUBS 0.007624f
C268 B.n228 VSUBS 0.007624f
C269 B.n229 VSUBS 0.007624f
C270 B.n230 VSUBS 0.007624f
C271 B.n231 VSUBS 0.007624f
C272 B.n232 VSUBS 0.007624f
C273 B.n233 VSUBS 0.017969f
C274 B.n234 VSUBS 0.017969f
C275 B.n235 VSUBS 0.018583f
C276 B.n236 VSUBS 0.007624f
C277 B.n237 VSUBS 0.007624f
C278 B.n238 VSUBS 0.007624f
C279 B.n239 VSUBS 0.007624f
C280 B.n240 VSUBS 0.007624f
C281 B.n241 VSUBS 0.007624f
C282 B.n242 VSUBS 0.007624f
C283 B.n243 VSUBS 0.007624f
C284 B.n244 VSUBS 0.007624f
C285 B.n245 VSUBS 0.007624f
C286 B.n246 VSUBS 0.007624f
C287 B.n247 VSUBS 0.007624f
C288 B.n248 VSUBS 0.007624f
C289 B.n249 VSUBS 0.007624f
C290 B.n250 VSUBS 0.007624f
C291 B.n251 VSUBS 0.007624f
C292 B.n252 VSUBS 0.007624f
C293 B.n253 VSUBS 0.007624f
C294 B.n254 VSUBS 0.007624f
C295 B.n255 VSUBS 0.007624f
C296 B.n256 VSUBS 0.007624f
C297 B.n257 VSUBS 0.007624f
C298 B.n258 VSUBS 0.007624f
C299 B.n259 VSUBS 0.007624f
C300 B.n260 VSUBS 0.007624f
C301 B.n261 VSUBS 0.007624f
C302 B.n262 VSUBS 0.007624f
C303 B.n263 VSUBS 0.007624f
C304 B.n264 VSUBS 0.007624f
C305 B.n265 VSUBS 0.007624f
C306 B.n266 VSUBS 0.007624f
C307 B.n267 VSUBS 0.007624f
C308 B.n268 VSUBS 0.007624f
C309 B.n269 VSUBS 0.007624f
C310 B.n270 VSUBS 0.007624f
C311 B.n271 VSUBS 0.007624f
C312 B.n272 VSUBS 0.007624f
C313 B.n273 VSUBS 0.007624f
C314 B.n274 VSUBS 0.007624f
C315 B.n275 VSUBS 0.007624f
C316 B.n276 VSUBS 0.007624f
C317 B.n277 VSUBS 0.007624f
C318 B.n278 VSUBS 0.007624f
C319 B.n279 VSUBS 0.007624f
C320 B.n280 VSUBS 0.00527f
C321 B.n281 VSUBS 0.017665f
C322 B.n282 VSUBS 0.006167f
C323 B.n283 VSUBS 0.007624f
C324 B.n284 VSUBS 0.007624f
C325 B.n285 VSUBS 0.007624f
C326 B.n286 VSUBS 0.007624f
C327 B.n287 VSUBS 0.007624f
C328 B.n288 VSUBS 0.007624f
C329 B.n289 VSUBS 0.007624f
C330 B.n290 VSUBS 0.007624f
C331 B.n291 VSUBS 0.007624f
C332 B.n292 VSUBS 0.007624f
C333 B.n293 VSUBS 0.007624f
C334 B.n294 VSUBS 0.006167f
C335 B.n295 VSUBS 0.007624f
C336 B.n296 VSUBS 0.007624f
C337 B.n297 VSUBS 0.00527f
C338 B.n298 VSUBS 0.007624f
C339 B.n299 VSUBS 0.007624f
C340 B.n300 VSUBS 0.007624f
C341 B.n301 VSUBS 0.007624f
C342 B.n302 VSUBS 0.007624f
C343 B.n303 VSUBS 0.007624f
C344 B.n304 VSUBS 0.007624f
C345 B.n305 VSUBS 0.007624f
C346 B.n306 VSUBS 0.007624f
C347 B.n307 VSUBS 0.007624f
C348 B.n308 VSUBS 0.007624f
C349 B.n309 VSUBS 0.007624f
C350 B.n310 VSUBS 0.007624f
C351 B.n311 VSUBS 0.007624f
C352 B.n312 VSUBS 0.007624f
C353 B.n313 VSUBS 0.007624f
C354 B.n314 VSUBS 0.007624f
C355 B.n315 VSUBS 0.007624f
C356 B.n316 VSUBS 0.007624f
C357 B.n317 VSUBS 0.007624f
C358 B.n318 VSUBS 0.007624f
C359 B.n319 VSUBS 0.007624f
C360 B.n320 VSUBS 0.007624f
C361 B.n321 VSUBS 0.007624f
C362 B.n322 VSUBS 0.007624f
C363 B.n323 VSUBS 0.007624f
C364 B.n324 VSUBS 0.007624f
C365 B.n325 VSUBS 0.007624f
C366 B.n326 VSUBS 0.007624f
C367 B.n327 VSUBS 0.007624f
C368 B.n328 VSUBS 0.007624f
C369 B.n329 VSUBS 0.007624f
C370 B.n330 VSUBS 0.007624f
C371 B.n331 VSUBS 0.007624f
C372 B.n332 VSUBS 0.007624f
C373 B.n333 VSUBS 0.007624f
C374 B.n334 VSUBS 0.007624f
C375 B.n335 VSUBS 0.007624f
C376 B.n336 VSUBS 0.007624f
C377 B.n337 VSUBS 0.007624f
C378 B.n338 VSUBS 0.007624f
C379 B.n339 VSUBS 0.007624f
C380 B.n340 VSUBS 0.007624f
C381 B.n341 VSUBS 0.018583f
C382 B.n342 VSUBS 0.018583f
C383 B.n343 VSUBS 0.017969f
C384 B.n344 VSUBS 0.007624f
C385 B.n345 VSUBS 0.007624f
C386 B.n346 VSUBS 0.007624f
C387 B.n347 VSUBS 0.007624f
C388 B.n348 VSUBS 0.007624f
C389 B.n349 VSUBS 0.007624f
C390 B.n350 VSUBS 0.007624f
C391 B.n351 VSUBS 0.007624f
C392 B.n352 VSUBS 0.007624f
C393 B.n353 VSUBS 0.007624f
C394 B.n354 VSUBS 0.007624f
C395 B.n355 VSUBS 0.007624f
C396 B.n356 VSUBS 0.007624f
C397 B.n357 VSUBS 0.007624f
C398 B.n358 VSUBS 0.007624f
C399 B.n359 VSUBS 0.007624f
C400 B.n360 VSUBS 0.007624f
C401 B.n361 VSUBS 0.007624f
C402 B.n362 VSUBS 0.007624f
C403 B.n363 VSUBS 0.007624f
C404 B.n364 VSUBS 0.007624f
C405 B.n365 VSUBS 0.007624f
C406 B.n366 VSUBS 0.007624f
C407 B.n367 VSUBS 0.007624f
C408 B.n368 VSUBS 0.007624f
C409 B.n369 VSUBS 0.007624f
C410 B.n370 VSUBS 0.007624f
C411 B.n371 VSUBS 0.007624f
C412 B.n372 VSUBS 0.007624f
C413 B.n373 VSUBS 0.007624f
C414 B.n374 VSUBS 0.007624f
C415 B.n375 VSUBS 0.007624f
C416 B.n376 VSUBS 0.007624f
C417 B.n377 VSUBS 0.007624f
C418 B.n378 VSUBS 0.007624f
C419 B.n379 VSUBS 0.007624f
C420 B.n380 VSUBS 0.007624f
C421 B.n381 VSUBS 0.007624f
C422 B.n382 VSUBS 0.007624f
C423 B.n383 VSUBS 0.007624f
C424 B.n384 VSUBS 0.007624f
C425 B.n385 VSUBS 0.007624f
C426 B.n386 VSUBS 0.007624f
C427 B.n387 VSUBS 0.007624f
C428 B.n388 VSUBS 0.007624f
C429 B.n389 VSUBS 0.007624f
C430 B.n390 VSUBS 0.007624f
C431 B.n391 VSUBS 0.007624f
C432 B.n392 VSUBS 0.007624f
C433 B.n393 VSUBS 0.007624f
C434 B.n394 VSUBS 0.007624f
C435 B.n395 VSUBS 0.007624f
C436 B.n396 VSUBS 0.007624f
C437 B.n397 VSUBS 0.007624f
C438 B.n398 VSUBS 0.007624f
C439 B.n399 VSUBS 0.007624f
C440 B.n400 VSUBS 0.007624f
C441 B.n401 VSUBS 0.007624f
C442 B.n402 VSUBS 0.007624f
C443 B.n403 VSUBS 0.007624f
C444 B.n404 VSUBS 0.007624f
C445 B.n405 VSUBS 0.007624f
C446 B.n406 VSUBS 0.007624f
C447 B.n407 VSUBS 0.007624f
C448 B.n408 VSUBS 0.007624f
C449 B.n409 VSUBS 0.007624f
C450 B.n410 VSUBS 0.007624f
C451 B.n411 VSUBS 0.007624f
C452 B.n412 VSUBS 0.007624f
C453 B.n413 VSUBS 0.007624f
C454 B.n414 VSUBS 0.007624f
C455 B.n415 VSUBS 0.007624f
C456 B.n416 VSUBS 0.007624f
C457 B.n417 VSUBS 0.007624f
C458 B.n418 VSUBS 0.007624f
C459 B.n419 VSUBS 0.007624f
C460 B.n420 VSUBS 0.007624f
C461 B.n421 VSUBS 0.007624f
C462 B.n422 VSUBS 0.007624f
C463 B.n423 VSUBS 0.007624f
C464 B.n424 VSUBS 0.007624f
C465 B.n425 VSUBS 0.007624f
C466 B.n426 VSUBS 0.007624f
C467 B.n427 VSUBS 0.007624f
C468 B.n428 VSUBS 0.007624f
C469 B.n429 VSUBS 0.007624f
C470 B.n430 VSUBS 0.007624f
C471 B.n431 VSUBS 0.007624f
C472 B.n432 VSUBS 0.007624f
C473 B.n433 VSUBS 0.007624f
C474 B.n434 VSUBS 0.007624f
C475 B.n435 VSUBS 0.007624f
C476 B.n436 VSUBS 0.007624f
C477 B.n437 VSUBS 0.007624f
C478 B.n438 VSUBS 0.007624f
C479 B.n439 VSUBS 0.007624f
C480 B.n440 VSUBS 0.007624f
C481 B.n441 VSUBS 0.007624f
C482 B.n442 VSUBS 0.007624f
C483 B.n443 VSUBS 0.007624f
C484 B.n444 VSUBS 0.007624f
C485 B.n445 VSUBS 0.007624f
C486 B.n446 VSUBS 0.007624f
C487 B.n447 VSUBS 0.007624f
C488 B.n448 VSUBS 0.007624f
C489 B.n449 VSUBS 0.007624f
C490 B.n450 VSUBS 0.007624f
C491 B.n451 VSUBS 0.007624f
C492 B.n452 VSUBS 0.007624f
C493 B.n453 VSUBS 0.007624f
C494 B.n454 VSUBS 0.007624f
C495 B.n455 VSUBS 0.007624f
C496 B.n456 VSUBS 0.007624f
C497 B.n457 VSUBS 0.007624f
C498 B.n458 VSUBS 0.007624f
C499 B.n459 VSUBS 0.007624f
C500 B.n460 VSUBS 0.007624f
C501 B.n461 VSUBS 0.007624f
C502 B.n462 VSUBS 0.007624f
C503 B.n463 VSUBS 0.007624f
C504 B.n464 VSUBS 0.007624f
C505 B.n465 VSUBS 0.007624f
C506 B.n466 VSUBS 0.007624f
C507 B.n467 VSUBS 0.007624f
C508 B.n468 VSUBS 0.007624f
C509 B.n469 VSUBS 0.007624f
C510 B.n470 VSUBS 0.007624f
C511 B.n471 VSUBS 0.007624f
C512 B.n472 VSUBS 0.007624f
C513 B.n473 VSUBS 0.007624f
C514 B.n474 VSUBS 0.007624f
C515 B.n475 VSUBS 0.017969f
C516 B.n476 VSUBS 0.018583f
C517 B.n477 VSUBS 0.017715f
C518 B.n478 VSUBS 0.007624f
C519 B.n479 VSUBS 0.007624f
C520 B.n480 VSUBS 0.007624f
C521 B.n481 VSUBS 0.007624f
C522 B.n482 VSUBS 0.007624f
C523 B.n483 VSUBS 0.007624f
C524 B.n484 VSUBS 0.007624f
C525 B.n485 VSUBS 0.007624f
C526 B.n486 VSUBS 0.007624f
C527 B.n487 VSUBS 0.007624f
C528 B.n488 VSUBS 0.007624f
C529 B.n489 VSUBS 0.007624f
C530 B.n490 VSUBS 0.007624f
C531 B.n491 VSUBS 0.007624f
C532 B.n492 VSUBS 0.007624f
C533 B.n493 VSUBS 0.007624f
C534 B.n494 VSUBS 0.007624f
C535 B.n495 VSUBS 0.007624f
C536 B.n496 VSUBS 0.007624f
C537 B.n497 VSUBS 0.007624f
C538 B.n498 VSUBS 0.007624f
C539 B.n499 VSUBS 0.007624f
C540 B.n500 VSUBS 0.007624f
C541 B.n501 VSUBS 0.007624f
C542 B.n502 VSUBS 0.007624f
C543 B.n503 VSUBS 0.007624f
C544 B.n504 VSUBS 0.007624f
C545 B.n505 VSUBS 0.007624f
C546 B.n506 VSUBS 0.007624f
C547 B.n507 VSUBS 0.007624f
C548 B.n508 VSUBS 0.007624f
C549 B.n509 VSUBS 0.007624f
C550 B.n510 VSUBS 0.007624f
C551 B.n511 VSUBS 0.007624f
C552 B.n512 VSUBS 0.007624f
C553 B.n513 VSUBS 0.007624f
C554 B.n514 VSUBS 0.007624f
C555 B.n515 VSUBS 0.007624f
C556 B.n516 VSUBS 0.007624f
C557 B.n517 VSUBS 0.007624f
C558 B.n518 VSUBS 0.007624f
C559 B.n519 VSUBS 0.007624f
C560 B.n520 VSUBS 0.007624f
C561 B.n521 VSUBS 0.00527f
C562 B.n522 VSUBS 0.007624f
C563 B.n523 VSUBS 0.007624f
C564 B.n524 VSUBS 0.006167f
C565 B.n525 VSUBS 0.007624f
C566 B.n526 VSUBS 0.007624f
C567 B.n527 VSUBS 0.007624f
C568 B.n528 VSUBS 0.007624f
C569 B.n529 VSUBS 0.007624f
C570 B.n530 VSUBS 0.007624f
C571 B.n531 VSUBS 0.007624f
C572 B.n532 VSUBS 0.007624f
C573 B.n533 VSUBS 0.007624f
C574 B.n534 VSUBS 0.007624f
C575 B.n535 VSUBS 0.007624f
C576 B.n536 VSUBS 0.006167f
C577 B.n537 VSUBS 0.017665f
C578 B.n538 VSUBS 0.00527f
C579 B.n539 VSUBS 0.007624f
C580 B.n540 VSUBS 0.007624f
C581 B.n541 VSUBS 0.007624f
C582 B.n542 VSUBS 0.007624f
C583 B.n543 VSUBS 0.007624f
C584 B.n544 VSUBS 0.007624f
C585 B.n545 VSUBS 0.007624f
C586 B.n546 VSUBS 0.007624f
C587 B.n547 VSUBS 0.007624f
C588 B.n548 VSUBS 0.007624f
C589 B.n549 VSUBS 0.007624f
C590 B.n550 VSUBS 0.007624f
C591 B.n551 VSUBS 0.007624f
C592 B.n552 VSUBS 0.007624f
C593 B.n553 VSUBS 0.007624f
C594 B.n554 VSUBS 0.007624f
C595 B.n555 VSUBS 0.007624f
C596 B.n556 VSUBS 0.007624f
C597 B.n557 VSUBS 0.007624f
C598 B.n558 VSUBS 0.007624f
C599 B.n559 VSUBS 0.007624f
C600 B.n560 VSUBS 0.007624f
C601 B.n561 VSUBS 0.007624f
C602 B.n562 VSUBS 0.007624f
C603 B.n563 VSUBS 0.007624f
C604 B.n564 VSUBS 0.007624f
C605 B.n565 VSUBS 0.007624f
C606 B.n566 VSUBS 0.007624f
C607 B.n567 VSUBS 0.007624f
C608 B.n568 VSUBS 0.007624f
C609 B.n569 VSUBS 0.007624f
C610 B.n570 VSUBS 0.007624f
C611 B.n571 VSUBS 0.007624f
C612 B.n572 VSUBS 0.007624f
C613 B.n573 VSUBS 0.007624f
C614 B.n574 VSUBS 0.007624f
C615 B.n575 VSUBS 0.007624f
C616 B.n576 VSUBS 0.007624f
C617 B.n577 VSUBS 0.007624f
C618 B.n578 VSUBS 0.007624f
C619 B.n579 VSUBS 0.007624f
C620 B.n580 VSUBS 0.007624f
C621 B.n581 VSUBS 0.007624f
C622 B.n582 VSUBS 0.007624f
C623 B.n583 VSUBS 0.018583f
C624 B.n584 VSUBS 0.017969f
C625 B.n585 VSUBS 0.017969f
C626 B.n586 VSUBS 0.007624f
C627 B.n587 VSUBS 0.007624f
C628 B.n588 VSUBS 0.007624f
C629 B.n589 VSUBS 0.007624f
C630 B.n590 VSUBS 0.007624f
C631 B.n591 VSUBS 0.007624f
C632 B.n592 VSUBS 0.007624f
C633 B.n593 VSUBS 0.007624f
C634 B.n594 VSUBS 0.007624f
C635 B.n595 VSUBS 0.007624f
C636 B.n596 VSUBS 0.007624f
C637 B.n597 VSUBS 0.007624f
C638 B.n598 VSUBS 0.007624f
C639 B.n599 VSUBS 0.007624f
C640 B.n600 VSUBS 0.007624f
C641 B.n601 VSUBS 0.007624f
C642 B.n602 VSUBS 0.007624f
C643 B.n603 VSUBS 0.007624f
C644 B.n604 VSUBS 0.007624f
C645 B.n605 VSUBS 0.007624f
C646 B.n606 VSUBS 0.007624f
C647 B.n607 VSUBS 0.007624f
C648 B.n608 VSUBS 0.007624f
C649 B.n609 VSUBS 0.007624f
C650 B.n610 VSUBS 0.007624f
C651 B.n611 VSUBS 0.007624f
C652 B.n612 VSUBS 0.007624f
C653 B.n613 VSUBS 0.007624f
C654 B.n614 VSUBS 0.007624f
C655 B.n615 VSUBS 0.007624f
C656 B.n616 VSUBS 0.007624f
C657 B.n617 VSUBS 0.007624f
C658 B.n618 VSUBS 0.007624f
C659 B.n619 VSUBS 0.007624f
C660 B.n620 VSUBS 0.007624f
C661 B.n621 VSUBS 0.007624f
C662 B.n622 VSUBS 0.007624f
C663 B.n623 VSUBS 0.007624f
C664 B.n624 VSUBS 0.007624f
C665 B.n625 VSUBS 0.007624f
C666 B.n626 VSUBS 0.007624f
C667 B.n627 VSUBS 0.007624f
C668 B.n628 VSUBS 0.007624f
C669 B.n629 VSUBS 0.007624f
C670 B.n630 VSUBS 0.007624f
C671 B.n631 VSUBS 0.007624f
C672 B.n632 VSUBS 0.007624f
C673 B.n633 VSUBS 0.007624f
C674 B.n634 VSUBS 0.007624f
C675 B.n635 VSUBS 0.007624f
C676 B.n636 VSUBS 0.007624f
C677 B.n637 VSUBS 0.007624f
C678 B.n638 VSUBS 0.007624f
C679 B.n639 VSUBS 0.007624f
C680 B.n640 VSUBS 0.007624f
C681 B.n641 VSUBS 0.007624f
C682 B.n642 VSUBS 0.007624f
C683 B.n643 VSUBS 0.007624f
C684 B.n644 VSUBS 0.007624f
C685 B.n645 VSUBS 0.007624f
C686 B.n646 VSUBS 0.007624f
C687 B.n647 VSUBS 0.007624f
C688 B.n648 VSUBS 0.007624f
C689 B.n649 VSUBS 0.007624f
C690 B.n650 VSUBS 0.007624f
C691 B.n651 VSUBS 0.017265f
C692 VDD2.t0 VSUBS 0.160496f
C693 VDD2.t6 VSUBS 0.160496f
C694 VDD2.n0 VSUBS 1.18339f
C695 VDD2.t1 VSUBS 0.160496f
C696 VDD2.t7 VSUBS 0.160496f
C697 VDD2.n1 VSUBS 1.18339f
C698 VDD2.n2 VSUBS 3.12107f
C699 VDD2.t3 VSUBS 0.160496f
C700 VDD2.t5 VSUBS 0.160496f
C701 VDD2.n3 VSUBS 1.17564f
C702 VDD2.n4 VSUBS 2.64555f
C703 VDD2.t2 VSUBS 0.160496f
C704 VDD2.t4 VSUBS 0.160496f
C705 VDD2.n5 VSUBS 1.18335f
C706 VN.n0 VSUBS 0.047196f
C707 VN.t0 VSUBS 1.69496f
C708 VN.n1 VSUBS 0.046098f
C709 VN.n2 VSUBS 0.0358f
C710 VN.t6 VSUBS 1.69496f
C711 VN.n3 VSUBS 0.052041f
C712 VN.n4 VSUBS 0.301606f
C713 VN.t1 VSUBS 1.69496f
C714 VN.t7 VSUBS 1.91029f
C715 VN.n5 VSUBS 0.696285f
C716 VN.n6 VSUBS 0.72586f
C717 VN.n7 VSUBS 0.064422f
C718 VN.n8 VSUBS 0.052041f
C719 VN.n9 VSUBS 0.0358f
C720 VN.n10 VSUBS 0.0358f
C721 VN.n11 VSUBS 0.0358f
C722 VN.n12 VSUBS 0.064422f
C723 VN.n13 VSUBS 0.621282f
C724 VN.n14 VSUBS 0.03558f
C725 VN.n15 VSUBS 0.066388f
C726 VN.n16 VSUBS 0.0358f
C727 VN.n17 VSUBS 0.0358f
C728 VN.n18 VSUBS 0.0358f
C729 VN.n19 VSUBS 0.057984f
C730 VN.n20 VSUBS 0.060489f
C731 VN.n21 VSUBS 0.736927f
C732 VN.n22 VSUBS 0.04379f
C733 VN.n23 VSUBS 0.047196f
C734 VN.t4 VSUBS 1.69496f
C735 VN.n24 VSUBS 0.046098f
C736 VN.n25 VSUBS 0.0358f
C737 VN.t2 VSUBS 1.69496f
C738 VN.n26 VSUBS 0.052041f
C739 VN.n27 VSUBS 0.301606f
C740 VN.t5 VSUBS 1.69496f
C741 VN.t3 VSUBS 1.91029f
C742 VN.n28 VSUBS 0.696285f
C743 VN.n29 VSUBS 0.72586f
C744 VN.n30 VSUBS 0.064422f
C745 VN.n31 VSUBS 0.052041f
C746 VN.n32 VSUBS 0.0358f
C747 VN.n33 VSUBS 0.0358f
C748 VN.n34 VSUBS 0.0358f
C749 VN.n35 VSUBS 0.064422f
C750 VN.n36 VSUBS 0.621282f
C751 VN.n37 VSUBS 0.03558f
C752 VN.n38 VSUBS 0.066388f
C753 VN.n39 VSUBS 0.0358f
C754 VN.n40 VSUBS 0.0358f
C755 VN.n41 VSUBS 0.0358f
C756 VN.n42 VSUBS 0.057984f
C757 VN.n43 VSUBS 0.060489f
C758 VN.n44 VSUBS 0.736927f
C759 VN.n45 VSUBS 1.7559f
C760 VDD1.t0 VSUBS 0.163153f
C761 VDD1.t6 VSUBS 0.163153f
C762 VDD1.n0 VSUBS 1.20397f
C763 VDD1.t5 VSUBS 0.163153f
C764 VDD1.t1 VSUBS 0.163153f
C765 VDD1.n1 VSUBS 1.20297f
C766 VDD1.t4 VSUBS 0.163153f
C767 VDD1.t7 VSUBS 0.163153f
C768 VDD1.n2 VSUBS 1.20297f
C769 VDD1.n3 VSUBS 3.22471f
C770 VDD1.t3 VSUBS 0.163153f
C771 VDD1.t2 VSUBS 0.163153f
C772 VDD1.n4 VSUBS 1.19509f
C773 VDD1.n5 VSUBS 2.71952f
C774 VTAIL.t7 VSUBS 0.173203f
C775 VTAIL.t1 VSUBS 0.173203f
C776 VTAIL.n0 VSUBS 1.16065f
C777 VTAIL.n1 VSUBS 0.701608f
C778 VTAIL.t3 VSUBS 1.55399f
C779 VTAIL.n2 VSUBS 0.815499f
C780 VTAIL.t14 VSUBS 1.55399f
C781 VTAIL.n3 VSUBS 0.815499f
C782 VTAIL.t15 VSUBS 0.173203f
C783 VTAIL.t10 VSUBS 0.173203f
C784 VTAIL.n4 VSUBS 1.16065f
C785 VTAIL.n5 VSUBS 0.874805f
C786 VTAIL.t13 VSUBS 1.55399f
C787 VTAIL.n6 VSUBS 1.91966f
C788 VTAIL.t4 VSUBS 1.554f
C789 VTAIL.n7 VSUBS 1.91965f
C790 VTAIL.t6 VSUBS 0.173203f
C791 VTAIL.t5 VSUBS 0.173203f
C792 VTAIL.n8 VSUBS 1.16065f
C793 VTAIL.n9 VSUBS 0.8748f
C794 VTAIL.t0 VSUBS 1.554f
C795 VTAIL.n10 VSUBS 0.815488f
C796 VTAIL.t9 VSUBS 1.554f
C797 VTAIL.n11 VSUBS 0.815488f
C798 VTAIL.t12 VSUBS 0.173203f
C799 VTAIL.t11 VSUBS 0.173203f
C800 VTAIL.n12 VSUBS 1.16065f
C801 VTAIL.n13 VSUBS 0.8748f
C802 VTAIL.t8 VSUBS 1.55399f
C803 VTAIL.n14 VSUBS 1.91966f
C804 VTAIL.t2 VSUBS 1.55399f
C805 VTAIL.n15 VSUBS 1.91474f
C806 VP.n0 VSUBS 0.048786f
C807 VP.t0 VSUBS 1.75204f
C808 VP.n1 VSUBS 0.047651f
C809 VP.n2 VSUBS 0.037006f
C810 VP.t3 VSUBS 1.75204f
C811 VP.n3 VSUBS 0.053793f
C812 VP.n4 VSUBS 0.037006f
C813 VP.t6 VSUBS 1.75204f
C814 VP.n5 VSUBS 0.068624f
C815 VP.n6 VSUBS 0.037006f
C816 VP.t2 VSUBS 1.75204f
C817 VP.n7 VSUBS 0.761744f
C818 VP.n8 VSUBS 0.048786f
C819 VP.t5 VSUBS 1.75204f
C820 VP.n9 VSUBS 0.047651f
C821 VP.n10 VSUBS 0.037006f
C822 VP.t4 VSUBS 1.75204f
C823 VP.n11 VSUBS 0.053793f
C824 VP.n12 VSUBS 0.311763f
C825 VP.t1 VSUBS 1.75204f
C826 VP.t7 VSUBS 1.97462f
C827 VP.n13 VSUBS 0.719734f
C828 VP.n14 VSUBS 0.750304f
C829 VP.n15 VSUBS 0.066591f
C830 VP.n16 VSUBS 0.053793f
C831 VP.n17 VSUBS 0.037006f
C832 VP.n18 VSUBS 0.037006f
C833 VP.n19 VSUBS 0.037006f
C834 VP.n20 VSUBS 0.066591f
C835 VP.n21 VSUBS 0.642204f
C836 VP.n22 VSUBS 0.036779f
C837 VP.n23 VSUBS 0.068624f
C838 VP.n24 VSUBS 0.037006f
C839 VP.n25 VSUBS 0.037006f
C840 VP.n26 VSUBS 0.037006f
C841 VP.n27 VSUBS 0.059937f
C842 VP.n28 VSUBS 0.062526f
C843 VP.n29 VSUBS 0.761744f
C844 VP.n30 VSUBS 1.79487f
C845 VP.n31 VSUBS 1.82394f
C846 VP.n32 VSUBS 0.048786f
C847 VP.n33 VSUBS 0.062526f
C848 VP.n34 VSUBS 0.059937f
C849 VP.n35 VSUBS 0.047651f
C850 VP.n36 VSUBS 0.037006f
C851 VP.n37 VSUBS 0.037006f
C852 VP.n38 VSUBS 0.037006f
C853 VP.n39 VSUBS 0.036779f
C854 VP.n40 VSUBS 0.642204f
C855 VP.n41 VSUBS 0.066591f
C856 VP.n42 VSUBS 0.053793f
C857 VP.n43 VSUBS 0.037006f
C858 VP.n44 VSUBS 0.037006f
C859 VP.n45 VSUBS 0.037006f
C860 VP.n46 VSUBS 0.066591f
C861 VP.n47 VSUBS 0.642204f
C862 VP.n48 VSUBS 0.036779f
C863 VP.n49 VSUBS 0.068624f
C864 VP.n50 VSUBS 0.037006f
C865 VP.n51 VSUBS 0.037006f
C866 VP.n52 VSUBS 0.037006f
C867 VP.n53 VSUBS 0.059937f
C868 VP.n54 VSUBS 0.062526f
C869 VP.n55 VSUBS 0.761744f
C870 VP.n56 VSUBS 0.045265f
.ends

