* NGSPICE file created from diff_pair_sample_0282.ext - technology: sky130A

.subckt diff_pair_sample_0282 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t4 VP.t0 VDD1.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=0.8736 pd=5.26 as=0.3696 ps=2.57 w=2.24 l=1.29
X1 B.t17 B.t15 B.t16 B.t5 sky130_fd_pr__nfet_01v8 ad=0.8736 pd=5.26 as=0 ps=0 w=2.24 l=1.29
X2 VTAIL.t3 VP.t1 VDD1.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=0.8736 pd=5.26 as=0.3696 ps=2.57 w=2.24 l=1.29
X3 VDD2.t3 VN.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.3696 pd=2.57 as=0.8736 ps=5.26 w=2.24 l=1.29
X4 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=0.8736 pd=5.26 as=0 ps=0 w=2.24 l=1.29
X5 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=0.8736 pd=5.26 as=0 ps=0 w=2.24 l=1.29
X6 VDD1.t2 VP.t2 VTAIL.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=0.3696 pd=2.57 as=0.8736 ps=5.26 w=2.24 l=1.29
X7 VDD1.t0 VP.t3 VTAIL.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=0.3696 pd=2.57 as=0.8736 ps=5.26 w=2.24 l=1.29
X8 VTAIL.t5 VN.t1 VDD2.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=0.8736 pd=5.26 as=0.3696 ps=2.57 w=2.24 l=1.29
X9 VDD2.t1 VN.t2 VTAIL.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=0.3696 pd=2.57 as=0.8736 ps=5.26 w=2.24 l=1.29
X10 VTAIL.t7 VN.t3 VDD2.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=0.8736 pd=5.26 as=0.3696 ps=2.57 w=2.24 l=1.29
X11 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=0.8736 pd=5.26 as=0 ps=0 w=2.24 l=1.29
R0 VP.n4 VP.n3 170.645
R1 VP.n10 VP.n9 170.645
R2 VP.n8 VP.n0 161.3
R3 VP.n7 VP.n6 161.3
R4 VP.n5 VP.n1 161.3
R5 VP.n2 VP.t0 79.2587
R6 VP.n2 VP.t3 79.0324
R7 VP.n4 VP.n2 52.8438
R8 VP.n3 VP.t1 41.8486
R9 VP.n9 VP.t2 41.8486
R10 VP.n7 VP.n1 40.577
R11 VP.n8 VP.n7 40.577
R12 VP.n3 VP.n1 15.2474
R13 VP.n9 VP.n8 15.2474
R14 VP.n5 VP.n4 0.189894
R15 VP.n6 VP.n5 0.189894
R16 VP.n6 VP.n0 0.189894
R17 VP.n10 VP.n0 0.189894
R18 VP VP.n10 0.0516364
R19 VDD1 VDD1.n1 124.992
R20 VDD1 VDD1.n0 94.6894
R21 VDD1.n0 VDD1.t1 8.83979
R22 VDD1.n0 VDD1.t0 8.83979
R23 VDD1.n1 VDD1.t3 8.83979
R24 VDD1.n1 VDD1.t2 8.83979
R25 VTAIL.n6 VTAIL.t1 86.7917
R26 VTAIL.n7 VTAIL.t0 86.7917
R27 VTAIL.n0 VTAIL.t5 86.7917
R28 VTAIL.n1 VTAIL.t2 86.7917
R29 VTAIL.n2 VTAIL.t3 86.7917
R30 VTAIL.n5 VTAIL.t4 86.7916
R31 VTAIL.n4 VTAIL.t6 86.7916
R32 VTAIL.n3 VTAIL.t7 86.7916
R33 VTAIL.n7 VTAIL.n6 15.6945
R34 VTAIL.n3 VTAIL.n2 15.6945
R35 VTAIL.n4 VTAIL.n3 1.39705
R36 VTAIL.n6 VTAIL.n5 1.39705
R37 VTAIL.n2 VTAIL.n1 1.39705
R38 VTAIL VTAIL.n0 0.756965
R39 VTAIL VTAIL.n7 0.640586
R40 VTAIL.n5 VTAIL.n4 0.470328
R41 VTAIL.n1 VTAIL.n0 0.470328
R42 B.n299 B.n66 585
R43 B.n66 B.n43 585
R44 B.n301 B.n300 585
R45 B.n303 B.n65 585
R46 B.n306 B.n305 585
R47 B.n307 B.n64 585
R48 B.n309 B.n308 585
R49 B.n311 B.n63 585
R50 B.n314 B.n313 585
R51 B.n315 B.n62 585
R52 B.n317 B.n316 585
R53 B.n319 B.n61 585
R54 B.n321 B.n320 585
R55 B.n323 B.n322 585
R56 B.n326 B.n325 585
R57 B.n327 B.n56 585
R58 B.n329 B.n328 585
R59 B.n331 B.n55 585
R60 B.n334 B.n333 585
R61 B.n335 B.n54 585
R62 B.n337 B.n336 585
R63 B.n339 B.n53 585
R64 B.n342 B.n341 585
R65 B.n344 B.n50 585
R66 B.n346 B.n345 585
R67 B.n348 B.n49 585
R68 B.n351 B.n350 585
R69 B.n352 B.n48 585
R70 B.n354 B.n353 585
R71 B.n356 B.n47 585
R72 B.n359 B.n358 585
R73 B.n360 B.n46 585
R74 B.n362 B.n361 585
R75 B.n364 B.n45 585
R76 B.n367 B.n366 585
R77 B.n368 B.n44 585
R78 B.n298 B.n42 585
R79 B.n371 B.n42 585
R80 B.n297 B.n41 585
R81 B.n372 B.n41 585
R82 B.n296 B.n40 585
R83 B.n373 B.n40 585
R84 B.n295 B.n294 585
R85 B.n294 B.n36 585
R86 B.n293 B.n35 585
R87 B.n379 B.n35 585
R88 B.n292 B.n34 585
R89 B.n380 B.n34 585
R90 B.n291 B.n33 585
R91 B.n381 B.n33 585
R92 B.n290 B.n289 585
R93 B.n289 B.n29 585
R94 B.n288 B.n28 585
R95 B.n387 B.n28 585
R96 B.n287 B.n27 585
R97 B.n388 B.n27 585
R98 B.n286 B.n26 585
R99 B.n389 B.n26 585
R100 B.n285 B.n284 585
R101 B.n284 B.n22 585
R102 B.n283 B.n21 585
R103 B.n395 B.n21 585
R104 B.n282 B.n20 585
R105 B.n396 B.n20 585
R106 B.n281 B.n19 585
R107 B.n397 B.n19 585
R108 B.n280 B.n279 585
R109 B.n279 B.n15 585
R110 B.n278 B.n14 585
R111 B.n403 B.n14 585
R112 B.n277 B.n13 585
R113 B.n404 B.n13 585
R114 B.n276 B.n12 585
R115 B.n405 B.n12 585
R116 B.n275 B.n274 585
R117 B.n274 B.n273 585
R118 B.n272 B.n271 585
R119 B.n272 B.n8 585
R120 B.n270 B.n7 585
R121 B.n412 B.n7 585
R122 B.n269 B.n6 585
R123 B.n413 B.n6 585
R124 B.n268 B.n5 585
R125 B.n414 B.n5 585
R126 B.n267 B.n266 585
R127 B.n266 B.n4 585
R128 B.n265 B.n67 585
R129 B.n265 B.n264 585
R130 B.n255 B.n68 585
R131 B.n69 B.n68 585
R132 B.n257 B.n256 585
R133 B.n258 B.n257 585
R134 B.n254 B.n74 585
R135 B.n74 B.n73 585
R136 B.n253 B.n252 585
R137 B.n252 B.n251 585
R138 B.n76 B.n75 585
R139 B.n77 B.n76 585
R140 B.n244 B.n243 585
R141 B.n245 B.n244 585
R142 B.n242 B.n81 585
R143 B.n85 B.n81 585
R144 B.n241 B.n240 585
R145 B.n240 B.n239 585
R146 B.n83 B.n82 585
R147 B.n84 B.n83 585
R148 B.n232 B.n231 585
R149 B.n233 B.n232 585
R150 B.n230 B.n90 585
R151 B.n90 B.n89 585
R152 B.n229 B.n228 585
R153 B.n228 B.n227 585
R154 B.n92 B.n91 585
R155 B.n93 B.n92 585
R156 B.n220 B.n219 585
R157 B.n221 B.n220 585
R158 B.n218 B.n97 585
R159 B.n101 B.n97 585
R160 B.n217 B.n216 585
R161 B.n216 B.n215 585
R162 B.n99 B.n98 585
R163 B.n100 B.n99 585
R164 B.n208 B.n207 585
R165 B.n209 B.n208 585
R166 B.n206 B.n106 585
R167 B.n106 B.n105 585
R168 B.n205 B.n204 585
R169 B.n204 B.n203 585
R170 B.n200 B.n110 585
R171 B.n199 B.n198 585
R172 B.n196 B.n111 585
R173 B.n196 B.n109 585
R174 B.n195 B.n194 585
R175 B.n193 B.n192 585
R176 B.n191 B.n113 585
R177 B.n189 B.n188 585
R178 B.n187 B.n114 585
R179 B.n186 B.n185 585
R180 B.n183 B.n115 585
R181 B.n181 B.n180 585
R182 B.n179 B.n116 585
R183 B.n178 B.n177 585
R184 B.n175 B.n174 585
R185 B.n173 B.n172 585
R186 B.n171 B.n121 585
R187 B.n169 B.n168 585
R188 B.n167 B.n122 585
R189 B.n166 B.n165 585
R190 B.n163 B.n123 585
R191 B.n161 B.n160 585
R192 B.n159 B.n124 585
R193 B.n157 B.n156 585
R194 B.n154 B.n127 585
R195 B.n152 B.n151 585
R196 B.n150 B.n128 585
R197 B.n149 B.n148 585
R198 B.n146 B.n129 585
R199 B.n144 B.n143 585
R200 B.n142 B.n130 585
R201 B.n141 B.n140 585
R202 B.n138 B.n131 585
R203 B.n136 B.n135 585
R204 B.n134 B.n133 585
R205 B.n108 B.n107 585
R206 B.n202 B.n201 585
R207 B.n203 B.n202 585
R208 B.n104 B.n103 585
R209 B.n105 B.n104 585
R210 B.n211 B.n210 585
R211 B.n210 B.n209 585
R212 B.n212 B.n102 585
R213 B.n102 B.n100 585
R214 B.n214 B.n213 585
R215 B.n215 B.n214 585
R216 B.n96 B.n95 585
R217 B.n101 B.n96 585
R218 B.n223 B.n222 585
R219 B.n222 B.n221 585
R220 B.n224 B.n94 585
R221 B.n94 B.n93 585
R222 B.n226 B.n225 585
R223 B.n227 B.n226 585
R224 B.n88 B.n87 585
R225 B.n89 B.n88 585
R226 B.n235 B.n234 585
R227 B.n234 B.n233 585
R228 B.n236 B.n86 585
R229 B.n86 B.n84 585
R230 B.n238 B.n237 585
R231 B.n239 B.n238 585
R232 B.n80 B.n79 585
R233 B.n85 B.n80 585
R234 B.n247 B.n246 585
R235 B.n246 B.n245 585
R236 B.n248 B.n78 585
R237 B.n78 B.n77 585
R238 B.n250 B.n249 585
R239 B.n251 B.n250 585
R240 B.n72 B.n71 585
R241 B.n73 B.n72 585
R242 B.n260 B.n259 585
R243 B.n259 B.n258 585
R244 B.n261 B.n70 585
R245 B.n70 B.n69 585
R246 B.n263 B.n262 585
R247 B.n264 B.n263 585
R248 B.n3 B.n0 585
R249 B.n4 B.n3 585
R250 B.n411 B.n1 585
R251 B.n412 B.n411 585
R252 B.n410 B.n409 585
R253 B.n410 B.n8 585
R254 B.n408 B.n9 585
R255 B.n273 B.n9 585
R256 B.n407 B.n406 585
R257 B.n406 B.n405 585
R258 B.n11 B.n10 585
R259 B.n404 B.n11 585
R260 B.n402 B.n401 585
R261 B.n403 B.n402 585
R262 B.n400 B.n16 585
R263 B.n16 B.n15 585
R264 B.n399 B.n398 585
R265 B.n398 B.n397 585
R266 B.n18 B.n17 585
R267 B.n396 B.n18 585
R268 B.n394 B.n393 585
R269 B.n395 B.n394 585
R270 B.n392 B.n23 585
R271 B.n23 B.n22 585
R272 B.n391 B.n390 585
R273 B.n390 B.n389 585
R274 B.n25 B.n24 585
R275 B.n388 B.n25 585
R276 B.n386 B.n385 585
R277 B.n387 B.n386 585
R278 B.n384 B.n30 585
R279 B.n30 B.n29 585
R280 B.n383 B.n382 585
R281 B.n382 B.n381 585
R282 B.n32 B.n31 585
R283 B.n380 B.n32 585
R284 B.n378 B.n377 585
R285 B.n379 B.n378 585
R286 B.n376 B.n37 585
R287 B.n37 B.n36 585
R288 B.n375 B.n374 585
R289 B.n374 B.n373 585
R290 B.n39 B.n38 585
R291 B.n372 B.n39 585
R292 B.n370 B.n369 585
R293 B.n371 B.n370 585
R294 B.n415 B.n414 585
R295 B.n413 B.n2 585
R296 B.n370 B.n44 516.524
R297 B.n66 B.n42 516.524
R298 B.n204 B.n108 516.524
R299 B.n202 B.n110 516.524
R300 B.n302 B.n43 256.663
R301 B.n304 B.n43 256.663
R302 B.n310 B.n43 256.663
R303 B.n312 B.n43 256.663
R304 B.n318 B.n43 256.663
R305 B.n60 B.n43 256.663
R306 B.n324 B.n43 256.663
R307 B.n330 B.n43 256.663
R308 B.n332 B.n43 256.663
R309 B.n338 B.n43 256.663
R310 B.n340 B.n43 256.663
R311 B.n347 B.n43 256.663
R312 B.n349 B.n43 256.663
R313 B.n355 B.n43 256.663
R314 B.n357 B.n43 256.663
R315 B.n363 B.n43 256.663
R316 B.n365 B.n43 256.663
R317 B.n197 B.n109 256.663
R318 B.n112 B.n109 256.663
R319 B.n190 B.n109 256.663
R320 B.n184 B.n109 256.663
R321 B.n182 B.n109 256.663
R322 B.n176 B.n109 256.663
R323 B.n120 B.n109 256.663
R324 B.n170 B.n109 256.663
R325 B.n164 B.n109 256.663
R326 B.n162 B.n109 256.663
R327 B.n155 B.n109 256.663
R328 B.n153 B.n109 256.663
R329 B.n147 B.n109 256.663
R330 B.n145 B.n109 256.663
R331 B.n139 B.n109 256.663
R332 B.n137 B.n109 256.663
R333 B.n132 B.n109 256.663
R334 B.n417 B.n416 256.663
R335 B.n51 B.t12 246.411
R336 B.n57 B.t8 246.411
R337 B.n125 B.t4 246.411
R338 B.n117 B.t15 246.411
R339 B.n203 B.n109 171.257
R340 B.n371 B.n43 171.257
R341 B.n366 B.n364 163.367
R342 B.n362 B.n46 163.367
R343 B.n358 B.n356 163.367
R344 B.n354 B.n48 163.367
R345 B.n350 B.n348 163.367
R346 B.n346 B.n50 163.367
R347 B.n341 B.n339 163.367
R348 B.n337 B.n54 163.367
R349 B.n333 B.n331 163.367
R350 B.n329 B.n56 163.367
R351 B.n325 B.n323 163.367
R352 B.n320 B.n319 163.367
R353 B.n317 B.n62 163.367
R354 B.n313 B.n311 163.367
R355 B.n309 B.n64 163.367
R356 B.n305 B.n303 163.367
R357 B.n301 B.n66 163.367
R358 B.n204 B.n106 163.367
R359 B.n208 B.n106 163.367
R360 B.n208 B.n99 163.367
R361 B.n216 B.n99 163.367
R362 B.n216 B.n97 163.367
R363 B.n220 B.n97 163.367
R364 B.n220 B.n92 163.367
R365 B.n228 B.n92 163.367
R366 B.n228 B.n90 163.367
R367 B.n232 B.n90 163.367
R368 B.n232 B.n83 163.367
R369 B.n240 B.n83 163.367
R370 B.n240 B.n81 163.367
R371 B.n244 B.n81 163.367
R372 B.n244 B.n76 163.367
R373 B.n252 B.n76 163.367
R374 B.n252 B.n74 163.367
R375 B.n257 B.n74 163.367
R376 B.n257 B.n68 163.367
R377 B.n265 B.n68 163.367
R378 B.n266 B.n265 163.367
R379 B.n266 B.n5 163.367
R380 B.n6 B.n5 163.367
R381 B.n7 B.n6 163.367
R382 B.n272 B.n7 163.367
R383 B.n274 B.n272 163.367
R384 B.n274 B.n12 163.367
R385 B.n13 B.n12 163.367
R386 B.n14 B.n13 163.367
R387 B.n279 B.n14 163.367
R388 B.n279 B.n19 163.367
R389 B.n20 B.n19 163.367
R390 B.n21 B.n20 163.367
R391 B.n284 B.n21 163.367
R392 B.n284 B.n26 163.367
R393 B.n27 B.n26 163.367
R394 B.n28 B.n27 163.367
R395 B.n289 B.n28 163.367
R396 B.n289 B.n33 163.367
R397 B.n34 B.n33 163.367
R398 B.n35 B.n34 163.367
R399 B.n294 B.n35 163.367
R400 B.n294 B.n40 163.367
R401 B.n41 B.n40 163.367
R402 B.n42 B.n41 163.367
R403 B.n198 B.n196 163.367
R404 B.n196 B.n195 163.367
R405 B.n192 B.n191 163.367
R406 B.n189 B.n114 163.367
R407 B.n185 B.n183 163.367
R408 B.n181 B.n116 163.367
R409 B.n177 B.n175 163.367
R410 B.n172 B.n171 163.367
R411 B.n169 B.n122 163.367
R412 B.n165 B.n163 163.367
R413 B.n161 B.n124 163.367
R414 B.n156 B.n154 163.367
R415 B.n152 B.n128 163.367
R416 B.n148 B.n146 163.367
R417 B.n144 B.n130 163.367
R418 B.n140 B.n138 163.367
R419 B.n136 B.n133 163.367
R420 B.n202 B.n104 163.367
R421 B.n210 B.n104 163.367
R422 B.n210 B.n102 163.367
R423 B.n214 B.n102 163.367
R424 B.n214 B.n96 163.367
R425 B.n222 B.n96 163.367
R426 B.n222 B.n94 163.367
R427 B.n226 B.n94 163.367
R428 B.n226 B.n88 163.367
R429 B.n234 B.n88 163.367
R430 B.n234 B.n86 163.367
R431 B.n238 B.n86 163.367
R432 B.n238 B.n80 163.367
R433 B.n246 B.n80 163.367
R434 B.n246 B.n78 163.367
R435 B.n250 B.n78 163.367
R436 B.n250 B.n72 163.367
R437 B.n259 B.n72 163.367
R438 B.n259 B.n70 163.367
R439 B.n263 B.n70 163.367
R440 B.n263 B.n3 163.367
R441 B.n415 B.n3 163.367
R442 B.n411 B.n2 163.367
R443 B.n411 B.n410 163.367
R444 B.n410 B.n9 163.367
R445 B.n406 B.n9 163.367
R446 B.n406 B.n11 163.367
R447 B.n402 B.n11 163.367
R448 B.n402 B.n16 163.367
R449 B.n398 B.n16 163.367
R450 B.n398 B.n18 163.367
R451 B.n394 B.n18 163.367
R452 B.n394 B.n23 163.367
R453 B.n390 B.n23 163.367
R454 B.n390 B.n25 163.367
R455 B.n386 B.n25 163.367
R456 B.n386 B.n30 163.367
R457 B.n382 B.n30 163.367
R458 B.n382 B.n32 163.367
R459 B.n378 B.n32 163.367
R460 B.n378 B.n37 163.367
R461 B.n374 B.n37 163.367
R462 B.n374 B.n39 163.367
R463 B.n370 B.n39 163.367
R464 B.n57 B.t10 117.742
R465 B.n125 B.t7 117.742
R466 B.n51 B.t13 117.74
R467 B.n117 B.t17 117.74
R468 B.n203 B.n105 99.5348
R469 B.n209 B.n105 99.5348
R470 B.n209 B.n100 99.5348
R471 B.n215 B.n100 99.5348
R472 B.n215 B.n101 99.5348
R473 B.n221 B.n93 99.5348
R474 B.n227 B.n93 99.5348
R475 B.n227 B.n89 99.5348
R476 B.n233 B.n89 99.5348
R477 B.n233 B.n84 99.5348
R478 B.n239 B.n84 99.5348
R479 B.n239 B.n85 99.5348
R480 B.n245 B.n77 99.5348
R481 B.n251 B.n77 99.5348
R482 B.n251 B.n73 99.5348
R483 B.n258 B.n73 99.5348
R484 B.n264 B.n69 99.5348
R485 B.n264 B.n4 99.5348
R486 B.n414 B.n4 99.5348
R487 B.n414 B.n413 99.5348
R488 B.n413 B.n412 99.5348
R489 B.n412 B.n8 99.5348
R490 B.n273 B.n8 99.5348
R491 B.n405 B.n404 99.5348
R492 B.n404 B.n403 99.5348
R493 B.n403 B.n15 99.5348
R494 B.n397 B.n15 99.5348
R495 B.n396 B.n395 99.5348
R496 B.n395 B.n22 99.5348
R497 B.n389 B.n22 99.5348
R498 B.n389 B.n388 99.5348
R499 B.n388 B.n387 99.5348
R500 B.n387 B.n29 99.5348
R501 B.n381 B.n29 99.5348
R502 B.n380 B.n379 99.5348
R503 B.n379 B.n36 99.5348
R504 B.n373 B.n36 99.5348
R505 B.n373 B.n372 99.5348
R506 B.n372 B.n371 99.5348
R507 B.n58 B.t11 86.3228
R508 B.n126 B.t6 86.3228
R509 B.n52 B.t14 86.3225
R510 B.n118 B.t16 86.3225
R511 B.n101 B.t5 77.5787
R512 B.t9 B.n380 77.5787
R513 B.n85 B.t2 74.6512
R514 B.t0 B.n396 74.6512
R515 B.n365 B.n44 71.676
R516 B.n364 B.n363 71.676
R517 B.n357 B.n46 71.676
R518 B.n356 B.n355 71.676
R519 B.n349 B.n48 71.676
R520 B.n348 B.n347 71.676
R521 B.n340 B.n50 71.676
R522 B.n339 B.n338 71.676
R523 B.n332 B.n54 71.676
R524 B.n331 B.n330 71.676
R525 B.n324 B.n56 71.676
R526 B.n323 B.n60 71.676
R527 B.n319 B.n318 71.676
R528 B.n312 B.n62 71.676
R529 B.n311 B.n310 71.676
R530 B.n304 B.n64 71.676
R531 B.n303 B.n302 71.676
R532 B.n302 B.n301 71.676
R533 B.n305 B.n304 71.676
R534 B.n310 B.n309 71.676
R535 B.n313 B.n312 71.676
R536 B.n318 B.n317 71.676
R537 B.n320 B.n60 71.676
R538 B.n325 B.n324 71.676
R539 B.n330 B.n329 71.676
R540 B.n333 B.n332 71.676
R541 B.n338 B.n337 71.676
R542 B.n341 B.n340 71.676
R543 B.n347 B.n346 71.676
R544 B.n350 B.n349 71.676
R545 B.n355 B.n354 71.676
R546 B.n358 B.n357 71.676
R547 B.n363 B.n362 71.676
R548 B.n366 B.n365 71.676
R549 B.n197 B.n110 71.676
R550 B.n195 B.n112 71.676
R551 B.n191 B.n190 71.676
R552 B.n184 B.n114 71.676
R553 B.n183 B.n182 71.676
R554 B.n176 B.n116 71.676
R555 B.n175 B.n120 71.676
R556 B.n171 B.n170 71.676
R557 B.n164 B.n122 71.676
R558 B.n163 B.n162 71.676
R559 B.n155 B.n124 71.676
R560 B.n154 B.n153 71.676
R561 B.n147 B.n128 71.676
R562 B.n146 B.n145 71.676
R563 B.n139 B.n130 71.676
R564 B.n138 B.n137 71.676
R565 B.n133 B.n132 71.676
R566 B.n198 B.n197 71.676
R567 B.n192 B.n112 71.676
R568 B.n190 B.n189 71.676
R569 B.n185 B.n184 71.676
R570 B.n182 B.n181 71.676
R571 B.n177 B.n176 71.676
R572 B.n172 B.n120 71.676
R573 B.n170 B.n169 71.676
R574 B.n165 B.n164 71.676
R575 B.n162 B.n161 71.676
R576 B.n156 B.n155 71.676
R577 B.n153 B.n152 71.676
R578 B.n148 B.n147 71.676
R579 B.n145 B.n144 71.676
R580 B.n140 B.n139 71.676
R581 B.n137 B.n136 71.676
R582 B.n132 B.n108 71.676
R583 B.n416 B.n415 71.676
R584 B.n416 B.n2 71.676
R585 B.n343 B.n52 59.5399
R586 B.n59 B.n58 59.5399
R587 B.n158 B.n126 59.5399
R588 B.n119 B.n118 59.5399
R589 B.n258 B.t1 51.2314
R590 B.n405 B.t3 51.2314
R591 B.t1 B.n69 48.3039
R592 B.n273 B.t3 48.3039
R593 B.n201 B.n200 33.5615
R594 B.n205 B.n107 33.5615
R595 B.n299 B.n298 33.5615
R596 B.n369 B.n368 33.5615
R597 B.n52 B.n51 31.4187
R598 B.n58 B.n57 31.4187
R599 B.n126 B.n125 31.4187
R600 B.n118 B.n117 31.4187
R601 B.n245 B.t2 24.8841
R602 B.n397 B.t0 24.8841
R603 B.n221 B.t5 21.9566
R604 B.n381 B.t9 21.9566
R605 B B.n417 18.0485
R606 B.n201 B.n103 10.6151
R607 B.n211 B.n103 10.6151
R608 B.n212 B.n211 10.6151
R609 B.n213 B.n212 10.6151
R610 B.n213 B.n95 10.6151
R611 B.n223 B.n95 10.6151
R612 B.n224 B.n223 10.6151
R613 B.n225 B.n224 10.6151
R614 B.n225 B.n87 10.6151
R615 B.n235 B.n87 10.6151
R616 B.n236 B.n235 10.6151
R617 B.n237 B.n236 10.6151
R618 B.n237 B.n79 10.6151
R619 B.n247 B.n79 10.6151
R620 B.n248 B.n247 10.6151
R621 B.n249 B.n248 10.6151
R622 B.n249 B.n71 10.6151
R623 B.n260 B.n71 10.6151
R624 B.n261 B.n260 10.6151
R625 B.n262 B.n261 10.6151
R626 B.n262 B.n0 10.6151
R627 B.n200 B.n199 10.6151
R628 B.n199 B.n111 10.6151
R629 B.n194 B.n111 10.6151
R630 B.n194 B.n193 10.6151
R631 B.n193 B.n113 10.6151
R632 B.n188 B.n113 10.6151
R633 B.n188 B.n187 10.6151
R634 B.n187 B.n186 10.6151
R635 B.n186 B.n115 10.6151
R636 B.n180 B.n115 10.6151
R637 B.n180 B.n179 10.6151
R638 B.n179 B.n178 10.6151
R639 B.n174 B.n173 10.6151
R640 B.n173 B.n121 10.6151
R641 B.n168 B.n121 10.6151
R642 B.n168 B.n167 10.6151
R643 B.n167 B.n166 10.6151
R644 B.n166 B.n123 10.6151
R645 B.n160 B.n123 10.6151
R646 B.n160 B.n159 10.6151
R647 B.n157 B.n127 10.6151
R648 B.n151 B.n127 10.6151
R649 B.n151 B.n150 10.6151
R650 B.n150 B.n149 10.6151
R651 B.n149 B.n129 10.6151
R652 B.n143 B.n129 10.6151
R653 B.n143 B.n142 10.6151
R654 B.n142 B.n141 10.6151
R655 B.n141 B.n131 10.6151
R656 B.n135 B.n131 10.6151
R657 B.n135 B.n134 10.6151
R658 B.n134 B.n107 10.6151
R659 B.n206 B.n205 10.6151
R660 B.n207 B.n206 10.6151
R661 B.n207 B.n98 10.6151
R662 B.n217 B.n98 10.6151
R663 B.n218 B.n217 10.6151
R664 B.n219 B.n218 10.6151
R665 B.n219 B.n91 10.6151
R666 B.n229 B.n91 10.6151
R667 B.n230 B.n229 10.6151
R668 B.n231 B.n230 10.6151
R669 B.n231 B.n82 10.6151
R670 B.n241 B.n82 10.6151
R671 B.n242 B.n241 10.6151
R672 B.n243 B.n242 10.6151
R673 B.n243 B.n75 10.6151
R674 B.n253 B.n75 10.6151
R675 B.n254 B.n253 10.6151
R676 B.n256 B.n254 10.6151
R677 B.n256 B.n255 10.6151
R678 B.n255 B.n67 10.6151
R679 B.n267 B.n67 10.6151
R680 B.n268 B.n267 10.6151
R681 B.n269 B.n268 10.6151
R682 B.n270 B.n269 10.6151
R683 B.n271 B.n270 10.6151
R684 B.n275 B.n271 10.6151
R685 B.n276 B.n275 10.6151
R686 B.n277 B.n276 10.6151
R687 B.n278 B.n277 10.6151
R688 B.n280 B.n278 10.6151
R689 B.n281 B.n280 10.6151
R690 B.n282 B.n281 10.6151
R691 B.n283 B.n282 10.6151
R692 B.n285 B.n283 10.6151
R693 B.n286 B.n285 10.6151
R694 B.n287 B.n286 10.6151
R695 B.n288 B.n287 10.6151
R696 B.n290 B.n288 10.6151
R697 B.n291 B.n290 10.6151
R698 B.n292 B.n291 10.6151
R699 B.n293 B.n292 10.6151
R700 B.n295 B.n293 10.6151
R701 B.n296 B.n295 10.6151
R702 B.n297 B.n296 10.6151
R703 B.n298 B.n297 10.6151
R704 B.n409 B.n1 10.6151
R705 B.n409 B.n408 10.6151
R706 B.n408 B.n407 10.6151
R707 B.n407 B.n10 10.6151
R708 B.n401 B.n10 10.6151
R709 B.n401 B.n400 10.6151
R710 B.n400 B.n399 10.6151
R711 B.n399 B.n17 10.6151
R712 B.n393 B.n17 10.6151
R713 B.n393 B.n392 10.6151
R714 B.n392 B.n391 10.6151
R715 B.n391 B.n24 10.6151
R716 B.n385 B.n24 10.6151
R717 B.n385 B.n384 10.6151
R718 B.n384 B.n383 10.6151
R719 B.n383 B.n31 10.6151
R720 B.n377 B.n31 10.6151
R721 B.n377 B.n376 10.6151
R722 B.n376 B.n375 10.6151
R723 B.n375 B.n38 10.6151
R724 B.n369 B.n38 10.6151
R725 B.n368 B.n367 10.6151
R726 B.n367 B.n45 10.6151
R727 B.n361 B.n45 10.6151
R728 B.n361 B.n360 10.6151
R729 B.n360 B.n359 10.6151
R730 B.n359 B.n47 10.6151
R731 B.n353 B.n47 10.6151
R732 B.n353 B.n352 10.6151
R733 B.n352 B.n351 10.6151
R734 B.n351 B.n49 10.6151
R735 B.n345 B.n49 10.6151
R736 B.n345 B.n344 10.6151
R737 B.n342 B.n53 10.6151
R738 B.n336 B.n53 10.6151
R739 B.n336 B.n335 10.6151
R740 B.n335 B.n334 10.6151
R741 B.n334 B.n55 10.6151
R742 B.n328 B.n55 10.6151
R743 B.n328 B.n327 10.6151
R744 B.n327 B.n326 10.6151
R745 B.n322 B.n321 10.6151
R746 B.n321 B.n61 10.6151
R747 B.n316 B.n61 10.6151
R748 B.n316 B.n315 10.6151
R749 B.n315 B.n314 10.6151
R750 B.n314 B.n63 10.6151
R751 B.n308 B.n63 10.6151
R752 B.n308 B.n307 10.6151
R753 B.n307 B.n306 10.6151
R754 B.n306 B.n65 10.6151
R755 B.n300 B.n65 10.6151
R756 B.n300 B.n299 10.6151
R757 B.n417 B.n0 8.11757
R758 B.n417 B.n1 8.11757
R759 B.n174 B.n119 6.5566
R760 B.n159 B.n158 6.5566
R761 B.n343 B.n342 6.5566
R762 B.n326 B.n59 6.5566
R763 B.n178 B.n119 4.05904
R764 B.n158 B.n157 4.05904
R765 B.n344 B.n343 4.05904
R766 B.n322 B.n59 4.05904
R767 VN.n0 VN.t1 79.2587
R768 VN.n1 VN.t2 79.2587
R769 VN.n0 VN.t0 79.0324
R770 VN.n1 VN.t3 79.0324
R771 VN VN.n1 53.2245
R772 VN VN.n0 18.0237
R773 VDD2.n2 VDD2.n0 124.466
R774 VDD2.n2 VDD2.n1 94.6313
R775 VDD2.n1 VDD2.t0 8.83979
R776 VDD2.n1 VDD2.t1 8.83979
R777 VDD2.n0 VDD2.t2 8.83979
R778 VDD2.n0 VDD2.t3 8.83979
R779 VDD2 VDD2.n2 0.0586897
C0 VN VP 3.44334f
C1 VDD2 VN 0.998039f
C2 VN VTAIL 1.22606f
C3 VDD1 VP 1.16073f
C4 VDD1 VDD2 0.706407f
C5 VDD1 VTAIL 2.52325f
C6 VDD1 VN 0.15349f
C7 VDD2 VP 0.317294f
C8 VP VTAIL 1.24016f
C9 VDD2 VTAIL 2.56867f
C10 VDD2 B 2.225195f
C11 VDD1 B 4.08701f
C12 VTAIL B 3.312985f
C13 VN B 6.69446f
C14 VP B 5.31068f
C15 VDD2.t2 B 0.035278f
C16 VDD2.t3 B 0.035278f
C17 VDD2.n0 B 0.407899f
C18 VDD2.t0 B 0.035278f
C19 VDD2.t1 B 0.035278f
C20 VDD2.n1 B 0.240498f
C21 VDD2.n2 B 1.71651f
C22 VN.t1 B 0.270439f
C23 VN.t0 B 0.269902f
C24 VN.n0 B 0.227411f
C25 VN.t2 B 0.270439f
C26 VN.t3 B 0.269902f
C27 VN.n1 B 0.835007f
C28 VTAIL.t5 B 0.221403f
C29 VTAIL.n0 B 0.203017f
C30 VTAIL.t2 B 0.221403f
C31 VTAIL.n1 B 0.235672f
C32 VTAIL.t3 B 0.221403f
C33 VTAIL.n2 B 0.596523f
C34 VTAIL.t7 B 0.221404f
C35 VTAIL.n3 B 0.596522f
C36 VTAIL.t6 B 0.221404f
C37 VTAIL.n4 B 0.23567f
C38 VTAIL.t4 B 0.221404f
C39 VTAIL.n5 B 0.23567f
C40 VTAIL.t1 B 0.221402f
C41 VTAIL.n6 B 0.596523f
C42 VTAIL.t0 B 0.221403f
C43 VTAIL.n7 B 0.557932f
C44 VDD1.t1 B 0.032987f
C45 VDD1.t0 B 0.032987f
C46 VDD1.n0 B 0.225024f
C47 VDD1.t3 B 0.032987f
C48 VDD1.t2 B 0.032987f
C49 VDD1.n1 B 0.392798f
C50 VP.n0 B 0.026767f
C51 VP.t2 B 0.184502f
C52 VP.n1 B 0.043607f
C53 VP.t0 B 0.273432f
C54 VP.t3 B 0.272888f
C55 VP.n2 B 0.830246f
C56 VP.t1 B 0.184502f
C57 VP.n3 B 0.148308f
C58 VP.n4 B 1.13216f
C59 VP.n5 B 0.026767f
C60 VP.n6 B 0.026767f
C61 VP.n7 B 0.021619f
C62 VP.n8 B 0.043607f
C63 VP.n9 B 0.148308f
C64 VP.n10 B 0.02373f
.ends

