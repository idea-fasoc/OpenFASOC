* NGSPICE file created from diff_pair_sample_1474.ext - technology: sky130A

.subckt diff_pair_sample_1474 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t1 VP.t0 VTAIL.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=4.8945 pd=25.88 as=4.8945 ps=25.88 w=12.55 l=2.93
X1 B.t15 B.t13 B.t14 B.t3 sky130_fd_pr__nfet_01v8 ad=4.8945 pd=25.88 as=0 ps=0 w=12.55 l=2.93
X2 VDD1.t0 VP.t1 VTAIL.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=4.8945 pd=25.88 as=4.8945 ps=25.88 w=12.55 l=2.93
X3 VDD2.t1 VN.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=4.8945 pd=25.88 as=4.8945 ps=25.88 w=12.55 l=2.93
X4 VDD2.t0 VN.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=4.8945 pd=25.88 as=4.8945 ps=25.88 w=12.55 l=2.93
X5 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=4.8945 pd=25.88 as=0 ps=0 w=12.55 l=2.93
X6 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=4.8945 pd=25.88 as=0 ps=0 w=12.55 l=2.93
X7 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=4.8945 pd=25.88 as=0 ps=0 w=12.55 l=2.93
R0 VP.n0 VP.t1 190.272
R1 VP.n0 VP.t0 144.323
R2 VP VP.n0 0.431811
R3 VTAIL.n1 VTAIL.t0 48.044
R4 VTAIL.n3 VTAIL.t1 48.0438
R5 VTAIL.n0 VTAIL.t3 48.0438
R6 VTAIL.n2 VTAIL.t2 48.0438
R7 VTAIL.n1 VTAIL.n0 28.8065
R8 VTAIL.n3 VTAIL.n2 25.9962
R9 VTAIL.n2 VTAIL.n1 1.8755
R10 VTAIL VTAIL.n0 1.2311
R11 VTAIL VTAIL.n3 0.644897
R12 VDD1 VDD1.t1 106.049
R13 VDD1 VDD1.t0 65.4834
R14 B.n706 B.n705 585
R15 B.n292 B.n100 585
R16 B.n291 B.n290 585
R17 B.n289 B.n288 585
R18 B.n287 B.n286 585
R19 B.n285 B.n284 585
R20 B.n283 B.n282 585
R21 B.n281 B.n280 585
R22 B.n279 B.n278 585
R23 B.n277 B.n276 585
R24 B.n275 B.n274 585
R25 B.n273 B.n272 585
R26 B.n271 B.n270 585
R27 B.n269 B.n268 585
R28 B.n267 B.n266 585
R29 B.n265 B.n264 585
R30 B.n263 B.n262 585
R31 B.n261 B.n260 585
R32 B.n259 B.n258 585
R33 B.n257 B.n256 585
R34 B.n255 B.n254 585
R35 B.n253 B.n252 585
R36 B.n251 B.n250 585
R37 B.n249 B.n248 585
R38 B.n247 B.n246 585
R39 B.n245 B.n244 585
R40 B.n243 B.n242 585
R41 B.n241 B.n240 585
R42 B.n239 B.n238 585
R43 B.n237 B.n236 585
R44 B.n235 B.n234 585
R45 B.n233 B.n232 585
R46 B.n231 B.n230 585
R47 B.n229 B.n228 585
R48 B.n227 B.n226 585
R49 B.n225 B.n224 585
R50 B.n223 B.n222 585
R51 B.n221 B.n220 585
R52 B.n219 B.n218 585
R53 B.n217 B.n216 585
R54 B.n215 B.n214 585
R55 B.n213 B.n212 585
R56 B.n211 B.n210 585
R57 B.n208 B.n207 585
R58 B.n206 B.n205 585
R59 B.n204 B.n203 585
R60 B.n202 B.n201 585
R61 B.n200 B.n199 585
R62 B.n198 B.n197 585
R63 B.n196 B.n195 585
R64 B.n194 B.n193 585
R65 B.n192 B.n191 585
R66 B.n190 B.n189 585
R67 B.n187 B.n186 585
R68 B.n185 B.n184 585
R69 B.n183 B.n182 585
R70 B.n181 B.n180 585
R71 B.n179 B.n178 585
R72 B.n177 B.n176 585
R73 B.n175 B.n174 585
R74 B.n173 B.n172 585
R75 B.n171 B.n170 585
R76 B.n169 B.n168 585
R77 B.n167 B.n166 585
R78 B.n165 B.n164 585
R79 B.n163 B.n162 585
R80 B.n161 B.n160 585
R81 B.n159 B.n158 585
R82 B.n157 B.n156 585
R83 B.n155 B.n154 585
R84 B.n153 B.n152 585
R85 B.n151 B.n150 585
R86 B.n149 B.n148 585
R87 B.n147 B.n146 585
R88 B.n145 B.n144 585
R89 B.n143 B.n142 585
R90 B.n141 B.n140 585
R91 B.n139 B.n138 585
R92 B.n137 B.n136 585
R93 B.n135 B.n134 585
R94 B.n133 B.n132 585
R95 B.n131 B.n130 585
R96 B.n129 B.n128 585
R97 B.n127 B.n126 585
R98 B.n125 B.n124 585
R99 B.n123 B.n122 585
R100 B.n121 B.n120 585
R101 B.n119 B.n118 585
R102 B.n117 B.n116 585
R103 B.n115 B.n114 585
R104 B.n113 B.n112 585
R105 B.n111 B.n110 585
R106 B.n109 B.n108 585
R107 B.n107 B.n106 585
R108 B.n53 B.n52 585
R109 B.n711 B.n710 585
R110 B.n704 B.n101 585
R111 B.n101 B.n50 585
R112 B.n703 B.n49 585
R113 B.n715 B.n49 585
R114 B.n702 B.n48 585
R115 B.n716 B.n48 585
R116 B.n701 B.n47 585
R117 B.n717 B.n47 585
R118 B.n700 B.n699 585
R119 B.n699 B.n43 585
R120 B.n698 B.n42 585
R121 B.n723 B.n42 585
R122 B.n697 B.n41 585
R123 B.n724 B.n41 585
R124 B.n696 B.n40 585
R125 B.n725 B.n40 585
R126 B.n695 B.n694 585
R127 B.n694 B.n36 585
R128 B.n693 B.n35 585
R129 B.n731 B.n35 585
R130 B.n692 B.n34 585
R131 B.n732 B.n34 585
R132 B.n691 B.n33 585
R133 B.n733 B.n33 585
R134 B.n690 B.n689 585
R135 B.n689 B.n29 585
R136 B.n688 B.n28 585
R137 B.n739 B.n28 585
R138 B.n687 B.n27 585
R139 B.n740 B.n27 585
R140 B.n686 B.n26 585
R141 B.n741 B.n26 585
R142 B.n685 B.n684 585
R143 B.n684 B.n22 585
R144 B.n683 B.n21 585
R145 B.n747 B.n21 585
R146 B.n682 B.n20 585
R147 B.n748 B.n20 585
R148 B.n681 B.n19 585
R149 B.n749 B.n19 585
R150 B.n680 B.n679 585
R151 B.n679 B.n18 585
R152 B.n678 B.n14 585
R153 B.n755 B.n14 585
R154 B.n677 B.n13 585
R155 B.n756 B.n13 585
R156 B.n676 B.n12 585
R157 B.n757 B.n12 585
R158 B.n675 B.n674 585
R159 B.n674 B.n8 585
R160 B.n673 B.n7 585
R161 B.n763 B.n7 585
R162 B.n672 B.n6 585
R163 B.n764 B.n6 585
R164 B.n671 B.n5 585
R165 B.n765 B.n5 585
R166 B.n670 B.n669 585
R167 B.n669 B.n4 585
R168 B.n668 B.n293 585
R169 B.n668 B.n667 585
R170 B.n658 B.n294 585
R171 B.n295 B.n294 585
R172 B.n660 B.n659 585
R173 B.n661 B.n660 585
R174 B.n657 B.n300 585
R175 B.n300 B.n299 585
R176 B.n656 B.n655 585
R177 B.n655 B.n654 585
R178 B.n302 B.n301 585
R179 B.n647 B.n302 585
R180 B.n646 B.n645 585
R181 B.n648 B.n646 585
R182 B.n644 B.n307 585
R183 B.n307 B.n306 585
R184 B.n643 B.n642 585
R185 B.n642 B.n641 585
R186 B.n309 B.n308 585
R187 B.n310 B.n309 585
R188 B.n634 B.n633 585
R189 B.n635 B.n634 585
R190 B.n632 B.n315 585
R191 B.n315 B.n314 585
R192 B.n631 B.n630 585
R193 B.n630 B.n629 585
R194 B.n317 B.n316 585
R195 B.n318 B.n317 585
R196 B.n622 B.n621 585
R197 B.n623 B.n622 585
R198 B.n620 B.n323 585
R199 B.n323 B.n322 585
R200 B.n619 B.n618 585
R201 B.n618 B.n617 585
R202 B.n325 B.n324 585
R203 B.n326 B.n325 585
R204 B.n610 B.n609 585
R205 B.n611 B.n610 585
R206 B.n608 B.n331 585
R207 B.n331 B.n330 585
R208 B.n607 B.n606 585
R209 B.n606 B.n605 585
R210 B.n333 B.n332 585
R211 B.n334 B.n333 585
R212 B.n598 B.n597 585
R213 B.n599 B.n598 585
R214 B.n596 B.n339 585
R215 B.n339 B.n338 585
R216 B.n595 B.n594 585
R217 B.n594 B.n593 585
R218 B.n341 B.n340 585
R219 B.n342 B.n341 585
R220 B.n589 B.n588 585
R221 B.n345 B.n344 585
R222 B.n585 B.n584 585
R223 B.n586 B.n585 585
R224 B.n583 B.n393 585
R225 B.n582 B.n581 585
R226 B.n580 B.n579 585
R227 B.n578 B.n577 585
R228 B.n576 B.n575 585
R229 B.n574 B.n573 585
R230 B.n572 B.n571 585
R231 B.n570 B.n569 585
R232 B.n568 B.n567 585
R233 B.n566 B.n565 585
R234 B.n564 B.n563 585
R235 B.n562 B.n561 585
R236 B.n560 B.n559 585
R237 B.n558 B.n557 585
R238 B.n556 B.n555 585
R239 B.n554 B.n553 585
R240 B.n552 B.n551 585
R241 B.n550 B.n549 585
R242 B.n548 B.n547 585
R243 B.n546 B.n545 585
R244 B.n544 B.n543 585
R245 B.n542 B.n541 585
R246 B.n540 B.n539 585
R247 B.n538 B.n537 585
R248 B.n536 B.n535 585
R249 B.n534 B.n533 585
R250 B.n532 B.n531 585
R251 B.n530 B.n529 585
R252 B.n528 B.n527 585
R253 B.n526 B.n525 585
R254 B.n524 B.n523 585
R255 B.n522 B.n521 585
R256 B.n520 B.n519 585
R257 B.n518 B.n517 585
R258 B.n516 B.n515 585
R259 B.n514 B.n513 585
R260 B.n512 B.n511 585
R261 B.n510 B.n509 585
R262 B.n508 B.n507 585
R263 B.n506 B.n505 585
R264 B.n504 B.n503 585
R265 B.n502 B.n501 585
R266 B.n500 B.n499 585
R267 B.n498 B.n497 585
R268 B.n496 B.n495 585
R269 B.n494 B.n493 585
R270 B.n492 B.n491 585
R271 B.n490 B.n489 585
R272 B.n488 B.n487 585
R273 B.n486 B.n485 585
R274 B.n484 B.n483 585
R275 B.n482 B.n481 585
R276 B.n480 B.n479 585
R277 B.n478 B.n477 585
R278 B.n476 B.n475 585
R279 B.n474 B.n473 585
R280 B.n472 B.n471 585
R281 B.n470 B.n469 585
R282 B.n468 B.n467 585
R283 B.n466 B.n465 585
R284 B.n464 B.n463 585
R285 B.n462 B.n461 585
R286 B.n460 B.n459 585
R287 B.n458 B.n457 585
R288 B.n456 B.n455 585
R289 B.n454 B.n453 585
R290 B.n452 B.n451 585
R291 B.n450 B.n449 585
R292 B.n448 B.n447 585
R293 B.n446 B.n445 585
R294 B.n444 B.n443 585
R295 B.n442 B.n441 585
R296 B.n440 B.n439 585
R297 B.n438 B.n437 585
R298 B.n436 B.n435 585
R299 B.n434 B.n433 585
R300 B.n432 B.n431 585
R301 B.n430 B.n429 585
R302 B.n428 B.n427 585
R303 B.n426 B.n425 585
R304 B.n424 B.n423 585
R305 B.n422 B.n421 585
R306 B.n420 B.n419 585
R307 B.n418 B.n417 585
R308 B.n416 B.n415 585
R309 B.n414 B.n413 585
R310 B.n412 B.n411 585
R311 B.n410 B.n409 585
R312 B.n408 B.n407 585
R313 B.n406 B.n405 585
R314 B.n404 B.n403 585
R315 B.n402 B.n401 585
R316 B.n400 B.n392 585
R317 B.n586 B.n392 585
R318 B.n590 B.n343 585
R319 B.n343 B.n342 585
R320 B.n592 B.n591 585
R321 B.n593 B.n592 585
R322 B.n337 B.n336 585
R323 B.n338 B.n337 585
R324 B.n601 B.n600 585
R325 B.n600 B.n599 585
R326 B.n602 B.n335 585
R327 B.n335 B.n334 585
R328 B.n604 B.n603 585
R329 B.n605 B.n604 585
R330 B.n329 B.n328 585
R331 B.n330 B.n329 585
R332 B.n613 B.n612 585
R333 B.n612 B.n611 585
R334 B.n614 B.n327 585
R335 B.n327 B.n326 585
R336 B.n616 B.n615 585
R337 B.n617 B.n616 585
R338 B.n321 B.n320 585
R339 B.n322 B.n321 585
R340 B.n625 B.n624 585
R341 B.n624 B.n623 585
R342 B.n626 B.n319 585
R343 B.n319 B.n318 585
R344 B.n628 B.n627 585
R345 B.n629 B.n628 585
R346 B.n313 B.n312 585
R347 B.n314 B.n313 585
R348 B.n637 B.n636 585
R349 B.n636 B.n635 585
R350 B.n638 B.n311 585
R351 B.n311 B.n310 585
R352 B.n640 B.n639 585
R353 B.n641 B.n640 585
R354 B.n305 B.n304 585
R355 B.n306 B.n305 585
R356 B.n650 B.n649 585
R357 B.n649 B.n648 585
R358 B.n651 B.n303 585
R359 B.n647 B.n303 585
R360 B.n653 B.n652 585
R361 B.n654 B.n653 585
R362 B.n298 B.n297 585
R363 B.n299 B.n298 585
R364 B.n663 B.n662 585
R365 B.n662 B.n661 585
R366 B.n664 B.n296 585
R367 B.n296 B.n295 585
R368 B.n666 B.n665 585
R369 B.n667 B.n666 585
R370 B.n2 B.n0 585
R371 B.n4 B.n2 585
R372 B.n3 B.n1 585
R373 B.n764 B.n3 585
R374 B.n762 B.n761 585
R375 B.n763 B.n762 585
R376 B.n760 B.n9 585
R377 B.n9 B.n8 585
R378 B.n759 B.n758 585
R379 B.n758 B.n757 585
R380 B.n11 B.n10 585
R381 B.n756 B.n11 585
R382 B.n754 B.n753 585
R383 B.n755 B.n754 585
R384 B.n752 B.n15 585
R385 B.n18 B.n15 585
R386 B.n751 B.n750 585
R387 B.n750 B.n749 585
R388 B.n17 B.n16 585
R389 B.n748 B.n17 585
R390 B.n746 B.n745 585
R391 B.n747 B.n746 585
R392 B.n744 B.n23 585
R393 B.n23 B.n22 585
R394 B.n743 B.n742 585
R395 B.n742 B.n741 585
R396 B.n25 B.n24 585
R397 B.n740 B.n25 585
R398 B.n738 B.n737 585
R399 B.n739 B.n738 585
R400 B.n736 B.n30 585
R401 B.n30 B.n29 585
R402 B.n735 B.n734 585
R403 B.n734 B.n733 585
R404 B.n32 B.n31 585
R405 B.n732 B.n32 585
R406 B.n730 B.n729 585
R407 B.n731 B.n730 585
R408 B.n728 B.n37 585
R409 B.n37 B.n36 585
R410 B.n727 B.n726 585
R411 B.n726 B.n725 585
R412 B.n39 B.n38 585
R413 B.n724 B.n39 585
R414 B.n722 B.n721 585
R415 B.n723 B.n722 585
R416 B.n720 B.n44 585
R417 B.n44 B.n43 585
R418 B.n719 B.n718 585
R419 B.n718 B.n717 585
R420 B.n46 B.n45 585
R421 B.n716 B.n46 585
R422 B.n714 B.n713 585
R423 B.n715 B.n714 585
R424 B.n712 B.n51 585
R425 B.n51 B.n50 585
R426 B.n767 B.n766 585
R427 B.n766 B.n765 585
R428 B.n588 B.n343 550.159
R429 B.n710 B.n51 550.159
R430 B.n392 B.n341 550.159
R431 B.n706 B.n101 550.159
R432 B.n397 B.t10 311.724
R433 B.n394 B.t6 311.724
R434 B.n104 B.t13 311.724
R435 B.n102 B.t2 311.724
R436 B.n708 B.n707 256.663
R437 B.n708 B.n99 256.663
R438 B.n708 B.n98 256.663
R439 B.n708 B.n97 256.663
R440 B.n708 B.n96 256.663
R441 B.n708 B.n95 256.663
R442 B.n708 B.n94 256.663
R443 B.n708 B.n93 256.663
R444 B.n708 B.n92 256.663
R445 B.n708 B.n91 256.663
R446 B.n708 B.n90 256.663
R447 B.n708 B.n89 256.663
R448 B.n708 B.n88 256.663
R449 B.n708 B.n87 256.663
R450 B.n708 B.n86 256.663
R451 B.n708 B.n85 256.663
R452 B.n708 B.n84 256.663
R453 B.n708 B.n83 256.663
R454 B.n708 B.n82 256.663
R455 B.n708 B.n81 256.663
R456 B.n708 B.n80 256.663
R457 B.n708 B.n79 256.663
R458 B.n708 B.n78 256.663
R459 B.n708 B.n77 256.663
R460 B.n708 B.n76 256.663
R461 B.n708 B.n75 256.663
R462 B.n708 B.n74 256.663
R463 B.n708 B.n73 256.663
R464 B.n708 B.n72 256.663
R465 B.n708 B.n71 256.663
R466 B.n708 B.n70 256.663
R467 B.n708 B.n69 256.663
R468 B.n708 B.n68 256.663
R469 B.n708 B.n67 256.663
R470 B.n708 B.n66 256.663
R471 B.n708 B.n65 256.663
R472 B.n708 B.n64 256.663
R473 B.n708 B.n63 256.663
R474 B.n708 B.n62 256.663
R475 B.n708 B.n61 256.663
R476 B.n708 B.n60 256.663
R477 B.n708 B.n59 256.663
R478 B.n708 B.n58 256.663
R479 B.n708 B.n57 256.663
R480 B.n708 B.n56 256.663
R481 B.n708 B.n55 256.663
R482 B.n708 B.n54 256.663
R483 B.n709 B.n708 256.663
R484 B.n587 B.n586 256.663
R485 B.n586 B.n346 256.663
R486 B.n586 B.n347 256.663
R487 B.n586 B.n348 256.663
R488 B.n586 B.n349 256.663
R489 B.n586 B.n350 256.663
R490 B.n586 B.n351 256.663
R491 B.n586 B.n352 256.663
R492 B.n586 B.n353 256.663
R493 B.n586 B.n354 256.663
R494 B.n586 B.n355 256.663
R495 B.n586 B.n356 256.663
R496 B.n586 B.n357 256.663
R497 B.n586 B.n358 256.663
R498 B.n586 B.n359 256.663
R499 B.n586 B.n360 256.663
R500 B.n586 B.n361 256.663
R501 B.n586 B.n362 256.663
R502 B.n586 B.n363 256.663
R503 B.n586 B.n364 256.663
R504 B.n586 B.n365 256.663
R505 B.n586 B.n366 256.663
R506 B.n586 B.n367 256.663
R507 B.n586 B.n368 256.663
R508 B.n586 B.n369 256.663
R509 B.n586 B.n370 256.663
R510 B.n586 B.n371 256.663
R511 B.n586 B.n372 256.663
R512 B.n586 B.n373 256.663
R513 B.n586 B.n374 256.663
R514 B.n586 B.n375 256.663
R515 B.n586 B.n376 256.663
R516 B.n586 B.n377 256.663
R517 B.n586 B.n378 256.663
R518 B.n586 B.n379 256.663
R519 B.n586 B.n380 256.663
R520 B.n586 B.n381 256.663
R521 B.n586 B.n382 256.663
R522 B.n586 B.n383 256.663
R523 B.n586 B.n384 256.663
R524 B.n586 B.n385 256.663
R525 B.n586 B.n386 256.663
R526 B.n586 B.n387 256.663
R527 B.n586 B.n388 256.663
R528 B.n586 B.n389 256.663
R529 B.n586 B.n390 256.663
R530 B.n586 B.n391 256.663
R531 B.n592 B.n343 163.367
R532 B.n592 B.n337 163.367
R533 B.n600 B.n337 163.367
R534 B.n600 B.n335 163.367
R535 B.n604 B.n335 163.367
R536 B.n604 B.n329 163.367
R537 B.n612 B.n329 163.367
R538 B.n612 B.n327 163.367
R539 B.n616 B.n327 163.367
R540 B.n616 B.n321 163.367
R541 B.n624 B.n321 163.367
R542 B.n624 B.n319 163.367
R543 B.n628 B.n319 163.367
R544 B.n628 B.n313 163.367
R545 B.n636 B.n313 163.367
R546 B.n636 B.n311 163.367
R547 B.n640 B.n311 163.367
R548 B.n640 B.n305 163.367
R549 B.n649 B.n305 163.367
R550 B.n649 B.n303 163.367
R551 B.n653 B.n303 163.367
R552 B.n653 B.n298 163.367
R553 B.n662 B.n298 163.367
R554 B.n662 B.n296 163.367
R555 B.n666 B.n296 163.367
R556 B.n666 B.n2 163.367
R557 B.n766 B.n2 163.367
R558 B.n766 B.n3 163.367
R559 B.n762 B.n3 163.367
R560 B.n762 B.n9 163.367
R561 B.n758 B.n9 163.367
R562 B.n758 B.n11 163.367
R563 B.n754 B.n11 163.367
R564 B.n754 B.n15 163.367
R565 B.n750 B.n15 163.367
R566 B.n750 B.n17 163.367
R567 B.n746 B.n17 163.367
R568 B.n746 B.n23 163.367
R569 B.n742 B.n23 163.367
R570 B.n742 B.n25 163.367
R571 B.n738 B.n25 163.367
R572 B.n738 B.n30 163.367
R573 B.n734 B.n30 163.367
R574 B.n734 B.n32 163.367
R575 B.n730 B.n32 163.367
R576 B.n730 B.n37 163.367
R577 B.n726 B.n37 163.367
R578 B.n726 B.n39 163.367
R579 B.n722 B.n39 163.367
R580 B.n722 B.n44 163.367
R581 B.n718 B.n44 163.367
R582 B.n718 B.n46 163.367
R583 B.n714 B.n46 163.367
R584 B.n714 B.n51 163.367
R585 B.n585 B.n345 163.367
R586 B.n585 B.n393 163.367
R587 B.n581 B.n580 163.367
R588 B.n577 B.n576 163.367
R589 B.n573 B.n572 163.367
R590 B.n569 B.n568 163.367
R591 B.n565 B.n564 163.367
R592 B.n561 B.n560 163.367
R593 B.n557 B.n556 163.367
R594 B.n553 B.n552 163.367
R595 B.n549 B.n548 163.367
R596 B.n545 B.n544 163.367
R597 B.n541 B.n540 163.367
R598 B.n537 B.n536 163.367
R599 B.n533 B.n532 163.367
R600 B.n529 B.n528 163.367
R601 B.n525 B.n524 163.367
R602 B.n521 B.n520 163.367
R603 B.n517 B.n516 163.367
R604 B.n513 B.n512 163.367
R605 B.n509 B.n508 163.367
R606 B.n505 B.n504 163.367
R607 B.n501 B.n500 163.367
R608 B.n497 B.n496 163.367
R609 B.n493 B.n492 163.367
R610 B.n489 B.n488 163.367
R611 B.n485 B.n484 163.367
R612 B.n481 B.n480 163.367
R613 B.n477 B.n476 163.367
R614 B.n473 B.n472 163.367
R615 B.n469 B.n468 163.367
R616 B.n465 B.n464 163.367
R617 B.n461 B.n460 163.367
R618 B.n457 B.n456 163.367
R619 B.n453 B.n452 163.367
R620 B.n449 B.n448 163.367
R621 B.n445 B.n444 163.367
R622 B.n441 B.n440 163.367
R623 B.n437 B.n436 163.367
R624 B.n433 B.n432 163.367
R625 B.n429 B.n428 163.367
R626 B.n425 B.n424 163.367
R627 B.n421 B.n420 163.367
R628 B.n417 B.n416 163.367
R629 B.n413 B.n412 163.367
R630 B.n409 B.n408 163.367
R631 B.n405 B.n404 163.367
R632 B.n401 B.n392 163.367
R633 B.n594 B.n341 163.367
R634 B.n594 B.n339 163.367
R635 B.n598 B.n339 163.367
R636 B.n598 B.n333 163.367
R637 B.n606 B.n333 163.367
R638 B.n606 B.n331 163.367
R639 B.n610 B.n331 163.367
R640 B.n610 B.n325 163.367
R641 B.n618 B.n325 163.367
R642 B.n618 B.n323 163.367
R643 B.n622 B.n323 163.367
R644 B.n622 B.n317 163.367
R645 B.n630 B.n317 163.367
R646 B.n630 B.n315 163.367
R647 B.n634 B.n315 163.367
R648 B.n634 B.n309 163.367
R649 B.n642 B.n309 163.367
R650 B.n642 B.n307 163.367
R651 B.n646 B.n307 163.367
R652 B.n646 B.n302 163.367
R653 B.n655 B.n302 163.367
R654 B.n655 B.n300 163.367
R655 B.n660 B.n300 163.367
R656 B.n660 B.n294 163.367
R657 B.n668 B.n294 163.367
R658 B.n669 B.n668 163.367
R659 B.n669 B.n5 163.367
R660 B.n6 B.n5 163.367
R661 B.n7 B.n6 163.367
R662 B.n674 B.n7 163.367
R663 B.n674 B.n12 163.367
R664 B.n13 B.n12 163.367
R665 B.n14 B.n13 163.367
R666 B.n679 B.n14 163.367
R667 B.n679 B.n19 163.367
R668 B.n20 B.n19 163.367
R669 B.n21 B.n20 163.367
R670 B.n684 B.n21 163.367
R671 B.n684 B.n26 163.367
R672 B.n27 B.n26 163.367
R673 B.n28 B.n27 163.367
R674 B.n689 B.n28 163.367
R675 B.n689 B.n33 163.367
R676 B.n34 B.n33 163.367
R677 B.n35 B.n34 163.367
R678 B.n694 B.n35 163.367
R679 B.n694 B.n40 163.367
R680 B.n41 B.n40 163.367
R681 B.n42 B.n41 163.367
R682 B.n699 B.n42 163.367
R683 B.n699 B.n47 163.367
R684 B.n48 B.n47 163.367
R685 B.n49 B.n48 163.367
R686 B.n101 B.n49 163.367
R687 B.n106 B.n53 163.367
R688 B.n110 B.n109 163.367
R689 B.n114 B.n113 163.367
R690 B.n118 B.n117 163.367
R691 B.n122 B.n121 163.367
R692 B.n126 B.n125 163.367
R693 B.n130 B.n129 163.367
R694 B.n134 B.n133 163.367
R695 B.n138 B.n137 163.367
R696 B.n142 B.n141 163.367
R697 B.n146 B.n145 163.367
R698 B.n150 B.n149 163.367
R699 B.n154 B.n153 163.367
R700 B.n158 B.n157 163.367
R701 B.n162 B.n161 163.367
R702 B.n166 B.n165 163.367
R703 B.n170 B.n169 163.367
R704 B.n174 B.n173 163.367
R705 B.n178 B.n177 163.367
R706 B.n182 B.n181 163.367
R707 B.n186 B.n185 163.367
R708 B.n191 B.n190 163.367
R709 B.n195 B.n194 163.367
R710 B.n199 B.n198 163.367
R711 B.n203 B.n202 163.367
R712 B.n207 B.n206 163.367
R713 B.n212 B.n211 163.367
R714 B.n216 B.n215 163.367
R715 B.n220 B.n219 163.367
R716 B.n224 B.n223 163.367
R717 B.n228 B.n227 163.367
R718 B.n232 B.n231 163.367
R719 B.n236 B.n235 163.367
R720 B.n240 B.n239 163.367
R721 B.n244 B.n243 163.367
R722 B.n248 B.n247 163.367
R723 B.n252 B.n251 163.367
R724 B.n256 B.n255 163.367
R725 B.n260 B.n259 163.367
R726 B.n264 B.n263 163.367
R727 B.n268 B.n267 163.367
R728 B.n272 B.n271 163.367
R729 B.n276 B.n275 163.367
R730 B.n280 B.n279 163.367
R731 B.n284 B.n283 163.367
R732 B.n288 B.n287 163.367
R733 B.n290 B.n100 163.367
R734 B.n397 B.t12 136.954
R735 B.n102 B.t4 136.954
R736 B.n394 B.t9 136.939
R737 B.n104 B.t14 136.939
R738 B.n586 B.n342 88.2473
R739 B.n708 B.n50 88.2473
R740 B.n398 B.t11 73.7302
R741 B.n103 B.t5 73.7302
R742 B.n395 B.t8 73.7145
R743 B.n105 B.t15 73.7145
R744 B.n588 B.n587 71.676
R745 B.n393 B.n346 71.676
R746 B.n580 B.n347 71.676
R747 B.n576 B.n348 71.676
R748 B.n572 B.n349 71.676
R749 B.n568 B.n350 71.676
R750 B.n564 B.n351 71.676
R751 B.n560 B.n352 71.676
R752 B.n556 B.n353 71.676
R753 B.n552 B.n354 71.676
R754 B.n548 B.n355 71.676
R755 B.n544 B.n356 71.676
R756 B.n540 B.n357 71.676
R757 B.n536 B.n358 71.676
R758 B.n532 B.n359 71.676
R759 B.n528 B.n360 71.676
R760 B.n524 B.n361 71.676
R761 B.n520 B.n362 71.676
R762 B.n516 B.n363 71.676
R763 B.n512 B.n364 71.676
R764 B.n508 B.n365 71.676
R765 B.n504 B.n366 71.676
R766 B.n500 B.n367 71.676
R767 B.n496 B.n368 71.676
R768 B.n492 B.n369 71.676
R769 B.n488 B.n370 71.676
R770 B.n484 B.n371 71.676
R771 B.n480 B.n372 71.676
R772 B.n476 B.n373 71.676
R773 B.n472 B.n374 71.676
R774 B.n468 B.n375 71.676
R775 B.n464 B.n376 71.676
R776 B.n460 B.n377 71.676
R777 B.n456 B.n378 71.676
R778 B.n452 B.n379 71.676
R779 B.n448 B.n380 71.676
R780 B.n444 B.n381 71.676
R781 B.n440 B.n382 71.676
R782 B.n436 B.n383 71.676
R783 B.n432 B.n384 71.676
R784 B.n428 B.n385 71.676
R785 B.n424 B.n386 71.676
R786 B.n420 B.n387 71.676
R787 B.n416 B.n388 71.676
R788 B.n412 B.n389 71.676
R789 B.n408 B.n390 71.676
R790 B.n404 B.n391 71.676
R791 B.n710 B.n709 71.676
R792 B.n106 B.n54 71.676
R793 B.n110 B.n55 71.676
R794 B.n114 B.n56 71.676
R795 B.n118 B.n57 71.676
R796 B.n122 B.n58 71.676
R797 B.n126 B.n59 71.676
R798 B.n130 B.n60 71.676
R799 B.n134 B.n61 71.676
R800 B.n138 B.n62 71.676
R801 B.n142 B.n63 71.676
R802 B.n146 B.n64 71.676
R803 B.n150 B.n65 71.676
R804 B.n154 B.n66 71.676
R805 B.n158 B.n67 71.676
R806 B.n162 B.n68 71.676
R807 B.n166 B.n69 71.676
R808 B.n170 B.n70 71.676
R809 B.n174 B.n71 71.676
R810 B.n178 B.n72 71.676
R811 B.n182 B.n73 71.676
R812 B.n186 B.n74 71.676
R813 B.n191 B.n75 71.676
R814 B.n195 B.n76 71.676
R815 B.n199 B.n77 71.676
R816 B.n203 B.n78 71.676
R817 B.n207 B.n79 71.676
R818 B.n212 B.n80 71.676
R819 B.n216 B.n81 71.676
R820 B.n220 B.n82 71.676
R821 B.n224 B.n83 71.676
R822 B.n228 B.n84 71.676
R823 B.n232 B.n85 71.676
R824 B.n236 B.n86 71.676
R825 B.n240 B.n87 71.676
R826 B.n244 B.n88 71.676
R827 B.n248 B.n89 71.676
R828 B.n252 B.n90 71.676
R829 B.n256 B.n91 71.676
R830 B.n260 B.n92 71.676
R831 B.n264 B.n93 71.676
R832 B.n268 B.n94 71.676
R833 B.n272 B.n95 71.676
R834 B.n276 B.n96 71.676
R835 B.n280 B.n97 71.676
R836 B.n284 B.n98 71.676
R837 B.n288 B.n99 71.676
R838 B.n707 B.n100 71.676
R839 B.n707 B.n706 71.676
R840 B.n290 B.n99 71.676
R841 B.n287 B.n98 71.676
R842 B.n283 B.n97 71.676
R843 B.n279 B.n96 71.676
R844 B.n275 B.n95 71.676
R845 B.n271 B.n94 71.676
R846 B.n267 B.n93 71.676
R847 B.n263 B.n92 71.676
R848 B.n259 B.n91 71.676
R849 B.n255 B.n90 71.676
R850 B.n251 B.n89 71.676
R851 B.n247 B.n88 71.676
R852 B.n243 B.n87 71.676
R853 B.n239 B.n86 71.676
R854 B.n235 B.n85 71.676
R855 B.n231 B.n84 71.676
R856 B.n227 B.n83 71.676
R857 B.n223 B.n82 71.676
R858 B.n219 B.n81 71.676
R859 B.n215 B.n80 71.676
R860 B.n211 B.n79 71.676
R861 B.n206 B.n78 71.676
R862 B.n202 B.n77 71.676
R863 B.n198 B.n76 71.676
R864 B.n194 B.n75 71.676
R865 B.n190 B.n74 71.676
R866 B.n185 B.n73 71.676
R867 B.n181 B.n72 71.676
R868 B.n177 B.n71 71.676
R869 B.n173 B.n70 71.676
R870 B.n169 B.n69 71.676
R871 B.n165 B.n68 71.676
R872 B.n161 B.n67 71.676
R873 B.n157 B.n66 71.676
R874 B.n153 B.n65 71.676
R875 B.n149 B.n64 71.676
R876 B.n145 B.n63 71.676
R877 B.n141 B.n62 71.676
R878 B.n137 B.n61 71.676
R879 B.n133 B.n60 71.676
R880 B.n129 B.n59 71.676
R881 B.n125 B.n58 71.676
R882 B.n121 B.n57 71.676
R883 B.n117 B.n56 71.676
R884 B.n113 B.n55 71.676
R885 B.n109 B.n54 71.676
R886 B.n709 B.n53 71.676
R887 B.n587 B.n345 71.676
R888 B.n581 B.n346 71.676
R889 B.n577 B.n347 71.676
R890 B.n573 B.n348 71.676
R891 B.n569 B.n349 71.676
R892 B.n565 B.n350 71.676
R893 B.n561 B.n351 71.676
R894 B.n557 B.n352 71.676
R895 B.n553 B.n353 71.676
R896 B.n549 B.n354 71.676
R897 B.n545 B.n355 71.676
R898 B.n541 B.n356 71.676
R899 B.n537 B.n357 71.676
R900 B.n533 B.n358 71.676
R901 B.n529 B.n359 71.676
R902 B.n525 B.n360 71.676
R903 B.n521 B.n361 71.676
R904 B.n517 B.n362 71.676
R905 B.n513 B.n363 71.676
R906 B.n509 B.n364 71.676
R907 B.n505 B.n365 71.676
R908 B.n501 B.n366 71.676
R909 B.n497 B.n367 71.676
R910 B.n493 B.n368 71.676
R911 B.n489 B.n369 71.676
R912 B.n485 B.n370 71.676
R913 B.n481 B.n371 71.676
R914 B.n477 B.n372 71.676
R915 B.n473 B.n373 71.676
R916 B.n469 B.n374 71.676
R917 B.n465 B.n375 71.676
R918 B.n461 B.n376 71.676
R919 B.n457 B.n377 71.676
R920 B.n453 B.n378 71.676
R921 B.n449 B.n379 71.676
R922 B.n445 B.n380 71.676
R923 B.n441 B.n381 71.676
R924 B.n437 B.n382 71.676
R925 B.n433 B.n383 71.676
R926 B.n429 B.n384 71.676
R927 B.n425 B.n385 71.676
R928 B.n421 B.n386 71.676
R929 B.n417 B.n387 71.676
R930 B.n413 B.n388 71.676
R931 B.n409 B.n389 71.676
R932 B.n405 B.n390 71.676
R933 B.n401 B.n391 71.676
R934 B.n398 B.n397 63.2247
R935 B.n395 B.n394 63.2247
R936 B.n105 B.n104 63.2247
R937 B.n103 B.n102 63.2247
R938 B.n399 B.n398 59.5399
R939 B.n396 B.n395 59.5399
R940 B.n188 B.n105 59.5399
R941 B.n209 B.n103 59.5399
R942 B.n593 B.n342 41.964
R943 B.n593 B.n338 41.964
R944 B.n599 B.n338 41.964
R945 B.n599 B.n334 41.964
R946 B.n605 B.n334 41.964
R947 B.n605 B.n330 41.964
R948 B.n611 B.n330 41.964
R949 B.n617 B.n326 41.964
R950 B.n617 B.n322 41.964
R951 B.n623 B.n322 41.964
R952 B.n623 B.n318 41.964
R953 B.n629 B.n318 41.964
R954 B.n629 B.n314 41.964
R955 B.n635 B.n314 41.964
R956 B.n635 B.n310 41.964
R957 B.n641 B.n310 41.964
R958 B.n641 B.n306 41.964
R959 B.n648 B.n306 41.964
R960 B.n648 B.n647 41.964
R961 B.n654 B.n299 41.964
R962 B.n661 B.n299 41.964
R963 B.n661 B.n295 41.964
R964 B.n667 B.n295 41.964
R965 B.n667 B.n4 41.964
R966 B.n765 B.n4 41.964
R967 B.n765 B.n764 41.964
R968 B.n764 B.n763 41.964
R969 B.n763 B.n8 41.964
R970 B.n757 B.n8 41.964
R971 B.n757 B.n756 41.964
R972 B.n756 B.n755 41.964
R973 B.n749 B.n18 41.964
R974 B.n749 B.n748 41.964
R975 B.n748 B.n747 41.964
R976 B.n747 B.n22 41.964
R977 B.n741 B.n22 41.964
R978 B.n741 B.n740 41.964
R979 B.n740 B.n739 41.964
R980 B.n739 B.n29 41.964
R981 B.n733 B.n29 41.964
R982 B.n733 B.n732 41.964
R983 B.n732 B.n731 41.964
R984 B.n731 B.n36 41.964
R985 B.n725 B.n724 41.964
R986 B.n724 B.n723 41.964
R987 B.n723 B.n43 41.964
R988 B.n717 B.n43 41.964
R989 B.n717 B.n716 41.964
R990 B.n716 B.n715 41.964
R991 B.n715 B.n50 41.964
R992 B.n712 B.n711 35.7468
R993 B.n705 B.n704 35.7468
R994 B.n400 B.n340 35.7468
R995 B.n590 B.n589 35.7468
R996 B.n611 B.t7 33.9416
R997 B.n725 B.t3 33.9416
R998 B.n647 B.t0 25.302
R999 B.n18 B.t1 25.302
R1000 B B.n767 18.0485
R1001 B.n654 B.t0 16.6625
R1002 B.n755 B.t1 16.6625
R1003 B.n711 B.n52 10.6151
R1004 B.n107 B.n52 10.6151
R1005 B.n108 B.n107 10.6151
R1006 B.n111 B.n108 10.6151
R1007 B.n112 B.n111 10.6151
R1008 B.n115 B.n112 10.6151
R1009 B.n116 B.n115 10.6151
R1010 B.n119 B.n116 10.6151
R1011 B.n120 B.n119 10.6151
R1012 B.n123 B.n120 10.6151
R1013 B.n124 B.n123 10.6151
R1014 B.n127 B.n124 10.6151
R1015 B.n128 B.n127 10.6151
R1016 B.n131 B.n128 10.6151
R1017 B.n132 B.n131 10.6151
R1018 B.n135 B.n132 10.6151
R1019 B.n136 B.n135 10.6151
R1020 B.n139 B.n136 10.6151
R1021 B.n140 B.n139 10.6151
R1022 B.n143 B.n140 10.6151
R1023 B.n144 B.n143 10.6151
R1024 B.n147 B.n144 10.6151
R1025 B.n148 B.n147 10.6151
R1026 B.n151 B.n148 10.6151
R1027 B.n152 B.n151 10.6151
R1028 B.n155 B.n152 10.6151
R1029 B.n156 B.n155 10.6151
R1030 B.n159 B.n156 10.6151
R1031 B.n160 B.n159 10.6151
R1032 B.n163 B.n160 10.6151
R1033 B.n164 B.n163 10.6151
R1034 B.n167 B.n164 10.6151
R1035 B.n168 B.n167 10.6151
R1036 B.n171 B.n168 10.6151
R1037 B.n172 B.n171 10.6151
R1038 B.n175 B.n172 10.6151
R1039 B.n176 B.n175 10.6151
R1040 B.n179 B.n176 10.6151
R1041 B.n180 B.n179 10.6151
R1042 B.n183 B.n180 10.6151
R1043 B.n184 B.n183 10.6151
R1044 B.n187 B.n184 10.6151
R1045 B.n192 B.n189 10.6151
R1046 B.n193 B.n192 10.6151
R1047 B.n196 B.n193 10.6151
R1048 B.n197 B.n196 10.6151
R1049 B.n200 B.n197 10.6151
R1050 B.n201 B.n200 10.6151
R1051 B.n204 B.n201 10.6151
R1052 B.n205 B.n204 10.6151
R1053 B.n208 B.n205 10.6151
R1054 B.n213 B.n210 10.6151
R1055 B.n214 B.n213 10.6151
R1056 B.n217 B.n214 10.6151
R1057 B.n218 B.n217 10.6151
R1058 B.n221 B.n218 10.6151
R1059 B.n222 B.n221 10.6151
R1060 B.n225 B.n222 10.6151
R1061 B.n226 B.n225 10.6151
R1062 B.n229 B.n226 10.6151
R1063 B.n230 B.n229 10.6151
R1064 B.n233 B.n230 10.6151
R1065 B.n234 B.n233 10.6151
R1066 B.n237 B.n234 10.6151
R1067 B.n238 B.n237 10.6151
R1068 B.n241 B.n238 10.6151
R1069 B.n242 B.n241 10.6151
R1070 B.n245 B.n242 10.6151
R1071 B.n246 B.n245 10.6151
R1072 B.n249 B.n246 10.6151
R1073 B.n250 B.n249 10.6151
R1074 B.n253 B.n250 10.6151
R1075 B.n254 B.n253 10.6151
R1076 B.n257 B.n254 10.6151
R1077 B.n258 B.n257 10.6151
R1078 B.n261 B.n258 10.6151
R1079 B.n262 B.n261 10.6151
R1080 B.n265 B.n262 10.6151
R1081 B.n266 B.n265 10.6151
R1082 B.n269 B.n266 10.6151
R1083 B.n270 B.n269 10.6151
R1084 B.n273 B.n270 10.6151
R1085 B.n274 B.n273 10.6151
R1086 B.n277 B.n274 10.6151
R1087 B.n278 B.n277 10.6151
R1088 B.n281 B.n278 10.6151
R1089 B.n282 B.n281 10.6151
R1090 B.n285 B.n282 10.6151
R1091 B.n286 B.n285 10.6151
R1092 B.n289 B.n286 10.6151
R1093 B.n291 B.n289 10.6151
R1094 B.n292 B.n291 10.6151
R1095 B.n705 B.n292 10.6151
R1096 B.n595 B.n340 10.6151
R1097 B.n596 B.n595 10.6151
R1098 B.n597 B.n596 10.6151
R1099 B.n597 B.n332 10.6151
R1100 B.n607 B.n332 10.6151
R1101 B.n608 B.n607 10.6151
R1102 B.n609 B.n608 10.6151
R1103 B.n609 B.n324 10.6151
R1104 B.n619 B.n324 10.6151
R1105 B.n620 B.n619 10.6151
R1106 B.n621 B.n620 10.6151
R1107 B.n621 B.n316 10.6151
R1108 B.n631 B.n316 10.6151
R1109 B.n632 B.n631 10.6151
R1110 B.n633 B.n632 10.6151
R1111 B.n633 B.n308 10.6151
R1112 B.n643 B.n308 10.6151
R1113 B.n644 B.n643 10.6151
R1114 B.n645 B.n644 10.6151
R1115 B.n645 B.n301 10.6151
R1116 B.n656 B.n301 10.6151
R1117 B.n657 B.n656 10.6151
R1118 B.n659 B.n657 10.6151
R1119 B.n659 B.n658 10.6151
R1120 B.n658 B.n293 10.6151
R1121 B.n670 B.n293 10.6151
R1122 B.n671 B.n670 10.6151
R1123 B.n672 B.n671 10.6151
R1124 B.n673 B.n672 10.6151
R1125 B.n675 B.n673 10.6151
R1126 B.n676 B.n675 10.6151
R1127 B.n677 B.n676 10.6151
R1128 B.n678 B.n677 10.6151
R1129 B.n680 B.n678 10.6151
R1130 B.n681 B.n680 10.6151
R1131 B.n682 B.n681 10.6151
R1132 B.n683 B.n682 10.6151
R1133 B.n685 B.n683 10.6151
R1134 B.n686 B.n685 10.6151
R1135 B.n687 B.n686 10.6151
R1136 B.n688 B.n687 10.6151
R1137 B.n690 B.n688 10.6151
R1138 B.n691 B.n690 10.6151
R1139 B.n692 B.n691 10.6151
R1140 B.n693 B.n692 10.6151
R1141 B.n695 B.n693 10.6151
R1142 B.n696 B.n695 10.6151
R1143 B.n697 B.n696 10.6151
R1144 B.n698 B.n697 10.6151
R1145 B.n700 B.n698 10.6151
R1146 B.n701 B.n700 10.6151
R1147 B.n702 B.n701 10.6151
R1148 B.n703 B.n702 10.6151
R1149 B.n704 B.n703 10.6151
R1150 B.n589 B.n344 10.6151
R1151 B.n584 B.n344 10.6151
R1152 B.n584 B.n583 10.6151
R1153 B.n583 B.n582 10.6151
R1154 B.n582 B.n579 10.6151
R1155 B.n579 B.n578 10.6151
R1156 B.n578 B.n575 10.6151
R1157 B.n575 B.n574 10.6151
R1158 B.n574 B.n571 10.6151
R1159 B.n571 B.n570 10.6151
R1160 B.n570 B.n567 10.6151
R1161 B.n567 B.n566 10.6151
R1162 B.n566 B.n563 10.6151
R1163 B.n563 B.n562 10.6151
R1164 B.n562 B.n559 10.6151
R1165 B.n559 B.n558 10.6151
R1166 B.n558 B.n555 10.6151
R1167 B.n555 B.n554 10.6151
R1168 B.n554 B.n551 10.6151
R1169 B.n551 B.n550 10.6151
R1170 B.n550 B.n547 10.6151
R1171 B.n547 B.n546 10.6151
R1172 B.n546 B.n543 10.6151
R1173 B.n543 B.n542 10.6151
R1174 B.n542 B.n539 10.6151
R1175 B.n539 B.n538 10.6151
R1176 B.n538 B.n535 10.6151
R1177 B.n535 B.n534 10.6151
R1178 B.n534 B.n531 10.6151
R1179 B.n531 B.n530 10.6151
R1180 B.n530 B.n527 10.6151
R1181 B.n527 B.n526 10.6151
R1182 B.n526 B.n523 10.6151
R1183 B.n523 B.n522 10.6151
R1184 B.n522 B.n519 10.6151
R1185 B.n519 B.n518 10.6151
R1186 B.n518 B.n515 10.6151
R1187 B.n515 B.n514 10.6151
R1188 B.n514 B.n511 10.6151
R1189 B.n511 B.n510 10.6151
R1190 B.n510 B.n507 10.6151
R1191 B.n507 B.n506 10.6151
R1192 B.n503 B.n502 10.6151
R1193 B.n502 B.n499 10.6151
R1194 B.n499 B.n498 10.6151
R1195 B.n498 B.n495 10.6151
R1196 B.n495 B.n494 10.6151
R1197 B.n494 B.n491 10.6151
R1198 B.n491 B.n490 10.6151
R1199 B.n490 B.n487 10.6151
R1200 B.n487 B.n486 10.6151
R1201 B.n483 B.n482 10.6151
R1202 B.n482 B.n479 10.6151
R1203 B.n479 B.n478 10.6151
R1204 B.n478 B.n475 10.6151
R1205 B.n475 B.n474 10.6151
R1206 B.n474 B.n471 10.6151
R1207 B.n471 B.n470 10.6151
R1208 B.n470 B.n467 10.6151
R1209 B.n467 B.n466 10.6151
R1210 B.n466 B.n463 10.6151
R1211 B.n463 B.n462 10.6151
R1212 B.n462 B.n459 10.6151
R1213 B.n459 B.n458 10.6151
R1214 B.n458 B.n455 10.6151
R1215 B.n455 B.n454 10.6151
R1216 B.n454 B.n451 10.6151
R1217 B.n451 B.n450 10.6151
R1218 B.n450 B.n447 10.6151
R1219 B.n447 B.n446 10.6151
R1220 B.n446 B.n443 10.6151
R1221 B.n443 B.n442 10.6151
R1222 B.n442 B.n439 10.6151
R1223 B.n439 B.n438 10.6151
R1224 B.n438 B.n435 10.6151
R1225 B.n435 B.n434 10.6151
R1226 B.n434 B.n431 10.6151
R1227 B.n431 B.n430 10.6151
R1228 B.n430 B.n427 10.6151
R1229 B.n427 B.n426 10.6151
R1230 B.n426 B.n423 10.6151
R1231 B.n423 B.n422 10.6151
R1232 B.n422 B.n419 10.6151
R1233 B.n419 B.n418 10.6151
R1234 B.n418 B.n415 10.6151
R1235 B.n415 B.n414 10.6151
R1236 B.n414 B.n411 10.6151
R1237 B.n411 B.n410 10.6151
R1238 B.n410 B.n407 10.6151
R1239 B.n407 B.n406 10.6151
R1240 B.n406 B.n403 10.6151
R1241 B.n403 B.n402 10.6151
R1242 B.n402 B.n400 10.6151
R1243 B.n591 B.n590 10.6151
R1244 B.n591 B.n336 10.6151
R1245 B.n601 B.n336 10.6151
R1246 B.n602 B.n601 10.6151
R1247 B.n603 B.n602 10.6151
R1248 B.n603 B.n328 10.6151
R1249 B.n613 B.n328 10.6151
R1250 B.n614 B.n613 10.6151
R1251 B.n615 B.n614 10.6151
R1252 B.n615 B.n320 10.6151
R1253 B.n625 B.n320 10.6151
R1254 B.n626 B.n625 10.6151
R1255 B.n627 B.n626 10.6151
R1256 B.n627 B.n312 10.6151
R1257 B.n637 B.n312 10.6151
R1258 B.n638 B.n637 10.6151
R1259 B.n639 B.n638 10.6151
R1260 B.n639 B.n304 10.6151
R1261 B.n650 B.n304 10.6151
R1262 B.n651 B.n650 10.6151
R1263 B.n652 B.n651 10.6151
R1264 B.n652 B.n297 10.6151
R1265 B.n663 B.n297 10.6151
R1266 B.n664 B.n663 10.6151
R1267 B.n665 B.n664 10.6151
R1268 B.n665 B.n0 10.6151
R1269 B.n761 B.n1 10.6151
R1270 B.n761 B.n760 10.6151
R1271 B.n760 B.n759 10.6151
R1272 B.n759 B.n10 10.6151
R1273 B.n753 B.n10 10.6151
R1274 B.n753 B.n752 10.6151
R1275 B.n752 B.n751 10.6151
R1276 B.n751 B.n16 10.6151
R1277 B.n745 B.n16 10.6151
R1278 B.n745 B.n744 10.6151
R1279 B.n744 B.n743 10.6151
R1280 B.n743 B.n24 10.6151
R1281 B.n737 B.n24 10.6151
R1282 B.n737 B.n736 10.6151
R1283 B.n736 B.n735 10.6151
R1284 B.n735 B.n31 10.6151
R1285 B.n729 B.n31 10.6151
R1286 B.n729 B.n728 10.6151
R1287 B.n728 B.n727 10.6151
R1288 B.n727 B.n38 10.6151
R1289 B.n721 B.n38 10.6151
R1290 B.n721 B.n720 10.6151
R1291 B.n720 B.n719 10.6151
R1292 B.n719 B.n45 10.6151
R1293 B.n713 B.n45 10.6151
R1294 B.n713 B.n712 10.6151
R1295 B.n188 B.n187 9.36635
R1296 B.n210 B.n209 9.36635
R1297 B.n506 B.n396 9.36635
R1298 B.n483 B.n399 9.36635
R1299 B.t7 B.n326 8.02294
R1300 B.t3 B.n36 8.02294
R1301 B.n767 B.n0 2.81026
R1302 B.n767 B.n1 2.81026
R1303 B.n189 B.n188 1.24928
R1304 B.n209 B.n208 1.24928
R1305 B.n503 B.n396 1.24928
R1306 B.n486 B.n399 1.24928
R1307 VN VN.t1 190.274
R1308 VN VN.t0 144.755
R1309 VDD2.n0 VDD2.t1 104.822
R1310 VDD2.n0 VDD2.t0 64.7226
R1311 VDD2 VDD2.n0 0.761276
C0 VN VTAIL 2.61599f
C1 VDD2 VP 0.346963f
C2 VN VDD1 0.148273f
C3 VDD1 VTAIL 5.26183f
C4 VN VP 5.71197f
C5 VN VDD2 2.94683f
C6 VTAIL VP 2.63026f
C7 VTAIL VDD2 5.31487f
C8 VDD1 VP 3.14306f
C9 VDD1 VDD2 0.714655f
C10 VDD2 B 4.643315f
C11 VDD1 B 7.880229f
C12 VTAIL B 7.748884f
C13 VN B 11.124599f
C14 VP B 6.843712f
C15 VDD2.t1 B 2.83935f
C16 VDD2.t0 B 2.27545f
C17 VDD2.n0 B 2.94426f
C18 VN.t0 B 3.19332f
C19 VN.t1 B 3.76639f
C20 VDD1.t0 B 2.31327f
C21 VDD1.t1 B 2.92134f
C22 VTAIL.t3 B 2.26694f
C23 VTAIL.n0 B 1.73384f
C24 VTAIL.t0 B 2.26696f
C25 VTAIL.n1 B 1.77684f
C26 VTAIL.t2 B 2.26694f
C27 VTAIL.n2 B 1.58926f
C28 VTAIL.t1 B 2.26694f
C29 VTAIL.n3 B 1.50711f
C30 VP.t0 B 3.25888f
C31 VP.t1 B 3.84565f
C32 VP.n0 B 4.21121f
.ends

