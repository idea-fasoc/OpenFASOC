* NGSPICE file created from diff_pair_sample_1036.ext - technology: sky130A

.subckt diff_pair_sample_1036 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t11 VN.t0 VDD2.t2 w_n4218_n3882# sky130_fd_pr__pfet_01v8 ad=2.40405 pd=14.9 as=2.40405 ps=14.9 w=14.57 l=3.73
X1 VDD2.t3 VN.t1 VTAIL.t10 w_n4218_n3882# sky130_fd_pr__pfet_01v8 ad=5.6823 pd=29.92 as=2.40405 ps=14.9 w=14.57 l=3.73
X2 B.t11 B.t9 B.t10 w_n4218_n3882# sky130_fd_pr__pfet_01v8 ad=5.6823 pd=29.92 as=0 ps=0 w=14.57 l=3.73
X3 B.t8 B.t6 B.t7 w_n4218_n3882# sky130_fd_pr__pfet_01v8 ad=5.6823 pd=29.92 as=0 ps=0 w=14.57 l=3.73
X4 VDD1.t5 VP.t0 VTAIL.t2 w_n4218_n3882# sky130_fd_pr__pfet_01v8 ad=5.6823 pd=29.92 as=2.40405 ps=14.9 w=14.57 l=3.73
X5 VDD1.t4 VP.t1 VTAIL.t0 w_n4218_n3882# sky130_fd_pr__pfet_01v8 ad=2.40405 pd=14.9 as=5.6823 ps=29.92 w=14.57 l=3.73
X6 VDD2.t5 VN.t2 VTAIL.t9 w_n4218_n3882# sky130_fd_pr__pfet_01v8 ad=2.40405 pd=14.9 as=5.6823 ps=29.92 w=14.57 l=3.73
X7 B.t5 B.t3 B.t4 w_n4218_n3882# sky130_fd_pr__pfet_01v8 ad=5.6823 pd=29.92 as=0 ps=0 w=14.57 l=3.73
X8 VDD1.t3 VP.t2 VTAIL.t1 w_n4218_n3882# sky130_fd_pr__pfet_01v8 ad=2.40405 pd=14.9 as=5.6823 ps=29.92 w=14.57 l=3.73
X9 VTAIL.t8 VN.t3 VDD2.t4 w_n4218_n3882# sky130_fd_pr__pfet_01v8 ad=2.40405 pd=14.9 as=2.40405 ps=14.9 w=14.57 l=3.73
X10 VTAIL.t4 VP.t3 VDD1.t2 w_n4218_n3882# sky130_fd_pr__pfet_01v8 ad=2.40405 pd=14.9 as=2.40405 ps=14.9 w=14.57 l=3.73
X11 VTAIL.t3 VP.t4 VDD1.t1 w_n4218_n3882# sky130_fd_pr__pfet_01v8 ad=2.40405 pd=14.9 as=2.40405 ps=14.9 w=14.57 l=3.73
X12 VDD2.t1 VN.t4 VTAIL.t7 w_n4218_n3882# sky130_fd_pr__pfet_01v8 ad=5.6823 pd=29.92 as=2.40405 ps=14.9 w=14.57 l=3.73
X13 B.t2 B.t0 B.t1 w_n4218_n3882# sky130_fd_pr__pfet_01v8 ad=5.6823 pd=29.92 as=0 ps=0 w=14.57 l=3.73
X14 VDD1.t0 VP.t5 VTAIL.t5 w_n4218_n3882# sky130_fd_pr__pfet_01v8 ad=5.6823 pd=29.92 as=2.40405 ps=14.9 w=14.57 l=3.73
X15 VDD2.t0 VN.t5 VTAIL.t6 w_n4218_n3882# sky130_fd_pr__pfet_01v8 ad=2.40405 pd=14.9 as=5.6823 ps=29.92 w=14.57 l=3.73
R0 VN.n38 VN.n37 161.3
R1 VN.n36 VN.n21 161.3
R2 VN.n35 VN.n34 161.3
R3 VN.n33 VN.n22 161.3
R4 VN.n32 VN.n31 161.3
R5 VN.n30 VN.n23 161.3
R6 VN.n29 VN.n28 161.3
R7 VN.n27 VN.n24 161.3
R8 VN.n18 VN.n17 161.3
R9 VN.n16 VN.n1 161.3
R10 VN.n15 VN.n14 161.3
R11 VN.n13 VN.n2 161.3
R12 VN.n12 VN.n11 161.3
R13 VN.n10 VN.n3 161.3
R14 VN.n9 VN.n8 161.3
R15 VN.n7 VN.n4 161.3
R16 VN.n26 VN.t2 127.058
R17 VN.n6 VN.t1 127.058
R18 VN.n5 VN.t3 94.1391
R19 VN.n0 VN.t5 94.1391
R20 VN.n25 VN.t0 94.1391
R21 VN.n20 VN.t4 94.1391
R22 VN.n19 VN.n0 87.1314
R23 VN.n39 VN.n20 87.1314
R24 VN VN.n39 55.2556
R25 VN.n6 VN.n5 50.484
R26 VN.n26 VN.n25 50.484
R27 VN.n11 VN.n2 43.4072
R28 VN.n31 VN.n22 43.4072
R29 VN.n11 VN.n10 37.5796
R30 VN.n31 VN.n30 37.5796
R31 VN.n5 VN.n4 24.4675
R32 VN.n9 VN.n4 24.4675
R33 VN.n10 VN.n9 24.4675
R34 VN.n15 VN.n2 24.4675
R35 VN.n16 VN.n15 24.4675
R36 VN.n17 VN.n16 24.4675
R37 VN.n30 VN.n29 24.4675
R38 VN.n29 VN.n24 24.4675
R39 VN.n25 VN.n24 24.4675
R40 VN.n37 VN.n36 24.4675
R41 VN.n36 VN.n35 24.4675
R42 VN.n35 VN.n22 24.4675
R43 VN.n17 VN.n0 2.93654
R44 VN.n37 VN.n20 2.93654
R45 VN.n27 VN.n26 2.46264
R46 VN.n7 VN.n6 2.46264
R47 VN.n39 VN.n38 0.354971
R48 VN.n19 VN.n18 0.354971
R49 VN VN.n19 0.26696
R50 VN.n38 VN.n21 0.189894
R51 VN.n34 VN.n21 0.189894
R52 VN.n34 VN.n33 0.189894
R53 VN.n33 VN.n32 0.189894
R54 VN.n32 VN.n23 0.189894
R55 VN.n28 VN.n23 0.189894
R56 VN.n28 VN.n27 0.189894
R57 VN.n8 VN.n7 0.189894
R58 VN.n8 VN.n3 0.189894
R59 VN.n12 VN.n3 0.189894
R60 VN.n13 VN.n12 0.189894
R61 VN.n14 VN.n13 0.189894
R62 VN.n14 VN.n1 0.189894
R63 VN.n18 VN.n1 0.189894
R64 VDD2.n1 VDD2.t3 74.7787
R65 VDD2.n2 VDD2.t1 72.2093
R66 VDD2.n1 VDD2.n0 70.798
R67 VDD2 VDD2.n3 70.7952
R68 VDD2.n2 VDD2.n1 47.6506
R69 VDD2 VDD2.n2 2.68369
R70 VDD2.n3 VDD2.t2 2.23145
R71 VDD2.n3 VDD2.t5 2.23145
R72 VDD2.n0 VDD2.t4 2.23145
R73 VDD2.n0 VDD2.t0 2.23145
R74 VTAIL.n7 VTAIL.t9 55.5305
R75 VTAIL.n10 VTAIL.t1 55.5305
R76 VTAIL.n11 VTAIL.t6 55.5303
R77 VTAIL.n2 VTAIL.t0 55.5303
R78 VTAIL.n9 VTAIL.n8 53.2996
R79 VTAIL.n6 VTAIL.n5 53.2996
R80 VTAIL.n1 VTAIL.n0 53.2995
R81 VTAIL.n4 VTAIL.n3 53.2995
R82 VTAIL.n6 VTAIL.n4 31.9272
R83 VTAIL.n11 VTAIL.n10 28.4272
R84 VTAIL.n7 VTAIL.n6 3.5005
R85 VTAIL.n10 VTAIL.n9 3.5005
R86 VTAIL.n4 VTAIL.n2 3.5005
R87 VTAIL VTAIL.n11 2.56731
R88 VTAIL.n0 VTAIL.t10 2.23145
R89 VTAIL.n0 VTAIL.t8 2.23145
R90 VTAIL.n3 VTAIL.t5 2.23145
R91 VTAIL.n3 VTAIL.t4 2.23145
R92 VTAIL.n8 VTAIL.t2 2.23145
R93 VTAIL.n8 VTAIL.t3 2.23145
R94 VTAIL.n5 VTAIL.t7 2.23145
R95 VTAIL.n5 VTAIL.t11 2.23145
R96 VTAIL.n9 VTAIL.n7 2.22033
R97 VTAIL.n2 VTAIL.n1 2.22033
R98 VTAIL VTAIL.n1 0.93369
R99 B.n648 B.n647 585
R100 B.n649 B.n88 585
R101 B.n651 B.n650 585
R102 B.n652 B.n87 585
R103 B.n654 B.n653 585
R104 B.n655 B.n86 585
R105 B.n657 B.n656 585
R106 B.n658 B.n85 585
R107 B.n660 B.n659 585
R108 B.n661 B.n84 585
R109 B.n663 B.n662 585
R110 B.n664 B.n83 585
R111 B.n666 B.n665 585
R112 B.n667 B.n82 585
R113 B.n669 B.n668 585
R114 B.n670 B.n81 585
R115 B.n672 B.n671 585
R116 B.n673 B.n80 585
R117 B.n675 B.n674 585
R118 B.n676 B.n79 585
R119 B.n678 B.n677 585
R120 B.n679 B.n78 585
R121 B.n681 B.n680 585
R122 B.n682 B.n77 585
R123 B.n684 B.n683 585
R124 B.n685 B.n76 585
R125 B.n687 B.n686 585
R126 B.n688 B.n75 585
R127 B.n690 B.n689 585
R128 B.n691 B.n74 585
R129 B.n693 B.n692 585
R130 B.n694 B.n73 585
R131 B.n696 B.n695 585
R132 B.n697 B.n72 585
R133 B.n699 B.n698 585
R134 B.n700 B.n71 585
R135 B.n702 B.n701 585
R136 B.n703 B.n70 585
R137 B.n705 B.n704 585
R138 B.n706 B.n69 585
R139 B.n708 B.n707 585
R140 B.n709 B.n68 585
R141 B.n711 B.n710 585
R142 B.n712 B.n67 585
R143 B.n714 B.n713 585
R144 B.n715 B.n66 585
R145 B.n717 B.n716 585
R146 B.n718 B.n65 585
R147 B.n720 B.n719 585
R148 B.n722 B.n62 585
R149 B.n724 B.n723 585
R150 B.n725 B.n61 585
R151 B.n727 B.n726 585
R152 B.n728 B.n60 585
R153 B.n730 B.n729 585
R154 B.n731 B.n59 585
R155 B.n733 B.n732 585
R156 B.n734 B.n55 585
R157 B.n736 B.n735 585
R158 B.n737 B.n54 585
R159 B.n739 B.n738 585
R160 B.n740 B.n53 585
R161 B.n742 B.n741 585
R162 B.n743 B.n52 585
R163 B.n745 B.n744 585
R164 B.n746 B.n51 585
R165 B.n748 B.n747 585
R166 B.n749 B.n50 585
R167 B.n751 B.n750 585
R168 B.n752 B.n49 585
R169 B.n754 B.n753 585
R170 B.n755 B.n48 585
R171 B.n757 B.n756 585
R172 B.n758 B.n47 585
R173 B.n760 B.n759 585
R174 B.n761 B.n46 585
R175 B.n763 B.n762 585
R176 B.n764 B.n45 585
R177 B.n766 B.n765 585
R178 B.n767 B.n44 585
R179 B.n769 B.n768 585
R180 B.n770 B.n43 585
R181 B.n772 B.n771 585
R182 B.n773 B.n42 585
R183 B.n775 B.n774 585
R184 B.n776 B.n41 585
R185 B.n778 B.n777 585
R186 B.n779 B.n40 585
R187 B.n781 B.n780 585
R188 B.n782 B.n39 585
R189 B.n784 B.n783 585
R190 B.n785 B.n38 585
R191 B.n787 B.n786 585
R192 B.n788 B.n37 585
R193 B.n790 B.n789 585
R194 B.n791 B.n36 585
R195 B.n793 B.n792 585
R196 B.n794 B.n35 585
R197 B.n796 B.n795 585
R198 B.n797 B.n34 585
R199 B.n799 B.n798 585
R200 B.n800 B.n33 585
R201 B.n802 B.n801 585
R202 B.n803 B.n32 585
R203 B.n805 B.n804 585
R204 B.n806 B.n31 585
R205 B.n808 B.n807 585
R206 B.n809 B.n30 585
R207 B.n646 B.n89 585
R208 B.n645 B.n644 585
R209 B.n643 B.n90 585
R210 B.n642 B.n641 585
R211 B.n640 B.n91 585
R212 B.n639 B.n638 585
R213 B.n637 B.n92 585
R214 B.n636 B.n635 585
R215 B.n634 B.n93 585
R216 B.n633 B.n632 585
R217 B.n631 B.n94 585
R218 B.n630 B.n629 585
R219 B.n628 B.n95 585
R220 B.n627 B.n626 585
R221 B.n625 B.n96 585
R222 B.n624 B.n623 585
R223 B.n622 B.n97 585
R224 B.n621 B.n620 585
R225 B.n619 B.n98 585
R226 B.n618 B.n617 585
R227 B.n616 B.n99 585
R228 B.n615 B.n614 585
R229 B.n613 B.n100 585
R230 B.n612 B.n611 585
R231 B.n610 B.n101 585
R232 B.n609 B.n608 585
R233 B.n607 B.n102 585
R234 B.n606 B.n605 585
R235 B.n604 B.n103 585
R236 B.n603 B.n602 585
R237 B.n601 B.n104 585
R238 B.n600 B.n599 585
R239 B.n598 B.n105 585
R240 B.n597 B.n596 585
R241 B.n595 B.n106 585
R242 B.n594 B.n593 585
R243 B.n592 B.n107 585
R244 B.n591 B.n590 585
R245 B.n589 B.n108 585
R246 B.n588 B.n587 585
R247 B.n586 B.n109 585
R248 B.n585 B.n584 585
R249 B.n583 B.n110 585
R250 B.n582 B.n581 585
R251 B.n580 B.n111 585
R252 B.n579 B.n578 585
R253 B.n577 B.n112 585
R254 B.n576 B.n575 585
R255 B.n574 B.n113 585
R256 B.n573 B.n572 585
R257 B.n571 B.n114 585
R258 B.n570 B.n569 585
R259 B.n568 B.n115 585
R260 B.n567 B.n566 585
R261 B.n565 B.n116 585
R262 B.n564 B.n563 585
R263 B.n562 B.n117 585
R264 B.n561 B.n560 585
R265 B.n559 B.n118 585
R266 B.n558 B.n557 585
R267 B.n556 B.n119 585
R268 B.n555 B.n554 585
R269 B.n553 B.n120 585
R270 B.n552 B.n551 585
R271 B.n550 B.n121 585
R272 B.n549 B.n548 585
R273 B.n547 B.n122 585
R274 B.n546 B.n545 585
R275 B.n544 B.n123 585
R276 B.n543 B.n542 585
R277 B.n541 B.n124 585
R278 B.n540 B.n539 585
R279 B.n538 B.n125 585
R280 B.n537 B.n536 585
R281 B.n535 B.n126 585
R282 B.n534 B.n533 585
R283 B.n532 B.n127 585
R284 B.n531 B.n530 585
R285 B.n529 B.n128 585
R286 B.n528 B.n527 585
R287 B.n526 B.n129 585
R288 B.n525 B.n524 585
R289 B.n523 B.n130 585
R290 B.n522 B.n521 585
R291 B.n520 B.n131 585
R292 B.n519 B.n518 585
R293 B.n517 B.n132 585
R294 B.n516 B.n515 585
R295 B.n514 B.n133 585
R296 B.n513 B.n512 585
R297 B.n511 B.n134 585
R298 B.n510 B.n509 585
R299 B.n508 B.n135 585
R300 B.n507 B.n506 585
R301 B.n505 B.n136 585
R302 B.n504 B.n503 585
R303 B.n502 B.n137 585
R304 B.n501 B.n500 585
R305 B.n499 B.n138 585
R306 B.n498 B.n497 585
R307 B.n496 B.n139 585
R308 B.n495 B.n494 585
R309 B.n493 B.n140 585
R310 B.n492 B.n491 585
R311 B.n490 B.n141 585
R312 B.n489 B.n488 585
R313 B.n487 B.n142 585
R314 B.n486 B.n485 585
R315 B.n484 B.n143 585
R316 B.n483 B.n482 585
R317 B.n481 B.n144 585
R318 B.n480 B.n479 585
R319 B.n478 B.n145 585
R320 B.n315 B.n314 585
R321 B.n316 B.n203 585
R322 B.n318 B.n317 585
R323 B.n319 B.n202 585
R324 B.n321 B.n320 585
R325 B.n322 B.n201 585
R326 B.n324 B.n323 585
R327 B.n325 B.n200 585
R328 B.n327 B.n326 585
R329 B.n328 B.n199 585
R330 B.n330 B.n329 585
R331 B.n331 B.n198 585
R332 B.n333 B.n332 585
R333 B.n334 B.n197 585
R334 B.n336 B.n335 585
R335 B.n337 B.n196 585
R336 B.n339 B.n338 585
R337 B.n340 B.n195 585
R338 B.n342 B.n341 585
R339 B.n343 B.n194 585
R340 B.n345 B.n344 585
R341 B.n346 B.n193 585
R342 B.n348 B.n347 585
R343 B.n349 B.n192 585
R344 B.n351 B.n350 585
R345 B.n352 B.n191 585
R346 B.n354 B.n353 585
R347 B.n355 B.n190 585
R348 B.n357 B.n356 585
R349 B.n358 B.n189 585
R350 B.n360 B.n359 585
R351 B.n361 B.n188 585
R352 B.n363 B.n362 585
R353 B.n364 B.n187 585
R354 B.n366 B.n365 585
R355 B.n367 B.n186 585
R356 B.n369 B.n368 585
R357 B.n370 B.n185 585
R358 B.n372 B.n371 585
R359 B.n373 B.n184 585
R360 B.n375 B.n374 585
R361 B.n376 B.n183 585
R362 B.n378 B.n377 585
R363 B.n379 B.n182 585
R364 B.n381 B.n380 585
R365 B.n382 B.n181 585
R366 B.n384 B.n383 585
R367 B.n385 B.n180 585
R368 B.n387 B.n386 585
R369 B.n389 B.n388 585
R370 B.n390 B.n176 585
R371 B.n392 B.n391 585
R372 B.n393 B.n175 585
R373 B.n395 B.n394 585
R374 B.n396 B.n174 585
R375 B.n398 B.n397 585
R376 B.n399 B.n173 585
R377 B.n401 B.n400 585
R378 B.n402 B.n170 585
R379 B.n405 B.n404 585
R380 B.n406 B.n169 585
R381 B.n408 B.n407 585
R382 B.n409 B.n168 585
R383 B.n411 B.n410 585
R384 B.n412 B.n167 585
R385 B.n414 B.n413 585
R386 B.n415 B.n166 585
R387 B.n417 B.n416 585
R388 B.n418 B.n165 585
R389 B.n420 B.n419 585
R390 B.n421 B.n164 585
R391 B.n423 B.n422 585
R392 B.n424 B.n163 585
R393 B.n426 B.n425 585
R394 B.n427 B.n162 585
R395 B.n429 B.n428 585
R396 B.n430 B.n161 585
R397 B.n432 B.n431 585
R398 B.n433 B.n160 585
R399 B.n435 B.n434 585
R400 B.n436 B.n159 585
R401 B.n438 B.n437 585
R402 B.n439 B.n158 585
R403 B.n441 B.n440 585
R404 B.n442 B.n157 585
R405 B.n444 B.n443 585
R406 B.n445 B.n156 585
R407 B.n447 B.n446 585
R408 B.n448 B.n155 585
R409 B.n450 B.n449 585
R410 B.n451 B.n154 585
R411 B.n453 B.n452 585
R412 B.n454 B.n153 585
R413 B.n456 B.n455 585
R414 B.n457 B.n152 585
R415 B.n459 B.n458 585
R416 B.n460 B.n151 585
R417 B.n462 B.n461 585
R418 B.n463 B.n150 585
R419 B.n465 B.n464 585
R420 B.n466 B.n149 585
R421 B.n468 B.n467 585
R422 B.n469 B.n148 585
R423 B.n471 B.n470 585
R424 B.n472 B.n147 585
R425 B.n474 B.n473 585
R426 B.n475 B.n146 585
R427 B.n477 B.n476 585
R428 B.n313 B.n204 585
R429 B.n312 B.n311 585
R430 B.n310 B.n205 585
R431 B.n309 B.n308 585
R432 B.n307 B.n206 585
R433 B.n306 B.n305 585
R434 B.n304 B.n207 585
R435 B.n303 B.n302 585
R436 B.n301 B.n208 585
R437 B.n300 B.n299 585
R438 B.n298 B.n209 585
R439 B.n297 B.n296 585
R440 B.n295 B.n210 585
R441 B.n294 B.n293 585
R442 B.n292 B.n211 585
R443 B.n291 B.n290 585
R444 B.n289 B.n212 585
R445 B.n288 B.n287 585
R446 B.n286 B.n213 585
R447 B.n285 B.n284 585
R448 B.n283 B.n214 585
R449 B.n282 B.n281 585
R450 B.n280 B.n215 585
R451 B.n279 B.n278 585
R452 B.n277 B.n216 585
R453 B.n276 B.n275 585
R454 B.n274 B.n217 585
R455 B.n273 B.n272 585
R456 B.n271 B.n218 585
R457 B.n270 B.n269 585
R458 B.n268 B.n219 585
R459 B.n267 B.n266 585
R460 B.n265 B.n220 585
R461 B.n264 B.n263 585
R462 B.n262 B.n221 585
R463 B.n261 B.n260 585
R464 B.n259 B.n222 585
R465 B.n258 B.n257 585
R466 B.n256 B.n223 585
R467 B.n255 B.n254 585
R468 B.n253 B.n224 585
R469 B.n252 B.n251 585
R470 B.n250 B.n225 585
R471 B.n249 B.n248 585
R472 B.n247 B.n226 585
R473 B.n246 B.n245 585
R474 B.n244 B.n227 585
R475 B.n243 B.n242 585
R476 B.n241 B.n228 585
R477 B.n240 B.n239 585
R478 B.n238 B.n229 585
R479 B.n237 B.n236 585
R480 B.n235 B.n230 585
R481 B.n234 B.n233 585
R482 B.n232 B.n231 585
R483 B.n2 B.n0 585
R484 B.n893 B.n1 585
R485 B.n892 B.n891 585
R486 B.n890 B.n3 585
R487 B.n889 B.n888 585
R488 B.n887 B.n4 585
R489 B.n886 B.n885 585
R490 B.n884 B.n5 585
R491 B.n883 B.n882 585
R492 B.n881 B.n6 585
R493 B.n880 B.n879 585
R494 B.n878 B.n7 585
R495 B.n877 B.n876 585
R496 B.n875 B.n8 585
R497 B.n874 B.n873 585
R498 B.n872 B.n9 585
R499 B.n871 B.n870 585
R500 B.n869 B.n10 585
R501 B.n868 B.n867 585
R502 B.n866 B.n11 585
R503 B.n865 B.n864 585
R504 B.n863 B.n12 585
R505 B.n862 B.n861 585
R506 B.n860 B.n13 585
R507 B.n859 B.n858 585
R508 B.n857 B.n14 585
R509 B.n856 B.n855 585
R510 B.n854 B.n15 585
R511 B.n853 B.n852 585
R512 B.n851 B.n16 585
R513 B.n850 B.n849 585
R514 B.n848 B.n17 585
R515 B.n847 B.n846 585
R516 B.n845 B.n18 585
R517 B.n844 B.n843 585
R518 B.n842 B.n19 585
R519 B.n841 B.n840 585
R520 B.n839 B.n20 585
R521 B.n838 B.n837 585
R522 B.n836 B.n21 585
R523 B.n835 B.n834 585
R524 B.n833 B.n22 585
R525 B.n832 B.n831 585
R526 B.n830 B.n23 585
R527 B.n829 B.n828 585
R528 B.n827 B.n24 585
R529 B.n826 B.n825 585
R530 B.n824 B.n25 585
R531 B.n823 B.n822 585
R532 B.n821 B.n26 585
R533 B.n820 B.n819 585
R534 B.n818 B.n27 585
R535 B.n817 B.n816 585
R536 B.n815 B.n28 585
R537 B.n814 B.n813 585
R538 B.n812 B.n29 585
R539 B.n811 B.n810 585
R540 B.n895 B.n894 585
R541 B.n315 B.n204 473.281
R542 B.n810 B.n809 473.281
R543 B.n478 B.n477 473.281
R544 B.n647 B.n646 473.281
R545 B.n171 B.t9 303.428
R546 B.n177 B.t0 303.428
R547 B.n56 B.t3 303.428
R548 B.n63 B.t6 303.428
R549 B.n171 B.t11 190.988
R550 B.n63 B.t7 190.988
R551 B.n177 B.t2 190.97
R552 B.n56 B.t4 190.97
R553 B.n311 B.n204 163.367
R554 B.n311 B.n310 163.367
R555 B.n310 B.n309 163.367
R556 B.n309 B.n206 163.367
R557 B.n305 B.n206 163.367
R558 B.n305 B.n304 163.367
R559 B.n304 B.n303 163.367
R560 B.n303 B.n208 163.367
R561 B.n299 B.n208 163.367
R562 B.n299 B.n298 163.367
R563 B.n298 B.n297 163.367
R564 B.n297 B.n210 163.367
R565 B.n293 B.n210 163.367
R566 B.n293 B.n292 163.367
R567 B.n292 B.n291 163.367
R568 B.n291 B.n212 163.367
R569 B.n287 B.n212 163.367
R570 B.n287 B.n286 163.367
R571 B.n286 B.n285 163.367
R572 B.n285 B.n214 163.367
R573 B.n281 B.n214 163.367
R574 B.n281 B.n280 163.367
R575 B.n280 B.n279 163.367
R576 B.n279 B.n216 163.367
R577 B.n275 B.n216 163.367
R578 B.n275 B.n274 163.367
R579 B.n274 B.n273 163.367
R580 B.n273 B.n218 163.367
R581 B.n269 B.n218 163.367
R582 B.n269 B.n268 163.367
R583 B.n268 B.n267 163.367
R584 B.n267 B.n220 163.367
R585 B.n263 B.n220 163.367
R586 B.n263 B.n262 163.367
R587 B.n262 B.n261 163.367
R588 B.n261 B.n222 163.367
R589 B.n257 B.n222 163.367
R590 B.n257 B.n256 163.367
R591 B.n256 B.n255 163.367
R592 B.n255 B.n224 163.367
R593 B.n251 B.n224 163.367
R594 B.n251 B.n250 163.367
R595 B.n250 B.n249 163.367
R596 B.n249 B.n226 163.367
R597 B.n245 B.n226 163.367
R598 B.n245 B.n244 163.367
R599 B.n244 B.n243 163.367
R600 B.n243 B.n228 163.367
R601 B.n239 B.n228 163.367
R602 B.n239 B.n238 163.367
R603 B.n238 B.n237 163.367
R604 B.n237 B.n230 163.367
R605 B.n233 B.n230 163.367
R606 B.n233 B.n232 163.367
R607 B.n232 B.n2 163.367
R608 B.n894 B.n2 163.367
R609 B.n894 B.n893 163.367
R610 B.n893 B.n892 163.367
R611 B.n892 B.n3 163.367
R612 B.n888 B.n3 163.367
R613 B.n888 B.n887 163.367
R614 B.n887 B.n886 163.367
R615 B.n886 B.n5 163.367
R616 B.n882 B.n5 163.367
R617 B.n882 B.n881 163.367
R618 B.n881 B.n880 163.367
R619 B.n880 B.n7 163.367
R620 B.n876 B.n7 163.367
R621 B.n876 B.n875 163.367
R622 B.n875 B.n874 163.367
R623 B.n874 B.n9 163.367
R624 B.n870 B.n9 163.367
R625 B.n870 B.n869 163.367
R626 B.n869 B.n868 163.367
R627 B.n868 B.n11 163.367
R628 B.n864 B.n11 163.367
R629 B.n864 B.n863 163.367
R630 B.n863 B.n862 163.367
R631 B.n862 B.n13 163.367
R632 B.n858 B.n13 163.367
R633 B.n858 B.n857 163.367
R634 B.n857 B.n856 163.367
R635 B.n856 B.n15 163.367
R636 B.n852 B.n15 163.367
R637 B.n852 B.n851 163.367
R638 B.n851 B.n850 163.367
R639 B.n850 B.n17 163.367
R640 B.n846 B.n17 163.367
R641 B.n846 B.n845 163.367
R642 B.n845 B.n844 163.367
R643 B.n844 B.n19 163.367
R644 B.n840 B.n19 163.367
R645 B.n840 B.n839 163.367
R646 B.n839 B.n838 163.367
R647 B.n838 B.n21 163.367
R648 B.n834 B.n21 163.367
R649 B.n834 B.n833 163.367
R650 B.n833 B.n832 163.367
R651 B.n832 B.n23 163.367
R652 B.n828 B.n23 163.367
R653 B.n828 B.n827 163.367
R654 B.n827 B.n826 163.367
R655 B.n826 B.n25 163.367
R656 B.n822 B.n25 163.367
R657 B.n822 B.n821 163.367
R658 B.n821 B.n820 163.367
R659 B.n820 B.n27 163.367
R660 B.n816 B.n27 163.367
R661 B.n816 B.n815 163.367
R662 B.n815 B.n814 163.367
R663 B.n814 B.n29 163.367
R664 B.n810 B.n29 163.367
R665 B.n316 B.n315 163.367
R666 B.n317 B.n316 163.367
R667 B.n317 B.n202 163.367
R668 B.n321 B.n202 163.367
R669 B.n322 B.n321 163.367
R670 B.n323 B.n322 163.367
R671 B.n323 B.n200 163.367
R672 B.n327 B.n200 163.367
R673 B.n328 B.n327 163.367
R674 B.n329 B.n328 163.367
R675 B.n329 B.n198 163.367
R676 B.n333 B.n198 163.367
R677 B.n334 B.n333 163.367
R678 B.n335 B.n334 163.367
R679 B.n335 B.n196 163.367
R680 B.n339 B.n196 163.367
R681 B.n340 B.n339 163.367
R682 B.n341 B.n340 163.367
R683 B.n341 B.n194 163.367
R684 B.n345 B.n194 163.367
R685 B.n346 B.n345 163.367
R686 B.n347 B.n346 163.367
R687 B.n347 B.n192 163.367
R688 B.n351 B.n192 163.367
R689 B.n352 B.n351 163.367
R690 B.n353 B.n352 163.367
R691 B.n353 B.n190 163.367
R692 B.n357 B.n190 163.367
R693 B.n358 B.n357 163.367
R694 B.n359 B.n358 163.367
R695 B.n359 B.n188 163.367
R696 B.n363 B.n188 163.367
R697 B.n364 B.n363 163.367
R698 B.n365 B.n364 163.367
R699 B.n365 B.n186 163.367
R700 B.n369 B.n186 163.367
R701 B.n370 B.n369 163.367
R702 B.n371 B.n370 163.367
R703 B.n371 B.n184 163.367
R704 B.n375 B.n184 163.367
R705 B.n376 B.n375 163.367
R706 B.n377 B.n376 163.367
R707 B.n377 B.n182 163.367
R708 B.n381 B.n182 163.367
R709 B.n382 B.n381 163.367
R710 B.n383 B.n382 163.367
R711 B.n383 B.n180 163.367
R712 B.n387 B.n180 163.367
R713 B.n388 B.n387 163.367
R714 B.n388 B.n176 163.367
R715 B.n392 B.n176 163.367
R716 B.n393 B.n392 163.367
R717 B.n394 B.n393 163.367
R718 B.n394 B.n174 163.367
R719 B.n398 B.n174 163.367
R720 B.n399 B.n398 163.367
R721 B.n400 B.n399 163.367
R722 B.n400 B.n170 163.367
R723 B.n405 B.n170 163.367
R724 B.n406 B.n405 163.367
R725 B.n407 B.n406 163.367
R726 B.n407 B.n168 163.367
R727 B.n411 B.n168 163.367
R728 B.n412 B.n411 163.367
R729 B.n413 B.n412 163.367
R730 B.n413 B.n166 163.367
R731 B.n417 B.n166 163.367
R732 B.n418 B.n417 163.367
R733 B.n419 B.n418 163.367
R734 B.n419 B.n164 163.367
R735 B.n423 B.n164 163.367
R736 B.n424 B.n423 163.367
R737 B.n425 B.n424 163.367
R738 B.n425 B.n162 163.367
R739 B.n429 B.n162 163.367
R740 B.n430 B.n429 163.367
R741 B.n431 B.n430 163.367
R742 B.n431 B.n160 163.367
R743 B.n435 B.n160 163.367
R744 B.n436 B.n435 163.367
R745 B.n437 B.n436 163.367
R746 B.n437 B.n158 163.367
R747 B.n441 B.n158 163.367
R748 B.n442 B.n441 163.367
R749 B.n443 B.n442 163.367
R750 B.n443 B.n156 163.367
R751 B.n447 B.n156 163.367
R752 B.n448 B.n447 163.367
R753 B.n449 B.n448 163.367
R754 B.n449 B.n154 163.367
R755 B.n453 B.n154 163.367
R756 B.n454 B.n453 163.367
R757 B.n455 B.n454 163.367
R758 B.n455 B.n152 163.367
R759 B.n459 B.n152 163.367
R760 B.n460 B.n459 163.367
R761 B.n461 B.n460 163.367
R762 B.n461 B.n150 163.367
R763 B.n465 B.n150 163.367
R764 B.n466 B.n465 163.367
R765 B.n467 B.n466 163.367
R766 B.n467 B.n148 163.367
R767 B.n471 B.n148 163.367
R768 B.n472 B.n471 163.367
R769 B.n473 B.n472 163.367
R770 B.n473 B.n146 163.367
R771 B.n477 B.n146 163.367
R772 B.n479 B.n478 163.367
R773 B.n479 B.n144 163.367
R774 B.n483 B.n144 163.367
R775 B.n484 B.n483 163.367
R776 B.n485 B.n484 163.367
R777 B.n485 B.n142 163.367
R778 B.n489 B.n142 163.367
R779 B.n490 B.n489 163.367
R780 B.n491 B.n490 163.367
R781 B.n491 B.n140 163.367
R782 B.n495 B.n140 163.367
R783 B.n496 B.n495 163.367
R784 B.n497 B.n496 163.367
R785 B.n497 B.n138 163.367
R786 B.n501 B.n138 163.367
R787 B.n502 B.n501 163.367
R788 B.n503 B.n502 163.367
R789 B.n503 B.n136 163.367
R790 B.n507 B.n136 163.367
R791 B.n508 B.n507 163.367
R792 B.n509 B.n508 163.367
R793 B.n509 B.n134 163.367
R794 B.n513 B.n134 163.367
R795 B.n514 B.n513 163.367
R796 B.n515 B.n514 163.367
R797 B.n515 B.n132 163.367
R798 B.n519 B.n132 163.367
R799 B.n520 B.n519 163.367
R800 B.n521 B.n520 163.367
R801 B.n521 B.n130 163.367
R802 B.n525 B.n130 163.367
R803 B.n526 B.n525 163.367
R804 B.n527 B.n526 163.367
R805 B.n527 B.n128 163.367
R806 B.n531 B.n128 163.367
R807 B.n532 B.n531 163.367
R808 B.n533 B.n532 163.367
R809 B.n533 B.n126 163.367
R810 B.n537 B.n126 163.367
R811 B.n538 B.n537 163.367
R812 B.n539 B.n538 163.367
R813 B.n539 B.n124 163.367
R814 B.n543 B.n124 163.367
R815 B.n544 B.n543 163.367
R816 B.n545 B.n544 163.367
R817 B.n545 B.n122 163.367
R818 B.n549 B.n122 163.367
R819 B.n550 B.n549 163.367
R820 B.n551 B.n550 163.367
R821 B.n551 B.n120 163.367
R822 B.n555 B.n120 163.367
R823 B.n556 B.n555 163.367
R824 B.n557 B.n556 163.367
R825 B.n557 B.n118 163.367
R826 B.n561 B.n118 163.367
R827 B.n562 B.n561 163.367
R828 B.n563 B.n562 163.367
R829 B.n563 B.n116 163.367
R830 B.n567 B.n116 163.367
R831 B.n568 B.n567 163.367
R832 B.n569 B.n568 163.367
R833 B.n569 B.n114 163.367
R834 B.n573 B.n114 163.367
R835 B.n574 B.n573 163.367
R836 B.n575 B.n574 163.367
R837 B.n575 B.n112 163.367
R838 B.n579 B.n112 163.367
R839 B.n580 B.n579 163.367
R840 B.n581 B.n580 163.367
R841 B.n581 B.n110 163.367
R842 B.n585 B.n110 163.367
R843 B.n586 B.n585 163.367
R844 B.n587 B.n586 163.367
R845 B.n587 B.n108 163.367
R846 B.n591 B.n108 163.367
R847 B.n592 B.n591 163.367
R848 B.n593 B.n592 163.367
R849 B.n593 B.n106 163.367
R850 B.n597 B.n106 163.367
R851 B.n598 B.n597 163.367
R852 B.n599 B.n598 163.367
R853 B.n599 B.n104 163.367
R854 B.n603 B.n104 163.367
R855 B.n604 B.n603 163.367
R856 B.n605 B.n604 163.367
R857 B.n605 B.n102 163.367
R858 B.n609 B.n102 163.367
R859 B.n610 B.n609 163.367
R860 B.n611 B.n610 163.367
R861 B.n611 B.n100 163.367
R862 B.n615 B.n100 163.367
R863 B.n616 B.n615 163.367
R864 B.n617 B.n616 163.367
R865 B.n617 B.n98 163.367
R866 B.n621 B.n98 163.367
R867 B.n622 B.n621 163.367
R868 B.n623 B.n622 163.367
R869 B.n623 B.n96 163.367
R870 B.n627 B.n96 163.367
R871 B.n628 B.n627 163.367
R872 B.n629 B.n628 163.367
R873 B.n629 B.n94 163.367
R874 B.n633 B.n94 163.367
R875 B.n634 B.n633 163.367
R876 B.n635 B.n634 163.367
R877 B.n635 B.n92 163.367
R878 B.n639 B.n92 163.367
R879 B.n640 B.n639 163.367
R880 B.n641 B.n640 163.367
R881 B.n641 B.n90 163.367
R882 B.n645 B.n90 163.367
R883 B.n646 B.n645 163.367
R884 B.n809 B.n808 163.367
R885 B.n808 B.n31 163.367
R886 B.n804 B.n31 163.367
R887 B.n804 B.n803 163.367
R888 B.n803 B.n802 163.367
R889 B.n802 B.n33 163.367
R890 B.n798 B.n33 163.367
R891 B.n798 B.n797 163.367
R892 B.n797 B.n796 163.367
R893 B.n796 B.n35 163.367
R894 B.n792 B.n35 163.367
R895 B.n792 B.n791 163.367
R896 B.n791 B.n790 163.367
R897 B.n790 B.n37 163.367
R898 B.n786 B.n37 163.367
R899 B.n786 B.n785 163.367
R900 B.n785 B.n784 163.367
R901 B.n784 B.n39 163.367
R902 B.n780 B.n39 163.367
R903 B.n780 B.n779 163.367
R904 B.n779 B.n778 163.367
R905 B.n778 B.n41 163.367
R906 B.n774 B.n41 163.367
R907 B.n774 B.n773 163.367
R908 B.n773 B.n772 163.367
R909 B.n772 B.n43 163.367
R910 B.n768 B.n43 163.367
R911 B.n768 B.n767 163.367
R912 B.n767 B.n766 163.367
R913 B.n766 B.n45 163.367
R914 B.n762 B.n45 163.367
R915 B.n762 B.n761 163.367
R916 B.n761 B.n760 163.367
R917 B.n760 B.n47 163.367
R918 B.n756 B.n47 163.367
R919 B.n756 B.n755 163.367
R920 B.n755 B.n754 163.367
R921 B.n754 B.n49 163.367
R922 B.n750 B.n49 163.367
R923 B.n750 B.n749 163.367
R924 B.n749 B.n748 163.367
R925 B.n748 B.n51 163.367
R926 B.n744 B.n51 163.367
R927 B.n744 B.n743 163.367
R928 B.n743 B.n742 163.367
R929 B.n742 B.n53 163.367
R930 B.n738 B.n53 163.367
R931 B.n738 B.n737 163.367
R932 B.n737 B.n736 163.367
R933 B.n736 B.n55 163.367
R934 B.n732 B.n55 163.367
R935 B.n732 B.n731 163.367
R936 B.n731 B.n730 163.367
R937 B.n730 B.n60 163.367
R938 B.n726 B.n60 163.367
R939 B.n726 B.n725 163.367
R940 B.n725 B.n724 163.367
R941 B.n724 B.n62 163.367
R942 B.n719 B.n62 163.367
R943 B.n719 B.n718 163.367
R944 B.n718 B.n717 163.367
R945 B.n717 B.n66 163.367
R946 B.n713 B.n66 163.367
R947 B.n713 B.n712 163.367
R948 B.n712 B.n711 163.367
R949 B.n711 B.n68 163.367
R950 B.n707 B.n68 163.367
R951 B.n707 B.n706 163.367
R952 B.n706 B.n705 163.367
R953 B.n705 B.n70 163.367
R954 B.n701 B.n70 163.367
R955 B.n701 B.n700 163.367
R956 B.n700 B.n699 163.367
R957 B.n699 B.n72 163.367
R958 B.n695 B.n72 163.367
R959 B.n695 B.n694 163.367
R960 B.n694 B.n693 163.367
R961 B.n693 B.n74 163.367
R962 B.n689 B.n74 163.367
R963 B.n689 B.n688 163.367
R964 B.n688 B.n687 163.367
R965 B.n687 B.n76 163.367
R966 B.n683 B.n76 163.367
R967 B.n683 B.n682 163.367
R968 B.n682 B.n681 163.367
R969 B.n681 B.n78 163.367
R970 B.n677 B.n78 163.367
R971 B.n677 B.n676 163.367
R972 B.n676 B.n675 163.367
R973 B.n675 B.n80 163.367
R974 B.n671 B.n80 163.367
R975 B.n671 B.n670 163.367
R976 B.n670 B.n669 163.367
R977 B.n669 B.n82 163.367
R978 B.n665 B.n82 163.367
R979 B.n665 B.n664 163.367
R980 B.n664 B.n663 163.367
R981 B.n663 B.n84 163.367
R982 B.n659 B.n84 163.367
R983 B.n659 B.n658 163.367
R984 B.n658 B.n657 163.367
R985 B.n657 B.n86 163.367
R986 B.n653 B.n86 163.367
R987 B.n653 B.n652 163.367
R988 B.n652 B.n651 163.367
R989 B.n651 B.n88 163.367
R990 B.n647 B.n88 163.367
R991 B.n172 B.t10 112.249
R992 B.n64 B.t8 112.249
R993 B.n178 B.t1 112.231
R994 B.n57 B.t5 112.231
R995 B.n172 B.n171 78.7399
R996 B.n178 B.n177 78.7399
R997 B.n57 B.n56 78.7399
R998 B.n64 B.n63 78.7399
R999 B.n403 B.n172 59.5399
R1000 B.n179 B.n178 59.5399
R1001 B.n58 B.n57 59.5399
R1002 B.n721 B.n64 59.5399
R1003 B.n811 B.n30 30.7517
R1004 B.n648 B.n89 30.7517
R1005 B.n476 B.n145 30.7517
R1006 B.n314 B.n313 30.7517
R1007 B B.n895 18.0485
R1008 B.n807 B.n30 10.6151
R1009 B.n807 B.n806 10.6151
R1010 B.n806 B.n805 10.6151
R1011 B.n805 B.n32 10.6151
R1012 B.n801 B.n32 10.6151
R1013 B.n801 B.n800 10.6151
R1014 B.n800 B.n799 10.6151
R1015 B.n799 B.n34 10.6151
R1016 B.n795 B.n34 10.6151
R1017 B.n795 B.n794 10.6151
R1018 B.n794 B.n793 10.6151
R1019 B.n793 B.n36 10.6151
R1020 B.n789 B.n36 10.6151
R1021 B.n789 B.n788 10.6151
R1022 B.n788 B.n787 10.6151
R1023 B.n787 B.n38 10.6151
R1024 B.n783 B.n38 10.6151
R1025 B.n783 B.n782 10.6151
R1026 B.n782 B.n781 10.6151
R1027 B.n781 B.n40 10.6151
R1028 B.n777 B.n40 10.6151
R1029 B.n777 B.n776 10.6151
R1030 B.n776 B.n775 10.6151
R1031 B.n775 B.n42 10.6151
R1032 B.n771 B.n42 10.6151
R1033 B.n771 B.n770 10.6151
R1034 B.n770 B.n769 10.6151
R1035 B.n769 B.n44 10.6151
R1036 B.n765 B.n44 10.6151
R1037 B.n765 B.n764 10.6151
R1038 B.n764 B.n763 10.6151
R1039 B.n763 B.n46 10.6151
R1040 B.n759 B.n46 10.6151
R1041 B.n759 B.n758 10.6151
R1042 B.n758 B.n757 10.6151
R1043 B.n757 B.n48 10.6151
R1044 B.n753 B.n48 10.6151
R1045 B.n753 B.n752 10.6151
R1046 B.n752 B.n751 10.6151
R1047 B.n751 B.n50 10.6151
R1048 B.n747 B.n50 10.6151
R1049 B.n747 B.n746 10.6151
R1050 B.n746 B.n745 10.6151
R1051 B.n745 B.n52 10.6151
R1052 B.n741 B.n52 10.6151
R1053 B.n741 B.n740 10.6151
R1054 B.n740 B.n739 10.6151
R1055 B.n739 B.n54 10.6151
R1056 B.n735 B.n734 10.6151
R1057 B.n734 B.n733 10.6151
R1058 B.n733 B.n59 10.6151
R1059 B.n729 B.n59 10.6151
R1060 B.n729 B.n728 10.6151
R1061 B.n728 B.n727 10.6151
R1062 B.n727 B.n61 10.6151
R1063 B.n723 B.n61 10.6151
R1064 B.n723 B.n722 10.6151
R1065 B.n720 B.n65 10.6151
R1066 B.n716 B.n65 10.6151
R1067 B.n716 B.n715 10.6151
R1068 B.n715 B.n714 10.6151
R1069 B.n714 B.n67 10.6151
R1070 B.n710 B.n67 10.6151
R1071 B.n710 B.n709 10.6151
R1072 B.n709 B.n708 10.6151
R1073 B.n708 B.n69 10.6151
R1074 B.n704 B.n69 10.6151
R1075 B.n704 B.n703 10.6151
R1076 B.n703 B.n702 10.6151
R1077 B.n702 B.n71 10.6151
R1078 B.n698 B.n71 10.6151
R1079 B.n698 B.n697 10.6151
R1080 B.n697 B.n696 10.6151
R1081 B.n696 B.n73 10.6151
R1082 B.n692 B.n73 10.6151
R1083 B.n692 B.n691 10.6151
R1084 B.n691 B.n690 10.6151
R1085 B.n690 B.n75 10.6151
R1086 B.n686 B.n75 10.6151
R1087 B.n686 B.n685 10.6151
R1088 B.n685 B.n684 10.6151
R1089 B.n684 B.n77 10.6151
R1090 B.n680 B.n77 10.6151
R1091 B.n680 B.n679 10.6151
R1092 B.n679 B.n678 10.6151
R1093 B.n678 B.n79 10.6151
R1094 B.n674 B.n79 10.6151
R1095 B.n674 B.n673 10.6151
R1096 B.n673 B.n672 10.6151
R1097 B.n672 B.n81 10.6151
R1098 B.n668 B.n81 10.6151
R1099 B.n668 B.n667 10.6151
R1100 B.n667 B.n666 10.6151
R1101 B.n666 B.n83 10.6151
R1102 B.n662 B.n83 10.6151
R1103 B.n662 B.n661 10.6151
R1104 B.n661 B.n660 10.6151
R1105 B.n660 B.n85 10.6151
R1106 B.n656 B.n85 10.6151
R1107 B.n656 B.n655 10.6151
R1108 B.n655 B.n654 10.6151
R1109 B.n654 B.n87 10.6151
R1110 B.n650 B.n87 10.6151
R1111 B.n650 B.n649 10.6151
R1112 B.n649 B.n648 10.6151
R1113 B.n480 B.n145 10.6151
R1114 B.n481 B.n480 10.6151
R1115 B.n482 B.n481 10.6151
R1116 B.n482 B.n143 10.6151
R1117 B.n486 B.n143 10.6151
R1118 B.n487 B.n486 10.6151
R1119 B.n488 B.n487 10.6151
R1120 B.n488 B.n141 10.6151
R1121 B.n492 B.n141 10.6151
R1122 B.n493 B.n492 10.6151
R1123 B.n494 B.n493 10.6151
R1124 B.n494 B.n139 10.6151
R1125 B.n498 B.n139 10.6151
R1126 B.n499 B.n498 10.6151
R1127 B.n500 B.n499 10.6151
R1128 B.n500 B.n137 10.6151
R1129 B.n504 B.n137 10.6151
R1130 B.n505 B.n504 10.6151
R1131 B.n506 B.n505 10.6151
R1132 B.n506 B.n135 10.6151
R1133 B.n510 B.n135 10.6151
R1134 B.n511 B.n510 10.6151
R1135 B.n512 B.n511 10.6151
R1136 B.n512 B.n133 10.6151
R1137 B.n516 B.n133 10.6151
R1138 B.n517 B.n516 10.6151
R1139 B.n518 B.n517 10.6151
R1140 B.n518 B.n131 10.6151
R1141 B.n522 B.n131 10.6151
R1142 B.n523 B.n522 10.6151
R1143 B.n524 B.n523 10.6151
R1144 B.n524 B.n129 10.6151
R1145 B.n528 B.n129 10.6151
R1146 B.n529 B.n528 10.6151
R1147 B.n530 B.n529 10.6151
R1148 B.n530 B.n127 10.6151
R1149 B.n534 B.n127 10.6151
R1150 B.n535 B.n534 10.6151
R1151 B.n536 B.n535 10.6151
R1152 B.n536 B.n125 10.6151
R1153 B.n540 B.n125 10.6151
R1154 B.n541 B.n540 10.6151
R1155 B.n542 B.n541 10.6151
R1156 B.n542 B.n123 10.6151
R1157 B.n546 B.n123 10.6151
R1158 B.n547 B.n546 10.6151
R1159 B.n548 B.n547 10.6151
R1160 B.n548 B.n121 10.6151
R1161 B.n552 B.n121 10.6151
R1162 B.n553 B.n552 10.6151
R1163 B.n554 B.n553 10.6151
R1164 B.n554 B.n119 10.6151
R1165 B.n558 B.n119 10.6151
R1166 B.n559 B.n558 10.6151
R1167 B.n560 B.n559 10.6151
R1168 B.n560 B.n117 10.6151
R1169 B.n564 B.n117 10.6151
R1170 B.n565 B.n564 10.6151
R1171 B.n566 B.n565 10.6151
R1172 B.n566 B.n115 10.6151
R1173 B.n570 B.n115 10.6151
R1174 B.n571 B.n570 10.6151
R1175 B.n572 B.n571 10.6151
R1176 B.n572 B.n113 10.6151
R1177 B.n576 B.n113 10.6151
R1178 B.n577 B.n576 10.6151
R1179 B.n578 B.n577 10.6151
R1180 B.n578 B.n111 10.6151
R1181 B.n582 B.n111 10.6151
R1182 B.n583 B.n582 10.6151
R1183 B.n584 B.n583 10.6151
R1184 B.n584 B.n109 10.6151
R1185 B.n588 B.n109 10.6151
R1186 B.n589 B.n588 10.6151
R1187 B.n590 B.n589 10.6151
R1188 B.n590 B.n107 10.6151
R1189 B.n594 B.n107 10.6151
R1190 B.n595 B.n594 10.6151
R1191 B.n596 B.n595 10.6151
R1192 B.n596 B.n105 10.6151
R1193 B.n600 B.n105 10.6151
R1194 B.n601 B.n600 10.6151
R1195 B.n602 B.n601 10.6151
R1196 B.n602 B.n103 10.6151
R1197 B.n606 B.n103 10.6151
R1198 B.n607 B.n606 10.6151
R1199 B.n608 B.n607 10.6151
R1200 B.n608 B.n101 10.6151
R1201 B.n612 B.n101 10.6151
R1202 B.n613 B.n612 10.6151
R1203 B.n614 B.n613 10.6151
R1204 B.n614 B.n99 10.6151
R1205 B.n618 B.n99 10.6151
R1206 B.n619 B.n618 10.6151
R1207 B.n620 B.n619 10.6151
R1208 B.n620 B.n97 10.6151
R1209 B.n624 B.n97 10.6151
R1210 B.n625 B.n624 10.6151
R1211 B.n626 B.n625 10.6151
R1212 B.n626 B.n95 10.6151
R1213 B.n630 B.n95 10.6151
R1214 B.n631 B.n630 10.6151
R1215 B.n632 B.n631 10.6151
R1216 B.n632 B.n93 10.6151
R1217 B.n636 B.n93 10.6151
R1218 B.n637 B.n636 10.6151
R1219 B.n638 B.n637 10.6151
R1220 B.n638 B.n91 10.6151
R1221 B.n642 B.n91 10.6151
R1222 B.n643 B.n642 10.6151
R1223 B.n644 B.n643 10.6151
R1224 B.n644 B.n89 10.6151
R1225 B.n314 B.n203 10.6151
R1226 B.n318 B.n203 10.6151
R1227 B.n319 B.n318 10.6151
R1228 B.n320 B.n319 10.6151
R1229 B.n320 B.n201 10.6151
R1230 B.n324 B.n201 10.6151
R1231 B.n325 B.n324 10.6151
R1232 B.n326 B.n325 10.6151
R1233 B.n326 B.n199 10.6151
R1234 B.n330 B.n199 10.6151
R1235 B.n331 B.n330 10.6151
R1236 B.n332 B.n331 10.6151
R1237 B.n332 B.n197 10.6151
R1238 B.n336 B.n197 10.6151
R1239 B.n337 B.n336 10.6151
R1240 B.n338 B.n337 10.6151
R1241 B.n338 B.n195 10.6151
R1242 B.n342 B.n195 10.6151
R1243 B.n343 B.n342 10.6151
R1244 B.n344 B.n343 10.6151
R1245 B.n344 B.n193 10.6151
R1246 B.n348 B.n193 10.6151
R1247 B.n349 B.n348 10.6151
R1248 B.n350 B.n349 10.6151
R1249 B.n350 B.n191 10.6151
R1250 B.n354 B.n191 10.6151
R1251 B.n355 B.n354 10.6151
R1252 B.n356 B.n355 10.6151
R1253 B.n356 B.n189 10.6151
R1254 B.n360 B.n189 10.6151
R1255 B.n361 B.n360 10.6151
R1256 B.n362 B.n361 10.6151
R1257 B.n362 B.n187 10.6151
R1258 B.n366 B.n187 10.6151
R1259 B.n367 B.n366 10.6151
R1260 B.n368 B.n367 10.6151
R1261 B.n368 B.n185 10.6151
R1262 B.n372 B.n185 10.6151
R1263 B.n373 B.n372 10.6151
R1264 B.n374 B.n373 10.6151
R1265 B.n374 B.n183 10.6151
R1266 B.n378 B.n183 10.6151
R1267 B.n379 B.n378 10.6151
R1268 B.n380 B.n379 10.6151
R1269 B.n380 B.n181 10.6151
R1270 B.n384 B.n181 10.6151
R1271 B.n385 B.n384 10.6151
R1272 B.n386 B.n385 10.6151
R1273 B.n390 B.n389 10.6151
R1274 B.n391 B.n390 10.6151
R1275 B.n391 B.n175 10.6151
R1276 B.n395 B.n175 10.6151
R1277 B.n396 B.n395 10.6151
R1278 B.n397 B.n396 10.6151
R1279 B.n397 B.n173 10.6151
R1280 B.n401 B.n173 10.6151
R1281 B.n402 B.n401 10.6151
R1282 B.n404 B.n169 10.6151
R1283 B.n408 B.n169 10.6151
R1284 B.n409 B.n408 10.6151
R1285 B.n410 B.n409 10.6151
R1286 B.n410 B.n167 10.6151
R1287 B.n414 B.n167 10.6151
R1288 B.n415 B.n414 10.6151
R1289 B.n416 B.n415 10.6151
R1290 B.n416 B.n165 10.6151
R1291 B.n420 B.n165 10.6151
R1292 B.n421 B.n420 10.6151
R1293 B.n422 B.n421 10.6151
R1294 B.n422 B.n163 10.6151
R1295 B.n426 B.n163 10.6151
R1296 B.n427 B.n426 10.6151
R1297 B.n428 B.n427 10.6151
R1298 B.n428 B.n161 10.6151
R1299 B.n432 B.n161 10.6151
R1300 B.n433 B.n432 10.6151
R1301 B.n434 B.n433 10.6151
R1302 B.n434 B.n159 10.6151
R1303 B.n438 B.n159 10.6151
R1304 B.n439 B.n438 10.6151
R1305 B.n440 B.n439 10.6151
R1306 B.n440 B.n157 10.6151
R1307 B.n444 B.n157 10.6151
R1308 B.n445 B.n444 10.6151
R1309 B.n446 B.n445 10.6151
R1310 B.n446 B.n155 10.6151
R1311 B.n450 B.n155 10.6151
R1312 B.n451 B.n450 10.6151
R1313 B.n452 B.n451 10.6151
R1314 B.n452 B.n153 10.6151
R1315 B.n456 B.n153 10.6151
R1316 B.n457 B.n456 10.6151
R1317 B.n458 B.n457 10.6151
R1318 B.n458 B.n151 10.6151
R1319 B.n462 B.n151 10.6151
R1320 B.n463 B.n462 10.6151
R1321 B.n464 B.n463 10.6151
R1322 B.n464 B.n149 10.6151
R1323 B.n468 B.n149 10.6151
R1324 B.n469 B.n468 10.6151
R1325 B.n470 B.n469 10.6151
R1326 B.n470 B.n147 10.6151
R1327 B.n474 B.n147 10.6151
R1328 B.n475 B.n474 10.6151
R1329 B.n476 B.n475 10.6151
R1330 B.n313 B.n312 10.6151
R1331 B.n312 B.n205 10.6151
R1332 B.n308 B.n205 10.6151
R1333 B.n308 B.n307 10.6151
R1334 B.n307 B.n306 10.6151
R1335 B.n306 B.n207 10.6151
R1336 B.n302 B.n207 10.6151
R1337 B.n302 B.n301 10.6151
R1338 B.n301 B.n300 10.6151
R1339 B.n300 B.n209 10.6151
R1340 B.n296 B.n209 10.6151
R1341 B.n296 B.n295 10.6151
R1342 B.n295 B.n294 10.6151
R1343 B.n294 B.n211 10.6151
R1344 B.n290 B.n211 10.6151
R1345 B.n290 B.n289 10.6151
R1346 B.n289 B.n288 10.6151
R1347 B.n288 B.n213 10.6151
R1348 B.n284 B.n213 10.6151
R1349 B.n284 B.n283 10.6151
R1350 B.n283 B.n282 10.6151
R1351 B.n282 B.n215 10.6151
R1352 B.n278 B.n215 10.6151
R1353 B.n278 B.n277 10.6151
R1354 B.n277 B.n276 10.6151
R1355 B.n276 B.n217 10.6151
R1356 B.n272 B.n217 10.6151
R1357 B.n272 B.n271 10.6151
R1358 B.n271 B.n270 10.6151
R1359 B.n270 B.n219 10.6151
R1360 B.n266 B.n219 10.6151
R1361 B.n266 B.n265 10.6151
R1362 B.n265 B.n264 10.6151
R1363 B.n264 B.n221 10.6151
R1364 B.n260 B.n221 10.6151
R1365 B.n260 B.n259 10.6151
R1366 B.n259 B.n258 10.6151
R1367 B.n258 B.n223 10.6151
R1368 B.n254 B.n223 10.6151
R1369 B.n254 B.n253 10.6151
R1370 B.n253 B.n252 10.6151
R1371 B.n252 B.n225 10.6151
R1372 B.n248 B.n225 10.6151
R1373 B.n248 B.n247 10.6151
R1374 B.n247 B.n246 10.6151
R1375 B.n246 B.n227 10.6151
R1376 B.n242 B.n227 10.6151
R1377 B.n242 B.n241 10.6151
R1378 B.n241 B.n240 10.6151
R1379 B.n240 B.n229 10.6151
R1380 B.n236 B.n229 10.6151
R1381 B.n236 B.n235 10.6151
R1382 B.n235 B.n234 10.6151
R1383 B.n234 B.n231 10.6151
R1384 B.n231 B.n0 10.6151
R1385 B.n891 B.n1 10.6151
R1386 B.n891 B.n890 10.6151
R1387 B.n890 B.n889 10.6151
R1388 B.n889 B.n4 10.6151
R1389 B.n885 B.n4 10.6151
R1390 B.n885 B.n884 10.6151
R1391 B.n884 B.n883 10.6151
R1392 B.n883 B.n6 10.6151
R1393 B.n879 B.n6 10.6151
R1394 B.n879 B.n878 10.6151
R1395 B.n878 B.n877 10.6151
R1396 B.n877 B.n8 10.6151
R1397 B.n873 B.n8 10.6151
R1398 B.n873 B.n872 10.6151
R1399 B.n872 B.n871 10.6151
R1400 B.n871 B.n10 10.6151
R1401 B.n867 B.n10 10.6151
R1402 B.n867 B.n866 10.6151
R1403 B.n866 B.n865 10.6151
R1404 B.n865 B.n12 10.6151
R1405 B.n861 B.n12 10.6151
R1406 B.n861 B.n860 10.6151
R1407 B.n860 B.n859 10.6151
R1408 B.n859 B.n14 10.6151
R1409 B.n855 B.n14 10.6151
R1410 B.n855 B.n854 10.6151
R1411 B.n854 B.n853 10.6151
R1412 B.n853 B.n16 10.6151
R1413 B.n849 B.n16 10.6151
R1414 B.n849 B.n848 10.6151
R1415 B.n848 B.n847 10.6151
R1416 B.n847 B.n18 10.6151
R1417 B.n843 B.n18 10.6151
R1418 B.n843 B.n842 10.6151
R1419 B.n842 B.n841 10.6151
R1420 B.n841 B.n20 10.6151
R1421 B.n837 B.n20 10.6151
R1422 B.n837 B.n836 10.6151
R1423 B.n836 B.n835 10.6151
R1424 B.n835 B.n22 10.6151
R1425 B.n831 B.n22 10.6151
R1426 B.n831 B.n830 10.6151
R1427 B.n830 B.n829 10.6151
R1428 B.n829 B.n24 10.6151
R1429 B.n825 B.n24 10.6151
R1430 B.n825 B.n824 10.6151
R1431 B.n824 B.n823 10.6151
R1432 B.n823 B.n26 10.6151
R1433 B.n819 B.n26 10.6151
R1434 B.n819 B.n818 10.6151
R1435 B.n818 B.n817 10.6151
R1436 B.n817 B.n28 10.6151
R1437 B.n813 B.n28 10.6151
R1438 B.n813 B.n812 10.6151
R1439 B.n812 B.n811 10.6151
R1440 B.n58 B.n54 9.36635
R1441 B.n721 B.n720 9.36635
R1442 B.n386 B.n179 9.36635
R1443 B.n404 B.n403 9.36635
R1444 B.n895 B.n0 2.81026
R1445 B.n895 B.n1 2.81026
R1446 B.n735 B.n58 1.24928
R1447 B.n722 B.n721 1.24928
R1448 B.n389 B.n179 1.24928
R1449 B.n403 B.n402 1.24928
R1450 VP.n16 VP.n13 161.3
R1451 VP.n18 VP.n17 161.3
R1452 VP.n19 VP.n12 161.3
R1453 VP.n21 VP.n20 161.3
R1454 VP.n22 VP.n11 161.3
R1455 VP.n24 VP.n23 161.3
R1456 VP.n25 VP.n10 161.3
R1457 VP.n27 VP.n26 161.3
R1458 VP.n56 VP.n55 161.3
R1459 VP.n54 VP.n1 161.3
R1460 VP.n53 VP.n52 161.3
R1461 VP.n51 VP.n2 161.3
R1462 VP.n50 VP.n49 161.3
R1463 VP.n48 VP.n3 161.3
R1464 VP.n47 VP.n46 161.3
R1465 VP.n45 VP.n4 161.3
R1466 VP.n44 VP.n43 161.3
R1467 VP.n42 VP.n5 161.3
R1468 VP.n41 VP.n40 161.3
R1469 VP.n39 VP.n6 161.3
R1470 VP.n38 VP.n37 161.3
R1471 VP.n36 VP.n7 161.3
R1472 VP.n35 VP.n34 161.3
R1473 VP.n33 VP.n8 161.3
R1474 VP.n32 VP.n31 161.3
R1475 VP.n15 VP.t0 127.058
R1476 VP.n43 VP.t3 94.1391
R1477 VP.n30 VP.t5 94.1391
R1478 VP.n0 VP.t1 94.1391
R1479 VP.n14 VP.t4 94.1391
R1480 VP.n9 VP.t2 94.1391
R1481 VP.n30 VP.n29 87.1314
R1482 VP.n57 VP.n0 87.1314
R1483 VP.n28 VP.n9 87.1314
R1484 VP.n29 VP.n28 55.0902
R1485 VP.n15 VP.n14 50.484
R1486 VP.n37 VP.n36 43.4072
R1487 VP.n49 VP.n2 43.4072
R1488 VP.n20 VP.n11 43.4072
R1489 VP.n37 VP.n6 37.5796
R1490 VP.n49 VP.n48 37.5796
R1491 VP.n20 VP.n19 37.5796
R1492 VP.n31 VP.n8 24.4675
R1493 VP.n35 VP.n8 24.4675
R1494 VP.n36 VP.n35 24.4675
R1495 VP.n41 VP.n6 24.4675
R1496 VP.n42 VP.n41 24.4675
R1497 VP.n43 VP.n42 24.4675
R1498 VP.n43 VP.n4 24.4675
R1499 VP.n47 VP.n4 24.4675
R1500 VP.n48 VP.n47 24.4675
R1501 VP.n53 VP.n2 24.4675
R1502 VP.n54 VP.n53 24.4675
R1503 VP.n55 VP.n54 24.4675
R1504 VP.n24 VP.n11 24.4675
R1505 VP.n25 VP.n24 24.4675
R1506 VP.n26 VP.n25 24.4675
R1507 VP.n14 VP.n13 24.4675
R1508 VP.n18 VP.n13 24.4675
R1509 VP.n19 VP.n18 24.4675
R1510 VP.n31 VP.n30 2.93654
R1511 VP.n55 VP.n0 2.93654
R1512 VP.n26 VP.n9 2.93654
R1513 VP.n16 VP.n15 2.46264
R1514 VP.n28 VP.n27 0.354971
R1515 VP.n32 VP.n29 0.354971
R1516 VP.n57 VP.n56 0.354971
R1517 VP VP.n57 0.26696
R1518 VP.n17 VP.n16 0.189894
R1519 VP.n17 VP.n12 0.189894
R1520 VP.n21 VP.n12 0.189894
R1521 VP.n22 VP.n21 0.189894
R1522 VP.n23 VP.n22 0.189894
R1523 VP.n23 VP.n10 0.189894
R1524 VP.n27 VP.n10 0.189894
R1525 VP.n33 VP.n32 0.189894
R1526 VP.n34 VP.n33 0.189894
R1527 VP.n34 VP.n7 0.189894
R1528 VP.n38 VP.n7 0.189894
R1529 VP.n39 VP.n38 0.189894
R1530 VP.n40 VP.n39 0.189894
R1531 VP.n40 VP.n5 0.189894
R1532 VP.n44 VP.n5 0.189894
R1533 VP.n45 VP.n44 0.189894
R1534 VP.n46 VP.n45 0.189894
R1535 VP.n46 VP.n3 0.189894
R1536 VP.n50 VP.n3 0.189894
R1537 VP.n51 VP.n50 0.189894
R1538 VP.n52 VP.n51 0.189894
R1539 VP.n52 VP.n1 0.189894
R1540 VP.n56 VP.n1 0.189894
R1541 VDD1 VDD1.t5 74.8925
R1542 VDD1.n1 VDD1.t0 74.7787
R1543 VDD1.n1 VDD1.n0 70.798
R1544 VDD1.n3 VDD1.n2 69.9783
R1545 VDD1.n3 VDD1.n1 49.9837
R1546 VDD1.n2 VDD1.t1 2.23145
R1547 VDD1.n2 VDD1.t3 2.23145
R1548 VDD1.n0 VDD1.t2 2.23145
R1549 VDD1.n0 VDD1.t4 2.23145
R1550 VDD1 VDD1.n3 0.81731
C0 B VDD2 2.6952f
C1 VDD2 VTAIL 9.00945f
C2 B VN 1.43582f
C3 VN VTAIL 8.88195f
C4 B VDD1 2.59401f
C5 VDD1 VTAIL 8.95053f
C6 B w_n4218_n3882# 11.9573f
C7 w_n4218_n3882# VTAIL 3.41433f
C8 VP B 2.35725f
C9 VP VTAIL 8.89663f
C10 VDD2 VN 8.573701f
C11 VDD2 VDD1 1.84709f
C12 w_n4218_n3882# VDD2 2.85778f
C13 VP VDD2 0.553725f
C14 VN VDD1 0.152134f
C15 w_n4218_n3882# VN 8.319519f
C16 w_n4218_n3882# VDD1 2.73658f
C17 VP VN 8.50287f
C18 VP VDD1 8.97235f
C19 B VTAIL 4.72523f
C20 VP w_n4218_n3882# 8.868f
C21 VDD2 VSUBS 2.28957f
C22 VDD1 VSUBS 2.87633f
C23 VTAIL VSUBS 1.497401f
C24 VN VSUBS 7.026299f
C25 VP VSUBS 3.900581f
C26 B VSUBS 5.970177f
C27 w_n4218_n3882# VSUBS 0.200895p
C28 VDD1.t5 VSUBS 3.40308f
C29 VDD1.t0 VSUBS 3.40141f
C30 VDD1.t2 VSUBS 0.322538f
C31 VDD1.t4 VSUBS 0.322538f
C32 VDD1.n0 VSUBS 2.59931f
C33 VDD1.n1 VSUBS 4.81024f
C34 VDD1.t1 VSUBS 0.322538f
C35 VDD1.t3 VSUBS 0.322538f
C36 VDD1.n2 VSUBS 2.58827f
C37 VDD1.n3 VSUBS 4.02128f
C38 VP.t1 VSUBS 3.86489f
C39 VP.n0 VSUBS 1.4382f
C40 VP.n1 VSUBS 0.025971f
C41 VP.n2 VSUBS 0.050694f
C42 VP.n3 VSUBS 0.025971f
C43 VP.n4 VSUBS 0.048402f
C44 VP.n5 VSUBS 0.025971f
C45 VP.t3 VSUBS 3.86489f
C46 VP.n6 VSUBS 0.052236f
C47 VP.n7 VSUBS 0.025971f
C48 VP.n8 VSUBS 0.048402f
C49 VP.t2 VSUBS 3.86489f
C50 VP.n9 VSUBS 1.4382f
C51 VP.n10 VSUBS 0.025971f
C52 VP.n11 VSUBS 0.050694f
C53 VP.n12 VSUBS 0.025971f
C54 VP.n13 VSUBS 0.048402f
C55 VP.t0 VSUBS 4.26585f
C56 VP.t4 VSUBS 3.86489f
C57 VP.n14 VSUBS 1.44883f
C58 VP.n15 VSUBS 1.37536f
C59 VP.n16 VSUBS 0.331573f
C60 VP.n17 VSUBS 0.025971f
C61 VP.n18 VSUBS 0.048402f
C62 VP.n19 VSUBS 0.052236f
C63 VP.n20 VSUBS 0.021296f
C64 VP.n21 VSUBS 0.025971f
C65 VP.n22 VSUBS 0.025971f
C66 VP.n23 VSUBS 0.025971f
C67 VP.n24 VSUBS 0.048402f
C68 VP.n25 VSUBS 0.048402f
C69 VP.n26 VSUBS 0.027373f
C70 VP.n27 VSUBS 0.041916f
C71 VP.n28 VSUBS 1.70898f
C72 VP.n29 VSUBS 1.72592f
C73 VP.t5 VSUBS 3.86489f
C74 VP.n30 VSUBS 1.4382f
C75 VP.n31 VSUBS 0.027373f
C76 VP.n32 VSUBS 0.041916f
C77 VP.n33 VSUBS 0.025971f
C78 VP.n34 VSUBS 0.025971f
C79 VP.n35 VSUBS 0.048402f
C80 VP.n36 VSUBS 0.050694f
C81 VP.n37 VSUBS 0.021296f
C82 VP.n38 VSUBS 0.025971f
C83 VP.n39 VSUBS 0.025971f
C84 VP.n40 VSUBS 0.025971f
C85 VP.n41 VSUBS 0.048402f
C86 VP.n42 VSUBS 0.048402f
C87 VP.n43 VSUBS 1.36686f
C88 VP.n44 VSUBS 0.025971f
C89 VP.n45 VSUBS 0.025971f
C90 VP.n46 VSUBS 0.025971f
C91 VP.n47 VSUBS 0.048402f
C92 VP.n48 VSUBS 0.052236f
C93 VP.n49 VSUBS 0.021296f
C94 VP.n50 VSUBS 0.025971f
C95 VP.n51 VSUBS 0.025971f
C96 VP.n52 VSUBS 0.025971f
C97 VP.n53 VSUBS 0.048402f
C98 VP.n54 VSUBS 0.048402f
C99 VP.n55 VSUBS 0.027373f
C100 VP.n56 VSUBS 0.041916f
C101 VP.n57 VSUBS 0.078731f
C102 B.n0 VSUBS 0.00493f
C103 B.n1 VSUBS 0.00493f
C104 B.n2 VSUBS 0.007796f
C105 B.n3 VSUBS 0.007796f
C106 B.n4 VSUBS 0.007796f
C107 B.n5 VSUBS 0.007796f
C108 B.n6 VSUBS 0.007796f
C109 B.n7 VSUBS 0.007796f
C110 B.n8 VSUBS 0.007796f
C111 B.n9 VSUBS 0.007796f
C112 B.n10 VSUBS 0.007796f
C113 B.n11 VSUBS 0.007796f
C114 B.n12 VSUBS 0.007796f
C115 B.n13 VSUBS 0.007796f
C116 B.n14 VSUBS 0.007796f
C117 B.n15 VSUBS 0.007796f
C118 B.n16 VSUBS 0.007796f
C119 B.n17 VSUBS 0.007796f
C120 B.n18 VSUBS 0.007796f
C121 B.n19 VSUBS 0.007796f
C122 B.n20 VSUBS 0.007796f
C123 B.n21 VSUBS 0.007796f
C124 B.n22 VSUBS 0.007796f
C125 B.n23 VSUBS 0.007796f
C126 B.n24 VSUBS 0.007796f
C127 B.n25 VSUBS 0.007796f
C128 B.n26 VSUBS 0.007796f
C129 B.n27 VSUBS 0.007796f
C130 B.n28 VSUBS 0.007796f
C131 B.n29 VSUBS 0.007796f
C132 B.n30 VSUBS 0.017936f
C133 B.n31 VSUBS 0.007796f
C134 B.n32 VSUBS 0.007796f
C135 B.n33 VSUBS 0.007796f
C136 B.n34 VSUBS 0.007796f
C137 B.n35 VSUBS 0.007796f
C138 B.n36 VSUBS 0.007796f
C139 B.n37 VSUBS 0.007796f
C140 B.n38 VSUBS 0.007796f
C141 B.n39 VSUBS 0.007796f
C142 B.n40 VSUBS 0.007796f
C143 B.n41 VSUBS 0.007796f
C144 B.n42 VSUBS 0.007796f
C145 B.n43 VSUBS 0.007796f
C146 B.n44 VSUBS 0.007796f
C147 B.n45 VSUBS 0.007796f
C148 B.n46 VSUBS 0.007796f
C149 B.n47 VSUBS 0.007796f
C150 B.n48 VSUBS 0.007796f
C151 B.n49 VSUBS 0.007796f
C152 B.n50 VSUBS 0.007796f
C153 B.n51 VSUBS 0.007796f
C154 B.n52 VSUBS 0.007796f
C155 B.n53 VSUBS 0.007796f
C156 B.n54 VSUBS 0.007338f
C157 B.n55 VSUBS 0.007796f
C158 B.t5 VSUBS 0.538881f
C159 B.t4 VSUBS 0.569483f
C160 B.t3 VSUBS 2.78989f
C161 B.n56 VSUBS 0.336758f
C162 B.n57 VSUBS 0.08534f
C163 B.n58 VSUBS 0.018063f
C164 B.n59 VSUBS 0.007796f
C165 B.n60 VSUBS 0.007796f
C166 B.n61 VSUBS 0.007796f
C167 B.n62 VSUBS 0.007796f
C168 B.t8 VSUBS 0.538867f
C169 B.t7 VSUBS 0.569472f
C170 B.t6 VSUBS 2.78989f
C171 B.n63 VSUBS 0.33677f
C172 B.n64 VSUBS 0.085354f
C173 B.n65 VSUBS 0.007796f
C174 B.n66 VSUBS 0.007796f
C175 B.n67 VSUBS 0.007796f
C176 B.n68 VSUBS 0.007796f
C177 B.n69 VSUBS 0.007796f
C178 B.n70 VSUBS 0.007796f
C179 B.n71 VSUBS 0.007796f
C180 B.n72 VSUBS 0.007796f
C181 B.n73 VSUBS 0.007796f
C182 B.n74 VSUBS 0.007796f
C183 B.n75 VSUBS 0.007796f
C184 B.n76 VSUBS 0.007796f
C185 B.n77 VSUBS 0.007796f
C186 B.n78 VSUBS 0.007796f
C187 B.n79 VSUBS 0.007796f
C188 B.n80 VSUBS 0.007796f
C189 B.n81 VSUBS 0.007796f
C190 B.n82 VSUBS 0.007796f
C191 B.n83 VSUBS 0.007796f
C192 B.n84 VSUBS 0.007796f
C193 B.n85 VSUBS 0.007796f
C194 B.n86 VSUBS 0.007796f
C195 B.n87 VSUBS 0.007796f
C196 B.n88 VSUBS 0.007796f
C197 B.n89 VSUBS 0.018126f
C198 B.n90 VSUBS 0.007796f
C199 B.n91 VSUBS 0.007796f
C200 B.n92 VSUBS 0.007796f
C201 B.n93 VSUBS 0.007796f
C202 B.n94 VSUBS 0.007796f
C203 B.n95 VSUBS 0.007796f
C204 B.n96 VSUBS 0.007796f
C205 B.n97 VSUBS 0.007796f
C206 B.n98 VSUBS 0.007796f
C207 B.n99 VSUBS 0.007796f
C208 B.n100 VSUBS 0.007796f
C209 B.n101 VSUBS 0.007796f
C210 B.n102 VSUBS 0.007796f
C211 B.n103 VSUBS 0.007796f
C212 B.n104 VSUBS 0.007796f
C213 B.n105 VSUBS 0.007796f
C214 B.n106 VSUBS 0.007796f
C215 B.n107 VSUBS 0.007796f
C216 B.n108 VSUBS 0.007796f
C217 B.n109 VSUBS 0.007796f
C218 B.n110 VSUBS 0.007796f
C219 B.n111 VSUBS 0.007796f
C220 B.n112 VSUBS 0.007796f
C221 B.n113 VSUBS 0.007796f
C222 B.n114 VSUBS 0.007796f
C223 B.n115 VSUBS 0.007796f
C224 B.n116 VSUBS 0.007796f
C225 B.n117 VSUBS 0.007796f
C226 B.n118 VSUBS 0.007796f
C227 B.n119 VSUBS 0.007796f
C228 B.n120 VSUBS 0.007796f
C229 B.n121 VSUBS 0.007796f
C230 B.n122 VSUBS 0.007796f
C231 B.n123 VSUBS 0.007796f
C232 B.n124 VSUBS 0.007796f
C233 B.n125 VSUBS 0.007796f
C234 B.n126 VSUBS 0.007796f
C235 B.n127 VSUBS 0.007796f
C236 B.n128 VSUBS 0.007796f
C237 B.n129 VSUBS 0.007796f
C238 B.n130 VSUBS 0.007796f
C239 B.n131 VSUBS 0.007796f
C240 B.n132 VSUBS 0.007796f
C241 B.n133 VSUBS 0.007796f
C242 B.n134 VSUBS 0.007796f
C243 B.n135 VSUBS 0.007796f
C244 B.n136 VSUBS 0.007796f
C245 B.n137 VSUBS 0.007796f
C246 B.n138 VSUBS 0.007796f
C247 B.n139 VSUBS 0.007796f
C248 B.n140 VSUBS 0.007796f
C249 B.n141 VSUBS 0.007796f
C250 B.n142 VSUBS 0.007796f
C251 B.n143 VSUBS 0.007796f
C252 B.n144 VSUBS 0.007796f
C253 B.n145 VSUBS 0.017148f
C254 B.n146 VSUBS 0.007796f
C255 B.n147 VSUBS 0.007796f
C256 B.n148 VSUBS 0.007796f
C257 B.n149 VSUBS 0.007796f
C258 B.n150 VSUBS 0.007796f
C259 B.n151 VSUBS 0.007796f
C260 B.n152 VSUBS 0.007796f
C261 B.n153 VSUBS 0.007796f
C262 B.n154 VSUBS 0.007796f
C263 B.n155 VSUBS 0.007796f
C264 B.n156 VSUBS 0.007796f
C265 B.n157 VSUBS 0.007796f
C266 B.n158 VSUBS 0.007796f
C267 B.n159 VSUBS 0.007796f
C268 B.n160 VSUBS 0.007796f
C269 B.n161 VSUBS 0.007796f
C270 B.n162 VSUBS 0.007796f
C271 B.n163 VSUBS 0.007796f
C272 B.n164 VSUBS 0.007796f
C273 B.n165 VSUBS 0.007796f
C274 B.n166 VSUBS 0.007796f
C275 B.n167 VSUBS 0.007796f
C276 B.n168 VSUBS 0.007796f
C277 B.n169 VSUBS 0.007796f
C278 B.n170 VSUBS 0.007796f
C279 B.t10 VSUBS 0.538867f
C280 B.t11 VSUBS 0.569472f
C281 B.t9 VSUBS 2.78989f
C282 B.n171 VSUBS 0.33677f
C283 B.n172 VSUBS 0.085354f
C284 B.n173 VSUBS 0.007796f
C285 B.n174 VSUBS 0.007796f
C286 B.n175 VSUBS 0.007796f
C287 B.n176 VSUBS 0.007796f
C288 B.t1 VSUBS 0.538881f
C289 B.t2 VSUBS 0.569483f
C290 B.t0 VSUBS 2.78989f
C291 B.n177 VSUBS 0.336758f
C292 B.n178 VSUBS 0.08534f
C293 B.n179 VSUBS 0.018063f
C294 B.n180 VSUBS 0.007796f
C295 B.n181 VSUBS 0.007796f
C296 B.n182 VSUBS 0.007796f
C297 B.n183 VSUBS 0.007796f
C298 B.n184 VSUBS 0.007796f
C299 B.n185 VSUBS 0.007796f
C300 B.n186 VSUBS 0.007796f
C301 B.n187 VSUBS 0.007796f
C302 B.n188 VSUBS 0.007796f
C303 B.n189 VSUBS 0.007796f
C304 B.n190 VSUBS 0.007796f
C305 B.n191 VSUBS 0.007796f
C306 B.n192 VSUBS 0.007796f
C307 B.n193 VSUBS 0.007796f
C308 B.n194 VSUBS 0.007796f
C309 B.n195 VSUBS 0.007796f
C310 B.n196 VSUBS 0.007796f
C311 B.n197 VSUBS 0.007796f
C312 B.n198 VSUBS 0.007796f
C313 B.n199 VSUBS 0.007796f
C314 B.n200 VSUBS 0.007796f
C315 B.n201 VSUBS 0.007796f
C316 B.n202 VSUBS 0.007796f
C317 B.n203 VSUBS 0.007796f
C318 B.n204 VSUBS 0.017148f
C319 B.n205 VSUBS 0.007796f
C320 B.n206 VSUBS 0.007796f
C321 B.n207 VSUBS 0.007796f
C322 B.n208 VSUBS 0.007796f
C323 B.n209 VSUBS 0.007796f
C324 B.n210 VSUBS 0.007796f
C325 B.n211 VSUBS 0.007796f
C326 B.n212 VSUBS 0.007796f
C327 B.n213 VSUBS 0.007796f
C328 B.n214 VSUBS 0.007796f
C329 B.n215 VSUBS 0.007796f
C330 B.n216 VSUBS 0.007796f
C331 B.n217 VSUBS 0.007796f
C332 B.n218 VSUBS 0.007796f
C333 B.n219 VSUBS 0.007796f
C334 B.n220 VSUBS 0.007796f
C335 B.n221 VSUBS 0.007796f
C336 B.n222 VSUBS 0.007796f
C337 B.n223 VSUBS 0.007796f
C338 B.n224 VSUBS 0.007796f
C339 B.n225 VSUBS 0.007796f
C340 B.n226 VSUBS 0.007796f
C341 B.n227 VSUBS 0.007796f
C342 B.n228 VSUBS 0.007796f
C343 B.n229 VSUBS 0.007796f
C344 B.n230 VSUBS 0.007796f
C345 B.n231 VSUBS 0.007796f
C346 B.n232 VSUBS 0.007796f
C347 B.n233 VSUBS 0.007796f
C348 B.n234 VSUBS 0.007796f
C349 B.n235 VSUBS 0.007796f
C350 B.n236 VSUBS 0.007796f
C351 B.n237 VSUBS 0.007796f
C352 B.n238 VSUBS 0.007796f
C353 B.n239 VSUBS 0.007796f
C354 B.n240 VSUBS 0.007796f
C355 B.n241 VSUBS 0.007796f
C356 B.n242 VSUBS 0.007796f
C357 B.n243 VSUBS 0.007796f
C358 B.n244 VSUBS 0.007796f
C359 B.n245 VSUBS 0.007796f
C360 B.n246 VSUBS 0.007796f
C361 B.n247 VSUBS 0.007796f
C362 B.n248 VSUBS 0.007796f
C363 B.n249 VSUBS 0.007796f
C364 B.n250 VSUBS 0.007796f
C365 B.n251 VSUBS 0.007796f
C366 B.n252 VSUBS 0.007796f
C367 B.n253 VSUBS 0.007796f
C368 B.n254 VSUBS 0.007796f
C369 B.n255 VSUBS 0.007796f
C370 B.n256 VSUBS 0.007796f
C371 B.n257 VSUBS 0.007796f
C372 B.n258 VSUBS 0.007796f
C373 B.n259 VSUBS 0.007796f
C374 B.n260 VSUBS 0.007796f
C375 B.n261 VSUBS 0.007796f
C376 B.n262 VSUBS 0.007796f
C377 B.n263 VSUBS 0.007796f
C378 B.n264 VSUBS 0.007796f
C379 B.n265 VSUBS 0.007796f
C380 B.n266 VSUBS 0.007796f
C381 B.n267 VSUBS 0.007796f
C382 B.n268 VSUBS 0.007796f
C383 B.n269 VSUBS 0.007796f
C384 B.n270 VSUBS 0.007796f
C385 B.n271 VSUBS 0.007796f
C386 B.n272 VSUBS 0.007796f
C387 B.n273 VSUBS 0.007796f
C388 B.n274 VSUBS 0.007796f
C389 B.n275 VSUBS 0.007796f
C390 B.n276 VSUBS 0.007796f
C391 B.n277 VSUBS 0.007796f
C392 B.n278 VSUBS 0.007796f
C393 B.n279 VSUBS 0.007796f
C394 B.n280 VSUBS 0.007796f
C395 B.n281 VSUBS 0.007796f
C396 B.n282 VSUBS 0.007796f
C397 B.n283 VSUBS 0.007796f
C398 B.n284 VSUBS 0.007796f
C399 B.n285 VSUBS 0.007796f
C400 B.n286 VSUBS 0.007796f
C401 B.n287 VSUBS 0.007796f
C402 B.n288 VSUBS 0.007796f
C403 B.n289 VSUBS 0.007796f
C404 B.n290 VSUBS 0.007796f
C405 B.n291 VSUBS 0.007796f
C406 B.n292 VSUBS 0.007796f
C407 B.n293 VSUBS 0.007796f
C408 B.n294 VSUBS 0.007796f
C409 B.n295 VSUBS 0.007796f
C410 B.n296 VSUBS 0.007796f
C411 B.n297 VSUBS 0.007796f
C412 B.n298 VSUBS 0.007796f
C413 B.n299 VSUBS 0.007796f
C414 B.n300 VSUBS 0.007796f
C415 B.n301 VSUBS 0.007796f
C416 B.n302 VSUBS 0.007796f
C417 B.n303 VSUBS 0.007796f
C418 B.n304 VSUBS 0.007796f
C419 B.n305 VSUBS 0.007796f
C420 B.n306 VSUBS 0.007796f
C421 B.n307 VSUBS 0.007796f
C422 B.n308 VSUBS 0.007796f
C423 B.n309 VSUBS 0.007796f
C424 B.n310 VSUBS 0.007796f
C425 B.n311 VSUBS 0.007796f
C426 B.n312 VSUBS 0.007796f
C427 B.n313 VSUBS 0.017148f
C428 B.n314 VSUBS 0.017936f
C429 B.n315 VSUBS 0.017936f
C430 B.n316 VSUBS 0.007796f
C431 B.n317 VSUBS 0.007796f
C432 B.n318 VSUBS 0.007796f
C433 B.n319 VSUBS 0.007796f
C434 B.n320 VSUBS 0.007796f
C435 B.n321 VSUBS 0.007796f
C436 B.n322 VSUBS 0.007796f
C437 B.n323 VSUBS 0.007796f
C438 B.n324 VSUBS 0.007796f
C439 B.n325 VSUBS 0.007796f
C440 B.n326 VSUBS 0.007796f
C441 B.n327 VSUBS 0.007796f
C442 B.n328 VSUBS 0.007796f
C443 B.n329 VSUBS 0.007796f
C444 B.n330 VSUBS 0.007796f
C445 B.n331 VSUBS 0.007796f
C446 B.n332 VSUBS 0.007796f
C447 B.n333 VSUBS 0.007796f
C448 B.n334 VSUBS 0.007796f
C449 B.n335 VSUBS 0.007796f
C450 B.n336 VSUBS 0.007796f
C451 B.n337 VSUBS 0.007796f
C452 B.n338 VSUBS 0.007796f
C453 B.n339 VSUBS 0.007796f
C454 B.n340 VSUBS 0.007796f
C455 B.n341 VSUBS 0.007796f
C456 B.n342 VSUBS 0.007796f
C457 B.n343 VSUBS 0.007796f
C458 B.n344 VSUBS 0.007796f
C459 B.n345 VSUBS 0.007796f
C460 B.n346 VSUBS 0.007796f
C461 B.n347 VSUBS 0.007796f
C462 B.n348 VSUBS 0.007796f
C463 B.n349 VSUBS 0.007796f
C464 B.n350 VSUBS 0.007796f
C465 B.n351 VSUBS 0.007796f
C466 B.n352 VSUBS 0.007796f
C467 B.n353 VSUBS 0.007796f
C468 B.n354 VSUBS 0.007796f
C469 B.n355 VSUBS 0.007796f
C470 B.n356 VSUBS 0.007796f
C471 B.n357 VSUBS 0.007796f
C472 B.n358 VSUBS 0.007796f
C473 B.n359 VSUBS 0.007796f
C474 B.n360 VSUBS 0.007796f
C475 B.n361 VSUBS 0.007796f
C476 B.n362 VSUBS 0.007796f
C477 B.n363 VSUBS 0.007796f
C478 B.n364 VSUBS 0.007796f
C479 B.n365 VSUBS 0.007796f
C480 B.n366 VSUBS 0.007796f
C481 B.n367 VSUBS 0.007796f
C482 B.n368 VSUBS 0.007796f
C483 B.n369 VSUBS 0.007796f
C484 B.n370 VSUBS 0.007796f
C485 B.n371 VSUBS 0.007796f
C486 B.n372 VSUBS 0.007796f
C487 B.n373 VSUBS 0.007796f
C488 B.n374 VSUBS 0.007796f
C489 B.n375 VSUBS 0.007796f
C490 B.n376 VSUBS 0.007796f
C491 B.n377 VSUBS 0.007796f
C492 B.n378 VSUBS 0.007796f
C493 B.n379 VSUBS 0.007796f
C494 B.n380 VSUBS 0.007796f
C495 B.n381 VSUBS 0.007796f
C496 B.n382 VSUBS 0.007796f
C497 B.n383 VSUBS 0.007796f
C498 B.n384 VSUBS 0.007796f
C499 B.n385 VSUBS 0.007796f
C500 B.n386 VSUBS 0.007338f
C501 B.n387 VSUBS 0.007796f
C502 B.n388 VSUBS 0.007796f
C503 B.n389 VSUBS 0.004357f
C504 B.n390 VSUBS 0.007796f
C505 B.n391 VSUBS 0.007796f
C506 B.n392 VSUBS 0.007796f
C507 B.n393 VSUBS 0.007796f
C508 B.n394 VSUBS 0.007796f
C509 B.n395 VSUBS 0.007796f
C510 B.n396 VSUBS 0.007796f
C511 B.n397 VSUBS 0.007796f
C512 B.n398 VSUBS 0.007796f
C513 B.n399 VSUBS 0.007796f
C514 B.n400 VSUBS 0.007796f
C515 B.n401 VSUBS 0.007796f
C516 B.n402 VSUBS 0.004357f
C517 B.n403 VSUBS 0.018063f
C518 B.n404 VSUBS 0.007338f
C519 B.n405 VSUBS 0.007796f
C520 B.n406 VSUBS 0.007796f
C521 B.n407 VSUBS 0.007796f
C522 B.n408 VSUBS 0.007796f
C523 B.n409 VSUBS 0.007796f
C524 B.n410 VSUBS 0.007796f
C525 B.n411 VSUBS 0.007796f
C526 B.n412 VSUBS 0.007796f
C527 B.n413 VSUBS 0.007796f
C528 B.n414 VSUBS 0.007796f
C529 B.n415 VSUBS 0.007796f
C530 B.n416 VSUBS 0.007796f
C531 B.n417 VSUBS 0.007796f
C532 B.n418 VSUBS 0.007796f
C533 B.n419 VSUBS 0.007796f
C534 B.n420 VSUBS 0.007796f
C535 B.n421 VSUBS 0.007796f
C536 B.n422 VSUBS 0.007796f
C537 B.n423 VSUBS 0.007796f
C538 B.n424 VSUBS 0.007796f
C539 B.n425 VSUBS 0.007796f
C540 B.n426 VSUBS 0.007796f
C541 B.n427 VSUBS 0.007796f
C542 B.n428 VSUBS 0.007796f
C543 B.n429 VSUBS 0.007796f
C544 B.n430 VSUBS 0.007796f
C545 B.n431 VSUBS 0.007796f
C546 B.n432 VSUBS 0.007796f
C547 B.n433 VSUBS 0.007796f
C548 B.n434 VSUBS 0.007796f
C549 B.n435 VSUBS 0.007796f
C550 B.n436 VSUBS 0.007796f
C551 B.n437 VSUBS 0.007796f
C552 B.n438 VSUBS 0.007796f
C553 B.n439 VSUBS 0.007796f
C554 B.n440 VSUBS 0.007796f
C555 B.n441 VSUBS 0.007796f
C556 B.n442 VSUBS 0.007796f
C557 B.n443 VSUBS 0.007796f
C558 B.n444 VSUBS 0.007796f
C559 B.n445 VSUBS 0.007796f
C560 B.n446 VSUBS 0.007796f
C561 B.n447 VSUBS 0.007796f
C562 B.n448 VSUBS 0.007796f
C563 B.n449 VSUBS 0.007796f
C564 B.n450 VSUBS 0.007796f
C565 B.n451 VSUBS 0.007796f
C566 B.n452 VSUBS 0.007796f
C567 B.n453 VSUBS 0.007796f
C568 B.n454 VSUBS 0.007796f
C569 B.n455 VSUBS 0.007796f
C570 B.n456 VSUBS 0.007796f
C571 B.n457 VSUBS 0.007796f
C572 B.n458 VSUBS 0.007796f
C573 B.n459 VSUBS 0.007796f
C574 B.n460 VSUBS 0.007796f
C575 B.n461 VSUBS 0.007796f
C576 B.n462 VSUBS 0.007796f
C577 B.n463 VSUBS 0.007796f
C578 B.n464 VSUBS 0.007796f
C579 B.n465 VSUBS 0.007796f
C580 B.n466 VSUBS 0.007796f
C581 B.n467 VSUBS 0.007796f
C582 B.n468 VSUBS 0.007796f
C583 B.n469 VSUBS 0.007796f
C584 B.n470 VSUBS 0.007796f
C585 B.n471 VSUBS 0.007796f
C586 B.n472 VSUBS 0.007796f
C587 B.n473 VSUBS 0.007796f
C588 B.n474 VSUBS 0.007796f
C589 B.n475 VSUBS 0.007796f
C590 B.n476 VSUBS 0.017936f
C591 B.n477 VSUBS 0.017936f
C592 B.n478 VSUBS 0.017148f
C593 B.n479 VSUBS 0.007796f
C594 B.n480 VSUBS 0.007796f
C595 B.n481 VSUBS 0.007796f
C596 B.n482 VSUBS 0.007796f
C597 B.n483 VSUBS 0.007796f
C598 B.n484 VSUBS 0.007796f
C599 B.n485 VSUBS 0.007796f
C600 B.n486 VSUBS 0.007796f
C601 B.n487 VSUBS 0.007796f
C602 B.n488 VSUBS 0.007796f
C603 B.n489 VSUBS 0.007796f
C604 B.n490 VSUBS 0.007796f
C605 B.n491 VSUBS 0.007796f
C606 B.n492 VSUBS 0.007796f
C607 B.n493 VSUBS 0.007796f
C608 B.n494 VSUBS 0.007796f
C609 B.n495 VSUBS 0.007796f
C610 B.n496 VSUBS 0.007796f
C611 B.n497 VSUBS 0.007796f
C612 B.n498 VSUBS 0.007796f
C613 B.n499 VSUBS 0.007796f
C614 B.n500 VSUBS 0.007796f
C615 B.n501 VSUBS 0.007796f
C616 B.n502 VSUBS 0.007796f
C617 B.n503 VSUBS 0.007796f
C618 B.n504 VSUBS 0.007796f
C619 B.n505 VSUBS 0.007796f
C620 B.n506 VSUBS 0.007796f
C621 B.n507 VSUBS 0.007796f
C622 B.n508 VSUBS 0.007796f
C623 B.n509 VSUBS 0.007796f
C624 B.n510 VSUBS 0.007796f
C625 B.n511 VSUBS 0.007796f
C626 B.n512 VSUBS 0.007796f
C627 B.n513 VSUBS 0.007796f
C628 B.n514 VSUBS 0.007796f
C629 B.n515 VSUBS 0.007796f
C630 B.n516 VSUBS 0.007796f
C631 B.n517 VSUBS 0.007796f
C632 B.n518 VSUBS 0.007796f
C633 B.n519 VSUBS 0.007796f
C634 B.n520 VSUBS 0.007796f
C635 B.n521 VSUBS 0.007796f
C636 B.n522 VSUBS 0.007796f
C637 B.n523 VSUBS 0.007796f
C638 B.n524 VSUBS 0.007796f
C639 B.n525 VSUBS 0.007796f
C640 B.n526 VSUBS 0.007796f
C641 B.n527 VSUBS 0.007796f
C642 B.n528 VSUBS 0.007796f
C643 B.n529 VSUBS 0.007796f
C644 B.n530 VSUBS 0.007796f
C645 B.n531 VSUBS 0.007796f
C646 B.n532 VSUBS 0.007796f
C647 B.n533 VSUBS 0.007796f
C648 B.n534 VSUBS 0.007796f
C649 B.n535 VSUBS 0.007796f
C650 B.n536 VSUBS 0.007796f
C651 B.n537 VSUBS 0.007796f
C652 B.n538 VSUBS 0.007796f
C653 B.n539 VSUBS 0.007796f
C654 B.n540 VSUBS 0.007796f
C655 B.n541 VSUBS 0.007796f
C656 B.n542 VSUBS 0.007796f
C657 B.n543 VSUBS 0.007796f
C658 B.n544 VSUBS 0.007796f
C659 B.n545 VSUBS 0.007796f
C660 B.n546 VSUBS 0.007796f
C661 B.n547 VSUBS 0.007796f
C662 B.n548 VSUBS 0.007796f
C663 B.n549 VSUBS 0.007796f
C664 B.n550 VSUBS 0.007796f
C665 B.n551 VSUBS 0.007796f
C666 B.n552 VSUBS 0.007796f
C667 B.n553 VSUBS 0.007796f
C668 B.n554 VSUBS 0.007796f
C669 B.n555 VSUBS 0.007796f
C670 B.n556 VSUBS 0.007796f
C671 B.n557 VSUBS 0.007796f
C672 B.n558 VSUBS 0.007796f
C673 B.n559 VSUBS 0.007796f
C674 B.n560 VSUBS 0.007796f
C675 B.n561 VSUBS 0.007796f
C676 B.n562 VSUBS 0.007796f
C677 B.n563 VSUBS 0.007796f
C678 B.n564 VSUBS 0.007796f
C679 B.n565 VSUBS 0.007796f
C680 B.n566 VSUBS 0.007796f
C681 B.n567 VSUBS 0.007796f
C682 B.n568 VSUBS 0.007796f
C683 B.n569 VSUBS 0.007796f
C684 B.n570 VSUBS 0.007796f
C685 B.n571 VSUBS 0.007796f
C686 B.n572 VSUBS 0.007796f
C687 B.n573 VSUBS 0.007796f
C688 B.n574 VSUBS 0.007796f
C689 B.n575 VSUBS 0.007796f
C690 B.n576 VSUBS 0.007796f
C691 B.n577 VSUBS 0.007796f
C692 B.n578 VSUBS 0.007796f
C693 B.n579 VSUBS 0.007796f
C694 B.n580 VSUBS 0.007796f
C695 B.n581 VSUBS 0.007796f
C696 B.n582 VSUBS 0.007796f
C697 B.n583 VSUBS 0.007796f
C698 B.n584 VSUBS 0.007796f
C699 B.n585 VSUBS 0.007796f
C700 B.n586 VSUBS 0.007796f
C701 B.n587 VSUBS 0.007796f
C702 B.n588 VSUBS 0.007796f
C703 B.n589 VSUBS 0.007796f
C704 B.n590 VSUBS 0.007796f
C705 B.n591 VSUBS 0.007796f
C706 B.n592 VSUBS 0.007796f
C707 B.n593 VSUBS 0.007796f
C708 B.n594 VSUBS 0.007796f
C709 B.n595 VSUBS 0.007796f
C710 B.n596 VSUBS 0.007796f
C711 B.n597 VSUBS 0.007796f
C712 B.n598 VSUBS 0.007796f
C713 B.n599 VSUBS 0.007796f
C714 B.n600 VSUBS 0.007796f
C715 B.n601 VSUBS 0.007796f
C716 B.n602 VSUBS 0.007796f
C717 B.n603 VSUBS 0.007796f
C718 B.n604 VSUBS 0.007796f
C719 B.n605 VSUBS 0.007796f
C720 B.n606 VSUBS 0.007796f
C721 B.n607 VSUBS 0.007796f
C722 B.n608 VSUBS 0.007796f
C723 B.n609 VSUBS 0.007796f
C724 B.n610 VSUBS 0.007796f
C725 B.n611 VSUBS 0.007796f
C726 B.n612 VSUBS 0.007796f
C727 B.n613 VSUBS 0.007796f
C728 B.n614 VSUBS 0.007796f
C729 B.n615 VSUBS 0.007796f
C730 B.n616 VSUBS 0.007796f
C731 B.n617 VSUBS 0.007796f
C732 B.n618 VSUBS 0.007796f
C733 B.n619 VSUBS 0.007796f
C734 B.n620 VSUBS 0.007796f
C735 B.n621 VSUBS 0.007796f
C736 B.n622 VSUBS 0.007796f
C737 B.n623 VSUBS 0.007796f
C738 B.n624 VSUBS 0.007796f
C739 B.n625 VSUBS 0.007796f
C740 B.n626 VSUBS 0.007796f
C741 B.n627 VSUBS 0.007796f
C742 B.n628 VSUBS 0.007796f
C743 B.n629 VSUBS 0.007796f
C744 B.n630 VSUBS 0.007796f
C745 B.n631 VSUBS 0.007796f
C746 B.n632 VSUBS 0.007796f
C747 B.n633 VSUBS 0.007796f
C748 B.n634 VSUBS 0.007796f
C749 B.n635 VSUBS 0.007796f
C750 B.n636 VSUBS 0.007796f
C751 B.n637 VSUBS 0.007796f
C752 B.n638 VSUBS 0.007796f
C753 B.n639 VSUBS 0.007796f
C754 B.n640 VSUBS 0.007796f
C755 B.n641 VSUBS 0.007796f
C756 B.n642 VSUBS 0.007796f
C757 B.n643 VSUBS 0.007796f
C758 B.n644 VSUBS 0.007796f
C759 B.n645 VSUBS 0.007796f
C760 B.n646 VSUBS 0.017148f
C761 B.n647 VSUBS 0.017936f
C762 B.n648 VSUBS 0.016957f
C763 B.n649 VSUBS 0.007796f
C764 B.n650 VSUBS 0.007796f
C765 B.n651 VSUBS 0.007796f
C766 B.n652 VSUBS 0.007796f
C767 B.n653 VSUBS 0.007796f
C768 B.n654 VSUBS 0.007796f
C769 B.n655 VSUBS 0.007796f
C770 B.n656 VSUBS 0.007796f
C771 B.n657 VSUBS 0.007796f
C772 B.n658 VSUBS 0.007796f
C773 B.n659 VSUBS 0.007796f
C774 B.n660 VSUBS 0.007796f
C775 B.n661 VSUBS 0.007796f
C776 B.n662 VSUBS 0.007796f
C777 B.n663 VSUBS 0.007796f
C778 B.n664 VSUBS 0.007796f
C779 B.n665 VSUBS 0.007796f
C780 B.n666 VSUBS 0.007796f
C781 B.n667 VSUBS 0.007796f
C782 B.n668 VSUBS 0.007796f
C783 B.n669 VSUBS 0.007796f
C784 B.n670 VSUBS 0.007796f
C785 B.n671 VSUBS 0.007796f
C786 B.n672 VSUBS 0.007796f
C787 B.n673 VSUBS 0.007796f
C788 B.n674 VSUBS 0.007796f
C789 B.n675 VSUBS 0.007796f
C790 B.n676 VSUBS 0.007796f
C791 B.n677 VSUBS 0.007796f
C792 B.n678 VSUBS 0.007796f
C793 B.n679 VSUBS 0.007796f
C794 B.n680 VSUBS 0.007796f
C795 B.n681 VSUBS 0.007796f
C796 B.n682 VSUBS 0.007796f
C797 B.n683 VSUBS 0.007796f
C798 B.n684 VSUBS 0.007796f
C799 B.n685 VSUBS 0.007796f
C800 B.n686 VSUBS 0.007796f
C801 B.n687 VSUBS 0.007796f
C802 B.n688 VSUBS 0.007796f
C803 B.n689 VSUBS 0.007796f
C804 B.n690 VSUBS 0.007796f
C805 B.n691 VSUBS 0.007796f
C806 B.n692 VSUBS 0.007796f
C807 B.n693 VSUBS 0.007796f
C808 B.n694 VSUBS 0.007796f
C809 B.n695 VSUBS 0.007796f
C810 B.n696 VSUBS 0.007796f
C811 B.n697 VSUBS 0.007796f
C812 B.n698 VSUBS 0.007796f
C813 B.n699 VSUBS 0.007796f
C814 B.n700 VSUBS 0.007796f
C815 B.n701 VSUBS 0.007796f
C816 B.n702 VSUBS 0.007796f
C817 B.n703 VSUBS 0.007796f
C818 B.n704 VSUBS 0.007796f
C819 B.n705 VSUBS 0.007796f
C820 B.n706 VSUBS 0.007796f
C821 B.n707 VSUBS 0.007796f
C822 B.n708 VSUBS 0.007796f
C823 B.n709 VSUBS 0.007796f
C824 B.n710 VSUBS 0.007796f
C825 B.n711 VSUBS 0.007796f
C826 B.n712 VSUBS 0.007796f
C827 B.n713 VSUBS 0.007796f
C828 B.n714 VSUBS 0.007796f
C829 B.n715 VSUBS 0.007796f
C830 B.n716 VSUBS 0.007796f
C831 B.n717 VSUBS 0.007796f
C832 B.n718 VSUBS 0.007796f
C833 B.n719 VSUBS 0.007796f
C834 B.n720 VSUBS 0.007338f
C835 B.n721 VSUBS 0.018063f
C836 B.n722 VSUBS 0.004357f
C837 B.n723 VSUBS 0.007796f
C838 B.n724 VSUBS 0.007796f
C839 B.n725 VSUBS 0.007796f
C840 B.n726 VSUBS 0.007796f
C841 B.n727 VSUBS 0.007796f
C842 B.n728 VSUBS 0.007796f
C843 B.n729 VSUBS 0.007796f
C844 B.n730 VSUBS 0.007796f
C845 B.n731 VSUBS 0.007796f
C846 B.n732 VSUBS 0.007796f
C847 B.n733 VSUBS 0.007796f
C848 B.n734 VSUBS 0.007796f
C849 B.n735 VSUBS 0.004357f
C850 B.n736 VSUBS 0.007796f
C851 B.n737 VSUBS 0.007796f
C852 B.n738 VSUBS 0.007796f
C853 B.n739 VSUBS 0.007796f
C854 B.n740 VSUBS 0.007796f
C855 B.n741 VSUBS 0.007796f
C856 B.n742 VSUBS 0.007796f
C857 B.n743 VSUBS 0.007796f
C858 B.n744 VSUBS 0.007796f
C859 B.n745 VSUBS 0.007796f
C860 B.n746 VSUBS 0.007796f
C861 B.n747 VSUBS 0.007796f
C862 B.n748 VSUBS 0.007796f
C863 B.n749 VSUBS 0.007796f
C864 B.n750 VSUBS 0.007796f
C865 B.n751 VSUBS 0.007796f
C866 B.n752 VSUBS 0.007796f
C867 B.n753 VSUBS 0.007796f
C868 B.n754 VSUBS 0.007796f
C869 B.n755 VSUBS 0.007796f
C870 B.n756 VSUBS 0.007796f
C871 B.n757 VSUBS 0.007796f
C872 B.n758 VSUBS 0.007796f
C873 B.n759 VSUBS 0.007796f
C874 B.n760 VSUBS 0.007796f
C875 B.n761 VSUBS 0.007796f
C876 B.n762 VSUBS 0.007796f
C877 B.n763 VSUBS 0.007796f
C878 B.n764 VSUBS 0.007796f
C879 B.n765 VSUBS 0.007796f
C880 B.n766 VSUBS 0.007796f
C881 B.n767 VSUBS 0.007796f
C882 B.n768 VSUBS 0.007796f
C883 B.n769 VSUBS 0.007796f
C884 B.n770 VSUBS 0.007796f
C885 B.n771 VSUBS 0.007796f
C886 B.n772 VSUBS 0.007796f
C887 B.n773 VSUBS 0.007796f
C888 B.n774 VSUBS 0.007796f
C889 B.n775 VSUBS 0.007796f
C890 B.n776 VSUBS 0.007796f
C891 B.n777 VSUBS 0.007796f
C892 B.n778 VSUBS 0.007796f
C893 B.n779 VSUBS 0.007796f
C894 B.n780 VSUBS 0.007796f
C895 B.n781 VSUBS 0.007796f
C896 B.n782 VSUBS 0.007796f
C897 B.n783 VSUBS 0.007796f
C898 B.n784 VSUBS 0.007796f
C899 B.n785 VSUBS 0.007796f
C900 B.n786 VSUBS 0.007796f
C901 B.n787 VSUBS 0.007796f
C902 B.n788 VSUBS 0.007796f
C903 B.n789 VSUBS 0.007796f
C904 B.n790 VSUBS 0.007796f
C905 B.n791 VSUBS 0.007796f
C906 B.n792 VSUBS 0.007796f
C907 B.n793 VSUBS 0.007796f
C908 B.n794 VSUBS 0.007796f
C909 B.n795 VSUBS 0.007796f
C910 B.n796 VSUBS 0.007796f
C911 B.n797 VSUBS 0.007796f
C912 B.n798 VSUBS 0.007796f
C913 B.n799 VSUBS 0.007796f
C914 B.n800 VSUBS 0.007796f
C915 B.n801 VSUBS 0.007796f
C916 B.n802 VSUBS 0.007796f
C917 B.n803 VSUBS 0.007796f
C918 B.n804 VSUBS 0.007796f
C919 B.n805 VSUBS 0.007796f
C920 B.n806 VSUBS 0.007796f
C921 B.n807 VSUBS 0.007796f
C922 B.n808 VSUBS 0.007796f
C923 B.n809 VSUBS 0.017936f
C924 B.n810 VSUBS 0.017148f
C925 B.n811 VSUBS 0.017148f
C926 B.n812 VSUBS 0.007796f
C927 B.n813 VSUBS 0.007796f
C928 B.n814 VSUBS 0.007796f
C929 B.n815 VSUBS 0.007796f
C930 B.n816 VSUBS 0.007796f
C931 B.n817 VSUBS 0.007796f
C932 B.n818 VSUBS 0.007796f
C933 B.n819 VSUBS 0.007796f
C934 B.n820 VSUBS 0.007796f
C935 B.n821 VSUBS 0.007796f
C936 B.n822 VSUBS 0.007796f
C937 B.n823 VSUBS 0.007796f
C938 B.n824 VSUBS 0.007796f
C939 B.n825 VSUBS 0.007796f
C940 B.n826 VSUBS 0.007796f
C941 B.n827 VSUBS 0.007796f
C942 B.n828 VSUBS 0.007796f
C943 B.n829 VSUBS 0.007796f
C944 B.n830 VSUBS 0.007796f
C945 B.n831 VSUBS 0.007796f
C946 B.n832 VSUBS 0.007796f
C947 B.n833 VSUBS 0.007796f
C948 B.n834 VSUBS 0.007796f
C949 B.n835 VSUBS 0.007796f
C950 B.n836 VSUBS 0.007796f
C951 B.n837 VSUBS 0.007796f
C952 B.n838 VSUBS 0.007796f
C953 B.n839 VSUBS 0.007796f
C954 B.n840 VSUBS 0.007796f
C955 B.n841 VSUBS 0.007796f
C956 B.n842 VSUBS 0.007796f
C957 B.n843 VSUBS 0.007796f
C958 B.n844 VSUBS 0.007796f
C959 B.n845 VSUBS 0.007796f
C960 B.n846 VSUBS 0.007796f
C961 B.n847 VSUBS 0.007796f
C962 B.n848 VSUBS 0.007796f
C963 B.n849 VSUBS 0.007796f
C964 B.n850 VSUBS 0.007796f
C965 B.n851 VSUBS 0.007796f
C966 B.n852 VSUBS 0.007796f
C967 B.n853 VSUBS 0.007796f
C968 B.n854 VSUBS 0.007796f
C969 B.n855 VSUBS 0.007796f
C970 B.n856 VSUBS 0.007796f
C971 B.n857 VSUBS 0.007796f
C972 B.n858 VSUBS 0.007796f
C973 B.n859 VSUBS 0.007796f
C974 B.n860 VSUBS 0.007796f
C975 B.n861 VSUBS 0.007796f
C976 B.n862 VSUBS 0.007796f
C977 B.n863 VSUBS 0.007796f
C978 B.n864 VSUBS 0.007796f
C979 B.n865 VSUBS 0.007796f
C980 B.n866 VSUBS 0.007796f
C981 B.n867 VSUBS 0.007796f
C982 B.n868 VSUBS 0.007796f
C983 B.n869 VSUBS 0.007796f
C984 B.n870 VSUBS 0.007796f
C985 B.n871 VSUBS 0.007796f
C986 B.n872 VSUBS 0.007796f
C987 B.n873 VSUBS 0.007796f
C988 B.n874 VSUBS 0.007796f
C989 B.n875 VSUBS 0.007796f
C990 B.n876 VSUBS 0.007796f
C991 B.n877 VSUBS 0.007796f
C992 B.n878 VSUBS 0.007796f
C993 B.n879 VSUBS 0.007796f
C994 B.n880 VSUBS 0.007796f
C995 B.n881 VSUBS 0.007796f
C996 B.n882 VSUBS 0.007796f
C997 B.n883 VSUBS 0.007796f
C998 B.n884 VSUBS 0.007796f
C999 B.n885 VSUBS 0.007796f
C1000 B.n886 VSUBS 0.007796f
C1001 B.n887 VSUBS 0.007796f
C1002 B.n888 VSUBS 0.007796f
C1003 B.n889 VSUBS 0.007796f
C1004 B.n890 VSUBS 0.007796f
C1005 B.n891 VSUBS 0.007796f
C1006 B.n892 VSUBS 0.007796f
C1007 B.n893 VSUBS 0.007796f
C1008 B.n894 VSUBS 0.007796f
C1009 B.n895 VSUBS 0.017654f
C1010 VTAIL.t10 VSUBS 0.335545f
C1011 VTAIL.t8 VSUBS 0.335545f
C1012 VTAIL.n0 VSUBS 2.51467f
C1013 VTAIL.n1 VSUBS 1.00873f
C1014 VTAIL.t0 VSUBS 3.30547f
C1015 VTAIL.n2 VSUBS 1.37409f
C1016 VTAIL.t5 VSUBS 0.335545f
C1017 VTAIL.t4 VSUBS 0.335545f
C1018 VTAIL.n3 VSUBS 2.51467f
C1019 VTAIL.n4 VSUBS 3.27402f
C1020 VTAIL.t7 VSUBS 0.335545f
C1021 VTAIL.t11 VSUBS 0.335545f
C1022 VTAIL.n5 VSUBS 2.51467f
C1023 VTAIL.n6 VSUBS 3.27402f
C1024 VTAIL.t9 VSUBS 3.30548f
C1025 VTAIL.n7 VSUBS 1.37407f
C1026 VTAIL.t2 VSUBS 0.335545f
C1027 VTAIL.t3 VSUBS 0.335545f
C1028 VTAIL.n8 VSUBS 2.51467f
C1029 VTAIL.n9 VSUBS 1.24976f
C1030 VTAIL.t1 VSUBS 3.30549f
C1031 VTAIL.n10 VSUBS 3.06965f
C1032 VTAIL.t6 VSUBS 3.30547f
C1033 VTAIL.n11 VSUBS 2.98204f
C1034 VDD2.t3 VSUBS 3.40191f
C1035 VDD2.t4 VSUBS 0.322586f
C1036 VDD2.t0 VSUBS 0.322586f
C1037 VDD2.n0 VSUBS 2.5997f
C1038 VDD2.n1 VSUBS 4.63552f
C1039 VDD2.t1 VSUBS 3.37124f
C1040 VDD2.n2 VSUBS 4.04355f
C1041 VDD2.t2 VSUBS 0.322586f
C1042 VDD2.t5 VSUBS 0.322586f
C1043 VDD2.n3 VSUBS 2.59965f
C1044 VN.t5 VSUBS 3.51293f
C1045 VN.n0 VSUBS 1.30723f
C1046 VN.n1 VSUBS 0.023605f
C1047 VN.n2 VSUBS 0.046078f
C1048 VN.n3 VSUBS 0.023605f
C1049 VN.n4 VSUBS 0.043995f
C1050 VN.t3 VSUBS 3.51293f
C1051 VN.n5 VSUBS 1.31689f
C1052 VN.t1 VSUBS 3.87738f
C1053 VN.n6 VSUBS 1.25011f
C1054 VN.n7 VSUBS 0.301378f
C1055 VN.n8 VSUBS 0.023605f
C1056 VN.n9 VSUBS 0.043995f
C1057 VN.n10 VSUBS 0.047479f
C1058 VN.n11 VSUBS 0.019357f
C1059 VN.n12 VSUBS 0.023605f
C1060 VN.n13 VSUBS 0.023605f
C1061 VN.n14 VSUBS 0.023605f
C1062 VN.n15 VSUBS 0.043995f
C1063 VN.n16 VSUBS 0.043995f
C1064 VN.n17 VSUBS 0.024881f
C1065 VN.n18 VSUBS 0.038099f
C1066 VN.n19 VSUBS 0.071561f
C1067 VN.t4 VSUBS 3.51293f
C1068 VN.n20 VSUBS 1.30723f
C1069 VN.n21 VSUBS 0.023605f
C1070 VN.n22 VSUBS 0.046078f
C1071 VN.n23 VSUBS 0.023605f
C1072 VN.n24 VSUBS 0.043995f
C1073 VN.t2 VSUBS 3.87738f
C1074 VN.t0 VSUBS 3.51293f
C1075 VN.n25 VSUBS 1.31689f
C1076 VN.n26 VSUBS 1.25011f
C1077 VN.n27 VSUBS 0.301378f
C1078 VN.n28 VSUBS 0.023605f
C1079 VN.n29 VSUBS 0.043995f
C1080 VN.n30 VSUBS 0.047479f
C1081 VN.n31 VSUBS 0.019357f
C1082 VN.n32 VSUBS 0.023605f
C1083 VN.n33 VSUBS 0.023605f
C1084 VN.n34 VSUBS 0.023605f
C1085 VN.n35 VSUBS 0.043995f
C1086 VN.n36 VSUBS 0.043995f
C1087 VN.n37 VSUBS 0.024881f
C1088 VN.n38 VSUBS 0.038099f
C1089 VN.n39 VSUBS 1.5627f
.ends

