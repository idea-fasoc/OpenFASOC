* NGSPICE file created from diff_pair_sample_0057.ext - technology: sky130A

.subckt diff_pair_sample_0057 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t11 VN.t0 VDD2.t0 w_n3178_n2648# sky130_fd_pr__pfet_01v8 ad=1.386 pd=8.73 as=1.386 ps=8.73 w=8.4 l=2.43
X1 VDD1.t5 VP.t0 VTAIL.t3 w_n3178_n2648# sky130_fd_pr__pfet_01v8 ad=3.276 pd=17.58 as=1.386 ps=8.73 w=8.4 l=2.43
X2 B.t11 B.t9 B.t10 w_n3178_n2648# sky130_fd_pr__pfet_01v8 ad=3.276 pd=17.58 as=0 ps=0 w=8.4 l=2.43
X3 VTAIL.t5 VP.t1 VDD1.t4 w_n3178_n2648# sky130_fd_pr__pfet_01v8 ad=1.386 pd=8.73 as=1.386 ps=8.73 w=8.4 l=2.43
X4 B.t8 B.t6 B.t7 w_n3178_n2648# sky130_fd_pr__pfet_01v8 ad=3.276 pd=17.58 as=0 ps=0 w=8.4 l=2.43
X5 VDD1.t3 VP.t2 VTAIL.t4 w_n3178_n2648# sky130_fd_pr__pfet_01v8 ad=3.276 pd=17.58 as=1.386 ps=8.73 w=8.4 l=2.43
X6 VDD2.t4 VN.t1 VTAIL.t10 w_n3178_n2648# sky130_fd_pr__pfet_01v8 ad=1.386 pd=8.73 as=3.276 ps=17.58 w=8.4 l=2.43
X7 VDD1.t2 VP.t3 VTAIL.t0 w_n3178_n2648# sky130_fd_pr__pfet_01v8 ad=1.386 pd=8.73 as=3.276 ps=17.58 w=8.4 l=2.43
X8 VDD2.t2 VN.t2 VTAIL.t9 w_n3178_n2648# sky130_fd_pr__pfet_01v8 ad=1.386 pd=8.73 as=3.276 ps=17.58 w=8.4 l=2.43
X9 VTAIL.t8 VN.t3 VDD2.t1 w_n3178_n2648# sky130_fd_pr__pfet_01v8 ad=1.386 pd=8.73 as=1.386 ps=8.73 w=8.4 l=2.43
X10 VDD1.t1 VP.t4 VTAIL.t1 w_n3178_n2648# sky130_fd_pr__pfet_01v8 ad=1.386 pd=8.73 as=3.276 ps=17.58 w=8.4 l=2.43
X11 B.t5 B.t3 B.t4 w_n3178_n2648# sky130_fd_pr__pfet_01v8 ad=3.276 pd=17.58 as=0 ps=0 w=8.4 l=2.43
X12 VTAIL.t2 VP.t5 VDD1.t0 w_n3178_n2648# sky130_fd_pr__pfet_01v8 ad=1.386 pd=8.73 as=1.386 ps=8.73 w=8.4 l=2.43
X13 VDD2.t5 VN.t4 VTAIL.t7 w_n3178_n2648# sky130_fd_pr__pfet_01v8 ad=3.276 pd=17.58 as=1.386 ps=8.73 w=8.4 l=2.43
X14 B.t2 B.t0 B.t1 w_n3178_n2648# sky130_fd_pr__pfet_01v8 ad=3.276 pd=17.58 as=0 ps=0 w=8.4 l=2.43
X15 VDD2.t3 VN.t5 VTAIL.t6 w_n3178_n2648# sky130_fd_pr__pfet_01v8 ad=3.276 pd=17.58 as=1.386 ps=8.73 w=8.4 l=2.43
R0 VN.n25 VN.n14 161.3
R1 VN.n24 VN.n23 161.3
R2 VN.n22 VN.n15 161.3
R3 VN.n21 VN.n20 161.3
R4 VN.n19 VN.n16 161.3
R5 VN.n11 VN.n0 161.3
R6 VN.n10 VN.n9 161.3
R7 VN.n8 VN.n1 161.3
R8 VN.n7 VN.n6 161.3
R9 VN.n5 VN.n2 161.3
R10 VN.n3 VN.t5 117.751
R11 VN.n17 VN.t1 117.751
R12 VN.n13 VN.n12 97.9476
R13 VN.n27 VN.n26 97.9476
R14 VN.n4 VN.t3 83.3091
R15 VN.n12 VN.t2 83.3091
R16 VN.n18 VN.t0 83.3091
R17 VN.n26 VN.t4 83.3091
R18 VN.n6 VN.n1 52.0954
R19 VN.n20 VN.n15 52.0954
R20 VN.n4 VN.n3 47.9149
R21 VN.n18 VN.n17 47.9149
R22 VN VN.n27 45.5815
R23 VN.n10 VN.n1 28.7258
R24 VN.n24 VN.n15 28.7258
R25 VN.n5 VN.n4 24.3439
R26 VN.n6 VN.n5 24.3439
R27 VN.n11 VN.n10 24.3439
R28 VN.n20 VN.n19 24.3439
R29 VN.n19 VN.n18 24.3439
R30 VN.n25 VN.n24 24.3439
R31 VN.n12 VN.n11 12.6591
R32 VN.n26 VN.n25 12.6591
R33 VN.n17 VN.n16 6.67718
R34 VN.n3 VN.n2 6.67718
R35 VN.n27 VN.n14 0.278398
R36 VN.n13 VN.n0 0.278398
R37 VN.n23 VN.n14 0.189894
R38 VN.n23 VN.n22 0.189894
R39 VN.n22 VN.n21 0.189894
R40 VN.n21 VN.n16 0.189894
R41 VN.n7 VN.n2 0.189894
R42 VN.n8 VN.n7 0.189894
R43 VN.n9 VN.n8 0.189894
R44 VN.n9 VN.n0 0.189894
R45 VN VN.n13 0.153422
R46 VDD2.n1 VDD2.t3 84.9705
R47 VDD2.n2 VDD2.t5 83.2416
R48 VDD2.n1 VDD2.n0 79.9114
R49 VDD2 VDD2.n3 79.9086
R50 VDD2.n2 VDD2.n1 38.6894
R51 VDD2.n3 VDD2.t0 3.87014
R52 VDD2.n3 VDD2.t4 3.87014
R53 VDD2.n0 VDD2.t1 3.87014
R54 VDD2.n0 VDD2.t2 3.87014
R55 VDD2 VDD2.n2 1.84317
R56 VTAIL.n7 VTAIL.t10 66.5628
R57 VTAIL.n10 VTAIL.t1 66.5628
R58 VTAIL.n11 VTAIL.t9 66.5626
R59 VTAIL.n2 VTAIL.t0 66.5626
R60 VTAIL.n9 VTAIL.n8 62.6932
R61 VTAIL.n6 VTAIL.n5 62.6932
R62 VTAIL.n1 VTAIL.n0 62.6931
R63 VTAIL.n4 VTAIL.n3 62.6931
R64 VTAIL.n6 VTAIL.n4 24.3669
R65 VTAIL.n11 VTAIL.n10 21.9876
R66 VTAIL.n0 VTAIL.t6 3.87014
R67 VTAIL.n0 VTAIL.t8 3.87014
R68 VTAIL.n3 VTAIL.t3 3.87014
R69 VTAIL.n3 VTAIL.t5 3.87014
R70 VTAIL.n8 VTAIL.t4 3.87014
R71 VTAIL.n8 VTAIL.t2 3.87014
R72 VTAIL.n5 VTAIL.t7 3.87014
R73 VTAIL.n5 VTAIL.t11 3.87014
R74 VTAIL.n7 VTAIL.n6 2.37981
R75 VTAIL.n10 VTAIL.n9 2.37981
R76 VTAIL.n4 VTAIL.n2 2.37981
R77 VTAIL VTAIL.n11 1.72679
R78 VTAIL.n9 VTAIL.n7 1.65998
R79 VTAIL.n2 VTAIL.n1 1.65998
R80 VTAIL VTAIL.n1 0.653517
R81 VP.n11 VP.n8 161.3
R82 VP.n13 VP.n12 161.3
R83 VP.n14 VP.n7 161.3
R84 VP.n16 VP.n15 161.3
R85 VP.n17 VP.n6 161.3
R86 VP.n37 VP.n0 161.3
R87 VP.n36 VP.n35 161.3
R88 VP.n34 VP.n1 161.3
R89 VP.n33 VP.n32 161.3
R90 VP.n31 VP.n2 161.3
R91 VP.n30 VP.n29 161.3
R92 VP.n28 VP.n3 161.3
R93 VP.n27 VP.n26 161.3
R94 VP.n25 VP.n4 161.3
R95 VP.n24 VP.n23 161.3
R96 VP.n22 VP.n5 161.3
R97 VP.n9 VP.t2 117.751
R98 VP.n21 VP.n20 97.9476
R99 VP.n39 VP.n38 97.9476
R100 VP.n19 VP.n18 97.9476
R101 VP.n30 VP.t1 83.3091
R102 VP.n20 VP.t0 83.3091
R103 VP.n38 VP.t3 83.3091
R104 VP.n10 VP.t5 83.3091
R105 VP.n18 VP.t4 83.3091
R106 VP.n26 VP.n25 52.0954
R107 VP.n32 VP.n1 52.0954
R108 VP.n12 VP.n7 52.0954
R109 VP.n10 VP.n9 47.9149
R110 VP.n21 VP.n19 45.3026
R111 VP.n25 VP.n24 28.7258
R112 VP.n36 VP.n1 28.7258
R113 VP.n16 VP.n7 28.7258
R114 VP.n24 VP.n5 24.3439
R115 VP.n26 VP.n3 24.3439
R116 VP.n30 VP.n3 24.3439
R117 VP.n31 VP.n30 24.3439
R118 VP.n32 VP.n31 24.3439
R119 VP.n37 VP.n36 24.3439
R120 VP.n17 VP.n16 24.3439
R121 VP.n11 VP.n10 24.3439
R122 VP.n12 VP.n11 24.3439
R123 VP.n20 VP.n5 12.6591
R124 VP.n38 VP.n37 12.6591
R125 VP.n18 VP.n17 12.6591
R126 VP.n9 VP.n8 6.67718
R127 VP.n19 VP.n6 0.278398
R128 VP.n22 VP.n21 0.278398
R129 VP.n39 VP.n0 0.278398
R130 VP.n13 VP.n8 0.189894
R131 VP.n14 VP.n13 0.189894
R132 VP.n15 VP.n14 0.189894
R133 VP.n15 VP.n6 0.189894
R134 VP.n23 VP.n22 0.189894
R135 VP.n23 VP.n4 0.189894
R136 VP.n27 VP.n4 0.189894
R137 VP.n28 VP.n27 0.189894
R138 VP.n29 VP.n28 0.189894
R139 VP.n29 VP.n2 0.189894
R140 VP.n33 VP.n2 0.189894
R141 VP.n34 VP.n33 0.189894
R142 VP.n35 VP.n34 0.189894
R143 VP.n35 VP.n0 0.189894
R144 VP VP.n39 0.153422
R145 VDD1 VDD1.t3 85.0843
R146 VDD1.n1 VDD1.t5 84.9705
R147 VDD1.n1 VDD1.n0 79.9114
R148 VDD1.n3 VDD1.n2 79.372
R149 VDD1.n3 VDD1.n1 40.4621
R150 VDD1.n2 VDD1.t0 3.87014
R151 VDD1.n2 VDD1.t1 3.87014
R152 VDD1.n0 VDD1.t4 3.87014
R153 VDD1.n0 VDD1.t2 3.87014
R154 VDD1 VDD1.n3 0.537138
R155 B.n331 B.n104 585
R156 B.n330 B.n329 585
R157 B.n328 B.n105 585
R158 B.n327 B.n326 585
R159 B.n325 B.n106 585
R160 B.n324 B.n323 585
R161 B.n322 B.n107 585
R162 B.n321 B.n320 585
R163 B.n319 B.n108 585
R164 B.n318 B.n317 585
R165 B.n316 B.n109 585
R166 B.n315 B.n314 585
R167 B.n313 B.n110 585
R168 B.n312 B.n311 585
R169 B.n310 B.n111 585
R170 B.n309 B.n308 585
R171 B.n307 B.n112 585
R172 B.n306 B.n305 585
R173 B.n304 B.n113 585
R174 B.n303 B.n302 585
R175 B.n301 B.n114 585
R176 B.n300 B.n299 585
R177 B.n298 B.n115 585
R178 B.n297 B.n296 585
R179 B.n295 B.n116 585
R180 B.n294 B.n293 585
R181 B.n292 B.n117 585
R182 B.n291 B.n290 585
R183 B.n289 B.n118 585
R184 B.n288 B.n287 585
R185 B.n286 B.n119 585
R186 B.n285 B.n284 585
R187 B.n280 B.n120 585
R188 B.n279 B.n278 585
R189 B.n277 B.n121 585
R190 B.n276 B.n275 585
R191 B.n274 B.n122 585
R192 B.n273 B.n272 585
R193 B.n271 B.n123 585
R194 B.n270 B.n269 585
R195 B.n268 B.n124 585
R196 B.n266 B.n265 585
R197 B.n264 B.n127 585
R198 B.n263 B.n262 585
R199 B.n261 B.n128 585
R200 B.n260 B.n259 585
R201 B.n258 B.n129 585
R202 B.n257 B.n256 585
R203 B.n255 B.n130 585
R204 B.n254 B.n253 585
R205 B.n252 B.n131 585
R206 B.n251 B.n250 585
R207 B.n249 B.n132 585
R208 B.n248 B.n247 585
R209 B.n246 B.n133 585
R210 B.n245 B.n244 585
R211 B.n243 B.n134 585
R212 B.n242 B.n241 585
R213 B.n240 B.n135 585
R214 B.n239 B.n238 585
R215 B.n237 B.n136 585
R216 B.n236 B.n235 585
R217 B.n234 B.n137 585
R218 B.n233 B.n232 585
R219 B.n231 B.n138 585
R220 B.n230 B.n229 585
R221 B.n228 B.n139 585
R222 B.n227 B.n226 585
R223 B.n225 B.n140 585
R224 B.n224 B.n223 585
R225 B.n222 B.n141 585
R226 B.n221 B.n220 585
R227 B.n333 B.n332 585
R228 B.n334 B.n103 585
R229 B.n336 B.n335 585
R230 B.n337 B.n102 585
R231 B.n339 B.n338 585
R232 B.n340 B.n101 585
R233 B.n342 B.n341 585
R234 B.n343 B.n100 585
R235 B.n345 B.n344 585
R236 B.n346 B.n99 585
R237 B.n348 B.n347 585
R238 B.n349 B.n98 585
R239 B.n351 B.n350 585
R240 B.n352 B.n97 585
R241 B.n354 B.n353 585
R242 B.n355 B.n96 585
R243 B.n357 B.n356 585
R244 B.n358 B.n95 585
R245 B.n360 B.n359 585
R246 B.n361 B.n94 585
R247 B.n363 B.n362 585
R248 B.n364 B.n93 585
R249 B.n366 B.n365 585
R250 B.n367 B.n92 585
R251 B.n369 B.n368 585
R252 B.n370 B.n91 585
R253 B.n372 B.n371 585
R254 B.n373 B.n90 585
R255 B.n375 B.n374 585
R256 B.n376 B.n89 585
R257 B.n378 B.n377 585
R258 B.n379 B.n88 585
R259 B.n381 B.n380 585
R260 B.n382 B.n87 585
R261 B.n384 B.n383 585
R262 B.n385 B.n86 585
R263 B.n387 B.n386 585
R264 B.n388 B.n85 585
R265 B.n390 B.n389 585
R266 B.n391 B.n84 585
R267 B.n393 B.n392 585
R268 B.n394 B.n83 585
R269 B.n396 B.n395 585
R270 B.n397 B.n82 585
R271 B.n399 B.n398 585
R272 B.n400 B.n81 585
R273 B.n402 B.n401 585
R274 B.n403 B.n80 585
R275 B.n405 B.n404 585
R276 B.n406 B.n79 585
R277 B.n408 B.n407 585
R278 B.n409 B.n78 585
R279 B.n411 B.n410 585
R280 B.n412 B.n77 585
R281 B.n414 B.n413 585
R282 B.n415 B.n76 585
R283 B.n417 B.n416 585
R284 B.n418 B.n75 585
R285 B.n420 B.n419 585
R286 B.n421 B.n74 585
R287 B.n423 B.n422 585
R288 B.n424 B.n73 585
R289 B.n426 B.n425 585
R290 B.n427 B.n72 585
R291 B.n429 B.n428 585
R292 B.n430 B.n71 585
R293 B.n432 B.n431 585
R294 B.n433 B.n70 585
R295 B.n435 B.n434 585
R296 B.n436 B.n69 585
R297 B.n438 B.n437 585
R298 B.n439 B.n68 585
R299 B.n441 B.n440 585
R300 B.n442 B.n67 585
R301 B.n444 B.n443 585
R302 B.n445 B.n66 585
R303 B.n447 B.n446 585
R304 B.n448 B.n65 585
R305 B.n450 B.n449 585
R306 B.n451 B.n64 585
R307 B.n453 B.n452 585
R308 B.n454 B.n63 585
R309 B.n563 B.n22 585
R310 B.n562 B.n561 585
R311 B.n560 B.n23 585
R312 B.n559 B.n558 585
R313 B.n557 B.n24 585
R314 B.n556 B.n555 585
R315 B.n554 B.n25 585
R316 B.n553 B.n552 585
R317 B.n551 B.n26 585
R318 B.n550 B.n549 585
R319 B.n548 B.n27 585
R320 B.n547 B.n546 585
R321 B.n545 B.n28 585
R322 B.n544 B.n543 585
R323 B.n542 B.n29 585
R324 B.n541 B.n540 585
R325 B.n539 B.n30 585
R326 B.n538 B.n537 585
R327 B.n536 B.n31 585
R328 B.n535 B.n534 585
R329 B.n533 B.n32 585
R330 B.n532 B.n531 585
R331 B.n530 B.n33 585
R332 B.n529 B.n528 585
R333 B.n527 B.n34 585
R334 B.n526 B.n525 585
R335 B.n524 B.n35 585
R336 B.n523 B.n522 585
R337 B.n521 B.n36 585
R338 B.n520 B.n519 585
R339 B.n518 B.n37 585
R340 B.n516 B.n515 585
R341 B.n514 B.n40 585
R342 B.n513 B.n512 585
R343 B.n511 B.n41 585
R344 B.n510 B.n509 585
R345 B.n508 B.n42 585
R346 B.n507 B.n506 585
R347 B.n505 B.n43 585
R348 B.n504 B.n503 585
R349 B.n502 B.n44 585
R350 B.n501 B.n500 585
R351 B.n499 B.n45 585
R352 B.n498 B.n497 585
R353 B.n496 B.n49 585
R354 B.n495 B.n494 585
R355 B.n493 B.n50 585
R356 B.n492 B.n491 585
R357 B.n490 B.n51 585
R358 B.n489 B.n488 585
R359 B.n487 B.n52 585
R360 B.n486 B.n485 585
R361 B.n484 B.n53 585
R362 B.n483 B.n482 585
R363 B.n481 B.n54 585
R364 B.n480 B.n479 585
R365 B.n478 B.n55 585
R366 B.n477 B.n476 585
R367 B.n475 B.n56 585
R368 B.n474 B.n473 585
R369 B.n472 B.n57 585
R370 B.n471 B.n470 585
R371 B.n469 B.n58 585
R372 B.n468 B.n467 585
R373 B.n466 B.n59 585
R374 B.n465 B.n464 585
R375 B.n463 B.n60 585
R376 B.n462 B.n461 585
R377 B.n460 B.n61 585
R378 B.n459 B.n458 585
R379 B.n457 B.n62 585
R380 B.n456 B.n455 585
R381 B.n565 B.n564 585
R382 B.n566 B.n21 585
R383 B.n568 B.n567 585
R384 B.n569 B.n20 585
R385 B.n571 B.n570 585
R386 B.n572 B.n19 585
R387 B.n574 B.n573 585
R388 B.n575 B.n18 585
R389 B.n577 B.n576 585
R390 B.n578 B.n17 585
R391 B.n580 B.n579 585
R392 B.n581 B.n16 585
R393 B.n583 B.n582 585
R394 B.n584 B.n15 585
R395 B.n586 B.n585 585
R396 B.n587 B.n14 585
R397 B.n589 B.n588 585
R398 B.n590 B.n13 585
R399 B.n592 B.n591 585
R400 B.n593 B.n12 585
R401 B.n595 B.n594 585
R402 B.n596 B.n11 585
R403 B.n598 B.n597 585
R404 B.n599 B.n10 585
R405 B.n601 B.n600 585
R406 B.n602 B.n9 585
R407 B.n604 B.n603 585
R408 B.n605 B.n8 585
R409 B.n607 B.n606 585
R410 B.n608 B.n7 585
R411 B.n610 B.n609 585
R412 B.n611 B.n6 585
R413 B.n613 B.n612 585
R414 B.n614 B.n5 585
R415 B.n616 B.n615 585
R416 B.n617 B.n4 585
R417 B.n619 B.n618 585
R418 B.n620 B.n3 585
R419 B.n622 B.n621 585
R420 B.n623 B.n0 585
R421 B.n2 B.n1 585
R422 B.n162 B.n161 585
R423 B.n164 B.n163 585
R424 B.n165 B.n160 585
R425 B.n167 B.n166 585
R426 B.n168 B.n159 585
R427 B.n170 B.n169 585
R428 B.n171 B.n158 585
R429 B.n173 B.n172 585
R430 B.n174 B.n157 585
R431 B.n176 B.n175 585
R432 B.n177 B.n156 585
R433 B.n179 B.n178 585
R434 B.n180 B.n155 585
R435 B.n182 B.n181 585
R436 B.n183 B.n154 585
R437 B.n185 B.n184 585
R438 B.n186 B.n153 585
R439 B.n188 B.n187 585
R440 B.n189 B.n152 585
R441 B.n191 B.n190 585
R442 B.n192 B.n151 585
R443 B.n194 B.n193 585
R444 B.n195 B.n150 585
R445 B.n197 B.n196 585
R446 B.n198 B.n149 585
R447 B.n200 B.n199 585
R448 B.n201 B.n148 585
R449 B.n203 B.n202 585
R450 B.n204 B.n147 585
R451 B.n206 B.n205 585
R452 B.n207 B.n146 585
R453 B.n209 B.n208 585
R454 B.n210 B.n145 585
R455 B.n212 B.n211 585
R456 B.n213 B.n144 585
R457 B.n215 B.n214 585
R458 B.n216 B.n143 585
R459 B.n218 B.n217 585
R460 B.n219 B.n142 585
R461 B.n221 B.n142 482.89
R462 B.n333 B.n104 482.89
R463 B.n455 B.n454 482.89
R464 B.n564 B.n563 482.89
R465 B.n125 B.t3 291.084
R466 B.n281 B.t6 291.084
R467 B.n46 B.t0 291.084
R468 B.n38 B.t9 291.084
R469 B.n625 B.n624 256.663
R470 B.n624 B.n623 235.042
R471 B.n624 B.n2 235.042
R472 B.n281 B.t7 166.613
R473 B.n46 B.t2 166.613
R474 B.n125 B.t4 166.605
R475 B.n38 B.t11 166.605
R476 B.n222 B.n221 163.367
R477 B.n223 B.n222 163.367
R478 B.n223 B.n140 163.367
R479 B.n227 B.n140 163.367
R480 B.n228 B.n227 163.367
R481 B.n229 B.n228 163.367
R482 B.n229 B.n138 163.367
R483 B.n233 B.n138 163.367
R484 B.n234 B.n233 163.367
R485 B.n235 B.n234 163.367
R486 B.n235 B.n136 163.367
R487 B.n239 B.n136 163.367
R488 B.n240 B.n239 163.367
R489 B.n241 B.n240 163.367
R490 B.n241 B.n134 163.367
R491 B.n245 B.n134 163.367
R492 B.n246 B.n245 163.367
R493 B.n247 B.n246 163.367
R494 B.n247 B.n132 163.367
R495 B.n251 B.n132 163.367
R496 B.n252 B.n251 163.367
R497 B.n253 B.n252 163.367
R498 B.n253 B.n130 163.367
R499 B.n257 B.n130 163.367
R500 B.n258 B.n257 163.367
R501 B.n259 B.n258 163.367
R502 B.n259 B.n128 163.367
R503 B.n263 B.n128 163.367
R504 B.n264 B.n263 163.367
R505 B.n265 B.n264 163.367
R506 B.n265 B.n124 163.367
R507 B.n270 B.n124 163.367
R508 B.n271 B.n270 163.367
R509 B.n272 B.n271 163.367
R510 B.n272 B.n122 163.367
R511 B.n276 B.n122 163.367
R512 B.n277 B.n276 163.367
R513 B.n278 B.n277 163.367
R514 B.n278 B.n120 163.367
R515 B.n285 B.n120 163.367
R516 B.n286 B.n285 163.367
R517 B.n287 B.n286 163.367
R518 B.n287 B.n118 163.367
R519 B.n291 B.n118 163.367
R520 B.n292 B.n291 163.367
R521 B.n293 B.n292 163.367
R522 B.n293 B.n116 163.367
R523 B.n297 B.n116 163.367
R524 B.n298 B.n297 163.367
R525 B.n299 B.n298 163.367
R526 B.n299 B.n114 163.367
R527 B.n303 B.n114 163.367
R528 B.n304 B.n303 163.367
R529 B.n305 B.n304 163.367
R530 B.n305 B.n112 163.367
R531 B.n309 B.n112 163.367
R532 B.n310 B.n309 163.367
R533 B.n311 B.n310 163.367
R534 B.n311 B.n110 163.367
R535 B.n315 B.n110 163.367
R536 B.n316 B.n315 163.367
R537 B.n317 B.n316 163.367
R538 B.n317 B.n108 163.367
R539 B.n321 B.n108 163.367
R540 B.n322 B.n321 163.367
R541 B.n323 B.n322 163.367
R542 B.n323 B.n106 163.367
R543 B.n327 B.n106 163.367
R544 B.n328 B.n327 163.367
R545 B.n329 B.n328 163.367
R546 B.n329 B.n104 163.367
R547 B.n454 B.n453 163.367
R548 B.n453 B.n64 163.367
R549 B.n449 B.n64 163.367
R550 B.n449 B.n448 163.367
R551 B.n448 B.n447 163.367
R552 B.n447 B.n66 163.367
R553 B.n443 B.n66 163.367
R554 B.n443 B.n442 163.367
R555 B.n442 B.n441 163.367
R556 B.n441 B.n68 163.367
R557 B.n437 B.n68 163.367
R558 B.n437 B.n436 163.367
R559 B.n436 B.n435 163.367
R560 B.n435 B.n70 163.367
R561 B.n431 B.n70 163.367
R562 B.n431 B.n430 163.367
R563 B.n430 B.n429 163.367
R564 B.n429 B.n72 163.367
R565 B.n425 B.n72 163.367
R566 B.n425 B.n424 163.367
R567 B.n424 B.n423 163.367
R568 B.n423 B.n74 163.367
R569 B.n419 B.n74 163.367
R570 B.n419 B.n418 163.367
R571 B.n418 B.n417 163.367
R572 B.n417 B.n76 163.367
R573 B.n413 B.n76 163.367
R574 B.n413 B.n412 163.367
R575 B.n412 B.n411 163.367
R576 B.n411 B.n78 163.367
R577 B.n407 B.n78 163.367
R578 B.n407 B.n406 163.367
R579 B.n406 B.n405 163.367
R580 B.n405 B.n80 163.367
R581 B.n401 B.n80 163.367
R582 B.n401 B.n400 163.367
R583 B.n400 B.n399 163.367
R584 B.n399 B.n82 163.367
R585 B.n395 B.n82 163.367
R586 B.n395 B.n394 163.367
R587 B.n394 B.n393 163.367
R588 B.n393 B.n84 163.367
R589 B.n389 B.n84 163.367
R590 B.n389 B.n388 163.367
R591 B.n388 B.n387 163.367
R592 B.n387 B.n86 163.367
R593 B.n383 B.n86 163.367
R594 B.n383 B.n382 163.367
R595 B.n382 B.n381 163.367
R596 B.n381 B.n88 163.367
R597 B.n377 B.n88 163.367
R598 B.n377 B.n376 163.367
R599 B.n376 B.n375 163.367
R600 B.n375 B.n90 163.367
R601 B.n371 B.n90 163.367
R602 B.n371 B.n370 163.367
R603 B.n370 B.n369 163.367
R604 B.n369 B.n92 163.367
R605 B.n365 B.n92 163.367
R606 B.n365 B.n364 163.367
R607 B.n364 B.n363 163.367
R608 B.n363 B.n94 163.367
R609 B.n359 B.n94 163.367
R610 B.n359 B.n358 163.367
R611 B.n358 B.n357 163.367
R612 B.n357 B.n96 163.367
R613 B.n353 B.n96 163.367
R614 B.n353 B.n352 163.367
R615 B.n352 B.n351 163.367
R616 B.n351 B.n98 163.367
R617 B.n347 B.n98 163.367
R618 B.n347 B.n346 163.367
R619 B.n346 B.n345 163.367
R620 B.n345 B.n100 163.367
R621 B.n341 B.n100 163.367
R622 B.n341 B.n340 163.367
R623 B.n340 B.n339 163.367
R624 B.n339 B.n102 163.367
R625 B.n335 B.n102 163.367
R626 B.n335 B.n334 163.367
R627 B.n334 B.n333 163.367
R628 B.n563 B.n562 163.367
R629 B.n562 B.n23 163.367
R630 B.n558 B.n23 163.367
R631 B.n558 B.n557 163.367
R632 B.n557 B.n556 163.367
R633 B.n556 B.n25 163.367
R634 B.n552 B.n25 163.367
R635 B.n552 B.n551 163.367
R636 B.n551 B.n550 163.367
R637 B.n550 B.n27 163.367
R638 B.n546 B.n27 163.367
R639 B.n546 B.n545 163.367
R640 B.n545 B.n544 163.367
R641 B.n544 B.n29 163.367
R642 B.n540 B.n29 163.367
R643 B.n540 B.n539 163.367
R644 B.n539 B.n538 163.367
R645 B.n538 B.n31 163.367
R646 B.n534 B.n31 163.367
R647 B.n534 B.n533 163.367
R648 B.n533 B.n532 163.367
R649 B.n532 B.n33 163.367
R650 B.n528 B.n33 163.367
R651 B.n528 B.n527 163.367
R652 B.n527 B.n526 163.367
R653 B.n526 B.n35 163.367
R654 B.n522 B.n35 163.367
R655 B.n522 B.n521 163.367
R656 B.n521 B.n520 163.367
R657 B.n520 B.n37 163.367
R658 B.n515 B.n37 163.367
R659 B.n515 B.n514 163.367
R660 B.n514 B.n513 163.367
R661 B.n513 B.n41 163.367
R662 B.n509 B.n41 163.367
R663 B.n509 B.n508 163.367
R664 B.n508 B.n507 163.367
R665 B.n507 B.n43 163.367
R666 B.n503 B.n43 163.367
R667 B.n503 B.n502 163.367
R668 B.n502 B.n501 163.367
R669 B.n501 B.n45 163.367
R670 B.n497 B.n45 163.367
R671 B.n497 B.n496 163.367
R672 B.n496 B.n495 163.367
R673 B.n495 B.n50 163.367
R674 B.n491 B.n50 163.367
R675 B.n491 B.n490 163.367
R676 B.n490 B.n489 163.367
R677 B.n489 B.n52 163.367
R678 B.n485 B.n52 163.367
R679 B.n485 B.n484 163.367
R680 B.n484 B.n483 163.367
R681 B.n483 B.n54 163.367
R682 B.n479 B.n54 163.367
R683 B.n479 B.n478 163.367
R684 B.n478 B.n477 163.367
R685 B.n477 B.n56 163.367
R686 B.n473 B.n56 163.367
R687 B.n473 B.n472 163.367
R688 B.n472 B.n471 163.367
R689 B.n471 B.n58 163.367
R690 B.n467 B.n58 163.367
R691 B.n467 B.n466 163.367
R692 B.n466 B.n465 163.367
R693 B.n465 B.n60 163.367
R694 B.n461 B.n60 163.367
R695 B.n461 B.n460 163.367
R696 B.n460 B.n459 163.367
R697 B.n459 B.n62 163.367
R698 B.n455 B.n62 163.367
R699 B.n564 B.n21 163.367
R700 B.n568 B.n21 163.367
R701 B.n569 B.n568 163.367
R702 B.n570 B.n569 163.367
R703 B.n570 B.n19 163.367
R704 B.n574 B.n19 163.367
R705 B.n575 B.n574 163.367
R706 B.n576 B.n575 163.367
R707 B.n576 B.n17 163.367
R708 B.n580 B.n17 163.367
R709 B.n581 B.n580 163.367
R710 B.n582 B.n581 163.367
R711 B.n582 B.n15 163.367
R712 B.n586 B.n15 163.367
R713 B.n587 B.n586 163.367
R714 B.n588 B.n587 163.367
R715 B.n588 B.n13 163.367
R716 B.n592 B.n13 163.367
R717 B.n593 B.n592 163.367
R718 B.n594 B.n593 163.367
R719 B.n594 B.n11 163.367
R720 B.n598 B.n11 163.367
R721 B.n599 B.n598 163.367
R722 B.n600 B.n599 163.367
R723 B.n600 B.n9 163.367
R724 B.n604 B.n9 163.367
R725 B.n605 B.n604 163.367
R726 B.n606 B.n605 163.367
R727 B.n606 B.n7 163.367
R728 B.n610 B.n7 163.367
R729 B.n611 B.n610 163.367
R730 B.n612 B.n611 163.367
R731 B.n612 B.n5 163.367
R732 B.n616 B.n5 163.367
R733 B.n617 B.n616 163.367
R734 B.n618 B.n617 163.367
R735 B.n618 B.n3 163.367
R736 B.n622 B.n3 163.367
R737 B.n623 B.n622 163.367
R738 B.n162 B.n2 163.367
R739 B.n163 B.n162 163.367
R740 B.n163 B.n160 163.367
R741 B.n167 B.n160 163.367
R742 B.n168 B.n167 163.367
R743 B.n169 B.n168 163.367
R744 B.n169 B.n158 163.367
R745 B.n173 B.n158 163.367
R746 B.n174 B.n173 163.367
R747 B.n175 B.n174 163.367
R748 B.n175 B.n156 163.367
R749 B.n179 B.n156 163.367
R750 B.n180 B.n179 163.367
R751 B.n181 B.n180 163.367
R752 B.n181 B.n154 163.367
R753 B.n185 B.n154 163.367
R754 B.n186 B.n185 163.367
R755 B.n187 B.n186 163.367
R756 B.n187 B.n152 163.367
R757 B.n191 B.n152 163.367
R758 B.n192 B.n191 163.367
R759 B.n193 B.n192 163.367
R760 B.n193 B.n150 163.367
R761 B.n197 B.n150 163.367
R762 B.n198 B.n197 163.367
R763 B.n199 B.n198 163.367
R764 B.n199 B.n148 163.367
R765 B.n203 B.n148 163.367
R766 B.n204 B.n203 163.367
R767 B.n205 B.n204 163.367
R768 B.n205 B.n146 163.367
R769 B.n209 B.n146 163.367
R770 B.n210 B.n209 163.367
R771 B.n211 B.n210 163.367
R772 B.n211 B.n144 163.367
R773 B.n215 B.n144 163.367
R774 B.n216 B.n215 163.367
R775 B.n217 B.n216 163.367
R776 B.n217 B.n142 163.367
R777 B.n282 B.t8 113.085
R778 B.n47 B.t1 113.085
R779 B.n126 B.t5 113.076
R780 B.n39 B.t10 113.076
R781 B.n267 B.n126 59.5399
R782 B.n283 B.n282 59.5399
R783 B.n48 B.n47 59.5399
R784 B.n517 B.n39 59.5399
R785 B.n126 B.n125 53.5278
R786 B.n282 B.n281 53.5278
R787 B.n47 B.n46 53.5278
R788 B.n39 B.n38 53.5278
R789 B.n565 B.n22 31.3761
R790 B.n456 B.n63 31.3761
R791 B.n332 B.n331 31.3761
R792 B.n220 B.n219 31.3761
R793 B B.n625 18.0485
R794 B.n566 B.n565 10.6151
R795 B.n567 B.n566 10.6151
R796 B.n567 B.n20 10.6151
R797 B.n571 B.n20 10.6151
R798 B.n572 B.n571 10.6151
R799 B.n573 B.n572 10.6151
R800 B.n573 B.n18 10.6151
R801 B.n577 B.n18 10.6151
R802 B.n578 B.n577 10.6151
R803 B.n579 B.n578 10.6151
R804 B.n579 B.n16 10.6151
R805 B.n583 B.n16 10.6151
R806 B.n584 B.n583 10.6151
R807 B.n585 B.n584 10.6151
R808 B.n585 B.n14 10.6151
R809 B.n589 B.n14 10.6151
R810 B.n590 B.n589 10.6151
R811 B.n591 B.n590 10.6151
R812 B.n591 B.n12 10.6151
R813 B.n595 B.n12 10.6151
R814 B.n596 B.n595 10.6151
R815 B.n597 B.n596 10.6151
R816 B.n597 B.n10 10.6151
R817 B.n601 B.n10 10.6151
R818 B.n602 B.n601 10.6151
R819 B.n603 B.n602 10.6151
R820 B.n603 B.n8 10.6151
R821 B.n607 B.n8 10.6151
R822 B.n608 B.n607 10.6151
R823 B.n609 B.n608 10.6151
R824 B.n609 B.n6 10.6151
R825 B.n613 B.n6 10.6151
R826 B.n614 B.n613 10.6151
R827 B.n615 B.n614 10.6151
R828 B.n615 B.n4 10.6151
R829 B.n619 B.n4 10.6151
R830 B.n620 B.n619 10.6151
R831 B.n621 B.n620 10.6151
R832 B.n621 B.n0 10.6151
R833 B.n561 B.n22 10.6151
R834 B.n561 B.n560 10.6151
R835 B.n560 B.n559 10.6151
R836 B.n559 B.n24 10.6151
R837 B.n555 B.n24 10.6151
R838 B.n555 B.n554 10.6151
R839 B.n554 B.n553 10.6151
R840 B.n553 B.n26 10.6151
R841 B.n549 B.n26 10.6151
R842 B.n549 B.n548 10.6151
R843 B.n548 B.n547 10.6151
R844 B.n547 B.n28 10.6151
R845 B.n543 B.n28 10.6151
R846 B.n543 B.n542 10.6151
R847 B.n542 B.n541 10.6151
R848 B.n541 B.n30 10.6151
R849 B.n537 B.n30 10.6151
R850 B.n537 B.n536 10.6151
R851 B.n536 B.n535 10.6151
R852 B.n535 B.n32 10.6151
R853 B.n531 B.n32 10.6151
R854 B.n531 B.n530 10.6151
R855 B.n530 B.n529 10.6151
R856 B.n529 B.n34 10.6151
R857 B.n525 B.n34 10.6151
R858 B.n525 B.n524 10.6151
R859 B.n524 B.n523 10.6151
R860 B.n523 B.n36 10.6151
R861 B.n519 B.n36 10.6151
R862 B.n519 B.n518 10.6151
R863 B.n516 B.n40 10.6151
R864 B.n512 B.n40 10.6151
R865 B.n512 B.n511 10.6151
R866 B.n511 B.n510 10.6151
R867 B.n510 B.n42 10.6151
R868 B.n506 B.n42 10.6151
R869 B.n506 B.n505 10.6151
R870 B.n505 B.n504 10.6151
R871 B.n504 B.n44 10.6151
R872 B.n500 B.n499 10.6151
R873 B.n499 B.n498 10.6151
R874 B.n498 B.n49 10.6151
R875 B.n494 B.n49 10.6151
R876 B.n494 B.n493 10.6151
R877 B.n493 B.n492 10.6151
R878 B.n492 B.n51 10.6151
R879 B.n488 B.n51 10.6151
R880 B.n488 B.n487 10.6151
R881 B.n487 B.n486 10.6151
R882 B.n486 B.n53 10.6151
R883 B.n482 B.n53 10.6151
R884 B.n482 B.n481 10.6151
R885 B.n481 B.n480 10.6151
R886 B.n480 B.n55 10.6151
R887 B.n476 B.n55 10.6151
R888 B.n476 B.n475 10.6151
R889 B.n475 B.n474 10.6151
R890 B.n474 B.n57 10.6151
R891 B.n470 B.n57 10.6151
R892 B.n470 B.n469 10.6151
R893 B.n469 B.n468 10.6151
R894 B.n468 B.n59 10.6151
R895 B.n464 B.n59 10.6151
R896 B.n464 B.n463 10.6151
R897 B.n463 B.n462 10.6151
R898 B.n462 B.n61 10.6151
R899 B.n458 B.n61 10.6151
R900 B.n458 B.n457 10.6151
R901 B.n457 B.n456 10.6151
R902 B.n452 B.n63 10.6151
R903 B.n452 B.n451 10.6151
R904 B.n451 B.n450 10.6151
R905 B.n450 B.n65 10.6151
R906 B.n446 B.n65 10.6151
R907 B.n446 B.n445 10.6151
R908 B.n445 B.n444 10.6151
R909 B.n444 B.n67 10.6151
R910 B.n440 B.n67 10.6151
R911 B.n440 B.n439 10.6151
R912 B.n439 B.n438 10.6151
R913 B.n438 B.n69 10.6151
R914 B.n434 B.n69 10.6151
R915 B.n434 B.n433 10.6151
R916 B.n433 B.n432 10.6151
R917 B.n432 B.n71 10.6151
R918 B.n428 B.n71 10.6151
R919 B.n428 B.n427 10.6151
R920 B.n427 B.n426 10.6151
R921 B.n426 B.n73 10.6151
R922 B.n422 B.n73 10.6151
R923 B.n422 B.n421 10.6151
R924 B.n421 B.n420 10.6151
R925 B.n420 B.n75 10.6151
R926 B.n416 B.n75 10.6151
R927 B.n416 B.n415 10.6151
R928 B.n415 B.n414 10.6151
R929 B.n414 B.n77 10.6151
R930 B.n410 B.n77 10.6151
R931 B.n410 B.n409 10.6151
R932 B.n409 B.n408 10.6151
R933 B.n408 B.n79 10.6151
R934 B.n404 B.n79 10.6151
R935 B.n404 B.n403 10.6151
R936 B.n403 B.n402 10.6151
R937 B.n402 B.n81 10.6151
R938 B.n398 B.n81 10.6151
R939 B.n398 B.n397 10.6151
R940 B.n397 B.n396 10.6151
R941 B.n396 B.n83 10.6151
R942 B.n392 B.n83 10.6151
R943 B.n392 B.n391 10.6151
R944 B.n391 B.n390 10.6151
R945 B.n390 B.n85 10.6151
R946 B.n386 B.n85 10.6151
R947 B.n386 B.n385 10.6151
R948 B.n385 B.n384 10.6151
R949 B.n384 B.n87 10.6151
R950 B.n380 B.n87 10.6151
R951 B.n380 B.n379 10.6151
R952 B.n379 B.n378 10.6151
R953 B.n378 B.n89 10.6151
R954 B.n374 B.n89 10.6151
R955 B.n374 B.n373 10.6151
R956 B.n373 B.n372 10.6151
R957 B.n372 B.n91 10.6151
R958 B.n368 B.n91 10.6151
R959 B.n368 B.n367 10.6151
R960 B.n367 B.n366 10.6151
R961 B.n366 B.n93 10.6151
R962 B.n362 B.n93 10.6151
R963 B.n362 B.n361 10.6151
R964 B.n361 B.n360 10.6151
R965 B.n360 B.n95 10.6151
R966 B.n356 B.n95 10.6151
R967 B.n356 B.n355 10.6151
R968 B.n355 B.n354 10.6151
R969 B.n354 B.n97 10.6151
R970 B.n350 B.n97 10.6151
R971 B.n350 B.n349 10.6151
R972 B.n349 B.n348 10.6151
R973 B.n348 B.n99 10.6151
R974 B.n344 B.n99 10.6151
R975 B.n344 B.n343 10.6151
R976 B.n343 B.n342 10.6151
R977 B.n342 B.n101 10.6151
R978 B.n338 B.n101 10.6151
R979 B.n338 B.n337 10.6151
R980 B.n337 B.n336 10.6151
R981 B.n336 B.n103 10.6151
R982 B.n332 B.n103 10.6151
R983 B.n161 B.n1 10.6151
R984 B.n164 B.n161 10.6151
R985 B.n165 B.n164 10.6151
R986 B.n166 B.n165 10.6151
R987 B.n166 B.n159 10.6151
R988 B.n170 B.n159 10.6151
R989 B.n171 B.n170 10.6151
R990 B.n172 B.n171 10.6151
R991 B.n172 B.n157 10.6151
R992 B.n176 B.n157 10.6151
R993 B.n177 B.n176 10.6151
R994 B.n178 B.n177 10.6151
R995 B.n178 B.n155 10.6151
R996 B.n182 B.n155 10.6151
R997 B.n183 B.n182 10.6151
R998 B.n184 B.n183 10.6151
R999 B.n184 B.n153 10.6151
R1000 B.n188 B.n153 10.6151
R1001 B.n189 B.n188 10.6151
R1002 B.n190 B.n189 10.6151
R1003 B.n190 B.n151 10.6151
R1004 B.n194 B.n151 10.6151
R1005 B.n195 B.n194 10.6151
R1006 B.n196 B.n195 10.6151
R1007 B.n196 B.n149 10.6151
R1008 B.n200 B.n149 10.6151
R1009 B.n201 B.n200 10.6151
R1010 B.n202 B.n201 10.6151
R1011 B.n202 B.n147 10.6151
R1012 B.n206 B.n147 10.6151
R1013 B.n207 B.n206 10.6151
R1014 B.n208 B.n207 10.6151
R1015 B.n208 B.n145 10.6151
R1016 B.n212 B.n145 10.6151
R1017 B.n213 B.n212 10.6151
R1018 B.n214 B.n213 10.6151
R1019 B.n214 B.n143 10.6151
R1020 B.n218 B.n143 10.6151
R1021 B.n219 B.n218 10.6151
R1022 B.n220 B.n141 10.6151
R1023 B.n224 B.n141 10.6151
R1024 B.n225 B.n224 10.6151
R1025 B.n226 B.n225 10.6151
R1026 B.n226 B.n139 10.6151
R1027 B.n230 B.n139 10.6151
R1028 B.n231 B.n230 10.6151
R1029 B.n232 B.n231 10.6151
R1030 B.n232 B.n137 10.6151
R1031 B.n236 B.n137 10.6151
R1032 B.n237 B.n236 10.6151
R1033 B.n238 B.n237 10.6151
R1034 B.n238 B.n135 10.6151
R1035 B.n242 B.n135 10.6151
R1036 B.n243 B.n242 10.6151
R1037 B.n244 B.n243 10.6151
R1038 B.n244 B.n133 10.6151
R1039 B.n248 B.n133 10.6151
R1040 B.n249 B.n248 10.6151
R1041 B.n250 B.n249 10.6151
R1042 B.n250 B.n131 10.6151
R1043 B.n254 B.n131 10.6151
R1044 B.n255 B.n254 10.6151
R1045 B.n256 B.n255 10.6151
R1046 B.n256 B.n129 10.6151
R1047 B.n260 B.n129 10.6151
R1048 B.n261 B.n260 10.6151
R1049 B.n262 B.n261 10.6151
R1050 B.n262 B.n127 10.6151
R1051 B.n266 B.n127 10.6151
R1052 B.n269 B.n268 10.6151
R1053 B.n269 B.n123 10.6151
R1054 B.n273 B.n123 10.6151
R1055 B.n274 B.n273 10.6151
R1056 B.n275 B.n274 10.6151
R1057 B.n275 B.n121 10.6151
R1058 B.n279 B.n121 10.6151
R1059 B.n280 B.n279 10.6151
R1060 B.n284 B.n280 10.6151
R1061 B.n288 B.n119 10.6151
R1062 B.n289 B.n288 10.6151
R1063 B.n290 B.n289 10.6151
R1064 B.n290 B.n117 10.6151
R1065 B.n294 B.n117 10.6151
R1066 B.n295 B.n294 10.6151
R1067 B.n296 B.n295 10.6151
R1068 B.n296 B.n115 10.6151
R1069 B.n300 B.n115 10.6151
R1070 B.n301 B.n300 10.6151
R1071 B.n302 B.n301 10.6151
R1072 B.n302 B.n113 10.6151
R1073 B.n306 B.n113 10.6151
R1074 B.n307 B.n306 10.6151
R1075 B.n308 B.n307 10.6151
R1076 B.n308 B.n111 10.6151
R1077 B.n312 B.n111 10.6151
R1078 B.n313 B.n312 10.6151
R1079 B.n314 B.n313 10.6151
R1080 B.n314 B.n109 10.6151
R1081 B.n318 B.n109 10.6151
R1082 B.n319 B.n318 10.6151
R1083 B.n320 B.n319 10.6151
R1084 B.n320 B.n107 10.6151
R1085 B.n324 B.n107 10.6151
R1086 B.n325 B.n324 10.6151
R1087 B.n326 B.n325 10.6151
R1088 B.n326 B.n105 10.6151
R1089 B.n330 B.n105 10.6151
R1090 B.n331 B.n330 10.6151
R1091 B.n518 B.n517 9.36635
R1092 B.n500 B.n48 9.36635
R1093 B.n267 B.n266 9.36635
R1094 B.n283 B.n119 9.36635
R1095 B.n625 B.n0 8.11757
R1096 B.n625 B.n1 8.11757
R1097 B.n517 B.n516 1.24928
R1098 B.n48 B.n44 1.24928
R1099 B.n268 B.n267 1.24928
R1100 B.n284 B.n283 1.24928
C0 VDD2 w_n3178_n2648# 2.07915f
C1 VP VDD1 5.04788f
C2 VDD2 B 1.83568f
C3 w_n3178_n2648# VN 5.91768f
C4 VTAIL VP 5.04685f
C5 B VN 1.08535f
C6 VDD2 VDD1 1.34028f
C7 VDD2 VTAIL 6.41817f
C8 VDD1 VN 0.150164f
C9 VTAIL VN 5.03261f
C10 w_n3178_n2648# B 8.4319f
C11 VDD2 VP 0.44327f
C12 VP VN 6.099299f
C13 w_n3178_n2648# VDD1 1.99949f
C14 w_n3178_n2648# VTAIL 2.45681f
C15 B VDD1 1.76566f
C16 B VTAIL 2.82698f
C17 VDD2 VN 4.75735f
C18 w_n3178_n2648# VP 6.32808f
C19 B VP 1.7697f
C20 VTAIL VDD1 6.36777f
C21 VDD2 VSUBS 1.662967f
C22 VDD1 VSUBS 1.987368f
C23 VTAIL VSUBS 1.03059f
C24 VN VSUBS 5.55328f
C25 VP VSUBS 2.672791f
C26 B VSUBS 4.161675f
C27 w_n3178_n2648# VSUBS 0.104302p
C28 B.n0 VSUBS 0.006096f
C29 B.n1 VSUBS 0.006096f
C30 B.n2 VSUBS 0.009015f
C31 B.n3 VSUBS 0.006909f
C32 B.n4 VSUBS 0.006909f
C33 B.n5 VSUBS 0.006909f
C34 B.n6 VSUBS 0.006909f
C35 B.n7 VSUBS 0.006909f
C36 B.n8 VSUBS 0.006909f
C37 B.n9 VSUBS 0.006909f
C38 B.n10 VSUBS 0.006909f
C39 B.n11 VSUBS 0.006909f
C40 B.n12 VSUBS 0.006909f
C41 B.n13 VSUBS 0.006909f
C42 B.n14 VSUBS 0.006909f
C43 B.n15 VSUBS 0.006909f
C44 B.n16 VSUBS 0.006909f
C45 B.n17 VSUBS 0.006909f
C46 B.n18 VSUBS 0.006909f
C47 B.n19 VSUBS 0.006909f
C48 B.n20 VSUBS 0.006909f
C49 B.n21 VSUBS 0.006909f
C50 B.n22 VSUBS 0.016338f
C51 B.n23 VSUBS 0.006909f
C52 B.n24 VSUBS 0.006909f
C53 B.n25 VSUBS 0.006909f
C54 B.n26 VSUBS 0.006909f
C55 B.n27 VSUBS 0.006909f
C56 B.n28 VSUBS 0.006909f
C57 B.n29 VSUBS 0.006909f
C58 B.n30 VSUBS 0.006909f
C59 B.n31 VSUBS 0.006909f
C60 B.n32 VSUBS 0.006909f
C61 B.n33 VSUBS 0.006909f
C62 B.n34 VSUBS 0.006909f
C63 B.n35 VSUBS 0.006909f
C64 B.n36 VSUBS 0.006909f
C65 B.n37 VSUBS 0.006909f
C66 B.t10 VSUBS 0.25781f
C67 B.t11 VSUBS 0.277087f
C68 B.t9 VSUBS 0.933044f
C69 B.n38 VSUBS 0.147264f
C70 B.n39 VSUBS 0.069854f
C71 B.n40 VSUBS 0.006909f
C72 B.n41 VSUBS 0.006909f
C73 B.n42 VSUBS 0.006909f
C74 B.n43 VSUBS 0.006909f
C75 B.n44 VSUBS 0.003861f
C76 B.n45 VSUBS 0.006909f
C77 B.t1 VSUBS 0.257808f
C78 B.t2 VSUBS 0.277085f
C79 B.t0 VSUBS 0.933044f
C80 B.n46 VSUBS 0.147267f
C81 B.n47 VSUBS 0.069857f
C82 B.n48 VSUBS 0.016007f
C83 B.n49 VSUBS 0.006909f
C84 B.n50 VSUBS 0.006909f
C85 B.n51 VSUBS 0.006909f
C86 B.n52 VSUBS 0.006909f
C87 B.n53 VSUBS 0.006909f
C88 B.n54 VSUBS 0.006909f
C89 B.n55 VSUBS 0.006909f
C90 B.n56 VSUBS 0.006909f
C91 B.n57 VSUBS 0.006909f
C92 B.n58 VSUBS 0.006909f
C93 B.n59 VSUBS 0.006909f
C94 B.n60 VSUBS 0.006909f
C95 B.n61 VSUBS 0.006909f
C96 B.n62 VSUBS 0.006909f
C97 B.n63 VSUBS 0.015157f
C98 B.n64 VSUBS 0.006909f
C99 B.n65 VSUBS 0.006909f
C100 B.n66 VSUBS 0.006909f
C101 B.n67 VSUBS 0.006909f
C102 B.n68 VSUBS 0.006909f
C103 B.n69 VSUBS 0.006909f
C104 B.n70 VSUBS 0.006909f
C105 B.n71 VSUBS 0.006909f
C106 B.n72 VSUBS 0.006909f
C107 B.n73 VSUBS 0.006909f
C108 B.n74 VSUBS 0.006909f
C109 B.n75 VSUBS 0.006909f
C110 B.n76 VSUBS 0.006909f
C111 B.n77 VSUBS 0.006909f
C112 B.n78 VSUBS 0.006909f
C113 B.n79 VSUBS 0.006909f
C114 B.n80 VSUBS 0.006909f
C115 B.n81 VSUBS 0.006909f
C116 B.n82 VSUBS 0.006909f
C117 B.n83 VSUBS 0.006909f
C118 B.n84 VSUBS 0.006909f
C119 B.n85 VSUBS 0.006909f
C120 B.n86 VSUBS 0.006909f
C121 B.n87 VSUBS 0.006909f
C122 B.n88 VSUBS 0.006909f
C123 B.n89 VSUBS 0.006909f
C124 B.n90 VSUBS 0.006909f
C125 B.n91 VSUBS 0.006909f
C126 B.n92 VSUBS 0.006909f
C127 B.n93 VSUBS 0.006909f
C128 B.n94 VSUBS 0.006909f
C129 B.n95 VSUBS 0.006909f
C130 B.n96 VSUBS 0.006909f
C131 B.n97 VSUBS 0.006909f
C132 B.n98 VSUBS 0.006909f
C133 B.n99 VSUBS 0.006909f
C134 B.n100 VSUBS 0.006909f
C135 B.n101 VSUBS 0.006909f
C136 B.n102 VSUBS 0.006909f
C137 B.n103 VSUBS 0.006909f
C138 B.n104 VSUBS 0.016338f
C139 B.n105 VSUBS 0.006909f
C140 B.n106 VSUBS 0.006909f
C141 B.n107 VSUBS 0.006909f
C142 B.n108 VSUBS 0.006909f
C143 B.n109 VSUBS 0.006909f
C144 B.n110 VSUBS 0.006909f
C145 B.n111 VSUBS 0.006909f
C146 B.n112 VSUBS 0.006909f
C147 B.n113 VSUBS 0.006909f
C148 B.n114 VSUBS 0.006909f
C149 B.n115 VSUBS 0.006909f
C150 B.n116 VSUBS 0.006909f
C151 B.n117 VSUBS 0.006909f
C152 B.n118 VSUBS 0.006909f
C153 B.n119 VSUBS 0.006502f
C154 B.n120 VSUBS 0.006909f
C155 B.n121 VSUBS 0.006909f
C156 B.n122 VSUBS 0.006909f
C157 B.n123 VSUBS 0.006909f
C158 B.n124 VSUBS 0.006909f
C159 B.t5 VSUBS 0.25781f
C160 B.t4 VSUBS 0.277087f
C161 B.t3 VSUBS 0.933044f
C162 B.n125 VSUBS 0.147264f
C163 B.n126 VSUBS 0.069854f
C164 B.n127 VSUBS 0.006909f
C165 B.n128 VSUBS 0.006909f
C166 B.n129 VSUBS 0.006909f
C167 B.n130 VSUBS 0.006909f
C168 B.n131 VSUBS 0.006909f
C169 B.n132 VSUBS 0.006909f
C170 B.n133 VSUBS 0.006909f
C171 B.n134 VSUBS 0.006909f
C172 B.n135 VSUBS 0.006909f
C173 B.n136 VSUBS 0.006909f
C174 B.n137 VSUBS 0.006909f
C175 B.n138 VSUBS 0.006909f
C176 B.n139 VSUBS 0.006909f
C177 B.n140 VSUBS 0.006909f
C178 B.n141 VSUBS 0.006909f
C179 B.n142 VSUBS 0.015157f
C180 B.n143 VSUBS 0.006909f
C181 B.n144 VSUBS 0.006909f
C182 B.n145 VSUBS 0.006909f
C183 B.n146 VSUBS 0.006909f
C184 B.n147 VSUBS 0.006909f
C185 B.n148 VSUBS 0.006909f
C186 B.n149 VSUBS 0.006909f
C187 B.n150 VSUBS 0.006909f
C188 B.n151 VSUBS 0.006909f
C189 B.n152 VSUBS 0.006909f
C190 B.n153 VSUBS 0.006909f
C191 B.n154 VSUBS 0.006909f
C192 B.n155 VSUBS 0.006909f
C193 B.n156 VSUBS 0.006909f
C194 B.n157 VSUBS 0.006909f
C195 B.n158 VSUBS 0.006909f
C196 B.n159 VSUBS 0.006909f
C197 B.n160 VSUBS 0.006909f
C198 B.n161 VSUBS 0.006909f
C199 B.n162 VSUBS 0.006909f
C200 B.n163 VSUBS 0.006909f
C201 B.n164 VSUBS 0.006909f
C202 B.n165 VSUBS 0.006909f
C203 B.n166 VSUBS 0.006909f
C204 B.n167 VSUBS 0.006909f
C205 B.n168 VSUBS 0.006909f
C206 B.n169 VSUBS 0.006909f
C207 B.n170 VSUBS 0.006909f
C208 B.n171 VSUBS 0.006909f
C209 B.n172 VSUBS 0.006909f
C210 B.n173 VSUBS 0.006909f
C211 B.n174 VSUBS 0.006909f
C212 B.n175 VSUBS 0.006909f
C213 B.n176 VSUBS 0.006909f
C214 B.n177 VSUBS 0.006909f
C215 B.n178 VSUBS 0.006909f
C216 B.n179 VSUBS 0.006909f
C217 B.n180 VSUBS 0.006909f
C218 B.n181 VSUBS 0.006909f
C219 B.n182 VSUBS 0.006909f
C220 B.n183 VSUBS 0.006909f
C221 B.n184 VSUBS 0.006909f
C222 B.n185 VSUBS 0.006909f
C223 B.n186 VSUBS 0.006909f
C224 B.n187 VSUBS 0.006909f
C225 B.n188 VSUBS 0.006909f
C226 B.n189 VSUBS 0.006909f
C227 B.n190 VSUBS 0.006909f
C228 B.n191 VSUBS 0.006909f
C229 B.n192 VSUBS 0.006909f
C230 B.n193 VSUBS 0.006909f
C231 B.n194 VSUBS 0.006909f
C232 B.n195 VSUBS 0.006909f
C233 B.n196 VSUBS 0.006909f
C234 B.n197 VSUBS 0.006909f
C235 B.n198 VSUBS 0.006909f
C236 B.n199 VSUBS 0.006909f
C237 B.n200 VSUBS 0.006909f
C238 B.n201 VSUBS 0.006909f
C239 B.n202 VSUBS 0.006909f
C240 B.n203 VSUBS 0.006909f
C241 B.n204 VSUBS 0.006909f
C242 B.n205 VSUBS 0.006909f
C243 B.n206 VSUBS 0.006909f
C244 B.n207 VSUBS 0.006909f
C245 B.n208 VSUBS 0.006909f
C246 B.n209 VSUBS 0.006909f
C247 B.n210 VSUBS 0.006909f
C248 B.n211 VSUBS 0.006909f
C249 B.n212 VSUBS 0.006909f
C250 B.n213 VSUBS 0.006909f
C251 B.n214 VSUBS 0.006909f
C252 B.n215 VSUBS 0.006909f
C253 B.n216 VSUBS 0.006909f
C254 B.n217 VSUBS 0.006909f
C255 B.n218 VSUBS 0.006909f
C256 B.n219 VSUBS 0.015157f
C257 B.n220 VSUBS 0.016338f
C258 B.n221 VSUBS 0.016338f
C259 B.n222 VSUBS 0.006909f
C260 B.n223 VSUBS 0.006909f
C261 B.n224 VSUBS 0.006909f
C262 B.n225 VSUBS 0.006909f
C263 B.n226 VSUBS 0.006909f
C264 B.n227 VSUBS 0.006909f
C265 B.n228 VSUBS 0.006909f
C266 B.n229 VSUBS 0.006909f
C267 B.n230 VSUBS 0.006909f
C268 B.n231 VSUBS 0.006909f
C269 B.n232 VSUBS 0.006909f
C270 B.n233 VSUBS 0.006909f
C271 B.n234 VSUBS 0.006909f
C272 B.n235 VSUBS 0.006909f
C273 B.n236 VSUBS 0.006909f
C274 B.n237 VSUBS 0.006909f
C275 B.n238 VSUBS 0.006909f
C276 B.n239 VSUBS 0.006909f
C277 B.n240 VSUBS 0.006909f
C278 B.n241 VSUBS 0.006909f
C279 B.n242 VSUBS 0.006909f
C280 B.n243 VSUBS 0.006909f
C281 B.n244 VSUBS 0.006909f
C282 B.n245 VSUBS 0.006909f
C283 B.n246 VSUBS 0.006909f
C284 B.n247 VSUBS 0.006909f
C285 B.n248 VSUBS 0.006909f
C286 B.n249 VSUBS 0.006909f
C287 B.n250 VSUBS 0.006909f
C288 B.n251 VSUBS 0.006909f
C289 B.n252 VSUBS 0.006909f
C290 B.n253 VSUBS 0.006909f
C291 B.n254 VSUBS 0.006909f
C292 B.n255 VSUBS 0.006909f
C293 B.n256 VSUBS 0.006909f
C294 B.n257 VSUBS 0.006909f
C295 B.n258 VSUBS 0.006909f
C296 B.n259 VSUBS 0.006909f
C297 B.n260 VSUBS 0.006909f
C298 B.n261 VSUBS 0.006909f
C299 B.n262 VSUBS 0.006909f
C300 B.n263 VSUBS 0.006909f
C301 B.n264 VSUBS 0.006909f
C302 B.n265 VSUBS 0.006909f
C303 B.n266 VSUBS 0.006502f
C304 B.n267 VSUBS 0.016007f
C305 B.n268 VSUBS 0.003861f
C306 B.n269 VSUBS 0.006909f
C307 B.n270 VSUBS 0.006909f
C308 B.n271 VSUBS 0.006909f
C309 B.n272 VSUBS 0.006909f
C310 B.n273 VSUBS 0.006909f
C311 B.n274 VSUBS 0.006909f
C312 B.n275 VSUBS 0.006909f
C313 B.n276 VSUBS 0.006909f
C314 B.n277 VSUBS 0.006909f
C315 B.n278 VSUBS 0.006909f
C316 B.n279 VSUBS 0.006909f
C317 B.n280 VSUBS 0.006909f
C318 B.t8 VSUBS 0.257808f
C319 B.t7 VSUBS 0.277085f
C320 B.t6 VSUBS 0.933044f
C321 B.n281 VSUBS 0.147267f
C322 B.n282 VSUBS 0.069857f
C323 B.n283 VSUBS 0.016007f
C324 B.n284 VSUBS 0.003861f
C325 B.n285 VSUBS 0.006909f
C326 B.n286 VSUBS 0.006909f
C327 B.n287 VSUBS 0.006909f
C328 B.n288 VSUBS 0.006909f
C329 B.n289 VSUBS 0.006909f
C330 B.n290 VSUBS 0.006909f
C331 B.n291 VSUBS 0.006909f
C332 B.n292 VSUBS 0.006909f
C333 B.n293 VSUBS 0.006909f
C334 B.n294 VSUBS 0.006909f
C335 B.n295 VSUBS 0.006909f
C336 B.n296 VSUBS 0.006909f
C337 B.n297 VSUBS 0.006909f
C338 B.n298 VSUBS 0.006909f
C339 B.n299 VSUBS 0.006909f
C340 B.n300 VSUBS 0.006909f
C341 B.n301 VSUBS 0.006909f
C342 B.n302 VSUBS 0.006909f
C343 B.n303 VSUBS 0.006909f
C344 B.n304 VSUBS 0.006909f
C345 B.n305 VSUBS 0.006909f
C346 B.n306 VSUBS 0.006909f
C347 B.n307 VSUBS 0.006909f
C348 B.n308 VSUBS 0.006909f
C349 B.n309 VSUBS 0.006909f
C350 B.n310 VSUBS 0.006909f
C351 B.n311 VSUBS 0.006909f
C352 B.n312 VSUBS 0.006909f
C353 B.n313 VSUBS 0.006909f
C354 B.n314 VSUBS 0.006909f
C355 B.n315 VSUBS 0.006909f
C356 B.n316 VSUBS 0.006909f
C357 B.n317 VSUBS 0.006909f
C358 B.n318 VSUBS 0.006909f
C359 B.n319 VSUBS 0.006909f
C360 B.n320 VSUBS 0.006909f
C361 B.n321 VSUBS 0.006909f
C362 B.n322 VSUBS 0.006909f
C363 B.n323 VSUBS 0.006909f
C364 B.n324 VSUBS 0.006909f
C365 B.n325 VSUBS 0.006909f
C366 B.n326 VSUBS 0.006909f
C367 B.n327 VSUBS 0.006909f
C368 B.n328 VSUBS 0.006909f
C369 B.n329 VSUBS 0.006909f
C370 B.n330 VSUBS 0.006909f
C371 B.n331 VSUBS 0.015489f
C372 B.n332 VSUBS 0.016007f
C373 B.n333 VSUBS 0.015157f
C374 B.n334 VSUBS 0.006909f
C375 B.n335 VSUBS 0.006909f
C376 B.n336 VSUBS 0.006909f
C377 B.n337 VSUBS 0.006909f
C378 B.n338 VSUBS 0.006909f
C379 B.n339 VSUBS 0.006909f
C380 B.n340 VSUBS 0.006909f
C381 B.n341 VSUBS 0.006909f
C382 B.n342 VSUBS 0.006909f
C383 B.n343 VSUBS 0.006909f
C384 B.n344 VSUBS 0.006909f
C385 B.n345 VSUBS 0.006909f
C386 B.n346 VSUBS 0.006909f
C387 B.n347 VSUBS 0.006909f
C388 B.n348 VSUBS 0.006909f
C389 B.n349 VSUBS 0.006909f
C390 B.n350 VSUBS 0.006909f
C391 B.n351 VSUBS 0.006909f
C392 B.n352 VSUBS 0.006909f
C393 B.n353 VSUBS 0.006909f
C394 B.n354 VSUBS 0.006909f
C395 B.n355 VSUBS 0.006909f
C396 B.n356 VSUBS 0.006909f
C397 B.n357 VSUBS 0.006909f
C398 B.n358 VSUBS 0.006909f
C399 B.n359 VSUBS 0.006909f
C400 B.n360 VSUBS 0.006909f
C401 B.n361 VSUBS 0.006909f
C402 B.n362 VSUBS 0.006909f
C403 B.n363 VSUBS 0.006909f
C404 B.n364 VSUBS 0.006909f
C405 B.n365 VSUBS 0.006909f
C406 B.n366 VSUBS 0.006909f
C407 B.n367 VSUBS 0.006909f
C408 B.n368 VSUBS 0.006909f
C409 B.n369 VSUBS 0.006909f
C410 B.n370 VSUBS 0.006909f
C411 B.n371 VSUBS 0.006909f
C412 B.n372 VSUBS 0.006909f
C413 B.n373 VSUBS 0.006909f
C414 B.n374 VSUBS 0.006909f
C415 B.n375 VSUBS 0.006909f
C416 B.n376 VSUBS 0.006909f
C417 B.n377 VSUBS 0.006909f
C418 B.n378 VSUBS 0.006909f
C419 B.n379 VSUBS 0.006909f
C420 B.n380 VSUBS 0.006909f
C421 B.n381 VSUBS 0.006909f
C422 B.n382 VSUBS 0.006909f
C423 B.n383 VSUBS 0.006909f
C424 B.n384 VSUBS 0.006909f
C425 B.n385 VSUBS 0.006909f
C426 B.n386 VSUBS 0.006909f
C427 B.n387 VSUBS 0.006909f
C428 B.n388 VSUBS 0.006909f
C429 B.n389 VSUBS 0.006909f
C430 B.n390 VSUBS 0.006909f
C431 B.n391 VSUBS 0.006909f
C432 B.n392 VSUBS 0.006909f
C433 B.n393 VSUBS 0.006909f
C434 B.n394 VSUBS 0.006909f
C435 B.n395 VSUBS 0.006909f
C436 B.n396 VSUBS 0.006909f
C437 B.n397 VSUBS 0.006909f
C438 B.n398 VSUBS 0.006909f
C439 B.n399 VSUBS 0.006909f
C440 B.n400 VSUBS 0.006909f
C441 B.n401 VSUBS 0.006909f
C442 B.n402 VSUBS 0.006909f
C443 B.n403 VSUBS 0.006909f
C444 B.n404 VSUBS 0.006909f
C445 B.n405 VSUBS 0.006909f
C446 B.n406 VSUBS 0.006909f
C447 B.n407 VSUBS 0.006909f
C448 B.n408 VSUBS 0.006909f
C449 B.n409 VSUBS 0.006909f
C450 B.n410 VSUBS 0.006909f
C451 B.n411 VSUBS 0.006909f
C452 B.n412 VSUBS 0.006909f
C453 B.n413 VSUBS 0.006909f
C454 B.n414 VSUBS 0.006909f
C455 B.n415 VSUBS 0.006909f
C456 B.n416 VSUBS 0.006909f
C457 B.n417 VSUBS 0.006909f
C458 B.n418 VSUBS 0.006909f
C459 B.n419 VSUBS 0.006909f
C460 B.n420 VSUBS 0.006909f
C461 B.n421 VSUBS 0.006909f
C462 B.n422 VSUBS 0.006909f
C463 B.n423 VSUBS 0.006909f
C464 B.n424 VSUBS 0.006909f
C465 B.n425 VSUBS 0.006909f
C466 B.n426 VSUBS 0.006909f
C467 B.n427 VSUBS 0.006909f
C468 B.n428 VSUBS 0.006909f
C469 B.n429 VSUBS 0.006909f
C470 B.n430 VSUBS 0.006909f
C471 B.n431 VSUBS 0.006909f
C472 B.n432 VSUBS 0.006909f
C473 B.n433 VSUBS 0.006909f
C474 B.n434 VSUBS 0.006909f
C475 B.n435 VSUBS 0.006909f
C476 B.n436 VSUBS 0.006909f
C477 B.n437 VSUBS 0.006909f
C478 B.n438 VSUBS 0.006909f
C479 B.n439 VSUBS 0.006909f
C480 B.n440 VSUBS 0.006909f
C481 B.n441 VSUBS 0.006909f
C482 B.n442 VSUBS 0.006909f
C483 B.n443 VSUBS 0.006909f
C484 B.n444 VSUBS 0.006909f
C485 B.n445 VSUBS 0.006909f
C486 B.n446 VSUBS 0.006909f
C487 B.n447 VSUBS 0.006909f
C488 B.n448 VSUBS 0.006909f
C489 B.n449 VSUBS 0.006909f
C490 B.n450 VSUBS 0.006909f
C491 B.n451 VSUBS 0.006909f
C492 B.n452 VSUBS 0.006909f
C493 B.n453 VSUBS 0.006909f
C494 B.n454 VSUBS 0.015157f
C495 B.n455 VSUBS 0.016338f
C496 B.n456 VSUBS 0.016338f
C497 B.n457 VSUBS 0.006909f
C498 B.n458 VSUBS 0.006909f
C499 B.n459 VSUBS 0.006909f
C500 B.n460 VSUBS 0.006909f
C501 B.n461 VSUBS 0.006909f
C502 B.n462 VSUBS 0.006909f
C503 B.n463 VSUBS 0.006909f
C504 B.n464 VSUBS 0.006909f
C505 B.n465 VSUBS 0.006909f
C506 B.n466 VSUBS 0.006909f
C507 B.n467 VSUBS 0.006909f
C508 B.n468 VSUBS 0.006909f
C509 B.n469 VSUBS 0.006909f
C510 B.n470 VSUBS 0.006909f
C511 B.n471 VSUBS 0.006909f
C512 B.n472 VSUBS 0.006909f
C513 B.n473 VSUBS 0.006909f
C514 B.n474 VSUBS 0.006909f
C515 B.n475 VSUBS 0.006909f
C516 B.n476 VSUBS 0.006909f
C517 B.n477 VSUBS 0.006909f
C518 B.n478 VSUBS 0.006909f
C519 B.n479 VSUBS 0.006909f
C520 B.n480 VSUBS 0.006909f
C521 B.n481 VSUBS 0.006909f
C522 B.n482 VSUBS 0.006909f
C523 B.n483 VSUBS 0.006909f
C524 B.n484 VSUBS 0.006909f
C525 B.n485 VSUBS 0.006909f
C526 B.n486 VSUBS 0.006909f
C527 B.n487 VSUBS 0.006909f
C528 B.n488 VSUBS 0.006909f
C529 B.n489 VSUBS 0.006909f
C530 B.n490 VSUBS 0.006909f
C531 B.n491 VSUBS 0.006909f
C532 B.n492 VSUBS 0.006909f
C533 B.n493 VSUBS 0.006909f
C534 B.n494 VSUBS 0.006909f
C535 B.n495 VSUBS 0.006909f
C536 B.n496 VSUBS 0.006909f
C537 B.n497 VSUBS 0.006909f
C538 B.n498 VSUBS 0.006909f
C539 B.n499 VSUBS 0.006909f
C540 B.n500 VSUBS 0.006502f
C541 B.n501 VSUBS 0.006909f
C542 B.n502 VSUBS 0.006909f
C543 B.n503 VSUBS 0.006909f
C544 B.n504 VSUBS 0.006909f
C545 B.n505 VSUBS 0.006909f
C546 B.n506 VSUBS 0.006909f
C547 B.n507 VSUBS 0.006909f
C548 B.n508 VSUBS 0.006909f
C549 B.n509 VSUBS 0.006909f
C550 B.n510 VSUBS 0.006909f
C551 B.n511 VSUBS 0.006909f
C552 B.n512 VSUBS 0.006909f
C553 B.n513 VSUBS 0.006909f
C554 B.n514 VSUBS 0.006909f
C555 B.n515 VSUBS 0.006909f
C556 B.n516 VSUBS 0.003861f
C557 B.n517 VSUBS 0.016007f
C558 B.n518 VSUBS 0.006502f
C559 B.n519 VSUBS 0.006909f
C560 B.n520 VSUBS 0.006909f
C561 B.n521 VSUBS 0.006909f
C562 B.n522 VSUBS 0.006909f
C563 B.n523 VSUBS 0.006909f
C564 B.n524 VSUBS 0.006909f
C565 B.n525 VSUBS 0.006909f
C566 B.n526 VSUBS 0.006909f
C567 B.n527 VSUBS 0.006909f
C568 B.n528 VSUBS 0.006909f
C569 B.n529 VSUBS 0.006909f
C570 B.n530 VSUBS 0.006909f
C571 B.n531 VSUBS 0.006909f
C572 B.n532 VSUBS 0.006909f
C573 B.n533 VSUBS 0.006909f
C574 B.n534 VSUBS 0.006909f
C575 B.n535 VSUBS 0.006909f
C576 B.n536 VSUBS 0.006909f
C577 B.n537 VSUBS 0.006909f
C578 B.n538 VSUBS 0.006909f
C579 B.n539 VSUBS 0.006909f
C580 B.n540 VSUBS 0.006909f
C581 B.n541 VSUBS 0.006909f
C582 B.n542 VSUBS 0.006909f
C583 B.n543 VSUBS 0.006909f
C584 B.n544 VSUBS 0.006909f
C585 B.n545 VSUBS 0.006909f
C586 B.n546 VSUBS 0.006909f
C587 B.n547 VSUBS 0.006909f
C588 B.n548 VSUBS 0.006909f
C589 B.n549 VSUBS 0.006909f
C590 B.n550 VSUBS 0.006909f
C591 B.n551 VSUBS 0.006909f
C592 B.n552 VSUBS 0.006909f
C593 B.n553 VSUBS 0.006909f
C594 B.n554 VSUBS 0.006909f
C595 B.n555 VSUBS 0.006909f
C596 B.n556 VSUBS 0.006909f
C597 B.n557 VSUBS 0.006909f
C598 B.n558 VSUBS 0.006909f
C599 B.n559 VSUBS 0.006909f
C600 B.n560 VSUBS 0.006909f
C601 B.n561 VSUBS 0.006909f
C602 B.n562 VSUBS 0.006909f
C603 B.n563 VSUBS 0.016338f
C604 B.n564 VSUBS 0.015157f
C605 B.n565 VSUBS 0.015157f
C606 B.n566 VSUBS 0.006909f
C607 B.n567 VSUBS 0.006909f
C608 B.n568 VSUBS 0.006909f
C609 B.n569 VSUBS 0.006909f
C610 B.n570 VSUBS 0.006909f
C611 B.n571 VSUBS 0.006909f
C612 B.n572 VSUBS 0.006909f
C613 B.n573 VSUBS 0.006909f
C614 B.n574 VSUBS 0.006909f
C615 B.n575 VSUBS 0.006909f
C616 B.n576 VSUBS 0.006909f
C617 B.n577 VSUBS 0.006909f
C618 B.n578 VSUBS 0.006909f
C619 B.n579 VSUBS 0.006909f
C620 B.n580 VSUBS 0.006909f
C621 B.n581 VSUBS 0.006909f
C622 B.n582 VSUBS 0.006909f
C623 B.n583 VSUBS 0.006909f
C624 B.n584 VSUBS 0.006909f
C625 B.n585 VSUBS 0.006909f
C626 B.n586 VSUBS 0.006909f
C627 B.n587 VSUBS 0.006909f
C628 B.n588 VSUBS 0.006909f
C629 B.n589 VSUBS 0.006909f
C630 B.n590 VSUBS 0.006909f
C631 B.n591 VSUBS 0.006909f
C632 B.n592 VSUBS 0.006909f
C633 B.n593 VSUBS 0.006909f
C634 B.n594 VSUBS 0.006909f
C635 B.n595 VSUBS 0.006909f
C636 B.n596 VSUBS 0.006909f
C637 B.n597 VSUBS 0.006909f
C638 B.n598 VSUBS 0.006909f
C639 B.n599 VSUBS 0.006909f
C640 B.n600 VSUBS 0.006909f
C641 B.n601 VSUBS 0.006909f
C642 B.n602 VSUBS 0.006909f
C643 B.n603 VSUBS 0.006909f
C644 B.n604 VSUBS 0.006909f
C645 B.n605 VSUBS 0.006909f
C646 B.n606 VSUBS 0.006909f
C647 B.n607 VSUBS 0.006909f
C648 B.n608 VSUBS 0.006909f
C649 B.n609 VSUBS 0.006909f
C650 B.n610 VSUBS 0.006909f
C651 B.n611 VSUBS 0.006909f
C652 B.n612 VSUBS 0.006909f
C653 B.n613 VSUBS 0.006909f
C654 B.n614 VSUBS 0.006909f
C655 B.n615 VSUBS 0.006909f
C656 B.n616 VSUBS 0.006909f
C657 B.n617 VSUBS 0.006909f
C658 B.n618 VSUBS 0.006909f
C659 B.n619 VSUBS 0.006909f
C660 B.n620 VSUBS 0.006909f
C661 B.n621 VSUBS 0.006909f
C662 B.n622 VSUBS 0.006909f
C663 B.n623 VSUBS 0.009015f
C664 B.n624 VSUBS 0.009604f
C665 B.n625 VSUBS 0.019098f
C666 VDD1.t3 VSUBS 1.39217f
C667 VDD1.t5 VSUBS 1.39123f
C668 VDD1.t4 VSUBS 0.145341f
C669 VDD1.t2 VSUBS 0.145341f
C670 VDD1.n0 VSUBS 1.04719f
C671 VDD1.n1 VSUBS 2.82187f
C672 VDD1.t0 VSUBS 0.145341f
C673 VDD1.t1 VSUBS 0.145341f
C674 VDD1.n2 VSUBS 1.04306f
C675 VDD1.n3 VSUBS 2.37355f
C676 VP.n0 VSUBS 0.047457f
C677 VP.t3 VSUBS 1.97728f
C678 VP.n1 VSUBS 0.036445f
C679 VP.n2 VSUBS 0.035994f
C680 VP.t1 VSUBS 1.97728f
C681 VP.n3 VSUBS 0.067419f
C682 VP.n4 VSUBS 0.035994f
C683 VP.n5 VSUBS 0.051441f
C684 VP.n6 VSUBS 0.047457f
C685 VP.t4 VSUBS 1.97728f
C686 VP.n7 VSUBS 0.036445f
C687 VP.n8 VSUBS 0.341811f
C688 VP.t5 VSUBS 1.97728f
C689 VP.t2 VSUBS 2.25129f
C690 VP.n9 VSUBS 0.791216f
C691 VP.n10 VSUBS 0.83957f
C692 VP.n11 VSUBS 0.067419f
C693 VP.n12 VSUBS 0.064937f
C694 VP.n13 VSUBS 0.035994f
C695 VP.n14 VSUBS 0.035994f
C696 VP.n15 VSUBS 0.035994f
C697 VP.n16 VSUBS 0.071583f
C698 VP.n17 VSUBS 0.051441f
C699 VP.n18 VSUBS 0.838262f
C700 VP.n19 VSUBS 1.7218f
C701 VP.t0 VSUBS 1.97728f
C702 VP.n20 VSUBS 0.838262f
C703 VP.n21 VSUBS 1.75028f
C704 VP.n22 VSUBS 0.047457f
C705 VP.n23 VSUBS 0.035994f
C706 VP.n24 VSUBS 0.071583f
C707 VP.n25 VSUBS 0.036445f
C708 VP.n26 VSUBS 0.064937f
C709 VP.n27 VSUBS 0.035994f
C710 VP.n28 VSUBS 0.035994f
C711 VP.n29 VSUBS 0.035994f
C712 VP.n30 VSUBS 0.753747f
C713 VP.n31 VSUBS 0.067419f
C714 VP.n32 VSUBS 0.064937f
C715 VP.n33 VSUBS 0.035994f
C716 VP.n34 VSUBS 0.035994f
C717 VP.n35 VSUBS 0.035994f
C718 VP.n36 VSUBS 0.071583f
C719 VP.n37 VSUBS 0.051441f
C720 VP.n38 VSUBS 0.838262f
C721 VP.n39 VSUBS 0.0542f
C722 VTAIL.t6 VSUBS 0.20348f
C723 VTAIL.t8 VSUBS 0.20348f
C724 VTAIL.n0 VSUBS 1.31451f
C725 VTAIL.n1 VSUBS 0.88639f
C726 VTAIL.t0 VSUBS 1.7726f
C727 VTAIL.n2 VSUBS 1.15376f
C728 VTAIL.t3 VSUBS 0.20348f
C729 VTAIL.t5 VSUBS 0.20348f
C730 VTAIL.n3 VSUBS 1.31451f
C731 VTAIL.n4 VSUBS 2.49468f
C732 VTAIL.t7 VSUBS 0.20348f
C733 VTAIL.t11 VSUBS 0.20348f
C734 VTAIL.n5 VSUBS 1.31451f
C735 VTAIL.n6 VSUBS 2.49468f
C736 VTAIL.t10 VSUBS 1.77261f
C737 VTAIL.n7 VSUBS 1.15375f
C738 VTAIL.t4 VSUBS 0.20348f
C739 VTAIL.t2 VSUBS 0.20348f
C740 VTAIL.n8 VSUBS 1.31451f
C741 VTAIL.n9 VSUBS 1.0569f
C742 VTAIL.t1 VSUBS 1.77261f
C743 VTAIL.n10 VSUBS 2.35651f
C744 VTAIL.t9 VSUBS 1.7726f
C745 VTAIL.n11 VSUBS 2.29202f
C746 VDD2.t3 VSUBS 1.63469f
C747 VDD2.t1 VSUBS 0.170776f
C748 VDD2.t2 VSUBS 0.170776f
C749 VDD2.n0 VSUBS 1.23045f
C750 VDD2.n1 VSUBS 3.19559f
C751 VDD2.t5 VSUBS 1.62067f
C752 VDD2.n2 VSUBS 2.79573f
C753 VDD2.t0 VSUBS 0.170776f
C754 VDD2.t4 VSUBS 0.170776f
C755 VDD2.n3 VSUBS 1.23042f
C756 VN.n0 VSUBS 0.046082f
C757 VN.t2 VSUBS 1.91998f
C758 VN.n1 VSUBS 0.035389f
C759 VN.n2 VSUBS 0.331905f
C760 VN.t3 VSUBS 1.91998f
C761 VN.t5 VSUBS 2.18605f
C762 VN.n3 VSUBS 0.768287f
C763 VN.n4 VSUBS 0.81524f
C764 VN.n5 VSUBS 0.065466f
C765 VN.n6 VSUBS 0.063055f
C766 VN.n7 VSUBS 0.034951f
C767 VN.n8 VSUBS 0.034951f
C768 VN.n9 VSUBS 0.034951f
C769 VN.n10 VSUBS 0.069509f
C770 VN.n11 VSUBS 0.049951f
C771 VN.n12 VSUBS 0.81397f
C772 VN.n13 VSUBS 0.052629f
C773 VN.n14 VSUBS 0.046082f
C774 VN.t4 VSUBS 1.91998f
C775 VN.n15 VSUBS 0.035389f
C776 VN.n16 VSUBS 0.331905f
C777 VN.t0 VSUBS 1.91998f
C778 VN.t1 VSUBS 2.18605f
C779 VN.n17 VSUBS 0.768287f
C780 VN.n18 VSUBS 0.81524f
C781 VN.n19 VSUBS 0.065466f
C782 VN.n20 VSUBS 0.063055f
C783 VN.n21 VSUBS 0.034951f
C784 VN.n22 VSUBS 0.034951f
C785 VN.n23 VSUBS 0.034951f
C786 VN.n24 VSUBS 0.069509f
C787 VN.n25 VSUBS 0.049951f
C788 VN.n26 VSUBS 0.81397f
C789 VN.n27 VSUBS 1.69099f
.ends

