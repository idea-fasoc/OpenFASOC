* NGSPICE file created from diff_pair_sample_1165.ext - technology: sky130A

.subckt diff_pair_sample_1165 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t7 VN.t0 VDD2.t0 w_n2674_n3956# sky130_fd_pr__pfet_01v8 ad=5.8266 pd=30.66 as=2.4651 ps=15.27 w=14.94 l=2.51
X1 B.t11 B.t9 B.t10 w_n2674_n3956# sky130_fd_pr__pfet_01v8 ad=5.8266 pd=30.66 as=0 ps=0 w=14.94 l=2.51
X2 B.t8 B.t6 B.t7 w_n2674_n3956# sky130_fd_pr__pfet_01v8 ad=5.8266 pd=30.66 as=0 ps=0 w=14.94 l=2.51
X3 VTAIL.t2 VP.t0 VDD1.t3 w_n2674_n3956# sky130_fd_pr__pfet_01v8 ad=5.8266 pd=30.66 as=2.4651 ps=15.27 w=14.94 l=2.51
X4 VTAIL.t3 VP.t1 VDD1.t2 w_n2674_n3956# sky130_fd_pr__pfet_01v8 ad=5.8266 pd=30.66 as=2.4651 ps=15.27 w=14.94 l=2.51
X5 VDD2.t1 VN.t1 VTAIL.t6 w_n2674_n3956# sky130_fd_pr__pfet_01v8 ad=2.4651 pd=15.27 as=5.8266 ps=30.66 w=14.94 l=2.51
X6 VDD2.t2 VN.t2 VTAIL.t5 w_n2674_n3956# sky130_fd_pr__pfet_01v8 ad=2.4651 pd=15.27 as=5.8266 ps=30.66 w=14.94 l=2.51
X7 VDD1.t1 VP.t2 VTAIL.t0 w_n2674_n3956# sky130_fd_pr__pfet_01v8 ad=2.4651 pd=15.27 as=5.8266 ps=30.66 w=14.94 l=2.51
X8 B.t5 B.t3 B.t4 w_n2674_n3956# sky130_fd_pr__pfet_01v8 ad=5.8266 pd=30.66 as=0 ps=0 w=14.94 l=2.51
X9 B.t2 B.t0 B.t1 w_n2674_n3956# sky130_fd_pr__pfet_01v8 ad=5.8266 pd=30.66 as=0 ps=0 w=14.94 l=2.51
X10 VDD1.t0 VP.t3 VTAIL.t1 w_n2674_n3956# sky130_fd_pr__pfet_01v8 ad=2.4651 pd=15.27 as=5.8266 ps=30.66 w=14.94 l=2.51
X11 VTAIL.t4 VN.t3 VDD2.t3 w_n2674_n3956# sky130_fd_pr__pfet_01v8 ad=5.8266 pd=30.66 as=2.4651 ps=15.27 w=14.94 l=2.51
R0 VN.n0 VN.t3 179.035
R1 VN.n1 VN.t1 179.035
R2 VN.n0 VN.t2 178.274
R3 VN.n1 VN.t0 178.274
R4 VN VN.n1 52.9915
R5 VN VN.n0 4.49533
R6 VDD2.n2 VDD2.n0 113.831
R7 VDD2.n2 VDD2.n1 69.892
R8 VDD2.n1 VDD2.t0 2.1762
R9 VDD2.n1 VDD2.t1 2.1762
R10 VDD2.n0 VDD2.t3 2.1762
R11 VDD2.n0 VDD2.t2 2.1762
R12 VDD2 VDD2.n2 0.0586897
R13 VTAIL.n650 VTAIL.n574 756.745
R14 VTAIL.n76 VTAIL.n0 756.745
R15 VTAIL.n158 VTAIL.n82 756.745
R16 VTAIL.n240 VTAIL.n164 756.745
R17 VTAIL.n568 VTAIL.n492 756.745
R18 VTAIL.n486 VTAIL.n410 756.745
R19 VTAIL.n404 VTAIL.n328 756.745
R20 VTAIL.n322 VTAIL.n246 756.745
R21 VTAIL.n601 VTAIL.n600 585
R22 VTAIL.n598 VTAIL.n597 585
R23 VTAIL.n607 VTAIL.n606 585
R24 VTAIL.n609 VTAIL.n608 585
R25 VTAIL.n594 VTAIL.n593 585
R26 VTAIL.n615 VTAIL.n614 585
R27 VTAIL.n618 VTAIL.n617 585
R28 VTAIL.n616 VTAIL.n590 585
R29 VTAIL.n623 VTAIL.n589 585
R30 VTAIL.n625 VTAIL.n624 585
R31 VTAIL.n627 VTAIL.n626 585
R32 VTAIL.n586 VTAIL.n585 585
R33 VTAIL.n633 VTAIL.n632 585
R34 VTAIL.n635 VTAIL.n634 585
R35 VTAIL.n582 VTAIL.n581 585
R36 VTAIL.n641 VTAIL.n640 585
R37 VTAIL.n643 VTAIL.n642 585
R38 VTAIL.n578 VTAIL.n577 585
R39 VTAIL.n649 VTAIL.n648 585
R40 VTAIL.n651 VTAIL.n650 585
R41 VTAIL.n27 VTAIL.n26 585
R42 VTAIL.n24 VTAIL.n23 585
R43 VTAIL.n33 VTAIL.n32 585
R44 VTAIL.n35 VTAIL.n34 585
R45 VTAIL.n20 VTAIL.n19 585
R46 VTAIL.n41 VTAIL.n40 585
R47 VTAIL.n44 VTAIL.n43 585
R48 VTAIL.n42 VTAIL.n16 585
R49 VTAIL.n49 VTAIL.n15 585
R50 VTAIL.n51 VTAIL.n50 585
R51 VTAIL.n53 VTAIL.n52 585
R52 VTAIL.n12 VTAIL.n11 585
R53 VTAIL.n59 VTAIL.n58 585
R54 VTAIL.n61 VTAIL.n60 585
R55 VTAIL.n8 VTAIL.n7 585
R56 VTAIL.n67 VTAIL.n66 585
R57 VTAIL.n69 VTAIL.n68 585
R58 VTAIL.n4 VTAIL.n3 585
R59 VTAIL.n75 VTAIL.n74 585
R60 VTAIL.n77 VTAIL.n76 585
R61 VTAIL.n109 VTAIL.n108 585
R62 VTAIL.n106 VTAIL.n105 585
R63 VTAIL.n115 VTAIL.n114 585
R64 VTAIL.n117 VTAIL.n116 585
R65 VTAIL.n102 VTAIL.n101 585
R66 VTAIL.n123 VTAIL.n122 585
R67 VTAIL.n126 VTAIL.n125 585
R68 VTAIL.n124 VTAIL.n98 585
R69 VTAIL.n131 VTAIL.n97 585
R70 VTAIL.n133 VTAIL.n132 585
R71 VTAIL.n135 VTAIL.n134 585
R72 VTAIL.n94 VTAIL.n93 585
R73 VTAIL.n141 VTAIL.n140 585
R74 VTAIL.n143 VTAIL.n142 585
R75 VTAIL.n90 VTAIL.n89 585
R76 VTAIL.n149 VTAIL.n148 585
R77 VTAIL.n151 VTAIL.n150 585
R78 VTAIL.n86 VTAIL.n85 585
R79 VTAIL.n157 VTAIL.n156 585
R80 VTAIL.n159 VTAIL.n158 585
R81 VTAIL.n191 VTAIL.n190 585
R82 VTAIL.n188 VTAIL.n187 585
R83 VTAIL.n197 VTAIL.n196 585
R84 VTAIL.n199 VTAIL.n198 585
R85 VTAIL.n184 VTAIL.n183 585
R86 VTAIL.n205 VTAIL.n204 585
R87 VTAIL.n208 VTAIL.n207 585
R88 VTAIL.n206 VTAIL.n180 585
R89 VTAIL.n213 VTAIL.n179 585
R90 VTAIL.n215 VTAIL.n214 585
R91 VTAIL.n217 VTAIL.n216 585
R92 VTAIL.n176 VTAIL.n175 585
R93 VTAIL.n223 VTAIL.n222 585
R94 VTAIL.n225 VTAIL.n224 585
R95 VTAIL.n172 VTAIL.n171 585
R96 VTAIL.n231 VTAIL.n230 585
R97 VTAIL.n233 VTAIL.n232 585
R98 VTAIL.n168 VTAIL.n167 585
R99 VTAIL.n239 VTAIL.n238 585
R100 VTAIL.n241 VTAIL.n240 585
R101 VTAIL.n569 VTAIL.n568 585
R102 VTAIL.n567 VTAIL.n566 585
R103 VTAIL.n496 VTAIL.n495 585
R104 VTAIL.n561 VTAIL.n560 585
R105 VTAIL.n559 VTAIL.n558 585
R106 VTAIL.n500 VTAIL.n499 585
R107 VTAIL.n553 VTAIL.n552 585
R108 VTAIL.n551 VTAIL.n550 585
R109 VTAIL.n504 VTAIL.n503 585
R110 VTAIL.n545 VTAIL.n544 585
R111 VTAIL.n543 VTAIL.n542 585
R112 VTAIL.n541 VTAIL.n507 585
R113 VTAIL.n511 VTAIL.n508 585
R114 VTAIL.n536 VTAIL.n535 585
R115 VTAIL.n534 VTAIL.n533 585
R116 VTAIL.n513 VTAIL.n512 585
R117 VTAIL.n528 VTAIL.n527 585
R118 VTAIL.n526 VTAIL.n525 585
R119 VTAIL.n517 VTAIL.n516 585
R120 VTAIL.n520 VTAIL.n519 585
R121 VTAIL.n487 VTAIL.n486 585
R122 VTAIL.n485 VTAIL.n484 585
R123 VTAIL.n414 VTAIL.n413 585
R124 VTAIL.n479 VTAIL.n478 585
R125 VTAIL.n477 VTAIL.n476 585
R126 VTAIL.n418 VTAIL.n417 585
R127 VTAIL.n471 VTAIL.n470 585
R128 VTAIL.n469 VTAIL.n468 585
R129 VTAIL.n422 VTAIL.n421 585
R130 VTAIL.n463 VTAIL.n462 585
R131 VTAIL.n461 VTAIL.n460 585
R132 VTAIL.n459 VTAIL.n425 585
R133 VTAIL.n429 VTAIL.n426 585
R134 VTAIL.n454 VTAIL.n453 585
R135 VTAIL.n452 VTAIL.n451 585
R136 VTAIL.n431 VTAIL.n430 585
R137 VTAIL.n446 VTAIL.n445 585
R138 VTAIL.n444 VTAIL.n443 585
R139 VTAIL.n435 VTAIL.n434 585
R140 VTAIL.n438 VTAIL.n437 585
R141 VTAIL.n405 VTAIL.n404 585
R142 VTAIL.n403 VTAIL.n402 585
R143 VTAIL.n332 VTAIL.n331 585
R144 VTAIL.n397 VTAIL.n396 585
R145 VTAIL.n395 VTAIL.n394 585
R146 VTAIL.n336 VTAIL.n335 585
R147 VTAIL.n389 VTAIL.n388 585
R148 VTAIL.n387 VTAIL.n386 585
R149 VTAIL.n340 VTAIL.n339 585
R150 VTAIL.n381 VTAIL.n380 585
R151 VTAIL.n379 VTAIL.n378 585
R152 VTAIL.n377 VTAIL.n343 585
R153 VTAIL.n347 VTAIL.n344 585
R154 VTAIL.n372 VTAIL.n371 585
R155 VTAIL.n370 VTAIL.n369 585
R156 VTAIL.n349 VTAIL.n348 585
R157 VTAIL.n364 VTAIL.n363 585
R158 VTAIL.n362 VTAIL.n361 585
R159 VTAIL.n353 VTAIL.n352 585
R160 VTAIL.n356 VTAIL.n355 585
R161 VTAIL.n323 VTAIL.n322 585
R162 VTAIL.n321 VTAIL.n320 585
R163 VTAIL.n250 VTAIL.n249 585
R164 VTAIL.n315 VTAIL.n314 585
R165 VTAIL.n313 VTAIL.n312 585
R166 VTAIL.n254 VTAIL.n253 585
R167 VTAIL.n307 VTAIL.n306 585
R168 VTAIL.n305 VTAIL.n304 585
R169 VTAIL.n258 VTAIL.n257 585
R170 VTAIL.n299 VTAIL.n298 585
R171 VTAIL.n297 VTAIL.n296 585
R172 VTAIL.n295 VTAIL.n261 585
R173 VTAIL.n265 VTAIL.n262 585
R174 VTAIL.n290 VTAIL.n289 585
R175 VTAIL.n288 VTAIL.n287 585
R176 VTAIL.n267 VTAIL.n266 585
R177 VTAIL.n282 VTAIL.n281 585
R178 VTAIL.n280 VTAIL.n279 585
R179 VTAIL.n271 VTAIL.n270 585
R180 VTAIL.n274 VTAIL.n273 585
R181 VTAIL.t5 VTAIL.n599 329.036
R182 VTAIL.t4 VTAIL.n25 329.036
R183 VTAIL.t0 VTAIL.n107 329.036
R184 VTAIL.t3 VTAIL.n189 329.036
R185 VTAIL.t1 VTAIL.n518 329.036
R186 VTAIL.t2 VTAIL.n436 329.036
R187 VTAIL.t6 VTAIL.n354 329.036
R188 VTAIL.t7 VTAIL.n272 329.036
R189 VTAIL.n600 VTAIL.n597 171.744
R190 VTAIL.n607 VTAIL.n597 171.744
R191 VTAIL.n608 VTAIL.n607 171.744
R192 VTAIL.n608 VTAIL.n593 171.744
R193 VTAIL.n615 VTAIL.n593 171.744
R194 VTAIL.n617 VTAIL.n615 171.744
R195 VTAIL.n617 VTAIL.n616 171.744
R196 VTAIL.n616 VTAIL.n589 171.744
R197 VTAIL.n625 VTAIL.n589 171.744
R198 VTAIL.n626 VTAIL.n625 171.744
R199 VTAIL.n626 VTAIL.n585 171.744
R200 VTAIL.n633 VTAIL.n585 171.744
R201 VTAIL.n634 VTAIL.n633 171.744
R202 VTAIL.n634 VTAIL.n581 171.744
R203 VTAIL.n641 VTAIL.n581 171.744
R204 VTAIL.n642 VTAIL.n641 171.744
R205 VTAIL.n642 VTAIL.n577 171.744
R206 VTAIL.n649 VTAIL.n577 171.744
R207 VTAIL.n650 VTAIL.n649 171.744
R208 VTAIL.n26 VTAIL.n23 171.744
R209 VTAIL.n33 VTAIL.n23 171.744
R210 VTAIL.n34 VTAIL.n33 171.744
R211 VTAIL.n34 VTAIL.n19 171.744
R212 VTAIL.n41 VTAIL.n19 171.744
R213 VTAIL.n43 VTAIL.n41 171.744
R214 VTAIL.n43 VTAIL.n42 171.744
R215 VTAIL.n42 VTAIL.n15 171.744
R216 VTAIL.n51 VTAIL.n15 171.744
R217 VTAIL.n52 VTAIL.n51 171.744
R218 VTAIL.n52 VTAIL.n11 171.744
R219 VTAIL.n59 VTAIL.n11 171.744
R220 VTAIL.n60 VTAIL.n59 171.744
R221 VTAIL.n60 VTAIL.n7 171.744
R222 VTAIL.n67 VTAIL.n7 171.744
R223 VTAIL.n68 VTAIL.n67 171.744
R224 VTAIL.n68 VTAIL.n3 171.744
R225 VTAIL.n75 VTAIL.n3 171.744
R226 VTAIL.n76 VTAIL.n75 171.744
R227 VTAIL.n108 VTAIL.n105 171.744
R228 VTAIL.n115 VTAIL.n105 171.744
R229 VTAIL.n116 VTAIL.n115 171.744
R230 VTAIL.n116 VTAIL.n101 171.744
R231 VTAIL.n123 VTAIL.n101 171.744
R232 VTAIL.n125 VTAIL.n123 171.744
R233 VTAIL.n125 VTAIL.n124 171.744
R234 VTAIL.n124 VTAIL.n97 171.744
R235 VTAIL.n133 VTAIL.n97 171.744
R236 VTAIL.n134 VTAIL.n133 171.744
R237 VTAIL.n134 VTAIL.n93 171.744
R238 VTAIL.n141 VTAIL.n93 171.744
R239 VTAIL.n142 VTAIL.n141 171.744
R240 VTAIL.n142 VTAIL.n89 171.744
R241 VTAIL.n149 VTAIL.n89 171.744
R242 VTAIL.n150 VTAIL.n149 171.744
R243 VTAIL.n150 VTAIL.n85 171.744
R244 VTAIL.n157 VTAIL.n85 171.744
R245 VTAIL.n158 VTAIL.n157 171.744
R246 VTAIL.n190 VTAIL.n187 171.744
R247 VTAIL.n197 VTAIL.n187 171.744
R248 VTAIL.n198 VTAIL.n197 171.744
R249 VTAIL.n198 VTAIL.n183 171.744
R250 VTAIL.n205 VTAIL.n183 171.744
R251 VTAIL.n207 VTAIL.n205 171.744
R252 VTAIL.n207 VTAIL.n206 171.744
R253 VTAIL.n206 VTAIL.n179 171.744
R254 VTAIL.n215 VTAIL.n179 171.744
R255 VTAIL.n216 VTAIL.n215 171.744
R256 VTAIL.n216 VTAIL.n175 171.744
R257 VTAIL.n223 VTAIL.n175 171.744
R258 VTAIL.n224 VTAIL.n223 171.744
R259 VTAIL.n224 VTAIL.n171 171.744
R260 VTAIL.n231 VTAIL.n171 171.744
R261 VTAIL.n232 VTAIL.n231 171.744
R262 VTAIL.n232 VTAIL.n167 171.744
R263 VTAIL.n239 VTAIL.n167 171.744
R264 VTAIL.n240 VTAIL.n239 171.744
R265 VTAIL.n568 VTAIL.n567 171.744
R266 VTAIL.n567 VTAIL.n495 171.744
R267 VTAIL.n560 VTAIL.n495 171.744
R268 VTAIL.n560 VTAIL.n559 171.744
R269 VTAIL.n559 VTAIL.n499 171.744
R270 VTAIL.n552 VTAIL.n499 171.744
R271 VTAIL.n552 VTAIL.n551 171.744
R272 VTAIL.n551 VTAIL.n503 171.744
R273 VTAIL.n544 VTAIL.n503 171.744
R274 VTAIL.n544 VTAIL.n543 171.744
R275 VTAIL.n543 VTAIL.n507 171.744
R276 VTAIL.n511 VTAIL.n507 171.744
R277 VTAIL.n535 VTAIL.n511 171.744
R278 VTAIL.n535 VTAIL.n534 171.744
R279 VTAIL.n534 VTAIL.n512 171.744
R280 VTAIL.n527 VTAIL.n512 171.744
R281 VTAIL.n527 VTAIL.n526 171.744
R282 VTAIL.n526 VTAIL.n516 171.744
R283 VTAIL.n519 VTAIL.n516 171.744
R284 VTAIL.n486 VTAIL.n485 171.744
R285 VTAIL.n485 VTAIL.n413 171.744
R286 VTAIL.n478 VTAIL.n413 171.744
R287 VTAIL.n478 VTAIL.n477 171.744
R288 VTAIL.n477 VTAIL.n417 171.744
R289 VTAIL.n470 VTAIL.n417 171.744
R290 VTAIL.n470 VTAIL.n469 171.744
R291 VTAIL.n469 VTAIL.n421 171.744
R292 VTAIL.n462 VTAIL.n421 171.744
R293 VTAIL.n462 VTAIL.n461 171.744
R294 VTAIL.n461 VTAIL.n425 171.744
R295 VTAIL.n429 VTAIL.n425 171.744
R296 VTAIL.n453 VTAIL.n429 171.744
R297 VTAIL.n453 VTAIL.n452 171.744
R298 VTAIL.n452 VTAIL.n430 171.744
R299 VTAIL.n445 VTAIL.n430 171.744
R300 VTAIL.n445 VTAIL.n444 171.744
R301 VTAIL.n444 VTAIL.n434 171.744
R302 VTAIL.n437 VTAIL.n434 171.744
R303 VTAIL.n404 VTAIL.n403 171.744
R304 VTAIL.n403 VTAIL.n331 171.744
R305 VTAIL.n396 VTAIL.n331 171.744
R306 VTAIL.n396 VTAIL.n395 171.744
R307 VTAIL.n395 VTAIL.n335 171.744
R308 VTAIL.n388 VTAIL.n335 171.744
R309 VTAIL.n388 VTAIL.n387 171.744
R310 VTAIL.n387 VTAIL.n339 171.744
R311 VTAIL.n380 VTAIL.n339 171.744
R312 VTAIL.n380 VTAIL.n379 171.744
R313 VTAIL.n379 VTAIL.n343 171.744
R314 VTAIL.n347 VTAIL.n343 171.744
R315 VTAIL.n371 VTAIL.n347 171.744
R316 VTAIL.n371 VTAIL.n370 171.744
R317 VTAIL.n370 VTAIL.n348 171.744
R318 VTAIL.n363 VTAIL.n348 171.744
R319 VTAIL.n363 VTAIL.n362 171.744
R320 VTAIL.n362 VTAIL.n352 171.744
R321 VTAIL.n355 VTAIL.n352 171.744
R322 VTAIL.n322 VTAIL.n321 171.744
R323 VTAIL.n321 VTAIL.n249 171.744
R324 VTAIL.n314 VTAIL.n249 171.744
R325 VTAIL.n314 VTAIL.n313 171.744
R326 VTAIL.n313 VTAIL.n253 171.744
R327 VTAIL.n306 VTAIL.n253 171.744
R328 VTAIL.n306 VTAIL.n305 171.744
R329 VTAIL.n305 VTAIL.n257 171.744
R330 VTAIL.n298 VTAIL.n257 171.744
R331 VTAIL.n298 VTAIL.n297 171.744
R332 VTAIL.n297 VTAIL.n261 171.744
R333 VTAIL.n265 VTAIL.n261 171.744
R334 VTAIL.n289 VTAIL.n265 171.744
R335 VTAIL.n289 VTAIL.n288 171.744
R336 VTAIL.n288 VTAIL.n266 171.744
R337 VTAIL.n281 VTAIL.n266 171.744
R338 VTAIL.n281 VTAIL.n280 171.744
R339 VTAIL.n280 VTAIL.n270 171.744
R340 VTAIL.n273 VTAIL.n270 171.744
R341 VTAIL.n600 VTAIL.t5 85.8723
R342 VTAIL.n26 VTAIL.t4 85.8723
R343 VTAIL.n108 VTAIL.t0 85.8723
R344 VTAIL.n190 VTAIL.t3 85.8723
R345 VTAIL.n519 VTAIL.t1 85.8723
R346 VTAIL.n437 VTAIL.t2 85.8723
R347 VTAIL.n355 VTAIL.t6 85.8723
R348 VTAIL.n273 VTAIL.t7 85.8723
R349 VTAIL.n655 VTAIL.n654 31.0217
R350 VTAIL.n81 VTAIL.n80 31.0217
R351 VTAIL.n163 VTAIL.n162 31.0217
R352 VTAIL.n245 VTAIL.n244 31.0217
R353 VTAIL.n573 VTAIL.n572 31.0217
R354 VTAIL.n491 VTAIL.n490 31.0217
R355 VTAIL.n409 VTAIL.n408 31.0217
R356 VTAIL.n327 VTAIL.n326 31.0217
R357 VTAIL.n655 VTAIL.n573 27.6945
R358 VTAIL.n327 VTAIL.n245 27.6945
R359 VTAIL.n624 VTAIL.n623 13.1884
R360 VTAIL.n50 VTAIL.n49 13.1884
R361 VTAIL.n132 VTAIL.n131 13.1884
R362 VTAIL.n214 VTAIL.n213 13.1884
R363 VTAIL.n542 VTAIL.n541 13.1884
R364 VTAIL.n460 VTAIL.n459 13.1884
R365 VTAIL.n378 VTAIL.n377 13.1884
R366 VTAIL.n296 VTAIL.n295 13.1884
R367 VTAIL.n622 VTAIL.n590 12.8005
R368 VTAIL.n627 VTAIL.n588 12.8005
R369 VTAIL.n48 VTAIL.n16 12.8005
R370 VTAIL.n53 VTAIL.n14 12.8005
R371 VTAIL.n130 VTAIL.n98 12.8005
R372 VTAIL.n135 VTAIL.n96 12.8005
R373 VTAIL.n212 VTAIL.n180 12.8005
R374 VTAIL.n217 VTAIL.n178 12.8005
R375 VTAIL.n545 VTAIL.n506 12.8005
R376 VTAIL.n540 VTAIL.n508 12.8005
R377 VTAIL.n463 VTAIL.n424 12.8005
R378 VTAIL.n458 VTAIL.n426 12.8005
R379 VTAIL.n381 VTAIL.n342 12.8005
R380 VTAIL.n376 VTAIL.n344 12.8005
R381 VTAIL.n299 VTAIL.n260 12.8005
R382 VTAIL.n294 VTAIL.n262 12.8005
R383 VTAIL.n619 VTAIL.n618 12.0247
R384 VTAIL.n628 VTAIL.n586 12.0247
R385 VTAIL.n45 VTAIL.n44 12.0247
R386 VTAIL.n54 VTAIL.n12 12.0247
R387 VTAIL.n127 VTAIL.n126 12.0247
R388 VTAIL.n136 VTAIL.n94 12.0247
R389 VTAIL.n209 VTAIL.n208 12.0247
R390 VTAIL.n218 VTAIL.n176 12.0247
R391 VTAIL.n546 VTAIL.n504 12.0247
R392 VTAIL.n537 VTAIL.n536 12.0247
R393 VTAIL.n464 VTAIL.n422 12.0247
R394 VTAIL.n455 VTAIL.n454 12.0247
R395 VTAIL.n382 VTAIL.n340 12.0247
R396 VTAIL.n373 VTAIL.n372 12.0247
R397 VTAIL.n300 VTAIL.n258 12.0247
R398 VTAIL.n291 VTAIL.n290 12.0247
R399 VTAIL.n614 VTAIL.n592 11.249
R400 VTAIL.n632 VTAIL.n631 11.249
R401 VTAIL.n40 VTAIL.n18 11.249
R402 VTAIL.n58 VTAIL.n57 11.249
R403 VTAIL.n122 VTAIL.n100 11.249
R404 VTAIL.n140 VTAIL.n139 11.249
R405 VTAIL.n204 VTAIL.n182 11.249
R406 VTAIL.n222 VTAIL.n221 11.249
R407 VTAIL.n550 VTAIL.n549 11.249
R408 VTAIL.n533 VTAIL.n510 11.249
R409 VTAIL.n468 VTAIL.n467 11.249
R410 VTAIL.n451 VTAIL.n428 11.249
R411 VTAIL.n386 VTAIL.n385 11.249
R412 VTAIL.n369 VTAIL.n346 11.249
R413 VTAIL.n304 VTAIL.n303 11.249
R414 VTAIL.n287 VTAIL.n264 11.249
R415 VTAIL.n601 VTAIL.n599 10.7239
R416 VTAIL.n27 VTAIL.n25 10.7239
R417 VTAIL.n109 VTAIL.n107 10.7239
R418 VTAIL.n191 VTAIL.n189 10.7239
R419 VTAIL.n520 VTAIL.n518 10.7239
R420 VTAIL.n438 VTAIL.n436 10.7239
R421 VTAIL.n356 VTAIL.n354 10.7239
R422 VTAIL.n274 VTAIL.n272 10.7239
R423 VTAIL.n613 VTAIL.n594 10.4732
R424 VTAIL.n635 VTAIL.n584 10.4732
R425 VTAIL.n39 VTAIL.n20 10.4732
R426 VTAIL.n61 VTAIL.n10 10.4732
R427 VTAIL.n121 VTAIL.n102 10.4732
R428 VTAIL.n143 VTAIL.n92 10.4732
R429 VTAIL.n203 VTAIL.n184 10.4732
R430 VTAIL.n225 VTAIL.n174 10.4732
R431 VTAIL.n553 VTAIL.n502 10.4732
R432 VTAIL.n532 VTAIL.n513 10.4732
R433 VTAIL.n471 VTAIL.n420 10.4732
R434 VTAIL.n450 VTAIL.n431 10.4732
R435 VTAIL.n389 VTAIL.n338 10.4732
R436 VTAIL.n368 VTAIL.n349 10.4732
R437 VTAIL.n307 VTAIL.n256 10.4732
R438 VTAIL.n286 VTAIL.n267 10.4732
R439 VTAIL.n610 VTAIL.n609 9.69747
R440 VTAIL.n636 VTAIL.n582 9.69747
R441 VTAIL.n36 VTAIL.n35 9.69747
R442 VTAIL.n62 VTAIL.n8 9.69747
R443 VTAIL.n118 VTAIL.n117 9.69747
R444 VTAIL.n144 VTAIL.n90 9.69747
R445 VTAIL.n200 VTAIL.n199 9.69747
R446 VTAIL.n226 VTAIL.n172 9.69747
R447 VTAIL.n554 VTAIL.n500 9.69747
R448 VTAIL.n529 VTAIL.n528 9.69747
R449 VTAIL.n472 VTAIL.n418 9.69747
R450 VTAIL.n447 VTAIL.n446 9.69747
R451 VTAIL.n390 VTAIL.n336 9.69747
R452 VTAIL.n365 VTAIL.n364 9.69747
R453 VTAIL.n308 VTAIL.n254 9.69747
R454 VTAIL.n283 VTAIL.n282 9.69747
R455 VTAIL.n654 VTAIL.n653 9.45567
R456 VTAIL.n80 VTAIL.n79 9.45567
R457 VTAIL.n162 VTAIL.n161 9.45567
R458 VTAIL.n244 VTAIL.n243 9.45567
R459 VTAIL.n572 VTAIL.n571 9.45567
R460 VTAIL.n490 VTAIL.n489 9.45567
R461 VTAIL.n408 VTAIL.n407 9.45567
R462 VTAIL.n326 VTAIL.n325 9.45567
R463 VTAIL.n647 VTAIL.n646 9.3005
R464 VTAIL.n576 VTAIL.n575 9.3005
R465 VTAIL.n653 VTAIL.n652 9.3005
R466 VTAIL.n580 VTAIL.n579 9.3005
R467 VTAIL.n639 VTAIL.n638 9.3005
R468 VTAIL.n637 VTAIL.n636 9.3005
R469 VTAIL.n584 VTAIL.n583 9.3005
R470 VTAIL.n631 VTAIL.n630 9.3005
R471 VTAIL.n629 VTAIL.n628 9.3005
R472 VTAIL.n588 VTAIL.n587 9.3005
R473 VTAIL.n603 VTAIL.n602 9.3005
R474 VTAIL.n605 VTAIL.n604 9.3005
R475 VTAIL.n596 VTAIL.n595 9.3005
R476 VTAIL.n611 VTAIL.n610 9.3005
R477 VTAIL.n613 VTAIL.n612 9.3005
R478 VTAIL.n592 VTAIL.n591 9.3005
R479 VTAIL.n620 VTAIL.n619 9.3005
R480 VTAIL.n622 VTAIL.n621 9.3005
R481 VTAIL.n645 VTAIL.n644 9.3005
R482 VTAIL.n73 VTAIL.n72 9.3005
R483 VTAIL.n2 VTAIL.n1 9.3005
R484 VTAIL.n79 VTAIL.n78 9.3005
R485 VTAIL.n6 VTAIL.n5 9.3005
R486 VTAIL.n65 VTAIL.n64 9.3005
R487 VTAIL.n63 VTAIL.n62 9.3005
R488 VTAIL.n10 VTAIL.n9 9.3005
R489 VTAIL.n57 VTAIL.n56 9.3005
R490 VTAIL.n55 VTAIL.n54 9.3005
R491 VTAIL.n14 VTAIL.n13 9.3005
R492 VTAIL.n29 VTAIL.n28 9.3005
R493 VTAIL.n31 VTAIL.n30 9.3005
R494 VTAIL.n22 VTAIL.n21 9.3005
R495 VTAIL.n37 VTAIL.n36 9.3005
R496 VTAIL.n39 VTAIL.n38 9.3005
R497 VTAIL.n18 VTAIL.n17 9.3005
R498 VTAIL.n46 VTAIL.n45 9.3005
R499 VTAIL.n48 VTAIL.n47 9.3005
R500 VTAIL.n71 VTAIL.n70 9.3005
R501 VTAIL.n155 VTAIL.n154 9.3005
R502 VTAIL.n84 VTAIL.n83 9.3005
R503 VTAIL.n161 VTAIL.n160 9.3005
R504 VTAIL.n88 VTAIL.n87 9.3005
R505 VTAIL.n147 VTAIL.n146 9.3005
R506 VTAIL.n145 VTAIL.n144 9.3005
R507 VTAIL.n92 VTAIL.n91 9.3005
R508 VTAIL.n139 VTAIL.n138 9.3005
R509 VTAIL.n137 VTAIL.n136 9.3005
R510 VTAIL.n96 VTAIL.n95 9.3005
R511 VTAIL.n111 VTAIL.n110 9.3005
R512 VTAIL.n113 VTAIL.n112 9.3005
R513 VTAIL.n104 VTAIL.n103 9.3005
R514 VTAIL.n119 VTAIL.n118 9.3005
R515 VTAIL.n121 VTAIL.n120 9.3005
R516 VTAIL.n100 VTAIL.n99 9.3005
R517 VTAIL.n128 VTAIL.n127 9.3005
R518 VTAIL.n130 VTAIL.n129 9.3005
R519 VTAIL.n153 VTAIL.n152 9.3005
R520 VTAIL.n237 VTAIL.n236 9.3005
R521 VTAIL.n166 VTAIL.n165 9.3005
R522 VTAIL.n243 VTAIL.n242 9.3005
R523 VTAIL.n170 VTAIL.n169 9.3005
R524 VTAIL.n229 VTAIL.n228 9.3005
R525 VTAIL.n227 VTAIL.n226 9.3005
R526 VTAIL.n174 VTAIL.n173 9.3005
R527 VTAIL.n221 VTAIL.n220 9.3005
R528 VTAIL.n219 VTAIL.n218 9.3005
R529 VTAIL.n178 VTAIL.n177 9.3005
R530 VTAIL.n193 VTAIL.n192 9.3005
R531 VTAIL.n195 VTAIL.n194 9.3005
R532 VTAIL.n186 VTAIL.n185 9.3005
R533 VTAIL.n201 VTAIL.n200 9.3005
R534 VTAIL.n203 VTAIL.n202 9.3005
R535 VTAIL.n182 VTAIL.n181 9.3005
R536 VTAIL.n210 VTAIL.n209 9.3005
R537 VTAIL.n212 VTAIL.n211 9.3005
R538 VTAIL.n235 VTAIL.n234 9.3005
R539 VTAIL.n494 VTAIL.n493 9.3005
R540 VTAIL.n565 VTAIL.n564 9.3005
R541 VTAIL.n563 VTAIL.n562 9.3005
R542 VTAIL.n498 VTAIL.n497 9.3005
R543 VTAIL.n557 VTAIL.n556 9.3005
R544 VTAIL.n555 VTAIL.n554 9.3005
R545 VTAIL.n502 VTAIL.n501 9.3005
R546 VTAIL.n549 VTAIL.n548 9.3005
R547 VTAIL.n547 VTAIL.n546 9.3005
R548 VTAIL.n506 VTAIL.n505 9.3005
R549 VTAIL.n540 VTAIL.n539 9.3005
R550 VTAIL.n538 VTAIL.n537 9.3005
R551 VTAIL.n510 VTAIL.n509 9.3005
R552 VTAIL.n532 VTAIL.n531 9.3005
R553 VTAIL.n530 VTAIL.n529 9.3005
R554 VTAIL.n515 VTAIL.n514 9.3005
R555 VTAIL.n524 VTAIL.n523 9.3005
R556 VTAIL.n522 VTAIL.n521 9.3005
R557 VTAIL.n571 VTAIL.n570 9.3005
R558 VTAIL.n440 VTAIL.n439 9.3005
R559 VTAIL.n442 VTAIL.n441 9.3005
R560 VTAIL.n433 VTAIL.n432 9.3005
R561 VTAIL.n448 VTAIL.n447 9.3005
R562 VTAIL.n450 VTAIL.n449 9.3005
R563 VTAIL.n428 VTAIL.n427 9.3005
R564 VTAIL.n456 VTAIL.n455 9.3005
R565 VTAIL.n458 VTAIL.n457 9.3005
R566 VTAIL.n412 VTAIL.n411 9.3005
R567 VTAIL.n489 VTAIL.n488 9.3005
R568 VTAIL.n483 VTAIL.n482 9.3005
R569 VTAIL.n481 VTAIL.n480 9.3005
R570 VTAIL.n416 VTAIL.n415 9.3005
R571 VTAIL.n475 VTAIL.n474 9.3005
R572 VTAIL.n473 VTAIL.n472 9.3005
R573 VTAIL.n420 VTAIL.n419 9.3005
R574 VTAIL.n467 VTAIL.n466 9.3005
R575 VTAIL.n465 VTAIL.n464 9.3005
R576 VTAIL.n424 VTAIL.n423 9.3005
R577 VTAIL.n358 VTAIL.n357 9.3005
R578 VTAIL.n360 VTAIL.n359 9.3005
R579 VTAIL.n351 VTAIL.n350 9.3005
R580 VTAIL.n366 VTAIL.n365 9.3005
R581 VTAIL.n368 VTAIL.n367 9.3005
R582 VTAIL.n346 VTAIL.n345 9.3005
R583 VTAIL.n374 VTAIL.n373 9.3005
R584 VTAIL.n376 VTAIL.n375 9.3005
R585 VTAIL.n330 VTAIL.n329 9.3005
R586 VTAIL.n407 VTAIL.n406 9.3005
R587 VTAIL.n401 VTAIL.n400 9.3005
R588 VTAIL.n399 VTAIL.n398 9.3005
R589 VTAIL.n334 VTAIL.n333 9.3005
R590 VTAIL.n393 VTAIL.n392 9.3005
R591 VTAIL.n391 VTAIL.n390 9.3005
R592 VTAIL.n338 VTAIL.n337 9.3005
R593 VTAIL.n385 VTAIL.n384 9.3005
R594 VTAIL.n383 VTAIL.n382 9.3005
R595 VTAIL.n342 VTAIL.n341 9.3005
R596 VTAIL.n276 VTAIL.n275 9.3005
R597 VTAIL.n278 VTAIL.n277 9.3005
R598 VTAIL.n269 VTAIL.n268 9.3005
R599 VTAIL.n284 VTAIL.n283 9.3005
R600 VTAIL.n286 VTAIL.n285 9.3005
R601 VTAIL.n264 VTAIL.n263 9.3005
R602 VTAIL.n292 VTAIL.n291 9.3005
R603 VTAIL.n294 VTAIL.n293 9.3005
R604 VTAIL.n248 VTAIL.n247 9.3005
R605 VTAIL.n325 VTAIL.n324 9.3005
R606 VTAIL.n319 VTAIL.n318 9.3005
R607 VTAIL.n317 VTAIL.n316 9.3005
R608 VTAIL.n252 VTAIL.n251 9.3005
R609 VTAIL.n311 VTAIL.n310 9.3005
R610 VTAIL.n309 VTAIL.n308 9.3005
R611 VTAIL.n256 VTAIL.n255 9.3005
R612 VTAIL.n303 VTAIL.n302 9.3005
R613 VTAIL.n301 VTAIL.n300 9.3005
R614 VTAIL.n260 VTAIL.n259 9.3005
R615 VTAIL.n606 VTAIL.n596 8.92171
R616 VTAIL.n640 VTAIL.n639 8.92171
R617 VTAIL.n654 VTAIL.n574 8.92171
R618 VTAIL.n32 VTAIL.n22 8.92171
R619 VTAIL.n66 VTAIL.n65 8.92171
R620 VTAIL.n80 VTAIL.n0 8.92171
R621 VTAIL.n114 VTAIL.n104 8.92171
R622 VTAIL.n148 VTAIL.n147 8.92171
R623 VTAIL.n162 VTAIL.n82 8.92171
R624 VTAIL.n196 VTAIL.n186 8.92171
R625 VTAIL.n230 VTAIL.n229 8.92171
R626 VTAIL.n244 VTAIL.n164 8.92171
R627 VTAIL.n572 VTAIL.n492 8.92171
R628 VTAIL.n558 VTAIL.n557 8.92171
R629 VTAIL.n525 VTAIL.n515 8.92171
R630 VTAIL.n490 VTAIL.n410 8.92171
R631 VTAIL.n476 VTAIL.n475 8.92171
R632 VTAIL.n443 VTAIL.n433 8.92171
R633 VTAIL.n408 VTAIL.n328 8.92171
R634 VTAIL.n394 VTAIL.n393 8.92171
R635 VTAIL.n361 VTAIL.n351 8.92171
R636 VTAIL.n326 VTAIL.n246 8.92171
R637 VTAIL.n312 VTAIL.n311 8.92171
R638 VTAIL.n279 VTAIL.n269 8.92171
R639 VTAIL.n605 VTAIL.n598 8.14595
R640 VTAIL.n643 VTAIL.n580 8.14595
R641 VTAIL.n652 VTAIL.n651 8.14595
R642 VTAIL.n31 VTAIL.n24 8.14595
R643 VTAIL.n69 VTAIL.n6 8.14595
R644 VTAIL.n78 VTAIL.n77 8.14595
R645 VTAIL.n113 VTAIL.n106 8.14595
R646 VTAIL.n151 VTAIL.n88 8.14595
R647 VTAIL.n160 VTAIL.n159 8.14595
R648 VTAIL.n195 VTAIL.n188 8.14595
R649 VTAIL.n233 VTAIL.n170 8.14595
R650 VTAIL.n242 VTAIL.n241 8.14595
R651 VTAIL.n570 VTAIL.n569 8.14595
R652 VTAIL.n561 VTAIL.n498 8.14595
R653 VTAIL.n524 VTAIL.n517 8.14595
R654 VTAIL.n488 VTAIL.n487 8.14595
R655 VTAIL.n479 VTAIL.n416 8.14595
R656 VTAIL.n442 VTAIL.n435 8.14595
R657 VTAIL.n406 VTAIL.n405 8.14595
R658 VTAIL.n397 VTAIL.n334 8.14595
R659 VTAIL.n360 VTAIL.n353 8.14595
R660 VTAIL.n324 VTAIL.n323 8.14595
R661 VTAIL.n315 VTAIL.n252 8.14595
R662 VTAIL.n278 VTAIL.n271 8.14595
R663 VTAIL.n602 VTAIL.n601 7.3702
R664 VTAIL.n644 VTAIL.n578 7.3702
R665 VTAIL.n648 VTAIL.n576 7.3702
R666 VTAIL.n28 VTAIL.n27 7.3702
R667 VTAIL.n70 VTAIL.n4 7.3702
R668 VTAIL.n74 VTAIL.n2 7.3702
R669 VTAIL.n110 VTAIL.n109 7.3702
R670 VTAIL.n152 VTAIL.n86 7.3702
R671 VTAIL.n156 VTAIL.n84 7.3702
R672 VTAIL.n192 VTAIL.n191 7.3702
R673 VTAIL.n234 VTAIL.n168 7.3702
R674 VTAIL.n238 VTAIL.n166 7.3702
R675 VTAIL.n566 VTAIL.n494 7.3702
R676 VTAIL.n562 VTAIL.n496 7.3702
R677 VTAIL.n521 VTAIL.n520 7.3702
R678 VTAIL.n484 VTAIL.n412 7.3702
R679 VTAIL.n480 VTAIL.n414 7.3702
R680 VTAIL.n439 VTAIL.n438 7.3702
R681 VTAIL.n402 VTAIL.n330 7.3702
R682 VTAIL.n398 VTAIL.n332 7.3702
R683 VTAIL.n357 VTAIL.n356 7.3702
R684 VTAIL.n320 VTAIL.n248 7.3702
R685 VTAIL.n316 VTAIL.n250 7.3702
R686 VTAIL.n275 VTAIL.n274 7.3702
R687 VTAIL.n647 VTAIL.n578 6.59444
R688 VTAIL.n648 VTAIL.n647 6.59444
R689 VTAIL.n73 VTAIL.n4 6.59444
R690 VTAIL.n74 VTAIL.n73 6.59444
R691 VTAIL.n155 VTAIL.n86 6.59444
R692 VTAIL.n156 VTAIL.n155 6.59444
R693 VTAIL.n237 VTAIL.n168 6.59444
R694 VTAIL.n238 VTAIL.n237 6.59444
R695 VTAIL.n566 VTAIL.n565 6.59444
R696 VTAIL.n565 VTAIL.n496 6.59444
R697 VTAIL.n484 VTAIL.n483 6.59444
R698 VTAIL.n483 VTAIL.n414 6.59444
R699 VTAIL.n402 VTAIL.n401 6.59444
R700 VTAIL.n401 VTAIL.n332 6.59444
R701 VTAIL.n320 VTAIL.n319 6.59444
R702 VTAIL.n319 VTAIL.n250 6.59444
R703 VTAIL.n602 VTAIL.n598 5.81868
R704 VTAIL.n644 VTAIL.n643 5.81868
R705 VTAIL.n651 VTAIL.n576 5.81868
R706 VTAIL.n28 VTAIL.n24 5.81868
R707 VTAIL.n70 VTAIL.n69 5.81868
R708 VTAIL.n77 VTAIL.n2 5.81868
R709 VTAIL.n110 VTAIL.n106 5.81868
R710 VTAIL.n152 VTAIL.n151 5.81868
R711 VTAIL.n159 VTAIL.n84 5.81868
R712 VTAIL.n192 VTAIL.n188 5.81868
R713 VTAIL.n234 VTAIL.n233 5.81868
R714 VTAIL.n241 VTAIL.n166 5.81868
R715 VTAIL.n569 VTAIL.n494 5.81868
R716 VTAIL.n562 VTAIL.n561 5.81868
R717 VTAIL.n521 VTAIL.n517 5.81868
R718 VTAIL.n487 VTAIL.n412 5.81868
R719 VTAIL.n480 VTAIL.n479 5.81868
R720 VTAIL.n439 VTAIL.n435 5.81868
R721 VTAIL.n405 VTAIL.n330 5.81868
R722 VTAIL.n398 VTAIL.n397 5.81868
R723 VTAIL.n357 VTAIL.n353 5.81868
R724 VTAIL.n323 VTAIL.n248 5.81868
R725 VTAIL.n316 VTAIL.n315 5.81868
R726 VTAIL.n275 VTAIL.n271 5.81868
R727 VTAIL.n606 VTAIL.n605 5.04292
R728 VTAIL.n640 VTAIL.n580 5.04292
R729 VTAIL.n652 VTAIL.n574 5.04292
R730 VTAIL.n32 VTAIL.n31 5.04292
R731 VTAIL.n66 VTAIL.n6 5.04292
R732 VTAIL.n78 VTAIL.n0 5.04292
R733 VTAIL.n114 VTAIL.n113 5.04292
R734 VTAIL.n148 VTAIL.n88 5.04292
R735 VTAIL.n160 VTAIL.n82 5.04292
R736 VTAIL.n196 VTAIL.n195 5.04292
R737 VTAIL.n230 VTAIL.n170 5.04292
R738 VTAIL.n242 VTAIL.n164 5.04292
R739 VTAIL.n570 VTAIL.n492 5.04292
R740 VTAIL.n558 VTAIL.n498 5.04292
R741 VTAIL.n525 VTAIL.n524 5.04292
R742 VTAIL.n488 VTAIL.n410 5.04292
R743 VTAIL.n476 VTAIL.n416 5.04292
R744 VTAIL.n443 VTAIL.n442 5.04292
R745 VTAIL.n406 VTAIL.n328 5.04292
R746 VTAIL.n394 VTAIL.n334 5.04292
R747 VTAIL.n361 VTAIL.n360 5.04292
R748 VTAIL.n324 VTAIL.n246 5.04292
R749 VTAIL.n312 VTAIL.n252 5.04292
R750 VTAIL.n279 VTAIL.n278 5.04292
R751 VTAIL.n609 VTAIL.n596 4.26717
R752 VTAIL.n639 VTAIL.n582 4.26717
R753 VTAIL.n35 VTAIL.n22 4.26717
R754 VTAIL.n65 VTAIL.n8 4.26717
R755 VTAIL.n117 VTAIL.n104 4.26717
R756 VTAIL.n147 VTAIL.n90 4.26717
R757 VTAIL.n199 VTAIL.n186 4.26717
R758 VTAIL.n229 VTAIL.n172 4.26717
R759 VTAIL.n557 VTAIL.n500 4.26717
R760 VTAIL.n528 VTAIL.n515 4.26717
R761 VTAIL.n475 VTAIL.n418 4.26717
R762 VTAIL.n446 VTAIL.n433 4.26717
R763 VTAIL.n393 VTAIL.n336 4.26717
R764 VTAIL.n364 VTAIL.n351 4.26717
R765 VTAIL.n311 VTAIL.n254 4.26717
R766 VTAIL.n282 VTAIL.n269 4.26717
R767 VTAIL.n610 VTAIL.n594 3.49141
R768 VTAIL.n636 VTAIL.n635 3.49141
R769 VTAIL.n36 VTAIL.n20 3.49141
R770 VTAIL.n62 VTAIL.n61 3.49141
R771 VTAIL.n118 VTAIL.n102 3.49141
R772 VTAIL.n144 VTAIL.n143 3.49141
R773 VTAIL.n200 VTAIL.n184 3.49141
R774 VTAIL.n226 VTAIL.n225 3.49141
R775 VTAIL.n554 VTAIL.n553 3.49141
R776 VTAIL.n529 VTAIL.n513 3.49141
R777 VTAIL.n472 VTAIL.n471 3.49141
R778 VTAIL.n447 VTAIL.n431 3.49141
R779 VTAIL.n390 VTAIL.n389 3.49141
R780 VTAIL.n365 VTAIL.n349 3.49141
R781 VTAIL.n308 VTAIL.n307 3.49141
R782 VTAIL.n283 VTAIL.n267 3.49141
R783 VTAIL.n614 VTAIL.n613 2.71565
R784 VTAIL.n632 VTAIL.n584 2.71565
R785 VTAIL.n40 VTAIL.n39 2.71565
R786 VTAIL.n58 VTAIL.n10 2.71565
R787 VTAIL.n122 VTAIL.n121 2.71565
R788 VTAIL.n140 VTAIL.n92 2.71565
R789 VTAIL.n204 VTAIL.n203 2.71565
R790 VTAIL.n222 VTAIL.n174 2.71565
R791 VTAIL.n550 VTAIL.n502 2.71565
R792 VTAIL.n533 VTAIL.n532 2.71565
R793 VTAIL.n468 VTAIL.n420 2.71565
R794 VTAIL.n451 VTAIL.n450 2.71565
R795 VTAIL.n386 VTAIL.n338 2.71565
R796 VTAIL.n369 VTAIL.n368 2.71565
R797 VTAIL.n304 VTAIL.n256 2.71565
R798 VTAIL.n287 VTAIL.n286 2.71565
R799 VTAIL.n409 VTAIL.n327 2.44878
R800 VTAIL.n573 VTAIL.n491 2.44878
R801 VTAIL.n245 VTAIL.n163 2.44878
R802 VTAIL.n522 VTAIL.n518 2.41282
R803 VTAIL.n440 VTAIL.n436 2.41282
R804 VTAIL.n358 VTAIL.n354 2.41282
R805 VTAIL.n276 VTAIL.n272 2.41282
R806 VTAIL.n603 VTAIL.n599 2.41282
R807 VTAIL.n29 VTAIL.n25 2.41282
R808 VTAIL.n111 VTAIL.n107 2.41282
R809 VTAIL.n193 VTAIL.n189 2.41282
R810 VTAIL.n618 VTAIL.n592 1.93989
R811 VTAIL.n631 VTAIL.n586 1.93989
R812 VTAIL.n44 VTAIL.n18 1.93989
R813 VTAIL.n57 VTAIL.n12 1.93989
R814 VTAIL.n126 VTAIL.n100 1.93989
R815 VTAIL.n139 VTAIL.n94 1.93989
R816 VTAIL.n208 VTAIL.n182 1.93989
R817 VTAIL.n221 VTAIL.n176 1.93989
R818 VTAIL.n549 VTAIL.n504 1.93989
R819 VTAIL.n536 VTAIL.n510 1.93989
R820 VTAIL.n467 VTAIL.n422 1.93989
R821 VTAIL.n454 VTAIL.n428 1.93989
R822 VTAIL.n385 VTAIL.n340 1.93989
R823 VTAIL.n372 VTAIL.n346 1.93989
R824 VTAIL.n303 VTAIL.n258 1.93989
R825 VTAIL.n290 VTAIL.n264 1.93989
R826 VTAIL VTAIL.n81 1.28283
R827 VTAIL VTAIL.n655 1.16645
R828 VTAIL.n619 VTAIL.n590 1.16414
R829 VTAIL.n628 VTAIL.n627 1.16414
R830 VTAIL.n45 VTAIL.n16 1.16414
R831 VTAIL.n54 VTAIL.n53 1.16414
R832 VTAIL.n127 VTAIL.n98 1.16414
R833 VTAIL.n136 VTAIL.n135 1.16414
R834 VTAIL.n209 VTAIL.n180 1.16414
R835 VTAIL.n218 VTAIL.n217 1.16414
R836 VTAIL.n546 VTAIL.n545 1.16414
R837 VTAIL.n537 VTAIL.n508 1.16414
R838 VTAIL.n464 VTAIL.n463 1.16414
R839 VTAIL.n455 VTAIL.n426 1.16414
R840 VTAIL.n382 VTAIL.n381 1.16414
R841 VTAIL.n373 VTAIL.n344 1.16414
R842 VTAIL.n300 VTAIL.n299 1.16414
R843 VTAIL.n291 VTAIL.n262 1.16414
R844 VTAIL.n491 VTAIL.n409 0.470328
R845 VTAIL.n163 VTAIL.n81 0.470328
R846 VTAIL.n623 VTAIL.n622 0.388379
R847 VTAIL.n624 VTAIL.n588 0.388379
R848 VTAIL.n49 VTAIL.n48 0.388379
R849 VTAIL.n50 VTAIL.n14 0.388379
R850 VTAIL.n131 VTAIL.n130 0.388379
R851 VTAIL.n132 VTAIL.n96 0.388379
R852 VTAIL.n213 VTAIL.n212 0.388379
R853 VTAIL.n214 VTAIL.n178 0.388379
R854 VTAIL.n542 VTAIL.n506 0.388379
R855 VTAIL.n541 VTAIL.n540 0.388379
R856 VTAIL.n460 VTAIL.n424 0.388379
R857 VTAIL.n459 VTAIL.n458 0.388379
R858 VTAIL.n378 VTAIL.n342 0.388379
R859 VTAIL.n377 VTAIL.n376 0.388379
R860 VTAIL.n296 VTAIL.n260 0.388379
R861 VTAIL.n295 VTAIL.n294 0.388379
R862 VTAIL.n604 VTAIL.n603 0.155672
R863 VTAIL.n604 VTAIL.n595 0.155672
R864 VTAIL.n611 VTAIL.n595 0.155672
R865 VTAIL.n612 VTAIL.n611 0.155672
R866 VTAIL.n612 VTAIL.n591 0.155672
R867 VTAIL.n620 VTAIL.n591 0.155672
R868 VTAIL.n621 VTAIL.n620 0.155672
R869 VTAIL.n621 VTAIL.n587 0.155672
R870 VTAIL.n629 VTAIL.n587 0.155672
R871 VTAIL.n630 VTAIL.n629 0.155672
R872 VTAIL.n630 VTAIL.n583 0.155672
R873 VTAIL.n637 VTAIL.n583 0.155672
R874 VTAIL.n638 VTAIL.n637 0.155672
R875 VTAIL.n638 VTAIL.n579 0.155672
R876 VTAIL.n645 VTAIL.n579 0.155672
R877 VTAIL.n646 VTAIL.n645 0.155672
R878 VTAIL.n646 VTAIL.n575 0.155672
R879 VTAIL.n653 VTAIL.n575 0.155672
R880 VTAIL.n30 VTAIL.n29 0.155672
R881 VTAIL.n30 VTAIL.n21 0.155672
R882 VTAIL.n37 VTAIL.n21 0.155672
R883 VTAIL.n38 VTAIL.n37 0.155672
R884 VTAIL.n38 VTAIL.n17 0.155672
R885 VTAIL.n46 VTAIL.n17 0.155672
R886 VTAIL.n47 VTAIL.n46 0.155672
R887 VTAIL.n47 VTAIL.n13 0.155672
R888 VTAIL.n55 VTAIL.n13 0.155672
R889 VTAIL.n56 VTAIL.n55 0.155672
R890 VTAIL.n56 VTAIL.n9 0.155672
R891 VTAIL.n63 VTAIL.n9 0.155672
R892 VTAIL.n64 VTAIL.n63 0.155672
R893 VTAIL.n64 VTAIL.n5 0.155672
R894 VTAIL.n71 VTAIL.n5 0.155672
R895 VTAIL.n72 VTAIL.n71 0.155672
R896 VTAIL.n72 VTAIL.n1 0.155672
R897 VTAIL.n79 VTAIL.n1 0.155672
R898 VTAIL.n112 VTAIL.n111 0.155672
R899 VTAIL.n112 VTAIL.n103 0.155672
R900 VTAIL.n119 VTAIL.n103 0.155672
R901 VTAIL.n120 VTAIL.n119 0.155672
R902 VTAIL.n120 VTAIL.n99 0.155672
R903 VTAIL.n128 VTAIL.n99 0.155672
R904 VTAIL.n129 VTAIL.n128 0.155672
R905 VTAIL.n129 VTAIL.n95 0.155672
R906 VTAIL.n137 VTAIL.n95 0.155672
R907 VTAIL.n138 VTAIL.n137 0.155672
R908 VTAIL.n138 VTAIL.n91 0.155672
R909 VTAIL.n145 VTAIL.n91 0.155672
R910 VTAIL.n146 VTAIL.n145 0.155672
R911 VTAIL.n146 VTAIL.n87 0.155672
R912 VTAIL.n153 VTAIL.n87 0.155672
R913 VTAIL.n154 VTAIL.n153 0.155672
R914 VTAIL.n154 VTAIL.n83 0.155672
R915 VTAIL.n161 VTAIL.n83 0.155672
R916 VTAIL.n194 VTAIL.n193 0.155672
R917 VTAIL.n194 VTAIL.n185 0.155672
R918 VTAIL.n201 VTAIL.n185 0.155672
R919 VTAIL.n202 VTAIL.n201 0.155672
R920 VTAIL.n202 VTAIL.n181 0.155672
R921 VTAIL.n210 VTAIL.n181 0.155672
R922 VTAIL.n211 VTAIL.n210 0.155672
R923 VTAIL.n211 VTAIL.n177 0.155672
R924 VTAIL.n219 VTAIL.n177 0.155672
R925 VTAIL.n220 VTAIL.n219 0.155672
R926 VTAIL.n220 VTAIL.n173 0.155672
R927 VTAIL.n227 VTAIL.n173 0.155672
R928 VTAIL.n228 VTAIL.n227 0.155672
R929 VTAIL.n228 VTAIL.n169 0.155672
R930 VTAIL.n235 VTAIL.n169 0.155672
R931 VTAIL.n236 VTAIL.n235 0.155672
R932 VTAIL.n236 VTAIL.n165 0.155672
R933 VTAIL.n243 VTAIL.n165 0.155672
R934 VTAIL.n571 VTAIL.n493 0.155672
R935 VTAIL.n564 VTAIL.n493 0.155672
R936 VTAIL.n564 VTAIL.n563 0.155672
R937 VTAIL.n563 VTAIL.n497 0.155672
R938 VTAIL.n556 VTAIL.n497 0.155672
R939 VTAIL.n556 VTAIL.n555 0.155672
R940 VTAIL.n555 VTAIL.n501 0.155672
R941 VTAIL.n548 VTAIL.n501 0.155672
R942 VTAIL.n548 VTAIL.n547 0.155672
R943 VTAIL.n547 VTAIL.n505 0.155672
R944 VTAIL.n539 VTAIL.n505 0.155672
R945 VTAIL.n539 VTAIL.n538 0.155672
R946 VTAIL.n538 VTAIL.n509 0.155672
R947 VTAIL.n531 VTAIL.n509 0.155672
R948 VTAIL.n531 VTAIL.n530 0.155672
R949 VTAIL.n530 VTAIL.n514 0.155672
R950 VTAIL.n523 VTAIL.n514 0.155672
R951 VTAIL.n523 VTAIL.n522 0.155672
R952 VTAIL.n489 VTAIL.n411 0.155672
R953 VTAIL.n482 VTAIL.n411 0.155672
R954 VTAIL.n482 VTAIL.n481 0.155672
R955 VTAIL.n481 VTAIL.n415 0.155672
R956 VTAIL.n474 VTAIL.n415 0.155672
R957 VTAIL.n474 VTAIL.n473 0.155672
R958 VTAIL.n473 VTAIL.n419 0.155672
R959 VTAIL.n466 VTAIL.n419 0.155672
R960 VTAIL.n466 VTAIL.n465 0.155672
R961 VTAIL.n465 VTAIL.n423 0.155672
R962 VTAIL.n457 VTAIL.n423 0.155672
R963 VTAIL.n457 VTAIL.n456 0.155672
R964 VTAIL.n456 VTAIL.n427 0.155672
R965 VTAIL.n449 VTAIL.n427 0.155672
R966 VTAIL.n449 VTAIL.n448 0.155672
R967 VTAIL.n448 VTAIL.n432 0.155672
R968 VTAIL.n441 VTAIL.n432 0.155672
R969 VTAIL.n441 VTAIL.n440 0.155672
R970 VTAIL.n407 VTAIL.n329 0.155672
R971 VTAIL.n400 VTAIL.n329 0.155672
R972 VTAIL.n400 VTAIL.n399 0.155672
R973 VTAIL.n399 VTAIL.n333 0.155672
R974 VTAIL.n392 VTAIL.n333 0.155672
R975 VTAIL.n392 VTAIL.n391 0.155672
R976 VTAIL.n391 VTAIL.n337 0.155672
R977 VTAIL.n384 VTAIL.n337 0.155672
R978 VTAIL.n384 VTAIL.n383 0.155672
R979 VTAIL.n383 VTAIL.n341 0.155672
R980 VTAIL.n375 VTAIL.n341 0.155672
R981 VTAIL.n375 VTAIL.n374 0.155672
R982 VTAIL.n374 VTAIL.n345 0.155672
R983 VTAIL.n367 VTAIL.n345 0.155672
R984 VTAIL.n367 VTAIL.n366 0.155672
R985 VTAIL.n366 VTAIL.n350 0.155672
R986 VTAIL.n359 VTAIL.n350 0.155672
R987 VTAIL.n359 VTAIL.n358 0.155672
R988 VTAIL.n325 VTAIL.n247 0.155672
R989 VTAIL.n318 VTAIL.n247 0.155672
R990 VTAIL.n318 VTAIL.n317 0.155672
R991 VTAIL.n317 VTAIL.n251 0.155672
R992 VTAIL.n310 VTAIL.n251 0.155672
R993 VTAIL.n310 VTAIL.n309 0.155672
R994 VTAIL.n309 VTAIL.n255 0.155672
R995 VTAIL.n302 VTAIL.n255 0.155672
R996 VTAIL.n302 VTAIL.n301 0.155672
R997 VTAIL.n301 VTAIL.n259 0.155672
R998 VTAIL.n293 VTAIL.n259 0.155672
R999 VTAIL.n293 VTAIL.n292 0.155672
R1000 VTAIL.n292 VTAIL.n263 0.155672
R1001 VTAIL.n285 VTAIL.n263 0.155672
R1002 VTAIL.n285 VTAIL.n284 0.155672
R1003 VTAIL.n284 VTAIL.n268 0.155672
R1004 VTAIL.n277 VTAIL.n268 0.155672
R1005 VTAIL.n277 VTAIL.n276 0.155672
R1006 B.n503 B.n78 585
R1007 B.n505 B.n504 585
R1008 B.n506 B.n77 585
R1009 B.n508 B.n507 585
R1010 B.n509 B.n76 585
R1011 B.n511 B.n510 585
R1012 B.n512 B.n75 585
R1013 B.n514 B.n513 585
R1014 B.n515 B.n74 585
R1015 B.n517 B.n516 585
R1016 B.n518 B.n73 585
R1017 B.n520 B.n519 585
R1018 B.n521 B.n72 585
R1019 B.n523 B.n522 585
R1020 B.n524 B.n71 585
R1021 B.n526 B.n525 585
R1022 B.n527 B.n70 585
R1023 B.n529 B.n528 585
R1024 B.n530 B.n69 585
R1025 B.n532 B.n531 585
R1026 B.n533 B.n68 585
R1027 B.n535 B.n534 585
R1028 B.n536 B.n67 585
R1029 B.n538 B.n537 585
R1030 B.n539 B.n66 585
R1031 B.n541 B.n540 585
R1032 B.n542 B.n65 585
R1033 B.n544 B.n543 585
R1034 B.n545 B.n64 585
R1035 B.n547 B.n546 585
R1036 B.n548 B.n63 585
R1037 B.n550 B.n549 585
R1038 B.n551 B.n62 585
R1039 B.n553 B.n552 585
R1040 B.n554 B.n61 585
R1041 B.n556 B.n555 585
R1042 B.n557 B.n60 585
R1043 B.n559 B.n558 585
R1044 B.n560 B.n59 585
R1045 B.n562 B.n561 585
R1046 B.n563 B.n58 585
R1047 B.n565 B.n564 585
R1048 B.n566 B.n57 585
R1049 B.n568 B.n567 585
R1050 B.n569 B.n56 585
R1051 B.n571 B.n570 585
R1052 B.n572 B.n55 585
R1053 B.n574 B.n573 585
R1054 B.n575 B.n51 585
R1055 B.n577 B.n576 585
R1056 B.n578 B.n50 585
R1057 B.n580 B.n579 585
R1058 B.n581 B.n49 585
R1059 B.n583 B.n582 585
R1060 B.n584 B.n48 585
R1061 B.n586 B.n585 585
R1062 B.n587 B.n47 585
R1063 B.n589 B.n588 585
R1064 B.n590 B.n46 585
R1065 B.n592 B.n591 585
R1066 B.n594 B.n43 585
R1067 B.n596 B.n595 585
R1068 B.n597 B.n42 585
R1069 B.n599 B.n598 585
R1070 B.n600 B.n41 585
R1071 B.n602 B.n601 585
R1072 B.n603 B.n40 585
R1073 B.n605 B.n604 585
R1074 B.n606 B.n39 585
R1075 B.n608 B.n607 585
R1076 B.n609 B.n38 585
R1077 B.n611 B.n610 585
R1078 B.n612 B.n37 585
R1079 B.n614 B.n613 585
R1080 B.n615 B.n36 585
R1081 B.n617 B.n616 585
R1082 B.n618 B.n35 585
R1083 B.n620 B.n619 585
R1084 B.n621 B.n34 585
R1085 B.n623 B.n622 585
R1086 B.n624 B.n33 585
R1087 B.n626 B.n625 585
R1088 B.n627 B.n32 585
R1089 B.n629 B.n628 585
R1090 B.n630 B.n31 585
R1091 B.n632 B.n631 585
R1092 B.n633 B.n30 585
R1093 B.n635 B.n634 585
R1094 B.n636 B.n29 585
R1095 B.n638 B.n637 585
R1096 B.n639 B.n28 585
R1097 B.n641 B.n640 585
R1098 B.n642 B.n27 585
R1099 B.n644 B.n643 585
R1100 B.n645 B.n26 585
R1101 B.n647 B.n646 585
R1102 B.n648 B.n25 585
R1103 B.n650 B.n649 585
R1104 B.n651 B.n24 585
R1105 B.n653 B.n652 585
R1106 B.n654 B.n23 585
R1107 B.n656 B.n655 585
R1108 B.n657 B.n22 585
R1109 B.n659 B.n658 585
R1110 B.n660 B.n21 585
R1111 B.n662 B.n661 585
R1112 B.n663 B.n20 585
R1113 B.n665 B.n664 585
R1114 B.n666 B.n19 585
R1115 B.n668 B.n667 585
R1116 B.n502 B.n501 585
R1117 B.n500 B.n79 585
R1118 B.n499 B.n498 585
R1119 B.n497 B.n80 585
R1120 B.n496 B.n495 585
R1121 B.n494 B.n81 585
R1122 B.n493 B.n492 585
R1123 B.n491 B.n82 585
R1124 B.n490 B.n489 585
R1125 B.n488 B.n83 585
R1126 B.n487 B.n486 585
R1127 B.n485 B.n84 585
R1128 B.n484 B.n483 585
R1129 B.n482 B.n85 585
R1130 B.n481 B.n480 585
R1131 B.n479 B.n86 585
R1132 B.n478 B.n477 585
R1133 B.n476 B.n87 585
R1134 B.n475 B.n474 585
R1135 B.n473 B.n88 585
R1136 B.n472 B.n471 585
R1137 B.n470 B.n89 585
R1138 B.n469 B.n468 585
R1139 B.n467 B.n90 585
R1140 B.n466 B.n465 585
R1141 B.n464 B.n91 585
R1142 B.n463 B.n462 585
R1143 B.n461 B.n92 585
R1144 B.n460 B.n459 585
R1145 B.n458 B.n93 585
R1146 B.n457 B.n456 585
R1147 B.n455 B.n94 585
R1148 B.n454 B.n453 585
R1149 B.n452 B.n95 585
R1150 B.n451 B.n450 585
R1151 B.n449 B.n96 585
R1152 B.n448 B.n447 585
R1153 B.n446 B.n97 585
R1154 B.n445 B.n444 585
R1155 B.n443 B.n98 585
R1156 B.n442 B.n441 585
R1157 B.n440 B.n99 585
R1158 B.n439 B.n438 585
R1159 B.n437 B.n100 585
R1160 B.n436 B.n435 585
R1161 B.n434 B.n101 585
R1162 B.n433 B.n432 585
R1163 B.n431 B.n102 585
R1164 B.n430 B.n429 585
R1165 B.n428 B.n103 585
R1166 B.n427 B.n426 585
R1167 B.n425 B.n104 585
R1168 B.n424 B.n423 585
R1169 B.n422 B.n105 585
R1170 B.n421 B.n420 585
R1171 B.n419 B.n106 585
R1172 B.n418 B.n417 585
R1173 B.n416 B.n107 585
R1174 B.n415 B.n414 585
R1175 B.n413 B.n108 585
R1176 B.n412 B.n411 585
R1177 B.n410 B.n109 585
R1178 B.n409 B.n408 585
R1179 B.n407 B.n110 585
R1180 B.n406 B.n405 585
R1181 B.n404 B.n111 585
R1182 B.n403 B.n402 585
R1183 B.n236 B.n171 585
R1184 B.n238 B.n237 585
R1185 B.n239 B.n170 585
R1186 B.n241 B.n240 585
R1187 B.n242 B.n169 585
R1188 B.n244 B.n243 585
R1189 B.n245 B.n168 585
R1190 B.n247 B.n246 585
R1191 B.n248 B.n167 585
R1192 B.n250 B.n249 585
R1193 B.n251 B.n166 585
R1194 B.n253 B.n252 585
R1195 B.n254 B.n165 585
R1196 B.n256 B.n255 585
R1197 B.n257 B.n164 585
R1198 B.n259 B.n258 585
R1199 B.n260 B.n163 585
R1200 B.n262 B.n261 585
R1201 B.n263 B.n162 585
R1202 B.n265 B.n264 585
R1203 B.n266 B.n161 585
R1204 B.n268 B.n267 585
R1205 B.n269 B.n160 585
R1206 B.n271 B.n270 585
R1207 B.n272 B.n159 585
R1208 B.n274 B.n273 585
R1209 B.n275 B.n158 585
R1210 B.n277 B.n276 585
R1211 B.n278 B.n157 585
R1212 B.n280 B.n279 585
R1213 B.n281 B.n156 585
R1214 B.n283 B.n282 585
R1215 B.n284 B.n155 585
R1216 B.n286 B.n285 585
R1217 B.n287 B.n154 585
R1218 B.n289 B.n288 585
R1219 B.n290 B.n153 585
R1220 B.n292 B.n291 585
R1221 B.n293 B.n152 585
R1222 B.n295 B.n294 585
R1223 B.n296 B.n151 585
R1224 B.n298 B.n297 585
R1225 B.n299 B.n150 585
R1226 B.n301 B.n300 585
R1227 B.n302 B.n149 585
R1228 B.n304 B.n303 585
R1229 B.n305 B.n148 585
R1230 B.n307 B.n306 585
R1231 B.n308 B.n147 585
R1232 B.n310 B.n309 585
R1233 B.n312 B.n144 585
R1234 B.n314 B.n313 585
R1235 B.n315 B.n143 585
R1236 B.n317 B.n316 585
R1237 B.n318 B.n142 585
R1238 B.n320 B.n319 585
R1239 B.n321 B.n141 585
R1240 B.n323 B.n322 585
R1241 B.n324 B.n140 585
R1242 B.n326 B.n325 585
R1243 B.n328 B.n327 585
R1244 B.n329 B.n136 585
R1245 B.n331 B.n330 585
R1246 B.n332 B.n135 585
R1247 B.n334 B.n333 585
R1248 B.n335 B.n134 585
R1249 B.n337 B.n336 585
R1250 B.n338 B.n133 585
R1251 B.n340 B.n339 585
R1252 B.n341 B.n132 585
R1253 B.n343 B.n342 585
R1254 B.n344 B.n131 585
R1255 B.n346 B.n345 585
R1256 B.n347 B.n130 585
R1257 B.n349 B.n348 585
R1258 B.n350 B.n129 585
R1259 B.n352 B.n351 585
R1260 B.n353 B.n128 585
R1261 B.n355 B.n354 585
R1262 B.n356 B.n127 585
R1263 B.n358 B.n357 585
R1264 B.n359 B.n126 585
R1265 B.n361 B.n360 585
R1266 B.n362 B.n125 585
R1267 B.n364 B.n363 585
R1268 B.n365 B.n124 585
R1269 B.n367 B.n366 585
R1270 B.n368 B.n123 585
R1271 B.n370 B.n369 585
R1272 B.n371 B.n122 585
R1273 B.n373 B.n372 585
R1274 B.n374 B.n121 585
R1275 B.n376 B.n375 585
R1276 B.n377 B.n120 585
R1277 B.n379 B.n378 585
R1278 B.n380 B.n119 585
R1279 B.n382 B.n381 585
R1280 B.n383 B.n118 585
R1281 B.n385 B.n384 585
R1282 B.n386 B.n117 585
R1283 B.n388 B.n387 585
R1284 B.n389 B.n116 585
R1285 B.n391 B.n390 585
R1286 B.n392 B.n115 585
R1287 B.n394 B.n393 585
R1288 B.n395 B.n114 585
R1289 B.n397 B.n396 585
R1290 B.n398 B.n113 585
R1291 B.n400 B.n399 585
R1292 B.n401 B.n112 585
R1293 B.n235 B.n234 585
R1294 B.n233 B.n172 585
R1295 B.n232 B.n231 585
R1296 B.n230 B.n173 585
R1297 B.n229 B.n228 585
R1298 B.n227 B.n174 585
R1299 B.n226 B.n225 585
R1300 B.n224 B.n175 585
R1301 B.n223 B.n222 585
R1302 B.n221 B.n176 585
R1303 B.n220 B.n219 585
R1304 B.n218 B.n177 585
R1305 B.n217 B.n216 585
R1306 B.n215 B.n178 585
R1307 B.n214 B.n213 585
R1308 B.n212 B.n179 585
R1309 B.n211 B.n210 585
R1310 B.n209 B.n180 585
R1311 B.n208 B.n207 585
R1312 B.n206 B.n181 585
R1313 B.n205 B.n204 585
R1314 B.n203 B.n182 585
R1315 B.n202 B.n201 585
R1316 B.n200 B.n183 585
R1317 B.n199 B.n198 585
R1318 B.n197 B.n184 585
R1319 B.n196 B.n195 585
R1320 B.n194 B.n185 585
R1321 B.n193 B.n192 585
R1322 B.n191 B.n186 585
R1323 B.n190 B.n189 585
R1324 B.n188 B.n187 585
R1325 B.n2 B.n0 585
R1326 B.n717 B.n1 585
R1327 B.n716 B.n715 585
R1328 B.n714 B.n3 585
R1329 B.n713 B.n712 585
R1330 B.n711 B.n4 585
R1331 B.n710 B.n709 585
R1332 B.n708 B.n5 585
R1333 B.n707 B.n706 585
R1334 B.n705 B.n6 585
R1335 B.n704 B.n703 585
R1336 B.n702 B.n7 585
R1337 B.n701 B.n700 585
R1338 B.n699 B.n8 585
R1339 B.n698 B.n697 585
R1340 B.n696 B.n9 585
R1341 B.n695 B.n694 585
R1342 B.n693 B.n10 585
R1343 B.n692 B.n691 585
R1344 B.n690 B.n11 585
R1345 B.n689 B.n688 585
R1346 B.n687 B.n12 585
R1347 B.n686 B.n685 585
R1348 B.n684 B.n13 585
R1349 B.n683 B.n682 585
R1350 B.n681 B.n14 585
R1351 B.n680 B.n679 585
R1352 B.n678 B.n15 585
R1353 B.n677 B.n676 585
R1354 B.n675 B.n16 585
R1355 B.n674 B.n673 585
R1356 B.n672 B.n17 585
R1357 B.n671 B.n670 585
R1358 B.n669 B.n18 585
R1359 B.n719 B.n718 585
R1360 B.n236 B.n235 535.745
R1361 B.n669 B.n668 535.745
R1362 B.n403 B.n112 535.745
R1363 B.n501 B.n78 535.745
R1364 B.n137 B.t2 483.865
R1365 B.n52 B.t7 483.865
R1366 B.n145 B.t11 483.865
R1367 B.n44 B.t4 483.865
R1368 B.n138 B.t1 428.786
R1369 B.n53 B.t8 428.786
R1370 B.n146 B.t10 428.786
R1371 B.n45 B.t5 428.786
R1372 B.n137 B.t0 351.354
R1373 B.n145 B.t9 351.354
R1374 B.n44 B.t3 351.354
R1375 B.n52 B.t6 351.354
R1376 B.n235 B.n172 163.367
R1377 B.n231 B.n172 163.367
R1378 B.n231 B.n230 163.367
R1379 B.n230 B.n229 163.367
R1380 B.n229 B.n174 163.367
R1381 B.n225 B.n174 163.367
R1382 B.n225 B.n224 163.367
R1383 B.n224 B.n223 163.367
R1384 B.n223 B.n176 163.367
R1385 B.n219 B.n176 163.367
R1386 B.n219 B.n218 163.367
R1387 B.n218 B.n217 163.367
R1388 B.n217 B.n178 163.367
R1389 B.n213 B.n178 163.367
R1390 B.n213 B.n212 163.367
R1391 B.n212 B.n211 163.367
R1392 B.n211 B.n180 163.367
R1393 B.n207 B.n180 163.367
R1394 B.n207 B.n206 163.367
R1395 B.n206 B.n205 163.367
R1396 B.n205 B.n182 163.367
R1397 B.n201 B.n182 163.367
R1398 B.n201 B.n200 163.367
R1399 B.n200 B.n199 163.367
R1400 B.n199 B.n184 163.367
R1401 B.n195 B.n184 163.367
R1402 B.n195 B.n194 163.367
R1403 B.n194 B.n193 163.367
R1404 B.n193 B.n186 163.367
R1405 B.n189 B.n186 163.367
R1406 B.n189 B.n188 163.367
R1407 B.n188 B.n2 163.367
R1408 B.n718 B.n2 163.367
R1409 B.n718 B.n717 163.367
R1410 B.n717 B.n716 163.367
R1411 B.n716 B.n3 163.367
R1412 B.n712 B.n3 163.367
R1413 B.n712 B.n711 163.367
R1414 B.n711 B.n710 163.367
R1415 B.n710 B.n5 163.367
R1416 B.n706 B.n5 163.367
R1417 B.n706 B.n705 163.367
R1418 B.n705 B.n704 163.367
R1419 B.n704 B.n7 163.367
R1420 B.n700 B.n7 163.367
R1421 B.n700 B.n699 163.367
R1422 B.n699 B.n698 163.367
R1423 B.n698 B.n9 163.367
R1424 B.n694 B.n9 163.367
R1425 B.n694 B.n693 163.367
R1426 B.n693 B.n692 163.367
R1427 B.n692 B.n11 163.367
R1428 B.n688 B.n11 163.367
R1429 B.n688 B.n687 163.367
R1430 B.n687 B.n686 163.367
R1431 B.n686 B.n13 163.367
R1432 B.n682 B.n13 163.367
R1433 B.n682 B.n681 163.367
R1434 B.n681 B.n680 163.367
R1435 B.n680 B.n15 163.367
R1436 B.n676 B.n15 163.367
R1437 B.n676 B.n675 163.367
R1438 B.n675 B.n674 163.367
R1439 B.n674 B.n17 163.367
R1440 B.n670 B.n17 163.367
R1441 B.n670 B.n669 163.367
R1442 B.n237 B.n236 163.367
R1443 B.n237 B.n170 163.367
R1444 B.n241 B.n170 163.367
R1445 B.n242 B.n241 163.367
R1446 B.n243 B.n242 163.367
R1447 B.n243 B.n168 163.367
R1448 B.n247 B.n168 163.367
R1449 B.n248 B.n247 163.367
R1450 B.n249 B.n248 163.367
R1451 B.n249 B.n166 163.367
R1452 B.n253 B.n166 163.367
R1453 B.n254 B.n253 163.367
R1454 B.n255 B.n254 163.367
R1455 B.n255 B.n164 163.367
R1456 B.n259 B.n164 163.367
R1457 B.n260 B.n259 163.367
R1458 B.n261 B.n260 163.367
R1459 B.n261 B.n162 163.367
R1460 B.n265 B.n162 163.367
R1461 B.n266 B.n265 163.367
R1462 B.n267 B.n266 163.367
R1463 B.n267 B.n160 163.367
R1464 B.n271 B.n160 163.367
R1465 B.n272 B.n271 163.367
R1466 B.n273 B.n272 163.367
R1467 B.n273 B.n158 163.367
R1468 B.n277 B.n158 163.367
R1469 B.n278 B.n277 163.367
R1470 B.n279 B.n278 163.367
R1471 B.n279 B.n156 163.367
R1472 B.n283 B.n156 163.367
R1473 B.n284 B.n283 163.367
R1474 B.n285 B.n284 163.367
R1475 B.n285 B.n154 163.367
R1476 B.n289 B.n154 163.367
R1477 B.n290 B.n289 163.367
R1478 B.n291 B.n290 163.367
R1479 B.n291 B.n152 163.367
R1480 B.n295 B.n152 163.367
R1481 B.n296 B.n295 163.367
R1482 B.n297 B.n296 163.367
R1483 B.n297 B.n150 163.367
R1484 B.n301 B.n150 163.367
R1485 B.n302 B.n301 163.367
R1486 B.n303 B.n302 163.367
R1487 B.n303 B.n148 163.367
R1488 B.n307 B.n148 163.367
R1489 B.n308 B.n307 163.367
R1490 B.n309 B.n308 163.367
R1491 B.n309 B.n144 163.367
R1492 B.n314 B.n144 163.367
R1493 B.n315 B.n314 163.367
R1494 B.n316 B.n315 163.367
R1495 B.n316 B.n142 163.367
R1496 B.n320 B.n142 163.367
R1497 B.n321 B.n320 163.367
R1498 B.n322 B.n321 163.367
R1499 B.n322 B.n140 163.367
R1500 B.n326 B.n140 163.367
R1501 B.n327 B.n326 163.367
R1502 B.n327 B.n136 163.367
R1503 B.n331 B.n136 163.367
R1504 B.n332 B.n331 163.367
R1505 B.n333 B.n332 163.367
R1506 B.n333 B.n134 163.367
R1507 B.n337 B.n134 163.367
R1508 B.n338 B.n337 163.367
R1509 B.n339 B.n338 163.367
R1510 B.n339 B.n132 163.367
R1511 B.n343 B.n132 163.367
R1512 B.n344 B.n343 163.367
R1513 B.n345 B.n344 163.367
R1514 B.n345 B.n130 163.367
R1515 B.n349 B.n130 163.367
R1516 B.n350 B.n349 163.367
R1517 B.n351 B.n350 163.367
R1518 B.n351 B.n128 163.367
R1519 B.n355 B.n128 163.367
R1520 B.n356 B.n355 163.367
R1521 B.n357 B.n356 163.367
R1522 B.n357 B.n126 163.367
R1523 B.n361 B.n126 163.367
R1524 B.n362 B.n361 163.367
R1525 B.n363 B.n362 163.367
R1526 B.n363 B.n124 163.367
R1527 B.n367 B.n124 163.367
R1528 B.n368 B.n367 163.367
R1529 B.n369 B.n368 163.367
R1530 B.n369 B.n122 163.367
R1531 B.n373 B.n122 163.367
R1532 B.n374 B.n373 163.367
R1533 B.n375 B.n374 163.367
R1534 B.n375 B.n120 163.367
R1535 B.n379 B.n120 163.367
R1536 B.n380 B.n379 163.367
R1537 B.n381 B.n380 163.367
R1538 B.n381 B.n118 163.367
R1539 B.n385 B.n118 163.367
R1540 B.n386 B.n385 163.367
R1541 B.n387 B.n386 163.367
R1542 B.n387 B.n116 163.367
R1543 B.n391 B.n116 163.367
R1544 B.n392 B.n391 163.367
R1545 B.n393 B.n392 163.367
R1546 B.n393 B.n114 163.367
R1547 B.n397 B.n114 163.367
R1548 B.n398 B.n397 163.367
R1549 B.n399 B.n398 163.367
R1550 B.n399 B.n112 163.367
R1551 B.n404 B.n403 163.367
R1552 B.n405 B.n404 163.367
R1553 B.n405 B.n110 163.367
R1554 B.n409 B.n110 163.367
R1555 B.n410 B.n409 163.367
R1556 B.n411 B.n410 163.367
R1557 B.n411 B.n108 163.367
R1558 B.n415 B.n108 163.367
R1559 B.n416 B.n415 163.367
R1560 B.n417 B.n416 163.367
R1561 B.n417 B.n106 163.367
R1562 B.n421 B.n106 163.367
R1563 B.n422 B.n421 163.367
R1564 B.n423 B.n422 163.367
R1565 B.n423 B.n104 163.367
R1566 B.n427 B.n104 163.367
R1567 B.n428 B.n427 163.367
R1568 B.n429 B.n428 163.367
R1569 B.n429 B.n102 163.367
R1570 B.n433 B.n102 163.367
R1571 B.n434 B.n433 163.367
R1572 B.n435 B.n434 163.367
R1573 B.n435 B.n100 163.367
R1574 B.n439 B.n100 163.367
R1575 B.n440 B.n439 163.367
R1576 B.n441 B.n440 163.367
R1577 B.n441 B.n98 163.367
R1578 B.n445 B.n98 163.367
R1579 B.n446 B.n445 163.367
R1580 B.n447 B.n446 163.367
R1581 B.n447 B.n96 163.367
R1582 B.n451 B.n96 163.367
R1583 B.n452 B.n451 163.367
R1584 B.n453 B.n452 163.367
R1585 B.n453 B.n94 163.367
R1586 B.n457 B.n94 163.367
R1587 B.n458 B.n457 163.367
R1588 B.n459 B.n458 163.367
R1589 B.n459 B.n92 163.367
R1590 B.n463 B.n92 163.367
R1591 B.n464 B.n463 163.367
R1592 B.n465 B.n464 163.367
R1593 B.n465 B.n90 163.367
R1594 B.n469 B.n90 163.367
R1595 B.n470 B.n469 163.367
R1596 B.n471 B.n470 163.367
R1597 B.n471 B.n88 163.367
R1598 B.n475 B.n88 163.367
R1599 B.n476 B.n475 163.367
R1600 B.n477 B.n476 163.367
R1601 B.n477 B.n86 163.367
R1602 B.n481 B.n86 163.367
R1603 B.n482 B.n481 163.367
R1604 B.n483 B.n482 163.367
R1605 B.n483 B.n84 163.367
R1606 B.n487 B.n84 163.367
R1607 B.n488 B.n487 163.367
R1608 B.n489 B.n488 163.367
R1609 B.n489 B.n82 163.367
R1610 B.n493 B.n82 163.367
R1611 B.n494 B.n493 163.367
R1612 B.n495 B.n494 163.367
R1613 B.n495 B.n80 163.367
R1614 B.n499 B.n80 163.367
R1615 B.n500 B.n499 163.367
R1616 B.n501 B.n500 163.367
R1617 B.n668 B.n19 163.367
R1618 B.n664 B.n19 163.367
R1619 B.n664 B.n663 163.367
R1620 B.n663 B.n662 163.367
R1621 B.n662 B.n21 163.367
R1622 B.n658 B.n21 163.367
R1623 B.n658 B.n657 163.367
R1624 B.n657 B.n656 163.367
R1625 B.n656 B.n23 163.367
R1626 B.n652 B.n23 163.367
R1627 B.n652 B.n651 163.367
R1628 B.n651 B.n650 163.367
R1629 B.n650 B.n25 163.367
R1630 B.n646 B.n25 163.367
R1631 B.n646 B.n645 163.367
R1632 B.n645 B.n644 163.367
R1633 B.n644 B.n27 163.367
R1634 B.n640 B.n27 163.367
R1635 B.n640 B.n639 163.367
R1636 B.n639 B.n638 163.367
R1637 B.n638 B.n29 163.367
R1638 B.n634 B.n29 163.367
R1639 B.n634 B.n633 163.367
R1640 B.n633 B.n632 163.367
R1641 B.n632 B.n31 163.367
R1642 B.n628 B.n31 163.367
R1643 B.n628 B.n627 163.367
R1644 B.n627 B.n626 163.367
R1645 B.n626 B.n33 163.367
R1646 B.n622 B.n33 163.367
R1647 B.n622 B.n621 163.367
R1648 B.n621 B.n620 163.367
R1649 B.n620 B.n35 163.367
R1650 B.n616 B.n35 163.367
R1651 B.n616 B.n615 163.367
R1652 B.n615 B.n614 163.367
R1653 B.n614 B.n37 163.367
R1654 B.n610 B.n37 163.367
R1655 B.n610 B.n609 163.367
R1656 B.n609 B.n608 163.367
R1657 B.n608 B.n39 163.367
R1658 B.n604 B.n39 163.367
R1659 B.n604 B.n603 163.367
R1660 B.n603 B.n602 163.367
R1661 B.n602 B.n41 163.367
R1662 B.n598 B.n41 163.367
R1663 B.n598 B.n597 163.367
R1664 B.n597 B.n596 163.367
R1665 B.n596 B.n43 163.367
R1666 B.n591 B.n43 163.367
R1667 B.n591 B.n590 163.367
R1668 B.n590 B.n589 163.367
R1669 B.n589 B.n47 163.367
R1670 B.n585 B.n47 163.367
R1671 B.n585 B.n584 163.367
R1672 B.n584 B.n583 163.367
R1673 B.n583 B.n49 163.367
R1674 B.n579 B.n49 163.367
R1675 B.n579 B.n578 163.367
R1676 B.n578 B.n577 163.367
R1677 B.n577 B.n51 163.367
R1678 B.n573 B.n51 163.367
R1679 B.n573 B.n572 163.367
R1680 B.n572 B.n571 163.367
R1681 B.n571 B.n56 163.367
R1682 B.n567 B.n56 163.367
R1683 B.n567 B.n566 163.367
R1684 B.n566 B.n565 163.367
R1685 B.n565 B.n58 163.367
R1686 B.n561 B.n58 163.367
R1687 B.n561 B.n560 163.367
R1688 B.n560 B.n559 163.367
R1689 B.n559 B.n60 163.367
R1690 B.n555 B.n60 163.367
R1691 B.n555 B.n554 163.367
R1692 B.n554 B.n553 163.367
R1693 B.n553 B.n62 163.367
R1694 B.n549 B.n62 163.367
R1695 B.n549 B.n548 163.367
R1696 B.n548 B.n547 163.367
R1697 B.n547 B.n64 163.367
R1698 B.n543 B.n64 163.367
R1699 B.n543 B.n542 163.367
R1700 B.n542 B.n541 163.367
R1701 B.n541 B.n66 163.367
R1702 B.n537 B.n66 163.367
R1703 B.n537 B.n536 163.367
R1704 B.n536 B.n535 163.367
R1705 B.n535 B.n68 163.367
R1706 B.n531 B.n68 163.367
R1707 B.n531 B.n530 163.367
R1708 B.n530 B.n529 163.367
R1709 B.n529 B.n70 163.367
R1710 B.n525 B.n70 163.367
R1711 B.n525 B.n524 163.367
R1712 B.n524 B.n523 163.367
R1713 B.n523 B.n72 163.367
R1714 B.n519 B.n72 163.367
R1715 B.n519 B.n518 163.367
R1716 B.n518 B.n517 163.367
R1717 B.n517 B.n74 163.367
R1718 B.n513 B.n74 163.367
R1719 B.n513 B.n512 163.367
R1720 B.n512 B.n511 163.367
R1721 B.n511 B.n76 163.367
R1722 B.n507 B.n76 163.367
R1723 B.n507 B.n506 163.367
R1724 B.n506 B.n505 163.367
R1725 B.n505 B.n78 163.367
R1726 B.n139 B.n138 59.5399
R1727 B.n311 B.n146 59.5399
R1728 B.n593 B.n45 59.5399
R1729 B.n54 B.n53 59.5399
R1730 B.n138 B.n137 55.0793
R1731 B.n146 B.n145 55.0793
R1732 B.n45 B.n44 55.0793
R1733 B.n53 B.n52 55.0793
R1734 B.n503 B.n502 34.8103
R1735 B.n667 B.n18 34.8103
R1736 B.n402 B.n401 34.8103
R1737 B.n234 B.n171 34.8103
R1738 B B.n719 18.0485
R1739 B.n667 B.n666 10.6151
R1740 B.n666 B.n665 10.6151
R1741 B.n665 B.n20 10.6151
R1742 B.n661 B.n20 10.6151
R1743 B.n661 B.n660 10.6151
R1744 B.n660 B.n659 10.6151
R1745 B.n659 B.n22 10.6151
R1746 B.n655 B.n22 10.6151
R1747 B.n655 B.n654 10.6151
R1748 B.n654 B.n653 10.6151
R1749 B.n653 B.n24 10.6151
R1750 B.n649 B.n24 10.6151
R1751 B.n649 B.n648 10.6151
R1752 B.n648 B.n647 10.6151
R1753 B.n647 B.n26 10.6151
R1754 B.n643 B.n26 10.6151
R1755 B.n643 B.n642 10.6151
R1756 B.n642 B.n641 10.6151
R1757 B.n641 B.n28 10.6151
R1758 B.n637 B.n28 10.6151
R1759 B.n637 B.n636 10.6151
R1760 B.n636 B.n635 10.6151
R1761 B.n635 B.n30 10.6151
R1762 B.n631 B.n30 10.6151
R1763 B.n631 B.n630 10.6151
R1764 B.n630 B.n629 10.6151
R1765 B.n629 B.n32 10.6151
R1766 B.n625 B.n32 10.6151
R1767 B.n625 B.n624 10.6151
R1768 B.n624 B.n623 10.6151
R1769 B.n623 B.n34 10.6151
R1770 B.n619 B.n34 10.6151
R1771 B.n619 B.n618 10.6151
R1772 B.n618 B.n617 10.6151
R1773 B.n617 B.n36 10.6151
R1774 B.n613 B.n36 10.6151
R1775 B.n613 B.n612 10.6151
R1776 B.n612 B.n611 10.6151
R1777 B.n611 B.n38 10.6151
R1778 B.n607 B.n38 10.6151
R1779 B.n607 B.n606 10.6151
R1780 B.n606 B.n605 10.6151
R1781 B.n605 B.n40 10.6151
R1782 B.n601 B.n40 10.6151
R1783 B.n601 B.n600 10.6151
R1784 B.n600 B.n599 10.6151
R1785 B.n599 B.n42 10.6151
R1786 B.n595 B.n42 10.6151
R1787 B.n595 B.n594 10.6151
R1788 B.n592 B.n46 10.6151
R1789 B.n588 B.n46 10.6151
R1790 B.n588 B.n587 10.6151
R1791 B.n587 B.n586 10.6151
R1792 B.n586 B.n48 10.6151
R1793 B.n582 B.n48 10.6151
R1794 B.n582 B.n581 10.6151
R1795 B.n581 B.n580 10.6151
R1796 B.n580 B.n50 10.6151
R1797 B.n576 B.n575 10.6151
R1798 B.n575 B.n574 10.6151
R1799 B.n574 B.n55 10.6151
R1800 B.n570 B.n55 10.6151
R1801 B.n570 B.n569 10.6151
R1802 B.n569 B.n568 10.6151
R1803 B.n568 B.n57 10.6151
R1804 B.n564 B.n57 10.6151
R1805 B.n564 B.n563 10.6151
R1806 B.n563 B.n562 10.6151
R1807 B.n562 B.n59 10.6151
R1808 B.n558 B.n59 10.6151
R1809 B.n558 B.n557 10.6151
R1810 B.n557 B.n556 10.6151
R1811 B.n556 B.n61 10.6151
R1812 B.n552 B.n61 10.6151
R1813 B.n552 B.n551 10.6151
R1814 B.n551 B.n550 10.6151
R1815 B.n550 B.n63 10.6151
R1816 B.n546 B.n63 10.6151
R1817 B.n546 B.n545 10.6151
R1818 B.n545 B.n544 10.6151
R1819 B.n544 B.n65 10.6151
R1820 B.n540 B.n65 10.6151
R1821 B.n540 B.n539 10.6151
R1822 B.n539 B.n538 10.6151
R1823 B.n538 B.n67 10.6151
R1824 B.n534 B.n67 10.6151
R1825 B.n534 B.n533 10.6151
R1826 B.n533 B.n532 10.6151
R1827 B.n532 B.n69 10.6151
R1828 B.n528 B.n69 10.6151
R1829 B.n528 B.n527 10.6151
R1830 B.n527 B.n526 10.6151
R1831 B.n526 B.n71 10.6151
R1832 B.n522 B.n71 10.6151
R1833 B.n522 B.n521 10.6151
R1834 B.n521 B.n520 10.6151
R1835 B.n520 B.n73 10.6151
R1836 B.n516 B.n73 10.6151
R1837 B.n516 B.n515 10.6151
R1838 B.n515 B.n514 10.6151
R1839 B.n514 B.n75 10.6151
R1840 B.n510 B.n75 10.6151
R1841 B.n510 B.n509 10.6151
R1842 B.n509 B.n508 10.6151
R1843 B.n508 B.n77 10.6151
R1844 B.n504 B.n77 10.6151
R1845 B.n504 B.n503 10.6151
R1846 B.n402 B.n111 10.6151
R1847 B.n406 B.n111 10.6151
R1848 B.n407 B.n406 10.6151
R1849 B.n408 B.n407 10.6151
R1850 B.n408 B.n109 10.6151
R1851 B.n412 B.n109 10.6151
R1852 B.n413 B.n412 10.6151
R1853 B.n414 B.n413 10.6151
R1854 B.n414 B.n107 10.6151
R1855 B.n418 B.n107 10.6151
R1856 B.n419 B.n418 10.6151
R1857 B.n420 B.n419 10.6151
R1858 B.n420 B.n105 10.6151
R1859 B.n424 B.n105 10.6151
R1860 B.n425 B.n424 10.6151
R1861 B.n426 B.n425 10.6151
R1862 B.n426 B.n103 10.6151
R1863 B.n430 B.n103 10.6151
R1864 B.n431 B.n430 10.6151
R1865 B.n432 B.n431 10.6151
R1866 B.n432 B.n101 10.6151
R1867 B.n436 B.n101 10.6151
R1868 B.n437 B.n436 10.6151
R1869 B.n438 B.n437 10.6151
R1870 B.n438 B.n99 10.6151
R1871 B.n442 B.n99 10.6151
R1872 B.n443 B.n442 10.6151
R1873 B.n444 B.n443 10.6151
R1874 B.n444 B.n97 10.6151
R1875 B.n448 B.n97 10.6151
R1876 B.n449 B.n448 10.6151
R1877 B.n450 B.n449 10.6151
R1878 B.n450 B.n95 10.6151
R1879 B.n454 B.n95 10.6151
R1880 B.n455 B.n454 10.6151
R1881 B.n456 B.n455 10.6151
R1882 B.n456 B.n93 10.6151
R1883 B.n460 B.n93 10.6151
R1884 B.n461 B.n460 10.6151
R1885 B.n462 B.n461 10.6151
R1886 B.n462 B.n91 10.6151
R1887 B.n466 B.n91 10.6151
R1888 B.n467 B.n466 10.6151
R1889 B.n468 B.n467 10.6151
R1890 B.n468 B.n89 10.6151
R1891 B.n472 B.n89 10.6151
R1892 B.n473 B.n472 10.6151
R1893 B.n474 B.n473 10.6151
R1894 B.n474 B.n87 10.6151
R1895 B.n478 B.n87 10.6151
R1896 B.n479 B.n478 10.6151
R1897 B.n480 B.n479 10.6151
R1898 B.n480 B.n85 10.6151
R1899 B.n484 B.n85 10.6151
R1900 B.n485 B.n484 10.6151
R1901 B.n486 B.n485 10.6151
R1902 B.n486 B.n83 10.6151
R1903 B.n490 B.n83 10.6151
R1904 B.n491 B.n490 10.6151
R1905 B.n492 B.n491 10.6151
R1906 B.n492 B.n81 10.6151
R1907 B.n496 B.n81 10.6151
R1908 B.n497 B.n496 10.6151
R1909 B.n498 B.n497 10.6151
R1910 B.n498 B.n79 10.6151
R1911 B.n502 B.n79 10.6151
R1912 B.n238 B.n171 10.6151
R1913 B.n239 B.n238 10.6151
R1914 B.n240 B.n239 10.6151
R1915 B.n240 B.n169 10.6151
R1916 B.n244 B.n169 10.6151
R1917 B.n245 B.n244 10.6151
R1918 B.n246 B.n245 10.6151
R1919 B.n246 B.n167 10.6151
R1920 B.n250 B.n167 10.6151
R1921 B.n251 B.n250 10.6151
R1922 B.n252 B.n251 10.6151
R1923 B.n252 B.n165 10.6151
R1924 B.n256 B.n165 10.6151
R1925 B.n257 B.n256 10.6151
R1926 B.n258 B.n257 10.6151
R1927 B.n258 B.n163 10.6151
R1928 B.n262 B.n163 10.6151
R1929 B.n263 B.n262 10.6151
R1930 B.n264 B.n263 10.6151
R1931 B.n264 B.n161 10.6151
R1932 B.n268 B.n161 10.6151
R1933 B.n269 B.n268 10.6151
R1934 B.n270 B.n269 10.6151
R1935 B.n270 B.n159 10.6151
R1936 B.n274 B.n159 10.6151
R1937 B.n275 B.n274 10.6151
R1938 B.n276 B.n275 10.6151
R1939 B.n276 B.n157 10.6151
R1940 B.n280 B.n157 10.6151
R1941 B.n281 B.n280 10.6151
R1942 B.n282 B.n281 10.6151
R1943 B.n282 B.n155 10.6151
R1944 B.n286 B.n155 10.6151
R1945 B.n287 B.n286 10.6151
R1946 B.n288 B.n287 10.6151
R1947 B.n288 B.n153 10.6151
R1948 B.n292 B.n153 10.6151
R1949 B.n293 B.n292 10.6151
R1950 B.n294 B.n293 10.6151
R1951 B.n294 B.n151 10.6151
R1952 B.n298 B.n151 10.6151
R1953 B.n299 B.n298 10.6151
R1954 B.n300 B.n299 10.6151
R1955 B.n300 B.n149 10.6151
R1956 B.n304 B.n149 10.6151
R1957 B.n305 B.n304 10.6151
R1958 B.n306 B.n305 10.6151
R1959 B.n306 B.n147 10.6151
R1960 B.n310 B.n147 10.6151
R1961 B.n313 B.n312 10.6151
R1962 B.n313 B.n143 10.6151
R1963 B.n317 B.n143 10.6151
R1964 B.n318 B.n317 10.6151
R1965 B.n319 B.n318 10.6151
R1966 B.n319 B.n141 10.6151
R1967 B.n323 B.n141 10.6151
R1968 B.n324 B.n323 10.6151
R1969 B.n325 B.n324 10.6151
R1970 B.n329 B.n328 10.6151
R1971 B.n330 B.n329 10.6151
R1972 B.n330 B.n135 10.6151
R1973 B.n334 B.n135 10.6151
R1974 B.n335 B.n334 10.6151
R1975 B.n336 B.n335 10.6151
R1976 B.n336 B.n133 10.6151
R1977 B.n340 B.n133 10.6151
R1978 B.n341 B.n340 10.6151
R1979 B.n342 B.n341 10.6151
R1980 B.n342 B.n131 10.6151
R1981 B.n346 B.n131 10.6151
R1982 B.n347 B.n346 10.6151
R1983 B.n348 B.n347 10.6151
R1984 B.n348 B.n129 10.6151
R1985 B.n352 B.n129 10.6151
R1986 B.n353 B.n352 10.6151
R1987 B.n354 B.n353 10.6151
R1988 B.n354 B.n127 10.6151
R1989 B.n358 B.n127 10.6151
R1990 B.n359 B.n358 10.6151
R1991 B.n360 B.n359 10.6151
R1992 B.n360 B.n125 10.6151
R1993 B.n364 B.n125 10.6151
R1994 B.n365 B.n364 10.6151
R1995 B.n366 B.n365 10.6151
R1996 B.n366 B.n123 10.6151
R1997 B.n370 B.n123 10.6151
R1998 B.n371 B.n370 10.6151
R1999 B.n372 B.n371 10.6151
R2000 B.n372 B.n121 10.6151
R2001 B.n376 B.n121 10.6151
R2002 B.n377 B.n376 10.6151
R2003 B.n378 B.n377 10.6151
R2004 B.n378 B.n119 10.6151
R2005 B.n382 B.n119 10.6151
R2006 B.n383 B.n382 10.6151
R2007 B.n384 B.n383 10.6151
R2008 B.n384 B.n117 10.6151
R2009 B.n388 B.n117 10.6151
R2010 B.n389 B.n388 10.6151
R2011 B.n390 B.n389 10.6151
R2012 B.n390 B.n115 10.6151
R2013 B.n394 B.n115 10.6151
R2014 B.n395 B.n394 10.6151
R2015 B.n396 B.n395 10.6151
R2016 B.n396 B.n113 10.6151
R2017 B.n400 B.n113 10.6151
R2018 B.n401 B.n400 10.6151
R2019 B.n234 B.n233 10.6151
R2020 B.n233 B.n232 10.6151
R2021 B.n232 B.n173 10.6151
R2022 B.n228 B.n173 10.6151
R2023 B.n228 B.n227 10.6151
R2024 B.n227 B.n226 10.6151
R2025 B.n226 B.n175 10.6151
R2026 B.n222 B.n175 10.6151
R2027 B.n222 B.n221 10.6151
R2028 B.n221 B.n220 10.6151
R2029 B.n220 B.n177 10.6151
R2030 B.n216 B.n177 10.6151
R2031 B.n216 B.n215 10.6151
R2032 B.n215 B.n214 10.6151
R2033 B.n214 B.n179 10.6151
R2034 B.n210 B.n179 10.6151
R2035 B.n210 B.n209 10.6151
R2036 B.n209 B.n208 10.6151
R2037 B.n208 B.n181 10.6151
R2038 B.n204 B.n181 10.6151
R2039 B.n204 B.n203 10.6151
R2040 B.n203 B.n202 10.6151
R2041 B.n202 B.n183 10.6151
R2042 B.n198 B.n183 10.6151
R2043 B.n198 B.n197 10.6151
R2044 B.n197 B.n196 10.6151
R2045 B.n196 B.n185 10.6151
R2046 B.n192 B.n185 10.6151
R2047 B.n192 B.n191 10.6151
R2048 B.n191 B.n190 10.6151
R2049 B.n190 B.n187 10.6151
R2050 B.n187 B.n0 10.6151
R2051 B.n715 B.n1 10.6151
R2052 B.n715 B.n714 10.6151
R2053 B.n714 B.n713 10.6151
R2054 B.n713 B.n4 10.6151
R2055 B.n709 B.n4 10.6151
R2056 B.n709 B.n708 10.6151
R2057 B.n708 B.n707 10.6151
R2058 B.n707 B.n6 10.6151
R2059 B.n703 B.n6 10.6151
R2060 B.n703 B.n702 10.6151
R2061 B.n702 B.n701 10.6151
R2062 B.n701 B.n8 10.6151
R2063 B.n697 B.n8 10.6151
R2064 B.n697 B.n696 10.6151
R2065 B.n696 B.n695 10.6151
R2066 B.n695 B.n10 10.6151
R2067 B.n691 B.n10 10.6151
R2068 B.n691 B.n690 10.6151
R2069 B.n690 B.n689 10.6151
R2070 B.n689 B.n12 10.6151
R2071 B.n685 B.n12 10.6151
R2072 B.n685 B.n684 10.6151
R2073 B.n684 B.n683 10.6151
R2074 B.n683 B.n14 10.6151
R2075 B.n679 B.n14 10.6151
R2076 B.n679 B.n678 10.6151
R2077 B.n678 B.n677 10.6151
R2078 B.n677 B.n16 10.6151
R2079 B.n673 B.n16 10.6151
R2080 B.n673 B.n672 10.6151
R2081 B.n672 B.n671 10.6151
R2082 B.n671 B.n18 10.6151
R2083 B.n594 B.n593 9.36635
R2084 B.n576 B.n54 9.36635
R2085 B.n311 B.n310 9.36635
R2086 B.n328 B.n139 9.36635
R2087 B.n719 B.n0 2.81026
R2088 B.n719 B.n1 2.81026
R2089 B.n593 B.n592 1.24928
R2090 B.n54 B.n50 1.24928
R2091 B.n312 B.n311 1.24928
R2092 B.n325 B.n139 1.24928
R2093 VP.n4 VP.t0 179.035
R2094 VP.n4 VP.t3 178.274
R2095 VP.n14 VP.n0 161.3
R2096 VP.n13 VP.n12 161.3
R2097 VP.n11 VP.n1 161.3
R2098 VP.n10 VP.n9 161.3
R2099 VP.n8 VP.n2 161.3
R2100 VP.n7 VP.n6 161.3
R2101 VP.n3 VP.t1 143.448
R2102 VP.n15 VP.t2 143.448
R2103 VP.n5 VP.n3 102.547
R2104 VP.n16 VP.n15 102.547
R2105 VP.n9 VP.n1 56.5617
R2106 VP.n5 VP.n4 52.7127
R2107 VP.n8 VP.n7 24.5923
R2108 VP.n9 VP.n8 24.5923
R2109 VP.n13 VP.n1 24.5923
R2110 VP.n14 VP.n13 24.5923
R2111 VP.n7 VP.n3 8.36172
R2112 VP.n15 VP.n14 8.36172
R2113 VP.n6 VP.n5 0.278335
R2114 VP.n16 VP.n0 0.278335
R2115 VP.n6 VP.n2 0.189894
R2116 VP.n10 VP.n2 0.189894
R2117 VP.n11 VP.n10 0.189894
R2118 VP.n12 VP.n11 0.189894
R2119 VP.n12 VP.n0 0.189894
R2120 VP VP.n16 0.153485
R2121 VDD1 VDD1.n1 114.356
R2122 VDD1 VDD1.n0 69.9502
R2123 VDD1.n0 VDD1.t3 2.1762
R2124 VDD1.n0 VDD1.t0 2.1762
R2125 VDD1.n1 VDD1.t2 2.1762
R2126 VDD1.n1 VDD1.t1 2.1762
C0 VTAIL VDD1 6.10319f
C1 VDD2 w_n2674_n3956# 1.57169f
C2 VP VDD1 6.03522f
C3 VN VDD1 0.149386f
C4 B w_n2674_n3956# 9.960099f
C5 VTAIL VP 5.58051f
C6 VTAIL VN 5.5664f
C7 VDD1 w_n2674_n3956# 1.51754f
C8 VN VP 6.66785f
C9 VDD2 B 1.37461f
C10 VTAIL w_n2674_n3956# 4.63651f
C11 VP w_n2674_n3956# 4.9068f
C12 VDD2 VDD1 1.01206f
C13 VN w_n2674_n3956# 4.56328f
C14 B VDD1 1.32396f
C15 VDD2 VTAIL 6.15679f
C16 B VTAIL 5.86541f
C17 VDD2 VP 0.389046f
C18 VDD2 VN 5.79628f
C19 B VP 1.69945f
C20 B VN 1.1298f
C21 VDD2 VSUBS 0.993058f
C22 VDD1 VSUBS 6.04188f
C23 VTAIL VSUBS 1.34267f
C24 VN VSUBS 5.52491f
C25 VP VSUBS 2.342796f
C26 B VSUBS 4.448296f
C27 w_n2674_n3956# VSUBS 0.129732p
C28 VDD1.t3 VSUBS 0.315502f
C29 VDD1.t0 VSUBS 0.315502f
C30 VDD1.n0 VSUBS 2.5427f
C31 VDD1.t2 VSUBS 0.315502f
C32 VDD1.t1 VSUBS 0.315502f
C33 VDD1.n1 VSUBS 3.40458f
C34 VP.n0 VSUBS 0.043013f
C35 VP.t2 VSUBS 3.35228f
C36 VP.n1 VSUBS 0.047428f
C37 VP.n2 VSUBS 0.032627f
C38 VP.t1 VSUBS 3.35228f
C39 VP.n3 VSUBS 1.27464f
C40 VP.t3 VSUBS 3.62014f
C41 VP.t0 VSUBS 3.62589f
C42 VP.n4 VSUBS 4.17589f
C43 VP.n5 VSUBS 1.91844f
C44 VP.n6 VSUBS 0.043013f
C45 VP.n7 VSUBS 0.04079f
C46 VP.n8 VSUBS 0.060503f
C47 VP.n9 VSUBS 0.047428f
C48 VP.n10 VSUBS 0.032627f
C49 VP.n11 VSUBS 0.032627f
C50 VP.n12 VSUBS 0.032627f
C51 VP.n13 VSUBS 0.060503f
C52 VP.n14 VSUBS 0.04079f
C53 VP.n15 VSUBS 1.27464f
C54 VP.n16 VSUBS 0.053442f
C55 B.n0 VSUBS 0.004059f
C56 B.n1 VSUBS 0.004059f
C57 B.n2 VSUBS 0.006419f
C58 B.n3 VSUBS 0.006419f
C59 B.n4 VSUBS 0.006419f
C60 B.n5 VSUBS 0.006419f
C61 B.n6 VSUBS 0.006419f
C62 B.n7 VSUBS 0.006419f
C63 B.n8 VSUBS 0.006419f
C64 B.n9 VSUBS 0.006419f
C65 B.n10 VSUBS 0.006419f
C66 B.n11 VSUBS 0.006419f
C67 B.n12 VSUBS 0.006419f
C68 B.n13 VSUBS 0.006419f
C69 B.n14 VSUBS 0.006419f
C70 B.n15 VSUBS 0.006419f
C71 B.n16 VSUBS 0.006419f
C72 B.n17 VSUBS 0.006419f
C73 B.n18 VSUBS 0.015262f
C74 B.n19 VSUBS 0.006419f
C75 B.n20 VSUBS 0.006419f
C76 B.n21 VSUBS 0.006419f
C77 B.n22 VSUBS 0.006419f
C78 B.n23 VSUBS 0.006419f
C79 B.n24 VSUBS 0.006419f
C80 B.n25 VSUBS 0.006419f
C81 B.n26 VSUBS 0.006419f
C82 B.n27 VSUBS 0.006419f
C83 B.n28 VSUBS 0.006419f
C84 B.n29 VSUBS 0.006419f
C85 B.n30 VSUBS 0.006419f
C86 B.n31 VSUBS 0.006419f
C87 B.n32 VSUBS 0.006419f
C88 B.n33 VSUBS 0.006419f
C89 B.n34 VSUBS 0.006419f
C90 B.n35 VSUBS 0.006419f
C91 B.n36 VSUBS 0.006419f
C92 B.n37 VSUBS 0.006419f
C93 B.n38 VSUBS 0.006419f
C94 B.n39 VSUBS 0.006419f
C95 B.n40 VSUBS 0.006419f
C96 B.n41 VSUBS 0.006419f
C97 B.n42 VSUBS 0.006419f
C98 B.n43 VSUBS 0.006419f
C99 B.t5 VSUBS 0.255334f
C100 B.t4 VSUBS 0.284598f
C101 B.t3 VSUBS 1.54055f
C102 B.n44 VSUBS 0.440593f
C103 B.n45 VSUBS 0.266233f
C104 B.n46 VSUBS 0.006419f
C105 B.n47 VSUBS 0.006419f
C106 B.n48 VSUBS 0.006419f
C107 B.n49 VSUBS 0.006419f
C108 B.n50 VSUBS 0.003587f
C109 B.n51 VSUBS 0.006419f
C110 B.t8 VSUBS 0.255337f
C111 B.t7 VSUBS 0.2846f
C112 B.t6 VSUBS 1.54055f
C113 B.n52 VSUBS 0.44059f
C114 B.n53 VSUBS 0.26623f
C115 B.n54 VSUBS 0.014872f
C116 B.n55 VSUBS 0.006419f
C117 B.n56 VSUBS 0.006419f
C118 B.n57 VSUBS 0.006419f
C119 B.n58 VSUBS 0.006419f
C120 B.n59 VSUBS 0.006419f
C121 B.n60 VSUBS 0.006419f
C122 B.n61 VSUBS 0.006419f
C123 B.n62 VSUBS 0.006419f
C124 B.n63 VSUBS 0.006419f
C125 B.n64 VSUBS 0.006419f
C126 B.n65 VSUBS 0.006419f
C127 B.n66 VSUBS 0.006419f
C128 B.n67 VSUBS 0.006419f
C129 B.n68 VSUBS 0.006419f
C130 B.n69 VSUBS 0.006419f
C131 B.n70 VSUBS 0.006419f
C132 B.n71 VSUBS 0.006419f
C133 B.n72 VSUBS 0.006419f
C134 B.n73 VSUBS 0.006419f
C135 B.n74 VSUBS 0.006419f
C136 B.n75 VSUBS 0.006419f
C137 B.n76 VSUBS 0.006419f
C138 B.n77 VSUBS 0.006419f
C139 B.n78 VSUBS 0.016078f
C140 B.n79 VSUBS 0.006419f
C141 B.n80 VSUBS 0.006419f
C142 B.n81 VSUBS 0.006419f
C143 B.n82 VSUBS 0.006419f
C144 B.n83 VSUBS 0.006419f
C145 B.n84 VSUBS 0.006419f
C146 B.n85 VSUBS 0.006419f
C147 B.n86 VSUBS 0.006419f
C148 B.n87 VSUBS 0.006419f
C149 B.n88 VSUBS 0.006419f
C150 B.n89 VSUBS 0.006419f
C151 B.n90 VSUBS 0.006419f
C152 B.n91 VSUBS 0.006419f
C153 B.n92 VSUBS 0.006419f
C154 B.n93 VSUBS 0.006419f
C155 B.n94 VSUBS 0.006419f
C156 B.n95 VSUBS 0.006419f
C157 B.n96 VSUBS 0.006419f
C158 B.n97 VSUBS 0.006419f
C159 B.n98 VSUBS 0.006419f
C160 B.n99 VSUBS 0.006419f
C161 B.n100 VSUBS 0.006419f
C162 B.n101 VSUBS 0.006419f
C163 B.n102 VSUBS 0.006419f
C164 B.n103 VSUBS 0.006419f
C165 B.n104 VSUBS 0.006419f
C166 B.n105 VSUBS 0.006419f
C167 B.n106 VSUBS 0.006419f
C168 B.n107 VSUBS 0.006419f
C169 B.n108 VSUBS 0.006419f
C170 B.n109 VSUBS 0.006419f
C171 B.n110 VSUBS 0.006419f
C172 B.n111 VSUBS 0.006419f
C173 B.n112 VSUBS 0.016078f
C174 B.n113 VSUBS 0.006419f
C175 B.n114 VSUBS 0.006419f
C176 B.n115 VSUBS 0.006419f
C177 B.n116 VSUBS 0.006419f
C178 B.n117 VSUBS 0.006419f
C179 B.n118 VSUBS 0.006419f
C180 B.n119 VSUBS 0.006419f
C181 B.n120 VSUBS 0.006419f
C182 B.n121 VSUBS 0.006419f
C183 B.n122 VSUBS 0.006419f
C184 B.n123 VSUBS 0.006419f
C185 B.n124 VSUBS 0.006419f
C186 B.n125 VSUBS 0.006419f
C187 B.n126 VSUBS 0.006419f
C188 B.n127 VSUBS 0.006419f
C189 B.n128 VSUBS 0.006419f
C190 B.n129 VSUBS 0.006419f
C191 B.n130 VSUBS 0.006419f
C192 B.n131 VSUBS 0.006419f
C193 B.n132 VSUBS 0.006419f
C194 B.n133 VSUBS 0.006419f
C195 B.n134 VSUBS 0.006419f
C196 B.n135 VSUBS 0.006419f
C197 B.n136 VSUBS 0.006419f
C198 B.t1 VSUBS 0.255337f
C199 B.t2 VSUBS 0.2846f
C200 B.t0 VSUBS 1.54055f
C201 B.n137 VSUBS 0.44059f
C202 B.n138 VSUBS 0.26623f
C203 B.n139 VSUBS 0.014872f
C204 B.n140 VSUBS 0.006419f
C205 B.n141 VSUBS 0.006419f
C206 B.n142 VSUBS 0.006419f
C207 B.n143 VSUBS 0.006419f
C208 B.n144 VSUBS 0.006419f
C209 B.t10 VSUBS 0.255334f
C210 B.t11 VSUBS 0.284598f
C211 B.t9 VSUBS 1.54055f
C212 B.n145 VSUBS 0.440593f
C213 B.n146 VSUBS 0.266233f
C214 B.n147 VSUBS 0.006419f
C215 B.n148 VSUBS 0.006419f
C216 B.n149 VSUBS 0.006419f
C217 B.n150 VSUBS 0.006419f
C218 B.n151 VSUBS 0.006419f
C219 B.n152 VSUBS 0.006419f
C220 B.n153 VSUBS 0.006419f
C221 B.n154 VSUBS 0.006419f
C222 B.n155 VSUBS 0.006419f
C223 B.n156 VSUBS 0.006419f
C224 B.n157 VSUBS 0.006419f
C225 B.n158 VSUBS 0.006419f
C226 B.n159 VSUBS 0.006419f
C227 B.n160 VSUBS 0.006419f
C228 B.n161 VSUBS 0.006419f
C229 B.n162 VSUBS 0.006419f
C230 B.n163 VSUBS 0.006419f
C231 B.n164 VSUBS 0.006419f
C232 B.n165 VSUBS 0.006419f
C233 B.n166 VSUBS 0.006419f
C234 B.n167 VSUBS 0.006419f
C235 B.n168 VSUBS 0.006419f
C236 B.n169 VSUBS 0.006419f
C237 B.n170 VSUBS 0.006419f
C238 B.n171 VSUBS 0.016078f
C239 B.n172 VSUBS 0.006419f
C240 B.n173 VSUBS 0.006419f
C241 B.n174 VSUBS 0.006419f
C242 B.n175 VSUBS 0.006419f
C243 B.n176 VSUBS 0.006419f
C244 B.n177 VSUBS 0.006419f
C245 B.n178 VSUBS 0.006419f
C246 B.n179 VSUBS 0.006419f
C247 B.n180 VSUBS 0.006419f
C248 B.n181 VSUBS 0.006419f
C249 B.n182 VSUBS 0.006419f
C250 B.n183 VSUBS 0.006419f
C251 B.n184 VSUBS 0.006419f
C252 B.n185 VSUBS 0.006419f
C253 B.n186 VSUBS 0.006419f
C254 B.n187 VSUBS 0.006419f
C255 B.n188 VSUBS 0.006419f
C256 B.n189 VSUBS 0.006419f
C257 B.n190 VSUBS 0.006419f
C258 B.n191 VSUBS 0.006419f
C259 B.n192 VSUBS 0.006419f
C260 B.n193 VSUBS 0.006419f
C261 B.n194 VSUBS 0.006419f
C262 B.n195 VSUBS 0.006419f
C263 B.n196 VSUBS 0.006419f
C264 B.n197 VSUBS 0.006419f
C265 B.n198 VSUBS 0.006419f
C266 B.n199 VSUBS 0.006419f
C267 B.n200 VSUBS 0.006419f
C268 B.n201 VSUBS 0.006419f
C269 B.n202 VSUBS 0.006419f
C270 B.n203 VSUBS 0.006419f
C271 B.n204 VSUBS 0.006419f
C272 B.n205 VSUBS 0.006419f
C273 B.n206 VSUBS 0.006419f
C274 B.n207 VSUBS 0.006419f
C275 B.n208 VSUBS 0.006419f
C276 B.n209 VSUBS 0.006419f
C277 B.n210 VSUBS 0.006419f
C278 B.n211 VSUBS 0.006419f
C279 B.n212 VSUBS 0.006419f
C280 B.n213 VSUBS 0.006419f
C281 B.n214 VSUBS 0.006419f
C282 B.n215 VSUBS 0.006419f
C283 B.n216 VSUBS 0.006419f
C284 B.n217 VSUBS 0.006419f
C285 B.n218 VSUBS 0.006419f
C286 B.n219 VSUBS 0.006419f
C287 B.n220 VSUBS 0.006419f
C288 B.n221 VSUBS 0.006419f
C289 B.n222 VSUBS 0.006419f
C290 B.n223 VSUBS 0.006419f
C291 B.n224 VSUBS 0.006419f
C292 B.n225 VSUBS 0.006419f
C293 B.n226 VSUBS 0.006419f
C294 B.n227 VSUBS 0.006419f
C295 B.n228 VSUBS 0.006419f
C296 B.n229 VSUBS 0.006419f
C297 B.n230 VSUBS 0.006419f
C298 B.n231 VSUBS 0.006419f
C299 B.n232 VSUBS 0.006419f
C300 B.n233 VSUBS 0.006419f
C301 B.n234 VSUBS 0.015262f
C302 B.n235 VSUBS 0.015262f
C303 B.n236 VSUBS 0.016078f
C304 B.n237 VSUBS 0.006419f
C305 B.n238 VSUBS 0.006419f
C306 B.n239 VSUBS 0.006419f
C307 B.n240 VSUBS 0.006419f
C308 B.n241 VSUBS 0.006419f
C309 B.n242 VSUBS 0.006419f
C310 B.n243 VSUBS 0.006419f
C311 B.n244 VSUBS 0.006419f
C312 B.n245 VSUBS 0.006419f
C313 B.n246 VSUBS 0.006419f
C314 B.n247 VSUBS 0.006419f
C315 B.n248 VSUBS 0.006419f
C316 B.n249 VSUBS 0.006419f
C317 B.n250 VSUBS 0.006419f
C318 B.n251 VSUBS 0.006419f
C319 B.n252 VSUBS 0.006419f
C320 B.n253 VSUBS 0.006419f
C321 B.n254 VSUBS 0.006419f
C322 B.n255 VSUBS 0.006419f
C323 B.n256 VSUBS 0.006419f
C324 B.n257 VSUBS 0.006419f
C325 B.n258 VSUBS 0.006419f
C326 B.n259 VSUBS 0.006419f
C327 B.n260 VSUBS 0.006419f
C328 B.n261 VSUBS 0.006419f
C329 B.n262 VSUBS 0.006419f
C330 B.n263 VSUBS 0.006419f
C331 B.n264 VSUBS 0.006419f
C332 B.n265 VSUBS 0.006419f
C333 B.n266 VSUBS 0.006419f
C334 B.n267 VSUBS 0.006419f
C335 B.n268 VSUBS 0.006419f
C336 B.n269 VSUBS 0.006419f
C337 B.n270 VSUBS 0.006419f
C338 B.n271 VSUBS 0.006419f
C339 B.n272 VSUBS 0.006419f
C340 B.n273 VSUBS 0.006419f
C341 B.n274 VSUBS 0.006419f
C342 B.n275 VSUBS 0.006419f
C343 B.n276 VSUBS 0.006419f
C344 B.n277 VSUBS 0.006419f
C345 B.n278 VSUBS 0.006419f
C346 B.n279 VSUBS 0.006419f
C347 B.n280 VSUBS 0.006419f
C348 B.n281 VSUBS 0.006419f
C349 B.n282 VSUBS 0.006419f
C350 B.n283 VSUBS 0.006419f
C351 B.n284 VSUBS 0.006419f
C352 B.n285 VSUBS 0.006419f
C353 B.n286 VSUBS 0.006419f
C354 B.n287 VSUBS 0.006419f
C355 B.n288 VSUBS 0.006419f
C356 B.n289 VSUBS 0.006419f
C357 B.n290 VSUBS 0.006419f
C358 B.n291 VSUBS 0.006419f
C359 B.n292 VSUBS 0.006419f
C360 B.n293 VSUBS 0.006419f
C361 B.n294 VSUBS 0.006419f
C362 B.n295 VSUBS 0.006419f
C363 B.n296 VSUBS 0.006419f
C364 B.n297 VSUBS 0.006419f
C365 B.n298 VSUBS 0.006419f
C366 B.n299 VSUBS 0.006419f
C367 B.n300 VSUBS 0.006419f
C368 B.n301 VSUBS 0.006419f
C369 B.n302 VSUBS 0.006419f
C370 B.n303 VSUBS 0.006419f
C371 B.n304 VSUBS 0.006419f
C372 B.n305 VSUBS 0.006419f
C373 B.n306 VSUBS 0.006419f
C374 B.n307 VSUBS 0.006419f
C375 B.n308 VSUBS 0.006419f
C376 B.n309 VSUBS 0.006419f
C377 B.n310 VSUBS 0.006041f
C378 B.n311 VSUBS 0.014872f
C379 B.n312 VSUBS 0.003587f
C380 B.n313 VSUBS 0.006419f
C381 B.n314 VSUBS 0.006419f
C382 B.n315 VSUBS 0.006419f
C383 B.n316 VSUBS 0.006419f
C384 B.n317 VSUBS 0.006419f
C385 B.n318 VSUBS 0.006419f
C386 B.n319 VSUBS 0.006419f
C387 B.n320 VSUBS 0.006419f
C388 B.n321 VSUBS 0.006419f
C389 B.n322 VSUBS 0.006419f
C390 B.n323 VSUBS 0.006419f
C391 B.n324 VSUBS 0.006419f
C392 B.n325 VSUBS 0.003587f
C393 B.n326 VSUBS 0.006419f
C394 B.n327 VSUBS 0.006419f
C395 B.n328 VSUBS 0.006041f
C396 B.n329 VSUBS 0.006419f
C397 B.n330 VSUBS 0.006419f
C398 B.n331 VSUBS 0.006419f
C399 B.n332 VSUBS 0.006419f
C400 B.n333 VSUBS 0.006419f
C401 B.n334 VSUBS 0.006419f
C402 B.n335 VSUBS 0.006419f
C403 B.n336 VSUBS 0.006419f
C404 B.n337 VSUBS 0.006419f
C405 B.n338 VSUBS 0.006419f
C406 B.n339 VSUBS 0.006419f
C407 B.n340 VSUBS 0.006419f
C408 B.n341 VSUBS 0.006419f
C409 B.n342 VSUBS 0.006419f
C410 B.n343 VSUBS 0.006419f
C411 B.n344 VSUBS 0.006419f
C412 B.n345 VSUBS 0.006419f
C413 B.n346 VSUBS 0.006419f
C414 B.n347 VSUBS 0.006419f
C415 B.n348 VSUBS 0.006419f
C416 B.n349 VSUBS 0.006419f
C417 B.n350 VSUBS 0.006419f
C418 B.n351 VSUBS 0.006419f
C419 B.n352 VSUBS 0.006419f
C420 B.n353 VSUBS 0.006419f
C421 B.n354 VSUBS 0.006419f
C422 B.n355 VSUBS 0.006419f
C423 B.n356 VSUBS 0.006419f
C424 B.n357 VSUBS 0.006419f
C425 B.n358 VSUBS 0.006419f
C426 B.n359 VSUBS 0.006419f
C427 B.n360 VSUBS 0.006419f
C428 B.n361 VSUBS 0.006419f
C429 B.n362 VSUBS 0.006419f
C430 B.n363 VSUBS 0.006419f
C431 B.n364 VSUBS 0.006419f
C432 B.n365 VSUBS 0.006419f
C433 B.n366 VSUBS 0.006419f
C434 B.n367 VSUBS 0.006419f
C435 B.n368 VSUBS 0.006419f
C436 B.n369 VSUBS 0.006419f
C437 B.n370 VSUBS 0.006419f
C438 B.n371 VSUBS 0.006419f
C439 B.n372 VSUBS 0.006419f
C440 B.n373 VSUBS 0.006419f
C441 B.n374 VSUBS 0.006419f
C442 B.n375 VSUBS 0.006419f
C443 B.n376 VSUBS 0.006419f
C444 B.n377 VSUBS 0.006419f
C445 B.n378 VSUBS 0.006419f
C446 B.n379 VSUBS 0.006419f
C447 B.n380 VSUBS 0.006419f
C448 B.n381 VSUBS 0.006419f
C449 B.n382 VSUBS 0.006419f
C450 B.n383 VSUBS 0.006419f
C451 B.n384 VSUBS 0.006419f
C452 B.n385 VSUBS 0.006419f
C453 B.n386 VSUBS 0.006419f
C454 B.n387 VSUBS 0.006419f
C455 B.n388 VSUBS 0.006419f
C456 B.n389 VSUBS 0.006419f
C457 B.n390 VSUBS 0.006419f
C458 B.n391 VSUBS 0.006419f
C459 B.n392 VSUBS 0.006419f
C460 B.n393 VSUBS 0.006419f
C461 B.n394 VSUBS 0.006419f
C462 B.n395 VSUBS 0.006419f
C463 B.n396 VSUBS 0.006419f
C464 B.n397 VSUBS 0.006419f
C465 B.n398 VSUBS 0.006419f
C466 B.n399 VSUBS 0.006419f
C467 B.n400 VSUBS 0.006419f
C468 B.n401 VSUBS 0.016078f
C469 B.n402 VSUBS 0.015262f
C470 B.n403 VSUBS 0.015262f
C471 B.n404 VSUBS 0.006419f
C472 B.n405 VSUBS 0.006419f
C473 B.n406 VSUBS 0.006419f
C474 B.n407 VSUBS 0.006419f
C475 B.n408 VSUBS 0.006419f
C476 B.n409 VSUBS 0.006419f
C477 B.n410 VSUBS 0.006419f
C478 B.n411 VSUBS 0.006419f
C479 B.n412 VSUBS 0.006419f
C480 B.n413 VSUBS 0.006419f
C481 B.n414 VSUBS 0.006419f
C482 B.n415 VSUBS 0.006419f
C483 B.n416 VSUBS 0.006419f
C484 B.n417 VSUBS 0.006419f
C485 B.n418 VSUBS 0.006419f
C486 B.n419 VSUBS 0.006419f
C487 B.n420 VSUBS 0.006419f
C488 B.n421 VSUBS 0.006419f
C489 B.n422 VSUBS 0.006419f
C490 B.n423 VSUBS 0.006419f
C491 B.n424 VSUBS 0.006419f
C492 B.n425 VSUBS 0.006419f
C493 B.n426 VSUBS 0.006419f
C494 B.n427 VSUBS 0.006419f
C495 B.n428 VSUBS 0.006419f
C496 B.n429 VSUBS 0.006419f
C497 B.n430 VSUBS 0.006419f
C498 B.n431 VSUBS 0.006419f
C499 B.n432 VSUBS 0.006419f
C500 B.n433 VSUBS 0.006419f
C501 B.n434 VSUBS 0.006419f
C502 B.n435 VSUBS 0.006419f
C503 B.n436 VSUBS 0.006419f
C504 B.n437 VSUBS 0.006419f
C505 B.n438 VSUBS 0.006419f
C506 B.n439 VSUBS 0.006419f
C507 B.n440 VSUBS 0.006419f
C508 B.n441 VSUBS 0.006419f
C509 B.n442 VSUBS 0.006419f
C510 B.n443 VSUBS 0.006419f
C511 B.n444 VSUBS 0.006419f
C512 B.n445 VSUBS 0.006419f
C513 B.n446 VSUBS 0.006419f
C514 B.n447 VSUBS 0.006419f
C515 B.n448 VSUBS 0.006419f
C516 B.n449 VSUBS 0.006419f
C517 B.n450 VSUBS 0.006419f
C518 B.n451 VSUBS 0.006419f
C519 B.n452 VSUBS 0.006419f
C520 B.n453 VSUBS 0.006419f
C521 B.n454 VSUBS 0.006419f
C522 B.n455 VSUBS 0.006419f
C523 B.n456 VSUBS 0.006419f
C524 B.n457 VSUBS 0.006419f
C525 B.n458 VSUBS 0.006419f
C526 B.n459 VSUBS 0.006419f
C527 B.n460 VSUBS 0.006419f
C528 B.n461 VSUBS 0.006419f
C529 B.n462 VSUBS 0.006419f
C530 B.n463 VSUBS 0.006419f
C531 B.n464 VSUBS 0.006419f
C532 B.n465 VSUBS 0.006419f
C533 B.n466 VSUBS 0.006419f
C534 B.n467 VSUBS 0.006419f
C535 B.n468 VSUBS 0.006419f
C536 B.n469 VSUBS 0.006419f
C537 B.n470 VSUBS 0.006419f
C538 B.n471 VSUBS 0.006419f
C539 B.n472 VSUBS 0.006419f
C540 B.n473 VSUBS 0.006419f
C541 B.n474 VSUBS 0.006419f
C542 B.n475 VSUBS 0.006419f
C543 B.n476 VSUBS 0.006419f
C544 B.n477 VSUBS 0.006419f
C545 B.n478 VSUBS 0.006419f
C546 B.n479 VSUBS 0.006419f
C547 B.n480 VSUBS 0.006419f
C548 B.n481 VSUBS 0.006419f
C549 B.n482 VSUBS 0.006419f
C550 B.n483 VSUBS 0.006419f
C551 B.n484 VSUBS 0.006419f
C552 B.n485 VSUBS 0.006419f
C553 B.n486 VSUBS 0.006419f
C554 B.n487 VSUBS 0.006419f
C555 B.n488 VSUBS 0.006419f
C556 B.n489 VSUBS 0.006419f
C557 B.n490 VSUBS 0.006419f
C558 B.n491 VSUBS 0.006419f
C559 B.n492 VSUBS 0.006419f
C560 B.n493 VSUBS 0.006419f
C561 B.n494 VSUBS 0.006419f
C562 B.n495 VSUBS 0.006419f
C563 B.n496 VSUBS 0.006419f
C564 B.n497 VSUBS 0.006419f
C565 B.n498 VSUBS 0.006419f
C566 B.n499 VSUBS 0.006419f
C567 B.n500 VSUBS 0.006419f
C568 B.n501 VSUBS 0.015262f
C569 B.n502 VSUBS 0.015973f
C570 B.n503 VSUBS 0.015366f
C571 B.n504 VSUBS 0.006419f
C572 B.n505 VSUBS 0.006419f
C573 B.n506 VSUBS 0.006419f
C574 B.n507 VSUBS 0.006419f
C575 B.n508 VSUBS 0.006419f
C576 B.n509 VSUBS 0.006419f
C577 B.n510 VSUBS 0.006419f
C578 B.n511 VSUBS 0.006419f
C579 B.n512 VSUBS 0.006419f
C580 B.n513 VSUBS 0.006419f
C581 B.n514 VSUBS 0.006419f
C582 B.n515 VSUBS 0.006419f
C583 B.n516 VSUBS 0.006419f
C584 B.n517 VSUBS 0.006419f
C585 B.n518 VSUBS 0.006419f
C586 B.n519 VSUBS 0.006419f
C587 B.n520 VSUBS 0.006419f
C588 B.n521 VSUBS 0.006419f
C589 B.n522 VSUBS 0.006419f
C590 B.n523 VSUBS 0.006419f
C591 B.n524 VSUBS 0.006419f
C592 B.n525 VSUBS 0.006419f
C593 B.n526 VSUBS 0.006419f
C594 B.n527 VSUBS 0.006419f
C595 B.n528 VSUBS 0.006419f
C596 B.n529 VSUBS 0.006419f
C597 B.n530 VSUBS 0.006419f
C598 B.n531 VSUBS 0.006419f
C599 B.n532 VSUBS 0.006419f
C600 B.n533 VSUBS 0.006419f
C601 B.n534 VSUBS 0.006419f
C602 B.n535 VSUBS 0.006419f
C603 B.n536 VSUBS 0.006419f
C604 B.n537 VSUBS 0.006419f
C605 B.n538 VSUBS 0.006419f
C606 B.n539 VSUBS 0.006419f
C607 B.n540 VSUBS 0.006419f
C608 B.n541 VSUBS 0.006419f
C609 B.n542 VSUBS 0.006419f
C610 B.n543 VSUBS 0.006419f
C611 B.n544 VSUBS 0.006419f
C612 B.n545 VSUBS 0.006419f
C613 B.n546 VSUBS 0.006419f
C614 B.n547 VSUBS 0.006419f
C615 B.n548 VSUBS 0.006419f
C616 B.n549 VSUBS 0.006419f
C617 B.n550 VSUBS 0.006419f
C618 B.n551 VSUBS 0.006419f
C619 B.n552 VSUBS 0.006419f
C620 B.n553 VSUBS 0.006419f
C621 B.n554 VSUBS 0.006419f
C622 B.n555 VSUBS 0.006419f
C623 B.n556 VSUBS 0.006419f
C624 B.n557 VSUBS 0.006419f
C625 B.n558 VSUBS 0.006419f
C626 B.n559 VSUBS 0.006419f
C627 B.n560 VSUBS 0.006419f
C628 B.n561 VSUBS 0.006419f
C629 B.n562 VSUBS 0.006419f
C630 B.n563 VSUBS 0.006419f
C631 B.n564 VSUBS 0.006419f
C632 B.n565 VSUBS 0.006419f
C633 B.n566 VSUBS 0.006419f
C634 B.n567 VSUBS 0.006419f
C635 B.n568 VSUBS 0.006419f
C636 B.n569 VSUBS 0.006419f
C637 B.n570 VSUBS 0.006419f
C638 B.n571 VSUBS 0.006419f
C639 B.n572 VSUBS 0.006419f
C640 B.n573 VSUBS 0.006419f
C641 B.n574 VSUBS 0.006419f
C642 B.n575 VSUBS 0.006419f
C643 B.n576 VSUBS 0.006041f
C644 B.n577 VSUBS 0.006419f
C645 B.n578 VSUBS 0.006419f
C646 B.n579 VSUBS 0.006419f
C647 B.n580 VSUBS 0.006419f
C648 B.n581 VSUBS 0.006419f
C649 B.n582 VSUBS 0.006419f
C650 B.n583 VSUBS 0.006419f
C651 B.n584 VSUBS 0.006419f
C652 B.n585 VSUBS 0.006419f
C653 B.n586 VSUBS 0.006419f
C654 B.n587 VSUBS 0.006419f
C655 B.n588 VSUBS 0.006419f
C656 B.n589 VSUBS 0.006419f
C657 B.n590 VSUBS 0.006419f
C658 B.n591 VSUBS 0.006419f
C659 B.n592 VSUBS 0.003587f
C660 B.n593 VSUBS 0.014872f
C661 B.n594 VSUBS 0.006041f
C662 B.n595 VSUBS 0.006419f
C663 B.n596 VSUBS 0.006419f
C664 B.n597 VSUBS 0.006419f
C665 B.n598 VSUBS 0.006419f
C666 B.n599 VSUBS 0.006419f
C667 B.n600 VSUBS 0.006419f
C668 B.n601 VSUBS 0.006419f
C669 B.n602 VSUBS 0.006419f
C670 B.n603 VSUBS 0.006419f
C671 B.n604 VSUBS 0.006419f
C672 B.n605 VSUBS 0.006419f
C673 B.n606 VSUBS 0.006419f
C674 B.n607 VSUBS 0.006419f
C675 B.n608 VSUBS 0.006419f
C676 B.n609 VSUBS 0.006419f
C677 B.n610 VSUBS 0.006419f
C678 B.n611 VSUBS 0.006419f
C679 B.n612 VSUBS 0.006419f
C680 B.n613 VSUBS 0.006419f
C681 B.n614 VSUBS 0.006419f
C682 B.n615 VSUBS 0.006419f
C683 B.n616 VSUBS 0.006419f
C684 B.n617 VSUBS 0.006419f
C685 B.n618 VSUBS 0.006419f
C686 B.n619 VSUBS 0.006419f
C687 B.n620 VSUBS 0.006419f
C688 B.n621 VSUBS 0.006419f
C689 B.n622 VSUBS 0.006419f
C690 B.n623 VSUBS 0.006419f
C691 B.n624 VSUBS 0.006419f
C692 B.n625 VSUBS 0.006419f
C693 B.n626 VSUBS 0.006419f
C694 B.n627 VSUBS 0.006419f
C695 B.n628 VSUBS 0.006419f
C696 B.n629 VSUBS 0.006419f
C697 B.n630 VSUBS 0.006419f
C698 B.n631 VSUBS 0.006419f
C699 B.n632 VSUBS 0.006419f
C700 B.n633 VSUBS 0.006419f
C701 B.n634 VSUBS 0.006419f
C702 B.n635 VSUBS 0.006419f
C703 B.n636 VSUBS 0.006419f
C704 B.n637 VSUBS 0.006419f
C705 B.n638 VSUBS 0.006419f
C706 B.n639 VSUBS 0.006419f
C707 B.n640 VSUBS 0.006419f
C708 B.n641 VSUBS 0.006419f
C709 B.n642 VSUBS 0.006419f
C710 B.n643 VSUBS 0.006419f
C711 B.n644 VSUBS 0.006419f
C712 B.n645 VSUBS 0.006419f
C713 B.n646 VSUBS 0.006419f
C714 B.n647 VSUBS 0.006419f
C715 B.n648 VSUBS 0.006419f
C716 B.n649 VSUBS 0.006419f
C717 B.n650 VSUBS 0.006419f
C718 B.n651 VSUBS 0.006419f
C719 B.n652 VSUBS 0.006419f
C720 B.n653 VSUBS 0.006419f
C721 B.n654 VSUBS 0.006419f
C722 B.n655 VSUBS 0.006419f
C723 B.n656 VSUBS 0.006419f
C724 B.n657 VSUBS 0.006419f
C725 B.n658 VSUBS 0.006419f
C726 B.n659 VSUBS 0.006419f
C727 B.n660 VSUBS 0.006419f
C728 B.n661 VSUBS 0.006419f
C729 B.n662 VSUBS 0.006419f
C730 B.n663 VSUBS 0.006419f
C731 B.n664 VSUBS 0.006419f
C732 B.n665 VSUBS 0.006419f
C733 B.n666 VSUBS 0.006419f
C734 B.n667 VSUBS 0.016078f
C735 B.n668 VSUBS 0.016078f
C736 B.n669 VSUBS 0.015262f
C737 B.n670 VSUBS 0.006419f
C738 B.n671 VSUBS 0.006419f
C739 B.n672 VSUBS 0.006419f
C740 B.n673 VSUBS 0.006419f
C741 B.n674 VSUBS 0.006419f
C742 B.n675 VSUBS 0.006419f
C743 B.n676 VSUBS 0.006419f
C744 B.n677 VSUBS 0.006419f
C745 B.n678 VSUBS 0.006419f
C746 B.n679 VSUBS 0.006419f
C747 B.n680 VSUBS 0.006419f
C748 B.n681 VSUBS 0.006419f
C749 B.n682 VSUBS 0.006419f
C750 B.n683 VSUBS 0.006419f
C751 B.n684 VSUBS 0.006419f
C752 B.n685 VSUBS 0.006419f
C753 B.n686 VSUBS 0.006419f
C754 B.n687 VSUBS 0.006419f
C755 B.n688 VSUBS 0.006419f
C756 B.n689 VSUBS 0.006419f
C757 B.n690 VSUBS 0.006419f
C758 B.n691 VSUBS 0.006419f
C759 B.n692 VSUBS 0.006419f
C760 B.n693 VSUBS 0.006419f
C761 B.n694 VSUBS 0.006419f
C762 B.n695 VSUBS 0.006419f
C763 B.n696 VSUBS 0.006419f
C764 B.n697 VSUBS 0.006419f
C765 B.n698 VSUBS 0.006419f
C766 B.n699 VSUBS 0.006419f
C767 B.n700 VSUBS 0.006419f
C768 B.n701 VSUBS 0.006419f
C769 B.n702 VSUBS 0.006419f
C770 B.n703 VSUBS 0.006419f
C771 B.n704 VSUBS 0.006419f
C772 B.n705 VSUBS 0.006419f
C773 B.n706 VSUBS 0.006419f
C774 B.n707 VSUBS 0.006419f
C775 B.n708 VSUBS 0.006419f
C776 B.n709 VSUBS 0.006419f
C777 B.n710 VSUBS 0.006419f
C778 B.n711 VSUBS 0.006419f
C779 B.n712 VSUBS 0.006419f
C780 B.n713 VSUBS 0.006419f
C781 B.n714 VSUBS 0.006419f
C782 B.n715 VSUBS 0.006419f
C783 B.n716 VSUBS 0.006419f
C784 B.n717 VSUBS 0.006419f
C785 B.n718 VSUBS 0.006419f
C786 B.n719 VSUBS 0.014535f
C787 VTAIL.n0 VSUBS 0.026f
C788 VTAIL.n1 VSUBS 0.022868f
C789 VTAIL.n2 VSUBS 0.012288f
C790 VTAIL.n3 VSUBS 0.029045f
C791 VTAIL.n4 VSUBS 0.013011f
C792 VTAIL.n5 VSUBS 0.022868f
C793 VTAIL.n6 VSUBS 0.012288f
C794 VTAIL.n7 VSUBS 0.029045f
C795 VTAIL.n8 VSUBS 0.013011f
C796 VTAIL.n9 VSUBS 0.022868f
C797 VTAIL.n10 VSUBS 0.012288f
C798 VTAIL.n11 VSUBS 0.029045f
C799 VTAIL.n12 VSUBS 0.013011f
C800 VTAIL.n13 VSUBS 0.022868f
C801 VTAIL.n14 VSUBS 0.012288f
C802 VTAIL.n15 VSUBS 0.029045f
C803 VTAIL.n16 VSUBS 0.013011f
C804 VTAIL.n17 VSUBS 0.022868f
C805 VTAIL.n18 VSUBS 0.012288f
C806 VTAIL.n19 VSUBS 0.029045f
C807 VTAIL.n20 VSUBS 0.013011f
C808 VTAIL.n21 VSUBS 0.022868f
C809 VTAIL.n22 VSUBS 0.012288f
C810 VTAIL.n23 VSUBS 0.029045f
C811 VTAIL.n24 VSUBS 0.013011f
C812 VTAIL.n25 VSUBS 0.210493f
C813 VTAIL.t4 VSUBS 0.062812f
C814 VTAIL.n26 VSUBS 0.021783f
C815 VTAIL.n27 VSUBS 0.021849f
C816 VTAIL.n28 VSUBS 0.012288f
C817 VTAIL.n29 VSUBS 1.41815f
C818 VTAIL.n30 VSUBS 0.022868f
C819 VTAIL.n31 VSUBS 0.012288f
C820 VTAIL.n32 VSUBS 0.013011f
C821 VTAIL.n33 VSUBS 0.029045f
C822 VTAIL.n34 VSUBS 0.029045f
C823 VTAIL.n35 VSUBS 0.013011f
C824 VTAIL.n36 VSUBS 0.012288f
C825 VTAIL.n37 VSUBS 0.022868f
C826 VTAIL.n38 VSUBS 0.022868f
C827 VTAIL.n39 VSUBS 0.012288f
C828 VTAIL.n40 VSUBS 0.013011f
C829 VTAIL.n41 VSUBS 0.029045f
C830 VTAIL.n42 VSUBS 0.029045f
C831 VTAIL.n43 VSUBS 0.029045f
C832 VTAIL.n44 VSUBS 0.013011f
C833 VTAIL.n45 VSUBS 0.012288f
C834 VTAIL.n46 VSUBS 0.022868f
C835 VTAIL.n47 VSUBS 0.022868f
C836 VTAIL.n48 VSUBS 0.012288f
C837 VTAIL.n49 VSUBS 0.012649f
C838 VTAIL.n50 VSUBS 0.012649f
C839 VTAIL.n51 VSUBS 0.029045f
C840 VTAIL.n52 VSUBS 0.029045f
C841 VTAIL.n53 VSUBS 0.013011f
C842 VTAIL.n54 VSUBS 0.012288f
C843 VTAIL.n55 VSUBS 0.022868f
C844 VTAIL.n56 VSUBS 0.022868f
C845 VTAIL.n57 VSUBS 0.012288f
C846 VTAIL.n58 VSUBS 0.013011f
C847 VTAIL.n59 VSUBS 0.029045f
C848 VTAIL.n60 VSUBS 0.029045f
C849 VTAIL.n61 VSUBS 0.013011f
C850 VTAIL.n62 VSUBS 0.012288f
C851 VTAIL.n63 VSUBS 0.022868f
C852 VTAIL.n64 VSUBS 0.022868f
C853 VTAIL.n65 VSUBS 0.012288f
C854 VTAIL.n66 VSUBS 0.013011f
C855 VTAIL.n67 VSUBS 0.029045f
C856 VTAIL.n68 VSUBS 0.029045f
C857 VTAIL.n69 VSUBS 0.013011f
C858 VTAIL.n70 VSUBS 0.012288f
C859 VTAIL.n71 VSUBS 0.022868f
C860 VTAIL.n72 VSUBS 0.022868f
C861 VTAIL.n73 VSUBS 0.012288f
C862 VTAIL.n74 VSUBS 0.013011f
C863 VTAIL.n75 VSUBS 0.029045f
C864 VTAIL.n76 VSUBS 0.07329f
C865 VTAIL.n77 VSUBS 0.013011f
C866 VTAIL.n78 VSUBS 0.012288f
C867 VTAIL.n79 VSUBS 0.050983f
C868 VTAIL.n80 VSUBS 0.03693f
C869 VTAIL.n81 VSUBS 0.147581f
C870 VTAIL.n82 VSUBS 0.026f
C871 VTAIL.n83 VSUBS 0.022868f
C872 VTAIL.n84 VSUBS 0.012288f
C873 VTAIL.n85 VSUBS 0.029045f
C874 VTAIL.n86 VSUBS 0.013011f
C875 VTAIL.n87 VSUBS 0.022868f
C876 VTAIL.n88 VSUBS 0.012288f
C877 VTAIL.n89 VSUBS 0.029045f
C878 VTAIL.n90 VSUBS 0.013011f
C879 VTAIL.n91 VSUBS 0.022868f
C880 VTAIL.n92 VSUBS 0.012288f
C881 VTAIL.n93 VSUBS 0.029045f
C882 VTAIL.n94 VSUBS 0.013011f
C883 VTAIL.n95 VSUBS 0.022868f
C884 VTAIL.n96 VSUBS 0.012288f
C885 VTAIL.n97 VSUBS 0.029045f
C886 VTAIL.n98 VSUBS 0.013011f
C887 VTAIL.n99 VSUBS 0.022868f
C888 VTAIL.n100 VSUBS 0.012288f
C889 VTAIL.n101 VSUBS 0.029045f
C890 VTAIL.n102 VSUBS 0.013011f
C891 VTAIL.n103 VSUBS 0.022868f
C892 VTAIL.n104 VSUBS 0.012288f
C893 VTAIL.n105 VSUBS 0.029045f
C894 VTAIL.n106 VSUBS 0.013011f
C895 VTAIL.n107 VSUBS 0.210493f
C896 VTAIL.t0 VSUBS 0.062812f
C897 VTAIL.n108 VSUBS 0.021783f
C898 VTAIL.n109 VSUBS 0.021849f
C899 VTAIL.n110 VSUBS 0.012288f
C900 VTAIL.n111 VSUBS 1.41815f
C901 VTAIL.n112 VSUBS 0.022868f
C902 VTAIL.n113 VSUBS 0.012288f
C903 VTAIL.n114 VSUBS 0.013011f
C904 VTAIL.n115 VSUBS 0.029045f
C905 VTAIL.n116 VSUBS 0.029045f
C906 VTAIL.n117 VSUBS 0.013011f
C907 VTAIL.n118 VSUBS 0.012288f
C908 VTAIL.n119 VSUBS 0.022868f
C909 VTAIL.n120 VSUBS 0.022868f
C910 VTAIL.n121 VSUBS 0.012288f
C911 VTAIL.n122 VSUBS 0.013011f
C912 VTAIL.n123 VSUBS 0.029045f
C913 VTAIL.n124 VSUBS 0.029045f
C914 VTAIL.n125 VSUBS 0.029045f
C915 VTAIL.n126 VSUBS 0.013011f
C916 VTAIL.n127 VSUBS 0.012288f
C917 VTAIL.n128 VSUBS 0.022868f
C918 VTAIL.n129 VSUBS 0.022868f
C919 VTAIL.n130 VSUBS 0.012288f
C920 VTAIL.n131 VSUBS 0.012649f
C921 VTAIL.n132 VSUBS 0.012649f
C922 VTAIL.n133 VSUBS 0.029045f
C923 VTAIL.n134 VSUBS 0.029045f
C924 VTAIL.n135 VSUBS 0.013011f
C925 VTAIL.n136 VSUBS 0.012288f
C926 VTAIL.n137 VSUBS 0.022868f
C927 VTAIL.n138 VSUBS 0.022868f
C928 VTAIL.n139 VSUBS 0.012288f
C929 VTAIL.n140 VSUBS 0.013011f
C930 VTAIL.n141 VSUBS 0.029045f
C931 VTAIL.n142 VSUBS 0.029045f
C932 VTAIL.n143 VSUBS 0.013011f
C933 VTAIL.n144 VSUBS 0.012288f
C934 VTAIL.n145 VSUBS 0.022868f
C935 VTAIL.n146 VSUBS 0.022868f
C936 VTAIL.n147 VSUBS 0.012288f
C937 VTAIL.n148 VSUBS 0.013011f
C938 VTAIL.n149 VSUBS 0.029045f
C939 VTAIL.n150 VSUBS 0.029045f
C940 VTAIL.n151 VSUBS 0.013011f
C941 VTAIL.n152 VSUBS 0.012288f
C942 VTAIL.n153 VSUBS 0.022868f
C943 VTAIL.n154 VSUBS 0.022868f
C944 VTAIL.n155 VSUBS 0.012288f
C945 VTAIL.n156 VSUBS 0.013011f
C946 VTAIL.n157 VSUBS 0.029045f
C947 VTAIL.n158 VSUBS 0.07329f
C948 VTAIL.n159 VSUBS 0.013011f
C949 VTAIL.n160 VSUBS 0.012288f
C950 VTAIL.n161 VSUBS 0.050983f
C951 VTAIL.n162 VSUBS 0.03693f
C952 VTAIL.n163 VSUBS 0.233493f
C953 VTAIL.n164 VSUBS 0.026f
C954 VTAIL.n165 VSUBS 0.022868f
C955 VTAIL.n166 VSUBS 0.012288f
C956 VTAIL.n167 VSUBS 0.029045f
C957 VTAIL.n168 VSUBS 0.013011f
C958 VTAIL.n169 VSUBS 0.022868f
C959 VTAIL.n170 VSUBS 0.012288f
C960 VTAIL.n171 VSUBS 0.029045f
C961 VTAIL.n172 VSUBS 0.013011f
C962 VTAIL.n173 VSUBS 0.022868f
C963 VTAIL.n174 VSUBS 0.012288f
C964 VTAIL.n175 VSUBS 0.029045f
C965 VTAIL.n176 VSUBS 0.013011f
C966 VTAIL.n177 VSUBS 0.022868f
C967 VTAIL.n178 VSUBS 0.012288f
C968 VTAIL.n179 VSUBS 0.029045f
C969 VTAIL.n180 VSUBS 0.013011f
C970 VTAIL.n181 VSUBS 0.022868f
C971 VTAIL.n182 VSUBS 0.012288f
C972 VTAIL.n183 VSUBS 0.029045f
C973 VTAIL.n184 VSUBS 0.013011f
C974 VTAIL.n185 VSUBS 0.022868f
C975 VTAIL.n186 VSUBS 0.012288f
C976 VTAIL.n187 VSUBS 0.029045f
C977 VTAIL.n188 VSUBS 0.013011f
C978 VTAIL.n189 VSUBS 0.210493f
C979 VTAIL.t3 VSUBS 0.062812f
C980 VTAIL.n190 VSUBS 0.021783f
C981 VTAIL.n191 VSUBS 0.021849f
C982 VTAIL.n192 VSUBS 0.012288f
C983 VTAIL.n193 VSUBS 1.41815f
C984 VTAIL.n194 VSUBS 0.022868f
C985 VTAIL.n195 VSUBS 0.012288f
C986 VTAIL.n196 VSUBS 0.013011f
C987 VTAIL.n197 VSUBS 0.029045f
C988 VTAIL.n198 VSUBS 0.029045f
C989 VTAIL.n199 VSUBS 0.013011f
C990 VTAIL.n200 VSUBS 0.012288f
C991 VTAIL.n201 VSUBS 0.022868f
C992 VTAIL.n202 VSUBS 0.022868f
C993 VTAIL.n203 VSUBS 0.012288f
C994 VTAIL.n204 VSUBS 0.013011f
C995 VTAIL.n205 VSUBS 0.029045f
C996 VTAIL.n206 VSUBS 0.029045f
C997 VTAIL.n207 VSUBS 0.029045f
C998 VTAIL.n208 VSUBS 0.013011f
C999 VTAIL.n209 VSUBS 0.012288f
C1000 VTAIL.n210 VSUBS 0.022868f
C1001 VTAIL.n211 VSUBS 0.022868f
C1002 VTAIL.n212 VSUBS 0.012288f
C1003 VTAIL.n213 VSUBS 0.012649f
C1004 VTAIL.n214 VSUBS 0.012649f
C1005 VTAIL.n215 VSUBS 0.029045f
C1006 VTAIL.n216 VSUBS 0.029045f
C1007 VTAIL.n217 VSUBS 0.013011f
C1008 VTAIL.n218 VSUBS 0.012288f
C1009 VTAIL.n219 VSUBS 0.022868f
C1010 VTAIL.n220 VSUBS 0.022868f
C1011 VTAIL.n221 VSUBS 0.012288f
C1012 VTAIL.n222 VSUBS 0.013011f
C1013 VTAIL.n223 VSUBS 0.029045f
C1014 VTAIL.n224 VSUBS 0.029045f
C1015 VTAIL.n225 VSUBS 0.013011f
C1016 VTAIL.n226 VSUBS 0.012288f
C1017 VTAIL.n227 VSUBS 0.022868f
C1018 VTAIL.n228 VSUBS 0.022868f
C1019 VTAIL.n229 VSUBS 0.012288f
C1020 VTAIL.n230 VSUBS 0.013011f
C1021 VTAIL.n231 VSUBS 0.029045f
C1022 VTAIL.n232 VSUBS 0.029045f
C1023 VTAIL.n233 VSUBS 0.013011f
C1024 VTAIL.n234 VSUBS 0.012288f
C1025 VTAIL.n235 VSUBS 0.022868f
C1026 VTAIL.n236 VSUBS 0.022868f
C1027 VTAIL.n237 VSUBS 0.012288f
C1028 VTAIL.n238 VSUBS 0.013011f
C1029 VTAIL.n239 VSUBS 0.029045f
C1030 VTAIL.n240 VSUBS 0.07329f
C1031 VTAIL.n241 VSUBS 0.013011f
C1032 VTAIL.n242 VSUBS 0.012288f
C1033 VTAIL.n243 VSUBS 0.050983f
C1034 VTAIL.n244 VSUBS 0.03693f
C1035 VTAIL.n245 VSUBS 1.63891f
C1036 VTAIL.n246 VSUBS 0.026f
C1037 VTAIL.n247 VSUBS 0.022868f
C1038 VTAIL.n248 VSUBS 0.012288f
C1039 VTAIL.n249 VSUBS 0.029045f
C1040 VTAIL.n250 VSUBS 0.013011f
C1041 VTAIL.n251 VSUBS 0.022868f
C1042 VTAIL.n252 VSUBS 0.012288f
C1043 VTAIL.n253 VSUBS 0.029045f
C1044 VTAIL.n254 VSUBS 0.013011f
C1045 VTAIL.n255 VSUBS 0.022868f
C1046 VTAIL.n256 VSUBS 0.012288f
C1047 VTAIL.n257 VSUBS 0.029045f
C1048 VTAIL.n258 VSUBS 0.013011f
C1049 VTAIL.n259 VSUBS 0.022868f
C1050 VTAIL.n260 VSUBS 0.012288f
C1051 VTAIL.n261 VSUBS 0.029045f
C1052 VTAIL.n262 VSUBS 0.013011f
C1053 VTAIL.n263 VSUBS 0.022868f
C1054 VTAIL.n264 VSUBS 0.012288f
C1055 VTAIL.n265 VSUBS 0.029045f
C1056 VTAIL.n266 VSUBS 0.029045f
C1057 VTAIL.n267 VSUBS 0.013011f
C1058 VTAIL.n268 VSUBS 0.022868f
C1059 VTAIL.n269 VSUBS 0.012288f
C1060 VTAIL.n270 VSUBS 0.029045f
C1061 VTAIL.n271 VSUBS 0.013011f
C1062 VTAIL.n272 VSUBS 0.210493f
C1063 VTAIL.t7 VSUBS 0.062812f
C1064 VTAIL.n273 VSUBS 0.021783f
C1065 VTAIL.n274 VSUBS 0.021849f
C1066 VTAIL.n275 VSUBS 0.012288f
C1067 VTAIL.n276 VSUBS 1.41815f
C1068 VTAIL.n277 VSUBS 0.022868f
C1069 VTAIL.n278 VSUBS 0.012288f
C1070 VTAIL.n279 VSUBS 0.013011f
C1071 VTAIL.n280 VSUBS 0.029045f
C1072 VTAIL.n281 VSUBS 0.029045f
C1073 VTAIL.n282 VSUBS 0.013011f
C1074 VTAIL.n283 VSUBS 0.012288f
C1075 VTAIL.n284 VSUBS 0.022868f
C1076 VTAIL.n285 VSUBS 0.022868f
C1077 VTAIL.n286 VSUBS 0.012288f
C1078 VTAIL.n287 VSUBS 0.013011f
C1079 VTAIL.n288 VSUBS 0.029045f
C1080 VTAIL.n289 VSUBS 0.029045f
C1081 VTAIL.n290 VSUBS 0.013011f
C1082 VTAIL.n291 VSUBS 0.012288f
C1083 VTAIL.n292 VSUBS 0.022868f
C1084 VTAIL.n293 VSUBS 0.022868f
C1085 VTAIL.n294 VSUBS 0.012288f
C1086 VTAIL.n295 VSUBS 0.012649f
C1087 VTAIL.n296 VSUBS 0.012649f
C1088 VTAIL.n297 VSUBS 0.029045f
C1089 VTAIL.n298 VSUBS 0.029045f
C1090 VTAIL.n299 VSUBS 0.013011f
C1091 VTAIL.n300 VSUBS 0.012288f
C1092 VTAIL.n301 VSUBS 0.022868f
C1093 VTAIL.n302 VSUBS 0.022868f
C1094 VTAIL.n303 VSUBS 0.012288f
C1095 VTAIL.n304 VSUBS 0.013011f
C1096 VTAIL.n305 VSUBS 0.029045f
C1097 VTAIL.n306 VSUBS 0.029045f
C1098 VTAIL.n307 VSUBS 0.013011f
C1099 VTAIL.n308 VSUBS 0.012288f
C1100 VTAIL.n309 VSUBS 0.022868f
C1101 VTAIL.n310 VSUBS 0.022868f
C1102 VTAIL.n311 VSUBS 0.012288f
C1103 VTAIL.n312 VSUBS 0.013011f
C1104 VTAIL.n313 VSUBS 0.029045f
C1105 VTAIL.n314 VSUBS 0.029045f
C1106 VTAIL.n315 VSUBS 0.013011f
C1107 VTAIL.n316 VSUBS 0.012288f
C1108 VTAIL.n317 VSUBS 0.022868f
C1109 VTAIL.n318 VSUBS 0.022868f
C1110 VTAIL.n319 VSUBS 0.012288f
C1111 VTAIL.n320 VSUBS 0.013011f
C1112 VTAIL.n321 VSUBS 0.029045f
C1113 VTAIL.n322 VSUBS 0.07329f
C1114 VTAIL.n323 VSUBS 0.013011f
C1115 VTAIL.n324 VSUBS 0.012288f
C1116 VTAIL.n325 VSUBS 0.050983f
C1117 VTAIL.n326 VSUBS 0.03693f
C1118 VTAIL.n327 VSUBS 1.63891f
C1119 VTAIL.n328 VSUBS 0.026f
C1120 VTAIL.n329 VSUBS 0.022868f
C1121 VTAIL.n330 VSUBS 0.012288f
C1122 VTAIL.n331 VSUBS 0.029045f
C1123 VTAIL.n332 VSUBS 0.013011f
C1124 VTAIL.n333 VSUBS 0.022868f
C1125 VTAIL.n334 VSUBS 0.012288f
C1126 VTAIL.n335 VSUBS 0.029045f
C1127 VTAIL.n336 VSUBS 0.013011f
C1128 VTAIL.n337 VSUBS 0.022868f
C1129 VTAIL.n338 VSUBS 0.012288f
C1130 VTAIL.n339 VSUBS 0.029045f
C1131 VTAIL.n340 VSUBS 0.013011f
C1132 VTAIL.n341 VSUBS 0.022868f
C1133 VTAIL.n342 VSUBS 0.012288f
C1134 VTAIL.n343 VSUBS 0.029045f
C1135 VTAIL.n344 VSUBS 0.013011f
C1136 VTAIL.n345 VSUBS 0.022868f
C1137 VTAIL.n346 VSUBS 0.012288f
C1138 VTAIL.n347 VSUBS 0.029045f
C1139 VTAIL.n348 VSUBS 0.029045f
C1140 VTAIL.n349 VSUBS 0.013011f
C1141 VTAIL.n350 VSUBS 0.022868f
C1142 VTAIL.n351 VSUBS 0.012288f
C1143 VTAIL.n352 VSUBS 0.029045f
C1144 VTAIL.n353 VSUBS 0.013011f
C1145 VTAIL.n354 VSUBS 0.210493f
C1146 VTAIL.t6 VSUBS 0.062812f
C1147 VTAIL.n355 VSUBS 0.021783f
C1148 VTAIL.n356 VSUBS 0.021849f
C1149 VTAIL.n357 VSUBS 0.012288f
C1150 VTAIL.n358 VSUBS 1.41815f
C1151 VTAIL.n359 VSUBS 0.022868f
C1152 VTAIL.n360 VSUBS 0.012288f
C1153 VTAIL.n361 VSUBS 0.013011f
C1154 VTAIL.n362 VSUBS 0.029045f
C1155 VTAIL.n363 VSUBS 0.029045f
C1156 VTAIL.n364 VSUBS 0.013011f
C1157 VTAIL.n365 VSUBS 0.012288f
C1158 VTAIL.n366 VSUBS 0.022868f
C1159 VTAIL.n367 VSUBS 0.022868f
C1160 VTAIL.n368 VSUBS 0.012288f
C1161 VTAIL.n369 VSUBS 0.013011f
C1162 VTAIL.n370 VSUBS 0.029045f
C1163 VTAIL.n371 VSUBS 0.029045f
C1164 VTAIL.n372 VSUBS 0.013011f
C1165 VTAIL.n373 VSUBS 0.012288f
C1166 VTAIL.n374 VSUBS 0.022868f
C1167 VTAIL.n375 VSUBS 0.022868f
C1168 VTAIL.n376 VSUBS 0.012288f
C1169 VTAIL.n377 VSUBS 0.012649f
C1170 VTAIL.n378 VSUBS 0.012649f
C1171 VTAIL.n379 VSUBS 0.029045f
C1172 VTAIL.n380 VSUBS 0.029045f
C1173 VTAIL.n381 VSUBS 0.013011f
C1174 VTAIL.n382 VSUBS 0.012288f
C1175 VTAIL.n383 VSUBS 0.022868f
C1176 VTAIL.n384 VSUBS 0.022868f
C1177 VTAIL.n385 VSUBS 0.012288f
C1178 VTAIL.n386 VSUBS 0.013011f
C1179 VTAIL.n387 VSUBS 0.029045f
C1180 VTAIL.n388 VSUBS 0.029045f
C1181 VTAIL.n389 VSUBS 0.013011f
C1182 VTAIL.n390 VSUBS 0.012288f
C1183 VTAIL.n391 VSUBS 0.022868f
C1184 VTAIL.n392 VSUBS 0.022868f
C1185 VTAIL.n393 VSUBS 0.012288f
C1186 VTAIL.n394 VSUBS 0.013011f
C1187 VTAIL.n395 VSUBS 0.029045f
C1188 VTAIL.n396 VSUBS 0.029045f
C1189 VTAIL.n397 VSUBS 0.013011f
C1190 VTAIL.n398 VSUBS 0.012288f
C1191 VTAIL.n399 VSUBS 0.022868f
C1192 VTAIL.n400 VSUBS 0.022868f
C1193 VTAIL.n401 VSUBS 0.012288f
C1194 VTAIL.n402 VSUBS 0.013011f
C1195 VTAIL.n403 VSUBS 0.029045f
C1196 VTAIL.n404 VSUBS 0.07329f
C1197 VTAIL.n405 VSUBS 0.013011f
C1198 VTAIL.n406 VSUBS 0.012288f
C1199 VTAIL.n407 VSUBS 0.050983f
C1200 VTAIL.n408 VSUBS 0.03693f
C1201 VTAIL.n409 VSUBS 0.233493f
C1202 VTAIL.n410 VSUBS 0.026f
C1203 VTAIL.n411 VSUBS 0.022868f
C1204 VTAIL.n412 VSUBS 0.012288f
C1205 VTAIL.n413 VSUBS 0.029045f
C1206 VTAIL.n414 VSUBS 0.013011f
C1207 VTAIL.n415 VSUBS 0.022868f
C1208 VTAIL.n416 VSUBS 0.012288f
C1209 VTAIL.n417 VSUBS 0.029045f
C1210 VTAIL.n418 VSUBS 0.013011f
C1211 VTAIL.n419 VSUBS 0.022868f
C1212 VTAIL.n420 VSUBS 0.012288f
C1213 VTAIL.n421 VSUBS 0.029045f
C1214 VTAIL.n422 VSUBS 0.013011f
C1215 VTAIL.n423 VSUBS 0.022868f
C1216 VTAIL.n424 VSUBS 0.012288f
C1217 VTAIL.n425 VSUBS 0.029045f
C1218 VTAIL.n426 VSUBS 0.013011f
C1219 VTAIL.n427 VSUBS 0.022868f
C1220 VTAIL.n428 VSUBS 0.012288f
C1221 VTAIL.n429 VSUBS 0.029045f
C1222 VTAIL.n430 VSUBS 0.029045f
C1223 VTAIL.n431 VSUBS 0.013011f
C1224 VTAIL.n432 VSUBS 0.022868f
C1225 VTAIL.n433 VSUBS 0.012288f
C1226 VTAIL.n434 VSUBS 0.029045f
C1227 VTAIL.n435 VSUBS 0.013011f
C1228 VTAIL.n436 VSUBS 0.210493f
C1229 VTAIL.t2 VSUBS 0.062812f
C1230 VTAIL.n437 VSUBS 0.021783f
C1231 VTAIL.n438 VSUBS 0.021849f
C1232 VTAIL.n439 VSUBS 0.012288f
C1233 VTAIL.n440 VSUBS 1.41815f
C1234 VTAIL.n441 VSUBS 0.022868f
C1235 VTAIL.n442 VSUBS 0.012288f
C1236 VTAIL.n443 VSUBS 0.013011f
C1237 VTAIL.n444 VSUBS 0.029045f
C1238 VTAIL.n445 VSUBS 0.029045f
C1239 VTAIL.n446 VSUBS 0.013011f
C1240 VTAIL.n447 VSUBS 0.012288f
C1241 VTAIL.n448 VSUBS 0.022868f
C1242 VTAIL.n449 VSUBS 0.022868f
C1243 VTAIL.n450 VSUBS 0.012288f
C1244 VTAIL.n451 VSUBS 0.013011f
C1245 VTAIL.n452 VSUBS 0.029045f
C1246 VTAIL.n453 VSUBS 0.029045f
C1247 VTAIL.n454 VSUBS 0.013011f
C1248 VTAIL.n455 VSUBS 0.012288f
C1249 VTAIL.n456 VSUBS 0.022868f
C1250 VTAIL.n457 VSUBS 0.022868f
C1251 VTAIL.n458 VSUBS 0.012288f
C1252 VTAIL.n459 VSUBS 0.012649f
C1253 VTAIL.n460 VSUBS 0.012649f
C1254 VTAIL.n461 VSUBS 0.029045f
C1255 VTAIL.n462 VSUBS 0.029045f
C1256 VTAIL.n463 VSUBS 0.013011f
C1257 VTAIL.n464 VSUBS 0.012288f
C1258 VTAIL.n465 VSUBS 0.022868f
C1259 VTAIL.n466 VSUBS 0.022868f
C1260 VTAIL.n467 VSUBS 0.012288f
C1261 VTAIL.n468 VSUBS 0.013011f
C1262 VTAIL.n469 VSUBS 0.029045f
C1263 VTAIL.n470 VSUBS 0.029045f
C1264 VTAIL.n471 VSUBS 0.013011f
C1265 VTAIL.n472 VSUBS 0.012288f
C1266 VTAIL.n473 VSUBS 0.022868f
C1267 VTAIL.n474 VSUBS 0.022868f
C1268 VTAIL.n475 VSUBS 0.012288f
C1269 VTAIL.n476 VSUBS 0.013011f
C1270 VTAIL.n477 VSUBS 0.029045f
C1271 VTAIL.n478 VSUBS 0.029045f
C1272 VTAIL.n479 VSUBS 0.013011f
C1273 VTAIL.n480 VSUBS 0.012288f
C1274 VTAIL.n481 VSUBS 0.022868f
C1275 VTAIL.n482 VSUBS 0.022868f
C1276 VTAIL.n483 VSUBS 0.012288f
C1277 VTAIL.n484 VSUBS 0.013011f
C1278 VTAIL.n485 VSUBS 0.029045f
C1279 VTAIL.n486 VSUBS 0.07329f
C1280 VTAIL.n487 VSUBS 0.013011f
C1281 VTAIL.n488 VSUBS 0.012288f
C1282 VTAIL.n489 VSUBS 0.050983f
C1283 VTAIL.n490 VSUBS 0.03693f
C1284 VTAIL.n491 VSUBS 0.233493f
C1285 VTAIL.n492 VSUBS 0.026f
C1286 VTAIL.n493 VSUBS 0.022868f
C1287 VTAIL.n494 VSUBS 0.012288f
C1288 VTAIL.n495 VSUBS 0.029045f
C1289 VTAIL.n496 VSUBS 0.013011f
C1290 VTAIL.n497 VSUBS 0.022868f
C1291 VTAIL.n498 VSUBS 0.012288f
C1292 VTAIL.n499 VSUBS 0.029045f
C1293 VTAIL.n500 VSUBS 0.013011f
C1294 VTAIL.n501 VSUBS 0.022868f
C1295 VTAIL.n502 VSUBS 0.012288f
C1296 VTAIL.n503 VSUBS 0.029045f
C1297 VTAIL.n504 VSUBS 0.013011f
C1298 VTAIL.n505 VSUBS 0.022868f
C1299 VTAIL.n506 VSUBS 0.012288f
C1300 VTAIL.n507 VSUBS 0.029045f
C1301 VTAIL.n508 VSUBS 0.013011f
C1302 VTAIL.n509 VSUBS 0.022868f
C1303 VTAIL.n510 VSUBS 0.012288f
C1304 VTAIL.n511 VSUBS 0.029045f
C1305 VTAIL.n512 VSUBS 0.029045f
C1306 VTAIL.n513 VSUBS 0.013011f
C1307 VTAIL.n514 VSUBS 0.022868f
C1308 VTAIL.n515 VSUBS 0.012288f
C1309 VTAIL.n516 VSUBS 0.029045f
C1310 VTAIL.n517 VSUBS 0.013011f
C1311 VTAIL.n518 VSUBS 0.210493f
C1312 VTAIL.t1 VSUBS 0.062812f
C1313 VTAIL.n519 VSUBS 0.021783f
C1314 VTAIL.n520 VSUBS 0.021849f
C1315 VTAIL.n521 VSUBS 0.012288f
C1316 VTAIL.n522 VSUBS 1.41815f
C1317 VTAIL.n523 VSUBS 0.022868f
C1318 VTAIL.n524 VSUBS 0.012288f
C1319 VTAIL.n525 VSUBS 0.013011f
C1320 VTAIL.n526 VSUBS 0.029045f
C1321 VTAIL.n527 VSUBS 0.029045f
C1322 VTAIL.n528 VSUBS 0.013011f
C1323 VTAIL.n529 VSUBS 0.012288f
C1324 VTAIL.n530 VSUBS 0.022868f
C1325 VTAIL.n531 VSUBS 0.022868f
C1326 VTAIL.n532 VSUBS 0.012288f
C1327 VTAIL.n533 VSUBS 0.013011f
C1328 VTAIL.n534 VSUBS 0.029045f
C1329 VTAIL.n535 VSUBS 0.029045f
C1330 VTAIL.n536 VSUBS 0.013011f
C1331 VTAIL.n537 VSUBS 0.012288f
C1332 VTAIL.n538 VSUBS 0.022868f
C1333 VTAIL.n539 VSUBS 0.022868f
C1334 VTAIL.n540 VSUBS 0.012288f
C1335 VTAIL.n541 VSUBS 0.012649f
C1336 VTAIL.n542 VSUBS 0.012649f
C1337 VTAIL.n543 VSUBS 0.029045f
C1338 VTAIL.n544 VSUBS 0.029045f
C1339 VTAIL.n545 VSUBS 0.013011f
C1340 VTAIL.n546 VSUBS 0.012288f
C1341 VTAIL.n547 VSUBS 0.022868f
C1342 VTAIL.n548 VSUBS 0.022868f
C1343 VTAIL.n549 VSUBS 0.012288f
C1344 VTAIL.n550 VSUBS 0.013011f
C1345 VTAIL.n551 VSUBS 0.029045f
C1346 VTAIL.n552 VSUBS 0.029045f
C1347 VTAIL.n553 VSUBS 0.013011f
C1348 VTAIL.n554 VSUBS 0.012288f
C1349 VTAIL.n555 VSUBS 0.022868f
C1350 VTAIL.n556 VSUBS 0.022868f
C1351 VTAIL.n557 VSUBS 0.012288f
C1352 VTAIL.n558 VSUBS 0.013011f
C1353 VTAIL.n559 VSUBS 0.029045f
C1354 VTAIL.n560 VSUBS 0.029045f
C1355 VTAIL.n561 VSUBS 0.013011f
C1356 VTAIL.n562 VSUBS 0.012288f
C1357 VTAIL.n563 VSUBS 0.022868f
C1358 VTAIL.n564 VSUBS 0.022868f
C1359 VTAIL.n565 VSUBS 0.012288f
C1360 VTAIL.n566 VSUBS 0.013011f
C1361 VTAIL.n567 VSUBS 0.029045f
C1362 VTAIL.n568 VSUBS 0.07329f
C1363 VTAIL.n569 VSUBS 0.013011f
C1364 VTAIL.n570 VSUBS 0.012288f
C1365 VTAIL.n571 VSUBS 0.050983f
C1366 VTAIL.n572 VSUBS 0.03693f
C1367 VTAIL.n573 VSUBS 1.63891f
C1368 VTAIL.n574 VSUBS 0.026f
C1369 VTAIL.n575 VSUBS 0.022868f
C1370 VTAIL.n576 VSUBS 0.012288f
C1371 VTAIL.n577 VSUBS 0.029045f
C1372 VTAIL.n578 VSUBS 0.013011f
C1373 VTAIL.n579 VSUBS 0.022868f
C1374 VTAIL.n580 VSUBS 0.012288f
C1375 VTAIL.n581 VSUBS 0.029045f
C1376 VTAIL.n582 VSUBS 0.013011f
C1377 VTAIL.n583 VSUBS 0.022868f
C1378 VTAIL.n584 VSUBS 0.012288f
C1379 VTAIL.n585 VSUBS 0.029045f
C1380 VTAIL.n586 VSUBS 0.013011f
C1381 VTAIL.n587 VSUBS 0.022868f
C1382 VTAIL.n588 VSUBS 0.012288f
C1383 VTAIL.n589 VSUBS 0.029045f
C1384 VTAIL.n590 VSUBS 0.013011f
C1385 VTAIL.n591 VSUBS 0.022868f
C1386 VTAIL.n592 VSUBS 0.012288f
C1387 VTAIL.n593 VSUBS 0.029045f
C1388 VTAIL.n594 VSUBS 0.013011f
C1389 VTAIL.n595 VSUBS 0.022868f
C1390 VTAIL.n596 VSUBS 0.012288f
C1391 VTAIL.n597 VSUBS 0.029045f
C1392 VTAIL.n598 VSUBS 0.013011f
C1393 VTAIL.n599 VSUBS 0.210493f
C1394 VTAIL.t5 VSUBS 0.062812f
C1395 VTAIL.n600 VSUBS 0.021783f
C1396 VTAIL.n601 VSUBS 0.021849f
C1397 VTAIL.n602 VSUBS 0.012288f
C1398 VTAIL.n603 VSUBS 1.41815f
C1399 VTAIL.n604 VSUBS 0.022868f
C1400 VTAIL.n605 VSUBS 0.012288f
C1401 VTAIL.n606 VSUBS 0.013011f
C1402 VTAIL.n607 VSUBS 0.029045f
C1403 VTAIL.n608 VSUBS 0.029045f
C1404 VTAIL.n609 VSUBS 0.013011f
C1405 VTAIL.n610 VSUBS 0.012288f
C1406 VTAIL.n611 VSUBS 0.022868f
C1407 VTAIL.n612 VSUBS 0.022868f
C1408 VTAIL.n613 VSUBS 0.012288f
C1409 VTAIL.n614 VSUBS 0.013011f
C1410 VTAIL.n615 VSUBS 0.029045f
C1411 VTAIL.n616 VSUBS 0.029045f
C1412 VTAIL.n617 VSUBS 0.029045f
C1413 VTAIL.n618 VSUBS 0.013011f
C1414 VTAIL.n619 VSUBS 0.012288f
C1415 VTAIL.n620 VSUBS 0.022868f
C1416 VTAIL.n621 VSUBS 0.022868f
C1417 VTAIL.n622 VSUBS 0.012288f
C1418 VTAIL.n623 VSUBS 0.012649f
C1419 VTAIL.n624 VSUBS 0.012649f
C1420 VTAIL.n625 VSUBS 0.029045f
C1421 VTAIL.n626 VSUBS 0.029045f
C1422 VTAIL.n627 VSUBS 0.013011f
C1423 VTAIL.n628 VSUBS 0.012288f
C1424 VTAIL.n629 VSUBS 0.022868f
C1425 VTAIL.n630 VSUBS 0.022868f
C1426 VTAIL.n631 VSUBS 0.012288f
C1427 VTAIL.n632 VSUBS 0.013011f
C1428 VTAIL.n633 VSUBS 0.029045f
C1429 VTAIL.n634 VSUBS 0.029045f
C1430 VTAIL.n635 VSUBS 0.013011f
C1431 VTAIL.n636 VSUBS 0.012288f
C1432 VTAIL.n637 VSUBS 0.022868f
C1433 VTAIL.n638 VSUBS 0.022868f
C1434 VTAIL.n639 VSUBS 0.012288f
C1435 VTAIL.n640 VSUBS 0.013011f
C1436 VTAIL.n641 VSUBS 0.029045f
C1437 VTAIL.n642 VSUBS 0.029045f
C1438 VTAIL.n643 VSUBS 0.013011f
C1439 VTAIL.n644 VSUBS 0.012288f
C1440 VTAIL.n645 VSUBS 0.022868f
C1441 VTAIL.n646 VSUBS 0.022868f
C1442 VTAIL.n647 VSUBS 0.012288f
C1443 VTAIL.n648 VSUBS 0.013011f
C1444 VTAIL.n649 VSUBS 0.029045f
C1445 VTAIL.n650 VSUBS 0.07329f
C1446 VTAIL.n651 VSUBS 0.013011f
C1447 VTAIL.n652 VSUBS 0.012288f
C1448 VTAIL.n653 VSUBS 0.050983f
C1449 VTAIL.n654 VSUBS 0.03693f
C1450 VTAIL.n655 VSUBS 1.54442f
C1451 VDD2.t3 VSUBS 0.315467f
C1452 VDD2.t2 VSUBS 0.315467f
C1453 VDD2.n0 VSUBS 3.37755f
C1454 VDD2.t0 VSUBS 0.315467f
C1455 VDD2.t1 VSUBS 0.315467f
C1456 VDD2.n1 VSUBS 2.5418f
C1457 VDD2.n2 VSUBS 4.602241f
C1458 VN.t3 VSUBS 3.54075f
C1459 VN.t2 VSUBS 3.53513f
C1460 VN.n0 VSUBS 2.28415f
C1461 VN.t1 VSUBS 3.54075f
C1462 VN.t0 VSUBS 3.53513f
C1463 VN.n1 VSUBS 4.09449f
.ends

