* NGSPICE file created from diff_pair_sample_0974.ext - technology: sky130A

.subckt diff_pair_sample_0974 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t6 VP.t0 VDD1.t3 w_n2740_n3454# sky130_fd_pr__pfet_01v8 ad=4.8477 pd=25.64 as=2.05095 ps=12.76 w=12.43 l=2.62
X1 VTAIL.t5 VP.t1 VDD1.t0 w_n2740_n3454# sky130_fd_pr__pfet_01v8 ad=4.8477 pd=25.64 as=2.05095 ps=12.76 w=12.43 l=2.62
X2 VDD2.t3 VN.t0 VTAIL.t2 w_n2740_n3454# sky130_fd_pr__pfet_01v8 ad=2.05095 pd=12.76 as=4.8477 ps=25.64 w=12.43 l=2.62
X3 B.t11 B.t9 B.t10 w_n2740_n3454# sky130_fd_pr__pfet_01v8 ad=4.8477 pd=25.64 as=0 ps=0 w=12.43 l=2.62
X4 VDD1.t2 VP.t2 VTAIL.t4 w_n2740_n3454# sky130_fd_pr__pfet_01v8 ad=2.05095 pd=12.76 as=4.8477 ps=25.64 w=12.43 l=2.62
X5 VDD1.t1 VP.t3 VTAIL.t3 w_n2740_n3454# sky130_fd_pr__pfet_01v8 ad=2.05095 pd=12.76 as=4.8477 ps=25.64 w=12.43 l=2.62
X6 VDD2.t2 VN.t1 VTAIL.t0 w_n2740_n3454# sky130_fd_pr__pfet_01v8 ad=2.05095 pd=12.76 as=4.8477 ps=25.64 w=12.43 l=2.62
X7 VTAIL.t1 VN.t2 VDD2.t1 w_n2740_n3454# sky130_fd_pr__pfet_01v8 ad=4.8477 pd=25.64 as=2.05095 ps=12.76 w=12.43 l=2.62
X8 B.t8 B.t6 B.t7 w_n2740_n3454# sky130_fd_pr__pfet_01v8 ad=4.8477 pd=25.64 as=0 ps=0 w=12.43 l=2.62
X9 B.t5 B.t3 B.t4 w_n2740_n3454# sky130_fd_pr__pfet_01v8 ad=4.8477 pd=25.64 as=0 ps=0 w=12.43 l=2.62
X10 VTAIL.t7 VN.t3 VDD2.t0 w_n2740_n3454# sky130_fd_pr__pfet_01v8 ad=4.8477 pd=25.64 as=2.05095 ps=12.76 w=12.43 l=2.62
X11 B.t2 B.t0 B.t1 w_n2740_n3454# sky130_fd_pr__pfet_01v8 ad=4.8477 pd=25.64 as=0 ps=0 w=12.43 l=2.62
R0 VP.n14 VP.n0 161.3
R1 VP.n13 VP.n12 161.3
R2 VP.n11 VP.n1 161.3
R3 VP.n10 VP.n9 161.3
R4 VP.n8 VP.n2 161.3
R5 VP.n7 VP.n6 161.3
R6 VP.n4 VP.t0 150.673
R7 VP.n4 VP.t3 149.894
R8 VP.n3 VP.t1 114.338
R9 VP.n15 VP.t2 114.338
R10 VP.n5 VP.n3 99.7463
R11 VP.n16 VP.n15 99.7463
R12 VP.n9 VP.n1 56.5193
R13 VP.n5 VP.n4 51.0251
R14 VP.n8 VP.n7 24.4675
R15 VP.n9 VP.n8 24.4675
R16 VP.n13 VP.n1 24.4675
R17 VP.n14 VP.n13 24.4675
R18 VP.n7 VP.n3 11.0107
R19 VP.n15 VP.n14 11.0107
R20 VP.n6 VP.n5 0.278367
R21 VP.n16 VP.n0 0.278367
R22 VP.n6 VP.n2 0.189894
R23 VP.n10 VP.n2 0.189894
R24 VP.n11 VP.n10 0.189894
R25 VP.n12 VP.n11 0.189894
R26 VP.n12 VP.n0 0.189894
R27 VP VP.n16 0.153454
R28 VDD1 VDD1.n1 115.026
R29 VDD1 VDD1.n0 72.5
R30 VDD1.n0 VDD1.t3 2.61554
R31 VDD1.n0 VDD1.t1 2.61554
R32 VDD1.n1 VDD1.t0 2.61554
R33 VDD1.n1 VDD1.t2 2.61554
R34 VTAIL.n5 VTAIL.t6 58.3783
R35 VTAIL.n4 VTAIL.t0 58.3783
R36 VTAIL.n3 VTAIL.t7 58.3783
R37 VTAIL.n7 VTAIL.t2 58.3781
R38 VTAIL.n0 VTAIL.t1 58.3781
R39 VTAIL.n1 VTAIL.t4 58.3781
R40 VTAIL.n2 VTAIL.t5 58.3781
R41 VTAIL.n6 VTAIL.t3 58.3781
R42 VTAIL.n7 VTAIL.n6 25.6255
R43 VTAIL.n3 VTAIL.n2 25.6255
R44 VTAIL.n4 VTAIL.n3 2.5436
R45 VTAIL.n6 VTAIL.n5 2.5436
R46 VTAIL.n2 VTAIL.n1 2.5436
R47 VTAIL VTAIL.n0 1.33024
R48 VTAIL VTAIL.n7 1.21386
R49 VTAIL.n5 VTAIL.n4 0.470328
R50 VTAIL.n1 VTAIL.n0 0.470328
R51 VN.n0 VN.t2 150.673
R52 VN.n1 VN.t1 150.673
R53 VN.n0 VN.t0 149.894
R54 VN.n1 VN.t3 149.894
R55 VN VN.n1 51.304
R56 VN VN.n0 4.29263
R57 VDD2.n2 VDD2.n0 114.501
R58 VDD2.n2 VDD2.n1 72.4419
R59 VDD2.n1 VDD2.t0 2.61554
R60 VDD2.n1 VDD2.t2 2.61554
R61 VDD2.n0 VDD2.t1 2.61554
R62 VDD2.n0 VDD2.t3 2.61554
R63 VDD2 VDD2.n2 0.0586897
R64 B.n472 B.n71 585
R65 B.n474 B.n473 585
R66 B.n475 B.n70 585
R67 B.n477 B.n476 585
R68 B.n478 B.n69 585
R69 B.n480 B.n479 585
R70 B.n481 B.n68 585
R71 B.n483 B.n482 585
R72 B.n484 B.n67 585
R73 B.n486 B.n485 585
R74 B.n487 B.n66 585
R75 B.n489 B.n488 585
R76 B.n490 B.n65 585
R77 B.n492 B.n491 585
R78 B.n493 B.n64 585
R79 B.n495 B.n494 585
R80 B.n496 B.n63 585
R81 B.n498 B.n497 585
R82 B.n499 B.n62 585
R83 B.n501 B.n500 585
R84 B.n502 B.n61 585
R85 B.n504 B.n503 585
R86 B.n505 B.n60 585
R87 B.n507 B.n506 585
R88 B.n508 B.n59 585
R89 B.n510 B.n509 585
R90 B.n511 B.n58 585
R91 B.n513 B.n512 585
R92 B.n514 B.n57 585
R93 B.n516 B.n515 585
R94 B.n517 B.n56 585
R95 B.n519 B.n518 585
R96 B.n520 B.n55 585
R97 B.n522 B.n521 585
R98 B.n523 B.n54 585
R99 B.n525 B.n524 585
R100 B.n526 B.n53 585
R101 B.n528 B.n527 585
R102 B.n529 B.n52 585
R103 B.n531 B.n530 585
R104 B.n532 B.n51 585
R105 B.n534 B.n533 585
R106 B.n535 B.n48 585
R107 B.n538 B.n537 585
R108 B.n539 B.n47 585
R109 B.n541 B.n540 585
R110 B.n542 B.n46 585
R111 B.n544 B.n543 585
R112 B.n545 B.n45 585
R113 B.n547 B.n546 585
R114 B.n548 B.n41 585
R115 B.n550 B.n549 585
R116 B.n551 B.n40 585
R117 B.n553 B.n552 585
R118 B.n554 B.n39 585
R119 B.n556 B.n555 585
R120 B.n557 B.n38 585
R121 B.n559 B.n558 585
R122 B.n560 B.n37 585
R123 B.n562 B.n561 585
R124 B.n563 B.n36 585
R125 B.n565 B.n564 585
R126 B.n566 B.n35 585
R127 B.n568 B.n567 585
R128 B.n569 B.n34 585
R129 B.n571 B.n570 585
R130 B.n572 B.n33 585
R131 B.n574 B.n573 585
R132 B.n575 B.n32 585
R133 B.n577 B.n576 585
R134 B.n578 B.n31 585
R135 B.n580 B.n579 585
R136 B.n581 B.n30 585
R137 B.n583 B.n582 585
R138 B.n584 B.n29 585
R139 B.n586 B.n585 585
R140 B.n587 B.n28 585
R141 B.n589 B.n588 585
R142 B.n590 B.n27 585
R143 B.n592 B.n591 585
R144 B.n593 B.n26 585
R145 B.n595 B.n594 585
R146 B.n596 B.n25 585
R147 B.n598 B.n597 585
R148 B.n599 B.n24 585
R149 B.n601 B.n600 585
R150 B.n602 B.n23 585
R151 B.n604 B.n603 585
R152 B.n605 B.n22 585
R153 B.n607 B.n606 585
R154 B.n608 B.n21 585
R155 B.n610 B.n609 585
R156 B.n611 B.n20 585
R157 B.n613 B.n612 585
R158 B.n614 B.n19 585
R159 B.n471 B.n470 585
R160 B.n469 B.n72 585
R161 B.n468 B.n467 585
R162 B.n466 B.n73 585
R163 B.n465 B.n464 585
R164 B.n463 B.n74 585
R165 B.n462 B.n461 585
R166 B.n460 B.n75 585
R167 B.n459 B.n458 585
R168 B.n457 B.n76 585
R169 B.n456 B.n455 585
R170 B.n454 B.n77 585
R171 B.n453 B.n452 585
R172 B.n451 B.n78 585
R173 B.n450 B.n449 585
R174 B.n448 B.n79 585
R175 B.n447 B.n446 585
R176 B.n445 B.n80 585
R177 B.n444 B.n443 585
R178 B.n442 B.n81 585
R179 B.n441 B.n440 585
R180 B.n439 B.n82 585
R181 B.n438 B.n437 585
R182 B.n436 B.n83 585
R183 B.n435 B.n434 585
R184 B.n433 B.n84 585
R185 B.n432 B.n431 585
R186 B.n430 B.n85 585
R187 B.n429 B.n428 585
R188 B.n427 B.n86 585
R189 B.n426 B.n425 585
R190 B.n424 B.n87 585
R191 B.n423 B.n422 585
R192 B.n421 B.n88 585
R193 B.n420 B.n419 585
R194 B.n418 B.n89 585
R195 B.n417 B.n416 585
R196 B.n415 B.n90 585
R197 B.n414 B.n413 585
R198 B.n412 B.n91 585
R199 B.n411 B.n410 585
R200 B.n409 B.n92 585
R201 B.n408 B.n407 585
R202 B.n406 B.n93 585
R203 B.n405 B.n404 585
R204 B.n403 B.n94 585
R205 B.n402 B.n401 585
R206 B.n400 B.n95 585
R207 B.n399 B.n398 585
R208 B.n397 B.n96 585
R209 B.n396 B.n395 585
R210 B.n394 B.n97 585
R211 B.n393 B.n392 585
R212 B.n391 B.n98 585
R213 B.n390 B.n389 585
R214 B.n388 B.n99 585
R215 B.n387 B.n386 585
R216 B.n385 B.n100 585
R217 B.n384 B.n383 585
R218 B.n382 B.n101 585
R219 B.n381 B.n380 585
R220 B.n379 B.n102 585
R221 B.n378 B.n377 585
R222 B.n376 B.n103 585
R223 B.n375 B.n374 585
R224 B.n373 B.n104 585
R225 B.n372 B.n371 585
R226 B.n370 B.n105 585
R227 B.n369 B.n368 585
R228 B.n222 B.n155 585
R229 B.n224 B.n223 585
R230 B.n225 B.n154 585
R231 B.n227 B.n226 585
R232 B.n228 B.n153 585
R233 B.n230 B.n229 585
R234 B.n231 B.n152 585
R235 B.n233 B.n232 585
R236 B.n234 B.n151 585
R237 B.n236 B.n235 585
R238 B.n237 B.n150 585
R239 B.n239 B.n238 585
R240 B.n240 B.n149 585
R241 B.n242 B.n241 585
R242 B.n243 B.n148 585
R243 B.n245 B.n244 585
R244 B.n246 B.n147 585
R245 B.n248 B.n247 585
R246 B.n249 B.n146 585
R247 B.n251 B.n250 585
R248 B.n252 B.n145 585
R249 B.n254 B.n253 585
R250 B.n255 B.n144 585
R251 B.n257 B.n256 585
R252 B.n258 B.n143 585
R253 B.n260 B.n259 585
R254 B.n261 B.n142 585
R255 B.n263 B.n262 585
R256 B.n264 B.n141 585
R257 B.n266 B.n265 585
R258 B.n267 B.n140 585
R259 B.n269 B.n268 585
R260 B.n270 B.n139 585
R261 B.n272 B.n271 585
R262 B.n273 B.n138 585
R263 B.n275 B.n274 585
R264 B.n276 B.n137 585
R265 B.n278 B.n277 585
R266 B.n279 B.n136 585
R267 B.n281 B.n280 585
R268 B.n282 B.n135 585
R269 B.n284 B.n283 585
R270 B.n285 B.n132 585
R271 B.n288 B.n287 585
R272 B.n289 B.n131 585
R273 B.n291 B.n290 585
R274 B.n292 B.n130 585
R275 B.n294 B.n293 585
R276 B.n295 B.n129 585
R277 B.n297 B.n296 585
R278 B.n298 B.n128 585
R279 B.n303 B.n302 585
R280 B.n304 B.n127 585
R281 B.n306 B.n305 585
R282 B.n307 B.n126 585
R283 B.n309 B.n308 585
R284 B.n310 B.n125 585
R285 B.n312 B.n311 585
R286 B.n313 B.n124 585
R287 B.n315 B.n314 585
R288 B.n316 B.n123 585
R289 B.n318 B.n317 585
R290 B.n319 B.n122 585
R291 B.n321 B.n320 585
R292 B.n322 B.n121 585
R293 B.n324 B.n323 585
R294 B.n325 B.n120 585
R295 B.n327 B.n326 585
R296 B.n328 B.n119 585
R297 B.n330 B.n329 585
R298 B.n331 B.n118 585
R299 B.n333 B.n332 585
R300 B.n334 B.n117 585
R301 B.n336 B.n335 585
R302 B.n337 B.n116 585
R303 B.n339 B.n338 585
R304 B.n340 B.n115 585
R305 B.n342 B.n341 585
R306 B.n343 B.n114 585
R307 B.n345 B.n344 585
R308 B.n346 B.n113 585
R309 B.n348 B.n347 585
R310 B.n349 B.n112 585
R311 B.n351 B.n350 585
R312 B.n352 B.n111 585
R313 B.n354 B.n353 585
R314 B.n355 B.n110 585
R315 B.n357 B.n356 585
R316 B.n358 B.n109 585
R317 B.n360 B.n359 585
R318 B.n361 B.n108 585
R319 B.n363 B.n362 585
R320 B.n364 B.n107 585
R321 B.n366 B.n365 585
R322 B.n367 B.n106 585
R323 B.n221 B.n220 585
R324 B.n219 B.n156 585
R325 B.n218 B.n217 585
R326 B.n216 B.n157 585
R327 B.n215 B.n214 585
R328 B.n213 B.n158 585
R329 B.n212 B.n211 585
R330 B.n210 B.n159 585
R331 B.n209 B.n208 585
R332 B.n207 B.n160 585
R333 B.n206 B.n205 585
R334 B.n204 B.n161 585
R335 B.n203 B.n202 585
R336 B.n201 B.n162 585
R337 B.n200 B.n199 585
R338 B.n198 B.n163 585
R339 B.n197 B.n196 585
R340 B.n195 B.n164 585
R341 B.n194 B.n193 585
R342 B.n192 B.n165 585
R343 B.n191 B.n190 585
R344 B.n189 B.n166 585
R345 B.n188 B.n187 585
R346 B.n186 B.n167 585
R347 B.n185 B.n184 585
R348 B.n183 B.n168 585
R349 B.n182 B.n181 585
R350 B.n180 B.n169 585
R351 B.n179 B.n178 585
R352 B.n177 B.n170 585
R353 B.n176 B.n175 585
R354 B.n174 B.n171 585
R355 B.n173 B.n172 585
R356 B.n2 B.n0 585
R357 B.n665 B.n1 585
R358 B.n664 B.n663 585
R359 B.n662 B.n3 585
R360 B.n661 B.n660 585
R361 B.n659 B.n4 585
R362 B.n658 B.n657 585
R363 B.n656 B.n5 585
R364 B.n655 B.n654 585
R365 B.n653 B.n6 585
R366 B.n652 B.n651 585
R367 B.n650 B.n7 585
R368 B.n649 B.n648 585
R369 B.n647 B.n8 585
R370 B.n646 B.n645 585
R371 B.n644 B.n9 585
R372 B.n643 B.n642 585
R373 B.n641 B.n10 585
R374 B.n640 B.n639 585
R375 B.n638 B.n11 585
R376 B.n637 B.n636 585
R377 B.n635 B.n12 585
R378 B.n634 B.n633 585
R379 B.n632 B.n13 585
R380 B.n631 B.n630 585
R381 B.n629 B.n14 585
R382 B.n628 B.n627 585
R383 B.n626 B.n15 585
R384 B.n625 B.n624 585
R385 B.n623 B.n16 585
R386 B.n622 B.n621 585
R387 B.n620 B.n17 585
R388 B.n619 B.n618 585
R389 B.n617 B.n18 585
R390 B.n616 B.n615 585
R391 B.n667 B.n666 585
R392 B.n222 B.n221 550.159
R393 B.n616 B.n19 550.159
R394 B.n369 B.n106 550.159
R395 B.n472 B.n471 550.159
R396 B.n299 B.t6 322.414
R397 B.n133 B.t0 322.414
R398 B.n42 B.t9 322.414
R399 B.n49 B.t3 322.414
R400 B.n299 B.t8 167.906
R401 B.n49 B.t4 167.906
R402 B.n133 B.t2 167.892
R403 B.n42 B.t10 167.892
R404 B.n221 B.n156 163.367
R405 B.n217 B.n156 163.367
R406 B.n217 B.n216 163.367
R407 B.n216 B.n215 163.367
R408 B.n215 B.n158 163.367
R409 B.n211 B.n158 163.367
R410 B.n211 B.n210 163.367
R411 B.n210 B.n209 163.367
R412 B.n209 B.n160 163.367
R413 B.n205 B.n160 163.367
R414 B.n205 B.n204 163.367
R415 B.n204 B.n203 163.367
R416 B.n203 B.n162 163.367
R417 B.n199 B.n162 163.367
R418 B.n199 B.n198 163.367
R419 B.n198 B.n197 163.367
R420 B.n197 B.n164 163.367
R421 B.n193 B.n164 163.367
R422 B.n193 B.n192 163.367
R423 B.n192 B.n191 163.367
R424 B.n191 B.n166 163.367
R425 B.n187 B.n166 163.367
R426 B.n187 B.n186 163.367
R427 B.n186 B.n185 163.367
R428 B.n185 B.n168 163.367
R429 B.n181 B.n168 163.367
R430 B.n181 B.n180 163.367
R431 B.n180 B.n179 163.367
R432 B.n179 B.n170 163.367
R433 B.n175 B.n170 163.367
R434 B.n175 B.n174 163.367
R435 B.n174 B.n173 163.367
R436 B.n173 B.n2 163.367
R437 B.n666 B.n2 163.367
R438 B.n666 B.n665 163.367
R439 B.n665 B.n664 163.367
R440 B.n664 B.n3 163.367
R441 B.n660 B.n3 163.367
R442 B.n660 B.n659 163.367
R443 B.n659 B.n658 163.367
R444 B.n658 B.n5 163.367
R445 B.n654 B.n5 163.367
R446 B.n654 B.n653 163.367
R447 B.n653 B.n652 163.367
R448 B.n652 B.n7 163.367
R449 B.n648 B.n7 163.367
R450 B.n648 B.n647 163.367
R451 B.n647 B.n646 163.367
R452 B.n646 B.n9 163.367
R453 B.n642 B.n9 163.367
R454 B.n642 B.n641 163.367
R455 B.n641 B.n640 163.367
R456 B.n640 B.n11 163.367
R457 B.n636 B.n11 163.367
R458 B.n636 B.n635 163.367
R459 B.n635 B.n634 163.367
R460 B.n634 B.n13 163.367
R461 B.n630 B.n13 163.367
R462 B.n630 B.n629 163.367
R463 B.n629 B.n628 163.367
R464 B.n628 B.n15 163.367
R465 B.n624 B.n15 163.367
R466 B.n624 B.n623 163.367
R467 B.n623 B.n622 163.367
R468 B.n622 B.n17 163.367
R469 B.n618 B.n17 163.367
R470 B.n618 B.n617 163.367
R471 B.n617 B.n616 163.367
R472 B.n223 B.n222 163.367
R473 B.n223 B.n154 163.367
R474 B.n227 B.n154 163.367
R475 B.n228 B.n227 163.367
R476 B.n229 B.n228 163.367
R477 B.n229 B.n152 163.367
R478 B.n233 B.n152 163.367
R479 B.n234 B.n233 163.367
R480 B.n235 B.n234 163.367
R481 B.n235 B.n150 163.367
R482 B.n239 B.n150 163.367
R483 B.n240 B.n239 163.367
R484 B.n241 B.n240 163.367
R485 B.n241 B.n148 163.367
R486 B.n245 B.n148 163.367
R487 B.n246 B.n245 163.367
R488 B.n247 B.n246 163.367
R489 B.n247 B.n146 163.367
R490 B.n251 B.n146 163.367
R491 B.n252 B.n251 163.367
R492 B.n253 B.n252 163.367
R493 B.n253 B.n144 163.367
R494 B.n257 B.n144 163.367
R495 B.n258 B.n257 163.367
R496 B.n259 B.n258 163.367
R497 B.n259 B.n142 163.367
R498 B.n263 B.n142 163.367
R499 B.n264 B.n263 163.367
R500 B.n265 B.n264 163.367
R501 B.n265 B.n140 163.367
R502 B.n269 B.n140 163.367
R503 B.n270 B.n269 163.367
R504 B.n271 B.n270 163.367
R505 B.n271 B.n138 163.367
R506 B.n275 B.n138 163.367
R507 B.n276 B.n275 163.367
R508 B.n277 B.n276 163.367
R509 B.n277 B.n136 163.367
R510 B.n281 B.n136 163.367
R511 B.n282 B.n281 163.367
R512 B.n283 B.n282 163.367
R513 B.n283 B.n132 163.367
R514 B.n288 B.n132 163.367
R515 B.n289 B.n288 163.367
R516 B.n290 B.n289 163.367
R517 B.n290 B.n130 163.367
R518 B.n294 B.n130 163.367
R519 B.n295 B.n294 163.367
R520 B.n296 B.n295 163.367
R521 B.n296 B.n128 163.367
R522 B.n303 B.n128 163.367
R523 B.n304 B.n303 163.367
R524 B.n305 B.n304 163.367
R525 B.n305 B.n126 163.367
R526 B.n309 B.n126 163.367
R527 B.n310 B.n309 163.367
R528 B.n311 B.n310 163.367
R529 B.n311 B.n124 163.367
R530 B.n315 B.n124 163.367
R531 B.n316 B.n315 163.367
R532 B.n317 B.n316 163.367
R533 B.n317 B.n122 163.367
R534 B.n321 B.n122 163.367
R535 B.n322 B.n321 163.367
R536 B.n323 B.n322 163.367
R537 B.n323 B.n120 163.367
R538 B.n327 B.n120 163.367
R539 B.n328 B.n327 163.367
R540 B.n329 B.n328 163.367
R541 B.n329 B.n118 163.367
R542 B.n333 B.n118 163.367
R543 B.n334 B.n333 163.367
R544 B.n335 B.n334 163.367
R545 B.n335 B.n116 163.367
R546 B.n339 B.n116 163.367
R547 B.n340 B.n339 163.367
R548 B.n341 B.n340 163.367
R549 B.n341 B.n114 163.367
R550 B.n345 B.n114 163.367
R551 B.n346 B.n345 163.367
R552 B.n347 B.n346 163.367
R553 B.n347 B.n112 163.367
R554 B.n351 B.n112 163.367
R555 B.n352 B.n351 163.367
R556 B.n353 B.n352 163.367
R557 B.n353 B.n110 163.367
R558 B.n357 B.n110 163.367
R559 B.n358 B.n357 163.367
R560 B.n359 B.n358 163.367
R561 B.n359 B.n108 163.367
R562 B.n363 B.n108 163.367
R563 B.n364 B.n363 163.367
R564 B.n365 B.n364 163.367
R565 B.n365 B.n106 163.367
R566 B.n370 B.n369 163.367
R567 B.n371 B.n370 163.367
R568 B.n371 B.n104 163.367
R569 B.n375 B.n104 163.367
R570 B.n376 B.n375 163.367
R571 B.n377 B.n376 163.367
R572 B.n377 B.n102 163.367
R573 B.n381 B.n102 163.367
R574 B.n382 B.n381 163.367
R575 B.n383 B.n382 163.367
R576 B.n383 B.n100 163.367
R577 B.n387 B.n100 163.367
R578 B.n388 B.n387 163.367
R579 B.n389 B.n388 163.367
R580 B.n389 B.n98 163.367
R581 B.n393 B.n98 163.367
R582 B.n394 B.n393 163.367
R583 B.n395 B.n394 163.367
R584 B.n395 B.n96 163.367
R585 B.n399 B.n96 163.367
R586 B.n400 B.n399 163.367
R587 B.n401 B.n400 163.367
R588 B.n401 B.n94 163.367
R589 B.n405 B.n94 163.367
R590 B.n406 B.n405 163.367
R591 B.n407 B.n406 163.367
R592 B.n407 B.n92 163.367
R593 B.n411 B.n92 163.367
R594 B.n412 B.n411 163.367
R595 B.n413 B.n412 163.367
R596 B.n413 B.n90 163.367
R597 B.n417 B.n90 163.367
R598 B.n418 B.n417 163.367
R599 B.n419 B.n418 163.367
R600 B.n419 B.n88 163.367
R601 B.n423 B.n88 163.367
R602 B.n424 B.n423 163.367
R603 B.n425 B.n424 163.367
R604 B.n425 B.n86 163.367
R605 B.n429 B.n86 163.367
R606 B.n430 B.n429 163.367
R607 B.n431 B.n430 163.367
R608 B.n431 B.n84 163.367
R609 B.n435 B.n84 163.367
R610 B.n436 B.n435 163.367
R611 B.n437 B.n436 163.367
R612 B.n437 B.n82 163.367
R613 B.n441 B.n82 163.367
R614 B.n442 B.n441 163.367
R615 B.n443 B.n442 163.367
R616 B.n443 B.n80 163.367
R617 B.n447 B.n80 163.367
R618 B.n448 B.n447 163.367
R619 B.n449 B.n448 163.367
R620 B.n449 B.n78 163.367
R621 B.n453 B.n78 163.367
R622 B.n454 B.n453 163.367
R623 B.n455 B.n454 163.367
R624 B.n455 B.n76 163.367
R625 B.n459 B.n76 163.367
R626 B.n460 B.n459 163.367
R627 B.n461 B.n460 163.367
R628 B.n461 B.n74 163.367
R629 B.n465 B.n74 163.367
R630 B.n466 B.n465 163.367
R631 B.n467 B.n466 163.367
R632 B.n467 B.n72 163.367
R633 B.n471 B.n72 163.367
R634 B.n612 B.n19 163.367
R635 B.n612 B.n611 163.367
R636 B.n611 B.n610 163.367
R637 B.n610 B.n21 163.367
R638 B.n606 B.n21 163.367
R639 B.n606 B.n605 163.367
R640 B.n605 B.n604 163.367
R641 B.n604 B.n23 163.367
R642 B.n600 B.n23 163.367
R643 B.n600 B.n599 163.367
R644 B.n599 B.n598 163.367
R645 B.n598 B.n25 163.367
R646 B.n594 B.n25 163.367
R647 B.n594 B.n593 163.367
R648 B.n593 B.n592 163.367
R649 B.n592 B.n27 163.367
R650 B.n588 B.n27 163.367
R651 B.n588 B.n587 163.367
R652 B.n587 B.n586 163.367
R653 B.n586 B.n29 163.367
R654 B.n582 B.n29 163.367
R655 B.n582 B.n581 163.367
R656 B.n581 B.n580 163.367
R657 B.n580 B.n31 163.367
R658 B.n576 B.n31 163.367
R659 B.n576 B.n575 163.367
R660 B.n575 B.n574 163.367
R661 B.n574 B.n33 163.367
R662 B.n570 B.n33 163.367
R663 B.n570 B.n569 163.367
R664 B.n569 B.n568 163.367
R665 B.n568 B.n35 163.367
R666 B.n564 B.n35 163.367
R667 B.n564 B.n563 163.367
R668 B.n563 B.n562 163.367
R669 B.n562 B.n37 163.367
R670 B.n558 B.n37 163.367
R671 B.n558 B.n557 163.367
R672 B.n557 B.n556 163.367
R673 B.n556 B.n39 163.367
R674 B.n552 B.n39 163.367
R675 B.n552 B.n551 163.367
R676 B.n551 B.n550 163.367
R677 B.n550 B.n41 163.367
R678 B.n546 B.n41 163.367
R679 B.n546 B.n545 163.367
R680 B.n545 B.n544 163.367
R681 B.n544 B.n46 163.367
R682 B.n540 B.n46 163.367
R683 B.n540 B.n539 163.367
R684 B.n539 B.n538 163.367
R685 B.n538 B.n48 163.367
R686 B.n533 B.n48 163.367
R687 B.n533 B.n532 163.367
R688 B.n532 B.n531 163.367
R689 B.n531 B.n52 163.367
R690 B.n527 B.n52 163.367
R691 B.n527 B.n526 163.367
R692 B.n526 B.n525 163.367
R693 B.n525 B.n54 163.367
R694 B.n521 B.n54 163.367
R695 B.n521 B.n520 163.367
R696 B.n520 B.n519 163.367
R697 B.n519 B.n56 163.367
R698 B.n515 B.n56 163.367
R699 B.n515 B.n514 163.367
R700 B.n514 B.n513 163.367
R701 B.n513 B.n58 163.367
R702 B.n509 B.n58 163.367
R703 B.n509 B.n508 163.367
R704 B.n508 B.n507 163.367
R705 B.n507 B.n60 163.367
R706 B.n503 B.n60 163.367
R707 B.n503 B.n502 163.367
R708 B.n502 B.n501 163.367
R709 B.n501 B.n62 163.367
R710 B.n497 B.n62 163.367
R711 B.n497 B.n496 163.367
R712 B.n496 B.n495 163.367
R713 B.n495 B.n64 163.367
R714 B.n491 B.n64 163.367
R715 B.n491 B.n490 163.367
R716 B.n490 B.n489 163.367
R717 B.n489 B.n66 163.367
R718 B.n485 B.n66 163.367
R719 B.n485 B.n484 163.367
R720 B.n484 B.n483 163.367
R721 B.n483 B.n68 163.367
R722 B.n479 B.n68 163.367
R723 B.n479 B.n478 163.367
R724 B.n478 B.n477 163.367
R725 B.n477 B.n70 163.367
R726 B.n473 B.n70 163.367
R727 B.n473 B.n472 163.367
R728 B.n300 B.t7 110.695
R729 B.n50 B.t5 110.695
R730 B.n134 B.t1 110.68
R731 B.n43 B.t11 110.68
R732 B.n301 B.n300 59.5399
R733 B.n286 B.n134 59.5399
R734 B.n44 B.n43 59.5399
R735 B.n536 B.n50 59.5399
R736 B.n300 B.n299 57.2126
R737 B.n134 B.n133 57.2126
R738 B.n43 B.n42 57.2126
R739 B.n50 B.n49 57.2126
R740 B.n615 B.n614 35.7468
R741 B.n368 B.n367 35.7468
R742 B.n220 B.n155 35.7468
R743 B.n470 B.n71 35.7468
R744 B B.n667 18.0485
R745 B.n614 B.n613 10.6151
R746 B.n613 B.n20 10.6151
R747 B.n609 B.n20 10.6151
R748 B.n609 B.n608 10.6151
R749 B.n608 B.n607 10.6151
R750 B.n607 B.n22 10.6151
R751 B.n603 B.n22 10.6151
R752 B.n603 B.n602 10.6151
R753 B.n602 B.n601 10.6151
R754 B.n601 B.n24 10.6151
R755 B.n597 B.n24 10.6151
R756 B.n597 B.n596 10.6151
R757 B.n596 B.n595 10.6151
R758 B.n595 B.n26 10.6151
R759 B.n591 B.n26 10.6151
R760 B.n591 B.n590 10.6151
R761 B.n590 B.n589 10.6151
R762 B.n589 B.n28 10.6151
R763 B.n585 B.n28 10.6151
R764 B.n585 B.n584 10.6151
R765 B.n584 B.n583 10.6151
R766 B.n583 B.n30 10.6151
R767 B.n579 B.n30 10.6151
R768 B.n579 B.n578 10.6151
R769 B.n578 B.n577 10.6151
R770 B.n577 B.n32 10.6151
R771 B.n573 B.n32 10.6151
R772 B.n573 B.n572 10.6151
R773 B.n572 B.n571 10.6151
R774 B.n571 B.n34 10.6151
R775 B.n567 B.n34 10.6151
R776 B.n567 B.n566 10.6151
R777 B.n566 B.n565 10.6151
R778 B.n565 B.n36 10.6151
R779 B.n561 B.n36 10.6151
R780 B.n561 B.n560 10.6151
R781 B.n560 B.n559 10.6151
R782 B.n559 B.n38 10.6151
R783 B.n555 B.n38 10.6151
R784 B.n555 B.n554 10.6151
R785 B.n554 B.n553 10.6151
R786 B.n553 B.n40 10.6151
R787 B.n549 B.n548 10.6151
R788 B.n548 B.n547 10.6151
R789 B.n547 B.n45 10.6151
R790 B.n543 B.n45 10.6151
R791 B.n543 B.n542 10.6151
R792 B.n542 B.n541 10.6151
R793 B.n541 B.n47 10.6151
R794 B.n537 B.n47 10.6151
R795 B.n535 B.n534 10.6151
R796 B.n534 B.n51 10.6151
R797 B.n530 B.n51 10.6151
R798 B.n530 B.n529 10.6151
R799 B.n529 B.n528 10.6151
R800 B.n528 B.n53 10.6151
R801 B.n524 B.n53 10.6151
R802 B.n524 B.n523 10.6151
R803 B.n523 B.n522 10.6151
R804 B.n522 B.n55 10.6151
R805 B.n518 B.n55 10.6151
R806 B.n518 B.n517 10.6151
R807 B.n517 B.n516 10.6151
R808 B.n516 B.n57 10.6151
R809 B.n512 B.n57 10.6151
R810 B.n512 B.n511 10.6151
R811 B.n511 B.n510 10.6151
R812 B.n510 B.n59 10.6151
R813 B.n506 B.n59 10.6151
R814 B.n506 B.n505 10.6151
R815 B.n505 B.n504 10.6151
R816 B.n504 B.n61 10.6151
R817 B.n500 B.n61 10.6151
R818 B.n500 B.n499 10.6151
R819 B.n499 B.n498 10.6151
R820 B.n498 B.n63 10.6151
R821 B.n494 B.n63 10.6151
R822 B.n494 B.n493 10.6151
R823 B.n493 B.n492 10.6151
R824 B.n492 B.n65 10.6151
R825 B.n488 B.n65 10.6151
R826 B.n488 B.n487 10.6151
R827 B.n487 B.n486 10.6151
R828 B.n486 B.n67 10.6151
R829 B.n482 B.n67 10.6151
R830 B.n482 B.n481 10.6151
R831 B.n481 B.n480 10.6151
R832 B.n480 B.n69 10.6151
R833 B.n476 B.n69 10.6151
R834 B.n476 B.n475 10.6151
R835 B.n475 B.n474 10.6151
R836 B.n474 B.n71 10.6151
R837 B.n368 B.n105 10.6151
R838 B.n372 B.n105 10.6151
R839 B.n373 B.n372 10.6151
R840 B.n374 B.n373 10.6151
R841 B.n374 B.n103 10.6151
R842 B.n378 B.n103 10.6151
R843 B.n379 B.n378 10.6151
R844 B.n380 B.n379 10.6151
R845 B.n380 B.n101 10.6151
R846 B.n384 B.n101 10.6151
R847 B.n385 B.n384 10.6151
R848 B.n386 B.n385 10.6151
R849 B.n386 B.n99 10.6151
R850 B.n390 B.n99 10.6151
R851 B.n391 B.n390 10.6151
R852 B.n392 B.n391 10.6151
R853 B.n392 B.n97 10.6151
R854 B.n396 B.n97 10.6151
R855 B.n397 B.n396 10.6151
R856 B.n398 B.n397 10.6151
R857 B.n398 B.n95 10.6151
R858 B.n402 B.n95 10.6151
R859 B.n403 B.n402 10.6151
R860 B.n404 B.n403 10.6151
R861 B.n404 B.n93 10.6151
R862 B.n408 B.n93 10.6151
R863 B.n409 B.n408 10.6151
R864 B.n410 B.n409 10.6151
R865 B.n410 B.n91 10.6151
R866 B.n414 B.n91 10.6151
R867 B.n415 B.n414 10.6151
R868 B.n416 B.n415 10.6151
R869 B.n416 B.n89 10.6151
R870 B.n420 B.n89 10.6151
R871 B.n421 B.n420 10.6151
R872 B.n422 B.n421 10.6151
R873 B.n422 B.n87 10.6151
R874 B.n426 B.n87 10.6151
R875 B.n427 B.n426 10.6151
R876 B.n428 B.n427 10.6151
R877 B.n428 B.n85 10.6151
R878 B.n432 B.n85 10.6151
R879 B.n433 B.n432 10.6151
R880 B.n434 B.n433 10.6151
R881 B.n434 B.n83 10.6151
R882 B.n438 B.n83 10.6151
R883 B.n439 B.n438 10.6151
R884 B.n440 B.n439 10.6151
R885 B.n440 B.n81 10.6151
R886 B.n444 B.n81 10.6151
R887 B.n445 B.n444 10.6151
R888 B.n446 B.n445 10.6151
R889 B.n446 B.n79 10.6151
R890 B.n450 B.n79 10.6151
R891 B.n451 B.n450 10.6151
R892 B.n452 B.n451 10.6151
R893 B.n452 B.n77 10.6151
R894 B.n456 B.n77 10.6151
R895 B.n457 B.n456 10.6151
R896 B.n458 B.n457 10.6151
R897 B.n458 B.n75 10.6151
R898 B.n462 B.n75 10.6151
R899 B.n463 B.n462 10.6151
R900 B.n464 B.n463 10.6151
R901 B.n464 B.n73 10.6151
R902 B.n468 B.n73 10.6151
R903 B.n469 B.n468 10.6151
R904 B.n470 B.n469 10.6151
R905 B.n224 B.n155 10.6151
R906 B.n225 B.n224 10.6151
R907 B.n226 B.n225 10.6151
R908 B.n226 B.n153 10.6151
R909 B.n230 B.n153 10.6151
R910 B.n231 B.n230 10.6151
R911 B.n232 B.n231 10.6151
R912 B.n232 B.n151 10.6151
R913 B.n236 B.n151 10.6151
R914 B.n237 B.n236 10.6151
R915 B.n238 B.n237 10.6151
R916 B.n238 B.n149 10.6151
R917 B.n242 B.n149 10.6151
R918 B.n243 B.n242 10.6151
R919 B.n244 B.n243 10.6151
R920 B.n244 B.n147 10.6151
R921 B.n248 B.n147 10.6151
R922 B.n249 B.n248 10.6151
R923 B.n250 B.n249 10.6151
R924 B.n250 B.n145 10.6151
R925 B.n254 B.n145 10.6151
R926 B.n255 B.n254 10.6151
R927 B.n256 B.n255 10.6151
R928 B.n256 B.n143 10.6151
R929 B.n260 B.n143 10.6151
R930 B.n261 B.n260 10.6151
R931 B.n262 B.n261 10.6151
R932 B.n262 B.n141 10.6151
R933 B.n266 B.n141 10.6151
R934 B.n267 B.n266 10.6151
R935 B.n268 B.n267 10.6151
R936 B.n268 B.n139 10.6151
R937 B.n272 B.n139 10.6151
R938 B.n273 B.n272 10.6151
R939 B.n274 B.n273 10.6151
R940 B.n274 B.n137 10.6151
R941 B.n278 B.n137 10.6151
R942 B.n279 B.n278 10.6151
R943 B.n280 B.n279 10.6151
R944 B.n280 B.n135 10.6151
R945 B.n284 B.n135 10.6151
R946 B.n285 B.n284 10.6151
R947 B.n287 B.n131 10.6151
R948 B.n291 B.n131 10.6151
R949 B.n292 B.n291 10.6151
R950 B.n293 B.n292 10.6151
R951 B.n293 B.n129 10.6151
R952 B.n297 B.n129 10.6151
R953 B.n298 B.n297 10.6151
R954 B.n302 B.n298 10.6151
R955 B.n306 B.n127 10.6151
R956 B.n307 B.n306 10.6151
R957 B.n308 B.n307 10.6151
R958 B.n308 B.n125 10.6151
R959 B.n312 B.n125 10.6151
R960 B.n313 B.n312 10.6151
R961 B.n314 B.n313 10.6151
R962 B.n314 B.n123 10.6151
R963 B.n318 B.n123 10.6151
R964 B.n319 B.n318 10.6151
R965 B.n320 B.n319 10.6151
R966 B.n320 B.n121 10.6151
R967 B.n324 B.n121 10.6151
R968 B.n325 B.n324 10.6151
R969 B.n326 B.n325 10.6151
R970 B.n326 B.n119 10.6151
R971 B.n330 B.n119 10.6151
R972 B.n331 B.n330 10.6151
R973 B.n332 B.n331 10.6151
R974 B.n332 B.n117 10.6151
R975 B.n336 B.n117 10.6151
R976 B.n337 B.n336 10.6151
R977 B.n338 B.n337 10.6151
R978 B.n338 B.n115 10.6151
R979 B.n342 B.n115 10.6151
R980 B.n343 B.n342 10.6151
R981 B.n344 B.n343 10.6151
R982 B.n344 B.n113 10.6151
R983 B.n348 B.n113 10.6151
R984 B.n349 B.n348 10.6151
R985 B.n350 B.n349 10.6151
R986 B.n350 B.n111 10.6151
R987 B.n354 B.n111 10.6151
R988 B.n355 B.n354 10.6151
R989 B.n356 B.n355 10.6151
R990 B.n356 B.n109 10.6151
R991 B.n360 B.n109 10.6151
R992 B.n361 B.n360 10.6151
R993 B.n362 B.n361 10.6151
R994 B.n362 B.n107 10.6151
R995 B.n366 B.n107 10.6151
R996 B.n367 B.n366 10.6151
R997 B.n220 B.n219 10.6151
R998 B.n219 B.n218 10.6151
R999 B.n218 B.n157 10.6151
R1000 B.n214 B.n157 10.6151
R1001 B.n214 B.n213 10.6151
R1002 B.n213 B.n212 10.6151
R1003 B.n212 B.n159 10.6151
R1004 B.n208 B.n159 10.6151
R1005 B.n208 B.n207 10.6151
R1006 B.n207 B.n206 10.6151
R1007 B.n206 B.n161 10.6151
R1008 B.n202 B.n161 10.6151
R1009 B.n202 B.n201 10.6151
R1010 B.n201 B.n200 10.6151
R1011 B.n200 B.n163 10.6151
R1012 B.n196 B.n163 10.6151
R1013 B.n196 B.n195 10.6151
R1014 B.n195 B.n194 10.6151
R1015 B.n194 B.n165 10.6151
R1016 B.n190 B.n165 10.6151
R1017 B.n190 B.n189 10.6151
R1018 B.n189 B.n188 10.6151
R1019 B.n188 B.n167 10.6151
R1020 B.n184 B.n167 10.6151
R1021 B.n184 B.n183 10.6151
R1022 B.n183 B.n182 10.6151
R1023 B.n182 B.n169 10.6151
R1024 B.n178 B.n169 10.6151
R1025 B.n178 B.n177 10.6151
R1026 B.n177 B.n176 10.6151
R1027 B.n176 B.n171 10.6151
R1028 B.n172 B.n171 10.6151
R1029 B.n172 B.n0 10.6151
R1030 B.n663 B.n1 10.6151
R1031 B.n663 B.n662 10.6151
R1032 B.n662 B.n661 10.6151
R1033 B.n661 B.n4 10.6151
R1034 B.n657 B.n4 10.6151
R1035 B.n657 B.n656 10.6151
R1036 B.n656 B.n655 10.6151
R1037 B.n655 B.n6 10.6151
R1038 B.n651 B.n6 10.6151
R1039 B.n651 B.n650 10.6151
R1040 B.n650 B.n649 10.6151
R1041 B.n649 B.n8 10.6151
R1042 B.n645 B.n8 10.6151
R1043 B.n645 B.n644 10.6151
R1044 B.n644 B.n643 10.6151
R1045 B.n643 B.n10 10.6151
R1046 B.n639 B.n10 10.6151
R1047 B.n639 B.n638 10.6151
R1048 B.n638 B.n637 10.6151
R1049 B.n637 B.n12 10.6151
R1050 B.n633 B.n12 10.6151
R1051 B.n633 B.n632 10.6151
R1052 B.n632 B.n631 10.6151
R1053 B.n631 B.n14 10.6151
R1054 B.n627 B.n14 10.6151
R1055 B.n627 B.n626 10.6151
R1056 B.n626 B.n625 10.6151
R1057 B.n625 B.n16 10.6151
R1058 B.n621 B.n16 10.6151
R1059 B.n621 B.n620 10.6151
R1060 B.n620 B.n619 10.6151
R1061 B.n619 B.n18 10.6151
R1062 B.n615 B.n18 10.6151
R1063 B.n549 B.n44 6.5566
R1064 B.n537 B.n536 6.5566
R1065 B.n287 B.n286 6.5566
R1066 B.n302 B.n301 6.5566
R1067 B.n44 B.n40 4.05904
R1068 B.n536 B.n535 4.05904
R1069 B.n286 B.n285 4.05904
R1070 B.n301 B.n127 4.05904
R1071 B.n667 B.n0 2.81026
R1072 B.n667 B.n1 2.81026
C0 VP VDD2 0.395714f
C1 w_n2740_n3454# VDD2 1.52792f
C2 VDD2 VN 4.91261f
C3 B VP 1.7022f
C4 B w_n2740_n3454# 9.39157f
C5 B VN 1.1175f
C6 VDD1 VP 5.15843f
C7 VDD1 w_n2740_n3454# 1.47136f
C8 VDD1 VN 0.149154f
C9 VTAIL VDD2 5.56687f
C10 B VTAIL 5.09693f
C11 VDD1 VTAIL 5.51253f
C12 VP w_n2740_n3454# 4.99646f
C13 VP VN 6.28264f
C14 w_n2740_n3454# VN 4.64417f
C15 B VDD2 1.3284f
C16 VDD1 VDD2 1.02554f
C17 VP VTAIL 4.82243f
C18 VDD1 B 1.27594f
C19 w_n2740_n3454# VTAIL 4.07238f
C20 VTAIL VN 4.80833f
C21 VDD2 VSUBS 0.968145f
C22 VDD1 VSUBS 5.82397f
C23 VTAIL VSUBS 1.235958f
C24 VN VSUBS 5.46595f
C25 VP VSUBS 2.310885f
C26 B VSUBS 4.330704f
C27 w_n2740_n3454# VSUBS 0.116428p
C28 B.n0 VSUBS 0.004203f
C29 B.n1 VSUBS 0.004203f
C30 B.n2 VSUBS 0.006647f
C31 B.n3 VSUBS 0.006647f
C32 B.n4 VSUBS 0.006647f
C33 B.n5 VSUBS 0.006647f
C34 B.n6 VSUBS 0.006647f
C35 B.n7 VSUBS 0.006647f
C36 B.n8 VSUBS 0.006647f
C37 B.n9 VSUBS 0.006647f
C38 B.n10 VSUBS 0.006647f
C39 B.n11 VSUBS 0.006647f
C40 B.n12 VSUBS 0.006647f
C41 B.n13 VSUBS 0.006647f
C42 B.n14 VSUBS 0.006647f
C43 B.n15 VSUBS 0.006647f
C44 B.n16 VSUBS 0.006647f
C45 B.n17 VSUBS 0.006647f
C46 B.n18 VSUBS 0.006647f
C47 B.n19 VSUBS 0.016843f
C48 B.n20 VSUBS 0.006647f
C49 B.n21 VSUBS 0.006647f
C50 B.n22 VSUBS 0.006647f
C51 B.n23 VSUBS 0.006647f
C52 B.n24 VSUBS 0.006647f
C53 B.n25 VSUBS 0.006647f
C54 B.n26 VSUBS 0.006647f
C55 B.n27 VSUBS 0.006647f
C56 B.n28 VSUBS 0.006647f
C57 B.n29 VSUBS 0.006647f
C58 B.n30 VSUBS 0.006647f
C59 B.n31 VSUBS 0.006647f
C60 B.n32 VSUBS 0.006647f
C61 B.n33 VSUBS 0.006647f
C62 B.n34 VSUBS 0.006647f
C63 B.n35 VSUBS 0.006647f
C64 B.n36 VSUBS 0.006647f
C65 B.n37 VSUBS 0.006647f
C66 B.n38 VSUBS 0.006647f
C67 B.n39 VSUBS 0.006647f
C68 B.n40 VSUBS 0.004594f
C69 B.n41 VSUBS 0.006647f
C70 B.t11 VSUBS 0.386066f
C71 B.t10 VSUBS 0.4061f
C72 B.t9 VSUBS 1.40613f
C73 B.n42 VSUBS 0.213827f
C74 B.n43 VSUBS 0.068272f
C75 B.n44 VSUBS 0.0154f
C76 B.n45 VSUBS 0.006647f
C77 B.n46 VSUBS 0.006647f
C78 B.n47 VSUBS 0.006647f
C79 B.n48 VSUBS 0.006647f
C80 B.t5 VSUBS 0.386058f
C81 B.t4 VSUBS 0.406093f
C82 B.t3 VSUBS 1.40613f
C83 B.n49 VSUBS 0.213834f
C84 B.n50 VSUBS 0.06828f
C85 B.n51 VSUBS 0.006647f
C86 B.n52 VSUBS 0.006647f
C87 B.n53 VSUBS 0.006647f
C88 B.n54 VSUBS 0.006647f
C89 B.n55 VSUBS 0.006647f
C90 B.n56 VSUBS 0.006647f
C91 B.n57 VSUBS 0.006647f
C92 B.n58 VSUBS 0.006647f
C93 B.n59 VSUBS 0.006647f
C94 B.n60 VSUBS 0.006647f
C95 B.n61 VSUBS 0.006647f
C96 B.n62 VSUBS 0.006647f
C97 B.n63 VSUBS 0.006647f
C98 B.n64 VSUBS 0.006647f
C99 B.n65 VSUBS 0.006647f
C100 B.n66 VSUBS 0.006647f
C101 B.n67 VSUBS 0.006647f
C102 B.n68 VSUBS 0.006647f
C103 B.n69 VSUBS 0.006647f
C104 B.n70 VSUBS 0.006647f
C105 B.n71 VSUBS 0.016125f
C106 B.n72 VSUBS 0.006647f
C107 B.n73 VSUBS 0.006647f
C108 B.n74 VSUBS 0.006647f
C109 B.n75 VSUBS 0.006647f
C110 B.n76 VSUBS 0.006647f
C111 B.n77 VSUBS 0.006647f
C112 B.n78 VSUBS 0.006647f
C113 B.n79 VSUBS 0.006647f
C114 B.n80 VSUBS 0.006647f
C115 B.n81 VSUBS 0.006647f
C116 B.n82 VSUBS 0.006647f
C117 B.n83 VSUBS 0.006647f
C118 B.n84 VSUBS 0.006647f
C119 B.n85 VSUBS 0.006647f
C120 B.n86 VSUBS 0.006647f
C121 B.n87 VSUBS 0.006647f
C122 B.n88 VSUBS 0.006647f
C123 B.n89 VSUBS 0.006647f
C124 B.n90 VSUBS 0.006647f
C125 B.n91 VSUBS 0.006647f
C126 B.n92 VSUBS 0.006647f
C127 B.n93 VSUBS 0.006647f
C128 B.n94 VSUBS 0.006647f
C129 B.n95 VSUBS 0.006647f
C130 B.n96 VSUBS 0.006647f
C131 B.n97 VSUBS 0.006647f
C132 B.n98 VSUBS 0.006647f
C133 B.n99 VSUBS 0.006647f
C134 B.n100 VSUBS 0.006647f
C135 B.n101 VSUBS 0.006647f
C136 B.n102 VSUBS 0.006647f
C137 B.n103 VSUBS 0.006647f
C138 B.n104 VSUBS 0.006647f
C139 B.n105 VSUBS 0.006647f
C140 B.n106 VSUBS 0.016843f
C141 B.n107 VSUBS 0.006647f
C142 B.n108 VSUBS 0.006647f
C143 B.n109 VSUBS 0.006647f
C144 B.n110 VSUBS 0.006647f
C145 B.n111 VSUBS 0.006647f
C146 B.n112 VSUBS 0.006647f
C147 B.n113 VSUBS 0.006647f
C148 B.n114 VSUBS 0.006647f
C149 B.n115 VSUBS 0.006647f
C150 B.n116 VSUBS 0.006647f
C151 B.n117 VSUBS 0.006647f
C152 B.n118 VSUBS 0.006647f
C153 B.n119 VSUBS 0.006647f
C154 B.n120 VSUBS 0.006647f
C155 B.n121 VSUBS 0.006647f
C156 B.n122 VSUBS 0.006647f
C157 B.n123 VSUBS 0.006647f
C158 B.n124 VSUBS 0.006647f
C159 B.n125 VSUBS 0.006647f
C160 B.n126 VSUBS 0.006647f
C161 B.n127 VSUBS 0.004594f
C162 B.n128 VSUBS 0.006647f
C163 B.n129 VSUBS 0.006647f
C164 B.n130 VSUBS 0.006647f
C165 B.n131 VSUBS 0.006647f
C166 B.n132 VSUBS 0.006647f
C167 B.t1 VSUBS 0.386066f
C168 B.t2 VSUBS 0.4061f
C169 B.t0 VSUBS 1.40613f
C170 B.n133 VSUBS 0.213827f
C171 B.n134 VSUBS 0.068272f
C172 B.n135 VSUBS 0.006647f
C173 B.n136 VSUBS 0.006647f
C174 B.n137 VSUBS 0.006647f
C175 B.n138 VSUBS 0.006647f
C176 B.n139 VSUBS 0.006647f
C177 B.n140 VSUBS 0.006647f
C178 B.n141 VSUBS 0.006647f
C179 B.n142 VSUBS 0.006647f
C180 B.n143 VSUBS 0.006647f
C181 B.n144 VSUBS 0.006647f
C182 B.n145 VSUBS 0.006647f
C183 B.n146 VSUBS 0.006647f
C184 B.n147 VSUBS 0.006647f
C185 B.n148 VSUBS 0.006647f
C186 B.n149 VSUBS 0.006647f
C187 B.n150 VSUBS 0.006647f
C188 B.n151 VSUBS 0.006647f
C189 B.n152 VSUBS 0.006647f
C190 B.n153 VSUBS 0.006647f
C191 B.n154 VSUBS 0.006647f
C192 B.n155 VSUBS 0.016843f
C193 B.n156 VSUBS 0.006647f
C194 B.n157 VSUBS 0.006647f
C195 B.n158 VSUBS 0.006647f
C196 B.n159 VSUBS 0.006647f
C197 B.n160 VSUBS 0.006647f
C198 B.n161 VSUBS 0.006647f
C199 B.n162 VSUBS 0.006647f
C200 B.n163 VSUBS 0.006647f
C201 B.n164 VSUBS 0.006647f
C202 B.n165 VSUBS 0.006647f
C203 B.n166 VSUBS 0.006647f
C204 B.n167 VSUBS 0.006647f
C205 B.n168 VSUBS 0.006647f
C206 B.n169 VSUBS 0.006647f
C207 B.n170 VSUBS 0.006647f
C208 B.n171 VSUBS 0.006647f
C209 B.n172 VSUBS 0.006647f
C210 B.n173 VSUBS 0.006647f
C211 B.n174 VSUBS 0.006647f
C212 B.n175 VSUBS 0.006647f
C213 B.n176 VSUBS 0.006647f
C214 B.n177 VSUBS 0.006647f
C215 B.n178 VSUBS 0.006647f
C216 B.n179 VSUBS 0.006647f
C217 B.n180 VSUBS 0.006647f
C218 B.n181 VSUBS 0.006647f
C219 B.n182 VSUBS 0.006647f
C220 B.n183 VSUBS 0.006647f
C221 B.n184 VSUBS 0.006647f
C222 B.n185 VSUBS 0.006647f
C223 B.n186 VSUBS 0.006647f
C224 B.n187 VSUBS 0.006647f
C225 B.n188 VSUBS 0.006647f
C226 B.n189 VSUBS 0.006647f
C227 B.n190 VSUBS 0.006647f
C228 B.n191 VSUBS 0.006647f
C229 B.n192 VSUBS 0.006647f
C230 B.n193 VSUBS 0.006647f
C231 B.n194 VSUBS 0.006647f
C232 B.n195 VSUBS 0.006647f
C233 B.n196 VSUBS 0.006647f
C234 B.n197 VSUBS 0.006647f
C235 B.n198 VSUBS 0.006647f
C236 B.n199 VSUBS 0.006647f
C237 B.n200 VSUBS 0.006647f
C238 B.n201 VSUBS 0.006647f
C239 B.n202 VSUBS 0.006647f
C240 B.n203 VSUBS 0.006647f
C241 B.n204 VSUBS 0.006647f
C242 B.n205 VSUBS 0.006647f
C243 B.n206 VSUBS 0.006647f
C244 B.n207 VSUBS 0.006647f
C245 B.n208 VSUBS 0.006647f
C246 B.n209 VSUBS 0.006647f
C247 B.n210 VSUBS 0.006647f
C248 B.n211 VSUBS 0.006647f
C249 B.n212 VSUBS 0.006647f
C250 B.n213 VSUBS 0.006647f
C251 B.n214 VSUBS 0.006647f
C252 B.n215 VSUBS 0.006647f
C253 B.n216 VSUBS 0.006647f
C254 B.n217 VSUBS 0.006647f
C255 B.n218 VSUBS 0.006647f
C256 B.n219 VSUBS 0.006647f
C257 B.n220 VSUBS 0.016195f
C258 B.n221 VSUBS 0.016195f
C259 B.n222 VSUBS 0.016843f
C260 B.n223 VSUBS 0.006647f
C261 B.n224 VSUBS 0.006647f
C262 B.n225 VSUBS 0.006647f
C263 B.n226 VSUBS 0.006647f
C264 B.n227 VSUBS 0.006647f
C265 B.n228 VSUBS 0.006647f
C266 B.n229 VSUBS 0.006647f
C267 B.n230 VSUBS 0.006647f
C268 B.n231 VSUBS 0.006647f
C269 B.n232 VSUBS 0.006647f
C270 B.n233 VSUBS 0.006647f
C271 B.n234 VSUBS 0.006647f
C272 B.n235 VSUBS 0.006647f
C273 B.n236 VSUBS 0.006647f
C274 B.n237 VSUBS 0.006647f
C275 B.n238 VSUBS 0.006647f
C276 B.n239 VSUBS 0.006647f
C277 B.n240 VSUBS 0.006647f
C278 B.n241 VSUBS 0.006647f
C279 B.n242 VSUBS 0.006647f
C280 B.n243 VSUBS 0.006647f
C281 B.n244 VSUBS 0.006647f
C282 B.n245 VSUBS 0.006647f
C283 B.n246 VSUBS 0.006647f
C284 B.n247 VSUBS 0.006647f
C285 B.n248 VSUBS 0.006647f
C286 B.n249 VSUBS 0.006647f
C287 B.n250 VSUBS 0.006647f
C288 B.n251 VSUBS 0.006647f
C289 B.n252 VSUBS 0.006647f
C290 B.n253 VSUBS 0.006647f
C291 B.n254 VSUBS 0.006647f
C292 B.n255 VSUBS 0.006647f
C293 B.n256 VSUBS 0.006647f
C294 B.n257 VSUBS 0.006647f
C295 B.n258 VSUBS 0.006647f
C296 B.n259 VSUBS 0.006647f
C297 B.n260 VSUBS 0.006647f
C298 B.n261 VSUBS 0.006647f
C299 B.n262 VSUBS 0.006647f
C300 B.n263 VSUBS 0.006647f
C301 B.n264 VSUBS 0.006647f
C302 B.n265 VSUBS 0.006647f
C303 B.n266 VSUBS 0.006647f
C304 B.n267 VSUBS 0.006647f
C305 B.n268 VSUBS 0.006647f
C306 B.n269 VSUBS 0.006647f
C307 B.n270 VSUBS 0.006647f
C308 B.n271 VSUBS 0.006647f
C309 B.n272 VSUBS 0.006647f
C310 B.n273 VSUBS 0.006647f
C311 B.n274 VSUBS 0.006647f
C312 B.n275 VSUBS 0.006647f
C313 B.n276 VSUBS 0.006647f
C314 B.n277 VSUBS 0.006647f
C315 B.n278 VSUBS 0.006647f
C316 B.n279 VSUBS 0.006647f
C317 B.n280 VSUBS 0.006647f
C318 B.n281 VSUBS 0.006647f
C319 B.n282 VSUBS 0.006647f
C320 B.n283 VSUBS 0.006647f
C321 B.n284 VSUBS 0.006647f
C322 B.n285 VSUBS 0.004594f
C323 B.n286 VSUBS 0.0154f
C324 B.n287 VSUBS 0.005376f
C325 B.n288 VSUBS 0.006647f
C326 B.n289 VSUBS 0.006647f
C327 B.n290 VSUBS 0.006647f
C328 B.n291 VSUBS 0.006647f
C329 B.n292 VSUBS 0.006647f
C330 B.n293 VSUBS 0.006647f
C331 B.n294 VSUBS 0.006647f
C332 B.n295 VSUBS 0.006647f
C333 B.n296 VSUBS 0.006647f
C334 B.n297 VSUBS 0.006647f
C335 B.n298 VSUBS 0.006647f
C336 B.t7 VSUBS 0.386058f
C337 B.t8 VSUBS 0.406093f
C338 B.t6 VSUBS 1.40613f
C339 B.n299 VSUBS 0.213834f
C340 B.n300 VSUBS 0.06828f
C341 B.n301 VSUBS 0.0154f
C342 B.n302 VSUBS 0.005376f
C343 B.n303 VSUBS 0.006647f
C344 B.n304 VSUBS 0.006647f
C345 B.n305 VSUBS 0.006647f
C346 B.n306 VSUBS 0.006647f
C347 B.n307 VSUBS 0.006647f
C348 B.n308 VSUBS 0.006647f
C349 B.n309 VSUBS 0.006647f
C350 B.n310 VSUBS 0.006647f
C351 B.n311 VSUBS 0.006647f
C352 B.n312 VSUBS 0.006647f
C353 B.n313 VSUBS 0.006647f
C354 B.n314 VSUBS 0.006647f
C355 B.n315 VSUBS 0.006647f
C356 B.n316 VSUBS 0.006647f
C357 B.n317 VSUBS 0.006647f
C358 B.n318 VSUBS 0.006647f
C359 B.n319 VSUBS 0.006647f
C360 B.n320 VSUBS 0.006647f
C361 B.n321 VSUBS 0.006647f
C362 B.n322 VSUBS 0.006647f
C363 B.n323 VSUBS 0.006647f
C364 B.n324 VSUBS 0.006647f
C365 B.n325 VSUBS 0.006647f
C366 B.n326 VSUBS 0.006647f
C367 B.n327 VSUBS 0.006647f
C368 B.n328 VSUBS 0.006647f
C369 B.n329 VSUBS 0.006647f
C370 B.n330 VSUBS 0.006647f
C371 B.n331 VSUBS 0.006647f
C372 B.n332 VSUBS 0.006647f
C373 B.n333 VSUBS 0.006647f
C374 B.n334 VSUBS 0.006647f
C375 B.n335 VSUBS 0.006647f
C376 B.n336 VSUBS 0.006647f
C377 B.n337 VSUBS 0.006647f
C378 B.n338 VSUBS 0.006647f
C379 B.n339 VSUBS 0.006647f
C380 B.n340 VSUBS 0.006647f
C381 B.n341 VSUBS 0.006647f
C382 B.n342 VSUBS 0.006647f
C383 B.n343 VSUBS 0.006647f
C384 B.n344 VSUBS 0.006647f
C385 B.n345 VSUBS 0.006647f
C386 B.n346 VSUBS 0.006647f
C387 B.n347 VSUBS 0.006647f
C388 B.n348 VSUBS 0.006647f
C389 B.n349 VSUBS 0.006647f
C390 B.n350 VSUBS 0.006647f
C391 B.n351 VSUBS 0.006647f
C392 B.n352 VSUBS 0.006647f
C393 B.n353 VSUBS 0.006647f
C394 B.n354 VSUBS 0.006647f
C395 B.n355 VSUBS 0.006647f
C396 B.n356 VSUBS 0.006647f
C397 B.n357 VSUBS 0.006647f
C398 B.n358 VSUBS 0.006647f
C399 B.n359 VSUBS 0.006647f
C400 B.n360 VSUBS 0.006647f
C401 B.n361 VSUBS 0.006647f
C402 B.n362 VSUBS 0.006647f
C403 B.n363 VSUBS 0.006647f
C404 B.n364 VSUBS 0.006647f
C405 B.n365 VSUBS 0.006647f
C406 B.n366 VSUBS 0.006647f
C407 B.n367 VSUBS 0.016843f
C408 B.n368 VSUBS 0.016195f
C409 B.n369 VSUBS 0.016195f
C410 B.n370 VSUBS 0.006647f
C411 B.n371 VSUBS 0.006647f
C412 B.n372 VSUBS 0.006647f
C413 B.n373 VSUBS 0.006647f
C414 B.n374 VSUBS 0.006647f
C415 B.n375 VSUBS 0.006647f
C416 B.n376 VSUBS 0.006647f
C417 B.n377 VSUBS 0.006647f
C418 B.n378 VSUBS 0.006647f
C419 B.n379 VSUBS 0.006647f
C420 B.n380 VSUBS 0.006647f
C421 B.n381 VSUBS 0.006647f
C422 B.n382 VSUBS 0.006647f
C423 B.n383 VSUBS 0.006647f
C424 B.n384 VSUBS 0.006647f
C425 B.n385 VSUBS 0.006647f
C426 B.n386 VSUBS 0.006647f
C427 B.n387 VSUBS 0.006647f
C428 B.n388 VSUBS 0.006647f
C429 B.n389 VSUBS 0.006647f
C430 B.n390 VSUBS 0.006647f
C431 B.n391 VSUBS 0.006647f
C432 B.n392 VSUBS 0.006647f
C433 B.n393 VSUBS 0.006647f
C434 B.n394 VSUBS 0.006647f
C435 B.n395 VSUBS 0.006647f
C436 B.n396 VSUBS 0.006647f
C437 B.n397 VSUBS 0.006647f
C438 B.n398 VSUBS 0.006647f
C439 B.n399 VSUBS 0.006647f
C440 B.n400 VSUBS 0.006647f
C441 B.n401 VSUBS 0.006647f
C442 B.n402 VSUBS 0.006647f
C443 B.n403 VSUBS 0.006647f
C444 B.n404 VSUBS 0.006647f
C445 B.n405 VSUBS 0.006647f
C446 B.n406 VSUBS 0.006647f
C447 B.n407 VSUBS 0.006647f
C448 B.n408 VSUBS 0.006647f
C449 B.n409 VSUBS 0.006647f
C450 B.n410 VSUBS 0.006647f
C451 B.n411 VSUBS 0.006647f
C452 B.n412 VSUBS 0.006647f
C453 B.n413 VSUBS 0.006647f
C454 B.n414 VSUBS 0.006647f
C455 B.n415 VSUBS 0.006647f
C456 B.n416 VSUBS 0.006647f
C457 B.n417 VSUBS 0.006647f
C458 B.n418 VSUBS 0.006647f
C459 B.n419 VSUBS 0.006647f
C460 B.n420 VSUBS 0.006647f
C461 B.n421 VSUBS 0.006647f
C462 B.n422 VSUBS 0.006647f
C463 B.n423 VSUBS 0.006647f
C464 B.n424 VSUBS 0.006647f
C465 B.n425 VSUBS 0.006647f
C466 B.n426 VSUBS 0.006647f
C467 B.n427 VSUBS 0.006647f
C468 B.n428 VSUBS 0.006647f
C469 B.n429 VSUBS 0.006647f
C470 B.n430 VSUBS 0.006647f
C471 B.n431 VSUBS 0.006647f
C472 B.n432 VSUBS 0.006647f
C473 B.n433 VSUBS 0.006647f
C474 B.n434 VSUBS 0.006647f
C475 B.n435 VSUBS 0.006647f
C476 B.n436 VSUBS 0.006647f
C477 B.n437 VSUBS 0.006647f
C478 B.n438 VSUBS 0.006647f
C479 B.n439 VSUBS 0.006647f
C480 B.n440 VSUBS 0.006647f
C481 B.n441 VSUBS 0.006647f
C482 B.n442 VSUBS 0.006647f
C483 B.n443 VSUBS 0.006647f
C484 B.n444 VSUBS 0.006647f
C485 B.n445 VSUBS 0.006647f
C486 B.n446 VSUBS 0.006647f
C487 B.n447 VSUBS 0.006647f
C488 B.n448 VSUBS 0.006647f
C489 B.n449 VSUBS 0.006647f
C490 B.n450 VSUBS 0.006647f
C491 B.n451 VSUBS 0.006647f
C492 B.n452 VSUBS 0.006647f
C493 B.n453 VSUBS 0.006647f
C494 B.n454 VSUBS 0.006647f
C495 B.n455 VSUBS 0.006647f
C496 B.n456 VSUBS 0.006647f
C497 B.n457 VSUBS 0.006647f
C498 B.n458 VSUBS 0.006647f
C499 B.n459 VSUBS 0.006647f
C500 B.n460 VSUBS 0.006647f
C501 B.n461 VSUBS 0.006647f
C502 B.n462 VSUBS 0.006647f
C503 B.n463 VSUBS 0.006647f
C504 B.n464 VSUBS 0.006647f
C505 B.n465 VSUBS 0.006647f
C506 B.n466 VSUBS 0.006647f
C507 B.n467 VSUBS 0.006647f
C508 B.n468 VSUBS 0.006647f
C509 B.n469 VSUBS 0.006647f
C510 B.n470 VSUBS 0.016913f
C511 B.n471 VSUBS 0.016195f
C512 B.n472 VSUBS 0.016843f
C513 B.n473 VSUBS 0.006647f
C514 B.n474 VSUBS 0.006647f
C515 B.n475 VSUBS 0.006647f
C516 B.n476 VSUBS 0.006647f
C517 B.n477 VSUBS 0.006647f
C518 B.n478 VSUBS 0.006647f
C519 B.n479 VSUBS 0.006647f
C520 B.n480 VSUBS 0.006647f
C521 B.n481 VSUBS 0.006647f
C522 B.n482 VSUBS 0.006647f
C523 B.n483 VSUBS 0.006647f
C524 B.n484 VSUBS 0.006647f
C525 B.n485 VSUBS 0.006647f
C526 B.n486 VSUBS 0.006647f
C527 B.n487 VSUBS 0.006647f
C528 B.n488 VSUBS 0.006647f
C529 B.n489 VSUBS 0.006647f
C530 B.n490 VSUBS 0.006647f
C531 B.n491 VSUBS 0.006647f
C532 B.n492 VSUBS 0.006647f
C533 B.n493 VSUBS 0.006647f
C534 B.n494 VSUBS 0.006647f
C535 B.n495 VSUBS 0.006647f
C536 B.n496 VSUBS 0.006647f
C537 B.n497 VSUBS 0.006647f
C538 B.n498 VSUBS 0.006647f
C539 B.n499 VSUBS 0.006647f
C540 B.n500 VSUBS 0.006647f
C541 B.n501 VSUBS 0.006647f
C542 B.n502 VSUBS 0.006647f
C543 B.n503 VSUBS 0.006647f
C544 B.n504 VSUBS 0.006647f
C545 B.n505 VSUBS 0.006647f
C546 B.n506 VSUBS 0.006647f
C547 B.n507 VSUBS 0.006647f
C548 B.n508 VSUBS 0.006647f
C549 B.n509 VSUBS 0.006647f
C550 B.n510 VSUBS 0.006647f
C551 B.n511 VSUBS 0.006647f
C552 B.n512 VSUBS 0.006647f
C553 B.n513 VSUBS 0.006647f
C554 B.n514 VSUBS 0.006647f
C555 B.n515 VSUBS 0.006647f
C556 B.n516 VSUBS 0.006647f
C557 B.n517 VSUBS 0.006647f
C558 B.n518 VSUBS 0.006647f
C559 B.n519 VSUBS 0.006647f
C560 B.n520 VSUBS 0.006647f
C561 B.n521 VSUBS 0.006647f
C562 B.n522 VSUBS 0.006647f
C563 B.n523 VSUBS 0.006647f
C564 B.n524 VSUBS 0.006647f
C565 B.n525 VSUBS 0.006647f
C566 B.n526 VSUBS 0.006647f
C567 B.n527 VSUBS 0.006647f
C568 B.n528 VSUBS 0.006647f
C569 B.n529 VSUBS 0.006647f
C570 B.n530 VSUBS 0.006647f
C571 B.n531 VSUBS 0.006647f
C572 B.n532 VSUBS 0.006647f
C573 B.n533 VSUBS 0.006647f
C574 B.n534 VSUBS 0.006647f
C575 B.n535 VSUBS 0.004594f
C576 B.n536 VSUBS 0.0154f
C577 B.n537 VSUBS 0.005376f
C578 B.n538 VSUBS 0.006647f
C579 B.n539 VSUBS 0.006647f
C580 B.n540 VSUBS 0.006647f
C581 B.n541 VSUBS 0.006647f
C582 B.n542 VSUBS 0.006647f
C583 B.n543 VSUBS 0.006647f
C584 B.n544 VSUBS 0.006647f
C585 B.n545 VSUBS 0.006647f
C586 B.n546 VSUBS 0.006647f
C587 B.n547 VSUBS 0.006647f
C588 B.n548 VSUBS 0.006647f
C589 B.n549 VSUBS 0.005376f
C590 B.n550 VSUBS 0.006647f
C591 B.n551 VSUBS 0.006647f
C592 B.n552 VSUBS 0.006647f
C593 B.n553 VSUBS 0.006647f
C594 B.n554 VSUBS 0.006647f
C595 B.n555 VSUBS 0.006647f
C596 B.n556 VSUBS 0.006647f
C597 B.n557 VSUBS 0.006647f
C598 B.n558 VSUBS 0.006647f
C599 B.n559 VSUBS 0.006647f
C600 B.n560 VSUBS 0.006647f
C601 B.n561 VSUBS 0.006647f
C602 B.n562 VSUBS 0.006647f
C603 B.n563 VSUBS 0.006647f
C604 B.n564 VSUBS 0.006647f
C605 B.n565 VSUBS 0.006647f
C606 B.n566 VSUBS 0.006647f
C607 B.n567 VSUBS 0.006647f
C608 B.n568 VSUBS 0.006647f
C609 B.n569 VSUBS 0.006647f
C610 B.n570 VSUBS 0.006647f
C611 B.n571 VSUBS 0.006647f
C612 B.n572 VSUBS 0.006647f
C613 B.n573 VSUBS 0.006647f
C614 B.n574 VSUBS 0.006647f
C615 B.n575 VSUBS 0.006647f
C616 B.n576 VSUBS 0.006647f
C617 B.n577 VSUBS 0.006647f
C618 B.n578 VSUBS 0.006647f
C619 B.n579 VSUBS 0.006647f
C620 B.n580 VSUBS 0.006647f
C621 B.n581 VSUBS 0.006647f
C622 B.n582 VSUBS 0.006647f
C623 B.n583 VSUBS 0.006647f
C624 B.n584 VSUBS 0.006647f
C625 B.n585 VSUBS 0.006647f
C626 B.n586 VSUBS 0.006647f
C627 B.n587 VSUBS 0.006647f
C628 B.n588 VSUBS 0.006647f
C629 B.n589 VSUBS 0.006647f
C630 B.n590 VSUBS 0.006647f
C631 B.n591 VSUBS 0.006647f
C632 B.n592 VSUBS 0.006647f
C633 B.n593 VSUBS 0.006647f
C634 B.n594 VSUBS 0.006647f
C635 B.n595 VSUBS 0.006647f
C636 B.n596 VSUBS 0.006647f
C637 B.n597 VSUBS 0.006647f
C638 B.n598 VSUBS 0.006647f
C639 B.n599 VSUBS 0.006647f
C640 B.n600 VSUBS 0.006647f
C641 B.n601 VSUBS 0.006647f
C642 B.n602 VSUBS 0.006647f
C643 B.n603 VSUBS 0.006647f
C644 B.n604 VSUBS 0.006647f
C645 B.n605 VSUBS 0.006647f
C646 B.n606 VSUBS 0.006647f
C647 B.n607 VSUBS 0.006647f
C648 B.n608 VSUBS 0.006647f
C649 B.n609 VSUBS 0.006647f
C650 B.n610 VSUBS 0.006647f
C651 B.n611 VSUBS 0.006647f
C652 B.n612 VSUBS 0.006647f
C653 B.n613 VSUBS 0.006647f
C654 B.n614 VSUBS 0.016843f
C655 B.n615 VSUBS 0.016195f
C656 B.n616 VSUBS 0.016195f
C657 B.n617 VSUBS 0.006647f
C658 B.n618 VSUBS 0.006647f
C659 B.n619 VSUBS 0.006647f
C660 B.n620 VSUBS 0.006647f
C661 B.n621 VSUBS 0.006647f
C662 B.n622 VSUBS 0.006647f
C663 B.n623 VSUBS 0.006647f
C664 B.n624 VSUBS 0.006647f
C665 B.n625 VSUBS 0.006647f
C666 B.n626 VSUBS 0.006647f
C667 B.n627 VSUBS 0.006647f
C668 B.n628 VSUBS 0.006647f
C669 B.n629 VSUBS 0.006647f
C670 B.n630 VSUBS 0.006647f
C671 B.n631 VSUBS 0.006647f
C672 B.n632 VSUBS 0.006647f
C673 B.n633 VSUBS 0.006647f
C674 B.n634 VSUBS 0.006647f
C675 B.n635 VSUBS 0.006647f
C676 B.n636 VSUBS 0.006647f
C677 B.n637 VSUBS 0.006647f
C678 B.n638 VSUBS 0.006647f
C679 B.n639 VSUBS 0.006647f
C680 B.n640 VSUBS 0.006647f
C681 B.n641 VSUBS 0.006647f
C682 B.n642 VSUBS 0.006647f
C683 B.n643 VSUBS 0.006647f
C684 B.n644 VSUBS 0.006647f
C685 B.n645 VSUBS 0.006647f
C686 B.n646 VSUBS 0.006647f
C687 B.n647 VSUBS 0.006647f
C688 B.n648 VSUBS 0.006647f
C689 B.n649 VSUBS 0.006647f
C690 B.n650 VSUBS 0.006647f
C691 B.n651 VSUBS 0.006647f
C692 B.n652 VSUBS 0.006647f
C693 B.n653 VSUBS 0.006647f
C694 B.n654 VSUBS 0.006647f
C695 B.n655 VSUBS 0.006647f
C696 B.n656 VSUBS 0.006647f
C697 B.n657 VSUBS 0.006647f
C698 B.n658 VSUBS 0.006647f
C699 B.n659 VSUBS 0.006647f
C700 B.n660 VSUBS 0.006647f
C701 B.n661 VSUBS 0.006647f
C702 B.n662 VSUBS 0.006647f
C703 B.n663 VSUBS 0.006647f
C704 B.n664 VSUBS 0.006647f
C705 B.n665 VSUBS 0.006647f
C706 B.n666 VSUBS 0.006647f
C707 B.n667 VSUBS 0.01505f
C708 VDD2.t1 VSUBS 0.263784f
C709 VDD2.t3 VSUBS 0.263784f
C710 VDD2.n0 VSUBS 2.79914f
C711 VDD2.t0 VSUBS 0.263784f
C712 VDD2.t2 VSUBS 0.263784f
C713 VDD2.n1 VSUBS 2.06615f
C714 VDD2.n2 VSUBS 4.35373f
C715 VN.t2 VSUBS 3.17497f
C716 VN.t0 VSUBS 3.16881f
C717 VN.n0 VSUBS 2.00711f
C718 VN.t1 VSUBS 3.17497f
C719 VN.t3 VSUBS 3.16881f
C720 VN.n1 VSUBS 3.78181f
C721 VTAIL.t1 VSUBS 2.21894f
C722 VTAIL.n0 VSUBS 0.780544f
C723 VTAIL.t4 VSUBS 2.21894f
C724 VTAIL.n1 VSUBS 0.872713f
C725 VTAIL.t5 VSUBS 2.21894f
C726 VTAIL.n2 VSUBS 2.1644f
C727 VTAIL.t7 VSUBS 2.21896f
C728 VTAIL.n3 VSUBS 2.16438f
C729 VTAIL.t0 VSUBS 2.21896f
C730 VTAIL.n4 VSUBS 0.872697f
C731 VTAIL.t6 VSUBS 2.21896f
C732 VTAIL.n5 VSUBS 0.872697f
C733 VTAIL.t3 VSUBS 2.21894f
C734 VTAIL.n6 VSUBS 2.1644f
C735 VTAIL.t2 VSUBS 2.21894f
C736 VTAIL.n7 VSUBS 2.06339f
C737 VDD1.t3 VSUBS 0.266293f
C738 VDD1.t1 VSUBS 0.266293f
C739 VDD1.n0 VSUBS 2.08641f
C740 VDD1.t0 VSUBS 0.266293f
C741 VDD1.t2 VSUBS 0.266293f
C742 VDD1.n1 VSUBS 2.85153f
C743 VP.n0 VSUBS 0.044281f
C744 VP.t2 VSUBS 2.98317f
C745 VP.n1 VSUBS 0.049031f
C746 VP.n2 VSUBS 0.033587f
C747 VP.t1 VSUBS 2.98317f
C748 VP.n3 VSUBS 1.1683f
C749 VP.t3 VSUBS 3.28375f
C750 VP.t0 VSUBS 3.29013f
C751 VP.n4 VSUBS 3.90134f
C752 VP.n5 VSUBS 1.8853f
C753 VP.n6 VSUBS 0.044281f
C754 VP.n7 VSUBS 0.045598f
C755 VP.n8 VSUBS 0.062597f
C756 VP.n9 VSUBS 0.049031f
C757 VP.n10 VSUBS 0.033587f
C758 VP.n11 VSUBS 0.033587f
C759 VP.n12 VSUBS 0.033587f
C760 VP.n13 VSUBS 0.062597f
C761 VP.n14 VSUBS 0.045598f
C762 VP.n15 VSUBS 1.1683f
C763 VP.n16 VSUBS 0.053931f
.ends

