* NGSPICE file created from diff_pair_sample_1737.ext - technology: sky130A

.subckt diff_pair_sample_1737 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t5 VP.t0 VTAIL.t6 w_n1706_n1414# sky130_fd_pr__pfet_01v8 ad=0.8697 pd=5.24 as=0.36795 ps=2.56 w=2.23 l=0.59
X1 VTAIL.t1 VN.t0 VDD2.t5 w_n1706_n1414# sky130_fd_pr__pfet_01v8 ad=0.36795 pd=2.56 as=0.36795 ps=2.56 w=2.23 l=0.59
X2 B.t11 B.t9 B.t10 w_n1706_n1414# sky130_fd_pr__pfet_01v8 ad=0.8697 pd=5.24 as=0 ps=0 w=2.23 l=0.59
X3 VDD2.t4 VN.t1 VTAIL.t5 w_n1706_n1414# sky130_fd_pr__pfet_01v8 ad=0.8697 pd=5.24 as=0.36795 ps=2.56 w=2.23 l=0.59
X4 VDD1.t4 VP.t1 VTAIL.t7 w_n1706_n1414# sky130_fd_pr__pfet_01v8 ad=0.8697 pd=5.24 as=0.36795 ps=2.56 w=2.23 l=0.59
X5 VDD1.t3 VP.t2 VTAIL.t8 w_n1706_n1414# sky130_fd_pr__pfet_01v8 ad=0.36795 pd=2.56 as=0.8697 ps=5.24 w=2.23 l=0.59
X6 VDD2.t3 VN.t2 VTAIL.t2 w_n1706_n1414# sky130_fd_pr__pfet_01v8 ad=0.36795 pd=2.56 as=0.8697 ps=5.24 w=2.23 l=0.59
X7 B.t8 B.t6 B.t7 w_n1706_n1414# sky130_fd_pr__pfet_01v8 ad=0.8697 pd=5.24 as=0 ps=0 w=2.23 l=0.59
X8 VTAIL.t4 VN.t3 VDD2.t2 w_n1706_n1414# sky130_fd_pr__pfet_01v8 ad=0.36795 pd=2.56 as=0.36795 ps=2.56 w=2.23 l=0.59
X9 B.t5 B.t3 B.t4 w_n1706_n1414# sky130_fd_pr__pfet_01v8 ad=0.8697 pd=5.24 as=0 ps=0 w=2.23 l=0.59
X10 VDD2.t1 VN.t4 VTAIL.t3 w_n1706_n1414# sky130_fd_pr__pfet_01v8 ad=0.36795 pd=2.56 as=0.8697 ps=5.24 w=2.23 l=0.59
X11 VDD1.t2 VP.t3 VTAIL.t9 w_n1706_n1414# sky130_fd_pr__pfet_01v8 ad=0.36795 pd=2.56 as=0.8697 ps=5.24 w=2.23 l=0.59
X12 VDD2.t0 VN.t5 VTAIL.t0 w_n1706_n1414# sky130_fd_pr__pfet_01v8 ad=0.8697 pd=5.24 as=0.36795 ps=2.56 w=2.23 l=0.59
X13 VTAIL.t10 VP.t4 VDD1.t1 w_n1706_n1414# sky130_fd_pr__pfet_01v8 ad=0.36795 pd=2.56 as=0.36795 ps=2.56 w=2.23 l=0.59
X14 VTAIL.t11 VP.t5 VDD1.t0 w_n1706_n1414# sky130_fd_pr__pfet_01v8 ad=0.36795 pd=2.56 as=0.36795 ps=2.56 w=2.23 l=0.59
X15 B.t2 B.t0 B.t1 w_n1706_n1414# sky130_fd_pr__pfet_01v8 ad=0.8697 pd=5.24 as=0 ps=0 w=2.23 l=0.59
R0 VP.n1 VP.t1 184.901
R1 VP.n9 VP.n8 161.3
R2 VP.n4 VP.n3 161.3
R3 VP.n6 VP.n5 161.3
R4 VP.n6 VP.t0 158.081
R5 VP.n7 VP.t4 158.081
R6 VP.n8 VP.t3 158.081
R7 VP.n3 VP.t2 158.081
R8 VP.n2 VP.t5 158.081
R9 VP.n7 VP.n0 80.6037
R10 VP.n7 VP.n6 48.2005
R11 VP.n8 VP.n7 48.2005
R12 VP.n3 VP.n2 48.2005
R13 VP.n4 VP.n1 45.1367
R14 VP.n5 VP.n4 33.4475
R15 VP.n2 VP.n1 13.3799
R16 VP.n5 VP.n0 0.285035
R17 VP.n9 VP.n0 0.285035
R18 VP VP.n9 0.0516364
R19 VTAIL.n11 VTAIL.t3 172.422
R20 VTAIL.n2 VTAIL.t9 172.422
R21 VTAIL.n10 VTAIL.t8 172.422
R22 VTAIL.n7 VTAIL.t2 172.422
R23 VTAIL.n9 VTAIL.n8 157.845
R24 VTAIL.n6 VTAIL.n5 157.845
R25 VTAIL.n1 VTAIL.n0 157.845
R26 VTAIL.n4 VTAIL.n3 157.845
R27 VTAIL.n6 VTAIL.n4 15.8755
R28 VTAIL.n11 VTAIL.n10 15.0824
R29 VTAIL.n0 VTAIL.t5 14.5767
R30 VTAIL.n0 VTAIL.t4 14.5767
R31 VTAIL.n3 VTAIL.t6 14.5767
R32 VTAIL.n3 VTAIL.t10 14.5767
R33 VTAIL.n8 VTAIL.t7 14.5767
R34 VTAIL.n8 VTAIL.t11 14.5767
R35 VTAIL.n5 VTAIL.t0 14.5767
R36 VTAIL.n5 VTAIL.t1 14.5767
R37 VTAIL.n9 VTAIL.n7 0.866879
R38 VTAIL.n2 VTAIL.n1 0.866879
R39 VTAIL.n7 VTAIL.n6 0.793603
R40 VTAIL.n10 VTAIL.n9 0.793603
R41 VTAIL.n4 VTAIL.n2 0.793603
R42 VTAIL VTAIL.n11 0.537138
R43 VTAIL VTAIL.n1 0.256966
R44 VDD1 VDD1.t4 189.754
R45 VDD1.n1 VDD1.t5 189.639
R46 VDD1.n1 VDD1.n0 174.667
R47 VDD1.n3 VDD1.n2 174.524
R48 VDD1.n3 VDD1.n1 29.1949
R49 VDD1.n2 VDD1.t0 14.5767
R50 VDD1.n2 VDD1.t3 14.5767
R51 VDD1.n0 VDD1.t1 14.5767
R52 VDD1.n0 VDD1.t2 14.5767
R53 VDD1 VDD1.n3 0.140586
R54 VN.n0 VN.t1 184.901
R55 VN.n4 VN.t2 184.901
R56 VN.n3 VN.n2 161.3
R57 VN.n7 VN.n6 161.3
R58 VN.n1 VN.t3 158.081
R59 VN.n2 VN.t4 158.081
R60 VN.n5 VN.t0 158.081
R61 VN.n6 VN.t5 158.081
R62 VN.n2 VN.n1 48.2005
R63 VN.n6 VN.n5 48.2005
R64 VN.n7 VN.n4 45.1367
R65 VN.n3 VN.n0 45.1367
R66 VN VN.n7 33.8282
R67 VN.n5 VN.n4 13.3799
R68 VN.n1 VN.n0 13.3799
R69 VN VN.n3 0.0516364
R70 VDD2.n1 VDD2.t4 189.639
R71 VDD2.n2 VDD2.t0 189.101
R72 VDD2.n1 VDD2.n0 174.667
R73 VDD2 VDD2.n3 174.665
R74 VDD2.n2 VDD2.n1 28.2153
R75 VDD2.n3 VDD2.t5 14.5767
R76 VDD2.n3 VDD2.t3 14.5767
R77 VDD2.n0 VDD2.t2 14.5767
R78 VDD2.n0 VDD2.t1 14.5767
R79 VDD2 VDD2.n2 0.653517
R80 B.n224 B.n33 585
R81 B.n226 B.n225 585
R82 B.n227 B.n32 585
R83 B.n229 B.n228 585
R84 B.n230 B.n31 585
R85 B.n232 B.n231 585
R86 B.n233 B.n30 585
R87 B.n235 B.n234 585
R88 B.n236 B.n29 585
R89 B.n238 B.n237 585
R90 B.n239 B.n28 585
R91 B.n241 B.n240 585
R92 B.n242 B.n25 585
R93 B.n245 B.n244 585
R94 B.n246 B.n24 585
R95 B.n248 B.n247 585
R96 B.n249 B.n23 585
R97 B.n251 B.n250 585
R98 B.n252 B.n22 585
R99 B.n254 B.n253 585
R100 B.n255 B.n21 585
R101 B.n257 B.n256 585
R102 B.n259 B.n258 585
R103 B.n260 B.n17 585
R104 B.n262 B.n261 585
R105 B.n263 B.n16 585
R106 B.n265 B.n264 585
R107 B.n266 B.n15 585
R108 B.n268 B.n267 585
R109 B.n269 B.n14 585
R110 B.n271 B.n270 585
R111 B.n272 B.n13 585
R112 B.n274 B.n273 585
R113 B.n275 B.n12 585
R114 B.n277 B.n276 585
R115 B.n223 B.n222 585
R116 B.n221 B.n34 585
R117 B.n220 B.n219 585
R118 B.n218 B.n35 585
R119 B.n217 B.n216 585
R120 B.n215 B.n36 585
R121 B.n214 B.n213 585
R122 B.n212 B.n37 585
R123 B.n211 B.n210 585
R124 B.n209 B.n38 585
R125 B.n208 B.n207 585
R126 B.n206 B.n39 585
R127 B.n205 B.n204 585
R128 B.n203 B.n40 585
R129 B.n202 B.n201 585
R130 B.n200 B.n41 585
R131 B.n199 B.n198 585
R132 B.n197 B.n42 585
R133 B.n196 B.n195 585
R134 B.n194 B.n43 585
R135 B.n193 B.n192 585
R136 B.n191 B.n44 585
R137 B.n190 B.n189 585
R138 B.n188 B.n45 585
R139 B.n187 B.n186 585
R140 B.n185 B.n46 585
R141 B.n184 B.n183 585
R142 B.n182 B.n47 585
R143 B.n181 B.n180 585
R144 B.n179 B.n48 585
R145 B.n178 B.n177 585
R146 B.n176 B.n49 585
R147 B.n175 B.n174 585
R148 B.n173 B.n50 585
R149 B.n172 B.n171 585
R150 B.n170 B.n51 585
R151 B.n169 B.n168 585
R152 B.n167 B.n52 585
R153 B.n166 B.n165 585
R154 B.n112 B.n111 585
R155 B.n113 B.n74 585
R156 B.n115 B.n114 585
R157 B.n116 B.n73 585
R158 B.n118 B.n117 585
R159 B.n119 B.n72 585
R160 B.n121 B.n120 585
R161 B.n122 B.n71 585
R162 B.n124 B.n123 585
R163 B.n125 B.n70 585
R164 B.n127 B.n126 585
R165 B.n128 B.n69 585
R166 B.n130 B.n129 585
R167 B.n132 B.n131 585
R168 B.n133 B.n65 585
R169 B.n135 B.n134 585
R170 B.n136 B.n64 585
R171 B.n138 B.n137 585
R172 B.n139 B.n63 585
R173 B.n141 B.n140 585
R174 B.n142 B.n62 585
R175 B.n144 B.n143 585
R176 B.n146 B.n59 585
R177 B.n148 B.n147 585
R178 B.n149 B.n58 585
R179 B.n151 B.n150 585
R180 B.n152 B.n57 585
R181 B.n154 B.n153 585
R182 B.n155 B.n56 585
R183 B.n157 B.n156 585
R184 B.n158 B.n55 585
R185 B.n160 B.n159 585
R186 B.n161 B.n54 585
R187 B.n163 B.n162 585
R188 B.n164 B.n53 585
R189 B.n110 B.n75 585
R190 B.n109 B.n108 585
R191 B.n107 B.n76 585
R192 B.n106 B.n105 585
R193 B.n104 B.n77 585
R194 B.n103 B.n102 585
R195 B.n101 B.n78 585
R196 B.n100 B.n99 585
R197 B.n98 B.n79 585
R198 B.n97 B.n96 585
R199 B.n95 B.n80 585
R200 B.n94 B.n93 585
R201 B.n92 B.n81 585
R202 B.n91 B.n90 585
R203 B.n89 B.n82 585
R204 B.n88 B.n87 585
R205 B.n86 B.n83 585
R206 B.n85 B.n84 585
R207 B.n2 B.n0 585
R208 B.n305 B.n1 585
R209 B.n304 B.n303 585
R210 B.n302 B.n3 585
R211 B.n301 B.n300 585
R212 B.n299 B.n4 585
R213 B.n298 B.n297 585
R214 B.n296 B.n5 585
R215 B.n295 B.n294 585
R216 B.n293 B.n6 585
R217 B.n292 B.n291 585
R218 B.n290 B.n7 585
R219 B.n289 B.n288 585
R220 B.n287 B.n8 585
R221 B.n286 B.n285 585
R222 B.n284 B.n9 585
R223 B.n283 B.n282 585
R224 B.n281 B.n10 585
R225 B.n280 B.n279 585
R226 B.n278 B.n11 585
R227 B.n307 B.n306 585
R228 B.n112 B.n75 516.524
R229 B.n276 B.n11 516.524
R230 B.n166 B.n53 516.524
R231 B.n222 B.n33 516.524
R232 B.n60 B.t3 295.659
R233 B.n66 B.t0 295.659
R234 B.n18 B.t6 295.659
R235 B.n26 B.t9 295.659
R236 B.n60 B.t5 191.073
R237 B.n26 B.t10 191.073
R238 B.n66 B.t2 191.073
R239 B.n18 B.t7 191.073
R240 B.n61 B.t4 173.232
R241 B.n27 B.t11 173.232
R242 B.n67 B.t1 173.231
R243 B.n19 B.t8 173.231
R244 B.n108 B.n75 163.367
R245 B.n108 B.n107 163.367
R246 B.n107 B.n106 163.367
R247 B.n106 B.n77 163.367
R248 B.n102 B.n77 163.367
R249 B.n102 B.n101 163.367
R250 B.n101 B.n100 163.367
R251 B.n100 B.n79 163.367
R252 B.n96 B.n79 163.367
R253 B.n96 B.n95 163.367
R254 B.n95 B.n94 163.367
R255 B.n94 B.n81 163.367
R256 B.n90 B.n81 163.367
R257 B.n90 B.n89 163.367
R258 B.n89 B.n88 163.367
R259 B.n88 B.n83 163.367
R260 B.n84 B.n83 163.367
R261 B.n84 B.n2 163.367
R262 B.n306 B.n2 163.367
R263 B.n306 B.n305 163.367
R264 B.n305 B.n304 163.367
R265 B.n304 B.n3 163.367
R266 B.n300 B.n3 163.367
R267 B.n300 B.n299 163.367
R268 B.n299 B.n298 163.367
R269 B.n298 B.n5 163.367
R270 B.n294 B.n5 163.367
R271 B.n294 B.n293 163.367
R272 B.n293 B.n292 163.367
R273 B.n292 B.n7 163.367
R274 B.n288 B.n7 163.367
R275 B.n288 B.n287 163.367
R276 B.n287 B.n286 163.367
R277 B.n286 B.n9 163.367
R278 B.n282 B.n9 163.367
R279 B.n282 B.n281 163.367
R280 B.n281 B.n280 163.367
R281 B.n280 B.n11 163.367
R282 B.n113 B.n112 163.367
R283 B.n114 B.n113 163.367
R284 B.n114 B.n73 163.367
R285 B.n118 B.n73 163.367
R286 B.n119 B.n118 163.367
R287 B.n120 B.n119 163.367
R288 B.n120 B.n71 163.367
R289 B.n124 B.n71 163.367
R290 B.n125 B.n124 163.367
R291 B.n126 B.n125 163.367
R292 B.n126 B.n69 163.367
R293 B.n130 B.n69 163.367
R294 B.n131 B.n130 163.367
R295 B.n131 B.n65 163.367
R296 B.n135 B.n65 163.367
R297 B.n136 B.n135 163.367
R298 B.n137 B.n136 163.367
R299 B.n137 B.n63 163.367
R300 B.n141 B.n63 163.367
R301 B.n142 B.n141 163.367
R302 B.n143 B.n142 163.367
R303 B.n143 B.n59 163.367
R304 B.n148 B.n59 163.367
R305 B.n149 B.n148 163.367
R306 B.n150 B.n149 163.367
R307 B.n150 B.n57 163.367
R308 B.n154 B.n57 163.367
R309 B.n155 B.n154 163.367
R310 B.n156 B.n155 163.367
R311 B.n156 B.n55 163.367
R312 B.n160 B.n55 163.367
R313 B.n161 B.n160 163.367
R314 B.n162 B.n161 163.367
R315 B.n162 B.n53 163.367
R316 B.n167 B.n166 163.367
R317 B.n168 B.n167 163.367
R318 B.n168 B.n51 163.367
R319 B.n172 B.n51 163.367
R320 B.n173 B.n172 163.367
R321 B.n174 B.n173 163.367
R322 B.n174 B.n49 163.367
R323 B.n178 B.n49 163.367
R324 B.n179 B.n178 163.367
R325 B.n180 B.n179 163.367
R326 B.n180 B.n47 163.367
R327 B.n184 B.n47 163.367
R328 B.n185 B.n184 163.367
R329 B.n186 B.n185 163.367
R330 B.n186 B.n45 163.367
R331 B.n190 B.n45 163.367
R332 B.n191 B.n190 163.367
R333 B.n192 B.n191 163.367
R334 B.n192 B.n43 163.367
R335 B.n196 B.n43 163.367
R336 B.n197 B.n196 163.367
R337 B.n198 B.n197 163.367
R338 B.n198 B.n41 163.367
R339 B.n202 B.n41 163.367
R340 B.n203 B.n202 163.367
R341 B.n204 B.n203 163.367
R342 B.n204 B.n39 163.367
R343 B.n208 B.n39 163.367
R344 B.n209 B.n208 163.367
R345 B.n210 B.n209 163.367
R346 B.n210 B.n37 163.367
R347 B.n214 B.n37 163.367
R348 B.n215 B.n214 163.367
R349 B.n216 B.n215 163.367
R350 B.n216 B.n35 163.367
R351 B.n220 B.n35 163.367
R352 B.n221 B.n220 163.367
R353 B.n222 B.n221 163.367
R354 B.n276 B.n275 163.367
R355 B.n275 B.n274 163.367
R356 B.n274 B.n13 163.367
R357 B.n270 B.n13 163.367
R358 B.n270 B.n269 163.367
R359 B.n269 B.n268 163.367
R360 B.n268 B.n15 163.367
R361 B.n264 B.n15 163.367
R362 B.n264 B.n263 163.367
R363 B.n263 B.n262 163.367
R364 B.n262 B.n17 163.367
R365 B.n258 B.n17 163.367
R366 B.n258 B.n257 163.367
R367 B.n257 B.n21 163.367
R368 B.n253 B.n21 163.367
R369 B.n253 B.n252 163.367
R370 B.n252 B.n251 163.367
R371 B.n251 B.n23 163.367
R372 B.n247 B.n23 163.367
R373 B.n247 B.n246 163.367
R374 B.n246 B.n245 163.367
R375 B.n245 B.n25 163.367
R376 B.n240 B.n25 163.367
R377 B.n240 B.n239 163.367
R378 B.n239 B.n238 163.367
R379 B.n238 B.n29 163.367
R380 B.n234 B.n29 163.367
R381 B.n234 B.n233 163.367
R382 B.n233 B.n232 163.367
R383 B.n232 B.n31 163.367
R384 B.n228 B.n31 163.367
R385 B.n228 B.n227 163.367
R386 B.n227 B.n226 163.367
R387 B.n226 B.n33 163.367
R388 B.n145 B.n61 59.5399
R389 B.n68 B.n67 59.5399
R390 B.n20 B.n19 59.5399
R391 B.n243 B.n27 59.5399
R392 B.n278 B.n277 33.5615
R393 B.n224 B.n223 33.5615
R394 B.n165 B.n164 33.5615
R395 B.n111 B.n110 33.5615
R396 B B.n307 18.0485
R397 B.n61 B.n60 17.8429
R398 B.n67 B.n66 17.8429
R399 B.n19 B.n18 17.8429
R400 B.n27 B.n26 17.8429
R401 B.n277 B.n12 10.6151
R402 B.n273 B.n12 10.6151
R403 B.n273 B.n272 10.6151
R404 B.n272 B.n271 10.6151
R405 B.n271 B.n14 10.6151
R406 B.n267 B.n14 10.6151
R407 B.n267 B.n266 10.6151
R408 B.n266 B.n265 10.6151
R409 B.n265 B.n16 10.6151
R410 B.n261 B.n16 10.6151
R411 B.n261 B.n260 10.6151
R412 B.n260 B.n259 10.6151
R413 B.n256 B.n255 10.6151
R414 B.n255 B.n254 10.6151
R415 B.n254 B.n22 10.6151
R416 B.n250 B.n22 10.6151
R417 B.n250 B.n249 10.6151
R418 B.n249 B.n248 10.6151
R419 B.n248 B.n24 10.6151
R420 B.n244 B.n24 10.6151
R421 B.n242 B.n241 10.6151
R422 B.n241 B.n28 10.6151
R423 B.n237 B.n28 10.6151
R424 B.n237 B.n236 10.6151
R425 B.n236 B.n235 10.6151
R426 B.n235 B.n30 10.6151
R427 B.n231 B.n30 10.6151
R428 B.n231 B.n230 10.6151
R429 B.n230 B.n229 10.6151
R430 B.n229 B.n32 10.6151
R431 B.n225 B.n32 10.6151
R432 B.n225 B.n224 10.6151
R433 B.n165 B.n52 10.6151
R434 B.n169 B.n52 10.6151
R435 B.n170 B.n169 10.6151
R436 B.n171 B.n170 10.6151
R437 B.n171 B.n50 10.6151
R438 B.n175 B.n50 10.6151
R439 B.n176 B.n175 10.6151
R440 B.n177 B.n176 10.6151
R441 B.n177 B.n48 10.6151
R442 B.n181 B.n48 10.6151
R443 B.n182 B.n181 10.6151
R444 B.n183 B.n182 10.6151
R445 B.n183 B.n46 10.6151
R446 B.n187 B.n46 10.6151
R447 B.n188 B.n187 10.6151
R448 B.n189 B.n188 10.6151
R449 B.n189 B.n44 10.6151
R450 B.n193 B.n44 10.6151
R451 B.n194 B.n193 10.6151
R452 B.n195 B.n194 10.6151
R453 B.n195 B.n42 10.6151
R454 B.n199 B.n42 10.6151
R455 B.n200 B.n199 10.6151
R456 B.n201 B.n200 10.6151
R457 B.n201 B.n40 10.6151
R458 B.n205 B.n40 10.6151
R459 B.n206 B.n205 10.6151
R460 B.n207 B.n206 10.6151
R461 B.n207 B.n38 10.6151
R462 B.n211 B.n38 10.6151
R463 B.n212 B.n211 10.6151
R464 B.n213 B.n212 10.6151
R465 B.n213 B.n36 10.6151
R466 B.n217 B.n36 10.6151
R467 B.n218 B.n217 10.6151
R468 B.n219 B.n218 10.6151
R469 B.n219 B.n34 10.6151
R470 B.n223 B.n34 10.6151
R471 B.n111 B.n74 10.6151
R472 B.n115 B.n74 10.6151
R473 B.n116 B.n115 10.6151
R474 B.n117 B.n116 10.6151
R475 B.n117 B.n72 10.6151
R476 B.n121 B.n72 10.6151
R477 B.n122 B.n121 10.6151
R478 B.n123 B.n122 10.6151
R479 B.n123 B.n70 10.6151
R480 B.n127 B.n70 10.6151
R481 B.n128 B.n127 10.6151
R482 B.n129 B.n128 10.6151
R483 B.n133 B.n132 10.6151
R484 B.n134 B.n133 10.6151
R485 B.n134 B.n64 10.6151
R486 B.n138 B.n64 10.6151
R487 B.n139 B.n138 10.6151
R488 B.n140 B.n139 10.6151
R489 B.n140 B.n62 10.6151
R490 B.n144 B.n62 10.6151
R491 B.n147 B.n146 10.6151
R492 B.n147 B.n58 10.6151
R493 B.n151 B.n58 10.6151
R494 B.n152 B.n151 10.6151
R495 B.n153 B.n152 10.6151
R496 B.n153 B.n56 10.6151
R497 B.n157 B.n56 10.6151
R498 B.n158 B.n157 10.6151
R499 B.n159 B.n158 10.6151
R500 B.n159 B.n54 10.6151
R501 B.n163 B.n54 10.6151
R502 B.n164 B.n163 10.6151
R503 B.n110 B.n109 10.6151
R504 B.n109 B.n76 10.6151
R505 B.n105 B.n76 10.6151
R506 B.n105 B.n104 10.6151
R507 B.n104 B.n103 10.6151
R508 B.n103 B.n78 10.6151
R509 B.n99 B.n78 10.6151
R510 B.n99 B.n98 10.6151
R511 B.n98 B.n97 10.6151
R512 B.n97 B.n80 10.6151
R513 B.n93 B.n80 10.6151
R514 B.n93 B.n92 10.6151
R515 B.n92 B.n91 10.6151
R516 B.n91 B.n82 10.6151
R517 B.n87 B.n82 10.6151
R518 B.n87 B.n86 10.6151
R519 B.n86 B.n85 10.6151
R520 B.n85 B.n0 10.6151
R521 B.n303 B.n1 10.6151
R522 B.n303 B.n302 10.6151
R523 B.n302 B.n301 10.6151
R524 B.n301 B.n4 10.6151
R525 B.n297 B.n4 10.6151
R526 B.n297 B.n296 10.6151
R527 B.n296 B.n295 10.6151
R528 B.n295 B.n6 10.6151
R529 B.n291 B.n6 10.6151
R530 B.n291 B.n290 10.6151
R531 B.n290 B.n289 10.6151
R532 B.n289 B.n8 10.6151
R533 B.n285 B.n8 10.6151
R534 B.n285 B.n284 10.6151
R535 B.n284 B.n283 10.6151
R536 B.n283 B.n10 10.6151
R537 B.n279 B.n10 10.6151
R538 B.n279 B.n278 10.6151
R539 B.n256 B.n20 6.5566
R540 B.n244 B.n243 6.5566
R541 B.n132 B.n68 6.5566
R542 B.n145 B.n144 6.5566
R543 B.n259 B.n20 4.05904
R544 B.n243 B.n242 4.05904
R545 B.n129 B.n68 4.05904
R546 B.n146 B.n145 4.05904
R547 B.n307 B.n0 2.81026
R548 B.n307 B.n1 2.81026
C0 VTAIL VN 1.14659f
C1 VP B 0.965352f
C2 VTAIL VDD1 3.42859f
C3 VTAIL w_n1706_n1414# 1.34083f
C4 VDD1 VN 0.154097f
C5 VN w_n1706_n1414# 2.52781f
C6 VTAIL VDD2 3.46727f
C7 VDD1 w_n1706_n1414# 1.05122f
C8 VDD2 VN 1.00533f
C9 VTAIL VP 1.1608f
C10 VTAIL B 0.898191f
C11 VDD2 VDD1 0.668928f
C12 VDD2 w_n1706_n1414# 1.07118f
C13 VN VP 3.17022f
C14 VN B 0.617236f
C15 VDD1 VP 1.14296f
C16 VDD1 B 0.819011f
C17 VP w_n1706_n1414# 2.73894f
C18 B w_n1706_n1414# 4.14934f
C19 VDD2 VP 0.293555f
C20 VDD2 B 0.845543f
C21 VDD2 VSUBS 0.709192f
C22 VDD1 VSUBS 0.930767f
C23 VTAIL VSUBS 0.302247f
C24 VN VSUBS 3.13192f
C25 VP VSUBS 0.926081f
C26 B VSUBS 1.734064f
C27 w_n1706_n1414# VSUBS 30.728498f
C28 B.n0 VSUBS 0.005374f
C29 B.n1 VSUBS 0.005374f
C30 B.n2 VSUBS 0.008498f
C31 B.n3 VSUBS 0.008498f
C32 B.n4 VSUBS 0.008498f
C33 B.n5 VSUBS 0.008498f
C34 B.n6 VSUBS 0.008498f
C35 B.n7 VSUBS 0.008498f
C36 B.n8 VSUBS 0.008498f
C37 B.n9 VSUBS 0.008498f
C38 B.n10 VSUBS 0.008498f
C39 B.n11 VSUBS 0.019971f
C40 B.n12 VSUBS 0.008498f
C41 B.n13 VSUBS 0.008498f
C42 B.n14 VSUBS 0.008498f
C43 B.n15 VSUBS 0.008498f
C44 B.n16 VSUBS 0.008498f
C45 B.n17 VSUBS 0.008498f
C46 B.t8 VSUBS 0.059841f
C47 B.t7 VSUBS 0.064604f
C48 B.t6 VSUBS 0.074495f
C49 B.n18 VSUBS 0.067851f
C50 B.n19 VSUBS 0.063132f
C51 B.n20 VSUBS 0.019689f
C52 B.n21 VSUBS 0.008498f
C53 B.n22 VSUBS 0.008498f
C54 B.n23 VSUBS 0.008498f
C55 B.n24 VSUBS 0.008498f
C56 B.n25 VSUBS 0.008498f
C57 B.t11 VSUBS 0.059841f
C58 B.t10 VSUBS 0.064604f
C59 B.t9 VSUBS 0.074495f
C60 B.n26 VSUBS 0.067851f
C61 B.n27 VSUBS 0.063132f
C62 B.n28 VSUBS 0.008498f
C63 B.n29 VSUBS 0.008498f
C64 B.n30 VSUBS 0.008498f
C65 B.n31 VSUBS 0.008498f
C66 B.n32 VSUBS 0.008498f
C67 B.n33 VSUBS 0.020519f
C68 B.n34 VSUBS 0.008498f
C69 B.n35 VSUBS 0.008498f
C70 B.n36 VSUBS 0.008498f
C71 B.n37 VSUBS 0.008498f
C72 B.n38 VSUBS 0.008498f
C73 B.n39 VSUBS 0.008498f
C74 B.n40 VSUBS 0.008498f
C75 B.n41 VSUBS 0.008498f
C76 B.n42 VSUBS 0.008498f
C77 B.n43 VSUBS 0.008498f
C78 B.n44 VSUBS 0.008498f
C79 B.n45 VSUBS 0.008498f
C80 B.n46 VSUBS 0.008498f
C81 B.n47 VSUBS 0.008498f
C82 B.n48 VSUBS 0.008498f
C83 B.n49 VSUBS 0.008498f
C84 B.n50 VSUBS 0.008498f
C85 B.n51 VSUBS 0.008498f
C86 B.n52 VSUBS 0.008498f
C87 B.n53 VSUBS 0.020519f
C88 B.n54 VSUBS 0.008498f
C89 B.n55 VSUBS 0.008498f
C90 B.n56 VSUBS 0.008498f
C91 B.n57 VSUBS 0.008498f
C92 B.n58 VSUBS 0.008498f
C93 B.n59 VSUBS 0.008498f
C94 B.t4 VSUBS 0.059841f
C95 B.t5 VSUBS 0.064604f
C96 B.t3 VSUBS 0.074495f
C97 B.n60 VSUBS 0.067851f
C98 B.n61 VSUBS 0.063132f
C99 B.n62 VSUBS 0.008498f
C100 B.n63 VSUBS 0.008498f
C101 B.n64 VSUBS 0.008498f
C102 B.n65 VSUBS 0.008498f
C103 B.t1 VSUBS 0.059841f
C104 B.t2 VSUBS 0.064604f
C105 B.t0 VSUBS 0.074495f
C106 B.n66 VSUBS 0.067851f
C107 B.n67 VSUBS 0.063132f
C108 B.n68 VSUBS 0.019689f
C109 B.n69 VSUBS 0.008498f
C110 B.n70 VSUBS 0.008498f
C111 B.n71 VSUBS 0.008498f
C112 B.n72 VSUBS 0.008498f
C113 B.n73 VSUBS 0.008498f
C114 B.n74 VSUBS 0.008498f
C115 B.n75 VSUBS 0.019971f
C116 B.n76 VSUBS 0.008498f
C117 B.n77 VSUBS 0.008498f
C118 B.n78 VSUBS 0.008498f
C119 B.n79 VSUBS 0.008498f
C120 B.n80 VSUBS 0.008498f
C121 B.n81 VSUBS 0.008498f
C122 B.n82 VSUBS 0.008498f
C123 B.n83 VSUBS 0.008498f
C124 B.n84 VSUBS 0.008498f
C125 B.n85 VSUBS 0.008498f
C126 B.n86 VSUBS 0.008498f
C127 B.n87 VSUBS 0.008498f
C128 B.n88 VSUBS 0.008498f
C129 B.n89 VSUBS 0.008498f
C130 B.n90 VSUBS 0.008498f
C131 B.n91 VSUBS 0.008498f
C132 B.n92 VSUBS 0.008498f
C133 B.n93 VSUBS 0.008498f
C134 B.n94 VSUBS 0.008498f
C135 B.n95 VSUBS 0.008498f
C136 B.n96 VSUBS 0.008498f
C137 B.n97 VSUBS 0.008498f
C138 B.n98 VSUBS 0.008498f
C139 B.n99 VSUBS 0.008498f
C140 B.n100 VSUBS 0.008498f
C141 B.n101 VSUBS 0.008498f
C142 B.n102 VSUBS 0.008498f
C143 B.n103 VSUBS 0.008498f
C144 B.n104 VSUBS 0.008498f
C145 B.n105 VSUBS 0.008498f
C146 B.n106 VSUBS 0.008498f
C147 B.n107 VSUBS 0.008498f
C148 B.n108 VSUBS 0.008498f
C149 B.n109 VSUBS 0.008498f
C150 B.n110 VSUBS 0.019971f
C151 B.n111 VSUBS 0.020519f
C152 B.n112 VSUBS 0.020519f
C153 B.n113 VSUBS 0.008498f
C154 B.n114 VSUBS 0.008498f
C155 B.n115 VSUBS 0.008498f
C156 B.n116 VSUBS 0.008498f
C157 B.n117 VSUBS 0.008498f
C158 B.n118 VSUBS 0.008498f
C159 B.n119 VSUBS 0.008498f
C160 B.n120 VSUBS 0.008498f
C161 B.n121 VSUBS 0.008498f
C162 B.n122 VSUBS 0.008498f
C163 B.n123 VSUBS 0.008498f
C164 B.n124 VSUBS 0.008498f
C165 B.n125 VSUBS 0.008498f
C166 B.n126 VSUBS 0.008498f
C167 B.n127 VSUBS 0.008498f
C168 B.n128 VSUBS 0.008498f
C169 B.n129 VSUBS 0.005873f
C170 B.n130 VSUBS 0.008498f
C171 B.n131 VSUBS 0.008498f
C172 B.n132 VSUBS 0.006873f
C173 B.n133 VSUBS 0.008498f
C174 B.n134 VSUBS 0.008498f
C175 B.n135 VSUBS 0.008498f
C176 B.n136 VSUBS 0.008498f
C177 B.n137 VSUBS 0.008498f
C178 B.n138 VSUBS 0.008498f
C179 B.n139 VSUBS 0.008498f
C180 B.n140 VSUBS 0.008498f
C181 B.n141 VSUBS 0.008498f
C182 B.n142 VSUBS 0.008498f
C183 B.n143 VSUBS 0.008498f
C184 B.n144 VSUBS 0.006873f
C185 B.n145 VSUBS 0.019689f
C186 B.n146 VSUBS 0.005873f
C187 B.n147 VSUBS 0.008498f
C188 B.n148 VSUBS 0.008498f
C189 B.n149 VSUBS 0.008498f
C190 B.n150 VSUBS 0.008498f
C191 B.n151 VSUBS 0.008498f
C192 B.n152 VSUBS 0.008498f
C193 B.n153 VSUBS 0.008498f
C194 B.n154 VSUBS 0.008498f
C195 B.n155 VSUBS 0.008498f
C196 B.n156 VSUBS 0.008498f
C197 B.n157 VSUBS 0.008498f
C198 B.n158 VSUBS 0.008498f
C199 B.n159 VSUBS 0.008498f
C200 B.n160 VSUBS 0.008498f
C201 B.n161 VSUBS 0.008498f
C202 B.n162 VSUBS 0.008498f
C203 B.n163 VSUBS 0.008498f
C204 B.n164 VSUBS 0.020519f
C205 B.n165 VSUBS 0.019971f
C206 B.n166 VSUBS 0.019971f
C207 B.n167 VSUBS 0.008498f
C208 B.n168 VSUBS 0.008498f
C209 B.n169 VSUBS 0.008498f
C210 B.n170 VSUBS 0.008498f
C211 B.n171 VSUBS 0.008498f
C212 B.n172 VSUBS 0.008498f
C213 B.n173 VSUBS 0.008498f
C214 B.n174 VSUBS 0.008498f
C215 B.n175 VSUBS 0.008498f
C216 B.n176 VSUBS 0.008498f
C217 B.n177 VSUBS 0.008498f
C218 B.n178 VSUBS 0.008498f
C219 B.n179 VSUBS 0.008498f
C220 B.n180 VSUBS 0.008498f
C221 B.n181 VSUBS 0.008498f
C222 B.n182 VSUBS 0.008498f
C223 B.n183 VSUBS 0.008498f
C224 B.n184 VSUBS 0.008498f
C225 B.n185 VSUBS 0.008498f
C226 B.n186 VSUBS 0.008498f
C227 B.n187 VSUBS 0.008498f
C228 B.n188 VSUBS 0.008498f
C229 B.n189 VSUBS 0.008498f
C230 B.n190 VSUBS 0.008498f
C231 B.n191 VSUBS 0.008498f
C232 B.n192 VSUBS 0.008498f
C233 B.n193 VSUBS 0.008498f
C234 B.n194 VSUBS 0.008498f
C235 B.n195 VSUBS 0.008498f
C236 B.n196 VSUBS 0.008498f
C237 B.n197 VSUBS 0.008498f
C238 B.n198 VSUBS 0.008498f
C239 B.n199 VSUBS 0.008498f
C240 B.n200 VSUBS 0.008498f
C241 B.n201 VSUBS 0.008498f
C242 B.n202 VSUBS 0.008498f
C243 B.n203 VSUBS 0.008498f
C244 B.n204 VSUBS 0.008498f
C245 B.n205 VSUBS 0.008498f
C246 B.n206 VSUBS 0.008498f
C247 B.n207 VSUBS 0.008498f
C248 B.n208 VSUBS 0.008498f
C249 B.n209 VSUBS 0.008498f
C250 B.n210 VSUBS 0.008498f
C251 B.n211 VSUBS 0.008498f
C252 B.n212 VSUBS 0.008498f
C253 B.n213 VSUBS 0.008498f
C254 B.n214 VSUBS 0.008498f
C255 B.n215 VSUBS 0.008498f
C256 B.n216 VSUBS 0.008498f
C257 B.n217 VSUBS 0.008498f
C258 B.n218 VSUBS 0.008498f
C259 B.n219 VSUBS 0.008498f
C260 B.n220 VSUBS 0.008498f
C261 B.n221 VSUBS 0.008498f
C262 B.n222 VSUBS 0.019971f
C263 B.n223 VSUBS 0.020948f
C264 B.n224 VSUBS 0.019542f
C265 B.n225 VSUBS 0.008498f
C266 B.n226 VSUBS 0.008498f
C267 B.n227 VSUBS 0.008498f
C268 B.n228 VSUBS 0.008498f
C269 B.n229 VSUBS 0.008498f
C270 B.n230 VSUBS 0.008498f
C271 B.n231 VSUBS 0.008498f
C272 B.n232 VSUBS 0.008498f
C273 B.n233 VSUBS 0.008498f
C274 B.n234 VSUBS 0.008498f
C275 B.n235 VSUBS 0.008498f
C276 B.n236 VSUBS 0.008498f
C277 B.n237 VSUBS 0.008498f
C278 B.n238 VSUBS 0.008498f
C279 B.n239 VSUBS 0.008498f
C280 B.n240 VSUBS 0.008498f
C281 B.n241 VSUBS 0.008498f
C282 B.n242 VSUBS 0.005873f
C283 B.n243 VSUBS 0.019689f
C284 B.n244 VSUBS 0.006873f
C285 B.n245 VSUBS 0.008498f
C286 B.n246 VSUBS 0.008498f
C287 B.n247 VSUBS 0.008498f
C288 B.n248 VSUBS 0.008498f
C289 B.n249 VSUBS 0.008498f
C290 B.n250 VSUBS 0.008498f
C291 B.n251 VSUBS 0.008498f
C292 B.n252 VSUBS 0.008498f
C293 B.n253 VSUBS 0.008498f
C294 B.n254 VSUBS 0.008498f
C295 B.n255 VSUBS 0.008498f
C296 B.n256 VSUBS 0.006873f
C297 B.n257 VSUBS 0.008498f
C298 B.n258 VSUBS 0.008498f
C299 B.n259 VSUBS 0.005873f
C300 B.n260 VSUBS 0.008498f
C301 B.n261 VSUBS 0.008498f
C302 B.n262 VSUBS 0.008498f
C303 B.n263 VSUBS 0.008498f
C304 B.n264 VSUBS 0.008498f
C305 B.n265 VSUBS 0.008498f
C306 B.n266 VSUBS 0.008498f
C307 B.n267 VSUBS 0.008498f
C308 B.n268 VSUBS 0.008498f
C309 B.n269 VSUBS 0.008498f
C310 B.n270 VSUBS 0.008498f
C311 B.n271 VSUBS 0.008498f
C312 B.n272 VSUBS 0.008498f
C313 B.n273 VSUBS 0.008498f
C314 B.n274 VSUBS 0.008498f
C315 B.n275 VSUBS 0.008498f
C316 B.n276 VSUBS 0.020519f
C317 B.n277 VSUBS 0.020519f
C318 B.n278 VSUBS 0.019971f
C319 B.n279 VSUBS 0.008498f
C320 B.n280 VSUBS 0.008498f
C321 B.n281 VSUBS 0.008498f
C322 B.n282 VSUBS 0.008498f
C323 B.n283 VSUBS 0.008498f
C324 B.n284 VSUBS 0.008498f
C325 B.n285 VSUBS 0.008498f
C326 B.n286 VSUBS 0.008498f
C327 B.n287 VSUBS 0.008498f
C328 B.n288 VSUBS 0.008498f
C329 B.n289 VSUBS 0.008498f
C330 B.n290 VSUBS 0.008498f
C331 B.n291 VSUBS 0.008498f
C332 B.n292 VSUBS 0.008498f
C333 B.n293 VSUBS 0.008498f
C334 B.n294 VSUBS 0.008498f
C335 B.n295 VSUBS 0.008498f
C336 B.n296 VSUBS 0.008498f
C337 B.n297 VSUBS 0.008498f
C338 B.n298 VSUBS 0.008498f
C339 B.n299 VSUBS 0.008498f
C340 B.n300 VSUBS 0.008498f
C341 B.n301 VSUBS 0.008498f
C342 B.n302 VSUBS 0.008498f
C343 B.n303 VSUBS 0.008498f
C344 B.n304 VSUBS 0.008498f
C345 B.n305 VSUBS 0.008498f
C346 B.n306 VSUBS 0.008498f
C347 B.n307 VSUBS 0.019242f
C348 VDD2.t4 VSUBS 0.226465f
C349 VDD2.t2 VSUBS 0.032961f
C350 VDD2.t1 VSUBS 0.032961f
C351 VDD2.n0 VSUBS 0.152139f
C352 VDD2.n1 VSUBS 1.17771f
C353 VDD2.t0 VSUBS 0.225709f
C354 VDD2.n2 VSUBS 1.11333f
C355 VDD2.t5 VSUBS 0.032961f
C356 VDD2.t3 VSUBS 0.032961f
C357 VDD2.n3 VSUBS 0.152132f
C358 VN.t1 VSUBS 0.241841f
C359 VN.n0 VSUBS 0.128102f
C360 VN.t3 VSUBS 0.220277f
C361 VN.n1 VSUBS 0.160879f
C362 VN.t4 VSUBS 0.220277f
C363 VN.n2 VSUBS 0.148506f
C364 VN.n3 VSUBS 0.219124f
C365 VN.t2 VSUBS 0.241841f
C366 VN.n4 VSUBS 0.128102f
C367 VN.t0 VSUBS 0.220277f
C368 VN.n5 VSUBS 0.160879f
C369 VN.t5 VSUBS 0.220277f
C370 VN.n6 VSUBS 0.148506f
C371 VN.n7 VSUBS 1.69886f
C372 VDD1.t4 VSUBS 0.215908f
C373 VDD1.t5 VSUBS 0.215737f
C374 VDD1.t1 VSUBS 0.031399f
C375 VDD1.t2 VSUBS 0.031399f
C376 VDD1.n0 VSUBS 0.144931f
C377 VDD1.n1 VSUBS 1.17186f
C378 VDD1.t0 VSUBS 0.031399f
C379 VDD1.t3 VSUBS 0.031399f
C380 VDD1.n2 VSUBS 0.144716f
C381 VDD1.n3 VSUBS 1.07721f
C382 VTAIL.t5 VSUBS 0.040129f
C383 VTAIL.t4 VSUBS 0.040129f
C384 VTAIL.n0 VSUBS 0.158481f
C385 VTAIL.n1 VSUBS 0.332736f
C386 VTAIL.t9 VSUBS 0.248666f
C387 VTAIL.n2 VSUBS 0.39137f
C388 VTAIL.t6 VSUBS 0.040129f
C389 VTAIL.t10 VSUBS 0.040129f
C390 VTAIL.n3 VSUBS 0.158481f
C391 VTAIL.n4 VSUBS 0.875321f
C392 VTAIL.t0 VSUBS 0.040129f
C393 VTAIL.t1 VSUBS 0.040129f
C394 VTAIL.n5 VSUBS 0.158482f
C395 VTAIL.n6 VSUBS 0.875321f
C396 VTAIL.t2 VSUBS 0.248667f
C397 VTAIL.n7 VSUBS 0.39137f
C398 VTAIL.t7 VSUBS 0.040129f
C399 VTAIL.t11 VSUBS 0.040129f
C400 VTAIL.n8 VSUBS 0.158482f
C401 VTAIL.n9 VSUBS 0.372112f
C402 VTAIL.t8 VSUBS 0.248666f
C403 VTAIL.n10 VSUBS 0.836384f
C404 VTAIL.t3 VSUBS 0.248666f
C405 VTAIL.n11 VSUBS 0.817565f
C406 VP.n0 VSUBS 0.076157f
C407 VP.t1 VSUBS 0.253739f
C408 VP.n1 VSUBS 0.134404f
C409 VP.t2 VSUBS 0.231114f
C410 VP.t5 VSUBS 0.231114f
C411 VP.n2 VSUBS 0.168793f
C412 VP.n3 VSUBS 0.155812f
C413 VP.n4 VSUBS 1.74428f
C414 VP.n5 VSUBS 1.63932f
C415 VP.t0 VSUBS 0.231114f
C416 VP.n6 VSUBS 0.155812f
C417 VP.t4 VSUBS 0.231114f
C418 VP.n7 VSUBS 0.168793f
C419 VP.t3 VSUBS 0.231114f
C420 VP.n8 VSUBS 0.155812f
C421 VP.n9 VSUBS 0.063462f
.ends

