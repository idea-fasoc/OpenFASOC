* NGSPICE file created from diff_pair_sample_0829.ext - technology: sky130A

.subckt diff_pair_sample_0829 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n1610_n1834# sky130_fd_pr__pfet_01v8 ad=1.6887 pd=9.44 as=0 ps=0 w=4.33 l=1.27
X1 VDD1.t1 VP.t0 VTAIL.t2 w_n1610_n1834# sky130_fd_pr__pfet_01v8 ad=1.6887 pd=9.44 as=1.6887 ps=9.44 w=4.33 l=1.27
X2 VDD2.t1 VN.t0 VTAIL.t0 w_n1610_n1834# sky130_fd_pr__pfet_01v8 ad=1.6887 pd=9.44 as=1.6887 ps=9.44 w=4.33 l=1.27
X3 VDD2.t0 VN.t1 VTAIL.t1 w_n1610_n1834# sky130_fd_pr__pfet_01v8 ad=1.6887 pd=9.44 as=1.6887 ps=9.44 w=4.33 l=1.27
X4 B.t8 B.t6 B.t7 w_n1610_n1834# sky130_fd_pr__pfet_01v8 ad=1.6887 pd=9.44 as=0 ps=0 w=4.33 l=1.27
X5 B.t5 B.t3 B.t4 w_n1610_n1834# sky130_fd_pr__pfet_01v8 ad=1.6887 pd=9.44 as=0 ps=0 w=4.33 l=1.27
X6 VDD1.t0 VP.t1 VTAIL.t3 w_n1610_n1834# sky130_fd_pr__pfet_01v8 ad=1.6887 pd=9.44 as=1.6887 ps=9.44 w=4.33 l=1.27
X7 B.t2 B.t0 B.t1 w_n1610_n1834# sky130_fd_pr__pfet_01v8 ad=1.6887 pd=9.44 as=0 ps=0 w=4.33 l=1.27
R0 B.n190 B.n57 585
R1 B.n189 B.n188 585
R2 B.n187 B.n58 585
R3 B.n186 B.n185 585
R4 B.n184 B.n59 585
R5 B.n183 B.n182 585
R6 B.n181 B.n60 585
R7 B.n180 B.n179 585
R8 B.n178 B.n61 585
R9 B.n177 B.n176 585
R10 B.n175 B.n62 585
R11 B.n174 B.n173 585
R12 B.n172 B.n63 585
R13 B.n171 B.n170 585
R14 B.n169 B.n64 585
R15 B.n168 B.n167 585
R16 B.n166 B.n65 585
R17 B.n165 B.n164 585
R18 B.n163 B.n66 585
R19 B.n162 B.n161 585
R20 B.n157 B.n67 585
R21 B.n156 B.n155 585
R22 B.n154 B.n68 585
R23 B.n153 B.n152 585
R24 B.n151 B.n69 585
R25 B.n150 B.n149 585
R26 B.n148 B.n70 585
R27 B.n147 B.n146 585
R28 B.n145 B.n71 585
R29 B.n143 B.n142 585
R30 B.n141 B.n74 585
R31 B.n140 B.n139 585
R32 B.n138 B.n75 585
R33 B.n137 B.n136 585
R34 B.n135 B.n76 585
R35 B.n134 B.n133 585
R36 B.n132 B.n77 585
R37 B.n131 B.n130 585
R38 B.n129 B.n78 585
R39 B.n128 B.n127 585
R40 B.n126 B.n79 585
R41 B.n125 B.n124 585
R42 B.n123 B.n80 585
R43 B.n122 B.n121 585
R44 B.n120 B.n81 585
R45 B.n119 B.n118 585
R46 B.n117 B.n82 585
R47 B.n116 B.n115 585
R48 B.n192 B.n191 585
R49 B.n193 B.n56 585
R50 B.n195 B.n194 585
R51 B.n196 B.n55 585
R52 B.n198 B.n197 585
R53 B.n199 B.n54 585
R54 B.n201 B.n200 585
R55 B.n202 B.n53 585
R56 B.n204 B.n203 585
R57 B.n205 B.n52 585
R58 B.n207 B.n206 585
R59 B.n208 B.n51 585
R60 B.n210 B.n209 585
R61 B.n211 B.n50 585
R62 B.n213 B.n212 585
R63 B.n214 B.n49 585
R64 B.n216 B.n215 585
R65 B.n217 B.n48 585
R66 B.n219 B.n218 585
R67 B.n220 B.n47 585
R68 B.n222 B.n221 585
R69 B.n223 B.n46 585
R70 B.n225 B.n224 585
R71 B.n226 B.n45 585
R72 B.n228 B.n227 585
R73 B.n229 B.n44 585
R74 B.n231 B.n230 585
R75 B.n232 B.n43 585
R76 B.n234 B.n233 585
R77 B.n235 B.n42 585
R78 B.n237 B.n236 585
R79 B.n238 B.n41 585
R80 B.n240 B.n239 585
R81 B.n241 B.n40 585
R82 B.n243 B.n242 585
R83 B.n244 B.n39 585
R84 B.n318 B.n317 585
R85 B.n316 B.n11 585
R86 B.n315 B.n314 585
R87 B.n313 B.n12 585
R88 B.n312 B.n311 585
R89 B.n310 B.n13 585
R90 B.n309 B.n308 585
R91 B.n307 B.n14 585
R92 B.n306 B.n305 585
R93 B.n304 B.n15 585
R94 B.n303 B.n302 585
R95 B.n301 B.n16 585
R96 B.n300 B.n299 585
R97 B.n298 B.n17 585
R98 B.n297 B.n296 585
R99 B.n295 B.n18 585
R100 B.n294 B.n293 585
R101 B.n292 B.n19 585
R102 B.n291 B.n290 585
R103 B.n289 B.n288 585
R104 B.n287 B.n23 585
R105 B.n286 B.n285 585
R106 B.n284 B.n24 585
R107 B.n283 B.n282 585
R108 B.n281 B.n25 585
R109 B.n280 B.n279 585
R110 B.n278 B.n26 585
R111 B.n277 B.n276 585
R112 B.n275 B.n27 585
R113 B.n273 B.n272 585
R114 B.n271 B.n30 585
R115 B.n270 B.n269 585
R116 B.n268 B.n31 585
R117 B.n267 B.n266 585
R118 B.n265 B.n32 585
R119 B.n264 B.n263 585
R120 B.n262 B.n33 585
R121 B.n261 B.n260 585
R122 B.n259 B.n34 585
R123 B.n258 B.n257 585
R124 B.n256 B.n35 585
R125 B.n255 B.n254 585
R126 B.n253 B.n36 585
R127 B.n252 B.n251 585
R128 B.n250 B.n37 585
R129 B.n249 B.n248 585
R130 B.n247 B.n38 585
R131 B.n246 B.n245 585
R132 B.n319 B.n10 585
R133 B.n321 B.n320 585
R134 B.n322 B.n9 585
R135 B.n324 B.n323 585
R136 B.n325 B.n8 585
R137 B.n327 B.n326 585
R138 B.n328 B.n7 585
R139 B.n330 B.n329 585
R140 B.n331 B.n6 585
R141 B.n333 B.n332 585
R142 B.n334 B.n5 585
R143 B.n336 B.n335 585
R144 B.n337 B.n4 585
R145 B.n339 B.n338 585
R146 B.n340 B.n3 585
R147 B.n342 B.n341 585
R148 B.n343 B.n0 585
R149 B.n2 B.n1 585
R150 B.n92 B.n91 585
R151 B.n93 B.n90 585
R152 B.n95 B.n94 585
R153 B.n96 B.n89 585
R154 B.n98 B.n97 585
R155 B.n99 B.n88 585
R156 B.n101 B.n100 585
R157 B.n102 B.n87 585
R158 B.n104 B.n103 585
R159 B.n105 B.n86 585
R160 B.n107 B.n106 585
R161 B.n108 B.n85 585
R162 B.n110 B.n109 585
R163 B.n111 B.n84 585
R164 B.n113 B.n112 585
R165 B.n114 B.n83 585
R166 B.n116 B.n83 478.086
R167 B.n192 B.n57 478.086
R168 B.n246 B.n39 478.086
R169 B.n319 B.n318 478.086
R170 B.n72 B.t6 286.635
R171 B.n158 B.t9 286.635
R172 B.n28 B.t0 286.635
R173 B.n20 B.t3 286.635
R174 B.n345 B.n344 256.663
R175 B.n344 B.n343 235.042
R176 B.n344 B.n2 235.042
R177 B.n117 B.n116 163.367
R178 B.n118 B.n117 163.367
R179 B.n118 B.n81 163.367
R180 B.n122 B.n81 163.367
R181 B.n123 B.n122 163.367
R182 B.n124 B.n123 163.367
R183 B.n124 B.n79 163.367
R184 B.n128 B.n79 163.367
R185 B.n129 B.n128 163.367
R186 B.n130 B.n129 163.367
R187 B.n130 B.n77 163.367
R188 B.n134 B.n77 163.367
R189 B.n135 B.n134 163.367
R190 B.n136 B.n135 163.367
R191 B.n136 B.n75 163.367
R192 B.n140 B.n75 163.367
R193 B.n141 B.n140 163.367
R194 B.n142 B.n141 163.367
R195 B.n142 B.n71 163.367
R196 B.n147 B.n71 163.367
R197 B.n148 B.n147 163.367
R198 B.n149 B.n148 163.367
R199 B.n149 B.n69 163.367
R200 B.n153 B.n69 163.367
R201 B.n154 B.n153 163.367
R202 B.n155 B.n154 163.367
R203 B.n155 B.n67 163.367
R204 B.n162 B.n67 163.367
R205 B.n163 B.n162 163.367
R206 B.n164 B.n163 163.367
R207 B.n164 B.n65 163.367
R208 B.n168 B.n65 163.367
R209 B.n169 B.n168 163.367
R210 B.n170 B.n169 163.367
R211 B.n170 B.n63 163.367
R212 B.n174 B.n63 163.367
R213 B.n175 B.n174 163.367
R214 B.n176 B.n175 163.367
R215 B.n176 B.n61 163.367
R216 B.n180 B.n61 163.367
R217 B.n181 B.n180 163.367
R218 B.n182 B.n181 163.367
R219 B.n182 B.n59 163.367
R220 B.n186 B.n59 163.367
R221 B.n187 B.n186 163.367
R222 B.n188 B.n187 163.367
R223 B.n188 B.n57 163.367
R224 B.n242 B.n39 163.367
R225 B.n242 B.n241 163.367
R226 B.n241 B.n240 163.367
R227 B.n240 B.n41 163.367
R228 B.n236 B.n41 163.367
R229 B.n236 B.n235 163.367
R230 B.n235 B.n234 163.367
R231 B.n234 B.n43 163.367
R232 B.n230 B.n43 163.367
R233 B.n230 B.n229 163.367
R234 B.n229 B.n228 163.367
R235 B.n228 B.n45 163.367
R236 B.n224 B.n45 163.367
R237 B.n224 B.n223 163.367
R238 B.n223 B.n222 163.367
R239 B.n222 B.n47 163.367
R240 B.n218 B.n47 163.367
R241 B.n218 B.n217 163.367
R242 B.n217 B.n216 163.367
R243 B.n216 B.n49 163.367
R244 B.n212 B.n49 163.367
R245 B.n212 B.n211 163.367
R246 B.n211 B.n210 163.367
R247 B.n210 B.n51 163.367
R248 B.n206 B.n51 163.367
R249 B.n206 B.n205 163.367
R250 B.n205 B.n204 163.367
R251 B.n204 B.n53 163.367
R252 B.n200 B.n53 163.367
R253 B.n200 B.n199 163.367
R254 B.n199 B.n198 163.367
R255 B.n198 B.n55 163.367
R256 B.n194 B.n55 163.367
R257 B.n194 B.n193 163.367
R258 B.n193 B.n192 163.367
R259 B.n318 B.n11 163.367
R260 B.n314 B.n11 163.367
R261 B.n314 B.n313 163.367
R262 B.n313 B.n312 163.367
R263 B.n312 B.n13 163.367
R264 B.n308 B.n13 163.367
R265 B.n308 B.n307 163.367
R266 B.n307 B.n306 163.367
R267 B.n306 B.n15 163.367
R268 B.n302 B.n15 163.367
R269 B.n302 B.n301 163.367
R270 B.n301 B.n300 163.367
R271 B.n300 B.n17 163.367
R272 B.n296 B.n17 163.367
R273 B.n296 B.n295 163.367
R274 B.n295 B.n294 163.367
R275 B.n294 B.n19 163.367
R276 B.n290 B.n19 163.367
R277 B.n290 B.n289 163.367
R278 B.n289 B.n23 163.367
R279 B.n285 B.n23 163.367
R280 B.n285 B.n284 163.367
R281 B.n284 B.n283 163.367
R282 B.n283 B.n25 163.367
R283 B.n279 B.n25 163.367
R284 B.n279 B.n278 163.367
R285 B.n278 B.n277 163.367
R286 B.n277 B.n27 163.367
R287 B.n272 B.n27 163.367
R288 B.n272 B.n271 163.367
R289 B.n271 B.n270 163.367
R290 B.n270 B.n31 163.367
R291 B.n266 B.n31 163.367
R292 B.n266 B.n265 163.367
R293 B.n265 B.n264 163.367
R294 B.n264 B.n33 163.367
R295 B.n260 B.n33 163.367
R296 B.n260 B.n259 163.367
R297 B.n259 B.n258 163.367
R298 B.n258 B.n35 163.367
R299 B.n254 B.n35 163.367
R300 B.n254 B.n253 163.367
R301 B.n253 B.n252 163.367
R302 B.n252 B.n37 163.367
R303 B.n248 B.n37 163.367
R304 B.n248 B.n247 163.367
R305 B.n247 B.n246 163.367
R306 B.n320 B.n319 163.367
R307 B.n320 B.n9 163.367
R308 B.n324 B.n9 163.367
R309 B.n325 B.n324 163.367
R310 B.n326 B.n325 163.367
R311 B.n326 B.n7 163.367
R312 B.n330 B.n7 163.367
R313 B.n331 B.n330 163.367
R314 B.n332 B.n331 163.367
R315 B.n332 B.n5 163.367
R316 B.n336 B.n5 163.367
R317 B.n337 B.n336 163.367
R318 B.n338 B.n337 163.367
R319 B.n338 B.n3 163.367
R320 B.n342 B.n3 163.367
R321 B.n343 B.n342 163.367
R322 B.n92 B.n2 163.367
R323 B.n93 B.n92 163.367
R324 B.n94 B.n93 163.367
R325 B.n94 B.n89 163.367
R326 B.n98 B.n89 163.367
R327 B.n99 B.n98 163.367
R328 B.n100 B.n99 163.367
R329 B.n100 B.n87 163.367
R330 B.n104 B.n87 163.367
R331 B.n105 B.n104 163.367
R332 B.n106 B.n105 163.367
R333 B.n106 B.n85 163.367
R334 B.n110 B.n85 163.367
R335 B.n111 B.n110 163.367
R336 B.n112 B.n111 163.367
R337 B.n112 B.n83 163.367
R338 B.n158 B.t10 154.51
R339 B.n28 B.t2 154.51
R340 B.n72 B.t7 154.506
R341 B.n20 B.t5 154.506
R342 B.n159 B.t11 123.48
R343 B.n29 B.t1 123.48
R344 B.n73 B.t8 123.475
R345 B.n21 B.t4 123.475
R346 B.n144 B.n73 59.5399
R347 B.n160 B.n159 59.5399
R348 B.n274 B.n29 59.5399
R349 B.n22 B.n21 59.5399
R350 B.n317 B.n10 31.0639
R351 B.n245 B.n244 31.0639
R352 B.n191 B.n190 31.0639
R353 B.n115 B.n114 31.0639
R354 B.n73 B.n72 31.0308
R355 B.n159 B.n158 31.0308
R356 B.n29 B.n28 31.0308
R357 B.n21 B.n20 31.0308
R358 B B.n345 18.0485
R359 B.n321 B.n10 10.6151
R360 B.n322 B.n321 10.6151
R361 B.n323 B.n322 10.6151
R362 B.n323 B.n8 10.6151
R363 B.n327 B.n8 10.6151
R364 B.n328 B.n327 10.6151
R365 B.n329 B.n328 10.6151
R366 B.n329 B.n6 10.6151
R367 B.n333 B.n6 10.6151
R368 B.n334 B.n333 10.6151
R369 B.n335 B.n334 10.6151
R370 B.n335 B.n4 10.6151
R371 B.n339 B.n4 10.6151
R372 B.n340 B.n339 10.6151
R373 B.n341 B.n340 10.6151
R374 B.n341 B.n0 10.6151
R375 B.n317 B.n316 10.6151
R376 B.n316 B.n315 10.6151
R377 B.n315 B.n12 10.6151
R378 B.n311 B.n12 10.6151
R379 B.n311 B.n310 10.6151
R380 B.n310 B.n309 10.6151
R381 B.n309 B.n14 10.6151
R382 B.n305 B.n14 10.6151
R383 B.n305 B.n304 10.6151
R384 B.n304 B.n303 10.6151
R385 B.n303 B.n16 10.6151
R386 B.n299 B.n16 10.6151
R387 B.n299 B.n298 10.6151
R388 B.n298 B.n297 10.6151
R389 B.n297 B.n18 10.6151
R390 B.n293 B.n18 10.6151
R391 B.n293 B.n292 10.6151
R392 B.n292 B.n291 10.6151
R393 B.n288 B.n287 10.6151
R394 B.n287 B.n286 10.6151
R395 B.n286 B.n24 10.6151
R396 B.n282 B.n24 10.6151
R397 B.n282 B.n281 10.6151
R398 B.n281 B.n280 10.6151
R399 B.n280 B.n26 10.6151
R400 B.n276 B.n26 10.6151
R401 B.n276 B.n275 10.6151
R402 B.n273 B.n30 10.6151
R403 B.n269 B.n30 10.6151
R404 B.n269 B.n268 10.6151
R405 B.n268 B.n267 10.6151
R406 B.n267 B.n32 10.6151
R407 B.n263 B.n32 10.6151
R408 B.n263 B.n262 10.6151
R409 B.n262 B.n261 10.6151
R410 B.n261 B.n34 10.6151
R411 B.n257 B.n34 10.6151
R412 B.n257 B.n256 10.6151
R413 B.n256 B.n255 10.6151
R414 B.n255 B.n36 10.6151
R415 B.n251 B.n36 10.6151
R416 B.n251 B.n250 10.6151
R417 B.n250 B.n249 10.6151
R418 B.n249 B.n38 10.6151
R419 B.n245 B.n38 10.6151
R420 B.n244 B.n243 10.6151
R421 B.n243 B.n40 10.6151
R422 B.n239 B.n40 10.6151
R423 B.n239 B.n238 10.6151
R424 B.n238 B.n237 10.6151
R425 B.n237 B.n42 10.6151
R426 B.n233 B.n42 10.6151
R427 B.n233 B.n232 10.6151
R428 B.n232 B.n231 10.6151
R429 B.n231 B.n44 10.6151
R430 B.n227 B.n44 10.6151
R431 B.n227 B.n226 10.6151
R432 B.n226 B.n225 10.6151
R433 B.n225 B.n46 10.6151
R434 B.n221 B.n46 10.6151
R435 B.n221 B.n220 10.6151
R436 B.n220 B.n219 10.6151
R437 B.n219 B.n48 10.6151
R438 B.n215 B.n48 10.6151
R439 B.n215 B.n214 10.6151
R440 B.n214 B.n213 10.6151
R441 B.n213 B.n50 10.6151
R442 B.n209 B.n50 10.6151
R443 B.n209 B.n208 10.6151
R444 B.n208 B.n207 10.6151
R445 B.n207 B.n52 10.6151
R446 B.n203 B.n52 10.6151
R447 B.n203 B.n202 10.6151
R448 B.n202 B.n201 10.6151
R449 B.n201 B.n54 10.6151
R450 B.n197 B.n54 10.6151
R451 B.n197 B.n196 10.6151
R452 B.n196 B.n195 10.6151
R453 B.n195 B.n56 10.6151
R454 B.n191 B.n56 10.6151
R455 B.n91 B.n1 10.6151
R456 B.n91 B.n90 10.6151
R457 B.n95 B.n90 10.6151
R458 B.n96 B.n95 10.6151
R459 B.n97 B.n96 10.6151
R460 B.n97 B.n88 10.6151
R461 B.n101 B.n88 10.6151
R462 B.n102 B.n101 10.6151
R463 B.n103 B.n102 10.6151
R464 B.n103 B.n86 10.6151
R465 B.n107 B.n86 10.6151
R466 B.n108 B.n107 10.6151
R467 B.n109 B.n108 10.6151
R468 B.n109 B.n84 10.6151
R469 B.n113 B.n84 10.6151
R470 B.n114 B.n113 10.6151
R471 B.n115 B.n82 10.6151
R472 B.n119 B.n82 10.6151
R473 B.n120 B.n119 10.6151
R474 B.n121 B.n120 10.6151
R475 B.n121 B.n80 10.6151
R476 B.n125 B.n80 10.6151
R477 B.n126 B.n125 10.6151
R478 B.n127 B.n126 10.6151
R479 B.n127 B.n78 10.6151
R480 B.n131 B.n78 10.6151
R481 B.n132 B.n131 10.6151
R482 B.n133 B.n132 10.6151
R483 B.n133 B.n76 10.6151
R484 B.n137 B.n76 10.6151
R485 B.n138 B.n137 10.6151
R486 B.n139 B.n138 10.6151
R487 B.n139 B.n74 10.6151
R488 B.n143 B.n74 10.6151
R489 B.n146 B.n145 10.6151
R490 B.n146 B.n70 10.6151
R491 B.n150 B.n70 10.6151
R492 B.n151 B.n150 10.6151
R493 B.n152 B.n151 10.6151
R494 B.n152 B.n68 10.6151
R495 B.n156 B.n68 10.6151
R496 B.n157 B.n156 10.6151
R497 B.n161 B.n157 10.6151
R498 B.n165 B.n66 10.6151
R499 B.n166 B.n165 10.6151
R500 B.n167 B.n166 10.6151
R501 B.n167 B.n64 10.6151
R502 B.n171 B.n64 10.6151
R503 B.n172 B.n171 10.6151
R504 B.n173 B.n172 10.6151
R505 B.n173 B.n62 10.6151
R506 B.n177 B.n62 10.6151
R507 B.n178 B.n177 10.6151
R508 B.n179 B.n178 10.6151
R509 B.n179 B.n60 10.6151
R510 B.n183 B.n60 10.6151
R511 B.n184 B.n183 10.6151
R512 B.n185 B.n184 10.6151
R513 B.n185 B.n58 10.6151
R514 B.n189 B.n58 10.6151
R515 B.n190 B.n189 10.6151
R516 B.n291 B.n22 9.36635
R517 B.n274 B.n273 9.36635
R518 B.n144 B.n143 9.36635
R519 B.n160 B.n66 9.36635
R520 B.n345 B.n0 8.11757
R521 B.n345 B.n1 8.11757
R522 B.n288 B.n22 1.24928
R523 B.n275 B.n274 1.24928
R524 B.n145 B.n144 1.24928
R525 B.n161 B.n160 1.24928
R526 VP.n0 VP.t0 229.212
R527 VP.n0 VP.t1 193.893
R528 VP VP.n0 0.146778
R529 VTAIL.n1 VTAIL.t0 101.736
R530 VTAIL.n3 VTAIL.t1 101.736
R531 VTAIL.n0 VTAIL.t3 101.736
R532 VTAIL.n2 VTAIL.t2 101.736
R533 VTAIL.n1 VTAIL.n0 18.8583
R534 VTAIL.n3 VTAIL.n2 17.4789
R535 VTAIL.n2 VTAIL.n1 1.15998
R536 VTAIL VTAIL.n0 0.873345
R537 VTAIL VTAIL.n3 0.287138
R538 VDD1 VDD1.t0 149.435
R539 VDD1 VDD1.t1 118.817
R540 VN VN.t0 229.498
R541 VN VN.t1 194.038
R542 VDD2.n0 VDD2.t0 148.565
R543 VDD2.n0 VDD2.t1 118.415
R544 VDD2 VDD2.n0 0.403517
C0 VDD2 VP 0.280828f
C1 B VTAIL 1.50819f
C2 B VN 0.730775f
C3 w_n1610_n1834# VTAIL 1.61844f
C4 VTAIL VDD1 2.76492f
C5 w_n1610_n1834# VN 1.95734f
C6 VN VDD1 0.151575f
C7 VDD2 VTAIL 2.80756f
C8 VDD2 VN 1.02095f
C9 VP VTAIL 1.00271f
C10 VP VN 3.41765f
C11 VN VTAIL 0.988477f
C12 B w_n1610_n1834# 5.22268f
C13 B VDD1 0.933485f
C14 B VDD2 0.952231f
C15 w_n1610_n1834# VDD1 1.07941f
C16 B VP 1.05775f
C17 w_n1610_n1834# VDD2 1.08941f
C18 VDD2 VDD1 0.519249f
C19 w_n1610_n1834# VP 2.15911f
C20 VP VDD1 1.14841f
C21 VDD2 VSUBS 0.509813f
C22 VDD1 VSUBS 2.411783f
C23 VTAIL VSUBS 0.396841f
C24 VN VSUBS 3.56601f
C25 VP VSUBS 0.90563f
C26 B VSUBS 2.160079f
C27 w_n1610_n1834# VSUBS 37.1137f
C28 VDD2.t0 VSUBS 0.595697f
C29 VDD2.t1 VSUBS 0.433612f
C30 VDD2.n0 VSUBS 1.71615f
C31 VN.t1 VSUBS 0.585922f
C32 VN.t0 VSUBS 0.755695f
C33 VDD1.t1 VSUBS 0.425912f
C34 VDD1.t0 VSUBS 0.595806f
C35 VTAIL.t3 VSUBS 0.452922f
C36 VTAIL.n0 VSUBS 0.970065f
C37 VTAIL.t0 VSUBS 0.452924f
C38 VTAIL.n1 VSUBS 0.986413f
C39 VTAIL.t2 VSUBS 0.452922f
C40 VTAIL.n2 VSUBS 0.907741f
C41 VTAIL.t1 VSUBS 0.452922f
C42 VTAIL.n3 VSUBS 0.857956f
C43 VP.t0 VSUBS 1.25395f
C44 VP.t1 VSUBS 0.97698f
C45 VP.n0 VSUBS 3.32411f
C46 B.n0 VSUBS 0.006252f
C47 B.n1 VSUBS 0.006252f
C48 B.n2 VSUBS 0.009247f
C49 B.n3 VSUBS 0.007086f
C50 B.n4 VSUBS 0.007086f
C51 B.n5 VSUBS 0.007086f
C52 B.n6 VSUBS 0.007086f
C53 B.n7 VSUBS 0.007086f
C54 B.n8 VSUBS 0.007086f
C55 B.n9 VSUBS 0.007086f
C56 B.n10 VSUBS 0.0155f
C57 B.n11 VSUBS 0.007086f
C58 B.n12 VSUBS 0.007086f
C59 B.n13 VSUBS 0.007086f
C60 B.n14 VSUBS 0.007086f
C61 B.n15 VSUBS 0.007086f
C62 B.n16 VSUBS 0.007086f
C63 B.n17 VSUBS 0.007086f
C64 B.n18 VSUBS 0.007086f
C65 B.n19 VSUBS 0.007086f
C66 B.t4 VSUBS 0.117573f
C67 B.t5 VSUBS 0.128533f
C68 B.t3 VSUBS 0.257639f
C69 B.n20 VSUBS 0.084458f
C70 B.n21 VSUBS 0.064679f
C71 B.n22 VSUBS 0.016417f
C72 B.n23 VSUBS 0.007086f
C73 B.n24 VSUBS 0.007086f
C74 B.n25 VSUBS 0.007086f
C75 B.n26 VSUBS 0.007086f
C76 B.n27 VSUBS 0.007086f
C77 B.t1 VSUBS 0.117573f
C78 B.t2 VSUBS 0.128532f
C79 B.t0 VSUBS 0.257639f
C80 B.n28 VSUBS 0.084458f
C81 B.n29 VSUBS 0.064679f
C82 B.n30 VSUBS 0.007086f
C83 B.n31 VSUBS 0.007086f
C84 B.n32 VSUBS 0.007086f
C85 B.n33 VSUBS 0.007086f
C86 B.n34 VSUBS 0.007086f
C87 B.n35 VSUBS 0.007086f
C88 B.n36 VSUBS 0.007086f
C89 B.n37 VSUBS 0.007086f
C90 B.n38 VSUBS 0.007086f
C91 B.n39 VSUBS 0.0155f
C92 B.n40 VSUBS 0.007086f
C93 B.n41 VSUBS 0.007086f
C94 B.n42 VSUBS 0.007086f
C95 B.n43 VSUBS 0.007086f
C96 B.n44 VSUBS 0.007086f
C97 B.n45 VSUBS 0.007086f
C98 B.n46 VSUBS 0.007086f
C99 B.n47 VSUBS 0.007086f
C100 B.n48 VSUBS 0.007086f
C101 B.n49 VSUBS 0.007086f
C102 B.n50 VSUBS 0.007086f
C103 B.n51 VSUBS 0.007086f
C104 B.n52 VSUBS 0.007086f
C105 B.n53 VSUBS 0.007086f
C106 B.n54 VSUBS 0.007086f
C107 B.n55 VSUBS 0.007086f
C108 B.n56 VSUBS 0.007086f
C109 B.n57 VSUBS 0.016595f
C110 B.n58 VSUBS 0.007086f
C111 B.n59 VSUBS 0.007086f
C112 B.n60 VSUBS 0.007086f
C113 B.n61 VSUBS 0.007086f
C114 B.n62 VSUBS 0.007086f
C115 B.n63 VSUBS 0.007086f
C116 B.n64 VSUBS 0.007086f
C117 B.n65 VSUBS 0.007086f
C118 B.n66 VSUBS 0.006669f
C119 B.n67 VSUBS 0.007086f
C120 B.n68 VSUBS 0.007086f
C121 B.n69 VSUBS 0.007086f
C122 B.n70 VSUBS 0.007086f
C123 B.n71 VSUBS 0.007086f
C124 B.t8 VSUBS 0.117573f
C125 B.t7 VSUBS 0.128533f
C126 B.t6 VSUBS 0.257639f
C127 B.n72 VSUBS 0.084458f
C128 B.n73 VSUBS 0.064679f
C129 B.n74 VSUBS 0.007086f
C130 B.n75 VSUBS 0.007086f
C131 B.n76 VSUBS 0.007086f
C132 B.n77 VSUBS 0.007086f
C133 B.n78 VSUBS 0.007086f
C134 B.n79 VSUBS 0.007086f
C135 B.n80 VSUBS 0.007086f
C136 B.n81 VSUBS 0.007086f
C137 B.n82 VSUBS 0.007086f
C138 B.n83 VSUBS 0.0155f
C139 B.n84 VSUBS 0.007086f
C140 B.n85 VSUBS 0.007086f
C141 B.n86 VSUBS 0.007086f
C142 B.n87 VSUBS 0.007086f
C143 B.n88 VSUBS 0.007086f
C144 B.n89 VSUBS 0.007086f
C145 B.n90 VSUBS 0.007086f
C146 B.n91 VSUBS 0.007086f
C147 B.n92 VSUBS 0.007086f
C148 B.n93 VSUBS 0.007086f
C149 B.n94 VSUBS 0.007086f
C150 B.n95 VSUBS 0.007086f
C151 B.n96 VSUBS 0.007086f
C152 B.n97 VSUBS 0.007086f
C153 B.n98 VSUBS 0.007086f
C154 B.n99 VSUBS 0.007086f
C155 B.n100 VSUBS 0.007086f
C156 B.n101 VSUBS 0.007086f
C157 B.n102 VSUBS 0.007086f
C158 B.n103 VSUBS 0.007086f
C159 B.n104 VSUBS 0.007086f
C160 B.n105 VSUBS 0.007086f
C161 B.n106 VSUBS 0.007086f
C162 B.n107 VSUBS 0.007086f
C163 B.n108 VSUBS 0.007086f
C164 B.n109 VSUBS 0.007086f
C165 B.n110 VSUBS 0.007086f
C166 B.n111 VSUBS 0.007086f
C167 B.n112 VSUBS 0.007086f
C168 B.n113 VSUBS 0.007086f
C169 B.n114 VSUBS 0.0155f
C170 B.n115 VSUBS 0.016595f
C171 B.n116 VSUBS 0.016595f
C172 B.n117 VSUBS 0.007086f
C173 B.n118 VSUBS 0.007086f
C174 B.n119 VSUBS 0.007086f
C175 B.n120 VSUBS 0.007086f
C176 B.n121 VSUBS 0.007086f
C177 B.n122 VSUBS 0.007086f
C178 B.n123 VSUBS 0.007086f
C179 B.n124 VSUBS 0.007086f
C180 B.n125 VSUBS 0.007086f
C181 B.n126 VSUBS 0.007086f
C182 B.n127 VSUBS 0.007086f
C183 B.n128 VSUBS 0.007086f
C184 B.n129 VSUBS 0.007086f
C185 B.n130 VSUBS 0.007086f
C186 B.n131 VSUBS 0.007086f
C187 B.n132 VSUBS 0.007086f
C188 B.n133 VSUBS 0.007086f
C189 B.n134 VSUBS 0.007086f
C190 B.n135 VSUBS 0.007086f
C191 B.n136 VSUBS 0.007086f
C192 B.n137 VSUBS 0.007086f
C193 B.n138 VSUBS 0.007086f
C194 B.n139 VSUBS 0.007086f
C195 B.n140 VSUBS 0.007086f
C196 B.n141 VSUBS 0.007086f
C197 B.n142 VSUBS 0.007086f
C198 B.n143 VSUBS 0.006669f
C199 B.n144 VSUBS 0.016417f
C200 B.n145 VSUBS 0.00396f
C201 B.n146 VSUBS 0.007086f
C202 B.n147 VSUBS 0.007086f
C203 B.n148 VSUBS 0.007086f
C204 B.n149 VSUBS 0.007086f
C205 B.n150 VSUBS 0.007086f
C206 B.n151 VSUBS 0.007086f
C207 B.n152 VSUBS 0.007086f
C208 B.n153 VSUBS 0.007086f
C209 B.n154 VSUBS 0.007086f
C210 B.n155 VSUBS 0.007086f
C211 B.n156 VSUBS 0.007086f
C212 B.n157 VSUBS 0.007086f
C213 B.t11 VSUBS 0.117573f
C214 B.t10 VSUBS 0.128532f
C215 B.t9 VSUBS 0.257639f
C216 B.n158 VSUBS 0.084458f
C217 B.n159 VSUBS 0.064679f
C218 B.n160 VSUBS 0.016417f
C219 B.n161 VSUBS 0.00396f
C220 B.n162 VSUBS 0.007086f
C221 B.n163 VSUBS 0.007086f
C222 B.n164 VSUBS 0.007086f
C223 B.n165 VSUBS 0.007086f
C224 B.n166 VSUBS 0.007086f
C225 B.n167 VSUBS 0.007086f
C226 B.n168 VSUBS 0.007086f
C227 B.n169 VSUBS 0.007086f
C228 B.n170 VSUBS 0.007086f
C229 B.n171 VSUBS 0.007086f
C230 B.n172 VSUBS 0.007086f
C231 B.n173 VSUBS 0.007086f
C232 B.n174 VSUBS 0.007086f
C233 B.n175 VSUBS 0.007086f
C234 B.n176 VSUBS 0.007086f
C235 B.n177 VSUBS 0.007086f
C236 B.n178 VSUBS 0.007086f
C237 B.n179 VSUBS 0.007086f
C238 B.n180 VSUBS 0.007086f
C239 B.n181 VSUBS 0.007086f
C240 B.n182 VSUBS 0.007086f
C241 B.n183 VSUBS 0.007086f
C242 B.n184 VSUBS 0.007086f
C243 B.n185 VSUBS 0.007086f
C244 B.n186 VSUBS 0.007086f
C245 B.n187 VSUBS 0.007086f
C246 B.n188 VSUBS 0.007086f
C247 B.n189 VSUBS 0.007086f
C248 B.n190 VSUBS 0.015715f
C249 B.n191 VSUBS 0.01638f
C250 B.n192 VSUBS 0.0155f
C251 B.n193 VSUBS 0.007086f
C252 B.n194 VSUBS 0.007086f
C253 B.n195 VSUBS 0.007086f
C254 B.n196 VSUBS 0.007086f
C255 B.n197 VSUBS 0.007086f
C256 B.n198 VSUBS 0.007086f
C257 B.n199 VSUBS 0.007086f
C258 B.n200 VSUBS 0.007086f
C259 B.n201 VSUBS 0.007086f
C260 B.n202 VSUBS 0.007086f
C261 B.n203 VSUBS 0.007086f
C262 B.n204 VSUBS 0.007086f
C263 B.n205 VSUBS 0.007086f
C264 B.n206 VSUBS 0.007086f
C265 B.n207 VSUBS 0.007086f
C266 B.n208 VSUBS 0.007086f
C267 B.n209 VSUBS 0.007086f
C268 B.n210 VSUBS 0.007086f
C269 B.n211 VSUBS 0.007086f
C270 B.n212 VSUBS 0.007086f
C271 B.n213 VSUBS 0.007086f
C272 B.n214 VSUBS 0.007086f
C273 B.n215 VSUBS 0.007086f
C274 B.n216 VSUBS 0.007086f
C275 B.n217 VSUBS 0.007086f
C276 B.n218 VSUBS 0.007086f
C277 B.n219 VSUBS 0.007086f
C278 B.n220 VSUBS 0.007086f
C279 B.n221 VSUBS 0.007086f
C280 B.n222 VSUBS 0.007086f
C281 B.n223 VSUBS 0.007086f
C282 B.n224 VSUBS 0.007086f
C283 B.n225 VSUBS 0.007086f
C284 B.n226 VSUBS 0.007086f
C285 B.n227 VSUBS 0.007086f
C286 B.n228 VSUBS 0.007086f
C287 B.n229 VSUBS 0.007086f
C288 B.n230 VSUBS 0.007086f
C289 B.n231 VSUBS 0.007086f
C290 B.n232 VSUBS 0.007086f
C291 B.n233 VSUBS 0.007086f
C292 B.n234 VSUBS 0.007086f
C293 B.n235 VSUBS 0.007086f
C294 B.n236 VSUBS 0.007086f
C295 B.n237 VSUBS 0.007086f
C296 B.n238 VSUBS 0.007086f
C297 B.n239 VSUBS 0.007086f
C298 B.n240 VSUBS 0.007086f
C299 B.n241 VSUBS 0.007086f
C300 B.n242 VSUBS 0.007086f
C301 B.n243 VSUBS 0.007086f
C302 B.n244 VSUBS 0.0155f
C303 B.n245 VSUBS 0.016595f
C304 B.n246 VSUBS 0.016595f
C305 B.n247 VSUBS 0.007086f
C306 B.n248 VSUBS 0.007086f
C307 B.n249 VSUBS 0.007086f
C308 B.n250 VSUBS 0.007086f
C309 B.n251 VSUBS 0.007086f
C310 B.n252 VSUBS 0.007086f
C311 B.n253 VSUBS 0.007086f
C312 B.n254 VSUBS 0.007086f
C313 B.n255 VSUBS 0.007086f
C314 B.n256 VSUBS 0.007086f
C315 B.n257 VSUBS 0.007086f
C316 B.n258 VSUBS 0.007086f
C317 B.n259 VSUBS 0.007086f
C318 B.n260 VSUBS 0.007086f
C319 B.n261 VSUBS 0.007086f
C320 B.n262 VSUBS 0.007086f
C321 B.n263 VSUBS 0.007086f
C322 B.n264 VSUBS 0.007086f
C323 B.n265 VSUBS 0.007086f
C324 B.n266 VSUBS 0.007086f
C325 B.n267 VSUBS 0.007086f
C326 B.n268 VSUBS 0.007086f
C327 B.n269 VSUBS 0.007086f
C328 B.n270 VSUBS 0.007086f
C329 B.n271 VSUBS 0.007086f
C330 B.n272 VSUBS 0.007086f
C331 B.n273 VSUBS 0.006669f
C332 B.n274 VSUBS 0.016417f
C333 B.n275 VSUBS 0.00396f
C334 B.n276 VSUBS 0.007086f
C335 B.n277 VSUBS 0.007086f
C336 B.n278 VSUBS 0.007086f
C337 B.n279 VSUBS 0.007086f
C338 B.n280 VSUBS 0.007086f
C339 B.n281 VSUBS 0.007086f
C340 B.n282 VSUBS 0.007086f
C341 B.n283 VSUBS 0.007086f
C342 B.n284 VSUBS 0.007086f
C343 B.n285 VSUBS 0.007086f
C344 B.n286 VSUBS 0.007086f
C345 B.n287 VSUBS 0.007086f
C346 B.n288 VSUBS 0.00396f
C347 B.n289 VSUBS 0.007086f
C348 B.n290 VSUBS 0.007086f
C349 B.n291 VSUBS 0.006669f
C350 B.n292 VSUBS 0.007086f
C351 B.n293 VSUBS 0.007086f
C352 B.n294 VSUBS 0.007086f
C353 B.n295 VSUBS 0.007086f
C354 B.n296 VSUBS 0.007086f
C355 B.n297 VSUBS 0.007086f
C356 B.n298 VSUBS 0.007086f
C357 B.n299 VSUBS 0.007086f
C358 B.n300 VSUBS 0.007086f
C359 B.n301 VSUBS 0.007086f
C360 B.n302 VSUBS 0.007086f
C361 B.n303 VSUBS 0.007086f
C362 B.n304 VSUBS 0.007086f
C363 B.n305 VSUBS 0.007086f
C364 B.n306 VSUBS 0.007086f
C365 B.n307 VSUBS 0.007086f
C366 B.n308 VSUBS 0.007086f
C367 B.n309 VSUBS 0.007086f
C368 B.n310 VSUBS 0.007086f
C369 B.n311 VSUBS 0.007086f
C370 B.n312 VSUBS 0.007086f
C371 B.n313 VSUBS 0.007086f
C372 B.n314 VSUBS 0.007086f
C373 B.n315 VSUBS 0.007086f
C374 B.n316 VSUBS 0.007086f
C375 B.n317 VSUBS 0.016595f
C376 B.n318 VSUBS 0.016595f
C377 B.n319 VSUBS 0.0155f
C378 B.n320 VSUBS 0.007086f
C379 B.n321 VSUBS 0.007086f
C380 B.n322 VSUBS 0.007086f
C381 B.n323 VSUBS 0.007086f
C382 B.n324 VSUBS 0.007086f
C383 B.n325 VSUBS 0.007086f
C384 B.n326 VSUBS 0.007086f
C385 B.n327 VSUBS 0.007086f
C386 B.n328 VSUBS 0.007086f
C387 B.n329 VSUBS 0.007086f
C388 B.n330 VSUBS 0.007086f
C389 B.n331 VSUBS 0.007086f
C390 B.n332 VSUBS 0.007086f
C391 B.n333 VSUBS 0.007086f
C392 B.n334 VSUBS 0.007086f
C393 B.n335 VSUBS 0.007086f
C394 B.n336 VSUBS 0.007086f
C395 B.n337 VSUBS 0.007086f
C396 B.n338 VSUBS 0.007086f
C397 B.n339 VSUBS 0.007086f
C398 B.n340 VSUBS 0.007086f
C399 B.n341 VSUBS 0.007086f
C400 B.n342 VSUBS 0.007086f
C401 B.n343 VSUBS 0.009247f
C402 B.n344 VSUBS 0.00985f
C403 B.n345 VSUBS 0.019588f
.ends

