* NGSPICE file created from diff_pair_sample_1792.ext - technology: sky130A

.subckt diff_pair_sample_1792 VTAIL VN VP B VDD2 VDD1
X0 B.t21 B.t19 B.t20 B.t9 sky130_fd_pr__nfet_01v8 ad=6.1269 pd=32.2 as=0 ps=0 w=15.71 l=3.98
X1 VDD2.t7 VN.t0 VTAIL.t9 B.t7 sky130_fd_pr__nfet_01v8 ad=2.59215 pd=16.04 as=2.59215 ps=16.04 w=15.71 l=3.98
X2 VTAIL.t3 VP.t0 VDD1.t7 B.t4 sky130_fd_pr__nfet_01v8 ad=2.59215 pd=16.04 as=2.59215 ps=16.04 w=15.71 l=3.98
X3 B.t18 B.t16 B.t17 B.t13 sky130_fd_pr__nfet_01v8 ad=6.1269 pd=32.2 as=0 ps=0 w=15.71 l=3.98
X4 VTAIL.t12 VN.t1 VDD2.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=6.1269 pd=32.2 as=2.59215 ps=16.04 w=15.71 l=3.98
X5 VTAIL.t7 VP.t1 VDD1.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=2.59215 pd=16.04 as=2.59215 ps=16.04 w=15.71 l=3.98
X6 VTAIL.t13 VN.t2 VDD2.t5 B.t4 sky130_fd_pr__nfet_01v8 ad=2.59215 pd=16.04 as=2.59215 ps=16.04 w=15.71 l=3.98
X7 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=6.1269 pd=32.2 as=0 ps=0 w=15.71 l=3.98
X8 VTAIL.t11 VN.t3 VDD2.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=2.59215 pd=16.04 as=2.59215 ps=16.04 w=15.71 l=3.98
X9 VTAIL.t5 VP.t2 VDD1.t5 B.t6 sky130_fd_pr__nfet_01v8 ad=6.1269 pd=32.2 as=2.59215 ps=16.04 w=15.71 l=3.98
X10 VDD1.t4 VP.t3 VTAIL.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=2.59215 pd=16.04 as=2.59215 ps=16.04 w=15.71 l=3.98
X11 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=6.1269 pd=32.2 as=0 ps=0 w=15.71 l=3.98
X12 VDD1.t3 VP.t4 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.59215 pd=16.04 as=6.1269 ps=32.2 w=15.71 l=3.98
X13 VDD2.t3 VN.t4 VTAIL.t10 B.t2 sky130_fd_pr__nfet_01v8 ad=2.59215 pd=16.04 as=6.1269 ps=32.2 w=15.71 l=3.98
X14 VDD1.t2 VP.t5 VTAIL.t6 B.t7 sky130_fd_pr__nfet_01v8 ad=2.59215 pd=16.04 as=2.59215 ps=16.04 w=15.71 l=3.98
X15 VDD2.t2 VN.t5 VTAIL.t14 B.t0 sky130_fd_pr__nfet_01v8 ad=2.59215 pd=16.04 as=6.1269 ps=32.2 w=15.71 l=3.98
X16 VDD2.t1 VN.t6 VTAIL.t8 B.t3 sky130_fd_pr__nfet_01v8 ad=2.59215 pd=16.04 as=2.59215 ps=16.04 w=15.71 l=3.98
X17 VDD1.t1 VP.t6 VTAIL.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=2.59215 pd=16.04 as=6.1269 ps=32.2 w=15.71 l=3.98
X18 VTAIL.t15 VN.t7 VDD2.t0 B.t6 sky130_fd_pr__nfet_01v8 ad=6.1269 pd=32.2 as=2.59215 ps=16.04 w=15.71 l=3.98
X19 VTAIL.t4 VP.t7 VDD1.t0 B.t5 sky130_fd_pr__nfet_01v8 ad=6.1269 pd=32.2 as=2.59215 ps=16.04 w=15.71 l=3.98
R0 B.n1157 B.n1156 585
R1 B.n1158 B.n1157 585
R2 B.n418 B.n188 585
R3 B.n417 B.n416 585
R4 B.n415 B.n414 585
R5 B.n413 B.n412 585
R6 B.n411 B.n410 585
R7 B.n409 B.n408 585
R8 B.n407 B.n406 585
R9 B.n405 B.n404 585
R10 B.n403 B.n402 585
R11 B.n401 B.n400 585
R12 B.n399 B.n398 585
R13 B.n397 B.n396 585
R14 B.n395 B.n394 585
R15 B.n393 B.n392 585
R16 B.n391 B.n390 585
R17 B.n389 B.n388 585
R18 B.n387 B.n386 585
R19 B.n385 B.n384 585
R20 B.n383 B.n382 585
R21 B.n381 B.n380 585
R22 B.n379 B.n378 585
R23 B.n377 B.n376 585
R24 B.n375 B.n374 585
R25 B.n373 B.n372 585
R26 B.n371 B.n370 585
R27 B.n369 B.n368 585
R28 B.n367 B.n366 585
R29 B.n365 B.n364 585
R30 B.n363 B.n362 585
R31 B.n361 B.n360 585
R32 B.n359 B.n358 585
R33 B.n357 B.n356 585
R34 B.n355 B.n354 585
R35 B.n353 B.n352 585
R36 B.n351 B.n350 585
R37 B.n349 B.n348 585
R38 B.n347 B.n346 585
R39 B.n345 B.n344 585
R40 B.n343 B.n342 585
R41 B.n341 B.n340 585
R42 B.n339 B.n338 585
R43 B.n337 B.n336 585
R44 B.n335 B.n334 585
R45 B.n333 B.n332 585
R46 B.n331 B.n330 585
R47 B.n329 B.n328 585
R48 B.n327 B.n326 585
R49 B.n325 B.n324 585
R50 B.n323 B.n322 585
R51 B.n321 B.n320 585
R52 B.n319 B.n318 585
R53 B.n317 B.n316 585
R54 B.n315 B.n314 585
R55 B.n313 B.n312 585
R56 B.n311 B.n310 585
R57 B.n309 B.n308 585
R58 B.n307 B.n306 585
R59 B.n305 B.n304 585
R60 B.n303 B.n302 585
R61 B.n301 B.n300 585
R62 B.n299 B.n298 585
R63 B.n296 B.n295 585
R64 B.n294 B.n293 585
R65 B.n292 B.n291 585
R66 B.n290 B.n289 585
R67 B.n288 B.n287 585
R68 B.n286 B.n285 585
R69 B.n284 B.n283 585
R70 B.n282 B.n281 585
R71 B.n280 B.n279 585
R72 B.n278 B.n277 585
R73 B.n276 B.n275 585
R74 B.n274 B.n273 585
R75 B.n272 B.n271 585
R76 B.n270 B.n269 585
R77 B.n268 B.n267 585
R78 B.n266 B.n265 585
R79 B.n264 B.n263 585
R80 B.n262 B.n261 585
R81 B.n260 B.n259 585
R82 B.n258 B.n257 585
R83 B.n256 B.n255 585
R84 B.n254 B.n253 585
R85 B.n252 B.n251 585
R86 B.n250 B.n249 585
R87 B.n248 B.n247 585
R88 B.n246 B.n245 585
R89 B.n244 B.n243 585
R90 B.n242 B.n241 585
R91 B.n240 B.n239 585
R92 B.n238 B.n237 585
R93 B.n236 B.n235 585
R94 B.n234 B.n233 585
R95 B.n232 B.n231 585
R96 B.n230 B.n229 585
R97 B.n228 B.n227 585
R98 B.n226 B.n225 585
R99 B.n224 B.n223 585
R100 B.n222 B.n221 585
R101 B.n220 B.n219 585
R102 B.n218 B.n217 585
R103 B.n216 B.n215 585
R104 B.n214 B.n213 585
R105 B.n212 B.n211 585
R106 B.n210 B.n209 585
R107 B.n208 B.n207 585
R108 B.n206 B.n205 585
R109 B.n204 B.n203 585
R110 B.n202 B.n201 585
R111 B.n200 B.n199 585
R112 B.n198 B.n197 585
R113 B.n196 B.n195 585
R114 B.n131 B.n130 585
R115 B.n1161 B.n1160 585
R116 B.n1155 B.n189 585
R117 B.n189 B.n128 585
R118 B.n1154 B.n127 585
R119 B.n1165 B.n127 585
R120 B.n1153 B.n126 585
R121 B.n1166 B.n126 585
R122 B.n1152 B.n125 585
R123 B.n1167 B.n125 585
R124 B.n1151 B.n1150 585
R125 B.n1150 B.n121 585
R126 B.n1149 B.n120 585
R127 B.n1173 B.n120 585
R128 B.n1148 B.n119 585
R129 B.n1174 B.n119 585
R130 B.n1147 B.n118 585
R131 B.n1175 B.n118 585
R132 B.n1146 B.n1145 585
R133 B.n1145 B.n114 585
R134 B.n1144 B.n113 585
R135 B.n1181 B.n113 585
R136 B.n1143 B.n112 585
R137 B.n1182 B.n112 585
R138 B.n1142 B.n111 585
R139 B.n1183 B.n111 585
R140 B.n1141 B.n1140 585
R141 B.n1140 B.n107 585
R142 B.n1139 B.n106 585
R143 B.n1189 B.n106 585
R144 B.n1138 B.n105 585
R145 B.n1190 B.n105 585
R146 B.n1137 B.n104 585
R147 B.n1191 B.n104 585
R148 B.n1136 B.n1135 585
R149 B.n1135 B.n100 585
R150 B.n1134 B.n99 585
R151 B.n1197 B.n99 585
R152 B.n1133 B.n98 585
R153 B.n1198 B.n98 585
R154 B.n1132 B.n97 585
R155 B.n1199 B.n97 585
R156 B.n1131 B.n1130 585
R157 B.n1130 B.n93 585
R158 B.n1129 B.n92 585
R159 B.n1205 B.n92 585
R160 B.n1128 B.n91 585
R161 B.n1206 B.n91 585
R162 B.n1127 B.n90 585
R163 B.n1207 B.n90 585
R164 B.n1126 B.n1125 585
R165 B.n1125 B.n86 585
R166 B.n1124 B.n85 585
R167 B.n1213 B.n85 585
R168 B.n1123 B.n84 585
R169 B.n1214 B.n84 585
R170 B.n1122 B.n83 585
R171 B.n1215 B.n83 585
R172 B.n1121 B.n1120 585
R173 B.n1120 B.n79 585
R174 B.n1119 B.n78 585
R175 B.n1221 B.n78 585
R176 B.n1118 B.n77 585
R177 B.n1222 B.n77 585
R178 B.n1117 B.n76 585
R179 B.n1223 B.n76 585
R180 B.n1116 B.n1115 585
R181 B.n1115 B.n72 585
R182 B.n1114 B.n71 585
R183 B.n1229 B.n71 585
R184 B.n1113 B.n70 585
R185 B.n1230 B.n70 585
R186 B.n1112 B.n69 585
R187 B.n1231 B.n69 585
R188 B.n1111 B.n1110 585
R189 B.n1110 B.n65 585
R190 B.n1109 B.n64 585
R191 B.n1237 B.n64 585
R192 B.n1108 B.n63 585
R193 B.n1238 B.n63 585
R194 B.n1107 B.n62 585
R195 B.n1239 B.n62 585
R196 B.n1106 B.n1105 585
R197 B.n1105 B.n58 585
R198 B.n1104 B.n57 585
R199 B.n1245 B.n57 585
R200 B.n1103 B.n56 585
R201 B.n1246 B.n56 585
R202 B.n1102 B.n55 585
R203 B.n1247 B.n55 585
R204 B.n1101 B.n1100 585
R205 B.n1100 B.n51 585
R206 B.n1099 B.n50 585
R207 B.n1253 B.n50 585
R208 B.n1098 B.n49 585
R209 B.n1254 B.n49 585
R210 B.n1097 B.n48 585
R211 B.n1255 B.n48 585
R212 B.n1096 B.n1095 585
R213 B.n1095 B.n44 585
R214 B.n1094 B.n43 585
R215 B.n1261 B.n43 585
R216 B.n1093 B.n42 585
R217 B.n1262 B.n42 585
R218 B.n1092 B.n41 585
R219 B.n1263 B.n41 585
R220 B.n1091 B.n1090 585
R221 B.n1090 B.n37 585
R222 B.n1089 B.n36 585
R223 B.n1269 B.n36 585
R224 B.n1088 B.n35 585
R225 B.n1270 B.n35 585
R226 B.n1087 B.n34 585
R227 B.n1271 B.n34 585
R228 B.n1086 B.n1085 585
R229 B.n1085 B.n30 585
R230 B.n1084 B.n29 585
R231 B.n1277 B.n29 585
R232 B.n1083 B.n28 585
R233 B.n1278 B.n28 585
R234 B.n1082 B.n27 585
R235 B.n1279 B.n27 585
R236 B.n1081 B.n1080 585
R237 B.n1080 B.n23 585
R238 B.n1079 B.n22 585
R239 B.n1285 B.n22 585
R240 B.n1078 B.n21 585
R241 B.n1286 B.n21 585
R242 B.n1077 B.n20 585
R243 B.n1287 B.n20 585
R244 B.n1076 B.n1075 585
R245 B.n1075 B.n16 585
R246 B.n1074 B.n15 585
R247 B.n1293 B.n15 585
R248 B.n1073 B.n14 585
R249 B.n1294 B.n14 585
R250 B.n1072 B.n13 585
R251 B.n1295 B.n13 585
R252 B.n1071 B.n1070 585
R253 B.n1070 B.n12 585
R254 B.n1069 B.n1068 585
R255 B.n1069 B.n8 585
R256 B.n1067 B.n7 585
R257 B.n1302 B.n7 585
R258 B.n1066 B.n6 585
R259 B.n1303 B.n6 585
R260 B.n1065 B.n5 585
R261 B.n1304 B.n5 585
R262 B.n1064 B.n1063 585
R263 B.n1063 B.n4 585
R264 B.n1062 B.n419 585
R265 B.n1062 B.n1061 585
R266 B.n1052 B.n420 585
R267 B.n421 B.n420 585
R268 B.n1054 B.n1053 585
R269 B.n1055 B.n1054 585
R270 B.n1051 B.n426 585
R271 B.n426 B.n425 585
R272 B.n1050 B.n1049 585
R273 B.n1049 B.n1048 585
R274 B.n428 B.n427 585
R275 B.n429 B.n428 585
R276 B.n1041 B.n1040 585
R277 B.n1042 B.n1041 585
R278 B.n1039 B.n434 585
R279 B.n434 B.n433 585
R280 B.n1038 B.n1037 585
R281 B.n1037 B.n1036 585
R282 B.n436 B.n435 585
R283 B.n437 B.n436 585
R284 B.n1029 B.n1028 585
R285 B.n1030 B.n1029 585
R286 B.n1027 B.n442 585
R287 B.n442 B.n441 585
R288 B.n1026 B.n1025 585
R289 B.n1025 B.n1024 585
R290 B.n444 B.n443 585
R291 B.n445 B.n444 585
R292 B.n1017 B.n1016 585
R293 B.n1018 B.n1017 585
R294 B.n1015 B.n450 585
R295 B.n450 B.n449 585
R296 B.n1014 B.n1013 585
R297 B.n1013 B.n1012 585
R298 B.n452 B.n451 585
R299 B.n453 B.n452 585
R300 B.n1005 B.n1004 585
R301 B.n1006 B.n1005 585
R302 B.n1003 B.n457 585
R303 B.n461 B.n457 585
R304 B.n1002 B.n1001 585
R305 B.n1001 B.n1000 585
R306 B.n459 B.n458 585
R307 B.n460 B.n459 585
R308 B.n993 B.n992 585
R309 B.n994 B.n993 585
R310 B.n991 B.n466 585
R311 B.n466 B.n465 585
R312 B.n990 B.n989 585
R313 B.n989 B.n988 585
R314 B.n468 B.n467 585
R315 B.n469 B.n468 585
R316 B.n981 B.n980 585
R317 B.n982 B.n981 585
R318 B.n979 B.n474 585
R319 B.n474 B.n473 585
R320 B.n978 B.n977 585
R321 B.n977 B.n976 585
R322 B.n476 B.n475 585
R323 B.n477 B.n476 585
R324 B.n969 B.n968 585
R325 B.n970 B.n969 585
R326 B.n967 B.n481 585
R327 B.n485 B.n481 585
R328 B.n966 B.n965 585
R329 B.n965 B.n964 585
R330 B.n483 B.n482 585
R331 B.n484 B.n483 585
R332 B.n957 B.n956 585
R333 B.n958 B.n957 585
R334 B.n955 B.n490 585
R335 B.n490 B.n489 585
R336 B.n954 B.n953 585
R337 B.n953 B.n952 585
R338 B.n492 B.n491 585
R339 B.n493 B.n492 585
R340 B.n945 B.n944 585
R341 B.n946 B.n945 585
R342 B.n943 B.n498 585
R343 B.n498 B.n497 585
R344 B.n942 B.n941 585
R345 B.n941 B.n940 585
R346 B.n500 B.n499 585
R347 B.n501 B.n500 585
R348 B.n933 B.n932 585
R349 B.n934 B.n933 585
R350 B.n931 B.n506 585
R351 B.n506 B.n505 585
R352 B.n930 B.n929 585
R353 B.n929 B.n928 585
R354 B.n508 B.n507 585
R355 B.n509 B.n508 585
R356 B.n921 B.n920 585
R357 B.n922 B.n921 585
R358 B.n919 B.n514 585
R359 B.n514 B.n513 585
R360 B.n918 B.n917 585
R361 B.n917 B.n916 585
R362 B.n516 B.n515 585
R363 B.n517 B.n516 585
R364 B.n909 B.n908 585
R365 B.n910 B.n909 585
R366 B.n907 B.n522 585
R367 B.n522 B.n521 585
R368 B.n906 B.n905 585
R369 B.n905 B.n904 585
R370 B.n524 B.n523 585
R371 B.n525 B.n524 585
R372 B.n897 B.n896 585
R373 B.n898 B.n897 585
R374 B.n895 B.n530 585
R375 B.n530 B.n529 585
R376 B.n894 B.n893 585
R377 B.n893 B.n892 585
R378 B.n532 B.n531 585
R379 B.n533 B.n532 585
R380 B.n885 B.n884 585
R381 B.n886 B.n885 585
R382 B.n883 B.n538 585
R383 B.n538 B.n537 585
R384 B.n882 B.n881 585
R385 B.n881 B.n880 585
R386 B.n540 B.n539 585
R387 B.n541 B.n540 585
R388 B.n873 B.n872 585
R389 B.n874 B.n873 585
R390 B.n871 B.n546 585
R391 B.n546 B.n545 585
R392 B.n870 B.n869 585
R393 B.n869 B.n868 585
R394 B.n548 B.n547 585
R395 B.n549 B.n548 585
R396 B.n861 B.n860 585
R397 B.n862 B.n861 585
R398 B.n859 B.n554 585
R399 B.n554 B.n553 585
R400 B.n858 B.n857 585
R401 B.n857 B.n856 585
R402 B.n556 B.n555 585
R403 B.n557 B.n556 585
R404 B.n852 B.n851 585
R405 B.n560 B.n559 585
R406 B.n848 B.n847 585
R407 B.n849 B.n848 585
R408 B.n846 B.n617 585
R409 B.n845 B.n844 585
R410 B.n843 B.n842 585
R411 B.n841 B.n840 585
R412 B.n839 B.n838 585
R413 B.n837 B.n836 585
R414 B.n835 B.n834 585
R415 B.n833 B.n832 585
R416 B.n831 B.n830 585
R417 B.n829 B.n828 585
R418 B.n827 B.n826 585
R419 B.n825 B.n824 585
R420 B.n823 B.n822 585
R421 B.n821 B.n820 585
R422 B.n819 B.n818 585
R423 B.n817 B.n816 585
R424 B.n815 B.n814 585
R425 B.n813 B.n812 585
R426 B.n811 B.n810 585
R427 B.n809 B.n808 585
R428 B.n807 B.n806 585
R429 B.n805 B.n804 585
R430 B.n803 B.n802 585
R431 B.n801 B.n800 585
R432 B.n799 B.n798 585
R433 B.n797 B.n796 585
R434 B.n795 B.n794 585
R435 B.n793 B.n792 585
R436 B.n791 B.n790 585
R437 B.n789 B.n788 585
R438 B.n787 B.n786 585
R439 B.n785 B.n784 585
R440 B.n783 B.n782 585
R441 B.n781 B.n780 585
R442 B.n779 B.n778 585
R443 B.n777 B.n776 585
R444 B.n775 B.n774 585
R445 B.n773 B.n772 585
R446 B.n771 B.n770 585
R447 B.n769 B.n768 585
R448 B.n767 B.n766 585
R449 B.n765 B.n764 585
R450 B.n763 B.n762 585
R451 B.n761 B.n760 585
R452 B.n759 B.n758 585
R453 B.n757 B.n756 585
R454 B.n755 B.n754 585
R455 B.n753 B.n752 585
R456 B.n751 B.n750 585
R457 B.n749 B.n748 585
R458 B.n747 B.n746 585
R459 B.n745 B.n744 585
R460 B.n743 B.n742 585
R461 B.n741 B.n740 585
R462 B.n739 B.n738 585
R463 B.n737 B.n736 585
R464 B.n735 B.n734 585
R465 B.n733 B.n732 585
R466 B.n731 B.n730 585
R467 B.n728 B.n727 585
R468 B.n726 B.n725 585
R469 B.n724 B.n723 585
R470 B.n722 B.n721 585
R471 B.n720 B.n719 585
R472 B.n718 B.n717 585
R473 B.n716 B.n715 585
R474 B.n714 B.n713 585
R475 B.n712 B.n711 585
R476 B.n710 B.n709 585
R477 B.n708 B.n707 585
R478 B.n706 B.n705 585
R479 B.n704 B.n703 585
R480 B.n702 B.n701 585
R481 B.n700 B.n699 585
R482 B.n698 B.n697 585
R483 B.n696 B.n695 585
R484 B.n694 B.n693 585
R485 B.n692 B.n691 585
R486 B.n690 B.n689 585
R487 B.n688 B.n687 585
R488 B.n686 B.n685 585
R489 B.n684 B.n683 585
R490 B.n682 B.n681 585
R491 B.n680 B.n679 585
R492 B.n678 B.n677 585
R493 B.n676 B.n675 585
R494 B.n674 B.n673 585
R495 B.n672 B.n671 585
R496 B.n670 B.n669 585
R497 B.n668 B.n667 585
R498 B.n666 B.n665 585
R499 B.n664 B.n663 585
R500 B.n662 B.n661 585
R501 B.n660 B.n659 585
R502 B.n658 B.n657 585
R503 B.n656 B.n655 585
R504 B.n654 B.n653 585
R505 B.n652 B.n651 585
R506 B.n650 B.n649 585
R507 B.n648 B.n647 585
R508 B.n646 B.n645 585
R509 B.n644 B.n643 585
R510 B.n642 B.n641 585
R511 B.n640 B.n639 585
R512 B.n638 B.n637 585
R513 B.n636 B.n635 585
R514 B.n634 B.n633 585
R515 B.n632 B.n631 585
R516 B.n630 B.n629 585
R517 B.n628 B.n627 585
R518 B.n626 B.n625 585
R519 B.n624 B.n623 585
R520 B.n853 B.n558 585
R521 B.n558 B.n557 585
R522 B.n855 B.n854 585
R523 B.n856 B.n855 585
R524 B.n552 B.n551 585
R525 B.n553 B.n552 585
R526 B.n864 B.n863 585
R527 B.n863 B.n862 585
R528 B.n865 B.n550 585
R529 B.n550 B.n549 585
R530 B.n867 B.n866 585
R531 B.n868 B.n867 585
R532 B.n544 B.n543 585
R533 B.n545 B.n544 585
R534 B.n876 B.n875 585
R535 B.n875 B.n874 585
R536 B.n877 B.n542 585
R537 B.n542 B.n541 585
R538 B.n879 B.n878 585
R539 B.n880 B.n879 585
R540 B.n536 B.n535 585
R541 B.n537 B.n536 585
R542 B.n888 B.n887 585
R543 B.n887 B.n886 585
R544 B.n889 B.n534 585
R545 B.n534 B.n533 585
R546 B.n891 B.n890 585
R547 B.n892 B.n891 585
R548 B.n528 B.n527 585
R549 B.n529 B.n528 585
R550 B.n900 B.n899 585
R551 B.n899 B.n898 585
R552 B.n901 B.n526 585
R553 B.n526 B.n525 585
R554 B.n903 B.n902 585
R555 B.n904 B.n903 585
R556 B.n520 B.n519 585
R557 B.n521 B.n520 585
R558 B.n912 B.n911 585
R559 B.n911 B.n910 585
R560 B.n913 B.n518 585
R561 B.n518 B.n517 585
R562 B.n915 B.n914 585
R563 B.n916 B.n915 585
R564 B.n512 B.n511 585
R565 B.n513 B.n512 585
R566 B.n924 B.n923 585
R567 B.n923 B.n922 585
R568 B.n925 B.n510 585
R569 B.n510 B.n509 585
R570 B.n927 B.n926 585
R571 B.n928 B.n927 585
R572 B.n504 B.n503 585
R573 B.n505 B.n504 585
R574 B.n936 B.n935 585
R575 B.n935 B.n934 585
R576 B.n937 B.n502 585
R577 B.n502 B.n501 585
R578 B.n939 B.n938 585
R579 B.n940 B.n939 585
R580 B.n496 B.n495 585
R581 B.n497 B.n496 585
R582 B.n948 B.n947 585
R583 B.n947 B.n946 585
R584 B.n949 B.n494 585
R585 B.n494 B.n493 585
R586 B.n951 B.n950 585
R587 B.n952 B.n951 585
R588 B.n488 B.n487 585
R589 B.n489 B.n488 585
R590 B.n960 B.n959 585
R591 B.n959 B.n958 585
R592 B.n961 B.n486 585
R593 B.n486 B.n484 585
R594 B.n963 B.n962 585
R595 B.n964 B.n963 585
R596 B.n480 B.n479 585
R597 B.n485 B.n480 585
R598 B.n972 B.n971 585
R599 B.n971 B.n970 585
R600 B.n973 B.n478 585
R601 B.n478 B.n477 585
R602 B.n975 B.n974 585
R603 B.n976 B.n975 585
R604 B.n472 B.n471 585
R605 B.n473 B.n472 585
R606 B.n984 B.n983 585
R607 B.n983 B.n982 585
R608 B.n985 B.n470 585
R609 B.n470 B.n469 585
R610 B.n987 B.n986 585
R611 B.n988 B.n987 585
R612 B.n464 B.n463 585
R613 B.n465 B.n464 585
R614 B.n996 B.n995 585
R615 B.n995 B.n994 585
R616 B.n997 B.n462 585
R617 B.n462 B.n460 585
R618 B.n999 B.n998 585
R619 B.n1000 B.n999 585
R620 B.n456 B.n455 585
R621 B.n461 B.n456 585
R622 B.n1008 B.n1007 585
R623 B.n1007 B.n1006 585
R624 B.n1009 B.n454 585
R625 B.n454 B.n453 585
R626 B.n1011 B.n1010 585
R627 B.n1012 B.n1011 585
R628 B.n448 B.n447 585
R629 B.n449 B.n448 585
R630 B.n1020 B.n1019 585
R631 B.n1019 B.n1018 585
R632 B.n1021 B.n446 585
R633 B.n446 B.n445 585
R634 B.n1023 B.n1022 585
R635 B.n1024 B.n1023 585
R636 B.n440 B.n439 585
R637 B.n441 B.n440 585
R638 B.n1032 B.n1031 585
R639 B.n1031 B.n1030 585
R640 B.n1033 B.n438 585
R641 B.n438 B.n437 585
R642 B.n1035 B.n1034 585
R643 B.n1036 B.n1035 585
R644 B.n432 B.n431 585
R645 B.n433 B.n432 585
R646 B.n1044 B.n1043 585
R647 B.n1043 B.n1042 585
R648 B.n1045 B.n430 585
R649 B.n430 B.n429 585
R650 B.n1047 B.n1046 585
R651 B.n1048 B.n1047 585
R652 B.n424 B.n423 585
R653 B.n425 B.n424 585
R654 B.n1057 B.n1056 585
R655 B.n1056 B.n1055 585
R656 B.n1058 B.n422 585
R657 B.n422 B.n421 585
R658 B.n1060 B.n1059 585
R659 B.n1061 B.n1060 585
R660 B.n3 B.n0 585
R661 B.n4 B.n3 585
R662 B.n1301 B.n1 585
R663 B.n1302 B.n1301 585
R664 B.n1300 B.n1299 585
R665 B.n1300 B.n8 585
R666 B.n1298 B.n9 585
R667 B.n12 B.n9 585
R668 B.n1297 B.n1296 585
R669 B.n1296 B.n1295 585
R670 B.n11 B.n10 585
R671 B.n1294 B.n11 585
R672 B.n1292 B.n1291 585
R673 B.n1293 B.n1292 585
R674 B.n1290 B.n17 585
R675 B.n17 B.n16 585
R676 B.n1289 B.n1288 585
R677 B.n1288 B.n1287 585
R678 B.n19 B.n18 585
R679 B.n1286 B.n19 585
R680 B.n1284 B.n1283 585
R681 B.n1285 B.n1284 585
R682 B.n1282 B.n24 585
R683 B.n24 B.n23 585
R684 B.n1281 B.n1280 585
R685 B.n1280 B.n1279 585
R686 B.n26 B.n25 585
R687 B.n1278 B.n26 585
R688 B.n1276 B.n1275 585
R689 B.n1277 B.n1276 585
R690 B.n1274 B.n31 585
R691 B.n31 B.n30 585
R692 B.n1273 B.n1272 585
R693 B.n1272 B.n1271 585
R694 B.n33 B.n32 585
R695 B.n1270 B.n33 585
R696 B.n1268 B.n1267 585
R697 B.n1269 B.n1268 585
R698 B.n1266 B.n38 585
R699 B.n38 B.n37 585
R700 B.n1265 B.n1264 585
R701 B.n1264 B.n1263 585
R702 B.n40 B.n39 585
R703 B.n1262 B.n40 585
R704 B.n1260 B.n1259 585
R705 B.n1261 B.n1260 585
R706 B.n1258 B.n45 585
R707 B.n45 B.n44 585
R708 B.n1257 B.n1256 585
R709 B.n1256 B.n1255 585
R710 B.n47 B.n46 585
R711 B.n1254 B.n47 585
R712 B.n1252 B.n1251 585
R713 B.n1253 B.n1252 585
R714 B.n1250 B.n52 585
R715 B.n52 B.n51 585
R716 B.n1249 B.n1248 585
R717 B.n1248 B.n1247 585
R718 B.n54 B.n53 585
R719 B.n1246 B.n54 585
R720 B.n1244 B.n1243 585
R721 B.n1245 B.n1244 585
R722 B.n1242 B.n59 585
R723 B.n59 B.n58 585
R724 B.n1241 B.n1240 585
R725 B.n1240 B.n1239 585
R726 B.n61 B.n60 585
R727 B.n1238 B.n61 585
R728 B.n1236 B.n1235 585
R729 B.n1237 B.n1236 585
R730 B.n1234 B.n66 585
R731 B.n66 B.n65 585
R732 B.n1233 B.n1232 585
R733 B.n1232 B.n1231 585
R734 B.n68 B.n67 585
R735 B.n1230 B.n68 585
R736 B.n1228 B.n1227 585
R737 B.n1229 B.n1228 585
R738 B.n1226 B.n73 585
R739 B.n73 B.n72 585
R740 B.n1225 B.n1224 585
R741 B.n1224 B.n1223 585
R742 B.n75 B.n74 585
R743 B.n1222 B.n75 585
R744 B.n1220 B.n1219 585
R745 B.n1221 B.n1220 585
R746 B.n1218 B.n80 585
R747 B.n80 B.n79 585
R748 B.n1217 B.n1216 585
R749 B.n1216 B.n1215 585
R750 B.n82 B.n81 585
R751 B.n1214 B.n82 585
R752 B.n1212 B.n1211 585
R753 B.n1213 B.n1212 585
R754 B.n1210 B.n87 585
R755 B.n87 B.n86 585
R756 B.n1209 B.n1208 585
R757 B.n1208 B.n1207 585
R758 B.n89 B.n88 585
R759 B.n1206 B.n89 585
R760 B.n1204 B.n1203 585
R761 B.n1205 B.n1204 585
R762 B.n1202 B.n94 585
R763 B.n94 B.n93 585
R764 B.n1201 B.n1200 585
R765 B.n1200 B.n1199 585
R766 B.n96 B.n95 585
R767 B.n1198 B.n96 585
R768 B.n1196 B.n1195 585
R769 B.n1197 B.n1196 585
R770 B.n1194 B.n101 585
R771 B.n101 B.n100 585
R772 B.n1193 B.n1192 585
R773 B.n1192 B.n1191 585
R774 B.n103 B.n102 585
R775 B.n1190 B.n103 585
R776 B.n1188 B.n1187 585
R777 B.n1189 B.n1188 585
R778 B.n1186 B.n108 585
R779 B.n108 B.n107 585
R780 B.n1185 B.n1184 585
R781 B.n1184 B.n1183 585
R782 B.n110 B.n109 585
R783 B.n1182 B.n110 585
R784 B.n1180 B.n1179 585
R785 B.n1181 B.n1180 585
R786 B.n1178 B.n115 585
R787 B.n115 B.n114 585
R788 B.n1177 B.n1176 585
R789 B.n1176 B.n1175 585
R790 B.n117 B.n116 585
R791 B.n1174 B.n117 585
R792 B.n1172 B.n1171 585
R793 B.n1173 B.n1172 585
R794 B.n1170 B.n122 585
R795 B.n122 B.n121 585
R796 B.n1169 B.n1168 585
R797 B.n1168 B.n1167 585
R798 B.n124 B.n123 585
R799 B.n1166 B.n124 585
R800 B.n1164 B.n1163 585
R801 B.n1165 B.n1164 585
R802 B.n1162 B.n129 585
R803 B.n129 B.n128 585
R804 B.n1305 B.n1304 585
R805 B.n1303 B.n2 585
R806 B.n1160 B.n129 468.476
R807 B.n1157 B.n189 468.476
R808 B.n623 B.n556 468.476
R809 B.n851 B.n558 468.476
R810 B.n193 B.t8 304.606
R811 B.n190 B.t19 304.606
R812 B.n621 B.t12 304.606
R813 B.n618 B.t16 304.606
R814 B.n1158 B.n187 256.663
R815 B.n1158 B.n186 256.663
R816 B.n1158 B.n185 256.663
R817 B.n1158 B.n184 256.663
R818 B.n1158 B.n183 256.663
R819 B.n1158 B.n182 256.663
R820 B.n1158 B.n181 256.663
R821 B.n1158 B.n180 256.663
R822 B.n1158 B.n179 256.663
R823 B.n1158 B.n178 256.663
R824 B.n1158 B.n177 256.663
R825 B.n1158 B.n176 256.663
R826 B.n1158 B.n175 256.663
R827 B.n1158 B.n174 256.663
R828 B.n1158 B.n173 256.663
R829 B.n1158 B.n172 256.663
R830 B.n1158 B.n171 256.663
R831 B.n1158 B.n170 256.663
R832 B.n1158 B.n169 256.663
R833 B.n1158 B.n168 256.663
R834 B.n1158 B.n167 256.663
R835 B.n1158 B.n166 256.663
R836 B.n1158 B.n165 256.663
R837 B.n1158 B.n164 256.663
R838 B.n1158 B.n163 256.663
R839 B.n1158 B.n162 256.663
R840 B.n1158 B.n161 256.663
R841 B.n1158 B.n160 256.663
R842 B.n1158 B.n159 256.663
R843 B.n1158 B.n158 256.663
R844 B.n1158 B.n157 256.663
R845 B.n1158 B.n156 256.663
R846 B.n1158 B.n155 256.663
R847 B.n1158 B.n154 256.663
R848 B.n1158 B.n153 256.663
R849 B.n1158 B.n152 256.663
R850 B.n1158 B.n151 256.663
R851 B.n1158 B.n150 256.663
R852 B.n1158 B.n149 256.663
R853 B.n1158 B.n148 256.663
R854 B.n1158 B.n147 256.663
R855 B.n1158 B.n146 256.663
R856 B.n1158 B.n145 256.663
R857 B.n1158 B.n144 256.663
R858 B.n1158 B.n143 256.663
R859 B.n1158 B.n142 256.663
R860 B.n1158 B.n141 256.663
R861 B.n1158 B.n140 256.663
R862 B.n1158 B.n139 256.663
R863 B.n1158 B.n138 256.663
R864 B.n1158 B.n137 256.663
R865 B.n1158 B.n136 256.663
R866 B.n1158 B.n135 256.663
R867 B.n1158 B.n134 256.663
R868 B.n1158 B.n133 256.663
R869 B.n1158 B.n132 256.663
R870 B.n1159 B.n1158 256.663
R871 B.n850 B.n849 256.663
R872 B.n849 B.n561 256.663
R873 B.n849 B.n562 256.663
R874 B.n849 B.n563 256.663
R875 B.n849 B.n564 256.663
R876 B.n849 B.n565 256.663
R877 B.n849 B.n566 256.663
R878 B.n849 B.n567 256.663
R879 B.n849 B.n568 256.663
R880 B.n849 B.n569 256.663
R881 B.n849 B.n570 256.663
R882 B.n849 B.n571 256.663
R883 B.n849 B.n572 256.663
R884 B.n849 B.n573 256.663
R885 B.n849 B.n574 256.663
R886 B.n849 B.n575 256.663
R887 B.n849 B.n576 256.663
R888 B.n849 B.n577 256.663
R889 B.n849 B.n578 256.663
R890 B.n849 B.n579 256.663
R891 B.n849 B.n580 256.663
R892 B.n849 B.n581 256.663
R893 B.n849 B.n582 256.663
R894 B.n849 B.n583 256.663
R895 B.n849 B.n584 256.663
R896 B.n849 B.n585 256.663
R897 B.n849 B.n586 256.663
R898 B.n849 B.n587 256.663
R899 B.n849 B.n588 256.663
R900 B.n849 B.n589 256.663
R901 B.n849 B.n590 256.663
R902 B.n849 B.n591 256.663
R903 B.n849 B.n592 256.663
R904 B.n849 B.n593 256.663
R905 B.n849 B.n594 256.663
R906 B.n849 B.n595 256.663
R907 B.n849 B.n596 256.663
R908 B.n849 B.n597 256.663
R909 B.n849 B.n598 256.663
R910 B.n849 B.n599 256.663
R911 B.n849 B.n600 256.663
R912 B.n849 B.n601 256.663
R913 B.n849 B.n602 256.663
R914 B.n849 B.n603 256.663
R915 B.n849 B.n604 256.663
R916 B.n849 B.n605 256.663
R917 B.n849 B.n606 256.663
R918 B.n849 B.n607 256.663
R919 B.n849 B.n608 256.663
R920 B.n849 B.n609 256.663
R921 B.n849 B.n610 256.663
R922 B.n849 B.n611 256.663
R923 B.n849 B.n612 256.663
R924 B.n849 B.n613 256.663
R925 B.n849 B.n614 256.663
R926 B.n849 B.n615 256.663
R927 B.n849 B.n616 256.663
R928 B.n1307 B.n1306 256.663
R929 B.n195 B.n131 163.367
R930 B.n199 B.n198 163.367
R931 B.n203 B.n202 163.367
R932 B.n207 B.n206 163.367
R933 B.n211 B.n210 163.367
R934 B.n215 B.n214 163.367
R935 B.n219 B.n218 163.367
R936 B.n223 B.n222 163.367
R937 B.n227 B.n226 163.367
R938 B.n231 B.n230 163.367
R939 B.n235 B.n234 163.367
R940 B.n239 B.n238 163.367
R941 B.n243 B.n242 163.367
R942 B.n247 B.n246 163.367
R943 B.n251 B.n250 163.367
R944 B.n255 B.n254 163.367
R945 B.n259 B.n258 163.367
R946 B.n263 B.n262 163.367
R947 B.n267 B.n266 163.367
R948 B.n271 B.n270 163.367
R949 B.n275 B.n274 163.367
R950 B.n279 B.n278 163.367
R951 B.n283 B.n282 163.367
R952 B.n287 B.n286 163.367
R953 B.n291 B.n290 163.367
R954 B.n295 B.n294 163.367
R955 B.n300 B.n299 163.367
R956 B.n304 B.n303 163.367
R957 B.n308 B.n307 163.367
R958 B.n312 B.n311 163.367
R959 B.n316 B.n315 163.367
R960 B.n320 B.n319 163.367
R961 B.n324 B.n323 163.367
R962 B.n328 B.n327 163.367
R963 B.n332 B.n331 163.367
R964 B.n336 B.n335 163.367
R965 B.n340 B.n339 163.367
R966 B.n344 B.n343 163.367
R967 B.n348 B.n347 163.367
R968 B.n352 B.n351 163.367
R969 B.n356 B.n355 163.367
R970 B.n360 B.n359 163.367
R971 B.n364 B.n363 163.367
R972 B.n368 B.n367 163.367
R973 B.n372 B.n371 163.367
R974 B.n376 B.n375 163.367
R975 B.n380 B.n379 163.367
R976 B.n384 B.n383 163.367
R977 B.n388 B.n387 163.367
R978 B.n392 B.n391 163.367
R979 B.n396 B.n395 163.367
R980 B.n400 B.n399 163.367
R981 B.n404 B.n403 163.367
R982 B.n408 B.n407 163.367
R983 B.n412 B.n411 163.367
R984 B.n416 B.n415 163.367
R985 B.n1157 B.n188 163.367
R986 B.n857 B.n556 163.367
R987 B.n857 B.n554 163.367
R988 B.n861 B.n554 163.367
R989 B.n861 B.n548 163.367
R990 B.n869 B.n548 163.367
R991 B.n869 B.n546 163.367
R992 B.n873 B.n546 163.367
R993 B.n873 B.n540 163.367
R994 B.n881 B.n540 163.367
R995 B.n881 B.n538 163.367
R996 B.n885 B.n538 163.367
R997 B.n885 B.n532 163.367
R998 B.n893 B.n532 163.367
R999 B.n893 B.n530 163.367
R1000 B.n897 B.n530 163.367
R1001 B.n897 B.n524 163.367
R1002 B.n905 B.n524 163.367
R1003 B.n905 B.n522 163.367
R1004 B.n909 B.n522 163.367
R1005 B.n909 B.n516 163.367
R1006 B.n917 B.n516 163.367
R1007 B.n917 B.n514 163.367
R1008 B.n921 B.n514 163.367
R1009 B.n921 B.n508 163.367
R1010 B.n929 B.n508 163.367
R1011 B.n929 B.n506 163.367
R1012 B.n933 B.n506 163.367
R1013 B.n933 B.n500 163.367
R1014 B.n941 B.n500 163.367
R1015 B.n941 B.n498 163.367
R1016 B.n945 B.n498 163.367
R1017 B.n945 B.n492 163.367
R1018 B.n953 B.n492 163.367
R1019 B.n953 B.n490 163.367
R1020 B.n957 B.n490 163.367
R1021 B.n957 B.n483 163.367
R1022 B.n965 B.n483 163.367
R1023 B.n965 B.n481 163.367
R1024 B.n969 B.n481 163.367
R1025 B.n969 B.n476 163.367
R1026 B.n977 B.n476 163.367
R1027 B.n977 B.n474 163.367
R1028 B.n981 B.n474 163.367
R1029 B.n981 B.n468 163.367
R1030 B.n989 B.n468 163.367
R1031 B.n989 B.n466 163.367
R1032 B.n993 B.n466 163.367
R1033 B.n993 B.n459 163.367
R1034 B.n1001 B.n459 163.367
R1035 B.n1001 B.n457 163.367
R1036 B.n1005 B.n457 163.367
R1037 B.n1005 B.n452 163.367
R1038 B.n1013 B.n452 163.367
R1039 B.n1013 B.n450 163.367
R1040 B.n1017 B.n450 163.367
R1041 B.n1017 B.n444 163.367
R1042 B.n1025 B.n444 163.367
R1043 B.n1025 B.n442 163.367
R1044 B.n1029 B.n442 163.367
R1045 B.n1029 B.n436 163.367
R1046 B.n1037 B.n436 163.367
R1047 B.n1037 B.n434 163.367
R1048 B.n1041 B.n434 163.367
R1049 B.n1041 B.n428 163.367
R1050 B.n1049 B.n428 163.367
R1051 B.n1049 B.n426 163.367
R1052 B.n1054 B.n426 163.367
R1053 B.n1054 B.n420 163.367
R1054 B.n1062 B.n420 163.367
R1055 B.n1063 B.n1062 163.367
R1056 B.n1063 B.n5 163.367
R1057 B.n6 B.n5 163.367
R1058 B.n7 B.n6 163.367
R1059 B.n1069 B.n7 163.367
R1060 B.n1070 B.n1069 163.367
R1061 B.n1070 B.n13 163.367
R1062 B.n14 B.n13 163.367
R1063 B.n15 B.n14 163.367
R1064 B.n1075 B.n15 163.367
R1065 B.n1075 B.n20 163.367
R1066 B.n21 B.n20 163.367
R1067 B.n22 B.n21 163.367
R1068 B.n1080 B.n22 163.367
R1069 B.n1080 B.n27 163.367
R1070 B.n28 B.n27 163.367
R1071 B.n29 B.n28 163.367
R1072 B.n1085 B.n29 163.367
R1073 B.n1085 B.n34 163.367
R1074 B.n35 B.n34 163.367
R1075 B.n36 B.n35 163.367
R1076 B.n1090 B.n36 163.367
R1077 B.n1090 B.n41 163.367
R1078 B.n42 B.n41 163.367
R1079 B.n43 B.n42 163.367
R1080 B.n1095 B.n43 163.367
R1081 B.n1095 B.n48 163.367
R1082 B.n49 B.n48 163.367
R1083 B.n50 B.n49 163.367
R1084 B.n1100 B.n50 163.367
R1085 B.n1100 B.n55 163.367
R1086 B.n56 B.n55 163.367
R1087 B.n57 B.n56 163.367
R1088 B.n1105 B.n57 163.367
R1089 B.n1105 B.n62 163.367
R1090 B.n63 B.n62 163.367
R1091 B.n64 B.n63 163.367
R1092 B.n1110 B.n64 163.367
R1093 B.n1110 B.n69 163.367
R1094 B.n70 B.n69 163.367
R1095 B.n71 B.n70 163.367
R1096 B.n1115 B.n71 163.367
R1097 B.n1115 B.n76 163.367
R1098 B.n77 B.n76 163.367
R1099 B.n78 B.n77 163.367
R1100 B.n1120 B.n78 163.367
R1101 B.n1120 B.n83 163.367
R1102 B.n84 B.n83 163.367
R1103 B.n85 B.n84 163.367
R1104 B.n1125 B.n85 163.367
R1105 B.n1125 B.n90 163.367
R1106 B.n91 B.n90 163.367
R1107 B.n92 B.n91 163.367
R1108 B.n1130 B.n92 163.367
R1109 B.n1130 B.n97 163.367
R1110 B.n98 B.n97 163.367
R1111 B.n99 B.n98 163.367
R1112 B.n1135 B.n99 163.367
R1113 B.n1135 B.n104 163.367
R1114 B.n105 B.n104 163.367
R1115 B.n106 B.n105 163.367
R1116 B.n1140 B.n106 163.367
R1117 B.n1140 B.n111 163.367
R1118 B.n112 B.n111 163.367
R1119 B.n113 B.n112 163.367
R1120 B.n1145 B.n113 163.367
R1121 B.n1145 B.n118 163.367
R1122 B.n119 B.n118 163.367
R1123 B.n120 B.n119 163.367
R1124 B.n1150 B.n120 163.367
R1125 B.n1150 B.n125 163.367
R1126 B.n126 B.n125 163.367
R1127 B.n127 B.n126 163.367
R1128 B.n189 B.n127 163.367
R1129 B.n848 B.n560 163.367
R1130 B.n848 B.n617 163.367
R1131 B.n844 B.n843 163.367
R1132 B.n840 B.n839 163.367
R1133 B.n836 B.n835 163.367
R1134 B.n832 B.n831 163.367
R1135 B.n828 B.n827 163.367
R1136 B.n824 B.n823 163.367
R1137 B.n820 B.n819 163.367
R1138 B.n816 B.n815 163.367
R1139 B.n812 B.n811 163.367
R1140 B.n808 B.n807 163.367
R1141 B.n804 B.n803 163.367
R1142 B.n800 B.n799 163.367
R1143 B.n796 B.n795 163.367
R1144 B.n792 B.n791 163.367
R1145 B.n788 B.n787 163.367
R1146 B.n784 B.n783 163.367
R1147 B.n780 B.n779 163.367
R1148 B.n776 B.n775 163.367
R1149 B.n772 B.n771 163.367
R1150 B.n768 B.n767 163.367
R1151 B.n764 B.n763 163.367
R1152 B.n760 B.n759 163.367
R1153 B.n756 B.n755 163.367
R1154 B.n752 B.n751 163.367
R1155 B.n748 B.n747 163.367
R1156 B.n744 B.n743 163.367
R1157 B.n740 B.n739 163.367
R1158 B.n736 B.n735 163.367
R1159 B.n732 B.n731 163.367
R1160 B.n727 B.n726 163.367
R1161 B.n723 B.n722 163.367
R1162 B.n719 B.n718 163.367
R1163 B.n715 B.n714 163.367
R1164 B.n711 B.n710 163.367
R1165 B.n707 B.n706 163.367
R1166 B.n703 B.n702 163.367
R1167 B.n699 B.n698 163.367
R1168 B.n695 B.n694 163.367
R1169 B.n691 B.n690 163.367
R1170 B.n687 B.n686 163.367
R1171 B.n683 B.n682 163.367
R1172 B.n679 B.n678 163.367
R1173 B.n675 B.n674 163.367
R1174 B.n671 B.n670 163.367
R1175 B.n667 B.n666 163.367
R1176 B.n663 B.n662 163.367
R1177 B.n659 B.n658 163.367
R1178 B.n655 B.n654 163.367
R1179 B.n651 B.n650 163.367
R1180 B.n647 B.n646 163.367
R1181 B.n643 B.n642 163.367
R1182 B.n639 B.n638 163.367
R1183 B.n635 B.n634 163.367
R1184 B.n631 B.n630 163.367
R1185 B.n627 B.n626 163.367
R1186 B.n855 B.n558 163.367
R1187 B.n855 B.n552 163.367
R1188 B.n863 B.n552 163.367
R1189 B.n863 B.n550 163.367
R1190 B.n867 B.n550 163.367
R1191 B.n867 B.n544 163.367
R1192 B.n875 B.n544 163.367
R1193 B.n875 B.n542 163.367
R1194 B.n879 B.n542 163.367
R1195 B.n879 B.n536 163.367
R1196 B.n887 B.n536 163.367
R1197 B.n887 B.n534 163.367
R1198 B.n891 B.n534 163.367
R1199 B.n891 B.n528 163.367
R1200 B.n899 B.n528 163.367
R1201 B.n899 B.n526 163.367
R1202 B.n903 B.n526 163.367
R1203 B.n903 B.n520 163.367
R1204 B.n911 B.n520 163.367
R1205 B.n911 B.n518 163.367
R1206 B.n915 B.n518 163.367
R1207 B.n915 B.n512 163.367
R1208 B.n923 B.n512 163.367
R1209 B.n923 B.n510 163.367
R1210 B.n927 B.n510 163.367
R1211 B.n927 B.n504 163.367
R1212 B.n935 B.n504 163.367
R1213 B.n935 B.n502 163.367
R1214 B.n939 B.n502 163.367
R1215 B.n939 B.n496 163.367
R1216 B.n947 B.n496 163.367
R1217 B.n947 B.n494 163.367
R1218 B.n951 B.n494 163.367
R1219 B.n951 B.n488 163.367
R1220 B.n959 B.n488 163.367
R1221 B.n959 B.n486 163.367
R1222 B.n963 B.n486 163.367
R1223 B.n963 B.n480 163.367
R1224 B.n971 B.n480 163.367
R1225 B.n971 B.n478 163.367
R1226 B.n975 B.n478 163.367
R1227 B.n975 B.n472 163.367
R1228 B.n983 B.n472 163.367
R1229 B.n983 B.n470 163.367
R1230 B.n987 B.n470 163.367
R1231 B.n987 B.n464 163.367
R1232 B.n995 B.n464 163.367
R1233 B.n995 B.n462 163.367
R1234 B.n999 B.n462 163.367
R1235 B.n999 B.n456 163.367
R1236 B.n1007 B.n456 163.367
R1237 B.n1007 B.n454 163.367
R1238 B.n1011 B.n454 163.367
R1239 B.n1011 B.n448 163.367
R1240 B.n1019 B.n448 163.367
R1241 B.n1019 B.n446 163.367
R1242 B.n1023 B.n446 163.367
R1243 B.n1023 B.n440 163.367
R1244 B.n1031 B.n440 163.367
R1245 B.n1031 B.n438 163.367
R1246 B.n1035 B.n438 163.367
R1247 B.n1035 B.n432 163.367
R1248 B.n1043 B.n432 163.367
R1249 B.n1043 B.n430 163.367
R1250 B.n1047 B.n430 163.367
R1251 B.n1047 B.n424 163.367
R1252 B.n1056 B.n424 163.367
R1253 B.n1056 B.n422 163.367
R1254 B.n1060 B.n422 163.367
R1255 B.n1060 B.n3 163.367
R1256 B.n1305 B.n3 163.367
R1257 B.n1301 B.n2 163.367
R1258 B.n1301 B.n1300 163.367
R1259 B.n1300 B.n9 163.367
R1260 B.n1296 B.n9 163.367
R1261 B.n1296 B.n11 163.367
R1262 B.n1292 B.n11 163.367
R1263 B.n1292 B.n17 163.367
R1264 B.n1288 B.n17 163.367
R1265 B.n1288 B.n19 163.367
R1266 B.n1284 B.n19 163.367
R1267 B.n1284 B.n24 163.367
R1268 B.n1280 B.n24 163.367
R1269 B.n1280 B.n26 163.367
R1270 B.n1276 B.n26 163.367
R1271 B.n1276 B.n31 163.367
R1272 B.n1272 B.n31 163.367
R1273 B.n1272 B.n33 163.367
R1274 B.n1268 B.n33 163.367
R1275 B.n1268 B.n38 163.367
R1276 B.n1264 B.n38 163.367
R1277 B.n1264 B.n40 163.367
R1278 B.n1260 B.n40 163.367
R1279 B.n1260 B.n45 163.367
R1280 B.n1256 B.n45 163.367
R1281 B.n1256 B.n47 163.367
R1282 B.n1252 B.n47 163.367
R1283 B.n1252 B.n52 163.367
R1284 B.n1248 B.n52 163.367
R1285 B.n1248 B.n54 163.367
R1286 B.n1244 B.n54 163.367
R1287 B.n1244 B.n59 163.367
R1288 B.n1240 B.n59 163.367
R1289 B.n1240 B.n61 163.367
R1290 B.n1236 B.n61 163.367
R1291 B.n1236 B.n66 163.367
R1292 B.n1232 B.n66 163.367
R1293 B.n1232 B.n68 163.367
R1294 B.n1228 B.n68 163.367
R1295 B.n1228 B.n73 163.367
R1296 B.n1224 B.n73 163.367
R1297 B.n1224 B.n75 163.367
R1298 B.n1220 B.n75 163.367
R1299 B.n1220 B.n80 163.367
R1300 B.n1216 B.n80 163.367
R1301 B.n1216 B.n82 163.367
R1302 B.n1212 B.n82 163.367
R1303 B.n1212 B.n87 163.367
R1304 B.n1208 B.n87 163.367
R1305 B.n1208 B.n89 163.367
R1306 B.n1204 B.n89 163.367
R1307 B.n1204 B.n94 163.367
R1308 B.n1200 B.n94 163.367
R1309 B.n1200 B.n96 163.367
R1310 B.n1196 B.n96 163.367
R1311 B.n1196 B.n101 163.367
R1312 B.n1192 B.n101 163.367
R1313 B.n1192 B.n103 163.367
R1314 B.n1188 B.n103 163.367
R1315 B.n1188 B.n108 163.367
R1316 B.n1184 B.n108 163.367
R1317 B.n1184 B.n110 163.367
R1318 B.n1180 B.n110 163.367
R1319 B.n1180 B.n115 163.367
R1320 B.n1176 B.n115 163.367
R1321 B.n1176 B.n117 163.367
R1322 B.n1172 B.n117 163.367
R1323 B.n1172 B.n122 163.367
R1324 B.n1168 B.n122 163.367
R1325 B.n1168 B.n124 163.367
R1326 B.n1164 B.n124 163.367
R1327 B.n1164 B.n129 163.367
R1328 B.n190 B.t20 152.351
R1329 B.n621 B.t15 152.351
R1330 B.n193 B.t10 152.331
R1331 B.n618 B.t18 152.331
R1332 B.n194 B.n193 83.5884
R1333 B.n191 B.n190 83.5884
R1334 B.n622 B.n621 83.5884
R1335 B.n619 B.n618 83.5884
R1336 B.n1160 B.n1159 71.676
R1337 B.n195 B.n132 71.676
R1338 B.n199 B.n133 71.676
R1339 B.n203 B.n134 71.676
R1340 B.n207 B.n135 71.676
R1341 B.n211 B.n136 71.676
R1342 B.n215 B.n137 71.676
R1343 B.n219 B.n138 71.676
R1344 B.n223 B.n139 71.676
R1345 B.n227 B.n140 71.676
R1346 B.n231 B.n141 71.676
R1347 B.n235 B.n142 71.676
R1348 B.n239 B.n143 71.676
R1349 B.n243 B.n144 71.676
R1350 B.n247 B.n145 71.676
R1351 B.n251 B.n146 71.676
R1352 B.n255 B.n147 71.676
R1353 B.n259 B.n148 71.676
R1354 B.n263 B.n149 71.676
R1355 B.n267 B.n150 71.676
R1356 B.n271 B.n151 71.676
R1357 B.n275 B.n152 71.676
R1358 B.n279 B.n153 71.676
R1359 B.n283 B.n154 71.676
R1360 B.n287 B.n155 71.676
R1361 B.n291 B.n156 71.676
R1362 B.n295 B.n157 71.676
R1363 B.n300 B.n158 71.676
R1364 B.n304 B.n159 71.676
R1365 B.n308 B.n160 71.676
R1366 B.n312 B.n161 71.676
R1367 B.n316 B.n162 71.676
R1368 B.n320 B.n163 71.676
R1369 B.n324 B.n164 71.676
R1370 B.n328 B.n165 71.676
R1371 B.n332 B.n166 71.676
R1372 B.n336 B.n167 71.676
R1373 B.n340 B.n168 71.676
R1374 B.n344 B.n169 71.676
R1375 B.n348 B.n170 71.676
R1376 B.n352 B.n171 71.676
R1377 B.n356 B.n172 71.676
R1378 B.n360 B.n173 71.676
R1379 B.n364 B.n174 71.676
R1380 B.n368 B.n175 71.676
R1381 B.n372 B.n176 71.676
R1382 B.n376 B.n177 71.676
R1383 B.n380 B.n178 71.676
R1384 B.n384 B.n179 71.676
R1385 B.n388 B.n180 71.676
R1386 B.n392 B.n181 71.676
R1387 B.n396 B.n182 71.676
R1388 B.n400 B.n183 71.676
R1389 B.n404 B.n184 71.676
R1390 B.n408 B.n185 71.676
R1391 B.n412 B.n186 71.676
R1392 B.n416 B.n187 71.676
R1393 B.n188 B.n187 71.676
R1394 B.n415 B.n186 71.676
R1395 B.n411 B.n185 71.676
R1396 B.n407 B.n184 71.676
R1397 B.n403 B.n183 71.676
R1398 B.n399 B.n182 71.676
R1399 B.n395 B.n181 71.676
R1400 B.n391 B.n180 71.676
R1401 B.n387 B.n179 71.676
R1402 B.n383 B.n178 71.676
R1403 B.n379 B.n177 71.676
R1404 B.n375 B.n176 71.676
R1405 B.n371 B.n175 71.676
R1406 B.n367 B.n174 71.676
R1407 B.n363 B.n173 71.676
R1408 B.n359 B.n172 71.676
R1409 B.n355 B.n171 71.676
R1410 B.n351 B.n170 71.676
R1411 B.n347 B.n169 71.676
R1412 B.n343 B.n168 71.676
R1413 B.n339 B.n167 71.676
R1414 B.n335 B.n166 71.676
R1415 B.n331 B.n165 71.676
R1416 B.n327 B.n164 71.676
R1417 B.n323 B.n163 71.676
R1418 B.n319 B.n162 71.676
R1419 B.n315 B.n161 71.676
R1420 B.n311 B.n160 71.676
R1421 B.n307 B.n159 71.676
R1422 B.n303 B.n158 71.676
R1423 B.n299 B.n157 71.676
R1424 B.n294 B.n156 71.676
R1425 B.n290 B.n155 71.676
R1426 B.n286 B.n154 71.676
R1427 B.n282 B.n153 71.676
R1428 B.n278 B.n152 71.676
R1429 B.n274 B.n151 71.676
R1430 B.n270 B.n150 71.676
R1431 B.n266 B.n149 71.676
R1432 B.n262 B.n148 71.676
R1433 B.n258 B.n147 71.676
R1434 B.n254 B.n146 71.676
R1435 B.n250 B.n145 71.676
R1436 B.n246 B.n144 71.676
R1437 B.n242 B.n143 71.676
R1438 B.n238 B.n142 71.676
R1439 B.n234 B.n141 71.676
R1440 B.n230 B.n140 71.676
R1441 B.n226 B.n139 71.676
R1442 B.n222 B.n138 71.676
R1443 B.n218 B.n137 71.676
R1444 B.n214 B.n136 71.676
R1445 B.n210 B.n135 71.676
R1446 B.n206 B.n134 71.676
R1447 B.n202 B.n133 71.676
R1448 B.n198 B.n132 71.676
R1449 B.n1159 B.n131 71.676
R1450 B.n851 B.n850 71.676
R1451 B.n617 B.n561 71.676
R1452 B.n843 B.n562 71.676
R1453 B.n839 B.n563 71.676
R1454 B.n835 B.n564 71.676
R1455 B.n831 B.n565 71.676
R1456 B.n827 B.n566 71.676
R1457 B.n823 B.n567 71.676
R1458 B.n819 B.n568 71.676
R1459 B.n815 B.n569 71.676
R1460 B.n811 B.n570 71.676
R1461 B.n807 B.n571 71.676
R1462 B.n803 B.n572 71.676
R1463 B.n799 B.n573 71.676
R1464 B.n795 B.n574 71.676
R1465 B.n791 B.n575 71.676
R1466 B.n787 B.n576 71.676
R1467 B.n783 B.n577 71.676
R1468 B.n779 B.n578 71.676
R1469 B.n775 B.n579 71.676
R1470 B.n771 B.n580 71.676
R1471 B.n767 B.n581 71.676
R1472 B.n763 B.n582 71.676
R1473 B.n759 B.n583 71.676
R1474 B.n755 B.n584 71.676
R1475 B.n751 B.n585 71.676
R1476 B.n747 B.n586 71.676
R1477 B.n743 B.n587 71.676
R1478 B.n739 B.n588 71.676
R1479 B.n735 B.n589 71.676
R1480 B.n731 B.n590 71.676
R1481 B.n726 B.n591 71.676
R1482 B.n722 B.n592 71.676
R1483 B.n718 B.n593 71.676
R1484 B.n714 B.n594 71.676
R1485 B.n710 B.n595 71.676
R1486 B.n706 B.n596 71.676
R1487 B.n702 B.n597 71.676
R1488 B.n698 B.n598 71.676
R1489 B.n694 B.n599 71.676
R1490 B.n690 B.n600 71.676
R1491 B.n686 B.n601 71.676
R1492 B.n682 B.n602 71.676
R1493 B.n678 B.n603 71.676
R1494 B.n674 B.n604 71.676
R1495 B.n670 B.n605 71.676
R1496 B.n666 B.n606 71.676
R1497 B.n662 B.n607 71.676
R1498 B.n658 B.n608 71.676
R1499 B.n654 B.n609 71.676
R1500 B.n650 B.n610 71.676
R1501 B.n646 B.n611 71.676
R1502 B.n642 B.n612 71.676
R1503 B.n638 B.n613 71.676
R1504 B.n634 B.n614 71.676
R1505 B.n630 B.n615 71.676
R1506 B.n626 B.n616 71.676
R1507 B.n850 B.n560 71.676
R1508 B.n844 B.n561 71.676
R1509 B.n840 B.n562 71.676
R1510 B.n836 B.n563 71.676
R1511 B.n832 B.n564 71.676
R1512 B.n828 B.n565 71.676
R1513 B.n824 B.n566 71.676
R1514 B.n820 B.n567 71.676
R1515 B.n816 B.n568 71.676
R1516 B.n812 B.n569 71.676
R1517 B.n808 B.n570 71.676
R1518 B.n804 B.n571 71.676
R1519 B.n800 B.n572 71.676
R1520 B.n796 B.n573 71.676
R1521 B.n792 B.n574 71.676
R1522 B.n788 B.n575 71.676
R1523 B.n784 B.n576 71.676
R1524 B.n780 B.n577 71.676
R1525 B.n776 B.n578 71.676
R1526 B.n772 B.n579 71.676
R1527 B.n768 B.n580 71.676
R1528 B.n764 B.n581 71.676
R1529 B.n760 B.n582 71.676
R1530 B.n756 B.n583 71.676
R1531 B.n752 B.n584 71.676
R1532 B.n748 B.n585 71.676
R1533 B.n744 B.n586 71.676
R1534 B.n740 B.n587 71.676
R1535 B.n736 B.n588 71.676
R1536 B.n732 B.n589 71.676
R1537 B.n727 B.n590 71.676
R1538 B.n723 B.n591 71.676
R1539 B.n719 B.n592 71.676
R1540 B.n715 B.n593 71.676
R1541 B.n711 B.n594 71.676
R1542 B.n707 B.n595 71.676
R1543 B.n703 B.n596 71.676
R1544 B.n699 B.n597 71.676
R1545 B.n695 B.n598 71.676
R1546 B.n691 B.n599 71.676
R1547 B.n687 B.n600 71.676
R1548 B.n683 B.n601 71.676
R1549 B.n679 B.n602 71.676
R1550 B.n675 B.n603 71.676
R1551 B.n671 B.n604 71.676
R1552 B.n667 B.n605 71.676
R1553 B.n663 B.n606 71.676
R1554 B.n659 B.n607 71.676
R1555 B.n655 B.n608 71.676
R1556 B.n651 B.n609 71.676
R1557 B.n647 B.n610 71.676
R1558 B.n643 B.n611 71.676
R1559 B.n639 B.n612 71.676
R1560 B.n635 B.n613 71.676
R1561 B.n631 B.n614 71.676
R1562 B.n627 B.n615 71.676
R1563 B.n623 B.n616 71.676
R1564 B.n1306 B.n1305 71.676
R1565 B.n1306 B.n2 71.676
R1566 B.n191 B.t21 68.7633
R1567 B.n622 B.t14 68.7633
R1568 B.n194 B.t11 68.7426
R1569 B.n619 B.t17 68.7426
R1570 B.n849 B.n557 64.4751
R1571 B.n1158 B.n128 64.4751
R1572 B.n297 B.n194 59.5399
R1573 B.n192 B.n191 59.5399
R1574 B.n729 B.n622 59.5399
R1575 B.n620 B.n619 59.5399
R1576 B.n856 B.n557 35.645
R1577 B.n856 B.n553 35.645
R1578 B.n862 B.n553 35.645
R1579 B.n862 B.n549 35.645
R1580 B.n868 B.n549 35.645
R1581 B.n868 B.n545 35.645
R1582 B.n874 B.n545 35.645
R1583 B.n874 B.n541 35.645
R1584 B.n880 B.n541 35.645
R1585 B.n886 B.n537 35.645
R1586 B.n886 B.n533 35.645
R1587 B.n892 B.n533 35.645
R1588 B.n892 B.n529 35.645
R1589 B.n898 B.n529 35.645
R1590 B.n898 B.n525 35.645
R1591 B.n904 B.n525 35.645
R1592 B.n904 B.n521 35.645
R1593 B.n910 B.n521 35.645
R1594 B.n910 B.n517 35.645
R1595 B.n916 B.n517 35.645
R1596 B.n916 B.n513 35.645
R1597 B.n922 B.n513 35.645
R1598 B.n922 B.n509 35.645
R1599 B.n928 B.n509 35.645
R1600 B.n934 B.n505 35.645
R1601 B.n934 B.n501 35.645
R1602 B.n940 B.n501 35.645
R1603 B.n940 B.n497 35.645
R1604 B.n946 B.n497 35.645
R1605 B.n946 B.n493 35.645
R1606 B.n952 B.n493 35.645
R1607 B.n952 B.n489 35.645
R1608 B.n958 B.n489 35.645
R1609 B.n958 B.n484 35.645
R1610 B.n964 B.n484 35.645
R1611 B.n964 B.n485 35.645
R1612 B.n970 B.n477 35.645
R1613 B.n976 B.n477 35.645
R1614 B.n976 B.n473 35.645
R1615 B.n982 B.n473 35.645
R1616 B.n982 B.n469 35.645
R1617 B.n988 B.n469 35.645
R1618 B.n988 B.n465 35.645
R1619 B.n994 B.n465 35.645
R1620 B.n994 B.n460 35.645
R1621 B.n1000 B.n460 35.645
R1622 B.n1000 B.n461 35.645
R1623 B.n1006 B.n453 35.645
R1624 B.n1012 B.n453 35.645
R1625 B.n1012 B.n449 35.645
R1626 B.n1018 B.n449 35.645
R1627 B.n1018 B.n445 35.645
R1628 B.n1024 B.n445 35.645
R1629 B.n1024 B.n441 35.645
R1630 B.n1030 B.n441 35.645
R1631 B.n1030 B.n437 35.645
R1632 B.n1036 B.n437 35.645
R1633 B.n1036 B.n433 35.645
R1634 B.n1042 B.n433 35.645
R1635 B.n1048 B.n429 35.645
R1636 B.n1048 B.n425 35.645
R1637 B.n1055 B.n425 35.645
R1638 B.n1055 B.n421 35.645
R1639 B.n1061 B.n421 35.645
R1640 B.n1061 B.n4 35.645
R1641 B.n1304 B.n4 35.645
R1642 B.n1304 B.n1303 35.645
R1643 B.n1303 B.n1302 35.645
R1644 B.n1302 B.n8 35.645
R1645 B.n12 B.n8 35.645
R1646 B.n1295 B.n12 35.645
R1647 B.n1295 B.n1294 35.645
R1648 B.n1294 B.n1293 35.645
R1649 B.n1293 B.n16 35.645
R1650 B.n1287 B.n1286 35.645
R1651 B.n1286 B.n1285 35.645
R1652 B.n1285 B.n23 35.645
R1653 B.n1279 B.n23 35.645
R1654 B.n1279 B.n1278 35.645
R1655 B.n1278 B.n1277 35.645
R1656 B.n1277 B.n30 35.645
R1657 B.n1271 B.n30 35.645
R1658 B.n1271 B.n1270 35.645
R1659 B.n1270 B.n1269 35.645
R1660 B.n1269 B.n37 35.645
R1661 B.n1263 B.n37 35.645
R1662 B.n1262 B.n1261 35.645
R1663 B.n1261 B.n44 35.645
R1664 B.n1255 B.n44 35.645
R1665 B.n1255 B.n1254 35.645
R1666 B.n1254 B.n1253 35.645
R1667 B.n1253 B.n51 35.645
R1668 B.n1247 B.n51 35.645
R1669 B.n1247 B.n1246 35.645
R1670 B.n1246 B.n1245 35.645
R1671 B.n1245 B.n58 35.645
R1672 B.n1239 B.n58 35.645
R1673 B.n1238 B.n1237 35.645
R1674 B.n1237 B.n65 35.645
R1675 B.n1231 B.n65 35.645
R1676 B.n1231 B.n1230 35.645
R1677 B.n1230 B.n1229 35.645
R1678 B.n1229 B.n72 35.645
R1679 B.n1223 B.n72 35.645
R1680 B.n1223 B.n1222 35.645
R1681 B.n1222 B.n1221 35.645
R1682 B.n1221 B.n79 35.645
R1683 B.n1215 B.n79 35.645
R1684 B.n1215 B.n1214 35.645
R1685 B.n1213 B.n86 35.645
R1686 B.n1207 B.n86 35.645
R1687 B.n1207 B.n1206 35.645
R1688 B.n1206 B.n1205 35.645
R1689 B.n1205 B.n93 35.645
R1690 B.n1199 B.n93 35.645
R1691 B.n1199 B.n1198 35.645
R1692 B.n1198 B.n1197 35.645
R1693 B.n1197 B.n100 35.645
R1694 B.n1191 B.n100 35.645
R1695 B.n1191 B.n1190 35.645
R1696 B.n1190 B.n1189 35.645
R1697 B.n1189 B.n107 35.645
R1698 B.n1183 B.n107 35.645
R1699 B.n1183 B.n1182 35.645
R1700 B.n1181 B.n114 35.645
R1701 B.n1175 B.n114 35.645
R1702 B.n1175 B.n1174 35.645
R1703 B.n1174 B.n1173 35.645
R1704 B.n1173 B.n121 35.645
R1705 B.n1167 B.n121 35.645
R1706 B.n1167 B.n1166 35.645
R1707 B.n1166 B.n1165 35.645
R1708 B.n1165 B.n128 35.645
R1709 B.n461 B.t1 31.4515
R1710 B.t7 B.n1262 31.4515
R1711 B.n853 B.n852 30.4395
R1712 B.n624 B.n555 30.4395
R1713 B.n1156 B.n1155 30.4395
R1714 B.n1162 B.n1161 30.4395
R1715 B.n970 B.t3 28.3064
R1716 B.n1239 B.t4 28.3064
R1717 B.n880 B.t13 23.0646
R1718 B.t9 B.n1181 23.0646
R1719 B.n1042 B.t2 19.9195
R1720 B.n1287 B.t6 19.9195
R1721 B.n928 B.t5 18.8711
R1722 B.t0 B.n1213 18.8711
R1723 B B.n1307 18.0485
R1724 B.t5 B.n505 16.7744
R1725 B.n1214 B.t0 16.7744
R1726 B.t2 B.n429 15.726
R1727 B.t6 B.n16 15.726
R1728 B.t13 B.n537 12.5809
R1729 B.n1182 B.t9 12.5809
R1730 B.n854 B.n853 10.6151
R1731 B.n854 B.n551 10.6151
R1732 B.n864 B.n551 10.6151
R1733 B.n865 B.n864 10.6151
R1734 B.n866 B.n865 10.6151
R1735 B.n866 B.n543 10.6151
R1736 B.n876 B.n543 10.6151
R1737 B.n877 B.n876 10.6151
R1738 B.n878 B.n877 10.6151
R1739 B.n878 B.n535 10.6151
R1740 B.n888 B.n535 10.6151
R1741 B.n889 B.n888 10.6151
R1742 B.n890 B.n889 10.6151
R1743 B.n890 B.n527 10.6151
R1744 B.n900 B.n527 10.6151
R1745 B.n901 B.n900 10.6151
R1746 B.n902 B.n901 10.6151
R1747 B.n902 B.n519 10.6151
R1748 B.n912 B.n519 10.6151
R1749 B.n913 B.n912 10.6151
R1750 B.n914 B.n913 10.6151
R1751 B.n914 B.n511 10.6151
R1752 B.n924 B.n511 10.6151
R1753 B.n925 B.n924 10.6151
R1754 B.n926 B.n925 10.6151
R1755 B.n926 B.n503 10.6151
R1756 B.n936 B.n503 10.6151
R1757 B.n937 B.n936 10.6151
R1758 B.n938 B.n937 10.6151
R1759 B.n938 B.n495 10.6151
R1760 B.n948 B.n495 10.6151
R1761 B.n949 B.n948 10.6151
R1762 B.n950 B.n949 10.6151
R1763 B.n950 B.n487 10.6151
R1764 B.n960 B.n487 10.6151
R1765 B.n961 B.n960 10.6151
R1766 B.n962 B.n961 10.6151
R1767 B.n962 B.n479 10.6151
R1768 B.n972 B.n479 10.6151
R1769 B.n973 B.n972 10.6151
R1770 B.n974 B.n973 10.6151
R1771 B.n974 B.n471 10.6151
R1772 B.n984 B.n471 10.6151
R1773 B.n985 B.n984 10.6151
R1774 B.n986 B.n985 10.6151
R1775 B.n986 B.n463 10.6151
R1776 B.n996 B.n463 10.6151
R1777 B.n997 B.n996 10.6151
R1778 B.n998 B.n997 10.6151
R1779 B.n998 B.n455 10.6151
R1780 B.n1008 B.n455 10.6151
R1781 B.n1009 B.n1008 10.6151
R1782 B.n1010 B.n1009 10.6151
R1783 B.n1010 B.n447 10.6151
R1784 B.n1020 B.n447 10.6151
R1785 B.n1021 B.n1020 10.6151
R1786 B.n1022 B.n1021 10.6151
R1787 B.n1022 B.n439 10.6151
R1788 B.n1032 B.n439 10.6151
R1789 B.n1033 B.n1032 10.6151
R1790 B.n1034 B.n1033 10.6151
R1791 B.n1034 B.n431 10.6151
R1792 B.n1044 B.n431 10.6151
R1793 B.n1045 B.n1044 10.6151
R1794 B.n1046 B.n1045 10.6151
R1795 B.n1046 B.n423 10.6151
R1796 B.n1057 B.n423 10.6151
R1797 B.n1058 B.n1057 10.6151
R1798 B.n1059 B.n1058 10.6151
R1799 B.n1059 B.n0 10.6151
R1800 B.n852 B.n559 10.6151
R1801 B.n847 B.n559 10.6151
R1802 B.n847 B.n846 10.6151
R1803 B.n846 B.n845 10.6151
R1804 B.n845 B.n842 10.6151
R1805 B.n842 B.n841 10.6151
R1806 B.n841 B.n838 10.6151
R1807 B.n838 B.n837 10.6151
R1808 B.n837 B.n834 10.6151
R1809 B.n834 B.n833 10.6151
R1810 B.n833 B.n830 10.6151
R1811 B.n830 B.n829 10.6151
R1812 B.n829 B.n826 10.6151
R1813 B.n826 B.n825 10.6151
R1814 B.n825 B.n822 10.6151
R1815 B.n822 B.n821 10.6151
R1816 B.n821 B.n818 10.6151
R1817 B.n818 B.n817 10.6151
R1818 B.n817 B.n814 10.6151
R1819 B.n814 B.n813 10.6151
R1820 B.n813 B.n810 10.6151
R1821 B.n810 B.n809 10.6151
R1822 B.n809 B.n806 10.6151
R1823 B.n806 B.n805 10.6151
R1824 B.n805 B.n802 10.6151
R1825 B.n802 B.n801 10.6151
R1826 B.n801 B.n798 10.6151
R1827 B.n798 B.n797 10.6151
R1828 B.n797 B.n794 10.6151
R1829 B.n794 B.n793 10.6151
R1830 B.n793 B.n790 10.6151
R1831 B.n790 B.n789 10.6151
R1832 B.n789 B.n786 10.6151
R1833 B.n786 B.n785 10.6151
R1834 B.n785 B.n782 10.6151
R1835 B.n782 B.n781 10.6151
R1836 B.n781 B.n778 10.6151
R1837 B.n778 B.n777 10.6151
R1838 B.n777 B.n774 10.6151
R1839 B.n774 B.n773 10.6151
R1840 B.n773 B.n770 10.6151
R1841 B.n770 B.n769 10.6151
R1842 B.n769 B.n766 10.6151
R1843 B.n766 B.n765 10.6151
R1844 B.n765 B.n762 10.6151
R1845 B.n762 B.n761 10.6151
R1846 B.n761 B.n758 10.6151
R1847 B.n758 B.n757 10.6151
R1848 B.n757 B.n754 10.6151
R1849 B.n754 B.n753 10.6151
R1850 B.n753 B.n750 10.6151
R1851 B.n750 B.n749 10.6151
R1852 B.n746 B.n745 10.6151
R1853 B.n745 B.n742 10.6151
R1854 B.n742 B.n741 10.6151
R1855 B.n741 B.n738 10.6151
R1856 B.n738 B.n737 10.6151
R1857 B.n737 B.n734 10.6151
R1858 B.n734 B.n733 10.6151
R1859 B.n733 B.n730 10.6151
R1860 B.n728 B.n725 10.6151
R1861 B.n725 B.n724 10.6151
R1862 B.n724 B.n721 10.6151
R1863 B.n721 B.n720 10.6151
R1864 B.n720 B.n717 10.6151
R1865 B.n717 B.n716 10.6151
R1866 B.n716 B.n713 10.6151
R1867 B.n713 B.n712 10.6151
R1868 B.n712 B.n709 10.6151
R1869 B.n709 B.n708 10.6151
R1870 B.n708 B.n705 10.6151
R1871 B.n705 B.n704 10.6151
R1872 B.n704 B.n701 10.6151
R1873 B.n701 B.n700 10.6151
R1874 B.n700 B.n697 10.6151
R1875 B.n697 B.n696 10.6151
R1876 B.n696 B.n693 10.6151
R1877 B.n693 B.n692 10.6151
R1878 B.n692 B.n689 10.6151
R1879 B.n689 B.n688 10.6151
R1880 B.n688 B.n685 10.6151
R1881 B.n685 B.n684 10.6151
R1882 B.n684 B.n681 10.6151
R1883 B.n681 B.n680 10.6151
R1884 B.n680 B.n677 10.6151
R1885 B.n677 B.n676 10.6151
R1886 B.n676 B.n673 10.6151
R1887 B.n673 B.n672 10.6151
R1888 B.n672 B.n669 10.6151
R1889 B.n669 B.n668 10.6151
R1890 B.n668 B.n665 10.6151
R1891 B.n665 B.n664 10.6151
R1892 B.n664 B.n661 10.6151
R1893 B.n661 B.n660 10.6151
R1894 B.n660 B.n657 10.6151
R1895 B.n657 B.n656 10.6151
R1896 B.n656 B.n653 10.6151
R1897 B.n653 B.n652 10.6151
R1898 B.n652 B.n649 10.6151
R1899 B.n649 B.n648 10.6151
R1900 B.n648 B.n645 10.6151
R1901 B.n645 B.n644 10.6151
R1902 B.n644 B.n641 10.6151
R1903 B.n641 B.n640 10.6151
R1904 B.n640 B.n637 10.6151
R1905 B.n637 B.n636 10.6151
R1906 B.n636 B.n633 10.6151
R1907 B.n633 B.n632 10.6151
R1908 B.n632 B.n629 10.6151
R1909 B.n629 B.n628 10.6151
R1910 B.n628 B.n625 10.6151
R1911 B.n625 B.n624 10.6151
R1912 B.n858 B.n555 10.6151
R1913 B.n859 B.n858 10.6151
R1914 B.n860 B.n859 10.6151
R1915 B.n860 B.n547 10.6151
R1916 B.n870 B.n547 10.6151
R1917 B.n871 B.n870 10.6151
R1918 B.n872 B.n871 10.6151
R1919 B.n872 B.n539 10.6151
R1920 B.n882 B.n539 10.6151
R1921 B.n883 B.n882 10.6151
R1922 B.n884 B.n883 10.6151
R1923 B.n884 B.n531 10.6151
R1924 B.n894 B.n531 10.6151
R1925 B.n895 B.n894 10.6151
R1926 B.n896 B.n895 10.6151
R1927 B.n896 B.n523 10.6151
R1928 B.n906 B.n523 10.6151
R1929 B.n907 B.n906 10.6151
R1930 B.n908 B.n907 10.6151
R1931 B.n908 B.n515 10.6151
R1932 B.n918 B.n515 10.6151
R1933 B.n919 B.n918 10.6151
R1934 B.n920 B.n919 10.6151
R1935 B.n920 B.n507 10.6151
R1936 B.n930 B.n507 10.6151
R1937 B.n931 B.n930 10.6151
R1938 B.n932 B.n931 10.6151
R1939 B.n932 B.n499 10.6151
R1940 B.n942 B.n499 10.6151
R1941 B.n943 B.n942 10.6151
R1942 B.n944 B.n943 10.6151
R1943 B.n944 B.n491 10.6151
R1944 B.n954 B.n491 10.6151
R1945 B.n955 B.n954 10.6151
R1946 B.n956 B.n955 10.6151
R1947 B.n956 B.n482 10.6151
R1948 B.n966 B.n482 10.6151
R1949 B.n967 B.n966 10.6151
R1950 B.n968 B.n967 10.6151
R1951 B.n968 B.n475 10.6151
R1952 B.n978 B.n475 10.6151
R1953 B.n979 B.n978 10.6151
R1954 B.n980 B.n979 10.6151
R1955 B.n980 B.n467 10.6151
R1956 B.n990 B.n467 10.6151
R1957 B.n991 B.n990 10.6151
R1958 B.n992 B.n991 10.6151
R1959 B.n992 B.n458 10.6151
R1960 B.n1002 B.n458 10.6151
R1961 B.n1003 B.n1002 10.6151
R1962 B.n1004 B.n1003 10.6151
R1963 B.n1004 B.n451 10.6151
R1964 B.n1014 B.n451 10.6151
R1965 B.n1015 B.n1014 10.6151
R1966 B.n1016 B.n1015 10.6151
R1967 B.n1016 B.n443 10.6151
R1968 B.n1026 B.n443 10.6151
R1969 B.n1027 B.n1026 10.6151
R1970 B.n1028 B.n1027 10.6151
R1971 B.n1028 B.n435 10.6151
R1972 B.n1038 B.n435 10.6151
R1973 B.n1039 B.n1038 10.6151
R1974 B.n1040 B.n1039 10.6151
R1975 B.n1040 B.n427 10.6151
R1976 B.n1050 B.n427 10.6151
R1977 B.n1051 B.n1050 10.6151
R1978 B.n1053 B.n1051 10.6151
R1979 B.n1053 B.n1052 10.6151
R1980 B.n1052 B.n419 10.6151
R1981 B.n1064 B.n419 10.6151
R1982 B.n1065 B.n1064 10.6151
R1983 B.n1066 B.n1065 10.6151
R1984 B.n1067 B.n1066 10.6151
R1985 B.n1068 B.n1067 10.6151
R1986 B.n1071 B.n1068 10.6151
R1987 B.n1072 B.n1071 10.6151
R1988 B.n1073 B.n1072 10.6151
R1989 B.n1074 B.n1073 10.6151
R1990 B.n1076 B.n1074 10.6151
R1991 B.n1077 B.n1076 10.6151
R1992 B.n1078 B.n1077 10.6151
R1993 B.n1079 B.n1078 10.6151
R1994 B.n1081 B.n1079 10.6151
R1995 B.n1082 B.n1081 10.6151
R1996 B.n1083 B.n1082 10.6151
R1997 B.n1084 B.n1083 10.6151
R1998 B.n1086 B.n1084 10.6151
R1999 B.n1087 B.n1086 10.6151
R2000 B.n1088 B.n1087 10.6151
R2001 B.n1089 B.n1088 10.6151
R2002 B.n1091 B.n1089 10.6151
R2003 B.n1092 B.n1091 10.6151
R2004 B.n1093 B.n1092 10.6151
R2005 B.n1094 B.n1093 10.6151
R2006 B.n1096 B.n1094 10.6151
R2007 B.n1097 B.n1096 10.6151
R2008 B.n1098 B.n1097 10.6151
R2009 B.n1099 B.n1098 10.6151
R2010 B.n1101 B.n1099 10.6151
R2011 B.n1102 B.n1101 10.6151
R2012 B.n1103 B.n1102 10.6151
R2013 B.n1104 B.n1103 10.6151
R2014 B.n1106 B.n1104 10.6151
R2015 B.n1107 B.n1106 10.6151
R2016 B.n1108 B.n1107 10.6151
R2017 B.n1109 B.n1108 10.6151
R2018 B.n1111 B.n1109 10.6151
R2019 B.n1112 B.n1111 10.6151
R2020 B.n1113 B.n1112 10.6151
R2021 B.n1114 B.n1113 10.6151
R2022 B.n1116 B.n1114 10.6151
R2023 B.n1117 B.n1116 10.6151
R2024 B.n1118 B.n1117 10.6151
R2025 B.n1119 B.n1118 10.6151
R2026 B.n1121 B.n1119 10.6151
R2027 B.n1122 B.n1121 10.6151
R2028 B.n1123 B.n1122 10.6151
R2029 B.n1124 B.n1123 10.6151
R2030 B.n1126 B.n1124 10.6151
R2031 B.n1127 B.n1126 10.6151
R2032 B.n1128 B.n1127 10.6151
R2033 B.n1129 B.n1128 10.6151
R2034 B.n1131 B.n1129 10.6151
R2035 B.n1132 B.n1131 10.6151
R2036 B.n1133 B.n1132 10.6151
R2037 B.n1134 B.n1133 10.6151
R2038 B.n1136 B.n1134 10.6151
R2039 B.n1137 B.n1136 10.6151
R2040 B.n1138 B.n1137 10.6151
R2041 B.n1139 B.n1138 10.6151
R2042 B.n1141 B.n1139 10.6151
R2043 B.n1142 B.n1141 10.6151
R2044 B.n1143 B.n1142 10.6151
R2045 B.n1144 B.n1143 10.6151
R2046 B.n1146 B.n1144 10.6151
R2047 B.n1147 B.n1146 10.6151
R2048 B.n1148 B.n1147 10.6151
R2049 B.n1149 B.n1148 10.6151
R2050 B.n1151 B.n1149 10.6151
R2051 B.n1152 B.n1151 10.6151
R2052 B.n1153 B.n1152 10.6151
R2053 B.n1154 B.n1153 10.6151
R2054 B.n1155 B.n1154 10.6151
R2055 B.n1299 B.n1 10.6151
R2056 B.n1299 B.n1298 10.6151
R2057 B.n1298 B.n1297 10.6151
R2058 B.n1297 B.n10 10.6151
R2059 B.n1291 B.n10 10.6151
R2060 B.n1291 B.n1290 10.6151
R2061 B.n1290 B.n1289 10.6151
R2062 B.n1289 B.n18 10.6151
R2063 B.n1283 B.n18 10.6151
R2064 B.n1283 B.n1282 10.6151
R2065 B.n1282 B.n1281 10.6151
R2066 B.n1281 B.n25 10.6151
R2067 B.n1275 B.n25 10.6151
R2068 B.n1275 B.n1274 10.6151
R2069 B.n1274 B.n1273 10.6151
R2070 B.n1273 B.n32 10.6151
R2071 B.n1267 B.n32 10.6151
R2072 B.n1267 B.n1266 10.6151
R2073 B.n1266 B.n1265 10.6151
R2074 B.n1265 B.n39 10.6151
R2075 B.n1259 B.n39 10.6151
R2076 B.n1259 B.n1258 10.6151
R2077 B.n1258 B.n1257 10.6151
R2078 B.n1257 B.n46 10.6151
R2079 B.n1251 B.n46 10.6151
R2080 B.n1251 B.n1250 10.6151
R2081 B.n1250 B.n1249 10.6151
R2082 B.n1249 B.n53 10.6151
R2083 B.n1243 B.n53 10.6151
R2084 B.n1243 B.n1242 10.6151
R2085 B.n1242 B.n1241 10.6151
R2086 B.n1241 B.n60 10.6151
R2087 B.n1235 B.n60 10.6151
R2088 B.n1235 B.n1234 10.6151
R2089 B.n1234 B.n1233 10.6151
R2090 B.n1233 B.n67 10.6151
R2091 B.n1227 B.n67 10.6151
R2092 B.n1227 B.n1226 10.6151
R2093 B.n1226 B.n1225 10.6151
R2094 B.n1225 B.n74 10.6151
R2095 B.n1219 B.n74 10.6151
R2096 B.n1219 B.n1218 10.6151
R2097 B.n1218 B.n1217 10.6151
R2098 B.n1217 B.n81 10.6151
R2099 B.n1211 B.n81 10.6151
R2100 B.n1211 B.n1210 10.6151
R2101 B.n1210 B.n1209 10.6151
R2102 B.n1209 B.n88 10.6151
R2103 B.n1203 B.n88 10.6151
R2104 B.n1203 B.n1202 10.6151
R2105 B.n1202 B.n1201 10.6151
R2106 B.n1201 B.n95 10.6151
R2107 B.n1195 B.n95 10.6151
R2108 B.n1195 B.n1194 10.6151
R2109 B.n1194 B.n1193 10.6151
R2110 B.n1193 B.n102 10.6151
R2111 B.n1187 B.n102 10.6151
R2112 B.n1187 B.n1186 10.6151
R2113 B.n1186 B.n1185 10.6151
R2114 B.n1185 B.n109 10.6151
R2115 B.n1179 B.n109 10.6151
R2116 B.n1179 B.n1178 10.6151
R2117 B.n1178 B.n1177 10.6151
R2118 B.n1177 B.n116 10.6151
R2119 B.n1171 B.n116 10.6151
R2120 B.n1171 B.n1170 10.6151
R2121 B.n1170 B.n1169 10.6151
R2122 B.n1169 B.n123 10.6151
R2123 B.n1163 B.n123 10.6151
R2124 B.n1163 B.n1162 10.6151
R2125 B.n1161 B.n130 10.6151
R2126 B.n196 B.n130 10.6151
R2127 B.n197 B.n196 10.6151
R2128 B.n200 B.n197 10.6151
R2129 B.n201 B.n200 10.6151
R2130 B.n204 B.n201 10.6151
R2131 B.n205 B.n204 10.6151
R2132 B.n208 B.n205 10.6151
R2133 B.n209 B.n208 10.6151
R2134 B.n212 B.n209 10.6151
R2135 B.n213 B.n212 10.6151
R2136 B.n216 B.n213 10.6151
R2137 B.n217 B.n216 10.6151
R2138 B.n220 B.n217 10.6151
R2139 B.n221 B.n220 10.6151
R2140 B.n224 B.n221 10.6151
R2141 B.n225 B.n224 10.6151
R2142 B.n228 B.n225 10.6151
R2143 B.n229 B.n228 10.6151
R2144 B.n232 B.n229 10.6151
R2145 B.n233 B.n232 10.6151
R2146 B.n236 B.n233 10.6151
R2147 B.n237 B.n236 10.6151
R2148 B.n240 B.n237 10.6151
R2149 B.n241 B.n240 10.6151
R2150 B.n244 B.n241 10.6151
R2151 B.n245 B.n244 10.6151
R2152 B.n248 B.n245 10.6151
R2153 B.n249 B.n248 10.6151
R2154 B.n252 B.n249 10.6151
R2155 B.n253 B.n252 10.6151
R2156 B.n256 B.n253 10.6151
R2157 B.n257 B.n256 10.6151
R2158 B.n260 B.n257 10.6151
R2159 B.n261 B.n260 10.6151
R2160 B.n264 B.n261 10.6151
R2161 B.n265 B.n264 10.6151
R2162 B.n268 B.n265 10.6151
R2163 B.n269 B.n268 10.6151
R2164 B.n272 B.n269 10.6151
R2165 B.n273 B.n272 10.6151
R2166 B.n276 B.n273 10.6151
R2167 B.n277 B.n276 10.6151
R2168 B.n280 B.n277 10.6151
R2169 B.n281 B.n280 10.6151
R2170 B.n284 B.n281 10.6151
R2171 B.n285 B.n284 10.6151
R2172 B.n288 B.n285 10.6151
R2173 B.n289 B.n288 10.6151
R2174 B.n292 B.n289 10.6151
R2175 B.n293 B.n292 10.6151
R2176 B.n296 B.n293 10.6151
R2177 B.n301 B.n298 10.6151
R2178 B.n302 B.n301 10.6151
R2179 B.n305 B.n302 10.6151
R2180 B.n306 B.n305 10.6151
R2181 B.n309 B.n306 10.6151
R2182 B.n310 B.n309 10.6151
R2183 B.n313 B.n310 10.6151
R2184 B.n314 B.n313 10.6151
R2185 B.n318 B.n317 10.6151
R2186 B.n321 B.n318 10.6151
R2187 B.n322 B.n321 10.6151
R2188 B.n325 B.n322 10.6151
R2189 B.n326 B.n325 10.6151
R2190 B.n329 B.n326 10.6151
R2191 B.n330 B.n329 10.6151
R2192 B.n333 B.n330 10.6151
R2193 B.n334 B.n333 10.6151
R2194 B.n337 B.n334 10.6151
R2195 B.n338 B.n337 10.6151
R2196 B.n341 B.n338 10.6151
R2197 B.n342 B.n341 10.6151
R2198 B.n345 B.n342 10.6151
R2199 B.n346 B.n345 10.6151
R2200 B.n349 B.n346 10.6151
R2201 B.n350 B.n349 10.6151
R2202 B.n353 B.n350 10.6151
R2203 B.n354 B.n353 10.6151
R2204 B.n357 B.n354 10.6151
R2205 B.n358 B.n357 10.6151
R2206 B.n361 B.n358 10.6151
R2207 B.n362 B.n361 10.6151
R2208 B.n365 B.n362 10.6151
R2209 B.n366 B.n365 10.6151
R2210 B.n369 B.n366 10.6151
R2211 B.n370 B.n369 10.6151
R2212 B.n373 B.n370 10.6151
R2213 B.n374 B.n373 10.6151
R2214 B.n377 B.n374 10.6151
R2215 B.n378 B.n377 10.6151
R2216 B.n381 B.n378 10.6151
R2217 B.n382 B.n381 10.6151
R2218 B.n385 B.n382 10.6151
R2219 B.n386 B.n385 10.6151
R2220 B.n389 B.n386 10.6151
R2221 B.n390 B.n389 10.6151
R2222 B.n393 B.n390 10.6151
R2223 B.n394 B.n393 10.6151
R2224 B.n397 B.n394 10.6151
R2225 B.n398 B.n397 10.6151
R2226 B.n401 B.n398 10.6151
R2227 B.n402 B.n401 10.6151
R2228 B.n405 B.n402 10.6151
R2229 B.n406 B.n405 10.6151
R2230 B.n409 B.n406 10.6151
R2231 B.n410 B.n409 10.6151
R2232 B.n413 B.n410 10.6151
R2233 B.n414 B.n413 10.6151
R2234 B.n417 B.n414 10.6151
R2235 B.n418 B.n417 10.6151
R2236 B.n1156 B.n418 10.6151
R2237 B.n1307 B.n0 8.11757
R2238 B.n1307 B.n1 8.11757
R2239 B.n485 B.t3 7.33908
R2240 B.t4 B.n1238 7.33908
R2241 B.n746 B.n620 6.5566
R2242 B.n730 B.n729 6.5566
R2243 B.n298 B.n297 6.5566
R2244 B.n314 B.n192 6.5566
R2245 B.n1006 B.t1 4.19397
R2246 B.n1263 B.t7 4.19397
R2247 B.n749 B.n620 4.05904
R2248 B.n729 B.n728 4.05904
R2249 B.n297 B.n296 4.05904
R2250 B.n317 B.n192 4.05904
R2251 VN.n75 VN.n39 161.3
R2252 VN.n74 VN.n73 161.3
R2253 VN.n72 VN.n40 161.3
R2254 VN.n71 VN.n70 161.3
R2255 VN.n69 VN.n41 161.3
R2256 VN.n68 VN.n67 161.3
R2257 VN.n66 VN.n42 161.3
R2258 VN.n65 VN.n64 161.3
R2259 VN.n62 VN.n43 161.3
R2260 VN.n61 VN.n60 161.3
R2261 VN.n59 VN.n44 161.3
R2262 VN.n58 VN.n57 161.3
R2263 VN.n56 VN.n45 161.3
R2264 VN.n55 VN.n54 161.3
R2265 VN.n53 VN.n46 161.3
R2266 VN.n52 VN.n51 161.3
R2267 VN.n50 VN.n47 161.3
R2268 VN.n36 VN.n0 161.3
R2269 VN.n35 VN.n34 161.3
R2270 VN.n33 VN.n1 161.3
R2271 VN.n32 VN.n31 161.3
R2272 VN.n30 VN.n2 161.3
R2273 VN.n29 VN.n28 161.3
R2274 VN.n27 VN.n3 161.3
R2275 VN.n26 VN.n25 161.3
R2276 VN.n23 VN.n4 161.3
R2277 VN.n22 VN.n21 161.3
R2278 VN.n20 VN.n5 161.3
R2279 VN.n19 VN.n18 161.3
R2280 VN.n17 VN.n6 161.3
R2281 VN.n16 VN.n15 161.3
R2282 VN.n14 VN.n7 161.3
R2283 VN.n13 VN.n12 161.3
R2284 VN.n11 VN.n8 161.3
R2285 VN.n9 VN.t7 127.237
R2286 VN.n48 VN.t4 127.237
R2287 VN.n10 VN.t0 95.1289
R2288 VN.n24 VN.t2 95.1289
R2289 VN.n37 VN.t5 95.1289
R2290 VN.n49 VN.t3 95.1289
R2291 VN.n63 VN.t6 95.1289
R2292 VN.n76 VN.t1 95.1289
R2293 VN.n10 VN.n9 67.569
R2294 VN.n49 VN.n48 67.569
R2295 VN VN.n77 60.4814
R2296 VN.n38 VN.n37 59.4275
R2297 VN.n77 VN.n76 59.4275
R2298 VN.n31 VN.n30 56.5193
R2299 VN.n70 VN.n69 56.5193
R2300 VN.n17 VN.n16 40.4934
R2301 VN.n18 VN.n17 40.4934
R2302 VN.n56 VN.n55 40.4934
R2303 VN.n57 VN.n56 40.4934
R2304 VN.n12 VN.n11 24.4675
R2305 VN.n12 VN.n7 24.4675
R2306 VN.n16 VN.n7 24.4675
R2307 VN.n18 VN.n5 24.4675
R2308 VN.n22 VN.n5 24.4675
R2309 VN.n23 VN.n22 24.4675
R2310 VN.n25 VN.n3 24.4675
R2311 VN.n29 VN.n3 24.4675
R2312 VN.n30 VN.n29 24.4675
R2313 VN.n31 VN.n1 24.4675
R2314 VN.n35 VN.n1 24.4675
R2315 VN.n36 VN.n35 24.4675
R2316 VN.n55 VN.n46 24.4675
R2317 VN.n51 VN.n46 24.4675
R2318 VN.n51 VN.n50 24.4675
R2319 VN.n69 VN.n68 24.4675
R2320 VN.n68 VN.n42 24.4675
R2321 VN.n64 VN.n42 24.4675
R2322 VN.n62 VN.n61 24.4675
R2323 VN.n61 VN.n44 24.4675
R2324 VN.n57 VN.n44 24.4675
R2325 VN.n75 VN.n74 24.4675
R2326 VN.n74 VN.n40 24.4675
R2327 VN.n70 VN.n40 24.4675
R2328 VN.n37 VN.n36 22.7548
R2329 VN.n76 VN.n75 22.7548
R2330 VN.n25 VN.n24 16.8827
R2331 VN.n64 VN.n63 16.8827
R2332 VN.n11 VN.n10 7.58527
R2333 VN.n24 VN.n23 7.58527
R2334 VN.n50 VN.n49 7.58527
R2335 VN.n63 VN.n62 7.58527
R2336 VN.n48 VN.n47 2.59903
R2337 VN.n9 VN.n8 2.59903
R2338 VN.n77 VN.n39 0.417535
R2339 VN.n38 VN.n0 0.417535
R2340 VN VN.n38 0.394291
R2341 VN.n73 VN.n39 0.189894
R2342 VN.n73 VN.n72 0.189894
R2343 VN.n72 VN.n71 0.189894
R2344 VN.n71 VN.n41 0.189894
R2345 VN.n67 VN.n41 0.189894
R2346 VN.n67 VN.n66 0.189894
R2347 VN.n66 VN.n65 0.189894
R2348 VN.n65 VN.n43 0.189894
R2349 VN.n60 VN.n43 0.189894
R2350 VN.n60 VN.n59 0.189894
R2351 VN.n59 VN.n58 0.189894
R2352 VN.n58 VN.n45 0.189894
R2353 VN.n54 VN.n45 0.189894
R2354 VN.n54 VN.n53 0.189894
R2355 VN.n53 VN.n52 0.189894
R2356 VN.n52 VN.n47 0.189894
R2357 VN.n13 VN.n8 0.189894
R2358 VN.n14 VN.n13 0.189894
R2359 VN.n15 VN.n14 0.189894
R2360 VN.n15 VN.n6 0.189894
R2361 VN.n19 VN.n6 0.189894
R2362 VN.n20 VN.n19 0.189894
R2363 VN.n21 VN.n20 0.189894
R2364 VN.n21 VN.n4 0.189894
R2365 VN.n26 VN.n4 0.189894
R2366 VN.n27 VN.n26 0.189894
R2367 VN.n28 VN.n27 0.189894
R2368 VN.n28 VN.n2 0.189894
R2369 VN.n32 VN.n2 0.189894
R2370 VN.n33 VN.n32 0.189894
R2371 VN.n34 VN.n33 0.189894
R2372 VN.n34 VN.n0 0.189894
R2373 VTAIL.n11 VTAIL.t5 45.1958
R2374 VTAIL.n10 VTAIL.t10 45.1958
R2375 VTAIL.n7 VTAIL.t12 45.1958
R2376 VTAIL.n15 VTAIL.t14 45.1957
R2377 VTAIL.n2 VTAIL.t15 45.1957
R2378 VTAIL.n3 VTAIL.t1 45.1957
R2379 VTAIL.n6 VTAIL.t4 45.1957
R2380 VTAIL.n14 VTAIL.t0 45.1957
R2381 VTAIL.n13 VTAIL.n12 43.9356
R2382 VTAIL.n9 VTAIL.n8 43.9356
R2383 VTAIL.n1 VTAIL.n0 43.9353
R2384 VTAIL.n5 VTAIL.n4 43.9353
R2385 VTAIL.n15 VTAIL.n14 29.6255
R2386 VTAIL.n7 VTAIL.n6 29.6255
R2387 VTAIL.n9 VTAIL.n7 3.71602
R2388 VTAIL.n10 VTAIL.n9 3.71602
R2389 VTAIL.n13 VTAIL.n11 3.71602
R2390 VTAIL.n14 VTAIL.n13 3.71602
R2391 VTAIL.n6 VTAIL.n5 3.71602
R2392 VTAIL.n5 VTAIL.n3 3.71602
R2393 VTAIL.n2 VTAIL.n1 3.71602
R2394 VTAIL VTAIL.n15 3.65783
R2395 VTAIL.n0 VTAIL.t9 1.26084
R2396 VTAIL.n0 VTAIL.t13 1.26084
R2397 VTAIL.n4 VTAIL.t2 1.26084
R2398 VTAIL.n4 VTAIL.t7 1.26084
R2399 VTAIL.n12 VTAIL.t6 1.26084
R2400 VTAIL.n12 VTAIL.t3 1.26084
R2401 VTAIL.n8 VTAIL.t8 1.26084
R2402 VTAIL.n8 VTAIL.t11 1.26084
R2403 VTAIL.n11 VTAIL.n10 0.470328
R2404 VTAIL.n3 VTAIL.n2 0.470328
R2405 VTAIL VTAIL.n1 0.0586897
R2406 VDD2.n2 VDD2.n1 62.4165
R2407 VDD2.n2 VDD2.n0 62.4165
R2408 VDD2 VDD2.n5 62.4137
R2409 VDD2.n4 VDD2.n3 60.6144
R2410 VDD2.n4 VDD2.n2 53.9782
R2411 VDD2 VDD2.n4 1.91645
R2412 VDD2.n5 VDD2.t4 1.26084
R2413 VDD2.n5 VDD2.t3 1.26084
R2414 VDD2.n3 VDD2.t6 1.26084
R2415 VDD2.n3 VDD2.t1 1.26084
R2416 VDD2.n1 VDD2.t5 1.26084
R2417 VDD2.n1 VDD2.t2 1.26084
R2418 VDD2.n0 VDD2.t0 1.26084
R2419 VDD2.n0 VDD2.t7 1.26084
R2420 VP.n24 VP.n21 161.3
R2421 VP.n26 VP.n25 161.3
R2422 VP.n27 VP.n20 161.3
R2423 VP.n29 VP.n28 161.3
R2424 VP.n30 VP.n19 161.3
R2425 VP.n32 VP.n31 161.3
R2426 VP.n33 VP.n18 161.3
R2427 VP.n35 VP.n34 161.3
R2428 VP.n36 VP.n17 161.3
R2429 VP.n39 VP.n38 161.3
R2430 VP.n40 VP.n16 161.3
R2431 VP.n42 VP.n41 161.3
R2432 VP.n43 VP.n15 161.3
R2433 VP.n45 VP.n44 161.3
R2434 VP.n46 VP.n14 161.3
R2435 VP.n48 VP.n47 161.3
R2436 VP.n49 VP.n13 161.3
R2437 VP.n92 VP.n0 161.3
R2438 VP.n91 VP.n90 161.3
R2439 VP.n89 VP.n1 161.3
R2440 VP.n88 VP.n87 161.3
R2441 VP.n86 VP.n2 161.3
R2442 VP.n85 VP.n84 161.3
R2443 VP.n83 VP.n3 161.3
R2444 VP.n82 VP.n81 161.3
R2445 VP.n79 VP.n4 161.3
R2446 VP.n78 VP.n77 161.3
R2447 VP.n76 VP.n5 161.3
R2448 VP.n75 VP.n74 161.3
R2449 VP.n73 VP.n6 161.3
R2450 VP.n72 VP.n71 161.3
R2451 VP.n70 VP.n7 161.3
R2452 VP.n69 VP.n68 161.3
R2453 VP.n67 VP.n8 161.3
R2454 VP.n65 VP.n64 161.3
R2455 VP.n63 VP.n9 161.3
R2456 VP.n62 VP.n61 161.3
R2457 VP.n60 VP.n10 161.3
R2458 VP.n59 VP.n58 161.3
R2459 VP.n57 VP.n11 161.3
R2460 VP.n56 VP.n55 161.3
R2461 VP.n54 VP.n12 161.3
R2462 VP.n22 VP.t2 127.237
R2463 VP.n53 VP.t7 95.1289
R2464 VP.n66 VP.t3 95.1289
R2465 VP.n80 VP.t1 95.1289
R2466 VP.n93 VP.t6 95.1289
R2467 VP.n50 VP.t4 95.1289
R2468 VP.n37 VP.t0 95.1289
R2469 VP.n23 VP.t5 95.1289
R2470 VP.n23 VP.n22 67.569
R2471 VP.n52 VP.n51 60.4434
R2472 VP.n53 VP.n52 59.4275
R2473 VP.n94 VP.n93 59.4275
R2474 VP.n51 VP.n50 59.4275
R2475 VP.n60 VP.n59 56.5193
R2476 VP.n87 VP.n86 56.5193
R2477 VP.n44 VP.n43 56.5193
R2478 VP.n73 VP.n72 40.4934
R2479 VP.n74 VP.n73 40.4934
R2480 VP.n31 VP.n30 40.4934
R2481 VP.n30 VP.n29 40.4934
R2482 VP.n55 VP.n54 24.4675
R2483 VP.n55 VP.n11 24.4675
R2484 VP.n59 VP.n11 24.4675
R2485 VP.n61 VP.n60 24.4675
R2486 VP.n61 VP.n9 24.4675
R2487 VP.n65 VP.n9 24.4675
R2488 VP.n68 VP.n67 24.4675
R2489 VP.n68 VP.n7 24.4675
R2490 VP.n72 VP.n7 24.4675
R2491 VP.n74 VP.n5 24.4675
R2492 VP.n78 VP.n5 24.4675
R2493 VP.n79 VP.n78 24.4675
R2494 VP.n81 VP.n3 24.4675
R2495 VP.n85 VP.n3 24.4675
R2496 VP.n86 VP.n85 24.4675
R2497 VP.n87 VP.n1 24.4675
R2498 VP.n91 VP.n1 24.4675
R2499 VP.n92 VP.n91 24.4675
R2500 VP.n44 VP.n14 24.4675
R2501 VP.n48 VP.n14 24.4675
R2502 VP.n49 VP.n48 24.4675
R2503 VP.n31 VP.n18 24.4675
R2504 VP.n35 VP.n18 24.4675
R2505 VP.n36 VP.n35 24.4675
R2506 VP.n38 VP.n16 24.4675
R2507 VP.n42 VP.n16 24.4675
R2508 VP.n43 VP.n42 24.4675
R2509 VP.n25 VP.n24 24.4675
R2510 VP.n25 VP.n20 24.4675
R2511 VP.n29 VP.n20 24.4675
R2512 VP.n54 VP.n53 22.7548
R2513 VP.n93 VP.n92 22.7548
R2514 VP.n50 VP.n49 22.7548
R2515 VP.n66 VP.n65 16.8827
R2516 VP.n81 VP.n80 16.8827
R2517 VP.n38 VP.n37 16.8827
R2518 VP.n67 VP.n66 7.58527
R2519 VP.n80 VP.n79 7.58527
R2520 VP.n37 VP.n36 7.58527
R2521 VP.n24 VP.n23 7.58527
R2522 VP.n22 VP.n21 2.599
R2523 VP.n51 VP.n13 0.417535
R2524 VP.n52 VP.n12 0.417535
R2525 VP.n94 VP.n0 0.417535
R2526 VP VP.n94 0.394291
R2527 VP.n26 VP.n21 0.189894
R2528 VP.n27 VP.n26 0.189894
R2529 VP.n28 VP.n27 0.189894
R2530 VP.n28 VP.n19 0.189894
R2531 VP.n32 VP.n19 0.189894
R2532 VP.n33 VP.n32 0.189894
R2533 VP.n34 VP.n33 0.189894
R2534 VP.n34 VP.n17 0.189894
R2535 VP.n39 VP.n17 0.189894
R2536 VP.n40 VP.n39 0.189894
R2537 VP.n41 VP.n40 0.189894
R2538 VP.n41 VP.n15 0.189894
R2539 VP.n45 VP.n15 0.189894
R2540 VP.n46 VP.n45 0.189894
R2541 VP.n47 VP.n46 0.189894
R2542 VP.n47 VP.n13 0.189894
R2543 VP.n56 VP.n12 0.189894
R2544 VP.n57 VP.n56 0.189894
R2545 VP.n58 VP.n57 0.189894
R2546 VP.n58 VP.n10 0.189894
R2547 VP.n62 VP.n10 0.189894
R2548 VP.n63 VP.n62 0.189894
R2549 VP.n64 VP.n63 0.189894
R2550 VP.n64 VP.n8 0.189894
R2551 VP.n69 VP.n8 0.189894
R2552 VP.n70 VP.n69 0.189894
R2553 VP.n71 VP.n70 0.189894
R2554 VP.n71 VP.n6 0.189894
R2555 VP.n75 VP.n6 0.189894
R2556 VP.n76 VP.n75 0.189894
R2557 VP.n77 VP.n76 0.189894
R2558 VP.n77 VP.n4 0.189894
R2559 VP.n82 VP.n4 0.189894
R2560 VP.n83 VP.n82 0.189894
R2561 VP.n84 VP.n83 0.189894
R2562 VP.n84 VP.n2 0.189894
R2563 VP.n88 VP.n2 0.189894
R2564 VP.n89 VP.n88 0.189894
R2565 VP.n90 VP.n89 0.189894
R2566 VP.n90 VP.n0 0.189894
R2567 VDD1 VDD1.n0 62.5303
R2568 VDD1.n3 VDD1.n2 62.4165
R2569 VDD1.n3 VDD1.n1 62.4165
R2570 VDD1.n5 VDD1.n4 60.6142
R2571 VDD1.n5 VDD1.n3 54.5612
R2572 VDD1 VDD1.n5 1.80007
R2573 VDD1.n4 VDD1.t7 1.26084
R2574 VDD1.n4 VDD1.t3 1.26084
R2575 VDD1.n0 VDD1.t5 1.26084
R2576 VDD1.n0 VDD1.t2 1.26084
R2577 VDD1.n2 VDD1.t6 1.26084
R2578 VDD1.n2 VDD1.t1 1.26084
R2579 VDD1.n1 VDD1.t0 1.26084
R2580 VDD1.n1 VDD1.t4 1.26084
C0 VDD2 VP 0.666672f
C1 VN VTAIL 12.7323f
C2 VDD1 VP 12.5542f
C3 VDD2 VN 12.044f
C4 VDD2 VTAIL 9.789481f
C5 VDD1 VN 0.154377f
C6 VDD1 VTAIL 9.725809f
C7 VDD1 VDD2 2.49528f
C8 VN VP 10.0387f
C9 VTAIL VP 12.7464f
C10 VDD2 B 7.05632f
C11 VDD1 B 7.643719f
C12 VTAIL B 13.650852f
C13 VN B 21.12767f
C14 VP B 19.773958f
C15 VDD1.t5 B 0.337069f
C16 VDD1.t2 B 0.337069f
C17 VDD1.n0 B 3.0751f
C18 VDD1.t0 B 0.337069f
C19 VDD1.t4 B 0.337069f
C20 VDD1.n1 B 3.07354f
C21 VDD1.t6 B 0.337069f
C22 VDD1.t1 B 0.337069f
C23 VDD1.n2 B 3.07354f
C24 VDD1.n3 B 4.73649f
C25 VDD1.t7 B 0.337069f
C26 VDD1.t3 B 0.337069f
C27 VDD1.n4 B 3.05281f
C28 VDD1.n5 B 4.06206f
C29 VP.n0 B 0.030652f
C30 VP.t6 B 2.79482f
C31 VP.n1 B 0.030371f
C32 VP.n2 B 0.016296f
C33 VP.n3 B 0.030371f
C34 VP.n4 B 0.016296f
C35 VP.t1 B 2.79482f
C36 VP.n5 B 0.030371f
C37 VP.n6 B 0.016296f
C38 VP.n7 B 0.030371f
C39 VP.n8 B 0.016296f
C40 VP.t3 B 2.79482f
C41 VP.n9 B 0.030371f
C42 VP.n10 B 0.016296f
C43 VP.n11 B 0.030371f
C44 VP.n12 B 0.030652f
C45 VP.t7 B 2.79482f
C46 VP.n13 B 0.030652f
C47 VP.t4 B 2.79482f
C48 VP.n14 B 0.030371f
C49 VP.n15 B 0.016296f
C50 VP.n16 B 0.030371f
C51 VP.n17 B 0.016296f
C52 VP.t0 B 2.79482f
C53 VP.n18 B 0.030371f
C54 VP.n19 B 0.016296f
C55 VP.n20 B 0.030371f
C56 VP.n21 B 0.215723f
C57 VP.t5 B 2.79482f
C58 VP.t2 B 3.07182f
C59 VP.n22 B 0.977146f
C60 VP.n23 B 1.02362f
C61 VP.n24 B 0.020024f
C62 VP.n25 B 0.030371f
C63 VP.n26 B 0.016296f
C64 VP.n27 B 0.016296f
C65 VP.n28 B 0.016296f
C66 VP.n29 B 0.032387f
C67 VP.n30 B 0.013173f
C68 VP.n31 B 0.032387f
C69 VP.n32 B 0.016296f
C70 VP.n33 B 0.016296f
C71 VP.n34 B 0.016296f
C72 VP.n35 B 0.030371f
C73 VP.n36 B 0.020024f
C74 VP.n37 B 0.966795f
C75 VP.n38 B 0.025722f
C76 VP.n39 B 0.016296f
C77 VP.n40 B 0.016296f
C78 VP.n41 B 0.016296f
C79 VP.n42 B 0.030371f
C80 VP.n43 B 0.026513f
C81 VP.n44 B 0.021064f
C82 VP.n45 B 0.016296f
C83 VP.n46 B 0.016296f
C84 VP.n47 B 0.016296f
C85 VP.n48 B 0.030371f
C86 VP.n49 B 0.02932f
C87 VP.n50 B 1.04138f
C88 VP.n51 B 1.22554f
C89 VP.n52 B 1.23523f
C90 VP.n53 B 1.04138f
C91 VP.n54 B 0.02932f
C92 VP.n55 B 0.030371f
C93 VP.n56 B 0.016296f
C94 VP.n57 B 0.016296f
C95 VP.n58 B 0.016296f
C96 VP.n59 B 0.021064f
C97 VP.n60 B 0.026513f
C98 VP.n61 B 0.030371f
C99 VP.n62 B 0.016296f
C100 VP.n63 B 0.016296f
C101 VP.n64 B 0.016296f
C102 VP.n65 B 0.025722f
C103 VP.n66 B 0.966795f
C104 VP.n67 B 0.020024f
C105 VP.n68 B 0.030371f
C106 VP.n69 B 0.016296f
C107 VP.n70 B 0.016296f
C108 VP.n71 B 0.016296f
C109 VP.n72 B 0.032387f
C110 VP.n73 B 0.013173f
C111 VP.n74 B 0.032387f
C112 VP.n75 B 0.016296f
C113 VP.n76 B 0.016296f
C114 VP.n77 B 0.016296f
C115 VP.n78 B 0.030371f
C116 VP.n79 B 0.020024f
C117 VP.n80 B 0.966795f
C118 VP.n81 B 0.025722f
C119 VP.n82 B 0.016296f
C120 VP.n83 B 0.016296f
C121 VP.n84 B 0.016296f
C122 VP.n85 B 0.030371f
C123 VP.n86 B 0.026513f
C124 VP.n87 B 0.021064f
C125 VP.n88 B 0.016296f
C126 VP.n89 B 0.016296f
C127 VP.n90 B 0.016296f
C128 VP.n91 B 0.030371f
C129 VP.n92 B 0.02932f
C130 VP.n93 B 1.04138f
C131 VP.n94 B 0.049631f
C132 VDD2.t0 B 0.331614f
C133 VDD2.t7 B 0.331614f
C134 VDD2.n0 B 3.0238f
C135 VDD2.t5 B 0.331614f
C136 VDD2.t2 B 0.331614f
C137 VDD2.n1 B 3.0238f
C138 VDD2.n2 B 4.60507f
C139 VDD2.t6 B 0.331614f
C140 VDD2.t1 B 0.331614f
C141 VDD2.n3 B 3.00341f
C142 VDD2.n4 B 3.96243f
C143 VDD2.t4 B 0.331614f
C144 VDD2.t3 B 0.331614f
C145 VDD2.n5 B 3.02374f
C146 VTAIL.t9 B 0.244876f
C147 VTAIL.t13 B 0.244876f
C148 VTAIL.n0 B 2.15761f
C149 VTAIL.n1 B 0.435654f
C150 VTAIL.t15 B 2.75348f
C151 VTAIL.n2 B 0.533788f
C152 VTAIL.t1 B 2.75348f
C153 VTAIL.n3 B 0.533788f
C154 VTAIL.t2 B 0.244876f
C155 VTAIL.t7 B 0.244876f
C156 VTAIL.n4 B 2.15761f
C157 VTAIL.n5 B 0.668107f
C158 VTAIL.t4 B 2.75348f
C159 VTAIL.n6 B 1.86879f
C160 VTAIL.t12 B 2.7535f
C161 VTAIL.n7 B 1.86878f
C162 VTAIL.t8 B 0.244876f
C163 VTAIL.t11 B 0.244876f
C164 VTAIL.n8 B 2.15761f
C165 VTAIL.n9 B 0.668104f
C166 VTAIL.t10 B 2.7535f
C167 VTAIL.n10 B 0.53377f
C168 VTAIL.t5 B 2.7535f
C169 VTAIL.n11 B 0.53377f
C170 VTAIL.t6 B 0.244876f
C171 VTAIL.t3 B 0.244876f
C172 VTAIL.n12 B 2.15761f
C173 VTAIL.n13 B 0.668104f
C174 VTAIL.t0 B 2.75348f
C175 VTAIL.n14 B 1.86879f
C176 VTAIL.t14 B 2.75348f
C177 VTAIL.n15 B 1.8651f
C178 VN.n0 B 0.030111f
C179 VN.t5 B 2.74554f
C180 VN.n1 B 0.029835f
C181 VN.n2 B 0.016008f
C182 VN.n3 B 0.029835f
C183 VN.n4 B 0.016008f
C184 VN.t2 B 2.74554f
C185 VN.n5 B 0.029835f
C186 VN.n6 B 0.016008f
C187 VN.n7 B 0.029835f
C188 VN.n8 B 0.211918f
C189 VN.t0 B 2.74554f
C190 VN.t7 B 3.01765f
C191 VN.n9 B 0.959911f
C192 VN.n10 B 1.00557f
C193 VN.n11 B 0.019671f
C194 VN.n12 B 0.029835f
C195 VN.n13 B 0.016008f
C196 VN.n14 B 0.016008f
C197 VN.n15 B 0.016008f
C198 VN.n16 B 0.031816f
C199 VN.n17 B 0.012941f
C200 VN.n18 B 0.031816f
C201 VN.n19 B 0.016008f
C202 VN.n20 B 0.016008f
C203 VN.n21 B 0.016008f
C204 VN.n22 B 0.029835f
C205 VN.n23 B 0.019671f
C206 VN.n24 B 0.949746f
C207 VN.n25 B 0.025268f
C208 VN.n26 B 0.016008f
C209 VN.n27 B 0.016008f
C210 VN.n28 B 0.016008f
C211 VN.n29 B 0.029835f
C212 VN.n30 B 0.026046f
C213 VN.n31 B 0.020692f
C214 VN.n32 B 0.016008f
C215 VN.n33 B 0.016008f
C216 VN.n34 B 0.016008f
C217 VN.n35 B 0.029835f
C218 VN.n36 B 0.028803f
C219 VN.n37 B 1.02302f
C220 VN.n38 B 0.048756f
C221 VN.n39 B 0.030111f
C222 VN.t1 B 2.74554f
C223 VN.n40 B 0.029835f
C224 VN.n41 B 0.016008f
C225 VN.n42 B 0.029835f
C226 VN.n43 B 0.016008f
C227 VN.t6 B 2.74554f
C228 VN.n44 B 0.029835f
C229 VN.n45 B 0.016008f
C230 VN.n46 B 0.029835f
C231 VN.n47 B 0.211918f
C232 VN.t3 B 2.74554f
C233 VN.t4 B 3.01765f
C234 VN.n48 B 0.959911f
C235 VN.n49 B 1.00557f
C236 VN.n50 B 0.019671f
C237 VN.n51 B 0.029835f
C238 VN.n52 B 0.016008f
C239 VN.n53 B 0.016008f
C240 VN.n54 B 0.016008f
C241 VN.n55 B 0.031816f
C242 VN.n56 B 0.012941f
C243 VN.n57 B 0.031816f
C244 VN.n58 B 0.016008f
C245 VN.n59 B 0.016008f
C246 VN.n60 B 0.016008f
C247 VN.n61 B 0.029835f
C248 VN.n62 B 0.019671f
C249 VN.n63 B 0.949746f
C250 VN.n64 B 0.025268f
C251 VN.n65 B 0.016008f
C252 VN.n66 B 0.016008f
C253 VN.n67 B 0.016008f
C254 VN.n68 B 0.029835f
C255 VN.n69 B 0.026046f
C256 VN.n70 B 0.020692f
C257 VN.n71 B 0.016008f
C258 VN.n72 B 0.016008f
C259 VN.n73 B 0.016008f
C260 VN.n74 B 0.029835f
C261 VN.n75 B 0.028803f
C262 VN.n76 B 1.02302f
C263 VN.n77 B 1.20756f
.ends

