* NGSPICE file created from diff_pair_sample_1063.ext - technology: sky130A

.subckt diff_pair_sample_1063 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t19 VP.t0 VDD1.t9 w_n2122_n3970# sky130_fd_pr__pfet_01v8 ad=2.47665 pd=15.34 as=2.47665 ps=15.34 w=15.01 l=0.63
X1 VDD2.t9 VN.t0 VTAIL.t4 w_n2122_n3970# sky130_fd_pr__pfet_01v8 ad=2.47665 pd=15.34 as=5.8539 ps=30.8 w=15.01 l=0.63
X2 B.t11 B.t9 B.t10 w_n2122_n3970# sky130_fd_pr__pfet_01v8 ad=5.8539 pd=30.8 as=0 ps=0 w=15.01 l=0.63
X3 B.t8 B.t6 B.t7 w_n2122_n3970# sky130_fd_pr__pfet_01v8 ad=5.8539 pd=30.8 as=0 ps=0 w=15.01 l=0.63
X4 VDD2.t8 VN.t1 VTAIL.t3 w_n2122_n3970# sky130_fd_pr__pfet_01v8 ad=2.47665 pd=15.34 as=2.47665 ps=15.34 w=15.01 l=0.63
X5 VDD1.t6 VP.t1 VTAIL.t18 w_n2122_n3970# sky130_fd_pr__pfet_01v8 ad=5.8539 pd=30.8 as=2.47665 ps=15.34 w=15.01 l=0.63
X6 B.t5 B.t3 B.t4 w_n2122_n3970# sky130_fd_pr__pfet_01v8 ad=5.8539 pd=30.8 as=0 ps=0 w=15.01 l=0.63
X7 VDD2.t7 VN.t2 VTAIL.t0 w_n2122_n3970# sky130_fd_pr__pfet_01v8 ad=2.47665 pd=15.34 as=5.8539 ps=30.8 w=15.01 l=0.63
X8 VTAIL.t7 VN.t3 VDD2.t6 w_n2122_n3970# sky130_fd_pr__pfet_01v8 ad=2.47665 pd=15.34 as=2.47665 ps=15.34 w=15.01 l=0.63
X9 VDD2.t5 VN.t4 VTAIL.t2 w_n2122_n3970# sky130_fd_pr__pfet_01v8 ad=2.47665 pd=15.34 as=2.47665 ps=15.34 w=15.01 l=0.63
X10 VDD2.t4 VN.t5 VTAIL.t5 w_n2122_n3970# sky130_fd_pr__pfet_01v8 ad=5.8539 pd=30.8 as=2.47665 ps=15.34 w=15.01 l=0.63
X11 B.t2 B.t0 B.t1 w_n2122_n3970# sky130_fd_pr__pfet_01v8 ad=5.8539 pd=30.8 as=0 ps=0 w=15.01 l=0.63
X12 VDD2.t3 VN.t6 VTAIL.t8 w_n2122_n3970# sky130_fd_pr__pfet_01v8 ad=5.8539 pd=30.8 as=2.47665 ps=15.34 w=15.01 l=0.63
X13 VTAIL.t1 VN.t7 VDD2.t2 w_n2122_n3970# sky130_fd_pr__pfet_01v8 ad=2.47665 pd=15.34 as=2.47665 ps=15.34 w=15.01 l=0.63
X14 VDD1.t2 VP.t2 VTAIL.t17 w_n2122_n3970# sky130_fd_pr__pfet_01v8 ad=2.47665 pd=15.34 as=2.47665 ps=15.34 w=15.01 l=0.63
X15 VDD1.t8 VP.t3 VTAIL.t16 w_n2122_n3970# sky130_fd_pr__pfet_01v8 ad=2.47665 pd=15.34 as=5.8539 ps=30.8 w=15.01 l=0.63
X16 VDD1.t5 VP.t4 VTAIL.t15 w_n2122_n3970# sky130_fd_pr__pfet_01v8 ad=2.47665 pd=15.34 as=5.8539 ps=30.8 w=15.01 l=0.63
X17 VTAIL.t14 VP.t5 VDD1.t7 w_n2122_n3970# sky130_fd_pr__pfet_01v8 ad=2.47665 pd=15.34 as=2.47665 ps=15.34 w=15.01 l=0.63
X18 VDD1.t3 VP.t6 VTAIL.t13 w_n2122_n3970# sky130_fd_pr__pfet_01v8 ad=2.47665 pd=15.34 as=2.47665 ps=15.34 w=15.01 l=0.63
X19 VDD1.t0 VP.t7 VTAIL.t12 w_n2122_n3970# sky130_fd_pr__pfet_01v8 ad=5.8539 pd=30.8 as=2.47665 ps=15.34 w=15.01 l=0.63
X20 VTAIL.t11 VP.t8 VDD1.t1 w_n2122_n3970# sky130_fd_pr__pfet_01v8 ad=2.47665 pd=15.34 as=2.47665 ps=15.34 w=15.01 l=0.63
X21 VTAIL.t6 VN.t8 VDD2.t1 w_n2122_n3970# sky130_fd_pr__pfet_01v8 ad=2.47665 pd=15.34 as=2.47665 ps=15.34 w=15.01 l=0.63
X22 VTAIL.t9 VN.t9 VDD2.t0 w_n2122_n3970# sky130_fd_pr__pfet_01v8 ad=2.47665 pd=15.34 as=2.47665 ps=15.34 w=15.01 l=0.63
X23 VTAIL.t10 VP.t9 VDD1.t4 w_n2122_n3970# sky130_fd_pr__pfet_01v8 ad=2.47665 pd=15.34 as=2.47665 ps=15.34 w=15.01 l=0.63
R0 VP.n4 VP.t7 663.75
R1 VP.n10 VP.t1 636.929
R2 VP.n1 VP.t9 636.929
R3 VP.n14 VP.t2 636.929
R4 VP.n15 VP.t0 636.929
R5 VP.n16 VP.t4 636.929
R6 VP.n8 VP.t3 636.929
R7 VP.n7 VP.t5 636.929
R8 VP.n6 VP.t6 636.929
R9 VP.n5 VP.t8 636.929
R10 VP.n17 VP.n16 161.3
R11 VP.n9 VP.n8 161.3
R12 VP.n11 VP.n10 161.3
R13 VP.n6 VP.n3 80.6037
R14 VP.n7 VP.n2 80.6037
R15 VP.n15 VP.n0 80.6037
R16 VP.n14 VP.n13 80.6037
R17 VP.n12 VP.n1 80.6037
R18 VP.n10 VP.n1 48.2005
R19 VP.n14 VP.n1 48.2005
R20 VP.n15 VP.n14 48.2005
R21 VP.n16 VP.n15 48.2005
R22 VP.n8 VP.n7 48.2005
R23 VP.n7 VP.n6 48.2005
R24 VP.n6 VP.n5 48.2005
R25 VP.n4 VP.n3 45.2318
R26 VP.n11 VP.n9 44.7505
R27 VP.n5 VP.n4 13.3799
R28 VP.n3 VP.n2 0.380177
R29 VP.n13 VP.n12 0.380177
R30 VP.n13 VP.n0 0.380177
R31 VP.n9 VP.n2 0.285035
R32 VP.n12 VP.n11 0.285035
R33 VP.n17 VP.n0 0.285035
R34 VP VP.n17 0.0516364
R35 VDD1.n1 VDD1.t0 73.6922
R36 VDD1.n3 VDD1.t6 73.692
R37 VDD1.n5 VDD1.n4 71.2642
R38 VDD1.n1 VDD1.n0 70.6991
R39 VDD1.n7 VDD1.n6 70.6989
R40 VDD1.n3 VDD1.n2 70.6988
R41 VDD1.n7 VDD1.n5 41.5828
R42 VDD1.n6 VDD1.t7 2.16606
R43 VDD1.n6 VDD1.t8 2.16606
R44 VDD1.n0 VDD1.t1 2.16606
R45 VDD1.n0 VDD1.t3 2.16606
R46 VDD1.n4 VDD1.t9 2.16606
R47 VDD1.n4 VDD1.t5 2.16606
R48 VDD1.n2 VDD1.t4 2.16606
R49 VDD1.n2 VDD1.t2 2.16606
R50 VDD1 VDD1.n7 0.563
R51 VDD1 VDD1.n1 0.265586
R52 VDD1.n5 VDD1.n3 0.152051
R53 VTAIL.n11 VTAIL.t0 56.1859
R54 VTAIL.n17 VTAIL.t4 56.1856
R55 VTAIL.n2 VTAIL.t15 56.1856
R56 VTAIL.n16 VTAIL.t16 56.1856
R57 VTAIL.n15 VTAIL.n14 54.0203
R58 VTAIL.n13 VTAIL.n12 54.0203
R59 VTAIL.n10 VTAIL.n9 54.0203
R60 VTAIL.n8 VTAIL.n7 54.0203
R61 VTAIL.n19 VTAIL.n18 54.0201
R62 VTAIL.n1 VTAIL.n0 54.0201
R63 VTAIL.n4 VTAIL.n3 54.0201
R64 VTAIL.n6 VTAIL.n5 54.0201
R65 VTAIL.n8 VTAIL.n6 26.9617
R66 VTAIL.n17 VTAIL.n16 26.1341
R67 VTAIL.n18 VTAIL.t3 2.16606
R68 VTAIL.n18 VTAIL.t6 2.16606
R69 VTAIL.n0 VTAIL.t8 2.16606
R70 VTAIL.n0 VTAIL.t9 2.16606
R71 VTAIL.n3 VTAIL.t17 2.16606
R72 VTAIL.n3 VTAIL.t19 2.16606
R73 VTAIL.n5 VTAIL.t18 2.16606
R74 VTAIL.n5 VTAIL.t10 2.16606
R75 VTAIL.n14 VTAIL.t13 2.16606
R76 VTAIL.n14 VTAIL.t14 2.16606
R77 VTAIL.n12 VTAIL.t12 2.16606
R78 VTAIL.n12 VTAIL.t11 2.16606
R79 VTAIL.n9 VTAIL.t2 2.16606
R80 VTAIL.n9 VTAIL.t7 2.16606
R81 VTAIL.n7 VTAIL.t5 2.16606
R82 VTAIL.n7 VTAIL.t1 2.16606
R83 VTAIL.n13 VTAIL.n11 0.884121
R84 VTAIL.n2 VTAIL.n1 0.884121
R85 VTAIL.n10 VTAIL.n8 0.828086
R86 VTAIL.n11 VTAIL.n10 0.828086
R87 VTAIL.n15 VTAIL.n13 0.828086
R88 VTAIL.n16 VTAIL.n15 0.828086
R89 VTAIL.n6 VTAIL.n4 0.828086
R90 VTAIL.n4 VTAIL.n2 0.828086
R91 VTAIL.n19 VTAIL.n17 0.828086
R92 VTAIL VTAIL.n1 0.679379
R93 VTAIL VTAIL.n19 0.149207
R94 VN.n2 VN.t6 663.75
R95 VN.n10 VN.t2 663.75
R96 VN.n1 VN.t9 636.929
R97 VN.n4 VN.t1 636.929
R98 VN.n5 VN.t8 636.929
R99 VN.n6 VN.t0 636.929
R100 VN.n9 VN.t3 636.929
R101 VN.n12 VN.t4 636.929
R102 VN.n13 VN.t7 636.929
R103 VN.n14 VN.t5 636.929
R104 VN.n7 VN.n6 161.3
R105 VN.n15 VN.n14 161.3
R106 VN.n13 VN.n8 80.6037
R107 VN.n12 VN.n11 80.6037
R108 VN.n5 VN.n0 80.6037
R109 VN.n4 VN.n3 80.6037
R110 VN.n4 VN.n1 48.2005
R111 VN.n5 VN.n4 48.2005
R112 VN.n6 VN.n5 48.2005
R113 VN.n12 VN.n9 48.2005
R114 VN.n13 VN.n12 48.2005
R115 VN.n14 VN.n13 48.2005
R116 VN.n11 VN.n10 45.2318
R117 VN.n3 VN.n2 45.2318
R118 VN VN.n15 45.1312
R119 VN.n10 VN.n9 13.3799
R120 VN.n2 VN.n1 13.3799
R121 VN.n11 VN.n8 0.380177
R122 VN.n3 VN.n0 0.380177
R123 VN.n15 VN.n8 0.285035
R124 VN.n7 VN.n0 0.285035
R125 VN VN.n7 0.0516364
R126 VDD2.n1 VDD2.t3 73.692
R127 VDD2.n4 VDD2.t4 72.8647
R128 VDD2.n3 VDD2.n2 71.2642
R129 VDD2 VDD2.n7 71.2614
R130 VDD2.n6 VDD2.n5 70.6991
R131 VDD2.n1 VDD2.n0 70.6988
R132 VDD2.n4 VDD2.n3 40.586
R133 VDD2.n7 VDD2.t6 2.16606
R134 VDD2.n7 VDD2.t7 2.16606
R135 VDD2.n5 VDD2.t2 2.16606
R136 VDD2.n5 VDD2.t5 2.16606
R137 VDD2.n2 VDD2.t1 2.16606
R138 VDD2.n2 VDD2.t9 2.16606
R139 VDD2.n0 VDD2.t0 2.16606
R140 VDD2.n0 VDD2.t8 2.16606
R141 VDD2.n6 VDD2.n4 0.828086
R142 VDD2 VDD2.n6 0.265586
R143 VDD2.n3 VDD2.n1 0.152051
R144 B.n125 B.t3 778.114
R145 B.n133 B.t6 778.114
R146 B.n40 B.t9 778.114
R147 B.n48 B.t0 778.114
R148 B.n451 B.n74 585
R149 B.n453 B.n452 585
R150 B.n454 B.n73 585
R151 B.n456 B.n455 585
R152 B.n457 B.n72 585
R153 B.n459 B.n458 585
R154 B.n460 B.n71 585
R155 B.n462 B.n461 585
R156 B.n463 B.n70 585
R157 B.n465 B.n464 585
R158 B.n466 B.n69 585
R159 B.n468 B.n467 585
R160 B.n469 B.n68 585
R161 B.n471 B.n470 585
R162 B.n472 B.n67 585
R163 B.n474 B.n473 585
R164 B.n475 B.n66 585
R165 B.n477 B.n476 585
R166 B.n478 B.n65 585
R167 B.n480 B.n479 585
R168 B.n481 B.n64 585
R169 B.n483 B.n482 585
R170 B.n484 B.n63 585
R171 B.n486 B.n485 585
R172 B.n487 B.n62 585
R173 B.n489 B.n488 585
R174 B.n490 B.n61 585
R175 B.n492 B.n491 585
R176 B.n493 B.n60 585
R177 B.n495 B.n494 585
R178 B.n496 B.n59 585
R179 B.n498 B.n497 585
R180 B.n499 B.n58 585
R181 B.n501 B.n500 585
R182 B.n502 B.n57 585
R183 B.n504 B.n503 585
R184 B.n505 B.n56 585
R185 B.n507 B.n506 585
R186 B.n508 B.n55 585
R187 B.n510 B.n509 585
R188 B.n511 B.n54 585
R189 B.n513 B.n512 585
R190 B.n514 B.n53 585
R191 B.n516 B.n515 585
R192 B.n517 B.n52 585
R193 B.n519 B.n518 585
R194 B.n520 B.n51 585
R195 B.n522 B.n521 585
R196 B.n523 B.n47 585
R197 B.n525 B.n524 585
R198 B.n526 B.n46 585
R199 B.n528 B.n527 585
R200 B.n529 B.n45 585
R201 B.n531 B.n530 585
R202 B.n532 B.n44 585
R203 B.n534 B.n533 585
R204 B.n535 B.n43 585
R205 B.n537 B.n536 585
R206 B.n538 B.n42 585
R207 B.n540 B.n539 585
R208 B.n542 B.n39 585
R209 B.n544 B.n543 585
R210 B.n545 B.n38 585
R211 B.n547 B.n546 585
R212 B.n548 B.n37 585
R213 B.n550 B.n549 585
R214 B.n551 B.n36 585
R215 B.n553 B.n552 585
R216 B.n554 B.n35 585
R217 B.n556 B.n555 585
R218 B.n557 B.n34 585
R219 B.n559 B.n558 585
R220 B.n560 B.n33 585
R221 B.n562 B.n561 585
R222 B.n563 B.n32 585
R223 B.n565 B.n564 585
R224 B.n566 B.n31 585
R225 B.n568 B.n567 585
R226 B.n569 B.n30 585
R227 B.n571 B.n570 585
R228 B.n572 B.n29 585
R229 B.n574 B.n573 585
R230 B.n575 B.n28 585
R231 B.n577 B.n576 585
R232 B.n578 B.n27 585
R233 B.n580 B.n579 585
R234 B.n581 B.n26 585
R235 B.n583 B.n582 585
R236 B.n584 B.n25 585
R237 B.n586 B.n585 585
R238 B.n587 B.n24 585
R239 B.n589 B.n588 585
R240 B.n590 B.n23 585
R241 B.n592 B.n591 585
R242 B.n593 B.n22 585
R243 B.n595 B.n594 585
R244 B.n596 B.n21 585
R245 B.n598 B.n597 585
R246 B.n599 B.n20 585
R247 B.n601 B.n600 585
R248 B.n602 B.n19 585
R249 B.n604 B.n603 585
R250 B.n605 B.n18 585
R251 B.n607 B.n606 585
R252 B.n608 B.n17 585
R253 B.n610 B.n609 585
R254 B.n611 B.n16 585
R255 B.n613 B.n612 585
R256 B.n614 B.n15 585
R257 B.n616 B.n615 585
R258 B.n450 B.n449 585
R259 B.n448 B.n75 585
R260 B.n447 B.n446 585
R261 B.n445 B.n76 585
R262 B.n444 B.n443 585
R263 B.n442 B.n77 585
R264 B.n441 B.n440 585
R265 B.n439 B.n78 585
R266 B.n438 B.n437 585
R267 B.n436 B.n79 585
R268 B.n435 B.n434 585
R269 B.n433 B.n80 585
R270 B.n432 B.n431 585
R271 B.n430 B.n81 585
R272 B.n429 B.n428 585
R273 B.n427 B.n82 585
R274 B.n426 B.n425 585
R275 B.n424 B.n83 585
R276 B.n423 B.n422 585
R277 B.n421 B.n84 585
R278 B.n420 B.n419 585
R279 B.n418 B.n85 585
R280 B.n417 B.n416 585
R281 B.n415 B.n86 585
R282 B.n414 B.n413 585
R283 B.n412 B.n87 585
R284 B.n411 B.n410 585
R285 B.n409 B.n88 585
R286 B.n408 B.n407 585
R287 B.n406 B.n89 585
R288 B.n405 B.n404 585
R289 B.n403 B.n90 585
R290 B.n402 B.n401 585
R291 B.n400 B.n91 585
R292 B.n399 B.n398 585
R293 B.n397 B.n92 585
R294 B.n396 B.n395 585
R295 B.n394 B.n93 585
R296 B.n393 B.n392 585
R297 B.n391 B.n94 585
R298 B.n390 B.n389 585
R299 B.n388 B.n95 585
R300 B.n387 B.n386 585
R301 B.n385 B.n96 585
R302 B.n384 B.n383 585
R303 B.n382 B.n97 585
R304 B.n381 B.n380 585
R305 B.n379 B.n98 585
R306 B.n378 B.n377 585
R307 B.n376 B.n99 585
R308 B.n375 B.n374 585
R309 B.n208 B.n159 585
R310 B.n210 B.n209 585
R311 B.n211 B.n158 585
R312 B.n213 B.n212 585
R313 B.n214 B.n157 585
R314 B.n216 B.n215 585
R315 B.n217 B.n156 585
R316 B.n219 B.n218 585
R317 B.n220 B.n155 585
R318 B.n222 B.n221 585
R319 B.n223 B.n154 585
R320 B.n225 B.n224 585
R321 B.n226 B.n153 585
R322 B.n228 B.n227 585
R323 B.n229 B.n152 585
R324 B.n231 B.n230 585
R325 B.n232 B.n151 585
R326 B.n234 B.n233 585
R327 B.n235 B.n150 585
R328 B.n237 B.n236 585
R329 B.n238 B.n149 585
R330 B.n240 B.n239 585
R331 B.n241 B.n148 585
R332 B.n243 B.n242 585
R333 B.n244 B.n147 585
R334 B.n246 B.n245 585
R335 B.n247 B.n146 585
R336 B.n249 B.n248 585
R337 B.n250 B.n145 585
R338 B.n252 B.n251 585
R339 B.n253 B.n144 585
R340 B.n255 B.n254 585
R341 B.n256 B.n143 585
R342 B.n258 B.n257 585
R343 B.n259 B.n142 585
R344 B.n261 B.n260 585
R345 B.n262 B.n141 585
R346 B.n264 B.n263 585
R347 B.n265 B.n140 585
R348 B.n267 B.n266 585
R349 B.n268 B.n139 585
R350 B.n270 B.n269 585
R351 B.n271 B.n138 585
R352 B.n273 B.n272 585
R353 B.n274 B.n137 585
R354 B.n276 B.n275 585
R355 B.n277 B.n136 585
R356 B.n279 B.n278 585
R357 B.n280 B.n135 585
R358 B.n282 B.n281 585
R359 B.n284 B.n132 585
R360 B.n286 B.n285 585
R361 B.n287 B.n131 585
R362 B.n289 B.n288 585
R363 B.n290 B.n130 585
R364 B.n292 B.n291 585
R365 B.n293 B.n129 585
R366 B.n295 B.n294 585
R367 B.n296 B.n128 585
R368 B.n298 B.n297 585
R369 B.n300 B.n299 585
R370 B.n301 B.n124 585
R371 B.n303 B.n302 585
R372 B.n304 B.n123 585
R373 B.n306 B.n305 585
R374 B.n307 B.n122 585
R375 B.n309 B.n308 585
R376 B.n310 B.n121 585
R377 B.n312 B.n311 585
R378 B.n313 B.n120 585
R379 B.n315 B.n314 585
R380 B.n316 B.n119 585
R381 B.n318 B.n317 585
R382 B.n319 B.n118 585
R383 B.n321 B.n320 585
R384 B.n322 B.n117 585
R385 B.n324 B.n323 585
R386 B.n325 B.n116 585
R387 B.n327 B.n326 585
R388 B.n328 B.n115 585
R389 B.n330 B.n329 585
R390 B.n331 B.n114 585
R391 B.n333 B.n332 585
R392 B.n334 B.n113 585
R393 B.n336 B.n335 585
R394 B.n337 B.n112 585
R395 B.n339 B.n338 585
R396 B.n340 B.n111 585
R397 B.n342 B.n341 585
R398 B.n343 B.n110 585
R399 B.n345 B.n344 585
R400 B.n346 B.n109 585
R401 B.n348 B.n347 585
R402 B.n349 B.n108 585
R403 B.n351 B.n350 585
R404 B.n352 B.n107 585
R405 B.n354 B.n353 585
R406 B.n355 B.n106 585
R407 B.n357 B.n356 585
R408 B.n358 B.n105 585
R409 B.n360 B.n359 585
R410 B.n361 B.n104 585
R411 B.n363 B.n362 585
R412 B.n364 B.n103 585
R413 B.n366 B.n365 585
R414 B.n367 B.n102 585
R415 B.n369 B.n368 585
R416 B.n370 B.n101 585
R417 B.n372 B.n371 585
R418 B.n373 B.n100 585
R419 B.n207 B.n206 585
R420 B.n205 B.n160 585
R421 B.n204 B.n203 585
R422 B.n202 B.n161 585
R423 B.n201 B.n200 585
R424 B.n199 B.n162 585
R425 B.n198 B.n197 585
R426 B.n196 B.n163 585
R427 B.n195 B.n194 585
R428 B.n193 B.n164 585
R429 B.n192 B.n191 585
R430 B.n190 B.n165 585
R431 B.n189 B.n188 585
R432 B.n187 B.n166 585
R433 B.n186 B.n185 585
R434 B.n184 B.n167 585
R435 B.n183 B.n182 585
R436 B.n181 B.n168 585
R437 B.n180 B.n179 585
R438 B.n178 B.n169 585
R439 B.n177 B.n176 585
R440 B.n175 B.n170 585
R441 B.n174 B.n173 585
R442 B.n172 B.n171 585
R443 B.n2 B.n0 585
R444 B.n653 B.n1 585
R445 B.n652 B.n651 585
R446 B.n650 B.n3 585
R447 B.n649 B.n648 585
R448 B.n647 B.n4 585
R449 B.n646 B.n645 585
R450 B.n644 B.n5 585
R451 B.n643 B.n642 585
R452 B.n641 B.n6 585
R453 B.n640 B.n639 585
R454 B.n638 B.n7 585
R455 B.n637 B.n636 585
R456 B.n635 B.n8 585
R457 B.n634 B.n633 585
R458 B.n632 B.n9 585
R459 B.n631 B.n630 585
R460 B.n629 B.n10 585
R461 B.n628 B.n627 585
R462 B.n626 B.n11 585
R463 B.n625 B.n624 585
R464 B.n623 B.n12 585
R465 B.n622 B.n621 585
R466 B.n620 B.n13 585
R467 B.n619 B.n618 585
R468 B.n617 B.n14 585
R469 B.n655 B.n654 585
R470 B.n208 B.n207 550.159
R471 B.n617 B.n616 550.159
R472 B.n375 B.n100 550.159
R473 B.n449 B.n74 550.159
R474 B.n207 B.n160 163.367
R475 B.n203 B.n160 163.367
R476 B.n203 B.n202 163.367
R477 B.n202 B.n201 163.367
R478 B.n201 B.n162 163.367
R479 B.n197 B.n162 163.367
R480 B.n197 B.n196 163.367
R481 B.n196 B.n195 163.367
R482 B.n195 B.n164 163.367
R483 B.n191 B.n164 163.367
R484 B.n191 B.n190 163.367
R485 B.n190 B.n189 163.367
R486 B.n189 B.n166 163.367
R487 B.n185 B.n166 163.367
R488 B.n185 B.n184 163.367
R489 B.n184 B.n183 163.367
R490 B.n183 B.n168 163.367
R491 B.n179 B.n168 163.367
R492 B.n179 B.n178 163.367
R493 B.n178 B.n177 163.367
R494 B.n177 B.n170 163.367
R495 B.n173 B.n170 163.367
R496 B.n173 B.n172 163.367
R497 B.n172 B.n2 163.367
R498 B.n654 B.n2 163.367
R499 B.n654 B.n653 163.367
R500 B.n653 B.n652 163.367
R501 B.n652 B.n3 163.367
R502 B.n648 B.n3 163.367
R503 B.n648 B.n647 163.367
R504 B.n647 B.n646 163.367
R505 B.n646 B.n5 163.367
R506 B.n642 B.n5 163.367
R507 B.n642 B.n641 163.367
R508 B.n641 B.n640 163.367
R509 B.n640 B.n7 163.367
R510 B.n636 B.n7 163.367
R511 B.n636 B.n635 163.367
R512 B.n635 B.n634 163.367
R513 B.n634 B.n9 163.367
R514 B.n630 B.n9 163.367
R515 B.n630 B.n629 163.367
R516 B.n629 B.n628 163.367
R517 B.n628 B.n11 163.367
R518 B.n624 B.n11 163.367
R519 B.n624 B.n623 163.367
R520 B.n623 B.n622 163.367
R521 B.n622 B.n13 163.367
R522 B.n618 B.n13 163.367
R523 B.n618 B.n617 163.367
R524 B.n209 B.n208 163.367
R525 B.n209 B.n158 163.367
R526 B.n213 B.n158 163.367
R527 B.n214 B.n213 163.367
R528 B.n215 B.n214 163.367
R529 B.n215 B.n156 163.367
R530 B.n219 B.n156 163.367
R531 B.n220 B.n219 163.367
R532 B.n221 B.n220 163.367
R533 B.n221 B.n154 163.367
R534 B.n225 B.n154 163.367
R535 B.n226 B.n225 163.367
R536 B.n227 B.n226 163.367
R537 B.n227 B.n152 163.367
R538 B.n231 B.n152 163.367
R539 B.n232 B.n231 163.367
R540 B.n233 B.n232 163.367
R541 B.n233 B.n150 163.367
R542 B.n237 B.n150 163.367
R543 B.n238 B.n237 163.367
R544 B.n239 B.n238 163.367
R545 B.n239 B.n148 163.367
R546 B.n243 B.n148 163.367
R547 B.n244 B.n243 163.367
R548 B.n245 B.n244 163.367
R549 B.n245 B.n146 163.367
R550 B.n249 B.n146 163.367
R551 B.n250 B.n249 163.367
R552 B.n251 B.n250 163.367
R553 B.n251 B.n144 163.367
R554 B.n255 B.n144 163.367
R555 B.n256 B.n255 163.367
R556 B.n257 B.n256 163.367
R557 B.n257 B.n142 163.367
R558 B.n261 B.n142 163.367
R559 B.n262 B.n261 163.367
R560 B.n263 B.n262 163.367
R561 B.n263 B.n140 163.367
R562 B.n267 B.n140 163.367
R563 B.n268 B.n267 163.367
R564 B.n269 B.n268 163.367
R565 B.n269 B.n138 163.367
R566 B.n273 B.n138 163.367
R567 B.n274 B.n273 163.367
R568 B.n275 B.n274 163.367
R569 B.n275 B.n136 163.367
R570 B.n279 B.n136 163.367
R571 B.n280 B.n279 163.367
R572 B.n281 B.n280 163.367
R573 B.n281 B.n132 163.367
R574 B.n286 B.n132 163.367
R575 B.n287 B.n286 163.367
R576 B.n288 B.n287 163.367
R577 B.n288 B.n130 163.367
R578 B.n292 B.n130 163.367
R579 B.n293 B.n292 163.367
R580 B.n294 B.n293 163.367
R581 B.n294 B.n128 163.367
R582 B.n298 B.n128 163.367
R583 B.n299 B.n298 163.367
R584 B.n299 B.n124 163.367
R585 B.n303 B.n124 163.367
R586 B.n304 B.n303 163.367
R587 B.n305 B.n304 163.367
R588 B.n305 B.n122 163.367
R589 B.n309 B.n122 163.367
R590 B.n310 B.n309 163.367
R591 B.n311 B.n310 163.367
R592 B.n311 B.n120 163.367
R593 B.n315 B.n120 163.367
R594 B.n316 B.n315 163.367
R595 B.n317 B.n316 163.367
R596 B.n317 B.n118 163.367
R597 B.n321 B.n118 163.367
R598 B.n322 B.n321 163.367
R599 B.n323 B.n322 163.367
R600 B.n323 B.n116 163.367
R601 B.n327 B.n116 163.367
R602 B.n328 B.n327 163.367
R603 B.n329 B.n328 163.367
R604 B.n329 B.n114 163.367
R605 B.n333 B.n114 163.367
R606 B.n334 B.n333 163.367
R607 B.n335 B.n334 163.367
R608 B.n335 B.n112 163.367
R609 B.n339 B.n112 163.367
R610 B.n340 B.n339 163.367
R611 B.n341 B.n340 163.367
R612 B.n341 B.n110 163.367
R613 B.n345 B.n110 163.367
R614 B.n346 B.n345 163.367
R615 B.n347 B.n346 163.367
R616 B.n347 B.n108 163.367
R617 B.n351 B.n108 163.367
R618 B.n352 B.n351 163.367
R619 B.n353 B.n352 163.367
R620 B.n353 B.n106 163.367
R621 B.n357 B.n106 163.367
R622 B.n358 B.n357 163.367
R623 B.n359 B.n358 163.367
R624 B.n359 B.n104 163.367
R625 B.n363 B.n104 163.367
R626 B.n364 B.n363 163.367
R627 B.n365 B.n364 163.367
R628 B.n365 B.n102 163.367
R629 B.n369 B.n102 163.367
R630 B.n370 B.n369 163.367
R631 B.n371 B.n370 163.367
R632 B.n371 B.n100 163.367
R633 B.n376 B.n375 163.367
R634 B.n377 B.n376 163.367
R635 B.n377 B.n98 163.367
R636 B.n381 B.n98 163.367
R637 B.n382 B.n381 163.367
R638 B.n383 B.n382 163.367
R639 B.n383 B.n96 163.367
R640 B.n387 B.n96 163.367
R641 B.n388 B.n387 163.367
R642 B.n389 B.n388 163.367
R643 B.n389 B.n94 163.367
R644 B.n393 B.n94 163.367
R645 B.n394 B.n393 163.367
R646 B.n395 B.n394 163.367
R647 B.n395 B.n92 163.367
R648 B.n399 B.n92 163.367
R649 B.n400 B.n399 163.367
R650 B.n401 B.n400 163.367
R651 B.n401 B.n90 163.367
R652 B.n405 B.n90 163.367
R653 B.n406 B.n405 163.367
R654 B.n407 B.n406 163.367
R655 B.n407 B.n88 163.367
R656 B.n411 B.n88 163.367
R657 B.n412 B.n411 163.367
R658 B.n413 B.n412 163.367
R659 B.n413 B.n86 163.367
R660 B.n417 B.n86 163.367
R661 B.n418 B.n417 163.367
R662 B.n419 B.n418 163.367
R663 B.n419 B.n84 163.367
R664 B.n423 B.n84 163.367
R665 B.n424 B.n423 163.367
R666 B.n425 B.n424 163.367
R667 B.n425 B.n82 163.367
R668 B.n429 B.n82 163.367
R669 B.n430 B.n429 163.367
R670 B.n431 B.n430 163.367
R671 B.n431 B.n80 163.367
R672 B.n435 B.n80 163.367
R673 B.n436 B.n435 163.367
R674 B.n437 B.n436 163.367
R675 B.n437 B.n78 163.367
R676 B.n441 B.n78 163.367
R677 B.n442 B.n441 163.367
R678 B.n443 B.n442 163.367
R679 B.n443 B.n76 163.367
R680 B.n447 B.n76 163.367
R681 B.n448 B.n447 163.367
R682 B.n449 B.n448 163.367
R683 B.n616 B.n15 163.367
R684 B.n612 B.n15 163.367
R685 B.n612 B.n611 163.367
R686 B.n611 B.n610 163.367
R687 B.n610 B.n17 163.367
R688 B.n606 B.n17 163.367
R689 B.n606 B.n605 163.367
R690 B.n605 B.n604 163.367
R691 B.n604 B.n19 163.367
R692 B.n600 B.n19 163.367
R693 B.n600 B.n599 163.367
R694 B.n599 B.n598 163.367
R695 B.n598 B.n21 163.367
R696 B.n594 B.n21 163.367
R697 B.n594 B.n593 163.367
R698 B.n593 B.n592 163.367
R699 B.n592 B.n23 163.367
R700 B.n588 B.n23 163.367
R701 B.n588 B.n587 163.367
R702 B.n587 B.n586 163.367
R703 B.n586 B.n25 163.367
R704 B.n582 B.n25 163.367
R705 B.n582 B.n581 163.367
R706 B.n581 B.n580 163.367
R707 B.n580 B.n27 163.367
R708 B.n576 B.n27 163.367
R709 B.n576 B.n575 163.367
R710 B.n575 B.n574 163.367
R711 B.n574 B.n29 163.367
R712 B.n570 B.n29 163.367
R713 B.n570 B.n569 163.367
R714 B.n569 B.n568 163.367
R715 B.n568 B.n31 163.367
R716 B.n564 B.n31 163.367
R717 B.n564 B.n563 163.367
R718 B.n563 B.n562 163.367
R719 B.n562 B.n33 163.367
R720 B.n558 B.n33 163.367
R721 B.n558 B.n557 163.367
R722 B.n557 B.n556 163.367
R723 B.n556 B.n35 163.367
R724 B.n552 B.n35 163.367
R725 B.n552 B.n551 163.367
R726 B.n551 B.n550 163.367
R727 B.n550 B.n37 163.367
R728 B.n546 B.n37 163.367
R729 B.n546 B.n545 163.367
R730 B.n545 B.n544 163.367
R731 B.n544 B.n39 163.367
R732 B.n539 B.n39 163.367
R733 B.n539 B.n538 163.367
R734 B.n538 B.n537 163.367
R735 B.n537 B.n43 163.367
R736 B.n533 B.n43 163.367
R737 B.n533 B.n532 163.367
R738 B.n532 B.n531 163.367
R739 B.n531 B.n45 163.367
R740 B.n527 B.n45 163.367
R741 B.n527 B.n526 163.367
R742 B.n526 B.n525 163.367
R743 B.n525 B.n47 163.367
R744 B.n521 B.n47 163.367
R745 B.n521 B.n520 163.367
R746 B.n520 B.n519 163.367
R747 B.n519 B.n52 163.367
R748 B.n515 B.n52 163.367
R749 B.n515 B.n514 163.367
R750 B.n514 B.n513 163.367
R751 B.n513 B.n54 163.367
R752 B.n509 B.n54 163.367
R753 B.n509 B.n508 163.367
R754 B.n508 B.n507 163.367
R755 B.n507 B.n56 163.367
R756 B.n503 B.n56 163.367
R757 B.n503 B.n502 163.367
R758 B.n502 B.n501 163.367
R759 B.n501 B.n58 163.367
R760 B.n497 B.n58 163.367
R761 B.n497 B.n496 163.367
R762 B.n496 B.n495 163.367
R763 B.n495 B.n60 163.367
R764 B.n491 B.n60 163.367
R765 B.n491 B.n490 163.367
R766 B.n490 B.n489 163.367
R767 B.n489 B.n62 163.367
R768 B.n485 B.n62 163.367
R769 B.n485 B.n484 163.367
R770 B.n484 B.n483 163.367
R771 B.n483 B.n64 163.367
R772 B.n479 B.n64 163.367
R773 B.n479 B.n478 163.367
R774 B.n478 B.n477 163.367
R775 B.n477 B.n66 163.367
R776 B.n473 B.n66 163.367
R777 B.n473 B.n472 163.367
R778 B.n472 B.n471 163.367
R779 B.n471 B.n68 163.367
R780 B.n467 B.n68 163.367
R781 B.n467 B.n466 163.367
R782 B.n466 B.n465 163.367
R783 B.n465 B.n70 163.367
R784 B.n461 B.n70 163.367
R785 B.n461 B.n460 163.367
R786 B.n460 B.n459 163.367
R787 B.n459 B.n72 163.367
R788 B.n455 B.n72 163.367
R789 B.n455 B.n454 163.367
R790 B.n454 B.n453 163.367
R791 B.n453 B.n74 163.367
R792 B.n125 B.t5 126.147
R793 B.n48 B.t1 126.147
R794 B.n133 B.t8 126.129
R795 B.n40 B.t10 126.129
R796 B.n126 B.t4 107.529
R797 B.n49 B.t2 107.529
R798 B.n134 B.t7 107.51
R799 B.n41 B.t11 107.51
R800 B.n127 B.n126 59.5399
R801 B.n283 B.n134 59.5399
R802 B.n541 B.n41 59.5399
R803 B.n50 B.n49 59.5399
R804 B.n615 B.n14 35.7468
R805 B.n451 B.n450 35.7468
R806 B.n374 B.n373 35.7468
R807 B.n206 B.n159 35.7468
R808 B.n126 B.n125 18.6187
R809 B.n134 B.n133 18.6187
R810 B.n41 B.n40 18.6187
R811 B.n49 B.n48 18.6187
R812 B B.n655 18.0485
R813 B.n615 B.n614 10.6151
R814 B.n614 B.n613 10.6151
R815 B.n613 B.n16 10.6151
R816 B.n609 B.n16 10.6151
R817 B.n609 B.n608 10.6151
R818 B.n608 B.n607 10.6151
R819 B.n607 B.n18 10.6151
R820 B.n603 B.n18 10.6151
R821 B.n603 B.n602 10.6151
R822 B.n602 B.n601 10.6151
R823 B.n601 B.n20 10.6151
R824 B.n597 B.n20 10.6151
R825 B.n597 B.n596 10.6151
R826 B.n596 B.n595 10.6151
R827 B.n595 B.n22 10.6151
R828 B.n591 B.n22 10.6151
R829 B.n591 B.n590 10.6151
R830 B.n590 B.n589 10.6151
R831 B.n589 B.n24 10.6151
R832 B.n585 B.n24 10.6151
R833 B.n585 B.n584 10.6151
R834 B.n584 B.n583 10.6151
R835 B.n583 B.n26 10.6151
R836 B.n579 B.n26 10.6151
R837 B.n579 B.n578 10.6151
R838 B.n578 B.n577 10.6151
R839 B.n577 B.n28 10.6151
R840 B.n573 B.n28 10.6151
R841 B.n573 B.n572 10.6151
R842 B.n572 B.n571 10.6151
R843 B.n571 B.n30 10.6151
R844 B.n567 B.n30 10.6151
R845 B.n567 B.n566 10.6151
R846 B.n566 B.n565 10.6151
R847 B.n565 B.n32 10.6151
R848 B.n561 B.n32 10.6151
R849 B.n561 B.n560 10.6151
R850 B.n560 B.n559 10.6151
R851 B.n559 B.n34 10.6151
R852 B.n555 B.n34 10.6151
R853 B.n555 B.n554 10.6151
R854 B.n554 B.n553 10.6151
R855 B.n553 B.n36 10.6151
R856 B.n549 B.n36 10.6151
R857 B.n549 B.n548 10.6151
R858 B.n548 B.n547 10.6151
R859 B.n547 B.n38 10.6151
R860 B.n543 B.n38 10.6151
R861 B.n543 B.n542 10.6151
R862 B.n540 B.n42 10.6151
R863 B.n536 B.n42 10.6151
R864 B.n536 B.n535 10.6151
R865 B.n535 B.n534 10.6151
R866 B.n534 B.n44 10.6151
R867 B.n530 B.n44 10.6151
R868 B.n530 B.n529 10.6151
R869 B.n529 B.n528 10.6151
R870 B.n528 B.n46 10.6151
R871 B.n524 B.n523 10.6151
R872 B.n523 B.n522 10.6151
R873 B.n522 B.n51 10.6151
R874 B.n518 B.n51 10.6151
R875 B.n518 B.n517 10.6151
R876 B.n517 B.n516 10.6151
R877 B.n516 B.n53 10.6151
R878 B.n512 B.n53 10.6151
R879 B.n512 B.n511 10.6151
R880 B.n511 B.n510 10.6151
R881 B.n510 B.n55 10.6151
R882 B.n506 B.n55 10.6151
R883 B.n506 B.n505 10.6151
R884 B.n505 B.n504 10.6151
R885 B.n504 B.n57 10.6151
R886 B.n500 B.n57 10.6151
R887 B.n500 B.n499 10.6151
R888 B.n499 B.n498 10.6151
R889 B.n498 B.n59 10.6151
R890 B.n494 B.n59 10.6151
R891 B.n494 B.n493 10.6151
R892 B.n493 B.n492 10.6151
R893 B.n492 B.n61 10.6151
R894 B.n488 B.n61 10.6151
R895 B.n488 B.n487 10.6151
R896 B.n487 B.n486 10.6151
R897 B.n486 B.n63 10.6151
R898 B.n482 B.n63 10.6151
R899 B.n482 B.n481 10.6151
R900 B.n481 B.n480 10.6151
R901 B.n480 B.n65 10.6151
R902 B.n476 B.n65 10.6151
R903 B.n476 B.n475 10.6151
R904 B.n475 B.n474 10.6151
R905 B.n474 B.n67 10.6151
R906 B.n470 B.n67 10.6151
R907 B.n470 B.n469 10.6151
R908 B.n469 B.n468 10.6151
R909 B.n468 B.n69 10.6151
R910 B.n464 B.n69 10.6151
R911 B.n464 B.n463 10.6151
R912 B.n463 B.n462 10.6151
R913 B.n462 B.n71 10.6151
R914 B.n458 B.n71 10.6151
R915 B.n458 B.n457 10.6151
R916 B.n457 B.n456 10.6151
R917 B.n456 B.n73 10.6151
R918 B.n452 B.n73 10.6151
R919 B.n452 B.n451 10.6151
R920 B.n374 B.n99 10.6151
R921 B.n378 B.n99 10.6151
R922 B.n379 B.n378 10.6151
R923 B.n380 B.n379 10.6151
R924 B.n380 B.n97 10.6151
R925 B.n384 B.n97 10.6151
R926 B.n385 B.n384 10.6151
R927 B.n386 B.n385 10.6151
R928 B.n386 B.n95 10.6151
R929 B.n390 B.n95 10.6151
R930 B.n391 B.n390 10.6151
R931 B.n392 B.n391 10.6151
R932 B.n392 B.n93 10.6151
R933 B.n396 B.n93 10.6151
R934 B.n397 B.n396 10.6151
R935 B.n398 B.n397 10.6151
R936 B.n398 B.n91 10.6151
R937 B.n402 B.n91 10.6151
R938 B.n403 B.n402 10.6151
R939 B.n404 B.n403 10.6151
R940 B.n404 B.n89 10.6151
R941 B.n408 B.n89 10.6151
R942 B.n409 B.n408 10.6151
R943 B.n410 B.n409 10.6151
R944 B.n410 B.n87 10.6151
R945 B.n414 B.n87 10.6151
R946 B.n415 B.n414 10.6151
R947 B.n416 B.n415 10.6151
R948 B.n416 B.n85 10.6151
R949 B.n420 B.n85 10.6151
R950 B.n421 B.n420 10.6151
R951 B.n422 B.n421 10.6151
R952 B.n422 B.n83 10.6151
R953 B.n426 B.n83 10.6151
R954 B.n427 B.n426 10.6151
R955 B.n428 B.n427 10.6151
R956 B.n428 B.n81 10.6151
R957 B.n432 B.n81 10.6151
R958 B.n433 B.n432 10.6151
R959 B.n434 B.n433 10.6151
R960 B.n434 B.n79 10.6151
R961 B.n438 B.n79 10.6151
R962 B.n439 B.n438 10.6151
R963 B.n440 B.n439 10.6151
R964 B.n440 B.n77 10.6151
R965 B.n444 B.n77 10.6151
R966 B.n445 B.n444 10.6151
R967 B.n446 B.n445 10.6151
R968 B.n446 B.n75 10.6151
R969 B.n450 B.n75 10.6151
R970 B.n210 B.n159 10.6151
R971 B.n211 B.n210 10.6151
R972 B.n212 B.n211 10.6151
R973 B.n212 B.n157 10.6151
R974 B.n216 B.n157 10.6151
R975 B.n217 B.n216 10.6151
R976 B.n218 B.n217 10.6151
R977 B.n218 B.n155 10.6151
R978 B.n222 B.n155 10.6151
R979 B.n223 B.n222 10.6151
R980 B.n224 B.n223 10.6151
R981 B.n224 B.n153 10.6151
R982 B.n228 B.n153 10.6151
R983 B.n229 B.n228 10.6151
R984 B.n230 B.n229 10.6151
R985 B.n230 B.n151 10.6151
R986 B.n234 B.n151 10.6151
R987 B.n235 B.n234 10.6151
R988 B.n236 B.n235 10.6151
R989 B.n236 B.n149 10.6151
R990 B.n240 B.n149 10.6151
R991 B.n241 B.n240 10.6151
R992 B.n242 B.n241 10.6151
R993 B.n242 B.n147 10.6151
R994 B.n246 B.n147 10.6151
R995 B.n247 B.n246 10.6151
R996 B.n248 B.n247 10.6151
R997 B.n248 B.n145 10.6151
R998 B.n252 B.n145 10.6151
R999 B.n253 B.n252 10.6151
R1000 B.n254 B.n253 10.6151
R1001 B.n254 B.n143 10.6151
R1002 B.n258 B.n143 10.6151
R1003 B.n259 B.n258 10.6151
R1004 B.n260 B.n259 10.6151
R1005 B.n260 B.n141 10.6151
R1006 B.n264 B.n141 10.6151
R1007 B.n265 B.n264 10.6151
R1008 B.n266 B.n265 10.6151
R1009 B.n266 B.n139 10.6151
R1010 B.n270 B.n139 10.6151
R1011 B.n271 B.n270 10.6151
R1012 B.n272 B.n271 10.6151
R1013 B.n272 B.n137 10.6151
R1014 B.n276 B.n137 10.6151
R1015 B.n277 B.n276 10.6151
R1016 B.n278 B.n277 10.6151
R1017 B.n278 B.n135 10.6151
R1018 B.n282 B.n135 10.6151
R1019 B.n285 B.n284 10.6151
R1020 B.n285 B.n131 10.6151
R1021 B.n289 B.n131 10.6151
R1022 B.n290 B.n289 10.6151
R1023 B.n291 B.n290 10.6151
R1024 B.n291 B.n129 10.6151
R1025 B.n295 B.n129 10.6151
R1026 B.n296 B.n295 10.6151
R1027 B.n297 B.n296 10.6151
R1028 B.n301 B.n300 10.6151
R1029 B.n302 B.n301 10.6151
R1030 B.n302 B.n123 10.6151
R1031 B.n306 B.n123 10.6151
R1032 B.n307 B.n306 10.6151
R1033 B.n308 B.n307 10.6151
R1034 B.n308 B.n121 10.6151
R1035 B.n312 B.n121 10.6151
R1036 B.n313 B.n312 10.6151
R1037 B.n314 B.n313 10.6151
R1038 B.n314 B.n119 10.6151
R1039 B.n318 B.n119 10.6151
R1040 B.n319 B.n318 10.6151
R1041 B.n320 B.n319 10.6151
R1042 B.n320 B.n117 10.6151
R1043 B.n324 B.n117 10.6151
R1044 B.n325 B.n324 10.6151
R1045 B.n326 B.n325 10.6151
R1046 B.n326 B.n115 10.6151
R1047 B.n330 B.n115 10.6151
R1048 B.n331 B.n330 10.6151
R1049 B.n332 B.n331 10.6151
R1050 B.n332 B.n113 10.6151
R1051 B.n336 B.n113 10.6151
R1052 B.n337 B.n336 10.6151
R1053 B.n338 B.n337 10.6151
R1054 B.n338 B.n111 10.6151
R1055 B.n342 B.n111 10.6151
R1056 B.n343 B.n342 10.6151
R1057 B.n344 B.n343 10.6151
R1058 B.n344 B.n109 10.6151
R1059 B.n348 B.n109 10.6151
R1060 B.n349 B.n348 10.6151
R1061 B.n350 B.n349 10.6151
R1062 B.n350 B.n107 10.6151
R1063 B.n354 B.n107 10.6151
R1064 B.n355 B.n354 10.6151
R1065 B.n356 B.n355 10.6151
R1066 B.n356 B.n105 10.6151
R1067 B.n360 B.n105 10.6151
R1068 B.n361 B.n360 10.6151
R1069 B.n362 B.n361 10.6151
R1070 B.n362 B.n103 10.6151
R1071 B.n366 B.n103 10.6151
R1072 B.n367 B.n366 10.6151
R1073 B.n368 B.n367 10.6151
R1074 B.n368 B.n101 10.6151
R1075 B.n372 B.n101 10.6151
R1076 B.n373 B.n372 10.6151
R1077 B.n206 B.n205 10.6151
R1078 B.n205 B.n204 10.6151
R1079 B.n204 B.n161 10.6151
R1080 B.n200 B.n161 10.6151
R1081 B.n200 B.n199 10.6151
R1082 B.n199 B.n198 10.6151
R1083 B.n198 B.n163 10.6151
R1084 B.n194 B.n163 10.6151
R1085 B.n194 B.n193 10.6151
R1086 B.n193 B.n192 10.6151
R1087 B.n192 B.n165 10.6151
R1088 B.n188 B.n165 10.6151
R1089 B.n188 B.n187 10.6151
R1090 B.n187 B.n186 10.6151
R1091 B.n186 B.n167 10.6151
R1092 B.n182 B.n167 10.6151
R1093 B.n182 B.n181 10.6151
R1094 B.n181 B.n180 10.6151
R1095 B.n180 B.n169 10.6151
R1096 B.n176 B.n169 10.6151
R1097 B.n176 B.n175 10.6151
R1098 B.n175 B.n174 10.6151
R1099 B.n174 B.n171 10.6151
R1100 B.n171 B.n0 10.6151
R1101 B.n651 B.n1 10.6151
R1102 B.n651 B.n650 10.6151
R1103 B.n650 B.n649 10.6151
R1104 B.n649 B.n4 10.6151
R1105 B.n645 B.n4 10.6151
R1106 B.n645 B.n644 10.6151
R1107 B.n644 B.n643 10.6151
R1108 B.n643 B.n6 10.6151
R1109 B.n639 B.n6 10.6151
R1110 B.n639 B.n638 10.6151
R1111 B.n638 B.n637 10.6151
R1112 B.n637 B.n8 10.6151
R1113 B.n633 B.n8 10.6151
R1114 B.n633 B.n632 10.6151
R1115 B.n632 B.n631 10.6151
R1116 B.n631 B.n10 10.6151
R1117 B.n627 B.n10 10.6151
R1118 B.n627 B.n626 10.6151
R1119 B.n626 B.n625 10.6151
R1120 B.n625 B.n12 10.6151
R1121 B.n621 B.n12 10.6151
R1122 B.n621 B.n620 10.6151
R1123 B.n620 B.n619 10.6151
R1124 B.n619 B.n14 10.6151
R1125 B.n542 B.n541 9.36635
R1126 B.n524 B.n50 9.36635
R1127 B.n283 B.n282 9.36635
R1128 B.n300 B.n127 9.36635
R1129 B.n655 B.n0 2.81026
R1130 B.n655 B.n1 2.81026
R1131 B.n541 B.n540 1.24928
R1132 B.n50 B.n46 1.24928
R1133 B.n284 B.n283 1.24928
R1134 B.n297 B.n127 1.24928
C0 VDD1 VP 7.96825f
C1 VTAIL VP 7.48654f
C2 VDD1 VTAIL 18.0123f
C3 w_n2122_n3970# VN 3.98533f
C4 B w_n2122_n3970# 8.08114f
C5 VDD2 w_n2122_n3970# 2.2765f
C6 B VN 0.815665f
C7 VDD2 VN 7.78981f
C8 VDD2 B 1.93215f
C9 w_n2122_n3970# VP 4.25552f
C10 VDD1 w_n2122_n3970# 2.23549f
C11 w_n2122_n3970# VTAIL 3.50042f
C12 VP VN 6.04974f
C13 B VP 1.25915f
C14 VDD1 VN 0.148984f
C15 VTAIL VN 7.47178f
C16 VDD1 B 1.89055f
C17 B VTAIL 3.21284f
C18 VDD2 VP 0.33328f
C19 VDD1 VDD2 0.930581f
C20 VDD2 VTAIL 18.044f
C21 VDD2 VSUBS 1.554574f
C22 VDD1 VSUBS 1.232318f
C23 VTAIL VSUBS 0.825859f
C24 VN VSUBS 5.09807f
C25 VP VSUBS 1.850631f
C26 B VSUBS 3.178122f
C27 w_n2122_n3970# VSUBS 0.103307p
C28 B.n0 VSUBS 0.004482f
C29 B.n1 VSUBS 0.004482f
C30 B.n2 VSUBS 0.007088f
C31 B.n3 VSUBS 0.007088f
C32 B.n4 VSUBS 0.007088f
C33 B.n5 VSUBS 0.007088f
C34 B.n6 VSUBS 0.007088f
C35 B.n7 VSUBS 0.007088f
C36 B.n8 VSUBS 0.007088f
C37 B.n9 VSUBS 0.007088f
C38 B.n10 VSUBS 0.007088f
C39 B.n11 VSUBS 0.007088f
C40 B.n12 VSUBS 0.007088f
C41 B.n13 VSUBS 0.007088f
C42 B.n14 VSUBS 0.017383f
C43 B.n15 VSUBS 0.007088f
C44 B.n16 VSUBS 0.007088f
C45 B.n17 VSUBS 0.007088f
C46 B.n18 VSUBS 0.007088f
C47 B.n19 VSUBS 0.007088f
C48 B.n20 VSUBS 0.007088f
C49 B.n21 VSUBS 0.007088f
C50 B.n22 VSUBS 0.007088f
C51 B.n23 VSUBS 0.007088f
C52 B.n24 VSUBS 0.007088f
C53 B.n25 VSUBS 0.007088f
C54 B.n26 VSUBS 0.007088f
C55 B.n27 VSUBS 0.007088f
C56 B.n28 VSUBS 0.007088f
C57 B.n29 VSUBS 0.007088f
C58 B.n30 VSUBS 0.007088f
C59 B.n31 VSUBS 0.007088f
C60 B.n32 VSUBS 0.007088f
C61 B.n33 VSUBS 0.007088f
C62 B.n34 VSUBS 0.007088f
C63 B.n35 VSUBS 0.007088f
C64 B.n36 VSUBS 0.007088f
C65 B.n37 VSUBS 0.007088f
C66 B.n38 VSUBS 0.007088f
C67 B.n39 VSUBS 0.007088f
C68 B.t11 VSUBS 0.505989f
C69 B.t10 VSUBS 0.514039f
C70 B.t9 VSUBS 0.387254f
C71 B.n40 VSUBS 0.153671f
C72 B.n41 VSUBS 0.064649f
C73 B.n42 VSUBS 0.007088f
C74 B.n43 VSUBS 0.007088f
C75 B.n44 VSUBS 0.007088f
C76 B.n45 VSUBS 0.007088f
C77 B.n46 VSUBS 0.003961f
C78 B.n47 VSUBS 0.007088f
C79 B.t2 VSUBS 0.505974f
C80 B.t1 VSUBS 0.514026f
C81 B.t0 VSUBS 0.387254f
C82 B.n48 VSUBS 0.153685f
C83 B.n49 VSUBS 0.064664f
C84 B.n50 VSUBS 0.016423f
C85 B.n51 VSUBS 0.007088f
C86 B.n52 VSUBS 0.007088f
C87 B.n53 VSUBS 0.007088f
C88 B.n54 VSUBS 0.007088f
C89 B.n55 VSUBS 0.007088f
C90 B.n56 VSUBS 0.007088f
C91 B.n57 VSUBS 0.007088f
C92 B.n58 VSUBS 0.007088f
C93 B.n59 VSUBS 0.007088f
C94 B.n60 VSUBS 0.007088f
C95 B.n61 VSUBS 0.007088f
C96 B.n62 VSUBS 0.007088f
C97 B.n63 VSUBS 0.007088f
C98 B.n64 VSUBS 0.007088f
C99 B.n65 VSUBS 0.007088f
C100 B.n66 VSUBS 0.007088f
C101 B.n67 VSUBS 0.007088f
C102 B.n68 VSUBS 0.007088f
C103 B.n69 VSUBS 0.007088f
C104 B.n70 VSUBS 0.007088f
C105 B.n71 VSUBS 0.007088f
C106 B.n72 VSUBS 0.007088f
C107 B.n73 VSUBS 0.007088f
C108 B.n74 VSUBS 0.01785f
C109 B.n75 VSUBS 0.007088f
C110 B.n76 VSUBS 0.007088f
C111 B.n77 VSUBS 0.007088f
C112 B.n78 VSUBS 0.007088f
C113 B.n79 VSUBS 0.007088f
C114 B.n80 VSUBS 0.007088f
C115 B.n81 VSUBS 0.007088f
C116 B.n82 VSUBS 0.007088f
C117 B.n83 VSUBS 0.007088f
C118 B.n84 VSUBS 0.007088f
C119 B.n85 VSUBS 0.007088f
C120 B.n86 VSUBS 0.007088f
C121 B.n87 VSUBS 0.007088f
C122 B.n88 VSUBS 0.007088f
C123 B.n89 VSUBS 0.007088f
C124 B.n90 VSUBS 0.007088f
C125 B.n91 VSUBS 0.007088f
C126 B.n92 VSUBS 0.007088f
C127 B.n93 VSUBS 0.007088f
C128 B.n94 VSUBS 0.007088f
C129 B.n95 VSUBS 0.007088f
C130 B.n96 VSUBS 0.007088f
C131 B.n97 VSUBS 0.007088f
C132 B.n98 VSUBS 0.007088f
C133 B.n99 VSUBS 0.007088f
C134 B.n100 VSUBS 0.01785f
C135 B.n101 VSUBS 0.007088f
C136 B.n102 VSUBS 0.007088f
C137 B.n103 VSUBS 0.007088f
C138 B.n104 VSUBS 0.007088f
C139 B.n105 VSUBS 0.007088f
C140 B.n106 VSUBS 0.007088f
C141 B.n107 VSUBS 0.007088f
C142 B.n108 VSUBS 0.007088f
C143 B.n109 VSUBS 0.007088f
C144 B.n110 VSUBS 0.007088f
C145 B.n111 VSUBS 0.007088f
C146 B.n112 VSUBS 0.007088f
C147 B.n113 VSUBS 0.007088f
C148 B.n114 VSUBS 0.007088f
C149 B.n115 VSUBS 0.007088f
C150 B.n116 VSUBS 0.007088f
C151 B.n117 VSUBS 0.007088f
C152 B.n118 VSUBS 0.007088f
C153 B.n119 VSUBS 0.007088f
C154 B.n120 VSUBS 0.007088f
C155 B.n121 VSUBS 0.007088f
C156 B.n122 VSUBS 0.007088f
C157 B.n123 VSUBS 0.007088f
C158 B.n124 VSUBS 0.007088f
C159 B.t4 VSUBS 0.505974f
C160 B.t5 VSUBS 0.514026f
C161 B.t3 VSUBS 0.387254f
C162 B.n125 VSUBS 0.153685f
C163 B.n126 VSUBS 0.064664f
C164 B.n127 VSUBS 0.016423f
C165 B.n128 VSUBS 0.007088f
C166 B.n129 VSUBS 0.007088f
C167 B.n130 VSUBS 0.007088f
C168 B.n131 VSUBS 0.007088f
C169 B.n132 VSUBS 0.007088f
C170 B.t7 VSUBS 0.505989f
C171 B.t8 VSUBS 0.514039f
C172 B.t6 VSUBS 0.387254f
C173 B.n133 VSUBS 0.153671f
C174 B.n134 VSUBS 0.064649f
C175 B.n135 VSUBS 0.007088f
C176 B.n136 VSUBS 0.007088f
C177 B.n137 VSUBS 0.007088f
C178 B.n138 VSUBS 0.007088f
C179 B.n139 VSUBS 0.007088f
C180 B.n140 VSUBS 0.007088f
C181 B.n141 VSUBS 0.007088f
C182 B.n142 VSUBS 0.007088f
C183 B.n143 VSUBS 0.007088f
C184 B.n144 VSUBS 0.007088f
C185 B.n145 VSUBS 0.007088f
C186 B.n146 VSUBS 0.007088f
C187 B.n147 VSUBS 0.007088f
C188 B.n148 VSUBS 0.007088f
C189 B.n149 VSUBS 0.007088f
C190 B.n150 VSUBS 0.007088f
C191 B.n151 VSUBS 0.007088f
C192 B.n152 VSUBS 0.007088f
C193 B.n153 VSUBS 0.007088f
C194 B.n154 VSUBS 0.007088f
C195 B.n155 VSUBS 0.007088f
C196 B.n156 VSUBS 0.007088f
C197 B.n157 VSUBS 0.007088f
C198 B.n158 VSUBS 0.007088f
C199 B.n159 VSUBS 0.01785f
C200 B.n160 VSUBS 0.007088f
C201 B.n161 VSUBS 0.007088f
C202 B.n162 VSUBS 0.007088f
C203 B.n163 VSUBS 0.007088f
C204 B.n164 VSUBS 0.007088f
C205 B.n165 VSUBS 0.007088f
C206 B.n166 VSUBS 0.007088f
C207 B.n167 VSUBS 0.007088f
C208 B.n168 VSUBS 0.007088f
C209 B.n169 VSUBS 0.007088f
C210 B.n170 VSUBS 0.007088f
C211 B.n171 VSUBS 0.007088f
C212 B.n172 VSUBS 0.007088f
C213 B.n173 VSUBS 0.007088f
C214 B.n174 VSUBS 0.007088f
C215 B.n175 VSUBS 0.007088f
C216 B.n176 VSUBS 0.007088f
C217 B.n177 VSUBS 0.007088f
C218 B.n178 VSUBS 0.007088f
C219 B.n179 VSUBS 0.007088f
C220 B.n180 VSUBS 0.007088f
C221 B.n181 VSUBS 0.007088f
C222 B.n182 VSUBS 0.007088f
C223 B.n183 VSUBS 0.007088f
C224 B.n184 VSUBS 0.007088f
C225 B.n185 VSUBS 0.007088f
C226 B.n186 VSUBS 0.007088f
C227 B.n187 VSUBS 0.007088f
C228 B.n188 VSUBS 0.007088f
C229 B.n189 VSUBS 0.007088f
C230 B.n190 VSUBS 0.007088f
C231 B.n191 VSUBS 0.007088f
C232 B.n192 VSUBS 0.007088f
C233 B.n193 VSUBS 0.007088f
C234 B.n194 VSUBS 0.007088f
C235 B.n195 VSUBS 0.007088f
C236 B.n196 VSUBS 0.007088f
C237 B.n197 VSUBS 0.007088f
C238 B.n198 VSUBS 0.007088f
C239 B.n199 VSUBS 0.007088f
C240 B.n200 VSUBS 0.007088f
C241 B.n201 VSUBS 0.007088f
C242 B.n202 VSUBS 0.007088f
C243 B.n203 VSUBS 0.007088f
C244 B.n204 VSUBS 0.007088f
C245 B.n205 VSUBS 0.007088f
C246 B.n206 VSUBS 0.017383f
C247 B.n207 VSUBS 0.017383f
C248 B.n208 VSUBS 0.01785f
C249 B.n209 VSUBS 0.007088f
C250 B.n210 VSUBS 0.007088f
C251 B.n211 VSUBS 0.007088f
C252 B.n212 VSUBS 0.007088f
C253 B.n213 VSUBS 0.007088f
C254 B.n214 VSUBS 0.007088f
C255 B.n215 VSUBS 0.007088f
C256 B.n216 VSUBS 0.007088f
C257 B.n217 VSUBS 0.007088f
C258 B.n218 VSUBS 0.007088f
C259 B.n219 VSUBS 0.007088f
C260 B.n220 VSUBS 0.007088f
C261 B.n221 VSUBS 0.007088f
C262 B.n222 VSUBS 0.007088f
C263 B.n223 VSUBS 0.007088f
C264 B.n224 VSUBS 0.007088f
C265 B.n225 VSUBS 0.007088f
C266 B.n226 VSUBS 0.007088f
C267 B.n227 VSUBS 0.007088f
C268 B.n228 VSUBS 0.007088f
C269 B.n229 VSUBS 0.007088f
C270 B.n230 VSUBS 0.007088f
C271 B.n231 VSUBS 0.007088f
C272 B.n232 VSUBS 0.007088f
C273 B.n233 VSUBS 0.007088f
C274 B.n234 VSUBS 0.007088f
C275 B.n235 VSUBS 0.007088f
C276 B.n236 VSUBS 0.007088f
C277 B.n237 VSUBS 0.007088f
C278 B.n238 VSUBS 0.007088f
C279 B.n239 VSUBS 0.007088f
C280 B.n240 VSUBS 0.007088f
C281 B.n241 VSUBS 0.007088f
C282 B.n242 VSUBS 0.007088f
C283 B.n243 VSUBS 0.007088f
C284 B.n244 VSUBS 0.007088f
C285 B.n245 VSUBS 0.007088f
C286 B.n246 VSUBS 0.007088f
C287 B.n247 VSUBS 0.007088f
C288 B.n248 VSUBS 0.007088f
C289 B.n249 VSUBS 0.007088f
C290 B.n250 VSUBS 0.007088f
C291 B.n251 VSUBS 0.007088f
C292 B.n252 VSUBS 0.007088f
C293 B.n253 VSUBS 0.007088f
C294 B.n254 VSUBS 0.007088f
C295 B.n255 VSUBS 0.007088f
C296 B.n256 VSUBS 0.007088f
C297 B.n257 VSUBS 0.007088f
C298 B.n258 VSUBS 0.007088f
C299 B.n259 VSUBS 0.007088f
C300 B.n260 VSUBS 0.007088f
C301 B.n261 VSUBS 0.007088f
C302 B.n262 VSUBS 0.007088f
C303 B.n263 VSUBS 0.007088f
C304 B.n264 VSUBS 0.007088f
C305 B.n265 VSUBS 0.007088f
C306 B.n266 VSUBS 0.007088f
C307 B.n267 VSUBS 0.007088f
C308 B.n268 VSUBS 0.007088f
C309 B.n269 VSUBS 0.007088f
C310 B.n270 VSUBS 0.007088f
C311 B.n271 VSUBS 0.007088f
C312 B.n272 VSUBS 0.007088f
C313 B.n273 VSUBS 0.007088f
C314 B.n274 VSUBS 0.007088f
C315 B.n275 VSUBS 0.007088f
C316 B.n276 VSUBS 0.007088f
C317 B.n277 VSUBS 0.007088f
C318 B.n278 VSUBS 0.007088f
C319 B.n279 VSUBS 0.007088f
C320 B.n280 VSUBS 0.007088f
C321 B.n281 VSUBS 0.007088f
C322 B.n282 VSUBS 0.006671f
C323 B.n283 VSUBS 0.016423f
C324 B.n284 VSUBS 0.003961f
C325 B.n285 VSUBS 0.007088f
C326 B.n286 VSUBS 0.007088f
C327 B.n287 VSUBS 0.007088f
C328 B.n288 VSUBS 0.007088f
C329 B.n289 VSUBS 0.007088f
C330 B.n290 VSUBS 0.007088f
C331 B.n291 VSUBS 0.007088f
C332 B.n292 VSUBS 0.007088f
C333 B.n293 VSUBS 0.007088f
C334 B.n294 VSUBS 0.007088f
C335 B.n295 VSUBS 0.007088f
C336 B.n296 VSUBS 0.007088f
C337 B.n297 VSUBS 0.003961f
C338 B.n298 VSUBS 0.007088f
C339 B.n299 VSUBS 0.007088f
C340 B.n300 VSUBS 0.006671f
C341 B.n301 VSUBS 0.007088f
C342 B.n302 VSUBS 0.007088f
C343 B.n303 VSUBS 0.007088f
C344 B.n304 VSUBS 0.007088f
C345 B.n305 VSUBS 0.007088f
C346 B.n306 VSUBS 0.007088f
C347 B.n307 VSUBS 0.007088f
C348 B.n308 VSUBS 0.007088f
C349 B.n309 VSUBS 0.007088f
C350 B.n310 VSUBS 0.007088f
C351 B.n311 VSUBS 0.007088f
C352 B.n312 VSUBS 0.007088f
C353 B.n313 VSUBS 0.007088f
C354 B.n314 VSUBS 0.007088f
C355 B.n315 VSUBS 0.007088f
C356 B.n316 VSUBS 0.007088f
C357 B.n317 VSUBS 0.007088f
C358 B.n318 VSUBS 0.007088f
C359 B.n319 VSUBS 0.007088f
C360 B.n320 VSUBS 0.007088f
C361 B.n321 VSUBS 0.007088f
C362 B.n322 VSUBS 0.007088f
C363 B.n323 VSUBS 0.007088f
C364 B.n324 VSUBS 0.007088f
C365 B.n325 VSUBS 0.007088f
C366 B.n326 VSUBS 0.007088f
C367 B.n327 VSUBS 0.007088f
C368 B.n328 VSUBS 0.007088f
C369 B.n329 VSUBS 0.007088f
C370 B.n330 VSUBS 0.007088f
C371 B.n331 VSUBS 0.007088f
C372 B.n332 VSUBS 0.007088f
C373 B.n333 VSUBS 0.007088f
C374 B.n334 VSUBS 0.007088f
C375 B.n335 VSUBS 0.007088f
C376 B.n336 VSUBS 0.007088f
C377 B.n337 VSUBS 0.007088f
C378 B.n338 VSUBS 0.007088f
C379 B.n339 VSUBS 0.007088f
C380 B.n340 VSUBS 0.007088f
C381 B.n341 VSUBS 0.007088f
C382 B.n342 VSUBS 0.007088f
C383 B.n343 VSUBS 0.007088f
C384 B.n344 VSUBS 0.007088f
C385 B.n345 VSUBS 0.007088f
C386 B.n346 VSUBS 0.007088f
C387 B.n347 VSUBS 0.007088f
C388 B.n348 VSUBS 0.007088f
C389 B.n349 VSUBS 0.007088f
C390 B.n350 VSUBS 0.007088f
C391 B.n351 VSUBS 0.007088f
C392 B.n352 VSUBS 0.007088f
C393 B.n353 VSUBS 0.007088f
C394 B.n354 VSUBS 0.007088f
C395 B.n355 VSUBS 0.007088f
C396 B.n356 VSUBS 0.007088f
C397 B.n357 VSUBS 0.007088f
C398 B.n358 VSUBS 0.007088f
C399 B.n359 VSUBS 0.007088f
C400 B.n360 VSUBS 0.007088f
C401 B.n361 VSUBS 0.007088f
C402 B.n362 VSUBS 0.007088f
C403 B.n363 VSUBS 0.007088f
C404 B.n364 VSUBS 0.007088f
C405 B.n365 VSUBS 0.007088f
C406 B.n366 VSUBS 0.007088f
C407 B.n367 VSUBS 0.007088f
C408 B.n368 VSUBS 0.007088f
C409 B.n369 VSUBS 0.007088f
C410 B.n370 VSUBS 0.007088f
C411 B.n371 VSUBS 0.007088f
C412 B.n372 VSUBS 0.007088f
C413 B.n373 VSUBS 0.01785f
C414 B.n374 VSUBS 0.017383f
C415 B.n375 VSUBS 0.017383f
C416 B.n376 VSUBS 0.007088f
C417 B.n377 VSUBS 0.007088f
C418 B.n378 VSUBS 0.007088f
C419 B.n379 VSUBS 0.007088f
C420 B.n380 VSUBS 0.007088f
C421 B.n381 VSUBS 0.007088f
C422 B.n382 VSUBS 0.007088f
C423 B.n383 VSUBS 0.007088f
C424 B.n384 VSUBS 0.007088f
C425 B.n385 VSUBS 0.007088f
C426 B.n386 VSUBS 0.007088f
C427 B.n387 VSUBS 0.007088f
C428 B.n388 VSUBS 0.007088f
C429 B.n389 VSUBS 0.007088f
C430 B.n390 VSUBS 0.007088f
C431 B.n391 VSUBS 0.007088f
C432 B.n392 VSUBS 0.007088f
C433 B.n393 VSUBS 0.007088f
C434 B.n394 VSUBS 0.007088f
C435 B.n395 VSUBS 0.007088f
C436 B.n396 VSUBS 0.007088f
C437 B.n397 VSUBS 0.007088f
C438 B.n398 VSUBS 0.007088f
C439 B.n399 VSUBS 0.007088f
C440 B.n400 VSUBS 0.007088f
C441 B.n401 VSUBS 0.007088f
C442 B.n402 VSUBS 0.007088f
C443 B.n403 VSUBS 0.007088f
C444 B.n404 VSUBS 0.007088f
C445 B.n405 VSUBS 0.007088f
C446 B.n406 VSUBS 0.007088f
C447 B.n407 VSUBS 0.007088f
C448 B.n408 VSUBS 0.007088f
C449 B.n409 VSUBS 0.007088f
C450 B.n410 VSUBS 0.007088f
C451 B.n411 VSUBS 0.007088f
C452 B.n412 VSUBS 0.007088f
C453 B.n413 VSUBS 0.007088f
C454 B.n414 VSUBS 0.007088f
C455 B.n415 VSUBS 0.007088f
C456 B.n416 VSUBS 0.007088f
C457 B.n417 VSUBS 0.007088f
C458 B.n418 VSUBS 0.007088f
C459 B.n419 VSUBS 0.007088f
C460 B.n420 VSUBS 0.007088f
C461 B.n421 VSUBS 0.007088f
C462 B.n422 VSUBS 0.007088f
C463 B.n423 VSUBS 0.007088f
C464 B.n424 VSUBS 0.007088f
C465 B.n425 VSUBS 0.007088f
C466 B.n426 VSUBS 0.007088f
C467 B.n427 VSUBS 0.007088f
C468 B.n428 VSUBS 0.007088f
C469 B.n429 VSUBS 0.007088f
C470 B.n430 VSUBS 0.007088f
C471 B.n431 VSUBS 0.007088f
C472 B.n432 VSUBS 0.007088f
C473 B.n433 VSUBS 0.007088f
C474 B.n434 VSUBS 0.007088f
C475 B.n435 VSUBS 0.007088f
C476 B.n436 VSUBS 0.007088f
C477 B.n437 VSUBS 0.007088f
C478 B.n438 VSUBS 0.007088f
C479 B.n439 VSUBS 0.007088f
C480 B.n440 VSUBS 0.007088f
C481 B.n441 VSUBS 0.007088f
C482 B.n442 VSUBS 0.007088f
C483 B.n443 VSUBS 0.007088f
C484 B.n444 VSUBS 0.007088f
C485 B.n445 VSUBS 0.007088f
C486 B.n446 VSUBS 0.007088f
C487 B.n447 VSUBS 0.007088f
C488 B.n448 VSUBS 0.007088f
C489 B.n449 VSUBS 0.017383f
C490 B.n450 VSUBS 0.018149f
C491 B.n451 VSUBS 0.017085f
C492 B.n452 VSUBS 0.007088f
C493 B.n453 VSUBS 0.007088f
C494 B.n454 VSUBS 0.007088f
C495 B.n455 VSUBS 0.007088f
C496 B.n456 VSUBS 0.007088f
C497 B.n457 VSUBS 0.007088f
C498 B.n458 VSUBS 0.007088f
C499 B.n459 VSUBS 0.007088f
C500 B.n460 VSUBS 0.007088f
C501 B.n461 VSUBS 0.007088f
C502 B.n462 VSUBS 0.007088f
C503 B.n463 VSUBS 0.007088f
C504 B.n464 VSUBS 0.007088f
C505 B.n465 VSUBS 0.007088f
C506 B.n466 VSUBS 0.007088f
C507 B.n467 VSUBS 0.007088f
C508 B.n468 VSUBS 0.007088f
C509 B.n469 VSUBS 0.007088f
C510 B.n470 VSUBS 0.007088f
C511 B.n471 VSUBS 0.007088f
C512 B.n472 VSUBS 0.007088f
C513 B.n473 VSUBS 0.007088f
C514 B.n474 VSUBS 0.007088f
C515 B.n475 VSUBS 0.007088f
C516 B.n476 VSUBS 0.007088f
C517 B.n477 VSUBS 0.007088f
C518 B.n478 VSUBS 0.007088f
C519 B.n479 VSUBS 0.007088f
C520 B.n480 VSUBS 0.007088f
C521 B.n481 VSUBS 0.007088f
C522 B.n482 VSUBS 0.007088f
C523 B.n483 VSUBS 0.007088f
C524 B.n484 VSUBS 0.007088f
C525 B.n485 VSUBS 0.007088f
C526 B.n486 VSUBS 0.007088f
C527 B.n487 VSUBS 0.007088f
C528 B.n488 VSUBS 0.007088f
C529 B.n489 VSUBS 0.007088f
C530 B.n490 VSUBS 0.007088f
C531 B.n491 VSUBS 0.007088f
C532 B.n492 VSUBS 0.007088f
C533 B.n493 VSUBS 0.007088f
C534 B.n494 VSUBS 0.007088f
C535 B.n495 VSUBS 0.007088f
C536 B.n496 VSUBS 0.007088f
C537 B.n497 VSUBS 0.007088f
C538 B.n498 VSUBS 0.007088f
C539 B.n499 VSUBS 0.007088f
C540 B.n500 VSUBS 0.007088f
C541 B.n501 VSUBS 0.007088f
C542 B.n502 VSUBS 0.007088f
C543 B.n503 VSUBS 0.007088f
C544 B.n504 VSUBS 0.007088f
C545 B.n505 VSUBS 0.007088f
C546 B.n506 VSUBS 0.007088f
C547 B.n507 VSUBS 0.007088f
C548 B.n508 VSUBS 0.007088f
C549 B.n509 VSUBS 0.007088f
C550 B.n510 VSUBS 0.007088f
C551 B.n511 VSUBS 0.007088f
C552 B.n512 VSUBS 0.007088f
C553 B.n513 VSUBS 0.007088f
C554 B.n514 VSUBS 0.007088f
C555 B.n515 VSUBS 0.007088f
C556 B.n516 VSUBS 0.007088f
C557 B.n517 VSUBS 0.007088f
C558 B.n518 VSUBS 0.007088f
C559 B.n519 VSUBS 0.007088f
C560 B.n520 VSUBS 0.007088f
C561 B.n521 VSUBS 0.007088f
C562 B.n522 VSUBS 0.007088f
C563 B.n523 VSUBS 0.007088f
C564 B.n524 VSUBS 0.006671f
C565 B.n525 VSUBS 0.007088f
C566 B.n526 VSUBS 0.007088f
C567 B.n527 VSUBS 0.007088f
C568 B.n528 VSUBS 0.007088f
C569 B.n529 VSUBS 0.007088f
C570 B.n530 VSUBS 0.007088f
C571 B.n531 VSUBS 0.007088f
C572 B.n532 VSUBS 0.007088f
C573 B.n533 VSUBS 0.007088f
C574 B.n534 VSUBS 0.007088f
C575 B.n535 VSUBS 0.007088f
C576 B.n536 VSUBS 0.007088f
C577 B.n537 VSUBS 0.007088f
C578 B.n538 VSUBS 0.007088f
C579 B.n539 VSUBS 0.007088f
C580 B.n540 VSUBS 0.003961f
C581 B.n541 VSUBS 0.016423f
C582 B.n542 VSUBS 0.006671f
C583 B.n543 VSUBS 0.007088f
C584 B.n544 VSUBS 0.007088f
C585 B.n545 VSUBS 0.007088f
C586 B.n546 VSUBS 0.007088f
C587 B.n547 VSUBS 0.007088f
C588 B.n548 VSUBS 0.007088f
C589 B.n549 VSUBS 0.007088f
C590 B.n550 VSUBS 0.007088f
C591 B.n551 VSUBS 0.007088f
C592 B.n552 VSUBS 0.007088f
C593 B.n553 VSUBS 0.007088f
C594 B.n554 VSUBS 0.007088f
C595 B.n555 VSUBS 0.007088f
C596 B.n556 VSUBS 0.007088f
C597 B.n557 VSUBS 0.007088f
C598 B.n558 VSUBS 0.007088f
C599 B.n559 VSUBS 0.007088f
C600 B.n560 VSUBS 0.007088f
C601 B.n561 VSUBS 0.007088f
C602 B.n562 VSUBS 0.007088f
C603 B.n563 VSUBS 0.007088f
C604 B.n564 VSUBS 0.007088f
C605 B.n565 VSUBS 0.007088f
C606 B.n566 VSUBS 0.007088f
C607 B.n567 VSUBS 0.007088f
C608 B.n568 VSUBS 0.007088f
C609 B.n569 VSUBS 0.007088f
C610 B.n570 VSUBS 0.007088f
C611 B.n571 VSUBS 0.007088f
C612 B.n572 VSUBS 0.007088f
C613 B.n573 VSUBS 0.007088f
C614 B.n574 VSUBS 0.007088f
C615 B.n575 VSUBS 0.007088f
C616 B.n576 VSUBS 0.007088f
C617 B.n577 VSUBS 0.007088f
C618 B.n578 VSUBS 0.007088f
C619 B.n579 VSUBS 0.007088f
C620 B.n580 VSUBS 0.007088f
C621 B.n581 VSUBS 0.007088f
C622 B.n582 VSUBS 0.007088f
C623 B.n583 VSUBS 0.007088f
C624 B.n584 VSUBS 0.007088f
C625 B.n585 VSUBS 0.007088f
C626 B.n586 VSUBS 0.007088f
C627 B.n587 VSUBS 0.007088f
C628 B.n588 VSUBS 0.007088f
C629 B.n589 VSUBS 0.007088f
C630 B.n590 VSUBS 0.007088f
C631 B.n591 VSUBS 0.007088f
C632 B.n592 VSUBS 0.007088f
C633 B.n593 VSUBS 0.007088f
C634 B.n594 VSUBS 0.007088f
C635 B.n595 VSUBS 0.007088f
C636 B.n596 VSUBS 0.007088f
C637 B.n597 VSUBS 0.007088f
C638 B.n598 VSUBS 0.007088f
C639 B.n599 VSUBS 0.007088f
C640 B.n600 VSUBS 0.007088f
C641 B.n601 VSUBS 0.007088f
C642 B.n602 VSUBS 0.007088f
C643 B.n603 VSUBS 0.007088f
C644 B.n604 VSUBS 0.007088f
C645 B.n605 VSUBS 0.007088f
C646 B.n606 VSUBS 0.007088f
C647 B.n607 VSUBS 0.007088f
C648 B.n608 VSUBS 0.007088f
C649 B.n609 VSUBS 0.007088f
C650 B.n610 VSUBS 0.007088f
C651 B.n611 VSUBS 0.007088f
C652 B.n612 VSUBS 0.007088f
C653 B.n613 VSUBS 0.007088f
C654 B.n614 VSUBS 0.007088f
C655 B.n615 VSUBS 0.01785f
C656 B.n616 VSUBS 0.01785f
C657 B.n617 VSUBS 0.017383f
C658 B.n618 VSUBS 0.007088f
C659 B.n619 VSUBS 0.007088f
C660 B.n620 VSUBS 0.007088f
C661 B.n621 VSUBS 0.007088f
C662 B.n622 VSUBS 0.007088f
C663 B.n623 VSUBS 0.007088f
C664 B.n624 VSUBS 0.007088f
C665 B.n625 VSUBS 0.007088f
C666 B.n626 VSUBS 0.007088f
C667 B.n627 VSUBS 0.007088f
C668 B.n628 VSUBS 0.007088f
C669 B.n629 VSUBS 0.007088f
C670 B.n630 VSUBS 0.007088f
C671 B.n631 VSUBS 0.007088f
C672 B.n632 VSUBS 0.007088f
C673 B.n633 VSUBS 0.007088f
C674 B.n634 VSUBS 0.007088f
C675 B.n635 VSUBS 0.007088f
C676 B.n636 VSUBS 0.007088f
C677 B.n637 VSUBS 0.007088f
C678 B.n638 VSUBS 0.007088f
C679 B.n639 VSUBS 0.007088f
C680 B.n640 VSUBS 0.007088f
C681 B.n641 VSUBS 0.007088f
C682 B.n642 VSUBS 0.007088f
C683 B.n643 VSUBS 0.007088f
C684 B.n644 VSUBS 0.007088f
C685 B.n645 VSUBS 0.007088f
C686 B.n646 VSUBS 0.007088f
C687 B.n647 VSUBS 0.007088f
C688 B.n648 VSUBS 0.007088f
C689 B.n649 VSUBS 0.007088f
C690 B.n650 VSUBS 0.007088f
C691 B.n651 VSUBS 0.007088f
C692 B.n652 VSUBS 0.007088f
C693 B.n653 VSUBS 0.007088f
C694 B.n654 VSUBS 0.007088f
C695 B.n655 VSUBS 0.016051f
C696 VDD2.t3 VSUBS 3.40096f
C697 VDD2.t0 VSUBS 0.321629f
C698 VDD2.t8 VSUBS 0.321629f
C699 VDD2.n0 VSUBS 2.61005f
C700 VDD2.n1 VSUBS 1.29777f
C701 VDD2.t1 VSUBS 0.321629f
C702 VDD2.t9 VSUBS 0.321629f
C703 VDD2.n2 VSUBS 2.61523f
C704 VDD2.n3 VSUBS 2.51801f
C705 VDD2.t4 VSUBS 3.39314f
C706 VDD2.n4 VSUBS 3.13295f
C707 VDD2.t2 VSUBS 0.321629f
C708 VDD2.t5 VSUBS 0.321629f
C709 VDD2.n5 VSUBS 2.61006f
C710 VDD2.n6 VSUBS 0.614757f
C711 VDD2.t6 VSUBS 0.321629f
C712 VDD2.t7 VSUBS 0.321629f
C713 VDD2.n7 VSUBS 2.61519f
C714 VN.n0 VSUBS 0.087314f
C715 VN.t9 VSUBS 1.40896f
C716 VN.n1 VSUBS 0.55782f
C717 VN.t6 VSUBS 1.43103f
C718 VN.n2 VSUBS 0.525455f
C719 VN.n3 VSUBS 0.275701f
C720 VN.t1 VSUBS 1.40896f
C721 VN.n4 VSUBS 0.55782f
C722 VN.t8 VSUBS 1.40896f
C723 VN.n5 VSUBS 0.55782f
C724 VN.t0 VSUBS 1.40896f
C725 VN.n6 VSUBS 0.545924f
C726 VN.n7 VSUBS 0.058153f
C727 VN.n8 VSUBS 0.087314f
C728 VN.t3 VSUBS 1.40896f
C729 VN.n9 VSUBS 0.55782f
C730 VN.t4 VSUBS 1.40896f
C731 VN.t2 VSUBS 1.43103f
C732 VN.n10 VSUBS 0.525455f
C733 VN.n11 VSUBS 0.275701f
C734 VN.n12 VSUBS 0.55782f
C735 VN.t7 VSUBS 1.40896f
C736 VN.n13 VSUBS 0.55782f
C737 VN.t5 VSUBS 1.40896f
C738 VN.n14 VSUBS 0.545924f
C739 VN.n15 VSUBS 2.45167f
C740 VTAIL.t8 VSUBS 0.345845f
C741 VTAIL.t9 VSUBS 0.345845f
C742 VTAIL.n0 VSUBS 2.63588f
C743 VTAIL.n1 VSUBS 0.836248f
C744 VTAIL.t15 VSUBS 3.45447f
C745 VTAIL.n2 VSUBS 0.974839f
C746 VTAIL.t17 VSUBS 0.345845f
C747 VTAIL.t19 VSUBS 0.345845f
C748 VTAIL.n3 VSUBS 2.63588f
C749 VTAIL.n4 VSUBS 0.844955f
C750 VTAIL.t18 VSUBS 0.345845f
C751 VTAIL.t10 VSUBS 0.345845f
C752 VTAIL.n5 VSUBS 2.63588f
C753 VTAIL.n6 VSUBS 2.53447f
C754 VTAIL.t5 VSUBS 0.345845f
C755 VTAIL.t1 VSUBS 0.345845f
C756 VTAIL.n7 VSUBS 2.63588f
C757 VTAIL.n8 VSUBS 2.53447f
C758 VTAIL.t2 VSUBS 0.345845f
C759 VTAIL.t7 VSUBS 0.345845f
C760 VTAIL.n9 VSUBS 2.63588f
C761 VTAIL.n10 VSUBS 0.84495f
C762 VTAIL.t0 VSUBS 3.45448f
C763 VTAIL.n11 VSUBS 0.974833f
C764 VTAIL.t12 VSUBS 0.345845f
C765 VTAIL.t11 VSUBS 0.345845f
C766 VTAIL.n12 VSUBS 2.63588f
C767 VTAIL.n13 VSUBS 0.850214f
C768 VTAIL.t13 VSUBS 0.345845f
C769 VTAIL.t14 VSUBS 0.345845f
C770 VTAIL.n14 VSUBS 2.63588f
C771 VTAIL.n15 VSUBS 0.84495f
C772 VTAIL.t16 VSUBS 3.45447f
C773 VTAIL.n16 VSUBS 2.58134f
C774 VTAIL.t4 VSUBS 3.45447f
C775 VTAIL.n17 VSUBS 2.58134f
C776 VTAIL.t3 VSUBS 0.345845f
C777 VTAIL.t6 VSUBS 0.345845f
C778 VTAIL.n18 VSUBS 2.63588f
C779 VTAIL.n19 VSUBS 0.781173f
C780 VDD1.t0 VSUBS 3.40095f
C781 VDD1.t1 VSUBS 0.321627f
C782 VDD1.t3 VSUBS 0.321627f
C783 VDD1.n0 VSUBS 2.61004f
C784 VDD1.n1 VSUBS 1.30353f
C785 VDD1.t6 VSUBS 3.40095f
C786 VDD1.t4 VSUBS 0.321627f
C787 VDD1.t2 VSUBS 0.321627f
C788 VDD1.n2 VSUBS 2.61004f
C789 VDD1.n3 VSUBS 1.29776f
C790 VDD1.t9 VSUBS 0.321627f
C791 VDD1.t5 VSUBS 0.321627f
C792 VDD1.n4 VSUBS 2.61522f
C793 VDD1.n5 VSUBS 2.6006f
C794 VDD1.t7 VSUBS 0.321627f
C795 VDD1.t8 VSUBS 0.321627f
C796 VDD1.n6 VSUBS 2.61003f
C797 VDD1.n7 VSUBS 3.10556f
C798 VP.n0 VSUBS 0.0893f
C799 VP.t9 VSUBS 1.441f
C800 VP.n1 VSUBS 0.570506f
C801 VP.n2 VSUBS 0.0893f
C802 VP.t3 VSUBS 1.441f
C803 VP.t5 VSUBS 1.441f
C804 VP.t6 VSUBS 1.441f
C805 VP.n3 VSUBS 0.28197f
C806 VP.t8 VSUBS 1.441f
C807 VP.t7 VSUBS 1.46357f
C808 VP.n4 VSUBS 0.537404f
C809 VP.n5 VSUBS 0.570506f
C810 VP.n6 VSUBS 0.570506f
C811 VP.n7 VSUBS 0.570506f
C812 VP.n8 VSUBS 0.55834f
C813 VP.n9 VSUBS 2.47236f
C814 VP.t1 VSUBS 1.441f
C815 VP.n10 VSUBS 0.55834f
C816 VP.n11 VSUBS 2.51542f
C817 VP.n12 VSUBS 0.0893f
C818 VP.n13 VSUBS 0.107227f
C819 VP.t2 VSUBS 1.441f
C820 VP.n14 VSUBS 0.570506f
C821 VP.t0 VSUBS 1.441f
C822 VP.n15 VSUBS 0.570506f
C823 VP.t4 VSUBS 1.441f
C824 VP.n16 VSUBS 0.55834f
C825 VP.n17 VSUBS 0.059475f
.ends

