* NGSPICE file created from diff_pair_sample_0323.ext - technology: sky130A

.subckt diff_pair_sample_0323 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t7 VP.t0 VTAIL.t10 w_n4410_n1380# sky130_fd_pr__pfet_01v8 ad=0.3399 pd=2.39 as=0.3399 ps=2.39 w=2.06 l=3.11
X1 B.t11 B.t9 B.t10 w_n4410_n1380# sky130_fd_pr__pfet_01v8 ad=0.8034 pd=4.9 as=0 ps=0 w=2.06 l=3.11
X2 VDD2.t7 VN.t0 VTAIL.t7 w_n4410_n1380# sky130_fd_pr__pfet_01v8 ad=0.3399 pd=2.39 as=0.3399 ps=2.39 w=2.06 l=3.11
X3 VTAIL.t2 VN.t1 VDD2.t6 w_n4410_n1380# sky130_fd_pr__pfet_01v8 ad=0.3399 pd=2.39 as=0.3399 ps=2.39 w=2.06 l=3.11
X4 VTAIL.t14 VP.t1 VDD1.t6 w_n4410_n1380# sky130_fd_pr__pfet_01v8 ad=0.8034 pd=4.9 as=0.3399 ps=2.39 w=2.06 l=3.11
X5 VTAIL.t8 VP.t2 VDD1.t5 w_n4410_n1380# sky130_fd_pr__pfet_01v8 ad=0.8034 pd=4.9 as=0.3399 ps=2.39 w=2.06 l=3.11
X6 VDD2.t5 VN.t2 VTAIL.t1 w_n4410_n1380# sky130_fd_pr__pfet_01v8 ad=0.3399 pd=2.39 as=0.8034 ps=4.9 w=2.06 l=3.11
X7 VTAIL.t0 VN.t3 VDD2.t4 w_n4410_n1380# sky130_fd_pr__pfet_01v8 ad=0.8034 pd=4.9 as=0.3399 ps=2.39 w=2.06 l=3.11
X8 VDD1.t4 VP.t3 VTAIL.t15 w_n4410_n1380# sky130_fd_pr__pfet_01v8 ad=0.3399 pd=2.39 as=0.8034 ps=4.9 w=2.06 l=3.11
X9 B.t8 B.t6 B.t7 w_n4410_n1380# sky130_fd_pr__pfet_01v8 ad=0.8034 pd=4.9 as=0 ps=0 w=2.06 l=3.11
X10 VDD2.t3 VN.t4 VTAIL.t6 w_n4410_n1380# sky130_fd_pr__pfet_01v8 ad=0.3399 pd=2.39 as=0.3399 ps=2.39 w=2.06 l=3.11
X11 VTAIL.t11 VP.t4 VDD1.t3 w_n4410_n1380# sky130_fd_pr__pfet_01v8 ad=0.3399 pd=2.39 as=0.3399 ps=2.39 w=2.06 l=3.11
X12 VTAIL.t4 VN.t5 VDD2.t2 w_n4410_n1380# sky130_fd_pr__pfet_01v8 ad=0.8034 pd=4.9 as=0.3399 ps=2.39 w=2.06 l=3.11
X13 B.t5 B.t3 B.t4 w_n4410_n1380# sky130_fd_pr__pfet_01v8 ad=0.8034 pd=4.9 as=0 ps=0 w=2.06 l=3.11
X14 B.t2 B.t0 B.t1 w_n4410_n1380# sky130_fd_pr__pfet_01v8 ad=0.8034 pd=4.9 as=0 ps=0 w=2.06 l=3.11
X15 VTAIL.t3 VN.t6 VDD2.t1 w_n4410_n1380# sky130_fd_pr__pfet_01v8 ad=0.3399 pd=2.39 as=0.3399 ps=2.39 w=2.06 l=3.11
X16 VDD1.t2 VP.t5 VTAIL.t13 w_n4410_n1380# sky130_fd_pr__pfet_01v8 ad=0.3399 pd=2.39 as=0.3399 ps=2.39 w=2.06 l=3.11
X17 VDD1.t1 VP.t6 VTAIL.t12 w_n4410_n1380# sky130_fd_pr__pfet_01v8 ad=0.3399 pd=2.39 as=0.8034 ps=4.9 w=2.06 l=3.11
X18 VDD2.t0 VN.t7 VTAIL.t5 w_n4410_n1380# sky130_fd_pr__pfet_01v8 ad=0.3399 pd=2.39 as=0.8034 ps=4.9 w=2.06 l=3.11
X19 VTAIL.t9 VP.t7 VDD1.t0 w_n4410_n1380# sky130_fd_pr__pfet_01v8 ad=0.3399 pd=2.39 as=0.3399 ps=2.39 w=2.06 l=3.11
R0 VP.n21 VP.n18 161.3
R1 VP.n23 VP.n22 161.3
R2 VP.n24 VP.n17 161.3
R3 VP.n26 VP.n25 161.3
R4 VP.n27 VP.n16 161.3
R5 VP.n29 VP.n28 161.3
R6 VP.n31 VP.n30 161.3
R7 VP.n32 VP.n14 161.3
R8 VP.n34 VP.n33 161.3
R9 VP.n35 VP.n13 161.3
R10 VP.n37 VP.n36 161.3
R11 VP.n38 VP.n12 161.3
R12 VP.n40 VP.n39 161.3
R13 VP.n75 VP.n74 161.3
R14 VP.n73 VP.n1 161.3
R15 VP.n72 VP.n71 161.3
R16 VP.n70 VP.n2 161.3
R17 VP.n69 VP.n68 161.3
R18 VP.n67 VP.n3 161.3
R19 VP.n66 VP.n65 161.3
R20 VP.n64 VP.n63 161.3
R21 VP.n62 VP.n5 161.3
R22 VP.n61 VP.n60 161.3
R23 VP.n59 VP.n6 161.3
R24 VP.n58 VP.n57 161.3
R25 VP.n56 VP.n7 161.3
R26 VP.n54 VP.n53 161.3
R27 VP.n52 VP.n8 161.3
R28 VP.n51 VP.n50 161.3
R29 VP.n49 VP.n9 161.3
R30 VP.n48 VP.n47 161.3
R31 VP.n46 VP.n10 161.3
R32 VP.n45 VP.n44 161.3
R33 VP.n43 VP.n42 69.9294
R34 VP.n76 VP.n0 69.9294
R35 VP.n41 VP.n11 69.9294
R36 VP.n49 VP.n48 56.4773
R37 VP.n72 VP.n2 56.4773
R38 VP.n37 VP.n13 56.4773
R39 VP.n61 VP.n6 56.4773
R40 VP.n26 VP.n17 56.4773
R41 VP.n20 VP.n19 50.754
R42 VP.n19 VP.t2 49.2866
R43 VP.n42 VP.n41 45.9006
R44 VP.n44 VP.n10 24.3439
R45 VP.n48 VP.n10 24.3439
R46 VP.n50 VP.n49 24.3439
R47 VP.n50 VP.n8 24.3439
R48 VP.n54 VP.n8 24.3439
R49 VP.n57 VP.n56 24.3439
R50 VP.n57 VP.n6 24.3439
R51 VP.n62 VP.n61 24.3439
R52 VP.n63 VP.n62 24.3439
R53 VP.n67 VP.n66 24.3439
R54 VP.n68 VP.n67 24.3439
R55 VP.n68 VP.n2 24.3439
R56 VP.n73 VP.n72 24.3439
R57 VP.n74 VP.n73 24.3439
R58 VP.n38 VP.n37 24.3439
R59 VP.n39 VP.n38 24.3439
R60 VP.n27 VP.n26 24.3439
R61 VP.n28 VP.n27 24.3439
R62 VP.n32 VP.n31 24.3439
R63 VP.n33 VP.n32 24.3439
R64 VP.n33 VP.n13 24.3439
R65 VP.n22 VP.n21 24.3439
R66 VP.n22 VP.n17 24.3439
R67 VP.n56 VP.n55 22.8833
R68 VP.n63 VP.n4 22.8833
R69 VP.n28 VP.n15 22.8833
R70 VP.n21 VP.n20 22.8833
R71 VP.n44 VP.n43 19.9621
R72 VP.n74 VP.n0 19.9621
R73 VP.n39 VP.n11 19.9621
R74 VP.n43 VP.t1 15.9638
R75 VP.n55 VP.t5 15.9638
R76 VP.n4 VP.t7 15.9638
R77 VP.n0 VP.t6 15.9638
R78 VP.n11 VP.t3 15.9638
R79 VP.n15 VP.t4 15.9638
R80 VP.n20 VP.t0 15.9638
R81 VP.n19 VP.n18 3.92639
R82 VP.n55 VP.n54 1.46111
R83 VP.n66 VP.n4 1.46111
R84 VP.n31 VP.n15 1.46111
R85 VP.n41 VP.n40 0.355081
R86 VP.n45 VP.n42 0.355081
R87 VP.n76 VP.n75 0.355081
R88 VP VP.n76 0.26685
R89 VP.n23 VP.n18 0.189894
R90 VP.n24 VP.n23 0.189894
R91 VP.n25 VP.n24 0.189894
R92 VP.n25 VP.n16 0.189894
R93 VP.n29 VP.n16 0.189894
R94 VP.n30 VP.n29 0.189894
R95 VP.n30 VP.n14 0.189894
R96 VP.n34 VP.n14 0.189894
R97 VP.n35 VP.n34 0.189894
R98 VP.n36 VP.n35 0.189894
R99 VP.n36 VP.n12 0.189894
R100 VP.n40 VP.n12 0.189894
R101 VP.n46 VP.n45 0.189894
R102 VP.n47 VP.n46 0.189894
R103 VP.n47 VP.n9 0.189894
R104 VP.n51 VP.n9 0.189894
R105 VP.n52 VP.n51 0.189894
R106 VP.n53 VP.n52 0.189894
R107 VP.n53 VP.n7 0.189894
R108 VP.n58 VP.n7 0.189894
R109 VP.n59 VP.n58 0.189894
R110 VP.n60 VP.n59 0.189894
R111 VP.n60 VP.n5 0.189894
R112 VP.n64 VP.n5 0.189894
R113 VP.n65 VP.n64 0.189894
R114 VP.n65 VP.n3 0.189894
R115 VP.n69 VP.n3 0.189894
R116 VP.n70 VP.n69 0.189894
R117 VP.n71 VP.n70 0.189894
R118 VP.n71 VP.n1 0.189894
R119 VP.n75 VP.n1 0.189894
R120 VTAIL.n15 VTAIL.t5 170.327
R121 VTAIL.n2 VTAIL.t0 170.327
R122 VTAIL.n3 VTAIL.t12 170.327
R123 VTAIL.n6 VTAIL.t14 170.327
R124 VTAIL.n14 VTAIL.t15 170.327
R125 VTAIL.n11 VTAIL.t8 170.327
R126 VTAIL.n10 VTAIL.t1 170.327
R127 VTAIL.n7 VTAIL.t4 170.327
R128 VTAIL.n13 VTAIL.n12 154.548
R129 VTAIL.n9 VTAIL.n8 154.548
R130 VTAIL.n1 VTAIL.n0 154.548
R131 VTAIL.n5 VTAIL.n4 154.548
R132 VTAIL.n15 VTAIL.n14 17.1083
R133 VTAIL.n7 VTAIL.n6 17.1083
R134 VTAIL.n0 VTAIL.t6 15.7796
R135 VTAIL.n0 VTAIL.t3 15.7796
R136 VTAIL.n4 VTAIL.t13 15.7796
R137 VTAIL.n4 VTAIL.t9 15.7796
R138 VTAIL.n12 VTAIL.t10 15.7796
R139 VTAIL.n12 VTAIL.t11 15.7796
R140 VTAIL.n8 VTAIL.t7 15.7796
R141 VTAIL.n8 VTAIL.t2 15.7796
R142 VTAIL.n9 VTAIL.n7 2.96602
R143 VTAIL.n10 VTAIL.n9 2.96602
R144 VTAIL.n13 VTAIL.n11 2.96602
R145 VTAIL.n14 VTAIL.n13 2.96602
R146 VTAIL.n6 VTAIL.n5 2.96602
R147 VTAIL.n5 VTAIL.n3 2.96602
R148 VTAIL.n2 VTAIL.n1 2.96602
R149 VTAIL VTAIL.n15 2.90783
R150 VTAIL.n11 VTAIL.n10 0.470328
R151 VTAIL.n3 VTAIL.n2 0.470328
R152 VTAIL VTAIL.n1 0.0586897
R153 VDD1 VDD1.n0 172.768
R154 VDD1.n3 VDD1.n2 172.655
R155 VDD1.n3 VDD1.n1 172.655
R156 VDD1.n5 VDD1.n4 171.227
R157 VDD1.n5 VDD1.n3 39.419
R158 VDD1.n4 VDD1.t3 15.7796
R159 VDD1.n4 VDD1.t4 15.7796
R160 VDD1.n0 VDD1.t5 15.7796
R161 VDD1.n0 VDD1.t7 15.7796
R162 VDD1.n2 VDD1.t0 15.7796
R163 VDD1.n2 VDD1.t1 15.7796
R164 VDD1.n1 VDD1.t6 15.7796
R165 VDD1.n1 VDD1.t2 15.7796
R166 VDD1 VDD1.n5 1.42507
R167 B.n299 B.n298 585
R168 B.n297 B.n112 585
R169 B.n296 B.n295 585
R170 B.n294 B.n113 585
R171 B.n293 B.n292 585
R172 B.n291 B.n114 585
R173 B.n290 B.n289 585
R174 B.n288 B.n115 585
R175 B.n287 B.n286 585
R176 B.n285 B.n116 585
R177 B.n284 B.n283 585
R178 B.n282 B.n117 585
R179 B.n280 B.n279 585
R180 B.n278 B.n120 585
R181 B.n277 B.n276 585
R182 B.n275 B.n121 585
R183 B.n274 B.n273 585
R184 B.n272 B.n122 585
R185 B.n271 B.n270 585
R186 B.n269 B.n123 585
R187 B.n268 B.n267 585
R188 B.n266 B.n124 585
R189 B.n265 B.n264 585
R190 B.n260 B.n125 585
R191 B.n259 B.n258 585
R192 B.n257 B.n126 585
R193 B.n256 B.n255 585
R194 B.n254 B.n127 585
R195 B.n253 B.n252 585
R196 B.n251 B.n128 585
R197 B.n250 B.n249 585
R198 B.n248 B.n129 585
R199 B.n247 B.n246 585
R200 B.n245 B.n130 585
R201 B.n300 B.n111 585
R202 B.n302 B.n301 585
R203 B.n303 B.n110 585
R204 B.n305 B.n304 585
R205 B.n306 B.n109 585
R206 B.n308 B.n307 585
R207 B.n309 B.n108 585
R208 B.n311 B.n310 585
R209 B.n312 B.n107 585
R210 B.n314 B.n313 585
R211 B.n315 B.n106 585
R212 B.n317 B.n316 585
R213 B.n318 B.n105 585
R214 B.n320 B.n319 585
R215 B.n321 B.n104 585
R216 B.n323 B.n322 585
R217 B.n324 B.n103 585
R218 B.n326 B.n325 585
R219 B.n327 B.n102 585
R220 B.n329 B.n328 585
R221 B.n330 B.n101 585
R222 B.n332 B.n331 585
R223 B.n333 B.n100 585
R224 B.n335 B.n334 585
R225 B.n336 B.n99 585
R226 B.n338 B.n337 585
R227 B.n339 B.n98 585
R228 B.n341 B.n340 585
R229 B.n342 B.n97 585
R230 B.n344 B.n343 585
R231 B.n345 B.n96 585
R232 B.n347 B.n346 585
R233 B.n348 B.n95 585
R234 B.n350 B.n349 585
R235 B.n351 B.n94 585
R236 B.n353 B.n352 585
R237 B.n354 B.n93 585
R238 B.n356 B.n355 585
R239 B.n357 B.n92 585
R240 B.n359 B.n358 585
R241 B.n360 B.n91 585
R242 B.n362 B.n361 585
R243 B.n363 B.n90 585
R244 B.n365 B.n364 585
R245 B.n366 B.n89 585
R246 B.n368 B.n367 585
R247 B.n369 B.n88 585
R248 B.n371 B.n370 585
R249 B.n372 B.n87 585
R250 B.n374 B.n373 585
R251 B.n375 B.n86 585
R252 B.n377 B.n376 585
R253 B.n378 B.n85 585
R254 B.n380 B.n379 585
R255 B.n381 B.n84 585
R256 B.n383 B.n382 585
R257 B.n384 B.n83 585
R258 B.n386 B.n385 585
R259 B.n387 B.n82 585
R260 B.n389 B.n388 585
R261 B.n390 B.n81 585
R262 B.n392 B.n391 585
R263 B.n393 B.n80 585
R264 B.n395 B.n394 585
R265 B.n396 B.n79 585
R266 B.n398 B.n397 585
R267 B.n399 B.n78 585
R268 B.n401 B.n400 585
R269 B.n402 B.n77 585
R270 B.n404 B.n403 585
R271 B.n405 B.n76 585
R272 B.n407 B.n406 585
R273 B.n408 B.n75 585
R274 B.n410 B.n409 585
R275 B.n411 B.n74 585
R276 B.n413 B.n412 585
R277 B.n414 B.n73 585
R278 B.n416 B.n415 585
R279 B.n417 B.n72 585
R280 B.n419 B.n418 585
R281 B.n420 B.n71 585
R282 B.n422 B.n421 585
R283 B.n423 B.n70 585
R284 B.n425 B.n424 585
R285 B.n426 B.n69 585
R286 B.n428 B.n427 585
R287 B.n429 B.n68 585
R288 B.n431 B.n430 585
R289 B.n432 B.n67 585
R290 B.n434 B.n433 585
R291 B.n435 B.n66 585
R292 B.n437 B.n436 585
R293 B.n438 B.n65 585
R294 B.n440 B.n439 585
R295 B.n441 B.n64 585
R296 B.n443 B.n442 585
R297 B.n444 B.n63 585
R298 B.n446 B.n445 585
R299 B.n447 B.n62 585
R300 B.n449 B.n448 585
R301 B.n450 B.n61 585
R302 B.n452 B.n451 585
R303 B.n453 B.n60 585
R304 B.n455 B.n454 585
R305 B.n456 B.n59 585
R306 B.n458 B.n457 585
R307 B.n459 B.n58 585
R308 B.n461 B.n460 585
R309 B.n462 B.n57 585
R310 B.n464 B.n463 585
R311 B.n465 B.n56 585
R312 B.n467 B.n466 585
R313 B.n468 B.n55 585
R314 B.n470 B.n469 585
R315 B.n471 B.n54 585
R316 B.n473 B.n472 585
R317 B.n474 B.n53 585
R318 B.n476 B.n475 585
R319 B.n528 B.n31 585
R320 B.n527 B.n526 585
R321 B.n525 B.n32 585
R322 B.n524 B.n523 585
R323 B.n522 B.n33 585
R324 B.n521 B.n520 585
R325 B.n519 B.n34 585
R326 B.n518 B.n517 585
R327 B.n516 B.n35 585
R328 B.n515 B.n514 585
R329 B.n513 B.n36 585
R330 B.n512 B.n511 585
R331 B.n509 B.n37 585
R332 B.n508 B.n507 585
R333 B.n506 B.n40 585
R334 B.n505 B.n504 585
R335 B.n503 B.n41 585
R336 B.n502 B.n501 585
R337 B.n500 B.n42 585
R338 B.n499 B.n498 585
R339 B.n497 B.n43 585
R340 B.n496 B.n495 585
R341 B.n494 B.n493 585
R342 B.n492 B.n47 585
R343 B.n491 B.n490 585
R344 B.n489 B.n48 585
R345 B.n488 B.n487 585
R346 B.n486 B.n49 585
R347 B.n485 B.n484 585
R348 B.n483 B.n50 585
R349 B.n482 B.n481 585
R350 B.n480 B.n51 585
R351 B.n479 B.n478 585
R352 B.n477 B.n52 585
R353 B.n530 B.n529 585
R354 B.n531 B.n30 585
R355 B.n533 B.n532 585
R356 B.n534 B.n29 585
R357 B.n536 B.n535 585
R358 B.n537 B.n28 585
R359 B.n539 B.n538 585
R360 B.n540 B.n27 585
R361 B.n542 B.n541 585
R362 B.n543 B.n26 585
R363 B.n545 B.n544 585
R364 B.n546 B.n25 585
R365 B.n548 B.n547 585
R366 B.n549 B.n24 585
R367 B.n551 B.n550 585
R368 B.n552 B.n23 585
R369 B.n554 B.n553 585
R370 B.n555 B.n22 585
R371 B.n557 B.n556 585
R372 B.n558 B.n21 585
R373 B.n560 B.n559 585
R374 B.n561 B.n20 585
R375 B.n563 B.n562 585
R376 B.n564 B.n19 585
R377 B.n566 B.n565 585
R378 B.n567 B.n18 585
R379 B.n569 B.n568 585
R380 B.n570 B.n17 585
R381 B.n572 B.n571 585
R382 B.n573 B.n16 585
R383 B.n575 B.n574 585
R384 B.n576 B.n15 585
R385 B.n578 B.n577 585
R386 B.n579 B.n14 585
R387 B.n581 B.n580 585
R388 B.n582 B.n13 585
R389 B.n584 B.n583 585
R390 B.n585 B.n12 585
R391 B.n587 B.n586 585
R392 B.n588 B.n11 585
R393 B.n590 B.n589 585
R394 B.n591 B.n10 585
R395 B.n593 B.n592 585
R396 B.n594 B.n9 585
R397 B.n596 B.n595 585
R398 B.n597 B.n8 585
R399 B.n599 B.n598 585
R400 B.n600 B.n7 585
R401 B.n602 B.n601 585
R402 B.n603 B.n6 585
R403 B.n605 B.n604 585
R404 B.n606 B.n5 585
R405 B.n608 B.n607 585
R406 B.n609 B.n4 585
R407 B.n611 B.n610 585
R408 B.n612 B.n3 585
R409 B.n614 B.n613 585
R410 B.n615 B.n0 585
R411 B.n2 B.n1 585
R412 B.n160 B.n159 585
R413 B.n161 B.n158 585
R414 B.n163 B.n162 585
R415 B.n164 B.n157 585
R416 B.n166 B.n165 585
R417 B.n167 B.n156 585
R418 B.n169 B.n168 585
R419 B.n170 B.n155 585
R420 B.n172 B.n171 585
R421 B.n173 B.n154 585
R422 B.n175 B.n174 585
R423 B.n176 B.n153 585
R424 B.n178 B.n177 585
R425 B.n179 B.n152 585
R426 B.n181 B.n180 585
R427 B.n182 B.n151 585
R428 B.n184 B.n183 585
R429 B.n185 B.n150 585
R430 B.n187 B.n186 585
R431 B.n188 B.n149 585
R432 B.n190 B.n189 585
R433 B.n191 B.n148 585
R434 B.n193 B.n192 585
R435 B.n194 B.n147 585
R436 B.n196 B.n195 585
R437 B.n197 B.n146 585
R438 B.n199 B.n198 585
R439 B.n200 B.n145 585
R440 B.n202 B.n201 585
R441 B.n203 B.n144 585
R442 B.n205 B.n204 585
R443 B.n206 B.n143 585
R444 B.n208 B.n207 585
R445 B.n209 B.n142 585
R446 B.n211 B.n210 585
R447 B.n212 B.n141 585
R448 B.n214 B.n213 585
R449 B.n215 B.n140 585
R450 B.n217 B.n216 585
R451 B.n218 B.n139 585
R452 B.n220 B.n219 585
R453 B.n221 B.n138 585
R454 B.n223 B.n222 585
R455 B.n224 B.n137 585
R456 B.n226 B.n225 585
R457 B.n227 B.n136 585
R458 B.n229 B.n228 585
R459 B.n230 B.n135 585
R460 B.n232 B.n231 585
R461 B.n233 B.n134 585
R462 B.n235 B.n234 585
R463 B.n236 B.n133 585
R464 B.n238 B.n237 585
R465 B.n239 B.n132 585
R466 B.n241 B.n240 585
R467 B.n242 B.n131 585
R468 B.n244 B.n243 585
R469 B.n245 B.n244 559.769
R470 B.n298 B.n111 559.769
R471 B.n477 B.n476 559.769
R472 B.n530 B.n31 559.769
R473 B.n617 B.n616 256.663
R474 B.n118 B.t1 237.852
R475 B.n44 B.t11 237.852
R476 B.n261 B.t7 237.851
R477 B.n38 B.t5 237.851
R478 B.n616 B.n615 235.042
R479 B.n616 B.n2 235.042
R480 B.n261 B.t6 224.669
R481 B.n118 B.t0 224.669
R482 B.n44 B.t9 224.669
R483 B.n38 B.t3 224.669
R484 B.n119 B.t2 171.137
R485 B.n45 B.t10 171.137
R486 B.n262 B.t8 171.137
R487 B.n39 B.t4 171.137
R488 B.n246 B.n245 163.367
R489 B.n246 B.n129 163.367
R490 B.n250 B.n129 163.367
R491 B.n251 B.n250 163.367
R492 B.n252 B.n251 163.367
R493 B.n252 B.n127 163.367
R494 B.n256 B.n127 163.367
R495 B.n257 B.n256 163.367
R496 B.n258 B.n257 163.367
R497 B.n258 B.n125 163.367
R498 B.n265 B.n125 163.367
R499 B.n266 B.n265 163.367
R500 B.n267 B.n266 163.367
R501 B.n267 B.n123 163.367
R502 B.n271 B.n123 163.367
R503 B.n272 B.n271 163.367
R504 B.n273 B.n272 163.367
R505 B.n273 B.n121 163.367
R506 B.n277 B.n121 163.367
R507 B.n278 B.n277 163.367
R508 B.n279 B.n278 163.367
R509 B.n279 B.n117 163.367
R510 B.n284 B.n117 163.367
R511 B.n285 B.n284 163.367
R512 B.n286 B.n285 163.367
R513 B.n286 B.n115 163.367
R514 B.n290 B.n115 163.367
R515 B.n291 B.n290 163.367
R516 B.n292 B.n291 163.367
R517 B.n292 B.n113 163.367
R518 B.n296 B.n113 163.367
R519 B.n297 B.n296 163.367
R520 B.n298 B.n297 163.367
R521 B.n476 B.n53 163.367
R522 B.n472 B.n53 163.367
R523 B.n472 B.n471 163.367
R524 B.n471 B.n470 163.367
R525 B.n470 B.n55 163.367
R526 B.n466 B.n55 163.367
R527 B.n466 B.n465 163.367
R528 B.n465 B.n464 163.367
R529 B.n464 B.n57 163.367
R530 B.n460 B.n57 163.367
R531 B.n460 B.n459 163.367
R532 B.n459 B.n458 163.367
R533 B.n458 B.n59 163.367
R534 B.n454 B.n59 163.367
R535 B.n454 B.n453 163.367
R536 B.n453 B.n452 163.367
R537 B.n452 B.n61 163.367
R538 B.n448 B.n61 163.367
R539 B.n448 B.n447 163.367
R540 B.n447 B.n446 163.367
R541 B.n446 B.n63 163.367
R542 B.n442 B.n63 163.367
R543 B.n442 B.n441 163.367
R544 B.n441 B.n440 163.367
R545 B.n440 B.n65 163.367
R546 B.n436 B.n65 163.367
R547 B.n436 B.n435 163.367
R548 B.n435 B.n434 163.367
R549 B.n434 B.n67 163.367
R550 B.n430 B.n67 163.367
R551 B.n430 B.n429 163.367
R552 B.n429 B.n428 163.367
R553 B.n428 B.n69 163.367
R554 B.n424 B.n69 163.367
R555 B.n424 B.n423 163.367
R556 B.n423 B.n422 163.367
R557 B.n422 B.n71 163.367
R558 B.n418 B.n71 163.367
R559 B.n418 B.n417 163.367
R560 B.n417 B.n416 163.367
R561 B.n416 B.n73 163.367
R562 B.n412 B.n73 163.367
R563 B.n412 B.n411 163.367
R564 B.n411 B.n410 163.367
R565 B.n410 B.n75 163.367
R566 B.n406 B.n75 163.367
R567 B.n406 B.n405 163.367
R568 B.n405 B.n404 163.367
R569 B.n404 B.n77 163.367
R570 B.n400 B.n77 163.367
R571 B.n400 B.n399 163.367
R572 B.n399 B.n398 163.367
R573 B.n398 B.n79 163.367
R574 B.n394 B.n79 163.367
R575 B.n394 B.n393 163.367
R576 B.n393 B.n392 163.367
R577 B.n392 B.n81 163.367
R578 B.n388 B.n81 163.367
R579 B.n388 B.n387 163.367
R580 B.n387 B.n386 163.367
R581 B.n386 B.n83 163.367
R582 B.n382 B.n83 163.367
R583 B.n382 B.n381 163.367
R584 B.n381 B.n380 163.367
R585 B.n380 B.n85 163.367
R586 B.n376 B.n85 163.367
R587 B.n376 B.n375 163.367
R588 B.n375 B.n374 163.367
R589 B.n374 B.n87 163.367
R590 B.n370 B.n87 163.367
R591 B.n370 B.n369 163.367
R592 B.n369 B.n368 163.367
R593 B.n368 B.n89 163.367
R594 B.n364 B.n89 163.367
R595 B.n364 B.n363 163.367
R596 B.n363 B.n362 163.367
R597 B.n362 B.n91 163.367
R598 B.n358 B.n91 163.367
R599 B.n358 B.n357 163.367
R600 B.n357 B.n356 163.367
R601 B.n356 B.n93 163.367
R602 B.n352 B.n93 163.367
R603 B.n352 B.n351 163.367
R604 B.n351 B.n350 163.367
R605 B.n350 B.n95 163.367
R606 B.n346 B.n95 163.367
R607 B.n346 B.n345 163.367
R608 B.n345 B.n344 163.367
R609 B.n344 B.n97 163.367
R610 B.n340 B.n97 163.367
R611 B.n340 B.n339 163.367
R612 B.n339 B.n338 163.367
R613 B.n338 B.n99 163.367
R614 B.n334 B.n99 163.367
R615 B.n334 B.n333 163.367
R616 B.n333 B.n332 163.367
R617 B.n332 B.n101 163.367
R618 B.n328 B.n101 163.367
R619 B.n328 B.n327 163.367
R620 B.n327 B.n326 163.367
R621 B.n326 B.n103 163.367
R622 B.n322 B.n103 163.367
R623 B.n322 B.n321 163.367
R624 B.n321 B.n320 163.367
R625 B.n320 B.n105 163.367
R626 B.n316 B.n105 163.367
R627 B.n316 B.n315 163.367
R628 B.n315 B.n314 163.367
R629 B.n314 B.n107 163.367
R630 B.n310 B.n107 163.367
R631 B.n310 B.n309 163.367
R632 B.n309 B.n308 163.367
R633 B.n308 B.n109 163.367
R634 B.n304 B.n109 163.367
R635 B.n304 B.n303 163.367
R636 B.n303 B.n302 163.367
R637 B.n302 B.n111 163.367
R638 B.n526 B.n31 163.367
R639 B.n526 B.n525 163.367
R640 B.n525 B.n524 163.367
R641 B.n524 B.n33 163.367
R642 B.n520 B.n33 163.367
R643 B.n520 B.n519 163.367
R644 B.n519 B.n518 163.367
R645 B.n518 B.n35 163.367
R646 B.n514 B.n35 163.367
R647 B.n514 B.n513 163.367
R648 B.n513 B.n512 163.367
R649 B.n512 B.n37 163.367
R650 B.n507 B.n37 163.367
R651 B.n507 B.n506 163.367
R652 B.n506 B.n505 163.367
R653 B.n505 B.n41 163.367
R654 B.n501 B.n41 163.367
R655 B.n501 B.n500 163.367
R656 B.n500 B.n499 163.367
R657 B.n499 B.n43 163.367
R658 B.n495 B.n43 163.367
R659 B.n495 B.n494 163.367
R660 B.n494 B.n47 163.367
R661 B.n490 B.n47 163.367
R662 B.n490 B.n489 163.367
R663 B.n489 B.n488 163.367
R664 B.n488 B.n49 163.367
R665 B.n484 B.n49 163.367
R666 B.n484 B.n483 163.367
R667 B.n483 B.n482 163.367
R668 B.n482 B.n51 163.367
R669 B.n478 B.n51 163.367
R670 B.n478 B.n477 163.367
R671 B.n531 B.n530 163.367
R672 B.n532 B.n531 163.367
R673 B.n532 B.n29 163.367
R674 B.n536 B.n29 163.367
R675 B.n537 B.n536 163.367
R676 B.n538 B.n537 163.367
R677 B.n538 B.n27 163.367
R678 B.n542 B.n27 163.367
R679 B.n543 B.n542 163.367
R680 B.n544 B.n543 163.367
R681 B.n544 B.n25 163.367
R682 B.n548 B.n25 163.367
R683 B.n549 B.n548 163.367
R684 B.n550 B.n549 163.367
R685 B.n550 B.n23 163.367
R686 B.n554 B.n23 163.367
R687 B.n555 B.n554 163.367
R688 B.n556 B.n555 163.367
R689 B.n556 B.n21 163.367
R690 B.n560 B.n21 163.367
R691 B.n561 B.n560 163.367
R692 B.n562 B.n561 163.367
R693 B.n562 B.n19 163.367
R694 B.n566 B.n19 163.367
R695 B.n567 B.n566 163.367
R696 B.n568 B.n567 163.367
R697 B.n568 B.n17 163.367
R698 B.n572 B.n17 163.367
R699 B.n573 B.n572 163.367
R700 B.n574 B.n573 163.367
R701 B.n574 B.n15 163.367
R702 B.n578 B.n15 163.367
R703 B.n579 B.n578 163.367
R704 B.n580 B.n579 163.367
R705 B.n580 B.n13 163.367
R706 B.n584 B.n13 163.367
R707 B.n585 B.n584 163.367
R708 B.n586 B.n585 163.367
R709 B.n586 B.n11 163.367
R710 B.n590 B.n11 163.367
R711 B.n591 B.n590 163.367
R712 B.n592 B.n591 163.367
R713 B.n592 B.n9 163.367
R714 B.n596 B.n9 163.367
R715 B.n597 B.n596 163.367
R716 B.n598 B.n597 163.367
R717 B.n598 B.n7 163.367
R718 B.n602 B.n7 163.367
R719 B.n603 B.n602 163.367
R720 B.n604 B.n603 163.367
R721 B.n604 B.n5 163.367
R722 B.n608 B.n5 163.367
R723 B.n609 B.n608 163.367
R724 B.n610 B.n609 163.367
R725 B.n610 B.n3 163.367
R726 B.n614 B.n3 163.367
R727 B.n615 B.n614 163.367
R728 B.n160 B.n2 163.367
R729 B.n161 B.n160 163.367
R730 B.n162 B.n161 163.367
R731 B.n162 B.n157 163.367
R732 B.n166 B.n157 163.367
R733 B.n167 B.n166 163.367
R734 B.n168 B.n167 163.367
R735 B.n168 B.n155 163.367
R736 B.n172 B.n155 163.367
R737 B.n173 B.n172 163.367
R738 B.n174 B.n173 163.367
R739 B.n174 B.n153 163.367
R740 B.n178 B.n153 163.367
R741 B.n179 B.n178 163.367
R742 B.n180 B.n179 163.367
R743 B.n180 B.n151 163.367
R744 B.n184 B.n151 163.367
R745 B.n185 B.n184 163.367
R746 B.n186 B.n185 163.367
R747 B.n186 B.n149 163.367
R748 B.n190 B.n149 163.367
R749 B.n191 B.n190 163.367
R750 B.n192 B.n191 163.367
R751 B.n192 B.n147 163.367
R752 B.n196 B.n147 163.367
R753 B.n197 B.n196 163.367
R754 B.n198 B.n197 163.367
R755 B.n198 B.n145 163.367
R756 B.n202 B.n145 163.367
R757 B.n203 B.n202 163.367
R758 B.n204 B.n203 163.367
R759 B.n204 B.n143 163.367
R760 B.n208 B.n143 163.367
R761 B.n209 B.n208 163.367
R762 B.n210 B.n209 163.367
R763 B.n210 B.n141 163.367
R764 B.n214 B.n141 163.367
R765 B.n215 B.n214 163.367
R766 B.n216 B.n215 163.367
R767 B.n216 B.n139 163.367
R768 B.n220 B.n139 163.367
R769 B.n221 B.n220 163.367
R770 B.n222 B.n221 163.367
R771 B.n222 B.n137 163.367
R772 B.n226 B.n137 163.367
R773 B.n227 B.n226 163.367
R774 B.n228 B.n227 163.367
R775 B.n228 B.n135 163.367
R776 B.n232 B.n135 163.367
R777 B.n233 B.n232 163.367
R778 B.n234 B.n233 163.367
R779 B.n234 B.n133 163.367
R780 B.n238 B.n133 163.367
R781 B.n239 B.n238 163.367
R782 B.n240 B.n239 163.367
R783 B.n240 B.n131 163.367
R784 B.n244 B.n131 163.367
R785 B.n262 B.n261 66.7156
R786 B.n119 B.n118 66.7156
R787 B.n45 B.n44 66.7156
R788 B.n39 B.n38 66.7156
R789 B.n263 B.n262 59.5399
R790 B.n281 B.n119 59.5399
R791 B.n46 B.n45 59.5399
R792 B.n510 B.n39 59.5399
R793 B.n529 B.n528 36.3712
R794 B.n475 B.n52 36.3712
R795 B.n300 B.n299 36.3712
R796 B.n243 B.n130 36.3712
R797 B B.n617 18.0485
R798 B.n529 B.n30 10.6151
R799 B.n533 B.n30 10.6151
R800 B.n534 B.n533 10.6151
R801 B.n535 B.n534 10.6151
R802 B.n535 B.n28 10.6151
R803 B.n539 B.n28 10.6151
R804 B.n540 B.n539 10.6151
R805 B.n541 B.n540 10.6151
R806 B.n541 B.n26 10.6151
R807 B.n545 B.n26 10.6151
R808 B.n546 B.n545 10.6151
R809 B.n547 B.n546 10.6151
R810 B.n547 B.n24 10.6151
R811 B.n551 B.n24 10.6151
R812 B.n552 B.n551 10.6151
R813 B.n553 B.n552 10.6151
R814 B.n553 B.n22 10.6151
R815 B.n557 B.n22 10.6151
R816 B.n558 B.n557 10.6151
R817 B.n559 B.n558 10.6151
R818 B.n559 B.n20 10.6151
R819 B.n563 B.n20 10.6151
R820 B.n564 B.n563 10.6151
R821 B.n565 B.n564 10.6151
R822 B.n565 B.n18 10.6151
R823 B.n569 B.n18 10.6151
R824 B.n570 B.n569 10.6151
R825 B.n571 B.n570 10.6151
R826 B.n571 B.n16 10.6151
R827 B.n575 B.n16 10.6151
R828 B.n576 B.n575 10.6151
R829 B.n577 B.n576 10.6151
R830 B.n577 B.n14 10.6151
R831 B.n581 B.n14 10.6151
R832 B.n582 B.n581 10.6151
R833 B.n583 B.n582 10.6151
R834 B.n583 B.n12 10.6151
R835 B.n587 B.n12 10.6151
R836 B.n588 B.n587 10.6151
R837 B.n589 B.n588 10.6151
R838 B.n589 B.n10 10.6151
R839 B.n593 B.n10 10.6151
R840 B.n594 B.n593 10.6151
R841 B.n595 B.n594 10.6151
R842 B.n595 B.n8 10.6151
R843 B.n599 B.n8 10.6151
R844 B.n600 B.n599 10.6151
R845 B.n601 B.n600 10.6151
R846 B.n601 B.n6 10.6151
R847 B.n605 B.n6 10.6151
R848 B.n606 B.n605 10.6151
R849 B.n607 B.n606 10.6151
R850 B.n607 B.n4 10.6151
R851 B.n611 B.n4 10.6151
R852 B.n612 B.n611 10.6151
R853 B.n613 B.n612 10.6151
R854 B.n613 B.n0 10.6151
R855 B.n528 B.n527 10.6151
R856 B.n527 B.n32 10.6151
R857 B.n523 B.n32 10.6151
R858 B.n523 B.n522 10.6151
R859 B.n522 B.n521 10.6151
R860 B.n521 B.n34 10.6151
R861 B.n517 B.n34 10.6151
R862 B.n517 B.n516 10.6151
R863 B.n516 B.n515 10.6151
R864 B.n515 B.n36 10.6151
R865 B.n511 B.n36 10.6151
R866 B.n509 B.n508 10.6151
R867 B.n508 B.n40 10.6151
R868 B.n504 B.n40 10.6151
R869 B.n504 B.n503 10.6151
R870 B.n503 B.n502 10.6151
R871 B.n502 B.n42 10.6151
R872 B.n498 B.n42 10.6151
R873 B.n498 B.n497 10.6151
R874 B.n497 B.n496 10.6151
R875 B.n493 B.n492 10.6151
R876 B.n492 B.n491 10.6151
R877 B.n491 B.n48 10.6151
R878 B.n487 B.n48 10.6151
R879 B.n487 B.n486 10.6151
R880 B.n486 B.n485 10.6151
R881 B.n485 B.n50 10.6151
R882 B.n481 B.n50 10.6151
R883 B.n481 B.n480 10.6151
R884 B.n480 B.n479 10.6151
R885 B.n479 B.n52 10.6151
R886 B.n475 B.n474 10.6151
R887 B.n474 B.n473 10.6151
R888 B.n473 B.n54 10.6151
R889 B.n469 B.n54 10.6151
R890 B.n469 B.n468 10.6151
R891 B.n468 B.n467 10.6151
R892 B.n467 B.n56 10.6151
R893 B.n463 B.n56 10.6151
R894 B.n463 B.n462 10.6151
R895 B.n462 B.n461 10.6151
R896 B.n461 B.n58 10.6151
R897 B.n457 B.n58 10.6151
R898 B.n457 B.n456 10.6151
R899 B.n456 B.n455 10.6151
R900 B.n455 B.n60 10.6151
R901 B.n451 B.n60 10.6151
R902 B.n451 B.n450 10.6151
R903 B.n450 B.n449 10.6151
R904 B.n449 B.n62 10.6151
R905 B.n445 B.n62 10.6151
R906 B.n445 B.n444 10.6151
R907 B.n444 B.n443 10.6151
R908 B.n443 B.n64 10.6151
R909 B.n439 B.n64 10.6151
R910 B.n439 B.n438 10.6151
R911 B.n438 B.n437 10.6151
R912 B.n437 B.n66 10.6151
R913 B.n433 B.n66 10.6151
R914 B.n433 B.n432 10.6151
R915 B.n432 B.n431 10.6151
R916 B.n431 B.n68 10.6151
R917 B.n427 B.n68 10.6151
R918 B.n427 B.n426 10.6151
R919 B.n426 B.n425 10.6151
R920 B.n425 B.n70 10.6151
R921 B.n421 B.n70 10.6151
R922 B.n421 B.n420 10.6151
R923 B.n420 B.n419 10.6151
R924 B.n419 B.n72 10.6151
R925 B.n415 B.n72 10.6151
R926 B.n415 B.n414 10.6151
R927 B.n414 B.n413 10.6151
R928 B.n413 B.n74 10.6151
R929 B.n409 B.n74 10.6151
R930 B.n409 B.n408 10.6151
R931 B.n408 B.n407 10.6151
R932 B.n407 B.n76 10.6151
R933 B.n403 B.n76 10.6151
R934 B.n403 B.n402 10.6151
R935 B.n402 B.n401 10.6151
R936 B.n401 B.n78 10.6151
R937 B.n397 B.n78 10.6151
R938 B.n397 B.n396 10.6151
R939 B.n396 B.n395 10.6151
R940 B.n395 B.n80 10.6151
R941 B.n391 B.n80 10.6151
R942 B.n391 B.n390 10.6151
R943 B.n390 B.n389 10.6151
R944 B.n389 B.n82 10.6151
R945 B.n385 B.n82 10.6151
R946 B.n385 B.n384 10.6151
R947 B.n384 B.n383 10.6151
R948 B.n383 B.n84 10.6151
R949 B.n379 B.n84 10.6151
R950 B.n379 B.n378 10.6151
R951 B.n378 B.n377 10.6151
R952 B.n377 B.n86 10.6151
R953 B.n373 B.n86 10.6151
R954 B.n373 B.n372 10.6151
R955 B.n372 B.n371 10.6151
R956 B.n371 B.n88 10.6151
R957 B.n367 B.n88 10.6151
R958 B.n367 B.n366 10.6151
R959 B.n366 B.n365 10.6151
R960 B.n365 B.n90 10.6151
R961 B.n361 B.n90 10.6151
R962 B.n361 B.n360 10.6151
R963 B.n360 B.n359 10.6151
R964 B.n359 B.n92 10.6151
R965 B.n355 B.n92 10.6151
R966 B.n355 B.n354 10.6151
R967 B.n354 B.n353 10.6151
R968 B.n353 B.n94 10.6151
R969 B.n349 B.n94 10.6151
R970 B.n349 B.n348 10.6151
R971 B.n348 B.n347 10.6151
R972 B.n347 B.n96 10.6151
R973 B.n343 B.n96 10.6151
R974 B.n343 B.n342 10.6151
R975 B.n342 B.n341 10.6151
R976 B.n341 B.n98 10.6151
R977 B.n337 B.n98 10.6151
R978 B.n337 B.n336 10.6151
R979 B.n336 B.n335 10.6151
R980 B.n335 B.n100 10.6151
R981 B.n331 B.n100 10.6151
R982 B.n331 B.n330 10.6151
R983 B.n330 B.n329 10.6151
R984 B.n329 B.n102 10.6151
R985 B.n325 B.n102 10.6151
R986 B.n325 B.n324 10.6151
R987 B.n324 B.n323 10.6151
R988 B.n323 B.n104 10.6151
R989 B.n319 B.n104 10.6151
R990 B.n319 B.n318 10.6151
R991 B.n318 B.n317 10.6151
R992 B.n317 B.n106 10.6151
R993 B.n313 B.n106 10.6151
R994 B.n313 B.n312 10.6151
R995 B.n312 B.n311 10.6151
R996 B.n311 B.n108 10.6151
R997 B.n307 B.n108 10.6151
R998 B.n307 B.n306 10.6151
R999 B.n306 B.n305 10.6151
R1000 B.n305 B.n110 10.6151
R1001 B.n301 B.n110 10.6151
R1002 B.n301 B.n300 10.6151
R1003 B.n159 B.n1 10.6151
R1004 B.n159 B.n158 10.6151
R1005 B.n163 B.n158 10.6151
R1006 B.n164 B.n163 10.6151
R1007 B.n165 B.n164 10.6151
R1008 B.n165 B.n156 10.6151
R1009 B.n169 B.n156 10.6151
R1010 B.n170 B.n169 10.6151
R1011 B.n171 B.n170 10.6151
R1012 B.n171 B.n154 10.6151
R1013 B.n175 B.n154 10.6151
R1014 B.n176 B.n175 10.6151
R1015 B.n177 B.n176 10.6151
R1016 B.n177 B.n152 10.6151
R1017 B.n181 B.n152 10.6151
R1018 B.n182 B.n181 10.6151
R1019 B.n183 B.n182 10.6151
R1020 B.n183 B.n150 10.6151
R1021 B.n187 B.n150 10.6151
R1022 B.n188 B.n187 10.6151
R1023 B.n189 B.n188 10.6151
R1024 B.n189 B.n148 10.6151
R1025 B.n193 B.n148 10.6151
R1026 B.n194 B.n193 10.6151
R1027 B.n195 B.n194 10.6151
R1028 B.n195 B.n146 10.6151
R1029 B.n199 B.n146 10.6151
R1030 B.n200 B.n199 10.6151
R1031 B.n201 B.n200 10.6151
R1032 B.n201 B.n144 10.6151
R1033 B.n205 B.n144 10.6151
R1034 B.n206 B.n205 10.6151
R1035 B.n207 B.n206 10.6151
R1036 B.n207 B.n142 10.6151
R1037 B.n211 B.n142 10.6151
R1038 B.n212 B.n211 10.6151
R1039 B.n213 B.n212 10.6151
R1040 B.n213 B.n140 10.6151
R1041 B.n217 B.n140 10.6151
R1042 B.n218 B.n217 10.6151
R1043 B.n219 B.n218 10.6151
R1044 B.n219 B.n138 10.6151
R1045 B.n223 B.n138 10.6151
R1046 B.n224 B.n223 10.6151
R1047 B.n225 B.n224 10.6151
R1048 B.n225 B.n136 10.6151
R1049 B.n229 B.n136 10.6151
R1050 B.n230 B.n229 10.6151
R1051 B.n231 B.n230 10.6151
R1052 B.n231 B.n134 10.6151
R1053 B.n235 B.n134 10.6151
R1054 B.n236 B.n235 10.6151
R1055 B.n237 B.n236 10.6151
R1056 B.n237 B.n132 10.6151
R1057 B.n241 B.n132 10.6151
R1058 B.n242 B.n241 10.6151
R1059 B.n243 B.n242 10.6151
R1060 B.n247 B.n130 10.6151
R1061 B.n248 B.n247 10.6151
R1062 B.n249 B.n248 10.6151
R1063 B.n249 B.n128 10.6151
R1064 B.n253 B.n128 10.6151
R1065 B.n254 B.n253 10.6151
R1066 B.n255 B.n254 10.6151
R1067 B.n255 B.n126 10.6151
R1068 B.n259 B.n126 10.6151
R1069 B.n260 B.n259 10.6151
R1070 B.n264 B.n260 10.6151
R1071 B.n268 B.n124 10.6151
R1072 B.n269 B.n268 10.6151
R1073 B.n270 B.n269 10.6151
R1074 B.n270 B.n122 10.6151
R1075 B.n274 B.n122 10.6151
R1076 B.n275 B.n274 10.6151
R1077 B.n276 B.n275 10.6151
R1078 B.n276 B.n120 10.6151
R1079 B.n280 B.n120 10.6151
R1080 B.n283 B.n282 10.6151
R1081 B.n283 B.n116 10.6151
R1082 B.n287 B.n116 10.6151
R1083 B.n288 B.n287 10.6151
R1084 B.n289 B.n288 10.6151
R1085 B.n289 B.n114 10.6151
R1086 B.n293 B.n114 10.6151
R1087 B.n294 B.n293 10.6151
R1088 B.n295 B.n294 10.6151
R1089 B.n295 B.n112 10.6151
R1090 B.n299 B.n112 10.6151
R1091 B.n511 B.n510 9.36635
R1092 B.n493 B.n46 9.36635
R1093 B.n264 B.n263 9.36635
R1094 B.n282 B.n281 9.36635
R1095 B.n617 B.n0 8.11757
R1096 B.n617 B.n1 8.11757
R1097 B.n510 B.n509 1.24928
R1098 B.n496 B.n46 1.24928
R1099 B.n263 B.n124 1.24928
R1100 B.n281 B.n280 1.24928
R1101 VN.n60 VN.n59 161.3
R1102 VN.n58 VN.n32 161.3
R1103 VN.n57 VN.n56 161.3
R1104 VN.n55 VN.n33 161.3
R1105 VN.n54 VN.n53 161.3
R1106 VN.n52 VN.n34 161.3
R1107 VN.n51 VN.n50 161.3
R1108 VN.n49 VN.n48 161.3
R1109 VN.n47 VN.n36 161.3
R1110 VN.n46 VN.n45 161.3
R1111 VN.n44 VN.n37 161.3
R1112 VN.n43 VN.n42 161.3
R1113 VN.n41 VN.n38 161.3
R1114 VN.n29 VN.n28 161.3
R1115 VN.n27 VN.n1 161.3
R1116 VN.n26 VN.n25 161.3
R1117 VN.n24 VN.n2 161.3
R1118 VN.n23 VN.n22 161.3
R1119 VN.n21 VN.n3 161.3
R1120 VN.n20 VN.n19 161.3
R1121 VN.n18 VN.n17 161.3
R1122 VN.n16 VN.n5 161.3
R1123 VN.n15 VN.n14 161.3
R1124 VN.n13 VN.n6 161.3
R1125 VN.n12 VN.n11 161.3
R1126 VN.n10 VN.n7 161.3
R1127 VN.n30 VN.n0 69.9294
R1128 VN.n61 VN.n31 69.9294
R1129 VN.n26 VN.n2 56.4773
R1130 VN.n57 VN.n33 56.4773
R1131 VN.n15 VN.n6 56.4773
R1132 VN.n46 VN.n37 56.4773
R1133 VN.n40 VN.n39 50.754
R1134 VN.n9 VN.n8 50.7539
R1135 VN.n39 VN.t2 49.2868
R1136 VN.n8 VN.t3 49.2868
R1137 VN VN.n61 46.0661
R1138 VN.n11 VN.n10 24.3439
R1139 VN.n11 VN.n6 24.3439
R1140 VN.n16 VN.n15 24.3439
R1141 VN.n17 VN.n16 24.3439
R1142 VN.n21 VN.n20 24.3439
R1143 VN.n22 VN.n21 24.3439
R1144 VN.n22 VN.n2 24.3439
R1145 VN.n27 VN.n26 24.3439
R1146 VN.n28 VN.n27 24.3439
R1147 VN.n42 VN.n37 24.3439
R1148 VN.n42 VN.n41 24.3439
R1149 VN.n53 VN.n33 24.3439
R1150 VN.n53 VN.n52 24.3439
R1151 VN.n52 VN.n51 24.3439
R1152 VN.n48 VN.n47 24.3439
R1153 VN.n47 VN.n46 24.3439
R1154 VN.n59 VN.n58 24.3439
R1155 VN.n58 VN.n57 24.3439
R1156 VN.n10 VN.n9 22.8833
R1157 VN.n17 VN.n4 22.8833
R1158 VN.n41 VN.n40 22.8833
R1159 VN.n48 VN.n35 22.8833
R1160 VN.n28 VN.n0 19.9621
R1161 VN.n59 VN.n31 19.9621
R1162 VN.n9 VN.t4 15.9638
R1163 VN.n4 VN.t6 15.9638
R1164 VN.n0 VN.t7 15.9638
R1165 VN.n40 VN.t1 15.9638
R1166 VN.n35 VN.t0 15.9638
R1167 VN.n31 VN.t5 15.9638
R1168 VN.n39 VN.n38 3.92641
R1169 VN.n8 VN.n7 3.92641
R1170 VN.n20 VN.n4 1.46111
R1171 VN.n51 VN.n35 1.46111
R1172 VN.n61 VN.n60 0.355081
R1173 VN.n30 VN.n29 0.355081
R1174 VN VN.n30 0.26685
R1175 VN.n60 VN.n32 0.189894
R1176 VN.n56 VN.n32 0.189894
R1177 VN.n56 VN.n55 0.189894
R1178 VN.n55 VN.n54 0.189894
R1179 VN.n54 VN.n34 0.189894
R1180 VN.n50 VN.n34 0.189894
R1181 VN.n50 VN.n49 0.189894
R1182 VN.n49 VN.n36 0.189894
R1183 VN.n45 VN.n36 0.189894
R1184 VN.n45 VN.n44 0.189894
R1185 VN.n44 VN.n43 0.189894
R1186 VN.n43 VN.n38 0.189894
R1187 VN.n12 VN.n7 0.189894
R1188 VN.n13 VN.n12 0.189894
R1189 VN.n14 VN.n13 0.189894
R1190 VN.n14 VN.n5 0.189894
R1191 VN.n18 VN.n5 0.189894
R1192 VN.n19 VN.n18 0.189894
R1193 VN.n19 VN.n3 0.189894
R1194 VN.n23 VN.n3 0.189894
R1195 VN.n24 VN.n23 0.189894
R1196 VN.n25 VN.n24 0.189894
R1197 VN.n25 VN.n1 0.189894
R1198 VN.n29 VN.n1 0.189894
R1199 VDD2.n2 VDD2.n1 172.655
R1200 VDD2.n2 VDD2.n0 172.655
R1201 VDD2 VDD2.n5 172.651
R1202 VDD2.n4 VDD2.n3 171.227
R1203 VDD2.n4 VDD2.n2 38.836
R1204 VDD2.n5 VDD2.t6 15.7796
R1205 VDD2.n5 VDD2.t5 15.7796
R1206 VDD2.n3 VDD2.t2 15.7796
R1207 VDD2.n3 VDD2.t7 15.7796
R1208 VDD2.n1 VDD2.t1 15.7796
R1209 VDD2.n1 VDD2.t0 15.7796
R1210 VDD2.n0 VDD2.t4 15.7796
R1211 VDD2.n0 VDD2.t3 15.7796
R1212 VDD2 VDD2.n4 1.54145
C0 VN VP 6.46027f
C1 VDD1 w_n4410_n1380# 1.85047f
C2 VDD1 VTAIL 5.19488f
C3 B VP 2.18996f
C4 VDD2 w_n4410_n1380# 1.98586f
C5 VDD2 VTAIL 5.25271f
C6 VDD1 VP 2.34508f
C7 VTAIL w_n4410_n1380# 2.01317f
C8 VN B 1.22573f
C9 VDD2 VP 0.580771f
C10 VDD1 VN 0.1582f
C11 VP w_n4410_n1380# 9.531839f
C12 VTAIL VP 3.28949f
C13 VDD1 B 1.53599f
C14 VDD2 VN 1.92578f
C15 VN w_n4410_n1380# 8.9622f
C16 VTAIL VN 3.27539f
C17 VDD2 B 1.64846f
C18 B w_n4410_n1380# 8.16916f
C19 VTAIL B 1.74278f
C20 VDD2 VDD1 2.04394f
C21 VDD2 VSUBS 1.49433f
C22 VDD1 VSUBS 2.46754f
C23 VTAIL VSUBS 0.634641f
C24 VN VSUBS 7.39103f
C25 VP VSUBS 3.491042f
C26 B VSUBS 4.440054f
C27 w_n4410_n1380# VSUBS 77.6336f
C28 VDD2.t4 VSUBS 0.039828f
C29 VDD2.t3 VSUBS 0.039828f
C30 VDD2.n0 VSUBS 0.186021f
C31 VDD2.t1 VSUBS 0.039828f
C32 VDD2.t0 VSUBS 0.039828f
C33 VDD2.n1 VSUBS 0.186021f
C34 VDD2.n2 VSUBS 3.03254f
C35 VDD2.t2 VSUBS 0.039828f
C36 VDD2.t7 VSUBS 0.039828f
C37 VDD2.n3 VSUBS 0.180921f
C38 VDD2.n4 VSUBS 2.36492f
C39 VDD2.t6 VSUBS 0.039828f
C40 VDD2.t5 VSUBS 0.039828f
C41 VDD2.n5 VSUBS 0.186005f
C42 VN.t7 VSUBS 0.689026f
C43 VN.n0 VSUBS 0.504495f
C44 VN.n1 VSUBS 0.045785f
C45 VN.n2 VSUBS 0.05942f
C46 VN.n3 VSUBS 0.045785f
C47 VN.t6 VSUBS 0.689026f
C48 VN.n4 VSUBS 0.316357f
C49 VN.n5 VSUBS 0.045785f
C50 VN.n6 VSUBS 0.067129f
C51 VN.n7 VSUBS 0.522833f
C52 VN.t4 VSUBS 0.689026f
C53 VN.t3 VSUBS 1.12508f
C54 VN.n8 VSUBS 0.477921f
C55 VN.n9 VSUBS 0.486289f
C56 VN.n10 VSUBS 0.083219f
C57 VN.n11 VSUBS 0.08576f
C58 VN.n12 VSUBS 0.045785f
C59 VN.n13 VSUBS 0.045785f
C60 VN.n14 VSUBS 0.045785f
C61 VN.n15 VSUBS 0.067129f
C62 VN.n16 VSUBS 0.08576f
C63 VN.n17 VSUBS 0.083219f
C64 VN.n18 VSUBS 0.045785f
C65 VN.n19 VSUBS 0.045785f
C66 VN.n20 VSUBS 0.045958f
C67 VN.n21 VSUBS 0.08576f
C68 VN.n22 VSUBS 0.08576f
C69 VN.n23 VSUBS 0.045785f
C70 VN.n24 VSUBS 0.045785f
C71 VN.n25 VSUBS 0.045785f
C72 VN.n26 VSUBS 0.074839f
C73 VN.n27 VSUBS 0.08576f
C74 VN.n28 VSUBS 0.078138f
C75 VN.n29 VSUBS 0.073908f
C76 VN.n30 VSUBS 0.096875f
C77 VN.t5 VSUBS 0.689026f
C78 VN.n31 VSUBS 0.504495f
C79 VN.n32 VSUBS 0.045785f
C80 VN.n33 VSUBS 0.05942f
C81 VN.n34 VSUBS 0.045785f
C82 VN.t0 VSUBS 0.689026f
C83 VN.n35 VSUBS 0.316357f
C84 VN.n36 VSUBS 0.045785f
C85 VN.n37 VSUBS 0.067129f
C86 VN.n38 VSUBS 0.522833f
C87 VN.t1 VSUBS 0.689026f
C88 VN.t2 VSUBS 1.12508f
C89 VN.n39 VSUBS 0.477921f
C90 VN.n40 VSUBS 0.486289f
C91 VN.n41 VSUBS 0.083219f
C92 VN.n42 VSUBS 0.08576f
C93 VN.n43 VSUBS 0.045785f
C94 VN.n44 VSUBS 0.045785f
C95 VN.n45 VSUBS 0.045785f
C96 VN.n46 VSUBS 0.067129f
C97 VN.n47 VSUBS 0.08576f
C98 VN.n48 VSUBS 0.083219f
C99 VN.n49 VSUBS 0.045785f
C100 VN.n50 VSUBS 0.045785f
C101 VN.n51 VSUBS 0.045958f
C102 VN.n52 VSUBS 0.08576f
C103 VN.n53 VSUBS 0.08576f
C104 VN.n54 VSUBS 0.045785f
C105 VN.n55 VSUBS 0.045785f
C106 VN.n56 VSUBS 0.045785f
C107 VN.n57 VSUBS 0.074839f
C108 VN.n58 VSUBS 0.08576f
C109 VN.n59 VSUBS 0.078138f
C110 VN.n60 VSUBS 0.073908f
C111 VN.n61 VSUBS 2.3038f
C112 B.n0 VSUBS 0.009564f
C113 B.n1 VSUBS 0.009564f
C114 B.n2 VSUBS 0.014144f
C115 B.n3 VSUBS 0.010839f
C116 B.n4 VSUBS 0.010839f
C117 B.n5 VSUBS 0.010839f
C118 B.n6 VSUBS 0.010839f
C119 B.n7 VSUBS 0.010839f
C120 B.n8 VSUBS 0.010839f
C121 B.n9 VSUBS 0.010839f
C122 B.n10 VSUBS 0.010839f
C123 B.n11 VSUBS 0.010839f
C124 B.n12 VSUBS 0.010839f
C125 B.n13 VSUBS 0.010839f
C126 B.n14 VSUBS 0.010839f
C127 B.n15 VSUBS 0.010839f
C128 B.n16 VSUBS 0.010839f
C129 B.n17 VSUBS 0.010839f
C130 B.n18 VSUBS 0.010839f
C131 B.n19 VSUBS 0.010839f
C132 B.n20 VSUBS 0.010839f
C133 B.n21 VSUBS 0.010839f
C134 B.n22 VSUBS 0.010839f
C135 B.n23 VSUBS 0.010839f
C136 B.n24 VSUBS 0.010839f
C137 B.n25 VSUBS 0.010839f
C138 B.n26 VSUBS 0.010839f
C139 B.n27 VSUBS 0.010839f
C140 B.n28 VSUBS 0.010839f
C141 B.n29 VSUBS 0.010839f
C142 B.n30 VSUBS 0.010839f
C143 B.n31 VSUBS 0.027831f
C144 B.n32 VSUBS 0.010839f
C145 B.n33 VSUBS 0.010839f
C146 B.n34 VSUBS 0.010839f
C147 B.n35 VSUBS 0.010839f
C148 B.n36 VSUBS 0.010839f
C149 B.n37 VSUBS 0.010839f
C150 B.t4 VSUBS 0.069458f
C151 B.t5 VSUBS 0.091499f
C152 B.t3 VSUBS 0.489647f
C153 B.n38 VSUBS 0.117628f
C154 B.n39 VSUBS 0.09404f
C155 B.n40 VSUBS 0.010839f
C156 B.n41 VSUBS 0.010839f
C157 B.n42 VSUBS 0.010839f
C158 B.n43 VSUBS 0.010839f
C159 B.t10 VSUBS 0.069458f
C160 B.t11 VSUBS 0.091499f
C161 B.t9 VSUBS 0.489647f
C162 B.n44 VSUBS 0.117628f
C163 B.n45 VSUBS 0.09404f
C164 B.n46 VSUBS 0.025112f
C165 B.n47 VSUBS 0.010839f
C166 B.n48 VSUBS 0.010839f
C167 B.n49 VSUBS 0.010839f
C168 B.n50 VSUBS 0.010839f
C169 B.n51 VSUBS 0.010839f
C170 B.n52 VSUBS 0.027831f
C171 B.n53 VSUBS 0.010839f
C172 B.n54 VSUBS 0.010839f
C173 B.n55 VSUBS 0.010839f
C174 B.n56 VSUBS 0.010839f
C175 B.n57 VSUBS 0.010839f
C176 B.n58 VSUBS 0.010839f
C177 B.n59 VSUBS 0.010839f
C178 B.n60 VSUBS 0.010839f
C179 B.n61 VSUBS 0.010839f
C180 B.n62 VSUBS 0.010839f
C181 B.n63 VSUBS 0.010839f
C182 B.n64 VSUBS 0.010839f
C183 B.n65 VSUBS 0.010839f
C184 B.n66 VSUBS 0.010839f
C185 B.n67 VSUBS 0.010839f
C186 B.n68 VSUBS 0.010839f
C187 B.n69 VSUBS 0.010839f
C188 B.n70 VSUBS 0.010839f
C189 B.n71 VSUBS 0.010839f
C190 B.n72 VSUBS 0.010839f
C191 B.n73 VSUBS 0.010839f
C192 B.n74 VSUBS 0.010839f
C193 B.n75 VSUBS 0.010839f
C194 B.n76 VSUBS 0.010839f
C195 B.n77 VSUBS 0.010839f
C196 B.n78 VSUBS 0.010839f
C197 B.n79 VSUBS 0.010839f
C198 B.n80 VSUBS 0.010839f
C199 B.n81 VSUBS 0.010839f
C200 B.n82 VSUBS 0.010839f
C201 B.n83 VSUBS 0.010839f
C202 B.n84 VSUBS 0.010839f
C203 B.n85 VSUBS 0.010839f
C204 B.n86 VSUBS 0.010839f
C205 B.n87 VSUBS 0.010839f
C206 B.n88 VSUBS 0.010839f
C207 B.n89 VSUBS 0.010839f
C208 B.n90 VSUBS 0.010839f
C209 B.n91 VSUBS 0.010839f
C210 B.n92 VSUBS 0.010839f
C211 B.n93 VSUBS 0.010839f
C212 B.n94 VSUBS 0.010839f
C213 B.n95 VSUBS 0.010839f
C214 B.n96 VSUBS 0.010839f
C215 B.n97 VSUBS 0.010839f
C216 B.n98 VSUBS 0.010839f
C217 B.n99 VSUBS 0.010839f
C218 B.n100 VSUBS 0.010839f
C219 B.n101 VSUBS 0.010839f
C220 B.n102 VSUBS 0.010839f
C221 B.n103 VSUBS 0.010839f
C222 B.n104 VSUBS 0.010839f
C223 B.n105 VSUBS 0.010839f
C224 B.n106 VSUBS 0.010839f
C225 B.n107 VSUBS 0.010839f
C226 B.n108 VSUBS 0.010839f
C227 B.n109 VSUBS 0.010839f
C228 B.n110 VSUBS 0.010839f
C229 B.n111 VSUBS 0.026681f
C230 B.n112 VSUBS 0.010839f
C231 B.n113 VSUBS 0.010839f
C232 B.n114 VSUBS 0.010839f
C233 B.n115 VSUBS 0.010839f
C234 B.n116 VSUBS 0.010839f
C235 B.n117 VSUBS 0.010839f
C236 B.t2 VSUBS 0.069458f
C237 B.t1 VSUBS 0.091499f
C238 B.t0 VSUBS 0.489647f
C239 B.n118 VSUBS 0.117628f
C240 B.n119 VSUBS 0.09404f
C241 B.n120 VSUBS 0.010839f
C242 B.n121 VSUBS 0.010839f
C243 B.n122 VSUBS 0.010839f
C244 B.n123 VSUBS 0.010839f
C245 B.n124 VSUBS 0.006057f
C246 B.n125 VSUBS 0.010839f
C247 B.n126 VSUBS 0.010839f
C248 B.n127 VSUBS 0.010839f
C249 B.n128 VSUBS 0.010839f
C250 B.n129 VSUBS 0.010839f
C251 B.n130 VSUBS 0.027831f
C252 B.n131 VSUBS 0.010839f
C253 B.n132 VSUBS 0.010839f
C254 B.n133 VSUBS 0.010839f
C255 B.n134 VSUBS 0.010839f
C256 B.n135 VSUBS 0.010839f
C257 B.n136 VSUBS 0.010839f
C258 B.n137 VSUBS 0.010839f
C259 B.n138 VSUBS 0.010839f
C260 B.n139 VSUBS 0.010839f
C261 B.n140 VSUBS 0.010839f
C262 B.n141 VSUBS 0.010839f
C263 B.n142 VSUBS 0.010839f
C264 B.n143 VSUBS 0.010839f
C265 B.n144 VSUBS 0.010839f
C266 B.n145 VSUBS 0.010839f
C267 B.n146 VSUBS 0.010839f
C268 B.n147 VSUBS 0.010839f
C269 B.n148 VSUBS 0.010839f
C270 B.n149 VSUBS 0.010839f
C271 B.n150 VSUBS 0.010839f
C272 B.n151 VSUBS 0.010839f
C273 B.n152 VSUBS 0.010839f
C274 B.n153 VSUBS 0.010839f
C275 B.n154 VSUBS 0.010839f
C276 B.n155 VSUBS 0.010839f
C277 B.n156 VSUBS 0.010839f
C278 B.n157 VSUBS 0.010839f
C279 B.n158 VSUBS 0.010839f
C280 B.n159 VSUBS 0.010839f
C281 B.n160 VSUBS 0.010839f
C282 B.n161 VSUBS 0.010839f
C283 B.n162 VSUBS 0.010839f
C284 B.n163 VSUBS 0.010839f
C285 B.n164 VSUBS 0.010839f
C286 B.n165 VSUBS 0.010839f
C287 B.n166 VSUBS 0.010839f
C288 B.n167 VSUBS 0.010839f
C289 B.n168 VSUBS 0.010839f
C290 B.n169 VSUBS 0.010839f
C291 B.n170 VSUBS 0.010839f
C292 B.n171 VSUBS 0.010839f
C293 B.n172 VSUBS 0.010839f
C294 B.n173 VSUBS 0.010839f
C295 B.n174 VSUBS 0.010839f
C296 B.n175 VSUBS 0.010839f
C297 B.n176 VSUBS 0.010839f
C298 B.n177 VSUBS 0.010839f
C299 B.n178 VSUBS 0.010839f
C300 B.n179 VSUBS 0.010839f
C301 B.n180 VSUBS 0.010839f
C302 B.n181 VSUBS 0.010839f
C303 B.n182 VSUBS 0.010839f
C304 B.n183 VSUBS 0.010839f
C305 B.n184 VSUBS 0.010839f
C306 B.n185 VSUBS 0.010839f
C307 B.n186 VSUBS 0.010839f
C308 B.n187 VSUBS 0.010839f
C309 B.n188 VSUBS 0.010839f
C310 B.n189 VSUBS 0.010839f
C311 B.n190 VSUBS 0.010839f
C312 B.n191 VSUBS 0.010839f
C313 B.n192 VSUBS 0.010839f
C314 B.n193 VSUBS 0.010839f
C315 B.n194 VSUBS 0.010839f
C316 B.n195 VSUBS 0.010839f
C317 B.n196 VSUBS 0.010839f
C318 B.n197 VSUBS 0.010839f
C319 B.n198 VSUBS 0.010839f
C320 B.n199 VSUBS 0.010839f
C321 B.n200 VSUBS 0.010839f
C322 B.n201 VSUBS 0.010839f
C323 B.n202 VSUBS 0.010839f
C324 B.n203 VSUBS 0.010839f
C325 B.n204 VSUBS 0.010839f
C326 B.n205 VSUBS 0.010839f
C327 B.n206 VSUBS 0.010839f
C328 B.n207 VSUBS 0.010839f
C329 B.n208 VSUBS 0.010839f
C330 B.n209 VSUBS 0.010839f
C331 B.n210 VSUBS 0.010839f
C332 B.n211 VSUBS 0.010839f
C333 B.n212 VSUBS 0.010839f
C334 B.n213 VSUBS 0.010839f
C335 B.n214 VSUBS 0.010839f
C336 B.n215 VSUBS 0.010839f
C337 B.n216 VSUBS 0.010839f
C338 B.n217 VSUBS 0.010839f
C339 B.n218 VSUBS 0.010839f
C340 B.n219 VSUBS 0.010839f
C341 B.n220 VSUBS 0.010839f
C342 B.n221 VSUBS 0.010839f
C343 B.n222 VSUBS 0.010839f
C344 B.n223 VSUBS 0.010839f
C345 B.n224 VSUBS 0.010839f
C346 B.n225 VSUBS 0.010839f
C347 B.n226 VSUBS 0.010839f
C348 B.n227 VSUBS 0.010839f
C349 B.n228 VSUBS 0.010839f
C350 B.n229 VSUBS 0.010839f
C351 B.n230 VSUBS 0.010839f
C352 B.n231 VSUBS 0.010839f
C353 B.n232 VSUBS 0.010839f
C354 B.n233 VSUBS 0.010839f
C355 B.n234 VSUBS 0.010839f
C356 B.n235 VSUBS 0.010839f
C357 B.n236 VSUBS 0.010839f
C358 B.n237 VSUBS 0.010839f
C359 B.n238 VSUBS 0.010839f
C360 B.n239 VSUBS 0.010839f
C361 B.n240 VSUBS 0.010839f
C362 B.n241 VSUBS 0.010839f
C363 B.n242 VSUBS 0.010839f
C364 B.n243 VSUBS 0.026681f
C365 B.n244 VSUBS 0.026681f
C366 B.n245 VSUBS 0.027831f
C367 B.n246 VSUBS 0.010839f
C368 B.n247 VSUBS 0.010839f
C369 B.n248 VSUBS 0.010839f
C370 B.n249 VSUBS 0.010839f
C371 B.n250 VSUBS 0.010839f
C372 B.n251 VSUBS 0.010839f
C373 B.n252 VSUBS 0.010839f
C374 B.n253 VSUBS 0.010839f
C375 B.n254 VSUBS 0.010839f
C376 B.n255 VSUBS 0.010839f
C377 B.n256 VSUBS 0.010839f
C378 B.n257 VSUBS 0.010839f
C379 B.n258 VSUBS 0.010839f
C380 B.n259 VSUBS 0.010839f
C381 B.n260 VSUBS 0.010839f
C382 B.t8 VSUBS 0.069458f
C383 B.t7 VSUBS 0.091499f
C384 B.t6 VSUBS 0.489647f
C385 B.n261 VSUBS 0.117628f
C386 B.n262 VSUBS 0.09404f
C387 B.n263 VSUBS 0.025112f
C388 B.n264 VSUBS 0.010201f
C389 B.n265 VSUBS 0.010839f
C390 B.n266 VSUBS 0.010839f
C391 B.n267 VSUBS 0.010839f
C392 B.n268 VSUBS 0.010839f
C393 B.n269 VSUBS 0.010839f
C394 B.n270 VSUBS 0.010839f
C395 B.n271 VSUBS 0.010839f
C396 B.n272 VSUBS 0.010839f
C397 B.n273 VSUBS 0.010839f
C398 B.n274 VSUBS 0.010839f
C399 B.n275 VSUBS 0.010839f
C400 B.n276 VSUBS 0.010839f
C401 B.n277 VSUBS 0.010839f
C402 B.n278 VSUBS 0.010839f
C403 B.n279 VSUBS 0.010839f
C404 B.n280 VSUBS 0.006057f
C405 B.n281 VSUBS 0.025112f
C406 B.n282 VSUBS 0.010201f
C407 B.n283 VSUBS 0.010839f
C408 B.n284 VSUBS 0.010839f
C409 B.n285 VSUBS 0.010839f
C410 B.n286 VSUBS 0.010839f
C411 B.n287 VSUBS 0.010839f
C412 B.n288 VSUBS 0.010839f
C413 B.n289 VSUBS 0.010839f
C414 B.n290 VSUBS 0.010839f
C415 B.n291 VSUBS 0.010839f
C416 B.n292 VSUBS 0.010839f
C417 B.n293 VSUBS 0.010839f
C418 B.n294 VSUBS 0.010839f
C419 B.n295 VSUBS 0.010839f
C420 B.n296 VSUBS 0.010839f
C421 B.n297 VSUBS 0.010839f
C422 B.n298 VSUBS 0.027831f
C423 B.n299 VSUBS 0.026681f
C424 B.n300 VSUBS 0.027831f
C425 B.n301 VSUBS 0.010839f
C426 B.n302 VSUBS 0.010839f
C427 B.n303 VSUBS 0.010839f
C428 B.n304 VSUBS 0.010839f
C429 B.n305 VSUBS 0.010839f
C430 B.n306 VSUBS 0.010839f
C431 B.n307 VSUBS 0.010839f
C432 B.n308 VSUBS 0.010839f
C433 B.n309 VSUBS 0.010839f
C434 B.n310 VSUBS 0.010839f
C435 B.n311 VSUBS 0.010839f
C436 B.n312 VSUBS 0.010839f
C437 B.n313 VSUBS 0.010839f
C438 B.n314 VSUBS 0.010839f
C439 B.n315 VSUBS 0.010839f
C440 B.n316 VSUBS 0.010839f
C441 B.n317 VSUBS 0.010839f
C442 B.n318 VSUBS 0.010839f
C443 B.n319 VSUBS 0.010839f
C444 B.n320 VSUBS 0.010839f
C445 B.n321 VSUBS 0.010839f
C446 B.n322 VSUBS 0.010839f
C447 B.n323 VSUBS 0.010839f
C448 B.n324 VSUBS 0.010839f
C449 B.n325 VSUBS 0.010839f
C450 B.n326 VSUBS 0.010839f
C451 B.n327 VSUBS 0.010839f
C452 B.n328 VSUBS 0.010839f
C453 B.n329 VSUBS 0.010839f
C454 B.n330 VSUBS 0.010839f
C455 B.n331 VSUBS 0.010839f
C456 B.n332 VSUBS 0.010839f
C457 B.n333 VSUBS 0.010839f
C458 B.n334 VSUBS 0.010839f
C459 B.n335 VSUBS 0.010839f
C460 B.n336 VSUBS 0.010839f
C461 B.n337 VSUBS 0.010839f
C462 B.n338 VSUBS 0.010839f
C463 B.n339 VSUBS 0.010839f
C464 B.n340 VSUBS 0.010839f
C465 B.n341 VSUBS 0.010839f
C466 B.n342 VSUBS 0.010839f
C467 B.n343 VSUBS 0.010839f
C468 B.n344 VSUBS 0.010839f
C469 B.n345 VSUBS 0.010839f
C470 B.n346 VSUBS 0.010839f
C471 B.n347 VSUBS 0.010839f
C472 B.n348 VSUBS 0.010839f
C473 B.n349 VSUBS 0.010839f
C474 B.n350 VSUBS 0.010839f
C475 B.n351 VSUBS 0.010839f
C476 B.n352 VSUBS 0.010839f
C477 B.n353 VSUBS 0.010839f
C478 B.n354 VSUBS 0.010839f
C479 B.n355 VSUBS 0.010839f
C480 B.n356 VSUBS 0.010839f
C481 B.n357 VSUBS 0.010839f
C482 B.n358 VSUBS 0.010839f
C483 B.n359 VSUBS 0.010839f
C484 B.n360 VSUBS 0.010839f
C485 B.n361 VSUBS 0.010839f
C486 B.n362 VSUBS 0.010839f
C487 B.n363 VSUBS 0.010839f
C488 B.n364 VSUBS 0.010839f
C489 B.n365 VSUBS 0.010839f
C490 B.n366 VSUBS 0.010839f
C491 B.n367 VSUBS 0.010839f
C492 B.n368 VSUBS 0.010839f
C493 B.n369 VSUBS 0.010839f
C494 B.n370 VSUBS 0.010839f
C495 B.n371 VSUBS 0.010839f
C496 B.n372 VSUBS 0.010839f
C497 B.n373 VSUBS 0.010839f
C498 B.n374 VSUBS 0.010839f
C499 B.n375 VSUBS 0.010839f
C500 B.n376 VSUBS 0.010839f
C501 B.n377 VSUBS 0.010839f
C502 B.n378 VSUBS 0.010839f
C503 B.n379 VSUBS 0.010839f
C504 B.n380 VSUBS 0.010839f
C505 B.n381 VSUBS 0.010839f
C506 B.n382 VSUBS 0.010839f
C507 B.n383 VSUBS 0.010839f
C508 B.n384 VSUBS 0.010839f
C509 B.n385 VSUBS 0.010839f
C510 B.n386 VSUBS 0.010839f
C511 B.n387 VSUBS 0.010839f
C512 B.n388 VSUBS 0.010839f
C513 B.n389 VSUBS 0.010839f
C514 B.n390 VSUBS 0.010839f
C515 B.n391 VSUBS 0.010839f
C516 B.n392 VSUBS 0.010839f
C517 B.n393 VSUBS 0.010839f
C518 B.n394 VSUBS 0.010839f
C519 B.n395 VSUBS 0.010839f
C520 B.n396 VSUBS 0.010839f
C521 B.n397 VSUBS 0.010839f
C522 B.n398 VSUBS 0.010839f
C523 B.n399 VSUBS 0.010839f
C524 B.n400 VSUBS 0.010839f
C525 B.n401 VSUBS 0.010839f
C526 B.n402 VSUBS 0.010839f
C527 B.n403 VSUBS 0.010839f
C528 B.n404 VSUBS 0.010839f
C529 B.n405 VSUBS 0.010839f
C530 B.n406 VSUBS 0.010839f
C531 B.n407 VSUBS 0.010839f
C532 B.n408 VSUBS 0.010839f
C533 B.n409 VSUBS 0.010839f
C534 B.n410 VSUBS 0.010839f
C535 B.n411 VSUBS 0.010839f
C536 B.n412 VSUBS 0.010839f
C537 B.n413 VSUBS 0.010839f
C538 B.n414 VSUBS 0.010839f
C539 B.n415 VSUBS 0.010839f
C540 B.n416 VSUBS 0.010839f
C541 B.n417 VSUBS 0.010839f
C542 B.n418 VSUBS 0.010839f
C543 B.n419 VSUBS 0.010839f
C544 B.n420 VSUBS 0.010839f
C545 B.n421 VSUBS 0.010839f
C546 B.n422 VSUBS 0.010839f
C547 B.n423 VSUBS 0.010839f
C548 B.n424 VSUBS 0.010839f
C549 B.n425 VSUBS 0.010839f
C550 B.n426 VSUBS 0.010839f
C551 B.n427 VSUBS 0.010839f
C552 B.n428 VSUBS 0.010839f
C553 B.n429 VSUBS 0.010839f
C554 B.n430 VSUBS 0.010839f
C555 B.n431 VSUBS 0.010839f
C556 B.n432 VSUBS 0.010839f
C557 B.n433 VSUBS 0.010839f
C558 B.n434 VSUBS 0.010839f
C559 B.n435 VSUBS 0.010839f
C560 B.n436 VSUBS 0.010839f
C561 B.n437 VSUBS 0.010839f
C562 B.n438 VSUBS 0.010839f
C563 B.n439 VSUBS 0.010839f
C564 B.n440 VSUBS 0.010839f
C565 B.n441 VSUBS 0.010839f
C566 B.n442 VSUBS 0.010839f
C567 B.n443 VSUBS 0.010839f
C568 B.n444 VSUBS 0.010839f
C569 B.n445 VSUBS 0.010839f
C570 B.n446 VSUBS 0.010839f
C571 B.n447 VSUBS 0.010839f
C572 B.n448 VSUBS 0.010839f
C573 B.n449 VSUBS 0.010839f
C574 B.n450 VSUBS 0.010839f
C575 B.n451 VSUBS 0.010839f
C576 B.n452 VSUBS 0.010839f
C577 B.n453 VSUBS 0.010839f
C578 B.n454 VSUBS 0.010839f
C579 B.n455 VSUBS 0.010839f
C580 B.n456 VSUBS 0.010839f
C581 B.n457 VSUBS 0.010839f
C582 B.n458 VSUBS 0.010839f
C583 B.n459 VSUBS 0.010839f
C584 B.n460 VSUBS 0.010839f
C585 B.n461 VSUBS 0.010839f
C586 B.n462 VSUBS 0.010839f
C587 B.n463 VSUBS 0.010839f
C588 B.n464 VSUBS 0.010839f
C589 B.n465 VSUBS 0.010839f
C590 B.n466 VSUBS 0.010839f
C591 B.n467 VSUBS 0.010839f
C592 B.n468 VSUBS 0.010839f
C593 B.n469 VSUBS 0.010839f
C594 B.n470 VSUBS 0.010839f
C595 B.n471 VSUBS 0.010839f
C596 B.n472 VSUBS 0.010839f
C597 B.n473 VSUBS 0.010839f
C598 B.n474 VSUBS 0.010839f
C599 B.n475 VSUBS 0.026681f
C600 B.n476 VSUBS 0.026681f
C601 B.n477 VSUBS 0.027831f
C602 B.n478 VSUBS 0.010839f
C603 B.n479 VSUBS 0.010839f
C604 B.n480 VSUBS 0.010839f
C605 B.n481 VSUBS 0.010839f
C606 B.n482 VSUBS 0.010839f
C607 B.n483 VSUBS 0.010839f
C608 B.n484 VSUBS 0.010839f
C609 B.n485 VSUBS 0.010839f
C610 B.n486 VSUBS 0.010839f
C611 B.n487 VSUBS 0.010839f
C612 B.n488 VSUBS 0.010839f
C613 B.n489 VSUBS 0.010839f
C614 B.n490 VSUBS 0.010839f
C615 B.n491 VSUBS 0.010839f
C616 B.n492 VSUBS 0.010839f
C617 B.n493 VSUBS 0.010201f
C618 B.n494 VSUBS 0.010839f
C619 B.n495 VSUBS 0.010839f
C620 B.n496 VSUBS 0.006057f
C621 B.n497 VSUBS 0.010839f
C622 B.n498 VSUBS 0.010839f
C623 B.n499 VSUBS 0.010839f
C624 B.n500 VSUBS 0.010839f
C625 B.n501 VSUBS 0.010839f
C626 B.n502 VSUBS 0.010839f
C627 B.n503 VSUBS 0.010839f
C628 B.n504 VSUBS 0.010839f
C629 B.n505 VSUBS 0.010839f
C630 B.n506 VSUBS 0.010839f
C631 B.n507 VSUBS 0.010839f
C632 B.n508 VSUBS 0.010839f
C633 B.n509 VSUBS 0.006057f
C634 B.n510 VSUBS 0.025112f
C635 B.n511 VSUBS 0.010201f
C636 B.n512 VSUBS 0.010839f
C637 B.n513 VSUBS 0.010839f
C638 B.n514 VSUBS 0.010839f
C639 B.n515 VSUBS 0.010839f
C640 B.n516 VSUBS 0.010839f
C641 B.n517 VSUBS 0.010839f
C642 B.n518 VSUBS 0.010839f
C643 B.n519 VSUBS 0.010839f
C644 B.n520 VSUBS 0.010839f
C645 B.n521 VSUBS 0.010839f
C646 B.n522 VSUBS 0.010839f
C647 B.n523 VSUBS 0.010839f
C648 B.n524 VSUBS 0.010839f
C649 B.n525 VSUBS 0.010839f
C650 B.n526 VSUBS 0.010839f
C651 B.n527 VSUBS 0.010839f
C652 B.n528 VSUBS 0.027831f
C653 B.n529 VSUBS 0.026681f
C654 B.n530 VSUBS 0.026681f
C655 B.n531 VSUBS 0.010839f
C656 B.n532 VSUBS 0.010839f
C657 B.n533 VSUBS 0.010839f
C658 B.n534 VSUBS 0.010839f
C659 B.n535 VSUBS 0.010839f
C660 B.n536 VSUBS 0.010839f
C661 B.n537 VSUBS 0.010839f
C662 B.n538 VSUBS 0.010839f
C663 B.n539 VSUBS 0.010839f
C664 B.n540 VSUBS 0.010839f
C665 B.n541 VSUBS 0.010839f
C666 B.n542 VSUBS 0.010839f
C667 B.n543 VSUBS 0.010839f
C668 B.n544 VSUBS 0.010839f
C669 B.n545 VSUBS 0.010839f
C670 B.n546 VSUBS 0.010839f
C671 B.n547 VSUBS 0.010839f
C672 B.n548 VSUBS 0.010839f
C673 B.n549 VSUBS 0.010839f
C674 B.n550 VSUBS 0.010839f
C675 B.n551 VSUBS 0.010839f
C676 B.n552 VSUBS 0.010839f
C677 B.n553 VSUBS 0.010839f
C678 B.n554 VSUBS 0.010839f
C679 B.n555 VSUBS 0.010839f
C680 B.n556 VSUBS 0.010839f
C681 B.n557 VSUBS 0.010839f
C682 B.n558 VSUBS 0.010839f
C683 B.n559 VSUBS 0.010839f
C684 B.n560 VSUBS 0.010839f
C685 B.n561 VSUBS 0.010839f
C686 B.n562 VSUBS 0.010839f
C687 B.n563 VSUBS 0.010839f
C688 B.n564 VSUBS 0.010839f
C689 B.n565 VSUBS 0.010839f
C690 B.n566 VSUBS 0.010839f
C691 B.n567 VSUBS 0.010839f
C692 B.n568 VSUBS 0.010839f
C693 B.n569 VSUBS 0.010839f
C694 B.n570 VSUBS 0.010839f
C695 B.n571 VSUBS 0.010839f
C696 B.n572 VSUBS 0.010839f
C697 B.n573 VSUBS 0.010839f
C698 B.n574 VSUBS 0.010839f
C699 B.n575 VSUBS 0.010839f
C700 B.n576 VSUBS 0.010839f
C701 B.n577 VSUBS 0.010839f
C702 B.n578 VSUBS 0.010839f
C703 B.n579 VSUBS 0.010839f
C704 B.n580 VSUBS 0.010839f
C705 B.n581 VSUBS 0.010839f
C706 B.n582 VSUBS 0.010839f
C707 B.n583 VSUBS 0.010839f
C708 B.n584 VSUBS 0.010839f
C709 B.n585 VSUBS 0.010839f
C710 B.n586 VSUBS 0.010839f
C711 B.n587 VSUBS 0.010839f
C712 B.n588 VSUBS 0.010839f
C713 B.n589 VSUBS 0.010839f
C714 B.n590 VSUBS 0.010839f
C715 B.n591 VSUBS 0.010839f
C716 B.n592 VSUBS 0.010839f
C717 B.n593 VSUBS 0.010839f
C718 B.n594 VSUBS 0.010839f
C719 B.n595 VSUBS 0.010839f
C720 B.n596 VSUBS 0.010839f
C721 B.n597 VSUBS 0.010839f
C722 B.n598 VSUBS 0.010839f
C723 B.n599 VSUBS 0.010839f
C724 B.n600 VSUBS 0.010839f
C725 B.n601 VSUBS 0.010839f
C726 B.n602 VSUBS 0.010839f
C727 B.n603 VSUBS 0.010839f
C728 B.n604 VSUBS 0.010839f
C729 B.n605 VSUBS 0.010839f
C730 B.n606 VSUBS 0.010839f
C731 B.n607 VSUBS 0.010839f
C732 B.n608 VSUBS 0.010839f
C733 B.n609 VSUBS 0.010839f
C734 B.n610 VSUBS 0.010839f
C735 B.n611 VSUBS 0.010839f
C736 B.n612 VSUBS 0.010839f
C737 B.n613 VSUBS 0.010839f
C738 B.n614 VSUBS 0.010839f
C739 B.n615 VSUBS 0.014144f
C740 B.n616 VSUBS 0.015067f
C741 B.n617 VSUBS 0.029962f
C742 VDD1.t5 VSUBS 0.051197f
C743 VDD1.t7 VSUBS 0.051197f
C744 VDD1.n0 VSUBS 0.239737f
C745 VDD1.t6 VSUBS 0.051197f
C746 VDD1.t2 VSUBS 0.051197f
C747 VDD1.n1 VSUBS 0.239122f
C748 VDD1.t0 VSUBS 0.051197f
C749 VDD1.t1 VSUBS 0.051197f
C750 VDD1.n2 VSUBS 0.239122f
C751 VDD1.n3 VSUBS 3.96361f
C752 VDD1.t3 VSUBS 0.051197f
C753 VDD1.t4 VSUBS 0.051197f
C754 VDD1.n4 VSUBS 0.232566f
C755 VDD1.n5 VSUBS 3.07895f
C756 VTAIL.t6 VSUBS 0.059447f
C757 VTAIL.t3 VSUBS 0.059447f
C758 VTAIL.n0 VSUBS 0.228862f
C759 VTAIL.n1 VSUBS 0.735867f
C760 VTAIL.t0 VSUBS 0.360276f
C761 VTAIL.n2 VSUBS 0.815019f
C762 VTAIL.t12 VSUBS 0.360276f
C763 VTAIL.n3 VSUBS 0.815019f
C764 VTAIL.t13 VSUBS 0.059447f
C765 VTAIL.t9 VSUBS 0.059447f
C766 VTAIL.n4 VSUBS 0.228862f
C767 VTAIL.n5 VSUBS 1.07797f
C768 VTAIL.t14 VSUBS 0.360276f
C769 VTAIL.n6 VSUBS 1.8137f
C770 VTAIL.t4 VSUBS 0.360277f
C771 VTAIL.n7 VSUBS 1.8137f
C772 VTAIL.t7 VSUBS 0.059447f
C773 VTAIL.t2 VSUBS 0.059447f
C774 VTAIL.n8 VSUBS 0.228863f
C775 VTAIL.n9 VSUBS 1.07797f
C776 VTAIL.t1 VSUBS 0.360277f
C777 VTAIL.n10 VSUBS 0.815017f
C778 VTAIL.t8 VSUBS 0.360277f
C779 VTAIL.n11 VSUBS 0.815017f
C780 VTAIL.t10 VSUBS 0.059447f
C781 VTAIL.t11 VSUBS 0.059447f
C782 VTAIL.n12 VSUBS 0.228863f
C783 VTAIL.n13 VSUBS 1.07797f
C784 VTAIL.t15 VSUBS 0.360276f
C785 VTAIL.n14 VSUBS 1.8137f
C786 VTAIL.t5 VSUBS 0.360276f
C787 VTAIL.n15 VSUBS 1.80686f
C788 VP.t6 VSUBS 0.875274f
C789 VP.n0 VSUBS 0.640862f
C790 VP.n1 VSUBS 0.058161f
C791 VP.n2 VSUBS 0.075481f
C792 VP.n3 VSUBS 0.058161f
C793 VP.t7 VSUBS 0.875274f
C794 VP.n4 VSUBS 0.401871f
C795 VP.n5 VSUBS 0.058161f
C796 VP.n6 VSUBS 0.085275f
C797 VP.n7 VSUBS 0.058161f
C798 VP.t5 VSUBS 0.875274f
C799 VP.n8 VSUBS 0.108941f
C800 VP.n9 VSUBS 0.058161f
C801 VP.n10 VSUBS 0.108941f
C802 VP.t3 VSUBS 0.875274f
C803 VP.n11 VSUBS 0.640862f
C804 VP.n12 VSUBS 0.058161f
C805 VP.n13 VSUBS 0.075481f
C806 VP.n14 VSUBS 0.058161f
C807 VP.t4 VSUBS 0.875274f
C808 VP.n15 VSUBS 0.401871f
C809 VP.n16 VSUBS 0.058161f
C810 VP.n17 VSUBS 0.085275f
C811 VP.n18 VSUBS 0.664159f
C812 VP.t0 VSUBS 0.875274f
C813 VP.t2 VSUBS 1.4292f
C814 VP.n19 VSUBS 0.607107f
C815 VP.n20 VSUBS 0.617736f
C816 VP.n21 VSUBS 0.105714f
C817 VP.n22 VSUBS 0.108941f
C818 VP.n23 VSUBS 0.058161f
C819 VP.n24 VSUBS 0.058161f
C820 VP.n25 VSUBS 0.058161f
C821 VP.n26 VSUBS 0.085275f
C822 VP.n27 VSUBS 0.108941f
C823 VP.n28 VSUBS 0.105714f
C824 VP.n29 VSUBS 0.058161f
C825 VP.n30 VSUBS 0.058161f
C826 VP.n31 VSUBS 0.05838f
C827 VP.n32 VSUBS 0.108941f
C828 VP.n33 VSUBS 0.108941f
C829 VP.n34 VSUBS 0.058161f
C830 VP.n35 VSUBS 0.058161f
C831 VP.n36 VSUBS 0.058161f
C832 VP.n37 VSUBS 0.095068f
C833 VP.n38 VSUBS 0.108941f
C834 VP.n39 VSUBS 0.09926f
C835 VP.n40 VSUBS 0.093886f
C836 VP.n41 VSUBS 2.902f
C837 VP.n42 VSUBS 2.94742f
C838 VP.t1 VSUBS 0.875274f
C839 VP.n43 VSUBS 0.640862f
C840 VP.n44 VSUBS 0.09926f
C841 VP.n45 VSUBS 0.093886f
C842 VP.n46 VSUBS 0.058161f
C843 VP.n47 VSUBS 0.058161f
C844 VP.n48 VSUBS 0.095068f
C845 VP.n49 VSUBS 0.075481f
C846 VP.n50 VSUBS 0.108941f
C847 VP.n51 VSUBS 0.058161f
C848 VP.n52 VSUBS 0.058161f
C849 VP.n53 VSUBS 0.058161f
C850 VP.n54 VSUBS 0.05838f
C851 VP.n55 VSUBS 0.401871f
C852 VP.n56 VSUBS 0.105714f
C853 VP.n57 VSUBS 0.108941f
C854 VP.n58 VSUBS 0.058161f
C855 VP.n59 VSUBS 0.058161f
C856 VP.n60 VSUBS 0.058161f
C857 VP.n61 VSUBS 0.085275f
C858 VP.n62 VSUBS 0.108941f
C859 VP.n63 VSUBS 0.105714f
C860 VP.n64 VSUBS 0.058161f
C861 VP.n65 VSUBS 0.058161f
C862 VP.n66 VSUBS 0.05838f
C863 VP.n67 VSUBS 0.108941f
C864 VP.n68 VSUBS 0.108941f
C865 VP.n69 VSUBS 0.058161f
C866 VP.n70 VSUBS 0.058161f
C867 VP.n71 VSUBS 0.058161f
C868 VP.n72 VSUBS 0.095068f
C869 VP.n73 VSUBS 0.108941f
C870 VP.n74 VSUBS 0.09926f
C871 VP.n75 VSUBS 0.093886f
C872 VP.n76 VSUBS 0.123061f
.ends

