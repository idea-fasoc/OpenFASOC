* NGSPICE file created from diff_pair_sample_1127.ext - technology: sky130A

.subckt diff_pair_sample_1127 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VN.t0 VDD2.t4 w_n3220_n1646# sky130_fd_pr__pfet_01v8 ad=1.3221 pd=7.56 as=0.55935 ps=3.72 w=3.39 l=1.92
X1 VDD1.t7 VP.t0 VTAIL.t4 w_n3220_n1646# sky130_fd_pr__pfet_01v8 ad=0.55935 pd=3.72 as=1.3221 ps=7.56 w=3.39 l=1.92
X2 B.t11 B.t9 B.t10 w_n3220_n1646# sky130_fd_pr__pfet_01v8 ad=1.3221 pd=7.56 as=0 ps=0 w=3.39 l=1.92
X3 B.t8 B.t6 B.t7 w_n3220_n1646# sky130_fd_pr__pfet_01v8 ad=1.3221 pd=7.56 as=0 ps=0 w=3.39 l=1.92
X4 VTAIL.t14 VN.t1 VDD2.t5 w_n3220_n1646# sky130_fd_pr__pfet_01v8 ad=0.55935 pd=3.72 as=0.55935 ps=3.72 w=3.39 l=1.92
X5 VTAIL.t3 VP.t1 VDD1.t6 w_n3220_n1646# sky130_fd_pr__pfet_01v8 ad=1.3221 pd=7.56 as=0.55935 ps=3.72 w=3.39 l=1.92
X6 VTAIL.t7 VP.t2 VDD1.t5 w_n3220_n1646# sky130_fd_pr__pfet_01v8 ad=0.55935 pd=3.72 as=0.55935 ps=3.72 w=3.39 l=1.92
X7 VTAIL.t5 VP.t3 VDD1.t4 w_n3220_n1646# sky130_fd_pr__pfet_01v8 ad=1.3221 pd=7.56 as=0.55935 ps=3.72 w=3.39 l=1.92
X8 VTAIL.t13 VN.t2 VDD2.t6 w_n3220_n1646# sky130_fd_pr__pfet_01v8 ad=1.3221 pd=7.56 as=0.55935 ps=3.72 w=3.39 l=1.92
X9 VDD2.t3 VN.t3 VTAIL.t12 w_n3220_n1646# sky130_fd_pr__pfet_01v8 ad=0.55935 pd=3.72 as=1.3221 ps=7.56 w=3.39 l=1.92
X10 B.t5 B.t3 B.t4 w_n3220_n1646# sky130_fd_pr__pfet_01v8 ad=1.3221 pd=7.56 as=0 ps=0 w=3.39 l=1.92
X11 VDD2.t1 VN.t4 VTAIL.t11 w_n3220_n1646# sky130_fd_pr__pfet_01v8 ad=0.55935 pd=3.72 as=0.55935 ps=3.72 w=3.39 l=1.92
X12 VTAIL.t1 VP.t4 VDD1.t3 w_n3220_n1646# sky130_fd_pr__pfet_01v8 ad=0.55935 pd=3.72 as=0.55935 ps=3.72 w=3.39 l=1.92
X13 VDD2.t2 VN.t5 VTAIL.t10 w_n3220_n1646# sky130_fd_pr__pfet_01v8 ad=0.55935 pd=3.72 as=1.3221 ps=7.56 w=3.39 l=1.92
X14 VDD1.t2 VP.t5 VTAIL.t2 w_n3220_n1646# sky130_fd_pr__pfet_01v8 ad=0.55935 pd=3.72 as=1.3221 ps=7.56 w=3.39 l=1.92
X15 VDD1.t1 VP.t6 VTAIL.t0 w_n3220_n1646# sky130_fd_pr__pfet_01v8 ad=0.55935 pd=3.72 as=0.55935 ps=3.72 w=3.39 l=1.92
X16 B.t2 B.t0 B.t1 w_n3220_n1646# sky130_fd_pr__pfet_01v8 ad=1.3221 pd=7.56 as=0 ps=0 w=3.39 l=1.92
X17 VDD2.t7 VN.t6 VTAIL.t9 w_n3220_n1646# sky130_fd_pr__pfet_01v8 ad=0.55935 pd=3.72 as=0.55935 ps=3.72 w=3.39 l=1.92
X18 VDD1.t0 VP.t7 VTAIL.t6 w_n3220_n1646# sky130_fd_pr__pfet_01v8 ad=0.55935 pd=3.72 as=0.55935 ps=3.72 w=3.39 l=1.92
X19 VTAIL.t8 VN.t7 VDD2.t0 w_n3220_n1646# sky130_fd_pr__pfet_01v8 ad=0.55935 pd=3.72 as=0.55935 ps=3.72 w=3.39 l=1.92
R0 VN.n43 VN.n23 161.3
R1 VN.n42 VN.n41 161.3
R2 VN.n40 VN.n24 161.3
R3 VN.n39 VN.n38 161.3
R4 VN.n36 VN.n25 161.3
R5 VN.n35 VN.n34 161.3
R6 VN.n33 VN.n26 161.3
R7 VN.n32 VN.n31 161.3
R8 VN.n30 VN.n27 161.3
R9 VN.n20 VN.n0 161.3
R10 VN.n19 VN.n18 161.3
R11 VN.n17 VN.n1 161.3
R12 VN.n16 VN.n15 161.3
R13 VN.n13 VN.n2 161.3
R14 VN.n12 VN.n11 161.3
R15 VN.n10 VN.n3 161.3
R16 VN.n9 VN.n8 161.3
R17 VN.n7 VN.n4 161.3
R18 VN.n22 VN.n21 92.4062
R19 VN.n45 VN.n44 92.4062
R20 VN.n5 VN.t0 72.5661
R21 VN.n28 VN.t3 72.5661
R22 VN.n6 VN.n5 63.4562
R23 VN.n29 VN.n28 63.4562
R24 VN.n19 VN.n1 56.5193
R25 VN.n42 VN.n24 56.5193
R26 VN.n6 VN.t4 42.5521
R27 VN.n14 VN.t1 42.5521
R28 VN.n21 VN.t5 42.5521
R29 VN.n29 VN.t7 42.5521
R30 VN.n37 VN.t6 42.5521
R31 VN.n44 VN.t2 42.5521
R32 VN VN.n45 41.4527
R33 VN.n8 VN.n3 40.4934
R34 VN.n12 VN.n3 40.4934
R35 VN.n31 VN.n26 40.4934
R36 VN.n35 VN.n26 40.4934
R37 VN.n8 VN.n7 24.4675
R38 VN.n13 VN.n12 24.4675
R39 VN.n15 VN.n1 24.4675
R40 VN.n20 VN.n19 24.4675
R41 VN.n31 VN.n30 24.4675
R42 VN.n38 VN.n24 24.4675
R43 VN.n36 VN.n35 24.4675
R44 VN.n43 VN.n42 24.4675
R45 VN.n15 VN.n14 18.3508
R46 VN.n21 VN.n20 18.3508
R47 VN.n38 VN.n37 18.3508
R48 VN.n44 VN.n43 18.3508
R49 VN.n28 VN.n27 13.5379
R50 VN.n5 VN.n4 13.5379
R51 VN.n7 VN.n6 6.11725
R52 VN.n14 VN.n13 6.11725
R53 VN.n30 VN.n29 6.11725
R54 VN.n37 VN.n36 6.11725
R55 VN.n45 VN.n23 0.278367
R56 VN.n22 VN.n0 0.278367
R57 VN.n41 VN.n23 0.189894
R58 VN.n41 VN.n40 0.189894
R59 VN.n40 VN.n39 0.189894
R60 VN.n39 VN.n25 0.189894
R61 VN.n34 VN.n25 0.189894
R62 VN.n34 VN.n33 0.189894
R63 VN.n33 VN.n32 0.189894
R64 VN.n32 VN.n27 0.189894
R65 VN.n9 VN.n4 0.189894
R66 VN.n10 VN.n9 0.189894
R67 VN.n11 VN.n10 0.189894
R68 VN.n11 VN.n2 0.189894
R69 VN.n16 VN.n2 0.189894
R70 VN.n17 VN.n16 0.189894
R71 VN.n18 VN.n17 0.189894
R72 VN.n18 VN.n0 0.189894
R73 VN VN.n22 0.153454
R74 VDD2.n2 VDD2.n1 128.087
R75 VDD2.n2 VDD2.n0 128.087
R76 VDD2 VDD2.n5 128.083
R77 VDD2.n4 VDD2.n3 127.172
R78 VDD2.n4 VDD2.n2 35.3662
R79 VDD2.n5 VDD2.t0 9.589
R80 VDD2.n5 VDD2.t3 9.589
R81 VDD2.n3 VDD2.t6 9.589
R82 VDD2.n3 VDD2.t7 9.589
R83 VDD2.n1 VDD2.t5 9.589
R84 VDD2.n1 VDD2.t2 9.589
R85 VDD2.n0 VDD2.t4 9.589
R86 VDD2.n0 VDD2.t1 9.589
R87 VDD2 VDD2.n4 1.02852
R88 VTAIL.n130 VTAIL.n120 756.745
R89 VTAIL.n12 VTAIL.n2 756.745
R90 VTAIL.n28 VTAIL.n18 756.745
R91 VTAIL.n46 VTAIL.n36 756.745
R92 VTAIL.n114 VTAIL.n104 756.745
R93 VTAIL.n96 VTAIL.n86 756.745
R94 VTAIL.n80 VTAIL.n70 756.745
R95 VTAIL.n62 VTAIL.n52 756.745
R96 VTAIL.n124 VTAIL.n123 585
R97 VTAIL.n129 VTAIL.n128 585
R98 VTAIL.n131 VTAIL.n130 585
R99 VTAIL.n6 VTAIL.n5 585
R100 VTAIL.n11 VTAIL.n10 585
R101 VTAIL.n13 VTAIL.n12 585
R102 VTAIL.n22 VTAIL.n21 585
R103 VTAIL.n27 VTAIL.n26 585
R104 VTAIL.n29 VTAIL.n28 585
R105 VTAIL.n40 VTAIL.n39 585
R106 VTAIL.n45 VTAIL.n44 585
R107 VTAIL.n47 VTAIL.n46 585
R108 VTAIL.n115 VTAIL.n114 585
R109 VTAIL.n113 VTAIL.n112 585
R110 VTAIL.n108 VTAIL.n107 585
R111 VTAIL.n97 VTAIL.n96 585
R112 VTAIL.n95 VTAIL.n94 585
R113 VTAIL.n90 VTAIL.n89 585
R114 VTAIL.n81 VTAIL.n80 585
R115 VTAIL.n79 VTAIL.n78 585
R116 VTAIL.n74 VTAIL.n73 585
R117 VTAIL.n63 VTAIL.n62 585
R118 VTAIL.n61 VTAIL.n60 585
R119 VTAIL.n56 VTAIL.n55 585
R120 VTAIL.n125 VTAIL.t10 338.558
R121 VTAIL.n7 VTAIL.t15 338.558
R122 VTAIL.n23 VTAIL.t2 338.558
R123 VTAIL.n41 VTAIL.t3 338.558
R124 VTAIL.n91 VTAIL.t5 338.558
R125 VTAIL.n75 VTAIL.t12 338.558
R126 VTAIL.n57 VTAIL.t13 338.558
R127 VTAIL.n109 VTAIL.t4 338.558
R128 VTAIL.n129 VTAIL.n123 171.744
R129 VTAIL.n130 VTAIL.n129 171.744
R130 VTAIL.n11 VTAIL.n5 171.744
R131 VTAIL.n12 VTAIL.n11 171.744
R132 VTAIL.n27 VTAIL.n21 171.744
R133 VTAIL.n28 VTAIL.n27 171.744
R134 VTAIL.n45 VTAIL.n39 171.744
R135 VTAIL.n46 VTAIL.n45 171.744
R136 VTAIL.n114 VTAIL.n113 171.744
R137 VTAIL.n113 VTAIL.n107 171.744
R138 VTAIL.n96 VTAIL.n95 171.744
R139 VTAIL.n95 VTAIL.n89 171.744
R140 VTAIL.n80 VTAIL.n79 171.744
R141 VTAIL.n79 VTAIL.n73 171.744
R142 VTAIL.n62 VTAIL.n61 171.744
R143 VTAIL.n61 VTAIL.n55 171.744
R144 VTAIL.n1 VTAIL.n0 110.493
R145 VTAIL.n35 VTAIL.n34 110.493
R146 VTAIL.n103 VTAIL.n102 110.493
R147 VTAIL.n69 VTAIL.n68 110.493
R148 VTAIL.t10 VTAIL.n123 85.8723
R149 VTAIL.t15 VTAIL.n5 85.8723
R150 VTAIL.t2 VTAIL.n21 85.8723
R151 VTAIL.t3 VTAIL.n39 85.8723
R152 VTAIL.t4 VTAIL.n107 85.8723
R153 VTAIL.t5 VTAIL.n89 85.8723
R154 VTAIL.t12 VTAIL.n73 85.8723
R155 VTAIL.t13 VTAIL.n55 85.8723
R156 VTAIL.n135 VTAIL.n134 30.4399
R157 VTAIL.n17 VTAIL.n16 30.4399
R158 VTAIL.n33 VTAIL.n32 30.4399
R159 VTAIL.n51 VTAIL.n50 30.4399
R160 VTAIL.n119 VTAIL.n118 30.4399
R161 VTAIL.n101 VTAIL.n100 30.4399
R162 VTAIL.n85 VTAIL.n84 30.4399
R163 VTAIL.n67 VTAIL.n66 30.4399
R164 VTAIL.n135 VTAIL.n119 17.2289
R165 VTAIL.n67 VTAIL.n51 17.2289
R166 VTAIL.n125 VTAIL.n124 10.6058
R167 VTAIL.n7 VTAIL.n6 10.6058
R168 VTAIL.n23 VTAIL.n22 10.6058
R169 VTAIL.n41 VTAIL.n40 10.6058
R170 VTAIL.n109 VTAIL.n108 10.6058
R171 VTAIL.n91 VTAIL.n90 10.6058
R172 VTAIL.n75 VTAIL.n74 10.6058
R173 VTAIL.n57 VTAIL.n56 10.6058
R174 VTAIL.n134 VTAIL.n120 9.69747
R175 VTAIL.n16 VTAIL.n2 9.69747
R176 VTAIL.n32 VTAIL.n18 9.69747
R177 VTAIL.n50 VTAIL.n36 9.69747
R178 VTAIL.n118 VTAIL.n104 9.69747
R179 VTAIL.n100 VTAIL.n86 9.69747
R180 VTAIL.n84 VTAIL.n70 9.69747
R181 VTAIL.n66 VTAIL.n52 9.69747
R182 VTAIL.n0 VTAIL.t11 9.589
R183 VTAIL.n0 VTAIL.t14 9.589
R184 VTAIL.n34 VTAIL.t0 9.589
R185 VTAIL.n34 VTAIL.t7 9.589
R186 VTAIL.n102 VTAIL.t6 9.589
R187 VTAIL.n102 VTAIL.t1 9.589
R188 VTAIL.n68 VTAIL.t9 9.589
R189 VTAIL.n68 VTAIL.t8 9.589
R190 VTAIL.n134 VTAIL.n133 9.45567
R191 VTAIL.n16 VTAIL.n15 9.45567
R192 VTAIL.n32 VTAIL.n31 9.45567
R193 VTAIL.n50 VTAIL.n49 9.45567
R194 VTAIL.n118 VTAIL.n117 9.45567
R195 VTAIL.n100 VTAIL.n99 9.45567
R196 VTAIL.n84 VTAIL.n83 9.45567
R197 VTAIL.n66 VTAIL.n65 9.45567
R198 VTAIL.n127 VTAIL.n126 9.3005
R199 VTAIL.n122 VTAIL.n121 9.3005
R200 VTAIL.n133 VTAIL.n132 9.3005
R201 VTAIL.n9 VTAIL.n8 9.3005
R202 VTAIL.n4 VTAIL.n3 9.3005
R203 VTAIL.n15 VTAIL.n14 9.3005
R204 VTAIL.n25 VTAIL.n24 9.3005
R205 VTAIL.n20 VTAIL.n19 9.3005
R206 VTAIL.n31 VTAIL.n30 9.3005
R207 VTAIL.n43 VTAIL.n42 9.3005
R208 VTAIL.n38 VTAIL.n37 9.3005
R209 VTAIL.n49 VTAIL.n48 9.3005
R210 VTAIL.n106 VTAIL.n105 9.3005
R211 VTAIL.n111 VTAIL.n110 9.3005
R212 VTAIL.n117 VTAIL.n116 9.3005
R213 VTAIL.n88 VTAIL.n87 9.3005
R214 VTAIL.n99 VTAIL.n98 9.3005
R215 VTAIL.n93 VTAIL.n92 9.3005
R216 VTAIL.n72 VTAIL.n71 9.3005
R217 VTAIL.n83 VTAIL.n82 9.3005
R218 VTAIL.n77 VTAIL.n76 9.3005
R219 VTAIL.n54 VTAIL.n53 9.3005
R220 VTAIL.n65 VTAIL.n64 9.3005
R221 VTAIL.n59 VTAIL.n58 9.3005
R222 VTAIL.n132 VTAIL.n131 8.92171
R223 VTAIL.n14 VTAIL.n13 8.92171
R224 VTAIL.n30 VTAIL.n29 8.92171
R225 VTAIL.n48 VTAIL.n47 8.92171
R226 VTAIL.n116 VTAIL.n115 8.92171
R227 VTAIL.n98 VTAIL.n97 8.92171
R228 VTAIL.n82 VTAIL.n81 8.92171
R229 VTAIL.n64 VTAIL.n63 8.92171
R230 VTAIL.n128 VTAIL.n122 8.14595
R231 VTAIL.n10 VTAIL.n4 8.14595
R232 VTAIL.n26 VTAIL.n20 8.14595
R233 VTAIL.n44 VTAIL.n38 8.14595
R234 VTAIL.n112 VTAIL.n106 8.14595
R235 VTAIL.n94 VTAIL.n88 8.14595
R236 VTAIL.n78 VTAIL.n72 8.14595
R237 VTAIL.n60 VTAIL.n54 8.14595
R238 VTAIL.n127 VTAIL.n124 7.3702
R239 VTAIL.n9 VTAIL.n6 7.3702
R240 VTAIL.n25 VTAIL.n22 7.3702
R241 VTAIL.n43 VTAIL.n40 7.3702
R242 VTAIL.n111 VTAIL.n108 7.3702
R243 VTAIL.n93 VTAIL.n90 7.3702
R244 VTAIL.n77 VTAIL.n74 7.3702
R245 VTAIL.n59 VTAIL.n56 7.3702
R246 VTAIL.n128 VTAIL.n127 5.81868
R247 VTAIL.n10 VTAIL.n9 5.81868
R248 VTAIL.n26 VTAIL.n25 5.81868
R249 VTAIL.n44 VTAIL.n43 5.81868
R250 VTAIL.n112 VTAIL.n111 5.81868
R251 VTAIL.n94 VTAIL.n93 5.81868
R252 VTAIL.n78 VTAIL.n77 5.81868
R253 VTAIL.n60 VTAIL.n59 5.81868
R254 VTAIL.n131 VTAIL.n122 5.04292
R255 VTAIL.n13 VTAIL.n4 5.04292
R256 VTAIL.n29 VTAIL.n20 5.04292
R257 VTAIL.n47 VTAIL.n38 5.04292
R258 VTAIL.n115 VTAIL.n106 5.04292
R259 VTAIL.n97 VTAIL.n88 5.04292
R260 VTAIL.n81 VTAIL.n72 5.04292
R261 VTAIL.n63 VTAIL.n54 5.04292
R262 VTAIL.n132 VTAIL.n120 4.26717
R263 VTAIL.n14 VTAIL.n2 4.26717
R264 VTAIL.n30 VTAIL.n18 4.26717
R265 VTAIL.n48 VTAIL.n36 4.26717
R266 VTAIL.n116 VTAIL.n104 4.26717
R267 VTAIL.n98 VTAIL.n86 4.26717
R268 VTAIL.n82 VTAIL.n70 4.26717
R269 VTAIL.n64 VTAIL.n52 4.26717
R270 VTAIL.n126 VTAIL.n125 2.5326
R271 VTAIL.n8 VTAIL.n7 2.5326
R272 VTAIL.n24 VTAIL.n23 2.5326
R273 VTAIL.n42 VTAIL.n41 2.5326
R274 VTAIL.n110 VTAIL.n109 2.5326
R275 VTAIL.n92 VTAIL.n91 2.5326
R276 VTAIL.n76 VTAIL.n75 2.5326
R277 VTAIL.n58 VTAIL.n57 2.5326
R278 VTAIL.n69 VTAIL.n67 1.94016
R279 VTAIL.n85 VTAIL.n69 1.94016
R280 VTAIL.n103 VTAIL.n101 1.94016
R281 VTAIL.n119 VTAIL.n103 1.94016
R282 VTAIL.n51 VTAIL.n35 1.94016
R283 VTAIL.n35 VTAIL.n33 1.94016
R284 VTAIL.n17 VTAIL.n1 1.94016
R285 VTAIL VTAIL.n135 1.88197
R286 VTAIL.n101 VTAIL.n85 0.470328
R287 VTAIL.n33 VTAIL.n17 0.470328
R288 VTAIL.n126 VTAIL.n121 0.155672
R289 VTAIL.n133 VTAIL.n121 0.155672
R290 VTAIL.n8 VTAIL.n3 0.155672
R291 VTAIL.n15 VTAIL.n3 0.155672
R292 VTAIL.n24 VTAIL.n19 0.155672
R293 VTAIL.n31 VTAIL.n19 0.155672
R294 VTAIL.n42 VTAIL.n37 0.155672
R295 VTAIL.n49 VTAIL.n37 0.155672
R296 VTAIL.n117 VTAIL.n105 0.155672
R297 VTAIL.n110 VTAIL.n105 0.155672
R298 VTAIL.n99 VTAIL.n87 0.155672
R299 VTAIL.n92 VTAIL.n87 0.155672
R300 VTAIL.n83 VTAIL.n71 0.155672
R301 VTAIL.n76 VTAIL.n71 0.155672
R302 VTAIL.n65 VTAIL.n53 0.155672
R303 VTAIL.n58 VTAIL.n53 0.155672
R304 VTAIL VTAIL.n1 0.0586897
R305 VP.n14 VP.n11 161.3
R306 VP.n16 VP.n15 161.3
R307 VP.n17 VP.n10 161.3
R308 VP.n19 VP.n18 161.3
R309 VP.n20 VP.n9 161.3
R310 VP.n23 VP.n22 161.3
R311 VP.n24 VP.n8 161.3
R312 VP.n26 VP.n25 161.3
R313 VP.n27 VP.n7 161.3
R314 VP.n52 VP.n0 161.3
R315 VP.n51 VP.n50 161.3
R316 VP.n49 VP.n1 161.3
R317 VP.n48 VP.n47 161.3
R318 VP.n45 VP.n2 161.3
R319 VP.n44 VP.n43 161.3
R320 VP.n42 VP.n3 161.3
R321 VP.n41 VP.n40 161.3
R322 VP.n39 VP.n4 161.3
R323 VP.n37 VP.n36 161.3
R324 VP.n35 VP.n5 161.3
R325 VP.n34 VP.n33 161.3
R326 VP.n32 VP.n6 161.3
R327 VP.n31 VP.n30 92.4062
R328 VP.n54 VP.n53 92.4062
R329 VP.n29 VP.n28 92.4062
R330 VP.n12 VP.t3 72.5661
R331 VP.n13 VP.n12 63.4562
R332 VP.n33 VP.n5 56.5193
R333 VP.n51 VP.n1 56.5193
R334 VP.n26 VP.n8 56.5193
R335 VP.n31 VP.t1 42.5521
R336 VP.n38 VP.t6 42.5521
R337 VP.n46 VP.t2 42.5521
R338 VP.n53 VP.t5 42.5521
R339 VP.n28 VP.t0 42.5521
R340 VP.n21 VP.t4 42.5521
R341 VP.n13 VP.t7 42.5521
R342 VP.n30 VP.n29 41.1738
R343 VP.n40 VP.n3 40.4934
R344 VP.n44 VP.n3 40.4934
R345 VP.n19 VP.n10 40.4934
R346 VP.n15 VP.n10 40.4934
R347 VP.n33 VP.n32 24.4675
R348 VP.n37 VP.n5 24.4675
R349 VP.n40 VP.n39 24.4675
R350 VP.n45 VP.n44 24.4675
R351 VP.n47 VP.n1 24.4675
R352 VP.n52 VP.n51 24.4675
R353 VP.n27 VP.n26 24.4675
R354 VP.n20 VP.n19 24.4675
R355 VP.n22 VP.n8 24.4675
R356 VP.n15 VP.n14 24.4675
R357 VP.n32 VP.n31 18.3508
R358 VP.n38 VP.n37 18.3508
R359 VP.n47 VP.n46 18.3508
R360 VP.n53 VP.n52 18.3508
R361 VP.n28 VP.n27 18.3508
R362 VP.n22 VP.n21 18.3508
R363 VP.n12 VP.n11 13.5379
R364 VP.n39 VP.n38 6.11725
R365 VP.n46 VP.n45 6.11725
R366 VP.n21 VP.n20 6.11725
R367 VP.n14 VP.n13 6.11725
R368 VP.n29 VP.n7 0.278367
R369 VP.n30 VP.n6 0.278367
R370 VP.n54 VP.n0 0.278367
R371 VP.n16 VP.n11 0.189894
R372 VP.n17 VP.n16 0.189894
R373 VP.n18 VP.n17 0.189894
R374 VP.n18 VP.n9 0.189894
R375 VP.n23 VP.n9 0.189894
R376 VP.n24 VP.n23 0.189894
R377 VP.n25 VP.n24 0.189894
R378 VP.n25 VP.n7 0.189894
R379 VP.n34 VP.n6 0.189894
R380 VP.n35 VP.n34 0.189894
R381 VP.n36 VP.n35 0.189894
R382 VP.n36 VP.n4 0.189894
R383 VP.n41 VP.n4 0.189894
R384 VP.n42 VP.n41 0.189894
R385 VP.n43 VP.n42 0.189894
R386 VP.n43 VP.n2 0.189894
R387 VP.n48 VP.n2 0.189894
R388 VP.n49 VP.n48 0.189894
R389 VP.n50 VP.n49 0.189894
R390 VP.n50 VP.n0 0.189894
R391 VP VP.n54 0.153454
R392 VDD1 VDD1.n0 128.201
R393 VDD1.n3 VDD1.n2 128.087
R394 VDD1.n3 VDD1.n1 128.087
R395 VDD1.n5 VDD1.n4 127.172
R396 VDD1.n5 VDD1.n3 35.9492
R397 VDD1.n4 VDD1.t3 9.589
R398 VDD1.n4 VDD1.t7 9.589
R399 VDD1.n0 VDD1.t4 9.589
R400 VDD1.n0 VDD1.t0 9.589
R401 VDD1.n2 VDD1.t5 9.589
R402 VDD1.n2 VDD1.t2 9.589
R403 VDD1.n1 VDD1.t6 9.589
R404 VDD1.n1 VDD1.t1 9.589
R405 VDD1 VDD1.n5 0.912138
R406 B.n385 B.n48 585
R407 B.n387 B.n386 585
R408 B.n388 B.n47 585
R409 B.n390 B.n389 585
R410 B.n391 B.n46 585
R411 B.n393 B.n392 585
R412 B.n394 B.n45 585
R413 B.n396 B.n395 585
R414 B.n397 B.n44 585
R415 B.n399 B.n398 585
R416 B.n400 B.n43 585
R417 B.n402 B.n401 585
R418 B.n403 B.n42 585
R419 B.n405 B.n404 585
R420 B.n406 B.n41 585
R421 B.n408 B.n407 585
R422 B.n410 B.n38 585
R423 B.n412 B.n411 585
R424 B.n413 B.n37 585
R425 B.n415 B.n414 585
R426 B.n416 B.n36 585
R427 B.n418 B.n417 585
R428 B.n419 B.n35 585
R429 B.n421 B.n420 585
R430 B.n422 B.n31 585
R431 B.n424 B.n423 585
R432 B.n425 B.n30 585
R433 B.n427 B.n426 585
R434 B.n428 B.n29 585
R435 B.n430 B.n429 585
R436 B.n431 B.n28 585
R437 B.n433 B.n432 585
R438 B.n434 B.n27 585
R439 B.n436 B.n435 585
R440 B.n437 B.n26 585
R441 B.n439 B.n438 585
R442 B.n440 B.n25 585
R443 B.n442 B.n441 585
R444 B.n443 B.n24 585
R445 B.n445 B.n444 585
R446 B.n446 B.n23 585
R447 B.n448 B.n447 585
R448 B.n384 B.n383 585
R449 B.n382 B.n49 585
R450 B.n381 B.n380 585
R451 B.n379 B.n50 585
R452 B.n378 B.n377 585
R453 B.n376 B.n51 585
R454 B.n375 B.n374 585
R455 B.n373 B.n52 585
R456 B.n372 B.n371 585
R457 B.n370 B.n53 585
R458 B.n369 B.n368 585
R459 B.n367 B.n54 585
R460 B.n366 B.n365 585
R461 B.n364 B.n55 585
R462 B.n363 B.n362 585
R463 B.n361 B.n56 585
R464 B.n360 B.n359 585
R465 B.n358 B.n57 585
R466 B.n357 B.n356 585
R467 B.n355 B.n58 585
R468 B.n354 B.n353 585
R469 B.n352 B.n59 585
R470 B.n351 B.n350 585
R471 B.n349 B.n60 585
R472 B.n348 B.n347 585
R473 B.n346 B.n61 585
R474 B.n345 B.n344 585
R475 B.n343 B.n62 585
R476 B.n342 B.n341 585
R477 B.n340 B.n63 585
R478 B.n339 B.n338 585
R479 B.n337 B.n64 585
R480 B.n336 B.n335 585
R481 B.n334 B.n65 585
R482 B.n333 B.n332 585
R483 B.n331 B.n66 585
R484 B.n330 B.n329 585
R485 B.n328 B.n67 585
R486 B.n327 B.n326 585
R487 B.n325 B.n68 585
R488 B.n324 B.n323 585
R489 B.n322 B.n69 585
R490 B.n321 B.n320 585
R491 B.n319 B.n70 585
R492 B.n318 B.n317 585
R493 B.n316 B.n71 585
R494 B.n315 B.n314 585
R495 B.n313 B.n72 585
R496 B.n312 B.n311 585
R497 B.n310 B.n73 585
R498 B.n309 B.n308 585
R499 B.n307 B.n74 585
R500 B.n306 B.n305 585
R501 B.n304 B.n75 585
R502 B.n303 B.n302 585
R503 B.n301 B.n76 585
R504 B.n300 B.n299 585
R505 B.n298 B.n77 585
R506 B.n297 B.n296 585
R507 B.n295 B.n78 585
R508 B.n294 B.n293 585
R509 B.n292 B.n79 585
R510 B.n291 B.n290 585
R511 B.n289 B.n80 585
R512 B.n288 B.n287 585
R513 B.n286 B.n81 585
R514 B.n285 B.n284 585
R515 B.n283 B.n82 585
R516 B.n282 B.n281 585
R517 B.n280 B.n83 585
R518 B.n279 B.n278 585
R519 B.n277 B.n84 585
R520 B.n276 B.n275 585
R521 B.n274 B.n85 585
R522 B.n273 B.n272 585
R523 B.n271 B.n86 585
R524 B.n270 B.n269 585
R525 B.n268 B.n87 585
R526 B.n267 B.n266 585
R527 B.n265 B.n88 585
R528 B.n264 B.n263 585
R529 B.n262 B.n89 585
R530 B.n261 B.n260 585
R531 B.n196 B.n115 585
R532 B.n198 B.n197 585
R533 B.n199 B.n114 585
R534 B.n201 B.n200 585
R535 B.n202 B.n113 585
R536 B.n204 B.n203 585
R537 B.n205 B.n112 585
R538 B.n207 B.n206 585
R539 B.n208 B.n111 585
R540 B.n210 B.n209 585
R541 B.n211 B.n110 585
R542 B.n213 B.n212 585
R543 B.n214 B.n109 585
R544 B.n216 B.n215 585
R545 B.n217 B.n108 585
R546 B.n219 B.n218 585
R547 B.n221 B.n220 585
R548 B.n222 B.n104 585
R549 B.n224 B.n223 585
R550 B.n225 B.n103 585
R551 B.n227 B.n226 585
R552 B.n228 B.n102 585
R553 B.n230 B.n229 585
R554 B.n231 B.n101 585
R555 B.n233 B.n232 585
R556 B.n234 B.n98 585
R557 B.n237 B.n236 585
R558 B.n238 B.n97 585
R559 B.n240 B.n239 585
R560 B.n241 B.n96 585
R561 B.n243 B.n242 585
R562 B.n244 B.n95 585
R563 B.n246 B.n245 585
R564 B.n247 B.n94 585
R565 B.n249 B.n248 585
R566 B.n250 B.n93 585
R567 B.n252 B.n251 585
R568 B.n253 B.n92 585
R569 B.n255 B.n254 585
R570 B.n256 B.n91 585
R571 B.n258 B.n257 585
R572 B.n259 B.n90 585
R573 B.n195 B.n194 585
R574 B.n193 B.n116 585
R575 B.n192 B.n191 585
R576 B.n190 B.n117 585
R577 B.n189 B.n188 585
R578 B.n187 B.n118 585
R579 B.n186 B.n185 585
R580 B.n184 B.n119 585
R581 B.n183 B.n182 585
R582 B.n181 B.n120 585
R583 B.n180 B.n179 585
R584 B.n178 B.n121 585
R585 B.n177 B.n176 585
R586 B.n175 B.n122 585
R587 B.n174 B.n173 585
R588 B.n172 B.n123 585
R589 B.n171 B.n170 585
R590 B.n169 B.n124 585
R591 B.n168 B.n167 585
R592 B.n166 B.n125 585
R593 B.n165 B.n164 585
R594 B.n163 B.n126 585
R595 B.n162 B.n161 585
R596 B.n160 B.n127 585
R597 B.n159 B.n158 585
R598 B.n157 B.n128 585
R599 B.n156 B.n155 585
R600 B.n154 B.n129 585
R601 B.n153 B.n152 585
R602 B.n151 B.n130 585
R603 B.n150 B.n149 585
R604 B.n148 B.n131 585
R605 B.n147 B.n146 585
R606 B.n145 B.n132 585
R607 B.n144 B.n143 585
R608 B.n142 B.n133 585
R609 B.n141 B.n140 585
R610 B.n139 B.n134 585
R611 B.n138 B.n137 585
R612 B.n136 B.n135 585
R613 B.n2 B.n0 585
R614 B.n509 B.n1 585
R615 B.n508 B.n507 585
R616 B.n506 B.n3 585
R617 B.n505 B.n504 585
R618 B.n503 B.n4 585
R619 B.n502 B.n501 585
R620 B.n500 B.n5 585
R621 B.n499 B.n498 585
R622 B.n497 B.n6 585
R623 B.n496 B.n495 585
R624 B.n494 B.n7 585
R625 B.n493 B.n492 585
R626 B.n491 B.n8 585
R627 B.n490 B.n489 585
R628 B.n488 B.n9 585
R629 B.n487 B.n486 585
R630 B.n485 B.n10 585
R631 B.n484 B.n483 585
R632 B.n482 B.n11 585
R633 B.n481 B.n480 585
R634 B.n479 B.n12 585
R635 B.n478 B.n477 585
R636 B.n476 B.n13 585
R637 B.n475 B.n474 585
R638 B.n473 B.n14 585
R639 B.n472 B.n471 585
R640 B.n470 B.n15 585
R641 B.n469 B.n468 585
R642 B.n467 B.n16 585
R643 B.n466 B.n465 585
R644 B.n464 B.n17 585
R645 B.n463 B.n462 585
R646 B.n461 B.n18 585
R647 B.n460 B.n459 585
R648 B.n458 B.n19 585
R649 B.n457 B.n456 585
R650 B.n455 B.n20 585
R651 B.n454 B.n453 585
R652 B.n452 B.n21 585
R653 B.n451 B.n450 585
R654 B.n449 B.n22 585
R655 B.n511 B.n510 585
R656 B.n196 B.n195 545.355
R657 B.n449 B.n448 545.355
R658 B.n261 B.n90 545.355
R659 B.n383 B.n48 545.355
R660 B.n99 B.t2 272.882
R661 B.n39 B.t7 272.882
R662 B.n105 B.t5 272.882
R663 B.n32 B.t10 272.882
R664 B.n99 B.t0 249.275
R665 B.n105 B.t3 249.275
R666 B.n32 B.t9 249.275
R667 B.n39 B.t6 249.275
R668 B.n100 B.t1 229.245
R669 B.n40 B.t8 229.245
R670 B.n106 B.t4 229.245
R671 B.n33 B.t11 229.245
R672 B.n195 B.n116 163.367
R673 B.n191 B.n116 163.367
R674 B.n191 B.n190 163.367
R675 B.n190 B.n189 163.367
R676 B.n189 B.n118 163.367
R677 B.n185 B.n118 163.367
R678 B.n185 B.n184 163.367
R679 B.n184 B.n183 163.367
R680 B.n183 B.n120 163.367
R681 B.n179 B.n120 163.367
R682 B.n179 B.n178 163.367
R683 B.n178 B.n177 163.367
R684 B.n177 B.n122 163.367
R685 B.n173 B.n122 163.367
R686 B.n173 B.n172 163.367
R687 B.n172 B.n171 163.367
R688 B.n171 B.n124 163.367
R689 B.n167 B.n124 163.367
R690 B.n167 B.n166 163.367
R691 B.n166 B.n165 163.367
R692 B.n165 B.n126 163.367
R693 B.n161 B.n126 163.367
R694 B.n161 B.n160 163.367
R695 B.n160 B.n159 163.367
R696 B.n159 B.n128 163.367
R697 B.n155 B.n128 163.367
R698 B.n155 B.n154 163.367
R699 B.n154 B.n153 163.367
R700 B.n153 B.n130 163.367
R701 B.n149 B.n130 163.367
R702 B.n149 B.n148 163.367
R703 B.n148 B.n147 163.367
R704 B.n147 B.n132 163.367
R705 B.n143 B.n132 163.367
R706 B.n143 B.n142 163.367
R707 B.n142 B.n141 163.367
R708 B.n141 B.n134 163.367
R709 B.n137 B.n134 163.367
R710 B.n137 B.n136 163.367
R711 B.n136 B.n2 163.367
R712 B.n510 B.n2 163.367
R713 B.n510 B.n509 163.367
R714 B.n509 B.n508 163.367
R715 B.n508 B.n3 163.367
R716 B.n504 B.n3 163.367
R717 B.n504 B.n503 163.367
R718 B.n503 B.n502 163.367
R719 B.n502 B.n5 163.367
R720 B.n498 B.n5 163.367
R721 B.n498 B.n497 163.367
R722 B.n497 B.n496 163.367
R723 B.n496 B.n7 163.367
R724 B.n492 B.n7 163.367
R725 B.n492 B.n491 163.367
R726 B.n491 B.n490 163.367
R727 B.n490 B.n9 163.367
R728 B.n486 B.n9 163.367
R729 B.n486 B.n485 163.367
R730 B.n485 B.n484 163.367
R731 B.n484 B.n11 163.367
R732 B.n480 B.n11 163.367
R733 B.n480 B.n479 163.367
R734 B.n479 B.n478 163.367
R735 B.n478 B.n13 163.367
R736 B.n474 B.n13 163.367
R737 B.n474 B.n473 163.367
R738 B.n473 B.n472 163.367
R739 B.n472 B.n15 163.367
R740 B.n468 B.n15 163.367
R741 B.n468 B.n467 163.367
R742 B.n467 B.n466 163.367
R743 B.n466 B.n17 163.367
R744 B.n462 B.n17 163.367
R745 B.n462 B.n461 163.367
R746 B.n461 B.n460 163.367
R747 B.n460 B.n19 163.367
R748 B.n456 B.n19 163.367
R749 B.n456 B.n455 163.367
R750 B.n455 B.n454 163.367
R751 B.n454 B.n21 163.367
R752 B.n450 B.n21 163.367
R753 B.n450 B.n449 163.367
R754 B.n197 B.n196 163.367
R755 B.n197 B.n114 163.367
R756 B.n201 B.n114 163.367
R757 B.n202 B.n201 163.367
R758 B.n203 B.n202 163.367
R759 B.n203 B.n112 163.367
R760 B.n207 B.n112 163.367
R761 B.n208 B.n207 163.367
R762 B.n209 B.n208 163.367
R763 B.n209 B.n110 163.367
R764 B.n213 B.n110 163.367
R765 B.n214 B.n213 163.367
R766 B.n215 B.n214 163.367
R767 B.n215 B.n108 163.367
R768 B.n219 B.n108 163.367
R769 B.n220 B.n219 163.367
R770 B.n220 B.n104 163.367
R771 B.n224 B.n104 163.367
R772 B.n225 B.n224 163.367
R773 B.n226 B.n225 163.367
R774 B.n226 B.n102 163.367
R775 B.n230 B.n102 163.367
R776 B.n231 B.n230 163.367
R777 B.n232 B.n231 163.367
R778 B.n232 B.n98 163.367
R779 B.n237 B.n98 163.367
R780 B.n238 B.n237 163.367
R781 B.n239 B.n238 163.367
R782 B.n239 B.n96 163.367
R783 B.n243 B.n96 163.367
R784 B.n244 B.n243 163.367
R785 B.n245 B.n244 163.367
R786 B.n245 B.n94 163.367
R787 B.n249 B.n94 163.367
R788 B.n250 B.n249 163.367
R789 B.n251 B.n250 163.367
R790 B.n251 B.n92 163.367
R791 B.n255 B.n92 163.367
R792 B.n256 B.n255 163.367
R793 B.n257 B.n256 163.367
R794 B.n257 B.n90 163.367
R795 B.n262 B.n261 163.367
R796 B.n263 B.n262 163.367
R797 B.n263 B.n88 163.367
R798 B.n267 B.n88 163.367
R799 B.n268 B.n267 163.367
R800 B.n269 B.n268 163.367
R801 B.n269 B.n86 163.367
R802 B.n273 B.n86 163.367
R803 B.n274 B.n273 163.367
R804 B.n275 B.n274 163.367
R805 B.n275 B.n84 163.367
R806 B.n279 B.n84 163.367
R807 B.n280 B.n279 163.367
R808 B.n281 B.n280 163.367
R809 B.n281 B.n82 163.367
R810 B.n285 B.n82 163.367
R811 B.n286 B.n285 163.367
R812 B.n287 B.n286 163.367
R813 B.n287 B.n80 163.367
R814 B.n291 B.n80 163.367
R815 B.n292 B.n291 163.367
R816 B.n293 B.n292 163.367
R817 B.n293 B.n78 163.367
R818 B.n297 B.n78 163.367
R819 B.n298 B.n297 163.367
R820 B.n299 B.n298 163.367
R821 B.n299 B.n76 163.367
R822 B.n303 B.n76 163.367
R823 B.n304 B.n303 163.367
R824 B.n305 B.n304 163.367
R825 B.n305 B.n74 163.367
R826 B.n309 B.n74 163.367
R827 B.n310 B.n309 163.367
R828 B.n311 B.n310 163.367
R829 B.n311 B.n72 163.367
R830 B.n315 B.n72 163.367
R831 B.n316 B.n315 163.367
R832 B.n317 B.n316 163.367
R833 B.n317 B.n70 163.367
R834 B.n321 B.n70 163.367
R835 B.n322 B.n321 163.367
R836 B.n323 B.n322 163.367
R837 B.n323 B.n68 163.367
R838 B.n327 B.n68 163.367
R839 B.n328 B.n327 163.367
R840 B.n329 B.n328 163.367
R841 B.n329 B.n66 163.367
R842 B.n333 B.n66 163.367
R843 B.n334 B.n333 163.367
R844 B.n335 B.n334 163.367
R845 B.n335 B.n64 163.367
R846 B.n339 B.n64 163.367
R847 B.n340 B.n339 163.367
R848 B.n341 B.n340 163.367
R849 B.n341 B.n62 163.367
R850 B.n345 B.n62 163.367
R851 B.n346 B.n345 163.367
R852 B.n347 B.n346 163.367
R853 B.n347 B.n60 163.367
R854 B.n351 B.n60 163.367
R855 B.n352 B.n351 163.367
R856 B.n353 B.n352 163.367
R857 B.n353 B.n58 163.367
R858 B.n357 B.n58 163.367
R859 B.n358 B.n357 163.367
R860 B.n359 B.n358 163.367
R861 B.n359 B.n56 163.367
R862 B.n363 B.n56 163.367
R863 B.n364 B.n363 163.367
R864 B.n365 B.n364 163.367
R865 B.n365 B.n54 163.367
R866 B.n369 B.n54 163.367
R867 B.n370 B.n369 163.367
R868 B.n371 B.n370 163.367
R869 B.n371 B.n52 163.367
R870 B.n375 B.n52 163.367
R871 B.n376 B.n375 163.367
R872 B.n377 B.n376 163.367
R873 B.n377 B.n50 163.367
R874 B.n381 B.n50 163.367
R875 B.n382 B.n381 163.367
R876 B.n383 B.n382 163.367
R877 B.n448 B.n23 163.367
R878 B.n444 B.n23 163.367
R879 B.n444 B.n443 163.367
R880 B.n443 B.n442 163.367
R881 B.n442 B.n25 163.367
R882 B.n438 B.n25 163.367
R883 B.n438 B.n437 163.367
R884 B.n437 B.n436 163.367
R885 B.n436 B.n27 163.367
R886 B.n432 B.n27 163.367
R887 B.n432 B.n431 163.367
R888 B.n431 B.n430 163.367
R889 B.n430 B.n29 163.367
R890 B.n426 B.n29 163.367
R891 B.n426 B.n425 163.367
R892 B.n425 B.n424 163.367
R893 B.n424 B.n31 163.367
R894 B.n420 B.n31 163.367
R895 B.n420 B.n419 163.367
R896 B.n419 B.n418 163.367
R897 B.n418 B.n36 163.367
R898 B.n414 B.n36 163.367
R899 B.n414 B.n413 163.367
R900 B.n413 B.n412 163.367
R901 B.n412 B.n38 163.367
R902 B.n407 B.n38 163.367
R903 B.n407 B.n406 163.367
R904 B.n406 B.n405 163.367
R905 B.n405 B.n42 163.367
R906 B.n401 B.n42 163.367
R907 B.n401 B.n400 163.367
R908 B.n400 B.n399 163.367
R909 B.n399 B.n44 163.367
R910 B.n395 B.n44 163.367
R911 B.n395 B.n394 163.367
R912 B.n394 B.n393 163.367
R913 B.n393 B.n46 163.367
R914 B.n389 B.n46 163.367
R915 B.n389 B.n388 163.367
R916 B.n388 B.n387 163.367
R917 B.n387 B.n48 163.367
R918 B.n235 B.n100 59.5399
R919 B.n107 B.n106 59.5399
R920 B.n34 B.n33 59.5399
R921 B.n409 B.n40 59.5399
R922 B.n100 B.n99 43.6369
R923 B.n106 B.n105 43.6369
R924 B.n33 B.n32 43.6369
R925 B.n40 B.n39 43.6369
R926 B.n385 B.n384 35.4346
R927 B.n447 B.n22 35.4346
R928 B.n260 B.n259 35.4346
R929 B.n194 B.n115 35.4346
R930 B B.n511 18.0485
R931 B.n447 B.n446 10.6151
R932 B.n446 B.n445 10.6151
R933 B.n445 B.n24 10.6151
R934 B.n441 B.n24 10.6151
R935 B.n441 B.n440 10.6151
R936 B.n440 B.n439 10.6151
R937 B.n439 B.n26 10.6151
R938 B.n435 B.n26 10.6151
R939 B.n435 B.n434 10.6151
R940 B.n434 B.n433 10.6151
R941 B.n433 B.n28 10.6151
R942 B.n429 B.n28 10.6151
R943 B.n429 B.n428 10.6151
R944 B.n428 B.n427 10.6151
R945 B.n427 B.n30 10.6151
R946 B.n423 B.n422 10.6151
R947 B.n422 B.n421 10.6151
R948 B.n421 B.n35 10.6151
R949 B.n417 B.n35 10.6151
R950 B.n417 B.n416 10.6151
R951 B.n416 B.n415 10.6151
R952 B.n415 B.n37 10.6151
R953 B.n411 B.n37 10.6151
R954 B.n411 B.n410 10.6151
R955 B.n408 B.n41 10.6151
R956 B.n404 B.n41 10.6151
R957 B.n404 B.n403 10.6151
R958 B.n403 B.n402 10.6151
R959 B.n402 B.n43 10.6151
R960 B.n398 B.n43 10.6151
R961 B.n398 B.n397 10.6151
R962 B.n397 B.n396 10.6151
R963 B.n396 B.n45 10.6151
R964 B.n392 B.n45 10.6151
R965 B.n392 B.n391 10.6151
R966 B.n391 B.n390 10.6151
R967 B.n390 B.n47 10.6151
R968 B.n386 B.n47 10.6151
R969 B.n386 B.n385 10.6151
R970 B.n260 B.n89 10.6151
R971 B.n264 B.n89 10.6151
R972 B.n265 B.n264 10.6151
R973 B.n266 B.n265 10.6151
R974 B.n266 B.n87 10.6151
R975 B.n270 B.n87 10.6151
R976 B.n271 B.n270 10.6151
R977 B.n272 B.n271 10.6151
R978 B.n272 B.n85 10.6151
R979 B.n276 B.n85 10.6151
R980 B.n277 B.n276 10.6151
R981 B.n278 B.n277 10.6151
R982 B.n278 B.n83 10.6151
R983 B.n282 B.n83 10.6151
R984 B.n283 B.n282 10.6151
R985 B.n284 B.n283 10.6151
R986 B.n284 B.n81 10.6151
R987 B.n288 B.n81 10.6151
R988 B.n289 B.n288 10.6151
R989 B.n290 B.n289 10.6151
R990 B.n290 B.n79 10.6151
R991 B.n294 B.n79 10.6151
R992 B.n295 B.n294 10.6151
R993 B.n296 B.n295 10.6151
R994 B.n296 B.n77 10.6151
R995 B.n300 B.n77 10.6151
R996 B.n301 B.n300 10.6151
R997 B.n302 B.n301 10.6151
R998 B.n302 B.n75 10.6151
R999 B.n306 B.n75 10.6151
R1000 B.n307 B.n306 10.6151
R1001 B.n308 B.n307 10.6151
R1002 B.n308 B.n73 10.6151
R1003 B.n312 B.n73 10.6151
R1004 B.n313 B.n312 10.6151
R1005 B.n314 B.n313 10.6151
R1006 B.n314 B.n71 10.6151
R1007 B.n318 B.n71 10.6151
R1008 B.n319 B.n318 10.6151
R1009 B.n320 B.n319 10.6151
R1010 B.n320 B.n69 10.6151
R1011 B.n324 B.n69 10.6151
R1012 B.n325 B.n324 10.6151
R1013 B.n326 B.n325 10.6151
R1014 B.n326 B.n67 10.6151
R1015 B.n330 B.n67 10.6151
R1016 B.n331 B.n330 10.6151
R1017 B.n332 B.n331 10.6151
R1018 B.n332 B.n65 10.6151
R1019 B.n336 B.n65 10.6151
R1020 B.n337 B.n336 10.6151
R1021 B.n338 B.n337 10.6151
R1022 B.n338 B.n63 10.6151
R1023 B.n342 B.n63 10.6151
R1024 B.n343 B.n342 10.6151
R1025 B.n344 B.n343 10.6151
R1026 B.n344 B.n61 10.6151
R1027 B.n348 B.n61 10.6151
R1028 B.n349 B.n348 10.6151
R1029 B.n350 B.n349 10.6151
R1030 B.n350 B.n59 10.6151
R1031 B.n354 B.n59 10.6151
R1032 B.n355 B.n354 10.6151
R1033 B.n356 B.n355 10.6151
R1034 B.n356 B.n57 10.6151
R1035 B.n360 B.n57 10.6151
R1036 B.n361 B.n360 10.6151
R1037 B.n362 B.n361 10.6151
R1038 B.n362 B.n55 10.6151
R1039 B.n366 B.n55 10.6151
R1040 B.n367 B.n366 10.6151
R1041 B.n368 B.n367 10.6151
R1042 B.n368 B.n53 10.6151
R1043 B.n372 B.n53 10.6151
R1044 B.n373 B.n372 10.6151
R1045 B.n374 B.n373 10.6151
R1046 B.n374 B.n51 10.6151
R1047 B.n378 B.n51 10.6151
R1048 B.n379 B.n378 10.6151
R1049 B.n380 B.n379 10.6151
R1050 B.n380 B.n49 10.6151
R1051 B.n384 B.n49 10.6151
R1052 B.n198 B.n115 10.6151
R1053 B.n199 B.n198 10.6151
R1054 B.n200 B.n199 10.6151
R1055 B.n200 B.n113 10.6151
R1056 B.n204 B.n113 10.6151
R1057 B.n205 B.n204 10.6151
R1058 B.n206 B.n205 10.6151
R1059 B.n206 B.n111 10.6151
R1060 B.n210 B.n111 10.6151
R1061 B.n211 B.n210 10.6151
R1062 B.n212 B.n211 10.6151
R1063 B.n212 B.n109 10.6151
R1064 B.n216 B.n109 10.6151
R1065 B.n217 B.n216 10.6151
R1066 B.n218 B.n217 10.6151
R1067 B.n222 B.n221 10.6151
R1068 B.n223 B.n222 10.6151
R1069 B.n223 B.n103 10.6151
R1070 B.n227 B.n103 10.6151
R1071 B.n228 B.n227 10.6151
R1072 B.n229 B.n228 10.6151
R1073 B.n229 B.n101 10.6151
R1074 B.n233 B.n101 10.6151
R1075 B.n234 B.n233 10.6151
R1076 B.n236 B.n97 10.6151
R1077 B.n240 B.n97 10.6151
R1078 B.n241 B.n240 10.6151
R1079 B.n242 B.n241 10.6151
R1080 B.n242 B.n95 10.6151
R1081 B.n246 B.n95 10.6151
R1082 B.n247 B.n246 10.6151
R1083 B.n248 B.n247 10.6151
R1084 B.n248 B.n93 10.6151
R1085 B.n252 B.n93 10.6151
R1086 B.n253 B.n252 10.6151
R1087 B.n254 B.n253 10.6151
R1088 B.n254 B.n91 10.6151
R1089 B.n258 B.n91 10.6151
R1090 B.n259 B.n258 10.6151
R1091 B.n194 B.n193 10.6151
R1092 B.n193 B.n192 10.6151
R1093 B.n192 B.n117 10.6151
R1094 B.n188 B.n117 10.6151
R1095 B.n188 B.n187 10.6151
R1096 B.n187 B.n186 10.6151
R1097 B.n186 B.n119 10.6151
R1098 B.n182 B.n119 10.6151
R1099 B.n182 B.n181 10.6151
R1100 B.n181 B.n180 10.6151
R1101 B.n180 B.n121 10.6151
R1102 B.n176 B.n121 10.6151
R1103 B.n176 B.n175 10.6151
R1104 B.n175 B.n174 10.6151
R1105 B.n174 B.n123 10.6151
R1106 B.n170 B.n123 10.6151
R1107 B.n170 B.n169 10.6151
R1108 B.n169 B.n168 10.6151
R1109 B.n168 B.n125 10.6151
R1110 B.n164 B.n125 10.6151
R1111 B.n164 B.n163 10.6151
R1112 B.n163 B.n162 10.6151
R1113 B.n162 B.n127 10.6151
R1114 B.n158 B.n127 10.6151
R1115 B.n158 B.n157 10.6151
R1116 B.n157 B.n156 10.6151
R1117 B.n156 B.n129 10.6151
R1118 B.n152 B.n129 10.6151
R1119 B.n152 B.n151 10.6151
R1120 B.n151 B.n150 10.6151
R1121 B.n150 B.n131 10.6151
R1122 B.n146 B.n131 10.6151
R1123 B.n146 B.n145 10.6151
R1124 B.n145 B.n144 10.6151
R1125 B.n144 B.n133 10.6151
R1126 B.n140 B.n133 10.6151
R1127 B.n140 B.n139 10.6151
R1128 B.n139 B.n138 10.6151
R1129 B.n138 B.n135 10.6151
R1130 B.n135 B.n0 10.6151
R1131 B.n507 B.n1 10.6151
R1132 B.n507 B.n506 10.6151
R1133 B.n506 B.n505 10.6151
R1134 B.n505 B.n4 10.6151
R1135 B.n501 B.n4 10.6151
R1136 B.n501 B.n500 10.6151
R1137 B.n500 B.n499 10.6151
R1138 B.n499 B.n6 10.6151
R1139 B.n495 B.n6 10.6151
R1140 B.n495 B.n494 10.6151
R1141 B.n494 B.n493 10.6151
R1142 B.n493 B.n8 10.6151
R1143 B.n489 B.n8 10.6151
R1144 B.n489 B.n488 10.6151
R1145 B.n488 B.n487 10.6151
R1146 B.n487 B.n10 10.6151
R1147 B.n483 B.n10 10.6151
R1148 B.n483 B.n482 10.6151
R1149 B.n482 B.n481 10.6151
R1150 B.n481 B.n12 10.6151
R1151 B.n477 B.n12 10.6151
R1152 B.n477 B.n476 10.6151
R1153 B.n476 B.n475 10.6151
R1154 B.n475 B.n14 10.6151
R1155 B.n471 B.n14 10.6151
R1156 B.n471 B.n470 10.6151
R1157 B.n470 B.n469 10.6151
R1158 B.n469 B.n16 10.6151
R1159 B.n465 B.n16 10.6151
R1160 B.n465 B.n464 10.6151
R1161 B.n464 B.n463 10.6151
R1162 B.n463 B.n18 10.6151
R1163 B.n459 B.n18 10.6151
R1164 B.n459 B.n458 10.6151
R1165 B.n458 B.n457 10.6151
R1166 B.n457 B.n20 10.6151
R1167 B.n453 B.n20 10.6151
R1168 B.n453 B.n452 10.6151
R1169 B.n452 B.n451 10.6151
R1170 B.n451 B.n22 10.6151
R1171 B.n34 B.n30 9.36635
R1172 B.n409 B.n408 9.36635
R1173 B.n218 B.n107 9.36635
R1174 B.n236 B.n235 9.36635
R1175 B.n511 B.n0 2.81026
R1176 B.n511 B.n1 2.81026
R1177 B.n423 B.n34 1.24928
R1178 B.n410 B.n409 1.24928
R1179 B.n221 B.n107 1.24928
R1180 B.n235 B.n234 1.24928
C0 B VDD1 1.21035f
C1 VTAIL VDD1 4.69712f
C2 VDD2 B 1.28514f
C3 VDD2 VTAIL 4.746971f
C4 B VTAIL 1.91124f
C5 VN w_n3220_n1646# 6.21454f
C6 VP w_n3220_n1646# 6.62884f
C7 VDD1 w_n3220_n1646# 1.50144f
C8 VDD2 w_n3220_n1646# 1.58718f
C9 VN VP 5.24658f
C10 B w_n3220_n1646# 6.67619f
C11 VTAIL w_n3220_n1646# 2.15015f
C12 VN VDD1 0.155262f
C13 VP VDD1 2.89707f
C14 VDD2 VN 2.60142f
C15 VDD2 VP 0.452705f
C16 B VN 0.979362f
C17 VN VTAIL 3.32182f
C18 B VP 1.6728f
C19 VTAIL VP 3.33592f
C20 VDD2 VDD1 1.42415f
C21 VDD2 VSUBS 1.2797f
C22 VDD1 VSUBS 1.819708f
C23 VTAIL VSUBS 0.535173f
C24 VN VSUBS 5.61419f
C25 VP VSUBS 2.372417f
C26 B VSUBS 3.313579f
C27 w_n3220_n1646# VSUBS 66.963104f
C28 B.n0 VSUBS 0.004721f
C29 B.n1 VSUBS 0.004721f
C30 B.n2 VSUBS 0.007466f
C31 B.n3 VSUBS 0.007466f
C32 B.n4 VSUBS 0.007466f
C33 B.n5 VSUBS 0.007466f
C34 B.n6 VSUBS 0.007466f
C35 B.n7 VSUBS 0.007466f
C36 B.n8 VSUBS 0.007466f
C37 B.n9 VSUBS 0.007466f
C38 B.n10 VSUBS 0.007466f
C39 B.n11 VSUBS 0.007466f
C40 B.n12 VSUBS 0.007466f
C41 B.n13 VSUBS 0.007466f
C42 B.n14 VSUBS 0.007466f
C43 B.n15 VSUBS 0.007466f
C44 B.n16 VSUBS 0.007466f
C45 B.n17 VSUBS 0.007466f
C46 B.n18 VSUBS 0.007466f
C47 B.n19 VSUBS 0.007466f
C48 B.n20 VSUBS 0.007466f
C49 B.n21 VSUBS 0.007466f
C50 B.n22 VSUBS 0.017979f
C51 B.n23 VSUBS 0.007466f
C52 B.n24 VSUBS 0.007466f
C53 B.n25 VSUBS 0.007466f
C54 B.n26 VSUBS 0.007466f
C55 B.n27 VSUBS 0.007466f
C56 B.n28 VSUBS 0.007466f
C57 B.n29 VSUBS 0.007466f
C58 B.n30 VSUBS 0.007027f
C59 B.n31 VSUBS 0.007466f
C60 B.t11 VSUBS 0.053712f
C61 B.t10 VSUBS 0.068789f
C62 B.t9 VSUBS 0.332513f
C63 B.n32 VSUBS 0.121f
C64 B.n33 VSUBS 0.104933f
C65 B.n34 VSUBS 0.017298f
C66 B.n35 VSUBS 0.007466f
C67 B.n36 VSUBS 0.007466f
C68 B.n37 VSUBS 0.007466f
C69 B.n38 VSUBS 0.007466f
C70 B.t8 VSUBS 0.053713f
C71 B.t7 VSUBS 0.06879f
C72 B.t6 VSUBS 0.332513f
C73 B.n39 VSUBS 0.120999f
C74 B.n40 VSUBS 0.104933f
C75 B.n41 VSUBS 0.007466f
C76 B.n42 VSUBS 0.007466f
C77 B.n43 VSUBS 0.007466f
C78 B.n44 VSUBS 0.007466f
C79 B.n45 VSUBS 0.007466f
C80 B.n46 VSUBS 0.007466f
C81 B.n47 VSUBS 0.007466f
C82 B.n48 VSUBS 0.018911f
C83 B.n49 VSUBS 0.007466f
C84 B.n50 VSUBS 0.007466f
C85 B.n51 VSUBS 0.007466f
C86 B.n52 VSUBS 0.007466f
C87 B.n53 VSUBS 0.007466f
C88 B.n54 VSUBS 0.007466f
C89 B.n55 VSUBS 0.007466f
C90 B.n56 VSUBS 0.007466f
C91 B.n57 VSUBS 0.007466f
C92 B.n58 VSUBS 0.007466f
C93 B.n59 VSUBS 0.007466f
C94 B.n60 VSUBS 0.007466f
C95 B.n61 VSUBS 0.007466f
C96 B.n62 VSUBS 0.007466f
C97 B.n63 VSUBS 0.007466f
C98 B.n64 VSUBS 0.007466f
C99 B.n65 VSUBS 0.007466f
C100 B.n66 VSUBS 0.007466f
C101 B.n67 VSUBS 0.007466f
C102 B.n68 VSUBS 0.007466f
C103 B.n69 VSUBS 0.007466f
C104 B.n70 VSUBS 0.007466f
C105 B.n71 VSUBS 0.007466f
C106 B.n72 VSUBS 0.007466f
C107 B.n73 VSUBS 0.007466f
C108 B.n74 VSUBS 0.007466f
C109 B.n75 VSUBS 0.007466f
C110 B.n76 VSUBS 0.007466f
C111 B.n77 VSUBS 0.007466f
C112 B.n78 VSUBS 0.007466f
C113 B.n79 VSUBS 0.007466f
C114 B.n80 VSUBS 0.007466f
C115 B.n81 VSUBS 0.007466f
C116 B.n82 VSUBS 0.007466f
C117 B.n83 VSUBS 0.007466f
C118 B.n84 VSUBS 0.007466f
C119 B.n85 VSUBS 0.007466f
C120 B.n86 VSUBS 0.007466f
C121 B.n87 VSUBS 0.007466f
C122 B.n88 VSUBS 0.007466f
C123 B.n89 VSUBS 0.007466f
C124 B.n90 VSUBS 0.018911f
C125 B.n91 VSUBS 0.007466f
C126 B.n92 VSUBS 0.007466f
C127 B.n93 VSUBS 0.007466f
C128 B.n94 VSUBS 0.007466f
C129 B.n95 VSUBS 0.007466f
C130 B.n96 VSUBS 0.007466f
C131 B.n97 VSUBS 0.007466f
C132 B.n98 VSUBS 0.007466f
C133 B.t1 VSUBS 0.053713f
C134 B.t2 VSUBS 0.06879f
C135 B.t0 VSUBS 0.332513f
C136 B.n99 VSUBS 0.120999f
C137 B.n100 VSUBS 0.104933f
C138 B.n101 VSUBS 0.007466f
C139 B.n102 VSUBS 0.007466f
C140 B.n103 VSUBS 0.007466f
C141 B.n104 VSUBS 0.007466f
C142 B.t4 VSUBS 0.053712f
C143 B.t5 VSUBS 0.068789f
C144 B.t3 VSUBS 0.332513f
C145 B.n105 VSUBS 0.121f
C146 B.n106 VSUBS 0.104933f
C147 B.n107 VSUBS 0.017298f
C148 B.n108 VSUBS 0.007466f
C149 B.n109 VSUBS 0.007466f
C150 B.n110 VSUBS 0.007466f
C151 B.n111 VSUBS 0.007466f
C152 B.n112 VSUBS 0.007466f
C153 B.n113 VSUBS 0.007466f
C154 B.n114 VSUBS 0.007466f
C155 B.n115 VSUBS 0.018911f
C156 B.n116 VSUBS 0.007466f
C157 B.n117 VSUBS 0.007466f
C158 B.n118 VSUBS 0.007466f
C159 B.n119 VSUBS 0.007466f
C160 B.n120 VSUBS 0.007466f
C161 B.n121 VSUBS 0.007466f
C162 B.n122 VSUBS 0.007466f
C163 B.n123 VSUBS 0.007466f
C164 B.n124 VSUBS 0.007466f
C165 B.n125 VSUBS 0.007466f
C166 B.n126 VSUBS 0.007466f
C167 B.n127 VSUBS 0.007466f
C168 B.n128 VSUBS 0.007466f
C169 B.n129 VSUBS 0.007466f
C170 B.n130 VSUBS 0.007466f
C171 B.n131 VSUBS 0.007466f
C172 B.n132 VSUBS 0.007466f
C173 B.n133 VSUBS 0.007466f
C174 B.n134 VSUBS 0.007466f
C175 B.n135 VSUBS 0.007466f
C176 B.n136 VSUBS 0.007466f
C177 B.n137 VSUBS 0.007466f
C178 B.n138 VSUBS 0.007466f
C179 B.n139 VSUBS 0.007466f
C180 B.n140 VSUBS 0.007466f
C181 B.n141 VSUBS 0.007466f
C182 B.n142 VSUBS 0.007466f
C183 B.n143 VSUBS 0.007466f
C184 B.n144 VSUBS 0.007466f
C185 B.n145 VSUBS 0.007466f
C186 B.n146 VSUBS 0.007466f
C187 B.n147 VSUBS 0.007466f
C188 B.n148 VSUBS 0.007466f
C189 B.n149 VSUBS 0.007466f
C190 B.n150 VSUBS 0.007466f
C191 B.n151 VSUBS 0.007466f
C192 B.n152 VSUBS 0.007466f
C193 B.n153 VSUBS 0.007466f
C194 B.n154 VSUBS 0.007466f
C195 B.n155 VSUBS 0.007466f
C196 B.n156 VSUBS 0.007466f
C197 B.n157 VSUBS 0.007466f
C198 B.n158 VSUBS 0.007466f
C199 B.n159 VSUBS 0.007466f
C200 B.n160 VSUBS 0.007466f
C201 B.n161 VSUBS 0.007466f
C202 B.n162 VSUBS 0.007466f
C203 B.n163 VSUBS 0.007466f
C204 B.n164 VSUBS 0.007466f
C205 B.n165 VSUBS 0.007466f
C206 B.n166 VSUBS 0.007466f
C207 B.n167 VSUBS 0.007466f
C208 B.n168 VSUBS 0.007466f
C209 B.n169 VSUBS 0.007466f
C210 B.n170 VSUBS 0.007466f
C211 B.n171 VSUBS 0.007466f
C212 B.n172 VSUBS 0.007466f
C213 B.n173 VSUBS 0.007466f
C214 B.n174 VSUBS 0.007466f
C215 B.n175 VSUBS 0.007466f
C216 B.n176 VSUBS 0.007466f
C217 B.n177 VSUBS 0.007466f
C218 B.n178 VSUBS 0.007466f
C219 B.n179 VSUBS 0.007466f
C220 B.n180 VSUBS 0.007466f
C221 B.n181 VSUBS 0.007466f
C222 B.n182 VSUBS 0.007466f
C223 B.n183 VSUBS 0.007466f
C224 B.n184 VSUBS 0.007466f
C225 B.n185 VSUBS 0.007466f
C226 B.n186 VSUBS 0.007466f
C227 B.n187 VSUBS 0.007466f
C228 B.n188 VSUBS 0.007466f
C229 B.n189 VSUBS 0.007466f
C230 B.n190 VSUBS 0.007466f
C231 B.n191 VSUBS 0.007466f
C232 B.n192 VSUBS 0.007466f
C233 B.n193 VSUBS 0.007466f
C234 B.n194 VSUBS 0.017979f
C235 B.n195 VSUBS 0.017979f
C236 B.n196 VSUBS 0.018911f
C237 B.n197 VSUBS 0.007466f
C238 B.n198 VSUBS 0.007466f
C239 B.n199 VSUBS 0.007466f
C240 B.n200 VSUBS 0.007466f
C241 B.n201 VSUBS 0.007466f
C242 B.n202 VSUBS 0.007466f
C243 B.n203 VSUBS 0.007466f
C244 B.n204 VSUBS 0.007466f
C245 B.n205 VSUBS 0.007466f
C246 B.n206 VSUBS 0.007466f
C247 B.n207 VSUBS 0.007466f
C248 B.n208 VSUBS 0.007466f
C249 B.n209 VSUBS 0.007466f
C250 B.n210 VSUBS 0.007466f
C251 B.n211 VSUBS 0.007466f
C252 B.n212 VSUBS 0.007466f
C253 B.n213 VSUBS 0.007466f
C254 B.n214 VSUBS 0.007466f
C255 B.n215 VSUBS 0.007466f
C256 B.n216 VSUBS 0.007466f
C257 B.n217 VSUBS 0.007466f
C258 B.n218 VSUBS 0.007027f
C259 B.n219 VSUBS 0.007466f
C260 B.n220 VSUBS 0.007466f
C261 B.n221 VSUBS 0.004172f
C262 B.n222 VSUBS 0.007466f
C263 B.n223 VSUBS 0.007466f
C264 B.n224 VSUBS 0.007466f
C265 B.n225 VSUBS 0.007466f
C266 B.n226 VSUBS 0.007466f
C267 B.n227 VSUBS 0.007466f
C268 B.n228 VSUBS 0.007466f
C269 B.n229 VSUBS 0.007466f
C270 B.n230 VSUBS 0.007466f
C271 B.n231 VSUBS 0.007466f
C272 B.n232 VSUBS 0.007466f
C273 B.n233 VSUBS 0.007466f
C274 B.n234 VSUBS 0.004172f
C275 B.n235 VSUBS 0.017298f
C276 B.n236 VSUBS 0.007027f
C277 B.n237 VSUBS 0.007466f
C278 B.n238 VSUBS 0.007466f
C279 B.n239 VSUBS 0.007466f
C280 B.n240 VSUBS 0.007466f
C281 B.n241 VSUBS 0.007466f
C282 B.n242 VSUBS 0.007466f
C283 B.n243 VSUBS 0.007466f
C284 B.n244 VSUBS 0.007466f
C285 B.n245 VSUBS 0.007466f
C286 B.n246 VSUBS 0.007466f
C287 B.n247 VSUBS 0.007466f
C288 B.n248 VSUBS 0.007466f
C289 B.n249 VSUBS 0.007466f
C290 B.n250 VSUBS 0.007466f
C291 B.n251 VSUBS 0.007466f
C292 B.n252 VSUBS 0.007466f
C293 B.n253 VSUBS 0.007466f
C294 B.n254 VSUBS 0.007466f
C295 B.n255 VSUBS 0.007466f
C296 B.n256 VSUBS 0.007466f
C297 B.n257 VSUBS 0.007466f
C298 B.n258 VSUBS 0.007466f
C299 B.n259 VSUBS 0.018911f
C300 B.n260 VSUBS 0.017979f
C301 B.n261 VSUBS 0.017979f
C302 B.n262 VSUBS 0.007466f
C303 B.n263 VSUBS 0.007466f
C304 B.n264 VSUBS 0.007466f
C305 B.n265 VSUBS 0.007466f
C306 B.n266 VSUBS 0.007466f
C307 B.n267 VSUBS 0.007466f
C308 B.n268 VSUBS 0.007466f
C309 B.n269 VSUBS 0.007466f
C310 B.n270 VSUBS 0.007466f
C311 B.n271 VSUBS 0.007466f
C312 B.n272 VSUBS 0.007466f
C313 B.n273 VSUBS 0.007466f
C314 B.n274 VSUBS 0.007466f
C315 B.n275 VSUBS 0.007466f
C316 B.n276 VSUBS 0.007466f
C317 B.n277 VSUBS 0.007466f
C318 B.n278 VSUBS 0.007466f
C319 B.n279 VSUBS 0.007466f
C320 B.n280 VSUBS 0.007466f
C321 B.n281 VSUBS 0.007466f
C322 B.n282 VSUBS 0.007466f
C323 B.n283 VSUBS 0.007466f
C324 B.n284 VSUBS 0.007466f
C325 B.n285 VSUBS 0.007466f
C326 B.n286 VSUBS 0.007466f
C327 B.n287 VSUBS 0.007466f
C328 B.n288 VSUBS 0.007466f
C329 B.n289 VSUBS 0.007466f
C330 B.n290 VSUBS 0.007466f
C331 B.n291 VSUBS 0.007466f
C332 B.n292 VSUBS 0.007466f
C333 B.n293 VSUBS 0.007466f
C334 B.n294 VSUBS 0.007466f
C335 B.n295 VSUBS 0.007466f
C336 B.n296 VSUBS 0.007466f
C337 B.n297 VSUBS 0.007466f
C338 B.n298 VSUBS 0.007466f
C339 B.n299 VSUBS 0.007466f
C340 B.n300 VSUBS 0.007466f
C341 B.n301 VSUBS 0.007466f
C342 B.n302 VSUBS 0.007466f
C343 B.n303 VSUBS 0.007466f
C344 B.n304 VSUBS 0.007466f
C345 B.n305 VSUBS 0.007466f
C346 B.n306 VSUBS 0.007466f
C347 B.n307 VSUBS 0.007466f
C348 B.n308 VSUBS 0.007466f
C349 B.n309 VSUBS 0.007466f
C350 B.n310 VSUBS 0.007466f
C351 B.n311 VSUBS 0.007466f
C352 B.n312 VSUBS 0.007466f
C353 B.n313 VSUBS 0.007466f
C354 B.n314 VSUBS 0.007466f
C355 B.n315 VSUBS 0.007466f
C356 B.n316 VSUBS 0.007466f
C357 B.n317 VSUBS 0.007466f
C358 B.n318 VSUBS 0.007466f
C359 B.n319 VSUBS 0.007466f
C360 B.n320 VSUBS 0.007466f
C361 B.n321 VSUBS 0.007466f
C362 B.n322 VSUBS 0.007466f
C363 B.n323 VSUBS 0.007466f
C364 B.n324 VSUBS 0.007466f
C365 B.n325 VSUBS 0.007466f
C366 B.n326 VSUBS 0.007466f
C367 B.n327 VSUBS 0.007466f
C368 B.n328 VSUBS 0.007466f
C369 B.n329 VSUBS 0.007466f
C370 B.n330 VSUBS 0.007466f
C371 B.n331 VSUBS 0.007466f
C372 B.n332 VSUBS 0.007466f
C373 B.n333 VSUBS 0.007466f
C374 B.n334 VSUBS 0.007466f
C375 B.n335 VSUBS 0.007466f
C376 B.n336 VSUBS 0.007466f
C377 B.n337 VSUBS 0.007466f
C378 B.n338 VSUBS 0.007466f
C379 B.n339 VSUBS 0.007466f
C380 B.n340 VSUBS 0.007466f
C381 B.n341 VSUBS 0.007466f
C382 B.n342 VSUBS 0.007466f
C383 B.n343 VSUBS 0.007466f
C384 B.n344 VSUBS 0.007466f
C385 B.n345 VSUBS 0.007466f
C386 B.n346 VSUBS 0.007466f
C387 B.n347 VSUBS 0.007466f
C388 B.n348 VSUBS 0.007466f
C389 B.n349 VSUBS 0.007466f
C390 B.n350 VSUBS 0.007466f
C391 B.n351 VSUBS 0.007466f
C392 B.n352 VSUBS 0.007466f
C393 B.n353 VSUBS 0.007466f
C394 B.n354 VSUBS 0.007466f
C395 B.n355 VSUBS 0.007466f
C396 B.n356 VSUBS 0.007466f
C397 B.n357 VSUBS 0.007466f
C398 B.n358 VSUBS 0.007466f
C399 B.n359 VSUBS 0.007466f
C400 B.n360 VSUBS 0.007466f
C401 B.n361 VSUBS 0.007466f
C402 B.n362 VSUBS 0.007466f
C403 B.n363 VSUBS 0.007466f
C404 B.n364 VSUBS 0.007466f
C405 B.n365 VSUBS 0.007466f
C406 B.n366 VSUBS 0.007466f
C407 B.n367 VSUBS 0.007466f
C408 B.n368 VSUBS 0.007466f
C409 B.n369 VSUBS 0.007466f
C410 B.n370 VSUBS 0.007466f
C411 B.n371 VSUBS 0.007466f
C412 B.n372 VSUBS 0.007466f
C413 B.n373 VSUBS 0.007466f
C414 B.n374 VSUBS 0.007466f
C415 B.n375 VSUBS 0.007466f
C416 B.n376 VSUBS 0.007466f
C417 B.n377 VSUBS 0.007466f
C418 B.n378 VSUBS 0.007466f
C419 B.n379 VSUBS 0.007466f
C420 B.n380 VSUBS 0.007466f
C421 B.n381 VSUBS 0.007466f
C422 B.n382 VSUBS 0.007466f
C423 B.n383 VSUBS 0.017979f
C424 B.n384 VSUBS 0.018792f
C425 B.n385 VSUBS 0.018098f
C426 B.n386 VSUBS 0.007466f
C427 B.n387 VSUBS 0.007466f
C428 B.n388 VSUBS 0.007466f
C429 B.n389 VSUBS 0.007466f
C430 B.n390 VSUBS 0.007466f
C431 B.n391 VSUBS 0.007466f
C432 B.n392 VSUBS 0.007466f
C433 B.n393 VSUBS 0.007466f
C434 B.n394 VSUBS 0.007466f
C435 B.n395 VSUBS 0.007466f
C436 B.n396 VSUBS 0.007466f
C437 B.n397 VSUBS 0.007466f
C438 B.n398 VSUBS 0.007466f
C439 B.n399 VSUBS 0.007466f
C440 B.n400 VSUBS 0.007466f
C441 B.n401 VSUBS 0.007466f
C442 B.n402 VSUBS 0.007466f
C443 B.n403 VSUBS 0.007466f
C444 B.n404 VSUBS 0.007466f
C445 B.n405 VSUBS 0.007466f
C446 B.n406 VSUBS 0.007466f
C447 B.n407 VSUBS 0.007466f
C448 B.n408 VSUBS 0.007027f
C449 B.n409 VSUBS 0.017298f
C450 B.n410 VSUBS 0.004172f
C451 B.n411 VSUBS 0.007466f
C452 B.n412 VSUBS 0.007466f
C453 B.n413 VSUBS 0.007466f
C454 B.n414 VSUBS 0.007466f
C455 B.n415 VSUBS 0.007466f
C456 B.n416 VSUBS 0.007466f
C457 B.n417 VSUBS 0.007466f
C458 B.n418 VSUBS 0.007466f
C459 B.n419 VSUBS 0.007466f
C460 B.n420 VSUBS 0.007466f
C461 B.n421 VSUBS 0.007466f
C462 B.n422 VSUBS 0.007466f
C463 B.n423 VSUBS 0.004172f
C464 B.n424 VSUBS 0.007466f
C465 B.n425 VSUBS 0.007466f
C466 B.n426 VSUBS 0.007466f
C467 B.n427 VSUBS 0.007466f
C468 B.n428 VSUBS 0.007466f
C469 B.n429 VSUBS 0.007466f
C470 B.n430 VSUBS 0.007466f
C471 B.n431 VSUBS 0.007466f
C472 B.n432 VSUBS 0.007466f
C473 B.n433 VSUBS 0.007466f
C474 B.n434 VSUBS 0.007466f
C475 B.n435 VSUBS 0.007466f
C476 B.n436 VSUBS 0.007466f
C477 B.n437 VSUBS 0.007466f
C478 B.n438 VSUBS 0.007466f
C479 B.n439 VSUBS 0.007466f
C480 B.n440 VSUBS 0.007466f
C481 B.n441 VSUBS 0.007466f
C482 B.n442 VSUBS 0.007466f
C483 B.n443 VSUBS 0.007466f
C484 B.n444 VSUBS 0.007466f
C485 B.n445 VSUBS 0.007466f
C486 B.n446 VSUBS 0.007466f
C487 B.n447 VSUBS 0.018911f
C488 B.n448 VSUBS 0.018911f
C489 B.n449 VSUBS 0.017979f
C490 B.n450 VSUBS 0.007466f
C491 B.n451 VSUBS 0.007466f
C492 B.n452 VSUBS 0.007466f
C493 B.n453 VSUBS 0.007466f
C494 B.n454 VSUBS 0.007466f
C495 B.n455 VSUBS 0.007466f
C496 B.n456 VSUBS 0.007466f
C497 B.n457 VSUBS 0.007466f
C498 B.n458 VSUBS 0.007466f
C499 B.n459 VSUBS 0.007466f
C500 B.n460 VSUBS 0.007466f
C501 B.n461 VSUBS 0.007466f
C502 B.n462 VSUBS 0.007466f
C503 B.n463 VSUBS 0.007466f
C504 B.n464 VSUBS 0.007466f
C505 B.n465 VSUBS 0.007466f
C506 B.n466 VSUBS 0.007466f
C507 B.n467 VSUBS 0.007466f
C508 B.n468 VSUBS 0.007466f
C509 B.n469 VSUBS 0.007466f
C510 B.n470 VSUBS 0.007466f
C511 B.n471 VSUBS 0.007466f
C512 B.n472 VSUBS 0.007466f
C513 B.n473 VSUBS 0.007466f
C514 B.n474 VSUBS 0.007466f
C515 B.n475 VSUBS 0.007466f
C516 B.n476 VSUBS 0.007466f
C517 B.n477 VSUBS 0.007466f
C518 B.n478 VSUBS 0.007466f
C519 B.n479 VSUBS 0.007466f
C520 B.n480 VSUBS 0.007466f
C521 B.n481 VSUBS 0.007466f
C522 B.n482 VSUBS 0.007466f
C523 B.n483 VSUBS 0.007466f
C524 B.n484 VSUBS 0.007466f
C525 B.n485 VSUBS 0.007466f
C526 B.n486 VSUBS 0.007466f
C527 B.n487 VSUBS 0.007466f
C528 B.n488 VSUBS 0.007466f
C529 B.n489 VSUBS 0.007466f
C530 B.n490 VSUBS 0.007466f
C531 B.n491 VSUBS 0.007466f
C532 B.n492 VSUBS 0.007466f
C533 B.n493 VSUBS 0.007466f
C534 B.n494 VSUBS 0.007466f
C535 B.n495 VSUBS 0.007466f
C536 B.n496 VSUBS 0.007466f
C537 B.n497 VSUBS 0.007466f
C538 B.n498 VSUBS 0.007466f
C539 B.n499 VSUBS 0.007466f
C540 B.n500 VSUBS 0.007466f
C541 B.n501 VSUBS 0.007466f
C542 B.n502 VSUBS 0.007466f
C543 B.n503 VSUBS 0.007466f
C544 B.n504 VSUBS 0.007466f
C545 B.n505 VSUBS 0.007466f
C546 B.n506 VSUBS 0.007466f
C547 B.n507 VSUBS 0.007466f
C548 B.n508 VSUBS 0.007466f
C549 B.n509 VSUBS 0.007466f
C550 B.n510 VSUBS 0.007466f
C551 B.n511 VSUBS 0.016905f
C552 VDD1.t4 VSUBS 0.066758f
C553 VDD1.t0 VSUBS 0.066758f
C554 VDD1.n0 VSUBS 0.358139f
C555 VDD1.t6 VSUBS 0.066758f
C556 VDD1.t1 VSUBS 0.066758f
C557 VDD1.n1 VSUBS 0.357555f
C558 VDD1.t5 VSUBS 0.066758f
C559 VDD1.t2 VSUBS 0.066758f
C560 VDD1.n2 VSUBS 0.357555f
C561 VDD1.n3 VSUBS 2.69158f
C562 VDD1.t3 VSUBS 0.066758f
C563 VDD1.t7 VSUBS 0.066758f
C564 VDD1.n4 VSUBS 0.353379f
C565 VDD1.n5 VSUBS 2.20316f
C566 VP.n0 VSUBS 0.067369f
C567 VP.t5 VSUBS 0.840435f
C568 VP.n1 VSUBS 0.074596f
C569 VP.n2 VSUBS 0.051099f
C570 VP.t2 VSUBS 0.840435f
C571 VP.n3 VSUBS 0.041309f
C572 VP.n4 VSUBS 0.051099f
C573 VP.t6 VSUBS 0.840435f
C574 VP.n5 VSUBS 0.074596f
C575 VP.n6 VSUBS 0.067369f
C576 VP.t1 VSUBS 0.840435f
C577 VP.n7 VSUBS 0.067369f
C578 VP.t0 VSUBS 0.840435f
C579 VP.n8 VSUBS 0.074596f
C580 VP.n9 VSUBS 0.051099f
C581 VP.t4 VSUBS 0.840435f
C582 VP.n10 VSUBS 0.041309f
C583 VP.n11 VSUBS 0.378621f
C584 VP.t7 VSUBS 0.840435f
C585 VP.t3 VSUBS 1.08732f
C586 VP.n12 VSUBS 0.475237f
C587 VP.n13 VSUBS 0.465068f
C588 VP.n14 VSUBS 0.05997f
C589 VP.n15 VSUBS 0.101559f
C590 VP.n16 VSUBS 0.051099f
C591 VP.n17 VSUBS 0.051099f
C592 VP.n18 VSUBS 0.051099f
C593 VP.n19 VSUBS 0.101559f
C594 VP.n20 VSUBS 0.05997f
C595 VP.n21 VSUBS 0.357709f
C596 VP.n22 VSUBS 0.083479f
C597 VP.n23 VSUBS 0.051099f
C598 VP.n24 VSUBS 0.051099f
C599 VP.n25 VSUBS 0.051099f
C600 VP.n26 VSUBS 0.074596f
C601 VP.n27 VSUBS 0.083479f
C602 VP.n28 VSUBS 0.50389f
C603 VP.n29 VSUBS 2.08297f
C604 VP.n30 VSUBS 2.12758f
C605 VP.n31 VSUBS 0.50389f
C606 VP.n32 VSUBS 0.083479f
C607 VP.n33 VSUBS 0.074596f
C608 VP.n34 VSUBS 0.051099f
C609 VP.n35 VSUBS 0.051099f
C610 VP.n36 VSUBS 0.051099f
C611 VP.n37 VSUBS 0.083479f
C612 VP.n38 VSUBS 0.357709f
C613 VP.n39 VSUBS 0.05997f
C614 VP.n40 VSUBS 0.101559f
C615 VP.n41 VSUBS 0.051099f
C616 VP.n42 VSUBS 0.051099f
C617 VP.n43 VSUBS 0.051099f
C618 VP.n44 VSUBS 0.101559f
C619 VP.n45 VSUBS 0.05997f
C620 VP.n46 VSUBS 0.357709f
C621 VP.n47 VSUBS 0.083479f
C622 VP.n48 VSUBS 0.051099f
C623 VP.n49 VSUBS 0.051099f
C624 VP.n50 VSUBS 0.051099f
C625 VP.n51 VSUBS 0.074596f
C626 VP.n52 VSUBS 0.083479f
C627 VP.n53 VSUBS 0.50389f
C628 VP.n54 VSUBS 0.063328f
C629 VTAIL.t11 VSUBS 0.078254f
C630 VTAIL.t14 VSUBS 0.078254f
C631 VTAIL.n0 VSUBS 0.353984f
C632 VTAIL.n1 VSUBS 0.613293f
C633 VTAIL.n2 VSUBS 0.033337f
C634 VTAIL.n3 VSUBS 0.029212f
C635 VTAIL.n4 VSUBS 0.015697f
C636 VTAIL.n5 VSUBS 0.027827f
C637 VTAIL.n6 VSUBS 0.02727f
C638 VTAIL.t15 VSUBS 0.085653f
C639 VTAIL.n7 VSUBS 0.118183f
C640 VTAIL.n8 VSUBS 0.325467f
C641 VTAIL.n9 VSUBS 0.015697f
C642 VTAIL.n10 VSUBS 0.01662f
C643 VTAIL.n11 VSUBS 0.037102f
C644 VTAIL.n12 VSUBS 0.094044f
C645 VTAIL.n13 VSUBS 0.01662f
C646 VTAIL.n14 VSUBS 0.015697f
C647 VTAIL.n15 VSUBS 0.06393f
C648 VTAIL.n16 VSUBS 0.047368f
C649 VTAIL.n17 VSUBS 0.24972f
C650 VTAIL.n18 VSUBS 0.033337f
C651 VTAIL.n19 VSUBS 0.029212f
C652 VTAIL.n20 VSUBS 0.015697f
C653 VTAIL.n21 VSUBS 0.027827f
C654 VTAIL.n22 VSUBS 0.02727f
C655 VTAIL.t2 VSUBS 0.085653f
C656 VTAIL.n23 VSUBS 0.118183f
C657 VTAIL.n24 VSUBS 0.325467f
C658 VTAIL.n25 VSUBS 0.015697f
C659 VTAIL.n26 VSUBS 0.01662f
C660 VTAIL.n27 VSUBS 0.037102f
C661 VTAIL.n28 VSUBS 0.094044f
C662 VTAIL.n29 VSUBS 0.01662f
C663 VTAIL.n30 VSUBS 0.015697f
C664 VTAIL.n31 VSUBS 0.06393f
C665 VTAIL.n32 VSUBS 0.047368f
C666 VTAIL.n33 VSUBS 0.24972f
C667 VTAIL.t0 VSUBS 0.078254f
C668 VTAIL.t7 VSUBS 0.078254f
C669 VTAIL.n34 VSUBS 0.353984f
C670 VTAIL.n35 VSUBS 0.790389f
C671 VTAIL.n36 VSUBS 0.033337f
C672 VTAIL.n37 VSUBS 0.029212f
C673 VTAIL.n38 VSUBS 0.015697f
C674 VTAIL.n39 VSUBS 0.027827f
C675 VTAIL.n40 VSUBS 0.02727f
C676 VTAIL.t3 VSUBS 0.085653f
C677 VTAIL.n41 VSUBS 0.118183f
C678 VTAIL.n42 VSUBS 0.325467f
C679 VTAIL.n43 VSUBS 0.015697f
C680 VTAIL.n44 VSUBS 0.01662f
C681 VTAIL.n45 VSUBS 0.037102f
C682 VTAIL.n46 VSUBS 0.094044f
C683 VTAIL.n47 VSUBS 0.01662f
C684 VTAIL.n48 VSUBS 0.015697f
C685 VTAIL.n49 VSUBS 0.06393f
C686 VTAIL.n50 VSUBS 0.047368f
C687 VTAIL.n51 VSUBS 1.05995f
C688 VTAIL.n52 VSUBS 0.033337f
C689 VTAIL.n53 VSUBS 0.029212f
C690 VTAIL.n54 VSUBS 0.015697f
C691 VTAIL.n55 VSUBS 0.027827f
C692 VTAIL.n56 VSUBS 0.02727f
C693 VTAIL.t13 VSUBS 0.085653f
C694 VTAIL.n57 VSUBS 0.118183f
C695 VTAIL.n58 VSUBS 0.325467f
C696 VTAIL.n59 VSUBS 0.015697f
C697 VTAIL.n60 VSUBS 0.01662f
C698 VTAIL.n61 VSUBS 0.037102f
C699 VTAIL.n62 VSUBS 0.094044f
C700 VTAIL.n63 VSUBS 0.01662f
C701 VTAIL.n64 VSUBS 0.015697f
C702 VTAIL.n65 VSUBS 0.06393f
C703 VTAIL.n66 VSUBS 0.047368f
C704 VTAIL.n67 VSUBS 1.05995f
C705 VTAIL.t9 VSUBS 0.078254f
C706 VTAIL.t8 VSUBS 0.078254f
C707 VTAIL.n68 VSUBS 0.353986f
C708 VTAIL.n69 VSUBS 0.790387f
C709 VTAIL.n70 VSUBS 0.033337f
C710 VTAIL.n71 VSUBS 0.029212f
C711 VTAIL.n72 VSUBS 0.015697f
C712 VTAIL.n73 VSUBS 0.027827f
C713 VTAIL.n74 VSUBS 0.02727f
C714 VTAIL.t12 VSUBS 0.085653f
C715 VTAIL.n75 VSUBS 0.118183f
C716 VTAIL.n76 VSUBS 0.325467f
C717 VTAIL.n77 VSUBS 0.015697f
C718 VTAIL.n78 VSUBS 0.01662f
C719 VTAIL.n79 VSUBS 0.037102f
C720 VTAIL.n80 VSUBS 0.094044f
C721 VTAIL.n81 VSUBS 0.01662f
C722 VTAIL.n82 VSUBS 0.015697f
C723 VTAIL.n83 VSUBS 0.06393f
C724 VTAIL.n84 VSUBS 0.047368f
C725 VTAIL.n85 VSUBS 0.24972f
C726 VTAIL.n86 VSUBS 0.033337f
C727 VTAIL.n87 VSUBS 0.029212f
C728 VTAIL.n88 VSUBS 0.015697f
C729 VTAIL.n89 VSUBS 0.027827f
C730 VTAIL.n90 VSUBS 0.02727f
C731 VTAIL.t5 VSUBS 0.085653f
C732 VTAIL.n91 VSUBS 0.118183f
C733 VTAIL.n92 VSUBS 0.325467f
C734 VTAIL.n93 VSUBS 0.015697f
C735 VTAIL.n94 VSUBS 0.01662f
C736 VTAIL.n95 VSUBS 0.037102f
C737 VTAIL.n96 VSUBS 0.094044f
C738 VTAIL.n97 VSUBS 0.01662f
C739 VTAIL.n98 VSUBS 0.015697f
C740 VTAIL.n99 VSUBS 0.06393f
C741 VTAIL.n100 VSUBS 0.047368f
C742 VTAIL.n101 VSUBS 0.24972f
C743 VTAIL.t6 VSUBS 0.078254f
C744 VTAIL.t1 VSUBS 0.078254f
C745 VTAIL.n102 VSUBS 0.353986f
C746 VTAIL.n103 VSUBS 0.790387f
C747 VTAIL.n104 VSUBS 0.033337f
C748 VTAIL.n105 VSUBS 0.029212f
C749 VTAIL.n106 VSUBS 0.015697f
C750 VTAIL.n107 VSUBS 0.027827f
C751 VTAIL.n108 VSUBS 0.02727f
C752 VTAIL.t4 VSUBS 0.085653f
C753 VTAIL.n109 VSUBS 0.118183f
C754 VTAIL.n110 VSUBS 0.325467f
C755 VTAIL.n111 VSUBS 0.015697f
C756 VTAIL.n112 VSUBS 0.01662f
C757 VTAIL.n113 VSUBS 0.037102f
C758 VTAIL.n114 VSUBS 0.094044f
C759 VTAIL.n115 VSUBS 0.01662f
C760 VTAIL.n116 VSUBS 0.015697f
C761 VTAIL.n117 VSUBS 0.06393f
C762 VTAIL.n118 VSUBS 0.047368f
C763 VTAIL.n119 VSUBS 1.05995f
C764 VTAIL.n120 VSUBS 0.033337f
C765 VTAIL.n121 VSUBS 0.029212f
C766 VTAIL.n122 VSUBS 0.015697f
C767 VTAIL.n123 VSUBS 0.027827f
C768 VTAIL.n124 VSUBS 0.02727f
C769 VTAIL.t10 VSUBS 0.085653f
C770 VTAIL.n125 VSUBS 0.118183f
C771 VTAIL.n126 VSUBS 0.325467f
C772 VTAIL.n127 VSUBS 0.015697f
C773 VTAIL.n128 VSUBS 0.01662f
C774 VTAIL.n129 VSUBS 0.037102f
C775 VTAIL.n130 VSUBS 0.094044f
C776 VTAIL.n131 VSUBS 0.01662f
C777 VTAIL.n132 VSUBS 0.015697f
C778 VTAIL.n133 VSUBS 0.06393f
C779 VTAIL.n134 VSUBS 0.047368f
C780 VTAIL.n135 VSUBS 1.05447f
C781 VDD2.t4 VSUBS 0.064909f
C782 VDD2.t1 VSUBS 0.064909f
C783 VDD2.n0 VSUBS 0.347651f
C784 VDD2.t5 VSUBS 0.064909f
C785 VDD2.t2 VSUBS 0.064909f
C786 VDD2.n1 VSUBS 0.347651f
C787 VDD2.n2 VSUBS 2.56594f
C788 VDD2.t6 VSUBS 0.064909f
C789 VDD2.t7 VSUBS 0.064909f
C790 VDD2.n3 VSUBS 0.343591f
C791 VDD2.n4 VSUBS 2.11281f
C792 VDD2.t0 VSUBS 0.064909f
C793 VDD2.t3 VSUBS 0.064909f
C794 VDD2.n5 VSUBS 0.347634f
C795 VN.n0 VSUBS 0.064492f
C796 VN.t5 VSUBS 0.804541f
C797 VN.n1 VSUBS 0.07141f
C798 VN.n2 VSUBS 0.048917f
C799 VN.t1 VSUBS 0.804541f
C800 VN.n3 VSUBS 0.039545f
C801 VN.n4 VSUBS 0.362451f
C802 VN.t4 VSUBS 0.804541f
C803 VN.t0 VSUBS 1.04088f
C804 VN.n5 VSUBS 0.454941f
C805 VN.n6 VSUBS 0.445205f
C806 VN.n7 VSUBS 0.057408f
C807 VN.n8 VSUBS 0.097222f
C808 VN.n9 VSUBS 0.048917f
C809 VN.n10 VSUBS 0.048917f
C810 VN.n11 VSUBS 0.048917f
C811 VN.n12 VSUBS 0.097222f
C812 VN.n13 VSUBS 0.057408f
C813 VN.n14 VSUBS 0.342432f
C814 VN.n15 VSUBS 0.079914f
C815 VN.n16 VSUBS 0.048917f
C816 VN.n17 VSUBS 0.048917f
C817 VN.n18 VSUBS 0.048917f
C818 VN.n19 VSUBS 0.07141f
C819 VN.n20 VSUBS 0.079914f
C820 VN.n21 VSUBS 0.482369f
C821 VN.n22 VSUBS 0.060623f
C822 VN.n23 VSUBS 0.064492f
C823 VN.t2 VSUBS 0.804541f
C824 VN.n24 VSUBS 0.07141f
C825 VN.n25 VSUBS 0.048917f
C826 VN.t6 VSUBS 0.804541f
C827 VN.n26 VSUBS 0.039545f
C828 VN.n27 VSUBS 0.362451f
C829 VN.t7 VSUBS 0.804541f
C830 VN.t3 VSUBS 1.04088f
C831 VN.n28 VSUBS 0.454941f
C832 VN.n29 VSUBS 0.445205f
C833 VN.n30 VSUBS 0.057408f
C834 VN.n31 VSUBS 0.097222f
C835 VN.n32 VSUBS 0.048917f
C836 VN.n33 VSUBS 0.048917f
C837 VN.n34 VSUBS 0.048917f
C838 VN.n35 VSUBS 0.097222f
C839 VN.n36 VSUBS 0.057408f
C840 VN.n37 VSUBS 0.342432f
C841 VN.n38 VSUBS 0.079914f
C842 VN.n39 VSUBS 0.048917f
C843 VN.n40 VSUBS 0.048917f
C844 VN.n41 VSUBS 0.048917f
C845 VN.n42 VSUBS 0.07141f
C846 VN.n43 VSUBS 0.079914f
C847 VN.n44 VSUBS 0.482369f
C848 VN.n45 VSUBS 2.02119f
.ends

