* NGSPICE file created from diff_pair_sample_1769.ext - technology: sky130A

.subckt diff_pair_sample_1769 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t11 VN.t0 VDD2.t0 w_n3810_n1262# sky130_fd_pr__pfet_01v8 ad=0.24255 pd=1.8 as=0.24255 ps=1.8 w=1.47 l=3.22
X1 VDD1.t5 VP.t0 VTAIL.t4 w_n3810_n1262# sky130_fd_pr__pfet_01v8 ad=0.5733 pd=3.72 as=0.24255 ps=1.8 w=1.47 l=3.22
X2 B.t11 B.t9 B.t10 w_n3810_n1262# sky130_fd_pr__pfet_01v8 ad=0.5733 pd=3.72 as=0 ps=0 w=1.47 l=3.22
X3 B.t8 B.t6 B.t7 w_n3810_n1262# sky130_fd_pr__pfet_01v8 ad=0.5733 pd=3.72 as=0 ps=0 w=1.47 l=3.22
X4 VDD2.t1 VN.t1 VTAIL.t10 w_n3810_n1262# sky130_fd_pr__pfet_01v8 ad=0.24255 pd=1.8 as=0.5733 ps=3.72 w=1.47 l=3.22
X5 VDD1.t4 VP.t1 VTAIL.t5 w_n3810_n1262# sky130_fd_pr__pfet_01v8 ad=0.24255 pd=1.8 as=0.5733 ps=3.72 w=1.47 l=3.22
X6 VDD2.t4 VN.t2 VTAIL.t9 w_n3810_n1262# sky130_fd_pr__pfet_01v8 ad=0.5733 pd=3.72 as=0.24255 ps=1.8 w=1.47 l=3.22
X7 VTAIL.t8 VN.t3 VDD2.t5 w_n3810_n1262# sky130_fd_pr__pfet_01v8 ad=0.24255 pd=1.8 as=0.24255 ps=1.8 w=1.47 l=3.22
X8 VDD2.t3 VN.t4 VTAIL.t7 w_n3810_n1262# sky130_fd_pr__pfet_01v8 ad=0.24255 pd=1.8 as=0.5733 ps=3.72 w=1.47 l=3.22
X9 B.t5 B.t3 B.t4 w_n3810_n1262# sky130_fd_pr__pfet_01v8 ad=0.5733 pd=3.72 as=0 ps=0 w=1.47 l=3.22
X10 B.t2 B.t0 B.t1 w_n3810_n1262# sky130_fd_pr__pfet_01v8 ad=0.5733 pd=3.72 as=0 ps=0 w=1.47 l=3.22
X11 VTAIL.t3 VP.t2 VDD1.t3 w_n3810_n1262# sky130_fd_pr__pfet_01v8 ad=0.24255 pd=1.8 as=0.24255 ps=1.8 w=1.47 l=3.22
X12 VDD2.t2 VN.t5 VTAIL.t6 w_n3810_n1262# sky130_fd_pr__pfet_01v8 ad=0.5733 pd=3.72 as=0.24255 ps=1.8 w=1.47 l=3.22
X13 VDD1.t2 VP.t3 VTAIL.t2 w_n3810_n1262# sky130_fd_pr__pfet_01v8 ad=0.24255 pd=1.8 as=0.5733 ps=3.72 w=1.47 l=3.22
X14 VTAIL.t0 VP.t4 VDD1.t1 w_n3810_n1262# sky130_fd_pr__pfet_01v8 ad=0.24255 pd=1.8 as=0.24255 ps=1.8 w=1.47 l=3.22
X15 VDD1.t0 VP.t5 VTAIL.t1 w_n3810_n1262# sky130_fd_pr__pfet_01v8 ad=0.5733 pd=3.72 as=0.24255 ps=1.8 w=1.47 l=3.22
R0 VN.n34 VN.n33 161.3
R1 VN.n32 VN.n19 161.3
R2 VN.n31 VN.n30 161.3
R3 VN.n29 VN.n20 161.3
R4 VN.n28 VN.n27 161.3
R5 VN.n26 VN.n21 161.3
R6 VN.n25 VN.n24 161.3
R7 VN.n16 VN.n15 161.3
R8 VN.n14 VN.n1 161.3
R9 VN.n13 VN.n12 161.3
R10 VN.n11 VN.n2 161.3
R11 VN.n10 VN.n9 161.3
R12 VN.n8 VN.n3 161.3
R13 VN.n7 VN.n6 161.3
R14 VN.n17 VN.n0 75.3872
R15 VN.n35 VN.n18 75.3872
R16 VN.n5 VN.n4 62.0451
R17 VN.n23 VN.n22 62.0451
R18 VN.n5 VN.t2 43.9548
R19 VN.n23 VN.t1 43.9548
R20 VN VN.n35 43.3882
R21 VN.n13 VN.n2 42.9216
R22 VN.n31 VN.n20 42.9216
R23 VN.n9 VN.n2 38.0652
R24 VN.n27 VN.n20 38.0652
R25 VN.n8 VN.n7 24.4675
R26 VN.n9 VN.n8 24.4675
R27 VN.n14 VN.n13 24.4675
R28 VN.n15 VN.n14 24.4675
R29 VN.n27 VN.n26 24.4675
R30 VN.n26 VN.n25 24.4675
R31 VN.n33 VN.n32 24.4675
R32 VN.n32 VN.n31 24.4675
R33 VN.n15 VN.n0 14.6807
R34 VN.n33 VN.n18 14.6807
R35 VN.n7 VN.n4 12.234
R36 VN.n25 VN.n22 12.234
R37 VN.n4 VN.t3 11.0027
R38 VN.n0 VN.t4 11.0027
R39 VN.n22 VN.t0 11.0027
R40 VN.n18 VN.t5 11.0027
R41 VN.n6 VN.n5 4.15861
R42 VN.n24 VN.n23 4.15861
R43 VN.n35 VN.n34 0.354971
R44 VN.n17 VN.n16 0.354971
R45 VN VN.n17 0.26696
R46 VN.n34 VN.n19 0.189894
R47 VN.n30 VN.n19 0.189894
R48 VN.n30 VN.n29 0.189894
R49 VN.n29 VN.n28 0.189894
R50 VN.n28 VN.n21 0.189894
R51 VN.n24 VN.n21 0.189894
R52 VN.n6 VN.n3 0.189894
R53 VN.n10 VN.n3 0.189894
R54 VN.n11 VN.n10 0.189894
R55 VN.n12 VN.n11 0.189894
R56 VN.n12 VN.n1 0.189894
R57 VN.n16 VN.n1 0.189894
R58 VDD2.n1 VDD2.t4 274.723
R59 VDD2.n2 VDD2.t2 272.483
R60 VDD2.n1 VDD2.n0 251.081
R61 VDD2 VDD2.n3 251.077
R62 VDD2.n2 VDD2.n1 34.9287
R63 VDD2.n3 VDD2.t0 22.1127
R64 VDD2.n3 VDD2.t1 22.1127
R65 VDD2.n0 VDD2.t5 22.1127
R66 VDD2.n0 VDD2.t3 22.1127
R67 VDD2 VDD2.n2 2.35395
R68 VTAIL.n7 VTAIL.t10 255.804
R69 VTAIL.n11 VTAIL.t7 255.804
R70 VTAIL.n2 VTAIL.t2 255.804
R71 VTAIL.n10 VTAIL.t5 255.804
R72 VTAIL.n9 VTAIL.n8 233.691
R73 VTAIL.n6 VTAIL.n5 233.691
R74 VTAIL.n1 VTAIL.n0 233.691
R75 VTAIL.n4 VTAIL.n3 233.691
R76 VTAIL.n0 VTAIL.t9 22.1127
R77 VTAIL.n0 VTAIL.t8 22.1127
R78 VTAIL.n3 VTAIL.t1 22.1127
R79 VTAIL.n3 VTAIL.t0 22.1127
R80 VTAIL.n8 VTAIL.t4 22.1127
R81 VTAIL.n8 VTAIL.t3 22.1127
R82 VTAIL.n5 VTAIL.t6 22.1127
R83 VTAIL.n5 VTAIL.t11 22.1127
R84 VTAIL.n6 VTAIL.n4 19.7548
R85 VTAIL.n11 VTAIL.n10 16.6945
R86 VTAIL.n7 VTAIL.n6 3.06084
R87 VTAIL.n10 VTAIL.n9 3.06084
R88 VTAIL.n4 VTAIL.n2 3.06084
R89 VTAIL VTAIL.n11 2.23757
R90 VTAIL.n9 VTAIL.n7 2.0005
R91 VTAIL.n2 VTAIL.n1 2.0005
R92 VTAIL VTAIL.n1 0.823776
R93 VP.n16 VP.n15 161.3
R94 VP.n17 VP.n12 161.3
R95 VP.n19 VP.n18 161.3
R96 VP.n20 VP.n11 161.3
R97 VP.n22 VP.n21 161.3
R98 VP.n23 VP.n10 161.3
R99 VP.n25 VP.n24 161.3
R100 VP.n49 VP.n48 161.3
R101 VP.n47 VP.n1 161.3
R102 VP.n46 VP.n45 161.3
R103 VP.n44 VP.n2 161.3
R104 VP.n43 VP.n42 161.3
R105 VP.n41 VP.n3 161.3
R106 VP.n40 VP.n39 161.3
R107 VP.n38 VP.n37 161.3
R108 VP.n36 VP.n5 161.3
R109 VP.n35 VP.n34 161.3
R110 VP.n33 VP.n6 161.3
R111 VP.n32 VP.n31 161.3
R112 VP.n30 VP.n7 161.3
R113 VP.n29 VP.n28 161.3
R114 VP.n27 VP.n8 75.3872
R115 VP.n50 VP.n0 75.3872
R116 VP.n26 VP.n9 75.3872
R117 VP.n14 VP.n13 62.0451
R118 VP.n14 VP.t0 43.9546
R119 VP.n27 VP.n26 43.2228
R120 VP.n31 VP.n6 42.9216
R121 VP.n46 VP.n2 42.9216
R122 VP.n22 VP.n11 42.9216
R123 VP.n35 VP.n6 38.0652
R124 VP.n42 VP.n2 38.0652
R125 VP.n18 VP.n11 38.0652
R126 VP.n30 VP.n29 24.4675
R127 VP.n31 VP.n30 24.4675
R128 VP.n36 VP.n35 24.4675
R129 VP.n37 VP.n36 24.4675
R130 VP.n41 VP.n40 24.4675
R131 VP.n42 VP.n41 24.4675
R132 VP.n47 VP.n46 24.4675
R133 VP.n48 VP.n47 24.4675
R134 VP.n23 VP.n22 24.4675
R135 VP.n24 VP.n23 24.4675
R136 VP.n17 VP.n16 24.4675
R137 VP.n18 VP.n17 24.4675
R138 VP.n29 VP.n8 14.6807
R139 VP.n48 VP.n0 14.6807
R140 VP.n24 VP.n9 14.6807
R141 VP.n37 VP.n4 12.234
R142 VP.n40 VP.n4 12.234
R143 VP.n16 VP.n13 12.234
R144 VP.n8 VP.t5 11.0027
R145 VP.n4 VP.t4 11.0027
R146 VP.n0 VP.t3 11.0027
R147 VP.n9 VP.t1 11.0027
R148 VP.n13 VP.t2 11.0027
R149 VP.n15 VP.n14 4.15859
R150 VP.n26 VP.n25 0.354971
R151 VP.n28 VP.n27 0.354971
R152 VP.n50 VP.n49 0.354971
R153 VP VP.n50 0.26696
R154 VP.n15 VP.n12 0.189894
R155 VP.n19 VP.n12 0.189894
R156 VP.n20 VP.n19 0.189894
R157 VP.n21 VP.n20 0.189894
R158 VP.n21 VP.n10 0.189894
R159 VP.n25 VP.n10 0.189894
R160 VP.n28 VP.n7 0.189894
R161 VP.n32 VP.n7 0.189894
R162 VP.n33 VP.n32 0.189894
R163 VP.n34 VP.n33 0.189894
R164 VP.n34 VP.n5 0.189894
R165 VP.n38 VP.n5 0.189894
R166 VP.n39 VP.n38 0.189894
R167 VP.n39 VP.n3 0.189894
R168 VP.n43 VP.n3 0.189894
R169 VP.n44 VP.n43 0.189894
R170 VP.n45 VP.n44 0.189894
R171 VP.n45 VP.n1 0.189894
R172 VP.n49 VP.n1 0.189894
R173 VDD1 VDD1.t5 274.837
R174 VDD1.n1 VDD1.t0 274.723
R175 VDD1.n1 VDD1.n0 251.081
R176 VDD1.n3 VDD1.n2 250.37
R177 VDD1.n3 VDD1.n1 37.0418
R178 VDD1.n2 VDD1.t3 22.1127
R179 VDD1.n2 VDD1.t4 22.1127
R180 VDD1.n0 VDD1.t1 22.1127
R181 VDD1.n0 VDD1.t2 22.1127
R182 VDD1 VDD1.n3 0.707397
R183 B.n416 B.n47 585
R184 B.n418 B.n417 585
R185 B.n419 B.n46 585
R186 B.n421 B.n420 585
R187 B.n422 B.n45 585
R188 B.n424 B.n423 585
R189 B.n425 B.n44 585
R190 B.n427 B.n426 585
R191 B.n428 B.n43 585
R192 B.n430 B.n429 585
R193 B.n431 B.n40 585
R194 B.n434 B.n433 585
R195 B.n435 B.n39 585
R196 B.n437 B.n436 585
R197 B.n438 B.n38 585
R198 B.n440 B.n439 585
R199 B.n441 B.n37 585
R200 B.n443 B.n442 585
R201 B.n444 B.n33 585
R202 B.n446 B.n445 585
R203 B.n447 B.n32 585
R204 B.n449 B.n448 585
R205 B.n450 B.n31 585
R206 B.n452 B.n451 585
R207 B.n453 B.n30 585
R208 B.n455 B.n454 585
R209 B.n456 B.n29 585
R210 B.n458 B.n457 585
R211 B.n459 B.n28 585
R212 B.n461 B.n460 585
R213 B.n462 B.n27 585
R214 B.n415 B.n414 585
R215 B.n413 B.n48 585
R216 B.n412 B.n411 585
R217 B.n410 B.n49 585
R218 B.n409 B.n408 585
R219 B.n407 B.n50 585
R220 B.n406 B.n405 585
R221 B.n404 B.n51 585
R222 B.n403 B.n402 585
R223 B.n401 B.n52 585
R224 B.n400 B.n399 585
R225 B.n398 B.n53 585
R226 B.n397 B.n396 585
R227 B.n395 B.n54 585
R228 B.n394 B.n393 585
R229 B.n392 B.n55 585
R230 B.n391 B.n390 585
R231 B.n389 B.n56 585
R232 B.n388 B.n387 585
R233 B.n386 B.n57 585
R234 B.n385 B.n384 585
R235 B.n383 B.n58 585
R236 B.n382 B.n381 585
R237 B.n380 B.n59 585
R238 B.n379 B.n378 585
R239 B.n377 B.n60 585
R240 B.n376 B.n375 585
R241 B.n374 B.n61 585
R242 B.n373 B.n372 585
R243 B.n371 B.n62 585
R244 B.n370 B.n369 585
R245 B.n368 B.n63 585
R246 B.n367 B.n366 585
R247 B.n365 B.n64 585
R248 B.n364 B.n363 585
R249 B.n362 B.n65 585
R250 B.n361 B.n360 585
R251 B.n359 B.n66 585
R252 B.n358 B.n357 585
R253 B.n356 B.n67 585
R254 B.n355 B.n354 585
R255 B.n353 B.n68 585
R256 B.n352 B.n351 585
R257 B.n350 B.n69 585
R258 B.n349 B.n348 585
R259 B.n347 B.n70 585
R260 B.n346 B.n345 585
R261 B.n344 B.n71 585
R262 B.n343 B.n342 585
R263 B.n341 B.n72 585
R264 B.n340 B.n339 585
R265 B.n338 B.n73 585
R266 B.n337 B.n336 585
R267 B.n335 B.n74 585
R268 B.n334 B.n333 585
R269 B.n332 B.n75 585
R270 B.n331 B.n330 585
R271 B.n329 B.n76 585
R272 B.n328 B.n327 585
R273 B.n326 B.n77 585
R274 B.n325 B.n324 585
R275 B.n323 B.n78 585
R276 B.n322 B.n321 585
R277 B.n320 B.n79 585
R278 B.n319 B.n318 585
R279 B.n317 B.n80 585
R280 B.n316 B.n315 585
R281 B.n314 B.n81 585
R282 B.n313 B.n312 585
R283 B.n311 B.n82 585
R284 B.n310 B.n309 585
R285 B.n308 B.n83 585
R286 B.n307 B.n306 585
R287 B.n305 B.n84 585
R288 B.n304 B.n303 585
R289 B.n302 B.n85 585
R290 B.n301 B.n300 585
R291 B.n299 B.n86 585
R292 B.n298 B.n297 585
R293 B.n296 B.n87 585
R294 B.n295 B.n294 585
R295 B.n293 B.n88 585
R296 B.n292 B.n291 585
R297 B.n290 B.n89 585
R298 B.n289 B.n288 585
R299 B.n287 B.n90 585
R300 B.n286 B.n285 585
R301 B.n284 B.n91 585
R302 B.n283 B.n282 585
R303 B.n281 B.n92 585
R304 B.n280 B.n279 585
R305 B.n278 B.n93 585
R306 B.n277 B.n276 585
R307 B.n275 B.n94 585
R308 B.n274 B.n273 585
R309 B.n272 B.n95 585
R310 B.n271 B.n270 585
R311 B.n269 B.n96 585
R312 B.n268 B.n267 585
R313 B.n266 B.n97 585
R314 B.n265 B.n264 585
R315 B.n214 B.n115 585
R316 B.n216 B.n215 585
R317 B.n217 B.n114 585
R318 B.n219 B.n218 585
R319 B.n220 B.n113 585
R320 B.n222 B.n221 585
R321 B.n223 B.n112 585
R322 B.n225 B.n224 585
R323 B.n226 B.n111 585
R324 B.n228 B.n227 585
R325 B.n229 B.n108 585
R326 B.n232 B.n231 585
R327 B.n233 B.n107 585
R328 B.n235 B.n234 585
R329 B.n236 B.n106 585
R330 B.n238 B.n237 585
R331 B.n239 B.n105 585
R332 B.n241 B.n240 585
R333 B.n242 B.n104 585
R334 B.n247 B.n246 585
R335 B.n248 B.n103 585
R336 B.n250 B.n249 585
R337 B.n251 B.n102 585
R338 B.n253 B.n252 585
R339 B.n254 B.n101 585
R340 B.n256 B.n255 585
R341 B.n257 B.n100 585
R342 B.n259 B.n258 585
R343 B.n260 B.n99 585
R344 B.n262 B.n261 585
R345 B.n263 B.n98 585
R346 B.n213 B.n212 585
R347 B.n211 B.n116 585
R348 B.n210 B.n209 585
R349 B.n208 B.n117 585
R350 B.n207 B.n206 585
R351 B.n205 B.n118 585
R352 B.n204 B.n203 585
R353 B.n202 B.n119 585
R354 B.n201 B.n200 585
R355 B.n199 B.n120 585
R356 B.n198 B.n197 585
R357 B.n196 B.n121 585
R358 B.n195 B.n194 585
R359 B.n193 B.n122 585
R360 B.n192 B.n191 585
R361 B.n190 B.n123 585
R362 B.n189 B.n188 585
R363 B.n187 B.n124 585
R364 B.n186 B.n185 585
R365 B.n184 B.n125 585
R366 B.n183 B.n182 585
R367 B.n181 B.n126 585
R368 B.n180 B.n179 585
R369 B.n178 B.n127 585
R370 B.n177 B.n176 585
R371 B.n175 B.n128 585
R372 B.n174 B.n173 585
R373 B.n172 B.n129 585
R374 B.n171 B.n170 585
R375 B.n169 B.n130 585
R376 B.n168 B.n167 585
R377 B.n166 B.n131 585
R378 B.n165 B.n164 585
R379 B.n163 B.n132 585
R380 B.n162 B.n161 585
R381 B.n160 B.n133 585
R382 B.n159 B.n158 585
R383 B.n157 B.n134 585
R384 B.n156 B.n155 585
R385 B.n154 B.n135 585
R386 B.n153 B.n152 585
R387 B.n151 B.n136 585
R388 B.n150 B.n149 585
R389 B.n148 B.n137 585
R390 B.n147 B.n146 585
R391 B.n145 B.n138 585
R392 B.n144 B.n143 585
R393 B.n142 B.n139 585
R394 B.n141 B.n140 585
R395 B.n2 B.n0 585
R396 B.n537 B.n1 585
R397 B.n536 B.n535 585
R398 B.n534 B.n3 585
R399 B.n533 B.n532 585
R400 B.n531 B.n4 585
R401 B.n530 B.n529 585
R402 B.n528 B.n5 585
R403 B.n527 B.n526 585
R404 B.n525 B.n6 585
R405 B.n524 B.n523 585
R406 B.n522 B.n7 585
R407 B.n521 B.n520 585
R408 B.n519 B.n8 585
R409 B.n518 B.n517 585
R410 B.n516 B.n9 585
R411 B.n515 B.n514 585
R412 B.n513 B.n10 585
R413 B.n512 B.n511 585
R414 B.n510 B.n11 585
R415 B.n509 B.n508 585
R416 B.n507 B.n12 585
R417 B.n506 B.n505 585
R418 B.n504 B.n13 585
R419 B.n503 B.n502 585
R420 B.n501 B.n14 585
R421 B.n500 B.n499 585
R422 B.n498 B.n15 585
R423 B.n497 B.n496 585
R424 B.n495 B.n16 585
R425 B.n494 B.n493 585
R426 B.n492 B.n17 585
R427 B.n491 B.n490 585
R428 B.n489 B.n18 585
R429 B.n488 B.n487 585
R430 B.n486 B.n19 585
R431 B.n485 B.n484 585
R432 B.n483 B.n20 585
R433 B.n482 B.n481 585
R434 B.n480 B.n21 585
R435 B.n479 B.n478 585
R436 B.n477 B.n22 585
R437 B.n476 B.n475 585
R438 B.n474 B.n23 585
R439 B.n473 B.n472 585
R440 B.n471 B.n24 585
R441 B.n470 B.n469 585
R442 B.n468 B.n25 585
R443 B.n467 B.n466 585
R444 B.n465 B.n26 585
R445 B.n464 B.n463 585
R446 B.n539 B.n538 585
R447 B.n214 B.n213 468.476
R448 B.n464 B.n27 468.476
R449 B.n265 B.n98 468.476
R450 B.n416 B.n415 468.476
R451 B.n243 B.t5 318.156
R452 B.n41 B.t7 318.156
R453 B.n109 B.t2 318.156
R454 B.n34 B.t10 318.156
R455 B.n244 B.t4 249.309
R456 B.n42 B.t8 249.309
R457 B.n110 B.t1 249.308
R458 B.n35 B.t11 249.308
R459 B.n243 B.t3 209.363
R460 B.n109 B.t0 209.363
R461 B.n34 B.t9 209.363
R462 B.n41 B.t6 209.363
R463 B.n213 B.n116 163.367
R464 B.n209 B.n116 163.367
R465 B.n209 B.n208 163.367
R466 B.n208 B.n207 163.367
R467 B.n207 B.n118 163.367
R468 B.n203 B.n118 163.367
R469 B.n203 B.n202 163.367
R470 B.n202 B.n201 163.367
R471 B.n201 B.n120 163.367
R472 B.n197 B.n120 163.367
R473 B.n197 B.n196 163.367
R474 B.n196 B.n195 163.367
R475 B.n195 B.n122 163.367
R476 B.n191 B.n122 163.367
R477 B.n191 B.n190 163.367
R478 B.n190 B.n189 163.367
R479 B.n189 B.n124 163.367
R480 B.n185 B.n124 163.367
R481 B.n185 B.n184 163.367
R482 B.n184 B.n183 163.367
R483 B.n183 B.n126 163.367
R484 B.n179 B.n126 163.367
R485 B.n179 B.n178 163.367
R486 B.n178 B.n177 163.367
R487 B.n177 B.n128 163.367
R488 B.n173 B.n128 163.367
R489 B.n173 B.n172 163.367
R490 B.n172 B.n171 163.367
R491 B.n171 B.n130 163.367
R492 B.n167 B.n130 163.367
R493 B.n167 B.n166 163.367
R494 B.n166 B.n165 163.367
R495 B.n165 B.n132 163.367
R496 B.n161 B.n132 163.367
R497 B.n161 B.n160 163.367
R498 B.n160 B.n159 163.367
R499 B.n159 B.n134 163.367
R500 B.n155 B.n134 163.367
R501 B.n155 B.n154 163.367
R502 B.n154 B.n153 163.367
R503 B.n153 B.n136 163.367
R504 B.n149 B.n136 163.367
R505 B.n149 B.n148 163.367
R506 B.n148 B.n147 163.367
R507 B.n147 B.n138 163.367
R508 B.n143 B.n138 163.367
R509 B.n143 B.n142 163.367
R510 B.n142 B.n141 163.367
R511 B.n141 B.n2 163.367
R512 B.n538 B.n2 163.367
R513 B.n538 B.n537 163.367
R514 B.n537 B.n536 163.367
R515 B.n536 B.n3 163.367
R516 B.n532 B.n3 163.367
R517 B.n532 B.n531 163.367
R518 B.n531 B.n530 163.367
R519 B.n530 B.n5 163.367
R520 B.n526 B.n5 163.367
R521 B.n526 B.n525 163.367
R522 B.n525 B.n524 163.367
R523 B.n524 B.n7 163.367
R524 B.n520 B.n7 163.367
R525 B.n520 B.n519 163.367
R526 B.n519 B.n518 163.367
R527 B.n518 B.n9 163.367
R528 B.n514 B.n9 163.367
R529 B.n514 B.n513 163.367
R530 B.n513 B.n512 163.367
R531 B.n512 B.n11 163.367
R532 B.n508 B.n11 163.367
R533 B.n508 B.n507 163.367
R534 B.n507 B.n506 163.367
R535 B.n506 B.n13 163.367
R536 B.n502 B.n13 163.367
R537 B.n502 B.n501 163.367
R538 B.n501 B.n500 163.367
R539 B.n500 B.n15 163.367
R540 B.n496 B.n15 163.367
R541 B.n496 B.n495 163.367
R542 B.n495 B.n494 163.367
R543 B.n494 B.n17 163.367
R544 B.n490 B.n17 163.367
R545 B.n490 B.n489 163.367
R546 B.n489 B.n488 163.367
R547 B.n488 B.n19 163.367
R548 B.n484 B.n19 163.367
R549 B.n484 B.n483 163.367
R550 B.n483 B.n482 163.367
R551 B.n482 B.n21 163.367
R552 B.n478 B.n21 163.367
R553 B.n478 B.n477 163.367
R554 B.n477 B.n476 163.367
R555 B.n476 B.n23 163.367
R556 B.n472 B.n23 163.367
R557 B.n472 B.n471 163.367
R558 B.n471 B.n470 163.367
R559 B.n470 B.n25 163.367
R560 B.n466 B.n25 163.367
R561 B.n466 B.n465 163.367
R562 B.n465 B.n464 163.367
R563 B.n215 B.n214 163.367
R564 B.n215 B.n114 163.367
R565 B.n219 B.n114 163.367
R566 B.n220 B.n219 163.367
R567 B.n221 B.n220 163.367
R568 B.n221 B.n112 163.367
R569 B.n225 B.n112 163.367
R570 B.n226 B.n225 163.367
R571 B.n227 B.n226 163.367
R572 B.n227 B.n108 163.367
R573 B.n232 B.n108 163.367
R574 B.n233 B.n232 163.367
R575 B.n234 B.n233 163.367
R576 B.n234 B.n106 163.367
R577 B.n238 B.n106 163.367
R578 B.n239 B.n238 163.367
R579 B.n240 B.n239 163.367
R580 B.n240 B.n104 163.367
R581 B.n247 B.n104 163.367
R582 B.n248 B.n247 163.367
R583 B.n249 B.n248 163.367
R584 B.n249 B.n102 163.367
R585 B.n253 B.n102 163.367
R586 B.n254 B.n253 163.367
R587 B.n255 B.n254 163.367
R588 B.n255 B.n100 163.367
R589 B.n259 B.n100 163.367
R590 B.n260 B.n259 163.367
R591 B.n261 B.n260 163.367
R592 B.n261 B.n98 163.367
R593 B.n266 B.n265 163.367
R594 B.n267 B.n266 163.367
R595 B.n267 B.n96 163.367
R596 B.n271 B.n96 163.367
R597 B.n272 B.n271 163.367
R598 B.n273 B.n272 163.367
R599 B.n273 B.n94 163.367
R600 B.n277 B.n94 163.367
R601 B.n278 B.n277 163.367
R602 B.n279 B.n278 163.367
R603 B.n279 B.n92 163.367
R604 B.n283 B.n92 163.367
R605 B.n284 B.n283 163.367
R606 B.n285 B.n284 163.367
R607 B.n285 B.n90 163.367
R608 B.n289 B.n90 163.367
R609 B.n290 B.n289 163.367
R610 B.n291 B.n290 163.367
R611 B.n291 B.n88 163.367
R612 B.n295 B.n88 163.367
R613 B.n296 B.n295 163.367
R614 B.n297 B.n296 163.367
R615 B.n297 B.n86 163.367
R616 B.n301 B.n86 163.367
R617 B.n302 B.n301 163.367
R618 B.n303 B.n302 163.367
R619 B.n303 B.n84 163.367
R620 B.n307 B.n84 163.367
R621 B.n308 B.n307 163.367
R622 B.n309 B.n308 163.367
R623 B.n309 B.n82 163.367
R624 B.n313 B.n82 163.367
R625 B.n314 B.n313 163.367
R626 B.n315 B.n314 163.367
R627 B.n315 B.n80 163.367
R628 B.n319 B.n80 163.367
R629 B.n320 B.n319 163.367
R630 B.n321 B.n320 163.367
R631 B.n321 B.n78 163.367
R632 B.n325 B.n78 163.367
R633 B.n326 B.n325 163.367
R634 B.n327 B.n326 163.367
R635 B.n327 B.n76 163.367
R636 B.n331 B.n76 163.367
R637 B.n332 B.n331 163.367
R638 B.n333 B.n332 163.367
R639 B.n333 B.n74 163.367
R640 B.n337 B.n74 163.367
R641 B.n338 B.n337 163.367
R642 B.n339 B.n338 163.367
R643 B.n339 B.n72 163.367
R644 B.n343 B.n72 163.367
R645 B.n344 B.n343 163.367
R646 B.n345 B.n344 163.367
R647 B.n345 B.n70 163.367
R648 B.n349 B.n70 163.367
R649 B.n350 B.n349 163.367
R650 B.n351 B.n350 163.367
R651 B.n351 B.n68 163.367
R652 B.n355 B.n68 163.367
R653 B.n356 B.n355 163.367
R654 B.n357 B.n356 163.367
R655 B.n357 B.n66 163.367
R656 B.n361 B.n66 163.367
R657 B.n362 B.n361 163.367
R658 B.n363 B.n362 163.367
R659 B.n363 B.n64 163.367
R660 B.n367 B.n64 163.367
R661 B.n368 B.n367 163.367
R662 B.n369 B.n368 163.367
R663 B.n369 B.n62 163.367
R664 B.n373 B.n62 163.367
R665 B.n374 B.n373 163.367
R666 B.n375 B.n374 163.367
R667 B.n375 B.n60 163.367
R668 B.n379 B.n60 163.367
R669 B.n380 B.n379 163.367
R670 B.n381 B.n380 163.367
R671 B.n381 B.n58 163.367
R672 B.n385 B.n58 163.367
R673 B.n386 B.n385 163.367
R674 B.n387 B.n386 163.367
R675 B.n387 B.n56 163.367
R676 B.n391 B.n56 163.367
R677 B.n392 B.n391 163.367
R678 B.n393 B.n392 163.367
R679 B.n393 B.n54 163.367
R680 B.n397 B.n54 163.367
R681 B.n398 B.n397 163.367
R682 B.n399 B.n398 163.367
R683 B.n399 B.n52 163.367
R684 B.n403 B.n52 163.367
R685 B.n404 B.n403 163.367
R686 B.n405 B.n404 163.367
R687 B.n405 B.n50 163.367
R688 B.n409 B.n50 163.367
R689 B.n410 B.n409 163.367
R690 B.n411 B.n410 163.367
R691 B.n411 B.n48 163.367
R692 B.n415 B.n48 163.367
R693 B.n460 B.n27 163.367
R694 B.n460 B.n459 163.367
R695 B.n459 B.n458 163.367
R696 B.n458 B.n29 163.367
R697 B.n454 B.n29 163.367
R698 B.n454 B.n453 163.367
R699 B.n453 B.n452 163.367
R700 B.n452 B.n31 163.367
R701 B.n448 B.n31 163.367
R702 B.n448 B.n447 163.367
R703 B.n447 B.n446 163.367
R704 B.n446 B.n33 163.367
R705 B.n442 B.n33 163.367
R706 B.n442 B.n441 163.367
R707 B.n441 B.n440 163.367
R708 B.n440 B.n38 163.367
R709 B.n436 B.n38 163.367
R710 B.n436 B.n435 163.367
R711 B.n435 B.n434 163.367
R712 B.n434 B.n40 163.367
R713 B.n429 B.n40 163.367
R714 B.n429 B.n428 163.367
R715 B.n428 B.n427 163.367
R716 B.n427 B.n44 163.367
R717 B.n423 B.n44 163.367
R718 B.n423 B.n422 163.367
R719 B.n422 B.n421 163.367
R720 B.n421 B.n46 163.367
R721 B.n417 B.n46 163.367
R722 B.n417 B.n416 163.367
R723 B.n244 B.n243 68.849
R724 B.n110 B.n109 68.849
R725 B.n35 B.n34 68.849
R726 B.n42 B.n41 68.849
R727 B.n245 B.n244 59.5399
R728 B.n230 B.n110 59.5399
R729 B.n36 B.n35 59.5399
R730 B.n432 B.n42 59.5399
R731 B.n463 B.n462 30.4395
R732 B.n414 B.n47 30.4395
R733 B.n264 B.n263 30.4395
R734 B.n212 B.n115 30.4395
R735 B B.n539 18.0485
R736 B.n462 B.n461 10.6151
R737 B.n461 B.n28 10.6151
R738 B.n457 B.n28 10.6151
R739 B.n457 B.n456 10.6151
R740 B.n456 B.n455 10.6151
R741 B.n455 B.n30 10.6151
R742 B.n451 B.n30 10.6151
R743 B.n451 B.n450 10.6151
R744 B.n450 B.n449 10.6151
R745 B.n449 B.n32 10.6151
R746 B.n445 B.n444 10.6151
R747 B.n444 B.n443 10.6151
R748 B.n443 B.n37 10.6151
R749 B.n439 B.n37 10.6151
R750 B.n439 B.n438 10.6151
R751 B.n438 B.n437 10.6151
R752 B.n437 B.n39 10.6151
R753 B.n433 B.n39 10.6151
R754 B.n431 B.n430 10.6151
R755 B.n430 B.n43 10.6151
R756 B.n426 B.n43 10.6151
R757 B.n426 B.n425 10.6151
R758 B.n425 B.n424 10.6151
R759 B.n424 B.n45 10.6151
R760 B.n420 B.n45 10.6151
R761 B.n420 B.n419 10.6151
R762 B.n419 B.n418 10.6151
R763 B.n418 B.n47 10.6151
R764 B.n264 B.n97 10.6151
R765 B.n268 B.n97 10.6151
R766 B.n269 B.n268 10.6151
R767 B.n270 B.n269 10.6151
R768 B.n270 B.n95 10.6151
R769 B.n274 B.n95 10.6151
R770 B.n275 B.n274 10.6151
R771 B.n276 B.n275 10.6151
R772 B.n276 B.n93 10.6151
R773 B.n280 B.n93 10.6151
R774 B.n281 B.n280 10.6151
R775 B.n282 B.n281 10.6151
R776 B.n282 B.n91 10.6151
R777 B.n286 B.n91 10.6151
R778 B.n287 B.n286 10.6151
R779 B.n288 B.n287 10.6151
R780 B.n288 B.n89 10.6151
R781 B.n292 B.n89 10.6151
R782 B.n293 B.n292 10.6151
R783 B.n294 B.n293 10.6151
R784 B.n294 B.n87 10.6151
R785 B.n298 B.n87 10.6151
R786 B.n299 B.n298 10.6151
R787 B.n300 B.n299 10.6151
R788 B.n300 B.n85 10.6151
R789 B.n304 B.n85 10.6151
R790 B.n305 B.n304 10.6151
R791 B.n306 B.n305 10.6151
R792 B.n306 B.n83 10.6151
R793 B.n310 B.n83 10.6151
R794 B.n311 B.n310 10.6151
R795 B.n312 B.n311 10.6151
R796 B.n312 B.n81 10.6151
R797 B.n316 B.n81 10.6151
R798 B.n317 B.n316 10.6151
R799 B.n318 B.n317 10.6151
R800 B.n318 B.n79 10.6151
R801 B.n322 B.n79 10.6151
R802 B.n323 B.n322 10.6151
R803 B.n324 B.n323 10.6151
R804 B.n324 B.n77 10.6151
R805 B.n328 B.n77 10.6151
R806 B.n329 B.n328 10.6151
R807 B.n330 B.n329 10.6151
R808 B.n330 B.n75 10.6151
R809 B.n334 B.n75 10.6151
R810 B.n335 B.n334 10.6151
R811 B.n336 B.n335 10.6151
R812 B.n336 B.n73 10.6151
R813 B.n340 B.n73 10.6151
R814 B.n341 B.n340 10.6151
R815 B.n342 B.n341 10.6151
R816 B.n342 B.n71 10.6151
R817 B.n346 B.n71 10.6151
R818 B.n347 B.n346 10.6151
R819 B.n348 B.n347 10.6151
R820 B.n348 B.n69 10.6151
R821 B.n352 B.n69 10.6151
R822 B.n353 B.n352 10.6151
R823 B.n354 B.n353 10.6151
R824 B.n354 B.n67 10.6151
R825 B.n358 B.n67 10.6151
R826 B.n359 B.n358 10.6151
R827 B.n360 B.n359 10.6151
R828 B.n360 B.n65 10.6151
R829 B.n364 B.n65 10.6151
R830 B.n365 B.n364 10.6151
R831 B.n366 B.n365 10.6151
R832 B.n366 B.n63 10.6151
R833 B.n370 B.n63 10.6151
R834 B.n371 B.n370 10.6151
R835 B.n372 B.n371 10.6151
R836 B.n372 B.n61 10.6151
R837 B.n376 B.n61 10.6151
R838 B.n377 B.n376 10.6151
R839 B.n378 B.n377 10.6151
R840 B.n378 B.n59 10.6151
R841 B.n382 B.n59 10.6151
R842 B.n383 B.n382 10.6151
R843 B.n384 B.n383 10.6151
R844 B.n384 B.n57 10.6151
R845 B.n388 B.n57 10.6151
R846 B.n389 B.n388 10.6151
R847 B.n390 B.n389 10.6151
R848 B.n390 B.n55 10.6151
R849 B.n394 B.n55 10.6151
R850 B.n395 B.n394 10.6151
R851 B.n396 B.n395 10.6151
R852 B.n396 B.n53 10.6151
R853 B.n400 B.n53 10.6151
R854 B.n401 B.n400 10.6151
R855 B.n402 B.n401 10.6151
R856 B.n402 B.n51 10.6151
R857 B.n406 B.n51 10.6151
R858 B.n407 B.n406 10.6151
R859 B.n408 B.n407 10.6151
R860 B.n408 B.n49 10.6151
R861 B.n412 B.n49 10.6151
R862 B.n413 B.n412 10.6151
R863 B.n414 B.n413 10.6151
R864 B.n216 B.n115 10.6151
R865 B.n217 B.n216 10.6151
R866 B.n218 B.n217 10.6151
R867 B.n218 B.n113 10.6151
R868 B.n222 B.n113 10.6151
R869 B.n223 B.n222 10.6151
R870 B.n224 B.n223 10.6151
R871 B.n224 B.n111 10.6151
R872 B.n228 B.n111 10.6151
R873 B.n229 B.n228 10.6151
R874 B.n231 B.n107 10.6151
R875 B.n235 B.n107 10.6151
R876 B.n236 B.n235 10.6151
R877 B.n237 B.n236 10.6151
R878 B.n237 B.n105 10.6151
R879 B.n241 B.n105 10.6151
R880 B.n242 B.n241 10.6151
R881 B.n246 B.n242 10.6151
R882 B.n250 B.n103 10.6151
R883 B.n251 B.n250 10.6151
R884 B.n252 B.n251 10.6151
R885 B.n252 B.n101 10.6151
R886 B.n256 B.n101 10.6151
R887 B.n257 B.n256 10.6151
R888 B.n258 B.n257 10.6151
R889 B.n258 B.n99 10.6151
R890 B.n262 B.n99 10.6151
R891 B.n263 B.n262 10.6151
R892 B.n212 B.n211 10.6151
R893 B.n211 B.n210 10.6151
R894 B.n210 B.n117 10.6151
R895 B.n206 B.n117 10.6151
R896 B.n206 B.n205 10.6151
R897 B.n205 B.n204 10.6151
R898 B.n204 B.n119 10.6151
R899 B.n200 B.n119 10.6151
R900 B.n200 B.n199 10.6151
R901 B.n199 B.n198 10.6151
R902 B.n198 B.n121 10.6151
R903 B.n194 B.n121 10.6151
R904 B.n194 B.n193 10.6151
R905 B.n193 B.n192 10.6151
R906 B.n192 B.n123 10.6151
R907 B.n188 B.n123 10.6151
R908 B.n188 B.n187 10.6151
R909 B.n187 B.n186 10.6151
R910 B.n186 B.n125 10.6151
R911 B.n182 B.n125 10.6151
R912 B.n182 B.n181 10.6151
R913 B.n181 B.n180 10.6151
R914 B.n180 B.n127 10.6151
R915 B.n176 B.n127 10.6151
R916 B.n176 B.n175 10.6151
R917 B.n175 B.n174 10.6151
R918 B.n174 B.n129 10.6151
R919 B.n170 B.n129 10.6151
R920 B.n170 B.n169 10.6151
R921 B.n169 B.n168 10.6151
R922 B.n168 B.n131 10.6151
R923 B.n164 B.n131 10.6151
R924 B.n164 B.n163 10.6151
R925 B.n163 B.n162 10.6151
R926 B.n162 B.n133 10.6151
R927 B.n158 B.n133 10.6151
R928 B.n158 B.n157 10.6151
R929 B.n157 B.n156 10.6151
R930 B.n156 B.n135 10.6151
R931 B.n152 B.n135 10.6151
R932 B.n152 B.n151 10.6151
R933 B.n151 B.n150 10.6151
R934 B.n150 B.n137 10.6151
R935 B.n146 B.n137 10.6151
R936 B.n146 B.n145 10.6151
R937 B.n145 B.n144 10.6151
R938 B.n144 B.n139 10.6151
R939 B.n140 B.n139 10.6151
R940 B.n140 B.n0 10.6151
R941 B.n535 B.n1 10.6151
R942 B.n535 B.n534 10.6151
R943 B.n534 B.n533 10.6151
R944 B.n533 B.n4 10.6151
R945 B.n529 B.n4 10.6151
R946 B.n529 B.n528 10.6151
R947 B.n528 B.n527 10.6151
R948 B.n527 B.n6 10.6151
R949 B.n523 B.n6 10.6151
R950 B.n523 B.n522 10.6151
R951 B.n522 B.n521 10.6151
R952 B.n521 B.n8 10.6151
R953 B.n517 B.n8 10.6151
R954 B.n517 B.n516 10.6151
R955 B.n516 B.n515 10.6151
R956 B.n515 B.n10 10.6151
R957 B.n511 B.n10 10.6151
R958 B.n511 B.n510 10.6151
R959 B.n510 B.n509 10.6151
R960 B.n509 B.n12 10.6151
R961 B.n505 B.n12 10.6151
R962 B.n505 B.n504 10.6151
R963 B.n504 B.n503 10.6151
R964 B.n503 B.n14 10.6151
R965 B.n499 B.n14 10.6151
R966 B.n499 B.n498 10.6151
R967 B.n498 B.n497 10.6151
R968 B.n497 B.n16 10.6151
R969 B.n493 B.n16 10.6151
R970 B.n493 B.n492 10.6151
R971 B.n492 B.n491 10.6151
R972 B.n491 B.n18 10.6151
R973 B.n487 B.n18 10.6151
R974 B.n487 B.n486 10.6151
R975 B.n486 B.n485 10.6151
R976 B.n485 B.n20 10.6151
R977 B.n481 B.n20 10.6151
R978 B.n481 B.n480 10.6151
R979 B.n480 B.n479 10.6151
R980 B.n479 B.n22 10.6151
R981 B.n475 B.n22 10.6151
R982 B.n475 B.n474 10.6151
R983 B.n474 B.n473 10.6151
R984 B.n473 B.n24 10.6151
R985 B.n469 B.n24 10.6151
R986 B.n469 B.n468 10.6151
R987 B.n468 B.n467 10.6151
R988 B.n467 B.n26 10.6151
R989 B.n463 B.n26 10.6151
R990 B.n445 B.n36 6.5566
R991 B.n433 B.n432 6.5566
R992 B.n231 B.n230 6.5566
R993 B.n246 B.n245 6.5566
R994 B.n36 B.n32 4.05904
R995 B.n432 B.n431 4.05904
R996 B.n230 B.n229 4.05904
R997 B.n245 B.n103 4.05904
R998 B.n539 B.n0 2.81026
R999 B.n539 B.n1 2.81026
C0 VDD1 VP 1.56828f
C1 VN VP 5.58981f
C2 VTAIL w_n3810_n1262# 1.52055f
C3 B VDD1 1.41116f
C4 VDD1 VDD2 1.64666f
C5 B VN 1.14238f
C6 VN VDD2 1.21157f
C7 VTAIL VP 2.3622f
C8 w_n3810_n1262# VP 7.6787f
C9 VTAIL B 1.33177f
C10 VTAIL VDD2 4.42507f
C11 B w_n3810_n1262# 7.65644f
C12 w_n3810_n1262# VDD2 1.81104f
C13 B VP 1.96981f
C14 VDD2 VP 0.518656f
C15 VN VDD1 0.158625f
C16 B VDD2 1.50067f
C17 VTAIL VDD1 4.36754f
C18 VTAIL VN 2.34808f
C19 w_n3810_n1262# VDD1 1.70705f
C20 w_n3810_n1262# VN 7.19065f
C21 VDD2 VSUBS 1.16161f
C22 VDD1 VSUBS 1.670686f
C23 VTAIL VSUBS 0.600287f
C24 VN VSUBS 6.58389f
C25 VP VSUBS 2.811989f
C26 B VSUBS 4.097774f
C27 w_n3810_n1262# VSUBS 61.676296f
C28 B.n0 VSUBS 0.006058f
C29 B.n1 VSUBS 0.006058f
C30 B.n2 VSUBS 0.009581f
C31 B.n3 VSUBS 0.009581f
C32 B.n4 VSUBS 0.009581f
C33 B.n5 VSUBS 0.009581f
C34 B.n6 VSUBS 0.009581f
C35 B.n7 VSUBS 0.009581f
C36 B.n8 VSUBS 0.009581f
C37 B.n9 VSUBS 0.009581f
C38 B.n10 VSUBS 0.009581f
C39 B.n11 VSUBS 0.009581f
C40 B.n12 VSUBS 0.009581f
C41 B.n13 VSUBS 0.009581f
C42 B.n14 VSUBS 0.009581f
C43 B.n15 VSUBS 0.009581f
C44 B.n16 VSUBS 0.009581f
C45 B.n17 VSUBS 0.009581f
C46 B.n18 VSUBS 0.009581f
C47 B.n19 VSUBS 0.009581f
C48 B.n20 VSUBS 0.009581f
C49 B.n21 VSUBS 0.009581f
C50 B.n22 VSUBS 0.009581f
C51 B.n23 VSUBS 0.009581f
C52 B.n24 VSUBS 0.009581f
C53 B.n25 VSUBS 0.009581f
C54 B.n26 VSUBS 0.009581f
C55 B.n27 VSUBS 0.021934f
C56 B.n28 VSUBS 0.009581f
C57 B.n29 VSUBS 0.009581f
C58 B.n30 VSUBS 0.009581f
C59 B.n31 VSUBS 0.009581f
C60 B.n32 VSUBS 0.006622f
C61 B.n33 VSUBS 0.009581f
C62 B.t11 VSUBS 0.040757f
C63 B.t10 VSUBS 0.054072f
C64 B.t9 VSUBS 0.326272f
C65 B.n34 VSUBS 0.095003f
C66 B.n35 VSUBS 0.075191f
C67 B.n36 VSUBS 0.022198f
C68 B.n37 VSUBS 0.009581f
C69 B.n38 VSUBS 0.009581f
C70 B.n39 VSUBS 0.009581f
C71 B.n40 VSUBS 0.009581f
C72 B.t8 VSUBS 0.040757f
C73 B.t7 VSUBS 0.054072f
C74 B.t6 VSUBS 0.326272f
C75 B.n41 VSUBS 0.095003f
C76 B.n42 VSUBS 0.075191f
C77 B.n43 VSUBS 0.009581f
C78 B.n44 VSUBS 0.009581f
C79 B.n45 VSUBS 0.009581f
C80 B.n46 VSUBS 0.009581f
C81 B.n47 VSUBS 0.02072f
C82 B.n48 VSUBS 0.009581f
C83 B.n49 VSUBS 0.009581f
C84 B.n50 VSUBS 0.009581f
C85 B.n51 VSUBS 0.009581f
C86 B.n52 VSUBS 0.009581f
C87 B.n53 VSUBS 0.009581f
C88 B.n54 VSUBS 0.009581f
C89 B.n55 VSUBS 0.009581f
C90 B.n56 VSUBS 0.009581f
C91 B.n57 VSUBS 0.009581f
C92 B.n58 VSUBS 0.009581f
C93 B.n59 VSUBS 0.009581f
C94 B.n60 VSUBS 0.009581f
C95 B.n61 VSUBS 0.009581f
C96 B.n62 VSUBS 0.009581f
C97 B.n63 VSUBS 0.009581f
C98 B.n64 VSUBS 0.009581f
C99 B.n65 VSUBS 0.009581f
C100 B.n66 VSUBS 0.009581f
C101 B.n67 VSUBS 0.009581f
C102 B.n68 VSUBS 0.009581f
C103 B.n69 VSUBS 0.009581f
C104 B.n70 VSUBS 0.009581f
C105 B.n71 VSUBS 0.009581f
C106 B.n72 VSUBS 0.009581f
C107 B.n73 VSUBS 0.009581f
C108 B.n74 VSUBS 0.009581f
C109 B.n75 VSUBS 0.009581f
C110 B.n76 VSUBS 0.009581f
C111 B.n77 VSUBS 0.009581f
C112 B.n78 VSUBS 0.009581f
C113 B.n79 VSUBS 0.009581f
C114 B.n80 VSUBS 0.009581f
C115 B.n81 VSUBS 0.009581f
C116 B.n82 VSUBS 0.009581f
C117 B.n83 VSUBS 0.009581f
C118 B.n84 VSUBS 0.009581f
C119 B.n85 VSUBS 0.009581f
C120 B.n86 VSUBS 0.009581f
C121 B.n87 VSUBS 0.009581f
C122 B.n88 VSUBS 0.009581f
C123 B.n89 VSUBS 0.009581f
C124 B.n90 VSUBS 0.009581f
C125 B.n91 VSUBS 0.009581f
C126 B.n92 VSUBS 0.009581f
C127 B.n93 VSUBS 0.009581f
C128 B.n94 VSUBS 0.009581f
C129 B.n95 VSUBS 0.009581f
C130 B.n96 VSUBS 0.009581f
C131 B.n97 VSUBS 0.009581f
C132 B.n98 VSUBS 0.021934f
C133 B.n99 VSUBS 0.009581f
C134 B.n100 VSUBS 0.009581f
C135 B.n101 VSUBS 0.009581f
C136 B.n102 VSUBS 0.009581f
C137 B.n103 VSUBS 0.006622f
C138 B.n104 VSUBS 0.009581f
C139 B.n105 VSUBS 0.009581f
C140 B.n106 VSUBS 0.009581f
C141 B.n107 VSUBS 0.009581f
C142 B.n108 VSUBS 0.009581f
C143 B.t1 VSUBS 0.040757f
C144 B.t2 VSUBS 0.054072f
C145 B.t0 VSUBS 0.326272f
C146 B.n109 VSUBS 0.095003f
C147 B.n110 VSUBS 0.075191f
C148 B.n111 VSUBS 0.009581f
C149 B.n112 VSUBS 0.009581f
C150 B.n113 VSUBS 0.009581f
C151 B.n114 VSUBS 0.009581f
C152 B.n115 VSUBS 0.021934f
C153 B.n116 VSUBS 0.009581f
C154 B.n117 VSUBS 0.009581f
C155 B.n118 VSUBS 0.009581f
C156 B.n119 VSUBS 0.009581f
C157 B.n120 VSUBS 0.009581f
C158 B.n121 VSUBS 0.009581f
C159 B.n122 VSUBS 0.009581f
C160 B.n123 VSUBS 0.009581f
C161 B.n124 VSUBS 0.009581f
C162 B.n125 VSUBS 0.009581f
C163 B.n126 VSUBS 0.009581f
C164 B.n127 VSUBS 0.009581f
C165 B.n128 VSUBS 0.009581f
C166 B.n129 VSUBS 0.009581f
C167 B.n130 VSUBS 0.009581f
C168 B.n131 VSUBS 0.009581f
C169 B.n132 VSUBS 0.009581f
C170 B.n133 VSUBS 0.009581f
C171 B.n134 VSUBS 0.009581f
C172 B.n135 VSUBS 0.009581f
C173 B.n136 VSUBS 0.009581f
C174 B.n137 VSUBS 0.009581f
C175 B.n138 VSUBS 0.009581f
C176 B.n139 VSUBS 0.009581f
C177 B.n140 VSUBS 0.009581f
C178 B.n141 VSUBS 0.009581f
C179 B.n142 VSUBS 0.009581f
C180 B.n143 VSUBS 0.009581f
C181 B.n144 VSUBS 0.009581f
C182 B.n145 VSUBS 0.009581f
C183 B.n146 VSUBS 0.009581f
C184 B.n147 VSUBS 0.009581f
C185 B.n148 VSUBS 0.009581f
C186 B.n149 VSUBS 0.009581f
C187 B.n150 VSUBS 0.009581f
C188 B.n151 VSUBS 0.009581f
C189 B.n152 VSUBS 0.009581f
C190 B.n153 VSUBS 0.009581f
C191 B.n154 VSUBS 0.009581f
C192 B.n155 VSUBS 0.009581f
C193 B.n156 VSUBS 0.009581f
C194 B.n157 VSUBS 0.009581f
C195 B.n158 VSUBS 0.009581f
C196 B.n159 VSUBS 0.009581f
C197 B.n160 VSUBS 0.009581f
C198 B.n161 VSUBS 0.009581f
C199 B.n162 VSUBS 0.009581f
C200 B.n163 VSUBS 0.009581f
C201 B.n164 VSUBS 0.009581f
C202 B.n165 VSUBS 0.009581f
C203 B.n166 VSUBS 0.009581f
C204 B.n167 VSUBS 0.009581f
C205 B.n168 VSUBS 0.009581f
C206 B.n169 VSUBS 0.009581f
C207 B.n170 VSUBS 0.009581f
C208 B.n171 VSUBS 0.009581f
C209 B.n172 VSUBS 0.009581f
C210 B.n173 VSUBS 0.009581f
C211 B.n174 VSUBS 0.009581f
C212 B.n175 VSUBS 0.009581f
C213 B.n176 VSUBS 0.009581f
C214 B.n177 VSUBS 0.009581f
C215 B.n178 VSUBS 0.009581f
C216 B.n179 VSUBS 0.009581f
C217 B.n180 VSUBS 0.009581f
C218 B.n181 VSUBS 0.009581f
C219 B.n182 VSUBS 0.009581f
C220 B.n183 VSUBS 0.009581f
C221 B.n184 VSUBS 0.009581f
C222 B.n185 VSUBS 0.009581f
C223 B.n186 VSUBS 0.009581f
C224 B.n187 VSUBS 0.009581f
C225 B.n188 VSUBS 0.009581f
C226 B.n189 VSUBS 0.009581f
C227 B.n190 VSUBS 0.009581f
C228 B.n191 VSUBS 0.009581f
C229 B.n192 VSUBS 0.009581f
C230 B.n193 VSUBS 0.009581f
C231 B.n194 VSUBS 0.009581f
C232 B.n195 VSUBS 0.009581f
C233 B.n196 VSUBS 0.009581f
C234 B.n197 VSUBS 0.009581f
C235 B.n198 VSUBS 0.009581f
C236 B.n199 VSUBS 0.009581f
C237 B.n200 VSUBS 0.009581f
C238 B.n201 VSUBS 0.009581f
C239 B.n202 VSUBS 0.009581f
C240 B.n203 VSUBS 0.009581f
C241 B.n204 VSUBS 0.009581f
C242 B.n205 VSUBS 0.009581f
C243 B.n206 VSUBS 0.009581f
C244 B.n207 VSUBS 0.009581f
C245 B.n208 VSUBS 0.009581f
C246 B.n209 VSUBS 0.009581f
C247 B.n210 VSUBS 0.009581f
C248 B.n211 VSUBS 0.009581f
C249 B.n212 VSUBS 0.020897f
C250 B.n213 VSUBS 0.020897f
C251 B.n214 VSUBS 0.021934f
C252 B.n215 VSUBS 0.009581f
C253 B.n216 VSUBS 0.009581f
C254 B.n217 VSUBS 0.009581f
C255 B.n218 VSUBS 0.009581f
C256 B.n219 VSUBS 0.009581f
C257 B.n220 VSUBS 0.009581f
C258 B.n221 VSUBS 0.009581f
C259 B.n222 VSUBS 0.009581f
C260 B.n223 VSUBS 0.009581f
C261 B.n224 VSUBS 0.009581f
C262 B.n225 VSUBS 0.009581f
C263 B.n226 VSUBS 0.009581f
C264 B.n227 VSUBS 0.009581f
C265 B.n228 VSUBS 0.009581f
C266 B.n229 VSUBS 0.006622f
C267 B.n230 VSUBS 0.022198f
C268 B.n231 VSUBS 0.007749f
C269 B.n232 VSUBS 0.009581f
C270 B.n233 VSUBS 0.009581f
C271 B.n234 VSUBS 0.009581f
C272 B.n235 VSUBS 0.009581f
C273 B.n236 VSUBS 0.009581f
C274 B.n237 VSUBS 0.009581f
C275 B.n238 VSUBS 0.009581f
C276 B.n239 VSUBS 0.009581f
C277 B.n240 VSUBS 0.009581f
C278 B.n241 VSUBS 0.009581f
C279 B.n242 VSUBS 0.009581f
C280 B.t4 VSUBS 0.040757f
C281 B.t5 VSUBS 0.054072f
C282 B.t3 VSUBS 0.326272f
C283 B.n243 VSUBS 0.095003f
C284 B.n244 VSUBS 0.075191f
C285 B.n245 VSUBS 0.022198f
C286 B.n246 VSUBS 0.007749f
C287 B.n247 VSUBS 0.009581f
C288 B.n248 VSUBS 0.009581f
C289 B.n249 VSUBS 0.009581f
C290 B.n250 VSUBS 0.009581f
C291 B.n251 VSUBS 0.009581f
C292 B.n252 VSUBS 0.009581f
C293 B.n253 VSUBS 0.009581f
C294 B.n254 VSUBS 0.009581f
C295 B.n255 VSUBS 0.009581f
C296 B.n256 VSUBS 0.009581f
C297 B.n257 VSUBS 0.009581f
C298 B.n258 VSUBS 0.009581f
C299 B.n259 VSUBS 0.009581f
C300 B.n260 VSUBS 0.009581f
C301 B.n261 VSUBS 0.009581f
C302 B.n262 VSUBS 0.009581f
C303 B.n263 VSUBS 0.021934f
C304 B.n264 VSUBS 0.020897f
C305 B.n265 VSUBS 0.020897f
C306 B.n266 VSUBS 0.009581f
C307 B.n267 VSUBS 0.009581f
C308 B.n268 VSUBS 0.009581f
C309 B.n269 VSUBS 0.009581f
C310 B.n270 VSUBS 0.009581f
C311 B.n271 VSUBS 0.009581f
C312 B.n272 VSUBS 0.009581f
C313 B.n273 VSUBS 0.009581f
C314 B.n274 VSUBS 0.009581f
C315 B.n275 VSUBS 0.009581f
C316 B.n276 VSUBS 0.009581f
C317 B.n277 VSUBS 0.009581f
C318 B.n278 VSUBS 0.009581f
C319 B.n279 VSUBS 0.009581f
C320 B.n280 VSUBS 0.009581f
C321 B.n281 VSUBS 0.009581f
C322 B.n282 VSUBS 0.009581f
C323 B.n283 VSUBS 0.009581f
C324 B.n284 VSUBS 0.009581f
C325 B.n285 VSUBS 0.009581f
C326 B.n286 VSUBS 0.009581f
C327 B.n287 VSUBS 0.009581f
C328 B.n288 VSUBS 0.009581f
C329 B.n289 VSUBS 0.009581f
C330 B.n290 VSUBS 0.009581f
C331 B.n291 VSUBS 0.009581f
C332 B.n292 VSUBS 0.009581f
C333 B.n293 VSUBS 0.009581f
C334 B.n294 VSUBS 0.009581f
C335 B.n295 VSUBS 0.009581f
C336 B.n296 VSUBS 0.009581f
C337 B.n297 VSUBS 0.009581f
C338 B.n298 VSUBS 0.009581f
C339 B.n299 VSUBS 0.009581f
C340 B.n300 VSUBS 0.009581f
C341 B.n301 VSUBS 0.009581f
C342 B.n302 VSUBS 0.009581f
C343 B.n303 VSUBS 0.009581f
C344 B.n304 VSUBS 0.009581f
C345 B.n305 VSUBS 0.009581f
C346 B.n306 VSUBS 0.009581f
C347 B.n307 VSUBS 0.009581f
C348 B.n308 VSUBS 0.009581f
C349 B.n309 VSUBS 0.009581f
C350 B.n310 VSUBS 0.009581f
C351 B.n311 VSUBS 0.009581f
C352 B.n312 VSUBS 0.009581f
C353 B.n313 VSUBS 0.009581f
C354 B.n314 VSUBS 0.009581f
C355 B.n315 VSUBS 0.009581f
C356 B.n316 VSUBS 0.009581f
C357 B.n317 VSUBS 0.009581f
C358 B.n318 VSUBS 0.009581f
C359 B.n319 VSUBS 0.009581f
C360 B.n320 VSUBS 0.009581f
C361 B.n321 VSUBS 0.009581f
C362 B.n322 VSUBS 0.009581f
C363 B.n323 VSUBS 0.009581f
C364 B.n324 VSUBS 0.009581f
C365 B.n325 VSUBS 0.009581f
C366 B.n326 VSUBS 0.009581f
C367 B.n327 VSUBS 0.009581f
C368 B.n328 VSUBS 0.009581f
C369 B.n329 VSUBS 0.009581f
C370 B.n330 VSUBS 0.009581f
C371 B.n331 VSUBS 0.009581f
C372 B.n332 VSUBS 0.009581f
C373 B.n333 VSUBS 0.009581f
C374 B.n334 VSUBS 0.009581f
C375 B.n335 VSUBS 0.009581f
C376 B.n336 VSUBS 0.009581f
C377 B.n337 VSUBS 0.009581f
C378 B.n338 VSUBS 0.009581f
C379 B.n339 VSUBS 0.009581f
C380 B.n340 VSUBS 0.009581f
C381 B.n341 VSUBS 0.009581f
C382 B.n342 VSUBS 0.009581f
C383 B.n343 VSUBS 0.009581f
C384 B.n344 VSUBS 0.009581f
C385 B.n345 VSUBS 0.009581f
C386 B.n346 VSUBS 0.009581f
C387 B.n347 VSUBS 0.009581f
C388 B.n348 VSUBS 0.009581f
C389 B.n349 VSUBS 0.009581f
C390 B.n350 VSUBS 0.009581f
C391 B.n351 VSUBS 0.009581f
C392 B.n352 VSUBS 0.009581f
C393 B.n353 VSUBS 0.009581f
C394 B.n354 VSUBS 0.009581f
C395 B.n355 VSUBS 0.009581f
C396 B.n356 VSUBS 0.009581f
C397 B.n357 VSUBS 0.009581f
C398 B.n358 VSUBS 0.009581f
C399 B.n359 VSUBS 0.009581f
C400 B.n360 VSUBS 0.009581f
C401 B.n361 VSUBS 0.009581f
C402 B.n362 VSUBS 0.009581f
C403 B.n363 VSUBS 0.009581f
C404 B.n364 VSUBS 0.009581f
C405 B.n365 VSUBS 0.009581f
C406 B.n366 VSUBS 0.009581f
C407 B.n367 VSUBS 0.009581f
C408 B.n368 VSUBS 0.009581f
C409 B.n369 VSUBS 0.009581f
C410 B.n370 VSUBS 0.009581f
C411 B.n371 VSUBS 0.009581f
C412 B.n372 VSUBS 0.009581f
C413 B.n373 VSUBS 0.009581f
C414 B.n374 VSUBS 0.009581f
C415 B.n375 VSUBS 0.009581f
C416 B.n376 VSUBS 0.009581f
C417 B.n377 VSUBS 0.009581f
C418 B.n378 VSUBS 0.009581f
C419 B.n379 VSUBS 0.009581f
C420 B.n380 VSUBS 0.009581f
C421 B.n381 VSUBS 0.009581f
C422 B.n382 VSUBS 0.009581f
C423 B.n383 VSUBS 0.009581f
C424 B.n384 VSUBS 0.009581f
C425 B.n385 VSUBS 0.009581f
C426 B.n386 VSUBS 0.009581f
C427 B.n387 VSUBS 0.009581f
C428 B.n388 VSUBS 0.009581f
C429 B.n389 VSUBS 0.009581f
C430 B.n390 VSUBS 0.009581f
C431 B.n391 VSUBS 0.009581f
C432 B.n392 VSUBS 0.009581f
C433 B.n393 VSUBS 0.009581f
C434 B.n394 VSUBS 0.009581f
C435 B.n395 VSUBS 0.009581f
C436 B.n396 VSUBS 0.009581f
C437 B.n397 VSUBS 0.009581f
C438 B.n398 VSUBS 0.009581f
C439 B.n399 VSUBS 0.009581f
C440 B.n400 VSUBS 0.009581f
C441 B.n401 VSUBS 0.009581f
C442 B.n402 VSUBS 0.009581f
C443 B.n403 VSUBS 0.009581f
C444 B.n404 VSUBS 0.009581f
C445 B.n405 VSUBS 0.009581f
C446 B.n406 VSUBS 0.009581f
C447 B.n407 VSUBS 0.009581f
C448 B.n408 VSUBS 0.009581f
C449 B.n409 VSUBS 0.009581f
C450 B.n410 VSUBS 0.009581f
C451 B.n411 VSUBS 0.009581f
C452 B.n412 VSUBS 0.009581f
C453 B.n413 VSUBS 0.009581f
C454 B.n414 VSUBS 0.022112f
C455 B.n415 VSUBS 0.020897f
C456 B.n416 VSUBS 0.021934f
C457 B.n417 VSUBS 0.009581f
C458 B.n418 VSUBS 0.009581f
C459 B.n419 VSUBS 0.009581f
C460 B.n420 VSUBS 0.009581f
C461 B.n421 VSUBS 0.009581f
C462 B.n422 VSUBS 0.009581f
C463 B.n423 VSUBS 0.009581f
C464 B.n424 VSUBS 0.009581f
C465 B.n425 VSUBS 0.009581f
C466 B.n426 VSUBS 0.009581f
C467 B.n427 VSUBS 0.009581f
C468 B.n428 VSUBS 0.009581f
C469 B.n429 VSUBS 0.009581f
C470 B.n430 VSUBS 0.009581f
C471 B.n431 VSUBS 0.006622f
C472 B.n432 VSUBS 0.022198f
C473 B.n433 VSUBS 0.007749f
C474 B.n434 VSUBS 0.009581f
C475 B.n435 VSUBS 0.009581f
C476 B.n436 VSUBS 0.009581f
C477 B.n437 VSUBS 0.009581f
C478 B.n438 VSUBS 0.009581f
C479 B.n439 VSUBS 0.009581f
C480 B.n440 VSUBS 0.009581f
C481 B.n441 VSUBS 0.009581f
C482 B.n442 VSUBS 0.009581f
C483 B.n443 VSUBS 0.009581f
C484 B.n444 VSUBS 0.009581f
C485 B.n445 VSUBS 0.007749f
C486 B.n446 VSUBS 0.009581f
C487 B.n447 VSUBS 0.009581f
C488 B.n448 VSUBS 0.009581f
C489 B.n449 VSUBS 0.009581f
C490 B.n450 VSUBS 0.009581f
C491 B.n451 VSUBS 0.009581f
C492 B.n452 VSUBS 0.009581f
C493 B.n453 VSUBS 0.009581f
C494 B.n454 VSUBS 0.009581f
C495 B.n455 VSUBS 0.009581f
C496 B.n456 VSUBS 0.009581f
C497 B.n457 VSUBS 0.009581f
C498 B.n458 VSUBS 0.009581f
C499 B.n459 VSUBS 0.009581f
C500 B.n460 VSUBS 0.009581f
C501 B.n461 VSUBS 0.009581f
C502 B.n462 VSUBS 0.021934f
C503 B.n463 VSUBS 0.020897f
C504 B.n464 VSUBS 0.020897f
C505 B.n465 VSUBS 0.009581f
C506 B.n466 VSUBS 0.009581f
C507 B.n467 VSUBS 0.009581f
C508 B.n468 VSUBS 0.009581f
C509 B.n469 VSUBS 0.009581f
C510 B.n470 VSUBS 0.009581f
C511 B.n471 VSUBS 0.009581f
C512 B.n472 VSUBS 0.009581f
C513 B.n473 VSUBS 0.009581f
C514 B.n474 VSUBS 0.009581f
C515 B.n475 VSUBS 0.009581f
C516 B.n476 VSUBS 0.009581f
C517 B.n477 VSUBS 0.009581f
C518 B.n478 VSUBS 0.009581f
C519 B.n479 VSUBS 0.009581f
C520 B.n480 VSUBS 0.009581f
C521 B.n481 VSUBS 0.009581f
C522 B.n482 VSUBS 0.009581f
C523 B.n483 VSUBS 0.009581f
C524 B.n484 VSUBS 0.009581f
C525 B.n485 VSUBS 0.009581f
C526 B.n486 VSUBS 0.009581f
C527 B.n487 VSUBS 0.009581f
C528 B.n488 VSUBS 0.009581f
C529 B.n489 VSUBS 0.009581f
C530 B.n490 VSUBS 0.009581f
C531 B.n491 VSUBS 0.009581f
C532 B.n492 VSUBS 0.009581f
C533 B.n493 VSUBS 0.009581f
C534 B.n494 VSUBS 0.009581f
C535 B.n495 VSUBS 0.009581f
C536 B.n496 VSUBS 0.009581f
C537 B.n497 VSUBS 0.009581f
C538 B.n498 VSUBS 0.009581f
C539 B.n499 VSUBS 0.009581f
C540 B.n500 VSUBS 0.009581f
C541 B.n501 VSUBS 0.009581f
C542 B.n502 VSUBS 0.009581f
C543 B.n503 VSUBS 0.009581f
C544 B.n504 VSUBS 0.009581f
C545 B.n505 VSUBS 0.009581f
C546 B.n506 VSUBS 0.009581f
C547 B.n507 VSUBS 0.009581f
C548 B.n508 VSUBS 0.009581f
C549 B.n509 VSUBS 0.009581f
C550 B.n510 VSUBS 0.009581f
C551 B.n511 VSUBS 0.009581f
C552 B.n512 VSUBS 0.009581f
C553 B.n513 VSUBS 0.009581f
C554 B.n514 VSUBS 0.009581f
C555 B.n515 VSUBS 0.009581f
C556 B.n516 VSUBS 0.009581f
C557 B.n517 VSUBS 0.009581f
C558 B.n518 VSUBS 0.009581f
C559 B.n519 VSUBS 0.009581f
C560 B.n520 VSUBS 0.009581f
C561 B.n521 VSUBS 0.009581f
C562 B.n522 VSUBS 0.009581f
C563 B.n523 VSUBS 0.009581f
C564 B.n524 VSUBS 0.009581f
C565 B.n525 VSUBS 0.009581f
C566 B.n526 VSUBS 0.009581f
C567 B.n527 VSUBS 0.009581f
C568 B.n528 VSUBS 0.009581f
C569 B.n529 VSUBS 0.009581f
C570 B.n530 VSUBS 0.009581f
C571 B.n531 VSUBS 0.009581f
C572 B.n532 VSUBS 0.009581f
C573 B.n533 VSUBS 0.009581f
C574 B.n534 VSUBS 0.009581f
C575 B.n535 VSUBS 0.009581f
C576 B.n536 VSUBS 0.009581f
C577 B.n537 VSUBS 0.009581f
C578 B.n538 VSUBS 0.009581f
C579 B.n539 VSUBS 0.021694f
C580 VDD1.t5 VSUBS 0.127535f
C581 VDD1.t0 VSUBS 0.127356f
C582 VDD1.t1 VSUBS 0.020496f
C583 VDD1.t2 VSUBS 0.020496f
C584 VDD1.n0 VSUBS 0.079269f
C585 VDD1.n1 VSUBS 1.89182f
C586 VDD1.t3 VSUBS 0.020496f
C587 VDD1.t4 VSUBS 0.020496f
C588 VDD1.n2 VSUBS 0.078185f
C589 VDD1.n3 VSUBS 1.53067f
C590 VP.t3 VSUBS 0.562812f
C591 VP.n0 VSUBS 0.504284f
C592 VP.n1 VSUBS 0.05487f
C593 VP.n2 VSUBS 0.044801f
C594 VP.n3 VSUBS 0.05487f
C595 VP.t4 VSUBS 0.562812f
C596 VP.n4 VSUBS 0.293108f
C597 VP.n5 VSUBS 0.05487f
C598 VP.n6 VSUBS 0.044801f
C599 VP.n7 VSUBS 0.05487f
C600 VP.t5 VSUBS 0.562812f
C601 VP.n8 VSUBS 0.504284f
C602 VP.t1 VSUBS 0.562812f
C603 VP.n9 VSUBS 0.504284f
C604 VP.n10 VSUBS 0.05487f
C605 VP.n11 VSUBS 0.044801f
C606 VP.n12 VSUBS 0.05487f
C607 VP.t2 VSUBS 0.562812f
C608 VP.n13 VSUBS 0.474163f
C609 VP.t0 VSUBS 1.0726f
C610 VP.n14 VSUBS 0.512113f
C611 VP.n15 VSUBS 0.639444f
C612 VP.n16 VSUBS 0.07702f
C613 VP.n17 VSUBS 0.102264f
C614 VP.n18 VSUBS 0.110199f
C615 VP.n19 VSUBS 0.05487f
C616 VP.n20 VSUBS 0.05487f
C617 VP.n21 VSUBS 0.05487f
C618 VP.n22 VSUBS 0.107473f
C619 VP.n23 VSUBS 0.102264f
C620 VP.n24 VSUBS 0.082068f
C621 VP.n25 VSUBS 0.088559f
C622 VP.n26 VSUBS 2.50996f
C623 VP.n27 VSUBS 2.55559f
C624 VP.n28 VSUBS 0.088559f
C625 VP.n29 VSUBS 0.082068f
C626 VP.n30 VSUBS 0.102264f
C627 VP.n31 VSUBS 0.107473f
C628 VP.n32 VSUBS 0.05487f
C629 VP.n33 VSUBS 0.05487f
C630 VP.n34 VSUBS 0.05487f
C631 VP.n35 VSUBS 0.110199f
C632 VP.n36 VSUBS 0.102264f
C633 VP.n37 VSUBS 0.07702f
C634 VP.n38 VSUBS 0.05487f
C635 VP.n39 VSUBS 0.05487f
C636 VP.n40 VSUBS 0.07702f
C637 VP.n41 VSUBS 0.102264f
C638 VP.n42 VSUBS 0.110199f
C639 VP.n43 VSUBS 0.05487f
C640 VP.n44 VSUBS 0.05487f
C641 VP.n45 VSUBS 0.05487f
C642 VP.n46 VSUBS 0.107473f
C643 VP.n47 VSUBS 0.102264f
C644 VP.n48 VSUBS 0.082068f
C645 VP.n49 VSUBS 0.088559f
C646 VP.n50 VSUBS 0.130972f
C647 VTAIL.t9 VSUBS 0.044253f
C648 VTAIL.t8 VSUBS 0.044253f
C649 VTAIL.n0 VSUBS 0.144404f
C650 VTAIL.n1 VSUBS 0.668385f
C651 VTAIL.t2 VSUBS 0.246003f
C652 VTAIL.n2 VSUBS 0.962078f
C653 VTAIL.t1 VSUBS 0.044253f
C654 VTAIL.t0 VSUBS 0.044253f
C655 VTAIL.n3 VSUBS 0.144404f
C656 VTAIL.n4 VSUBS 2.12184f
C657 VTAIL.t6 VSUBS 0.044253f
C658 VTAIL.t11 VSUBS 0.044253f
C659 VTAIL.n5 VSUBS 0.144404f
C660 VTAIL.n6 VSUBS 2.12184f
C661 VTAIL.t10 VSUBS 0.246004f
C662 VTAIL.n7 VSUBS 0.962077f
C663 VTAIL.t4 VSUBS 0.044253f
C664 VTAIL.t3 VSUBS 0.044253f
C665 VTAIL.n8 VSUBS 0.144404f
C666 VTAIL.n9 VSUBS 0.942987f
C667 VTAIL.t5 VSUBS 0.246003f
C668 VTAIL.n10 VSUBS 1.76527f
C669 VTAIL.t7 VSUBS 0.246003f
C670 VTAIL.n11 VSUBS 1.66421f
C671 VDD2.t4 VSUBS 0.129271f
C672 VDD2.t5 VSUBS 0.020804f
C673 VDD2.t3 VSUBS 0.020804f
C674 VDD2.n0 VSUBS 0.080461f
C675 VDD2.n1 VSUBS 1.82865f
C676 VDD2.t2 VSUBS 0.126742f
C677 VDD2.n2 VSUBS 1.50692f
C678 VDD2.t0 VSUBS 0.020804f
C679 VDD2.t1 VSUBS 0.020804f
C680 VDD2.n3 VSUBS 0.080455f
C681 VN.t4 VSUBS 0.538657f
C682 VN.n0 VSUBS 0.482641f
C683 VN.n1 VSUBS 0.052515f
C684 VN.n2 VSUBS 0.042879f
C685 VN.n3 VSUBS 0.052515f
C686 VN.t3 VSUBS 0.538657f
C687 VN.n4 VSUBS 0.453813f
C688 VN.t2 VSUBS 1.02657f
C689 VN.n5 VSUBS 0.490133f
C690 VN.n6 VSUBS 0.611999f
C691 VN.n7 VSUBS 0.073714f
C692 VN.n8 VSUBS 0.097875f
C693 VN.n9 VSUBS 0.10547f
C694 VN.n10 VSUBS 0.052515f
C695 VN.n11 VSUBS 0.052515f
C696 VN.n12 VSUBS 0.052515f
C697 VN.n13 VSUBS 0.102861f
C698 VN.n14 VSUBS 0.097875f
C699 VN.n15 VSUBS 0.078546f
C700 VN.n16 VSUBS 0.084758f
C701 VN.n17 VSUBS 0.125351f
C702 VN.t5 VSUBS 0.538657f
C703 VN.n18 VSUBS 0.482641f
C704 VN.n19 VSUBS 0.052515f
C705 VN.n20 VSUBS 0.042879f
C706 VN.n21 VSUBS 0.052515f
C707 VN.t0 VSUBS 0.538657f
C708 VN.n22 VSUBS 0.453813f
C709 VN.t1 VSUBS 1.02657f
C710 VN.n23 VSUBS 0.490133f
C711 VN.n24 VSUBS 0.611999f
C712 VN.n25 VSUBS 0.073714f
C713 VN.n26 VSUBS 0.097875f
C714 VN.n27 VSUBS 0.10547f
C715 VN.n28 VSUBS 0.052515f
C716 VN.n29 VSUBS 0.052515f
C717 VN.n30 VSUBS 0.052515f
C718 VN.n31 VSUBS 0.102861f
C719 VN.n32 VSUBS 0.097875f
C720 VN.n33 VSUBS 0.078546f
C721 VN.n34 VSUBS 0.084758f
C722 VN.n35 VSUBS 2.42488f
.ends

