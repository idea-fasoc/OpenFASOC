* NGSPICE file created from diff_pair_sample_0290.ext - technology: sky130A

.subckt diff_pair_sample_0290 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t5 VP.t0 VTAIL.t9 w_n3658_n4352# sky130_fd_pr__pfet_01v8 ad=2.7918 pd=17.25 as=6.5988 ps=34.62 w=16.92 l=3.03
X1 VDD2.t5 VN.t0 VTAIL.t4 w_n3658_n4352# sky130_fd_pr__pfet_01v8 ad=2.7918 pd=17.25 as=6.5988 ps=34.62 w=16.92 l=3.03
X2 VDD2.t4 VN.t1 VTAIL.t0 w_n3658_n4352# sky130_fd_pr__pfet_01v8 ad=6.5988 pd=34.62 as=2.7918 ps=17.25 w=16.92 l=3.03
X3 VTAIL.t3 VN.t2 VDD2.t3 w_n3658_n4352# sky130_fd_pr__pfet_01v8 ad=2.7918 pd=17.25 as=2.7918 ps=17.25 w=16.92 l=3.03
X4 VDD1.t4 VP.t1 VTAIL.t8 w_n3658_n4352# sky130_fd_pr__pfet_01v8 ad=6.5988 pd=34.62 as=2.7918 ps=17.25 w=16.92 l=3.03
X5 VTAIL.t7 VP.t2 VDD1.t3 w_n3658_n4352# sky130_fd_pr__pfet_01v8 ad=2.7918 pd=17.25 as=2.7918 ps=17.25 w=16.92 l=3.03
X6 VDD2.t2 VN.t3 VTAIL.t2 w_n3658_n4352# sky130_fd_pr__pfet_01v8 ad=2.7918 pd=17.25 as=6.5988 ps=34.62 w=16.92 l=3.03
X7 VTAIL.t1 VN.t4 VDD2.t1 w_n3658_n4352# sky130_fd_pr__pfet_01v8 ad=2.7918 pd=17.25 as=2.7918 ps=17.25 w=16.92 l=3.03
X8 VTAIL.t11 VP.t3 VDD1.t2 w_n3658_n4352# sky130_fd_pr__pfet_01v8 ad=2.7918 pd=17.25 as=2.7918 ps=17.25 w=16.92 l=3.03
X9 B.t11 B.t9 B.t10 w_n3658_n4352# sky130_fd_pr__pfet_01v8 ad=6.5988 pd=34.62 as=0 ps=0 w=16.92 l=3.03
X10 B.t8 B.t6 B.t7 w_n3658_n4352# sky130_fd_pr__pfet_01v8 ad=6.5988 pd=34.62 as=0 ps=0 w=16.92 l=3.03
X11 VDD1.t1 VP.t4 VTAIL.t10 w_n3658_n4352# sky130_fd_pr__pfet_01v8 ad=6.5988 pd=34.62 as=2.7918 ps=17.25 w=16.92 l=3.03
X12 B.t5 B.t3 B.t4 w_n3658_n4352# sky130_fd_pr__pfet_01v8 ad=6.5988 pd=34.62 as=0 ps=0 w=16.92 l=3.03
X13 B.t2 B.t0 B.t1 w_n3658_n4352# sky130_fd_pr__pfet_01v8 ad=6.5988 pd=34.62 as=0 ps=0 w=16.92 l=3.03
X14 VDD2.t0 VN.t5 VTAIL.t5 w_n3658_n4352# sky130_fd_pr__pfet_01v8 ad=6.5988 pd=34.62 as=2.7918 ps=17.25 w=16.92 l=3.03
X15 VDD1.t0 VP.t5 VTAIL.t6 w_n3658_n4352# sky130_fd_pr__pfet_01v8 ad=2.7918 pd=17.25 as=6.5988 ps=34.62 w=16.92 l=3.03
R0 VP.n11 VP.t4 167.808
R1 VP.n13 VP.n10 161.3
R2 VP.n15 VP.n14 161.3
R3 VP.n16 VP.n9 161.3
R4 VP.n18 VP.n17 161.3
R5 VP.n19 VP.n8 161.3
R6 VP.n21 VP.n20 161.3
R7 VP.n44 VP.n43 161.3
R8 VP.n42 VP.n1 161.3
R9 VP.n41 VP.n40 161.3
R10 VP.n39 VP.n2 161.3
R11 VP.n38 VP.n37 161.3
R12 VP.n36 VP.n3 161.3
R13 VP.n35 VP.n34 161.3
R14 VP.n33 VP.n4 161.3
R15 VP.n32 VP.n31 161.3
R16 VP.n30 VP.n5 161.3
R17 VP.n29 VP.n28 161.3
R18 VP.n27 VP.n6 161.3
R19 VP.n26 VP.n25 161.3
R20 VP.n35 VP.t2 134.578
R21 VP.n24 VP.t1 134.578
R22 VP.n0 VP.t5 134.578
R23 VP.n12 VP.t3 134.578
R24 VP.n7 VP.t0 134.578
R25 VP.n24 VP.n23 72.3637
R26 VP.n45 VP.n0 72.3637
R27 VP.n22 VP.n7 72.3637
R28 VP.n30 VP.n29 56.4773
R29 VP.n41 VP.n2 56.4773
R30 VP.n18 VP.n9 56.4773
R31 VP.n23 VP.n22 54.1809
R32 VP.n12 VP.n11 49.1756
R33 VP.n25 VP.n6 24.3439
R34 VP.n29 VP.n6 24.3439
R35 VP.n31 VP.n30 24.3439
R36 VP.n31 VP.n4 24.3439
R37 VP.n35 VP.n4 24.3439
R38 VP.n36 VP.n35 24.3439
R39 VP.n37 VP.n36 24.3439
R40 VP.n37 VP.n2 24.3439
R41 VP.n42 VP.n41 24.3439
R42 VP.n43 VP.n42 24.3439
R43 VP.n19 VP.n18 24.3439
R44 VP.n20 VP.n19 24.3439
R45 VP.n13 VP.n12 24.3439
R46 VP.n14 VP.n13 24.3439
R47 VP.n14 VP.n9 24.3439
R48 VP.n25 VP.n24 17.5278
R49 VP.n43 VP.n0 17.5278
R50 VP.n20 VP.n7 17.5278
R51 VP.n11 VP.n10 4.04421
R52 VP.n22 VP.n21 0.355081
R53 VP.n26 VP.n23 0.355081
R54 VP.n45 VP.n44 0.355081
R55 VP VP.n45 0.26685
R56 VP.n15 VP.n10 0.189894
R57 VP.n16 VP.n15 0.189894
R58 VP.n17 VP.n16 0.189894
R59 VP.n17 VP.n8 0.189894
R60 VP.n21 VP.n8 0.189894
R61 VP.n27 VP.n26 0.189894
R62 VP.n28 VP.n27 0.189894
R63 VP.n28 VP.n5 0.189894
R64 VP.n32 VP.n5 0.189894
R65 VP.n33 VP.n32 0.189894
R66 VP.n34 VP.n33 0.189894
R67 VP.n34 VP.n3 0.189894
R68 VP.n38 VP.n3 0.189894
R69 VP.n39 VP.n38 0.189894
R70 VP.n40 VP.n39 0.189894
R71 VP.n40 VP.n1 0.189894
R72 VP.n44 VP.n1 0.189894
R73 VTAIL.n378 VTAIL.n290 756.745
R74 VTAIL.n90 VTAIL.n2 756.745
R75 VTAIL.n284 VTAIL.n196 756.745
R76 VTAIL.n188 VTAIL.n100 756.745
R77 VTAIL.n321 VTAIL.n320 585
R78 VTAIL.n318 VTAIL.n317 585
R79 VTAIL.n327 VTAIL.n326 585
R80 VTAIL.n329 VTAIL.n328 585
R81 VTAIL.n314 VTAIL.n313 585
R82 VTAIL.n335 VTAIL.n334 585
R83 VTAIL.n337 VTAIL.n336 585
R84 VTAIL.n310 VTAIL.n309 585
R85 VTAIL.n343 VTAIL.n342 585
R86 VTAIL.n345 VTAIL.n344 585
R87 VTAIL.n306 VTAIL.n305 585
R88 VTAIL.n351 VTAIL.n350 585
R89 VTAIL.n353 VTAIL.n352 585
R90 VTAIL.n302 VTAIL.n301 585
R91 VTAIL.n359 VTAIL.n358 585
R92 VTAIL.n362 VTAIL.n361 585
R93 VTAIL.n360 VTAIL.n298 585
R94 VTAIL.n367 VTAIL.n297 585
R95 VTAIL.n369 VTAIL.n368 585
R96 VTAIL.n371 VTAIL.n370 585
R97 VTAIL.n294 VTAIL.n293 585
R98 VTAIL.n377 VTAIL.n376 585
R99 VTAIL.n379 VTAIL.n378 585
R100 VTAIL.n33 VTAIL.n32 585
R101 VTAIL.n30 VTAIL.n29 585
R102 VTAIL.n39 VTAIL.n38 585
R103 VTAIL.n41 VTAIL.n40 585
R104 VTAIL.n26 VTAIL.n25 585
R105 VTAIL.n47 VTAIL.n46 585
R106 VTAIL.n49 VTAIL.n48 585
R107 VTAIL.n22 VTAIL.n21 585
R108 VTAIL.n55 VTAIL.n54 585
R109 VTAIL.n57 VTAIL.n56 585
R110 VTAIL.n18 VTAIL.n17 585
R111 VTAIL.n63 VTAIL.n62 585
R112 VTAIL.n65 VTAIL.n64 585
R113 VTAIL.n14 VTAIL.n13 585
R114 VTAIL.n71 VTAIL.n70 585
R115 VTAIL.n74 VTAIL.n73 585
R116 VTAIL.n72 VTAIL.n10 585
R117 VTAIL.n79 VTAIL.n9 585
R118 VTAIL.n81 VTAIL.n80 585
R119 VTAIL.n83 VTAIL.n82 585
R120 VTAIL.n6 VTAIL.n5 585
R121 VTAIL.n89 VTAIL.n88 585
R122 VTAIL.n91 VTAIL.n90 585
R123 VTAIL.n285 VTAIL.n284 585
R124 VTAIL.n283 VTAIL.n282 585
R125 VTAIL.n200 VTAIL.n199 585
R126 VTAIL.n277 VTAIL.n276 585
R127 VTAIL.n275 VTAIL.n274 585
R128 VTAIL.n273 VTAIL.n203 585
R129 VTAIL.n207 VTAIL.n204 585
R130 VTAIL.n268 VTAIL.n267 585
R131 VTAIL.n266 VTAIL.n265 585
R132 VTAIL.n209 VTAIL.n208 585
R133 VTAIL.n260 VTAIL.n259 585
R134 VTAIL.n258 VTAIL.n257 585
R135 VTAIL.n213 VTAIL.n212 585
R136 VTAIL.n252 VTAIL.n251 585
R137 VTAIL.n250 VTAIL.n249 585
R138 VTAIL.n217 VTAIL.n216 585
R139 VTAIL.n244 VTAIL.n243 585
R140 VTAIL.n242 VTAIL.n241 585
R141 VTAIL.n221 VTAIL.n220 585
R142 VTAIL.n236 VTAIL.n235 585
R143 VTAIL.n234 VTAIL.n233 585
R144 VTAIL.n225 VTAIL.n224 585
R145 VTAIL.n228 VTAIL.n227 585
R146 VTAIL.n189 VTAIL.n188 585
R147 VTAIL.n187 VTAIL.n186 585
R148 VTAIL.n104 VTAIL.n103 585
R149 VTAIL.n181 VTAIL.n180 585
R150 VTAIL.n179 VTAIL.n178 585
R151 VTAIL.n177 VTAIL.n107 585
R152 VTAIL.n111 VTAIL.n108 585
R153 VTAIL.n172 VTAIL.n171 585
R154 VTAIL.n170 VTAIL.n169 585
R155 VTAIL.n113 VTAIL.n112 585
R156 VTAIL.n164 VTAIL.n163 585
R157 VTAIL.n162 VTAIL.n161 585
R158 VTAIL.n117 VTAIL.n116 585
R159 VTAIL.n156 VTAIL.n155 585
R160 VTAIL.n154 VTAIL.n153 585
R161 VTAIL.n121 VTAIL.n120 585
R162 VTAIL.n148 VTAIL.n147 585
R163 VTAIL.n146 VTAIL.n145 585
R164 VTAIL.n125 VTAIL.n124 585
R165 VTAIL.n140 VTAIL.n139 585
R166 VTAIL.n138 VTAIL.n137 585
R167 VTAIL.n129 VTAIL.n128 585
R168 VTAIL.n132 VTAIL.n131 585
R169 VTAIL.t9 VTAIL.n226 327.466
R170 VTAIL.t2 VTAIL.n130 327.466
R171 VTAIL.t4 VTAIL.n319 327.466
R172 VTAIL.t6 VTAIL.n31 327.466
R173 VTAIL.n320 VTAIL.n317 171.744
R174 VTAIL.n327 VTAIL.n317 171.744
R175 VTAIL.n328 VTAIL.n327 171.744
R176 VTAIL.n328 VTAIL.n313 171.744
R177 VTAIL.n335 VTAIL.n313 171.744
R178 VTAIL.n336 VTAIL.n335 171.744
R179 VTAIL.n336 VTAIL.n309 171.744
R180 VTAIL.n343 VTAIL.n309 171.744
R181 VTAIL.n344 VTAIL.n343 171.744
R182 VTAIL.n344 VTAIL.n305 171.744
R183 VTAIL.n351 VTAIL.n305 171.744
R184 VTAIL.n352 VTAIL.n351 171.744
R185 VTAIL.n352 VTAIL.n301 171.744
R186 VTAIL.n359 VTAIL.n301 171.744
R187 VTAIL.n361 VTAIL.n359 171.744
R188 VTAIL.n361 VTAIL.n360 171.744
R189 VTAIL.n360 VTAIL.n297 171.744
R190 VTAIL.n369 VTAIL.n297 171.744
R191 VTAIL.n370 VTAIL.n369 171.744
R192 VTAIL.n370 VTAIL.n293 171.744
R193 VTAIL.n377 VTAIL.n293 171.744
R194 VTAIL.n378 VTAIL.n377 171.744
R195 VTAIL.n32 VTAIL.n29 171.744
R196 VTAIL.n39 VTAIL.n29 171.744
R197 VTAIL.n40 VTAIL.n39 171.744
R198 VTAIL.n40 VTAIL.n25 171.744
R199 VTAIL.n47 VTAIL.n25 171.744
R200 VTAIL.n48 VTAIL.n47 171.744
R201 VTAIL.n48 VTAIL.n21 171.744
R202 VTAIL.n55 VTAIL.n21 171.744
R203 VTAIL.n56 VTAIL.n55 171.744
R204 VTAIL.n56 VTAIL.n17 171.744
R205 VTAIL.n63 VTAIL.n17 171.744
R206 VTAIL.n64 VTAIL.n63 171.744
R207 VTAIL.n64 VTAIL.n13 171.744
R208 VTAIL.n71 VTAIL.n13 171.744
R209 VTAIL.n73 VTAIL.n71 171.744
R210 VTAIL.n73 VTAIL.n72 171.744
R211 VTAIL.n72 VTAIL.n9 171.744
R212 VTAIL.n81 VTAIL.n9 171.744
R213 VTAIL.n82 VTAIL.n81 171.744
R214 VTAIL.n82 VTAIL.n5 171.744
R215 VTAIL.n89 VTAIL.n5 171.744
R216 VTAIL.n90 VTAIL.n89 171.744
R217 VTAIL.n284 VTAIL.n283 171.744
R218 VTAIL.n283 VTAIL.n199 171.744
R219 VTAIL.n276 VTAIL.n199 171.744
R220 VTAIL.n276 VTAIL.n275 171.744
R221 VTAIL.n275 VTAIL.n203 171.744
R222 VTAIL.n207 VTAIL.n203 171.744
R223 VTAIL.n267 VTAIL.n207 171.744
R224 VTAIL.n267 VTAIL.n266 171.744
R225 VTAIL.n266 VTAIL.n208 171.744
R226 VTAIL.n259 VTAIL.n208 171.744
R227 VTAIL.n259 VTAIL.n258 171.744
R228 VTAIL.n258 VTAIL.n212 171.744
R229 VTAIL.n251 VTAIL.n212 171.744
R230 VTAIL.n251 VTAIL.n250 171.744
R231 VTAIL.n250 VTAIL.n216 171.744
R232 VTAIL.n243 VTAIL.n216 171.744
R233 VTAIL.n243 VTAIL.n242 171.744
R234 VTAIL.n242 VTAIL.n220 171.744
R235 VTAIL.n235 VTAIL.n220 171.744
R236 VTAIL.n235 VTAIL.n234 171.744
R237 VTAIL.n234 VTAIL.n224 171.744
R238 VTAIL.n227 VTAIL.n224 171.744
R239 VTAIL.n188 VTAIL.n187 171.744
R240 VTAIL.n187 VTAIL.n103 171.744
R241 VTAIL.n180 VTAIL.n103 171.744
R242 VTAIL.n180 VTAIL.n179 171.744
R243 VTAIL.n179 VTAIL.n107 171.744
R244 VTAIL.n111 VTAIL.n107 171.744
R245 VTAIL.n171 VTAIL.n111 171.744
R246 VTAIL.n171 VTAIL.n170 171.744
R247 VTAIL.n170 VTAIL.n112 171.744
R248 VTAIL.n163 VTAIL.n112 171.744
R249 VTAIL.n163 VTAIL.n162 171.744
R250 VTAIL.n162 VTAIL.n116 171.744
R251 VTAIL.n155 VTAIL.n116 171.744
R252 VTAIL.n155 VTAIL.n154 171.744
R253 VTAIL.n154 VTAIL.n120 171.744
R254 VTAIL.n147 VTAIL.n120 171.744
R255 VTAIL.n147 VTAIL.n146 171.744
R256 VTAIL.n146 VTAIL.n124 171.744
R257 VTAIL.n139 VTAIL.n124 171.744
R258 VTAIL.n139 VTAIL.n138 171.744
R259 VTAIL.n138 VTAIL.n128 171.744
R260 VTAIL.n131 VTAIL.n128 171.744
R261 VTAIL.n320 VTAIL.t4 85.8723
R262 VTAIL.n32 VTAIL.t6 85.8723
R263 VTAIL.n227 VTAIL.t9 85.8723
R264 VTAIL.n131 VTAIL.t2 85.8723
R265 VTAIL.n195 VTAIL.n194 55.0405
R266 VTAIL.n99 VTAIL.n98 55.0405
R267 VTAIL.n1 VTAIL.n0 55.0403
R268 VTAIL.n97 VTAIL.n96 55.0403
R269 VTAIL.n383 VTAIL.n382 34.5126
R270 VTAIL.n95 VTAIL.n94 34.5126
R271 VTAIL.n289 VTAIL.n288 34.5126
R272 VTAIL.n193 VTAIL.n192 34.5126
R273 VTAIL.n99 VTAIL.n97 32.7462
R274 VTAIL.n383 VTAIL.n289 29.8496
R275 VTAIL.n321 VTAIL.n319 16.3895
R276 VTAIL.n33 VTAIL.n31 16.3895
R277 VTAIL.n228 VTAIL.n226 16.3895
R278 VTAIL.n132 VTAIL.n130 16.3895
R279 VTAIL.n368 VTAIL.n367 13.1884
R280 VTAIL.n80 VTAIL.n79 13.1884
R281 VTAIL.n274 VTAIL.n273 13.1884
R282 VTAIL.n178 VTAIL.n177 13.1884
R283 VTAIL.n322 VTAIL.n318 12.8005
R284 VTAIL.n366 VTAIL.n298 12.8005
R285 VTAIL.n371 VTAIL.n296 12.8005
R286 VTAIL.n34 VTAIL.n30 12.8005
R287 VTAIL.n78 VTAIL.n10 12.8005
R288 VTAIL.n83 VTAIL.n8 12.8005
R289 VTAIL.n277 VTAIL.n202 12.8005
R290 VTAIL.n272 VTAIL.n204 12.8005
R291 VTAIL.n229 VTAIL.n225 12.8005
R292 VTAIL.n181 VTAIL.n106 12.8005
R293 VTAIL.n176 VTAIL.n108 12.8005
R294 VTAIL.n133 VTAIL.n129 12.8005
R295 VTAIL.n326 VTAIL.n325 12.0247
R296 VTAIL.n363 VTAIL.n362 12.0247
R297 VTAIL.n372 VTAIL.n294 12.0247
R298 VTAIL.n38 VTAIL.n37 12.0247
R299 VTAIL.n75 VTAIL.n74 12.0247
R300 VTAIL.n84 VTAIL.n6 12.0247
R301 VTAIL.n278 VTAIL.n200 12.0247
R302 VTAIL.n269 VTAIL.n268 12.0247
R303 VTAIL.n233 VTAIL.n232 12.0247
R304 VTAIL.n182 VTAIL.n104 12.0247
R305 VTAIL.n173 VTAIL.n172 12.0247
R306 VTAIL.n137 VTAIL.n136 12.0247
R307 VTAIL.n329 VTAIL.n316 11.249
R308 VTAIL.n358 VTAIL.n300 11.249
R309 VTAIL.n376 VTAIL.n375 11.249
R310 VTAIL.n41 VTAIL.n28 11.249
R311 VTAIL.n70 VTAIL.n12 11.249
R312 VTAIL.n88 VTAIL.n87 11.249
R313 VTAIL.n282 VTAIL.n281 11.249
R314 VTAIL.n265 VTAIL.n206 11.249
R315 VTAIL.n236 VTAIL.n223 11.249
R316 VTAIL.n186 VTAIL.n185 11.249
R317 VTAIL.n169 VTAIL.n110 11.249
R318 VTAIL.n140 VTAIL.n127 11.249
R319 VTAIL.n330 VTAIL.n314 10.4732
R320 VTAIL.n357 VTAIL.n302 10.4732
R321 VTAIL.n379 VTAIL.n292 10.4732
R322 VTAIL.n42 VTAIL.n26 10.4732
R323 VTAIL.n69 VTAIL.n14 10.4732
R324 VTAIL.n91 VTAIL.n4 10.4732
R325 VTAIL.n285 VTAIL.n198 10.4732
R326 VTAIL.n264 VTAIL.n209 10.4732
R327 VTAIL.n237 VTAIL.n221 10.4732
R328 VTAIL.n189 VTAIL.n102 10.4732
R329 VTAIL.n168 VTAIL.n113 10.4732
R330 VTAIL.n141 VTAIL.n125 10.4732
R331 VTAIL.n334 VTAIL.n333 9.69747
R332 VTAIL.n354 VTAIL.n353 9.69747
R333 VTAIL.n380 VTAIL.n290 9.69747
R334 VTAIL.n46 VTAIL.n45 9.69747
R335 VTAIL.n66 VTAIL.n65 9.69747
R336 VTAIL.n92 VTAIL.n2 9.69747
R337 VTAIL.n286 VTAIL.n196 9.69747
R338 VTAIL.n261 VTAIL.n260 9.69747
R339 VTAIL.n241 VTAIL.n240 9.69747
R340 VTAIL.n190 VTAIL.n100 9.69747
R341 VTAIL.n165 VTAIL.n164 9.69747
R342 VTAIL.n145 VTAIL.n144 9.69747
R343 VTAIL.n382 VTAIL.n381 9.45567
R344 VTAIL.n94 VTAIL.n93 9.45567
R345 VTAIL.n288 VTAIL.n287 9.45567
R346 VTAIL.n192 VTAIL.n191 9.45567
R347 VTAIL.n381 VTAIL.n380 9.3005
R348 VTAIL.n292 VTAIL.n291 9.3005
R349 VTAIL.n375 VTAIL.n374 9.3005
R350 VTAIL.n373 VTAIL.n372 9.3005
R351 VTAIL.n296 VTAIL.n295 9.3005
R352 VTAIL.n341 VTAIL.n340 9.3005
R353 VTAIL.n339 VTAIL.n338 9.3005
R354 VTAIL.n312 VTAIL.n311 9.3005
R355 VTAIL.n333 VTAIL.n332 9.3005
R356 VTAIL.n331 VTAIL.n330 9.3005
R357 VTAIL.n316 VTAIL.n315 9.3005
R358 VTAIL.n325 VTAIL.n324 9.3005
R359 VTAIL.n323 VTAIL.n322 9.3005
R360 VTAIL.n308 VTAIL.n307 9.3005
R361 VTAIL.n347 VTAIL.n346 9.3005
R362 VTAIL.n349 VTAIL.n348 9.3005
R363 VTAIL.n304 VTAIL.n303 9.3005
R364 VTAIL.n355 VTAIL.n354 9.3005
R365 VTAIL.n357 VTAIL.n356 9.3005
R366 VTAIL.n300 VTAIL.n299 9.3005
R367 VTAIL.n364 VTAIL.n363 9.3005
R368 VTAIL.n366 VTAIL.n365 9.3005
R369 VTAIL.n93 VTAIL.n92 9.3005
R370 VTAIL.n4 VTAIL.n3 9.3005
R371 VTAIL.n87 VTAIL.n86 9.3005
R372 VTAIL.n85 VTAIL.n84 9.3005
R373 VTAIL.n8 VTAIL.n7 9.3005
R374 VTAIL.n53 VTAIL.n52 9.3005
R375 VTAIL.n51 VTAIL.n50 9.3005
R376 VTAIL.n24 VTAIL.n23 9.3005
R377 VTAIL.n45 VTAIL.n44 9.3005
R378 VTAIL.n43 VTAIL.n42 9.3005
R379 VTAIL.n28 VTAIL.n27 9.3005
R380 VTAIL.n37 VTAIL.n36 9.3005
R381 VTAIL.n35 VTAIL.n34 9.3005
R382 VTAIL.n20 VTAIL.n19 9.3005
R383 VTAIL.n59 VTAIL.n58 9.3005
R384 VTAIL.n61 VTAIL.n60 9.3005
R385 VTAIL.n16 VTAIL.n15 9.3005
R386 VTAIL.n67 VTAIL.n66 9.3005
R387 VTAIL.n69 VTAIL.n68 9.3005
R388 VTAIL.n12 VTAIL.n11 9.3005
R389 VTAIL.n76 VTAIL.n75 9.3005
R390 VTAIL.n78 VTAIL.n77 9.3005
R391 VTAIL.n254 VTAIL.n253 9.3005
R392 VTAIL.n256 VTAIL.n255 9.3005
R393 VTAIL.n211 VTAIL.n210 9.3005
R394 VTAIL.n262 VTAIL.n261 9.3005
R395 VTAIL.n264 VTAIL.n263 9.3005
R396 VTAIL.n206 VTAIL.n205 9.3005
R397 VTAIL.n270 VTAIL.n269 9.3005
R398 VTAIL.n272 VTAIL.n271 9.3005
R399 VTAIL.n287 VTAIL.n286 9.3005
R400 VTAIL.n198 VTAIL.n197 9.3005
R401 VTAIL.n281 VTAIL.n280 9.3005
R402 VTAIL.n279 VTAIL.n278 9.3005
R403 VTAIL.n202 VTAIL.n201 9.3005
R404 VTAIL.n215 VTAIL.n214 9.3005
R405 VTAIL.n248 VTAIL.n247 9.3005
R406 VTAIL.n246 VTAIL.n245 9.3005
R407 VTAIL.n219 VTAIL.n218 9.3005
R408 VTAIL.n240 VTAIL.n239 9.3005
R409 VTAIL.n238 VTAIL.n237 9.3005
R410 VTAIL.n223 VTAIL.n222 9.3005
R411 VTAIL.n232 VTAIL.n231 9.3005
R412 VTAIL.n230 VTAIL.n229 9.3005
R413 VTAIL.n158 VTAIL.n157 9.3005
R414 VTAIL.n160 VTAIL.n159 9.3005
R415 VTAIL.n115 VTAIL.n114 9.3005
R416 VTAIL.n166 VTAIL.n165 9.3005
R417 VTAIL.n168 VTAIL.n167 9.3005
R418 VTAIL.n110 VTAIL.n109 9.3005
R419 VTAIL.n174 VTAIL.n173 9.3005
R420 VTAIL.n176 VTAIL.n175 9.3005
R421 VTAIL.n191 VTAIL.n190 9.3005
R422 VTAIL.n102 VTAIL.n101 9.3005
R423 VTAIL.n185 VTAIL.n184 9.3005
R424 VTAIL.n183 VTAIL.n182 9.3005
R425 VTAIL.n106 VTAIL.n105 9.3005
R426 VTAIL.n119 VTAIL.n118 9.3005
R427 VTAIL.n152 VTAIL.n151 9.3005
R428 VTAIL.n150 VTAIL.n149 9.3005
R429 VTAIL.n123 VTAIL.n122 9.3005
R430 VTAIL.n144 VTAIL.n143 9.3005
R431 VTAIL.n142 VTAIL.n141 9.3005
R432 VTAIL.n127 VTAIL.n126 9.3005
R433 VTAIL.n136 VTAIL.n135 9.3005
R434 VTAIL.n134 VTAIL.n133 9.3005
R435 VTAIL.n337 VTAIL.n312 8.92171
R436 VTAIL.n350 VTAIL.n304 8.92171
R437 VTAIL.n49 VTAIL.n24 8.92171
R438 VTAIL.n62 VTAIL.n16 8.92171
R439 VTAIL.n257 VTAIL.n211 8.92171
R440 VTAIL.n244 VTAIL.n219 8.92171
R441 VTAIL.n161 VTAIL.n115 8.92171
R442 VTAIL.n148 VTAIL.n123 8.92171
R443 VTAIL.n338 VTAIL.n310 8.14595
R444 VTAIL.n349 VTAIL.n306 8.14595
R445 VTAIL.n50 VTAIL.n22 8.14595
R446 VTAIL.n61 VTAIL.n18 8.14595
R447 VTAIL.n256 VTAIL.n213 8.14595
R448 VTAIL.n245 VTAIL.n217 8.14595
R449 VTAIL.n160 VTAIL.n117 8.14595
R450 VTAIL.n149 VTAIL.n121 8.14595
R451 VTAIL.n342 VTAIL.n341 7.3702
R452 VTAIL.n346 VTAIL.n345 7.3702
R453 VTAIL.n54 VTAIL.n53 7.3702
R454 VTAIL.n58 VTAIL.n57 7.3702
R455 VTAIL.n253 VTAIL.n252 7.3702
R456 VTAIL.n249 VTAIL.n248 7.3702
R457 VTAIL.n157 VTAIL.n156 7.3702
R458 VTAIL.n153 VTAIL.n152 7.3702
R459 VTAIL.n342 VTAIL.n308 6.59444
R460 VTAIL.n345 VTAIL.n308 6.59444
R461 VTAIL.n54 VTAIL.n20 6.59444
R462 VTAIL.n57 VTAIL.n20 6.59444
R463 VTAIL.n252 VTAIL.n215 6.59444
R464 VTAIL.n249 VTAIL.n215 6.59444
R465 VTAIL.n156 VTAIL.n119 6.59444
R466 VTAIL.n153 VTAIL.n119 6.59444
R467 VTAIL.n341 VTAIL.n310 5.81868
R468 VTAIL.n346 VTAIL.n306 5.81868
R469 VTAIL.n53 VTAIL.n22 5.81868
R470 VTAIL.n58 VTAIL.n18 5.81868
R471 VTAIL.n253 VTAIL.n213 5.81868
R472 VTAIL.n248 VTAIL.n217 5.81868
R473 VTAIL.n157 VTAIL.n117 5.81868
R474 VTAIL.n152 VTAIL.n121 5.81868
R475 VTAIL.n338 VTAIL.n337 5.04292
R476 VTAIL.n350 VTAIL.n349 5.04292
R477 VTAIL.n50 VTAIL.n49 5.04292
R478 VTAIL.n62 VTAIL.n61 5.04292
R479 VTAIL.n257 VTAIL.n256 5.04292
R480 VTAIL.n245 VTAIL.n244 5.04292
R481 VTAIL.n161 VTAIL.n160 5.04292
R482 VTAIL.n149 VTAIL.n148 5.04292
R483 VTAIL.n334 VTAIL.n312 4.26717
R484 VTAIL.n353 VTAIL.n304 4.26717
R485 VTAIL.n382 VTAIL.n290 4.26717
R486 VTAIL.n46 VTAIL.n24 4.26717
R487 VTAIL.n65 VTAIL.n16 4.26717
R488 VTAIL.n94 VTAIL.n2 4.26717
R489 VTAIL.n288 VTAIL.n196 4.26717
R490 VTAIL.n260 VTAIL.n211 4.26717
R491 VTAIL.n241 VTAIL.n219 4.26717
R492 VTAIL.n192 VTAIL.n100 4.26717
R493 VTAIL.n164 VTAIL.n115 4.26717
R494 VTAIL.n145 VTAIL.n123 4.26717
R495 VTAIL.n323 VTAIL.n319 3.70982
R496 VTAIL.n35 VTAIL.n31 3.70982
R497 VTAIL.n230 VTAIL.n226 3.70982
R498 VTAIL.n134 VTAIL.n130 3.70982
R499 VTAIL.n333 VTAIL.n314 3.49141
R500 VTAIL.n354 VTAIL.n302 3.49141
R501 VTAIL.n380 VTAIL.n379 3.49141
R502 VTAIL.n45 VTAIL.n26 3.49141
R503 VTAIL.n66 VTAIL.n14 3.49141
R504 VTAIL.n92 VTAIL.n91 3.49141
R505 VTAIL.n286 VTAIL.n285 3.49141
R506 VTAIL.n261 VTAIL.n209 3.49141
R507 VTAIL.n240 VTAIL.n221 3.49141
R508 VTAIL.n190 VTAIL.n189 3.49141
R509 VTAIL.n165 VTAIL.n113 3.49141
R510 VTAIL.n144 VTAIL.n125 3.49141
R511 VTAIL.n193 VTAIL.n99 2.89705
R512 VTAIL.n289 VTAIL.n195 2.89705
R513 VTAIL.n97 VTAIL.n95 2.89705
R514 VTAIL.n330 VTAIL.n329 2.71565
R515 VTAIL.n358 VTAIL.n357 2.71565
R516 VTAIL.n376 VTAIL.n292 2.71565
R517 VTAIL.n42 VTAIL.n41 2.71565
R518 VTAIL.n70 VTAIL.n69 2.71565
R519 VTAIL.n88 VTAIL.n4 2.71565
R520 VTAIL.n282 VTAIL.n198 2.71565
R521 VTAIL.n265 VTAIL.n264 2.71565
R522 VTAIL.n237 VTAIL.n236 2.71565
R523 VTAIL.n186 VTAIL.n102 2.71565
R524 VTAIL.n169 VTAIL.n168 2.71565
R525 VTAIL.n141 VTAIL.n140 2.71565
R526 VTAIL VTAIL.n383 2.11472
R527 VTAIL.n326 VTAIL.n316 1.93989
R528 VTAIL.n362 VTAIL.n300 1.93989
R529 VTAIL.n375 VTAIL.n294 1.93989
R530 VTAIL.n38 VTAIL.n28 1.93989
R531 VTAIL.n74 VTAIL.n12 1.93989
R532 VTAIL.n87 VTAIL.n6 1.93989
R533 VTAIL.n281 VTAIL.n200 1.93989
R534 VTAIL.n268 VTAIL.n206 1.93989
R535 VTAIL.n233 VTAIL.n223 1.93989
R536 VTAIL.n185 VTAIL.n104 1.93989
R537 VTAIL.n172 VTAIL.n110 1.93989
R538 VTAIL.n137 VTAIL.n127 1.93989
R539 VTAIL.n0 VTAIL.t5 1.9216
R540 VTAIL.n0 VTAIL.t3 1.9216
R541 VTAIL.n96 VTAIL.t8 1.9216
R542 VTAIL.n96 VTAIL.t7 1.9216
R543 VTAIL.n194 VTAIL.t10 1.9216
R544 VTAIL.n194 VTAIL.t11 1.9216
R545 VTAIL.n98 VTAIL.t0 1.9216
R546 VTAIL.n98 VTAIL.t1 1.9216
R547 VTAIL.n195 VTAIL.n193 1.9186
R548 VTAIL.n95 VTAIL.n1 1.9186
R549 VTAIL.n325 VTAIL.n318 1.16414
R550 VTAIL.n363 VTAIL.n298 1.16414
R551 VTAIL.n372 VTAIL.n371 1.16414
R552 VTAIL.n37 VTAIL.n30 1.16414
R553 VTAIL.n75 VTAIL.n10 1.16414
R554 VTAIL.n84 VTAIL.n83 1.16414
R555 VTAIL.n278 VTAIL.n277 1.16414
R556 VTAIL.n269 VTAIL.n204 1.16414
R557 VTAIL.n232 VTAIL.n225 1.16414
R558 VTAIL.n182 VTAIL.n181 1.16414
R559 VTAIL.n173 VTAIL.n108 1.16414
R560 VTAIL.n136 VTAIL.n129 1.16414
R561 VTAIL VTAIL.n1 0.782828
R562 VTAIL.n322 VTAIL.n321 0.388379
R563 VTAIL.n367 VTAIL.n366 0.388379
R564 VTAIL.n368 VTAIL.n296 0.388379
R565 VTAIL.n34 VTAIL.n33 0.388379
R566 VTAIL.n79 VTAIL.n78 0.388379
R567 VTAIL.n80 VTAIL.n8 0.388379
R568 VTAIL.n274 VTAIL.n202 0.388379
R569 VTAIL.n273 VTAIL.n272 0.388379
R570 VTAIL.n229 VTAIL.n228 0.388379
R571 VTAIL.n178 VTAIL.n106 0.388379
R572 VTAIL.n177 VTAIL.n176 0.388379
R573 VTAIL.n133 VTAIL.n132 0.388379
R574 VTAIL.n324 VTAIL.n323 0.155672
R575 VTAIL.n324 VTAIL.n315 0.155672
R576 VTAIL.n331 VTAIL.n315 0.155672
R577 VTAIL.n332 VTAIL.n331 0.155672
R578 VTAIL.n332 VTAIL.n311 0.155672
R579 VTAIL.n339 VTAIL.n311 0.155672
R580 VTAIL.n340 VTAIL.n339 0.155672
R581 VTAIL.n340 VTAIL.n307 0.155672
R582 VTAIL.n347 VTAIL.n307 0.155672
R583 VTAIL.n348 VTAIL.n347 0.155672
R584 VTAIL.n348 VTAIL.n303 0.155672
R585 VTAIL.n355 VTAIL.n303 0.155672
R586 VTAIL.n356 VTAIL.n355 0.155672
R587 VTAIL.n356 VTAIL.n299 0.155672
R588 VTAIL.n364 VTAIL.n299 0.155672
R589 VTAIL.n365 VTAIL.n364 0.155672
R590 VTAIL.n365 VTAIL.n295 0.155672
R591 VTAIL.n373 VTAIL.n295 0.155672
R592 VTAIL.n374 VTAIL.n373 0.155672
R593 VTAIL.n374 VTAIL.n291 0.155672
R594 VTAIL.n381 VTAIL.n291 0.155672
R595 VTAIL.n36 VTAIL.n35 0.155672
R596 VTAIL.n36 VTAIL.n27 0.155672
R597 VTAIL.n43 VTAIL.n27 0.155672
R598 VTAIL.n44 VTAIL.n43 0.155672
R599 VTAIL.n44 VTAIL.n23 0.155672
R600 VTAIL.n51 VTAIL.n23 0.155672
R601 VTAIL.n52 VTAIL.n51 0.155672
R602 VTAIL.n52 VTAIL.n19 0.155672
R603 VTAIL.n59 VTAIL.n19 0.155672
R604 VTAIL.n60 VTAIL.n59 0.155672
R605 VTAIL.n60 VTAIL.n15 0.155672
R606 VTAIL.n67 VTAIL.n15 0.155672
R607 VTAIL.n68 VTAIL.n67 0.155672
R608 VTAIL.n68 VTAIL.n11 0.155672
R609 VTAIL.n76 VTAIL.n11 0.155672
R610 VTAIL.n77 VTAIL.n76 0.155672
R611 VTAIL.n77 VTAIL.n7 0.155672
R612 VTAIL.n85 VTAIL.n7 0.155672
R613 VTAIL.n86 VTAIL.n85 0.155672
R614 VTAIL.n86 VTAIL.n3 0.155672
R615 VTAIL.n93 VTAIL.n3 0.155672
R616 VTAIL.n287 VTAIL.n197 0.155672
R617 VTAIL.n280 VTAIL.n197 0.155672
R618 VTAIL.n280 VTAIL.n279 0.155672
R619 VTAIL.n279 VTAIL.n201 0.155672
R620 VTAIL.n271 VTAIL.n201 0.155672
R621 VTAIL.n271 VTAIL.n270 0.155672
R622 VTAIL.n270 VTAIL.n205 0.155672
R623 VTAIL.n263 VTAIL.n205 0.155672
R624 VTAIL.n263 VTAIL.n262 0.155672
R625 VTAIL.n262 VTAIL.n210 0.155672
R626 VTAIL.n255 VTAIL.n210 0.155672
R627 VTAIL.n255 VTAIL.n254 0.155672
R628 VTAIL.n254 VTAIL.n214 0.155672
R629 VTAIL.n247 VTAIL.n214 0.155672
R630 VTAIL.n247 VTAIL.n246 0.155672
R631 VTAIL.n246 VTAIL.n218 0.155672
R632 VTAIL.n239 VTAIL.n218 0.155672
R633 VTAIL.n239 VTAIL.n238 0.155672
R634 VTAIL.n238 VTAIL.n222 0.155672
R635 VTAIL.n231 VTAIL.n222 0.155672
R636 VTAIL.n231 VTAIL.n230 0.155672
R637 VTAIL.n191 VTAIL.n101 0.155672
R638 VTAIL.n184 VTAIL.n101 0.155672
R639 VTAIL.n184 VTAIL.n183 0.155672
R640 VTAIL.n183 VTAIL.n105 0.155672
R641 VTAIL.n175 VTAIL.n105 0.155672
R642 VTAIL.n175 VTAIL.n174 0.155672
R643 VTAIL.n174 VTAIL.n109 0.155672
R644 VTAIL.n167 VTAIL.n109 0.155672
R645 VTAIL.n167 VTAIL.n166 0.155672
R646 VTAIL.n166 VTAIL.n114 0.155672
R647 VTAIL.n159 VTAIL.n114 0.155672
R648 VTAIL.n159 VTAIL.n158 0.155672
R649 VTAIL.n158 VTAIL.n118 0.155672
R650 VTAIL.n151 VTAIL.n118 0.155672
R651 VTAIL.n151 VTAIL.n150 0.155672
R652 VTAIL.n150 VTAIL.n122 0.155672
R653 VTAIL.n143 VTAIL.n122 0.155672
R654 VTAIL.n143 VTAIL.n142 0.155672
R655 VTAIL.n142 VTAIL.n126 0.155672
R656 VTAIL.n135 VTAIL.n126 0.155672
R657 VTAIL.n135 VTAIL.n134 0.155672
R658 VDD1.n88 VDD1.n0 756.745
R659 VDD1.n181 VDD1.n93 756.745
R660 VDD1.n89 VDD1.n88 585
R661 VDD1.n87 VDD1.n86 585
R662 VDD1.n4 VDD1.n3 585
R663 VDD1.n81 VDD1.n80 585
R664 VDD1.n79 VDD1.n78 585
R665 VDD1.n77 VDD1.n7 585
R666 VDD1.n11 VDD1.n8 585
R667 VDD1.n72 VDD1.n71 585
R668 VDD1.n70 VDD1.n69 585
R669 VDD1.n13 VDD1.n12 585
R670 VDD1.n64 VDD1.n63 585
R671 VDD1.n62 VDD1.n61 585
R672 VDD1.n17 VDD1.n16 585
R673 VDD1.n56 VDD1.n55 585
R674 VDD1.n54 VDD1.n53 585
R675 VDD1.n21 VDD1.n20 585
R676 VDD1.n48 VDD1.n47 585
R677 VDD1.n46 VDD1.n45 585
R678 VDD1.n25 VDD1.n24 585
R679 VDD1.n40 VDD1.n39 585
R680 VDD1.n38 VDD1.n37 585
R681 VDD1.n29 VDD1.n28 585
R682 VDD1.n32 VDD1.n31 585
R683 VDD1.n124 VDD1.n123 585
R684 VDD1.n121 VDD1.n120 585
R685 VDD1.n130 VDD1.n129 585
R686 VDD1.n132 VDD1.n131 585
R687 VDD1.n117 VDD1.n116 585
R688 VDD1.n138 VDD1.n137 585
R689 VDD1.n140 VDD1.n139 585
R690 VDD1.n113 VDD1.n112 585
R691 VDD1.n146 VDD1.n145 585
R692 VDD1.n148 VDD1.n147 585
R693 VDD1.n109 VDD1.n108 585
R694 VDD1.n154 VDD1.n153 585
R695 VDD1.n156 VDD1.n155 585
R696 VDD1.n105 VDD1.n104 585
R697 VDD1.n162 VDD1.n161 585
R698 VDD1.n165 VDD1.n164 585
R699 VDD1.n163 VDD1.n101 585
R700 VDD1.n170 VDD1.n100 585
R701 VDD1.n172 VDD1.n171 585
R702 VDD1.n174 VDD1.n173 585
R703 VDD1.n97 VDD1.n96 585
R704 VDD1.n180 VDD1.n179 585
R705 VDD1.n182 VDD1.n181 585
R706 VDD1.t1 VDD1.n30 327.466
R707 VDD1.t4 VDD1.n122 327.466
R708 VDD1.n88 VDD1.n87 171.744
R709 VDD1.n87 VDD1.n3 171.744
R710 VDD1.n80 VDD1.n3 171.744
R711 VDD1.n80 VDD1.n79 171.744
R712 VDD1.n79 VDD1.n7 171.744
R713 VDD1.n11 VDD1.n7 171.744
R714 VDD1.n71 VDD1.n11 171.744
R715 VDD1.n71 VDD1.n70 171.744
R716 VDD1.n70 VDD1.n12 171.744
R717 VDD1.n63 VDD1.n12 171.744
R718 VDD1.n63 VDD1.n62 171.744
R719 VDD1.n62 VDD1.n16 171.744
R720 VDD1.n55 VDD1.n16 171.744
R721 VDD1.n55 VDD1.n54 171.744
R722 VDD1.n54 VDD1.n20 171.744
R723 VDD1.n47 VDD1.n20 171.744
R724 VDD1.n47 VDD1.n46 171.744
R725 VDD1.n46 VDD1.n24 171.744
R726 VDD1.n39 VDD1.n24 171.744
R727 VDD1.n39 VDD1.n38 171.744
R728 VDD1.n38 VDD1.n28 171.744
R729 VDD1.n31 VDD1.n28 171.744
R730 VDD1.n123 VDD1.n120 171.744
R731 VDD1.n130 VDD1.n120 171.744
R732 VDD1.n131 VDD1.n130 171.744
R733 VDD1.n131 VDD1.n116 171.744
R734 VDD1.n138 VDD1.n116 171.744
R735 VDD1.n139 VDD1.n138 171.744
R736 VDD1.n139 VDD1.n112 171.744
R737 VDD1.n146 VDD1.n112 171.744
R738 VDD1.n147 VDD1.n146 171.744
R739 VDD1.n147 VDD1.n108 171.744
R740 VDD1.n154 VDD1.n108 171.744
R741 VDD1.n155 VDD1.n154 171.744
R742 VDD1.n155 VDD1.n104 171.744
R743 VDD1.n162 VDD1.n104 171.744
R744 VDD1.n164 VDD1.n162 171.744
R745 VDD1.n164 VDD1.n163 171.744
R746 VDD1.n163 VDD1.n100 171.744
R747 VDD1.n172 VDD1.n100 171.744
R748 VDD1.n173 VDD1.n172 171.744
R749 VDD1.n173 VDD1.n96 171.744
R750 VDD1.n180 VDD1.n96 171.744
R751 VDD1.n181 VDD1.n180 171.744
R752 VDD1.n31 VDD1.t1 85.8723
R753 VDD1.n123 VDD1.t4 85.8723
R754 VDD1.n187 VDD1.n186 72.3879
R755 VDD1.n189 VDD1.n188 71.7191
R756 VDD1 VDD1.n92 53.422
R757 VDD1.n187 VDD1.n185 53.3085
R758 VDD1.n189 VDD1.n187 49.7466
R759 VDD1.n32 VDD1.n30 16.3895
R760 VDD1.n124 VDD1.n122 16.3895
R761 VDD1.n78 VDD1.n77 13.1884
R762 VDD1.n171 VDD1.n170 13.1884
R763 VDD1.n81 VDD1.n6 12.8005
R764 VDD1.n76 VDD1.n8 12.8005
R765 VDD1.n33 VDD1.n29 12.8005
R766 VDD1.n125 VDD1.n121 12.8005
R767 VDD1.n169 VDD1.n101 12.8005
R768 VDD1.n174 VDD1.n99 12.8005
R769 VDD1.n82 VDD1.n4 12.0247
R770 VDD1.n73 VDD1.n72 12.0247
R771 VDD1.n37 VDD1.n36 12.0247
R772 VDD1.n129 VDD1.n128 12.0247
R773 VDD1.n166 VDD1.n165 12.0247
R774 VDD1.n175 VDD1.n97 12.0247
R775 VDD1.n86 VDD1.n85 11.249
R776 VDD1.n69 VDD1.n10 11.249
R777 VDD1.n40 VDD1.n27 11.249
R778 VDD1.n132 VDD1.n119 11.249
R779 VDD1.n161 VDD1.n103 11.249
R780 VDD1.n179 VDD1.n178 11.249
R781 VDD1.n89 VDD1.n2 10.4732
R782 VDD1.n68 VDD1.n13 10.4732
R783 VDD1.n41 VDD1.n25 10.4732
R784 VDD1.n133 VDD1.n117 10.4732
R785 VDD1.n160 VDD1.n105 10.4732
R786 VDD1.n182 VDD1.n95 10.4732
R787 VDD1.n90 VDD1.n0 9.69747
R788 VDD1.n65 VDD1.n64 9.69747
R789 VDD1.n45 VDD1.n44 9.69747
R790 VDD1.n137 VDD1.n136 9.69747
R791 VDD1.n157 VDD1.n156 9.69747
R792 VDD1.n183 VDD1.n93 9.69747
R793 VDD1.n92 VDD1.n91 9.45567
R794 VDD1.n185 VDD1.n184 9.45567
R795 VDD1.n58 VDD1.n57 9.3005
R796 VDD1.n60 VDD1.n59 9.3005
R797 VDD1.n15 VDD1.n14 9.3005
R798 VDD1.n66 VDD1.n65 9.3005
R799 VDD1.n68 VDD1.n67 9.3005
R800 VDD1.n10 VDD1.n9 9.3005
R801 VDD1.n74 VDD1.n73 9.3005
R802 VDD1.n76 VDD1.n75 9.3005
R803 VDD1.n91 VDD1.n90 9.3005
R804 VDD1.n2 VDD1.n1 9.3005
R805 VDD1.n85 VDD1.n84 9.3005
R806 VDD1.n83 VDD1.n82 9.3005
R807 VDD1.n6 VDD1.n5 9.3005
R808 VDD1.n19 VDD1.n18 9.3005
R809 VDD1.n52 VDD1.n51 9.3005
R810 VDD1.n50 VDD1.n49 9.3005
R811 VDD1.n23 VDD1.n22 9.3005
R812 VDD1.n44 VDD1.n43 9.3005
R813 VDD1.n42 VDD1.n41 9.3005
R814 VDD1.n27 VDD1.n26 9.3005
R815 VDD1.n36 VDD1.n35 9.3005
R816 VDD1.n34 VDD1.n33 9.3005
R817 VDD1.n184 VDD1.n183 9.3005
R818 VDD1.n95 VDD1.n94 9.3005
R819 VDD1.n178 VDD1.n177 9.3005
R820 VDD1.n176 VDD1.n175 9.3005
R821 VDD1.n99 VDD1.n98 9.3005
R822 VDD1.n144 VDD1.n143 9.3005
R823 VDD1.n142 VDD1.n141 9.3005
R824 VDD1.n115 VDD1.n114 9.3005
R825 VDD1.n136 VDD1.n135 9.3005
R826 VDD1.n134 VDD1.n133 9.3005
R827 VDD1.n119 VDD1.n118 9.3005
R828 VDD1.n128 VDD1.n127 9.3005
R829 VDD1.n126 VDD1.n125 9.3005
R830 VDD1.n111 VDD1.n110 9.3005
R831 VDD1.n150 VDD1.n149 9.3005
R832 VDD1.n152 VDD1.n151 9.3005
R833 VDD1.n107 VDD1.n106 9.3005
R834 VDD1.n158 VDD1.n157 9.3005
R835 VDD1.n160 VDD1.n159 9.3005
R836 VDD1.n103 VDD1.n102 9.3005
R837 VDD1.n167 VDD1.n166 9.3005
R838 VDD1.n169 VDD1.n168 9.3005
R839 VDD1.n61 VDD1.n15 8.92171
R840 VDD1.n48 VDD1.n23 8.92171
R841 VDD1.n140 VDD1.n115 8.92171
R842 VDD1.n153 VDD1.n107 8.92171
R843 VDD1.n60 VDD1.n17 8.14595
R844 VDD1.n49 VDD1.n21 8.14595
R845 VDD1.n141 VDD1.n113 8.14595
R846 VDD1.n152 VDD1.n109 8.14595
R847 VDD1.n57 VDD1.n56 7.3702
R848 VDD1.n53 VDD1.n52 7.3702
R849 VDD1.n145 VDD1.n144 7.3702
R850 VDD1.n149 VDD1.n148 7.3702
R851 VDD1.n56 VDD1.n19 6.59444
R852 VDD1.n53 VDD1.n19 6.59444
R853 VDD1.n145 VDD1.n111 6.59444
R854 VDD1.n148 VDD1.n111 6.59444
R855 VDD1.n57 VDD1.n17 5.81868
R856 VDD1.n52 VDD1.n21 5.81868
R857 VDD1.n144 VDD1.n113 5.81868
R858 VDD1.n149 VDD1.n109 5.81868
R859 VDD1.n61 VDD1.n60 5.04292
R860 VDD1.n49 VDD1.n48 5.04292
R861 VDD1.n141 VDD1.n140 5.04292
R862 VDD1.n153 VDD1.n152 5.04292
R863 VDD1.n92 VDD1.n0 4.26717
R864 VDD1.n64 VDD1.n15 4.26717
R865 VDD1.n45 VDD1.n23 4.26717
R866 VDD1.n137 VDD1.n115 4.26717
R867 VDD1.n156 VDD1.n107 4.26717
R868 VDD1.n185 VDD1.n93 4.26717
R869 VDD1.n34 VDD1.n30 3.70982
R870 VDD1.n126 VDD1.n122 3.70982
R871 VDD1.n90 VDD1.n89 3.49141
R872 VDD1.n65 VDD1.n13 3.49141
R873 VDD1.n44 VDD1.n25 3.49141
R874 VDD1.n136 VDD1.n117 3.49141
R875 VDD1.n157 VDD1.n105 3.49141
R876 VDD1.n183 VDD1.n182 3.49141
R877 VDD1.n86 VDD1.n2 2.71565
R878 VDD1.n69 VDD1.n68 2.71565
R879 VDD1.n41 VDD1.n40 2.71565
R880 VDD1.n133 VDD1.n132 2.71565
R881 VDD1.n161 VDD1.n160 2.71565
R882 VDD1.n179 VDD1.n95 2.71565
R883 VDD1.n85 VDD1.n4 1.93989
R884 VDD1.n72 VDD1.n10 1.93989
R885 VDD1.n37 VDD1.n27 1.93989
R886 VDD1.n129 VDD1.n119 1.93989
R887 VDD1.n165 VDD1.n103 1.93989
R888 VDD1.n178 VDD1.n97 1.93989
R889 VDD1.n188 VDD1.t2 1.9216
R890 VDD1.n188 VDD1.t5 1.9216
R891 VDD1.n186 VDD1.t3 1.9216
R892 VDD1.n186 VDD1.t0 1.9216
R893 VDD1.n82 VDD1.n81 1.16414
R894 VDD1.n73 VDD1.n8 1.16414
R895 VDD1.n36 VDD1.n29 1.16414
R896 VDD1.n128 VDD1.n121 1.16414
R897 VDD1.n166 VDD1.n101 1.16414
R898 VDD1.n175 VDD1.n174 1.16414
R899 VDD1 VDD1.n189 0.666448
R900 VDD1.n78 VDD1.n6 0.388379
R901 VDD1.n77 VDD1.n76 0.388379
R902 VDD1.n33 VDD1.n32 0.388379
R903 VDD1.n125 VDD1.n124 0.388379
R904 VDD1.n170 VDD1.n169 0.388379
R905 VDD1.n171 VDD1.n99 0.388379
R906 VDD1.n91 VDD1.n1 0.155672
R907 VDD1.n84 VDD1.n1 0.155672
R908 VDD1.n84 VDD1.n83 0.155672
R909 VDD1.n83 VDD1.n5 0.155672
R910 VDD1.n75 VDD1.n5 0.155672
R911 VDD1.n75 VDD1.n74 0.155672
R912 VDD1.n74 VDD1.n9 0.155672
R913 VDD1.n67 VDD1.n9 0.155672
R914 VDD1.n67 VDD1.n66 0.155672
R915 VDD1.n66 VDD1.n14 0.155672
R916 VDD1.n59 VDD1.n14 0.155672
R917 VDD1.n59 VDD1.n58 0.155672
R918 VDD1.n58 VDD1.n18 0.155672
R919 VDD1.n51 VDD1.n18 0.155672
R920 VDD1.n51 VDD1.n50 0.155672
R921 VDD1.n50 VDD1.n22 0.155672
R922 VDD1.n43 VDD1.n22 0.155672
R923 VDD1.n43 VDD1.n42 0.155672
R924 VDD1.n42 VDD1.n26 0.155672
R925 VDD1.n35 VDD1.n26 0.155672
R926 VDD1.n35 VDD1.n34 0.155672
R927 VDD1.n127 VDD1.n126 0.155672
R928 VDD1.n127 VDD1.n118 0.155672
R929 VDD1.n134 VDD1.n118 0.155672
R930 VDD1.n135 VDD1.n134 0.155672
R931 VDD1.n135 VDD1.n114 0.155672
R932 VDD1.n142 VDD1.n114 0.155672
R933 VDD1.n143 VDD1.n142 0.155672
R934 VDD1.n143 VDD1.n110 0.155672
R935 VDD1.n150 VDD1.n110 0.155672
R936 VDD1.n151 VDD1.n150 0.155672
R937 VDD1.n151 VDD1.n106 0.155672
R938 VDD1.n158 VDD1.n106 0.155672
R939 VDD1.n159 VDD1.n158 0.155672
R940 VDD1.n159 VDD1.n102 0.155672
R941 VDD1.n167 VDD1.n102 0.155672
R942 VDD1.n168 VDD1.n167 0.155672
R943 VDD1.n168 VDD1.n98 0.155672
R944 VDD1.n176 VDD1.n98 0.155672
R945 VDD1.n177 VDD1.n176 0.155672
R946 VDD1.n177 VDD1.n94 0.155672
R947 VDD1.n184 VDD1.n94 0.155672
R948 VN.n20 VN.t3 167.808
R949 VN.n4 VN.t5 167.808
R950 VN.n30 VN.n29 161.3
R951 VN.n28 VN.n17 161.3
R952 VN.n27 VN.n26 161.3
R953 VN.n25 VN.n18 161.3
R954 VN.n24 VN.n23 161.3
R955 VN.n22 VN.n19 161.3
R956 VN.n14 VN.n13 161.3
R957 VN.n12 VN.n1 161.3
R958 VN.n11 VN.n10 161.3
R959 VN.n9 VN.n2 161.3
R960 VN.n8 VN.n7 161.3
R961 VN.n6 VN.n3 161.3
R962 VN.n5 VN.t2 134.578
R963 VN.n0 VN.t0 134.578
R964 VN.n21 VN.t4 134.578
R965 VN.n16 VN.t1 134.578
R966 VN.n15 VN.n0 72.3637
R967 VN.n31 VN.n16 72.3637
R968 VN.n11 VN.n2 56.4773
R969 VN.n27 VN.n18 56.4773
R970 VN VN.n31 54.3464
R971 VN.n5 VN.n4 49.1755
R972 VN.n21 VN.n20 49.1755
R973 VN.n6 VN.n5 24.3439
R974 VN.n7 VN.n6 24.3439
R975 VN.n7 VN.n2 24.3439
R976 VN.n12 VN.n11 24.3439
R977 VN.n13 VN.n12 24.3439
R978 VN.n23 VN.n18 24.3439
R979 VN.n23 VN.n22 24.3439
R980 VN.n22 VN.n21 24.3439
R981 VN.n29 VN.n28 24.3439
R982 VN.n28 VN.n27 24.3439
R983 VN.n13 VN.n0 17.5278
R984 VN.n29 VN.n16 17.5278
R985 VN.n20 VN.n19 4.04423
R986 VN.n4 VN.n3 4.04423
R987 VN.n31 VN.n30 0.355081
R988 VN.n15 VN.n14 0.355081
R989 VN VN.n15 0.26685
R990 VN.n30 VN.n17 0.189894
R991 VN.n26 VN.n17 0.189894
R992 VN.n26 VN.n25 0.189894
R993 VN.n25 VN.n24 0.189894
R994 VN.n24 VN.n19 0.189894
R995 VN.n8 VN.n3 0.189894
R996 VN.n9 VN.n8 0.189894
R997 VN.n10 VN.n9 0.189894
R998 VN.n10 VN.n1 0.189894
R999 VN.n14 VN.n1 0.189894
R1000 VDD2.n183 VDD2.n95 756.745
R1001 VDD2.n88 VDD2.n0 756.745
R1002 VDD2.n184 VDD2.n183 585
R1003 VDD2.n182 VDD2.n181 585
R1004 VDD2.n99 VDD2.n98 585
R1005 VDD2.n176 VDD2.n175 585
R1006 VDD2.n174 VDD2.n173 585
R1007 VDD2.n172 VDD2.n102 585
R1008 VDD2.n106 VDD2.n103 585
R1009 VDD2.n167 VDD2.n166 585
R1010 VDD2.n165 VDD2.n164 585
R1011 VDD2.n108 VDD2.n107 585
R1012 VDD2.n159 VDD2.n158 585
R1013 VDD2.n157 VDD2.n156 585
R1014 VDD2.n112 VDD2.n111 585
R1015 VDD2.n151 VDD2.n150 585
R1016 VDD2.n149 VDD2.n148 585
R1017 VDD2.n116 VDD2.n115 585
R1018 VDD2.n143 VDD2.n142 585
R1019 VDD2.n141 VDD2.n140 585
R1020 VDD2.n120 VDD2.n119 585
R1021 VDD2.n135 VDD2.n134 585
R1022 VDD2.n133 VDD2.n132 585
R1023 VDD2.n124 VDD2.n123 585
R1024 VDD2.n127 VDD2.n126 585
R1025 VDD2.n31 VDD2.n30 585
R1026 VDD2.n28 VDD2.n27 585
R1027 VDD2.n37 VDD2.n36 585
R1028 VDD2.n39 VDD2.n38 585
R1029 VDD2.n24 VDD2.n23 585
R1030 VDD2.n45 VDD2.n44 585
R1031 VDD2.n47 VDD2.n46 585
R1032 VDD2.n20 VDD2.n19 585
R1033 VDD2.n53 VDD2.n52 585
R1034 VDD2.n55 VDD2.n54 585
R1035 VDD2.n16 VDD2.n15 585
R1036 VDD2.n61 VDD2.n60 585
R1037 VDD2.n63 VDD2.n62 585
R1038 VDD2.n12 VDD2.n11 585
R1039 VDD2.n69 VDD2.n68 585
R1040 VDD2.n72 VDD2.n71 585
R1041 VDD2.n70 VDD2.n8 585
R1042 VDD2.n77 VDD2.n7 585
R1043 VDD2.n79 VDD2.n78 585
R1044 VDD2.n81 VDD2.n80 585
R1045 VDD2.n4 VDD2.n3 585
R1046 VDD2.n87 VDD2.n86 585
R1047 VDD2.n89 VDD2.n88 585
R1048 VDD2.t4 VDD2.n125 327.466
R1049 VDD2.t0 VDD2.n29 327.466
R1050 VDD2.n183 VDD2.n182 171.744
R1051 VDD2.n182 VDD2.n98 171.744
R1052 VDD2.n175 VDD2.n98 171.744
R1053 VDD2.n175 VDD2.n174 171.744
R1054 VDD2.n174 VDD2.n102 171.744
R1055 VDD2.n106 VDD2.n102 171.744
R1056 VDD2.n166 VDD2.n106 171.744
R1057 VDD2.n166 VDD2.n165 171.744
R1058 VDD2.n165 VDD2.n107 171.744
R1059 VDD2.n158 VDD2.n107 171.744
R1060 VDD2.n158 VDD2.n157 171.744
R1061 VDD2.n157 VDD2.n111 171.744
R1062 VDD2.n150 VDD2.n111 171.744
R1063 VDD2.n150 VDD2.n149 171.744
R1064 VDD2.n149 VDD2.n115 171.744
R1065 VDD2.n142 VDD2.n115 171.744
R1066 VDD2.n142 VDD2.n141 171.744
R1067 VDD2.n141 VDD2.n119 171.744
R1068 VDD2.n134 VDD2.n119 171.744
R1069 VDD2.n134 VDD2.n133 171.744
R1070 VDD2.n133 VDD2.n123 171.744
R1071 VDD2.n126 VDD2.n123 171.744
R1072 VDD2.n30 VDD2.n27 171.744
R1073 VDD2.n37 VDD2.n27 171.744
R1074 VDD2.n38 VDD2.n37 171.744
R1075 VDD2.n38 VDD2.n23 171.744
R1076 VDD2.n45 VDD2.n23 171.744
R1077 VDD2.n46 VDD2.n45 171.744
R1078 VDD2.n46 VDD2.n19 171.744
R1079 VDD2.n53 VDD2.n19 171.744
R1080 VDD2.n54 VDD2.n53 171.744
R1081 VDD2.n54 VDD2.n15 171.744
R1082 VDD2.n61 VDD2.n15 171.744
R1083 VDD2.n62 VDD2.n61 171.744
R1084 VDD2.n62 VDD2.n11 171.744
R1085 VDD2.n69 VDD2.n11 171.744
R1086 VDD2.n71 VDD2.n69 171.744
R1087 VDD2.n71 VDD2.n70 171.744
R1088 VDD2.n70 VDD2.n7 171.744
R1089 VDD2.n79 VDD2.n7 171.744
R1090 VDD2.n80 VDD2.n79 171.744
R1091 VDD2.n80 VDD2.n3 171.744
R1092 VDD2.n87 VDD2.n3 171.744
R1093 VDD2.n88 VDD2.n87 171.744
R1094 VDD2.n126 VDD2.t4 85.8723
R1095 VDD2.n30 VDD2.t0 85.8723
R1096 VDD2.n94 VDD2.n93 72.3879
R1097 VDD2 VDD2.n189 72.3851
R1098 VDD2.n94 VDD2.n92 53.3085
R1099 VDD2.n188 VDD2.n187 51.1914
R1100 VDD2.n188 VDD2.n94 47.7153
R1101 VDD2.n127 VDD2.n125 16.3895
R1102 VDD2.n31 VDD2.n29 16.3895
R1103 VDD2.n173 VDD2.n172 13.1884
R1104 VDD2.n78 VDD2.n77 13.1884
R1105 VDD2.n176 VDD2.n101 12.8005
R1106 VDD2.n171 VDD2.n103 12.8005
R1107 VDD2.n128 VDD2.n124 12.8005
R1108 VDD2.n32 VDD2.n28 12.8005
R1109 VDD2.n76 VDD2.n8 12.8005
R1110 VDD2.n81 VDD2.n6 12.8005
R1111 VDD2.n177 VDD2.n99 12.0247
R1112 VDD2.n168 VDD2.n167 12.0247
R1113 VDD2.n132 VDD2.n131 12.0247
R1114 VDD2.n36 VDD2.n35 12.0247
R1115 VDD2.n73 VDD2.n72 12.0247
R1116 VDD2.n82 VDD2.n4 12.0247
R1117 VDD2.n181 VDD2.n180 11.249
R1118 VDD2.n164 VDD2.n105 11.249
R1119 VDD2.n135 VDD2.n122 11.249
R1120 VDD2.n39 VDD2.n26 11.249
R1121 VDD2.n68 VDD2.n10 11.249
R1122 VDD2.n86 VDD2.n85 11.249
R1123 VDD2.n184 VDD2.n97 10.4732
R1124 VDD2.n163 VDD2.n108 10.4732
R1125 VDD2.n136 VDD2.n120 10.4732
R1126 VDD2.n40 VDD2.n24 10.4732
R1127 VDD2.n67 VDD2.n12 10.4732
R1128 VDD2.n89 VDD2.n2 10.4732
R1129 VDD2.n185 VDD2.n95 9.69747
R1130 VDD2.n160 VDD2.n159 9.69747
R1131 VDD2.n140 VDD2.n139 9.69747
R1132 VDD2.n44 VDD2.n43 9.69747
R1133 VDD2.n64 VDD2.n63 9.69747
R1134 VDD2.n90 VDD2.n0 9.69747
R1135 VDD2.n187 VDD2.n186 9.45567
R1136 VDD2.n92 VDD2.n91 9.45567
R1137 VDD2.n153 VDD2.n152 9.3005
R1138 VDD2.n155 VDD2.n154 9.3005
R1139 VDD2.n110 VDD2.n109 9.3005
R1140 VDD2.n161 VDD2.n160 9.3005
R1141 VDD2.n163 VDD2.n162 9.3005
R1142 VDD2.n105 VDD2.n104 9.3005
R1143 VDD2.n169 VDD2.n168 9.3005
R1144 VDD2.n171 VDD2.n170 9.3005
R1145 VDD2.n186 VDD2.n185 9.3005
R1146 VDD2.n97 VDD2.n96 9.3005
R1147 VDD2.n180 VDD2.n179 9.3005
R1148 VDD2.n178 VDD2.n177 9.3005
R1149 VDD2.n101 VDD2.n100 9.3005
R1150 VDD2.n114 VDD2.n113 9.3005
R1151 VDD2.n147 VDD2.n146 9.3005
R1152 VDD2.n145 VDD2.n144 9.3005
R1153 VDD2.n118 VDD2.n117 9.3005
R1154 VDD2.n139 VDD2.n138 9.3005
R1155 VDD2.n137 VDD2.n136 9.3005
R1156 VDD2.n122 VDD2.n121 9.3005
R1157 VDD2.n131 VDD2.n130 9.3005
R1158 VDD2.n129 VDD2.n128 9.3005
R1159 VDD2.n91 VDD2.n90 9.3005
R1160 VDD2.n2 VDD2.n1 9.3005
R1161 VDD2.n85 VDD2.n84 9.3005
R1162 VDD2.n83 VDD2.n82 9.3005
R1163 VDD2.n6 VDD2.n5 9.3005
R1164 VDD2.n51 VDD2.n50 9.3005
R1165 VDD2.n49 VDD2.n48 9.3005
R1166 VDD2.n22 VDD2.n21 9.3005
R1167 VDD2.n43 VDD2.n42 9.3005
R1168 VDD2.n41 VDD2.n40 9.3005
R1169 VDD2.n26 VDD2.n25 9.3005
R1170 VDD2.n35 VDD2.n34 9.3005
R1171 VDD2.n33 VDD2.n32 9.3005
R1172 VDD2.n18 VDD2.n17 9.3005
R1173 VDD2.n57 VDD2.n56 9.3005
R1174 VDD2.n59 VDD2.n58 9.3005
R1175 VDD2.n14 VDD2.n13 9.3005
R1176 VDD2.n65 VDD2.n64 9.3005
R1177 VDD2.n67 VDD2.n66 9.3005
R1178 VDD2.n10 VDD2.n9 9.3005
R1179 VDD2.n74 VDD2.n73 9.3005
R1180 VDD2.n76 VDD2.n75 9.3005
R1181 VDD2.n156 VDD2.n110 8.92171
R1182 VDD2.n143 VDD2.n118 8.92171
R1183 VDD2.n47 VDD2.n22 8.92171
R1184 VDD2.n60 VDD2.n14 8.92171
R1185 VDD2.n155 VDD2.n112 8.14595
R1186 VDD2.n144 VDD2.n116 8.14595
R1187 VDD2.n48 VDD2.n20 8.14595
R1188 VDD2.n59 VDD2.n16 8.14595
R1189 VDD2.n152 VDD2.n151 7.3702
R1190 VDD2.n148 VDD2.n147 7.3702
R1191 VDD2.n52 VDD2.n51 7.3702
R1192 VDD2.n56 VDD2.n55 7.3702
R1193 VDD2.n151 VDD2.n114 6.59444
R1194 VDD2.n148 VDD2.n114 6.59444
R1195 VDD2.n52 VDD2.n18 6.59444
R1196 VDD2.n55 VDD2.n18 6.59444
R1197 VDD2.n152 VDD2.n112 5.81868
R1198 VDD2.n147 VDD2.n116 5.81868
R1199 VDD2.n51 VDD2.n20 5.81868
R1200 VDD2.n56 VDD2.n16 5.81868
R1201 VDD2.n156 VDD2.n155 5.04292
R1202 VDD2.n144 VDD2.n143 5.04292
R1203 VDD2.n48 VDD2.n47 5.04292
R1204 VDD2.n60 VDD2.n59 5.04292
R1205 VDD2.n187 VDD2.n95 4.26717
R1206 VDD2.n159 VDD2.n110 4.26717
R1207 VDD2.n140 VDD2.n118 4.26717
R1208 VDD2.n44 VDD2.n22 4.26717
R1209 VDD2.n63 VDD2.n14 4.26717
R1210 VDD2.n92 VDD2.n0 4.26717
R1211 VDD2.n129 VDD2.n125 3.70982
R1212 VDD2.n33 VDD2.n29 3.70982
R1213 VDD2.n185 VDD2.n184 3.49141
R1214 VDD2.n160 VDD2.n108 3.49141
R1215 VDD2.n139 VDD2.n120 3.49141
R1216 VDD2.n43 VDD2.n24 3.49141
R1217 VDD2.n64 VDD2.n12 3.49141
R1218 VDD2.n90 VDD2.n89 3.49141
R1219 VDD2.n181 VDD2.n97 2.71565
R1220 VDD2.n164 VDD2.n163 2.71565
R1221 VDD2.n136 VDD2.n135 2.71565
R1222 VDD2.n40 VDD2.n39 2.71565
R1223 VDD2.n68 VDD2.n67 2.71565
R1224 VDD2.n86 VDD2.n2 2.71565
R1225 VDD2 VDD2.n188 2.2311
R1226 VDD2.n180 VDD2.n99 1.93989
R1227 VDD2.n167 VDD2.n105 1.93989
R1228 VDD2.n132 VDD2.n122 1.93989
R1229 VDD2.n36 VDD2.n26 1.93989
R1230 VDD2.n72 VDD2.n10 1.93989
R1231 VDD2.n85 VDD2.n4 1.93989
R1232 VDD2.n189 VDD2.t1 1.9216
R1233 VDD2.n189 VDD2.t2 1.9216
R1234 VDD2.n93 VDD2.t3 1.9216
R1235 VDD2.n93 VDD2.t5 1.9216
R1236 VDD2.n177 VDD2.n176 1.16414
R1237 VDD2.n168 VDD2.n103 1.16414
R1238 VDD2.n131 VDD2.n124 1.16414
R1239 VDD2.n35 VDD2.n28 1.16414
R1240 VDD2.n73 VDD2.n8 1.16414
R1241 VDD2.n82 VDD2.n81 1.16414
R1242 VDD2.n173 VDD2.n101 0.388379
R1243 VDD2.n172 VDD2.n171 0.388379
R1244 VDD2.n128 VDD2.n127 0.388379
R1245 VDD2.n32 VDD2.n31 0.388379
R1246 VDD2.n77 VDD2.n76 0.388379
R1247 VDD2.n78 VDD2.n6 0.388379
R1248 VDD2.n186 VDD2.n96 0.155672
R1249 VDD2.n179 VDD2.n96 0.155672
R1250 VDD2.n179 VDD2.n178 0.155672
R1251 VDD2.n178 VDD2.n100 0.155672
R1252 VDD2.n170 VDD2.n100 0.155672
R1253 VDD2.n170 VDD2.n169 0.155672
R1254 VDD2.n169 VDD2.n104 0.155672
R1255 VDD2.n162 VDD2.n104 0.155672
R1256 VDD2.n162 VDD2.n161 0.155672
R1257 VDD2.n161 VDD2.n109 0.155672
R1258 VDD2.n154 VDD2.n109 0.155672
R1259 VDD2.n154 VDD2.n153 0.155672
R1260 VDD2.n153 VDD2.n113 0.155672
R1261 VDD2.n146 VDD2.n113 0.155672
R1262 VDD2.n146 VDD2.n145 0.155672
R1263 VDD2.n145 VDD2.n117 0.155672
R1264 VDD2.n138 VDD2.n117 0.155672
R1265 VDD2.n138 VDD2.n137 0.155672
R1266 VDD2.n137 VDD2.n121 0.155672
R1267 VDD2.n130 VDD2.n121 0.155672
R1268 VDD2.n130 VDD2.n129 0.155672
R1269 VDD2.n34 VDD2.n33 0.155672
R1270 VDD2.n34 VDD2.n25 0.155672
R1271 VDD2.n41 VDD2.n25 0.155672
R1272 VDD2.n42 VDD2.n41 0.155672
R1273 VDD2.n42 VDD2.n21 0.155672
R1274 VDD2.n49 VDD2.n21 0.155672
R1275 VDD2.n50 VDD2.n49 0.155672
R1276 VDD2.n50 VDD2.n17 0.155672
R1277 VDD2.n57 VDD2.n17 0.155672
R1278 VDD2.n58 VDD2.n57 0.155672
R1279 VDD2.n58 VDD2.n13 0.155672
R1280 VDD2.n65 VDD2.n13 0.155672
R1281 VDD2.n66 VDD2.n65 0.155672
R1282 VDD2.n66 VDD2.n9 0.155672
R1283 VDD2.n74 VDD2.n9 0.155672
R1284 VDD2.n75 VDD2.n74 0.155672
R1285 VDD2.n75 VDD2.n5 0.155672
R1286 VDD2.n83 VDD2.n5 0.155672
R1287 VDD2.n84 VDD2.n83 0.155672
R1288 VDD2.n84 VDD2.n1 0.155672
R1289 VDD2.n91 VDD2.n1 0.155672
R1290 B.n481 B.n480 585
R1291 B.n479 B.n140 585
R1292 B.n478 B.n477 585
R1293 B.n476 B.n141 585
R1294 B.n475 B.n474 585
R1295 B.n473 B.n142 585
R1296 B.n472 B.n471 585
R1297 B.n470 B.n143 585
R1298 B.n469 B.n468 585
R1299 B.n467 B.n144 585
R1300 B.n466 B.n465 585
R1301 B.n464 B.n145 585
R1302 B.n463 B.n462 585
R1303 B.n461 B.n146 585
R1304 B.n460 B.n459 585
R1305 B.n458 B.n147 585
R1306 B.n457 B.n456 585
R1307 B.n455 B.n148 585
R1308 B.n454 B.n453 585
R1309 B.n452 B.n149 585
R1310 B.n451 B.n450 585
R1311 B.n449 B.n150 585
R1312 B.n448 B.n447 585
R1313 B.n446 B.n151 585
R1314 B.n445 B.n444 585
R1315 B.n443 B.n152 585
R1316 B.n442 B.n441 585
R1317 B.n440 B.n153 585
R1318 B.n439 B.n438 585
R1319 B.n437 B.n154 585
R1320 B.n436 B.n435 585
R1321 B.n434 B.n155 585
R1322 B.n433 B.n432 585
R1323 B.n431 B.n156 585
R1324 B.n430 B.n429 585
R1325 B.n428 B.n157 585
R1326 B.n427 B.n426 585
R1327 B.n425 B.n158 585
R1328 B.n424 B.n423 585
R1329 B.n422 B.n159 585
R1330 B.n421 B.n420 585
R1331 B.n419 B.n160 585
R1332 B.n418 B.n417 585
R1333 B.n416 B.n161 585
R1334 B.n415 B.n414 585
R1335 B.n413 B.n162 585
R1336 B.n412 B.n411 585
R1337 B.n410 B.n163 585
R1338 B.n409 B.n408 585
R1339 B.n407 B.n164 585
R1340 B.n406 B.n405 585
R1341 B.n404 B.n165 585
R1342 B.n403 B.n402 585
R1343 B.n401 B.n166 585
R1344 B.n400 B.n399 585
R1345 B.n398 B.n167 585
R1346 B.n397 B.n396 585
R1347 B.n392 B.n168 585
R1348 B.n391 B.n390 585
R1349 B.n389 B.n169 585
R1350 B.n388 B.n387 585
R1351 B.n386 B.n170 585
R1352 B.n385 B.n384 585
R1353 B.n383 B.n171 585
R1354 B.n382 B.n381 585
R1355 B.n380 B.n172 585
R1356 B.n378 B.n377 585
R1357 B.n376 B.n175 585
R1358 B.n375 B.n374 585
R1359 B.n373 B.n176 585
R1360 B.n372 B.n371 585
R1361 B.n370 B.n177 585
R1362 B.n369 B.n368 585
R1363 B.n367 B.n178 585
R1364 B.n366 B.n365 585
R1365 B.n364 B.n179 585
R1366 B.n363 B.n362 585
R1367 B.n361 B.n180 585
R1368 B.n360 B.n359 585
R1369 B.n358 B.n181 585
R1370 B.n357 B.n356 585
R1371 B.n355 B.n182 585
R1372 B.n354 B.n353 585
R1373 B.n352 B.n183 585
R1374 B.n351 B.n350 585
R1375 B.n349 B.n184 585
R1376 B.n348 B.n347 585
R1377 B.n346 B.n185 585
R1378 B.n345 B.n344 585
R1379 B.n343 B.n186 585
R1380 B.n342 B.n341 585
R1381 B.n340 B.n187 585
R1382 B.n339 B.n338 585
R1383 B.n337 B.n188 585
R1384 B.n336 B.n335 585
R1385 B.n334 B.n189 585
R1386 B.n333 B.n332 585
R1387 B.n331 B.n190 585
R1388 B.n330 B.n329 585
R1389 B.n328 B.n191 585
R1390 B.n327 B.n326 585
R1391 B.n325 B.n192 585
R1392 B.n324 B.n323 585
R1393 B.n322 B.n193 585
R1394 B.n321 B.n320 585
R1395 B.n319 B.n194 585
R1396 B.n318 B.n317 585
R1397 B.n316 B.n195 585
R1398 B.n315 B.n314 585
R1399 B.n313 B.n196 585
R1400 B.n312 B.n311 585
R1401 B.n310 B.n197 585
R1402 B.n309 B.n308 585
R1403 B.n307 B.n198 585
R1404 B.n306 B.n305 585
R1405 B.n304 B.n199 585
R1406 B.n303 B.n302 585
R1407 B.n301 B.n200 585
R1408 B.n300 B.n299 585
R1409 B.n298 B.n201 585
R1410 B.n297 B.n296 585
R1411 B.n295 B.n202 585
R1412 B.n482 B.n139 585
R1413 B.n484 B.n483 585
R1414 B.n485 B.n138 585
R1415 B.n487 B.n486 585
R1416 B.n488 B.n137 585
R1417 B.n490 B.n489 585
R1418 B.n491 B.n136 585
R1419 B.n493 B.n492 585
R1420 B.n494 B.n135 585
R1421 B.n496 B.n495 585
R1422 B.n497 B.n134 585
R1423 B.n499 B.n498 585
R1424 B.n500 B.n133 585
R1425 B.n502 B.n501 585
R1426 B.n503 B.n132 585
R1427 B.n505 B.n504 585
R1428 B.n506 B.n131 585
R1429 B.n508 B.n507 585
R1430 B.n509 B.n130 585
R1431 B.n511 B.n510 585
R1432 B.n512 B.n129 585
R1433 B.n514 B.n513 585
R1434 B.n515 B.n128 585
R1435 B.n517 B.n516 585
R1436 B.n518 B.n127 585
R1437 B.n520 B.n519 585
R1438 B.n521 B.n126 585
R1439 B.n523 B.n522 585
R1440 B.n524 B.n125 585
R1441 B.n526 B.n525 585
R1442 B.n527 B.n124 585
R1443 B.n529 B.n528 585
R1444 B.n530 B.n123 585
R1445 B.n532 B.n531 585
R1446 B.n533 B.n122 585
R1447 B.n535 B.n534 585
R1448 B.n536 B.n121 585
R1449 B.n538 B.n537 585
R1450 B.n539 B.n120 585
R1451 B.n541 B.n540 585
R1452 B.n542 B.n119 585
R1453 B.n544 B.n543 585
R1454 B.n545 B.n118 585
R1455 B.n547 B.n546 585
R1456 B.n548 B.n117 585
R1457 B.n550 B.n549 585
R1458 B.n551 B.n116 585
R1459 B.n553 B.n552 585
R1460 B.n554 B.n115 585
R1461 B.n556 B.n555 585
R1462 B.n557 B.n114 585
R1463 B.n559 B.n558 585
R1464 B.n560 B.n113 585
R1465 B.n562 B.n561 585
R1466 B.n563 B.n112 585
R1467 B.n565 B.n564 585
R1468 B.n566 B.n111 585
R1469 B.n568 B.n567 585
R1470 B.n569 B.n110 585
R1471 B.n571 B.n570 585
R1472 B.n572 B.n109 585
R1473 B.n574 B.n573 585
R1474 B.n575 B.n108 585
R1475 B.n577 B.n576 585
R1476 B.n578 B.n107 585
R1477 B.n580 B.n579 585
R1478 B.n581 B.n106 585
R1479 B.n583 B.n582 585
R1480 B.n584 B.n105 585
R1481 B.n586 B.n585 585
R1482 B.n587 B.n104 585
R1483 B.n589 B.n588 585
R1484 B.n590 B.n103 585
R1485 B.n592 B.n591 585
R1486 B.n593 B.n102 585
R1487 B.n595 B.n594 585
R1488 B.n596 B.n101 585
R1489 B.n598 B.n597 585
R1490 B.n599 B.n100 585
R1491 B.n601 B.n600 585
R1492 B.n602 B.n99 585
R1493 B.n604 B.n603 585
R1494 B.n605 B.n98 585
R1495 B.n607 B.n606 585
R1496 B.n608 B.n97 585
R1497 B.n610 B.n609 585
R1498 B.n611 B.n96 585
R1499 B.n613 B.n612 585
R1500 B.n614 B.n95 585
R1501 B.n616 B.n615 585
R1502 B.n617 B.n94 585
R1503 B.n619 B.n618 585
R1504 B.n620 B.n93 585
R1505 B.n622 B.n621 585
R1506 B.n623 B.n92 585
R1507 B.n625 B.n624 585
R1508 B.n809 B.n808 585
R1509 B.n807 B.n26 585
R1510 B.n806 B.n805 585
R1511 B.n804 B.n27 585
R1512 B.n803 B.n802 585
R1513 B.n801 B.n28 585
R1514 B.n800 B.n799 585
R1515 B.n798 B.n29 585
R1516 B.n797 B.n796 585
R1517 B.n795 B.n30 585
R1518 B.n794 B.n793 585
R1519 B.n792 B.n31 585
R1520 B.n791 B.n790 585
R1521 B.n789 B.n32 585
R1522 B.n788 B.n787 585
R1523 B.n786 B.n33 585
R1524 B.n785 B.n784 585
R1525 B.n783 B.n34 585
R1526 B.n782 B.n781 585
R1527 B.n780 B.n35 585
R1528 B.n779 B.n778 585
R1529 B.n777 B.n36 585
R1530 B.n776 B.n775 585
R1531 B.n774 B.n37 585
R1532 B.n773 B.n772 585
R1533 B.n771 B.n38 585
R1534 B.n770 B.n769 585
R1535 B.n768 B.n39 585
R1536 B.n767 B.n766 585
R1537 B.n765 B.n40 585
R1538 B.n764 B.n763 585
R1539 B.n762 B.n41 585
R1540 B.n761 B.n760 585
R1541 B.n759 B.n42 585
R1542 B.n758 B.n757 585
R1543 B.n756 B.n43 585
R1544 B.n755 B.n754 585
R1545 B.n753 B.n44 585
R1546 B.n752 B.n751 585
R1547 B.n750 B.n45 585
R1548 B.n749 B.n748 585
R1549 B.n747 B.n46 585
R1550 B.n746 B.n745 585
R1551 B.n744 B.n47 585
R1552 B.n743 B.n742 585
R1553 B.n741 B.n48 585
R1554 B.n740 B.n739 585
R1555 B.n738 B.n49 585
R1556 B.n737 B.n736 585
R1557 B.n735 B.n50 585
R1558 B.n734 B.n733 585
R1559 B.n732 B.n51 585
R1560 B.n731 B.n730 585
R1561 B.n729 B.n52 585
R1562 B.n728 B.n727 585
R1563 B.n726 B.n53 585
R1564 B.n724 B.n723 585
R1565 B.n722 B.n56 585
R1566 B.n721 B.n720 585
R1567 B.n719 B.n57 585
R1568 B.n718 B.n717 585
R1569 B.n716 B.n58 585
R1570 B.n715 B.n714 585
R1571 B.n713 B.n59 585
R1572 B.n712 B.n711 585
R1573 B.n710 B.n60 585
R1574 B.n709 B.n708 585
R1575 B.n707 B.n61 585
R1576 B.n706 B.n705 585
R1577 B.n704 B.n65 585
R1578 B.n703 B.n702 585
R1579 B.n701 B.n66 585
R1580 B.n700 B.n699 585
R1581 B.n698 B.n67 585
R1582 B.n697 B.n696 585
R1583 B.n695 B.n68 585
R1584 B.n694 B.n693 585
R1585 B.n692 B.n69 585
R1586 B.n691 B.n690 585
R1587 B.n689 B.n70 585
R1588 B.n688 B.n687 585
R1589 B.n686 B.n71 585
R1590 B.n685 B.n684 585
R1591 B.n683 B.n72 585
R1592 B.n682 B.n681 585
R1593 B.n680 B.n73 585
R1594 B.n679 B.n678 585
R1595 B.n677 B.n74 585
R1596 B.n676 B.n675 585
R1597 B.n674 B.n75 585
R1598 B.n673 B.n672 585
R1599 B.n671 B.n76 585
R1600 B.n670 B.n669 585
R1601 B.n668 B.n77 585
R1602 B.n667 B.n666 585
R1603 B.n665 B.n78 585
R1604 B.n664 B.n663 585
R1605 B.n662 B.n79 585
R1606 B.n661 B.n660 585
R1607 B.n659 B.n80 585
R1608 B.n658 B.n657 585
R1609 B.n656 B.n81 585
R1610 B.n655 B.n654 585
R1611 B.n653 B.n82 585
R1612 B.n652 B.n651 585
R1613 B.n650 B.n83 585
R1614 B.n649 B.n648 585
R1615 B.n647 B.n84 585
R1616 B.n646 B.n645 585
R1617 B.n644 B.n85 585
R1618 B.n643 B.n642 585
R1619 B.n641 B.n86 585
R1620 B.n640 B.n639 585
R1621 B.n638 B.n87 585
R1622 B.n637 B.n636 585
R1623 B.n635 B.n88 585
R1624 B.n634 B.n633 585
R1625 B.n632 B.n89 585
R1626 B.n631 B.n630 585
R1627 B.n629 B.n90 585
R1628 B.n628 B.n627 585
R1629 B.n626 B.n91 585
R1630 B.n810 B.n25 585
R1631 B.n812 B.n811 585
R1632 B.n813 B.n24 585
R1633 B.n815 B.n814 585
R1634 B.n816 B.n23 585
R1635 B.n818 B.n817 585
R1636 B.n819 B.n22 585
R1637 B.n821 B.n820 585
R1638 B.n822 B.n21 585
R1639 B.n824 B.n823 585
R1640 B.n825 B.n20 585
R1641 B.n827 B.n826 585
R1642 B.n828 B.n19 585
R1643 B.n830 B.n829 585
R1644 B.n831 B.n18 585
R1645 B.n833 B.n832 585
R1646 B.n834 B.n17 585
R1647 B.n836 B.n835 585
R1648 B.n837 B.n16 585
R1649 B.n839 B.n838 585
R1650 B.n840 B.n15 585
R1651 B.n842 B.n841 585
R1652 B.n843 B.n14 585
R1653 B.n845 B.n844 585
R1654 B.n846 B.n13 585
R1655 B.n848 B.n847 585
R1656 B.n849 B.n12 585
R1657 B.n851 B.n850 585
R1658 B.n852 B.n11 585
R1659 B.n854 B.n853 585
R1660 B.n855 B.n10 585
R1661 B.n857 B.n856 585
R1662 B.n858 B.n9 585
R1663 B.n860 B.n859 585
R1664 B.n861 B.n8 585
R1665 B.n863 B.n862 585
R1666 B.n864 B.n7 585
R1667 B.n866 B.n865 585
R1668 B.n867 B.n6 585
R1669 B.n869 B.n868 585
R1670 B.n870 B.n5 585
R1671 B.n872 B.n871 585
R1672 B.n873 B.n4 585
R1673 B.n875 B.n874 585
R1674 B.n876 B.n3 585
R1675 B.n878 B.n877 585
R1676 B.n879 B.n0 585
R1677 B.n2 B.n1 585
R1678 B.n226 B.n225 585
R1679 B.n228 B.n227 585
R1680 B.n229 B.n224 585
R1681 B.n231 B.n230 585
R1682 B.n232 B.n223 585
R1683 B.n234 B.n233 585
R1684 B.n235 B.n222 585
R1685 B.n237 B.n236 585
R1686 B.n238 B.n221 585
R1687 B.n240 B.n239 585
R1688 B.n241 B.n220 585
R1689 B.n243 B.n242 585
R1690 B.n244 B.n219 585
R1691 B.n246 B.n245 585
R1692 B.n247 B.n218 585
R1693 B.n249 B.n248 585
R1694 B.n250 B.n217 585
R1695 B.n252 B.n251 585
R1696 B.n253 B.n216 585
R1697 B.n255 B.n254 585
R1698 B.n256 B.n215 585
R1699 B.n258 B.n257 585
R1700 B.n259 B.n214 585
R1701 B.n261 B.n260 585
R1702 B.n262 B.n213 585
R1703 B.n264 B.n263 585
R1704 B.n265 B.n212 585
R1705 B.n267 B.n266 585
R1706 B.n268 B.n211 585
R1707 B.n270 B.n269 585
R1708 B.n271 B.n210 585
R1709 B.n273 B.n272 585
R1710 B.n274 B.n209 585
R1711 B.n276 B.n275 585
R1712 B.n277 B.n208 585
R1713 B.n279 B.n278 585
R1714 B.n280 B.n207 585
R1715 B.n282 B.n281 585
R1716 B.n283 B.n206 585
R1717 B.n285 B.n284 585
R1718 B.n286 B.n205 585
R1719 B.n288 B.n287 585
R1720 B.n289 B.n204 585
R1721 B.n291 B.n290 585
R1722 B.n292 B.n203 585
R1723 B.n294 B.n293 585
R1724 B.n393 B.t10 529.532
R1725 B.n62 B.t2 529.532
R1726 B.n173 B.t7 529.532
R1727 B.n54 B.t5 529.532
R1728 B.n293 B.n202 502.111
R1729 B.n482 B.n481 502.111
R1730 B.n626 B.n625 502.111
R1731 B.n808 B.n25 502.111
R1732 B.n394 B.t11 464.368
R1733 B.n63 B.t1 464.368
R1734 B.n174 B.t8 464.368
R1735 B.n55 B.t4 464.368
R1736 B.n173 B.t6 343.193
R1737 B.n393 B.t9 343.193
R1738 B.n62 B.t0 343.193
R1739 B.n54 B.t3 343.193
R1740 B.n881 B.n880 256.663
R1741 B.n880 B.n879 235.042
R1742 B.n880 B.n2 235.042
R1743 B.n297 B.n202 163.367
R1744 B.n298 B.n297 163.367
R1745 B.n299 B.n298 163.367
R1746 B.n299 B.n200 163.367
R1747 B.n303 B.n200 163.367
R1748 B.n304 B.n303 163.367
R1749 B.n305 B.n304 163.367
R1750 B.n305 B.n198 163.367
R1751 B.n309 B.n198 163.367
R1752 B.n310 B.n309 163.367
R1753 B.n311 B.n310 163.367
R1754 B.n311 B.n196 163.367
R1755 B.n315 B.n196 163.367
R1756 B.n316 B.n315 163.367
R1757 B.n317 B.n316 163.367
R1758 B.n317 B.n194 163.367
R1759 B.n321 B.n194 163.367
R1760 B.n322 B.n321 163.367
R1761 B.n323 B.n322 163.367
R1762 B.n323 B.n192 163.367
R1763 B.n327 B.n192 163.367
R1764 B.n328 B.n327 163.367
R1765 B.n329 B.n328 163.367
R1766 B.n329 B.n190 163.367
R1767 B.n333 B.n190 163.367
R1768 B.n334 B.n333 163.367
R1769 B.n335 B.n334 163.367
R1770 B.n335 B.n188 163.367
R1771 B.n339 B.n188 163.367
R1772 B.n340 B.n339 163.367
R1773 B.n341 B.n340 163.367
R1774 B.n341 B.n186 163.367
R1775 B.n345 B.n186 163.367
R1776 B.n346 B.n345 163.367
R1777 B.n347 B.n346 163.367
R1778 B.n347 B.n184 163.367
R1779 B.n351 B.n184 163.367
R1780 B.n352 B.n351 163.367
R1781 B.n353 B.n352 163.367
R1782 B.n353 B.n182 163.367
R1783 B.n357 B.n182 163.367
R1784 B.n358 B.n357 163.367
R1785 B.n359 B.n358 163.367
R1786 B.n359 B.n180 163.367
R1787 B.n363 B.n180 163.367
R1788 B.n364 B.n363 163.367
R1789 B.n365 B.n364 163.367
R1790 B.n365 B.n178 163.367
R1791 B.n369 B.n178 163.367
R1792 B.n370 B.n369 163.367
R1793 B.n371 B.n370 163.367
R1794 B.n371 B.n176 163.367
R1795 B.n375 B.n176 163.367
R1796 B.n376 B.n375 163.367
R1797 B.n377 B.n376 163.367
R1798 B.n377 B.n172 163.367
R1799 B.n382 B.n172 163.367
R1800 B.n383 B.n382 163.367
R1801 B.n384 B.n383 163.367
R1802 B.n384 B.n170 163.367
R1803 B.n388 B.n170 163.367
R1804 B.n389 B.n388 163.367
R1805 B.n390 B.n389 163.367
R1806 B.n390 B.n168 163.367
R1807 B.n397 B.n168 163.367
R1808 B.n398 B.n397 163.367
R1809 B.n399 B.n398 163.367
R1810 B.n399 B.n166 163.367
R1811 B.n403 B.n166 163.367
R1812 B.n404 B.n403 163.367
R1813 B.n405 B.n404 163.367
R1814 B.n405 B.n164 163.367
R1815 B.n409 B.n164 163.367
R1816 B.n410 B.n409 163.367
R1817 B.n411 B.n410 163.367
R1818 B.n411 B.n162 163.367
R1819 B.n415 B.n162 163.367
R1820 B.n416 B.n415 163.367
R1821 B.n417 B.n416 163.367
R1822 B.n417 B.n160 163.367
R1823 B.n421 B.n160 163.367
R1824 B.n422 B.n421 163.367
R1825 B.n423 B.n422 163.367
R1826 B.n423 B.n158 163.367
R1827 B.n427 B.n158 163.367
R1828 B.n428 B.n427 163.367
R1829 B.n429 B.n428 163.367
R1830 B.n429 B.n156 163.367
R1831 B.n433 B.n156 163.367
R1832 B.n434 B.n433 163.367
R1833 B.n435 B.n434 163.367
R1834 B.n435 B.n154 163.367
R1835 B.n439 B.n154 163.367
R1836 B.n440 B.n439 163.367
R1837 B.n441 B.n440 163.367
R1838 B.n441 B.n152 163.367
R1839 B.n445 B.n152 163.367
R1840 B.n446 B.n445 163.367
R1841 B.n447 B.n446 163.367
R1842 B.n447 B.n150 163.367
R1843 B.n451 B.n150 163.367
R1844 B.n452 B.n451 163.367
R1845 B.n453 B.n452 163.367
R1846 B.n453 B.n148 163.367
R1847 B.n457 B.n148 163.367
R1848 B.n458 B.n457 163.367
R1849 B.n459 B.n458 163.367
R1850 B.n459 B.n146 163.367
R1851 B.n463 B.n146 163.367
R1852 B.n464 B.n463 163.367
R1853 B.n465 B.n464 163.367
R1854 B.n465 B.n144 163.367
R1855 B.n469 B.n144 163.367
R1856 B.n470 B.n469 163.367
R1857 B.n471 B.n470 163.367
R1858 B.n471 B.n142 163.367
R1859 B.n475 B.n142 163.367
R1860 B.n476 B.n475 163.367
R1861 B.n477 B.n476 163.367
R1862 B.n477 B.n140 163.367
R1863 B.n481 B.n140 163.367
R1864 B.n625 B.n92 163.367
R1865 B.n621 B.n92 163.367
R1866 B.n621 B.n620 163.367
R1867 B.n620 B.n619 163.367
R1868 B.n619 B.n94 163.367
R1869 B.n615 B.n94 163.367
R1870 B.n615 B.n614 163.367
R1871 B.n614 B.n613 163.367
R1872 B.n613 B.n96 163.367
R1873 B.n609 B.n96 163.367
R1874 B.n609 B.n608 163.367
R1875 B.n608 B.n607 163.367
R1876 B.n607 B.n98 163.367
R1877 B.n603 B.n98 163.367
R1878 B.n603 B.n602 163.367
R1879 B.n602 B.n601 163.367
R1880 B.n601 B.n100 163.367
R1881 B.n597 B.n100 163.367
R1882 B.n597 B.n596 163.367
R1883 B.n596 B.n595 163.367
R1884 B.n595 B.n102 163.367
R1885 B.n591 B.n102 163.367
R1886 B.n591 B.n590 163.367
R1887 B.n590 B.n589 163.367
R1888 B.n589 B.n104 163.367
R1889 B.n585 B.n104 163.367
R1890 B.n585 B.n584 163.367
R1891 B.n584 B.n583 163.367
R1892 B.n583 B.n106 163.367
R1893 B.n579 B.n106 163.367
R1894 B.n579 B.n578 163.367
R1895 B.n578 B.n577 163.367
R1896 B.n577 B.n108 163.367
R1897 B.n573 B.n108 163.367
R1898 B.n573 B.n572 163.367
R1899 B.n572 B.n571 163.367
R1900 B.n571 B.n110 163.367
R1901 B.n567 B.n110 163.367
R1902 B.n567 B.n566 163.367
R1903 B.n566 B.n565 163.367
R1904 B.n565 B.n112 163.367
R1905 B.n561 B.n112 163.367
R1906 B.n561 B.n560 163.367
R1907 B.n560 B.n559 163.367
R1908 B.n559 B.n114 163.367
R1909 B.n555 B.n114 163.367
R1910 B.n555 B.n554 163.367
R1911 B.n554 B.n553 163.367
R1912 B.n553 B.n116 163.367
R1913 B.n549 B.n116 163.367
R1914 B.n549 B.n548 163.367
R1915 B.n548 B.n547 163.367
R1916 B.n547 B.n118 163.367
R1917 B.n543 B.n118 163.367
R1918 B.n543 B.n542 163.367
R1919 B.n542 B.n541 163.367
R1920 B.n541 B.n120 163.367
R1921 B.n537 B.n120 163.367
R1922 B.n537 B.n536 163.367
R1923 B.n536 B.n535 163.367
R1924 B.n535 B.n122 163.367
R1925 B.n531 B.n122 163.367
R1926 B.n531 B.n530 163.367
R1927 B.n530 B.n529 163.367
R1928 B.n529 B.n124 163.367
R1929 B.n525 B.n124 163.367
R1930 B.n525 B.n524 163.367
R1931 B.n524 B.n523 163.367
R1932 B.n523 B.n126 163.367
R1933 B.n519 B.n126 163.367
R1934 B.n519 B.n518 163.367
R1935 B.n518 B.n517 163.367
R1936 B.n517 B.n128 163.367
R1937 B.n513 B.n128 163.367
R1938 B.n513 B.n512 163.367
R1939 B.n512 B.n511 163.367
R1940 B.n511 B.n130 163.367
R1941 B.n507 B.n130 163.367
R1942 B.n507 B.n506 163.367
R1943 B.n506 B.n505 163.367
R1944 B.n505 B.n132 163.367
R1945 B.n501 B.n132 163.367
R1946 B.n501 B.n500 163.367
R1947 B.n500 B.n499 163.367
R1948 B.n499 B.n134 163.367
R1949 B.n495 B.n134 163.367
R1950 B.n495 B.n494 163.367
R1951 B.n494 B.n493 163.367
R1952 B.n493 B.n136 163.367
R1953 B.n489 B.n136 163.367
R1954 B.n489 B.n488 163.367
R1955 B.n488 B.n487 163.367
R1956 B.n487 B.n138 163.367
R1957 B.n483 B.n138 163.367
R1958 B.n483 B.n482 163.367
R1959 B.n808 B.n807 163.367
R1960 B.n807 B.n806 163.367
R1961 B.n806 B.n27 163.367
R1962 B.n802 B.n27 163.367
R1963 B.n802 B.n801 163.367
R1964 B.n801 B.n800 163.367
R1965 B.n800 B.n29 163.367
R1966 B.n796 B.n29 163.367
R1967 B.n796 B.n795 163.367
R1968 B.n795 B.n794 163.367
R1969 B.n794 B.n31 163.367
R1970 B.n790 B.n31 163.367
R1971 B.n790 B.n789 163.367
R1972 B.n789 B.n788 163.367
R1973 B.n788 B.n33 163.367
R1974 B.n784 B.n33 163.367
R1975 B.n784 B.n783 163.367
R1976 B.n783 B.n782 163.367
R1977 B.n782 B.n35 163.367
R1978 B.n778 B.n35 163.367
R1979 B.n778 B.n777 163.367
R1980 B.n777 B.n776 163.367
R1981 B.n776 B.n37 163.367
R1982 B.n772 B.n37 163.367
R1983 B.n772 B.n771 163.367
R1984 B.n771 B.n770 163.367
R1985 B.n770 B.n39 163.367
R1986 B.n766 B.n39 163.367
R1987 B.n766 B.n765 163.367
R1988 B.n765 B.n764 163.367
R1989 B.n764 B.n41 163.367
R1990 B.n760 B.n41 163.367
R1991 B.n760 B.n759 163.367
R1992 B.n759 B.n758 163.367
R1993 B.n758 B.n43 163.367
R1994 B.n754 B.n43 163.367
R1995 B.n754 B.n753 163.367
R1996 B.n753 B.n752 163.367
R1997 B.n752 B.n45 163.367
R1998 B.n748 B.n45 163.367
R1999 B.n748 B.n747 163.367
R2000 B.n747 B.n746 163.367
R2001 B.n746 B.n47 163.367
R2002 B.n742 B.n47 163.367
R2003 B.n742 B.n741 163.367
R2004 B.n741 B.n740 163.367
R2005 B.n740 B.n49 163.367
R2006 B.n736 B.n49 163.367
R2007 B.n736 B.n735 163.367
R2008 B.n735 B.n734 163.367
R2009 B.n734 B.n51 163.367
R2010 B.n730 B.n51 163.367
R2011 B.n730 B.n729 163.367
R2012 B.n729 B.n728 163.367
R2013 B.n728 B.n53 163.367
R2014 B.n723 B.n53 163.367
R2015 B.n723 B.n722 163.367
R2016 B.n722 B.n721 163.367
R2017 B.n721 B.n57 163.367
R2018 B.n717 B.n57 163.367
R2019 B.n717 B.n716 163.367
R2020 B.n716 B.n715 163.367
R2021 B.n715 B.n59 163.367
R2022 B.n711 B.n59 163.367
R2023 B.n711 B.n710 163.367
R2024 B.n710 B.n709 163.367
R2025 B.n709 B.n61 163.367
R2026 B.n705 B.n61 163.367
R2027 B.n705 B.n704 163.367
R2028 B.n704 B.n703 163.367
R2029 B.n703 B.n66 163.367
R2030 B.n699 B.n66 163.367
R2031 B.n699 B.n698 163.367
R2032 B.n698 B.n697 163.367
R2033 B.n697 B.n68 163.367
R2034 B.n693 B.n68 163.367
R2035 B.n693 B.n692 163.367
R2036 B.n692 B.n691 163.367
R2037 B.n691 B.n70 163.367
R2038 B.n687 B.n70 163.367
R2039 B.n687 B.n686 163.367
R2040 B.n686 B.n685 163.367
R2041 B.n685 B.n72 163.367
R2042 B.n681 B.n72 163.367
R2043 B.n681 B.n680 163.367
R2044 B.n680 B.n679 163.367
R2045 B.n679 B.n74 163.367
R2046 B.n675 B.n74 163.367
R2047 B.n675 B.n674 163.367
R2048 B.n674 B.n673 163.367
R2049 B.n673 B.n76 163.367
R2050 B.n669 B.n76 163.367
R2051 B.n669 B.n668 163.367
R2052 B.n668 B.n667 163.367
R2053 B.n667 B.n78 163.367
R2054 B.n663 B.n78 163.367
R2055 B.n663 B.n662 163.367
R2056 B.n662 B.n661 163.367
R2057 B.n661 B.n80 163.367
R2058 B.n657 B.n80 163.367
R2059 B.n657 B.n656 163.367
R2060 B.n656 B.n655 163.367
R2061 B.n655 B.n82 163.367
R2062 B.n651 B.n82 163.367
R2063 B.n651 B.n650 163.367
R2064 B.n650 B.n649 163.367
R2065 B.n649 B.n84 163.367
R2066 B.n645 B.n84 163.367
R2067 B.n645 B.n644 163.367
R2068 B.n644 B.n643 163.367
R2069 B.n643 B.n86 163.367
R2070 B.n639 B.n86 163.367
R2071 B.n639 B.n638 163.367
R2072 B.n638 B.n637 163.367
R2073 B.n637 B.n88 163.367
R2074 B.n633 B.n88 163.367
R2075 B.n633 B.n632 163.367
R2076 B.n632 B.n631 163.367
R2077 B.n631 B.n90 163.367
R2078 B.n627 B.n90 163.367
R2079 B.n627 B.n626 163.367
R2080 B.n812 B.n25 163.367
R2081 B.n813 B.n812 163.367
R2082 B.n814 B.n813 163.367
R2083 B.n814 B.n23 163.367
R2084 B.n818 B.n23 163.367
R2085 B.n819 B.n818 163.367
R2086 B.n820 B.n819 163.367
R2087 B.n820 B.n21 163.367
R2088 B.n824 B.n21 163.367
R2089 B.n825 B.n824 163.367
R2090 B.n826 B.n825 163.367
R2091 B.n826 B.n19 163.367
R2092 B.n830 B.n19 163.367
R2093 B.n831 B.n830 163.367
R2094 B.n832 B.n831 163.367
R2095 B.n832 B.n17 163.367
R2096 B.n836 B.n17 163.367
R2097 B.n837 B.n836 163.367
R2098 B.n838 B.n837 163.367
R2099 B.n838 B.n15 163.367
R2100 B.n842 B.n15 163.367
R2101 B.n843 B.n842 163.367
R2102 B.n844 B.n843 163.367
R2103 B.n844 B.n13 163.367
R2104 B.n848 B.n13 163.367
R2105 B.n849 B.n848 163.367
R2106 B.n850 B.n849 163.367
R2107 B.n850 B.n11 163.367
R2108 B.n854 B.n11 163.367
R2109 B.n855 B.n854 163.367
R2110 B.n856 B.n855 163.367
R2111 B.n856 B.n9 163.367
R2112 B.n860 B.n9 163.367
R2113 B.n861 B.n860 163.367
R2114 B.n862 B.n861 163.367
R2115 B.n862 B.n7 163.367
R2116 B.n866 B.n7 163.367
R2117 B.n867 B.n866 163.367
R2118 B.n868 B.n867 163.367
R2119 B.n868 B.n5 163.367
R2120 B.n872 B.n5 163.367
R2121 B.n873 B.n872 163.367
R2122 B.n874 B.n873 163.367
R2123 B.n874 B.n3 163.367
R2124 B.n878 B.n3 163.367
R2125 B.n879 B.n878 163.367
R2126 B.n226 B.n2 163.367
R2127 B.n227 B.n226 163.367
R2128 B.n227 B.n224 163.367
R2129 B.n231 B.n224 163.367
R2130 B.n232 B.n231 163.367
R2131 B.n233 B.n232 163.367
R2132 B.n233 B.n222 163.367
R2133 B.n237 B.n222 163.367
R2134 B.n238 B.n237 163.367
R2135 B.n239 B.n238 163.367
R2136 B.n239 B.n220 163.367
R2137 B.n243 B.n220 163.367
R2138 B.n244 B.n243 163.367
R2139 B.n245 B.n244 163.367
R2140 B.n245 B.n218 163.367
R2141 B.n249 B.n218 163.367
R2142 B.n250 B.n249 163.367
R2143 B.n251 B.n250 163.367
R2144 B.n251 B.n216 163.367
R2145 B.n255 B.n216 163.367
R2146 B.n256 B.n255 163.367
R2147 B.n257 B.n256 163.367
R2148 B.n257 B.n214 163.367
R2149 B.n261 B.n214 163.367
R2150 B.n262 B.n261 163.367
R2151 B.n263 B.n262 163.367
R2152 B.n263 B.n212 163.367
R2153 B.n267 B.n212 163.367
R2154 B.n268 B.n267 163.367
R2155 B.n269 B.n268 163.367
R2156 B.n269 B.n210 163.367
R2157 B.n273 B.n210 163.367
R2158 B.n274 B.n273 163.367
R2159 B.n275 B.n274 163.367
R2160 B.n275 B.n208 163.367
R2161 B.n279 B.n208 163.367
R2162 B.n280 B.n279 163.367
R2163 B.n281 B.n280 163.367
R2164 B.n281 B.n206 163.367
R2165 B.n285 B.n206 163.367
R2166 B.n286 B.n285 163.367
R2167 B.n287 B.n286 163.367
R2168 B.n287 B.n204 163.367
R2169 B.n291 B.n204 163.367
R2170 B.n292 B.n291 163.367
R2171 B.n293 B.n292 163.367
R2172 B.n174 B.n173 65.1641
R2173 B.n394 B.n393 65.1641
R2174 B.n63 B.n62 65.1641
R2175 B.n55 B.n54 65.1641
R2176 B.n379 B.n174 59.5399
R2177 B.n395 B.n394 59.5399
R2178 B.n64 B.n63 59.5399
R2179 B.n725 B.n55 59.5399
R2180 B.n810 B.n809 32.6249
R2181 B.n624 B.n91 32.6249
R2182 B.n480 B.n139 32.6249
R2183 B.n295 B.n294 32.6249
R2184 B B.n881 18.0485
R2185 B.n811 B.n810 10.6151
R2186 B.n811 B.n24 10.6151
R2187 B.n815 B.n24 10.6151
R2188 B.n816 B.n815 10.6151
R2189 B.n817 B.n816 10.6151
R2190 B.n817 B.n22 10.6151
R2191 B.n821 B.n22 10.6151
R2192 B.n822 B.n821 10.6151
R2193 B.n823 B.n822 10.6151
R2194 B.n823 B.n20 10.6151
R2195 B.n827 B.n20 10.6151
R2196 B.n828 B.n827 10.6151
R2197 B.n829 B.n828 10.6151
R2198 B.n829 B.n18 10.6151
R2199 B.n833 B.n18 10.6151
R2200 B.n834 B.n833 10.6151
R2201 B.n835 B.n834 10.6151
R2202 B.n835 B.n16 10.6151
R2203 B.n839 B.n16 10.6151
R2204 B.n840 B.n839 10.6151
R2205 B.n841 B.n840 10.6151
R2206 B.n841 B.n14 10.6151
R2207 B.n845 B.n14 10.6151
R2208 B.n846 B.n845 10.6151
R2209 B.n847 B.n846 10.6151
R2210 B.n847 B.n12 10.6151
R2211 B.n851 B.n12 10.6151
R2212 B.n852 B.n851 10.6151
R2213 B.n853 B.n852 10.6151
R2214 B.n853 B.n10 10.6151
R2215 B.n857 B.n10 10.6151
R2216 B.n858 B.n857 10.6151
R2217 B.n859 B.n858 10.6151
R2218 B.n859 B.n8 10.6151
R2219 B.n863 B.n8 10.6151
R2220 B.n864 B.n863 10.6151
R2221 B.n865 B.n864 10.6151
R2222 B.n865 B.n6 10.6151
R2223 B.n869 B.n6 10.6151
R2224 B.n870 B.n869 10.6151
R2225 B.n871 B.n870 10.6151
R2226 B.n871 B.n4 10.6151
R2227 B.n875 B.n4 10.6151
R2228 B.n876 B.n875 10.6151
R2229 B.n877 B.n876 10.6151
R2230 B.n877 B.n0 10.6151
R2231 B.n809 B.n26 10.6151
R2232 B.n805 B.n26 10.6151
R2233 B.n805 B.n804 10.6151
R2234 B.n804 B.n803 10.6151
R2235 B.n803 B.n28 10.6151
R2236 B.n799 B.n28 10.6151
R2237 B.n799 B.n798 10.6151
R2238 B.n798 B.n797 10.6151
R2239 B.n797 B.n30 10.6151
R2240 B.n793 B.n30 10.6151
R2241 B.n793 B.n792 10.6151
R2242 B.n792 B.n791 10.6151
R2243 B.n791 B.n32 10.6151
R2244 B.n787 B.n32 10.6151
R2245 B.n787 B.n786 10.6151
R2246 B.n786 B.n785 10.6151
R2247 B.n785 B.n34 10.6151
R2248 B.n781 B.n34 10.6151
R2249 B.n781 B.n780 10.6151
R2250 B.n780 B.n779 10.6151
R2251 B.n779 B.n36 10.6151
R2252 B.n775 B.n36 10.6151
R2253 B.n775 B.n774 10.6151
R2254 B.n774 B.n773 10.6151
R2255 B.n773 B.n38 10.6151
R2256 B.n769 B.n38 10.6151
R2257 B.n769 B.n768 10.6151
R2258 B.n768 B.n767 10.6151
R2259 B.n767 B.n40 10.6151
R2260 B.n763 B.n40 10.6151
R2261 B.n763 B.n762 10.6151
R2262 B.n762 B.n761 10.6151
R2263 B.n761 B.n42 10.6151
R2264 B.n757 B.n42 10.6151
R2265 B.n757 B.n756 10.6151
R2266 B.n756 B.n755 10.6151
R2267 B.n755 B.n44 10.6151
R2268 B.n751 B.n44 10.6151
R2269 B.n751 B.n750 10.6151
R2270 B.n750 B.n749 10.6151
R2271 B.n749 B.n46 10.6151
R2272 B.n745 B.n46 10.6151
R2273 B.n745 B.n744 10.6151
R2274 B.n744 B.n743 10.6151
R2275 B.n743 B.n48 10.6151
R2276 B.n739 B.n48 10.6151
R2277 B.n739 B.n738 10.6151
R2278 B.n738 B.n737 10.6151
R2279 B.n737 B.n50 10.6151
R2280 B.n733 B.n50 10.6151
R2281 B.n733 B.n732 10.6151
R2282 B.n732 B.n731 10.6151
R2283 B.n731 B.n52 10.6151
R2284 B.n727 B.n52 10.6151
R2285 B.n727 B.n726 10.6151
R2286 B.n724 B.n56 10.6151
R2287 B.n720 B.n56 10.6151
R2288 B.n720 B.n719 10.6151
R2289 B.n719 B.n718 10.6151
R2290 B.n718 B.n58 10.6151
R2291 B.n714 B.n58 10.6151
R2292 B.n714 B.n713 10.6151
R2293 B.n713 B.n712 10.6151
R2294 B.n712 B.n60 10.6151
R2295 B.n708 B.n707 10.6151
R2296 B.n707 B.n706 10.6151
R2297 B.n706 B.n65 10.6151
R2298 B.n702 B.n65 10.6151
R2299 B.n702 B.n701 10.6151
R2300 B.n701 B.n700 10.6151
R2301 B.n700 B.n67 10.6151
R2302 B.n696 B.n67 10.6151
R2303 B.n696 B.n695 10.6151
R2304 B.n695 B.n694 10.6151
R2305 B.n694 B.n69 10.6151
R2306 B.n690 B.n69 10.6151
R2307 B.n690 B.n689 10.6151
R2308 B.n689 B.n688 10.6151
R2309 B.n688 B.n71 10.6151
R2310 B.n684 B.n71 10.6151
R2311 B.n684 B.n683 10.6151
R2312 B.n683 B.n682 10.6151
R2313 B.n682 B.n73 10.6151
R2314 B.n678 B.n73 10.6151
R2315 B.n678 B.n677 10.6151
R2316 B.n677 B.n676 10.6151
R2317 B.n676 B.n75 10.6151
R2318 B.n672 B.n75 10.6151
R2319 B.n672 B.n671 10.6151
R2320 B.n671 B.n670 10.6151
R2321 B.n670 B.n77 10.6151
R2322 B.n666 B.n77 10.6151
R2323 B.n666 B.n665 10.6151
R2324 B.n665 B.n664 10.6151
R2325 B.n664 B.n79 10.6151
R2326 B.n660 B.n79 10.6151
R2327 B.n660 B.n659 10.6151
R2328 B.n659 B.n658 10.6151
R2329 B.n658 B.n81 10.6151
R2330 B.n654 B.n81 10.6151
R2331 B.n654 B.n653 10.6151
R2332 B.n653 B.n652 10.6151
R2333 B.n652 B.n83 10.6151
R2334 B.n648 B.n83 10.6151
R2335 B.n648 B.n647 10.6151
R2336 B.n647 B.n646 10.6151
R2337 B.n646 B.n85 10.6151
R2338 B.n642 B.n85 10.6151
R2339 B.n642 B.n641 10.6151
R2340 B.n641 B.n640 10.6151
R2341 B.n640 B.n87 10.6151
R2342 B.n636 B.n87 10.6151
R2343 B.n636 B.n635 10.6151
R2344 B.n635 B.n634 10.6151
R2345 B.n634 B.n89 10.6151
R2346 B.n630 B.n89 10.6151
R2347 B.n630 B.n629 10.6151
R2348 B.n629 B.n628 10.6151
R2349 B.n628 B.n91 10.6151
R2350 B.n624 B.n623 10.6151
R2351 B.n623 B.n622 10.6151
R2352 B.n622 B.n93 10.6151
R2353 B.n618 B.n93 10.6151
R2354 B.n618 B.n617 10.6151
R2355 B.n617 B.n616 10.6151
R2356 B.n616 B.n95 10.6151
R2357 B.n612 B.n95 10.6151
R2358 B.n612 B.n611 10.6151
R2359 B.n611 B.n610 10.6151
R2360 B.n610 B.n97 10.6151
R2361 B.n606 B.n97 10.6151
R2362 B.n606 B.n605 10.6151
R2363 B.n605 B.n604 10.6151
R2364 B.n604 B.n99 10.6151
R2365 B.n600 B.n99 10.6151
R2366 B.n600 B.n599 10.6151
R2367 B.n599 B.n598 10.6151
R2368 B.n598 B.n101 10.6151
R2369 B.n594 B.n101 10.6151
R2370 B.n594 B.n593 10.6151
R2371 B.n593 B.n592 10.6151
R2372 B.n592 B.n103 10.6151
R2373 B.n588 B.n103 10.6151
R2374 B.n588 B.n587 10.6151
R2375 B.n587 B.n586 10.6151
R2376 B.n586 B.n105 10.6151
R2377 B.n582 B.n105 10.6151
R2378 B.n582 B.n581 10.6151
R2379 B.n581 B.n580 10.6151
R2380 B.n580 B.n107 10.6151
R2381 B.n576 B.n107 10.6151
R2382 B.n576 B.n575 10.6151
R2383 B.n575 B.n574 10.6151
R2384 B.n574 B.n109 10.6151
R2385 B.n570 B.n109 10.6151
R2386 B.n570 B.n569 10.6151
R2387 B.n569 B.n568 10.6151
R2388 B.n568 B.n111 10.6151
R2389 B.n564 B.n111 10.6151
R2390 B.n564 B.n563 10.6151
R2391 B.n563 B.n562 10.6151
R2392 B.n562 B.n113 10.6151
R2393 B.n558 B.n113 10.6151
R2394 B.n558 B.n557 10.6151
R2395 B.n557 B.n556 10.6151
R2396 B.n556 B.n115 10.6151
R2397 B.n552 B.n115 10.6151
R2398 B.n552 B.n551 10.6151
R2399 B.n551 B.n550 10.6151
R2400 B.n550 B.n117 10.6151
R2401 B.n546 B.n117 10.6151
R2402 B.n546 B.n545 10.6151
R2403 B.n545 B.n544 10.6151
R2404 B.n544 B.n119 10.6151
R2405 B.n540 B.n119 10.6151
R2406 B.n540 B.n539 10.6151
R2407 B.n539 B.n538 10.6151
R2408 B.n538 B.n121 10.6151
R2409 B.n534 B.n121 10.6151
R2410 B.n534 B.n533 10.6151
R2411 B.n533 B.n532 10.6151
R2412 B.n532 B.n123 10.6151
R2413 B.n528 B.n123 10.6151
R2414 B.n528 B.n527 10.6151
R2415 B.n527 B.n526 10.6151
R2416 B.n526 B.n125 10.6151
R2417 B.n522 B.n125 10.6151
R2418 B.n522 B.n521 10.6151
R2419 B.n521 B.n520 10.6151
R2420 B.n520 B.n127 10.6151
R2421 B.n516 B.n127 10.6151
R2422 B.n516 B.n515 10.6151
R2423 B.n515 B.n514 10.6151
R2424 B.n514 B.n129 10.6151
R2425 B.n510 B.n129 10.6151
R2426 B.n510 B.n509 10.6151
R2427 B.n509 B.n508 10.6151
R2428 B.n508 B.n131 10.6151
R2429 B.n504 B.n131 10.6151
R2430 B.n504 B.n503 10.6151
R2431 B.n503 B.n502 10.6151
R2432 B.n502 B.n133 10.6151
R2433 B.n498 B.n133 10.6151
R2434 B.n498 B.n497 10.6151
R2435 B.n497 B.n496 10.6151
R2436 B.n496 B.n135 10.6151
R2437 B.n492 B.n135 10.6151
R2438 B.n492 B.n491 10.6151
R2439 B.n491 B.n490 10.6151
R2440 B.n490 B.n137 10.6151
R2441 B.n486 B.n137 10.6151
R2442 B.n486 B.n485 10.6151
R2443 B.n485 B.n484 10.6151
R2444 B.n484 B.n139 10.6151
R2445 B.n225 B.n1 10.6151
R2446 B.n228 B.n225 10.6151
R2447 B.n229 B.n228 10.6151
R2448 B.n230 B.n229 10.6151
R2449 B.n230 B.n223 10.6151
R2450 B.n234 B.n223 10.6151
R2451 B.n235 B.n234 10.6151
R2452 B.n236 B.n235 10.6151
R2453 B.n236 B.n221 10.6151
R2454 B.n240 B.n221 10.6151
R2455 B.n241 B.n240 10.6151
R2456 B.n242 B.n241 10.6151
R2457 B.n242 B.n219 10.6151
R2458 B.n246 B.n219 10.6151
R2459 B.n247 B.n246 10.6151
R2460 B.n248 B.n247 10.6151
R2461 B.n248 B.n217 10.6151
R2462 B.n252 B.n217 10.6151
R2463 B.n253 B.n252 10.6151
R2464 B.n254 B.n253 10.6151
R2465 B.n254 B.n215 10.6151
R2466 B.n258 B.n215 10.6151
R2467 B.n259 B.n258 10.6151
R2468 B.n260 B.n259 10.6151
R2469 B.n260 B.n213 10.6151
R2470 B.n264 B.n213 10.6151
R2471 B.n265 B.n264 10.6151
R2472 B.n266 B.n265 10.6151
R2473 B.n266 B.n211 10.6151
R2474 B.n270 B.n211 10.6151
R2475 B.n271 B.n270 10.6151
R2476 B.n272 B.n271 10.6151
R2477 B.n272 B.n209 10.6151
R2478 B.n276 B.n209 10.6151
R2479 B.n277 B.n276 10.6151
R2480 B.n278 B.n277 10.6151
R2481 B.n278 B.n207 10.6151
R2482 B.n282 B.n207 10.6151
R2483 B.n283 B.n282 10.6151
R2484 B.n284 B.n283 10.6151
R2485 B.n284 B.n205 10.6151
R2486 B.n288 B.n205 10.6151
R2487 B.n289 B.n288 10.6151
R2488 B.n290 B.n289 10.6151
R2489 B.n290 B.n203 10.6151
R2490 B.n294 B.n203 10.6151
R2491 B.n296 B.n295 10.6151
R2492 B.n296 B.n201 10.6151
R2493 B.n300 B.n201 10.6151
R2494 B.n301 B.n300 10.6151
R2495 B.n302 B.n301 10.6151
R2496 B.n302 B.n199 10.6151
R2497 B.n306 B.n199 10.6151
R2498 B.n307 B.n306 10.6151
R2499 B.n308 B.n307 10.6151
R2500 B.n308 B.n197 10.6151
R2501 B.n312 B.n197 10.6151
R2502 B.n313 B.n312 10.6151
R2503 B.n314 B.n313 10.6151
R2504 B.n314 B.n195 10.6151
R2505 B.n318 B.n195 10.6151
R2506 B.n319 B.n318 10.6151
R2507 B.n320 B.n319 10.6151
R2508 B.n320 B.n193 10.6151
R2509 B.n324 B.n193 10.6151
R2510 B.n325 B.n324 10.6151
R2511 B.n326 B.n325 10.6151
R2512 B.n326 B.n191 10.6151
R2513 B.n330 B.n191 10.6151
R2514 B.n331 B.n330 10.6151
R2515 B.n332 B.n331 10.6151
R2516 B.n332 B.n189 10.6151
R2517 B.n336 B.n189 10.6151
R2518 B.n337 B.n336 10.6151
R2519 B.n338 B.n337 10.6151
R2520 B.n338 B.n187 10.6151
R2521 B.n342 B.n187 10.6151
R2522 B.n343 B.n342 10.6151
R2523 B.n344 B.n343 10.6151
R2524 B.n344 B.n185 10.6151
R2525 B.n348 B.n185 10.6151
R2526 B.n349 B.n348 10.6151
R2527 B.n350 B.n349 10.6151
R2528 B.n350 B.n183 10.6151
R2529 B.n354 B.n183 10.6151
R2530 B.n355 B.n354 10.6151
R2531 B.n356 B.n355 10.6151
R2532 B.n356 B.n181 10.6151
R2533 B.n360 B.n181 10.6151
R2534 B.n361 B.n360 10.6151
R2535 B.n362 B.n361 10.6151
R2536 B.n362 B.n179 10.6151
R2537 B.n366 B.n179 10.6151
R2538 B.n367 B.n366 10.6151
R2539 B.n368 B.n367 10.6151
R2540 B.n368 B.n177 10.6151
R2541 B.n372 B.n177 10.6151
R2542 B.n373 B.n372 10.6151
R2543 B.n374 B.n373 10.6151
R2544 B.n374 B.n175 10.6151
R2545 B.n378 B.n175 10.6151
R2546 B.n381 B.n380 10.6151
R2547 B.n381 B.n171 10.6151
R2548 B.n385 B.n171 10.6151
R2549 B.n386 B.n385 10.6151
R2550 B.n387 B.n386 10.6151
R2551 B.n387 B.n169 10.6151
R2552 B.n391 B.n169 10.6151
R2553 B.n392 B.n391 10.6151
R2554 B.n396 B.n392 10.6151
R2555 B.n400 B.n167 10.6151
R2556 B.n401 B.n400 10.6151
R2557 B.n402 B.n401 10.6151
R2558 B.n402 B.n165 10.6151
R2559 B.n406 B.n165 10.6151
R2560 B.n407 B.n406 10.6151
R2561 B.n408 B.n407 10.6151
R2562 B.n408 B.n163 10.6151
R2563 B.n412 B.n163 10.6151
R2564 B.n413 B.n412 10.6151
R2565 B.n414 B.n413 10.6151
R2566 B.n414 B.n161 10.6151
R2567 B.n418 B.n161 10.6151
R2568 B.n419 B.n418 10.6151
R2569 B.n420 B.n419 10.6151
R2570 B.n420 B.n159 10.6151
R2571 B.n424 B.n159 10.6151
R2572 B.n425 B.n424 10.6151
R2573 B.n426 B.n425 10.6151
R2574 B.n426 B.n157 10.6151
R2575 B.n430 B.n157 10.6151
R2576 B.n431 B.n430 10.6151
R2577 B.n432 B.n431 10.6151
R2578 B.n432 B.n155 10.6151
R2579 B.n436 B.n155 10.6151
R2580 B.n437 B.n436 10.6151
R2581 B.n438 B.n437 10.6151
R2582 B.n438 B.n153 10.6151
R2583 B.n442 B.n153 10.6151
R2584 B.n443 B.n442 10.6151
R2585 B.n444 B.n443 10.6151
R2586 B.n444 B.n151 10.6151
R2587 B.n448 B.n151 10.6151
R2588 B.n449 B.n448 10.6151
R2589 B.n450 B.n449 10.6151
R2590 B.n450 B.n149 10.6151
R2591 B.n454 B.n149 10.6151
R2592 B.n455 B.n454 10.6151
R2593 B.n456 B.n455 10.6151
R2594 B.n456 B.n147 10.6151
R2595 B.n460 B.n147 10.6151
R2596 B.n461 B.n460 10.6151
R2597 B.n462 B.n461 10.6151
R2598 B.n462 B.n145 10.6151
R2599 B.n466 B.n145 10.6151
R2600 B.n467 B.n466 10.6151
R2601 B.n468 B.n467 10.6151
R2602 B.n468 B.n143 10.6151
R2603 B.n472 B.n143 10.6151
R2604 B.n473 B.n472 10.6151
R2605 B.n474 B.n473 10.6151
R2606 B.n474 B.n141 10.6151
R2607 B.n478 B.n141 10.6151
R2608 B.n479 B.n478 10.6151
R2609 B.n480 B.n479 10.6151
R2610 B.n726 B.n725 9.36635
R2611 B.n708 B.n64 9.36635
R2612 B.n379 B.n378 9.36635
R2613 B.n395 B.n167 9.36635
R2614 B.n881 B.n0 8.11757
R2615 B.n881 B.n1 8.11757
R2616 B.n725 B.n724 1.24928
R2617 B.n64 B.n60 1.24928
R2618 B.n380 B.n379 1.24928
R2619 B.n396 B.n395 1.24928
C0 w_n3658_n4352# B 11.6496f
C1 VP VDD1 9.92008f
C2 VDD2 B 2.68251f
C3 VN VDD1 0.151081f
C4 VTAIL VDD1 9.52513f
C5 VP VN 8.264549f
C6 VP VTAIL 9.63331f
C7 VN VTAIL 9.619f
C8 B VDD1 2.5981f
C9 VP B 2.10523f
C10 VN B 1.31146f
C11 B VTAIL 4.99536f
C12 VDD2 w_n3658_n4352# 2.83516f
C13 w_n3658_n4352# VDD1 2.73636f
C14 VP w_n3658_n4352# 7.613451f
C15 VDD2 VDD1 1.57577f
C16 VDD2 VP 0.494878f
C17 VN w_n3658_n4352# 7.13932f
C18 w_n3658_n4352# VTAIL 3.68976f
C19 VDD2 VN 9.58014f
C20 VDD2 VTAIL 9.578279f
C21 VDD2 VSUBS 2.14656f
C22 VDD1 VSUBS 2.110301f
C23 VTAIL VSUBS 1.457729f
C24 VN VSUBS 6.44128f
C25 VP VSUBS 3.457886f
C26 B VSUBS 5.478882f
C27 w_n3658_n4352# VSUBS 0.194854p
C28 B.n0 VSUBS 0.006785f
C29 B.n1 VSUBS 0.006785f
C30 B.n2 VSUBS 0.010034f
C31 B.n3 VSUBS 0.007689f
C32 B.n4 VSUBS 0.007689f
C33 B.n5 VSUBS 0.007689f
C34 B.n6 VSUBS 0.007689f
C35 B.n7 VSUBS 0.007689f
C36 B.n8 VSUBS 0.007689f
C37 B.n9 VSUBS 0.007689f
C38 B.n10 VSUBS 0.007689f
C39 B.n11 VSUBS 0.007689f
C40 B.n12 VSUBS 0.007689f
C41 B.n13 VSUBS 0.007689f
C42 B.n14 VSUBS 0.007689f
C43 B.n15 VSUBS 0.007689f
C44 B.n16 VSUBS 0.007689f
C45 B.n17 VSUBS 0.007689f
C46 B.n18 VSUBS 0.007689f
C47 B.n19 VSUBS 0.007689f
C48 B.n20 VSUBS 0.007689f
C49 B.n21 VSUBS 0.007689f
C50 B.n22 VSUBS 0.007689f
C51 B.n23 VSUBS 0.007689f
C52 B.n24 VSUBS 0.007689f
C53 B.n25 VSUBS 0.017347f
C54 B.n26 VSUBS 0.007689f
C55 B.n27 VSUBS 0.007689f
C56 B.n28 VSUBS 0.007689f
C57 B.n29 VSUBS 0.007689f
C58 B.n30 VSUBS 0.007689f
C59 B.n31 VSUBS 0.007689f
C60 B.n32 VSUBS 0.007689f
C61 B.n33 VSUBS 0.007689f
C62 B.n34 VSUBS 0.007689f
C63 B.n35 VSUBS 0.007689f
C64 B.n36 VSUBS 0.007689f
C65 B.n37 VSUBS 0.007689f
C66 B.n38 VSUBS 0.007689f
C67 B.n39 VSUBS 0.007689f
C68 B.n40 VSUBS 0.007689f
C69 B.n41 VSUBS 0.007689f
C70 B.n42 VSUBS 0.007689f
C71 B.n43 VSUBS 0.007689f
C72 B.n44 VSUBS 0.007689f
C73 B.n45 VSUBS 0.007689f
C74 B.n46 VSUBS 0.007689f
C75 B.n47 VSUBS 0.007689f
C76 B.n48 VSUBS 0.007689f
C77 B.n49 VSUBS 0.007689f
C78 B.n50 VSUBS 0.007689f
C79 B.n51 VSUBS 0.007689f
C80 B.n52 VSUBS 0.007689f
C81 B.n53 VSUBS 0.007689f
C82 B.t4 VSUBS 0.357243f
C83 B.t5 VSUBS 0.398786f
C84 B.t3 VSUBS 2.53649f
C85 B.n54 VSUBS 0.624072f
C86 B.n55 VSUBS 0.348553f
C87 B.n56 VSUBS 0.007689f
C88 B.n57 VSUBS 0.007689f
C89 B.n58 VSUBS 0.007689f
C90 B.n59 VSUBS 0.007689f
C91 B.n60 VSUBS 0.004297f
C92 B.n61 VSUBS 0.007689f
C93 B.t1 VSUBS 0.357247f
C94 B.t2 VSUBS 0.398789f
C95 B.t0 VSUBS 2.53649f
C96 B.n62 VSUBS 0.624069f
C97 B.n63 VSUBS 0.348549f
C98 B.n64 VSUBS 0.017815f
C99 B.n65 VSUBS 0.007689f
C100 B.n66 VSUBS 0.007689f
C101 B.n67 VSUBS 0.007689f
C102 B.n68 VSUBS 0.007689f
C103 B.n69 VSUBS 0.007689f
C104 B.n70 VSUBS 0.007689f
C105 B.n71 VSUBS 0.007689f
C106 B.n72 VSUBS 0.007689f
C107 B.n73 VSUBS 0.007689f
C108 B.n74 VSUBS 0.007689f
C109 B.n75 VSUBS 0.007689f
C110 B.n76 VSUBS 0.007689f
C111 B.n77 VSUBS 0.007689f
C112 B.n78 VSUBS 0.007689f
C113 B.n79 VSUBS 0.007689f
C114 B.n80 VSUBS 0.007689f
C115 B.n81 VSUBS 0.007689f
C116 B.n82 VSUBS 0.007689f
C117 B.n83 VSUBS 0.007689f
C118 B.n84 VSUBS 0.007689f
C119 B.n85 VSUBS 0.007689f
C120 B.n86 VSUBS 0.007689f
C121 B.n87 VSUBS 0.007689f
C122 B.n88 VSUBS 0.007689f
C123 B.n89 VSUBS 0.007689f
C124 B.n90 VSUBS 0.007689f
C125 B.n91 VSUBS 0.018612f
C126 B.n92 VSUBS 0.007689f
C127 B.n93 VSUBS 0.007689f
C128 B.n94 VSUBS 0.007689f
C129 B.n95 VSUBS 0.007689f
C130 B.n96 VSUBS 0.007689f
C131 B.n97 VSUBS 0.007689f
C132 B.n98 VSUBS 0.007689f
C133 B.n99 VSUBS 0.007689f
C134 B.n100 VSUBS 0.007689f
C135 B.n101 VSUBS 0.007689f
C136 B.n102 VSUBS 0.007689f
C137 B.n103 VSUBS 0.007689f
C138 B.n104 VSUBS 0.007689f
C139 B.n105 VSUBS 0.007689f
C140 B.n106 VSUBS 0.007689f
C141 B.n107 VSUBS 0.007689f
C142 B.n108 VSUBS 0.007689f
C143 B.n109 VSUBS 0.007689f
C144 B.n110 VSUBS 0.007689f
C145 B.n111 VSUBS 0.007689f
C146 B.n112 VSUBS 0.007689f
C147 B.n113 VSUBS 0.007689f
C148 B.n114 VSUBS 0.007689f
C149 B.n115 VSUBS 0.007689f
C150 B.n116 VSUBS 0.007689f
C151 B.n117 VSUBS 0.007689f
C152 B.n118 VSUBS 0.007689f
C153 B.n119 VSUBS 0.007689f
C154 B.n120 VSUBS 0.007689f
C155 B.n121 VSUBS 0.007689f
C156 B.n122 VSUBS 0.007689f
C157 B.n123 VSUBS 0.007689f
C158 B.n124 VSUBS 0.007689f
C159 B.n125 VSUBS 0.007689f
C160 B.n126 VSUBS 0.007689f
C161 B.n127 VSUBS 0.007689f
C162 B.n128 VSUBS 0.007689f
C163 B.n129 VSUBS 0.007689f
C164 B.n130 VSUBS 0.007689f
C165 B.n131 VSUBS 0.007689f
C166 B.n132 VSUBS 0.007689f
C167 B.n133 VSUBS 0.007689f
C168 B.n134 VSUBS 0.007689f
C169 B.n135 VSUBS 0.007689f
C170 B.n136 VSUBS 0.007689f
C171 B.n137 VSUBS 0.007689f
C172 B.n138 VSUBS 0.007689f
C173 B.n139 VSUBS 0.018257f
C174 B.n140 VSUBS 0.007689f
C175 B.n141 VSUBS 0.007689f
C176 B.n142 VSUBS 0.007689f
C177 B.n143 VSUBS 0.007689f
C178 B.n144 VSUBS 0.007689f
C179 B.n145 VSUBS 0.007689f
C180 B.n146 VSUBS 0.007689f
C181 B.n147 VSUBS 0.007689f
C182 B.n148 VSUBS 0.007689f
C183 B.n149 VSUBS 0.007689f
C184 B.n150 VSUBS 0.007689f
C185 B.n151 VSUBS 0.007689f
C186 B.n152 VSUBS 0.007689f
C187 B.n153 VSUBS 0.007689f
C188 B.n154 VSUBS 0.007689f
C189 B.n155 VSUBS 0.007689f
C190 B.n156 VSUBS 0.007689f
C191 B.n157 VSUBS 0.007689f
C192 B.n158 VSUBS 0.007689f
C193 B.n159 VSUBS 0.007689f
C194 B.n160 VSUBS 0.007689f
C195 B.n161 VSUBS 0.007689f
C196 B.n162 VSUBS 0.007689f
C197 B.n163 VSUBS 0.007689f
C198 B.n164 VSUBS 0.007689f
C199 B.n165 VSUBS 0.007689f
C200 B.n166 VSUBS 0.007689f
C201 B.n167 VSUBS 0.007237f
C202 B.n168 VSUBS 0.007689f
C203 B.n169 VSUBS 0.007689f
C204 B.n170 VSUBS 0.007689f
C205 B.n171 VSUBS 0.007689f
C206 B.n172 VSUBS 0.007689f
C207 B.t8 VSUBS 0.357243f
C208 B.t7 VSUBS 0.398786f
C209 B.t6 VSUBS 2.53649f
C210 B.n173 VSUBS 0.624072f
C211 B.n174 VSUBS 0.348553f
C212 B.n175 VSUBS 0.007689f
C213 B.n176 VSUBS 0.007689f
C214 B.n177 VSUBS 0.007689f
C215 B.n178 VSUBS 0.007689f
C216 B.n179 VSUBS 0.007689f
C217 B.n180 VSUBS 0.007689f
C218 B.n181 VSUBS 0.007689f
C219 B.n182 VSUBS 0.007689f
C220 B.n183 VSUBS 0.007689f
C221 B.n184 VSUBS 0.007689f
C222 B.n185 VSUBS 0.007689f
C223 B.n186 VSUBS 0.007689f
C224 B.n187 VSUBS 0.007689f
C225 B.n188 VSUBS 0.007689f
C226 B.n189 VSUBS 0.007689f
C227 B.n190 VSUBS 0.007689f
C228 B.n191 VSUBS 0.007689f
C229 B.n192 VSUBS 0.007689f
C230 B.n193 VSUBS 0.007689f
C231 B.n194 VSUBS 0.007689f
C232 B.n195 VSUBS 0.007689f
C233 B.n196 VSUBS 0.007689f
C234 B.n197 VSUBS 0.007689f
C235 B.n198 VSUBS 0.007689f
C236 B.n199 VSUBS 0.007689f
C237 B.n200 VSUBS 0.007689f
C238 B.n201 VSUBS 0.007689f
C239 B.n202 VSUBS 0.018612f
C240 B.n203 VSUBS 0.007689f
C241 B.n204 VSUBS 0.007689f
C242 B.n205 VSUBS 0.007689f
C243 B.n206 VSUBS 0.007689f
C244 B.n207 VSUBS 0.007689f
C245 B.n208 VSUBS 0.007689f
C246 B.n209 VSUBS 0.007689f
C247 B.n210 VSUBS 0.007689f
C248 B.n211 VSUBS 0.007689f
C249 B.n212 VSUBS 0.007689f
C250 B.n213 VSUBS 0.007689f
C251 B.n214 VSUBS 0.007689f
C252 B.n215 VSUBS 0.007689f
C253 B.n216 VSUBS 0.007689f
C254 B.n217 VSUBS 0.007689f
C255 B.n218 VSUBS 0.007689f
C256 B.n219 VSUBS 0.007689f
C257 B.n220 VSUBS 0.007689f
C258 B.n221 VSUBS 0.007689f
C259 B.n222 VSUBS 0.007689f
C260 B.n223 VSUBS 0.007689f
C261 B.n224 VSUBS 0.007689f
C262 B.n225 VSUBS 0.007689f
C263 B.n226 VSUBS 0.007689f
C264 B.n227 VSUBS 0.007689f
C265 B.n228 VSUBS 0.007689f
C266 B.n229 VSUBS 0.007689f
C267 B.n230 VSUBS 0.007689f
C268 B.n231 VSUBS 0.007689f
C269 B.n232 VSUBS 0.007689f
C270 B.n233 VSUBS 0.007689f
C271 B.n234 VSUBS 0.007689f
C272 B.n235 VSUBS 0.007689f
C273 B.n236 VSUBS 0.007689f
C274 B.n237 VSUBS 0.007689f
C275 B.n238 VSUBS 0.007689f
C276 B.n239 VSUBS 0.007689f
C277 B.n240 VSUBS 0.007689f
C278 B.n241 VSUBS 0.007689f
C279 B.n242 VSUBS 0.007689f
C280 B.n243 VSUBS 0.007689f
C281 B.n244 VSUBS 0.007689f
C282 B.n245 VSUBS 0.007689f
C283 B.n246 VSUBS 0.007689f
C284 B.n247 VSUBS 0.007689f
C285 B.n248 VSUBS 0.007689f
C286 B.n249 VSUBS 0.007689f
C287 B.n250 VSUBS 0.007689f
C288 B.n251 VSUBS 0.007689f
C289 B.n252 VSUBS 0.007689f
C290 B.n253 VSUBS 0.007689f
C291 B.n254 VSUBS 0.007689f
C292 B.n255 VSUBS 0.007689f
C293 B.n256 VSUBS 0.007689f
C294 B.n257 VSUBS 0.007689f
C295 B.n258 VSUBS 0.007689f
C296 B.n259 VSUBS 0.007689f
C297 B.n260 VSUBS 0.007689f
C298 B.n261 VSUBS 0.007689f
C299 B.n262 VSUBS 0.007689f
C300 B.n263 VSUBS 0.007689f
C301 B.n264 VSUBS 0.007689f
C302 B.n265 VSUBS 0.007689f
C303 B.n266 VSUBS 0.007689f
C304 B.n267 VSUBS 0.007689f
C305 B.n268 VSUBS 0.007689f
C306 B.n269 VSUBS 0.007689f
C307 B.n270 VSUBS 0.007689f
C308 B.n271 VSUBS 0.007689f
C309 B.n272 VSUBS 0.007689f
C310 B.n273 VSUBS 0.007689f
C311 B.n274 VSUBS 0.007689f
C312 B.n275 VSUBS 0.007689f
C313 B.n276 VSUBS 0.007689f
C314 B.n277 VSUBS 0.007689f
C315 B.n278 VSUBS 0.007689f
C316 B.n279 VSUBS 0.007689f
C317 B.n280 VSUBS 0.007689f
C318 B.n281 VSUBS 0.007689f
C319 B.n282 VSUBS 0.007689f
C320 B.n283 VSUBS 0.007689f
C321 B.n284 VSUBS 0.007689f
C322 B.n285 VSUBS 0.007689f
C323 B.n286 VSUBS 0.007689f
C324 B.n287 VSUBS 0.007689f
C325 B.n288 VSUBS 0.007689f
C326 B.n289 VSUBS 0.007689f
C327 B.n290 VSUBS 0.007689f
C328 B.n291 VSUBS 0.007689f
C329 B.n292 VSUBS 0.007689f
C330 B.n293 VSUBS 0.017347f
C331 B.n294 VSUBS 0.017347f
C332 B.n295 VSUBS 0.018612f
C333 B.n296 VSUBS 0.007689f
C334 B.n297 VSUBS 0.007689f
C335 B.n298 VSUBS 0.007689f
C336 B.n299 VSUBS 0.007689f
C337 B.n300 VSUBS 0.007689f
C338 B.n301 VSUBS 0.007689f
C339 B.n302 VSUBS 0.007689f
C340 B.n303 VSUBS 0.007689f
C341 B.n304 VSUBS 0.007689f
C342 B.n305 VSUBS 0.007689f
C343 B.n306 VSUBS 0.007689f
C344 B.n307 VSUBS 0.007689f
C345 B.n308 VSUBS 0.007689f
C346 B.n309 VSUBS 0.007689f
C347 B.n310 VSUBS 0.007689f
C348 B.n311 VSUBS 0.007689f
C349 B.n312 VSUBS 0.007689f
C350 B.n313 VSUBS 0.007689f
C351 B.n314 VSUBS 0.007689f
C352 B.n315 VSUBS 0.007689f
C353 B.n316 VSUBS 0.007689f
C354 B.n317 VSUBS 0.007689f
C355 B.n318 VSUBS 0.007689f
C356 B.n319 VSUBS 0.007689f
C357 B.n320 VSUBS 0.007689f
C358 B.n321 VSUBS 0.007689f
C359 B.n322 VSUBS 0.007689f
C360 B.n323 VSUBS 0.007689f
C361 B.n324 VSUBS 0.007689f
C362 B.n325 VSUBS 0.007689f
C363 B.n326 VSUBS 0.007689f
C364 B.n327 VSUBS 0.007689f
C365 B.n328 VSUBS 0.007689f
C366 B.n329 VSUBS 0.007689f
C367 B.n330 VSUBS 0.007689f
C368 B.n331 VSUBS 0.007689f
C369 B.n332 VSUBS 0.007689f
C370 B.n333 VSUBS 0.007689f
C371 B.n334 VSUBS 0.007689f
C372 B.n335 VSUBS 0.007689f
C373 B.n336 VSUBS 0.007689f
C374 B.n337 VSUBS 0.007689f
C375 B.n338 VSUBS 0.007689f
C376 B.n339 VSUBS 0.007689f
C377 B.n340 VSUBS 0.007689f
C378 B.n341 VSUBS 0.007689f
C379 B.n342 VSUBS 0.007689f
C380 B.n343 VSUBS 0.007689f
C381 B.n344 VSUBS 0.007689f
C382 B.n345 VSUBS 0.007689f
C383 B.n346 VSUBS 0.007689f
C384 B.n347 VSUBS 0.007689f
C385 B.n348 VSUBS 0.007689f
C386 B.n349 VSUBS 0.007689f
C387 B.n350 VSUBS 0.007689f
C388 B.n351 VSUBS 0.007689f
C389 B.n352 VSUBS 0.007689f
C390 B.n353 VSUBS 0.007689f
C391 B.n354 VSUBS 0.007689f
C392 B.n355 VSUBS 0.007689f
C393 B.n356 VSUBS 0.007689f
C394 B.n357 VSUBS 0.007689f
C395 B.n358 VSUBS 0.007689f
C396 B.n359 VSUBS 0.007689f
C397 B.n360 VSUBS 0.007689f
C398 B.n361 VSUBS 0.007689f
C399 B.n362 VSUBS 0.007689f
C400 B.n363 VSUBS 0.007689f
C401 B.n364 VSUBS 0.007689f
C402 B.n365 VSUBS 0.007689f
C403 B.n366 VSUBS 0.007689f
C404 B.n367 VSUBS 0.007689f
C405 B.n368 VSUBS 0.007689f
C406 B.n369 VSUBS 0.007689f
C407 B.n370 VSUBS 0.007689f
C408 B.n371 VSUBS 0.007689f
C409 B.n372 VSUBS 0.007689f
C410 B.n373 VSUBS 0.007689f
C411 B.n374 VSUBS 0.007689f
C412 B.n375 VSUBS 0.007689f
C413 B.n376 VSUBS 0.007689f
C414 B.n377 VSUBS 0.007689f
C415 B.n378 VSUBS 0.007237f
C416 B.n379 VSUBS 0.017815f
C417 B.n380 VSUBS 0.004297f
C418 B.n381 VSUBS 0.007689f
C419 B.n382 VSUBS 0.007689f
C420 B.n383 VSUBS 0.007689f
C421 B.n384 VSUBS 0.007689f
C422 B.n385 VSUBS 0.007689f
C423 B.n386 VSUBS 0.007689f
C424 B.n387 VSUBS 0.007689f
C425 B.n388 VSUBS 0.007689f
C426 B.n389 VSUBS 0.007689f
C427 B.n390 VSUBS 0.007689f
C428 B.n391 VSUBS 0.007689f
C429 B.n392 VSUBS 0.007689f
C430 B.t11 VSUBS 0.357247f
C431 B.t10 VSUBS 0.398789f
C432 B.t9 VSUBS 2.53649f
C433 B.n393 VSUBS 0.624069f
C434 B.n394 VSUBS 0.348549f
C435 B.n395 VSUBS 0.017815f
C436 B.n396 VSUBS 0.004297f
C437 B.n397 VSUBS 0.007689f
C438 B.n398 VSUBS 0.007689f
C439 B.n399 VSUBS 0.007689f
C440 B.n400 VSUBS 0.007689f
C441 B.n401 VSUBS 0.007689f
C442 B.n402 VSUBS 0.007689f
C443 B.n403 VSUBS 0.007689f
C444 B.n404 VSUBS 0.007689f
C445 B.n405 VSUBS 0.007689f
C446 B.n406 VSUBS 0.007689f
C447 B.n407 VSUBS 0.007689f
C448 B.n408 VSUBS 0.007689f
C449 B.n409 VSUBS 0.007689f
C450 B.n410 VSUBS 0.007689f
C451 B.n411 VSUBS 0.007689f
C452 B.n412 VSUBS 0.007689f
C453 B.n413 VSUBS 0.007689f
C454 B.n414 VSUBS 0.007689f
C455 B.n415 VSUBS 0.007689f
C456 B.n416 VSUBS 0.007689f
C457 B.n417 VSUBS 0.007689f
C458 B.n418 VSUBS 0.007689f
C459 B.n419 VSUBS 0.007689f
C460 B.n420 VSUBS 0.007689f
C461 B.n421 VSUBS 0.007689f
C462 B.n422 VSUBS 0.007689f
C463 B.n423 VSUBS 0.007689f
C464 B.n424 VSUBS 0.007689f
C465 B.n425 VSUBS 0.007689f
C466 B.n426 VSUBS 0.007689f
C467 B.n427 VSUBS 0.007689f
C468 B.n428 VSUBS 0.007689f
C469 B.n429 VSUBS 0.007689f
C470 B.n430 VSUBS 0.007689f
C471 B.n431 VSUBS 0.007689f
C472 B.n432 VSUBS 0.007689f
C473 B.n433 VSUBS 0.007689f
C474 B.n434 VSUBS 0.007689f
C475 B.n435 VSUBS 0.007689f
C476 B.n436 VSUBS 0.007689f
C477 B.n437 VSUBS 0.007689f
C478 B.n438 VSUBS 0.007689f
C479 B.n439 VSUBS 0.007689f
C480 B.n440 VSUBS 0.007689f
C481 B.n441 VSUBS 0.007689f
C482 B.n442 VSUBS 0.007689f
C483 B.n443 VSUBS 0.007689f
C484 B.n444 VSUBS 0.007689f
C485 B.n445 VSUBS 0.007689f
C486 B.n446 VSUBS 0.007689f
C487 B.n447 VSUBS 0.007689f
C488 B.n448 VSUBS 0.007689f
C489 B.n449 VSUBS 0.007689f
C490 B.n450 VSUBS 0.007689f
C491 B.n451 VSUBS 0.007689f
C492 B.n452 VSUBS 0.007689f
C493 B.n453 VSUBS 0.007689f
C494 B.n454 VSUBS 0.007689f
C495 B.n455 VSUBS 0.007689f
C496 B.n456 VSUBS 0.007689f
C497 B.n457 VSUBS 0.007689f
C498 B.n458 VSUBS 0.007689f
C499 B.n459 VSUBS 0.007689f
C500 B.n460 VSUBS 0.007689f
C501 B.n461 VSUBS 0.007689f
C502 B.n462 VSUBS 0.007689f
C503 B.n463 VSUBS 0.007689f
C504 B.n464 VSUBS 0.007689f
C505 B.n465 VSUBS 0.007689f
C506 B.n466 VSUBS 0.007689f
C507 B.n467 VSUBS 0.007689f
C508 B.n468 VSUBS 0.007689f
C509 B.n469 VSUBS 0.007689f
C510 B.n470 VSUBS 0.007689f
C511 B.n471 VSUBS 0.007689f
C512 B.n472 VSUBS 0.007689f
C513 B.n473 VSUBS 0.007689f
C514 B.n474 VSUBS 0.007689f
C515 B.n475 VSUBS 0.007689f
C516 B.n476 VSUBS 0.007689f
C517 B.n477 VSUBS 0.007689f
C518 B.n478 VSUBS 0.007689f
C519 B.n479 VSUBS 0.007689f
C520 B.n480 VSUBS 0.017702f
C521 B.n481 VSUBS 0.018612f
C522 B.n482 VSUBS 0.017347f
C523 B.n483 VSUBS 0.007689f
C524 B.n484 VSUBS 0.007689f
C525 B.n485 VSUBS 0.007689f
C526 B.n486 VSUBS 0.007689f
C527 B.n487 VSUBS 0.007689f
C528 B.n488 VSUBS 0.007689f
C529 B.n489 VSUBS 0.007689f
C530 B.n490 VSUBS 0.007689f
C531 B.n491 VSUBS 0.007689f
C532 B.n492 VSUBS 0.007689f
C533 B.n493 VSUBS 0.007689f
C534 B.n494 VSUBS 0.007689f
C535 B.n495 VSUBS 0.007689f
C536 B.n496 VSUBS 0.007689f
C537 B.n497 VSUBS 0.007689f
C538 B.n498 VSUBS 0.007689f
C539 B.n499 VSUBS 0.007689f
C540 B.n500 VSUBS 0.007689f
C541 B.n501 VSUBS 0.007689f
C542 B.n502 VSUBS 0.007689f
C543 B.n503 VSUBS 0.007689f
C544 B.n504 VSUBS 0.007689f
C545 B.n505 VSUBS 0.007689f
C546 B.n506 VSUBS 0.007689f
C547 B.n507 VSUBS 0.007689f
C548 B.n508 VSUBS 0.007689f
C549 B.n509 VSUBS 0.007689f
C550 B.n510 VSUBS 0.007689f
C551 B.n511 VSUBS 0.007689f
C552 B.n512 VSUBS 0.007689f
C553 B.n513 VSUBS 0.007689f
C554 B.n514 VSUBS 0.007689f
C555 B.n515 VSUBS 0.007689f
C556 B.n516 VSUBS 0.007689f
C557 B.n517 VSUBS 0.007689f
C558 B.n518 VSUBS 0.007689f
C559 B.n519 VSUBS 0.007689f
C560 B.n520 VSUBS 0.007689f
C561 B.n521 VSUBS 0.007689f
C562 B.n522 VSUBS 0.007689f
C563 B.n523 VSUBS 0.007689f
C564 B.n524 VSUBS 0.007689f
C565 B.n525 VSUBS 0.007689f
C566 B.n526 VSUBS 0.007689f
C567 B.n527 VSUBS 0.007689f
C568 B.n528 VSUBS 0.007689f
C569 B.n529 VSUBS 0.007689f
C570 B.n530 VSUBS 0.007689f
C571 B.n531 VSUBS 0.007689f
C572 B.n532 VSUBS 0.007689f
C573 B.n533 VSUBS 0.007689f
C574 B.n534 VSUBS 0.007689f
C575 B.n535 VSUBS 0.007689f
C576 B.n536 VSUBS 0.007689f
C577 B.n537 VSUBS 0.007689f
C578 B.n538 VSUBS 0.007689f
C579 B.n539 VSUBS 0.007689f
C580 B.n540 VSUBS 0.007689f
C581 B.n541 VSUBS 0.007689f
C582 B.n542 VSUBS 0.007689f
C583 B.n543 VSUBS 0.007689f
C584 B.n544 VSUBS 0.007689f
C585 B.n545 VSUBS 0.007689f
C586 B.n546 VSUBS 0.007689f
C587 B.n547 VSUBS 0.007689f
C588 B.n548 VSUBS 0.007689f
C589 B.n549 VSUBS 0.007689f
C590 B.n550 VSUBS 0.007689f
C591 B.n551 VSUBS 0.007689f
C592 B.n552 VSUBS 0.007689f
C593 B.n553 VSUBS 0.007689f
C594 B.n554 VSUBS 0.007689f
C595 B.n555 VSUBS 0.007689f
C596 B.n556 VSUBS 0.007689f
C597 B.n557 VSUBS 0.007689f
C598 B.n558 VSUBS 0.007689f
C599 B.n559 VSUBS 0.007689f
C600 B.n560 VSUBS 0.007689f
C601 B.n561 VSUBS 0.007689f
C602 B.n562 VSUBS 0.007689f
C603 B.n563 VSUBS 0.007689f
C604 B.n564 VSUBS 0.007689f
C605 B.n565 VSUBS 0.007689f
C606 B.n566 VSUBS 0.007689f
C607 B.n567 VSUBS 0.007689f
C608 B.n568 VSUBS 0.007689f
C609 B.n569 VSUBS 0.007689f
C610 B.n570 VSUBS 0.007689f
C611 B.n571 VSUBS 0.007689f
C612 B.n572 VSUBS 0.007689f
C613 B.n573 VSUBS 0.007689f
C614 B.n574 VSUBS 0.007689f
C615 B.n575 VSUBS 0.007689f
C616 B.n576 VSUBS 0.007689f
C617 B.n577 VSUBS 0.007689f
C618 B.n578 VSUBS 0.007689f
C619 B.n579 VSUBS 0.007689f
C620 B.n580 VSUBS 0.007689f
C621 B.n581 VSUBS 0.007689f
C622 B.n582 VSUBS 0.007689f
C623 B.n583 VSUBS 0.007689f
C624 B.n584 VSUBS 0.007689f
C625 B.n585 VSUBS 0.007689f
C626 B.n586 VSUBS 0.007689f
C627 B.n587 VSUBS 0.007689f
C628 B.n588 VSUBS 0.007689f
C629 B.n589 VSUBS 0.007689f
C630 B.n590 VSUBS 0.007689f
C631 B.n591 VSUBS 0.007689f
C632 B.n592 VSUBS 0.007689f
C633 B.n593 VSUBS 0.007689f
C634 B.n594 VSUBS 0.007689f
C635 B.n595 VSUBS 0.007689f
C636 B.n596 VSUBS 0.007689f
C637 B.n597 VSUBS 0.007689f
C638 B.n598 VSUBS 0.007689f
C639 B.n599 VSUBS 0.007689f
C640 B.n600 VSUBS 0.007689f
C641 B.n601 VSUBS 0.007689f
C642 B.n602 VSUBS 0.007689f
C643 B.n603 VSUBS 0.007689f
C644 B.n604 VSUBS 0.007689f
C645 B.n605 VSUBS 0.007689f
C646 B.n606 VSUBS 0.007689f
C647 B.n607 VSUBS 0.007689f
C648 B.n608 VSUBS 0.007689f
C649 B.n609 VSUBS 0.007689f
C650 B.n610 VSUBS 0.007689f
C651 B.n611 VSUBS 0.007689f
C652 B.n612 VSUBS 0.007689f
C653 B.n613 VSUBS 0.007689f
C654 B.n614 VSUBS 0.007689f
C655 B.n615 VSUBS 0.007689f
C656 B.n616 VSUBS 0.007689f
C657 B.n617 VSUBS 0.007689f
C658 B.n618 VSUBS 0.007689f
C659 B.n619 VSUBS 0.007689f
C660 B.n620 VSUBS 0.007689f
C661 B.n621 VSUBS 0.007689f
C662 B.n622 VSUBS 0.007689f
C663 B.n623 VSUBS 0.007689f
C664 B.n624 VSUBS 0.017347f
C665 B.n625 VSUBS 0.017347f
C666 B.n626 VSUBS 0.018612f
C667 B.n627 VSUBS 0.007689f
C668 B.n628 VSUBS 0.007689f
C669 B.n629 VSUBS 0.007689f
C670 B.n630 VSUBS 0.007689f
C671 B.n631 VSUBS 0.007689f
C672 B.n632 VSUBS 0.007689f
C673 B.n633 VSUBS 0.007689f
C674 B.n634 VSUBS 0.007689f
C675 B.n635 VSUBS 0.007689f
C676 B.n636 VSUBS 0.007689f
C677 B.n637 VSUBS 0.007689f
C678 B.n638 VSUBS 0.007689f
C679 B.n639 VSUBS 0.007689f
C680 B.n640 VSUBS 0.007689f
C681 B.n641 VSUBS 0.007689f
C682 B.n642 VSUBS 0.007689f
C683 B.n643 VSUBS 0.007689f
C684 B.n644 VSUBS 0.007689f
C685 B.n645 VSUBS 0.007689f
C686 B.n646 VSUBS 0.007689f
C687 B.n647 VSUBS 0.007689f
C688 B.n648 VSUBS 0.007689f
C689 B.n649 VSUBS 0.007689f
C690 B.n650 VSUBS 0.007689f
C691 B.n651 VSUBS 0.007689f
C692 B.n652 VSUBS 0.007689f
C693 B.n653 VSUBS 0.007689f
C694 B.n654 VSUBS 0.007689f
C695 B.n655 VSUBS 0.007689f
C696 B.n656 VSUBS 0.007689f
C697 B.n657 VSUBS 0.007689f
C698 B.n658 VSUBS 0.007689f
C699 B.n659 VSUBS 0.007689f
C700 B.n660 VSUBS 0.007689f
C701 B.n661 VSUBS 0.007689f
C702 B.n662 VSUBS 0.007689f
C703 B.n663 VSUBS 0.007689f
C704 B.n664 VSUBS 0.007689f
C705 B.n665 VSUBS 0.007689f
C706 B.n666 VSUBS 0.007689f
C707 B.n667 VSUBS 0.007689f
C708 B.n668 VSUBS 0.007689f
C709 B.n669 VSUBS 0.007689f
C710 B.n670 VSUBS 0.007689f
C711 B.n671 VSUBS 0.007689f
C712 B.n672 VSUBS 0.007689f
C713 B.n673 VSUBS 0.007689f
C714 B.n674 VSUBS 0.007689f
C715 B.n675 VSUBS 0.007689f
C716 B.n676 VSUBS 0.007689f
C717 B.n677 VSUBS 0.007689f
C718 B.n678 VSUBS 0.007689f
C719 B.n679 VSUBS 0.007689f
C720 B.n680 VSUBS 0.007689f
C721 B.n681 VSUBS 0.007689f
C722 B.n682 VSUBS 0.007689f
C723 B.n683 VSUBS 0.007689f
C724 B.n684 VSUBS 0.007689f
C725 B.n685 VSUBS 0.007689f
C726 B.n686 VSUBS 0.007689f
C727 B.n687 VSUBS 0.007689f
C728 B.n688 VSUBS 0.007689f
C729 B.n689 VSUBS 0.007689f
C730 B.n690 VSUBS 0.007689f
C731 B.n691 VSUBS 0.007689f
C732 B.n692 VSUBS 0.007689f
C733 B.n693 VSUBS 0.007689f
C734 B.n694 VSUBS 0.007689f
C735 B.n695 VSUBS 0.007689f
C736 B.n696 VSUBS 0.007689f
C737 B.n697 VSUBS 0.007689f
C738 B.n698 VSUBS 0.007689f
C739 B.n699 VSUBS 0.007689f
C740 B.n700 VSUBS 0.007689f
C741 B.n701 VSUBS 0.007689f
C742 B.n702 VSUBS 0.007689f
C743 B.n703 VSUBS 0.007689f
C744 B.n704 VSUBS 0.007689f
C745 B.n705 VSUBS 0.007689f
C746 B.n706 VSUBS 0.007689f
C747 B.n707 VSUBS 0.007689f
C748 B.n708 VSUBS 0.007237f
C749 B.n709 VSUBS 0.007689f
C750 B.n710 VSUBS 0.007689f
C751 B.n711 VSUBS 0.007689f
C752 B.n712 VSUBS 0.007689f
C753 B.n713 VSUBS 0.007689f
C754 B.n714 VSUBS 0.007689f
C755 B.n715 VSUBS 0.007689f
C756 B.n716 VSUBS 0.007689f
C757 B.n717 VSUBS 0.007689f
C758 B.n718 VSUBS 0.007689f
C759 B.n719 VSUBS 0.007689f
C760 B.n720 VSUBS 0.007689f
C761 B.n721 VSUBS 0.007689f
C762 B.n722 VSUBS 0.007689f
C763 B.n723 VSUBS 0.007689f
C764 B.n724 VSUBS 0.004297f
C765 B.n725 VSUBS 0.017815f
C766 B.n726 VSUBS 0.007237f
C767 B.n727 VSUBS 0.007689f
C768 B.n728 VSUBS 0.007689f
C769 B.n729 VSUBS 0.007689f
C770 B.n730 VSUBS 0.007689f
C771 B.n731 VSUBS 0.007689f
C772 B.n732 VSUBS 0.007689f
C773 B.n733 VSUBS 0.007689f
C774 B.n734 VSUBS 0.007689f
C775 B.n735 VSUBS 0.007689f
C776 B.n736 VSUBS 0.007689f
C777 B.n737 VSUBS 0.007689f
C778 B.n738 VSUBS 0.007689f
C779 B.n739 VSUBS 0.007689f
C780 B.n740 VSUBS 0.007689f
C781 B.n741 VSUBS 0.007689f
C782 B.n742 VSUBS 0.007689f
C783 B.n743 VSUBS 0.007689f
C784 B.n744 VSUBS 0.007689f
C785 B.n745 VSUBS 0.007689f
C786 B.n746 VSUBS 0.007689f
C787 B.n747 VSUBS 0.007689f
C788 B.n748 VSUBS 0.007689f
C789 B.n749 VSUBS 0.007689f
C790 B.n750 VSUBS 0.007689f
C791 B.n751 VSUBS 0.007689f
C792 B.n752 VSUBS 0.007689f
C793 B.n753 VSUBS 0.007689f
C794 B.n754 VSUBS 0.007689f
C795 B.n755 VSUBS 0.007689f
C796 B.n756 VSUBS 0.007689f
C797 B.n757 VSUBS 0.007689f
C798 B.n758 VSUBS 0.007689f
C799 B.n759 VSUBS 0.007689f
C800 B.n760 VSUBS 0.007689f
C801 B.n761 VSUBS 0.007689f
C802 B.n762 VSUBS 0.007689f
C803 B.n763 VSUBS 0.007689f
C804 B.n764 VSUBS 0.007689f
C805 B.n765 VSUBS 0.007689f
C806 B.n766 VSUBS 0.007689f
C807 B.n767 VSUBS 0.007689f
C808 B.n768 VSUBS 0.007689f
C809 B.n769 VSUBS 0.007689f
C810 B.n770 VSUBS 0.007689f
C811 B.n771 VSUBS 0.007689f
C812 B.n772 VSUBS 0.007689f
C813 B.n773 VSUBS 0.007689f
C814 B.n774 VSUBS 0.007689f
C815 B.n775 VSUBS 0.007689f
C816 B.n776 VSUBS 0.007689f
C817 B.n777 VSUBS 0.007689f
C818 B.n778 VSUBS 0.007689f
C819 B.n779 VSUBS 0.007689f
C820 B.n780 VSUBS 0.007689f
C821 B.n781 VSUBS 0.007689f
C822 B.n782 VSUBS 0.007689f
C823 B.n783 VSUBS 0.007689f
C824 B.n784 VSUBS 0.007689f
C825 B.n785 VSUBS 0.007689f
C826 B.n786 VSUBS 0.007689f
C827 B.n787 VSUBS 0.007689f
C828 B.n788 VSUBS 0.007689f
C829 B.n789 VSUBS 0.007689f
C830 B.n790 VSUBS 0.007689f
C831 B.n791 VSUBS 0.007689f
C832 B.n792 VSUBS 0.007689f
C833 B.n793 VSUBS 0.007689f
C834 B.n794 VSUBS 0.007689f
C835 B.n795 VSUBS 0.007689f
C836 B.n796 VSUBS 0.007689f
C837 B.n797 VSUBS 0.007689f
C838 B.n798 VSUBS 0.007689f
C839 B.n799 VSUBS 0.007689f
C840 B.n800 VSUBS 0.007689f
C841 B.n801 VSUBS 0.007689f
C842 B.n802 VSUBS 0.007689f
C843 B.n803 VSUBS 0.007689f
C844 B.n804 VSUBS 0.007689f
C845 B.n805 VSUBS 0.007689f
C846 B.n806 VSUBS 0.007689f
C847 B.n807 VSUBS 0.007689f
C848 B.n808 VSUBS 0.018612f
C849 B.n809 VSUBS 0.018612f
C850 B.n810 VSUBS 0.017347f
C851 B.n811 VSUBS 0.007689f
C852 B.n812 VSUBS 0.007689f
C853 B.n813 VSUBS 0.007689f
C854 B.n814 VSUBS 0.007689f
C855 B.n815 VSUBS 0.007689f
C856 B.n816 VSUBS 0.007689f
C857 B.n817 VSUBS 0.007689f
C858 B.n818 VSUBS 0.007689f
C859 B.n819 VSUBS 0.007689f
C860 B.n820 VSUBS 0.007689f
C861 B.n821 VSUBS 0.007689f
C862 B.n822 VSUBS 0.007689f
C863 B.n823 VSUBS 0.007689f
C864 B.n824 VSUBS 0.007689f
C865 B.n825 VSUBS 0.007689f
C866 B.n826 VSUBS 0.007689f
C867 B.n827 VSUBS 0.007689f
C868 B.n828 VSUBS 0.007689f
C869 B.n829 VSUBS 0.007689f
C870 B.n830 VSUBS 0.007689f
C871 B.n831 VSUBS 0.007689f
C872 B.n832 VSUBS 0.007689f
C873 B.n833 VSUBS 0.007689f
C874 B.n834 VSUBS 0.007689f
C875 B.n835 VSUBS 0.007689f
C876 B.n836 VSUBS 0.007689f
C877 B.n837 VSUBS 0.007689f
C878 B.n838 VSUBS 0.007689f
C879 B.n839 VSUBS 0.007689f
C880 B.n840 VSUBS 0.007689f
C881 B.n841 VSUBS 0.007689f
C882 B.n842 VSUBS 0.007689f
C883 B.n843 VSUBS 0.007689f
C884 B.n844 VSUBS 0.007689f
C885 B.n845 VSUBS 0.007689f
C886 B.n846 VSUBS 0.007689f
C887 B.n847 VSUBS 0.007689f
C888 B.n848 VSUBS 0.007689f
C889 B.n849 VSUBS 0.007689f
C890 B.n850 VSUBS 0.007689f
C891 B.n851 VSUBS 0.007689f
C892 B.n852 VSUBS 0.007689f
C893 B.n853 VSUBS 0.007689f
C894 B.n854 VSUBS 0.007689f
C895 B.n855 VSUBS 0.007689f
C896 B.n856 VSUBS 0.007689f
C897 B.n857 VSUBS 0.007689f
C898 B.n858 VSUBS 0.007689f
C899 B.n859 VSUBS 0.007689f
C900 B.n860 VSUBS 0.007689f
C901 B.n861 VSUBS 0.007689f
C902 B.n862 VSUBS 0.007689f
C903 B.n863 VSUBS 0.007689f
C904 B.n864 VSUBS 0.007689f
C905 B.n865 VSUBS 0.007689f
C906 B.n866 VSUBS 0.007689f
C907 B.n867 VSUBS 0.007689f
C908 B.n868 VSUBS 0.007689f
C909 B.n869 VSUBS 0.007689f
C910 B.n870 VSUBS 0.007689f
C911 B.n871 VSUBS 0.007689f
C912 B.n872 VSUBS 0.007689f
C913 B.n873 VSUBS 0.007689f
C914 B.n874 VSUBS 0.007689f
C915 B.n875 VSUBS 0.007689f
C916 B.n876 VSUBS 0.007689f
C917 B.n877 VSUBS 0.007689f
C918 B.n878 VSUBS 0.007689f
C919 B.n879 VSUBS 0.010034f
C920 B.n880 VSUBS 0.010689f
C921 B.n881 VSUBS 0.021256f
C922 VDD2.n0 VSUBS 0.030337f
C923 VDD2.n1 VSUBS 0.027292f
C924 VDD2.n2 VSUBS 0.014665f
C925 VDD2.n3 VSUBS 0.034664f
C926 VDD2.n4 VSUBS 0.015528f
C927 VDD2.n5 VSUBS 0.027292f
C928 VDD2.n6 VSUBS 0.014665f
C929 VDD2.n7 VSUBS 0.034664f
C930 VDD2.n8 VSUBS 0.015528f
C931 VDD2.n9 VSUBS 0.027292f
C932 VDD2.n10 VSUBS 0.014665f
C933 VDD2.n11 VSUBS 0.034664f
C934 VDD2.n12 VSUBS 0.015528f
C935 VDD2.n13 VSUBS 0.027292f
C936 VDD2.n14 VSUBS 0.014665f
C937 VDD2.n15 VSUBS 0.034664f
C938 VDD2.n16 VSUBS 0.015528f
C939 VDD2.n17 VSUBS 0.027292f
C940 VDD2.n18 VSUBS 0.014665f
C941 VDD2.n19 VSUBS 0.034664f
C942 VDD2.n20 VSUBS 0.015528f
C943 VDD2.n21 VSUBS 0.027292f
C944 VDD2.n22 VSUBS 0.014665f
C945 VDD2.n23 VSUBS 0.034664f
C946 VDD2.n24 VSUBS 0.015528f
C947 VDD2.n25 VSUBS 0.027292f
C948 VDD2.n26 VSUBS 0.014665f
C949 VDD2.n27 VSUBS 0.034664f
C950 VDD2.n28 VSUBS 0.015528f
C951 VDD2.n29 VSUBS 0.207839f
C952 VDD2.t0 VSUBS 0.074338f
C953 VDD2.n30 VSUBS 0.025998f
C954 VDD2.n31 VSUBS 0.022051f
C955 VDD2.n32 VSUBS 0.014665f
C956 VDD2.n33 VSUBS 1.98052f
C957 VDD2.n34 VSUBS 0.027292f
C958 VDD2.n35 VSUBS 0.014665f
C959 VDD2.n36 VSUBS 0.015528f
C960 VDD2.n37 VSUBS 0.034664f
C961 VDD2.n38 VSUBS 0.034664f
C962 VDD2.n39 VSUBS 0.015528f
C963 VDD2.n40 VSUBS 0.014665f
C964 VDD2.n41 VSUBS 0.027292f
C965 VDD2.n42 VSUBS 0.027292f
C966 VDD2.n43 VSUBS 0.014665f
C967 VDD2.n44 VSUBS 0.015528f
C968 VDD2.n45 VSUBS 0.034664f
C969 VDD2.n46 VSUBS 0.034664f
C970 VDD2.n47 VSUBS 0.015528f
C971 VDD2.n48 VSUBS 0.014665f
C972 VDD2.n49 VSUBS 0.027292f
C973 VDD2.n50 VSUBS 0.027292f
C974 VDD2.n51 VSUBS 0.014665f
C975 VDD2.n52 VSUBS 0.015528f
C976 VDD2.n53 VSUBS 0.034664f
C977 VDD2.n54 VSUBS 0.034664f
C978 VDD2.n55 VSUBS 0.015528f
C979 VDD2.n56 VSUBS 0.014665f
C980 VDD2.n57 VSUBS 0.027292f
C981 VDD2.n58 VSUBS 0.027292f
C982 VDD2.n59 VSUBS 0.014665f
C983 VDD2.n60 VSUBS 0.015528f
C984 VDD2.n61 VSUBS 0.034664f
C985 VDD2.n62 VSUBS 0.034664f
C986 VDD2.n63 VSUBS 0.015528f
C987 VDD2.n64 VSUBS 0.014665f
C988 VDD2.n65 VSUBS 0.027292f
C989 VDD2.n66 VSUBS 0.027292f
C990 VDD2.n67 VSUBS 0.014665f
C991 VDD2.n68 VSUBS 0.015528f
C992 VDD2.n69 VSUBS 0.034664f
C993 VDD2.n70 VSUBS 0.034664f
C994 VDD2.n71 VSUBS 0.034664f
C995 VDD2.n72 VSUBS 0.015528f
C996 VDD2.n73 VSUBS 0.014665f
C997 VDD2.n74 VSUBS 0.027292f
C998 VDD2.n75 VSUBS 0.027292f
C999 VDD2.n76 VSUBS 0.014665f
C1000 VDD2.n77 VSUBS 0.015097f
C1001 VDD2.n78 VSUBS 0.015097f
C1002 VDD2.n79 VSUBS 0.034664f
C1003 VDD2.n80 VSUBS 0.034664f
C1004 VDD2.n81 VSUBS 0.015528f
C1005 VDD2.n82 VSUBS 0.014665f
C1006 VDD2.n83 VSUBS 0.027292f
C1007 VDD2.n84 VSUBS 0.027292f
C1008 VDD2.n85 VSUBS 0.014665f
C1009 VDD2.n86 VSUBS 0.015528f
C1010 VDD2.n87 VSUBS 0.034664f
C1011 VDD2.n88 VSUBS 0.085105f
C1012 VDD2.n89 VSUBS 0.015528f
C1013 VDD2.n90 VSUBS 0.014665f
C1014 VDD2.n91 VSUBS 0.067558f
C1015 VDD2.n92 VSUBS 0.07139f
C1016 VDD2.t3 VSUBS 0.36491f
C1017 VDD2.t5 VSUBS 0.36491f
C1018 VDD2.n93 VSUBS 3.02621f
C1019 VDD2.n94 VSUBS 3.76127f
C1020 VDD2.n95 VSUBS 0.030337f
C1021 VDD2.n96 VSUBS 0.027292f
C1022 VDD2.n97 VSUBS 0.014665f
C1023 VDD2.n98 VSUBS 0.034664f
C1024 VDD2.n99 VSUBS 0.015528f
C1025 VDD2.n100 VSUBS 0.027292f
C1026 VDD2.n101 VSUBS 0.014665f
C1027 VDD2.n102 VSUBS 0.034664f
C1028 VDD2.n103 VSUBS 0.015528f
C1029 VDD2.n104 VSUBS 0.027292f
C1030 VDD2.n105 VSUBS 0.014665f
C1031 VDD2.n106 VSUBS 0.034664f
C1032 VDD2.n107 VSUBS 0.034664f
C1033 VDD2.n108 VSUBS 0.015528f
C1034 VDD2.n109 VSUBS 0.027292f
C1035 VDD2.n110 VSUBS 0.014665f
C1036 VDD2.n111 VSUBS 0.034664f
C1037 VDD2.n112 VSUBS 0.015528f
C1038 VDD2.n113 VSUBS 0.027292f
C1039 VDD2.n114 VSUBS 0.014665f
C1040 VDD2.n115 VSUBS 0.034664f
C1041 VDD2.n116 VSUBS 0.015528f
C1042 VDD2.n117 VSUBS 0.027292f
C1043 VDD2.n118 VSUBS 0.014665f
C1044 VDD2.n119 VSUBS 0.034664f
C1045 VDD2.n120 VSUBS 0.015528f
C1046 VDD2.n121 VSUBS 0.027292f
C1047 VDD2.n122 VSUBS 0.014665f
C1048 VDD2.n123 VSUBS 0.034664f
C1049 VDD2.n124 VSUBS 0.015528f
C1050 VDD2.n125 VSUBS 0.207839f
C1051 VDD2.t4 VSUBS 0.074338f
C1052 VDD2.n126 VSUBS 0.025998f
C1053 VDD2.n127 VSUBS 0.022051f
C1054 VDD2.n128 VSUBS 0.014665f
C1055 VDD2.n129 VSUBS 1.98052f
C1056 VDD2.n130 VSUBS 0.027292f
C1057 VDD2.n131 VSUBS 0.014665f
C1058 VDD2.n132 VSUBS 0.015528f
C1059 VDD2.n133 VSUBS 0.034664f
C1060 VDD2.n134 VSUBS 0.034664f
C1061 VDD2.n135 VSUBS 0.015528f
C1062 VDD2.n136 VSUBS 0.014665f
C1063 VDD2.n137 VSUBS 0.027292f
C1064 VDD2.n138 VSUBS 0.027292f
C1065 VDD2.n139 VSUBS 0.014665f
C1066 VDD2.n140 VSUBS 0.015528f
C1067 VDD2.n141 VSUBS 0.034664f
C1068 VDD2.n142 VSUBS 0.034664f
C1069 VDD2.n143 VSUBS 0.015528f
C1070 VDD2.n144 VSUBS 0.014665f
C1071 VDD2.n145 VSUBS 0.027292f
C1072 VDD2.n146 VSUBS 0.027292f
C1073 VDD2.n147 VSUBS 0.014665f
C1074 VDD2.n148 VSUBS 0.015528f
C1075 VDD2.n149 VSUBS 0.034664f
C1076 VDD2.n150 VSUBS 0.034664f
C1077 VDD2.n151 VSUBS 0.015528f
C1078 VDD2.n152 VSUBS 0.014665f
C1079 VDD2.n153 VSUBS 0.027292f
C1080 VDD2.n154 VSUBS 0.027292f
C1081 VDD2.n155 VSUBS 0.014665f
C1082 VDD2.n156 VSUBS 0.015528f
C1083 VDD2.n157 VSUBS 0.034664f
C1084 VDD2.n158 VSUBS 0.034664f
C1085 VDD2.n159 VSUBS 0.015528f
C1086 VDD2.n160 VSUBS 0.014665f
C1087 VDD2.n161 VSUBS 0.027292f
C1088 VDD2.n162 VSUBS 0.027292f
C1089 VDD2.n163 VSUBS 0.014665f
C1090 VDD2.n164 VSUBS 0.015528f
C1091 VDD2.n165 VSUBS 0.034664f
C1092 VDD2.n166 VSUBS 0.034664f
C1093 VDD2.n167 VSUBS 0.015528f
C1094 VDD2.n168 VSUBS 0.014665f
C1095 VDD2.n169 VSUBS 0.027292f
C1096 VDD2.n170 VSUBS 0.027292f
C1097 VDD2.n171 VSUBS 0.014665f
C1098 VDD2.n172 VSUBS 0.015097f
C1099 VDD2.n173 VSUBS 0.015097f
C1100 VDD2.n174 VSUBS 0.034664f
C1101 VDD2.n175 VSUBS 0.034664f
C1102 VDD2.n176 VSUBS 0.015528f
C1103 VDD2.n177 VSUBS 0.014665f
C1104 VDD2.n178 VSUBS 0.027292f
C1105 VDD2.n179 VSUBS 0.027292f
C1106 VDD2.n180 VSUBS 0.014665f
C1107 VDD2.n181 VSUBS 0.015528f
C1108 VDD2.n182 VSUBS 0.034664f
C1109 VDD2.n183 VSUBS 0.085105f
C1110 VDD2.n184 VSUBS 0.015528f
C1111 VDD2.n185 VSUBS 0.014665f
C1112 VDD2.n186 VSUBS 0.067558f
C1113 VDD2.n187 VSUBS 0.061796f
C1114 VDD2.n188 VSUBS 3.33726f
C1115 VDD2.t1 VSUBS 0.36491f
C1116 VDD2.t2 VSUBS 0.36491f
C1117 VDD2.n189 VSUBS 3.02617f
C1118 VN.t0 VSUBS 3.57914f
C1119 VN.n0 VSUBS 1.33837f
C1120 VN.n1 VSUBS 0.025412f
C1121 VN.n2 VSUBS 0.032266f
C1122 VN.n3 VSUBS 0.289176f
C1123 VN.t2 VSUBS 3.57914f
C1124 VN.t5 VSUBS 3.85979f
C1125 VN.n4 VSUBS 1.27912f
C1126 VN.n5 VSUBS 1.33559f
C1127 VN.n6 VSUBS 0.047599f
C1128 VN.n7 VSUBS 0.047599f
C1129 VN.n8 VSUBS 0.025412f
C1130 VN.n9 VSUBS 0.025412f
C1131 VN.n10 VSUBS 0.025412f
C1132 VN.n11 VSUBS 0.04225f
C1133 VN.n12 VSUBS 0.047599f
C1134 VN.n13 VSUBS 0.041018f
C1135 VN.n14 VSUBS 0.041021f
C1136 VN.n15 VSUBS 0.05582f
C1137 VN.t1 VSUBS 3.57914f
C1138 VN.n16 VSUBS 1.33837f
C1139 VN.n17 VSUBS 0.025412f
C1140 VN.n18 VSUBS 0.032266f
C1141 VN.n19 VSUBS 0.289176f
C1142 VN.t4 VSUBS 3.57914f
C1143 VN.t3 VSUBS 3.85979f
C1144 VN.n20 VSUBS 1.27912f
C1145 VN.n21 VSUBS 1.33559f
C1146 VN.n22 VSUBS 0.047599f
C1147 VN.n23 VSUBS 0.047599f
C1148 VN.n24 VSUBS 0.025412f
C1149 VN.n25 VSUBS 0.025412f
C1150 VN.n26 VSUBS 0.025412f
C1151 VN.n27 VSUBS 0.04225f
C1152 VN.n28 VSUBS 0.047599f
C1153 VN.n29 VSUBS 0.041018f
C1154 VN.n30 VSUBS 0.041021f
C1155 VN.n31 VSUBS 1.62254f
C1156 VDD1.n0 VSUBS 0.030213f
C1157 VDD1.n1 VSUBS 0.027181f
C1158 VDD1.n2 VSUBS 0.014606f
C1159 VDD1.n3 VSUBS 0.034523f
C1160 VDD1.n4 VSUBS 0.015465f
C1161 VDD1.n5 VSUBS 0.027181f
C1162 VDD1.n6 VSUBS 0.014606f
C1163 VDD1.n7 VSUBS 0.034523f
C1164 VDD1.n8 VSUBS 0.015465f
C1165 VDD1.n9 VSUBS 0.027181f
C1166 VDD1.n10 VSUBS 0.014606f
C1167 VDD1.n11 VSUBS 0.034523f
C1168 VDD1.n12 VSUBS 0.034523f
C1169 VDD1.n13 VSUBS 0.015465f
C1170 VDD1.n14 VSUBS 0.027181f
C1171 VDD1.n15 VSUBS 0.014606f
C1172 VDD1.n16 VSUBS 0.034523f
C1173 VDD1.n17 VSUBS 0.015465f
C1174 VDD1.n18 VSUBS 0.027181f
C1175 VDD1.n19 VSUBS 0.014606f
C1176 VDD1.n20 VSUBS 0.034523f
C1177 VDD1.n21 VSUBS 0.015465f
C1178 VDD1.n22 VSUBS 0.027181f
C1179 VDD1.n23 VSUBS 0.014606f
C1180 VDD1.n24 VSUBS 0.034523f
C1181 VDD1.n25 VSUBS 0.015465f
C1182 VDD1.n26 VSUBS 0.027181f
C1183 VDD1.n27 VSUBS 0.014606f
C1184 VDD1.n28 VSUBS 0.034523f
C1185 VDD1.n29 VSUBS 0.015465f
C1186 VDD1.n30 VSUBS 0.206994f
C1187 VDD1.t1 VSUBS 0.074036f
C1188 VDD1.n31 VSUBS 0.025892f
C1189 VDD1.n32 VSUBS 0.021962f
C1190 VDD1.n33 VSUBS 0.014606f
C1191 VDD1.n34 VSUBS 1.97247f
C1192 VDD1.n35 VSUBS 0.027181f
C1193 VDD1.n36 VSUBS 0.014606f
C1194 VDD1.n37 VSUBS 0.015465f
C1195 VDD1.n38 VSUBS 0.034523f
C1196 VDD1.n39 VSUBS 0.034523f
C1197 VDD1.n40 VSUBS 0.015465f
C1198 VDD1.n41 VSUBS 0.014606f
C1199 VDD1.n42 VSUBS 0.027181f
C1200 VDD1.n43 VSUBS 0.027181f
C1201 VDD1.n44 VSUBS 0.014606f
C1202 VDD1.n45 VSUBS 0.015465f
C1203 VDD1.n46 VSUBS 0.034523f
C1204 VDD1.n47 VSUBS 0.034523f
C1205 VDD1.n48 VSUBS 0.015465f
C1206 VDD1.n49 VSUBS 0.014606f
C1207 VDD1.n50 VSUBS 0.027181f
C1208 VDD1.n51 VSUBS 0.027181f
C1209 VDD1.n52 VSUBS 0.014606f
C1210 VDD1.n53 VSUBS 0.015465f
C1211 VDD1.n54 VSUBS 0.034523f
C1212 VDD1.n55 VSUBS 0.034523f
C1213 VDD1.n56 VSUBS 0.015465f
C1214 VDD1.n57 VSUBS 0.014606f
C1215 VDD1.n58 VSUBS 0.027181f
C1216 VDD1.n59 VSUBS 0.027181f
C1217 VDD1.n60 VSUBS 0.014606f
C1218 VDD1.n61 VSUBS 0.015465f
C1219 VDD1.n62 VSUBS 0.034523f
C1220 VDD1.n63 VSUBS 0.034523f
C1221 VDD1.n64 VSUBS 0.015465f
C1222 VDD1.n65 VSUBS 0.014606f
C1223 VDD1.n66 VSUBS 0.027181f
C1224 VDD1.n67 VSUBS 0.027181f
C1225 VDD1.n68 VSUBS 0.014606f
C1226 VDD1.n69 VSUBS 0.015465f
C1227 VDD1.n70 VSUBS 0.034523f
C1228 VDD1.n71 VSUBS 0.034523f
C1229 VDD1.n72 VSUBS 0.015465f
C1230 VDD1.n73 VSUBS 0.014606f
C1231 VDD1.n74 VSUBS 0.027181f
C1232 VDD1.n75 VSUBS 0.027181f
C1233 VDD1.n76 VSUBS 0.014606f
C1234 VDD1.n77 VSUBS 0.015035f
C1235 VDD1.n78 VSUBS 0.015035f
C1236 VDD1.n79 VSUBS 0.034523f
C1237 VDD1.n80 VSUBS 0.034523f
C1238 VDD1.n81 VSUBS 0.015465f
C1239 VDD1.n82 VSUBS 0.014606f
C1240 VDD1.n83 VSUBS 0.027181f
C1241 VDD1.n84 VSUBS 0.027181f
C1242 VDD1.n85 VSUBS 0.014606f
C1243 VDD1.n86 VSUBS 0.015465f
C1244 VDD1.n87 VSUBS 0.034523f
C1245 VDD1.n88 VSUBS 0.084759f
C1246 VDD1.n89 VSUBS 0.015465f
C1247 VDD1.n90 VSUBS 0.014606f
C1248 VDD1.n91 VSUBS 0.067283f
C1249 VDD1.n92 VSUBS 0.071994f
C1250 VDD1.n93 VSUBS 0.030213f
C1251 VDD1.n94 VSUBS 0.027181f
C1252 VDD1.n95 VSUBS 0.014606f
C1253 VDD1.n96 VSUBS 0.034523f
C1254 VDD1.n97 VSUBS 0.015465f
C1255 VDD1.n98 VSUBS 0.027181f
C1256 VDD1.n99 VSUBS 0.014606f
C1257 VDD1.n100 VSUBS 0.034523f
C1258 VDD1.n101 VSUBS 0.015465f
C1259 VDD1.n102 VSUBS 0.027181f
C1260 VDD1.n103 VSUBS 0.014606f
C1261 VDD1.n104 VSUBS 0.034523f
C1262 VDD1.n105 VSUBS 0.015465f
C1263 VDD1.n106 VSUBS 0.027181f
C1264 VDD1.n107 VSUBS 0.014606f
C1265 VDD1.n108 VSUBS 0.034523f
C1266 VDD1.n109 VSUBS 0.015465f
C1267 VDD1.n110 VSUBS 0.027181f
C1268 VDD1.n111 VSUBS 0.014606f
C1269 VDD1.n112 VSUBS 0.034523f
C1270 VDD1.n113 VSUBS 0.015465f
C1271 VDD1.n114 VSUBS 0.027181f
C1272 VDD1.n115 VSUBS 0.014606f
C1273 VDD1.n116 VSUBS 0.034523f
C1274 VDD1.n117 VSUBS 0.015465f
C1275 VDD1.n118 VSUBS 0.027181f
C1276 VDD1.n119 VSUBS 0.014606f
C1277 VDD1.n120 VSUBS 0.034523f
C1278 VDD1.n121 VSUBS 0.015465f
C1279 VDD1.n122 VSUBS 0.206994f
C1280 VDD1.t4 VSUBS 0.074036f
C1281 VDD1.n123 VSUBS 0.025892f
C1282 VDD1.n124 VSUBS 0.021962f
C1283 VDD1.n125 VSUBS 0.014606f
C1284 VDD1.n126 VSUBS 1.97247f
C1285 VDD1.n127 VSUBS 0.027181f
C1286 VDD1.n128 VSUBS 0.014606f
C1287 VDD1.n129 VSUBS 0.015465f
C1288 VDD1.n130 VSUBS 0.034523f
C1289 VDD1.n131 VSUBS 0.034523f
C1290 VDD1.n132 VSUBS 0.015465f
C1291 VDD1.n133 VSUBS 0.014606f
C1292 VDD1.n134 VSUBS 0.027181f
C1293 VDD1.n135 VSUBS 0.027181f
C1294 VDD1.n136 VSUBS 0.014606f
C1295 VDD1.n137 VSUBS 0.015465f
C1296 VDD1.n138 VSUBS 0.034523f
C1297 VDD1.n139 VSUBS 0.034523f
C1298 VDD1.n140 VSUBS 0.015465f
C1299 VDD1.n141 VSUBS 0.014606f
C1300 VDD1.n142 VSUBS 0.027181f
C1301 VDD1.n143 VSUBS 0.027181f
C1302 VDD1.n144 VSUBS 0.014606f
C1303 VDD1.n145 VSUBS 0.015465f
C1304 VDD1.n146 VSUBS 0.034523f
C1305 VDD1.n147 VSUBS 0.034523f
C1306 VDD1.n148 VSUBS 0.015465f
C1307 VDD1.n149 VSUBS 0.014606f
C1308 VDD1.n150 VSUBS 0.027181f
C1309 VDD1.n151 VSUBS 0.027181f
C1310 VDD1.n152 VSUBS 0.014606f
C1311 VDD1.n153 VSUBS 0.015465f
C1312 VDD1.n154 VSUBS 0.034523f
C1313 VDD1.n155 VSUBS 0.034523f
C1314 VDD1.n156 VSUBS 0.015465f
C1315 VDD1.n157 VSUBS 0.014606f
C1316 VDD1.n158 VSUBS 0.027181f
C1317 VDD1.n159 VSUBS 0.027181f
C1318 VDD1.n160 VSUBS 0.014606f
C1319 VDD1.n161 VSUBS 0.015465f
C1320 VDD1.n162 VSUBS 0.034523f
C1321 VDD1.n163 VSUBS 0.034523f
C1322 VDD1.n164 VSUBS 0.034523f
C1323 VDD1.n165 VSUBS 0.015465f
C1324 VDD1.n166 VSUBS 0.014606f
C1325 VDD1.n167 VSUBS 0.027181f
C1326 VDD1.n168 VSUBS 0.027181f
C1327 VDD1.n169 VSUBS 0.014606f
C1328 VDD1.n170 VSUBS 0.015035f
C1329 VDD1.n171 VSUBS 0.015035f
C1330 VDD1.n172 VSUBS 0.034523f
C1331 VDD1.n173 VSUBS 0.034523f
C1332 VDD1.n174 VSUBS 0.015465f
C1333 VDD1.n175 VSUBS 0.014606f
C1334 VDD1.n176 VSUBS 0.027181f
C1335 VDD1.n177 VSUBS 0.027181f
C1336 VDD1.n178 VSUBS 0.014606f
C1337 VDD1.n179 VSUBS 0.015465f
C1338 VDD1.n180 VSUBS 0.034523f
C1339 VDD1.n181 VSUBS 0.084759f
C1340 VDD1.n182 VSUBS 0.015465f
C1341 VDD1.n183 VSUBS 0.014606f
C1342 VDD1.n184 VSUBS 0.067283f
C1343 VDD1.n185 VSUBS 0.0711f
C1344 VDD1.t3 VSUBS 0.363427f
C1345 VDD1.t0 VSUBS 0.363427f
C1346 VDD1.n186 VSUBS 3.01391f
C1347 VDD1.n187 VSUBS 3.89721f
C1348 VDD1.t2 VSUBS 0.363427f
C1349 VDD1.t5 VSUBS 0.363427f
C1350 VDD1.n188 VSUBS 3.0061f
C1351 VDD1.n189 VSUBS 3.86669f
C1352 VTAIL.t5 VSUBS 0.374545f
C1353 VTAIL.t3 VSUBS 0.374545f
C1354 VTAIL.n0 VSUBS 2.93694f
C1355 VTAIL.n1 VSUBS 0.90387f
C1356 VTAIL.n2 VSUBS 0.031137f
C1357 VTAIL.n3 VSUBS 0.028012f
C1358 VTAIL.n4 VSUBS 0.015053f
C1359 VTAIL.n5 VSUBS 0.035579f
C1360 VTAIL.n6 VSUBS 0.015938f
C1361 VTAIL.n7 VSUBS 0.028012f
C1362 VTAIL.n8 VSUBS 0.015053f
C1363 VTAIL.n9 VSUBS 0.035579f
C1364 VTAIL.n10 VSUBS 0.015938f
C1365 VTAIL.n11 VSUBS 0.028012f
C1366 VTAIL.n12 VSUBS 0.015053f
C1367 VTAIL.n13 VSUBS 0.035579f
C1368 VTAIL.n14 VSUBS 0.015938f
C1369 VTAIL.n15 VSUBS 0.028012f
C1370 VTAIL.n16 VSUBS 0.015053f
C1371 VTAIL.n17 VSUBS 0.035579f
C1372 VTAIL.n18 VSUBS 0.015938f
C1373 VTAIL.n19 VSUBS 0.028012f
C1374 VTAIL.n20 VSUBS 0.015053f
C1375 VTAIL.n21 VSUBS 0.035579f
C1376 VTAIL.n22 VSUBS 0.015938f
C1377 VTAIL.n23 VSUBS 0.028012f
C1378 VTAIL.n24 VSUBS 0.015053f
C1379 VTAIL.n25 VSUBS 0.035579f
C1380 VTAIL.n26 VSUBS 0.015938f
C1381 VTAIL.n27 VSUBS 0.028012f
C1382 VTAIL.n28 VSUBS 0.015053f
C1383 VTAIL.n29 VSUBS 0.035579f
C1384 VTAIL.n30 VSUBS 0.015938f
C1385 VTAIL.n31 VSUBS 0.213327f
C1386 VTAIL.t6 VSUBS 0.076301f
C1387 VTAIL.n32 VSUBS 0.026684f
C1388 VTAIL.n33 VSUBS 0.022634f
C1389 VTAIL.n34 VSUBS 0.015053f
C1390 VTAIL.n35 VSUBS 2.03281f
C1391 VTAIL.n36 VSUBS 0.028012f
C1392 VTAIL.n37 VSUBS 0.015053f
C1393 VTAIL.n38 VSUBS 0.015938f
C1394 VTAIL.n39 VSUBS 0.035579f
C1395 VTAIL.n40 VSUBS 0.035579f
C1396 VTAIL.n41 VSUBS 0.015938f
C1397 VTAIL.n42 VSUBS 0.015053f
C1398 VTAIL.n43 VSUBS 0.028012f
C1399 VTAIL.n44 VSUBS 0.028012f
C1400 VTAIL.n45 VSUBS 0.015053f
C1401 VTAIL.n46 VSUBS 0.015938f
C1402 VTAIL.n47 VSUBS 0.035579f
C1403 VTAIL.n48 VSUBS 0.035579f
C1404 VTAIL.n49 VSUBS 0.015938f
C1405 VTAIL.n50 VSUBS 0.015053f
C1406 VTAIL.n51 VSUBS 0.028012f
C1407 VTAIL.n52 VSUBS 0.028012f
C1408 VTAIL.n53 VSUBS 0.015053f
C1409 VTAIL.n54 VSUBS 0.015938f
C1410 VTAIL.n55 VSUBS 0.035579f
C1411 VTAIL.n56 VSUBS 0.035579f
C1412 VTAIL.n57 VSUBS 0.015938f
C1413 VTAIL.n58 VSUBS 0.015053f
C1414 VTAIL.n59 VSUBS 0.028012f
C1415 VTAIL.n60 VSUBS 0.028012f
C1416 VTAIL.n61 VSUBS 0.015053f
C1417 VTAIL.n62 VSUBS 0.015938f
C1418 VTAIL.n63 VSUBS 0.035579f
C1419 VTAIL.n64 VSUBS 0.035579f
C1420 VTAIL.n65 VSUBS 0.015938f
C1421 VTAIL.n66 VSUBS 0.015053f
C1422 VTAIL.n67 VSUBS 0.028012f
C1423 VTAIL.n68 VSUBS 0.028012f
C1424 VTAIL.n69 VSUBS 0.015053f
C1425 VTAIL.n70 VSUBS 0.015938f
C1426 VTAIL.n71 VSUBS 0.035579f
C1427 VTAIL.n72 VSUBS 0.035579f
C1428 VTAIL.n73 VSUBS 0.035579f
C1429 VTAIL.n74 VSUBS 0.015938f
C1430 VTAIL.n75 VSUBS 0.015053f
C1431 VTAIL.n76 VSUBS 0.028012f
C1432 VTAIL.n77 VSUBS 0.028012f
C1433 VTAIL.n78 VSUBS 0.015053f
C1434 VTAIL.n79 VSUBS 0.015495f
C1435 VTAIL.n80 VSUBS 0.015495f
C1436 VTAIL.n81 VSUBS 0.035579f
C1437 VTAIL.n82 VSUBS 0.035579f
C1438 VTAIL.n83 VSUBS 0.015938f
C1439 VTAIL.n84 VSUBS 0.015053f
C1440 VTAIL.n85 VSUBS 0.028012f
C1441 VTAIL.n86 VSUBS 0.028012f
C1442 VTAIL.n87 VSUBS 0.015053f
C1443 VTAIL.n88 VSUBS 0.015938f
C1444 VTAIL.n89 VSUBS 0.035579f
C1445 VTAIL.n90 VSUBS 0.087352f
C1446 VTAIL.n91 VSUBS 0.015938f
C1447 VTAIL.n92 VSUBS 0.015053f
C1448 VTAIL.n93 VSUBS 0.069341f
C1449 VTAIL.n94 VSUBS 0.044119f
C1450 VTAIL.n95 VSUBS 0.461102f
C1451 VTAIL.t8 VSUBS 0.374545f
C1452 VTAIL.t7 VSUBS 0.374545f
C1453 VTAIL.n96 VSUBS 2.93694f
C1454 VTAIL.n97 VSUBS 3.14157f
C1455 VTAIL.t0 VSUBS 0.374545f
C1456 VTAIL.t1 VSUBS 0.374545f
C1457 VTAIL.n98 VSUBS 2.93696f
C1458 VTAIL.n99 VSUBS 3.14155f
C1459 VTAIL.n100 VSUBS 0.031137f
C1460 VTAIL.n101 VSUBS 0.028012f
C1461 VTAIL.n102 VSUBS 0.015053f
C1462 VTAIL.n103 VSUBS 0.035579f
C1463 VTAIL.n104 VSUBS 0.015938f
C1464 VTAIL.n105 VSUBS 0.028012f
C1465 VTAIL.n106 VSUBS 0.015053f
C1466 VTAIL.n107 VSUBS 0.035579f
C1467 VTAIL.n108 VSUBS 0.015938f
C1468 VTAIL.n109 VSUBS 0.028012f
C1469 VTAIL.n110 VSUBS 0.015053f
C1470 VTAIL.n111 VSUBS 0.035579f
C1471 VTAIL.n112 VSUBS 0.035579f
C1472 VTAIL.n113 VSUBS 0.015938f
C1473 VTAIL.n114 VSUBS 0.028012f
C1474 VTAIL.n115 VSUBS 0.015053f
C1475 VTAIL.n116 VSUBS 0.035579f
C1476 VTAIL.n117 VSUBS 0.015938f
C1477 VTAIL.n118 VSUBS 0.028012f
C1478 VTAIL.n119 VSUBS 0.015053f
C1479 VTAIL.n120 VSUBS 0.035579f
C1480 VTAIL.n121 VSUBS 0.015938f
C1481 VTAIL.n122 VSUBS 0.028012f
C1482 VTAIL.n123 VSUBS 0.015053f
C1483 VTAIL.n124 VSUBS 0.035579f
C1484 VTAIL.n125 VSUBS 0.015938f
C1485 VTAIL.n126 VSUBS 0.028012f
C1486 VTAIL.n127 VSUBS 0.015053f
C1487 VTAIL.n128 VSUBS 0.035579f
C1488 VTAIL.n129 VSUBS 0.015938f
C1489 VTAIL.n130 VSUBS 0.213327f
C1490 VTAIL.t2 VSUBS 0.076301f
C1491 VTAIL.n131 VSUBS 0.026684f
C1492 VTAIL.n132 VSUBS 0.022634f
C1493 VTAIL.n133 VSUBS 0.015053f
C1494 VTAIL.n134 VSUBS 2.03281f
C1495 VTAIL.n135 VSUBS 0.028012f
C1496 VTAIL.n136 VSUBS 0.015053f
C1497 VTAIL.n137 VSUBS 0.015938f
C1498 VTAIL.n138 VSUBS 0.035579f
C1499 VTAIL.n139 VSUBS 0.035579f
C1500 VTAIL.n140 VSUBS 0.015938f
C1501 VTAIL.n141 VSUBS 0.015053f
C1502 VTAIL.n142 VSUBS 0.028012f
C1503 VTAIL.n143 VSUBS 0.028012f
C1504 VTAIL.n144 VSUBS 0.015053f
C1505 VTAIL.n145 VSUBS 0.015938f
C1506 VTAIL.n146 VSUBS 0.035579f
C1507 VTAIL.n147 VSUBS 0.035579f
C1508 VTAIL.n148 VSUBS 0.015938f
C1509 VTAIL.n149 VSUBS 0.015053f
C1510 VTAIL.n150 VSUBS 0.028012f
C1511 VTAIL.n151 VSUBS 0.028012f
C1512 VTAIL.n152 VSUBS 0.015053f
C1513 VTAIL.n153 VSUBS 0.015938f
C1514 VTAIL.n154 VSUBS 0.035579f
C1515 VTAIL.n155 VSUBS 0.035579f
C1516 VTAIL.n156 VSUBS 0.015938f
C1517 VTAIL.n157 VSUBS 0.015053f
C1518 VTAIL.n158 VSUBS 0.028012f
C1519 VTAIL.n159 VSUBS 0.028012f
C1520 VTAIL.n160 VSUBS 0.015053f
C1521 VTAIL.n161 VSUBS 0.015938f
C1522 VTAIL.n162 VSUBS 0.035579f
C1523 VTAIL.n163 VSUBS 0.035579f
C1524 VTAIL.n164 VSUBS 0.015938f
C1525 VTAIL.n165 VSUBS 0.015053f
C1526 VTAIL.n166 VSUBS 0.028012f
C1527 VTAIL.n167 VSUBS 0.028012f
C1528 VTAIL.n168 VSUBS 0.015053f
C1529 VTAIL.n169 VSUBS 0.015938f
C1530 VTAIL.n170 VSUBS 0.035579f
C1531 VTAIL.n171 VSUBS 0.035579f
C1532 VTAIL.n172 VSUBS 0.015938f
C1533 VTAIL.n173 VSUBS 0.015053f
C1534 VTAIL.n174 VSUBS 0.028012f
C1535 VTAIL.n175 VSUBS 0.028012f
C1536 VTAIL.n176 VSUBS 0.015053f
C1537 VTAIL.n177 VSUBS 0.015495f
C1538 VTAIL.n178 VSUBS 0.015495f
C1539 VTAIL.n179 VSUBS 0.035579f
C1540 VTAIL.n180 VSUBS 0.035579f
C1541 VTAIL.n181 VSUBS 0.015938f
C1542 VTAIL.n182 VSUBS 0.015053f
C1543 VTAIL.n183 VSUBS 0.028012f
C1544 VTAIL.n184 VSUBS 0.028012f
C1545 VTAIL.n185 VSUBS 0.015053f
C1546 VTAIL.n186 VSUBS 0.015938f
C1547 VTAIL.n187 VSUBS 0.035579f
C1548 VTAIL.n188 VSUBS 0.087352f
C1549 VTAIL.n189 VSUBS 0.015938f
C1550 VTAIL.n190 VSUBS 0.015053f
C1551 VTAIL.n191 VSUBS 0.069341f
C1552 VTAIL.n192 VSUBS 0.044119f
C1553 VTAIL.n193 VSUBS 0.461102f
C1554 VTAIL.t10 VSUBS 0.374545f
C1555 VTAIL.t11 VSUBS 0.374545f
C1556 VTAIL.n194 VSUBS 2.93696f
C1557 VTAIL.n195 VSUBS 1.09469f
C1558 VTAIL.n196 VSUBS 0.031137f
C1559 VTAIL.n197 VSUBS 0.028012f
C1560 VTAIL.n198 VSUBS 0.015053f
C1561 VTAIL.n199 VSUBS 0.035579f
C1562 VTAIL.n200 VSUBS 0.015938f
C1563 VTAIL.n201 VSUBS 0.028012f
C1564 VTAIL.n202 VSUBS 0.015053f
C1565 VTAIL.n203 VSUBS 0.035579f
C1566 VTAIL.n204 VSUBS 0.015938f
C1567 VTAIL.n205 VSUBS 0.028012f
C1568 VTAIL.n206 VSUBS 0.015053f
C1569 VTAIL.n207 VSUBS 0.035579f
C1570 VTAIL.n208 VSUBS 0.035579f
C1571 VTAIL.n209 VSUBS 0.015938f
C1572 VTAIL.n210 VSUBS 0.028012f
C1573 VTAIL.n211 VSUBS 0.015053f
C1574 VTAIL.n212 VSUBS 0.035579f
C1575 VTAIL.n213 VSUBS 0.015938f
C1576 VTAIL.n214 VSUBS 0.028012f
C1577 VTAIL.n215 VSUBS 0.015053f
C1578 VTAIL.n216 VSUBS 0.035579f
C1579 VTAIL.n217 VSUBS 0.015938f
C1580 VTAIL.n218 VSUBS 0.028012f
C1581 VTAIL.n219 VSUBS 0.015053f
C1582 VTAIL.n220 VSUBS 0.035579f
C1583 VTAIL.n221 VSUBS 0.015938f
C1584 VTAIL.n222 VSUBS 0.028012f
C1585 VTAIL.n223 VSUBS 0.015053f
C1586 VTAIL.n224 VSUBS 0.035579f
C1587 VTAIL.n225 VSUBS 0.015938f
C1588 VTAIL.n226 VSUBS 0.213327f
C1589 VTAIL.t9 VSUBS 0.076301f
C1590 VTAIL.n227 VSUBS 0.026684f
C1591 VTAIL.n228 VSUBS 0.022634f
C1592 VTAIL.n229 VSUBS 0.015053f
C1593 VTAIL.n230 VSUBS 2.03281f
C1594 VTAIL.n231 VSUBS 0.028012f
C1595 VTAIL.n232 VSUBS 0.015053f
C1596 VTAIL.n233 VSUBS 0.015938f
C1597 VTAIL.n234 VSUBS 0.035579f
C1598 VTAIL.n235 VSUBS 0.035579f
C1599 VTAIL.n236 VSUBS 0.015938f
C1600 VTAIL.n237 VSUBS 0.015053f
C1601 VTAIL.n238 VSUBS 0.028012f
C1602 VTAIL.n239 VSUBS 0.028012f
C1603 VTAIL.n240 VSUBS 0.015053f
C1604 VTAIL.n241 VSUBS 0.015938f
C1605 VTAIL.n242 VSUBS 0.035579f
C1606 VTAIL.n243 VSUBS 0.035579f
C1607 VTAIL.n244 VSUBS 0.015938f
C1608 VTAIL.n245 VSUBS 0.015053f
C1609 VTAIL.n246 VSUBS 0.028012f
C1610 VTAIL.n247 VSUBS 0.028012f
C1611 VTAIL.n248 VSUBS 0.015053f
C1612 VTAIL.n249 VSUBS 0.015938f
C1613 VTAIL.n250 VSUBS 0.035579f
C1614 VTAIL.n251 VSUBS 0.035579f
C1615 VTAIL.n252 VSUBS 0.015938f
C1616 VTAIL.n253 VSUBS 0.015053f
C1617 VTAIL.n254 VSUBS 0.028012f
C1618 VTAIL.n255 VSUBS 0.028012f
C1619 VTAIL.n256 VSUBS 0.015053f
C1620 VTAIL.n257 VSUBS 0.015938f
C1621 VTAIL.n258 VSUBS 0.035579f
C1622 VTAIL.n259 VSUBS 0.035579f
C1623 VTAIL.n260 VSUBS 0.015938f
C1624 VTAIL.n261 VSUBS 0.015053f
C1625 VTAIL.n262 VSUBS 0.028012f
C1626 VTAIL.n263 VSUBS 0.028012f
C1627 VTAIL.n264 VSUBS 0.015053f
C1628 VTAIL.n265 VSUBS 0.015938f
C1629 VTAIL.n266 VSUBS 0.035579f
C1630 VTAIL.n267 VSUBS 0.035579f
C1631 VTAIL.n268 VSUBS 0.015938f
C1632 VTAIL.n269 VSUBS 0.015053f
C1633 VTAIL.n270 VSUBS 0.028012f
C1634 VTAIL.n271 VSUBS 0.028012f
C1635 VTAIL.n272 VSUBS 0.015053f
C1636 VTAIL.n273 VSUBS 0.015495f
C1637 VTAIL.n274 VSUBS 0.015495f
C1638 VTAIL.n275 VSUBS 0.035579f
C1639 VTAIL.n276 VSUBS 0.035579f
C1640 VTAIL.n277 VSUBS 0.015938f
C1641 VTAIL.n278 VSUBS 0.015053f
C1642 VTAIL.n279 VSUBS 0.028012f
C1643 VTAIL.n280 VSUBS 0.028012f
C1644 VTAIL.n281 VSUBS 0.015053f
C1645 VTAIL.n282 VSUBS 0.015938f
C1646 VTAIL.n283 VSUBS 0.035579f
C1647 VTAIL.n284 VSUBS 0.087352f
C1648 VTAIL.n285 VSUBS 0.015938f
C1649 VTAIL.n286 VSUBS 0.015053f
C1650 VTAIL.n287 VSUBS 0.069341f
C1651 VTAIL.n288 VSUBS 0.044119f
C1652 VTAIL.n289 VSUBS 2.24652f
C1653 VTAIL.n290 VSUBS 0.031137f
C1654 VTAIL.n291 VSUBS 0.028012f
C1655 VTAIL.n292 VSUBS 0.015053f
C1656 VTAIL.n293 VSUBS 0.035579f
C1657 VTAIL.n294 VSUBS 0.015938f
C1658 VTAIL.n295 VSUBS 0.028012f
C1659 VTAIL.n296 VSUBS 0.015053f
C1660 VTAIL.n297 VSUBS 0.035579f
C1661 VTAIL.n298 VSUBS 0.015938f
C1662 VTAIL.n299 VSUBS 0.028012f
C1663 VTAIL.n300 VSUBS 0.015053f
C1664 VTAIL.n301 VSUBS 0.035579f
C1665 VTAIL.n302 VSUBS 0.015938f
C1666 VTAIL.n303 VSUBS 0.028012f
C1667 VTAIL.n304 VSUBS 0.015053f
C1668 VTAIL.n305 VSUBS 0.035579f
C1669 VTAIL.n306 VSUBS 0.015938f
C1670 VTAIL.n307 VSUBS 0.028012f
C1671 VTAIL.n308 VSUBS 0.015053f
C1672 VTAIL.n309 VSUBS 0.035579f
C1673 VTAIL.n310 VSUBS 0.015938f
C1674 VTAIL.n311 VSUBS 0.028012f
C1675 VTAIL.n312 VSUBS 0.015053f
C1676 VTAIL.n313 VSUBS 0.035579f
C1677 VTAIL.n314 VSUBS 0.015938f
C1678 VTAIL.n315 VSUBS 0.028012f
C1679 VTAIL.n316 VSUBS 0.015053f
C1680 VTAIL.n317 VSUBS 0.035579f
C1681 VTAIL.n318 VSUBS 0.015938f
C1682 VTAIL.n319 VSUBS 0.213327f
C1683 VTAIL.t4 VSUBS 0.076301f
C1684 VTAIL.n320 VSUBS 0.026684f
C1685 VTAIL.n321 VSUBS 0.022634f
C1686 VTAIL.n322 VSUBS 0.015053f
C1687 VTAIL.n323 VSUBS 2.03281f
C1688 VTAIL.n324 VSUBS 0.028012f
C1689 VTAIL.n325 VSUBS 0.015053f
C1690 VTAIL.n326 VSUBS 0.015938f
C1691 VTAIL.n327 VSUBS 0.035579f
C1692 VTAIL.n328 VSUBS 0.035579f
C1693 VTAIL.n329 VSUBS 0.015938f
C1694 VTAIL.n330 VSUBS 0.015053f
C1695 VTAIL.n331 VSUBS 0.028012f
C1696 VTAIL.n332 VSUBS 0.028012f
C1697 VTAIL.n333 VSUBS 0.015053f
C1698 VTAIL.n334 VSUBS 0.015938f
C1699 VTAIL.n335 VSUBS 0.035579f
C1700 VTAIL.n336 VSUBS 0.035579f
C1701 VTAIL.n337 VSUBS 0.015938f
C1702 VTAIL.n338 VSUBS 0.015053f
C1703 VTAIL.n339 VSUBS 0.028012f
C1704 VTAIL.n340 VSUBS 0.028012f
C1705 VTAIL.n341 VSUBS 0.015053f
C1706 VTAIL.n342 VSUBS 0.015938f
C1707 VTAIL.n343 VSUBS 0.035579f
C1708 VTAIL.n344 VSUBS 0.035579f
C1709 VTAIL.n345 VSUBS 0.015938f
C1710 VTAIL.n346 VSUBS 0.015053f
C1711 VTAIL.n347 VSUBS 0.028012f
C1712 VTAIL.n348 VSUBS 0.028012f
C1713 VTAIL.n349 VSUBS 0.015053f
C1714 VTAIL.n350 VSUBS 0.015938f
C1715 VTAIL.n351 VSUBS 0.035579f
C1716 VTAIL.n352 VSUBS 0.035579f
C1717 VTAIL.n353 VSUBS 0.015938f
C1718 VTAIL.n354 VSUBS 0.015053f
C1719 VTAIL.n355 VSUBS 0.028012f
C1720 VTAIL.n356 VSUBS 0.028012f
C1721 VTAIL.n357 VSUBS 0.015053f
C1722 VTAIL.n358 VSUBS 0.015938f
C1723 VTAIL.n359 VSUBS 0.035579f
C1724 VTAIL.n360 VSUBS 0.035579f
C1725 VTAIL.n361 VSUBS 0.035579f
C1726 VTAIL.n362 VSUBS 0.015938f
C1727 VTAIL.n363 VSUBS 0.015053f
C1728 VTAIL.n364 VSUBS 0.028012f
C1729 VTAIL.n365 VSUBS 0.028012f
C1730 VTAIL.n366 VSUBS 0.015053f
C1731 VTAIL.n367 VSUBS 0.015495f
C1732 VTAIL.n368 VSUBS 0.015495f
C1733 VTAIL.n369 VSUBS 0.035579f
C1734 VTAIL.n370 VSUBS 0.035579f
C1735 VTAIL.n371 VSUBS 0.015938f
C1736 VTAIL.n372 VSUBS 0.015053f
C1737 VTAIL.n373 VSUBS 0.028012f
C1738 VTAIL.n374 VSUBS 0.028012f
C1739 VTAIL.n375 VSUBS 0.015053f
C1740 VTAIL.n376 VSUBS 0.015938f
C1741 VTAIL.n377 VSUBS 0.035579f
C1742 VTAIL.n378 VSUBS 0.087352f
C1743 VTAIL.n379 VSUBS 0.015938f
C1744 VTAIL.n380 VSUBS 0.015053f
C1745 VTAIL.n381 VSUBS 0.069341f
C1746 VTAIL.n382 VSUBS 0.044119f
C1747 VTAIL.n383 VSUBS 2.1759f
C1748 VP.t5 VSUBS 3.88313f
C1749 VP.n0 VSUBS 1.45204f
C1750 VP.n1 VSUBS 0.02757f
C1751 VP.n2 VSUBS 0.035007f
C1752 VP.n3 VSUBS 0.02757f
C1753 VP.t2 VSUBS 3.88313f
C1754 VP.n4 VSUBS 0.051641f
C1755 VP.n5 VSUBS 0.02757f
C1756 VP.n6 VSUBS 0.051641f
C1757 VP.t0 VSUBS 3.88313f
C1758 VP.n7 VSUBS 1.45204f
C1759 VP.n8 VSUBS 0.02757f
C1760 VP.n9 VSUBS 0.035007f
C1761 VP.n10 VSUBS 0.313738f
C1762 VP.t3 VSUBS 3.88313f
C1763 VP.t4 VSUBS 4.18762f
C1764 VP.n11 VSUBS 1.38777f
C1765 VP.n12 VSUBS 1.44903f
C1766 VP.n13 VSUBS 0.051641f
C1767 VP.n14 VSUBS 0.051641f
C1768 VP.n15 VSUBS 0.02757f
C1769 VP.n16 VSUBS 0.02757f
C1770 VP.n17 VSUBS 0.02757f
C1771 VP.n18 VSUBS 0.045839f
C1772 VP.n19 VSUBS 0.051641f
C1773 VP.n20 VSUBS 0.044502f
C1774 VP.n21 VSUBS 0.044505f
C1775 VP.n22 VSUBS 1.74936f
C1776 VP.n23 VSUBS 1.7676f
C1777 VP.t1 VSUBS 3.88313f
C1778 VP.n24 VSUBS 1.45204f
C1779 VP.n25 VSUBS 0.044502f
C1780 VP.n26 VSUBS 0.044505f
C1781 VP.n27 VSUBS 0.02757f
C1782 VP.n28 VSUBS 0.02757f
C1783 VP.n29 VSUBS 0.045839f
C1784 VP.n30 VSUBS 0.035007f
C1785 VP.n31 VSUBS 0.051641f
C1786 VP.n32 VSUBS 0.02757f
C1787 VP.n33 VSUBS 0.02757f
C1788 VP.n34 VSUBS 0.02757f
C1789 VP.n35 VSUBS 1.37203f
C1790 VP.n36 VSUBS 0.051641f
C1791 VP.n37 VSUBS 0.051641f
C1792 VP.n38 VSUBS 0.02757f
C1793 VP.n39 VSUBS 0.02757f
C1794 VP.n40 VSUBS 0.02757f
C1795 VP.n41 VSUBS 0.045839f
C1796 VP.n42 VSUBS 0.051641f
C1797 VP.n43 VSUBS 0.044502f
C1798 VP.n44 VSUBS 0.044505f
C1799 VP.n45 VSUBS 0.060561f
.ends

