* NGSPICE file created from diff_pair_sample_1061.ext - technology: sky130A

.subckt diff_pair_sample_1061 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t7 VP.t0 VTAIL.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=1.1154 pd=7.09 as=2.6364 ps=14.3 w=6.76 l=0.81
X1 B.t21 B.t19 B.t20 B.t9 sky130_fd_pr__nfet_01v8 ad=2.6364 pd=14.3 as=0 ps=0 w=6.76 l=0.81
X2 VDD1.t6 VP.t1 VTAIL.t10 B.t0 sky130_fd_pr__nfet_01v8 ad=1.1154 pd=7.09 as=2.6364 ps=14.3 w=6.76 l=0.81
X3 B.t18 B.t16 B.t17 B.t13 sky130_fd_pr__nfet_01v8 ad=2.6364 pd=14.3 as=0 ps=0 w=6.76 l=0.81
X4 VDD2.t7 VN.t0 VTAIL.t12 B.t5 sky130_fd_pr__nfet_01v8 ad=1.1154 pd=7.09 as=1.1154 ps=7.09 w=6.76 l=0.81
X5 VTAIL.t3 VN.t1 VDD2.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=1.1154 pd=7.09 as=1.1154 ps=7.09 w=6.76 l=0.81
X6 VTAIL.t9 VP.t2 VDD1.t5 B.t1 sky130_fd_pr__nfet_01v8 ad=2.6364 pd=14.3 as=1.1154 ps=7.09 w=6.76 l=0.81
X7 VDD2.t5 VN.t2 VTAIL.t13 B.t6 sky130_fd_pr__nfet_01v8 ad=1.1154 pd=7.09 as=1.1154 ps=7.09 w=6.76 l=0.81
X8 VDD1.t4 VP.t3 VTAIL.t7 B.t6 sky130_fd_pr__nfet_01v8 ad=1.1154 pd=7.09 as=1.1154 ps=7.09 w=6.76 l=0.81
X9 VTAIL.t1 VN.t3 VDD2.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=2.6364 pd=14.3 as=1.1154 ps=7.09 w=6.76 l=0.81
X10 VDD2.t3 VN.t4 VTAIL.t14 B.t7 sky130_fd_pr__nfet_01v8 ad=1.1154 pd=7.09 as=2.6364 ps=14.3 w=6.76 l=0.81
X11 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=2.6364 pd=14.3 as=0 ps=0 w=6.76 l=0.81
X12 VDD1.t3 VP.t4 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=1.1154 pd=7.09 as=1.1154 ps=7.09 w=6.76 l=0.81
X13 VTAIL.t15 VN.t5 VDD2.t2 B.t4 sky130_fd_pr__nfet_01v8 ad=2.6364 pd=14.3 as=1.1154 ps=7.09 w=6.76 l=0.81
X14 VTAIL.t4 VP.t5 VDD1.t2 B.t4 sky130_fd_pr__nfet_01v8 ad=2.6364 pd=14.3 as=1.1154 ps=7.09 w=6.76 l=0.81
X15 VTAIL.t8 VP.t6 VDD1.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=1.1154 pd=7.09 as=1.1154 ps=7.09 w=6.76 l=0.81
X16 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=2.6364 pd=14.3 as=0 ps=0 w=6.76 l=0.81
X17 VTAIL.t6 VP.t7 VDD1.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=1.1154 pd=7.09 as=1.1154 ps=7.09 w=6.76 l=0.81
X18 VTAIL.t2 VN.t6 VDD2.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=1.1154 pd=7.09 as=1.1154 ps=7.09 w=6.76 l=0.81
X19 VDD2.t0 VN.t7 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.1154 pd=7.09 as=2.6364 ps=14.3 w=6.76 l=0.81
R0 VP.n4 VP.t2 270.652
R1 VP.n11 VP.t5 249.629
R2 VP.n1 VP.t4 249.629
R3 VP.n16 VP.t6 249.629
R4 VP.n18 VP.t0 249.629
R5 VP.n8 VP.t1 249.629
R6 VP.n6 VP.t7 249.629
R7 VP.n5 VP.t3 249.629
R8 VP.n19 VP.n18 161.3
R9 VP.n7 VP.n2 161.3
R10 VP.n9 VP.n8 161.3
R11 VP.n17 VP.n0 161.3
R12 VP.n13 VP.n12 161.3
R13 VP.n11 VP.n10 161.3
R14 VP.n6 VP.n3 80.6037
R15 VP.n16 VP.n15 80.6037
R16 VP.n14 VP.n1 80.6037
R17 VP.n16 VP.n1 48.2005
R18 VP.n6 VP.n5 48.2005
R19 VP.n12 VP.n1 40.1672
R20 VP.n17 VP.n16 40.1672
R21 VP.n7 VP.n6 40.1672
R22 VP.n10 VP.n9 38.5005
R23 VP.n4 VP.n3 31.6481
R24 VP.n5 VP.n4 17.444
R25 VP.n12 VP.n11 8.03383
R26 VP.n18 VP.n17 8.03383
R27 VP.n8 VP.n7 8.03383
R28 VP.n15 VP.n14 0.380177
R29 VP.n3 VP.n2 0.285035
R30 VP.n14 VP.n13 0.285035
R31 VP.n15 VP.n0 0.285035
R32 VP.n9 VP.n2 0.189894
R33 VP.n13 VP.n10 0.189894
R34 VP.n19 VP.n0 0.189894
R35 VP VP.n19 0.0516364
R36 VTAIL.n290 VTAIL.n260 289.615
R37 VTAIL.n32 VTAIL.n2 289.615
R38 VTAIL.n68 VTAIL.n38 289.615
R39 VTAIL.n106 VTAIL.n76 289.615
R40 VTAIL.n254 VTAIL.n224 289.615
R41 VTAIL.n216 VTAIL.n186 289.615
R42 VTAIL.n180 VTAIL.n150 289.615
R43 VTAIL.n142 VTAIL.n112 289.615
R44 VTAIL.n273 VTAIL.n272 185
R45 VTAIL.n275 VTAIL.n274 185
R46 VTAIL.n268 VTAIL.n267 185
R47 VTAIL.n281 VTAIL.n280 185
R48 VTAIL.n283 VTAIL.n282 185
R49 VTAIL.n264 VTAIL.n263 185
R50 VTAIL.n289 VTAIL.n288 185
R51 VTAIL.n291 VTAIL.n290 185
R52 VTAIL.n15 VTAIL.n14 185
R53 VTAIL.n17 VTAIL.n16 185
R54 VTAIL.n10 VTAIL.n9 185
R55 VTAIL.n23 VTAIL.n22 185
R56 VTAIL.n25 VTAIL.n24 185
R57 VTAIL.n6 VTAIL.n5 185
R58 VTAIL.n31 VTAIL.n30 185
R59 VTAIL.n33 VTAIL.n32 185
R60 VTAIL.n51 VTAIL.n50 185
R61 VTAIL.n53 VTAIL.n52 185
R62 VTAIL.n46 VTAIL.n45 185
R63 VTAIL.n59 VTAIL.n58 185
R64 VTAIL.n61 VTAIL.n60 185
R65 VTAIL.n42 VTAIL.n41 185
R66 VTAIL.n67 VTAIL.n66 185
R67 VTAIL.n69 VTAIL.n68 185
R68 VTAIL.n89 VTAIL.n88 185
R69 VTAIL.n91 VTAIL.n90 185
R70 VTAIL.n84 VTAIL.n83 185
R71 VTAIL.n97 VTAIL.n96 185
R72 VTAIL.n99 VTAIL.n98 185
R73 VTAIL.n80 VTAIL.n79 185
R74 VTAIL.n105 VTAIL.n104 185
R75 VTAIL.n107 VTAIL.n106 185
R76 VTAIL.n255 VTAIL.n254 185
R77 VTAIL.n253 VTAIL.n252 185
R78 VTAIL.n228 VTAIL.n227 185
R79 VTAIL.n247 VTAIL.n246 185
R80 VTAIL.n245 VTAIL.n244 185
R81 VTAIL.n232 VTAIL.n231 185
R82 VTAIL.n239 VTAIL.n238 185
R83 VTAIL.n237 VTAIL.n236 185
R84 VTAIL.n217 VTAIL.n216 185
R85 VTAIL.n215 VTAIL.n214 185
R86 VTAIL.n190 VTAIL.n189 185
R87 VTAIL.n209 VTAIL.n208 185
R88 VTAIL.n207 VTAIL.n206 185
R89 VTAIL.n194 VTAIL.n193 185
R90 VTAIL.n201 VTAIL.n200 185
R91 VTAIL.n199 VTAIL.n198 185
R92 VTAIL.n181 VTAIL.n180 185
R93 VTAIL.n179 VTAIL.n178 185
R94 VTAIL.n154 VTAIL.n153 185
R95 VTAIL.n173 VTAIL.n172 185
R96 VTAIL.n171 VTAIL.n170 185
R97 VTAIL.n158 VTAIL.n157 185
R98 VTAIL.n165 VTAIL.n164 185
R99 VTAIL.n163 VTAIL.n162 185
R100 VTAIL.n143 VTAIL.n142 185
R101 VTAIL.n141 VTAIL.n140 185
R102 VTAIL.n116 VTAIL.n115 185
R103 VTAIL.n135 VTAIL.n134 185
R104 VTAIL.n133 VTAIL.n132 185
R105 VTAIL.n120 VTAIL.n119 185
R106 VTAIL.n127 VTAIL.n126 185
R107 VTAIL.n125 VTAIL.n124 185
R108 VTAIL.n271 VTAIL.t0 147.659
R109 VTAIL.n13 VTAIL.t1 147.659
R110 VTAIL.n49 VTAIL.t11 147.659
R111 VTAIL.n87 VTAIL.t4 147.659
R112 VTAIL.n235 VTAIL.t10 147.659
R113 VTAIL.n197 VTAIL.t9 147.659
R114 VTAIL.n161 VTAIL.t14 147.659
R115 VTAIL.n123 VTAIL.t15 147.659
R116 VTAIL.n274 VTAIL.n273 104.615
R117 VTAIL.n274 VTAIL.n267 104.615
R118 VTAIL.n281 VTAIL.n267 104.615
R119 VTAIL.n282 VTAIL.n281 104.615
R120 VTAIL.n282 VTAIL.n263 104.615
R121 VTAIL.n289 VTAIL.n263 104.615
R122 VTAIL.n290 VTAIL.n289 104.615
R123 VTAIL.n16 VTAIL.n15 104.615
R124 VTAIL.n16 VTAIL.n9 104.615
R125 VTAIL.n23 VTAIL.n9 104.615
R126 VTAIL.n24 VTAIL.n23 104.615
R127 VTAIL.n24 VTAIL.n5 104.615
R128 VTAIL.n31 VTAIL.n5 104.615
R129 VTAIL.n32 VTAIL.n31 104.615
R130 VTAIL.n52 VTAIL.n51 104.615
R131 VTAIL.n52 VTAIL.n45 104.615
R132 VTAIL.n59 VTAIL.n45 104.615
R133 VTAIL.n60 VTAIL.n59 104.615
R134 VTAIL.n60 VTAIL.n41 104.615
R135 VTAIL.n67 VTAIL.n41 104.615
R136 VTAIL.n68 VTAIL.n67 104.615
R137 VTAIL.n90 VTAIL.n89 104.615
R138 VTAIL.n90 VTAIL.n83 104.615
R139 VTAIL.n97 VTAIL.n83 104.615
R140 VTAIL.n98 VTAIL.n97 104.615
R141 VTAIL.n98 VTAIL.n79 104.615
R142 VTAIL.n105 VTAIL.n79 104.615
R143 VTAIL.n106 VTAIL.n105 104.615
R144 VTAIL.n254 VTAIL.n253 104.615
R145 VTAIL.n253 VTAIL.n227 104.615
R146 VTAIL.n246 VTAIL.n227 104.615
R147 VTAIL.n246 VTAIL.n245 104.615
R148 VTAIL.n245 VTAIL.n231 104.615
R149 VTAIL.n238 VTAIL.n231 104.615
R150 VTAIL.n238 VTAIL.n237 104.615
R151 VTAIL.n216 VTAIL.n215 104.615
R152 VTAIL.n215 VTAIL.n189 104.615
R153 VTAIL.n208 VTAIL.n189 104.615
R154 VTAIL.n208 VTAIL.n207 104.615
R155 VTAIL.n207 VTAIL.n193 104.615
R156 VTAIL.n200 VTAIL.n193 104.615
R157 VTAIL.n200 VTAIL.n199 104.615
R158 VTAIL.n180 VTAIL.n179 104.615
R159 VTAIL.n179 VTAIL.n153 104.615
R160 VTAIL.n172 VTAIL.n153 104.615
R161 VTAIL.n172 VTAIL.n171 104.615
R162 VTAIL.n171 VTAIL.n157 104.615
R163 VTAIL.n164 VTAIL.n157 104.615
R164 VTAIL.n164 VTAIL.n163 104.615
R165 VTAIL.n142 VTAIL.n141 104.615
R166 VTAIL.n141 VTAIL.n115 104.615
R167 VTAIL.n134 VTAIL.n115 104.615
R168 VTAIL.n134 VTAIL.n133 104.615
R169 VTAIL.n133 VTAIL.n119 104.615
R170 VTAIL.n126 VTAIL.n119 104.615
R171 VTAIL.n126 VTAIL.n125 104.615
R172 VTAIL.n273 VTAIL.t0 52.3082
R173 VTAIL.n15 VTAIL.t1 52.3082
R174 VTAIL.n51 VTAIL.t11 52.3082
R175 VTAIL.n89 VTAIL.t4 52.3082
R176 VTAIL.n237 VTAIL.t10 52.3082
R177 VTAIL.n199 VTAIL.t9 52.3082
R178 VTAIL.n163 VTAIL.t14 52.3082
R179 VTAIL.n125 VTAIL.t15 52.3082
R180 VTAIL.n223 VTAIL.n222 50.1711
R181 VTAIL.n149 VTAIL.n148 50.1711
R182 VTAIL.n1 VTAIL.n0 50.1709
R183 VTAIL.n75 VTAIL.n74 50.1709
R184 VTAIL.n295 VTAIL.n294 32.9611
R185 VTAIL.n37 VTAIL.n36 32.9611
R186 VTAIL.n73 VTAIL.n72 32.9611
R187 VTAIL.n111 VTAIL.n110 32.9611
R188 VTAIL.n259 VTAIL.n258 32.9611
R189 VTAIL.n221 VTAIL.n220 32.9611
R190 VTAIL.n185 VTAIL.n184 32.9611
R191 VTAIL.n147 VTAIL.n146 32.9611
R192 VTAIL.n295 VTAIL.n259 19.1772
R193 VTAIL.n147 VTAIL.n111 19.1772
R194 VTAIL.n272 VTAIL.n271 15.6676
R195 VTAIL.n14 VTAIL.n13 15.6676
R196 VTAIL.n50 VTAIL.n49 15.6676
R197 VTAIL.n88 VTAIL.n87 15.6676
R198 VTAIL.n236 VTAIL.n235 15.6676
R199 VTAIL.n198 VTAIL.n197 15.6676
R200 VTAIL.n162 VTAIL.n161 15.6676
R201 VTAIL.n124 VTAIL.n123 15.6676
R202 VTAIL.n275 VTAIL.n270 12.8005
R203 VTAIL.n17 VTAIL.n12 12.8005
R204 VTAIL.n53 VTAIL.n48 12.8005
R205 VTAIL.n91 VTAIL.n86 12.8005
R206 VTAIL.n239 VTAIL.n234 12.8005
R207 VTAIL.n201 VTAIL.n196 12.8005
R208 VTAIL.n165 VTAIL.n160 12.8005
R209 VTAIL.n127 VTAIL.n122 12.8005
R210 VTAIL.n276 VTAIL.n268 12.0247
R211 VTAIL.n18 VTAIL.n10 12.0247
R212 VTAIL.n54 VTAIL.n46 12.0247
R213 VTAIL.n92 VTAIL.n84 12.0247
R214 VTAIL.n240 VTAIL.n232 12.0247
R215 VTAIL.n202 VTAIL.n194 12.0247
R216 VTAIL.n166 VTAIL.n158 12.0247
R217 VTAIL.n128 VTAIL.n120 12.0247
R218 VTAIL.n280 VTAIL.n279 11.249
R219 VTAIL.n22 VTAIL.n21 11.249
R220 VTAIL.n58 VTAIL.n57 11.249
R221 VTAIL.n96 VTAIL.n95 11.249
R222 VTAIL.n244 VTAIL.n243 11.249
R223 VTAIL.n206 VTAIL.n205 11.249
R224 VTAIL.n170 VTAIL.n169 11.249
R225 VTAIL.n132 VTAIL.n131 11.249
R226 VTAIL.n283 VTAIL.n266 10.4732
R227 VTAIL.n25 VTAIL.n8 10.4732
R228 VTAIL.n61 VTAIL.n44 10.4732
R229 VTAIL.n99 VTAIL.n82 10.4732
R230 VTAIL.n247 VTAIL.n230 10.4732
R231 VTAIL.n209 VTAIL.n192 10.4732
R232 VTAIL.n173 VTAIL.n156 10.4732
R233 VTAIL.n135 VTAIL.n118 10.4732
R234 VTAIL.n284 VTAIL.n264 9.69747
R235 VTAIL.n26 VTAIL.n6 9.69747
R236 VTAIL.n62 VTAIL.n42 9.69747
R237 VTAIL.n100 VTAIL.n80 9.69747
R238 VTAIL.n248 VTAIL.n228 9.69747
R239 VTAIL.n210 VTAIL.n190 9.69747
R240 VTAIL.n174 VTAIL.n154 9.69747
R241 VTAIL.n136 VTAIL.n116 9.69747
R242 VTAIL.n294 VTAIL.n293 9.45567
R243 VTAIL.n36 VTAIL.n35 9.45567
R244 VTAIL.n72 VTAIL.n71 9.45567
R245 VTAIL.n110 VTAIL.n109 9.45567
R246 VTAIL.n258 VTAIL.n257 9.45567
R247 VTAIL.n220 VTAIL.n219 9.45567
R248 VTAIL.n184 VTAIL.n183 9.45567
R249 VTAIL.n146 VTAIL.n145 9.45567
R250 VTAIL.n262 VTAIL.n261 9.3005
R251 VTAIL.n287 VTAIL.n286 9.3005
R252 VTAIL.n285 VTAIL.n284 9.3005
R253 VTAIL.n266 VTAIL.n265 9.3005
R254 VTAIL.n279 VTAIL.n278 9.3005
R255 VTAIL.n277 VTAIL.n276 9.3005
R256 VTAIL.n270 VTAIL.n269 9.3005
R257 VTAIL.n293 VTAIL.n292 9.3005
R258 VTAIL.n4 VTAIL.n3 9.3005
R259 VTAIL.n29 VTAIL.n28 9.3005
R260 VTAIL.n27 VTAIL.n26 9.3005
R261 VTAIL.n8 VTAIL.n7 9.3005
R262 VTAIL.n21 VTAIL.n20 9.3005
R263 VTAIL.n19 VTAIL.n18 9.3005
R264 VTAIL.n12 VTAIL.n11 9.3005
R265 VTAIL.n35 VTAIL.n34 9.3005
R266 VTAIL.n40 VTAIL.n39 9.3005
R267 VTAIL.n65 VTAIL.n64 9.3005
R268 VTAIL.n63 VTAIL.n62 9.3005
R269 VTAIL.n44 VTAIL.n43 9.3005
R270 VTAIL.n57 VTAIL.n56 9.3005
R271 VTAIL.n55 VTAIL.n54 9.3005
R272 VTAIL.n48 VTAIL.n47 9.3005
R273 VTAIL.n71 VTAIL.n70 9.3005
R274 VTAIL.n78 VTAIL.n77 9.3005
R275 VTAIL.n103 VTAIL.n102 9.3005
R276 VTAIL.n101 VTAIL.n100 9.3005
R277 VTAIL.n82 VTAIL.n81 9.3005
R278 VTAIL.n95 VTAIL.n94 9.3005
R279 VTAIL.n93 VTAIL.n92 9.3005
R280 VTAIL.n86 VTAIL.n85 9.3005
R281 VTAIL.n109 VTAIL.n108 9.3005
R282 VTAIL.n257 VTAIL.n256 9.3005
R283 VTAIL.n226 VTAIL.n225 9.3005
R284 VTAIL.n251 VTAIL.n250 9.3005
R285 VTAIL.n249 VTAIL.n248 9.3005
R286 VTAIL.n230 VTAIL.n229 9.3005
R287 VTAIL.n243 VTAIL.n242 9.3005
R288 VTAIL.n241 VTAIL.n240 9.3005
R289 VTAIL.n234 VTAIL.n233 9.3005
R290 VTAIL.n219 VTAIL.n218 9.3005
R291 VTAIL.n188 VTAIL.n187 9.3005
R292 VTAIL.n213 VTAIL.n212 9.3005
R293 VTAIL.n211 VTAIL.n210 9.3005
R294 VTAIL.n192 VTAIL.n191 9.3005
R295 VTAIL.n205 VTAIL.n204 9.3005
R296 VTAIL.n203 VTAIL.n202 9.3005
R297 VTAIL.n196 VTAIL.n195 9.3005
R298 VTAIL.n183 VTAIL.n182 9.3005
R299 VTAIL.n152 VTAIL.n151 9.3005
R300 VTAIL.n177 VTAIL.n176 9.3005
R301 VTAIL.n175 VTAIL.n174 9.3005
R302 VTAIL.n156 VTAIL.n155 9.3005
R303 VTAIL.n169 VTAIL.n168 9.3005
R304 VTAIL.n167 VTAIL.n166 9.3005
R305 VTAIL.n160 VTAIL.n159 9.3005
R306 VTAIL.n145 VTAIL.n144 9.3005
R307 VTAIL.n114 VTAIL.n113 9.3005
R308 VTAIL.n139 VTAIL.n138 9.3005
R309 VTAIL.n137 VTAIL.n136 9.3005
R310 VTAIL.n118 VTAIL.n117 9.3005
R311 VTAIL.n131 VTAIL.n130 9.3005
R312 VTAIL.n129 VTAIL.n128 9.3005
R313 VTAIL.n122 VTAIL.n121 9.3005
R314 VTAIL.n288 VTAIL.n287 8.92171
R315 VTAIL.n30 VTAIL.n29 8.92171
R316 VTAIL.n66 VTAIL.n65 8.92171
R317 VTAIL.n104 VTAIL.n103 8.92171
R318 VTAIL.n252 VTAIL.n251 8.92171
R319 VTAIL.n214 VTAIL.n213 8.92171
R320 VTAIL.n178 VTAIL.n177 8.92171
R321 VTAIL.n140 VTAIL.n139 8.92171
R322 VTAIL.n291 VTAIL.n262 8.14595
R323 VTAIL.n33 VTAIL.n4 8.14595
R324 VTAIL.n69 VTAIL.n40 8.14595
R325 VTAIL.n107 VTAIL.n78 8.14595
R326 VTAIL.n255 VTAIL.n226 8.14595
R327 VTAIL.n217 VTAIL.n188 8.14595
R328 VTAIL.n181 VTAIL.n152 8.14595
R329 VTAIL.n143 VTAIL.n114 8.14595
R330 VTAIL.n292 VTAIL.n260 7.3702
R331 VTAIL.n34 VTAIL.n2 7.3702
R332 VTAIL.n70 VTAIL.n38 7.3702
R333 VTAIL.n108 VTAIL.n76 7.3702
R334 VTAIL.n256 VTAIL.n224 7.3702
R335 VTAIL.n218 VTAIL.n186 7.3702
R336 VTAIL.n182 VTAIL.n150 7.3702
R337 VTAIL.n144 VTAIL.n112 7.3702
R338 VTAIL.n294 VTAIL.n260 6.59444
R339 VTAIL.n36 VTAIL.n2 6.59444
R340 VTAIL.n72 VTAIL.n38 6.59444
R341 VTAIL.n110 VTAIL.n76 6.59444
R342 VTAIL.n258 VTAIL.n224 6.59444
R343 VTAIL.n220 VTAIL.n186 6.59444
R344 VTAIL.n184 VTAIL.n150 6.59444
R345 VTAIL.n146 VTAIL.n112 6.59444
R346 VTAIL.n292 VTAIL.n291 5.81868
R347 VTAIL.n34 VTAIL.n33 5.81868
R348 VTAIL.n70 VTAIL.n69 5.81868
R349 VTAIL.n108 VTAIL.n107 5.81868
R350 VTAIL.n256 VTAIL.n255 5.81868
R351 VTAIL.n218 VTAIL.n217 5.81868
R352 VTAIL.n182 VTAIL.n181 5.81868
R353 VTAIL.n144 VTAIL.n143 5.81868
R354 VTAIL.n288 VTAIL.n262 5.04292
R355 VTAIL.n30 VTAIL.n4 5.04292
R356 VTAIL.n66 VTAIL.n40 5.04292
R357 VTAIL.n104 VTAIL.n78 5.04292
R358 VTAIL.n252 VTAIL.n226 5.04292
R359 VTAIL.n214 VTAIL.n188 5.04292
R360 VTAIL.n178 VTAIL.n152 5.04292
R361 VTAIL.n140 VTAIL.n114 5.04292
R362 VTAIL.n271 VTAIL.n269 4.38571
R363 VTAIL.n13 VTAIL.n11 4.38571
R364 VTAIL.n49 VTAIL.n47 4.38571
R365 VTAIL.n87 VTAIL.n85 4.38571
R366 VTAIL.n235 VTAIL.n233 4.38571
R367 VTAIL.n197 VTAIL.n195 4.38571
R368 VTAIL.n161 VTAIL.n159 4.38571
R369 VTAIL.n123 VTAIL.n121 4.38571
R370 VTAIL.n287 VTAIL.n264 4.26717
R371 VTAIL.n29 VTAIL.n6 4.26717
R372 VTAIL.n65 VTAIL.n42 4.26717
R373 VTAIL.n103 VTAIL.n80 4.26717
R374 VTAIL.n251 VTAIL.n228 4.26717
R375 VTAIL.n213 VTAIL.n190 4.26717
R376 VTAIL.n177 VTAIL.n154 4.26717
R377 VTAIL.n139 VTAIL.n116 4.26717
R378 VTAIL.n284 VTAIL.n283 3.49141
R379 VTAIL.n26 VTAIL.n25 3.49141
R380 VTAIL.n62 VTAIL.n61 3.49141
R381 VTAIL.n100 VTAIL.n99 3.49141
R382 VTAIL.n248 VTAIL.n247 3.49141
R383 VTAIL.n210 VTAIL.n209 3.49141
R384 VTAIL.n174 VTAIL.n173 3.49141
R385 VTAIL.n136 VTAIL.n135 3.49141
R386 VTAIL.n0 VTAIL.t13 2.92949
R387 VTAIL.n0 VTAIL.t3 2.92949
R388 VTAIL.n74 VTAIL.t5 2.92949
R389 VTAIL.n74 VTAIL.t8 2.92949
R390 VTAIL.n222 VTAIL.t7 2.92949
R391 VTAIL.n222 VTAIL.t6 2.92949
R392 VTAIL.n148 VTAIL.t12 2.92949
R393 VTAIL.n148 VTAIL.t2 2.92949
R394 VTAIL.n280 VTAIL.n266 2.71565
R395 VTAIL.n22 VTAIL.n8 2.71565
R396 VTAIL.n58 VTAIL.n44 2.71565
R397 VTAIL.n96 VTAIL.n82 2.71565
R398 VTAIL.n244 VTAIL.n230 2.71565
R399 VTAIL.n206 VTAIL.n192 2.71565
R400 VTAIL.n170 VTAIL.n156 2.71565
R401 VTAIL.n132 VTAIL.n118 2.71565
R402 VTAIL.n279 VTAIL.n268 1.93989
R403 VTAIL.n21 VTAIL.n10 1.93989
R404 VTAIL.n57 VTAIL.n46 1.93989
R405 VTAIL.n95 VTAIL.n84 1.93989
R406 VTAIL.n243 VTAIL.n232 1.93989
R407 VTAIL.n205 VTAIL.n194 1.93989
R408 VTAIL.n169 VTAIL.n158 1.93989
R409 VTAIL.n131 VTAIL.n120 1.93989
R410 VTAIL.n276 VTAIL.n275 1.16414
R411 VTAIL.n18 VTAIL.n17 1.16414
R412 VTAIL.n54 VTAIL.n53 1.16414
R413 VTAIL.n92 VTAIL.n91 1.16414
R414 VTAIL.n240 VTAIL.n239 1.16414
R415 VTAIL.n202 VTAIL.n201 1.16414
R416 VTAIL.n166 VTAIL.n165 1.16414
R417 VTAIL.n128 VTAIL.n127 1.16414
R418 VTAIL.n149 VTAIL.n147 0.983259
R419 VTAIL.n185 VTAIL.n149 0.983259
R420 VTAIL.n223 VTAIL.n221 0.983259
R421 VTAIL.n259 VTAIL.n223 0.983259
R422 VTAIL.n111 VTAIL.n75 0.983259
R423 VTAIL.n75 VTAIL.n73 0.983259
R424 VTAIL.n37 VTAIL.n1 0.983259
R425 VTAIL VTAIL.n295 0.925069
R426 VTAIL.n221 VTAIL.n185 0.470328
R427 VTAIL.n73 VTAIL.n37 0.470328
R428 VTAIL.n272 VTAIL.n270 0.388379
R429 VTAIL.n14 VTAIL.n12 0.388379
R430 VTAIL.n50 VTAIL.n48 0.388379
R431 VTAIL.n88 VTAIL.n86 0.388379
R432 VTAIL.n236 VTAIL.n234 0.388379
R433 VTAIL.n198 VTAIL.n196 0.388379
R434 VTAIL.n162 VTAIL.n160 0.388379
R435 VTAIL.n124 VTAIL.n122 0.388379
R436 VTAIL.n277 VTAIL.n269 0.155672
R437 VTAIL.n278 VTAIL.n277 0.155672
R438 VTAIL.n278 VTAIL.n265 0.155672
R439 VTAIL.n285 VTAIL.n265 0.155672
R440 VTAIL.n286 VTAIL.n285 0.155672
R441 VTAIL.n286 VTAIL.n261 0.155672
R442 VTAIL.n293 VTAIL.n261 0.155672
R443 VTAIL.n19 VTAIL.n11 0.155672
R444 VTAIL.n20 VTAIL.n19 0.155672
R445 VTAIL.n20 VTAIL.n7 0.155672
R446 VTAIL.n27 VTAIL.n7 0.155672
R447 VTAIL.n28 VTAIL.n27 0.155672
R448 VTAIL.n28 VTAIL.n3 0.155672
R449 VTAIL.n35 VTAIL.n3 0.155672
R450 VTAIL.n55 VTAIL.n47 0.155672
R451 VTAIL.n56 VTAIL.n55 0.155672
R452 VTAIL.n56 VTAIL.n43 0.155672
R453 VTAIL.n63 VTAIL.n43 0.155672
R454 VTAIL.n64 VTAIL.n63 0.155672
R455 VTAIL.n64 VTAIL.n39 0.155672
R456 VTAIL.n71 VTAIL.n39 0.155672
R457 VTAIL.n93 VTAIL.n85 0.155672
R458 VTAIL.n94 VTAIL.n93 0.155672
R459 VTAIL.n94 VTAIL.n81 0.155672
R460 VTAIL.n101 VTAIL.n81 0.155672
R461 VTAIL.n102 VTAIL.n101 0.155672
R462 VTAIL.n102 VTAIL.n77 0.155672
R463 VTAIL.n109 VTAIL.n77 0.155672
R464 VTAIL.n257 VTAIL.n225 0.155672
R465 VTAIL.n250 VTAIL.n225 0.155672
R466 VTAIL.n250 VTAIL.n249 0.155672
R467 VTAIL.n249 VTAIL.n229 0.155672
R468 VTAIL.n242 VTAIL.n229 0.155672
R469 VTAIL.n242 VTAIL.n241 0.155672
R470 VTAIL.n241 VTAIL.n233 0.155672
R471 VTAIL.n219 VTAIL.n187 0.155672
R472 VTAIL.n212 VTAIL.n187 0.155672
R473 VTAIL.n212 VTAIL.n211 0.155672
R474 VTAIL.n211 VTAIL.n191 0.155672
R475 VTAIL.n204 VTAIL.n191 0.155672
R476 VTAIL.n204 VTAIL.n203 0.155672
R477 VTAIL.n203 VTAIL.n195 0.155672
R478 VTAIL.n183 VTAIL.n151 0.155672
R479 VTAIL.n176 VTAIL.n151 0.155672
R480 VTAIL.n176 VTAIL.n175 0.155672
R481 VTAIL.n175 VTAIL.n155 0.155672
R482 VTAIL.n168 VTAIL.n155 0.155672
R483 VTAIL.n168 VTAIL.n167 0.155672
R484 VTAIL.n167 VTAIL.n159 0.155672
R485 VTAIL.n145 VTAIL.n113 0.155672
R486 VTAIL.n138 VTAIL.n113 0.155672
R487 VTAIL.n138 VTAIL.n137 0.155672
R488 VTAIL.n137 VTAIL.n117 0.155672
R489 VTAIL.n130 VTAIL.n117 0.155672
R490 VTAIL.n130 VTAIL.n129 0.155672
R491 VTAIL.n129 VTAIL.n121 0.155672
R492 VTAIL VTAIL.n1 0.0586897
R493 VDD1 VDD1.n0 67.3994
R494 VDD1.n3 VDD1.n2 67.2857
R495 VDD1.n3 VDD1.n1 67.2857
R496 VDD1.n5 VDD1.n4 66.8497
R497 VDD1.n5 VDD1.n3 34.5483
R498 VDD1.n4 VDD1.t0 2.92949
R499 VDD1.n4 VDD1.t6 2.92949
R500 VDD1.n0 VDD1.t5 2.92949
R501 VDD1.n0 VDD1.t4 2.92949
R502 VDD1.n2 VDD1.t1 2.92949
R503 VDD1.n2 VDD1.t7 2.92949
R504 VDD1.n1 VDD1.t2 2.92949
R505 VDD1.n1 VDD1.t3 2.92949
R506 VDD1 VDD1.n5 0.43369
R507 B.n523 B.n522 585
R508 B.n206 B.n79 585
R509 B.n205 B.n204 585
R510 B.n203 B.n202 585
R511 B.n201 B.n200 585
R512 B.n199 B.n198 585
R513 B.n197 B.n196 585
R514 B.n195 B.n194 585
R515 B.n193 B.n192 585
R516 B.n191 B.n190 585
R517 B.n189 B.n188 585
R518 B.n187 B.n186 585
R519 B.n185 B.n184 585
R520 B.n183 B.n182 585
R521 B.n181 B.n180 585
R522 B.n179 B.n178 585
R523 B.n177 B.n176 585
R524 B.n175 B.n174 585
R525 B.n173 B.n172 585
R526 B.n171 B.n170 585
R527 B.n169 B.n168 585
R528 B.n167 B.n166 585
R529 B.n165 B.n164 585
R530 B.n163 B.n162 585
R531 B.n161 B.n160 585
R532 B.n159 B.n158 585
R533 B.n157 B.n156 585
R534 B.n155 B.n154 585
R535 B.n153 B.n152 585
R536 B.n151 B.n150 585
R537 B.n149 B.n148 585
R538 B.n147 B.n146 585
R539 B.n145 B.n144 585
R540 B.n143 B.n142 585
R541 B.n141 B.n140 585
R542 B.n139 B.n138 585
R543 B.n137 B.n136 585
R544 B.n135 B.n134 585
R545 B.n133 B.n132 585
R546 B.n131 B.n130 585
R547 B.n129 B.n128 585
R548 B.n127 B.n126 585
R549 B.n125 B.n124 585
R550 B.n123 B.n122 585
R551 B.n121 B.n120 585
R552 B.n119 B.n118 585
R553 B.n117 B.n116 585
R554 B.n115 B.n114 585
R555 B.n113 B.n112 585
R556 B.n111 B.n110 585
R557 B.n109 B.n108 585
R558 B.n107 B.n106 585
R559 B.n105 B.n104 585
R560 B.n103 B.n102 585
R561 B.n101 B.n100 585
R562 B.n99 B.n98 585
R563 B.n97 B.n96 585
R564 B.n95 B.n94 585
R565 B.n93 B.n92 585
R566 B.n91 B.n90 585
R567 B.n89 B.n88 585
R568 B.n87 B.n86 585
R569 B.n521 B.n48 585
R570 B.n526 B.n48 585
R571 B.n520 B.n47 585
R572 B.n527 B.n47 585
R573 B.n519 B.n518 585
R574 B.n518 B.n43 585
R575 B.n517 B.n42 585
R576 B.n533 B.n42 585
R577 B.n516 B.n41 585
R578 B.n534 B.n41 585
R579 B.n515 B.n40 585
R580 B.n535 B.n40 585
R581 B.n514 B.n513 585
R582 B.n513 B.n36 585
R583 B.n512 B.n35 585
R584 B.n541 B.n35 585
R585 B.n511 B.n34 585
R586 B.n542 B.n34 585
R587 B.n510 B.n33 585
R588 B.n543 B.n33 585
R589 B.n509 B.n508 585
R590 B.n508 B.n29 585
R591 B.n507 B.n28 585
R592 B.n549 B.n28 585
R593 B.n506 B.n27 585
R594 B.n550 B.n27 585
R595 B.n505 B.n26 585
R596 B.n551 B.n26 585
R597 B.n504 B.n503 585
R598 B.n503 B.n22 585
R599 B.n502 B.n21 585
R600 B.n557 B.n21 585
R601 B.n501 B.n20 585
R602 B.n558 B.n20 585
R603 B.n500 B.n19 585
R604 B.n559 B.n19 585
R605 B.n499 B.n498 585
R606 B.n498 B.n18 585
R607 B.n497 B.n14 585
R608 B.n565 B.n14 585
R609 B.n496 B.n13 585
R610 B.n566 B.n13 585
R611 B.n495 B.n12 585
R612 B.n567 B.n12 585
R613 B.n494 B.n493 585
R614 B.n493 B.n8 585
R615 B.n492 B.n7 585
R616 B.n573 B.n7 585
R617 B.n491 B.n6 585
R618 B.n574 B.n6 585
R619 B.n490 B.n5 585
R620 B.n575 B.n5 585
R621 B.n489 B.n488 585
R622 B.n488 B.n4 585
R623 B.n487 B.n207 585
R624 B.n487 B.n486 585
R625 B.n477 B.n208 585
R626 B.n209 B.n208 585
R627 B.n479 B.n478 585
R628 B.n480 B.n479 585
R629 B.n476 B.n214 585
R630 B.n214 B.n213 585
R631 B.n475 B.n474 585
R632 B.n474 B.n473 585
R633 B.n216 B.n215 585
R634 B.n466 B.n216 585
R635 B.n465 B.n464 585
R636 B.n467 B.n465 585
R637 B.n463 B.n221 585
R638 B.n221 B.n220 585
R639 B.n462 B.n461 585
R640 B.n461 B.n460 585
R641 B.n223 B.n222 585
R642 B.n224 B.n223 585
R643 B.n453 B.n452 585
R644 B.n454 B.n453 585
R645 B.n451 B.n229 585
R646 B.n229 B.n228 585
R647 B.n450 B.n449 585
R648 B.n449 B.n448 585
R649 B.n231 B.n230 585
R650 B.n232 B.n231 585
R651 B.n441 B.n440 585
R652 B.n442 B.n441 585
R653 B.n439 B.n237 585
R654 B.n237 B.n236 585
R655 B.n438 B.n437 585
R656 B.n437 B.n436 585
R657 B.n239 B.n238 585
R658 B.n240 B.n239 585
R659 B.n429 B.n428 585
R660 B.n430 B.n429 585
R661 B.n427 B.n245 585
R662 B.n245 B.n244 585
R663 B.n426 B.n425 585
R664 B.n425 B.n424 585
R665 B.n247 B.n246 585
R666 B.n248 B.n247 585
R667 B.n417 B.n416 585
R668 B.n418 B.n417 585
R669 B.n415 B.n253 585
R670 B.n253 B.n252 585
R671 B.n410 B.n409 585
R672 B.n408 B.n286 585
R673 B.n407 B.n285 585
R674 B.n412 B.n285 585
R675 B.n406 B.n405 585
R676 B.n404 B.n403 585
R677 B.n402 B.n401 585
R678 B.n400 B.n399 585
R679 B.n398 B.n397 585
R680 B.n396 B.n395 585
R681 B.n394 B.n393 585
R682 B.n392 B.n391 585
R683 B.n390 B.n389 585
R684 B.n388 B.n387 585
R685 B.n386 B.n385 585
R686 B.n384 B.n383 585
R687 B.n382 B.n381 585
R688 B.n380 B.n379 585
R689 B.n378 B.n377 585
R690 B.n376 B.n375 585
R691 B.n374 B.n373 585
R692 B.n372 B.n371 585
R693 B.n370 B.n369 585
R694 B.n368 B.n367 585
R695 B.n366 B.n365 585
R696 B.n364 B.n363 585
R697 B.n362 B.n361 585
R698 B.n359 B.n358 585
R699 B.n357 B.n356 585
R700 B.n355 B.n354 585
R701 B.n353 B.n352 585
R702 B.n351 B.n350 585
R703 B.n349 B.n348 585
R704 B.n347 B.n346 585
R705 B.n345 B.n344 585
R706 B.n343 B.n342 585
R707 B.n341 B.n340 585
R708 B.n338 B.n337 585
R709 B.n336 B.n335 585
R710 B.n334 B.n333 585
R711 B.n332 B.n331 585
R712 B.n330 B.n329 585
R713 B.n328 B.n327 585
R714 B.n326 B.n325 585
R715 B.n324 B.n323 585
R716 B.n322 B.n321 585
R717 B.n320 B.n319 585
R718 B.n318 B.n317 585
R719 B.n316 B.n315 585
R720 B.n314 B.n313 585
R721 B.n312 B.n311 585
R722 B.n310 B.n309 585
R723 B.n308 B.n307 585
R724 B.n306 B.n305 585
R725 B.n304 B.n303 585
R726 B.n302 B.n301 585
R727 B.n300 B.n299 585
R728 B.n298 B.n297 585
R729 B.n296 B.n295 585
R730 B.n294 B.n293 585
R731 B.n292 B.n291 585
R732 B.n255 B.n254 585
R733 B.n414 B.n413 585
R734 B.n413 B.n412 585
R735 B.n251 B.n250 585
R736 B.n252 B.n251 585
R737 B.n420 B.n419 585
R738 B.n419 B.n418 585
R739 B.n421 B.n249 585
R740 B.n249 B.n248 585
R741 B.n423 B.n422 585
R742 B.n424 B.n423 585
R743 B.n243 B.n242 585
R744 B.n244 B.n243 585
R745 B.n432 B.n431 585
R746 B.n431 B.n430 585
R747 B.n433 B.n241 585
R748 B.n241 B.n240 585
R749 B.n435 B.n434 585
R750 B.n436 B.n435 585
R751 B.n235 B.n234 585
R752 B.n236 B.n235 585
R753 B.n444 B.n443 585
R754 B.n443 B.n442 585
R755 B.n445 B.n233 585
R756 B.n233 B.n232 585
R757 B.n447 B.n446 585
R758 B.n448 B.n447 585
R759 B.n227 B.n226 585
R760 B.n228 B.n227 585
R761 B.n456 B.n455 585
R762 B.n455 B.n454 585
R763 B.n457 B.n225 585
R764 B.n225 B.n224 585
R765 B.n459 B.n458 585
R766 B.n460 B.n459 585
R767 B.n219 B.n218 585
R768 B.n220 B.n219 585
R769 B.n469 B.n468 585
R770 B.n468 B.n467 585
R771 B.n470 B.n217 585
R772 B.n466 B.n217 585
R773 B.n472 B.n471 585
R774 B.n473 B.n472 585
R775 B.n212 B.n211 585
R776 B.n213 B.n212 585
R777 B.n482 B.n481 585
R778 B.n481 B.n480 585
R779 B.n483 B.n210 585
R780 B.n210 B.n209 585
R781 B.n485 B.n484 585
R782 B.n486 B.n485 585
R783 B.n2 B.n0 585
R784 B.n4 B.n2 585
R785 B.n3 B.n1 585
R786 B.n574 B.n3 585
R787 B.n572 B.n571 585
R788 B.n573 B.n572 585
R789 B.n570 B.n9 585
R790 B.n9 B.n8 585
R791 B.n569 B.n568 585
R792 B.n568 B.n567 585
R793 B.n11 B.n10 585
R794 B.n566 B.n11 585
R795 B.n564 B.n563 585
R796 B.n565 B.n564 585
R797 B.n562 B.n15 585
R798 B.n18 B.n15 585
R799 B.n561 B.n560 585
R800 B.n560 B.n559 585
R801 B.n17 B.n16 585
R802 B.n558 B.n17 585
R803 B.n556 B.n555 585
R804 B.n557 B.n556 585
R805 B.n554 B.n23 585
R806 B.n23 B.n22 585
R807 B.n553 B.n552 585
R808 B.n552 B.n551 585
R809 B.n25 B.n24 585
R810 B.n550 B.n25 585
R811 B.n548 B.n547 585
R812 B.n549 B.n548 585
R813 B.n546 B.n30 585
R814 B.n30 B.n29 585
R815 B.n545 B.n544 585
R816 B.n544 B.n543 585
R817 B.n32 B.n31 585
R818 B.n542 B.n32 585
R819 B.n540 B.n539 585
R820 B.n541 B.n540 585
R821 B.n538 B.n37 585
R822 B.n37 B.n36 585
R823 B.n537 B.n536 585
R824 B.n536 B.n535 585
R825 B.n39 B.n38 585
R826 B.n534 B.n39 585
R827 B.n532 B.n531 585
R828 B.n533 B.n532 585
R829 B.n530 B.n44 585
R830 B.n44 B.n43 585
R831 B.n529 B.n528 585
R832 B.n528 B.n527 585
R833 B.n46 B.n45 585
R834 B.n526 B.n46 585
R835 B.n577 B.n576 585
R836 B.n576 B.n575 585
R837 B.n410 B.n251 478.086
R838 B.n86 B.n46 478.086
R839 B.n413 B.n253 478.086
R840 B.n523 B.n48 478.086
R841 B.n289 B.t16 402.928
R842 B.n287 B.t12 402.928
R843 B.n83 B.t19 402.928
R844 B.n80 B.t8 402.928
R845 B.n525 B.n524 256.663
R846 B.n525 B.n78 256.663
R847 B.n525 B.n77 256.663
R848 B.n525 B.n76 256.663
R849 B.n525 B.n75 256.663
R850 B.n525 B.n74 256.663
R851 B.n525 B.n73 256.663
R852 B.n525 B.n72 256.663
R853 B.n525 B.n71 256.663
R854 B.n525 B.n70 256.663
R855 B.n525 B.n69 256.663
R856 B.n525 B.n68 256.663
R857 B.n525 B.n67 256.663
R858 B.n525 B.n66 256.663
R859 B.n525 B.n65 256.663
R860 B.n525 B.n64 256.663
R861 B.n525 B.n63 256.663
R862 B.n525 B.n62 256.663
R863 B.n525 B.n61 256.663
R864 B.n525 B.n60 256.663
R865 B.n525 B.n59 256.663
R866 B.n525 B.n58 256.663
R867 B.n525 B.n57 256.663
R868 B.n525 B.n56 256.663
R869 B.n525 B.n55 256.663
R870 B.n525 B.n54 256.663
R871 B.n525 B.n53 256.663
R872 B.n525 B.n52 256.663
R873 B.n525 B.n51 256.663
R874 B.n525 B.n50 256.663
R875 B.n525 B.n49 256.663
R876 B.n412 B.n411 256.663
R877 B.n412 B.n256 256.663
R878 B.n412 B.n257 256.663
R879 B.n412 B.n258 256.663
R880 B.n412 B.n259 256.663
R881 B.n412 B.n260 256.663
R882 B.n412 B.n261 256.663
R883 B.n412 B.n262 256.663
R884 B.n412 B.n263 256.663
R885 B.n412 B.n264 256.663
R886 B.n412 B.n265 256.663
R887 B.n412 B.n266 256.663
R888 B.n412 B.n267 256.663
R889 B.n412 B.n268 256.663
R890 B.n412 B.n269 256.663
R891 B.n412 B.n270 256.663
R892 B.n412 B.n271 256.663
R893 B.n412 B.n272 256.663
R894 B.n412 B.n273 256.663
R895 B.n412 B.n274 256.663
R896 B.n412 B.n275 256.663
R897 B.n412 B.n276 256.663
R898 B.n412 B.n277 256.663
R899 B.n412 B.n278 256.663
R900 B.n412 B.n279 256.663
R901 B.n412 B.n280 256.663
R902 B.n412 B.n281 256.663
R903 B.n412 B.n282 256.663
R904 B.n412 B.n283 256.663
R905 B.n412 B.n284 256.663
R906 B.n289 B.t18 214.326
R907 B.n80 B.t10 214.326
R908 B.n287 B.t15 214.326
R909 B.n83 B.t20 214.326
R910 B.n290 B.t17 192.216
R911 B.n81 B.t11 192.216
R912 B.n288 B.t14 192.216
R913 B.n84 B.t21 192.216
R914 B.n419 B.n251 163.367
R915 B.n419 B.n249 163.367
R916 B.n423 B.n249 163.367
R917 B.n423 B.n243 163.367
R918 B.n431 B.n243 163.367
R919 B.n431 B.n241 163.367
R920 B.n435 B.n241 163.367
R921 B.n435 B.n235 163.367
R922 B.n443 B.n235 163.367
R923 B.n443 B.n233 163.367
R924 B.n447 B.n233 163.367
R925 B.n447 B.n227 163.367
R926 B.n455 B.n227 163.367
R927 B.n455 B.n225 163.367
R928 B.n459 B.n225 163.367
R929 B.n459 B.n219 163.367
R930 B.n468 B.n219 163.367
R931 B.n468 B.n217 163.367
R932 B.n472 B.n217 163.367
R933 B.n472 B.n212 163.367
R934 B.n481 B.n212 163.367
R935 B.n481 B.n210 163.367
R936 B.n485 B.n210 163.367
R937 B.n485 B.n2 163.367
R938 B.n576 B.n2 163.367
R939 B.n576 B.n3 163.367
R940 B.n572 B.n3 163.367
R941 B.n572 B.n9 163.367
R942 B.n568 B.n9 163.367
R943 B.n568 B.n11 163.367
R944 B.n564 B.n11 163.367
R945 B.n564 B.n15 163.367
R946 B.n560 B.n15 163.367
R947 B.n560 B.n17 163.367
R948 B.n556 B.n17 163.367
R949 B.n556 B.n23 163.367
R950 B.n552 B.n23 163.367
R951 B.n552 B.n25 163.367
R952 B.n548 B.n25 163.367
R953 B.n548 B.n30 163.367
R954 B.n544 B.n30 163.367
R955 B.n544 B.n32 163.367
R956 B.n540 B.n32 163.367
R957 B.n540 B.n37 163.367
R958 B.n536 B.n37 163.367
R959 B.n536 B.n39 163.367
R960 B.n532 B.n39 163.367
R961 B.n532 B.n44 163.367
R962 B.n528 B.n44 163.367
R963 B.n528 B.n46 163.367
R964 B.n286 B.n285 163.367
R965 B.n405 B.n285 163.367
R966 B.n403 B.n402 163.367
R967 B.n399 B.n398 163.367
R968 B.n395 B.n394 163.367
R969 B.n391 B.n390 163.367
R970 B.n387 B.n386 163.367
R971 B.n383 B.n382 163.367
R972 B.n379 B.n378 163.367
R973 B.n375 B.n374 163.367
R974 B.n371 B.n370 163.367
R975 B.n367 B.n366 163.367
R976 B.n363 B.n362 163.367
R977 B.n358 B.n357 163.367
R978 B.n354 B.n353 163.367
R979 B.n350 B.n349 163.367
R980 B.n346 B.n345 163.367
R981 B.n342 B.n341 163.367
R982 B.n337 B.n336 163.367
R983 B.n333 B.n332 163.367
R984 B.n329 B.n328 163.367
R985 B.n325 B.n324 163.367
R986 B.n321 B.n320 163.367
R987 B.n317 B.n316 163.367
R988 B.n313 B.n312 163.367
R989 B.n309 B.n308 163.367
R990 B.n305 B.n304 163.367
R991 B.n301 B.n300 163.367
R992 B.n297 B.n296 163.367
R993 B.n293 B.n292 163.367
R994 B.n413 B.n255 163.367
R995 B.n417 B.n253 163.367
R996 B.n417 B.n247 163.367
R997 B.n425 B.n247 163.367
R998 B.n425 B.n245 163.367
R999 B.n429 B.n245 163.367
R1000 B.n429 B.n239 163.367
R1001 B.n437 B.n239 163.367
R1002 B.n437 B.n237 163.367
R1003 B.n441 B.n237 163.367
R1004 B.n441 B.n231 163.367
R1005 B.n449 B.n231 163.367
R1006 B.n449 B.n229 163.367
R1007 B.n453 B.n229 163.367
R1008 B.n453 B.n223 163.367
R1009 B.n461 B.n223 163.367
R1010 B.n461 B.n221 163.367
R1011 B.n465 B.n221 163.367
R1012 B.n465 B.n216 163.367
R1013 B.n474 B.n216 163.367
R1014 B.n474 B.n214 163.367
R1015 B.n479 B.n214 163.367
R1016 B.n479 B.n208 163.367
R1017 B.n487 B.n208 163.367
R1018 B.n488 B.n487 163.367
R1019 B.n488 B.n5 163.367
R1020 B.n6 B.n5 163.367
R1021 B.n7 B.n6 163.367
R1022 B.n493 B.n7 163.367
R1023 B.n493 B.n12 163.367
R1024 B.n13 B.n12 163.367
R1025 B.n14 B.n13 163.367
R1026 B.n498 B.n14 163.367
R1027 B.n498 B.n19 163.367
R1028 B.n20 B.n19 163.367
R1029 B.n21 B.n20 163.367
R1030 B.n503 B.n21 163.367
R1031 B.n503 B.n26 163.367
R1032 B.n27 B.n26 163.367
R1033 B.n28 B.n27 163.367
R1034 B.n508 B.n28 163.367
R1035 B.n508 B.n33 163.367
R1036 B.n34 B.n33 163.367
R1037 B.n35 B.n34 163.367
R1038 B.n513 B.n35 163.367
R1039 B.n513 B.n40 163.367
R1040 B.n41 B.n40 163.367
R1041 B.n42 B.n41 163.367
R1042 B.n518 B.n42 163.367
R1043 B.n518 B.n47 163.367
R1044 B.n48 B.n47 163.367
R1045 B.n90 B.n89 163.367
R1046 B.n94 B.n93 163.367
R1047 B.n98 B.n97 163.367
R1048 B.n102 B.n101 163.367
R1049 B.n106 B.n105 163.367
R1050 B.n110 B.n109 163.367
R1051 B.n114 B.n113 163.367
R1052 B.n118 B.n117 163.367
R1053 B.n122 B.n121 163.367
R1054 B.n126 B.n125 163.367
R1055 B.n130 B.n129 163.367
R1056 B.n134 B.n133 163.367
R1057 B.n138 B.n137 163.367
R1058 B.n142 B.n141 163.367
R1059 B.n146 B.n145 163.367
R1060 B.n150 B.n149 163.367
R1061 B.n154 B.n153 163.367
R1062 B.n158 B.n157 163.367
R1063 B.n162 B.n161 163.367
R1064 B.n166 B.n165 163.367
R1065 B.n170 B.n169 163.367
R1066 B.n174 B.n173 163.367
R1067 B.n178 B.n177 163.367
R1068 B.n182 B.n181 163.367
R1069 B.n186 B.n185 163.367
R1070 B.n190 B.n189 163.367
R1071 B.n194 B.n193 163.367
R1072 B.n198 B.n197 163.367
R1073 B.n202 B.n201 163.367
R1074 B.n204 B.n79 163.367
R1075 B.n412 B.n252 105.111
R1076 B.n526 B.n525 105.111
R1077 B.n411 B.n410 71.676
R1078 B.n405 B.n256 71.676
R1079 B.n402 B.n257 71.676
R1080 B.n398 B.n258 71.676
R1081 B.n394 B.n259 71.676
R1082 B.n390 B.n260 71.676
R1083 B.n386 B.n261 71.676
R1084 B.n382 B.n262 71.676
R1085 B.n378 B.n263 71.676
R1086 B.n374 B.n264 71.676
R1087 B.n370 B.n265 71.676
R1088 B.n366 B.n266 71.676
R1089 B.n362 B.n267 71.676
R1090 B.n357 B.n268 71.676
R1091 B.n353 B.n269 71.676
R1092 B.n349 B.n270 71.676
R1093 B.n345 B.n271 71.676
R1094 B.n341 B.n272 71.676
R1095 B.n336 B.n273 71.676
R1096 B.n332 B.n274 71.676
R1097 B.n328 B.n275 71.676
R1098 B.n324 B.n276 71.676
R1099 B.n320 B.n277 71.676
R1100 B.n316 B.n278 71.676
R1101 B.n312 B.n279 71.676
R1102 B.n308 B.n280 71.676
R1103 B.n304 B.n281 71.676
R1104 B.n300 B.n282 71.676
R1105 B.n296 B.n283 71.676
R1106 B.n292 B.n284 71.676
R1107 B.n86 B.n49 71.676
R1108 B.n90 B.n50 71.676
R1109 B.n94 B.n51 71.676
R1110 B.n98 B.n52 71.676
R1111 B.n102 B.n53 71.676
R1112 B.n106 B.n54 71.676
R1113 B.n110 B.n55 71.676
R1114 B.n114 B.n56 71.676
R1115 B.n118 B.n57 71.676
R1116 B.n122 B.n58 71.676
R1117 B.n126 B.n59 71.676
R1118 B.n130 B.n60 71.676
R1119 B.n134 B.n61 71.676
R1120 B.n138 B.n62 71.676
R1121 B.n142 B.n63 71.676
R1122 B.n146 B.n64 71.676
R1123 B.n150 B.n65 71.676
R1124 B.n154 B.n66 71.676
R1125 B.n158 B.n67 71.676
R1126 B.n162 B.n68 71.676
R1127 B.n166 B.n69 71.676
R1128 B.n170 B.n70 71.676
R1129 B.n174 B.n71 71.676
R1130 B.n178 B.n72 71.676
R1131 B.n182 B.n73 71.676
R1132 B.n186 B.n74 71.676
R1133 B.n190 B.n75 71.676
R1134 B.n194 B.n76 71.676
R1135 B.n198 B.n77 71.676
R1136 B.n202 B.n78 71.676
R1137 B.n524 B.n79 71.676
R1138 B.n524 B.n523 71.676
R1139 B.n204 B.n78 71.676
R1140 B.n201 B.n77 71.676
R1141 B.n197 B.n76 71.676
R1142 B.n193 B.n75 71.676
R1143 B.n189 B.n74 71.676
R1144 B.n185 B.n73 71.676
R1145 B.n181 B.n72 71.676
R1146 B.n177 B.n71 71.676
R1147 B.n173 B.n70 71.676
R1148 B.n169 B.n69 71.676
R1149 B.n165 B.n68 71.676
R1150 B.n161 B.n67 71.676
R1151 B.n157 B.n66 71.676
R1152 B.n153 B.n65 71.676
R1153 B.n149 B.n64 71.676
R1154 B.n145 B.n63 71.676
R1155 B.n141 B.n62 71.676
R1156 B.n137 B.n61 71.676
R1157 B.n133 B.n60 71.676
R1158 B.n129 B.n59 71.676
R1159 B.n125 B.n58 71.676
R1160 B.n121 B.n57 71.676
R1161 B.n117 B.n56 71.676
R1162 B.n113 B.n55 71.676
R1163 B.n109 B.n54 71.676
R1164 B.n105 B.n53 71.676
R1165 B.n101 B.n52 71.676
R1166 B.n97 B.n51 71.676
R1167 B.n93 B.n50 71.676
R1168 B.n89 B.n49 71.676
R1169 B.n411 B.n286 71.676
R1170 B.n403 B.n256 71.676
R1171 B.n399 B.n257 71.676
R1172 B.n395 B.n258 71.676
R1173 B.n391 B.n259 71.676
R1174 B.n387 B.n260 71.676
R1175 B.n383 B.n261 71.676
R1176 B.n379 B.n262 71.676
R1177 B.n375 B.n263 71.676
R1178 B.n371 B.n264 71.676
R1179 B.n367 B.n265 71.676
R1180 B.n363 B.n266 71.676
R1181 B.n358 B.n267 71.676
R1182 B.n354 B.n268 71.676
R1183 B.n350 B.n269 71.676
R1184 B.n346 B.n270 71.676
R1185 B.n342 B.n271 71.676
R1186 B.n337 B.n272 71.676
R1187 B.n333 B.n273 71.676
R1188 B.n329 B.n274 71.676
R1189 B.n325 B.n275 71.676
R1190 B.n321 B.n276 71.676
R1191 B.n317 B.n277 71.676
R1192 B.n313 B.n278 71.676
R1193 B.n309 B.n279 71.676
R1194 B.n305 B.n280 71.676
R1195 B.n301 B.n281 71.676
R1196 B.n297 B.n282 71.676
R1197 B.n293 B.n283 71.676
R1198 B.n284 B.n255 71.676
R1199 B.n418 B.n252 62.1526
R1200 B.n418 B.n248 62.1526
R1201 B.n424 B.n248 62.1526
R1202 B.n424 B.n244 62.1526
R1203 B.n430 B.n244 62.1526
R1204 B.n436 B.n240 62.1526
R1205 B.n436 B.n236 62.1526
R1206 B.n442 B.n236 62.1526
R1207 B.n442 B.n232 62.1526
R1208 B.n448 B.n232 62.1526
R1209 B.n454 B.n228 62.1526
R1210 B.n454 B.n224 62.1526
R1211 B.n460 B.n224 62.1526
R1212 B.n467 B.n220 62.1526
R1213 B.n467 B.n466 62.1526
R1214 B.n473 B.n213 62.1526
R1215 B.n480 B.n213 62.1526
R1216 B.n486 B.n209 62.1526
R1217 B.n486 B.n4 62.1526
R1218 B.n575 B.n4 62.1526
R1219 B.n575 B.n574 62.1526
R1220 B.n574 B.n573 62.1526
R1221 B.n573 B.n8 62.1526
R1222 B.n567 B.n566 62.1526
R1223 B.n566 B.n565 62.1526
R1224 B.n559 B.n18 62.1526
R1225 B.n559 B.n558 62.1526
R1226 B.n557 B.n22 62.1526
R1227 B.n551 B.n22 62.1526
R1228 B.n551 B.n550 62.1526
R1229 B.n549 B.n29 62.1526
R1230 B.n543 B.n29 62.1526
R1231 B.n543 B.n542 62.1526
R1232 B.n542 B.n541 62.1526
R1233 B.n541 B.n36 62.1526
R1234 B.n535 B.n534 62.1526
R1235 B.n534 B.n533 62.1526
R1236 B.n533 B.n43 62.1526
R1237 B.n527 B.n43 62.1526
R1238 B.n527 B.n526 62.1526
R1239 B.t5 B.n220 61.2386
R1240 B.n558 B.t3 61.2386
R1241 B.n339 B.n290 59.5399
R1242 B.n360 B.n288 59.5399
R1243 B.n85 B.n84 59.5399
R1244 B.n82 B.n81 59.5399
R1245 B.t13 B.n240 55.7546
R1246 B.t9 B.n36 55.7546
R1247 B.n480 B.t7 44.7865
R1248 B.n567 B.t1 44.7865
R1249 B.n448 B.t4 41.1305
R1250 B.t0 B.n549 41.1305
R1251 B.n473 B.t2 39.3025
R1252 B.n565 B.t6 39.3025
R1253 B.n87 B.n45 31.0639
R1254 B.n522 B.n521 31.0639
R1255 B.n415 B.n414 31.0639
R1256 B.n409 B.n250 31.0639
R1257 B.n466 B.t2 22.8505
R1258 B.n18 B.t6 22.8505
R1259 B.n290 B.n289 22.1096
R1260 B.n288 B.n287 22.1096
R1261 B.n84 B.n83 22.1096
R1262 B.n81 B.n80 22.1096
R1263 B.t4 B.n228 21.0225
R1264 B.n550 B.t0 21.0225
R1265 B B.n577 18.0485
R1266 B.t7 B.n209 17.3665
R1267 B.t1 B.n8 17.3665
R1268 B.n88 B.n87 10.6151
R1269 B.n91 B.n88 10.6151
R1270 B.n92 B.n91 10.6151
R1271 B.n95 B.n92 10.6151
R1272 B.n96 B.n95 10.6151
R1273 B.n99 B.n96 10.6151
R1274 B.n100 B.n99 10.6151
R1275 B.n103 B.n100 10.6151
R1276 B.n104 B.n103 10.6151
R1277 B.n107 B.n104 10.6151
R1278 B.n108 B.n107 10.6151
R1279 B.n111 B.n108 10.6151
R1280 B.n112 B.n111 10.6151
R1281 B.n115 B.n112 10.6151
R1282 B.n116 B.n115 10.6151
R1283 B.n119 B.n116 10.6151
R1284 B.n120 B.n119 10.6151
R1285 B.n123 B.n120 10.6151
R1286 B.n124 B.n123 10.6151
R1287 B.n127 B.n124 10.6151
R1288 B.n128 B.n127 10.6151
R1289 B.n131 B.n128 10.6151
R1290 B.n132 B.n131 10.6151
R1291 B.n135 B.n132 10.6151
R1292 B.n136 B.n135 10.6151
R1293 B.n140 B.n139 10.6151
R1294 B.n143 B.n140 10.6151
R1295 B.n144 B.n143 10.6151
R1296 B.n147 B.n144 10.6151
R1297 B.n148 B.n147 10.6151
R1298 B.n151 B.n148 10.6151
R1299 B.n152 B.n151 10.6151
R1300 B.n155 B.n152 10.6151
R1301 B.n156 B.n155 10.6151
R1302 B.n160 B.n159 10.6151
R1303 B.n163 B.n160 10.6151
R1304 B.n164 B.n163 10.6151
R1305 B.n167 B.n164 10.6151
R1306 B.n168 B.n167 10.6151
R1307 B.n171 B.n168 10.6151
R1308 B.n172 B.n171 10.6151
R1309 B.n175 B.n172 10.6151
R1310 B.n176 B.n175 10.6151
R1311 B.n179 B.n176 10.6151
R1312 B.n180 B.n179 10.6151
R1313 B.n183 B.n180 10.6151
R1314 B.n184 B.n183 10.6151
R1315 B.n187 B.n184 10.6151
R1316 B.n188 B.n187 10.6151
R1317 B.n191 B.n188 10.6151
R1318 B.n192 B.n191 10.6151
R1319 B.n195 B.n192 10.6151
R1320 B.n196 B.n195 10.6151
R1321 B.n199 B.n196 10.6151
R1322 B.n200 B.n199 10.6151
R1323 B.n203 B.n200 10.6151
R1324 B.n205 B.n203 10.6151
R1325 B.n206 B.n205 10.6151
R1326 B.n522 B.n206 10.6151
R1327 B.n416 B.n415 10.6151
R1328 B.n416 B.n246 10.6151
R1329 B.n426 B.n246 10.6151
R1330 B.n427 B.n426 10.6151
R1331 B.n428 B.n427 10.6151
R1332 B.n428 B.n238 10.6151
R1333 B.n438 B.n238 10.6151
R1334 B.n439 B.n438 10.6151
R1335 B.n440 B.n439 10.6151
R1336 B.n440 B.n230 10.6151
R1337 B.n450 B.n230 10.6151
R1338 B.n451 B.n450 10.6151
R1339 B.n452 B.n451 10.6151
R1340 B.n452 B.n222 10.6151
R1341 B.n462 B.n222 10.6151
R1342 B.n463 B.n462 10.6151
R1343 B.n464 B.n463 10.6151
R1344 B.n464 B.n215 10.6151
R1345 B.n475 B.n215 10.6151
R1346 B.n476 B.n475 10.6151
R1347 B.n478 B.n476 10.6151
R1348 B.n478 B.n477 10.6151
R1349 B.n477 B.n207 10.6151
R1350 B.n489 B.n207 10.6151
R1351 B.n490 B.n489 10.6151
R1352 B.n491 B.n490 10.6151
R1353 B.n492 B.n491 10.6151
R1354 B.n494 B.n492 10.6151
R1355 B.n495 B.n494 10.6151
R1356 B.n496 B.n495 10.6151
R1357 B.n497 B.n496 10.6151
R1358 B.n499 B.n497 10.6151
R1359 B.n500 B.n499 10.6151
R1360 B.n501 B.n500 10.6151
R1361 B.n502 B.n501 10.6151
R1362 B.n504 B.n502 10.6151
R1363 B.n505 B.n504 10.6151
R1364 B.n506 B.n505 10.6151
R1365 B.n507 B.n506 10.6151
R1366 B.n509 B.n507 10.6151
R1367 B.n510 B.n509 10.6151
R1368 B.n511 B.n510 10.6151
R1369 B.n512 B.n511 10.6151
R1370 B.n514 B.n512 10.6151
R1371 B.n515 B.n514 10.6151
R1372 B.n516 B.n515 10.6151
R1373 B.n517 B.n516 10.6151
R1374 B.n519 B.n517 10.6151
R1375 B.n520 B.n519 10.6151
R1376 B.n521 B.n520 10.6151
R1377 B.n409 B.n408 10.6151
R1378 B.n408 B.n407 10.6151
R1379 B.n407 B.n406 10.6151
R1380 B.n406 B.n404 10.6151
R1381 B.n404 B.n401 10.6151
R1382 B.n401 B.n400 10.6151
R1383 B.n400 B.n397 10.6151
R1384 B.n397 B.n396 10.6151
R1385 B.n396 B.n393 10.6151
R1386 B.n393 B.n392 10.6151
R1387 B.n392 B.n389 10.6151
R1388 B.n389 B.n388 10.6151
R1389 B.n388 B.n385 10.6151
R1390 B.n385 B.n384 10.6151
R1391 B.n384 B.n381 10.6151
R1392 B.n381 B.n380 10.6151
R1393 B.n380 B.n377 10.6151
R1394 B.n377 B.n376 10.6151
R1395 B.n376 B.n373 10.6151
R1396 B.n373 B.n372 10.6151
R1397 B.n372 B.n369 10.6151
R1398 B.n369 B.n368 10.6151
R1399 B.n368 B.n365 10.6151
R1400 B.n365 B.n364 10.6151
R1401 B.n364 B.n361 10.6151
R1402 B.n359 B.n356 10.6151
R1403 B.n356 B.n355 10.6151
R1404 B.n355 B.n352 10.6151
R1405 B.n352 B.n351 10.6151
R1406 B.n351 B.n348 10.6151
R1407 B.n348 B.n347 10.6151
R1408 B.n347 B.n344 10.6151
R1409 B.n344 B.n343 10.6151
R1410 B.n343 B.n340 10.6151
R1411 B.n338 B.n335 10.6151
R1412 B.n335 B.n334 10.6151
R1413 B.n334 B.n331 10.6151
R1414 B.n331 B.n330 10.6151
R1415 B.n330 B.n327 10.6151
R1416 B.n327 B.n326 10.6151
R1417 B.n326 B.n323 10.6151
R1418 B.n323 B.n322 10.6151
R1419 B.n322 B.n319 10.6151
R1420 B.n319 B.n318 10.6151
R1421 B.n318 B.n315 10.6151
R1422 B.n315 B.n314 10.6151
R1423 B.n314 B.n311 10.6151
R1424 B.n311 B.n310 10.6151
R1425 B.n310 B.n307 10.6151
R1426 B.n307 B.n306 10.6151
R1427 B.n306 B.n303 10.6151
R1428 B.n303 B.n302 10.6151
R1429 B.n302 B.n299 10.6151
R1430 B.n299 B.n298 10.6151
R1431 B.n298 B.n295 10.6151
R1432 B.n295 B.n294 10.6151
R1433 B.n294 B.n291 10.6151
R1434 B.n291 B.n254 10.6151
R1435 B.n414 B.n254 10.6151
R1436 B.n420 B.n250 10.6151
R1437 B.n421 B.n420 10.6151
R1438 B.n422 B.n421 10.6151
R1439 B.n422 B.n242 10.6151
R1440 B.n432 B.n242 10.6151
R1441 B.n433 B.n432 10.6151
R1442 B.n434 B.n433 10.6151
R1443 B.n434 B.n234 10.6151
R1444 B.n444 B.n234 10.6151
R1445 B.n445 B.n444 10.6151
R1446 B.n446 B.n445 10.6151
R1447 B.n446 B.n226 10.6151
R1448 B.n456 B.n226 10.6151
R1449 B.n457 B.n456 10.6151
R1450 B.n458 B.n457 10.6151
R1451 B.n458 B.n218 10.6151
R1452 B.n469 B.n218 10.6151
R1453 B.n470 B.n469 10.6151
R1454 B.n471 B.n470 10.6151
R1455 B.n471 B.n211 10.6151
R1456 B.n482 B.n211 10.6151
R1457 B.n483 B.n482 10.6151
R1458 B.n484 B.n483 10.6151
R1459 B.n484 B.n0 10.6151
R1460 B.n571 B.n1 10.6151
R1461 B.n571 B.n570 10.6151
R1462 B.n570 B.n569 10.6151
R1463 B.n569 B.n10 10.6151
R1464 B.n563 B.n10 10.6151
R1465 B.n563 B.n562 10.6151
R1466 B.n562 B.n561 10.6151
R1467 B.n561 B.n16 10.6151
R1468 B.n555 B.n16 10.6151
R1469 B.n555 B.n554 10.6151
R1470 B.n554 B.n553 10.6151
R1471 B.n553 B.n24 10.6151
R1472 B.n547 B.n24 10.6151
R1473 B.n547 B.n546 10.6151
R1474 B.n546 B.n545 10.6151
R1475 B.n545 B.n31 10.6151
R1476 B.n539 B.n31 10.6151
R1477 B.n539 B.n538 10.6151
R1478 B.n538 B.n537 10.6151
R1479 B.n537 B.n38 10.6151
R1480 B.n531 B.n38 10.6151
R1481 B.n531 B.n530 10.6151
R1482 B.n530 B.n529 10.6151
R1483 B.n529 B.n45 10.6151
R1484 B.n136 B.n85 9.36635
R1485 B.n159 B.n82 9.36635
R1486 B.n361 B.n360 9.36635
R1487 B.n339 B.n338 9.36635
R1488 B.n430 B.t13 6.39851
R1489 B.n535 B.t9 6.39851
R1490 B.n577 B.n0 2.81026
R1491 B.n577 B.n1 2.81026
R1492 B.n139 B.n85 1.24928
R1493 B.n156 B.n82 1.24928
R1494 B.n360 B.n359 1.24928
R1495 B.n340 B.n339 1.24928
R1496 B.n460 B.t5 0.914501
R1497 B.t3 B.n557 0.914501
R1498 VN.n2 VN.t3 270.652
R1499 VN.n10 VN.t4 270.652
R1500 VN.n1 VN.t2 249.629
R1501 VN.n4 VN.t1 249.629
R1502 VN.n6 VN.t7 249.629
R1503 VN.n9 VN.t6 249.629
R1504 VN.n12 VN.t0 249.629
R1505 VN.n14 VN.t5 249.629
R1506 VN.n7 VN.n6 161.3
R1507 VN.n15 VN.n14 161.3
R1508 VN.n13 VN.n8 161.3
R1509 VN.n5 VN.n0 161.3
R1510 VN.n12 VN.n11 80.6037
R1511 VN.n4 VN.n3 80.6037
R1512 VN.n4 VN.n1 48.2005
R1513 VN.n12 VN.n9 48.2005
R1514 VN.n5 VN.n4 40.1672
R1515 VN.n13 VN.n12 40.1672
R1516 VN VN.n15 38.8812
R1517 VN.n11 VN.n10 31.6481
R1518 VN.n3 VN.n2 31.6481
R1519 VN.n2 VN.n1 17.444
R1520 VN.n10 VN.n9 17.444
R1521 VN.n6 VN.n5 8.03383
R1522 VN.n14 VN.n13 8.03383
R1523 VN.n11 VN.n8 0.285035
R1524 VN.n3 VN.n0 0.285035
R1525 VN.n15 VN.n8 0.189894
R1526 VN.n7 VN.n0 0.189894
R1527 VN VN.n7 0.0516364
R1528 VDD2.n2 VDD2.n1 67.2857
R1529 VDD2.n2 VDD2.n0 67.2857
R1530 VDD2 VDD2.n5 67.2829
R1531 VDD2.n4 VDD2.n3 66.8499
R1532 VDD2.n4 VDD2.n2 33.9653
R1533 VDD2.n5 VDD2.t1 2.92949
R1534 VDD2.n5 VDD2.t3 2.92949
R1535 VDD2.n3 VDD2.t2 2.92949
R1536 VDD2.n3 VDD2.t7 2.92949
R1537 VDD2.n1 VDD2.t6 2.92949
R1538 VDD2.n1 VDD2.t0 2.92949
R1539 VDD2.n0 VDD2.t4 2.92949
R1540 VDD2.n0 VDD2.t5 2.92949
R1541 VDD2 VDD2.n4 0.550069
C0 VN VDD1 0.148659f
C1 VDD2 VDD1 0.879662f
C2 VN VDD2 3.50913f
C3 VP VDD1 3.68934f
C4 VP VN 4.50197f
C5 VTAIL VDD1 6.83249f
C6 VP VDD2 0.329363f
C7 VN VTAIL 3.57871f
C8 VDD2 VTAIL 6.87491f
C9 VP VTAIL 3.59281f
C10 VDD2 B 3.182562f
C11 VDD1 B 3.427642f
C12 VTAIL B 5.921696f
C13 VN B 8.28264f
C14 VP B 6.623445f
C15 VDD2.t4 B 0.141245f
C16 VDD2.t5 B 0.141245f
C17 VDD2.n0 B 1.19693f
C18 VDD2.t6 B 0.141245f
C19 VDD2.t0 B 0.141245f
C20 VDD2.n1 B 1.19693f
C21 VDD2.n2 B 2.02984f
C22 VDD2.t2 B 0.141245f
C23 VDD2.t7 B 0.141245f
C24 VDD2.n3 B 1.19467f
C25 VDD2.n4 B 2.0254f
C26 VDD2.t1 B 0.141245f
C27 VDD2.t3 B 0.141245f
C28 VDD2.n5 B 1.19691f
C29 VN.n0 B 0.056932f
C30 VN.t2 B 0.675051f
C31 VN.n1 B 0.310944f
C32 VN.t3 B 0.698522f
C33 VN.n2 B 0.282518f
C34 VN.n3 B 0.245225f
C35 VN.t1 B 0.675051f
C36 VN.n4 B 0.310084f
C37 VN.n5 B 0.009682f
C38 VN.t7 B 0.675051f
C39 VN.n6 B 0.294615f
C40 VN.n7 B 0.033064f
C41 VN.n8 B 0.056932f
C42 VN.t6 B 0.675051f
C43 VN.n9 B 0.310944f
C44 VN.t0 B 0.675051f
C45 VN.t4 B 0.698522f
C46 VN.n10 B 0.282518f
C47 VN.n11 B 0.245225f
C48 VN.n12 B 0.310084f
C49 VN.n13 B 0.009682f
C50 VN.t5 B 0.675051f
C51 VN.n14 B 0.294615f
C52 VN.n15 B 1.54453f
C53 VDD1.t5 B 0.141276f
C54 VDD1.t4 B 0.141276f
C55 VDD1.n0 B 1.19786f
C56 VDD1.t2 B 0.141276f
C57 VDD1.t3 B 0.141276f
C58 VDD1.n1 B 1.1972f
C59 VDD1.t1 B 0.141276f
C60 VDD1.t7 B 0.141276f
C61 VDD1.n2 B 1.1972f
C62 VDD1.n3 B 2.08686f
C63 VDD1.t0 B 0.141276f
C64 VDD1.t6 B 0.141276f
C65 VDD1.n4 B 1.19493f
C66 VDD1.n5 B 2.05705f
C67 VTAIL.t13 B 0.113659f
C68 VTAIL.t3 B 0.113659f
C69 VTAIL.n0 B 0.904748f
C70 VTAIL.n1 B 0.273315f
C71 VTAIL.n2 B 0.031055f
C72 VTAIL.n3 B 0.021277f
C73 VTAIL.n4 B 0.011433f
C74 VTAIL.n5 B 0.027024f
C75 VTAIL.n6 B 0.012106f
C76 VTAIL.n7 B 0.021277f
C77 VTAIL.n8 B 0.011433f
C78 VTAIL.n9 B 0.027024f
C79 VTAIL.n10 B 0.012106f
C80 VTAIL.n11 B 0.580545f
C81 VTAIL.n12 B 0.011433f
C82 VTAIL.t1 B 0.044039f
C83 VTAIL.n13 B 0.094982f
C84 VTAIL.n14 B 0.015963f
C85 VTAIL.n15 B 0.020268f
C86 VTAIL.n16 B 0.027024f
C87 VTAIL.n17 B 0.012106f
C88 VTAIL.n18 B 0.011433f
C89 VTAIL.n19 B 0.021277f
C90 VTAIL.n20 B 0.021277f
C91 VTAIL.n21 B 0.011433f
C92 VTAIL.n22 B 0.012106f
C93 VTAIL.n23 B 0.027024f
C94 VTAIL.n24 B 0.027024f
C95 VTAIL.n25 B 0.012106f
C96 VTAIL.n26 B 0.011433f
C97 VTAIL.n27 B 0.021277f
C98 VTAIL.n28 B 0.021277f
C99 VTAIL.n29 B 0.011433f
C100 VTAIL.n30 B 0.012106f
C101 VTAIL.n31 B 0.027024f
C102 VTAIL.n32 B 0.060533f
C103 VTAIL.n33 B 0.012106f
C104 VTAIL.n34 B 0.011433f
C105 VTAIL.n35 B 0.050342f
C106 VTAIL.n36 B 0.034114f
C107 VTAIL.n37 B 0.118414f
C108 VTAIL.n38 B 0.031055f
C109 VTAIL.n39 B 0.021277f
C110 VTAIL.n40 B 0.011433f
C111 VTAIL.n41 B 0.027024f
C112 VTAIL.n42 B 0.012106f
C113 VTAIL.n43 B 0.021277f
C114 VTAIL.n44 B 0.011433f
C115 VTAIL.n45 B 0.027024f
C116 VTAIL.n46 B 0.012106f
C117 VTAIL.n47 B 0.580545f
C118 VTAIL.n48 B 0.011433f
C119 VTAIL.t11 B 0.044039f
C120 VTAIL.n49 B 0.094982f
C121 VTAIL.n50 B 0.015963f
C122 VTAIL.n51 B 0.020268f
C123 VTAIL.n52 B 0.027024f
C124 VTAIL.n53 B 0.012106f
C125 VTAIL.n54 B 0.011433f
C126 VTAIL.n55 B 0.021277f
C127 VTAIL.n56 B 0.021277f
C128 VTAIL.n57 B 0.011433f
C129 VTAIL.n58 B 0.012106f
C130 VTAIL.n59 B 0.027024f
C131 VTAIL.n60 B 0.027024f
C132 VTAIL.n61 B 0.012106f
C133 VTAIL.n62 B 0.011433f
C134 VTAIL.n63 B 0.021277f
C135 VTAIL.n64 B 0.021277f
C136 VTAIL.n65 B 0.011433f
C137 VTAIL.n66 B 0.012106f
C138 VTAIL.n67 B 0.027024f
C139 VTAIL.n68 B 0.060533f
C140 VTAIL.n69 B 0.012106f
C141 VTAIL.n70 B 0.011433f
C142 VTAIL.n71 B 0.050342f
C143 VTAIL.n72 B 0.034114f
C144 VTAIL.n73 B 0.118414f
C145 VTAIL.t5 B 0.113659f
C146 VTAIL.t8 B 0.113659f
C147 VTAIL.n74 B 0.904748f
C148 VTAIL.n75 B 0.336702f
C149 VTAIL.n76 B 0.031055f
C150 VTAIL.n77 B 0.021277f
C151 VTAIL.n78 B 0.011433f
C152 VTAIL.n79 B 0.027024f
C153 VTAIL.n80 B 0.012106f
C154 VTAIL.n81 B 0.021277f
C155 VTAIL.n82 B 0.011433f
C156 VTAIL.n83 B 0.027024f
C157 VTAIL.n84 B 0.012106f
C158 VTAIL.n85 B 0.580545f
C159 VTAIL.n86 B 0.011433f
C160 VTAIL.t4 B 0.044039f
C161 VTAIL.n87 B 0.094982f
C162 VTAIL.n88 B 0.015963f
C163 VTAIL.n89 B 0.020268f
C164 VTAIL.n90 B 0.027024f
C165 VTAIL.n91 B 0.012106f
C166 VTAIL.n92 B 0.011433f
C167 VTAIL.n93 B 0.021277f
C168 VTAIL.n94 B 0.021277f
C169 VTAIL.n95 B 0.011433f
C170 VTAIL.n96 B 0.012106f
C171 VTAIL.n97 B 0.027024f
C172 VTAIL.n98 B 0.027024f
C173 VTAIL.n99 B 0.012106f
C174 VTAIL.n100 B 0.011433f
C175 VTAIL.n101 B 0.021277f
C176 VTAIL.n102 B 0.021277f
C177 VTAIL.n103 B 0.011433f
C178 VTAIL.n104 B 0.012106f
C179 VTAIL.n105 B 0.027024f
C180 VTAIL.n106 B 0.060533f
C181 VTAIL.n107 B 0.012106f
C182 VTAIL.n108 B 0.011433f
C183 VTAIL.n109 B 0.050342f
C184 VTAIL.n110 B 0.034114f
C185 VTAIL.n111 B 0.842124f
C186 VTAIL.n112 B 0.031055f
C187 VTAIL.n113 B 0.021277f
C188 VTAIL.n114 B 0.011433f
C189 VTAIL.n115 B 0.027024f
C190 VTAIL.n116 B 0.012106f
C191 VTAIL.n117 B 0.021277f
C192 VTAIL.n118 B 0.011433f
C193 VTAIL.n119 B 0.027024f
C194 VTAIL.n120 B 0.012106f
C195 VTAIL.n121 B 0.580545f
C196 VTAIL.n122 B 0.011433f
C197 VTAIL.t15 B 0.044039f
C198 VTAIL.n123 B 0.094982f
C199 VTAIL.n124 B 0.015963f
C200 VTAIL.n125 B 0.020268f
C201 VTAIL.n126 B 0.027024f
C202 VTAIL.n127 B 0.012106f
C203 VTAIL.n128 B 0.011433f
C204 VTAIL.n129 B 0.021277f
C205 VTAIL.n130 B 0.021277f
C206 VTAIL.n131 B 0.011433f
C207 VTAIL.n132 B 0.012106f
C208 VTAIL.n133 B 0.027024f
C209 VTAIL.n134 B 0.027024f
C210 VTAIL.n135 B 0.012106f
C211 VTAIL.n136 B 0.011433f
C212 VTAIL.n137 B 0.021277f
C213 VTAIL.n138 B 0.021277f
C214 VTAIL.n139 B 0.011433f
C215 VTAIL.n140 B 0.012106f
C216 VTAIL.n141 B 0.027024f
C217 VTAIL.n142 B 0.060533f
C218 VTAIL.n143 B 0.012106f
C219 VTAIL.n144 B 0.011433f
C220 VTAIL.n145 B 0.050342f
C221 VTAIL.n146 B 0.034114f
C222 VTAIL.n147 B 0.842124f
C223 VTAIL.t12 B 0.113659f
C224 VTAIL.t2 B 0.113659f
C225 VTAIL.n148 B 0.904754f
C226 VTAIL.n149 B 0.336696f
C227 VTAIL.n150 B 0.031055f
C228 VTAIL.n151 B 0.021277f
C229 VTAIL.n152 B 0.011433f
C230 VTAIL.n153 B 0.027024f
C231 VTAIL.n154 B 0.012106f
C232 VTAIL.n155 B 0.021277f
C233 VTAIL.n156 B 0.011433f
C234 VTAIL.n157 B 0.027024f
C235 VTAIL.n158 B 0.012106f
C236 VTAIL.n159 B 0.580545f
C237 VTAIL.n160 B 0.011433f
C238 VTAIL.t14 B 0.044039f
C239 VTAIL.n161 B 0.094982f
C240 VTAIL.n162 B 0.015963f
C241 VTAIL.n163 B 0.020268f
C242 VTAIL.n164 B 0.027024f
C243 VTAIL.n165 B 0.012106f
C244 VTAIL.n166 B 0.011433f
C245 VTAIL.n167 B 0.021277f
C246 VTAIL.n168 B 0.021277f
C247 VTAIL.n169 B 0.011433f
C248 VTAIL.n170 B 0.012106f
C249 VTAIL.n171 B 0.027024f
C250 VTAIL.n172 B 0.027024f
C251 VTAIL.n173 B 0.012106f
C252 VTAIL.n174 B 0.011433f
C253 VTAIL.n175 B 0.021277f
C254 VTAIL.n176 B 0.021277f
C255 VTAIL.n177 B 0.011433f
C256 VTAIL.n178 B 0.012106f
C257 VTAIL.n179 B 0.027024f
C258 VTAIL.n180 B 0.060533f
C259 VTAIL.n181 B 0.012106f
C260 VTAIL.n182 B 0.011433f
C261 VTAIL.n183 B 0.050342f
C262 VTAIL.n184 B 0.034114f
C263 VTAIL.n185 B 0.118414f
C264 VTAIL.n186 B 0.031055f
C265 VTAIL.n187 B 0.021277f
C266 VTAIL.n188 B 0.011433f
C267 VTAIL.n189 B 0.027024f
C268 VTAIL.n190 B 0.012106f
C269 VTAIL.n191 B 0.021277f
C270 VTAIL.n192 B 0.011433f
C271 VTAIL.n193 B 0.027024f
C272 VTAIL.n194 B 0.012106f
C273 VTAIL.n195 B 0.580545f
C274 VTAIL.n196 B 0.011433f
C275 VTAIL.t9 B 0.044039f
C276 VTAIL.n197 B 0.094982f
C277 VTAIL.n198 B 0.015963f
C278 VTAIL.n199 B 0.020268f
C279 VTAIL.n200 B 0.027024f
C280 VTAIL.n201 B 0.012106f
C281 VTAIL.n202 B 0.011433f
C282 VTAIL.n203 B 0.021277f
C283 VTAIL.n204 B 0.021277f
C284 VTAIL.n205 B 0.011433f
C285 VTAIL.n206 B 0.012106f
C286 VTAIL.n207 B 0.027024f
C287 VTAIL.n208 B 0.027024f
C288 VTAIL.n209 B 0.012106f
C289 VTAIL.n210 B 0.011433f
C290 VTAIL.n211 B 0.021277f
C291 VTAIL.n212 B 0.021277f
C292 VTAIL.n213 B 0.011433f
C293 VTAIL.n214 B 0.012106f
C294 VTAIL.n215 B 0.027024f
C295 VTAIL.n216 B 0.060533f
C296 VTAIL.n217 B 0.012106f
C297 VTAIL.n218 B 0.011433f
C298 VTAIL.n219 B 0.050342f
C299 VTAIL.n220 B 0.034114f
C300 VTAIL.n221 B 0.118414f
C301 VTAIL.t7 B 0.113659f
C302 VTAIL.t6 B 0.113659f
C303 VTAIL.n222 B 0.904754f
C304 VTAIL.n223 B 0.336696f
C305 VTAIL.n224 B 0.031055f
C306 VTAIL.n225 B 0.021277f
C307 VTAIL.n226 B 0.011433f
C308 VTAIL.n227 B 0.027024f
C309 VTAIL.n228 B 0.012106f
C310 VTAIL.n229 B 0.021277f
C311 VTAIL.n230 B 0.011433f
C312 VTAIL.n231 B 0.027024f
C313 VTAIL.n232 B 0.012106f
C314 VTAIL.n233 B 0.580545f
C315 VTAIL.n234 B 0.011433f
C316 VTAIL.t10 B 0.044039f
C317 VTAIL.n235 B 0.094982f
C318 VTAIL.n236 B 0.015963f
C319 VTAIL.n237 B 0.020268f
C320 VTAIL.n238 B 0.027024f
C321 VTAIL.n239 B 0.012106f
C322 VTAIL.n240 B 0.011433f
C323 VTAIL.n241 B 0.021277f
C324 VTAIL.n242 B 0.021277f
C325 VTAIL.n243 B 0.011433f
C326 VTAIL.n244 B 0.012106f
C327 VTAIL.n245 B 0.027024f
C328 VTAIL.n246 B 0.027024f
C329 VTAIL.n247 B 0.012106f
C330 VTAIL.n248 B 0.011433f
C331 VTAIL.n249 B 0.021277f
C332 VTAIL.n250 B 0.021277f
C333 VTAIL.n251 B 0.011433f
C334 VTAIL.n252 B 0.012106f
C335 VTAIL.n253 B 0.027024f
C336 VTAIL.n254 B 0.060533f
C337 VTAIL.n255 B 0.012106f
C338 VTAIL.n256 B 0.011433f
C339 VTAIL.n257 B 0.050342f
C340 VTAIL.n258 B 0.034114f
C341 VTAIL.n259 B 0.842124f
C342 VTAIL.n260 B 0.031055f
C343 VTAIL.n261 B 0.021277f
C344 VTAIL.n262 B 0.011433f
C345 VTAIL.n263 B 0.027024f
C346 VTAIL.n264 B 0.012106f
C347 VTAIL.n265 B 0.021277f
C348 VTAIL.n266 B 0.011433f
C349 VTAIL.n267 B 0.027024f
C350 VTAIL.n268 B 0.012106f
C351 VTAIL.n269 B 0.580545f
C352 VTAIL.n270 B 0.011433f
C353 VTAIL.t0 B 0.044039f
C354 VTAIL.n271 B 0.094982f
C355 VTAIL.n272 B 0.015963f
C356 VTAIL.n273 B 0.020268f
C357 VTAIL.n274 B 0.027024f
C358 VTAIL.n275 B 0.012106f
C359 VTAIL.n276 B 0.011433f
C360 VTAIL.n277 B 0.021277f
C361 VTAIL.n278 B 0.021277f
C362 VTAIL.n279 B 0.011433f
C363 VTAIL.n280 B 0.012106f
C364 VTAIL.n281 B 0.027024f
C365 VTAIL.n282 B 0.027024f
C366 VTAIL.n283 B 0.012106f
C367 VTAIL.n284 B 0.011433f
C368 VTAIL.n285 B 0.021277f
C369 VTAIL.n286 B 0.021277f
C370 VTAIL.n287 B 0.011433f
C371 VTAIL.n288 B 0.012106f
C372 VTAIL.n289 B 0.027024f
C373 VTAIL.n290 B 0.060533f
C374 VTAIL.n291 B 0.012106f
C375 VTAIL.n292 B 0.011433f
C376 VTAIL.n293 B 0.050342f
C377 VTAIL.n294 B 0.034114f
C378 VTAIL.n295 B 0.838134f
C379 VP.n0 B 0.058215f
C380 VP.t4 B 0.690259f
C381 VP.n1 B 0.317069f
C382 VP.n2 B 0.058215f
C383 VP.t1 B 0.690259f
C384 VP.t7 B 0.690259f
C385 VP.n3 B 0.25075f
C386 VP.t3 B 0.690259f
C387 VP.t2 B 0.714258f
C388 VP.n4 B 0.288882f
C389 VP.n5 B 0.317949f
C390 VP.n6 B 0.317069f
C391 VP.n7 B 0.0099f
C392 VP.n8 B 0.301252f
C393 VP.n9 B 1.55052f
C394 VP.n10 B 1.59137f
C395 VP.t5 B 0.690259f
C396 VP.n11 B 0.301252f
C397 VP.n12 B 0.0099f
C398 VP.n13 B 0.058215f
C399 VP.n14 B 0.072666f
C400 VP.n15 B 0.072666f
C401 VP.t6 B 0.690259f
C402 VP.n16 B 0.317069f
C403 VP.n17 B 0.0099f
C404 VP.t0 B 0.690259f
C405 VP.n18 B 0.301252f
C406 VP.n19 B 0.033809f
.ends

