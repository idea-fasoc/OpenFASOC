* NGSPICE file created from diff_pair_sample_1713.ext - technology: sky130A

.subckt diff_pair_sample_1713 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n1542_n3676# sky130_fd_pr__pfet_01v8 ad=5.2728 pd=27.82 as=0 ps=0 w=13.52 l=1.1
X1 VDD2.t1 VN.t0 VTAIL.t2 w_n1542_n3676# sky130_fd_pr__pfet_01v8 ad=5.2728 pd=27.82 as=5.2728 ps=27.82 w=13.52 l=1.1
X2 B.t8 B.t6 B.t7 w_n1542_n3676# sky130_fd_pr__pfet_01v8 ad=5.2728 pd=27.82 as=0 ps=0 w=13.52 l=1.1
X3 VDD1.t1 VP.t0 VTAIL.t0 w_n1542_n3676# sky130_fd_pr__pfet_01v8 ad=5.2728 pd=27.82 as=5.2728 ps=27.82 w=13.52 l=1.1
X4 VDD1.t0 VP.t1 VTAIL.t1 w_n1542_n3676# sky130_fd_pr__pfet_01v8 ad=5.2728 pd=27.82 as=5.2728 ps=27.82 w=13.52 l=1.1
X5 B.t5 B.t3 B.t4 w_n1542_n3676# sky130_fd_pr__pfet_01v8 ad=5.2728 pd=27.82 as=0 ps=0 w=13.52 l=1.1
X6 VDD2.t0 VN.t1 VTAIL.t3 w_n1542_n3676# sky130_fd_pr__pfet_01v8 ad=5.2728 pd=27.82 as=5.2728 ps=27.82 w=13.52 l=1.1
X7 B.t2 B.t0 B.t1 w_n1542_n3676# sky130_fd_pr__pfet_01v8 ad=5.2728 pd=27.82 as=0 ps=0 w=13.52 l=1.1
R0 B.n322 B.n321 585
R1 B.n320 B.n83 585
R2 B.n319 B.n318 585
R3 B.n317 B.n84 585
R4 B.n316 B.n315 585
R5 B.n314 B.n85 585
R6 B.n313 B.n312 585
R7 B.n311 B.n86 585
R8 B.n310 B.n309 585
R9 B.n308 B.n87 585
R10 B.n307 B.n306 585
R11 B.n305 B.n88 585
R12 B.n304 B.n303 585
R13 B.n302 B.n89 585
R14 B.n301 B.n300 585
R15 B.n299 B.n90 585
R16 B.n298 B.n297 585
R17 B.n296 B.n91 585
R18 B.n295 B.n294 585
R19 B.n293 B.n92 585
R20 B.n292 B.n291 585
R21 B.n290 B.n93 585
R22 B.n289 B.n288 585
R23 B.n287 B.n94 585
R24 B.n286 B.n285 585
R25 B.n284 B.n95 585
R26 B.n283 B.n282 585
R27 B.n281 B.n96 585
R28 B.n280 B.n279 585
R29 B.n278 B.n97 585
R30 B.n277 B.n276 585
R31 B.n275 B.n98 585
R32 B.n274 B.n273 585
R33 B.n272 B.n99 585
R34 B.n271 B.n270 585
R35 B.n269 B.n100 585
R36 B.n268 B.n267 585
R37 B.n266 B.n101 585
R38 B.n265 B.n264 585
R39 B.n263 B.n102 585
R40 B.n262 B.n261 585
R41 B.n260 B.n103 585
R42 B.n259 B.n258 585
R43 B.n257 B.n104 585
R44 B.n256 B.n255 585
R45 B.n254 B.n105 585
R46 B.n252 B.n251 585
R47 B.n250 B.n108 585
R48 B.n249 B.n248 585
R49 B.n247 B.n109 585
R50 B.n246 B.n245 585
R51 B.n244 B.n110 585
R52 B.n243 B.n242 585
R53 B.n241 B.n111 585
R54 B.n240 B.n239 585
R55 B.n238 B.n112 585
R56 B.n237 B.n236 585
R57 B.n232 B.n113 585
R58 B.n231 B.n230 585
R59 B.n229 B.n114 585
R60 B.n228 B.n227 585
R61 B.n226 B.n115 585
R62 B.n225 B.n224 585
R63 B.n223 B.n116 585
R64 B.n222 B.n221 585
R65 B.n220 B.n117 585
R66 B.n219 B.n218 585
R67 B.n217 B.n118 585
R68 B.n216 B.n215 585
R69 B.n214 B.n119 585
R70 B.n213 B.n212 585
R71 B.n211 B.n120 585
R72 B.n210 B.n209 585
R73 B.n208 B.n121 585
R74 B.n207 B.n206 585
R75 B.n205 B.n122 585
R76 B.n204 B.n203 585
R77 B.n202 B.n123 585
R78 B.n201 B.n200 585
R79 B.n199 B.n124 585
R80 B.n198 B.n197 585
R81 B.n196 B.n125 585
R82 B.n195 B.n194 585
R83 B.n193 B.n126 585
R84 B.n192 B.n191 585
R85 B.n190 B.n127 585
R86 B.n189 B.n188 585
R87 B.n187 B.n128 585
R88 B.n186 B.n185 585
R89 B.n184 B.n129 585
R90 B.n183 B.n182 585
R91 B.n181 B.n130 585
R92 B.n180 B.n179 585
R93 B.n178 B.n131 585
R94 B.n177 B.n176 585
R95 B.n175 B.n132 585
R96 B.n174 B.n173 585
R97 B.n172 B.n133 585
R98 B.n171 B.n170 585
R99 B.n169 B.n134 585
R100 B.n168 B.n167 585
R101 B.n166 B.n135 585
R102 B.n323 B.n82 585
R103 B.n325 B.n324 585
R104 B.n326 B.n81 585
R105 B.n328 B.n327 585
R106 B.n329 B.n80 585
R107 B.n331 B.n330 585
R108 B.n332 B.n79 585
R109 B.n334 B.n333 585
R110 B.n335 B.n78 585
R111 B.n337 B.n336 585
R112 B.n338 B.n77 585
R113 B.n340 B.n339 585
R114 B.n341 B.n76 585
R115 B.n343 B.n342 585
R116 B.n344 B.n75 585
R117 B.n346 B.n345 585
R118 B.n347 B.n74 585
R119 B.n349 B.n348 585
R120 B.n350 B.n73 585
R121 B.n352 B.n351 585
R122 B.n353 B.n72 585
R123 B.n355 B.n354 585
R124 B.n356 B.n71 585
R125 B.n358 B.n357 585
R126 B.n359 B.n70 585
R127 B.n361 B.n360 585
R128 B.n362 B.n69 585
R129 B.n364 B.n363 585
R130 B.n365 B.n68 585
R131 B.n367 B.n366 585
R132 B.n368 B.n67 585
R133 B.n370 B.n369 585
R134 B.n371 B.n66 585
R135 B.n373 B.n372 585
R136 B.n527 B.n10 585
R137 B.n526 B.n525 585
R138 B.n524 B.n11 585
R139 B.n523 B.n522 585
R140 B.n521 B.n12 585
R141 B.n520 B.n519 585
R142 B.n518 B.n13 585
R143 B.n517 B.n516 585
R144 B.n515 B.n14 585
R145 B.n514 B.n513 585
R146 B.n512 B.n15 585
R147 B.n511 B.n510 585
R148 B.n509 B.n16 585
R149 B.n508 B.n507 585
R150 B.n506 B.n17 585
R151 B.n505 B.n504 585
R152 B.n503 B.n18 585
R153 B.n502 B.n501 585
R154 B.n500 B.n19 585
R155 B.n499 B.n498 585
R156 B.n497 B.n20 585
R157 B.n496 B.n495 585
R158 B.n494 B.n21 585
R159 B.n493 B.n492 585
R160 B.n491 B.n22 585
R161 B.n490 B.n489 585
R162 B.n488 B.n23 585
R163 B.n487 B.n486 585
R164 B.n485 B.n24 585
R165 B.n484 B.n483 585
R166 B.n482 B.n25 585
R167 B.n481 B.n480 585
R168 B.n479 B.n26 585
R169 B.n478 B.n477 585
R170 B.n476 B.n27 585
R171 B.n475 B.n474 585
R172 B.n473 B.n28 585
R173 B.n472 B.n471 585
R174 B.n470 B.n29 585
R175 B.n469 B.n468 585
R176 B.n467 B.n30 585
R177 B.n466 B.n465 585
R178 B.n464 B.n31 585
R179 B.n463 B.n462 585
R180 B.n461 B.n32 585
R181 B.n460 B.n459 585
R182 B.n457 B.n33 585
R183 B.n456 B.n455 585
R184 B.n454 B.n36 585
R185 B.n453 B.n452 585
R186 B.n451 B.n37 585
R187 B.n450 B.n449 585
R188 B.n448 B.n38 585
R189 B.n447 B.n446 585
R190 B.n445 B.n39 585
R191 B.n444 B.n443 585
R192 B.n442 B.n441 585
R193 B.n440 B.n43 585
R194 B.n439 B.n438 585
R195 B.n437 B.n44 585
R196 B.n436 B.n435 585
R197 B.n434 B.n45 585
R198 B.n433 B.n432 585
R199 B.n431 B.n46 585
R200 B.n430 B.n429 585
R201 B.n428 B.n47 585
R202 B.n427 B.n426 585
R203 B.n425 B.n48 585
R204 B.n424 B.n423 585
R205 B.n422 B.n49 585
R206 B.n421 B.n420 585
R207 B.n419 B.n50 585
R208 B.n418 B.n417 585
R209 B.n416 B.n51 585
R210 B.n415 B.n414 585
R211 B.n413 B.n52 585
R212 B.n412 B.n411 585
R213 B.n410 B.n53 585
R214 B.n409 B.n408 585
R215 B.n407 B.n54 585
R216 B.n406 B.n405 585
R217 B.n404 B.n55 585
R218 B.n403 B.n402 585
R219 B.n401 B.n56 585
R220 B.n400 B.n399 585
R221 B.n398 B.n57 585
R222 B.n397 B.n396 585
R223 B.n395 B.n58 585
R224 B.n394 B.n393 585
R225 B.n392 B.n59 585
R226 B.n391 B.n390 585
R227 B.n389 B.n60 585
R228 B.n388 B.n387 585
R229 B.n386 B.n61 585
R230 B.n385 B.n384 585
R231 B.n383 B.n62 585
R232 B.n382 B.n381 585
R233 B.n380 B.n63 585
R234 B.n379 B.n378 585
R235 B.n377 B.n64 585
R236 B.n376 B.n375 585
R237 B.n374 B.n65 585
R238 B.n529 B.n528 585
R239 B.n530 B.n9 585
R240 B.n532 B.n531 585
R241 B.n533 B.n8 585
R242 B.n535 B.n534 585
R243 B.n536 B.n7 585
R244 B.n538 B.n537 585
R245 B.n539 B.n6 585
R246 B.n541 B.n540 585
R247 B.n542 B.n5 585
R248 B.n544 B.n543 585
R249 B.n545 B.n4 585
R250 B.n547 B.n546 585
R251 B.n548 B.n3 585
R252 B.n550 B.n549 585
R253 B.n551 B.n0 585
R254 B.n2 B.n1 585
R255 B.n144 B.n143 585
R256 B.n145 B.n142 585
R257 B.n147 B.n146 585
R258 B.n148 B.n141 585
R259 B.n150 B.n149 585
R260 B.n151 B.n140 585
R261 B.n153 B.n152 585
R262 B.n154 B.n139 585
R263 B.n156 B.n155 585
R264 B.n157 B.n138 585
R265 B.n159 B.n158 585
R266 B.n160 B.n137 585
R267 B.n162 B.n161 585
R268 B.n163 B.n136 585
R269 B.n165 B.n164 585
R270 B.n233 B.t3 499.772
R271 B.n106 B.t6 499.772
R272 B.n40 B.t0 499.772
R273 B.n34 B.t9 499.772
R274 B.n164 B.n135 492.5
R275 B.n323 B.n322 492.5
R276 B.n372 B.n65 492.5
R277 B.n528 B.n527 492.5
R278 B.n106 B.t7 430.861
R279 B.n40 B.t2 430.861
R280 B.n233 B.t4 430.861
R281 B.n34 B.t11 430.861
R282 B.n107 B.t8 403.127
R283 B.n41 B.t1 403.127
R284 B.n234 B.t5 403.127
R285 B.n35 B.t10 403.127
R286 B.n553 B.n552 256.663
R287 B.n552 B.n551 235.042
R288 B.n552 B.n2 235.042
R289 B.n168 B.n135 163.367
R290 B.n169 B.n168 163.367
R291 B.n170 B.n169 163.367
R292 B.n170 B.n133 163.367
R293 B.n174 B.n133 163.367
R294 B.n175 B.n174 163.367
R295 B.n176 B.n175 163.367
R296 B.n176 B.n131 163.367
R297 B.n180 B.n131 163.367
R298 B.n181 B.n180 163.367
R299 B.n182 B.n181 163.367
R300 B.n182 B.n129 163.367
R301 B.n186 B.n129 163.367
R302 B.n187 B.n186 163.367
R303 B.n188 B.n187 163.367
R304 B.n188 B.n127 163.367
R305 B.n192 B.n127 163.367
R306 B.n193 B.n192 163.367
R307 B.n194 B.n193 163.367
R308 B.n194 B.n125 163.367
R309 B.n198 B.n125 163.367
R310 B.n199 B.n198 163.367
R311 B.n200 B.n199 163.367
R312 B.n200 B.n123 163.367
R313 B.n204 B.n123 163.367
R314 B.n205 B.n204 163.367
R315 B.n206 B.n205 163.367
R316 B.n206 B.n121 163.367
R317 B.n210 B.n121 163.367
R318 B.n211 B.n210 163.367
R319 B.n212 B.n211 163.367
R320 B.n212 B.n119 163.367
R321 B.n216 B.n119 163.367
R322 B.n217 B.n216 163.367
R323 B.n218 B.n217 163.367
R324 B.n218 B.n117 163.367
R325 B.n222 B.n117 163.367
R326 B.n223 B.n222 163.367
R327 B.n224 B.n223 163.367
R328 B.n224 B.n115 163.367
R329 B.n228 B.n115 163.367
R330 B.n229 B.n228 163.367
R331 B.n230 B.n229 163.367
R332 B.n230 B.n113 163.367
R333 B.n237 B.n113 163.367
R334 B.n238 B.n237 163.367
R335 B.n239 B.n238 163.367
R336 B.n239 B.n111 163.367
R337 B.n243 B.n111 163.367
R338 B.n244 B.n243 163.367
R339 B.n245 B.n244 163.367
R340 B.n245 B.n109 163.367
R341 B.n249 B.n109 163.367
R342 B.n250 B.n249 163.367
R343 B.n251 B.n250 163.367
R344 B.n251 B.n105 163.367
R345 B.n256 B.n105 163.367
R346 B.n257 B.n256 163.367
R347 B.n258 B.n257 163.367
R348 B.n258 B.n103 163.367
R349 B.n262 B.n103 163.367
R350 B.n263 B.n262 163.367
R351 B.n264 B.n263 163.367
R352 B.n264 B.n101 163.367
R353 B.n268 B.n101 163.367
R354 B.n269 B.n268 163.367
R355 B.n270 B.n269 163.367
R356 B.n270 B.n99 163.367
R357 B.n274 B.n99 163.367
R358 B.n275 B.n274 163.367
R359 B.n276 B.n275 163.367
R360 B.n276 B.n97 163.367
R361 B.n280 B.n97 163.367
R362 B.n281 B.n280 163.367
R363 B.n282 B.n281 163.367
R364 B.n282 B.n95 163.367
R365 B.n286 B.n95 163.367
R366 B.n287 B.n286 163.367
R367 B.n288 B.n287 163.367
R368 B.n288 B.n93 163.367
R369 B.n292 B.n93 163.367
R370 B.n293 B.n292 163.367
R371 B.n294 B.n293 163.367
R372 B.n294 B.n91 163.367
R373 B.n298 B.n91 163.367
R374 B.n299 B.n298 163.367
R375 B.n300 B.n299 163.367
R376 B.n300 B.n89 163.367
R377 B.n304 B.n89 163.367
R378 B.n305 B.n304 163.367
R379 B.n306 B.n305 163.367
R380 B.n306 B.n87 163.367
R381 B.n310 B.n87 163.367
R382 B.n311 B.n310 163.367
R383 B.n312 B.n311 163.367
R384 B.n312 B.n85 163.367
R385 B.n316 B.n85 163.367
R386 B.n317 B.n316 163.367
R387 B.n318 B.n317 163.367
R388 B.n318 B.n83 163.367
R389 B.n322 B.n83 163.367
R390 B.n372 B.n371 163.367
R391 B.n371 B.n370 163.367
R392 B.n370 B.n67 163.367
R393 B.n366 B.n67 163.367
R394 B.n366 B.n365 163.367
R395 B.n365 B.n364 163.367
R396 B.n364 B.n69 163.367
R397 B.n360 B.n69 163.367
R398 B.n360 B.n359 163.367
R399 B.n359 B.n358 163.367
R400 B.n358 B.n71 163.367
R401 B.n354 B.n71 163.367
R402 B.n354 B.n353 163.367
R403 B.n353 B.n352 163.367
R404 B.n352 B.n73 163.367
R405 B.n348 B.n73 163.367
R406 B.n348 B.n347 163.367
R407 B.n347 B.n346 163.367
R408 B.n346 B.n75 163.367
R409 B.n342 B.n75 163.367
R410 B.n342 B.n341 163.367
R411 B.n341 B.n340 163.367
R412 B.n340 B.n77 163.367
R413 B.n336 B.n77 163.367
R414 B.n336 B.n335 163.367
R415 B.n335 B.n334 163.367
R416 B.n334 B.n79 163.367
R417 B.n330 B.n79 163.367
R418 B.n330 B.n329 163.367
R419 B.n329 B.n328 163.367
R420 B.n328 B.n81 163.367
R421 B.n324 B.n81 163.367
R422 B.n324 B.n323 163.367
R423 B.n527 B.n526 163.367
R424 B.n526 B.n11 163.367
R425 B.n522 B.n11 163.367
R426 B.n522 B.n521 163.367
R427 B.n521 B.n520 163.367
R428 B.n520 B.n13 163.367
R429 B.n516 B.n13 163.367
R430 B.n516 B.n515 163.367
R431 B.n515 B.n514 163.367
R432 B.n514 B.n15 163.367
R433 B.n510 B.n15 163.367
R434 B.n510 B.n509 163.367
R435 B.n509 B.n508 163.367
R436 B.n508 B.n17 163.367
R437 B.n504 B.n17 163.367
R438 B.n504 B.n503 163.367
R439 B.n503 B.n502 163.367
R440 B.n502 B.n19 163.367
R441 B.n498 B.n19 163.367
R442 B.n498 B.n497 163.367
R443 B.n497 B.n496 163.367
R444 B.n496 B.n21 163.367
R445 B.n492 B.n21 163.367
R446 B.n492 B.n491 163.367
R447 B.n491 B.n490 163.367
R448 B.n490 B.n23 163.367
R449 B.n486 B.n23 163.367
R450 B.n486 B.n485 163.367
R451 B.n485 B.n484 163.367
R452 B.n484 B.n25 163.367
R453 B.n480 B.n25 163.367
R454 B.n480 B.n479 163.367
R455 B.n479 B.n478 163.367
R456 B.n478 B.n27 163.367
R457 B.n474 B.n27 163.367
R458 B.n474 B.n473 163.367
R459 B.n473 B.n472 163.367
R460 B.n472 B.n29 163.367
R461 B.n468 B.n29 163.367
R462 B.n468 B.n467 163.367
R463 B.n467 B.n466 163.367
R464 B.n466 B.n31 163.367
R465 B.n462 B.n31 163.367
R466 B.n462 B.n461 163.367
R467 B.n461 B.n460 163.367
R468 B.n460 B.n33 163.367
R469 B.n455 B.n33 163.367
R470 B.n455 B.n454 163.367
R471 B.n454 B.n453 163.367
R472 B.n453 B.n37 163.367
R473 B.n449 B.n37 163.367
R474 B.n449 B.n448 163.367
R475 B.n448 B.n447 163.367
R476 B.n447 B.n39 163.367
R477 B.n443 B.n39 163.367
R478 B.n443 B.n442 163.367
R479 B.n442 B.n43 163.367
R480 B.n438 B.n43 163.367
R481 B.n438 B.n437 163.367
R482 B.n437 B.n436 163.367
R483 B.n436 B.n45 163.367
R484 B.n432 B.n45 163.367
R485 B.n432 B.n431 163.367
R486 B.n431 B.n430 163.367
R487 B.n430 B.n47 163.367
R488 B.n426 B.n47 163.367
R489 B.n426 B.n425 163.367
R490 B.n425 B.n424 163.367
R491 B.n424 B.n49 163.367
R492 B.n420 B.n49 163.367
R493 B.n420 B.n419 163.367
R494 B.n419 B.n418 163.367
R495 B.n418 B.n51 163.367
R496 B.n414 B.n51 163.367
R497 B.n414 B.n413 163.367
R498 B.n413 B.n412 163.367
R499 B.n412 B.n53 163.367
R500 B.n408 B.n53 163.367
R501 B.n408 B.n407 163.367
R502 B.n407 B.n406 163.367
R503 B.n406 B.n55 163.367
R504 B.n402 B.n55 163.367
R505 B.n402 B.n401 163.367
R506 B.n401 B.n400 163.367
R507 B.n400 B.n57 163.367
R508 B.n396 B.n57 163.367
R509 B.n396 B.n395 163.367
R510 B.n395 B.n394 163.367
R511 B.n394 B.n59 163.367
R512 B.n390 B.n59 163.367
R513 B.n390 B.n389 163.367
R514 B.n389 B.n388 163.367
R515 B.n388 B.n61 163.367
R516 B.n384 B.n61 163.367
R517 B.n384 B.n383 163.367
R518 B.n383 B.n382 163.367
R519 B.n382 B.n63 163.367
R520 B.n378 B.n63 163.367
R521 B.n378 B.n377 163.367
R522 B.n377 B.n376 163.367
R523 B.n376 B.n65 163.367
R524 B.n528 B.n9 163.367
R525 B.n532 B.n9 163.367
R526 B.n533 B.n532 163.367
R527 B.n534 B.n533 163.367
R528 B.n534 B.n7 163.367
R529 B.n538 B.n7 163.367
R530 B.n539 B.n538 163.367
R531 B.n540 B.n539 163.367
R532 B.n540 B.n5 163.367
R533 B.n544 B.n5 163.367
R534 B.n545 B.n544 163.367
R535 B.n546 B.n545 163.367
R536 B.n546 B.n3 163.367
R537 B.n550 B.n3 163.367
R538 B.n551 B.n550 163.367
R539 B.n144 B.n2 163.367
R540 B.n145 B.n144 163.367
R541 B.n146 B.n145 163.367
R542 B.n146 B.n141 163.367
R543 B.n150 B.n141 163.367
R544 B.n151 B.n150 163.367
R545 B.n152 B.n151 163.367
R546 B.n152 B.n139 163.367
R547 B.n156 B.n139 163.367
R548 B.n157 B.n156 163.367
R549 B.n158 B.n157 163.367
R550 B.n158 B.n137 163.367
R551 B.n162 B.n137 163.367
R552 B.n163 B.n162 163.367
R553 B.n164 B.n163 163.367
R554 B.n235 B.n234 59.5399
R555 B.n253 B.n107 59.5399
R556 B.n42 B.n41 59.5399
R557 B.n458 B.n35 59.5399
R558 B.n529 B.n10 32.0005
R559 B.n374 B.n373 32.0005
R560 B.n321 B.n82 32.0005
R561 B.n166 B.n165 32.0005
R562 B.n234 B.n233 27.7338
R563 B.n107 B.n106 27.7338
R564 B.n41 B.n40 27.7338
R565 B.n35 B.n34 27.7338
R566 B B.n553 18.0485
R567 B.n530 B.n529 10.6151
R568 B.n531 B.n530 10.6151
R569 B.n531 B.n8 10.6151
R570 B.n535 B.n8 10.6151
R571 B.n536 B.n535 10.6151
R572 B.n537 B.n536 10.6151
R573 B.n537 B.n6 10.6151
R574 B.n541 B.n6 10.6151
R575 B.n542 B.n541 10.6151
R576 B.n543 B.n542 10.6151
R577 B.n543 B.n4 10.6151
R578 B.n547 B.n4 10.6151
R579 B.n548 B.n547 10.6151
R580 B.n549 B.n548 10.6151
R581 B.n549 B.n0 10.6151
R582 B.n525 B.n10 10.6151
R583 B.n525 B.n524 10.6151
R584 B.n524 B.n523 10.6151
R585 B.n523 B.n12 10.6151
R586 B.n519 B.n12 10.6151
R587 B.n519 B.n518 10.6151
R588 B.n518 B.n517 10.6151
R589 B.n517 B.n14 10.6151
R590 B.n513 B.n14 10.6151
R591 B.n513 B.n512 10.6151
R592 B.n512 B.n511 10.6151
R593 B.n511 B.n16 10.6151
R594 B.n507 B.n16 10.6151
R595 B.n507 B.n506 10.6151
R596 B.n506 B.n505 10.6151
R597 B.n505 B.n18 10.6151
R598 B.n501 B.n18 10.6151
R599 B.n501 B.n500 10.6151
R600 B.n500 B.n499 10.6151
R601 B.n499 B.n20 10.6151
R602 B.n495 B.n20 10.6151
R603 B.n495 B.n494 10.6151
R604 B.n494 B.n493 10.6151
R605 B.n493 B.n22 10.6151
R606 B.n489 B.n22 10.6151
R607 B.n489 B.n488 10.6151
R608 B.n488 B.n487 10.6151
R609 B.n487 B.n24 10.6151
R610 B.n483 B.n24 10.6151
R611 B.n483 B.n482 10.6151
R612 B.n482 B.n481 10.6151
R613 B.n481 B.n26 10.6151
R614 B.n477 B.n26 10.6151
R615 B.n477 B.n476 10.6151
R616 B.n476 B.n475 10.6151
R617 B.n475 B.n28 10.6151
R618 B.n471 B.n28 10.6151
R619 B.n471 B.n470 10.6151
R620 B.n470 B.n469 10.6151
R621 B.n469 B.n30 10.6151
R622 B.n465 B.n30 10.6151
R623 B.n465 B.n464 10.6151
R624 B.n464 B.n463 10.6151
R625 B.n463 B.n32 10.6151
R626 B.n459 B.n32 10.6151
R627 B.n457 B.n456 10.6151
R628 B.n456 B.n36 10.6151
R629 B.n452 B.n36 10.6151
R630 B.n452 B.n451 10.6151
R631 B.n451 B.n450 10.6151
R632 B.n450 B.n38 10.6151
R633 B.n446 B.n38 10.6151
R634 B.n446 B.n445 10.6151
R635 B.n445 B.n444 10.6151
R636 B.n441 B.n440 10.6151
R637 B.n440 B.n439 10.6151
R638 B.n439 B.n44 10.6151
R639 B.n435 B.n44 10.6151
R640 B.n435 B.n434 10.6151
R641 B.n434 B.n433 10.6151
R642 B.n433 B.n46 10.6151
R643 B.n429 B.n46 10.6151
R644 B.n429 B.n428 10.6151
R645 B.n428 B.n427 10.6151
R646 B.n427 B.n48 10.6151
R647 B.n423 B.n48 10.6151
R648 B.n423 B.n422 10.6151
R649 B.n422 B.n421 10.6151
R650 B.n421 B.n50 10.6151
R651 B.n417 B.n50 10.6151
R652 B.n417 B.n416 10.6151
R653 B.n416 B.n415 10.6151
R654 B.n415 B.n52 10.6151
R655 B.n411 B.n52 10.6151
R656 B.n411 B.n410 10.6151
R657 B.n410 B.n409 10.6151
R658 B.n409 B.n54 10.6151
R659 B.n405 B.n54 10.6151
R660 B.n405 B.n404 10.6151
R661 B.n404 B.n403 10.6151
R662 B.n403 B.n56 10.6151
R663 B.n399 B.n56 10.6151
R664 B.n399 B.n398 10.6151
R665 B.n398 B.n397 10.6151
R666 B.n397 B.n58 10.6151
R667 B.n393 B.n58 10.6151
R668 B.n393 B.n392 10.6151
R669 B.n392 B.n391 10.6151
R670 B.n391 B.n60 10.6151
R671 B.n387 B.n60 10.6151
R672 B.n387 B.n386 10.6151
R673 B.n386 B.n385 10.6151
R674 B.n385 B.n62 10.6151
R675 B.n381 B.n62 10.6151
R676 B.n381 B.n380 10.6151
R677 B.n380 B.n379 10.6151
R678 B.n379 B.n64 10.6151
R679 B.n375 B.n64 10.6151
R680 B.n375 B.n374 10.6151
R681 B.n373 B.n66 10.6151
R682 B.n369 B.n66 10.6151
R683 B.n369 B.n368 10.6151
R684 B.n368 B.n367 10.6151
R685 B.n367 B.n68 10.6151
R686 B.n363 B.n68 10.6151
R687 B.n363 B.n362 10.6151
R688 B.n362 B.n361 10.6151
R689 B.n361 B.n70 10.6151
R690 B.n357 B.n70 10.6151
R691 B.n357 B.n356 10.6151
R692 B.n356 B.n355 10.6151
R693 B.n355 B.n72 10.6151
R694 B.n351 B.n72 10.6151
R695 B.n351 B.n350 10.6151
R696 B.n350 B.n349 10.6151
R697 B.n349 B.n74 10.6151
R698 B.n345 B.n74 10.6151
R699 B.n345 B.n344 10.6151
R700 B.n344 B.n343 10.6151
R701 B.n343 B.n76 10.6151
R702 B.n339 B.n76 10.6151
R703 B.n339 B.n338 10.6151
R704 B.n338 B.n337 10.6151
R705 B.n337 B.n78 10.6151
R706 B.n333 B.n78 10.6151
R707 B.n333 B.n332 10.6151
R708 B.n332 B.n331 10.6151
R709 B.n331 B.n80 10.6151
R710 B.n327 B.n80 10.6151
R711 B.n327 B.n326 10.6151
R712 B.n326 B.n325 10.6151
R713 B.n325 B.n82 10.6151
R714 B.n143 B.n1 10.6151
R715 B.n143 B.n142 10.6151
R716 B.n147 B.n142 10.6151
R717 B.n148 B.n147 10.6151
R718 B.n149 B.n148 10.6151
R719 B.n149 B.n140 10.6151
R720 B.n153 B.n140 10.6151
R721 B.n154 B.n153 10.6151
R722 B.n155 B.n154 10.6151
R723 B.n155 B.n138 10.6151
R724 B.n159 B.n138 10.6151
R725 B.n160 B.n159 10.6151
R726 B.n161 B.n160 10.6151
R727 B.n161 B.n136 10.6151
R728 B.n165 B.n136 10.6151
R729 B.n167 B.n166 10.6151
R730 B.n167 B.n134 10.6151
R731 B.n171 B.n134 10.6151
R732 B.n172 B.n171 10.6151
R733 B.n173 B.n172 10.6151
R734 B.n173 B.n132 10.6151
R735 B.n177 B.n132 10.6151
R736 B.n178 B.n177 10.6151
R737 B.n179 B.n178 10.6151
R738 B.n179 B.n130 10.6151
R739 B.n183 B.n130 10.6151
R740 B.n184 B.n183 10.6151
R741 B.n185 B.n184 10.6151
R742 B.n185 B.n128 10.6151
R743 B.n189 B.n128 10.6151
R744 B.n190 B.n189 10.6151
R745 B.n191 B.n190 10.6151
R746 B.n191 B.n126 10.6151
R747 B.n195 B.n126 10.6151
R748 B.n196 B.n195 10.6151
R749 B.n197 B.n196 10.6151
R750 B.n197 B.n124 10.6151
R751 B.n201 B.n124 10.6151
R752 B.n202 B.n201 10.6151
R753 B.n203 B.n202 10.6151
R754 B.n203 B.n122 10.6151
R755 B.n207 B.n122 10.6151
R756 B.n208 B.n207 10.6151
R757 B.n209 B.n208 10.6151
R758 B.n209 B.n120 10.6151
R759 B.n213 B.n120 10.6151
R760 B.n214 B.n213 10.6151
R761 B.n215 B.n214 10.6151
R762 B.n215 B.n118 10.6151
R763 B.n219 B.n118 10.6151
R764 B.n220 B.n219 10.6151
R765 B.n221 B.n220 10.6151
R766 B.n221 B.n116 10.6151
R767 B.n225 B.n116 10.6151
R768 B.n226 B.n225 10.6151
R769 B.n227 B.n226 10.6151
R770 B.n227 B.n114 10.6151
R771 B.n231 B.n114 10.6151
R772 B.n232 B.n231 10.6151
R773 B.n236 B.n232 10.6151
R774 B.n240 B.n112 10.6151
R775 B.n241 B.n240 10.6151
R776 B.n242 B.n241 10.6151
R777 B.n242 B.n110 10.6151
R778 B.n246 B.n110 10.6151
R779 B.n247 B.n246 10.6151
R780 B.n248 B.n247 10.6151
R781 B.n248 B.n108 10.6151
R782 B.n252 B.n108 10.6151
R783 B.n255 B.n254 10.6151
R784 B.n255 B.n104 10.6151
R785 B.n259 B.n104 10.6151
R786 B.n260 B.n259 10.6151
R787 B.n261 B.n260 10.6151
R788 B.n261 B.n102 10.6151
R789 B.n265 B.n102 10.6151
R790 B.n266 B.n265 10.6151
R791 B.n267 B.n266 10.6151
R792 B.n267 B.n100 10.6151
R793 B.n271 B.n100 10.6151
R794 B.n272 B.n271 10.6151
R795 B.n273 B.n272 10.6151
R796 B.n273 B.n98 10.6151
R797 B.n277 B.n98 10.6151
R798 B.n278 B.n277 10.6151
R799 B.n279 B.n278 10.6151
R800 B.n279 B.n96 10.6151
R801 B.n283 B.n96 10.6151
R802 B.n284 B.n283 10.6151
R803 B.n285 B.n284 10.6151
R804 B.n285 B.n94 10.6151
R805 B.n289 B.n94 10.6151
R806 B.n290 B.n289 10.6151
R807 B.n291 B.n290 10.6151
R808 B.n291 B.n92 10.6151
R809 B.n295 B.n92 10.6151
R810 B.n296 B.n295 10.6151
R811 B.n297 B.n296 10.6151
R812 B.n297 B.n90 10.6151
R813 B.n301 B.n90 10.6151
R814 B.n302 B.n301 10.6151
R815 B.n303 B.n302 10.6151
R816 B.n303 B.n88 10.6151
R817 B.n307 B.n88 10.6151
R818 B.n308 B.n307 10.6151
R819 B.n309 B.n308 10.6151
R820 B.n309 B.n86 10.6151
R821 B.n313 B.n86 10.6151
R822 B.n314 B.n313 10.6151
R823 B.n315 B.n314 10.6151
R824 B.n315 B.n84 10.6151
R825 B.n319 B.n84 10.6151
R826 B.n320 B.n319 10.6151
R827 B.n321 B.n320 10.6151
R828 B.n459 B.n458 8.74196
R829 B.n441 B.n42 8.74196
R830 B.n236 B.n235 8.74196
R831 B.n254 B.n253 8.74196
R832 B.n553 B.n0 8.11757
R833 B.n553 B.n1 8.11757
R834 B.n458 B.n457 1.87367
R835 B.n444 B.n42 1.87367
R836 B.n235 B.n112 1.87367
R837 B.n253 B.n252 1.87367
R838 VN VN.t1 535.448
R839 VN VN.t0 493.274
R840 VTAIL.n290 VTAIL.n222 756.745
R841 VTAIL.n68 VTAIL.n0 756.745
R842 VTAIL.n216 VTAIL.n148 756.745
R843 VTAIL.n142 VTAIL.n74 756.745
R844 VTAIL.n247 VTAIL.n246 585
R845 VTAIL.n249 VTAIL.n248 585
R846 VTAIL.n242 VTAIL.n241 585
R847 VTAIL.n255 VTAIL.n254 585
R848 VTAIL.n257 VTAIL.n256 585
R849 VTAIL.n238 VTAIL.n237 585
R850 VTAIL.n264 VTAIL.n263 585
R851 VTAIL.n265 VTAIL.n236 585
R852 VTAIL.n267 VTAIL.n266 585
R853 VTAIL.n234 VTAIL.n233 585
R854 VTAIL.n273 VTAIL.n272 585
R855 VTAIL.n275 VTAIL.n274 585
R856 VTAIL.n230 VTAIL.n229 585
R857 VTAIL.n281 VTAIL.n280 585
R858 VTAIL.n283 VTAIL.n282 585
R859 VTAIL.n226 VTAIL.n225 585
R860 VTAIL.n289 VTAIL.n288 585
R861 VTAIL.n291 VTAIL.n290 585
R862 VTAIL.n25 VTAIL.n24 585
R863 VTAIL.n27 VTAIL.n26 585
R864 VTAIL.n20 VTAIL.n19 585
R865 VTAIL.n33 VTAIL.n32 585
R866 VTAIL.n35 VTAIL.n34 585
R867 VTAIL.n16 VTAIL.n15 585
R868 VTAIL.n42 VTAIL.n41 585
R869 VTAIL.n43 VTAIL.n14 585
R870 VTAIL.n45 VTAIL.n44 585
R871 VTAIL.n12 VTAIL.n11 585
R872 VTAIL.n51 VTAIL.n50 585
R873 VTAIL.n53 VTAIL.n52 585
R874 VTAIL.n8 VTAIL.n7 585
R875 VTAIL.n59 VTAIL.n58 585
R876 VTAIL.n61 VTAIL.n60 585
R877 VTAIL.n4 VTAIL.n3 585
R878 VTAIL.n67 VTAIL.n66 585
R879 VTAIL.n69 VTAIL.n68 585
R880 VTAIL.n217 VTAIL.n216 585
R881 VTAIL.n215 VTAIL.n214 585
R882 VTAIL.n152 VTAIL.n151 585
R883 VTAIL.n209 VTAIL.n208 585
R884 VTAIL.n207 VTAIL.n206 585
R885 VTAIL.n156 VTAIL.n155 585
R886 VTAIL.n201 VTAIL.n200 585
R887 VTAIL.n199 VTAIL.n198 585
R888 VTAIL.n160 VTAIL.n159 585
R889 VTAIL.n164 VTAIL.n162 585
R890 VTAIL.n193 VTAIL.n192 585
R891 VTAIL.n191 VTAIL.n190 585
R892 VTAIL.n166 VTAIL.n165 585
R893 VTAIL.n185 VTAIL.n184 585
R894 VTAIL.n183 VTAIL.n182 585
R895 VTAIL.n170 VTAIL.n169 585
R896 VTAIL.n177 VTAIL.n176 585
R897 VTAIL.n175 VTAIL.n174 585
R898 VTAIL.n143 VTAIL.n142 585
R899 VTAIL.n141 VTAIL.n140 585
R900 VTAIL.n78 VTAIL.n77 585
R901 VTAIL.n135 VTAIL.n134 585
R902 VTAIL.n133 VTAIL.n132 585
R903 VTAIL.n82 VTAIL.n81 585
R904 VTAIL.n127 VTAIL.n126 585
R905 VTAIL.n125 VTAIL.n124 585
R906 VTAIL.n86 VTAIL.n85 585
R907 VTAIL.n90 VTAIL.n88 585
R908 VTAIL.n119 VTAIL.n118 585
R909 VTAIL.n117 VTAIL.n116 585
R910 VTAIL.n92 VTAIL.n91 585
R911 VTAIL.n111 VTAIL.n110 585
R912 VTAIL.n109 VTAIL.n108 585
R913 VTAIL.n96 VTAIL.n95 585
R914 VTAIL.n103 VTAIL.n102 585
R915 VTAIL.n101 VTAIL.n100 585
R916 VTAIL.n245 VTAIL.t2 329.036
R917 VTAIL.n23 VTAIL.t0 329.036
R918 VTAIL.n173 VTAIL.t1 329.036
R919 VTAIL.n99 VTAIL.t3 329.036
R920 VTAIL.n248 VTAIL.n247 171.744
R921 VTAIL.n248 VTAIL.n241 171.744
R922 VTAIL.n255 VTAIL.n241 171.744
R923 VTAIL.n256 VTAIL.n255 171.744
R924 VTAIL.n256 VTAIL.n237 171.744
R925 VTAIL.n264 VTAIL.n237 171.744
R926 VTAIL.n265 VTAIL.n264 171.744
R927 VTAIL.n266 VTAIL.n265 171.744
R928 VTAIL.n266 VTAIL.n233 171.744
R929 VTAIL.n273 VTAIL.n233 171.744
R930 VTAIL.n274 VTAIL.n273 171.744
R931 VTAIL.n274 VTAIL.n229 171.744
R932 VTAIL.n281 VTAIL.n229 171.744
R933 VTAIL.n282 VTAIL.n281 171.744
R934 VTAIL.n282 VTAIL.n225 171.744
R935 VTAIL.n289 VTAIL.n225 171.744
R936 VTAIL.n290 VTAIL.n289 171.744
R937 VTAIL.n26 VTAIL.n25 171.744
R938 VTAIL.n26 VTAIL.n19 171.744
R939 VTAIL.n33 VTAIL.n19 171.744
R940 VTAIL.n34 VTAIL.n33 171.744
R941 VTAIL.n34 VTAIL.n15 171.744
R942 VTAIL.n42 VTAIL.n15 171.744
R943 VTAIL.n43 VTAIL.n42 171.744
R944 VTAIL.n44 VTAIL.n43 171.744
R945 VTAIL.n44 VTAIL.n11 171.744
R946 VTAIL.n51 VTAIL.n11 171.744
R947 VTAIL.n52 VTAIL.n51 171.744
R948 VTAIL.n52 VTAIL.n7 171.744
R949 VTAIL.n59 VTAIL.n7 171.744
R950 VTAIL.n60 VTAIL.n59 171.744
R951 VTAIL.n60 VTAIL.n3 171.744
R952 VTAIL.n67 VTAIL.n3 171.744
R953 VTAIL.n68 VTAIL.n67 171.744
R954 VTAIL.n216 VTAIL.n215 171.744
R955 VTAIL.n215 VTAIL.n151 171.744
R956 VTAIL.n208 VTAIL.n151 171.744
R957 VTAIL.n208 VTAIL.n207 171.744
R958 VTAIL.n207 VTAIL.n155 171.744
R959 VTAIL.n200 VTAIL.n155 171.744
R960 VTAIL.n200 VTAIL.n199 171.744
R961 VTAIL.n199 VTAIL.n159 171.744
R962 VTAIL.n164 VTAIL.n159 171.744
R963 VTAIL.n192 VTAIL.n164 171.744
R964 VTAIL.n192 VTAIL.n191 171.744
R965 VTAIL.n191 VTAIL.n165 171.744
R966 VTAIL.n184 VTAIL.n165 171.744
R967 VTAIL.n184 VTAIL.n183 171.744
R968 VTAIL.n183 VTAIL.n169 171.744
R969 VTAIL.n176 VTAIL.n169 171.744
R970 VTAIL.n176 VTAIL.n175 171.744
R971 VTAIL.n142 VTAIL.n141 171.744
R972 VTAIL.n141 VTAIL.n77 171.744
R973 VTAIL.n134 VTAIL.n77 171.744
R974 VTAIL.n134 VTAIL.n133 171.744
R975 VTAIL.n133 VTAIL.n81 171.744
R976 VTAIL.n126 VTAIL.n81 171.744
R977 VTAIL.n126 VTAIL.n125 171.744
R978 VTAIL.n125 VTAIL.n85 171.744
R979 VTAIL.n90 VTAIL.n85 171.744
R980 VTAIL.n118 VTAIL.n90 171.744
R981 VTAIL.n118 VTAIL.n117 171.744
R982 VTAIL.n117 VTAIL.n91 171.744
R983 VTAIL.n110 VTAIL.n91 171.744
R984 VTAIL.n110 VTAIL.n109 171.744
R985 VTAIL.n109 VTAIL.n95 171.744
R986 VTAIL.n102 VTAIL.n95 171.744
R987 VTAIL.n102 VTAIL.n101 171.744
R988 VTAIL.n247 VTAIL.t2 85.8723
R989 VTAIL.n25 VTAIL.t0 85.8723
R990 VTAIL.n175 VTAIL.t1 85.8723
R991 VTAIL.n101 VTAIL.t3 85.8723
R992 VTAIL.n295 VTAIL.n294 31.4096
R993 VTAIL.n73 VTAIL.n72 31.4096
R994 VTAIL.n221 VTAIL.n220 31.4096
R995 VTAIL.n147 VTAIL.n146 31.4096
R996 VTAIL.n147 VTAIL.n73 26.5048
R997 VTAIL.n295 VTAIL.n221 25.2721
R998 VTAIL.n267 VTAIL.n234 13.1884
R999 VTAIL.n45 VTAIL.n12 13.1884
R1000 VTAIL.n162 VTAIL.n160 13.1884
R1001 VTAIL.n88 VTAIL.n86 13.1884
R1002 VTAIL.n268 VTAIL.n236 12.8005
R1003 VTAIL.n272 VTAIL.n271 12.8005
R1004 VTAIL.n46 VTAIL.n14 12.8005
R1005 VTAIL.n50 VTAIL.n49 12.8005
R1006 VTAIL.n198 VTAIL.n197 12.8005
R1007 VTAIL.n194 VTAIL.n193 12.8005
R1008 VTAIL.n124 VTAIL.n123 12.8005
R1009 VTAIL.n120 VTAIL.n119 12.8005
R1010 VTAIL.n263 VTAIL.n262 12.0247
R1011 VTAIL.n275 VTAIL.n232 12.0247
R1012 VTAIL.n41 VTAIL.n40 12.0247
R1013 VTAIL.n53 VTAIL.n10 12.0247
R1014 VTAIL.n201 VTAIL.n158 12.0247
R1015 VTAIL.n190 VTAIL.n163 12.0247
R1016 VTAIL.n127 VTAIL.n84 12.0247
R1017 VTAIL.n116 VTAIL.n89 12.0247
R1018 VTAIL.n261 VTAIL.n238 11.249
R1019 VTAIL.n276 VTAIL.n230 11.249
R1020 VTAIL.n39 VTAIL.n16 11.249
R1021 VTAIL.n54 VTAIL.n8 11.249
R1022 VTAIL.n202 VTAIL.n156 11.249
R1023 VTAIL.n189 VTAIL.n166 11.249
R1024 VTAIL.n128 VTAIL.n82 11.249
R1025 VTAIL.n115 VTAIL.n92 11.249
R1026 VTAIL.n246 VTAIL.n245 10.7239
R1027 VTAIL.n24 VTAIL.n23 10.7239
R1028 VTAIL.n174 VTAIL.n173 10.7239
R1029 VTAIL.n100 VTAIL.n99 10.7239
R1030 VTAIL.n258 VTAIL.n257 10.4732
R1031 VTAIL.n280 VTAIL.n279 10.4732
R1032 VTAIL.n36 VTAIL.n35 10.4732
R1033 VTAIL.n58 VTAIL.n57 10.4732
R1034 VTAIL.n206 VTAIL.n205 10.4732
R1035 VTAIL.n186 VTAIL.n185 10.4732
R1036 VTAIL.n132 VTAIL.n131 10.4732
R1037 VTAIL.n112 VTAIL.n111 10.4732
R1038 VTAIL.n254 VTAIL.n240 9.69747
R1039 VTAIL.n283 VTAIL.n228 9.69747
R1040 VTAIL.n32 VTAIL.n18 9.69747
R1041 VTAIL.n61 VTAIL.n6 9.69747
R1042 VTAIL.n209 VTAIL.n154 9.69747
R1043 VTAIL.n182 VTAIL.n168 9.69747
R1044 VTAIL.n135 VTAIL.n80 9.69747
R1045 VTAIL.n108 VTAIL.n94 9.69747
R1046 VTAIL.n294 VTAIL.n293 9.45567
R1047 VTAIL.n72 VTAIL.n71 9.45567
R1048 VTAIL.n220 VTAIL.n219 9.45567
R1049 VTAIL.n146 VTAIL.n145 9.45567
R1050 VTAIL.n293 VTAIL.n292 9.3005
R1051 VTAIL.n287 VTAIL.n286 9.3005
R1052 VTAIL.n285 VTAIL.n284 9.3005
R1053 VTAIL.n228 VTAIL.n227 9.3005
R1054 VTAIL.n279 VTAIL.n278 9.3005
R1055 VTAIL.n277 VTAIL.n276 9.3005
R1056 VTAIL.n232 VTAIL.n231 9.3005
R1057 VTAIL.n271 VTAIL.n270 9.3005
R1058 VTAIL.n244 VTAIL.n243 9.3005
R1059 VTAIL.n251 VTAIL.n250 9.3005
R1060 VTAIL.n253 VTAIL.n252 9.3005
R1061 VTAIL.n240 VTAIL.n239 9.3005
R1062 VTAIL.n259 VTAIL.n258 9.3005
R1063 VTAIL.n261 VTAIL.n260 9.3005
R1064 VTAIL.n262 VTAIL.n235 9.3005
R1065 VTAIL.n269 VTAIL.n268 9.3005
R1066 VTAIL.n224 VTAIL.n223 9.3005
R1067 VTAIL.n71 VTAIL.n70 9.3005
R1068 VTAIL.n65 VTAIL.n64 9.3005
R1069 VTAIL.n63 VTAIL.n62 9.3005
R1070 VTAIL.n6 VTAIL.n5 9.3005
R1071 VTAIL.n57 VTAIL.n56 9.3005
R1072 VTAIL.n55 VTAIL.n54 9.3005
R1073 VTAIL.n10 VTAIL.n9 9.3005
R1074 VTAIL.n49 VTAIL.n48 9.3005
R1075 VTAIL.n22 VTAIL.n21 9.3005
R1076 VTAIL.n29 VTAIL.n28 9.3005
R1077 VTAIL.n31 VTAIL.n30 9.3005
R1078 VTAIL.n18 VTAIL.n17 9.3005
R1079 VTAIL.n37 VTAIL.n36 9.3005
R1080 VTAIL.n39 VTAIL.n38 9.3005
R1081 VTAIL.n40 VTAIL.n13 9.3005
R1082 VTAIL.n47 VTAIL.n46 9.3005
R1083 VTAIL.n2 VTAIL.n1 9.3005
R1084 VTAIL.n172 VTAIL.n171 9.3005
R1085 VTAIL.n179 VTAIL.n178 9.3005
R1086 VTAIL.n181 VTAIL.n180 9.3005
R1087 VTAIL.n168 VTAIL.n167 9.3005
R1088 VTAIL.n187 VTAIL.n186 9.3005
R1089 VTAIL.n189 VTAIL.n188 9.3005
R1090 VTAIL.n163 VTAIL.n161 9.3005
R1091 VTAIL.n195 VTAIL.n194 9.3005
R1092 VTAIL.n219 VTAIL.n218 9.3005
R1093 VTAIL.n150 VTAIL.n149 9.3005
R1094 VTAIL.n213 VTAIL.n212 9.3005
R1095 VTAIL.n211 VTAIL.n210 9.3005
R1096 VTAIL.n154 VTAIL.n153 9.3005
R1097 VTAIL.n205 VTAIL.n204 9.3005
R1098 VTAIL.n203 VTAIL.n202 9.3005
R1099 VTAIL.n158 VTAIL.n157 9.3005
R1100 VTAIL.n197 VTAIL.n196 9.3005
R1101 VTAIL.n98 VTAIL.n97 9.3005
R1102 VTAIL.n105 VTAIL.n104 9.3005
R1103 VTAIL.n107 VTAIL.n106 9.3005
R1104 VTAIL.n94 VTAIL.n93 9.3005
R1105 VTAIL.n113 VTAIL.n112 9.3005
R1106 VTAIL.n115 VTAIL.n114 9.3005
R1107 VTAIL.n89 VTAIL.n87 9.3005
R1108 VTAIL.n121 VTAIL.n120 9.3005
R1109 VTAIL.n145 VTAIL.n144 9.3005
R1110 VTAIL.n76 VTAIL.n75 9.3005
R1111 VTAIL.n139 VTAIL.n138 9.3005
R1112 VTAIL.n137 VTAIL.n136 9.3005
R1113 VTAIL.n80 VTAIL.n79 9.3005
R1114 VTAIL.n131 VTAIL.n130 9.3005
R1115 VTAIL.n129 VTAIL.n128 9.3005
R1116 VTAIL.n84 VTAIL.n83 9.3005
R1117 VTAIL.n123 VTAIL.n122 9.3005
R1118 VTAIL.n253 VTAIL.n242 8.92171
R1119 VTAIL.n284 VTAIL.n226 8.92171
R1120 VTAIL.n31 VTAIL.n20 8.92171
R1121 VTAIL.n62 VTAIL.n4 8.92171
R1122 VTAIL.n210 VTAIL.n152 8.92171
R1123 VTAIL.n181 VTAIL.n170 8.92171
R1124 VTAIL.n136 VTAIL.n78 8.92171
R1125 VTAIL.n107 VTAIL.n96 8.92171
R1126 VTAIL.n250 VTAIL.n249 8.14595
R1127 VTAIL.n288 VTAIL.n287 8.14595
R1128 VTAIL.n28 VTAIL.n27 8.14595
R1129 VTAIL.n66 VTAIL.n65 8.14595
R1130 VTAIL.n214 VTAIL.n213 8.14595
R1131 VTAIL.n178 VTAIL.n177 8.14595
R1132 VTAIL.n140 VTAIL.n139 8.14595
R1133 VTAIL.n104 VTAIL.n103 8.14595
R1134 VTAIL.n246 VTAIL.n244 7.3702
R1135 VTAIL.n291 VTAIL.n224 7.3702
R1136 VTAIL.n294 VTAIL.n222 7.3702
R1137 VTAIL.n24 VTAIL.n22 7.3702
R1138 VTAIL.n69 VTAIL.n2 7.3702
R1139 VTAIL.n72 VTAIL.n0 7.3702
R1140 VTAIL.n220 VTAIL.n148 7.3702
R1141 VTAIL.n217 VTAIL.n150 7.3702
R1142 VTAIL.n174 VTAIL.n172 7.3702
R1143 VTAIL.n146 VTAIL.n74 7.3702
R1144 VTAIL.n143 VTAIL.n76 7.3702
R1145 VTAIL.n100 VTAIL.n98 7.3702
R1146 VTAIL.n292 VTAIL.n291 6.59444
R1147 VTAIL.n292 VTAIL.n222 6.59444
R1148 VTAIL.n70 VTAIL.n69 6.59444
R1149 VTAIL.n70 VTAIL.n0 6.59444
R1150 VTAIL.n218 VTAIL.n148 6.59444
R1151 VTAIL.n218 VTAIL.n217 6.59444
R1152 VTAIL.n144 VTAIL.n74 6.59444
R1153 VTAIL.n144 VTAIL.n143 6.59444
R1154 VTAIL.n249 VTAIL.n244 5.81868
R1155 VTAIL.n288 VTAIL.n224 5.81868
R1156 VTAIL.n27 VTAIL.n22 5.81868
R1157 VTAIL.n66 VTAIL.n2 5.81868
R1158 VTAIL.n214 VTAIL.n150 5.81868
R1159 VTAIL.n177 VTAIL.n172 5.81868
R1160 VTAIL.n140 VTAIL.n76 5.81868
R1161 VTAIL.n103 VTAIL.n98 5.81868
R1162 VTAIL.n250 VTAIL.n242 5.04292
R1163 VTAIL.n287 VTAIL.n226 5.04292
R1164 VTAIL.n28 VTAIL.n20 5.04292
R1165 VTAIL.n65 VTAIL.n4 5.04292
R1166 VTAIL.n213 VTAIL.n152 5.04292
R1167 VTAIL.n178 VTAIL.n170 5.04292
R1168 VTAIL.n139 VTAIL.n78 5.04292
R1169 VTAIL.n104 VTAIL.n96 5.04292
R1170 VTAIL.n254 VTAIL.n253 4.26717
R1171 VTAIL.n284 VTAIL.n283 4.26717
R1172 VTAIL.n32 VTAIL.n31 4.26717
R1173 VTAIL.n62 VTAIL.n61 4.26717
R1174 VTAIL.n210 VTAIL.n209 4.26717
R1175 VTAIL.n182 VTAIL.n181 4.26717
R1176 VTAIL.n136 VTAIL.n135 4.26717
R1177 VTAIL.n108 VTAIL.n107 4.26717
R1178 VTAIL.n257 VTAIL.n240 3.49141
R1179 VTAIL.n280 VTAIL.n228 3.49141
R1180 VTAIL.n35 VTAIL.n18 3.49141
R1181 VTAIL.n58 VTAIL.n6 3.49141
R1182 VTAIL.n206 VTAIL.n154 3.49141
R1183 VTAIL.n185 VTAIL.n168 3.49141
R1184 VTAIL.n132 VTAIL.n80 3.49141
R1185 VTAIL.n111 VTAIL.n94 3.49141
R1186 VTAIL.n258 VTAIL.n238 2.71565
R1187 VTAIL.n279 VTAIL.n230 2.71565
R1188 VTAIL.n36 VTAIL.n16 2.71565
R1189 VTAIL.n57 VTAIL.n8 2.71565
R1190 VTAIL.n205 VTAIL.n156 2.71565
R1191 VTAIL.n186 VTAIL.n166 2.71565
R1192 VTAIL.n131 VTAIL.n82 2.71565
R1193 VTAIL.n112 VTAIL.n92 2.71565
R1194 VTAIL.n245 VTAIL.n243 2.41282
R1195 VTAIL.n23 VTAIL.n21 2.41282
R1196 VTAIL.n173 VTAIL.n171 2.41282
R1197 VTAIL.n99 VTAIL.n97 2.41282
R1198 VTAIL.n263 VTAIL.n261 1.93989
R1199 VTAIL.n276 VTAIL.n275 1.93989
R1200 VTAIL.n41 VTAIL.n39 1.93989
R1201 VTAIL.n54 VTAIL.n53 1.93989
R1202 VTAIL.n202 VTAIL.n201 1.93989
R1203 VTAIL.n190 VTAIL.n189 1.93989
R1204 VTAIL.n128 VTAIL.n127 1.93989
R1205 VTAIL.n116 VTAIL.n115 1.93989
R1206 VTAIL.n262 VTAIL.n236 1.16414
R1207 VTAIL.n272 VTAIL.n232 1.16414
R1208 VTAIL.n40 VTAIL.n14 1.16414
R1209 VTAIL.n50 VTAIL.n10 1.16414
R1210 VTAIL.n198 VTAIL.n158 1.16414
R1211 VTAIL.n193 VTAIL.n163 1.16414
R1212 VTAIL.n124 VTAIL.n84 1.16414
R1213 VTAIL.n119 VTAIL.n89 1.16414
R1214 VTAIL.n221 VTAIL.n147 1.08671
R1215 VTAIL VTAIL.n73 0.836707
R1216 VTAIL.n268 VTAIL.n267 0.388379
R1217 VTAIL.n271 VTAIL.n234 0.388379
R1218 VTAIL.n46 VTAIL.n45 0.388379
R1219 VTAIL.n49 VTAIL.n12 0.388379
R1220 VTAIL.n197 VTAIL.n160 0.388379
R1221 VTAIL.n194 VTAIL.n162 0.388379
R1222 VTAIL.n123 VTAIL.n86 0.388379
R1223 VTAIL.n120 VTAIL.n88 0.388379
R1224 VTAIL VTAIL.n295 0.2505
R1225 VTAIL.n251 VTAIL.n243 0.155672
R1226 VTAIL.n252 VTAIL.n251 0.155672
R1227 VTAIL.n252 VTAIL.n239 0.155672
R1228 VTAIL.n259 VTAIL.n239 0.155672
R1229 VTAIL.n260 VTAIL.n259 0.155672
R1230 VTAIL.n260 VTAIL.n235 0.155672
R1231 VTAIL.n269 VTAIL.n235 0.155672
R1232 VTAIL.n270 VTAIL.n269 0.155672
R1233 VTAIL.n270 VTAIL.n231 0.155672
R1234 VTAIL.n277 VTAIL.n231 0.155672
R1235 VTAIL.n278 VTAIL.n277 0.155672
R1236 VTAIL.n278 VTAIL.n227 0.155672
R1237 VTAIL.n285 VTAIL.n227 0.155672
R1238 VTAIL.n286 VTAIL.n285 0.155672
R1239 VTAIL.n286 VTAIL.n223 0.155672
R1240 VTAIL.n293 VTAIL.n223 0.155672
R1241 VTAIL.n29 VTAIL.n21 0.155672
R1242 VTAIL.n30 VTAIL.n29 0.155672
R1243 VTAIL.n30 VTAIL.n17 0.155672
R1244 VTAIL.n37 VTAIL.n17 0.155672
R1245 VTAIL.n38 VTAIL.n37 0.155672
R1246 VTAIL.n38 VTAIL.n13 0.155672
R1247 VTAIL.n47 VTAIL.n13 0.155672
R1248 VTAIL.n48 VTAIL.n47 0.155672
R1249 VTAIL.n48 VTAIL.n9 0.155672
R1250 VTAIL.n55 VTAIL.n9 0.155672
R1251 VTAIL.n56 VTAIL.n55 0.155672
R1252 VTAIL.n56 VTAIL.n5 0.155672
R1253 VTAIL.n63 VTAIL.n5 0.155672
R1254 VTAIL.n64 VTAIL.n63 0.155672
R1255 VTAIL.n64 VTAIL.n1 0.155672
R1256 VTAIL.n71 VTAIL.n1 0.155672
R1257 VTAIL.n219 VTAIL.n149 0.155672
R1258 VTAIL.n212 VTAIL.n149 0.155672
R1259 VTAIL.n212 VTAIL.n211 0.155672
R1260 VTAIL.n211 VTAIL.n153 0.155672
R1261 VTAIL.n204 VTAIL.n153 0.155672
R1262 VTAIL.n204 VTAIL.n203 0.155672
R1263 VTAIL.n203 VTAIL.n157 0.155672
R1264 VTAIL.n196 VTAIL.n157 0.155672
R1265 VTAIL.n196 VTAIL.n195 0.155672
R1266 VTAIL.n195 VTAIL.n161 0.155672
R1267 VTAIL.n188 VTAIL.n161 0.155672
R1268 VTAIL.n188 VTAIL.n187 0.155672
R1269 VTAIL.n187 VTAIL.n167 0.155672
R1270 VTAIL.n180 VTAIL.n167 0.155672
R1271 VTAIL.n180 VTAIL.n179 0.155672
R1272 VTAIL.n179 VTAIL.n171 0.155672
R1273 VTAIL.n145 VTAIL.n75 0.155672
R1274 VTAIL.n138 VTAIL.n75 0.155672
R1275 VTAIL.n138 VTAIL.n137 0.155672
R1276 VTAIL.n137 VTAIL.n79 0.155672
R1277 VTAIL.n130 VTAIL.n79 0.155672
R1278 VTAIL.n130 VTAIL.n129 0.155672
R1279 VTAIL.n129 VTAIL.n83 0.155672
R1280 VTAIL.n122 VTAIL.n83 0.155672
R1281 VTAIL.n122 VTAIL.n121 0.155672
R1282 VTAIL.n121 VTAIL.n87 0.155672
R1283 VTAIL.n114 VTAIL.n87 0.155672
R1284 VTAIL.n114 VTAIL.n113 0.155672
R1285 VTAIL.n113 VTAIL.n93 0.155672
R1286 VTAIL.n106 VTAIL.n93 0.155672
R1287 VTAIL.n106 VTAIL.n105 0.155672
R1288 VTAIL.n105 VTAIL.n97 0.155672
R1289 VDD2.n141 VDD2.n73 756.745
R1290 VDD2.n68 VDD2.n0 756.745
R1291 VDD2.n142 VDD2.n141 585
R1292 VDD2.n140 VDD2.n139 585
R1293 VDD2.n77 VDD2.n76 585
R1294 VDD2.n134 VDD2.n133 585
R1295 VDD2.n132 VDD2.n131 585
R1296 VDD2.n81 VDD2.n80 585
R1297 VDD2.n126 VDD2.n125 585
R1298 VDD2.n124 VDD2.n123 585
R1299 VDD2.n85 VDD2.n84 585
R1300 VDD2.n89 VDD2.n87 585
R1301 VDD2.n118 VDD2.n117 585
R1302 VDD2.n116 VDD2.n115 585
R1303 VDD2.n91 VDD2.n90 585
R1304 VDD2.n110 VDD2.n109 585
R1305 VDD2.n108 VDD2.n107 585
R1306 VDD2.n95 VDD2.n94 585
R1307 VDD2.n102 VDD2.n101 585
R1308 VDD2.n100 VDD2.n99 585
R1309 VDD2.n25 VDD2.n24 585
R1310 VDD2.n27 VDD2.n26 585
R1311 VDD2.n20 VDD2.n19 585
R1312 VDD2.n33 VDD2.n32 585
R1313 VDD2.n35 VDD2.n34 585
R1314 VDD2.n16 VDD2.n15 585
R1315 VDD2.n42 VDD2.n41 585
R1316 VDD2.n43 VDD2.n14 585
R1317 VDD2.n45 VDD2.n44 585
R1318 VDD2.n12 VDD2.n11 585
R1319 VDD2.n51 VDD2.n50 585
R1320 VDD2.n53 VDD2.n52 585
R1321 VDD2.n8 VDD2.n7 585
R1322 VDD2.n59 VDD2.n58 585
R1323 VDD2.n61 VDD2.n60 585
R1324 VDD2.n4 VDD2.n3 585
R1325 VDD2.n67 VDD2.n66 585
R1326 VDD2.n69 VDD2.n68 585
R1327 VDD2.n98 VDD2.t0 329.036
R1328 VDD2.n23 VDD2.t1 329.036
R1329 VDD2.n141 VDD2.n140 171.744
R1330 VDD2.n140 VDD2.n76 171.744
R1331 VDD2.n133 VDD2.n76 171.744
R1332 VDD2.n133 VDD2.n132 171.744
R1333 VDD2.n132 VDD2.n80 171.744
R1334 VDD2.n125 VDD2.n80 171.744
R1335 VDD2.n125 VDD2.n124 171.744
R1336 VDD2.n124 VDD2.n84 171.744
R1337 VDD2.n89 VDD2.n84 171.744
R1338 VDD2.n117 VDD2.n89 171.744
R1339 VDD2.n117 VDD2.n116 171.744
R1340 VDD2.n116 VDD2.n90 171.744
R1341 VDD2.n109 VDD2.n90 171.744
R1342 VDD2.n109 VDD2.n108 171.744
R1343 VDD2.n108 VDD2.n94 171.744
R1344 VDD2.n101 VDD2.n94 171.744
R1345 VDD2.n101 VDD2.n100 171.744
R1346 VDD2.n26 VDD2.n25 171.744
R1347 VDD2.n26 VDD2.n19 171.744
R1348 VDD2.n33 VDD2.n19 171.744
R1349 VDD2.n34 VDD2.n33 171.744
R1350 VDD2.n34 VDD2.n15 171.744
R1351 VDD2.n42 VDD2.n15 171.744
R1352 VDD2.n43 VDD2.n42 171.744
R1353 VDD2.n44 VDD2.n43 171.744
R1354 VDD2.n44 VDD2.n11 171.744
R1355 VDD2.n51 VDD2.n11 171.744
R1356 VDD2.n52 VDD2.n51 171.744
R1357 VDD2.n52 VDD2.n7 171.744
R1358 VDD2.n59 VDD2.n7 171.744
R1359 VDD2.n60 VDD2.n59 171.744
R1360 VDD2.n60 VDD2.n3 171.744
R1361 VDD2.n67 VDD2.n3 171.744
R1362 VDD2.n68 VDD2.n67 171.744
R1363 VDD2.n146 VDD2.n72 85.8858
R1364 VDD2.n100 VDD2.t0 85.8723
R1365 VDD2.n25 VDD2.t1 85.8723
R1366 VDD2.n146 VDD2.n145 48.0884
R1367 VDD2.n87 VDD2.n85 13.1884
R1368 VDD2.n45 VDD2.n12 13.1884
R1369 VDD2.n123 VDD2.n122 12.8005
R1370 VDD2.n119 VDD2.n118 12.8005
R1371 VDD2.n46 VDD2.n14 12.8005
R1372 VDD2.n50 VDD2.n49 12.8005
R1373 VDD2.n126 VDD2.n83 12.0247
R1374 VDD2.n115 VDD2.n88 12.0247
R1375 VDD2.n41 VDD2.n40 12.0247
R1376 VDD2.n53 VDD2.n10 12.0247
R1377 VDD2.n127 VDD2.n81 11.249
R1378 VDD2.n114 VDD2.n91 11.249
R1379 VDD2.n39 VDD2.n16 11.249
R1380 VDD2.n54 VDD2.n8 11.249
R1381 VDD2.n99 VDD2.n98 10.7239
R1382 VDD2.n24 VDD2.n23 10.7239
R1383 VDD2.n131 VDD2.n130 10.4732
R1384 VDD2.n111 VDD2.n110 10.4732
R1385 VDD2.n36 VDD2.n35 10.4732
R1386 VDD2.n58 VDD2.n57 10.4732
R1387 VDD2.n134 VDD2.n79 9.69747
R1388 VDD2.n107 VDD2.n93 9.69747
R1389 VDD2.n32 VDD2.n18 9.69747
R1390 VDD2.n61 VDD2.n6 9.69747
R1391 VDD2.n145 VDD2.n144 9.45567
R1392 VDD2.n72 VDD2.n71 9.45567
R1393 VDD2.n97 VDD2.n96 9.3005
R1394 VDD2.n104 VDD2.n103 9.3005
R1395 VDD2.n106 VDD2.n105 9.3005
R1396 VDD2.n93 VDD2.n92 9.3005
R1397 VDD2.n112 VDD2.n111 9.3005
R1398 VDD2.n114 VDD2.n113 9.3005
R1399 VDD2.n88 VDD2.n86 9.3005
R1400 VDD2.n120 VDD2.n119 9.3005
R1401 VDD2.n144 VDD2.n143 9.3005
R1402 VDD2.n75 VDD2.n74 9.3005
R1403 VDD2.n138 VDD2.n137 9.3005
R1404 VDD2.n136 VDD2.n135 9.3005
R1405 VDD2.n79 VDD2.n78 9.3005
R1406 VDD2.n130 VDD2.n129 9.3005
R1407 VDD2.n128 VDD2.n127 9.3005
R1408 VDD2.n83 VDD2.n82 9.3005
R1409 VDD2.n122 VDD2.n121 9.3005
R1410 VDD2.n71 VDD2.n70 9.3005
R1411 VDD2.n65 VDD2.n64 9.3005
R1412 VDD2.n63 VDD2.n62 9.3005
R1413 VDD2.n6 VDD2.n5 9.3005
R1414 VDD2.n57 VDD2.n56 9.3005
R1415 VDD2.n55 VDD2.n54 9.3005
R1416 VDD2.n10 VDD2.n9 9.3005
R1417 VDD2.n49 VDD2.n48 9.3005
R1418 VDD2.n22 VDD2.n21 9.3005
R1419 VDD2.n29 VDD2.n28 9.3005
R1420 VDD2.n31 VDD2.n30 9.3005
R1421 VDD2.n18 VDD2.n17 9.3005
R1422 VDD2.n37 VDD2.n36 9.3005
R1423 VDD2.n39 VDD2.n38 9.3005
R1424 VDD2.n40 VDD2.n13 9.3005
R1425 VDD2.n47 VDD2.n46 9.3005
R1426 VDD2.n2 VDD2.n1 9.3005
R1427 VDD2.n135 VDD2.n77 8.92171
R1428 VDD2.n106 VDD2.n95 8.92171
R1429 VDD2.n31 VDD2.n20 8.92171
R1430 VDD2.n62 VDD2.n4 8.92171
R1431 VDD2.n139 VDD2.n138 8.14595
R1432 VDD2.n103 VDD2.n102 8.14595
R1433 VDD2.n28 VDD2.n27 8.14595
R1434 VDD2.n66 VDD2.n65 8.14595
R1435 VDD2.n145 VDD2.n73 7.3702
R1436 VDD2.n142 VDD2.n75 7.3702
R1437 VDD2.n99 VDD2.n97 7.3702
R1438 VDD2.n24 VDD2.n22 7.3702
R1439 VDD2.n69 VDD2.n2 7.3702
R1440 VDD2.n72 VDD2.n0 7.3702
R1441 VDD2.n143 VDD2.n73 6.59444
R1442 VDD2.n143 VDD2.n142 6.59444
R1443 VDD2.n70 VDD2.n69 6.59444
R1444 VDD2.n70 VDD2.n0 6.59444
R1445 VDD2.n139 VDD2.n75 5.81868
R1446 VDD2.n102 VDD2.n97 5.81868
R1447 VDD2.n27 VDD2.n22 5.81868
R1448 VDD2.n66 VDD2.n2 5.81868
R1449 VDD2.n138 VDD2.n77 5.04292
R1450 VDD2.n103 VDD2.n95 5.04292
R1451 VDD2.n28 VDD2.n20 5.04292
R1452 VDD2.n65 VDD2.n4 5.04292
R1453 VDD2.n135 VDD2.n134 4.26717
R1454 VDD2.n107 VDD2.n106 4.26717
R1455 VDD2.n32 VDD2.n31 4.26717
R1456 VDD2.n62 VDD2.n61 4.26717
R1457 VDD2.n131 VDD2.n79 3.49141
R1458 VDD2.n110 VDD2.n93 3.49141
R1459 VDD2.n35 VDD2.n18 3.49141
R1460 VDD2.n58 VDD2.n6 3.49141
R1461 VDD2.n130 VDD2.n81 2.71565
R1462 VDD2.n111 VDD2.n91 2.71565
R1463 VDD2.n36 VDD2.n16 2.71565
R1464 VDD2.n57 VDD2.n8 2.71565
R1465 VDD2.n98 VDD2.n96 2.41282
R1466 VDD2.n23 VDD2.n21 2.41282
R1467 VDD2.n127 VDD2.n126 1.93989
R1468 VDD2.n115 VDD2.n114 1.93989
R1469 VDD2.n41 VDD2.n39 1.93989
R1470 VDD2.n54 VDD2.n53 1.93989
R1471 VDD2.n123 VDD2.n83 1.16414
R1472 VDD2.n118 VDD2.n88 1.16414
R1473 VDD2.n40 VDD2.n14 1.16414
R1474 VDD2.n50 VDD2.n10 1.16414
R1475 VDD2.n122 VDD2.n85 0.388379
R1476 VDD2.n119 VDD2.n87 0.388379
R1477 VDD2.n46 VDD2.n45 0.388379
R1478 VDD2.n49 VDD2.n12 0.388379
R1479 VDD2 VDD2.n146 0.366879
R1480 VDD2.n144 VDD2.n74 0.155672
R1481 VDD2.n137 VDD2.n74 0.155672
R1482 VDD2.n137 VDD2.n136 0.155672
R1483 VDD2.n136 VDD2.n78 0.155672
R1484 VDD2.n129 VDD2.n78 0.155672
R1485 VDD2.n129 VDD2.n128 0.155672
R1486 VDD2.n128 VDD2.n82 0.155672
R1487 VDD2.n121 VDD2.n82 0.155672
R1488 VDD2.n121 VDD2.n120 0.155672
R1489 VDD2.n120 VDD2.n86 0.155672
R1490 VDD2.n113 VDD2.n86 0.155672
R1491 VDD2.n113 VDD2.n112 0.155672
R1492 VDD2.n112 VDD2.n92 0.155672
R1493 VDD2.n105 VDD2.n92 0.155672
R1494 VDD2.n105 VDD2.n104 0.155672
R1495 VDD2.n104 VDD2.n96 0.155672
R1496 VDD2.n29 VDD2.n21 0.155672
R1497 VDD2.n30 VDD2.n29 0.155672
R1498 VDD2.n30 VDD2.n17 0.155672
R1499 VDD2.n37 VDD2.n17 0.155672
R1500 VDD2.n38 VDD2.n37 0.155672
R1501 VDD2.n38 VDD2.n13 0.155672
R1502 VDD2.n47 VDD2.n13 0.155672
R1503 VDD2.n48 VDD2.n47 0.155672
R1504 VDD2.n48 VDD2.n9 0.155672
R1505 VDD2.n55 VDD2.n9 0.155672
R1506 VDD2.n56 VDD2.n55 0.155672
R1507 VDD2.n56 VDD2.n5 0.155672
R1508 VDD2.n63 VDD2.n5 0.155672
R1509 VDD2.n64 VDD2.n63 0.155672
R1510 VDD2.n64 VDD2.n1 0.155672
R1511 VDD2.n71 VDD2.n1 0.155672
R1512 VP.n0 VP.t1 535.067
R1513 VP.n0 VP.t0 493.224
R1514 VP VP.n0 0.0516364
R1515 VDD1.n68 VDD1.n0 756.745
R1516 VDD1.n141 VDD1.n73 756.745
R1517 VDD1.n69 VDD1.n68 585
R1518 VDD1.n67 VDD1.n66 585
R1519 VDD1.n4 VDD1.n3 585
R1520 VDD1.n61 VDD1.n60 585
R1521 VDD1.n59 VDD1.n58 585
R1522 VDD1.n8 VDD1.n7 585
R1523 VDD1.n53 VDD1.n52 585
R1524 VDD1.n51 VDD1.n50 585
R1525 VDD1.n12 VDD1.n11 585
R1526 VDD1.n16 VDD1.n14 585
R1527 VDD1.n45 VDD1.n44 585
R1528 VDD1.n43 VDD1.n42 585
R1529 VDD1.n18 VDD1.n17 585
R1530 VDD1.n37 VDD1.n36 585
R1531 VDD1.n35 VDD1.n34 585
R1532 VDD1.n22 VDD1.n21 585
R1533 VDD1.n29 VDD1.n28 585
R1534 VDD1.n27 VDD1.n26 585
R1535 VDD1.n98 VDD1.n97 585
R1536 VDD1.n100 VDD1.n99 585
R1537 VDD1.n93 VDD1.n92 585
R1538 VDD1.n106 VDD1.n105 585
R1539 VDD1.n108 VDD1.n107 585
R1540 VDD1.n89 VDD1.n88 585
R1541 VDD1.n115 VDD1.n114 585
R1542 VDD1.n116 VDD1.n87 585
R1543 VDD1.n118 VDD1.n117 585
R1544 VDD1.n85 VDD1.n84 585
R1545 VDD1.n124 VDD1.n123 585
R1546 VDD1.n126 VDD1.n125 585
R1547 VDD1.n81 VDD1.n80 585
R1548 VDD1.n132 VDD1.n131 585
R1549 VDD1.n134 VDD1.n133 585
R1550 VDD1.n77 VDD1.n76 585
R1551 VDD1.n140 VDD1.n139 585
R1552 VDD1.n142 VDD1.n141 585
R1553 VDD1.n25 VDD1.t0 329.036
R1554 VDD1.n96 VDD1.t1 329.036
R1555 VDD1.n68 VDD1.n67 171.744
R1556 VDD1.n67 VDD1.n3 171.744
R1557 VDD1.n60 VDD1.n3 171.744
R1558 VDD1.n60 VDD1.n59 171.744
R1559 VDD1.n59 VDD1.n7 171.744
R1560 VDD1.n52 VDD1.n7 171.744
R1561 VDD1.n52 VDD1.n51 171.744
R1562 VDD1.n51 VDD1.n11 171.744
R1563 VDD1.n16 VDD1.n11 171.744
R1564 VDD1.n44 VDD1.n16 171.744
R1565 VDD1.n44 VDD1.n43 171.744
R1566 VDD1.n43 VDD1.n17 171.744
R1567 VDD1.n36 VDD1.n17 171.744
R1568 VDD1.n36 VDD1.n35 171.744
R1569 VDD1.n35 VDD1.n21 171.744
R1570 VDD1.n28 VDD1.n21 171.744
R1571 VDD1.n28 VDD1.n27 171.744
R1572 VDD1.n99 VDD1.n98 171.744
R1573 VDD1.n99 VDD1.n92 171.744
R1574 VDD1.n106 VDD1.n92 171.744
R1575 VDD1.n107 VDD1.n106 171.744
R1576 VDD1.n107 VDD1.n88 171.744
R1577 VDD1.n115 VDD1.n88 171.744
R1578 VDD1.n116 VDD1.n115 171.744
R1579 VDD1.n117 VDD1.n116 171.744
R1580 VDD1.n117 VDD1.n84 171.744
R1581 VDD1.n124 VDD1.n84 171.744
R1582 VDD1.n125 VDD1.n124 171.744
R1583 VDD1.n125 VDD1.n80 171.744
R1584 VDD1.n132 VDD1.n80 171.744
R1585 VDD1.n133 VDD1.n132 171.744
R1586 VDD1.n133 VDD1.n76 171.744
R1587 VDD1.n140 VDD1.n76 171.744
R1588 VDD1.n141 VDD1.n140 171.744
R1589 VDD1 VDD1.n145 86.7188
R1590 VDD1.n27 VDD1.t0 85.8723
R1591 VDD1.n98 VDD1.t1 85.8723
R1592 VDD1 VDD1.n72 48.4548
R1593 VDD1.n14 VDD1.n12 13.1884
R1594 VDD1.n118 VDD1.n85 13.1884
R1595 VDD1.n50 VDD1.n49 12.8005
R1596 VDD1.n46 VDD1.n45 12.8005
R1597 VDD1.n119 VDD1.n87 12.8005
R1598 VDD1.n123 VDD1.n122 12.8005
R1599 VDD1.n53 VDD1.n10 12.0247
R1600 VDD1.n42 VDD1.n15 12.0247
R1601 VDD1.n114 VDD1.n113 12.0247
R1602 VDD1.n126 VDD1.n83 12.0247
R1603 VDD1.n54 VDD1.n8 11.249
R1604 VDD1.n41 VDD1.n18 11.249
R1605 VDD1.n112 VDD1.n89 11.249
R1606 VDD1.n127 VDD1.n81 11.249
R1607 VDD1.n26 VDD1.n25 10.7239
R1608 VDD1.n97 VDD1.n96 10.7239
R1609 VDD1.n58 VDD1.n57 10.4732
R1610 VDD1.n38 VDD1.n37 10.4732
R1611 VDD1.n109 VDD1.n108 10.4732
R1612 VDD1.n131 VDD1.n130 10.4732
R1613 VDD1.n61 VDD1.n6 9.69747
R1614 VDD1.n34 VDD1.n20 9.69747
R1615 VDD1.n105 VDD1.n91 9.69747
R1616 VDD1.n134 VDD1.n79 9.69747
R1617 VDD1.n72 VDD1.n71 9.45567
R1618 VDD1.n145 VDD1.n144 9.45567
R1619 VDD1.n24 VDD1.n23 9.3005
R1620 VDD1.n31 VDD1.n30 9.3005
R1621 VDD1.n33 VDD1.n32 9.3005
R1622 VDD1.n20 VDD1.n19 9.3005
R1623 VDD1.n39 VDD1.n38 9.3005
R1624 VDD1.n41 VDD1.n40 9.3005
R1625 VDD1.n15 VDD1.n13 9.3005
R1626 VDD1.n47 VDD1.n46 9.3005
R1627 VDD1.n71 VDD1.n70 9.3005
R1628 VDD1.n2 VDD1.n1 9.3005
R1629 VDD1.n65 VDD1.n64 9.3005
R1630 VDD1.n63 VDD1.n62 9.3005
R1631 VDD1.n6 VDD1.n5 9.3005
R1632 VDD1.n57 VDD1.n56 9.3005
R1633 VDD1.n55 VDD1.n54 9.3005
R1634 VDD1.n10 VDD1.n9 9.3005
R1635 VDD1.n49 VDD1.n48 9.3005
R1636 VDD1.n144 VDD1.n143 9.3005
R1637 VDD1.n138 VDD1.n137 9.3005
R1638 VDD1.n136 VDD1.n135 9.3005
R1639 VDD1.n79 VDD1.n78 9.3005
R1640 VDD1.n130 VDD1.n129 9.3005
R1641 VDD1.n128 VDD1.n127 9.3005
R1642 VDD1.n83 VDD1.n82 9.3005
R1643 VDD1.n122 VDD1.n121 9.3005
R1644 VDD1.n95 VDD1.n94 9.3005
R1645 VDD1.n102 VDD1.n101 9.3005
R1646 VDD1.n104 VDD1.n103 9.3005
R1647 VDD1.n91 VDD1.n90 9.3005
R1648 VDD1.n110 VDD1.n109 9.3005
R1649 VDD1.n112 VDD1.n111 9.3005
R1650 VDD1.n113 VDD1.n86 9.3005
R1651 VDD1.n120 VDD1.n119 9.3005
R1652 VDD1.n75 VDD1.n74 9.3005
R1653 VDD1.n62 VDD1.n4 8.92171
R1654 VDD1.n33 VDD1.n22 8.92171
R1655 VDD1.n104 VDD1.n93 8.92171
R1656 VDD1.n135 VDD1.n77 8.92171
R1657 VDD1.n66 VDD1.n65 8.14595
R1658 VDD1.n30 VDD1.n29 8.14595
R1659 VDD1.n101 VDD1.n100 8.14595
R1660 VDD1.n139 VDD1.n138 8.14595
R1661 VDD1.n72 VDD1.n0 7.3702
R1662 VDD1.n69 VDD1.n2 7.3702
R1663 VDD1.n26 VDD1.n24 7.3702
R1664 VDD1.n97 VDD1.n95 7.3702
R1665 VDD1.n142 VDD1.n75 7.3702
R1666 VDD1.n145 VDD1.n73 7.3702
R1667 VDD1.n70 VDD1.n0 6.59444
R1668 VDD1.n70 VDD1.n69 6.59444
R1669 VDD1.n143 VDD1.n142 6.59444
R1670 VDD1.n143 VDD1.n73 6.59444
R1671 VDD1.n66 VDD1.n2 5.81868
R1672 VDD1.n29 VDD1.n24 5.81868
R1673 VDD1.n100 VDD1.n95 5.81868
R1674 VDD1.n139 VDD1.n75 5.81868
R1675 VDD1.n65 VDD1.n4 5.04292
R1676 VDD1.n30 VDD1.n22 5.04292
R1677 VDD1.n101 VDD1.n93 5.04292
R1678 VDD1.n138 VDD1.n77 5.04292
R1679 VDD1.n62 VDD1.n61 4.26717
R1680 VDD1.n34 VDD1.n33 4.26717
R1681 VDD1.n105 VDD1.n104 4.26717
R1682 VDD1.n135 VDD1.n134 4.26717
R1683 VDD1.n58 VDD1.n6 3.49141
R1684 VDD1.n37 VDD1.n20 3.49141
R1685 VDD1.n108 VDD1.n91 3.49141
R1686 VDD1.n131 VDD1.n79 3.49141
R1687 VDD1.n57 VDD1.n8 2.71565
R1688 VDD1.n38 VDD1.n18 2.71565
R1689 VDD1.n109 VDD1.n89 2.71565
R1690 VDD1.n130 VDD1.n81 2.71565
R1691 VDD1.n25 VDD1.n23 2.41282
R1692 VDD1.n96 VDD1.n94 2.41282
R1693 VDD1.n54 VDD1.n53 1.93989
R1694 VDD1.n42 VDD1.n41 1.93989
R1695 VDD1.n114 VDD1.n112 1.93989
R1696 VDD1.n127 VDD1.n126 1.93989
R1697 VDD1.n50 VDD1.n10 1.16414
R1698 VDD1.n45 VDD1.n15 1.16414
R1699 VDD1.n113 VDD1.n87 1.16414
R1700 VDD1.n123 VDD1.n83 1.16414
R1701 VDD1.n49 VDD1.n12 0.388379
R1702 VDD1.n46 VDD1.n14 0.388379
R1703 VDD1.n119 VDD1.n118 0.388379
R1704 VDD1.n122 VDD1.n85 0.388379
R1705 VDD1.n71 VDD1.n1 0.155672
R1706 VDD1.n64 VDD1.n1 0.155672
R1707 VDD1.n64 VDD1.n63 0.155672
R1708 VDD1.n63 VDD1.n5 0.155672
R1709 VDD1.n56 VDD1.n5 0.155672
R1710 VDD1.n56 VDD1.n55 0.155672
R1711 VDD1.n55 VDD1.n9 0.155672
R1712 VDD1.n48 VDD1.n9 0.155672
R1713 VDD1.n48 VDD1.n47 0.155672
R1714 VDD1.n47 VDD1.n13 0.155672
R1715 VDD1.n40 VDD1.n13 0.155672
R1716 VDD1.n40 VDD1.n39 0.155672
R1717 VDD1.n39 VDD1.n19 0.155672
R1718 VDD1.n32 VDD1.n19 0.155672
R1719 VDD1.n32 VDD1.n31 0.155672
R1720 VDD1.n31 VDD1.n23 0.155672
R1721 VDD1.n102 VDD1.n94 0.155672
R1722 VDD1.n103 VDD1.n102 0.155672
R1723 VDD1.n103 VDD1.n90 0.155672
R1724 VDD1.n110 VDD1.n90 0.155672
R1725 VDD1.n111 VDD1.n110 0.155672
R1726 VDD1.n111 VDD1.n86 0.155672
R1727 VDD1.n120 VDD1.n86 0.155672
R1728 VDD1.n121 VDD1.n120 0.155672
R1729 VDD1.n121 VDD1.n82 0.155672
R1730 VDD1.n128 VDD1.n82 0.155672
R1731 VDD1.n129 VDD1.n128 0.155672
R1732 VDD1.n129 VDD1.n78 0.155672
R1733 VDD1.n136 VDD1.n78 0.155672
R1734 VDD1.n137 VDD1.n136 0.155672
R1735 VDD1.n137 VDD1.n74 0.155672
R1736 VDD1.n144 VDD1.n74 0.155672
C0 VTAIL w_n1542_n3676# 3.09788f
C1 VN VDD2 2.56197f
C2 VDD2 VP 0.272168f
C3 VDD1 w_n1542_n3676# 1.72503f
C4 VN B 0.816494f
C5 VP B 1.12808f
C6 VDD1 VTAIL 5.71987f
C7 w_n1542_n3676# VDD2 1.73371f
C8 VTAIL VDD2 5.75707f
C9 w_n1542_n3676# B 7.6192f
C10 VTAIL B 3.22819f
C11 VDD1 VDD2 0.502912f
C12 VDD1 B 1.59854f
C13 VN VP 5.02158f
C14 VDD2 B 1.61592f
C15 VN w_n1542_n3676# 2.0164f
C16 w_n1542_n3676# VP 2.20958f
C17 VTAIL VN 2.04736f
C18 VTAIL VP 2.06191f
C19 VDD1 VN 0.149104f
C20 VDD1 VP 2.68082f
C21 VDD2 VSUBS 0.825942f
C22 VDD1 VSUBS 3.410294f
C23 VTAIL VSUBS 0.876028f
C24 VN VSUBS 7.75289f
C25 VP VSUBS 1.287219f
C26 B VSUBS 2.91795f
C27 w_n1542_n3676# VSUBS 69.6305f
C28 VDD1.n0 VSUBS 0.022622f
C29 VDD1.n1 VSUBS 0.020352f
C30 VDD1.n2 VSUBS 0.010936f
C31 VDD1.n3 VSUBS 0.025849f
C32 VDD1.n4 VSUBS 0.011579f
C33 VDD1.n5 VSUBS 0.020352f
C34 VDD1.n6 VSUBS 0.010936f
C35 VDD1.n7 VSUBS 0.025849f
C36 VDD1.n8 VSUBS 0.011579f
C37 VDD1.n9 VSUBS 0.020352f
C38 VDD1.n10 VSUBS 0.010936f
C39 VDD1.n11 VSUBS 0.025849f
C40 VDD1.n12 VSUBS 0.011258f
C41 VDD1.n13 VSUBS 0.020352f
C42 VDD1.n14 VSUBS 0.011258f
C43 VDD1.n15 VSUBS 0.010936f
C44 VDD1.n16 VSUBS 0.025849f
C45 VDD1.n17 VSUBS 0.025849f
C46 VDD1.n18 VSUBS 0.011579f
C47 VDD1.n19 VSUBS 0.020352f
C48 VDD1.n20 VSUBS 0.010936f
C49 VDD1.n21 VSUBS 0.025849f
C50 VDD1.n22 VSUBS 0.011579f
C51 VDD1.n23 VSUBS 1.13549f
C52 VDD1.n24 VSUBS 0.010936f
C53 VDD1.t0 VSUBS 0.055804f
C54 VDD1.n25 VSUBS 0.174267f
C55 VDD1.n26 VSUBS 0.019445f
C56 VDD1.n27 VSUBS 0.019387f
C57 VDD1.n28 VSUBS 0.025849f
C58 VDD1.n29 VSUBS 0.011579f
C59 VDD1.n30 VSUBS 0.010936f
C60 VDD1.n31 VSUBS 0.020352f
C61 VDD1.n32 VSUBS 0.020352f
C62 VDD1.n33 VSUBS 0.010936f
C63 VDD1.n34 VSUBS 0.011579f
C64 VDD1.n35 VSUBS 0.025849f
C65 VDD1.n36 VSUBS 0.025849f
C66 VDD1.n37 VSUBS 0.011579f
C67 VDD1.n38 VSUBS 0.010936f
C68 VDD1.n39 VSUBS 0.020352f
C69 VDD1.n40 VSUBS 0.020352f
C70 VDD1.n41 VSUBS 0.010936f
C71 VDD1.n42 VSUBS 0.011579f
C72 VDD1.n43 VSUBS 0.025849f
C73 VDD1.n44 VSUBS 0.025849f
C74 VDD1.n45 VSUBS 0.011579f
C75 VDD1.n46 VSUBS 0.010936f
C76 VDD1.n47 VSUBS 0.020352f
C77 VDD1.n48 VSUBS 0.020352f
C78 VDD1.n49 VSUBS 0.010936f
C79 VDD1.n50 VSUBS 0.011579f
C80 VDD1.n51 VSUBS 0.025849f
C81 VDD1.n52 VSUBS 0.025849f
C82 VDD1.n53 VSUBS 0.011579f
C83 VDD1.n54 VSUBS 0.010936f
C84 VDD1.n55 VSUBS 0.020352f
C85 VDD1.n56 VSUBS 0.020352f
C86 VDD1.n57 VSUBS 0.010936f
C87 VDD1.n58 VSUBS 0.011579f
C88 VDD1.n59 VSUBS 0.025849f
C89 VDD1.n60 VSUBS 0.025849f
C90 VDD1.n61 VSUBS 0.011579f
C91 VDD1.n62 VSUBS 0.010936f
C92 VDD1.n63 VSUBS 0.020352f
C93 VDD1.n64 VSUBS 0.020352f
C94 VDD1.n65 VSUBS 0.010936f
C95 VDD1.n66 VSUBS 0.011579f
C96 VDD1.n67 VSUBS 0.025849f
C97 VDD1.n68 VSUBS 0.063463f
C98 VDD1.n69 VSUBS 0.011579f
C99 VDD1.n70 VSUBS 0.010936f
C100 VDD1.n71 VSUBS 0.04593f
C101 VDD1.n72 VSUBS 0.046455f
C102 VDD1.n73 VSUBS 0.022622f
C103 VDD1.n74 VSUBS 0.020352f
C104 VDD1.n75 VSUBS 0.010936f
C105 VDD1.n76 VSUBS 0.025849f
C106 VDD1.n77 VSUBS 0.011579f
C107 VDD1.n78 VSUBS 0.020352f
C108 VDD1.n79 VSUBS 0.010936f
C109 VDD1.n80 VSUBS 0.025849f
C110 VDD1.n81 VSUBS 0.011579f
C111 VDD1.n82 VSUBS 0.020352f
C112 VDD1.n83 VSUBS 0.010936f
C113 VDD1.n84 VSUBS 0.025849f
C114 VDD1.n85 VSUBS 0.011258f
C115 VDD1.n86 VSUBS 0.020352f
C116 VDD1.n87 VSUBS 0.011579f
C117 VDD1.n88 VSUBS 0.025849f
C118 VDD1.n89 VSUBS 0.011579f
C119 VDD1.n90 VSUBS 0.020352f
C120 VDD1.n91 VSUBS 0.010936f
C121 VDD1.n92 VSUBS 0.025849f
C122 VDD1.n93 VSUBS 0.011579f
C123 VDD1.n94 VSUBS 1.13549f
C124 VDD1.n95 VSUBS 0.010936f
C125 VDD1.t1 VSUBS 0.055804f
C126 VDD1.n96 VSUBS 0.174267f
C127 VDD1.n97 VSUBS 0.019445f
C128 VDD1.n98 VSUBS 0.019387f
C129 VDD1.n99 VSUBS 0.025849f
C130 VDD1.n100 VSUBS 0.011579f
C131 VDD1.n101 VSUBS 0.010936f
C132 VDD1.n102 VSUBS 0.020352f
C133 VDD1.n103 VSUBS 0.020352f
C134 VDD1.n104 VSUBS 0.010936f
C135 VDD1.n105 VSUBS 0.011579f
C136 VDD1.n106 VSUBS 0.025849f
C137 VDD1.n107 VSUBS 0.025849f
C138 VDD1.n108 VSUBS 0.011579f
C139 VDD1.n109 VSUBS 0.010936f
C140 VDD1.n110 VSUBS 0.020352f
C141 VDD1.n111 VSUBS 0.020352f
C142 VDD1.n112 VSUBS 0.010936f
C143 VDD1.n113 VSUBS 0.010936f
C144 VDD1.n114 VSUBS 0.011579f
C145 VDD1.n115 VSUBS 0.025849f
C146 VDD1.n116 VSUBS 0.025849f
C147 VDD1.n117 VSUBS 0.025849f
C148 VDD1.n118 VSUBS 0.011258f
C149 VDD1.n119 VSUBS 0.010936f
C150 VDD1.n120 VSUBS 0.020352f
C151 VDD1.n121 VSUBS 0.020352f
C152 VDD1.n122 VSUBS 0.010936f
C153 VDD1.n123 VSUBS 0.011579f
C154 VDD1.n124 VSUBS 0.025849f
C155 VDD1.n125 VSUBS 0.025849f
C156 VDD1.n126 VSUBS 0.011579f
C157 VDD1.n127 VSUBS 0.010936f
C158 VDD1.n128 VSUBS 0.020352f
C159 VDD1.n129 VSUBS 0.020352f
C160 VDD1.n130 VSUBS 0.010936f
C161 VDD1.n131 VSUBS 0.011579f
C162 VDD1.n132 VSUBS 0.025849f
C163 VDD1.n133 VSUBS 0.025849f
C164 VDD1.n134 VSUBS 0.011579f
C165 VDD1.n135 VSUBS 0.010936f
C166 VDD1.n136 VSUBS 0.020352f
C167 VDD1.n137 VSUBS 0.020352f
C168 VDD1.n138 VSUBS 0.010936f
C169 VDD1.n139 VSUBS 0.011579f
C170 VDD1.n140 VSUBS 0.025849f
C171 VDD1.n141 VSUBS 0.063463f
C172 VDD1.n142 VSUBS 0.011579f
C173 VDD1.n143 VSUBS 0.010936f
C174 VDD1.n144 VSUBS 0.04593f
C175 VDD1.n145 VSUBS 0.598705f
C176 VP.t1 VSUBS 3.09143f
C177 VP.t0 VSUBS 2.84688f
C178 VP.n0 VSUBS 6.02613f
C179 VDD2.n0 VSUBS 0.022826f
C180 VDD2.n1 VSUBS 0.020536f
C181 VDD2.n2 VSUBS 0.011035f
C182 VDD2.n3 VSUBS 0.026082f
C183 VDD2.n4 VSUBS 0.011684f
C184 VDD2.n5 VSUBS 0.020536f
C185 VDD2.n6 VSUBS 0.011035f
C186 VDD2.n7 VSUBS 0.026082f
C187 VDD2.n8 VSUBS 0.011684f
C188 VDD2.n9 VSUBS 0.020536f
C189 VDD2.n10 VSUBS 0.011035f
C190 VDD2.n11 VSUBS 0.026082f
C191 VDD2.n12 VSUBS 0.011359f
C192 VDD2.n13 VSUBS 0.020536f
C193 VDD2.n14 VSUBS 0.011684f
C194 VDD2.n15 VSUBS 0.026082f
C195 VDD2.n16 VSUBS 0.011684f
C196 VDD2.n17 VSUBS 0.020536f
C197 VDD2.n18 VSUBS 0.011035f
C198 VDD2.n19 VSUBS 0.026082f
C199 VDD2.n20 VSUBS 0.011684f
C200 VDD2.n21 VSUBS 1.14574f
C201 VDD2.n22 VSUBS 0.011035f
C202 VDD2.t1 VSUBS 0.056308f
C203 VDD2.n23 VSUBS 0.175841f
C204 VDD2.n24 VSUBS 0.019621f
C205 VDD2.n25 VSUBS 0.019562f
C206 VDD2.n26 VSUBS 0.026082f
C207 VDD2.n27 VSUBS 0.011684f
C208 VDD2.n28 VSUBS 0.011035f
C209 VDD2.n29 VSUBS 0.020536f
C210 VDD2.n30 VSUBS 0.020536f
C211 VDD2.n31 VSUBS 0.011035f
C212 VDD2.n32 VSUBS 0.011684f
C213 VDD2.n33 VSUBS 0.026082f
C214 VDD2.n34 VSUBS 0.026082f
C215 VDD2.n35 VSUBS 0.011684f
C216 VDD2.n36 VSUBS 0.011035f
C217 VDD2.n37 VSUBS 0.020536f
C218 VDD2.n38 VSUBS 0.020536f
C219 VDD2.n39 VSUBS 0.011035f
C220 VDD2.n40 VSUBS 0.011035f
C221 VDD2.n41 VSUBS 0.011684f
C222 VDD2.n42 VSUBS 0.026082f
C223 VDD2.n43 VSUBS 0.026082f
C224 VDD2.n44 VSUBS 0.026082f
C225 VDD2.n45 VSUBS 0.011359f
C226 VDD2.n46 VSUBS 0.011035f
C227 VDD2.n47 VSUBS 0.020536f
C228 VDD2.n48 VSUBS 0.020536f
C229 VDD2.n49 VSUBS 0.011035f
C230 VDD2.n50 VSUBS 0.011684f
C231 VDD2.n51 VSUBS 0.026082f
C232 VDD2.n52 VSUBS 0.026082f
C233 VDD2.n53 VSUBS 0.011684f
C234 VDD2.n54 VSUBS 0.011035f
C235 VDD2.n55 VSUBS 0.020536f
C236 VDD2.n56 VSUBS 0.020536f
C237 VDD2.n57 VSUBS 0.011035f
C238 VDD2.n58 VSUBS 0.011684f
C239 VDD2.n59 VSUBS 0.026082f
C240 VDD2.n60 VSUBS 0.026082f
C241 VDD2.n61 VSUBS 0.011684f
C242 VDD2.n62 VSUBS 0.011035f
C243 VDD2.n63 VSUBS 0.020536f
C244 VDD2.n64 VSUBS 0.020536f
C245 VDD2.n65 VSUBS 0.011035f
C246 VDD2.n66 VSUBS 0.011684f
C247 VDD2.n67 VSUBS 0.026082f
C248 VDD2.n68 VSUBS 0.064036f
C249 VDD2.n69 VSUBS 0.011684f
C250 VDD2.n70 VSUBS 0.011035f
C251 VDD2.n71 VSUBS 0.046345f
C252 VDD2.n72 VSUBS 0.573145f
C253 VDD2.n73 VSUBS 0.022826f
C254 VDD2.n74 VSUBS 0.020536f
C255 VDD2.n75 VSUBS 0.011035f
C256 VDD2.n76 VSUBS 0.026082f
C257 VDD2.n77 VSUBS 0.011684f
C258 VDD2.n78 VSUBS 0.020536f
C259 VDD2.n79 VSUBS 0.011035f
C260 VDD2.n80 VSUBS 0.026082f
C261 VDD2.n81 VSUBS 0.011684f
C262 VDD2.n82 VSUBS 0.020536f
C263 VDD2.n83 VSUBS 0.011035f
C264 VDD2.n84 VSUBS 0.026082f
C265 VDD2.n85 VSUBS 0.011359f
C266 VDD2.n86 VSUBS 0.020536f
C267 VDD2.n87 VSUBS 0.011359f
C268 VDD2.n88 VSUBS 0.011035f
C269 VDD2.n89 VSUBS 0.026082f
C270 VDD2.n90 VSUBS 0.026082f
C271 VDD2.n91 VSUBS 0.011684f
C272 VDD2.n92 VSUBS 0.020536f
C273 VDD2.n93 VSUBS 0.011035f
C274 VDD2.n94 VSUBS 0.026082f
C275 VDD2.n95 VSUBS 0.011684f
C276 VDD2.n96 VSUBS 1.14574f
C277 VDD2.n97 VSUBS 0.011035f
C278 VDD2.t0 VSUBS 0.056308f
C279 VDD2.n98 VSUBS 0.175841f
C280 VDD2.n99 VSUBS 0.019621f
C281 VDD2.n100 VSUBS 0.019562f
C282 VDD2.n101 VSUBS 0.026082f
C283 VDD2.n102 VSUBS 0.011684f
C284 VDD2.n103 VSUBS 0.011035f
C285 VDD2.n104 VSUBS 0.020536f
C286 VDD2.n105 VSUBS 0.020536f
C287 VDD2.n106 VSUBS 0.011035f
C288 VDD2.n107 VSUBS 0.011684f
C289 VDD2.n108 VSUBS 0.026082f
C290 VDD2.n109 VSUBS 0.026082f
C291 VDD2.n110 VSUBS 0.011684f
C292 VDD2.n111 VSUBS 0.011035f
C293 VDD2.n112 VSUBS 0.020536f
C294 VDD2.n113 VSUBS 0.020536f
C295 VDD2.n114 VSUBS 0.011035f
C296 VDD2.n115 VSUBS 0.011684f
C297 VDD2.n116 VSUBS 0.026082f
C298 VDD2.n117 VSUBS 0.026082f
C299 VDD2.n118 VSUBS 0.011684f
C300 VDD2.n119 VSUBS 0.011035f
C301 VDD2.n120 VSUBS 0.020536f
C302 VDD2.n121 VSUBS 0.020536f
C303 VDD2.n122 VSUBS 0.011035f
C304 VDD2.n123 VSUBS 0.011684f
C305 VDD2.n124 VSUBS 0.026082f
C306 VDD2.n125 VSUBS 0.026082f
C307 VDD2.n126 VSUBS 0.011684f
C308 VDD2.n127 VSUBS 0.011035f
C309 VDD2.n128 VSUBS 0.020536f
C310 VDD2.n129 VSUBS 0.020536f
C311 VDD2.n130 VSUBS 0.011035f
C312 VDD2.n131 VSUBS 0.011684f
C313 VDD2.n132 VSUBS 0.026082f
C314 VDD2.n133 VSUBS 0.026082f
C315 VDD2.n134 VSUBS 0.011684f
C316 VDD2.n135 VSUBS 0.011035f
C317 VDD2.n136 VSUBS 0.020536f
C318 VDD2.n137 VSUBS 0.020536f
C319 VDD2.n138 VSUBS 0.011035f
C320 VDD2.n139 VSUBS 0.011684f
C321 VDD2.n140 VSUBS 0.026082f
C322 VDD2.n141 VSUBS 0.064036f
C323 VDD2.n142 VSUBS 0.011684f
C324 VDD2.n143 VSUBS 0.011035f
C325 VDD2.n144 VSUBS 0.046345f
C326 VDD2.n145 VSUBS 0.046397f
C327 VDD2.n146 VSUBS 2.39245f
C328 VTAIL.n0 VSUBS 0.031592f
C329 VTAIL.n1 VSUBS 0.028421f
C330 VTAIL.n2 VSUBS 0.015272f
C331 VTAIL.n3 VSUBS 0.036099f
C332 VTAIL.n4 VSUBS 0.016171f
C333 VTAIL.n5 VSUBS 0.028421f
C334 VTAIL.n6 VSUBS 0.015272f
C335 VTAIL.n7 VSUBS 0.036099f
C336 VTAIL.n8 VSUBS 0.016171f
C337 VTAIL.n9 VSUBS 0.028421f
C338 VTAIL.n10 VSUBS 0.015272f
C339 VTAIL.n11 VSUBS 0.036099f
C340 VTAIL.n12 VSUBS 0.015722f
C341 VTAIL.n13 VSUBS 0.028421f
C342 VTAIL.n14 VSUBS 0.016171f
C343 VTAIL.n15 VSUBS 0.036099f
C344 VTAIL.n16 VSUBS 0.016171f
C345 VTAIL.n17 VSUBS 0.028421f
C346 VTAIL.n18 VSUBS 0.015272f
C347 VTAIL.n19 VSUBS 0.036099f
C348 VTAIL.n20 VSUBS 0.016171f
C349 VTAIL.n21 VSUBS 1.58574f
C350 VTAIL.n22 VSUBS 0.015272f
C351 VTAIL.t0 VSUBS 0.077932f
C352 VTAIL.n23 VSUBS 0.243367f
C353 VTAIL.n24 VSUBS 0.027155f
C354 VTAIL.n25 VSUBS 0.027074f
C355 VTAIL.n26 VSUBS 0.036099f
C356 VTAIL.n27 VSUBS 0.016171f
C357 VTAIL.n28 VSUBS 0.015272f
C358 VTAIL.n29 VSUBS 0.028421f
C359 VTAIL.n30 VSUBS 0.028421f
C360 VTAIL.n31 VSUBS 0.015272f
C361 VTAIL.n32 VSUBS 0.016171f
C362 VTAIL.n33 VSUBS 0.036099f
C363 VTAIL.n34 VSUBS 0.036099f
C364 VTAIL.n35 VSUBS 0.016171f
C365 VTAIL.n36 VSUBS 0.015272f
C366 VTAIL.n37 VSUBS 0.028421f
C367 VTAIL.n38 VSUBS 0.028421f
C368 VTAIL.n39 VSUBS 0.015272f
C369 VTAIL.n40 VSUBS 0.015272f
C370 VTAIL.n41 VSUBS 0.016171f
C371 VTAIL.n42 VSUBS 0.036099f
C372 VTAIL.n43 VSUBS 0.036099f
C373 VTAIL.n44 VSUBS 0.036099f
C374 VTAIL.n45 VSUBS 0.015722f
C375 VTAIL.n46 VSUBS 0.015272f
C376 VTAIL.n47 VSUBS 0.028421f
C377 VTAIL.n48 VSUBS 0.028421f
C378 VTAIL.n49 VSUBS 0.015272f
C379 VTAIL.n50 VSUBS 0.016171f
C380 VTAIL.n51 VSUBS 0.036099f
C381 VTAIL.n52 VSUBS 0.036099f
C382 VTAIL.n53 VSUBS 0.016171f
C383 VTAIL.n54 VSUBS 0.015272f
C384 VTAIL.n55 VSUBS 0.028421f
C385 VTAIL.n56 VSUBS 0.028421f
C386 VTAIL.n57 VSUBS 0.015272f
C387 VTAIL.n58 VSUBS 0.016171f
C388 VTAIL.n59 VSUBS 0.036099f
C389 VTAIL.n60 VSUBS 0.036099f
C390 VTAIL.n61 VSUBS 0.016171f
C391 VTAIL.n62 VSUBS 0.015272f
C392 VTAIL.n63 VSUBS 0.028421f
C393 VTAIL.n64 VSUBS 0.028421f
C394 VTAIL.n65 VSUBS 0.015272f
C395 VTAIL.n66 VSUBS 0.016171f
C396 VTAIL.n67 VSUBS 0.036099f
C397 VTAIL.n68 VSUBS 0.088628f
C398 VTAIL.n69 VSUBS 0.016171f
C399 VTAIL.n70 VSUBS 0.015272f
C400 VTAIL.n71 VSUBS 0.064142f
C401 VTAIL.n72 VSUBS 0.044577f
C402 VTAIL.n73 VSUBS 1.78081f
C403 VTAIL.n74 VSUBS 0.031592f
C404 VTAIL.n75 VSUBS 0.028421f
C405 VTAIL.n76 VSUBS 0.015272f
C406 VTAIL.n77 VSUBS 0.036099f
C407 VTAIL.n78 VSUBS 0.016171f
C408 VTAIL.n79 VSUBS 0.028421f
C409 VTAIL.n80 VSUBS 0.015272f
C410 VTAIL.n81 VSUBS 0.036099f
C411 VTAIL.n82 VSUBS 0.016171f
C412 VTAIL.n83 VSUBS 0.028421f
C413 VTAIL.n84 VSUBS 0.015272f
C414 VTAIL.n85 VSUBS 0.036099f
C415 VTAIL.n86 VSUBS 0.015722f
C416 VTAIL.n87 VSUBS 0.028421f
C417 VTAIL.n88 VSUBS 0.015722f
C418 VTAIL.n89 VSUBS 0.015272f
C419 VTAIL.n90 VSUBS 0.036099f
C420 VTAIL.n91 VSUBS 0.036099f
C421 VTAIL.n92 VSUBS 0.016171f
C422 VTAIL.n93 VSUBS 0.028421f
C423 VTAIL.n94 VSUBS 0.015272f
C424 VTAIL.n95 VSUBS 0.036099f
C425 VTAIL.n96 VSUBS 0.016171f
C426 VTAIL.n97 VSUBS 1.58574f
C427 VTAIL.n98 VSUBS 0.015272f
C428 VTAIL.t3 VSUBS 0.077932f
C429 VTAIL.n99 VSUBS 0.243367f
C430 VTAIL.n100 VSUBS 0.027155f
C431 VTAIL.n101 VSUBS 0.027074f
C432 VTAIL.n102 VSUBS 0.036099f
C433 VTAIL.n103 VSUBS 0.016171f
C434 VTAIL.n104 VSUBS 0.015272f
C435 VTAIL.n105 VSUBS 0.028421f
C436 VTAIL.n106 VSUBS 0.028421f
C437 VTAIL.n107 VSUBS 0.015272f
C438 VTAIL.n108 VSUBS 0.016171f
C439 VTAIL.n109 VSUBS 0.036099f
C440 VTAIL.n110 VSUBS 0.036099f
C441 VTAIL.n111 VSUBS 0.016171f
C442 VTAIL.n112 VSUBS 0.015272f
C443 VTAIL.n113 VSUBS 0.028421f
C444 VTAIL.n114 VSUBS 0.028421f
C445 VTAIL.n115 VSUBS 0.015272f
C446 VTAIL.n116 VSUBS 0.016171f
C447 VTAIL.n117 VSUBS 0.036099f
C448 VTAIL.n118 VSUBS 0.036099f
C449 VTAIL.n119 VSUBS 0.016171f
C450 VTAIL.n120 VSUBS 0.015272f
C451 VTAIL.n121 VSUBS 0.028421f
C452 VTAIL.n122 VSUBS 0.028421f
C453 VTAIL.n123 VSUBS 0.015272f
C454 VTAIL.n124 VSUBS 0.016171f
C455 VTAIL.n125 VSUBS 0.036099f
C456 VTAIL.n126 VSUBS 0.036099f
C457 VTAIL.n127 VSUBS 0.016171f
C458 VTAIL.n128 VSUBS 0.015272f
C459 VTAIL.n129 VSUBS 0.028421f
C460 VTAIL.n130 VSUBS 0.028421f
C461 VTAIL.n131 VSUBS 0.015272f
C462 VTAIL.n132 VSUBS 0.016171f
C463 VTAIL.n133 VSUBS 0.036099f
C464 VTAIL.n134 VSUBS 0.036099f
C465 VTAIL.n135 VSUBS 0.016171f
C466 VTAIL.n136 VSUBS 0.015272f
C467 VTAIL.n137 VSUBS 0.028421f
C468 VTAIL.n138 VSUBS 0.028421f
C469 VTAIL.n139 VSUBS 0.015272f
C470 VTAIL.n140 VSUBS 0.016171f
C471 VTAIL.n141 VSUBS 0.036099f
C472 VTAIL.n142 VSUBS 0.088628f
C473 VTAIL.n143 VSUBS 0.016171f
C474 VTAIL.n144 VSUBS 0.015272f
C475 VTAIL.n145 VSUBS 0.064142f
C476 VTAIL.n146 VSUBS 0.044577f
C477 VTAIL.n147 VSUBS 1.80371f
C478 VTAIL.n148 VSUBS 0.031592f
C479 VTAIL.n149 VSUBS 0.028421f
C480 VTAIL.n150 VSUBS 0.015272f
C481 VTAIL.n151 VSUBS 0.036099f
C482 VTAIL.n152 VSUBS 0.016171f
C483 VTAIL.n153 VSUBS 0.028421f
C484 VTAIL.n154 VSUBS 0.015272f
C485 VTAIL.n155 VSUBS 0.036099f
C486 VTAIL.n156 VSUBS 0.016171f
C487 VTAIL.n157 VSUBS 0.028421f
C488 VTAIL.n158 VSUBS 0.015272f
C489 VTAIL.n159 VSUBS 0.036099f
C490 VTAIL.n160 VSUBS 0.015722f
C491 VTAIL.n161 VSUBS 0.028421f
C492 VTAIL.n162 VSUBS 0.015722f
C493 VTAIL.n163 VSUBS 0.015272f
C494 VTAIL.n164 VSUBS 0.036099f
C495 VTAIL.n165 VSUBS 0.036099f
C496 VTAIL.n166 VSUBS 0.016171f
C497 VTAIL.n167 VSUBS 0.028421f
C498 VTAIL.n168 VSUBS 0.015272f
C499 VTAIL.n169 VSUBS 0.036099f
C500 VTAIL.n170 VSUBS 0.016171f
C501 VTAIL.n171 VSUBS 1.58574f
C502 VTAIL.n172 VSUBS 0.015272f
C503 VTAIL.t1 VSUBS 0.077932f
C504 VTAIL.n173 VSUBS 0.243367f
C505 VTAIL.n174 VSUBS 0.027155f
C506 VTAIL.n175 VSUBS 0.027074f
C507 VTAIL.n176 VSUBS 0.036099f
C508 VTAIL.n177 VSUBS 0.016171f
C509 VTAIL.n178 VSUBS 0.015272f
C510 VTAIL.n179 VSUBS 0.028421f
C511 VTAIL.n180 VSUBS 0.028421f
C512 VTAIL.n181 VSUBS 0.015272f
C513 VTAIL.n182 VSUBS 0.016171f
C514 VTAIL.n183 VSUBS 0.036099f
C515 VTAIL.n184 VSUBS 0.036099f
C516 VTAIL.n185 VSUBS 0.016171f
C517 VTAIL.n186 VSUBS 0.015272f
C518 VTAIL.n187 VSUBS 0.028421f
C519 VTAIL.n188 VSUBS 0.028421f
C520 VTAIL.n189 VSUBS 0.015272f
C521 VTAIL.n190 VSUBS 0.016171f
C522 VTAIL.n191 VSUBS 0.036099f
C523 VTAIL.n192 VSUBS 0.036099f
C524 VTAIL.n193 VSUBS 0.016171f
C525 VTAIL.n194 VSUBS 0.015272f
C526 VTAIL.n195 VSUBS 0.028421f
C527 VTAIL.n196 VSUBS 0.028421f
C528 VTAIL.n197 VSUBS 0.015272f
C529 VTAIL.n198 VSUBS 0.016171f
C530 VTAIL.n199 VSUBS 0.036099f
C531 VTAIL.n200 VSUBS 0.036099f
C532 VTAIL.n201 VSUBS 0.016171f
C533 VTAIL.n202 VSUBS 0.015272f
C534 VTAIL.n203 VSUBS 0.028421f
C535 VTAIL.n204 VSUBS 0.028421f
C536 VTAIL.n205 VSUBS 0.015272f
C537 VTAIL.n206 VSUBS 0.016171f
C538 VTAIL.n207 VSUBS 0.036099f
C539 VTAIL.n208 VSUBS 0.036099f
C540 VTAIL.n209 VSUBS 0.016171f
C541 VTAIL.n210 VSUBS 0.015272f
C542 VTAIL.n211 VSUBS 0.028421f
C543 VTAIL.n212 VSUBS 0.028421f
C544 VTAIL.n213 VSUBS 0.015272f
C545 VTAIL.n214 VSUBS 0.016171f
C546 VTAIL.n215 VSUBS 0.036099f
C547 VTAIL.n216 VSUBS 0.088628f
C548 VTAIL.n217 VSUBS 0.016171f
C549 VTAIL.n218 VSUBS 0.015272f
C550 VTAIL.n219 VSUBS 0.064142f
C551 VTAIL.n220 VSUBS 0.044577f
C552 VTAIL.n221 VSUBS 1.69081f
C553 VTAIL.n222 VSUBS 0.031592f
C554 VTAIL.n223 VSUBS 0.028421f
C555 VTAIL.n224 VSUBS 0.015272f
C556 VTAIL.n225 VSUBS 0.036099f
C557 VTAIL.n226 VSUBS 0.016171f
C558 VTAIL.n227 VSUBS 0.028421f
C559 VTAIL.n228 VSUBS 0.015272f
C560 VTAIL.n229 VSUBS 0.036099f
C561 VTAIL.n230 VSUBS 0.016171f
C562 VTAIL.n231 VSUBS 0.028421f
C563 VTAIL.n232 VSUBS 0.015272f
C564 VTAIL.n233 VSUBS 0.036099f
C565 VTAIL.n234 VSUBS 0.015722f
C566 VTAIL.n235 VSUBS 0.028421f
C567 VTAIL.n236 VSUBS 0.016171f
C568 VTAIL.n237 VSUBS 0.036099f
C569 VTAIL.n238 VSUBS 0.016171f
C570 VTAIL.n239 VSUBS 0.028421f
C571 VTAIL.n240 VSUBS 0.015272f
C572 VTAIL.n241 VSUBS 0.036099f
C573 VTAIL.n242 VSUBS 0.016171f
C574 VTAIL.n243 VSUBS 1.58574f
C575 VTAIL.n244 VSUBS 0.015272f
C576 VTAIL.t2 VSUBS 0.077932f
C577 VTAIL.n245 VSUBS 0.243367f
C578 VTAIL.n246 VSUBS 0.027155f
C579 VTAIL.n247 VSUBS 0.027074f
C580 VTAIL.n248 VSUBS 0.036099f
C581 VTAIL.n249 VSUBS 0.016171f
C582 VTAIL.n250 VSUBS 0.015272f
C583 VTAIL.n251 VSUBS 0.028421f
C584 VTAIL.n252 VSUBS 0.028421f
C585 VTAIL.n253 VSUBS 0.015272f
C586 VTAIL.n254 VSUBS 0.016171f
C587 VTAIL.n255 VSUBS 0.036099f
C588 VTAIL.n256 VSUBS 0.036099f
C589 VTAIL.n257 VSUBS 0.016171f
C590 VTAIL.n258 VSUBS 0.015272f
C591 VTAIL.n259 VSUBS 0.028421f
C592 VTAIL.n260 VSUBS 0.028421f
C593 VTAIL.n261 VSUBS 0.015272f
C594 VTAIL.n262 VSUBS 0.015272f
C595 VTAIL.n263 VSUBS 0.016171f
C596 VTAIL.n264 VSUBS 0.036099f
C597 VTAIL.n265 VSUBS 0.036099f
C598 VTAIL.n266 VSUBS 0.036099f
C599 VTAIL.n267 VSUBS 0.015722f
C600 VTAIL.n268 VSUBS 0.015272f
C601 VTAIL.n269 VSUBS 0.028421f
C602 VTAIL.n270 VSUBS 0.028421f
C603 VTAIL.n271 VSUBS 0.015272f
C604 VTAIL.n272 VSUBS 0.016171f
C605 VTAIL.n273 VSUBS 0.036099f
C606 VTAIL.n274 VSUBS 0.036099f
C607 VTAIL.n275 VSUBS 0.016171f
C608 VTAIL.n276 VSUBS 0.015272f
C609 VTAIL.n277 VSUBS 0.028421f
C610 VTAIL.n278 VSUBS 0.028421f
C611 VTAIL.n279 VSUBS 0.015272f
C612 VTAIL.n280 VSUBS 0.016171f
C613 VTAIL.n281 VSUBS 0.036099f
C614 VTAIL.n282 VSUBS 0.036099f
C615 VTAIL.n283 VSUBS 0.016171f
C616 VTAIL.n284 VSUBS 0.015272f
C617 VTAIL.n285 VSUBS 0.028421f
C618 VTAIL.n286 VSUBS 0.028421f
C619 VTAIL.n287 VSUBS 0.015272f
C620 VTAIL.n288 VSUBS 0.016171f
C621 VTAIL.n289 VSUBS 0.036099f
C622 VTAIL.n290 VSUBS 0.088628f
C623 VTAIL.n291 VSUBS 0.016171f
C624 VTAIL.n292 VSUBS 0.015272f
C625 VTAIL.n293 VSUBS 0.064142f
C626 VTAIL.n294 VSUBS 0.044577f
C627 VTAIL.n295 VSUBS 1.61423f
C628 VN.t0 VSUBS 2.73293f
C629 VN.t1 VSUBS 2.97255f
C630 B.n0 VSUBS 0.005995f
C631 B.n1 VSUBS 0.005995f
C632 B.n2 VSUBS 0.008866f
C633 B.n3 VSUBS 0.006794f
C634 B.n4 VSUBS 0.006794f
C635 B.n5 VSUBS 0.006794f
C636 B.n6 VSUBS 0.006794f
C637 B.n7 VSUBS 0.006794f
C638 B.n8 VSUBS 0.006794f
C639 B.n9 VSUBS 0.006794f
C640 B.n10 VSUBS 0.016136f
C641 B.n11 VSUBS 0.006794f
C642 B.n12 VSUBS 0.006794f
C643 B.n13 VSUBS 0.006794f
C644 B.n14 VSUBS 0.006794f
C645 B.n15 VSUBS 0.006794f
C646 B.n16 VSUBS 0.006794f
C647 B.n17 VSUBS 0.006794f
C648 B.n18 VSUBS 0.006794f
C649 B.n19 VSUBS 0.006794f
C650 B.n20 VSUBS 0.006794f
C651 B.n21 VSUBS 0.006794f
C652 B.n22 VSUBS 0.006794f
C653 B.n23 VSUBS 0.006794f
C654 B.n24 VSUBS 0.006794f
C655 B.n25 VSUBS 0.006794f
C656 B.n26 VSUBS 0.006794f
C657 B.n27 VSUBS 0.006794f
C658 B.n28 VSUBS 0.006794f
C659 B.n29 VSUBS 0.006794f
C660 B.n30 VSUBS 0.006794f
C661 B.n31 VSUBS 0.006794f
C662 B.n32 VSUBS 0.006794f
C663 B.n33 VSUBS 0.006794f
C664 B.t10 VSUBS 0.238267f
C665 B.t11 VSUBS 0.254268f
C666 B.t9 VSUBS 0.611029f
C667 B.n34 VSUBS 0.3632f
C668 B.n35 VSUBS 0.258283f
C669 B.n36 VSUBS 0.006794f
C670 B.n37 VSUBS 0.006794f
C671 B.n38 VSUBS 0.006794f
C672 B.n39 VSUBS 0.006794f
C673 B.t1 VSUBS 0.23827f
C674 B.t2 VSUBS 0.254271f
C675 B.t0 VSUBS 0.611029f
C676 B.n40 VSUBS 0.363197f
C677 B.n41 VSUBS 0.25828f
C678 B.n42 VSUBS 0.015741f
C679 B.n43 VSUBS 0.006794f
C680 B.n44 VSUBS 0.006794f
C681 B.n45 VSUBS 0.006794f
C682 B.n46 VSUBS 0.006794f
C683 B.n47 VSUBS 0.006794f
C684 B.n48 VSUBS 0.006794f
C685 B.n49 VSUBS 0.006794f
C686 B.n50 VSUBS 0.006794f
C687 B.n51 VSUBS 0.006794f
C688 B.n52 VSUBS 0.006794f
C689 B.n53 VSUBS 0.006794f
C690 B.n54 VSUBS 0.006794f
C691 B.n55 VSUBS 0.006794f
C692 B.n56 VSUBS 0.006794f
C693 B.n57 VSUBS 0.006794f
C694 B.n58 VSUBS 0.006794f
C695 B.n59 VSUBS 0.006794f
C696 B.n60 VSUBS 0.006794f
C697 B.n61 VSUBS 0.006794f
C698 B.n62 VSUBS 0.006794f
C699 B.n63 VSUBS 0.006794f
C700 B.n64 VSUBS 0.006794f
C701 B.n65 VSUBS 0.016136f
C702 B.n66 VSUBS 0.006794f
C703 B.n67 VSUBS 0.006794f
C704 B.n68 VSUBS 0.006794f
C705 B.n69 VSUBS 0.006794f
C706 B.n70 VSUBS 0.006794f
C707 B.n71 VSUBS 0.006794f
C708 B.n72 VSUBS 0.006794f
C709 B.n73 VSUBS 0.006794f
C710 B.n74 VSUBS 0.006794f
C711 B.n75 VSUBS 0.006794f
C712 B.n76 VSUBS 0.006794f
C713 B.n77 VSUBS 0.006794f
C714 B.n78 VSUBS 0.006794f
C715 B.n79 VSUBS 0.006794f
C716 B.n80 VSUBS 0.006794f
C717 B.n81 VSUBS 0.006794f
C718 B.n82 VSUBS 0.016056f
C719 B.n83 VSUBS 0.006794f
C720 B.n84 VSUBS 0.006794f
C721 B.n85 VSUBS 0.006794f
C722 B.n86 VSUBS 0.006794f
C723 B.n87 VSUBS 0.006794f
C724 B.n88 VSUBS 0.006794f
C725 B.n89 VSUBS 0.006794f
C726 B.n90 VSUBS 0.006794f
C727 B.n91 VSUBS 0.006794f
C728 B.n92 VSUBS 0.006794f
C729 B.n93 VSUBS 0.006794f
C730 B.n94 VSUBS 0.006794f
C731 B.n95 VSUBS 0.006794f
C732 B.n96 VSUBS 0.006794f
C733 B.n97 VSUBS 0.006794f
C734 B.n98 VSUBS 0.006794f
C735 B.n99 VSUBS 0.006794f
C736 B.n100 VSUBS 0.006794f
C737 B.n101 VSUBS 0.006794f
C738 B.n102 VSUBS 0.006794f
C739 B.n103 VSUBS 0.006794f
C740 B.n104 VSUBS 0.006794f
C741 B.n105 VSUBS 0.006794f
C742 B.t8 VSUBS 0.23827f
C743 B.t7 VSUBS 0.254271f
C744 B.t6 VSUBS 0.611029f
C745 B.n106 VSUBS 0.363197f
C746 B.n107 VSUBS 0.25828f
C747 B.n108 VSUBS 0.006794f
C748 B.n109 VSUBS 0.006794f
C749 B.n110 VSUBS 0.006794f
C750 B.n111 VSUBS 0.006794f
C751 B.n112 VSUBS 0.003997f
C752 B.n113 VSUBS 0.006794f
C753 B.n114 VSUBS 0.006794f
C754 B.n115 VSUBS 0.006794f
C755 B.n116 VSUBS 0.006794f
C756 B.n117 VSUBS 0.006794f
C757 B.n118 VSUBS 0.006794f
C758 B.n119 VSUBS 0.006794f
C759 B.n120 VSUBS 0.006794f
C760 B.n121 VSUBS 0.006794f
C761 B.n122 VSUBS 0.006794f
C762 B.n123 VSUBS 0.006794f
C763 B.n124 VSUBS 0.006794f
C764 B.n125 VSUBS 0.006794f
C765 B.n126 VSUBS 0.006794f
C766 B.n127 VSUBS 0.006794f
C767 B.n128 VSUBS 0.006794f
C768 B.n129 VSUBS 0.006794f
C769 B.n130 VSUBS 0.006794f
C770 B.n131 VSUBS 0.006794f
C771 B.n132 VSUBS 0.006794f
C772 B.n133 VSUBS 0.006794f
C773 B.n134 VSUBS 0.006794f
C774 B.n135 VSUBS 0.016136f
C775 B.n136 VSUBS 0.006794f
C776 B.n137 VSUBS 0.006794f
C777 B.n138 VSUBS 0.006794f
C778 B.n139 VSUBS 0.006794f
C779 B.n140 VSUBS 0.006794f
C780 B.n141 VSUBS 0.006794f
C781 B.n142 VSUBS 0.006794f
C782 B.n143 VSUBS 0.006794f
C783 B.n144 VSUBS 0.006794f
C784 B.n145 VSUBS 0.006794f
C785 B.n146 VSUBS 0.006794f
C786 B.n147 VSUBS 0.006794f
C787 B.n148 VSUBS 0.006794f
C788 B.n149 VSUBS 0.006794f
C789 B.n150 VSUBS 0.006794f
C790 B.n151 VSUBS 0.006794f
C791 B.n152 VSUBS 0.006794f
C792 B.n153 VSUBS 0.006794f
C793 B.n154 VSUBS 0.006794f
C794 B.n155 VSUBS 0.006794f
C795 B.n156 VSUBS 0.006794f
C796 B.n157 VSUBS 0.006794f
C797 B.n158 VSUBS 0.006794f
C798 B.n159 VSUBS 0.006794f
C799 B.n160 VSUBS 0.006794f
C800 B.n161 VSUBS 0.006794f
C801 B.n162 VSUBS 0.006794f
C802 B.n163 VSUBS 0.006794f
C803 B.n164 VSUBS 0.015237f
C804 B.n165 VSUBS 0.015237f
C805 B.n166 VSUBS 0.016136f
C806 B.n167 VSUBS 0.006794f
C807 B.n168 VSUBS 0.006794f
C808 B.n169 VSUBS 0.006794f
C809 B.n170 VSUBS 0.006794f
C810 B.n171 VSUBS 0.006794f
C811 B.n172 VSUBS 0.006794f
C812 B.n173 VSUBS 0.006794f
C813 B.n174 VSUBS 0.006794f
C814 B.n175 VSUBS 0.006794f
C815 B.n176 VSUBS 0.006794f
C816 B.n177 VSUBS 0.006794f
C817 B.n178 VSUBS 0.006794f
C818 B.n179 VSUBS 0.006794f
C819 B.n180 VSUBS 0.006794f
C820 B.n181 VSUBS 0.006794f
C821 B.n182 VSUBS 0.006794f
C822 B.n183 VSUBS 0.006794f
C823 B.n184 VSUBS 0.006794f
C824 B.n185 VSUBS 0.006794f
C825 B.n186 VSUBS 0.006794f
C826 B.n187 VSUBS 0.006794f
C827 B.n188 VSUBS 0.006794f
C828 B.n189 VSUBS 0.006794f
C829 B.n190 VSUBS 0.006794f
C830 B.n191 VSUBS 0.006794f
C831 B.n192 VSUBS 0.006794f
C832 B.n193 VSUBS 0.006794f
C833 B.n194 VSUBS 0.006794f
C834 B.n195 VSUBS 0.006794f
C835 B.n196 VSUBS 0.006794f
C836 B.n197 VSUBS 0.006794f
C837 B.n198 VSUBS 0.006794f
C838 B.n199 VSUBS 0.006794f
C839 B.n200 VSUBS 0.006794f
C840 B.n201 VSUBS 0.006794f
C841 B.n202 VSUBS 0.006794f
C842 B.n203 VSUBS 0.006794f
C843 B.n204 VSUBS 0.006794f
C844 B.n205 VSUBS 0.006794f
C845 B.n206 VSUBS 0.006794f
C846 B.n207 VSUBS 0.006794f
C847 B.n208 VSUBS 0.006794f
C848 B.n209 VSUBS 0.006794f
C849 B.n210 VSUBS 0.006794f
C850 B.n211 VSUBS 0.006794f
C851 B.n212 VSUBS 0.006794f
C852 B.n213 VSUBS 0.006794f
C853 B.n214 VSUBS 0.006794f
C854 B.n215 VSUBS 0.006794f
C855 B.n216 VSUBS 0.006794f
C856 B.n217 VSUBS 0.006794f
C857 B.n218 VSUBS 0.006794f
C858 B.n219 VSUBS 0.006794f
C859 B.n220 VSUBS 0.006794f
C860 B.n221 VSUBS 0.006794f
C861 B.n222 VSUBS 0.006794f
C862 B.n223 VSUBS 0.006794f
C863 B.n224 VSUBS 0.006794f
C864 B.n225 VSUBS 0.006794f
C865 B.n226 VSUBS 0.006794f
C866 B.n227 VSUBS 0.006794f
C867 B.n228 VSUBS 0.006794f
C868 B.n229 VSUBS 0.006794f
C869 B.n230 VSUBS 0.006794f
C870 B.n231 VSUBS 0.006794f
C871 B.n232 VSUBS 0.006794f
C872 B.t5 VSUBS 0.238267f
C873 B.t4 VSUBS 0.254268f
C874 B.t3 VSUBS 0.611029f
C875 B.n233 VSUBS 0.3632f
C876 B.n234 VSUBS 0.258283f
C877 B.n235 VSUBS 0.015741f
C878 B.n236 VSUBS 0.006195f
C879 B.n237 VSUBS 0.006794f
C880 B.n238 VSUBS 0.006794f
C881 B.n239 VSUBS 0.006794f
C882 B.n240 VSUBS 0.006794f
C883 B.n241 VSUBS 0.006794f
C884 B.n242 VSUBS 0.006794f
C885 B.n243 VSUBS 0.006794f
C886 B.n244 VSUBS 0.006794f
C887 B.n245 VSUBS 0.006794f
C888 B.n246 VSUBS 0.006794f
C889 B.n247 VSUBS 0.006794f
C890 B.n248 VSUBS 0.006794f
C891 B.n249 VSUBS 0.006794f
C892 B.n250 VSUBS 0.006794f
C893 B.n251 VSUBS 0.006794f
C894 B.n252 VSUBS 0.003997f
C895 B.n253 VSUBS 0.015741f
C896 B.n254 VSUBS 0.006195f
C897 B.n255 VSUBS 0.006794f
C898 B.n256 VSUBS 0.006794f
C899 B.n257 VSUBS 0.006794f
C900 B.n258 VSUBS 0.006794f
C901 B.n259 VSUBS 0.006794f
C902 B.n260 VSUBS 0.006794f
C903 B.n261 VSUBS 0.006794f
C904 B.n262 VSUBS 0.006794f
C905 B.n263 VSUBS 0.006794f
C906 B.n264 VSUBS 0.006794f
C907 B.n265 VSUBS 0.006794f
C908 B.n266 VSUBS 0.006794f
C909 B.n267 VSUBS 0.006794f
C910 B.n268 VSUBS 0.006794f
C911 B.n269 VSUBS 0.006794f
C912 B.n270 VSUBS 0.006794f
C913 B.n271 VSUBS 0.006794f
C914 B.n272 VSUBS 0.006794f
C915 B.n273 VSUBS 0.006794f
C916 B.n274 VSUBS 0.006794f
C917 B.n275 VSUBS 0.006794f
C918 B.n276 VSUBS 0.006794f
C919 B.n277 VSUBS 0.006794f
C920 B.n278 VSUBS 0.006794f
C921 B.n279 VSUBS 0.006794f
C922 B.n280 VSUBS 0.006794f
C923 B.n281 VSUBS 0.006794f
C924 B.n282 VSUBS 0.006794f
C925 B.n283 VSUBS 0.006794f
C926 B.n284 VSUBS 0.006794f
C927 B.n285 VSUBS 0.006794f
C928 B.n286 VSUBS 0.006794f
C929 B.n287 VSUBS 0.006794f
C930 B.n288 VSUBS 0.006794f
C931 B.n289 VSUBS 0.006794f
C932 B.n290 VSUBS 0.006794f
C933 B.n291 VSUBS 0.006794f
C934 B.n292 VSUBS 0.006794f
C935 B.n293 VSUBS 0.006794f
C936 B.n294 VSUBS 0.006794f
C937 B.n295 VSUBS 0.006794f
C938 B.n296 VSUBS 0.006794f
C939 B.n297 VSUBS 0.006794f
C940 B.n298 VSUBS 0.006794f
C941 B.n299 VSUBS 0.006794f
C942 B.n300 VSUBS 0.006794f
C943 B.n301 VSUBS 0.006794f
C944 B.n302 VSUBS 0.006794f
C945 B.n303 VSUBS 0.006794f
C946 B.n304 VSUBS 0.006794f
C947 B.n305 VSUBS 0.006794f
C948 B.n306 VSUBS 0.006794f
C949 B.n307 VSUBS 0.006794f
C950 B.n308 VSUBS 0.006794f
C951 B.n309 VSUBS 0.006794f
C952 B.n310 VSUBS 0.006794f
C953 B.n311 VSUBS 0.006794f
C954 B.n312 VSUBS 0.006794f
C955 B.n313 VSUBS 0.006794f
C956 B.n314 VSUBS 0.006794f
C957 B.n315 VSUBS 0.006794f
C958 B.n316 VSUBS 0.006794f
C959 B.n317 VSUBS 0.006794f
C960 B.n318 VSUBS 0.006794f
C961 B.n319 VSUBS 0.006794f
C962 B.n320 VSUBS 0.006794f
C963 B.n321 VSUBS 0.015317f
C964 B.n322 VSUBS 0.016136f
C965 B.n323 VSUBS 0.015237f
C966 B.n324 VSUBS 0.006794f
C967 B.n325 VSUBS 0.006794f
C968 B.n326 VSUBS 0.006794f
C969 B.n327 VSUBS 0.006794f
C970 B.n328 VSUBS 0.006794f
C971 B.n329 VSUBS 0.006794f
C972 B.n330 VSUBS 0.006794f
C973 B.n331 VSUBS 0.006794f
C974 B.n332 VSUBS 0.006794f
C975 B.n333 VSUBS 0.006794f
C976 B.n334 VSUBS 0.006794f
C977 B.n335 VSUBS 0.006794f
C978 B.n336 VSUBS 0.006794f
C979 B.n337 VSUBS 0.006794f
C980 B.n338 VSUBS 0.006794f
C981 B.n339 VSUBS 0.006794f
C982 B.n340 VSUBS 0.006794f
C983 B.n341 VSUBS 0.006794f
C984 B.n342 VSUBS 0.006794f
C985 B.n343 VSUBS 0.006794f
C986 B.n344 VSUBS 0.006794f
C987 B.n345 VSUBS 0.006794f
C988 B.n346 VSUBS 0.006794f
C989 B.n347 VSUBS 0.006794f
C990 B.n348 VSUBS 0.006794f
C991 B.n349 VSUBS 0.006794f
C992 B.n350 VSUBS 0.006794f
C993 B.n351 VSUBS 0.006794f
C994 B.n352 VSUBS 0.006794f
C995 B.n353 VSUBS 0.006794f
C996 B.n354 VSUBS 0.006794f
C997 B.n355 VSUBS 0.006794f
C998 B.n356 VSUBS 0.006794f
C999 B.n357 VSUBS 0.006794f
C1000 B.n358 VSUBS 0.006794f
C1001 B.n359 VSUBS 0.006794f
C1002 B.n360 VSUBS 0.006794f
C1003 B.n361 VSUBS 0.006794f
C1004 B.n362 VSUBS 0.006794f
C1005 B.n363 VSUBS 0.006794f
C1006 B.n364 VSUBS 0.006794f
C1007 B.n365 VSUBS 0.006794f
C1008 B.n366 VSUBS 0.006794f
C1009 B.n367 VSUBS 0.006794f
C1010 B.n368 VSUBS 0.006794f
C1011 B.n369 VSUBS 0.006794f
C1012 B.n370 VSUBS 0.006794f
C1013 B.n371 VSUBS 0.006794f
C1014 B.n372 VSUBS 0.015237f
C1015 B.n373 VSUBS 0.015237f
C1016 B.n374 VSUBS 0.016136f
C1017 B.n375 VSUBS 0.006794f
C1018 B.n376 VSUBS 0.006794f
C1019 B.n377 VSUBS 0.006794f
C1020 B.n378 VSUBS 0.006794f
C1021 B.n379 VSUBS 0.006794f
C1022 B.n380 VSUBS 0.006794f
C1023 B.n381 VSUBS 0.006794f
C1024 B.n382 VSUBS 0.006794f
C1025 B.n383 VSUBS 0.006794f
C1026 B.n384 VSUBS 0.006794f
C1027 B.n385 VSUBS 0.006794f
C1028 B.n386 VSUBS 0.006794f
C1029 B.n387 VSUBS 0.006794f
C1030 B.n388 VSUBS 0.006794f
C1031 B.n389 VSUBS 0.006794f
C1032 B.n390 VSUBS 0.006794f
C1033 B.n391 VSUBS 0.006794f
C1034 B.n392 VSUBS 0.006794f
C1035 B.n393 VSUBS 0.006794f
C1036 B.n394 VSUBS 0.006794f
C1037 B.n395 VSUBS 0.006794f
C1038 B.n396 VSUBS 0.006794f
C1039 B.n397 VSUBS 0.006794f
C1040 B.n398 VSUBS 0.006794f
C1041 B.n399 VSUBS 0.006794f
C1042 B.n400 VSUBS 0.006794f
C1043 B.n401 VSUBS 0.006794f
C1044 B.n402 VSUBS 0.006794f
C1045 B.n403 VSUBS 0.006794f
C1046 B.n404 VSUBS 0.006794f
C1047 B.n405 VSUBS 0.006794f
C1048 B.n406 VSUBS 0.006794f
C1049 B.n407 VSUBS 0.006794f
C1050 B.n408 VSUBS 0.006794f
C1051 B.n409 VSUBS 0.006794f
C1052 B.n410 VSUBS 0.006794f
C1053 B.n411 VSUBS 0.006794f
C1054 B.n412 VSUBS 0.006794f
C1055 B.n413 VSUBS 0.006794f
C1056 B.n414 VSUBS 0.006794f
C1057 B.n415 VSUBS 0.006794f
C1058 B.n416 VSUBS 0.006794f
C1059 B.n417 VSUBS 0.006794f
C1060 B.n418 VSUBS 0.006794f
C1061 B.n419 VSUBS 0.006794f
C1062 B.n420 VSUBS 0.006794f
C1063 B.n421 VSUBS 0.006794f
C1064 B.n422 VSUBS 0.006794f
C1065 B.n423 VSUBS 0.006794f
C1066 B.n424 VSUBS 0.006794f
C1067 B.n425 VSUBS 0.006794f
C1068 B.n426 VSUBS 0.006794f
C1069 B.n427 VSUBS 0.006794f
C1070 B.n428 VSUBS 0.006794f
C1071 B.n429 VSUBS 0.006794f
C1072 B.n430 VSUBS 0.006794f
C1073 B.n431 VSUBS 0.006794f
C1074 B.n432 VSUBS 0.006794f
C1075 B.n433 VSUBS 0.006794f
C1076 B.n434 VSUBS 0.006794f
C1077 B.n435 VSUBS 0.006794f
C1078 B.n436 VSUBS 0.006794f
C1079 B.n437 VSUBS 0.006794f
C1080 B.n438 VSUBS 0.006794f
C1081 B.n439 VSUBS 0.006794f
C1082 B.n440 VSUBS 0.006794f
C1083 B.n441 VSUBS 0.006195f
C1084 B.n442 VSUBS 0.006794f
C1085 B.n443 VSUBS 0.006794f
C1086 B.n444 VSUBS 0.003997f
C1087 B.n445 VSUBS 0.006794f
C1088 B.n446 VSUBS 0.006794f
C1089 B.n447 VSUBS 0.006794f
C1090 B.n448 VSUBS 0.006794f
C1091 B.n449 VSUBS 0.006794f
C1092 B.n450 VSUBS 0.006794f
C1093 B.n451 VSUBS 0.006794f
C1094 B.n452 VSUBS 0.006794f
C1095 B.n453 VSUBS 0.006794f
C1096 B.n454 VSUBS 0.006794f
C1097 B.n455 VSUBS 0.006794f
C1098 B.n456 VSUBS 0.006794f
C1099 B.n457 VSUBS 0.003997f
C1100 B.n458 VSUBS 0.015741f
C1101 B.n459 VSUBS 0.006195f
C1102 B.n460 VSUBS 0.006794f
C1103 B.n461 VSUBS 0.006794f
C1104 B.n462 VSUBS 0.006794f
C1105 B.n463 VSUBS 0.006794f
C1106 B.n464 VSUBS 0.006794f
C1107 B.n465 VSUBS 0.006794f
C1108 B.n466 VSUBS 0.006794f
C1109 B.n467 VSUBS 0.006794f
C1110 B.n468 VSUBS 0.006794f
C1111 B.n469 VSUBS 0.006794f
C1112 B.n470 VSUBS 0.006794f
C1113 B.n471 VSUBS 0.006794f
C1114 B.n472 VSUBS 0.006794f
C1115 B.n473 VSUBS 0.006794f
C1116 B.n474 VSUBS 0.006794f
C1117 B.n475 VSUBS 0.006794f
C1118 B.n476 VSUBS 0.006794f
C1119 B.n477 VSUBS 0.006794f
C1120 B.n478 VSUBS 0.006794f
C1121 B.n479 VSUBS 0.006794f
C1122 B.n480 VSUBS 0.006794f
C1123 B.n481 VSUBS 0.006794f
C1124 B.n482 VSUBS 0.006794f
C1125 B.n483 VSUBS 0.006794f
C1126 B.n484 VSUBS 0.006794f
C1127 B.n485 VSUBS 0.006794f
C1128 B.n486 VSUBS 0.006794f
C1129 B.n487 VSUBS 0.006794f
C1130 B.n488 VSUBS 0.006794f
C1131 B.n489 VSUBS 0.006794f
C1132 B.n490 VSUBS 0.006794f
C1133 B.n491 VSUBS 0.006794f
C1134 B.n492 VSUBS 0.006794f
C1135 B.n493 VSUBS 0.006794f
C1136 B.n494 VSUBS 0.006794f
C1137 B.n495 VSUBS 0.006794f
C1138 B.n496 VSUBS 0.006794f
C1139 B.n497 VSUBS 0.006794f
C1140 B.n498 VSUBS 0.006794f
C1141 B.n499 VSUBS 0.006794f
C1142 B.n500 VSUBS 0.006794f
C1143 B.n501 VSUBS 0.006794f
C1144 B.n502 VSUBS 0.006794f
C1145 B.n503 VSUBS 0.006794f
C1146 B.n504 VSUBS 0.006794f
C1147 B.n505 VSUBS 0.006794f
C1148 B.n506 VSUBS 0.006794f
C1149 B.n507 VSUBS 0.006794f
C1150 B.n508 VSUBS 0.006794f
C1151 B.n509 VSUBS 0.006794f
C1152 B.n510 VSUBS 0.006794f
C1153 B.n511 VSUBS 0.006794f
C1154 B.n512 VSUBS 0.006794f
C1155 B.n513 VSUBS 0.006794f
C1156 B.n514 VSUBS 0.006794f
C1157 B.n515 VSUBS 0.006794f
C1158 B.n516 VSUBS 0.006794f
C1159 B.n517 VSUBS 0.006794f
C1160 B.n518 VSUBS 0.006794f
C1161 B.n519 VSUBS 0.006794f
C1162 B.n520 VSUBS 0.006794f
C1163 B.n521 VSUBS 0.006794f
C1164 B.n522 VSUBS 0.006794f
C1165 B.n523 VSUBS 0.006794f
C1166 B.n524 VSUBS 0.006794f
C1167 B.n525 VSUBS 0.006794f
C1168 B.n526 VSUBS 0.006794f
C1169 B.n527 VSUBS 0.016136f
C1170 B.n528 VSUBS 0.015237f
C1171 B.n529 VSUBS 0.015237f
C1172 B.n530 VSUBS 0.006794f
C1173 B.n531 VSUBS 0.006794f
C1174 B.n532 VSUBS 0.006794f
C1175 B.n533 VSUBS 0.006794f
C1176 B.n534 VSUBS 0.006794f
C1177 B.n535 VSUBS 0.006794f
C1178 B.n536 VSUBS 0.006794f
C1179 B.n537 VSUBS 0.006794f
C1180 B.n538 VSUBS 0.006794f
C1181 B.n539 VSUBS 0.006794f
C1182 B.n540 VSUBS 0.006794f
C1183 B.n541 VSUBS 0.006794f
C1184 B.n542 VSUBS 0.006794f
C1185 B.n543 VSUBS 0.006794f
C1186 B.n544 VSUBS 0.006794f
C1187 B.n545 VSUBS 0.006794f
C1188 B.n546 VSUBS 0.006794f
C1189 B.n547 VSUBS 0.006794f
C1190 B.n548 VSUBS 0.006794f
C1191 B.n549 VSUBS 0.006794f
C1192 B.n550 VSUBS 0.006794f
C1193 B.n551 VSUBS 0.008866f
C1194 B.n552 VSUBS 0.009444f
C1195 B.n553 VSUBS 0.018781f
.ends

