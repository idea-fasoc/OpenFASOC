* NGSPICE file created from diff_pair_sample_0335.ext - technology: sky130A

.subckt diff_pair_sample_0335 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t10 VP.t0 VDD1.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=2.9964 pd=18.49 as=2.9964 ps=18.49 w=18.16 l=1.44
X1 B.t19 B.t17 B.t18 B.t14 sky130_fd_pr__nfet_01v8 ad=7.0824 pd=37.1 as=0 ps=0 w=18.16 l=1.44
X2 VTAIL.t9 VP.t1 VDD1.t5 B.t4 sky130_fd_pr__nfet_01v8 ad=2.9964 pd=18.49 as=2.9964 ps=18.49 w=18.16 l=1.44
X3 VTAIL.t4 VN.t0 VDD2.t5 B.t4 sky130_fd_pr__nfet_01v8 ad=2.9964 pd=18.49 as=2.9964 ps=18.49 w=18.16 l=1.44
X4 B.t16 B.t13 B.t15 B.t14 sky130_fd_pr__nfet_01v8 ad=7.0824 pd=37.1 as=0 ps=0 w=18.16 l=1.44
X5 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=7.0824 pd=37.1 as=0 ps=0 w=18.16 l=1.44
X6 VDD1.t4 VP.t2 VTAIL.t8 B.t1 sky130_fd_pr__nfet_01v8 ad=7.0824 pd=37.1 as=2.9964 ps=18.49 w=18.16 l=1.44
X7 VDD1.t1 VP.t3 VTAIL.t7 B.t2 sky130_fd_pr__nfet_01v8 ad=7.0824 pd=37.1 as=2.9964 ps=18.49 w=18.16 l=1.44
X8 VDD2.t4 VN.t1 VTAIL.t11 B.t5 sky130_fd_pr__nfet_01v8 ad=2.9964 pd=18.49 as=7.0824 ps=37.1 w=18.16 l=1.44
X9 VDD2.t3 VN.t2 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.9964 pd=18.49 as=7.0824 ps=37.1 w=18.16 l=1.44
X10 VDD1.t0 VP.t4 VTAIL.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=2.9964 pd=18.49 as=7.0824 ps=37.1 w=18.16 l=1.44
X11 VDD1.t3 VP.t5 VTAIL.t5 B.t3 sky130_fd_pr__nfet_01v8 ad=2.9964 pd=18.49 as=7.0824 ps=37.1 w=18.16 l=1.44
X12 VDD2.t2 VN.t3 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=7.0824 pd=37.1 as=2.9964 ps=18.49 w=18.16 l=1.44
X13 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=7.0824 pd=37.1 as=0 ps=0 w=18.16 l=1.44
X14 VDD2.t1 VN.t4 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=7.0824 pd=37.1 as=2.9964 ps=18.49 w=18.16 l=1.44
X15 VTAIL.t0 VN.t5 VDD2.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.9964 pd=18.49 as=2.9964 ps=18.49 w=18.16 l=1.44
R0 VP.n7 VP.t3 340.046
R1 VP.n20 VP.t1 303.928
R2 VP.n14 VP.t2 303.928
R3 VP.n26 VP.t5 303.928
R4 VP.n6 VP.t0 303.928
R5 VP.n12 VP.t4 303.928
R6 VP.n15 VP.n14 172.613
R7 VP.n27 VP.n26 172.613
R8 VP.n13 VP.n12 172.613
R9 VP.n8 VP.n5 161.3
R10 VP.n10 VP.n9 161.3
R11 VP.n11 VP.n4 161.3
R12 VP.n25 VP.n0 161.3
R13 VP.n24 VP.n23 161.3
R14 VP.n22 VP.n1 161.3
R15 VP.n21 VP.n20 161.3
R16 VP.n19 VP.n2 161.3
R17 VP.n18 VP.n17 161.3
R18 VP.n16 VP.n3 161.3
R19 VP.n19 VP.n18 51.7179
R20 VP.n24 VP.n1 51.7179
R21 VP.n10 VP.n5 51.7179
R22 VP.n15 VP.n13 48.7543
R23 VP.n7 VP.n6 41.9337
R24 VP.n18 VP.n3 29.4362
R25 VP.n25 VP.n24 29.4362
R26 VP.n11 VP.n10 29.4362
R27 VP.n20 VP.n19 24.5923
R28 VP.n20 VP.n1 24.5923
R29 VP.n6 VP.n5 24.5923
R30 VP.n8 VP.n7 17.4039
R31 VP.n14 VP.n3 13.2801
R32 VP.n26 VP.n25 13.2801
R33 VP.n12 VP.n11 13.2801
R34 VP.n9 VP.n8 0.189894
R35 VP.n9 VP.n4 0.189894
R36 VP.n13 VP.n4 0.189894
R37 VP.n16 VP.n15 0.189894
R38 VP.n17 VP.n16 0.189894
R39 VP.n17 VP.n2 0.189894
R40 VP.n21 VP.n2 0.189894
R41 VP.n22 VP.n21 0.189894
R42 VP.n23 VP.n22 0.189894
R43 VP.n23 VP.n0 0.189894
R44 VP.n27 VP.n0 0.189894
R45 VP VP.n27 0.0516364
R46 VDD1.n96 VDD1.n0 289.615
R47 VDD1.n197 VDD1.n101 289.615
R48 VDD1.n97 VDD1.n96 185
R49 VDD1.n95 VDD1.n94 185
R50 VDD1.n4 VDD1.n3 185
R51 VDD1.n89 VDD1.n88 185
R52 VDD1.n87 VDD1.n86 185
R53 VDD1.n8 VDD1.n7 185
R54 VDD1.n81 VDD1.n80 185
R55 VDD1.n79 VDD1.n10 185
R56 VDD1.n78 VDD1.n77 185
R57 VDD1.n13 VDD1.n11 185
R58 VDD1.n72 VDD1.n71 185
R59 VDD1.n70 VDD1.n69 185
R60 VDD1.n17 VDD1.n16 185
R61 VDD1.n64 VDD1.n63 185
R62 VDD1.n62 VDD1.n61 185
R63 VDD1.n21 VDD1.n20 185
R64 VDD1.n56 VDD1.n55 185
R65 VDD1.n54 VDD1.n53 185
R66 VDD1.n25 VDD1.n24 185
R67 VDD1.n48 VDD1.n47 185
R68 VDD1.n46 VDD1.n45 185
R69 VDD1.n29 VDD1.n28 185
R70 VDD1.n40 VDD1.n39 185
R71 VDD1.n38 VDD1.n37 185
R72 VDD1.n33 VDD1.n32 185
R73 VDD1.n133 VDD1.n132 185
R74 VDD1.n138 VDD1.n137 185
R75 VDD1.n140 VDD1.n139 185
R76 VDD1.n129 VDD1.n128 185
R77 VDD1.n146 VDD1.n145 185
R78 VDD1.n148 VDD1.n147 185
R79 VDD1.n125 VDD1.n124 185
R80 VDD1.n154 VDD1.n153 185
R81 VDD1.n156 VDD1.n155 185
R82 VDD1.n121 VDD1.n120 185
R83 VDD1.n162 VDD1.n161 185
R84 VDD1.n164 VDD1.n163 185
R85 VDD1.n117 VDD1.n116 185
R86 VDD1.n170 VDD1.n169 185
R87 VDD1.n172 VDD1.n171 185
R88 VDD1.n113 VDD1.n112 185
R89 VDD1.n179 VDD1.n178 185
R90 VDD1.n180 VDD1.n111 185
R91 VDD1.n182 VDD1.n181 185
R92 VDD1.n109 VDD1.n108 185
R93 VDD1.n188 VDD1.n187 185
R94 VDD1.n190 VDD1.n189 185
R95 VDD1.n105 VDD1.n104 185
R96 VDD1.n196 VDD1.n195 185
R97 VDD1.n198 VDD1.n197 185
R98 VDD1.n34 VDD1.t1 147.659
R99 VDD1.n134 VDD1.t4 147.659
R100 VDD1.n96 VDD1.n95 104.615
R101 VDD1.n95 VDD1.n3 104.615
R102 VDD1.n88 VDD1.n3 104.615
R103 VDD1.n88 VDD1.n87 104.615
R104 VDD1.n87 VDD1.n7 104.615
R105 VDD1.n80 VDD1.n7 104.615
R106 VDD1.n80 VDD1.n79 104.615
R107 VDD1.n79 VDD1.n78 104.615
R108 VDD1.n78 VDD1.n11 104.615
R109 VDD1.n71 VDD1.n11 104.615
R110 VDD1.n71 VDD1.n70 104.615
R111 VDD1.n70 VDD1.n16 104.615
R112 VDD1.n63 VDD1.n16 104.615
R113 VDD1.n63 VDD1.n62 104.615
R114 VDD1.n62 VDD1.n20 104.615
R115 VDD1.n55 VDD1.n20 104.615
R116 VDD1.n55 VDD1.n54 104.615
R117 VDD1.n54 VDD1.n24 104.615
R118 VDD1.n47 VDD1.n24 104.615
R119 VDD1.n47 VDD1.n46 104.615
R120 VDD1.n46 VDD1.n28 104.615
R121 VDD1.n39 VDD1.n28 104.615
R122 VDD1.n39 VDD1.n38 104.615
R123 VDD1.n38 VDD1.n32 104.615
R124 VDD1.n138 VDD1.n132 104.615
R125 VDD1.n139 VDD1.n138 104.615
R126 VDD1.n139 VDD1.n128 104.615
R127 VDD1.n146 VDD1.n128 104.615
R128 VDD1.n147 VDD1.n146 104.615
R129 VDD1.n147 VDD1.n124 104.615
R130 VDD1.n154 VDD1.n124 104.615
R131 VDD1.n155 VDD1.n154 104.615
R132 VDD1.n155 VDD1.n120 104.615
R133 VDD1.n162 VDD1.n120 104.615
R134 VDD1.n163 VDD1.n162 104.615
R135 VDD1.n163 VDD1.n116 104.615
R136 VDD1.n170 VDD1.n116 104.615
R137 VDD1.n171 VDD1.n170 104.615
R138 VDD1.n171 VDD1.n112 104.615
R139 VDD1.n179 VDD1.n112 104.615
R140 VDD1.n180 VDD1.n179 104.615
R141 VDD1.n181 VDD1.n180 104.615
R142 VDD1.n181 VDD1.n108 104.615
R143 VDD1.n188 VDD1.n108 104.615
R144 VDD1.n189 VDD1.n188 104.615
R145 VDD1.n189 VDD1.n104 104.615
R146 VDD1.n196 VDD1.n104 104.615
R147 VDD1.n197 VDD1.n196 104.615
R148 VDD1.n203 VDD1.n202 59.4227
R149 VDD1.n205 VDD1.n204 59.0966
R150 VDD1.t1 VDD1.n32 52.3082
R151 VDD1.t4 VDD1.n132 52.3082
R152 VDD1 VDD1.n100 48.5152
R153 VDD1.n203 VDD1.n201 48.4017
R154 VDD1.n205 VDD1.n203 45.6755
R155 VDD1.n34 VDD1.n33 15.6677
R156 VDD1.n134 VDD1.n133 15.6677
R157 VDD1.n81 VDD1.n10 13.1884
R158 VDD1.n182 VDD1.n111 13.1884
R159 VDD1.n82 VDD1.n8 12.8005
R160 VDD1.n77 VDD1.n12 12.8005
R161 VDD1.n37 VDD1.n36 12.8005
R162 VDD1.n137 VDD1.n136 12.8005
R163 VDD1.n178 VDD1.n177 12.8005
R164 VDD1.n183 VDD1.n109 12.8005
R165 VDD1.n86 VDD1.n85 12.0247
R166 VDD1.n76 VDD1.n13 12.0247
R167 VDD1.n40 VDD1.n31 12.0247
R168 VDD1.n140 VDD1.n131 12.0247
R169 VDD1.n176 VDD1.n113 12.0247
R170 VDD1.n187 VDD1.n186 12.0247
R171 VDD1.n89 VDD1.n6 11.249
R172 VDD1.n73 VDD1.n72 11.249
R173 VDD1.n41 VDD1.n29 11.249
R174 VDD1.n141 VDD1.n129 11.249
R175 VDD1.n173 VDD1.n172 11.249
R176 VDD1.n190 VDD1.n107 11.249
R177 VDD1.n90 VDD1.n4 10.4732
R178 VDD1.n69 VDD1.n15 10.4732
R179 VDD1.n45 VDD1.n44 10.4732
R180 VDD1.n145 VDD1.n144 10.4732
R181 VDD1.n169 VDD1.n115 10.4732
R182 VDD1.n191 VDD1.n105 10.4732
R183 VDD1.n94 VDD1.n93 9.69747
R184 VDD1.n68 VDD1.n17 9.69747
R185 VDD1.n48 VDD1.n27 9.69747
R186 VDD1.n148 VDD1.n127 9.69747
R187 VDD1.n168 VDD1.n117 9.69747
R188 VDD1.n195 VDD1.n194 9.69747
R189 VDD1.n100 VDD1.n99 9.45567
R190 VDD1.n201 VDD1.n200 9.45567
R191 VDD1.n60 VDD1.n59 9.3005
R192 VDD1.n19 VDD1.n18 9.3005
R193 VDD1.n66 VDD1.n65 9.3005
R194 VDD1.n68 VDD1.n67 9.3005
R195 VDD1.n15 VDD1.n14 9.3005
R196 VDD1.n74 VDD1.n73 9.3005
R197 VDD1.n76 VDD1.n75 9.3005
R198 VDD1.n12 VDD1.n9 9.3005
R199 VDD1.n99 VDD1.n98 9.3005
R200 VDD1.n2 VDD1.n1 9.3005
R201 VDD1.n93 VDD1.n92 9.3005
R202 VDD1.n91 VDD1.n90 9.3005
R203 VDD1.n6 VDD1.n5 9.3005
R204 VDD1.n85 VDD1.n84 9.3005
R205 VDD1.n83 VDD1.n82 9.3005
R206 VDD1.n58 VDD1.n57 9.3005
R207 VDD1.n23 VDD1.n22 9.3005
R208 VDD1.n52 VDD1.n51 9.3005
R209 VDD1.n50 VDD1.n49 9.3005
R210 VDD1.n27 VDD1.n26 9.3005
R211 VDD1.n44 VDD1.n43 9.3005
R212 VDD1.n42 VDD1.n41 9.3005
R213 VDD1.n31 VDD1.n30 9.3005
R214 VDD1.n36 VDD1.n35 9.3005
R215 VDD1.n200 VDD1.n199 9.3005
R216 VDD1.n103 VDD1.n102 9.3005
R217 VDD1.n194 VDD1.n193 9.3005
R218 VDD1.n192 VDD1.n191 9.3005
R219 VDD1.n107 VDD1.n106 9.3005
R220 VDD1.n186 VDD1.n185 9.3005
R221 VDD1.n184 VDD1.n183 9.3005
R222 VDD1.n123 VDD1.n122 9.3005
R223 VDD1.n152 VDD1.n151 9.3005
R224 VDD1.n150 VDD1.n149 9.3005
R225 VDD1.n127 VDD1.n126 9.3005
R226 VDD1.n144 VDD1.n143 9.3005
R227 VDD1.n142 VDD1.n141 9.3005
R228 VDD1.n131 VDD1.n130 9.3005
R229 VDD1.n136 VDD1.n135 9.3005
R230 VDD1.n158 VDD1.n157 9.3005
R231 VDD1.n160 VDD1.n159 9.3005
R232 VDD1.n119 VDD1.n118 9.3005
R233 VDD1.n166 VDD1.n165 9.3005
R234 VDD1.n168 VDD1.n167 9.3005
R235 VDD1.n115 VDD1.n114 9.3005
R236 VDD1.n174 VDD1.n173 9.3005
R237 VDD1.n176 VDD1.n175 9.3005
R238 VDD1.n177 VDD1.n110 9.3005
R239 VDD1.n97 VDD1.n2 8.92171
R240 VDD1.n65 VDD1.n64 8.92171
R241 VDD1.n49 VDD1.n25 8.92171
R242 VDD1.n149 VDD1.n125 8.92171
R243 VDD1.n165 VDD1.n164 8.92171
R244 VDD1.n198 VDD1.n103 8.92171
R245 VDD1.n98 VDD1.n0 8.14595
R246 VDD1.n61 VDD1.n19 8.14595
R247 VDD1.n53 VDD1.n52 8.14595
R248 VDD1.n153 VDD1.n152 8.14595
R249 VDD1.n161 VDD1.n119 8.14595
R250 VDD1.n199 VDD1.n101 8.14595
R251 VDD1.n60 VDD1.n21 7.3702
R252 VDD1.n56 VDD1.n23 7.3702
R253 VDD1.n156 VDD1.n123 7.3702
R254 VDD1.n160 VDD1.n121 7.3702
R255 VDD1.n57 VDD1.n21 6.59444
R256 VDD1.n57 VDD1.n56 6.59444
R257 VDD1.n157 VDD1.n156 6.59444
R258 VDD1.n157 VDD1.n121 6.59444
R259 VDD1.n100 VDD1.n0 5.81868
R260 VDD1.n61 VDD1.n60 5.81868
R261 VDD1.n53 VDD1.n23 5.81868
R262 VDD1.n153 VDD1.n123 5.81868
R263 VDD1.n161 VDD1.n160 5.81868
R264 VDD1.n201 VDD1.n101 5.81868
R265 VDD1.n98 VDD1.n97 5.04292
R266 VDD1.n64 VDD1.n19 5.04292
R267 VDD1.n52 VDD1.n25 5.04292
R268 VDD1.n152 VDD1.n125 5.04292
R269 VDD1.n164 VDD1.n119 5.04292
R270 VDD1.n199 VDD1.n198 5.04292
R271 VDD1.n35 VDD1.n34 4.38563
R272 VDD1.n135 VDD1.n134 4.38563
R273 VDD1.n94 VDD1.n2 4.26717
R274 VDD1.n65 VDD1.n17 4.26717
R275 VDD1.n49 VDD1.n48 4.26717
R276 VDD1.n149 VDD1.n148 4.26717
R277 VDD1.n165 VDD1.n117 4.26717
R278 VDD1.n195 VDD1.n103 4.26717
R279 VDD1.n93 VDD1.n4 3.49141
R280 VDD1.n69 VDD1.n68 3.49141
R281 VDD1.n45 VDD1.n27 3.49141
R282 VDD1.n145 VDD1.n127 3.49141
R283 VDD1.n169 VDD1.n168 3.49141
R284 VDD1.n194 VDD1.n105 3.49141
R285 VDD1.n90 VDD1.n89 2.71565
R286 VDD1.n72 VDD1.n15 2.71565
R287 VDD1.n44 VDD1.n29 2.71565
R288 VDD1.n144 VDD1.n129 2.71565
R289 VDD1.n172 VDD1.n115 2.71565
R290 VDD1.n191 VDD1.n190 2.71565
R291 VDD1.n86 VDD1.n6 1.93989
R292 VDD1.n73 VDD1.n13 1.93989
R293 VDD1.n41 VDD1.n40 1.93989
R294 VDD1.n141 VDD1.n140 1.93989
R295 VDD1.n173 VDD1.n113 1.93989
R296 VDD1.n187 VDD1.n107 1.93989
R297 VDD1.n85 VDD1.n8 1.16414
R298 VDD1.n77 VDD1.n76 1.16414
R299 VDD1.n37 VDD1.n31 1.16414
R300 VDD1.n137 VDD1.n131 1.16414
R301 VDD1.n178 VDD1.n176 1.16414
R302 VDD1.n186 VDD1.n109 1.16414
R303 VDD1.n204 VDD1.t2 1.09081
R304 VDD1.n204 VDD1.t0 1.09081
R305 VDD1.n202 VDD1.t5 1.09081
R306 VDD1.n202 VDD1.t3 1.09081
R307 VDD1.n82 VDD1.n81 0.388379
R308 VDD1.n12 VDD1.n10 0.388379
R309 VDD1.n36 VDD1.n33 0.388379
R310 VDD1.n136 VDD1.n133 0.388379
R311 VDD1.n177 VDD1.n111 0.388379
R312 VDD1.n183 VDD1.n182 0.388379
R313 VDD1 VDD1.n205 0.323776
R314 VDD1.n99 VDD1.n1 0.155672
R315 VDD1.n92 VDD1.n1 0.155672
R316 VDD1.n92 VDD1.n91 0.155672
R317 VDD1.n91 VDD1.n5 0.155672
R318 VDD1.n84 VDD1.n5 0.155672
R319 VDD1.n84 VDD1.n83 0.155672
R320 VDD1.n83 VDD1.n9 0.155672
R321 VDD1.n75 VDD1.n9 0.155672
R322 VDD1.n75 VDD1.n74 0.155672
R323 VDD1.n74 VDD1.n14 0.155672
R324 VDD1.n67 VDD1.n14 0.155672
R325 VDD1.n67 VDD1.n66 0.155672
R326 VDD1.n66 VDD1.n18 0.155672
R327 VDD1.n59 VDD1.n18 0.155672
R328 VDD1.n59 VDD1.n58 0.155672
R329 VDD1.n58 VDD1.n22 0.155672
R330 VDD1.n51 VDD1.n22 0.155672
R331 VDD1.n51 VDD1.n50 0.155672
R332 VDD1.n50 VDD1.n26 0.155672
R333 VDD1.n43 VDD1.n26 0.155672
R334 VDD1.n43 VDD1.n42 0.155672
R335 VDD1.n42 VDD1.n30 0.155672
R336 VDD1.n35 VDD1.n30 0.155672
R337 VDD1.n135 VDD1.n130 0.155672
R338 VDD1.n142 VDD1.n130 0.155672
R339 VDD1.n143 VDD1.n142 0.155672
R340 VDD1.n143 VDD1.n126 0.155672
R341 VDD1.n150 VDD1.n126 0.155672
R342 VDD1.n151 VDD1.n150 0.155672
R343 VDD1.n151 VDD1.n122 0.155672
R344 VDD1.n158 VDD1.n122 0.155672
R345 VDD1.n159 VDD1.n158 0.155672
R346 VDD1.n159 VDD1.n118 0.155672
R347 VDD1.n166 VDD1.n118 0.155672
R348 VDD1.n167 VDD1.n166 0.155672
R349 VDD1.n167 VDD1.n114 0.155672
R350 VDD1.n174 VDD1.n114 0.155672
R351 VDD1.n175 VDD1.n174 0.155672
R352 VDD1.n175 VDD1.n110 0.155672
R353 VDD1.n184 VDD1.n110 0.155672
R354 VDD1.n185 VDD1.n184 0.155672
R355 VDD1.n185 VDD1.n106 0.155672
R356 VDD1.n192 VDD1.n106 0.155672
R357 VDD1.n193 VDD1.n192 0.155672
R358 VDD1.n193 VDD1.n102 0.155672
R359 VDD1.n200 VDD1.n102 0.155672
R360 VTAIL.n410 VTAIL.n314 289.615
R361 VTAIL.n98 VTAIL.n2 289.615
R362 VTAIL.n308 VTAIL.n212 289.615
R363 VTAIL.n204 VTAIL.n108 289.615
R364 VTAIL.n346 VTAIL.n345 185
R365 VTAIL.n351 VTAIL.n350 185
R366 VTAIL.n353 VTAIL.n352 185
R367 VTAIL.n342 VTAIL.n341 185
R368 VTAIL.n359 VTAIL.n358 185
R369 VTAIL.n361 VTAIL.n360 185
R370 VTAIL.n338 VTAIL.n337 185
R371 VTAIL.n367 VTAIL.n366 185
R372 VTAIL.n369 VTAIL.n368 185
R373 VTAIL.n334 VTAIL.n333 185
R374 VTAIL.n375 VTAIL.n374 185
R375 VTAIL.n377 VTAIL.n376 185
R376 VTAIL.n330 VTAIL.n329 185
R377 VTAIL.n383 VTAIL.n382 185
R378 VTAIL.n385 VTAIL.n384 185
R379 VTAIL.n326 VTAIL.n325 185
R380 VTAIL.n392 VTAIL.n391 185
R381 VTAIL.n393 VTAIL.n324 185
R382 VTAIL.n395 VTAIL.n394 185
R383 VTAIL.n322 VTAIL.n321 185
R384 VTAIL.n401 VTAIL.n400 185
R385 VTAIL.n403 VTAIL.n402 185
R386 VTAIL.n318 VTAIL.n317 185
R387 VTAIL.n409 VTAIL.n408 185
R388 VTAIL.n411 VTAIL.n410 185
R389 VTAIL.n34 VTAIL.n33 185
R390 VTAIL.n39 VTAIL.n38 185
R391 VTAIL.n41 VTAIL.n40 185
R392 VTAIL.n30 VTAIL.n29 185
R393 VTAIL.n47 VTAIL.n46 185
R394 VTAIL.n49 VTAIL.n48 185
R395 VTAIL.n26 VTAIL.n25 185
R396 VTAIL.n55 VTAIL.n54 185
R397 VTAIL.n57 VTAIL.n56 185
R398 VTAIL.n22 VTAIL.n21 185
R399 VTAIL.n63 VTAIL.n62 185
R400 VTAIL.n65 VTAIL.n64 185
R401 VTAIL.n18 VTAIL.n17 185
R402 VTAIL.n71 VTAIL.n70 185
R403 VTAIL.n73 VTAIL.n72 185
R404 VTAIL.n14 VTAIL.n13 185
R405 VTAIL.n80 VTAIL.n79 185
R406 VTAIL.n81 VTAIL.n12 185
R407 VTAIL.n83 VTAIL.n82 185
R408 VTAIL.n10 VTAIL.n9 185
R409 VTAIL.n89 VTAIL.n88 185
R410 VTAIL.n91 VTAIL.n90 185
R411 VTAIL.n6 VTAIL.n5 185
R412 VTAIL.n97 VTAIL.n96 185
R413 VTAIL.n99 VTAIL.n98 185
R414 VTAIL.n309 VTAIL.n308 185
R415 VTAIL.n307 VTAIL.n306 185
R416 VTAIL.n216 VTAIL.n215 185
R417 VTAIL.n301 VTAIL.n300 185
R418 VTAIL.n299 VTAIL.n298 185
R419 VTAIL.n220 VTAIL.n219 185
R420 VTAIL.n293 VTAIL.n292 185
R421 VTAIL.n291 VTAIL.n222 185
R422 VTAIL.n290 VTAIL.n289 185
R423 VTAIL.n225 VTAIL.n223 185
R424 VTAIL.n284 VTAIL.n283 185
R425 VTAIL.n282 VTAIL.n281 185
R426 VTAIL.n229 VTAIL.n228 185
R427 VTAIL.n276 VTAIL.n275 185
R428 VTAIL.n274 VTAIL.n273 185
R429 VTAIL.n233 VTAIL.n232 185
R430 VTAIL.n268 VTAIL.n267 185
R431 VTAIL.n266 VTAIL.n265 185
R432 VTAIL.n237 VTAIL.n236 185
R433 VTAIL.n260 VTAIL.n259 185
R434 VTAIL.n258 VTAIL.n257 185
R435 VTAIL.n241 VTAIL.n240 185
R436 VTAIL.n252 VTAIL.n251 185
R437 VTAIL.n250 VTAIL.n249 185
R438 VTAIL.n245 VTAIL.n244 185
R439 VTAIL.n205 VTAIL.n204 185
R440 VTAIL.n203 VTAIL.n202 185
R441 VTAIL.n112 VTAIL.n111 185
R442 VTAIL.n197 VTAIL.n196 185
R443 VTAIL.n195 VTAIL.n194 185
R444 VTAIL.n116 VTAIL.n115 185
R445 VTAIL.n189 VTAIL.n188 185
R446 VTAIL.n187 VTAIL.n118 185
R447 VTAIL.n186 VTAIL.n185 185
R448 VTAIL.n121 VTAIL.n119 185
R449 VTAIL.n180 VTAIL.n179 185
R450 VTAIL.n178 VTAIL.n177 185
R451 VTAIL.n125 VTAIL.n124 185
R452 VTAIL.n172 VTAIL.n171 185
R453 VTAIL.n170 VTAIL.n169 185
R454 VTAIL.n129 VTAIL.n128 185
R455 VTAIL.n164 VTAIL.n163 185
R456 VTAIL.n162 VTAIL.n161 185
R457 VTAIL.n133 VTAIL.n132 185
R458 VTAIL.n156 VTAIL.n155 185
R459 VTAIL.n154 VTAIL.n153 185
R460 VTAIL.n137 VTAIL.n136 185
R461 VTAIL.n148 VTAIL.n147 185
R462 VTAIL.n146 VTAIL.n145 185
R463 VTAIL.n141 VTAIL.n140 185
R464 VTAIL.n347 VTAIL.t11 147.659
R465 VTAIL.n35 VTAIL.t5 147.659
R466 VTAIL.n246 VTAIL.t6 147.659
R467 VTAIL.n142 VTAIL.t3 147.659
R468 VTAIL.n351 VTAIL.n345 104.615
R469 VTAIL.n352 VTAIL.n351 104.615
R470 VTAIL.n352 VTAIL.n341 104.615
R471 VTAIL.n359 VTAIL.n341 104.615
R472 VTAIL.n360 VTAIL.n359 104.615
R473 VTAIL.n360 VTAIL.n337 104.615
R474 VTAIL.n367 VTAIL.n337 104.615
R475 VTAIL.n368 VTAIL.n367 104.615
R476 VTAIL.n368 VTAIL.n333 104.615
R477 VTAIL.n375 VTAIL.n333 104.615
R478 VTAIL.n376 VTAIL.n375 104.615
R479 VTAIL.n376 VTAIL.n329 104.615
R480 VTAIL.n383 VTAIL.n329 104.615
R481 VTAIL.n384 VTAIL.n383 104.615
R482 VTAIL.n384 VTAIL.n325 104.615
R483 VTAIL.n392 VTAIL.n325 104.615
R484 VTAIL.n393 VTAIL.n392 104.615
R485 VTAIL.n394 VTAIL.n393 104.615
R486 VTAIL.n394 VTAIL.n321 104.615
R487 VTAIL.n401 VTAIL.n321 104.615
R488 VTAIL.n402 VTAIL.n401 104.615
R489 VTAIL.n402 VTAIL.n317 104.615
R490 VTAIL.n409 VTAIL.n317 104.615
R491 VTAIL.n410 VTAIL.n409 104.615
R492 VTAIL.n39 VTAIL.n33 104.615
R493 VTAIL.n40 VTAIL.n39 104.615
R494 VTAIL.n40 VTAIL.n29 104.615
R495 VTAIL.n47 VTAIL.n29 104.615
R496 VTAIL.n48 VTAIL.n47 104.615
R497 VTAIL.n48 VTAIL.n25 104.615
R498 VTAIL.n55 VTAIL.n25 104.615
R499 VTAIL.n56 VTAIL.n55 104.615
R500 VTAIL.n56 VTAIL.n21 104.615
R501 VTAIL.n63 VTAIL.n21 104.615
R502 VTAIL.n64 VTAIL.n63 104.615
R503 VTAIL.n64 VTAIL.n17 104.615
R504 VTAIL.n71 VTAIL.n17 104.615
R505 VTAIL.n72 VTAIL.n71 104.615
R506 VTAIL.n72 VTAIL.n13 104.615
R507 VTAIL.n80 VTAIL.n13 104.615
R508 VTAIL.n81 VTAIL.n80 104.615
R509 VTAIL.n82 VTAIL.n81 104.615
R510 VTAIL.n82 VTAIL.n9 104.615
R511 VTAIL.n89 VTAIL.n9 104.615
R512 VTAIL.n90 VTAIL.n89 104.615
R513 VTAIL.n90 VTAIL.n5 104.615
R514 VTAIL.n97 VTAIL.n5 104.615
R515 VTAIL.n98 VTAIL.n97 104.615
R516 VTAIL.n308 VTAIL.n307 104.615
R517 VTAIL.n307 VTAIL.n215 104.615
R518 VTAIL.n300 VTAIL.n215 104.615
R519 VTAIL.n300 VTAIL.n299 104.615
R520 VTAIL.n299 VTAIL.n219 104.615
R521 VTAIL.n292 VTAIL.n219 104.615
R522 VTAIL.n292 VTAIL.n291 104.615
R523 VTAIL.n291 VTAIL.n290 104.615
R524 VTAIL.n290 VTAIL.n223 104.615
R525 VTAIL.n283 VTAIL.n223 104.615
R526 VTAIL.n283 VTAIL.n282 104.615
R527 VTAIL.n282 VTAIL.n228 104.615
R528 VTAIL.n275 VTAIL.n228 104.615
R529 VTAIL.n275 VTAIL.n274 104.615
R530 VTAIL.n274 VTAIL.n232 104.615
R531 VTAIL.n267 VTAIL.n232 104.615
R532 VTAIL.n267 VTAIL.n266 104.615
R533 VTAIL.n266 VTAIL.n236 104.615
R534 VTAIL.n259 VTAIL.n236 104.615
R535 VTAIL.n259 VTAIL.n258 104.615
R536 VTAIL.n258 VTAIL.n240 104.615
R537 VTAIL.n251 VTAIL.n240 104.615
R538 VTAIL.n251 VTAIL.n250 104.615
R539 VTAIL.n250 VTAIL.n244 104.615
R540 VTAIL.n204 VTAIL.n203 104.615
R541 VTAIL.n203 VTAIL.n111 104.615
R542 VTAIL.n196 VTAIL.n111 104.615
R543 VTAIL.n196 VTAIL.n195 104.615
R544 VTAIL.n195 VTAIL.n115 104.615
R545 VTAIL.n188 VTAIL.n115 104.615
R546 VTAIL.n188 VTAIL.n187 104.615
R547 VTAIL.n187 VTAIL.n186 104.615
R548 VTAIL.n186 VTAIL.n119 104.615
R549 VTAIL.n179 VTAIL.n119 104.615
R550 VTAIL.n179 VTAIL.n178 104.615
R551 VTAIL.n178 VTAIL.n124 104.615
R552 VTAIL.n171 VTAIL.n124 104.615
R553 VTAIL.n171 VTAIL.n170 104.615
R554 VTAIL.n170 VTAIL.n128 104.615
R555 VTAIL.n163 VTAIL.n128 104.615
R556 VTAIL.n163 VTAIL.n162 104.615
R557 VTAIL.n162 VTAIL.n132 104.615
R558 VTAIL.n155 VTAIL.n132 104.615
R559 VTAIL.n155 VTAIL.n154 104.615
R560 VTAIL.n154 VTAIL.n136 104.615
R561 VTAIL.n147 VTAIL.n136 104.615
R562 VTAIL.n147 VTAIL.n146 104.615
R563 VTAIL.n146 VTAIL.n140 104.615
R564 VTAIL.t11 VTAIL.n345 52.3082
R565 VTAIL.t5 VTAIL.n33 52.3082
R566 VTAIL.t6 VTAIL.n244 52.3082
R567 VTAIL.t3 VTAIL.n140 52.3082
R568 VTAIL.n211 VTAIL.n210 42.418
R569 VTAIL.n107 VTAIL.n106 42.418
R570 VTAIL.n1 VTAIL.n0 42.4178
R571 VTAIL.n105 VTAIL.n104 42.4178
R572 VTAIL.n107 VTAIL.n105 31.0738
R573 VTAIL.n415 VTAIL.n414 30.6338
R574 VTAIL.n103 VTAIL.n102 30.6338
R575 VTAIL.n313 VTAIL.n312 30.6338
R576 VTAIL.n209 VTAIL.n208 30.6338
R577 VTAIL.n415 VTAIL.n313 29.5479
R578 VTAIL.n347 VTAIL.n346 15.6677
R579 VTAIL.n35 VTAIL.n34 15.6677
R580 VTAIL.n246 VTAIL.n245 15.6677
R581 VTAIL.n142 VTAIL.n141 15.6677
R582 VTAIL.n395 VTAIL.n324 13.1884
R583 VTAIL.n83 VTAIL.n12 13.1884
R584 VTAIL.n293 VTAIL.n222 13.1884
R585 VTAIL.n189 VTAIL.n118 13.1884
R586 VTAIL.n350 VTAIL.n349 12.8005
R587 VTAIL.n391 VTAIL.n390 12.8005
R588 VTAIL.n396 VTAIL.n322 12.8005
R589 VTAIL.n38 VTAIL.n37 12.8005
R590 VTAIL.n79 VTAIL.n78 12.8005
R591 VTAIL.n84 VTAIL.n10 12.8005
R592 VTAIL.n294 VTAIL.n220 12.8005
R593 VTAIL.n289 VTAIL.n224 12.8005
R594 VTAIL.n249 VTAIL.n248 12.8005
R595 VTAIL.n190 VTAIL.n116 12.8005
R596 VTAIL.n185 VTAIL.n120 12.8005
R597 VTAIL.n145 VTAIL.n144 12.8005
R598 VTAIL.n353 VTAIL.n344 12.0247
R599 VTAIL.n389 VTAIL.n326 12.0247
R600 VTAIL.n400 VTAIL.n399 12.0247
R601 VTAIL.n41 VTAIL.n32 12.0247
R602 VTAIL.n77 VTAIL.n14 12.0247
R603 VTAIL.n88 VTAIL.n87 12.0247
R604 VTAIL.n298 VTAIL.n297 12.0247
R605 VTAIL.n288 VTAIL.n225 12.0247
R606 VTAIL.n252 VTAIL.n243 12.0247
R607 VTAIL.n194 VTAIL.n193 12.0247
R608 VTAIL.n184 VTAIL.n121 12.0247
R609 VTAIL.n148 VTAIL.n139 12.0247
R610 VTAIL.n354 VTAIL.n342 11.249
R611 VTAIL.n386 VTAIL.n385 11.249
R612 VTAIL.n403 VTAIL.n320 11.249
R613 VTAIL.n42 VTAIL.n30 11.249
R614 VTAIL.n74 VTAIL.n73 11.249
R615 VTAIL.n91 VTAIL.n8 11.249
R616 VTAIL.n301 VTAIL.n218 11.249
R617 VTAIL.n285 VTAIL.n284 11.249
R618 VTAIL.n253 VTAIL.n241 11.249
R619 VTAIL.n197 VTAIL.n114 11.249
R620 VTAIL.n181 VTAIL.n180 11.249
R621 VTAIL.n149 VTAIL.n137 11.249
R622 VTAIL.n358 VTAIL.n357 10.4732
R623 VTAIL.n382 VTAIL.n328 10.4732
R624 VTAIL.n404 VTAIL.n318 10.4732
R625 VTAIL.n46 VTAIL.n45 10.4732
R626 VTAIL.n70 VTAIL.n16 10.4732
R627 VTAIL.n92 VTAIL.n6 10.4732
R628 VTAIL.n302 VTAIL.n216 10.4732
R629 VTAIL.n281 VTAIL.n227 10.4732
R630 VTAIL.n257 VTAIL.n256 10.4732
R631 VTAIL.n198 VTAIL.n112 10.4732
R632 VTAIL.n177 VTAIL.n123 10.4732
R633 VTAIL.n153 VTAIL.n152 10.4732
R634 VTAIL.n361 VTAIL.n340 9.69747
R635 VTAIL.n381 VTAIL.n330 9.69747
R636 VTAIL.n408 VTAIL.n407 9.69747
R637 VTAIL.n49 VTAIL.n28 9.69747
R638 VTAIL.n69 VTAIL.n18 9.69747
R639 VTAIL.n96 VTAIL.n95 9.69747
R640 VTAIL.n306 VTAIL.n305 9.69747
R641 VTAIL.n280 VTAIL.n229 9.69747
R642 VTAIL.n260 VTAIL.n239 9.69747
R643 VTAIL.n202 VTAIL.n201 9.69747
R644 VTAIL.n176 VTAIL.n125 9.69747
R645 VTAIL.n156 VTAIL.n135 9.69747
R646 VTAIL.n414 VTAIL.n413 9.45567
R647 VTAIL.n102 VTAIL.n101 9.45567
R648 VTAIL.n312 VTAIL.n311 9.45567
R649 VTAIL.n208 VTAIL.n207 9.45567
R650 VTAIL.n413 VTAIL.n412 9.3005
R651 VTAIL.n316 VTAIL.n315 9.3005
R652 VTAIL.n407 VTAIL.n406 9.3005
R653 VTAIL.n405 VTAIL.n404 9.3005
R654 VTAIL.n320 VTAIL.n319 9.3005
R655 VTAIL.n399 VTAIL.n398 9.3005
R656 VTAIL.n397 VTAIL.n396 9.3005
R657 VTAIL.n336 VTAIL.n335 9.3005
R658 VTAIL.n365 VTAIL.n364 9.3005
R659 VTAIL.n363 VTAIL.n362 9.3005
R660 VTAIL.n340 VTAIL.n339 9.3005
R661 VTAIL.n357 VTAIL.n356 9.3005
R662 VTAIL.n355 VTAIL.n354 9.3005
R663 VTAIL.n344 VTAIL.n343 9.3005
R664 VTAIL.n349 VTAIL.n348 9.3005
R665 VTAIL.n371 VTAIL.n370 9.3005
R666 VTAIL.n373 VTAIL.n372 9.3005
R667 VTAIL.n332 VTAIL.n331 9.3005
R668 VTAIL.n379 VTAIL.n378 9.3005
R669 VTAIL.n381 VTAIL.n380 9.3005
R670 VTAIL.n328 VTAIL.n327 9.3005
R671 VTAIL.n387 VTAIL.n386 9.3005
R672 VTAIL.n389 VTAIL.n388 9.3005
R673 VTAIL.n390 VTAIL.n323 9.3005
R674 VTAIL.n101 VTAIL.n100 9.3005
R675 VTAIL.n4 VTAIL.n3 9.3005
R676 VTAIL.n95 VTAIL.n94 9.3005
R677 VTAIL.n93 VTAIL.n92 9.3005
R678 VTAIL.n8 VTAIL.n7 9.3005
R679 VTAIL.n87 VTAIL.n86 9.3005
R680 VTAIL.n85 VTAIL.n84 9.3005
R681 VTAIL.n24 VTAIL.n23 9.3005
R682 VTAIL.n53 VTAIL.n52 9.3005
R683 VTAIL.n51 VTAIL.n50 9.3005
R684 VTAIL.n28 VTAIL.n27 9.3005
R685 VTAIL.n45 VTAIL.n44 9.3005
R686 VTAIL.n43 VTAIL.n42 9.3005
R687 VTAIL.n32 VTAIL.n31 9.3005
R688 VTAIL.n37 VTAIL.n36 9.3005
R689 VTAIL.n59 VTAIL.n58 9.3005
R690 VTAIL.n61 VTAIL.n60 9.3005
R691 VTAIL.n20 VTAIL.n19 9.3005
R692 VTAIL.n67 VTAIL.n66 9.3005
R693 VTAIL.n69 VTAIL.n68 9.3005
R694 VTAIL.n16 VTAIL.n15 9.3005
R695 VTAIL.n75 VTAIL.n74 9.3005
R696 VTAIL.n77 VTAIL.n76 9.3005
R697 VTAIL.n78 VTAIL.n11 9.3005
R698 VTAIL.n272 VTAIL.n271 9.3005
R699 VTAIL.n231 VTAIL.n230 9.3005
R700 VTAIL.n278 VTAIL.n277 9.3005
R701 VTAIL.n280 VTAIL.n279 9.3005
R702 VTAIL.n227 VTAIL.n226 9.3005
R703 VTAIL.n286 VTAIL.n285 9.3005
R704 VTAIL.n288 VTAIL.n287 9.3005
R705 VTAIL.n224 VTAIL.n221 9.3005
R706 VTAIL.n311 VTAIL.n310 9.3005
R707 VTAIL.n214 VTAIL.n213 9.3005
R708 VTAIL.n305 VTAIL.n304 9.3005
R709 VTAIL.n303 VTAIL.n302 9.3005
R710 VTAIL.n218 VTAIL.n217 9.3005
R711 VTAIL.n297 VTAIL.n296 9.3005
R712 VTAIL.n295 VTAIL.n294 9.3005
R713 VTAIL.n270 VTAIL.n269 9.3005
R714 VTAIL.n235 VTAIL.n234 9.3005
R715 VTAIL.n264 VTAIL.n263 9.3005
R716 VTAIL.n262 VTAIL.n261 9.3005
R717 VTAIL.n239 VTAIL.n238 9.3005
R718 VTAIL.n256 VTAIL.n255 9.3005
R719 VTAIL.n254 VTAIL.n253 9.3005
R720 VTAIL.n243 VTAIL.n242 9.3005
R721 VTAIL.n248 VTAIL.n247 9.3005
R722 VTAIL.n168 VTAIL.n167 9.3005
R723 VTAIL.n127 VTAIL.n126 9.3005
R724 VTAIL.n174 VTAIL.n173 9.3005
R725 VTAIL.n176 VTAIL.n175 9.3005
R726 VTAIL.n123 VTAIL.n122 9.3005
R727 VTAIL.n182 VTAIL.n181 9.3005
R728 VTAIL.n184 VTAIL.n183 9.3005
R729 VTAIL.n120 VTAIL.n117 9.3005
R730 VTAIL.n207 VTAIL.n206 9.3005
R731 VTAIL.n110 VTAIL.n109 9.3005
R732 VTAIL.n201 VTAIL.n200 9.3005
R733 VTAIL.n199 VTAIL.n198 9.3005
R734 VTAIL.n114 VTAIL.n113 9.3005
R735 VTAIL.n193 VTAIL.n192 9.3005
R736 VTAIL.n191 VTAIL.n190 9.3005
R737 VTAIL.n166 VTAIL.n165 9.3005
R738 VTAIL.n131 VTAIL.n130 9.3005
R739 VTAIL.n160 VTAIL.n159 9.3005
R740 VTAIL.n158 VTAIL.n157 9.3005
R741 VTAIL.n135 VTAIL.n134 9.3005
R742 VTAIL.n152 VTAIL.n151 9.3005
R743 VTAIL.n150 VTAIL.n149 9.3005
R744 VTAIL.n139 VTAIL.n138 9.3005
R745 VTAIL.n144 VTAIL.n143 9.3005
R746 VTAIL.n362 VTAIL.n338 8.92171
R747 VTAIL.n378 VTAIL.n377 8.92171
R748 VTAIL.n411 VTAIL.n316 8.92171
R749 VTAIL.n50 VTAIL.n26 8.92171
R750 VTAIL.n66 VTAIL.n65 8.92171
R751 VTAIL.n99 VTAIL.n4 8.92171
R752 VTAIL.n309 VTAIL.n214 8.92171
R753 VTAIL.n277 VTAIL.n276 8.92171
R754 VTAIL.n261 VTAIL.n237 8.92171
R755 VTAIL.n205 VTAIL.n110 8.92171
R756 VTAIL.n173 VTAIL.n172 8.92171
R757 VTAIL.n157 VTAIL.n133 8.92171
R758 VTAIL.n366 VTAIL.n365 8.14595
R759 VTAIL.n374 VTAIL.n332 8.14595
R760 VTAIL.n412 VTAIL.n314 8.14595
R761 VTAIL.n54 VTAIL.n53 8.14595
R762 VTAIL.n62 VTAIL.n20 8.14595
R763 VTAIL.n100 VTAIL.n2 8.14595
R764 VTAIL.n310 VTAIL.n212 8.14595
R765 VTAIL.n273 VTAIL.n231 8.14595
R766 VTAIL.n265 VTAIL.n264 8.14595
R767 VTAIL.n206 VTAIL.n108 8.14595
R768 VTAIL.n169 VTAIL.n127 8.14595
R769 VTAIL.n161 VTAIL.n160 8.14595
R770 VTAIL.n369 VTAIL.n336 7.3702
R771 VTAIL.n373 VTAIL.n334 7.3702
R772 VTAIL.n57 VTAIL.n24 7.3702
R773 VTAIL.n61 VTAIL.n22 7.3702
R774 VTAIL.n272 VTAIL.n233 7.3702
R775 VTAIL.n268 VTAIL.n235 7.3702
R776 VTAIL.n168 VTAIL.n129 7.3702
R777 VTAIL.n164 VTAIL.n131 7.3702
R778 VTAIL.n370 VTAIL.n369 6.59444
R779 VTAIL.n370 VTAIL.n334 6.59444
R780 VTAIL.n58 VTAIL.n57 6.59444
R781 VTAIL.n58 VTAIL.n22 6.59444
R782 VTAIL.n269 VTAIL.n233 6.59444
R783 VTAIL.n269 VTAIL.n268 6.59444
R784 VTAIL.n165 VTAIL.n129 6.59444
R785 VTAIL.n165 VTAIL.n164 6.59444
R786 VTAIL.n366 VTAIL.n336 5.81868
R787 VTAIL.n374 VTAIL.n373 5.81868
R788 VTAIL.n414 VTAIL.n314 5.81868
R789 VTAIL.n54 VTAIL.n24 5.81868
R790 VTAIL.n62 VTAIL.n61 5.81868
R791 VTAIL.n102 VTAIL.n2 5.81868
R792 VTAIL.n312 VTAIL.n212 5.81868
R793 VTAIL.n273 VTAIL.n272 5.81868
R794 VTAIL.n265 VTAIL.n235 5.81868
R795 VTAIL.n208 VTAIL.n108 5.81868
R796 VTAIL.n169 VTAIL.n168 5.81868
R797 VTAIL.n161 VTAIL.n131 5.81868
R798 VTAIL.n365 VTAIL.n338 5.04292
R799 VTAIL.n377 VTAIL.n332 5.04292
R800 VTAIL.n412 VTAIL.n411 5.04292
R801 VTAIL.n53 VTAIL.n26 5.04292
R802 VTAIL.n65 VTAIL.n20 5.04292
R803 VTAIL.n100 VTAIL.n99 5.04292
R804 VTAIL.n310 VTAIL.n309 5.04292
R805 VTAIL.n276 VTAIL.n231 5.04292
R806 VTAIL.n264 VTAIL.n237 5.04292
R807 VTAIL.n206 VTAIL.n205 5.04292
R808 VTAIL.n172 VTAIL.n127 5.04292
R809 VTAIL.n160 VTAIL.n133 5.04292
R810 VTAIL.n348 VTAIL.n347 4.38563
R811 VTAIL.n36 VTAIL.n35 4.38563
R812 VTAIL.n247 VTAIL.n246 4.38563
R813 VTAIL.n143 VTAIL.n142 4.38563
R814 VTAIL.n362 VTAIL.n361 4.26717
R815 VTAIL.n378 VTAIL.n330 4.26717
R816 VTAIL.n408 VTAIL.n316 4.26717
R817 VTAIL.n50 VTAIL.n49 4.26717
R818 VTAIL.n66 VTAIL.n18 4.26717
R819 VTAIL.n96 VTAIL.n4 4.26717
R820 VTAIL.n306 VTAIL.n214 4.26717
R821 VTAIL.n277 VTAIL.n229 4.26717
R822 VTAIL.n261 VTAIL.n260 4.26717
R823 VTAIL.n202 VTAIL.n110 4.26717
R824 VTAIL.n173 VTAIL.n125 4.26717
R825 VTAIL.n157 VTAIL.n156 4.26717
R826 VTAIL.n358 VTAIL.n340 3.49141
R827 VTAIL.n382 VTAIL.n381 3.49141
R828 VTAIL.n407 VTAIL.n318 3.49141
R829 VTAIL.n46 VTAIL.n28 3.49141
R830 VTAIL.n70 VTAIL.n69 3.49141
R831 VTAIL.n95 VTAIL.n6 3.49141
R832 VTAIL.n305 VTAIL.n216 3.49141
R833 VTAIL.n281 VTAIL.n280 3.49141
R834 VTAIL.n257 VTAIL.n239 3.49141
R835 VTAIL.n201 VTAIL.n112 3.49141
R836 VTAIL.n177 VTAIL.n176 3.49141
R837 VTAIL.n153 VTAIL.n135 3.49141
R838 VTAIL.n357 VTAIL.n342 2.71565
R839 VTAIL.n385 VTAIL.n328 2.71565
R840 VTAIL.n404 VTAIL.n403 2.71565
R841 VTAIL.n45 VTAIL.n30 2.71565
R842 VTAIL.n73 VTAIL.n16 2.71565
R843 VTAIL.n92 VTAIL.n91 2.71565
R844 VTAIL.n302 VTAIL.n301 2.71565
R845 VTAIL.n284 VTAIL.n227 2.71565
R846 VTAIL.n256 VTAIL.n241 2.71565
R847 VTAIL.n198 VTAIL.n197 2.71565
R848 VTAIL.n180 VTAIL.n123 2.71565
R849 VTAIL.n152 VTAIL.n137 2.71565
R850 VTAIL.n354 VTAIL.n353 1.93989
R851 VTAIL.n386 VTAIL.n326 1.93989
R852 VTAIL.n400 VTAIL.n320 1.93989
R853 VTAIL.n42 VTAIL.n41 1.93989
R854 VTAIL.n74 VTAIL.n14 1.93989
R855 VTAIL.n88 VTAIL.n8 1.93989
R856 VTAIL.n298 VTAIL.n218 1.93989
R857 VTAIL.n285 VTAIL.n225 1.93989
R858 VTAIL.n253 VTAIL.n252 1.93989
R859 VTAIL.n194 VTAIL.n114 1.93989
R860 VTAIL.n181 VTAIL.n121 1.93989
R861 VTAIL.n149 VTAIL.n148 1.93989
R862 VTAIL.n209 VTAIL.n107 1.52636
R863 VTAIL.n313 VTAIL.n211 1.52636
R864 VTAIL.n105 VTAIL.n103 1.52636
R865 VTAIL.n211 VTAIL.n209 1.23326
R866 VTAIL.n103 VTAIL.n1 1.23326
R867 VTAIL.n350 VTAIL.n344 1.16414
R868 VTAIL.n391 VTAIL.n389 1.16414
R869 VTAIL.n399 VTAIL.n322 1.16414
R870 VTAIL.n38 VTAIL.n32 1.16414
R871 VTAIL.n79 VTAIL.n77 1.16414
R872 VTAIL.n87 VTAIL.n10 1.16414
R873 VTAIL.n297 VTAIL.n220 1.16414
R874 VTAIL.n289 VTAIL.n288 1.16414
R875 VTAIL.n249 VTAIL.n243 1.16414
R876 VTAIL.n193 VTAIL.n116 1.16414
R877 VTAIL.n185 VTAIL.n184 1.16414
R878 VTAIL.n145 VTAIL.n139 1.16414
R879 VTAIL.n0 VTAIL.t2 1.09081
R880 VTAIL.n0 VTAIL.t0 1.09081
R881 VTAIL.n104 VTAIL.t8 1.09081
R882 VTAIL.n104 VTAIL.t9 1.09081
R883 VTAIL.n210 VTAIL.t7 1.09081
R884 VTAIL.n210 VTAIL.t10 1.09081
R885 VTAIL.n106 VTAIL.t1 1.09081
R886 VTAIL.n106 VTAIL.t4 1.09081
R887 VTAIL VTAIL.n415 1.08671
R888 VTAIL VTAIL.n1 0.440155
R889 VTAIL.n349 VTAIL.n346 0.388379
R890 VTAIL.n390 VTAIL.n324 0.388379
R891 VTAIL.n396 VTAIL.n395 0.388379
R892 VTAIL.n37 VTAIL.n34 0.388379
R893 VTAIL.n78 VTAIL.n12 0.388379
R894 VTAIL.n84 VTAIL.n83 0.388379
R895 VTAIL.n294 VTAIL.n293 0.388379
R896 VTAIL.n224 VTAIL.n222 0.388379
R897 VTAIL.n248 VTAIL.n245 0.388379
R898 VTAIL.n190 VTAIL.n189 0.388379
R899 VTAIL.n120 VTAIL.n118 0.388379
R900 VTAIL.n144 VTAIL.n141 0.388379
R901 VTAIL.n348 VTAIL.n343 0.155672
R902 VTAIL.n355 VTAIL.n343 0.155672
R903 VTAIL.n356 VTAIL.n355 0.155672
R904 VTAIL.n356 VTAIL.n339 0.155672
R905 VTAIL.n363 VTAIL.n339 0.155672
R906 VTAIL.n364 VTAIL.n363 0.155672
R907 VTAIL.n364 VTAIL.n335 0.155672
R908 VTAIL.n371 VTAIL.n335 0.155672
R909 VTAIL.n372 VTAIL.n371 0.155672
R910 VTAIL.n372 VTAIL.n331 0.155672
R911 VTAIL.n379 VTAIL.n331 0.155672
R912 VTAIL.n380 VTAIL.n379 0.155672
R913 VTAIL.n380 VTAIL.n327 0.155672
R914 VTAIL.n387 VTAIL.n327 0.155672
R915 VTAIL.n388 VTAIL.n387 0.155672
R916 VTAIL.n388 VTAIL.n323 0.155672
R917 VTAIL.n397 VTAIL.n323 0.155672
R918 VTAIL.n398 VTAIL.n397 0.155672
R919 VTAIL.n398 VTAIL.n319 0.155672
R920 VTAIL.n405 VTAIL.n319 0.155672
R921 VTAIL.n406 VTAIL.n405 0.155672
R922 VTAIL.n406 VTAIL.n315 0.155672
R923 VTAIL.n413 VTAIL.n315 0.155672
R924 VTAIL.n36 VTAIL.n31 0.155672
R925 VTAIL.n43 VTAIL.n31 0.155672
R926 VTAIL.n44 VTAIL.n43 0.155672
R927 VTAIL.n44 VTAIL.n27 0.155672
R928 VTAIL.n51 VTAIL.n27 0.155672
R929 VTAIL.n52 VTAIL.n51 0.155672
R930 VTAIL.n52 VTAIL.n23 0.155672
R931 VTAIL.n59 VTAIL.n23 0.155672
R932 VTAIL.n60 VTAIL.n59 0.155672
R933 VTAIL.n60 VTAIL.n19 0.155672
R934 VTAIL.n67 VTAIL.n19 0.155672
R935 VTAIL.n68 VTAIL.n67 0.155672
R936 VTAIL.n68 VTAIL.n15 0.155672
R937 VTAIL.n75 VTAIL.n15 0.155672
R938 VTAIL.n76 VTAIL.n75 0.155672
R939 VTAIL.n76 VTAIL.n11 0.155672
R940 VTAIL.n85 VTAIL.n11 0.155672
R941 VTAIL.n86 VTAIL.n85 0.155672
R942 VTAIL.n86 VTAIL.n7 0.155672
R943 VTAIL.n93 VTAIL.n7 0.155672
R944 VTAIL.n94 VTAIL.n93 0.155672
R945 VTAIL.n94 VTAIL.n3 0.155672
R946 VTAIL.n101 VTAIL.n3 0.155672
R947 VTAIL.n311 VTAIL.n213 0.155672
R948 VTAIL.n304 VTAIL.n213 0.155672
R949 VTAIL.n304 VTAIL.n303 0.155672
R950 VTAIL.n303 VTAIL.n217 0.155672
R951 VTAIL.n296 VTAIL.n217 0.155672
R952 VTAIL.n296 VTAIL.n295 0.155672
R953 VTAIL.n295 VTAIL.n221 0.155672
R954 VTAIL.n287 VTAIL.n221 0.155672
R955 VTAIL.n287 VTAIL.n286 0.155672
R956 VTAIL.n286 VTAIL.n226 0.155672
R957 VTAIL.n279 VTAIL.n226 0.155672
R958 VTAIL.n279 VTAIL.n278 0.155672
R959 VTAIL.n278 VTAIL.n230 0.155672
R960 VTAIL.n271 VTAIL.n230 0.155672
R961 VTAIL.n271 VTAIL.n270 0.155672
R962 VTAIL.n270 VTAIL.n234 0.155672
R963 VTAIL.n263 VTAIL.n234 0.155672
R964 VTAIL.n263 VTAIL.n262 0.155672
R965 VTAIL.n262 VTAIL.n238 0.155672
R966 VTAIL.n255 VTAIL.n238 0.155672
R967 VTAIL.n255 VTAIL.n254 0.155672
R968 VTAIL.n254 VTAIL.n242 0.155672
R969 VTAIL.n247 VTAIL.n242 0.155672
R970 VTAIL.n207 VTAIL.n109 0.155672
R971 VTAIL.n200 VTAIL.n109 0.155672
R972 VTAIL.n200 VTAIL.n199 0.155672
R973 VTAIL.n199 VTAIL.n113 0.155672
R974 VTAIL.n192 VTAIL.n113 0.155672
R975 VTAIL.n192 VTAIL.n191 0.155672
R976 VTAIL.n191 VTAIL.n117 0.155672
R977 VTAIL.n183 VTAIL.n117 0.155672
R978 VTAIL.n183 VTAIL.n182 0.155672
R979 VTAIL.n182 VTAIL.n122 0.155672
R980 VTAIL.n175 VTAIL.n122 0.155672
R981 VTAIL.n175 VTAIL.n174 0.155672
R982 VTAIL.n174 VTAIL.n126 0.155672
R983 VTAIL.n167 VTAIL.n126 0.155672
R984 VTAIL.n167 VTAIL.n166 0.155672
R985 VTAIL.n166 VTAIL.n130 0.155672
R986 VTAIL.n159 VTAIL.n130 0.155672
R987 VTAIL.n159 VTAIL.n158 0.155672
R988 VTAIL.n158 VTAIL.n134 0.155672
R989 VTAIL.n151 VTAIL.n134 0.155672
R990 VTAIL.n151 VTAIL.n150 0.155672
R991 VTAIL.n150 VTAIL.n138 0.155672
R992 VTAIL.n143 VTAIL.n138 0.155672
R993 B.n891 B.n890 585
R994 B.n892 B.n891 585
R995 B.n381 B.n120 585
R996 B.n380 B.n379 585
R997 B.n378 B.n377 585
R998 B.n376 B.n375 585
R999 B.n374 B.n373 585
R1000 B.n372 B.n371 585
R1001 B.n370 B.n369 585
R1002 B.n368 B.n367 585
R1003 B.n366 B.n365 585
R1004 B.n364 B.n363 585
R1005 B.n362 B.n361 585
R1006 B.n360 B.n359 585
R1007 B.n358 B.n357 585
R1008 B.n356 B.n355 585
R1009 B.n354 B.n353 585
R1010 B.n352 B.n351 585
R1011 B.n350 B.n349 585
R1012 B.n348 B.n347 585
R1013 B.n346 B.n345 585
R1014 B.n344 B.n343 585
R1015 B.n342 B.n341 585
R1016 B.n340 B.n339 585
R1017 B.n338 B.n337 585
R1018 B.n336 B.n335 585
R1019 B.n334 B.n333 585
R1020 B.n332 B.n331 585
R1021 B.n330 B.n329 585
R1022 B.n328 B.n327 585
R1023 B.n326 B.n325 585
R1024 B.n324 B.n323 585
R1025 B.n322 B.n321 585
R1026 B.n320 B.n319 585
R1027 B.n318 B.n317 585
R1028 B.n316 B.n315 585
R1029 B.n314 B.n313 585
R1030 B.n312 B.n311 585
R1031 B.n310 B.n309 585
R1032 B.n308 B.n307 585
R1033 B.n306 B.n305 585
R1034 B.n304 B.n303 585
R1035 B.n302 B.n301 585
R1036 B.n300 B.n299 585
R1037 B.n298 B.n297 585
R1038 B.n296 B.n295 585
R1039 B.n294 B.n293 585
R1040 B.n292 B.n291 585
R1041 B.n290 B.n289 585
R1042 B.n288 B.n287 585
R1043 B.n286 B.n285 585
R1044 B.n284 B.n283 585
R1045 B.n282 B.n281 585
R1046 B.n280 B.n279 585
R1047 B.n278 B.n277 585
R1048 B.n276 B.n275 585
R1049 B.n274 B.n273 585
R1050 B.n272 B.n271 585
R1051 B.n270 B.n269 585
R1052 B.n268 B.n267 585
R1053 B.n266 B.n265 585
R1054 B.n263 B.n262 585
R1055 B.n261 B.n260 585
R1056 B.n259 B.n258 585
R1057 B.n257 B.n256 585
R1058 B.n255 B.n254 585
R1059 B.n253 B.n252 585
R1060 B.n251 B.n250 585
R1061 B.n249 B.n248 585
R1062 B.n247 B.n246 585
R1063 B.n245 B.n244 585
R1064 B.n243 B.n242 585
R1065 B.n241 B.n240 585
R1066 B.n239 B.n238 585
R1067 B.n237 B.n236 585
R1068 B.n235 B.n234 585
R1069 B.n233 B.n232 585
R1070 B.n231 B.n230 585
R1071 B.n229 B.n228 585
R1072 B.n227 B.n226 585
R1073 B.n225 B.n224 585
R1074 B.n223 B.n222 585
R1075 B.n221 B.n220 585
R1076 B.n219 B.n218 585
R1077 B.n217 B.n216 585
R1078 B.n215 B.n214 585
R1079 B.n213 B.n212 585
R1080 B.n211 B.n210 585
R1081 B.n209 B.n208 585
R1082 B.n207 B.n206 585
R1083 B.n205 B.n204 585
R1084 B.n203 B.n202 585
R1085 B.n201 B.n200 585
R1086 B.n199 B.n198 585
R1087 B.n197 B.n196 585
R1088 B.n195 B.n194 585
R1089 B.n193 B.n192 585
R1090 B.n191 B.n190 585
R1091 B.n189 B.n188 585
R1092 B.n187 B.n186 585
R1093 B.n185 B.n184 585
R1094 B.n183 B.n182 585
R1095 B.n181 B.n180 585
R1096 B.n179 B.n178 585
R1097 B.n177 B.n176 585
R1098 B.n175 B.n174 585
R1099 B.n173 B.n172 585
R1100 B.n171 B.n170 585
R1101 B.n169 B.n168 585
R1102 B.n167 B.n166 585
R1103 B.n165 B.n164 585
R1104 B.n163 B.n162 585
R1105 B.n161 B.n160 585
R1106 B.n159 B.n158 585
R1107 B.n157 B.n156 585
R1108 B.n155 B.n154 585
R1109 B.n153 B.n152 585
R1110 B.n151 B.n150 585
R1111 B.n149 B.n148 585
R1112 B.n147 B.n146 585
R1113 B.n145 B.n144 585
R1114 B.n143 B.n142 585
R1115 B.n141 B.n140 585
R1116 B.n139 B.n138 585
R1117 B.n137 B.n136 585
R1118 B.n135 B.n134 585
R1119 B.n133 B.n132 585
R1120 B.n131 B.n130 585
R1121 B.n129 B.n128 585
R1122 B.n127 B.n126 585
R1123 B.n889 B.n55 585
R1124 B.n893 B.n55 585
R1125 B.n888 B.n54 585
R1126 B.n894 B.n54 585
R1127 B.n887 B.n886 585
R1128 B.n886 B.n50 585
R1129 B.n885 B.n49 585
R1130 B.n900 B.n49 585
R1131 B.n884 B.n48 585
R1132 B.n901 B.n48 585
R1133 B.n883 B.n47 585
R1134 B.n902 B.n47 585
R1135 B.n882 B.n881 585
R1136 B.n881 B.n43 585
R1137 B.n880 B.n42 585
R1138 B.n908 B.n42 585
R1139 B.n879 B.n41 585
R1140 B.n909 B.n41 585
R1141 B.n878 B.n40 585
R1142 B.n910 B.n40 585
R1143 B.n877 B.n876 585
R1144 B.n876 B.n36 585
R1145 B.n875 B.n35 585
R1146 B.n916 B.n35 585
R1147 B.n874 B.n34 585
R1148 B.n917 B.n34 585
R1149 B.n873 B.n33 585
R1150 B.n918 B.n33 585
R1151 B.n872 B.n871 585
R1152 B.n871 B.n32 585
R1153 B.n870 B.n28 585
R1154 B.n924 B.n28 585
R1155 B.n869 B.n27 585
R1156 B.n925 B.n27 585
R1157 B.n868 B.n26 585
R1158 B.n926 B.n26 585
R1159 B.n867 B.n866 585
R1160 B.n866 B.n22 585
R1161 B.n865 B.n21 585
R1162 B.n932 B.n21 585
R1163 B.n864 B.n20 585
R1164 B.n933 B.n20 585
R1165 B.n863 B.n19 585
R1166 B.n934 B.n19 585
R1167 B.n862 B.n861 585
R1168 B.n861 B.n15 585
R1169 B.n860 B.n14 585
R1170 B.n940 B.n14 585
R1171 B.n859 B.n13 585
R1172 B.n941 B.n13 585
R1173 B.n858 B.n12 585
R1174 B.n942 B.n12 585
R1175 B.n857 B.n856 585
R1176 B.n856 B.n8 585
R1177 B.n855 B.n7 585
R1178 B.n948 B.n7 585
R1179 B.n854 B.n6 585
R1180 B.n949 B.n6 585
R1181 B.n853 B.n5 585
R1182 B.n950 B.n5 585
R1183 B.n852 B.n851 585
R1184 B.n851 B.n4 585
R1185 B.n850 B.n382 585
R1186 B.n850 B.n849 585
R1187 B.n840 B.n383 585
R1188 B.n384 B.n383 585
R1189 B.n842 B.n841 585
R1190 B.n843 B.n842 585
R1191 B.n839 B.n388 585
R1192 B.n392 B.n388 585
R1193 B.n838 B.n837 585
R1194 B.n837 B.n836 585
R1195 B.n390 B.n389 585
R1196 B.n391 B.n390 585
R1197 B.n829 B.n828 585
R1198 B.n830 B.n829 585
R1199 B.n827 B.n397 585
R1200 B.n397 B.n396 585
R1201 B.n826 B.n825 585
R1202 B.n825 B.n824 585
R1203 B.n399 B.n398 585
R1204 B.n400 B.n399 585
R1205 B.n817 B.n816 585
R1206 B.n818 B.n817 585
R1207 B.n815 B.n405 585
R1208 B.n405 B.n404 585
R1209 B.n814 B.n813 585
R1210 B.n813 B.n812 585
R1211 B.n407 B.n406 585
R1212 B.n805 B.n407 585
R1213 B.n804 B.n803 585
R1214 B.n806 B.n804 585
R1215 B.n802 B.n412 585
R1216 B.n412 B.n411 585
R1217 B.n801 B.n800 585
R1218 B.n800 B.n799 585
R1219 B.n414 B.n413 585
R1220 B.n415 B.n414 585
R1221 B.n792 B.n791 585
R1222 B.n793 B.n792 585
R1223 B.n790 B.n420 585
R1224 B.n420 B.n419 585
R1225 B.n789 B.n788 585
R1226 B.n788 B.n787 585
R1227 B.n422 B.n421 585
R1228 B.n423 B.n422 585
R1229 B.n780 B.n779 585
R1230 B.n781 B.n780 585
R1231 B.n778 B.n428 585
R1232 B.n428 B.n427 585
R1233 B.n777 B.n776 585
R1234 B.n776 B.n775 585
R1235 B.n430 B.n429 585
R1236 B.n431 B.n430 585
R1237 B.n768 B.n767 585
R1238 B.n769 B.n768 585
R1239 B.n766 B.n436 585
R1240 B.n436 B.n435 585
R1241 B.n760 B.n759 585
R1242 B.n758 B.n502 585
R1243 B.n757 B.n501 585
R1244 B.n762 B.n501 585
R1245 B.n756 B.n755 585
R1246 B.n754 B.n753 585
R1247 B.n752 B.n751 585
R1248 B.n750 B.n749 585
R1249 B.n748 B.n747 585
R1250 B.n746 B.n745 585
R1251 B.n744 B.n743 585
R1252 B.n742 B.n741 585
R1253 B.n740 B.n739 585
R1254 B.n738 B.n737 585
R1255 B.n736 B.n735 585
R1256 B.n734 B.n733 585
R1257 B.n732 B.n731 585
R1258 B.n730 B.n729 585
R1259 B.n728 B.n727 585
R1260 B.n726 B.n725 585
R1261 B.n724 B.n723 585
R1262 B.n722 B.n721 585
R1263 B.n720 B.n719 585
R1264 B.n718 B.n717 585
R1265 B.n716 B.n715 585
R1266 B.n714 B.n713 585
R1267 B.n712 B.n711 585
R1268 B.n710 B.n709 585
R1269 B.n708 B.n707 585
R1270 B.n706 B.n705 585
R1271 B.n704 B.n703 585
R1272 B.n702 B.n701 585
R1273 B.n700 B.n699 585
R1274 B.n698 B.n697 585
R1275 B.n696 B.n695 585
R1276 B.n694 B.n693 585
R1277 B.n692 B.n691 585
R1278 B.n690 B.n689 585
R1279 B.n688 B.n687 585
R1280 B.n686 B.n685 585
R1281 B.n684 B.n683 585
R1282 B.n682 B.n681 585
R1283 B.n680 B.n679 585
R1284 B.n678 B.n677 585
R1285 B.n676 B.n675 585
R1286 B.n674 B.n673 585
R1287 B.n672 B.n671 585
R1288 B.n670 B.n669 585
R1289 B.n668 B.n667 585
R1290 B.n666 B.n665 585
R1291 B.n664 B.n663 585
R1292 B.n662 B.n661 585
R1293 B.n660 B.n659 585
R1294 B.n658 B.n657 585
R1295 B.n656 B.n655 585
R1296 B.n654 B.n653 585
R1297 B.n652 B.n651 585
R1298 B.n650 B.n649 585
R1299 B.n648 B.n647 585
R1300 B.n646 B.n645 585
R1301 B.n644 B.n643 585
R1302 B.n641 B.n640 585
R1303 B.n639 B.n638 585
R1304 B.n637 B.n636 585
R1305 B.n635 B.n634 585
R1306 B.n633 B.n632 585
R1307 B.n631 B.n630 585
R1308 B.n629 B.n628 585
R1309 B.n627 B.n626 585
R1310 B.n625 B.n624 585
R1311 B.n623 B.n622 585
R1312 B.n621 B.n620 585
R1313 B.n619 B.n618 585
R1314 B.n617 B.n616 585
R1315 B.n615 B.n614 585
R1316 B.n613 B.n612 585
R1317 B.n611 B.n610 585
R1318 B.n609 B.n608 585
R1319 B.n607 B.n606 585
R1320 B.n605 B.n604 585
R1321 B.n603 B.n602 585
R1322 B.n601 B.n600 585
R1323 B.n599 B.n598 585
R1324 B.n597 B.n596 585
R1325 B.n595 B.n594 585
R1326 B.n593 B.n592 585
R1327 B.n591 B.n590 585
R1328 B.n589 B.n588 585
R1329 B.n587 B.n586 585
R1330 B.n585 B.n584 585
R1331 B.n583 B.n582 585
R1332 B.n581 B.n580 585
R1333 B.n579 B.n578 585
R1334 B.n577 B.n576 585
R1335 B.n575 B.n574 585
R1336 B.n573 B.n572 585
R1337 B.n571 B.n570 585
R1338 B.n569 B.n568 585
R1339 B.n567 B.n566 585
R1340 B.n565 B.n564 585
R1341 B.n563 B.n562 585
R1342 B.n561 B.n560 585
R1343 B.n559 B.n558 585
R1344 B.n557 B.n556 585
R1345 B.n555 B.n554 585
R1346 B.n553 B.n552 585
R1347 B.n551 B.n550 585
R1348 B.n549 B.n548 585
R1349 B.n547 B.n546 585
R1350 B.n545 B.n544 585
R1351 B.n543 B.n542 585
R1352 B.n541 B.n540 585
R1353 B.n539 B.n538 585
R1354 B.n537 B.n536 585
R1355 B.n535 B.n534 585
R1356 B.n533 B.n532 585
R1357 B.n531 B.n530 585
R1358 B.n529 B.n528 585
R1359 B.n527 B.n526 585
R1360 B.n525 B.n524 585
R1361 B.n523 B.n522 585
R1362 B.n521 B.n520 585
R1363 B.n519 B.n518 585
R1364 B.n517 B.n516 585
R1365 B.n515 B.n514 585
R1366 B.n513 B.n512 585
R1367 B.n511 B.n510 585
R1368 B.n509 B.n508 585
R1369 B.n438 B.n437 585
R1370 B.n765 B.n764 585
R1371 B.n434 B.n433 585
R1372 B.n435 B.n434 585
R1373 B.n771 B.n770 585
R1374 B.n770 B.n769 585
R1375 B.n772 B.n432 585
R1376 B.n432 B.n431 585
R1377 B.n774 B.n773 585
R1378 B.n775 B.n774 585
R1379 B.n426 B.n425 585
R1380 B.n427 B.n426 585
R1381 B.n783 B.n782 585
R1382 B.n782 B.n781 585
R1383 B.n784 B.n424 585
R1384 B.n424 B.n423 585
R1385 B.n786 B.n785 585
R1386 B.n787 B.n786 585
R1387 B.n418 B.n417 585
R1388 B.n419 B.n418 585
R1389 B.n795 B.n794 585
R1390 B.n794 B.n793 585
R1391 B.n796 B.n416 585
R1392 B.n416 B.n415 585
R1393 B.n798 B.n797 585
R1394 B.n799 B.n798 585
R1395 B.n410 B.n409 585
R1396 B.n411 B.n410 585
R1397 B.n808 B.n807 585
R1398 B.n807 B.n806 585
R1399 B.n809 B.n408 585
R1400 B.n805 B.n408 585
R1401 B.n811 B.n810 585
R1402 B.n812 B.n811 585
R1403 B.n403 B.n402 585
R1404 B.n404 B.n403 585
R1405 B.n820 B.n819 585
R1406 B.n819 B.n818 585
R1407 B.n821 B.n401 585
R1408 B.n401 B.n400 585
R1409 B.n823 B.n822 585
R1410 B.n824 B.n823 585
R1411 B.n395 B.n394 585
R1412 B.n396 B.n395 585
R1413 B.n832 B.n831 585
R1414 B.n831 B.n830 585
R1415 B.n833 B.n393 585
R1416 B.n393 B.n391 585
R1417 B.n835 B.n834 585
R1418 B.n836 B.n835 585
R1419 B.n387 B.n386 585
R1420 B.n392 B.n387 585
R1421 B.n845 B.n844 585
R1422 B.n844 B.n843 585
R1423 B.n846 B.n385 585
R1424 B.n385 B.n384 585
R1425 B.n848 B.n847 585
R1426 B.n849 B.n848 585
R1427 B.n2 B.n0 585
R1428 B.n4 B.n2 585
R1429 B.n3 B.n1 585
R1430 B.n949 B.n3 585
R1431 B.n947 B.n946 585
R1432 B.n948 B.n947 585
R1433 B.n945 B.n9 585
R1434 B.n9 B.n8 585
R1435 B.n944 B.n943 585
R1436 B.n943 B.n942 585
R1437 B.n11 B.n10 585
R1438 B.n941 B.n11 585
R1439 B.n939 B.n938 585
R1440 B.n940 B.n939 585
R1441 B.n937 B.n16 585
R1442 B.n16 B.n15 585
R1443 B.n936 B.n935 585
R1444 B.n935 B.n934 585
R1445 B.n18 B.n17 585
R1446 B.n933 B.n18 585
R1447 B.n931 B.n930 585
R1448 B.n932 B.n931 585
R1449 B.n929 B.n23 585
R1450 B.n23 B.n22 585
R1451 B.n928 B.n927 585
R1452 B.n927 B.n926 585
R1453 B.n25 B.n24 585
R1454 B.n925 B.n25 585
R1455 B.n923 B.n922 585
R1456 B.n924 B.n923 585
R1457 B.n921 B.n29 585
R1458 B.n32 B.n29 585
R1459 B.n920 B.n919 585
R1460 B.n919 B.n918 585
R1461 B.n31 B.n30 585
R1462 B.n917 B.n31 585
R1463 B.n915 B.n914 585
R1464 B.n916 B.n915 585
R1465 B.n913 B.n37 585
R1466 B.n37 B.n36 585
R1467 B.n912 B.n911 585
R1468 B.n911 B.n910 585
R1469 B.n39 B.n38 585
R1470 B.n909 B.n39 585
R1471 B.n907 B.n906 585
R1472 B.n908 B.n907 585
R1473 B.n905 B.n44 585
R1474 B.n44 B.n43 585
R1475 B.n904 B.n903 585
R1476 B.n903 B.n902 585
R1477 B.n46 B.n45 585
R1478 B.n901 B.n46 585
R1479 B.n899 B.n898 585
R1480 B.n900 B.n899 585
R1481 B.n897 B.n51 585
R1482 B.n51 B.n50 585
R1483 B.n896 B.n895 585
R1484 B.n895 B.n894 585
R1485 B.n53 B.n52 585
R1486 B.n893 B.n53 585
R1487 B.n952 B.n951 585
R1488 B.n951 B.n950 585
R1489 B.n505 B.t6 509.137
R1490 B.n503 B.t10 509.137
R1491 B.n123 B.t17 509.137
R1492 B.n121 B.t13 509.137
R1493 B.n760 B.n434 492.5
R1494 B.n126 B.n53 492.5
R1495 B.n764 B.n436 492.5
R1496 B.n891 B.n55 492.5
R1497 B.n505 B.t9 422.522
R1498 B.n503 B.t12 422.522
R1499 B.n123 B.t18 422.522
R1500 B.n121 B.t15 422.522
R1501 B.n506 B.t8 388.195
R1502 B.n122 B.t16 388.195
R1503 B.n504 B.t11 388.195
R1504 B.n124 B.t19 388.195
R1505 B.n892 B.n119 256.663
R1506 B.n892 B.n118 256.663
R1507 B.n892 B.n117 256.663
R1508 B.n892 B.n116 256.663
R1509 B.n892 B.n115 256.663
R1510 B.n892 B.n114 256.663
R1511 B.n892 B.n113 256.663
R1512 B.n892 B.n112 256.663
R1513 B.n892 B.n111 256.663
R1514 B.n892 B.n110 256.663
R1515 B.n892 B.n109 256.663
R1516 B.n892 B.n108 256.663
R1517 B.n892 B.n107 256.663
R1518 B.n892 B.n106 256.663
R1519 B.n892 B.n105 256.663
R1520 B.n892 B.n104 256.663
R1521 B.n892 B.n103 256.663
R1522 B.n892 B.n102 256.663
R1523 B.n892 B.n101 256.663
R1524 B.n892 B.n100 256.663
R1525 B.n892 B.n99 256.663
R1526 B.n892 B.n98 256.663
R1527 B.n892 B.n97 256.663
R1528 B.n892 B.n96 256.663
R1529 B.n892 B.n95 256.663
R1530 B.n892 B.n94 256.663
R1531 B.n892 B.n93 256.663
R1532 B.n892 B.n92 256.663
R1533 B.n892 B.n91 256.663
R1534 B.n892 B.n90 256.663
R1535 B.n892 B.n89 256.663
R1536 B.n892 B.n88 256.663
R1537 B.n892 B.n87 256.663
R1538 B.n892 B.n86 256.663
R1539 B.n892 B.n85 256.663
R1540 B.n892 B.n84 256.663
R1541 B.n892 B.n83 256.663
R1542 B.n892 B.n82 256.663
R1543 B.n892 B.n81 256.663
R1544 B.n892 B.n80 256.663
R1545 B.n892 B.n79 256.663
R1546 B.n892 B.n78 256.663
R1547 B.n892 B.n77 256.663
R1548 B.n892 B.n76 256.663
R1549 B.n892 B.n75 256.663
R1550 B.n892 B.n74 256.663
R1551 B.n892 B.n73 256.663
R1552 B.n892 B.n72 256.663
R1553 B.n892 B.n71 256.663
R1554 B.n892 B.n70 256.663
R1555 B.n892 B.n69 256.663
R1556 B.n892 B.n68 256.663
R1557 B.n892 B.n67 256.663
R1558 B.n892 B.n66 256.663
R1559 B.n892 B.n65 256.663
R1560 B.n892 B.n64 256.663
R1561 B.n892 B.n63 256.663
R1562 B.n892 B.n62 256.663
R1563 B.n892 B.n61 256.663
R1564 B.n892 B.n60 256.663
R1565 B.n892 B.n59 256.663
R1566 B.n892 B.n58 256.663
R1567 B.n892 B.n57 256.663
R1568 B.n892 B.n56 256.663
R1569 B.n762 B.n761 256.663
R1570 B.n762 B.n439 256.663
R1571 B.n762 B.n440 256.663
R1572 B.n762 B.n441 256.663
R1573 B.n762 B.n442 256.663
R1574 B.n762 B.n443 256.663
R1575 B.n762 B.n444 256.663
R1576 B.n762 B.n445 256.663
R1577 B.n762 B.n446 256.663
R1578 B.n762 B.n447 256.663
R1579 B.n762 B.n448 256.663
R1580 B.n762 B.n449 256.663
R1581 B.n762 B.n450 256.663
R1582 B.n762 B.n451 256.663
R1583 B.n762 B.n452 256.663
R1584 B.n762 B.n453 256.663
R1585 B.n762 B.n454 256.663
R1586 B.n762 B.n455 256.663
R1587 B.n762 B.n456 256.663
R1588 B.n762 B.n457 256.663
R1589 B.n762 B.n458 256.663
R1590 B.n762 B.n459 256.663
R1591 B.n762 B.n460 256.663
R1592 B.n762 B.n461 256.663
R1593 B.n762 B.n462 256.663
R1594 B.n762 B.n463 256.663
R1595 B.n762 B.n464 256.663
R1596 B.n762 B.n465 256.663
R1597 B.n762 B.n466 256.663
R1598 B.n762 B.n467 256.663
R1599 B.n762 B.n468 256.663
R1600 B.n762 B.n469 256.663
R1601 B.n762 B.n470 256.663
R1602 B.n762 B.n471 256.663
R1603 B.n762 B.n472 256.663
R1604 B.n762 B.n473 256.663
R1605 B.n762 B.n474 256.663
R1606 B.n762 B.n475 256.663
R1607 B.n762 B.n476 256.663
R1608 B.n762 B.n477 256.663
R1609 B.n762 B.n478 256.663
R1610 B.n762 B.n479 256.663
R1611 B.n762 B.n480 256.663
R1612 B.n762 B.n481 256.663
R1613 B.n762 B.n482 256.663
R1614 B.n762 B.n483 256.663
R1615 B.n762 B.n484 256.663
R1616 B.n762 B.n485 256.663
R1617 B.n762 B.n486 256.663
R1618 B.n762 B.n487 256.663
R1619 B.n762 B.n488 256.663
R1620 B.n762 B.n489 256.663
R1621 B.n762 B.n490 256.663
R1622 B.n762 B.n491 256.663
R1623 B.n762 B.n492 256.663
R1624 B.n762 B.n493 256.663
R1625 B.n762 B.n494 256.663
R1626 B.n762 B.n495 256.663
R1627 B.n762 B.n496 256.663
R1628 B.n762 B.n497 256.663
R1629 B.n762 B.n498 256.663
R1630 B.n762 B.n499 256.663
R1631 B.n762 B.n500 256.663
R1632 B.n763 B.n762 256.663
R1633 B.n770 B.n434 163.367
R1634 B.n770 B.n432 163.367
R1635 B.n774 B.n432 163.367
R1636 B.n774 B.n426 163.367
R1637 B.n782 B.n426 163.367
R1638 B.n782 B.n424 163.367
R1639 B.n786 B.n424 163.367
R1640 B.n786 B.n418 163.367
R1641 B.n794 B.n418 163.367
R1642 B.n794 B.n416 163.367
R1643 B.n798 B.n416 163.367
R1644 B.n798 B.n410 163.367
R1645 B.n807 B.n410 163.367
R1646 B.n807 B.n408 163.367
R1647 B.n811 B.n408 163.367
R1648 B.n811 B.n403 163.367
R1649 B.n819 B.n403 163.367
R1650 B.n819 B.n401 163.367
R1651 B.n823 B.n401 163.367
R1652 B.n823 B.n395 163.367
R1653 B.n831 B.n395 163.367
R1654 B.n831 B.n393 163.367
R1655 B.n835 B.n393 163.367
R1656 B.n835 B.n387 163.367
R1657 B.n844 B.n387 163.367
R1658 B.n844 B.n385 163.367
R1659 B.n848 B.n385 163.367
R1660 B.n848 B.n2 163.367
R1661 B.n951 B.n2 163.367
R1662 B.n951 B.n3 163.367
R1663 B.n947 B.n3 163.367
R1664 B.n947 B.n9 163.367
R1665 B.n943 B.n9 163.367
R1666 B.n943 B.n11 163.367
R1667 B.n939 B.n11 163.367
R1668 B.n939 B.n16 163.367
R1669 B.n935 B.n16 163.367
R1670 B.n935 B.n18 163.367
R1671 B.n931 B.n18 163.367
R1672 B.n931 B.n23 163.367
R1673 B.n927 B.n23 163.367
R1674 B.n927 B.n25 163.367
R1675 B.n923 B.n25 163.367
R1676 B.n923 B.n29 163.367
R1677 B.n919 B.n29 163.367
R1678 B.n919 B.n31 163.367
R1679 B.n915 B.n31 163.367
R1680 B.n915 B.n37 163.367
R1681 B.n911 B.n37 163.367
R1682 B.n911 B.n39 163.367
R1683 B.n907 B.n39 163.367
R1684 B.n907 B.n44 163.367
R1685 B.n903 B.n44 163.367
R1686 B.n903 B.n46 163.367
R1687 B.n899 B.n46 163.367
R1688 B.n899 B.n51 163.367
R1689 B.n895 B.n51 163.367
R1690 B.n895 B.n53 163.367
R1691 B.n502 B.n501 163.367
R1692 B.n755 B.n501 163.367
R1693 B.n753 B.n752 163.367
R1694 B.n749 B.n748 163.367
R1695 B.n745 B.n744 163.367
R1696 B.n741 B.n740 163.367
R1697 B.n737 B.n736 163.367
R1698 B.n733 B.n732 163.367
R1699 B.n729 B.n728 163.367
R1700 B.n725 B.n724 163.367
R1701 B.n721 B.n720 163.367
R1702 B.n717 B.n716 163.367
R1703 B.n713 B.n712 163.367
R1704 B.n709 B.n708 163.367
R1705 B.n705 B.n704 163.367
R1706 B.n701 B.n700 163.367
R1707 B.n697 B.n696 163.367
R1708 B.n693 B.n692 163.367
R1709 B.n689 B.n688 163.367
R1710 B.n685 B.n684 163.367
R1711 B.n681 B.n680 163.367
R1712 B.n677 B.n676 163.367
R1713 B.n673 B.n672 163.367
R1714 B.n669 B.n668 163.367
R1715 B.n665 B.n664 163.367
R1716 B.n661 B.n660 163.367
R1717 B.n657 B.n656 163.367
R1718 B.n653 B.n652 163.367
R1719 B.n649 B.n648 163.367
R1720 B.n645 B.n644 163.367
R1721 B.n640 B.n639 163.367
R1722 B.n636 B.n635 163.367
R1723 B.n632 B.n631 163.367
R1724 B.n628 B.n627 163.367
R1725 B.n624 B.n623 163.367
R1726 B.n620 B.n619 163.367
R1727 B.n616 B.n615 163.367
R1728 B.n612 B.n611 163.367
R1729 B.n608 B.n607 163.367
R1730 B.n604 B.n603 163.367
R1731 B.n600 B.n599 163.367
R1732 B.n596 B.n595 163.367
R1733 B.n592 B.n591 163.367
R1734 B.n588 B.n587 163.367
R1735 B.n584 B.n583 163.367
R1736 B.n580 B.n579 163.367
R1737 B.n576 B.n575 163.367
R1738 B.n572 B.n571 163.367
R1739 B.n568 B.n567 163.367
R1740 B.n564 B.n563 163.367
R1741 B.n560 B.n559 163.367
R1742 B.n556 B.n555 163.367
R1743 B.n552 B.n551 163.367
R1744 B.n548 B.n547 163.367
R1745 B.n544 B.n543 163.367
R1746 B.n540 B.n539 163.367
R1747 B.n536 B.n535 163.367
R1748 B.n532 B.n531 163.367
R1749 B.n528 B.n527 163.367
R1750 B.n524 B.n523 163.367
R1751 B.n520 B.n519 163.367
R1752 B.n516 B.n515 163.367
R1753 B.n512 B.n511 163.367
R1754 B.n508 B.n438 163.367
R1755 B.n768 B.n436 163.367
R1756 B.n768 B.n430 163.367
R1757 B.n776 B.n430 163.367
R1758 B.n776 B.n428 163.367
R1759 B.n780 B.n428 163.367
R1760 B.n780 B.n422 163.367
R1761 B.n788 B.n422 163.367
R1762 B.n788 B.n420 163.367
R1763 B.n792 B.n420 163.367
R1764 B.n792 B.n414 163.367
R1765 B.n800 B.n414 163.367
R1766 B.n800 B.n412 163.367
R1767 B.n804 B.n412 163.367
R1768 B.n804 B.n407 163.367
R1769 B.n813 B.n407 163.367
R1770 B.n813 B.n405 163.367
R1771 B.n817 B.n405 163.367
R1772 B.n817 B.n399 163.367
R1773 B.n825 B.n399 163.367
R1774 B.n825 B.n397 163.367
R1775 B.n829 B.n397 163.367
R1776 B.n829 B.n390 163.367
R1777 B.n837 B.n390 163.367
R1778 B.n837 B.n388 163.367
R1779 B.n842 B.n388 163.367
R1780 B.n842 B.n383 163.367
R1781 B.n850 B.n383 163.367
R1782 B.n851 B.n850 163.367
R1783 B.n851 B.n5 163.367
R1784 B.n6 B.n5 163.367
R1785 B.n7 B.n6 163.367
R1786 B.n856 B.n7 163.367
R1787 B.n856 B.n12 163.367
R1788 B.n13 B.n12 163.367
R1789 B.n14 B.n13 163.367
R1790 B.n861 B.n14 163.367
R1791 B.n861 B.n19 163.367
R1792 B.n20 B.n19 163.367
R1793 B.n21 B.n20 163.367
R1794 B.n866 B.n21 163.367
R1795 B.n866 B.n26 163.367
R1796 B.n27 B.n26 163.367
R1797 B.n28 B.n27 163.367
R1798 B.n871 B.n28 163.367
R1799 B.n871 B.n33 163.367
R1800 B.n34 B.n33 163.367
R1801 B.n35 B.n34 163.367
R1802 B.n876 B.n35 163.367
R1803 B.n876 B.n40 163.367
R1804 B.n41 B.n40 163.367
R1805 B.n42 B.n41 163.367
R1806 B.n881 B.n42 163.367
R1807 B.n881 B.n47 163.367
R1808 B.n48 B.n47 163.367
R1809 B.n49 B.n48 163.367
R1810 B.n886 B.n49 163.367
R1811 B.n886 B.n54 163.367
R1812 B.n55 B.n54 163.367
R1813 B.n130 B.n129 163.367
R1814 B.n134 B.n133 163.367
R1815 B.n138 B.n137 163.367
R1816 B.n142 B.n141 163.367
R1817 B.n146 B.n145 163.367
R1818 B.n150 B.n149 163.367
R1819 B.n154 B.n153 163.367
R1820 B.n158 B.n157 163.367
R1821 B.n162 B.n161 163.367
R1822 B.n166 B.n165 163.367
R1823 B.n170 B.n169 163.367
R1824 B.n174 B.n173 163.367
R1825 B.n178 B.n177 163.367
R1826 B.n182 B.n181 163.367
R1827 B.n186 B.n185 163.367
R1828 B.n190 B.n189 163.367
R1829 B.n194 B.n193 163.367
R1830 B.n198 B.n197 163.367
R1831 B.n202 B.n201 163.367
R1832 B.n206 B.n205 163.367
R1833 B.n210 B.n209 163.367
R1834 B.n214 B.n213 163.367
R1835 B.n218 B.n217 163.367
R1836 B.n222 B.n221 163.367
R1837 B.n226 B.n225 163.367
R1838 B.n230 B.n229 163.367
R1839 B.n234 B.n233 163.367
R1840 B.n238 B.n237 163.367
R1841 B.n242 B.n241 163.367
R1842 B.n246 B.n245 163.367
R1843 B.n250 B.n249 163.367
R1844 B.n254 B.n253 163.367
R1845 B.n258 B.n257 163.367
R1846 B.n262 B.n261 163.367
R1847 B.n267 B.n266 163.367
R1848 B.n271 B.n270 163.367
R1849 B.n275 B.n274 163.367
R1850 B.n279 B.n278 163.367
R1851 B.n283 B.n282 163.367
R1852 B.n287 B.n286 163.367
R1853 B.n291 B.n290 163.367
R1854 B.n295 B.n294 163.367
R1855 B.n299 B.n298 163.367
R1856 B.n303 B.n302 163.367
R1857 B.n307 B.n306 163.367
R1858 B.n311 B.n310 163.367
R1859 B.n315 B.n314 163.367
R1860 B.n319 B.n318 163.367
R1861 B.n323 B.n322 163.367
R1862 B.n327 B.n326 163.367
R1863 B.n331 B.n330 163.367
R1864 B.n335 B.n334 163.367
R1865 B.n339 B.n338 163.367
R1866 B.n343 B.n342 163.367
R1867 B.n347 B.n346 163.367
R1868 B.n351 B.n350 163.367
R1869 B.n355 B.n354 163.367
R1870 B.n359 B.n358 163.367
R1871 B.n363 B.n362 163.367
R1872 B.n367 B.n366 163.367
R1873 B.n371 B.n370 163.367
R1874 B.n375 B.n374 163.367
R1875 B.n379 B.n378 163.367
R1876 B.n891 B.n120 163.367
R1877 B.n761 B.n760 71.676
R1878 B.n755 B.n439 71.676
R1879 B.n752 B.n440 71.676
R1880 B.n748 B.n441 71.676
R1881 B.n744 B.n442 71.676
R1882 B.n740 B.n443 71.676
R1883 B.n736 B.n444 71.676
R1884 B.n732 B.n445 71.676
R1885 B.n728 B.n446 71.676
R1886 B.n724 B.n447 71.676
R1887 B.n720 B.n448 71.676
R1888 B.n716 B.n449 71.676
R1889 B.n712 B.n450 71.676
R1890 B.n708 B.n451 71.676
R1891 B.n704 B.n452 71.676
R1892 B.n700 B.n453 71.676
R1893 B.n696 B.n454 71.676
R1894 B.n692 B.n455 71.676
R1895 B.n688 B.n456 71.676
R1896 B.n684 B.n457 71.676
R1897 B.n680 B.n458 71.676
R1898 B.n676 B.n459 71.676
R1899 B.n672 B.n460 71.676
R1900 B.n668 B.n461 71.676
R1901 B.n664 B.n462 71.676
R1902 B.n660 B.n463 71.676
R1903 B.n656 B.n464 71.676
R1904 B.n652 B.n465 71.676
R1905 B.n648 B.n466 71.676
R1906 B.n644 B.n467 71.676
R1907 B.n639 B.n468 71.676
R1908 B.n635 B.n469 71.676
R1909 B.n631 B.n470 71.676
R1910 B.n627 B.n471 71.676
R1911 B.n623 B.n472 71.676
R1912 B.n619 B.n473 71.676
R1913 B.n615 B.n474 71.676
R1914 B.n611 B.n475 71.676
R1915 B.n607 B.n476 71.676
R1916 B.n603 B.n477 71.676
R1917 B.n599 B.n478 71.676
R1918 B.n595 B.n479 71.676
R1919 B.n591 B.n480 71.676
R1920 B.n587 B.n481 71.676
R1921 B.n583 B.n482 71.676
R1922 B.n579 B.n483 71.676
R1923 B.n575 B.n484 71.676
R1924 B.n571 B.n485 71.676
R1925 B.n567 B.n486 71.676
R1926 B.n563 B.n487 71.676
R1927 B.n559 B.n488 71.676
R1928 B.n555 B.n489 71.676
R1929 B.n551 B.n490 71.676
R1930 B.n547 B.n491 71.676
R1931 B.n543 B.n492 71.676
R1932 B.n539 B.n493 71.676
R1933 B.n535 B.n494 71.676
R1934 B.n531 B.n495 71.676
R1935 B.n527 B.n496 71.676
R1936 B.n523 B.n497 71.676
R1937 B.n519 B.n498 71.676
R1938 B.n515 B.n499 71.676
R1939 B.n511 B.n500 71.676
R1940 B.n763 B.n438 71.676
R1941 B.n126 B.n56 71.676
R1942 B.n130 B.n57 71.676
R1943 B.n134 B.n58 71.676
R1944 B.n138 B.n59 71.676
R1945 B.n142 B.n60 71.676
R1946 B.n146 B.n61 71.676
R1947 B.n150 B.n62 71.676
R1948 B.n154 B.n63 71.676
R1949 B.n158 B.n64 71.676
R1950 B.n162 B.n65 71.676
R1951 B.n166 B.n66 71.676
R1952 B.n170 B.n67 71.676
R1953 B.n174 B.n68 71.676
R1954 B.n178 B.n69 71.676
R1955 B.n182 B.n70 71.676
R1956 B.n186 B.n71 71.676
R1957 B.n190 B.n72 71.676
R1958 B.n194 B.n73 71.676
R1959 B.n198 B.n74 71.676
R1960 B.n202 B.n75 71.676
R1961 B.n206 B.n76 71.676
R1962 B.n210 B.n77 71.676
R1963 B.n214 B.n78 71.676
R1964 B.n218 B.n79 71.676
R1965 B.n222 B.n80 71.676
R1966 B.n226 B.n81 71.676
R1967 B.n230 B.n82 71.676
R1968 B.n234 B.n83 71.676
R1969 B.n238 B.n84 71.676
R1970 B.n242 B.n85 71.676
R1971 B.n246 B.n86 71.676
R1972 B.n250 B.n87 71.676
R1973 B.n254 B.n88 71.676
R1974 B.n258 B.n89 71.676
R1975 B.n262 B.n90 71.676
R1976 B.n267 B.n91 71.676
R1977 B.n271 B.n92 71.676
R1978 B.n275 B.n93 71.676
R1979 B.n279 B.n94 71.676
R1980 B.n283 B.n95 71.676
R1981 B.n287 B.n96 71.676
R1982 B.n291 B.n97 71.676
R1983 B.n295 B.n98 71.676
R1984 B.n299 B.n99 71.676
R1985 B.n303 B.n100 71.676
R1986 B.n307 B.n101 71.676
R1987 B.n311 B.n102 71.676
R1988 B.n315 B.n103 71.676
R1989 B.n319 B.n104 71.676
R1990 B.n323 B.n105 71.676
R1991 B.n327 B.n106 71.676
R1992 B.n331 B.n107 71.676
R1993 B.n335 B.n108 71.676
R1994 B.n339 B.n109 71.676
R1995 B.n343 B.n110 71.676
R1996 B.n347 B.n111 71.676
R1997 B.n351 B.n112 71.676
R1998 B.n355 B.n113 71.676
R1999 B.n359 B.n114 71.676
R2000 B.n363 B.n115 71.676
R2001 B.n367 B.n116 71.676
R2002 B.n371 B.n117 71.676
R2003 B.n375 B.n118 71.676
R2004 B.n379 B.n119 71.676
R2005 B.n120 B.n119 71.676
R2006 B.n378 B.n118 71.676
R2007 B.n374 B.n117 71.676
R2008 B.n370 B.n116 71.676
R2009 B.n366 B.n115 71.676
R2010 B.n362 B.n114 71.676
R2011 B.n358 B.n113 71.676
R2012 B.n354 B.n112 71.676
R2013 B.n350 B.n111 71.676
R2014 B.n346 B.n110 71.676
R2015 B.n342 B.n109 71.676
R2016 B.n338 B.n108 71.676
R2017 B.n334 B.n107 71.676
R2018 B.n330 B.n106 71.676
R2019 B.n326 B.n105 71.676
R2020 B.n322 B.n104 71.676
R2021 B.n318 B.n103 71.676
R2022 B.n314 B.n102 71.676
R2023 B.n310 B.n101 71.676
R2024 B.n306 B.n100 71.676
R2025 B.n302 B.n99 71.676
R2026 B.n298 B.n98 71.676
R2027 B.n294 B.n97 71.676
R2028 B.n290 B.n96 71.676
R2029 B.n286 B.n95 71.676
R2030 B.n282 B.n94 71.676
R2031 B.n278 B.n93 71.676
R2032 B.n274 B.n92 71.676
R2033 B.n270 B.n91 71.676
R2034 B.n266 B.n90 71.676
R2035 B.n261 B.n89 71.676
R2036 B.n257 B.n88 71.676
R2037 B.n253 B.n87 71.676
R2038 B.n249 B.n86 71.676
R2039 B.n245 B.n85 71.676
R2040 B.n241 B.n84 71.676
R2041 B.n237 B.n83 71.676
R2042 B.n233 B.n82 71.676
R2043 B.n229 B.n81 71.676
R2044 B.n225 B.n80 71.676
R2045 B.n221 B.n79 71.676
R2046 B.n217 B.n78 71.676
R2047 B.n213 B.n77 71.676
R2048 B.n209 B.n76 71.676
R2049 B.n205 B.n75 71.676
R2050 B.n201 B.n74 71.676
R2051 B.n197 B.n73 71.676
R2052 B.n193 B.n72 71.676
R2053 B.n189 B.n71 71.676
R2054 B.n185 B.n70 71.676
R2055 B.n181 B.n69 71.676
R2056 B.n177 B.n68 71.676
R2057 B.n173 B.n67 71.676
R2058 B.n169 B.n66 71.676
R2059 B.n165 B.n65 71.676
R2060 B.n161 B.n64 71.676
R2061 B.n157 B.n63 71.676
R2062 B.n153 B.n62 71.676
R2063 B.n149 B.n61 71.676
R2064 B.n145 B.n60 71.676
R2065 B.n141 B.n59 71.676
R2066 B.n137 B.n58 71.676
R2067 B.n133 B.n57 71.676
R2068 B.n129 B.n56 71.676
R2069 B.n761 B.n502 71.676
R2070 B.n753 B.n439 71.676
R2071 B.n749 B.n440 71.676
R2072 B.n745 B.n441 71.676
R2073 B.n741 B.n442 71.676
R2074 B.n737 B.n443 71.676
R2075 B.n733 B.n444 71.676
R2076 B.n729 B.n445 71.676
R2077 B.n725 B.n446 71.676
R2078 B.n721 B.n447 71.676
R2079 B.n717 B.n448 71.676
R2080 B.n713 B.n449 71.676
R2081 B.n709 B.n450 71.676
R2082 B.n705 B.n451 71.676
R2083 B.n701 B.n452 71.676
R2084 B.n697 B.n453 71.676
R2085 B.n693 B.n454 71.676
R2086 B.n689 B.n455 71.676
R2087 B.n685 B.n456 71.676
R2088 B.n681 B.n457 71.676
R2089 B.n677 B.n458 71.676
R2090 B.n673 B.n459 71.676
R2091 B.n669 B.n460 71.676
R2092 B.n665 B.n461 71.676
R2093 B.n661 B.n462 71.676
R2094 B.n657 B.n463 71.676
R2095 B.n653 B.n464 71.676
R2096 B.n649 B.n465 71.676
R2097 B.n645 B.n466 71.676
R2098 B.n640 B.n467 71.676
R2099 B.n636 B.n468 71.676
R2100 B.n632 B.n469 71.676
R2101 B.n628 B.n470 71.676
R2102 B.n624 B.n471 71.676
R2103 B.n620 B.n472 71.676
R2104 B.n616 B.n473 71.676
R2105 B.n612 B.n474 71.676
R2106 B.n608 B.n475 71.676
R2107 B.n604 B.n476 71.676
R2108 B.n600 B.n477 71.676
R2109 B.n596 B.n478 71.676
R2110 B.n592 B.n479 71.676
R2111 B.n588 B.n480 71.676
R2112 B.n584 B.n481 71.676
R2113 B.n580 B.n482 71.676
R2114 B.n576 B.n483 71.676
R2115 B.n572 B.n484 71.676
R2116 B.n568 B.n485 71.676
R2117 B.n564 B.n486 71.676
R2118 B.n560 B.n487 71.676
R2119 B.n556 B.n488 71.676
R2120 B.n552 B.n489 71.676
R2121 B.n548 B.n490 71.676
R2122 B.n544 B.n491 71.676
R2123 B.n540 B.n492 71.676
R2124 B.n536 B.n493 71.676
R2125 B.n532 B.n494 71.676
R2126 B.n528 B.n495 71.676
R2127 B.n524 B.n496 71.676
R2128 B.n520 B.n497 71.676
R2129 B.n516 B.n498 71.676
R2130 B.n512 B.n499 71.676
R2131 B.n508 B.n500 71.676
R2132 B.n764 B.n763 71.676
R2133 B.n507 B.n506 59.5399
R2134 B.n642 B.n504 59.5399
R2135 B.n125 B.n124 59.5399
R2136 B.n264 B.n122 59.5399
R2137 B.n762 B.n435 55.8571
R2138 B.n893 B.n892 55.8571
R2139 B.n506 B.n505 34.3278
R2140 B.n504 B.n503 34.3278
R2141 B.n124 B.n123 34.3278
R2142 B.n122 B.n121 34.3278
R2143 B.n127 B.n52 32.0005
R2144 B.n890 B.n889 32.0005
R2145 B.n766 B.n765 32.0005
R2146 B.n759 B.n433 32.0005
R2147 B.n769 B.n435 31.9186
R2148 B.n769 B.n431 31.9186
R2149 B.n775 B.n431 31.9186
R2150 B.n775 B.n427 31.9186
R2151 B.n781 B.n427 31.9186
R2152 B.n787 B.n423 31.9186
R2153 B.n787 B.n419 31.9186
R2154 B.n793 B.n419 31.9186
R2155 B.n793 B.n415 31.9186
R2156 B.n799 B.n415 31.9186
R2157 B.n799 B.n411 31.9186
R2158 B.n806 B.n411 31.9186
R2159 B.n806 B.n805 31.9186
R2160 B.n812 B.n404 31.9186
R2161 B.n818 B.n404 31.9186
R2162 B.n818 B.n400 31.9186
R2163 B.n824 B.n400 31.9186
R2164 B.n830 B.n396 31.9186
R2165 B.n830 B.n391 31.9186
R2166 B.n836 B.n391 31.9186
R2167 B.n836 B.n392 31.9186
R2168 B.n843 B.n384 31.9186
R2169 B.n849 B.n384 31.9186
R2170 B.n849 B.n4 31.9186
R2171 B.n950 B.n4 31.9186
R2172 B.n950 B.n949 31.9186
R2173 B.n949 B.n948 31.9186
R2174 B.n948 B.n8 31.9186
R2175 B.n942 B.n8 31.9186
R2176 B.n941 B.n940 31.9186
R2177 B.n940 B.n15 31.9186
R2178 B.n934 B.n15 31.9186
R2179 B.n934 B.n933 31.9186
R2180 B.n932 B.n22 31.9186
R2181 B.n926 B.n22 31.9186
R2182 B.n926 B.n925 31.9186
R2183 B.n925 B.n924 31.9186
R2184 B.n918 B.n32 31.9186
R2185 B.n918 B.n917 31.9186
R2186 B.n917 B.n916 31.9186
R2187 B.n916 B.n36 31.9186
R2188 B.n910 B.n36 31.9186
R2189 B.n910 B.n909 31.9186
R2190 B.n909 B.n908 31.9186
R2191 B.n908 B.n43 31.9186
R2192 B.n902 B.n901 31.9186
R2193 B.n901 B.n900 31.9186
R2194 B.n900 B.n50 31.9186
R2195 B.n894 B.n50 31.9186
R2196 B.n894 B.n893 31.9186
R2197 B.n781 B.t7 30.9798
R2198 B.n902 B.t14 30.9798
R2199 B.n392 B.t3 25.3472
R2200 B.t2 B.n941 25.3472
R2201 B.n812 B.t1 19.7146
R2202 B.n924 B.t5 19.7146
R2203 B.n824 B.t4 18.7758
R2204 B.t0 B.n932 18.7758
R2205 B B.n952 18.0485
R2206 B.t4 B.n396 13.1432
R2207 B.n933 B.t0 13.1432
R2208 B.n805 B.t1 12.2045
R2209 B.n32 B.t5 12.2045
R2210 B.n128 B.n127 10.6151
R2211 B.n131 B.n128 10.6151
R2212 B.n132 B.n131 10.6151
R2213 B.n135 B.n132 10.6151
R2214 B.n136 B.n135 10.6151
R2215 B.n139 B.n136 10.6151
R2216 B.n140 B.n139 10.6151
R2217 B.n143 B.n140 10.6151
R2218 B.n144 B.n143 10.6151
R2219 B.n147 B.n144 10.6151
R2220 B.n148 B.n147 10.6151
R2221 B.n151 B.n148 10.6151
R2222 B.n152 B.n151 10.6151
R2223 B.n155 B.n152 10.6151
R2224 B.n156 B.n155 10.6151
R2225 B.n159 B.n156 10.6151
R2226 B.n160 B.n159 10.6151
R2227 B.n163 B.n160 10.6151
R2228 B.n164 B.n163 10.6151
R2229 B.n167 B.n164 10.6151
R2230 B.n168 B.n167 10.6151
R2231 B.n171 B.n168 10.6151
R2232 B.n172 B.n171 10.6151
R2233 B.n175 B.n172 10.6151
R2234 B.n176 B.n175 10.6151
R2235 B.n179 B.n176 10.6151
R2236 B.n180 B.n179 10.6151
R2237 B.n183 B.n180 10.6151
R2238 B.n184 B.n183 10.6151
R2239 B.n187 B.n184 10.6151
R2240 B.n188 B.n187 10.6151
R2241 B.n191 B.n188 10.6151
R2242 B.n192 B.n191 10.6151
R2243 B.n195 B.n192 10.6151
R2244 B.n196 B.n195 10.6151
R2245 B.n199 B.n196 10.6151
R2246 B.n200 B.n199 10.6151
R2247 B.n203 B.n200 10.6151
R2248 B.n204 B.n203 10.6151
R2249 B.n207 B.n204 10.6151
R2250 B.n208 B.n207 10.6151
R2251 B.n211 B.n208 10.6151
R2252 B.n212 B.n211 10.6151
R2253 B.n215 B.n212 10.6151
R2254 B.n216 B.n215 10.6151
R2255 B.n219 B.n216 10.6151
R2256 B.n220 B.n219 10.6151
R2257 B.n223 B.n220 10.6151
R2258 B.n224 B.n223 10.6151
R2259 B.n227 B.n224 10.6151
R2260 B.n228 B.n227 10.6151
R2261 B.n231 B.n228 10.6151
R2262 B.n232 B.n231 10.6151
R2263 B.n235 B.n232 10.6151
R2264 B.n236 B.n235 10.6151
R2265 B.n239 B.n236 10.6151
R2266 B.n240 B.n239 10.6151
R2267 B.n243 B.n240 10.6151
R2268 B.n244 B.n243 10.6151
R2269 B.n248 B.n247 10.6151
R2270 B.n251 B.n248 10.6151
R2271 B.n252 B.n251 10.6151
R2272 B.n255 B.n252 10.6151
R2273 B.n256 B.n255 10.6151
R2274 B.n259 B.n256 10.6151
R2275 B.n260 B.n259 10.6151
R2276 B.n263 B.n260 10.6151
R2277 B.n268 B.n265 10.6151
R2278 B.n269 B.n268 10.6151
R2279 B.n272 B.n269 10.6151
R2280 B.n273 B.n272 10.6151
R2281 B.n276 B.n273 10.6151
R2282 B.n277 B.n276 10.6151
R2283 B.n280 B.n277 10.6151
R2284 B.n281 B.n280 10.6151
R2285 B.n284 B.n281 10.6151
R2286 B.n285 B.n284 10.6151
R2287 B.n288 B.n285 10.6151
R2288 B.n289 B.n288 10.6151
R2289 B.n292 B.n289 10.6151
R2290 B.n293 B.n292 10.6151
R2291 B.n296 B.n293 10.6151
R2292 B.n297 B.n296 10.6151
R2293 B.n300 B.n297 10.6151
R2294 B.n301 B.n300 10.6151
R2295 B.n304 B.n301 10.6151
R2296 B.n305 B.n304 10.6151
R2297 B.n308 B.n305 10.6151
R2298 B.n309 B.n308 10.6151
R2299 B.n312 B.n309 10.6151
R2300 B.n313 B.n312 10.6151
R2301 B.n316 B.n313 10.6151
R2302 B.n317 B.n316 10.6151
R2303 B.n320 B.n317 10.6151
R2304 B.n321 B.n320 10.6151
R2305 B.n324 B.n321 10.6151
R2306 B.n325 B.n324 10.6151
R2307 B.n328 B.n325 10.6151
R2308 B.n329 B.n328 10.6151
R2309 B.n332 B.n329 10.6151
R2310 B.n333 B.n332 10.6151
R2311 B.n336 B.n333 10.6151
R2312 B.n337 B.n336 10.6151
R2313 B.n340 B.n337 10.6151
R2314 B.n341 B.n340 10.6151
R2315 B.n344 B.n341 10.6151
R2316 B.n345 B.n344 10.6151
R2317 B.n348 B.n345 10.6151
R2318 B.n349 B.n348 10.6151
R2319 B.n352 B.n349 10.6151
R2320 B.n353 B.n352 10.6151
R2321 B.n356 B.n353 10.6151
R2322 B.n357 B.n356 10.6151
R2323 B.n360 B.n357 10.6151
R2324 B.n361 B.n360 10.6151
R2325 B.n364 B.n361 10.6151
R2326 B.n365 B.n364 10.6151
R2327 B.n368 B.n365 10.6151
R2328 B.n369 B.n368 10.6151
R2329 B.n372 B.n369 10.6151
R2330 B.n373 B.n372 10.6151
R2331 B.n376 B.n373 10.6151
R2332 B.n377 B.n376 10.6151
R2333 B.n380 B.n377 10.6151
R2334 B.n381 B.n380 10.6151
R2335 B.n890 B.n381 10.6151
R2336 B.n767 B.n766 10.6151
R2337 B.n767 B.n429 10.6151
R2338 B.n777 B.n429 10.6151
R2339 B.n778 B.n777 10.6151
R2340 B.n779 B.n778 10.6151
R2341 B.n779 B.n421 10.6151
R2342 B.n789 B.n421 10.6151
R2343 B.n790 B.n789 10.6151
R2344 B.n791 B.n790 10.6151
R2345 B.n791 B.n413 10.6151
R2346 B.n801 B.n413 10.6151
R2347 B.n802 B.n801 10.6151
R2348 B.n803 B.n802 10.6151
R2349 B.n803 B.n406 10.6151
R2350 B.n814 B.n406 10.6151
R2351 B.n815 B.n814 10.6151
R2352 B.n816 B.n815 10.6151
R2353 B.n816 B.n398 10.6151
R2354 B.n826 B.n398 10.6151
R2355 B.n827 B.n826 10.6151
R2356 B.n828 B.n827 10.6151
R2357 B.n828 B.n389 10.6151
R2358 B.n838 B.n389 10.6151
R2359 B.n839 B.n838 10.6151
R2360 B.n841 B.n839 10.6151
R2361 B.n841 B.n840 10.6151
R2362 B.n840 B.n382 10.6151
R2363 B.n852 B.n382 10.6151
R2364 B.n853 B.n852 10.6151
R2365 B.n854 B.n853 10.6151
R2366 B.n855 B.n854 10.6151
R2367 B.n857 B.n855 10.6151
R2368 B.n858 B.n857 10.6151
R2369 B.n859 B.n858 10.6151
R2370 B.n860 B.n859 10.6151
R2371 B.n862 B.n860 10.6151
R2372 B.n863 B.n862 10.6151
R2373 B.n864 B.n863 10.6151
R2374 B.n865 B.n864 10.6151
R2375 B.n867 B.n865 10.6151
R2376 B.n868 B.n867 10.6151
R2377 B.n869 B.n868 10.6151
R2378 B.n870 B.n869 10.6151
R2379 B.n872 B.n870 10.6151
R2380 B.n873 B.n872 10.6151
R2381 B.n874 B.n873 10.6151
R2382 B.n875 B.n874 10.6151
R2383 B.n877 B.n875 10.6151
R2384 B.n878 B.n877 10.6151
R2385 B.n879 B.n878 10.6151
R2386 B.n880 B.n879 10.6151
R2387 B.n882 B.n880 10.6151
R2388 B.n883 B.n882 10.6151
R2389 B.n884 B.n883 10.6151
R2390 B.n885 B.n884 10.6151
R2391 B.n887 B.n885 10.6151
R2392 B.n888 B.n887 10.6151
R2393 B.n889 B.n888 10.6151
R2394 B.n759 B.n758 10.6151
R2395 B.n758 B.n757 10.6151
R2396 B.n757 B.n756 10.6151
R2397 B.n756 B.n754 10.6151
R2398 B.n754 B.n751 10.6151
R2399 B.n751 B.n750 10.6151
R2400 B.n750 B.n747 10.6151
R2401 B.n747 B.n746 10.6151
R2402 B.n746 B.n743 10.6151
R2403 B.n743 B.n742 10.6151
R2404 B.n742 B.n739 10.6151
R2405 B.n739 B.n738 10.6151
R2406 B.n738 B.n735 10.6151
R2407 B.n735 B.n734 10.6151
R2408 B.n734 B.n731 10.6151
R2409 B.n731 B.n730 10.6151
R2410 B.n730 B.n727 10.6151
R2411 B.n727 B.n726 10.6151
R2412 B.n726 B.n723 10.6151
R2413 B.n723 B.n722 10.6151
R2414 B.n722 B.n719 10.6151
R2415 B.n719 B.n718 10.6151
R2416 B.n718 B.n715 10.6151
R2417 B.n715 B.n714 10.6151
R2418 B.n714 B.n711 10.6151
R2419 B.n711 B.n710 10.6151
R2420 B.n710 B.n707 10.6151
R2421 B.n707 B.n706 10.6151
R2422 B.n706 B.n703 10.6151
R2423 B.n703 B.n702 10.6151
R2424 B.n702 B.n699 10.6151
R2425 B.n699 B.n698 10.6151
R2426 B.n698 B.n695 10.6151
R2427 B.n695 B.n694 10.6151
R2428 B.n694 B.n691 10.6151
R2429 B.n691 B.n690 10.6151
R2430 B.n690 B.n687 10.6151
R2431 B.n687 B.n686 10.6151
R2432 B.n686 B.n683 10.6151
R2433 B.n683 B.n682 10.6151
R2434 B.n682 B.n679 10.6151
R2435 B.n679 B.n678 10.6151
R2436 B.n678 B.n675 10.6151
R2437 B.n675 B.n674 10.6151
R2438 B.n674 B.n671 10.6151
R2439 B.n671 B.n670 10.6151
R2440 B.n670 B.n667 10.6151
R2441 B.n667 B.n666 10.6151
R2442 B.n666 B.n663 10.6151
R2443 B.n663 B.n662 10.6151
R2444 B.n662 B.n659 10.6151
R2445 B.n659 B.n658 10.6151
R2446 B.n658 B.n655 10.6151
R2447 B.n655 B.n654 10.6151
R2448 B.n654 B.n651 10.6151
R2449 B.n651 B.n650 10.6151
R2450 B.n650 B.n647 10.6151
R2451 B.n647 B.n646 10.6151
R2452 B.n646 B.n643 10.6151
R2453 B.n641 B.n638 10.6151
R2454 B.n638 B.n637 10.6151
R2455 B.n637 B.n634 10.6151
R2456 B.n634 B.n633 10.6151
R2457 B.n633 B.n630 10.6151
R2458 B.n630 B.n629 10.6151
R2459 B.n629 B.n626 10.6151
R2460 B.n626 B.n625 10.6151
R2461 B.n622 B.n621 10.6151
R2462 B.n621 B.n618 10.6151
R2463 B.n618 B.n617 10.6151
R2464 B.n617 B.n614 10.6151
R2465 B.n614 B.n613 10.6151
R2466 B.n613 B.n610 10.6151
R2467 B.n610 B.n609 10.6151
R2468 B.n609 B.n606 10.6151
R2469 B.n606 B.n605 10.6151
R2470 B.n605 B.n602 10.6151
R2471 B.n602 B.n601 10.6151
R2472 B.n601 B.n598 10.6151
R2473 B.n598 B.n597 10.6151
R2474 B.n597 B.n594 10.6151
R2475 B.n594 B.n593 10.6151
R2476 B.n593 B.n590 10.6151
R2477 B.n590 B.n589 10.6151
R2478 B.n589 B.n586 10.6151
R2479 B.n586 B.n585 10.6151
R2480 B.n585 B.n582 10.6151
R2481 B.n582 B.n581 10.6151
R2482 B.n581 B.n578 10.6151
R2483 B.n578 B.n577 10.6151
R2484 B.n577 B.n574 10.6151
R2485 B.n574 B.n573 10.6151
R2486 B.n573 B.n570 10.6151
R2487 B.n570 B.n569 10.6151
R2488 B.n569 B.n566 10.6151
R2489 B.n566 B.n565 10.6151
R2490 B.n565 B.n562 10.6151
R2491 B.n562 B.n561 10.6151
R2492 B.n561 B.n558 10.6151
R2493 B.n558 B.n557 10.6151
R2494 B.n557 B.n554 10.6151
R2495 B.n554 B.n553 10.6151
R2496 B.n553 B.n550 10.6151
R2497 B.n550 B.n549 10.6151
R2498 B.n549 B.n546 10.6151
R2499 B.n546 B.n545 10.6151
R2500 B.n545 B.n542 10.6151
R2501 B.n542 B.n541 10.6151
R2502 B.n541 B.n538 10.6151
R2503 B.n538 B.n537 10.6151
R2504 B.n537 B.n534 10.6151
R2505 B.n534 B.n533 10.6151
R2506 B.n533 B.n530 10.6151
R2507 B.n530 B.n529 10.6151
R2508 B.n529 B.n526 10.6151
R2509 B.n526 B.n525 10.6151
R2510 B.n525 B.n522 10.6151
R2511 B.n522 B.n521 10.6151
R2512 B.n521 B.n518 10.6151
R2513 B.n518 B.n517 10.6151
R2514 B.n517 B.n514 10.6151
R2515 B.n514 B.n513 10.6151
R2516 B.n513 B.n510 10.6151
R2517 B.n510 B.n509 10.6151
R2518 B.n509 B.n437 10.6151
R2519 B.n765 B.n437 10.6151
R2520 B.n771 B.n433 10.6151
R2521 B.n772 B.n771 10.6151
R2522 B.n773 B.n772 10.6151
R2523 B.n773 B.n425 10.6151
R2524 B.n783 B.n425 10.6151
R2525 B.n784 B.n783 10.6151
R2526 B.n785 B.n784 10.6151
R2527 B.n785 B.n417 10.6151
R2528 B.n795 B.n417 10.6151
R2529 B.n796 B.n795 10.6151
R2530 B.n797 B.n796 10.6151
R2531 B.n797 B.n409 10.6151
R2532 B.n808 B.n409 10.6151
R2533 B.n809 B.n808 10.6151
R2534 B.n810 B.n809 10.6151
R2535 B.n810 B.n402 10.6151
R2536 B.n820 B.n402 10.6151
R2537 B.n821 B.n820 10.6151
R2538 B.n822 B.n821 10.6151
R2539 B.n822 B.n394 10.6151
R2540 B.n832 B.n394 10.6151
R2541 B.n833 B.n832 10.6151
R2542 B.n834 B.n833 10.6151
R2543 B.n834 B.n386 10.6151
R2544 B.n845 B.n386 10.6151
R2545 B.n846 B.n845 10.6151
R2546 B.n847 B.n846 10.6151
R2547 B.n847 B.n0 10.6151
R2548 B.n946 B.n1 10.6151
R2549 B.n946 B.n945 10.6151
R2550 B.n945 B.n944 10.6151
R2551 B.n944 B.n10 10.6151
R2552 B.n938 B.n10 10.6151
R2553 B.n938 B.n937 10.6151
R2554 B.n937 B.n936 10.6151
R2555 B.n936 B.n17 10.6151
R2556 B.n930 B.n17 10.6151
R2557 B.n930 B.n929 10.6151
R2558 B.n929 B.n928 10.6151
R2559 B.n928 B.n24 10.6151
R2560 B.n922 B.n24 10.6151
R2561 B.n922 B.n921 10.6151
R2562 B.n921 B.n920 10.6151
R2563 B.n920 B.n30 10.6151
R2564 B.n914 B.n30 10.6151
R2565 B.n914 B.n913 10.6151
R2566 B.n913 B.n912 10.6151
R2567 B.n912 B.n38 10.6151
R2568 B.n906 B.n38 10.6151
R2569 B.n906 B.n905 10.6151
R2570 B.n905 B.n904 10.6151
R2571 B.n904 B.n45 10.6151
R2572 B.n898 B.n45 10.6151
R2573 B.n898 B.n897 10.6151
R2574 B.n897 B.n896 10.6151
R2575 B.n896 B.n52 10.6151
R2576 B.n843 B.t3 6.57187
R2577 B.n942 B.t2 6.57187
R2578 B.n247 B.n125 6.5566
R2579 B.n264 B.n263 6.5566
R2580 B.n642 B.n641 6.5566
R2581 B.n625 B.n507 6.5566
R2582 B.n244 B.n125 4.05904
R2583 B.n265 B.n264 4.05904
R2584 B.n643 B.n642 4.05904
R2585 B.n622 B.n507 4.05904
R2586 B.n952 B.n0 2.81026
R2587 B.n952 B.n1 2.81026
R2588 B.t7 B.n423 0.939267
R2589 B.t14 B.n43 0.939267
R2590 VN.n3 VN.t3 340.046
R2591 VN.n13 VN.t2 340.046
R2592 VN.n2 VN.t5 303.928
R2593 VN.n8 VN.t1 303.928
R2594 VN.n12 VN.t0 303.928
R2595 VN.n18 VN.t4 303.928
R2596 VN.n9 VN.n8 172.613
R2597 VN.n19 VN.n18 172.613
R2598 VN.n17 VN.n10 161.3
R2599 VN.n16 VN.n15 161.3
R2600 VN.n14 VN.n11 161.3
R2601 VN.n7 VN.n0 161.3
R2602 VN.n6 VN.n5 161.3
R2603 VN.n4 VN.n1 161.3
R2604 VN.n6 VN.n1 51.7179
R2605 VN.n16 VN.n11 51.7179
R2606 VN VN.n19 49.135
R2607 VN.n3 VN.n2 41.9337
R2608 VN.n13 VN.n12 41.9337
R2609 VN.n7 VN.n6 29.4362
R2610 VN.n17 VN.n16 29.4362
R2611 VN.n2 VN.n1 24.5923
R2612 VN.n12 VN.n11 24.5923
R2613 VN.n14 VN.n13 17.4039
R2614 VN.n4 VN.n3 17.4039
R2615 VN.n8 VN.n7 13.2801
R2616 VN.n18 VN.n17 13.2801
R2617 VN.n19 VN.n10 0.189894
R2618 VN.n15 VN.n10 0.189894
R2619 VN.n15 VN.n14 0.189894
R2620 VN.n5 VN.n4 0.189894
R2621 VN.n5 VN.n0 0.189894
R2622 VN.n9 VN.n0 0.189894
R2623 VN VN.n9 0.0516364
R2624 VDD2.n199 VDD2.n103 289.615
R2625 VDD2.n96 VDD2.n0 289.615
R2626 VDD2.n200 VDD2.n199 185
R2627 VDD2.n198 VDD2.n197 185
R2628 VDD2.n107 VDD2.n106 185
R2629 VDD2.n192 VDD2.n191 185
R2630 VDD2.n190 VDD2.n189 185
R2631 VDD2.n111 VDD2.n110 185
R2632 VDD2.n184 VDD2.n183 185
R2633 VDD2.n182 VDD2.n113 185
R2634 VDD2.n181 VDD2.n180 185
R2635 VDD2.n116 VDD2.n114 185
R2636 VDD2.n175 VDD2.n174 185
R2637 VDD2.n173 VDD2.n172 185
R2638 VDD2.n120 VDD2.n119 185
R2639 VDD2.n167 VDD2.n166 185
R2640 VDD2.n165 VDD2.n164 185
R2641 VDD2.n124 VDD2.n123 185
R2642 VDD2.n159 VDD2.n158 185
R2643 VDD2.n157 VDD2.n156 185
R2644 VDD2.n128 VDD2.n127 185
R2645 VDD2.n151 VDD2.n150 185
R2646 VDD2.n149 VDD2.n148 185
R2647 VDD2.n132 VDD2.n131 185
R2648 VDD2.n143 VDD2.n142 185
R2649 VDD2.n141 VDD2.n140 185
R2650 VDD2.n136 VDD2.n135 185
R2651 VDD2.n32 VDD2.n31 185
R2652 VDD2.n37 VDD2.n36 185
R2653 VDD2.n39 VDD2.n38 185
R2654 VDD2.n28 VDD2.n27 185
R2655 VDD2.n45 VDD2.n44 185
R2656 VDD2.n47 VDD2.n46 185
R2657 VDD2.n24 VDD2.n23 185
R2658 VDD2.n53 VDD2.n52 185
R2659 VDD2.n55 VDD2.n54 185
R2660 VDD2.n20 VDD2.n19 185
R2661 VDD2.n61 VDD2.n60 185
R2662 VDD2.n63 VDD2.n62 185
R2663 VDD2.n16 VDD2.n15 185
R2664 VDD2.n69 VDD2.n68 185
R2665 VDD2.n71 VDD2.n70 185
R2666 VDD2.n12 VDD2.n11 185
R2667 VDD2.n78 VDD2.n77 185
R2668 VDD2.n79 VDD2.n10 185
R2669 VDD2.n81 VDD2.n80 185
R2670 VDD2.n8 VDD2.n7 185
R2671 VDD2.n87 VDD2.n86 185
R2672 VDD2.n89 VDD2.n88 185
R2673 VDD2.n4 VDD2.n3 185
R2674 VDD2.n95 VDD2.n94 185
R2675 VDD2.n97 VDD2.n96 185
R2676 VDD2.n137 VDD2.t1 147.659
R2677 VDD2.n33 VDD2.t2 147.659
R2678 VDD2.n199 VDD2.n198 104.615
R2679 VDD2.n198 VDD2.n106 104.615
R2680 VDD2.n191 VDD2.n106 104.615
R2681 VDD2.n191 VDD2.n190 104.615
R2682 VDD2.n190 VDD2.n110 104.615
R2683 VDD2.n183 VDD2.n110 104.615
R2684 VDD2.n183 VDD2.n182 104.615
R2685 VDD2.n182 VDD2.n181 104.615
R2686 VDD2.n181 VDD2.n114 104.615
R2687 VDD2.n174 VDD2.n114 104.615
R2688 VDD2.n174 VDD2.n173 104.615
R2689 VDD2.n173 VDD2.n119 104.615
R2690 VDD2.n166 VDD2.n119 104.615
R2691 VDD2.n166 VDD2.n165 104.615
R2692 VDD2.n165 VDD2.n123 104.615
R2693 VDD2.n158 VDD2.n123 104.615
R2694 VDD2.n158 VDD2.n157 104.615
R2695 VDD2.n157 VDD2.n127 104.615
R2696 VDD2.n150 VDD2.n127 104.615
R2697 VDD2.n150 VDD2.n149 104.615
R2698 VDD2.n149 VDD2.n131 104.615
R2699 VDD2.n142 VDD2.n131 104.615
R2700 VDD2.n142 VDD2.n141 104.615
R2701 VDD2.n141 VDD2.n135 104.615
R2702 VDD2.n37 VDD2.n31 104.615
R2703 VDD2.n38 VDD2.n37 104.615
R2704 VDD2.n38 VDD2.n27 104.615
R2705 VDD2.n45 VDD2.n27 104.615
R2706 VDD2.n46 VDD2.n45 104.615
R2707 VDD2.n46 VDD2.n23 104.615
R2708 VDD2.n53 VDD2.n23 104.615
R2709 VDD2.n54 VDD2.n53 104.615
R2710 VDD2.n54 VDD2.n19 104.615
R2711 VDD2.n61 VDD2.n19 104.615
R2712 VDD2.n62 VDD2.n61 104.615
R2713 VDD2.n62 VDD2.n15 104.615
R2714 VDD2.n69 VDD2.n15 104.615
R2715 VDD2.n70 VDD2.n69 104.615
R2716 VDD2.n70 VDD2.n11 104.615
R2717 VDD2.n78 VDD2.n11 104.615
R2718 VDD2.n79 VDD2.n78 104.615
R2719 VDD2.n80 VDD2.n79 104.615
R2720 VDD2.n80 VDD2.n7 104.615
R2721 VDD2.n87 VDD2.n7 104.615
R2722 VDD2.n88 VDD2.n87 104.615
R2723 VDD2.n88 VDD2.n3 104.615
R2724 VDD2.n95 VDD2.n3 104.615
R2725 VDD2.n96 VDD2.n95 104.615
R2726 VDD2.n102 VDD2.n101 59.4227
R2727 VDD2 VDD2.n205 59.4199
R2728 VDD2.t1 VDD2.n135 52.3082
R2729 VDD2.t2 VDD2.n31 52.3082
R2730 VDD2.n102 VDD2.n100 48.4017
R2731 VDD2.n204 VDD2.n203 47.3126
R2732 VDD2.n204 VDD2.n102 44.3295
R2733 VDD2.n137 VDD2.n136 15.6677
R2734 VDD2.n33 VDD2.n32 15.6677
R2735 VDD2.n184 VDD2.n113 13.1884
R2736 VDD2.n81 VDD2.n10 13.1884
R2737 VDD2.n185 VDD2.n111 12.8005
R2738 VDD2.n180 VDD2.n115 12.8005
R2739 VDD2.n140 VDD2.n139 12.8005
R2740 VDD2.n36 VDD2.n35 12.8005
R2741 VDD2.n77 VDD2.n76 12.8005
R2742 VDD2.n82 VDD2.n8 12.8005
R2743 VDD2.n189 VDD2.n188 12.0247
R2744 VDD2.n179 VDD2.n116 12.0247
R2745 VDD2.n143 VDD2.n134 12.0247
R2746 VDD2.n39 VDD2.n30 12.0247
R2747 VDD2.n75 VDD2.n12 12.0247
R2748 VDD2.n86 VDD2.n85 12.0247
R2749 VDD2.n192 VDD2.n109 11.249
R2750 VDD2.n176 VDD2.n175 11.249
R2751 VDD2.n144 VDD2.n132 11.249
R2752 VDD2.n40 VDD2.n28 11.249
R2753 VDD2.n72 VDD2.n71 11.249
R2754 VDD2.n89 VDD2.n6 11.249
R2755 VDD2.n193 VDD2.n107 10.4732
R2756 VDD2.n172 VDD2.n118 10.4732
R2757 VDD2.n148 VDD2.n147 10.4732
R2758 VDD2.n44 VDD2.n43 10.4732
R2759 VDD2.n68 VDD2.n14 10.4732
R2760 VDD2.n90 VDD2.n4 10.4732
R2761 VDD2.n197 VDD2.n196 9.69747
R2762 VDD2.n171 VDD2.n120 9.69747
R2763 VDD2.n151 VDD2.n130 9.69747
R2764 VDD2.n47 VDD2.n26 9.69747
R2765 VDD2.n67 VDD2.n16 9.69747
R2766 VDD2.n94 VDD2.n93 9.69747
R2767 VDD2.n203 VDD2.n202 9.45567
R2768 VDD2.n100 VDD2.n99 9.45567
R2769 VDD2.n163 VDD2.n162 9.3005
R2770 VDD2.n122 VDD2.n121 9.3005
R2771 VDD2.n169 VDD2.n168 9.3005
R2772 VDD2.n171 VDD2.n170 9.3005
R2773 VDD2.n118 VDD2.n117 9.3005
R2774 VDD2.n177 VDD2.n176 9.3005
R2775 VDD2.n179 VDD2.n178 9.3005
R2776 VDD2.n115 VDD2.n112 9.3005
R2777 VDD2.n202 VDD2.n201 9.3005
R2778 VDD2.n105 VDD2.n104 9.3005
R2779 VDD2.n196 VDD2.n195 9.3005
R2780 VDD2.n194 VDD2.n193 9.3005
R2781 VDD2.n109 VDD2.n108 9.3005
R2782 VDD2.n188 VDD2.n187 9.3005
R2783 VDD2.n186 VDD2.n185 9.3005
R2784 VDD2.n161 VDD2.n160 9.3005
R2785 VDD2.n126 VDD2.n125 9.3005
R2786 VDD2.n155 VDD2.n154 9.3005
R2787 VDD2.n153 VDD2.n152 9.3005
R2788 VDD2.n130 VDD2.n129 9.3005
R2789 VDD2.n147 VDD2.n146 9.3005
R2790 VDD2.n145 VDD2.n144 9.3005
R2791 VDD2.n134 VDD2.n133 9.3005
R2792 VDD2.n139 VDD2.n138 9.3005
R2793 VDD2.n99 VDD2.n98 9.3005
R2794 VDD2.n2 VDD2.n1 9.3005
R2795 VDD2.n93 VDD2.n92 9.3005
R2796 VDD2.n91 VDD2.n90 9.3005
R2797 VDD2.n6 VDD2.n5 9.3005
R2798 VDD2.n85 VDD2.n84 9.3005
R2799 VDD2.n83 VDD2.n82 9.3005
R2800 VDD2.n22 VDD2.n21 9.3005
R2801 VDD2.n51 VDD2.n50 9.3005
R2802 VDD2.n49 VDD2.n48 9.3005
R2803 VDD2.n26 VDD2.n25 9.3005
R2804 VDD2.n43 VDD2.n42 9.3005
R2805 VDD2.n41 VDD2.n40 9.3005
R2806 VDD2.n30 VDD2.n29 9.3005
R2807 VDD2.n35 VDD2.n34 9.3005
R2808 VDD2.n57 VDD2.n56 9.3005
R2809 VDD2.n59 VDD2.n58 9.3005
R2810 VDD2.n18 VDD2.n17 9.3005
R2811 VDD2.n65 VDD2.n64 9.3005
R2812 VDD2.n67 VDD2.n66 9.3005
R2813 VDD2.n14 VDD2.n13 9.3005
R2814 VDD2.n73 VDD2.n72 9.3005
R2815 VDD2.n75 VDD2.n74 9.3005
R2816 VDD2.n76 VDD2.n9 9.3005
R2817 VDD2.n200 VDD2.n105 8.92171
R2818 VDD2.n168 VDD2.n167 8.92171
R2819 VDD2.n152 VDD2.n128 8.92171
R2820 VDD2.n48 VDD2.n24 8.92171
R2821 VDD2.n64 VDD2.n63 8.92171
R2822 VDD2.n97 VDD2.n2 8.92171
R2823 VDD2.n201 VDD2.n103 8.14595
R2824 VDD2.n164 VDD2.n122 8.14595
R2825 VDD2.n156 VDD2.n155 8.14595
R2826 VDD2.n52 VDD2.n51 8.14595
R2827 VDD2.n60 VDD2.n18 8.14595
R2828 VDD2.n98 VDD2.n0 8.14595
R2829 VDD2.n163 VDD2.n124 7.3702
R2830 VDD2.n159 VDD2.n126 7.3702
R2831 VDD2.n55 VDD2.n22 7.3702
R2832 VDD2.n59 VDD2.n20 7.3702
R2833 VDD2.n160 VDD2.n124 6.59444
R2834 VDD2.n160 VDD2.n159 6.59444
R2835 VDD2.n56 VDD2.n55 6.59444
R2836 VDD2.n56 VDD2.n20 6.59444
R2837 VDD2.n203 VDD2.n103 5.81868
R2838 VDD2.n164 VDD2.n163 5.81868
R2839 VDD2.n156 VDD2.n126 5.81868
R2840 VDD2.n52 VDD2.n22 5.81868
R2841 VDD2.n60 VDD2.n59 5.81868
R2842 VDD2.n100 VDD2.n0 5.81868
R2843 VDD2.n201 VDD2.n200 5.04292
R2844 VDD2.n167 VDD2.n122 5.04292
R2845 VDD2.n155 VDD2.n128 5.04292
R2846 VDD2.n51 VDD2.n24 5.04292
R2847 VDD2.n63 VDD2.n18 5.04292
R2848 VDD2.n98 VDD2.n97 5.04292
R2849 VDD2.n138 VDD2.n137 4.38563
R2850 VDD2.n34 VDD2.n33 4.38563
R2851 VDD2.n197 VDD2.n105 4.26717
R2852 VDD2.n168 VDD2.n120 4.26717
R2853 VDD2.n152 VDD2.n151 4.26717
R2854 VDD2.n48 VDD2.n47 4.26717
R2855 VDD2.n64 VDD2.n16 4.26717
R2856 VDD2.n94 VDD2.n2 4.26717
R2857 VDD2.n196 VDD2.n107 3.49141
R2858 VDD2.n172 VDD2.n171 3.49141
R2859 VDD2.n148 VDD2.n130 3.49141
R2860 VDD2.n44 VDD2.n26 3.49141
R2861 VDD2.n68 VDD2.n67 3.49141
R2862 VDD2.n93 VDD2.n4 3.49141
R2863 VDD2.n193 VDD2.n192 2.71565
R2864 VDD2.n175 VDD2.n118 2.71565
R2865 VDD2.n147 VDD2.n132 2.71565
R2866 VDD2.n43 VDD2.n28 2.71565
R2867 VDD2.n71 VDD2.n14 2.71565
R2868 VDD2.n90 VDD2.n89 2.71565
R2869 VDD2.n189 VDD2.n109 1.93989
R2870 VDD2.n176 VDD2.n116 1.93989
R2871 VDD2.n144 VDD2.n143 1.93989
R2872 VDD2.n40 VDD2.n39 1.93989
R2873 VDD2.n72 VDD2.n12 1.93989
R2874 VDD2.n86 VDD2.n6 1.93989
R2875 VDD2 VDD2.n204 1.20309
R2876 VDD2.n188 VDD2.n111 1.16414
R2877 VDD2.n180 VDD2.n179 1.16414
R2878 VDD2.n140 VDD2.n134 1.16414
R2879 VDD2.n36 VDD2.n30 1.16414
R2880 VDD2.n77 VDD2.n75 1.16414
R2881 VDD2.n85 VDD2.n8 1.16414
R2882 VDD2.n205 VDD2.t5 1.09081
R2883 VDD2.n205 VDD2.t3 1.09081
R2884 VDD2.n101 VDD2.t0 1.09081
R2885 VDD2.n101 VDD2.t4 1.09081
R2886 VDD2.n185 VDD2.n184 0.388379
R2887 VDD2.n115 VDD2.n113 0.388379
R2888 VDD2.n139 VDD2.n136 0.388379
R2889 VDD2.n35 VDD2.n32 0.388379
R2890 VDD2.n76 VDD2.n10 0.388379
R2891 VDD2.n82 VDD2.n81 0.388379
R2892 VDD2.n202 VDD2.n104 0.155672
R2893 VDD2.n195 VDD2.n104 0.155672
R2894 VDD2.n195 VDD2.n194 0.155672
R2895 VDD2.n194 VDD2.n108 0.155672
R2896 VDD2.n187 VDD2.n108 0.155672
R2897 VDD2.n187 VDD2.n186 0.155672
R2898 VDD2.n186 VDD2.n112 0.155672
R2899 VDD2.n178 VDD2.n112 0.155672
R2900 VDD2.n178 VDD2.n177 0.155672
R2901 VDD2.n177 VDD2.n117 0.155672
R2902 VDD2.n170 VDD2.n117 0.155672
R2903 VDD2.n170 VDD2.n169 0.155672
R2904 VDD2.n169 VDD2.n121 0.155672
R2905 VDD2.n162 VDD2.n121 0.155672
R2906 VDD2.n162 VDD2.n161 0.155672
R2907 VDD2.n161 VDD2.n125 0.155672
R2908 VDD2.n154 VDD2.n125 0.155672
R2909 VDD2.n154 VDD2.n153 0.155672
R2910 VDD2.n153 VDD2.n129 0.155672
R2911 VDD2.n146 VDD2.n129 0.155672
R2912 VDD2.n146 VDD2.n145 0.155672
R2913 VDD2.n145 VDD2.n133 0.155672
R2914 VDD2.n138 VDD2.n133 0.155672
R2915 VDD2.n34 VDD2.n29 0.155672
R2916 VDD2.n41 VDD2.n29 0.155672
R2917 VDD2.n42 VDD2.n41 0.155672
R2918 VDD2.n42 VDD2.n25 0.155672
R2919 VDD2.n49 VDD2.n25 0.155672
R2920 VDD2.n50 VDD2.n49 0.155672
R2921 VDD2.n50 VDD2.n21 0.155672
R2922 VDD2.n57 VDD2.n21 0.155672
R2923 VDD2.n58 VDD2.n57 0.155672
R2924 VDD2.n58 VDD2.n17 0.155672
R2925 VDD2.n65 VDD2.n17 0.155672
R2926 VDD2.n66 VDD2.n65 0.155672
R2927 VDD2.n66 VDD2.n13 0.155672
R2928 VDD2.n73 VDD2.n13 0.155672
R2929 VDD2.n74 VDD2.n73 0.155672
R2930 VDD2.n74 VDD2.n9 0.155672
R2931 VDD2.n83 VDD2.n9 0.155672
R2932 VDD2.n84 VDD2.n83 0.155672
R2933 VDD2.n84 VDD2.n5 0.155672
R2934 VDD2.n91 VDD2.n5 0.155672
R2935 VDD2.n92 VDD2.n91 0.155672
R2936 VDD2.n92 VDD2.n1 0.155672
R2937 VDD2.n99 VDD2.n1 0.155672
C0 VDD1 VTAIL 10.9275f
C1 VDD2 VTAIL 10.9664f
C2 VN VTAIL 8.24406f
C3 VDD1 VP 8.806769f
C4 VDD2 VP 0.361123f
C5 VP VN 6.93508f
C6 VDD1 VDD2 0.985495f
C7 VP VTAIL 8.25865f
C8 VDD1 VN 0.149455f
C9 VDD2 VN 8.600441f
C10 VDD2 B 6.171988f
C11 VDD1 B 6.232189f
C12 VTAIL B 9.355778f
C13 VN B 10.227839f
C14 VP B 8.406188f
C15 VDD2.n0 B 0.029328f
C16 VDD2.n1 B 0.021699f
C17 VDD2.n2 B 0.01166f
C18 VDD2.n3 B 0.02756f
C19 VDD2.n4 B 0.012346f
C20 VDD2.n5 B 0.021699f
C21 VDD2.n6 B 0.01166f
C22 VDD2.n7 B 0.02756f
C23 VDD2.n8 B 0.012346f
C24 VDD2.n9 B 0.021699f
C25 VDD2.n10 B 0.012003f
C26 VDD2.n11 B 0.02756f
C27 VDD2.n12 B 0.012346f
C28 VDD2.n13 B 0.021699f
C29 VDD2.n14 B 0.01166f
C30 VDD2.n15 B 0.02756f
C31 VDD2.n16 B 0.012346f
C32 VDD2.n17 B 0.021699f
C33 VDD2.n18 B 0.01166f
C34 VDD2.n19 B 0.02756f
C35 VDD2.n20 B 0.012346f
C36 VDD2.n21 B 0.021699f
C37 VDD2.n22 B 0.01166f
C38 VDD2.n23 B 0.02756f
C39 VDD2.n24 B 0.012346f
C40 VDD2.n25 B 0.021699f
C41 VDD2.n26 B 0.01166f
C42 VDD2.n27 B 0.02756f
C43 VDD2.n28 B 0.012346f
C44 VDD2.n29 B 0.021699f
C45 VDD2.n30 B 0.01166f
C46 VDD2.n31 B 0.02067f
C47 VDD2.n32 B 0.016281f
C48 VDD2.t2 B 0.045678f
C49 VDD2.n33 B 0.158716f
C50 VDD2.n34 B 1.72601f
C51 VDD2.n35 B 0.01166f
C52 VDD2.n36 B 0.012346f
C53 VDD2.n37 B 0.02756f
C54 VDD2.n38 B 0.02756f
C55 VDD2.n39 B 0.012346f
C56 VDD2.n40 B 0.01166f
C57 VDD2.n41 B 0.021699f
C58 VDD2.n42 B 0.021699f
C59 VDD2.n43 B 0.01166f
C60 VDD2.n44 B 0.012346f
C61 VDD2.n45 B 0.02756f
C62 VDD2.n46 B 0.02756f
C63 VDD2.n47 B 0.012346f
C64 VDD2.n48 B 0.01166f
C65 VDD2.n49 B 0.021699f
C66 VDD2.n50 B 0.021699f
C67 VDD2.n51 B 0.01166f
C68 VDD2.n52 B 0.012346f
C69 VDD2.n53 B 0.02756f
C70 VDD2.n54 B 0.02756f
C71 VDD2.n55 B 0.012346f
C72 VDD2.n56 B 0.01166f
C73 VDD2.n57 B 0.021699f
C74 VDD2.n58 B 0.021699f
C75 VDD2.n59 B 0.01166f
C76 VDD2.n60 B 0.012346f
C77 VDD2.n61 B 0.02756f
C78 VDD2.n62 B 0.02756f
C79 VDD2.n63 B 0.012346f
C80 VDD2.n64 B 0.01166f
C81 VDD2.n65 B 0.021699f
C82 VDD2.n66 B 0.021699f
C83 VDD2.n67 B 0.01166f
C84 VDD2.n68 B 0.012346f
C85 VDD2.n69 B 0.02756f
C86 VDD2.n70 B 0.02756f
C87 VDD2.n71 B 0.012346f
C88 VDD2.n72 B 0.01166f
C89 VDD2.n73 B 0.021699f
C90 VDD2.n74 B 0.021699f
C91 VDD2.n75 B 0.01166f
C92 VDD2.n76 B 0.01166f
C93 VDD2.n77 B 0.012346f
C94 VDD2.n78 B 0.02756f
C95 VDD2.n79 B 0.02756f
C96 VDD2.n80 B 0.02756f
C97 VDD2.n81 B 0.012003f
C98 VDD2.n82 B 0.01166f
C99 VDD2.n83 B 0.021699f
C100 VDD2.n84 B 0.021699f
C101 VDD2.n85 B 0.01166f
C102 VDD2.n86 B 0.012346f
C103 VDD2.n87 B 0.02756f
C104 VDD2.n88 B 0.02756f
C105 VDD2.n89 B 0.012346f
C106 VDD2.n90 B 0.01166f
C107 VDD2.n91 B 0.021699f
C108 VDD2.n92 B 0.021699f
C109 VDD2.n93 B 0.01166f
C110 VDD2.n94 B 0.012346f
C111 VDD2.n95 B 0.02756f
C112 VDD2.n96 B 0.057592f
C113 VDD2.n97 B 0.012346f
C114 VDD2.n98 B 0.01166f
C115 VDD2.n99 B 0.047784f
C116 VDD2.n100 B 0.049573f
C117 VDD2.t0 B 0.311391f
C118 VDD2.t4 B 0.311391f
C119 VDD2.n101 B 2.83738f
C120 VDD2.n102 B 2.22237f
C121 VDD2.n103 B 0.029328f
C122 VDD2.n104 B 0.021699f
C123 VDD2.n105 B 0.01166f
C124 VDD2.n106 B 0.02756f
C125 VDD2.n107 B 0.012346f
C126 VDD2.n108 B 0.021699f
C127 VDD2.n109 B 0.01166f
C128 VDD2.n110 B 0.02756f
C129 VDD2.n111 B 0.012346f
C130 VDD2.n112 B 0.021699f
C131 VDD2.n113 B 0.012003f
C132 VDD2.n114 B 0.02756f
C133 VDD2.n115 B 0.01166f
C134 VDD2.n116 B 0.012346f
C135 VDD2.n117 B 0.021699f
C136 VDD2.n118 B 0.01166f
C137 VDD2.n119 B 0.02756f
C138 VDD2.n120 B 0.012346f
C139 VDD2.n121 B 0.021699f
C140 VDD2.n122 B 0.01166f
C141 VDD2.n123 B 0.02756f
C142 VDD2.n124 B 0.012346f
C143 VDD2.n125 B 0.021699f
C144 VDD2.n126 B 0.01166f
C145 VDD2.n127 B 0.02756f
C146 VDD2.n128 B 0.012346f
C147 VDD2.n129 B 0.021699f
C148 VDD2.n130 B 0.01166f
C149 VDD2.n131 B 0.02756f
C150 VDD2.n132 B 0.012346f
C151 VDD2.n133 B 0.021699f
C152 VDD2.n134 B 0.01166f
C153 VDD2.n135 B 0.02067f
C154 VDD2.n136 B 0.016281f
C155 VDD2.t1 B 0.045678f
C156 VDD2.n137 B 0.158716f
C157 VDD2.n138 B 1.72601f
C158 VDD2.n139 B 0.01166f
C159 VDD2.n140 B 0.012346f
C160 VDD2.n141 B 0.02756f
C161 VDD2.n142 B 0.02756f
C162 VDD2.n143 B 0.012346f
C163 VDD2.n144 B 0.01166f
C164 VDD2.n145 B 0.021699f
C165 VDD2.n146 B 0.021699f
C166 VDD2.n147 B 0.01166f
C167 VDD2.n148 B 0.012346f
C168 VDD2.n149 B 0.02756f
C169 VDD2.n150 B 0.02756f
C170 VDD2.n151 B 0.012346f
C171 VDD2.n152 B 0.01166f
C172 VDD2.n153 B 0.021699f
C173 VDD2.n154 B 0.021699f
C174 VDD2.n155 B 0.01166f
C175 VDD2.n156 B 0.012346f
C176 VDD2.n157 B 0.02756f
C177 VDD2.n158 B 0.02756f
C178 VDD2.n159 B 0.012346f
C179 VDD2.n160 B 0.01166f
C180 VDD2.n161 B 0.021699f
C181 VDD2.n162 B 0.021699f
C182 VDD2.n163 B 0.01166f
C183 VDD2.n164 B 0.012346f
C184 VDD2.n165 B 0.02756f
C185 VDD2.n166 B 0.02756f
C186 VDD2.n167 B 0.012346f
C187 VDD2.n168 B 0.01166f
C188 VDD2.n169 B 0.021699f
C189 VDD2.n170 B 0.021699f
C190 VDD2.n171 B 0.01166f
C191 VDD2.n172 B 0.012346f
C192 VDD2.n173 B 0.02756f
C193 VDD2.n174 B 0.02756f
C194 VDD2.n175 B 0.012346f
C195 VDD2.n176 B 0.01166f
C196 VDD2.n177 B 0.021699f
C197 VDD2.n178 B 0.021699f
C198 VDD2.n179 B 0.01166f
C199 VDD2.n180 B 0.012346f
C200 VDD2.n181 B 0.02756f
C201 VDD2.n182 B 0.02756f
C202 VDD2.n183 B 0.02756f
C203 VDD2.n184 B 0.012003f
C204 VDD2.n185 B 0.01166f
C205 VDD2.n186 B 0.021699f
C206 VDD2.n187 B 0.021699f
C207 VDD2.n188 B 0.01166f
C208 VDD2.n189 B 0.012346f
C209 VDD2.n190 B 0.02756f
C210 VDD2.n191 B 0.02756f
C211 VDD2.n192 B 0.012346f
C212 VDD2.n193 B 0.01166f
C213 VDD2.n194 B 0.021699f
C214 VDD2.n195 B 0.021699f
C215 VDD2.n196 B 0.01166f
C216 VDD2.n197 B 0.012346f
C217 VDD2.n198 B 0.02756f
C218 VDD2.n199 B 0.057592f
C219 VDD2.n200 B 0.012346f
C220 VDD2.n201 B 0.01166f
C221 VDD2.n202 B 0.047784f
C222 VDD2.n203 B 0.04694f
C223 VDD2.n204 B 2.35778f
C224 VDD2.t5 B 0.311391f
C225 VDD2.t3 B 0.311391f
C226 VDD2.n205 B 2.83736f
C227 VN.n0 B 0.032232f
C228 VN.t1 B 2.31877f
C229 VN.n1 B 0.057914f
C230 VN.t3 B 2.41853f
C231 VN.t5 B 2.31877f
C232 VN.n2 B 0.890846f
C233 VN.n3 B 0.884335f
C234 VN.n4 B 0.204092f
C235 VN.n5 B 0.032232f
C236 VN.n6 B 0.03191f
C237 VN.n7 B 0.050082f
C238 VN.n8 B 0.884319f
C239 VN.n9 B 0.029708f
C240 VN.n10 B 0.032232f
C241 VN.t4 B 2.31877f
C242 VN.n11 B 0.057914f
C243 VN.t2 B 2.41853f
C244 VN.t0 B 2.31877f
C245 VN.n12 B 0.890846f
C246 VN.n13 B 0.884335f
C247 VN.n14 B 0.204092f
C248 VN.n15 B 0.032232f
C249 VN.n16 B 0.03191f
C250 VN.n17 B 0.050082f
C251 VN.n18 B 0.884319f
C252 VN.n19 B 1.71237f
C253 VTAIL.t2 B 0.321496f
C254 VTAIL.t0 B 0.321496f
C255 VTAIL.n0 B 2.85521f
C256 VTAIL.n1 B 0.351151f
C257 VTAIL.n2 B 0.03028f
C258 VTAIL.n3 B 0.022403f
C259 VTAIL.n4 B 0.012038f
C260 VTAIL.n5 B 0.028454f
C261 VTAIL.n6 B 0.012746f
C262 VTAIL.n7 B 0.022403f
C263 VTAIL.n8 B 0.012038f
C264 VTAIL.n9 B 0.028454f
C265 VTAIL.n10 B 0.012746f
C266 VTAIL.n11 B 0.022403f
C267 VTAIL.n12 B 0.012392f
C268 VTAIL.n13 B 0.028454f
C269 VTAIL.n14 B 0.012746f
C270 VTAIL.n15 B 0.022403f
C271 VTAIL.n16 B 0.012038f
C272 VTAIL.n17 B 0.028454f
C273 VTAIL.n18 B 0.012746f
C274 VTAIL.n19 B 0.022403f
C275 VTAIL.n20 B 0.012038f
C276 VTAIL.n21 B 0.028454f
C277 VTAIL.n22 B 0.012746f
C278 VTAIL.n23 B 0.022403f
C279 VTAIL.n24 B 0.012038f
C280 VTAIL.n25 B 0.028454f
C281 VTAIL.n26 B 0.012746f
C282 VTAIL.n27 B 0.022403f
C283 VTAIL.n28 B 0.012038f
C284 VTAIL.n29 B 0.028454f
C285 VTAIL.n30 B 0.012746f
C286 VTAIL.n31 B 0.022403f
C287 VTAIL.n32 B 0.012038f
C288 VTAIL.n33 B 0.021341f
C289 VTAIL.n34 B 0.016809f
C290 VTAIL.t5 B 0.047161f
C291 VTAIL.n35 B 0.163867f
C292 VTAIL.n36 B 1.78202f
C293 VTAIL.n37 B 0.012038f
C294 VTAIL.n38 B 0.012746f
C295 VTAIL.n39 B 0.028454f
C296 VTAIL.n40 B 0.028454f
C297 VTAIL.n41 B 0.012746f
C298 VTAIL.n42 B 0.012038f
C299 VTAIL.n43 B 0.022403f
C300 VTAIL.n44 B 0.022403f
C301 VTAIL.n45 B 0.012038f
C302 VTAIL.n46 B 0.012746f
C303 VTAIL.n47 B 0.028454f
C304 VTAIL.n48 B 0.028454f
C305 VTAIL.n49 B 0.012746f
C306 VTAIL.n50 B 0.012038f
C307 VTAIL.n51 B 0.022403f
C308 VTAIL.n52 B 0.022403f
C309 VTAIL.n53 B 0.012038f
C310 VTAIL.n54 B 0.012746f
C311 VTAIL.n55 B 0.028454f
C312 VTAIL.n56 B 0.028454f
C313 VTAIL.n57 B 0.012746f
C314 VTAIL.n58 B 0.012038f
C315 VTAIL.n59 B 0.022403f
C316 VTAIL.n60 B 0.022403f
C317 VTAIL.n61 B 0.012038f
C318 VTAIL.n62 B 0.012746f
C319 VTAIL.n63 B 0.028454f
C320 VTAIL.n64 B 0.028454f
C321 VTAIL.n65 B 0.012746f
C322 VTAIL.n66 B 0.012038f
C323 VTAIL.n67 B 0.022403f
C324 VTAIL.n68 B 0.022403f
C325 VTAIL.n69 B 0.012038f
C326 VTAIL.n70 B 0.012746f
C327 VTAIL.n71 B 0.028454f
C328 VTAIL.n72 B 0.028454f
C329 VTAIL.n73 B 0.012746f
C330 VTAIL.n74 B 0.012038f
C331 VTAIL.n75 B 0.022403f
C332 VTAIL.n76 B 0.022403f
C333 VTAIL.n77 B 0.012038f
C334 VTAIL.n78 B 0.012038f
C335 VTAIL.n79 B 0.012746f
C336 VTAIL.n80 B 0.028454f
C337 VTAIL.n81 B 0.028454f
C338 VTAIL.n82 B 0.028454f
C339 VTAIL.n83 B 0.012392f
C340 VTAIL.n84 B 0.012038f
C341 VTAIL.n85 B 0.022403f
C342 VTAIL.n86 B 0.022403f
C343 VTAIL.n87 B 0.012038f
C344 VTAIL.n88 B 0.012746f
C345 VTAIL.n89 B 0.028454f
C346 VTAIL.n90 B 0.028454f
C347 VTAIL.n91 B 0.012746f
C348 VTAIL.n92 B 0.012038f
C349 VTAIL.n93 B 0.022403f
C350 VTAIL.n94 B 0.022403f
C351 VTAIL.n95 B 0.012038f
C352 VTAIL.n96 B 0.012746f
C353 VTAIL.n97 B 0.028454f
C354 VTAIL.n98 B 0.059461f
C355 VTAIL.n99 B 0.012746f
C356 VTAIL.n100 B 0.012038f
C357 VTAIL.n101 B 0.049335f
C358 VTAIL.n102 B 0.032974f
C359 VTAIL.n103 B 0.216891f
C360 VTAIL.t8 B 0.321496f
C361 VTAIL.t9 B 0.321496f
C362 VTAIL.n104 B 2.85521f
C363 VTAIL.n105 B 1.99529f
C364 VTAIL.t1 B 0.321496f
C365 VTAIL.t4 B 0.321496f
C366 VTAIL.n106 B 2.85522f
C367 VTAIL.n107 B 1.99528f
C368 VTAIL.n108 B 0.03028f
C369 VTAIL.n109 B 0.022403f
C370 VTAIL.n110 B 0.012038f
C371 VTAIL.n111 B 0.028454f
C372 VTAIL.n112 B 0.012746f
C373 VTAIL.n113 B 0.022403f
C374 VTAIL.n114 B 0.012038f
C375 VTAIL.n115 B 0.028454f
C376 VTAIL.n116 B 0.012746f
C377 VTAIL.n117 B 0.022403f
C378 VTAIL.n118 B 0.012392f
C379 VTAIL.n119 B 0.028454f
C380 VTAIL.n120 B 0.012038f
C381 VTAIL.n121 B 0.012746f
C382 VTAIL.n122 B 0.022403f
C383 VTAIL.n123 B 0.012038f
C384 VTAIL.n124 B 0.028454f
C385 VTAIL.n125 B 0.012746f
C386 VTAIL.n126 B 0.022403f
C387 VTAIL.n127 B 0.012038f
C388 VTAIL.n128 B 0.028454f
C389 VTAIL.n129 B 0.012746f
C390 VTAIL.n130 B 0.022403f
C391 VTAIL.n131 B 0.012038f
C392 VTAIL.n132 B 0.028454f
C393 VTAIL.n133 B 0.012746f
C394 VTAIL.n134 B 0.022403f
C395 VTAIL.n135 B 0.012038f
C396 VTAIL.n136 B 0.028454f
C397 VTAIL.n137 B 0.012746f
C398 VTAIL.n138 B 0.022403f
C399 VTAIL.n139 B 0.012038f
C400 VTAIL.n140 B 0.021341f
C401 VTAIL.n141 B 0.016809f
C402 VTAIL.t3 B 0.047161f
C403 VTAIL.n142 B 0.163867f
C404 VTAIL.n143 B 1.78202f
C405 VTAIL.n144 B 0.012038f
C406 VTAIL.n145 B 0.012746f
C407 VTAIL.n146 B 0.028454f
C408 VTAIL.n147 B 0.028454f
C409 VTAIL.n148 B 0.012746f
C410 VTAIL.n149 B 0.012038f
C411 VTAIL.n150 B 0.022403f
C412 VTAIL.n151 B 0.022403f
C413 VTAIL.n152 B 0.012038f
C414 VTAIL.n153 B 0.012746f
C415 VTAIL.n154 B 0.028454f
C416 VTAIL.n155 B 0.028454f
C417 VTAIL.n156 B 0.012746f
C418 VTAIL.n157 B 0.012038f
C419 VTAIL.n158 B 0.022403f
C420 VTAIL.n159 B 0.022403f
C421 VTAIL.n160 B 0.012038f
C422 VTAIL.n161 B 0.012746f
C423 VTAIL.n162 B 0.028454f
C424 VTAIL.n163 B 0.028454f
C425 VTAIL.n164 B 0.012746f
C426 VTAIL.n165 B 0.012038f
C427 VTAIL.n166 B 0.022403f
C428 VTAIL.n167 B 0.022403f
C429 VTAIL.n168 B 0.012038f
C430 VTAIL.n169 B 0.012746f
C431 VTAIL.n170 B 0.028454f
C432 VTAIL.n171 B 0.028454f
C433 VTAIL.n172 B 0.012746f
C434 VTAIL.n173 B 0.012038f
C435 VTAIL.n174 B 0.022403f
C436 VTAIL.n175 B 0.022403f
C437 VTAIL.n176 B 0.012038f
C438 VTAIL.n177 B 0.012746f
C439 VTAIL.n178 B 0.028454f
C440 VTAIL.n179 B 0.028454f
C441 VTAIL.n180 B 0.012746f
C442 VTAIL.n181 B 0.012038f
C443 VTAIL.n182 B 0.022403f
C444 VTAIL.n183 B 0.022403f
C445 VTAIL.n184 B 0.012038f
C446 VTAIL.n185 B 0.012746f
C447 VTAIL.n186 B 0.028454f
C448 VTAIL.n187 B 0.028454f
C449 VTAIL.n188 B 0.028454f
C450 VTAIL.n189 B 0.012392f
C451 VTAIL.n190 B 0.012038f
C452 VTAIL.n191 B 0.022403f
C453 VTAIL.n192 B 0.022403f
C454 VTAIL.n193 B 0.012038f
C455 VTAIL.n194 B 0.012746f
C456 VTAIL.n195 B 0.028454f
C457 VTAIL.n196 B 0.028454f
C458 VTAIL.n197 B 0.012746f
C459 VTAIL.n198 B 0.012038f
C460 VTAIL.n199 B 0.022403f
C461 VTAIL.n200 B 0.022403f
C462 VTAIL.n201 B 0.012038f
C463 VTAIL.n202 B 0.012746f
C464 VTAIL.n203 B 0.028454f
C465 VTAIL.n204 B 0.059461f
C466 VTAIL.n205 B 0.012746f
C467 VTAIL.n206 B 0.012038f
C468 VTAIL.n207 B 0.049335f
C469 VTAIL.n208 B 0.032974f
C470 VTAIL.n209 B 0.216891f
C471 VTAIL.t7 B 0.321496f
C472 VTAIL.t10 B 0.321496f
C473 VTAIL.n210 B 2.85522f
C474 VTAIL.n211 B 0.429548f
C475 VTAIL.n212 B 0.03028f
C476 VTAIL.n213 B 0.022403f
C477 VTAIL.n214 B 0.012038f
C478 VTAIL.n215 B 0.028454f
C479 VTAIL.n216 B 0.012746f
C480 VTAIL.n217 B 0.022403f
C481 VTAIL.n218 B 0.012038f
C482 VTAIL.n219 B 0.028454f
C483 VTAIL.n220 B 0.012746f
C484 VTAIL.n221 B 0.022403f
C485 VTAIL.n222 B 0.012392f
C486 VTAIL.n223 B 0.028454f
C487 VTAIL.n224 B 0.012038f
C488 VTAIL.n225 B 0.012746f
C489 VTAIL.n226 B 0.022403f
C490 VTAIL.n227 B 0.012038f
C491 VTAIL.n228 B 0.028454f
C492 VTAIL.n229 B 0.012746f
C493 VTAIL.n230 B 0.022403f
C494 VTAIL.n231 B 0.012038f
C495 VTAIL.n232 B 0.028454f
C496 VTAIL.n233 B 0.012746f
C497 VTAIL.n234 B 0.022403f
C498 VTAIL.n235 B 0.012038f
C499 VTAIL.n236 B 0.028454f
C500 VTAIL.n237 B 0.012746f
C501 VTAIL.n238 B 0.022403f
C502 VTAIL.n239 B 0.012038f
C503 VTAIL.n240 B 0.028454f
C504 VTAIL.n241 B 0.012746f
C505 VTAIL.n242 B 0.022403f
C506 VTAIL.n243 B 0.012038f
C507 VTAIL.n244 B 0.021341f
C508 VTAIL.n245 B 0.016809f
C509 VTAIL.t6 B 0.047161f
C510 VTAIL.n246 B 0.163867f
C511 VTAIL.n247 B 1.78202f
C512 VTAIL.n248 B 0.012038f
C513 VTAIL.n249 B 0.012746f
C514 VTAIL.n250 B 0.028454f
C515 VTAIL.n251 B 0.028454f
C516 VTAIL.n252 B 0.012746f
C517 VTAIL.n253 B 0.012038f
C518 VTAIL.n254 B 0.022403f
C519 VTAIL.n255 B 0.022403f
C520 VTAIL.n256 B 0.012038f
C521 VTAIL.n257 B 0.012746f
C522 VTAIL.n258 B 0.028454f
C523 VTAIL.n259 B 0.028454f
C524 VTAIL.n260 B 0.012746f
C525 VTAIL.n261 B 0.012038f
C526 VTAIL.n262 B 0.022403f
C527 VTAIL.n263 B 0.022403f
C528 VTAIL.n264 B 0.012038f
C529 VTAIL.n265 B 0.012746f
C530 VTAIL.n266 B 0.028454f
C531 VTAIL.n267 B 0.028454f
C532 VTAIL.n268 B 0.012746f
C533 VTAIL.n269 B 0.012038f
C534 VTAIL.n270 B 0.022403f
C535 VTAIL.n271 B 0.022403f
C536 VTAIL.n272 B 0.012038f
C537 VTAIL.n273 B 0.012746f
C538 VTAIL.n274 B 0.028454f
C539 VTAIL.n275 B 0.028454f
C540 VTAIL.n276 B 0.012746f
C541 VTAIL.n277 B 0.012038f
C542 VTAIL.n278 B 0.022403f
C543 VTAIL.n279 B 0.022403f
C544 VTAIL.n280 B 0.012038f
C545 VTAIL.n281 B 0.012746f
C546 VTAIL.n282 B 0.028454f
C547 VTAIL.n283 B 0.028454f
C548 VTAIL.n284 B 0.012746f
C549 VTAIL.n285 B 0.012038f
C550 VTAIL.n286 B 0.022403f
C551 VTAIL.n287 B 0.022403f
C552 VTAIL.n288 B 0.012038f
C553 VTAIL.n289 B 0.012746f
C554 VTAIL.n290 B 0.028454f
C555 VTAIL.n291 B 0.028454f
C556 VTAIL.n292 B 0.028454f
C557 VTAIL.n293 B 0.012392f
C558 VTAIL.n294 B 0.012038f
C559 VTAIL.n295 B 0.022403f
C560 VTAIL.n296 B 0.022403f
C561 VTAIL.n297 B 0.012038f
C562 VTAIL.n298 B 0.012746f
C563 VTAIL.n299 B 0.028454f
C564 VTAIL.n300 B 0.028454f
C565 VTAIL.n301 B 0.012746f
C566 VTAIL.n302 B 0.012038f
C567 VTAIL.n303 B 0.022403f
C568 VTAIL.n304 B 0.022403f
C569 VTAIL.n305 B 0.012038f
C570 VTAIL.n306 B 0.012746f
C571 VTAIL.n307 B 0.028454f
C572 VTAIL.n308 B 0.059461f
C573 VTAIL.n309 B 0.012746f
C574 VTAIL.n310 B 0.012038f
C575 VTAIL.n311 B 0.049335f
C576 VTAIL.n312 B 0.032974f
C577 VTAIL.n313 B 1.67247f
C578 VTAIL.n314 B 0.03028f
C579 VTAIL.n315 B 0.022403f
C580 VTAIL.n316 B 0.012038f
C581 VTAIL.n317 B 0.028454f
C582 VTAIL.n318 B 0.012746f
C583 VTAIL.n319 B 0.022403f
C584 VTAIL.n320 B 0.012038f
C585 VTAIL.n321 B 0.028454f
C586 VTAIL.n322 B 0.012746f
C587 VTAIL.n323 B 0.022403f
C588 VTAIL.n324 B 0.012392f
C589 VTAIL.n325 B 0.028454f
C590 VTAIL.n326 B 0.012746f
C591 VTAIL.n327 B 0.022403f
C592 VTAIL.n328 B 0.012038f
C593 VTAIL.n329 B 0.028454f
C594 VTAIL.n330 B 0.012746f
C595 VTAIL.n331 B 0.022403f
C596 VTAIL.n332 B 0.012038f
C597 VTAIL.n333 B 0.028454f
C598 VTAIL.n334 B 0.012746f
C599 VTAIL.n335 B 0.022403f
C600 VTAIL.n336 B 0.012038f
C601 VTAIL.n337 B 0.028454f
C602 VTAIL.n338 B 0.012746f
C603 VTAIL.n339 B 0.022403f
C604 VTAIL.n340 B 0.012038f
C605 VTAIL.n341 B 0.028454f
C606 VTAIL.n342 B 0.012746f
C607 VTAIL.n343 B 0.022403f
C608 VTAIL.n344 B 0.012038f
C609 VTAIL.n345 B 0.021341f
C610 VTAIL.n346 B 0.016809f
C611 VTAIL.t11 B 0.047161f
C612 VTAIL.n347 B 0.163867f
C613 VTAIL.n348 B 1.78202f
C614 VTAIL.n349 B 0.012038f
C615 VTAIL.n350 B 0.012746f
C616 VTAIL.n351 B 0.028454f
C617 VTAIL.n352 B 0.028454f
C618 VTAIL.n353 B 0.012746f
C619 VTAIL.n354 B 0.012038f
C620 VTAIL.n355 B 0.022403f
C621 VTAIL.n356 B 0.022403f
C622 VTAIL.n357 B 0.012038f
C623 VTAIL.n358 B 0.012746f
C624 VTAIL.n359 B 0.028454f
C625 VTAIL.n360 B 0.028454f
C626 VTAIL.n361 B 0.012746f
C627 VTAIL.n362 B 0.012038f
C628 VTAIL.n363 B 0.022403f
C629 VTAIL.n364 B 0.022403f
C630 VTAIL.n365 B 0.012038f
C631 VTAIL.n366 B 0.012746f
C632 VTAIL.n367 B 0.028454f
C633 VTAIL.n368 B 0.028454f
C634 VTAIL.n369 B 0.012746f
C635 VTAIL.n370 B 0.012038f
C636 VTAIL.n371 B 0.022403f
C637 VTAIL.n372 B 0.022403f
C638 VTAIL.n373 B 0.012038f
C639 VTAIL.n374 B 0.012746f
C640 VTAIL.n375 B 0.028454f
C641 VTAIL.n376 B 0.028454f
C642 VTAIL.n377 B 0.012746f
C643 VTAIL.n378 B 0.012038f
C644 VTAIL.n379 B 0.022403f
C645 VTAIL.n380 B 0.022403f
C646 VTAIL.n381 B 0.012038f
C647 VTAIL.n382 B 0.012746f
C648 VTAIL.n383 B 0.028454f
C649 VTAIL.n384 B 0.028454f
C650 VTAIL.n385 B 0.012746f
C651 VTAIL.n386 B 0.012038f
C652 VTAIL.n387 B 0.022403f
C653 VTAIL.n388 B 0.022403f
C654 VTAIL.n389 B 0.012038f
C655 VTAIL.n390 B 0.012038f
C656 VTAIL.n391 B 0.012746f
C657 VTAIL.n392 B 0.028454f
C658 VTAIL.n393 B 0.028454f
C659 VTAIL.n394 B 0.028454f
C660 VTAIL.n395 B 0.012392f
C661 VTAIL.n396 B 0.012038f
C662 VTAIL.n397 B 0.022403f
C663 VTAIL.n398 B 0.022403f
C664 VTAIL.n399 B 0.012038f
C665 VTAIL.n400 B 0.012746f
C666 VTAIL.n401 B 0.028454f
C667 VTAIL.n402 B 0.028454f
C668 VTAIL.n403 B 0.012746f
C669 VTAIL.n404 B 0.012038f
C670 VTAIL.n405 B 0.022403f
C671 VTAIL.n406 B 0.022403f
C672 VTAIL.n407 B 0.012038f
C673 VTAIL.n408 B 0.012746f
C674 VTAIL.n409 B 0.028454f
C675 VTAIL.n410 B 0.059461f
C676 VTAIL.n411 B 0.012746f
C677 VTAIL.n412 B 0.012038f
C678 VTAIL.n413 B 0.049335f
C679 VTAIL.n414 B 0.032974f
C680 VTAIL.n415 B 1.64074f
C681 VDD1.n0 B 0.029358f
C682 VDD1.n1 B 0.021721f
C683 VDD1.n2 B 0.011672f
C684 VDD1.n3 B 0.027588f
C685 VDD1.n4 B 0.012358f
C686 VDD1.n5 B 0.021721f
C687 VDD1.n6 B 0.011672f
C688 VDD1.n7 B 0.027588f
C689 VDD1.n8 B 0.012358f
C690 VDD1.n9 B 0.021721f
C691 VDD1.n10 B 0.012015f
C692 VDD1.n11 B 0.027588f
C693 VDD1.n12 B 0.011672f
C694 VDD1.n13 B 0.012358f
C695 VDD1.n14 B 0.021721f
C696 VDD1.n15 B 0.011672f
C697 VDD1.n16 B 0.027588f
C698 VDD1.n17 B 0.012358f
C699 VDD1.n18 B 0.021721f
C700 VDD1.n19 B 0.011672f
C701 VDD1.n20 B 0.027588f
C702 VDD1.n21 B 0.012358f
C703 VDD1.n22 B 0.021721f
C704 VDD1.n23 B 0.011672f
C705 VDD1.n24 B 0.027588f
C706 VDD1.n25 B 0.012358f
C707 VDD1.n26 B 0.021721f
C708 VDD1.n27 B 0.011672f
C709 VDD1.n28 B 0.027588f
C710 VDD1.n29 B 0.012358f
C711 VDD1.n30 B 0.021721f
C712 VDD1.n31 B 0.011672f
C713 VDD1.n32 B 0.020691f
C714 VDD1.n33 B 0.016297f
C715 VDD1.t1 B 0.045724f
C716 VDD1.n34 B 0.158876f
C717 VDD1.n35 B 1.72775f
C718 VDD1.n36 B 0.011672f
C719 VDD1.n37 B 0.012358f
C720 VDD1.n38 B 0.027588f
C721 VDD1.n39 B 0.027588f
C722 VDD1.n40 B 0.012358f
C723 VDD1.n41 B 0.011672f
C724 VDD1.n42 B 0.021721f
C725 VDD1.n43 B 0.021721f
C726 VDD1.n44 B 0.011672f
C727 VDD1.n45 B 0.012358f
C728 VDD1.n46 B 0.027588f
C729 VDD1.n47 B 0.027588f
C730 VDD1.n48 B 0.012358f
C731 VDD1.n49 B 0.011672f
C732 VDD1.n50 B 0.021721f
C733 VDD1.n51 B 0.021721f
C734 VDD1.n52 B 0.011672f
C735 VDD1.n53 B 0.012358f
C736 VDD1.n54 B 0.027588f
C737 VDD1.n55 B 0.027588f
C738 VDD1.n56 B 0.012358f
C739 VDD1.n57 B 0.011672f
C740 VDD1.n58 B 0.021721f
C741 VDD1.n59 B 0.021721f
C742 VDD1.n60 B 0.011672f
C743 VDD1.n61 B 0.012358f
C744 VDD1.n62 B 0.027588f
C745 VDD1.n63 B 0.027588f
C746 VDD1.n64 B 0.012358f
C747 VDD1.n65 B 0.011672f
C748 VDD1.n66 B 0.021721f
C749 VDD1.n67 B 0.021721f
C750 VDD1.n68 B 0.011672f
C751 VDD1.n69 B 0.012358f
C752 VDD1.n70 B 0.027588f
C753 VDD1.n71 B 0.027588f
C754 VDD1.n72 B 0.012358f
C755 VDD1.n73 B 0.011672f
C756 VDD1.n74 B 0.021721f
C757 VDD1.n75 B 0.021721f
C758 VDD1.n76 B 0.011672f
C759 VDD1.n77 B 0.012358f
C760 VDD1.n78 B 0.027588f
C761 VDD1.n79 B 0.027588f
C762 VDD1.n80 B 0.027588f
C763 VDD1.n81 B 0.012015f
C764 VDD1.n82 B 0.011672f
C765 VDD1.n83 B 0.021721f
C766 VDD1.n84 B 0.021721f
C767 VDD1.n85 B 0.011672f
C768 VDD1.n86 B 0.012358f
C769 VDD1.n87 B 0.027588f
C770 VDD1.n88 B 0.027588f
C771 VDD1.n89 B 0.012358f
C772 VDD1.n90 B 0.011672f
C773 VDD1.n91 B 0.021721f
C774 VDD1.n92 B 0.021721f
C775 VDD1.n93 B 0.011672f
C776 VDD1.n94 B 0.012358f
C777 VDD1.n95 B 0.027588f
C778 VDD1.n96 B 0.05765f
C779 VDD1.n97 B 0.012358f
C780 VDD1.n98 B 0.011672f
C781 VDD1.n99 B 0.047833f
C782 VDD1.n100 B 0.050077f
C783 VDD1.n101 B 0.029358f
C784 VDD1.n102 B 0.021721f
C785 VDD1.n103 B 0.011672f
C786 VDD1.n104 B 0.027588f
C787 VDD1.n105 B 0.012358f
C788 VDD1.n106 B 0.021721f
C789 VDD1.n107 B 0.011672f
C790 VDD1.n108 B 0.027588f
C791 VDD1.n109 B 0.012358f
C792 VDD1.n110 B 0.021721f
C793 VDD1.n111 B 0.012015f
C794 VDD1.n112 B 0.027588f
C795 VDD1.n113 B 0.012358f
C796 VDD1.n114 B 0.021721f
C797 VDD1.n115 B 0.011672f
C798 VDD1.n116 B 0.027588f
C799 VDD1.n117 B 0.012358f
C800 VDD1.n118 B 0.021721f
C801 VDD1.n119 B 0.011672f
C802 VDD1.n120 B 0.027588f
C803 VDD1.n121 B 0.012358f
C804 VDD1.n122 B 0.021721f
C805 VDD1.n123 B 0.011672f
C806 VDD1.n124 B 0.027588f
C807 VDD1.n125 B 0.012358f
C808 VDD1.n126 B 0.021721f
C809 VDD1.n127 B 0.011672f
C810 VDD1.n128 B 0.027588f
C811 VDD1.n129 B 0.012358f
C812 VDD1.n130 B 0.021721f
C813 VDD1.n131 B 0.011672f
C814 VDD1.n132 B 0.020691f
C815 VDD1.n133 B 0.016297f
C816 VDD1.t4 B 0.045724f
C817 VDD1.n134 B 0.158876f
C818 VDD1.n135 B 1.72775f
C819 VDD1.n136 B 0.011672f
C820 VDD1.n137 B 0.012358f
C821 VDD1.n138 B 0.027588f
C822 VDD1.n139 B 0.027588f
C823 VDD1.n140 B 0.012358f
C824 VDD1.n141 B 0.011672f
C825 VDD1.n142 B 0.021721f
C826 VDD1.n143 B 0.021721f
C827 VDD1.n144 B 0.011672f
C828 VDD1.n145 B 0.012358f
C829 VDD1.n146 B 0.027588f
C830 VDD1.n147 B 0.027588f
C831 VDD1.n148 B 0.012358f
C832 VDD1.n149 B 0.011672f
C833 VDD1.n150 B 0.021721f
C834 VDD1.n151 B 0.021721f
C835 VDD1.n152 B 0.011672f
C836 VDD1.n153 B 0.012358f
C837 VDD1.n154 B 0.027588f
C838 VDD1.n155 B 0.027588f
C839 VDD1.n156 B 0.012358f
C840 VDD1.n157 B 0.011672f
C841 VDD1.n158 B 0.021721f
C842 VDD1.n159 B 0.021721f
C843 VDD1.n160 B 0.011672f
C844 VDD1.n161 B 0.012358f
C845 VDD1.n162 B 0.027588f
C846 VDD1.n163 B 0.027588f
C847 VDD1.n164 B 0.012358f
C848 VDD1.n165 B 0.011672f
C849 VDD1.n166 B 0.021721f
C850 VDD1.n167 B 0.021721f
C851 VDD1.n168 B 0.011672f
C852 VDD1.n169 B 0.012358f
C853 VDD1.n170 B 0.027588f
C854 VDD1.n171 B 0.027588f
C855 VDD1.n172 B 0.012358f
C856 VDD1.n173 B 0.011672f
C857 VDD1.n174 B 0.021721f
C858 VDD1.n175 B 0.021721f
C859 VDD1.n176 B 0.011672f
C860 VDD1.n177 B 0.011672f
C861 VDD1.n178 B 0.012358f
C862 VDD1.n179 B 0.027588f
C863 VDD1.n180 B 0.027588f
C864 VDD1.n181 B 0.027588f
C865 VDD1.n182 B 0.012015f
C866 VDD1.n183 B 0.011672f
C867 VDD1.n184 B 0.021721f
C868 VDD1.n185 B 0.021721f
C869 VDD1.n186 B 0.011672f
C870 VDD1.n187 B 0.012358f
C871 VDD1.n188 B 0.027588f
C872 VDD1.n189 B 0.027588f
C873 VDD1.n190 B 0.012358f
C874 VDD1.n191 B 0.011672f
C875 VDD1.n192 B 0.021721f
C876 VDD1.n193 B 0.021721f
C877 VDD1.n194 B 0.011672f
C878 VDD1.n195 B 0.012358f
C879 VDD1.n196 B 0.027588f
C880 VDD1.n197 B 0.05765f
C881 VDD1.n198 B 0.012358f
C882 VDD1.n199 B 0.011672f
C883 VDD1.n200 B 0.047833f
C884 VDD1.n201 B 0.049623f
C885 VDD1.t5 B 0.311705f
C886 VDD1.t3 B 0.311705f
C887 VDD1.n202 B 2.84025f
C888 VDD1.n203 B 2.30933f
C889 VDD1.t2 B 0.311705f
C890 VDD1.t0 B 0.311705f
C891 VDD1.n204 B 2.83848f
C892 VDD1.n205 B 2.55191f
C893 VP.n0 B 0.032702f
C894 VP.t5 B 2.35262f
C895 VP.n1 B 0.058759f
C896 VP.n2 B 0.032702f
C897 VP.t1 B 2.35262f
C898 VP.n3 B 0.050813f
C899 VP.n4 B 0.032702f
C900 VP.t4 B 2.35262f
C901 VP.n5 B 0.058759f
C902 VP.t3 B 2.45384f
C903 VP.t0 B 2.35262f
C904 VP.n6 B 0.90385f
C905 VP.n7 B 0.897244f
C906 VP.n8 B 0.207072f
C907 VP.n9 B 0.032702f
C908 VP.n10 B 0.032375f
C909 VP.n11 B 0.050813f
C910 VP.n12 B 0.897228f
C911 VP.n13 B 1.71608f
C912 VP.t2 B 2.35262f
C913 VP.n14 B 0.897228f
C914 VP.n15 B 1.74026f
C915 VP.n16 B 0.032702f
C916 VP.n17 B 0.032702f
C917 VP.n18 B 0.032375f
C918 VP.n19 B 0.058759f
C919 VP.n20 B 0.859515f
C920 VP.n21 B 0.032702f
C921 VP.n22 B 0.032702f
C922 VP.n23 B 0.032702f
C923 VP.n24 B 0.032375f
C924 VP.n25 B 0.050813f
C925 VP.n26 B 0.897228f
C926 VP.n27 B 0.030141f
.ends

