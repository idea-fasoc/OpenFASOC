* NGSPICE file created from diff_pair_sample_0521.ext - technology: sky130A

.subckt diff_pair_sample_0521 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t7 VP.t0 VTAIL.t8 B.t4 sky130_fd_pr__nfet_01v8 ad=1.0362 pd=6.61 as=2.4492 ps=13.34 w=6.28 l=2.9
X1 VTAIL.t10 VP.t1 VDD1.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=2.4492 pd=13.34 as=1.0362 ps=6.61 w=6.28 l=2.9
X2 VTAIL.t6 VN.t0 VDD2.t7 B.t6 sky130_fd_pr__nfet_01v8 ad=2.4492 pd=13.34 as=1.0362 ps=6.61 w=6.28 l=2.9
X3 VDD2.t6 VN.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.0362 pd=6.61 as=2.4492 ps=13.34 w=6.28 l=2.9
X4 VDD1.t5 VP.t2 VTAIL.t13 B.t1 sky130_fd_pr__nfet_01v8 ad=1.0362 pd=6.61 as=1.0362 ps=6.61 w=6.28 l=2.9
X5 VTAIL.t7 VN.t2 VDD2.t5 B.t7 sky130_fd_pr__nfet_01v8 ad=2.4492 pd=13.34 as=1.0362 ps=6.61 w=6.28 l=2.9
X6 VDD1.t4 VP.t3 VTAIL.t12 B.t3 sky130_fd_pr__nfet_01v8 ad=1.0362 pd=6.61 as=1.0362 ps=6.61 w=6.28 l=2.9
X7 VDD2.t4 VN.t3 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.0362 pd=6.61 as=1.0362 ps=6.61 w=6.28 l=2.9
X8 B.t21 B.t19 B.t20 B.t13 sky130_fd_pr__nfet_01v8 ad=2.4492 pd=13.34 as=0 ps=0 w=6.28 l=2.9
X9 B.t18 B.t16 B.t17 B.t9 sky130_fd_pr__nfet_01v8 ad=2.4492 pd=13.34 as=0 ps=0 w=6.28 l=2.9
X10 VTAIL.t15 VP.t4 VDD1.t3 B.t5 sky130_fd_pr__nfet_01v8 ad=1.0362 pd=6.61 as=1.0362 ps=6.61 w=6.28 l=2.9
X11 VDD2.t3 VN.t4 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.0362 pd=6.61 as=2.4492 ps=13.34 w=6.28 l=2.9
X12 VTAIL.t5 VN.t5 VDD2.t2 B.t5 sky130_fd_pr__nfet_01v8 ad=1.0362 pd=6.61 as=1.0362 ps=6.61 w=6.28 l=2.9
X13 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=2.4492 pd=13.34 as=0 ps=0 w=6.28 l=2.9
X14 VTAIL.t11 VP.t5 VDD1.t2 B.t7 sky130_fd_pr__nfet_01v8 ad=2.4492 pd=13.34 as=1.0362 ps=6.61 w=6.28 l=2.9
X15 VTAIL.t14 VP.t6 VDD1.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=1.0362 pd=6.61 as=1.0362 ps=6.61 w=6.28 l=2.9
X16 VDD1.t0 VP.t7 VTAIL.t9 B.t0 sky130_fd_pr__nfet_01v8 ad=1.0362 pd=6.61 as=2.4492 ps=13.34 w=6.28 l=2.9
X17 VTAIL.t2 VN.t6 VDD2.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=1.0362 pd=6.61 as=1.0362 ps=6.61 w=6.28 l=2.9
X18 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=2.4492 pd=13.34 as=0 ps=0 w=6.28 l=2.9
X19 VDD2.t0 VN.t7 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.0362 pd=6.61 as=1.0362 ps=6.61 w=6.28 l=2.9
R0 VP.n19 VP.n16 161.3
R1 VP.n21 VP.n20 161.3
R2 VP.n22 VP.n15 161.3
R3 VP.n24 VP.n23 161.3
R4 VP.n25 VP.n14 161.3
R5 VP.n28 VP.n27 161.3
R6 VP.n29 VP.n13 161.3
R7 VP.n31 VP.n30 161.3
R8 VP.n32 VP.n12 161.3
R9 VP.n34 VP.n33 161.3
R10 VP.n35 VP.n11 161.3
R11 VP.n37 VP.n36 161.3
R12 VP.n38 VP.n10 161.3
R13 VP.n74 VP.n0 161.3
R14 VP.n73 VP.n72 161.3
R15 VP.n71 VP.n1 161.3
R16 VP.n70 VP.n69 161.3
R17 VP.n68 VP.n2 161.3
R18 VP.n67 VP.n66 161.3
R19 VP.n65 VP.n3 161.3
R20 VP.n64 VP.n63 161.3
R21 VP.n61 VP.n4 161.3
R22 VP.n60 VP.n59 161.3
R23 VP.n58 VP.n5 161.3
R24 VP.n57 VP.n56 161.3
R25 VP.n55 VP.n6 161.3
R26 VP.n53 VP.n52 161.3
R27 VP.n51 VP.n7 161.3
R28 VP.n50 VP.n49 161.3
R29 VP.n48 VP.n8 161.3
R30 VP.n47 VP.n46 161.3
R31 VP.n45 VP.n9 161.3
R32 VP.n44 VP.n43 161.3
R33 VP.n42 VP.n41 106.236
R34 VP.n76 VP.n75 106.236
R35 VP.n40 VP.n39 106.236
R36 VP.n17 VP.t1 86.0624
R37 VP.n60 VP.n5 56.5617
R38 VP.n24 VP.n15 56.5617
R39 VP.n18 VP.n17 55.9508
R40 VP.n42 VP.t5 52.1895
R41 VP.n54 VP.t2 52.1895
R42 VP.n62 VP.t6 52.1895
R43 VP.n75 VP.t0 52.1895
R44 VP.n39 VP.t7 52.1895
R45 VP.n26 VP.t4 52.1895
R46 VP.n18 VP.t3 52.1895
R47 VP.n41 VP.n40 47.9769
R48 VP.n49 VP.n48 42.5146
R49 VP.n69 VP.n68 42.5146
R50 VP.n33 VP.n32 42.5146
R51 VP.n48 VP.n47 38.6395
R52 VP.n69 VP.n1 38.6395
R53 VP.n33 VP.n11 38.6395
R54 VP.n43 VP.n9 24.5923
R55 VP.n47 VP.n9 24.5923
R56 VP.n49 VP.n7 24.5923
R57 VP.n53 VP.n7 24.5923
R58 VP.n56 VP.n55 24.5923
R59 VP.n56 VP.n5 24.5923
R60 VP.n61 VP.n60 24.5923
R61 VP.n63 VP.n61 24.5923
R62 VP.n67 VP.n3 24.5923
R63 VP.n68 VP.n67 24.5923
R64 VP.n73 VP.n1 24.5923
R65 VP.n74 VP.n73 24.5923
R66 VP.n37 VP.n11 24.5923
R67 VP.n38 VP.n37 24.5923
R68 VP.n25 VP.n24 24.5923
R69 VP.n27 VP.n25 24.5923
R70 VP.n31 VP.n13 24.5923
R71 VP.n32 VP.n31 24.5923
R72 VP.n20 VP.n19 24.5923
R73 VP.n20 VP.n15 24.5923
R74 VP.n55 VP.n54 17.9525
R75 VP.n63 VP.n62 17.9525
R76 VP.n27 VP.n26 17.9525
R77 VP.n19 VP.n18 17.9525
R78 VP.n54 VP.n53 6.6403
R79 VP.n62 VP.n3 6.6403
R80 VP.n26 VP.n13 6.6403
R81 VP.n17 VP.n16 4.9785
R82 VP.n43 VP.n42 4.67295
R83 VP.n75 VP.n74 4.67295
R84 VP.n39 VP.n38 4.67295
R85 VP.n40 VP.n10 0.278335
R86 VP.n44 VP.n41 0.278335
R87 VP.n76 VP.n0 0.278335
R88 VP.n21 VP.n16 0.189894
R89 VP.n22 VP.n21 0.189894
R90 VP.n23 VP.n22 0.189894
R91 VP.n23 VP.n14 0.189894
R92 VP.n28 VP.n14 0.189894
R93 VP.n29 VP.n28 0.189894
R94 VP.n30 VP.n29 0.189894
R95 VP.n30 VP.n12 0.189894
R96 VP.n34 VP.n12 0.189894
R97 VP.n35 VP.n34 0.189894
R98 VP.n36 VP.n35 0.189894
R99 VP.n36 VP.n10 0.189894
R100 VP.n45 VP.n44 0.189894
R101 VP.n46 VP.n45 0.189894
R102 VP.n46 VP.n8 0.189894
R103 VP.n50 VP.n8 0.189894
R104 VP.n51 VP.n50 0.189894
R105 VP.n52 VP.n51 0.189894
R106 VP.n52 VP.n6 0.189894
R107 VP.n57 VP.n6 0.189894
R108 VP.n58 VP.n57 0.189894
R109 VP.n59 VP.n58 0.189894
R110 VP.n59 VP.n4 0.189894
R111 VP.n64 VP.n4 0.189894
R112 VP.n65 VP.n64 0.189894
R113 VP.n66 VP.n65 0.189894
R114 VP.n66 VP.n2 0.189894
R115 VP.n70 VP.n2 0.189894
R116 VP.n71 VP.n70 0.189894
R117 VP.n72 VP.n71 0.189894
R118 VP.n72 VP.n0 0.189894
R119 VP VP.n76 0.153485
R120 VTAIL.n11 VTAIL.t10 51.5186
R121 VTAIL.n10 VTAIL.t4 51.5186
R122 VTAIL.n7 VTAIL.t7 51.5186
R123 VTAIL.n15 VTAIL.t0 51.5185
R124 VTAIL.n2 VTAIL.t6 51.5185
R125 VTAIL.n3 VTAIL.t8 51.5185
R126 VTAIL.n6 VTAIL.t11 51.5185
R127 VTAIL.n14 VTAIL.t9 51.5185
R128 VTAIL.n13 VTAIL.n12 48.3657
R129 VTAIL.n9 VTAIL.n8 48.3657
R130 VTAIL.n1 VTAIL.n0 48.3655
R131 VTAIL.n5 VTAIL.n4 48.3655
R132 VTAIL.n15 VTAIL.n14 20.5652
R133 VTAIL.n7 VTAIL.n6 20.5652
R134 VTAIL.n0 VTAIL.t3 3.15337
R135 VTAIL.n0 VTAIL.t5 3.15337
R136 VTAIL.n4 VTAIL.t13 3.15337
R137 VTAIL.n4 VTAIL.t14 3.15337
R138 VTAIL.n12 VTAIL.t12 3.15337
R139 VTAIL.n12 VTAIL.t15 3.15337
R140 VTAIL.n8 VTAIL.t1 3.15337
R141 VTAIL.n8 VTAIL.t2 3.15337
R142 VTAIL.n9 VTAIL.n7 2.78498
R143 VTAIL.n10 VTAIL.n9 2.78498
R144 VTAIL.n13 VTAIL.n11 2.78498
R145 VTAIL.n14 VTAIL.n13 2.78498
R146 VTAIL.n6 VTAIL.n5 2.78498
R147 VTAIL.n5 VTAIL.n3 2.78498
R148 VTAIL.n2 VTAIL.n1 2.78498
R149 VTAIL VTAIL.n15 2.72679
R150 VTAIL.n11 VTAIL.n10 0.470328
R151 VTAIL.n3 VTAIL.n2 0.470328
R152 VTAIL VTAIL.n1 0.0586897
R153 VDD1 VDD1.n0 66.495
R154 VDD1.n3 VDD1.n2 66.3812
R155 VDD1.n3 VDD1.n1 66.3812
R156 VDD1.n5 VDD1.n4 65.0444
R157 VDD1.n5 VDD1.n3 42.2423
R158 VDD1.n4 VDD1.t3 3.15337
R159 VDD1.n4 VDD1.t0 3.15337
R160 VDD1.n0 VDD1.t6 3.15337
R161 VDD1.n0 VDD1.t4 3.15337
R162 VDD1.n2 VDD1.t1 3.15337
R163 VDD1.n2 VDD1.t7 3.15337
R164 VDD1.n1 VDD1.t2 3.15337
R165 VDD1.n1 VDD1.t5 3.15337
R166 VDD1 VDD1.n5 1.33455
R167 B.n749 B.n748 585
R168 B.n750 B.n749 585
R169 B.n250 B.n132 585
R170 B.n249 B.n248 585
R171 B.n247 B.n246 585
R172 B.n245 B.n244 585
R173 B.n243 B.n242 585
R174 B.n241 B.n240 585
R175 B.n239 B.n238 585
R176 B.n237 B.n236 585
R177 B.n235 B.n234 585
R178 B.n233 B.n232 585
R179 B.n231 B.n230 585
R180 B.n229 B.n228 585
R181 B.n227 B.n226 585
R182 B.n225 B.n224 585
R183 B.n223 B.n222 585
R184 B.n221 B.n220 585
R185 B.n219 B.n218 585
R186 B.n217 B.n216 585
R187 B.n215 B.n214 585
R188 B.n213 B.n212 585
R189 B.n211 B.n210 585
R190 B.n209 B.n208 585
R191 B.n207 B.n206 585
R192 B.n205 B.n204 585
R193 B.n203 B.n202 585
R194 B.n201 B.n200 585
R195 B.n199 B.n198 585
R196 B.n197 B.n196 585
R197 B.n195 B.n194 585
R198 B.n193 B.n192 585
R199 B.n191 B.n190 585
R200 B.n189 B.n188 585
R201 B.n187 B.n186 585
R202 B.n184 B.n183 585
R203 B.n182 B.n181 585
R204 B.n180 B.n179 585
R205 B.n178 B.n177 585
R206 B.n176 B.n175 585
R207 B.n174 B.n173 585
R208 B.n172 B.n171 585
R209 B.n170 B.n169 585
R210 B.n168 B.n167 585
R211 B.n166 B.n165 585
R212 B.n164 B.n163 585
R213 B.n162 B.n161 585
R214 B.n160 B.n159 585
R215 B.n158 B.n157 585
R216 B.n156 B.n155 585
R217 B.n154 B.n153 585
R218 B.n152 B.n151 585
R219 B.n150 B.n149 585
R220 B.n148 B.n147 585
R221 B.n146 B.n145 585
R222 B.n144 B.n143 585
R223 B.n142 B.n141 585
R224 B.n140 B.n139 585
R225 B.n103 B.n102 585
R226 B.n753 B.n752 585
R227 B.n747 B.n133 585
R228 B.n133 B.n100 585
R229 B.n746 B.n99 585
R230 B.n757 B.n99 585
R231 B.n745 B.n98 585
R232 B.n758 B.n98 585
R233 B.n744 B.n97 585
R234 B.n759 B.n97 585
R235 B.n743 B.n742 585
R236 B.n742 B.n93 585
R237 B.n741 B.n92 585
R238 B.n765 B.n92 585
R239 B.n740 B.n91 585
R240 B.n766 B.n91 585
R241 B.n739 B.n90 585
R242 B.n767 B.n90 585
R243 B.n738 B.n737 585
R244 B.n737 B.n86 585
R245 B.n736 B.n85 585
R246 B.n773 B.n85 585
R247 B.n735 B.n84 585
R248 B.n774 B.n84 585
R249 B.n734 B.n83 585
R250 B.n775 B.n83 585
R251 B.n733 B.n732 585
R252 B.n732 B.n79 585
R253 B.n731 B.n78 585
R254 B.n781 B.n78 585
R255 B.n730 B.n77 585
R256 B.n782 B.n77 585
R257 B.n729 B.n76 585
R258 B.n783 B.n76 585
R259 B.n728 B.n727 585
R260 B.n727 B.n72 585
R261 B.n726 B.n71 585
R262 B.n789 B.n71 585
R263 B.n725 B.n70 585
R264 B.n790 B.n70 585
R265 B.n724 B.n69 585
R266 B.n791 B.n69 585
R267 B.n723 B.n722 585
R268 B.n722 B.n68 585
R269 B.n721 B.n64 585
R270 B.n797 B.n64 585
R271 B.n720 B.n63 585
R272 B.n798 B.n63 585
R273 B.n719 B.n62 585
R274 B.n799 B.n62 585
R275 B.n718 B.n717 585
R276 B.n717 B.n58 585
R277 B.n716 B.n57 585
R278 B.n805 B.n57 585
R279 B.n715 B.n56 585
R280 B.n806 B.n56 585
R281 B.n714 B.n55 585
R282 B.n807 B.n55 585
R283 B.n713 B.n712 585
R284 B.n712 B.n51 585
R285 B.n711 B.n50 585
R286 B.n813 B.n50 585
R287 B.n710 B.n49 585
R288 B.n814 B.n49 585
R289 B.n709 B.n48 585
R290 B.n815 B.n48 585
R291 B.n708 B.n707 585
R292 B.n707 B.n44 585
R293 B.n706 B.n43 585
R294 B.n821 B.n43 585
R295 B.n705 B.n42 585
R296 B.n822 B.n42 585
R297 B.n704 B.n41 585
R298 B.n823 B.n41 585
R299 B.n703 B.n702 585
R300 B.n702 B.n37 585
R301 B.n701 B.n36 585
R302 B.n829 B.n36 585
R303 B.n700 B.n35 585
R304 B.n830 B.n35 585
R305 B.n699 B.n34 585
R306 B.n831 B.n34 585
R307 B.n698 B.n697 585
R308 B.n697 B.n30 585
R309 B.n696 B.n29 585
R310 B.n837 B.n29 585
R311 B.n695 B.n28 585
R312 B.n838 B.n28 585
R313 B.n694 B.n27 585
R314 B.n839 B.n27 585
R315 B.n693 B.n692 585
R316 B.n692 B.n23 585
R317 B.n691 B.n22 585
R318 B.n845 B.n22 585
R319 B.n690 B.n21 585
R320 B.n846 B.n21 585
R321 B.n689 B.n20 585
R322 B.n847 B.n20 585
R323 B.n688 B.n687 585
R324 B.n687 B.n16 585
R325 B.n686 B.n15 585
R326 B.n853 B.n15 585
R327 B.n685 B.n14 585
R328 B.n854 B.n14 585
R329 B.n684 B.n13 585
R330 B.n855 B.n13 585
R331 B.n683 B.n682 585
R332 B.n682 B.n12 585
R333 B.n681 B.n680 585
R334 B.n681 B.n8 585
R335 B.n679 B.n7 585
R336 B.n862 B.n7 585
R337 B.n678 B.n6 585
R338 B.n863 B.n6 585
R339 B.n677 B.n5 585
R340 B.n864 B.n5 585
R341 B.n676 B.n675 585
R342 B.n675 B.n4 585
R343 B.n674 B.n251 585
R344 B.n674 B.n673 585
R345 B.n664 B.n252 585
R346 B.n253 B.n252 585
R347 B.n666 B.n665 585
R348 B.n667 B.n666 585
R349 B.n663 B.n258 585
R350 B.n258 B.n257 585
R351 B.n662 B.n661 585
R352 B.n661 B.n660 585
R353 B.n260 B.n259 585
R354 B.n261 B.n260 585
R355 B.n653 B.n652 585
R356 B.n654 B.n653 585
R357 B.n651 B.n266 585
R358 B.n266 B.n265 585
R359 B.n650 B.n649 585
R360 B.n649 B.n648 585
R361 B.n268 B.n267 585
R362 B.n269 B.n268 585
R363 B.n641 B.n640 585
R364 B.n642 B.n641 585
R365 B.n639 B.n274 585
R366 B.n274 B.n273 585
R367 B.n638 B.n637 585
R368 B.n637 B.n636 585
R369 B.n276 B.n275 585
R370 B.n277 B.n276 585
R371 B.n629 B.n628 585
R372 B.n630 B.n629 585
R373 B.n627 B.n282 585
R374 B.n282 B.n281 585
R375 B.n626 B.n625 585
R376 B.n625 B.n624 585
R377 B.n284 B.n283 585
R378 B.n285 B.n284 585
R379 B.n617 B.n616 585
R380 B.n618 B.n617 585
R381 B.n615 B.n290 585
R382 B.n290 B.n289 585
R383 B.n614 B.n613 585
R384 B.n613 B.n612 585
R385 B.n292 B.n291 585
R386 B.n293 B.n292 585
R387 B.n605 B.n604 585
R388 B.n606 B.n605 585
R389 B.n603 B.n297 585
R390 B.n301 B.n297 585
R391 B.n602 B.n601 585
R392 B.n601 B.n600 585
R393 B.n299 B.n298 585
R394 B.n300 B.n299 585
R395 B.n593 B.n592 585
R396 B.n594 B.n593 585
R397 B.n591 B.n306 585
R398 B.n306 B.n305 585
R399 B.n590 B.n589 585
R400 B.n589 B.n588 585
R401 B.n308 B.n307 585
R402 B.n309 B.n308 585
R403 B.n581 B.n580 585
R404 B.n582 B.n581 585
R405 B.n579 B.n314 585
R406 B.n314 B.n313 585
R407 B.n578 B.n577 585
R408 B.n577 B.n576 585
R409 B.n316 B.n315 585
R410 B.n569 B.n316 585
R411 B.n568 B.n567 585
R412 B.n570 B.n568 585
R413 B.n566 B.n321 585
R414 B.n321 B.n320 585
R415 B.n565 B.n564 585
R416 B.n564 B.n563 585
R417 B.n323 B.n322 585
R418 B.n324 B.n323 585
R419 B.n556 B.n555 585
R420 B.n557 B.n556 585
R421 B.n554 B.n329 585
R422 B.n329 B.n328 585
R423 B.n553 B.n552 585
R424 B.n552 B.n551 585
R425 B.n331 B.n330 585
R426 B.n332 B.n331 585
R427 B.n544 B.n543 585
R428 B.n545 B.n544 585
R429 B.n542 B.n337 585
R430 B.n337 B.n336 585
R431 B.n541 B.n540 585
R432 B.n540 B.n539 585
R433 B.n339 B.n338 585
R434 B.n340 B.n339 585
R435 B.n532 B.n531 585
R436 B.n533 B.n532 585
R437 B.n530 B.n345 585
R438 B.n345 B.n344 585
R439 B.n529 B.n528 585
R440 B.n528 B.n527 585
R441 B.n347 B.n346 585
R442 B.n348 B.n347 585
R443 B.n520 B.n519 585
R444 B.n521 B.n520 585
R445 B.n518 B.n353 585
R446 B.n353 B.n352 585
R447 B.n517 B.n516 585
R448 B.n516 B.n515 585
R449 B.n355 B.n354 585
R450 B.n356 B.n355 585
R451 B.n511 B.n510 585
R452 B.n359 B.n358 585
R453 B.n507 B.n506 585
R454 B.n508 B.n507 585
R455 B.n505 B.n388 585
R456 B.n504 B.n503 585
R457 B.n502 B.n501 585
R458 B.n500 B.n499 585
R459 B.n498 B.n497 585
R460 B.n496 B.n495 585
R461 B.n494 B.n493 585
R462 B.n492 B.n491 585
R463 B.n490 B.n489 585
R464 B.n488 B.n487 585
R465 B.n486 B.n485 585
R466 B.n484 B.n483 585
R467 B.n482 B.n481 585
R468 B.n480 B.n479 585
R469 B.n478 B.n477 585
R470 B.n476 B.n475 585
R471 B.n474 B.n473 585
R472 B.n472 B.n471 585
R473 B.n470 B.n469 585
R474 B.n468 B.n467 585
R475 B.n466 B.n465 585
R476 B.n464 B.n463 585
R477 B.n462 B.n461 585
R478 B.n460 B.n459 585
R479 B.n458 B.n457 585
R480 B.n456 B.n455 585
R481 B.n454 B.n453 585
R482 B.n452 B.n451 585
R483 B.n450 B.n449 585
R484 B.n448 B.n447 585
R485 B.n446 B.n445 585
R486 B.n443 B.n442 585
R487 B.n441 B.n440 585
R488 B.n439 B.n438 585
R489 B.n437 B.n436 585
R490 B.n435 B.n434 585
R491 B.n433 B.n432 585
R492 B.n431 B.n430 585
R493 B.n429 B.n428 585
R494 B.n427 B.n426 585
R495 B.n425 B.n424 585
R496 B.n423 B.n422 585
R497 B.n421 B.n420 585
R498 B.n419 B.n418 585
R499 B.n417 B.n416 585
R500 B.n415 B.n414 585
R501 B.n413 B.n412 585
R502 B.n411 B.n410 585
R503 B.n409 B.n408 585
R504 B.n407 B.n406 585
R505 B.n405 B.n404 585
R506 B.n403 B.n402 585
R507 B.n401 B.n400 585
R508 B.n399 B.n398 585
R509 B.n397 B.n396 585
R510 B.n395 B.n394 585
R511 B.n512 B.n357 585
R512 B.n357 B.n356 585
R513 B.n514 B.n513 585
R514 B.n515 B.n514 585
R515 B.n351 B.n350 585
R516 B.n352 B.n351 585
R517 B.n523 B.n522 585
R518 B.n522 B.n521 585
R519 B.n524 B.n349 585
R520 B.n349 B.n348 585
R521 B.n526 B.n525 585
R522 B.n527 B.n526 585
R523 B.n343 B.n342 585
R524 B.n344 B.n343 585
R525 B.n535 B.n534 585
R526 B.n534 B.n533 585
R527 B.n536 B.n341 585
R528 B.n341 B.n340 585
R529 B.n538 B.n537 585
R530 B.n539 B.n538 585
R531 B.n335 B.n334 585
R532 B.n336 B.n335 585
R533 B.n547 B.n546 585
R534 B.n546 B.n545 585
R535 B.n548 B.n333 585
R536 B.n333 B.n332 585
R537 B.n550 B.n549 585
R538 B.n551 B.n550 585
R539 B.n327 B.n326 585
R540 B.n328 B.n327 585
R541 B.n559 B.n558 585
R542 B.n558 B.n557 585
R543 B.n560 B.n325 585
R544 B.n325 B.n324 585
R545 B.n562 B.n561 585
R546 B.n563 B.n562 585
R547 B.n319 B.n318 585
R548 B.n320 B.n319 585
R549 B.n572 B.n571 585
R550 B.n571 B.n570 585
R551 B.n573 B.n317 585
R552 B.n569 B.n317 585
R553 B.n575 B.n574 585
R554 B.n576 B.n575 585
R555 B.n312 B.n311 585
R556 B.n313 B.n312 585
R557 B.n584 B.n583 585
R558 B.n583 B.n582 585
R559 B.n585 B.n310 585
R560 B.n310 B.n309 585
R561 B.n587 B.n586 585
R562 B.n588 B.n587 585
R563 B.n304 B.n303 585
R564 B.n305 B.n304 585
R565 B.n596 B.n595 585
R566 B.n595 B.n594 585
R567 B.n597 B.n302 585
R568 B.n302 B.n300 585
R569 B.n599 B.n598 585
R570 B.n600 B.n599 585
R571 B.n296 B.n295 585
R572 B.n301 B.n296 585
R573 B.n608 B.n607 585
R574 B.n607 B.n606 585
R575 B.n609 B.n294 585
R576 B.n294 B.n293 585
R577 B.n611 B.n610 585
R578 B.n612 B.n611 585
R579 B.n288 B.n287 585
R580 B.n289 B.n288 585
R581 B.n620 B.n619 585
R582 B.n619 B.n618 585
R583 B.n621 B.n286 585
R584 B.n286 B.n285 585
R585 B.n623 B.n622 585
R586 B.n624 B.n623 585
R587 B.n280 B.n279 585
R588 B.n281 B.n280 585
R589 B.n632 B.n631 585
R590 B.n631 B.n630 585
R591 B.n633 B.n278 585
R592 B.n278 B.n277 585
R593 B.n635 B.n634 585
R594 B.n636 B.n635 585
R595 B.n272 B.n271 585
R596 B.n273 B.n272 585
R597 B.n644 B.n643 585
R598 B.n643 B.n642 585
R599 B.n645 B.n270 585
R600 B.n270 B.n269 585
R601 B.n647 B.n646 585
R602 B.n648 B.n647 585
R603 B.n264 B.n263 585
R604 B.n265 B.n264 585
R605 B.n656 B.n655 585
R606 B.n655 B.n654 585
R607 B.n657 B.n262 585
R608 B.n262 B.n261 585
R609 B.n659 B.n658 585
R610 B.n660 B.n659 585
R611 B.n256 B.n255 585
R612 B.n257 B.n256 585
R613 B.n669 B.n668 585
R614 B.n668 B.n667 585
R615 B.n670 B.n254 585
R616 B.n254 B.n253 585
R617 B.n672 B.n671 585
R618 B.n673 B.n672 585
R619 B.n3 B.n0 585
R620 B.n4 B.n3 585
R621 B.n861 B.n1 585
R622 B.n862 B.n861 585
R623 B.n860 B.n859 585
R624 B.n860 B.n8 585
R625 B.n858 B.n9 585
R626 B.n12 B.n9 585
R627 B.n857 B.n856 585
R628 B.n856 B.n855 585
R629 B.n11 B.n10 585
R630 B.n854 B.n11 585
R631 B.n852 B.n851 585
R632 B.n853 B.n852 585
R633 B.n850 B.n17 585
R634 B.n17 B.n16 585
R635 B.n849 B.n848 585
R636 B.n848 B.n847 585
R637 B.n19 B.n18 585
R638 B.n846 B.n19 585
R639 B.n844 B.n843 585
R640 B.n845 B.n844 585
R641 B.n842 B.n24 585
R642 B.n24 B.n23 585
R643 B.n841 B.n840 585
R644 B.n840 B.n839 585
R645 B.n26 B.n25 585
R646 B.n838 B.n26 585
R647 B.n836 B.n835 585
R648 B.n837 B.n836 585
R649 B.n834 B.n31 585
R650 B.n31 B.n30 585
R651 B.n833 B.n832 585
R652 B.n832 B.n831 585
R653 B.n33 B.n32 585
R654 B.n830 B.n33 585
R655 B.n828 B.n827 585
R656 B.n829 B.n828 585
R657 B.n826 B.n38 585
R658 B.n38 B.n37 585
R659 B.n825 B.n824 585
R660 B.n824 B.n823 585
R661 B.n40 B.n39 585
R662 B.n822 B.n40 585
R663 B.n820 B.n819 585
R664 B.n821 B.n820 585
R665 B.n818 B.n45 585
R666 B.n45 B.n44 585
R667 B.n817 B.n816 585
R668 B.n816 B.n815 585
R669 B.n47 B.n46 585
R670 B.n814 B.n47 585
R671 B.n812 B.n811 585
R672 B.n813 B.n812 585
R673 B.n810 B.n52 585
R674 B.n52 B.n51 585
R675 B.n809 B.n808 585
R676 B.n808 B.n807 585
R677 B.n54 B.n53 585
R678 B.n806 B.n54 585
R679 B.n804 B.n803 585
R680 B.n805 B.n804 585
R681 B.n802 B.n59 585
R682 B.n59 B.n58 585
R683 B.n801 B.n800 585
R684 B.n800 B.n799 585
R685 B.n61 B.n60 585
R686 B.n798 B.n61 585
R687 B.n796 B.n795 585
R688 B.n797 B.n796 585
R689 B.n794 B.n65 585
R690 B.n68 B.n65 585
R691 B.n793 B.n792 585
R692 B.n792 B.n791 585
R693 B.n67 B.n66 585
R694 B.n790 B.n67 585
R695 B.n788 B.n787 585
R696 B.n789 B.n788 585
R697 B.n786 B.n73 585
R698 B.n73 B.n72 585
R699 B.n785 B.n784 585
R700 B.n784 B.n783 585
R701 B.n75 B.n74 585
R702 B.n782 B.n75 585
R703 B.n780 B.n779 585
R704 B.n781 B.n780 585
R705 B.n778 B.n80 585
R706 B.n80 B.n79 585
R707 B.n777 B.n776 585
R708 B.n776 B.n775 585
R709 B.n82 B.n81 585
R710 B.n774 B.n82 585
R711 B.n772 B.n771 585
R712 B.n773 B.n772 585
R713 B.n770 B.n87 585
R714 B.n87 B.n86 585
R715 B.n769 B.n768 585
R716 B.n768 B.n767 585
R717 B.n89 B.n88 585
R718 B.n766 B.n89 585
R719 B.n764 B.n763 585
R720 B.n765 B.n764 585
R721 B.n762 B.n94 585
R722 B.n94 B.n93 585
R723 B.n761 B.n760 585
R724 B.n760 B.n759 585
R725 B.n96 B.n95 585
R726 B.n758 B.n96 585
R727 B.n756 B.n755 585
R728 B.n757 B.n756 585
R729 B.n754 B.n101 585
R730 B.n101 B.n100 585
R731 B.n865 B.n864 585
R732 B.n863 B.n2 585
R733 B.n752 B.n101 530.939
R734 B.n749 B.n133 530.939
R735 B.n394 B.n355 530.939
R736 B.n510 B.n357 530.939
R737 B.n137 B.t16 260.647
R738 B.n134 B.t8 260.647
R739 B.n392 B.t12 260.647
R740 B.n389 B.t19 260.647
R741 B.n750 B.n131 256.663
R742 B.n750 B.n130 256.663
R743 B.n750 B.n129 256.663
R744 B.n750 B.n128 256.663
R745 B.n750 B.n127 256.663
R746 B.n750 B.n126 256.663
R747 B.n750 B.n125 256.663
R748 B.n750 B.n124 256.663
R749 B.n750 B.n123 256.663
R750 B.n750 B.n122 256.663
R751 B.n750 B.n121 256.663
R752 B.n750 B.n120 256.663
R753 B.n750 B.n119 256.663
R754 B.n750 B.n118 256.663
R755 B.n750 B.n117 256.663
R756 B.n750 B.n116 256.663
R757 B.n750 B.n115 256.663
R758 B.n750 B.n114 256.663
R759 B.n750 B.n113 256.663
R760 B.n750 B.n112 256.663
R761 B.n750 B.n111 256.663
R762 B.n750 B.n110 256.663
R763 B.n750 B.n109 256.663
R764 B.n750 B.n108 256.663
R765 B.n750 B.n107 256.663
R766 B.n750 B.n106 256.663
R767 B.n750 B.n105 256.663
R768 B.n750 B.n104 256.663
R769 B.n751 B.n750 256.663
R770 B.n509 B.n508 256.663
R771 B.n508 B.n360 256.663
R772 B.n508 B.n361 256.663
R773 B.n508 B.n362 256.663
R774 B.n508 B.n363 256.663
R775 B.n508 B.n364 256.663
R776 B.n508 B.n365 256.663
R777 B.n508 B.n366 256.663
R778 B.n508 B.n367 256.663
R779 B.n508 B.n368 256.663
R780 B.n508 B.n369 256.663
R781 B.n508 B.n370 256.663
R782 B.n508 B.n371 256.663
R783 B.n508 B.n372 256.663
R784 B.n508 B.n373 256.663
R785 B.n508 B.n374 256.663
R786 B.n508 B.n375 256.663
R787 B.n508 B.n376 256.663
R788 B.n508 B.n377 256.663
R789 B.n508 B.n378 256.663
R790 B.n508 B.n379 256.663
R791 B.n508 B.n380 256.663
R792 B.n508 B.n381 256.663
R793 B.n508 B.n382 256.663
R794 B.n508 B.n383 256.663
R795 B.n508 B.n384 256.663
R796 B.n508 B.n385 256.663
R797 B.n508 B.n386 256.663
R798 B.n508 B.n387 256.663
R799 B.n867 B.n866 256.663
R800 B.n139 B.n103 163.367
R801 B.n143 B.n142 163.367
R802 B.n147 B.n146 163.367
R803 B.n151 B.n150 163.367
R804 B.n155 B.n154 163.367
R805 B.n159 B.n158 163.367
R806 B.n163 B.n162 163.367
R807 B.n167 B.n166 163.367
R808 B.n171 B.n170 163.367
R809 B.n175 B.n174 163.367
R810 B.n179 B.n178 163.367
R811 B.n183 B.n182 163.367
R812 B.n188 B.n187 163.367
R813 B.n192 B.n191 163.367
R814 B.n196 B.n195 163.367
R815 B.n200 B.n199 163.367
R816 B.n204 B.n203 163.367
R817 B.n208 B.n207 163.367
R818 B.n212 B.n211 163.367
R819 B.n216 B.n215 163.367
R820 B.n220 B.n219 163.367
R821 B.n224 B.n223 163.367
R822 B.n228 B.n227 163.367
R823 B.n232 B.n231 163.367
R824 B.n236 B.n235 163.367
R825 B.n240 B.n239 163.367
R826 B.n244 B.n243 163.367
R827 B.n248 B.n247 163.367
R828 B.n749 B.n132 163.367
R829 B.n516 B.n355 163.367
R830 B.n516 B.n353 163.367
R831 B.n520 B.n353 163.367
R832 B.n520 B.n347 163.367
R833 B.n528 B.n347 163.367
R834 B.n528 B.n345 163.367
R835 B.n532 B.n345 163.367
R836 B.n532 B.n339 163.367
R837 B.n540 B.n339 163.367
R838 B.n540 B.n337 163.367
R839 B.n544 B.n337 163.367
R840 B.n544 B.n331 163.367
R841 B.n552 B.n331 163.367
R842 B.n552 B.n329 163.367
R843 B.n556 B.n329 163.367
R844 B.n556 B.n323 163.367
R845 B.n564 B.n323 163.367
R846 B.n564 B.n321 163.367
R847 B.n568 B.n321 163.367
R848 B.n568 B.n316 163.367
R849 B.n577 B.n316 163.367
R850 B.n577 B.n314 163.367
R851 B.n581 B.n314 163.367
R852 B.n581 B.n308 163.367
R853 B.n589 B.n308 163.367
R854 B.n589 B.n306 163.367
R855 B.n593 B.n306 163.367
R856 B.n593 B.n299 163.367
R857 B.n601 B.n299 163.367
R858 B.n601 B.n297 163.367
R859 B.n605 B.n297 163.367
R860 B.n605 B.n292 163.367
R861 B.n613 B.n292 163.367
R862 B.n613 B.n290 163.367
R863 B.n617 B.n290 163.367
R864 B.n617 B.n284 163.367
R865 B.n625 B.n284 163.367
R866 B.n625 B.n282 163.367
R867 B.n629 B.n282 163.367
R868 B.n629 B.n276 163.367
R869 B.n637 B.n276 163.367
R870 B.n637 B.n274 163.367
R871 B.n641 B.n274 163.367
R872 B.n641 B.n268 163.367
R873 B.n649 B.n268 163.367
R874 B.n649 B.n266 163.367
R875 B.n653 B.n266 163.367
R876 B.n653 B.n260 163.367
R877 B.n661 B.n260 163.367
R878 B.n661 B.n258 163.367
R879 B.n666 B.n258 163.367
R880 B.n666 B.n252 163.367
R881 B.n674 B.n252 163.367
R882 B.n675 B.n674 163.367
R883 B.n675 B.n5 163.367
R884 B.n6 B.n5 163.367
R885 B.n7 B.n6 163.367
R886 B.n681 B.n7 163.367
R887 B.n682 B.n681 163.367
R888 B.n682 B.n13 163.367
R889 B.n14 B.n13 163.367
R890 B.n15 B.n14 163.367
R891 B.n687 B.n15 163.367
R892 B.n687 B.n20 163.367
R893 B.n21 B.n20 163.367
R894 B.n22 B.n21 163.367
R895 B.n692 B.n22 163.367
R896 B.n692 B.n27 163.367
R897 B.n28 B.n27 163.367
R898 B.n29 B.n28 163.367
R899 B.n697 B.n29 163.367
R900 B.n697 B.n34 163.367
R901 B.n35 B.n34 163.367
R902 B.n36 B.n35 163.367
R903 B.n702 B.n36 163.367
R904 B.n702 B.n41 163.367
R905 B.n42 B.n41 163.367
R906 B.n43 B.n42 163.367
R907 B.n707 B.n43 163.367
R908 B.n707 B.n48 163.367
R909 B.n49 B.n48 163.367
R910 B.n50 B.n49 163.367
R911 B.n712 B.n50 163.367
R912 B.n712 B.n55 163.367
R913 B.n56 B.n55 163.367
R914 B.n57 B.n56 163.367
R915 B.n717 B.n57 163.367
R916 B.n717 B.n62 163.367
R917 B.n63 B.n62 163.367
R918 B.n64 B.n63 163.367
R919 B.n722 B.n64 163.367
R920 B.n722 B.n69 163.367
R921 B.n70 B.n69 163.367
R922 B.n71 B.n70 163.367
R923 B.n727 B.n71 163.367
R924 B.n727 B.n76 163.367
R925 B.n77 B.n76 163.367
R926 B.n78 B.n77 163.367
R927 B.n732 B.n78 163.367
R928 B.n732 B.n83 163.367
R929 B.n84 B.n83 163.367
R930 B.n85 B.n84 163.367
R931 B.n737 B.n85 163.367
R932 B.n737 B.n90 163.367
R933 B.n91 B.n90 163.367
R934 B.n92 B.n91 163.367
R935 B.n742 B.n92 163.367
R936 B.n742 B.n97 163.367
R937 B.n98 B.n97 163.367
R938 B.n99 B.n98 163.367
R939 B.n133 B.n99 163.367
R940 B.n507 B.n359 163.367
R941 B.n507 B.n388 163.367
R942 B.n503 B.n502 163.367
R943 B.n499 B.n498 163.367
R944 B.n495 B.n494 163.367
R945 B.n491 B.n490 163.367
R946 B.n487 B.n486 163.367
R947 B.n483 B.n482 163.367
R948 B.n479 B.n478 163.367
R949 B.n475 B.n474 163.367
R950 B.n471 B.n470 163.367
R951 B.n467 B.n466 163.367
R952 B.n463 B.n462 163.367
R953 B.n459 B.n458 163.367
R954 B.n455 B.n454 163.367
R955 B.n451 B.n450 163.367
R956 B.n447 B.n446 163.367
R957 B.n442 B.n441 163.367
R958 B.n438 B.n437 163.367
R959 B.n434 B.n433 163.367
R960 B.n430 B.n429 163.367
R961 B.n426 B.n425 163.367
R962 B.n422 B.n421 163.367
R963 B.n418 B.n417 163.367
R964 B.n414 B.n413 163.367
R965 B.n410 B.n409 163.367
R966 B.n406 B.n405 163.367
R967 B.n402 B.n401 163.367
R968 B.n398 B.n397 163.367
R969 B.n514 B.n357 163.367
R970 B.n514 B.n351 163.367
R971 B.n522 B.n351 163.367
R972 B.n522 B.n349 163.367
R973 B.n526 B.n349 163.367
R974 B.n526 B.n343 163.367
R975 B.n534 B.n343 163.367
R976 B.n534 B.n341 163.367
R977 B.n538 B.n341 163.367
R978 B.n538 B.n335 163.367
R979 B.n546 B.n335 163.367
R980 B.n546 B.n333 163.367
R981 B.n550 B.n333 163.367
R982 B.n550 B.n327 163.367
R983 B.n558 B.n327 163.367
R984 B.n558 B.n325 163.367
R985 B.n562 B.n325 163.367
R986 B.n562 B.n319 163.367
R987 B.n571 B.n319 163.367
R988 B.n571 B.n317 163.367
R989 B.n575 B.n317 163.367
R990 B.n575 B.n312 163.367
R991 B.n583 B.n312 163.367
R992 B.n583 B.n310 163.367
R993 B.n587 B.n310 163.367
R994 B.n587 B.n304 163.367
R995 B.n595 B.n304 163.367
R996 B.n595 B.n302 163.367
R997 B.n599 B.n302 163.367
R998 B.n599 B.n296 163.367
R999 B.n607 B.n296 163.367
R1000 B.n607 B.n294 163.367
R1001 B.n611 B.n294 163.367
R1002 B.n611 B.n288 163.367
R1003 B.n619 B.n288 163.367
R1004 B.n619 B.n286 163.367
R1005 B.n623 B.n286 163.367
R1006 B.n623 B.n280 163.367
R1007 B.n631 B.n280 163.367
R1008 B.n631 B.n278 163.367
R1009 B.n635 B.n278 163.367
R1010 B.n635 B.n272 163.367
R1011 B.n643 B.n272 163.367
R1012 B.n643 B.n270 163.367
R1013 B.n647 B.n270 163.367
R1014 B.n647 B.n264 163.367
R1015 B.n655 B.n264 163.367
R1016 B.n655 B.n262 163.367
R1017 B.n659 B.n262 163.367
R1018 B.n659 B.n256 163.367
R1019 B.n668 B.n256 163.367
R1020 B.n668 B.n254 163.367
R1021 B.n672 B.n254 163.367
R1022 B.n672 B.n3 163.367
R1023 B.n865 B.n3 163.367
R1024 B.n861 B.n2 163.367
R1025 B.n861 B.n860 163.367
R1026 B.n860 B.n9 163.367
R1027 B.n856 B.n9 163.367
R1028 B.n856 B.n11 163.367
R1029 B.n852 B.n11 163.367
R1030 B.n852 B.n17 163.367
R1031 B.n848 B.n17 163.367
R1032 B.n848 B.n19 163.367
R1033 B.n844 B.n19 163.367
R1034 B.n844 B.n24 163.367
R1035 B.n840 B.n24 163.367
R1036 B.n840 B.n26 163.367
R1037 B.n836 B.n26 163.367
R1038 B.n836 B.n31 163.367
R1039 B.n832 B.n31 163.367
R1040 B.n832 B.n33 163.367
R1041 B.n828 B.n33 163.367
R1042 B.n828 B.n38 163.367
R1043 B.n824 B.n38 163.367
R1044 B.n824 B.n40 163.367
R1045 B.n820 B.n40 163.367
R1046 B.n820 B.n45 163.367
R1047 B.n816 B.n45 163.367
R1048 B.n816 B.n47 163.367
R1049 B.n812 B.n47 163.367
R1050 B.n812 B.n52 163.367
R1051 B.n808 B.n52 163.367
R1052 B.n808 B.n54 163.367
R1053 B.n804 B.n54 163.367
R1054 B.n804 B.n59 163.367
R1055 B.n800 B.n59 163.367
R1056 B.n800 B.n61 163.367
R1057 B.n796 B.n61 163.367
R1058 B.n796 B.n65 163.367
R1059 B.n792 B.n65 163.367
R1060 B.n792 B.n67 163.367
R1061 B.n788 B.n67 163.367
R1062 B.n788 B.n73 163.367
R1063 B.n784 B.n73 163.367
R1064 B.n784 B.n75 163.367
R1065 B.n780 B.n75 163.367
R1066 B.n780 B.n80 163.367
R1067 B.n776 B.n80 163.367
R1068 B.n776 B.n82 163.367
R1069 B.n772 B.n82 163.367
R1070 B.n772 B.n87 163.367
R1071 B.n768 B.n87 163.367
R1072 B.n768 B.n89 163.367
R1073 B.n764 B.n89 163.367
R1074 B.n764 B.n94 163.367
R1075 B.n760 B.n94 163.367
R1076 B.n760 B.n96 163.367
R1077 B.n756 B.n96 163.367
R1078 B.n756 B.n101 163.367
R1079 B.n134 B.t10 135.042
R1080 B.n392 B.t15 135.042
R1081 B.n137 B.t17 135.035
R1082 B.n389 B.t21 135.035
R1083 B.n508 B.n356 124.709
R1084 B.n750 B.n100 124.709
R1085 B.n135 B.t11 72.399
R1086 B.n393 B.t14 72.399
R1087 B.n138 B.t18 72.3922
R1088 B.n390 B.t20 72.3922
R1089 B.n752 B.n751 71.676
R1090 B.n139 B.n104 71.676
R1091 B.n143 B.n105 71.676
R1092 B.n147 B.n106 71.676
R1093 B.n151 B.n107 71.676
R1094 B.n155 B.n108 71.676
R1095 B.n159 B.n109 71.676
R1096 B.n163 B.n110 71.676
R1097 B.n167 B.n111 71.676
R1098 B.n171 B.n112 71.676
R1099 B.n175 B.n113 71.676
R1100 B.n179 B.n114 71.676
R1101 B.n183 B.n115 71.676
R1102 B.n188 B.n116 71.676
R1103 B.n192 B.n117 71.676
R1104 B.n196 B.n118 71.676
R1105 B.n200 B.n119 71.676
R1106 B.n204 B.n120 71.676
R1107 B.n208 B.n121 71.676
R1108 B.n212 B.n122 71.676
R1109 B.n216 B.n123 71.676
R1110 B.n220 B.n124 71.676
R1111 B.n224 B.n125 71.676
R1112 B.n228 B.n126 71.676
R1113 B.n232 B.n127 71.676
R1114 B.n236 B.n128 71.676
R1115 B.n240 B.n129 71.676
R1116 B.n244 B.n130 71.676
R1117 B.n248 B.n131 71.676
R1118 B.n132 B.n131 71.676
R1119 B.n247 B.n130 71.676
R1120 B.n243 B.n129 71.676
R1121 B.n239 B.n128 71.676
R1122 B.n235 B.n127 71.676
R1123 B.n231 B.n126 71.676
R1124 B.n227 B.n125 71.676
R1125 B.n223 B.n124 71.676
R1126 B.n219 B.n123 71.676
R1127 B.n215 B.n122 71.676
R1128 B.n211 B.n121 71.676
R1129 B.n207 B.n120 71.676
R1130 B.n203 B.n119 71.676
R1131 B.n199 B.n118 71.676
R1132 B.n195 B.n117 71.676
R1133 B.n191 B.n116 71.676
R1134 B.n187 B.n115 71.676
R1135 B.n182 B.n114 71.676
R1136 B.n178 B.n113 71.676
R1137 B.n174 B.n112 71.676
R1138 B.n170 B.n111 71.676
R1139 B.n166 B.n110 71.676
R1140 B.n162 B.n109 71.676
R1141 B.n158 B.n108 71.676
R1142 B.n154 B.n107 71.676
R1143 B.n150 B.n106 71.676
R1144 B.n146 B.n105 71.676
R1145 B.n142 B.n104 71.676
R1146 B.n751 B.n103 71.676
R1147 B.n510 B.n509 71.676
R1148 B.n388 B.n360 71.676
R1149 B.n502 B.n361 71.676
R1150 B.n498 B.n362 71.676
R1151 B.n494 B.n363 71.676
R1152 B.n490 B.n364 71.676
R1153 B.n486 B.n365 71.676
R1154 B.n482 B.n366 71.676
R1155 B.n478 B.n367 71.676
R1156 B.n474 B.n368 71.676
R1157 B.n470 B.n369 71.676
R1158 B.n466 B.n370 71.676
R1159 B.n462 B.n371 71.676
R1160 B.n458 B.n372 71.676
R1161 B.n454 B.n373 71.676
R1162 B.n450 B.n374 71.676
R1163 B.n446 B.n375 71.676
R1164 B.n441 B.n376 71.676
R1165 B.n437 B.n377 71.676
R1166 B.n433 B.n378 71.676
R1167 B.n429 B.n379 71.676
R1168 B.n425 B.n380 71.676
R1169 B.n421 B.n381 71.676
R1170 B.n417 B.n382 71.676
R1171 B.n413 B.n383 71.676
R1172 B.n409 B.n384 71.676
R1173 B.n405 B.n385 71.676
R1174 B.n401 B.n386 71.676
R1175 B.n397 B.n387 71.676
R1176 B.n509 B.n359 71.676
R1177 B.n503 B.n360 71.676
R1178 B.n499 B.n361 71.676
R1179 B.n495 B.n362 71.676
R1180 B.n491 B.n363 71.676
R1181 B.n487 B.n364 71.676
R1182 B.n483 B.n365 71.676
R1183 B.n479 B.n366 71.676
R1184 B.n475 B.n367 71.676
R1185 B.n471 B.n368 71.676
R1186 B.n467 B.n369 71.676
R1187 B.n463 B.n370 71.676
R1188 B.n459 B.n371 71.676
R1189 B.n455 B.n372 71.676
R1190 B.n451 B.n373 71.676
R1191 B.n447 B.n374 71.676
R1192 B.n442 B.n375 71.676
R1193 B.n438 B.n376 71.676
R1194 B.n434 B.n377 71.676
R1195 B.n430 B.n378 71.676
R1196 B.n426 B.n379 71.676
R1197 B.n422 B.n380 71.676
R1198 B.n418 B.n381 71.676
R1199 B.n414 B.n382 71.676
R1200 B.n410 B.n383 71.676
R1201 B.n406 B.n384 71.676
R1202 B.n402 B.n385 71.676
R1203 B.n398 B.n386 71.676
R1204 B.n394 B.n387 71.676
R1205 B.n866 B.n865 71.676
R1206 B.n866 B.n2 71.676
R1207 B.n515 B.n356 64.7344
R1208 B.n515 B.n352 64.7344
R1209 B.n521 B.n352 64.7344
R1210 B.n521 B.n348 64.7344
R1211 B.n527 B.n348 64.7344
R1212 B.n527 B.n344 64.7344
R1213 B.n533 B.n344 64.7344
R1214 B.n539 B.n340 64.7344
R1215 B.n539 B.n336 64.7344
R1216 B.n545 B.n336 64.7344
R1217 B.n545 B.n332 64.7344
R1218 B.n551 B.n332 64.7344
R1219 B.n551 B.n328 64.7344
R1220 B.n557 B.n328 64.7344
R1221 B.n557 B.n324 64.7344
R1222 B.n563 B.n324 64.7344
R1223 B.n563 B.n320 64.7344
R1224 B.n570 B.n320 64.7344
R1225 B.n570 B.n569 64.7344
R1226 B.n576 B.n313 64.7344
R1227 B.n582 B.n313 64.7344
R1228 B.n582 B.n309 64.7344
R1229 B.n588 B.n309 64.7344
R1230 B.n588 B.n305 64.7344
R1231 B.n594 B.n305 64.7344
R1232 B.n594 B.n300 64.7344
R1233 B.n600 B.n300 64.7344
R1234 B.n600 B.n301 64.7344
R1235 B.n606 B.n293 64.7344
R1236 B.n612 B.n293 64.7344
R1237 B.n612 B.n289 64.7344
R1238 B.n618 B.n289 64.7344
R1239 B.n618 B.n285 64.7344
R1240 B.n624 B.n285 64.7344
R1241 B.n624 B.n281 64.7344
R1242 B.n630 B.n281 64.7344
R1243 B.n636 B.n277 64.7344
R1244 B.n636 B.n273 64.7344
R1245 B.n642 B.n273 64.7344
R1246 B.n642 B.n269 64.7344
R1247 B.n648 B.n269 64.7344
R1248 B.n648 B.n265 64.7344
R1249 B.n654 B.n265 64.7344
R1250 B.n654 B.n261 64.7344
R1251 B.n660 B.n261 64.7344
R1252 B.n667 B.n257 64.7344
R1253 B.n667 B.n253 64.7344
R1254 B.n673 B.n253 64.7344
R1255 B.n673 B.n4 64.7344
R1256 B.n864 B.n4 64.7344
R1257 B.n864 B.n863 64.7344
R1258 B.n863 B.n862 64.7344
R1259 B.n862 B.n8 64.7344
R1260 B.n12 B.n8 64.7344
R1261 B.n855 B.n12 64.7344
R1262 B.n855 B.n854 64.7344
R1263 B.n853 B.n16 64.7344
R1264 B.n847 B.n16 64.7344
R1265 B.n847 B.n846 64.7344
R1266 B.n846 B.n845 64.7344
R1267 B.n845 B.n23 64.7344
R1268 B.n839 B.n23 64.7344
R1269 B.n839 B.n838 64.7344
R1270 B.n838 B.n837 64.7344
R1271 B.n837 B.n30 64.7344
R1272 B.n831 B.n830 64.7344
R1273 B.n830 B.n829 64.7344
R1274 B.n829 B.n37 64.7344
R1275 B.n823 B.n37 64.7344
R1276 B.n823 B.n822 64.7344
R1277 B.n822 B.n821 64.7344
R1278 B.n821 B.n44 64.7344
R1279 B.n815 B.n44 64.7344
R1280 B.n814 B.n813 64.7344
R1281 B.n813 B.n51 64.7344
R1282 B.n807 B.n51 64.7344
R1283 B.n807 B.n806 64.7344
R1284 B.n806 B.n805 64.7344
R1285 B.n805 B.n58 64.7344
R1286 B.n799 B.n58 64.7344
R1287 B.n799 B.n798 64.7344
R1288 B.n798 B.n797 64.7344
R1289 B.n791 B.n68 64.7344
R1290 B.n791 B.n790 64.7344
R1291 B.n790 B.n789 64.7344
R1292 B.n789 B.n72 64.7344
R1293 B.n783 B.n72 64.7344
R1294 B.n783 B.n782 64.7344
R1295 B.n782 B.n781 64.7344
R1296 B.n781 B.n79 64.7344
R1297 B.n775 B.n79 64.7344
R1298 B.n775 B.n774 64.7344
R1299 B.n774 B.n773 64.7344
R1300 B.n773 B.n86 64.7344
R1301 B.n767 B.n766 64.7344
R1302 B.n766 B.n765 64.7344
R1303 B.n765 B.n93 64.7344
R1304 B.n759 B.n93 64.7344
R1305 B.n759 B.n758 64.7344
R1306 B.n758 B.n757 64.7344
R1307 B.n757 B.n100 64.7344
R1308 B.n138 B.n137 62.6429
R1309 B.n135 B.n134 62.6429
R1310 B.n393 B.n392 62.6429
R1311 B.n390 B.n389 62.6429
R1312 B.n533 B.t13 60.9265
R1313 B.n767 B.t9 60.9265
R1314 B.n185 B.n138 59.5399
R1315 B.n136 B.n135 59.5399
R1316 B.n444 B.n393 59.5399
R1317 B.n391 B.n390 59.5399
R1318 B.n606 B.t1 55.2147
R1319 B.t4 B.n257 55.2147
R1320 B.n854 B.t6 55.2147
R1321 B.n815 B.t5 55.2147
R1322 B.n569 B.t7 41.8871
R1323 B.n630 B.t2 41.8871
R1324 B.n831 B.t3 41.8871
R1325 B.n68 B.t0 41.8871
R1326 B.n512 B.n511 34.4981
R1327 B.n395 B.n354 34.4981
R1328 B.n748 B.n747 34.4981
R1329 B.n754 B.n753 34.4981
R1330 B.n576 B.t7 22.8478
R1331 B.t2 B.n277 22.8478
R1332 B.t3 B.n30 22.8478
R1333 B.n797 B.t0 22.8478
R1334 B B.n867 18.0485
R1335 B.n513 B.n512 10.6151
R1336 B.n513 B.n350 10.6151
R1337 B.n523 B.n350 10.6151
R1338 B.n524 B.n523 10.6151
R1339 B.n525 B.n524 10.6151
R1340 B.n525 B.n342 10.6151
R1341 B.n535 B.n342 10.6151
R1342 B.n536 B.n535 10.6151
R1343 B.n537 B.n536 10.6151
R1344 B.n537 B.n334 10.6151
R1345 B.n547 B.n334 10.6151
R1346 B.n548 B.n547 10.6151
R1347 B.n549 B.n548 10.6151
R1348 B.n549 B.n326 10.6151
R1349 B.n559 B.n326 10.6151
R1350 B.n560 B.n559 10.6151
R1351 B.n561 B.n560 10.6151
R1352 B.n561 B.n318 10.6151
R1353 B.n572 B.n318 10.6151
R1354 B.n573 B.n572 10.6151
R1355 B.n574 B.n573 10.6151
R1356 B.n574 B.n311 10.6151
R1357 B.n584 B.n311 10.6151
R1358 B.n585 B.n584 10.6151
R1359 B.n586 B.n585 10.6151
R1360 B.n586 B.n303 10.6151
R1361 B.n596 B.n303 10.6151
R1362 B.n597 B.n596 10.6151
R1363 B.n598 B.n597 10.6151
R1364 B.n598 B.n295 10.6151
R1365 B.n608 B.n295 10.6151
R1366 B.n609 B.n608 10.6151
R1367 B.n610 B.n609 10.6151
R1368 B.n610 B.n287 10.6151
R1369 B.n620 B.n287 10.6151
R1370 B.n621 B.n620 10.6151
R1371 B.n622 B.n621 10.6151
R1372 B.n622 B.n279 10.6151
R1373 B.n632 B.n279 10.6151
R1374 B.n633 B.n632 10.6151
R1375 B.n634 B.n633 10.6151
R1376 B.n634 B.n271 10.6151
R1377 B.n644 B.n271 10.6151
R1378 B.n645 B.n644 10.6151
R1379 B.n646 B.n645 10.6151
R1380 B.n646 B.n263 10.6151
R1381 B.n656 B.n263 10.6151
R1382 B.n657 B.n656 10.6151
R1383 B.n658 B.n657 10.6151
R1384 B.n658 B.n255 10.6151
R1385 B.n669 B.n255 10.6151
R1386 B.n670 B.n669 10.6151
R1387 B.n671 B.n670 10.6151
R1388 B.n671 B.n0 10.6151
R1389 B.n511 B.n358 10.6151
R1390 B.n506 B.n358 10.6151
R1391 B.n506 B.n505 10.6151
R1392 B.n505 B.n504 10.6151
R1393 B.n504 B.n501 10.6151
R1394 B.n501 B.n500 10.6151
R1395 B.n500 B.n497 10.6151
R1396 B.n497 B.n496 10.6151
R1397 B.n496 B.n493 10.6151
R1398 B.n493 B.n492 10.6151
R1399 B.n492 B.n489 10.6151
R1400 B.n489 B.n488 10.6151
R1401 B.n488 B.n485 10.6151
R1402 B.n485 B.n484 10.6151
R1403 B.n484 B.n481 10.6151
R1404 B.n481 B.n480 10.6151
R1405 B.n480 B.n477 10.6151
R1406 B.n477 B.n476 10.6151
R1407 B.n476 B.n473 10.6151
R1408 B.n473 B.n472 10.6151
R1409 B.n472 B.n469 10.6151
R1410 B.n469 B.n468 10.6151
R1411 B.n468 B.n465 10.6151
R1412 B.n465 B.n464 10.6151
R1413 B.n461 B.n460 10.6151
R1414 B.n460 B.n457 10.6151
R1415 B.n457 B.n456 10.6151
R1416 B.n456 B.n453 10.6151
R1417 B.n453 B.n452 10.6151
R1418 B.n452 B.n449 10.6151
R1419 B.n449 B.n448 10.6151
R1420 B.n448 B.n445 10.6151
R1421 B.n443 B.n440 10.6151
R1422 B.n440 B.n439 10.6151
R1423 B.n439 B.n436 10.6151
R1424 B.n436 B.n435 10.6151
R1425 B.n435 B.n432 10.6151
R1426 B.n432 B.n431 10.6151
R1427 B.n431 B.n428 10.6151
R1428 B.n428 B.n427 10.6151
R1429 B.n427 B.n424 10.6151
R1430 B.n424 B.n423 10.6151
R1431 B.n423 B.n420 10.6151
R1432 B.n420 B.n419 10.6151
R1433 B.n419 B.n416 10.6151
R1434 B.n416 B.n415 10.6151
R1435 B.n415 B.n412 10.6151
R1436 B.n412 B.n411 10.6151
R1437 B.n411 B.n408 10.6151
R1438 B.n408 B.n407 10.6151
R1439 B.n407 B.n404 10.6151
R1440 B.n404 B.n403 10.6151
R1441 B.n403 B.n400 10.6151
R1442 B.n400 B.n399 10.6151
R1443 B.n399 B.n396 10.6151
R1444 B.n396 B.n395 10.6151
R1445 B.n517 B.n354 10.6151
R1446 B.n518 B.n517 10.6151
R1447 B.n519 B.n518 10.6151
R1448 B.n519 B.n346 10.6151
R1449 B.n529 B.n346 10.6151
R1450 B.n530 B.n529 10.6151
R1451 B.n531 B.n530 10.6151
R1452 B.n531 B.n338 10.6151
R1453 B.n541 B.n338 10.6151
R1454 B.n542 B.n541 10.6151
R1455 B.n543 B.n542 10.6151
R1456 B.n543 B.n330 10.6151
R1457 B.n553 B.n330 10.6151
R1458 B.n554 B.n553 10.6151
R1459 B.n555 B.n554 10.6151
R1460 B.n555 B.n322 10.6151
R1461 B.n565 B.n322 10.6151
R1462 B.n566 B.n565 10.6151
R1463 B.n567 B.n566 10.6151
R1464 B.n567 B.n315 10.6151
R1465 B.n578 B.n315 10.6151
R1466 B.n579 B.n578 10.6151
R1467 B.n580 B.n579 10.6151
R1468 B.n580 B.n307 10.6151
R1469 B.n590 B.n307 10.6151
R1470 B.n591 B.n590 10.6151
R1471 B.n592 B.n591 10.6151
R1472 B.n592 B.n298 10.6151
R1473 B.n602 B.n298 10.6151
R1474 B.n603 B.n602 10.6151
R1475 B.n604 B.n603 10.6151
R1476 B.n604 B.n291 10.6151
R1477 B.n614 B.n291 10.6151
R1478 B.n615 B.n614 10.6151
R1479 B.n616 B.n615 10.6151
R1480 B.n616 B.n283 10.6151
R1481 B.n626 B.n283 10.6151
R1482 B.n627 B.n626 10.6151
R1483 B.n628 B.n627 10.6151
R1484 B.n628 B.n275 10.6151
R1485 B.n638 B.n275 10.6151
R1486 B.n639 B.n638 10.6151
R1487 B.n640 B.n639 10.6151
R1488 B.n640 B.n267 10.6151
R1489 B.n650 B.n267 10.6151
R1490 B.n651 B.n650 10.6151
R1491 B.n652 B.n651 10.6151
R1492 B.n652 B.n259 10.6151
R1493 B.n662 B.n259 10.6151
R1494 B.n663 B.n662 10.6151
R1495 B.n665 B.n663 10.6151
R1496 B.n665 B.n664 10.6151
R1497 B.n664 B.n251 10.6151
R1498 B.n676 B.n251 10.6151
R1499 B.n677 B.n676 10.6151
R1500 B.n678 B.n677 10.6151
R1501 B.n679 B.n678 10.6151
R1502 B.n680 B.n679 10.6151
R1503 B.n683 B.n680 10.6151
R1504 B.n684 B.n683 10.6151
R1505 B.n685 B.n684 10.6151
R1506 B.n686 B.n685 10.6151
R1507 B.n688 B.n686 10.6151
R1508 B.n689 B.n688 10.6151
R1509 B.n690 B.n689 10.6151
R1510 B.n691 B.n690 10.6151
R1511 B.n693 B.n691 10.6151
R1512 B.n694 B.n693 10.6151
R1513 B.n695 B.n694 10.6151
R1514 B.n696 B.n695 10.6151
R1515 B.n698 B.n696 10.6151
R1516 B.n699 B.n698 10.6151
R1517 B.n700 B.n699 10.6151
R1518 B.n701 B.n700 10.6151
R1519 B.n703 B.n701 10.6151
R1520 B.n704 B.n703 10.6151
R1521 B.n705 B.n704 10.6151
R1522 B.n706 B.n705 10.6151
R1523 B.n708 B.n706 10.6151
R1524 B.n709 B.n708 10.6151
R1525 B.n710 B.n709 10.6151
R1526 B.n711 B.n710 10.6151
R1527 B.n713 B.n711 10.6151
R1528 B.n714 B.n713 10.6151
R1529 B.n715 B.n714 10.6151
R1530 B.n716 B.n715 10.6151
R1531 B.n718 B.n716 10.6151
R1532 B.n719 B.n718 10.6151
R1533 B.n720 B.n719 10.6151
R1534 B.n721 B.n720 10.6151
R1535 B.n723 B.n721 10.6151
R1536 B.n724 B.n723 10.6151
R1537 B.n725 B.n724 10.6151
R1538 B.n726 B.n725 10.6151
R1539 B.n728 B.n726 10.6151
R1540 B.n729 B.n728 10.6151
R1541 B.n730 B.n729 10.6151
R1542 B.n731 B.n730 10.6151
R1543 B.n733 B.n731 10.6151
R1544 B.n734 B.n733 10.6151
R1545 B.n735 B.n734 10.6151
R1546 B.n736 B.n735 10.6151
R1547 B.n738 B.n736 10.6151
R1548 B.n739 B.n738 10.6151
R1549 B.n740 B.n739 10.6151
R1550 B.n741 B.n740 10.6151
R1551 B.n743 B.n741 10.6151
R1552 B.n744 B.n743 10.6151
R1553 B.n745 B.n744 10.6151
R1554 B.n746 B.n745 10.6151
R1555 B.n747 B.n746 10.6151
R1556 B.n859 B.n1 10.6151
R1557 B.n859 B.n858 10.6151
R1558 B.n858 B.n857 10.6151
R1559 B.n857 B.n10 10.6151
R1560 B.n851 B.n10 10.6151
R1561 B.n851 B.n850 10.6151
R1562 B.n850 B.n849 10.6151
R1563 B.n849 B.n18 10.6151
R1564 B.n843 B.n18 10.6151
R1565 B.n843 B.n842 10.6151
R1566 B.n842 B.n841 10.6151
R1567 B.n841 B.n25 10.6151
R1568 B.n835 B.n25 10.6151
R1569 B.n835 B.n834 10.6151
R1570 B.n834 B.n833 10.6151
R1571 B.n833 B.n32 10.6151
R1572 B.n827 B.n32 10.6151
R1573 B.n827 B.n826 10.6151
R1574 B.n826 B.n825 10.6151
R1575 B.n825 B.n39 10.6151
R1576 B.n819 B.n39 10.6151
R1577 B.n819 B.n818 10.6151
R1578 B.n818 B.n817 10.6151
R1579 B.n817 B.n46 10.6151
R1580 B.n811 B.n46 10.6151
R1581 B.n811 B.n810 10.6151
R1582 B.n810 B.n809 10.6151
R1583 B.n809 B.n53 10.6151
R1584 B.n803 B.n53 10.6151
R1585 B.n803 B.n802 10.6151
R1586 B.n802 B.n801 10.6151
R1587 B.n801 B.n60 10.6151
R1588 B.n795 B.n60 10.6151
R1589 B.n795 B.n794 10.6151
R1590 B.n794 B.n793 10.6151
R1591 B.n793 B.n66 10.6151
R1592 B.n787 B.n66 10.6151
R1593 B.n787 B.n786 10.6151
R1594 B.n786 B.n785 10.6151
R1595 B.n785 B.n74 10.6151
R1596 B.n779 B.n74 10.6151
R1597 B.n779 B.n778 10.6151
R1598 B.n778 B.n777 10.6151
R1599 B.n777 B.n81 10.6151
R1600 B.n771 B.n81 10.6151
R1601 B.n771 B.n770 10.6151
R1602 B.n770 B.n769 10.6151
R1603 B.n769 B.n88 10.6151
R1604 B.n763 B.n88 10.6151
R1605 B.n763 B.n762 10.6151
R1606 B.n762 B.n761 10.6151
R1607 B.n761 B.n95 10.6151
R1608 B.n755 B.n95 10.6151
R1609 B.n755 B.n754 10.6151
R1610 B.n753 B.n102 10.6151
R1611 B.n140 B.n102 10.6151
R1612 B.n141 B.n140 10.6151
R1613 B.n144 B.n141 10.6151
R1614 B.n145 B.n144 10.6151
R1615 B.n148 B.n145 10.6151
R1616 B.n149 B.n148 10.6151
R1617 B.n152 B.n149 10.6151
R1618 B.n153 B.n152 10.6151
R1619 B.n156 B.n153 10.6151
R1620 B.n157 B.n156 10.6151
R1621 B.n160 B.n157 10.6151
R1622 B.n161 B.n160 10.6151
R1623 B.n164 B.n161 10.6151
R1624 B.n165 B.n164 10.6151
R1625 B.n168 B.n165 10.6151
R1626 B.n169 B.n168 10.6151
R1627 B.n172 B.n169 10.6151
R1628 B.n173 B.n172 10.6151
R1629 B.n176 B.n173 10.6151
R1630 B.n177 B.n176 10.6151
R1631 B.n180 B.n177 10.6151
R1632 B.n181 B.n180 10.6151
R1633 B.n184 B.n181 10.6151
R1634 B.n189 B.n186 10.6151
R1635 B.n190 B.n189 10.6151
R1636 B.n193 B.n190 10.6151
R1637 B.n194 B.n193 10.6151
R1638 B.n197 B.n194 10.6151
R1639 B.n198 B.n197 10.6151
R1640 B.n201 B.n198 10.6151
R1641 B.n202 B.n201 10.6151
R1642 B.n206 B.n205 10.6151
R1643 B.n209 B.n206 10.6151
R1644 B.n210 B.n209 10.6151
R1645 B.n213 B.n210 10.6151
R1646 B.n214 B.n213 10.6151
R1647 B.n217 B.n214 10.6151
R1648 B.n218 B.n217 10.6151
R1649 B.n221 B.n218 10.6151
R1650 B.n222 B.n221 10.6151
R1651 B.n225 B.n222 10.6151
R1652 B.n226 B.n225 10.6151
R1653 B.n229 B.n226 10.6151
R1654 B.n230 B.n229 10.6151
R1655 B.n233 B.n230 10.6151
R1656 B.n234 B.n233 10.6151
R1657 B.n237 B.n234 10.6151
R1658 B.n238 B.n237 10.6151
R1659 B.n241 B.n238 10.6151
R1660 B.n242 B.n241 10.6151
R1661 B.n245 B.n242 10.6151
R1662 B.n246 B.n245 10.6151
R1663 B.n249 B.n246 10.6151
R1664 B.n250 B.n249 10.6151
R1665 B.n748 B.n250 10.6151
R1666 B.n301 B.t1 9.52019
R1667 B.n660 B.t4 9.52019
R1668 B.t6 B.n853 9.52019
R1669 B.t5 B.n814 9.52019
R1670 B.n867 B.n0 8.11757
R1671 B.n867 B.n1 8.11757
R1672 B.n461 B.n391 6.5566
R1673 B.n445 B.n444 6.5566
R1674 B.n186 B.n185 6.5566
R1675 B.n202 B.n136 6.5566
R1676 B.n464 B.n391 4.05904
R1677 B.n444 B.n443 4.05904
R1678 B.n185 B.n184 4.05904
R1679 B.n205 B.n136 4.05904
R1680 B.t13 B.n340 3.80838
R1681 B.t9 B.n86 3.80838
R1682 VN.n59 VN.n31 161.3
R1683 VN.n58 VN.n57 161.3
R1684 VN.n56 VN.n32 161.3
R1685 VN.n55 VN.n54 161.3
R1686 VN.n53 VN.n33 161.3
R1687 VN.n52 VN.n51 161.3
R1688 VN.n50 VN.n34 161.3
R1689 VN.n49 VN.n48 161.3
R1690 VN.n47 VN.n35 161.3
R1691 VN.n46 VN.n45 161.3
R1692 VN.n44 VN.n37 161.3
R1693 VN.n43 VN.n42 161.3
R1694 VN.n41 VN.n38 161.3
R1695 VN.n28 VN.n0 161.3
R1696 VN.n27 VN.n26 161.3
R1697 VN.n25 VN.n1 161.3
R1698 VN.n24 VN.n23 161.3
R1699 VN.n22 VN.n2 161.3
R1700 VN.n21 VN.n20 161.3
R1701 VN.n19 VN.n3 161.3
R1702 VN.n18 VN.n17 161.3
R1703 VN.n15 VN.n4 161.3
R1704 VN.n14 VN.n13 161.3
R1705 VN.n12 VN.n5 161.3
R1706 VN.n11 VN.n10 161.3
R1707 VN.n9 VN.n6 161.3
R1708 VN.n30 VN.n29 106.236
R1709 VN.n61 VN.n60 106.236
R1710 VN.n7 VN.t0 86.0624
R1711 VN.n39 VN.t4 86.0624
R1712 VN.n14 VN.n5 56.5617
R1713 VN.n46 VN.n37 56.5617
R1714 VN.n8 VN.n7 55.9508
R1715 VN.n40 VN.n39 55.9508
R1716 VN.n8 VN.t7 52.1895
R1717 VN.n16 VN.t5 52.1895
R1718 VN.n29 VN.t1 52.1895
R1719 VN.n40 VN.t6 52.1895
R1720 VN.n36 VN.t3 52.1895
R1721 VN.n60 VN.t2 52.1895
R1722 VN VN.n61 48.2558
R1723 VN.n23 VN.n22 42.5146
R1724 VN.n54 VN.n53 42.5146
R1725 VN.n23 VN.n1 38.6395
R1726 VN.n54 VN.n32 38.6395
R1727 VN.n10 VN.n9 24.5923
R1728 VN.n10 VN.n5 24.5923
R1729 VN.n15 VN.n14 24.5923
R1730 VN.n17 VN.n15 24.5923
R1731 VN.n21 VN.n3 24.5923
R1732 VN.n22 VN.n21 24.5923
R1733 VN.n27 VN.n1 24.5923
R1734 VN.n28 VN.n27 24.5923
R1735 VN.n42 VN.n37 24.5923
R1736 VN.n42 VN.n41 24.5923
R1737 VN.n53 VN.n52 24.5923
R1738 VN.n52 VN.n34 24.5923
R1739 VN.n48 VN.n47 24.5923
R1740 VN.n47 VN.n46 24.5923
R1741 VN.n59 VN.n58 24.5923
R1742 VN.n58 VN.n32 24.5923
R1743 VN.n9 VN.n8 17.9525
R1744 VN.n17 VN.n16 17.9525
R1745 VN.n41 VN.n40 17.9525
R1746 VN.n48 VN.n36 17.9525
R1747 VN.n16 VN.n3 6.6403
R1748 VN.n36 VN.n34 6.6403
R1749 VN.n39 VN.n38 4.9785
R1750 VN.n7 VN.n6 4.9785
R1751 VN.n29 VN.n28 4.67295
R1752 VN.n60 VN.n59 4.67295
R1753 VN.n61 VN.n31 0.278335
R1754 VN.n30 VN.n0 0.278335
R1755 VN.n57 VN.n31 0.189894
R1756 VN.n57 VN.n56 0.189894
R1757 VN.n56 VN.n55 0.189894
R1758 VN.n55 VN.n33 0.189894
R1759 VN.n51 VN.n33 0.189894
R1760 VN.n51 VN.n50 0.189894
R1761 VN.n50 VN.n49 0.189894
R1762 VN.n49 VN.n35 0.189894
R1763 VN.n45 VN.n35 0.189894
R1764 VN.n45 VN.n44 0.189894
R1765 VN.n44 VN.n43 0.189894
R1766 VN.n43 VN.n38 0.189894
R1767 VN.n11 VN.n6 0.189894
R1768 VN.n12 VN.n11 0.189894
R1769 VN.n13 VN.n12 0.189894
R1770 VN.n13 VN.n4 0.189894
R1771 VN.n18 VN.n4 0.189894
R1772 VN.n19 VN.n18 0.189894
R1773 VN.n20 VN.n19 0.189894
R1774 VN.n20 VN.n2 0.189894
R1775 VN.n24 VN.n2 0.189894
R1776 VN.n25 VN.n24 0.189894
R1777 VN.n26 VN.n25 0.189894
R1778 VN.n26 VN.n0 0.189894
R1779 VN VN.n30 0.153485
R1780 VDD2.n2 VDD2.n1 66.3812
R1781 VDD2.n2 VDD2.n0 66.3812
R1782 VDD2 VDD2.n5 66.3784
R1783 VDD2.n4 VDD2.n3 65.0445
R1784 VDD2.n4 VDD2.n2 41.6593
R1785 VDD2.n5 VDD2.t1 3.15337
R1786 VDD2.n5 VDD2.t3 3.15337
R1787 VDD2.n3 VDD2.t5 3.15337
R1788 VDD2.n3 VDD2.t4 3.15337
R1789 VDD2.n1 VDD2.t2 3.15337
R1790 VDD2.n1 VDD2.t6 3.15337
R1791 VDD2.n0 VDD2.t7 3.15337
R1792 VDD2.n0 VDD2.t0 3.15337
R1793 VDD2 VDD2.n4 1.45093
C0 VDD1 VP 5.27009f
C1 VN VDD1 0.15219f
C2 VTAIL VDD2 6.39862f
C3 VN VP 6.96152f
C4 VTAIL VDD1 6.3422f
C5 VDD2 VDD1 1.93074f
C6 VTAIL VP 5.818181f
C7 VDD2 VP 0.551514f
C8 VTAIL VN 5.80408f
C9 VDD2 VN 4.87231f
C10 VDD2 B 5.179432f
C11 VDD1 B 5.652213f
C12 VTAIL B 6.850551f
C13 VN B 16.02875f
C14 VP B 14.658257f
C15 VDD2.t7 B 0.120317f
C16 VDD2.t0 B 0.120317f
C17 VDD2.n0 B 1.01889f
C18 VDD2.t2 B 0.120317f
C19 VDD2.t6 B 0.120317f
C20 VDD2.n1 B 1.01889f
C21 VDD2.n2 B 3.00236f
C22 VDD2.t5 B 0.120317f
C23 VDD2.t4 B 0.120317f
C24 VDD2.n3 B 1.00821f
C25 VDD2.n4 B 2.53355f
C26 VDD2.t1 B 0.120317f
C27 VDD2.t3 B 0.120317f
C28 VDD2.n5 B 1.01885f
C29 VN.n0 B 0.030639f
C30 VN.t1 B 1.12321f
C31 VN.n1 B 0.046346f
C32 VN.n2 B 0.023241f
C33 VN.n3 B 0.027566f
C34 VN.n4 B 0.023241f
C35 VN.n5 B 0.033784f
C36 VN.n6 B 0.246375f
C37 VN.t7 B 1.12321f
C38 VN.t0 B 1.34947f
C39 VN.n7 B 0.465399f
C40 VN.n8 B 0.493701f
C41 VN.n9 B 0.037353f
C42 VN.n10 B 0.043097f
C43 VN.n11 B 0.023241f
C44 VN.n12 B 0.023241f
C45 VN.n13 B 0.023241f
C46 VN.n14 B 0.033784f
C47 VN.n15 B 0.043097f
C48 VN.t5 B 1.12321f
C49 VN.n16 B 0.416664f
C50 VN.n17 B 0.037353f
C51 VN.n18 B 0.023241f
C52 VN.n19 B 0.023241f
C53 VN.n20 B 0.023241f
C54 VN.n21 B 0.043097f
C55 VN.n22 B 0.04543f
C56 VN.n23 B 0.018889f
C57 VN.n24 B 0.023241f
C58 VN.n25 B 0.023241f
C59 VN.n26 B 0.023241f
C60 VN.n27 B 0.043097f
C61 VN.n28 B 0.025864f
C62 VN.n29 B 0.496481f
C63 VN.n30 B 0.043298f
C64 VN.n31 B 0.030639f
C65 VN.t2 B 1.12321f
C66 VN.n32 B 0.046346f
C67 VN.n33 B 0.023241f
C68 VN.n34 B 0.027566f
C69 VN.n35 B 0.023241f
C70 VN.t3 B 1.12321f
C71 VN.n36 B 0.416664f
C72 VN.n37 B 0.033784f
C73 VN.n38 B 0.246375f
C74 VN.t6 B 1.12321f
C75 VN.t4 B 1.34947f
C76 VN.n39 B 0.465399f
C77 VN.n40 B 0.493701f
C78 VN.n41 B 0.037353f
C79 VN.n42 B 0.043097f
C80 VN.n43 B 0.023241f
C81 VN.n44 B 0.023241f
C82 VN.n45 B 0.023241f
C83 VN.n46 B 0.033784f
C84 VN.n47 B 0.043097f
C85 VN.n48 B 0.037353f
C86 VN.n49 B 0.023241f
C87 VN.n50 B 0.023241f
C88 VN.n51 B 0.023241f
C89 VN.n52 B 0.043097f
C90 VN.n53 B 0.04543f
C91 VN.n54 B 0.018889f
C92 VN.n55 B 0.023241f
C93 VN.n56 B 0.023241f
C94 VN.n57 B 0.023241f
C95 VN.n58 B 0.043097f
C96 VN.n59 B 0.025864f
C97 VN.n60 B 0.496481f
C98 VN.n61 B 1.23476f
C99 VDD1.t6 B 0.12254f
C100 VDD1.t4 B 0.12254f
C101 VDD1.n0 B 1.03881f
C102 VDD1.t2 B 0.12254f
C103 VDD1.t5 B 0.12254f
C104 VDD1.n1 B 1.03771f
C105 VDD1.t1 B 0.12254f
C106 VDD1.t7 B 0.12254f
C107 VDD1.n2 B 1.03771f
C108 VDD1.n3 B 3.10927f
C109 VDD1.t3 B 0.12254f
C110 VDD1.t0 B 0.12254f
C111 VDD1.n4 B 1.02683f
C112 VDD1.n5 B 2.61088f
C113 VTAIL.t3 B 0.116126f
C114 VTAIL.t5 B 0.116126f
C115 VTAIL.n0 B 0.908614f
C116 VTAIL.n1 B 0.43842f
C117 VTAIL.t6 B 1.15744f
C118 VTAIL.n2 B 0.537341f
C119 VTAIL.t8 B 1.15744f
C120 VTAIL.n3 B 0.537341f
C121 VTAIL.t13 B 0.116126f
C122 VTAIL.t14 B 0.116126f
C123 VTAIL.n4 B 0.908614f
C124 VTAIL.n5 B 0.643984f
C125 VTAIL.t11 B 1.15744f
C126 VTAIL.n6 B 1.43793f
C127 VTAIL.t7 B 1.15745f
C128 VTAIL.n7 B 1.43792f
C129 VTAIL.t1 B 0.116126f
C130 VTAIL.t2 B 0.116126f
C131 VTAIL.n8 B 0.908619f
C132 VTAIL.n9 B 0.643978f
C133 VTAIL.t4 B 1.15745f
C134 VTAIL.n10 B 0.537334f
C135 VTAIL.t10 B 1.15745f
C136 VTAIL.n11 B 0.537334f
C137 VTAIL.t12 B 0.116126f
C138 VTAIL.t15 B 0.116126f
C139 VTAIL.n12 B 0.908619f
C140 VTAIL.n13 B 0.643978f
C141 VTAIL.t9 B 1.15744f
C142 VTAIL.n14 B 1.43793f
C143 VTAIL.t0 B 1.15744f
C144 VTAIL.n15 B 1.43354f
C145 VP.n0 B 0.031389f
C146 VP.t0 B 1.15071f
C147 VP.n1 B 0.047481f
C148 VP.n2 B 0.02381f
C149 VP.n3 B 0.028241f
C150 VP.n4 B 0.02381f
C151 VP.n5 B 0.034611f
C152 VP.n6 B 0.02381f
C153 VP.t2 B 1.15071f
C154 VP.n7 B 0.044153f
C155 VP.n8 B 0.02381f
C156 VP.n9 B 0.044153f
C157 VP.n10 B 0.031389f
C158 VP.t7 B 1.15071f
C159 VP.n11 B 0.047481f
C160 VP.n12 B 0.02381f
C161 VP.n13 B 0.028241f
C162 VP.n14 B 0.02381f
C163 VP.n15 B 0.034611f
C164 VP.n16 B 0.252409f
C165 VP.t3 B 1.15071f
C166 VP.t1 B 1.38252f
C167 VP.n17 B 0.476796f
C168 VP.n18 B 0.505791f
C169 VP.n19 B 0.038268f
C170 VP.n20 B 0.044153f
C171 VP.n21 B 0.02381f
C172 VP.n22 B 0.02381f
C173 VP.n23 B 0.02381f
C174 VP.n24 B 0.034611f
C175 VP.n25 B 0.044153f
C176 VP.t4 B 1.15071f
C177 VP.n26 B 0.426869f
C178 VP.n27 B 0.038268f
C179 VP.n28 B 0.02381f
C180 VP.n29 B 0.02381f
C181 VP.n30 B 0.02381f
C182 VP.n31 B 0.044153f
C183 VP.n32 B 0.046542f
C184 VP.n33 B 0.019352f
C185 VP.n34 B 0.02381f
C186 VP.n35 B 0.02381f
C187 VP.n36 B 0.02381f
C188 VP.n37 B 0.044153f
C189 VP.n38 B 0.026497f
C190 VP.n39 B 0.50864f
C191 VP.n40 B 1.25212f
C192 VP.n41 B 1.27001f
C193 VP.t5 B 1.15071f
C194 VP.n42 B 0.50864f
C195 VP.n43 B 0.026497f
C196 VP.n44 B 0.031389f
C197 VP.n45 B 0.02381f
C198 VP.n46 B 0.02381f
C199 VP.n47 B 0.047481f
C200 VP.n48 B 0.019352f
C201 VP.n49 B 0.046542f
C202 VP.n50 B 0.02381f
C203 VP.n51 B 0.02381f
C204 VP.n52 B 0.02381f
C205 VP.n53 B 0.028241f
C206 VP.n54 B 0.426869f
C207 VP.n55 B 0.038268f
C208 VP.n56 B 0.044153f
C209 VP.n57 B 0.02381f
C210 VP.n58 B 0.02381f
C211 VP.n59 B 0.02381f
C212 VP.n60 B 0.034611f
C213 VP.n61 B 0.044153f
C214 VP.t6 B 1.15071f
C215 VP.n62 B 0.426869f
C216 VP.n63 B 0.038268f
C217 VP.n64 B 0.02381f
C218 VP.n65 B 0.02381f
C219 VP.n66 B 0.02381f
C220 VP.n67 B 0.044153f
C221 VP.n68 B 0.046542f
C222 VP.n69 B 0.019352f
C223 VP.n70 B 0.02381f
C224 VP.n71 B 0.02381f
C225 VP.n72 B 0.02381f
C226 VP.n73 B 0.044153f
C227 VP.n74 B 0.026497f
C228 VP.n75 B 0.50864f
C229 VP.n76 B 0.044358f
.ends

