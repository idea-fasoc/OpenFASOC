* NGSPICE file created from diff_pair_sample_0087.ext - technology: sky130A

.subckt diff_pair_sample_0087 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n1554_n2238# sky130_fd_pr__pfet_01v8 ad=2.4765 pd=13.48 as=0 ps=0 w=6.35 l=0.4
X1 VTAIL.t11 VP.t0 VDD1.t0 w_n1554_n2238# sky130_fd_pr__pfet_01v8 ad=1.04775 pd=6.68 as=1.04775 ps=6.68 w=6.35 l=0.4
X2 VDD2.t5 VN.t0 VTAIL.t1 w_n1554_n2238# sky130_fd_pr__pfet_01v8 ad=2.4765 pd=13.48 as=1.04775 ps=6.68 w=6.35 l=0.4
X3 VTAIL.t0 VN.t1 VDD2.t4 w_n1554_n2238# sky130_fd_pr__pfet_01v8 ad=1.04775 pd=6.68 as=1.04775 ps=6.68 w=6.35 l=0.4
X4 VDD1.t2 VP.t1 VTAIL.t10 w_n1554_n2238# sky130_fd_pr__pfet_01v8 ad=1.04775 pd=6.68 as=2.4765 ps=13.48 w=6.35 l=0.4
X5 VTAIL.t9 VP.t2 VDD1.t1 w_n1554_n2238# sky130_fd_pr__pfet_01v8 ad=1.04775 pd=6.68 as=1.04775 ps=6.68 w=6.35 l=0.4
X6 VDD1.t5 VP.t3 VTAIL.t8 w_n1554_n2238# sky130_fd_pr__pfet_01v8 ad=2.4765 pd=13.48 as=1.04775 ps=6.68 w=6.35 l=0.4
X7 B.t8 B.t6 B.t7 w_n1554_n2238# sky130_fd_pr__pfet_01v8 ad=2.4765 pd=13.48 as=0 ps=0 w=6.35 l=0.4
X8 VDD2.t3 VN.t2 VTAIL.t5 w_n1554_n2238# sky130_fd_pr__pfet_01v8 ad=1.04775 pd=6.68 as=2.4765 ps=13.48 w=6.35 l=0.4
X9 B.t5 B.t3 B.t4 w_n1554_n2238# sky130_fd_pr__pfet_01v8 ad=2.4765 pd=13.48 as=0 ps=0 w=6.35 l=0.4
X10 B.t2 B.t0 B.t1 w_n1554_n2238# sky130_fd_pr__pfet_01v8 ad=2.4765 pd=13.48 as=0 ps=0 w=6.35 l=0.4
X11 VDD1.t4 VP.t4 VTAIL.t7 w_n1554_n2238# sky130_fd_pr__pfet_01v8 ad=2.4765 pd=13.48 as=1.04775 ps=6.68 w=6.35 l=0.4
X12 VDD2.t2 VN.t3 VTAIL.t4 w_n1554_n2238# sky130_fd_pr__pfet_01v8 ad=2.4765 pd=13.48 as=1.04775 ps=6.68 w=6.35 l=0.4
X13 VTAIL.t3 VN.t4 VDD2.t1 w_n1554_n2238# sky130_fd_pr__pfet_01v8 ad=1.04775 pd=6.68 as=1.04775 ps=6.68 w=6.35 l=0.4
X14 VDD1.t3 VP.t5 VTAIL.t6 w_n1554_n2238# sky130_fd_pr__pfet_01v8 ad=1.04775 pd=6.68 as=2.4765 ps=13.48 w=6.35 l=0.4
X15 VDD2.t0 VN.t5 VTAIL.t2 w_n1554_n2238# sky130_fd_pr__pfet_01v8 ad=1.04775 pd=6.68 as=2.4765 ps=13.48 w=6.35 l=0.4
R0 B.n160 B.t0 592.009
R1 B.n75 B.t9 592.009
R2 B.n31 B.t6 592.009
R3 B.n24 B.t3 592.009
R4 B.n217 B.n62 585
R5 B.n216 B.n215 585
R6 B.n214 B.n63 585
R7 B.n213 B.n212 585
R8 B.n211 B.n64 585
R9 B.n210 B.n209 585
R10 B.n208 B.n65 585
R11 B.n207 B.n206 585
R12 B.n205 B.n66 585
R13 B.n204 B.n203 585
R14 B.n202 B.n67 585
R15 B.n201 B.n200 585
R16 B.n199 B.n68 585
R17 B.n198 B.n197 585
R18 B.n196 B.n69 585
R19 B.n195 B.n194 585
R20 B.n193 B.n70 585
R21 B.n192 B.n191 585
R22 B.n190 B.n71 585
R23 B.n189 B.n188 585
R24 B.n187 B.n72 585
R25 B.n186 B.n185 585
R26 B.n184 B.n73 585
R27 B.n183 B.n182 585
R28 B.n181 B.n74 585
R29 B.n179 B.n178 585
R30 B.n177 B.n77 585
R31 B.n176 B.n175 585
R32 B.n174 B.n78 585
R33 B.n173 B.n172 585
R34 B.n171 B.n79 585
R35 B.n170 B.n169 585
R36 B.n168 B.n80 585
R37 B.n167 B.n166 585
R38 B.n165 B.n81 585
R39 B.n164 B.n163 585
R40 B.n159 B.n82 585
R41 B.n158 B.n157 585
R42 B.n156 B.n83 585
R43 B.n155 B.n154 585
R44 B.n153 B.n84 585
R45 B.n152 B.n151 585
R46 B.n150 B.n85 585
R47 B.n149 B.n148 585
R48 B.n147 B.n86 585
R49 B.n146 B.n145 585
R50 B.n144 B.n87 585
R51 B.n143 B.n142 585
R52 B.n141 B.n88 585
R53 B.n140 B.n139 585
R54 B.n138 B.n89 585
R55 B.n137 B.n136 585
R56 B.n135 B.n90 585
R57 B.n134 B.n133 585
R58 B.n132 B.n91 585
R59 B.n131 B.n130 585
R60 B.n129 B.n92 585
R61 B.n128 B.n127 585
R62 B.n126 B.n93 585
R63 B.n125 B.n124 585
R64 B.n219 B.n218 585
R65 B.n220 B.n61 585
R66 B.n222 B.n221 585
R67 B.n223 B.n60 585
R68 B.n225 B.n224 585
R69 B.n226 B.n59 585
R70 B.n228 B.n227 585
R71 B.n229 B.n58 585
R72 B.n231 B.n230 585
R73 B.n232 B.n57 585
R74 B.n234 B.n233 585
R75 B.n235 B.n56 585
R76 B.n237 B.n236 585
R77 B.n238 B.n55 585
R78 B.n240 B.n239 585
R79 B.n241 B.n54 585
R80 B.n243 B.n242 585
R81 B.n244 B.n53 585
R82 B.n246 B.n245 585
R83 B.n247 B.n52 585
R84 B.n249 B.n248 585
R85 B.n250 B.n51 585
R86 B.n252 B.n251 585
R87 B.n253 B.n50 585
R88 B.n255 B.n254 585
R89 B.n256 B.n49 585
R90 B.n258 B.n257 585
R91 B.n259 B.n48 585
R92 B.n261 B.n260 585
R93 B.n262 B.n47 585
R94 B.n264 B.n263 585
R95 B.n265 B.n46 585
R96 B.n267 B.n266 585
R97 B.n268 B.n45 585
R98 B.n359 B.n10 585
R99 B.n358 B.n357 585
R100 B.n356 B.n11 585
R101 B.n355 B.n354 585
R102 B.n353 B.n12 585
R103 B.n352 B.n351 585
R104 B.n350 B.n13 585
R105 B.n349 B.n348 585
R106 B.n347 B.n14 585
R107 B.n346 B.n345 585
R108 B.n344 B.n15 585
R109 B.n343 B.n342 585
R110 B.n341 B.n16 585
R111 B.n340 B.n339 585
R112 B.n338 B.n17 585
R113 B.n337 B.n336 585
R114 B.n335 B.n18 585
R115 B.n334 B.n333 585
R116 B.n332 B.n19 585
R117 B.n331 B.n330 585
R118 B.n329 B.n20 585
R119 B.n328 B.n327 585
R120 B.n326 B.n21 585
R121 B.n325 B.n324 585
R122 B.n323 B.n22 585
R123 B.n322 B.n321 585
R124 B.n320 B.n23 585
R125 B.n319 B.n318 585
R126 B.n317 B.n27 585
R127 B.n316 B.n315 585
R128 B.n314 B.n28 585
R129 B.n313 B.n312 585
R130 B.n311 B.n29 585
R131 B.n310 B.n309 585
R132 B.n308 B.n30 585
R133 B.n306 B.n305 585
R134 B.n304 B.n33 585
R135 B.n303 B.n302 585
R136 B.n301 B.n34 585
R137 B.n300 B.n299 585
R138 B.n298 B.n35 585
R139 B.n297 B.n296 585
R140 B.n295 B.n36 585
R141 B.n294 B.n293 585
R142 B.n292 B.n37 585
R143 B.n291 B.n290 585
R144 B.n289 B.n38 585
R145 B.n288 B.n287 585
R146 B.n286 B.n39 585
R147 B.n285 B.n284 585
R148 B.n283 B.n40 585
R149 B.n282 B.n281 585
R150 B.n280 B.n41 585
R151 B.n279 B.n278 585
R152 B.n277 B.n42 585
R153 B.n276 B.n275 585
R154 B.n274 B.n43 585
R155 B.n273 B.n272 585
R156 B.n271 B.n44 585
R157 B.n270 B.n269 585
R158 B.n361 B.n360 585
R159 B.n362 B.n9 585
R160 B.n364 B.n363 585
R161 B.n365 B.n8 585
R162 B.n367 B.n366 585
R163 B.n368 B.n7 585
R164 B.n370 B.n369 585
R165 B.n371 B.n6 585
R166 B.n373 B.n372 585
R167 B.n374 B.n5 585
R168 B.n376 B.n375 585
R169 B.n377 B.n4 585
R170 B.n379 B.n378 585
R171 B.n380 B.n3 585
R172 B.n382 B.n381 585
R173 B.n383 B.n0 585
R174 B.n2 B.n1 585
R175 B.n102 B.n101 585
R176 B.n104 B.n103 585
R177 B.n105 B.n100 585
R178 B.n107 B.n106 585
R179 B.n108 B.n99 585
R180 B.n110 B.n109 585
R181 B.n111 B.n98 585
R182 B.n113 B.n112 585
R183 B.n114 B.n97 585
R184 B.n116 B.n115 585
R185 B.n117 B.n96 585
R186 B.n119 B.n118 585
R187 B.n120 B.n95 585
R188 B.n122 B.n121 585
R189 B.n123 B.n94 585
R190 B.n125 B.n94 497.305
R191 B.n219 B.n62 497.305
R192 B.n269 B.n268 497.305
R193 B.n360 B.n359 497.305
R194 B.n385 B.n384 256.663
R195 B.n384 B.n383 235.042
R196 B.n384 B.n2 235.042
R197 B.n126 B.n125 163.367
R198 B.n127 B.n126 163.367
R199 B.n127 B.n92 163.367
R200 B.n131 B.n92 163.367
R201 B.n132 B.n131 163.367
R202 B.n133 B.n132 163.367
R203 B.n133 B.n90 163.367
R204 B.n137 B.n90 163.367
R205 B.n138 B.n137 163.367
R206 B.n139 B.n138 163.367
R207 B.n139 B.n88 163.367
R208 B.n143 B.n88 163.367
R209 B.n144 B.n143 163.367
R210 B.n145 B.n144 163.367
R211 B.n145 B.n86 163.367
R212 B.n149 B.n86 163.367
R213 B.n150 B.n149 163.367
R214 B.n151 B.n150 163.367
R215 B.n151 B.n84 163.367
R216 B.n155 B.n84 163.367
R217 B.n156 B.n155 163.367
R218 B.n157 B.n156 163.367
R219 B.n157 B.n82 163.367
R220 B.n164 B.n82 163.367
R221 B.n165 B.n164 163.367
R222 B.n166 B.n165 163.367
R223 B.n166 B.n80 163.367
R224 B.n170 B.n80 163.367
R225 B.n171 B.n170 163.367
R226 B.n172 B.n171 163.367
R227 B.n172 B.n78 163.367
R228 B.n176 B.n78 163.367
R229 B.n177 B.n176 163.367
R230 B.n178 B.n177 163.367
R231 B.n178 B.n74 163.367
R232 B.n183 B.n74 163.367
R233 B.n184 B.n183 163.367
R234 B.n185 B.n184 163.367
R235 B.n185 B.n72 163.367
R236 B.n189 B.n72 163.367
R237 B.n190 B.n189 163.367
R238 B.n191 B.n190 163.367
R239 B.n191 B.n70 163.367
R240 B.n195 B.n70 163.367
R241 B.n196 B.n195 163.367
R242 B.n197 B.n196 163.367
R243 B.n197 B.n68 163.367
R244 B.n201 B.n68 163.367
R245 B.n202 B.n201 163.367
R246 B.n203 B.n202 163.367
R247 B.n203 B.n66 163.367
R248 B.n207 B.n66 163.367
R249 B.n208 B.n207 163.367
R250 B.n209 B.n208 163.367
R251 B.n209 B.n64 163.367
R252 B.n213 B.n64 163.367
R253 B.n214 B.n213 163.367
R254 B.n215 B.n214 163.367
R255 B.n215 B.n62 163.367
R256 B.n268 B.n267 163.367
R257 B.n267 B.n46 163.367
R258 B.n263 B.n46 163.367
R259 B.n263 B.n262 163.367
R260 B.n262 B.n261 163.367
R261 B.n261 B.n48 163.367
R262 B.n257 B.n48 163.367
R263 B.n257 B.n256 163.367
R264 B.n256 B.n255 163.367
R265 B.n255 B.n50 163.367
R266 B.n251 B.n50 163.367
R267 B.n251 B.n250 163.367
R268 B.n250 B.n249 163.367
R269 B.n249 B.n52 163.367
R270 B.n245 B.n52 163.367
R271 B.n245 B.n244 163.367
R272 B.n244 B.n243 163.367
R273 B.n243 B.n54 163.367
R274 B.n239 B.n54 163.367
R275 B.n239 B.n238 163.367
R276 B.n238 B.n237 163.367
R277 B.n237 B.n56 163.367
R278 B.n233 B.n56 163.367
R279 B.n233 B.n232 163.367
R280 B.n232 B.n231 163.367
R281 B.n231 B.n58 163.367
R282 B.n227 B.n58 163.367
R283 B.n227 B.n226 163.367
R284 B.n226 B.n225 163.367
R285 B.n225 B.n60 163.367
R286 B.n221 B.n60 163.367
R287 B.n221 B.n220 163.367
R288 B.n220 B.n219 163.367
R289 B.n359 B.n358 163.367
R290 B.n358 B.n11 163.367
R291 B.n354 B.n11 163.367
R292 B.n354 B.n353 163.367
R293 B.n353 B.n352 163.367
R294 B.n352 B.n13 163.367
R295 B.n348 B.n13 163.367
R296 B.n348 B.n347 163.367
R297 B.n347 B.n346 163.367
R298 B.n346 B.n15 163.367
R299 B.n342 B.n15 163.367
R300 B.n342 B.n341 163.367
R301 B.n341 B.n340 163.367
R302 B.n340 B.n17 163.367
R303 B.n336 B.n17 163.367
R304 B.n336 B.n335 163.367
R305 B.n335 B.n334 163.367
R306 B.n334 B.n19 163.367
R307 B.n330 B.n19 163.367
R308 B.n330 B.n329 163.367
R309 B.n329 B.n328 163.367
R310 B.n328 B.n21 163.367
R311 B.n324 B.n21 163.367
R312 B.n324 B.n323 163.367
R313 B.n323 B.n322 163.367
R314 B.n322 B.n23 163.367
R315 B.n318 B.n23 163.367
R316 B.n318 B.n317 163.367
R317 B.n317 B.n316 163.367
R318 B.n316 B.n28 163.367
R319 B.n312 B.n28 163.367
R320 B.n312 B.n311 163.367
R321 B.n311 B.n310 163.367
R322 B.n310 B.n30 163.367
R323 B.n305 B.n30 163.367
R324 B.n305 B.n304 163.367
R325 B.n304 B.n303 163.367
R326 B.n303 B.n34 163.367
R327 B.n299 B.n34 163.367
R328 B.n299 B.n298 163.367
R329 B.n298 B.n297 163.367
R330 B.n297 B.n36 163.367
R331 B.n293 B.n36 163.367
R332 B.n293 B.n292 163.367
R333 B.n292 B.n291 163.367
R334 B.n291 B.n38 163.367
R335 B.n287 B.n38 163.367
R336 B.n287 B.n286 163.367
R337 B.n286 B.n285 163.367
R338 B.n285 B.n40 163.367
R339 B.n281 B.n40 163.367
R340 B.n281 B.n280 163.367
R341 B.n280 B.n279 163.367
R342 B.n279 B.n42 163.367
R343 B.n275 B.n42 163.367
R344 B.n275 B.n274 163.367
R345 B.n274 B.n273 163.367
R346 B.n273 B.n44 163.367
R347 B.n269 B.n44 163.367
R348 B.n360 B.n9 163.367
R349 B.n364 B.n9 163.367
R350 B.n365 B.n364 163.367
R351 B.n366 B.n365 163.367
R352 B.n366 B.n7 163.367
R353 B.n370 B.n7 163.367
R354 B.n371 B.n370 163.367
R355 B.n372 B.n371 163.367
R356 B.n372 B.n5 163.367
R357 B.n376 B.n5 163.367
R358 B.n377 B.n376 163.367
R359 B.n378 B.n377 163.367
R360 B.n378 B.n3 163.367
R361 B.n382 B.n3 163.367
R362 B.n383 B.n382 163.367
R363 B.n102 B.n2 163.367
R364 B.n103 B.n102 163.367
R365 B.n103 B.n100 163.367
R366 B.n107 B.n100 163.367
R367 B.n108 B.n107 163.367
R368 B.n109 B.n108 163.367
R369 B.n109 B.n98 163.367
R370 B.n113 B.n98 163.367
R371 B.n114 B.n113 163.367
R372 B.n115 B.n114 163.367
R373 B.n115 B.n96 163.367
R374 B.n119 B.n96 163.367
R375 B.n120 B.n119 163.367
R376 B.n121 B.n120 163.367
R377 B.n121 B.n94 163.367
R378 B.n75 B.t10 129.198
R379 B.n31 B.t8 129.198
R380 B.n160 B.t1 129.192
R381 B.n24 B.t5 129.192
R382 B.n76 B.t11 115.041
R383 B.n32 B.t7 115.041
R384 B.n161 B.t2 115.034
R385 B.n25 B.t4 115.034
R386 B.n162 B.n161 59.5399
R387 B.n180 B.n76 59.5399
R388 B.n307 B.n32 59.5399
R389 B.n26 B.n25 59.5399
R390 B.n361 B.n10 32.3127
R391 B.n270 B.n45 32.3127
R392 B.n218 B.n217 32.3127
R393 B.n124 B.n123 32.3127
R394 B B.n385 18.0485
R395 B.n161 B.n160 14.1581
R396 B.n76 B.n75 14.1581
R397 B.n32 B.n31 14.1581
R398 B.n25 B.n24 14.1581
R399 B.n362 B.n361 10.6151
R400 B.n363 B.n362 10.6151
R401 B.n363 B.n8 10.6151
R402 B.n367 B.n8 10.6151
R403 B.n368 B.n367 10.6151
R404 B.n369 B.n368 10.6151
R405 B.n369 B.n6 10.6151
R406 B.n373 B.n6 10.6151
R407 B.n374 B.n373 10.6151
R408 B.n375 B.n374 10.6151
R409 B.n375 B.n4 10.6151
R410 B.n379 B.n4 10.6151
R411 B.n380 B.n379 10.6151
R412 B.n381 B.n380 10.6151
R413 B.n381 B.n0 10.6151
R414 B.n357 B.n10 10.6151
R415 B.n357 B.n356 10.6151
R416 B.n356 B.n355 10.6151
R417 B.n355 B.n12 10.6151
R418 B.n351 B.n12 10.6151
R419 B.n351 B.n350 10.6151
R420 B.n350 B.n349 10.6151
R421 B.n349 B.n14 10.6151
R422 B.n345 B.n14 10.6151
R423 B.n345 B.n344 10.6151
R424 B.n344 B.n343 10.6151
R425 B.n343 B.n16 10.6151
R426 B.n339 B.n16 10.6151
R427 B.n339 B.n338 10.6151
R428 B.n338 B.n337 10.6151
R429 B.n337 B.n18 10.6151
R430 B.n333 B.n18 10.6151
R431 B.n333 B.n332 10.6151
R432 B.n332 B.n331 10.6151
R433 B.n331 B.n20 10.6151
R434 B.n327 B.n20 10.6151
R435 B.n327 B.n326 10.6151
R436 B.n326 B.n325 10.6151
R437 B.n325 B.n22 10.6151
R438 B.n321 B.n320 10.6151
R439 B.n320 B.n319 10.6151
R440 B.n319 B.n27 10.6151
R441 B.n315 B.n27 10.6151
R442 B.n315 B.n314 10.6151
R443 B.n314 B.n313 10.6151
R444 B.n313 B.n29 10.6151
R445 B.n309 B.n29 10.6151
R446 B.n309 B.n308 10.6151
R447 B.n306 B.n33 10.6151
R448 B.n302 B.n33 10.6151
R449 B.n302 B.n301 10.6151
R450 B.n301 B.n300 10.6151
R451 B.n300 B.n35 10.6151
R452 B.n296 B.n35 10.6151
R453 B.n296 B.n295 10.6151
R454 B.n295 B.n294 10.6151
R455 B.n294 B.n37 10.6151
R456 B.n290 B.n37 10.6151
R457 B.n290 B.n289 10.6151
R458 B.n289 B.n288 10.6151
R459 B.n288 B.n39 10.6151
R460 B.n284 B.n39 10.6151
R461 B.n284 B.n283 10.6151
R462 B.n283 B.n282 10.6151
R463 B.n282 B.n41 10.6151
R464 B.n278 B.n41 10.6151
R465 B.n278 B.n277 10.6151
R466 B.n277 B.n276 10.6151
R467 B.n276 B.n43 10.6151
R468 B.n272 B.n43 10.6151
R469 B.n272 B.n271 10.6151
R470 B.n271 B.n270 10.6151
R471 B.n266 B.n45 10.6151
R472 B.n266 B.n265 10.6151
R473 B.n265 B.n264 10.6151
R474 B.n264 B.n47 10.6151
R475 B.n260 B.n47 10.6151
R476 B.n260 B.n259 10.6151
R477 B.n259 B.n258 10.6151
R478 B.n258 B.n49 10.6151
R479 B.n254 B.n49 10.6151
R480 B.n254 B.n253 10.6151
R481 B.n253 B.n252 10.6151
R482 B.n252 B.n51 10.6151
R483 B.n248 B.n51 10.6151
R484 B.n248 B.n247 10.6151
R485 B.n247 B.n246 10.6151
R486 B.n246 B.n53 10.6151
R487 B.n242 B.n53 10.6151
R488 B.n242 B.n241 10.6151
R489 B.n241 B.n240 10.6151
R490 B.n240 B.n55 10.6151
R491 B.n236 B.n55 10.6151
R492 B.n236 B.n235 10.6151
R493 B.n235 B.n234 10.6151
R494 B.n234 B.n57 10.6151
R495 B.n230 B.n57 10.6151
R496 B.n230 B.n229 10.6151
R497 B.n229 B.n228 10.6151
R498 B.n228 B.n59 10.6151
R499 B.n224 B.n59 10.6151
R500 B.n224 B.n223 10.6151
R501 B.n223 B.n222 10.6151
R502 B.n222 B.n61 10.6151
R503 B.n218 B.n61 10.6151
R504 B.n101 B.n1 10.6151
R505 B.n104 B.n101 10.6151
R506 B.n105 B.n104 10.6151
R507 B.n106 B.n105 10.6151
R508 B.n106 B.n99 10.6151
R509 B.n110 B.n99 10.6151
R510 B.n111 B.n110 10.6151
R511 B.n112 B.n111 10.6151
R512 B.n112 B.n97 10.6151
R513 B.n116 B.n97 10.6151
R514 B.n117 B.n116 10.6151
R515 B.n118 B.n117 10.6151
R516 B.n118 B.n95 10.6151
R517 B.n122 B.n95 10.6151
R518 B.n123 B.n122 10.6151
R519 B.n124 B.n93 10.6151
R520 B.n128 B.n93 10.6151
R521 B.n129 B.n128 10.6151
R522 B.n130 B.n129 10.6151
R523 B.n130 B.n91 10.6151
R524 B.n134 B.n91 10.6151
R525 B.n135 B.n134 10.6151
R526 B.n136 B.n135 10.6151
R527 B.n136 B.n89 10.6151
R528 B.n140 B.n89 10.6151
R529 B.n141 B.n140 10.6151
R530 B.n142 B.n141 10.6151
R531 B.n142 B.n87 10.6151
R532 B.n146 B.n87 10.6151
R533 B.n147 B.n146 10.6151
R534 B.n148 B.n147 10.6151
R535 B.n148 B.n85 10.6151
R536 B.n152 B.n85 10.6151
R537 B.n153 B.n152 10.6151
R538 B.n154 B.n153 10.6151
R539 B.n154 B.n83 10.6151
R540 B.n158 B.n83 10.6151
R541 B.n159 B.n158 10.6151
R542 B.n163 B.n159 10.6151
R543 B.n167 B.n81 10.6151
R544 B.n168 B.n167 10.6151
R545 B.n169 B.n168 10.6151
R546 B.n169 B.n79 10.6151
R547 B.n173 B.n79 10.6151
R548 B.n174 B.n173 10.6151
R549 B.n175 B.n174 10.6151
R550 B.n175 B.n77 10.6151
R551 B.n179 B.n77 10.6151
R552 B.n182 B.n181 10.6151
R553 B.n182 B.n73 10.6151
R554 B.n186 B.n73 10.6151
R555 B.n187 B.n186 10.6151
R556 B.n188 B.n187 10.6151
R557 B.n188 B.n71 10.6151
R558 B.n192 B.n71 10.6151
R559 B.n193 B.n192 10.6151
R560 B.n194 B.n193 10.6151
R561 B.n194 B.n69 10.6151
R562 B.n198 B.n69 10.6151
R563 B.n199 B.n198 10.6151
R564 B.n200 B.n199 10.6151
R565 B.n200 B.n67 10.6151
R566 B.n204 B.n67 10.6151
R567 B.n205 B.n204 10.6151
R568 B.n206 B.n205 10.6151
R569 B.n206 B.n65 10.6151
R570 B.n210 B.n65 10.6151
R571 B.n211 B.n210 10.6151
R572 B.n212 B.n211 10.6151
R573 B.n212 B.n63 10.6151
R574 B.n216 B.n63 10.6151
R575 B.n217 B.n216 10.6151
R576 B.n26 B.n22 9.36635
R577 B.n307 B.n306 9.36635
R578 B.n163 B.n162 9.36635
R579 B.n181 B.n180 9.36635
R580 B.n385 B.n0 8.11757
R581 B.n385 B.n1 8.11757
R582 B.n321 B.n26 1.24928
R583 B.n308 B.n307 1.24928
R584 B.n162 B.n81 1.24928
R585 B.n180 B.n179 1.24928
R586 VP.n1 VP.t4 505.082
R587 VP.n8 VP.t5 485.779
R588 VP.n6 VP.t3 485.779
R589 VP.n3 VP.t1 485.779
R590 VP.n7 VP.t0 481.397
R591 VP.n2 VP.t2 481.397
R592 VP.n9 VP.n8 161.3
R593 VP.n4 VP.n3 161.3
R594 VP.n7 VP.n0 161.3
R595 VP.n6 VP.n5 161.3
R596 VP.n4 VP.n1 71.2425
R597 VP.n7 VP.n6 43.8187
R598 VP.n8 VP.n7 43.8187
R599 VP.n3 VP.n2 43.8187
R600 VP.n5 VP.n4 35.8225
R601 VP.n2 VP.n1 19.2801
R602 VP.n5 VP.n0 0.189894
R603 VP.n9 VP.n0 0.189894
R604 VP VP.n9 0.0516364
R605 VDD1 VDD1.t4 95.6835
R606 VDD1.n1 VDD1.t5 95.5699
R607 VDD1.n1 VDD1.n0 90.1363
R608 VDD1.n3 VDD1.n2 90.0343
R609 VDD1.n3 VDD1.n1 32.1324
R610 VDD1.n2 VDD1.t1 5.1194
R611 VDD1.n2 VDD1.t2 5.1194
R612 VDD1.n0 VDD1.t0 5.1194
R613 VDD1.n0 VDD1.t3 5.1194
R614 VDD1 VDD1.n3 0.0996379
R615 VTAIL.n7 VTAIL.t5 78.4746
R616 VTAIL.n11 VTAIL.t2 78.4745
R617 VTAIL.n2 VTAIL.t6 78.4745
R618 VTAIL.n10 VTAIL.t10 78.4744
R619 VTAIL.n9 VTAIL.n8 73.3557
R620 VTAIL.n6 VTAIL.n5 73.3557
R621 VTAIL.n1 VTAIL.n0 73.3555
R622 VTAIL.n4 VTAIL.n3 73.3555
R623 VTAIL.n6 VTAIL.n4 19.0996
R624 VTAIL.n11 VTAIL.n10 18.4703
R625 VTAIL.n0 VTAIL.t4 5.1194
R626 VTAIL.n0 VTAIL.t3 5.1194
R627 VTAIL.n3 VTAIL.t8 5.1194
R628 VTAIL.n3 VTAIL.t11 5.1194
R629 VTAIL.n8 VTAIL.t7 5.1194
R630 VTAIL.n8 VTAIL.t9 5.1194
R631 VTAIL.n5 VTAIL.t1 5.1194
R632 VTAIL.n5 VTAIL.t0 5.1194
R633 VTAIL.n9 VTAIL.n7 0.784983
R634 VTAIL.n2 VTAIL.n1 0.784983
R635 VTAIL.n7 VTAIL.n6 0.62981
R636 VTAIL.n10 VTAIL.n9 0.62981
R637 VTAIL.n4 VTAIL.n2 0.62981
R638 VTAIL VTAIL.n11 0.414293
R639 VTAIL VTAIL.n1 0.216017
R640 VN.n0 VN.t3 505.082
R641 VN.n4 VN.t2 505.082
R642 VN.n2 VN.t5 485.779
R643 VN.n6 VN.t0 485.779
R644 VN.n1 VN.t4 481.397
R645 VN.n5 VN.t1 481.397
R646 VN.n3 VN.n2 161.3
R647 VN.n7 VN.n6 161.3
R648 VN.n7 VN.n4 71.2425
R649 VN.n3 VN.n0 71.2425
R650 VN.n2 VN.n1 43.8187
R651 VN.n6 VN.n5 43.8187
R652 VN VN.n7 36.2031
R653 VN.n5 VN.n4 19.2801
R654 VN.n1 VN.n0 19.2801
R655 VN VN.n3 0.0516364
R656 VDD2.n1 VDD2.t2 95.5699
R657 VDD2.n2 VDD2.t5 95.1534
R658 VDD2.n1 VDD2.n0 90.1363
R659 VDD2 VDD2.n3 90.1335
R660 VDD2.n2 VDD2.n1 31.2347
R661 VDD2.n3 VDD2.t4 5.1194
R662 VDD2.n3 VDD2.t3 5.1194
R663 VDD2.n0 VDD2.t1 5.1194
R664 VDD2.n0 VDD2.t0 5.1194
R665 VDD2 VDD2.n2 0.530672
C0 VDD2 VN 1.84634f
C1 VDD1 VTAIL 7.34455f
C2 VP B 0.945668f
C3 VDD1 B 1.06418f
C4 VTAIL w_n1554_n2238# 2.03832f
C5 VDD1 VP 1.96725f
C6 VTAIL VN 1.70497f
C7 w_n1554_n2238# B 5.058661f
C8 VDD2 VTAIL 7.37904f
C9 VN B 0.631539f
C10 VDD2 B 1.08643f
C11 VP w_n1554_n2238# 2.49716f
C12 VN VP 3.74236f
C13 VDD1 w_n1554_n2238# 1.30168f
C14 VDD2 VP 0.271377f
C15 VDD1 VN 0.147724f
C16 VDD2 VDD1 0.602802f
C17 VTAIL B 1.55338f
C18 VN w_n1554_n2238# 2.30238f
C19 VTAIL VP 1.7194f
C20 VDD2 w_n1554_n2238# 1.31662f
C21 VDD2 VSUBS 0.955522f
C22 VDD1 VSUBS 1.173635f
C23 VTAIL VSUBS 0.38336f
C24 VN VSUBS 2.99642f
C25 VP VSUBS 0.972546f
C26 B VSUBS 1.968528f
C27 w_n1554_n2238# VSUBS 43.3566f
C28 VDD2.t2 VSUBS 0.934842f
C29 VDD2.t1 VSUBS 0.103691f
C30 VDD2.t0 VSUBS 0.103691f
C31 VDD2.n0 VSUBS 0.697797f
C32 VDD2.n1 VSUBS 1.67391f
C33 VDD2.t5 VSUBS 0.932988f
C34 VDD2.n2 VSUBS 1.60776f
C35 VDD2.t4 VSUBS 0.103691f
C36 VDD2.t3 VSUBS 0.103691f
C37 VDD2.n3 VSUBS 0.697779f
C38 VN.t3 VSUBS 0.335512f
C39 VN.n0 VSUBS 0.148322f
C40 VN.t4 VSUBS 0.328321f
C41 VN.n1 VSUBS 0.161789f
C42 VN.t5 VSUBS 0.329629f
C43 VN.n2 VSUBS 0.153878f
C44 VN.n3 VSUBS 0.133409f
C45 VN.t2 VSUBS 0.335512f
C46 VN.n4 VSUBS 0.148322f
C47 VN.t0 VSUBS 0.329629f
C48 VN.t1 VSUBS 0.328321f
C49 VN.n5 VSUBS 0.161789f
C50 VN.n6 VSUBS 0.153878f
C51 VN.n7 VSUBS 1.5184f
C52 VTAIL.t4 VSUBS 0.128976f
C53 VTAIL.t3 VSUBS 0.128976f
C54 VTAIL.n0 VSUBS 0.771815f
C55 VTAIL.n1 VSUBS 0.568701f
C56 VTAIL.t6 VSUBS 1.05869f
C57 VTAIL.n2 VSUBS 0.66785f
C58 VTAIL.t8 VSUBS 0.128976f
C59 VTAIL.t11 VSUBS 0.128976f
C60 VTAIL.n3 VSUBS 0.771815f
C61 VTAIL.n4 VSUBS 1.44475f
C62 VTAIL.t1 VSUBS 0.128976f
C63 VTAIL.t0 VSUBS 0.128976f
C64 VTAIL.n5 VSUBS 0.771819f
C65 VTAIL.n6 VSUBS 1.44475f
C66 VTAIL.t5 VSUBS 1.0587f
C67 VTAIL.n7 VSUBS 0.667844f
C68 VTAIL.t7 VSUBS 0.128976f
C69 VTAIL.t9 VSUBS 0.128976f
C70 VTAIL.n8 VSUBS 0.771819f
C71 VTAIL.n9 VSUBS 0.602966f
C72 VTAIL.t10 VSUBS 1.05869f
C73 VTAIL.n10 VSUBS 1.45751f
C74 VTAIL.t2 VSUBS 1.05869f
C75 VTAIL.n11 VSUBS 1.43966f
C76 VDD1.t4 VSUBS 0.913325f
C77 VDD1.t5 VSUBS 0.912795f
C78 VDD1.t0 VSUBS 0.101245f
C79 VDD1.t3 VSUBS 0.101245f
C80 VDD1.n0 VSUBS 0.68134f
C81 VDD1.n1 VSUBS 1.68976f
C82 VDD1.t1 VSUBS 0.101245f
C83 VDD1.t2 VSUBS 0.101245f
C84 VDD1.n2 VSUBS 0.680894f
C85 VDD1.n3 VSUBS 1.55589f
C86 VP.n0 VSUBS 0.046599f
C87 VP.t3 VSUBS 0.344216f
C88 VP.t4 VSUBS 0.350359f
C89 VP.n1 VSUBS 0.154885f
C90 VP.t2 VSUBS 0.342849f
C91 VP.n2 VSUBS 0.168948f
C92 VP.t1 VSUBS 0.344216f
C93 VP.n3 VSUBS 0.160687f
C94 VP.n4 VSUBS 1.55468f
C95 VP.n5 VSUBS 1.49824f
C96 VP.n6 VSUBS 0.160687f
C97 VP.t0 VSUBS 0.342849f
C98 VP.n7 VSUBS 0.168948f
C99 VP.t5 VSUBS 0.344216f
C100 VP.n8 VSUBS 0.160687f
C101 VP.n9 VSUBS 0.036113f
C102 B.n0 VSUBS 0.005882f
C103 B.n1 VSUBS 0.005882f
C104 B.n2 VSUBS 0.008698f
C105 B.n3 VSUBS 0.006666f
C106 B.n4 VSUBS 0.006666f
C107 B.n5 VSUBS 0.006666f
C108 B.n6 VSUBS 0.006666f
C109 B.n7 VSUBS 0.006666f
C110 B.n8 VSUBS 0.006666f
C111 B.n9 VSUBS 0.006666f
C112 B.n10 VSUBS 0.016139f
C113 B.n11 VSUBS 0.006666f
C114 B.n12 VSUBS 0.006666f
C115 B.n13 VSUBS 0.006666f
C116 B.n14 VSUBS 0.006666f
C117 B.n15 VSUBS 0.006666f
C118 B.n16 VSUBS 0.006666f
C119 B.n17 VSUBS 0.006666f
C120 B.n18 VSUBS 0.006666f
C121 B.n19 VSUBS 0.006666f
C122 B.n20 VSUBS 0.006666f
C123 B.n21 VSUBS 0.006666f
C124 B.n22 VSUBS 0.006274f
C125 B.n23 VSUBS 0.006666f
C126 B.t4 VSUBS 0.17857f
C127 B.t5 VSUBS 0.183993f
C128 B.t3 VSUBS 0.100011f
C129 B.n24 VSUBS 0.076468f
C130 B.n25 VSUBS 0.058987f
C131 B.n26 VSUBS 0.015444f
C132 B.n27 VSUBS 0.006666f
C133 B.n28 VSUBS 0.006666f
C134 B.n29 VSUBS 0.006666f
C135 B.n30 VSUBS 0.006666f
C136 B.t7 VSUBS 0.17857f
C137 B.t8 VSUBS 0.183992f
C138 B.t6 VSUBS 0.100011f
C139 B.n31 VSUBS 0.076469f
C140 B.n32 VSUBS 0.058988f
C141 B.n33 VSUBS 0.006666f
C142 B.n34 VSUBS 0.006666f
C143 B.n35 VSUBS 0.006666f
C144 B.n36 VSUBS 0.006666f
C145 B.n37 VSUBS 0.006666f
C146 B.n38 VSUBS 0.006666f
C147 B.n39 VSUBS 0.006666f
C148 B.n40 VSUBS 0.006666f
C149 B.n41 VSUBS 0.006666f
C150 B.n42 VSUBS 0.006666f
C151 B.n43 VSUBS 0.006666f
C152 B.n44 VSUBS 0.006666f
C153 B.n45 VSUBS 0.014838f
C154 B.n46 VSUBS 0.006666f
C155 B.n47 VSUBS 0.006666f
C156 B.n48 VSUBS 0.006666f
C157 B.n49 VSUBS 0.006666f
C158 B.n50 VSUBS 0.006666f
C159 B.n51 VSUBS 0.006666f
C160 B.n52 VSUBS 0.006666f
C161 B.n53 VSUBS 0.006666f
C162 B.n54 VSUBS 0.006666f
C163 B.n55 VSUBS 0.006666f
C164 B.n56 VSUBS 0.006666f
C165 B.n57 VSUBS 0.006666f
C166 B.n58 VSUBS 0.006666f
C167 B.n59 VSUBS 0.006666f
C168 B.n60 VSUBS 0.006666f
C169 B.n61 VSUBS 0.006666f
C170 B.n62 VSUBS 0.016139f
C171 B.n63 VSUBS 0.006666f
C172 B.n64 VSUBS 0.006666f
C173 B.n65 VSUBS 0.006666f
C174 B.n66 VSUBS 0.006666f
C175 B.n67 VSUBS 0.006666f
C176 B.n68 VSUBS 0.006666f
C177 B.n69 VSUBS 0.006666f
C178 B.n70 VSUBS 0.006666f
C179 B.n71 VSUBS 0.006666f
C180 B.n72 VSUBS 0.006666f
C181 B.n73 VSUBS 0.006666f
C182 B.n74 VSUBS 0.006666f
C183 B.t11 VSUBS 0.17857f
C184 B.t10 VSUBS 0.183992f
C185 B.t9 VSUBS 0.100011f
C186 B.n75 VSUBS 0.076469f
C187 B.n76 VSUBS 0.058988f
C188 B.n77 VSUBS 0.006666f
C189 B.n78 VSUBS 0.006666f
C190 B.n79 VSUBS 0.006666f
C191 B.n80 VSUBS 0.006666f
C192 B.n81 VSUBS 0.003725f
C193 B.n82 VSUBS 0.006666f
C194 B.n83 VSUBS 0.006666f
C195 B.n84 VSUBS 0.006666f
C196 B.n85 VSUBS 0.006666f
C197 B.n86 VSUBS 0.006666f
C198 B.n87 VSUBS 0.006666f
C199 B.n88 VSUBS 0.006666f
C200 B.n89 VSUBS 0.006666f
C201 B.n90 VSUBS 0.006666f
C202 B.n91 VSUBS 0.006666f
C203 B.n92 VSUBS 0.006666f
C204 B.n93 VSUBS 0.006666f
C205 B.n94 VSUBS 0.014838f
C206 B.n95 VSUBS 0.006666f
C207 B.n96 VSUBS 0.006666f
C208 B.n97 VSUBS 0.006666f
C209 B.n98 VSUBS 0.006666f
C210 B.n99 VSUBS 0.006666f
C211 B.n100 VSUBS 0.006666f
C212 B.n101 VSUBS 0.006666f
C213 B.n102 VSUBS 0.006666f
C214 B.n103 VSUBS 0.006666f
C215 B.n104 VSUBS 0.006666f
C216 B.n105 VSUBS 0.006666f
C217 B.n106 VSUBS 0.006666f
C218 B.n107 VSUBS 0.006666f
C219 B.n108 VSUBS 0.006666f
C220 B.n109 VSUBS 0.006666f
C221 B.n110 VSUBS 0.006666f
C222 B.n111 VSUBS 0.006666f
C223 B.n112 VSUBS 0.006666f
C224 B.n113 VSUBS 0.006666f
C225 B.n114 VSUBS 0.006666f
C226 B.n115 VSUBS 0.006666f
C227 B.n116 VSUBS 0.006666f
C228 B.n117 VSUBS 0.006666f
C229 B.n118 VSUBS 0.006666f
C230 B.n119 VSUBS 0.006666f
C231 B.n120 VSUBS 0.006666f
C232 B.n121 VSUBS 0.006666f
C233 B.n122 VSUBS 0.006666f
C234 B.n123 VSUBS 0.014838f
C235 B.n124 VSUBS 0.016139f
C236 B.n125 VSUBS 0.016139f
C237 B.n126 VSUBS 0.006666f
C238 B.n127 VSUBS 0.006666f
C239 B.n128 VSUBS 0.006666f
C240 B.n129 VSUBS 0.006666f
C241 B.n130 VSUBS 0.006666f
C242 B.n131 VSUBS 0.006666f
C243 B.n132 VSUBS 0.006666f
C244 B.n133 VSUBS 0.006666f
C245 B.n134 VSUBS 0.006666f
C246 B.n135 VSUBS 0.006666f
C247 B.n136 VSUBS 0.006666f
C248 B.n137 VSUBS 0.006666f
C249 B.n138 VSUBS 0.006666f
C250 B.n139 VSUBS 0.006666f
C251 B.n140 VSUBS 0.006666f
C252 B.n141 VSUBS 0.006666f
C253 B.n142 VSUBS 0.006666f
C254 B.n143 VSUBS 0.006666f
C255 B.n144 VSUBS 0.006666f
C256 B.n145 VSUBS 0.006666f
C257 B.n146 VSUBS 0.006666f
C258 B.n147 VSUBS 0.006666f
C259 B.n148 VSUBS 0.006666f
C260 B.n149 VSUBS 0.006666f
C261 B.n150 VSUBS 0.006666f
C262 B.n151 VSUBS 0.006666f
C263 B.n152 VSUBS 0.006666f
C264 B.n153 VSUBS 0.006666f
C265 B.n154 VSUBS 0.006666f
C266 B.n155 VSUBS 0.006666f
C267 B.n156 VSUBS 0.006666f
C268 B.n157 VSUBS 0.006666f
C269 B.n158 VSUBS 0.006666f
C270 B.n159 VSUBS 0.006666f
C271 B.t2 VSUBS 0.17857f
C272 B.t1 VSUBS 0.183993f
C273 B.t0 VSUBS 0.100011f
C274 B.n160 VSUBS 0.076468f
C275 B.n161 VSUBS 0.058987f
C276 B.n162 VSUBS 0.015444f
C277 B.n163 VSUBS 0.006274f
C278 B.n164 VSUBS 0.006666f
C279 B.n165 VSUBS 0.006666f
C280 B.n166 VSUBS 0.006666f
C281 B.n167 VSUBS 0.006666f
C282 B.n168 VSUBS 0.006666f
C283 B.n169 VSUBS 0.006666f
C284 B.n170 VSUBS 0.006666f
C285 B.n171 VSUBS 0.006666f
C286 B.n172 VSUBS 0.006666f
C287 B.n173 VSUBS 0.006666f
C288 B.n174 VSUBS 0.006666f
C289 B.n175 VSUBS 0.006666f
C290 B.n176 VSUBS 0.006666f
C291 B.n177 VSUBS 0.006666f
C292 B.n178 VSUBS 0.006666f
C293 B.n179 VSUBS 0.003725f
C294 B.n180 VSUBS 0.015444f
C295 B.n181 VSUBS 0.006274f
C296 B.n182 VSUBS 0.006666f
C297 B.n183 VSUBS 0.006666f
C298 B.n184 VSUBS 0.006666f
C299 B.n185 VSUBS 0.006666f
C300 B.n186 VSUBS 0.006666f
C301 B.n187 VSUBS 0.006666f
C302 B.n188 VSUBS 0.006666f
C303 B.n189 VSUBS 0.006666f
C304 B.n190 VSUBS 0.006666f
C305 B.n191 VSUBS 0.006666f
C306 B.n192 VSUBS 0.006666f
C307 B.n193 VSUBS 0.006666f
C308 B.n194 VSUBS 0.006666f
C309 B.n195 VSUBS 0.006666f
C310 B.n196 VSUBS 0.006666f
C311 B.n197 VSUBS 0.006666f
C312 B.n198 VSUBS 0.006666f
C313 B.n199 VSUBS 0.006666f
C314 B.n200 VSUBS 0.006666f
C315 B.n201 VSUBS 0.006666f
C316 B.n202 VSUBS 0.006666f
C317 B.n203 VSUBS 0.006666f
C318 B.n204 VSUBS 0.006666f
C319 B.n205 VSUBS 0.006666f
C320 B.n206 VSUBS 0.006666f
C321 B.n207 VSUBS 0.006666f
C322 B.n208 VSUBS 0.006666f
C323 B.n209 VSUBS 0.006666f
C324 B.n210 VSUBS 0.006666f
C325 B.n211 VSUBS 0.006666f
C326 B.n212 VSUBS 0.006666f
C327 B.n213 VSUBS 0.006666f
C328 B.n214 VSUBS 0.006666f
C329 B.n215 VSUBS 0.006666f
C330 B.n216 VSUBS 0.006666f
C331 B.n217 VSUBS 0.015343f
C332 B.n218 VSUBS 0.015634f
C333 B.n219 VSUBS 0.014838f
C334 B.n220 VSUBS 0.006666f
C335 B.n221 VSUBS 0.006666f
C336 B.n222 VSUBS 0.006666f
C337 B.n223 VSUBS 0.006666f
C338 B.n224 VSUBS 0.006666f
C339 B.n225 VSUBS 0.006666f
C340 B.n226 VSUBS 0.006666f
C341 B.n227 VSUBS 0.006666f
C342 B.n228 VSUBS 0.006666f
C343 B.n229 VSUBS 0.006666f
C344 B.n230 VSUBS 0.006666f
C345 B.n231 VSUBS 0.006666f
C346 B.n232 VSUBS 0.006666f
C347 B.n233 VSUBS 0.006666f
C348 B.n234 VSUBS 0.006666f
C349 B.n235 VSUBS 0.006666f
C350 B.n236 VSUBS 0.006666f
C351 B.n237 VSUBS 0.006666f
C352 B.n238 VSUBS 0.006666f
C353 B.n239 VSUBS 0.006666f
C354 B.n240 VSUBS 0.006666f
C355 B.n241 VSUBS 0.006666f
C356 B.n242 VSUBS 0.006666f
C357 B.n243 VSUBS 0.006666f
C358 B.n244 VSUBS 0.006666f
C359 B.n245 VSUBS 0.006666f
C360 B.n246 VSUBS 0.006666f
C361 B.n247 VSUBS 0.006666f
C362 B.n248 VSUBS 0.006666f
C363 B.n249 VSUBS 0.006666f
C364 B.n250 VSUBS 0.006666f
C365 B.n251 VSUBS 0.006666f
C366 B.n252 VSUBS 0.006666f
C367 B.n253 VSUBS 0.006666f
C368 B.n254 VSUBS 0.006666f
C369 B.n255 VSUBS 0.006666f
C370 B.n256 VSUBS 0.006666f
C371 B.n257 VSUBS 0.006666f
C372 B.n258 VSUBS 0.006666f
C373 B.n259 VSUBS 0.006666f
C374 B.n260 VSUBS 0.006666f
C375 B.n261 VSUBS 0.006666f
C376 B.n262 VSUBS 0.006666f
C377 B.n263 VSUBS 0.006666f
C378 B.n264 VSUBS 0.006666f
C379 B.n265 VSUBS 0.006666f
C380 B.n266 VSUBS 0.006666f
C381 B.n267 VSUBS 0.006666f
C382 B.n268 VSUBS 0.014838f
C383 B.n269 VSUBS 0.016139f
C384 B.n270 VSUBS 0.016139f
C385 B.n271 VSUBS 0.006666f
C386 B.n272 VSUBS 0.006666f
C387 B.n273 VSUBS 0.006666f
C388 B.n274 VSUBS 0.006666f
C389 B.n275 VSUBS 0.006666f
C390 B.n276 VSUBS 0.006666f
C391 B.n277 VSUBS 0.006666f
C392 B.n278 VSUBS 0.006666f
C393 B.n279 VSUBS 0.006666f
C394 B.n280 VSUBS 0.006666f
C395 B.n281 VSUBS 0.006666f
C396 B.n282 VSUBS 0.006666f
C397 B.n283 VSUBS 0.006666f
C398 B.n284 VSUBS 0.006666f
C399 B.n285 VSUBS 0.006666f
C400 B.n286 VSUBS 0.006666f
C401 B.n287 VSUBS 0.006666f
C402 B.n288 VSUBS 0.006666f
C403 B.n289 VSUBS 0.006666f
C404 B.n290 VSUBS 0.006666f
C405 B.n291 VSUBS 0.006666f
C406 B.n292 VSUBS 0.006666f
C407 B.n293 VSUBS 0.006666f
C408 B.n294 VSUBS 0.006666f
C409 B.n295 VSUBS 0.006666f
C410 B.n296 VSUBS 0.006666f
C411 B.n297 VSUBS 0.006666f
C412 B.n298 VSUBS 0.006666f
C413 B.n299 VSUBS 0.006666f
C414 B.n300 VSUBS 0.006666f
C415 B.n301 VSUBS 0.006666f
C416 B.n302 VSUBS 0.006666f
C417 B.n303 VSUBS 0.006666f
C418 B.n304 VSUBS 0.006666f
C419 B.n305 VSUBS 0.006666f
C420 B.n306 VSUBS 0.006274f
C421 B.n307 VSUBS 0.015444f
C422 B.n308 VSUBS 0.003725f
C423 B.n309 VSUBS 0.006666f
C424 B.n310 VSUBS 0.006666f
C425 B.n311 VSUBS 0.006666f
C426 B.n312 VSUBS 0.006666f
C427 B.n313 VSUBS 0.006666f
C428 B.n314 VSUBS 0.006666f
C429 B.n315 VSUBS 0.006666f
C430 B.n316 VSUBS 0.006666f
C431 B.n317 VSUBS 0.006666f
C432 B.n318 VSUBS 0.006666f
C433 B.n319 VSUBS 0.006666f
C434 B.n320 VSUBS 0.006666f
C435 B.n321 VSUBS 0.003725f
C436 B.n322 VSUBS 0.006666f
C437 B.n323 VSUBS 0.006666f
C438 B.n324 VSUBS 0.006666f
C439 B.n325 VSUBS 0.006666f
C440 B.n326 VSUBS 0.006666f
C441 B.n327 VSUBS 0.006666f
C442 B.n328 VSUBS 0.006666f
C443 B.n329 VSUBS 0.006666f
C444 B.n330 VSUBS 0.006666f
C445 B.n331 VSUBS 0.006666f
C446 B.n332 VSUBS 0.006666f
C447 B.n333 VSUBS 0.006666f
C448 B.n334 VSUBS 0.006666f
C449 B.n335 VSUBS 0.006666f
C450 B.n336 VSUBS 0.006666f
C451 B.n337 VSUBS 0.006666f
C452 B.n338 VSUBS 0.006666f
C453 B.n339 VSUBS 0.006666f
C454 B.n340 VSUBS 0.006666f
C455 B.n341 VSUBS 0.006666f
C456 B.n342 VSUBS 0.006666f
C457 B.n343 VSUBS 0.006666f
C458 B.n344 VSUBS 0.006666f
C459 B.n345 VSUBS 0.006666f
C460 B.n346 VSUBS 0.006666f
C461 B.n347 VSUBS 0.006666f
C462 B.n348 VSUBS 0.006666f
C463 B.n349 VSUBS 0.006666f
C464 B.n350 VSUBS 0.006666f
C465 B.n351 VSUBS 0.006666f
C466 B.n352 VSUBS 0.006666f
C467 B.n353 VSUBS 0.006666f
C468 B.n354 VSUBS 0.006666f
C469 B.n355 VSUBS 0.006666f
C470 B.n356 VSUBS 0.006666f
C471 B.n357 VSUBS 0.006666f
C472 B.n358 VSUBS 0.006666f
C473 B.n359 VSUBS 0.016139f
C474 B.n360 VSUBS 0.014838f
C475 B.n361 VSUBS 0.014838f
C476 B.n362 VSUBS 0.006666f
C477 B.n363 VSUBS 0.006666f
C478 B.n364 VSUBS 0.006666f
C479 B.n365 VSUBS 0.006666f
C480 B.n366 VSUBS 0.006666f
C481 B.n367 VSUBS 0.006666f
C482 B.n368 VSUBS 0.006666f
C483 B.n369 VSUBS 0.006666f
C484 B.n370 VSUBS 0.006666f
C485 B.n371 VSUBS 0.006666f
C486 B.n372 VSUBS 0.006666f
C487 B.n373 VSUBS 0.006666f
C488 B.n374 VSUBS 0.006666f
C489 B.n375 VSUBS 0.006666f
C490 B.n376 VSUBS 0.006666f
C491 B.n377 VSUBS 0.006666f
C492 B.n378 VSUBS 0.006666f
C493 B.n379 VSUBS 0.006666f
C494 B.n380 VSUBS 0.006666f
C495 B.n381 VSUBS 0.006666f
C496 B.n382 VSUBS 0.006666f
C497 B.n383 VSUBS 0.008698f
C498 B.n384 VSUBS 0.009266f
C499 B.n385 VSUBS 0.018427f
.ends

