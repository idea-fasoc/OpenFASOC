* NGSPICE file created from diff_pair_sample_1106.ext - technology: sky130A

.subckt diff_pair_sample_1106 VTAIL VN VP B VDD2 VDD1
X0 B.t21 B.t19 B.t20 B.t9 sky130_fd_pr__nfet_01v8 ad=1.3338 pd=7.62 as=0 ps=0 w=3.42 l=0.45
X1 VTAIL.t14 VN.t0 VDD2.t3 B.t4 sky130_fd_pr__nfet_01v8 ad=0.5643 pd=3.75 as=0.5643 ps=3.75 w=3.42 l=0.45
X2 VDD1.t7 VP.t0 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.5643 pd=3.75 as=1.3338 ps=7.62 w=3.42 l=0.45
X3 VDD1.t6 VP.t1 VTAIL.t4 B.t5 sky130_fd_pr__nfet_01v8 ad=0.5643 pd=3.75 as=0.5643 ps=3.75 w=3.42 l=0.45
X4 VTAIL.t1 VP.t2 VDD1.t5 B.t0 sky130_fd_pr__nfet_01v8 ad=1.3338 pd=7.62 as=0.5643 ps=3.75 w=3.42 l=0.45
X5 VTAIL.t15 VP.t3 VDD1.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=0.5643 pd=3.75 as=0.5643 ps=3.75 w=3.42 l=0.45
X6 B.t18 B.t16 B.t17 B.t13 sky130_fd_pr__nfet_01v8 ad=1.3338 pd=7.62 as=0 ps=0 w=3.42 l=0.45
X7 VDD1.t3 VP.t4 VTAIL.t3 B.t7 sky130_fd_pr__nfet_01v8 ad=0.5643 pd=3.75 as=1.3338 ps=7.62 w=3.42 l=0.45
X8 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=1.3338 pd=7.62 as=0 ps=0 w=3.42 l=0.45
X9 VTAIL.t0 VP.t5 VDD1.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=1.3338 pd=7.62 as=0.5643 ps=3.75 w=3.42 l=0.45
X10 VTAIL.t13 VN.t1 VDD2.t7 B.t0 sky130_fd_pr__nfet_01v8 ad=1.3338 pd=7.62 as=0.5643 ps=3.75 w=3.42 l=0.45
X11 VDD2.t5 VN.t2 VTAIL.t12 B.t2 sky130_fd_pr__nfet_01v8 ad=0.5643 pd=3.75 as=1.3338 ps=7.62 w=3.42 l=0.45
X12 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=1.3338 pd=7.62 as=0 ps=0 w=3.42 l=0.45
X13 VDD2.t0 VN.t3 VTAIL.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=0.5643 pd=3.75 as=1.3338 ps=7.62 w=3.42 l=0.45
X14 VTAIL.t5 VP.t6 VDD1.t1 B.t6 sky130_fd_pr__nfet_01v8 ad=0.5643 pd=3.75 as=0.5643 ps=3.75 w=3.42 l=0.45
X15 VTAIL.t10 VN.t4 VDD2.t4 B.t6 sky130_fd_pr__nfet_01v8 ad=0.5643 pd=3.75 as=0.5643 ps=3.75 w=3.42 l=0.45
X16 VDD2.t6 VN.t5 VTAIL.t9 B.t3 sky130_fd_pr__nfet_01v8 ad=0.5643 pd=3.75 as=0.5643 ps=3.75 w=3.42 l=0.45
X17 VTAIL.t8 VN.t6 VDD2.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=1.3338 pd=7.62 as=0.5643 ps=3.75 w=3.42 l=0.45
X18 VDD2.t1 VN.t7 VTAIL.t7 B.t5 sky130_fd_pr__nfet_01v8 ad=0.5643 pd=3.75 as=0.5643 ps=3.75 w=3.42 l=0.45
X19 VDD1.t0 VP.t7 VTAIL.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=0.5643 pd=3.75 as=0.5643 ps=3.75 w=3.42 l=0.45
R0 B.n375 B.n374 585
R1 B.n144 B.n60 585
R2 B.n143 B.n142 585
R3 B.n141 B.n140 585
R4 B.n139 B.n138 585
R5 B.n137 B.n136 585
R6 B.n135 B.n134 585
R7 B.n133 B.n132 585
R8 B.n131 B.n130 585
R9 B.n129 B.n128 585
R10 B.n127 B.n126 585
R11 B.n125 B.n124 585
R12 B.n123 B.n122 585
R13 B.n121 B.n120 585
R14 B.n119 B.n118 585
R15 B.n117 B.n116 585
R16 B.n115 B.n114 585
R17 B.n113 B.n112 585
R18 B.n111 B.n110 585
R19 B.n109 B.n108 585
R20 B.n107 B.n106 585
R21 B.n105 B.n104 585
R22 B.n103 B.n102 585
R23 B.n101 B.n100 585
R24 B.n99 B.n98 585
R25 B.n97 B.n96 585
R26 B.n95 B.n94 585
R27 B.n93 B.n92 585
R28 B.n91 B.n90 585
R29 B.n89 B.n88 585
R30 B.n87 B.n86 585
R31 B.n85 B.n84 585
R32 B.n83 B.n82 585
R33 B.n81 B.n80 585
R34 B.n79 B.n78 585
R35 B.n77 B.n76 585
R36 B.n75 B.n74 585
R37 B.n73 B.n72 585
R38 B.n71 B.n70 585
R39 B.n69 B.n68 585
R40 B.n40 B.n39 585
R41 B.n380 B.n379 585
R42 B.n373 B.n61 585
R43 B.n61 B.n37 585
R44 B.n372 B.n36 585
R45 B.n384 B.n36 585
R46 B.n371 B.n35 585
R47 B.n385 B.n35 585
R48 B.n370 B.n34 585
R49 B.n386 B.n34 585
R50 B.n369 B.n368 585
R51 B.n368 B.n33 585
R52 B.n367 B.n29 585
R53 B.n392 B.n29 585
R54 B.n366 B.n28 585
R55 B.n393 B.n28 585
R56 B.n365 B.n27 585
R57 B.n394 B.n27 585
R58 B.n364 B.n363 585
R59 B.n363 B.n23 585
R60 B.n362 B.n22 585
R61 B.n400 B.n22 585
R62 B.n361 B.n21 585
R63 B.n401 B.n21 585
R64 B.n360 B.n20 585
R65 B.n402 B.n20 585
R66 B.n359 B.n358 585
R67 B.n358 B.n19 585
R68 B.n357 B.n15 585
R69 B.n408 B.n15 585
R70 B.n356 B.n14 585
R71 B.n409 B.n14 585
R72 B.n355 B.n13 585
R73 B.n410 B.n13 585
R74 B.n354 B.n353 585
R75 B.n353 B.n12 585
R76 B.n352 B.n351 585
R77 B.n352 B.n8 585
R78 B.n350 B.n7 585
R79 B.n417 B.n7 585
R80 B.n349 B.n6 585
R81 B.n418 B.n6 585
R82 B.n348 B.n5 585
R83 B.n419 B.n5 585
R84 B.n347 B.n346 585
R85 B.n346 B.n4 585
R86 B.n345 B.n145 585
R87 B.n345 B.n344 585
R88 B.n334 B.n146 585
R89 B.n337 B.n146 585
R90 B.n336 B.n335 585
R91 B.n338 B.n336 585
R92 B.n333 B.n150 585
R93 B.n153 B.n150 585
R94 B.n332 B.n331 585
R95 B.n331 B.n330 585
R96 B.n152 B.n151 585
R97 B.n323 B.n152 585
R98 B.n322 B.n321 585
R99 B.n324 B.n322 585
R100 B.n320 B.n158 585
R101 B.n158 B.n157 585
R102 B.n319 B.n318 585
R103 B.n318 B.n317 585
R104 B.n160 B.n159 585
R105 B.n161 B.n160 585
R106 B.n310 B.n309 585
R107 B.n311 B.n310 585
R108 B.n308 B.n166 585
R109 B.n166 B.n165 585
R110 B.n307 B.n306 585
R111 B.n306 B.n305 585
R112 B.n168 B.n167 585
R113 B.n298 B.n168 585
R114 B.n297 B.n296 585
R115 B.n299 B.n297 585
R116 B.n295 B.n173 585
R117 B.n173 B.n172 585
R118 B.n294 B.n293 585
R119 B.n293 B.n292 585
R120 B.n175 B.n174 585
R121 B.n176 B.n175 585
R122 B.n288 B.n287 585
R123 B.n179 B.n178 585
R124 B.n284 B.n283 585
R125 B.n285 B.n284 585
R126 B.n282 B.n200 585
R127 B.n281 B.n280 585
R128 B.n279 B.n278 585
R129 B.n277 B.n276 585
R130 B.n275 B.n274 585
R131 B.n273 B.n272 585
R132 B.n271 B.n270 585
R133 B.n269 B.n268 585
R134 B.n267 B.n266 585
R135 B.n265 B.n264 585
R136 B.n263 B.n262 585
R137 B.n261 B.n260 585
R138 B.n259 B.n258 585
R139 B.n256 B.n255 585
R140 B.n254 B.n253 585
R141 B.n252 B.n251 585
R142 B.n250 B.n249 585
R143 B.n248 B.n247 585
R144 B.n246 B.n245 585
R145 B.n244 B.n243 585
R146 B.n242 B.n241 585
R147 B.n240 B.n239 585
R148 B.n238 B.n237 585
R149 B.n235 B.n234 585
R150 B.n233 B.n232 585
R151 B.n231 B.n230 585
R152 B.n229 B.n228 585
R153 B.n227 B.n226 585
R154 B.n225 B.n224 585
R155 B.n223 B.n222 585
R156 B.n221 B.n220 585
R157 B.n219 B.n218 585
R158 B.n217 B.n216 585
R159 B.n215 B.n214 585
R160 B.n213 B.n212 585
R161 B.n211 B.n210 585
R162 B.n209 B.n208 585
R163 B.n207 B.n206 585
R164 B.n205 B.n199 585
R165 B.n285 B.n199 585
R166 B.n289 B.n177 585
R167 B.n177 B.n176 585
R168 B.n291 B.n290 585
R169 B.n292 B.n291 585
R170 B.n171 B.n170 585
R171 B.n172 B.n171 585
R172 B.n301 B.n300 585
R173 B.n300 B.n299 585
R174 B.n302 B.n169 585
R175 B.n298 B.n169 585
R176 B.n304 B.n303 585
R177 B.n305 B.n304 585
R178 B.n164 B.n163 585
R179 B.n165 B.n164 585
R180 B.n313 B.n312 585
R181 B.n312 B.n311 585
R182 B.n314 B.n162 585
R183 B.n162 B.n161 585
R184 B.n316 B.n315 585
R185 B.n317 B.n316 585
R186 B.n156 B.n155 585
R187 B.n157 B.n156 585
R188 B.n326 B.n325 585
R189 B.n325 B.n324 585
R190 B.n327 B.n154 585
R191 B.n323 B.n154 585
R192 B.n329 B.n328 585
R193 B.n330 B.n329 585
R194 B.n149 B.n148 585
R195 B.n153 B.n149 585
R196 B.n340 B.n339 585
R197 B.n339 B.n338 585
R198 B.n341 B.n147 585
R199 B.n337 B.n147 585
R200 B.n343 B.n342 585
R201 B.n344 B.n343 585
R202 B.n3 B.n0 585
R203 B.n4 B.n3 585
R204 B.n416 B.n1 585
R205 B.n417 B.n416 585
R206 B.n415 B.n414 585
R207 B.n415 B.n8 585
R208 B.n413 B.n9 585
R209 B.n12 B.n9 585
R210 B.n412 B.n411 585
R211 B.n411 B.n410 585
R212 B.n11 B.n10 585
R213 B.n409 B.n11 585
R214 B.n407 B.n406 585
R215 B.n408 B.n407 585
R216 B.n405 B.n16 585
R217 B.n19 B.n16 585
R218 B.n404 B.n403 585
R219 B.n403 B.n402 585
R220 B.n18 B.n17 585
R221 B.n401 B.n18 585
R222 B.n399 B.n398 585
R223 B.n400 B.n399 585
R224 B.n397 B.n24 585
R225 B.n24 B.n23 585
R226 B.n396 B.n395 585
R227 B.n395 B.n394 585
R228 B.n26 B.n25 585
R229 B.n393 B.n26 585
R230 B.n391 B.n390 585
R231 B.n392 B.n391 585
R232 B.n389 B.n30 585
R233 B.n33 B.n30 585
R234 B.n388 B.n387 585
R235 B.n387 B.n386 585
R236 B.n32 B.n31 585
R237 B.n385 B.n32 585
R238 B.n383 B.n382 585
R239 B.n384 B.n383 585
R240 B.n381 B.n38 585
R241 B.n38 B.n37 585
R242 B.n420 B.n419 585
R243 B.n418 B.n2 585
R244 B.n379 B.n38 540.549
R245 B.n375 B.n61 540.549
R246 B.n199 B.n175 540.549
R247 B.n287 B.n177 540.549
R248 B.n65 B.t16 390.906
R249 B.n62 B.t12 390.906
R250 B.n203 B.t19 390.906
R251 B.n201 B.t8 390.906
R252 B.n377 B.n376 256.663
R253 B.n377 B.n59 256.663
R254 B.n377 B.n58 256.663
R255 B.n377 B.n57 256.663
R256 B.n377 B.n56 256.663
R257 B.n377 B.n55 256.663
R258 B.n377 B.n54 256.663
R259 B.n377 B.n53 256.663
R260 B.n377 B.n52 256.663
R261 B.n377 B.n51 256.663
R262 B.n377 B.n50 256.663
R263 B.n377 B.n49 256.663
R264 B.n377 B.n48 256.663
R265 B.n377 B.n47 256.663
R266 B.n377 B.n46 256.663
R267 B.n377 B.n45 256.663
R268 B.n377 B.n44 256.663
R269 B.n377 B.n43 256.663
R270 B.n377 B.n42 256.663
R271 B.n377 B.n41 256.663
R272 B.n378 B.n377 256.663
R273 B.n286 B.n285 256.663
R274 B.n285 B.n180 256.663
R275 B.n285 B.n181 256.663
R276 B.n285 B.n182 256.663
R277 B.n285 B.n183 256.663
R278 B.n285 B.n184 256.663
R279 B.n285 B.n185 256.663
R280 B.n285 B.n186 256.663
R281 B.n285 B.n187 256.663
R282 B.n285 B.n188 256.663
R283 B.n285 B.n189 256.663
R284 B.n285 B.n190 256.663
R285 B.n285 B.n191 256.663
R286 B.n285 B.n192 256.663
R287 B.n285 B.n193 256.663
R288 B.n285 B.n194 256.663
R289 B.n285 B.n195 256.663
R290 B.n285 B.n196 256.663
R291 B.n285 B.n197 256.663
R292 B.n285 B.n198 256.663
R293 B.n422 B.n421 256.663
R294 B.n68 B.n40 163.367
R295 B.n72 B.n71 163.367
R296 B.n76 B.n75 163.367
R297 B.n80 B.n79 163.367
R298 B.n84 B.n83 163.367
R299 B.n88 B.n87 163.367
R300 B.n92 B.n91 163.367
R301 B.n96 B.n95 163.367
R302 B.n100 B.n99 163.367
R303 B.n104 B.n103 163.367
R304 B.n108 B.n107 163.367
R305 B.n112 B.n111 163.367
R306 B.n116 B.n115 163.367
R307 B.n120 B.n119 163.367
R308 B.n124 B.n123 163.367
R309 B.n128 B.n127 163.367
R310 B.n132 B.n131 163.367
R311 B.n136 B.n135 163.367
R312 B.n140 B.n139 163.367
R313 B.n142 B.n60 163.367
R314 B.n293 B.n175 163.367
R315 B.n293 B.n173 163.367
R316 B.n297 B.n173 163.367
R317 B.n297 B.n168 163.367
R318 B.n306 B.n168 163.367
R319 B.n306 B.n166 163.367
R320 B.n310 B.n166 163.367
R321 B.n310 B.n160 163.367
R322 B.n318 B.n160 163.367
R323 B.n318 B.n158 163.367
R324 B.n322 B.n158 163.367
R325 B.n322 B.n152 163.367
R326 B.n331 B.n152 163.367
R327 B.n331 B.n150 163.367
R328 B.n336 B.n150 163.367
R329 B.n336 B.n146 163.367
R330 B.n345 B.n146 163.367
R331 B.n346 B.n345 163.367
R332 B.n346 B.n5 163.367
R333 B.n6 B.n5 163.367
R334 B.n7 B.n6 163.367
R335 B.n352 B.n7 163.367
R336 B.n353 B.n352 163.367
R337 B.n353 B.n13 163.367
R338 B.n14 B.n13 163.367
R339 B.n15 B.n14 163.367
R340 B.n358 B.n15 163.367
R341 B.n358 B.n20 163.367
R342 B.n21 B.n20 163.367
R343 B.n22 B.n21 163.367
R344 B.n363 B.n22 163.367
R345 B.n363 B.n27 163.367
R346 B.n28 B.n27 163.367
R347 B.n29 B.n28 163.367
R348 B.n368 B.n29 163.367
R349 B.n368 B.n34 163.367
R350 B.n35 B.n34 163.367
R351 B.n36 B.n35 163.367
R352 B.n61 B.n36 163.367
R353 B.n284 B.n179 163.367
R354 B.n284 B.n200 163.367
R355 B.n280 B.n279 163.367
R356 B.n276 B.n275 163.367
R357 B.n272 B.n271 163.367
R358 B.n268 B.n267 163.367
R359 B.n264 B.n263 163.367
R360 B.n260 B.n259 163.367
R361 B.n255 B.n254 163.367
R362 B.n251 B.n250 163.367
R363 B.n247 B.n246 163.367
R364 B.n243 B.n242 163.367
R365 B.n239 B.n238 163.367
R366 B.n234 B.n233 163.367
R367 B.n230 B.n229 163.367
R368 B.n226 B.n225 163.367
R369 B.n222 B.n221 163.367
R370 B.n218 B.n217 163.367
R371 B.n214 B.n213 163.367
R372 B.n210 B.n209 163.367
R373 B.n206 B.n199 163.367
R374 B.n291 B.n177 163.367
R375 B.n291 B.n171 163.367
R376 B.n300 B.n171 163.367
R377 B.n300 B.n169 163.367
R378 B.n304 B.n169 163.367
R379 B.n304 B.n164 163.367
R380 B.n312 B.n164 163.367
R381 B.n312 B.n162 163.367
R382 B.n316 B.n162 163.367
R383 B.n316 B.n156 163.367
R384 B.n325 B.n156 163.367
R385 B.n325 B.n154 163.367
R386 B.n329 B.n154 163.367
R387 B.n329 B.n149 163.367
R388 B.n339 B.n149 163.367
R389 B.n339 B.n147 163.367
R390 B.n343 B.n147 163.367
R391 B.n343 B.n3 163.367
R392 B.n420 B.n3 163.367
R393 B.n416 B.n2 163.367
R394 B.n416 B.n415 163.367
R395 B.n415 B.n9 163.367
R396 B.n411 B.n9 163.367
R397 B.n411 B.n11 163.367
R398 B.n407 B.n11 163.367
R399 B.n407 B.n16 163.367
R400 B.n403 B.n16 163.367
R401 B.n403 B.n18 163.367
R402 B.n399 B.n18 163.367
R403 B.n399 B.n24 163.367
R404 B.n395 B.n24 163.367
R405 B.n395 B.n26 163.367
R406 B.n391 B.n26 163.367
R407 B.n391 B.n30 163.367
R408 B.n387 B.n30 163.367
R409 B.n387 B.n32 163.367
R410 B.n383 B.n32 163.367
R411 B.n383 B.n38 163.367
R412 B.n285 B.n176 163.197
R413 B.n377 B.n37 163.197
R414 B.n62 B.t14 88.2662
R415 B.n203 B.t21 88.2662
R416 B.n65 B.t17 88.2633
R417 B.n201 B.t11 88.2633
R418 B.n292 B.n176 86.027
R419 B.n292 B.n172 86.027
R420 B.n299 B.n172 86.027
R421 B.n299 B.n298 86.027
R422 B.n305 B.n165 86.027
R423 B.n311 B.n165 86.027
R424 B.n311 B.n161 86.027
R425 B.n317 B.n161 86.027
R426 B.n324 B.n157 86.027
R427 B.n324 B.n323 86.027
R428 B.n330 B.n153 86.027
R429 B.n338 B.n337 86.027
R430 B.n344 B.n4 86.027
R431 B.n419 B.n4 86.027
R432 B.n419 B.n418 86.027
R433 B.n418 B.n417 86.027
R434 B.n417 B.n8 86.027
R435 B.n410 B.n12 86.027
R436 B.n409 B.n408 86.027
R437 B.n402 B.n19 86.027
R438 B.n402 B.n401 86.027
R439 B.n400 B.n23 86.027
R440 B.n394 B.n23 86.027
R441 B.n394 B.n393 86.027
R442 B.n393 B.n392 86.027
R443 B.n386 B.n33 86.027
R444 B.n386 B.n385 86.027
R445 B.n385 B.n384 86.027
R446 B.n384 B.n37 86.027
R447 B.n317 B.t0 74.6411
R448 B.t2 B.n400 74.6411
R449 B.n63 B.t15 73.1389
R450 B.n204 B.t20 73.1389
R451 B.n66 B.t18 73.136
R452 B.n202 B.t10 73.136
R453 B.n330 B.t5 72.1109
R454 B.n408 B.t6 72.1109
R455 B.n379 B.n378 71.676
R456 B.n68 B.n41 71.676
R457 B.n72 B.n42 71.676
R458 B.n76 B.n43 71.676
R459 B.n80 B.n44 71.676
R460 B.n84 B.n45 71.676
R461 B.n88 B.n46 71.676
R462 B.n92 B.n47 71.676
R463 B.n96 B.n48 71.676
R464 B.n100 B.n49 71.676
R465 B.n104 B.n50 71.676
R466 B.n108 B.n51 71.676
R467 B.n112 B.n52 71.676
R468 B.n116 B.n53 71.676
R469 B.n120 B.n54 71.676
R470 B.n124 B.n55 71.676
R471 B.n128 B.n56 71.676
R472 B.n132 B.n57 71.676
R473 B.n136 B.n58 71.676
R474 B.n140 B.n59 71.676
R475 B.n376 B.n60 71.676
R476 B.n376 B.n375 71.676
R477 B.n142 B.n59 71.676
R478 B.n139 B.n58 71.676
R479 B.n135 B.n57 71.676
R480 B.n131 B.n56 71.676
R481 B.n127 B.n55 71.676
R482 B.n123 B.n54 71.676
R483 B.n119 B.n53 71.676
R484 B.n115 B.n52 71.676
R485 B.n111 B.n51 71.676
R486 B.n107 B.n50 71.676
R487 B.n103 B.n49 71.676
R488 B.n99 B.n48 71.676
R489 B.n95 B.n47 71.676
R490 B.n91 B.n46 71.676
R491 B.n87 B.n45 71.676
R492 B.n83 B.n44 71.676
R493 B.n79 B.n43 71.676
R494 B.n75 B.n42 71.676
R495 B.n71 B.n41 71.676
R496 B.n378 B.n40 71.676
R497 B.n287 B.n286 71.676
R498 B.n200 B.n180 71.676
R499 B.n279 B.n181 71.676
R500 B.n275 B.n182 71.676
R501 B.n271 B.n183 71.676
R502 B.n267 B.n184 71.676
R503 B.n263 B.n185 71.676
R504 B.n259 B.n186 71.676
R505 B.n254 B.n187 71.676
R506 B.n250 B.n188 71.676
R507 B.n246 B.n189 71.676
R508 B.n242 B.n190 71.676
R509 B.n238 B.n191 71.676
R510 B.n233 B.n192 71.676
R511 B.n229 B.n193 71.676
R512 B.n225 B.n194 71.676
R513 B.n221 B.n195 71.676
R514 B.n217 B.n196 71.676
R515 B.n213 B.n197 71.676
R516 B.n209 B.n198 71.676
R517 B.n286 B.n179 71.676
R518 B.n280 B.n180 71.676
R519 B.n276 B.n181 71.676
R520 B.n272 B.n182 71.676
R521 B.n268 B.n183 71.676
R522 B.n264 B.n184 71.676
R523 B.n260 B.n185 71.676
R524 B.n255 B.n186 71.676
R525 B.n251 B.n187 71.676
R526 B.n247 B.n188 71.676
R527 B.n243 B.n189 71.676
R528 B.n239 B.n190 71.676
R529 B.n234 B.n191 71.676
R530 B.n230 B.n192 71.676
R531 B.n226 B.n193 71.676
R532 B.n222 B.n194 71.676
R533 B.n218 B.n195 71.676
R534 B.n214 B.n196 71.676
R535 B.n210 B.n197 71.676
R536 B.n206 B.n198 71.676
R537 B.n421 B.n420 71.676
R538 B.n421 B.n2 71.676
R539 B.n337 B.t7 64.5203
R540 B.n12 B.t1 64.5203
R541 B.n67 B.n66 59.5399
R542 B.n64 B.n63 59.5399
R543 B.n236 B.n204 59.5399
R544 B.n257 B.n202 59.5399
R545 B.n305 B.t9 54.3996
R546 B.n392 B.t13 54.3996
R547 B.n338 B.t4 46.809
R548 B.n410 B.t3 46.809
R549 B.n153 B.t4 39.2184
R550 B.t3 B.n409 39.2184
R551 B.n289 B.n288 35.1225
R552 B.n205 B.n174 35.1225
R553 B.n381 B.n380 35.1225
R554 B.n374 B.n373 35.1224
R555 B.n298 B.t9 31.6279
R556 B.n33 B.t13 31.6279
R557 B.n344 B.t7 21.5071
R558 B.t1 B.n8 21.5071
R559 B B.n422 18.0485
R560 B.n66 B.n65 15.1278
R561 B.n63 B.n62 15.1278
R562 B.n204 B.n203 15.1278
R563 B.n202 B.n201 15.1278
R564 B.n323 B.t5 13.9165
R565 B.n19 B.t6 13.9165
R566 B.t0 B.n157 11.3864
R567 B.n401 B.t2 11.3864
R568 B.n290 B.n289 10.6151
R569 B.n290 B.n170 10.6151
R570 B.n301 B.n170 10.6151
R571 B.n302 B.n301 10.6151
R572 B.n303 B.n302 10.6151
R573 B.n303 B.n163 10.6151
R574 B.n313 B.n163 10.6151
R575 B.n314 B.n313 10.6151
R576 B.n315 B.n314 10.6151
R577 B.n315 B.n155 10.6151
R578 B.n326 B.n155 10.6151
R579 B.n327 B.n326 10.6151
R580 B.n328 B.n327 10.6151
R581 B.n328 B.n148 10.6151
R582 B.n340 B.n148 10.6151
R583 B.n341 B.n340 10.6151
R584 B.n342 B.n341 10.6151
R585 B.n342 B.n0 10.6151
R586 B.n288 B.n178 10.6151
R587 B.n283 B.n178 10.6151
R588 B.n283 B.n282 10.6151
R589 B.n282 B.n281 10.6151
R590 B.n281 B.n278 10.6151
R591 B.n278 B.n277 10.6151
R592 B.n277 B.n274 10.6151
R593 B.n274 B.n273 10.6151
R594 B.n273 B.n270 10.6151
R595 B.n270 B.n269 10.6151
R596 B.n269 B.n266 10.6151
R597 B.n266 B.n265 10.6151
R598 B.n265 B.n262 10.6151
R599 B.n262 B.n261 10.6151
R600 B.n261 B.n258 10.6151
R601 B.n256 B.n253 10.6151
R602 B.n253 B.n252 10.6151
R603 B.n252 B.n249 10.6151
R604 B.n249 B.n248 10.6151
R605 B.n248 B.n245 10.6151
R606 B.n245 B.n244 10.6151
R607 B.n244 B.n241 10.6151
R608 B.n241 B.n240 10.6151
R609 B.n240 B.n237 10.6151
R610 B.n235 B.n232 10.6151
R611 B.n232 B.n231 10.6151
R612 B.n231 B.n228 10.6151
R613 B.n228 B.n227 10.6151
R614 B.n227 B.n224 10.6151
R615 B.n224 B.n223 10.6151
R616 B.n223 B.n220 10.6151
R617 B.n220 B.n219 10.6151
R618 B.n219 B.n216 10.6151
R619 B.n216 B.n215 10.6151
R620 B.n215 B.n212 10.6151
R621 B.n212 B.n211 10.6151
R622 B.n211 B.n208 10.6151
R623 B.n208 B.n207 10.6151
R624 B.n207 B.n205 10.6151
R625 B.n294 B.n174 10.6151
R626 B.n295 B.n294 10.6151
R627 B.n296 B.n295 10.6151
R628 B.n296 B.n167 10.6151
R629 B.n307 B.n167 10.6151
R630 B.n308 B.n307 10.6151
R631 B.n309 B.n308 10.6151
R632 B.n309 B.n159 10.6151
R633 B.n319 B.n159 10.6151
R634 B.n320 B.n319 10.6151
R635 B.n321 B.n320 10.6151
R636 B.n321 B.n151 10.6151
R637 B.n332 B.n151 10.6151
R638 B.n333 B.n332 10.6151
R639 B.n335 B.n333 10.6151
R640 B.n335 B.n334 10.6151
R641 B.n334 B.n145 10.6151
R642 B.n347 B.n145 10.6151
R643 B.n348 B.n347 10.6151
R644 B.n349 B.n348 10.6151
R645 B.n350 B.n349 10.6151
R646 B.n351 B.n350 10.6151
R647 B.n354 B.n351 10.6151
R648 B.n355 B.n354 10.6151
R649 B.n356 B.n355 10.6151
R650 B.n357 B.n356 10.6151
R651 B.n359 B.n357 10.6151
R652 B.n360 B.n359 10.6151
R653 B.n361 B.n360 10.6151
R654 B.n362 B.n361 10.6151
R655 B.n364 B.n362 10.6151
R656 B.n365 B.n364 10.6151
R657 B.n366 B.n365 10.6151
R658 B.n367 B.n366 10.6151
R659 B.n369 B.n367 10.6151
R660 B.n370 B.n369 10.6151
R661 B.n371 B.n370 10.6151
R662 B.n372 B.n371 10.6151
R663 B.n373 B.n372 10.6151
R664 B.n414 B.n1 10.6151
R665 B.n414 B.n413 10.6151
R666 B.n413 B.n412 10.6151
R667 B.n412 B.n10 10.6151
R668 B.n406 B.n10 10.6151
R669 B.n406 B.n405 10.6151
R670 B.n405 B.n404 10.6151
R671 B.n404 B.n17 10.6151
R672 B.n398 B.n17 10.6151
R673 B.n398 B.n397 10.6151
R674 B.n397 B.n396 10.6151
R675 B.n396 B.n25 10.6151
R676 B.n390 B.n25 10.6151
R677 B.n390 B.n389 10.6151
R678 B.n389 B.n388 10.6151
R679 B.n388 B.n31 10.6151
R680 B.n382 B.n31 10.6151
R681 B.n382 B.n381 10.6151
R682 B.n380 B.n39 10.6151
R683 B.n69 B.n39 10.6151
R684 B.n70 B.n69 10.6151
R685 B.n73 B.n70 10.6151
R686 B.n74 B.n73 10.6151
R687 B.n77 B.n74 10.6151
R688 B.n78 B.n77 10.6151
R689 B.n81 B.n78 10.6151
R690 B.n82 B.n81 10.6151
R691 B.n85 B.n82 10.6151
R692 B.n86 B.n85 10.6151
R693 B.n89 B.n86 10.6151
R694 B.n90 B.n89 10.6151
R695 B.n93 B.n90 10.6151
R696 B.n94 B.n93 10.6151
R697 B.n98 B.n97 10.6151
R698 B.n101 B.n98 10.6151
R699 B.n102 B.n101 10.6151
R700 B.n105 B.n102 10.6151
R701 B.n106 B.n105 10.6151
R702 B.n109 B.n106 10.6151
R703 B.n110 B.n109 10.6151
R704 B.n113 B.n110 10.6151
R705 B.n114 B.n113 10.6151
R706 B.n118 B.n117 10.6151
R707 B.n121 B.n118 10.6151
R708 B.n122 B.n121 10.6151
R709 B.n125 B.n122 10.6151
R710 B.n126 B.n125 10.6151
R711 B.n129 B.n126 10.6151
R712 B.n130 B.n129 10.6151
R713 B.n133 B.n130 10.6151
R714 B.n134 B.n133 10.6151
R715 B.n137 B.n134 10.6151
R716 B.n138 B.n137 10.6151
R717 B.n141 B.n138 10.6151
R718 B.n143 B.n141 10.6151
R719 B.n144 B.n143 10.6151
R720 B.n374 B.n144 10.6151
R721 B.n258 B.n257 9.36635
R722 B.n236 B.n235 9.36635
R723 B.n94 B.n67 9.36635
R724 B.n117 B.n64 9.36635
R725 B.n422 B.n0 8.11757
R726 B.n422 B.n1 8.11757
R727 B.n257 B.n256 1.24928
R728 B.n237 B.n236 1.24928
R729 B.n97 B.n67 1.24928
R730 B.n114 B.n64 1.24928
R731 VN.n2 VN.t6 291.438
R732 VN.n10 VN.t3 291.438
R733 VN.n1 VN.t5 270.457
R734 VN.n5 VN.t4 270.457
R735 VN.n6 VN.t2 270.457
R736 VN.n9 VN.t0 270.457
R737 VN.n13 VN.t7 270.457
R738 VN.n14 VN.t1 270.457
R739 VN.n7 VN.n6 161.3
R740 VN.n15 VN.n14 161.3
R741 VN.n13 VN.n8 161.3
R742 VN.n12 VN.n11 161.3
R743 VN.n5 VN.n0 161.3
R744 VN.n4 VN.n3 161.3
R745 VN.n11 VN.n10 70.4033
R746 VN.n3 VN.n2 70.4033
R747 VN.n6 VN.n5 48.2005
R748 VN.n14 VN.n13 48.2005
R749 VN VN.n15 34.7372
R750 VN.n4 VN.n1 24.1005
R751 VN.n5 VN.n4 24.1005
R752 VN.n13 VN.n12 24.1005
R753 VN.n12 VN.n9 24.1005
R754 VN.n10 VN.n9 20.9576
R755 VN.n2 VN.n1 20.9576
R756 VN.n15 VN.n8 0.189894
R757 VN.n11 VN.n8 0.189894
R758 VN.n3 VN.n0 0.189894
R759 VN.n7 VN.n0 0.189894
R760 VN VN.n7 0.0516364
R761 VDD2.n2 VDD2.n1 74.4776
R762 VDD2.n2 VDD2.n0 74.4776
R763 VDD2 VDD2.n5 74.4749
R764 VDD2.n4 VDD2.n3 74.197
R765 VDD2.n4 VDD2.n2 29.6894
R766 VDD2.n5 VDD2.t3 5.78997
R767 VDD2.n5 VDD2.t0 5.78997
R768 VDD2.n3 VDD2.t7 5.78997
R769 VDD2.n3 VDD2.t1 5.78997
R770 VDD2.n1 VDD2.t4 5.78997
R771 VDD2.n1 VDD2.t5 5.78997
R772 VDD2.n0 VDD2.t2 5.78997
R773 VDD2.n0 VDD2.t6 5.78997
R774 VDD2 VDD2.n4 0.394897
R775 VTAIL.n11 VTAIL.t0 63.3076
R776 VTAIL.n10 VTAIL.t11 63.3076
R777 VTAIL.n7 VTAIL.t13 63.3076
R778 VTAIL.n15 VTAIL.t12 63.3076
R779 VTAIL.n2 VTAIL.t8 63.3076
R780 VTAIL.n3 VTAIL.t3 63.3076
R781 VTAIL.n6 VTAIL.t1 63.3076
R782 VTAIL.n14 VTAIL.t2 63.3076
R783 VTAIL.n13 VTAIL.n12 57.5182
R784 VTAIL.n9 VTAIL.n8 57.5182
R785 VTAIL.n1 VTAIL.n0 57.518
R786 VTAIL.n5 VTAIL.n4 57.518
R787 VTAIL.n15 VTAIL.n14 15.9876
R788 VTAIL.n7 VTAIL.n6 15.9876
R789 VTAIL.n0 VTAIL.t9 5.78997
R790 VTAIL.n0 VTAIL.t10 5.78997
R791 VTAIL.n4 VTAIL.t4 5.78997
R792 VTAIL.n4 VTAIL.t15 5.78997
R793 VTAIL.n12 VTAIL.t6 5.78997
R794 VTAIL.n12 VTAIL.t5 5.78997
R795 VTAIL.n8 VTAIL.t7 5.78997
R796 VTAIL.n8 VTAIL.t14 5.78997
R797 VTAIL.n9 VTAIL.n7 0.672914
R798 VTAIL.n10 VTAIL.n9 0.672914
R799 VTAIL.n13 VTAIL.n11 0.672914
R800 VTAIL.n14 VTAIL.n13 0.672914
R801 VTAIL.n6 VTAIL.n5 0.672914
R802 VTAIL.n5 VTAIL.n3 0.672914
R803 VTAIL.n2 VTAIL.n1 0.672914
R804 VTAIL VTAIL.n15 0.614724
R805 VTAIL.n11 VTAIL.n10 0.470328
R806 VTAIL.n3 VTAIL.n2 0.470328
R807 VTAIL VTAIL.n1 0.0586897
R808 VP.n4 VP.t5 291.438
R809 VP.n10 VP.t2 270.457
R810 VP.n1 VP.t1 270.457
R811 VP.n15 VP.t3 270.457
R812 VP.n16 VP.t4 270.457
R813 VP.n8 VP.t0 270.457
R814 VP.n7 VP.t6 270.457
R815 VP.n3 VP.t7 270.457
R816 VP.n17 VP.n16 161.3
R817 VP.n6 VP.n5 161.3
R818 VP.n7 VP.n2 161.3
R819 VP.n9 VP.n8 161.3
R820 VP.n15 VP.n0 161.3
R821 VP.n14 VP.n13 161.3
R822 VP.n12 VP.n1 161.3
R823 VP.n11 VP.n10 161.3
R824 VP.n5 VP.n4 70.4033
R825 VP.n10 VP.n1 48.2005
R826 VP.n16 VP.n15 48.2005
R827 VP.n8 VP.n7 48.2005
R828 VP.n11 VP.n9 34.3566
R829 VP.n14 VP.n1 24.1005
R830 VP.n15 VP.n14 24.1005
R831 VP.n6 VP.n3 24.1005
R832 VP.n7 VP.n6 24.1005
R833 VP.n4 VP.n3 20.9576
R834 VP.n5 VP.n2 0.189894
R835 VP.n9 VP.n2 0.189894
R836 VP.n12 VP.n11 0.189894
R837 VP.n13 VP.n12 0.189894
R838 VP.n13 VP.n0 0.189894
R839 VP.n17 VP.n0 0.189894
R840 VP VP.n17 0.0516364
R841 VDD1 VDD1.n0 74.5914
R842 VDD1.n3 VDD1.n2 74.4776
R843 VDD1.n3 VDD1.n1 74.4776
R844 VDD1.n5 VDD1.n4 74.1969
R845 VDD1.n5 VDD1.n3 30.2724
R846 VDD1.n4 VDD1.t1 5.78997
R847 VDD1.n4 VDD1.t7 5.78997
R848 VDD1.n0 VDD1.t2 5.78997
R849 VDD1.n0 VDD1.t0 5.78997
R850 VDD1.n2 VDD1.t4 5.78997
R851 VDD1.n2 VDD1.t3 5.78997
R852 VDD1.n1 VDD1.t5 5.78997
R853 VDD1.n1 VDD1.t6 5.78997
R854 VDD1 VDD1.n5 0.278517
C0 VN VDD1 0.152873f
C1 VDD2 VDD1 0.704224f
C2 VP VDD1 1.62495f
C3 VN VTAIL 1.5571f
C4 VDD2 VTAIL 5.2678f
C5 VP VTAIL 1.5712f
C6 VTAIL VDD1 5.2278f
C7 VN VDD2 1.48221f
C8 VN VP 3.44862f
C9 VDD2 VP 0.296344f
C10 VDD2 B 2.474351f
C11 VDD1 B 2.671213f
C12 VTAIL B 3.761444f
C13 VN B 5.860798f
C14 VP B 4.951251f
C15 VDD1.t2 B 0.058337f
C16 VDD1.t0 B 0.058337f
C17 VDD1.n0 B 0.447754f
C18 VDD1.t5 B 0.058337f
C19 VDD1.t6 B 0.058337f
C20 VDD1.n1 B 0.447355f
C21 VDD1.t4 B 0.058337f
C22 VDD1.t3 B 0.058337f
C23 VDD1.n2 B 0.447355f
C24 VDD1.n3 B 1.33183f
C25 VDD1.t1 B 0.058337f
C26 VDD1.t7 B 0.058337f
C27 VDD1.n4 B 0.446448f
C28 VDD1.n5 B 1.32064f
C29 VP.n0 B 0.027116f
C30 VP.t1 B 0.124133f
C31 VP.n1 B 0.073999f
C32 VP.n2 B 0.027116f
C33 VP.t0 B 0.124133f
C34 VP.t6 B 0.124133f
C35 VP.t7 B 0.124133f
C36 VP.n3 B 0.073999f
C37 VP.t5 B 0.129265f
C38 VP.n4 B 0.066305f
C39 VP.n5 B 0.086f
C40 VP.n6 B 0.006153f
C41 VP.n7 B 0.073999f
C42 VP.n8 B 0.07124f
C43 VP.n9 B 0.779296f
C44 VP.t2 B 0.124133f
C45 VP.n10 B 0.07124f
C46 VP.n11 B 0.807749f
C47 VP.n12 B 0.027116f
C48 VP.n13 B 0.027116f
C49 VP.n14 B 0.006153f
C50 VP.t3 B 0.124133f
C51 VP.n15 B 0.073999f
C52 VP.t4 B 0.124133f
C53 VP.n16 B 0.07124f
C54 VP.n17 B 0.021014f
C55 VTAIL.t9 B 0.052057f
C56 VTAIL.t10 B 0.052057f
C57 VTAIL.n0 B 0.357124f
C58 VTAIL.n1 B 0.20638f
C59 VTAIL.t8 B 0.458214f
C60 VTAIL.n2 B 0.272811f
C61 VTAIL.t3 B 0.458214f
C62 VTAIL.n3 B 0.272811f
C63 VTAIL.t4 B 0.052057f
C64 VTAIL.t15 B 0.052057f
C65 VTAIL.n4 B 0.357124f
C66 VTAIL.n5 B 0.244502f
C67 VTAIL.t1 B 0.458214f
C68 VTAIL.n6 B 0.730021f
C69 VTAIL.t13 B 0.458217f
C70 VTAIL.n7 B 0.730017f
C71 VTAIL.t7 B 0.052057f
C72 VTAIL.t14 B 0.052057f
C73 VTAIL.n8 B 0.357126f
C74 VTAIL.n9 B 0.2445f
C75 VTAIL.t11 B 0.458217f
C76 VTAIL.n10 B 0.272808f
C77 VTAIL.t0 B 0.458217f
C78 VTAIL.n11 B 0.272808f
C79 VTAIL.t6 B 0.052057f
C80 VTAIL.t5 B 0.052057f
C81 VTAIL.n12 B 0.357126f
C82 VTAIL.n13 B 0.2445f
C83 VTAIL.t2 B 0.458214f
C84 VTAIL.n14 B 0.730021f
C85 VTAIL.t12 B 0.458214f
C86 VTAIL.n15 B 0.726409f
C87 VDD2.t2 B 0.060385f
C88 VDD2.t6 B 0.060385f
C89 VDD2.n0 B 0.463058f
C90 VDD2.t4 B 0.060385f
C91 VDD2.t5 B 0.060385f
C92 VDD2.n1 B 0.463058f
C93 VDD2.n2 B 1.33049f
C94 VDD2.t7 B 0.060385f
C95 VDD2.t1 B 0.060385f
C96 VDD2.n3 B 0.462121f
C97 VDD2.n4 B 1.34093f
C98 VDD2.t3 B 0.060385f
C99 VDD2.t0 B 0.060385f
C100 VDD2.n5 B 0.46304f
C101 VN.n0 B 0.026816f
C102 VN.t5 B 0.122757f
C103 VN.n1 B 0.073179f
C104 VN.t6 B 0.127832f
C105 VN.n2 B 0.06557f
C106 VN.n3 B 0.085047f
C107 VN.n4 B 0.006085f
C108 VN.t4 B 0.122757f
C109 VN.n5 B 0.073179f
C110 VN.t2 B 0.122757f
C111 VN.n6 B 0.070451f
C112 VN.n7 B 0.020781f
C113 VN.n8 B 0.026816f
C114 VN.t0 B 0.122757f
C115 VN.n9 B 0.073179f
C116 VN.t3 B 0.127832f
C117 VN.n10 B 0.06557f
C118 VN.n11 B 0.085047f
C119 VN.n12 B 0.006085f
C120 VN.t7 B 0.122757f
C121 VN.n13 B 0.073179f
C122 VN.t1 B 0.122757f
C123 VN.n14 B 0.070451f
C124 VN.n15 B 0.788505f
.ends

