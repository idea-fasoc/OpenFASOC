* NGSPICE file created from diff_pair_sample_1291.ext - technology: sky130A

.subckt diff_pair_sample_1291 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VN.t0 VDD2.t7 w_n5240_n3990# sky130_fd_pr__pfet_01v8 ad=2.49315 pd=15.44 as=2.49315 ps=15.44 w=15.11 l=3.94
X1 B.t11 B.t9 B.t10 w_n5240_n3990# sky130_fd_pr__pfet_01v8 ad=5.8929 pd=31 as=0 ps=0 w=15.11 l=3.94
X2 B.t8 B.t6 B.t7 w_n5240_n3990# sky130_fd_pr__pfet_01v8 ad=5.8929 pd=31 as=0 ps=0 w=15.11 l=3.94
X3 B.t5 B.t3 B.t4 w_n5240_n3990# sky130_fd_pr__pfet_01v8 ad=5.8929 pd=31 as=0 ps=0 w=15.11 l=3.94
X4 VDD1.t7 VP.t0 VTAIL.t2 w_n5240_n3990# sky130_fd_pr__pfet_01v8 ad=2.49315 pd=15.44 as=2.49315 ps=15.44 w=15.11 l=3.94
X5 VTAIL.t14 VN.t1 VDD2.t6 w_n5240_n3990# sky130_fd_pr__pfet_01v8 ad=5.8929 pd=31 as=2.49315 ps=15.44 w=15.11 l=3.94
X6 VTAIL.t1 VP.t1 VDD1.t6 w_n5240_n3990# sky130_fd_pr__pfet_01v8 ad=5.8929 pd=31 as=2.49315 ps=15.44 w=15.11 l=3.94
X7 VDD2.t5 VN.t2 VTAIL.t13 w_n5240_n3990# sky130_fd_pr__pfet_01v8 ad=2.49315 pd=15.44 as=5.8929 ps=31 w=15.11 l=3.94
X8 VTAIL.t12 VN.t3 VDD2.t4 w_n5240_n3990# sky130_fd_pr__pfet_01v8 ad=2.49315 pd=15.44 as=2.49315 ps=15.44 w=15.11 l=3.94
X9 VDD2.t1 VN.t4 VTAIL.t11 w_n5240_n3990# sky130_fd_pr__pfet_01v8 ad=2.49315 pd=15.44 as=5.8929 ps=31 w=15.11 l=3.94
X10 B.t2 B.t0 B.t1 w_n5240_n3990# sky130_fd_pr__pfet_01v8 ad=5.8929 pd=31 as=0 ps=0 w=15.11 l=3.94
X11 VTAIL.t5 VP.t2 VDD1.t5 w_n5240_n3990# sky130_fd_pr__pfet_01v8 ad=2.49315 pd=15.44 as=2.49315 ps=15.44 w=15.11 l=3.94
X12 VDD1.t4 VP.t3 VTAIL.t0 w_n5240_n3990# sky130_fd_pr__pfet_01v8 ad=2.49315 pd=15.44 as=5.8929 ps=31 w=15.11 l=3.94
X13 VDD1.t3 VP.t4 VTAIL.t6 w_n5240_n3990# sky130_fd_pr__pfet_01v8 ad=2.49315 pd=15.44 as=5.8929 ps=31 w=15.11 l=3.94
X14 VDD1.t2 VP.t5 VTAIL.t4 w_n5240_n3990# sky130_fd_pr__pfet_01v8 ad=2.49315 pd=15.44 as=2.49315 ps=15.44 w=15.11 l=3.94
X15 VDD2.t0 VN.t5 VTAIL.t10 w_n5240_n3990# sky130_fd_pr__pfet_01v8 ad=2.49315 pd=15.44 as=2.49315 ps=15.44 w=15.11 l=3.94
X16 VTAIL.t3 VP.t6 VDD1.t1 w_n5240_n3990# sky130_fd_pr__pfet_01v8 ad=2.49315 pd=15.44 as=2.49315 ps=15.44 w=15.11 l=3.94
X17 VTAIL.t7 VP.t7 VDD1.t0 w_n5240_n3990# sky130_fd_pr__pfet_01v8 ad=5.8929 pd=31 as=2.49315 ps=15.44 w=15.11 l=3.94
X18 VTAIL.t9 VN.t6 VDD2.t3 w_n5240_n3990# sky130_fd_pr__pfet_01v8 ad=5.8929 pd=31 as=2.49315 ps=15.44 w=15.11 l=3.94
X19 VDD2.t2 VN.t7 VTAIL.t8 w_n5240_n3990# sky130_fd_pr__pfet_01v8 ad=2.49315 pd=15.44 as=2.49315 ps=15.44 w=15.11 l=3.94
R0 VN.n75 VN.n39 161.3
R1 VN.n74 VN.n73 161.3
R2 VN.n72 VN.n40 161.3
R3 VN.n71 VN.n70 161.3
R4 VN.n69 VN.n41 161.3
R5 VN.n68 VN.n67 161.3
R6 VN.n66 VN.n42 161.3
R7 VN.n65 VN.n64 161.3
R8 VN.n62 VN.n43 161.3
R9 VN.n61 VN.n60 161.3
R10 VN.n59 VN.n44 161.3
R11 VN.n58 VN.n57 161.3
R12 VN.n56 VN.n45 161.3
R13 VN.n55 VN.n54 161.3
R14 VN.n53 VN.n46 161.3
R15 VN.n52 VN.n51 161.3
R16 VN.n50 VN.n47 161.3
R17 VN.n36 VN.n0 161.3
R18 VN.n35 VN.n34 161.3
R19 VN.n33 VN.n1 161.3
R20 VN.n32 VN.n31 161.3
R21 VN.n30 VN.n2 161.3
R22 VN.n29 VN.n28 161.3
R23 VN.n27 VN.n3 161.3
R24 VN.n26 VN.n25 161.3
R25 VN.n23 VN.n4 161.3
R26 VN.n22 VN.n21 161.3
R27 VN.n20 VN.n5 161.3
R28 VN.n19 VN.n18 161.3
R29 VN.n17 VN.n6 161.3
R30 VN.n16 VN.n15 161.3
R31 VN.n14 VN.n7 161.3
R32 VN.n13 VN.n12 161.3
R33 VN.n11 VN.n8 161.3
R34 VN.n9 VN.t1 124.704
R35 VN.n48 VN.t2 124.704
R36 VN.n10 VN.t7 92.4246
R37 VN.n24 VN.t0 92.4246
R38 VN.n37 VN.t4 92.4246
R39 VN.n49 VN.t3 92.4246
R40 VN.n63 VN.t5 92.4246
R41 VN.n76 VN.t6 92.4246
R42 VN.n10 VN.n9 68.4464
R43 VN.n49 VN.n48 68.4464
R44 VN.n38 VN.n37 62.3635
R45 VN.n77 VN.n76 62.3635
R46 VN VN.n77 59.7845
R47 VN.n31 VN.n30 56.5193
R48 VN.n70 VN.n69 56.5193
R49 VN.n17 VN.n16 40.4934
R50 VN.n18 VN.n17 40.4934
R51 VN.n56 VN.n55 40.4934
R52 VN.n57 VN.n56 40.4934
R53 VN.n12 VN.n11 24.4675
R54 VN.n12 VN.n7 24.4675
R55 VN.n16 VN.n7 24.4675
R56 VN.n18 VN.n5 24.4675
R57 VN.n22 VN.n5 24.4675
R58 VN.n23 VN.n22 24.4675
R59 VN.n25 VN.n3 24.4675
R60 VN.n29 VN.n3 24.4675
R61 VN.n30 VN.n29 24.4675
R62 VN.n31 VN.n1 24.4675
R63 VN.n35 VN.n1 24.4675
R64 VN.n36 VN.n35 24.4675
R65 VN.n55 VN.n46 24.4675
R66 VN.n51 VN.n46 24.4675
R67 VN.n51 VN.n50 24.4675
R68 VN.n69 VN.n68 24.4675
R69 VN.n68 VN.n42 24.4675
R70 VN.n64 VN.n42 24.4675
R71 VN.n62 VN.n61 24.4675
R72 VN.n61 VN.n44 24.4675
R73 VN.n57 VN.n44 24.4675
R74 VN.n75 VN.n74 24.4675
R75 VN.n74 VN.n40 24.4675
R76 VN.n70 VN.n40 24.4675
R77 VN.n37 VN.n36 19.8188
R78 VN.n76 VN.n75 19.8188
R79 VN.n25 VN.n24 17.8614
R80 VN.n64 VN.n63 17.8614
R81 VN.n11 VN.n10 6.60659
R82 VN.n24 VN.n23 6.60659
R83 VN.n50 VN.n49 6.60659
R84 VN.n63 VN.n62 6.60659
R85 VN.n48 VN.n47 2.70028
R86 VN.n9 VN.n8 2.70028
R87 VN.n77 VN.n39 0.417535
R88 VN.n38 VN.n0 0.417535
R89 VN VN.n38 0.394291
R90 VN.n73 VN.n39 0.189894
R91 VN.n73 VN.n72 0.189894
R92 VN.n72 VN.n71 0.189894
R93 VN.n71 VN.n41 0.189894
R94 VN.n67 VN.n41 0.189894
R95 VN.n67 VN.n66 0.189894
R96 VN.n66 VN.n65 0.189894
R97 VN.n65 VN.n43 0.189894
R98 VN.n60 VN.n43 0.189894
R99 VN.n60 VN.n59 0.189894
R100 VN.n59 VN.n58 0.189894
R101 VN.n58 VN.n45 0.189894
R102 VN.n54 VN.n45 0.189894
R103 VN.n54 VN.n53 0.189894
R104 VN.n53 VN.n52 0.189894
R105 VN.n52 VN.n47 0.189894
R106 VN.n13 VN.n8 0.189894
R107 VN.n14 VN.n13 0.189894
R108 VN.n15 VN.n14 0.189894
R109 VN.n15 VN.n6 0.189894
R110 VN.n19 VN.n6 0.189894
R111 VN.n20 VN.n19 0.189894
R112 VN.n21 VN.n20 0.189894
R113 VN.n21 VN.n4 0.189894
R114 VN.n26 VN.n4 0.189894
R115 VN.n27 VN.n26 0.189894
R116 VN.n28 VN.n27 0.189894
R117 VN.n28 VN.n2 0.189894
R118 VN.n32 VN.n2 0.189894
R119 VN.n33 VN.n32 0.189894
R120 VN.n34 VN.n33 0.189894
R121 VN.n34 VN.n0 0.189894
R122 VDD2.n2 VDD2.n1 74.4234
R123 VDD2.n2 VDD2.n0 74.4234
R124 VDD2 VDD2.n5 74.4206
R125 VDD2.n4 VDD2.n3 72.6385
R126 VDD2.n4 VDD2.n2 53.3058
R127 VDD2.n5 VDD2.t4 2.15172
R128 VDD2.n5 VDD2.t5 2.15172
R129 VDD2.n3 VDD2.t3 2.15172
R130 VDD2.n3 VDD2.t0 2.15172
R131 VDD2.n1 VDD2.t7 2.15172
R132 VDD2.n1 VDD2.t1 2.15172
R133 VDD2.n0 VDD2.t6 2.15172
R134 VDD2.n0 VDD2.t2 2.15172
R135 VDD2 VDD2.n4 1.89921
R136 VTAIL.n11 VTAIL.t7 58.1109
R137 VTAIL.n10 VTAIL.t13 58.1109
R138 VTAIL.n7 VTAIL.t9 58.1109
R139 VTAIL.n15 VTAIL.t11 58.1107
R140 VTAIL.n2 VTAIL.t14 58.1107
R141 VTAIL.n3 VTAIL.t6 58.1107
R142 VTAIL.n6 VTAIL.t1 58.1107
R143 VTAIL.n14 VTAIL.t0 58.1107
R144 VTAIL.n13 VTAIL.n12 55.9597
R145 VTAIL.n9 VTAIL.n8 55.9597
R146 VTAIL.n1 VTAIL.n0 55.9594
R147 VTAIL.n5 VTAIL.n4 55.9594
R148 VTAIL.n15 VTAIL.n14 29.0738
R149 VTAIL.n7 VTAIL.n6 29.0738
R150 VTAIL.n9 VTAIL.n7 3.68153
R151 VTAIL.n10 VTAIL.n9 3.68153
R152 VTAIL.n13 VTAIL.n11 3.68153
R153 VTAIL.n14 VTAIL.n13 3.68153
R154 VTAIL.n6 VTAIL.n5 3.68153
R155 VTAIL.n5 VTAIL.n3 3.68153
R156 VTAIL.n2 VTAIL.n1 3.68153
R157 VTAIL VTAIL.n15 3.62334
R158 VTAIL.n0 VTAIL.t8 2.15172
R159 VTAIL.n0 VTAIL.t15 2.15172
R160 VTAIL.n4 VTAIL.t2 2.15172
R161 VTAIL.n4 VTAIL.t5 2.15172
R162 VTAIL.n12 VTAIL.t4 2.15172
R163 VTAIL.n12 VTAIL.t3 2.15172
R164 VTAIL.n8 VTAIL.t10 2.15172
R165 VTAIL.n8 VTAIL.t12 2.15172
R166 VTAIL.n11 VTAIL.n10 0.470328
R167 VTAIL.n3 VTAIL.n2 0.470328
R168 VTAIL VTAIL.n1 0.0586897
R169 B.n752 B.n751 585
R170 B.n753 B.n96 585
R171 B.n755 B.n754 585
R172 B.n756 B.n95 585
R173 B.n758 B.n757 585
R174 B.n759 B.n94 585
R175 B.n761 B.n760 585
R176 B.n762 B.n93 585
R177 B.n764 B.n763 585
R178 B.n765 B.n92 585
R179 B.n767 B.n766 585
R180 B.n768 B.n91 585
R181 B.n770 B.n769 585
R182 B.n771 B.n90 585
R183 B.n773 B.n772 585
R184 B.n774 B.n89 585
R185 B.n776 B.n775 585
R186 B.n777 B.n88 585
R187 B.n779 B.n778 585
R188 B.n780 B.n87 585
R189 B.n782 B.n781 585
R190 B.n783 B.n86 585
R191 B.n785 B.n784 585
R192 B.n786 B.n85 585
R193 B.n788 B.n787 585
R194 B.n789 B.n84 585
R195 B.n791 B.n790 585
R196 B.n792 B.n83 585
R197 B.n794 B.n793 585
R198 B.n795 B.n82 585
R199 B.n797 B.n796 585
R200 B.n798 B.n81 585
R201 B.n800 B.n799 585
R202 B.n801 B.n80 585
R203 B.n803 B.n802 585
R204 B.n804 B.n79 585
R205 B.n806 B.n805 585
R206 B.n807 B.n78 585
R207 B.n809 B.n808 585
R208 B.n810 B.n77 585
R209 B.n812 B.n811 585
R210 B.n813 B.n76 585
R211 B.n815 B.n814 585
R212 B.n816 B.n75 585
R213 B.n818 B.n817 585
R214 B.n819 B.n74 585
R215 B.n821 B.n820 585
R216 B.n822 B.n73 585
R217 B.n824 B.n823 585
R218 B.n825 B.n72 585
R219 B.n827 B.n826 585
R220 B.n829 B.n69 585
R221 B.n831 B.n830 585
R222 B.n832 B.n68 585
R223 B.n834 B.n833 585
R224 B.n835 B.n67 585
R225 B.n837 B.n836 585
R226 B.n838 B.n66 585
R227 B.n840 B.n839 585
R228 B.n841 B.n63 585
R229 B.n844 B.n843 585
R230 B.n845 B.n62 585
R231 B.n847 B.n846 585
R232 B.n848 B.n61 585
R233 B.n850 B.n849 585
R234 B.n851 B.n60 585
R235 B.n853 B.n852 585
R236 B.n854 B.n59 585
R237 B.n856 B.n855 585
R238 B.n857 B.n58 585
R239 B.n859 B.n858 585
R240 B.n860 B.n57 585
R241 B.n862 B.n861 585
R242 B.n863 B.n56 585
R243 B.n865 B.n864 585
R244 B.n866 B.n55 585
R245 B.n868 B.n867 585
R246 B.n869 B.n54 585
R247 B.n871 B.n870 585
R248 B.n872 B.n53 585
R249 B.n874 B.n873 585
R250 B.n875 B.n52 585
R251 B.n877 B.n876 585
R252 B.n878 B.n51 585
R253 B.n880 B.n879 585
R254 B.n881 B.n50 585
R255 B.n883 B.n882 585
R256 B.n884 B.n49 585
R257 B.n886 B.n885 585
R258 B.n887 B.n48 585
R259 B.n889 B.n888 585
R260 B.n890 B.n47 585
R261 B.n892 B.n891 585
R262 B.n893 B.n46 585
R263 B.n895 B.n894 585
R264 B.n896 B.n45 585
R265 B.n898 B.n897 585
R266 B.n899 B.n44 585
R267 B.n901 B.n900 585
R268 B.n902 B.n43 585
R269 B.n904 B.n903 585
R270 B.n905 B.n42 585
R271 B.n907 B.n906 585
R272 B.n908 B.n41 585
R273 B.n910 B.n909 585
R274 B.n911 B.n40 585
R275 B.n913 B.n912 585
R276 B.n914 B.n39 585
R277 B.n916 B.n915 585
R278 B.n917 B.n38 585
R279 B.n919 B.n918 585
R280 B.n750 B.n97 585
R281 B.n749 B.n748 585
R282 B.n747 B.n98 585
R283 B.n746 B.n745 585
R284 B.n744 B.n99 585
R285 B.n743 B.n742 585
R286 B.n741 B.n100 585
R287 B.n740 B.n739 585
R288 B.n738 B.n101 585
R289 B.n737 B.n736 585
R290 B.n735 B.n102 585
R291 B.n734 B.n733 585
R292 B.n732 B.n103 585
R293 B.n731 B.n730 585
R294 B.n729 B.n104 585
R295 B.n728 B.n727 585
R296 B.n726 B.n105 585
R297 B.n725 B.n724 585
R298 B.n723 B.n106 585
R299 B.n722 B.n721 585
R300 B.n720 B.n107 585
R301 B.n719 B.n718 585
R302 B.n717 B.n108 585
R303 B.n716 B.n715 585
R304 B.n714 B.n109 585
R305 B.n713 B.n712 585
R306 B.n711 B.n110 585
R307 B.n710 B.n709 585
R308 B.n708 B.n111 585
R309 B.n707 B.n706 585
R310 B.n705 B.n112 585
R311 B.n704 B.n703 585
R312 B.n702 B.n113 585
R313 B.n701 B.n700 585
R314 B.n699 B.n114 585
R315 B.n698 B.n697 585
R316 B.n696 B.n115 585
R317 B.n695 B.n694 585
R318 B.n693 B.n116 585
R319 B.n692 B.n691 585
R320 B.n690 B.n117 585
R321 B.n689 B.n688 585
R322 B.n687 B.n118 585
R323 B.n686 B.n685 585
R324 B.n684 B.n119 585
R325 B.n683 B.n682 585
R326 B.n681 B.n120 585
R327 B.n680 B.n679 585
R328 B.n678 B.n121 585
R329 B.n677 B.n676 585
R330 B.n675 B.n122 585
R331 B.n674 B.n673 585
R332 B.n672 B.n123 585
R333 B.n671 B.n670 585
R334 B.n669 B.n124 585
R335 B.n668 B.n667 585
R336 B.n666 B.n125 585
R337 B.n665 B.n664 585
R338 B.n663 B.n126 585
R339 B.n662 B.n661 585
R340 B.n660 B.n127 585
R341 B.n659 B.n658 585
R342 B.n657 B.n128 585
R343 B.n656 B.n655 585
R344 B.n654 B.n129 585
R345 B.n653 B.n652 585
R346 B.n651 B.n130 585
R347 B.n650 B.n649 585
R348 B.n648 B.n131 585
R349 B.n647 B.n646 585
R350 B.n645 B.n132 585
R351 B.n644 B.n643 585
R352 B.n642 B.n133 585
R353 B.n641 B.n640 585
R354 B.n639 B.n134 585
R355 B.n638 B.n637 585
R356 B.n636 B.n135 585
R357 B.n635 B.n634 585
R358 B.n633 B.n136 585
R359 B.n632 B.n631 585
R360 B.n630 B.n137 585
R361 B.n629 B.n628 585
R362 B.n627 B.n138 585
R363 B.n626 B.n625 585
R364 B.n624 B.n139 585
R365 B.n623 B.n622 585
R366 B.n621 B.n140 585
R367 B.n620 B.n619 585
R368 B.n618 B.n141 585
R369 B.n617 B.n616 585
R370 B.n615 B.n142 585
R371 B.n614 B.n613 585
R372 B.n612 B.n143 585
R373 B.n611 B.n610 585
R374 B.n609 B.n144 585
R375 B.n608 B.n607 585
R376 B.n606 B.n145 585
R377 B.n605 B.n604 585
R378 B.n603 B.n146 585
R379 B.n602 B.n601 585
R380 B.n600 B.n147 585
R381 B.n599 B.n598 585
R382 B.n597 B.n148 585
R383 B.n596 B.n595 585
R384 B.n594 B.n149 585
R385 B.n593 B.n592 585
R386 B.n591 B.n150 585
R387 B.n590 B.n589 585
R388 B.n588 B.n151 585
R389 B.n587 B.n586 585
R390 B.n585 B.n152 585
R391 B.n584 B.n583 585
R392 B.n582 B.n153 585
R393 B.n581 B.n580 585
R394 B.n579 B.n154 585
R395 B.n578 B.n577 585
R396 B.n576 B.n155 585
R397 B.n575 B.n574 585
R398 B.n573 B.n156 585
R399 B.n572 B.n571 585
R400 B.n570 B.n157 585
R401 B.n569 B.n568 585
R402 B.n567 B.n158 585
R403 B.n566 B.n565 585
R404 B.n564 B.n159 585
R405 B.n563 B.n562 585
R406 B.n561 B.n160 585
R407 B.n560 B.n559 585
R408 B.n558 B.n161 585
R409 B.n557 B.n556 585
R410 B.n555 B.n162 585
R411 B.n554 B.n553 585
R412 B.n552 B.n163 585
R413 B.n551 B.n550 585
R414 B.n549 B.n164 585
R415 B.n548 B.n547 585
R416 B.n546 B.n165 585
R417 B.n545 B.n544 585
R418 B.n543 B.n166 585
R419 B.n542 B.n541 585
R420 B.n540 B.n167 585
R421 B.n539 B.n538 585
R422 B.n537 B.n168 585
R423 B.n369 B.n228 585
R424 B.n371 B.n370 585
R425 B.n372 B.n227 585
R426 B.n374 B.n373 585
R427 B.n375 B.n226 585
R428 B.n377 B.n376 585
R429 B.n378 B.n225 585
R430 B.n380 B.n379 585
R431 B.n381 B.n224 585
R432 B.n383 B.n382 585
R433 B.n384 B.n223 585
R434 B.n386 B.n385 585
R435 B.n387 B.n222 585
R436 B.n389 B.n388 585
R437 B.n390 B.n221 585
R438 B.n392 B.n391 585
R439 B.n393 B.n220 585
R440 B.n395 B.n394 585
R441 B.n396 B.n219 585
R442 B.n398 B.n397 585
R443 B.n399 B.n218 585
R444 B.n401 B.n400 585
R445 B.n402 B.n217 585
R446 B.n404 B.n403 585
R447 B.n405 B.n216 585
R448 B.n407 B.n406 585
R449 B.n408 B.n215 585
R450 B.n410 B.n409 585
R451 B.n411 B.n214 585
R452 B.n413 B.n412 585
R453 B.n414 B.n213 585
R454 B.n416 B.n415 585
R455 B.n417 B.n212 585
R456 B.n419 B.n418 585
R457 B.n420 B.n211 585
R458 B.n422 B.n421 585
R459 B.n423 B.n210 585
R460 B.n425 B.n424 585
R461 B.n426 B.n209 585
R462 B.n428 B.n427 585
R463 B.n429 B.n208 585
R464 B.n431 B.n430 585
R465 B.n432 B.n207 585
R466 B.n434 B.n433 585
R467 B.n435 B.n206 585
R468 B.n437 B.n436 585
R469 B.n438 B.n205 585
R470 B.n440 B.n439 585
R471 B.n441 B.n204 585
R472 B.n443 B.n442 585
R473 B.n444 B.n201 585
R474 B.n447 B.n446 585
R475 B.n448 B.n200 585
R476 B.n450 B.n449 585
R477 B.n451 B.n199 585
R478 B.n453 B.n452 585
R479 B.n454 B.n198 585
R480 B.n456 B.n455 585
R481 B.n457 B.n197 585
R482 B.n459 B.n458 585
R483 B.n461 B.n460 585
R484 B.n462 B.n193 585
R485 B.n464 B.n463 585
R486 B.n465 B.n192 585
R487 B.n467 B.n466 585
R488 B.n468 B.n191 585
R489 B.n470 B.n469 585
R490 B.n471 B.n190 585
R491 B.n473 B.n472 585
R492 B.n474 B.n189 585
R493 B.n476 B.n475 585
R494 B.n477 B.n188 585
R495 B.n479 B.n478 585
R496 B.n480 B.n187 585
R497 B.n482 B.n481 585
R498 B.n483 B.n186 585
R499 B.n485 B.n484 585
R500 B.n486 B.n185 585
R501 B.n488 B.n487 585
R502 B.n489 B.n184 585
R503 B.n491 B.n490 585
R504 B.n492 B.n183 585
R505 B.n494 B.n493 585
R506 B.n495 B.n182 585
R507 B.n497 B.n496 585
R508 B.n498 B.n181 585
R509 B.n500 B.n499 585
R510 B.n501 B.n180 585
R511 B.n503 B.n502 585
R512 B.n504 B.n179 585
R513 B.n506 B.n505 585
R514 B.n507 B.n178 585
R515 B.n509 B.n508 585
R516 B.n510 B.n177 585
R517 B.n512 B.n511 585
R518 B.n513 B.n176 585
R519 B.n515 B.n514 585
R520 B.n516 B.n175 585
R521 B.n518 B.n517 585
R522 B.n519 B.n174 585
R523 B.n521 B.n520 585
R524 B.n522 B.n173 585
R525 B.n524 B.n523 585
R526 B.n525 B.n172 585
R527 B.n527 B.n526 585
R528 B.n528 B.n171 585
R529 B.n530 B.n529 585
R530 B.n531 B.n170 585
R531 B.n533 B.n532 585
R532 B.n534 B.n169 585
R533 B.n536 B.n535 585
R534 B.n368 B.n367 585
R535 B.n366 B.n229 585
R536 B.n365 B.n364 585
R537 B.n363 B.n230 585
R538 B.n362 B.n361 585
R539 B.n360 B.n231 585
R540 B.n359 B.n358 585
R541 B.n357 B.n232 585
R542 B.n356 B.n355 585
R543 B.n354 B.n233 585
R544 B.n353 B.n352 585
R545 B.n351 B.n234 585
R546 B.n350 B.n349 585
R547 B.n348 B.n235 585
R548 B.n347 B.n346 585
R549 B.n345 B.n236 585
R550 B.n344 B.n343 585
R551 B.n342 B.n237 585
R552 B.n341 B.n340 585
R553 B.n339 B.n238 585
R554 B.n338 B.n337 585
R555 B.n336 B.n239 585
R556 B.n335 B.n334 585
R557 B.n333 B.n240 585
R558 B.n332 B.n331 585
R559 B.n330 B.n241 585
R560 B.n329 B.n328 585
R561 B.n327 B.n242 585
R562 B.n326 B.n325 585
R563 B.n324 B.n243 585
R564 B.n323 B.n322 585
R565 B.n321 B.n244 585
R566 B.n320 B.n319 585
R567 B.n318 B.n245 585
R568 B.n317 B.n316 585
R569 B.n315 B.n246 585
R570 B.n314 B.n313 585
R571 B.n312 B.n247 585
R572 B.n311 B.n310 585
R573 B.n309 B.n248 585
R574 B.n308 B.n307 585
R575 B.n306 B.n249 585
R576 B.n305 B.n304 585
R577 B.n303 B.n250 585
R578 B.n302 B.n301 585
R579 B.n300 B.n251 585
R580 B.n299 B.n298 585
R581 B.n297 B.n252 585
R582 B.n296 B.n295 585
R583 B.n294 B.n253 585
R584 B.n293 B.n292 585
R585 B.n291 B.n254 585
R586 B.n290 B.n289 585
R587 B.n288 B.n255 585
R588 B.n287 B.n286 585
R589 B.n285 B.n256 585
R590 B.n284 B.n283 585
R591 B.n282 B.n257 585
R592 B.n281 B.n280 585
R593 B.n279 B.n258 585
R594 B.n278 B.n277 585
R595 B.n276 B.n259 585
R596 B.n275 B.n274 585
R597 B.n273 B.n260 585
R598 B.n272 B.n271 585
R599 B.n270 B.n261 585
R600 B.n269 B.n268 585
R601 B.n267 B.n262 585
R602 B.n266 B.n265 585
R603 B.n264 B.n263 585
R604 B.n2 B.n0 585
R605 B.n1025 B.n1 585
R606 B.n1024 B.n1023 585
R607 B.n1022 B.n3 585
R608 B.n1021 B.n1020 585
R609 B.n1019 B.n4 585
R610 B.n1018 B.n1017 585
R611 B.n1016 B.n5 585
R612 B.n1015 B.n1014 585
R613 B.n1013 B.n6 585
R614 B.n1012 B.n1011 585
R615 B.n1010 B.n7 585
R616 B.n1009 B.n1008 585
R617 B.n1007 B.n8 585
R618 B.n1006 B.n1005 585
R619 B.n1004 B.n9 585
R620 B.n1003 B.n1002 585
R621 B.n1001 B.n10 585
R622 B.n1000 B.n999 585
R623 B.n998 B.n11 585
R624 B.n997 B.n996 585
R625 B.n995 B.n12 585
R626 B.n994 B.n993 585
R627 B.n992 B.n13 585
R628 B.n991 B.n990 585
R629 B.n989 B.n14 585
R630 B.n988 B.n987 585
R631 B.n986 B.n15 585
R632 B.n985 B.n984 585
R633 B.n983 B.n16 585
R634 B.n982 B.n981 585
R635 B.n980 B.n17 585
R636 B.n979 B.n978 585
R637 B.n977 B.n18 585
R638 B.n976 B.n975 585
R639 B.n974 B.n19 585
R640 B.n973 B.n972 585
R641 B.n971 B.n20 585
R642 B.n970 B.n969 585
R643 B.n968 B.n21 585
R644 B.n967 B.n966 585
R645 B.n965 B.n22 585
R646 B.n964 B.n963 585
R647 B.n962 B.n23 585
R648 B.n961 B.n960 585
R649 B.n959 B.n24 585
R650 B.n958 B.n957 585
R651 B.n956 B.n25 585
R652 B.n955 B.n954 585
R653 B.n953 B.n26 585
R654 B.n952 B.n951 585
R655 B.n950 B.n27 585
R656 B.n949 B.n948 585
R657 B.n947 B.n28 585
R658 B.n946 B.n945 585
R659 B.n944 B.n29 585
R660 B.n943 B.n942 585
R661 B.n941 B.n30 585
R662 B.n940 B.n939 585
R663 B.n938 B.n31 585
R664 B.n937 B.n936 585
R665 B.n935 B.n32 585
R666 B.n934 B.n933 585
R667 B.n932 B.n33 585
R668 B.n931 B.n930 585
R669 B.n929 B.n34 585
R670 B.n928 B.n927 585
R671 B.n926 B.n35 585
R672 B.n925 B.n924 585
R673 B.n923 B.n36 585
R674 B.n922 B.n921 585
R675 B.n920 B.n37 585
R676 B.n1027 B.n1026 585
R677 B.n369 B.n368 492.5
R678 B.n918 B.n37 492.5
R679 B.n537 B.n536 492.5
R680 B.n752 B.n97 492.5
R681 B.n194 B.t9 301.873
R682 B.n202 B.t3 301.873
R683 B.n64 B.t6 301.873
R684 B.n70 B.t0 301.873
R685 B.n194 B.t11 192.267
R686 B.n70 B.t1 192.267
R687 B.n202 B.t5 192.248
R688 B.n64 B.t7 192.248
R689 B.n368 B.n229 163.367
R690 B.n364 B.n229 163.367
R691 B.n364 B.n363 163.367
R692 B.n363 B.n362 163.367
R693 B.n362 B.n231 163.367
R694 B.n358 B.n231 163.367
R695 B.n358 B.n357 163.367
R696 B.n357 B.n356 163.367
R697 B.n356 B.n233 163.367
R698 B.n352 B.n233 163.367
R699 B.n352 B.n351 163.367
R700 B.n351 B.n350 163.367
R701 B.n350 B.n235 163.367
R702 B.n346 B.n235 163.367
R703 B.n346 B.n345 163.367
R704 B.n345 B.n344 163.367
R705 B.n344 B.n237 163.367
R706 B.n340 B.n237 163.367
R707 B.n340 B.n339 163.367
R708 B.n339 B.n338 163.367
R709 B.n338 B.n239 163.367
R710 B.n334 B.n239 163.367
R711 B.n334 B.n333 163.367
R712 B.n333 B.n332 163.367
R713 B.n332 B.n241 163.367
R714 B.n328 B.n241 163.367
R715 B.n328 B.n327 163.367
R716 B.n327 B.n326 163.367
R717 B.n326 B.n243 163.367
R718 B.n322 B.n243 163.367
R719 B.n322 B.n321 163.367
R720 B.n321 B.n320 163.367
R721 B.n320 B.n245 163.367
R722 B.n316 B.n245 163.367
R723 B.n316 B.n315 163.367
R724 B.n315 B.n314 163.367
R725 B.n314 B.n247 163.367
R726 B.n310 B.n247 163.367
R727 B.n310 B.n309 163.367
R728 B.n309 B.n308 163.367
R729 B.n308 B.n249 163.367
R730 B.n304 B.n249 163.367
R731 B.n304 B.n303 163.367
R732 B.n303 B.n302 163.367
R733 B.n302 B.n251 163.367
R734 B.n298 B.n251 163.367
R735 B.n298 B.n297 163.367
R736 B.n297 B.n296 163.367
R737 B.n296 B.n253 163.367
R738 B.n292 B.n253 163.367
R739 B.n292 B.n291 163.367
R740 B.n291 B.n290 163.367
R741 B.n290 B.n255 163.367
R742 B.n286 B.n255 163.367
R743 B.n286 B.n285 163.367
R744 B.n285 B.n284 163.367
R745 B.n284 B.n257 163.367
R746 B.n280 B.n257 163.367
R747 B.n280 B.n279 163.367
R748 B.n279 B.n278 163.367
R749 B.n278 B.n259 163.367
R750 B.n274 B.n259 163.367
R751 B.n274 B.n273 163.367
R752 B.n273 B.n272 163.367
R753 B.n272 B.n261 163.367
R754 B.n268 B.n261 163.367
R755 B.n268 B.n267 163.367
R756 B.n267 B.n266 163.367
R757 B.n266 B.n263 163.367
R758 B.n263 B.n2 163.367
R759 B.n1026 B.n2 163.367
R760 B.n1026 B.n1025 163.367
R761 B.n1025 B.n1024 163.367
R762 B.n1024 B.n3 163.367
R763 B.n1020 B.n3 163.367
R764 B.n1020 B.n1019 163.367
R765 B.n1019 B.n1018 163.367
R766 B.n1018 B.n5 163.367
R767 B.n1014 B.n5 163.367
R768 B.n1014 B.n1013 163.367
R769 B.n1013 B.n1012 163.367
R770 B.n1012 B.n7 163.367
R771 B.n1008 B.n7 163.367
R772 B.n1008 B.n1007 163.367
R773 B.n1007 B.n1006 163.367
R774 B.n1006 B.n9 163.367
R775 B.n1002 B.n9 163.367
R776 B.n1002 B.n1001 163.367
R777 B.n1001 B.n1000 163.367
R778 B.n1000 B.n11 163.367
R779 B.n996 B.n11 163.367
R780 B.n996 B.n995 163.367
R781 B.n995 B.n994 163.367
R782 B.n994 B.n13 163.367
R783 B.n990 B.n13 163.367
R784 B.n990 B.n989 163.367
R785 B.n989 B.n988 163.367
R786 B.n988 B.n15 163.367
R787 B.n984 B.n15 163.367
R788 B.n984 B.n983 163.367
R789 B.n983 B.n982 163.367
R790 B.n982 B.n17 163.367
R791 B.n978 B.n17 163.367
R792 B.n978 B.n977 163.367
R793 B.n977 B.n976 163.367
R794 B.n976 B.n19 163.367
R795 B.n972 B.n19 163.367
R796 B.n972 B.n971 163.367
R797 B.n971 B.n970 163.367
R798 B.n970 B.n21 163.367
R799 B.n966 B.n21 163.367
R800 B.n966 B.n965 163.367
R801 B.n965 B.n964 163.367
R802 B.n964 B.n23 163.367
R803 B.n960 B.n23 163.367
R804 B.n960 B.n959 163.367
R805 B.n959 B.n958 163.367
R806 B.n958 B.n25 163.367
R807 B.n954 B.n25 163.367
R808 B.n954 B.n953 163.367
R809 B.n953 B.n952 163.367
R810 B.n952 B.n27 163.367
R811 B.n948 B.n27 163.367
R812 B.n948 B.n947 163.367
R813 B.n947 B.n946 163.367
R814 B.n946 B.n29 163.367
R815 B.n942 B.n29 163.367
R816 B.n942 B.n941 163.367
R817 B.n941 B.n940 163.367
R818 B.n940 B.n31 163.367
R819 B.n936 B.n31 163.367
R820 B.n936 B.n935 163.367
R821 B.n935 B.n934 163.367
R822 B.n934 B.n33 163.367
R823 B.n930 B.n33 163.367
R824 B.n930 B.n929 163.367
R825 B.n929 B.n928 163.367
R826 B.n928 B.n35 163.367
R827 B.n924 B.n35 163.367
R828 B.n924 B.n923 163.367
R829 B.n923 B.n922 163.367
R830 B.n922 B.n37 163.367
R831 B.n370 B.n369 163.367
R832 B.n370 B.n227 163.367
R833 B.n374 B.n227 163.367
R834 B.n375 B.n374 163.367
R835 B.n376 B.n375 163.367
R836 B.n376 B.n225 163.367
R837 B.n380 B.n225 163.367
R838 B.n381 B.n380 163.367
R839 B.n382 B.n381 163.367
R840 B.n382 B.n223 163.367
R841 B.n386 B.n223 163.367
R842 B.n387 B.n386 163.367
R843 B.n388 B.n387 163.367
R844 B.n388 B.n221 163.367
R845 B.n392 B.n221 163.367
R846 B.n393 B.n392 163.367
R847 B.n394 B.n393 163.367
R848 B.n394 B.n219 163.367
R849 B.n398 B.n219 163.367
R850 B.n399 B.n398 163.367
R851 B.n400 B.n399 163.367
R852 B.n400 B.n217 163.367
R853 B.n404 B.n217 163.367
R854 B.n405 B.n404 163.367
R855 B.n406 B.n405 163.367
R856 B.n406 B.n215 163.367
R857 B.n410 B.n215 163.367
R858 B.n411 B.n410 163.367
R859 B.n412 B.n411 163.367
R860 B.n412 B.n213 163.367
R861 B.n416 B.n213 163.367
R862 B.n417 B.n416 163.367
R863 B.n418 B.n417 163.367
R864 B.n418 B.n211 163.367
R865 B.n422 B.n211 163.367
R866 B.n423 B.n422 163.367
R867 B.n424 B.n423 163.367
R868 B.n424 B.n209 163.367
R869 B.n428 B.n209 163.367
R870 B.n429 B.n428 163.367
R871 B.n430 B.n429 163.367
R872 B.n430 B.n207 163.367
R873 B.n434 B.n207 163.367
R874 B.n435 B.n434 163.367
R875 B.n436 B.n435 163.367
R876 B.n436 B.n205 163.367
R877 B.n440 B.n205 163.367
R878 B.n441 B.n440 163.367
R879 B.n442 B.n441 163.367
R880 B.n442 B.n201 163.367
R881 B.n447 B.n201 163.367
R882 B.n448 B.n447 163.367
R883 B.n449 B.n448 163.367
R884 B.n449 B.n199 163.367
R885 B.n453 B.n199 163.367
R886 B.n454 B.n453 163.367
R887 B.n455 B.n454 163.367
R888 B.n455 B.n197 163.367
R889 B.n459 B.n197 163.367
R890 B.n460 B.n459 163.367
R891 B.n460 B.n193 163.367
R892 B.n464 B.n193 163.367
R893 B.n465 B.n464 163.367
R894 B.n466 B.n465 163.367
R895 B.n466 B.n191 163.367
R896 B.n470 B.n191 163.367
R897 B.n471 B.n470 163.367
R898 B.n472 B.n471 163.367
R899 B.n472 B.n189 163.367
R900 B.n476 B.n189 163.367
R901 B.n477 B.n476 163.367
R902 B.n478 B.n477 163.367
R903 B.n478 B.n187 163.367
R904 B.n482 B.n187 163.367
R905 B.n483 B.n482 163.367
R906 B.n484 B.n483 163.367
R907 B.n484 B.n185 163.367
R908 B.n488 B.n185 163.367
R909 B.n489 B.n488 163.367
R910 B.n490 B.n489 163.367
R911 B.n490 B.n183 163.367
R912 B.n494 B.n183 163.367
R913 B.n495 B.n494 163.367
R914 B.n496 B.n495 163.367
R915 B.n496 B.n181 163.367
R916 B.n500 B.n181 163.367
R917 B.n501 B.n500 163.367
R918 B.n502 B.n501 163.367
R919 B.n502 B.n179 163.367
R920 B.n506 B.n179 163.367
R921 B.n507 B.n506 163.367
R922 B.n508 B.n507 163.367
R923 B.n508 B.n177 163.367
R924 B.n512 B.n177 163.367
R925 B.n513 B.n512 163.367
R926 B.n514 B.n513 163.367
R927 B.n514 B.n175 163.367
R928 B.n518 B.n175 163.367
R929 B.n519 B.n518 163.367
R930 B.n520 B.n519 163.367
R931 B.n520 B.n173 163.367
R932 B.n524 B.n173 163.367
R933 B.n525 B.n524 163.367
R934 B.n526 B.n525 163.367
R935 B.n526 B.n171 163.367
R936 B.n530 B.n171 163.367
R937 B.n531 B.n530 163.367
R938 B.n532 B.n531 163.367
R939 B.n532 B.n169 163.367
R940 B.n536 B.n169 163.367
R941 B.n538 B.n537 163.367
R942 B.n538 B.n167 163.367
R943 B.n542 B.n167 163.367
R944 B.n543 B.n542 163.367
R945 B.n544 B.n543 163.367
R946 B.n544 B.n165 163.367
R947 B.n548 B.n165 163.367
R948 B.n549 B.n548 163.367
R949 B.n550 B.n549 163.367
R950 B.n550 B.n163 163.367
R951 B.n554 B.n163 163.367
R952 B.n555 B.n554 163.367
R953 B.n556 B.n555 163.367
R954 B.n556 B.n161 163.367
R955 B.n560 B.n161 163.367
R956 B.n561 B.n560 163.367
R957 B.n562 B.n561 163.367
R958 B.n562 B.n159 163.367
R959 B.n566 B.n159 163.367
R960 B.n567 B.n566 163.367
R961 B.n568 B.n567 163.367
R962 B.n568 B.n157 163.367
R963 B.n572 B.n157 163.367
R964 B.n573 B.n572 163.367
R965 B.n574 B.n573 163.367
R966 B.n574 B.n155 163.367
R967 B.n578 B.n155 163.367
R968 B.n579 B.n578 163.367
R969 B.n580 B.n579 163.367
R970 B.n580 B.n153 163.367
R971 B.n584 B.n153 163.367
R972 B.n585 B.n584 163.367
R973 B.n586 B.n585 163.367
R974 B.n586 B.n151 163.367
R975 B.n590 B.n151 163.367
R976 B.n591 B.n590 163.367
R977 B.n592 B.n591 163.367
R978 B.n592 B.n149 163.367
R979 B.n596 B.n149 163.367
R980 B.n597 B.n596 163.367
R981 B.n598 B.n597 163.367
R982 B.n598 B.n147 163.367
R983 B.n602 B.n147 163.367
R984 B.n603 B.n602 163.367
R985 B.n604 B.n603 163.367
R986 B.n604 B.n145 163.367
R987 B.n608 B.n145 163.367
R988 B.n609 B.n608 163.367
R989 B.n610 B.n609 163.367
R990 B.n610 B.n143 163.367
R991 B.n614 B.n143 163.367
R992 B.n615 B.n614 163.367
R993 B.n616 B.n615 163.367
R994 B.n616 B.n141 163.367
R995 B.n620 B.n141 163.367
R996 B.n621 B.n620 163.367
R997 B.n622 B.n621 163.367
R998 B.n622 B.n139 163.367
R999 B.n626 B.n139 163.367
R1000 B.n627 B.n626 163.367
R1001 B.n628 B.n627 163.367
R1002 B.n628 B.n137 163.367
R1003 B.n632 B.n137 163.367
R1004 B.n633 B.n632 163.367
R1005 B.n634 B.n633 163.367
R1006 B.n634 B.n135 163.367
R1007 B.n638 B.n135 163.367
R1008 B.n639 B.n638 163.367
R1009 B.n640 B.n639 163.367
R1010 B.n640 B.n133 163.367
R1011 B.n644 B.n133 163.367
R1012 B.n645 B.n644 163.367
R1013 B.n646 B.n645 163.367
R1014 B.n646 B.n131 163.367
R1015 B.n650 B.n131 163.367
R1016 B.n651 B.n650 163.367
R1017 B.n652 B.n651 163.367
R1018 B.n652 B.n129 163.367
R1019 B.n656 B.n129 163.367
R1020 B.n657 B.n656 163.367
R1021 B.n658 B.n657 163.367
R1022 B.n658 B.n127 163.367
R1023 B.n662 B.n127 163.367
R1024 B.n663 B.n662 163.367
R1025 B.n664 B.n663 163.367
R1026 B.n664 B.n125 163.367
R1027 B.n668 B.n125 163.367
R1028 B.n669 B.n668 163.367
R1029 B.n670 B.n669 163.367
R1030 B.n670 B.n123 163.367
R1031 B.n674 B.n123 163.367
R1032 B.n675 B.n674 163.367
R1033 B.n676 B.n675 163.367
R1034 B.n676 B.n121 163.367
R1035 B.n680 B.n121 163.367
R1036 B.n681 B.n680 163.367
R1037 B.n682 B.n681 163.367
R1038 B.n682 B.n119 163.367
R1039 B.n686 B.n119 163.367
R1040 B.n687 B.n686 163.367
R1041 B.n688 B.n687 163.367
R1042 B.n688 B.n117 163.367
R1043 B.n692 B.n117 163.367
R1044 B.n693 B.n692 163.367
R1045 B.n694 B.n693 163.367
R1046 B.n694 B.n115 163.367
R1047 B.n698 B.n115 163.367
R1048 B.n699 B.n698 163.367
R1049 B.n700 B.n699 163.367
R1050 B.n700 B.n113 163.367
R1051 B.n704 B.n113 163.367
R1052 B.n705 B.n704 163.367
R1053 B.n706 B.n705 163.367
R1054 B.n706 B.n111 163.367
R1055 B.n710 B.n111 163.367
R1056 B.n711 B.n710 163.367
R1057 B.n712 B.n711 163.367
R1058 B.n712 B.n109 163.367
R1059 B.n716 B.n109 163.367
R1060 B.n717 B.n716 163.367
R1061 B.n718 B.n717 163.367
R1062 B.n718 B.n107 163.367
R1063 B.n722 B.n107 163.367
R1064 B.n723 B.n722 163.367
R1065 B.n724 B.n723 163.367
R1066 B.n724 B.n105 163.367
R1067 B.n728 B.n105 163.367
R1068 B.n729 B.n728 163.367
R1069 B.n730 B.n729 163.367
R1070 B.n730 B.n103 163.367
R1071 B.n734 B.n103 163.367
R1072 B.n735 B.n734 163.367
R1073 B.n736 B.n735 163.367
R1074 B.n736 B.n101 163.367
R1075 B.n740 B.n101 163.367
R1076 B.n741 B.n740 163.367
R1077 B.n742 B.n741 163.367
R1078 B.n742 B.n99 163.367
R1079 B.n746 B.n99 163.367
R1080 B.n747 B.n746 163.367
R1081 B.n748 B.n747 163.367
R1082 B.n748 B.n97 163.367
R1083 B.n918 B.n917 163.367
R1084 B.n917 B.n916 163.367
R1085 B.n916 B.n39 163.367
R1086 B.n912 B.n39 163.367
R1087 B.n912 B.n911 163.367
R1088 B.n911 B.n910 163.367
R1089 B.n910 B.n41 163.367
R1090 B.n906 B.n41 163.367
R1091 B.n906 B.n905 163.367
R1092 B.n905 B.n904 163.367
R1093 B.n904 B.n43 163.367
R1094 B.n900 B.n43 163.367
R1095 B.n900 B.n899 163.367
R1096 B.n899 B.n898 163.367
R1097 B.n898 B.n45 163.367
R1098 B.n894 B.n45 163.367
R1099 B.n894 B.n893 163.367
R1100 B.n893 B.n892 163.367
R1101 B.n892 B.n47 163.367
R1102 B.n888 B.n47 163.367
R1103 B.n888 B.n887 163.367
R1104 B.n887 B.n886 163.367
R1105 B.n886 B.n49 163.367
R1106 B.n882 B.n49 163.367
R1107 B.n882 B.n881 163.367
R1108 B.n881 B.n880 163.367
R1109 B.n880 B.n51 163.367
R1110 B.n876 B.n51 163.367
R1111 B.n876 B.n875 163.367
R1112 B.n875 B.n874 163.367
R1113 B.n874 B.n53 163.367
R1114 B.n870 B.n53 163.367
R1115 B.n870 B.n869 163.367
R1116 B.n869 B.n868 163.367
R1117 B.n868 B.n55 163.367
R1118 B.n864 B.n55 163.367
R1119 B.n864 B.n863 163.367
R1120 B.n863 B.n862 163.367
R1121 B.n862 B.n57 163.367
R1122 B.n858 B.n57 163.367
R1123 B.n858 B.n857 163.367
R1124 B.n857 B.n856 163.367
R1125 B.n856 B.n59 163.367
R1126 B.n852 B.n59 163.367
R1127 B.n852 B.n851 163.367
R1128 B.n851 B.n850 163.367
R1129 B.n850 B.n61 163.367
R1130 B.n846 B.n61 163.367
R1131 B.n846 B.n845 163.367
R1132 B.n845 B.n844 163.367
R1133 B.n844 B.n63 163.367
R1134 B.n839 B.n63 163.367
R1135 B.n839 B.n838 163.367
R1136 B.n838 B.n837 163.367
R1137 B.n837 B.n67 163.367
R1138 B.n833 B.n67 163.367
R1139 B.n833 B.n832 163.367
R1140 B.n832 B.n831 163.367
R1141 B.n831 B.n69 163.367
R1142 B.n826 B.n69 163.367
R1143 B.n826 B.n825 163.367
R1144 B.n825 B.n824 163.367
R1145 B.n824 B.n73 163.367
R1146 B.n820 B.n73 163.367
R1147 B.n820 B.n819 163.367
R1148 B.n819 B.n818 163.367
R1149 B.n818 B.n75 163.367
R1150 B.n814 B.n75 163.367
R1151 B.n814 B.n813 163.367
R1152 B.n813 B.n812 163.367
R1153 B.n812 B.n77 163.367
R1154 B.n808 B.n77 163.367
R1155 B.n808 B.n807 163.367
R1156 B.n807 B.n806 163.367
R1157 B.n806 B.n79 163.367
R1158 B.n802 B.n79 163.367
R1159 B.n802 B.n801 163.367
R1160 B.n801 B.n800 163.367
R1161 B.n800 B.n81 163.367
R1162 B.n796 B.n81 163.367
R1163 B.n796 B.n795 163.367
R1164 B.n795 B.n794 163.367
R1165 B.n794 B.n83 163.367
R1166 B.n790 B.n83 163.367
R1167 B.n790 B.n789 163.367
R1168 B.n789 B.n788 163.367
R1169 B.n788 B.n85 163.367
R1170 B.n784 B.n85 163.367
R1171 B.n784 B.n783 163.367
R1172 B.n783 B.n782 163.367
R1173 B.n782 B.n87 163.367
R1174 B.n778 B.n87 163.367
R1175 B.n778 B.n777 163.367
R1176 B.n777 B.n776 163.367
R1177 B.n776 B.n89 163.367
R1178 B.n772 B.n89 163.367
R1179 B.n772 B.n771 163.367
R1180 B.n771 B.n770 163.367
R1181 B.n770 B.n91 163.367
R1182 B.n766 B.n91 163.367
R1183 B.n766 B.n765 163.367
R1184 B.n765 B.n764 163.367
R1185 B.n764 B.n93 163.367
R1186 B.n760 B.n93 163.367
R1187 B.n760 B.n759 163.367
R1188 B.n759 B.n758 163.367
R1189 B.n758 B.n95 163.367
R1190 B.n754 B.n95 163.367
R1191 B.n754 B.n753 163.367
R1192 B.n753 B.n752 163.367
R1193 B.n195 B.t10 109.454
R1194 B.n71 B.t2 109.454
R1195 B.n203 B.t4 109.436
R1196 B.n65 B.t8 109.436
R1197 B.n195 B.n194 82.8126
R1198 B.n203 B.n202 82.8126
R1199 B.n65 B.n64 82.8126
R1200 B.n71 B.n70 82.8126
R1201 B.n196 B.n195 59.5399
R1202 B.n445 B.n203 59.5399
R1203 B.n842 B.n65 59.5399
R1204 B.n828 B.n71 59.5399
R1205 B.n920 B.n919 32.0005
R1206 B.n751 B.n750 32.0005
R1207 B.n535 B.n168 32.0005
R1208 B.n367 B.n228 32.0005
R1209 B B.n1027 18.0485
R1210 B.n919 B.n38 10.6151
R1211 B.n915 B.n38 10.6151
R1212 B.n915 B.n914 10.6151
R1213 B.n914 B.n913 10.6151
R1214 B.n913 B.n40 10.6151
R1215 B.n909 B.n40 10.6151
R1216 B.n909 B.n908 10.6151
R1217 B.n908 B.n907 10.6151
R1218 B.n907 B.n42 10.6151
R1219 B.n903 B.n42 10.6151
R1220 B.n903 B.n902 10.6151
R1221 B.n902 B.n901 10.6151
R1222 B.n901 B.n44 10.6151
R1223 B.n897 B.n44 10.6151
R1224 B.n897 B.n896 10.6151
R1225 B.n896 B.n895 10.6151
R1226 B.n895 B.n46 10.6151
R1227 B.n891 B.n46 10.6151
R1228 B.n891 B.n890 10.6151
R1229 B.n890 B.n889 10.6151
R1230 B.n889 B.n48 10.6151
R1231 B.n885 B.n48 10.6151
R1232 B.n885 B.n884 10.6151
R1233 B.n884 B.n883 10.6151
R1234 B.n883 B.n50 10.6151
R1235 B.n879 B.n50 10.6151
R1236 B.n879 B.n878 10.6151
R1237 B.n878 B.n877 10.6151
R1238 B.n877 B.n52 10.6151
R1239 B.n873 B.n52 10.6151
R1240 B.n873 B.n872 10.6151
R1241 B.n872 B.n871 10.6151
R1242 B.n871 B.n54 10.6151
R1243 B.n867 B.n54 10.6151
R1244 B.n867 B.n866 10.6151
R1245 B.n866 B.n865 10.6151
R1246 B.n865 B.n56 10.6151
R1247 B.n861 B.n56 10.6151
R1248 B.n861 B.n860 10.6151
R1249 B.n860 B.n859 10.6151
R1250 B.n859 B.n58 10.6151
R1251 B.n855 B.n58 10.6151
R1252 B.n855 B.n854 10.6151
R1253 B.n854 B.n853 10.6151
R1254 B.n853 B.n60 10.6151
R1255 B.n849 B.n60 10.6151
R1256 B.n849 B.n848 10.6151
R1257 B.n848 B.n847 10.6151
R1258 B.n847 B.n62 10.6151
R1259 B.n843 B.n62 10.6151
R1260 B.n841 B.n840 10.6151
R1261 B.n840 B.n66 10.6151
R1262 B.n836 B.n66 10.6151
R1263 B.n836 B.n835 10.6151
R1264 B.n835 B.n834 10.6151
R1265 B.n834 B.n68 10.6151
R1266 B.n830 B.n68 10.6151
R1267 B.n830 B.n829 10.6151
R1268 B.n827 B.n72 10.6151
R1269 B.n823 B.n72 10.6151
R1270 B.n823 B.n822 10.6151
R1271 B.n822 B.n821 10.6151
R1272 B.n821 B.n74 10.6151
R1273 B.n817 B.n74 10.6151
R1274 B.n817 B.n816 10.6151
R1275 B.n816 B.n815 10.6151
R1276 B.n815 B.n76 10.6151
R1277 B.n811 B.n76 10.6151
R1278 B.n811 B.n810 10.6151
R1279 B.n810 B.n809 10.6151
R1280 B.n809 B.n78 10.6151
R1281 B.n805 B.n78 10.6151
R1282 B.n805 B.n804 10.6151
R1283 B.n804 B.n803 10.6151
R1284 B.n803 B.n80 10.6151
R1285 B.n799 B.n80 10.6151
R1286 B.n799 B.n798 10.6151
R1287 B.n798 B.n797 10.6151
R1288 B.n797 B.n82 10.6151
R1289 B.n793 B.n82 10.6151
R1290 B.n793 B.n792 10.6151
R1291 B.n792 B.n791 10.6151
R1292 B.n791 B.n84 10.6151
R1293 B.n787 B.n84 10.6151
R1294 B.n787 B.n786 10.6151
R1295 B.n786 B.n785 10.6151
R1296 B.n785 B.n86 10.6151
R1297 B.n781 B.n86 10.6151
R1298 B.n781 B.n780 10.6151
R1299 B.n780 B.n779 10.6151
R1300 B.n779 B.n88 10.6151
R1301 B.n775 B.n88 10.6151
R1302 B.n775 B.n774 10.6151
R1303 B.n774 B.n773 10.6151
R1304 B.n773 B.n90 10.6151
R1305 B.n769 B.n90 10.6151
R1306 B.n769 B.n768 10.6151
R1307 B.n768 B.n767 10.6151
R1308 B.n767 B.n92 10.6151
R1309 B.n763 B.n92 10.6151
R1310 B.n763 B.n762 10.6151
R1311 B.n762 B.n761 10.6151
R1312 B.n761 B.n94 10.6151
R1313 B.n757 B.n94 10.6151
R1314 B.n757 B.n756 10.6151
R1315 B.n756 B.n755 10.6151
R1316 B.n755 B.n96 10.6151
R1317 B.n751 B.n96 10.6151
R1318 B.n539 B.n168 10.6151
R1319 B.n540 B.n539 10.6151
R1320 B.n541 B.n540 10.6151
R1321 B.n541 B.n166 10.6151
R1322 B.n545 B.n166 10.6151
R1323 B.n546 B.n545 10.6151
R1324 B.n547 B.n546 10.6151
R1325 B.n547 B.n164 10.6151
R1326 B.n551 B.n164 10.6151
R1327 B.n552 B.n551 10.6151
R1328 B.n553 B.n552 10.6151
R1329 B.n553 B.n162 10.6151
R1330 B.n557 B.n162 10.6151
R1331 B.n558 B.n557 10.6151
R1332 B.n559 B.n558 10.6151
R1333 B.n559 B.n160 10.6151
R1334 B.n563 B.n160 10.6151
R1335 B.n564 B.n563 10.6151
R1336 B.n565 B.n564 10.6151
R1337 B.n565 B.n158 10.6151
R1338 B.n569 B.n158 10.6151
R1339 B.n570 B.n569 10.6151
R1340 B.n571 B.n570 10.6151
R1341 B.n571 B.n156 10.6151
R1342 B.n575 B.n156 10.6151
R1343 B.n576 B.n575 10.6151
R1344 B.n577 B.n576 10.6151
R1345 B.n577 B.n154 10.6151
R1346 B.n581 B.n154 10.6151
R1347 B.n582 B.n581 10.6151
R1348 B.n583 B.n582 10.6151
R1349 B.n583 B.n152 10.6151
R1350 B.n587 B.n152 10.6151
R1351 B.n588 B.n587 10.6151
R1352 B.n589 B.n588 10.6151
R1353 B.n589 B.n150 10.6151
R1354 B.n593 B.n150 10.6151
R1355 B.n594 B.n593 10.6151
R1356 B.n595 B.n594 10.6151
R1357 B.n595 B.n148 10.6151
R1358 B.n599 B.n148 10.6151
R1359 B.n600 B.n599 10.6151
R1360 B.n601 B.n600 10.6151
R1361 B.n601 B.n146 10.6151
R1362 B.n605 B.n146 10.6151
R1363 B.n606 B.n605 10.6151
R1364 B.n607 B.n606 10.6151
R1365 B.n607 B.n144 10.6151
R1366 B.n611 B.n144 10.6151
R1367 B.n612 B.n611 10.6151
R1368 B.n613 B.n612 10.6151
R1369 B.n613 B.n142 10.6151
R1370 B.n617 B.n142 10.6151
R1371 B.n618 B.n617 10.6151
R1372 B.n619 B.n618 10.6151
R1373 B.n619 B.n140 10.6151
R1374 B.n623 B.n140 10.6151
R1375 B.n624 B.n623 10.6151
R1376 B.n625 B.n624 10.6151
R1377 B.n625 B.n138 10.6151
R1378 B.n629 B.n138 10.6151
R1379 B.n630 B.n629 10.6151
R1380 B.n631 B.n630 10.6151
R1381 B.n631 B.n136 10.6151
R1382 B.n635 B.n136 10.6151
R1383 B.n636 B.n635 10.6151
R1384 B.n637 B.n636 10.6151
R1385 B.n637 B.n134 10.6151
R1386 B.n641 B.n134 10.6151
R1387 B.n642 B.n641 10.6151
R1388 B.n643 B.n642 10.6151
R1389 B.n643 B.n132 10.6151
R1390 B.n647 B.n132 10.6151
R1391 B.n648 B.n647 10.6151
R1392 B.n649 B.n648 10.6151
R1393 B.n649 B.n130 10.6151
R1394 B.n653 B.n130 10.6151
R1395 B.n654 B.n653 10.6151
R1396 B.n655 B.n654 10.6151
R1397 B.n655 B.n128 10.6151
R1398 B.n659 B.n128 10.6151
R1399 B.n660 B.n659 10.6151
R1400 B.n661 B.n660 10.6151
R1401 B.n661 B.n126 10.6151
R1402 B.n665 B.n126 10.6151
R1403 B.n666 B.n665 10.6151
R1404 B.n667 B.n666 10.6151
R1405 B.n667 B.n124 10.6151
R1406 B.n671 B.n124 10.6151
R1407 B.n672 B.n671 10.6151
R1408 B.n673 B.n672 10.6151
R1409 B.n673 B.n122 10.6151
R1410 B.n677 B.n122 10.6151
R1411 B.n678 B.n677 10.6151
R1412 B.n679 B.n678 10.6151
R1413 B.n679 B.n120 10.6151
R1414 B.n683 B.n120 10.6151
R1415 B.n684 B.n683 10.6151
R1416 B.n685 B.n684 10.6151
R1417 B.n685 B.n118 10.6151
R1418 B.n689 B.n118 10.6151
R1419 B.n690 B.n689 10.6151
R1420 B.n691 B.n690 10.6151
R1421 B.n691 B.n116 10.6151
R1422 B.n695 B.n116 10.6151
R1423 B.n696 B.n695 10.6151
R1424 B.n697 B.n696 10.6151
R1425 B.n697 B.n114 10.6151
R1426 B.n701 B.n114 10.6151
R1427 B.n702 B.n701 10.6151
R1428 B.n703 B.n702 10.6151
R1429 B.n703 B.n112 10.6151
R1430 B.n707 B.n112 10.6151
R1431 B.n708 B.n707 10.6151
R1432 B.n709 B.n708 10.6151
R1433 B.n709 B.n110 10.6151
R1434 B.n713 B.n110 10.6151
R1435 B.n714 B.n713 10.6151
R1436 B.n715 B.n714 10.6151
R1437 B.n715 B.n108 10.6151
R1438 B.n719 B.n108 10.6151
R1439 B.n720 B.n719 10.6151
R1440 B.n721 B.n720 10.6151
R1441 B.n721 B.n106 10.6151
R1442 B.n725 B.n106 10.6151
R1443 B.n726 B.n725 10.6151
R1444 B.n727 B.n726 10.6151
R1445 B.n727 B.n104 10.6151
R1446 B.n731 B.n104 10.6151
R1447 B.n732 B.n731 10.6151
R1448 B.n733 B.n732 10.6151
R1449 B.n733 B.n102 10.6151
R1450 B.n737 B.n102 10.6151
R1451 B.n738 B.n737 10.6151
R1452 B.n739 B.n738 10.6151
R1453 B.n739 B.n100 10.6151
R1454 B.n743 B.n100 10.6151
R1455 B.n744 B.n743 10.6151
R1456 B.n745 B.n744 10.6151
R1457 B.n745 B.n98 10.6151
R1458 B.n749 B.n98 10.6151
R1459 B.n750 B.n749 10.6151
R1460 B.n371 B.n228 10.6151
R1461 B.n372 B.n371 10.6151
R1462 B.n373 B.n372 10.6151
R1463 B.n373 B.n226 10.6151
R1464 B.n377 B.n226 10.6151
R1465 B.n378 B.n377 10.6151
R1466 B.n379 B.n378 10.6151
R1467 B.n379 B.n224 10.6151
R1468 B.n383 B.n224 10.6151
R1469 B.n384 B.n383 10.6151
R1470 B.n385 B.n384 10.6151
R1471 B.n385 B.n222 10.6151
R1472 B.n389 B.n222 10.6151
R1473 B.n390 B.n389 10.6151
R1474 B.n391 B.n390 10.6151
R1475 B.n391 B.n220 10.6151
R1476 B.n395 B.n220 10.6151
R1477 B.n396 B.n395 10.6151
R1478 B.n397 B.n396 10.6151
R1479 B.n397 B.n218 10.6151
R1480 B.n401 B.n218 10.6151
R1481 B.n402 B.n401 10.6151
R1482 B.n403 B.n402 10.6151
R1483 B.n403 B.n216 10.6151
R1484 B.n407 B.n216 10.6151
R1485 B.n408 B.n407 10.6151
R1486 B.n409 B.n408 10.6151
R1487 B.n409 B.n214 10.6151
R1488 B.n413 B.n214 10.6151
R1489 B.n414 B.n413 10.6151
R1490 B.n415 B.n414 10.6151
R1491 B.n415 B.n212 10.6151
R1492 B.n419 B.n212 10.6151
R1493 B.n420 B.n419 10.6151
R1494 B.n421 B.n420 10.6151
R1495 B.n421 B.n210 10.6151
R1496 B.n425 B.n210 10.6151
R1497 B.n426 B.n425 10.6151
R1498 B.n427 B.n426 10.6151
R1499 B.n427 B.n208 10.6151
R1500 B.n431 B.n208 10.6151
R1501 B.n432 B.n431 10.6151
R1502 B.n433 B.n432 10.6151
R1503 B.n433 B.n206 10.6151
R1504 B.n437 B.n206 10.6151
R1505 B.n438 B.n437 10.6151
R1506 B.n439 B.n438 10.6151
R1507 B.n439 B.n204 10.6151
R1508 B.n443 B.n204 10.6151
R1509 B.n444 B.n443 10.6151
R1510 B.n446 B.n200 10.6151
R1511 B.n450 B.n200 10.6151
R1512 B.n451 B.n450 10.6151
R1513 B.n452 B.n451 10.6151
R1514 B.n452 B.n198 10.6151
R1515 B.n456 B.n198 10.6151
R1516 B.n457 B.n456 10.6151
R1517 B.n458 B.n457 10.6151
R1518 B.n462 B.n461 10.6151
R1519 B.n463 B.n462 10.6151
R1520 B.n463 B.n192 10.6151
R1521 B.n467 B.n192 10.6151
R1522 B.n468 B.n467 10.6151
R1523 B.n469 B.n468 10.6151
R1524 B.n469 B.n190 10.6151
R1525 B.n473 B.n190 10.6151
R1526 B.n474 B.n473 10.6151
R1527 B.n475 B.n474 10.6151
R1528 B.n475 B.n188 10.6151
R1529 B.n479 B.n188 10.6151
R1530 B.n480 B.n479 10.6151
R1531 B.n481 B.n480 10.6151
R1532 B.n481 B.n186 10.6151
R1533 B.n485 B.n186 10.6151
R1534 B.n486 B.n485 10.6151
R1535 B.n487 B.n486 10.6151
R1536 B.n487 B.n184 10.6151
R1537 B.n491 B.n184 10.6151
R1538 B.n492 B.n491 10.6151
R1539 B.n493 B.n492 10.6151
R1540 B.n493 B.n182 10.6151
R1541 B.n497 B.n182 10.6151
R1542 B.n498 B.n497 10.6151
R1543 B.n499 B.n498 10.6151
R1544 B.n499 B.n180 10.6151
R1545 B.n503 B.n180 10.6151
R1546 B.n504 B.n503 10.6151
R1547 B.n505 B.n504 10.6151
R1548 B.n505 B.n178 10.6151
R1549 B.n509 B.n178 10.6151
R1550 B.n510 B.n509 10.6151
R1551 B.n511 B.n510 10.6151
R1552 B.n511 B.n176 10.6151
R1553 B.n515 B.n176 10.6151
R1554 B.n516 B.n515 10.6151
R1555 B.n517 B.n516 10.6151
R1556 B.n517 B.n174 10.6151
R1557 B.n521 B.n174 10.6151
R1558 B.n522 B.n521 10.6151
R1559 B.n523 B.n522 10.6151
R1560 B.n523 B.n172 10.6151
R1561 B.n527 B.n172 10.6151
R1562 B.n528 B.n527 10.6151
R1563 B.n529 B.n528 10.6151
R1564 B.n529 B.n170 10.6151
R1565 B.n533 B.n170 10.6151
R1566 B.n534 B.n533 10.6151
R1567 B.n535 B.n534 10.6151
R1568 B.n367 B.n366 10.6151
R1569 B.n366 B.n365 10.6151
R1570 B.n365 B.n230 10.6151
R1571 B.n361 B.n230 10.6151
R1572 B.n361 B.n360 10.6151
R1573 B.n360 B.n359 10.6151
R1574 B.n359 B.n232 10.6151
R1575 B.n355 B.n232 10.6151
R1576 B.n355 B.n354 10.6151
R1577 B.n354 B.n353 10.6151
R1578 B.n353 B.n234 10.6151
R1579 B.n349 B.n234 10.6151
R1580 B.n349 B.n348 10.6151
R1581 B.n348 B.n347 10.6151
R1582 B.n347 B.n236 10.6151
R1583 B.n343 B.n236 10.6151
R1584 B.n343 B.n342 10.6151
R1585 B.n342 B.n341 10.6151
R1586 B.n341 B.n238 10.6151
R1587 B.n337 B.n238 10.6151
R1588 B.n337 B.n336 10.6151
R1589 B.n336 B.n335 10.6151
R1590 B.n335 B.n240 10.6151
R1591 B.n331 B.n240 10.6151
R1592 B.n331 B.n330 10.6151
R1593 B.n330 B.n329 10.6151
R1594 B.n329 B.n242 10.6151
R1595 B.n325 B.n242 10.6151
R1596 B.n325 B.n324 10.6151
R1597 B.n324 B.n323 10.6151
R1598 B.n323 B.n244 10.6151
R1599 B.n319 B.n244 10.6151
R1600 B.n319 B.n318 10.6151
R1601 B.n318 B.n317 10.6151
R1602 B.n317 B.n246 10.6151
R1603 B.n313 B.n246 10.6151
R1604 B.n313 B.n312 10.6151
R1605 B.n312 B.n311 10.6151
R1606 B.n311 B.n248 10.6151
R1607 B.n307 B.n248 10.6151
R1608 B.n307 B.n306 10.6151
R1609 B.n306 B.n305 10.6151
R1610 B.n305 B.n250 10.6151
R1611 B.n301 B.n250 10.6151
R1612 B.n301 B.n300 10.6151
R1613 B.n300 B.n299 10.6151
R1614 B.n299 B.n252 10.6151
R1615 B.n295 B.n252 10.6151
R1616 B.n295 B.n294 10.6151
R1617 B.n294 B.n293 10.6151
R1618 B.n293 B.n254 10.6151
R1619 B.n289 B.n254 10.6151
R1620 B.n289 B.n288 10.6151
R1621 B.n288 B.n287 10.6151
R1622 B.n287 B.n256 10.6151
R1623 B.n283 B.n256 10.6151
R1624 B.n283 B.n282 10.6151
R1625 B.n282 B.n281 10.6151
R1626 B.n281 B.n258 10.6151
R1627 B.n277 B.n258 10.6151
R1628 B.n277 B.n276 10.6151
R1629 B.n276 B.n275 10.6151
R1630 B.n275 B.n260 10.6151
R1631 B.n271 B.n260 10.6151
R1632 B.n271 B.n270 10.6151
R1633 B.n270 B.n269 10.6151
R1634 B.n269 B.n262 10.6151
R1635 B.n265 B.n262 10.6151
R1636 B.n265 B.n264 10.6151
R1637 B.n264 B.n0 10.6151
R1638 B.n1023 B.n1 10.6151
R1639 B.n1023 B.n1022 10.6151
R1640 B.n1022 B.n1021 10.6151
R1641 B.n1021 B.n4 10.6151
R1642 B.n1017 B.n4 10.6151
R1643 B.n1017 B.n1016 10.6151
R1644 B.n1016 B.n1015 10.6151
R1645 B.n1015 B.n6 10.6151
R1646 B.n1011 B.n6 10.6151
R1647 B.n1011 B.n1010 10.6151
R1648 B.n1010 B.n1009 10.6151
R1649 B.n1009 B.n8 10.6151
R1650 B.n1005 B.n8 10.6151
R1651 B.n1005 B.n1004 10.6151
R1652 B.n1004 B.n1003 10.6151
R1653 B.n1003 B.n10 10.6151
R1654 B.n999 B.n10 10.6151
R1655 B.n999 B.n998 10.6151
R1656 B.n998 B.n997 10.6151
R1657 B.n997 B.n12 10.6151
R1658 B.n993 B.n12 10.6151
R1659 B.n993 B.n992 10.6151
R1660 B.n992 B.n991 10.6151
R1661 B.n991 B.n14 10.6151
R1662 B.n987 B.n14 10.6151
R1663 B.n987 B.n986 10.6151
R1664 B.n986 B.n985 10.6151
R1665 B.n985 B.n16 10.6151
R1666 B.n981 B.n16 10.6151
R1667 B.n981 B.n980 10.6151
R1668 B.n980 B.n979 10.6151
R1669 B.n979 B.n18 10.6151
R1670 B.n975 B.n18 10.6151
R1671 B.n975 B.n974 10.6151
R1672 B.n974 B.n973 10.6151
R1673 B.n973 B.n20 10.6151
R1674 B.n969 B.n20 10.6151
R1675 B.n969 B.n968 10.6151
R1676 B.n968 B.n967 10.6151
R1677 B.n967 B.n22 10.6151
R1678 B.n963 B.n22 10.6151
R1679 B.n963 B.n962 10.6151
R1680 B.n962 B.n961 10.6151
R1681 B.n961 B.n24 10.6151
R1682 B.n957 B.n24 10.6151
R1683 B.n957 B.n956 10.6151
R1684 B.n956 B.n955 10.6151
R1685 B.n955 B.n26 10.6151
R1686 B.n951 B.n26 10.6151
R1687 B.n951 B.n950 10.6151
R1688 B.n950 B.n949 10.6151
R1689 B.n949 B.n28 10.6151
R1690 B.n945 B.n28 10.6151
R1691 B.n945 B.n944 10.6151
R1692 B.n944 B.n943 10.6151
R1693 B.n943 B.n30 10.6151
R1694 B.n939 B.n30 10.6151
R1695 B.n939 B.n938 10.6151
R1696 B.n938 B.n937 10.6151
R1697 B.n937 B.n32 10.6151
R1698 B.n933 B.n32 10.6151
R1699 B.n933 B.n932 10.6151
R1700 B.n932 B.n931 10.6151
R1701 B.n931 B.n34 10.6151
R1702 B.n927 B.n34 10.6151
R1703 B.n927 B.n926 10.6151
R1704 B.n926 B.n925 10.6151
R1705 B.n925 B.n36 10.6151
R1706 B.n921 B.n36 10.6151
R1707 B.n921 B.n920 10.6151
R1708 B.n842 B.n841 6.5566
R1709 B.n829 B.n828 6.5566
R1710 B.n446 B.n445 6.5566
R1711 B.n458 B.n196 6.5566
R1712 B.n843 B.n842 4.05904
R1713 B.n828 B.n827 4.05904
R1714 B.n445 B.n444 4.05904
R1715 B.n461 B.n196 4.05904
R1716 B.n1027 B.n0 2.81026
R1717 B.n1027 B.n1 2.81026
R1718 VP.n24 VP.n21 161.3
R1719 VP.n26 VP.n25 161.3
R1720 VP.n27 VP.n20 161.3
R1721 VP.n29 VP.n28 161.3
R1722 VP.n30 VP.n19 161.3
R1723 VP.n32 VP.n31 161.3
R1724 VP.n33 VP.n18 161.3
R1725 VP.n35 VP.n34 161.3
R1726 VP.n36 VP.n17 161.3
R1727 VP.n39 VP.n38 161.3
R1728 VP.n40 VP.n16 161.3
R1729 VP.n42 VP.n41 161.3
R1730 VP.n43 VP.n15 161.3
R1731 VP.n45 VP.n44 161.3
R1732 VP.n46 VP.n14 161.3
R1733 VP.n48 VP.n47 161.3
R1734 VP.n49 VP.n13 161.3
R1735 VP.n92 VP.n0 161.3
R1736 VP.n91 VP.n90 161.3
R1737 VP.n89 VP.n1 161.3
R1738 VP.n88 VP.n87 161.3
R1739 VP.n86 VP.n2 161.3
R1740 VP.n85 VP.n84 161.3
R1741 VP.n83 VP.n3 161.3
R1742 VP.n82 VP.n81 161.3
R1743 VP.n79 VP.n4 161.3
R1744 VP.n78 VP.n77 161.3
R1745 VP.n76 VP.n5 161.3
R1746 VP.n75 VP.n74 161.3
R1747 VP.n73 VP.n6 161.3
R1748 VP.n72 VP.n71 161.3
R1749 VP.n70 VP.n7 161.3
R1750 VP.n69 VP.n68 161.3
R1751 VP.n67 VP.n8 161.3
R1752 VP.n65 VP.n64 161.3
R1753 VP.n63 VP.n9 161.3
R1754 VP.n62 VP.n61 161.3
R1755 VP.n60 VP.n10 161.3
R1756 VP.n59 VP.n58 161.3
R1757 VP.n57 VP.n11 161.3
R1758 VP.n56 VP.n55 161.3
R1759 VP.n54 VP.n12 161.3
R1760 VP.n22 VP.t7 124.704
R1761 VP.n53 VP.t1 92.4246
R1762 VP.n66 VP.t0 92.4246
R1763 VP.n80 VP.t2 92.4246
R1764 VP.n93 VP.t4 92.4246
R1765 VP.n50 VP.t3 92.4246
R1766 VP.n37 VP.t6 92.4246
R1767 VP.n23 VP.t5 92.4246
R1768 VP.n23 VP.n22 68.4464
R1769 VP.n53 VP.n52 62.3635
R1770 VP.n94 VP.n93 62.3635
R1771 VP.n51 VP.n50 62.3635
R1772 VP.n52 VP.n51 59.7464
R1773 VP.n60 VP.n59 56.5193
R1774 VP.n87 VP.n86 56.5193
R1775 VP.n44 VP.n43 56.5193
R1776 VP.n73 VP.n72 40.4934
R1777 VP.n74 VP.n73 40.4934
R1778 VP.n31 VP.n30 40.4934
R1779 VP.n30 VP.n29 40.4934
R1780 VP.n55 VP.n54 24.4675
R1781 VP.n55 VP.n11 24.4675
R1782 VP.n59 VP.n11 24.4675
R1783 VP.n61 VP.n60 24.4675
R1784 VP.n61 VP.n9 24.4675
R1785 VP.n65 VP.n9 24.4675
R1786 VP.n68 VP.n67 24.4675
R1787 VP.n68 VP.n7 24.4675
R1788 VP.n72 VP.n7 24.4675
R1789 VP.n74 VP.n5 24.4675
R1790 VP.n78 VP.n5 24.4675
R1791 VP.n79 VP.n78 24.4675
R1792 VP.n81 VP.n3 24.4675
R1793 VP.n85 VP.n3 24.4675
R1794 VP.n86 VP.n85 24.4675
R1795 VP.n87 VP.n1 24.4675
R1796 VP.n91 VP.n1 24.4675
R1797 VP.n92 VP.n91 24.4675
R1798 VP.n44 VP.n14 24.4675
R1799 VP.n48 VP.n14 24.4675
R1800 VP.n49 VP.n48 24.4675
R1801 VP.n31 VP.n18 24.4675
R1802 VP.n35 VP.n18 24.4675
R1803 VP.n36 VP.n35 24.4675
R1804 VP.n38 VP.n16 24.4675
R1805 VP.n42 VP.n16 24.4675
R1806 VP.n43 VP.n42 24.4675
R1807 VP.n25 VP.n24 24.4675
R1808 VP.n25 VP.n20 24.4675
R1809 VP.n29 VP.n20 24.4675
R1810 VP.n54 VP.n53 19.8188
R1811 VP.n93 VP.n92 19.8188
R1812 VP.n50 VP.n49 19.8188
R1813 VP.n66 VP.n65 17.8614
R1814 VP.n81 VP.n80 17.8614
R1815 VP.n38 VP.n37 17.8614
R1816 VP.n67 VP.n66 6.60659
R1817 VP.n80 VP.n79 6.60659
R1818 VP.n37 VP.n36 6.60659
R1819 VP.n24 VP.n23 6.60659
R1820 VP.n22 VP.n21 2.70025
R1821 VP.n51 VP.n13 0.417535
R1822 VP.n52 VP.n12 0.417535
R1823 VP.n94 VP.n0 0.417535
R1824 VP VP.n94 0.394291
R1825 VP.n26 VP.n21 0.189894
R1826 VP.n27 VP.n26 0.189894
R1827 VP.n28 VP.n27 0.189894
R1828 VP.n28 VP.n19 0.189894
R1829 VP.n32 VP.n19 0.189894
R1830 VP.n33 VP.n32 0.189894
R1831 VP.n34 VP.n33 0.189894
R1832 VP.n34 VP.n17 0.189894
R1833 VP.n39 VP.n17 0.189894
R1834 VP.n40 VP.n39 0.189894
R1835 VP.n41 VP.n40 0.189894
R1836 VP.n41 VP.n15 0.189894
R1837 VP.n45 VP.n15 0.189894
R1838 VP.n46 VP.n45 0.189894
R1839 VP.n47 VP.n46 0.189894
R1840 VP.n47 VP.n13 0.189894
R1841 VP.n56 VP.n12 0.189894
R1842 VP.n57 VP.n56 0.189894
R1843 VP.n58 VP.n57 0.189894
R1844 VP.n58 VP.n10 0.189894
R1845 VP.n62 VP.n10 0.189894
R1846 VP.n63 VP.n62 0.189894
R1847 VP.n64 VP.n63 0.189894
R1848 VP.n64 VP.n8 0.189894
R1849 VP.n69 VP.n8 0.189894
R1850 VP.n70 VP.n69 0.189894
R1851 VP.n71 VP.n70 0.189894
R1852 VP.n71 VP.n6 0.189894
R1853 VP.n75 VP.n6 0.189894
R1854 VP.n76 VP.n75 0.189894
R1855 VP.n77 VP.n76 0.189894
R1856 VP.n77 VP.n4 0.189894
R1857 VP.n82 VP.n4 0.189894
R1858 VP.n83 VP.n82 0.189894
R1859 VP.n84 VP.n83 0.189894
R1860 VP.n84 VP.n2 0.189894
R1861 VP.n88 VP.n2 0.189894
R1862 VP.n89 VP.n88 0.189894
R1863 VP.n90 VP.n89 0.189894
R1864 VP.n90 VP.n0 0.189894
R1865 VDD1 VDD1.n0 74.5372
R1866 VDD1.n3 VDD1.n2 74.4234
R1867 VDD1.n3 VDD1.n1 74.4234
R1868 VDD1.n5 VDD1.n4 72.6383
R1869 VDD1.n5 VDD1.n3 53.8888
R1870 VDD1.n4 VDD1.t1 2.15172
R1871 VDD1.n4 VDD1.t4 2.15172
R1872 VDD1.n0 VDD1.t0 2.15172
R1873 VDD1.n0 VDD1.t2 2.15172
R1874 VDD1.n2 VDD1.t5 2.15172
R1875 VDD1.n2 VDD1.t3 2.15172
R1876 VDD1.n1 VDD1.t6 2.15172
R1877 VDD1.n1 VDD1.t7 2.15172
R1878 VDD1 VDD1.n5 1.78283
C0 VDD1 VDD2 2.4744f
C1 B w_n5240_n3990# 13.0383f
C2 VP w_n5240_n3990# 11.7877f
C3 B VN 1.57361f
C4 VP VN 9.881289f
C5 VTAIL B 6.60662f
C6 VTAIL VP 12.3046f
C7 B VDD2 2.28088f
C8 VP VDD2 0.662414f
C9 VN w_n5240_n3990# 11.1035f
C10 VTAIL w_n5240_n3990# 4.99055f
C11 VDD2 w_n5240_n3990# 2.64122f
C12 VDD1 B 2.1427f
C13 VDD1 VP 12.0925f
C14 VTAIL VN 12.2905f
C15 VN VDD2 11.5864f
C16 VTAIL VDD2 9.604401f
C17 VDD1 w_n5240_n3990# 2.4703f
C18 VDD1 VN 0.154303f
C19 B VP 2.72773f
C20 VDD1 VTAIL 9.541f
C21 VDD2 VSUBS 2.60176f
C22 VDD1 VSUBS 3.478f
C23 VTAIL VSUBS 1.725632f
C24 VN VSUBS 8.649639f
C25 VP VSUBS 5.086952f
C26 B VSUBS 6.759576f
C27 w_n5240_n3990# VSUBS 0.256362p
C28 VDD1.t0 VSUBS 0.386584f
C29 VDD1.t2 VSUBS 0.386584f
C30 VDD1.n0 VSUBS 3.18077f
C31 VDD1.t6 VSUBS 0.386584f
C32 VDD1.t7 VSUBS 0.386584f
C33 VDD1.n1 VSUBS 3.1787f
C34 VDD1.t5 VSUBS 0.386584f
C35 VDD1.t3 VSUBS 0.386584f
C36 VDD1.n2 VSUBS 3.1787f
C37 VDD1.n3 VSUBS 6.24823f
C38 VDD1.t1 VSUBS 0.386584f
C39 VDD1.t4 VSUBS 0.386584f
C40 VDD1.n4 VSUBS 3.15003f
C41 VDD1.n5 VSUBS 5.11173f
C42 VP.n0 VSUBS 0.044271f
C43 VP.t4 VSUBS 3.84009f
C44 VP.n1 VSUBS 0.043865f
C45 VP.n2 VSUBS 0.023536f
C46 VP.n3 VSUBS 0.043865f
C47 VP.n4 VSUBS 0.023536f
C48 VP.t2 VSUBS 3.84009f
C49 VP.n5 VSUBS 0.043865f
C50 VP.n6 VSUBS 0.023536f
C51 VP.n7 VSUBS 0.043865f
C52 VP.n8 VSUBS 0.023536f
C53 VP.t0 VSUBS 3.84009f
C54 VP.n9 VSUBS 0.043865f
C55 VP.n10 VSUBS 0.023536f
C56 VP.n11 VSUBS 0.043865f
C57 VP.n12 VSUBS 0.044271f
C58 VP.t1 VSUBS 3.84009f
C59 VP.n13 VSUBS 0.044271f
C60 VP.t3 VSUBS 3.84009f
C61 VP.n14 VSUBS 0.043865f
C62 VP.n15 VSUBS 0.023536f
C63 VP.n16 VSUBS 0.043865f
C64 VP.n17 VSUBS 0.023536f
C65 VP.t6 VSUBS 3.84009f
C66 VP.n18 VSUBS 0.043865f
C67 VP.n19 VSUBS 0.023536f
C68 VP.n20 VSUBS 0.043865f
C69 VP.n21 VSUBS 0.313376f
C70 VP.t5 VSUBS 3.84009f
C71 VP.t7 VSUBS 4.23227f
C72 VP.n22 VSUBS 1.34449f
C73 VP.n23 VSUBS 1.41135f
C74 VP.n24 VSUBS 0.028055f
C75 VP.n25 VSUBS 0.043865f
C76 VP.n26 VSUBS 0.023536f
C77 VP.n27 VSUBS 0.023536f
C78 VP.n28 VSUBS 0.023536f
C79 VP.n29 VSUBS 0.046777f
C80 VP.n30 VSUBS 0.019026f
C81 VP.n31 VSUBS 0.046777f
C82 VP.n32 VSUBS 0.023536f
C83 VP.n33 VSUBS 0.023536f
C84 VP.n34 VSUBS 0.023536f
C85 VP.n35 VSUBS 0.043865f
C86 VP.n36 VSUBS 0.028055f
C87 VP.n37 VSUBS 1.33056f
C88 VP.n38 VSUBS 0.038016f
C89 VP.n39 VSUBS 0.023536f
C90 VP.n40 VSUBS 0.023536f
C91 VP.n41 VSUBS 0.023536f
C92 VP.n42 VSUBS 0.043865f
C93 VP.n43 VSUBS 0.03567f
C94 VP.n44 VSUBS 0.033046f
C95 VP.n45 VSUBS 0.023536f
C96 VP.n46 VSUBS 0.023536f
C97 VP.n47 VSUBS 0.023536f
C98 VP.n48 VSUBS 0.043865f
C99 VP.n49 VSUBS 0.039749f
C100 VP.n50 VSUBS 1.43246f
C101 VP.n51 VSUBS 1.74477f
C102 VP.n52 VSUBS 1.75893f
C103 VP.n53 VSUBS 1.43246f
C104 VP.n54 VSUBS 0.039749f
C105 VP.n55 VSUBS 0.043865f
C106 VP.n56 VSUBS 0.023536f
C107 VP.n57 VSUBS 0.023536f
C108 VP.n58 VSUBS 0.023536f
C109 VP.n59 VSUBS 0.033046f
C110 VP.n60 VSUBS 0.03567f
C111 VP.n61 VSUBS 0.043865f
C112 VP.n62 VSUBS 0.023536f
C113 VP.n63 VSUBS 0.023536f
C114 VP.n64 VSUBS 0.023536f
C115 VP.n65 VSUBS 0.038016f
C116 VP.n66 VSUBS 1.33056f
C117 VP.n67 VSUBS 0.028055f
C118 VP.n68 VSUBS 0.043865f
C119 VP.n69 VSUBS 0.023536f
C120 VP.n70 VSUBS 0.023536f
C121 VP.n71 VSUBS 0.023536f
C122 VP.n72 VSUBS 0.046777f
C123 VP.n73 VSUBS 0.019026f
C124 VP.n74 VSUBS 0.046777f
C125 VP.n75 VSUBS 0.023536f
C126 VP.n76 VSUBS 0.023536f
C127 VP.n77 VSUBS 0.023536f
C128 VP.n78 VSUBS 0.043865f
C129 VP.n79 VSUBS 0.028055f
C130 VP.n80 VSUBS 1.33056f
C131 VP.n81 VSUBS 0.038016f
C132 VP.n82 VSUBS 0.023536f
C133 VP.n83 VSUBS 0.023536f
C134 VP.n84 VSUBS 0.023536f
C135 VP.n85 VSUBS 0.043865f
C136 VP.n86 VSUBS 0.03567f
C137 VP.n87 VSUBS 0.033046f
C138 VP.n88 VSUBS 0.023536f
C139 VP.n89 VSUBS 0.023536f
C140 VP.n90 VSUBS 0.023536f
C141 VP.n91 VSUBS 0.043865f
C142 VP.n92 VSUBS 0.039749f
C143 VP.n93 VSUBS 1.43246f
C144 VP.n94 VSUBS 0.075196f
C145 B.n0 VSUBS 0.004914f
C146 B.n1 VSUBS 0.004914f
C147 B.n2 VSUBS 0.007771f
C148 B.n3 VSUBS 0.007771f
C149 B.n4 VSUBS 0.007771f
C150 B.n5 VSUBS 0.007771f
C151 B.n6 VSUBS 0.007771f
C152 B.n7 VSUBS 0.007771f
C153 B.n8 VSUBS 0.007771f
C154 B.n9 VSUBS 0.007771f
C155 B.n10 VSUBS 0.007771f
C156 B.n11 VSUBS 0.007771f
C157 B.n12 VSUBS 0.007771f
C158 B.n13 VSUBS 0.007771f
C159 B.n14 VSUBS 0.007771f
C160 B.n15 VSUBS 0.007771f
C161 B.n16 VSUBS 0.007771f
C162 B.n17 VSUBS 0.007771f
C163 B.n18 VSUBS 0.007771f
C164 B.n19 VSUBS 0.007771f
C165 B.n20 VSUBS 0.007771f
C166 B.n21 VSUBS 0.007771f
C167 B.n22 VSUBS 0.007771f
C168 B.n23 VSUBS 0.007771f
C169 B.n24 VSUBS 0.007771f
C170 B.n25 VSUBS 0.007771f
C171 B.n26 VSUBS 0.007771f
C172 B.n27 VSUBS 0.007771f
C173 B.n28 VSUBS 0.007771f
C174 B.n29 VSUBS 0.007771f
C175 B.n30 VSUBS 0.007771f
C176 B.n31 VSUBS 0.007771f
C177 B.n32 VSUBS 0.007771f
C178 B.n33 VSUBS 0.007771f
C179 B.n34 VSUBS 0.007771f
C180 B.n35 VSUBS 0.007771f
C181 B.n36 VSUBS 0.007771f
C182 B.n37 VSUBS 0.017611f
C183 B.n38 VSUBS 0.007771f
C184 B.n39 VSUBS 0.007771f
C185 B.n40 VSUBS 0.007771f
C186 B.n41 VSUBS 0.007771f
C187 B.n42 VSUBS 0.007771f
C188 B.n43 VSUBS 0.007771f
C189 B.n44 VSUBS 0.007771f
C190 B.n45 VSUBS 0.007771f
C191 B.n46 VSUBS 0.007771f
C192 B.n47 VSUBS 0.007771f
C193 B.n48 VSUBS 0.007771f
C194 B.n49 VSUBS 0.007771f
C195 B.n50 VSUBS 0.007771f
C196 B.n51 VSUBS 0.007771f
C197 B.n52 VSUBS 0.007771f
C198 B.n53 VSUBS 0.007771f
C199 B.n54 VSUBS 0.007771f
C200 B.n55 VSUBS 0.007771f
C201 B.n56 VSUBS 0.007771f
C202 B.n57 VSUBS 0.007771f
C203 B.n58 VSUBS 0.007771f
C204 B.n59 VSUBS 0.007771f
C205 B.n60 VSUBS 0.007771f
C206 B.n61 VSUBS 0.007771f
C207 B.n62 VSUBS 0.007771f
C208 B.n63 VSUBS 0.007771f
C209 B.t8 VSUBS 0.558773f
C210 B.t7 VSUBS 0.591076f
C211 B.t6 VSUBS 3.05032f
C212 B.n64 VSUBS 0.356574f
C213 B.n65 VSUBS 0.086075f
C214 B.n66 VSUBS 0.007771f
C215 B.n67 VSUBS 0.007771f
C216 B.n68 VSUBS 0.007771f
C217 B.n69 VSUBS 0.007771f
C218 B.t2 VSUBS 0.558758f
C219 B.t1 VSUBS 0.591064f
C220 B.t0 VSUBS 3.05032f
C221 B.n70 VSUBS 0.356586f
C222 B.n71 VSUBS 0.086091f
C223 B.n72 VSUBS 0.007771f
C224 B.n73 VSUBS 0.007771f
C225 B.n74 VSUBS 0.007771f
C226 B.n75 VSUBS 0.007771f
C227 B.n76 VSUBS 0.007771f
C228 B.n77 VSUBS 0.007771f
C229 B.n78 VSUBS 0.007771f
C230 B.n79 VSUBS 0.007771f
C231 B.n80 VSUBS 0.007771f
C232 B.n81 VSUBS 0.007771f
C233 B.n82 VSUBS 0.007771f
C234 B.n83 VSUBS 0.007771f
C235 B.n84 VSUBS 0.007771f
C236 B.n85 VSUBS 0.007771f
C237 B.n86 VSUBS 0.007771f
C238 B.n87 VSUBS 0.007771f
C239 B.n88 VSUBS 0.007771f
C240 B.n89 VSUBS 0.007771f
C241 B.n90 VSUBS 0.007771f
C242 B.n91 VSUBS 0.007771f
C243 B.n92 VSUBS 0.007771f
C244 B.n93 VSUBS 0.007771f
C245 B.n94 VSUBS 0.007771f
C246 B.n95 VSUBS 0.007771f
C247 B.n96 VSUBS 0.007771f
C248 B.n97 VSUBS 0.017611f
C249 B.n98 VSUBS 0.007771f
C250 B.n99 VSUBS 0.007771f
C251 B.n100 VSUBS 0.007771f
C252 B.n101 VSUBS 0.007771f
C253 B.n102 VSUBS 0.007771f
C254 B.n103 VSUBS 0.007771f
C255 B.n104 VSUBS 0.007771f
C256 B.n105 VSUBS 0.007771f
C257 B.n106 VSUBS 0.007771f
C258 B.n107 VSUBS 0.007771f
C259 B.n108 VSUBS 0.007771f
C260 B.n109 VSUBS 0.007771f
C261 B.n110 VSUBS 0.007771f
C262 B.n111 VSUBS 0.007771f
C263 B.n112 VSUBS 0.007771f
C264 B.n113 VSUBS 0.007771f
C265 B.n114 VSUBS 0.007771f
C266 B.n115 VSUBS 0.007771f
C267 B.n116 VSUBS 0.007771f
C268 B.n117 VSUBS 0.007771f
C269 B.n118 VSUBS 0.007771f
C270 B.n119 VSUBS 0.007771f
C271 B.n120 VSUBS 0.007771f
C272 B.n121 VSUBS 0.007771f
C273 B.n122 VSUBS 0.007771f
C274 B.n123 VSUBS 0.007771f
C275 B.n124 VSUBS 0.007771f
C276 B.n125 VSUBS 0.007771f
C277 B.n126 VSUBS 0.007771f
C278 B.n127 VSUBS 0.007771f
C279 B.n128 VSUBS 0.007771f
C280 B.n129 VSUBS 0.007771f
C281 B.n130 VSUBS 0.007771f
C282 B.n131 VSUBS 0.007771f
C283 B.n132 VSUBS 0.007771f
C284 B.n133 VSUBS 0.007771f
C285 B.n134 VSUBS 0.007771f
C286 B.n135 VSUBS 0.007771f
C287 B.n136 VSUBS 0.007771f
C288 B.n137 VSUBS 0.007771f
C289 B.n138 VSUBS 0.007771f
C290 B.n139 VSUBS 0.007771f
C291 B.n140 VSUBS 0.007771f
C292 B.n141 VSUBS 0.007771f
C293 B.n142 VSUBS 0.007771f
C294 B.n143 VSUBS 0.007771f
C295 B.n144 VSUBS 0.007771f
C296 B.n145 VSUBS 0.007771f
C297 B.n146 VSUBS 0.007771f
C298 B.n147 VSUBS 0.007771f
C299 B.n148 VSUBS 0.007771f
C300 B.n149 VSUBS 0.007771f
C301 B.n150 VSUBS 0.007771f
C302 B.n151 VSUBS 0.007771f
C303 B.n152 VSUBS 0.007771f
C304 B.n153 VSUBS 0.007771f
C305 B.n154 VSUBS 0.007771f
C306 B.n155 VSUBS 0.007771f
C307 B.n156 VSUBS 0.007771f
C308 B.n157 VSUBS 0.007771f
C309 B.n158 VSUBS 0.007771f
C310 B.n159 VSUBS 0.007771f
C311 B.n160 VSUBS 0.007771f
C312 B.n161 VSUBS 0.007771f
C313 B.n162 VSUBS 0.007771f
C314 B.n163 VSUBS 0.007771f
C315 B.n164 VSUBS 0.007771f
C316 B.n165 VSUBS 0.007771f
C317 B.n166 VSUBS 0.007771f
C318 B.n167 VSUBS 0.007771f
C319 B.n168 VSUBS 0.017611f
C320 B.n169 VSUBS 0.007771f
C321 B.n170 VSUBS 0.007771f
C322 B.n171 VSUBS 0.007771f
C323 B.n172 VSUBS 0.007771f
C324 B.n173 VSUBS 0.007771f
C325 B.n174 VSUBS 0.007771f
C326 B.n175 VSUBS 0.007771f
C327 B.n176 VSUBS 0.007771f
C328 B.n177 VSUBS 0.007771f
C329 B.n178 VSUBS 0.007771f
C330 B.n179 VSUBS 0.007771f
C331 B.n180 VSUBS 0.007771f
C332 B.n181 VSUBS 0.007771f
C333 B.n182 VSUBS 0.007771f
C334 B.n183 VSUBS 0.007771f
C335 B.n184 VSUBS 0.007771f
C336 B.n185 VSUBS 0.007771f
C337 B.n186 VSUBS 0.007771f
C338 B.n187 VSUBS 0.007771f
C339 B.n188 VSUBS 0.007771f
C340 B.n189 VSUBS 0.007771f
C341 B.n190 VSUBS 0.007771f
C342 B.n191 VSUBS 0.007771f
C343 B.n192 VSUBS 0.007771f
C344 B.n193 VSUBS 0.007771f
C345 B.t10 VSUBS 0.558758f
C346 B.t11 VSUBS 0.591064f
C347 B.t9 VSUBS 3.05032f
C348 B.n194 VSUBS 0.356586f
C349 B.n195 VSUBS 0.086091f
C350 B.n196 VSUBS 0.018005f
C351 B.n197 VSUBS 0.007771f
C352 B.n198 VSUBS 0.007771f
C353 B.n199 VSUBS 0.007771f
C354 B.n200 VSUBS 0.007771f
C355 B.n201 VSUBS 0.007771f
C356 B.t4 VSUBS 0.558773f
C357 B.t5 VSUBS 0.591076f
C358 B.t3 VSUBS 3.05032f
C359 B.n202 VSUBS 0.356574f
C360 B.n203 VSUBS 0.086075f
C361 B.n204 VSUBS 0.007771f
C362 B.n205 VSUBS 0.007771f
C363 B.n206 VSUBS 0.007771f
C364 B.n207 VSUBS 0.007771f
C365 B.n208 VSUBS 0.007771f
C366 B.n209 VSUBS 0.007771f
C367 B.n210 VSUBS 0.007771f
C368 B.n211 VSUBS 0.007771f
C369 B.n212 VSUBS 0.007771f
C370 B.n213 VSUBS 0.007771f
C371 B.n214 VSUBS 0.007771f
C372 B.n215 VSUBS 0.007771f
C373 B.n216 VSUBS 0.007771f
C374 B.n217 VSUBS 0.007771f
C375 B.n218 VSUBS 0.007771f
C376 B.n219 VSUBS 0.007771f
C377 B.n220 VSUBS 0.007771f
C378 B.n221 VSUBS 0.007771f
C379 B.n222 VSUBS 0.007771f
C380 B.n223 VSUBS 0.007771f
C381 B.n224 VSUBS 0.007771f
C382 B.n225 VSUBS 0.007771f
C383 B.n226 VSUBS 0.007771f
C384 B.n227 VSUBS 0.007771f
C385 B.n228 VSUBS 0.018274f
C386 B.n229 VSUBS 0.007771f
C387 B.n230 VSUBS 0.007771f
C388 B.n231 VSUBS 0.007771f
C389 B.n232 VSUBS 0.007771f
C390 B.n233 VSUBS 0.007771f
C391 B.n234 VSUBS 0.007771f
C392 B.n235 VSUBS 0.007771f
C393 B.n236 VSUBS 0.007771f
C394 B.n237 VSUBS 0.007771f
C395 B.n238 VSUBS 0.007771f
C396 B.n239 VSUBS 0.007771f
C397 B.n240 VSUBS 0.007771f
C398 B.n241 VSUBS 0.007771f
C399 B.n242 VSUBS 0.007771f
C400 B.n243 VSUBS 0.007771f
C401 B.n244 VSUBS 0.007771f
C402 B.n245 VSUBS 0.007771f
C403 B.n246 VSUBS 0.007771f
C404 B.n247 VSUBS 0.007771f
C405 B.n248 VSUBS 0.007771f
C406 B.n249 VSUBS 0.007771f
C407 B.n250 VSUBS 0.007771f
C408 B.n251 VSUBS 0.007771f
C409 B.n252 VSUBS 0.007771f
C410 B.n253 VSUBS 0.007771f
C411 B.n254 VSUBS 0.007771f
C412 B.n255 VSUBS 0.007771f
C413 B.n256 VSUBS 0.007771f
C414 B.n257 VSUBS 0.007771f
C415 B.n258 VSUBS 0.007771f
C416 B.n259 VSUBS 0.007771f
C417 B.n260 VSUBS 0.007771f
C418 B.n261 VSUBS 0.007771f
C419 B.n262 VSUBS 0.007771f
C420 B.n263 VSUBS 0.007771f
C421 B.n264 VSUBS 0.007771f
C422 B.n265 VSUBS 0.007771f
C423 B.n266 VSUBS 0.007771f
C424 B.n267 VSUBS 0.007771f
C425 B.n268 VSUBS 0.007771f
C426 B.n269 VSUBS 0.007771f
C427 B.n270 VSUBS 0.007771f
C428 B.n271 VSUBS 0.007771f
C429 B.n272 VSUBS 0.007771f
C430 B.n273 VSUBS 0.007771f
C431 B.n274 VSUBS 0.007771f
C432 B.n275 VSUBS 0.007771f
C433 B.n276 VSUBS 0.007771f
C434 B.n277 VSUBS 0.007771f
C435 B.n278 VSUBS 0.007771f
C436 B.n279 VSUBS 0.007771f
C437 B.n280 VSUBS 0.007771f
C438 B.n281 VSUBS 0.007771f
C439 B.n282 VSUBS 0.007771f
C440 B.n283 VSUBS 0.007771f
C441 B.n284 VSUBS 0.007771f
C442 B.n285 VSUBS 0.007771f
C443 B.n286 VSUBS 0.007771f
C444 B.n287 VSUBS 0.007771f
C445 B.n288 VSUBS 0.007771f
C446 B.n289 VSUBS 0.007771f
C447 B.n290 VSUBS 0.007771f
C448 B.n291 VSUBS 0.007771f
C449 B.n292 VSUBS 0.007771f
C450 B.n293 VSUBS 0.007771f
C451 B.n294 VSUBS 0.007771f
C452 B.n295 VSUBS 0.007771f
C453 B.n296 VSUBS 0.007771f
C454 B.n297 VSUBS 0.007771f
C455 B.n298 VSUBS 0.007771f
C456 B.n299 VSUBS 0.007771f
C457 B.n300 VSUBS 0.007771f
C458 B.n301 VSUBS 0.007771f
C459 B.n302 VSUBS 0.007771f
C460 B.n303 VSUBS 0.007771f
C461 B.n304 VSUBS 0.007771f
C462 B.n305 VSUBS 0.007771f
C463 B.n306 VSUBS 0.007771f
C464 B.n307 VSUBS 0.007771f
C465 B.n308 VSUBS 0.007771f
C466 B.n309 VSUBS 0.007771f
C467 B.n310 VSUBS 0.007771f
C468 B.n311 VSUBS 0.007771f
C469 B.n312 VSUBS 0.007771f
C470 B.n313 VSUBS 0.007771f
C471 B.n314 VSUBS 0.007771f
C472 B.n315 VSUBS 0.007771f
C473 B.n316 VSUBS 0.007771f
C474 B.n317 VSUBS 0.007771f
C475 B.n318 VSUBS 0.007771f
C476 B.n319 VSUBS 0.007771f
C477 B.n320 VSUBS 0.007771f
C478 B.n321 VSUBS 0.007771f
C479 B.n322 VSUBS 0.007771f
C480 B.n323 VSUBS 0.007771f
C481 B.n324 VSUBS 0.007771f
C482 B.n325 VSUBS 0.007771f
C483 B.n326 VSUBS 0.007771f
C484 B.n327 VSUBS 0.007771f
C485 B.n328 VSUBS 0.007771f
C486 B.n329 VSUBS 0.007771f
C487 B.n330 VSUBS 0.007771f
C488 B.n331 VSUBS 0.007771f
C489 B.n332 VSUBS 0.007771f
C490 B.n333 VSUBS 0.007771f
C491 B.n334 VSUBS 0.007771f
C492 B.n335 VSUBS 0.007771f
C493 B.n336 VSUBS 0.007771f
C494 B.n337 VSUBS 0.007771f
C495 B.n338 VSUBS 0.007771f
C496 B.n339 VSUBS 0.007771f
C497 B.n340 VSUBS 0.007771f
C498 B.n341 VSUBS 0.007771f
C499 B.n342 VSUBS 0.007771f
C500 B.n343 VSUBS 0.007771f
C501 B.n344 VSUBS 0.007771f
C502 B.n345 VSUBS 0.007771f
C503 B.n346 VSUBS 0.007771f
C504 B.n347 VSUBS 0.007771f
C505 B.n348 VSUBS 0.007771f
C506 B.n349 VSUBS 0.007771f
C507 B.n350 VSUBS 0.007771f
C508 B.n351 VSUBS 0.007771f
C509 B.n352 VSUBS 0.007771f
C510 B.n353 VSUBS 0.007771f
C511 B.n354 VSUBS 0.007771f
C512 B.n355 VSUBS 0.007771f
C513 B.n356 VSUBS 0.007771f
C514 B.n357 VSUBS 0.007771f
C515 B.n358 VSUBS 0.007771f
C516 B.n359 VSUBS 0.007771f
C517 B.n360 VSUBS 0.007771f
C518 B.n361 VSUBS 0.007771f
C519 B.n362 VSUBS 0.007771f
C520 B.n363 VSUBS 0.007771f
C521 B.n364 VSUBS 0.007771f
C522 B.n365 VSUBS 0.007771f
C523 B.n366 VSUBS 0.007771f
C524 B.n367 VSUBS 0.017611f
C525 B.n368 VSUBS 0.017611f
C526 B.n369 VSUBS 0.018274f
C527 B.n370 VSUBS 0.007771f
C528 B.n371 VSUBS 0.007771f
C529 B.n372 VSUBS 0.007771f
C530 B.n373 VSUBS 0.007771f
C531 B.n374 VSUBS 0.007771f
C532 B.n375 VSUBS 0.007771f
C533 B.n376 VSUBS 0.007771f
C534 B.n377 VSUBS 0.007771f
C535 B.n378 VSUBS 0.007771f
C536 B.n379 VSUBS 0.007771f
C537 B.n380 VSUBS 0.007771f
C538 B.n381 VSUBS 0.007771f
C539 B.n382 VSUBS 0.007771f
C540 B.n383 VSUBS 0.007771f
C541 B.n384 VSUBS 0.007771f
C542 B.n385 VSUBS 0.007771f
C543 B.n386 VSUBS 0.007771f
C544 B.n387 VSUBS 0.007771f
C545 B.n388 VSUBS 0.007771f
C546 B.n389 VSUBS 0.007771f
C547 B.n390 VSUBS 0.007771f
C548 B.n391 VSUBS 0.007771f
C549 B.n392 VSUBS 0.007771f
C550 B.n393 VSUBS 0.007771f
C551 B.n394 VSUBS 0.007771f
C552 B.n395 VSUBS 0.007771f
C553 B.n396 VSUBS 0.007771f
C554 B.n397 VSUBS 0.007771f
C555 B.n398 VSUBS 0.007771f
C556 B.n399 VSUBS 0.007771f
C557 B.n400 VSUBS 0.007771f
C558 B.n401 VSUBS 0.007771f
C559 B.n402 VSUBS 0.007771f
C560 B.n403 VSUBS 0.007771f
C561 B.n404 VSUBS 0.007771f
C562 B.n405 VSUBS 0.007771f
C563 B.n406 VSUBS 0.007771f
C564 B.n407 VSUBS 0.007771f
C565 B.n408 VSUBS 0.007771f
C566 B.n409 VSUBS 0.007771f
C567 B.n410 VSUBS 0.007771f
C568 B.n411 VSUBS 0.007771f
C569 B.n412 VSUBS 0.007771f
C570 B.n413 VSUBS 0.007771f
C571 B.n414 VSUBS 0.007771f
C572 B.n415 VSUBS 0.007771f
C573 B.n416 VSUBS 0.007771f
C574 B.n417 VSUBS 0.007771f
C575 B.n418 VSUBS 0.007771f
C576 B.n419 VSUBS 0.007771f
C577 B.n420 VSUBS 0.007771f
C578 B.n421 VSUBS 0.007771f
C579 B.n422 VSUBS 0.007771f
C580 B.n423 VSUBS 0.007771f
C581 B.n424 VSUBS 0.007771f
C582 B.n425 VSUBS 0.007771f
C583 B.n426 VSUBS 0.007771f
C584 B.n427 VSUBS 0.007771f
C585 B.n428 VSUBS 0.007771f
C586 B.n429 VSUBS 0.007771f
C587 B.n430 VSUBS 0.007771f
C588 B.n431 VSUBS 0.007771f
C589 B.n432 VSUBS 0.007771f
C590 B.n433 VSUBS 0.007771f
C591 B.n434 VSUBS 0.007771f
C592 B.n435 VSUBS 0.007771f
C593 B.n436 VSUBS 0.007771f
C594 B.n437 VSUBS 0.007771f
C595 B.n438 VSUBS 0.007771f
C596 B.n439 VSUBS 0.007771f
C597 B.n440 VSUBS 0.007771f
C598 B.n441 VSUBS 0.007771f
C599 B.n442 VSUBS 0.007771f
C600 B.n443 VSUBS 0.007771f
C601 B.n444 VSUBS 0.005371f
C602 B.n445 VSUBS 0.018005f
C603 B.n446 VSUBS 0.006286f
C604 B.n447 VSUBS 0.007771f
C605 B.n448 VSUBS 0.007771f
C606 B.n449 VSUBS 0.007771f
C607 B.n450 VSUBS 0.007771f
C608 B.n451 VSUBS 0.007771f
C609 B.n452 VSUBS 0.007771f
C610 B.n453 VSUBS 0.007771f
C611 B.n454 VSUBS 0.007771f
C612 B.n455 VSUBS 0.007771f
C613 B.n456 VSUBS 0.007771f
C614 B.n457 VSUBS 0.007771f
C615 B.n458 VSUBS 0.006286f
C616 B.n459 VSUBS 0.007771f
C617 B.n460 VSUBS 0.007771f
C618 B.n461 VSUBS 0.005371f
C619 B.n462 VSUBS 0.007771f
C620 B.n463 VSUBS 0.007771f
C621 B.n464 VSUBS 0.007771f
C622 B.n465 VSUBS 0.007771f
C623 B.n466 VSUBS 0.007771f
C624 B.n467 VSUBS 0.007771f
C625 B.n468 VSUBS 0.007771f
C626 B.n469 VSUBS 0.007771f
C627 B.n470 VSUBS 0.007771f
C628 B.n471 VSUBS 0.007771f
C629 B.n472 VSUBS 0.007771f
C630 B.n473 VSUBS 0.007771f
C631 B.n474 VSUBS 0.007771f
C632 B.n475 VSUBS 0.007771f
C633 B.n476 VSUBS 0.007771f
C634 B.n477 VSUBS 0.007771f
C635 B.n478 VSUBS 0.007771f
C636 B.n479 VSUBS 0.007771f
C637 B.n480 VSUBS 0.007771f
C638 B.n481 VSUBS 0.007771f
C639 B.n482 VSUBS 0.007771f
C640 B.n483 VSUBS 0.007771f
C641 B.n484 VSUBS 0.007771f
C642 B.n485 VSUBS 0.007771f
C643 B.n486 VSUBS 0.007771f
C644 B.n487 VSUBS 0.007771f
C645 B.n488 VSUBS 0.007771f
C646 B.n489 VSUBS 0.007771f
C647 B.n490 VSUBS 0.007771f
C648 B.n491 VSUBS 0.007771f
C649 B.n492 VSUBS 0.007771f
C650 B.n493 VSUBS 0.007771f
C651 B.n494 VSUBS 0.007771f
C652 B.n495 VSUBS 0.007771f
C653 B.n496 VSUBS 0.007771f
C654 B.n497 VSUBS 0.007771f
C655 B.n498 VSUBS 0.007771f
C656 B.n499 VSUBS 0.007771f
C657 B.n500 VSUBS 0.007771f
C658 B.n501 VSUBS 0.007771f
C659 B.n502 VSUBS 0.007771f
C660 B.n503 VSUBS 0.007771f
C661 B.n504 VSUBS 0.007771f
C662 B.n505 VSUBS 0.007771f
C663 B.n506 VSUBS 0.007771f
C664 B.n507 VSUBS 0.007771f
C665 B.n508 VSUBS 0.007771f
C666 B.n509 VSUBS 0.007771f
C667 B.n510 VSUBS 0.007771f
C668 B.n511 VSUBS 0.007771f
C669 B.n512 VSUBS 0.007771f
C670 B.n513 VSUBS 0.007771f
C671 B.n514 VSUBS 0.007771f
C672 B.n515 VSUBS 0.007771f
C673 B.n516 VSUBS 0.007771f
C674 B.n517 VSUBS 0.007771f
C675 B.n518 VSUBS 0.007771f
C676 B.n519 VSUBS 0.007771f
C677 B.n520 VSUBS 0.007771f
C678 B.n521 VSUBS 0.007771f
C679 B.n522 VSUBS 0.007771f
C680 B.n523 VSUBS 0.007771f
C681 B.n524 VSUBS 0.007771f
C682 B.n525 VSUBS 0.007771f
C683 B.n526 VSUBS 0.007771f
C684 B.n527 VSUBS 0.007771f
C685 B.n528 VSUBS 0.007771f
C686 B.n529 VSUBS 0.007771f
C687 B.n530 VSUBS 0.007771f
C688 B.n531 VSUBS 0.007771f
C689 B.n532 VSUBS 0.007771f
C690 B.n533 VSUBS 0.007771f
C691 B.n534 VSUBS 0.007771f
C692 B.n535 VSUBS 0.018274f
C693 B.n536 VSUBS 0.018274f
C694 B.n537 VSUBS 0.017611f
C695 B.n538 VSUBS 0.007771f
C696 B.n539 VSUBS 0.007771f
C697 B.n540 VSUBS 0.007771f
C698 B.n541 VSUBS 0.007771f
C699 B.n542 VSUBS 0.007771f
C700 B.n543 VSUBS 0.007771f
C701 B.n544 VSUBS 0.007771f
C702 B.n545 VSUBS 0.007771f
C703 B.n546 VSUBS 0.007771f
C704 B.n547 VSUBS 0.007771f
C705 B.n548 VSUBS 0.007771f
C706 B.n549 VSUBS 0.007771f
C707 B.n550 VSUBS 0.007771f
C708 B.n551 VSUBS 0.007771f
C709 B.n552 VSUBS 0.007771f
C710 B.n553 VSUBS 0.007771f
C711 B.n554 VSUBS 0.007771f
C712 B.n555 VSUBS 0.007771f
C713 B.n556 VSUBS 0.007771f
C714 B.n557 VSUBS 0.007771f
C715 B.n558 VSUBS 0.007771f
C716 B.n559 VSUBS 0.007771f
C717 B.n560 VSUBS 0.007771f
C718 B.n561 VSUBS 0.007771f
C719 B.n562 VSUBS 0.007771f
C720 B.n563 VSUBS 0.007771f
C721 B.n564 VSUBS 0.007771f
C722 B.n565 VSUBS 0.007771f
C723 B.n566 VSUBS 0.007771f
C724 B.n567 VSUBS 0.007771f
C725 B.n568 VSUBS 0.007771f
C726 B.n569 VSUBS 0.007771f
C727 B.n570 VSUBS 0.007771f
C728 B.n571 VSUBS 0.007771f
C729 B.n572 VSUBS 0.007771f
C730 B.n573 VSUBS 0.007771f
C731 B.n574 VSUBS 0.007771f
C732 B.n575 VSUBS 0.007771f
C733 B.n576 VSUBS 0.007771f
C734 B.n577 VSUBS 0.007771f
C735 B.n578 VSUBS 0.007771f
C736 B.n579 VSUBS 0.007771f
C737 B.n580 VSUBS 0.007771f
C738 B.n581 VSUBS 0.007771f
C739 B.n582 VSUBS 0.007771f
C740 B.n583 VSUBS 0.007771f
C741 B.n584 VSUBS 0.007771f
C742 B.n585 VSUBS 0.007771f
C743 B.n586 VSUBS 0.007771f
C744 B.n587 VSUBS 0.007771f
C745 B.n588 VSUBS 0.007771f
C746 B.n589 VSUBS 0.007771f
C747 B.n590 VSUBS 0.007771f
C748 B.n591 VSUBS 0.007771f
C749 B.n592 VSUBS 0.007771f
C750 B.n593 VSUBS 0.007771f
C751 B.n594 VSUBS 0.007771f
C752 B.n595 VSUBS 0.007771f
C753 B.n596 VSUBS 0.007771f
C754 B.n597 VSUBS 0.007771f
C755 B.n598 VSUBS 0.007771f
C756 B.n599 VSUBS 0.007771f
C757 B.n600 VSUBS 0.007771f
C758 B.n601 VSUBS 0.007771f
C759 B.n602 VSUBS 0.007771f
C760 B.n603 VSUBS 0.007771f
C761 B.n604 VSUBS 0.007771f
C762 B.n605 VSUBS 0.007771f
C763 B.n606 VSUBS 0.007771f
C764 B.n607 VSUBS 0.007771f
C765 B.n608 VSUBS 0.007771f
C766 B.n609 VSUBS 0.007771f
C767 B.n610 VSUBS 0.007771f
C768 B.n611 VSUBS 0.007771f
C769 B.n612 VSUBS 0.007771f
C770 B.n613 VSUBS 0.007771f
C771 B.n614 VSUBS 0.007771f
C772 B.n615 VSUBS 0.007771f
C773 B.n616 VSUBS 0.007771f
C774 B.n617 VSUBS 0.007771f
C775 B.n618 VSUBS 0.007771f
C776 B.n619 VSUBS 0.007771f
C777 B.n620 VSUBS 0.007771f
C778 B.n621 VSUBS 0.007771f
C779 B.n622 VSUBS 0.007771f
C780 B.n623 VSUBS 0.007771f
C781 B.n624 VSUBS 0.007771f
C782 B.n625 VSUBS 0.007771f
C783 B.n626 VSUBS 0.007771f
C784 B.n627 VSUBS 0.007771f
C785 B.n628 VSUBS 0.007771f
C786 B.n629 VSUBS 0.007771f
C787 B.n630 VSUBS 0.007771f
C788 B.n631 VSUBS 0.007771f
C789 B.n632 VSUBS 0.007771f
C790 B.n633 VSUBS 0.007771f
C791 B.n634 VSUBS 0.007771f
C792 B.n635 VSUBS 0.007771f
C793 B.n636 VSUBS 0.007771f
C794 B.n637 VSUBS 0.007771f
C795 B.n638 VSUBS 0.007771f
C796 B.n639 VSUBS 0.007771f
C797 B.n640 VSUBS 0.007771f
C798 B.n641 VSUBS 0.007771f
C799 B.n642 VSUBS 0.007771f
C800 B.n643 VSUBS 0.007771f
C801 B.n644 VSUBS 0.007771f
C802 B.n645 VSUBS 0.007771f
C803 B.n646 VSUBS 0.007771f
C804 B.n647 VSUBS 0.007771f
C805 B.n648 VSUBS 0.007771f
C806 B.n649 VSUBS 0.007771f
C807 B.n650 VSUBS 0.007771f
C808 B.n651 VSUBS 0.007771f
C809 B.n652 VSUBS 0.007771f
C810 B.n653 VSUBS 0.007771f
C811 B.n654 VSUBS 0.007771f
C812 B.n655 VSUBS 0.007771f
C813 B.n656 VSUBS 0.007771f
C814 B.n657 VSUBS 0.007771f
C815 B.n658 VSUBS 0.007771f
C816 B.n659 VSUBS 0.007771f
C817 B.n660 VSUBS 0.007771f
C818 B.n661 VSUBS 0.007771f
C819 B.n662 VSUBS 0.007771f
C820 B.n663 VSUBS 0.007771f
C821 B.n664 VSUBS 0.007771f
C822 B.n665 VSUBS 0.007771f
C823 B.n666 VSUBS 0.007771f
C824 B.n667 VSUBS 0.007771f
C825 B.n668 VSUBS 0.007771f
C826 B.n669 VSUBS 0.007771f
C827 B.n670 VSUBS 0.007771f
C828 B.n671 VSUBS 0.007771f
C829 B.n672 VSUBS 0.007771f
C830 B.n673 VSUBS 0.007771f
C831 B.n674 VSUBS 0.007771f
C832 B.n675 VSUBS 0.007771f
C833 B.n676 VSUBS 0.007771f
C834 B.n677 VSUBS 0.007771f
C835 B.n678 VSUBS 0.007771f
C836 B.n679 VSUBS 0.007771f
C837 B.n680 VSUBS 0.007771f
C838 B.n681 VSUBS 0.007771f
C839 B.n682 VSUBS 0.007771f
C840 B.n683 VSUBS 0.007771f
C841 B.n684 VSUBS 0.007771f
C842 B.n685 VSUBS 0.007771f
C843 B.n686 VSUBS 0.007771f
C844 B.n687 VSUBS 0.007771f
C845 B.n688 VSUBS 0.007771f
C846 B.n689 VSUBS 0.007771f
C847 B.n690 VSUBS 0.007771f
C848 B.n691 VSUBS 0.007771f
C849 B.n692 VSUBS 0.007771f
C850 B.n693 VSUBS 0.007771f
C851 B.n694 VSUBS 0.007771f
C852 B.n695 VSUBS 0.007771f
C853 B.n696 VSUBS 0.007771f
C854 B.n697 VSUBS 0.007771f
C855 B.n698 VSUBS 0.007771f
C856 B.n699 VSUBS 0.007771f
C857 B.n700 VSUBS 0.007771f
C858 B.n701 VSUBS 0.007771f
C859 B.n702 VSUBS 0.007771f
C860 B.n703 VSUBS 0.007771f
C861 B.n704 VSUBS 0.007771f
C862 B.n705 VSUBS 0.007771f
C863 B.n706 VSUBS 0.007771f
C864 B.n707 VSUBS 0.007771f
C865 B.n708 VSUBS 0.007771f
C866 B.n709 VSUBS 0.007771f
C867 B.n710 VSUBS 0.007771f
C868 B.n711 VSUBS 0.007771f
C869 B.n712 VSUBS 0.007771f
C870 B.n713 VSUBS 0.007771f
C871 B.n714 VSUBS 0.007771f
C872 B.n715 VSUBS 0.007771f
C873 B.n716 VSUBS 0.007771f
C874 B.n717 VSUBS 0.007771f
C875 B.n718 VSUBS 0.007771f
C876 B.n719 VSUBS 0.007771f
C877 B.n720 VSUBS 0.007771f
C878 B.n721 VSUBS 0.007771f
C879 B.n722 VSUBS 0.007771f
C880 B.n723 VSUBS 0.007771f
C881 B.n724 VSUBS 0.007771f
C882 B.n725 VSUBS 0.007771f
C883 B.n726 VSUBS 0.007771f
C884 B.n727 VSUBS 0.007771f
C885 B.n728 VSUBS 0.007771f
C886 B.n729 VSUBS 0.007771f
C887 B.n730 VSUBS 0.007771f
C888 B.n731 VSUBS 0.007771f
C889 B.n732 VSUBS 0.007771f
C890 B.n733 VSUBS 0.007771f
C891 B.n734 VSUBS 0.007771f
C892 B.n735 VSUBS 0.007771f
C893 B.n736 VSUBS 0.007771f
C894 B.n737 VSUBS 0.007771f
C895 B.n738 VSUBS 0.007771f
C896 B.n739 VSUBS 0.007771f
C897 B.n740 VSUBS 0.007771f
C898 B.n741 VSUBS 0.007771f
C899 B.n742 VSUBS 0.007771f
C900 B.n743 VSUBS 0.007771f
C901 B.n744 VSUBS 0.007771f
C902 B.n745 VSUBS 0.007771f
C903 B.n746 VSUBS 0.007771f
C904 B.n747 VSUBS 0.007771f
C905 B.n748 VSUBS 0.007771f
C906 B.n749 VSUBS 0.007771f
C907 B.n750 VSUBS 0.018548f
C908 B.n751 VSUBS 0.017337f
C909 B.n752 VSUBS 0.018274f
C910 B.n753 VSUBS 0.007771f
C911 B.n754 VSUBS 0.007771f
C912 B.n755 VSUBS 0.007771f
C913 B.n756 VSUBS 0.007771f
C914 B.n757 VSUBS 0.007771f
C915 B.n758 VSUBS 0.007771f
C916 B.n759 VSUBS 0.007771f
C917 B.n760 VSUBS 0.007771f
C918 B.n761 VSUBS 0.007771f
C919 B.n762 VSUBS 0.007771f
C920 B.n763 VSUBS 0.007771f
C921 B.n764 VSUBS 0.007771f
C922 B.n765 VSUBS 0.007771f
C923 B.n766 VSUBS 0.007771f
C924 B.n767 VSUBS 0.007771f
C925 B.n768 VSUBS 0.007771f
C926 B.n769 VSUBS 0.007771f
C927 B.n770 VSUBS 0.007771f
C928 B.n771 VSUBS 0.007771f
C929 B.n772 VSUBS 0.007771f
C930 B.n773 VSUBS 0.007771f
C931 B.n774 VSUBS 0.007771f
C932 B.n775 VSUBS 0.007771f
C933 B.n776 VSUBS 0.007771f
C934 B.n777 VSUBS 0.007771f
C935 B.n778 VSUBS 0.007771f
C936 B.n779 VSUBS 0.007771f
C937 B.n780 VSUBS 0.007771f
C938 B.n781 VSUBS 0.007771f
C939 B.n782 VSUBS 0.007771f
C940 B.n783 VSUBS 0.007771f
C941 B.n784 VSUBS 0.007771f
C942 B.n785 VSUBS 0.007771f
C943 B.n786 VSUBS 0.007771f
C944 B.n787 VSUBS 0.007771f
C945 B.n788 VSUBS 0.007771f
C946 B.n789 VSUBS 0.007771f
C947 B.n790 VSUBS 0.007771f
C948 B.n791 VSUBS 0.007771f
C949 B.n792 VSUBS 0.007771f
C950 B.n793 VSUBS 0.007771f
C951 B.n794 VSUBS 0.007771f
C952 B.n795 VSUBS 0.007771f
C953 B.n796 VSUBS 0.007771f
C954 B.n797 VSUBS 0.007771f
C955 B.n798 VSUBS 0.007771f
C956 B.n799 VSUBS 0.007771f
C957 B.n800 VSUBS 0.007771f
C958 B.n801 VSUBS 0.007771f
C959 B.n802 VSUBS 0.007771f
C960 B.n803 VSUBS 0.007771f
C961 B.n804 VSUBS 0.007771f
C962 B.n805 VSUBS 0.007771f
C963 B.n806 VSUBS 0.007771f
C964 B.n807 VSUBS 0.007771f
C965 B.n808 VSUBS 0.007771f
C966 B.n809 VSUBS 0.007771f
C967 B.n810 VSUBS 0.007771f
C968 B.n811 VSUBS 0.007771f
C969 B.n812 VSUBS 0.007771f
C970 B.n813 VSUBS 0.007771f
C971 B.n814 VSUBS 0.007771f
C972 B.n815 VSUBS 0.007771f
C973 B.n816 VSUBS 0.007771f
C974 B.n817 VSUBS 0.007771f
C975 B.n818 VSUBS 0.007771f
C976 B.n819 VSUBS 0.007771f
C977 B.n820 VSUBS 0.007771f
C978 B.n821 VSUBS 0.007771f
C979 B.n822 VSUBS 0.007771f
C980 B.n823 VSUBS 0.007771f
C981 B.n824 VSUBS 0.007771f
C982 B.n825 VSUBS 0.007771f
C983 B.n826 VSUBS 0.007771f
C984 B.n827 VSUBS 0.005371f
C985 B.n828 VSUBS 0.018005f
C986 B.n829 VSUBS 0.006286f
C987 B.n830 VSUBS 0.007771f
C988 B.n831 VSUBS 0.007771f
C989 B.n832 VSUBS 0.007771f
C990 B.n833 VSUBS 0.007771f
C991 B.n834 VSUBS 0.007771f
C992 B.n835 VSUBS 0.007771f
C993 B.n836 VSUBS 0.007771f
C994 B.n837 VSUBS 0.007771f
C995 B.n838 VSUBS 0.007771f
C996 B.n839 VSUBS 0.007771f
C997 B.n840 VSUBS 0.007771f
C998 B.n841 VSUBS 0.006286f
C999 B.n842 VSUBS 0.018005f
C1000 B.n843 VSUBS 0.005371f
C1001 B.n844 VSUBS 0.007771f
C1002 B.n845 VSUBS 0.007771f
C1003 B.n846 VSUBS 0.007771f
C1004 B.n847 VSUBS 0.007771f
C1005 B.n848 VSUBS 0.007771f
C1006 B.n849 VSUBS 0.007771f
C1007 B.n850 VSUBS 0.007771f
C1008 B.n851 VSUBS 0.007771f
C1009 B.n852 VSUBS 0.007771f
C1010 B.n853 VSUBS 0.007771f
C1011 B.n854 VSUBS 0.007771f
C1012 B.n855 VSUBS 0.007771f
C1013 B.n856 VSUBS 0.007771f
C1014 B.n857 VSUBS 0.007771f
C1015 B.n858 VSUBS 0.007771f
C1016 B.n859 VSUBS 0.007771f
C1017 B.n860 VSUBS 0.007771f
C1018 B.n861 VSUBS 0.007771f
C1019 B.n862 VSUBS 0.007771f
C1020 B.n863 VSUBS 0.007771f
C1021 B.n864 VSUBS 0.007771f
C1022 B.n865 VSUBS 0.007771f
C1023 B.n866 VSUBS 0.007771f
C1024 B.n867 VSUBS 0.007771f
C1025 B.n868 VSUBS 0.007771f
C1026 B.n869 VSUBS 0.007771f
C1027 B.n870 VSUBS 0.007771f
C1028 B.n871 VSUBS 0.007771f
C1029 B.n872 VSUBS 0.007771f
C1030 B.n873 VSUBS 0.007771f
C1031 B.n874 VSUBS 0.007771f
C1032 B.n875 VSUBS 0.007771f
C1033 B.n876 VSUBS 0.007771f
C1034 B.n877 VSUBS 0.007771f
C1035 B.n878 VSUBS 0.007771f
C1036 B.n879 VSUBS 0.007771f
C1037 B.n880 VSUBS 0.007771f
C1038 B.n881 VSUBS 0.007771f
C1039 B.n882 VSUBS 0.007771f
C1040 B.n883 VSUBS 0.007771f
C1041 B.n884 VSUBS 0.007771f
C1042 B.n885 VSUBS 0.007771f
C1043 B.n886 VSUBS 0.007771f
C1044 B.n887 VSUBS 0.007771f
C1045 B.n888 VSUBS 0.007771f
C1046 B.n889 VSUBS 0.007771f
C1047 B.n890 VSUBS 0.007771f
C1048 B.n891 VSUBS 0.007771f
C1049 B.n892 VSUBS 0.007771f
C1050 B.n893 VSUBS 0.007771f
C1051 B.n894 VSUBS 0.007771f
C1052 B.n895 VSUBS 0.007771f
C1053 B.n896 VSUBS 0.007771f
C1054 B.n897 VSUBS 0.007771f
C1055 B.n898 VSUBS 0.007771f
C1056 B.n899 VSUBS 0.007771f
C1057 B.n900 VSUBS 0.007771f
C1058 B.n901 VSUBS 0.007771f
C1059 B.n902 VSUBS 0.007771f
C1060 B.n903 VSUBS 0.007771f
C1061 B.n904 VSUBS 0.007771f
C1062 B.n905 VSUBS 0.007771f
C1063 B.n906 VSUBS 0.007771f
C1064 B.n907 VSUBS 0.007771f
C1065 B.n908 VSUBS 0.007771f
C1066 B.n909 VSUBS 0.007771f
C1067 B.n910 VSUBS 0.007771f
C1068 B.n911 VSUBS 0.007771f
C1069 B.n912 VSUBS 0.007771f
C1070 B.n913 VSUBS 0.007771f
C1071 B.n914 VSUBS 0.007771f
C1072 B.n915 VSUBS 0.007771f
C1073 B.n916 VSUBS 0.007771f
C1074 B.n917 VSUBS 0.007771f
C1075 B.n918 VSUBS 0.018274f
C1076 B.n919 VSUBS 0.018274f
C1077 B.n920 VSUBS 0.017611f
C1078 B.n921 VSUBS 0.007771f
C1079 B.n922 VSUBS 0.007771f
C1080 B.n923 VSUBS 0.007771f
C1081 B.n924 VSUBS 0.007771f
C1082 B.n925 VSUBS 0.007771f
C1083 B.n926 VSUBS 0.007771f
C1084 B.n927 VSUBS 0.007771f
C1085 B.n928 VSUBS 0.007771f
C1086 B.n929 VSUBS 0.007771f
C1087 B.n930 VSUBS 0.007771f
C1088 B.n931 VSUBS 0.007771f
C1089 B.n932 VSUBS 0.007771f
C1090 B.n933 VSUBS 0.007771f
C1091 B.n934 VSUBS 0.007771f
C1092 B.n935 VSUBS 0.007771f
C1093 B.n936 VSUBS 0.007771f
C1094 B.n937 VSUBS 0.007771f
C1095 B.n938 VSUBS 0.007771f
C1096 B.n939 VSUBS 0.007771f
C1097 B.n940 VSUBS 0.007771f
C1098 B.n941 VSUBS 0.007771f
C1099 B.n942 VSUBS 0.007771f
C1100 B.n943 VSUBS 0.007771f
C1101 B.n944 VSUBS 0.007771f
C1102 B.n945 VSUBS 0.007771f
C1103 B.n946 VSUBS 0.007771f
C1104 B.n947 VSUBS 0.007771f
C1105 B.n948 VSUBS 0.007771f
C1106 B.n949 VSUBS 0.007771f
C1107 B.n950 VSUBS 0.007771f
C1108 B.n951 VSUBS 0.007771f
C1109 B.n952 VSUBS 0.007771f
C1110 B.n953 VSUBS 0.007771f
C1111 B.n954 VSUBS 0.007771f
C1112 B.n955 VSUBS 0.007771f
C1113 B.n956 VSUBS 0.007771f
C1114 B.n957 VSUBS 0.007771f
C1115 B.n958 VSUBS 0.007771f
C1116 B.n959 VSUBS 0.007771f
C1117 B.n960 VSUBS 0.007771f
C1118 B.n961 VSUBS 0.007771f
C1119 B.n962 VSUBS 0.007771f
C1120 B.n963 VSUBS 0.007771f
C1121 B.n964 VSUBS 0.007771f
C1122 B.n965 VSUBS 0.007771f
C1123 B.n966 VSUBS 0.007771f
C1124 B.n967 VSUBS 0.007771f
C1125 B.n968 VSUBS 0.007771f
C1126 B.n969 VSUBS 0.007771f
C1127 B.n970 VSUBS 0.007771f
C1128 B.n971 VSUBS 0.007771f
C1129 B.n972 VSUBS 0.007771f
C1130 B.n973 VSUBS 0.007771f
C1131 B.n974 VSUBS 0.007771f
C1132 B.n975 VSUBS 0.007771f
C1133 B.n976 VSUBS 0.007771f
C1134 B.n977 VSUBS 0.007771f
C1135 B.n978 VSUBS 0.007771f
C1136 B.n979 VSUBS 0.007771f
C1137 B.n980 VSUBS 0.007771f
C1138 B.n981 VSUBS 0.007771f
C1139 B.n982 VSUBS 0.007771f
C1140 B.n983 VSUBS 0.007771f
C1141 B.n984 VSUBS 0.007771f
C1142 B.n985 VSUBS 0.007771f
C1143 B.n986 VSUBS 0.007771f
C1144 B.n987 VSUBS 0.007771f
C1145 B.n988 VSUBS 0.007771f
C1146 B.n989 VSUBS 0.007771f
C1147 B.n990 VSUBS 0.007771f
C1148 B.n991 VSUBS 0.007771f
C1149 B.n992 VSUBS 0.007771f
C1150 B.n993 VSUBS 0.007771f
C1151 B.n994 VSUBS 0.007771f
C1152 B.n995 VSUBS 0.007771f
C1153 B.n996 VSUBS 0.007771f
C1154 B.n997 VSUBS 0.007771f
C1155 B.n998 VSUBS 0.007771f
C1156 B.n999 VSUBS 0.007771f
C1157 B.n1000 VSUBS 0.007771f
C1158 B.n1001 VSUBS 0.007771f
C1159 B.n1002 VSUBS 0.007771f
C1160 B.n1003 VSUBS 0.007771f
C1161 B.n1004 VSUBS 0.007771f
C1162 B.n1005 VSUBS 0.007771f
C1163 B.n1006 VSUBS 0.007771f
C1164 B.n1007 VSUBS 0.007771f
C1165 B.n1008 VSUBS 0.007771f
C1166 B.n1009 VSUBS 0.007771f
C1167 B.n1010 VSUBS 0.007771f
C1168 B.n1011 VSUBS 0.007771f
C1169 B.n1012 VSUBS 0.007771f
C1170 B.n1013 VSUBS 0.007771f
C1171 B.n1014 VSUBS 0.007771f
C1172 B.n1015 VSUBS 0.007771f
C1173 B.n1016 VSUBS 0.007771f
C1174 B.n1017 VSUBS 0.007771f
C1175 B.n1018 VSUBS 0.007771f
C1176 B.n1019 VSUBS 0.007771f
C1177 B.n1020 VSUBS 0.007771f
C1178 B.n1021 VSUBS 0.007771f
C1179 B.n1022 VSUBS 0.007771f
C1180 B.n1023 VSUBS 0.007771f
C1181 B.n1024 VSUBS 0.007771f
C1182 B.n1025 VSUBS 0.007771f
C1183 B.n1026 VSUBS 0.007771f
C1184 B.n1027 VSUBS 0.017597f
C1185 VTAIL.t8 VSUBS 0.300255f
C1186 VTAIL.t15 VSUBS 0.300255f
C1187 VTAIL.n0 VSUBS 2.30664f
C1188 VTAIL.n1 VSUBS 0.883111f
C1189 VTAIL.t14 VSUBS 3.02093f
C1190 VTAIL.n2 VSUBS 1.02106f
C1191 VTAIL.t6 VSUBS 3.02093f
C1192 VTAIL.n3 VSUBS 1.02106f
C1193 VTAIL.t2 VSUBS 0.300255f
C1194 VTAIL.t5 VSUBS 0.300255f
C1195 VTAIL.n4 VSUBS 2.30664f
C1196 VTAIL.n5 VSUBS 1.17666f
C1197 VTAIL.t1 VSUBS 3.02093f
C1198 VTAIL.n6 VSUBS 2.67827f
C1199 VTAIL.t9 VSUBS 3.02094f
C1200 VTAIL.n7 VSUBS 2.67827f
C1201 VTAIL.t10 VSUBS 0.300255f
C1202 VTAIL.t12 VSUBS 0.300255f
C1203 VTAIL.n8 VSUBS 2.30665f
C1204 VTAIL.n9 VSUBS 1.17665f
C1205 VTAIL.t13 VSUBS 3.02094f
C1206 VTAIL.n10 VSUBS 1.02105f
C1207 VTAIL.t7 VSUBS 3.02094f
C1208 VTAIL.n11 VSUBS 1.02105f
C1209 VTAIL.t4 VSUBS 0.300255f
C1210 VTAIL.t3 VSUBS 0.300255f
C1211 VTAIL.n12 VSUBS 2.30665f
C1212 VTAIL.n13 VSUBS 1.17665f
C1213 VTAIL.t0 VSUBS 3.02093f
C1214 VTAIL.n14 VSUBS 2.67827f
C1215 VTAIL.t11 VSUBS 3.02093f
C1216 VTAIL.n15 VSUBS 2.67356f
C1217 VDD2.t6 VSUBS 0.386849f
C1218 VDD2.t2 VSUBS 0.386849f
C1219 VDD2.n0 VSUBS 3.18087f
C1220 VDD2.t7 VSUBS 0.386849f
C1221 VDD2.t1 VSUBS 0.386849f
C1222 VDD2.n1 VSUBS 3.18087f
C1223 VDD2.n2 VSUBS 6.18604f
C1224 VDD2.t3 VSUBS 0.386849f
C1225 VDD2.t0 VSUBS 0.386849f
C1226 VDD2.n3 VSUBS 3.15221f
C1227 VDD2.n4 VSUBS 5.07418f
C1228 VDD2.t4 VSUBS 0.386849f
C1229 VDD2.t5 VSUBS 0.386849f
C1230 VDD2.n5 VSUBS 3.1808f
C1231 VN.n0 VSUBS 0.040705f
C1232 VN.t4 VSUBS 3.5308f
C1233 VN.n1 VSUBS 0.040332f
C1234 VN.n2 VSUBS 0.02164f
C1235 VN.n3 VSUBS 0.040332f
C1236 VN.n4 VSUBS 0.02164f
C1237 VN.t0 VSUBS 3.5308f
C1238 VN.n5 VSUBS 0.040332f
C1239 VN.n6 VSUBS 0.02164f
C1240 VN.n7 VSUBS 0.040332f
C1241 VN.n8 VSUBS 0.288136f
C1242 VN.t7 VSUBS 3.5308f
C1243 VN.t1 VSUBS 3.8914f
C1244 VN.n9 VSUBS 1.2362f
C1245 VN.n10 VSUBS 1.29767f
C1246 VN.n11 VSUBS 0.025795f
C1247 VN.n12 VSUBS 0.040332f
C1248 VN.n13 VSUBS 0.02164f
C1249 VN.n14 VSUBS 0.02164f
C1250 VN.n15 VSUBS 0.02164f
C1251 VN.n16 VSUBS 0.043009f
C1252 VN.n17 VSUBS 0.017494f
C1253 VN.n18 VSUBS 0.043009f
C1254 VN.n19 VSUBS 0.02164f
C1255 VN.n20 VSUBS 0.02164f
C1256 VN.n21 VSUBS 0.02164f
C1257 VN.n22 VSUBS 0.040332f
C1258 VN.n23 VSUBS 0.025795f
C1259 VN.n24 VSUBS 1.22339f
C1260 VN.n25 VSUBS 0.034954f
C1261 VN.n26 VSUBS 0.02164f
C1262 VN.n27 VSUBS 0.02164f
C1263 VN.n28 VSUBS 0.02164f
C1264 VN.n29 VSUBS 0.040332f
C1265 VN.n30 VSUBS 0.032797f
C1266 VN.n31 VSUBS 0.030385f
C1267 VN.n32 VSUBS 0.02164f
C1268 VN.n33 VSUBS 0.02164f
C1269 VN.n34 VSUBS 0.02164f
C1270 VN.n35 VSUBS 0.040332f
C1271 VN.n36 VSUBS 0.036548f
C1272 VN.n37 VSUBS 1.31709f
C1273 VN.n38 VSUBS 0.06914f
C1274 VN.n39 VSUBS 0.040705f
C1275 VN.t6 VSUBS 3.5308f
C1276 VN.n40 VSUBS 0.040332f
C1277 VN.n41 VSUBS 0.02164f
C1278 VN.n42 VSUBS 0.040332f
C1279 VN.n43 VSUBS 0.02164f
C1280 VN.t5 VSUBS 3.5308f
C1281 VN.n44 VSUBS 0.040332f
C1282 VN.n45 VSUBS 0.02164f
C1283 VN.n46 VSUBS 0.040332f
C1284 VN.n47 VSUBS 0.288136f
C1285 VN.t3 VSUBS 3.5308f
C1286 VN.t2 VSUBS 3.8914f
C1287 VN.n48 VSUBS 1.2362f
C1288 VN.n49 VSUBS 1.29767f
C1289 VN.n50 VSUBS 0.025795f
C1290 VN.n51 VSUBS 0.040332f
C1291 VN.n52 VSUBS 0.02164f
C1292 VN.n53 VSUBS 0.02164f
C1293 VN.n54 VSUBS 0.02164f
C1294 VN.n55 VSUBS 0.043009f
C1295 VN.n56 VSUBS 0.017494f
C1296 VN.n57 VSUBS 0.043009f
C1297 VN.n58 VSUBS 0.02164f
C1298 VN.n59 VSUBS 0.02164f
C1299 VN.n60 VSUBS 0.02164f
C1300 VN.n61 VSUBS 0.040332f
C1301 VN.n62 VSUBS 0.025795f
C1302 VN.n63 VSUBS 1.22339f
C1303 VN.n64 VSUBS 0.034954f
C1304 VN.n65 VSUBS 0.02164f
C1305 VN.n66 VSUBS 0.02164f
C1306 VN.n67 VSUBS 0.02164f
C1307 VN.n68 VSUBS 0.040332f
C1308 VN.n69 VSUBS 0.032797f
C1309 VN.n70 VSUBS 0.030385f
C1310 VN.n71 VSUBS 0.02164f
C1311 VN.n72 VSUBS 0.02164f
C1312 VN.n73 VSUBS 0.02164f
C1313 VN.n74 VSUBS 0.040332f
C1314 VN.n75 VSUBS 0.036548f
C1315 VN.n76 VSUBS 1.31709f
C1316 VN.n77 VSUBS 1.60921f
.ends

