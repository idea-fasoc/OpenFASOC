* NGSPICE file created from diff_pair_sample_1460.ext - technology: sky130A

.subckt diff_pair_sample_1460 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VN.t0 VDD2.t4 B.t7 sky130_fd_pr__nfet_01v8 ad=1.023 pd=6.53 as=1.023 ps=6.53 w=6.2 l=3.07
X1 VDD1.t7 VP.t0 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.023 pd=6.53 as=2.418 ps=13.18 w=6.2 l=3.07
X2 B.t21 B.t19 B.t20 B.t13 sky130_fd_pr__nfet_01v8 ad=2.418 pd=13.18 as=0 ps=0 w=6.2 l=3.07
X3 VTAIL.t5 VP.t1 VDD1.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=2.418 pd=13.18 as=1.023 ps=6.53 w=6.2 l=3.07
X4 B.t18 B.t16 B.t17 B.t9 sky130_fd_pr__nfet_01v8 ad=2.418 pd=13.18 as=0 ps=0 w=6.2 l=3.07
X5 VDD2.t5 VN.t1 VTAIL.t14 B.t1 sky130_fd_pr__nfet_01v8 ad=1.023 pd=6.53 as=1.023 ps=6.53 w=6.2 l=3.07
X6 VTAIL.t13 VN.t2 VDD2.t2 B.t5 sky130_fd_pr__nfet_01v8 ad=2.418 pd=13.18 as=1.023 ps=6.53 w=6.2 l=3.07
X7 VDD2.t6 VN.t3 VTAIL.t12 B.t0 sky130_fd_pr__nfet_01v8 ad=1.023 pd=6.53 as=2.418 ps=13.18 w=6.2 l=3.07
X8 VTAIL.t11 VN.t4 VDD2.t7 B.t6 sky130_fd_pr__nfet_01v8 ad=2.418 pd=13.18 as=1.023 ps=6.53 w=6.2 l=3.07
X9 VDD1.t5 VP.t2 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.023 pd=6.53 as=1.023 ps=6.53 w=6.2 l=3.07
X10 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=2.418 pd=13.18 as=0 ps=0 w=6.2 l=3.07
X11 VDD2.t0 VN.t5 VTAIL.t10 B.t2 sky130_fd_pr__nfet_01v8 ad=1.023 pd=6.53 as=1.023 ps=6.53 w=6.2 l=3.07
X12 VDD1.t4 VP.t3 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.023 pd=6.53 as=1.023 ps=6.53 w=6.2 l=3.07
X13 VDD2.t3 VN.t6 VTAIL.t9 B.t3 sky130_fd_pr__nfet_01v8 ad=1.023 pd=6.53 as=2.418 ps=13.18 w=6.2 l=3.07
X14 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=2.418 pd=13.18 as=0 ps=0 w=6.2 l=3.07
X15 VTAIL.t4 VP.t4 VDD1.t3 B.t4 sky130_fd_pr__nfet_01v8 ad=1.023 pd=6.53 as=1.023 ps=6.53 w=6.2 l=3.07
X16 VDD1.t2 VP.t5 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.023 pd=6.53 as=2.418 ps=13.18 w=6.2 l=3.07
X17 VTAIL.t7 VP.t6 VDD1.t1 B.t7 sky130_fd_pr__nfet_01v8 ad=1.023 pd=6.53 as=1.023 ps=6.53 w=6.2 l=3.07
X18 VTAIL.t8 VN.t7 VDD2.t1 B.t4 sky130_fd_pr__nfet_01v8 ad=1.023 pd=6.53 as=1.023 ps=6.53 w=6.2 l=3.07
X19 VTAIL.t6 VP.t7 VDD1.t0 B.t6 sky130_fd_pr__nfet_01v8 ad=2.418 pd=13.18 as=1.023 ps=6.53 w=6.2 l=3.07
R0 VN.n60 VN.n59 161.3
R1 VN.n58 VN.n32 161.3
R2 VN.n57 VN.n56 161.3
R3 VN.n55 VN.n33 161.3
R4 VN.n54 VN.n53 161.3
R5 VN.n52 VN.n34 161.3
R6 VN.n51 VN.n50 161.3
R7 VN.n49 VN.n48 161.3
R8 VN.n47 VN.n36 161.3
R9 VN.n46 VN.n45 161.3
R10 VN.n44 VN.n37 161.3
R11 VN.n43 VN.n42 161.3
R12 VN.n41 VN.n38 161.3
R13 VN.n29 VN.n28 161.3
R14 VN.n27 VN.n1 161.3
R15 VN.n26 VN.n25 161.3
R16 VN.n24 VN.n2 161.3
R17 VN.n23 VN.n22 161.3
R18 VN.n21 VN.n3 161.3
R19 VN.n20 VN.n19 161.3
R20 VN.n18 VN.n17 161.3
R21 VN.n16 VN.n5 161.3
R22 VN.n15 VN.n14 161.3
R23 VN.n13 VN.n6 161.3
R24 VN.n12 VN.n11 161.3
R25 VN.n10 VN.n7 161.3
R26 VN.n39 VN.t6 82.0222
R27 VN.n8 VN.t2 82.0222
R28 VN.n30 VN.n0 73.0313
R29 VN.n61 VN.n31 73.0313
R30 VN.n15 VN.n6 56.5617
R31 VN.n46 VN.n37 56.5617
R32 VN.n26 VN.n2 55.1086
R33 VN.n57 VN.n33 55.1086
R34 VN.n40 VN.n39 51.9074
R35 VN.n9 VN.n8 51.9074
R36 VN VN.n61 48.9603
R37 VN.n9 VN.t1 48.6715
R38 VN.n4 VN.t7 48.6715
R39 VN.n0 VN.t3 48.6715
R40 VN.n40 VN.t0 48.6715
R41 VN.n35 VN.t5 48.6715
R42 VN.n31 VN.t4 48.6715
R43 VN.n22 VN.n2 26.0455
R44 VN.n53 VN.n33 26.0455
R45 VN.n11 VN.n10 24.5923
R46 VN.n11 VN.n6 24.5923
R47 VN.n16 VN.n15 24.5923
R48 VN.n17 VN.n16 24.5923
R49 VN.n21 VN.n20 24.5923
R50 VN.n22 VN.n21 24.5923
R51 VN.n27 VN.n26 24.5923
R52 VN.n28 VN.n27 24.5923
R53 VN.n42 VN.n37 24.5923
R54 VN.n42 VN.n41 24.5923
R55 VN.n53 VN.n52 24.5923
R56 VN.n52 VN.n51 24.5923
R57 VN.n48 VN.n47 24.5923
R58 VN.n47 VN.n46 24.5923
R59 VN.n59 VN.n58 24.5923
R60 VN.n58 VN.n57 24.5923
R61 VN.n10 VN.n9 22.1332
R62 VN.n17 VN.n4 22.1332
R63 VN.n41 VN.n40 22.1332
R64 VN.n48 VN.n35 22.1332
R65 VN.n28 VN.n0 17.2148
R66 VN.n59 VN.n31 17.2148
R67 VN.n39 VN.n38 4.03539
R68 VN.n8 VN.n7 4.03539
R69 VN.n20 VN.n4 2.45968
R70 VN.n51 VN.n35 2.45968
R71 VN.n61 VN.n60 0.354861
R72 VN.n30 VN.n29 0.354861
R73 VN VN.n30 0.267071
R74 VN.n60 VN.n32 0.189894
R75 VN.n56 VN.n32 0.189894
R76 VN.n56 VN.n55 0.189894
R77 VN.n55 VN.n54 0.189894
R78 VN.n54 VN.n34 0.189894
R79 VN.n50 VN.n34 0.189894
R80 VN.n50 VN.n49 0.189894
R81 VN.n49 VN.n36 0.189894
R82 VN.n45 VN.n36 0.189894
R83 VN.n45 VN.n44 0.189894
R84 VN.n44 VN.n43 0.189894
R85 VN.n43 VN.n38 0.189894
R86 VN.n12 VN.n7 0.189894
R87 VN.n13 VN.n12 0.189894
R88 VN.n14 VN.n13 0.189894
R89 VN.n14 VN.n5 0.189894
R90 VN.n18 VN.n5 0.189894
R91 VN.n19 VN.n18 0.189894
R92 VN.n19 VN.n3 0.189894
R93 VN.n23 VN.n3 0.189894
R94 VN.n24 VN.n23 0.189894
R95 VN.n25 VN.n24 0.189894
R96 VN.n25 VN.n1 0.189894
R97 VN.n29 VN.n1 0.189894
R98 VDD2.n2 VDD2.n1 71.1509
R99 VDD2.n2 VDD2.n0 71.1509
R100 VDD2 VDD2.n5 71.1472
R101 VDD2.n4 VDD2.n3 69.7408
R102 VDD2.n4 VDD2.n2 42.2498
R103 VDD2.n5 VDD2.t4 3.19405
R104 VDD2.n5 VDD2.t3 3.19405
R105 VDD2.n3 VDD2.t7 3.19405
R106 VDD2.n3 VDD2.t0 3.19405
R107 VDD2.n1 VDD2.t1 3.19405
R108 VDD2.n1 VDD2.t6 3.19405
R109 VDD2.n0 VDD2.t2 3.19405
R110 VDD2.n0 VDD2.t5 3.19405
R111 VDD2 VDD2.n4 1.52421
R112 VTAIL.n11 VTAIL.t5 56.2556
R113 VTAIL.n10 VTAIL.t9 56.2556
R114 VTAIL.n7 VTAIL.t11 56.2556
R115 VTAIL.n14 VTAIL.t0 56.2547
R116 VTAIL.n15 VTAIL.t12 56.2546
R117 VTAIL.n2 VTAIL.t13 56.2546
R118 VTAIL.n3 VTAIL.t3 56.2546
R119 VTAIL.n6 VTAIL.t6 56.2546
R120 VTAIL.n13 VTAIL.n12 53.062
R121 VTAIL.n9 VTAIL.n8 53.062
R122 VTAIL.n1 VTAIL.n0 53.0619
R123 VTAIL.n5 VTAIL.n4 53.0619
R124 VTAIL.n15 VTAIL.n14 20.6427
R125 VTAIL.n7 VTAIL.n6 20.6427
R126 VTAIL.n0 VTAIL.t14 3.19405
R127 VTAIL.n0 VTAIL.t8 3.19405
R128 VTAIL.n4 VTAIL.t2 3.19405
R129 VTAIL.n4 VTAIL.t7 3.19405
R130 VTAIL.n12 VTAIL.t1 3.19405
R131 VTAIL.n12 VTAIL.t4 3.19405
R132 VTAIL.n8 VTAIL.t10 3.19405
R133 VTAIL.n8 VTAIL.t15 3.19405
R134 VTAIL.n9 VTAIL.n7 2.93153
R135 VTAIL.n10 VTAIL.n9 2.93153
R136 VTAIL.n13 VTAIL.n11 2.93153
R137 VTAIL.n14 VTAIL.n13 2.93153
R138 VTAIL.n6 VTAIL.n5 2.93153
R139 VTAIL.n5 VTAIL.n3 2.93153
R140 VTAIL.n2 VTAIL.n1 2.93153
R141 VTAIL VTAIL.n15 2.87334
R142 VTAIL.n11 VTAIL.n10 0.470328
R143 VTAIL.n3 VTAIL.n2 0.470328
R144 VTAIL VTAIL.n1 0.0586897
R145 B.n656 B.n141 585
R146 B.n141 B.n106 585
R147 B.n658 B.n657 585
R148 B.n660 B.n140 585
R149 B.n663 B.n662 585
R150 B.n664 B.n139 585
R151 B.n666 B.n665 585
R152 B.n668 B.n138 585
R153 B.n671 B.n670 585
R154 B.n672 B.n137 585
R155 B.n674 B.n673 585
R156 B.n676 B.n136 585
R157 B.n679 B.n678 585
R158 B.n680 B.n135 585
R159 B.n682 B.n681 585
R160 B.n684 B.n134 585
R161 B.n687 B.n686 585
R162 B.n688 B.n133 585
R163 B.n690 B.n689 585
R164 B.n692 B.n132 585
R165 B.n695 B.n694 585
R166 B.n696 B.n131 585
R167 B.n698 B.n697 585
R168 B.n700 B.n130 585
R169 B.n702 B.n701 585
R170 B.n704 B.n703 585
R171 B.n707 B.n706 585
R172 B.n708 B.n125 585
R173 B.n710 B.n709 585
R174 B.n712 B.n124 585
R175 B.n715 B.n714 585
R176 B.n716 B.n123 585
R177 B.n718 B.n717 585
R178 B.n720 B.n122 585
R179 B.n723 B.n722 585
R180 B.n725 B.n119 585
R181 B.n727 B.n726 585
R182 B.n729 B.n118 585
R183 B.n732 B.n731 585
R184 B.n733 B.n117 585
R185 B.n735 B.n734 585
R186 B.n737 B.n116 585
R187 B.n740 B.n739 585
R188 B.n741 B.n115 585
R189 B.n743 B.n742 585
R190 B.n745 B.n114 585
R191 B.n748 B.n747 585
R192 B.n749 B.n113 585
R193 B.n751 B.n750 585
R194 B.n753 B.n112 585
R195 B.n756 B.n755 585
R196 B.n757 B.n111 585
R197 B.n759 B.n758 585
R198 B.n761 B.n110 585
R199 B.n764 B.n763 585
R200 B.n765 B.n109 585
R201 B.n767 B.n766 585
R202 B.n769 B.n108 585
R203 B.n772 B.n771 585
R204 B.n773 B.n107 585
R205 B.n655 B.n105 585
R206 B.n776 B.n105 585
R207 B.n654 B.n104 585
R208 B.n777 B.n104 585
R209 B.n653 B.n103 585
R210 B.n778 B.n103 585
R211 B.n652 B.n651 585
R212 B.n651 B.n99 585
R213 B.n650 B.n98 585
R214 B.n784 B.n98 585
R215 B.n649 B.n97 585
R216 B.n785 B.n97 585
R217 B.n648 B.n96 585
R218 B.n786 B.n96 585
R219 B.n647 B.n646 585
R220 B.n646 B.n92 585
R221 B.n645 B.n91 585
R222 B.n792 B.n91 585
R223 B.n644 B.n90 585
R224 B.n793 B.n90 585
R225 B.n643 B.n89 585
R226 B.n794 B.n89 585
R227 B.n642 B.n641 585
R228 B.n641 B.n85 585
R229 B.n640 B.n84 585
R230 B.n800 B.n84 585
R231 B.n639 B.n83 585
R232 B.n801 B.n83 585
R233 B.n638 B.n82 585
R234 B.n802 B.n82 585
R235 B.n637 B.n636 585
R236 B.n636 B.n78 585
R237 B.n635 B.n77 585
R238 B.n808 B.n77 585
R239 B.n634 B.n76 585
R240 B.n809 B.n76 585
R241 B.n633 B.n75 585
R242 B.n810 B.n75 585
R243 B.n632 B.n631 585
R244 B.n631 B.n71 585
R245 B.n630 B.n70 585
R246 B.n816 B.n70 585
R247 B.n629 B.n69 585
R248 B.n817 B.n69 585
R249 B.n628 B.n68 585
R250 B.n818 B.n68 585
R251 B.n627 B.n626 585
R252 B.n626 B.n64 585
R253 B.n625 B.n63 585
R254 B.n824 B.n63 585
R255 B.n624 B.n62 585
R256 B.n825 B.n62 585
R257 B.n623 B.n61 585
R258 B.n826 B.n61 585
R259 B.n622 B.n621 585
R260 B.n621 B.n57 585
R261 B.n620 B.n56 585
R262 B.n832 B.n56 585
R263 B.n619 B.n55 585
R264 B.n833 B.n55 585
R265 B.n618 B.n54 585
R266 B.n834 B.n54 585
R267 B.n617 B.n616 585
R268 B.n616 B.n53 585
R269 B.n615 B.n49 585
R270 B.n840 B.n49 585
R271 B.n614 B.n48 585
R272 B.n841 B.n48 585
R273 B.n613 B.n47 585
R274 B.n842 B.n47 585
R275 B.n612 B.n611 585
R276 B.n611 B.n43 585
R277 B.n610 B.n42 585
R278 B.n848 B.n42 585
R279 B.n609 B.n41 585
R280 B.n849 B.n41 585
R281 B.n608 B.n40 585
R282 B.n850 B.n40 585
R283 B.n607 B.n606 585
R284 B.n606 B.n36 585
R285 B.n605 B.n35 585
R286 B.n856 B.n35 585
R287 B.n604 B.n34 585
R288 B.n857 B.n34 585
R289 B.n603 B.n33 585
R290 B.n858 B.n33 585
R291 B.n602 B.n601 585
R292 B.n601 B.n29 585
R293 B.n600 B.n28 585
R294 B.n864 B.n28 585
R295 B.n599 B.n27 585
R296 B.n865 B.n27 585
R297 B.n598 B.n26 585
R298 B.n866 B.n26 585
R299 B.n597 B.n596 585
R300 B.n596 B.n22 585
R301 B.n595 B.n21 585
R302 B.n872 B.n21 585
R303 B.n594 B.n20 585
R304 B.n873 B.n20 585
R305 B.n593 B.n19 585
R306 B.n874 B.n19 585
R307 B.n592 B.n591 585
R308 B.n591 B.n18 585
R309 B.n590 B.n14 585
R310 B.n880 B.n14 585
R311 B.n589 B.n13 585
R312 B.n881 B.n13 585
R313 B.n588 B.n12 585
R314 B.n882 B.n12 585
R315 B.n587 B.n586 585
R316 B.n586 B.n8 585
R317 B.n585 B.n7 585
R318 B.n888 B.n7 585
R319 B.n584 B.n6 585
R320 B.n889 B.n6 585
R321 B.n583 B.n5 585
R322 B.n890 B.n5 585
R323 B.n582 B.n581 585
R324 B.n581 B.n4 585
R325 B.n580 B.n142 585
R326 B.n580 B.n579 585
R327 B.n570 B.n143 585
R328 B.n144 B.n143 585
R329 B.n572 B.n571 585
R330 B.n573 B.n572 585
R331 B.n569 B.n149 585
R332 B.n149 B.n148 585
R333 B.n568 B.n567 585
R334 B.n567 B.n566 585
R335 B.n151 B.n150 585
R336 B.n559 B.n151 585
R337 B.n558 B.n557 585
R338 B.n560 B.n558 585
R339 B.n556 B.n156 585
R340 B.n156 B.n155 585
R341 B.n555 B.n554 585
R342 B.n554 B.n553 585
R343 B.n158 B.n157 585
R344 B.n159 B.n158 585
R345 B.n546 B.n545 585
R346 B.n547 B.n546 585
R347 B.n544 B.n164 585
R348 B.n164 B.n163 585
R349 B.n543 B.n542 585
R350 B.n542 B.n541 585
R351 B.n166 B.n165 585
R352 B.n167 B.n166 585
R353 B.n534 B.n533 585
R354 B.n535 B.n534 585
R355 B.n532 B.n171 585
R356 B.n175 B.n171 585
R357 B.n531 B.n530 585
R358 B.n530 B.n529 585
R359 B.n173 B.n172 585
R360 B.n174 B.n173 585
R361 B.n522 B.n521 585
R362 B.n523 B.n522 585
R363 B.n520 B.n180 585
R364 B.n180 B.n179 585
R365 B.n519 B.n518 585
R366 B.n518 B.n517 585
R367 B.n182 B.n181 585
R368 B.n183 B.n182 585
R369 B.n510 B.n509 585
R370 B.n511 B.n510 585
R371 B.n508 B.n188 585
R372 B.n188 B.n187 585
R373 B.n507 B.n506 585
R374 B.n506 B.n505 585
R375 B.n190 B.n189 585
R376 B.n498 B.n190 585
R377 B.n497 B.n496 585
R378 B.n499 B.n497 585
R379 B.n495 B.n195 585
R380 B.n195 B.n194 585
R381 B.n494 B.n493 585
R382 B.n493 B.n492 585
R383 B.n197 B.n196 585
R384 B.n198 B.n197 585
R385 B.n485 B.n484 585
R386 B.n486 B.n485 585
R387 B.n483 B.n203 585
R388 B.n203 B.n202 585
R389 B.n482 B.n481 585
R390 B.n481 B.n480 585
R391 B.n205 B.n204 585
R392 B.n206 B.n205 585
R393 B.n473 B.n472 585
R394 B.n474 B.n473 585
R395 B.n471 B.n210 585
R396 B.n214 B.n210 585
R397 B.n470 B.n469 585
R398 B.n469 B.n468 585
R399 B.n212 B.n211 585
R400 B.n213 B.n212 585
R401 B.n461 B.n460 585
R402 B.n462 B.n461 585
R403 B.n459 B.n219 585
R404 B.n219 B.n218 585
R405 B.n458 B.n457 585
R406 B.n457 B.n456 585
R407 B.n221 B.n220 585
R408 B.n222 B.n221 585
R409 B.n449 B.n448 585
R410 B.n450 B.n449 585
R411 B.n447 B.n227 585
R412 B.n227 B.n226 585
R413 B.n446 B.n445 585
R414 B.n445 B.n444 585
R415 B.n229 B.n228 585
R416 B.n230 B.n229 585
R417 B.n437 B.n436 585
R418 B.n438 B.n437 585
R419 B.n435 B.n235 585
R420 B.n235 B.n234 585
R421 B.n434 B.n433 585
R422 B.n433 B.n432 585
R423 B.n237 B.n236 585
R424 B.n238 B.n237 585
R425 B.n425 B.n424 585
R426 B.n426 B.n425 585
R427 B.n423 B.n243 585
R428 B.n243 B.n242 585
R429 B.n422 B.n421 585
R430 B.n421 B.n420 585
R431 B.n245 B.n244 585
R432 B.n246 B.n245 585
R433 B.n413 B.n412 585
R434 B.n414 B.n413 585
R435 B.n411 B.n251 585
R436 B.n251 B.n250 585
R437 B.n410 B.n409 585
R438 B.n409 B.n408 585
R439 B.n405 B.n255 585
R440 B.n404 B.n403 585
R441 B.n401 B.n256 585
R442 B.n401 B.n254 585
R443 B.n400 B.n399 585
R444 B.n398 B.n397 585
R445 B.n396 B.n258 585
R446 B.n394 B.n393 585
R447 B.n392 B.n259 585
R448 B.n391 B.n390 585
R449 B.n388 B.n260 585
R450 B.n386 B.n385 585
R451 B.n384 B.n261 585
R452 B.n383 B.n382 585
R453 B.n380 B.n262 585
R454 B.n378 B.n377 585
R455 B.n376 B.n263 585
R456 B.n375 B.n374 585
R457 B.n372 B.n264 585
R458 B.n370 B.n369 585
R459 B.n368 B.n265 585
R460 B.n367 B.n366 585
R461 B.n364 B.n266 585
R462 B.n362 B.n361 585
R463 B.n360 B.n267 585
R464 B.n359 B.n358 585
R465 B.n356 B.n355 585
R466 B.n354 B.n353 585
R467 B.n352 B.n272 585
R468 B.n350 B.n349 585
R469 B.n348 B.n273 585
R470 B.n347 B.n346 585
R471 B.n344 B.n274 585
R472 B.n342 B.n341 585
R473 B.n340 B.n275 585
R474 B.n338 B.n337 585
R475 B.n335 B.n278 585
R476 B.n333 B.n332 585
R477 B.n331 B.n279 585
R478 B.n330 B.n329 585
R479 B.n327 B.n280 585
R480 B.n325 B.n324 585
R481 B.n323 B.n281 585
R482 B.n322 B.n321 585
R483 B.n319 B.n282 585
R484 B.n317 B.n316 585
R485 B.n315 B.n283 585
R486 B.n314 B.n313 585
R487 B.n311 B.n284 585
R488 B.n309 B.n308 585
R489 B.n307 B.n285 585
R490 B.n306 B.n305 585
R491 B.n303 B.n286 585
R492 B.n301 B.n300 585
R493 B.n299 B.n287 585
R494 B.n298 B.n297 585
R495 B.n295 B.n288 585
R496 B.n293 B.n292 585
R497 B.n291 B.n290 585
R498 B.n253 B.n252 585
R499 B.n407 B.n406 585
R500 B.n408 B.n407 585
R501 B.n249 B.n248 585
R502 B.n250 B.n249 585
R503 B.n416 B.n415 585
R504 B.n415 B.n414 585
R505 B.n417 B.n247 585
R506 B.n247 B.n246 585
R507 B.n419 B.n418 585
R508 B.n420 B.n419 585
R509 B.n241 B.n240 585
R510 B.n242 B.n241 585
R511 B.n428 B.n427 585
R512 B.n427 B.n426 585
R513 B.n429 B.n239 585
R514 B.n239 B.n238 585
R515 B.n431 B.n430 585
R516 B.n432 B.n431 585
R517 B.n233 B.n232 585
R518 B.n234 B.n233 585
R519 B.n440 B.n439 585
R520 B.n439 B.n438 585
R521 B.n441 B.n231 585
R522 B.n231 B.n230 585
R523 B.n443 B.n442 585
R524 B.n444 B.n443 585
R525 B.n225 B.n224 585
R526 B.n226 B.n225 585
R527 B.n452 B.n451 585
R528 B.n451 B.n450 585
R529 B.n453 B.n223 585
R530 B.n223 B.n222 585
R531 B.n455 B.n454 585
R532 B.n456 B.n455 585
R533 B.n217 B.n216 585
R534 B.n218 B.n217 585
R535 B.n464 B.n463 585
R536 B.n463 B.n462 585
R537 B.n465 B.n215 585
R538 B.n215 B.n213 585
R539 B.n467 B.n466 585
R540 B.n468 B.n467 585
R541 B.n209 B.n208 585
R542 B.n214 B.n209 585
R543 B.n476 B.n475 585
R544 B.n475 B.n474 585
R545 B.n477 B.n207 585
R546 B.n207 B.n206 585
R547 B.n479 B.n478 585
R548 B.n480 B.n479 585
R549 B.n201 B.n200 585
R550 B.n202 B.n201 585
R551 B.n488 B.n487 585
R552 B.n487 B.n486 585
R553 B.n489 B.n199 585
R554 B.n199 B.n198 585
R555 B.n491 B.n490 585
R556 B.n492 B.n491 585
R557 B.n193 B.n192 585
R558 B.n194 B.n193 585
R559 B.n501 B.n500 585
R560 B.n500 B.n499 585
R561 B.n502 B.n191 585
R562 B.n498 B.n191 585
R563 B.n504 B.n503 585
R564 B.n505 B.n504 585
R565 B.n186 B.n185 585
R566 B.n187 B.n186 585
R567 B.n513 B.n512 585
R568 B.n512 B.n511 585
R569 B.n514 B.n184 585
R570 B.n184 B.n183 585
R571 B.n516 B.n515 585
R572 B.n517 B.n516 585
R573 B.n178 B.n177 585
R574 B.n179 B.n178 585
R575 B.n525 B.n524 585
R576 B.n524 B.n523 585
R577 B.n526 B.n176 585
R578 B.n176 B.n174 585
R579 B.n528 B.n527 585
R580 B.n529 B.n528 585
R581 B.n170 B.n169 585
R582 B.n175 B.n170 585
R583 B.n537 B.n536 585
R584 B.n536 B.n535 585
R585 B.n538 B.n168 585
R586 B.n168 B.n167 585
R587 B.n540 B.n539 585
R588 B.n541 B.n540 585
R589 B.n162 B.n161 585
R590 B.n163 B.n162 585
R591 B.n549 B.n548 585
R592 B.n548 B.n547 585
R593 B.n550 B.n160 585
R594 B.n160 B.n159 585
R595 B.n552 B.n551 585
R596 B.n553 B.n552 585
R597 B.n154 B.n153 585
R598 B.n155 B.n154 585
R599 B.n562 B.n561 585
R600 B.n561 B.n560 585
R601 B.n563 B.n152 585
R602 B.n559 B.n152 585
R603 B.n565 B.n564 585
R604 B.n566 B.n565 585
R605 B.n147 B.n146 585
R606 B.n148 B.n147 585
R607 B.n575 B.n574 585
R608 B.n574 B.n573 585
R609 B.n576 B.n145 585
R610 B.n145 B.n144 585
R611 B.n578 B.n577 585
R612 B.n579 B.n578 585
R613 B.n2 B.n0 585
R614 B.n4 B.n2 585
R615 B.n3 B.n1 585
R616 B.n889 B.n3 585
R617 B.n887 B.n886 585
R618 B.n888 B.n887 585
R619 B.n885 B.n9 585
R620 B.n9 B.n8 585
R621 B.n884 B.n883 585
R622 B.n883 B.n882 585
R623 B.n11 B.n10 585
R624 B.n881 B.n11 585
R625 B.n879 B.n878 585
R626 B.n880 B.n879 585
R627 B.n877 B.n15 585
R628 B.n18 B.n15 585
R629 B.n876 B.n875 585
R630 B.n875 B.n874 585
R631 B.n17 B.n16 585
R632 B.n873 B.n17 585
R633 B.n871 B.n870 585
R634 B.n872 B.n871 585
R635 B.n869 B.n23 585
R636 B.n23 B.n22 585
R637 B.n868 B.n867 585
R638 B.n867 B.n866 585
R639 B.n25 B.n24 585
R640 B.n865 B.n25 585
R641 B.n863 B.n862 585
R642 B.n864 B.n863 585
R643 B.n861 B.n30 585
R644 B.n30 B.n29 585
R645 B.n860 B.n859 585
R646 B.n859 B.n858 585
R647 B.n32 B.n31 585
R648 B.n857 B.n32 585
R649 B.n855 B.n854 585
R650 B.n856 B.n855 585
R651 B.n853 B.n37 585
R652 B.n37 B.n36 585
R653 B.n852 B.n851 585
R654 B.n851 B.n850 585
R655 B.n39 B.n38 585
R656 B.n849 B.n39 585
R657 B.n847 B.n846 585
R658 B.n848 B.n847 585
R659 B.n845 B.n44 585
R660 B.n44 B.n43 585
R661 B.n844 B.n843 585
R662 B.n843 B.n842 585
R663 B.n46 B.n45 585
R664 B.n841 B.n46 585
R665 B.n839 B.n838 585
R666 B.n840 B.n839 585
R667 B.n837 B.n50 585
R668 B.n53 B.n50 585
R669 B.n836 B.n835 585
R670 B.n835 B.n834 585
R671 B.n52 B.n51 585
R672 B.n833 B.n52 585
R673 B.n831 B.n830 585
R674 B.n832 B.n831 585
R675 B.n829 B.n58 585
R676 B.n58 B.n57 585
R677 B.n828 B.n827 585
R678 B.n827 B.n826 585
R679 B.n60 B.n59 585
R680 B.n825 B.n60 585
R681 B.n823 B.n822 585
R682 B.n824 B.n823 585
R683 B.n821 B.n65 585
R684 B.n65 B.n64 585
R685 B.n820 B.n819 585
R686 B.n819 B.n818 585
R687 B.n67 B.n66 585
R688 B.n817 B.n67 585
R689 B.n815 B.n814 585
R690 B.n816 B.n815 585
R691 B.n813 B.n72 585
R692 B.n72 B.n71 585
R693 B.n812 B.n811 585
R694 B.n811 B.n810 585
R695 B.n74 B.n73 585
R696 B.n809 B.n74 585
R697 B.n807 B.n806 585
R698 B.n808 B.n807 585
R699 B.n805 B.n79 585
R700 B.n79 B.n78 585
R701 B.n804 B.n803 585
R702 B.n803 B.n802 585
R703 B.n81 B.n80 585
R704 B.n801 B.n81 585
R705 B.n799 B.n798 585
R706 B.n800 B.n799 585
R707 B.n797 B.n86 585
R708 B.n86 B.n85 585
R709 B.n796 B.n795 585
R710 B.n795 B.n794 585
R711 B.n88 B.n87 585
R712 B.n793 B.n88 585
R713 B.n791 B.n790 585
R714 B.n792 B.n791 585
R715 B.n789 B.n93 585
R716 B.n93 B.n92 585
R717 B.n788 B.n787 585
R718 B.n787 B.n786 585
R719 B.n95 B.n94 585
R720 B.n785 B.n95 585
R721 B.n783 B.n782 585
R722 B.n784 B.n783 585
R723 B.n781 B.n100 585
R724 B.n100 B.n99 585
R725 B.n780 B.n779 585
R726 B.n779 B.n778 585
R727 B.n102 B.n101 585
R728 B.n777 B.n102 585
R729 B.n775 B.n774 585
R730 B.n776 B.n775 585
R731 B.n892 B.n891 585
R732 B.n891 B.n890 585
R733 B.n407 B.n255 492.5
R734 B.n775 B.n107 492.5
R735 B.n409 B.n253 492.5
R736 B.n141 B.n105 492.5
R737 B.n276 B.t8 257.332
R738 B.n268 B.t16 257.332
R739 B.n120 B.t12 257.332
R740 B.n126 B.t19 257.332
R741 B.n659 B.n106 256.663
R742 B.n661 B.n106 256.663
R743 B.n667 B.n106 256.663
R744 B.n669 B.n106 256.663
R745 B.n675 B.n106 256.663
R746 B.n677 B.n106 256.663
R747 B.n683 B.n106 256.663
R748 B.n685 B.n106 256.663
R749 B.n691 B.n106 256.663
R750 B.n693 B.n106 256.663
R751 B.n699 B.n106 256.663
R752 B.n129 B.n106 256.663
R753 B.n705 B.n106 256.663
R754 B.n711 B.n106 256.663
R755 B.n713 B.n106 256.663
R756 B.n719 B.n106 256.663
R757 B.n721 B.n106 256.663
R758 B.n728 B.n106 256.663
R759 B.n730 B.n106 256.663
R760 B.n736 B.n106 256.663
R761 B.n738 B.n106 256.663
R762 B.n744 B.n106 256.663
R763 B.n746 B.n106 256.663
R764 B.n752 B.n106 256.663
R765 B.n754 B.n106 256.663
R766 B.n760 B.n106 256.663
R767 B.n762 B.n106 256.663
R768 B.n768 B.n106 256.663
R769 B.n770 B.n106 256.663
R770 B.n402 B.n254 256.663
R771 B.n257 B.n254 256.663
R772 B.n395 B.n254 256.663
R773 B.n389 B.n254 256.663
R774 B.n387 B.n254 256.663
R775 B.n381 B.n254 256.663
R776 B.n379 B.n254 256.663
R777 B.n373 B.n254 256.663
R778 B.n371 B.n254 256.663
R779 B.n365 B.n254 256.663
R780 B.n363 B.n254 256.663
R781 B.n357 B.n254 256.663
R782 B.n271 B.n254 256.663
R783 B.n351 B.n254 256.663
R784 B.n345 B.n254 256.663
R785 B.n343 B.n254 256.663
R786 B.n336 B.n254 256.663
R787 B.n334 B.n254 256.663
R788 B.n328 B.n254 256.663
R789 B.n326 B.n254 256.663
R790 B.n320 B.n254 256.663
R791 B.n318 B.n254 256.663
R792 B.n312 B.n254 256.663
R793 B.n310 B.n254 256.663
R794 B.n304 B.n254 256.663
R795 B.n302 B.n254 256.663
R796 B.n296 B.n254 256.663
R797 B.n294 B.n254 256.663
R798 B.n289 B.n254 256.663
R799 B.n407 B.n249 163.367
R800 B.n415 B.n249 163.367
R801 B.n415 B.n247 163.367
R802 B.n419 B.n247 163.367
R803 B.n419 B.n241 163.367
R804 B.n427 B.n241 163.367
R805 B.n427 B.n239 163.367
R806 B.n431 B.n239 163.367
R807 B.n431 B.n233 163.367
R808 B.n439 B.n233 163.367
R809 B.n439 B.n231 163.367
R810 B.n443 B.n231 163.367
R811 B.n443 B.n225 163.367
R812 B.n451 B.n225 163.367
R813 B.n451 B.n223 163.367
R814 B.n455 B.n223 163.367
R815 B.n455 B.n217 163.367
R816 B.n463 B.n217 163.367
R817 B.n463 B.n215 163.367
R818 B.n467 B.n215 163.367
R819 B.n467 B.n209 163.367
R820 B.n475 B.n209 163.367
R821 B.n475 B.n207 163.367
R822 B.n479 B.n207 163.367
R823 B.n479 B.n201 163.367
R824 B.n487 B.n201 163.367
R825 B.n487 B.n199 163.367
R826 B.n491 B.n199 163.367
R827 B.n491 B.n193 163.367
R828 B.n500 B.n193 163.367
R829 B.n500 B.n191 163.367
R830 B.n504 B.n191 163.367
R831 B.n504 B.n186 163.367
R832 B.n512 B.n186 163.367
R833 B.n512 B.n184 163.367
R834 B.n516 B.n184 163.367
R835 B.n516 B.n178 163.367
R836 B.n524 B.n178 163.367
R837 B.n524 B.n176 163.367
R838 B.n528 B.n176 163.367
R839 B.n528 B.n170 163.367
R840 B.n536 B.n170 163.367
R841 B.n536 B.n168 163.367
R842 B.n540 B.n168 163.367
R843 B.n540 B.n162 163.367
R844 B.n548 B.n162 163.367
R845 B.n548 B.n160 163.367
R846 B.n552 B.n160 163.367
R847 B.n552 B.n154 163.367
R848 B.n561 B.n154 163.367
R849 B.n561 B.n152 163.367
R850 B.n565 B.n152 163.367
R851 B.n565 B.n147 163.367
R852 B.n574 B.n147 163.367
R853 B.n574 B.n145 163.367
R854 B.n578 B.n145 163.367
R855 B.n578 B.n2 163.367
R856 B.n891 B.n2 163.367
R857 B.n891 B.n3 163.367
R858 B.n887 B.n3 163.367
R859 B.n887 B.n9 163.367
R860 B.n883 B.n9 163.367
R861 B.n883 B.n11 163.367
R862 B.n879 B.n11 163.367
R863 B.n879 B.n15 163.367
R864 B.n875 B.n15 163.367
R865 B.n875 B.n17 163.367
R866 B.n871 B.n17 163.367
R867 B.n871 B.n23 163.367
R868 B.n867 B.n23 163.367
R869 B.n867 B.n25 163.367
R870 B.n863 B.n25 163.367
R871 B.n863 B.n30 163.367
R872 B.n859 B.n30 163.367
R873 B.n859 B.n32 163.367
R874 B.n855 B.n32 163.367
R875 B.n855 B.n37 163.367
R876 B.n851 B.n37 163.367
R877 B.n851 B.n39 163.367
R878 B.n847 B.n39 163.367
R879 B.n847 B.n44 163.367
R880 B.n843 B.n44 163.367
R881 B.n843 B.n46 163.367
R882 B.n839 B.n46 163.367
R883 B.n839 B.n50 163.367
R884 B.n835 B.n50 163.367
R885 B.n835 B.n52 163.367
R886 B.n831 B.n52 163.367
R887 B.n831 B.n58 163.367
R888 B.n827 B.n58 163.367
R889 B.n827 B.n60 163.367
R890 B.n823 B.n60 163.367
R891 B.n823 B.n65 163.367
R892 B.n819 B.n65 163.367
R893 B.n819 B.n67 163.367
R894 B.n815 B.n67 163.367
R895 B.n815 B.n72 163.367
R896 B.n811 B.n72 163.367
R897 B.n811 B.n74 163.367
R898 B.n807 B.n74 163.367
R899 B.n807 B.n79 163.367
R900 B.n803 B.n79 163.367
R901 B.n803 B.n81 163.367
R902 B.n799 B.n81 163.367
R903 B.n799 B.n86 163.367
R904 B.n795 B.n86 163.367
R905 B.n795 B.n88 163.367
R906 B.n791 B.n88 163.367
R907 B.n791 B.n93 163.367
R908 B.n787 B.n93 163.367
R909 B.n787 B.n95 163.367
R910 B.n783 B.n95 163.367
R911 B.n783 B.n100 163.367
R912 B.n779 B.n100 163.367
R913 B.n779 B.n102 163.367
R914 B.n775 B.n102 163.367
R915 B.n403 B.n401 163.367
R916 B.n401 B.n400 163.367
R917 B.n397 B.n396 163.367
R918 B.n394 B.n259 163.367
R919 B.n390 B.n388 163.367
R920 B.n386 B.n261 163.367
R921 B.n382 B.n380 163.367
R922 B.n378 B.n263 163.367
R923 B.n374 B.n372 163.367
R924 B.n370 B.n265 163.367
R925 B.n366 B.n364 163.367
R926 B.n362 B.n267 163.367
R927 B.n358 B.n356 163.367
R928 B.n353 B.n352 163.367
R929 B.n350 B.n273 163.367
R930 B.n346 B.n344 163.367
R931 B.n342 B.n275 163.367
R932 B.n337 B.n335 163.367
R933 B.n333 B.n279 163.367
R934 B.n329 B.n327 163.367
R935 B.n325 B.n281 163.367
R936 B.n321 B.n319 163.367
R937 B.n317 B.n283 163.367
R938 B.n313 B.n311 163.367
R939 B.n309 B.n285 163.367
R940 B.n305 B.n303 163.367
R941 B.n301 B.n287 163.367
R942 B.n297 B.n295 163.367
R943 B.n293 B.n290 163.367
R944 B.n409 B.n251 163.367
R945 B.n413 B.n251 163.367
R946 B.n413 B.n245 163.367
R947 B.n421 B.n245 163.367
R948 B.n421 B.n243 163.367
R949 B.n425 B.n243 163.367
R950 B.n425 B.n237 163.367
R951 B.n433 B.n237 163.367
R952 B.n433 B.n235 163.367
R953 B.n437 B.n235 163.367
R954 B.n437 B.n229 163.367
R955 B.n445 B.n229 163.367
R956 B.n445 B.n227 163.367
R957 B.n449 B.n227 163.367
R958 B.n449 B.n221 163.367
R959 B.n457 B.n221 163.367
R960 B.n457 B.n219 163.367
R961 B.n461 B.n219 163.367
R962 B.n461 B.n212 163.367
R963 B.n469 B.n212 163.367
R964 B.n469 B.n210 163.367
R965 B.n473 B.n210 163.367
R966 B.n473 B.n205 163.367
R967 B.n481 B.n205 163.367
R968 B.n481 B.n203 163.367
R969 B.n485 B.n203 163.367
R970 B.n485 B.n197 163.367
R971 B.n493 B.n197 163.367
R972 B.n493 B.n195 163.367
R973 B.n497 B.n195 163.367
R974 B.n497 B.n190 163.367
R975 B.n506 B.n190 163.367
R976 B.n506 B.n188 163.367
R977 B.n510 B.n188 163.367
R978 B.n510 B.n182 163.367
R979 B.n518 B.n182 163.367
R980 B.n518 B.n180 163.367
R981 B.n522 B.n180 163.367
R982 B.n522 B.n173 163.367
R983 B.n530 B.n173 163.367
R984 B.n530 B.n171 163.367
R985 B.n534 B.n171 163.367
R986 B.n534 B.n166 163.367
R987 B.n542 B.n166 163.367
R988 B.n542 B.n164 163.367
R989 B.n546 B.n164 163.367
R990 B.n546 B.n158 163.367
R991 B.n554 B.n158 163.367
R992 B.n554 B.n156 163.367
R993 B.n558 B.n156 163.367
R994 B.n558 B.n151 163.367
R995 B.n567 B.n151 163.367
R996 B.n567 B.n149 163.367
R997 B.n572 B.n149 163.367
R998 B.n572 B.n143 163.367
R999 B.n580 B.n143 163.367
R1000 B.n581 B.n580 163.367
R1001 B.n581 B.n5 163.367
R1002 B.n6 B.n5 163.367
R1003 B.n7 B.n6 163.367
R1004 B.n586 B.n7 163.367
R1005 B.n586 B.n12 163.367
R1006 B.n13 B.n12 163.367
R1007 B.n14 B.n13 163.367
R1008 B.n591 B.n14 163.367
R1009 B.n591 B.n19 163.367
R1010 B.n20 B.n19 163.367
R1011 B.n21 B.n20 163.367
R1012 B.n596 B.n21 163.367
R1013 B.n596 B.n26 163.367
R1014 B.n27 B.n26 163.367
R1015 B.n28 B.n27 163.367
R1016 B.n601 B.n28 163.367
R1017 B.n601 B.n33 163.367
R1018 B.n34 B.n33 163.367
R1019 B.n35 B.n34 163.367
R1020 B.n606 B.n35 163.367
R1021 B.n606 B.n40 163.367
R1022 B.n41 B.n40 163.367
R1023 B.n42 B.n41 163.367
R1024 B.n611 B.n42 163.367
R1025 B.n611 B.n47 163.367
R1026 B.n48 B.n47 163.367
R1027 B.n49 B.n48 163.367
R1028 B.n616 B.n49 163.367
R1029 B.n616 B.n54 163.367
R1030 B.n55 B.n54 163.367
R1031 B.n56 B.n55 163.367
R1032 B.n621 B.n56 163.367
R1033 B.n621 B.n61 163.367
R1034 B.n62 B.n61 163.367
R1035 B.n63 B.n62 163.367
R1036 B.n626 B.n63 163.367
R1037 B.n626 B.n68 163.367
R1038 B.n69 B.n68 163.367
R1039 B.n70 B.n69 163.367
R1040 B.n631 B.n70 163.367
R1041 B.n631 B.n75 163.367
R1042 B.n76 B.n75 163.367
R1043 B.n77 B.n76 163.367
R1044 B.n636 B.n77 163.367
R1045 B.n636 B.n82 163.367
R1046 B.n83 B.n82 163.367
R1047 B.n84 B.n83 163.367
R1048 B.n641 B.n84 163.367
R1049 B.n641 B.n89 163.367
R1050 B.n90 B.n89 163.367
R1051 B.n91 B.n90 163.367
R1052 B.n646 B.n91 163.367
R1053 B.n646 B.n96 163.367
R1054 B.n97 B.n96 163.367
R1055 B.n98 B.n97 163.367
R1056 B.n651 B.n98 163.367
R1057 B.n651 B.n103 163.367
R1058 B.n104 B.n103 163.367
R1059 B.n105 B.n104 163.367
R1060 B.n771 B.n769 163.367
R1061 B.n767 B.n109 163.367
R1062 B.n763 B.n761 163.367
R1063 B.n759 B.n111 163.367
R1064 B.n755 B.n753 163.367
R1065 B.n751 B.n113 163.367
R1066 B.n747 B.n745 163.367
R1067 B.n743 B.n115 163.367
R1068 B.n739 B.n737 163.367
R1069 B.n735 B.n117 163.367
R1070 B.n731 B.n729 163.367
R1071 B.n727 B.n119 163.367
R1072 B.n722 B.n720 163.367
R1073 B.n718 B.n123 163.367
R1074 B.n714 B.n712 163.367
R1075 B.n710 B.n125 163.367
R1076 B.n706 B.n704 163.367
R1077 B.n701 B.n700 163.367
R1078 B.n698 B.n131 163.367
R1079 B.n694 B.n692 163.367
R1080 B.n690 B.n133 163.367
R1081 B.n686 B.n684 163.367
R1082 B.n682 B.n135 163.367
R1083 B.n678 B.n676 163.367
R1084 B.n674 B.n137 163.367
R1085 B.n670 B.n668 163.367
R1086 B.n666 B.n139 163.367
R1087 B.n662 B.n660 163.367
R1088 B.n658 B.n141 163.367
R1089 B.n276 B.t11 136.827
R1090 B.n126 B.t20 136.827
R1091 B.n268 B.t18 136.821
R1092 B.n120 B.t14 136.821
R1093 B.n408 B.n254 125.578
R1094 B.n776 B.n106 125.578
R1095 B.n402 B.n255 71.676
R1096 B.n400 B.n257 71.676
R1097 B.n396 B.n395 71.676
R1098 B.n389 B.n259 71.676
R1099 B.n388 B.n387 71.676
R1100 B.n381 B.n261 71.676
R1101 B.n380 B.n379 71.676
R1102 B.n373 B.n263 71.676
R1103 B.n372 B.n371 71.676
R1104 B.n365 B.n265 71.676
R1105 B.n364 B.n363 71.676
R1106 B.n357 B.n267 71.676
R1107 B.n356 B.n271 71.676
R1108 B.n352 B.n351 71.676
R1109 B.n345 B.n273 71.676
R1110 B.n344 B.n343 71.676
R1111 B.n336 B.n275 71.676
R1112 B.n335 B.n334 71.676
R1113 B.n328 B.n279 71.676
R1114 B.n327 B.n326 71.676
R1115 B.n320 B.n281 71.676
R1116 B.n319 B.n318 71.676
R1117 B.n312 B.n283 71.676
R1118 B.n311 B.n310 71.676
R1119 B.n304 B.n285 71.676
R1120 B.n303 B.n302 71.676
R1121 B.n296 B.n287 71.676
R1122 B.n295 B.n294 71.676
R1123 B.n290 B.n289 71.676
R1124 B.n770 B.n107 71.676
R1125 B.n769 B.n768 71.676
R1126 B.n762 B.n109 71.676
R1127 B.n761 B.n760 71.676
R1128 B.n754 B.n111 71.676
R1129 B.n753 B.n752 71.676
R1130 B.n746 B.n113 71.676
R1131 B.n745 B.n744 71.676
R1132 B.n738 B.n115 71.676
R1133 B.n737 B.n736 71.676
R1134 B.n730 B.n117 71.676
R1135 B.n729 B.n728 71.676
R1136 B.n721 B.n119 71.676
R1137 B.n720 B.n719 71.676
R1138 B.n713 B.n123 71.676
R1139 B.n712 B.n711 71.676
R1140 B.n705 B.n125 71.676
R1141 B.n704 B.n129 71.676
R1142 B.n700 B.n699 71.676
R1143 B.n693 B.n131 71.676
R1144 B.n692 B.n691 71.676
R1145 B.n685 B.n133 71.676
R1146 B.n684 B.n683 71.676
R1147 B.n677 B.n135 71.676
R1148 B.n676 B.n675 71.676
R1149 B.n669 B.n137 71.676
R1150 B.n668 B.n667 71.676
R1151 B.n661 B.n139 71.676
R1152 B.n660 B.n659 71.676
R1153 B.n659 B.n658 71.676
R1154 B.n662 B.n661 71.676
R1155 B.n667 B.n666 71.676
R1156 B.n670 B.n669 71.676
R1157 B.n675 B.n674 71.676
R1158 B.n678 B.n677 71.676
R1159 B.n683 B.n682 71.676
R1160 B.n686 B.n685 71.676
R1161 B.n691 B.n690 71.676
R1162 B.n694 B.n693 71.676
R1163 B.n699 B.n698 71.676
R1164 B.n701 B.n129 71.676
R1165 B.n706 B.n705 71.676
R1166 B.n711 B.n710 71.676
R1167 B.n714 B.n713 71.676
R1168 B.n719 B.n718 71.676
R1169 B.n722 B.n721 71.676
R1170 B.n728 B.n727 71.676
R1171 B.n731 B.n730 71.676
R1172 B.n736 B.n735 71.676
R1173 B.n739 B.n738 71.676
R1174 B.n744 B.n743 71.676
R1175 B.n747 B.n746 71.676
R1176 B.n752 B.n751 71.676
R1177 B.n755 B.n754 71.676
R1178 B.n760 B.n759 71.676
R1179 B.n763 B.n762 71.676
R1180 B.n768 B.n767 71.676
R1181 B.n771 B.n770 71.676
R1182 B.n403 B.n402 71.676
R1183 B.n397 B.n257 71.676
R1184 B.n395 B.n394 71.676
R1185 B.n390 B.n389 71.676
R1186 B.n387 B.n386 71.676
R1187 B.n382 B.n381 71.676
R1188 B.n379 B.n378 71.676
R1189 B.n374 B.n373 71.676
R1190 B.n371 B.n370 71.676
R1191 B.n366 B.n365 71.676
R1192 B.n363 B.n362 71.676
R1193 B.n358 B.n357 71.676
R1194 B.n353 B.n271 71.676
R1195 B.n351 B.n350 71.676
R1196 B.n346 B.n345 71.676
R1197 B.n343 B.n342 71.676
R1198 B.n337 B.n336 71.676
R1199 B.n334 B.n333 71.676
R1200 B.n329 B.n328 71.676
R1201 B.n326 B.n325 71.676
R1202 B.n321 B.n320 71.676
R1203 B.n318 B.n317 71.676
R1204 B.n313 B.n312 71.676
R1205 B.n310 B.n309 71.676
R1206 B.n305 B.n304 71.676
R1207 B.n302 B.n301 71.676
R1208 B.n297 B.n296 71.676
R1209 B.n294 B.n293 71.676
R1210 B.n289 B.n253 71.676
R1211 B.n277 B.t10 70.8882
R1212 B.n127 B.t21 70.8882
R1213 B.n269 B.t17 70.8814
R1214 B.n121 B.t15 70.8814
R1215 B.n277 B.n276 65.9399
R1216 B.n269 B.n268 65.9399
R1217 B.n121 B.n120 65.9399
R1218 B.n127 B.n126 65.9399
R1219 B.n408 B.n250 65.1857
R1220 B.n414 B.n250 65.1857
R1221 B.n414 B.n246 65.1857
R1222 B.n420 B.n246 65.1857
R1223 B.n420 B.n242 65.1857
R1224 B.n426 B.n242 65.1857
R1225 B.n426 B.n238 65.1857
R1226 B.n432 B.n238 65.1857
R1227 B.n438 B.n234 65.1857
R1228 B.n438 B.n230 65.1857
R1229 B.n444 B.n230 65.1857
R1230 B.n444 B.n226 65.1857
R1231 B.n450 B.n226 65.1857
R1232 B.n450 B.n222 65.1857
R1233 B.n456 B.n222 65.1857
R1234 B.n456 B.n218 65.1857
R1235 B.n462 B.n218 65.1857
R1236 B.n462 B.n213 65.1857
R1237 B.n468 B.n213 65.1857
R1238 B.n468 B.n214 65.1857
R1239 B.n474 B.n206 65.1857
R1240 B.n480 B.n206 65.1857
R1241 B.n480 B.n202 65.1857
R1242 B.n486 B.n202 65.1857
R1243 B.n486 B.n198 65.1857
R1244 B.n492 B.n198 65.1857
R1245 B.n492 B.n194 65.1857
R1246 B.n499 B.n194 65.1857
R1247 B.n499 B.n498 65.1857
R1248 B.n505 B.n187 65.1857
R1249 B.n511 B.n187 65.1857
R1250 B.n511 B.n183 65.1857
R1251 B.n517 B.n183 65.1857
R1252 B.n517 B.n179 65.1857
R1253 B.n523 B.n179 65.1857
R1254 B.n523 B.n174 65.1857
R1255 B.n529 B.n174 65.1857
R1256 B.n529 B.n175 65.1857
R1257 B.n535 B.n167 65.1857
R1258 B.n541 B.n167 65.1857
R1259 B.n541 B.n163 65.1857
R1260 B.n547 B.n163 65.1857
R1261 B.n547 B.n159 65.1857
R1262 B.n553 B.n159 65.1857
R1263 B.n553 B.n155 65.1857
R1264 B.n560 B.n155 65.1857
R1265 B.n560 B.n559 65.1857
R1266 B.n566 B.n148 65.1857
R1267 B.n573 B.n148 65.1857
R1268 B.n573 B.n144 65.1857
R1269 B.n579 B.n144 65.1857
R1270 B.n579 B.n4 65.1857
R1271 B.n890 B.n4 65.1857
R1272 B.n890 B.n889 65.1857
R1273 B.n889 B.n888 65.1857
R1274 B.n888 B.n8 65.1857
R1275 B.n882 B.n8 65.1857
R1276 B.n882 B.n881 65.1857
R1277 B.n881 B.n880 65.1857
R1278 B.n874 B.n18 65.1857
R1279 B.n874 B.n873 65.1857
R1280 B.n873 B.n872 65.1857
R1281 B.n872 B.n22 65.1857
R1282 B.n866 B.n22 65.1857
R1283 B.n866 B.n865 65.1857
R1284 B.n865 B.n864 65.1857
R1285 B.n864 B.n29 65.1857
R1286 B.n858 B.n29 65.1857
R1287 B.n857 B.n856 65.1857
R1288 B.n856 B.n36 65.1857
R1289 B.n850 B.n36 65.1857
R1290 B.n850 B.n849 65.1857
R1291 B.n849 B.n848 65.1857
R1292 B.n848 B.n43 65.1857
R1293 B.n842 B.n43 65.1857
R1294 B.n842 B.n841 65.1857
R1295 B.n841 B.n840 65.1857
R1296 B.n834 B.n53 65.1857
R1297 B.n834 B.n833 65.1857
R1298 B.n833 B.n832 65.1857
R1299 B.n832 B.n57 65.1857
R1300 B.n826 B.n57 65.1857
R1301 B.n826 B.n825 65.1857
R1302 B.n825 B.n824 65.1857
R1303 B.n824 B.n64 65.1857
R1304 B.n818 B.n64 65.1857
R1305 B.n817 B.n816 65.1857
R1306 B.n816 B.n71 65.1857
R1307 B.n810 B.n71 65.1857
R1308 B.n810 B.n809 65.1857
R1309 B.n809 B.n808 65.1857
R1310 B.n808 B.n78 65.1857
R1311 B.n802 B.n78 65.1857
R1312 B.n802 B.n801 65.1857
R1313 B.n801 B.n800 65.1857
R1314 B.n800 B.n85 65.1857
R1315 B.n794 B.n85 65.1857
R1316 B.n794 B.n793 65.1857
R1317 B.n792 B.n92 65.1857
R1318 B.n786 B.n92 65.1857
R1319 B.n786 B.n785 65.1857
R1320 B.n785 B.n784 65.1857
R1321 B.n784 B.n99 65.1857
R1322 B.n778 B.n99 65.1857
R1323 B.n778 B.n777 65.1857
R1324 B.n777 B.n776 65.1857
R1325 B.n339 B.n277 59.5399
R1326 B.n270 B.n269 59.5399
R1327 B.n724 B.n121 59.5399
R1328 B.n128 B.n127 59.5399
R1329 B.t9 B.n234 52.7238
R1330 B.n793 B.t13 52.7238
R1331 B.n474 B.t6 39.3033
R1332 B.n505 B.t2 39.3033
R1333 B.n535 B.t7 39.3033
R1334 B.n566 B.t3 39.3033
R1335 B.n880 B.t5 39.3033
R1336 B.n858 B.t1 39.3033
R1337 B.n840 B.t4 39.3033
R1338 B.n818 B.t0 39.3033
R1339 B.n774 B.n773 32.0005
R1340 B.n656 B.n655 32.0005
R1341 B.n410 B.n252 32.0005
R1342 B.n406 B.n405 32.0005
R1343 B.n214 B.t6 25.8829
R1344 B.n498 B.t2 25.8829
R1345 B.n175 B.t7 25.8829
R1346 B.n559 B.t3 25.8829
R1347 B.n18 B.t5 25.8829
R1348 B.t1 B.n857 25.8829
R1349 B.n53 B.t4 25.8829
R1350 B.t0 B.n817 25.8829
R1351 B B.n892 18.0485
R1352 B.n432 B.t9 12.4624
R1353 B.t13 B.n792 12.4624
R1354 B.n773 B.n772 10.6151
R1355 B.n772 B.n108 10.6151
R1356 B.n766 B.n108 10.6151
R1357 B.n766 B.n765 10.6151
R1358 B.n765 B.n764 10.6151
R1359 B.n764 B.n110 10.6151
R1360 B.n758 B.n110 10.6151
R1361 B.n758 B.n757 10.6151
R1362 B.n757 B.n756 10.6151
R1363 B.n756 B.n112 10.6151
R1364 B.n750 B.n112 10.6151
R1365 B.n750 B.n749 10.6151
R1366 B.n749 B.n748 10.6151
R1367 B.n748 B.n114 10.6151
R1368 B.n742 B.n114 10.6151
R1369 B.n742 B.n741 10.6151
R1370 B.n741 B.n740 10.6151
R1371 B.n740 B.n116 10.6151
R1372 B.n734 B.n116 10.6151
R1373 B.n734 B.n733 10.6151
R1374 B.n733 B.n732 10.6151
R1375 B.n732 B.n118 10.6151
R1376 B.n726 B.n118 10.6151
R1377 B.n726 B.n725 10.6151
R1378 B.n723 B.n122 10.6151
R1379 B.n717 B.n122 10.6151
R1380 B.n717 B.n716 10.6151
R1381 B.n716 B.n715 10.6151
R1382 B.n715 B.n124 10.6151
R1383 B.n709 B.n124 10.6151
R1384 B.n709 B.n708 10.6151
R1385 B.n708 B.n707 10.6151
R1386 B.n703 B.n702 10.6151
R1387 B.n702 B.n130 10.6151
R1388 B.n697 B.n130 10.6151
R1389 B.n697 B.n696 10.6151
R1390 B.n696 B.n695 10.6151
R1391 B.n695 B.n132 10.6151
R1392 B.n689 B.n132 10.6151
R1393 B.n689 B.n688 10.6151
R1394 B.n688 B.n687 10.6151
R1395 B.n687 B.n134 10.6151
R1396 B.n681 B.n134 10.6151
R1397 B.n681 B.n680 10.6151
R1398 B.n680 B.n679 10.6151
R1399 B.n679 B.n136 10.6151
R1400 B.n673 B.n136 10.6151
R1401 B.n673 B.n672 10.6151
R1402 B.n672 B.n671 10.6151
R1403 B.n671 B.n138 10.6151
R1404 B.n665 B.n138 10.6151
R1405 B.n665 B.n664 10.6151
R1406 B.n664 B.n663 10.6151
R1407 B.n663 B.n140 10.6151
R1408 B.n657 B.n140 10.6151
R1409 B.n657 B.n656 10.6151
R1410 B.n411 B.n410 10.6151
R1411 B.n412 B.n411 10.6151
R1412 B.n412 B.n244 10.6151
R1413 B.n422 B.n244 10.6151
R1414 B.n423 B.n422 10.6151
R1415 B.n424 B.n423 10.6151
R1416 B.n424 B.n236 10.6151
R1417 B.n434 B.n236 10.6151
R1418 B.n435 B.n434 10.6151
R1419 B.n436 B.n435 10.6151
R1420 B.n436 B.n228 10.6151
R1421 B.n446 B.n228 10.6151
R1422 B.n447 B.n446 10.6151
R1423 B.n448 B.n447 10.6151
R1424 B.n448 B.n220 10.6151
R1425 B.n458 B.n220 10.6151
R1426 B.n459 B.n458 10.6151
R1427 B.n460 B.n459 10.6151
R1428 B.n460 B.n211 10.6151
R1429 B.n470 B.n211 10.6151
R1430 B.n471 B.n470 10.6151
R1431 B.n472 B.n471 10.6151
R1432 B.n472 B.n204 10.6151
R1433 B.n482 B.n204 10.6151
R1434 B.n483 B.n482 10.6151
R1435 B.n484 B.n483 10.6151
R1436 B.n484 B.n196 10.6151
R1437 B.n494 B.n196 10.6151
R1438 B.n495 B.n494 10.6151
R1439 B.n496 B.n495 10.6151
R1440 B.n496 B.n189 10.6151
R1441 B.n507 B.n189 10.6151
R1442 B.n508 B.n507 10.6151
R1443 B.n509 B.n508 10.6151
R1444 B.n509 B.n181 10.6151
R1445 B.n519 B.n181 10.6151
R1446 B.n520 B.n519 10.6151
R1447 B.n521 B.n520 10.6151
R1448 B.n521 B.n172 10.6151
R1449 B.n531 B.n172 10.6151
R1450 B.n532 B.n531 10.6151
R1451 B.n533 B.n532 10.6151
R1452 B.n533 B.n165 10.6151
R1453 B.n543 B.n165 10.6151
R1454 B.n544 B.n543 10.6151
R1455 B.n545 B.n544 10.6151
R1456 B.n545 B.n157 10.6151
R1457 B.n555 B.n157 10.6151
R1458 B.n556 B.n555 10.6151
R1459 B.n557 B.n556 10.6151
R1460 B.n557 B.n150 10.6151
R1461 B.n568 B.n150 10.6151
R1462 B.n569 B.n568 10.6151
R1463 B.n571 B.n569 10.6151
R1464 B.n571 B.n570 10.6151
R1465 B.n570 B.n142 10.6151
R1466 B.n582 B.n142 10.6151
R1467 B.n583 B.n582 10.6151
R1468 B.n584 B.n583 10.6151
R1469 B.n585 B.n584 10.6151
R1470 B.n587 B.n585 10.6151
R1471 B.n588 B.n587 10.6151
R1472 B.n589 B.n588 10.6151
R1473 B.n590 B.n589 10.6151
R1474 B.n592 B.n590 10.6151
R1475 B.n593 B.n592 10.6151
R1476 B.n594 B.n593 10.6151
R1477 B.n595 B.n594 10.6151
R1478 B.n597 B.n595 10.6151
R1479 B.n598 B.n597 10.6151
R1480 B.n599 B.n598 10.6151
R1481 B.n600 B.n599 10.6151
R1482 B.n602 B.n600 10.6151
R1483 B.n603 B.n602 10.6151
R1484 B.n604 B.n603 10.6151
R1485 B.n605 B.n604 10.6151
R1486 B.n607 B.n605 10.6151
R1487 B.n608 B.n607 10.6151
R1488 B.n609 B.n608 10.6151
R1489 B.n610 B.n609 10.6151
R1490 B.n612 B.n610 10.6151
R1491 B.n613 B.n612 10.6151
R1492 B.n614 B.n613 10.6151
R1493 B.n615 B.n614 10.6151
R1494 B.n617 B.n615 10.6151
R1495 B.n618 B.n617 10.6151
R1496 B.n619 B.n618 10.6151
R1497 B.n620 B.n619 10.6151
R1498 B.n622 B.n620 10.6151
R1499 B.n623 B.n622 10.6151
R1500 B.n624 B.n623 10.6151
R1501 B.n625 B.n624 10.6151
R1502 B.n627 B.n625 10.6151
R1503 B.n628 B.n627 10.6151
R1504 B.n629 B.n628 10.6151
R1505 B.n630 B.n629 10.6151
R1506 B.n632 B.n630 10.6151
R1507 B.n633 B.n632 10.6151
R1508 B.n634 B.n633 10.6151
R1509 B.n635 B.n634 10.6151
R1510 B.n637 B.n635 10.6151
R1511 B.n638 B.n637 10.6151
R1512 B.n639 B.n638 10.6151
R1513 B.n640 B.n639 10.6151
R1514 B.n642 B.n640 10.6151
R1515 B.n643 B.n642 10.6151
R1516 B.n644 B.n643 10.6151
R1517 B.n645 B.n644 10.6151
R1518 B.n647 B.n645 10.6151
R1519 B.n648 B.n647 10.6151
R1520 B.n649 B.n648 10.6151
R1521 B.n650 B.n649 10.6151
R1522 B.n652 B.n650 10.6151
R1523 B.n653 B.n652 10.6151
R1524 B.n654 B.n653 10.6151
R1525 B.n655 B.n654 10.6151
R1526 B.n405 B.n404 10.6151
R1527 B.n404 B.n256 10.6151
R1528 B.n399 B.n256 10.6151
R1529 B.n399 B.n398 10.6151
R1530 B.n398 B.n258 10.6151
R1531 B.n393 B.n258 10.6151
R1532 B.n393 B.n392 10.6151
R1533 B.n392 B.n391 10.6151
R1534 B.n391 B.n260 10.6151
R1535 B.n385 B.n260 10.6151
R1536 B.n385 B.n384 10.6151
R1537 B.n384 B.n383 10.6151
R1538 B.n383 B.n262 10.6151
R1539 B.n377 B.n262 10.6151
R1540 B.n377 B.n376 10.6151
R1541 B.n376 B.n375 10.6151
R1542 B.n375 B.n264 10.6151
R1543 B.n369 B.n264 10.6151
R1544 B.n369 B.n368 10.6151
R1545 B.n368 B.n367 10.6151
R1546 B.n367 B.n266 10.6151
R1547 B.n361 B.n266 10.6151
R1548 B.n361 B.n360 10.6151
R1549 B.n360 B.n359 10.6151
R1550 B.n355 B.n354 10.6151
R1551 B.n354 B.n272 10.6151
R1552 B.n349 B.n272 10.6151
R1553 B.n349 B.n348 10.6151
R1554 B.n348 B.n347 10.6151
R1555 B.n347 B.n274 10.6151
R1556 B.n341 B.n274 10.6151
R1557 B.n341 B.n340 10.6151
R1558 B.n338 B.n278 10.6151
R1559 B.n332 B.n278 10.6151
R1560 B.n332 B.n331 10.6151
R1561 B.n331 B.n330 10.6151
R1562 B.n330 B.n280 10.6151
R1563 B.n324 B.n280 10.6151
R1564 B.n324 B.n323 10.6151
R1565 B.n323 B.n322 10.6151
R1566 B.n322 B.n282 10.6151
R1567 B.n316 B.n282 10.6151
R1568 B.n316 B.n315 10.6151
R1569 B.n315 B.n314 10.6151
R1570 B.n314 B.n284 10.6151
R1571 B.n308 B.n284 10.6151
R1572 B.n308 B.n307 10.6151
R1573 B.n307 B.n306 10.6151
R1574 B.n306 B.n286 10.6151
R1575 B.n300 B.n286 10.6151
R1576 B.n300 B.n299 10.6151
R1577 B.n299 B.n298 10.6151
R1578 B.n298 B.n288 10.6151
R1579 B.n292 B.n288 10.6151
R1580 B.n292 B.n291 10.6151
R1581 B.n291 B.n252 10.6151
R1582 B.n406 B.n248 10.6151
R1583 B.n416 B.n248 10.6151
R1584 B.n417 B.n416 10.6151
R1585 B.n418 B.n417 10.6151
R1586 B.n418 B.n240 10.6151
R1587 B.n428 B.n240 10.6151
R1588 B.n429 B.n428 10.6151
R1589 B.n430 B.n429 10.6151
R1590 B.n430 B.n232 10.6151
R1591 B.n440 B.n232 10.6151
R1592 B.n441 B.n440 10.6151
R1593 B.n442 B.n441 10.6151
R1594 B.n442 B.n224 10.6151
R1595 B.n452 B.n224 10.6151
R1596 B.n453 B.n452 10.6151
R1597 B.n454 B.n453 10.6151
R1598 B.n454 B.n216 10.6151
R1599 B.n464 B.n216 10.6151
R1600 B.n465 B.n464 10.6151
R1601 B.n466 B.n465 10.6151
R1602 B.n466 B.n208 10.6151
R1603 B.n476 B.n208 10.6151
R1604 B.n477 B.n476 10.6151
R1605 B.n478 B.n477 10.6151
R1606 B.n478 B.n200 10.6151
R1607 B.n488 B.n200 10.6151
R1608 B.n489 B.n488 10.6151
R1609 B.n490 B.n489 10.6151
R1610 B.n490 B.n192 10.6151
R1611 B.n501 B.n192 10.6151
R1612 B.n502 B.n501 10.6151
R1613 B.n503 B.n502 10.6151
R1614 B.n503 B.n185 10.6151
R1615 B.n513 B.n185 10.6151
R1616 B.n514 B.n513 10.6151
R1617 B.n515 B.n514 10.6151
R1618 B.n515 B.n177 10.6151
R1619 B.n525 B.n177 10.6151
R1620 B.n526 B.n525 10.6151
R1621 B.n527 B.n526 10.6151
R1622 B.n527 B.n169 10.6151
R1623 B.n537 B.n169 10.6151
R1624 B.n538 B.n537 10.6151
R1625 B.n539 B.n538 10.6151
R1626 B.n539 B.n161 10.6151
R1627 B.n549 B.n161 10.6151
R1628 B.n550 B.n549 10.6151
R1629 B.n551 B.n550 10.6151
R1630 B.n551 B.n153 10.6151
R1631 B.n562 B.n153 10.6151
R1632 B.n563 B.n562 10.6151
R1633 B.n564 B.n563 10.6151
R1634 B.n564 B.n146 10.6151
R1635 B.n575 B.n146 10.6151
R1636 B.n576 B.n575 10.6151
R1637 B.n577 B.n576 10.6151
R1638 B.n577 B.n0 10.6151
R1639 B.n886 B.n1 10.6151
R1640 B.n886 B.n885 10.6151
R1641 B.n885 B.n884 10.6151
R1642 B.n884 B.n10 10.6151
R1643 B.n878 B.n10 10.6151
R1644 B.n878 B.n877 10.6151
R1645 B.n877 B.n876 10.6151
R1646 B.n876 B.n16 10.6151
R1647 B.n870 B.n16 10.6151
R1648 B.n870 B.n869 10.6151
R1649 B.n869 B.n868 10.6151
R1650 B.n868 B.n24 10.6151
R1651 B.n862 B.n24 10.6151
R1652 B.n862 B.n861 10.6151
R1653 B.n861 B.n860 10.6151
R1654 B.n860 B.n31 10.6151
R1655 B.n854 B.n31 10.6151
R1656 B.n854 B.n853 10.6151
R1657 B.n853 B.n852 10.6151
R1658 B.n852 B.n38 10.6151
R1659 B.n846 B.n38 10.6151
R1660 B.n846 B.n845 10.6151
R1661 B.n845 B.n844 10.6151
R1662 B.n844 B.n45 10.6151
R1663 B.n838 B.n45 10.6151
R1664 B.n838 B.n837 10.6151
R1665 B.n837 B.n836 10.6151
R1666 B.n836 B.n51 10.6151
R1667 B.n830 B.n51 10.6151
R1668 B.n830 B.n829 10.6151
R1669 B.n829 B.n828 10.6151
R1670 B.n828 B.n59 10.6151
R1671 B.n822 B.n59 10.6151
R1672 B.n822 B.n821 10.6151
R1673 B.n821 B.n820 10.6151
R1674 B.n820 B.n66 10.6151
R1675 B.n814 B.n66 10.6151
R1676 B.n814 B.n813 10.6151
R1677 B.n813 B.n812 10.6151
R1678 B.n812 B.n73 10.6151
R1679 B.n806 B.n73 10.6151
R1680 B.n806 B.n805 10.6151
R1681 B.n805 B.n804 10.6151
R1682 B.n804 B.n80 10.6151
R1683 B.n798 B.n80 10.6151
R1684 B.n798 B.n797 10.6151
R1685 B.n797 B.n796 10.6151
R1686 B.n796 B.n87 10.6151
R1687 B.n790 B.n87 10.6151
R1688 B.n790 B.n789 10.6151
R1689 B.n789 B.n788 10.6151
R1690 B.n788 B.n94 10.6151
R1691 B.n782 B.n94 10.6151
R1692 B.n782 B.n781 10.6151
R1693 B.n781 B.n780 10.6151
R1694 B.n780 B.n101 10.6151
R1695 B.n774 B.n101 10.6151
R1696 B.n724 B.n723 6.5566
R1697 B.n707 B.n128 6.5566
R1698 B.n355 B.n270 6.5566
R1699 B.n340 B.n339 6.5566
R1700 B.n725 B.n724 4.05904
R1701 B.n703 B.n128 4.05904
R1702 B.n359 B.n270 4.05904
R1703 B.n339 B.n338 4.05904
R1704 B.n892 B.n0 2.81026
R1705 B.n892 B.n1 2.81026
R1706 VP.n21 VP.n18 161.3
R1707 VP.n23 VP.n22 161.3
R1708 VP.n24 VP.n17 161.3
R1709 VP.n26 VP.n25 161.3
R1710 VP.n27 VP.n16 161.3
R1711 VP.n29 VP.n28 161.3
R1712 VP.n31 VP.n30 161.3
R1713 VP.n32 VP.n14 161.3
R1714 VP.n34 VP.n33 161.3
R1715 VP.n35 VP.n13 161.3
R1716 VP.n37 VP.n36 161.3
R1717 VP.n38 VP.n12 161.3
R1718 VP.n40 VP.n39 161.3
R1719 VP.n75 VP.n74 161.3
R1720 VP.n73 VP.n1 161.3
R1721 VP.n72 VP.n71 161.3
R1722 VP.n70 VP.n2 161.3
R1723 VP.n69 VP.n68 161.3
R1724 VP.n67 VP.n3 161.3
R1725 VP.n66 VP.n65 161.3
R1726 VP.n64 VP.n63 161.3
R1727 VP.n62 VP.n5 161.3
R1728 VP.n61 VP.n60 161.3
R1729 VP.n59 VP.n6 161.3
R1730 VP.n58 VP.n57 161.3
R1731 VP.n56 VP.n7 161.3
R1732 VP.n54 VP.n53 161.3
R1733 VP.n52 VP.n8 161.3
R1734 VP.n51 VP.n50 161.3
R1735 VP.n49 VP.n9 161.3
R1736 VP.n48 VP.n47 161.3
R1737 VP.n46 VP.n10 161.3
R1738 VP.n45 VP.n44 161.3
R1739 VP.n19 VP.t1 82.0219
R1740 VP.n43 VP.n42 73.0313
R1741 VP.n76 VP.n0 73.0313
R1742 VP.n41 VP.n11 73.0313
R1743 VP.n61 VP.n6 56.5617
R1744 VP.n26 VP.n17 56.5617
R1745 VP.n49 VP.n48 55.1086
R1746 VP.n72 VP.n2 55.1086
R1747 VP.n37 VP.n13 55.1086
R1748 VP.n20 VP.n19 51.9075
R1749 VP.n42 VP.n41 48.795
R1750 VP.n43 VP.t7 48.6715
R1751 VP.n55 VP.t3 48.6715
R1752 VP.n4 VP.t6 48.6715
R1753 VP.n0 VP.t0 48.6715
R1754 VP.n11 VP.t5 48.6715
R1755 VP.n15 VP.t4 48.6715
R1756 VP.n20 VP.t2 48.6715
R1757 VP.n50 VP.n49 26.0455
R1758 VP.n68 VP.n2 26.0455
R1759 VP.n33 VP.n13 26.0455
R1760 VP.n44 VP.n10 24.5923
R1761 VP.n48 VP.n10 24.5923
R1762 VP.n50 VP.n8 24.5923
R1763 VP.n54 VP.n8 24.5923
R1764 VP.n57 VP.n56 24.5923
R1765 VP.n57 VP.n6 24.5923
R1766 VP.n62 VP.n61 24.5923
R1767 VP.n63 VP.n62 24.5923
R1768 VP.n67 VP.n66 24.5923
R1769 VP.n68 VP.n67 24.5923
R1770 VP.n73 VP.n72 24.5923
R1771 VP.n74 VP.n73 24.5923
R1772 VP.n38 VP.n37 24.5923
R1773 VP.n39 VP.n38 24.5923
R1774 VP.n27 VP.n26 24.5923
R1775 VP.n28 VP.n27 24.5923
R1776 VP.n32 VP.n31 24.5923
R1777 VP.n33 VP.n32 24.5923
R1778 VP.n22 VP.n21 24.5923
R1779 VP.n22 VP.n17 24.5923
R1780 VP.n56 VP.n55 22.1332
R1781 VP.n63 VP.n4 22.1332
R1782 VP.n28 VP.n15 22.1332
R1783 VP.n21 VP.n20 22.1332
R1784 VP.n44 VP.n43 17.2148
R1785 VP.n74 VP.n0 17.2148
R1786 VP.n39 VP.n11 17.2148
R1787 VP.n19 VP.n18 4.03537
R1788 VP.n55 VP.n54 2.45968
R1789 VP.n66 VP.n4 2.45968
R1790 VP.n31 VP.n15 2.45968
R1791 VP.n41 VP.n40 0.354861
R1792 VP.n45 VP.n42 0.354861
R1793 VP.n76 VP.n75 0.354861
R1794 VP VP.n76 0.267071
R1795 VP.n23 VP.n18 0.189894
R1796 VP.n24 VP.n23 0.189894
R1797 VP.n25 VP.n24 0.189894
R1798 VP.n25 VP.n16 0.189894
R1799 VP.n29 VP.n16 0.189894
R1800 VP.n30 VP.n29 0.189894
R1801 VP.n30 VP.n14 0.189894
R1802 VP.n34 VP.n14 0.189894
R1803 VP.n35 VP.n34 0.189894
R1804 VP.n36 VP.n35 0.189894
R1805 VP.n36 VP.n12 0.189894
R1806 VP.n40 VP.n12 0.189894
R1807 VP.n46 VP.n45 0.189894
R1808 VP.n47 VP.n46 0.189894
R1809 VP.n47 VP.n9 0.189894
R1810 VP.n51 VP.n9 0.189894
R1811 VP.n52 VP.n51 0.189894
R1812 VP.n53 VP.n52 0.189894
R1813 VP.n53 VP.n7 0.189894
R1814 VP.n58 VP.n7 0.189894
R1815 VP.n59 VP.n58 0.189894
R1816 VP.n60 VP.n59 0.189894
R1817 VP.n60 VP.n5 0.189894
R1818 VP.n64 VP.n5 0.189894
R1819 VP.n65 VP.n64 0.189894
R1820 VP.n65 VP.n3 0.189894
R1821 VP.n69 VP.n3 0.189894
R1822 VP.n70 VP.n69 0.189894
R1823 VP.n71 VP.n70 0.189894
R1824 VP.n71 VP.n1 0.189894
R1825 VP.n75 VP.n1 0.189894
R1826 VDD1 VDD1.n0 71.2645
R1827 VDD1.n3 VDD1.n2 71.1509
R1828 VDD1.n3 VDD1.n1 71.1509
R1829 VDD1.n5 VDD1.n4 69.7399
R1830 VDD1.n5 VDD1.n3 42.8328
R1831 VDD1.n4 VDD1.t3 3.19405
R1832 VDD1.n4 VDD1.t2 3.19405
R1833 VDD1.n0 VDD1.t6 3.19405
R1834 VDD1.n0 VDD1.t5 3.19405
R1835 VDD1.n2 VDD1.t1 3.19405
R1836 VDD1.n2 VDD1.t7 3.19405
R1837 VDD1.n1 VDD1.t0 3.19405
R1838 VDD1.n1 VDD1.t4 3.19405
R1839 VDD1 VDD1.n5 1.40783
C0 VTAIL VP 5.8829f
C1 VDD1 VN 0.152962f
C2 VDD2 VP 0.570068f
C3 VDD1 VTAIL 6.43458f
C4 VTAIL VN 5.8688f
C5 VDD1 VDD2 2.02259f
C6 VN VDD2 4.852109f
C7 VTAIL VDD2 6.49214f
C8 VDD1 VP 5.26758f
C9 VN VP 7.15978f
C10 VDD2 B 5.465888f
C11 VDD1 B 5.956802f
C12 VTAIL B 6.890757f
C13 VN B 16.70669f
C14 VP B 15.333453f
C15 VDD1.t6 B 0.141615f
C16 VDD1.t5 B 0.141615f
C17 VDD1.n0 B 1.21196f
C18 VDD1.t0 B 0.141615f
C19 VDD1.t4 B 0.141615f
C20 VDD1.n1 B 1.21074f
C21 VDD1.t1 B 0.141615f
C22 VDD1.t7 B 0.141615f
C23 VDD1.n2 B 1.21074f
C24 VDD1.n3 B 3.72228f
C25 VDD1.t3 B 0.141615f
C26 VDD1.t2 B 0.141615f
C27 VDD1.n4 B 1.19807f
C28 VDD1.n5 B 3.10469f
C29 VP.t0 B 1.16954f
C30 VP.n0 B 0.52159f
C31 VP.n1 B 0.023171f
C32 VP.n2 B 0.026338f
C33 VP.n3 B 0.023171f
C34 VP.t6 B 1.16954f
C35 VP.n4 B 0.433209f
C36 VP.n5 B 0.023171f
C37 VP.n6 B 0.033682f
C38 VP.n7 B 0.023171f
C39 VP.t3 B 1.16954f
C40 VP.n8 B 0.042968f
C41 VP.n9 B 0.023171f
C42 VP.n10 B 0.042968f
C43 VP.t5 B 1.16954f
C44 VP.n11 B 0.52159f
C45 VP.n12 B 0.023171f
C46 VP.n13 B 0.026338f
C47 VP.n14 B 0.023171f
C48 VP.t4 B 1.16954f
C49 VP.n15 B 0.433209f
C50 VP.n16 B 0.023171f
C51 VP.n17 B 0.033682f
C52 VP.n18 B 0.264696f
C53 VP.t2 B 1.16954f
C54 VP.t1 B 1.41077f
C55 VP.n19 B 0.485007f
C56 VP.n20 B 0.516487f
C57 VP.n21 B 0.040847f
C58 VP.n22 B 0.042968f
C59 VP.n23 B 0.023171f
C60 VP.n24 B 0.023171f
C61 VP.n25 B 0.023171f
C62 VP.n26 B 0.033682f
C63 VP.n27 B 0.042968f
C64 VP.n28 B 0.040847f
C65 VP.n29 B 0.023171f
C66 VP.n30 B 0.023171f
C67 VP.n31 B 0.023877f
C68 VP.n32 B 0.042968f
C69 VP.n33 B 0.044081f
C70 VP.n34 B 0.023171f
C71 VP.n35 B 0.023171f
C72 VP.n36 B 0.023171f
C73 VP.n37 B 0.039914f
C74 VP.n38 B 0.042968f
C75 VP.n39 B 0.036605f
C76 VP.n40 B 0.037391f
C77 VP.n41 B 1.26705f
C78 VP.n42 B 1.28417f
C79 VP.t7 B 1.16954f
C80 VP.n43 B 0.52159f
C81 VP.n44 B 0.036605f
C82 VP.n45 B 0.037391f
C83 VP.n46 B 0.023171f
C84 VP.n47 B 0.023171f
C85 VP.n48 B 0.039914f
C86 VP.n49 B 0.026338f
C87 VP.n50 B 0.044081f
C88 VP.n51 B 0.023171f
C89 VP.n52 B 0.023171f
C90 VP.n53 B 0.023171f
C91 VP.n54 B 0.023877f
C92 VP.n55 B 0.433209f
C93 VP.n56 B 0.040847f
C94 VP.n57 B 0.042968f
C95 VP.n58 B 0.023171f
C96 VP.n59 B 0.023171f
C97 VP.n60 B 0.023171f
C98 VP.n61 B 0.033682f
C99 VP.n62 B 0.042968f
C100 VP.n63 B 0.040847f
C101 VP.n64 B 0.023171f
C102 VP.n65 B 0.023171f
C103 VP.n66 B 0.023877f
C104 VP.n67 B 0.042968f
C105 VP.n68 B 0.044081f
C106 VP.n69 B 0.023171f
C107 VP.n70 B 0.023171f
C108 VP.n71 B 0.023171f
C109 VP.n72 B 0.039914f
C110 VP.n73 B 0.042968f
C111 VP.n74 B 0.036605f
C112 VP.n75 B 0.037391f
C113 VP.n76 B 0.051626f
C114 VTAIL.t14 B 0.116596f
C115 VTAIL.t8 B 0.116596f
C116 VTAIL.n0 B 0.930126f
C117 VTAIL.n1 B 0.436728f
C118 VTAIL.t13 B 1.18388f
C119 VTAIL.n2 B 0.532524f
C120 VTAIL.t3 B 1.18388f
C121 VTAIL.n3 B 0.532524f
C122 VTAIL.t2 B 0.116596f
C123 VTAIL.t7 B 0.116596f
C124 VTAIL.n4 B 0.930126f
C125 VTAIL.n5 B 0.657023f
C126 VTAIL.t6 B 1.18388f
C127 VTAIL.n6 B 1.45437f
C128 VTAIL.t11 B 1.18388f
C129 VTAIL.n7 B 1.45437f
C130 VTAIL.t10 B 0.116596f
C131 VTAIL.t15 B 0.116596f
C132 VTAIL.n8 B 0.93013f
C133 VTAIL.n9 B 0.657019f
C134 VTAIL.t9 B 1.18388f
C135 VTAIL.n10 B 0.532524f
C136 VTAIL.t5 B 1.18388f
C137 VTAIL.n11 B 0.532524f
C138 VTAIL.t1 B 0.116596f
C139 VTAIL.t4 B 0.116596f
C140 VTAIL.n12 B 0.93013f
C141 VTAIL.n13 B 0.657019f
C142 VTAIL.t0 B 1.18388f
C143 VTAIL.n14 B 1.45438f
C144 VTAIL.t12 B 1.18388f
C145 VTAIL.n15 B 1.44991f
C146 VDD2.t2 B 0.139602f
C147 VDD2.t5 B 0.139602f
C148 VDD2.n0 B 1.19353f
C149 VDD2.t1 B 0.139602f
C150 VDD2.t6 B 0.139602f
C151 VDD2.n1 B 1.19353f
C152 VDD2.n2 B 3.61012f
C153 VDD2.t7 B 0.139602f
C154 VDD2.t0 B 0.139602f
C155 VDD2.n3 B 1.18104f
C156 VDD2.n4 B 3.02524f
C157 VDD2.t4 B 0.139602f
C158 VDD2.t3 B 0.139602f
C159 VDD2.n5 B 1.19349f
C160 VN.t3 B 1.14209f
C161 VN.n0 B 0.509349f
C162 VN.n1 B 0.022627f
C163 VN.n2 B 0.02572f
C164 VN.n3 B 0.022627f
C165 VN.t7 B 1.14209f
C166 VN.n4 B 0.423042f
C167 VN.n5 B 0.022627f
C168 VN.n6 B 0.032892f
C169 VN.n7 B 0.258484f
C170 VN.t1 B 1.14209f
C171 VN.t2 B 1.37766f
C172 VN.n8 B 0.473624f
C173 VN.n9 B 0.504366f
C174 VN.n10 B 0.039888f
C175 VN.n11 B 0.04196f
C176 VN.n12 B 0.022627f
C177 VN.n13 B 0.022627f
C178 VN.n14 B 0.022627f
C179 VN.n15 B 0.032892f
C180 VN.n16 B 0.04196f
C181 VN.n17 B 0.039888f
C182 VN.n18 B 0.022627f
C183 VN.n19 B 0.022627f
C184 VN.n20 B 0.023317f
C185 VN.n21 B 0.04196f
C186 VN.n22 B 0.043046f
C187 VN.n23 B 0.022627f
C188 VN.n24 B 0.022627f
C189 VN.n25 B 0.022627f
C190 VN.n26 B 0.038978f
C191 VN.n27 B 0.04196f
C192 VN.n28 B 0.035746f
C193 VN.n29 B 0.036514f
C194 VN.n30 B 0.050414f
C195 VN.t4 B 1.14209f
C196 VN.n31 B 0.509349f
C197 VN.n32 B 0.022627f
C198 VN.n33 B 0.02572f
C199 VN.n34 B 0.022627f
C200 VN.t5 B 1.14209f
C201 VN.n35 B 0.423042f
C202 VN.n36 B 0.022627f
C203 VN.n37 B 0.032892f
C204 VN.n38 B 0.258484f
C205 VN.t0 B 1.14209f
C206 VN.t6 B 1.37766f
C207 VN.n39 B 0.473624f
C208 VN.n40 B 0.504366f
C209 VN.n41 B 0.039888f
C210 VN.n42 B 0.04196f
C211 VN.n43 B 0.022627f
C212 VN.n44 B 0.022627f
C213 VN.n45 B 0.022627f
C214 VN.n46 B 0.032892f
C215 VN.n47 B 0.04196f
C216 VN.n48 B 0.039888f
C217 VN.n49 B 0.022627f
C218 VN.n50 B 0.022627f
C219 VN.n51 B 0.023317f
C220 VN.n52 B 0.04196f
C221 VN.n53 B 0.043046f
C222 VN.n54 B 0.022627f
C223 VN.n55 B 0.022627f
C224 VN.n56 B 0.022627f
C225 VN.n57 B 0.038978f
C226 VN.n58 B 0.04196f
C227 VN.n59 B 0.035746f
C228 VN.n60 B 0.036514f
C229 VN.n61 B 1.24666f
.ends

