* NGSPICE file created from diff_pair_sample_0447.ext - technology: sky130A

.subckt diff_pair_sample_0447 VTAIL VN VP B VDD2 VDD1
X0 B.t21 B.t19 B.t20 B.t13 sky130_fd_pr__nfet_01v8 ad=3.9468 pd=21.02 as=0 ps=0 w=10.12 l=2.17
X1 VTAIL.t15 VN.t0 VDD2.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=1.6698 pd=10.45 as=1.6698 ps=10.45 w=10.12 l=2.17
X2 VTAIL.t4 VP.t0 VDD1.t7 B.t5 sky130_fd_pr__nfet_01v8 ad=1.6698 pd=10.45 as=1.6698 ps=10.45 w=10.12 l=2.17
X3 VTAIL.t14 VN.t1 VDD2.t4 B.t7 sky130_fd_pr__nfet_01v8 ad=3.9468 pd=21.02 as=1.6698 ps=10.45 w=10.12 l=2.17
X4 VTAIL.t7 VP.t1 VDD1.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=3.9468 pd=21.02 as=1.6698 ps=10.45 w=10.12 l=2.17
X5 VTAIL.t6 VP.t2 VDD1.t5 B.t7 sky130_fd_pr__nfet_01v8 ad=3.9468 pd=21.02 as=1.6698 ps=10.45 w=10.12 l=2.17
X6 VDD2.t0 VN.t2 VTAIL.t13 B.t4 sky130_fd_pr__nfet_01v8 ad=1.6698 pd=10.45 as=3.9468 ps=21.02 w=10.12 l=2.17
X7 VDD2.t5 VN.t3 VTAIL.t12 B.t2 sky130_fd_pr__nfet_01v8 ad=1.6698 pd=10.45 as=1.6698 ps=10.45 w=10.12 l=2.17
X8 VDD1.t4 VP.t3 VTAIL.t3 B.t4 sky130_fd_pr__nfet_01v8 ad=1.6698 pd=10.45 as=3.9468 ps=21.02 w=10.12 l=2.17
X9 VTAIL.t1 VP.t4 VDD1.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=1.6698 pd=10.45 as=1.6698 ps=10.45 w=10.12 l=2.17
X10 B.t18 B.t16 B.t17 B.t9 sky130_fd_pr__nfet_01v8 ad=3.9468 pd=21.02 as=0 ps=0 w=10.12 l=2.17
X11 VDD2.t6 VN.t4 VTAIL.t11 B.t0 sky130_fd_pr__nfet_01v8 ad=1.6698 pd=10.45 as=3.9468 ps=21.02 w=10.12 l=2.17
X12 VDD1.t2 VP.t5 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.6698 pd=10.45 as=1.6698 ps=10.45 w=10.12 l=2.17
X13 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=3.9468 pd=21.02 as=0 ps=0 w=10.12 l=2.17
X14 VDD2.t2 VN.t5 VTAIL.t10 B.t6 sky130_fd_pr__nfet_01v8 ad=1.6698 pd=10.45 as=1.6698 ps=10.45 w=10.12 l=2.17
X15 VDD1.t1 VP.t6 VTAIL.t5 B.t6 sky130_fd_pr__nfet_01v8 ad=1.6698 pd=10.45 as=1.6698 ps=10.45 w=10.12 l=2.17
X16 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=3.9468 pd=21.02 as=0 ps=0 w=10.12 l=2.17
X17 VTAIL.t9 VN.t6 VDD2.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=3.9468 pd=21.02 as=1.6698 ps=10.45 w=10.12 l=2.17
X18 VDD1.t0 VP.t7 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.6698 pd=10.45 as=3.9468 ps=21.02 w=10.12 l=2.17
X19 VTAIL.t8 VN.t7 VDD2.t7 B.t5 sky130_fd_pr__nfet_01v8 ad=1.6698 pd=10.45 as=1.6698 ps=10.45 w=10.12 l=2.17
R0 B.n783 B.n782 585
R1 B.n291 B.n124 585
R2 B.n290 B.n289 585
R3 B.n288 B.n287 585
R4 B.n286 B.n285 585
R5 B.n284 B.n283 585
R6 B.n282 B.n281 585
R7 B.n280 B.n279 585
R8 B.n278 B.n277 585
R9 B.n276 B.n275 585
R10 B.n274 B.n273 585
R11 B.n272 B.n271 585
R12 B.n270 B.n269 585
R13 B.n268 B.n267 585
R14 B.n266 B.n265 585
R15 B.n264 B.n263 585
R16 B.n262 B.n261 585
R17 B.n260 B.n259 585
R18 B.n258 B.n257 585
R19 B.n256 B.n255 585
R20 B.n254 B.n253 585
R21 B.n252 B.n251 585
R22 B.n250 B.n249 585
R23 B.n248 B.n247 585
R24 B.n246 B.n245 585
R25 B.n244 B.n243 585
R26 B.n242 B.n241 585
R27 B.n240 B.n239 585
R28 B.n238 B.n237 585
R29 B.n236 B.n235 585
R30 B.n234 B.n233 585
R31 B.n232 B.n231 585
R32 B.n230 B.n229 585
R33 B.n228 B.n227 585
R34 B.n226 B.n225 585
R35 B.n224 B.n223 585
R36 B.n222 B.n221 585
R37 B.n220 B.n219 585
R38 B.n218 B.n217 585
R39 B.n216 B.n215 585
R40 B.n214 B.n213 585
R41 B.n212 B.n211 585
R42 B.n210 B.n209 585
R43 B.n208 B.n207 585
R44 B.n206 B.n205 585
R45 B.n204 B.n203 585
R46 B.n202 B.n201 585
R47 B.n200 B.n199 585
R48 B.n198 B.n197 585
R49 B.n196 B.n195 585
R50 B.n194 B.n193 585
R51 B.n192 B.n191 585
R52 B.n190 B.n189 585
R53 B.n188 B.n187 585
R54 B.n186 B.n185 585
R55 B.n184 B.n183 585
R56 B.n182 B.n181 585
R57 B.n180 B.n179 585
R58 B.n178 B.n177 585
R59 B.n176 B.n175 585
R60 B.n174 B.n173 585
R61 B.n172 B.n171 585
R62 B.n170 B.n169 585
R63 B.n168 B.n167 585
R64 B.n166 B.n165 585
R65 B.n164 B.n163 585
R66 B.n162 B.n161 585
R67 B.n160 B.n159 585
R68 B.n158 B.n157 585
R69 B.n156 B.n155 585
R70 B.n154 B.n153 585
R71 B.n152 B.n151 585
R72 B.n150 B.n149 585
R73 B.n148 B.n147 585
R74 B.n146 B.n145 585
R75 B.n144 B.n143 585
R76 B.n142 B.n141 585
R77 B.n140 B.n139 585
R78 B.n138 B.n137 585
R79 B.n136 B.n135 585
R80 B.n134 B.n133 585
R81 B.n132 B.n131 585
R82 B.n781 B.n83 585
R83 B.n786 B.n83 585
R84 B.n780 B.n82 585
R85 B.n787 B.n82 585
R86 B.n779 B.n778 585
R87 B.n778 B.n78 585
R88 B.n777 B.n77 585
R89 B.n793 B.n77 585
R90 B.n776 B.n76 585
R91 B.n794 B.n76 585
R92 B.n775 B.n75 585
R93 B.n795 B.n75 585
R94 B.n774 B.n773 585
R95 B.n773 B.n71 585
R96 B.n772 B.n70 585
R97 B.n801 B.n70 585
R98 B.n771 B.n69 585
R99 B.n802 B.n69 585
R100 B.n770 B.n68 585
R101 B.n803 B.n68 585
R102 B.n769 B.n768 585
R103 B.n768 B.n64 585
R104 B.n767 B.n63 585
R105 B.n809 B.n63 585
R106 B.n766 B.n62 585
R107 B.n810 B.n62 585
R108 B.n765 B.n61 585
R109 B.n811 B.n61 585
R110 B.n764 B.n763 585
R111 B.n763 B.n57 585
R112 B.n762 B.n56 585
R113 B.n817 B.n56 585
R114 B.n761 B.n55 585
R115 B.n818 B.n55 585
R116 B.n760 B.n54 585
R117 B.n819 B.n54 585
R118 B.n759 B.n758 585
R119 B.n758 B.n50 585
R120 B.n757 B.n49 585
R121 B.n825 B.n49 585
R122 B.n756 B.n48 585
R123 B.n826 B.n48 585
R124 B.n755 B.n47 585
R125 B.n827 B.n47 585
R126 B.n754 B.n753 585
R127 B.n753 B.n43 585
R128 B.n752 B.n42 585
R129 B.n833 B.n42 585
R130 B.n751 B.n41 585
R131 B.n834 B.n41 585
R132 B.n750 B.n40 585
R133 B.n835 B.n40 585
R134 B.n749 B.n748 585
R135 B.n748 B.n36 585
R136 B.n747 B.n35 585
R137 B.n841 B.n35 585
R138 B.n746 B.n34 585
R139 B.n842 B.n34 585
R140 B.n745 B.n33 585
R141 B.n843 B.n33 585
R142 B.n744 B.n743 585
R143 B.n743 B.n29 585
R144 B.n742 B.n28 585
R145 B.n849 B.n28 585
R146 B.n741 B.n27 585
R147 B.n850 B.n27 585
R148 B.n740 B.n26 585
R149 B.n851 B.n26 585
R150 B.n739 B.n738 585
R151 B.n738 B.n22 585
R152 B.n737 B.n21 585
R153 B.n857 B.n21 585
R154 B.n736 B.n20 585
R155 B.n858 B.n20 585
R156 B.n735 B.n19 585
R157 B.n859 B.n19 585
R158 B.n734 B.n733 585
R159 B.n733 B.n15 585
R160 B.n732 B.n14 585
R161 B.n865 B.n14 585
R162 B.n731 B.n13 585
R163 B.n866 B.n13 585
R164 B.n730 B.n12 585
R165 B.n867 B.n12 585
R166 B.n729 B.n728 585
R167 B.n728 B.n8 585
R168 B.n727 B.n7 585
R169 B.n873 B.n7 585
R170 B.n726 B.n6 585
R171 B.n874 B.n6 585
R172 B.n725 B.n5 585
R173 B.n875 B.n5 585
R174 B.n724 B.n723 585
R175 B.n723 B.n4 585
R176 B.n722 B.n292 585
R177 B.n722 B.n721 585
R178 B.n712 B.n293 585
R179 B.n294 B.n293 585
R180 B.n714 B.n713 585
R181 B.n715 B.n714 585
R182 B.n711 B.n299 585
R183 B.n299 B.n298 585
R184 B.n710 B.n709 585
R185 B.n709 B.n708 585
R186 B.n301 B.n300 585
R187 B.n302 B.n301 585
R188 B.n701 B.n700 585
R189 B.n702 B.n701 585
R190 B.n699 B.n307 585
R191 B.n307 B.n306 585
R192 B.n698 B.n697 585
R193 B.n697 B.n696 585
R194 B.n309 B.n308 585
R195 B.n310 B.n309 585
R196 B.n689 B.n688 585
R197 B.n690 B.n689 585
R198 B.n687 B.n314 585
R199 B.n318 B.n314 585
R200 B.n686 B.n685 585
R201 B.n685 B.n684 585
R202 B.n316 B.n315 585
R203 B.n317 B.n316 585
R204 B.n677 B.n676 585
R205 B.n678 B.n677 585
R206 B.n675 B.n323 585
R207 B.n323 B.n322 585
R208 B.n674 B.n673 585
R209 B.n673 B.n672 585
R210 B.n325 B.n324 585
R211 B.n326 B.n325 585
R212 B.n665 B.n664 585
R213 B.n666 B.n665 585
R214 B.n663 B.n331 585
R215 B.n331 B.n330 585
R216 B.n662 B.n661 585
R217 B.n661 B.n660 585
R218 B.n333 B.n332 585
R219 B.n334 B.n333 585
R220 B.n653 B.n652 585
R221 B.n654 B.n653 585
R222 B.n651 B.n339 585
R223 B.n339 B.n338 585
R224 B.n650 B.n649 585
R225 B.n649 B.n648 585
R226 B.n341 B.n340 585
R227 B.n342 B.n341 585
R228 B.n641 B.n640 585
R229 B.n642 B.n641 585
R230 B.n639 B.n347 585
R231 B.n347 B.n346 585
R232 B.n638 B.n637 585
R233 B.n637 B.n636 585
R234 B.n349 B.n348 585
R235 B.n350 B.n349 585
R236 B.n629 B.n628 585
R237 B.n630 B.n629 585
R238 B.n627 B.n355 585
R239 B.n355 B.n354 585
R240 B.n626 B.n625 585
R241 B.n625 B.n624 585
R242 B.n357 B.n356 585
R243 B.n358 B.n357 585
R244 B.n617 B.n616 585
R245 B.n618 B.n617 585
R246 B.n615 B.n363 585
R247 B.n363 B.n362 585
R248 B.n614 B.n613 585
R249 B.n613 B.n612 585
R250 B.n365 B.n364 585
R251 B.n366 B.n365 585
R252 B.n605 B.n604 585
R253 B.n606 B.n605 585
R254 B.n603 B.n371 585
R255 B.n371 B.n370 585
R256 B.n602 B.n601 585
R257 B.n601 B.n600 585
R258 B.n373 B.n372 585
R259 B.n374 B.n373 585
R260 B.n593 B.n592 585
R261 B.n594 B.n593 585
R262 B.n591 B.n379 585
R263 B.n379 B.n378 585
R264 B.n586 B.n585 585
R265 B.n584 B.n422 585
R266 B.n583 B.n421 585
R267 B.n588 B.n421 585
R268 B.n582 B.n581 585
R269 B.n580 B.n579 585
R270 B.n578 B.n577 585
R271 B.n576 B.n575 585
R272 B.n574 B.n573 585
R273 B.n572 B.n571 585
R274 B.n570 B.n569 585
R275 B.n568 B.n567 585
R276 B.n566 B.n565 585
R277 B.n564 B.n563 585
R278 B.n562 B.n561 585
R279 B.n560 B.n559 585
R280 B.n558 B.n557 585
R281 B.n556 B.n555 585
R282 B.n554 B.n553 585
R283 B.n552 B.n551 585
R284 B.n550 B.n549 585
R285 B.n548 B.n547 585
R286 B.n546 B.n545 585
R287 B.n544 B.n543 585
R288 B.n542 B.n541 585
R289 B.n540 B.n539 585
R290 B.n538 B.n537 585
R291 B.n536 B.n535 585
R292 B.n534 B.n533 585
R293 B.n532 B.n531 585
R294 B.n530 B.n529 585
R295 B.n528 B.n527 585
R296 B.n526 B.n525 585
R297 B.n524 B.n523 585
R298 B.n522 B.n521 585
R299 B.n520 B.n519 585
R300 B.n518 B.n517 585
R301 B.n515 B.n514 585
R302 B.n513 B.n512 585
R303 B.n511 B.n510 585
R304 B.n509 B.n508 585
R305 B.n507 B.n506 585
R306 B.n505 B.n504 585
R307 B.n503 B.n502 585
R308 B.n501 B.n500 585
R309 B.n499 B.n498 585
R310 B.n497 B.n496 585
R311 B.n494 B.n493 585
R312 B.n492 B.n491 585
R313 B.n490 B.n489 585
R314 B.n488 B.n487 585
R315 B.n486 B.n485 585
R316 B.n484 B.n483 585
R317 B.n482 B.n481 585
R318 B.n480 B.n479 585
R319 B.n478 B.n477 585
R320 B.n476 B.n475 585
R321 B.n474 B.n473 585
R322 B.n472 B.n471 585
R323 B.n470 B.n469 585
R324 B.n468 B.n467 585
R325 B.n466 B.n465 585
R326 B.n464 B.n463 585
R327 B.n462 B.n461 585
R328 B.n460 B.n459 585
R329 B.n458 B.n457 585
R330 B.n456 B.n455 585
R331 B.n454 B.n453 585
R332 B.n452 B.n451 585
R333 B.n450 B.n449 585
R334 B.n448 B.n447 585
R335 B.n446 B.n445 585
R336 B.n444 B.n443 585
R337 B.n442 B.n441 585
R338 B.n440 B.n439 585
R339 B.n438 B.n437 585
R340 B.n436 B.n435 585
R341 B.n434 B.n433 585
R342 B.n432 B.n431 585
R343 B.n430 B.n429 585
R344 B.n428 B.n427 585
R345 B.n381 B.n380 585
R346 B.n590 B.n589 585
R347 B.n589 B.n588 585
R348 B.n377 B.n376 585
R349 B.n378 B.n377 585
R350 B.n596 B.n595 585
R351 B.n595 B.n594 585
R352 B.n597 B.n375 585
R353 B.n375 B.n374 585
R354 B.n599 B.n598 585
R355 B.n600 B.n599 585
R356 B.n369 B.n368 585
R357 B.n370 B.n369 585
R358 B.n608 B.n607 585
R359 B.n607 B.n606 585
R360 B.n609 B.n367 585
R361 B.n367 B.n366 585
R362 B.n611 B.n610 585
R363 B.n612 B.n611 585
R364 B.n361 B.n360 585
R365 B.n362 B.n361 585
R366 B.n620 B.n619 585
R367 B.n619 B.n618 585
R368 B.n621 B.n359 585
R369 B.n359 B.n358 585
R370 B.n623 B.n622 585
R371 B.n624 B.n623 585
R372 B.n353 B.n352 585
R373 B.n354 B.n353 585
R374 B.n632 B.n631 585
R375 B.n631 B.n630 585
R376 B.n633 B.n351 585
R377 B.n351 B.n350 585
R378 B.n635 B.n634 585
R379 B.n636 B.n635 585
R380 B.n345 B.n344 585
R381 B.n346 B.n345 585
R382 B.n644 B.n643 585
R383 B.n643 B.n642 585
R384 B.n645 B.n343 585
R385 B.n343 B.n342 585
R386 B.n647 B.n646 585
R387 B.n648 B.n647 585
R388 B.n337 B.n336 585
R389 B.n338 B.n337 585
R390 B.n656 B.n655 585
R391 B.n655 B.n654 585
R392 B.n657 B.n335 585
R393 B.n335 B.n334 585
R394 B.n659 B.n658 585
R395 B.n660 B.n659 585
R396 B.n329 B.n328 585
R397 B.n330 B.n329 585
R398 B.n668 B.n667 585
R399 B.n667 B.n666 585
R400 B.n669 B.n327 585
R401 B.n327 B.n326 585
R402 B.n671 B.n670 585
R403 B.n672 B.n671 585
R404 B.n321 B.n320 585
R405 B.n322 B.n321 585
R406 B.n680 B.n679 585
R407 B.n679 B.n678 585
R408 B.n681 B.n319 585
R409 B.n319 B.n317 585
R410 B.n683 B.n682 585
R411 B.n684 B.n683 585
R412 B.n313 B.n312 585
R413 B.n318 B.n313 585
R414 B.n692 B.n691 585
R415 B.n691 B.n690 585
R416 B.n693 B.n311 585
R417 B.n311 B.n310 585
R418 B.n695 B.n694 585
R419 B.n696 B.n695 585
R420 B.n305 B.n304 585
R421 B.n306 B.n305 585
R422 B.n704 B.n703 585
R423 B.n703 B.n702 585
R424 B.n705 B.n303 585
R425 B.n303 B.n302 585
R426 B.n707 B.n706 585
R427 B.n708 B.n707 585
R428 B.n297 B.n296 585
R429 B.n298 B.n297 585
R430 B.n717 B.n716 585
R431 B.n716 B.n715 585
R432 B.n718 B.n295 585
R433 B.n295 B.n294 585
R434 B.n720 B.n719 585
R435 B.n721 B.n720 585
R436 B.n2 B.n0 585
R437 B.n4 B.n2 585
R438 B.n3 B.n1 585
R439 B.n874 B.n3 585
R440 B.n872 B.n871 585
R441 B.n873 B.n872 585
R442 B.n870 B.n9 585
R443 B.n9 B.n8 585
R444 B.n869 B.n868 585
R445 B.n868 B.n867 585
R446 B.n11 B.n10 585
R447 B.n866 B.n11 585
R448 B.n864 B.n863 585
R449 B.n865 B.n864 585
R450 B.n862 B.n16 585
R451 B.n16 B.n15 585
R452 B.n861 B.n860 585
R453 B.n860 B.n859 585
R454 B.n18 B.n17 585
R455 B.n858 B.n18 585
R456 B.n856 B.n855 585
R457 B.n857 B.n856 585
R458 B.n854 B.n23 585
R459 B.n23 B.n22 585
R460 B.n853 B.n852 585
R461 B.n852 B.n851 585
R462 B.n25 B.n24 585
R463 B.n850 B.n25 585
R464 B.n848 B.n847 585
R465 B.n849 B.n848 585
R466 B.n846 B.n30 585
R467 B.n30 B.n29 585
R468 B.n845 B.n844 585
R469 B.n844 B.n843 585
R470 B.n32 B.n31 585
R471 B.n842 B.n32 585
R472 B.n840 B.n839 585
R473 B.n841 B.n840 585
R474 B.n838 B.n37 585
R475 B.n37 B.n36 585
R476 B.n837 B.n836 585
R477 B.n836 B.n835 585
R478 B.n39 B.n38 585
R479 B.n834 B.n39 585
R480 B.n832 B.n831 585
R481 B.n833 B.n832 585
R482 B.n830 B.n44 585
R483 B.n44 B.n43 585
R484 B.n829 B.n828 585
R485 B.n828 B.n827 585
R486 B.n46 B.n45 585
R487 B.n826 B.n46 585
R488 B.n824 B.n823 585
R489 B.n825 B.n824 585
R490 B.n822 B.n51 585
R491 B.n51 B.n50 585
R492 B.n821 B.n820 585
R493 B.n820 B.n819 585
R494 B.n53 B.n52 585
R495 B.n818 B.n53 585
R496 B.n816 B.n815 585
R497 B.n817 B.n816 585
R498 B.n814 B.n58 585
R499 B.n58 B.n57 585
R500 B.n813 B.n812 585
R501 B.n812 B.n811 585
R502 B.n60 B.n59 585
R503 B.n810 B.n60 585
R504 B.n808 B.n807 585
R505 B.n809 B.n808 585
R506 B.n806 B.n65 585
R507 B.n65 B.n64 585
R508 B.n805 B.n804 585
R509 B.n804 B.n803 585
R510 B.n67 B.n66 585
R511 B.n802 B.n67 585
R512 B.n800 B.n799 585
R513 B.n801 B.n800 585
R514 B.n798 B.n72 585
R515 B.n72 B.n71 585
R516 B.n797 B.n796 585
R517 B.n796 B.n795 585
R518 B.n74 B.n73 585
R519 B.n794 B.n74 585
R520 B.n792 B.n791 585
R521 B.n793 B.n792 585
R522 B.n790 B.n79 585
R523 B.n79 B.n78 585
R524 B.n789 B.n788 585
R525 B.n788 B.n787 585
R526 B.n81 B.n80 585
R527 B.n786 B.n81 585
R528 B.n877 B.n876 585
R529 B.n876 B.n875 585
R530 B.n586 B.n377 458.866
R531 B.n131 B.n81 458.866
R532 B.n589 B.n379 458.866
R533 B.n783 B.n83 458.866
R534 B.n425 B.t12 319.683
R535 B.n423 B.t19 319.683
R536 B.n128 B.t16 319.683
R537 B.n125 B.t8 319.683
R538 B.n425 B.t15 298.459
R539 B.n125 B.t10 298.459
R540 B.n423 B.t21 298.459
R541 B.n128 B.t17 298.459
R542 B.n785 B.n784 256.663
R543 B.n785 B.n123 256.663
R544 B.n785 B.n122 256.663
R545 B.n785 B.n121 256.663
R546 B.n785 B.n120 256.663
R547 B.n785 B.n119 256.663
R548 B.n785 B.n118 256.663
R549 B.n785 B.n117 256.663
R550 B.n785 B.n116 256.663
R551 B.n785 B.n115 256.663
R552 B.n785 B.n114 256.663
R553 B.n785 B.n113 256.663
R554 B.n785 B.n112 256.663
R555 B.n785 B.n111 256.663
R556 B.n785 B.n110 256.663
R557 B.n785 B.n109 256.663
R558 B.n785 B.n108 256.663
R559 B.n785 B.n107 256.663
R560 B.n785 B.n106 256.663
R561 B.n785 B.n105 256.663
R562 B.n785 B.n104 256.663
R563 B.n785 B.n103 256.663
R564 B.n785 B.n102 256.663
R565 B.n785 B.n101 256.663
R566 B.n785 B.n100 256.663
R567 B.n785 B.n99 256.663
R568 B.n785 B.n98 256.663
R569 B.n785 B.n97 256.663
R570 B.n785 B.n96 256.663
R571 B.n785 B.n95 256.663
R572 B.n785 B.n94 256.663
R573 B.n785 B.n93 256.663
R574 B.n785 B.n92 256.663
R575 B.n785 B.n91 256.663
R576 B.n785 B.n90 256.663
R577 B.n785 B.n89 256.663
R578 B.n785 B.n88 256.663
R579 B.n785 B.n87 256.663
R580 B.n785 B.n86 256.663
R581 B.n785 B.n85 256.663
R582 B.n785 B.n84 256.663
R583 B.n588 B.n587 256.663
R584 B.n588 B.n382 256.663
R585 B.n588 B.n383 256.663
R586 B.n588 B.n384 256.663
R587 B.n588 B.n385 256.663
R588 B.n588 B.n386 256.663
R589 B.n588 B.n387 256.663
R590 B.n588 B.n388 256.663
R591 B.n588 B.n389 256.663
R592 B.n588 B.n390 256.663
R593 B.n588 B.n391 256.663
R594 B.n588 B.n392 256.663
R595 B.n588 B.n393 256.663
R596 B.n588 B.n394 256.663
R597 B.n588 B.n395 256.663
R598 B.n588 B.n396 256.663
R599 B.n588 B.n397 256.663
R600 B.n588 B.n398 256.663
R601 B.n588 B.n399 256.663
R602 B.n588 B.n400 256.663
R603 B.n588 B.n401 256.663
R604 B.n588 B.n402 256.663
R605 B.n588 B.n403 256.663
R606 B.n588 B.n404 256.663
R607 B.n588 B.n405 256.663
R608 B.n588 B.n406 256.663
R609 B.n588 B.n407 256.663
R610 B.n588 B.n408 256.663
R611 B.n588 B.n409 256.663
R612 B.n588 B.n410 256.663
R613 B.n588 B.n411 256.663
R614 B.n588 B.n412 256.663
R615 B.n588 B.n413 256.663
R616 B.n588 B.n414 256.663
R617 B.n588 B.n415 256.663
R618 B.n588 B.n416 256.663
R619 B.n588 B.n417 256.663
R620 B.n588 B.n418 256.663
R621 B.n588 B.n419 256.663
R622 B.n588 B.n420 256.663
R623 B.n426 B.t14 249.975
R624 B.n126 B.t11 249.975
R625 B.n424 B.t20 249.975
R626 B.n129 B.t18 249.975
R627 B.n595 B.n377 163.367
R628 B.n595 B.n375 163.367
R629 B.n599 B.n375 163.367
R630 B.n599 B.n369 163.367
R631 B.n607 B.n369 163.367
R632 B.n607 B.n367 163.367
R633 B.n611 B.n367 163.367
R634 B.n611 B.n361 163.367
R635 B.n619 B.n361 163.367
R636 B.n619 B.n359 163.367
R637 B.n623 B.n359 163.367
R638 B.n623 B.n353 163.367
R639 B.n631 B.n353 163.367
R640 B.n631 B.n351 163.367
R641 B.n635 B.n351 163.367
R642 B.n635 B.n345 163.367
R643 B.n643 B.n345 163.367
R644 B.n643 B.n343 163.367
R645 B.n647 B.n343 163.367
R646 B.n647 B.n337 163.367
R647 B.n655 B.n337 163.367
R648 B.n655 B.n335 163.367
R649 B.n659 B.n335 163.367
R650 B.n659 B.n329 163.367
R651 B.n667 B.n329 163.367
R652 B.n667 B.n327 163.367
R653 B.n671 B.n327 163.367
R654 B.n671 B.n321 163.367
R655 B.n679 B.n321 163.367
R656 B.n679 B.n319 163.367
R657 B.n683 B.n319 163.367
R658 B.n683 B.n313 163.367
R659 B.n691 B.n313 163.367
R660 B.n691 B.n311 163.367
R661 B.n695 B.n311 163.367
R662 B.n695 B.n305 163.367
R663 B.n703 B.n305 163.367
R664 B.n703 B.n303 163.367
R665 B.n707 B.n303 163.367
R666 B.n707 B.n297 163.367
R667 B.n716 B.n297 163.367
R668 B.n716 B.n295 163.367
R669 B.n720 B.n295 163.367
R670 B.n720 B.n2 163.367
R671 B.n876 B.n2 163.367
R672 B.n876 B.n3 163.367
R673 B.n872 B.n3 163.367
R674 B.n872 B.n9 163.367
R675 B.n868 B.n9 163.367
R676 B.n868 B.n11 163.367
R677 B.n864 B.n11 163.367
R678 B.n864 B.n16 163.367
R679 B.n860 B.n16 163.367
R680 B.n860 B.n18 163.367
R681 B.n856 B.n18 163.367
R682 B.n856 B.n23 163.367
R683 B.n852 B.n23 163.367
R684 B.n852 B.n25 163.367
R685 B.n848 B.n25 163.367
R686 B.n848 B.n30 163.367
R687 B.n844 B.n30 163.367
R688 B.n844 B.n32 163.367
R689 B.n840 B.n32 163.367
R690 B.n840 B.n37 163.367
R691 B.n836 B.n37 163.367
R692 B.n836 B.n39 163.367
R693 B.n832 B.n39 163.367
R694 B.n832 B.n44 163.367
R695 B.n828 B.n44 163.367
R696 B.n828 B.n46 163.367
R697 B.n824 B.n46 163.367
R698 B.n824 B.n51 163.367
R699 B.n820 B.n51 163.367
R700 B.n820 B.n53 163.367
R701 B.n816 B.n53 163.367
R702 B.n816 B.n58 163.367
R703 B.n812 B.n58 163.367
R704 B.n812 B.n60 163.367
R705 B.n808 B.n60 163.367
R706 B.n808 B.n65 163.367
R707 B.n804 B.n65 163.367
R708 B.n804 B.n67 163.367
R709 B.n800 B.n67 163.367
R710 B.n800 B.n72 163.367
R711 B.n796 B.n72 163.367
R712 B.n796 B.n74 163.367
R713 B.n792 B.n74 163.367
R714 B.n792 B.n79 163.367
R715 B.n788 B.n79 163.367
R716 B.n788 B.n81 163.367
R717 B.n422 B.n421 163.367
R718 B.n581 B.n421 163.367
R719 B.n579 B.n578 163.367
R720 B.n575 B.n574 163.367
R721 B.n571 B.n570 163.367
R722 B.n567 B.n566 163.367
R723 B.n563 B.n562 163.367
R724 B.n559 B.n558 163.367
R725 B.n555 B.n554 163.367
R726 B.n551 B.n550 163.367
R727 B.n547 B.n546 163.367
R728 B.n543 B.n542 163.367
R729 B.n539 B.n538 163.367
R730 B.n535 B.n534 163.367
R731 B.n531 B.n530 163.367
R732 B.n527 B.n526 163.367
R733 B.n523 B.n522 163.367
R734 B.n519 B.n518 163.367
R735 B.n514 B.n513 163.367
R736 B.n510 B.n509 163.367
R737 B.n506 B.n505 163.367
R738 B.n502 B.n501 163.367
R739 B.n498 B.n497 163.367
R740 B.n493 B.n492 163.367
R741 B.n489 B.n488 163.367
R742 B.n485 B.n484 163.367
R743 B.n481 B.n480 163.367
R744 B.n477 B.n476 163.367
R745 B.n473 B.n472 163.367
R746 B.n469 B.n468 163.367
R747 B.n465 B.n464 163.367
R748 B.n461 B.n460 163.367
R749 B.n457 B.n456 163.367
R750 B.n453 B.n452 163.367
R751 B.n449 B.n448 163.367
R752 B.n445 B.n444 163.367
R753 B.n441 B.n440 163.367
R754 B.n437 B.n436 163.367
R755 B.n433 B.n432 163.367
R756 B.n429 B.n428 163.367
R757 B.n589 B.n381 163.367
R758 B.n593 B.n379 163.367
R759 B.n593 B.n373 163.367
R760 B.n601 B.n373 163.367
R761 B.n601 B.n371 163.367
R762 B.n605 B.n371 163.367
R763 B.n605 B.n365 163.367
R764 B.n613 B.n365 163.367
R765 B.n613 B.n363 163.367
R766 B.n617 B.n363 163.367
R767 B.n617 B.n357 163.367
R768 B.n625 B.n357 163.367
R769 B.n625 B.n355 163.367
R770 B.n629 B.n355 163.367
R771 B.n629 B.n349 163.367
R772 B.n637 B.n349 163.367
R773 B.n637 B.n347 163.367
R774 B.n641 B.n347 163.367
R775 B.n641 B.n341 163.367
R776 B.n649 B.n341 163.367
R777 B.n649 B.n339 163.367
R778 B.n653 B.n339 163.367
R779 B.n653 B.n333 163.367
R780 B.n661 B.n333 163.367
R781 B.n661 B.n331 163.367
R782 B.n665 B.n331 163.367
R783 B.n665 B.n325 163.367
R784 B.n673 B.n325 163.367
R785 B.n673 B.n323 163.367
R786 B.n677 B.n323 163.367
R787 B.n677 B.n316 163.367
R788 B.n685 B.n316 163.367
R789 B.n685 B.n314 163.367
R790 B.n689 B.n314 163.367
R791 B.n689 B.n309 163.367
R792 B.n697 B.n309 163.367
R793 B.n697 B.n307 163.367
R794 B.n701 B.n307 163.367
R795 B.n701 B.n301 163.367
R796 B.n709 B.n301 163.367
R797 B.n709 B.n299 163.367
R798 B.n714 B.n299 163.367
R799 B.n714 B.n293 163.367
R800 B.n722 B.n293 163.367
R801 B.n723 B.n722 163.367
R802 B.n723 B.n5 163.367
R803 B.n6 B.n5 163.367
R804 B.n7 B.n6 163.367
R805 B.n728 B.n7 163.367
R806 B.n728 B.n12 163.367
R807 B.n13 B.n12 163.367
R808 B.n14 B.n13 163.367
R809 B.n733 B.n14 163.367
R810 B.n733 B.n19 163.367
R811 B.n20 B.n19 163.367
R812 B.n21 B.n20 163.367
R813 B.n738 B.n21 163.367
R814 B.n738 B.n26 163.367
R815 B.n27 B.n26 163.367
R816 B.n28 B.n27 163.367
R817 B.n743 B.n28 163.367
R818 B.n743 B.n33 163.367
R819 B.n34 B.n33 163.367
R820 B.n35 B.n34 163.367
R821 B.n748 B.n35 163.367
R822 B.n748 B.n40 163.367
R823 B.n41 B.n40 163.367
R824 B.n42 B.n41 163.367
R825 B.n753 B.n42 163.367
R826 B.n753 B.n47 163.367
R827 B.n48 B.n47 163.367
R828 B.n49 B.n48 163.367
R829 B.n758 B.n49 163.367
R830 B.n758 B.n54 163.367
R831 B.n55 B.n54 163.367
R832 B.n56 B.n55 163.367
R833 B.n763 B.n56 163.367
R834 B.n763 B.n61 163.367
R835 B.n62 B.n61 163.367
R836 B.n63 B.n62 163.367
R837 B.n768 B.n63 163.367
R838 B.n768 B.n68 163.367
R839 B.n69 B.n68 163.367
R840 B.n70 B.n69 163.367
R841 B.n773 B.n70 163.367
R842 B.n773 B.n75 163.367
R843 B.n76 B.n75 163.367
R844 B.n77 B.n76 163.367
R845 B.n778 B.n77 163.367
R846 B.n778 B.n82 163.367
R847 B.n83 B.n82 163.367
R848 B.n135 B.n134 163.367
R849 B.n139 B.n138 163.367
R850 B.n143 B.n142 163.367
R851 B.n147 B.n146 163.367
R852 B.n151 B.n150 163.367
R853 B.n155 B.n154 163.367
R854 B.n159 B.n158 163.367
R855 B.n163 B.n162 163.367
R856 B.n167 B.n166 163.367
R857 B.n171 B.n170 163.367
R858 B.n175 B.n174 163.367
R859 B.n179 B.n178 163.367
R860 B.n183 B.n182 163.367
R861 B.n187 B.n186 163.367
R862 B.n191 B.n190 163.367
R863 B.n195 B.n194 163.367
R864 B.n199 B.n198 163.367
R865 B.n203 B.n202 163.367
R866 B.n207 B.n206 163.367
R867 B.n211 B.n210 163.367
R868 B.n215 B.n214 163.367
R869 B.n219 B.n218 163.367
R870 B.n223 B.n222 163.367
R871 B.n227 B.n226 163.367
R872 B.n231 B.n230 163.367
R873 B.n235 B.n234 163.367
R874 B.n239 B.n238 163.367
R875 B.n243 B.n242 163.367
R876 B.n247 B.n246 163.367
R877 B.n251 B.n250 163.367
R878 B.n255 B.n254 163.367
R879 B.n259 B.n258 163.367
R880 B.n263 B.n262 163.367
R881 B.n267 B.n266 163.367
R882 B.n271 B.n270 163.367
R883 B.n275 B.n274 163.367
R884 B.n279 B.n278 163.367
R885 B.n283 B.n282 163.367
R886 B.n287 B.n286 163.367
R887 B.n289 B.n124 163.367
R888 B.n588 B.n378 82.17
R889 B.n786 B.n785 82.17
R890 B.n587 B.n586 71.676
R891 B.n581 B.n382 71.676
R892 B.n578 B.n383 71.676
R893 B.n574 B.n384 71.676
R894 B.n570 B.n385 71.676
R895 B.n566 B.n386 71.676
R896 B.n562 B.n387 71.676
R897 B.n558 B.n388 71.676
R898 B.n554 B.n389 71.676
R899 B.n550 B.n390 71.676
R900 B.n546 B.n391 71.676
R901 B.n542 B.n392 71.676
R902 B.n538 B.n393 71.676
R903 B.n534 B.n394 71.676
R904 B.n530 B.n395 71.676
R905 B.n526 B.n396 71.676
R906 B.n522 B.n397 71.676
R907 B.n518 B.n398 71.676
R908 B.n513 B.n399 71.676
R909 B.n509 B.n400 71.676
R910 B.n505 B.n401 71.676
R911 B.n501 B.n402 71.676
R912 B.n497 B.n403 71.676
R913 B.n492 B.n404 71.676
R914 B.n488 B.n405 71.676
R915 B.n484 B.n406 71.676
R916 B.n480 B.n407 71.676
R917 B.n476 B.n408 71.676
R918 B.n472 B.n409 71.676
R919 B.n468 B.n410 71.676
R920 B.n464 B.n411 71.676
R921 B.n460 B.n412 71.676
R922 B.n456 B.n413 71.676
R923 B.n452 B.n414 71.676
R924 B.n448 B.n415 71.676
R925 B.n444 B.n416 71.676
R926 B.n440 B.n417 71.676
R927 B.n436 B.n418 71.676
R928 B.n432 B.n419 71.676
R929 B.n428 B.n420 71.676
R930 B.n131 B.n84 71.676
R931 B.n135 B.n85 71.676
R932 B.n139 B.n86 71.676
R933 B.n143 B.n87 71.676
R934 B.n147 B.n88 71.676
R935 B.n151 B.n89 71.676
R936 B.n155 B.n90 71.676
R937 B.n159 B.n91 71.676
R938 B.n163 B.n92 71.676
R939 B.n167 B.n93 71.676
R940 B.n171 B.n94 71.676
R941 B.n175 B.n95 71.676
R942 B.n179 B.n96 71.676
R943 B.n183 B.n97 71.676
R944 B.n187 B.n98 71.676
R945 B.n191 B.n99 71.676
R946 B.n195 B.n100 71.676
R947 B.n199 B.n101 71.676
R948 B.n203 B.n102 71.676
R949 B.n207 B.n103 71.676
R950 B.n211 B.n104 71.676
R951 B.n215 B.n105 71.676
R952 B.n219 B.n106 71.676
R953 B.n223 B.n107 71.676
R954 B.n227 B.n108 71.676
R955 B.n231 B.n109 71.676
R956 B.n235 B.n110 71.676
R957 B.n239 B.n111 71.676
R958 B.n243 B.n112 71.676
R959 B.n247 B.n113 71.676
R960 B.n251 B.n114 71.676
R961 B.n255 B.n115 71.676
R962 B.n259 B.n116 71.676
R963 B.n263 B.n117 71.676
R964 B.n267 B.n118 71.676
R965 B.n271 B.n119 71.676
R966 B.n275 B.n120 71.676
R967 B.n279 B.n121 71.676
R968 B.n283 B.n122 71.676
R969 B.n287 B.n123 71.676
R970 B.n784 B.n124 71.676
R971 B.n784 B.n783 71.676
R972 B.n289 B.n123 71.676
R973 B.n286 B.n122 71.676
R974 B.n282 B.n121 71.676
R975 B.n278 B.n120 71.676
R976 B.n274 B.n119 71.676
R977 B.n270 B.n118 71.676
R978 B.n266 B.n117 71.676
R979 B.n262 B.n116 71.676
R980 B.n258 B.n115 71.676
R981 B.n254 B.n114 71.676
R982 B.n250 B.n113 71.676
R983 B.n246 B.n112 71.676
R984 B.n242 B.n111 71.676
R985 B.n238 B.n110 71.676
R986 B.n234 B.n109 71.676
R987 B.n230 B.n108 71.676
R988 B.n226 B.n107 71.676
R989 B.n222 B.n106 71.676
R990 B.n218 B.n105 71.676
R991 B.n214 B.n104 71.676
R992 B.n210 B.n103 71.676
R993 B.n206 B.n102 71.676
R994 B.n202 B.n101 71.676
R995 B.n198 B.n100 71.676
R996 B.n194 B.n99 71.676
R997 B.n190 B.n98 71.676
R998 B.n186 B.n97 71.676
R999 B.n182 B.n96 71.676
R1000 B.n178 B.n95 71.676
R1001 B.n174 B.n94 71.676
R1002 B.n170 B.n93 71.676
R1003 B.n166 B.n92 71.676
R1004 B.n162 B.n91 71.676
R1005 B.n158 B.n90 71.676
R1006 B.n154 B.n89 71.676
R1007 B.n150 B.n88 71.676
R1008 B.n146 B.n87 71.676
R1009 B.n142 B.n86 71.676
R1010 B.n138 B.n85 71.676
R1011 B.n134 B.n84 71.676
R1012 B.n587 B.n422 71.676
R1013 B.n579 B.n382 71.676
R1014 B.n575 B.n383 71.676
R1015 B.n571 B.n384 71.676
R1016 B.n567 B.n385 71.676
R1017 B.n563 B.n386 71.676
R1018 B.n559 B.n387 71.676
R1019 B.n555 B.n388 71.676
R1020 B.n551 B.n389 71.676
R1021 B.n547 B.n390 71.676
R1022 B.n543 B.n391 71.676
R1023 B.n539 B.n392 71.676
R1024 B.n535 B.n393 71.676
R1025 B.n531 B.n394 71.676
R1026 B.n527 B.n395 71.676
R1027 B.n523 B.n396 71.676
R1028 B.n519 B.n397 71.676
R1029 B.n514 B.n398 71.676
R1030 B.n510 B.n399 71.676
R1031 B.n506 B.n400 71.676
R1032 B.n502 B.n401 71.676
R1033 B.n498 B.n402 71.676
R1034 B.n493 B.n403 71.676
R1035 B.n489 B.n404 71.676
R1036 B.n485 B.n405 71.676
R1037 B.n481 B.n406 71.676
R1038 B.n477 B.n407 71.676
R1039 B.n473 B.n408 71.676
R1040 B.n469 B.n409 71.676
R1041 B.n465 B.n410 71.676
R1042 B.n461 B.n411 71.676
R1043 B.n457 B.n412 71.676
R1044 B.n453 B.n413 71.676
R1045 B.n449 B.n414 71.676
R1046 B.n445 B.n415 71.676
R1047 B.n441 B.n416 71.676
R1048 B.n437 B.n417 71.676
R1049 B.n433 B.n418 71.676
R1050 B.n429 B.n419 71.676
R1051 B.n420 B.n381 71.676
R1052 B.n495 B.n426 59.5399
R1053 B.n516 B.n424 59.5399
R1054 B.n130 B.n129 59.5399
R1055 B.n127 B.n126 59.5399
R1056 B.n594 B.n378 48.5877
R1057 B.n594 B.n374 48.5877
R1058 B.n600 B.n374 48.5877
R1059 B.n600 B.n370 48.5877
R1060 B.n606 B.n370 48.5877
R1061 B.n606 B.n366 48.5877
R1062 B.n612 B.n366 48.5877
R1063 B.n618 B.n362 48.5877
R1064 B.n618 B.n358 48.5877
R1065 B.n624 B.n358 48.5877
R1066 B.n624 B.n354 48.5877
R1067 B.n630 B.n354 48.5877
R1068 B.n630 B.n350 48.5877
R1069 B.n636 B.n350 48.5877
R1070 B.n636 B.n346 48.5877
R1071 B.n642 B.n346 48.5877
R1072 B.n648 B.n342 48.5877
R1073 B.n648 B.n338 48.5877
R1074 B.n654 B.n338 48.5877
R1075 B.n654 B.n334 48.5877
R1076 B.n660 B.n334 48.5877
R1077 B.n660 B.n330 48.5877
R1078 B.n666 B.n330 48.5877
R1079 B.n672 B.n326 48.5877
R1080 B.n672 B.n322 48.5877
R1081 B.n678 B.n322 48.5877
R1082 B.n678 B.n317 48.5877
R1083 B.n684 B.n317 48.5877
R1084 B.n684 B.n318 48.5877
R1085 B.n690 B.n310 48.5877
R1086 B.n696 B.n310 48.5877
R1087 B.n696 B.n306 48.5877
R1088 B.n702 B.n306 48.5877
R1089 B.n702 B.n302 48.5877
R1090 B.n708 B.n302 48.5877
R1091 B.n715 B.n298 48.5877
R1092 B.n715 B.n294 48.5877
R1093 B.n721 B.n294 48.5877
R1094 B.n721 B.n4 48.5877
R1095 B.n875 B.n4 48.5877
R1096 B.n875 B.n874 48.5877
R1097 B.n874 B.n873 48.5877
R1098 B.n873 B.n8 48.5877
R1099 B.n867 B.n8 48.5877
R1100 B.n867 B.n866 48.5877
R1101 B.n865 B.n15 48.5877
R1102 B.n859 B.n15 48.5877
R1103 B.n859 B.n858 48.5877
R1104 B.n858 B.n857 48.5877
R1105 B.n857 B.n22 48.5877
R1106 B.n851 B.n22 48.5877
R1107 B.n850 B.n849 48.5877
R1108 B.n849 B.n29 48.5877
R1109 B.n843 B.n29 48.5877
R1110 B.n843 B.n842 48.5877
R1111 B.n842 B.n841 48.5877
R1112 B.n841 B.n36 48.5877
R1113 B.n835 B.n834 48.5877
R1114 B.n834 B.n833 48.5877
R1115 B.n833 B.n43 48.5877
R1116 B.n827 B.n43 48.5877
R1117 B.n827 B.n826 48.5877
R1118 B.n826 B.n825 48.5877
R1119 B.n825 B.n50 48.5877
R1120 B.n819 B.n818 48.5877
R1121 B.n818 B.n817 48.5877
R1122 B.n817 B.n57 48.5877
R1123 B.n811 B.n57 48.5877
R1124 B.n811 B.n810 48.5877
R1125 B.n810 B.n809 48.5877
R1126 B.n809 B.n64 48.5877
R1127 B.n803 B.n64 48.5877
R1128 B.n803 B.n802 48.5877
R1129 B.n801 B.n71 48.5877
R1130 B.n795 B.n71 48.5877
R1131 B.n795 B.n794 48.5877
R1132 B.n794 B.n793 48.5877
R1133 B.n793 B.n78 48.5877
R1134 B.n787 B.n78 48.5877
R1135 B.n787 B.n786 48.5877
R1136 B.n426 B.n425 48.4853
R1137 B.n424 B.n423 48.4853
R1138 B.n129 B.n128 48.4853
R1139 B.n126 B.n125 48.4853
R1140 B.t6 B.n326 47.8732
R1141 B.t5 B.n36 47.8732
R1142 B.t13 B.n362 43.5861
R1143 B.n802 B.t9 43.5861
R1144 B.n708 B.t0 35.0119
R1145 B.t3 B.n865 35.0119
R1146 B.n642 B.t7 32.1538
R1147 B.n819 B.t4 32.1538
R1148 B.n690 B.t1 30.7248
R1149 B.n851 B.t2 30.7248
R1150 B.n132 B.n80 29.8151
R1151 B.n782 B.n781 29.8151
R1152 B.n591 B.n590 29.8151
R1153 B.n585 B.n376 29.8151
R1154 B B.n877 18.0485
R1155 B.n318 B.t1 17.8634
R1156 B.t2 B.n850 17.8634
R1157 B.t7 B.n342 16.4344
R1158 B.t4 B.n50 16.4344
R1159 B.t0 B.n298 13.5763
R1160 B.n866 B.t3 13.5763
R1161 B.n133 B.n132 10.6151
R1162 B.n136 B.n133 10.6151
R1163 B.n137 B.n136 10.6151
R1164 B.n140 B.n137 10.6151
R1165 B.n141 B.n140 10.6151
R1166 B.n144 B.n141 10.6151
R1167 B.n145 B.n144 10.6151
R1168 B.n148 B.n145 10.6151
R1169 B.n149 B.n148 10.6151
R1170 B.n152 B.n149 10.6151
R1171 B.n153 B.n152 10.6151
R1172 B.n156 B.n153 10.6151
R1173 B.n157 B.n156 10.6151
R1174 B.n160 B.n157 10.6151
R1175 B.n161 B.n160 10.6151
R1176 B.n164 B.n161 10.6151
R1177 B.n165 B.n164 10.6151
R1178 B.n168 B.n165 10.6151
R1179 B.n169 B.n168 10.6151
R1180 B.n172 B.n169 10.6151
R1181 B.n173 B.n172 10.6151
R1182 B.n176 B.n173 10.6151
R1183 B.n177 B.n176 10.6151
R1184 B.n180 B.n177 10.6151
R1185 B.n181 B.n180 10.6151
R1186 B.n184 B.n181 10.6151
R1187 B.n185 B.n184 10.6151
R1188 B.n188 B.n185 10.6151
R1189 B.n189 B.n188 10.6151
R1190 B.n192 B.n189 10.6151
R1191 B.n193 B.n192 10.6151
R1192 B.n196 B.n193 10.6151
R1193 B.n197 B.n196 10.6151
R1194 B.n200 B.n197 10.6151
R1195 B.n201 B.n200 10.6151
R1196 B.n205 B.n204 10.6151
R1197 B.n208 B.n205 10.6151
R1198 B.n209 B.n208 10.6151
R1199 B.n212 B.n209 10.6151
R1200 B.n213 B.n212 10.6151
R1201 B.n216 B.n213 10.6151
R1202 B.n217 B.n216 10.6151
R1203 B.n220 B.n217 10.6151
R1204 B.n221 B.n220 10.6151
R1205 B.n225 B.n224 10.6151
R1206 B.n228 B.n225 10.6151
R1207 B.n229 B.n228 10.6151
R1208 B.n232 B.n229 10.6151
R1209 B.n233 B.n232 10.6151
R1210 B.n236 B.n233 10.6151
R1211 B.n237 B.n236 10.6151
R1212 B.n240 B.n237 10.6151
R1213 B.n241 B.n240 10.6151
R1214 B.n244 B.n241 10.6151
R1215 B.n245 B.n244 10.6151
R1216 B.n248 B.n245 10.6151
R1217 B.n249 B.n248 10.6151
R1218 B.n252 B.n249 10.6151
R1219 B.n253 B.n252 10.6151
R1220 B.n256 B.n253 10.6151
R1221 B.n257 B.n256 10.6151
R1222 B.n260 B.n257 10.6151
R1223 B.n261 B.n260 10.6151
R1224 B.n264 B.n261 10.6151
R1225 B.n265 B.n264 10.6151
R1226 B.n268 B.n265 10.6151
R1227 B.n269 B.n268 10.6151
R1228 B.n272 B.n269 10.6151
R1229 B.n273 B.n272 10.6151
R1230 B.n276 B.n273 10.6151
R1231 B.n277 B.n276 10.6151
R1232 B.n280 B.n277 10.6151
R1233 B.n281 B.n280 10.6151
R1234 B.n284 B.n281 10.6151
R1235 B.n285 B.n284 10.6151
R1236 B.n288 B.n285 10.6151
R1237 B.n290 B.n288 10.6151
R1238 B.n291 B.n290 10.6151
R1239 B.n782 B.n291 10.6151
R1240 B.n592 B.n591 10.6151
R1241 B.n592 B.n372 10.6151
R1242 B.n602 B.n372 10.6151
R1243 B.n603 B.n602 10.6151
R1244 B.n604 B.n603 10.6151
R1245 B.n604 B.n364 10.6151
R1246 B.n614 B.n364 10.6151
R1247 B.n615 B.n614 10.6151
R1248 B.n616 B.n615 10.6151
R1249 B.n616 B.n356 10.6151
R1250 B.n626 B.n356 10.6151
R1251 B.n627 B.n626 10.6151
R1252 B.n628 B.n627 10.6151
R1253 B.n628 B.n348 10.6151
R1254 B.n638 B.n348 10.6151
R1255 B.n639 B.n638 10.6151
R1256 B.n640 B.n639 10.6151
R1257 B.n640 B.n340 10.6151
R1258 B.n650 B.n340 10.6151
R1259 B.n651 B.n650 10.6151
R1260 B.n652 B.n651 10.6151
R1261 B.n652 B.n332 10.6151
R1262 B.n662 B.n332 10.6151
R1263 B.n663 B.n662 10.6151
R1264 B.n664 B.n663 10.6151
R1265 B.n664 B.n324 10.6151
R1266 B.n674 B.n324 10.6151
R1267 B.n675 B.n674 10.6151
R1268 B.n676 B.n675 10.6151
R1269 B.n676 B.n315 10.6151
R1270 B.n686 B.n315 10.6151
R1271 B.n687 B.n686 10.6151
R1272 B.n688 B.n687 10.6151
R1273 B.n688 B.n308 10.6151
R1274 B.n698 B.n308 10.6151
R1275 B.n699 B.n698 10.6151
R1276 B.n700 B.n699 10.6151
R1277 B.n700 B.n300 10.6151
R1278 B.n710 B.n300 10.6151
R1279 B.n711 B.n710 10.6151
R1280 B.n713 B.n711 10.6151
R1281 B.n713 B.n712 10.6151
R1282 B.n712 B.n292 10.6151
R1283 B.n724 B.n292 10.6151
R1284 B.n725 B.n724 10.6151
R1285 B.n726 B.n725 10.6151
R1286 B.n727 B.n726 10.6151
R1287 B.n729 B.n727 10.6151
R1288 B.n730 B.n729 10.6151
R1289 B.n731 B.n730 10.6151
R1290 B.n732 B.n731 10.6151
R1291 B.n734 B.n732 10.6151
R1292 B.n735 B.n734 10.6151
R1293 B.n736 B.n735 10.6151
R1294 B.n737 B.n736 10.6151
R1295 B.n739 B.n737 10.6151
R1296 B.n740 B.n739 10.6151
R1297 B.n741 B.n740 10.6151
R1298 B.n742 B.n741 10.6151
R1299 B.n744 B.n742 10.6151
R1300 B.n745 B.n744 10.6151
R1301 B.n746 B.n745 10.6151
R1302 B.n747 B.n746 10.6151
R1303 B.n749 B.n747 10.6151
R1304 B.n750 B.n749 10.6151
R1305 B.n751 B.n750 10.6151
R1306 B.n752 B.n751 10.6151
R1307 B.n754 B.n752 10.6151
R1308 B.n755 B.n754 10.6151
R1309 B.n756 B.n755 10.6151
R1310 B.n757 B.n756 10.6151
R1311 B.n759 B.n757 10.6151
R1312 B.n760 B.n759 10.6151
R1313 B.n761 B.n760 10.6151
R1314 B.n762 B.n761 10.6151
R1315 B.n764 B.n762 10.6151
R1316 B.n765 B.n764 10.6151
R1317 B.n766 B.n765 10.6151
R1318 B.n767 B.n766 10.6151
R1319 B.n769 B.n767 10.6151
R1320 B.n770 B.n769 10.6151
R1321 B.n771 B.n770 10.6151
R1322 B.n772 B.n771 10.6151
R1323 B.n774 B.n772 10.6151
R1324 B.n775 B.n774 10.6151
R1325 B.n776 B.n775 10.6151
R1326 B.n777 B.n776 10.6151
R1327 B.n779 B.n777 10.6151
R1328 B.n780 B.n779 10.6151
R1329 B.n781 B.n780 10.6151
R1330 B.n585 B.n584 10.6151
R1331 B.n584 B.n583 10.6151
R1332 B.n583 B.n582 10.6151
R1333 B.n582 B.n580 10.6151
R1334 B.n580 B.n577 10.6151
R1335 B.n577 B.n576 10.6151
R1336 B.n576 B.n573 10.6151
R1337 B.n573 B.n572 10.6151
R1338 B.n572 B.n569 10.6151
R1339 B.n569 B.n568 10.6151
R1340 B.n568 B.n565 10.6151
R1341 B.n565 B.n564 10.6151
R1342 B.n564 B.n561 10.6151
R1343 B.n561 B.n560 10.6151
R1344 B.n560 B.n557 10.6151
R1345 B.n557 B.n556 10.6151
R1346 B.n556 B.n553 10.6151
R1347 B.n553 B.n552 10.6151
R1348 B.n552 B.n549 10.6151
R1349 B.n549 B.n548 10.6151
R1350 B.n548 B.n545 10.6151
R1351 B.n545 B.n544 10.6151
R1352 B.n544 B.n541 10.6151
R1353 B.n541 B.n540 10.6151
R1354 B.n540 B.n537 10.6151
R1355 B.n537 B.n536 10.6151
R1356 B.n536 B.n533 10.6151
R1357 B.n533 B.n532 10.6151
R1358 B.n532 B.n529 10.6151
R1359 B.n529 B.n528 10.6151
R1360 B.n528 B.n525 10.6151
R1361 B.n525 B.n524 10.6151
R1362 B.n524 B.n521 10.6151
R1363 B.n521 B.n520 10.6151
R1364 B.n520 B.n517 10.6151
R1365 B.n515 B.n512 10.6151
R1366 B.n512 B.n511 10.6151
R1367 B.n511 B.n508 10.6151
R1368 B.n508 B.n507 10.6151
R1369 B.n507 B.n504 10.6151
R1370 B.n504 B.n503 10.6151
R1371 B.n503 B.n500 10.6151
R1372 B.n500 B.n499 10.6151
R1373 B.n499 B.n496 10.6151
R1374 B.n494 B.n491 10.6151
R1375 B.n491 B.n490 10.6151
R1376 B.n490 B.n487 10.6151
R1377 B.n487 B.n486 10.6151
R1378 B.n486 B.n483 10.6151
R1379 B.n483 B.n482 10.6151
R1380 B.n482 B.n479 10.6151
R1381 B.n479 B.n478 10.6151
R1382 B.n478 B.n475 10.6151
R1383 B.n475 B.n474 10.6151
R1384 B.n474 B.n471 10.6151
R1385 B.n471 B.n470 10.6151
R1386 B.n470 B.n467 10.6151
R1387 B.n467 B.n466 10.6151
R1388 B.n466 B.n463 10.6151
R1389 B.n463 B.n462 10.6151
R1390 B.n462 B.n459 10.6151
R1391 B.n459 B.n458 10.6151
R1392 B.n458 B.n455 10.6151
R1393 B.n455 B.n454 10.6151
R1394 B.n454 B.n451 10.6151
R1395 B.n451 B.n450 10.6151
R1396 B.n450 B.n447 10.6151
R1397 B.n447 B.n446 10.6151
R1398 B.n446 B.n443 10.6151
R1399 B.n443 B.n442 10.6151
R1400 B.n442 B.n439 10.6151
R1401 B.n439 B.n438 10.6151
R1402 B.n438 B.n435 10.6151
R1403 B.n435 B.n434 10.6151
R1404 B.n434 B.n431 10.6151
R1405 B.n431 B.n430 10.6151
R1406 B.n430 B.n427 10.6151
R1407 B.n427 B.n380 10.6151
R1408 B.n590 B.n380 10.6151
R1409 B.n596 B.n376 10.6151
R1410 B.n597 B.n596 10.6151
R1411 B.n598 B.n597 10.6151
R1412 B.n598 B.n368 10.6151
R1413 B.n608 B.n368 10.6151
R1414 B.n609 B.n608 10.6151
R1415 B.n610 B.n609 10.6151
R1416 B.n610 B.n360 10.6151
R1417 B.n620 B.n360 10.6151
R1418 B.n621 B.n620 10.6151
R1419 B.n622 B.n621 10.6151
R1420 B.n622 B.n352 10.6151
R1421 B.n632 B.n352 10.6151
R1422 B.n633 B.n632 10.6151
R1423 B.n634 B.n633 10.6151
R1424 B.n634 B.n344 10.6151
R1425 B.n644 B.n344 10.6151
R1426 B.n645 B.n644 10.6151
R1427 B.n646 B.n645 10.6151
R1428 B.n646 B.n336 10.6151
R1429 B.n656 B.n336 10.6151
R1430 B.n657 B.n656 10.6151
R1431 B.n658 B.n657 10.6151
R1432 B.n658 B.n328 10.6151
R1433 B.n668 B.n328 10.6151
R1434 B.n669 B.n668 10.6151
R1435 B.n670 B.n669 10.6151
R1436 B.n670 B.n320 10.6151
R1437 B.n680 B.n320 10.6151
R1438 B.n681 B.n680 10.6151
R1439 B.n682 B.n681 10.6151
R1440 B.n682 B.n312 10.6151
R1441 B.n692 B.n312 10.6151
R1442 B.n693 B.n692 10.6151
R1443 B.n694 B.n693 10.6151
R1444 B.n694 B.n304 10.6151
R1445 B.n704 B.n304 10.6151
R1446 B.n705 B.n704 10.6151
R1447 B.n706 B.n705 10.6151
R1448 B.n706 B.n296 10.6151
R1449 B.n717 B.n296 10.6151
R1450 B.n718 B.n717 10.6151
R1451 B.n719 B.n718 10.6151
R1452 B.n719 B.n0 10.6151
R1453 B.n871 B.n1 10.6151
R1454 B.n871 B.n870 10.6151
R1455 B.n870 B.n869 10.6151
R1456 B.n869 B.n10 10.6151
R1457 B.n863 B.n10 10.6151
R1458 B.n863 B.n862 10.6151
R1459 B.n862 B.n861 10.6151
R1460 B.n861 B.n17 10.6151
R1461 B.n855 B.n17 10.6151
R1462 B.n855 B.n854 10.6151
R1463 B.n854 B.n853 10.6151
R1464 B.n853 B.n24 10.6151
R1465 B.n847 B.n24 10.6151
R1466 B.n847 B.n846 10.6151
R1467 B.n846 B.n845 10.6151
R1468 B.n845 B.n31 10.6151
R1469 B.n839 B.n31 10.6151
R1470 B.n839 B.n838 10.6151
R1471 B.n838 B.n837 10.6151
R1472 B.n837 B.n38 10.6151
R1473 B.n831 B.n38 10.6151
R1474 B.n831 B.n830 10.6151
R1475 B.n830 B.n829 10.6151
R1476 B.n829 B.n45 10.6151
R1477 B.n823 B.n45 10.6151
R1478 B.n823 B.n822 10.6151
R1479 B.n822 B.n821 10.6151
R1480 B.n821 B.n52 10.6151
R1481 B.n815 B.n52 10.6151
R1482 B.n815 B.n814 10.6151
R1483 B.n814 B.n813 10.6151
R1484 B.n813 B.n59 10.6151
R1485 B.n807 B.n59 10.6151
R1486 B.n807 B.n806 10.6151
R1487 B.n806 B.n805 10.6151
R1488 B.n805 B.n66 10.6151
R1489 B.n799 B.n66 10.6151
R1490 B.n799 B.n798 10.6151
R1491 B.n798 B.n797 10.6151
R1492 B.n797 B.n73 10.6151
R1493 B.n791 B.n73 10.6151
R1494 B.n791 B.n790 10.6151
R1495 B.n790 B.n789 10.6151
R1496 B.n789 B.n80 10.6151
R1497 B.n201 B.n130 9.36635
R1498 B.n224 B.n127 9.36635
R1499 B.n517 B.n516 9.36635
R1500 B.n495 B.n494 9.36635
R1501 B.n612 B.t13 5.00212
R1502 B.t9 B.n801 5.00212
R1503 B.n877 B.n0 2.81026
R1504 B.n877 B.n1 2.81026
R1505 B.n204 B.n130 1.24928
R1506 B.n221 B.n127 1.24928
R1507 B.n516 B.n515 1.24928
R1508 B.n496 B.n495 1.24928
R1509 B.n666 B.t6 0.715018
R1510 B.n835 B.t5 0.715018
R1511 VN.n47 VN.n25 161.3
R1512 VN.n46 VN.n45 161.3
R1513 VN.n44 VN.n26 161.3
R1514 VN.n43 VN.n42 161.3
R1515 VN.n41 VN.n27 161.3
R1516 VN.n39 VN.n38 161.3
R1517 VN.n37 VN.n28 161.3
R1518 VN.n36 VN.n35 161.3
R1519 VN.n34 VN.n29 161.3
R1520 VN.n33 VN.n32 161.3
R1521 VN.n22 VN.n0 161.3
R1522 VN.n21 VN.n20 161.3
R1523 VN.n19 VN.n1 161.3
R1524 VN.n18 VN.n17 161.3
R1525 VN.n16 VN.n2 161.3
R1526 VN.n14 VN.n13 161.3
R1527 VN.n12 VN.n3 161.3
R1528 VN.n11 VN.n10 161.3
R1529 VN.n9 VN.n4 161.3
R1530 VN.n8 VN.n7 161.3
R1531 VN.n6 VN.t6 144.47
R1532 VN.n31 VN.t4 144.47
R1533 VN.n5 VN.t3 112.394
R1534 VN.n15 VN.t7 112.394
R1535 VN.n23 VN.t2 112.394
R1536 VN.n30 VN.t0 112.394
R1537 VN.n40 VN.t5 112.394
R1538 VN.n48 VN.t1 112.394
R1539 VN.n24 VN.n23 98.6123
R1540 VN.n49 VN.n48 98.6123
R1541 VN.n6 VN.n5 59.4159
R1542 VN.n31 VN.n30 59.4159
R1543 VN VN.n49 47.6876
R1544 VN.n10 VN.n9 40.577
R1545 VN.n10 VN.n3 40.577
R1546 VN.n17 VN.n1 40.577
R1547 VN.n21 VN.n1 40.577
R1548 VN.n35 VN.n34 40.577
R1549 VN.n35 VN.n28 40.577
R1550 VN.n42 VN.n26 40.577
R1551 VN.n46 VN.n26 40.577
R1552 VN.n9 VN.n8 24.5923
R1553 VN.n14 VN.n3 24.5923
R1554 VN.n17 VN.n16 24.5923
R1555 VN.n22 VN.n21 24.5923
R1556 VN.n34 VN.n33 24.5923
R1557 VN.n42 VN.n41 24.5923
R1558 VN.n39 VN.n28 24.5923
R1559 VN.n47 VN.n46 24.5923
R1560 VN.n8 VN.n5 12.2964
R1561 VN.n15 VN.n14 12.2964
R1562 VN.n16 VN.n15 12.2964
R1563 VN.n23 VN.n22 12.2964
R1564 VN.n33 VN.n30 12.2964
R1565 VN.n41 VN.n40 12.2964
R1566 VN.n40 VN.n39 12.2964
R1567 VN.n48 VN.n47 12.2964
R1568 VN.n32 VN.n31 9.706
R1569 VN.n7 VN.n6 9.706
R1570 VN.n49 VN.n25 0.278335
R1571 VN.n24 VN.n0 0.278335
R1572 VN.n45 VN.n25 0.189894
R1573 VN.n45 VN.n44 0.189894
R1574 VN.n44 VN.n43 0.189894
R1575 VN.n43 VN.n27 0.189894
R1576 VN.n38 VN.n27 0.189894
R1577 VN.n38 VN.n37 0.189894
R1578 VN.n37 VN.n36 0.189894
R1579 VN.n36 VN.n29 0.189894
R1580 VN.n32 VN.n29 0.189894
R1581 VN.n7 VN.n4 0.189894
R1582 VN.n11 VN.n4 0.189894
R1583 VN.n12 VN.n11 0.189894
R1584 VN.n13 VN.n12 0.189894
R1585 VN.n13 VN.n2 0.189894
R1586 VN.n18 VN.n2 0.189894
R1587 VN.n19 VN.n18 0.189894
R1588 VN.n20 VN.n19 0.189894
R1589 VN.n20 VN.n0 0.189894
R1590 VN VN.n24 0.153485
R1591 VDD2.n2 VDD2.n1 66.7654
R1592 VDD2.n2 VDD2.n0 66.7654
R1593 VDD2 VDD2.n5 66.7626
R1594 VDD2.n4 VDD2.n3 65.7434
R1595 VDD2.n4 VDD2.n2 42.1377
R1596 VDD2.n5 VDD2.t3 1.95702
R1597 VDD2.n5 VDD2.t6 1.95702
R1598 VDD2.n3 VDD2.t4 1.95702
R1599 VDD2.n3 VDD2.t2 1.95702
R1600 VDD2.n1 VDD2.t7 1.95702
R1601 VDD2.n1 VDD2.t0 1.95702
R1602 VDD2.n0 VDD2.t1 1.95702
R1603 VDD2.n0 VDD2.t5 1.95702
R1604 VDD2 VDD2.n4 1.13628
R1605 VTAIL.n434 VTAIL.n386 289.615
R1606 VTAIL.n50 VTAIL.n2 289.615
R1607 VTAIL.n104 VTAIL.n56 289.615
R1608 VTAIL.n160 VTAIL.n112 289.615
R1609 VTAIL.n380 VTAIL.n332 289.615
R1610 VTAIL.n324 VTAIL.n276 289.615
R1611 VTAIL.n270 VTAIL.n222 289.615
R1612 VTAIL.n214 VTAIL.n166 289.615
R1613 VTAIL.n402 VTAIL.n401 185
R1614 VTAIL.n407 VTAIL.n406 185
R1615 VTAIL.n409 VTAIL.n408 185
R1616 VTAIL.n398 VTAIL.n397 185
R1617 VTAIL.n415 VTAIL.n414 185
R1618 VTAIL.n417 VTAIL.n416 185
R1619 VTAIL.n394 VTAIL.n393 185
R1620 VTAIL.n424 VTAIL.n423 185
R1621 VTAIL.n425 VTAIL.n392 185
R1622 VTAIL.n427 VTAIL.n426 185
R1623 VTAIL.n390 VTAIL.n389 185
R1624 VTAIL.n433 VTAIL.n432 185
R1625 VTAIL.n435 VTAIL.n434 185
R1626 VTAIL.n18 VTAIL.n17 185
R1627 VTAIL.n23 VTAIL.n22 185
R1628 VTAIL.n25 VTAIL.n24 185
R1629 VTAIL.n14 VTAIL.n13 185
R1630 VTAIL.n31 VTAIL.n30 185
R1631 VTAIL.n33 VTAIL.n32 185
R1632 VTAIL.n10 VTAIL.n9 185
R1633 VTAIL.n40 VTAIL.n39 185
R1634 VTAIL.n41 VTAIL.n8 185
R1635 VTAIL.n43 VTAIL.n42 185
R1636 VTAIL.n6 VTAIL.n5 185
R1637 VTAIL.n49 VTAIL.n48 185
R1638 VTAIL.n51 VTAIL.n50 185
R1639 VTAIL.n72 VTAIL.n71 185
R1640 VTAIL.n77 VTAIL.n76 185
R1641 VTAIL.n79 VTAIL.n78 185
R1642 VTAIL.n68 VTAIL.n67 185
R1643 VTAIL.n85 VTAIL.n84 185
R1644 VTAIL.n87 VTAIL.n86 185
R1645 VTAIL.n64 VTAIL.n63 185
R1646 VTAIL.n94 VTAIL.n93 185
R1647 VTAIL.n95 VTAIL.n62 185
R1648 VTAIL.n97 VTAIL.n96 185
R1649 VTAIL.n60 VTAIL.n59 185
R1650 VTAIL.n103 VTAIL.n102 185
R1651 VTAIL.n105 VTAIL.n104 185
R1652 VTAIL.n128 VTAIL.n127 185
R1653 VTAIL.n133 VTAIL.n132 185
R1654 VTAIL.n135 VTAIL.n134 185
R1655 VTAIL.n124 VTAIL.n123 185
R1656 VTAIL.n141 VTAIL.n140 185
R1657 VTAIL.n143 VTAIL.n142 185
R1658 VTAIL.n120 VTAIL.n119 185
R1659 VTAIL.n150 VTAIL.n149 185
R1660 VTAIL.n151 VTAIL.n118 185
R1661 VTAIL.n153 VTAIL.n152 185
R1662 VTAIL.n116 VTAIL.n115 185
R1663 VTAIL.n159 VTAIL.n158 185
R1664 VTAIL.n161 VTAIL.n160 185
R1665 VTAIL.n381 VTAIL.n380 185
R1666 VTAIL.n379 VTAIL.n378 185
R1667 VTAIL.n336 VTAIL.n335 185
R1668 VTAIL.n373 VTAIL.n372 185
R1669 VTAIL.n371 VTAIL.n338 185
R1670 VTAIL.n370 VTAIL.n369 185
R1671 VTAIL.n341 VTAIL.n339 185
R1672 VTAIL.n364 VTAIL.n363 185
R1673 VTAIL.n362 VTAIL.n361 185
R1674 VTAIL.n345 VTAIL.n344 185
R1675 VTAIL.n356 VTAIL.n355 185
R1676 VTAIL.n354 VTAIL.n353 185
R1677 VTAIL.n349 VTAIL.n348 185
R1678 VTAIL.n325 VTAIL.n324 185
R1679 VTAIL.n323 VTAIL.n322 185
R1680 VTAIL.n280 VTAIL.n279 185
R1681 VTAIL.n317 VTAIL.n316 185
R1682 VTAIL.n315 VTAIL.n282 185
R1683 VTAIL.n314 VTAIL.n313 185
R1684 VTAIL.n285 VTAIL.n283 185
R1685 VTAIL.n308 VTAIL.n307 185
R1686 VTAIL.n306 VTAIL.n305 185
R1687 VTAIL.n289 VTAIL.n288 185
R1688 VTAIL.n300 VTAIL.n299 185
R1689 VTAIL.n298 VTAIL.n297 185
R1690 VTAIL.n293 VTAIL.n292 185
R1691 VTAIL.n271 VTAIL.n270 185
R1692 VTAIL.n269 VTAIL.n268 185
R1693 VTAIL.n226 VTAIL.n225 185
R1694 VTAIL.n263 VTAIL.n262 185
R1695 VTAIL.n261 VTAIL.n228 185
R1696 VTAIL.n260 VTAIL.n259 185
R1697 VTAIL.n231 VTAIL.n229 185
R1698 VTAIL.n254 VTAIL.n253 185
R1699 VTAIL.n252 VTAIL.n251 185
R1700 VTAIL.n235 VTAIL.n234 185
R1701 VTAIL.n246 VTAIL.n245 185
R1702 VTAIL.n244 VTAIL.n243 185
R1703 VTAIL.n239 VTAIL.n238 185
R1704 VTAIL.n215 VTAIL.n214 185
R1705 VTAIL.n213 VTAIL.n212 185
R1706 VTAIL.n170 VTAIL.n169 185
R1707 VTAIL.n207 VTAIL.n206 185
R1708 VTAIL.n205 VTAIL.n172 185
R1709 VTAIL.n204 VTAIL.n203 185
R1710 VTAIL.n175 VTAIL.n173 185
R1711 VTAIL.n198 VTAIL.n197 185
R1712 VTAIL.n196 VTAIL.n195 185
R1713 VTAIL.n179 VTAIL.n178 185
R1714 VTAIL.n190 VTAIL.n189 185
R1715 VTAIL.n188 VTAIL.n187 185
R1716 VTAIL.n183 VTAIL.n182 185
R1717 VTAIL.n403 VTAIL.t13 149.524
R1718 VTAIL.n19 VTAIL.t9 149.524
R1719 VTAIL.n73 VTAIL.t0 149.524
R1720 VTAIL.n129 VTAIL.t6 149.524
R1721 VTAIL.n350 VTAIL.t3 149.524
R1722 VTAIL.n294 VTAIL.t7 149.524
R1723 VTAIL.n240 VTAIL.t11 149.524
R1724 VTAIL.n184 VTAIL.t14 149.524
R1725 VTAIL.n407 VTAIL.n401 104.615
R1726 VTAIL.n408 VTAIL.n407 104.615
R1727 VTAIL.n408 VTAIL.n397 104.615
R1728 VTAIL.n415 VTAIL.n397 104.615
R1729 VTAIL.n416 VTAIL.n415 104.615
R1730 VTAIL.n416 VTAIL.n393 104.615
R1731 VTAIL.n424 VTAIL.n393 104.615
R1732 VTAIL.n425 VTAIL.n424 104.615
R1733 VTAIL.n426 VTAIL.n425 104.615
R1734 VTAIL.n426 VTAIL.n389 104.615
R1735 VTAIL.n433 VTAIL.n389 104.615
R1736 VTAIL.n434 VTAIL.n433 104.615
R1737 VTAIL.n23 VTAIL.n17 104.615
R1738 VTAIL.n24 VTAIL.n23 104.615
R1739 VTAIL.n24 VTAIL.n13 104.615
R1740 VTAIL.n31 VTAIL.n13 104.615
R1741 VTAIL.n32 VTAIL.n31 104.615
R1742 VTAIL.n32 VTAIL.n9 104.615
R1743 VTAIL.n40 VTAIL.n9 104.615
R1744 VTAIL.n41 VTAIL.n40 104.615
R1745 VTAIL.n42 VTAIL.n41 104.615
R1746 VTAIL.n42 VTAIL.n5 104.615
R1747 VTAIL.n49 VTAIL.n5 104.615
R1748 VTAIL.n50 VTAIL.n49 104.615
R1749 VTAIL.n77 VTAIL.n71 104.615
R1750 VTAIL.n78 VTAIL.n77 104.615
R1751 VTAIL.n78 VTAIL.n67 104.615
R1752 VTAIL.n85 VTAIL.n67 104.615
R1753 VTAIL.n86 VTAIL.n85 104.615
R1754 VTAIL.n86 VTAIL.n63 104.615
R1755 VTAIL.n94 VTAIL.n63 104.615
R1756 VTAIL.n95 VTAIL.n94 104.615
R1757 VTAIL.n96 VTAIL.n95 104.615
R1758 VTAIL.n96 VTAIL.n59 104.615
R1759 VTAIL.n103 VTAIL.n59 104.615
R1760 VTAIL.n104 VTAIL.n103 104.615
R1761 VTAIL.n133 VTAIL.n127 104.615
R1762 VTAIL.n134 VTAIL.n133 104.615
R1763 VTAIL.n134 VTAIL.n123 104.615
R1764 VTAIL.n141 VTAIL.n123 104.615
R1765 VTAIL.n142 VTAIL.n141 104.615
R1766 VTAIL.n142 VTAIL.n119 104.615
R1767 VTAIL.n150 VTAIL.n119 104.615
R1768 VTAIL.n151 VTAIL.n150 104.615
R1769 VTAIL.n152 VTAIL.n151 104.615
R1770 VTAIL.n152 VTAIL.n115 104.615
R1771 VTAIL.n159 VTAIL.n115 104.615
R1772 VTAIL.n160 VTAIL.n159 104.615
R1773 VTAIL.n380 VTAIL.n379 104.615
R1774 VTAIL.n379 VTAIL.n335 104.615
R1775 VTAIL.n372 VTAIL.n335 104.615
R1776 VTAIL.n372 VTAIL.n371 104.615
R1777 VTAIL.n371 VTAIL.n370 104.615
R1778 VTAIL.n370 VTAIL.n339 104.615
R1779 VTAIL.n363 VTAIL.n339 104.615
R1780 VTAIL.n363 VTAIL.n362 104.615
R1781 VTAIL.n362 VTAIL.n344 104.615
R1782 VTAIL.n355 VTAIL.n344 104.615
R1783 VTAIL.n355 VTAIL.n354 104.615
R1784 VTAIL.n354 VTAIL.n348 104.615
R1785 VTAIL.n324 VTAIL.n323 104.615
R1786 VTAIL.n323 VTAIL.n279 104.615
R1787 VTAIL.n316 VTAIL.n279 104.615
R1788 VTAIL.n316 VTAIL.n315 104.615
R1789 VTAIL.n315 VTAIL.n314 104.615
R1790 VTAIL.n314 VTAIL.n283 104.615
R1791 VTAIL.n307 VTAIL.n283 104.615
R1792 VTAIL.n307 VTAIL.n306 104.615
R1793 VTAIL.n306 VTAIL.n288 104.615
R1794 VTAIL.n299 VTAIL.n288 104.615
R1795 VTAIL.n299 VTAIL.n298 104.615
R1796 VTAIL.n298 VTAIL.n292 104.615
R1797 VTAIL.n270 VTAIL.n269 104.615
R1798 VTAIL.n269 VTAIL.n225 104.615
R1799 VTAIL.n262 VTAIL.n225 104.615
R1800 VTAIL.n262 VTAIL.n261 104.615
R1801 VTAIL.n261 VTAIL.n260 104.615
R1802 VTAIL.n260 VTAIL.n229 104.615
R1803 VTAIL.n253 VTAIL.n229 104.615
R1804 VTAIL.n253 VTAIL.n252 104.615
R1805 VTAIL.n252 VTAIL.n234 104.615
R1806 VTAIL.n245 VTAIL.n234 104.615
R1807 VTAIL.n245 VTAIL.n244 104.615
R1808 VTAIL.n244 VTAIL.n238 104.615
R1809 VTAIL.n214 VTAIL.n213 104.615
R1810 VTAIL.n213 VTAIL.n169 104.615
R1811 VTAIL.n206 VTAIL.n169 104.615
R1812 VTAIL.n206 VTAIL.n205 104.615
R1813 VTAIL.n205 VTAIL.n204 104.615
R1814 VTAIL.n204 VTAIL.n173 104.615
R1815 VTAIL.n197 VTAIL.n173 104.615
R1816 VTAIL.n197 VTAIL.n196 104.615
R1817 VTAIL.n196 VTAIL.n178 104.615
R1818 VTAIL.n189 VTAIL.n178 104.615
R1819 VTAIL.n189 VTAIL.n188 104.615
R1820 VTAIL.n188 VTAIL.n182 104.615
R1821 VTAIL.t13 VTAIL.n401 52.3082
R1822 VTAIL.t9 VTAIL.n17 52.3082
R1823 VTAIL.t0 VTAIL.n71 52.3082
R1824 VTAIL.t6 VTAIL.n127 52.3082
R1825 VTAIL.t3 VTAIL.n348 52.3082
R1826 VTAIL.t7 VTAIL.n292 52.3082
R1827 VTAIL.t11 VTAIL.n238 52.3082
R1828 VTAIL.t14 VTAIL.n182 52.3082
R1829 VTAIL.n331 VTAIL.n330 49.0646
R1830 VTAIL.n221 VTAIL.n220 49.0646
R1831 VTAIL.n1 VTAIL.n0 49.0644
R1832 VTAIL.n111 VTAIL.n110 49.0644
R1833 VTAIL.n439 VTAIL.n438 35.2884
R1834 VTAIL.n55 VTAIL.n54 35.2884
R1835 VTAIL.n109 VTAIL.n108 35.2884
R1836 VTAIL.n165 VTAIL.n164 35.2884
R1837 VTAIL.n385 VTAIL.n384 35.2884
R1838 VTAIL.n329 VTAIL.n328 35.2884
R1839 VTAIL.n275 VTAIL.n274 35.2884
R1840 VTAIL.n219 VTAIL.n218 35.2884
R1841 VTAIL.n439 VTAIL.n385 23.2462
R1842 VTAIL.n219 VTAIL.n165 23.2462
R1843 VTAIL.n427 VTAIL.n392 13.1884
R1844 VTAIL.n43 VTAIL.n8 13.1884
R1845 VTAIL.n97 VTAIL.n62 13.1884
R1846 VTAIL.n153 VTAIL.n118 13.1884
R1847 VTAIL.n373 VTAIL.n338 13.1884
R1848 VTAIL.n317 VTAIL.n282 13.1884
R1849 VTAIL.n263 VTAIL.n228 13.1884
R1850 VTAIL.n207 VTAIL.n172 13.1884
R1851 VTAIL.n423 VTAIL.n422 12.8005
R1852 VTAIL.n428 VTAIL.n390 12.8005
R1853 VTAIL.n39 VTAIL.n38 12.8005
R1854 VTAIL.n44 VTAIL.n6 12.8005
R1855 VTAIL.n93 VTAIL.n92 12.8005
R1856 VTAIL.n98 VTAIL.n60 12.8005
R1857 VTAIL.n149 VTAIL.n148 12.8005
R1858 VTAIL.n154 VTAIL.n116 12.8005
R1859 VTAIL.n374 VTAIL.n336 12.8005
R1860 VTAIL.n369 VTAIL.n340 12.8005
R1861 VTAIL.n318 VTAIL.n280 12.8005
R1862 VTAIL.n313 VTAIL.n284 12.8005
R1863 VTAIL.n264 VTAIL.n226 12.8005
R1864 VTAIL.n259 VTAIL.n230 12.8005
R1865 VTAIL.n208 VTAIL.n170 12.8005
R1866 VTAIL.n203 VTAIL.n174 12.8005
R1867 VTAIL.n421 VTAIL.n394 12.0247
R1868 VTAIL.n432 VTAIL.n431 12.0247
R1869 VTAIL.n37 VTAIL.n10 12.0247
R1870 VTAIL.n48 VTAIL.n47 12.0247
R1871 VTAIL.n91 VTAIL.n64 12.0247
R1872 VTAIL.n102 VTAIL.n101 12.0247
R1873 VTAIL.n147 VTAIL.n120 12.0247
R1874 VTAIL.n158 VTAIL.n157 12.0247
R1875 VTAIL.n378 VTAIL.n377 12.0247
R1876 VTAIL.n368 VTAIL.n341 12.0247
R1877 VTAIL.n322 VTAIL.n321 12.0247
R1878 VTAIL.n312 VTAIL.n285 12.0247
R1879 VTAIL.n268 VTAIL.n267 12.0247
R1880 VTAIL.n258 VTAIL.n231 12.0247
R1881 VTAIL.n212 VTAIL.n211 12.0247
R1882 VTAIL.n202 VTAIL.n175 12.0247
R1883 VTAIL.n418 VTAIL.n417 11.249
R1884 VTAIL.n435 VTAIL.n388 11.249
R1885 VTAIL.n34 VTAIL.n33 11.249
R1886 VTAIL.n51 VTAIL.n4 11.249
R1887 VTAIL.n88 VTAIL.n87 11.249
R1888 VTAIL.n105 VTAIL.n58 11.249
R1889 VTAIL.n144 VTAIL.n143 11.249
R1890 VTAIL.n161 VTAIL.n114 11.249
R1891 VTAIL.n381 VTAIL.n334 11.249
R1892 VTAIL.n365 VTAIL.n364 11.249
R1893 VTAIL.n325 VTAIL.n278 11.249
R1894 VTAIL.n309 VTAIL.n308 11.249
R1895 VTAIL.n271 VTAIL.n224 11.249
R1896 VTAIL.n255 VTAIL.n254 11.249
R1897 VTAIL.n215 VTAIL.n168 11.249
R1898 VTAIL.n199 VTAIL.n198 11.249
R1899 VTAIL.n414 VTAIL.n396 10.4732
R1900 VTAIL.n436 VTAIL.n386 10.4732
R1901 VTAIL.n30 VTAIL.n12 10.4732
R1902 VTAIL.n52 VTAIL.n2 10.4732
R1903 VTAIL.n84 VTAIL.n66 10.4732
R1904 VTAIL.n106 VTAIL.n56 10.4732
R1905 VTAIL.n140 VTAIL.n122 10.4732
R1906 VTAIL.n162 VTAIL.n112 10.4732
R1907 VTAIL.n382 VTAIL.n332 10.4732
R1908 VTAIL.n361 VTAIL.n343 10.4732
R1909 VTAIL.n326 VTAIL.n276 10.4732
R1910 VTAIL.n305 VTAIL.n287 10.4732
R1911 VTAIL.n272 VTAIL.n222 10.4732
R1912 VTAIL.n251 VTAIL.n233 10.4732
R1913 VTAIL.n216 VTAIL.n166 10.4732
R1914 VTAIL.n195 VTAIL.n177 10.4732
R1915 VTAIL.n403 VTAIL.n402 10.2747
R1916 VTAIL.n19 VTAIL.n18 10.2747
R1917 VTAIL.n73 VTAIL.n72 10.2747
R1918 VTAIL.n129 VTAIL.n128 10.2747
R1919 VTAIL.n350 VTAIL.n349 10.2747
R1920 VTAIL.n294 VTAIL.n293 10.2747
R1921 VTAIL.n240 VTAIL.n239 10.2747
R1922 VTAIL.n184 VTAIL.n183 10.2747
R1923 VTAIL.n413 VTAIL.n398 9.69747
R1924 VTAIL.n29 VTAIL.n14 9.69747
R1925 VTAIL.n83 VTAIL.n68 9.69747
R1926 VTAIL.n139 VTAIL.n124 9.69747
R1927 VTAIL.n360 VTAIL.n345 9.69747
R1928 VTAIL.n304 VTAIL.n289 9.69747
R1929 VTAIL.n250 VTAIL.n235 9.69747
R1930 VTAIL.n194 VTAIL.n179 9.69747
R1931 VTAIL.n438 VTAIL.n437 9.45567
R1932 VTAIL.n54 VTAIL.n53 9.45567
R1933 VTAIL.n108 VTAIL.n107 9.45567
R1934 VTAIL.n164 VTAIL.n163 9.45567
R1935 VTAIL.n384 VTAIL.n383 9.45567
R1936 VTAIL.n328 VTAIL.n327 9.45567
R1937 VTAIL.n274 VTAIL.n273 9.45567
R1938 VTAIL.n218 VTAIL.n217 9.45567
R1939 VTAIL.n437 VTAIL.n436 9.3005
R1940 VTAIL.n388 VTAIL.n387 9.3005
R1941 VTAIL.n431 VTAIL.n430 9.3005
R1942 VTAIL.n429 VTAIL.n428 9.3005
R1943 VTAIL.n405 VTAIL.n404 9.3005
R1944 VTAIL.n400 VTAIL.n399 9.3005
R1945 VTAIL.n411 VTAIL.n410 9.3005
R1946 VTAIL.n413 VTAIL.n412 9.3005
R1947 VTAIL.n396 VTAIL.n395 9.3005
R1948 VTAIL.n419 VTAIL.n418 9.3005
R1949 VTAIL.n421 VTAIL.n420 9.3005
R1950 VTAIL.n422 VTAIL.n391 9.3005
R1951 VTAIL.n53 VTAIL.n52 9.3005
R1952 VTAIL.n4 VTAIL.n3 9.3005
R1953 VTAIL.n47 VTAIL.n46 9.3005
R1954 VTAIL.n45 VTAIL.n44 9.3005
R1955 VTAIL.n21 VTAIL.n20 9.3005
R1956 VTAIL.n16 VTAIL.n15 9.3005
R1957 VTAIL.n27 VTAIL.n26 9.3005
R1958 VTAIL.n29 VTAIL.n28 9.3005
R1959 VTAIL.n12 VTAIL.n11 9.3005
R1960 VTAIL.n35 VTAIL.n34 9.3005
R1961 VTAIL.n37 VTAIL.n36 9.3005
R1962 VTAIL.n38 VTAIL.n7 9.3005
R1963 VTAIL.n107 VTAIL.n106 9.3005
R1964 VTAIL.n58 VTAIL.n57 9.3005
R1965 VTAIL.n101 VTAIL.n100 9.3005
R1966 VTAIL.n99 VTAIL.n98 9.3005
R1967 VTAIL.n75 VTAIL.n74 9.3005
R1968 VTAIL.n70 VTAIL.n69 9.3005
R1969 VTAIL.n81 VTAIL.n80 9.3005
R1970 VTAIL.n83 VTAIL.n82 9.3005
R1971 VTAIL.n66 VTAIL.n65 9.3005
R1972 VTAIL.n89 VTAIL.n88 9.3005
R1973 VTAIL.n91 VTAIL.n90 9.3005
R1974 VTAIL.n92 VTAIL.n61 9.3005
R1975 VTAIL.n163 VTAIL.n162 9.3005
R1976 VTAIL.n114 VTAIL.n113 9.3005
R1977 VTAIL.n157 VTAIL.n156 9.3005
R1978 VTAIL.n155 VTAIL.n154 9.3005
R1979 VTAIL.n131 VTAIL.n130 9.3005
R1980 VTAIL.n126 VTAIL.n125 9.3005
R1981 VTAIL.n137 VTAIL.n136 9.3005
R1982 VTAIL.n139 VTAIL.n138 9.3005
R1983 VTAIL.n122 VTAIL.n121 9.3005
R1984 VTAIL.n145 VTAIL.n144 9.3005
R1985 VTAIL.n147 VTAIL.n146 9.3005
R1986 VTAIL.n148 VTAIL.n117 9.3005
R1987 VTAIL.n352 VTAIL.n351 9.3005
R1988 VTAIL.n347 VTAIL.n346 9.3005
R1989 VTAIL.n358 VTAIL.n357 9.3005
R1990 VTAIL.n360 VTAIL.n359 9.3005
R1991 VTAIL.n343 VTAIL.n342 9.3005
R1992 VTAIL.n366 VTAIL.n365 9.3005
R1993 VTAIL.n368 VTAIL.n367 9.3005
R1994 VTAIL.n340 VTAIL.n337 9.3005
R1995 VTAIL.n383 VTAIL.n382 9.3005
R1996 VTAIL.n334 VTAIL.n333 9.3005
R1997 VTAIL.n377 VTAIL.n376 9.3005
R1998 VTAIL.n375 VTAIL.n374 9.3005
R1999 VTAIL.n296 VTAIL.n295 9.3005
R2000 VTAIL.n291 VTAIL.n290 9.3005
R2001 VTAIL.n302 VTAIL.n301 9.3005
R2002 VTAIL.n304 VTAIL.n303 9.3005
R2003 VTAIL.n287 VTAIL.n286 9.3005
R2004 VTAIL.n310 VTAIL.n309 9.3005
R2005 VTAIL.n312 VTAIL.n311 9.3005
R2006 VTAIL.n284 VTAIL.n281 9.3005
R2007 VTAIL.n327 VTAIL.n326 9.3005
R2008 VTAIL.n278 VTAIL.n277 9.3005
R2009 VTAIL.n321 VTAIL.n320 9.3005
R2010 VTAIL.n319 VTAIL.n318 9.3005
R2011 VTAIL.n242 VTAIL.n241 9.3005
R2012 VTAIL.n237 VTAIL.n236 9.3005
R2013 VTAIL.n248 VTAIL.n247 9.3005
R2014 VTAIL.n250 VTAIL.n249 9.3005
R2015 VTAIL.n233 VTAIL.n232 9.3005
R2016 VTAIL.n256 VTAIL.n255 9.3005
R2017 VTAIL.n258 VTAIL.n257 9.3005
R2018 VTAIL.n230 VTAIL.n227 9.3005
R2019 VTAIL.n273 VTAIL.n272 9.3005
R2020 VTAIL.n224 VTAIL.n223 9.3005
R2021 VTAIL.n267 VTAIL.n266 9.3005
R2022 VTAIL.n265 VTAIL.n264 9.3005
R2023 VTAIL.n186 VTAIL.n185 9.3005
R2024 VTAIL.n181 VTAIL.n180 9.3005
R2025 VTAIL.n192 VTAIL.n191 9.3005
R2026 VTAIL.n194 VTAIL.n193 9.3005
R2027 VTAIL.n177 VTAIL.n176 9.3005
R2028 VTAIL.n200 VTAIL.n199 9.3005
R2029 VTAIL.n202 VTAIL.n201 9.3005
R2030 VTAIL.n174 VTAIL.n171 9.3005
R2031 VTAIL.n217 VTAIL.n216 9.3005
R2032 VTAIL.n168 VTAIL.n167 9.3005
R2033 VTAIL.n211 VTAIL.n210 9.3005
R2034 VTAIL.n209 VTAIL.n208 9.3005
R2035 VTAIL.n410 VTAIL.n409 8.92171
R2036 VTAIL.n26 VTAIL.n25 8.92171
R2037 VTAIL.n80 VTAIL.n79 8.92171
R2038 VTAIL.n136 VTAIL.n135 8.92171
R2039 VTAIL.n357 VTAIL.n356 8.92171
R2040 VTAIL.n301 VTAIL.n300 8.92171
R2041 VTAIL.n247 VTAIL.n246 8.92171
R2042 VTAIL.n191 VTAIL.n190 8.92171
R2043 VTAIL.n406 VTAIL.n400 8.14595
R2044 VTAIL.n22 VTAIL.n16 8.14595
R2045 VTAIL.n76 VTAIL.n70 8.14595
R2046 VTAIL.n132 VTAIL.n126 8.14595
R2047 VTAIL.n353 VTAIL.n347 8.14595
R2048 VTAIL.n297 VTAIL.n291 8.14595
R2049 VTAIL.n243 VTAIL.n237 8.14595
R2050 VTAIL.n187 VTAIL.n181 8.14595
R2051 VTAIL.n405 VTAIL.n402 7.3702
R2052 VTAIL.n21 VTAIL.n18 7.3702
R2053 VTAIL.n75 VTAIL.n72 7.3702
R2054 VTAIL.n131 VTAIL.n128 7.3702
R2055 VTAIL.n352 VTAIL.n349 7.3702
R2056 VTAIL.n296 VTAIL.n293 7.3702
R2057 VTAIL.n242 VTAIL.n239 7.3702
R2058 VTAIL.n186 VTAIL.n183 7.3702
R2059 VTAIL.n406 VTAIL.n405 5.81868
R2060 VTAIL.n22 VTAIL.n21 5.81868
R2061 VTAIL.n76 VTAIL.n75 5.81868
R2062 VTAIL.n132 VTAIL.n131 5.81868
R2063 VTAIL.n353 VTAIL.n352 5.81868
R2064 VTAIL.n297 VTAIL.n296 5.81868
R2065 VTAIL.n243 VTAIL.n242 5.81868
R2066 VTAIL.n187 VTAIL.n186 5.81868
R2067 VTAIL.n409 VTAIL.n400 5.04292
R2068 VTAIL.n25 VTAIL.n16 5.04292
R2069 VTAIL.n79 VTAIL.n70 5.04292
R2070 VTAIL.n135 VTAIL.n126 5.04292
R2071 VTAIL.n356 VTAIL.n347 5.04292
R2072 VTAIL.n300 VTAIL.n291 5.04292
R2073 VTAIL.n246 VTAIL.n237 5.04292
R2074 VTAIL.n190 VTAIL.n181 5.04292
R2075 VTAIL.n410 VTAIL.n398 4.26717
R2076 VTAIL.n26 VTAIL.n14 4.26717
R2077 VTAIL.n80 VTAIL.n68 4.26717
R2078 VTAIL.n136 VTAIL.n124 4.26717
R2079 VTAIL.n357 VTAIL.n345 4.26717
R2080 VTAIL.n301 VTAIL.n289 4.26717
R2081 VTAIL.n247 VTAIL.n235 4.26717
R2082 VTAIL.n191 VTAIL.n179 4.26717
R2083 VTAIL.n414 VTAIL.n413 3.49141
R2084 VTAIL.n438 VTAIL.n386 3.49141
R2085 VTAIL.n30 VTAIL.n29 3.49141
R2086 VTAIL.n54 VTAIL.n2 3.49141
R2087 VTAIL.n84 VTAIL.n83 3.49141
R2088 VTAIL.n108 VTAIL.n56 3.49141
R2089 VTAIL.n140 VTAIL.n139 3.49141
R2090 VTAIL.n164 VTAIL.n112 3.49141
R2091 VTAIL.n384 VTAIL.n332 3.49141
R2092 VTAIL.n361 VTAIL.n360 3.49141
R2093 VTAIL.n328 VTAIL.n276 3.49141
R2094 VTAIL.n305 VTAIL.n304 3.49141
R2095 VTAIL.n274 VTAIL.n222 3.49141
R2096 VTAIL.n251 VTAIL.n250 3.49141
R2097 VTAIL.n218 VTAIL.n166 3.49141
R2098 VTAIL.n195 VTAIL.n194 3.49141
R2099 VTAIL.n404 VTAIL.n403 2.84303
R2100 VTAIL.n20 VTAIL.n19 2.84303
R2101 VTAIL.n74 VTAIL.n73 2.84303
R2102 VTAIL.n130 VTAIL.n129 2.84303
R2103 VTAIL.n351 VTAIL.n350 2.84303
R2104 VTAIL.n295 VTAIL.n294 2.84303
R2105 VTAIL.n241 VTAIL.n240 2.84303
R2106 VTAIL.n185 VTAIL.n184 2.84303
R2107 VTAIL.n417 VTAIL.n396 2.71565
R2108 VTAIL.n436 VTAIL.n435 2.71565
R2109 VTAIL.n33 VTAIL.n12 2.71565
R2110 VTAIL.n52 VTAIL.n51 2.71565
R2111 VTAIL.n87 VTAIL.n66 2.71565
R2112 VTAIL.n106 VTAIL.n105 2.71565
R2113 VTAIL.n143 VTAIL.n122 2.71565
R2114 VTAIL.n162 VTAIL.n161 2.71565
R2115 VTAIL.n382 VTAIL.n381 2.71565
R2116 VTAIL.n364 VTAIL.n343 2.71565
R2117 VTAIL.n326 VTAIL.n325 2.71565
R2118 VTAIL.n308 VTAIL.n287 2.71565
R2119 VTAIL.n272 VTAIL.n271 2.71565
R2120 VTAIL.n254 VTAIL.n233 2.71565
R2121 VTAIL.n216 VTAIL.n215 2.71565
R2122 VTAIL.n198 VTAIL.n177 2.71565
R2123 VTAIL.n221 VTAIL.n219 2.15567
R2124 VTAIL.n275 VTAIL.n221 2.15567
R2125 VTAIL.n331 VTAIL.n329 2.15567
R2126 VTAIL.n385 VTAIL.n331 2.15567
R2127 VTAIL.n165 VTAIL.n111 2.15567
R2128 VTAIL.n111 VTAIL.n109 2.15567
R2129 VTAIL.n55 VTAIL.n1 2.15567
R2130 VTAIL VTAIL.n439 2.09748
R2131 VTAIL.n0 VTAIL.t12 1.95702
R2132 VTAIL.n0 VTAIL.t8 1.95702
R2133 VTAIL.n110 VTAIL.t5 1.95702
R2134 VTAIL.n110 VTAIL.t1 1.95702
R2135 VTAIL.n330 VTAIL.t2 1.95702
R2136 VTAIL.n330 VTAIL.t4 1.95702
R2137 VTAIL.n220 VTAIL.t10 1.95702
R2138 VTAIL.n220 VTAIL.t15 1.95702
R2139 VTAIL.n418 VTAIL.n394 1.93989
R2140 VTAIL.n432 VTAIL.n388 1.93989
R2141 VTAIL.n34 VTAIL.n10 1.93989
R2142 VTAIL.n48 VTAIL.n4 1.93989
R2143 VTAIL.n88 VTAIL.n64 1.93989
R2144 VTAIL.n102 VTAIL.n58 1.93989
R2145 VTAIL.n144 VTAIL.n120 1.93989
R2146 VTAIL.n158 VTAIL.n114 1.93989
R2147 VTAIL.n378 VTAIL.n334 1.93989
R2148 VTAIL.n365 VTAIL.n341 1.93989
R2149 VTAIL.n322 VTAIL.n278 1.93989
R2150 VTAIL.n309 VTAIL.n285 1.93989
R2151 VTAIL.n268 VTAIL.n224 1.93989
R2152 VTAIL.n255 VTAIL.n231 1.93989
R2153 VTAIL.n212 VTAIL.n168 1.93989
R2154 VTAIL.n199 VTAIL.n175 1.93989
R2155 VTAIL.n423 VTAIL.n421 1.16414
R2156 VTAIL.n431 VTAIL.n390 1.16414
R2157 VTAIL.n39 VTAIL.n37 1.16414
R2158 VTAIL.n47 VTAIL.n6 1.16414
R2159 VTAIL.n93 VTAIL.n91 1.16414
R2160 VTAIL.n101 VTAIL.n60 1.16414
R2161 VTAIL.n149 VTAIL.n147 1.16414
R2162 VTAIL.n157 VTAIL.n116 1.16414
R2163 VTAIL.n377 VTAIL.n336 1.16414
R2164 VTAIL.n369 VTAIL.n368 1.16414
R2165 VTAIL.n321 VTAIL.n280 1.16414
R2166 VTAIL.n313 VTAIL.n312 1.16414
R2167 VTAIL.n267 VTAIL.n226 1.16414
R2168 VTAIL.n259 VTAIL.n258 1.16414
R2169 VTAIL.n211 VTAIL.n170 1.16414
R2170 VTAIL.n203 VTAIL.n202 1.16414
R2171 VTAIL.n329 VTAIL.n275 0.470328
R2172 VTAIL.n109 VTAIL.n55 0.470328
R2173 VTAIL.n422 VTAIL.n392 0.388379
R2174 VTAIL.n428 VTAIL.n427 0.388379
R2175 VTAIL.n38 VTAIL.n8 0.388379
R2176 VTAIL.n44 VTAIL.n43 0.388379
R2177 VTAIL.n92 VTAIL.n62 0.388379
R2178 VTAIL.n98 VTAIL.n97 0.388379
R2179 VTAIL.n148 VTAIL.n118 0.388379
R2180 VTAIL.n154 VTAIL.n153 0.388379
R2181 VTAIL.n374 VTAIL.n373 0.388379
R2182 VTAIL.n340 VTAIL.n338 0.388379
R2183 VTAIL.n318 VTAIL.n317 0.388379
R2184 VTAIL.n284 VTAIL.n282 0.388379
R2185 VTAIL.n264 VTAIL.n263 0.388379
R2186 VTAIL.n230 VTAIL.n228 0.388379
R2187 VTAIL.n208 VTAIL.n207 0.388379
R2188 VTAIL.n174 VTAIL.n172 0.388379
R2189 VTAIL.n404 VTAIL.n399 0.155672
R2190 VTAIL.n411 VTAIL.n399 0.155672
R2191 VTAIL.n412 VTAIL.n411 0.155672
R2192 VTAIL.n412 VTAIL.n395 0.155672
R2193 VTAIL.n419 VTAIL.n395 0.155672
R2194 VTAIL.n420 VTAIL.n419 0.155672
R2195 VTAIL.n420 VTAIL.n391 0.155672
R2196 VTAIL.n429 VTAIL.n391 0.155672
R2197 VTAIL.n430 VTAIL.n429 0.155672
R2198 VTAIL.n430 VTAIL.n387 0.155672
R2199 VTAIL.n437 VTAIL.n387 0.155672
R2200 VTAIL.n20 VTAIL.n15 0.155672
R2201 VTAIL.n27 VTAIL.n15 0.155672
R2202 VTAIL.n28 VTAIL.n27 0.155672
R2203 VTAIL.n28 VTAIL.n11 0.155672
R2204 VTAIL.n35 VTAIL.n11 0.155672
R2205 VTAIL.n36 VTAIL.n35 0.155672
R2206 VTAIL.n36 VTAIL.n7 0.155672
R2207 VTAIL.n45 VTAIL.n7 0.155672
R2208 VTAIL.n46 VTAIL.n45 0.155672
R2209 VTAIL.n46 VTAIL.n3 0.155672
R2210 VTAIL.n53 VTAIL.n3 0.155672
R2211 VTAIL.n74 VTAIL.n69 0.155672
R2212 VTAIL.n81 VTAIL.n69 0.155672
R2213 VTAIL.n82 VTAIL.n81 0.155672
R2214 VTAIL.n82 VTAIL.n65 0.155672
R2215 VTAIL.n89 VTAIL.n65 0.155672
R2216 VTAIL.n90 VTAIL.n89 0.155672
R2217 VTAIL.n90 VTAIL.n61 0.155672
R2218 VTAIL.n99 VTAIL.n61 0.155672
R2219 VTAIL.n100 VTAIL.n99 0.155672
R2220 VTAIL.n100 VTAIL.n57 0.155672
R2221 VTAIL.n107 VTAIL.n57 0.155672
R2222 VTAIL.n130 VTAIL.n125 0.155672
R2223 VTAIL.n137 VTAIL.n125 0.155672
R2224 VTAIL.n138 VTAIL.n137 0.155672
R2225 VTAIL.n138 VTAIL.n121 0.155672
R2226 VTAIL.n145 VTAIL.n121 0.155672
R2227 VTAIL.n146 VTAIL.n145 0.155672
R2228 VTAIL.n146 VTAIL.n117 0.155672
R2229 VTAIL.n155 VTAIL.n117 0.155672
R2230 VTAIL.n156 VTAIL.n155 0.155672
R2231 VTAIL.n156 VTAIL.n113 0.155672
R2232 VTAIL.n163 VTAIL.n113 0.155672
R2233 VTAIL.n383 VTAIL.n333 0.155672
R2234 VTAIL.n376 VTAIL.n333 0.155672
R2235 VTAIL.n376 VTAIL.n375 0.155672
R2236 VTAIL.n375 VTAIL.n337 0.155672
R2237 VTAIL.n367 VTAIL.n337 0.155672
R2238 VTAIL.n367 VTAIL.n366 0.155672
R2239 VTAIL.n366 VTAIL.n342 0.155672
R2240 VTAIL.n359 VTAIL.n342 0.155672
R2241 VTAIL.n359 VTAIL.n358 0.155672
R2242 VTAIL.n358 VTAIL.n346 0.155672
R2243 VTAIL.n351 VTAIL.n346 0.155672
R2244 VTAIL.n327 VTAIL.n277 0.155672
R2245 VTAIL.n320 VTAIL.n277 0.155672
R2246 VTAIL.n320 VTAIL.n319 0.155672
R2247 VTAIL.n319 VTAIL.n281 0.155672
R2248 VTAIL.n311 VTAIL.n281 0.155672
R2249 VTAIL.n311 VTAIL.n310 0.155672
R2250 VTAIL.n310 VTAIL.n286 0.155672
R2251 VTAIL.n303 VTAIL.n286 0.155672
R2252 VTAIL.n303 VTAIL.n302 0.155672
R2253 VTAIL.n302 VTAIL.n290 0.155672
R2254 VTAIL.n295 VTAIL.n290 0.155672
R2255 VTAIL.n273 VTAIL.n223 0.155672
R2256 VTAIL.n266 VTAIL.n223 0.155672
R2257 VTAIL.n266 VTAIL.n265 0.155672
R2258 VTAIL.n265 VTAIL.n227 0.155672
R2259 VTAIL.n257 VTAIL.n227 0.155672
R2260 VTAIL.n257 VTAIL.n256 0.155672
R2261 VTAIL.n256 VTAIL.n232 0.155672
R2262 VTAIL.n249 VTAIL.n232 0.155672
R2263 VTAIL.n249 VTAIL.n248 0.155672
R2264 VTAIL.n248 VTAIL.n236 0.155672
R2265 VTAIL.n241 VTAIL.n236 0.155672
R2266 VTAIL.n217 VTAIL.n167 0.155672
R2267 VTAIL.n210 VTAIL.n167 0.155672
R2268 VTAIL.n210 VTAIL.n209 0.155672
R2269 VTAIL.n209 VTAIL.n171 0.155672
R2270 VTAIL.n201 VTAIL.n171 0.155672
R2271 VTAIL.n201 VTAIL.n200 0.155672
R2272 VTAIL.n200 VTAIL.n176 0.155672
R2273 VTAIL.n193 VTAIL.n176 0.155672
R2274 VTAIL.n193 VTAIL.n192 0.155672
R2275 VTAIL.n192 VTAIL.n180 0.155672
R2276 VTAIL.n185 VTAIL.n180 0.155672
R2277 VTAIL VTAIL.n1 0.0586897
R2278 VP.n16 VP.n15 161.3
R2279 VP.n17 VP.n12 161.3
R2280 VP.n19 VP.n18 161.3
R2281 VP.n20 VP.n11 161.3
R2282 VP.n22 VP.n21 161.3
R2283 VP.n24 VP.n10 161.3
R2284 VP.n26 VP.n25 161.3
R2285 VP.n27 VP.n9 161.3
R2286 VP.n29 VP.n28 161.3
R2287 VP.n30 VP.n8 161.3
R2288 VP.n58 VP.n0 161.3
R2289 VP.n57 VP.n56 161.3
R2290 VP.n55 VP.n1 161.3
R2291 VP.n54 VP.n53 161.3
R2292 VP.n52 VP.n2 161.3
R2293 VP.n50 VP.n49 161.3
R2294 VP.n48 VP.n3 161.3
R2295 VP.n47 VP.n46 161.3
R2296 VP.n45 VP.n4 161.3
R2297 VP.n44 VP.n43 161.3
R2298 VP.n42 VP.n41 161.3
R2299 VP.n40 VP.n6 161.3
R2300 VP.n39 VP.n38 161.3
R2301 VP.n37 VP.n7 161.3
R2302 VP.n36 VP.n35 161.3
R2303 VP.n14 VP.t1 144.47
R2304 VP.n34 VP.t2 112.394
R2305 VP.n5 VP.t6 112.394
R2306 VP.n51 VP.t4 112.394
R2307 VP.n59 VP.t7 112.394
R2308 VP.n31 VP.t3 112.394
R2309 VP.n23 VP.t0 112.394
R2310 VP.n13 VP.t5 112.394
R2311 VP.n34 VP.n33 98.6123
R2312 VP.n60 VP.n59 98.6123
R2313 VP.n32 VP.n31 98.6123
R2314 VP.n14 VP.n13 59.4159
R2315 VP.n33 VP.n32 47.4087
R2316 VP.n39 VP.n7 40.577
R2317 VP.n40 VP.n39 40.577
R2318 VP.n46 VP.n45 40.577
R2319 VP.n46 VP.n3 40.577
R2320 VP.n53 VP.n1 40.577
R2321 VP.n57 VP.n1 40.577
R2322 VP.n29 VP.n9 40.577
R2323 VP.n25 VP.n9 40.577
R2324 VP.n18 VP.n11 40.577
R2325 VP.n18 VP.n17 40.577
R2326 VP.n35 VP.n7 24.5923
R2327 VP.n41 VP.n40 24.5923
R2328 VP.n45 VP.n44 24.5923
R2329 VP.n50 VP.n3 24.5923
R2330 VP.n53 VP.n52 24.5923
R2331 VP.n58 VP.n57 24.5923
R2332 VP.n30 VP.n29 24.5923
R2333 VP.n22 VP.n11 24.5923
R2334 VP.n25 VP.n24 24.5923
R2335 VP.n17 VP.n16 24.5923
R2336 VP.n35 VP.n34 12.2964
R2337 VP.n41 VP.n5 12.2964
R2338 VP.n44 VP.n5 12.2964
R2339 VP.n51 VP.n50 12.2964
R2340 VP.n52 VP.n51 12.2964
R2341 VP.n59 VP.n58 12.2964
R2342 VP.n31 VP.n30 12.2964
R2343 VP.n23 VP.n22 12.2964
R2344 VP.n24 VP.n23 12.2964
R2345 VP.n16 VP.n13 12.2964
R2346 VP.n15 VP.n14 9.706
R2347 VP.n32 VP.n8 0.278335
R2348 VP.n36 VP.n33 0.278335
R2349 VP.n60 VP.n0 0.278335
R2350 VP.n15 VP.n12 0.189894
R2351 VP.n19 VP.n12 0.189894
R2352 VP.n20 VP.n19 0.189894
R2353 VP.n21 VP.n20 0.189894
R2354 VP.n21 VP.n10 0.189894
R2355 VP.n26 VP.n10 0.189894
R2356 VP.n27 VP.n26 0.189894
R2357 VP.n28 VP.n27 0.189894
R2358 VP.n28 VP.n8 0.189894
R2359 VP.n37 VP.n36 0.189894
R2360 VP.n38 VP.n37 0.189894
R2361 VP.n38 VP.n6 0.189894
R2362 VP.n42 VP.n6 0.189894
R2363 VP.n43 VP.n42 0.189894
R2364 VP.n43 VP.n4 0.189894
R2365 VP.n47 VP.n4 0.189894
R2366 VP.n48 VP.n47 0.189894
R2367 VP.n49 VP.n48 0.189894
R2368 VP.n49 VP.n2 0.189894
R2369 VP.n54 VP.n2 0.189894
R2370 VP.n55 VP.n54 0.189894
R2371 VP.n56 VP.n55 0.189894
R2372 VP.n56 VP.n0 0.189894
R2373 VP VP.n60 0.153485
R2374 VDD1 VDD1.n0 66.8791
R2375 VDD1.n3 VDD1.n2 66.7654
R2376 VDD1.n3 VDD1.n1 66.7654
R2377 VDD1.n5 VDD1.n4 65.7432
R2378 VDD1.n5 VDD1.n3 42.7207
R2379 VDD1.n4 VDD1.t7 1.95702
R2380 VDD1.n4 VDD1.t4 1.95702
R2381 VDD1.n0 VDD1.t6 1.95702
R2382 VDD1.n0 VDD1.t2 1.95702
R2383 VDD1.n2 VDD1.t3 1.95702
R2384 VDD1.n2 VDD1.t0 1.95702
R2385 VDD1.n1 VDD1.t5 1.95702
R2386 VDD1.n1 VDD1.t1 1.95702
R2387 VDD1 VDD1.n5 1.0199
C0 VN VDD2 7.13239f
C1 VTAIL VDD2 7.41598f
C2 VDD1 VDD2 1.55004f
C3 VN VTAIL 7.46368f
C4 VN VDD1 0.150774f
C5 VTAIL VDD1 7.36445f
C6 VP VDD2 0.473738f
C7 VP VN 6.78734f
C8 VP VTAIL 7.47778f
C9 VP VDD1 7.45418f
C10 VDD2 B 4.775568f
C11 VDD1 B 5.172893f
C12 VTAIL B 9.06145f
C13 VN B 13.72334f
C14 VP B 12.286482f
C15 VDD1.t6 B 0.199114f
C16 VDD1.t2 B 0.199114f
C17 VDD1.n0 B 1.76527f
C18 VDD1.t5 B 0.199114f
C19 VDD1.t1 B 0.199114f
C20 VDD1.n1 B 1.76434f
C21 VDD1.t3 B 0.199114f
C22 VDD1.t0 B 0.199114f
C23 VDD1.n2 B 1.76434f
C24 VDD1.n3 B 2.94474f
C25 VDD1.t7 B 0.199114f
C26 VDD1.t4 B 0.199114f
C27 VDD1.n4 B 1.7572f
C28 VDD1.n5 B 2.67157f
C29 VP.n0 B 0.034063f
C30 VP.t7 B 1.53779f
C31 VP.n1 B 0.020869f
C32 VP.n2 B 0.025838f
C33 VP.t4 B 1.53779f
C34 VP.n3 B 0.051083f
C35 VP.n4 B 0.025838f
C36 VP.t6 B 1.53779f
C37 VP.n5 B 0.55371f
C38 VP.n6 B 0.025838f
C39 VP.n7 B 0.051083f
C40 VP.n8 B 0.034063f
C41 VP.t3 B 1.53779f
C42 VP.n9 B 0.020869f
C43 VP.n10 B 0.025838f
C44 VP.t0 B 1.53779f
C45 VP.n11 B 0.051083f
C46 VP.n12 B 0.025838f
C47 VP.t5 B 1.53779f
C48 VP.n13 B 0.619425f
C49 VP.t1 B 1.69073f
C50 VP.n14 B 0.612745f
C51 VP.n15 B 0.21898f
C52 VP.n16 B 0.036087f
C53 VP.n17 B 0.051083f
C54 VP.n18 B 0.020869f
C55 VP.n19 B 0.025838f
C56 VP.n20 B 0.025838f
C57 VP.n21 B 0.025838f
C58 VP.n22 B 0.036087f
C59 VP.n23 B 0.55371f
C60 VP.n24 B 0.036087f
C61 VP.n25 B 0.051083f
C62 VP.n26 B 0.025838f
C63 VP.n27 B 0.025838f
C64 VP.n28 B 0.025838f
C65 VP.n29 B 0.051083f
C66 VP.n30 B 0.036087f
C67 VP.n31 B 0.627798f
C68 VP.n32 B 1.32223f
C69 VP.n33 B 1.34188f
C70 VP.t2 B 1.53779f
C71 VP.n34 B 0.627798f
C72 VP.n35 B 0.036087f
C73 VP.n36 B 0.034063f
C74 VP.n37 B 0.025838f
C75 VP.n38 B 0.025838f
C76 VP.n39 B 0.020869f
C77 VP.n40 B 0.051083f
C78 VP.n41 B 0.036087f
C79 VP.n42 B 0.025838f
C80 VP.n43 B 0.025838f
C81 VP.n44 B 0.036087f
C82 VP.n45 B 0.051083f
C83 VP.n46 B 0.020869f
C84 VP.n47 B 0.025838f
C85 VP.n48 B 0.025838f
C86 VP.n49 B 0.025838f
C87 VP.n50 B 0.036087f
C88 VP.n51 B 0.55371f
C89 VP.n52 B 0.036087f
C90 VP.n53 B 0.051083f
C91 VP.n54 B 0.025838f
C92 VP.n55 B 0.025838f
C93 VP.n56 B 0.025838f
C94 VP.n57 B 0.051083f
C95 VP.n58 B 0.036087f
C96 VP.n59 B 0.627798f
C97 VP.n60 B 0.037335f
C98 VTAIL.t12 B 0.161292f
C99 VTAIL.t8 B 0.161292f
C100 VTAIL.n0 B 1.36944f
C101 VTAIL.n1 B 0.333028f
C102 VTAIL.n2 B 0.028893f
C103 VTAIL.n3 B 0.020169f
C104 VTAIL.n4 B 0.010838f
C105 VTAIL.n5 B 0.025617f
C106 VTAIL.n6 B 0.011475f
C107 VTAIL.n7 B 0.020169f
C108 VTAIL.n8 B 0.011157f
C109 VTAIL.n9 B 0.025617f
C110 VTAIL.n10 B 0.011475f
C111 VTAIL.n11 B 0.020169f
C112 VTAIL.n12 B 0.010838f
C113 VTAIL.n13 B 0.025617f
C114 VTAIL.n14 B 0.011475f
C115 VTAIL.n15 B 0.020169f
C116 VTAIL.n16 B 0.010838f
C117 VTAIL.n17 B 0.019212f
C118 VTAIL.n18 B 0.018109f
C119 VTAIL.t9 B 0.043063f
C120 VTAIL.n19 B 0.130861f
C121 VTAIL.n20 B 0.848822f
C122 VTAIL.n21 B 0.010838f
C123 VTAIL.n22 B 0.011475f
C124 VTAIL.n23 B 0.025617f
C125 VTAIL.n24 B 0.025617f
C126 VTAIL.n25 B 0.011475f
C127 VTAIL.n26 B 0.010838f
C128 VTAIL.n27 B 0.020169f
C129 VTAIL.n28 B 0.020169f
C130 VTAIL.n29 B 0.010838f
C131 VTAIL.n30 B 0.011475f
C132 VTAIL.n31 B 0.025617f
C133 VTAIL.n32 B 0.025617f
C134 VTAIL.n33 B 0.011475f
C135 VTAIL.n34 B 0.010838f
C136 VTAIL.n35 B 0.020169f
C137 VTAIL.n36 B 0.020169f
C138 VTAIL.n37 B 0.010838f
C139 VTAIL.n38 B 0.010838f
C140 VTAIL.n39 B 0.011475f
C141 VTAIL.n40 B 0.025617f
C142 VTAIL.n41 B 0.025617f
C143 VTAIL.n42 B 0.025617f
C144 VTAIL.n43 B 0.011157f
C145 VTAIL.n44 B 0.010838f
C146 VTAIL.n45 B 0.020169f
C147 VTAIL.n46 B 0.020169f
C148 VTAIL.n47 B 0.010838f
C149 VTAIL.n48 B 0.011475f
C150 VTAIL.n49 B 0.025617f
C151 VTAIL.n50 B 0.056418f
C152 VTAIL.n51 B 0.011475f
C153 VTAIL.n52 B 0.010838f
C154 VTAIL.n53 B 0.051027f
C155 VTAIL.n54 B 0.031797f
C156 VTAIL.n55 B 0.190313f
C157 VTAIL.n56 B 0.028893f
C158 VTAIL.n57 B 0.020169f
C159 VTAIL.n58 B 0.010838f
C160 VTAIL.n59 B 0.025617f
C161 VTAIL.n60 B 0.011475f
C162 VTAIL.n61 B 0.020169f
C163 VTAIL.n62 B 0.011157f
C164 VTAIL.n63 B 0.025617f
C165 VTAIL.n64 B 0.011475f
C166 VTAIL.n65 B 0.020169f
C167 VTAIL.n66 B 0.010838f
C168 VTAIL.n67 B 0.025617f
C169 VTAIL.n68 B 0.011475f
C170 VTAIL.n69 B 0.020169f
C171 VTAIL.n70 B 0.010838f
C172 VTAIL.n71 B 0.019212f
C173 VTAIL.n72 B 0.018109f
C174 VTAIL.t0 B 0.043063f
C175 VTAIL.n73 B 0.130861f
C176 VTAIL.n74 B 0.848822f
C177 VTAIL.n75 B 0.010838f
C178 VTAIL.n76 B 0.011475f
C179 VTAIL.n77 B 0.025617f
C180 VTAIL.n78 B 0.025617f
C181 VTAIL.n79 B 0.011475f
C182 VTAIL.n80 B 0.010838f
C183 VTAIL.n81 B 0.020169f
C184 VTAIL.n82 B 0.020169f
C185 VTAIL.n83 B 0.010838f
C186 VTAIL.n84 B 0.011475f
C187 VTAIL.n85 B 0.025617f
C188 VTAIL.n86 B 0.025617f
C189 VTAIL.n87 B 0.011475f
C190 VTAIL.n88 B 0.010838f
C191 VTAIL.n89 B 0.020169f
C192 VTAIL.n90 B 0.020169f
C193 VTAIL.n91 B 0.010838f
C194 VTAIL.n92 B 0.010838f
C195 VTAIL.n93 B 0.011475f
C196 VTAIL.n94 B 0.025617f
C197 VTAIL.n95 B 0.025617f
C198 VTAIL.n96 B 0.025617f
C199 VTAIL.n97 B 0.011157f
C200 VTAIL.n98 B 0.010838f
C201 VTAIL.n99 B 0.020169f
C202 VTAIL.n100 B 0.020169f
C203 VTAIL.n101 B 0.010838f
C204 VTAIL.n102 B 0.011475f
C205 VTAIL.n103 B 0.025617f
C206 VTAIL.n104 B 0.056418f
C207 VTAIL.n105 B 0.011475f
C208 VTAIL.n106 B 0.010838f
C209 VTAIL.n107 B 0.051027f
C210 VTAIL.n108 B 0.031797f
C211 VTAIL.n109 B 0.190313f
C212 VTAIL.t5 B 0.161292f
C213 VTAIL.t1 B 0.161292f
C214 VTAIL.n110 B 1.36944f
C215 VTAIL.n111 B 0.469307f
C216 VTAIL.n112 B 0.028893f
C217 VTAIL.n113 B 0.020169f
C218 VTAIL.n114 B 0.010838f
C219 VTAIL.n115 B 0.025617f
C220 VTAIL.n116 B 0.011475f
C221 VTAIL.n117 B 0.020169f
C222 VTAIL.n118 B 0.011157f
C223 VTAIL.n119 B 0.025617f
C224 VTAIL.n120 B 0.011475f
C225 VTAIL.n121 B 0.020169f
C226 VTAIL.n122 B 0.010838f
C227 VTAIL.n123 B 0.025617f
C228 VTAIL.n124 B 0.011475f
C229 VTAIL.n125 B 0.020169f
C230 VTAIL.n126 B 0.010838f
C231 VTAIL.n127 B 0.019212f
C232 VTAIL.n128 B 0.018109f
C233 VTAIL.t6 B 0.043063f
C234 VTAIL.n129 B 0.130861f
C235 VTAIL.n130 B 0.848822f
C236 VTAIL.n131 B 0.010838f
C237 VTAIL.n132 B 0.011475f
C238 VTAIL.n133 B 0.025617f
C239 VTAIL.n134 B 0.025617f
C240 VTAIL.n135 B 0.011475f
C241 VTAIL.n136 B 0.010838f
C242 VTAIL.n137 B 0.020169f
C243 VTAIL.n138 B 0.020169f
C244 VTAIL.n139 B 0.010838f
C245 VTAIL.n140 B 0.011475f
C246 VTAIL.n141 B 0.025617f
C247 VTAIL.n142 B 0.025617f
C248 VTAIL.n143 B 0.011475f
C249 VTAIL.n144 B 0.010838f
C250 VTAIL.n145 B 0.020169f
C251 VTAIL.n146 B 0.020169f
C252 VTAIL.n147 B 0.010838f
C253 VTAIL.n148 B 0.010838f
C254 VTAIL.n149 B 0.011475f
C255 VTAIL.n150 B 0.025617f
C256 VTAIL.n151 B 0.025617f
C257 VTAIL.n152 B 0.025617f
C258 VTAIL.n153 B 0.011157f
C259 VTAIL.n154 B 0.010838f
C260 VTAIL.n155 B 0.020169f
C261 VTAIL.n156 B 0.020169f
C262 VTAIL.n157 B 0.010838f
C263 VTAIL.n158 B 0.011475f
C264 VTAIL.n159 B 0.025617f
C265 VTAIL.n160 B 0.056418f
C266 VTAIL.n161 B 0.011475f
C267 VTAIL.n162 B 0.010838f
C268 VTAIL.n163 B 0.051027f
C269 VTAIL.n164 B 0.031797f
C270 VTAIL.n165 B 1.14077f
C271 VTAIL.n166 B 0.028893f
C272 VTAIL.n167 B 0.020169f
C273 VTAIL.n168 B 0.010838f
C274 VTAIL.n169 B 0.025617f
C275 VTAIL.n170 B 0.011475f
C276 VTAIL.n171 B 0.020169f
C277 VTAIL.n172 B 0.011157f
C278 VTAIL.n173 B 0.025617f
C279 VTAIL.n174 B 0.010838f
C280 VTAIL.n175 B 0.011475f
C281 VTAIL.n176 B 0.020169f
C282 VTAIL.n177 B 0.010838f
C283 VTAIL.n178 B 0.025617f
C284 VTAIL.n179 B 0.011475f
C285 VTAIL.n180 B 0.020169f
C286 VTAIL.n181 B 0.010838f
C287 VTAIL.n182 B 0.019212f
C288 VTAIL.n183 B 0.018109f
C289 VTAIL.t14 B 0.043063f
C290 VTAIL.n184 B 0.130861f
C291 VTAIL.n185 B 0.848822f
C292 VTAIL.n186 B 0.010838f
C293 VTAIL.n187 B 0.011475f
C294 VTAIL.n188 B 0.025617f
C295 VTAIL.n189 B 0.025617f
C296 VTAIL.n190 B 0.011475f
C297 VTAIL.n191 B 0.010838f
C298 VTAIL.n192 B 0.020169f
C299 VTAIL.n193 B 0.020169f
C300 VTAIL.n194 B 0.010838f
C301 VTAIL.n195 B 0.011475f
C302 VTAIL.n196 B 0.025617f
C303 VTAIL.n197 B 0.025617f
C304 VTAIL.n198 B 0.011475f
C305 VTAIL.n199 B 0.010838f
C306 VTAIL.n200 B 0.020169f
C307 VTAIL.n201 B 0.020169f
C308 VTAIL.n202 B 0.010838f
C309 VTAIL.n203 B 0.011475f
C310 VTAIL.n204 B 0.025617f
C311 VTAIL.n205 B 0.025617f
C312 VTAIL.n206 B 0.025617f
C313 VTAIL.n207 B 0.011157f
C314 VTAIL.n208 B 0.010838f
C315 VTAIL.n209 B 0.020169f
C316 VTAIL.n210 B 0.020169f
C317 VTAIL.n211 B 0.010838f
C318 VTAIL.n212 B 0.011475f
C319 VTAIL.n213 B 0.025617f
C320 VTAIL.n214 B 0.056418f
C321 VTAIL.n215 B 0.011475f
C322 VTAIL.n216 B 0.010838f
C323 VTAIL.n217 B 0.051027f
C324 VTAIL.n218 B 0.031797f
C325 VTAIL.n219 B 1.14077f
C326 VTAIL.t10 B 0.161292f
C327 VTAIL.t15 B 0.161292f
C328 VTAIL.n220 B 1.36945f
C329 VTAIL.n221 B 0.469299f
C330 VTAIL.n222 B 0.028893f
C331 VTAIL.n223 B 0.020169f
C332 VTAIL.n224 B 0.010838f
C333 VTAIL.n225 B 0.025617f
C334 VTAIL.n226 B 0.011475f
C335 VTAIL.n227 B 0.020169f
C336 VTAIL.n228 B 0.011157f
C337 VTAIL.n229 B 0.025617f
C338 VTAIL.n230 B 0.010838f
C339 VTAIL.n231 B 0.011475f
C340 VTAIL.n232 B 0.020169f
C341 VTAIL.n233 B 0.010838f
C342 VTAIL.n234 B 0.025617f
C343 VTAIL.n235 B 0.011475f
C344 VTAIL.n236 B 0.020169f
C345 VTAIL.n237 B 0.010838f
C346 VTAIL.n238 B 0.019212f
C347 VTAIL.n239 B 0.018109f
C348 VTAIL.t11 B 0.043063f
C349 VTAIL.n240 B 0.130861f
C350 VTAIL.n241 B 0.848822f
C351 VTAIL.n242 B 0.010838f
C352 VTAIL.n243 B 0.011475f
C353 VTAIL.n244 B 0.025617f
C354 VTAIL.n245 B 0.025617f
C355 VTAIL.n246 B 0.011475f
C356 VTAIL.n247 B 0.010838f
C357 VTAIL.n248 B 0.020169f
C358 VTAIL.n249 B 0.020169f
C359 VTAIL.n250 B 0.010838f
C360 VTAIL.n251 B 0.011475f
C361 VTAIL.n252 B 0.025617f
C362 VTAIL.n253 B 0.025617f
C363 VTAIL.n254 B 0.011475f
C364 VTAIL.n255 B 0.010838f
C365 VTAIL.n256 B 0.020169f
C366 VTAIL.n257 B 0.020169f
C367 VTAIL.n258 B 0.010838f
C368 VTAIL.n259 B 0.011475f
C369 VTAIL.n260 B 0.025617f
C370 VTAIL.n261 B 0.025617f
C371 VTAIL.n262 B 0.025617f
C372 VTAIL.n263 B 0.011157f
C373 VTAIL.n264 B 0.010838f
C374 VTAIL.n265 B 0.020169f
C375 VTAIL.n266 B 0.020169f
C376 VTAIL.n267 B 0.010838f
C377 VTAIL.n268 B 0.011475f
C378 VTAIL.n269 B 0.025617f
C379 VTAIL.n270 B 0.056418f
C380 VTAIL.n271 B 0.011475f
C381 VTAIL.n272 B 0.010838f
C382 VTAIL.n273 B 0.051027f
C383 VTAIL.n274 B 0.031797f
C384 VTAIL.n275 B 0.190313f
C385 VTAIL.n276 B 0.028893f
C386 VTAIL.n277 B 0.020169f
C387 VTAIL.n278 B 0.010838f
C388 VTAIL.n279 B 0.025617f
C389 VTAIL.n280 B 0.011475f
C390 VTAIL.n281 B 0.020169f
C391 VTAIL.n282 B 0.011157f
C392 VTAIL.n283 B 0.025617f
C393 VTAIL.n284 B 0.010838f
C394 VTAIL.n285 B 0.011475f
C395 VTAIL.n286 B 0.020169f
C396 VTAIL.n287 B 0.010838f
C397 VTAIL.n288 B 0.025617f
C398 VTAIL.n289 B 0.011475f
C399 VTAIL.n290 B 0.020169f
C400 VTAIL.n291 B 0.010838f
C401 VTAIL.n292 B 0.019212f
C402 VTAIL.n293 B 0.018109f
C403 VTAIL.t7 B 0.043063f
C404 VTAIL.n294 B 0.130861f
C405 VTAIL.n295 B 0.848822f
C406 VTAIL.n296 B 0.010838f
C407 VTAIL.n297 B 0.011475f
C408 VTAIL.n298 B 0.025617f
C409 VTAIL.n299 B 0.025617f
C410 VTAIL.n300 B 0.011475f
C411 VTAIL.n301 B 0.010838f
C412 VTAIL.n302 B 0.020169f
C413 VTAIL.n303 B 0.020169f
C414 VTAIL.n304 B 0.010838f
C415 VTAIL.n305 B 0.011475f
C416 VTAIL.n306 B 0.025617f
C417 VTAIL.n307 B 0.025617f
C418 VTAIL.n308 B 0.011475f
C419 VTAIL.n309 B 0.010838f
C420 VTAIL.n310 B 0.020169f
C421 VTAIL.n311 B 0.020169f
C422 VTAIL.n312 B 0.010838f
C423 VTAIL.n313 B 0.011475f
C424 VTAIL.n314 B 0.025617f
C425 VTAIL.n315 B 0.025617f
C426 VTAIL.n316 B 0.025617f
C427 VTAIL.n317 B 0.011157f
C428 VTAIL.n318 B 0.010838f
C429 VTAIL.n319 B 0.020169f
C430 VTAIL.n320 B 0.020169f
C431 VTAIL.n321 B 0.010838f
C432 VTAIL.n322 B 0.011475f
C433 VTAIL.n323 B 0.025617f
C434 VTAIL.n324 B 0.056418f
C435 VTAIL.n325 B 0.011475f
C436 VTAIL.n326 B 0.010838f
C437 VTAIL.n327 B 0.051027f
C438 VTAIL.n328 B 0.031797f
C439 VTAIL.n329 B 0.190313f
C440 VTAIL.t2 B 0.161292f
C441 VTAIL.t4 B 0.161292f
C442 VTAIL.n330 B 1.36945f
C443 VTAIL.n331 B 0.469299f
C444 VTAIL.n332 B 0.028893f
C445 VTAIL.n333 B 0.020169f
C446 VTAIL.n334 B 0.010838f
C447 VTAIL.n335 B 0.025617f
C448 VTAIL.n336 B 0.011475f
C449 VTAIL.n337 B 0.020169f
C450 VTAIL.n338 B 0.011157f
C451 VTAIL.n339 B 0.025617f
C452 VTAIL.n340 B 0.010838f
C453 VTAIL.n341 B 0.011475f
C454 VTAIL.n342 B 0.020169f
C455 VTAIL.n343 B 0.010838f
C456 VTAIL.n344 B 0.025617f
C457 VTAIL.n345 B 0.011475f
C458 VTAIL.n346 B 0.020169f
C459 VTAIL.n347 B 0.010838f
C460 VTAIL.n348 B 0.019212f
C461 VTAIL.n349 B 0.018109f
C462 VTAIL.t3 B 0.043063f
C463 VTAIL.n350 B 0.130861f
C464 VTAIL.n351 B 0.848822f
C465 VTAIL.n352 B 0.010838f
C466 VTAIL.n353 B 0.011475f
C467 VTAIL.n354 B 0.025617f
C468 VTAIL.n355 B 0.025617f
C469 VTAIL.n356 B 0.011475f
C470 VTAIL.n357 B 0.010838f
C471 VTAIL.n358 B 0.020169f
C472 VTAIL.n359 B 0.020169f
C473 VTAIL.n360 B 0.010838f
C474 VTAIL.n361 B 0.011475f
C475 VTAIL.n362 B 0.025617f
C476 VTAIL.n363 B 0.025617f
C477 VTAIL.n364 B 0.011475f
C478 VTAIL.n365 B 0.010838f
C479 VTAIL.n366 B 0.020169f
C480 VTAIL.n367 B 0.020169f
C481 VTAIL.n368 B 0.010838f
C482 VTAIL.n369 B 0.011475f
C483 VTAIL.n370 B 0.025617f
C484 VTAIL.n371 B 0.025617f
C485 VTAIL.n372 B 0.025617f
C486 VTAIL.n373 B 0.011157f
C487 VTAIL.n374 B 0.010838f
C488 VTAIL.n375 B 0.020169f
C489 VTAIL.n376 B 0.020169f
C490 VTAIL.n377 B 0.010838f
C491 VTAIL.n378 B 0.011475f
C492 VTAIL.n379 B 0.025617f
C493 VTAIL.n380 B 0.056418f
C494 VTAIL.n381 B 0.011475f
C495 VTAIL.n382 B 0.010838f
C496 VTAIL.n383 B 0.051027f
C497 VTAIL.n384 B 0.031797f
C498 VTAIL.n385 B 1.14077f
C499 VTAIL.n386 B 0.028893f
C500 VTAIL.n387 B 0.020169f
C501 VTAIL.n388 B 0.010838f
C502 VTAIL.n389 B 0.025617f
C503 VTAIL.n390 B 0.011475f
C504 VTAIL.n391 B 0.020169f
C505 VTAIL.n392 B 0.011157f
C506 VTAIL.n393 B 0.025617f
C507 VTAIL.n394 B 0.011475f
C508 VTAIL.n395 B 0.020169f
C509 VTAIL.n396 B 0.010838f
C510 VTAIL.n397 B 0.025617f
C511 VTAIL.n398 B 0.011475f
C512 VTAIL.n399 B 0.020169f
C513 VTAIL.n400 B 0.010838f
C514 VTAIL.n401 B 0.019212f
C515 VTAIL.n402 B 0.018109f
C516 VTAIL.t13 B 0.043063f
C517 VTAIL.n403 B 0.130861f
C518 VTAIL.n404 B 0.848822f
C519 VTAIL.n405 B 0.010838f
C520 VTAIL.n406 B 0.011475f
C521 VTAIL.n407 B 0.025617f
C522 VTAIL.n408 B 0.025617f
C523 VTAIL.n409 B 0.011475f
C524 VTAIL.n410 B 0.010838f
C525 VTAIL.n411 B 0.020169f
C526 VTAIL.n412 B 0.020169f
C527 VTAIL.n413 B 0.010838f
C528 VTAIL.n414 B 0.011475f
C529 VTAIL.n415 B 0.025617f
C530 VTAIL.n416 B 0.025617f
C531 VTAIL.n417 B 0.011475f
C532 VTAIL.n418 B 0.010838f
C533 VTAIL.n419 B 0.020169f
C534 VTAIL.n420 B 0.020169f
C535 VTAIL.n421 B 0.010838f
C536 VTAIL.n422 B 0.010838f
C537 VTAIL.n423 B 0.011475f
C538 VTAIL.n424 B 0.025617f
C539 VTAIL.n425 B 0.025617f
C540 VTAIL.n426 B 0.025617f
C541 VTAIL.n427 B 0.011157f
C542 VTAIL.n428 B 0.010838f
C543 VTAIL.n429 B 0.020169f
C544 VTAIL.n430 B 0.020169f
C545 VTAIL.n431 B 0.010838f
C546 VTAIL.n432 B 0.011475f
C547 VTAIL.n433 B 0.025617f
C548 VTAIL.n434 B 0.056418f
C549 VTAIL.n435 B 0.011475f
C550 VTAIL.n436 B 0.010838f
C551 VTAIL.n437 B 0.051027f
C552 VTAIL.n438 B 0.031797f
C553 VTAIL.n439 B 1.13699f
C554 VDD2.t1 B 0.194972f
C555 VDD2.t5 B 0.194972f
C556 VDD2.n0 B 1.72764f
C557 VDD2.t7 B 0.194972f
C558 VDD2.t0 B 0.194972f
C559 VDD2.n1 B 1.72764f
C560 VDD2.n2 B 2.83238f
C561 VDD2.t4 B 0.194972f
C562 VDD2.t2 B 0.194972f
C563 VDD2.n3 B 1.72065f
C564 VDD2.n4 B 2.58618f
C565 VDD2.t3 B 0.194972f
C566 VDD2.t6 B 0.194972f
C567 VDD2.n5 B 1.7276f
C568 VN.n0 B 0.033382f
C569 VN.t2 B 1.50706f
C570 VN.n1 B 0.020452f
C571 VN.n2 B 0.025322f
C572 VN.t7 B 1.50706f
C573 VN.n3 B 0.050062f
C574 VN.n4 B 0.025322f
C575 VN.t3 B 1.50706f
C576 VN.n5 B 0.607048f
C577 VN.t6 B 1.65695f
C578 VN.n6 B 0.600502f
C579 VN.n7 B 0.214604f
C580 VN.n8 B 0.035366f
C581 VN.n9 B 0.050062f
C582 VN.n10 B 0.020452f
C583 VN.n11 B 0.025322f
C584 VN.n12 B 0.025322f
C585 VN.n13 B 0.025322f
C586 VN.n14 B 0.035366f
C587 VN.n15 B 0.542646f
C588 VN.n16 B 0.035366f
C589 VN.n17 B 0.050062f
C590 VN.n18 B 0.025322f
C591 VN.n19 B 0.025322f
C592 VN.n20 B 0.025322f
C593 VN.n21 B 0.050062f
C594 VN.n22 B 0.035366f
C595 VN.n23 B 0.615254f
C596 VN.n24 B 0.036589f
C597 VN.n25 B 0.033382f
C598 VN.t1 B 1.50706f
C599 VN.n26 B 0.020452f
C600 VN.n27 B 0.025322f
C601 VN.t5 B 1.50706f
C602 VN.n28 B 0.050062f
C603 VN.n29 B 0.025322f
C604 VN.t0 B 1.50706f
C605 VN.n30 B 0.607048f
C606 VN.t4 B 1.65695f
C607 VN.n31 B 0.600502f
C608 VN.n32 B 0.214604f
C609 VN.n33 B 0.035366f
C610 VN.n34 B 0.050062f
C611 VN.n35 B 0.020452f
C612 VN.n36 B 0.025322f
C613 VN.n37 B 0.025322f
C614 VN.n38 B 0.025322f
C615 VN.n39 B 0.035366f
C616 VN.n40 B 0.542646f
C617 VN.n41 B 0.035366f
C618 VN.n42 B 0.050062f
C619 VN.n43 B 0.025322f
C620 VN.n44 B 0.025322f
C621 VN.n45 B 0.025322f
C622 VN.n46 B 0.050062f
C623 VN.n47 B 0.035366f
C624 VN.n48 B 0.615254f
C625 VN.n49 B 1.30953f
.ends

