* NGSPICE file created from diff_pair_sample_0322.ext - technology: sky130A

.subckt diff_pair_sample_0322 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VP.t0 VDD1.t3 w_n4170_n3652# sky130_fd_pr__pfet_01v8 ad=5.2338 pd=27.62 as=2.2143 ps=13.75 w=13.42 l=2.87
X1 B.t11 B.t9 B.t10 w_n4170_n3652# sky130_fd_pr__pfet_01v8 ad=5.2338 pd=27.62 as=0 ps=0 w=13.42 l=2.87
X2 VTAIL.t3 VN.t0 VDD2.t7 w_n4170_n3652# sky130_fd_pr__pfet_01v8 ad=5.2338 pd=27.62 as=2.2143 ps=13.75 w=13.42 l=2.87
X3 VDD1.t5 VP.t1 VTAIL.t14 w_n4170_n3652# sky130_fd_pr__pfet_01v8 ad=2.2143 pd=13.75 as=5.2338 ps=27.62 w=13.42 l=2.87
X4 VDD1.t6 VP.t2 VTAIL.t13 w_n4170_n3652# sky130_fd_pr__pfet_01v8 ad=2.2143 pd=13.75 as=2.2143 ps=13.75 w=13.42 l=2.87
X5 VDD2.t6 VN.t1 VTAIL.t6 w_n4170_n3652# sky130_fd_pr__pfet_01v8 ad=2.2143 pd=13.75 as=2.2143 ps=13.75 w=13.42 l=2.87
X6 VDD1.t0 VP.t3 VTAIL.t12 w_n4170_n3652# sky130_fd_pr__pfet_01v8 ad=2.2143 pd=13.75 as=2.2143 ps=13.75 w=13.42 l=2.87
X7 VTAIL.t11 VP.t4 VDD1.t1 w_n4170_n3652# sky130_fd_pr__pfet_01v8 ad=2.2143 pd=13.75 as=2.2143 ps=13.75 w=13.42 l=2.87
X8 B.t8 B.t6 B.t7 w_n4170_n3652# sky130_fd_pr__pfet_01v8 ad=5.2338 pd=27.62 as=0 ps=0 w=13.42 l=2.87
X9 VTAIL.t7 VN.t2 VDD2.t5 w_n4170_n3652# sky130_fd_pr__pfet_01v8 ad=2.2143 pd=13.75 as=2.2143 ps=13.75 w=13.42 l=2.87
X10 B.t5 B.t3 B.t4 w_n4170_n3652# sky130_fd_pr__pfet_01v8 ad=5.2338 pd=27.62 as=0 ps=0 w=13.42 l=2.87
X11 VTAIL.t5 VN.t3 VDD2.t4 w_n4170_n3652# sky130_fd_pr__pfet_01v8 ad=5.2338 pd=27.62 as=2.2143 ps=13.75 w=13.42 l=2.87
X12 VDD2.t3 VN.t4 VTAIL.t2 w_n4170_n3652# sky130_fd_pr__pfet_01v8 ad=2.2143 pd=13.75 as=5.2338 ps=27.62 w=13.42 l=2.87
X13 VDD1.t2 VP.t5 VTAIL.t10 w_n4170_n3652# sky130_fd_pr__pfet_01v8 ad=2.2143 pd=13.75 as=5.2338 ps=27.62 w=13.42 l=2.87
X14 VTAIL.t9 VP.t6 VDD1.t4 w_n4170_n3652# sky130_fd_pr__pfet_01v8 ad=2.2143 pd=13.75 as=2.2143 ps=13.75 w=13.42 l=2.87
X15 VTAIL.t8 VP.t7 VDD1.t7 w_n4170_n3652# sky130_fd_pr__pfet_01v8 ad=5.2338 pd=27.62 as=2.2143 ps=13.75 w=13.42 l=2.87
X16 VTAIL.t4 VN.t5 VDD2.t2 w_n4170_n3652# sky130_fd_pr__pfet_01v8 ad=2.2143 pd=13.75 as=2.2143 ps=13.75 w=13.42 l=2.87
X17 VDD2.t1 VN.t6 VTAIL.t1 w_n4170_n3652# sky130_fd_pr__pfet_01v8 ad=2.2143 pd=13.75 as=2.2143 ps=13.75 w=13.42 l=2.87
X18 B.t2 B.t0 B.t1 w_n4170_n3652# sky130_fd_pr__pfet_01v8 ad=5.2338 pd=27.62 as=0 ps=0 w=13.42 l=2.87
X19 VDD2.t0 VN.t7 VTAIL.t0 w_n4170_n3652# sky130_fd_pr__pfet_01v8 ad=2.2143 pd=13.75 as=5.2338 ps=27.62 w=13.42 l=2.87
R0 VP.n19 VP.n16 161.3
R1 VP.n21 VP.n20 161.3
R2 VP.n22 VP.n15 161.3
R3 VP.n24 VP.n23 161.3
R4 VP.n25 VP.n14 161.3
R5 VP.n28 VP.n27 161.3
R6 VP.n29 VP.n13 161.3
R7 VP.n31 VP.n30 161.3
R8 VP.n32 VP.n12 161.3
R9 VP.n34 VP.n33 161.3
R10 VP.n35 VP.n11 161.3
R11 VP.n37 VP.n36 161.3
R12 VP.n38 VP.n10 161.3
R13 VP.n74 VP.n0 161.3
R14 VP.n73 VP.n72 161.3
R15 VP.n71 VP.n1 161.3
R16 VP.n70 VP.n69 161.3
R17 VP.n68 VP.n2 161.3
R18 VP.n67 VP.n66 161.3
R19 VP.n65 VP.n3 161.3
R20 VP.n64 VP.n63 161.3
R21 VP.n61 VP.n4 161.3
R22 VP.n60 VP.n59 161.3
R23 VP.n58 VP.n5 161.3
R24 VP.n57 VP.n56 161.3
R25 VP.n55 VP.n6 161.3
R26 VP.n53 VP.n52 161.3
R27 VP.n51 VP.n7 161.3
R28 VP.n50 VP.n49 161.3
R29 VP.n48 VP.n8 161.3
R30 VP.n47 VP.n46 161.3
R31 VP.n45 VP.n9 161.3
R32 VP.n44 VP.n43 161.3
R33 VP.n17 VP.t0 145.733
R34 VP.n42 VP.t7 112.692
R35 VP.n54 VP.t3 112.692
R36 VP.n62 VP.t6 112.692
R37 VP.n75 VP.t1 112.692
R38 VP.n39 VP.t5 112.692
R39 VP.n26 VP.t4 112.692
R40 VP.n18 VP.t2 112.692
R41 VP.n42 VP.n41 108.45
R42 VP.n76 VP.n75 108.45
R43 VP.n40 VP.n39 108.45
R44 VP.n18 VP.n17 56.7106
R45 VP.n60 VP.n5 56.5617
R46 VP.n24 VP.n15 56.5617
R47 VP.n41 VP.n40 53.2042
R48 VP.n49 VP.n48 45.4209
R49 VP.n69 VP.n68 45.4209
R50 VP.n33 VP.n32 45.4209
R51 VP.n48 VP.n47 35.7332
R52 VP.n69 VP.n1 35.7332
R53 VP.n33 VP.n11 35.7332
R54 VP.n43 VP.n9 24.5923
R55 VP.n47 VP.n9 24.5923
R56 VP.n49 VP.n7 24.5923
R57 VP.n53 VP.n7 24.5923
R58 VP.n56 VP.n55 24.5923
R59 VP.n56 VP.n5 24.5923
R60 VP.n61 VP.n60 24.5923
R61 VP.n63 VP.n61 24.5923
R62 VP.n67 VP.n3 24.5923
R63 VP.n68 VP.n67 24.5923
R64 VP.n73 VP.n1 24.5923
R65 VP.n74 VP.n73 24.5923
R66 VP.n37 VP.n11 24.5923
R67 VP.n38 VP.n37 24.5923
R68 VP.n25 VP.n24 24.5923
R69 VP.n27 VP.n25 24.5923
R70 VP.n31 VP.n13 24.5923
R71 VP.n32 VP.n31 24.5923
R72 VP.n20 VP.n19 24.5923
R73 VP.n20 VP.n15 24.5923
R74 VP.n55 VP.n54 17.2148
R75 VP.n63 VP.n62 17.2148
R76 VP.n27 VP.n26 17.2148
R77 VP.n19 VP.n18 17.2148
R78 VP.n54 VP.n53 7.37805
R79 VP.n62 VP.n3 7.37805
R80 VP.n26 VP.n13 7.37805
R81 VP.n17 VP.n16 5.07592
R82 VP.n43 VP.n42 2.45968
R83 VP.n75 VP.n74 2.45968
R84 VP.n39 VP.n38 2.45968
R85 VP.n40 VP.n10 0.278335
R86 VP.n44 VP.n41 0.278335
R87 VP.n76 VP.n0 0.278335
R88 VP.n21 VP.n16 0.189894
R89 VP.n22 VP.n21 0.189894
R90 VP.n23 VP.n22 0.189894
R91 VP.n23 VP.n14 0.189894
R92 VP.n28 VP.n14 0.189894
R93 VP.n29 VP.n28 0.189894
R94 VP.n30 VP.n29 0.189894
R95 VP.n30 VP.n12 0.189894
R96 VP.n34 VP.n12 0.189894
R97 VP.n35 VP.n34 0.189894
R98 VP.n36 VP.n35 0.189894
R99 VP.n36 VP.n10 0.189894
R100 VP.n45 VP.n44 0.189894
R101 VP.n46 VP.n45 0.189894
R102 VP.n46 VP.n8 0.189894
R103 VP.n50 VP.n8 0.189894
R104 VP.n51 VP.n50 0.189894
R105 VP.n52 VP.n51 0.189894
R106 VP.n52 VP.n6 0.189894
R107 VP.n57 VP.n6 0.189894
R108 VP.n58 VP.n57 0.189894
R109 VP.n59 VP.n58 0.189894
R110 VP.n59 VP.n4 0.189894
R111 VP.n64 VP.n4 0.189894
R112 VP.n65 VP.n64 0.189894
R113 VP.n66 VP.n65 0.189894
R114 VP.n66 VP.n2 0.189894
R115 VP.n70 VP.n2 0.189894
R116 VP.n71 VP.n70 0.189894
R117 VP.n72 VP.n71 0.189894
R118 VP.n72 VP.n0 0.189894
R119 VP VP.n76 0.153485
R120 VDD1 VDD1.n0 77.6707
R121 VDD1.n3 VDD1.n2 77.557
R122 VDD1.n3 VDD1.n1 77.557
R123 VDD1.n5 VDD1.n4 76.2331
R124 VDD1.n5 VDD1.n3 48.2811
R125 VDD1.n4 VDD1.t1 2.42263
R126 VDD1.n4 VDD1.t2 2.42263
R127 VDD1.n0 VDD1.t3 2.42263
R128 VDD1.n0 VDD1.t6 2.42263
R129 VDD1.n2 VDD1.t4 2.42263
R130 VDD1.n2 VDD1.t5 2.42263
R131 VDD1.n1 VDD1.t7 2.42263
R132 VDD1.n1 VDD1.t0 2.42263
R133 VDD1 VDD1.n5 1.32162
R134 VTAIL.n537 VTAIL.n536 585
R135 VTAIL.n539 VTAIL.n538 585
R136 VTAIL.n532 VTAIL.n531 585
R137 VTAIL.n545 VTAIL.n544 585
R138 VTAIL.n547 VTAIL.n546 585
R139 VTAIL.n528 VTAIL.n527 585
R140 VTAIL.n553 VTAIL.n552 585
R141 VTAIL.n555 VTAIL.n554 585
R142 VTAIL.n524 VTAIL.n523 585
R143 VTAIL.n561 VTAIL.n560 585
R144 VTAIL.n563 VTAIL.n562 585
R145 VTAIL.n520 VTAIL.n519 585
R146 VTAIL.n569 VTAIL.n568 585
R147 VTAIL.n571 VTAIL.n570 585
R148 VTAIL.n516 VTAIL.n515 585
R149 VTAIL.n577 VTAIL.n576 585
R150 VTAIL.n579 VTAIL.n578 585
R151 VTAIL.n27 VTAIL.n26 585
R152 VTAIL.n29 VTAIL.n28 585
R153 VTAIL.n22 VTAIL.n21 585
R154 VTAIL.n35 VTAIL.n34 585
R155 VTAIL.n37 VTAIL.n36 585
R156 VTAIL.n18 VTAIL.n17 585
R157 VTAIL.n43 VTAIL.n42 585
R158 VTAIL.n45 VTAIL.n44 585
R159 VTAIL.n14 VTAIL.n13 585
R160 VTAIL.n51 VTAIL.n50 585
R161 VTAIL.n53 VTAIL.n52 585
R162 VTAIL.n10 VTAIL.n9 585
R163 VTAIL.n59 VTAIL.n58 585
R164 VTAIL.n61 VTAIL.n60 585
R165 VTAIL.n6 VTAIL.n5 585
R166 VTAIL.n67 VTAIL.n66 585
R167 VTAIL.n69 VTAIL.n68 585
R168 VTAIL.n99 VTAIL.n98 585
R169 VTAIL.n101 VTAIL.n100 585
R170 VTAIL.n94 VTAIL.n93 585
R171 VTAIL.n107 VTAIL.n106 585
R172 VTAIL.n109 VTAIL.n108 585
R173 VTAIL.n90 VTAIL.n89 585
R174 VTAIL.n115 VTAIL.n114 585
R175 VTAIL.n117 VTAIL.n116 585
R176 VTAIL.n86 VTAIL.n85 585
R177 VTAIL.n123 VTAIL.n122 585
R178 VTAIL.n125 VTAIL.n124 585
R179 VTAIL.n82 VTAIL.n81 585
R180 VTAIL.n131 VTAIL.n130 585
R181 VTAIL.n133 VTAIL.n132 585
R182 VTAIL.n78 VTAIL.n77 585
R183 VTAIL.n139 VTAIL.n138 585
R184 VTAIL.n141 VTAIL.n140 585
R185 VTAIL.n173 VTAIL.n172 585
R186 VTAIL.n175 VTAIL.n174 585
R187 VTAIL.n168 VTAIL.n167 585
R188 VTAIL.n181 VTAIL.n180 585
R189 VTAIL.n183 VTAIL.n182 585
R190 VTAIL.n164 VTAIL.n163 585
R191 VTAIL.n189 VTAIL.n188 585
R192 VTAIL.n191 VTAIL.n190 585
R193 VTAIL.n160 VTAIL.n159 585
R194 VTAIL.n197 VTAIL.n196 585
R195 VTAIL.n199 VTAIL.n198 585
R196 VTAIL.n156 VTAIL.n155 585
R197 VTAIL.n205 VTAIL.n204 585
R198 VTAIL.n207 VTAIL.n206 585
R199 VTAIL.n152 VTAIL.n151 585
R200 VTAIL.n213 VTAIL.n212 585
R201 VTAIL.n215 VTAIL.n214 585
R202 VTAIL.n507 VTAIL.n506 585
R203 VTAIL.n505 VTAIL.n504 585
R204 VTAIL.n444 VTAIL.n443 585
R205 VTAIL.n499 VTAIL.n498 585
R206 VTAIL.n497 VTAIL.n496 585
R207 VTAIL.n448 VTAIL.n447 585
R208 VTAIL.n491 VTAIL.n490 585
R209 VTAIL.n489 VTAIL.n488 585
R210 VTAIL.n452 VTAIL.n451 585
R211 VTAIL.n483 VTAIL.n482 585
R212 VTAIL.n481 VTAIL.n480 585
R213 VTAIL.n456 VTAIL.n455 585
R214 VTAIL.n475 VTAIL.n474 585
R215 VTAIL.n473 VTAIL.n472 585
R216 VTAIL.n460 VTAIL.n459 585
R217 VTAIL.n467 VTAIL.n466 585
R218 VTAIL.n465 VTAIL.n464 585
R219 VTAIL.n433 VTAIL.n432 585
R220 VTAIL.n431 VTAIL.n430 585
R221 VTAIL.n370 VTAIL.n369 585
R222 VTAIL.n425 VTAIL.n424 585
R223 VTAIL.n423 VTAIL.n422 585
R224 VTAIL.n374 VTAIL.n373 585
R225 VTAIL.n417 VTAIL.n416 585
R226 VTAIL.n415 VTAIL.n414 585
R227 VTAIL.n378 VTAIL.n377 585
R228 VTAIL.n409 VTAIL.n408 585
R229 VTAIL.n407 VTAIL.n406 585
R230 VTAIL.n382 VTAIL.n381 585
R231 VTAIL.n401 VTAIL.n400 585
R232 VTAIL.n399 VTAIL.n398 585
R233 VTAIL.n386 VTAIL.n385 585
R234 VTAIL.n393 VTAIL.n392 585
R235 VTAIL.n391 VTAIL.n390 585
R236 VTAIL.n361 VTAIL.n360 585
R237 VTAIL.n359 VTAIL.n358 585
R238 VTAIL.n298 VTAIL.n297 585
R239 VTAIL.n353 VTAIL.n352 585
R240 VTAIL.n351 VTAIL.n350 585
R241 VTAIL.n302 VTAIL.n301 585
R242 VTAIL.n345 VTAIL.n344 585
R243 VTAIL.n343 VTAIL.n342 585
R244 VTAIL.n306 VTAIL.n305 585
R245 VTAIL.n337 VTAIL.n336 585
R246 VTAIL.n335 VTAIL.n334 585
R247 VTAIL.n310 VTAIL.n309 585
R248 VTAIL.n329 VTAIL.n328 585
R249 VTAIL.n327 VTAIL.n326 585
R250 VTAIL.n314 VTAIL.n313 585
R251 VTAIL.n321 VTAIL.n320 585
R252 VTAIL.n319 VTAIL.n318 585
R253 VTAIL.n287 VTAIL.n286 585
R254 VTAIL.n285 VTAIL.n284 585
R255 VTAIL.n224 VTAIL.n223 585
R256 VTAIL.n279 VTAIL.n278 585
R257 VTAIL.n277 VTAIL.n276 585
R258 VTAIL.n228 VTAIL.n227 585
R259 VTAIL.n271 VTAIL.n270 585
R260 VTAIL.n269 VTAIL.n268 585
R261 VTAIL.n232 VTAIL.n231 585
R262 VTAIL.n263 VTAIL.n262 585
R263 VTAIL.n261 VTAIL.n260 585
R264 VTAIL.n236 VTAIL.n235 585
R265 VTAIL.n255 VTAIL.n254 585
R266 VTAIL.n253 VTAIL.n252 585
R267 VTAIL.n240 VTAIL.n239 585
R268 VTAIL.n247 VTAIL.n246 585
R269 VTAIL.n245 VTAIL.n244 585
R270 VTAIL.n578 VTAIL.n512 498.474
R271 VTAIL.n68 VTAIL.n2 498.474
R272 VTAIL.n140 VTAIL.n74 498.474
R273 VTAIL.n214 VTAIL.n148 498.474
R274 VTAIL.n506 VTAIL.n440 498.474
R275 VTAIL.n432 VTAIL.n366 498.474
R276 VTAIL.n360 VTAIL.n294 498.474
R277 VTAIL.n286 VTAIL.n220 498.474
R278 VTAIL.n535 VTAIL.t0 327.466
R279 VTAIL.n25 VTAIL.t5 327.466
R280 VTAIL.n97 VTAIL.t14 327.466
R281 VTAIL.n171 VTAIL.t8 327.466
R282 VTAIL.n463 VTAIL.t10 327.466
R283 VTAIL.n389 VTAIL.t15 327.466
R284 VTAIL.n317 VTAIL.t2 327.466
R285 VTAIL.n243 VTAIL.t3 327.466
R286 VTAIL.n538 VTAIL.n537 171.744
R287 VTAIL.n538 VTAIL.n531 171.744
R288 VTAIL.n545 VTAIL.n531 171.744
R289 VTAIL.n546 VTAIL.n545 171.744
R290 VTAIL.n546 VTAIL.n527 171.744
R291 VTAIL.n553 VTAIL.n527 171.744
R292 VTAIL.n554 VTAIL.n553 171.744
R293 VTAIL.n554 VTAIL.n523 171.744
R294 VTAIL.n561 VTAIL.n523 171.744
R295 VTAIL.n562 VTAIL.n561 171.744
R296 VTAIL.n562 VTAIL.n519 171.744
R297 VTAIL.n569 VTAIL.n519 171.744
R298 VTAIL.n570 VTAIL.n569 171.744
R299 VTAIL.n570 VTAIL.n515 171.744
R300 VTAIL.n577 VTAIL.n515 171.744
R301 VTAIL.n578 VTAIL.n577 171.744
R302 VTAIL.n28 VTAIL.n27 171.744
R303 VTAIL.n28 VTAIL.n21 171.744
R304 VTAIL.n35 VTAIL.n21 171.744
R305 VTAIL.n36 VTAIL.n35 171.744
R306 VTAIL.n36 VTAIL.n17 171.744
R307 VTAIL.n43 VTAIL.n17 171.744
R308 VTAIL.n44 VTAIL.n43 171.744
R309 VTAIL.n44 VTAIL.n13 171.744
R310 VTAIL.n51 VTAIL.n13 171.744
R311 VTAIL.n52 VTAIL.n51 171.744
R312 VTAIL.n52 VTAIL.n9 171.744
R313 VTAIL.n59 VTAIL.n9 171.744
R314 VTAIL.n60 VTAIL.n59 171.744
R315 VTAIL.n60 VTAIL.n5 171.744
R316 VTAIL.n67 VTAIL.n5 171.744
R317 VTAIL.n68 VTAIL.n67 171.744
R318 VTAIL.n100 VTAIL.n99 171.744
R319 VTAIL.n100 VTAIL.n93 171.744
R320 VTAIL.n107 VTAIL.n93 171.744
R321 VTAIL.n108 VTAIL.n107 171.744
R322 VTAIL.n108 VTAIL.n89 171.744
R323 VTAIL.n115 VTAIL.n89 171.744
R324 VTAIL.n116 VTAIL.n115 171.744
R325 VTAIL.n116 VTAIL.n85 171.744
R326 VTAIL.n123 VTAIL.n85 171.744
R327 VTAIL.n124 VTAIL.n123 171.744
R328 VTAIL.n124 VTAIL.n81 171.744
R329 VTAIL.n131 VTAIL.n81 171.744
R330 VTAIL.n132 VTAIL.n131 171.744
R331 VTAIL.n132 VTAIL.n77 171.744
R332 VTAIL.n139 VTAIL.n77 171.744
R333 VTAIL.n140 VTAIL.n139 171.744
R334 VTAIL.n174 VTAIL.n173 171.744
R335 VTAIL.n174 VTAIL.n167 171.744
R336 VTAIL.n181 VTAIL.n167 171.744
R337 VTAIL.n182 VTAIL.n181 171.744
R338 VTAIL.n182 VTAIL.n163 171.744
R339 VTAIL.n189 VTAIL.n163 171.744
R340 VTAIL.n190 VTAIL.n189 171.744
R341 VTAIL.n190 VTAIL.n159 171.744
R342 VTAIL.n197 VTAIL.n159 171.744
R343 VTAIL.n198 VTAIL.n197 171.744
R344 VTAIL.n198 VTAIL.n155 171.744
R345 VTAIL.n205 VTAIL.n155 171.744
R346 VTAIL.n206 VTAIL.n205 171.744
R347 VTAIL.n206 VTAIL.n151 171.744
R348 VTAIL.n213 VTAIL.n151 171.744
R349 VTAIL.n214 VTAIL.n213 171.744
R350 VTAIL.n506 VTAIL.n505 171.744
R351 VTAIL.n505 VTAIL.n443 171.744
R352 VTAIL.n498 VTAIL.n443 171.744
R353 VTAIL.n498 VTAIL.n497 171.744
R354 VTAIL.n497 VTAIL.n447 171.744
R355 VTAIL.n490 VTAIL.n447 171.744
R356 VTAIL.n490 VTAIL.n489 171.744
R357 VTAIL.n489 VTAIL.n451 171.744
R358 VTAIL.n482 VTAIL.n451 171.744
R359 VTAIL.n482 VTAIL.n481 171.744
R360 VTAIL.n481 VTAIL.n455 171.744
R361 VTAIL.n474 VTAIL.n455 171.744
R362 VTAIL.n474 VTAIL.n473 171.744
R363 VTAIL.n473 VTAIL.n459 171.744
R364 VTAIL.n466 VTAIL.n459 171.744
R365 VTAIL.n466 VTAIL.n465 171.744
R366 VTAIL.n432 VTAIL.n431 171.744
R367 VTAIL.n431 VTAIL.n369 171.744
R368 VTAIL.n424 VTAIL.n369 171.744
R369 VTAIL.n424 VTAIL.n423 171.744
R370 VTAIL.n423 VTAIL.n373 171.744
R371 VTAIL.n416 VTAIL.n373 171.744
R372 VTAIL.n416 VTAIL.n415 171.744
R373 VTAIL.n415 VTAIL.n377 171.744
R374 VTAIL.n408 VTAIL.n377 171.744
R375 VTAIL.n408 VTAIL.n407 171.744
R376 VTAIL.n407 VTAIL.n381 171.744
R377 VTAIL.n400 VTAIL.n381 171.744
R378 VTAIL.n400 VTAIL.n399 171.744
R379 VTAIL.n399 VTAIL.n385 171.744
R380 VTAIL.n392 VTAIL.n385 171.744
R381 VTAIL.n392 VTAIL.n391 171.744
R382 VTAIL.n360 VTAIL.n359 171.744
R383 VTAIL.n359 VTAIL.n297 171.744
R384 VTAIL.n352 VTAIL.n297 171.744
R385 VTAIL.n352 VTAIL.n351 171.744
R386 VTAIL.n351 VTAIL.n301 171.744
R387 VTAIL.n344 VTAIL.n301 171.744
R388 VTAIL.n344 VTAIL.n343 171.744
R389 VTAIL.n343 VTAIL.n305 171.744
R390 VTAIL.n336 VTAIL.n305 171.744
R391 VTAIL.n336 VTAIL.n335 171.744
R392 VTAIL.n335 VTAIL.n309 171.744
R393 VTAIL.n328 VTAIL.n309 171.744
R394 VTAIL.n328 VTAIL.n327 171.744
R395 VTAIL.n327 VTAIL.n313 171.744
R396 VTAIL.n320 VTAIL.n313 171.744
R397 VTAIL.n320 VTAIL.n319 171.744
R398 VTAIL.n286 VTAIL.n285 171.744
R399 VTAIL.n285 VTAIL.n223 171.744
R400 VTAIL.n278 VTAIL.n223 171.744
R401 VTAIL.n278 VTAIL.n277 171.744
R402 VTAIL.n277 VTAIL.n227 171.744
R403 VTAIL.n270 VTAIL.n227 171.744
R404 VTAIL.n270 VTAIL.n269 171.744
R405 VTAIL.n269 VTAIL.n231 171.744
R406 VTAIL.n262 VTAIL.n231 171.744
R407 VTAIL.n262 VTAIL.n261 171.744
R408 VTAIL.n261 VTAIL.n235 171.744
R409 VTAIL.n254 VTAIL.n235 171.744
R410 VTAIL.n254 VTAIL.n253 171.744
R411 VTAIL.n253 VTAIL.n239 171.744
R412 VTAIL.n246 VTAIL.n239 171.744
R413 VTAIL.n246 VTAIL.n245 171.744
R414 VTAIL.n537 VTAIL.t0 85.8723
R415 VTAIL.n27 VTAIL.t5 85.8723
R416 VTAIL.n99 VTAIL.t14 85.8723
R417 VTAIL.n173 VTAIL.t8 85.8723
R418 VTAIL.n465 VTAIL.t10 85.8723
R419 VTAIL.n391 VTAIL.t15 85.8723
R420 VTAIL.n319 VTAIL.t2 85.8723
R421 VTAIL.n245 VTAIL.t3 85.8723
R422 VTAIL.n439 VTAIL.n438 59.5544
R423 VTAIL.n293 VTAIL.n292 59.5544
R424 VTAIL.n1 VTAIL.n0 59.5543
R425 VTAIL.n147 VTAIL.n146 59.5543
R426 VTAIL.n583 VTAIL.n582 36.452
R427 VTAIL.n73 VTAIL.n72 36.452
R428 VTAIL.n145 VTAIL.n144 36.452
R429 VTAIL.n219 VTAIL.n218 36.452
R430 VTAIL.n511 VTAIL.n510 36.452
R431 VTAIL.n437 VTAIL.n436 36.452
R432 VTAIL.n365 VTAIL.n364 36.452
R433 VTAIL.n291 VTAIL.n290 36.452
R434 VTAIL.n583 VTAIL.n511 26.6945
R435 VTAIL.n291 VTAIL.n219 26.6945
R436 VTAIL.n536 VTAIL.n535 16.3895
R437 VTAIL.n26 VTAIL.n25 16.3895
R438 VTAIL.n98 VTAIL.n97 16.3895
R439 VTAIL.n172 VTAIL.n171 16.3895
R440 VTAIL.n464 VTAIL.n463 16.3895
R441 VTAIL.n390 VTAIL.n389 16.3895
R442 VTAIL.n318 VTAIL.n317 16.3895
R443 VTAIL.n244 VTAIL.n243 16.3895
R444 VTAIL.n539 VTAIL.n534 12.8005
R445 VTAIL.n580 VTAIL.n579 12.8005
R446 VTAIL.n29 VTAIL.n24 12.8005
R447 VTAIL.n70 VTAIL.n69 12.8005
R448 VTAIL.n101 VTAIL.n96 12.8005
R449 VTAIL.n142 VTAIL.n141 12.8005
R450 VTAIL.n175 VTAIL.n170 12.8005
R451 VTAIL.n216 VTAIL.n215 12.8005
R452 VTAIL.n508 VTAIL.n507 12.8005
R453 VTAIL.n467 VTAIL.n462 12.8005
R454 VTAIL.n434 VTAIL.n433 12.8005
R455 VTAIL.n393 VTAIL.n388 12.8005
R456 VTAIL.n362 VTAIL.n361 12.8005
R457 VTAIL.n321 VTAIL.n316 12.8005
R458 VTAIL.n288 VTAIL.n287 12.8005
R459 VTAIL.n247 VTAIL.n242 12.8005
R460 VTAIL.n540 VTAIL.n532 12.0247
R461 VTAIL.n576 VTAIL.n514 12.0247
R462 VTAIL.n30 VTAIL.n22 12.0247
R463 VTAIL.n66 VTAIL.n4 12.0247
R464 VTAIL.n102 VTAIL.n94 12.0247
R465 VTAIL.n138 VTAIL.n76 12.0247
R466 VTAIL.n176 VTAIL.n168 12.0247
R467 VTAIL.n212 VTAIL.n150 12.0247
R468 VTAIL.n504 VTAIL.n442 12.0247
R469 VTAIL.n468 VTAIL.n460 12.0247
R470 VTAIL.n430 VTAIL.n368 12.0247
R471 VTAIL.n394 VTAIL.n386 12.0247
R472 VTAIL.n358 VTAIL.n296 12.0247
R473 VTAIL.n322 VTAIL.n314 12.0247
R474 VTAIL.n284 VTAIL.n222 12.0247
R475 VTAIL.n248 VTAIL.n240 12.0247
R476 VTAIL.n544 VTAIL.n543 11.249
R477 VTAIL.n575 VTAIL.n516 11.249
R478 VTAIL.n34 VTAIL.n33 11.249
R479 VTAIL.n65 VTAIL.n6 11.249
R480 VTAIL.n106 VTAIL.n105 11.249
R481 VTAIL.n137 VTAIL.n78 11.249
R482 VTAIL.n180 VTAIL.n179 11.249
R483 VTAIL.n211 VTAIL.n152 11.249
R484 VTAIL.n503 VTAIL.n444 11.249
R485 VTAIL.n472 VTAIL.n471 11.249
R486 VTAIL.n429 VTAIL.n370 11.249
R487 VTAIL.n398 VTAIL.n397 11.249
R488 VTAIL.n357 VTAIL.n298 11.249
R489 VTAIL.n326 VTAIL.n325 11.249
R490 VTAIL.n283 VTAIL.n224 11.249
R491 VTAIL.n252 VTAIL.n251 11.249
R492 VTAIL.n547 VTAIL.n530 10.4732
R493 VTAIL.n572 VTAIL.n571 10.4732
R494 VTAIL.n37 VTAIL.n20 10.4732
R495 VTAIL.n62 VTAIL.n61 10.4732
R496 VTAIL.n109 VTAIL.n92 10.4732
R497 VTAIL.n134 VTAIL.n133 10.4732
R498 VTAIL.n183 VTAIL.n166 10.4732
R499 VTAIL.n208 VTAIL.n207 10.4732
R500 VTAIL.n500 VTAIL.n499 10.4732
R501 VTAIL.n475 VTAIL.n458 10.4732
R502 VTAIL.n426 VTAIL.n425 10.4732
R503 VTAIL.n401 VTAIL.n384 10.4732
R504 VTAIL.n354 VTAIL.n353 10.4732
R505 VTAIL.n329 VTAIL.n312 10.4732
R506 VTAIL.n280 VTAIL.n279 10.4732
R507 VTAIL.n255 VTAIL.n238 10.4732
R508 VTAIL.n548 VTAIL.n528 9.69747
R509 VTAIL.n568 VTAIL.n518 9.69747
R510 VTAIL.n38 VTAIL.n18 9.69747
R511 VTAIL.n58 VTAIL.n8 9.69747
R512 VTAIL.n110 VTAIL.n90 9.69747
R513 VTAIL.n130 VTAIL.n80 9.69747
R514 VTAIL.n184 VTAIL.n164 9.69747
R515 VTAIL.n204 VTAIL.n154 9.69747
R516 VTAIL.n496 VTAIL.n446 9.69747
R517 VTAIL.n476 VTAIL.n456 9.69747
R518 VTAIL.n422 VTAIL.n372 9.69747
R519 VTAIL.n402 VTAIL.n382 9.69747
R520 VTAIL.n350 VTAIL.n300 9.69747
R521 VTAIL.n330 VTAIL.n310 9.69747
R522 VTAIL.n276 VTAIL.n226 9.69747
R523 VTAIL.n256 VTAIL.n236 9.69747
R524 VTAIL.n582 VTAIL.n581 9.45567
R525 VTAIL.n72 VTAIL.n71 9.45567
R526 VTAIL.n144 VTAIL.n143 9.45567
R527 VTAIL.n218 VTAIL.n217 9.45567
R528 VTAIL.n510 VTAIL.n509 9.45567
R529 VTAIL.n436 VTAIL.n435 9.45567
R530 VTAIL.n364 VTAIL.n363 9.45567
R531 VTAIL.n290 VTAIL.n289 9.45567
R532 VTAIL.n557 VTAIL.n556 9.3005
R533 VTAIL.n526 VTAIL.n525 9.3005
R534 VTAIL.n551 VTAIL.n550 9.3005
R535 VTAIL.n549 VTAIL.n548 9.3005
R536 VTAIL.n530 VTAIL.n529 9.3005
R537 VTAIL.n543 VTAIL.n542 9.3005
R538 VTAIL.n541 VTAIL.n540 9.3005
R539 VTAIL.n534 VTAIL.n533 9.3005
R540 VTAIL.n559 VTAIL.n558 9.3005
R541 VTAIL.n522 VTAIL.n521 9.3005
R542 VTAIL.n565 VTAIL.n564 9.3005
R543 VTAIL.n567 VTAIL.n566 9.3005
R544 VTAIL.n518 VTAIL.n517 9.3005
R545 VTAIL.n573 VTAIL.n572 9.3005
R546 VTAIL.n575 VTAIL.n574 9.3005
R547 VTAIL.n514 VTAIL.n513 9.3005
R548 VTAIL.n581 VTAIL.n580 9.3005
R549 VTAIL.n47 VTAIL.n46 9.3005
R550 VTAIL.n16 VTAIL.n15 9.3005
R551 VTAIL.n41 VTAIL.n40 9.3005
R552 VTAIL.n39 VTAIL.n38 9.3005
R553 VTAIL.n20 VTAIL.n19 9.3005
R554 VTAIL.n33 VTAIL.n32 9.3005
R555 VTAIL.n31 VTAIL.n30 9.3005
R556 VTAIL.n24 VTAIL.n23 9.3005
R557 VTAIL.n49 VTAIL.n48 9.3005
R558 VTAIL.n12 VTAIL.n11 9.3005
R559 VTAIL.n55 VTAIL.n54 9.3005
R560 VTAIL.n57 VTAIL.n56 9.3005
R561 VTAIL.n8 VTAIL.n7 9.3005
R562 VTAIL.n63 VTAIL.n62 9.3005
R563 VTAIL.n65 VTAIL.n64 9.3005
R564 VTAIL.n4 VTAIL.n3 9.3005
R565 VTAIL.n71 VTAIL.n70 9.3005
R566 VTAIL.n119 VTAIL.n118 9.3005
R567 VTAIL.n88 VTAIL.n87 9.3005
R568 VTAIL.n113 VTAIL.n112 9.3005
R569 VTAIL.n111 VTAIL.n110 9.3005
R570 VTAIL.n92 VTAIL.n91 9.3005
R571 VTAIL.n105 VTAIL.n104 9.3005
R572 VTAIL.n103 VTAIL.n102 9.3005
R573 VTAIL.n96 VTAIL.n95 9.3005
R574 VTAIL.n121 VTAIL.n120 9.3005
R575 VTAIL.n84 VTAIL.n83 9.3005
R576 VTAIL.n127 VTAIL.n126 9.3005
R577 VTAIL.n129 VTAIL.n128 9.3005
R578 VTAIL.n80 VTAIL.n79 9.3005
R579 VTAIL.n135 VTAIL.n134 9.3005
R580 VTAIL.n137 VTAIL.n136 9.3005
R581 VTAIL.n76 VTAIL.n75 9.3005
R582 VTAIL.n143 VTAIL.n142 9.3005
R583 VTAIL.n193 VTAIL.n192 9.3005
R584 VTAIL.n162 VTAIL.n161 9.3005
R585 VTAIL.n187 VTAIL.n186 9.3005
R586 VTAIL.n185 VTAIL.n184 9.3005
R587 VTAIL.n166 VTAIL.n165 9.3005
R588 VTAIL.n179 VTAIL.n178 9.3005
R589 VTAIL.n177 VTAIL.n176 9.3005
R590 VTAIL.n170 VTAIL.n169 9.3005
R591 VTAIL.n195 VTAIL.n194 9.3005
R592 VTAIL.n158 VTAIL.n157 9.3005
R593 VTAIL.n201 VTAIL.n200 9.3005
R594 VTAIL.n203 VTAIL.n202 9.3005
R595 VTAIL.n154 VTAIL.n153 9.3005
R596 VTAIL.n209 VTAIL.n208 9.3005
R597 VTAIL.n211 VTAIL.n210 9.3005
R598 VTAIL.n150 VTAIL.n149 9.3005
R599 VTAIL.n217 VTAIL.n216 9.3005
R600 VTAIL.n450 VTAIL.n449 9.3005
R601 VTAIL.n493 VTAIL.n492 9.3005
R602 VTAIL.n495 VTAIL.n494 9.3005
R603 VTAIL.n446 VTAIL.n445 9.3005
R604 VTAIL.n501 VTAIL.n500 9.3005
R605 VTAIL.n503 VTAIL.n502 9.3005
R606 VTAIL.n442 VTAIL.n441 9.3005
R607 VTAIL.n509 VTAIL.n508 9.3005
R608 VTAIL.n487 VTAIL.n486 9.3005
R609 VTAIL.n485 VTAIL.n484 9.3005
R610 VTAIL.n454 VTAIL.n453 9.3005
R611 VTAIL.n479 VTAIL.n478 9.3005
R612 VTAIL.n477 VTAIL.n476 9.3005
R613 VTAIL.n458 VTAIL.n457 9.3005
R614 VTAIL.n471 VTAIL.n470 9.3005
R615 VTAIL.n469 VTAIL.n468 9.3005
R616 VTAIL.n462 VTAIL.n461 9.3005
R617 VTAIL.n376 VTAIL.n375 9.3005
R618 VTAIL.n419 VTAIL.n418 9.3005
R619 VTAIL.n421 VTAIL.n420 9.3005
R620 VTAIL.n372 VTAIL.n371 9.3005
R621 VTAIL.n427 VTAIL.n426 9.3005
R622 VTAIL.n429 VTAIL.n428 9.3005
R623 VTAIL.n368 VTAIL.n367 9.3005
R624 VTAIL.n435 VTAIL.n434 9.3005
R625 VTAIL.n413 VTAIL.n412 9.3005
R626 VTAIL.n411 VTAIL.n410 9.3005
R627 VTAIL.n380 VTAIL.n379 9.3005
R628 VTAIL.n405 VTAIL.n404 9.3005
R629 VTAIL.n403 VTAIL.n402 9.3005
R630 VTAIL.n384 VTAIL.n383 9.3005
R631 VTAIL.n397 VTAIL.n396 9.3005
R632 VTAIL.n395 VTAIL.n394 9.3005
R633 VTAIL.n388 VTAIL.n387 9.3005
R634 VTAIL.n304 VTAIL.n303 9.3005
R635 VTAIL.n347 VTAIL.n346 9.3005
R636 VTAIL.n349 VTAIL.n348 9.3005
R637 VTAIL.n300 VTAIL.n299 9.3005
R638 VTAIL.n355 VTAIL.n354 9.3005
R639 VTAIL.n357 VTAIL.n356 9.3005
R640 VTAIL.n296 VTAIL.n295 9.3005
R641 VTAIL.n363 VTAIL.n362 9.3005
R642 VTAIL.n341 VTAIL.n340 9.3005
R643 VTAIL.n339 VTAIL.n338 9.3005
R644 VTAIL.n308 VTAIL.n307 9.3005
R645 VTAIL.n333 VTAIL.n332 9.3005
R646 VTAIL.n331 VTAIL.n330 9.3005
R647 VTAIL.n312 VTAIL.n311 9.3005
R648 VTAIL.n325 VTAIL.n324 9.3005
R649 VTAIL.n323 VTAIL.n322 9.3005
R650 VTAIL.n316 VTAIL.n315 9.3005
R651 VTAIL.n230 VTAIL.n229 9.3005
R652 VTAIL.n273 VTAIL.n272 9.3005
R653 VTAIL.n275 VTAIL.n274 9.3005
R654 VTAIL.n226 VTAIL.n225 9.3005
R655 VTAIL.n281 VTAIL.n280 9.3005
R656 VTAIL.n283 VTAIL.n282 9.3005
R657 VTAIL.n222 VTAIL.n221 9.3005
R658 VTAIL.n289 VTAIL.n288 9.3005
R659 VTAIL.n267 VTAIL.n266 9.3005
R660 VTAIL.n265 VTAIL.n264 9.3005
R661 VTAIL.n234 VTAIL.n233 9.3005
R662 VTAIL.n259 VTAIL.n258 9.3005
R663 VTAIL.n257 VTAIL.n256 9.3005
R664 VTAIL.n238 VTAIL.n237 9.3005
R665 VTAIL.n251 VTAIL.n250 9.3005
R666 VTAIL.n249 VTAIL.n248 9.3005
R667 VTAIL.n242 VTAIL.n241 9.3005
R668 VTAIL.n552 VTAIL.n551 8.92171
R669 VTAIL.n567 VTAIL.n520 8.92171
R670 VTAIL.n42 VTAIL.n41 8.92171
R671 VTAIL.n57 VTAIL.n10 8.92171
R672 VTAIL.n114 VTAIL.n113 8.92171
R673 VTAIL.n129 VTAIL.n82 8.92171
R674 VTAIL.n188 VTAIL.n187 8.92171
R675 VTAIL.n203 VTAIL.n156 8.92171
R676 VTAIL.n495 VTAIL.n448 8.92171
R677 VTAIL.n480 VTAIL.n479 8.92171
R678 VTAIL.n421 VTAIL.n374 8.92171
R679 VTAIL.n406 VTAIL.n405 8.92171
R680 VTAIL.n349 VTAIL.n302 8.92171
R681 VTAIL.n334 VTAIL.n333 8.92171
R682 VTAIL.n275 VTAIL.n228 8.92171
R683 VTAIL.n260 VTAIL.n259 8.92171
R684 VTAIL.n555 VTAIL.n526 8.14595
R685 VTAIL.n564 VTAIL.n563 8.14595
R686 VTAIL.n45 VTAIL.n16 8.14595
R687 VTAIL.n54 VTAIL.n53 8.14595
R688 VTAIL.n117 VTAIL.n88 8.14595
R689 VTAIL.n126 VTAIL.n125 8.14595
R690 VTAIL.n191 VTAIL.n162 8.14595
R691 VTAIL.n200 VTAIL.n199 8.14595
R692 VTAIL.n492 VTAIL.n491 8.14595
R693 VTAIL.n483 VTAIL.n454 8.14595
R694 VTAIL.n418 VTAIL.n417 8.14595
R695 VTAIL.n409 VTAIL.n380 8.14595
R696 VTAIL.n346 VTAIL.n345 8.14595
R697 VTAIL.n337 VTAIL.n308 8.14595
R698 VTAIL.n272 VTAIL.n271 8.14595
R699 VTAIL.n263 VTAIL.n234 8.14595
R700 VTAIL.n582 VTAIL.n512 7.75445
R701 VTAIL.n72 VTAIL.n2 7.75445
R702 VTAIL.n144 VTAIL.n74 7.75445
R703 VTAIL.n218 VTAIL.n148 7.75445
R704 VTAIL.n510 VTAIL.n440 7.75445
R705 VTAIL.n436 VTAIL.n366 7.75445
R706 VTAIL.n364 VTAIL.n294 7.75445
R707 VTAIL.n290 VTAIL.n220 7.75445
R708 VTAIL.n556 VTAIL.n524 7.3702
R709 VTAIL.n560 VTAIL.n522 7.3702
R710 VTAIL.n46 VTAIL.n14 7.3702
R711 VTAIL.n50 VTAIL.n12 7.3702
R712 VTAIL.n118 VTAIL.n86 7.3702
R713 VTAIL.n122 VTAIL.n84 7.3702
R714 VTAIL.n192 VTAIL.n160 7.3702
R715 VTAIL.n196 VTAIL.n158 7.3702
R716 VTAIL.n488 VTAIL.n450 7.3702
R717 VTAIL.n484 VTAIL.n452 7.3702
R718 VTAIL.n414 VTAIL.n376 7.3702
R719 VTAIL.n410 VTAIL.n378 7.3702
R720 VTAIL.n342 VTAIL.n304 7.3702
R721 VTAIL.n338 VTAIL.n306 7.3702
R722 VTAIL.n268 VTAIL.n230 7.3702
R723 VTAIL.n264 VTAIL.n232 7.3702
R724 VTAIL.n559 VTAIL.n524 6.59444
R725 VTAIL.n560 VTAIL.n559 6.59444
R726 VTAIL.n49 VTAIL.n14 6.59444
R727 VTAIL.n50 VTAIL.n49 6.59444
R728 VTAIL.n121 VTAIL.n86 6.59444
R729 VTAIL.n122 VTAIL.n121 6.59444
R730 VTAIL.n195 VTAIL.n160 6.59444
R731 VTAIL.n196 VTAIL.n195 6.59444
R732 VTAIL.n488 VTAIL.n487 6.59444
R733 VTAIL.n487 VTAIL.n452 6.59444
R734 VTAIL.n414 VTAIL.n413 6.59444
R735 VTAIL.n413 VTAIL.n378 6.59444
R736 VTAIL.n342 VTAIL.n341 6.59444
R737 VTAIL.n341 VTAIL.n306 6.59444
R738 VTAIL.n268 VTAIL.n267 6.59444
R739 VTAIL.n267 VTAIL.n232 6.59444
R740 VTAIL.n580 VTAIL.n512 6.08283
R741 VTAIL.n70 VTAIL.n2 6.08283
R742 VTAIL.n142 VTAIL.n74 6.08283
R743 VTAIL.n216 VTAIL.n148 6.08283
R744 VTAIL.n508 VTAIL.n440 6.08283
R745 VTAIL.n434 VTAIL.n366 6.08283
R746 VTAIL.n362 VTAIL.n294 6.08283
R747 VTAIL.n288 VTAIL.n220 6.08283
R748 VTAIL.n556 VTAIL.n555 5.81868
R749 VTAIL.n563 VTAIL.n522 5.81868
R750 VTAIL.n46 VTAIL.n45 5.81868
R751 VTAIL.n53 VTAIL.n12 5.81868
R752 VTAIL.n118 VTAIL.n117 5.81868
R753 VTAIL.n125 VTAIL.n84 5.81868
R754 VTAIL.n192 VTAIL.n191 5.81868
R755 VTAIL.n199 VTAIL.n158 5.81868
R756 VTAIL.n491 VTAIL.n450 5.81868
R757 VTAIL.n484 VTAIL.n483 5.81868
R758 VTAIL.n417 VTAIL.n376 5.81868
R759 VTAIL.n410 VTAIL.n409 5.81868
R760 VTAIL.n345 VTAIL.n304 5.81868
R761 VTAIL.n338 VTAIL.n337 5.81868
R762 VTAIL.n271 VTAIL.n230 5.81868
R763 VTAIL.n264 VTAIL.n263 5.81868
R764 VTAIL.n552 VTAIL.n526 5.04292
R765 VTAIL.n564 VTAIL.n520 5.04292
R766 VTAIL.n42 VTAIL.n16 5.04292
R767 VTAIL.n54 VTAIL.n10 5.04292
R768 VTAIL.n114 VTAIL.n88 5.04292
R769 VTAIL.n126 VTAIL.n82 5.04292
R770 VTAIL.n188 VTAIL.n162 5.04292
R771 VTAIL.n200 VTAIL.n156 5.04292
R772 VTAIL.n492 VTAIL.n448 5.04292
R773 VTAIL.n480 VTAIL.n454 5.04292
R774 VTAIL.n418 VTAIL.n374 5.04292
R775 VTAIL.n406 VTAIL.n380 5.04292
R776 VTAIL.n346 VTAIL.n302 5.04292
R777 VTAIL.n334 VTAIL.n308 5.04292
R778 VTAIL.n272 VTAIL.n228 5.04292
R779 VTAIL.n260 VTAIL.n234 5.04292
R780 VTAIL.n551 VTAIL.n528 4.26717
R781 VTAIL.n568 VTAIL.n567 4.26717
R782 VTAIL.n41 VTAIL.n18 4.26717
R783 VTAIL.n58 VTAIL.n57 4.26717
R784 VTAIL.n113 VTAIL.n90 4.26717
R785 VTAIL.n130 VTAIL.n129 4.26717
R786 VTAIL.n187 VTAIL.n164 4.26717
R787 VTAIL.n204 VTAIL.n203 4.26717
R788 VTAIL.n496 VTAIL.n495 4.26717
R789 VTAIL.n479 VTAIL.n456 4.26717
R790 VTAIL.n422 VTAIL.n421 4.26717
R791 VTAIL.n405 VTAIL.n382 4.26717
R792 VTAIL.n350 VTAIL.n349 4.26717
R793 VTAIL.n333 VTAIL.n310 4.26717
R794 VTAIL.n276 VTAIL.n275 4.26717
R795 VTAIL.n259 VTAIL.n236 4.26717
R796 VTAIL.n535 VTAIL.n533 3.70982
R797 VTAIL.n25 VTAIL.n23 3.70982
R798 VTAIL.n97 VTAIL.n95 3.70982
R799 VTAIL.n171 VTAIL.n169 3.70982
R800 VTAIL.n463 VTAIL.n461 3.70982
R801 VTAIL.n389 VTAIL.n387 3.70982
R802 VTAIL.n317 VTAIL.n315 3.70982
R803 VTAIL.n243 VTAIL.n241 3.70982
R804 VTAIL.n548 VTAIL.n547 3.49141
R805 VTAIL.n571 VTAIL.n518 3.49141
R806 VTAIL.n38 VTAIL.n37 3.49141
R807 VTAIL.n61 VTAIL.n8 3.49141
R808 VTAIL.n110 VTAIL.n109 3.49141
R809 VTAIL.n133 VTAIL.n80 3.49141
R810 VTAIL.n184 VTAIL.n183 3.49141
R811 VTAIL.n207 VTAIL.n154 3.49141
R812 VTAIL.n499 VTAIL.n446 3.49141
R813 VTAIL.n476 VTAIL.n475 3.49141
R814 VTAIL.n425 VTAIL.n372 3.49141
R815 VTAIL.n402 VTAIL.n401 3.49141
R816 VTAIL.n353 VTAIL.n300 3.49141
R817 VTAIL.n330 VTAIL.n329 3.49141
R818 VTAIL.n279 VTAIL.n226 3.49141
R819 VTAIL.n256 VTAIL.n255 3.49141
R820 VTAIL.n293 VTAIL.n291 2.75912
R821 VTAIL.n365 VTAIL.n293 2.75912
R822 VTAIL.n439 VTAIL.n437 2.75912
R823 VTAIL.n511 VTAIL.n439 2.75912
R824 VTAIL.n219 VTAIL.n147 2.75912
R825 VTAIL.n147 VTAIL.n145 2.75912
R826 VTAIL.n73 VTAIL.n1 2.75912
R827 VTAIL.n544 VTAIL.n530 2.71565
R828 VTAIL.n572 VTAIL.n516 2.71565
R829 VTAIL.n34 VTAIL.n20 2.71565
R830 VTAIL.n62 VTAIL.n6 2.71565
R831 VTAIL.n106 VTAIL.n92 2.71565
R832 VTAIL.n134 VTAIL.n78 2.71565
R833 VTAIL.n180 VTAIL.n166 2.71565
R834 VTAIL.n208 VTAIL.n152 2.71565
R835 VTAIL.n500 VTAIL.n444 2.71565
R836 VTAIL.n472 VTAIL.n458 2.71565
R837 VTAIL.n426 VTAIL.n370 2.71565
R838 VTAIL.n398 VTAIL.n384 2.71565
R839 VTAIL.n354 VTAIL.n298 2.71565
R840 VTAIL.n326 VTAIL.n312 2.71565
R841 VTAIL.n280 VTAIL.n224 2.71565
R842 VTAIL.n252 VTAIL.n238 2.71565
R843 VTAIL VTAIL.n583 2.70093
R844 VTAIL.n0 VTAIL.t1 2.42263
R845 VTAIL.n0 VTAIL.t7 2.42263
R846 VTAIL.n146 VTAIL.t12 2.42263
R847 VTAIL.n146 VTAIL.t9 2.42263
R848 VTAIL.n438 VTAIL.t13 2.42263
R849 VTAIL.n438 VTAIL.t11 2.42263
R850 VTAIL.n292 VTAIL.t6 2.42263
R851 VTAIL.n292 VTAIL.t4 2.42263
R852 VTAIL.n543 VTAIL.n532 1.93989
R853 VTAIL.n576 VTAIL.n575 1.93989
R854 VTAIL.n33 VTAIL.n22 1.93989
R855 VTAIL.n66 VTAIL.n65 1.93989
R856 VTAIL.n105 VTAIL.n94 1.93989
R857 VTAIL.n138 VTAIL.n137 1.93989
R858 VTAIL.n179 VTAIL.n168 1.93989
R859 VTAIL.n212 VTAIL.n211 1.93989
R860 VTAIL.n504 VTAIL.n503 1.93989
R861 VTAIL.n471 VTAIL.n460 1.93989
R862 VTAIL.n430 VTAIL.n429 1.93989
R863 VTAIL.n397 VTAIL.n386 1.93989
R864 VTAIL.n358 VTAIL.n357 1.93989
R865 VTAIL.n325 VTAIL.n314 1.93989
R866 VTAIL.n284 VTAIL.n283 1.93989
R867 VTAIL.n251 VTAIL.n240 1.93989
R868 VTAIL.n540 VTAIL.n539 1.16414
R869 VTAIL.n579 VTAIL.n514 1.16414
R870 VTAIL.n30 VTAIL.n29 1.16414
R871 VTAIL.n69 VTAIL.n4 1.16414
R872 VTAIL.n102 VTAIL.n101 1.16414
R873 VTAIL.n141 VTAIL.n76 1.16414
R874 VTAIL.n176 VTAIL.n175 1.16414
R875 VTAIL.n215 VTAIL.n150 1.16414
R876 VTAIL.n507 VTAIL.n442 1.16414
R877 VTAIL.n468 VTAIL.n467 1.16414
R878 VTAIL.n433 VTAIL.n368 1.16414
R879 VTAIL.n394 VTAIL.n393 1.16414
R880 VTAIL.n361 VTAIL.n296 1.16414
R881 VTAIL.n322 VTAIL.n321 1.16414
R882 VTAIL.n287 VTAIL.n222 1.16414
R883 VTAIL.n248 VTAIL.n247 1.16414
R884 VTAIL.n437 VTAIL.n365 0.470328
R885 VTAIL.n145 VTAIL.n73 0.470328
R886 VTAIL.n536 VTAIL.n534 0.388379
R887 VTAIL.n26 VTAIL.n24 0.388379
R888 VTAIL.n98 VTAIL.n96 0.388379
R889 VTAIL.n172 VTAIL.n170 0.388379
R890 VTAIL.n464 VTAIL.n462 0.388379
R891 VTAIL.n390 VTAIL.n388 0.388379
R892 VTAIL.n318 VTAIL.n316 0.388379
R893 VTAIL.n244 VTAIL.n242 0.388379
R894 VTAIL.n541 VTAIL.n533 0.155672
R895 VTAIL.n542 VTAIL.n541 0.155672
R896 VTAIL.n542 VTAIL.n529 0.155672
R897 VTAIL.n549 VTAIL.n529 0.155672
R898 VTAIL.n550 VTAIL.n549 0.155672
R899 VTAIL.n550 VTAIL.n525 0.155672
R900 VTAIL.n557 VTAIL.n525 0.155672
R901 VTAIL.n558 VTAIL.n557 0.155672
R902 VTAIL.n558 VTAIL.n521 0.155672
R903 VTAIL.n565 VTAIL.n521 0.155672
R904 VTAIL.n566 VTAIL.n565 0.155672
R905 VTAIL.n566 VTAIL.n517 0.155672
R906 VTAIL.n573 VTAIL.n517 0.155672
R907 VTAIL.n574 VTAIL.n573 0.155672
R908 VTAIL.n574 VTAIL.n513 0.155672
R909 VTAIL.n581 VTAIL.n513 0.155672
R910 VTAIL.n31 VTAIL.n23 0.155672
R911 VTAIL.n32 VTAIL.n31 0.155672
R912 VTAIL.n32 VTAIL.n19 0.155672
R913 VTAIL.n39 VTAIL.n19 0.155672
R914 VTAIL.n40 VTAIL.n39 0.155672
R915 VTAIL.n40 VTAIL.n15 0.155672
R916 VTAIL.n47 VTAIL.n15 0.155672
R917 VTAIL.n48 VTAIL.n47 0.155672
R918 VTAIL.n48 VTAIL.n11 0.155672
R919 VTAIL.n55 VTAIL.n11 0.155672
R920 VTAIL.n56 VTAIL.n55 0.155672
R921 VTAIL.n56 VTAIL.n7 0.155672
R922 VTAIL.n63 VTAIL.n7 0.155672
R923 VTAIL.n64 VTAIL.n63 0.155672
R924 VTAIL.n64 VTAIL.n3 0.155672
R925 VTAIL.n71 VTAIL.n3 0.155672
R926 VTAIL.n103 VTAIL.n95 0.155672
R927 VTAIL.n104 VTAIL.n103 0.155672
R928 VTAIL.n104 VTAIL.n91 0.155672
R929 VTAIL.n111 VTAIL.n91 0.155672
R930 VTAIL.n112 VTAIL.n111 0.155672
R931 VTAIL.n112 VTAIL.n87 0.155672
R932 VTAIL.n119 VTAIL.n87 0.155672
R933 VTAIL.n120 VTAIL.n119 0.155672
R934 VTAIL.n120 VTAIL.n83 0.155672
R935 VTAIL.n127 VTAIL.n83 0.155672
R936 VTAIL.n128 VTAIL.n127 0.155672
R937 VTAIL.n128 VTAIL.n79 0.155672
R938 VTAIL.n135 VTAIL.n79 0.155672
R939 VTAIL.n136 VTAIL.n135 0.155672
R940 VTAIL.n136 VTAIL.n75 0.155672
R941 VTAIL.n143 VTAIL.n75 0.155672
R942 VTAIL.n177 VTAIL.n169 0.155672
R943 VTAIL.n178 VTAIL.n177 0.155672
R944 VTAIL.n178 VTAIL.n165 0.155672
R945 VTAIL.n185 VTAIL.n165 0.155672
R946 VTAIL.n186 VTAIL.n185 0.155672
R947 VTAIL.n186 VTAIL.n161 0.155672
R948 VTAIL.n193 VTAIL.n161 0.155672
R949 VTAIL.n194 VTAIL.n193 0.155672
R950 VTAIL.n194 VTAIL.n157 0.155672
R951 VTAIL.n201 VTAIL.n157 0.155672
R952 VTAIL.n202 VTAIL.n201 0.155672
R953 VTAIL.n202 VTAIL.n153 0.155672
R954 VTAIL.n209 VTAIL.n153 0.155672
R955 VTAIL.n210 VTAIL.n209 0.155672
R956 VTAIL.n210 VTAIL.n149 0.155672
R957 VTAIL.n217 VTAIL.n149 0.155672
R958 VTAIL.n509 VTAIL.n441 0.155672
R959 VTAIL.n502 VTAIL.n441 0.155672
R960 VTAIL.n502 VTAIL.n501 0.155672
R961 VTAIL.n501 VTAIL.n445 0.155672
R962 VTAIL.n494 VTAIL.n445 0.155672
R963 VTAIL.n494 VTAIL.n493 0.155672
R964 VTAIL.n493 VTAIL.n449 0.155672
R965 VTAIL.n486 VTAIL.n449 0.155672
R966 VTAIL.n486 VTAIL.n485 0.155672
R967 VTAIL.n485 VTAIL.n453 0.155672
R968 VTAIL.n478 VTAIL.n453 0.155672
R969 VTAIL.n478 VTAIL.n477 0.155672
R970 VTAIL.n477 VTAIL.n457 0.155672
R971 VTAIL.n470 VTAIL.n457 0.155672
R972 VTAIL.n470 VTAIL.n469 0.155672
R973 VTAIL.n469 VTAIL.n461 0.155672
R974 VTAIL.n435 VTAIL.n367 0.155672
R975 VTAIL.n428 VTAIL.n367 0.155672
R976 VTAIL.n428 VTAIL.n427 0.155672
R977 VTAIL.n427 VTAIL.n371 0.155672
R978 VTAIL.n420 VTAIL.n371 0.155672
R979 VTAIL.n420 VTAIL.n419 0.155672
R980 VTAIL.n419 VTAIL.n375 0.155672
R981 VTAIL.n412 VTAIL.n375 0.155672
R982 VTAIL.n412 VTAIL.n411 0.155672
R983 VTAIL.n411 VTAIL.n379 0.155672
R984 VTAIL.n404 VTAIL.n379 0.155672
R985 VTAIL.n404 VTAIL.n403 0.155672
R986 VTAIL.n403 VTAIL.n383 0.155672
R987 VTAIL.n396 VTAIL.n383 0.155672
R988 VTAIL.n396 VTAIL.n395 0.155672
R989 VTAIL.n395 VTAIL.n387 0.155672
R990 VTAIL.n363 VTAIL.n295 0.155672
R991 VTAIL.n356 VTAIL.n295 0.155672
R992 VTAIL.n356 VTAIL.n355 0.155672
R993 VTAIL.n355 VTAIL.n299 0.155672
R994 VTAIL.n348 VTAIL.n299 0.155672
R995 VTAIL.n348 VTAIL.n347 0.155672
R996 VTAIL.n347 VTAIL.n303 0.155672
R997 VTAIL.n340 VTAIL.n303 0.155672
R998 VTAIL.n340 VTAIL.n339 0.155672
R999 VTAIL.n339 VTAIL.n307 0.155672
R1000 VTAIL.n332 VTAIL.n307 0.155672
R1001 VTAIL.n332 VTAIL.n331 0.155672
R1002 VTAIL.n331 VTAIL.n311 0.155672
R1003 VTAIL.n324 VTAIL.n311 0.155672
R1004 VTAIL.n324 VTAIL.n323 0.155672
R1005 VTAIL.n323 VTAIL.n315 0.155672
R1006 VTAIL.n289 VTAIL.n221 0.155672
R1007 VTAIL.n282 VTAIL.n221 0.155672
R1008 VTAIL.n282 VTAIL.n281 0.155672
R1009 VTAIL.n281 VTAIL.n225 0.155672
R1010 VTAIL.n274 VTAIL.n225 0.155672
R1011 VTAIL.n274 VTAIL.n273 0.155672
R1012 VTAIL.n273 VTAIL.n229 0.155672
R1013 VTAIL.n266 VTAIL.n229 0.155672
R1014 VTAIL.n266 VTAIL.n265 0.155672
R1015 VTAIL.n265 VTAIL.n233 0.155672
R1016 VTAIL.n258 VTAIL.n233 0.155672
R1017 VTAIL.n258 VTAIL.n257 0.155672
R1018 VTAIL.n257 VTAIL.n237 0.155672
R1019 VTAIL.n250 VTAIL.n237 0.155672
R1020 VTAIL.n250 VTAIL.n249 0.155672
R1021 VTAIL.n249 VTAIL.n241 0.155672
R1022 VTAIL VTAIL.n1 0.0586897
R1023 B.n624 B.n623 585
R1024 B.n625 B.n84 585
R1025 B.n627 B.n626 585
R1026 B.n628 B.n83 585
R1027 B.n630 B.n629 585
R1028 B.n631 B.n82 585
R1029 B.n633 B.n632 585
R1030 B.n634 B.n81 585
R1031 B.n636 B.n635 585
R1032 B.n637 B.n80 585
R1033 B.n639 B.n638 585
R1034 B.n640 B.n79 585
R1035 B.n642 B.n641 585
R1036 B.n643 B.n78 585
R1037 B.n645 B.n644 585
R1038 B.n646 B.n77 585
R1039 B.n648 B.n647 585
R1040 B.n649 B.n76 585
R1041 B.n651 B.n650 585
R1042 B.n652 B.n75 585
R1043 B.n654 B.n653 585
R1044 B.n655 B.n74 585
R1045 B.n657 B.n656 585
R1046 B.n658 B.n73 585
R1047 B.n660 B.n659 585
R1048 B.n661 B.n72 585
R1049 B.n663 B.n662 585
R1050 B.n664 B.n71 585
R1051 B.n666 B.n665 585
R1052 B.n667 B.n70 585
R1053 B.n669 B.n668 585
R1054 B.n670 B.n69 585
R1055 B.n672 B.n671 585
R1056 B.n673 B.n68 585
R1057 B.n675 B.n674 585
R1058 B.n676 B.n67 585
R1059 B.n678 B.n677 585
R1060 B.n679 B.n66 585
R1061 B.n681 B.n680 585
R1062 B.n682 B.n65 585
R1063 B.n684 B.n683 585
R1064 B.n685 B.n64 585
R1065 B.n687 B.n686 585
R1066 B.n688 B.n63 585
R1067 B.n690 B.n689 585
R1068 B.n691 B.n60 585
R1069 B.n694 B.n693 585
R1070 B.n695 B.n59 585
R1071 B.n697 B.n696 585
R1072 B.n698 B.n58 585
R1073 B.n700 B.n699 585
R1074 B.n701 B.n57 585
R1075 B.n703 B.n702 585
R1076 B.n704 B.n53 585
R1077 B.n706 B.n705 585
R1078 B.n707 B.n52 585
R1079 B.n709 B.n708 585
R1080 B.n710 B.n51 585
R1081 B.n712 B.n711 585
R1082 B.n713 B.n50 585
R1083 B.n715 B.n714 585
R1084 B.n716 B.n49 585
R1085 B.n718 B.n717 585
R1086 B.n719 B.n48 585
R1087 B.n721 B.n720 585
R1088 B.n722 B.n47 585
R1089 B.n724 B.n723 585
R1090 B.n725 B.n46 585
R1091 B.n727 B.n726 585
R1092 B.n728 B.n45 585
R1093 B.n730 B.n729 585
R1094 B.n731 B.n44 585
R1095 B.n733 B.n732 585
R1096 B.n734 B.n43 585
R1097 B.n736 B.n735 585
R1098 B.n737 B.n42 585
R1099 B.n739 B.n738 585
R1100 B.n740 B.n41 585
R1101 B.n742 B.n741 585
R1102 B.n743 B.n40 585
R1103 B.n745 B.n744 585
R1104 B.n746 B.n39 585
R1105 B.n748 B.n747 585
R1106 B.n749 B.n38 585
R1107 B.n751 B.n750 585
R1108 B.n752 B.n37 585
R1109 B.n754 B.n753 585
R1110 B.n755 B.n36 585
R1111 B.n757 B.n756 585
R1112 B.n758 B.n35 585
R1113 B.n760 B.n759 585
R1114 B.n761 B.n34 585
R1115 B.n763 B.n762 585
R1116 B.n764 B.n33 585
R1117 B.n766 B.n765 585
R1118 B.n767 B.n32 585
R1119 B.n769 B.n768 585
R1120 B.n770 B.n31 585
R1121 B.n772 B.n771 585
R1122 B.n773 B.n30 585
R1123 B.n775 B.n774 585
R1124 B.n622 B.n85 585
R1125 B.n621 B.n620 585
R1126 B.n619 B.n86 585
R1127 B.n618 B.n617 585
R1128 B.n616 B.n87 585
R1129 B.n615 B.n614 585
R1130 B.n613 B.n88 585
R1131 B.n612 B.n611 585
R1132 B.n610 B.n89 585
R1133 B.n609 B.n608 585
R1134 B.n607 B.n90 585
R1135 B.n606 B.n605 585
R1136 B.n604 B.n91 585
R1137 B.n603 B.n602 585
R1138 B.n601 B.n92 585
R1139 B.n600 B.n599 585
R1140 B.n598 B.n93 585
R1141 B.n597 B.n596 585
R1142 B.n595 B.n94 585
R1143 B.n594 B.n593 585
R1144 B.n592 B.n95 585
R1145 B.n591 B.n590 585
R1146 B.n589 B.n96 585
R1147 B.n588 B.n587 585
R1148 B.n586 B.n97 585
R1149 B.n585 B.n584 585
R1150 B.n583 B.n98 585
R1151 B.n582 B.n581 585
R1152 B.n580 B.n99 585
R1153 B.n579 B.n578 585
R1154 B.n577 B.n100 585
R1155 B.n576 B.n575 585
R1156 B.n574 B.n101 585
R1157 B.n573 B.n572 585
R1158 B.n571 B.n102 585
R1159 B.n570 B.n569 585
R1160 B.n568 B.n103 585
R1161 B.n567 B.n566 585
R1162 B.n565 B.n104 585
R1163 B.n564 B.n563 585
R1164 B.n562 B.n105 585
R1165 B.n561 B.n560 585
R1166 B.n559 B.n106 585
R1167 B.n558 B.n557 585
R1168 B.n556 B.n107 585
R1169 B.n555 B.n554 585
R1170 B.n553 B.n108 585
R1171 B.n552 B.n551 585
R1172 B.n550 B.n109 585
R1173 B.n549 B.n548 585
R1174 B.n547 B.n110 585
R1175 B.n546 B.n545 585
R1176 B.n544 B.n111 585
R1177 B.n543 B.n542 585
R1178 B.n541 B.n112 585
R1179 B.n540 B.n539 585
R1180 B.n538 B.n113 585
R1181 B.n537 B.n536 585
R1182 B.n535 B.n114 585
R1183 B.n534 B.n533 585
R1184 B.n532 B.n115 585
R1185 B.n531 B.n530 585
R1186 B.n529 B.n116 585
R1187 B.n528 B.n527 585
R1188 B.n526 B.n117 585
R1189 B.n525 B.n524 585
R1190 B.n523 B.n118 585
R1191 B.n522 B.n521 585
R1192 B.n520 B.n119 585
R1193 B.n519 B.n518 585
R1194 B.n517 B.n120 585
R1195 B.n516 B.n515 585
R1196 B.n514 B.n121 585
R1197 B.n513 B.n512 585
R1198 B.n511 B.n122 585
R1199 B.n510 B.n509 585
R1200 B.n508 B.n123 585
R1201 B.n507 B.n506 585
R1202 B.n505 B.n124 585
R1203 B.n504 B.n503 585
R1204 B.n502 B.n125 585
R1205 B.n501 B.n500 585
R1206 B.n499 B.n126 585
R1207 B.n498 B.n497 585
R1208 B.n496 B.n127 585
R1209 B.n495 B.n494 585
R1210 B.n493 B.n128 585
R1211 B.n492 B.n491 585
R1212 B.n490 B.n129 585
R1213 B.n489 B.n488 585
R1214 B.n487 B.n130 585
R1215 B.n486 B.n485 585
R1216 B.n484 B.n131 585
R1217 B.n483 B.n482 585
R1218 B.n481 B.n132 585
R1219 B.n480 B.n479 585
R1220 B.n478 B.n133 585
R1221 B.n477 B.n476 585
R1222 B.n475 B.n134 585
R1223 B.n474 B.n473 585
R1224 B.n472 B.n135 585
R1225 B.n471 B.n470 585
R1226 B.n469 B.n136 585
R1227 B.n468 B.n467 585
R1228 B.n466 B.n137 585
R1229 B.n465 B.n464 585
R1230 B.n463 B.n138 585
R1231 B.n462 B.n461 585
R1232 B.n460 B.n139 585
R1233 B.n459 B.n458 585
R1234 B.n457 B.n140 585
R1235 B.n302 B.n301 585
R1236 B.n303 B.n192 585
R1237 B.n305 B.n304 585
R1238 B.n306 B.n191 585
R1239 B.n308 B.n307 585
R1240 B.n309 B.n190 585
R1241 B.n311 B.n310 585
R1242 B.n312 B.n189 585
R1243 B.n314 B.n313 585
R1244 B.n315 B.n188 585
R1245 B.n317 B.n316 585
R1246 B.n318 B.n187 585
R1247 B.n320 B.n319 585
R1248 B.n321 B.n186 585
R1249 B.n323 B.n322 585
R1250 B.n324 B.n185 585
R1251 B.n326 B.n325 585
R1252 B.n327 B.n184 585
R1253 B.n329 B.n328 585
R1254 B.n330 B.n183 585
R1255 B.n332 B.n331 585
R1256 B.n333 B.n182 585
R1257 B.n335 B.n334 585
R1258 B.n336 B.n181 585
R1259 B.n338 B.n337 585
R1260 B.n339 B.n180 585
R1261 B.n341 B.n340 585
R1262 B.n342 B.n179 585
R1263 B.n344 B.n343 585
R1264 B.n345 B.n178 585
R1265 B.n347 B.n346 585
R1266 B.n348 B.n177 585
R1267 B.n350 B.n349 585
R1268 B.n351 B.n176 585
R1269 B.n353 B.n352 585
R1270 B.n354 B.n175 585
R1271 B.n356 B.n355 585
R1272 B.n357 B.n174 585
R1273 B.n359 B.n358 585
R1274 B.n360 B.n173 585
R1275 B.n362 B.n361 585
R1276 B.n363 B.n172 585
R1277 B.n365 B.n364 585
R1278 B.n366 B.n171 585
R1279 B.n368 B.n367 585
R1280 B.n369 B.n168 585
R1281 B.n372 B.n371 585
R1282 B.n373 B.n167 585
R1283 B.n375 B.n374 585
R1284 B.n376 B.n166 585
R1285 B.n378 B.n377 585
R1286 B.n379 B.n165 585
R1287 B.n381 B.n380 585
R1288 B.n382 B.n164 585
R1289 B.n387 B.n386 585
R1290 B.n388 B.n163 585
R1291 B.n390 B.n389 585
R1292 B.n391 B.n162 585
R1293 B.n393 B.n392 585
R1294 B.n394 B.n161 585
R1295 B.n396 B.n395 585
R1296 B.n397 B.n160 585
R1297 B.n399 B.n398 585
R1298 B.n400 B.n159 585
R1299 B.n402 B.n401 585
R1300 B.n403 B.n158 585
R1301 B.n405 B.n404 585
R1302 B.n406 B.n157 585
R1303 B.n408 B.n407 585
R1304 B.n409 B.n156 585
R1305 B.n411 B.n410 585
R1306 B.n412 B.n155 585
R1307 B.n414 B.n413 585
R1308 B.n415 B.n154 585
R1309 B.n417 B.n416 585
R1310 B.n418 B.n153 585
R1311 B.n420 B.n419 585
R1312 B.n421 B.n152 585
R1313 B.n423 B.n422 585
R1314 B.n424 B.n151 585
R1315 B.n426 B.n425 585
R1316 B.n427 B.n150 585
R1317 B.n429 B.n428 585
R1318 B.n430 B.n149 585
R1319 B.n432 B.n431 585
R1320 B.n433 B.n148 585
R1321 B.n435 B.n434 585
R1322 B.n436 B.n147 585
R1323 B.n438 B.n437 585
R1324 B.n439 B.n146 585
R1325 B.n441 B.n440 585
R1326 B.n442 B.n145 585
R1327 B.n444 B.n443 585
R1328 B.n445 B.n144 585
R1329 B.n447 B.n446 585
R1330 B.n448 B.n143 585
R1331 B.n450 B.n449 585
R1332 B.n451 B.n142 585
R1333 B.n453 B.n452 585
R1334 B.n454 B.n141 585
R1335 B.n456 B.n455 585
R1336 B.n300 B.n193 585
R1337 B.n299 B.n298 585
R1338 B.n297 B.n194 585
R1339 B.n296 B.n295 585
R1340 B.n294 B.n195 585
R1341 B.n293 B.n292 585
R1342 B.n291 B.n196 585
R1343 B.n290 B.n289 585
R1344 B.n288 B.n197 585
R1345 B.n287 B.n286 585
R1346 B.n285 B.n198 585
R1347 B.n284 B.n283 585
R1348 B.n282 B.n199 585
R1349 B.n281 B.n280 585
R1350 B.n279 B.n200 585
R1351 B.n278 B.n277 585
R1352 B.n276 B.n201 585
R1353 B.n275 B.n274 585
R1354 B.n273 B.n202 585
R1355 B.n272 B.n271 585
R1356 B.n270 B.n203 585
R1357 B.n269 B.n268 585
R1358 B.n267 B.n204 585
R1359 B.n266 B.n265 585
R1360 B.n264 B.n205 585
R1361 B.n263 B.n262 585
R1362 B.n261 B.n206 585
R1363 B.n260 B.n259 585
R1364 B.n258 B.n207 585
R1365 B.n257 B.n256 585
R1366 B.n255 B.n208 585
R1367 B.n254 B.n253 585
R1368 B.n252 B.n209 585
R1369 B.n251 B.n250 585
R1370 B.n249 B.n210 585
R1371 B.n248 B.n247 585
R1372 B.n246 B.n211 585
R1373 B.n245 B.n244 585
R1374 B.n243 B.n212 585
R1375 B.n242 B.n241 585
R1376 B.n240 B.n213 585
R1377 B.n239 B.n238 585
R1378 B.n237 B.n214 585
R1379 B.n236 B.n235 585
R1380 B.n234 B.n215 585
R1381 B.n233 B.n232 585
R1382 B.n231 B.n216 585
R1383 B.n230 B.n229 585
R1384 B.n228 B.n217 585
R1385 B.n227 B.n226 585
R1386 B.n225 B.n218 585
R1387 B.n224 B.n223 585
R1388 B.n222 B.n219 585
R1389 B.n221 B.n220 585
R1390 B.n2 B.n0 585
R1391 B.n857 B.n1 585
R1392 B.n856 B.n855 585
R1393 B.n854 B.n3 585
R1394 B.n853 B.n852 585
R1395 B.n851 B.n4 585
R1396 B.n850 B.n849 585
R1397 B.n848 B.n5 585
R1398 B.n847 B.n846 585
R1399 B.n845 B.n6 585
R1400 B.n844 B.n843 585
R1401 B.n842 B.n7 585
R1402 B.n841 B.n840 585
R1403 B.n839 B.n8 585
R1404 B.n838 B.n837 585
R1405 B.n836 B.n9 585
R1406 B.n835 B.n834 585
R1407 B.n833 B.n10 585
R1408 B.n832 B.n831 585
R1409 B.n830 B.n11 585
R1410 B.n829 B.n828 585
R1411 B.n827 B.n12 585
R1412 B.n826 B.n825 585
R1413 B.n824 B.n13 585
R1414 B.n823 B.n822 585
R1415 B.n821 B.n14 585
R1416 B.n820 B.n819 585
R1417 B.n818 B.n15 585
R1418 B.n817 B.n816 585
R1419 B.n815 B.n16 585
R1420 B.n814 B.n813 585
R1421 B.n812 B.n17 585
R1422 B.n811 B.n810 585
R1423 B.n809 B.n18 585
R1424 B.n808 B.n807 585
R1425 B.n806 B.n19 585
R1426 B.n805 B.n804 585
R1427 B.n803 B.n20 585
R1428 B.n802 B.n801 585
R1429 B.n800 B.n21 585
R1430 B.n799 B.n798 585
R1431 B.n797 B.n22 585
R1432 B.n796 B.n795 585
R1433 B.n794 B.n23 585
R1434 B.n793 B.n792 585
R1435 B.n791 B.n24 585
R1436 B.n790 B.n789 585
R1437 B.n788 B.n25 585
R1438 B.n787 B.n786 585
R1439 B.n785 B.n26 585
R1440 B.n784 B.n783 585
R1441 B.n782 B.n27 585
R1442 B.n781 B.n780 585
R1443 B.n779 B.n28 585
R1444 B.n778 B.n777 585
R1445 B.n776 B.n29 585
R1446 B.n859 B.n858 585
R1447 B.n301 B.n300 540.549
R1448 B.n774 B.n29 540.549
R1449 B.n455 B.n140 540.549
R1450 B.n623 B.n622 540.549
R1451 B.n383 B.t5 463.248
R1452 B.n61 B.t7 463.248
R1453 B.n169 B.t11 463.248
R1454 B.n54 B.t1 463.248
R1455 B.n384 B.t4 401.188
R1456 B.n62 B.t8 401.188
R1457 B.n170 B.t10 401.188
R1458 B.n55 B.t2 401.188
R1459 B.n383 B.t3 321.111
R1460 B.n169 B.t9 321.111
R1461 B.n54 B.t0 321.111
R1462 B.n61 B.t6 321.111
R1463 B.n300 B.n299 163.367
R1464 B.n299 B.n194 163.367
R1465 B.n295 B.n194 163.367
R1466 B.n295 B.n294 163.367
R1467 B.n294 B.n293 163.367
R1468 B.n293 B.n196 163.367
R1469 B.n289 B.n196 163.367
R1470 B.n289 B.n288 163.367
R1471 B.n288 B.n287 163.367
R1472 B.n287 B.n198 163.367
R1473 B.n283 B.n198 163.367
R1474 B.n283 B.n282 163.367
R1475 B.n282 B.n281 163.367
R1476 B.n281 B.n200 163.367
R1477 B.n277 B.n200 163.367
R1478 B.n277 B.n276 163.367
R1479 B.n276 B.n275 163.367
R1480 B.n275 B.n202 163.367
R1481 B.n271 B.n202 163.367
R1482 B.n271 B.n270 163.367
R1483 B.n270 B.n269 163.367
R1484 B.n269 B.n204 163.367
R1485 B.n265 B.n204 163.367
R1486 B.n265 B.n264 163.367
R1487 B.n264 B.n263 163.367
R1488 B.n263 B.n206 163.367
R1489 B.n259 B.n206 163.367
R1490 B.n259 B.n258 163.367
R1491 B.n258 B.n257 163.367
R1492 B.n257 B.n208 163.367
R1493 B.n253 B.n208 163.367
R1494 B.n253 B.n252 163.367
R1495 B.n252 B.n251 163.367
R1496 B.n251 B.n210 163.367
R1497 B.n247 B.n210 163.367
R1498 B.n247 B.n246 163.367
R1499 B.n246 B.n245 163.367
R1500 B.n245 B.n212 163.367
R1501 B.n241 B.n212 163.367
R1502 B.n241 B.n240 163.367
R1503 B.n240 B.n239 163.367
R1504 B.n239 B.n214 163.367
R1505 B.n235 B.n214 163.367
R1506 B.n235 B.n234 163.367
R1507 B.n234 B.n233 163.367
R1508 B.n233 B.n216 163.367
R1509 B.n229 B.n216 163.367
R1510 B.n229 B.n228 163.367
R1511 B.n228 B.n227 163.367
R1512 B.n227 B.n218 163.367
R1513 B.n223 B.n218 163.367
R1514 B.n223 B.n222 163.367
R1515 B.n222 B.n221 163.367
R1516 B.n221 B.n2 163.367
R1517 B.n858 B.n2 163.367
R1518 B.n858 B.n857 163.367
R1519 B.n857 B.n856 163.367
R1520 B.n856 B.n3 163.367
R1521 B.n852 B.n3 163.367
R1522 B.n852 B.n851 163.367
R1523 B.n851 B.n850 163.367
R1524 B.n850 B.n5 163.367
R1525 B.n846 B.n5 163.367
R1526 B.n846 B.n845 163.367
R1527 B.n845 B.n844 163.367
R1528 B.n844 B.n7 163.367
R1529 B.n840 B.n7 163.367
R1530 B.n840 B.n839 163.367
R1531 B.n839 B.n838 163.367
R1532 B.n838 B.n9 163.367
R1533 B.n834 B.n9 163.367
R1534 B.n834 B.n833 163.367
R1535 B.n833 B.n832 163.367
R1536 B.n832 B.n11 163.367
R1537 B.n828 B.n11 163.367
R1538 B.n828 B.n827 163.367
R1539 B.n827 B.n826 163.367
R1540 B.n826 B.n13 163.367
R1541 B.n822 B.n13 163.367
R1542 B.n822 B.n821 163.367
R1543 B.n821 B.n820 163.367
R1544 B.n820 B.n15 163.367
R1545 B.n816 B.n15 163.367
R1546 B.n816 B.n815 163.367
R1547 B.n815 B.n814 163.367
R1548 B.n814 B.n17 163.367
R1549 B.n810 B.n17 163.367
R1550 B.n810 B.n809 163.367
R1551 B.n809 B.n808 163.367
R1552 B.n808 B.n19 163.367
R1553 B.n804 B.n19 163.367
R1554 B.n804 B.n803 163.367
R1555 B.n803 B.n802 163.367
R1556 B.n802 B.n21 163.367
R1557 B.n798 B.n21 163.367
R1558 B.n798 B.n797 163.367
R1559 B.n797 B.n796 163.367
R1560 B.n796 B.n23 163.367
R1561 B.n792 B.n23 163.367
R1562 B.n792 B.n791 163.367
R1563 B.n791 B.n790 163.367
R1564 B.n790 B.n25 163.367
R1565 B.n786 B.n25 163.367
R1566 B.n786 B.n785 163.367
R1567 B.n785 B.n784 163.367
R1568 B.n784 B.n27 163.367
R1569 B.n780 B.n27 163.367
R1570 B.n780 B.n779 163.367
R1571 B.n779 B.n778 163.367
R1572 B.n778 B.n29 163.367
R1573 B.n301 B.n192 163.367
R1574 B.n305 B.n192 163.367
R1575 B.n306 B.n305 163.367
R1576 B.n307 B.n306 163.367
R1577 B.n307 B.n190 163.367
R1578 B.n311 B.n190 163.367
R1579 B.n312 B.n311 163.367
R1580 B.n313 B.n312 163.367
R1581 B.n313 B.n188 163.367
R1582 B.n317 B.n188 163.367
R1583 B.n318 B.n317 163.367
R1584 B.n319 B.n318 163.367
R1585 B.n319 B.n186 163.367
R1586 B.n323 B.n186 163.367
R1587 B.n324 B.n323 163.367
R1588 B.n325 B.n324 163.367
R1589 B.n325 B.n184 163.367
R1590 B.n329 B.n184 163.367
R1591 B.n330 B.n329 163.367
R1592 B.n331 B.n330 163.367
R1593 B.n331 B.n182 163.367
R1594 B.n335 B.n182 163.367
R1595 B.n336 B.n335 163.367
R1596 B.n337 B.n336 163.367
R1597 B.n337 B.n180 163.367
R1598 B.n341 B.n180 163.367
R1599 B.n342 B.n341 163.367
R1600 B.n343 B.n342 163.367
R1601 B.n343 B.n178 163.367
R1602 B.n347 B.n178 163.367
R1603 B.n348 B.n347 163.367
R1604 B.n349 B.n348 163.367
R1605 B.n349 B.n176 163.367
R1606 B.n353 B.n176 163.367
R1607 B.n354 B.n353 163.367
R1608 B.n355 B.n354 163.367
R1609 B.n355 B.n174 163.367
R1610 B.n359 B.n174 163.367
R1611 B.n360 B.n359 163.367
R1612 B.n361 B.n360 163.367
R1613 B.n361 B.n172 163.367
R1614 B.n365 B.n172 163.367
R1615 B.n366 B.n365 163.367
R1616 B.n367 B.n366 163.367
R1617 B.n367 B.n168 163.367
R1618 B.n372 B.n168 163.367
R1619 B.n373 B.n372 163.367
R1620 B.n374 B.n373 163.367
R1621 B.n374 B.n166 163.367
R1622 B.n378 B.n166 163.367
R1623 B.n379 B.n378 163.367
R1624 B.n380 B.n379 163.367
R1625 B.n380 B.n164 163.367
R1626 B.n387 B.n164 163.367
R1627 B.n388 B.n387 163.367
R1628 B.n389 B.n388 163.367
R1629 B.n389 B.n162 163.367
R1630 B.n393 B.n162 163.367
R1631 B.n394 B.n393 163.367
R1632 B.n395 B.n394 163.367
R1633 B.n395 B.n160 163.367
R1634 B.n399 B.n160 163.367
R1635 B.n400 B.n399 163.367
R1636 B.n401 B.n400 163.367
R1637 B.n401 B.n158 163.367
R1638 B.n405 B.n158 163.367
R1639 B.n406 B.n405 163.367
R1640 B.n407 B.n406 163.367
R1641 B.n407 B.n156 163.367
R1642 B.n411 B.n156 163.367
R1643 B.n412 B.n411 163.367
R1644 B.n413 B.n412 163.367
R1645 B.n413 B.n154 163.367
R1646 B.n417 B.n154 163.367
R1647 B.n418 B.n417 163.367
R1648 B.n419 B.n418 163.367
R1649 B.n419 B.n152 163.367
R1650 B.n423 B.n152 163.367
R1651 B.n424 B.n423 163.367
R1652 B.n425 B.n424 163.367
R1653 B.n425 B.n150 163.367
R1654 B.n429 B.n150 163.367
R1655 B.n430 B.n429 163.367
R1656 B.n431 B.n430 163.367
R1657 B.n431 B.n148 163.367
R1658 B.n435 B.n148 163.367
R1659 B.n436 B.n435 163.367
R1660 B.n437 B.n436 163.367
R1661 B.n437 B.n146 163.367
R1662 B.n441 B.n146 163.367
R1663 B.n442 B.n441 163.367
R1664 B.n443 B.n442 163.367
R1665 B.n443 B.n144 163.367
R1666 B.n447 B.n144 163.367
R1667 B.n448 B.n447 163.367
R1668 B.n449 B.n448 163.367
R1669 B.n449 B.n142 163.367
R1670 B.n453 B.n142 163.367
R1671 B.n454 B.n453 163.367
R1672 B.n455 B.n454 163.367
R1673 B.n459 B.n140 163.367
R1674 B.n460 B.n459 163.367
R1675 B.n461 B.n460 163.367
R1676 B.n461 B.n138 163.367
R1677 B.n465 B.n138 163.367
R1678 B.n466 B.n465 163.367
R1679 B.n467 B.n466 163.367
R1680 B.n467 B.n136 163.367
R1681 B.n471 B.n136 163.367
R1682 B.n472 B.n471 163.367
R1683 B.n473 B.n472 163.367
R1684 B.n473 B.n134 163.367
R1685 B.n477 B.n134 163.367
R1686 B.n478 B.n477 163.367
R1687 B.n479 B.n478 163.367
R1688 B.n479 B.n132 163.367
R1689 B.n483 B.n132 163.367
R1690 B.n484 B.n483 163.367
R1691 B.n485 B.n484 163.367
R1692 B.n485 B.n130 163.367
R1693 B.n489 B.n130 163.367
R1694 B.n490 B.n489 163.367
R1695 B.n491 B.n490 163.367
R1696 B.n491 B.n128 163.367
R1697 B.n495 B.n128 163.367
R1698 B.n496 B.n495 163.367
R1699 B.n497 B.n496 163.367
R1700 B.n497 B.n126 163.367
R1701 B.n501 B.n126 163.367
R1702 B.n502 B.n501 163.367
R1703 B.n503 B.n502 163.367
R1704 B.n503 B.n124 163.367
R1705 B.n507 B.n124 163.367
R1706 B.n508 B.n507 163.367
R1707 B.n509 B.n508 163.367
R1708 B.n509 B.n122 163.367
R1709 B.n513 B.n122 163.367
R1710 B.n514 B.n513 163.367
R1711 B.n515 B.n514 163.367
R1712 B.n515 B.n120 163.367
R1713 B.n519 B.n120 163.367
R1714 B.n520 B.n519 163.367
R1715 B.n521 B.n520 163.367
R1716 B.n521 B.n118 163.367
R1717 B.n525 B.n118 163.367
R1718 B.n526 B.n525 163.367
R1719 B.n527 B.n526 163.367
R1720 B.n527 B.n116 163.367
R1721 B.n531 B.n116 163.367
R1722 B.n532 B.n531 163.367
R1723 B.n533 B.n532 163.367
R1724 B.n533 B.n114 163.367
R1725 B.n537 B.n114 163.367
R1726 B.n538 B.n537 163.367
R1727 B.n539 B.n538 163.367
R1728 B.n539 B.n112 163.367
R1729 B.n543 B.n112 163.367
R1730 B.n544 B.n543 163.367
R1731 B.n545 B.n544 163.367
R1732 B.n545 B.n110 163.367
R1733 B.n549 B.n110 163.367
R1734 B.n550 B.n549 163.367
R1735 B.n551 B.n550 163.367
R1736 B.n551 B.n108 163.367
R1737 B.n555 B.n108 163.367
R1738 B.n556 B.n555 163.367
R1739 B.n557 B.n556 163.367
R1740 B.n557 B.n106 163.367
R1741 B.n561 B.n106 163.367
R1742 B.n562 B.n561 163.367
R1743 B.n563 B.n562 163.367
R1744 B.n563 B.n104 163.367
R1745 B.n567 B.n104 163.367
R1746 B.n568 B.n567 163.367
R1747 B.n569 B.n568 163.367
R1748 B.n569 B.n102 163.367
R1749 B.n573 B.n102 163.367
R1750 B.n574 B.n573 163.367
R1751 B.n575 B.n574 163.367
R1752 B.n575 B.n100 163.367
R1753 B.n579 B.n100 163.367
R1754 B.n580 B.n579 163.367
R1755 B.n581 B.n580 163.367
R1756 B.n581 B.n98 163.367
R1757 B.n585 B.n98 163.367
R1758 B.n586 B.n585 163.367
R1759 B.n587 B.n586 163.367
R1760 B.n587 B.n96 163.367
R1761 B.n591 B.n96 163.367
R1762 B.n592 B.n591 163.367
R1763 B.n593 B.n592 163.367
R1764 B.n593 B.n94 163.367
R1765 B.n597 B.n94 163.367
R1766 B.n598 B.n597 163.367
R1767 B.n599 B.n598 163.367
R1768 B.n599 B.n92 163.367
R1769 B.n603 B.n92 163.367
R1770 B.n604 B.n603 163.367
R1771 B.n605 B.n604 163.367
R1772 B.n605 B.n90 163.367
R1773 B.n609 B.n90 163.367
R1774 B.n610 B.n609 163.367
R1775 B.n611 B.n610 163.367
R1776 B.n611 B.n88 163.367
R1777 B.n615 B.n88 163.367
R1778 B.n616 B.n615 163.367
R1779 B.n617 B.n616 163.367
R1780 B.n617 B.n86 163.367
R1781 B.n621 B.n86 163.367
R1782 B.n622 B.n621 163.367
R1783 B.n774 B.n773 163.367
R1784 B.n773 B.n772 163.367
R1785 B.n772 B.n31 163.367
R1786 B.n768 B.n31 163.367
R1787 B.n768 B.n767 163.367
R1788 B.n767 B.n766 163.367
R1789 B.n766 B.n33 163.367
R1790 B.n762 B.n33 163.367
R1791 B.n762 B.n761 163.367
R1792 B.n761 B.n760 163.367
R1793 B.n760 B.n35 163.367
R1794 B.n756 B.n35 163.367
R1795 B.n756 B.n755 163.367
R1796 B.n755 B.n754 163.367
R1797 B.n754 B.n37 163.367
R1798 B.n750 B.n37 163.367
R1799 B.n750 B.n749 163.367
R1800 B.n749 B.n748 163.367
R1801 B.n748 B.n39 163.367
R1802 B.n744 B.n39 163.367
R1803 B.n744 B.n743 163.367
R1804 B.n743 B.n742 163.367
R1805 B.n742 B.n41 163.367
R1806 B.n738 B.n41 163.367
R1807 B.n738 B.n737 163.367
R1808 B.n737 B.n736 163.367
R1809 B.n736 B.n43 163.367
R1810 B.n732 B.n43 163.367
R1811 B.n732 B.n731 163.367
R1812 B.n731 B.n730 163.367
R1813 B.n730 B.n45 163.367
R1814 B.n726 B.n45 163.367
R1815 B.n726 B.n725 163.367
R1816 B.n725 B.n724 163.367
R1817 B.n724 B.n47 163.367
R1818 B.n720 B.n47 163.367
R1819 B.n720 B.n719 163.367
R1820 B.n719 B.n718 163.367
R1821 B.n718 B.n49 163.367
R1822 B.n714 B.n49 163.367
R1823 B.n714 B.n713 163.367
R1824 B.n713 B.n712 163.367
R1825 B.n712 B.n51 163.367
R1826 B.n708 B.n51 163.367
R1827 B.n708 B.n707 163.367
R1828 B.n707 B.n706 163.367
R1829 B.n706 B.n53 163.367
R1830 B.n702 B.n53 163.367
R1831 B.n702 B.n701 163.367
R1832 B.n701 B.n700 163.367
R1833 B.n700 B.n58 163.367
R1834 B.n696 B.n58 163.367
R1835 B.n696 B.n695 163.367
R1836 B.n695 B.n694 163.367
R1837 B.n694 B.n60 163.367
R1838 B.n689 B.n60 163.367
R1839 B.n689 B.n688 163.367
R1840 B.n688 B.n687 163.367
R1841 B.n687 B.n64 163.367
R1842 B.n683 B.n64 163.367
R1843 B.n683 B.n682 163.367
R1844 B.n682 B.n681 163.367
R1845 B.n681 B.n66 163.367
R1846 B.n677 B.n66 163.367
R1847 B.n677 B.n676 163.367
R1848 B.n676 B.n675 163.367
R1849 B.n675 B.n68 163.367
R1850 B.n671 B.n68 163.367
R1851 B.n671 B.n670 163.367
R1852 B.n670 B.n669 163.367
R1853 B.n669 B.n70 163.367
R1854 B.n665 B.n70 163.367
R1855 B.n665 B.n664 163.367
R1856 B.n664 B.n663 163.367
R1857 B.n663 B.n72 163.367
R1858 B.n659 B.n72 163.367
R1859 B.n659 B.n658 163.367
R1860 B.n658 B.n657 163.367
R1861 B.n657 B.n74 163.367
R1862 B.n653 B.n74 163.367
R1863 B.n653 B.n652 163.367
R1864 B.n652 B.n651 163.367
R1865 B.n651 B.n76 163.367
R1866 B.n647 B.n76 163.367
R1867 B.n647 B.n646 163.367
R1868 B.n646 B.n645 163.367
R1869 B.n645 B.n78 163.367
R1870 B.n641 B.n78 163.367
R1871 B.n641 B.n640 163.367
R1872 B.n640 B.n639 163.367
R1873 B.n639 B.n80 163.367
R1874 B.n635 B.n80 163.367
R1875 B.n635 B.n634 163.367
R1876 B.n634 B.n633 163.367
R1877 B.n633 B.n82 163.367
R1878 B.n629 B.n82 163.367
R1879 B.n629 B.n628 163.367
R1880 B.n628 B.n627 163.367
R1881 B.n627 B.n84 163.367
R1882 B.n623 B.n84 163.367
R1883 B.n384 B.n383 62.0611
R1884 B.n170 B.n169 62.0611
R1885 B.n55 B.n54 62.0611
R1886 B.n62 B.n61 62.0611
R1887 B.n385 B.n384 59.5399
R1888 B.n370 B.n170 59.5399
R1889 B.n56 B.n55 59.5399
R1890 B.n692 B.n62 59.5399
R1891 B.n624 B.n85 35.1225
R1892 B.n776 B.n775 35.1224
R1893 B.n457 B.n456 35.1224
R1894 B.n302 B.n193 35.1224
R1895 B B.n859 18.0485
R1896 B.n775 B.n30 10.6151
R1897 B.n771 B.n30 10.6151
R1898 B.n771 B.n770 10.6151
R1899 B.n770 B.n769 10.6151
R1900 B.n769 B.n32 10.6151
R1901 B.n765 B.n32 10.6151
R1902 B.n765 B.n764 10.6151
R1903 B.n764 B.n763 10.6151
R1904 B.n763 B.n34 10.6151
R1905 B.n759 B.n34 10.6151
R1906 B.n759 B.n758 10.6151
R1907 B.n758 B.n757 10.6151
R1908 B.n757 B.n36 10.6151
R1909 B.n753 B.n36 10.6151
R1910 B.n753 B.n752 10.6151
R1911 B.n752 B.n751 10.6151
R1912 B.n751 B.n38 10.6151
R1913 B.n747 B.n38 10.6151
R1914 B.n747 B.n746 10.6151
R1915 B.n746 B.n745 10.6151
R1916 B.n745 B.n40 10.6151
R1917 B.n741 B.n40 10.6151
R1918 B.n741 B.n740 10.6151
R1919 B.n740 B.n739 10.6151
R1920 B.n739 B.n42 10.6151
R1921 B.n735 B.n42 10.6151
R1922 B.n735 B.n734 10.6151
R1923 B.n734 B.n733 10.6151
R1924 B.n733 B.n44 10.6151
R1925 B.n729 B.n44 10.6151
R1926 B.n729 B.n728 10.6151
R1927 B.n728 B.n727 10.6151
R1928 B.n727 B.n46 10.6151
R1929 B.n723 B.n46 10.6151
R1930 B.n723 B.n722 10.6151
R1931 B.n722 B.n721 10.6151
R1932 B.n721 B.n48 10.6151
R1933 B.n717 B.n48 10.6151
R1934 B.n717 B.n716 10.6151
R1935 B.n716 B.n715 10.6151
R1936 B.n715 B.n50 10.6151
R1937 B.n711 B.n50 10.6151
R1938 B.n711 B.n710 10.6151
R1939 B.n710 B.n709 10.6151
R1940 B.n709 B.n52 10.6151
R1941 B.n705 B.n704 10.6151
R1942 B.n704 B.n703 10.6151
R1943 B.n703 B.n57 10.6151
R1944 B.n699 B.n57 10.6151
R1945 B.n699 B.n698 10.6151
R1946 B.n698 B.n697 10.6151
R1947 B.n697 B.n59 10.6151
R1948 B.n693 B.n59 10.6151
R1949 B.n691 B.n690 10.6151
R1950 B.n690 B.n63 10.6151
R1951 B.n686 B.n63 10.6151
R1952 B.n686 B.n685 10.6151
R1953 B.n685 B.n684 10.6151
R1954 B.n684 B.n65 10.6151
R1955 B.n680 B.n65 10.6151
R1956 B.n680 B.n679 10.6151
R1957 B.n679 B.n678 10.6151
R1958 B.n678 B.n67 10.6151
R1959 B.n674 B.n67 10.6151
R1960 B.n674 B.n673 10.6151
R1961 B.n673 B.n672 10.6151
R1962 B.n672 B.n69 10.6151
R1963 B.n668 B.n69 10.6151
R1964 B.n668 B.n667 10.6151
R1965 B.n667 B.n666 10.6151
R1966 B.n666 B.n71 10.6151
R1967 B.n662 B.n71 10.6151
R1968 B.n662 B.n661 10.6151
R1969 B.n661 B.n660 10.6151
R1970 B.n660 B.n73 10.6151
R1971 B.n656 B.n73 10.6151
R1972 B.n656 B.n655 10.6151
R1973 B.n655 B.n654 10.6151
R1974 B.n654 B.n75 10.6151
R1975 B.n650 B.n75 10.6151
R1976 B.n650 B.n649 10.6151
R1977 B.n649 B.n648 10.6151
R1978 B.n648 B.n77 10.6151
R1979 B.n644 B.n77 10.6151
R1980 B.n644 B.n643 10.6151
R1981 B.n643 B.n642 10.6151
R1982 B.n642 B.n79 10.6151
R1983 B.n638 B.n79 10.6151
R1984 B.n638 B.n637 10.6151
R1985 B.n637 B.n636 10.6151
R1986 B.n636 B.n81 10.6151
R1987 B.n632 B.n81 10.6151
R1988 B.n632 B.n631 10.6151
R1989 B.n631 B.n630 10.6151
R1990 B.n630 B.n83 10.6151
R1991 B.n626 B.n83 10.6151
R1992 B.n626 B.n625 10.6151
R1993 B.n625 B.n624 10.6151
R1994 B.n458 B.n457 10.6151
R1995 B.n458 B.n139 10.6151
R1996 B.n462 B.n139 10.6151
R1997 B.n463 B.n462 10.6151
R1998 B.n464 B.n463 10.6151
R1999 B.n464 B.n137 10.6151
R2000 B.n468 B.n137 10.6151
R2001 B.n469 B.n468 10.6151
R2002 B.n470 B.n469 10.6151
R2003 B.n470 B.n135 10.6151
R2004 B.n474 B.n135 10.6151
R2005 B.n475 B.n474 10.6151
R2006 B.n476 B.n475 10.6151
R2007 B.n476 B.n133 10.6151
R2008 B.n480 B.n133 10.6151
R2009 B.n481 B.n480 10.6151
R2010 B.n482 B.n481 10.6151
R2011 B.n482 B.n131 10.6151
R2012 B.n486 B.n131 10.6151
R2013 B.n487 B.n486 10.6151
R2014 B.n488 B.n487 10.6151
R2015 B.n488 B.n129 10.6151
R2016 B.n492 B.n129 10.6151
R2017 B.n493 B.n492 10.6151
R2018 B.n494 B.n493 10.6151
R2019 B.n494 B.n127 10.6151
R2020 B.n498 B.n127 10.6151
R2021 B.n499 B.n498 10.6151
R2022 B.n500 B.n499 10.6151
R2023 B.n500 B.n125 10.6151
R2024 B.n504 B.n125 10.6151
R2025 B.n505 B.n504 10.6151
R2026 B.n506 B.n505 10.6151
R2027 B.n506 B.n123 10.6151
R2028 B.n510 B.n123 10.6151
R2029 B.n511 B.n510 10.6151
R2030 B.n512 B.n511 10.6151
R2031 B.n512 B.n121 10.6151
R2032 B.n516 B.n121 10.6151
R2033 B.n517 B.n516 10.6151
R2034 B.n518 B.n517 10.6151
R2035 B.n518 B.n119 10.6151
R2036 B.n522 B.n119 10.6151
R2037 B.n523 B.n522 10.6151
R2038 B.n524 B.n523 10.6151
R2039 B.n524 B.n117 10.6151
R2040 B.n528 B.n117 10.6151
R2041 B.n529 B.n528 10.6151
R2042 B.n530 B.n529 10.6151
R2043 B.n530 B.n115 10.6151
R2044 B.n534 B.n115 10.6151
R2045 B.n535 B.n534 10.6151
R2046 B.n536 B.n535 10.6151
R2047 B.n536 B.n113 10.6151
R2048 B.n540 B.n113 10.6151
R2049 B.n541 B.n540 10.6151
R2050 B.n542 B.n541 10.6151
R2051 B.n542 B.n111 10.6151
R2052 B.n546 B.n111 10.6151
R2053 B.n547 B.n546 10.6151
R2054 B.n548 B.n547 10.6151
R2055 B.n548 B.n109 10.6151
R2056 B.n552 B.n109 10.6151
R2057 B.n553 B.n552 10.6151
R2058 B.n554 B.n553 10.6151
R2059 B.n554 B.n107 10.6151
R2060 B.n558 B.n107 10.6151
R2061 B.n559 B.n558 10.6151
R2062 B.n560 B.n559 10.6151
R2063 B.n560 B.n105 10.6151
R2064 B.n564 B.n105 10.6151
R2065 B.n565 B.n564 10.6151
R2066 B.n566 B.n565 10.6151
R2067 B.n566 B.n103 10.6151
R2068 B.n570 B.n103 10.6151
R2069 B.n571 B.n570 10.6151
R2070 B.n572 B.n571 10.6151
R2071 B.n572 B.n101 10.6151
R2072 B.n576 B.n101 10.6151
R2073 B.n577 B.n576 10.6151
R2074 B.n578 B.n577 10.6151
R2075 B.n578 B.n99 10.6151
R2076 B.n582 B.n99 10.6151
R2077 B.n583 B.n582 10.6151
R2078 B.n584 B.n583 10.6151
R2079 B.n584 B.n97 10.6151
R2080 B.n588 B.n97 10.6151
R2081 B.n589 B.n588 10.6151
R2082 B.n590 B.n589 10.6151
R2083 B.n590 B.n95 10.6151
R2084 B.n594 B.n95 10.6151
R2085 B.n595 B.n594 10.6151
R2086 B.n596 B.n595 10.6151
R2087 B.n596 B.n93 10.6151
R2088 B.n600 B.n93 10.6151
R2089 B.n601 B.n600 10.6151
R2090 B.n602 B.n601 10.6151
R2091 B.n602 B.n91 10.6151
R2092 B.n606 B.n91 10.6151
R2093 B.n607 B.n606 10.6151
R2094 B.n608 B.n607 10.6151
R2095 B.n608 B.n89 10.6151
R2096 B.n612 B.n89 10.6151
R2097 B.n613 B.n612 10.6151
R2098 B.n614 B.n613 10.6151
R2099 B.n614 B.n87 10.6151
R2100 B.n618 B.n87 10.6151
R2101 B.n619 B.n618 10.6151
R2102 B.n620 B.n619 10.6151
R2103 B.n620 B.n85 10.6151
R2104 B.n303 B.n302 10.6151
R2105 B.n304 B.n303 10.6151
R2106 B.n304 B.n191 10.6151
R2107 B.n308 B.n191 10.6151
R2108 B.n309 B.n308 10.6151
R2109 B.n310 B.n309 10.6151
R2110 B.n310 B.n189 10.6151
R2111 B.n314 B.n189 10.6151
R2112 B.n315 B.n314 10.6151
R2113 B.n316 B.n315 10.6151
R2114 B.n316 B.n187 10.6151
R2115 B.n320 B.n187 10.6151
R2116 B.n321 B.n320 10.6151
R2117 B.n322 B.n321 10.6151
R2118 B.n322 B.n185 10.6151
R2119 B.n326 B.n185 10.6151
R2120 B.n327 B.n326 10.6151
R2121 B.n328 B.n327 10.6151
R2122 B.n328 B.n183 10.6151
R2123 B.n332 B.n183 10.6151
R2124 B.n333 B.n332 10.6151
R2125 B.n334 B.n333 10.6151
R2126 B.n334 B.n181 10.6151
R2127 B.n338 B.n181 10.6151
R2128 B.n339 B.n338 10.6151
R2129 B.n340 B.n339 10.6151
R2130 B.n340 B.n179 10.6151
R2131 B.n344 B.n179 10.6151
R2132 B.n345 B.n344 10.6151
R2133 B.n346 B.n345 10.6151
R2134 B.n346 B.n177 10.6151
R2135 B.n350 B.n177 10.6151
R2136 B.n351 B.n350 10.6151
R2137 B.n352 B.n351 10.6151
R2138 B.n352 B.n175 10.6151
R2139 B.n356 B.n175 10.6151
R2140 B.n357 B.n356 10.6151
R2141 B.n358 B.n357 10.6151
R2142 B.n358 B.n173 10.6151
R2143 B.n362 B.n173 10.6151
R2144 B.n363 B.n362 10.6151
R2145 B.n364 B.n363 10.6151
R2146 B.n364 B.n171 10.6151
R2147 B.n368 B.n171 10.6151
R2148 B.n369 B.n368 10.6151
R2149 B.n371 B.n167 10.6151
R2150 B.n375 B.n167 10.6151
R2151 B.n376 B.n375 10.6151
R2152 B.n377 B.n376 10.6151
R2153 B.n377 B.n165 10.6151
R2154 B.n381 B.n165 10.6151
R2155 B.n382 B.n381 10.6151
R2156 B.n386 B.n382 10.6151
R2157 B.n390 B.n163 10.6151
R2158 B.n391 B.n390 10.6151
R2159 B.n392 B.n391 10.6151
R2160 B.n392 B.n161 10.6151
R2161 B.n396 B.n161 10.6151
R2162 B.n397 B.n396 10.6151
R2163 B.n398 B.n397 10.6151
R2164 B.n398 B.n159 10.6151
R2165 B.n402 B.n159 10.6151
R2166 B.n403 B.n402 10.6151
R2167 B.n404 B.n403 10.6151
R2168 B.n404 B.n157 10.6151
R2169 B.n408 B.n157 10.6151
R2170 B.n409 B.n408 10.6151
R2171 B.n410 B.n409 10.6151
R2172 B.n410 B.n155 10.6151
R2173 B.n414 B.n155 10.6151
R2174 B.n415 B.n414 10.6151
R2175 B.n416 B.n415 10.6151
R2176 B.n416 B.n153 10.6151
R2177 B.n420 B.n153 10.6151
R2178 B.n421 B.n420 10.6151
R2179 B.n422 B.n421 10.6151
R2180 B.n422 B.n151 10.6151
R2181 B.n426 B.n151 10.6151
R2182 B.n427 B.n426 10.6151
R2183 B.n428 B.n427 10.6151
R2184 B.n428 B.n149 10.6151
R2185 B.n432 B.n149 10.6151
R2186 B.n433 B.n432 10.6151
R2187 B.n434 B.n433 10.6151
R2188 B.n434 B.n147 10.6151
R2189 B.n438 B.n147 10.6151
R2190 B.n439 B.n438 10.6151
R2191 B.n440 B.n439 10.6151
R2192 B.n440 B.n145 10.6151
R2193 B.n444 B.n145 10.6151
R2194 B.n445 B.n444 10.6151
R2195 B.n446 B.n445 10.6151
R2196 B.n446 B.n143 10.6151
R2197 B.n450 B.n143 10.6151
R2198 B.n451 B.n450 10.6151
R2199 B.n452 B.n451 10.6151
R2200 B.n452 B.n141 10.6151
R2201 B.n456 B.n141 10.6151
R2202 B.n298 B.n193 10.6151
R2203 B.n298 B.n297 10.6151
R2204 B.n297 B.n296 10.6151
R2205 B.n296 B.n195 10.6151
R2206 B.n292 B.n195 10.6151
R2207 B.n292 B.n291 10.6151
R2208 B.n291 B.n290 10.6151
R2209 B.n290 B.n197 10.6151
R2210 B.n286 B.n197 10.6151
R2211 B.n286 B.n285 10.6151
R2212 B.n285 B.n284 10.6151
R2213 B.n284 B.n199 10.6151
R2214 B.n280 B.n199 10.6151
R2215 B.n280 B.n279 10.6151
R2216 B.n279 B.n278 10.6151
R2217 B.n278 B.n201 10.6151
R2218 B.n274 B.n201 10.6151
R2219 B.n274 B.n273 10.6151
R2220 B.n273 B.n272 10.6151
R2221 B.n272 B.n203 10.6151
R2222 B.n268 B.n203 10.6151
R2223 B.n268 B.n267 10.6151
R2224 B.n267 B.n266 10.6151
R2225 B.n266 B.n205 10.6151
R2226 B.n262 B.n205 10.6151
R2227 B.n262 B.n261 10.6151
R2228 B.n261 B.n260 10.6151
R2229 B.n260 B.n207 10.6151
R2230 B.n256 B.n207 10.6151
R2231 B.n256 B.n255 10.6151
R2232 B.n255 B.n254 10.6151
R2233 B.n254 B.n209 10.6151
R2234 B.n250 B.n209 10.6151
R2235 B.n250 B.n249 10.6151
R2236 B.n249 B.n248 10.6151
R2237 B.n248 B.n211 10.6151
R2238 B.n244 B.n211 10.6151
R2239 B.n244 B.n243 10.6151
R2240 B.n243 B.n242 10.6151
R2241 B.n242 B.n213 10.6151
R2242 B.n238 B.n213 10.6151
R2243 B.n238 B.n237 10.6151
R2244 B.n237 B.n236 10.6151
R2245 B.n236 B.n215 10.6151
R2246 B.n232 B.n215 10.6151
R2247 B.n232 B.n231 10.6151
R2248 B.n231 B.n230 10.6151
R2249 B.n230 B.n217 10.6151
R2250 B.n226 B.n217 10.6151
R2251 B.n226 B.n225 10.6151
R2252 B.n225 B.n224 10.6151
R2253 B.n224 B.n219 10.6151
R2254 B.n220 B.n219 10.6151
R2255 B.n220 B.n0 10.6151
R2256 B.n855 B.n1 10.6151
R2257 B.n855 B.n854 10.6151
R2258 B.n854 B.n853 10.6151
R2259 B.n853 B.n4 10.6151
R2260 B.n849 B.n4 10.6151
R2261 B.n849 B.n848 10.6151
R2262 B.n848 B.n847 10.6151
R2263 B.n847 B.n6 10.6151
R2264 B.n843 B.n6 10.6151
R2265 B.n843 B.n842 10.6151
R2266 B.n842 B.n841 10.6151
R2267 B.n841 B.n8 10.6151
R2268 B.n837 B.n8 10.6151
R2269 B.n837 B.n836 10.6151
R2270 B.n836 B.n835 10.6151
R2271 B.n835 B.n10 10.6151
R2272 B.n831 B.n10 10.6151
R2273 B.n831 B.n830 10.6151
R2274 B.n830 B.n829 10.6151
R2275 B.n829 B.n12 10.6151
R2276 B.n825 B.n12 10.6151
R2277 B.n825 B.n824 10.6151
R2278 B.n824 B.n823 10.6151
R2279 B.n823 B.n14 10.6151
R2280 B.n819 B.n14 10.6151
R2281 B.n819 B.n818 10.6151
R2282 B.n818 B.n817 10.6151
R2283 B.n817 B.n16 10.6151
R2284 B.n813 B.n16 10.6151
R2285 B.n813 B.n812 10.6151
R2286 B.n812 B.n811 10.6151
R2287 B.n811 B.n18 10.6151
R2288 B.n807 B.n18 10.6151
R2289 B.n807 B.n806 10.6151
R2290 B.n806 B.n805 10.6151
R2291 B.n805 B.n20 10.6151
R2292 B.n801 B.n20 10.6151
R2293 B.n801 B.n800 10.6151
R2294 B.n800 B.n799 10.6151
R2295 B.n799 B.n22 10.6151
R2296 B.n795 B.n22 10.6151
R2297 B.n795 B.n794 10.6151
R2298 B.n794 B.n793 10.6151
R2299 B.n793 B.n24 10.6151
R2300 B.n789 B.n24 10.6151
R2301 B.n789 B.n788 10.6151
R2302 B.n788 B.n787 10.6151
R2303 B.n787 B.n26 10.6151
R2304 B.n783 B.n26 10.6151
R2305 B.n783 B.n782 10.6151
R2306 B.n782 B.n781 10.6151
R2307 B.n781 B.n28 10.6151
R2308 B.n777 B.n28 10.6151
R2309 B.n777 B.n776 10.6151
R2310 B.n705 B.n56 6.5566
R2311 B.n693 B.n692 6.5566
R2312 B.n371 B.n370 6.5566
R2313 B.n386 B.n385 6.5566
R2314 B.n56 B.n52 4.05904
R2315 B.n692 B.n691 4.05904
R2316 B.n370 B.n369 4.05904
R2317 B.n385 B.n163 4.05904
R2318 B.n859 B.n0 2.81026
R2319 B.n859 B.n1 2.81026
R2320 VN.n59 VN.n31 161.3
R2321 VN.n58 VN.n57 161.3
R2322 VN.n56 VN.n32 161.3
R2323 VN.n55 VN.n54 161.3
R2324 VN.n53 VN.n33 161.3
R2325 VN.n52 VN.n51 161.3
R2326 VN.n50 VN.n34 161.3
R2327 VN.n49 VN.n48 161.3
R2328 VN.n47 VN.n35 161.3
R2329 VN.n46 VN.n45 161.3
R2330 VN.n44 VN.n37 161.3
R2331 VN.n43 VN.n42 161.3
R2332 VN.n41 VN.n38 161.3
R2333 VN.n28 VN.n0 161.3
R2334 VN.n27 VN.n26 161.3
R2335 VN.n25 VN.n1 161.3
R2336 VN.n24 VN.n23 161.3
R2337 VN.n22 VN.n2 161.3
R2338 VN.n21 VN.n20 161.3
R2339 VN.n19 VN.n3 161.3
R2340 VN.n18 VN.n17 161.3
R2341 VN.n15 VN.n4 161.3
R2342 VN.n14 VN.n13 161.3
R2343 VN.n12 VN.n5 161.3
R2344 VN.n11 VN.n10 161.3
R2345 VN.n9 VN.n6 161.3
R2346 VN.n7 VN.t3 145.733
R2347 VN.n39 VN.t4 145.733
R2348 VN.n8 VN.t6 112.692
R2349 VN.n16 VN.t2 112.692
R2350 VN.n29 VN.t7 112.692
R2351 VN.n40 VN.t5 112.692
R2352 VN.n36 VN.t1 112.692
R2353 VN.n60 VN.t0 112.692
R2354 VN.n30 VN.n29 108.45
R2355 VN.n61 VN.n60 108.45
R2356 VN.n8 VN.n7 56.7106
R2357 VN.n40 VN.n39 56.7106
R2358 VN.n14 VN.n5 56.5617
R2359 VN.n46 VN.n37 56.5617
R2360 VN VN.n61 53.483
R2361 VN.n23 VN.n22 45.4209
R2362 VN.n54 VN.n53 45.4209
R2363 VN.n23 VN.n1 35.7332
R2364 VN.n54 VN.n32 35.7332
R2365 VN.n10 VN.n9 24.5923
R2366 VN.n10 VN.n5 24.5923
R2367 VN.n15 VN.n14 24.5923
R2368 VN.n17 VN.n15 24.5923
R2369 VN.n21 VN.n3 24.5923
R2370 VN.n22 VN.n21 24.5923
R2371 VN.n27 VN.n1 24.5923
R2372 VN.n28 VN.n27 24.5923
R2373 VN.n42 VN.n37 24.5923
R2374 VN.n42 VN.n41 24.5923
R2375 VN.n53 VN.n52 24.5923
R2376 VN.n52 VN.n34 24.5923
R2377 VN.n48 VN.n47 24.5923
R2378 VN.n47 VN.n46 24.5923
R2379 VN.n59 VN.n58 24.5923
R2380 VN.n58 VN.n32 24.5923
R2381 VN.n9 VN.n8 17.2148
R2382 VN.n17 VN.n16 17.2148
R2383 VN.n41 VN.n40 17.2148
R2384 VN.n48 VN.n36 17.2148
R2385 VN.n16 VN.n3 7.37805
R2386 VN.n36 VN.n34 7.37805
R2387 VN.n39 VN.n38 5.07592
R2388 VN.n7 VN.n6 5.07592
R2389 VN.n29 VN.n28 2.45968
R2390 VN.n60 VN.n59 2.45968
R2391 VN.n61 VN.n31 0.278335
R2392 VN.n30 VN.n0 0.278335
R2393 VN.n57 VN.n31 0.189894
R2394 VN.n57 VN.n56 0.189894
R2395 VN.n56 VN.n55 0.189894
R2396 VN.n55 VN.n33 0.189894
R2397 VN.n51 VN.n33 0.189894
R2398 VN.n51 VN.n50 0.189894
R2399 VN.n50 VN.n49 0.189894
R2400 VN.n49 VN.n35 0.189894
R2401 VN.n45 VN.n35 0.189894
R2402 VN.n45 VN.n44 0.189894
R2403 VN.n44 VN.n43 0.189894
R2404 VN.n43 VN.n38 0.189894
R2405 VN.n11 VN.n6 0.189894
R2406 VN.n12 VN.n11 0.189894
R2407 VN.n13 VN.n12 0.189894
R2408 VN.n13 VN.n4 0.189894
R2409 VN.n18 VN.n4 0.189894
R2410 VN.n19 VN.n18 0.189894
R2411 VN.n20 VN.n19 0.189894
R2412 VN.n20 VN.n2 0.189894
R2413 VN.n24 VN.n2 0.189894
R2414 VN.n25 VN.n24 0.189894
R2415 VN.n26 VN.n25 0.189894
R2416 VN.n26 VN.n0 0.189894
R2417 VN VN.n30 0.153485
R2418 VDD2.n2 VDD2.n1 77.557
R2419 VDD2.n2 VDD2.n0 77.557
R2420 VDD2 VDD2.n5 77.5542
R2421 VDD2.n4 VDD2.n3 76.2332
R2422 VDD2.n4 VDD2.n2 47.6981
R2423 VDD2.n5 VDD2.t2 2.42263
R2424 VDD2.n5 VDD2.t3 2.42263
R2425 VDD2.n3 VDD2.t7 2.42263
R2426 VDD2.n3 VDD2.t6 2.42263
R2427 VDD2.n1 VDD2.t5 2.42263
R2428 VDD2.n1 VDD2.t0 2.42263
R2429 VDD2.n0 VDD2.t4 2.42263
R2430 VDD2.n0 VDD2.t1 2.42263
R2431 VDD2 VDD2.n4 1.438
C0 VDD2 B 1.87376f
C1 VTAIL B 5.57638f
C2 VN VDD1 0.152241f
C3 w_n4170_n3652# VP 9.11901f
C4 VN VDD2 9.85667f
C5 VN VTAIL 10.2722f
C6 VDD1 VDD2 1.91584f
C7 VTAIL VDD1 8.59979f
C8 B VP 2.219f
C9 w_n4170_n3652# B 10.9273f
C10 VTAIL VDD2 8.656019f
C11 VN VP 8.249081f
C12 w_n4170_n3652# VN 8.57686f
C13 VDD1 VP 10.2513f
C14 w_n4170_n3652# VDD1 2.07548f
C15 VDD2 VP 0.548426f
C16 VTAIL VP 10.2863f
C17 w_n4170_n3652# VDD2 2.20151f
C18 VN B 1.30873f
C19 w_n4170_n3652# VTAIL 4.55192f
C20 VDD1 B 1.76924f
C21 VDD2 VSUBS 1.990705f
C22 VDD1 VSUBS 2.68317f
C23 VTAIL VSUBS 1.447601f
C24 VN VSUBS 7.13236f
C25 VP VSUBS 3.906621f
C26 B VSUBS 5.426089f
C27 w_n4170_n3652# VSUBS 0.1871p
C28 VDD2.t4 VSUBS 0.288605f
C29 VDD2.t1 VSUBS 0.288605f
C30 VDD2.n0 VSUBS 2.33518f
C31 VDD2.t5 VSUBS 0.288605f
C32 VDD2.t0 VSUBS 0.288605f
C33 VDD2.n1 VSUBS 2.33518f
C34 VDD2.n2 VSUBS 4.37253f
C35 VDD2.t7 VSUBS 0.288605f
C36 VDD2.t6 VSUBS 0.288605f
C37 VDD2.n3 VSUBS 2.32043f
C38 VDD2.n4 VSUBS 3.70185f
C39 VDD2.t2 VSUBS 0.288605f
C40 VDD2.t3 VSUBS 0.288605f
C41 VDD2.n5 VSUBS 2.33513f
C42 VN.n0 VSUBS 0.035225f
C43 VN.t7 VSUBS 2.81245f
C44 VN.n1 VSUBS 0.053668f
C45 VN.n2 VSUBS 0.02672f
C46 VN.n3 VSUBS 0.032426f
C47 VN.n4 VSUBS 0.02672f
C48 VN.n5 VSUBS 0.038841f
C49 VN.n6 VSUBS 0.282461f
C50 VN.t6 VSUBS 2.81245f
C51 VN.t3 VSUBS 3.07671f
C52 VN.n7 VSUBS 1.03254f
C53 VN.n8 VSUBS 1.07326f
C54 VN.n9 VSUBS 0.042211f
C55 VN.n10 VSUBS 0.049549f
C56 VN.n11 VSUBS 0.02672f
C57 VN.n12 VSUBS 0.02672f
C58 VN.n13 VSUBS 0.02672f
C59 VN.n14 VSUBS 0.038841f
C60 VN.n15 VSUBS 0.049549f
C61 VN.t2 VSUBS 2.81245f
C62 VN.n16 VSUBS 0.985822f
C63 VN.n17 VSUBS 0.042211f
C64 VN.n18 VSUBS 0.02672f
C65 VN.n19 VSUBS 0.02672f
C66 VN.n20 VSUBS 0.02672f
C67 VN.n21 VSUBS 0.049549f
C68 VN.n22 VSUBS 0.05112f
C69 VN.n23 VSUBS 0.022444f
C70 VN.n24 VSUBS 0.02672f
C71 VN.n25 VSUBS 0.02672f
C72 VN.n26 VSUBS 0.02672f
C73 VN.n27 VSUBS 0.049549f
C74 VN.n28 VSUBS 0.027534f
C75 VN.n29 VSUBS 1.07341f
C76 VN.n30 VSUBS 0.050803f
C77 VN.n31 VSUBS 0.035225f
C78 VN.t0 VSUBS 2.81245f
C79 VN.n32 VSUBS 0.053668f
C80 VN.n33 VSUBS 0.02672f
C81 VN.n34 VSUBS 0.032426f
C82 VN.n35 VSUBS 0.02672f
C83 VN.t1 VSUBS 2.81245f
C84 VN.n36 VSUBS 0.985822f
C85 VN.n37 VSUBS 0.038841f
C86 VN.n38 VSUBS 0.282461f
C87 VN.t5 VSUBS 2.81245f
C88 VN.t4 VSUBS 3.07671f
C89 VN.n39 VSUBS 1.03254f
C90 VN.n40 VSUBS 1.07326f
C91 VN.n41 VSUBS 0.042211f
C92 VN.n42 VSUBS 0.049549f
C93 VN.n43 VSUBS 0.02672f
C94 VN.n44 VSUBS 0.02672f
C95 VN.n45 VSUBS 0.02672f
C96 VN.n46 VSUBS 0.038841f
C97 VN.n47 VSUBS 0.049549f
C98 VN.n48 VSUBS 0.042211f
C99 VN.n49 VSUBS 0.02672f
C100 VN.n50 VSUBS 0.02672f
C101 VN.n51 VSUBS 0.02672f
C102 VN.n52 VSUBS 0.049549f
C103 VN.n53 VSUBS 0.05112f
C104 VN.n54 VSUBS 0.022444f
C105 VN.n55 VSUBS 0.02672f
C106 VN.n56 VSUBS 0.02672f
C107 VN.n57 VSUBS 0.02672f
C108 VN.n58 VSUBS 0.049549f
C109 VN.n59 VSUBS 0.027534f
C110 VN.n60 VSUBS 1.07341f
C111 VN.n61 VSUBS 1.6482f
C112 B.n0 VSUBS 0.004571f
C113 B.n1 VSUBS 0.004571f
C114 B.n2 VSUBS 0.007228f
C115 B.n3 VSUBS 0.007228f
C116 B.n4 VSUBS 0.007228f
C117 B.n5 VSUBS 0.007228f
C118 B.n6 VSUBS 0.007228f
C119 B.n7 VSUBS 0.007228f
C120 B.n8 VSUBS 0.007228f
C121 B.n9 VSUBS 0.007228f
C122 B.n10 VSUBS 0.007228f
C123 B.n11 VSUBS 0.007228f
C124 B.n12 VSUBS 0.007228f
C125 B.n13 VSUBS 0.007228f
C126 B.n14 VSUBS 0.007228f
C127 B.n15 VSUBS 0.007228f
C128 B.n16 VSUBS 0.007228f
C129 B.n17 VSUBS 0.007228f
C130 B.n18 VSUBS 0.007228f
C131 B.n19 VSUBS 0.007228f
C132 B.n20 VSUBS 0.007228f
C133 B.n21 VSUBS 0.007228f
C134 B.n22 VSUBS 0.007228f
C135 B.n23 VSUBS 0.007228f
C136 B.n24 VSUBS 0.007228f
C137 B.n25 VSUBS 0.007228f
C138 B.n26 VSUBS 0.007228f
C139 B.n27 VSUBS 0.007228f
C140 B.n28 VSUBS 0.007228f
C141 B.n29 VSUBS 0.017316f
C142 B.n30 VSUBS 0.007228f
C143 B.n31 VSUBS 0.007228f
C144 B.n32 VSUBS 0.007228f
C145 B.n33 VSUBS 0.007228f
C146 B.n34 VSUBS 0.007228f
C147 B.n35 VSUBS 0.007228f
C148 B.n36 VSUBS 0.007228f
C149 B.n37 VSUBS 0.007228f
C150 B.n38 VSUBS 0.007228f
C151 B.n39 VSUBS 0.007228f
C152 B.n40 VSUBS 0.007228f
C153 B.n41 VSUBS 0.007228f
C154 B.n42 VSUBS 0.007228f
C155 B.n43 VSUBS 0.007228f
C156 B.n44 VSUBS 0.007228f
C157 B.n45 VSUBS 0.007228f
C158 B.n46 VSUBS 0.007228f
C159 B.n47 VSUBS 0.007228f
C160 B.n48 VSUBS 0.007228f
C161 B.n49 VSUBS 0.007228f
C162 B.n50 VSUBS 0.007228f
C163 B.n51 VSUBS 0.007228f
C164 B.n52 VSUBS 0.004996f
C165 B.n53 VSUBS 0.007228f
C166 B.t2 VSUBS 0.250972f
C167 B.t1 VSUBS 0.287257f
C168 B.t0 VSUBS 1.81109f
C169 B.n54 VSUBS 0.453645f
C170 B.n55 VSUBS 0.281155f
C171 B.n56 VSUBS 0.016747f
C172 B.n57 VSUBS 0.007228f
C173 B.n58 VSUBS 0.007228f
C174 B.n59 VSUBS 0.007228f
C175 B.n60 VSUBS 0.007228f
C176 B.t8 VSUBS 0.250976f
C177 B.t7 VSUBS 0.28726f
C178 B.t6 VSUBS 1.81109f
C179 B.n61 VSUBS 0.453642f
C180 B.n62 VSUBS 0.281152f
C181 B.n63 VSUBS 0.007228f
C182 B.n64 VSUBS 0.007228f
C183 B.n65 VSUBS 0.007228f
C184 B.n66 VSUBS 0.007228f
C185 B.n67 VSUBS 0.007228f
C186 B.n68 VSUBS 0.007228f
C187 B.n69 VSUBS 0.007228f
C188 B.n70 VSUBS 0.007228f
C189 B.n71 VSUBS 0.007228f
C190 B.n72 VSUBS 0.007228f
C191 B.n73 VSUBS 0.007228f
C192 B.n74 VSUBS 0.007228f
C193 B.n75 VSUBS 0.007228f
C194 B.n76 VSUBS 0.007228f
C195 B.n77 VSUBS 0.007228f
C196 B.n78 VSUBS 0.007228f
C197 B.n79 VSUBS 0.007228f
C198 B.n80 VSUBS 0.007228f
C199 B.n81 VSUBS 0.007228f
C200 B.n82 VSUBS 0.007228f
C201 B.n83 VSUBS 0.007228f
C202 B.n84 VSUBS 0.007228f
C203 B.n85 VSUBS 0.01811f
C204 B.n86 VSUBS 0.007228f
C205 B.n87 VSUBS 0.007228f
C206 B.n88 VSUBS 0.007228f
C207 B.n89 VSUBS 0.007228f
C208 B.n90 VSUBS 0.007228f
C209 B.n91 VSUBS 0.007228f
C210 B.n92 VSUBS 0.007228f
C211 B.n93 VSUBS 0.007228f
C212 B.n94 VSUBS 0.007228f
C213 B.n95 VSUBS 0.007228f
C214 B.n96 VSUBS 0.007228f
C215 B.n97 VSUBS 0.007228f
C216 B.n98 VSUBS 0.007228f
C217 B.n99 VSUBS 0.007228f
C218 B.n100 VSUBS 0.007228f
C219 B.n101 VSUBS 0.007228f
C220 B.n102 VSUBS 0.007228f
C221 B.n103 VSUBS 0.007228f
C222 B.n104 VSUBS 0.007228f
C223 B.n105 VSUBS 0.007228f
C224 B.n106 VSUBS 0.007228f
C225 B.n107 VSUBS 0.007228f
C226 B.n108 VSUBS 0.007228f
C227 B.n109 VSUBS 0.007228f
C228 B.n110 VSUBS 0.007228f
C229 B.n111 VSUBS 0.007228f
C230 B.n112 VSUBS 0.007228f
C231 B.n113 VSUBS 0.007228f
C232 B.n114 VSUBS 0.007228f
C233 B.n115 VSUBS 0.007228f
C234 B.n116 VSUBS 0.007228f
C235 B.n117 VSUBS 0.007228f
C236 B.n118 VSUBS 0.007228f
C237 B.n119 VSUBS 0.007228f
C238 B.n120 VSUBS 0.007228f
C239 B.n121 VSUBS 0.007228f
C240 B.n122 VSUBS 0.007228f
C241 B.n123 VSUBS 0.007228f
C242 B.n124 VSUBS 0.007228f
C243 B.n125 VSUBS 0.007228f
C244 B.n126 VSUBS 0.007228f
C245 B.n127 VSUBS 0.007228f
C246 B.n128 VSUBS 0.007228f
C247 B.n129 VSUBS 0.007228f
C248 B.n130 VSUBS 0.007228f
C249 B.n131 VSUBS 0.007228f
C250 B.n132 VSUBS 0.007228f
C251 B.n133 VSUBS 0.007228f
C252 B.n134 VSUBS 0.007228f
C253 B.n135 VSUBS 0.007228f
C254 B.n136 VSUBS 0.007228f
C255 B.n137 VSUBS 0.007228f
C256 B.n138 VSUBS 0.007228f
C257 B.n139 VSUBS 0.007228f
C258 B.n140 VSUBS 0.017316f
C259 B.n141 VSUBS 0.007228f
C260 B.n142 VSUBS 0.007228f
C261 B.n143 VSUBS 0.007228f
C262 B.n144 VSUBS 0.007228f
C263 B.n145 VSUBS 0.007228f
C264 B.n146 VSUBS 0.007228f
C265 B.n147 VSUBS 0.007228f
C266 B.n148 VSUBS 0.007228f
C267 B.n149 VSUBS 0.007228f
C268 B.n150 VSUBS 0.007228f
C269 B.n151 VSUBS 0.007228f
C270 B.n152 VSUBS 0.007228f
C271 B.n153 VSUBS 0.007228f
C272 B.n154 VSUBS 0.007228f
C273 B.n155 VSUBS 0.007228f
C274 B.n156 VSUBS 0.007228f
C275 B.n157 VSUBS 0.007228f
C276 B.n158 VSUBS 0.007228f
C277 B.n159 VSUBS 0.007228f
C278 B.n160 VSUBS 0.007228f
C279 B.n161 VSUBS 0.007228f
C280 B.n162 VSUBS 0.007228f
C281 B.n163 VSUBS 0.004996f
C282 B.n164 VSUBS 0.007228f
C283 B.n165 VSUBS 0.007228f
C284 B.n166 VSUBS 0.007228f
C285 B.n167 VSUBS 0.007228f
C286 B.n168 VSUBS 0.007228f
C287 B.t10 VSUBS 0.250972f
C288 B.t11 VSUBS 0.287257f
C289 B.t9 VSUBS 1.81109f
C290 B.n169 VSUBS 0.453645f
C291 B.n170 VSUBS 0.281155f
C292 B.n171 VSUBS 0.007228f
C293 B.n172 VSUBS 0.007228f
C294 B.n173 VSUBS 0.007228f
C295 B.n174 VSUBS 0.007228f
C296 B.n175 VSUBS 0.007228f
C297 B.n176 VSUBS 0.007228f
C298 B.n177 VSUBS 0.007228f
C299 B.n178 VSUBS 0.007228f
C300 B.n179 VSUBS 0.007228f
C301 B.n180 VSUBS 0.007228f
C302 B.n181 VSUBS 0.007228f
C303 B.n182 VSUBS 0.007228f
C304 B.n183 VSUBS 0.007228f
C305 B.n184 VSUBS 0.007228f
C306 B.n185 VSUBS 0.007228f
C307 B.n186 VSUBS 0.007228f
C308 B.n187 VSUBS 0.007228f
C309 B.n188 VSUBS 0.007228f
C310 B.n189 VSUBS 0.007228f
C311 B.n190 VSUBS 0.007228f
C312 B.n191 VSUBS 0.007228f
C313 B.n192 VSUBS 0.007228f
C314 B.n193 VSUBS 0.017316f
C315 B.n194 VSUBS 0.007228f
C316 B.n195 VSUBS 0.007228f
C317 B.n196 VSUBS 0.007228f
C318 B.n197 VSUBS 0.007228f
C319 B.n198 VSUBS 0.007228f
C320 B.n199 VSUBS 0.007228f
C321 B.n200 VSUBS 0.007228f
C322 B.n201 VSUBS 0.007228f
C323 B.n202 VSUBS 0.007228f
C324 B.n203 VSUBS 0.007228f
C325 B.n204 VSUBS 0.007228f
C326 B.n205 VSUBS 0.007228f
C327 B.n206 VSUBS 0.007228f
C328 B.n207 VSUBS 0.007228f
C329 B.n208 VSUBS 0.007228f
C330 B.n209 VSUBS 0.007228f
C331 B.n210 VSUBS 0.007228f
C332 B.n211 VSUBS 0.007228f
C333 B.n212 VSUBS 0.007228f
C334 B.n213 VSUBS 0.007228f
C335 B.n214 VSUBS 0.007228f
C336 B.n215 VSUBS 0.007228f
C337 B.n216 VSUBS 0.007228f
C338 B.n217 VSUBS 0.007228f
C339 B.n218 VSUBS 0.007228f
C340 B.n219 VSUBS 0.007228f
C341 B.n220 VSUBS 0.007228f
C342 B.n221 VSUBS 0.007228f
C343 B.n222 VSUBS 0.007228f
C344 B.n223 VSUBS 0.007228f
C345 B.n224 VSUBS 0.007228f
C346 B.n225 VSUBS 0.007228f
C347 B.n226 VSUBS 0.007228f
C348 B.n227 VSUBS 0.007228f
C349 B.n228 VSUBS 0.007228f
C350 B.n229 VSUBS 0.007228f
C351 B.n230 VSUBS 0.007228f
C352 B.n231 VSUBS 0.007228f
C353 B.n232 VSUBS 0.007228f
C354 B.n233 VSUBS 0.007228f
C355 B.n234 VSUBS 0.007228f
C356 B.n235 VSUBS 0.007228f
C357 B.n236 VSUBS 0.007228f
C358 B.n237 VSUBS 0.007228f
C359 B.n238 VSUBS 0.007228f
C360 B.n239 VSUBS 0.007228f
C361 B.n240 VSUBS 0.007228f
C362 B.n241 VSUBS 0.007228f
C363 B.n242 VSUBS 0.007228f
C364 B.n243 VSUBS 0.007228f
C365 B.n244 VSUBS 0.007228f
C366 B.n245 VSUBS 0.007228f
C367 B.n246 VSUBS 0.007228f
C368 B.n247 VSUBS 0.007228f
C369 B.n248 VSUBS 0.007228f
C370 B.n249 VSUBS 0.007228f
C371 B.n250 VSUBS 0.007228f
C372 B.n251 VSUBS 0.007228f
C373 B.n252 VSUBS 0.007228f
C374 B.n253 VSUBS 0.007228f
C375 B.n254 VSUBS 0.007228f
C376 B.n255 VSUBS 0.007228f
C377 B.n256 VSUBS 0.007228f
C378 B.n257 VSUBS 0.007228f
C379 B.n258 VSUBS 0.007228f
C380 B.n259 VSUBS 0.007228f
C381 B.n260 VSUBS 0.007228f
C382 B.n261 VSUBS 0.007228f
C383 B.n262 VSUBS 0.007228f
C384 B.n263 VSUBS 0.007228f
C385 B.n264 VSUBS 0.007228f
C386 B.n265 VSUBS 0.007228f
C387 B.n266 VSUBS 0.007228f
C388 B.n267 VSUBS 0.007228f
C389 B.n268 VSUBS 0.007228f
C390 B.n269 VSUBS 0.007228f
C391 B.n270 VSUBS 0.007228f
C392 B.n271 VSUBS 0.007228f
C393 B.n272 VSUBS 0.007228f
C394 B.n273 VSUBS 0.007228f
C395 B.n274 VSUBS 0.007228f
C396 B.n275 VSUBS 0.007228f
C397 B.n276 VSUBS 0.007228f
C398 B.n277 VSUBS 0.007228f
C399 B.n278 VSUBS 0.007228f
C400 B.n279 VSUBS 0.007228f
C401 B.n280 VSUBS 0.007228f
C402 B.n281 VSUBS 0.007228f
C403 B.n282 VSUBS 0.007228f
C404 B.n283 VSUBS 0.007228f
C405 B.n284 VSUBS 0.007228f
C406 B.n285 VSUBS 0.007228f
C407 B.n286 VSUBS 0.007228f
C408 B.n287 VSUBS 0.007228f
C409 B.n288 VSUBS 0.007228f
C410 B.n289 VSUBS 0.007228f
C411 B.n290 VSUBS 0.007228f
C412 B.n291 VSUBS 0.007228f
C413 B.n292 VSUBS 0.007228f
C414 B.n293 VSUBS 0.007228f
C415 B.n294 VSUBS 0.007228f
C416 B.n295 VSUBS 0.007228f
C417 B.n296 VSUBS 0.007228f
C418 B.n297 VSUBS 0.007228f
C419 B.n298 VSUBS 0.007228f
C420 B.n299 VSUBS 0.007228f
C421 B.n300 VSUBS 0.017316f
C422 B.n301 VSUBS 0.018188f
C423 B.n302 VSUBS 0.018188f
C424 B.n303 VSUBS 0.007228f
C425 B.n304 VSUBS 0.007228f
C426 B.n305 VSUBS 0.007228f
C427 B.n306 VSUBS 0.007228f
C428 B.n307 VSUBS 0.007228f
C429 B.n308 VSUBS 0.007228f
C430 B.n309 VSUBS 0.007228f
C431 B.n310 VSUBS 0.007228f
C432 B.n311 VSUBS 0.007228f
C433 B.n312 VSUBS 0.007228f
C434 B.n313 VSUBS 0.007228f
C435 B.n314 VSUBS 0.007228f
C436 B.n315 VSUBS 0.007228f
C437 B.n316 VSUBS 0.007228f
C438 B.n317 VSUBS 0.007228f
C439 B.n318 VSUBS 0.007228f
C440 B.n319 VSUBS 0.007228f
C441 B.n320 VSUBS 0.007228f
C442 B.n321 VSUBS 0.007228f
C443 B.n322 VSUBS 0.007228f
C444 B.n323 VSUBS 0.007228f
C445 B.n324 VSUBS 0.007228f
C446 B.n325 VSUBS 0.007228f
C447 B.n326 VSUBS 0.007228f
C448 B.n327 VSUBS 0.007228f
C449 B.n328 VSUBS 0.007228f
C450 B.n329 VSUBS 0.007228f
C451 B.n330 VSUBS 0.007228f
C452 B.n331 VSUBS 0.007228f
C453 B.n332 VSUBS 0.007228f
C454 B.n333 VSUBS 0.007228f
C455 B.n334 VSUBS 0.007228f
C456 B.n335 VSUBS 0.007228f
C457 B.n336 VSUBS 0.007228f
C458 B.n337 VSUBS 0.007228f
C459 B.n338 VSUBS 0.007228f
C460 B.n339 VSUBS 0.007228f
C461 B.n340 VSUBS 0.007228f
C462 B.n341 VSUBS 0.007228f
C463 B.n342 VSUBS 0.007228f
C464 B.n343 VSUBS 0.007228f
C465 B.n344 VSUBS 0.007228f
C466 B.n345 VSUBS 0.007228f
C467 B.n346 VSUBS 0.007228f
C468 B.n347 VSUBS 0.007228f
C469 B.n348 VSUBS 0.007228f
C470 B.n349 VSUBS 0.007228f
C471 B.n350 VSUBS 0.007228f
C472 B.n351 VSUBS 0.007228f
C473 B.n352 VSUBS 0.007228f
C474 B.n353 VSUBS 0.007228f
C475 B.n354 VSUBS 0.007228f
C476 B.n355 VSUBS 0.007228f
C477 B.n356 VSUBS 0.007228f
C478 B.n357 VSUBS 0.007228f
C479 B.n358 VSUBS 0.007228f
C480 B.n359 VSUBS 0.007228f
C481 B.n360 VSUBS 0.007228f
C482 B.n361 VSUBS 0.007228f
C483 B.n362 VSUBS 0.007228f
C484 B.n363 VSUBS 0.007228f
C485 B.n364 VSUBS 0.007228f
C486 B.n365 VSUBS 0.007228f
C487 B.n366 VSUBS 0.007228f
C488 B.n367 VSUBS 0.007228f
C489 B.n368 VSUBS 0.007228f
C490 B.n369 VSUBS 0.004996f
C491 B.n370 VSUBS 0.016747f
C492 B.n371 VSUBS 0.005846f
C493 B.n372 VSUBS 0.007228f
C494 B.n373 VSUBS 0.007228f
C495 B.n374 VSUBS 0.007228f
C496 B.n375 VSUBS 0.007228f
C497 B.n376 VSUBS 0.007228f
C498 B.n377 VSUBS 0.007228f
C499 B.n378 VSUBS 0.007228f
C500 B.n379 VSUBS 0.007228f
C501 B.n380 VSUBS 0.007228f
C502 B.n381 VSUBS 0.007228f
C503 B.n382 VSUBS 0.007228f
C504 B.t4 VSUBS 0.250976f
C505 B.t5 VSUBS 0.28726f
C506 B.t3 VSUBS 1.81109f
C507 B.n383 VSUBS 0.453642f
C508 B.n384 VSUBS 0.281152f
C509 B.n385 VSUBS 0.016747f
C510 B.n386 VSUBS 0.005846f
C511 B.n387 VSUBS 0.007228f
C512 B.n388 VSUBS 0.007228f
C513 B.n389 VSUBS 0.007228f
C514 B.n390 VSUBS 0.007228f
C515 B.n391 VSUBS 0.007228f
C516 B.n392 VSUBS 0.007228f
C517 B.n393 VSUBS 0.007228f
C518 B.n394 VSUBS 0.007228f
C519 B.n395 VSUBS 0.007228f
C520 B.n396 VSUBS 0.007228f
C521 B.n397 VSUBS 0.007228f
C522 B.n398 VSUBS 0.007228f
C523 B.n399 VSUBS 0.007228f
C524 B.n400 VSUBS 0.007228f
C525 B.n401 VSUBS 0.007228f
C526 B.n402 VSUBS 0.007228f
C527 B.n403 VSUBS 0.007228f
C528 B.n404 VSUBS 0.007228f
C529 B.n405 VSUBS 0.007228f
C530 B.n406 VSUBS 0.007228f
C531 B.n407 VSUBS 0.007228f
C532 B.n408 VSUBS 0.007228f
C533 B.n409 VSUBS 0.007228f
C534 B.n410 VSUBS 0.007228f
C535 B.n411 VSUBS 0.007228f
C536 B.n412 VSUBS 0.007228f
C537 B.n413 VSUBS 0.007228f
C538 B.n414 VSUBS 0.007228f
C539 B.n415 VSUBS 0.007228f
C540 B.n416 VSUBS 0.007228f
C541 B.n417 VSUBS 0.007228f
C542 B.n418 VSUBS 0.007228f
C543 B.n419 VSUBS 0.007228f
C544 B.n420 VSUBS 0.007228f
C545 B.n421 VSUBS 0.007228f
C546 B.n422 VSUBS 0.007228f
C547 B.n423 VSUBS 0.007228f
C548 B.n424 VSUBS 0.007228f
C549 B.n425 VSUBS 0.007228f
C550 B.n426 VSUBS 0.007228f
C551 B.n427 VSUBS 0.007228f
C552 B.n428 VSUBS 0.007228f
C553 B.n429 VSUBS 0.007228f
C554 B.n430 VSUBS 0.007228f
C555 B.n431 VSUBS 0.007228f
C556 B.n432 VSUBS 0.007228f
C557 B.n433 VSUBS 0.007228f
C558 B.n434 VSUBS 0.007228f
C559 B.n435 VSUBS 0.007228f
C560 B.n436 VSUBS 0.007228f
C561 B.n437 VSUBS 0.007228f
C562 B.n438 VSUBS 0.007228f
C563 B.n439 VSUBS 0.007228f
C564 B.n440 VSUBS 0.007228f
C565 B.n441 VSUBS 0.007228f
C566 B.n442 VSUBS 0.007228f
C567 B.n443 VSUBS 0.007228f
C568 B.n444 VSUBS 0.007228f
C569 B.n445 VSUBS 0.007228f
C570 B.n446 VSUBS 0.007228f
C571 B.n447 VSUBS 0.007228f
C572 B.n448 VSUBS 0.007228f
C573 B.n449 VSUBS 0.007228f
C574 B.n450 VSUBS 0.007228f
C575 B.n451 VSUBS 0.007228f
C576 B.n452 VSUBS 0.007228f
C577 B.n453 VSUBS 0.007228f
C578 B.n454 VSUBS 0.007228f
C579 B.n455 VSUBS 0.018188f
C580 B.n456 VSUBS 0.018188f
C581 B.n457 VSUBS 0.017316f
C582 B.n458 VSUBS 0.007228f
C583 B.n459 VSUBS 0.007228f
C584 B.n460 VSUBS 0.007228f
C585 B.n461 VSUBS 0.007228f
C586 B.n462 VSUBS 0.007228f
C587 B.n463 VSUBS 0.007228f
C588 B.n464 VSUBS 0.007228f
C589 B.n465 VSUBS 0.007228f
C590 B.n466 VSUBS 0.007228f
C591 B.n467 VSUBS 0.007228f
C592 B.n468 VSUBS 0.007228f
C593 B.n469 VSUBS 0.007228f
C594 B.n470 VSUBS 0.007228f
C595 B.n471 VSUBS 0.007228f
C596 B.n472 VSUBS 0.007228f
C597 B.n473 VSUBS 0.007228f
C598 B.n474 VSUBS 0.007228f
C599 B.n475 VSUBS 0.007228f
C600 B.n476 VSUBS 0.007228f
C601 B.n477 VSUBS 0.007228f
C602 B.n478 VSUBS 0.007228f
C603 B.n479 VSUBS 0.007228f
C604 B.n480 VSUBS 0.007228f
C605 B.n481 VSUBS 0.007228f
C606 B.n482 VSUBS 0.007228f
C607 B.n483 VSUBS 0.007228f
C608 B.n484 VSUBS 0.007228f
C609 B.n485 VSUBS 0.007228f
C610 B.n486 VSUBS 0.007228f
C611 B.n487 VSUBS 0.007228f
C612 B.n488 VSUBS 0.007228f
C613 B.n489 VSUBS 0.007228f
C614 B.n490 VSUBS 0.007228f
C615 B.n491 VSUBS 0.007228f
C616 B.n492 VSUBS 0.007228f
C617 B.n493 VSUBS 0.007228f
C618 B.n494 VSUBS 0.007228f
C619 B.n495 VSUBS 0.007228f
C620 B.n496 VSUBS 0.007228f
C621 B.n497 VSUBS 0.007228f
C622 B.n498 VSUBS 0.007228f
C623 B.n499 VSUBS 0.007228f
C624 B.n500 VSUBS 0.007228f
C625 B.n501 VSUBS 0.007228f
C626 B.n502 VSUBS 0.007228f
C627 B.n503 VSUBS 0.007228f
C628 B.n504 VSUBS 0.007228f
C629 B.n505 VSUBS 0.007228f
C630 B.n506 VSUBS 0.007228f
C631 B.n507 VSUBS 0.007228f
C632 B.n508 VSUBS 0.007228f
C633 B.n509 VSUBS 0.007228f
C634 B.n510 VSUBS 0.007228f
C635 B.n511 VSUBS 0.007228f
C636 B.n512 VSUBS 0.007228f
C637 B.n513 VSUBS 0.007228f
C638 B.n514 VSUBS 0.007228f
C639 B.n515 VSUBS 0.007228f
C640 B.n516 VSUBS 0.007228f
C641 B.n517 VSUBS 0.007228f
C642 B.n518 VSUBS 0.007228f
C643 B.n519 VSUBS 0.007228f
C644 B.n520 VSUBS 0.007228f
C645 B.n521 VSUBS 0.007228f
C646 B.n522 VSUBS 0.007228f
C647 B.n523 VSUBS 0.007228f
C648 B.n524 VSUBS 0.007228f
C649 B.n525 VSUBS 0.007228f
C650 B.n526 VSUBS 0.007228f
C651 B.n527 VSUBS 0.007228f
C652 B.n528 VSUBS 0.007228f
C653 B.n529 VSUBS 0.007228f
C654 B.n530 VSUBS 0.007228f
C655 B.n531 VSUBS 0.007228f
C656 B.n532 VSUBS 0.007228f
C657 B.n533 VSUBS 0.007228f
C658 B.n534 VSUBS 0.007228f
C659 B.n535 VSUBS 0.007228f
C660 B.n536 VSUBS 0.007228f
C661 B.n537 VSUBS 0.007228f
C662 B.n538 VSUBS 0.007228f
C663 B.n539 VSUBS 0.007228f
C664 B.n540 VSUBS 0.007228f
C665 B.n541 VSUBS 0.007228f
C666 B.n542 VSUBS 0.007228f
C667 B.n543 VSUBS 0.007228f
C668 B.n544 VSUBS 0.007228f
C669 B.n545 VSUBS 0.007228f
C670 B.n546 VSUBS 0.007228f
C671 B.n547 VSUBS 0.007228f
C672 B.n548 VSUBS 0.007228f
C673 B.n549 VSUBS 0.007228f
C674 B.n550 VSUBS 0.007228f
C675 B.n551 VSUBS 0.007228f
C676 B.n552 VSUBS 0.007228f
C677 B.n553 VSUBS 0.007228f
C678 B.n554 VSUBS 0.007228f
C679 B.n555 VSUBS 0.007228f
C680 B.n556 VSUBS 0.007228f
C681 B.n557 VSUBS 0.007228f
C682 B.n558 VSUBS 0.007228f
C683 B.n559 VSUBS 0.007228f
C684 B.n560 VSUBS 0.007228f
C685 B.n561 VSUBS 0.007228f
C686 B.n562 VSUBS 0.007228f
C687 B.n563 VSUBS 0.007228f
C688 B.n564 VSUBS 0.007228f
C689 B.n565 VSUBS 0.007228f
C690 B.n566 VSUBS 0.007228f
C691 B.n567 VSUBS 0.007228f
C692 B.n568 VSUBS 0.007228f
C693 B.n569 VSUBS 0.007228f
C694 B.n570 VSUBS 0.007228f
C695 B.n571 VSUBS 0.007228f
C696 B.n572 VSUBS 0.007228f
C697 B.n573 VSUBS 0.007228f
C698 B.n574 VSUBS 0.007228f
C699 B.n575 VSUBS 0.007228f
C700 B.n576 VSUBS 0.007228f
C701 B.n577 VSUBS 0.007228f
C702 B.n578 VSUBS 0.007228f
C703 B.n579 VSUBS 0.007228f
C704 B.n580 VSUBS 0.007228f
C705 B.n581 VSUBS 0.007228f
C706 B.n582 VSUBS 0.007228f
C707 B.n583 VSUBS 0.007228f
C708 B.n584 VSUBS 0.007228f
C709 B.n585 VSUBS 0.007228f
C710 B.n586 VSUBS 0.007228f
C711 B.n587 VSUBS 0.007228f
C712 B.n588 VSUBS 0.007228f
C713 B.n589 VSUBS 0.007228f
C714 B.n590 VSUBS 0.007228f
C715 B.n591 VSUBS 0.007228f
C716 B.n592 VSUBS 0.007228f
C717 B.n593 VSUBS 0.007228f
C718 B.n594 VSUBS 0.007228f
C719 B.n595 VSUBS 0.007228f
C720 B.n596 VSUBS 0.007228f
C721 B.n597 VSUBS 0.007228f
C722 B.n598 VSUBS 0.007228f
C723 B.n599 VSUBS 0.007228f
C724 B.n600 VSUBS 0.007228f
C725 B.n601 VSUBS 0.007228f
C726 B.n602 VSUBS 0.007228f
C727 B.n603 VSUBS 0.007228f
C728 B.n604 VSUBS 0.007228f
C729 B.n605 VSUBS 0.007228f
C730 B.n606 VSUBS 0.007228f
C731 B.n607 VSUBS 0.007228f
C732 B.n608 VSUBS 0.007228f
C733 B.n609 VSUBS 0.007228f
C734 B.n610 VSUBS 0.007228f
C735 B.n611 VSUBS 0.007228f
C736 B.n612 VSUBS 0.007228f
C737 B.n613 VSUBS 0.007228f
C738 B.n614 VSUBS 0.007228f
C739 B.n615 VSUBS 0.007228f
C740 B.n616 VSUBS 0.007228f
C741 B.n617 VSUBS 0.007228f
C742 B.n618 VSUBS 0.007228f
C743 B.n619 VSUBS 0.007228f
C744 B.n620 VSUBS 0.007228f
C745 B.n621 VSUBS 0.007228f
C746 B.n622 VSUBS 0.017316f
C747 B.n623 VSUBS 0.018188f
C748 B.n624 VSUBS 0.017394f
C749 B.n625 VSUBS 0.007228f
C750 B.n626 VSUBS 0.007228f
C751 B.n627 VSUBS 0.007228f
C752 B.n628 VSUBS 0.007228f
C753 B.n629 VSUBS 0.007228f
C754 B.n630 VSUBS 0.007228f
C755 B.n631 VSUBS 0.007228f
C756 B.n632 VSUBS 0.007228f
C757 B.n633 VSUBS 0.007228f
C758 B.n634 VSUBS 0.007228f
C759 B.n635 VSUBS 0.007228f
C760 B.n636 VSUBS 0.007228f
C761 B.n637 VSUBS 0.007228f
C762 B.n638 VSUBS 0.007228f
C763 B.n639 VSUBS 0.007228f
C764 B.n640 VSUBS 0.007228f
C765 B.n641 VSUBS 0.007228f
C766 B.n642 VSUBS 0.007228f
C767 B.n643 VSUBS 0.007228f
C768 B.n644 VSUBS 0.007228f
C769 B.n645 VSUBS 0.007228f
C770 B.n646 VSUBS 0.007228f
C771 B.n647 VSUBS 0.007228f
C772 B.n648 VSUBS 0.007228f
C773 B.n649 VSUBS 0.007228f
C774 B.n650 VSUBS 0.007228f
C775 B.n651 VSUBS 0.007228f
C776 B.n652 VSUBS 0.007228f
C777 B.n653 VSUBS 0.007228f
C778 B.n654 VSUBS 0.007228f
C779 B.n655 VSUBS 0.007228f
C780 B.n656 VSUBS 0.007228f
C781 B.n657 VSUBS 0.007228f
C782 B.n658 VSUBS 0.007228f
C783 B.n659 VSUBS 0.007228f
C784 B.n660 VSUBS 0.007228f
C785 B.n661 VSUBS 0.007228f
C786 B.n662 VSUBS 0.007228f
C787 B.n663 VSUBS 0.007228f
C788 B.n664 VSUBS 0.007228f
C789 B.n665 VSUBS 0.007228f
C790 B.n666 VSUBS 0.007228f
C791 B.n667 VSUBS 0.007228f
C792 B.n668 VSUBS 0.007228f
C793 B.n669 VSUBS 0.007228f
C794 B.n670 VSUBS 0.007228f
C795 B.n671 VSUBS 0.007228f
C796 B.n672 VSUBS 0.007228f
C797 B.n673 VSUBS 0.007228f
C798 B.n674 VSUBS 0.007228f
C799 B.n675 VSUBS 0.007228f
C800 B.n676 VSUBS 0.007228f
C801 B.n677 VSUBS 0.007228f
C802 B.n678 VSUBS 0.007228f
C803 B.n679 VSUBS 0.007228f
C804 B.n680 VSUBS 0.007228f
C805 B.n681 VSUBS 0.007228f
C806 B.n682 VSUBS 0.007228f
C807 B.n683 VSUBS 0.007228f
C808 B.n684 VSUBS 0.007228f
C809 B.n685 VSUBS 0.007228f
C810 B.n686 VSUBS 0.007228f
C811 B.n687 VSUBS 0.007228f
C812 B.n688 VSUBS 0.007228f
C813 B.n689 VSUBS 0.007228f
C814 B.n690 VSUBS 0.007228f
C815 B.n691 VSUBS 0.004996f
C816 B.n692 VSUBS 0.016747f
C817 B.n693 VSUBS 0.005846f
C818 B.n694 VSUBS 0.007228f
C819 B.n695 VSUBS 0.007228f
C820 B.n696 VSUBS 0.007228f
C821 B.n697 VSUBS 0.007228f
C822 B.n698 VSUBS 0.007228f
C823 B.n699 VSUBS 0.007228f
C824 B.n700 VSUBS 0.007228f
C825 B.n701 VSUBS 0.007228f
C826 B.n702 VSUBS 0.007228f
C827 B.n703 VSUBS 0.007228f
C828 B.n704 VSUBS 0.007228f
C829 B.n705 VSUBS 0.005846f
C830 B.n706 VSUBS 0.007228f
C831 B.n707 VSUBS 0.007228f
C832 B.n708 VSUBS 0.007228f
C833 B.n709 VSUBS 0.007228f
C834 B.n710 VSUBS 0.007228f
C835 B.n711 VSUBS 0.007228f
C836 B.n712 VSUBS 0.007228f
C837 B.n713 VSUBS 0.007228f
C838 B.n714 VSUBS 0.007228f
C839 B.n715 VSUBS 0.007228f
C840 B.n716 VSUBS 0.007228f
C841 B.n717 VSUBS 0.007228f
C842 B.n718 VSUBS 0.007228f
C843 B.n719 VSUBS 0.007228f
C844 B.n720 VSUBS 0.007228f
C845 B.n721 VSUBS 0.007228f
C846 B.n722 VSUBS 0.007228f
C847 B.n723 VSUBS 0.007228f
C848 B.n724 VSUBS 0.007228f
C849 B.n725 VSUBS 0.007228f
C850 B.n726 VSUBS 0.007228f
C851 B.n727 VSUBS 0.007228f
C852 B.n728 VSUBS 0.007228f
C853 B.n729 VSUBS 0.007228f
C854 B.n730 VSUBS 0.007228f
C855 B.n731 VSUBS 0.007228f
C856 B.n732 VSUBS 0.007228f
C857 B.n733 VSUBS 0.007228f
C858 B.n734 VSUBS 0.007228f
C859 B.n735 VSUBS 0.007228f
C860 B.n736 VSUBS 0.007228f
C861 B.n737 VSUBS 0.007228f
C862 B.n738 VSUBS 0.007228f
C863 B.n739 VSUBS 0.007228f
C864 B.n740 VSUBS 0.007228f
C865 B.n741 VSUBS 0.007228f
C866 B.n742 VSUBS 0.007228f
C867 B.n743 VSUBS 0.007228f
C868 B.n744 VSUBS 0.007228f
C869 B.n745 VSUBS 0.007228f
C870 B.n746 VSUBS 0.007228f
C871 B.n747 VSUBS 0.007228f
C872 B.n748 VSUBS 0.007228f
C873 B.n749 VSUBS 0.007228f
C874 B.n750 VSUBS 0.007228f
C875 B.n751 VSUBS 0.007228f
C876 B.n752 VSUBS 0.007228f
C877 B.n753 VSUBS 0.007228f
C878 B.n754 VSUBS 0.007228f
C879 B.n755 VSUBS 0.007228f
C880 B.n756 VSUBS 0.007228f
C881 B.n757 VSUBS 0.007228f
C882 B.n758 VSUBS 0.007228f
C883 B.n759 VSUBS 0.007228f
C884 B.n760 VSUBS 0.007228f
C885 B.n761 VSUBS 0.007228f
C886 B.n762 VSUBS 0.007228f
C887 B.n763 VSUBS 0.007228f
C888 B.n764 VSUBS 0.007228f
C889 B.n765 VSUBS 0.007228f
C890 B.n766 VSUBS 0.007228f
C891 B.n767 VSUBS 0.007228f
C892 B.n768 VSUBS 0.007228f
C893 B.n769 VSUBS 0.007228f
C894 B.n770 VSUBS 0.007228f
C895 B.n771 VSUBS 0.007228f
C896 B.n772 VSUBS 0.007228f
C897 B.n773 VSUBS 0.007228f
C898 B.n774 VSUBS 0.018188f
C899 B.n775 VSUBS 0.018188f
C900 B.n776 VSUBS 0.017316f
C901 B.n777 VSUBS 0.007228f
C902 B.n778 VSUBS 0.007228f
C903 B.n779 VSUBS 0.007228f
C904 B.n780 VSUBS 0.007228f
C905 B.n781 VSUBS 0.007228f
C906 B.n782 VSUBS 0.007228f
C907 B.n783 VSUBS 0.007228f
C908 B.n784 VSUBS 0.007228f
C909 B.n785 VSUBS 0.007228f
C910 B.n786 VSUBS 0.007228f
C911 B.n787 VSUBS 0.007228f
C912 B.n788 VSUBS 0.007228f
C913 B.n789 VSUBS 0.007228f
C914 B.n790 VSUBS 0.007228f
C915 B.n791 VSUBS 0.007228f
C916 B.n792 VSUBS 0.007228f
C917 B.n793 VSUBS 0.007228f
C918 B.n794 VSUBS 0.007228f
C919 B.n795 VSUBS 0.007228f
C920 B.n796 VSUBS 0.007228f
C921 B.n797 VSUBS 0.007228f
C922 B.n798 VSUBS 0.007228f
C923 B.n799 VSUBS 0.007228f
C924 B.n800 VSUBS 0.007228f
C925 B.n801 VSUBS 0.007228f
C926 B.n802 VSUBS 0.007228f
C927 B.n803 VSUBS 0.007228f
C928 B.n804 VSUBS 0.007228f
C929 B.n805 VSUBS 0.007228f
C930 B.n806 VSUBS 0.007228f
C931 B.n807 VSUBS 0.007228f
C932 B.n808 VSUBS 0.007228f
C933 B.n809 VSUBS 0.007228f
C934 B.n810 VSUBS 0.007228f
C935 B.n811 VSUBS 0.007228f
C936 B.n812 VSUBS 0.007228f
C937 B.n813 VSUBS 0.007228f
C938 B.n814 VSUBS 0.007228f
C939 B.n815 VSUBS 0.007228f
C940 B.n816 VSUBS 0.007228f
C941 B.n817 VSUBS 0.007228f
C942 B.n818 VSUBS 0.007228f
C943 B.n819 VSUBS 0.007228f
C944 B.n820 VSUBS 0.007228f
C945 B.n821 VSUBS 0.007228f
C946 B.n822 VSUBS 0.007228f
C947 B.n823 VSUBS 0.007228f
C948 B.n824 VSUBS 0.007228f
C949 B.n825 VSUBS 0.007228f
C950 B.n826 VSUBS 0.007228f
C951 B.n827 VSUBS 0.007228f
C952 B.n828 VSUBS 0.007228f
C953 B.n829 VSUBS 0.007228f
C954 B.n830 VSUBS 0.007228f
C955 B.n831 VSUBS 0.007228f
C956 B.n832 VSUBS 0.007228f
C957 B.n833 VSUBS 0.007228f
C958 B.n834 VSUBS 0.007228f
C959 B.n835 VSUBS 0.007228f
C960 B.n836 VSUBS 0.007228f
C961 B.n837 VSUBS 0.007228f
C962 B.n838 VSUBS 0.007228f
C963 B.n839 VSUBS 0.007228f
C964 B.n840 VSUBS 0.007228f
C965 B.n841 VSUBS 0.007228f
C966 B.n842 VSUBS 0.007228f
C967 B.n843 VSUBS 0.007228f
C968 B.n844 VSUBS 0.007228f
C969 B.n845 VSUBS 0.007228f
C970 B.n846 VSUBS 0.007228f
C971 B.n847 VSUBS 0.007228f
C972 B.n848 VSUBS 0.007228f
C973 B.n849 VSUBS 0.007228f
C974 B.n850 VSUBS 0.007228f
C975 B.n851 VSUBS 0.007228f
C976 B.n852 VSUBS 0.007228f
C977 B.n853 VSUBS 0.007228f
C978 B.n854 VSUBS 0.007228f
C979 B.n855 VSUBS 0.007228f
C980 B.n856 VSUBS 0.007228f
C981 B.n857 VSUBS 0.007228f
C982 B.n858 VSUBS 0.007228f
C983 B.n859 VSUBS 0.016368f
C984 VTAIL.t1 VSUBS 0.264489f
C985 VTAIL.t7 VSUBS 0.264489f
C986 VTAIL.n0 VSUBS 2.00082f
C987 VTAIL.n1 VSUBS 0.77176f
C988 VTAIL.n2 VSUBS 0.027749f
C989 VTAIL.n3 VSUBS 0.02494f
C990 VTAIL.n4 VSUBS 0.013402f
C991 VTAIL.n5 VSUBS 0.031677f
C992 VTAIL.n6 VSUBS 0.01419f
C993 VTAIL.n7 VSUBS 0.02494f
C994 VTAIL.n8 VSUBS 0.013402f
C995 VTAIL.n9 VSUBS 0.031677f
C996 VTAIL.n10 VSUBS 0.01419f
C997 VTAIL.n11 VSUBS 0.02494f
C998 VTAIL.n12 VSUBS 0.013402f
C999 VTAIL.n13 VSUBS 0.031677f
C1000 VTAIL.n14 VSUBS 0.01419f
C1001 VTAIL.n15 VSUBS 0.02494f
C1002 VTAIL.n16 VSUBS 0.013402f
C1003 VTAIL.n17 VSUBS 0.031677f
C1004 VTAIL.n18 VSUBS 0.01419f
C1005 VTAIL.n19 VSUBS 0.02494f
C1006 VTAIL.n20 VSUBS 0.013402f
C1007 VTAIL.n21 VSUBS 0.031677f
C1008 VTAIL.n22 VSUBS 0.01419f
C1009 VTAIL.n23 VSUBS 1.41359f
C1010 VTAIL.n24 VSUBS 0.013402f
C1011 VTAIL.t5 VSUBS 0.067718f
C1012 VTAIL.n25 VSUBS 0.164186f
C1013 VTAIL.n26 VSUBS 0.020152f
C1014 VTAIL.n27 VSUBS 0.023758f
C1015 VTAIL.n28 VSUBS 0.031677f
C1016 VTAIL.n29 VSUBS 0.01419f
C1017 VTAIL.n30 VSUBS 0.013402f
C1018 VTAIL.n31 VSUBS 0.02494f
C1019 VTAIL.n32 VSUBS 0.02494f
C1020 VTAIL.n33 VSUBS 0.013402f
C1021 VTAIL.n34 VSUBS 0.01419f
C1022 VTAIL.n35 VSUBS 0.031677f
C1023 VTAIL.n36 VSUBS 0.031677f
C1024 VTAIL.n37 VSUBS 0.01419f
C1025 VTAIL.n38 VSUBS 0.013402f
C1026 VTAIL.n39 VSUBS 0.02494f
C1027 VTAIL.n40 VSUBS 0.02494f
C1028 VTAIL.n41 VSUBS 0.013402f
C1029 VTAIL.n42 VSUBS 0.01419f
C1030 VTAIL.n43 VSUBS 0.031677f
C1031 VTAIL.n44 VSUBS 0.031677f
C1032 VTAIL.n45 VSUBS 0.01419f
C1033 VTAIL.n46 VSUBS 0.013402f
C1034 VTAIL.n47 VSUBS 0.02494f
C1035 VTAIL.n48 VSUBS 0.02494f
C1036 VTAIL.n49 VSUBS 0.013402f
C1037 VTAIL.n50 VSUBS 0.01419f
C1038 VTAIL.n51 VSUBS 0.031677f
C1039 VTAIL.n52 VSUBS 0.031677f
C1040 VTAIL.n53 VSUBS 0.01419f
C1041 VTAIL.n54 VSUBS 0.013402f
C1042 VTAIL.n55 VSUBS 0.02494f
C1043 VTAIL.n56 VSUBS 0.02494f
C1044 VTAIL.n57 VSUBS 0.013402f
C1045 VTAIL.n58 VSUBS 0.01419f
C1046 VTAIL.n59 VSUBS 0.031677f
C1047 VTAIL.n60 VSUBS 0.031677f
C1048 VTAIL.n61 VSUBS 0.01419f
C1049 VTAIL.n62 VSUBS 0.013402f
C1050 VTAIL.n63 VSUBS 0.02494f
C1051 VTAIL.n64 VSUBS 0.02494f
C1052 VTAIL.n65 VSUBS 0.013402f
C1053 VTAIL.n66 VSUBS 0.01419f
C1054 VTAIL.n67 VSUBS 0.031677f
C1055 VTAIL.n68 VSUBS 0.080293f
C1056 VTAIL.n69 VSUBS 0.01419f
C1057 VTAIL.n70 VSUBS 0.026318f
C1058 VTAIL.n71 VSUBS 0.065144f
C1059 VTAIL.n72 VSUBS 0.062363f
C1060 VTAIL.n73 VSUBS 0.284992f
C1061 VTAIL.n74 VSUBS 0.027749f
C1062 VTAIL.n75 VSUBS 0.02494f
C1063 VTAIL.n76 VSUBS 0.013402f
C1064 VTAIL.n77 VSUBS 0.031677f
C1065 VTAIL.n78 VSUBS 0.01419f
C1066 VTAIL.n79 VSUBS 0.02494f
C1067 VTAIL.n80 VSUBS 0.013402f
C1068 VTAIL.n81 VSUBS 0.031677f
C1069 VTAIL.n82 VSUBS 0.01419f
C1070 VTAIL.n83 VSUBS 0.02494f
C1071 VTAIL.n84 VSUBS 0.013402f
C1072 VTAIL.n85 VSUBS 0.031677f
C1073 VTAIL.n86 VSUBS 0.01419f
C1074 VTAIL.n87 VSUBS 0.02494f
C1075 VTAIL.n88 VSUBS 0.013402f
C1076 VTAIL.n89 VSUBS 0.031677f
C1077 VTAIL.n90 VSUBS 0.01419f
C1078 VTAIL.n91 VSUBS 0.02494f
C1079 VTAIL.n92 VSUBS 0.013402f
C1080 VTAIL.n93 VSUBS 0.031677f
C1081 VTAIL.n94 VSUBS 0.01419f
C1082 VTAIL.n95 VSUBS 1.41359f
C1083 VTAIL.n96 VSUBS 0.013402f
C1084 VTAIL.t14 VSUBS 0.067718f
C1085 VTAIL.n97 VSUBS 0.164186f
C1086 VTAIL.n98 VSUBS 0.020152f
C1087 VTAIL.n99 VSUBS 0.023758f
C1088 VTAIL.n100 VSUBS 0.031677f
C1089 VTAIL.n101 VSUBS 0.01419f
C1090 VTAIL.n102 VSUBS 0.013402f
C1091 VTAIL.n103 VSUBS 0.02494f
C1092 VTAIL.n104 VSUBS 0.02494f
C1093 VTAIL.n105 VSUBS 0.013402f
C1094 VTAIL.n106 VSUBS 0.01419f
C1095 VTAIL.n107 VSUBS 0.031677f
C1096 VTAIL.n108 VSUBS 0.031677f
C1097 VTAIL.n109 VSUBS 0.01419f
C1098 VTAIL.n110 VSUBS 0.013402f
C1099 VTAIL.n111 VSUBS 0.02494f
C1100 VTAIL.n112 VSUBS 0.02494f
C1101 VTAIL.n113 VSUBS 0.013402f
C1102 VTAIL.n114 VSUBS 0.01419f
C1103 VTAIL.n115 VSUBS 0.031677f
C1104 VTAIL.n116 VSUBS 0.031677f
C1105 VTAIL.n117 VSUBS 0.01419f
C1106 VTAIL.n118 VSUBS 0.013402f
C1107 VTAIL.n119 VSUBS 0.02494f
C1108 VTAIL.n120 VSUBS 0.02494f
C1109 VTAIL.n121 VSUBS 0.013402f
C1110 VTAIL.n122 VSUBS 0.01419f
C1111 VTAIL.n123 VSUBS 0.031677f
C1112 VTAIL.n124 VSUBS 0.031677f
C1113 VTAIL.n125 VSUBS 0.01419f
C1114 VTAIL.n126 VSUBS 0.013402f
C1115 VTAIL.n127 VSUBS 0.02494f
C1116 VTAIL.n128 VSUBS 0.02494f
C1117 VTAIL.n129 VSUBS 0.013402f
C1118 VTAIL.n130 VSUBS 0.01419f
C1119 VTAIL.n131 VSUBS 0.031677f
C1120 VTAIL.n132 VSUBS 0.031677f
C1121 VTAIL.n133 VSUBS 0.01419f
C1122 VTAIL.n134 VSUBS 0.013402f
C1123 VTAIL.n135 VSUBS 0.02494f
C1124 VTAIL.n136 VSUBS 0.02494f
C1125 VTAIL.n137 VSUBS 0.013402f
C1126 VTAIL.n138 VSUBS 0.01419f
C1127 VTAIL.n139 VSUBS 0.031677f
C1128 VTAIL.n140 VSUBS 0.080293f
C1129 VTAIL.n141 VSUBS 0.01419f
C1130 VTAIL.n142 VSUBS 0.026318f
C1131 VTAIL.n143 VSUBS 0.065144f
C1132 VTAIL.n144 VSUBS 0.062363f
C1133 VTAIL.n145 VSUBS 0.284992f
C1134 VTAIL.t12 VSUBS 0.264489f
C1135 VTAIL.t9 VSUBS 0.264489f
C1136 VTAIL.n146 VSUBS 2.00082f
C1137 VTAIL.n147 VSUBS 0.988776f
C1138 VTAIL.n148 VSUBS 0.027749f
C1139 VTAIL.n149 VSUBS 0.02494f
C1140 VTAIL.n150 VSUBS 0.013402f
C1141 VTAIL.n151 VSUBS 0.031677f
C1142 VTAIL.n152 VSUBS 0.01419f
C1143 VTAIL.n153 VSUBS 0.02494f
C1144 VTAIL.n154 VSUBS 0.013402f
C1145 VTAIL.n155 VSUBS 0.031677f
C1146 VTAIL.n156 VSUBS 0.01419f
C1147 VTAIL.n157 VSUBS 0.02494f
C1148 VTAIL.n158 VSUBS 0.013402f
C1149 VTAIL.n159 VSUBS 0.031677f
C1150 VTAIL.n160 VSUBS 0.01419f
C1151 VTAIL.n161 VSUBS 0.02494f
C1152 VTAIL.n162 VSUBS 0.013402f
C1153 VTAIL.n163 VSUBS 0.031677f
C1154 VTAIL.n164 VSUBS 0.01419f
C1155 VTAIL.n165 VSUBS 0.02494f
C1156 VTAIL.n166 VSUBS 0.013402f
C1157 VTAIL.n167 VSUBS 0.031677f
C1158 VTAIL.n168 VSUBS 0.01419f
C1159 VTAIL.n169 VSUBS 1.41359f
C1160 VTAIL.n170 VSUBS 0.013402f
C1161 VTAIL.t8 VSUBS 0.067718f
C1162 VTAIL.n171 VSUBS 0.164186f
C1163 VTAIL.n172 VSUBS 0.020152f
C1164 VTAIL.n173 VSUBS 0.023758f
C1165 VTAIL.n174 VSUBS 0.031677f
C1166 VTAIL.n175 VSUBS 0.01419f
C1167 VTAIL.n176 VSUBS 0.013402f
C1168 VTAIL.n177 VSUBS 0.02494f
C1169 VTAIL.n178 VSUBS 0.02494f
C1170 VTAIL.n179 VSUBS 0.013402f
C1171 VTAIL.n180 VSUBS 0.01419f
C1172 VTAIL.n181 VSUBS 0.031677f
C1173 VTAIL.n182 VSUBS 0.031677f
C1174 VTAIL.n183 VSUBS 0.01419f
C1175 VTAIL.n184 VSUBS 0.013402f
C1176 VTAIL.n185 VSUBS 0.02494f
C1177 VTAIL.n186 VSUBS 0.02494f
C1178 VTAIL.n187 VSUBS 0.013402f
C1179 VTAIL.n188 VSUBS 0.01419f
C1180 VTAIL.n189 VSUBS 0.031677f
C1181 VTAIL.n190 VSUBS 0.031677f
C1182 VTAIL.n191 VSUBS 0.01419f
C1183 VTAIL.n192 VSUBS 0.013402f
C1184 VTAIL.n193 VSUBS 0.02494f
C1185 VTAIL.n194 VSUBS 0.02494f
C1186 VTAIL.n195 VSUBS 0.013402f
C1187 VTAIL.n196 VSUBS 0.01419f
C1188 VTAIL.n197 VSUBS 0.031677f
C1189 VTAIL.n198 VSUBS 0.031677f
C1190 VTAIL.n199 VSUBS 0.01419f
C1191 VTAIL.n200 VSUBS 0.013402f
C1192 VTAIL.n201 VSUBS 0.02494f
C1193 VTAIL.n202 VSUBS 0.02494f
C1194 VTAIL.n203 VSUBS 0.013402f
C1195 VTAIL.n204 VSUBS 0.01419f
C1196 VTAIL.n205 VSUBS 0.031677f
C1197 VTAIL.n206 VSUBS 0.031677f
C1198 VTAIL.n207 VSUBS 0.01419f
C1199 VTAIL.n208 VSUBS 0.013402f
C1200 VTAIL.n209 VSUBS 0.02494f
C1201 VTAIL.n210 VSUBS 0.02494f
C1202 VTAIL.n211 VSUBS 0.013402f
C1203 VTAIL.n212 VSUBS 0.01419f
C1204 VTAIL.n213 VSUBS 0.031677f
C1205 VTAIL.n214 VSUBS 0.080293f
C1206 VTAIL.n215 VSUBS 0.01419f
C1207 VTAIL.n216 VSUBS 0.026318f
C1208 VTAIL.n217 VSUBS 0.065144f
C1209 VTAIL.n218 VSUBS 0.062363f
C1210 VTAIL.n219 VSUBS 1.73743f
C1211 VTAIL.n220 VSUBS 0.027749f
C1212 VTAIL.n221 VSUBS 0.02494f
C1213 VTAIL.n222 VSUBS 0.013402f
C1214 VTAIL.n223 VSUBS 0.031677f
C1215 VTAIL.n224 VSUBS 0.01419f
C1216 VTAIL.n225 VSUBS 0.02494f
C1217 VTAIL.n226 VSUBS 0.013402f
C1218 VTAIL.n227 VSUBS 0.031677f
C1219 VTAIL.n228 VSUBS 0.01419f
C1220 VTAIL.n229 VSUBS 0.02494f
C1221 VTAIL.n230 VSUBS 0.013402f
C1222 VTAIL.n231 VSUBS 0.031677f
C1223 VTAIL.n232 VSUBS 0.01419f
C1224 VTAIL.n233 VSUBS 0.02494f
C1225 VTAIL.n234 VSUBS 0.013402f
C1226 VTAIL.n235 VSUBS 0.031677f
C1227 VTAIL.n236 VSUBS 0.01419f
C1228 VTAIL.n237 VSUBS 0.02494f
C1229 VTAIL.n238 VSUBS 0.013402f
C1230 VTAIL.n239 VSUBS 0.031677f
C1231 VTAIL.n240 VSUBS 0.01419f
C1232 VTAIL.n241 VSUBS 1.41359f
C1233 VTAIL.n242 VSUBS 0.013402f
C1234 VTAIL.t3 VSUBS 0.067718f
C1235 VTAIL.n243 VSUBS 0.164186f
C1236 VTAIL.n244 VSUBS 0.020152f
C1237 VTAIL.n245 VSUBS 0.023758f
C1238 VTAIL.n246 VSUBS 0.031677f
C1239 VTAIL.n247 VSUBS 0.01419f
C1240 VTAIL.n248 VSUBS 0.013402f
C1241 VTAIL.n249 VSUBS 0.02494f
C1242 VTAIL.n250 VSUBS 0.02494f
C1243 VTAIL.n251 VSUBS 0.013402f
C1244 VTAIL.n252 VSUBS 0.01419f
C1245 VTAIL.n253 VSUBS 0.031677f
C1246 VTAIL.n254 VSUBS 0.031677f
C1247 VTAIL.n255 VSUBS 0.01419f
C1248 VTAIL.n256 VSUBS 0.013402f
C1249 VTAIL.n257 VSUBS 0.02494f
C1250 VTAIL.n258 VSUBS 0.02494f
C1251 VTAIL.n259 VSUBS 0.013402f
C1252 VTAIL.n260 VSUBS 0.01419f
C1253 VTAIL.n261 VSUBS 0.031677f
C1254 VTAIL.n262 VSUBS 0.031677f
C1255 VTAIL.n263 VSUBS 0.01419f
C1256 VTAIL.n264 VSUBS 0.013402f
C1257 VTAIL.n265 VSUBS 0.02494f
C1258 VTAIL.n266 VSUBS 0.02494f
C1259 VTAIL.n267 VSUBS 0.013402f
C1260 VTAIL.n268 VSUBS 0.01419f
C1261 VTAIL.n269 VSUBS 0.031677f
C1262 VTAIL.n270 VSUBS 0.031677f
C1263 VTAIL.n271 VSUBS 0.01419f
C1264 VTAIL.n272 VSUBS 0.013402f
C1265 VTAIL.n273 VSUBS 0.02494f
C1266 VTAIL.n274 VSUBS 0.02494f
C1267 VTAIL.n275 VSUBS 0.013402f
C1268 VTAIL.n276 VSUBS 0.01419f
C1269 VTAIL.n277 VSUBS 0.031677f
C1270 VTAIL.n278 VSUBS 0.031677f
C1271 VTAIL.n279 VSUBS 0.01419f
C1272 VTAIL.n280 VSUBS 0.013402f
C1273 VTAIL.n281 VSUBS 0.02494f
C1274 VTAIL.n282 VSUBS 0.02494f
C1275 VTAIL.n283 VSUBS 0.013402f
C1276 VTAIL.n284 VSUBS 0.01419f
C1277 VTAIL.n285 VSUBS 0.031677f
C1278 VTAIL.n286 VSUBS 0.080293f
C1279 VTAIL.n287 VSUBS 0.01419f
C1280 VTAIL.n288 VSUBS 0.026318f
C1281 VTAIL.n289 VSUBS 0.065144f
C1282 VTAIL.n290 VSUBS 0.062363f
C1283 VTAIL.n291 VSUBS 1.73743f
C1284 VTAIL.t6 VSUBS 0.264489f
C1285 VTAIL.t4 VSUBS 0.264489f
C1286 VTAIL.n292 VSUBS 2.00084f
C1287 VTAIL.n293 VSUBS 0.988762f
C1288 VTAIL.n294 VSUBS 0.027749f
C1289 VTAIL.n295 VSUBS 0.02494f
C1290 VTAIL.n296 VSUBS 0.013402f
C1291 VTAIL.n297 VSUBS 0.031677f
C1292 VTAIL.n298 VSUBS 0.01419f
C1293 VTAIL.n299 VSUBS 0.02494f
C1294 VTAIL.n300 VSUBS 0.013402f
C1295 VTAIL.n301 VSUBS 0.031677f
C1296 VTAIL.n302 VSUBS 0.01419f
C1297 VTAIL.n303 VSUBS 0.02494f
C1298 VTAIL.n304 VSUBS 0.013402f
C1299 VTAIL.n305 VSUBS 0.031677f
C1300 VTAIL.n306 VSUBS 0.01419f
C1301 VTAIL.n307 VSUBS 0.02494f
C1302 VTAIL.n308 VSUBS 0.013402f
C1303 VTAIL.n309 VSUBS 0.031677f
C1304 VTAIL.n310 VSUBS 0.01419f
C1305 VTAIL.n311 VSUBS 0.02494f
C1306 VTAIL.n312 VSUBS 0.013402f
C1307 VTAIL.n313 VSUBS 0.031677f
C1308 VTAIL.n314 VSUBS 0.01419f
C1309 VTAIL.n315 VSUBS 1.41359f
C1310 VTAIL.n316 VSUBS 0.013402f
C1311 VTAIL.t2 VSUBS 0.067718f
C1312 VTAIL.n317 VSUBS 0.164186f
C1313 VTAIL.n318 VSUBS 0.020152f
C1314 VTAIL.n319 VSUBS 0.023758f
C1315 VTAIL.n320 VSUBS 0.031677f
C1316 VTAIL.n321 VSUBS 0.01419f
C1317 VTAIL.n322 VSUBS 0.013402f
C1318 VTAIL.n323 VSUBS 0.02494f
C1319 VTAIL.n324 VSUBS 0.02494f
C1320 VTAIL.n325 VSUBS 0.013402f
C1321 VTAIL.n326 VSUBS 0.01419f
C1322 VTAIL.n327 VSUBS 0.031677f
C1323 VTAIL.n328 VSUBS 0.031677f
C1324 VTAIL.n329 VSUBS 0.01419f
C1325 VTAIL.n330 VSUBS 0.013402f
C1326 VTAIL.n331 VSUBS 0.02494f
C1327 VTAIL.n332 VSUBS 0.02494f
C1328 VTAIL.n333 VSUBS 0.013402f
C1329 VTAIL.n334 VSUBS 0.01419f
C1330 VTAIL.n335 VSUBS 0.031677f
C1331 VTAIL.n336 VSUBS 0.031677f
C1332 VTAIL.n337 VSUBS 0.01419f
C1333 VTAIL.n338 VSUBS 0.013402f
C1334 VTAIL.n339 VSUBS 0.02494f
C1335 VTAIL.n340 VSUBS 0.02494f
C1336 VTAIL.n341 VSUBS 0.013402f
C1337 VTAIL.n342 VSUBS 0.01419f
C1338 VTAIL.n343 VSUBS 0.031677f
C1339 VTAIL.n344 VSUBS 0.031677f
C1340 VTAIL.n345 VSUBS 0.01419f
C1341 VTAIL.n346 VSUBS 0.013402f
C1342 VTAIL.n347 VSUBS 0.02494f
C1343 VTAIL.n348 VSUBS 0.02494f
C1344 VTAIL.n349 VSUBS 0.013402f
C1345 VTAIL.n350 VSUBS 0.01419f
C1346 VTAIL.n351 VSUBS 0.031677f
C1347 VTAIL.n352 VSUBS 0.031677f
C1348 VTAIL.n353 VSUBS 0.01419f
C1349 VTAIL.n354 VSUBS 0.013402f
C1350 VTAIL.n355 VSUBS 0.02494f
C1351 VTAIL.n356 VSUBS 0.02494f
C1352 VTAIL.n357 VSUBS 0.013402f
C1353 VTAIL.n358 VSUBS 0.01419f
C1354 VTAIL.n359 VSUBS 0.031677f
C1355 VTAIL.n360 VSUBS 0.080293f
C1356 VTAIL.n361 VSUBS 0.01419f
C1357 VTAIL.n362 VSUBS 0.026318f
C1358 VTAIL.n363 VSUBS 0.065144f
C1359 VTAIL.n364 VSUBS 0.062363f
C1360 VTAIL.n365 VSUBS 0.284992f
C1361 VTAIL.n366 VSUBS 0.027749f
C1362 VTAIL.n367 VSUBS 0.02494f
C1363 VTAIL.n368 VSUBS 0.013402f
C1364 VTAIL.n369 VSUBS 0.031677f
C1365 VTAIL.n370 VSUBS 0.01419f
C1366 VTAIL.n371 VSUBS 0.02494f
C1367 VTAIL.n372 VSUBS 0.013402f
C1368 VTAIL.n373 VSUBS 0.031677f
C1369 VTAIL.n374 VSUBS 0.01419f
C1370 VTAIL.n375 VSUBS 0.02494f
C1371 VTAIL.n376 VSUBS 0.013402f
C1372 VTAIL.n377 VSUBS 0.031677f
C1373 VTAIL.n378 VSUBS 0.01419f
C1374 VTAIL.n379 VSUBS 0.02494f
C1375 VTAIL.n380 VSUBS 0.013402f
C1376 VTAIL.n381 VSUBS 0.031677f
C1377 VTAIL.n382 VSUBS 0.01419f
C1378 VTAIL.n383 VSUBS 0.02494f
C1379 VTAIL.n384 VSUBS 0.013402f
C1380 VTAIL.n385 VSUBS 0.031677f
C1381 VTAIL.n386 VSUBS 0.01419f
C1382 VTAIL.n387 VSUBS 1.41359f
C1383 VTAIL.n388 VSUBS 0.013402f
C1384 VTAIL.t15 VSUBS 0.067718f
C1385 VTAIL.n389 VSUBS 0.164186f
C1386 VTAIL.n390 VSUBS 0.020152f
C1387 VTAIL.n391 VSUBS 0.023758f
C1388 VTAIL.n392 VSUBS 0.031677f
C1389 VTAIL.n393 VSUBS 0.01419f
C1390 VTAIL.n394 VSUBS 0.013402f
C1391 VTAIL.n395 VSUBS 0.02494f
C1392 VTAIL.n396 VSUBS 0.02494f
C1393 VTAIL.n397 VSUBS 0.013402f
C1394 VTAIL.n398 VSUBS 0.01419f
C1395 VTAIL.n399 VSUBS 0.031677f
C1396 VTAIL.n400 VSUBS 0.031677f
C1397 VTAIL.n401 VSUBS 0.01419f
C1398 VTAIL.n402 VSUBS 0.013402f
C1399 VTAIL.n403 VSUBS 0.02494f
C1400 VTAIL.n404 VSUBS 0.02494f
C1401 VTAIL.n405 VSUBS 0.013402f
C1402 VTAIL.n406 VSUBS 0.01419f
C1403 VTAIL.n407 VSUBS 0.031677f
C1404 VTAIL.n408 VSUBS 0.031677f
C1405 VTAIL.n409 VSUBS 0.01419f
C1406 VTAIL.n410 VSUBS 0.013402f
C1407 VTAIL.n411 VSUBS 0.02494f
C1408 VTAIL.n412 VSUBS 0.02494f
C1409 VTAIL.n413 VSUBS 0.013402f
C1410 VTAIL.n414 VSUBS 0.01419f
C1411 VTAIL.n415 VSUBS 0.031677f
C1412 VTAIL.n416 VSUBS 0.031677f
C1413 VTAIL.n417 VSUBS 0.01419f
C1414 VTAIL.n418 VSUBS 0.013402f
C1415 VTAIL.n419 VSUBS 0.02494f
C1416 VTAIL.n420 VSUBS 0.02494f
C1417 VTAIL.n421 VSUBS 0.013402f
C1418 VTAIL.n422 VSUBS 0.01419f
C1419 VTAIL.n423 VSUBS 0.031677f
C1420 VTAIL.n424 VSUBS 0.031677f
C1421 VTAIL.n425 VSUBS 0.01419f
C1422 VTAIL.n426 VSUBS 0.013402f
C1423 VTAIL.n427 VSUBS 0.02494f
C1424 VTAIL.n428 VSUBS 0.02494f
C1425 VTAIL.n429 VSUBS 0.013402f
C1426 VTAIL.n430 VSUBS 0.01419f
C1427 VTAIL.n431 VSUBS 0.031677f
C1428 VTAIL.n432 VSUBS 0.080293f
C1429 VTAIL.n433 VSUBS 0.01419f
C1430 VTAIL.n434 VSUBS 0.026318f
C1431 VTAIL.n435 VSUBS 0.065144f
C1432 VTAIL.n436 VSUBS 0.062363f
C1433 VTAIL.n437 VSUBS 0.284992f
C1434 VTAIL.t13 VSUBS 0.264489f
C1435 VTAIL.t11 VSUBS 0.264489f
C1436 VTAIL.n438 VSUBS 2.00084f
C1437 VTAIL.n439 VSUBS 0.988762f
C1438 VTAIL.n440 VSUBS 0.027749f
C1439 VTAIL.n441 VSUBS 0.02494f
C1440 VTAIL.n442 VSUBS 0.013402f
C1441 VTAIL.n443 VSUBS 0.031677f
C1442 VTAIL.n444 VSUBS 0.01419f
C1443 VTAIL.n445 VSUBS 0.02494f
C1444 VTAIL.n446 VSUBS 0.013402f
C1445 VTAIL.n447 VSUBS 0.031677f
C1446 VTAIL.n448 VSUBS 0.01419f
C1447 VTAIL.n449 VSUBS 0.02494f
C1448 VTAIL.n450 VSUBS 0.013402f
C1449 VTAIL.n451 VSUBS 0.031677f
C1450 VTAIL.n452 VSUBS 0.01419f
C1451 VTAIL.n453 VSUBS 0.02494f
C1452 VTAIL.n454 VSUBS 0.013402f
C1453 VTAIL.n455 VSUBS 0.031677f
C1454 VTAIL.n456 VSUBS 0.01419f
C1455 VTAIL.n457 VSUBS 0.02494f
C1456 VTAIL.n458 VSUBS 0.013402f
C1457 VTAIL.n459 VSUBS 0.031677f
C1458 VTAIL.n460 VSUBS 0.01419f
C1459 VTAIL.n461 VSUBS 1.41359f
C1460 VTAIL.n462 VSUBS 0.013402f
C1461 VTAIL.t10 VSUBS 0.067718f
C1462 VTAIL.n463 VSUBS 0.164186f
C1463 VTAIL.n464 VSUBS 0.020152f
C1464 VTAIL.n465 VSUBS 0.023758f
C1465 VTAIL.n466 VSUBS 0.031677f
C1466 VTAIL.n467 VSUBS 0.01419f
C1467 VTAIL.n468 VSUBS 0.013402f
C1468 VTAIL.n469 VSUBS 0.02494f
C1469 VTAIL.n470 VSUBS 0.02494f
C1470 VTAIL.n471 VSUBS 0.013402f
C1471 VTAIL.n472 VSUBS 0.01419f
C1472 VTAIL.n473 VSUBS 0.031677f
C1473 VTAIL.n474 VSUBS 0.031677f
C1474 VTAIL.n475 VSUBS 0.01419f
C1475 VTAIL.n476 VSUBS 0.013402f
C1476 VTAIL.n477 VSUBS 0.02494f
C1477 VTAIL.n478 VSUBS 0.02494f
C1478 VTAIL.n479 VSUBS 0.013402f
C1479 VTAIL.n480 VSUBS 0.01419f
C1480 VTAIL.n481 VSUBS 0.031677f
C1481 VTAIL.n482 VSUBS 0.031677f
C1482 VTAIL.n483 VSUBS 0.01419f
C1483 VTAIL.n484 VSUBS 0.013402f
C1484 VTAIL.n485 VSUBS 0.02494f
C1485 VTAIL.n486 VSUBS 0.02494f
C1486 VTAIL.n487 VSUBS 0.013402f
C1487 VTAIL.n488 VSUBS 0.01419f
C1488 VTAIL.n489 VSUBS 0.031677f
C1489 VTAIL.n490 VSUBS 0.031677f
C1490 VTAIL.n491 VSUBS 0.01419f
C1491 VTAIL.n492 VSUBS 0.013402f
C1492 VTAIL.n493 VSUBS 0.02494f
C1493 VTAIL.n494 VSUBS 0.02494f
C1494 VTAIL.n495 VSUBS 0.013402f
C1495 VTAIL.n496 VSUBS 0.01419f
C1496 VTAIL.n497 VSUBS 0.031677f
C1497 VTAIL.n498 VSUBS 0.031677f
C1498 VTAIL.n499 VSUBS 0.01419f
C1499 VTAIL.n500 VSUBS 0.013402f
C1500 VTAIL.n501 VSUBS 0.02494f
C1501 VTAIL.n502 VSUBS 0.02494f
C1502 VTAIL.n503 VSUBS 0.013402f
C1503 VTAIL.n504 VSUBS 0.01419f
C1504 VTAIL.n505 VSUBS 0.031677f
C1505 VTAIL.n506 VSUBS 0.080293f
C1506 VTAIL.n507 VSUBS 0.01419f
C1507 VTAIL.n508 VSUBS 0.026318f
C1508 VTAIL.n509 VSUBS 0.065144f
C1509 VTAIL.n510 VSUBS 0.062363f
C1510 VTAIL.n511 VSUBS 1.73743f
C1511 VTAIL.n512 VSUBS 0.027749f
C1512 VTAIL.n513 VSUBS 0.02494f
C1513 VTAIL.n514 VSUBS 0.013402f
C1514 VTAIL.n515 VSUBS 0.031677f
C1515 VTAIL.n516 VSUBS 0.01419f
C1516 VTAIL.n517 VSUBS 0.02494f
C1517 VTAIL.n518 VSUBS 0.013402f
C1518 VTAIL.n519 VSUBS 0.031677f
C1519 VTAIL.n520 VSUBS 0.01419f
C1520 VTAIL.n521 VSUBS 0.02494f
C1521 VTAIL.n522 VSUBS 0.013402f
C1522 VTAIL.n523 VSUBS 0.031677f
C1523 VTAIL.n524 VSUBS 0.01419f
C1524 VTAIL.n525 VSUBS 0.02494f
C1525 VTAIL.n526 VSUBS 0.013402f
C1526 VTAIL.n527 VSUBS 0.031677f
C1527 VTAIL.n528 VSUBS 0.01419f
C1528 VTAIL.n529 VSUBS 0.02494f
C1529 VTAIL.n530 VSUBS 0.013402f
C1530 VTAIL.n531 VSUBS 0.031677f
C1531 VTAIL.n532 VSUBS 0.01419f
C1532 VTAIL.n533 VSUBS 1.41359f
C1533 VTAIL.n534 VSUBS 0.013402f
C1534 VTAIL.t0 VSUBS 0.067718f
C1535 VTAIL.n535 VSUBS 0.164186f
C1536 VTAIL.n536 VSUBS 0.020152f
C1537 VTAIL.n537 VSUBS 0.023758f
C1538 VTAIL.n538 VSUBS 0.031677f
C1539 VTAIL.n539 VSUBS 0.01419f
C1540 VTAIL.n540 VSUBS 0.013402f
C1541 VTAIL.n541 VSUBS 0.02494f
C1542 VTAIL.n542 VSUBS 0.02494f
C1543 VTAIL.n543 VSUBS 0.013402f
C1544 VTAIL.n544 VSUBS 0.01419f
C1545 VTAIL.n545 VSUBS 0.031677f
C1546 VTAIL.n546 VSUBS 0.031677f
C1547 VTAIL.n547 VSUBS 0.01419f
C1548 VTAIL.n548 VSUBS 0.013402f
C1549 VTAIL.n549 VSUBS 0.02494f
C1550 VTAIL.n550 VSUBS 0.02494f
C1551 VTAIL.n551 VSUBS 0.013402f
C1552 VTAIL.n552 VSUBS 0.01419f
C1553 VTAIL.n553 VSUBS 0.031677f
C1554 VTAIL.n554 VSUBS 0.031677f
C1555 VTAIL.n555 VSUBS 0.01419f
C1556 VTAIL.n556 VSUBS 0.013402f
C1557 VTAIL.n557 VSUBS 0.02494f
C1558 VTAIL.n558 VSUBS 0.02494f
C1559 VTAIL.n559 VSUBS 0.013402f
C1560 VTAIL.n560 VSUBS 0.01419f
C1561 VTAIL.n561 VSUBS 0.031677f
C1562 VTAIL.n562 VSUBS 0.031677f
C1563 VTAIL.n563 VSUBS 0.01419f
C1564 VTAIL.n564 VSUBS 0.013402f
C1565 VTAIL.n565 VSUBS 0.02494f
C1566 VTAIL.n566 VSUBS 0.02494f
C1567 VTAIL.n567 VSUBS 0.013402f
C1568 VTAIL.n568 VSUBS 0.01419f
C1569 VTAIL.n569 VSUBS 0.031677f
C1570 VTAIL.n570 VSUBS 0.031677f
C1571 VTAIL.n571 VSUBS 0.01419f
C1572 VTAIL.n572 VSUBS 0.013402f
C1573 VTAIL.n573 VSUBS 0.02494f
C1574 VTAIL.n574 VSUBS 0.02494f
C1575 VTAIL.n575 VSUBS 0.013402f
C1576 VTAIL.n576 VSUBS 0.01419f
C1577 VTAIL.n577 VSUBS 0.031677f
C1578 VTAIL.n578 VSUBS 0.080293f
C1579 VTAIL.n579 VSUBS 0.01419f
C1580 VTAIL.n580 VSUBS 0.026318f
C1581 VTAIL.n581 VSUBS 0.065144f
C1582 VTAIL.n582 VSUBS 0.062363f
C1583 VTAIL.n583 VSUBS 1.73275f
C1584 VDD1.t3 VSUBS 0.289979f
C1585 VDD1.t6 VSUBS 0.289979f
C1586 VDD1.n0 VSUBS 2.34773f
C1587 VDD1.t7 VSUBS 0.289979f
C1588 VDD1.t0 VSUBS 0.289979f
C1589 VDD1.n1 VSUBS 2.34629f
C1590 VDD1.t4 VSUBS 0.289979f
C1591 VDD1.t5 VSUBS 0.289979f
C1592 VDD1.n2 VSUBS 2.34629f
C1593 VDD1.n3 VSUBS 4.45008f
C1594 VDD1.t1 VSUBS 0.289979f
C1595 VDD1.t2 VSUBS 0.289979f
C1596 VDD1.n4 VSUBS 2.33147f
C1597 VDD1.n5 VSUBS 3.75349f
C1598 VP.n0 VSUBS 0.038215f
C1599 VP.t1 VSUBS 3.05118f
C1600 VP.n1 VSUBS 0.058223f
C1601 VP.n2 VSUBS 0.028988f
C1602 VP.n3 VSUBS 0.035179f
C1603 VP.n4 VSUBS 0.028988f
C1604 VP.n5 VSUBS 0.042138f
C1605 VP.n6 VSUBS 0.028988f
C1606 VP.t3 VSUBS 3.05118f
C1607 VP.n7 VSUBS 0.053755f
C1608 VP.n8 VSUBS 0.028988f
C1609 VP.n9 VSUBS 0.053755f
C1610 VP.n10 VSUBS 0.038215f
C1611 VP.t5 VSUBS 3.05118f
C1612 VP.n11 VSUBS 0.058223f
C1613 VP.n12 VSUBS 0.028988f
C1614 VP.n13 VSUBS 0.035179f
C1615 VP.n14 VSUBS 0.028988f
C1616 VP.n15 VSUBS 0.042138f
C1617 VP.n16 VSUBS 0.306438f
C1618 VP.t2 VSUBS 3.05118f
C1619 VP.t0 VSUBS 3.33787f
C1620 VP.n17 VSUBS 1.12019f
C1621 VP.n18 VSUBS 1.16436f
C1622 VP.n19 VSUBS 0.045794f
C1623 VP.n20 VSUBS 0.053755f
C1624 VP.n21 VSUBS 0.028988f
C1625 VP.n22 VSUBS 0.028988f
C1626 VP.n23 VSUBS 0.028988f
C1627 VP.n24 VSUBS 0.042138f
C1628 VP.n25 VSUBS 0.053755f
C1629 VP.t4 VSUBS 3.05118f
C1630 VP.n26 VSUBS 1.0695f
C1631 VP.n27 VSUBS 0.045794f
C1632 VP.n28 VSUBS 0.028988f
C1633 VP.n29 VSUBS 0.028988f
C1634 VP.n30 VSUBS 0.028988f
C1635 VP.n31 VSUBS 0.053755f
C1636 VP.n32 VSUBS 0.055459f
C1637 VP.n33 VSUBS 0.02435f
C1638 VP.n34 VSUBS 0.028988f
C1639 VP.n35 VSUBS 0.028988f
C1640 VP.n36 VSUBS 0.028988f
C1641 VP.n37 VSUBS 0.053755f
C1642 VP.n38 VSUBS 0.029872f
C1643 VP.n39 VSUBS 1.16453f
C1644 VP.n40 VSUBS 1.77269f
C1645 VP.n41 VSUBS 1.79233f
C1646 VP.t7 VSUBS 3.05118f
C1647 VP.n42 VSUBS 1.16453f
C1648 VP.n43 VSUBS 0.029872f
C1649 VP.n44 VSUBS 0.038215f
C1650 VP.n45 VSUBS 0.028988f
C1651 VP.n46 VSUBS 0.028988f
C1652 VP.n47 VSUBS 0.058223f
C1653 VP.n48 VSUBS 0.02435f
C1654 VP.n49 VSUBS 0.055459f
C1655 VP.n50 VSUBS 0.028988f
C1656 VP.n51 VSUBS 0.028988f
C1657 VP.n52 VSUBS 0.028988f
C1658 VP.n53 VSUBS 0.035179f
C1659 VP.n54 VSUBS 1.0695f
C1660 VP.n55 VSUBS 0.045794f
C1661 VP.n56 VSUBS 0.053755f
C1662 VP.n57 VSUBS 0.028988f
C1663 VP.n58 VSUBS 0.028988f
C1664 VP.n59 VSUBS 0.028988f
C1665 VP.n60 VSUBS 0.042138f
C1666 VP.n61 VSUBS 0.053755f
C1667 VP.t6 VSUBS 3.05118f
C1668 VP.n62 VSUBS 1.0695f
C1669 VP.n63 VSUBS 0.045794f
C1670 VP.n64 VSUBS 0.028988f
C1671 VP.n65 VSUBS 0.028988f
C1672 VP.n66 VSUBS 0.028988f
C1673 VP.n67 VSUBS 0.053755f
C1674 VP.n68 VSUBS 0.055459f
C1675 VP.n69 VSUBS 0.02435f
C1676 VP.n70 VSUBS 0.028988f
C1677 VP.n71 VSUBS 0.028988f
C1678 VP.n72 VSUBS 0.028988f
C1679 VP.n73 VSUBS 0.053755f
C1680 VP.n74 VSUBS 0.029872f
C1681 VP.n75 VSUBS 1.16453f
C1682 VP.n76 VSUBS 0.055115f
.ends

