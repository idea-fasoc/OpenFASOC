* NGSPICE file created from diff_pair_sample_0285.ext - technology: sky130A

.subckt diff_pair_sample_0285 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n2662_n3362# sky130_fd_pr__pfet_01v8 ad=4.6683 pd=24.72 as=0 ps=0 w=11.97 l=2.49
X1 VDD2.t3 VN.t0 VTAIL.t5 w_n2662_n3362# sky130_fd_pr__pfet_01v8 ad=1.97505 pd=12.3 as=4.6683 ps=24.72 w=11.97 l=2.49
X2 VDD1.t3 VP.t0 VTAIL.t3 w_n2662_n3362# sky130_fd_pr__pfet_01v8 ad=1.97505 pd=12.3 as=4.6683 ps=24.72 w=11.97 l=2.49
X3 VTAIL.t7 VN.t1 VDD2.t2 w_n2662_n3362# sky130_fd_pr__pfet_01v8 ad=4.6683 pd=24.72 as=1.97505 ps=12.3 w=11.97 l=2.49
X4 VTAIL.t4 VN.t2 VDD2.t1 w_n2662_n3362# sky130_fd_pr__pfet_01v8 ad=4.6683 pd=24.72 as=1.97505 ps=12.3 w=11.97 l=2.49
X5 VDD2.t0 VN.t3 VTAIL.t6 w_n2662_n3362# sky130_fd_pr__pfet_01v8 ad=1.97505 pd=12.3 as=4.6683 ps=24.72 w=11.97 l=2.49
X6 B.t8 B.t6 B.t7 w_n2662_n3362# sky130_fd_pr__pfet_01v8 ad=4.6683 pd=24.72 as=0 ps=0 w=11.97 l=2.49
X7 VTAIL.t1 VP.t1 VDD1.t2 w_n2662_n3362# sky130_fd_pr__pfet_01v8 ad=4.6683 pd=24.72 as=1.97505 ps=12.3 w=11.97 l=2.49
X8 B.t5 B.t3 B.t4 w_n2662_n3362# sky130_fd_pr__pfet_01v8 ad=4.6683 pd=24.72 as=0 ps=0 w=11.97 l=2.49
X9 VDD1.t1 VP.t2 VTAIL.t0 w_n2662_n3362# sky130_fd_pr__pfet_01v8 ad=1.97505 pd=12.3 as=4.6683 ps=24.72 w=11.97 l=2.49
X10 B.t2 B.t0 B.t1 w_n2662_n3362# sky130_fd_pr__pfet_01v8 ad=4.6683 pd=24.72 as=0 ps=0 w=11.97 l=2.49
X11 VTAIL.t2 VP.t3 VDD1.t0 w_n2662_n3362# sky130_fd_pr__pfet_01v8 ad=4.6683 pd=24.72 as=1.97505 ps=12.3 w=11.97 l=2.49
R0 B.n460 B.n69 585
R1 B.n462 B.n461 585
R2 B.n463 B.n68 585
R3 B.n465 B.n464 585
R4 B.n466 B.n67 585
R5 B.n468 B.n467 585
R6 B.n469 B.n66 585
R7 B.n471 B.n470 585
R8 B.n472 B.n65 585
R9 B.n474 B.n473 585
R10 B.n475 B.n64 585
R11 B.n477 B.n476 585
R12 B.n478 B.n63 585
R13 B.n480 B.n479 585
R14 B.n481 B.n62 585
R15 B.n483 B.n482 585
R16 B.n484 B.n61 585
R17 B.n486 B.n485 585
R18 B.n487 B.n60 585
R19 B.n489 B.n488 585
R20 B.n490 B.n59 585
R21 B.n492 B.n491 585
R22 B.n493 B.n58 585
R23 B.n495 B.n494 585
R24 B.n496 B.n57 585
R25 B.n498 B.n497 585
R26 B.n499 B.n56 585
R27 B.n501 B.n500 585
R28 B.n502 B.n55 585
R29 B.n504 B.n503 585
R30 B.n505 B.n54 585
R31 B.n507 B.n506 585
R32 B.n508 B.n53 585
R33 B.n510 B.n509 585
R34 B.n511 B.n52 585
R35 B.n513 B.n512 585
R36 B.n514 B.n51 585
R37 B.n516 B.n515 585
R38 B.n517 B.n50 585
R39 B.n519 B.n518 585
R40 B.n520 B.n49 585
R41 B.n522 B.n521 585
R42 B.n524 B.n523 585
R43 B.n525 B.n45 585
R44 B.n527 B.n526 585
R45 B.n528 B.n44 585
R46 B.n530 B.n529 585
R47 B.n531 B.n43 585
R48 B.n533 B.n532 585
R49 B.n534 B.n42 585
R50 B.n536 B.n535 585
R51 B.n538 B.n39 585
R52 B.n540 B.n539 585
R53 B.n541 B.n38 585
R54 B.n543 B.n542 585
R55 B.n544 B.n37 585
R56 B.n546 B.n545 585
R57 B.n547 B.n36 585
R58 B.n549 B.n548 585
R59 B.n550 B.n35 585
R60 B.n552 B.n551 585
R61 B.n553 B.n34 585
R62 B.n555 B.n554 585
R63 B.n556 B.n33 585
R64 B.n558 B.n557 585
R65 B.n559 B.n32 585
R66 B.n561 B.n560 585
R67 B.n562 B.n31 585
R68 B.n564 B.n563 585
R69 B.n565 B.n30 585
R70 B.n567 B.n566 585
R71 B.n568 B.n29 585
R72 B.n570 B.n569 585
R73 B.n571 B.n28 585
R74 B.n573 B.n572 585
R75 B.n574 B.n27 585
R76 B.n576 B.n575 585
R77 B.n577 B.n26 585
R78 B.n579 B.n578 585
R79 B.n580 B.n25 585
R80 B.n582 B.n581 585
R81 B.n583 B.n24 585
R82 B.n585 B.n584 585
R83 B.n586 B.n23 585
R84 B.n588 B.n587 585
R85 B.n589 B.n22 585
R86 B.n591 B.n590 585
R87 B.n592 B.n21 585
R88 B.n594 B.n593 585
R89 B.n595 B.n20 585
R90 B.n597 B.n596 585
R91 B.n598 B.n19 585
R92 B.n600 B.n599 585
R93 B.n459 B.n458 585
R94 B.n457 B.n70 585
R95 B.n456 B.n455 585
R96 B.n454 B.n71 585
R97 B.n453 B.n452 585
R98 B.n451 B.n72 585
R99 B.n450 B.n449 585
R100 B.n448 B.n73 585
R101 B.n447 B.n446 585
R102 B.n445 B.n74 585
R103 B.n444 B.n443 585
R104 B.n442 B.n75 585
R105 B.n441 B.n440 585
R106 B.n439 B.n76 585
R107 B.n438 B.n437 585
R108 B.n436 B.n77 585
R109 B.n435 B.n434 585
R110 B.n433 B.n78 585
R111 B.n432 B.n431 585
R112 B.n430 B.n79 585
R113 B.n429 B.n428 585
R114 B.n427 B.n80 585
R115 B.n426 B.n425 585
R116 B.n424 B.n81 585
R117 B.n423 B.n422 585
R118 B.n421 B.n82 585
R119 B.n420 B.n419 585
R120 B.n418 B.n83 585
R121 B.n417 B.n416 585
R122 B.n415 B.n84 585
R123 B.n414 B.n413 585
R124 B.n412 B.n85 585
R125 B.n411 B.n410 585
R126 B.n409 B.n86 585
R127 B.n408 B.n407 585
R128 B.n406 B.n87 585
R129 B.n405 B.n404 585
R130 B.n403 B.n88 585
R131 B.n402 B.n401 585
R132 B.n400 B.n89 585
R133 B.n399 B.n398 585
R134 B.n397 B.n90 585
R135 B.n396 B.n395 585
R136 B.n394 B.n91 585
R137 B.n393 B.n392 585
R138 B.n391 B.n92 585
R139 B.n390 B.n389 585
R140 B.n388 B.n93 585
R141 B.n387 B.n386 585
R142 B.n385 B.n94 585
R143 B.n384 B.n383 585
R144 B.n382 B.n95 585
R145 B.n381 B.n380 585
R146 B.n379 B.n96 585
R147 B.n378 B.n377 585
R148 B.n376 B.n97 585
R149 B.n375 B.n374 585
R150 B.n373 B.n98 585
R151 B.n372 B.n371 585
R152 B.n370 B.n99 585
R153 B.n369 B.n368 585
R154 B.n367 B.n100 585
R155 B.n366 B.n365 585
R156 B.n364 B.n101 585
R157 B.n363 B.n362 585
R158 B.n361 B.n102 585
R159 B.n360 B.n359 585
R160 B.n219 B.n218 585
R161 B.n220 B.n153 585
R162 B.n222 B.n221 585
R163 B.n223 B.n152 585
R164 B.n225 B.n224 585
R165 B.n226 B.n151 585
R166 B.n228 B.n227 585
R167 B.n229 B.n150 585
R168 B.n231 B.n230 585
R169 B.n232 B.n149 585
R170 B.n234 B.n233 585
R171 B.n235 B.n148 585
R172 B.n237 B.n236 585
R173 B.n238 B.n147 585
R174 B.n240 B.n239 585
R175 B.n241 B.n146 585
R176 B.n243 B.n242 585
R177 B.n244 B.n145 585
R178 B.n246 B.n245 585
R179 B.n247 B.n144 585
R180 B.n249 B.n248 585
R181 B.n250 B.n143 585
R182 B.n252 B.n251 585
R183 B.n253 B.n142 585
R184 B.n255 B.n254 585
R185 B.n256 B.n141 585
R186 B.n258 B.n257 585
R187 B.n259 B.n140 585
R188 B.n261 B.n260 585
R189 B.n262 B.n139 585
R190 B.n264 B.n263 585
R191 B.n265 B.n138 585
R192 B.n267 B.n266 585
R193 B.n268 B.n137 585
R194 B.n270 B.n269 585
R195 B.n271 B.n136 585
R196 B.n273 B.n272 585
R197 B.n274 B.n135 585
R198 B.n276 B.n275 585
R199 B.n277 B.n134 585
R200 B.n279 B.n278 585
R201 B.n280 B.n131 585
R202 B.n283 B.n282 585
R203 B.n284 B.n130 585
R204 B.n286 B.n285 585
R205 B.n287 B.n129 585
R206 B.n289 B.n288 585
R207 B.n290 B.n128 585
R208 B.n292 B.n291 585
R209 B.n293 B.n127 585
R210 B.n295 B.n294 585
R211 B.n297 B.n296 585
R212 B.n298 B.n123 585
R213 B.n300 B.n299 585
R214 B.n301 B.n122 585
R215 B.n303 B.n302 585
R216 B.n304 B.n121 585
R217 B.n306 B.n305 585
R218 B.n307 B.n120 585
R219 B.n309 B.n308 585
R220 B.n310 B.n119 585
R221 B.n312 B.n311 585
R222 B.n313 B.n118 585
R223 B.n315 B.n314 585
R224 B.n316 B.n117 585
R225 B.n318 B.n317 585
R226 B.n319 B.n116 585
R227 B.n321 B.n320 585
R228 B.n322 B.n115 585
R229 B.n324 B.n323 585
R230 B.n325 B.n114 585
R231 B.n327 B.n326 585
R232 B.n328 B.n113 585
R233 B.n330 B.n329 585
R234 B.n331 B.n112 585
R235 B.n333 B.n332 585
R236 B.n334 B.n111 585
R237 B.n336 B.n335 585
R238 B.n337 B.n110 585
R239 B.n339 B.n338 585
R240 B.n340 B.n109 585
R241 B.n342 B.n341 585
R242 B.n343 B.n108 585
R243 B.n345 B.n344 585
R244 B.n346 B.n107 585
R245 B.n348 B.n347 585
R246 B.n349 B.n106 585
R247 B.n351 B.n350 585
R248 B.n352 B.n105 585
R249 B.n354 B.n353 585
R250 B.n355 B.n104 585
R251 B.n357 B.n356 585
R252 B.n358 B.n103 585
R253 B.n217 B.n154 585
R254 B.n216 B.n215 585
R255 B.n214 B.n155 585
R256 B.n213 B.n212 585
R257 B.n211 B.n156 585
R258 B.n210 B.n209 585
R259 B.n208 B.n157 585
R260 B.n207 B.n206 585
R261 B.n205 B.n158 585
R262 B.n204 B.n203 585
R263 B.n202 B.n159 585
R264 B.n201 B.n200 585
R265 B.n199 B.n160 585
R266 B.n198 B.n197 585
R267 B.n196 B.n161 585
R268 B.n195 B.n194 585
R269 B.n193 B.n162 585
R270 B.n192 B.n191 585
R271 B.n190 B.n163 585
R272 B.n189 B.n188 585
R273 B.n187 B.n164 585
R274 B.n186 B.n185 585
R275 B.n184 B.n165 585
R276 B.n183 B.n182 585
R277 B.n181 B.n166 585
R278 B.n180 B.n179 585
R279 B.n178 B.n167 585
R280 B.n177 B.n176 585
R281 B.n175 B.n168 585
R282 B.n174 B.n173 585
R283 B.n172 B.n169 585
R284 B.n171 B.n170 585
R285 B.n2 B.n0 585
R286 B.n649 B.n1 585
R287 B.n648 B.n647 585
R288 B.n646 B.n3 585
R289 B.n645 B.n644 585
R290 B.n643 B.n4 585
R291 B.n642 B.n641 585
R292 B.n640 B.n5 585
R293 B.n639 B.n638 585
R294 B.n637 B.n6 585
R295 B.n636 B.n635 585
R296 B.n634 B.n7 585
R297 B.n633 B.n632 585
R298 B.n631 B.n8 585
R299 B.n630 B.n629 585
R300 B.n628 B.n9 585
R301 B.n627 B.n626 585
R302 B.n625 B.n10 585
R303 B.n624 B.n623 585
R304 B.n622 B.n11 585
R305 B.n621 B.n620 585
R306 B.n619 B.n12 585
R307 B.n618 B.n617 585
R308 B.n616 B.n13 585
R309 B.n615 B.n614 585
R310 B.n613 B.n14 585
R311 B.n612 B.n611 585
R312 B.n610 B.n15 585
R313 B.n609 B.n608 585
R314 B.n607 B.n16 585
R315 B.n606 B.n605 585
R316 B.n604 B.n17 585
R317 B.n603 B.n602 585
R318 B.n601 B.n18 585
R319 B.n651 B.n650 585
R320 B.n218 B.n217 468.476
R321 B.n601 B.n600 468.476
R322 B.n360 B.n103 468.476
R323 B.n458 B.n69 468.476
R324 B.n124 B.t8 429.639
R325 B.n46 B.t10 429.639
R326 B.n132 B.t2 429.639
R327 B.n40 B.t4 429.639
R328 B.n125 B.t7 374.949
R329 B.n47 B.t11 374.949
R330 B.n133 B.t1 374.949
R331 B.n41 B.t5 374.949
R332 B.n124 B.t6 323.729
R333 B.n132 B.t0 323.729
R334 B.n40 B.t3 323.729
R335 B.n46 B.t9 323.729
R336 B.n217 B.n216 163.367
R337 B.n216 B.n155 163.367
R338 B.n212 B.n155 163.367
R339 B.n212 B.n211 163.367
R340 B.n211 B.n210 163.367
R341 B.n210 B.n157 163.367
R342 B.n206 B.n157 163.367
R343 B.n206 B.n205 163.367
R344 B.n205 B.n204 163.367
R345 B.n204 B.n159 163.367
R346 B.n200 B.n159 163.367
R347 B.n200 B.n199 163.367
R348 B.n199 B.n198 163.367
R349 B.n198 B.n161 163.367
R350 B.n194 B.n161 163.367
R351 B.n194 B.n193 163.367
R352 B.n193 B.n192 163.367
R353 B.n192 B.n163 163.367
R354 B.n188 B.n163 163.367
R355 B.n188 B.n187 163.367
R356 B.n187 B.n186 163.367
R357 B.n186 B.n165 163.367
R358 B.n182 B.n165 163.367
R359 B.n182 B.n181 163.367
R360 B.n181 B.n180 163.367
R361 B.n180 B.n167 163.367
R362 B.n176 B.n167 163.367
R363 B.n176 B.n175 163.367
R364 B.n175 B.n174 163.367
R365 B.n174 B.n169 163.367
R366 B.n170 B.n169 163.367
R367 B.n170 B.n2 163.367
R368 B.n650 B.n2 163.367
R369 B.n650 B.n649 163.367
R370 B.n649 B.n648 163.367
R371 B.n648 B.n3 163.367
R372 B.n644 B.n3 163.367
R373 B.n644 B.n643 163.367
R374 B.n643 B.n642 163.367
R375 B.n642 B.n5 163.367
R376 B.n638 B.n5 163.367
R377 B.n638 B.n637 163.367
R378 B.n637 B.n636 163.367
R379 B.n636 B.n7 163.367
R380 B.n632 B.n7 163.367
R381 B.n632 B.n631 163.367
R382 B.n631 B.n630 163.367
R383 B.n630 B.n9 163.367
R384 B.n626 B.n9 163.367
R385 B.n626 B.n625 163.367
R386 B.n625 B.n624 163.367
R387 B.n624 B.n11 163.367
R388 B.n620 B.n11 163.367
R389 B.n620 B.n619 163.367
R390 B.n619 B.n618 163.367
R391 B.n618 B.n13 163.367
R392 B.n614 B.n13 163.367
R393 B.n614 B.n613 163.367
R394 B.n613 B.n612 163.367
R395 B.n612 B.n15 163.367
R396 B.n608 B.n15 163.367
R397 B.n608 B.n607 163.367
R398 B.n607 B.n606 163.367
R399 B.n606 B.n17 163.367
R400 B.n602 B.n17 163.367
R401 B.n602 B.n601 163.367
R402 B.n218 B.n153 163.367
R403 B.n222 B.n153 163.367
R404 B.n223 B.n222 163.367
R405 B.n224 B.n223 163.367
R406 B.n224 B.n151 163.367
R407 B.n228 B.n151 163.367
R408 B.n229 B.n228 163.367
R409 B.n230 B.n229 163.367
R410 B.n230 B.n149 163.367
R411 B.n234 B.n149 163.367
R412 B.n235 B.n234 163.367
R413 B.n236 B.n235 163.367
R414 B.n236 B.n147 163.367
R415 B.n240 B.n147 163.367
R416 B.n241 B.n240 163.367
R417 B.n242 B.n241 163.367
R418 B.n242 B.n145 163.367
R419 B.n246 B.n145 163.367
R420 B.n247 B.n246 163.367
R421 B.n248 B.n247 163.367
R422 B.n248 B.n143 163.367
R423 B.n252 B.n143 163.367
R424 B.n253 B.n252 163.367
R425 B.n254 B.n253 163.367
R426 B.n254 B.n141 163.367
R427 B.n258 B.n141 163.367
R428 B.n259 B.n258 163.367
R429 B.n260 B.n259 163.367
R430 B.n260 B.n139 163.367
R431 B.n264 B.n139 163.367
R432 B.n265 B.n264 163.367
R433 B.n266 B.n265 163.367
R434 B.n266 B.n137 163.367
R435 B.n270 B.n137 163.367
R436 B.n271 B.n270 163.367
R437 B.n272 B.n271 163.367
R438 B.n272 B.n135 163.367
R439 B.n276 B.n135 163.367
R440 B.n277 B.n276 163.367
R441 B.n278 B.n277 163.367
R442 B.n278 B.n131 163.367
R443 B.n283 B.n131 163.367
R444 B.n284 B.n283 163.367
R445 B.n285 B.n284 163.367
R446 B.n285 B.n129 163.367
R447 B.n289 B.n129 163.367
R448 B.n290 B.n289 163.367
R449 B.n291 B.n290 163.367
R450 B.n291 B.n127 163.367
R451 B.n295 B.n127 163.367
R452 B.n296 B.n295 163.367
R453 B.n296 B.n123 163.367
R454 B.n300 B.n123 163.367
R455 B.n301 B.n300 163.367
R456 B.n302 B.n301 163.367
R457 B.n302 B.n121 163.367
R458 B.n306 B.n121 163.367
R459 B.n307 B.n306 163.367
R460 B.n308 B.n307 163.367
R461 B.n308 B.n119 163.367
R462 B.n312 B.n119 163.367
R463 B.n313 B.n312 163.367
R464 B.n314 B.n313 163.367
R465 B.n314 B.n117 163.367
R466 B.n318 B.n117 163.367
R467 B.n319 B.n318 163.367
R468 B.n320 B.n319 163.367
R469 B.n320 B.n115 163.367
R470 B.n324 B.n115 163.367
R471 B.n325 B.n324 163.367
R472 B.n326 B.n325 163.367
R473 B.n326 B.n113 163.367
R474 B.n330 B.n113 163.367
R475 B.n331 B.n330 163.367
R476 B.n332 B.n331 163.367
R477 B.n332 B.n111 163.367
R478 B.n336 B.n111 163.367
R479 B.n337 B.n336 163.367
R480 B.n338 B.n337 163.367
R481 B.n338 B.n109 163.367
R482 B.n342 B.n109 163.367
R483 B.n343 B.n342 163.367
R484 B.n344 B.n343 163.367
R485 B.n344 B.n107 163.367
R486 B.n348 B.n107 163.367
R487 B.n349 B.n348 163.367
R488 B.n350 B.n349 163.367
R489 B.n350 B.n105 163.367
R490 B.n354 B.n105 163.367
R491 B.n355 B.n354 163.367
R492 B.n356 B.n355 163.367
R493 B.n356 B.n103 163.367
R494 B.n361 B.n360 163.367
R495 B.n362 B.n361 163.367
R496 B.n362 B.n101 163.367
R497 B.n366 B.n101 163.367
R498 B.n367 B.n366 163.367
R499 B.n368 B.n367 163.367
R500 B.n368 B.n99 163.367
R501 B.n372 B.n99 163.367
R502 B.n373 B.n372 163.367
R503 B.n374 B.n373 163.367
R504 B.n374 B.n97 163.367
R505 B.n378 B.n97 163.367
R506 B.n379 B.n378 163.367
R507 B.n380 B.n379 163.367
R508 B.n380 B.n95 163.367
R509 B.n384 B.n95 163.367
R510 B.n385 B.n384 163.367
R511 B.n386 B.n385 163.367
R512 B.n386 B.n93 163.367
R513 B.n390 B.n93 163.367
R514 B.n391 B.n390 163.367
R515 B.n392 B.n391 163.367
R516 B.n392 B.n91 163.367
R517 B.n396 B.n91 163.367
R518 B.n397 B.n396 163.367
R519 B.n398 B.n397 163.367
R520 B.n398 B.n89 163.367
R521 B.n402 B.n89 163.367
R522 B.n403 B.n402 163.367
R523 B.n404 B.n403 163.367
R524 B.n404 B.n87 163.367
R525 B.n408 B.n87 163.367
R526 B.n409 B.n408 163.367
R527 B.n410 B.n409 163.367
R528 B.n410 B.n85 163.367
R529 B.n414 B.n85 163.367
R530 B.n415 B.n414 163.367
R531 B.n416 B.n415 163.367
R532 B.n416 B.n83 163.367
R533 B.n420 B.n83 163.367
R534 B.n421 B.n420 163.367
R535 B.n422 B.n421 163.367
R536 B.n422 B.n81 163.367
R537 B.n426 B.n81 163.367
R538 B.n427 B.n426 163.367
R539 B.n428 B.n427 163.367
R540 B.n428 B.n79 163.367
R541 B.n432 B.n79 163.367
R542 B.n433 B.n432 163.367
R543 B.n434 B.n433 163.367
R544 B.n434 B.n77 163.367
R545 B.n438 B.n77 163.367
R546 B.n439 B.n438 163.367
R547 B.n440 B.n439 163.367
R548 B.n440 B.n75 163.367
R549 B.n444 B.n75 163.367
R550 B.n445 B.n444 163.367
R551 B.n446 B.n445 163.367
R552 B.n446 B.n73 163.367
R553 B.n450 B.n73 163.367
R554 B.n451 B.n450 163.367
R555 B.n452 B.n451 163.367
R556 B.n452 B.n71 163.367
R557 B.n456 B.n71 163.367
R558 B.n457 B.n456 163.367
R559 B.n458 B.n457 163.367
R560 B.n600 B.n19 163.367
R561 B.n596 B.n19 163.367
R562 B.n596 B.n595 163.367
R563 B.n595 B.n594 163.367
R564 B.n594 B.n21 163.367
R565 B.n590 B.n21 163.367
R566 B.n590 B.n589 163.367
R567 B.n589 B.n588 163.367
R568 B.n588 B.n23 163.367
R569 B.n584 B.n23 163.367
R570 B.n584 B.n583 163.367
R571 B.n583 B.n582 163.367
R572 B.n582 B.n25 163.367
R573 B.n578 B.n25 163.367
R574 B.n578 B.n577 163.367
R575 B.n577 B.n576 163.367
R576 B.n576 B.n27 163.367
R577 B.n572 B.n27 163.367
R578 B.n572 B.n571 163.367
R579 B.n571 B.n570 163.367
R580 B.n570 B.n29 163.367
R581 B.n566 B.n29 163.367
R582 B.n566 B.n565 163.367
R583 B.n565 B.n564 163.367
R584 B.n564 B.n31 163.367
R585 B.n560 B.n31 163.367
R586 B.n560 B.n559 163.367
R587 B.n559 B.n558 163.367
R588 B.n558 B.n33 163.367
R589 B.n554 B.n33 163.367
R590 B.n554 B.n553 163.367
R591 B.n553 B.n552 163.367
R592 B.n552 B.n35 163.367
R593 B.n548 B.n35 163.367
R594 B.n548 B.n547 163.367
R595 B.n547 B.n546 163.367
R596 B.n546 B.n37 163.367
R597 B.n542 B.n37 163.367
R598 B.n542 B.n541 163.367
R599 B.n541 B.n540 163.367
R600 B.n540 B.n39 163.367
R601 B.n535 B.n39 163.367
R602 B.n535 B.n534 163.367
R603 B.n534 B.n533 163.367
R604 B.n533 B.n43 163.367
R605 B.n529 B.n43 163.367
R606 B.n529 B.n528 163.367
R607 B.n528 B.n527 163.367
R608 B.n527 B.n45 163.367
R609 B.n523 B.n45 163.367
R610 B.n523 B.n522 163.367
R611 B.n522 B.n49 163.367
R612 B.n518 B.n49 163.367
R613 B.n518 B.n517 163.367
R614 B.n517 B.n516 163.367
R615 B.n516 B.n51 163.367
R616 B.n512 B.n51 163.367
R617 B.n512 B.n511 163.367
R618 B.n511 B.n510 163.367
R619 B.n510 B.n53 163.367
R620 B.n506 B.n53 163.367
R621 B.n506 B.n505 163.367
R622 B.n505 B.n504 163.367
R623 B.n504 B.n55 163.367
R624 B.n500 B.n55 163.367
R625 B.n500 B.n499 163.367
R626 B.n499 B.n498 163.367
R627 B.n498 B.n57 163.367
R628 B.n494 B.n57 163.367
R629 B.n494 B.n493 163.367
R630 B.n493 B.n492 163.367
R631 B.n492 B.n59 163.367
R632 B.n488 B.n59 163.367
R633 B.n488 B.n487 163.367
R634 B.n487 B.n486 163.367
R635 B.n486 B.n61 163.367
R636 B.n482 B.n61 163.367
R637 B.n482 B.n481 163.367
R638 B.n481 B.n480 163.367
R639 B.n480 B.n63 163.367
R640 B.n476 B.n63 163.367
R641 B.n476 B.n475 163.367
R642 B.n475 B.n474 163.367
R643 B.n474 B.n65 163.367
R644 B.n470 B.n65 163.367
R645 B.n470 B.n469 163.367
R646 B.n469 B.n468 163.367
R647 B.n468 B.n67 163.367
R648 B.n464 B.n67 163.367
R649 B.n464 B.n463 163.367
R650 B.n463 B.n462 163.367
R651 B.n462 B.n69 163.367
R652 B.n126 B.n125 59.5399
R653 B.n281 B.n133 59.5399
R654 B.n537 B.n41 59.5399
R655 B.n48 B.n47 59.5399
R656 B.n125 B.n124 54.6914
R657 B.n133 B.n132 54.6914
R658 B.n41 B.n40 54.6914
R659 B.n47 B.n46 54.6914
R660 B.n599 B.n18 30.4395
R661 B.n460 B.n459 30.4395
R662 B.n359 B.n358 30.4395
R663 B.n219 B.n154 30.4395
R664 B B.n651 18.0485
R665 B.n599 B.n598 10.6151
R666 B.n598 B.n597 10.6151
R667 B.n597 B.n20 10.6151
R668 B.n593 B.n20 10.6151
R669 B.n593 B.n592 10.6151
R670 B.n592 B.n591 10.6151
R671 B.n591 B.n22 10.6151
R672 B.n587 B.n22 10.6151
R673 B.n587 B.n586 10.6151
R674 B.n586 B.n585 10.6151
R675 B.n585 B.n24 10.6151
R676 B.n581 B.n24 10.6151
R677 B.n581 B.n580 10.6151
R678 B.n580 B.n579 10.6151
R679 B.n579 B.n26 10.6151
R680 B.n575 B.n26 10.6151
R681 B.n575 B.n574 10.6151
R682 B.n574 B.n573 10.6151
R683 B.n573 B.n28 10.6151
R684 B.n569 B.n28 10.6151
R685 B.n569 B.n568 10.6151
R686 B.n568 B.n567 10.6151
R687 B.n567 B.n30 10.6151
R688 B.n563 B.n30 10.6151
R689 B.n563 B.n562 10.6151
R690 B.n562 B.n561 10.6151
R691 B.n561 B.n32 10.6151
R692 B.n557 B.n32 10.6151
R693 B.n557 B.n556 10.6151
R694 B.n556 B.n555 10.6151
R695 B.n555 B.n34 10.6151
R696 B.n551 B.n34 10.6151
R697 B.n551 B.n550 10.6151
R698 B.n550 B.n549 10.6151
R699 B.n549 B.n36 10.6151
R700 B.n545 B.n36 10.6151
R701 B.n545 B.n544 10.6151
R702 B.n544 B.n543 10.6151
R703 B.n543 B.n38 10.6151
R704 B.n539 B.n38 10.6151
R705 B.n539 B.n538 10.6151
R706 B.n536 B.n42 10.6151
R707 B.n532 B.n42 10.6151
R708 B.n532 B.n531 10.6151
R709 B.n531 B.n530 10.6151
R710 B.n530 B.n44 10.6151
R711 B.n526 B.n44 10.6151
R712 B.n526 B.n525 10.6151
R713 B.n525 B.n524 10.6151
R714 B.n521 B.n520 10.6151
R715 B.n520 B.n519 10.6151
R716 B.n519 B.n50 10.6151
R717 B.n515 B.n50 10.6151
R718 B.n515 B.n514 10.6151
R719 B.n514 B.n513 10.6151
R720 B.n513 B.n52 10.6151
R721 B.n509 B.n52 10.6151
R722 B.n509 B.n508 10.6151
R723 B.n508 B.n507 10.6151
R724 B.n507 B.n54 10.6151
R725 B.n503 B.n54 10.6151
R726 B.n503 B.n502 10.6151
R727 B.n502 B.n501 10.6151
R728 B.n501 B.n56 10.6151
R729 B.n497 B.n56 10.6151
R730 B.n497 B.n496 10.6151
R731 B.n496 B.n495 10.6151
R732 B.n495 B.n58 10.6151
R733 B.n491 B.n58 10.6151
R734 B.n491 B.n490 10.6151
R735 B.n490 B.n489 10.6151
R736 B.n489 B.n60 10.6151
R737 B.n485 B.n60 10.6151
R738 B.n485 B.n484 10.6151
R739 B.n484 B.n483 10.6151
R740 B.n483 B.n62 10.6151
R741 B.n479 B.n62 10.6151
R742 B.n479 B.n478 10.6151
R743 B.n478 B.n477 10.6151
R744 B.n477 B.n64 10.6151
R745 B.n473 B.n64 10.6151
R746 B.n473 B.n472 10.6151
R747 B.n472 B.n471 10.6151
R748 B.n471 B.n66 10.6151
R749 B.n467 B.n66 10.6151
R750 B.n467 B.n466 10.6151
R751 B.n466 B.n465 10.6151
R752 B.n465 B.n68 10.6151
R753 B.n461 B.n68 10.6151
R754 B.n461 B.n460 10.6151
R755 B.n359 B.n102 10.6151
R756 B.n363 B.n102 10.6151
R757 B.n364 B.n363 10.6151
R758 B.n365 B.n364 10.6151
R759 B.n365 B.n100 10.6151
R760 B.n369 B.n100 10.6151
R761 B.n370 B.n369 10.6151
R762 B.n371 B.n370 10.6151
R763 B.n371 B.n98 10.6151
R764 B.n375 B.n98 10.6151
R765 B.n376 B.n375 10.6151
R766 B.n377 B.n376 10.6151
R767 B.n377 B.n96 10.6151
R768 B.n381 B.n96 10.6151
R769 B.n382 B.n381 10.6151
R770 B.n383 B.n382 10.6151
R771 B.n383 B.n94 10.6151
R772 B.n387 B.n94 10.6151
R773 B.n388 B.n387 10.6151
R774 B.n389 B.n388 10.6151
R775 B.n389 B.n92 10.6151
R776 B.n393 B.n92 10.6151
R777 B.n394 B.n393 10.6151
R778 B.n395 B.n394 10.6151
R779 B.n395 B.n90 10.6151
R780 B.n399 B.n90 10.6151
R781 B.n400 B.n399 10.6151
R782 B.n401 B.n400 10.6151
R783 B.n401 B.n88 10.6151
R784 B.n405 B.n88 10.6151
R785 B.n406 B.n405 10.6151
R786 B.n407 B.n406 10.6151
R787 B.n407 B.n86 10.6151
R788 B.n411 B.n86 10.6151
R789 B.n412 B.n411 10.6151
R790 B.n413 B.n412 10.6151
R791 B.n413 B.n84 10.6151
R792 B.n417 B.n84 10.6151
R793 B.n418 B.n417 10.6151
R794 B.n419 B.n418 10.6151
R795 B.n419 B.n82 10.6151
R796 B.n423 B.n82 10.6151
R797 B.n424 B.n423 10.6151
R798 B.n425 B.n424 10.6151
R799 B.n425 B.n80 10.6151
R800 B.n429 B.n80 10.6151
R801 B.n430 B.n429 10.6151
R802 B.n431 B.n430 10.6151
R803 B.n431 B.n78 10.6151
R804 B.n435 B.n78 10.6151
R805 B.n436 B.n435 10.6151
R806 B.n437 B.n436 10.6151
R807 B.n437 B.n76 10.6151
R808 B.n441 B.n76 10.6151
R809 B.n442 B.n441 10.6151
R810 B.n443 B.n442 10.6151
R811 B.n443 B.n74 10.6151
R812 B.n447 B.n74 10.6151
R813 B.n448 B.n447 10.6151
R814 B.n449 B.n448 10.6151
R815 B.n449 B.n72 10.6151
R816 B.n453 B.n72 10.6151
R817 B.n454 B.n453 10.6151
R818 B.n455 B.n454 10.6151
R819 B.n455 B.n70 10.6151
R820 B.n459 B.n70 10.6151
R821 B.n220 B.n219 10.6151
R822 B.n221 B.n220 10.6151
R823 B.n221 B.n152 10.6151
R824 B.n225 B.n152 10.6151
R825 B.n226 B.n225 10.6151
R826 B.n227 B.n226 10.6151
R827 B.n227 B.n150 10.6151
R828 B.n231 B.n150 10.6151
R829 B.n232 B.n231 10.6151
R830 B.n233 B.n232 10.6151
R831 B.n233 B.n148 10.6151
R832 B.n237 B.n148 10.6151
R833 B.n238 B.n237 10.6151
R834 B.n239 B.n238 10.6151
R835 B.n239 B.n146 10.6151
R836 B.n243 B.n146 10.6151
R837 B.n244 B.n243 10.6151
R838 B.n245 B.n244 10.6151
R839 B.n245 B.n144 10.6151
R840 B.n249 B.n144 10.6151
R841 B.n250 B.n249 10.6151
R842 B.n251 B.n250 10.6151
R843 B.n251 B.n142 10.6151
R844 B.n255 B.n142 10.6151
R845 B.n256 B.n255 10.6151
R846 B.n257 B.n256 10.6151
R847 B.n257 B.n140 10.6151
R848 B.n261 B.n140 10.6151
R849 B.n262 B.n261 10.6151
R850 B.n263 B.n262 10.6151
R851 B.n263 B.n138 10.6151
R852 B.n267 B.n138 10.6151
R853 B.n268 B.n267 10.6151
R854 B.n269 B.n268 10.6151
R855 B.n269 B.n136 10.6151
R856 B.n273 B.n136 10.6151
R857 B.n274 B.n273 10.6151
R858 B.n275 B.n274 10.6151
R859 B.n275 B.n134 10.6151
R860 B.n279 B.n134 10.6151
R861 B.n280 B.n279 10.6151
R862 B.n282 B.n130 10.6151
R863 B.n286 B.n130 10.6151
R864 B.n287 B.n286 10.6151
R865 B.n288 B.n287 10.6151
R866 B.n288 B.n128 10.6151
R867 B.n292 B.n128 10.6151
R868 B.n293 B.n292 10.6151
R869 B.n294 B.n293 10.6151
R870 B.n298 B.n297 10.6151
R871 B.n299 B.n298 10.6151
R872 B.n299 B.n122 10.6151
R873 B.n303 B.n122 10.6151
R874 B.n304 B.n303 10.6151
R875 B.n305 B.n304 10.6151
R876 B.n305 B.n120 10.6151
R877 B.n309 B.n120 10.6151
R878 B.n310 B.n309 10.6151
R879 B.n311 B.n310 10.6151
R880 B.n311 B.n118 10.6151
R881 B.n315 B.n118 10.6151
R882 B.n316 B.n315 10.6151
R883 B.n317 B.n316 10.6151
R884 B.n317 B.n116 10.6151
R885 B.n321 B.n116 10.6151
R886 B.n322 B.n321 10.6151
R887 B.n323 B.n322 10.6151
R888 B.n323 B.n114 10.6151
R889 B.n327 B.n114 10.6151
R890 B.n328 B.n327 10.6151
R891 B.n329 B.n328 10.6151
R892 B.n329 B.n112 10.6151
R893 B.n333 B.n112 10.6151
R894 B.n334 B.n333 10.6151
R895 B.n335 B.n334 10.6151
R896 B.n335 B.n110 10.6151
R897 B.n339 B.n110 10.6151
R898 B.n340 B.n339 10.6151
R899 B.n341 B.n340 10.6151
R900 B.n341 B.n108 10.6151
R901 B.n345 B.n108 10.6151
R902 B.n346 B.n345 10.6151
R903 B.n347 B.n346 10.6151
R904 B.n347 B.n106 10.6151
R905 B.n351 B.n106 10.6151
R906 B.n352 B.n351 10.6151
R907 B.n353 B.n352 10.6151
R908 B.n353 B.n104 10.6151
R909 B.n357 B.n104 10.6151
R910 B.n358 B.n357 10.6151
R911 B.n215 B.n154 10.6151
R912 B.n215 B.n214 10.6151
R913 B.n214 B.n213 10.6151
R914 B.n213 B.n156 10.6151
R915 B.n209 B.n156 10.6151
R916 B.n209 B.n208 10.6151
R917 B.n208 B.n207 10.6151
R918 B.n207 B.n158 10.6151
R919 B.n203 B.n158 10.6151
R920 B.n203 B.n202 10.6151
R921 B.n202 B.n201 10.6151
R922 B.n201 B.n160 10.6151
R923 B.n197 B.n160 10.6151
R924 B.n197 B.n196 10.6151
R925 B.n196 B.n195 10.6151
R926 B.n195 B.n162 10.6151
R927 B.n191 B.n162 10.6151
R928 B.n191 B.n190 10.6151
R929 B.n190 B.n189 10.6151
R930 B.n189 B.n164 10.6151
R931 B.n185 B.n164 10.6151
R932 B.n185 B.n184 10.6151
R933 B.n184 B.n183 10.6151
R934 B.n183 B.n166 10.6151
R935 B.n179 B.n166 10.6151
R936 B.n179 B.n178 10.6151
R937 B.n178 B.n177 10.6151
R938 B.n177 B.n168 10.6151
R939 B.n173 B.n168 10.6151
R940 B.n173 B.n172 10.6151
R941 B.n172 B.n171 10.6151
R942 B.n171 B.n0 10.6151
R943 B.n647 B.n1 10.6151
R944 B.n647 B.n646 10.6151
R945 B.n646 B.n645 10.6151
R946 B.n645 B.n4 10.6151
R947 B.n641 B.n4 10.6151
R948 B.n641 B.n640 10.6151
R949 B.n640 B.n639 10.6151
R950 B.n639 B.n6 10.6151
R951 B.n635 B.n6 10.6151
R952 B.n635 B.n634 10.6151
R953 B.n634 B.n633 10.6151
R954 B.n633 B.n8 10.6151
R955 B.n629 B.n8 10.6151
R956 B.n629 B.n628 10.6151
R957 B.n628 B.n627 10.6151
R958 B.n627 B.n10 10.6151
R959 B.n623 B.n10 10.6151
R960 B.n623 B.n622 10.6151
R961 B.n622 B.n621 10.6151
R962 B.n621 B.n12 10.6151
R963 B.n617 B.n12 10.6151
R964 B.n617 B.n616 10.6151
R965 B.n616 B.n615 10.6151
R966 B.n615 B.n14 10.6151
R967 B.n611 B.n14 10.6151
R968 B.n611 B.n610 10.6151
R969 B.n610 B.n609 10.6151
R970 B.n609 B.n16 10.6151
R971 B.n605 B.n16 10.6151
R972 B.n605 B.n604 10.6151
R973 B.n604 B.n603 10.6151
R974 B.n603 B.n18 10.6151
R975 B.n537 B.n536 6.5566
R976 B.n524 B.n48 6.5566
R977 B.n282 B.n281 6.5566
R978 B.n294 B.n126 6.5566
R979 B.n538 B.n537 4.05904
R980 B.n521 B.n48 4.05904
R981 B.n281 B.n280 4.05904
R982 B.n297 B.n126 4.05904
R983 B.n651 B.n0 2.81026
R984 B.n651 B.n1 2.81026
R985 VN.n0 VN.t1 151.201
R986 VN.n1 VN.t3 151.201
R987 VN.n0 VN.t0 150.445
R988 VN.n1 VN.t2 150.445
R989 VN VN.n1 50.7193
R990 VN VN.n0 4.54889
R991 VTAIL.n526 VTAIL.n525 756.745
R992 VTAIL.n64 VTAIL.n63 756.745
R993 VTAIL.n130 VTAIL.n129 756.745
R994 VTAIL.n196 VTAIL.n195 756.745
R995 VTAIL.n460 VTAIL.n459 756.745
R996 VTAIL.n394 VTAIL.n393 756.745
R997 VTAIL.n328 VTAIL.n327 756.745
R998 VTAIL.n262 VTAIL.n261 756.745
R999 VTAIL.n485 VTAIL.n484 585
R1000 VTAIL.n487 VTAIL.n486 585
R1001 VTAIL.n480 VTAIL.n479 585
R1002 VTAIL.n493 VTAIL.n492 585
R1003 VTAIL.n495 VTAIL.n494 585
R1004 VTAIL.n476 VTAIL.n475 585
R1005 VTAIL.n501 VTAIL.n500 585
R1006 VTAIL.n503 VTAIL.n502 585
R1007 VTAIL.n472 VTAIL.n471 585
R1008 VTAIL.n509 VTAIL.n508 585
R1009 VTAIL.n511 VTAIL.n510 585
R1010 VTAIL.n468 VTAIL.n467 585
R1011 VTAIL.n517 VTAIL.n516 585
R1012 VTAIL.n519 VTAIL.n518 585
R1013 VTAIL.n464 VTAIL.n463 585
R1014 VTAIL.n525 VTAIL.n524 585
R1015 VTAIL.n23 VTAIL.n22 585
R1016 VTAIL.n25 VTAIL.n24 585
R1017 VTAIL.n18 VTAIL.n17 585
R1018 VTAIL.n31 VTAIL.n30 585
R1019 VTAIL.n33 VTAIL.n32 585
R1020 VTAIL.n14 VTAIL.n13 585
R1021 VTAIL.n39 VTAIL.n38 585
R1022 VTAIL.n41 VTAIL.n40 585
R1023 VTAIL.n10 VTAIL.n9 585
R1024 VTAIL.n47 VTAIL.n46 585
R1025 VTAIL.n49 VTAIL.n48 585
R1026 VTAIL.n6 VTAIL.n5 585
R1027 VTAIL.n55 VTAIL.n54 585
R1028 VTAIL.n57 VTAIL.n56 585
R1029 VTAIL.n2 VTAIL.n1 585
R1030 VTAIL.n63 VTAIL.n62 585
R1031 VTAIL.n89 VTAIL.n88 585
R1032 VTAIL.n91 VTAIL.n90 585
R1033 VTAIL.n84 VTAIL.n83 585
R1034 VTAIL.n97 VTAIL.n96 585
R1035 VTAIL.n99 VTAIL.n98 585
R1036 VTAIL.n80 VTAIL.n79 585
R1037 VTAIL.n105 VTAIL.n104 585
R1038 VTAIL.n107 VTAIL.n106 585
R1039 VTAIL.n76 VTAIL.n75 585
R1040 VTAIL.n113 VTAIL.n112 585
R1041 VTAIL.n115 VTAIL.n114 585
R1042 VTAIL.n72 VTAIL.n71 585
R1043 VTAIL.n121 VTAIL.n120 585
R1044 VTAIL.n123 VTAIL.n122 585
R1045 VTAIL.n68 VTAIL.n67 585
R1046 VTAIL.n129 VTAIL.n128 585
R1047 VTAIL.n155 VTAIL.n154 585
R1048 VTAIL.n157 VTAIL.n156 585
R1049 VTAIL.n150 VTAIL.n149 585
R1050 VTAIL.n163 VTAIL.n162 585
R1051 VTAIL.n165 VTAIL.n164 585
R1052 VTAIL.n146 VTAIL.n145 585
R1053 VTAIL.n171 VTAIL.n170 585
R1054 VTAIL.n173 VTAIL.n172 585
R1055 VTAIL.n142 VTAIL.n141 585
R1056 VTAIL.n179 VTAIL.n178 585
R1057 VTAIL.n181 VTAIL.n180 585
R1058 VTAIL.n138 VTAIL.n137 585
R1059 VTAIL.n187 VTAIL.n186 585
R1060 VTAIL.n189 VTAIL.n188 585
R1061 VTAIL.n134 VTAIL.n133 585
R1062 VTAIL.n195 VTAIL.n194 585
R1063 VTAIL.n459 VTAIL.n458 585
R1064 VTAIL.n398 VTAIL.n397 585
R1065 VTAIL.n453 VTAIL.n452 585
R1066 VTAIL.n451 VTAIL.n450 585
R1067 VTAIL.n402 VTAIL.n401 585
R1068 VTAIL.n445 VTAIL.n444 585
R1069 VTAIL.n443 VTAIL.n442 585
R1070 VTAIL.n406 VTAIL.n405 585
R1071 VTAIL.n437 VTAIL.n436 585
R1072 VTAIL.n435 VTAIL.n434 585
R1073 VTAIL.n410 VTAIL.n409 585
R1074 VTAIL.n429 VTAIL.n428 585
R1075 VTAIL.n427 VTAIL.n426 585
R1076 VTAIL.n414 VTAIL.n413 585
R1077 VTAIL.n421 VTAIL.n420 585
R1078 VTAIL.n419 VTAIL.n418 585
R1079 VTAIL.n393 VTAIL.n392 585
R1080 VTAIL.n332 VTAIL.n331 585
R1081 VTAIL.n387 VTAIL.n386 585
R1082 VTAIL.n385 VTAIL.n384 585
R1083 VTAIL.n336 VTAIL.n335 585
R1084 VTAIL.n379 VTAIL.n378 585
R1085 VTAIL.n377 VTAIL.n376 585
R1086 VTAIL.n340 VTAIL.n339 585
R1087 VTAIL.n371 VTAIL.n370 585
R1088 VTAIL.n369 VTAIL.n368 585
R1089 VTAIL.n344 VTAIL.n343 585
R1090 VTAIL.n363 VTAIL.n362 585
R1091 VTAIL.n361 VTAIL.n360 585
R1092 VTAIL.n348 VTAIL.n347 585
R1093 VTAIL.n355 VTAIL.n354 585
R1094 VTAIL.n353 VTAIL.n352 585
R1095 VTAIL.n327 VTAIL.n326 585
R1096 VTAIL.n266 VTAIL.n265 585
R1097 VTAIL.n321 VTAIL.n320 585
R1098 VTAIL.n319 VTAIL.n318 585
R1099 VTAIL.n270 VTAIL.n269 585
R1100 VTAIL.n313 VTAIL.n312 585
R1101 VTAIL.n311 VTAIL.n310 585
R1102 VTAIL.n274 VTAIL.n273 585
R1103 VTAIL.n305 VTAIL.n304 585
R1104 VTAIL.n303 VTAIL.n302 585
R1105 VTAIL.n278 VTAIL.n277 585
R1106 VTAIL.n297 VTAIL.n296 585
R1107 VTAIL.n295 VTAIL.n294 585
R1108 VTAIL.n282 VTAIL.n281 585
R1109 VTAIL.n289 VTAIL.n288 585
R1110 VTAIL.n287 VTAIL.n286 585
R1111 VTAIL.n261 VTAIL.n260 585
R1112 VTAIL.n200 VTAIL.n199 585
R1113 VTAIL.n255 VTAIL.n254 585
R1114 VTAIL.n253 VTAIL.n252 585
R1115 VTAIL.n204 VTAIL.n203 585
R1116 VTAIL.n247 VTAIL.n246 585
R1117 VTAIL.n245 VTAIL.n244 585
R1118 VTAIL.n208 VTAIL.n207 585
R1119 VTAIL.n239 VTAIL.n238 585
R1120 VTAIL.n237 VTAIL.n236 585
R1121 VTAIL.n212 VTAIL.n211 585
R1122 VTAIL.n231 VTAIL.n230 585
R1123 VTAIL.n229 VTAIL.n228 585
R1124 VTAIL.n216 VTAIL.n215 585
R1125 VTAIL.n223 VTAIL.n222 585
R1126 VTAIL.n221 VTAIL.n220 585
R1127 VTAIL.n417 VTAIL.t3 327.466
R1128 VTAIL.n351 VTAIL.t1 327.466
R1129 VTAIL.n285 VTAIL.t6 327.466
R1130 VTAIL.n219 VTAIL.t4 327.466
R1131 VTAIL.n483 VTAIL.t5 327.466
R1132 VTAIL.n21 VTAIL.t7 327.466
R1133 VTAIL.n87 VTAIL.t0 327.466
R1134 VTAIL.n153 VTAIL.t2 327.466
R1135 VTAIL.n486 VTAIL.n485 171.744
R1136 VTAIL.n486 VTAIL.n479 171.744
R1137 VTAIL.n493 VTAIL.n479 171.744
R1138 VTAIL.n494 VTAIL.n493 171.744
R1139 VTAIL.n494 VTAIL.n475 171.744
R1140 VTAIL.n501 VTAIL.n475 171.744
R1141 VTAIL.n502 VTAIL.n501 171.744
R1142 VTAIL.n502 VTAIL.n471 171.744
R1143 VTAIL.n509 VTAIL.n471 171.744
R1144 VTAIL.n510 VTAIL.n509 171.744
R1145 VTAIL.n510 VTAIL.n467 171.744
R1146 VTAIL.n517 VTAIL.n467 171.744
R1147 VTAIL.n518 VTAIL.n517 171.744
R1148 VTAIL.n518 VTAIL.n463 171.744
R1149 VTAIL.n525 VTAIL.n463 171.744
R1150 VTAIL.n24 VTAIL.n23 171.744
R1151 VTAIL.n24 VTAIL.n17 171.744
R1152 VTAIL.n31 VTAIL.n17 171.744
R1153 VTAIL.n32 VTAIL.n31 171.744
R1154 VTAIL.n32 VTAIL.n13 171.744
R1155 VTAIL.n39 VTAIL.n13 171.744
R1156 VTAIL.n40 VTAIL.n39 171.744
R1157 VTAIL.n40 VTAIL.n9 171.744
R1158 VTAIL.n47 VTAIL.n9 171.744
R1159 VTAIL.n48 VTAIL.n47 171.744
R1160 VTAIL.n48 VTAIL.n5 171.744
R1161 VTAIL.n55 VTAIL.n5 171.744
R1162 VTAIL.n56 VTAIL.n55 171.744
R1163 VTAIL.n56 VTAIL.n1 171.744
R1164 VTAIL.n63 VTAIL.n1 171.744
R1165 VTAIL.n90 VTAIL.n89 171.744
R1166 VTAIL.n90 VTAIL.n83 171.744
R1167 VTAIL.n97 VTAIL.n83 171.744
R1168 VTAIL.n98 VTAIL.n97 171.744
R1169 VTAIL.n98 VTAIL.n79 171.744
R1170 VTAIL.n105 VTAIL.n79 171.744
R1171 VTAIL.n106 VTAIL.n105 171.744
R1172 VTAIL.n106 VTAIL.n75 171.744
R1173 VTAIL.n113 VTAIL.n75 171.744
R1174 VTAIL.n114 VTAIL.n113 171.744
R1175 VTAIL.n114 VTAIL.n71 171.744
R1176 VTAIL.n121 VTAIL.n71 171.744
R1177 VTAIL.n122 VTAIL.n121 171.744
R1178 VTAIL.n122 VTAIL.n67 171.744
R1179 VTAIL.n129 VTAIL.n67 171.744
R1180 VTAIL.n156 VTAIL.n155 171.744
R1181 VTAIL.n156 VTAIL.n149 171.744
R1182 VTAIL.n163 VTAIL.n149 171.744
R1183 VTAIL.n164 VTAIL.n163 171.744
R1184 VTAIL.n164 VTAIL.n145 171.744
R1185 VTAIL.n171 VTAIL.n145 171.744
R1186 VTAIL.n172 VTAIL.n171 171.744
R1187 VTAIL.n172 VTAIL.n141 171.744
R1188 VTAIL.n179 VTAIL.n141 171.744
R1189 VTAIL.n180 VTAIL.n179 171.744
R1190 VTAIL.n180 VTAIL.n137 171.744
R1191 VTAIL.n187 VTAIL.n137 171.744
R1192 VTAIL.n188 VTAIL.n187 171.744
R1193 VTAIL.n188 VTAIL.n133 171.744
R1194 VTAIL.n195 VTAIL.n133 171.744
R1195 VTAIL.n459 VTAIL.n397 171.744
R1196 VTAIL.n452 VTAIL.n397 171.744
R1197 VTAIL.n452 VTAIL.n451 171.744
R1198 VTAIL.n451 VTAIL.n401 171.744
R1199 VTAIL.n444 VTAIL.n401 171.744
R1200 VTAIL.n444 VTAIL.n443 171.744
R1201 VTAIL.n443 VTAIL.n405 171.744
R1202 VTAIL.n436 VTAIL.n405 171.744
R1203 VTAIL.n436 VTAIL.n435 171.744
R1204 VTAIL.n435 VTAIL.n409 171.744
R1205 VTAIL.n428 VTAIL.n409 171.744
R1206 VTAIL.n428 VTAIL.n427 171.744
R1207 VTAIL.n427 VTAIL.n413 171.744
R1208 VTAIL.n420 VTAIL.n413 171.744
R1209 VTAIL.n420 VTAIL.n419 171.744
R1210 VTAIL.n393 VTAIL.n331 171.744
R1211 VTAIL.n386 VTAIL.n331 171.744
R1212 VTAIL.n386 VTAIL.n385 171.744
R1213 VTAIL.n385 VTAIL.n335 171.744
R1214 VTAIL.n378 VTAIL.n335 171.744
R1215 VTAIL.n378 VTAIL.n377 171.744
R1216 VTAIL.n377 VTAIL.n339 171.744
R1217 VTAIL.n370 VTAIL.n339 171.744
R1218 VTAIL.n370 VTAIL.n369 171.744
R1219 VTAIL.n369 VTAIL.n343 171.744
R1220 VTAIL.n362 VTAIL.n343 171.744
R1221 VTAIL.n362 VTAIL.n361 171.744
R1222 VTAIL.n361 VTAIL.n347 171.744
R1223 VTAIL.n354 VTAIL.n347 171.744
R1224 VTAIL.n354 VTAIL.n353 171.744
R1225 VTAIL.n327 VTAIL.n265 171.744
R1226 VTAIL.n320 VTAIL.n265 171.744
R1227 VTAIL.n320 VTAIL.n319 171.744
R1228 VTAIL.n319 VTAIL.n269 171.744
R1229 VTAIL.n312 VTAIL.n269 171.744
R1230 VTAIL.n312 VTAIL.n311 171.744
R1231 VTAIL.n311 VTAIL.n273 171.744
R1232 VTAIL.n304 VTAIL.n273 171.744
R1233 VTAIL.n304 VTAIL.n303 171.744
R1234 VTAIL.n303 VTAIL.n277 171.744
R1235 VTAIL.n296 VTAIL.n277 171.744
R1236 VTAIL.n296 VTAIL.n295 171.744
R1237 VTAIL.n295 VTAIL.n281 171.744
R1238 VTAIL.n288 VTAIL.n281 171.744
R1239 VTAIL.n288 VTAIL.n287 171.744
R1240 VTAIL.n261 VTAIL.n199 171.744
R1241 VTAIL.n254 VTAIL.n199 171.744
R1242 VTAIL.n254 VTAIL.n253 171.744
R1243 VTAIL.n253 VTAIL.n203 171.744
R1244 VTAIL.n246 VTAIL.n203 171.744
R1245 VTAIL.n246 VTAIL.n245 171.744
R1246 VTAIL.n245 VTAIL.n207 171.744
R1247 VTAIL.n238 VTAIL.n207 171.744
R1248 VTAIL.n238 VTAIL.n237 171.744
R1249 VTAIL.n237 VTAIL.n211 171.744
R1250 VTAIL.n230 VTAIL.n211 171.744
R1251 VTAIL.n230 VTAIL.n229 171.744
R1252 VTAIL.n229 VTAIL.n215 171.744
R1253 VTAIL.n222 VTAIL.n215 171.744
R1254 VTAIL.n222 VTAIL.n221 171.744
R1255 VTAIL.n485 VTAIL.t5 85.8723
R1256 VTAIL.n23 VTAIL.t7 85.8723
R1257 VTAIL.n89 VTAIL.t0 85.8723
R1258 VTAIL.n155 VTAIL.t2 85.8723
R1259 VTAIL.n419 VTAIL.t3 85.8723
R1260 VTAIL.n353 VTAIL.t1 85.8723
R1261 VTAIL.n287 VTAIL.t6 85.8723
R1262 VTAIL.n221 VTAIL.t4 85.8723
R1263 VTAIL.n527 VTAIL.n526 35.0944
R1264 VTAIL.n65 VTAIL.n64 35.0944
R1265 VTAIL.n131 VTAIL.n130 35.0944
R1266 VTAIL.n197 VTAIL.n196 35.0944
R1267 VTAIL.n461 VTAIL.n460 35.0944
R1268 VTAIL.n395 VTAIL.n394 35.0944
R1269 VTAIL.n329 VTAIL.n328 35.0944
R1270 VTAIL.n263 VTAIL.n262 35.0944
R1271 VTAIL.n527 VTAIL.n461 25.1169
R1272 VTAIL.n263 VTAIL.n197 25.1169
R1273 VTAIL.n484 VTAIL.n483 16.3895
R1274 VTAIL.n22 VTAIL.n21 16.3895
R1275 VTAIL.n88 VTAIL.n87 16.3895
R1276 VTAIL.n154 VTAIL.n153 16.3895
R1277 VTAIL.n418 VTAIL.n417 16.3895
R1278 VTAIL.n352 VTAIL.n351 16.3895
R1279 VTAIL.n286 VTAIL.n285 16.3895
R1280 VTAIL.n220 VTAIL.n219 16.3895
R1281 VTAIL.n487 VTAIL.n482 12.8005
R1282 VTAIL.n25 VTAIL.n20 12.8005
R1283 VTAIL.n91 VTAIL.n86 12.8005
R1284 VTAIL.n157 VTAIL.n152 12.8005
R1285 VTAIL.n421 VTAIL.n416 12.8005
R1286 VTAIL.n355 VTAIL.n350 12.8005
R1287 VTAIL.n289 VTAIL.n284 12.8005
R1288 VTAIL.n223 VTAIL.n218 12.8005
R1289 VTAIL.n488 VTAIL.n480 12.0247
R1290 VTAIL.n524 VTAIL.n462 12.0247
R1291 VTAIL.n26 VTAIL.n18 12.0247
R1292 VTAIL.n62 VTAIL.n0 12.0247
R1293 VTAIL.n92 VTAIL.n84 12.0247
R1294 VTAIL.n128 VTAIL.n66 12.0247
R1295 VTAIL.n158 VTAIL.n150 12.0247
R1296 VTAIL.n194 VTAIL.n132 12.0247
R1297 VTAIL.n458 VTAIL.n396 12.0247
R1298 VTAIL.n422 VTAIL.n414 12.0247
R1299 VTAIL.n392 VTAIL.n330 12.0247
R1300 VTAIL.n356 VTAIL.n348 12.0247
R1301 VTAIL.n326 VTAIL.n264 12.0247
R1302 VTAIL.n290 VTAIL.n282 12.0247
R1303 VTAIL.n260 VTAIL.n198 12.0247
R1304 VTAIL.n224 VTAIL.n216 12.0247
R1305 VTAIL.n492 VTAIL.n491 11.249
R1306 VTAIL.n523 VTAIL.n464 11.249
R1307 VTAIL.n30 VTAIL.n29 11.249
R1308 VTAIL.n61 VTAIL.n2 11.249
R1309 VTAIL.n96 VTAIL.n95 11.249
R1310 VTAIL.n127 VTAIL.n68 11.249
R1311 VTAIL.n162 VTAIL.n161 11.249
R1312 VTAIL.n193 VTAIL.n134 11.249
R1313 VTAIL.n457 VTAIL.n398 11.249
R1314 VTAIL.n426 VTAIL.n425 11.249
R1315 VTAIL.n391 VTAIL.n332 11.249
R1316 VTAIL.n360 VTAIL.n359 11.249
R1317 VTAIL.n325 VTAIL.n266 11.249
R1318 VTAIL.n294 VTAIL.n293 11.249
R1319 VTAIL.n259 VTAIL.n200 11.249
R1320 VTAIL.n228 VTAIL.n227 11.249
R1321 VTAIL.n495 VTAIL.n478 10.4732
R1322 VTAIL.n520 VTAIL.n519 10.4732
R1323 VTAIL.n33 VTAIL.n16 10.4732
R1324 VTAIL.n58 VTAIL.n57 10.4732
R1325 VTAIL.n99 VTAIL.n82 10.4732
R1326 VTAIL.n124 VTAIL.n123 10.4732
R1327 VTAIL.n165 VTAIL.n148 10.4732
R1328 VTAIL.n190 VTAIL.n189 10.4732
R1329 VTAIL.n454 VTAIL.n453 10.4732
R1330 VTAIL.n429 VTAIL.n412 10.4732
R1331 VTAIL.n388 VTAIL.n387 10.4732
R1332 VTAIL.n363 VTAIL.n346 10.4732
R1333 VTAIL.n322 VTAIL.n321 10.4732
R1334 VTAIL.n297 VTAIL.n280 10.4732
R1335 VTAIL.n256 VTAIL.n255 10.4732
R1336 VTAIL.n231 VTAIL.n214 10.4732
R1337 VTAIL.n496 VTAIL.n476 9.69747
R1338 VTAIL.n516 VTAIL.n466 9.69747
R1339 VTAIL.n34 VTAIL.n14 9.69747
R1340 VTAIL.n54 VTAIL.n4 9.69747
R1341 VTAIL.n100 VTAIL.n80 9.69747
R1342 VTAIL.n120 VTAIL.n70 9.69747
R1343 VTAIL.n166 VTAIL.n146 9.69747
R1344 VTAIL.n186 VTAIL.n136 9.69747
R1345 VTAIL.n450 VTAIL.n400 9.69747
R1346 VTAIL.n430 VTAIL.n410 9.69747
R1347 VTAIL.n384 VTAIL.n334 9.69747
R1348 VTAIL.n364 VTAIL.n344 9.69747
R1349 VTAIL.n318 VTAIL.n268 9.69747
R1350 VTAIL.n298 VTAIL.n278 9.69747
R1351 VTAIL.n252 VTAIL.n202 9.69747
R1352 VTAIL.n232 VTAIL.n212 9.69747
R1353 VTAIL.n522 VTAIL.n462 9.45567
R1354 VTAIL.n60 VTAIL.n0 9.45567
R1355 VTAIL.n126 VTAIL.n66 9.45567
R1356 VTAIL.n192 VTAIL.n132 9.45567
R1357 VTAIL.n456 VTAIL.n396 9.45567
R1358 VTAIL.n390 VTAIL.n330 9.45567
R1359 VTAIL.n324 VTAIL.n264 9.45567
R1360 VTAIL.n258 VTAIL.n198 9.45567
R1361 VTAIL.n507 VTAIL.n506 9.3005
R1362 VTAIL.n470 VTAIL.n469 9.3005
R1363 VTAIL.n513 VTAIL.n512 9.3005
R1364 VTAIL.n515 VTAIL.n514 9.3005
R1365 VTAIL.n466 VTAIL.n465 9.3005
R1366 VTAIL.n521 VTAIL.n520 9.3005
R1367 VTAIL.n523 VTAIL.n522 9.3005
R1368 VTAIL.n474 VTAIL.n473 9.3005
R1369 VTAIL.n499 VTAIL.n498 9.3005
R1370 VTAIL.n497 VTAIL.n496 9.3005
R1371 VTAIL.n478 VTAIL.n477 9.3005
R1372 VTAIL.n491 VTAIL.n490 9.3005
R1373 VTAIL.n489 VTAIL.n488 9.3005
R1374 VTAIL.n482 VTAIL.n481 9.3005
R1375 VTAIL.n505 VTAIL.n504 9.3005
R1376 VTAIL.n45 VTAIL.n44 9.3005
R1377 VTAIL.n8 VTAIL.n7 9.3005
R1378 VTAIL.n51 VTAIL.n50 9.3005
R1379 VTAIL.n53 VTAIL.n52 9.3005
R1380 VTAIL.n4 VTAIL.n3 9.3005
R1381 VTAIL.n59 VTAIL.n58 9.3005
R1382 VTAIL.n61 VTAIL.n60 9.3005
R1383 VTAIL.n12 VTAIL.n11 9.3005
R1384 VTAIL.n37 VTAIL.n36 9.3005
R1385 VTAIL.n35 VTAIL.n34 9.3005
R1386 VTAIL.n16 VTAIL.n15 9.3005
R1387 VTAIL.n29 VTAIL.n28 9.3005
R1388 VTAIL.n27 VTAIL.n26 9.3005
R1389 VTAIL.n20 VTAIL.n19 9.3005
R1390 VTAIL.n43 VTAIL.n42 9.3005
R1391 VTAIL.n111 VTAIL.n110 9.3005
R1392 VTAIL.n74 VTAIL.n73 9.3005
R1393 VTAIL.n117 VTAIL.n116 9.3005
R1394 VTAIL.n119 VTAIL.n118 9.3005
R1395 VTAIL.n70 VTAIL.n69 9.3005
R1396 VTAIL.n125 VTAIL.n124 9.3005
R1397 VTAIL.n127 VTAIL.n126 9.3005
R1398 VTAIL.n78 VTAIL.n77 9.3005
R1399 VTAIL.n103 VTAIL.n102 9.3005
R1400 VTAIL.n101 VTAIL.n100 9.3005
R1401 VTAIL.n82 VTAIL.n81 9.3005
R1402 VTAIL.n95 VTAIL.n94 9.3005
R1403 VTAIL.n93 VTAIL.n92 9.3005
R1404 VTAIL.n86 VTAIL.n85 9.3005
R1405 VTAIL.n109 VTAIL.n108 9.3005
R1406 VTAIL.n177 VTAIL.n176 9.3005
R1407 VTAIL.n140 VTAIL.n139 9.3005
R1408 VTAIL.n183 VTAIL.n182 9.3005
R1409 VTAIL.n185 VTAIL.n184 9.3005
R1410 VTAIL.n136 VTAIL.n135 9.3005
R1411 VTAIL.n191 VTAIL.n190 9.3005
R1412 VTAIL.n193 VTAIL.n192 9.3005
R1413 VTAIL.n144 VTAIL.n143 9.3005
R1414 VTAIL.n169 VTAIL.n168 9.3005
R1415 VTAIL.n167 VTAIL.n166 9.3005
R1416 VTAIL.n148 VTAIL.n147 9.3005
R1417 VTAIL.n161 VTAIL.n160 9.3005
R1418 VTAIL.n159 VTAIL.n158 9.3005
R1419 VTAIL.n152 VTAIL.n151 9.3005
R1420 VTAIL.n175 VTAIL.n174 9.3005
R1421 VTAIL.n457 VTAIL.n456 9.3005
R1422 VTAIL.n455 VTAIL.n454 9.3005
R1423 VTAIL.n400 VTAIL.n399 9.3005
R1424 VTAIL.n449 VTAIL.n448 9.3005
R1425 VTAIL.n447 VTAIL.n446 9.3005
R1426 VTAIL.n404 VTAIL.n403 9.3005
R1427 VTAIL.n441 VTAIL.n440 9.3005
R1428 VTAIL.n439 VTAIL.n438 9.3005
R1429 VTAIL.n408 VTAIL.n407 9.3005
R1430 VTAIL.n433 VTAIL.n432 9.3005
R1431 VTAIL.n431 VTAIL.n430 9.3005
R1432 VTAIL.n412 VTAIL.n411 9.3005
R1433 VTAIL.n425 VTAIL.n424 9.3005
R1434 VTAIL.n423 VTAIL.n422 9.3005
R1435 VTAIL.n416 VTAIL.n415 9.3005
R1436 VTAIL.n338 VTAIL.n337 9.3005
R1437 VTAIL.n381 VTAIL.n380 9.3005
R1438 VTAIL.n383 VTAIL.n382 9.3005
R1439 VTAIL.n334 VTAIL.n333 9.3005
R1440 VTAIL.n389 VTAIL.n388 9.3005
R1441 VTAIL.n391 VTAIL.n390 9.3005
R1442 VTAIL.n375 VTAIL.n374 9.3005
R1443 VTAIL.n373 VTAIL.n372 9.3005
R1444 VTAIL.n342 VTAIL.n341 9.3005
R1445 VTAIL.n367 VTAIL.n366 9.3005
R1446 VTAIL.n365 VTAIL.n364 9.3005
R1447 VTAIL.n346 VTAIL.n345 9.3005
R1448 VTAIL.n359 VTAIL.n358 9.3005
R1449 VTAIL.n357 VTAIL.n356 9.3005
R1450 VTAIL.n350 VTAIL.n349 9.3005
R1451 VTAIL.n272 VTAIL.n271 9.3005
R1452 VTAIL.n315 VTAIL.n314 9.3005
R1453 VTAIL.n317 VTAIL.n316 9.3005
R1454 VTAIL.n268 VTAIL.n267 9.3005
R1455 VTAIL.n323 VTAIL.n322 9.3005
R1456 VTAIL.n325 VTAIL.n324 9.3005
R1457 VTAIL.n309 VTAIL.n308 9.3005
R1458 VTAIL.n307 VTAIL.n306 9.3005
R1459 VTAIL.n276 VTAIL.n275 9.3005
R1460 VTAIL.n301 VTAIL.n300 9.3005
R1461 VTAIL.n299 VTAIL.n298 9.3005
R1462 VTAIL.n280 VTAIL.n279 9.3005
R1463 VTAIL.n293 VTAIL.n292 9.3005
R1464 VTAIL.n291 VTAIL.n290 9.3005
R1465 VTAIL.n284 VTAIL.n283 9.3005
R1466 VTAIL.n206 VTAIL.n205 9.3005
R1467 VTAIL.n249 VTAIL.n248 9.3005
R1468 VTAIL.n251 VTAIL.n250 9.3005
R1469 VTAIL.n202 VTAIL.n201 9.3005
R1470 VTAIL.n257 VTAIL.n256 9.3005
R1471 VTAIL.n259 VTAIL.n258 9.3005
R1472 VTAIL.n243 VTAIL.n242 9.3005
R1473 VTAIL.n241 VTAIL.n240 9.3005
R1474 VTAIL.n210 VTAIL.n209 9.3005
R1475 VTAIL.n235 VTAIL.n234 9.3005
R1476 VTAIL.n233 VTAIL.n232 9.3005
R1477 VTAIL.n214 VTAIL.n213 9.3005
R1478 VTAIL.n227 VTAIL.n226 9.3005
R1479 VTAIL.n225 VTAIL.n224 9.3005
R1480 VTAIL.n218 VTAIL.n217 9.3005
R1481 VTAIL.n500 VTAIL.n499 8.92171
R1482 VTAIL.n515 VTAIL.n468 8.92171
R1483 VTAIL.n38 VTAIL.n37 8.92171
R1484 VTAIL.n53 VTAIL.n6 8.92171
R1485 VTAIL.n104 VTAIL.n103 8.92171
R1486 VTAIL.n119 VTAIL.n72 8.92171
R1487 VTAIL.n170 VTAIL.n169 8.92171
R1488 VTAIL.n185 VTAIL.n138 8.92171
R1489 VTAIL.n449 VTAIL.n402 8.92171
R1490 VTAIL.n434 VTAIL.n433 8.92171
R1491 VTAIL.n383 VTAIL.n336 8.92171
R1492 VTAIL.n368 VTAIL.n367 8.92171
R1493 VTAIL.n317 VTAIL.n270 8.92171
R1494 VTAIL.n302 VTAIL.n301 8.92171
R1495 VTAIL.n251 VTAIL.n204 8.92171
R1496 VTAIL.n236 VTAIL.n235 8.92171
R1497 VTAIL.n503 VTAIL.n474 8.14595
R1498 VTAIL.n512 VTAIL.n511 8.14595
R1499 VTAIL.n41 VTAIL.n12 8.14595
R1500 VTAIL.n50 VTAIL.n49 8.14595
R1501 VTAIL.n107 VTAIL.n78 8.14595
R1502 VTAIL.n116 VTAIL.n115 8.14595
R1503 VTAIL.n173 VTAIL.n144 8.14595
R1504 VTAIL.n182 VTAIL.n181 8.14595
R1505 VTAIL.n446 VTAIL.n445 8.14595
R1506 VTAIL.n437 VTAIL.n408 8.14595
R1507 VTAIL.n380 VTAIL.n379 8.14595
R1508 VTAIL.n371 VTAIL.n342 8.14595
R1509 VTAIL.n314 VTAIL.n313 8.14595
R1510 VTAIL.n305 VTAIL.n276 8.14595
R1511 VTAIL.n248 VTAIL.n247 8.14595
R1512 VTAIL.n239 VTAIL.n210 8.14595
R1513 VTAIL.n504 VTAIL.n472 7.3702
R1514 VTAIL.n508 VTAIL.n470 7.3702
R1515 VTAIL.n42 VTAIL.n10 7.3702
R1516 VTAIL.n46 VTAIL.n8 7.3702
R1517 VTAIL.n108 VTAIL.n76 7.3702
R1518 VTAIL.n112 VTAIL.n74 7.3702
R1519 VTAIL.n174 VTAIL.n142 7.3702
R1520 VTAIL.n178 VTAIL.n140 7.3702
R1521 VTAIL.n442 VTAIL.n404 7.3702
R1522 VTAIL.n438 VTAIL.n406 7.3702
R1523 VTAIL.n376 VTAIL.n338 7.3702
R1524 VTAIL.n372 VTAIL.n340 7.3702
R1525 VTAIL.n310 VTAIL.n272 7.3702
R1526 VTAIL.n306 VTAIL.n274 7.3702
R1527 VTAIL.n244 VTAIL.n206 7.3702
R1528 VTAIL.n240 VTAIL.n208 7.3702
R1529 VTAIL.n507 VTAIL.n472 6.59444
R1530 VTAIL.n508 VTAIL.n507 6.59444
R1531 VTAIL.n45 VTAIL.n10 6.59444
R1532 VTAIL.n46 VTAIL.n45 6.59444
R1533 VTAIL.n111 VTAIL.n76 6.59444
R1534 VTAIL.n112 VTAIL.n111 6.59444
R1535 VTAIL.n177 VTAIL.n142 6.59444
R1536 VTAIL.n178 VTAIL.n177 6.59444
R1537 VTAIL.n442 VTAIL.n441 6.59444
R1538 VTAIL.n441 VTAIL.n406 6.59444
R1539 VTAIL.n376 VTAIL.n375 6.59444
R1540 VTAIL.n375 VTAIL.n340 6.59444
R1541 VTAIL.n310 VTAIL.n309 6.59444
R1542 VTAIL.n309 VTAIL.n274 6.59444
R1543 VTAIL.n244 VTAIL.n243 6.59444
R1544 VTAIL.n243 VTAIL.n208 6.59444
R1545 VTAIL.n504 VTAIL.n503 5.81868
R1546 VTAIL.n511 VTAIL.n470 5.81868
R1547 VTAIL.n42 VTAIL.n41 5.81868
R1548 VTAIL.n49 VTAIL.n8 5.81868
R1549 VTAIL.n108 VTAIL.n107 5.81868
R1550 VTAIL.n115 VTAIL.n74 5.81868
R1551 VTAIL.n174 VTAIL.n173 5.81868
R1552 VTAIL.n181 VTAIL.n140 5.81868
R1553 VTAIL.n445 VTAIL.n404 5.81868
R1554 VTAIL.n438 VTAIL.n437 5.81868
R1555 VTAIL.n379 VTAIL.n338 5.81868
R1556 VTAIL.n372 VTAIL.n371 5.81868
R1557 VTAIL.n313 VTAIL.n272 5.81868
R1558 VTAIL.n306 VTAIL.n305 5.81868
R1559 VTAIL.n247 VTAIL.n206 5.81868
R1560 VTAIL.n240 VTAIL.n239 5.81868
R1561 VTAIL.n500 VTAIL.n474 5.04292
R1562 VTAIL.n512 VTAIL.n468 5.04292
R1563 VTAIL.n38 VTAIL.n12 5.04292
R1564 VTAIL.n50 VTAIL.n6 5.04292
R1565 VTAIL.n104 VTAIL.n78 5.04292
R1566 VTAIL.n116 VTAIL.n72 5.04292
R1567 VTAIL.n170 VTAIL.n144 5.04292
R1568 VTAIL.n182 VTAIL.n138 5.04292
R1569 VTAIL.n446 VTAIL.n402 5.04292
R1570 VTAIL.n434 VTAIL.n408 5.04292
R1571 VTAIL.n380 VTAIL.n336 5.04292
R1572 VTAIL.n368 VTAIL.n342 5.04292
R1573 VTAIL.n314 VTAIL.n270 5.04292
R1574 VTAIL.n302 VTAIL.n276 5.04292
R1575 VTAIL.n248 VTAIL.n204 5.04292
R1576 VTAIL.n236 VTAIL.n210 5.04292
R1577 VTAIL.n499 VTAIL.n476 4.26717
R1578 VTAIL.n516 VTAIL.n515 4.26717
R1579 VTAIL.n37 VTAIL.n14 4.26717
R1580 VTAIL.n54 VTAIL.n53 4.26717
R1581 VTAIL.n103 VTAIL.n80 4.26717
R1582 VTAIL.n120 VTAIL.n119 4.26717
R1583 VTAIL.n169 VTAIL.n146 4.26717
R1584 VTAIL.n186 VTAIL.n185 4.26717
R1585 VTAIL.n450 VTAIL.n449 4.26717
R1586 VTAIL.n433 VTAIL.n410 4.26717
R1587 VTAIL.n384 VTAIL.n383 4.26717
R1588 VTAIL.n367 VTAIL.n344 4.26717
R1589 VTAIL.n318 VTAIL.n317 4.26717
R1590 VTAIL.n301 VTAIL.n278 4.26717
R1591 VTAIL.n252 VTAIL.n251 4.26717
R1592 VTAIL.n235 VTAIL.n212 4.26717
R1593 VTAIL.n417 VTAIL.n415 3.70982
R1594 VTAIL.n351 VTAIL.n349 3.70982
R1595 VTAIL.n285 VTAIL.n283 3.70982
R1596 VTAIL.n219 VTAIL.n217 3.70982
R1597 VTAIL.n483 VTAIL.n481 3.70982
R1598 VTAIL.n21 VTAIL.n19 3.70982
R1599 VTAIL.n87 VTAIL.n85 3.70982
R1600 VTAIL.n153 VTAIL.n151 3.70982
R1601 VTAIL.n496 VTAIL.n495 3.49141
R1602 VTAIL.n519 VTAIL.n466 3.49141
R1603 VTAIL.n34 VTAIL.n33 3.49141
R1604 VTAIL.n57 VTAIL.n4 3.49141
R1605 VTAIL.n100 VTAIL.n99 3.49141
R1606 VTAIL.n123 VTAIL.n70 3.49141
R1607 VTAIL.n166 VTAIL.n165 3.49141
R1608 VTAIL.n189 VTAIL.n136 3.49141
R1609 VTAIL.n453 VTAIL.n400 3.49141
R1610 VTAIL.n430 VTAIL.n429 3.49141
R1611 VTAIL.n387 VTAIL.n334 3.49141
R1612 VTAIL.n364 VTAIL.n363 3.49141
R1613 VTAIL.n321 VTAIL.n268 3.49141
R1614 VTAIL.n298 VTAIL.n297 3.49141
R1615 VTAIL.n255 VTAIL.n202 3.49141
R1616 VTAIL.n232 VTAIL.n231 3.49141
R1617 VTAIL.n492 VTAIL.n478 2.71565
R1618 VTAIL.n520 VTAIL.n464 2.71565
R1619 VTAIL.n30 VTAIL.n16 2.71565
R1620 VTAIL.n58 VTAIL.n2 2.71565
R1621 VTAIL.n96 VTAIL.n82 2.71565
R1622 VTAIL.n124 VTAIL.n68 2.71565
R1623 VTAIL.n162 VTAIL.n148 2.71565
R1624 VTAIL.n190 VTAIL.n134 2.71565
R1625 VTAIL.n454 VTAIL.n398 2.71565
R1626 VTAIL.n426 VTAIL.n412 2.71565
R1627 VTAIL.n388 VTAIL.n332 2.71565
R1628 VTAIL.n360 VTAIL.n346 2.71565
R1629 VTAIL.n322 VTAIL.n266 2.71565
R1630 VTAIL.n294 VTAIL.n280 2.71565
R1631 VTAIL.n256 VTAIL.n200 2.71565
R1632 VTAIL.n228 VTAIL.n214 2.71565
R1633 VTAIL.n329 VTAIL.n263 2.43153
R1634 VTAIL.n461 VTAIL.n395 2.43153
R1635 VTAIL.n197 VTAIL.n131 2.43153
R1636 VTAIL.n491 VTAIL.n480 1.93989
R1637 VTAIL.n524 VTAIL.n523 1.93989
R1638 VTAIL.n29 VTAIL.n18 1.93989
R1639 VTAIL.n62 VTAIL.n61 1.93989
R1640 VTAIL.n95 VTAIL.n84 1.93989
R1641 VTAIL.n128 VTAIL.n127 1.93989
R1642 VTAIL.n161 VTAIL.n150 1.93989
R1643 VTAIL.n194 VTAIL.n193 1.93989
R1644 VTAIL.n458 VTAIL.n457 1.93989
R1645 VTAIL.n425 VTAIL.n414 1.93989
R1646 VTAIL.n392 VTAIL.n391 1.93989
R1647 VTAIL.n359 VTAIL.n348 1.93989
R1648 VTAIL.n326 VTAIL.n325 1.93989
R1649 VTAIL.n293 VTAIL.n282 1.93989
R1650 VTAIL.n260 VTAIL.n259 1.93989
R1651 VTAIL.n227 VTAIL.n216 1.93989
R1652 VTAIL VTAIL.n65 1.27421
R1653 VTAIL.n488 VTAIL.n487 1.16414
R1654 VTAIL.n526 VTAIL.n462 1.16414
R1655 VTAIL.n26 VTAIL.n25 1.16414
R1656 VTAIL.n64 VTAIL.n0 1.16414
R1657 VTAIL.n92 VTAIL.n91 1.16414
R1658 VTAIL.n130 VTAIL.n66 1.16414
R1659 VTAIL.n158 VTAIL.n157 1.16414
R1660 VTAIL.n196 VTAIL.n132 1.16414
R1661 VTAIL.n460 VTAIL.n396 1.16414
R1662 VTAIL.n422 VTAIL.n421 1.16414
R1663 VTAIL.n394 VTAIL.n330 1.16414
R1664 VTAIL.n356 VTAIL.n355 1.16414
R1665 VTAIL.n328 VTAIL.n264 1.16414
R1666 VTAIL.n290 VTAIL.n289 1.16414
R1667 VTAIL.n262 VTAIL.n198 1.16414
R1668 VTAIL.n224 VTAIL.n223 1.16414
R1669 VTAIL VTAIL.n527 1.15783
R1670 VTAIL.n395 VTAIL.n329 0.470328
R1671 VTAIL.n131 VTAIL.n65 0.470328
R1672 VTAIL.n484 VTAIL.n482 0.388379
R1673 VTAIL.n22 VTAIL.n20 0.388379
R1674 VTAIL.n88 VTAIL.n86 0.388379
R1675 VTAIL.n154 VTAIL.n152 0.388379
R1676 VTAIL.n418 VTAIL.n416 0.388379
R1677 VTAIL.n352 VTAIL.n350 0.388379
R1678 VTAIL.n286 VTAIL.n284 0.388379
R1679 VTAIL.n220 VTAIL.n218 0.388379
R1680 VTAIL.n489 VTAIL.n481 0.155672
R1681 VTAIL.n490 VTAIL.n489 0.155672
R1682 VTAIL.n490 VTAIL.n477 0.155672
R1683 VTAIL.n497 VTAIL.n477 0.155672
R1684 VTAIL.n498 VTAIL.n497 0.155672
R1685 VTAIL.n498 VTAIL.n473 0.155672
R1686 VTAIL.n505 VTAIL.n473 0.155672
R1687 VTAIL.n506 VTAIL.n505 0.155672
R1688 VTAIL.n506 VTAIL.n469 0.155672
R1689 VTAIL.n513 VTAIL.n469 0.155672
R1690 VTAIL.n514 VTAIL.n513 0.155672
R1691 VTAIL.n514 VTAIL.n465 0.155672
R1692 VTAIL.n521 VTAIL.n465 0.155672
R1693 VTAIL.n522 VTAIL.n521 0.155672
R1694 VTAIL.n27 VTAIL.n19 0.155672
R1695 VTAIL.n28 VTAIL.n27 0.155672
R1696 VTAIL.n28 VTAIL.n15 0.155672
R1697 VTAIL.n35 VTAIL.n15 0.155672
R1698 VTAIL.n36 VTAIL.n35 0.155672
R1699 VTAIL.n36 VTAIL.n11 0.155672
R1700 VTAIL.n43 VTAIL.n11 0.155672
R1701 VTAIL.n44 VTAIL.n43 0.155672
R1702 VTAIL.n44 VTAIL.n7 0.155672
R1703 VTAIL.n51 VTAIL.n7 0.155672
R1704 VTAIL.n52 VTAIL.n51 0.155672
R1705 VTAIL.n52 VTAIL.n3 0.155672
R1706 VTAIL.n59 VTAIL.n3 0.155672
R1707 VTAIL.n60 VTAIL.n59 0.155672
R1708 VTAIL.n93 VTAIL.n85 0.155672
R1709 VTAIL.n94 VTAIL.n93 0.155672
R1710 VTAIL.n94 VTAIL.n81 0.155672
R1711 VTAIL.n101 VTAIL.n81 0.155672
R1712 VTAIL.n102 VTAIL.n101 0.155672
R1713 VTAIL.n102 VTAIL.n77 0.155672
R1714 VTAIL.n109 VTAIL.n77 0.155672
R1715 VTAIL.n110 VTAIL.n109 0.155672
R1716 VTAIL.n110 VTAIL.n73 0.155672
R1717 VTAIL.n117 VTAIL.n73 0.155672
R1718 VTAIL.n118 VTAIL.n117 0.155672
R1719 VTAIL.n118 VTAIL.n69 0.155672
R1720 VTAIL.n125 VTAIL.n69 0.155672
R1721 VTAIL.n126 VTAIL.n125 0.155672
R1722 VTAIL.n159 VTAIL.n151 0.155672
R1723 VTAIL.n160 VTAIL.n159 0.155672
R1724 VTAIL.n160 VTAIL.n147 0.155672
R1725 VTAIL.n167 VTAIL.n147 0.155672
R1726 VTAIL.n168 VTAIL.n167 0.155672
R1727 VTAIL.n168 VTAIL.n143 0.155672
R1728 VTAIL.n175 VTAIL.n143 0.155672
R1729 VTAIL.n176 VTAIL.n175 0.155672
R1730 VTAIL.n176 VTAIL.n139 0.155672
R1731 VTAIL.n183 VTAIL.n139 0.155672
R1732 VTAIL.n184 VTAIL.n183 0.155672
R1733 VTAIL.n184 VTAIL.n135 0.155672
R1734 VTAIL.n191 VTAIL.n135 0.155672
R1735 VTAIL.n192 VTAIL.n191 0.155672
R1736 VTAIL.n456 VTAIL.n455 0.155672
R1737 VTAIL.n455 VTAIL.n399 0.155672
R1738 VTAIL.n448 VTAIL.n399 0.155672
R1739 VTAIL.n448 VTAIL.n447 0.155672
R1740 VTAIL.n447 VTAIL.n403 0.155672
R1741 VTAIL.n440 VTAIL.n403 0.155672
R1742 VTAIL.n440 VTAIL.n439 0.155672
R1743 VTAIL.n439 VTAIL.n407 0.155672
R1744 VTAIL.n432 VTAIL.n407 0.155672
R1745 VTAIL.n432 VTAIL.n431 0.155672
R1746 VTAIL.n431 VTAIL.n411 0.155672
R1747 VTAIL.n424 VTAIL.n411 0.155672
R1748 VTAIL.n424 VTAIL.n423 0.155672
R1749 VTAIL.n423 VTAIL.n415 0.155672
R1750 VTAIL.n390 VTAIL.n389 0.155672
R1751 VTAIL.n389 VTAIL.n333 0.155672
R1752 VTAIL.n382 VTAIL.n333 0.155672
R1753 VTAIL.n382 VTAIL.n381 0.155672
R1754 VTAIL.n381 VTAIL.n337 0.155672
R1755 VTAIL.n374 VTAIL.n337 0.155672
R1756 VTAIL.n374 VTAIL.n373 0.155672
R1757 VTAIL.n373 VTAIL.n341 0.155672
R1758 VTAIL.n366 VTAIL.n341 0.155672
R1759 VTAIL.n366 VTAIL.n365 0.155672
R1760 VTAIL.n365 VTAIL.n345 0.155672
R1761 VTAIL.n358 VTAIL.n345 0.155672
R1762 VTAIL.n358 VTAIL.n357 0.155672
R1763 VTAIL.n357 VTAIL.n349 0.155672
R1764 VTAIL.n324 VTAIL.n323 0.155672
R1765 VTAIL.n323 VTAIL.n267 0.155672
R1766 VTAIL.n316 VTAIL.n267 0.155672
R1767 VTAIL.n316 VTAIL.n315 0.155672
R1768 VTAIL.n315 VTAIL.n271 0.155672
R1769 VTAIL.n308 VTAIL.n271 0.155672
R1770 VTAIL.n308 VTAIL.n307 0.155672
R1771 VTAIL.n307 VTAIL.n275 0.155672
R1772 VTAIL.n300 VTAIL.n275 0.155672
R1773 VTAIL.n300 VTAIL.n299 0.155672
R1774 VTAIL.n299 VTAIL.n279 0.155672
R1775 VTAIL.n292 VTAIL.n279 0.155672
R1776 VTAIL.n292 VTAIL.n291 0.155672
R1777 VTAIL.n291 VTAIL.n283 0.155672
R1778 VTAIL.n258 VTAIL.n257 0.155672
R1779 VTAIL.n257 VTAIL.n201 0.155672
R1780 VTAIL.n250 VTAIL.n201 0.155672
R1781 VTAIL.n250 VTAIL.n249 0.155672
R1782 VTAIL.n249 VTAIL.n205 0.155672
R1783 VTAIL.n242 VTAIL.n205 0.155672
R1784 VTAIL.n242 VTAIL.n241 0.155672
R1785 VTAIL.n241 VTAIL.n209 0.155672
R1786 VTAIL.n234 VTAIL.n209 0.155672
R1787 VTAIL.n234 VTAIL.n233 0.155672
R1788 VTAIL.n233 VTAIL.n213 0.155672
R1789 VTAIL.n226 VTAIL.n213 0.155672
R1790 VTAIL.n226 VTAIL.n225 0.155672
R1791 VTAIL.n225 VTAIL.n217 0.155672
R1792 VDD2.n2 VDD2.n0 118.816
R1793 VDD2.n2 VDD2.n1 77.4875
R1794 VDD2.n1 VDD2.t1 2.71604
R1795 VDD2.n1 VDD2.t0 2.71604
R1796 VDD2.n0 VDD2.t2 2.71604
R1797 VDD2.n0 VDD2.t3 2.71604
R1798 VDD2 VDD2.n2 0.0586897
R1799 VP.n14 VP.n0 161.3
R1800 VP.n13 VP.n12 161.3
R1801 VP.n11 VP.n1 161.3
R1802 VP.n10 VP.n9 161.3
R1803 VP.n8 VP.n2 161.3
R1804 VP.n7 VP.n6 161.3
R1805 VP.n4 VP.t1 151.201
R1806 VP.n4 VP.t0 150.445
R1807 VP.n3 VP.t3 115.855
R1808 VP.n15 VP.t2 115.855
R1809 VP.n5 VP.n3 102.927
R1810 VP.n16 VP.n15 102.927
R1811 VP.n9 VP.n1 56.5193
R1812 VP.n5 VP.n4 50.4405
R1813 VP.n8 VP.n7 24.4675
R1814 VP.n9 VP.n8 24.4675
R1815 VP.n13 VP.n1 24.4675
R1816 VP.n14 VP.n13 24.4675
R1817 VP.n7 VP.n3 7.82994
R1818 VP.n15 VP.n14 7.82994
R1819 VP.n6 VP.n5 0.278367
R1820 VP.n16 VP.n0 0.278367
R1821 VP.n6 VP.n2 0.189894
R1822 VP.n10 VP.n2 0.189894
R1823 VP.n11 VP.n10 0.189894
R1824 VP.n12 VP.n11 0.189894
R1825 VP.n12 VP.n0 0.189894
R1826 VP VP.n16 0.153454
R1827 VDD1 VDD1.n1 119.341
R1828 VDD1 VDD1.n0 77.5457
R1829 VDD1.n0 VDD1.t2 2.71604
R1830 VDD1.n0 VDD1.t3 2.71604
R1831 VDD1.n1 VDD1.t0 2.71604
R1832 VDD1.n1 VDD1.t1 2.71604
C0 VTAIL B 4.88672f
C1 VP B 1.65434f
C2 VN w_n2662_n3362# 4.49048f
C3 VDD1 B 1.24038f
C4 VDD2 w_n2662_n3362# 1.48778f
C5 VTAIL w_n2662_n3362# 3.96688f
C6 VP w_n2662_n3362# 4.83241f
C7 VDD1 w_n2662_n3362# 1.43407f
C8 VN VDD2 4.69841f
C9 VTAIL VN 4.5967f
C10 VN VP 6.10803f
C11 VN VDD1 0.149034f
C12 w_n2662_n3362# B 9.10279f
C13 VTAIL VDD2 5.43803f
C14 VDD2 VP 0.387439f
C15 VDD2 VDD1 1.00702f
C16 VN B 1.08743f
C17 VTAIL VP 4.61081f
C18 VTAIL VDD1 5.38456f
C19 VDD1 VP 4.93611f
C20 VDD2 B 1.29069f
C21 VDD2 VSUBS 0.917933f
C22 VDD1 VSUBS 5.62896f
C23 VTAIL VSUBS 1.198391f
C24 VN VSUBS 5.39798f
C25 VP VSUBS 2.223042f
C26 B VSUBS 4.180214f
C27 w_n2662_n3362# VSUBS 0.110175p
C28 VDD1.t2 VSUBS 0.25508f
C29 VDD1.t3 VSUBS 0.25508f
C30 VDD1.n0 VSUBS 2.01563f
C31 VDD1.t0 VSUBS 0.25508f
C32 VDD1.t1 VSUBS 0.25508f
C33 VDD1.n1 VSUBS 2.71094f
C34 VP.n0 VSUBS 0.045708f
C35 VP.t2 VSUBS 2.81522f
C36 VP.n1 VSUBS 0.050611f
C37 VP.n2 VSUBS 0.034669f
C38 VP.t3 VSUBS 2.81522f
C39 VP.n3 VSUBS 1.10423f
C40 VP.t0 VSUBS 3.09289f
C41 VP.t1 VSUBS 3.09887f
C42 VP.n4 VSUBS 3.81974f
C43 VP.n5 VSUBS 1.90653f
C44 VP.n6 VSUBS 0.045708f
C45 VP.n7 VSUBS 0.042922f
C46 VP.n8 VSUBS 0.064615f
C47 VP.n9 VSUBS 0.050611f
C48 VP.n10 VSUBS 0.034669f
C49 VP.n11 VSUBS 0.034669f
C50 VP.n12 VSUBS 0.034669f
C51 VP.n13 VSUBS 0.064615f
C52 VP.n14 VSUBS 0.042922f
C53 VP.n15 VSUBS 1.10423f
C54 VP.n16 VSUBS 0.056968f
C55 VDD2.t2 VSUBS 0.25257f
C56 VDD2.t3 VSUBS 0.25257f
C57 VDD2.n0 VSUBS 2.66012f
C58 VDD2.t1 VSUBS 0.25257f
C59 VDD2.t0 VSUBS 0.25257f
C60 VDD2.n1 VSUBS 1.99527f
C61 VDD2.n2 VSUBS 4.21942f
C62 VTAIL.n0 VSUBS 0.013325f
C63 VTAIL.n1 VSUBS 0.030006f
C64 VTAIL.n2 VSUBS 0.013442f
C65 VTAIL.n3 VSUBS 0.023625f
C66 VTAIL.n4 VSUBS 0.012695f
C67 VTAIL.n5 VSUBS 0.030006f
C68 VTAIL.n6 VSUBS 0.013442f
C69 VTAIL.n7 VSUBS 0.023625f
C70 VTAIL.n8 VSUBS 0.012695f
C71 VTAIL.n9 VSUBS 0.030006f
C72 VTAIL.n10 VSUBS 0.013442f
C73 VTAIL.n11 VSUBS 0.023625f
C74 VTAIL.n12 VSUBS 0.012695f
C75 VTAIL.n13 VSUBS 0.030006f
C76 VTAIL.n14 VSUBS 0.013442f
C77 VTAIL.n15 VSUBS 0.023625f
C78 VTAIL.n16 VSUBS 0.012695f
C79 VTAIL.n17 VSUBS 0.030006f
C80 VTAIL.n18 VSUBS 0.013442f
C81 VTAIL.n19 VSUBS 1.18352f
C82 VTAIL.n20 VSUBS 0.012695f
C83 VTAIL.t7 VSUBS 0.064063f
C84 VTAIL.n21 VSUBS 0.145425f
C85 VTAIL.n22 VSUBS 0.019089f
C86 VTAIL.n23 VSUBS 0.022505f
C87 VTAIL.n24 VSUBS 0.030006f
C88 VTAIL.n25 VSUBS 0.013442f
C89 VTAIL.n26 VSUBS 0.012695f
C90 VTAIL.n27 VSUBS 0.023625f
C91 VTAIL.n28 VSUBS 0.023625f
C92 VTAIL.n29 VSUBS 0.012695f
C93 VTAIL.n30 VSUBS 0.013442f
C94 VTAIL.n31 VSUBS 0.030006f
C95 VTAIL.n32 VSUBS 0.030006f
C96 VTAIL.n33 VSUBS 0.013442f
C97 VTAIL.n34 VSUBS 0.012695f
C98 VTAIL.n35 VSUBS 0.023625f
C99 VTAIL.n36 VSUBS 0.023625f
C100 VTAIL.n37 VSUBS 0.012695f
C101 VTAIL.n38 VSUBS 0.013442f
C102 VTAIL.n39 VSUBS 0.030006f
C103 VTAIL.n40 VSUBS 0.030006f
C104 VTAIL.n41 VSUBS 0.013442f
C105 VTAIL.n42 VSUBS 0.012695f
C106 VTAIL.n43 VSUBS 0.023625f
C107 VTAIL.n44 VSUBS 0.023625f
C108 VTAIL.n45 VSUBS 0.012695f
C109 VTAIL.n46 VSUBS 0.013442f
C110 VTAIL.n47 VSUBS 0.030006f
C111 VTAIL.n48 VSUBS 0.030006f
C112 VTAIL.n49 VSUBS 0.013442f
C113 VTAIL.n50 VSUBS 0.012695f
C114 VTAIL.n51 VSUBS 0.023625f
C115 VTAIL.n52 VSUBS 0.023625f
C116 VTAIL.n53 VSUBS 0.012695f
C117 VTAIL.n54 VSUBS 0.013442f
C118 VTAIL.n55 VSUBS 0.030006f
C119 VTAIL.n56 VSUBS 0.030006f
C120 VTAIL.n57 VSUBS 0.013442f
C121 VTAIL.n58 VSUBS 0.012695f
C122 VTAIL.n59 VSUBS 0.023625f
C123 VTAIL.n60 VSUBS 0.061385f
C124 VTAIL.n61 VSUBS 0.012695f
C125 VTAIL.n62 VSUBS 0.013442f
C126 VTAIL.n63 VSUBS 0.067189f
C127 VTAIL.n64 VSUBS 0.045128f
C128 VTAIL.n65 VSUBS 0.155641f
C129 VTAIL.n66 VSUBS 0.013325f
C130 VTAIL.n67 VSUBS 0.030006f
C131 VTAIL.n68 VSUBS 0.013442f
C132 VTAIL.n69 VSUBS 0.023625f
C133 VTAIL.n70 VSUBS 0.012695f
C134 VTAIL.n71 VSUBS 0.030006f
C135 VTAIL.n72 VSUBS 0.013442f
C136 VTAIL.n73 VSUBS 0.023625f
C137 VTAIL.n74 VSUBS 0.012695f
C138 VTAIL.n75 VSUBS 0.030006f
C139 VTAIL.n76 VSUBS 0.013442f
C140 VTAIL.n77 VSUBS 0.023625f
C141 VTAIL.n78 VSUBS 0.012695f
C142 VTAIL.n79 VSUBS 0.030006f
C143 VTAIL.n80 VSUBS 0.013442f
C144 VTAIL.n81 VSUBS 0.023625f
C145 VTAIL.n82 VSUBS 0.012695f
C146 VTAIL.n83 VSUBS 0.030006f
C147 VTAIL.n84 VSUBS 0.013442f
C148 VTAIL.n85 VSUBS 1.18352f
C149 VTAIL.n86 VSUBS 0.012695f
C150 VTAIL.t0 VSUBS 0.064063f
C151 VTAIL.n87 VSUBS 0.145425f
C152 VTAIL.n88 VSUBS 0.019089f
C153 VTAIL.n89 VSUBS 0.022505f
C154 VTAIL.n90 VSUBS 0.030006f
C155 VTAIL.n91 VSUBS 0.013442f
C156 VTAIL.n92 VSUBS 0.012695f
C157 VTAIL.n93 VSUBS 0.023625f
C158 VTAIL.n94 VSUBS 0.023625f
C159 VTAIL.n95 VSUBS 0.012695f
C160 VTAIL.n96 VSUBS 0.013442f
C161 VTAIL.n97 VSUBS 0.030006f
C162 VTAIL.n98 VSUBS 0.030006f
C163 VTAIL.n99 VSUBS 0.013442f
C164 VTAIL.n100 VSUBS 0.012695f
C165 VTAIL.n101 VSUBS 0.023625f
C166 VTAIL.n102 VSUBS 0.023625f
C167 VTAIL.n103 VSUBS 0.012695f
C168 VTAIL.n104 VSUBS 0.013442f
C169 VTAIL.n105 VSUBS 0.030006f
C170 VTAIL.n106 VSUBS 0.030006f
C171 VTAIL.n107 VSUBS 0.013442f
C172 VTAIL.n108 VSUBS 0.012695f
C173 VTAIL.n109 VSUBS 0.023625f
C174 VTAIL.n110 VSUBS 0.023625f
C175 VTAIL.n111 VSUBS 0.012695f
C176 VTAIL.n112 VSUBS 0.013442f
C177 VTAIL.n113 VSUBS 0.030006f
C178 VTAIL.n114 VSUBS 0.030006f
C179 VTAIL.n115 VSUBS 0.013442f
C180 VTAIL.n116 VSUBS 0.012695f
C181 VTAIL.n117 VSUBS 0.023625f
C182 VTAIL.n118 VSUBS 0.023625f
C183 VTAIL.n119 VSUBS 0.012695f
C184 VTAIL.n120 VSUBS 0.013442f
C185 VTAIL.n121 VSUBS 0.030006f
C186 VTAIL.n122 VSUBS 0.030006f
C187 VTAIL.n123 VSUBS 0.013442f
C188 VTAIL.n124 VSUBS 0.012695f
C189 VTAIL.n125 VSUBS 0.023625f
C190 VTAIL.n126 VSUBS 0.061385f
C191 VTAIL.n127 VSUBS 0.012695f
C192 VTAIL.n128 VSUBS 0.013442f
C193 VTAIL.n129 VSUBS 0.067189f
C194 VTAIL.n130 VSUBS 0.045128f
C195 VTAIL.n131 VSUBS 0.243742f
C196 VTAIL.n132 VSUBS 0.013325f
C197 VTAIL.n133 VSUBS 0.030006f
C198 VTAIL.n134 VSUBS 0.013442f
C199 VTAIL.n135 VSUBS 0.023625f
C200 VTAIL.n136 VSUBS 0.012695f
C201 VTAIL.n137 VSUBS 0.030006f
C202 VTAIL.n138 VSUBS 0.013442f
C203 VTAIL.n139 VSUBS 0.023625f
C204 VTAIL.n140 VSUBS 0.012695f
C205 VTAIL.n141 VSUBS 0.030006f
C206 VTAIL.n142 VSUBS 0.013442f
C207 VTAIL.n143 VSUBS 0.023625f
C208 VTAIL.n144 VSUBS 0.012695f
C209 VTAIL.n145 VSUBS 0.030006f
C210 VTAIL.n146 VSUBS 0.013442f
C211 VTAIL.n147 VSUBS 0.023625f
C212 VTAIL.n148 VSUBS 0.012695f
C213 VTAIL.n149 VSUBS 0.030006f
C214 VTAIL.n150 VSUBS 0.013442f
C215 VTAIL.n151 VSUBS 1.18352f
C216 VTAIL.n152 VSUBS 0.012695f
C217 VTAIL.t2 VSUBS 0.064063f
C218 VTAIL.n153 VSUBS 0.145425f
C219 VTAIL.n154 VSUBS 0.019089f
C220 VTAIL.n155 VSUBS 0.022505f
C221 VTAIL.n156 VSUBS 0.030006f
C222 VTAIL.n157 VSUBS 0.013442f
C223 VTAIL.n158 VSUBS 0.012695f
C224 VTAIL.n159 VSUBS 0.023625f
C225 VTAIL.n160 VSUBS 0.023625f
C226 VTAIL.n161 VSUBS 0.012695f
C227 VTAIL.n162 VSUBS 0.013442f
C228 VTAIL.n163 VSUBS 0.030006f
C229 VTAIL.n164 VSUBS 0.030006f
C230 VTAIL.n165 VSUBS 0.013442f
C231 VTAIL.n166 VSUBS 0.012695f
C232 VTAIL.n167 VSUBS 0.023625f
C233 VTAIL.n168 VSUBS 0.023625f
C234 VTAIL.n169 VSUBS 0.012695f
C235 VTAIL.n170 VSUBS 0.013442f
C236 VTAIL.n171 VSUBS 0.030006f
C237 VTAIL.n172 VSUBS 0.030006f
C238 VTAIL.n173 VSUBS 0.013442f
C239 VTAIL.n174 VSUBS 0.012695f
C240 VTAIL.n175 VSUBS 0.023625f
C241 VTAIL.n176 VSUBS 0.023625f
C242 VTAIL.n177 VSUBS 0.012695f
C243 VTAIL.n178 VSUBS 0.013442f
C244 VTAIL.n179 VSUBS 0.030006f
C245 VTAIL.n180 VSUBS 0.030006f
C246 VTAIL.n181 VSUBS 0.013442f
C247 VTAIL.n182 VSUBS 0.012695f
C248 VTAIL.n183 VSUBS 0.023625f
C249 VTAIL.n184 VSUBS 0.023625f
C250 VTAIL.n185 VSUBS 0.012695f
C251 VTAIL.n186 VSUBS 0.013442f
C252 VTAIL.n187 VSUBS 0.030006f
C253 VTAIL.n188 VSUBS 0.030006f
C254 VTAIL.n189 VSUBS 0.013442f
C255 VTAIL.n190 VSUBS 0.012695f
C256 VTAIL.n191 VSUBS 0.023625f
C257 VTAIL.n192 VSUBS 0.061385f
C258 VTAIL.n193 VSUBS 0.012695f
C259 VTAIL.n194 VSUBS 0.013442f
C260 VTAIL.n195 VSUBS 0.067189f
C261 VTAIL.n196 VSUBS 0.045128f
C262 VTAIL.n197 VSUBS 1.49948f
C263 VTAIL.n198 VSUBS 0.013325f
C264 VTAIL.n199 VSUBS 0.030006f
C265 VTAIL.n200 VSUBS 0.013442f
C266 VTAIL.n201 VSUBS 0.023625f
C267 VTAIL.n202 VSUBS 0.012695f
C268 VTAIL.n203 VSUBS 0.030006f
C269 VTAIL.n204 VSUBS 0.013442f
C270 VTAIL.n205 VSUBS 0.023625f
C271 VTAIL.n206 VSUBS 0.012695f
C272 VTAIL.n207 VSUBS 0.030006f
C273 VTAIL.n208 VSUBS 0.013442f
C274 VTAIL.n209 VSUBS 0.023625f
C275 VTAIL.n210 VSUBS 0.012695f
C276 VTAIL.n211 VSUBS 0.030006f
C277 VTAIL.n212 VSUBS 0.013442f
C278 VTAIL.n213 VSUBS 0.023625f
C279 VTAIL.n214 VSUBS 0.012695f
C280 VTAIL.n215 VSUBS 0.030006f
C281 VTAIL.n216 VSUBS 0.013442f
C282 VTAIL.n217 VSUBS 1.18352f
C283 VTAIL.n218 VSUBS 0.012695f
C284 VTAIL.t4 VSUBS 0.064063f
C285 VTAIL.n219 VSUBS 0.145425f
C286 VTAIL.n220 VSUBS 0.019089f
C287 VTAIL.n221 VSUBS 0.022505f
C288 VTAIL.n222 VSUBS 0.030006f
C289 VTAIL.n223 VSUBS 0.013442f
C290 VTAIL.n224 VSUBS 0.012695f
C291 VTAIL.n225 VSUBS 0.023625f
C292 VTAIL.n226 VSUBS 0.023625f
C293 VTAIL.n227 VSUBS 0.012695f
C294 VTAIL.n228 VSUBS 0.013442f
C295 VTAIL.n229 VSUBS 0.030006f
C296 VTAIL.n230 VSUBS 0.030006f
C297 VTAIL.n231 VSUBS 0.013442f
C298 VTAIL.n232 VSUBS 0.012695f
C299 VTAIL.n233 VSUBS 0.023625f
C300 VTAIL.n234 VSUBS 0.023625f
C301 VTAIL.n235 VSUBS 0.012695f
C302 VTAIL.n236 VSUBS 0.013442f
C303 VTAIL.n237 VSUBS 0.030006f
C304 VTAIL.n238 VSUBS 0.030006f
C305 VTAIL.n239 VSUBS 0.013442f
C306 VTAIL.n240 VSUBS 0.012695f
C307 VTAIL.n241 VSUBS 0.023625f
C308 VTAIL.n242 VSUBS 0.023625f
C309 VTAIL.n243 VSUBS 0.012695f
C310 VTAIL.n244 VSUBS 0.013442f
C311 VTAIL.n245 VSUBS 0.030006f
C312 VTAIL.n246 VSUBS 0.030006f
C313 VTAIL.n247 VSUBS 0.013442f
C314 VTAIL.n248 VSUBS 0.012695f
C315 VTAIL.n249 VSUBS 0.023625f
C316 VTAIL.n250 VSUBS 0.023625f
C317 VTAIL.n251 VSUBS 0.012695f
C318 VTAIL.n252 VSUBS 0.013442f
C319 VTAIL.n253 VSUBS 0.030006f
C320 VTAIL.n254 VSUBS 0.030006f
C321 VTAIL.n255 VSUBS 0.013442f
C322 VTAIL.n256 VSUBS 0.012695f
C323 VTAIL.n257 VSUBS 0.023625f
C324 VTAIL.n258 VSUBS 0.061385f
C325 VTAIL.n259 VSUBS 0.012695f
C326 VTAIL.n260 VSUBS 0.013442f
C327 VTAIL.n261 VSUBS 0.067189f
C328 VTAIL.n262 VSUBS 0.045128f
C329 VTAIL.n263 VSUBS 1.49948f
C330 VTAIL.n264 VSUBS 0.013325f
C331 VTAIL.n265 VSUBS 0.030006f
C332 VTAIL.n266 VSUBS 0.013442f
C333 VTAIL.n267 VSUBS 0.023625f
C334 VTAIL.n268 VSUBS 0.012695f
C335 VTAIL.n269 VSUBS 0.030006f
C336 VTAIL.n270 VSUBS 0.013442f
C337 VTAIL.n271 VSUBS 0.023625f
C338 VTAIL.n272 VSUBS 0.012695f
C339 VTAIL.n273 VSUBS 0.030006f
C340 VTAIL.n274 VSUBS 0.013442f
C341 VTAIL.n275 VSUBS 0.023625f
C342 VTAIL.n276 VSUBS 0.012695f
C343 VTAIL.n277 VSUBS 0.030006f
C344 VTAIL.n278 VSUBS 0.013442f
C345 VTAIL.n279 VSUBS 0.023625f
C346 VTAIL.n280 VSUBS 0.012695f
C347 VTAIL.n281 VSUBS 0.030006f
C348 VTAIL.n282 VSUBS 0.013442f
C349 VTAIL.n283 VSUBS 1.18352f
C350 VTAIL.n284 VSUBS 0.012695f
C351 VTAIL.t6 VSUBS 0.064063f
C352 VTAIL.n285 VSUBS 0.145425f
C353 VTAIL.n286 VSUBS 0.019089f
C354 VTAIL.n287 VSUBS 0.022505f
C355 VTAIL.n288 VSUBS 0.030006f
C356 VTAIL.n289 VSUBS 0.013442f
C357 VTAIL.n290 VSUBS 0.012695f
C358 VTAIL.n291 VSUBS 0.023625f
C359 VTAIL.n292 VSUBS 0.023625f
C360 VTAIL.n293 VSUBS 0.012695f
C361 VTAIL.n294 VSUBS 0.013442f
C362 VTAIL.n295 VSUBS 0.030006f
C363 VTAIL.n296 VSUBS 0.030006f
C364 VTAIL.n297 VSUBS 0.013442f
C365 VTAIL.n298 VSUBS 0.012695f
C366 VTAIL.n299 VSUBS 0.023625f
C367 VTAIL.n300 VSUBS 0.023625f
C368 VTAIL.n301 VSUBS 0.012695f
C369 VTAIL.n302 VSUBS 0.013442f
C370 VTAIL.n303 VSUBS 0.030006f
C371 VTAIL.n304 VSUBS 0.030006f
C372 VTAIL.n305 VSUBS 0.013442f
C373 VTAIL.n306 VSUBS 0.012695f
C374 VTAIL.n307 VSUBS 0.023625f
C375 VTAIL.n308 VSUBS 0.023625f
C376 VTAIL.n309 VSUBS 0.012695f
C377 VTAIL.n310 VSUBS 0.013442f
C378 VTAIL.n311 VSUBS 0.030006f
C379 VTAIL.n312 VSUBS 0.030006f
C380 VTAIL.n313 VSUBS 0.013442f
C381 VTAIL.n314 VSUBS 0.012695f
C382 VTAIL.n315 VSUBS 0.023625f
C383 VTAIL.n316 VSUBS 0.023625f
C384 VTAIL.n317 VSUBS 0.012695f
C385 VTAIL.n318 VSUBS 0.013442f
C386 VTAIL.n319 VSUBS 0.030006f
C387 VTAIL.n320 VSUBS 0.030006f
C388 VTAIL.n321 VSUBS 0.013442f
C389 VTAIL.n322 VSUBS 0.012695f
C390 VTAIL.n323 VSUBS 0.023625f
C391 VTAIL.n324 VSUBS 0.061385f
C392 VTAIL.n325 VSUBS 0.012695f
C393 VTAIL.n326 VSUBS 0.013442f
C394 VTAIL.n327 VSUBS 0.067189f
C395 VTAIL.n328 VSUBS 0.045128f
C396 VTAIL.n329 VSUBS 0.243742f
C397 VTAIL.n330 VSUBS 0.013325f
C398 VTAIL.n331 VSUBS 0.030006f
C399 VTAIL.n332 VSUBS 0.013442f
C400 VTAIL.n333 VSUBS 0.023625f
C401 VTAIL.n334 VSUBS 0.012695f
C402 VTAIL.n335 VSUBS 0.030006f
C403 VTAIL.n336 VSUBS 0.013442f
C404 VTAIL.n337 VSUBS 0.023625f
C405 VTAIL.n338 VSUBS 0.012695f
C406 VTAIL.n339 VSUBS 0.030006f
C407 VTAIL.n340 VSUBS 0.013442f
C408 VTAIL.n341 VSUBS 0.023625f
C409 VTAIL.n342 VSUBS 0.012695f
C410 VTAIL.n343 VSUBS 0.030006f
C411 VTAIL.n344 VSUBS 0.013442f
C412 VTAIL.n345 VSUBS 0.023625f
C413 VTAIL.n346 VSUBS 0.012695f
C414 VTAIL.n347 VSUBS 0.030006f
C415 VTAIL.n348 VSUBS 0.013442f
C416 VTAIL.n349 VSUBS 1.18352f
C417 VTAIL.n350 VSUBS 0.012695f
C418 VTAIL.t1 VSUBS 0.064063f
C419 VTAIL.n351 VSUBS 0.145425f
C420 VTAIL.n352 VSUBS 0.019089f
C421 VTAIL.n353 VSUBS 0.022505f
C422 VTAIL.n354 VSUBS 0.030006f
C423 VTAIL.n355 VSUBS 0.013442f
C424 VTAIL.n356 VSUBS 0.012695f
C425 VTAIL.n357 VSUBS 0.023625f
C426 VTAIL.n358 VSUBS 0.023625f
C427 VTAIL.n359 VSUBS 0.012695f
C428 VTAIL.n360 VSUBS 0.013442f
C429 VTAIL.n361 VSUBS 0.030006f
C430 VTAIL.n362 VSUBS 0.030006f
C431 VTAIL.n363 VSUBS 0.013442f
C432 VTAIL.n364 VSUBS 0.012695f
C433 VTAIL.n365 VSUBS 0.023625f
C434 VTAIL.n366 VSUBS 0.023625f
C435 VTAIL.n367 VSUBS 0.012695f
C436 VTAIL.n368 VSUBS 0.013442f
C437 VTAIL.n369 VSUBS 0.030006f
C438 VTAIL.n370 VSUBS 0.030006f
C439 VTAIL.n371 VSUBS 0.013442f
C440 VTAIL.n372 VSUBS 0.012695f
C441 VTAIL.n373 VSUBS 0.023625f
C442 VTAIL.n374 VSUBS 0.023625f
C443 VTAIL.n375 VSUBS 0.012695f
C444 VTAIL.n376 VSUBS 0.013442f
C445 VTAIL.n377 VSUBS 0.030006f
C446 VTAIL.n378 VSUBS 0.030006f
C447 VTAIL.n379 VSUBS 0.013442f
C448 VTAIL.n380 VSUBS 0.012695f
C449 VTAIL.n381 VSUBS 0.023625f
C450 VTAIL.n382 VSUBS 0.023625f
C451 VTAIL.n383 VSUBS 0.012695f
C452 VTAIL.n384 VSUBS 0.013442f
C453 VTAIL.n385 VSUBS 0.030006f
C454 VTAIL.n386 VSUBS 0.030006f
C455 VTAIL.n387 VSUBS 0.013442f
C456 VTAIL.n388 VSUBS 0.012695f
C457 VTAIL.n389 VSUBS 0.023625f
C458 VTAIL.n390 VSUBS 0.061385f
C459 VTAIL.n391 VSUBS 0.012695f
C460 VTAIL.n392 VSUBS 0.013442f
C461 VTAIL.n393 VSUBS 0.067189f
C462 VTAIL.n394 VSUBS 0.045128f
C463 VTAIL.n395 VSUBS 0.243742f
C464 VTAIL.n396 VSUBS 0.013325f
C465 VTAIL.n397 VSUBS 0.030006f
C466 VTAIL.n398 VSUBS 0.013442f
C467 VTAIL.n399 VSUBS 0.023625f
C468 VTAIL.n400 VSUBS 0.012695f
C469 VTAIL.n401 VSUBS 0.030006f
C470 VTAIL.n402 VSUBS 0.013442f
C471 VTAIL.n403 VSUBS 0.023625f
C472 VTAIL.n404 VSUBS 0.012695f
C473 VTAIL.n405 VSUBS 0.030006f
C474 VTAIL.n406 VSUBS 0.013442f
C475 VTAIL.n407 VSUBS 0.023625f
C476 VTAIL.n408 VSUBS 0.012695f
C477 VTAIL.n409 VSUBS 0.030006f
C478 VTAIL.n410 VSUBS 0.013442f
C479 VTAIL.n411 VSUBS 0.023625f
C480 VTAIL.n412 VSUBS 0.012695f
C481 VTAIL.n413 VSUBS 0.030006f
C482 VTAIL.n414 VSUBS 0.013442f
C483 VTAIL.n415 VSUBS 1.18352f
C484 VTAIL.n416 VSUBS 0.012695f
C485 VTAIL.t3 VSUBS 0.064063f
C486 VTAIL.n417 VSUBS 0.145425f
C487 VTAIL.n418 VSUBS 0.019089f
C488 VTAIL.n419 VSUBS 0.022505f
C489 VTAIL.n420 VSUBS 0.030006f
C490 VTAIL.n421 VSUBS 0.013442f
C491 VTAIL.n422 VSUBS 0.012695f
C492 VTAIL.n423 VSUBS 0.023625f
C493 VTAIL.n424 VSUBS 0.023625f
C494 VTAIL.n425 VSUBS 0.012695f
C495 VTAIL.n426 VSUBS 0.013442f
C496 VTAIL.n427 VSUBS 0.030006f
C497 VTAIL.n428 VSUBS 0.030006f
C498 VTAIL.n429 VSUBS 0.013442f
C499 VTAIL.n430 VSUBS 0.012695f
C500 VTAIL.n431 VSUBS 0.023625f
C501 VTAIL.n432 VSUBS 0.023625f
C502 VTAIL.n433 VSUBS 0.012695f
C503 VTAIL.n434 VSUBS 0.013442f
C504 VTAIL.n435 VSUBS 0.030006f
C505 VTAIL.n436 VSUBS 0.030006f
C506 VTAIL.n437 VSUBS 0.013442f
C507 VTAIL.n438 VSUBS 0.012695f
C508 VTAIL.n439 VSUBS 0.023625f
C509 VTAIL.n440 VSUBS 0.023625f
C510 VTAIL.n441 VSUBS 0.012695f
C511 VTAIL.n442 VSUBS 0.013442f
C512 VTAIL.n443 VSUBS 0.030006f
C513 VTAIL.n444 VSUBS 0.030006f
C514 VTAIL.n445 VSUBS 0.013442f
C515 VTAIL.n446 VSUBS 0.012695f
C516 VTAIL.n447 VSUBS 0.023625f
C517 VTAIL.n448 VSUBS 0.023625f
C518 VTAIL.n449 VSUBS 0.012695f
C519 VTAIL.n450 VSUBS 0.013442f
C520 VTAIL.n451 VSUBS 0.030006f
C521 VTAIL.n452 VSUBS 0.030006f
C522 VTAIL.n453 VSUBS 0.013442f
C523 VTAIL.n454 VSUBS 0.012695f
C524 VTAIL.n455 VSUBS 0.023625f
C525 VTAIL.n456 VSUBS 0.061385f
C526 VTAIL.n457 VSUBS 0.012695f
C527 VTAIL.n458 VSUBS 0.013442f
C528 VTAIL.n459 VSUBS 0.067189f
C529 VTAIL.n460 VSUBS 0.045128f
C530 VTAIL.n461 VSUBS 1.49948f
C531 VTAIL.n462 VSUBS 0.013325f
C532 VTAIL.n463 VSUBS 0.030006f
C533 VTAIL.n464 VSUBS 0.013442f
C534 VTAIL.n465 VSUBS 0.023625f
C535 VTAIL.n466 VSUBS 0.012695f
C536 VTAIL.n467 VSUBS 0.030006f
C537 VTAIL.n468 VSUBS 0.013442f
C538 VTAIL.n469 VSUBS 0.023625f
C539 VTAIL.n470 VSUBS 0.012695f
C540 VTAIL.n471 VSUBS 0.030006f
C541 VTAIL.n472 VSUBS 0.013442f
C542 VTAIL.n473 VSUBS 0.023625f
C543 VTAIL.n474 VSUBS 0.012695f
C544 VTAIL.n475 VSUBS 0.030006f
C545 VTAIL.n476 VSUBS 0.013442f
C546 VTAIL.n477 VSUBS 0.023625f
C547 VTAIL.n478 VSUBS 0.012695f
C548 VTAIL.n479 VSUBS 0.030006f
C549 VTAIL.n480 VSUBS 0.013442f
C550 VTAIL.n481 VSUBS 1.18352f
C551 VTAIL.n482 VSUBS 0.012695f
C552 VTAIL.t5 VSUBS 0.064063f
C553 VTAIL.n483 VSUBS 0.145425f
C554 VTAIL.n484 VSUBS 0.019089f
C555 VTAIL.n485 VSUBS 0.022505f
C556 VTAIL.n486 VSUBS 0.030006f
C557 VTAIL.n487 VSUBS 0.013442f
C558 VTAIL.n488 VSUBS 0.012695f
C559 VTAIL.n489 VSUBS 0.023625f
C560 VTAIL.n490 VSUBS 0.023625f
C561 VTAIL.n491 VSUBS 0.012695f
C562 VTAIL.n492 VSUBS 0.013442f
C563 VTAIL.n493 VSUBS 0.030006f
C564 VTAIL.n494 VSUBS 0.030006f
C565 VTAIL.n495 VSUBS 0.013442f
C566 VTAIL.n496 VSUBS 0.012695f
C567 VTAIL.n497 VSUBS 0.023625f
C568 VTAIL.n498 VSUBS 0.023625f
C569 VTAIL.n499 VSUBS 0.012695f
C570 VTAIL.n500 VSUBS 0.013442f
C571 VTAIL.n501 VSUBS 0.030006f
C572 VTAIL.n502 VSUBS 0.030006f
C573 VTAIL.n503 VSUBS 0.013442f
C574 VTAIL.n504 VSUBS 0.012695f
C575 VTAIL.n505 VSUBS 0.023625f
C576 VTAIL.n506 VSUBS 0.023625f
C577 VTAIL.n507 VSUBS 0.012695f
C578 VTAIL.n508 VSUBS 0.013442f
C579 VTAIL.n509 VSUBS 0.030006f
C580 VTAIL.n510 VSUBS 0.030006f
C581 VTAIL.n511 VSUBS 0.013442f
C582 VTAIL.n512 VSUBS 0.012695f
C583 VTAIL.n513 VSUBS 0.023625f
C584 VTAIL.n514 VSUBS 0.023625f
C585 VTAIL.n515 VSUBS 0.012695f
C586 VTAIL.n516 VSUBS 0.013442f
C587 VTAIL.n517 VSUBS 0.030006f
C588 VTAIL.n518 VSUBS 0.030006f
C589 VTAIL.n519 VSUBS 0.013442f
C590 VTAIL.n520 VSUBS 0.012695f
C591 VTAIL.n521 VSUBS 0.023625f
C592 VTAIL.n522 VSUBS 0.061385f
C593 VTAIL.n523 VSUBS 0.012695f
C594 VTAIL.n524 VSUBS 0.013442f
C595 VTAIL.n525 VSUBS 0.067189f
C596 VTAIL.n526 VSUBS 0.045128f
C597 VTAIL.n527 VSUBS 1.40252f
C598 VN.t1 VSUBS 3.01571f
C599 VN.t0 VSUBS 3.0099f
C600 VN.n0 VSUBS 1.94536f
C601 VN.t3 VSUBS 3.01571f
C602 VN.t2 VSUBS 3.0099f
C603 VN.n1 VSUBS 3.73496f
C604 B.n0 VSUBS 0.004293f
C605 B.n1 VSUBS 0.004293f
C606 B.n2 VSUBS 0.006789f
C607 B.n3 VSUBS 0.006789f
C608 B.n4 VSUBS 0.006789f
C609 B.n5 VSUBS 0.006789f
C610 B.n6 VSUBS 0.006789f
C611 B.n7 VSUBS 0.006789f
C612 B.n8 VSUBS 0.006789f
C613 B.n9 VSUBS 0.006789f
C614 B.n10 VSUBS 0.006789f
C615 B.n11 VSUBS 0.006789f
C616 B.n12 VSUBS 0.006789f
C617 B.n13 VSUBS 0.006789f
C618 B.n14 VSUBS 0.006789f
C619 B.n15 VSUBS 0.006789f
C620 B.n16 VSUBS 0.006789f
C621 B.n17 VSUBS 0.006789f
C622 B.n18 VSUBS 0.014641f
C623 B.n19 VSUBS 0.006789f
C624 B.n20 VSUBS 0.006789f
C625 B.n21 VSUBS 0.006789f
C626 B.n22 VSUBS 0.006789f
C627 B.n23 VSUBS 0.006789f
C628 B.n24 VSUBS 0.006789f
C629 B.n25 VSUBS 0.006789f
C630 B.n26 VSUBS 0.006789f
C631 B.n27 VSUBS 0.006789f
C632 B.n28 VSUBS 0.006789f
C633 B.n29 VSUBS 0.006789f
C634 B.n30 VSUBS 0.006789f
C635 B.n31 VSUBS 0.006789f
C636 B.n32 VSUBS 0.006789f
C637 B.n33 VSUBS 0.006789f
C638 B.n34 VSUBS 0.006789f
C639 B.n35 VSUBS 0.006789f
C640 B.n36 VSUBS 0.006789f
C641 B.n37 VSUBS 0.006789f
C642 B.n38 VSUBS 0.006789f
C643 B.n39 VSUBS 0.006789f
C644 B.t5 VSUBS 0.203864f
C645 B.t4 VSUBS 0.233637f
C646 B.t3 VSUBS 1.31304f
C647 B.n40 VSUBS 0.370673f
C648 B.n41 VSUBS 0.24357f
C649 B.n42 VSUBS 0.006789f
C650 B.n43 VSUBS 0.006789f
C651 B.n44 VSUBS 0.006789f
C652 B.n45 VSUBS 0.006789f
C653 B.t11 VSUBS 0.203867f
C654 B.t10 VSUBS 0.233639f
C655 B.t9 VSUBS 1.31304f
C656 B.n46 VSUBS 0.37067f
C657 B.n47 VSUBS 0.243567f
C658 B.n48 VSUBS 0.01573f
C659 B.n49 VSUBS 0.006789f
C660 B.n50 VSUBS 0.006789f
C661 B.n51 VSUBS 0.006789f
C662 B.n52 VSUBS 0.006789f
C663 B.n53 VSUBS 0.006789f
C664 B.n54 VSUBS 0.006789f
C665 B.n55 VSUBS 0.006789f
C666 B.n56 VSUBS 0.006789f
C667 B.n57 VSUBS 0.006789f
C668 B.n58 VSUBS 0.006789f
C669 B.n59 VSUBS 0.006789f
C670 B.n60 VSUBS 0.006789f
C671 B.n61 VSUBS 0.006789f
C672 B.n62 VSUBS 0.006789f
C673 B.n63 VSUBS 0.006789f
C674 B.n64 VSUBS 0.006789f
C675 B.n65 VSUBS 0.006789f
C676 B.n66 VSUBS 0.006789f
C677 B.n67 VSUBS 0.006789f
C678 B.n68 VSUBS 0.006789f
C679 B.n69 VSUBS 0.015711f
C680 B.n70 VSUBS 0.006789f
C681 B.n71 VSUBS 0.006789f
C682 B.n72 VSUBS 0.006789f
C683 B.n73 VSUBS 0.006789f
C684 B.n74 VSUBS 0.006789f
C685 B.n75 VSUBS 0.006789f
C686 B.n76 VSUBS 0.006789f
C687 B.n77 VSUBS 0.006789f
C688 B.n78 VSUBS 0.006789f
C689 B.n79 VSUBS 0.006789f
C690 B.n80 VSUBS 0.006789f
C691 B.n81 VSUBS 0.006789f
C692 B.n82 VSUBS 0.006789f
C693 B.n83 VSUBS 0.006789f
C694 B.n84 VSUBS 0.006789f
C695 B.n85 VSUBS 0.006789f
C696 B.n86 VSUBS 0.006789f
C697 B.n87 VSUBS 0.006789f
C698 B.n88 VSUBS 0.006789f
C699 B.n89 VSUBS 0.006789f
C700 B.n90 VSUBS 0.006789f
C701 B.n91 VSUBS 0.006789f
C702 B.n92 VSUBS 0.006789f
C703 B.n93 VSUBS 0.006789f
C704 B.n94 VSUBS 0.006789f
C705 B.n95 VSUBS 0.006789f
C706 B.n96 VSUBS 0.006789f
C707 B.n97 VSUBS 0.006789f
C708 B.n98 VSUBS 0.006789f
C709 B.n99 VSUBS 0.006789f
C710 B.n100 VSUBS 0.006789f
C711 B.n101 VSUBS 0.006789f
C712 B.n102 VSUBS 0.006789f
C713 B.n103 VSUBS 0.015711f
C714 B.n104 VSUBS 0.006789f
C715 B.n105 VSUBS 0.006789f
C716 B.n106 VSUBS 0.006789f
C717 B.n107 VSUBS 0.006789f
C718 B.n108 VSUBS 0.006789f
C719 B.n109 VSUBS 0.006789f
C720 B.n110 VSUBS 0.006789f
C721 B.n111 VSUBS 0.006789f
C722 B.n112 VSUBS 0.006789f
C723 B.n113 VSUBS 0.006789f
C724 B.n114 VSUBS 0.006789f
C725 B.n115 VSUBS 0.006789f
C726 B.n116 VSUBS 0.006789f
C727 B.n117 VSUBS 0.006789f
C728 B.n118 VSUBS 0.006789f
C729 B.n119 VSUBS 0.006789f
C730 B.n120 VSUBS 0.006789f
C731 B.n121 VSUBS 0.006789f
C732 B.n122 VSUBS 0.006789f
C733 B.n123 VSUBS 0.006789f
C734 B.t7 VSUBS 0.203867f
C735 B.t8 VSUBS 0.233639f
C736 B.t6 VSUBS 1.31304f
C737 B.n124 VSUBS 0.37067f
C738 B.n125 VSUBS 0.243567f
C739 B.n126 VSUBS 0.01573f
C740 B.n127 VSUBS 0.006789f
C741 B.n128 VSUBS 0.006789f
C742 B.n129 VSUBS 0.006789f
C743 B.n130 VSUBS 0.006789f
C744 B.n131 VSUBS 0.006789f
C745 B.t1 VSUBS 0.203864f
C746 B.t2 VSUBS 0.233637f
C747 B.t0 VSUBS 1.31304f
C748 B.n132 VSUBS 0.370673f
C749 B.n133 VSUBS 0.24357f
C750 B.n134 VSUBS 0.006789f
C751 B.n135 VSUBS 0.006789f
C752 B.n136 VSUBS 0.006789f
C753 B.n137 VSUBS 0.006789f
C754 B.n138 VSUBS 0.006789f
C755 B.n139 VSUBS 0.006789f
C756 B.n140 VSUBS 0.006789f
C757 B.n141 VSUBS 0.006789f
C758 B.n142 VSUBS 0.006789f
C759 B.n143 VSUBS 0.006789f
C760 B.n144 VSUBS 0.006789f
C761 B.n145 VSUBS 0.006789f
C762 B.n146 VSUBS 0.006789f
C763 B.n147 VSUBS 0.006789f
C764 B.n148 VSUBS 0.006789f
C765 B.n149 VSUBS 0.006789f
C766 B.n150 VSUBS 0.006789f
C767 B.n151 VSUBS 0.006789f
C768 B.n152 VSUBS 0.006789f
C769 B.n153 VSUBS 0.006789f
C770 B.n154 VSUBS 0.014641f
C771 B.n155 VSUBS 0.006789f
C772 B.n156 VSUBS 0.006789f
C773 B.n157 VSUBS 0.006789f
C774 B.n158 VSUBS 0.006789f
C775 B.n159 VSUBS 0.006789f
C776 B.n160 VSUBS 0.006789f
C777 B.n161 VSUBS 0.006789f
C778 B.n162 VSUBS 0.006789f
C779 B.n163 VSUBS 0.006789f
C780 B.n164 VSUBS 0.006789f
C781 B.n165 VSUBS 0.006789f
C782 B.n166 VSUBS 0.006789f
C783 B.n167 VSUBS 0.006789f
C784 B.n168 VSUBS 0.006789f
C785 B.n169 VSUBS 0.006789f
C786 B.n170 VSUBS 0.006789f
C787 B.n171 VSUBS 0.006789f
C788 B.n172 VSUBS 0.006789f
C789 B.n173 VSUBS 0.006789f
C790 B.n174 VSUBS 0.006789f
C791 B.n175 VSUBS 0.006789f
C792 B.n176 VSUBS 0.006789f
C793 B.n177 VSUBS 0.006789f
C794 B.n178 VSUBS 0.006789f
C795 B.n179 VSUBS 0.006789f
C796 B.n180 VSUBS 0.006789f
C797 B.n181 VSUBS 0.006789f
C798 B.n182 VSUBS 0.006789f
C799 B.n183 VSUBS 0.006789f
C800 B.n184 VSUBS 0.006789f
C801 B.n185 VSUBS 0.006789f
C802 B.n186 VSUBS 0.006789f
C803 B.n187 VSUBS 0.006789f
C804 B.n188 VSUBS 0.006789f
C805 B.n189 VSUBS 0.006789f
C806 B.n190 VSUBS 0.006789f
C807 B.n191 VSUBS 0.006789f
C808 B.n192 VSUBS 0.006789f
C809 B.n193 VSUBS 0.006789f
C810 B.n194 VSUBS 0.006789f
C811 B.n195 VSUBS 0.006789f
C812 B.n196 VSUBS 0.006789f
C813 B.n197 VSUBS 0.006789f
C814 B.n198 VSUBS 0.006789f
C815 B.n199 VSUBS 0.006789f
C816 B.n200 VSUBS 0.006789f
C817 B.n201 VSUBS 0.006789f
C818 B.n202 VSUBS 0.006789f
C819 B.n203 VSUBS 0.006789f
C820 B.n204 VSUBS 0.006789f
C821 B.n205 VSUBS 0.006789f
C822 B.n206 VSUBS 0.006789f
C823 B.n207 VSUBS 0.006789f
C824 B.n208 VSUBS 0.006789f
C825 B.n209 VSUBS 0.006789f
C826 B.n210 VSUBS 0.006789f
C827 B.n211 VSUBS 0.006789f
C828 B.n212 VSUBS 0.006789f
C829 B.n213 VSUBS 0.006789f
C830 B.n214 VSUBS 0.006789f
C831 B.n215 VSUBS 0.006789f
C832 B.n216 VSUBS 0.006789f
C833 B.n217 VSUBS 0.014641f
C834 B.n218 VSUBS 0.015711f
C835 B.n219 VSUBS 0.015711f
C836 B.n220 VSUBS 0.006789f
C837 B.n221 VSUBS 0.006789f
C838 B.n222 VSUBS 0.006789f
C839 B.n223 VSUBS 0.006789f
C840 B.n224 VSUBS 0.006789f
C841 B.n225 VSUBS 0.006789f
C842 B.n226 VSUBS 0.006789f
C843 B.n227 VSUBS 0.006789f
C844 B.n228 VSUBS 0.006789f
C845 B.n229 VSUBS 0.006789f
C846 B.n230 VSUBS 0.006789f
C847 B.n231 VSUBS 0.006789f
C848 B.n232 VSUBS 0.006789f
C849 B.n233 VSUBS 0.006789f
C850 B.n234 VSUBS 0.006789f
C851 B.n235 VSUBS 0.006789f
C852 B.n236 VSUBS 0.006789f
C853 B.n237 VSUBS 0.006789f
C854 B.n238 VSUBS 0.006789f
C855 B.n239 VSUBS 0.006789f
C856 B.n240 VSUBS 0.006789f
C857 B.n241 VSUBS 0.006789f
C858 B.n242 VSUBS 0.006789f
C859 B.n243 VSUBS 0.006789f
C860 B.n244 VSUBS 0.006789f
C861 B.n245 VSUBS 0.006789f
C862 B.n246 VSUBS 0.006789f
C863 B.n247 VSUBS 0.006789f
C864 B.n248 VSUBS 0.006789f
C865 B.n249 VSUBS 0.006789f
C866 B.n250 VSUBS 0.006789f
C867 B.n251 VSUBS 0.006789f
C868 B.n252 VSUBS 0.006789f
C869 B.n253 VSUBS 0.006789f
C870 B.n254 VSUBS 0.006789f
C871 B.n255 VSUBS 0.006789f
C872 B.n256 VSUBS 0.006789f
C873 B.n257 VSUBS 0.006789f
C874 B.n258 VSUBS 0.006789f
C875 B.n259 VSUBS 0.006789f
C876 B.n260 VSUBS 0.006789f
C877 B.n261 VSUBS 0.006789f
C878 B.n262 VSUBS 0.006789f
C879 B.n263 VSUBS 0.006789f
C880 B.n264 VSUBS 0.006789f
C881 B.n265 VSUBS 0.006789f
C882 B.n266 VSUBS 0.006789f
C883 B.n267 VSUBS 0.006789f
C884 B.n268 VSUBS 0.006789f
C885 B.n269 VSUBS 0.006789f
C886 B.n270 VSUBS 0.006789f
C887 B.n271 VSUBS 0.006789f
C888 B.n272 VSUBS 0.006789f
C889 B.n273 VSUBS 0.006789f
C890 B.n274 VSUBS 0.006789f
C891 B.n275 VSUBS 0.006789f
C892 B.n276 VSUBS 0.006789f
C893 B.n277 VSUBS 0.006789f
C894 B.n278 VSUBS 0.006789f
C895 B.n279 VSUBS 0.006789f
C896 B.n280 VSUBS 0.004693f
C897 B.n281 VSUBS 0.01573f
C898 B.n282 VSUBS 0.005491f
C899 B.n283 VSUBS 0.006789f
C900 B.n284 VSUBS 0.006789f
C901 B.n285 VSUBS 0.006789f
C902 B.n286 VSUBS 0.006789f
C903 B.n287 VSUBS 0.006789f
C904 B.n288 VSUBS 0.006789f
C905 B.n289 VSUBS 0.006789f
C906 B.n290 VSUBS 0.006789f
C907 B.n291 VSUBS 0.006789f
C908 B.n292 VSUBS 0.006789f
C909 B.n293 VSUBS 0.006789f
C910 B.n294 VSUBS 0.005491f
C911 B.n295 VSUBS 0.006789f
C912 B.n296 VSUBS 0.006789f
C913 B.n297 VSUBS 0.004693f
C914 B.n298 VSUBS 0.006789f
C915 B.n299 VSUBS 0.006789f
C916 B.n300 VSUBS 0.006789f
C917 B.n301 VSUBS 0.006789f
C918 B.n302 VSUBS 0.006789f
C919 B.n303 VSUBS 0.006789f
C920 B.n304 VSUBS 0.006789f
C921 B.n305 VSUBS 0.006789f
C922 B.n306 VSUBS 0.006789f
C923 B.n307 VSUBS 0.006789f
C924 B.n308 VSUBS 0.006789f
C925 B.n309 VSUBS 0.006789f
C926 B.n310 VSUBS 0.006789f
C927 B.n311 VSUBS 0.006789f
C928 B.n312 VSUBS 0.006789f
C929 B.n313 VSUBS 0.006789f
C930 B.n314 VSUBS 0.006789f
C931 B.n315 VSUBS 0.006789f
C932 B.n316 VSUBS 0.006789f
C933 B.n317 VSUBS 0.006789f
C934 B.n318 VSUBS 0.006789f
C935 B.n319 VSUBS 0.006789f
C936 B.n320 VSUBS 0.006789f
C937 B.n321 VSUBS 0.006789f
C938 B.n322 VSUBS 0.006789f
C939 B.n323 VSUBS 0.006789f
C940 B.n324 VSUBS 0.006789f
C941 B.n325 VSUBS 0.006789f
C942 B.n326 VSUBS 0.006789f
C943 B.n327 VSUBS 0.006789f
C944 B.n328 VSUBS 0.006789f
C945 B.n329 VSUBS 0.006789f
C946 B.n330 VSUBS 0.006789f
C947 B.n331 VSUBS 0.006789f
C948 B.n332 VSUBS 0.006789f
C949 B.n333 VSUBS 0.006789f
C950 B.n334 VSUBS 0.006789f
C951 B.n335 VSUBS 0.006789f
C952 B.n336 VSUBS 0.006789f
C953 B.n337 VSUBS 0.006789f
C954 B.n338 VSUBS 0.006789f
C955 B.n339 VSUBS 0.006789f
C956 B.n340 VSUBS 0.006789f
C957 B.n341 VSUBS 0.006789f
C958 B.n342 VSUBS 0.006789f
C959 B.n343 VSUBS 0.006789f
C960 B.n344 VSUBS 0.006789f
C961 B.n345 VSUBS 0.006789f
C962 B.n346 VSUBS 0.006789f
C963 B.n347 VSUBS 0.006789f
C964 B.n348 VSUBS 0.006789f
C965 B.n349 VSUBS 0.006789f
C966 B.n350 VSUBS 0.006789f
C967 B.n351 VSUBS 0.006789f
C968 B.n352 VSUBS 0.006789f
C969 B.n353 VSUBS 0.006789f
C970 B.n354 VSUBS 0.006789f
C971 B.n355 VSUBS 0.006789f
C972 B.n356 VSUBS 0.006789f
C973 B.n357 VSUBS 0.006789f
C974 B.n358 VSUBS 0.015711f
C975 B.n359 VSUBS 0.014641f
C976 B.n360 VSUBS 0.014641f
C977 B.n361 VSUBS 0.006789f
C978 B.n362 VSUBS 0.006789f
C979 B.n363 VSUBS 0.006789f
C980 B.n364 VSUBS 0.006789f
C981 B.n365 VSUBS 0.006789f
C982 B.n366 VSUBS 0.006789f
C983 B.n367 VSUBS 0.006789f
C984 B.n368 VSUBS 0.006789f
C985 B.n369 VSUBS 0.006789f
C986 B.n370 VSUBS 0.006789f
C987 B.n371 VSUBS 0.006789f
C988 B.n372 VSUBS 0.006789f
C989 B.n373 VSUBS 0.006789f
C990 B.n374 VSUBS 0.006789f
C991 B.n375 VSUBS 0.006789f
C992 B.n376 VSUBS 0.006789f
C993 B.n377 VSUBS 0.006789f
C994 B.n378 VSUBS 0.006789f
C995 B.n379 VSUBS 0.006789f
C996 B.n380 VSUBS 0.006789f
C997 B.n381 VSUBS 0.006789f
C998 B.n382 VSUBS 0.006789f
C999 B.n383 VSUBS 0.006789f
C1000 B.n384 VSUBS 0.006789f
C1001 B.n385 VSUBS 0.006789f
C1002 B.n386 VSUBS 0.006789f
C1003 B.n387 VSUBS 0.006789f
C1004 B.n388 VSUBS 0.006789f
C1005 B.n389 VSUBS 0.006789f
C1006 B.n390 VSUBS 0.006789f
C1007 B.n391 VSUBS 0.006789f
C1008 B.n392 VSUBS 0.006789f
C1009 B.n393 VSUBS 0.006789f
C1010 B.n394 VSUBS 0.006789f
C1011 B.n395 VSUBS 0.006789f
C1012 B.n396 VSUBS 0.006789f
C1013 B.n397 VSUBS 0.006789f
C1014 B.n398 VSUBS 0.006789f
C1015 B.n399 VSUBS 0.006789f
C1016 B.n400 VSUBS 0.006789f
C1017 B.n401 VSUBS 0.006789f
C1018 B.n402 VSUBS 0.006789f
C1019 B.n403 VSUBS 0.006789f
C1020 B.n404 VSUBS 0.006789f
C1021 B.n405 VSUBS 0.006789f
C1022 B.n406 VSUBS 0.006789f
C1023 B.n407 VSUBS 0.006789f
C1024 B.n408 VSUBS 0.006789f
C1025 B.n409 VSUBS 0.006789f
C1026 B.n410 VSUBS 0.006789f
C1027 B.n411 VSUBS 0.006789f
C1028 B.n412 VSUBS 0.006789f
C1029 B.n413 VSUBS 0.006789f
C1030 B.n414 VSUBS 0.006789f
C1031 B.n415 VSUBS 0.006789f
C1032 B.n416 VSUBS 0.006789f
C1033 B.n417 VSUBS 0.006789f
C1034 B.n418 VSUBS 0.006789f
C1035 B.n419 VSUBS 0.006789f
C1036 B.n420 VSUBS 0.006789f
C1037 B.n421 VSUBS 0.006789f
C1038 B.n422 VSUBS 0.006789f
C1039 B.n423 VSUBS 0.006789f
C1040 B.n424 VSUBS 0.006789f
C1041 B.n425 VSUBS 0.006789f
C1042 B.n426 VSUBS 0.006789f
C1043 B.n427 VSUBS 0.006789f
C1044 B.n428 VSUBS 0.006789f
C1045 B.n429 VSUBS 0.006789f
C1046 B.n430 VSUBS 0.006789f
C1047 B.n431 VSUBS 0.006789f
C1048 B.n432 VSUBS 0.006789f
C1049 B.n433 VSUBS 0.006789f
C1050 B.n434 VSUBS 0.006789f
C1051 B.n435 VSUBS 0.006789f
C1052 B.n436 VSUBS 0.006789f
C1053 B.n437 VSUBS 0.006789f
C1054 B.n438 VSUBS 0.006789f
C1055 B.n439 VSUBS 0.006789f
C1056 B.n440 VSUBS 0.006789f
C1057 B.n441 VSUBS 0.006789f
C1058 B.n442 VSUBS 0.006789f
C1059 B.n443 VSUBS 0.006789f
C1060 B.n444 VSUBS 0.006789f
C1061 B.n445 VSUBS 0.006789f
C1062 B.n446 VSUBS 0.006789f
C1063 B.n447 VSUBS 0.006789f
C1064 B.n448 VSUBS 0.006789f
C1065 B.n449 VSUBS 0.006789f
C1066 B.n450 VSUBS 0.006789f
C1067 B.n451 VSUBS 0.006789f
C1068 B.n452 VSUBS 0.006789f
C1069 B.n453 VSUBS 0.006789f
C1070 B.n454 VSUBS 0.006789f
C1071 B.n455 VSUBS 0.006789f
C1072 B.n456 VSUBS 0.006789f
C1073 B.n457 VSUBS 0.006789f
C1074 B.n458 VSUBS 0.014641f
C1075 B.n459 VSUBS 0.015502f
C1076 B.n460 VSUBS 0.014851f
C1077 B.n461 VSUBS 0.006789f
C1078 B.n462 VSUBS 0.006789f
C1079 B.n463 VSUBS 0.006789f
C1080 B.n464 VSUBS 0.006789f
C1081 B.n465 VSUBS 0.006789f
C1082 B.n466 VSUBS 0.006789f
C1083 B.n467 VSUBS 0.006789f
C1084 B.n468 VSUBS 0.006789f
C1085 B.n469 VSUBS 0.006789f
C1086 B.n470 VSUBS 0.006789f
C1087 B.n471 VSUBS 0.006789f
C1088 B.n472 VSUBS 0.006789f
C1089 B.n473 VSUBS 0.006789f
C1090 B.n474 VSUBS 0.006789f
C1091 B.n475 VSUBS 0.006789f
C1092 B.n476 VSUBS 0.006789f
C1093 B.n477 VSUBS 0.006789f
C1094 B.n478 VSUBS 0.006789f
C1095 B.n479 VSUBS 0.006789f
C1096 B.n480 VSUBS 0.006789f
C1097 B.n481 VSUBS 0.006789f
C1098 B.n482 VSUBS 0.006789f
C1099 B.n483 VSUBS 0.006789f
C1100 B.n484 VSUBS 0.006789f
C1101 B.n485 VSUBS 0.006789f
C1102 B.n486 VSUBS 0.006789f
C1103 B.n487 VSUBS 0.006789f
C1104 B.n488 VSUBS 0.006789f
C1105 B.n489 VSUBS 0.006789f
C1106 B.n490 VSUBS 0.006789f
C1107 B.n491 VSUBS 0.006789f
C1108 B.n492 VSUBS 0.006789f
C1109 B.n493 VSUBS 0.006789f
C1110 B.n494 VSUBS 0.006789f
C1111 B.n495 VSUBS 0.006789f
C1112 B.n496 VSUBS 0.006789f
C1113 B.n497 VSUBS 0.006789f
C1114 B.n498 VSUBS 0.006789f
C1115 B.n499 VSUBS 0.006789f
C1116 B.n500 VSUBS 0.006789f
C1117 B.n501 VSUBS 0.006789f
C1118 B.n502 VSUBS 0.006789f
C1119 B.n503 VSUBS 0.006789f
C1120 B.n504 VSUBS 0.006789f
C1121 B.n505 VSUBS 0.006789f
C1122 B.n506 VSUBS 0.006789f
C1123 B.n507 VSUBS 0.006789f
C1124 B.n508 VSUBS 0.006789f
C1125 B.n509 VSUBS 0.006789f
C1126 B.n510 VSUBS 0.006789f
C1127 B.n511 VSUBS 0.006789f
C1128 B.n512 VSUBS 0.006789f
C1129 B.n513 VSUBS 0.006789f
C1130 B.n514 VSUBS 0.006789f
C1131 B.n515 VSUBS 0.006789f
C1132 B.n516 VSUBS 0.006789f
C1133 B.n517 VSUBS 0.006789f
C1134 B.n518 VSUBS 0.006789f
C1135 B.n519 VSUBS 0.006789f
C1136 B.n520 VSUBS 0.006789f
C1137 B.n521 VSUBS 0.004693f
C1138 B.n522 VSUBS 0.006789f
C1139 B.n523 VSUBS 0.006789f
C1140 B.n524 VSUBS 0.005491f
C1141 B.n525 VSUBS 0.006789f
C1142 B.n526 VSUBS 0.006789f
C1143 B.n527 VSUBS 0.006789f
C1144 B.n528 VSUBS 0.006789f
C1145 B.n529 VSUBS 0.006789f
C1146 B.n530 VSUBS 0.006789f
C1147 B.n531 VSUBS 0.006789f
C1148 B.n532 VSUBS 0.006789f
C1149 B.n533 VSUBS 0.006789f
C1150 B.n534 VSUBS 0.006789f
C1151 B.n535 VSUBS 0.006789f
C1152 B.n536 VSUBS 0.005491f
C1153 B.n537 VSUBS 0.01573f
C1154 B.n538 VSUBS 0.004693f
C1155 B.n539 VSUBS 0.006789f
C1156 B.n540 VSUBS 0.006789f
C1157 B.n541 VSUBS 0.006789f
C1158 B.n542 VSUBS 0.006789f
C1159 B.n543 VSUBS 0.006789f
C1160 B.n544 VSUBS 0.006789f
C1161 B.n545 VSUBS 0.006789f
C1162 B.n546 VSUBS 0.006789f
C1163 B.n547 VSUBS 0.006789f
C1164 B.n548 VSUBS 0.006789f
C1165 B.n549 VSUBS 0.006789f
C1166 B.n550 VSUBS 0.006789f
C1167 B.n551 VSUBS 0.006789f
C1168 B.n552 VSUBS 0.006789f
C1169 B.n553 VSUBS 0.006789f
C1170 B.n554 VSUBS 0.006789f
C1171 B.n555 VSUBS 0.006789f
C1172 B.n556 VSUBS 0.006789f
C1173 B.n557 VSUBS 0.006789f
C1174 B.n558 VSUBS 0.006789f
C1175 B.n559 VSUBS 0.006789f
C1176 B.n560 VSUBS 0.006789f
C1177 B.n561 VSUBS 0.006789f
C1178 B.n562 VSUBS 0.006789f
C1179 B.n563 VSUBS 0.006789f
C1180 B.n564 VSUBS 0.006789f
C1181 B.n565 VSUBS 0.006789f
C1182 B.n566 VSUBS 0.006789f
C1183 B.n567 VSUBS 0.006789f
C1184 B.n568 VSUBS 0.006789f
C1185 B.n569 VSUBS 0.006789f
C1186 B.n570 VSUBS 0.006789f
C1187 B.n571 VSUBS 0.006789f
C1188 B.n572 VSUBS 0.006789f
C1189 B.n573 VSUBS 0.006789f
C1190 B.n574 VSUBS 0.006789f
C1191 B.n575 VSUBS 0.006789f
C1192 B.n576 VSUBS 0.006789f
C1193 B.n577 VSUBS 0.006789f
C1194 B.n578 VSUBS 0.006789f
C1195 B.n579 VSUBS 0.006789f
C1196 B.n580 VSUBS 0.006789f
C1197 B.n581 VSUBS 0.006789f
C1198 B.n582 VSUBS 0.006789f
C1199 B.n583 VSUBS 0.006789f
C1200 B.n584 VSUBS 0.006789f
C1201 B.n585 VSUBS 0.006789f
C1202 B.n586 VSUBS 0.006789f
C1203 B.n587 VSUBS 0.006789f
C1204 B.n588 VSUBS 0.006789f
C1205 B.n589 VSUBS 0.006789f
C1206 B.n590 VSUBS 0.006789f
C1207 B.n591 VSUBS 0.006789f
C1208 B.n592 VSUBS 0.006789f
C1209 B.n593 VSUBS 0.006789f
C1210 B.n594 VSUBS 0.006789f
C1211 B.n595 VSUBS 0.006789f
C1212 B.n596 VSUBS 0.006789f
C1213 B.n597 VSUBS 0.006789f
C1214 B.n598 VSUBS 0.006789f
C1215 B.n599 VSUBS 0.015711f
C1216 B.n600 VSUBS 0.015711f
C1217 B.n601 VSUBS 0.014641f
C1218 B.n602 VSUBS 0.006789f
C1219 B.n603 VSUBS 0.006789f
C1220 B.n604 VSUBS 0.006789f
C1221 B.n605 VSUBS 0.006789f
C1222 B.n606 VSUBS 0.006789f
C1223 B.n607 VSUBS 0.006789f
C1224 B.n608 VSUBS 0.006789f
C1225 B.n609 VSUBS 0.006789f
C1226 B.n610 VSUBS 0.006789f
C1227 B.n611 VSUBS 0.006789f
C1228 B.n612 VSUBS 0.006789f
C1229 B.n613 VSUBS 0.006789f
C1230 B.n614 VSUBS 0.006789f
C1231 B.n615 VSUBS 0.006789f
C1232 B.n616 VSUBS 0.006789f
C1233 B.n617 VSUBS 0.006789f
C1234 B.n618 VSUBS 0.006789f
C1235 B.n619 VSUBS 0.006789f
C1236 B.n620 VSUBS 0.006789f
C1237 B.n621 VSUBS 0.006789f
C1238 B.n622 VSUBS 0.006789f
C1239 B.n623 VSUBS 0.006789f
C1240 B.n624 VSUBS 0.006789f
C1241 B.n625 VSUBS 0.006789f
C1242 B.n626 VSUBS 0.006789f
C1243 B.n627 VSUBS 0.006789f
C1244 B.n628 VSUBS 0.006789f
C1245 B.n629 VSUBS 0.006789f
C1246 B.n630 VSUBS 0.006789f
C1247 B.n631 VSUBS 0.006789f
C1248 B.n632 VSUBS 0.006789f
C1249 B.n633 VSUBS 0.006789f
C1250 B.n634 VSUBS 0.006789f
C1251 B.n635 VSUBS 0.006789f
C1252 B.n636 VSUBS 0.006789f
C1253 B.n637 VSUBS 0.006789f
C1254 B.n638 VSUBS 0.006789f
C1255 B.n639 VSUBS 0.006789f
C1256 B.n640 VSUBS 0.006789f
C1257 B.n641 VSUBS 0.006789f
C1258 B.n642 VSUBS 0.006789f
C1259 B.n643 VSUBS 0.006789f
C1260 B.n644 VSUBS 0.006789f
C1261 B.n645 VSUBS 0.006789f
C1262 B.n646 VSUBS 0.006789f
C1263 B.n647 VSUBS 0.006789f
C1264 B.n648 VSUBS 0.006789f
C1265 B.n649 VSUBS 0.006789f
C1266 B.n650 VSUBS 0.006789f
C1267 B.n651 VSUBS 0.015373f
.ends

