* NGSPICE file created from diff_pair_sample_1101.ext - technology: sky130A

.subckt diff_pair_sample_1101 VTAIL VN VP B VDD2 VDD1
X0 B.t23 B.t21 B.t22 B.t15 sky130_fd_pr__nfet_01v8 ad=2.8158 pd=15.22 as=0 ps=0 w=7.22 l=1.19
X1 VDD2.t9 VN.t0 VTAIL.t13 B.t6 sky130_fd_pr__nfet_01v8 ad=2.8158 pd=15.22 as=1.1913 ps=7.55 w=7.22 l=1.19
X2 VDD1.t9 VP.t0 VTAIL.t3 B.t7 sky130_fd_pr__nfet_01v8 ad=1.1913 pd=7.55 as=2.8158 ps=15.22 w=7.22 l=1.19
X3 VTAIL.t18 VN.t1 VDD2.t8 B.t4 sky130_fd_pr__nfet_01v8 ad=1.1913 pd=7.55 as=1.1913 ps=7.55 w=7.22 l=1.19
X4 VTAIL.t10 VN.t2 VDD2.t7 B.t2 sky130_fd_pr__nfet_01v8 ad=1.1913 pd=7.55 as=1.1913 ps=7.55 w=7.22 l=1.19
X5 VDD1.t8 VP.t1 VTAIL.t5 B.t8 sky130_fd_pr__nfet_01v8 ad=1.1913 pd=7.55 as=1.1913 ps=7.55 w=7.22 l=1.19
X6 VDD2.t6 VN.t3 VTAIL.t14 B.t5 sky130_fd_pr__nfet_01v8 ad=1.1913 pd=7.55 as=1.1913 ps=7.55 w=7.22 l=1.19
X7 B.t20 B.t18 B.t19 B.t11 sky130_fd_pr__nfet_01v8 ad=2.8158 pd=15.22 as=0 ps=0 w=7.22 l=1.19
X8 VTAIL.t2 VP.t2 VDD1.t7 B.t4 sky130_fd_pr__nfet_01v8 ad=1.1913 pd=7.55 as=1.1913 ps=7.55 w=7.22 l=1.19
X9 VTAIL.t9 VP.t3 VDD1.t6 B.t9 sky130_fd_pr__nfet_01v8 ad=1.1913 pd=7.55 as=1.1913 ps=7.55 w=7.22 l=1.19
X10 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=2.8158 pd=15.22 as=0 ps=0 w=7.22 l=1.19
X11 VTAIL.t11 VN.t4 VDD2.t5 B.t9 sky130_fd_pr__nfet_01v8 ad=1.1913 pd=7.55 as=1.1913 ps=7.55 w=7.22 l=1.19
X12 VTAIL.t15 VN.t5 VDD2.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=1.1913 pd=7.55 as=1.1913 ps=7.55 w=7.22 l=1.19
X13 VDD1.t5 VP.t4 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=2.8158 pd=15.22 as=1.1913 ps=7.55 w=7.22 l=1.19
X14 VTAIL.t1 VP.t5 VDD1.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=1.1913 pd=7.55 as=1.1913 ps=7.55 w=7.22 l=1.19
X15 VDD2.t3 VN.t6 VTAIL.t12 B.t7 sky130_fd_pr__nfet_01v8 ad=1.1913 pd=7.55 as=2.8158 ps=15.22 w=7.22 l=1.19
X16 VDD2.t2 VN.t7 VTAIL.t19 B.t3 sky130_fd_pr__nfet_01v8 ad=1.1913 pd=7.55 as=2.8158 ps=15.22 w=7.22 l=1.19
X17 VDD1.t3 VP.t6 VTAIL.t8 B.t3 sky130_fd_pr__nfet_01v8 ad=1.1913 pd=7.55 as=2.8158 ps=15.22 w=7.22 l=1.19
X18 VDD1.t2 VP.t7 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.8158 pd=15.22 as=1.1913 ps=7.55 w=7.22 l=1.19
X19 VTAIL.t7 VP.t8 VDD1.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=1.1913 pd=7.55 as=1.1913 ps=7.55 w=7.22 l=1.19
X20 VDD2.t1 VN.t8 VTAIL.t17 B.t8 sky130_fd_pr__nfet_01v8 ad=1.1913 pd=7.55 as=1.1913 ps=7.55 w=7.22 l=1.19
X21 VDD1.t0 VP.t9 VTAIL.t4 B.t5 sky130_fd_pr__nfet_01v8 ad=1.1913 pd=7.55 as=1.1913 ps=7.55 w=7.22 l=1.19
X22 VDD2.t0 VN.t9 VTAIL.t16 B.t0 sky130_fd_pr__nfet_01v8 ad=2.8158 pd=15.22 as=1.1913 ps=7.55 w=7.22 l=1.19
X23 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=2.8158 pd=15.22 as=0 ps=0 w=7.22 l=1.19
R0 B.n616 B.n615 585
R1 B.n617 B.n616 585
R2 B.n229 B.n99 585
R3 B.n228 B.n227 585
R4 B.n226 B.n225 585
R5 B.n224 B.n223 585
R6 B.n222 B.n221 585
R7 B.n220 B.n219 585
R8 B.n218 B.n217 585
R9 B.n216 B.n215 585
R10 B.n214 B.n213 585
R11 B.n212 B.n211 585
R12 B.n210 B.n209 585
R13 B.n208 B.n207 585
R14 B.n206 B.n205 585
R15 B.n204 B.n203 585
R16 B.n202 B.n201 585
R17 B.n200 B.n199 585
R18 B.n198 B.n197 585
R19 B.n196 B.n195 585
R20 B.n194 B.n193 585
R21 B.n192 B.n191 585
R22 B.n190 B.n189 585
R23 B.n188 B.n187 585
R24 B.n186 B.n185 585
R25 B.n184 B.n183 585
R26 B.n182 B.n181 585
R27 B.n180 B.n179 585
R28 B.n178 B.n177 585
R29 B.n175 B.n174 585
R30 B.n173 B.n172 585
R31 B.n171 B.n170 585
R32 B.n169 B.n168 585
R33 B.n167 B.n166 585
R34 B.n165 B.n164 585
R35 B.n163 B.n162 585
R36 B.n161 B.n160 585
R37 B.n159 B.n158 585
R38 B.n157 B.n156 585
R39 B.n155 B.n154 585
R40 B.n153 B.n152 585
R41 B.n151 B.n150 585
R42 B.n149 B.n148 585
R43 B.n147 B.n146 585
R44 B.n145 B.n144 585
R45 B.n143 B.n142 585
R46 B.n141 B.n140 585
R47 B.n139 B.n138 585
R48 B.n137 B.n136 585
R49 B.n135 B.n134 585
R50 B.n133 B.n132 585
R51 B.n131 B.n130 585
R52 B.n129 B.n128 585
R53 B.n127 B.n126 585
R54 B.n125 B.n124 585
R55 B.n123 B.n122 585
R56 B.n121 B.n120 585
R57 B.n119 B.n118 585
R58 B.n117 B.n116 585
R59 B.n115 B.n114 585
R60 B.n113 B.n112 585
R61 B.n111 B.n110 585
R62 B.n109 B.n108 585
R63 B.n107 B.n106 585
R64 B.n67 B.n66 585
R65 B.n620 B.n619 585
R66 B.n614 B.n100 585
R67 B.n100 B.n64 585
R68 B.n613 B.n63 585
R69 B.n624 B.n63 585
R70 B.n612 B.n62 585
R71 B.n625 B.n62 585
R72 B.n611 B.n61 585
R73 B.n626 B.n61 585
R74 B.n610 B.n609 585
R75 B.n609 B.n57 585
R76 B.n608 B.n56 585
R77 B.n632 B.n56 585
R78 B.n607 B.n55 585
R79 B.n633 B.n55 585
R80 B.n606 B.n54 585
R81 B.n634 B.n54 585
R82 B.n605 B.n604 585
R83 B.n604 B.n50 585
R84 B.n603 B.n49 585
R85 B.n640 B.n49 585
R86 B.n602 B.n48 585
R87 B.n641 B.n48 585
R88 B.n601 B.n47 585
R89 B.n642 B.n47 585
R90 B.n600 B.n599 585
R91 B.n599 B.n43 585
R92 B.n598 B.n42 585
R93 B.n648 B.n42 585
R94 B.n597 B.n41 585
R95 B.n649 B.n41 585
R96 B.n596 B.n40 585
R97 B.n650 B.n40 585
R98 B.n595 B.n594 585
R99 B.n594 B.n36 585
R100 B.n593 B.n35 585
R101 B.n656 B.n35 585
R102 B.n592 B.n34 585
R103 B.n657 B.n34 585
R104 B.n591 B.n33 585
R105 B.n658 B.n33 585
R106 B.n590 B.n589 585
R107 B.n589 B.n29 585
R108 B.n588 B.n28 585
R109 B.n664 B.n28 585
R110 B.n587 B.n27 585
R111 B.n665 B.n27 585
R112 B.n586 B.n26 585
R113 B.n666 B.n26 585
R114 B.n585 B.n584 585
R115 B.n584 B.n22 585
R116 B.n583 B.n21 585
R117 B.n672 B.n21 585
R118 B.n582 B.n20 585
R119 B.n673 B.n20 585
R120 B.n581 B.n19 585
R121 B.n674 B.n19 585
R122 B.n580 B.n579 585
R123 B.n579 B.n15 585
R124 B.n578 B.n14 585
R125 B.n680 B.n14 585
R126 B.n577 B.n13 585
R127 B.n681 B.n13 585
R128 B.n576 B.n12 585
R129 B.n682 B.n12 585
R130 B.n575 B.n574 585
R131 B.n574 B.n8 585
R132 B.n573 B.n7 585
R133 B.n688 B.n7 585
R134 B.n572 B.n6 585
R135 B.n689 B.n6 585
R136 B.n571 B.n5 585
R137 B.n690 B.n5 585
R138 B.n570 B.n569 585
R139 B.n569 B.n4 585
R140 B.n568 B.n230 585
R141 B.n568 B.n567 585
R142 B.n558 B.n231 585
R143 B.n232 B.n231 585
R144 B.n560 B.n559 585
R145 B.n561 B.n560 585
R146 B.n557 B.n237 585
R147 B.n237 B.n236 585
R148 B.n556 B.n555 585
R149 B.n555 B.n554 585
R150 B.n239 B.n238 585
R151 B.n240 B.n239 585
R152 B.n547 B.n546 585
R153 B.n548 B.n547 585
R154 B.n545 B.n244 585
R155 B.n248 B.n244 585
R156 B.n544 B.n543 585
R157 B.n543 B.n542 585
R158 B.n246 B.n245 585
R159 B.n247 B.n246 585
R160 B.n535 B.n534 585
R161 B.n536 B.n535 585
R162 B.n533 B.n252 585
R163 B.n256 B.n252 585
R164 B.n532 B.n531 585
R165 B.n531 B.n530 585
R166 B.n254 B.n253 585
R167 B.n255 B.n254 585
R168 B.n523 B.n522 585
R169 B.n524 B.n523 585
R170 B.n521 B.n261 585
R171 B.n261 B.n260 585
R172 B.n520 B.n519 585
R173 B.n519 B.n518 585
R174 B.n263 B.n262 585
R175 B.n264 B.n263 585
R176 B.n511 B.n510 585
R177 B.n512 B.n511 585
R178 B.n509 B.n269 585
R179 B.n269 B.n268 585
R180 B.n508 B.n507 585
R181 B.n507 B.n506 585
R182 B.n271 B.n270 585
R183 B.n272 B.n271 585
R184 B.n499 B.n498 585
R185 B.n500 B.n499 585
R186 B.n497 B.n277 585
R187 B.n277 B.n276 585
R188 B.n496 B.n495 585
R189 B.n495 B.n494 585
R190 B.n279 B.n278 585
R191 B.n280 B.n279 585
R192 B.n487 B.n486 585
R193 B.n488 B.n487 585
R194 B.n485 B.n285 585
R195 B.n285 B.n284 585
R196 B.n484 B.n483 585
R197 B.n483 B.n482 585
R198 B.n287 B.n286 585
R199 B.n288 B.n287 585
R200 B.n475 B.n474 585
R201 B.n476 B.n475 585
R202 B.n473 B.n293 585
R203 B.n293 B.n292 585
R204 B.n472 B.n471 585
R205 B.n471 B.n470 585
R206 B.n295 B.n294 585
R207 B.n296 B.n295 585
R208 B.n466 B.n465 585
R209 B.n299 B.n298 585
R210 B.n462 B.n461 585
R211 B.n463 B.n462 585
R212 B.n460 B.n331 585
R213 B.n459 B.n458 585
R214 B.n457 B.n456 585
R215 B.n455 B.n454 585
R216 B.n453 B.n452 585
R217 B.n451 B.n450 585
R218 B.n449 B.n448 585
R219 B.n447 B.n446 585
R220 B.n445 B.n444 585
R221 B.n443 B.n442 585
R222 B.n441 B.n440 585
R223 B.n439 B.n438 585
R224 B.n437 B.n436 585
R225 B.n435 B.n434 585
R226 B.n433 B.n432 585
R227 B.n431 B.n430 585
R228 B.n429 B.n428 585
R229 B.n427 B.n426 585
R230 B.n425 B.n424 585
R231 B.n423 B.n422 585
R232 B.n421 B.n420 585
R233 B.n419 B.n418 585
R234 B.n417 B.n416 585
R235 B.n415 B.n414 585
R236 B.n413 B.n412 585
R237 B.n410 B.n409 585
R238 B.n408 B.n407 585
R239 B.n406 B.n405 585
R240 B.n404 B.n403 585
R241 B.n402 B.n401 585
R242 B.n400 B.n399 585
R243 B.n398 B.n397 585
R244 B.n396 B.n395 585
R245 B.n394 B.n393 585
R246 B.n392 B.n391 585
R247 B.n390 B.n389 585
R248 B.n388 B.n387 585
R249 B.n386 B.n385 585
R250 B.n384 B.n383 585
R251 B.n382 B.n381 585
R252 B.n380 B.n379 585
R253 B.n378 B.n377 585
R254 B.n376 B.n375 585
R255 B.n374 B.n373 585
R256 B.n372 B.n371 585
R257 B.n370 B.n369 585
R258 B.n368 B.n367 585
R259 B.n366 B.n365 585
R260 B.n364 B.n363 585
R261 B.n362 B.n361 585
R262 B.n360 B.n359 585
R263 B.n358 B.n357 585
R264 B.n356 B.n355 585
R265 B.n354 B.n353 585
R266 B.n352 B.n351 585
R267 B.n350 B.n349 585
R268 B.n348 B.n347 585
R269 B.n346 B.n345 585
R270 B.n344 B.n343 585
R271 B.n342 B.n341 585
R272 B.n340 B.n339 585
R273 B.n338 B.n337 585
R274 B.n467 B.n297 585
R275 B.n297 B.n296 585
R276 B.n469 B.n468 585
R277 B.n470 B.n469 585
R278 B.n291 B.n290 585
R279 B.n292 B.n291 585
R280 B.n478 B.n477 585
R281 B.n477 B.n476 585
R282 B.n479 B.n289 585
R283 B.n289 B.n288 585
R284 B.n481 B.n480 585
R285 B.n482 B.n481 585
R286 B.n283 B.n282 585
R287 B.n284 B.n283 585
R288 B.n490 B.n489 585
R289 B.n489 B.n488 585
R290 B.n491 B.n281 585
R291 B.n281 B.n280 585
R292 B.n493 B.n492 585
R293 B.n494 B.n493 585
R294 B.n275 B.n274 585
R295 B.n276 B.n275 585
R296 B.n502 B.n501 585
R297 B.n501 B.n500 585
R298 B.n503 B.n273 585
R299 B.n273 B.n272 585
R300 B.n505 B.n504 585
R301 B.n506 B.n505 585
R302 B.n267 B.n266 585
R303 B.n268 B.n267 585
R304 B.n514 B.n513 585
R305 B.n513 B.n512 585
R306 B.n515 B.n265 585
R307 B.n265 B.n264 585
R308 B.n517 B.n516 585
R309 B.n518 B.n517 585
R310 B.n259 B.n258 585
R311 B.n260 B.n259 585
R312 B.n526 B.n525 585
R313 B.n525 B.n524 585
R314 B.n527 B.n257 585
R315 B.n257 B.n255 585
R316 B.n529 B.n528 585
R317 B.n530 B.n529 585
R318 B.n251 B.n250 585
R319 B.n256 B.n251 585
R320 B.n538 B.n537 585
R321 B.n537 B.n536 585
R322 B.n539 B.n249 585
R323 B.n249 B.n247 585
R324 B.n541 B.n540 585
R325 B.n542 B.n541 585
R326 B.n243 B.n242 585
R327 B.n248 B.n243 585
R328 B.n550 B.n549 585
R329 B.n549 B.n548 585
R330 B.n551 B.n241 585
R331 B.n241 B.n240 585
R332 B.n553 B.n552 585
R333 B.n554 B.n553 585
R334 B.n235 B.n234 585
R335 B.n236 B.n235 585
R336 B.n563 B.n562 585
R337 B.n562 B.n561 585
R338 B.n564 B.n233 585
R339 B.n233 B.n232 585
R340 B.n566 B.n565 585
R341 B.n567 B.n566 585
R342 B.n2 B.n0 585
R343 B.n4 B.n2 585
R344 B.n3 B.n1 585
R345 B.n689 B.n3 585
R346 B.n687 B.n686 585
R347 B.n688 B.n687 585
R348 B.n685 B.n9 585
R349 B.n9 B.n8 585
R350 B.n684 B.n683 585
R351 B.n683 B.n682 585
R352 B.n11 B.n10 585
R353 B.n681 B.n11 585
R354 B.n679 B.n678 585
R355 B.n680 B.n679 585
R356 B.n677 B.n16 585
R357 B.n16 B.n15 585
R358 B.n676 B.n675 585
R359 B.n675 B.n674 585
R360 B.n18 B.n17 585
R361 B.n673 B.n18 585
R362 B.n671 B.n670 585
R363 B.n672 B.n671 585
R364 B.n669 B.n23 585
R365 B.n23 B.n22 585
R366 B.n668 B.n667 585
R367 B.n667 B.n666 585
R368 B.n25 B.n24 585
R369 B.n665 B.n25 585
R370 B.n663 B.n662 585
R371 B.n664 B.n663 585
R372 B.n661 B.n30 585
R373 B.n30 B.n29 585
R374 B.n660 B.n659 585
R375 B.n659 B.n658 585
R376 B.n32 B.n31 585
R377 B.n657 B.n32 585
R378 B.n655 B.n654 585
R379 B.n656 B.n655 585
R380 B.n653 B.n37 585
R381 B.n37 B.n36 585
R382 B.n652 B.n651 585
R383 B.n651 B.n650 585
R384 B.n39 B.n38 585
R385 B.n649 B.n39 585
R386 B.n647 B.n646 585
R387 B.n648 B.n647 585
R388 B.n645 B.n44 585
R389 B.n44 B.n43 585
R390 B.n644 B.n643 585
R391 B.n643 B.n642 585
R392 B.n46 B.n45 585
R393 B.n641 B.n46 585
R394 B.n639 B.n638 585
R395 B.n640 B.n639 585
R396 B.n637 B.n51 585
R397 B.n51 B.n50 585
R398 B.n636 B.n635 585
R399 B.n635 B.n634 585
R400 B.n53 B.n52 585
R401 B.n633 B.n53 585
R402 B.n631 B.n630 585
R403 B.n632 B.n631 585
R404 B.n629 B.n58 585
R405 B.n58 B.n57 585
R406 B.n628 B.n627 585
R407 B.n627 B.n626 585
R408 B.n60 B.n59 585
R409 B.n625 B.n60 585
R410 B.n623 B.n622 585
R411 B.n624 B.n623 585
R412 B.n621 B.n65 585
R413 B.n65 B.n64 585
R414 B.n692 B.n691 585
R415 B.n691 B.n690 585
R416 B.n465 B.n297 463.671
R417 B.n619 B.n65 463.671
R418 B.n337 B.n295 463.671
R419 B.n616 B.n100 463.671
R420 B.n334 B.t10 350.286
R421 B.n332 B.t18 350.286
R422 B.n103 B.t21 350.286
R423 B.n101 B.t14 350.286
R424 B.n617 B.n98 256.663
R425 B.n617 B.n97 256.663
R426 B.n617 B.n96 256.663
R427 B.n617 B.n95 256.663
R428 B.n617 B.n94 256.663
R429 B.n617 B.n93 256.663
R430 B.n617 B.n92 256.663
R431 B.n617 B.n91 256.663
R432 B.n617 B.n90 256.663
R433 B.n617 B.n89 256.663
R434 B.n617 B.n88 256.663
R435 B.n617 B.n87 256.663
R436 B.n617 B.n86 256.663
R437 B.n617 B.n85 256.663
R438 B.n617 B.n84 256.663
R439 B.n617 B.n83 256.663
R440 B.n617 B.n82 256.663
R441 B.n617 B.n81 256.663
R442 B.n617 B.n80 256.663
R443 B.n617 B.n79 256.663
R444 B.n617 B.n78 256.663
R445 B.n617 B.n77 256.663
R446 B.n617 B.n76 256.663
R447 B.n617 B.n75 256.663
R448 B.n617 B.n74 256.663
R449 B.n617 B.n73 256.663
R450 B.n617 B.n72 256.663
R451 B.n617 B.n71 256.663
R452 B.n617 B.n70 256.663
R453 B.n617 B.n69 256.663
R454 B.n617 B.n68 256.663
R455 B.n618 B.n617 256.663
R456 B.n464 B.n463 256.663
R457 B.n463 B.n300 256.663
R458 B.n463 B.n301 256.663
R459 B.n463 B.n302 256.663
R460 B.n463 B.n303 256.663
R461 B.n463 B.n304 256.663
R462 B.n463 B.n305 256.663
R463 B.n463 B.n306 256.663
R464 B.n463 B.n307 256.663
R465 B.n463 B.n308 256.663
R466 B.n463 B.n309 256.663
R467 B.n463 B.n310 256.663
R468 B.n463 B.n311 256.663
R469 B.n463 B.n312 256.663
R470 B.n463 B.n313 256.663
R471 B.n463 B.n314 256.663
R472 B.n463 B.n315 256.663
R473 B.n463 B.n316 256.663
R474 B.n463 B.n317 256.663
R475 B.n463 B.n318 256.663
R476 B.n463 B.n319 256.663
R477 B.n463 B.n320 256.663
R478 B.n463 B.n321 256.663
R479 B.n463 B.n322 256.663
R480 B.n463 B.n323 256.663
R481 B.n463 B.n324 256.663
R482 B.n463 B.n325 256.663
R483 B.n463 B.n326 256.663
R484 B.n463 B.n327 256.663
R485 B.n463 B.n328 256.663
R486 B.n463 B.n329 256.663
R487 B.n463 B.n330 256.663
R488 B.n334 B.t13 229.125
R489 B.n101 B.t16 229.125
R490 B.n332 B.t20 229.125
R491 B.n103 B.t22 229.125
R492 B.n335 B.t12 199.647
R493 B.n102 B.t17 199.647
R494 B.n333 B.t19 199.647
R495 B.n104 B.t23 199.647
R496 B.n469 B.n297 163.367
R497 B.n469 B.n291 163.367
R498 B.n477 B.n291 163.367
R499 B.n477 B.n289 163.367
R500 B.n481 B.n289 163.367
R501 B.n481 B.n283 163.367
R502 B.n489 B.n283 163.367
R503 B.n489 B.n281 163.367
R504 B.n493 B.n281 163.367
R505 B.n493 B.n275 163.367
R506 B.n501 B.n275 163.367
R507 B.n501 B.n273 163.367
R508 B.n505 B.n273 163.367
R509 B.n505 B.n267 163.367
R510 B.n513 B.n267 163.367
R511 B.n513 B.n265 163.367
R512 B.n517 B.n265 163.367
R513 B.n517 B.n259 163.367
R514 B.n525 B.n259 163.367
R515 B.n525 B.n257 163.367
R516 B.n529 B.n257 163.367
R517 B.n529 B.n251 163.367
R518 B.n537 B.n251 163.367
R519 B.n537 B.n249 163.367
R520 B.n541 B.n249 163.367
R521 B.n541 B.n243 163.367
R522 B.n549 B.n243 163.367
R523 B.n549 B.n241 163.367
R524 B.n553 B.n241 163.367
R525 B.n553 B.n235 163.367
R526 B.n562 B.n235 163.367
R527 B.n562 B.n233 163.367
R528 B.n566 B.n233 163.367
R529 B.n566 B.n2 163.367
R530 B.n691 B.n2 163.367
R531 B.n691 B.n3 163.367
R532 B.n687 B.n3 163.367
R533 B.n687 B.n9 163.367
R534 B.n683 B.n9 163.367
R535 B.n683 B.n11 163.367
R536 B.n679 B.n11 163.367
R537 B.n679 B.n16 163.367
R538 B.n675 B.n16 163.367
R539 B.n675 B.n18 163.367
R540 B.n671 B.n18 163.367
R541 B.n671 B.n23 163.367
R542 B.n667 B.n23 163.367
R543 B.n667 B.n25 163.367
R544 B.n663 B.n25 163.367
R545 B.n663 B.n30 163.367
R546 B.n659 B.n30 163.367
R547 B.n659 B.n32 163.367
R548 B.n655 B.n32 163.367
R549 B.n655 B.n37 163.367
R550 B.n651 B.n37 163.367
R551 B.n651 B.n39 163.367
R552 B.n647 B.n39 163.367
R553 B.n647 B.n44 163.367
R554 B.n643 B.n44 163.367
R555 B.n643 B.n46 163.367
R556 B.n639 B.n46 163.367
R557 B.n639 B.n51 163.367
R558 B.n635 B.n51 163.367
R559 B.n635 B.n53 163.367
R560 B.n631 B.n53 163.367
R561 B.n631 B.n58 163.367
R562 B.n627 B.n58 163.367
R563 B.n627 B.n60 163.367
R564 B.n623 B.n60 163.367
R565 B.n623 B.n65 163.367
R566 B.n462 B.n299 163.367
R567 B.n462 B.n331 163.367
R568 B.n458 B.n457 163.367
R569 B.n454 B.n453 163.367
R570 B.n450 B.n449 163.367
R571 B.n446 B.n445 163.367
R572 B.n442 B.n441 163.367
R573 B.n438 B.n437 163.367
R574 B.n434 B.n433 163.367
R575 B.n430 B.n429 163.367
R576 B.n426 B.n425 163.367
R577 B.n422 B.n421 163.367
R578 B.n418 B.n417 163.367
R579 B.n414 B.n413 163.367
R580 B.n409 B.n408 163.367
R581 B.n405 B.n404 163.367
R582 B.n401 B.n400 163.367
R583 B.n397 B.n396 163.367
R584 B.n393 B.n392 163.367
R585 B.n389 B.n388 163.367
R586 B.n385 B.n384 163.367
R587 B.n381 B.n380 163.367
R588 B.n377 B.n376 163.367
R589 B.n373 B.n372 163.367
R590 B.n369 B.n368 163.367
R591 B.n365 B.n364 163.367
R592 B.n361 B.n360 163.367
R593 B.n357 B.n356 163.367
R594 B.n353 B.n352 163.367
R595 B.n349 B.n348 163.367
R596 B.n345 B.n344 163.367
R597 B.n341 B.n340 163.367
R598 B.n471 B.n295 163.367
R599 B.n471 B.n293 163.367
R600 B.n475 B.n293 163.367
R601 B.n475 B.n287 163.367
R602 B.n483 B.n287 163.367
R603 B.n483 B.n285 163.367
R604 B.n487 B.n285 163.367
R605 B.n487 B.n279 163.367
R606 B.n495 B.n279 163.367
R607 B.n495 B.n277 163.367
R608 B.n499 B.n277 163.367
R609 B.n499 B.n271 163.367
R610 B.n507 B.n271 163.367
R611 B.n507 B.n269 163.367
R612 B.n511 B.n269 163.367
R613 B.n511 B.n263 163.367
R614 B.n519 B.n263 163.367
R615 B.n519 B.n261 163.367
R616 B.n523 B.n261 163.367
R617 B.n523 B.n254 163.367
R618 B.n531 B.n254 163.367
R619 B.n531 B.n252 163.367
R620 B.n535 B.n252 163.367
R621 B.n535 B.n246 163.367
R622 B.n543 B.n246 163.367
R623 B.n543 B.n244 163.367
R624 B.n547 B.n244 163.367
R625 B.n547 B.n239 163.367
R626 B.n555 B.n239 163.367
R627 B.n555 B.n237 163.367
R628 B.n560 B.n237 163.367
R629 B.n560 B.n231 163.367
R630 B.n568 B.n231 163.367
R631 B.n569 B.n568 163.367
R632 B.n569 B.n5 163.367
R633 B.n6 B.n5 163.367
R634 B.n7 B.n6 163.367
R635 B.n574 B.n7 163.367
R636 B.n574 B.n12 163.367
R637 B.n13 B.n12 163.367
R638 B.n14 B.n13 163.367
R639 B.n579 B.n14 163.367
R640 B.n579 B.n19 163.367
R641 B.n20 B.n19 163.367
R642 B.n21 B.n20 163.367
R643 B.n584 B.n21 163.367
R644 B.n584 B.n26 163.367
R645 B.n27 B.n26 163.367
R646 B.n28 B.n27 163.367
R647 B.n589 B.n28 163.367
R648 B.n589 B.n33 163.367
R649 B.n34 B.n33 163.367
R650 B.n35 B.n34 163.367
R651 B.n594 B.n35 163.367
R652 B.n594 B.n40 163.367
R653 B.n41 B.n40 163.367
R654 B.n42 B.n41 163.367
R655 B.n599 B.n42 163.367
R656 B.n599 B.n47 163.367
R657 B.n48 B.n47 163.367
R658 B.n49 B.n48 163.367
R659 B.n604 B.n49 163.367
R660 B.n604 B.n54 163.367
R661 B.n55 B.n54 163.367
R662 B.n56 B.n55 163.367
R663 B.n609 B.n56 163.367
R664 B.n609 B.n61 163.367
R665 B.n62 B.n61 163.367
R666 B.n63 B.n62 163.367
R667 B.n100 B.n63 163.367
R668 B.n106 B.n67 163.367
R669 B.n110 B.n109 163.367
R670 B.n114 B.n113 163.367
R671 B.n118 B.n117 163.367
R672 B.n122 B.n121 163.367
R673 B.n126 B.n125 163.367
R674 B.n130 B.n129 163.367
R675 B.n134 B.n133 163.367
R676 B.n138 B.n137 163.367
R677 B.n142 B.n141 163.367
R678 B.n146 B.n145 163.367
R679 B.n150 B.n149 163.367
R680 B.n154 B.n153 163.367
R681 B.n158 B.n157 163.367
R682 B.n162 B.n161 163.367
R683 B.n166 B.n165 163.367
R684 B.n170 B.n169 163.367
R685 B.n174 B.n173 163.367
R686 B.n179 B.n178 163.367
R687 B.n183 B.n182 163.367
R688 B.n187 B.n186 163.367
R689 B.n191 B.n190 163.367
R690 B.n195 B.n194 163.367
R691 B.n199 B.n198 163.367
R692 B.n203 B.n202 163.367
R693 B.n207 B.n206 163.367
R694 B.n211 B.n210 163.367
R695 B.n215 B.n214 163.367
R696 B.n219 B.n218 163.367
R697 B.n223 B.n222 163.367
R698 B.n227 B.n226 163.367
R699 B.n616 B.n99 163.367
R700 B.n463 B.n296 104.763
R701 B.n617 B.n64 104.763
R702 B.n465 B.n464 71.676
R703 B.n331 B.n300 71.676
R704 B.n457 B.n301 71.676
R705 B.n453 B.n302 71.676
R706 B.n449 B.n303 71.676
R707 B.n445 B.n304 71.676
R708 B.n441 B.n305 71.676
R709 B.n437 B.n306 71.676
R710 B.n433 B.n307 71.676
R711 B.n429 B.n308 71.676
R712 B.n425 B.n309 71.676
R713 B.n421 B.n310 71.676
R714 B.n417 B.n311 71.676
R715 B.n413 B.n312 71.676
R716 B.n408 B.n313 71.676
R717 B.n404 B.n314 71.676
R718 B.n400 B.n315 71.676
R719 B.n396 B.n316 71.676
R720 B.n392 B.n317 71.676
R721 B.n388 B.n318 71.676
R722 B.n384 B.n319 71.676
R723 B.n380 B.n320 71.676
R724 B.n376 B.n321 71.676
R725 B.n372 B.n322 71.676
R726 B.n368 B.n323 71.676
R727 B.n364 B.n324 71.676
R728 B.n360 B.n325 71.676
R729 B.n356 B.n326 71.676
R730 B.n352 B.n327 71.676
R731 B.n348 B.n328 71.676
R732 B.n344 B.n329 71.676
R733 B.n340 B.n330 71.676
R734 B.n619 B.n618 71.676
R735 B.n106 B.n68 71.676
R736 B.n110 B.n69 71.676
R737 B.n114 B.n70 71.676
R738 B.n118 B.n71 71.676
R739 B.n122 B.n72 71.676
R740 B.n126 B.n73 71.676
R741 B.n130 B.n74 71.676
R742 B.n134 B.n75 71.676
R743 B.n138 B.n76 71.676
R744 B.n142 B.n77 71.676
R745 B.n146 B.n78 71.676
R746 B.n150 B.n79 71.676
R747 B.n154 B.n80 71.676
R748 B.n158 B.n81 71.676
R749 B.n162 B.n82 71.676
R750 B.n166 B.n83 71.676
R751 B.n170 B.n84 71.676
R752 B.n174 B.n85 71.676
R753 B.n179 B.n86 71.676
R754 B.n183 B.n87 71.676
R755 B.n187 B.n88 71.676
R756 B.n191 B.n89 71.676
R757 B.n195 B.n90 71.676
R758 B.n199 B.n91 71.676
R759 B.n203 B.n92 71.676
R760 B.n207 B.n93 71.676
R761 B.n211 B.n94 71.676
R762 B.n215 B.n95 71.676
R763 B.n219 B.n96 71.676
R764 B.n223 B.n97 71.676
R765 B.n227 B.n98 71.676
R766 B.n99 B.n98 71.676
R767 B.n226 B.n97 71.676
R768 B.n222 B.n96 71.676
R769 B.n218 B.n95 71.676
R770 B.n214 B.n94 71.676
R771 B.n210 B.n93 71.676
R772 B.n206 B.n92 71.676
R773 B.n202 B.n91 71.676
R774 B.n198 B.n90 71.676
R775 B.n194 B.n89 71.676
R776 B.n190 B.n88 71.676
R777 B.n186 B.n87 71.676
R778 B.n182 B.n86 71.676
R779 B.n178 B.n85 71.676
R780 B.n173 B.n84 71.676
R781 B.n169 B.n83 71.676
R782 B.n165 B.n82 71.676
R783 B.n161 B.n81 71.676
R784 B.n157 B.n80 71.676
R785 B.n153 B.n79 71.676
R786 B.n149 B.n78 71.676
R787 B.n145 B.n77 71.676
R788 B.n141 B.n76 71.676
R789 B.n137 B.n75 71.676
R790 B.n133 B.n74 71.676
R791 B.n129 B.n73 71.676
R792 B.n125 B.n72 71.676
R793 B.n121 B.n71 71.676
R794 B.n117 B.n70 71.676
R795 B.n113 B.n69 71.676
R796 B.n109 B.n68 71.676
R797 B.n618 B.n67 71.676
R798 B.n464 B.n299 71.676
R799 B.n458 B.n300 71.676
R800 B.n454 B.n301 71.676
R801 B.n450 B.n302 71.676
R802 B.n446 B.n303 71.676
R803 B.n442 B.n304 71.676
R804 B.n438 B.n305 71.676
R805 B.n434 B.n306 71.676
R806 B.n430 B.n307 71.676
R807 B.n426 B.n308 71.676
R808 B.n422 B.n309 71.676
R809 B.n418 B.n310 71.676
R810 B.n414 B.n311 71.676
R811 B.n409 B.n312 71.676
R812 B.n405 B.n313 71.676
R813 B.n401 B.n314 71.676
R814 B.n397 B.n315 71.676
R815 B.n393 B.n316 71.676
R816 B.n389 B.n317 71.676
R817 B.n385 B.n318 71.676
R818 B.n381 B.n319 71.676
R819 B.n377 B.n320 71.676
R820 B.n373 B.n321 71.676
R821 B.n369 B.n322 71.676
R822 B.n365 B.n323 71.676
R823 B.n361 B.n324 71.676
R824 B.n357 B.n325 71.676
R825 B.n353 B.n326 71.676
R826 B.n349 B.n327 71.676
R827 B.n345 B.n328 71.676
R828 B.n341 B.n329 71.676
R829 B.n337 B.n330 71.676
R830 B.n470 B.n296 59.8644
R831 B.n470 B.n292 59.8644
R832 B.n476 B.n292 59.8644
R833 B.n476 B.n288 59.8644
R834 B.n482 B.n288 59.8644
R835 B.n488 B.n284 59.8644
R836 B.n488 B.n280 59.8644
R837 B.n494 B.n280 59.8644
R838 B.n494 B.n276 59.8644
R839 B.n500 B.n276 59.8644
R840 B.n500 B.n272 59.8644
R841 B.n506 B.n272 59.8644
R842 B.n512 B.n268 59.8644
R843 B.n512 B.n264 59.8644
R844 B.n518 B.n264 59.8644
R845 B.n524 B.n260 59.8644
R846 B.n524 B.n255 59.8644
R847 B.n530 B.n255 59.8644
R848 B.n530 B.n256 59.8644
R849 B.n536 B.n247 59.8644
R850 B.n542 B.n247 59.8644
R851 B.n542 B.n248 59.8644
R852 B.n548 B.n240 59.8644
R853 B.n554 B.n240 59.8644
R854 B.n554 B.n236 59.8644
R855 B.n561 B.n236 59.8644
R856 B.n567 B.n232 59.8644
R857 B.n567 B.n4 59.8644
R858 B.n690 B.n4 59.8644
R859 B.n690 B.n689 59.8644
R860 B.n689 B.n688 59.8644
R861 B.n688 B.n8 59.8644
R862 B.n682 B.n681 59.8644
R863 B.n681 B.n680 59.8644
R864 B.n680 B.n15 59.8644
R865 B.n674 B.n15 59.8644
R866 B.n673 B.n672 59.8644
R867 B.n672 B.n22 59.8644
R868 B.n666 B.n22 59.8644
R869 B.n665 B.n664 59.8644
R870 B.n664 B.n29 59.8644
R871 B.n658 B.n29 59.8644
R872 B.n658 B.n657 59.8644
R873 B.n656 B.n36 59.8644
R874 B.n650 B.n36 59.8644
R875 B.n650 B.n649 59.8644
R876 B.n648 B.n43 59.8644
R877 B.n642 B.n43 59.8644
R878 B.n642 B.n641 59.8644
R879 B.n641 B.n640 59.8644
R880 B.n640 B.n50 59.8644
R881 B.n634 B.n50 59.8644
R882 B.n634 B.n633 59.8644
R883 B.n632 B.n57 59.8644
R884 B.n626 B.n57 59.8644
R885 B.n626 B.n625 59.8644
R886 B.n625 B.n624 59.8644
R887 B.n624 B.n64 59.8644
R888 B.n336 B.n335 59.5399
R889 B.n411 B.n333 59.5399
R890 B.n105 B.n104 59.5399
R891 B.n176 B.n102 59.5399
R892 B.t7 B.n232 50.1806
R893 B.t6 B.n8 50.1806
R894 B.n536 B.t5 46.6592
R895 B.n666 B.t8 46.6592
R896 B.n518 B.t4 44.8985
R897 B.t2 B.n656 44.8985
R898 B.t0 B.n268 43.1378
R899 B.n649 B.t3 43.1378
R900 B.n248 B.t1 41.3771
R901 B.t9 B.n673 41.3771
R902 B.n482 B.t11 36.0949
R903 B.t15 B.n632 36.0949
R904 B.n621 B.n620 30.1273
R905 B.n615 B.n614 30.1273
R906 B.n338 B.n294 30.1273
R907 B.n467 B.n466 30.1273
R908 B.n335 B.n334 29.4793
R909 B.n333 B.n332 29.4793
R910 B.n104 B.n103 29.4793
R911 B.n102 B.n101 29.4793
R912 B.t11 B.n284 23.77
R913 B.n633 B.t15 23.77
R914 B.n548 B.t1 18.4879
R915 B.n674 B.t9 18.4879
R916 B B.n692 18.0485
R917 B.n506 B.t0 16.7272
R918 B.t3 B.n648 16.7272
R919 B.t4 B.n260 14.9665
R920 B.n657 B.t2 14.9665
R921 B.n256 B.t5 13.2058
R922 B.t8 B.n665 13.2058
R923 B.n620 B.n66 10.6151
R924 B.n107 B.n66 10.6151
R925 B.n108 B.n107 10.6151
R926 B.n111 B.n108 10.6151
R927 B.n112 B.n111 10.6151
R928 B.n115 B.n112 10.6151
R929 B.n116 B.n115 10.6151
R930 B.n119 B.n116 10.6151
R931 B.n120 B.n119 10.6151
R932 B.n123 B.n120 10.6151
R933 B.n124 B.n123 10.6151
R934 B.n127 B.n124 10.6151
R935 B.n128 B.n127 10.6151
R936 B.n131 B.n128 10.6151
R937 B.n132 B.n131 10.6151
R938 B.n135 B.n132 10.6151
R939 B.n136 B.n135 10.6151
R940 B.n139 B.n136 10.6151
R941 B.n140 B.n139 10.6151
R942 B.n143 B.n140 10.6151
R943 B.n144 B.n143 10.6151
R944 B.n147 B.n144 10.6151
R945 B.n148 B.n147 10.6151
R946 B.n151 B.n148 10.6151
R947 B.n152 B.n151 10.6151
R948 B.n155 B.n152 10.6151
R949 B.n156 B.n155 10.6151
R950 B.n160 B.n159 10.6151
R951 B.n163 B.n160 10.6151
R952 B.n164 B.n163 10.6151
R953 B.n167 B.n164 10.6151
R954 B.n168 B.n167 10.6151
R955 B.n171 B.n168 10.6151
R956 B.n172 B.n171 10.6151
R957 B.n175 B.n172 10.6151
R958 B.n180 B.n177 10.6151
R959 B.n181 B.n180 10.6151
R960 B.n184 B.n181 10.6151
R961 B.n185 B.n184 10.6151
R962 B.n188 B.n185 10.6151
R963 B.n189 B.n188 10.6151
R964 B.n192 B.n189 10.6151
R965 B.n193 B.n192 10.6151
R966 B.n196 B.n193 10.6151
R967 B.n197 B.n196 10.6151
R968 B.n200 B.n197 10.6151
R969 B.n201 B.n200 10.6151
R970 B.n204 B.n201 10.6151
R971 B.n205 B.n204 10.6151
R972 B.n208 B.n205 10.6151
R973 B.n209 B.n208 10.6151
R974 B.n212 B.n209 10.6151
R975 B.n213 B.n212 10.6151
R976 B.n216 B.n213 10.6151
R977 B.n217 B.n216 10.6151
R978 B.n220 B.n217 10.6151
R979 B.n221 B.n220 10.6151
R980 B.n224 B.n221 10.6151
R981 B.n225 B.n224 10.6151
R982 B.n228 B.n225 10.6151
R983 B.n229 B.n228 10.6151
R984 B.n615 B.n229 10.6151
R985 B.n472 B.n294 10.6151
R986 B.n473 B.n472 10.6151
R987 B.n474 B.n473 10.6151
R988 B.n474 B.n286 10.6151
R989 B.n484 B.n286 10.6151
R990 B.n485 B.n484 10.6151
R991 B.n486 B.n485 10.6151
R992 B.n486 B.n278 10.6151
R993 B.n496 B.n278 10.6151
R994 B.n497 B.n496 10.6151
R995 B.n498 B.n497 10.6151
R996 B.n498 B.n270 10.6151
R997 B.n508 B.n270 10.6151
R998 B.n509 B.n508 10.6151
R999 B.n510 B.n509 10.6151
R1000 B.n510 B.n262 10.6151
R1001 B.n520 B.n262 10.6151
R1002 B.n521 B.n520 10.6151
R1003 B.n522 B.n521 10.6151
R1004 B.n522 B.n253 10.6151
R1005 B.n532 B.n253 10.6151
R1006 B.n533 B.n532 10.6151
R1007 B.n534 B.n533 10.6151
R1008 B.n534 B.n245 10.6151
R1009 B.n544 B.n245 10.6151
R1010 B.n545 B.n544 10.6151
R1011 B.n546 B.n545 10.6151
R1012 B.n546 B.n238 10.6151
R1013 B.n556 B.n238 10.6151
R1014 B.n557 B.n556 10.6151
R1015 B.n559 B.n557 10.6151
R1016 B.n559 B.n558 10.6151
R1017 B.n558 B.n230 10.6151
R1018 B.n570 B.n230 10.6151
R1019 B.n571 B.n570 10.6151
R1020 B.n572 B.n571 10.6151
R1021 B.n573 B.n572 10.6151
R1022 B.n575 B.n573 10.6151
R1023 B.n576 B.n575 10.6151
R1024 B.n577 B.n576 10.6151
R1025 B.n578 B.n577 10.6151
R1026 B.n580 B.n578 10.6151
R1027 B.n581 B.n580 10.6151
R1028 B.n582 B.n581 10.6151
R1029 B.n583 B.n582 10.6151
R1030 B.n585 B.n583 10.6151
R1031 B.n586 B.n585 10.6151
R1032 B.n587 B.n586 10.6151
R1033 B.n588 B.n587 10.6151
R1034 B.n590 B.n588 10.6151
R1035 B.n591 B.n590 10.6151
R1036 B.n592 B.n591 10.6151
R1037 B.n593 B.n592 10.6151
R1038 B.n595 B.n593 10.6151
R1039 B.n596 B.n595 10.6151
R1040 B.n597 B.n596 10.6151
R1041 B.n598 B.n597 10.6151
R1042 B.n600 B.n598 10.6151
R1043 B.n601 B.n600 10.6151
R1044 B.n602 B.n601 10.6151
R1045 B.n603 B.n602 10.6151
R1046 B.n605 B.n603 10.6151
R1047 B.n606 B.n605 10.6151
R1048 B.n607 B.n606 10.6151
R1049 B.n608 B.n607 10.6151
R1050 B.n610 B.n608 10.6151
R1051 B.n611 B.n610 10.6151
R1052 B.n612 B.n611 10.6151
R1053 B.n613 B.n612 10.6151
R1054 B.n614 B.n613 10.6151
R1055 B.n466 B.n298 10.6151
R1056 B.n461 B.n298 10.6151
R1057 B.n461 B.n460 10.6151
R1058 B.n460 B.n459 10.6151
R1059 B.n459 B.n456 10.6151
R1060 B.n456 B.n455 10.6151
R1061 B.n455 B.n452 10.6151
R1062 B.n452 B.n451 10.6151
R1063 B.n451 B.n448 10.6151
R1064 B.n448 B.n447 10.6151
R1065 B.n447 B.n444 10.6151
R1066 B.n444 B.n443 10.6151
R1067 B.n443 B.n440 10.6151
R1068 B.n440 B.n439 10.6151
R1069 B.n439 B.n436 10.6151
R1070 B.n436 B.n435 10.6151
R1071 B.n435 B.n432 10.6151
R1072 B.n432 B.n431 10.6151
R1073 B.n431 B.n428 10.6151
R1074 B.n428 B.n427 10.6151
R1075 B.n427 B.n424 10.6151
R1076 B.n424 B.n423 10.6151
R1077 B.n423 B.n420 10.6151
R1078 B.n420 B.n419 10.6151
R1079 B.n419 B.n416 10.6151
R1080 B.n416 B.n415 10.6151
R1081 B.n415 B.n412 10.6151
R1082 B.n410 B.n407 10.6151
R1083 B.n407 B.n406 10.6151
R1084 B.n406 B.n403 10.6151
R1085 B.n403 B.n402 10.6151
R1086 B.n402 B.n399 10.6151
R1087 B.n399 B.n398 10.6151
R1088 B.n398 B.n395 10.6151
R1089 B.n395 B.n394 10.6151
R1090 B.n391 B.n390 10.6151
R1091 B.n390 B.n387 10.6151
R1092 B.n387 B.n386 10.6151
R1093 B.n386 B.n383 10.6151
R1094 B.n383 B.n382 10.6151
R1095 B.n382 B.n379 10.6151
R1096 B.n379 B.n378 10.6151
R1097 B.n378 B.n375 10.6151
R1098 B.n375 B.n374 10.6151
R1099 B.n374 B.n371 10.6151
R1100 B.n371 B.n370 10.6151
R1101 B.n370 B.n367 10.6151
R1102 B.n367 B.n366 10.6151
R1103 B.n366 B.n363 10.6151
R1104 B.n363 B.n362 10.6151
R1105 B.n362 B.n359 10.6151
R1106 B.n359 B.n358 10.6151
R1107 B.n358 B.n355 10.6151
R1108 B.n355 B.n354 10.6151
R1109 B.n354 B.n351 10.6151
R1110 B.n351 B.n350 10.6151
R1111 B.n350 B.n347 10.6151
R1112 B.n347 B.n346 10.6151
R1113 B.n346 B.n343 10.6151
R1114 B.n343 B.n342 10.6151
R1115 B.n342 B.n339 10.6151
R1116 B.n339 B.n338 10.6151
R1117 B.n468 B.n467 10.6151
R1118 B.n468 B.n290 10.6151
R1119 B.n478 B.n290 10.6151
R1120 B.n479 B.n478 10.6151
R1121 B.n480 B.n479 10.6151
R1122 B.n480 B.n282 10.6151
R1123 B.n490 B.n282 10.6151
R1124 B.n491 B.n490 10.6151
R1125 B.n492 B.n491 10.6151
R1126 B.n492 B.n274 10.6151
R1127 B.n502 B.n274 10.6151
R1128 B.n503 B.n502 10.6151
R1129 B.n504 B.n503 10.6151
R1130 B.n504 B.n266 10.6151
R1131 B.n514 B.n266 10.6151
R1132 B.n515 B.n514 10.6151
R1133 B.n516 B.n515 10.6151
R1134 B.n516 B.n258 10.6151
R1135 B.n526 B.n258 10.6151
R1136 B.n527 B.n526 10.6151
R1137 B.n528 B.n527 10.6151
R1138 B.n528 B.n250 10.6151
R1139 B.n538 B.n250 10.6151
R1140 B.n539 B.n538 10.6151
R1141 B.n540 B.n539 10.6151
R1142 B.n540 B.n242 10.6151
R1143 B.n550 B.n242 10.6151
R1144 B.n551 B.n550 10.6151
R1145 B.n552 B.n551 10.6151
R1146 B.n552 B.n234 10.6151
R1147 B.n563 B.n234 10.6151
R1148 B.n564 B.n563 10.6151
R1149 B.n565 B.n564 10.6151
R1150 B.n565 B.n0 10.6151
R1151 B.n686 B.n1 10.6151
R1152 B.n686 B.n685 10.6151
R1153 B.n685 B.n684 10.6151
R1154 B.n684 B.n10 10.6151
R1155 B.n678 B.n10 10.6151
R1156 B.n678 B.n677 10.6151
R1157 B.n677 B.n676 10.6151
R1158 B.n676 B.n17 10.6151
R1159 B.n670 B.n17 10.6151
R1160 B.n670 B.n669 10.6151
R1161 B.n669 B.n668 10.6151
R1162 B.n668 B.n24 10.6151
R1163 B.n662 B.n24 10.6151
R1164 B.n662 B.n661 10.6151
R1165 B.n661 B.n660 10.6151
R1166 B.n660 B.n31 10.6151
R1167 B.n654 B.n31 10.6151
R1168 B.n654 B.n653 10.6151
R1169 B.n653 B.n652 10.6151
R1170 B.n652 B.n38 10.6151
R1171 B.n646 B.n38 10.6151
R1172 B.n646 B.n645 10.6151
R1173 B.n645 B.n644 10.6151
R1174 B.n644 B.n45 10.6151
R1175 B.n638 B.n45 10.6151
R1176 B.n638 B.n637 10.6151
R1177 B.n637 B.n636 10.6151
R1178 B.n636 B.n52 10.6151
R1179 B.n630 B.n52 10.6151
R1180 B.n630 B.n629 10.6151
R1181 B.n629 B.n628 10.6151
R1182 B.n628 B.n59 10.6151
R1183 B.n622 B.n59 10.6151
R1184 B.n622 B.n621 10.6151
R1185 B.n561 B.t7 9.68437
R1186 B.n682 B.t6 9.68437
R1187 B.n159 B.n105 6.5566
R1188 B.n176 B.n175 6.5566
R1189 B.n411 B.n410 6.5566
R1190 B.n394 B.n336 6.5566
R1191 B.n156 B.n105 4.05904
R1192 B.n177 B.n176 4.05904
R1193 B.n412 B.n411 4.05904
R1194 B.n391 B.n336 4.05904
R1195 B.n692 B.n0 2.81026
R1196 B.n692 B.n1 2.81026
R1197 VN.n6 VN.t0 197.749
R1198 VN.n28 VN.t6 197.749
R1199 VN.n20 VN.t7 179.232
R1200 VN.n42 VN.t9 179.232
R1201 VN.n41 VN.n22 161.3
R1202 VN.n40 VN.n39 161.3
R1203 VN.n38 VN.n37 161.3
R1204 VN.n36 VN.n24 161.3
R1205 VN.n35 VN.n34 161.3
R1206 VN.n33 VN.n32 161.3
R1207 VN.n31 VN.n26 161.3
R1208 VN.n30 VN.n29 161.3
R1209 VN.n19 VN.n0 161.3
R1210 VN.n18 VN.n17 161.3
R1211 VN.n16 VN.n15 161.3
R1212 VN.n14 VN.n2 161.3
R1213 VN.n13 VN.n12 161.3
R1214 VN.n11 VN.n10 161.3
R1215 VN.n9 VN.n4 161.3
R1216 VN.n8 VN.n7 161.3
R1217 VN.n5 VN.t4 146.22
R1218 VN.n3 VN.t8 146.22
R1219 VN.n1 VN.t2 146.22
R1220 VN.n27 VN.t5 146.22
R1221 VN.n25 VN.t3 146.22
R1222 VN.n23 VN.t1 146.22
R1223 VN.n43 VN.n42 80.6037
R1224 VN.n21 VN.n20 80.6037
R1225 VN.n6 VN.n5 44.6572
R1226 VN.n28 VN.n27 44.6572
R1227 VN VN.n43 42.2187
R1228 VN.n9 VN.n8 41.5458
R1229 VN.n15 VN.n14 41.5458
R1230 VN.n31 VN.n30 41.5458
R1231 VN.n37 VN.n36 41.5458
R1232 VN.n10 VN.n9 39.6083
R1233 VN.n14 VN.n13 39.6083
R1234 VN.n32 VN.n31 39.6083
R1235 VN.n36 VN.n35 39.6083
R1236 VN.n19 VN.n18 37.6707
R1237 VN.n41 VN.n40 37.6707
R1238 VN.n29 VN.n28 29.7202
R1239 VN.n7 VN.n6 29.7202
R1240 VN.n20 VN.n19 28.4823
R1241 VN.n42 VN.n41 28.4823
R1242 VN.n8 VN.n5 13.2801
R1243 VN.n15 VN.n1 13.2801
R1244 VN.n30 VN.n27 13.2801
R1245 VN.n37 VN.n23 13.2801
R1246 VN.n10 VN.n3 12.2964
R1247 VN.n13 VN.n3 12.2964
R1248 VN.n35 VN.n25 12.2964
R1249 VN.n32 VN.n25 12.2964
R1250 VN.n18 VN.n1 11.3127
R1251 VN.n40 VN.n23 11.3127
R1252 VN.n43 VN.n22 0.285035
R1253 VN.n21 VN.n0 0.285035
R1254 VN.n39 VN.n22 0.189894
R1255 VN.n39 VN.n38 0.189894
R1256 VN.n38 VN.n24 0.189894
R1257 VN.n34 VN.n24 0.189894
R1258 VN.n34 VN.n33 0.189894
R1259 VN.n33 VN.n26 0.189894
R1260 VN.n29 VN.n26 0.189894
R1261 VN.n7 VN.n4 0.189894
R1262 VN.n11 VN.n4 0.189894
R1263 VN.n12 VN.n11 0.189894
R1264 VN.n12 VN.n2 0.189894
R1265 VN.n16 VN.n2 0.189894
R1266 VN.n17 VN.n16 0.189894
R1267 VN.n17 VN.n0 0.189894
R1268 VN VN.n21 0.146778
R1269 VTAIL.n152 VTAIL.n122 214.453
R1270 VTAIL.n32 VTAIL.n2 214.453
R1271 VTAIL.n116 VTAIL.n86 214.453
R1272 VTAIL.n76 VTAIL.n46 214.453
R1273 VTAIL.n135 VTAIL.n134 185
R1274 VTAIL.n137 VTAIL.n136 185
R1275 VTAIL.n130 VTAIL.n129 185
R1276 VTAIL.n143 VTAIL.n142 185
R1277 VTAIL.n145 VTAIL.n144 185
R1278 VTAIL.n126 VTAIL.n125 185
R1279 VTAIL.n151 VTAIL.n150 185
R1280 VTAIL.n153 VTAIL.n152 185
R1281 VTAIL.n15 VTAIL.n14 185
R1282 VTAIL.n17 VTAIL.n16 185
R1283 VTAIL.n10 VTAIL.n9 185
R1284 VTAIL.n23 VTAIL.n22 185
R1285 VTAIL.n25 VTAIL.n24 185
R1286 VTAIL.n6 VTAIL.n5 185
R1287 VTAIL.n31 VTAIL.n30 185
R1288 VTAIL.n33 VTAIL.n32 185
R1289 VTAIL.n117 VTAIL.n116 185
R1290 VTAIL.n115 VTAIL.n114 185
R1291 VTAIL.n90 VTAIL.n89 185
R1292 VTAIL.n109 VTAIL.n108 185
R1293 VTAIL.n107 VTAIL.n106 185
R1294 VTAIL.n94 VTAIL.n93 185
R1295 VTAIL.n101 VTAIL.n100 185
R1296 VTAIL.n99 VTAIL.n98 185
R1297 VTAIL.n77 VTAIL.n76 185
R1298 VTAIL.n75 VTAIL.n74 185
R1299 VTAIL.n50 VTAIL.n49 185
R1300 VTAIL.n69 VTAIL.n68 185
R1301 VTAIL.n67 VTAIL.n66 185
R1302 VTAIL.n54 VTAIL.n53 185
R1303 VTAIL.n61 VTAIL.n60 185
R1304 VTAIL.n59 VTAIL.n58 185
R1305 VTAIL.n133 VTAIL.t19 149.524
R1306 VTAIL.n13 VTAIL.t3 149.524
R1307 VTAIL.n97 VTAIL.t8 149.524
R1308 VTAIL.n57 VTAIL.t12 149.524
R1309 VTAIL.n136 VTAIL.n135 104.615
R1310 VTAIL.n136 VTAIL.n129 104.615
R1311 VTAIL.n143 VTAIL.n129 104.615
R1312 VTAIL.n144 VTAIL.n143 104.615
R1313 VTAIL.n144 VTAIL.n125 104.615
R1314 VTAIL.n151 VTAIL.n125 104.615
R1315 VTAIL.n152 VTAIL.n151 104.615
R1316 VTAIL.n16 VTAIL.n15 104.615
R1317 VTAIL.n16 VTAIL.n9 104.615
R1318 VTAIL.n23 VTAIL.n9 104.615
R1319 VTAIL.n24 VTAIL.n23 104.615
R1320 VTAIL.n24 VTAIL.n5 104.615
R1321 VTAIL.n31 VTAIL.n5 104.615
R1322 VTAIL.n32 VTAIL.n31 104.615
R1323 VTAIL.n116 VTAIL.n115 104.615
R1324 VTAIL.n115 VTAIL.n89 104.615
R1325 VTAIL.n108 VTAIL.n89 104.615
R1326 VTAIL.n108 VTAIL.n107 104.615
R1327 VTAIL.n107 VTAIL.n93 104.615
R1328 VTAIL.n100 VTAIL.n93 104.615
R1329 VTAIL.n100 VTAIL.n99 104.615
R1330 VTAIL.n76 VTAIL.n75 104.615
R1331 VTAIL.n75 VTAIL.n49 104.615
R1332 VTAIL.n68 VTAIL.n49 104.615
R1333 VTAIL.n68 VTAIL.n67 104.615
R1334 VTAIL.n67 VTAIL.n53 104.615
R1335 VTAIL.n60 VTAIL.n53 104.615
R1336 VTAIL.n60 VTAIL.n59 104.615
R1337 VTAIL.n135 VTAIL.t19 52.3082
R1338 VTAIL.n15 VTAIL.t3 52.3082
R1339 VTAIL.n99 VTAIL.t8 52.3082
R1340 VTAIL.n59 VTAIL.t12 52.3082
R1341 VTAIL.n85 VTAIL.n84 50.6713
R1342 VTAIL.n83 VTAIL.n82 50.6713
R1343 VTAIL.n45 VTAIL.n44 50.6713
R1344 VTAIL.n43 VTAIL.n42 50.6713
R1345 VTAIL.n159 VTAIL.n158 50.6712
R1346 VTAIL.n1 VTAIL.n0 50.6712
R1347 VTAIL.n39 VTAIL.n38 50.6712
R1348 VTAIL.n41 VTAIL.n40 50.6712
R1349 VTAIL.n157 VTAIL.n156 34.9005
R1350 VTAIL.n37 VTAIL.n36 34.9005
R1351 VTAIL.n121 VTAIL.n120 34.9005
R1352 VTAIL.n81 VTAIL.n80 34.9005
R1353 VTAIL.n43 VTAIL.n41 21.2117
R1354 VTAIL.n157 VTAIL.n121 19.9014
R1355 VTAIL.n154 VTAIL.n153 12.8005
R1356 VTAIL.n34 VTAIL.n33 12.8005
R1357 VTAIL.n118 VTAIL.n117 12.8005
R1358 VTAIL.n78 VTAIL.n77 12.8005
R1359 VTAIL.n150 VTAIL.n124 12.0247
R1360 VTAIL.n30 VTAIL.n4 12.0247
R1361 VTAIL.n114 VTAIL.n88 12.0247
R1362 VTAIL.n74 VTAIL.n48 12.0247
R1363 VTAIL.n149 VTAIL.n126 11.249
R1364 VTAIL.n29 VTAIL.n6 11.249
R1365 VTAIL.n113 VTAIL.n90 11.249
R1366 VTAIL.n73 VTAIL.n50 11.249
R1367 VTAIL.n146 VTAIL.n145 10.4732
R1368 VTAIL.n26 VTAIL.n25 10.4732
R1369 VTAIL.n110 VTAIL.n109 10.4732
R1370 VTAIL.n70 VTAIL.n69 10.4732
R1371 VTAIL.n134 VTAIL.n133 10.2747
R1372 VTAIL.n14 VTAIL.n13 10.2747
R1373 VTAIL.n98 VTAIL.n97 10.2747
R1374 VTAIL.n58 VTAIL.n57 10.2747
R1375 VTAIL.n142 VTAIL.n128 9.69747
R1376 VTAIL.n22 VTAIL.n8 9.69747
R1377 VTAIL.n106 VTAIL.n92 9.69747
R1378 VTAIL.n66 VTAIL.n52 9.69747
R1379 VTAIL.n156 VTAIL.n155 9.45567
R1380 VTAIL.n36 VTAIL.n35 9.45567
R1381 VTAIL.n120 VTAIL.n119 9.45567
R1382 VTAIL.n80 VTAIL.n79 9.45567
R1383 VTAIL.n132 VTAIL.n131 9.3005
R1384 VTAIL.n139 VTAIL.n138 9.3005
R1385 VTAIL.n141 VTAIL.n140 9.3005
R1386 VTAIL.n128 VTAIL.n127 9.3005
R1387 VTAIL.n147 VTAIL.n146 9.3005
R1388 VTAIL.n149 VTAIL.n148 9.3005
R1389 VTAIL.n124 VTAIL.n123 9.3005
R1390 VTAIL.n155 VTAIL.n154 9.3005
R1391 VTAIL.n12 VTAIL.n11 9.3005
R1392 VTAIL.n19 VTAIL.n18 9.3005
R1393 VTAIL.n21 VTAIL.n20 9.3005
R1394 VTAIL.n8 VTAIL.n7 9.3005
R1395 VTAIL.n27 VTAIL.n26 9.3005
R1396 VTAIL.n29 VTAIL.n28 9.3005
R1397 VTAIL.n4 VTAIL.n3 9.3005
R1398 VTAIL.n35 VTAIL.n34 9.3005
R1399 VTAIL.n96 VTAIL.n95 9.3005
R1400 VTAIL.n103 VTAIL.n102 9.3005
R1401 VTAIL.n105 VTAIL.n104 9.3005
R1402 VTAIL.n92 VTAIL.n91 9.3005
R1403 VTAIL.n111 VTAIL.n110 9.3005
R1404 VTAIL.n113 VTAIL.n112 9.3005
R1405 VTAIL.n88 VTAIL.n87 9.3005
R1406 VTAIL.n119 VTAIL.n118 9.3005
R1407 VTAIL.n56 VTAIL.n55 9.3005
R1408 VTAIL.n63 VTAIL.n62 9.3005
R1409 VTAIL.n65 VTAIL.n64 9.3005
R1410 VTAIL.n52 VTAIL.n51 9.3005
R1411 VTAIL.n71 VTAIL.n70 9.3005
R1412 VTAIL.n73 VTAIL.n72 9.3005
R1413 VTAIL.n48 VTAIL.n47 9.3005
R1414 VTAIL.n79 VTAIL.n78 9.3005
R1415 VTAIL.n141 VTAIL.n130 8.92171
R1416 VTAIL.n21 VTAIL.n10 8.92171
R1417 VTAIL.n105 VTAIL.n94 8.92171
R1418 VTAIL.n65 VTAIL.n54 8.92171
R1419 VTAIL.n156 VTAIL.n122 8.2187
R1420 VTAIL.n36 VTAIL.n2 8.2187
R1421 VTAIL.n120 VTAIL.n86 8.2187
R1422 VTAIL.n80 VTAIL.n46 8.2187
R1423 VTAIL.n138 VTAIL.n137 8.14595
R1424 VTAIL.n18 VTAIL.n17 8.14595
R1425 VTAIL.n102 VTAIL.n101 8.14595
R1426 VTAIL.n62 VTAIL.n61 8.14595
R1427 VTAIL.n134 VTAIL.n132 7.3702
R1428 VTAIL.n14 VTAIL.n12 7.3702
R1429 VTAIL.n98 VTAIL.n96 7.3702
R1430 VTAIL.n58 VTAIL.n56 7.3702
R1431 VTAIL.n137 VTAIL.n132 5.81868
R1432 VTAIL.n17 VTAIL.n12 5.81868
R1433 VTAIL.n101 VTAIL.n96 5.81868
R1434 VTAIL.n61 VTAIL.n56 5.81868
R1435 VTAIL.n154 VTAIL.n122 5.3904
R1436 VTAIL.n34 VTAIL.n2 5.3904
R1437 VTAIL.n118 VTAIL.n86 5.3904
R1438 VTAIL.n78 VTAIL.n46 5.3904
R1439 VTAIL.n138 VTAIL.n130 5.04292
R1440 VTAIL.n18 VTAIL.n10 5.04292
R1441 VTAIL.n102 VTAIL.n94 5.04292
R1442 VTAIL.n62 VTAIL.n54 5.04292
R1443 VTAIL.n142 VTAIL.n141 4.26717
R1444 VTAIL.n22 VTAIL.n21 4.26717
R1445 VTAIL.n106 VTAIL.n105 4.26717
R1446 VTAIL.n66 VTAIL.n65 4.26717
R1447 VTAIL.n145 VTAIL.n128 3.49141
R1448 VTAIL.n25 VTAIL.n8 3.49141
R1449 VTAIL.n109 VTAIL.n92 3.49141
R1450 VTAIL.n69 VTAIL.n52 3.49141
R1451 VTAIL.n133 VTAIL.n131 2.84305
R1452 VTAIL.n13 VTAIL.n11 2.84305
R1453 VTAIL.n97 VTAIL.n95 2.84305
R1454 VTAIL.n57 VTAIL.n55 2.84305
R1455 VTAIL.n158 VTAIL.t17 2.74288
R1456 VTAIL.n158 VTAIL.t10 2.74288
R1457 VTAIL.n0 VTAIL.t13 2.74288
R1458 VTAIL.n0 VTAIL.t11 2.74288
R1459 VTAIL.n38 VTAIL.t4 2.74288
R1460 VTAIL.n38 VTAIL.t1 2.74288
R1461 VTAIL.n40 VTAIL.t0 2.74288
R1462 VTAIL.n40 VTAIL.t2 2.74288
R1463 VTAIL.n84 VTAIL.t5 2.74288
R1464 VTAIL.n84 VTAIL.t7 2.74288
R1465 VTAIL.n82 VTAIL.t6 2.74288
R1466 VTAIL.n82 VTAIL.t9 2.74288
R1467 VTAIL.n44 VTAIL.t14 2.74288
R1468 VTAIL.n44 VTAIL.t15 2.74288
R1469 VTAIL.n42 VTAIL.t16 2.74288
R1470 VTAIL.n42 VTAIL.t18 2.74288
R1471 VTAIL.n146 VTAIL.n126 2.71565
R1472 VTAIL.n26 VTAIL.n6 2.71565
R1473 VTAIL.n110 VTAIL.n90 2.71565
R1474 VTAIL.n70 VTAIL.n50 2.71565
R1475 VTAIL.n150 VTAIL.n149 1.93989
R1476 VTAIL.n30 VTAIL.n29 1.93989
R1477 VTAIL.n114 VTAIL.n113 1.93989
R1478 VTAIL.n74 VTAIL.n73 1.93989
R1479 VTAIL.n45 VTAIL.n43 1.31084
R1480 VTAIL.n81 VTAIL.n45 1.31084
R1481 VTAIL.n85 VTAIL.n83 1.31084
R1482 VTAIL.n121 VTAIL.n85 1.31084
R1483 VTAIL.n41 VTAIL.n39 1.31084
R1484 VTAIL.n39 VTAIL.n37 1.31084
R1485 VTAIL.n159 VTAIL.n157 1.31084
R1486 VTAIL.n153 VTAIL.n124 1.16414
R1487 VTAIL.n33 VTAIL.n4 1.16414
R1488 VTAIL.n117 VTAIL.n88 1.16414
R1489 VTAIL.n77 VTAIL.n48 1.16414
R1490 VTAIL.n83 VTAIL.n81 1.1255
R1491 VTAIL.n37 VTAIL.n1 1.1255
R1492 VTAIL VTAIL.n1 1.04145
R1493 VTAIL VTAIL.n159 0.269897
R1494 VTAIL.n139 VTAIL.n131 0.155672
R1495 VTAIL.n140 VTAIL.n139 0.155672
R1496 VTAIL.n140 VTAIL.n127 0.155672
R1497 VTAIL.n147 VTAIL.n127 0.155672
R1498 VTAIL.n148 VTAIL.n147 0.155672
R1499 VTAIL.n148 VTAIL.n123 0.155672
R1500 VTAIL.n155 VTAIL.n123 0.155672
R1501 VTAIL.n19 VTAIL.n11 0.155672
R1502 VTAIL.n20 VTAIL.n19 0.155672
R1503 VTAIL.n20 VTAIL.n7 0.155672
R1504 VTAIL.n27 VTAIL.n7 0.155672
R1505 VTAIL.n28 VTAIL.n27 0.155672
R1506 VTAIL.n28 VTAIL.n3 0.155672
R1507 VTAIL.n35 VTAIL.n3 0.155672
R1508 VTAIL.n119 VTAIL.n87 0.155672
R1509 VTAIL.n112 VTAIL.n87 0.155672
R1510 VTAIL.n112 VTAIL.n111 0.155672
R1511 VTAIL.n111 VTAIL.n91 0.155672
R1512 VTAIL.n104 VTAIL.n91 0.155672
R1513 VTAIL.n104 VTAIL.n103 0.155672
R1514 VTAIL.n103 VTAIL.n95 0.155672
R1515 VTAIL.n79 VTAIL.n47 0.155672
R1516 VTAIL.n72 VTAIL.n47 0.155672
R1517 VTAIL.n72 VTAIL.n71 0.155672
R1518 VTAIL.n71 VTAIL.n51 0.155672
R1519 VTAIL.n64 VTAIL.n51 0.155672
R1520 VTAIL.n64 VTAIL.n63 0.155672
R1521 VTAIL.n63 VTAIL.n55 0.155672
R1522 VDD2.n69 VDD2.n39 214.453
R1523 VDD2.n30 VDD2.n0 214.453
R1524 VDD2.n70 VDD2.n69 185
R1525 VDD2.n68 VDD2.n67 185
R1526 VDD2.n43 VDD2.n42 185
R1527 VDD2.n62 VDD2.n61 185
R1528 VDD2.n60 VDD2.n59 185
R1529 VDD2.n47 VDD2.n46 185
R1530 VDD2.n54 VDD2.n53 185
R1531 VDD2.n52 VDD2.n51 185
R1532 VDD2.n13 VDD2.n12 185
R1533 VDD2.n15 VDD2.n14 185
R1534 VDD2.n8 VDD2.n7 185
R1535 VDD2.n21 VDD2.n20 185
R1536 VDD2.n23 VDD2.n22 185
R1537 VDD2.n4 VDD2.n3 185
R1538 VDD2.n29 VDD2.n28 185
R1539 VDD2.n31 VDD2.n30 185
R1540 VDD2.n11 VDD2.t9 149.524
R1541 VDD2.n50 VDD2.t0 149.524
R1542 VDD2.n69 VDD2.n68 104.615
R1543 VDD2.n68 VDD2.n42 104.615
R1544 VDD2.n61 VDD2.n42 104.615
R1545 VDD2.n61 VDD2.n60 104.615
R1546 VDD2.n60 VDD2.n46 104.615
R1547 VDD2.n53 VDD2.n46 104.615
R1548 VDD2.n53 VDD2.n52 104.615
R1549 VDD2.n14 VDD2.n13 104.615
R1550 VDD2.n14 VDD2.n7 104.615
R1551 VDD2.n21 VDD2.n7 104.615
R1552 VDD2.n22 VDD2.n21 104.615
R1553 VDD2.n22 VDD2.n3 104.615
R1554 VDD2.n29 VDD2.n3 104.615
R1555 VDD2.n30 VDD2.n29 104.615
R1556 VDD2.n38 VDD2.n37 68.2774
R1557 VDD2 VDD2.n77 68.2745
R1558 VDD2.n76 VDD2.n75 67.3501
R1559 VDD2.n36 VDD2.n35 67.3499
R1560 VDD2.n36 VDD2.n34 52.8896
R1561 VDD2.n52 VDD2.t0 52.3082
R1562 VDD2.n13 VDD2.t9 52.3082
R1563 VDD2.n74 VDD2.n73 51.5793
R1564 VDD2.n74 VDD2.n38 36.1636
R1565 VDD2.n71 VDD2.n70 12.8005
R1566 VDD2.n32 VDD2.n31 12.8005
R1567 VDD2.n67 VDD2.n41 12.0247
R1568 VDD2.n28 VDD2.n2 12.0247
R1569 VDD2.n66 VDD2.n43 11.249
R1570 VDD2.n27 VDD2.n4 11.249
R1571 VDD2.n63 VDD2.n62 10.4732
R1572 VDD2.n24 VDD2.n23 10.4732
R1573 VDD2.n51 VDD2.n50 10.2747
R1574 VDD2.n12 VDD2.n11 10.2747
R1575 VDD2.n59 VDD2.n45 9.69747
R1576 VDD2.n20 VDD2.n6 9.69747
R1577 VDD2.n73 VDD2.n72 9.45567
R1578 VDD2.n34 VDD2.n33 9.45567
R1579 VDD2.n49 VDD2.n48 9.3005
R1580 VDD2.n56 VDD2.n55 9.3005
R1581 VDD2.n58 VDD2.n57 9.3005
R1582 VDD2.n45 VDD2.n44 9.3005
R1583 VDD2.n64 VDD2.n63 9.3005
R1584 VDD2.n66 VDD2.n65 9.3005
R1585 VDD2.n41 VDD2.n40 9.3005
R1586 VDD2.n72 VDD2.n71 9.3005
R1587 VDD2.n10 VDD2.n9 9.3005
R1588 VDD2.n17 VDD2.n16 9.3005
R1589 VDD2.n19 VDD2.n18 9.3005
R1590 VDD2.n6 VDD2.n5 9.3005
R1591 VDD2.n25 VDD2.n24 9.3005
R1592 VDD2.n27 VDD2.n26 9.3005
R1593 VDD2.n2 VDD2.n1 9.3005
R1594 VDD2.n33 VDD2.n32 9.3005
R1595 VDD2.n58 VDD2.n47 8.92171
R1596 VDD2.n19 VDD2.n8 8.92171
R1597 VDD2.n73 VDD2.n39 8.2187
R1598 VDD2.n34 VDD2.n0 8.2187
R1599 VDD2.n55 VDD2.n54 8.14595
R1600 VDD2.n16 VDD2.n15 8.14595
R1601 VDD2.n51 VDD2.n49 7.3702
R1602 VDD2.n12 VDD2.n10 7.3702
R1603 VDD2.n54 VDD2.n49 5.81868
R1604 VDD2.n15 VDD2.n10 5.81868
R1605 VDD2.n71 VDD2.n39 5.3904
R1606 VDD2.n32 VDD2.n0 5.3904
R1607 VDD2.n55 VDD2.n47 5.04292
R1608 VDD2.n16 VDD2.n8 5.04292
R1609 VDD2.n59 VDD2.n58 4.26717
R1610 VDD2.n20 VDD2.n19 4.26717
R1611 VDD2.n62 VDD2.n45 3.49141
R1612 VDD2.n23 VDD2.n6 3.49141
R1613 VDD2.n50 VDD2.n48 2.84305
R1614 VDD2.n11 VDD2.n9 2.84305
R1615 VDD2.n77 VDD2.t4 2.74288
R1616 VDD2.n77 VDD2.t3 2.74288
R1617 VDD2.n75 VDD2.t8 2.74288
R1618 VDD2.n75 VDD2.t6 2.74288
R1619 VDD2.n37 VDD2.t7 2.74288
R1620 VDD2.n37 VDD2.t2 2.74288
R1621 VDD2.n35 VDD2.t5 2.74288
R1622 VDD2.n35 VDD2.t1 2.74288
R1623 VDD2.n63 VDD2.n43 2.71565
R1624 VDD2.n24 VDD2.n4 2.71565
R1625 VDD2.n67 VDD2.n66 1.93989
R1626 VDD2.n28 VDD2.n27 1.93989
R1627 VDD2.n76 VDD2.n74 1.31084
R1628 VDD2.n70 VDD2.n41 1.16414
R1629 VDD2.n31 VDD2.n2 1.16414
R1630 VDD2 VDD2.n76 0.386276
R1631 VDD2.n38 VDD2.n36 0.27274
R1632 VDD2.n72 VDD2.n40 0.155672
R1633 VDD2.n65 VDD2.n40 0.155672
R1634 VDD2.n65 VDD2.n64 0.155672
R1635 VDD2.n64 VDD2.n44 0.155672
R1636 VDD2.n57 VDD2.n44 0.155672
R1637 VDD2.n57 VDD2.n56 0.155672
R1638 VDD2.n56 VDD2.n48 0.155672
R1639 VDD2.n17 VDD2.n9 0.155672
R1640 VDD2.n18 VDD2.n17 0.155672
R1641 VDD2.n18 VDD2.n5 0.155672
R1642 VDD2.n25 VDD2.n5 0.155672
R1643 VDD2.n26 VDD2.n25 0.155672
R1644 VDD2.n26 VDD2.n1 0.155672
R1645 VDD2.n33 VDD2.n1 0.155672
R1646 VP.n13 VP.t4 197.749
R1647 VP.n30 VP.t7 179.232
R1648 VP.n47 VP.t0 179.232
R1649 VP.n27 VP.t6 179.232
R1650 VP.n15 VP.n14 161.3
R1651 VP.n16 VP.n11 161.3
R1652 VP.n18 VP.n17 161.3
R1653 VP.n20 VP.n19 161.3
R1654 VP.n21 VP.n9 161.3
R1655 VP.n23 VP.n22 161.3
R1656 VP.n25 VP.n24 161.3
R1657 VP.n26 VP.n7 161.3
R1658 VP.n46 VP.n0 161.3
R1659 VP.n45 VP.n44 161.3
R1660 VP.n43 VP.n42 161.3
R1661 VP.n41 VP.n2 161.3
R1662 VP.n40 VP.n39 161.3
R1663 VP.n38 VP.n37 161.3
R1664 VP.n36 VP.n4 161.3
R1665 VP.n35 VP.n34 161.3
R1666 VP.n33 VP.n32 161.3
R1667 VP.n31 VP.n6 161.3
R1668 VP.n5 VP.t2 146.22
R1669 VP.n3 VP.t9 146.22
R1670 VP.n1 VP.t5 146.22
R1671 VP.n8 VP.t8 146.22
R1672 VP.n10 VP.t1 146.22
R1673 VP.n12 VP.t3 146.22
R1674 VP.n28 VP.n27 80.6037
R1675 VP.n48 VP.n47 80.6037
R1676 VP.n30 VP.n29 80.6037
R1677 VP.n13 VP.n12 44.6572
R1678 VP.n29 VP.n28 41.9332
R1679 VP.n36 VP.n35 41.5458
R1680 VP.n42 VP.n41 41.5458
R1681 VP.n22 VP.n21 41.5458
R1682 VP.n16 VP.n15 41.5458
R1683 VP.n37 VP.n36 39.6083
R1684 VP.n41 VP.n40 39.6083
R1685 VP.n21 VP.n20 39.6083
R1686 VP.n17 VP.n16 39.6083
R1687 VP.n32 VP.n31 37.6707
R1688 VP.n46 VP.n45 37.6707
R1689 VP.n26 VP.n25 37.6707
R1690 VP.n14 VP.n13 29.7202
R1691 VP.n31 VP.n30 28.4823
R1692 VP.n47 VP.n46 28.4823
R1693 VP.n27 VP.n26 28.4823
R1694 VP.n35 VP.n5 13.2801
R1695 VP.n42 VP.n1 13.2801
R1696 VP.n22 VP.n8 13.2801
R1697 VP.n15 VP.n12 13.2801
R1698 VP.n37 VP.n3 12.2964
R1699 VP.n40 VP.n3 12.2964
R1700 VP.n17 VP.n10 12.2964
R1701 VP.n20 VP.n10 12.2964
R1702 VP.n32 VP.n5 11.3127
R1703 VP.n45 VP.n1 11.3127
R1704 VP.n25 VP.n8 11.3127
R1705 VP.n28 VP.n7 0.285035
R1706 VP.n29 VP.n6 0.285035
R1707 VP.n48 VP.n0 0.285035
R1708 VP.n14 VP.n11 0.189894
R1709 VP.n18 VP.n11 0.189894
R1710 VP.n19 VP.n18 0.189894
R1711 VP.n19 VP.n9 0.189894
R1712 VP.n23 VP.n9 0.189894
R1713 VP.n24 VP.n23 0.189894
R1714 VP.n24 VP.n7 0.189894
R1715 VP.n33 VP.n6 0.189894
R1716 VP.n34 VP.n33 0.189894
R1717 VP.n34 VP.n4 0.189894
R1718 VP.n38 VP.n4 0.189894
R1719 VP.n39 VP.n38 0.189894
R1720 VP.n39 VP.n2 0.189894
R1721 VP.n43 VP.n2 0.189894
R1722 VP.n44 VP.n43 0.189894
R1723 VP.n44 VP.n0 0.189894
R1724 VP VP.n48 0.146778
R1725 VDD1.n30 VDD1.n0 214.453
R1726 VDD1.n67 VDD1.n37 214.453
R1727 VDD1.n31 VDD1.n30 185
R1728 VDD1.n29 VDD1.n28 185
R1729 VDD1.n4 VDD1.n3 185
R1730 VDD1.n23 VDD1.n22 185
R1731 VDD1.n21 VDD1.n20 185
R1732 VDD1.n8 VDD1.n7 185
R1733 VDD1.n15 VDD1.n14 185
R1734 VDD1.n13 VDD1.n12 185
R1735 VDD1.n50 VDD1.n49 185
R1736 VDD1.n52 VDD1.n51 185
R1737 VDD1.n45 VDD1.n44 185
R1738 VDD1.n58 VDD1.n57 185
R1739 VDD1.n60 VDD1.n59 185
R1740 VDD1.n41 VDD1.n40 185
R1741 VDD1.n66 VDD1.n65 185
R1742 VDD1.n68 VDD1.n67 185
R1743 VDD1.n48 VDD1.t2 149.524
R1744 VDD1.n11 VDD1.t5 149.524
R1745 VDD1.n30 VDD1.n29 104.615
R1746 VDD1.n29 VDD1.n3 104.615
R1747 VDD1.n22 VDD1.n3 104.615
R1748 VDD1.n22 VDD1.n21 104.615
R1749 VDD1.n21 VDD1.n7 104.615
R1750 VDD1.n14 VDD1.n7 104.615
R1751 VDD1.n14 VDD1.n13 104.615
R1752 VDD1.n51 VDD1.n50 104.615
R1753 VDD1.n51 VDD1.n44 104.615
R1754 VDD1.n58 VDD1.n44 104.615
R1755 VDD1.n59 VDD1.n58 104.615
R1756 VDD1.n59 VDD1.n40 104.615
R1757 VDD1.n66 VDD1.n40 104.615
R1758 VDD1.n67 VDD1.n66 104.615
R1759 VDD1.n75 VDD1.n74 68.2774
R1760 VDD1.n36 VDD1.n35 67.3501
R1761 VDD1.n77 VDD1.n76 67.3499
R1762 VDD1.n73 VDD1.n72 67.3499
R1763 VDD1.n36 VDD1.n34 52.8896
R1764 VDD1.n73 VDD1.n71 52.8896
R1765 VDD1.n13 VDD1.t5 52.3082
R1766 VDD1.n50 VDD1.t2 52.3082
R1767 VDD1.n77 VDD1.n75 37.4018
R1768 VDD1.n32 VDD1.n31 12.8005
R1769 VDD1.n69 VDD1.n68 12.8005
R1770 VDD1.n28 VDD1.n2 12.0247
R1771 VDD1.n65 VDD1.n39 12.0247
R1772 VDD1.n27 VDD1.n4 11.249
R1773 VDD1.n64 VDD1.n41 11.249
R1774 VDD1.n24 VDD1.n23 10.4732
R1775 VDD1.n61 VDD1.n60 10.4732
R1776 VDD1.n12 VDD1.n11 10.2747
R1777 VDD1.n49 VDD1.n48 10.2747
R1778 VDD1.n20 VDD1.n6 9.69747
R1779 VDD1.n57 VDD1.n43 9.69747
R1780 VDD1.n34 VDD1.n33 9.45567
R1781 VDD1.n71 VDD1.n70 9.45567
R1782 VDD1.n10 VDD1.n9 9.3005
R1783 VDD1.n17 VDD1.n16 9.3005
R1784 VDD1.n19 VDD1.n18 9.3005
R1785 VDD1.n6 VDD1.n5 9.3005
R1786 VDD1.n25 VDD1.n24 9.3005
R1787 VDD1.n27 VDD1.n26 9.3005
R1788 VDD1.n2 VDD1.n1 9.3005
R1789 VDD1.n33 VDD1.n32 9.3005
R1790 VDD1.n47 VDD1.n46 9.3005
R1791 VDD1.n54 VDD1.n53 9.3005
R1792 VDD1.n56 VDD1.n55 9.3005
R1793 VDD1.n43 VDD1.n42 9.3005
R1794 VDD1.n62 VDD1.n61 9.3005
R1795 VDD1.n64 VDD1.n63 9.3005
R1796 VDD1.n39 VDD1.n38 9.3005
R1797 VDD1.n70 VDD1.n69 9.3005
R1798 VDD1.n19 VDD1.n8 8.92171
R1799 VDD1.n56 VDD1.n45 8.92171
R1800 VDD1.n34 VDD1.n0 8.2187
R1801 VDD1.n71 VDD1.n37 8.2187
R1802 VDD1.n16 VDD1.n15 8.14595
R1803 VDD1.n53 VDD1.n52 8.14595
R1804 VDD1.n12 VDD1.n10 7.3702
R1805 VDD1.n49 VDD1.n47 7.3702
R1806 VDD1.n15 VDD1.n10 5.81868
R1807 VDD1.n52 VDD1.n47 5.81868
R1808 VDD1.n32 VDD1.n0 5.3904
R1809 VDD1.n69 VDD1.n37 5.3904
R1810 VDD1.n16 VDD1.n8 5.04292
R1811 VDD1.n53 VDD1.n45 5.04292
R1812 VDD1.n20 VDD1.n19 4.26717
R1813 VDD1.n57 VDD1.n56 4.26717
R1814 VDD1.n23 VDD1.n6 3.49141
R1815 VDD1.n60 VDD1.n43 3.49141
R1816 VDD1.n11 VDD1.n9 2.84305
R1817 VDD1.n48 VDD1.n46 2.84305
R1818 VDD1.n76 VDD1.t1 2.74288
R1819 VDD1.n76 VDD1.t3 2.74288
R1820 VDD1.n35 VDD1.t6 2.74288
R1821 VDD1.n35 VDD1.t8 2.74288
R1822 VDD1.n74 VDD1.t4 2.74288
R1823 VDD1.n74 VDD1.t9 2.74288
R1824 VDD1.n72 VDD1.t7 2.74288
R1825 VDD1.n72 VDD1.t0 2.74288
R1826 VDD1.n24 VDD1.n4 2.71565
R1827 VDD1.n61 VDD1.n41 2.71565
R1828 VDD1.n28 VDD1.n27 1.93989
R1829 VDD1.n65 VDD1.n64 1.93989
R1830 VDD1.n31 VDD1.n2 1.16414
R1831 VDD1.n68 VDD1.n39 1.16414
R1832 VDD1 VDD1.n77 0.925069
R1833 VDD1 VDD1.n36 0.386276
R1834 VDD1.n75 VDD1.n73 0.27274
R1835 VDD1.n33 VDD1.n1 0.155672
R1836 VDD1.n26 VDD1.n1 0.155672
R1837 VDD1.n26 VDD1.n25 0.155672
R1838 VDD1.n25 VDD1.n5 0.155672
R1839 VDD1.n18 VDD1.n5 0.155672
R1840 VDD1.n18 VDD1.n17 0.155672
R1841 VDD1.n17 VDD1.n9 0.155672
R1842 VDD1.n54 VDD1.n46 0.155672
R1843 VDD1.n55 VDD1.n54 0.155672
R1844 VDD1.n55 VDD1.n42 0.155672
R1845 VDD1.n62 VDD1.n42 0.155672
R1846 VDD1.n63 VDD1.n62 0.155672
R1847 VDD1.n63 VDD1.n38 0.155672
R1848 VDD1.n70 VDD1.n38 0.155672
C0 VDD1 VN 0.150075f
C1 VTAIL VN 5.56854f
C2 VN VDD2 5.3238f
C3 VN VP 5.43207f
C4 VDD1 VTAIL 8.22763f
C5 VDD1 VDD2 1.26987f
C6 VDD1 VP 5.57405f
C7 VTAIL VDD2 8.26875f
C8 VTAIL VP 5.58287f
C9 VDD2 VP 0.403236f
C10 VDD2 B 4.687274f
C11 VDD1 B 4.649414f
C12 VTAIL B 5.193105f
C13 VN B 11.1369f
C14 VP B 9.55302f
C15 VDD1.n0 B 0.031679f
C16 VDD1.n1 B 0.02328f
C17 VDD1.n2 B 0.01251f
C18 VDD1.n3 B 0.029569f
C19 VDD1.n4 B 0.013246f
C20 VDD1.n5 B 0.02328f
C21 VDD1.n6 B 0.01251f
C22 VDD1.n7 B 0.029569f
C23 VDD1.n8 B 0.013246f
C24 VDD1.n9 B 0.679405f
C25 VDD1.n10 B 0.01251f
C26 VDD1.t5 B 0.049371f
C27 VDD1.n11 B 0.125179f
C28 VDD1.n12 B 0.020903f
C29 VDD1.n13 B 0.022176f
C30 VDD1.n14 B 0.029569f
C31 VDD1.n15 B 0.013246f
C32 VDD1.n16 B 0.01251f
C33 VDD1.n17 B 0.02328f
C34 VDD1.n18 B 0.02328f
C35 VDD1.n19 B 0.01251f
C36 VDD1.n20 B 0.013246f
C37 VDD1.n21 B 0.029569f
C38 VDD1.n22 B 0.029569f
C39 VDD1.n23 B 0.013246f
C40 VDD1.n24 B 0.01251f
C41 VDD1.n25 B 0.02328f
C42 VDD1.n26 B 0.02328f
C43 VDD1.n27 B 0.01251f
C44 VDD1.n28 B 0.013246f
C45 VDD1.n29 B 0.029569f
C46 VDD1.n30 B 0.060362f
C47 VDD1.n31 B 0.013246f
C48 VDD1.n32 B 0.024461f
C49 VDD1.n33 B 0.058263f
C50 VDD1.n34 B 0.081757f
C51 VDD1.t6 B 0.132824f
C52 VDD1.t8 B 0.132824f
C53 VDD1.n35 B 1.14036f
C54 VDD1.n36 B 0.452013f
C55 VDD1.n37 B 0.031679f
C56 VDD1.n38 B 0.02328f
C57 VDD1.n39 B 0.01251f
C58 VDD1.n40 B 0.029569f
C59 VDD1.n41 B 0.013246f
C60 VDD1.n42 B 0.02328f
C61 VDD1.n43 B 0.01251f
C62 VDD1.n44 B 0.029569f
C63 VDD1.n45 B 0.013246f
C64 VDD1.n46 B 0.679405f
C65 VDD1.n47 B 0.01251f
C66 VDD1.t2 B 0.049371f
C67 VDD1.n48 B 0.125179f
C68 VDD1.n49 B 0.020903f
C69 VDD1.n50 B 0.022176f
C70 VDD1.n51 B 0.029569f
C71 VDD1.n52 B 0.013246f
C72 VDD1.n53 B 0.01251f
C73 VDD1.n54 B 0.02328f
C74 VDD1.n55 B 0.02328f
C75 VDD1.n56 B 0.01251f
C76 VDD1.n57 B 0.013246f
C77 VDD1.n58 B 0.029569f
C78 VDD1.n59 B 0.029569f
C79 VDD1.n60 B 0.013246f
C80 VDD1.n61 B 0.01251f
C81 VDD1.n62 B 0.02328f
C82 VDD1.n63 B 0.02328f
C83 VDD1.n64 B 0.01251f
C84 VDD1.n65 B 0.013246f
C85 VDD1.n66 B 0.029569f
C86 VDD1.n67 B 0.060362f
C87 VDD1.n68 B 0.013246f
C88 VDD1.n69 B 0.024461f
C89 VDD1.n70 B 0.058263f
C90 VDD1.n71 B 0.081757f
C91 VDD1.t7 B 0.132824f
C92 VDD1.t0 B 0.132824f
C93 VDD1.n72 B 1.14036f
C94 VDD1.n73 B 0.445484f
C95 VDD1.t4 B 0.132824f
C96 VDD1.t9 B 0.132824f
C97 VDD1.n74 B 1.14525f
C98 VDD1.n75 B 1.81921f
C99 VDD1.t1 B 0.132824f
C100 VDD1.t3 B 0.132824f
C101 VDD1.n76 B 1.14036f
C102 VDD1.n77 B 2.0542f
C103 VP.n0 B 0.047501f
C104 VP.t5 B 0.81756f
C105 VP.n1 B 0.318299f
C106 VP.n2 B 0.035598f
C107 VP.t9 B 0.81756f
C108 VP.n3 B 0.318299f
C109 VP.n4 B 0.035598f
C110 VP.t2 B 0.81756f
C111 VP.n5 B 0.318299f
C112 VP.n6 B 0.047501f
C113 VP.n7 B 0.047501f
C114 VP.t6 B 0.882062f
C115 VP.t8 B 0.81756f
C116 VP.n8 B 0.318299f
C117 VP.n9 B 0.035598f
C118 VP.t1 B 0.81756f
C119 VP.n10 B 0.318299f
C120 VP.n11 B 0.035598f
C121 VP.t3 B 0.81756f
C122 VP.n12 B 0.363167f
C123 VP.t4 B 0.918628f
C124 VP.n13 B 0.376905f
C125 VP.n14 B 0.182304f
C126 VP.n15 B 0.055011f
C127 VP.n16 B 0.028796f
C128 VP.n17 B 0.054413f
C129 VP.n18 B 0.035598f
C130 VP.n19 B 0.035598f
C131 VP.n20 B 0.054413f
C132 VP.n21 B 0.028796f
C133 VP.n22 B 0.055011f
C134 VP.n23 B 0.035598f
C135 VP.n24 B 0.035598f
C136 VP.n25 B 0.053619f
C137 VP.n26 B 0.020827f
C138 VP.n27 B 0.382281f
C139 VP.n28 B 1.4781f
C140 VP.n29 B 1.5087f
C141 VP.t7 B 0.882062f
C142 VP.n30 B 0.382281f
C143 VP.n31 B 0.020827f
C144 VP.n32 B 0.053619f
C145 VP.n33 B 0.035598f
C146 VP.n34 B 0.035598f
C147 VP.n35 B 0.055011f
C148 VP.n36 B 0.028796f
C149 VP.n37 B 0.054413f
C150 VP.n38 B 0.035598f
C151 VP.n39 B 0.035598f
C152 VP.n40 B 0.054413f
C153 VP.n41 B 0.028796f
C154 VP.n42 B 0.055011f
C155 VP.n43 B 0.035598f
C156 VP.n44 B 0.035598f
C157 VP.n45 B 0.053619f
C158 VP.n46 B 0.020827f
C159 VP.t0 B 0.882062f
C160 VP.n47 B 0.382281f
C161 VP.n48 B 0.033339f
C162 VDD2.n0 B 0.031416f
C163 VDD2.n1 B 0.023087f
C164 VDD2.n2 B 0.012406f
C165 VDD2.n3 B 0.029323f
C166 VDD2.n4 B 0.013136f
C167 VDD2.n5 B 0.023087f
C168 VDD2.n6 B 0.012406f
C169 VDD2.n7 B 0.029323f
C170 VDD2.n8 B 0.013136f
C171 VDD2.n9 B 0.673757f
C172 VDD2.n10 B 0.012406f
C173 VDD2.t9 B 0.04896f
C174 VDD2.n11 B 0.124139f
C175 VDD2.n12 B 0.020729f
C176 VDD2.n13 B 0.021992f
C177 VDD2.n14 B 0.029323f
C178 VDD2.n15 B 0.013136f
C179 VDD2.n16 B 0.012406f
C180 VDD2.n17 B 0.023087f
C181 VDD2.n18 B 0.023087f
C182 VDD2.n19 B 0.012406f
C183 VDD2.n20 B 0.013136f
C184 VDD2.n21 B 0.029323f
C185 VDD2.n22 B 0.029323f
C186 VDD2.n23 B 0.013136f
C187 VDD2.n24 B 0.012406f
C188 VDD2.n25 B 0.023087f
C189 VDD2.n26 B 0.023087f
C190 VDD2.n27 B 0.012406f
C191 VDD2.n28 B 0.013136f
C192 VDD2.n29 B 0.029323f
C193 VDD2.n30 B 0.05986f
C194 VDD2.n31 B 0.013136f
C195 VDD2.n32 B 0.024257f
C196 VDD2.n33 B 0.057779f
C197 VDD2.n34 B 0.081077f
C198 VDD2.t5 B 0.13172f
C199 VDD2.t1 B 0.13172f
C200 VDD2.n35 B 1.13088f
C201 VDD2.n36 B 0.44178f
C202 VDD2.t7 B 0.13172f
C203 VDD2.t2 B 0.13172f
C204 VDD2.n37 B 1.13573f
C205 VDD2.n38 B 1.72444f
C206 VDD2.n39 B 0.031416f
C207 VDD2.n40 B 0.023087f
C208 VDD2.n41 B 0.012406f
C209 VDD2.n42 B 0.029323f
C210 VDD2.n43 B 0.013136f
C211 VDD2.n44 B 0.023087f
C212 VDD2.n45 B 0.012406f
C213 VDD2.n46 B 0.029323f
C214 VDD2.n47 B 0.013136f
C215 VDD2.n48 B 0.673757f
C216 VDD2.n49 B 0.012406f
C217 VDD2.t0 B 0.04896f
C218 VDD2.n50 B 0.124139f
C219 VDD2.n51 B 0.020729f
C220 VDD2.n52 B 0.021992f
C221 VDD2.n53 B 0.029323f
C222 VDD2.n54 B 0.013136f
C223 VDD2.n55 B 0.012406f
C224 VDD2.n56 B 0.023087f
C225 VDD2.n57 B 0.023087f
C226 VDD2.n58 B 0.012406f
C227 VDD2.n59 B 0.013136f
C228 VDD2.n60 B 0.029323f
C229 VDD2.n61 B 0.029323f
C230 VDD2.n62 B 0.013136f
C231 VDD2.n63 B 0.012406f
C232 VDD2.n64 B 0.023087f
C233 VDD2.n65 B 0.023087f
C234 VDD2.n66 B 0.012406f
C235 VDD2.n67 B 0.013136f
C236 VDD2.n68 B 0.029323f
C237 VDD2.n69 B 0.05986f
C238 VDD2.n70 B 0.013136f
C239 VDD2.n71 B 0.024257f
C240 VDD2.n72 B 0.057779f
C241 VDD2.n73 B 0.077498f
C242 VDD2.n74 B 1.8192f
C243 VDD2.t8 B 0.13172f
C244 VDD2.t6 B 0.13172f
C245 VDD2.n75 B 1.13088f
C246 VDD2.n76 B 0.307373f
C247 VDD2.t4 B 0.13172f
C248 VDD2.t3 B 0.13172f
C249 VDD2.n77 B 1.13571f
C250 VTAIL.t13 B 0.148933f
C251 VTAIL.t11 B 0.148933f
C252 VTAIL.n0 B 1.21285f
C253 VTAIL.n1 B 0.417388f
C254 VTAIL.n2 B 0.035521f
C255 VTAIL.n3 B 0.026104f
C256 VTAIL.n4 B 0.014027f
C257 VTAIL.n5 B 0.033154f
C258 VTAIL.n6 B 0.014852f
C259 VTAIL.n7 B 0.026104f
C260 VTAIL.n8 B 0.014027f
C261 VTAIL.n9 B 0.033154f
C262 VTAIL.n10 B 0.014852f
C263 VTAIL.n11 B 0.761801f
C264 VTAIL.n12 B 0.014027f
C265 VTAIL.t3 B 0.055358f
C266 VTAIL.n13 B 0.140361f
C267 VTAIL.n14 B 0.023438f
C268 VTAIL.n15 B 0.024866f
C269 VTAIL.n16 B 0.033154f
C270 VTAIL.n17 B 0.014852f
C271 VTAIL.n18 B 0.014027f
C272 VTAIL.n19 B 0.026104f
C273 VTAIL.n20 B 0.026104f
C274 VTAIL.n21 B 0.014027f
C275 VTAIL.n22 B 0.014852f
C276 VTAIL.n23 B 0.033154f
C277 VTAIL.n24 B 0.033154f
C278 VTAIL.n25 B 0.014852f
C279 VTAIL.n26 B 0.014027f
C280 VTAIL.n27 B 0.026104f
C281 VTAIL.n28 B 0.026104f
C282 VTAIL.n29 B 0.014027f
C283 VTAIL.n30 B 0.014852f
C284 VTAIL.n31 B 0.033154f
C285 VTAIL.n32 B 0.067682f
C286 VTAIL.n33 B 0.014852f
C287 VTAIL.n34 B 0.027427f
C288 VTAIL.n35 B 0.065329f
C289 VTAIL.n36 B 0.069637f
C290 VTAIL.n37 B 0.229958f
C291 VTAIL.t4 B 0.148933f
C292 VTAIL.t1 B 0.148933f
C293 VTAIL.n38 B 1.21285f
C294 VTAIL.n39 B 0.455637f
C295 VTAIL.t0 B 0.148933f
C296 VTAIL.t2 B 0.148933f
C297 VTAIL.n40 B 1.21285f
C298 VTAIL.n41 B 1.44396f
C299 VTAIL.t16 B 0.148933f
C300 VTAIL.t18 B 0.148933f
C301 VTAIL.n42 B 1.21286f
C302 VTAIL.n43 B 1.44395f
C303 VTAIL.t14 B 0.148933f
C304 VTAIL.t15 B 0.148933f
C305 VTAIL.n44 B 1.21286f
C306 VTAIL.n45 B 0.455628f
C307 VTAIL.n46 B 0.035521f
C308 VTAIL.n47 B 0.026104f
C309 VTAIL.n48 B 0.014027f
C310 VTAIL.n49 B 0.033154f
C311 VTAIL.n50 B 0.014852f
C312 VTAIL.n51 B 0.026104f
C313 VTAIL.n52 B 0.014027f
C314 VTAIL.n53 B 0.033154f
C315 VTAIL.n54 B 0.014852f
C316 VTAIL.n55 B 0.761801f
C317 VTAIL.n56 B 0.014027f
C318 VTAIL.t12 B 0.055358f
C319 VTAIL.n57 B 0.140361f
C320 VTAIL.n58 B 0.023438f
C321 VTAIL.n59 B 0.024866f
C322 VTAIL.n60 B 0.033154f
C323 VTAIL.n61 B 0.014852f
C324 VTAIL.n62 B 0.014027f
C325 VTAIL.n63 B 0.026104f
C326 VTAIL.n64 B 0.026104f
C327 VTAIL.n65 B 0.014027f
C328 VTAIL.n66 B 0.014852f
C329 VTAIL.n67 B 0.033154f
C330 VTAIL.n68 B 0.033154f
C331 VTAIL.n69 B 0.014852f
C332 VTAIL.n70 B 0.014027f
C333 VTAIL.n71 B 0.026104f
C334 VTAIL.n72 B 0.026104f
C335 VTAIL.n73 B 0.014027f
C336 VTAIL.n74 B 0.014852f
C337 VTAIL.n75 B 0.033154f
C338 VTAIL.n76 B 0.067682f
C339 VTAIL.n77 B 0.014852f
C340 VTAIL.n78 B 0.027427f
C341 VTAIL.n79 B 0.065329f
C342 VTAIL.n80 B 0.069637f
C343 VTAIL.n81 B 0.229958f
C344 VTAIL.t6 B 0.148933f
C345 VTAIL.t9 B 0.148933f
C346 VTAIL.n82 B 1.21286f
C347 VTAIL.n83 B 0.440038f
C348 VTAIL.t5 B 0.148933f
C349 VTAIL.t7 B 0.148933f
C350 VTAIL.n84 B 1.21286f
C351 VTAIL.n85 B 0.455628f
C352 VTAIL.n86 B 0.035521f
C353 VTAIL.n87 B 0.026104f
C354 VTAIL.n88 B 0.014027f
C355 VTAIL.n89 B 0.033154f
C356 VTAIL.n90 B 0.014852f
C357 VTAIL.n91 B 0.026104f
C358 VTAIL.n92 B 0.014027f
C359 VTAIL.n93 B 0.033154f
C360 VTAIL.n94 B 0.014852f
C361 VTAIL.n95 B 0.761801f
C362 VTAIL.n96 B 0.014027f
C363 VTAIL.t8 B 0.055358f
C364 VTAIL.n97 B 0.140361f
C365 VTAIL.n98 B 0.023438f
C366 VTAIL.n99 B 0.024866f
C367 VTAIL.n100 B 0.033154f
C368 VTAIL.n101 B 0.014852f
C369 VTAIL.n102 B 0.014027f
C370 VTAIL.n103 B 0.026104f
C371 VTAIL.n104 B 0.026104f
C372 VTAIL.n105 B 0.014027f
C373 VTAIL.n106 B 0.014852f
C374 VTAIL.n107 B 0.033154f
C375 VTAIL.n108 B 0.033154f
C376 VTAIL.n109 B 0.014852f
C377 VTAIL.n110 B 0.014027f
C378 VTAIL.n111 B 0.026104f
C379 VTAIL.n112 B 0.026104f
C380 VTAIL.n113 B 0.014027f
C381 VTAIL.n114 B 0.014852f
C382 VTAIL.n115 B 0.033154f
C383 VTAIL.n116 B 0.067682f
C384 VTAIL.n117 B 0.014852f
C385 VTAIL.n118 B 0.027427f
C386 VTAIL.n119 B 0.065329f
C387 VTAIL.n120 B 0.069637f
C388 VTAIL.n121 B 1.12365f
C389 VTAIL.n122 B 0.035521f
C390 VTAIL.n123 B 0.026104f
C391 VTAIL.n124 B 0.014027f
C392 VTAIL.n125 B 0.033154f
C393 VTAIL.n126 B 0.014852f
C394 VTAIL.n127 B 0.026104f
C395 VTAIL.n128 B 0.014027f
C396 VTAIL.n129 B 0.033154f
C397 VTAIL.n130 B 0.014852f
C398 VTAIL.n131 B 0.761801f
C399 VTAIL.n132 B 0.014027f
C400 VTAIL.t19 B 0.055358f
C401 VTAIL.n133 B 0.140361f
C402 VTAIL.n134 B 0.023438f
C403 VTAIL.n135 B 0.024866f
C404 VTAIL.n136 B 0.033154f
C405 VTAIL.n137 B 0.014852f
C406 VTAIL.n138 B 0.014027f
C407 VTAIL.n139 B 0.026104f
C408 VTAIL.n140 B 0.026104f
C409 VTAIL.n141 B 0.014027f
C410 VTAIL.n142 B 0.014852f
C411 VTAIL.n143 B 0.033154f
C412 VTAIL.n144 B 0.033154f
C413 VTAIL.n145 B 0.014852f
C414 VTAIL.n146 B 0.014027f
C415 VTAIL.n147 B 0.026104f
C416 VTAIL.n148 B 0.026104f
C417 VTAIL.n149 B 0.014027f
C418 VTAIL.n150 B 0.014852f
C419 VTAIL.n151 B 0.033154f
C420 VTAIL.n152 B 0.067682f
C421 VTAIL.n153 B 0.014852f
C422 VTAIL.n154 B 0.027427f
C423 VTAIL.n155 B 0.065329f
C424 VTAIL.n156 B 0.069637f
C425 VTAIL.n157 B 1.12365f
C426 VTAIL.t17 B 0.148933f
C427 VTAIL.t10 B 0.148933f
C428 VTAIL.n158 B 1.21285f
C429 VTAIL.n159 B 0.368081f
C430 VN.n0 B 0.046502f
C431 VN.t2 B 0.800372f
C432 VN.n1 B 0.311608f
C433 VN.n2 B 0.034849f
C434 VN.t8 B 0.800372f
C435 VN.n3 B 0.311608f
C436 VN.n4 B 0.034849f
C437 VN.t4 B 0.800372f
C438 VN.n5 B 0.355532f
C439 VN.t0 B 0.899315f
C440 VN.n6 B 0.368981f
C441 VN.n7 B 0.178471f
C442 VN.n8 B 0.053855f
C443 VN.n9 B 0.028191f
C444 VN.n10 B 0.053269f
C445 VN.n11 B 0.034849f
C446 VN.n12 B 0.034849f
C447 VN.n13 B 0.053269f
C448 VN.n14 B 0.028191f
C449 VN.n15 B 0.053855f
C450 VN.n16 B 0.034849f
C451 VN.n17 B 0.034849f
C452 VN.n18 B 0.052492f
C453 VN.n19 B 0.020389f
C454 VN.t7 B 0.863518f
C455 VN.n20 B 0.374244f
C456 VN.n21 B 0.032638f
C457 VN.n22 B 0.046502f
C458 VN.t1 B 0.800372f
C459 VN.n23 B 0.311608f
C460 VN.n24 B 0.034849f
C461 VN.t3 B 0.800372f
C462 VN.n25 B 0.311608f
C463 VN.n26 B 0.034849f
C464 VN.t5 B 0.800372f
C465 VN.n27 B 0.355532f
C466 VN.t6 B 0.899315f
C467 VN.n28 B 0.368981f
C468 VN.n29 B 0.178471f
C469 VN.n30 B 0.053855f
C470 VN.n31 B 0.028191f
C471 VN.n32 B 0.053269f
C472 VN.n33 B 0.034849f
C473 VN.n34 B 0.034849f
C474 VN.n35 B 0.053269f
C475 VN.n36 B 0.028191f
C476 VN.n37 B 0.053855f
C477 VN.n38 B 0.034849f
C478 VN.n39 B 0.034849f
C479 VN.n40 B 0.052492f
C480 VN.n41 B 0.020389f
C481 VN.t9 B 0.863518f
C482 VN.n42 B 0.374244f
C483 VN.n43 B 1.46658f
.ends

