* NGSPICE file created from diff_pair_sample_1499.ext - technology: sky130A

.subckt diff_pair_sample_1499 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n4910_n4582# sky130_fd_pr__pfet_01v8 ad=7.0473 pd=36.92 as=0 ps=0 w=18.07 l=3.61
X1 VDD1.t7 VP.t0 VTAIL.t10 w_n4910_n4582# sky130_fd_pr__pfet_01v8 ad=2.98155 pd=18.4 as=7.0473 ps=36.92 w=18.07 l=3.61
X2 VTAIL.t12 VP.t1 VDD1.t6 w_n4910_n4582# sky130_fd_pr__pfet_01v8 ad=7.0473 pd=36.92 as=2.98155 ps=18.4 w=18.07 l=3.61
X3 VDD2.t7 VN.t0 VTAIL.t15 w_n4910_n4582# sky130_fd_pr__pfet_01v8 ad=2.98155 pd=18.4 as=7.0473 ps=36.92 w=18.07 l=3.61
X4 VTAIL.t4 VN.t1 VDD2.t6 w_n4910_n4582# sky130_fd_pr__pfet_01v8 ad=2.98155 pd=18.4 as=2.98155 ps=18.4 w=18.07 l=3.61
X5 VDD1.t5 VP.t2 VTAIL.t8 w_n4910_n4582# sky130_fd_pr__pfet_01v8 ad=2.98155 pd=18.4 as=7.0473 ps=36.92 w=18.07 l=3.61
X6 VTAIL.t7 VP.t3 VDD1.t4 w_n4910_n4582# sky130_fd_pr__pfet_01v8 ad=2.98155 pd=18.4 as=2.98155 ps=18.4 w=18.07 l=3.61
X7 B.t8 B.t6 B.t7 w_n4910_n4582# sky130_fd_pr__pfet_01v8 ad=7.0473 pd=36.92 as=0 ps=0 w=18.07 l=3.61
X8 VDD2.t5 VN.t2 VTAIL.t6 w_n4910_n4582# sky130_fd_pr__pfet_01v8 ad=2.98155 pd=18.4 as=7.0473 ps=36.92 w=18.07 l=3.61
X9 VDD1.t3 VP.t4 VTAIL.t9 w_n4910_n4582# sky130_fd_pr__pfet_01v8 ad=2.98155 pd=18.4 as=2.98155 ps=18.4 w=18.07 l=3.61
X10 VTAIL.t13 VP.t5 VDD1.t2 w_n4910_n4582# sky130_fd_pr__pfet_01v8 ad=7.0473 pd=36.92 as=2.98155 ps=18.4 w=18.07 l=3.61
X11 VDD1.t1 VP.t6 VTAIL.t14 w_n4910_n4582# sky130_fd_pr__pfet_01v8 ad=2.98155 pd=18.4 as=2.98155 ps=18.4 w=18.07 l=3.61
X12 VDD2.t4 VN.t3 VTAIL.t3 w_n4910_n4582# sky130_fd_pr__pfet_01v8 ad=2.98155 pd=18.4 as=2.98155 ps=18.4 w=18.07 l=3.61
X13 B.t5 B.t3 B.t4 w_n4910_n4582# sky130_fd_pr__pfet_01v8 ad=7.0473 pd=36.92 as=0 ps=0 w=18.07 l=3.61
X14 VTAIL.t2 VN.t4 VDD2.t3 w_n4910_n4582# sky130_fd_pr__pfet_01v8 ad=7.0473 pd=36.92 as=2.98155 ps=18.4 w=18.07 l=3.61
X15 VTAIL.t11 VP.t7 VDD1.t0 w_n4910_n4582# sky130_fd_pr__pfet_01v8 ad=2.98155 pd=18.4 as=2.98155 ps=18.4 w=18.07 l=3.61
X16 B.t2 B.t0 B.t1 w_n4910_n4582# sky130_fd_pr__pfet_01v8 ad=7.0473 pd=36.92 as=0 ps=0 w=18.07 l=3.61
X17 VTAIL.t1 VN.t5 VDD2.t2 w_n4910_n4582# sky130_fd_pr__pfet_01v8 ad=7.0473 pd=36.92 as=2.98155 ps=18.4 w=18.07 l=3.61
X18 VDD2.t1 VN.t6 VTAIL.t5 w_n4910_n4582# sky130_fd_pr__pfet_01v8 ad=2.98155 pd=18.4 as=2.98155 ps=18.4 w=18.07 l=3.61
X19 VTAIL.t0 VN.t7 VDD2.t0 w_n4910_n4582# sky130_fd_pr__pfet_01v8 ad=2.98155 pd=18.4 as=2.98155 ps=18.4 w=18.07 l=3.61
R0 B.n764 B.n103 585
R1 B.n766 B.n765 585
R2 B.n767 B.n102 585
R3 B.n769 B.n768 585
R4 B.n770 B.n101 585
R5 B.n772 B.n771 585
R6 B.n773 B.n100 585
R7 B.n775 B.n774 585
R8 B.n776 B.n99 585
R9 B.n778 B.n777 585
R10 B.n779 B.n98 585
R11 B.n781 B.n780 585
R12 B.n782 B.n97 585
R13 B.n784 B.n783 585
R14 B.n785 B.n96 585
R15 B.n787 B.n786 585
R16 B.n788 B.n95 585
R17 B.n790 B.n789 585
R18 B.n791 B.n94 585
R19 B.n793 B.n792 585
R20 B.n794 B.n93 585
R21 B.n796 B.n795 585
R22 B.n797 B.n92 585
R23 B.n799 B.n798 585
R24 B.n800 B.n91 585
R25 B.n802 B.n801 585
R26 B.n803 B.n90 585
R27 B.n805 B.n804 585
R28 B.n806 B.n89 585
R29 B.n808 B.n807 585
R30 B.n809 B.n88 585
R31 B.n811 B.n810 585
R32 B.n812 B.n87 585
R33 B.n814 B.n813 585
R34 B.n815 B.n86 585
R35 B.n817 B.n816 585
R36 B.n818 B.n85 585
R37 B.n820 B.n819 585
R38 B.n821 B.n84 585
R39 B.n823 B.n822 585
R40 B.n824 B.n83 585
R41 B.n826 B.n825 585
R42 B.n827 B.n82 585
R43 B.n829 B.n828 585
R44 B.n830 B.n81 585
R45 B.n832 B.n831 585
R46 B.n833 B.n80 585
R47 B.n835 B.n834 585
R48 B.n836 B.n79 585
R49 B.n838 B.n837 585
R50 B.n839 B.n78 585
R51 B.n841 B.n840 585
R52 B.n842 B.n77 585
R53 B.n844 B.n843 585
R54 B.n845 B.n76 585
R55 B.n847 B.n846 585
R56 B.n848 B.n75 585
R57 B.n850 B.n849 585
R58 B.n851 B.n74 585
R59 B.n853 B.n852 585
R60 B.n855 B.n71 585
R61 B.n857 B.n856 585
R62 B.n858 B.n70 585
R63 B.n860 B.n859 585
R64 B.n861 B.n69 585
R65 B.n863 B.n862 585
R66 B.n864 B.n68 585
R67 B.n866 B.n865 585
R68 B.n867 B.n65 585
R69 B.n870 B.n869 585
R70 B.n871 B.n64 585
R71 B.n873 B.n872 585
R72 B.n874 B.n63 585
R73 B.n876 B.n875 585
R74 B.n877 B.n62 585
R75 B.n879 B.n878 585
R76 B.n880 B.n61 585
R77 B.n882 B.n881 585
R78 B.n883 B.n60 585
R79 B.n885 B.n884 585
R80 B.n886 B.n59 585
R81 B.n888 B.n887 585
R82 B.n889 B.n58 585
R83 B.n891 B.n890 585
R84 B.n892 B.n57 585
R85 B.n894 B.n893 585
R86 B.n895 B.n56 585
R87 B.n897 B.n896 585
R88 B.n898 B.n55 585
R89 B.n900 B.n899 585
R90 B.n901 B.n54 585
R91 B.n903 B.n902 585
R92 B.n904 B.n53 585
R93 B.n906 B.n905 585
R94 B.n907 B.n52 585
R95 B.n909 B.n908 585
R96 B.n910 B.n51 585
R97 B.n912 B.n911 585
R98 B.n913 B.n50 585
R99 B.n915 B.n914 585
R100 B.n916 B.n49 585
R101 B.n918 B.n917 585
R102 B.n919 B.n48 585
R103 B.n921 B.n920 585
R104 B.n922 B.n47 585
R105 B.n924 B.n923 585
R106 B.n925 B.n46 585
R107 B.n927 B.n926 585
R108 B.n928 B.n45 585
R109 B.n930 B.n929 585
R110 B.n931 B.n44 585
R111 B.n933 B.n932 585
R112 B.n934 B.n43 585
R113 B.n936 B.n935 585
R114 B.n937 B.n42 585
R115 B.n939 B.n938 585
R116 B.n940 B.n41 585
R117 B.n942 B.n941 585
R118 B.n943 B.n40 585
R119 B.n945 B.n944 585
R120 B.n946 B.n39 585
R121 B.n948 B.n947 585
R122 B.n949 B.n38 585
R123 B.n951 B.n950 585
R124 B.n952 B.n37 585
R125 B.n954 B.n953 585
R126 B.n955 B.n36 585
R127 B.n957 B.n956 585
R128 B.n958 B.n35 585
R129 B.n763 B.n762 585
R130 B.n761 B.n104 585
R131 B.n760 B.n759 585
R132 B.n758 B.n105 585
R133 B.n757 B.n756 585
R134 B.n755 B.n106 585
R135 B.n754 B.n753 585
R136 B.n752 B.n107 585
R137 B.n751 B.n750 585
R138 B.n749 B.n108 585
R139 B.n748 B.n747 585
R140 B.n746 B.n109 585
R141 B.n745 B.n744 585
R142 B.n743 B.n110 585
R143 B.n742 B.n741 585
R144 B.n740 B.n111 585
R145 B.n739 B.n738 585
R146 B.n737 B.n112 585
R147 B.n736 B.n735 585
R148 B.n734 B.n113 585
R149 B.n733 B.n732 585
R150 B.n731 B.n114 585
R151 B.n730 B.n729 585
R152 B.n728 B.n115 585
R153 B.n727 B.n726 585
R154 B.n725 B.n116 585
R155 B.n724 B.n723 585
R156 B.n722 B.n117 585
R157 B.n721 B.n720 585
R158 B.n719 B.n118 585
R159 B.n718 B.n717 585
R160 B.n716 B.n119 585
R161 B.n715 B.n714 585
R162 B.n713 B.n120 585
R163 B.n712 B.n711 585
R164 B.n710 B.n121 585
R165 B.n709 B.n708 585
R166 B.n707 B.n122 585
R167 B.n706 B.n705 585
R168 B.n704 B.n123 585
R169 B.n703 B.n702 585
R170 B.n701 B.n124 585
R171 B.n700 B.n699 585
R172 B.n698 B.n125 585
R173 B.n697 B.n696 585
R174 B.n695 B.n126 585
R175 B.n694 B.n693 585
R176 B.n692 B.n127 585
R177 B.n691 B.n690 585
R178 B.n689 B.n128 585
R179 B.n688 B.n687 585
R180 B.n686 B.n129 585
R181 B.n685 B.n684 585
R182 B.n683 B.n130 585
R183 B.n682 B.n681 585
R184 B.n680 B.n131 585
R185 B.n679 B.n678 585
R186 B.n677 B.n132 585
R187 B.n676 B.n675 585
R188 B.n674 B.n133 585
R189 B.n673 B.n672 585
R190 B.n671 B.n134 585
R191 B.n670 B.n669 585
R192 B.n668 B.n135 585
R193 B.n667 B.n666 585
R194 B.n665 B.n136 585
R195 B.n664 B.n663 585
R196 B.n662 B.n137 585
R197 B.n661 B.n660 585
R198 B.n659 B.n138 585
R199 B.n658 B.n657 585
R200 B.n656 B.n139 585
R201 B.n655 B.n654 585
R202 B.n653 B.n140 585
R203 B.n652 B.n651 585
R204 B.n650 B.n141 585
R205 B.n649 B.n648 585
R206 B.n647 B.n142 585
R207 B.n646 B.n645 585
R208 B.n644 B.n143 585
R209 B.n643 B.n642 585
R210 B.n641 B.n144 585
R211 B.n640 B.n639 585
R212 B.n638 B.n145 585
R213 B.n637 B.n636 585
R214 B.n635 B.n146 585
R215 B.n634 B.n633 585
R216 B.n632 B.n147 585
R217 B.n631 B.n630 585
R218 B.n629 B.n148 585
R219 B.n628 B.n627 585
R220 B.n626 B.n149 585
R221 B.n625 B.n624 585
R222 B.n623 B.n150 585
R223 B.n622 B.n621 585
R224 B.n620 B.n151 585
R225 B.n619 B.n618 585
R226 B.n617 B.n152 585
R227 B.n616 B.n615 585
R228 B.n614 B.n153 585
R229 B.n613 B.n612 585
R230 B.n611 B.n154 585
R231 B.n610 B.n609 585
R232 B.n608 B.n155 585
R233 B.n607 B.n606 585
R234 B.n605 B.n156 585
R235 B.n604 B.n603 585
R236 B.n602 B.n157 585
R237 B.n601 B.n600 585
R238 B.n599 B.n158 585
R239 B.n598 B.n597 585
R240 B.n596 B.n159 585
R241 B.n595 B.n594 585
R242 B.n593 B.n160 585
R243 B.n592 B.n591 585
R244 B.n590 B.n161 585
R245 B.n589 B.n588 585
R246 B.n587 B.n162 585
R247 B.n586 B.n585 585
R248 B.n584 B.n163 585
R249 B.n583 B.n582 585
R250 B.n581 B.n164 585
R251 B.n580 B.n579 585
R252 B.n578 B.n165 585
R253 B.n577 B.n576 585
R254 B.n575 B.n166 585
R255 B.n574 B.n573 585
R256 B.n572 B.n167 585
R257 B.n571 B.n570 585
R258 B.n569 B.n168 585
R259 B.n568 B.n567 585
R260 B.n566 B.n169 585
R261 B.n565 B.n564 585
R262 B.n370 B.n369 585
R263 B.n371 B.n238 585
R264 B.n373 B.n372 585
R265 B.n374 B.n237 585
R266 B.n376 B.n375 585
R267 B.n377 B.n236 585
R268 B.n379 B.n378 585
R269 B.n380 B.n235 585
R270 B.n382 B.n381 585
R271 B.n383 B.n234 585
R272 B.n385 B.n384 585
R273 B.n386 B.n233 585
R274 B.n388 B.n387 585
R275 B.n389 B.n232 585
R276 B.n391 B.n390 585
R277 B.n392 B.n231 585
R278 B.n394 B.n393 585
R279 B.n395 B.n230 585
R280 B.n397 B.n396 585
R281 B.n398 B.n229 585
R282 B.n400 B.n399 585
R283 B.n401 B.n228 585
R284 B.n403 B.n402 585
R285 B.n404 B.n227 585
R286 B.n406 B.n405 585
R287 B.n407 B.n226 585
R288 B.n409 B.n408 585
R289 B.n410 B.n225 585
R290 B.n412 B.n411 585
R291 B.n413 B.n224 585
R292 B.n415 B.n414 585
R293 B.n416 B.n223 585
R294 B.n418 B.n417 585
R295 B.n419 B.n222 585
R296 B.n421 B.n420 585
R297 B.n422 B.n221 585
R298 B.n424 B.n423 585
R299 B.n425 B.n220 585
R300 B.n427 B.n426 585
R301 B.n428 B.n219 585
R302 B.n430 B.n429 585
R303 B.n431 B.n218 585
R304 B.n433 B.n432 585
R305 B.n434 B.n217 585
R306 B.n436 B.n435 585
R307 B.n437 B.n216 585
R308 B.n439 B.n438 585
R309 B.n440 B.n215 585
R310 B.n442 B.n441 585
R311 B.n443 B.n214 585
R312 B.n445 B.n444 585
R313 B.n446 B.n213 585
R314 B.n448 B.n447 585
R315 B.n449 B.n212 585
R316 B.n451 B.n450 585
R317 B.n452 B.n211 585
R318 B.n454 B.n453 585
R319 B.n455 B.n210 585
R320 B.n457 B.n456 585
R321 B.n458 B.n207 585
R322 B.n461 B.n460 585
R323 B.n462 B.n206 585
R324 B.n464 B.n463 585
R325 B.n465 B.n205 585
R326 B.n467 B.n466 585
R327 B.n468 B.n204 585
R328 B.n470 B.n469 585
R329 B.n471 B.n203 585
R330 B.n473 B.n472 585
R331 B.n475 B.n474 585
R332 B.n476 B.n199 585
R333 B.n478 B.n477 585
R334 B.n479 B.n198 585
R335 B.n481 B.n480 585
R336 B.n482 B.n197 585
R337 B.n484 B.n483 585
R338 B.n485 B.n196 585
R339 B.n487 B.n486 585
R340 B.n488 B.n195 585
R341 B.n490 B.n489 585
R342 B.n491 B.n194 585
R343 B.n493 B.n492 585
R344 B.n494 B.n193 585
R345 B.n496 B.n495 585
R346 B.n497 B.n192 585
R347 B.n499 B.n498 585
R348 B.n500 B.n191 585
R349 B.n502 B.n501 585
R350 B.n503 B.n190 585
R351 B.n505 B.n504 585
R352 B.n506 B.n189 585
R353 B.n508 B.n507 585
R354 B.n509 B.n188 585
R355 B.n511 B.n510 585
R356 B.n512 B.n187 585
R357 B.n514 B.n513 585
R358 B.n515 B.n186 585
R359 B.n517 B.n516 585
R360 B.n518 B.n185 585
R361 B.n520 B.n519 585
R362 B.n521 B.n184 585
R363 B.n523 B.n522 585
R364 B.n524 B.n183 585
R365 B.n526 B.n525 585
R366 B.n527 B.n182 585
R367 B.n529 B.n528 585
R368 B.n530 B.n181 585
R369 B.n532 B.n531 585
R370 B.n533 B.n180 585
R371 B.n535 B.n534 585
R372 B.n536 B.n179 585
R373 B.n538 B.n537 585
R374 B.n539 B.n178 585
R375 B.n541 B.n540 585
R376 B.n542 B.n177 585
R377 B.n544 B.n543 585
R378 B.n545 B.n176 585
R379 B.n547 B.n546 585
R380 B.n548 B.n175 585
R381 B.n550 B.n549 585
R382 B.n551 B.n174 585
R383 B.n553 B.n552 585
R384 B.n554 B.n173 585
R385 B.n556 B.n555 585
R386 B.n557 B.n172 585
R387 B.n559 B.n558 585
R388 B.n560 B.n171 585
R389 B.n562 B.n561 585
R390 B.n563 B.n170 585
R391 B.n368 B.n239 585
R392 B.n367 B.n366 585
R393 B.n365 B.n240 585
R394 B.n364 B.n363 585
R395 B.n362 B.n241 585
R396 B.n361 B.n360 585
R397 B.n359 B.n242 585
R398 B.n358 B.n357 585
R399 B.n356 B.n243 585
R400 B.n355 B.n354 585
R401 B.n353 B.n244 585
R402 B.n352 B.n351 585
R403 B.n350 B.n245 585
R404 B.n349 B.n348 585
R405 B.n347 B.n246 585
R406 B.n346 B.n345 585
R407 B.n344 B.n247 585
R408 B.n343 B.n342 585
R409 B.n341 B.n248 585
R410 B.n340 B.n339 585
R411 B.n338 B.n249 585
R412 B.n337 B.n336 585
R413 B.n335 B.n250 585
R414 B.n334 B.n333 585
R415 B.n332 B.n251 585
R416 B.n331 B.n330 585
R417 B.n329 B.n252 585
R418 B.n328 B.n327 585
R419 B.n326 B.n253 585
R420 B.n325 B.n324 585
R421 B.n323 B.n254 585
R422 B.n322 B.n321 585
R423 B.n320 B.n255 585
R424 B.n319 B.n318 585
R425 B.n317 B.n256 585
R426 B.n316 B.n315 585
R427 B.n314 B.n257 585
R428 B.n313 B.n312 585
R429 B.n311 B.n258 585
R430 B.n310 B.n309 585
R431 B.n308 B.n259 585
R432 B.n307 B.n306 585
R433 B.n305 B.n260 585
R434 B.n304 B.n303 585
R435 B.n302 B.n261 585
R436 B.n301 B.n300 585
R437 B.n299 B.n262 585
R438 B.n298 B.n297 585
R439 B.n296 B.n263 585
R440 B.n295 B.n294 585
R441 B.n293 B.n264 585
R442 B.n292 B.n291 585
R443 B.n290 B.n265 585
R444 B.n289 B.n288 585
R445 B.n287 B.n266 585
R446 B.n286 B.n285 585
R447 B.n284 B.n267 585
R448 B.n283 B.n282 585
R449 B.n281 B.n268 585
R450 B.n280 B.n279 585
R451 B.n278 B.n269 585
R452 B.n277 B.n276 585
R453 B.n275 B.n270 585
R454 B.n274 B.n273 585
R455 B.n272 B.n271 585
R456 B.n2 B.n0 585
R457 B.n1057 B.n1 585
R458 B.n1056 B.n1055 585
R459 B.n1054 B.n3 585
R460 B.n1053 B.n1052 585
R461 B.n1051 B.n4 585
R462 B.n1050 B.n1049 585
R463 B.n1048 B.n5 585
R464 B.n1047 B.n1046 585
R465 B.n1045 B.n6 585
R466 B.n1044 B.n1043 585
R467 B.n1042 B.n7 585
R468 B.n1041 B.n1040 585
R469 B.n1039 B.n8 585
R470 B.n1038 B.n1037 585
R471 B.n1036 B.n9 585
R472 B.n1035 B.n1034 585
R473 B.n1033 B.n10 585
R474 B.n1032 B.n1031 585
R475 B.n1030 B.n11 585
R476 B.n1029 B.n1028 585
R477 B.n1027 B.n12 585
R478 B.n1026 B.n1025 585
R479 B.n1024 B.n13 585
R480 B.n1023 B.n1022 585
R481 B.n1021 B.n14 585
R482 B.n1020 B.n1019 585
R483 B.n1018 B.n15 585
R484 B.n1017 B.n1016 585
R485 B.n1015 B.n16 585
R486 B.n1014 B.n1013 585
R487 B.n1012 B.n17 585
R488 B.n1011 B.n1010 585
R489 B.n1009 B.n18 585
R490 B.n1008 B.n1007 585
R491 B.n1006 B.n19 585
R492 B.n1005 B.n1004 585
R493 B.n1003 B.n20 585
R494 B.n1002 B.n1001 585
R495 B.n1000 B.n21 585
R496 B.n999 B.n998 585
R497 B.n997 B.n22 585
R498 B.n996 B.n995 585
R499 B.n994 B.n23 585
R500 B.n993 B.n992 585
R501 B.n991 B.n24 585
R502 B.n990 B.n989 585
R503 B.n988 B.n25 585
R504 B.n987 B.n986 585
R505 B.n985 B.n26 585
R506 B.n984 B.n983 585
R507 B.n982 B.n27 585
R508 B.n981 B.n980 585
R509 B.n979 B.n28 585
R510 B.n978 B.n977 585
R511 B.n976 B.n29 585
R512 B.n975 B.n974 585
R513 B.n973 B.n30 585
R514 B.n972 B.n971 585
R515 B.n970 B.n31 585
R516 B.n969 B.n968 585
R517 B.n967 B.n32 585
R518 B.n966 B.n965 585
R519 B.n964 B.n33 585
R520 B.n963 B.n962 585
R521 B.n961 B.n34 585
R522 B.n960 B.n959 585
R523 B.n1059 B.n1058 585
R524 B.n200 B.t8 561.205
R525 B.n72 B.t10 561.205
R526 B.n208 B.t5 561.203
R527 B.n66 B.t1 561.203
R528 B.n201 B.t7 484.791
R529 B.n73 B.t11 484.791
R530 B.n209 B.t4 484.791
R531 B.n67 B.t2 484.791
R532 B.n370 B.n239 468.476
R533 B.n960 B.n35 468.476
R534 B.n564 B.n563 468.476
R535 B.n762 B.n103 468.476
R536 B.n200 B.t6 329.824
R537 B.n208 B.t3 329.824
R538 B.n66 B.t0 329.824
R539 B.n72 B.t9 329.824
R540 B.n366 B.n239 163.367
R541 B.n366 B.n365 163.367
R542 B.n365 B.n364 163.367
R543 B.n364 B.n241 163.367
R544 B.n360 B.n241 163.367
R545 B.n360 B.n359 163.367
R546 B.n359 B.n358 163.367
R547 B.n358 B.n243 163.367
R548 B.n354 B.n243 163.367
R549 B.n354 B.n353 163.367
R550 B.n353 B.n352 163.367
R551 B.n352 B.n245 163.367
R552 B.n348 B.n245 163.367
R553 B.n348 B.n347 163.367
R554 B.n347 B.n346 163.367
R555 B.n346 B.n247 163.367
R556 B.n342 B.n247 163.367
R557 B.n342 B.n341 163.367
R558 B.n341 B.n340 163.367
R559 B.n340 B.n249 163.367
R560 B.n336 B.n249 163.367
R561 B.n336 B.n335 163.367
R562 B.n335 B.n334 163.367
R563 B.n334 B.n251 163.367
R564 B.n330 B.n251 163.367
R565 B.n330 B.n329 163.367
R566 B.n329 B.n328 163.367
R567 B.n328 B.n253 163.367
R568 B.n324 B.n253 163.367
R569 B.n324 B.n323 163.367
R570 B.n323 B.n322 163.367
R571 B.n322 B.n255 163.367
R572 B.n318 B.n255 163.367
R573 B.n318 B.n317 163.367
R574 B.n317 B.n316 163.367
R575 B.n316 B.n257 163.367
R576 B.n312 B.n257 163.367
R577 B.n312 B.n311 163.367
R578 B.n311 B.n310 163.367
R579 B.n310 B.n259 163.367
R580 B.n306 B.n259 163.367
R581 B.n306 B.n305 163.367
R582 B.n305 B.n304 163.367
R583 B.n304 B.n261 163.367
R584 B.n300 B.n261 163.367
R585 B.n300 B.n299 163.367
R586 B.n299 B.n298 163.367
R587 B.n298 B.n263 163.367
R588 B.n294 B.n263 163.367
R589 B.n294 B.n293 163.367
R590 B.n293 B.n292 163.367
R591 B.n292 B.n265 163.367
R592 B.n288 B.n265 163.367
R593 B.n288 B.n287 163.367
R594 B.n287 B.n286 163.367
R595 B.n286 B.n267 163.367
R596 B.n282 B.n267 163.367
R597 B.n282 B.n281 163.367
R598 B.n281 B.n280 163.367
R599 B.n280 B.n269 163.367
R600 B.n276 B.n269 163.367
R601 B.n276 B.n275 163.367
R602 B.n275 B.n274 163.367
R603 B.n274 B.n271 163.367
R604 B.n271 B.n2 163.367
R605 B.n1058 B.n2 163.367
R606 B.n1058 B.n1057 163.367
R607 B.n1057 B.n1056 163.367
R608 B.n1056 B.n3 163.367
R609 B.n1052 B.n3 163.367
R610 B.n1052 B.n1051 163.367
R611 B.n1051 B.n1050 163.367
R612 B.n1050 B.n5 163.367
R613 B.n1046 B.n5 163.367
R614 B.n1046 B.n1045 163.367
R615 B.n1045 B.n1044 163.367
R616 B.n1044 B.n7 163.367
R617 B.n1040 B.n7 163.367
R618 B.n1040 B.n1039 163.367
R619 B.n1039 B.n1038 163.367
R620 B.n1038 B.n9 163.367
R621 B.n1034 B.n9 163.367
R622 B.n1034 B.n1033 163.367
R623 B.n1033 B.n1032 163.367
R624 B.n1032 B.n11 163.367
R625 B.n1028 B.n11 163.367
R626 B.n1028 B.n1027 163.367
R627 B.n1027 B.n1026 163.367
R628 B.n1026 B.n13 163.367
R629 B.n1022 B.n13 163.367
R630 B.n1022 B.n1021 163.367
R631 B.n1021 B.n1020 163.367
R632 B.n1020 B.n15 163.367
R633 B.n1016 B.n15 163.367
R634 B.n1016 B.n1015 163.367
R635 B.n1015 B.n1014 163.367
R636 B.n1014 B.n17 163.367
R637 B.n1010 B.n17 163.367
R638 B.n1010 B.n1009 163.367
R639 B.n1009 B.n1008 163.367
R640 B.n1008 B.n19 163.367
R641 B.n1004 B.n19 163.367
R642 B.n1004 B.n1003 163.367
R643 B.n1003 B.n1002 163.367
R644 B.n1002 B.n21 163.367
R645 B.n998 B.n21 163.367
R646 B.n998 B.n997 163.367
R647 B.n997 B.n996 163.367
R648 B.n996 B.n23 163.367
R649 B.n992 B.n23 163.367
R650 B.n992 B.n991 163.367
R651 B.n991 B.n990 163.367
R652 B.n990 B.n25 163.367
R653 B.n986 B.n25 163.367
R654 B.n986 B.n985 163.367
R655 B.n985 B.n984 163.367
R656 B.n984 B.n27 163.367
R657 B.n980 B.n27 163.367
R658 B.n980 B.n979 163.367
R659 B.n979 B.n978 163.367
R660 B.n978 B.n29 163.367
R661 B.n974 B.n29 163.367
R662 B.n974 B.n973 163.367
R663 B.n973 B.n972 163.367
R664 B.n972 B.n31 163.367
R665 B.n968 B.n31 163.367
R666 B.n968 B.n967 163.367
R667 B.n967 B.n966 163.367
R668 B.n966 B.n33 163.367
R669 B.n962 B.n33 163.367
R670 B.n962 B.n961 163.367
R671 B.n961 B.n960 163.367
R672 B.n371 B.n370 163.367
R673 B.n372 B.n371 163.367
R674 B.n372 B.n237 163.367
R675 B.n376 B.n237 163.367
R676 B.n377 B.n376 163.367
R677 B.n378 B.n377 163.367
R678 B.n378 B.n235 163.367
R679 B.n382 B.n235 163.367
R680 B.n383 B.n382 163.367
R681 B.n384 B.n383 163.367
R682 B.n384 B.n233 163.367
R683 B.n388 B.n233 163.367
R684 B.n389 B.n388 163.367
R685 B.n390 B.n389 163.367
R686 B.n390 B.n231 163.367
R687 B.n394 B.n231 163.367
R688 B.n395 B.n394 163.367
R689 B.n396 B.n395 163.367
R690 B.n396 B.n229 163.367
R691 B.n400 B.n229 163.367
R692 B.n401 B.n400 163.367
R693 B.n402 B.n401 163.367
R694 B.n402 B.n227 163.367
R695 B.n406 B.n227 163.367
R696 B.n407 B.n406 163.367
R697 B.n408 B.n407 163.367
R698 B.n408 B.n225 163.367
R699 B.n412 B.n225 163.367
R700 B.n413 B.n412 163.367
R701 B.n414 B.n413 163.367
R702 B.n414 B.n223 163.367
R703 B.n418 B.n223 163.367
R704 B.n419 B.n418 163.367
R705 B.n420 B.n419 163.367
R706 B.n420 B.n221 163.367
R707 B.n424 B.n221 163.367
R708 B.n425 B.n424 163.367
R709 B.n426 B.n425 163.367
R710 B.n426 B.n219 163.367
R711 B.n430 B.n219 163.367
R712 B.n431 B.n430 163.367
R713 B.n432 B.n431 163.367
R714 B.n432 B.n217 163.367
R715 B.n436 B.n217 163.367
R716 B.n437 B.n436 163.367
R717 B.n438 B.n437 163.367
R718 B.n438 B.n215 163.367
R719 B.n442 B.n215 163.367
R720 B.n443 B.n442 163.367
R721 B.n444 B.n443 163.367
R722 B.n444 B.n213 163.367
R723 B.n448 B.n213 163.367
R724 B.n449 B.n448 163.367
R725 B.n450 B.n449 163.367
R726 B.n450 B.n211 163.367
R727 B.n454 B.n211 163.367
R728 B.n455 B.n454 163.367
R729 B.n456 B.n455 163.367
R730 B.n456 B.n207 163.367
R731 B.n461 B.n207 163.367
R732 B.n462 B.n461 163.367
R733 B.n463 B.n462 163.367
R734 B.n463 B.n205 163.367
R735 B.n467 B.n205 163.367
R736 B.n468 B.n467 163.367
R737 B.n469 B.n468 163.367
R738 B.n469 B.n203 163.367
R739 B.n473 B.n203 163.367
R740 B.n474 B.n473 163.367
R741 B.n474 B.n199 163.367
R742 B.n478 B.n199 163.367
R743 B.n479 B.n478 163.367
R744 B.n480 B.n479 163.367
R745 B.n480 B.n197 163.367
R746 B.n484 B.n197 163.367
R747 B.n485 B.n484 163.367
R748 B.n486 B.n485 163.367
R749 B.n486 B.n195 163.367
R750 B.n490 B.n195 163.367
R751 B.n491 B.n490 163.367
R752 B.n492 B.n491 163.367
R753 B.n492 B.n193 163.367
R754 B.n496 B.n193 163.367
R755 B.n497 B.n496 163.367
R756 B.n498 B.n497 163.367
R757 B.n498 B.n191 163.367
R758 B.n502 B.n191 163.367
R759 B.n503 B.n502 163.367
R760 B.n504 B.n503 163.367
R761 B.n504 B.n189 163.367
R762 B.n508 B.n189 163.367
R763 B.n509 B.n508 163.367
R764 B.n510 B.n509 163.367
R765 B.n510 B.n187 163.367
R766 B.n514 B.n187 163.367
R767 B.n515 B.n514 163.367
R768 B.n516 B.n515 163.367
R769 B.n516 B.n185 163.367
R770 B.n520 B.n185 163.367
R771 B.n521 B.n520 163.367
R772 B.n522 B.n521 163.367
R773 B.n522 B.n183 163.367
R774 B.n526 B.n183 163.367
R775 B.n527 B.n526 163.367
R776 B.n528 B.n527 163.367
R777 B.n528 B.n181 163.367
R778 B.n532 B.n181 163.367
R779 B.n533 B.n532 163.367
R780 B.n534 B.n533 163.367
R781 B.n534 B.n179 163.367
R782 B.n538 B.n179 163.367
R783 B.n539 B.n538 163.367
R784 B.n540 B.n539 163.367
R785 B.n540 B.n177 163.367
R786 B.n544 B.n177 163.367
R787 B.n545 B.n544 163.367
R788 B.n546 B.n545 163.367
R789 B.n546 B.n175 163.367
R790 B.n550 B.n175 163.367
R791 B.n551 B.n550 163.367
R792 B.n552 B.n551 163.367
R793 B.n552 B.n173 163.367
R794 B.n556 B.n173 163.367
R795 B.n557 B.n556 163.367
R796 B.n558 B.n557 163.367
R797 B.n558 B.n171 163.367
R798 B.n562 B.n171 163.367
R799 B.n563 B.n562 163.367
R800 B.n564 B.n169 163.367
R801 B.n568 B.n169 163.367
R802 B.n569 B.n568 163.367
R803 B.n570 B.n569 163.367
R804 B.n570 B.n167 163.367
R805 B.n574 B.n167 163.367
R806 B.n575 B.n574 163.367
R807 B.n576 B.n575 163.367
R808 B.n576 B.n165 163.367
R809 B.n580 B.n165 163.367
R810 B.n581 B.n580 163.367
R811 B.n582 B.n581 163.367
R812 B.n582 B.n163 163.367
R813 B.n586 B.n163 163.367
R814 B.n587 B.n586 163.367
R815 B.n588 B.n587 163.367
R816 B.n588 B.n161 163.367
R817 B.n592 B.n161 163.367
R818 B.n593 B.n592 163.367
R819 B.n594 B.n593 163.367
R820 B.n594 B.n159 163.367
R821 B.n598 B.n159 163.367
R822 B.n599 B.n598 163.367
R823 B.n600 B.n599 163.367
R824 B.n600 B.n157 163.367
R825 B.n604 B.n157 163.367
R826 B.n605 B.n604 163.367
R827 B.n606 B.n605 163.367
R828 B.n606 B.n155 163.367
R829 B.n610 B.n155 163.367
R830 B.n611 B.n610 163.367
R831 B.n612 B.n611 163.367
R832 B.n612 B.n153 163.367
R833 B.n616 B.n153 163.367
R834 B.n617 B.n616 163.367
R835 B.n618 B.n617 163.367
R836 B.n618 B.n151 163.367
R837 B.n622 B.n151 163.367
R838 B.n623 B.n622 163.367
R839 B.n624 B.n623 163.367
R840 B.n624 B.n149 163.367
R841 B.n628 B.n149 163.367
R842 B.n629 B.n628 163.367
R843 B.n630 B.n629 163.367
R844 B.n630 B.n147 163.367
R845 B.n634 B.n147 163.367
R846 B.n635 B.n634 163.367
R847 B.n636 B.n635 163.367
R848 B.n636 B.n145 163.367
R849 B.n640 B.n145 163.367
R850 B.n641 B.n640 163.367
R851 B.n642 B.n641 163.367
R852 B.n642 B.n143 163.367
R853 B.n646 B.n143 163.367
R854 B.n647 B.n646 163.367
R855 B.n648 B.n647 163.367
R856 B.n648 B.n141 163.367
R857 B.n652 B.n141 163.367
R858 B.n653 B.n652 163.367
R859 B.n654 B.n653 163.367
R860 B.n654 B.n139 163.367
R861 B.n658 B.n139 163.367
R862 B.n659 B.n658 163.367
R863 B.n660 B.n659 163.367
R864 B.n660 B.n137 163.367
R865 B.n664 B.n137 163.367
R866 B.n665 B.n664 163.367
R867 B.n666 B.n665 163.367
R868 B.n666 B.n135 163.367
R869 B.n670 B.n135 163.367
R870 B.n671 B.n670 163.367
R871 B.n672 B.n671 163.367
R872 B.n672 B.n133 163.367
R873 B.n676 B.n133 163.367
R874 B.n677 B.n676 163.367
R875 B.n678 B.n677 163.367
R876 B.n678 B.n131 163.367
R877 B.n682 B.n131 163.367
R878 B.n683 B.n682 163.367
R879 B.n684 B.n683 163.367
R880 B.n684 B.n129 163.367
R881 B.n688 B.n129 163.367
R882 B.n689 B.n688 163.367
R883 B.n690 B.n689 163.367
R884 B.n690 B.n127 163.367
R885 B.n694 B.n127 163.367
R886 B.n695 B.n694 163.367
R887 B.n696 B.n695 163.367
R888 B.n696 B.n125 163.367
R889 B.n700 B.n125 163.367
R890 B.n701 B.n700 163.367
R891 B.n702 B.n701 163.367
R892 B.n702 B.n123 163.367
R893 B.n706 B.n123 163.367
R894 B.n707 B.n706 163.367
R895 B.n708 B.n707 163.367
R896 B.n708 B.n121 163.367
R897 B.n712 B.n121 163.367
R898 B.n713 B.n712 163.367
R899 B.n714 B.n713 163.367
R900 B.n714 B.n119 163.367
R901 B.n718 B.n119 163.367
R902 B.n719 B.n718 163.367
R903 B.n720 B.n719 163.367
R904 B.n720 B.n117 163.367
R905 B.n724 B.n117 163.367
R906 B.n725 B.n724 163.367
R907 B.n726 B.n725 163.367
R908 B.n726 B.n115 163.367
R909 B.n730 B.n115 163.367
R910 B.n731 B.n730 163.367
R911 B.n732 B.n731 163.367
R912 B.n732 B.n113 163.367
R913 B.n736 B.n113 163.367
R914 B.n737 B.n736 163.367
R915 B.n738 B.n737 163.367
R916 B.n738 B.n111 163.367
R917 B.n742 B.n111 163.367
R918 B.n743 B.n742 163.367
R919 B.n744 B.n743 163.367
R920 B.n744 B.n109 163.367
R921 B.n748 B.n109 163.367
R922 B.n749 B.n748 163.367
R923 B.n750 B.n749 163.367
R924 B.n750 B.n107 163.367
R925 B.n754 B.n107 163.367
R926 B.n755 B.n754 163.367
R927 B.n756 B.n755 163.367
R928 B.n756 B.n105 163.367
R929 B.n760 B.n105 163.367
R930 B.n761 B.n760 163.367
R931 B.n762 B.n761 163.367
R932 B.n956 B.n35 163.367
R933 B.n956 B.n955 163.367
R934 B.n955 B.n954 163.367
R935 B.n954 B.n37 163.367
R936 B.n950 B.n37 163.367
R937 B.n950 B.n949 163.367
R938 B.n949 B.n948 163.367
R939 B.n948 B.n39 163.367
R940 B.n944 B.n39 163.367
R941 B.n944 B.n943 163.367
R942 B.n943 B.n942 163.367
R943 B.n942 B.n41 163.367
R944 B.n938 B.n41 163.367
R945 B.n938 B.n937 163.367
R946 B.n937 B.n936 163.367
R947 B.n936 B.n43 163.367
R948 B.n932 B.n43 163.367
R949 B.n932 B.n931 163.367
R950 B.n931 B.n930 163.367
R951 B.n930 B.n45 163.367
R952 B.n926 B.n45 163.367
R953 B.n926 B.n925 163.367
R954 B.n925 B.n924 163.367
R955 B.n924 B.n47 163.367
R956 B.n920 B.n47 163.367
R957 B.n920 B.n919 163.367
R958 B.n919 B.n918 163.367
R959 B.n918 B.n49 163.367
R960 B.n914 B.n49 163.367
R961 B.n914 B.n913 163.367
R962 B.n913 B.n912 163.367
R963 B.n912 B.n51 163.367
R964 B.n908 B.n51 163.367
R965 B.n908 B.n907 163.367
R966 B.n907 B.n906 163.367
R967 B.n906 B.n53 163.367
R968 B.n902 B.n53 163.367
R969 B.n902 B.n901 163.367
R970 B.n901 B.n900 163.367
R971 B.n900 B.n55 163.367
R972 B.n896 B.n55 163.367
R973 B.n896 B.n895 163.367
R974 B.n895 B.n894 163.367
R975 B.n894 B.n57 163.367
R976 B.n890 B.n57 163.367
R977 B.n890 B.n889 163.367
R978 B.n889 B.n888 163.367
R979 B.n888 B.n59 163.367
R980 B.n884 B.n59 163.367
R981 B.n884 B.n883 163.367
R982 B.n883 B.n882 163.367
R983 B.n882 B.n61 163.367
R984 B.n878 B.n61 163.367
R985 B.n878 B.n877 163.367
R986 B.n877 B.n876 163.367
R987 B.n876 B.n63 163.367
R988 B.n872 B.n63 163.367
R989 B.n872 B.n871 163.367
R990 B.n871 B.n870 163.367
R991 B.n870 B.n65 163.367
R992 B.n865 B.n65 163.367
R993 B.n865 B.n864 163.367
R994 B.n864 B.n863 163.367
R995 B.n863 B.n69 163.367
R996 B.n859 B.n69 163.367
R997 B.n859 B.n858 163.367
R998 B.n858 B.n857 163.367
R999 B.n857 B.n71 163.367
R1000 B.n852 B.n71 163.367
R1001 B.n852 B.n851 163.367
R1002 B.n851 B.n850 163.367
R1003 B.n850 B.n75 163.367
R1004 B.n846 B.n75 163.367
R1005 B.n846 B.n845 163.367
R1006 B.n845 B.n844 163.367
R1007 B.n844 B.n77 163.367
R1008 B.n840 B.n77 163.367
R1009 B.n840 B.n839 163.367
R1010 B.n839 B.n838 163.367
R1011 B.n838 B.n79 163.367
R1012 B.n834 B.n79 163.367
R1013 B.n834 B.n833 163.367
R1014 B.n833 B.n832 163.367
R1015 B.n832 B.n81 163.367
R1016 B.n828 B.n81 163.367
R1017 B.n828 B.n827 163.367
R1018 B.n827 B.n826 163.367
R1019 B.n826 B.n83 163.367
R1020 B.n822 B.n83 163.367
R1021 B.n822 B.n821 163.367
R1022 B.n821 B.n820 163.367
R1023 B.n820 B.n85 163.367
R1024 B.n816 B.n85 163.367
R1025 B.n816 B.n815 163.367
R1026 B.n815 B.n814 163.367
R1027 B.n814 B.n87 163.367
R1028 B.n810 B.n87 163.367
R1029 B.n810 B.n809 163.367
R1030 B.n809 B.n808 163.367
R1031 B.n808 B.n89 163.367
R1032 B.n804 B.n89 163.367
R1033 B.n804 B.n803 163.367
R1034 B.n803 B.n802 163.367
R1035 B.n802 B.n91 163.367
R1036 B.n798 B.n91 163.367
R1037 B.n798 B.n797 163.367
R1038 B.n797 B.n796 163.367
R1039 B.n796 B.n93 163.367
R1040 B.n792 B.n93 163.367
R1041 B.n792 B.n791 163.367
R1042 B.n791 B.n790 163.367
R1043 B.n790 B.n95 163.367
R1044 B.n786 B.n95 163.367
R1045 B.n786 B.n785 163.367
R1046 B.n785 B.n784 163.367
R1047 B.n784 B.n97 163.367
R1048 B.n780 B.n97 163.367
R1049 B.n780 B.n779 163.367
R1050 B.n779 B.n778 163.367
R1051 B.n778 B.n99 163.367
R1052 B.n774 B.n99 163.367
R1053 B.n774 B.n773 163.367
R1054 B.n773 B.n772 163.367
R1055 B.n772 B.n101 163.367
R1056 B.n768 B.n101 163.367
R1057 B.n768 B.n767 163.367
R1058 B.n767 B.n766 163.367
R1059 B.n766 B.n103 163.367
R1060 B.n201 B.n200 76.4126
R1061 B.n209 B.n208 76.4126
R1062 B.n67 B.n66 76.4126
R1063 B.n73 B.n72 76.4126
R1064 B.n202 B.n201 59.5399
R1065 B.n459 B.n209 59.5399
R1066 B.n868 B.n67 59.5399
R1067 B.n854 B.n73 59.5399
R1068 B.n764 B.n763 30.4395
R1069 B.n959 B.n958 30.4395
R1070 B.n565 B.n170 30.4395
R1071 B.n369 B.n368 30.4395
R1072 B B.n1059 18.0485
R1073 B.n958 B.n957 10.6151
R1074 B.n957 B.n36 10.6151
R1075 B.n953 B.n36 10.6151
R1076 B.n953 B.n952 10.6151
R1077 B.n952 B.n951 10.6151
R1078 B.n951 B.n38 10.6151
R1079 B.n947 B.n38 10.6151
R1080 B.n947 B.n946 10.6151
R1081 B.n946 B.n945 10.6151
R1082 B.n945 B.n40 10.6151
R1083 B.n941 B.n40 10.6151
R1084 B.n941 B.n940 10.6151
R1085 B.n940 B.n939 10.6151
R1086 B.n939 B.n42 10.6151
R1087 B.n935 B.n42 10.6151
R1088 B.n935 B.n934 10.6151
R1089 B.n934 B.n933 10.6151
R1090 B.n933 B.n44 10.6151
R1091 B.n929 B.n44 10.6151
R1092 B.n929 B.n928 10.6151
R1093 B.n928 B.n927 10.6151
R1094 B.n927 B.n46 10.6151
R1095 B.n923 B.n46 10.6151
R1096 B.n923 B.n922 10.6151
R1097 B.n922 B.n921 10.6151
R1098 B.n921 B.n48 10.6151
R1099 B.n917 B.n48 10.6151
R1100 B.n917 B.n916 10.6151
R1101 B.n916 B.n915 10.6151
R1102 B.n915 B.n50 10.6151
R1103 B.n911 B.n50 10.6151
R1104 B.n911 B.n910 10.6151
R1105 B.n910 B.n909 10.6151
R1106 B.n909 B.n52 10.6151
R1107 B.n905 B.n52 10.6151
R1108 B.n905 B.n904 10.6151
R1109 B.n904 B.n903 10.6151
R1110 B.n903 B.n54 10.6151
R1111 B.n899 B.n54 10.6151
R1112 B.n899 B.n898 10.6151
R1113 B.n898 B.n897 10.6151
R1114 B.n897 B.n56 10.6151
R1115 B.n893 B.n56 10.6151
R1116 B.n893 B.n892 10.6151
R1117 B.n892 B.n891 10.6151
R1118 B.n891 B.n58 10.6151
R1119 B.n887 B.n58 10.6151
R1120 B.n887 B.n886 10.6151
R1121 B.n886 B.n885 10.6151
R1122 B.n885 B.n60 10.6151
R1123 B.n881 B.n60 10.6151
R1124 B.n881 B.n880 10.6151
R1125 B.n880 B.n879 10.6151
R1126 B.n879 B.n62 10.6151
R1127 B.n875 B.n62 10.6151
R1128 B.n875 B.n874 10.6151
R1129 B.n874 B.n873 10.6151
R1130 B.n873 B.n64 10.6151
R1131 B.n869 B.n64 10.6151
R1132 B.n867 B.n866 10.6151
R1133 B.n866 B.n68 10.6151
R1134 B.n862 B.n68 10.6151
R1135 B.n862 B.n861 10.6151
R1136 B.n861 B.n860 10.6151
R1137 B.n860 B.n70 10.6151
R1138 B.n856 B.n70 10.6151
R1139 B.n856 B.n855 10.6151
R1140 B.n853 B.n74 10.6151
R1141 B.n849 B.n74 10.6151
R1142 B.n849 B.n848 10.6151
R1143 B.n848 B.n847 10.6151
R1144 B.n847 B.n76 10.6151
R1145 B.n843 B.n76 10.6151
R1146 B.n843 B.n842 10.6151
R1147 B.n842 B.n841 10.6151
R1148 B.n841 B.n78 10.6151
R1149 B.n837 B.n78 10.6151
R1150 B.n837 B.n836 10.6151
R1151 B.n836 B.n835 10.6151
R1152 B.n835 B.n80 10.6151
R1153 B.n831 B.n80 10.6151
R1154 B.n831 B.n830 10.6151
R1155 B.n830 B.n829 10.6151
R1156 B.n829 B.n82 10.6151
R1157 B.n825 B.n82 10.6151
R1158 B.n825 B.n824 10.6151
R1159 B.n824 B.n823 10.6151
R1160 B.n823 B.n84 10.6151
R1161 B.n819 B.n84 10.6151
R1162 B.n819 B.n818 10.6151
R1163 B.n818 B.n817 10.6151
R1164 B.n817 B.n86 10.6151
R1165 B.n813 B.n86 10.6151
R1166 B.n813 B.n812 10.6151
R1167 B.n812 B.n811 10.6151
R1168 B.n811 B.n88 10.6151
R1169 B.n807 B.n88 10.6151
R1170 B.n807 B.n806 10.6151
R1171 B.n806 B.n805 10.6151
R1172 B.n805 B.n90 10.6151
R1173 B.n801 B.n90 10.6151
R1174 B.n801 B.n800 10.6151
R1175 B.n800 B.n799 10.6151
R1176 B.n799 B.n92 10.6151
R1177 B.n795 B.n92 10.6151
R1178 B.n795 B.n794 10.6151
R1179 B.n794 B.n793 10.6151
R1180 B.n793 B.n94 10.6151
R1181 B.n789 B.n94 10.6151
R1182 B.n789 B.n788 10.6151
R1183 B.n788 B.n787 10.6151
R1184 B.n787 B.n96 10.6151
R1185 B.n783 B.n96 10.6151
R1186 B.n783 B.n782 10.6151
R1187 B.n782 B.n781 10.6151
R1188 B.n781 B.n98 10.6151
R1189 B.n777 B.n98 10.6151
R1190 B.n777 B.n776 10.6151
R1191 B.n776 B.n775 10.6151
R1192 B.n775 B.n100 10.6151
R1193 B.n771 B.n100 10.6151
R1194 B.n771 B.n770 10.6151
R1195 B.n770 B.n769 10.6151
R1196 B.n769 B.n102 10.6151
R1197 B.n765 B.n102 10.6151
R1198 B.n765 B.n764 10.6151
R1199 B.n566 B.n565 10.6151
R1200 B.n567 B.n566 10.6151
R1201 B.n567 B.n168 10.6151
R1202 B.n571 B.n168 10.6151
R1203 B.n572 B.n571 10.6151
R1204 B.n573 B.n572 10.6151
R1205 B.n573 B.n166 10.6151
R1206 B.n577 B.n166 10.6151
R1207 B.n578 B.n577 10.6151
R1208 B.n579 B.n578 10.6151
R1209 B.n579 B.n164 10.6151
R1210 B.n583 B.n164 10.6151
R1211 B.n584 B.n583 10.6151
R1212 B.n585 B.n584 10.6151
R1213 B.n585 B.n162 10.6151
R1214 B.n589 B.n162 10.6151
R1215 B.n590 B.n589 10.6151
R1216 B.n591 B.n590 10.6151
R1217 B.n591 B.n160 10.6151
R1218 B.n595 B.n160 10.6151
R1219 B.n596 B.n595 10.6151
R1220 B.n597 B.n596 10.6151
R1221 B.n597 B.n158 10.6151
R1222 B.n601 B.n158 10.6151
R1223 B.n602 B.n601 10.6151
R1224 B.n603 B.n602 10.6151
R1225 B.n603 B.n156 10.6151
R1226 B.n607 B.n156 10.6151
R1227 B.n608 B.n607 10.6151
R1228 B.n609 B.n608 10.6151
R1229 B.n609 B.n154 10.6151
R1230 B.n613 B.n154 10.6151
R1231 B.n614 B.n613 10.6151
R1232 B.n615 B.n614 10.6151
R1233 B.n615 B.n152 10.6151
R1234 B.n619 B.n152 10.6151
R1235 B.n620 B.n619 10.6151
R1236 B.n621 B.n620 10.6151
R1237 B.n621 B.n150 10.6151
R1238 B.n625 B.n150 10.6151
R1239 B.n626 B.n625 10.6151
R1240 B.n627 B.n626 10.6151
R1241 B.n627 B.n148 10.6151
R1242 B.n631 B.n148 10.6151
R1243 B.n632 B.n631 10.6151
R1244 B.n633 B.n632 10.6151
R1245 B.n633 B.n146 10.6151
R1246 B.n637 B.n146 10.6151
R1247 B.n638 B.n637 10.6151
R1248 B.n639 B.n638 10.6151
R1249 B.n639 B.n144 10.6151
R1250 B.n643 B.n144 10.6151
R1251 B.n644 B.n643 10.6151
R1252 B.n645 B.n644 10.6151
R1253 B.n645 B.n142 10.6151
R1254 B.n649 B.n142 10.6151
R1255 B.n650 B.n649 10.6151
R1256 B.n651 B.n650 10.6151
R1257 B.n651 B.n140 10.6151
R1258 B.n655 B.n140 10.6151
R1259 B.n656 B.n655 10.6151
R1260 B.n657 B.n656 10.6151
R1261 B.n657 B.n138 10.6151
R1262 B.n661 B.n138 10.6151
R1263 B.n662 B.n661 10.6151
R1264 B.n663 B.n662 10.6151
R1265 B.n663 B.n136 10.6151
R1266 B.n667 B.n136 10.6151
R1267 B.n668 B.n667 10.6151
R1268 B.n669 B.n668 10.6151
R1269 B.n669 B.n134 10.6151
R1270 B.n673 B.n134 10.6151
R1271 B.n674 B.n673 10.6151
R1272 B.n675 B.n674 10.6151
R1273 B.n675 B.n132 10.6151
R1274 B.n679 B.n132 10.6151
R1275 B.n680 B.n679 10.6151
R1276 B.n681 B.n680 10.6151
R1277 B.n681 B.n130 10.6151
R1278 B.n685 B.n130 10.6151
R1279 B.n686 B.n685 10.6151
R1280 B.n687 B.n686 10.6151
R1281 B.n687 B.n128 10.6151
R1282 B.n691 B.n128 10.6151
R1283 B.n692 B.n691 10.6151
R1284 B.n693 B.n692 10.6151
R1285 B.n693 B.n126 10.6151
R1286 B.n697 B.n126 10.6151
R1287 B.n698 B.n697 10.6151
R1288 B.n699 B.n698 10.6151
R1289 B.n699 B.n124 10.6151
R1290 B.n703 B.n124 10.6151
R1291 B.n704 B.n703 10.6151
R1292 B.n705 B.n704 10.6151
R1293 B.n705 B.n122 10.6151
R1294 B.n709 B.n122 10.6151
R1295 B.n710 B.n709 10.6151
R1296 B.n711 B.n710 10.6151
R1297 B.n711 B.n120 10.6151
R1298 B.n715 B.n120 10.6151
R1299 B.n716 B.n715 10.6151
R1300 B.n717 B.n716 10.6151
R1301 B.n717 B.n118 10.6151
R1302 B.n721 B.n118 10.6151
R1303 B.n722 B.n721 10.6151
R1304 B.n723 B.n722 10.6151
R1305 B.n723 B.n116 10.6151
R1306 B.n727 B.n116 10.6151
R1307 B.n728 B.n727 10.6151
R1308 B.n729 B.n728 10.6151
R1309 B.n729 B.n114 10.6151
R1310 B.n733 B.n114 10.6151
R1311 B.n734 B.n733 10.6151
R1312 B.n735 B.n734 10.6151
R1313 B.n735 B.n112 10.6151
R1314 B.n739 B.n112 10.6151
R1315 B.n740 B.n739 10.6151
R1316 B.n741 B.n740 10.6151
R1317 B.n741 B.n110 10.6151
R1318 B.n745 B.n110 10.6151
R1319 B.n746 B.n745 10.6151
R1320 B.n747 B.n746 10.6151
R1321 B.n747 B.n108 10.6151
R1322 B.n751 B.n108 10.6151
R1323 B.n752 B.n751 10.6151
R1324 B.n753 B.n752 10.6151
R1325 B.n753 B.n106 10.6151
R1326 B.n757 B.n106 10.6151
R1327 B.n758 B.n757 10.6151
R1328 B.n759 B.n758 10.6151
R1329 B.n759 B.n104 10.6151
R1330 B.n763 B.n104 10.6151
R1331 B.n369 B.n238 10.6151
R1332 B.n373 B.n238 10.6151
R1333 B.n374 B.n373 10.6151
R1334 B.n375 B.n374 10.6151
R1335 B.n375 B.n236 10.6151
R1336 B.n379 B.n236 10.6151
R1337 B.n380 B.n379 10.6151
R1338 B.n381 B.n380 10.6151
R1339 B.n381 B.n234 10.6151
R1340 B.n385 B.n234 10.6151
R1341 B.n386 B.n385 10.6151
R1342 B.n387 B.n386 10.6151
R1343 B.n387 B.n232 10.6151
R1344 B.n391 B.n232 10.6151
R1345 B.n392 B.n391 10.6151
R1346 B.n393 B.n392 10.6151
R1347 B.n393 B.n230 10.6151
R1348 B.n397 B.n230 10.6151
R1349 B.n398 B.n397 10.6151
R1350 B.n399 B.n398 10.6151
R1351 B.n399 B.n228 10.6151
R1352 B.n403 B.n228 10.6151
R1353 B.n404 B.n403 10.6151
R1354 B.n405 B.n404 10.6151
R1355 B.n405 B.n226 10.6151
R1356 B.n409 B.n226 10.6151
R1357 B.n410 B.n409 10.6151
R1358 B.n411 B.n410 10.6151
R1359 B.n411 B.n224 10.6151
R1360 B.n415 B.n224 10.6151
R1361 B.n416 B.n415 10.6151
R1362 B.n417 B.n416 10.6151
R1363 B.n417 B.n222 10.6151
R1364 B.n421 B.n222 10.6151
R1365 B.n422 B.n421 10.6151
R1366 B.n423 B.n422 10.6151
R1367 B.n423 B.n220 10.6151
R1368 B.n427 B.n220 10.6151
R1369 B.n428 B.n427 10.6151
R1370 B.n429 B.n428 10.6151
R1371 B.n429 B.n218 10.6151
R1372 B.n433 B.n218 10.6151
R1373 B.n434 B.n433 10.6151
R1374 B.n435 B.n434 10.6151
R1375 B.n435 B.n216 10.6151
R1376 B.n439 B.n216 10.6151
R1377 B.n440 B.n439 10.6151
R1378 B.n441 B.n440 10.6151
R1379 B.n441 B.n214 10.6151
R1380 B.n445 B.n214 10.6151
R1381 B.n446 B.n445 10.6151
R1382 B.n447 B.n446 10.6151
R1383 B.n447 B.n212 10.6151
R1384 B.n451 B.n212 10.6151
R1385 B.n452 B.n451 10.6151
R1386 B.n453 B.n452 10.6151
R1387 B.n453 B.n210 10.6151
R1388 B.n457 B.n210 10.6151
R1389 B.n458 B.n457 10.6151
R1390 B.n460 B.n206 10.6151
R1391 B.n464 B.n206 10.6151
R1392 B.n465 B.n464 10.6151
R1393 B.n466 B.n465 10.6151
R1394 B.n466 B.n204 10.6151
R1395 B.n470 B.n204 10.6151
R1396 B.n471 B.n470 10.6151
R1397 B.n472 B.n471 10.6151
R1398 B.n476 B.n475 10.6151
R1399 B.n477 B.n476 10.6151
R1400 B.n477 B.n198 10.6151
R1401 B.n481 B.n198 10.6151
R1402 B.n482 B.n481 10.6151
R1403 B.n483 B.n482 10.6151
R1404 B.n483 B.n196 10.6151
R1405 B.n487 B.n196 10.6151
R1406 B.n488 B.n487 10.6151
R1407 B.n489 B.n488 10.6151
R1408 B.n489 B.n194 10.6151
R1409 B.n493 B.n194 10.6151
R1410 B.n494 B.n493 10.6151
R1411 B.n495 B.n494 10.6151
R1412 B.n495 B.n192 10.6151
R1413 B.n499 B.n192 10.6151
R1414 B.n500 B.n499 10.6151
R1415 B.n501 B.n500 10.6151
R1416 B.n501 B.n190 10.6151
R1417 B.n505 B.n190 10.6151
R1418 B.n506 B.n505 10.6151
R1419 B.n507 B.n506 10.6151
R1420 B.n507 B.n188 10.6151
R1421 B.n511 B.n188 10.6151
R1422 B.n512 B.n511 10.6151
R1423 B.n513 B.n512 10.6151
R1424 B.n513 B.n186 10.6151
R1425 B.n517 B.n186 10.6151
R1426 B.n518 B.n517 10.6151
R1427 B.n519 B.n518 10.6151
R1428 B.n519 B.n184 10.6151
R1429 B.n523 B.n184 10.6151
R1430 B.n524 B.n523 10.6151
R1431 B.n525 B.n524 10.6151
R1432 B.n525 B.n182 10.6151
R1433 B.n529 B.n182 10.6151
R1434 B.n530 B.n529 10.6151
R1435 B.n531 B.n530 10.6151
R1436 B.n531 B.n180 10.6151
R1437 B.n535 B.n180 10.6151
R1438 B.n536 B.n535 10.6151
R1439 B.n537 B.n536 10.6151
R1440 B.n537 B.n178 10.6151
R1441 B.n541 B.n178 10.6151
R1442 B.n542 B.n541 10.6151
R1443 B.n543 B.n542 10.6151
R1444 B.n543 B.n176 10.6151
R1445 B.n547 B.n176 10.6151
R1446 B.n548 B.n547 10.6151
R1447 B.n549 B.n548 10.6151
R1448 B.n549 B.n174 10.6151
R1449 B.n553 B.n174 10.6151
R1450 B.n554 B.n553 10.6151
R1451 B.n555 B.n554 10.6151
R1452 B.n555 B.n172 10.6151
R1453 B.n559 B.n172 10.6151
R1454 B.n560 B.n559 10.6151
R1455 B.n561 B.n560 10.6151
R1456 B.n561 B.n170 10.6151
R1457 B.n368 B.n367 10.6151
R1458 B.n367 B.n240 10.6151
R1459 B.n363 B.n240 10.6151
R1460 B.n363 B.n362 10.6151
R1461 B.n362 B.n361 10.6151
R1462 B.n361 B.n242 10.6151
R1463 B.n357 B.n242 10.6151
R1464 B.n357 B.n356 10.6151
R1465 B.n356 B.n355 10.6151
R1466 B.n355 B.n244 10.6151
R1467 B.n351 B.n244 10.6151
R1468 B.n351 B.n350 10.6151
R1469 B.n350 B.n349 10.6151
R1470 B.n349 B.n246 10.6151
R1471 B.n345 B.n246 10.6151
R1472 B.n345 B.n344 10.6151
R1473 B.n344 B.n343 10.6151
R1474 B.n343 B.n248 10.6151
R1475 B.n339 B.n248 10.6151
R1476 B.n339 B.n338 10.6151
R1477 B.n338 B.n337 10.6151
R1478 B.n337 B.n250 10.6151
R1479 B.n333 B.n250 10.6151
R1480 B.n333 B.n332 10.6151
R1481 B.n332 B.n331 10.6151
R1482 B.n331 B.n252 10.6151
R1483 B.n327 B.n252 10.6151
R1484 B.n327 B.n326 10.6151
R1485 B.n326 B.n325 10.6151
R1486 B.n325 B.n254 10.6151
R1487 B.n321 B.n254 10.6151
R1488 B.n321 B.n320 10.6151
R1489 B.n320 B.n319 10.6151
R1490 B.n319 B.n256 10.6151
R1491 B.n315 B.n256 10.6151
R1492 B.n315 B.n314 10.6151
R1493 B.n314 B.n313 10.6151
R1494 B.n313 B.n258 10.6151
R1495 B.n309 B.n258 10.6151
R1496 B.n309 B.n308 10.6151
R1497 B.n308 B.n307 10.6151
R1498 B.n307 B.n260 10.6151
R1499 B.n303 B.n260 10.6151
R1500 B.n303 B.n302 10.6151
R1501 B.n302 B.n301 10.6151
R1502 B.n301 B.n262 10.6151
R1503 B.n297 B.n262 10.6151
R1504 B.n297 B.n296 10.6151
R1505 B.n296 B.n295 10.6151
R1506 B.n295 B.n264 10.6151
R1507 B.n291 B.n264 10.6151
R1508 B.n291 B.n290 10.6151
R1509 B.n290 B.n289 10.6151
R1510 B.n289 B.n266 10.6151
R1511 B.n285 B.n266 10.6151
R1512 B.n285 B.n284 10.6151
R1513 B.n284 B.n283 10.6151
R1514 B.n283 B.n268 10.6151
R1515 B.n279 B.n268 10.6151
R1516 B.n279 B.n278 10.6151
R1517 B.n278 B.n277 10.6151
R1518 B.n277 B.n270 10.6151
R1519 B.n273 B.n270 10.6151
R1520 B.n273 B.n272 10.6151
R1521 B.n272 B.n0 10.6151
R1522 B.n1055 B.n1 10.6151
R1523 B.n1055 B.n1054 10.6151
R1524 B.n1054 B.n1053 10.6151
R1525 B.n1053 B.n4 10.6151
R1526 B.n1049 B.n4 10.6151
R1527 B.n1049 B.n1048 10.6151
R1528 B.n1048 B.n1047 10.6151
R1529 B.n1047 B.n6 10.6151
R1530 B.n1043 B.n6 10.6151
R1531 B.n1043 B.n1042 10.6151
R1532 B.n1042 B.n1041 10.6151
R1533 B.n1041 B.n8 10.6151
R1534 B.n1037 B.n8 10.6151
R1535 B.n1037 B.n1036 10.6151
R1536 B.n1036 B.n1035 10.6151
R1537 B.n1035 B.n10 10.6151
R1538 B.n1031 B.n10 10.6151
R1539 B.n1031 B.n1030 10.6151
R1540 B.n1030 B.n1029 10.6151
R1541 B.n1029 B.n12 10.6151
R1542 B.n1025 B.n12 10.6151
R1543 B.n1025 B.n1024 10.6151
R1544 B.n1024 B.n1023 10.6151
R1545 B.n1023 B.n14 10.6151
R1546 B.n1019 B.n14 10.6151
R1547 B.n1019 B.n1018 10.6151
R1548 B.n1018 B.n1017 10.6151
R1549 B.n1017 B.n16 10.6151
R1550 B.n1013 B.n16 10.6151
R1551 B.n1013 B.n1012 10.6151
R1552 B.n1012 B.n1011 10.6151
R1553 B.n1011 B.n18 10.6151
R1554 B.n1007 B.n18 10.6151
R1555 B.n1007 B.n1006 10.6151
R1556 B.n1006 B.n1005 10.6151
R1557 B.n1005 B.n20 10.6151
R1558 B.n1001 B.n20 10.6151
R1559 B.n1001 B.n1000 10.6151
R1560 B.n1000 B.n999 10.6151
R1561 B.n999 B.n22 10.6151
R1562 B.n995 B.n22 10.6151
R1563 B.n995 B.n994 10.6151
R1564 B.n994 B.n993 10.6151
R1565 B.n993 B.n24 10.6151
R1566 B.n989 B.n24 10.6151
R1567 B.n989 B.n988 10.6151
R1568 B.n988 B.n987 10.6151
R1569 B.n987 B.n26 10.6151
R1570 B.n983 B.n26 10.6151
R1571 B.n983 B.n982 10.6151
R1572 B.n982 B.n981 10.6151
R1573 B.n981 B.n28 10.6151
R1574 B.n977 B.n28 10.6151
R1575 B.n977 B.n976 10.6151
R1576 B.n976 B.n975 10.6151
R1577 B.n975 B.n30 10.6151
R1578 B.n971 B.n30 10.6151
R1579 B.n971 B.n970 10.6151
R1580 B.n970 B.n969 10.6151
R1581 B.n969 B.n32 10.6151
R1582 B.n965 B.n32 10.6151
R1583 B.n965 B.n964 10.6151
R1584 B.n964 B.n963 10.6151
R1585 B.n963 B.n34 10.6151
R1586 B.n959 B.n34 10.6151
R1587 B.n868 B.n867 6.5566
R1588 B.n855 B.n854 6.5566
R1589 B.n460 B.n459 6.5566
R1590 B.n472 B.n202 6.5566
R1591 B.n869 B.n868 4.05904
R1592 B.n854 B.n853 4.05904
R1593 B.n459 B.n458 4.05904
R1594 B.n475 B.n202 4.05904
R1595 B.n1059 B.n0 2.81026
R1596 B.n1059 B.n1 2.81026
R1597 VP.n24 VP.n21 161.3
R1598 VP.n26 VP.n25 161.3
R1599 VP.n27 VP.n20 161.3
R1600 VP.n29 VP.n28 161.3
R1601 VP.n30 VP.n19 161.3
R1602 VP.n32 VP.n31 161.3
R1603 VP.n33 VP.n18 161.3
R1604 VP.n36 VP.n35 161.3
R1605 VP.n37 VP.n17 161.3
R1606 VP.n39 VP.n38 161.3
R1607 VP.n40 VP.n16 161.3
R1608 VP.n42 VP.n41 161.3
R1609 VP.n43 VP.n15 161.3
R1610 VP.n45 VP.n44 161.3
R1611 VP.n46 VP.n14 161.3
R1612 VP.n48 VP.n47 161.3
R1613 VP.n89 VP.n88 161.3
R1614 VP.n87 VP.n1 161.3
R1615 VP.n86 VP.n85 161.3
R1616 VP.n84 VP.n2 161.3
R1617 VP.n83 VP.n82 161.3
R1618 VP.n81 VP.n3 161.3
R1619 VP.n80 VP.n79 161.3
R1620 VP.n78 VP.n4 161.3
R1621 VP.n77 VP.n76 161.3
R1622 VP.n74 VP.n5 161.3
R1623 VP.n73 VP.n72 161.3
R1624 VP.n71 VP.n6 161.3
R1625 VP.n70 VP.n69 161.3
R1626 VP.n68 VP.n7 161.3
R1627 VP.n67 VP.n66 161.3
R1628 VP.n65 VP.n8 161.3
R1629 VP.n64 VP.n63 161.3
R1630 VP.n61 VP.n9 161.3
R1631 VP.n60 VP.n59 161.3
R1632 VP.n58 VP.n10 161.3
R1633 VP.n57 VP.n56 161.3
R1634 VP.n55 VP.n11 161.3
R1635 VP.n54 VP.n53 161.3
R1636 VP.n52 VP.n12 161.3
R1637 VP.n23 VP.t1 153.655
R1638 VP.n50 VP.t5 120.635
R1639 VP.n62 VP.t4 120.635
R1640 VP.n75 VP.t3 120.635
R1641 VP.n0 VP.t2 120.635
R1642 VP.n13 VP.t0 120.635
R1643 VP.n34 VP.t7 120.635
R1644 VP.n22 VP.t6 120.635
R1645 VP.n51 VP.n50 82.238
R1646 VP.n90 VP.n0 82.238
R1647 VP.n49 VP.n13 82.238
R1648 VP.n23 VP.n22 63.7683
R1649 VP.n51 VP.n49 60.3024
R1650 VP.n56 VP.n10 56.5193
R1651 VP.n69 VP.n6 56.5193
R1652 VP.n82 VP.n2 56.5193
R1653 VP.n41 VP.n15 56.5193
R1654 VP.n28 VP.n19 56.5193
R1655 VP.n54 VP.n12 24.4675
R1656 VP.n55 VP.n54 24.4675
R1657 VP.n56 VP.n55 24.4675
R1658 VP.n60 VP.n10 24.4675
R1659 VP.n61 VP.n60 24.4675
R1660 VP.n63 VP.n61 24.4675
R1661 VP.n67 VP.n8 24.4675
R1662 VP.n68 VP.n67 24.4675
R1663 VP.n69 VP.n68 24.4675
R1664 VP.n73 VP.n6 24.4675
R1665 VP.n74 VP.n73 24.4675
R1666 VP.n76 VP.n74 24.4675
R1667 VP.n80 VP.n4 24.4675
R1668 VP.n81 VP.n80 24.4675
R1669 VP.n82 VP.n81 24.4675
R1670 VP.n86 VP.n2 24.4675
R1671 VP.n87 VP.n86 24.4675
R1672 VP.n88 VP.n87 24.4675
R1673 VP.n45 VP.n15 24.4675
R1674 VP.n46 VP.n45 24.4675
R1675 VP.n47 VP.n46 24.4675
R1676 VP.n32 VP.n19 24.4675
R1677 VP.n33 VP.n32 24.4675
R1678 VP.n35 VP.n33 24.4675
R1679 VP.n39 VP.n17 24.4675
R1680 VP.n40 VP.n39 24.4675
R1681 VP.n41 VP.n40 24.4675
R1682 VP.n26 VP.n21 24.4675
R1683 VP.n27 VP.n26 24.4675
R1684 VP.n28 VP.n27 24.4675
R1685 VP.n63 VP.n62 13.702
R1686 VP.n75 VP.n4 13.702
R1687 VP.n34 VP.n17 13.702
R1688 VP.n62 VP.n8 10.766
R1689 VP.n76 VP.n75 10.766
R1690 VP.n35 VP.n34 10.766
R1691 VP.n22 VP.n21 10.766
R1692 VP.n50 VP.n12 7.82994
R1693 VP.n88 VP.n0 7.82994
R1694 VP.n47 VP.n13 7.82994
R1695 VP.n24 VP.n23 3.22778
R1696 VP.n49 VP.n48 0.354971
R1697 VP.n52 VP.n51 0.354971
R1698 VP.n90 VP.n89 0.354971
R1699 VP VP.n90 0.26696
R1700 VP.n25 VP.n24 0.189894
R1701 VP.n25 VP.n20 0.189894
R1702 VP.n29 VP.n20 0.189894
R1703 VP.n30 VP.n29 0.189894
R1704 VP.n31 VP.n30 0.189894
R1705 VP.n31 VP.n18 0.189894
R1706 VP.n36 VP.n18 0.189894
R1707 VP.n37 VP.n36 0.189894
R1708 VP.n38 VP.n37 0.189894
R1709 VP.n38 VP.n16 0.189894
R1710 VP.n42 VP.n16 0.189894
R1711 VP.n43 VP.n42 0.189894
R1712 VP.n44 VP.n43 0.189894
R1713 VP.n44 VP.n14 0.189894
R1714 VP.n48 VP.n14 0.189894
R1715 VP.n53 VP.n52 0.189894
R1716 VP.n53 VP.n11 0.189894
R1717 VP.n57 VP.n11 0.189894
R1718 VP.n58 VP.n57 0.189894
R1719 VP.n59 VP.n58 0.189894
R1720 VP.n59 VP.n9 0.189894
R1721 VP.n64 VP.n9 0.189894
R1722 VP.n65 VP.n64 0.189894
R1723 VP.n66 VP.n65 0.189894
R1724 VP.n66 VP.n7 0.189894
R1725 VP.n70 VP.n7 0.189894
R1726 VP.n71 VP.n70 0.189894
R1727 VP.n72 VP.n71 0.189894
R1728 VP.n72 VP.n5 0.189894
R1729 VP.n77 VP.n5 0.189894
R1730 VP.n78 VP.n77 0.189894
R1731 VP.n79 VP.n78 0.189894
R1732 VP.n79 VP.n3 0.189894
R1733 VP.n83 VP.n3 0.189894
R1734 VP.n84 VP.n83 0.189894
R1735 VP.n85 VP.n84 0.189894
R1736 VP.n85 VP.n1 0.189894
R1737 VP.n89 VP.n1 0.189894
R1738 VTAIL.n806 VTAIL.n805 756.745
R1739 VTAIL.n100 VTAIL.n99 756.745
R1740 VTAIL.n200 VTAIL.n199 756.745
R1741 VTAIL.n302 VTAIL.n301 756.745
R1742 VTAIL.n706 VTAIL.n705 756.745
R1743 VTAIL.n604 VTAIL.n603 756.745
R1744 VTAIL.n504 VTAIL.n503 756.745
R1745 VTAIL.n402 VTAIL.n401 756.745
R1746 VTAIL.n741 VTAIL.n740 585
R1747 VTAIL.n738 VTAIL.n737 585
R1748 VTAIL.n747 VTAIL.n746 585
R1749 VTAIL.n749 VTAIL.n748 585
R1750 VTAIL.n734 VTAIL.n733 585
R1751 VTAIL.n755 VTAIL.n754 585
R1752 VTAIL.n758 VTAIL.n757 585
R1753 VTAIL.n756 VTAIL.n730 585
R1754 VTAIL.n763 VTAIL.n729 585
R1755 VTAIL.n765 VTAIL.n764 585
R1756 VTAIL.n767 VTAIL.n766 585
R1757 VTAIL.n726 VTAIL.n725 585
R1758 VTAIL.n773 VTAIL.n772 585
R1759 VTAIL.n775 VTAIL.n774 585
R1760 VTAIL.n722 VTAIL.n721 585
R1761 VTAIL.n781 VTAIL.n780 585
R1762 VTAIL.n783 VTAIL.n782 585
R1763 VTAIL.n718 VTAIL.n717 585
R1764 VTAIL.n789 VTAIL.n788 585
R1765 VTAIL.n791 VTAIL.n790 585
R1766 VTAIL.n714 VTAIL.n713 585
R1767 VTAIL.n797 VTAIL.n796 585
R1768 VTAIL.n799 VTAIL.n798 585
R1769 VTAIL.n710 VTAIL.n709 585
R1770 VTAIL.n805 VTAIL.n804 585
R1771 VTAIL.n35 VTAIL.n34 585
R1772 VTAIL.n32 VTAIL.n31 585
R1773 VTAIL.n41 VTAIL.n40 585
R1774 VTAIL.n43 VTAIL.n42 585
R1775 VTAIL.n28 VTAIL.n27 585
R1776 VTAIL.n49 VTAIL.n48 585
R1777 VTAIL.n52 VTAIL.n51 585
R1778 VTAIL.n50 VTAIL.n24 585
R1779 VTAIL.n57 VTAIL.n23 585
R1780 VTAIL.n59 VTAIL.n58 585
R1781 VTAIL.n61 VTAIL.n60 585
R1782 VTAIL.n20 VTAIL.n19 585
R1783 VTAIL.n67 VTAIL.n66 585
R1784 VTAIL.n69 VTAIL.n68 585
R1785 VTAIL.n16 VTAIL.n15 585
R1786 VTAIL.n75 VTAIL.n74 585
R1787 VTAIL.n77 VTAIL.n76 585
R1788 VTAIL.n12 VTAIL.n11 585
R1789 VTAIL.n83 VTAIL.n82 585
R1790 VTAIL.n85 VTAIL.n84 585
R1791 VTAIL.n8 VTAIL.n7 585
R1792 VTAIL.n91 VTAIL.n90 585
R1793 VTAIL.n93 VTAIL.n92 585
R1794 VTAIL.n4 VTAIL.n3 585
R1795 VTAIL.n99 VTAIL.n98 585
R1796 VTAIL.n135 VTAIL.n134 585
R1797 VTAIL.n132 VTAIL.n131 585
R1798 VTAIL.n141 VTAIL.n140 585
R1799 VTAIL.n143 VTAIL.n142 585
R1800 VTAIL.n128 VTAIL.n127 585
R1801 VTAIL.n149 VTAIL.n148 585
R1802 VTAIL.n152 VTAIL.n151 585
R1803 VTAIL.n150 VTAIL.n124 585
R1804 VTAIL.n157 VTAIL.n123 585
R1805 VTAIL.n159 VTAIL.n158 585
R1806 VTAIL.n161 VTAIL.n160 585
R1807 VTAIL.n120 VTAIL.n119 585
R1808 VTAIL.n167 VTAIL.n166 585
R1809 VTAIL.n169 VTAIL.n168 585
R1810 VTAIL.n116 VTAIL.n115 585
R1811 VTAIL.n175 VTAIL.n174 585
R1812 VTAIL.n177 VTAIL.n176 585
R1813 VTAIL.n112 VTAIL.n111 585
R1814 VTAIL.n183 VTAIL.n182 585
R1815 VTAIL.n185 VTAIL.n184 585
R1816 VTAIL.n108 VTAIL.n107 585
R1817 VTAIL.n191 VTAIL.n190 585
R1818 VTAIL.n193 VTAIL.n192 585
R1819 VTAIL.n104 VTAIL.n103 585
R1820 VTAIL.n199 VTAIL.n198 585
R1821 VTAIL.n237 VTAIL.n236 585
R1822 VTAIL.n234 VTAIL.n233 585
R1823 VTAIL.n243 VTAIL.n242 585
R1824 VTAIL.n245 VTAIL.n244 585
R1825 VTAIL.n230 VTAIL.n229 585
R1826 VTAIL.n251 VTAIL.n250 585
R1827 VTAIL.n254 VTAIL.n253 585
R1828 VTAIL.n252 VTAIL.n226 585
R1829 VTAIL.n259 VTAIL.n225 585
R1830 VTAIL.n261 VTAIL.n260 585
R1831 VTAIL.n263 VTAIL.n262 585
R1832 VTAIL.n222 VTAIL.n221 585
R1833 VTAIL.n269 VTAIL.n268 585
R1834 VTAIL.n271 VTAIL.n270 585
R1835 VTAIL.n218 VTAIL.n217 585
R1836 VTAIL.n277 VTAIL.n276 585
R1837 VTAIL.n279 VTAIL.n278 585
R1838 VTAIL.n214 VTAIL.n213 585
R1839 VTAIL.n285 VTAIL.n284 585
R1840 VTAIL.n287 VTAIL.n286 585
R1841 VTAIL.n210 VTAIL.n209 585
R1842 VTAIL.n293 VTAIL.n292 585
R1843 VTAIL.n295 VTAIL.n294 585
R1844 VTAIL.n206 VTAIL.n205 585
R1845 VTAIL.n301 VTAIL.n300 585
R1846 VTAIL.n705 VTAIL.n704 585
R1847 VTAIL.n610 VTAIL.n609 585
R1848 VTAIL.n699 VTAIL.n698 585
R1849 VTAIL.n697 VTAIL.n696 585
R1850 VTAIL.n614 VTAIL.n613 585
R1851 VTAIL.n691 VTAIL.n690 585
R1852 VTAIL.n689 VTAIL.n688 585
R1853 VTAIL.n618 VTAIL.n617 585
R1854 VTAIL.n683 VTAIL.n682 585
R1855 VTAIL.n681 VTAIL.n680 585
R1856 VTAIL.n622 VTAIL.n621 585
R1857 VTAIL.n675 VTAIL.n674 585
R1858 VTAIL.n673 VTAIL.n672 585
R1859 VTAIL.n626 VTAIL.n625 585
R1860 VTAIL.n667 VTAIL.n666 585
R1861 VTAIL.n665 VTAIL.n664 585
R1862 VTAIL.n663 VTAIL.n629 585
R1863 VTAIL.n633 VTAIL.n630 585
R1864 VTAIL.n658 VTAIL.n657 585
R1865 VTAIL.n656 VTAIL.n655 585
R1866 VTAIL.n635 VTAIL.n634 585
R1867 VTAIL.n650 VTAIL.n649 585
R1868 VTAIL.n648 VTAIL.n647 585
R1869 VTAIL.n639 VTAIL.n638 585
R1870 VTAIL.n642 VTAIL.n641 585
R1871 VTAIL.n603 VTAIL.n602 585
R1872 VTAIL.n508 VTAIL.n507 585
R1873 VTAIL.n597 VTAIL.n596 585
R1874 VTAIL.n595 VTAIL.n594 585
R1875 VTAIL.n512 VTAIL.n511 585
R1876 VTAIL.n589 VTAIL.n588 585
R1877 VTAIL.n587 VTAIL.n586 585
R1878 VTAIL.n516 VTAIL.n515 585
R1879 VTAIL.n581 VTAIL.n580 585
R1880 VTAIL.n579 VTAIL.n578 585
R1881 VTAIL.n520 VTAIL.n519 585
R1882 VTAIL.n573 VTAIL.n572 585
R1883 VTAIL.n571 VTAIL.n570 585
R1884 VTAIL.n524 VTAIL.n523 585
R1885 VTAIL.n565 VTAIL.n564 585
R1886 VTAIL.n563 VTAIL.n562 585
R1887 VTAIL.n561 VTAIL.n527 585
R1888 VTAIL.n531 VTAIL.n528 585
R1889 VTAIL.n556 VTAIL.n555 585
R1890 VTAIL.n554 VTAIL.n553 585
R1891 VTAIL.n533 VTAIL.n532 585
R1892 VTAIL.n548 VTAIL.n547 585
R1893 VTAIL.n546 VTAIL.n545 585
R1894 VTAIL.n537 VTAIL.n536 585
R1895 VTAIL.n540 VTAIL.n539 585
R1896 VTAIL.n503 VTAIL.n502 585
R1897 VTAIL.n408 VTAIL.n407 585
R1898 VTAIL.n497 VTAIL.n496 585
R1899 VTAIL.n495 VTAIL.n494 585
R1900 VTAIL.n412 VTAIL.n411 585
R1901 VTAIL.n489 VTAIL.n488 585
R1902 VTAIL.n487 VTAIL.n486 585
R1903 VTAIL.n416 VTAIL.n415 585
R1904 VTAIL.n481 VTAIL.n480 585
R1905 VTAIL.n479 VTAIL.n478 585
R1906 VTAIL.n420 VTAIL.n419 585
R1907 VTAIL.n473 VTAIL.n472 585
R1908 VTAIL.n471 VTAIL.n470 585
R1909 VTAIL.n424 VTAIL.n423 585
R1910 VTAIL.n465 VTAIL.n464 585
R1911 VTAIL.n463 VTAIL.n462 585
R1912 VTAIL.n461 VTAIL.n427 585
R1913 VTAIL.n431 VTAIL.n428 585
R1914 VTAIL.n456 VTAIL.n455 585
R1915 VTAIL.n454 VTAIL.n453 585
R1916 VTAIL.n433 VTAIL.n432 585
R1917 VTAIL.n448 VTAIL.n447 585
R1918 VTAIL.n446 VTAIL.n445 585
R1919 VTAIL.n437 VTAIL.n436 585
R1920 VTAIL.n440 VTAIL.n439 585
R1921 VTAIL.n401 VTAIL.n400 585
R1922 VTAIL.n306 VTAIL.n305 585
R1923 VTAIL.n395 VTAIL.n394 585
R1924 VTAIL.n393 VTAIL.n392 585
R1925 VTAIL.n310 VTAIL.n309 585
R1926 VTAIL.n387 VTAIL.n386 585
R1927 VTAIL.n385 VTAIL.n384 585
R1928 VTAIL.n314 VTAIL.n313 585
R1929 VTAIL.n379 VTAIL.n378 585
R1930 VTAIL.n377 VTAIL.n376 585
R1931 VTAIL.n318 VTAIL.n317 585
R1932 VTAIL.n371 VTAIL.n370 585
R1933 VTAIL.n369 VTAIL.n368 585
R1934 VTAIL.n322 VTAIL.n321 585
R1935 VTAIL.n363 VTAIL.n362 585
R1936 VTAIL.n361 VTAIL.n360 585
R1937 VTAIL.n359 VTAIL.n325 585
R1938 VTAIL.n329 VTAIL.n326 585
R1939 VTAIL.n354 VTAIL.n353 585
R1940 VTAIL.n352 VTAIL.n351 585
R1941 VTAIL.n331 VTAIL.n330 585
R1942 VTAIL.n346 VTAIL.n345 585
R1943 VTAIL.n344 VTAIL.n343 585
R1944 VTAIL.n335 VTAIL.n334 585
R1945 VTAIL.n338 VTAIL.n337 585
R1946 VTAIL.t15 VTAIL.n739 329.036
R1947 VTAIL.t2 VTAIL.n33 329.036
R1948 VTAIL.t8 VTAIL.n133 329.036
R1949 VTAIL.t13 VTAIL.n235 329.036
R1950 VTAIL.t12 VTAIL.n538 329.036
R1951 VTAIL.t6 VTAIL.n438 329.036
R1952 VTAIL.t1 VTAIL.n336 329.036
R1953 VTAIL.t10 VTAIL.n640 329.036
R1954 VTAIL.n740 VTAIL.n737 171.744
R1955 VTAIL.n747 VTAIL.n737 171.744
R1956 VTAIL.n748 VTAIL.n747 171.744
R1957 VTAIL.n748 VTAIL.n733 171.744
R1958 VTAIL.n755 VTAIL.n733 171.744
R1959 VTAIL.n757 VTAIL.n755 171.744
R1960 VTAIL.n757 VTAIL.n756 171.744
R1961 VTAIL.n756 VTAIL.n729 171.744
R1962 VTAIL.n765 VTAIL.n729 171.744
R1963 VTAIL.n766 VTAIL.n765 171.744
R1964 VTAIL.n766 VTAIL.n725 171.744
R1965 VTAIL.n773 VTAIL.n725 171.744
R1966 VTAIL.n774 VTAIL.n773 171.744
R1967 VTAIL.n774 VTAIL.n721 171.744
R1968 VTAIL.n781 VTAIL.n721 171.744
R1969 VTAIL.n782 VTAIL.n781 171.744
R1970 VTAIL.n782 VTAIL.n717 171.744
R1971 VTAIL.n789 VTAIL.n717 171.744
R1972 VTAIL.n790 VTAIL.n789 171.744
R1973 VTAIL.n790 VTAIL.n713 171.744
R1974 VTAIL.n797 VTAIL.n713 171.744
R1975 VTAIL.n798 VTAIL.n797 171.744
R1976 VTAIL.n798 VTAIL.n709 171.744
R1977 VTAIL.n805 VTAIL.n709 171.744
R1978 VTAIL.n34 VTAIL.n31 171.744
R1979 VTAIL.n41 VTAIL.n31 171.744
R1980 VTAIL.n42 VTAIL.n41 171.744
R1981 VTAIL.n42 VTAIL.n27 171.744
R1982 VTAIL.n49 VTAIL.n27 171.744
R1983 VTAIL.n51 VTAIL.n49 171.744
R1984 VTAIL.n51 VTAIL.n50 171.744
R1985 VTAIL.n50 VTAIL.n23 171.744
R1986 VTAIL.n59 VTAIL.n23 171.744
R1987 VTAIL.n60 VTAIL.n59 171.744
R1988 VTAIL.n60 VTAIL.n19 171.744
R1989 VTAIL.n67 VTAIL.n19 171.744
R1990 VTAIL.n68 VTAIL.n67 171.744
R1991 VTAIL.n68 VTAIL.n15 171.744
R1992 VTAIL.n75 VTAIL.n15 171.744
R1993 VTAIL.n76 VTAIL.n75 171.744
R1994 VTAIL.n76 VTAIL.n11 171.744
R1995 VTAIL.n83 VTAIL.n11 171.744
R1996 VTAIL.n84 VTAIL.n83 171.744
R1997 VTAIL.n84 VTAIL.n7 171.744
R1998 VTAIL.n91 VTAIL.n7 171.744
R1999 VTAIL.n92 VTAIL.n91 171.744
R2000 VTAIL.n92 VTAIL.n3 171.744
R2001 VTAIL.n99 VTAIL.n3 171.744
R2002 VTAIL.n134 VTAIL.n131 171.744
R2003 VTAIL.n141 VTAIL.n131 171.744
R2004 VTAIL.n142 VTAIL.n141 171.744
R2005 VTAIL.n142 VTAIL.n127 171.744
R2006 VTAIL.n149 VTAIL.n127 171.744
R2007 VTAIL.n151 VTAIL.n149 171.744
R2008 VTAIL.n151 VTAIL.n150 171.744
R2009 VTAIL.n150 VTAIL.n123 171.744
R2010 VTAIL.n159 VTAIL.n123 171.744
R2011 VTAIL.n160 VTAIL.n159 171.744
R2012 VTAIL.n160 VTAIL.n119 171.744
R2013 VTAIL.n167 VTAIL.n119 171.744
R2014 VTAIL.n168 VTAIL.n167 171.744
R2015 VTAIL.n168 VTAIL.n115 171.744
R2016 VTAIL.n175 VTAIL.n115 171.744
R2017 VTAIL.n176 VTAIL.n175 171.744
R2018 VTAIL.n176 VTAIL.n111 171.744
R2019 VTAIL.n183 VTAIL.n111 171.744
R2020 VTAIL.n184 VTAIL.n183 171.744
R2021 VTAIL.n184 VTAIL.n107 171.744
R2022 VTAIL.n191 VTAIL.n107 171.744
R2023 VTAIL.n192 VTAIL.n191 171.744
R2024 VTAIL.n192 VTAIL.n103 171.744
R2025 VTAIL.n199 VTAIL.n103 171.744
R2026 VTAIL.n236 VTAIL.n233 171.744
R2027 VTAIL.n243 VTAIL.n233 171.744
R2028 VTAIL.n244 VTAIL.n243 171.744
R2029 VTAIL.n244 VTAIL.n229 171.744
R2030 VTAIL.n251 VTAIL.n229 171.744
R2031 VTAIL.n253 VTAIL.n251 171.744
R2032 VTAIL.n253 VTAIL.n252 171.744
R2033 VTAIL.n252 VTAIL.n225 171.744
R2034 VTAIL.n261 VTAIL.n225 171.744
R2035 VTAIL.n262 VTAIL.n261 171.744
R2036 VTAIL.n262 VTAIL.n221 171.744
R2037 VTAIL.n269 VTAIL.n221 171.744
R2038 VTAIL.n270 VTAIL.n269 171.744
R2039 VTAIL.n270 VTAIL.n217 171.744
R2040 VTAIL.n277 VTAIL.n217 171.744
R2041 VTAIL.n278 VTAIL.n277 171.744
R2042 VTAIL.n278 VTAIL.n213 171.744
R2043 VTAIL.n285 VTAIL.n213 171.744
R2044 VTAIL.n286 VTAIL.n285 171.744
R2045 VTAIL.n286 VTAIL.n209 171.744
R2046 VTAIL.n293 VTAIL.n209 171.744
R2047 VTAIL.n294 VTAIL.n293 171.744
R2048 VTAIL.n294 VTAIL.n205 171.744
R2049 VTAIL.n301 VTAIL.n205 171.744
R2050 VTAIL.n705 VTAIL.n609 171.744
R2051 VTAIL.n698 VTAIL.n609 171.744
R2052 VTAIL.n698 VTAIL.n697 171.744
R2053 VTAIL.n697 VTAIL.n613 171.744
R2054 VTAIL.n690 VTAIL.n613 171.744
R2055 VTAIL.n690 VTAIL.n689 171.744
R2056 VTAIL.n689 VTAIL.n617 171.744
R2057 VTAIL.n682 VTAIL.n617 171.744
R2058 VTAIL.n682 VTAIL.n681 171.744
R2059 VTAIL.n681 VTAIL.n621 171.744
R2060 VTAIL.n674 VTAIL.n621 171.744
R2061 VTAIL.n674 VTAIL.n673 171.744
R2062 VTAIL.n673 VTAIL.n625 171.744
R2063 VTAIL.n666 VTAIL.n625 171.744
R2064 VTAIL.n666 VTAIL.n665 171.744
R2065 VTAIL.n665 VTAIL.n629 171.744
R2066 VTAIL.n633 VTAIL.n629 171.744
R2067 VTAIL.n657 VTAIL.n633 171.744
R2068 VTAIL.n657 VTAIL.n656 171.744
R2069 VTAIL.n656 VTAIL.n634 171.744
R2070 VTAIL.n649 VTAIL.n634 171.744
R2071 VTAIL.n649 VTAIL.n648 171.744
R2072 VTAIL.n648 VTAIL.n638 171.744
R2073 VTAIL.n641 VTAIL.n638 171.744
R2074 VTAIL.n603 VTAIL.n507 171.744
R2075 VTAIL.n596 VTAIL.n507 171.744
R2076 VTAIL.n596 VTAIL.n595 171.744
R2077 VTAIL.n595 VTAIL.n511 171.744
R2078 VTAIL.n588 VTAIL.n511 171.744
R2079 VTAIL.n588 VTAIL.n587 171.744
R2080 VTAIL.n587 VTAIL.n515 171.744
R2081 VTAIL.n580 VTAIL.n515 171.744
R2082 VTAIL.n580 VTAIL.n579 171.744
R2083 VTAIL.n579 VTAIL.n519 171.744
R2084 VTAIL.n572 VTAIL.n519 171.744
R2085 VTAIL.n572 VTAIL.n571 171.744
R2086 VTAIL.n571 VTAIL.n523 171.744
R2087 VTAIL.n564 VTAIL.n523 171.744
R2088 VTAIL.n564 VTAIL.n563 171.744
R2089 VTAIL.n563 VTAIL.n527 171.744
R2090 VTAIL.n531 VTAIL.n527 171.744
R2091 VTAIL.n555 VTAIL.n531 171.744
R2092 VTAIL.n555 VTAIL.n554 171.744
R2093 VTAIL.n554 VTAIL.n532 171.744
R2094 VTAIL.n547 VTAIL.n532 171.744
R2095 VTAIL.n547 VTAIL.n546 171.744
R2096 VTAIL.n546 VTAIL.n536 171.744
R2097 VTAIL.n539 VTAIL.n536 171.744
R2098 VTAIL.n503 VTAIL.n407 171.744
R2099 VTAIL.n496 VTAIL.n407 171.744
R2100 VTAIL.n496 VTAIL.n495 171.744
R2101 VTAIL.n495 VTAIL.n411 171.744
R2102 VTAIL.n488 VTAIL.n411 171.744
R2103 VTAIL.n488 VTAIL.n487 171.744
R2104 VTAIL.n487 VTAIL.n415 171.744
R2105 VTAIL.n480 VTAIL.n415 171.744
R2106 VTAIL.n480 VTAIL.n479 171.744
R2107 VTAIL.n479 VTAIL.n419 171.744
R2108 VTAIL.n472 VTAIL.n419 171.744
R2109 VTAIL.n472 VTAIL.n471 171.744
R2110 VTAIL.n471 VTAIL.n423 171.744
R2111 VTAIL.n464 VTAIL.n423 171.744
R2112 VTAIL.n464 VTAIL.n463 171.744
R2113 VTAIL.n463 VTAIL.n427 171.744
R2114 VTAIL.n431 VTAIL.n427 171.744
R2115 VTAIL.n455 VTAIL.n431 171.744
R2116 VTAIL.n455 VTAIL.n454 171.744
R2117 VTAIL.n454 VTAIL.n432 171.744
R2118 VTAIL.n447 VTAIL.n432 171.744
R2119 VTAIL.n447 VTAIL.n446 171.744
R2120 VTAIL.n446 VTAIL.n436 171.744
R2121 VTAIL.n439 VTAIL.n436 171.744
R2122 VTAIL.n401 VTAIL.n305 171.744
R2123 VTAIL.n394 VTAIL.n305 171.744
R2124 VTAIL.n394 VTAIL.n393 171.744
R2125 VTAIL.n393 VTAIL.n309 171.744
R2126 VTAIL.n386 VTAIL.n309 171.744
R2127 VTAIL.n386 VTAIL.n385 171.744
R2128 VTAIL.n385 VTAIL.n313 171.744
R2129 VTAIL.n378 VTAIL.n313 171.744
R2130 VTAIL.n378 VTAIL.n377 171.744
R2131 VTAIL.n377 VTAIL.n317 171.744
R2132 VTAIL.n370 VTAIL.n317 171.744
R2133 VTAIL.n370 VTAIL.n369 171.744
R2134 VTAIL.n369 VTAIL.n321 171.744
R2135 VTAIL.n362 VTAIL.n321 171.744
R2136 VTAIL.n362 VTAIL.n361 171.744
R2137 VTAIL.n361 VTAIL.n325 171.744
R2138 VTAIL.n329 VTAIL.n325 171.744
R2139 VTAIL.n353 VTAIL.n329 171.744
R2140 VTAIL.n353 VTAIL.n352 171.744
R2141 VTAIL.n352 VTAIL.n330 171.744
R2142 VTAIL.n345 VTAIL.n330 171.744
R2143 VTAIL.n345 VTAIL.n344 171.744
R2144 VTAIL.n344 VTAIL.n334 171.744
R2145 VTAIL.n337 VTAIL.n334 171.744
R2146 VTAIL.n740 VTAIL.t15 85.8723
R2147 VTAIL.n34 VTAIL.t2 85.8723
R2148 VTAIL.n134 VTAIL.t8 85.8723
R2149 VTAIL.n236 VTAIL.t13 85.8723
R2150 VTAIL.n641 VTAIL.t10 85.8723
R2151 VTAIL.n539 VTAIL.t12 85.8723
R2152 VTAIL.n439 VTAIL.t6 85.8723
R2153 VTAIL.n337 VTAIL.t1 85.8723
R2154 VTAIL.n607 VTAIL.n606 55.3449
R2155 VTAIL.n405 VTAIL.n404 55.3449
R2156 VTAIL.n1 VTAIL.n0 55.3447
R2157 VTAIL.n203 VTAIL.n202 55.3447
R2158 VTAIL.n807 VTAIL.n806 34.7066
R2159 VTAIL.n101 VTAIL.n100 34.7066
R2160 VTAIL.n201 VTAIL.n200 34.7066
R2161 VTAIL.n303 VTAIL.n302 34.7066
R2162 VTAIL.n707 VTAIL.n706 34.7066
R2163 VTAIL.n605 VTAIL.n604 34.7066
R2164 VTAIL.n505 VTAIL.n504 34.7066
R2165 VTAIL.n403 VTAIL.n402 34.7066
R2166 VTAIL.n807 VTAIL.n707 31.341
R2167 VTAIL.n403 VTAIL.n303 31.341
R2168 VTAIL.n764 VTAIL.n763 13.1884
R2169 VTAIL.n58 VTAIL.n57 13.1884
R2170 VTAIL.n158 VTAIL.n157 13.1884
R2171 VTAIL.n260 VTAIL.n259 13.1884
R2172 VTAIL.n664 VTAIL.n663 13.1884
R2173 VTAIL.n562 VTAIL.n561 13.1884
R2174 VTAIL.n462 VTAIL.n461 13.1884
R2175 VTAIL.n360 VTAIL.n359 13.1884
R2176 VTAIL.n762 VTAIL.n730 12.8005
R2177 VTAIL.n767 VTAIL.n728 12.8005
R2178 VTAIL.n56 VTAIL.n24 12.8005
R2179 VTAIL.n61 VTAIL.n22 12.8005
R2180 VTAIL.n156 VTAIL.n124 12.8005
R2181 VTAIL.n161 VTAIL.n122 12.8005
R2182 VTAIL.n258 VTAIL.n226 12.8005
R2183 VTAIL.n263 VTAIL.n224 12.8005
R2184 VTAIL.n667 VTAIL.n628 12.8005
R2185 VTAIL.n662 VTAIL.n630 12.8005
R2186 VTAIL.n565 VTAIL.n526 12.8005
R2187 VTAIL.n560 VTAIL.n528 12.8005
R2188 VTAIL.n465 VTAIL.n426 12.8005
R2189 VTAIL.n460 VTAIL.n428 12.8005
R2190 VTAIL.n363 VTAIL.n324 12.8005
R2191 VTAIL.n358 VTAIL.n326 12.8005
R2192 VTAIL.n759 VTAIL.n758 12.0247
R2193 VTAIL.n768 VTAIL.n726 12.0247
R2194 VTAIL.n804 VTAIL.n708 12.0247
R2195 VTAIL.n53 VTAIL.n52 12.0247
R2196 VTAIL.n62 VTAIL.n20 12.0247
R2197 VTAIL.n98 VTAIL.n2 12.0247
R2198 VTAIL.n153 VTAIL.n152 12.0247
R2199 VTAIL.n162 VTAIL.n120 12.0247
R2200 VTAIL.n198 VTAIL.n102 12.0247
R2201 VTAIL.n255 VTAIL.n254 12.0247
R2202 VTAIL.n264 VTAIL.n222 12.0247
R2203 VTAIL.n300 VTAIL.n204 12.0247
R2204 VTAIL.n704 VTAIL.n608 12.0247
R2205 VTAIL.n668 VTAIL.n626 12.0247
R2206 VTAIL.n659 VTAIL.n658 12.0247
R2207 VTAIL.n602 VTAIL.n506 12.0247
R2208 VTAIL.n566 VTAIL.n524 12.0247
R2209 VTAIL.n557 VTAIL.n556 12.0247
R2210 VTAIL.n502 VTAIL.n406 12.0247
R2211 VTAIL.n466 VTAIL.n424 12.0247
R2212 VTAIL.n457 VTAIL.n456 12.0247
R2213 VTAIL.n400 VTAIL.n304 12.0247
R2214 VTAIL.n364 VTAIL.n322 12.0247
R2215 VTAIL.n355 VTAIL.n354 12.0247
R2216 VTAIL.n754 VTAIL.n732 11.249
R2217 VTAIL.n772 VTAIL.n771 11.249
R2218 VTAIL.n803 VTAIL.n710 11.249
R2219 VTAIL.n48 VTAIL.n26 11.249
R2220 VTAIL.n66 VTAIL.n65 11.249
R2221 VTAIL.n97 VTAIL.n4 11.249
R2222 VTAIL.n148 VTAIL.n126 11.249
R2223 VTAIL.n166 VTAIL.n165 11.249
R2224 VTAIL.n197 VTAIL.n104 11.249
R2225 VTAIL.n250 VTAIL.n228 11.249
R2226 VTAIL.n268 VTAIL.n267 11.249
R2227 VTAIL.n299 VTAIL.n206 11.249
R2228 VTAIL.n703 VTAIL.n610 11.249
R2229 VTAIL.n672 VTAIL.n671 11.249
R2230 VTAIL.n655 VTAIL.n632 11.249
R2231 VTAIL.n601 VTAIL.n508 11.249
R2232 VTAIL.n570 VTAIL.n569 11.249
R2233 VTAIL.n553 VTAIL.n530 11.249
R2234 VTAIL.n501 VTAIL.n408 11.249
R2235 VTAIL.n470 VTAIL.n469 11.249
R2236 VTAIL.n453 VTAIL.n430 11.249
R2237 VTAIL.n399 VTAIL.n306 11.249
R2238 VTAIL.n368 VTAIL.n367 11.249
R2239 VTAIL.n351 VTAIL.n328 11.249
R2240 VTAIL.n741 VTAIL.n739 10.7239
R2241 VTAIL.n35 VTAIL.n33 10.7239
R2242 VTAIL.n135 VTAIL.n133 10.7239
R2243 VTAIL.n237 VTAIL.n235 10.7239
R2244 VTAIL.n642 VTAIL.n640 10.7239
R2245 VTAIL.n540 VTAIL.n538 10.7239
R2246 VTAIL.n440 VTAIL.n438 10.7239
R2247 VTAIL.n338 VTAIL.n336 10.7239
R2248 VTAIL.n753 VTAIL.n734 10.4732
R2249 VTAIL.n775 VTAIL.n724 10.4732
R2250 VTAIL.n800 VTAIL.n799 10.4732
R2251 VTAIL.n47 VTAIL.n28 10.4732
R2252 VTAIL.n69 VTAIL.n18 10.4732
R2253 VTAIL.n94 VTAIL.n93 10.4732
R2254 VTAIL.n147 VTAIL.n128 10.4732
R2255 VTAIL.n169 VTAIL.n118 10.4732
R2256 VTAIL.n194 VTAIL.n193 10.4732
R2257 VTAIL.n249 VTAIL.n230 10.4732
R2258 VTAIL.n271 VTAIL.n220 10.4732
R2259 VTAIL.n296 VTAIL.n295 10.4732
R2260 VTAIL.n700 VTAIL.n699 10.4732
R2261 VTAIL.n675 VTAIL.n624 10.4732
R2262 VTAIL.n654 VTAIL.n635 10.4732
R2263 VTAIL.n598 VTAIL.n597 10.4732
R2264 VTAIL.n573 VTAIL.n522 10.4732
R2265 VTAIL.n552 VTAIL.n533 10.4732
R2266 VTAIL.n498 VTAIL.n497 10.4732
R2267 VTAIL.n473 VTAIL.n422 10.4732
R2268 VTAIL.n452 VTAIL.n433 10.4732
R2269 VTAIL.n396 VTAIL.n395 10.4732
R2270 VTAIL.n371 VTAIL.n320 10.4732
R2271 VTAIL.n350 VTAIL.n331 10.4732
R2272 VTAIL.n750 VTAIL.n749 9.69747
R2273 VTAIL.n776 VTAIL.n722 9.69747
R2274 VTAIL.n796 VTAIL.n712 9.69747
R2275 VTAIL.n44 VTAIL.n43 9.69747
R2276 VTAIL.n70 VTAIL.n16 9.69747
R2277 VTAIL.n90 VTAIL.n6 9.69747
R2278 VTAIL.n144 VTAIL.n143 9.69747
R2279 VTAIL.n170 VTAIL.n116 9.69747
R2280 VTAIL.n190 VTAIL.n106 9.69747
R2281 VTAIL.n246 VTAIL.n245 9.69747
R2282 VTAIL.n272 VTAIL.n218 9.69747
R2283 VTAIL.n292 VTAIL.n208 9.69747
R2284 VTAIL.n696 VTAIL.n612 9.69747
R2285 VTAIL.n676 VTAIL.n622 9.69747
R2286 VTAIL.n651 VTAIL.n650 9.69747
R2287 VTAIL.n594 VTAIL.n510 9.69747
R2288 VTAIL.n574 VTAIL.n520 9.69747
R2289 VTAIL.n549 VTAIL.n548 9.69747
R2290 VTAIL.n494 VTAIL.n410 9.69747
R2291 VTAIL.n474 VTAIL.n420 9.69747
R2292 VTAIL.n449 VTAIL.n448 9.69747
R2293 VTAIL.n392 VTAIL.n308 9.69747
R2294 VTAIL.n372 VTAIL.n318 9.69747
R2295 VTAIL.n347 VTAIL.n346 9.69747
R2296 VTAIL.n802 VTAIL.n708 9.45567
R2297 VTAIL.n96 VTAIL.n2 9.45567
R2298 VTAIL.n196 VTAIL.n102 9.45567
R2299 VTAIL.n298 VTAIL.n204 9.45567
R2300 VTAIL.n702 VTAIL.n608 9.45567
R2301 VTAIL.n600 VTAIL.n506 9.45567
R2302 VTAIL.n500 VTAIL.n406 9.45567
R2303 VTAIL.n398 VTAIL.n304 9.45567
R2304 VTAIL.n787 VTAIL.n786 9.3005
R2305 VTAIL.n716 VTAIL.n715 9.3005
R2306 VTAIL.n793 VTAIL.n792 9.3005
R2307 VTAIL.n795 VTAIL.n794 9.3005
R2308 VTAIL.n712 VTAIL.n711 9.3005
R2309 VTAIL.n801 VTAIL.n800 9.3005
R2310 VTAIL.n803 VTAIL.n802 9.3005
R2311 VTAIL.n720 VTAIL.n719 9.3005
R2312 VTAIL.n779 VTAIL.n778 9.3005
R2313 VTAIL.n777 VTAIL.n776 9.3005
R2314 VTAIL.n724 VTAIL.n723 9.3005
R2315 VTAIL.n771 VTAIL.n770 9.3005
R2316 VTAIL.n769 VTAIL.n768 9.3005
R2317 VTAIL.n728 VTAIL.n727 9.3005
R2318 VTAIL.n743 VTAIL.n742 9.3005
R2319 VTAIL.n745 VTAIL.n744 9.3005
R2320 VTAIL.n736 VTAIL.n735 9.3005
R2321 VTAIL.n751 VTAIL.n750 9.3005
R2322 VTAIL.n753 VTAIL.n752 9.3005
R2323 VTAIL.n732 VTAIL.n731 9.3005
R2324 VTAIL.n760 VTAIL.n759 9.3005
R2325 VTAIL.n762 VTAIL.n761 9.3005
R2326 VTAIL.n785 VTAIL.n784 9.3005
R2327 VTAIL.n81 VTAIL.n80 9.3005
R2328 VTAIL.n10 VTAIL.n9 9.3005
R2329 VTAIL.n87 VTAIL.n86 9.3005
R2330 VTAIL.n89 VTAIL.n88 9.3005
R2331 VTAIL.n6 VTAIL.n5 9.3005
R2332 VTAIL.n95 VTAIL.n94 9.3005
R2333 VTAIL.n97 VTAIL.n96 9.3005
R2334 VTAIL.n14 VTAIL.n13 9.3005
R2335 VTAIL.n73 VTAIL.n72 9.3005
R2336 VTAIL.n71 VTAIL.n70 9.3005
R2337 VTAIL.n18 VTAIL.n17 9.3005
R2338 VTAIL.n65 VTAIL.n64 9.3005
R2339 VTAIL.n63 VTAIL.n62 9.3005
R2340 VTAIL.n22 VTAIL.n21 9.3005
R2341 VTAIL.n37 VTAIL.n36 9.3005
R2342 VTAIL.n39 VTAIL.n38 9.3005
R2343 VTAIL.n30 VTAIL.n29 9.3005
R2344 VTAIL.n45 VTAIL.n44 9.3005
R2345 VTAIL.n47 VTAIL.n46 9.3005
R2346 VTAIL.n26 VTAIL.n25 9.3005
R2347 VTAIL.n54 VTAIL.n53 9.3005
R2348 VTAIL.n56 VTAIL.n55 9.3005
R2349 VTAIL.n79 VTAIL.n78 9.3005
R2350 VTAIL.n181 VTAIL.n180 9.3005
R2351 VTAIL.n110 VTAIL.n109 9.3005
R2352 VTAIL.n187 VTAIL.n186 9.3005
R2353 VTAIL.n189 VTAIL.n188 9.3005
R2354 VTAIL.n106 VTAIL.n105 9.3005
R2355 VTAIL.n195 VTAIL.n194 9.3005
R2356 VTAIL.n197 VTAIL.n196 9.3005
R2357 VTAIL.n114 VTAIL.n113 9.3005
R2358 VTAIL.n173 VTAIL.n172 9.3005
R2359 VTAIL.n171 VTAIL.n170 9.3005
R2360 VTAIL.n118 VTAIL.n117 9.3005
R2361 VTAIL.n165 VTAIL.n164 9.3005
R2362 VTAIL.n163 VTAIL.n162 9.3005
R2363 VTAIL.n122 VTAIL.n121 9.3005
R2364 VTAIL.n137 VTAIL.n136 9.3005
R2365 VTAIL.n139 VTAIL.n138 9.3005
R2366 VTAIL.n130 VTAIL.n129 9.3005
R2367 VTAIL.n145 VTAIL.n144 9.3005
R2368 VTAIL.n147 VTAIL.n146 9.3005
R2369 VTAIL.n126 VTAIL.n125 9.3005
R2370 VTAIL.n154 VTAIL.n153 9.3005
R2371 VTAIL.n156 VTAIL.n155 9.3005
R2372 VTAIL.n179 VTAIL.n178 9.3005
R2373 VTAIL.n283 VTAIL.n282 9.3005
R2374 VTAIL.n212 VTAIL.n211 9.3005
R2375 VTAIL.n289 VTAIL.n288 9.3005
R2376 VTAIL.n291 VTAIL.n290 9.3005
R2377 VTAIL.n208 VTAIL.n207 9.3005
R2378 VTAIL.n297 VTAIL.n296 9.3005
R2379 VTAIL.n299 VTAIL.n298 9.3005
R2380 VTAIL.n216 VTAIL.n215 9.3005
R2381 VTAIL.n275 VTAIL.n274 9.3005
R2382 VTAIL.n273 VTAIL.n272 9.3005
R2383 VTAIL.n220 VTAIL.n219 9.3005
R2384 VTAIL.n267 VTAIL.n266 9.3005
R2385 VTAIL.n265 VTAIL.n264 9.3005
R2386 VTAIL.n224 VTAIL.n223 9.3005
R2387 VTAIL.n239 VTAIL.n238 9.3005
R2388 VTAIL.n241 VTAIL.n240 9.3005
R2389 VTAIL.n232 VTAIL.n231 9.3005
R2390 VTAIL.n247 VTAIL.n246 9.3005
R2391 VTAIL.n249 VTAIL.n248 9.3005
R2392 VTAIL.n228 VTAIL.n227 9.3005
R2393 VTAIL.n256 VTAIL.n255 9.3005
R2394 VTAIL.n258 VTAIL.n257 9.3005
R2395 VTAIL.n281 VTAIL.n280 9.3005
R2396 VTAIL.n703 VTAIL.n702 9.3005
R2397 VTAIL.n701 VTAIL.n700 9.3005
R2398 VTAIL.n612 VTAIL.n611 9.3005
R2399 VTAIL.n695 VTAIL.n694 9.3005
R2400 VTAIL.n693 VTAIL.n692 9.3005
R2401 VTAIL.n616 VTAIL.n615 9.3005
R2402 VTAIL.n687 VTAIL.n686 9.3005
R2403 VTAIL.n685 VTAIL.n684 9.3005
R2404 VTAIL.n620 VTAIL.n619 9.3005
R2405 VTAIL.n679 VTAIL.n678 9.3005
R2406 VTAIL.n677 VTAIL.n676 9.3005
R2407 VTAIL.n624 VTAIL.n623 9.3005
R2408 VTAIL.n671 VTAIL.n670 9.3005
R2409 VTAIL.n669 VTAIL.n668 9.3005
R2410 VTAIL.n628 VTAIL.n627 9.3005
R2411 VTAIL.n662 VTAIL.n661 9.3005
R2412 VTAIL.n660 VTAIL.n659 9.3005
R2413 VTAIL.n632 VTAIL.n631 9.3005
R2414 VTAIL.n654 VTAIL.n653 9.3005
R2415 VTAIL.n652 VTAIL.n651 9.3005
R2416 VTAIL.n637 VTAIL.n636 9.3005
R2417 VTAIL.n646 VTAIL.n645 9.3005
R2418 VTAIL.n644 VTAIL.n643 9.3005
R2419 VTAIL.n542 VTAIL.n541 9.3005
R2420 VTAIL.n544 VTAIL.n543 9.3005
R2421 VTAIL.n535 VTAIL.n534 9.3005
R2422 VTAIL.n550 VTAIL.n549 9.3005
R2423 VTAIL.n552 VTAIL.n551 9.3005
R2424 VTAIL.n530 VTAIL.n529 9.3005
R2425 VTAIL.n558 VTAIL.n557 9.3005
R2426 VTAIL.n560 VTAIL.n559 9.3005
R2427 VTAIL.n514 VTAIL.n513 9.3005
R2428 VTAIL.n591 VTAIL.n590 9.3005
R2429 VTAIL.n593 VTAIL.n592 9.3005
R2430 VTAIL.n510 VTAIL.n509 9.3005
R2431 VTAIL.n599 VTAIL.n598 9.3005
R2432 VTAIL.n601 VTAIL.n600 9.3005
R2433 VTAIL.n585 VTAIL.n584 9.3005
R2434 VTAIL.n583 VTAIL.n582 9.3005
R2435 VTAIL.n518 VTAIL.n517 9.3005
R2436 VTAIL.n577 VTAIL.n576 9.3005
R2437 VTAIL.n575 VTAIL.n574 9.3005
R2438 VTAIL.n522 VTAIL.n521 9.3005
R2439 VTAIL.n569 VTAIL.n568 9.3005
R2440 VTAIL.n567 VTAIL.n566 9.3005
R2441 VTAIL.n526 VTAIL.n525 9.3005
R2442 VTAIL.n442 VTAIL.n441 9.3005
R2443 VTAIL.n444 VTAIL.n443 9.3005
R2444 VTAIL.n435 VTAIL.n434 9.3005
R2445 VTAIL.n450 VTAIL.n449 9.3005
R2446 VTAIL.n452 VTAIL.n451 9.3005
R2447 VTAIL.n430 VTAIL.n429 9.3005
R2448 VTAIL.n458 VTAIL.n457 9.3005
R2449 VTAIL.n460 VTAIL.n459 9.3005
R2450 VTAIL.n414 VTAIL.n413 9.3005
R2451 VTAIL.n491 VTAIL.n490 9.3005
R2452 VTAIL.n493 VTAIL.n492 9.3005
R2453 VTAIL.n410 VTAIL.n409 9.3005
R2454 VTAIL.n499 VTAIL.n498 9.3005
R2455 VTAIL.n501 VTAIL.n500 9.3005
R2456 VTAIL.n485 VTAIL.n484 9.3005
R2457 VTAIL.n483 VTAIL.n482 9.3005
R2458 VTAIL.n418 VTAIL.n417 9.3005
R2459 VTAIL.n477 VTAIL.n476 9.3005
R2460 VTAIL.n475 VTAIL.n474 9.3005
R2461 VTAIL.n422 VTAIL.n421 9.3005
R2462 VTAIL.n469 VTAIL.n468 9.3005
R2463 VTAIL.n467 VTAIL.n466 9.3005
R2464 VTAIL.n426 VTAIL.n425 9.3005
R2465 VTAIL.n340 VTAIL.n339 9.3005
R2466 VTAIL.n342 VTAIL.n341 9.3005
R2467 VTAIL.n333 VTAIL.n332 9.3005
R2468 VTAIL.n348 VTAIL.n347 9.3005
R2469 VTAIL.n350 VTAIL.n349 9.3005
R2470 VTAIL.n328 VTAIL.n327 9.3005
R2471 VTAIL.n356 VTAIL.n355 9.3005
R2472 VTAIL.n358 VTAIL.n357 9.3005
R2473 VTAIL.n312 VTAIL.n311 9.3005
R2474 VTAIL.n389 VTAIL.n388 9.3005
R2475 VTAIL.n391 VTAIL.n390 9.3005
R2476 VTAIL.n308 VTAIL.n307 9.3005
R2477 VTAIL.n397 VTAIL.n396 9.3005
R2478 VTAIL.n399 VTAIL.n398 9.3005
R2479 VTAIL.n383 VTAIL.n382 9.3005
R2480 VTAIL.n381 VTAIL.n380 9.3005
R2481 VTAIL.n316 VTAIL.n315 9.3005
R2482 VTAIL.n375 VTAIL.n374 9.3005
R2483 VTAIL.n373 VTAIL.n372 9.3005
R2484 VTAIL.n320 VTAIL.n319 9.3005
R2485 VTAIL.n367 VTAIL.n366 9.3005
R2486 VTAIL.n365 VTAIL.n364 9.3005
R2487 VTAIL.n324 VTAIL.n323 9.3005
R2488 VTAIL.n746 VTAIL.n736 8.92171
R2489 VTAIL.n780 VTAIL.n779 8.92171
R2490 VTAIL.n795 VTAIL.n714 8.92171
R2491 VTAIL.n40 VTAIL.n30 8.92171
R2492 VTAIL.n74 VTAIL.n73 8.92171
R2493 VTAIL.n89 VTAIL.n8 8.92171
R2494 VTAIL.n140 VTAIL.n130 8.92171
R2495 VTAIL.n174 VTAIL.n173 8.92171
R2496 VTAIL.n189 VTAIL.n108 8.92171
R2497 VTAIL.n242 VTAIL.n232 8.92171
R2498 VTAIL.n276 VTAIL.n275 8.92171
R2499 VTAIL.n291 VTAIL.n210 8.92171
R2500 VTAIL.n695 VTAIL.n614 8.92171
R2501 VTAIL.n680 VTAIL.n679 8.92171
R2502 VTAIL.n647 VTAIL.n637 8.92171
R2503 VTAIL.n593 VTAIL.n512 8.92171
R2504 VTAIL.n578 VTAIL.n577 8.92171
R2505 VTAIL.n545 VTAIL.n535 8.92171
R2506 VTAIL.n493 VTAIL.n412 8.92171
R2507 VTAIL.n478 VTAIL.n477 8.92171
R2508 VTAIL.n445 VTAIL.n435 8.92171
R2509 VTAIL.n391 VTAIL.n310 8.92171
R2510 VTAIL.n376 VTAIL.n375 8.92171
R2511 VTAIL.n343 VTAIL.n333 8.92171
R2512 VTAIL.n745 VTAIL.n738 8.14595
R2513 VTAIL.n783 VTAIL.n720 8.14595
R2514 VTAIL.n792 VTAIL.n791 8.14595
R2515 VTAIL.n39 VTAIL.n32 8.14595
R2516 VTAIL.n77 VTAIL.n14 8.14595
R2517 VTAIL.n86 VTAIL.n85 8.14595
R2518 VTAIL.n139 VTAIL.n132 8.14595
R2519 VTAIL.n177 VTAIL.n114 8.14595
R2520 VTAIL.n186 VTAIL.n185 8.14595
R2521 VTAIL.n241 VTAIL.n234 8.14595
R2522 VTAIL.n279 VTAIL.n216 8.14595
R2523 VTAIL.n288 VTAIL.n287 8.14595
R2524 VTAIL.n692 VTAIL.n691 8.14595
R2525 VTAIL.n683 VTAIL.n620 8.14595
R2526 VTAIL.n646 VTAIL.n639 8.14595
R2527 VTAIL.n590 VTAIL.n589 8.14595
R2528 VTAIL.n581 VTAIL.n518 8.14595
R2529 VTAIL.n544 VTAIL.n537 8.14595
R2530 VTAIL.n490 VTAIL.n489 8.14595
R2531 VTAIL.n481 VTAIL.n418 8.14595
R2532 VTAIL.n444 VTAIL.n437 8.14595
R2533 VTAIL.n388 VTAIL.n387 8.14595
R2534 VTAIL.n379 VTAIL.n316 8.14595
R2535 VTAIL.n342 VTAIL.n335 8.14595
R2536 VTAIL.n742 VTAIL.n741 7.3702
R2537 VTAIL.n784 VTAIL.n718 7.3702
R2538 VTAIL.n788 VTAIL.n716 7.3702
R2539 VTAIL.n36 VTAIL.n35 7.3702
R2540 VTAIL.n78 VTAIL.n12 7.3702
R2541 VTAIL.n82 VTAIL.n10 7.3702
R2542 VTAIL.n136 VTAIL.n135 7.3702
R2543 VTAIL.n178 VTAIL.n112 7.3702
R2544 VTAIL.n182 VTAIL.n110 7.3702
R2545 VTAIL.n238 VTAIL.n237 7.3702
R2546 VTAIL.n280 VTAIL.n214 7.3702
R2547 VTAIL.n284 VTAIL.n212 7.3702
R2548 VTAIL.n688 VTAIL.n616 7.3702
R2549 VTAIL.n684 VTAIL.n618 7.3702
R2550 VTAIL.n643 VTAIL.n642 7.3702
R2551 VTAIL.n586 VTAIL.n514 7.3702
R2552 VTAIL.n582 VTAIL.n516 7.3702
R2553 VTAIL.n541 VTAIL.n540 7.3702
R2554 VTAIL.n486 VTAIL.n414 7.3702
R2555 VTAIL.n482 VTAIL.n416 7.3702
R2556 VTAIL.n441 VTAIL.n440 7.3702
R2557 VTAIL.n384 VTAIL.n312 7.3702
R2558 VTAIL.n380 VTAIL.n314 7.3702
R2559 VTAIL.n339 VTAIL.n338 7.3702
R2560 VTAIL.n787 VTAIL.n718 6.59444
R2561 VTAIL.n788 VTAIL.n787 6.59444
R2562 VTAIL.n81 VTAIL.n12 6.59444
R2563 VTAIL.n82 VTAIL.n81 6.59444
R2564 VTAIL.n181 VTAIL.n112 6.59444
R2565 VTAIL.n182 VTAIL.n181 6.59444
R2566 VTAIL.n283 VTAIL.n214 6.59444
R2567 VTAIL.n284 VTAIL.n283 6.59444
R2568 VTAIL.n688 VTAIL.n687 6.59444
R2569 VTAIL.n687 VTAIL.n618 6.59444
R2570 VTAIL.n586 VTAIL.n585 6.59444
R2571 VTAIL.n585 VTAIL.n516 6.59444
R2572 VTAIL.n486 VTAIL.n485 6.59444
R2573 VTAIL.n485 VTAIL.n416 6.59444
R2574 VTAIL.n384 VTAIL.n383 6.59444
R2575 VTAIL.n383 VTAIL.n314 6.59444
R2576 VTAIL.n742 VTAIL.n738 5.81868
R2577 VTAIL.n784 VTAIL.n783 5.81868
R2578 VTAIL.n791 VTAIL.n716 5.81868
R2579 VTAIL.n36 VTAIL.n32 5.81868
R2580 VTAIL.n78 VTAIL.n77 5.81868
R2581 VTAIL.n85 VTAIL.n10 5.81868
R2582 VTAIL.n136 VTAIL.n132 5.81868
R2583 VTAIL.n178 VTAIL.n177 5.81868
R2584 VTAIL.n185 VTAIL.n110 5.81868
R2585 VTAIL.n238 VTAIL.n234 5.81868
R2586 VTAIL.n280 VTAIL.n279 5.81868
R2587 VTAIL.n287 VTAIL.n212 5.81868
R2588 VTAIL.n691 VTAIL.n616 5.81868
R2589 VTAIL.n684 VTAIL.n683 5.81868
R2590 VTAIL.n643 VTAIL.n639 5.81868
R2591 VTAIL.n589 VTAIL.n514 5.81868
R2592 VTAIL.n582 VTAIL.n581 5.81868
R2593 VTAIL.n541 VTAIL.n537 5.81868
R2594 VTAIL.n489 VTAIL.n414 5.81868
R2595 VTAIL.n482 VTAIL.n481 5.81868
R2596 VTAIL.n441 VTAIL.n437 5.81868
R2597 VTAIL.n387 VTAIL.n312 5.81868
R2598 VTAIL.n380 VTAIL.n379 5.81868
R2599 VTAIL.n339 VTAIL.n335 5.81868
R2600 VTAIL.n746 VTAIL.n745 5.04292
R2601 VTAIL.n780 VTAIL.n720 5.04292
R2602 VTAIL.n792 VTAIL.n714 5.04292
R2603 VTAIL.n40 VTAIL.n39 5.04292
R2604 VTAIL.n74 VTAIL.n14 5.04292
R2605 VTAIL.n86 VTAIL.n8 5.04292
R2606 VTAIL.n140 VTAIL.n139 5.04292
R2607 VTAIL.n174 VTAIL.n114 5.04292
R2608 VTAIL.n186 VTAIL.n108 5.04292
R2609 VTAIL.n242 VTAIL.n241 5.04292
R2610 VTAIL.n276 VTAIL.n216 5.04292
R2611 VTAIL.n288 VTAIL.n210 5.04292
R2612 VTAIL.n692 VTAIL.n614 5.04292
R2613 VTAIL.n680 VTAIL.n620 5.04292
R2614 VTAIL.n647 VTAIL.n646 5.04292
R2615 VTAIL.n590 VTAIL.n512 5.04292
R2616 VTAIL.n578 VTAIL.n518 5.04292
R2617 VTAIL.n545 VTAIL.n544 5.04292
R2618 VTAIL.n490 VTAIL.n412 5.04292
R2619 VTAIL.n478 VTAIL.n418 5.04292
R2620 VTAIL.n445 VTAIL.n444 5.04292
R2621 VTAIL.n388 VTAIL.n310 5.04292
R2622 VTAIL.n376 VTAIL.n316 5.04292
R2623 VTAIL.n343 VTAIL.n342 5.04292
R2624 VTAIL.n749 VTAIL.n736 4.26717
R2625 VTAIL.n779 VTAIL.n722 4.26717
R2626 VTAIL.n796 VTAIL.n795 4.26717
R2627 VTAIL.n43 VTAIL.n30 4.26717
R2628 VTAIL.n73 VTAIL.n16 4.26717
R2629 VTAIL.n90 VTAIL.n89 4.26717
R2630 VTAIL.n143 VTAIL.n130 4.26717
R2631 VTAIL.n173 VTAIL.n116 4.26717
R2632 VTAIL.n190 VTAIL.n189 4.26717
R2633 VTAIL.n245 VTAIL.n232 4.26717
R2634 VTAIL.n275 VTAIL.n218 4.26717
R2635 VTAIL.n292 VTAIL.n291 4.26717
R2636 VTAIL.n696 VTAIL.n695 4.26717
R2637 VTAIL.n679 VTAIL.n622 4.26717
R2638 VTAIL.n650 VTAIL.n637 4.26717
R2639 VTAIL.n594 VTAIL.n593 4.26717
R2640 VTAIL.n577 VTAIL.n520 4.26717
R2641 VTAIL.n548 VTAIL.n535 4.26717
R2642 VTAIL.n494 VTAIL.n493 4.26717
R2643 VTAIL.n477 VTAIL.n420 4.26717
R2644 VTAIL.n448 VTAIL.n435 4.26717
R2645 VTAIL.n392 VTAIL.n391 4.26717
R2646 VTAIL.n375 VTAIL.n318 4.26717
R2647 VTAIL.n346 VTAIL.n333 4.26717
R2648 VTAIL.n750 VTAIL.n734 3.49141
R2649 VTAIL.n776 VTAIL.n775 3.49141
R2650 VTAIL.n799 VTAIL.n712 3.49141
R2651 VTAIL.n44 VTAIL.n28 3.49141
R2652 VTAIL.n70 VTAIL.n69 3.49141
R2653 VTAIL.n93 VTAIL.n6 3.49141
R2654 VTAIL.n144 VTAIL.n128 3.49141
R2655 VTAIL.n170 VTAIL.n169 3.49141
R2656 VTAIL.n193 VTAIL.n106 3.49141
R2657 VTAIL.n246 VTAIL.n230 3.49141
R2658 VTAIL.n272 VTAIL.n271 3.49141
R2659 VTAIL.n295 VTAIL.n208 3.49141
R2660 VTAIL.n699 VTAIL.n612 3.49141
R2661 VTAIL.n676 VTAIL.n675 3.49141
R2662 VTAIL.n651 VTAIL.n635 3.49141
R2663 VTAIL.n597 VTAIL.n510 3.49141
R2664 VTAIL.n574 VTAIL.n573 3.49141
R2665 VTAIL.n549 VTAIL.n533 3.49141
R2666 VTAIL.n497 VTAIL.n410 3.49141
R2667 VTAIL.n474 VTAIL.n473 3.49141
R2668 VTAIL.n449 VTAIL.n433 3.49141
R2669 VTAIL.n395 VTAIL.n308 3.49141
R2670 VTAIL.n372 VTAIL.n371 3.49141
R2671 VTAIL.n347 VTAIL.n331 3.49141
R2672 VTAIL.n405 VTAIL.n403 3.39705
R2673 VTAIL.n505 VTAIL.n405 3.39705
R2674 VTAIL.n607 VTAIL.n605 3.39705
R2675 VTAIL.n707 VTAIL.n607 3.39705
R2676 VTAIL.n303 VTAIL.n203 3.39705
R2677 VTAIL.n203 VTAIL.n201 3.39705
R2678 VTAIL.n101 VTAIL.n1 3.39705
R2679 VTAIL VTAIL.n807 3.33886
R2680 VTAIL.n754 VTAIL.n753 2.71565
R2681 VTAIL.n772 VTAIL.n724 2.71565
R2682 VTAIL.n800 VTAIL.n710 2.71565
R2683 VTAIL.n48 VTAIL.n47 2.71565
R2684 VTAIL.n66 VTAIL.n18 2.71565
R2685 VTAIL.n94 VTAIL.n4 2.71565
R2686 VTAIL.n148 VTAIL.n147 2.71565
R2687 VTAIL.n166 VTAIL.n118 2.71565
R2688 VTAIL.n194 VTAIL.n104 2.71565
R2689 VTAIL.n250 VTAIL.n249 2.71565
R2690 VTAIL.n268 VTAIL.n220 2.71565
R2691 VTAIL.n296 VTAIL.n206 2.71565
R2692 VTAIL.n700 VTAIL.n610 2.71565
R2693 VTAIL.n672 VTAIL.n624 2.71565
R2694 VTAIL.n655 VTAIL.n654 2.71565
R2695 VTAIL.n598 VTAIL.n508 2.71565
R2696 VTAIL.n570 VTAIL.n522 2.71565
R2697 VTAIL.n553 VTAIL.n552 2.71565
R2698 VTAIL.n498 VTAIL.n408 2.71565
R2699 VTAIL.n470 VTAIL.n422 2.71565
R2700 VTAIL.n453 VTAIL.n452 2.71565
R2701 VTAIL.n396 VTAIL.n306 2.71565
R2702 VTAIL.n368 VTAIL.n320 2.71565
R2703 VTAIL.n351 VTAIL.n350 2.71565
R2704 VTAIL.n743 VTAIL.n739 2.41282
R2705 VTAIL.n37 VTAIL.n33 2.41282
R2706 VTAIL.n137 VTAIL.n133 2.41282
R2707 VTAIL.n239 VTAIL.n235 2.41282
R2708 VTAIL.n644 VTAIL.n640 2.41282
R2709 VTAIL.n542 VTAIL.n538 2.41282
R2710 VTAIL.n442 VTAIL.n438 2.41282
R2711 VTAIL.n340 VTAIL.n336 2.41282
R2712 VTAIL.n758 VTAIL.n732 1.93989
R2713 VTAIL.n771 VTAIL.n726 1.93989
R2714 VTAIL.n804 VTAIL.n803 1.93989
R2715 VTAIL.n52 VTAIL.n26 1.93989
R2716 VTAIL.n65 VTAIL.n20 1.93989
R2717 VTAIL.n98 VTAIL.n97 1.93989
R2718 VTAIL.n152 VTAIL.n126 1.93989
R2719 VTAIL.n165 VTAIL.n120 1.93989
R2720 VTAIL.n198 VTAIL.n197 1.93989
R2721 VTAIL.n254 VTAIL.n228 1.93989
R2722 VTAIL.n267 VTAIL.n222 1.93989
R2723 VTAIL.n300 VTAIL.n299 1.93989
R2724 VTAIL.n704 VTAIL.n703 1.93989
R2725 VTAIL.n671 VTAIL.n626 1.93989
R2726 VTAIL.n658 VTAIL.n632 1.93989
R2727 VTAIL.n602 VTAIL.n601 1.93989
R2728 VTAIL.n569 VTAIL.n524 1.93989
R2729 VTAIL.n556 VTAIL.n530 1.93989
R2730 VTAIL.n502 VTAIL.n501 1.93989
R2731 VTAIL.n469 VTAIL.n424 1.93989
R2732 VTAIL.n456 VTAIL.n430 1.93989
R2733 VTAIL.n400 VTAIL.n399 1.93989
R2734 VTAIL.n367 VTAIL.n322 1.93989
R2735 VTAIL.n354 VTAIL.n328 1.93989
R2736 VTAIL.n0 VTAIL.t5 1.79934
R2737 VTAIL.n0 VTAIL.t4 1.79934
R2738 VTAIL.n202 VTAIL.t9 1.79934
R2739 VTAIL.n202 VTAIL.t7 1.79934
R2740 VTAIL.n606 VTAIL.t14 1.79934
R2741 VTAIL.n606 VTAIL.t11 1.79934
R2742 VTAIL.n404 VTAIL.t3 1.79934
R2743 VTAIL.n404 VTAIL.t0 1.79934
R2744 VTAIL.n759 VTAIL.n730 1.16414
R2745 VTAIL.n768 VTAIL.n767 1.16414
R2746 VTAIL.n806 VTAIL.n708 1.16414
R2747 VTAIL.n53 VTAIL.n24 1.16414
R2748 VTAIL.n62 VTAIL.n61 1.16414
R2749 VTAIL.n100 VTAIL.n2 1.16414
R2750 VTAIL.n153 VTAIL.n124 1.16414
R2751 VTAIL.n162 VTAIL.n161 1.16414
R2752 VTAIL.n200 VTAIL.n102 1.16414
R2753 VTAIL.n255 VTAIL.n226 1.16414
R2754 VTAIL.n264 VTAIL.n263 1.16414
R2755 VTAIL.n302 VTAIL.n204 1.16414
R2756 VTAIL.n706 VTAIL.n608 1.16414
R2757 VTAIL.n668 VTAIL.n667 1.16414
R2758 VTAIL.n659 VTAIL.n630 1.16414
R2759 VTAIL.n604 VTAIL.n506 1.16414
R2760 VTAIL.n566 VTAIL.n565 1.16414
R2761 VTAIL.n557 VTAIL.n528 1.16414
R2762 VTAIL.n504 VTAIL.n406 1.16414
R2763 VTAIL.n466 VTAIL.n465 1.16414
R2764 VTAIL.n457 VTAIL.n428 1.16414
R2765 VTAIL.n402 VTAIL.n304 1.16414
R2766 VTAIL.n364 VTAIL.n363 1.16414
R2767 VTAIL.n355 VTAIL.n326 1.16414
R2768 VTAIL.n605 VTAIL.n505 0.470328
R2769 VTAIL.n201 VTAIL.n101 0.470328
R2770 VTAIL.n763 VTAIL.n762 0.388379
R2771 VTAIL.n764 VTAIL.n728 0.388379
R2772 VTAIL.n57 VTAIL.n56 0.388379
R2773 VTAIL.n58 VTAIL.n22 0.388379
R2774 VTAIL.n157 VTAIL.n156 0.388379
R2775 VTAIL.n158 VTAIL.n122 0.388379
R2776 VTAIL.n259 VTAIL.n258 0.388379
R2777 VTAIL.n260 VTAIL.n224 0.388379
R2778 VTAIL.n664 VTAIL.n628 0.388379
R2779 VTAIL.n663 VTAIL.n662 0.388379
R2780 VTAIL.n562 VTAIL.n526 0.388379
R2781 VTAIL.n561 VTAIL.n560 0.388379
R2782 VTAIL.n462 VTAIL.n426 0.388379
R2783 VTAIL.n461 VTAIL.n460 0.388379
R2784 VTAIL.n360 VTAIL.n324 0.388379
R2785 VTAIL.n359 VTAIL.n358 0.388379
R2786 VTAIL.n744 VTAIL.n743 0.155672
R2787 VTAIL.n744 VTAIL.n735 0.155672
R2788 VTAIL.n751 VTAIL.n735 0.155672
R2789 VTAIL.n752 VTAIL.n751 0.155672
R2790 VTAIL.n752 VTAIL.n731 0.155672
R2791 VTAIL.n760 VTAIL.n731 0.155672
R2792 VTAIL.n761 VTAIL.n760 0.155672
R2793 VTAIL.n761 VTAIL.n727 0.155672
R2794 VTAIL.n769 VTAIL.n727 0.155672
R2795 VTAIL.n770 VTAIL.n769 0.155672
R2796 VTAIL.n770 VTAIL.n723 0.155672
R2797 VTAIL.n777 VTAIL.n723 0.155672
R2798 VTAIL.n778 VTAIL.n777 0.155672
R2799 VTAIL.n778 VTAIL.n719 0.155672
R2800 VTAIL.n785 VTAIL.n719 0.155672
R2801 VTAIL.n786 VTAIL.n785 0.155672
R2802 VTAIL.n786 VTAIL.n715 0.155672
R2803 VTAIL.n793 VTAIL.n715 0.155672
R2804 VTAIL.n794 VTAIL.n793 0.155672
R2805 VTAIL.n794 VTAIL.n711 0.155672
R2806 VTAIL.n801 VTAIL.n711 0.155672
R2807 VTAIL.n802 VTAIL.n801 0.155672
R2808 VTAIL.n38 VTAIL.n37 0.155672
R2809 VTAIL.n38 VTAIL.n29 0.155672
R2810 VTAIL.n45 VTAIL.n29 0.155672
R2811 VTAIL.n46 VTAIL.n45 0.155672
R2812 VTAIL.n46 VTAIL.n25 0.155672
R2813 VTAIL.n54 VTAIL.n25 0.155672
R2814 VTAIL.n55 VTAIL.n54 0.155672
R2815 VTAIL.n55 VTAIL.n21 0.155672
R2816 VTAIL.n63 VTAIL.n21 0.155672
R2817 VTAIL.n64 VTAIL.n63 0.155672
R2818 VTAIL.n64 VTAIL.n17 0.155672
R2819 VTAIL.n71 VTAIL.n17 0.155672
R2820 VTAIL.n72 VTAIL.n71 0.155672
R2821 VTAIL.n72 VTAIL.n13 0.155672
R2822 VTAIL.n79 VTAIL.n13 0.155672
R2823 VTAIL.n80 VTAIL.n79 0.155672
R2824 VTAIL.n80 VTAIL.n9 0.155672
R2825 VTAIL.n87 VTAIL.n9 0.155672
R2826 VTAIL.n88 VTAIL.n87 0.155672
R2827 VTAIL.n88 VTAIL.n5 0.155672
R2828 VTAIL.n95 VTAIL.n5 0.155672
R2829 VTAIL.n96 VTAIL.n95 0.155672
R2830 VTAIL.n138 VTAIL.n137 0.155672
R2831 VTAIL.n138 VTAIL.n129 0.155672
R2832 VTAIL.n145 VTAIL.n129 0.155672
R2833 VTAIL.n146 VTAIL.n145 0.155672
R2834 VTAIL.n146 VTAIL.n125 0.155672
R2835 VTAIL.n154 VTAIL.n125 0.155672
R2836 VTAIL.n155 VTAIL.n154 0.155672
R2837 VTAIL.n155 VTAIL.n121 0.155672
R2838 VTAIL.n163 VTAIL.n121 0.155672
R2839 VTAIL.n164 VTAIL.n163 0.155672
R2840 VTAIL.n164 VTAIL.n117 0.155672
R2841 VTAIL.n171 VTAIL.n117 0.155672
R2842 VTAIL.n172 VTAIL.n171 0.155672
R2843 VTAIL.n172 VTAIL.n113 0.155672
R2844 VTAIL.n179 VTAIL.n113 0.155672
R2845 VTAIL.n180 VTAIL.n179 0.155672
R2846 VTAIL.n180 VTAIL.n109 0.155672
R2847 VTAIL.n187 VTAIL.n109 0.155672
R2848 VTAIL.n188 VTAIL.n187 0.155672
R2849 VTAIL.n188 VTAIL.n105 0.155672
R2850 VTAIL.n195 VTAIL.n105 0.155672
R2851 VTAIL.n196 VTAIL.n195 0.155672
R2852 VTAIL.n240 VTAIL.n239 0.155672
R2853 VTAIL.n240 VTAIL.n231 0.155672
R2854 VTAIL.n247 VTAIL.n231 0.155672
R2855 VTAIL.n248 VTAIL.n247 0.155672
R2856 VTAIL.n248 VTAIL.n227 0.155672
R2857 VTAIL.n256 VTAIL.n227 0.155672
R2858 VTAIL.n257 VTAIL.n256 0.155672
R2859 VTAIL.n257 VTAIL.n223 0.155672
R2860 VTAIL.n265 VTAIL.n223 0.155672
R2861 VTAIL.n266 VTAIL.n265 0.155672
R2862 VTAIL.n266 VTAIL.n219 0.155672
R2863 VTAIL.n273 VTAIL.n219 0.155672
R2864 VTAIL.n274 VTAIL.n273 0.155672
R2865 VTAIL.n274 VTAIL.n215 0.155672
R2866 VTAIL.n281 VTAIL.n215 0.155672
R2867 VTAIL.n282 VTAIL.n281 0.155672
R2868 VTAIL.n282 VTAIL.n211 0.155672
R2869 VTAIL.n289 VTAIL.n211 0.155672
R2870 VTAIL.n290 VTAIL.n289 0.155672
R2871 VTAIL.n290 VTAIL.n207 0.155672
R2872 VTAIL.n297 VTAIL.n207 0.155672
R2873 VTAIL.n298 VTAIL.n297 0.155672
R2874 VTAIL.n702 VTAIL.n701 0.155672
R2875 VTAIL.n701 VTAIL.n611 0.155672
R2876 VTAIL.n694 VTAIL.n611 0.155672
R2877 VTAIL.n694 VTAIL.n693 0.155672
R2878 VTAIL.n693 VTAIL.n615 0.155672
R2879 VTAIL.n686 VTAIL.n615 0.155672
R2880 VTAIL.n686 VTAIL.n685 0.155672
R2881 VTAIL.n685 VTAIL.n619 0.155672
R2882 VTAIL.n678 VTAIL.n619 0.155672
R2883 VTAIL.n678 VTAIL.n677 0.155672
R2884 VTAIL.n677 VTAIL.n623 0.155672
R2885 VTAIL.n670 VTAIL.n623 0.155672
R2886 VTAIL.n670 VTAIL.n669 0.155672
R2887 VTAIL.n669 VTAIL.n627 0.155672
R2888 VTAIL.n661 VTAIL.n627 0.155672
R2889 VTAIL.n661 VTAIL.n660 0.155672
R2890 VTAIL.n660 VTAIL.n631 0.155672
R2891 VTAIL.n653 VTAIL.n631 0.155672
R2892 VTAIL.n653 VTAIL.n652 0.155672
R2893 VTAIL.n652 VTAIL.n636 0.155672
R2894 VTAIL.n645 VTAIL.n636 0.155672
R2895 VTAIL.n645 VTAIL.n644 0.155672
R2896 VTAIL.n600 VTAIL.n599 0.155672
R2897 VTAIL.n599 VTAIL.n509 0.155672
R2898 VTAIL.n592 VTAIL.n509 0.155672
R2899 VTAIL.n592 VTAIL.n591 0.155672
R2900 VTAIL.n591 VTAIL.n513 0.155672
R2901 VTAIL.n584 VTAIL.n513 0.155672
R2902 VTAIL.n584 VTAIL.n583 0.155672
R2903 VTAIL.n583 VTAIL.n517 0.155672
R2904 VTAIL.n576 VTAIL.n517 0.155672
R2905 VTAIL.n576 VTAIL.n575 0.155672
R2906 VTAIL.n575 VTAIL.n521 0.155672
R2907 VTAIL.n568 VTAIL.n521 0.155672
R2908 VTAIL.n568 VTAIL.n567 0.155672
R2909 VTAIL.n567 VTAIL.n525 0.155672
R2910 VTAIL.n559 VTAIL.n525 0.155672
R2911 VTAIL.n559 VTAIL.n558 0.155672
R2912 VTAIL.n558 VTAIL.n529 0.155672
R2913 VTAIL.n551 VTAIL.n529 0.155672
R2914 VTAIL.n551 VTAIL.n550 0.155672
R2915 VTAIL.n550 VTAIL.n534 0.155672
R2916 VTAIL.n543 VTAIL.n534 0.155672
R2917 VTAIL.n543 VTAIL.n542 0.155672
R2918 VTAIL.n500 VTAIL.n499 0.155672
R2919 VTAIL.n499 VTAIL.n409 0.155672
R2920 VTAIL.n492 VTAIL.n409 0.155672
R2921 VTAIL.n492 VTAIL.n491 0.155672
R2922 VTAIL.n491 VTAIL.n413 0.155672
R2923 VTAIL.n484 VTAIL.n413 0.155672
R2924 VTAIL.n484 VTAIL.n483 0.155672
R2925 VTAIL.n483 VTAIL.n417 0.155672
R2926 VTAIL.n476 VTAIL.n417 0.155672
R2927 VTAIL.n476 VTAIL.n475 0.155672
R2928 VTAIL.n475 VTAIL.n421 0.155672
R2929 VTAIL.n468 VTAIL.n421 0.155672
R2930 VTAIL.n468 VTAIL.n467 0.155672
R2931 VTAIL.n467 VTAIL.n425 0.155672
R2932 VTAIL.n459 VTAIL.n425 0.155672
R2933 VTAIL.n459 VTAIL.n458 0.155672
R2934 VTAIL.n458 VTAIL.n429 0.155672
R2935 VTAIL.n451 VTAIL.n429 0.155672
R2936 VTAIL.n451 VTAIL.n450 0.155672
R2937 VTAIL.n450 VTAIL.n434 0.155672
R2938 VTAIL.n443 VTAIL.n434 0.155672
R2939 VTAIL.n443 VTAIL.n442 0.155672
R2940 VTAIL.n398 VTAIL.n397 0.155672
R2941 VTAIL.n397 VTAIL.n307 0.155672
R2942 VTAIL.n390 VTAIL.n307 0.155672
R2943 VTAIL.n390 VTAIL.n389 0.155672
R2944 VTAIL.n389 VTAIL.n311 0.155672
R2945 VTAIL.n382 VTAIL.n311 0.155672
R2946 VTAIL.n382 VTAIL.n381 0.155672
R2947 VTAIL.n381 VTAIL.n315 0.155672
R2948 VTAIL.n374 VTAIL.n315 0.155672
R2949 VTAIL.n374 VTAIL.n373 0.155672
R2950 VTAIL.n373 VTAIL.n319 0.155672
R2951 VTAIL.n366 VTAIL.n319 0.155672
R2952 VTAIL.n366 VTAIL.n365 0.155672
R2953 VTAIL.n365 VTAIL.n323 0.155672
R2954 VTAIL.n357 VTAIL.n323 0.155672
R2955 VTAIL.n357 VTAIL.n356 0.155672
R2956 VTAIL.n356 VTAIL.n327 0.155672
R2957 VTAIL.n349 VTAIL.n327 0.155672
R2958 VTAIL.n349 VTAIL.n348 0.155672
R2959 VTAIL.n348 VTAIL.n332 0.155672
R2960 VTAIL.n341 VTAIL.n332 0.155672
R2961 VTAIL.n341 VTAIL.n340 0.155672
R2962 VTAIL VTAIL.n1 0.0586897
R2963 VDD1 VDD1.n0 73.7801
R2964 VDD1.n3 VDD1.n2 73.6664
R2965 VDD1.n3 VDD1.n1 73.6664
R2966 VDD1.n5 VDD1.n4 72.0225
R2967 VDD1.n5 VDD1.n3 55.1604
R2968 VDD1.n4 VDD1.t0 1.79934
R2969 VDD1.n4 VDD1.t7 1.79934
R2970 VDD1.n0 VDD1.t6 1.79934
R2971 VDD1.n0 VDD1.t1 1.79934
R2972 VDD1.n2 VDD1.t4 1.79934
R2973 VDD1.n2 VDD1.t5 1.79934
R2974 VDD1.n1 VDD1.t2 1.79934
R2975 VDD1.n1 VDD1.t3 1.79934
R2976 VDD1 VDD1.n5 1.64059
R2977 VN.n72 VN.n71 161.3
R2978 VN.n70 VN.n38 161.3
R2979 VN.n69 VN.n68 161.3
R2980 VN.n67 VN.n39 161.3
R2981 VN.n66 VN.n65 161.3
R2982 VN.n64 VN.n40 161.3
R2983 VN.n63 VN.n62 161.3
R2984 VN.n61 VN.n41 161.3
R2985 VN.n60 VN.n59 161.3
R2986 VN.n58 VN.n42 161.3
R2987 VN.n57 VN.n56 161.3
R2988 VN.n55 VN.n44 161.3
R2989 VN.n54 VN.n53 161.3
R2990 VN.n52 VN.n45 161.3
R2991 VN.n51 VN.n50 161.3
R2992 VN.n49 VN.n46 161.3
R2993 VN.n35 VN.n34 161.3
R2994 VN.n33 VN.n1 161.3
R2995 VN.n32 VN.n31 161.3
R2996 VN.n30 VN.n2 161.3
R2997 VN.n29 VN.n28 161.3
R2998 VN.n27 VN.n3 161.3
R2999 VN.n26 VN.n25 161.3
R3000 VN.n24 VN.n4 161.3
R3001 VN.n23 VN.n22 161.3
R3002 VN.n20 VN.n5 161.3
R3003 VN.n19 VN.n18 161.3
R3004 VN.n17 VN.n6 161.3
R3005 VN.n16 VN.n15 161.3
R3006 VN.n14 VN.n7 161.3
R3007 VN.n13 VN.n12 161.3
R3008 VN.n11 VN.n8 161.3
R3009 VN.n48 VN.t2 153.656
R3010 VN.n10 VN.t4 153.656
R3011 VN.n9 VN.t6 120.635
R3012 VN.n21 VN.t1 120.635
R3013 VN.n0 VN.t0 120.635
R3014 VN.n47 VN.t7 120.635
R3015 VN.n43 VN.t3 120.635
R3016 VN.n37 VN.t5 120.635
R3017 VN.n36 VN.n0 82.238
R3018 VN.n73 VN.n37 82.238
R3019 VN.n48 VN.n47 63.7683
R3020 VN.n10 VN.n9 63.7683
R3021 VN VN.n73 60.4677
R3022 VN.n15 VN.n6 56.5193
R3023 VN.n28 VN.n2 56.5193
R3024 VN.n53 VN.n44 56.5193
R3025 VN.n65 VN.n39 56.5193
R3026 VN.n13 VN.n8 24.4675
R3027 VN.n14 VN.n13 24.4675
R3028 VN.n15 VN.n14 24.4675
R3029 VN.n19 VN.n6 24.4675
R3030 VN.n20 VN.n19 24.4675
R3031 VN.n22 VN.n20 24.4675
R3032 VN.n26 VN.n4 24.4675
R3033 VN.n27 VN.n26 24.4675
R3034 VN.n28 VN.n27 24.4675
R3035 VN.n32 VN.n2 24.4675
R3036 VN.n33 VN.n32 24.4675
R3037 VN.n34 VN.n33 24.4675
R3038 VN.n53 VN.n52 24.4675
R3039 VN.n52 VN.n51 24.4675
R3040 VN.n51 VN.n46 24.4675
R3041 VN.n65 VN.n64 24.4675
R3042 VN.n64 VN.n63 24.4675
R3043 VN.n63 VN.n41 24.4675
R3044 VN.n59 VN.n58 24.4675
R3045 VN.n58 VN.n57 24.4675
R3046 VN.n57 VN.n44 24.4675
R3047 VN.n71 VN.n70 24.4675
R3048 VN.n70 VN.n69 24.4675
R3049 VN.n69 VN.n39 24.4675
R3050 VN.n21 VN.n4 13.702
R3051 VN.n43 VN.n41 13.702
R3052 VN.n9 VN.n8 10.766
R3053 VN.n22 VN.n21 10.766
R3054 VN.n47 VN.n46 10.766
R3055 VN.n59 VN.n43 10.766
R3056 VN.n34 VN.n0 7.82994
R3057 VN.n71 VN.n37 7.82994
R3058 VN.n49 VN.n48 3.22779
R3059 VN.n11 VN.n10 3.22779
R3060 VN.n73 VN.n72 0.354971
R3061 VN.n36 VN.n35 0.354971
R3062 VN VN.n36 0.26696
R3063 VN.n72 VN.n38 0.189894
R3064 VN.n68 VN.n38 0.189894
R3065 VN.n68 VN.n67 0.189894
R3066 VN.n67 VN.n66 0.189894
R3067 VN.n66 VN.n40 0.189894
R3068 VN.n62 VN.n40 0.189894
R3069 VN.n62 VN.n61 0.189894
R3070 VN.n61 VN.n60 0.189894
R3071 VN.n60 VN.n42 0.189894
R3072 VN.n56 VN.n42 0.189894
R3073 VN.n56 VN.n55 0.189894
R3074 VN.n55 VN.n54 0.189894
R3075 VN.n54 VN.n45 0.189894
R3076 VN.n50 VN.n45 0.189894
R3077 VN.n50 VN.n49 0.189894
R3078 VN.n12 VN.n11 0.189894
R3079 VN.n12 VN.n7 0.189894
R3080 VN.n16 VN.n7 0.189894
R3081 VN.n17 VN.n16 0.189894
R3082 VN.n18 VN.n17 0.189894
R3083 VN.n18 VN.n5 0.189894
R3084 VN.n23 VN.n5 0.189894
R3085 VN.n24 VN.n23 0.189894
R3086 VN.n25 VN.n24 0.189894
R3087 VN.n25 VN.n3 0.189894
R3088 VN.n29 VN.n3 0.189894
R3089 VN.n30 VN.n29 0.189894
R3090 VN.n31 VN.n30 0.189894
R3091 VN.n31 VN.n1 0.189894
R3092 VN.n35 VN.n1 0.189894
R3093 VDD2.n2 VDD2.n1 73.6664
R3094 VDD2.n2 VDD2.n0 73.6664
R3095 VDD2 VDD2.n5 73.6625
R3096 VDD2.n4 VDD2.n3 72.0236
R3097 VDD2.n4 VDD2.n2 54.5774
R3098 VDD2.n5 VDD2.t0 1.79934
R3099 VDD2.n5 VDD2.t5 1.79934
R3100 VDD2.n3 VDD2.t2 1.79934
R3101 VDD2.n3 VDD2.t4 1.79934
R3102 VDD2.n1 VDD2.t6 1.79934
R3103 VDD2.n1 VDD2.t7 1.79934
R3104 VDD2.n0 VDD2.t3 1.79934
R3105 VDD2.n0 VDD2.t1 1.79934
R3106 VDD2 VDD2.n4 1.75697
C0 VTAIL VP 14.0607f
C1 VP B 2.6105f
C2 VDD1 VP 14.0693f
C3 VTAIL VN 14.046599f
C4 VN B 1.53159f
C5 VDD2 w_n4910_n4582# 2.60183f
C6 VDD1 VN 0.153695f
C7 VTAIL B 7.49116f
C8 VDD2 VP 0.627287f
C9 VTAIL VDD1 10.2157f
C10 VDD1 B 2.12131f
C11 VDD2 VN 13.597599f
C12 VP w_n4910_n4582# 11.0238f
C13 VN w_n4910_n4582# 10.3834f
C14 VDD2 VTAIL 10.2769f
C15 VDD2 B 2.24911f
C16 VDD2 VDD1 2.30213f
C17 VP VN 10.022599f
C18 VTAIL w_n4910_n4582# 5.62845f
C19 w_n4910_n4582# B 13.363099f
C20 VDD1 w_n4910_n4582# 2.44476f
C21 VDD2 VSUBS 2.50535f
C22 VDD1 VSUBS 3.32344f
C23 VTAIL VSUBS 1.782008f
C24 VN VSUBS 8.28979f
C25 VP VSUBS 4.843283f
C26 B VSUBS 6.642685f
C27 w_n4910_n4582# VSUBS 0.275097p
C28 VDD2.t3 VSUBS 0.446108f
C29 VDD2.t1 VSUBS 0.446108f
C30 VDD2.n0 VSUBS 3.76233f
C31 VDD2.t6 VSUBS 0.446108f
C32 VDD2.t7 VSUBS 0.446108f
C33 VDD2.n1 VSUBS 3.76233f
C34 VDD2.n2 VSUBS 5.95832f
C35 VDD2.t2 VSUBS 0.446108f
C36 VDD2.t4 VSUBS 0.446108f
C37 VDD2.n3 VSUBS 3.73765f
C38 VDD2.n4 VSUBS 5.02472f
C39 VDD2.t0 VSUBS 0.446108f
C40 VDD2.t5 VSUBS 0.446108f
C41 VDD2.n5 VSUBS 3.76227f
C42 VN.t0 VSUBS 3.85429f
C43 VN.n0 VSUBS 1.41121f
C44 VN.n1 VSUBS 0.02148f
C45 VN.n2 VSUBS 0.034947f
C46 VN.n3 VSUBS 0.02148f
C47 VN.n4 VSUBS 0.031336f
C48 VN.n5 VSUBS 0.02148f
C49 VN.n6 VSUBS 0.031356f
C50 VN.n7 VSUBS 0.02148f
C51 VN.n8 VSUBS 0.028964f
C52 VN.t6 VSUBS 3.85429f
C53 VN.n9 VSUBS 1.40216f
C54 VN.t4 VSUBS 4.17485f
C55 VN.n10 VSUBS 1.34057f
C56 VN.n11 VSUBS 0.269044f
C57 VN.n12 VSUBS 0.02148f
C58 VN.n13 VSUBS 0.040032f
C59 VN.n14 VSUBS 0.040032f
C60 VN.n15 VSUBS 0.031356f
C61 VN.n16 VSUBS 0.02148f
C62 VN.n17 VSUBS 0.02148f
C63 VN.n18 VSUBS 0.02148f
C64 VN.n19 VSUBS 0.040032f
C65 VN.n20 VSUBS 0.040032f
C66 VN.t1 VSUBS 3.85429f
C67 VN.n21 VSUBS 1.32867f
C68 VN.n22 VSUBS 0.028964f
C69 VN.n23 VSUBS 0.02148f
C70 VN.n24 VSUBS 0.02148f
C71 VN.n25 VSUBS 0.02148f
C72 VN.n26 VSUBS 0.040032f
C73 VN.n27 VSUBS 0.040032f
C74 VN.n28 VSUBS 0.027765f
C75 VN.n29 VSUBS 0.02148f
C76 VN.n30 VSUBS 0.02148f
C77 VN.n31 VSUBS 0.02148f
C78 VN.n32 VSUBS 0.040032f
C79 VN.n33 VSUBS 0.040032f
C80 VN.n34 VSUBS 0.026593f
C81 VN.n35 VSUBS 0.034667f
C82 VN.n36 VSUBS 0.06046f
C83 VN.t5 VSUBS 3.85429f
C84 VN.n37 VSUBS 1.41121f
C85 VN.n38 VSUBS 0.02148f
C86 VN.n39 VSUBS 0.034947f
C87 VN.n40 VSUBS 0.02148f
C88 VN.n41 VSUBS 0.031336f
C89 VN.n42 VSUBS 0.02148f
C90 VN.t3 VSUBS 3.85429f
C91 VN.n43 VSUBS 1.32867f
C92 VN.n44 VSUBS 0.031356f
C93 VN.n45 VSUBS 0.02148f
C94 VN.n46 VSUBS 0.028964f
C95 VN.t2 VSUBS 4.17485f
C96 VN.t7 VSUBS 3.85429f
C97 VN.n47 VSUBS 1.40216f
C98 VN.n48 VSUBS 1.34057f
C99 VN.n49 VSUBS 0.269044f
C100 VN.n50 VSUBS 0.02148f
C101 VN.n51 VSUBS 0.040032f
C102 VN.n52 VSUBS 0.040032f
C103 VN.n53 VSUBS 0.031356f
C104 VN.n54 VSUBS 0.02148f
C105 VN.n55 VSUBS 0.02148f
C106 VN.n56 VSUBS 0.02148f
C107 VN.n57 VSUBS 0.040032f
C108 VN.n58 VSUBS 0.040032f
C109 VN.n59 VSUBS 0.028964f
C110 VN.n60 VSUBS 0.02148f
C111 VN.n61 VSUBS 0.02148f
C112 VN.n62 VSUBS 0.02148f
C113 VN.n63 VSUBS 0.040032f
C114 VN.n64 VSUBS 0.040032f
C115 VN.n65 VSUBS 0.027765f
C116 VN.n66 VSUBS 0.02148f
C117 VN.n67 VSUBS 0.02148f
C118 VN.n68 VSUBS 0.02148f
C119 VN.n69 VSUBS 0.040032f
C120 VN.n70 VSUBS 0.040032f
C121 VN.n71 VSUBS 0.026593f
C122 VN.n72 VSUBS 0.034667f
C123 VN.n73 VSUBS 1.60049f
C124 VDD1.t6 VSUBS 0.445887f
C125 VDD1.t1 VSUBS 0.445887f
C126 VDD1.n0 VSUBS 3.7624f
C127 VDD1.t2 VSUBS 0.445887f
C128 VDD1.t3 VSUBS 0.445887f
C129 VDD1.n1 VSUBS 3.76046f
C130 VDD1.t4 VSUBS 0.445887f
C131 VDD1.t5 VSUBS 0.445887f
C132 VDD1.n2 VSUBS 3.76046f
C133 VDD1.n3 VSUBS 6.01948f
C134 VDD1.t0 VSUBS 0.445887f
C135 VDD1.t7 VSUBS 0.445887f
C136 VDD1.n4 VSUBS 3.73579f
C137 VDD1.n5 VSUBS 5.061759f
C138 VTAIL.t5 VSUBS 0.345436f
C139 VTAIL.t4 VSUBS 0.345436f
C140 VTAIL.n0 VSUBS 2.75866f
C141 VTAIL.n1 VSUBS 0.82618f
C142 VTAIL.n2 VSUBS 0.013633f
C143 VTAIL.n3 VSUBS 0.030726f
C144 VTAIL.n4 VSUBS 0.013764f
C145 VTAIL.n5 VSUBS 0.024191f
C146 VTAIL.n6 VSUBS 0.012999f
C147 VTAIL.n7 VSUBS 0.030726f
C148 VTAIL.n8 VSUBS 0.013764f
C149 VTAIL.n9 VSUBS 0.024191f
C150 VTAIL.n10 VSUBS 0.012999f
C151 VTAIL.n11 VSUBS 0.030726f
C152 VTAIL.n12 VSUBS 0.013764f
C153 VTAIL.n13 VSUBS 0.024191f
C154 VTAIL.n14 VSUBS 0.012999f
C155 VTAIL.n15 VSUBS 0.030726f
C156 VTAIL.n16 VSUBS 0.013764f
C157 VTAIL.n17 VSUBS 0.024191f
C158 VTAIL.n18 VSUBS 0.012999f
C159 VTAIL.n19 VSUBS 0.030726f
C160 VTAIL.n20 VSUBS 0.013764f
C161 VTAIL.n21 VSUBS 0.024191f
C162 VTAIL.n22 VSUBS 0.012999f
C163 VTAIL.n23 VSUBS 0.030726f
C164 VTAIL.n24 VSUBS 0.013764f
C165 VTAIL.n25 VSUBS 0.024191f
C166 VTAIL.n26 VSUBS 0.012999f
C167 VTAIL.n27 VSUBS 0.030726f
C168 VTAIL.n28 VSUBS 0.013764f
C169 VTAIL.n29 VSUBS 0.024191f
C170 VTAIL.n30 VSUBS 0.012999f
C171 VTAIL.n31 VSUBS 0.030726f
C172 VTAIL.n32 VSUBS 0.013764f
C173 VTAIL.n33 VSUBS 0.256913f
C174 VTAIL.t2 VSUBS 0.066705f
C175 VTAIL.n34 VSUBS 0.023044f
C176 VTAIL.n35 VSUBS 0.023113f
C177 VTAIL.n36 VSUBS 0.012999f
C178 VTAIL.n37 VSUBS 1.83199f
C179 VTAIL.n38 VSUBS 0.024191f
C180 VTAIL.n39 VSUBS 0.012999f
C181 VTAIL.n40 VSUBS 0.013764f
C182 VTAIL.n41 VSUBS 0.030726f
C183 VTAIL.n42 VSUBS 0.030726f
C184 VTAIL.n43 VSUBS 0.013764f
C185 VTAIL.n44 VSUBS 0.012999f
C186 VTAIL.n45 VSUBS 0.024191f
C187 VTAIL.n46 VSUBS 0.024191f
C188 VTAIL.n47 VSUBS 0.012999f
C189 VTAIL.n48 VSUBS 0.013764f
C190 VTAIL.n49 VSUBS 0.030726f
C191 VTAIL.n50 VSUBS 0.030726f
C192 VTAIL.n51 VSUBS 0.030726f
C193 VTAIL.n52 VSUBS 0.013764f
C194 VTAIL.n53 VSUBS 0.012999f
C195 VTAIL.n54 VSUBS 0.024191f
C196 VTAIL.n55 VSUBS 0.024191f
C197 VTAIL.n56 VSUBS 0.012999f
C198 VTAIL.n57 VSUBS 0.013382f
C199 VTAIL.n58 VSUBS 0.013382f
C200 VTAIL.n59 VSUBS 0.030726f
C201 VTAIL.n60 VSUBS 0.030726f
C202 VTAIL.n61 VSUBS 0.013764f
C203 VTAIL.n62 VSUBS 0.012999f
C204 VTAIL.n63 VSUBS 0.024191f
C205 VTAIL.n64 VSUBS 0.024191f
C206 VTAIL.n65 VSUBS 0.012999f
C207 VTAIL.n66 VSUBS 0.013764f
C208 VTAIL.n67 VSUBS 0.030726f
C209 VTAIL.n68 VSUBS 0.030726f
C210 VTAIL.n69 VSUBS 0.013764f
C211 VTAIL.n70 VSUBS 0.012999f
C212 VTAIL.n71 VSUBS 0.024191f
C213 VTAIL.n72 VSUBS 0.024191f
C214 VTAIL.n73 VSUBS 0.012999f
C215 VTAIL.n74 VSUBS 0.013764f
C216 VTAIL.n75 VSUBS 0.030726f
C217 VTAIL.n76 VSUBS 0.030726f
C218 VTAIL.n77 VSUBS 0.013764f
C219 VTAIL.n78 VSUBS 0.012999f
C220 VTAIL.n79 VSUBS 0.024191f
C221 VTAIL.n80 VSUBS 0.024191f
C222 VTAIL.n81 VSUBS 0.012999f
C223 VTAIL.n82 VSUBS 0.013764f
C224 VTAIL.n83 VSUBS 0.030726f
C225 VTAIL.n84 VSUBS 0.030726f
C226 VTAIL.n85 VSUBS 0.013764f
C227 VTAIL.n86 VSUBS 0.012999f
C228 VTAIL.n87 VSUBS 0.024191f
C229 VTAIL.n88 VSUBS 0.024191f
C230 VTAIL.n89 VSUBS 0.012999f
C231 VTAIL.n90 VSUBS 0.013764f
C232 VTAIL.n91 VSUBS 0.030726f
C233 VTAIL.n92 VSUBS 0.030726f
C234 VTAIL.n93 VSUBS 0.013764f
C235 VTAIL.n94 VSUBS 0.012999f
C236 VTAIL.n95 VSUBS 0.024191f
C237 VTAIL.n96 VSUBS 0.062196f
C238 VTAIL.n97 VSUBS 0.012999f
C239 VTAIL.n98 VSUBS 0.013764f
C240 VTAIL.n99 VSUBS 0.068101f
C241 VTAIL.n100 VSUBS 0.045614f
C242 VTAIL.n101 VSUBS 0.324471f
C243 VTAIL.n102 VSUBS 0.013633f
C244 VTAIL.n103 VSUBS 0.030726f
C245 VTAIL.n104 VSUBS 0.013764f
C246 VTAIL.n105 VSUBS 0.024191f
C247 VTAIL.n106 VSUBS 0.012999f
C248 VTAIL.n107 VSUBS 0.030726f
C249 VTAIL.n108 VSUBS 0.013764f
C250 VTAIL.n109 VSUBS 0.024191f
C251 VTAIL.n110 VSUBS 0.012999f
C252 VTAIL.n111 VSUBS 0.030726f
C253 VTAIL.n112 VSUBS 0.013764f
C254 VTAIL.n113 VSUBS 0.024191f
C255 VTAIL.n114 VSUBS 0.012999f
C256 VTAIL.n115 VSUBS 0.030726f
C257 VTAIL.n116 VSUBS 0.013764f
C258 VTAIL.n117 VSUBS 0.024191f
C259 VTAIL.n118 VSUBS 0.012999f
C260 VTAIL.n119 VSUBS 0.030726f
C261 VTAIL.n120 VSUBS 0.013764f
C262 VTAIL.n121 VSUBS 0.024191f
C263 VTAIL.n122 VSUBS 0.012999f
C264 VTAIL.n123 VSUBS 0.030726f
C265 VTAIL.n124 VSUBS 0.013764f
C266 VTAIL.n125 VSUBS 0.024191f
C267 VTAIL.n126 VSUBS 0.012999f
C268 VTAIL.n127 VSUBS 0.030726f
C269 VTAIL.n128 VSUBS 0.013764f
C270 VTAIL.n129 VSUBS 0.024191f
C271 VTAIL.n130 VSUBS 0.012999f
C272 VTAIL.n131 VSUBS 0.030726f
C273 VTAIL.n132 VSUBS 0.013764f
C274 VTAIL.n133 VSUBS 0.256913f
C275 VTAIL.t8 VSUBS 0.066705f
C276 VTAIL.n134 VSUBS 0.023044f
C277 VTAIL.n135 VSUBS 0.023113f
C278 VTAIL.n136 VSUBS 0.012999f
C279 VTAIL.n137 VSUBS 1.83199f
C280 VTAIL.n138 VSUBS 0.024191f
C281 VTAIL.n139 VSUBS 0.012999f
C282 VTAIL.n140 VSUBS 0.013764f
C283 VTAIL.n141 VSUBS 0.030726f
C284 VTAIL.n142 VSUBS 0.030726f
C285 VTAIL.n143 VSUBS 0.013764f
C286 VTAIL.n144 VSUBS 0.012999f
C287 VTAIL.n145 VSUBS 0.024191f
C288 VTAIL.n146 VSUBS 0.024191f
C289 VTAIL.n147 VSUBS 0.012999f
C290 VTAIL.n148 VSUBS 0.013764f
C291 VTAIL.n149 VSUBS 0.030726f
C292 VTAIL.n150 VSUBS 0.030726f
C293 VTAIL.n151 VSUBS 0.030726f
C294 VTAIL.n152 VSUBS 0.013764f
C295 VTAIL.n153 VSUBS 0.012999f
C296 VTAIL.n154 VSUBS 0.024191f
C297 VTAIL.n155 VSUBS 0.024191f
C298 VTAIL.n156 VSUBS 0.012999f
C299 VTAIL.n157 VSUBS 0.013382f
C300 VTAIL.n158 VSUBS 0.013382f
C301 VTAIL.n159 VSUBS 0.030726f
C302 VTAIL.n160 VSUBS 0.030726f
C303 VTAIL.n161 VSUBS 0.013764f
C304 VTAIL.n162 VSUBS 0.012999f
C305 VTAIL.n163 VSUBS 0.024191f
C306 VTAIL.n164 VSUBS 0.024191f
C307 VTAIL.n165 VSUBS 0.012999f
C308 VTAIL.n166 VSUBS 0.013764f
C309 VTAIL.n167 VSUBS 0.030726f
C310 VTAIL.n168 VSUBS 0.030726f
C311 VTAIL.n169 VSUBS 0.013764f
C312 VTAIL.n170 VSUBS 0.012999f
C313 VTAIL.n171 VSUBS 0.024191f
C314 VTAIL.n172 VSUBS 0.024191f
C315 VTAIL.n173 VSUBS 0.012999f
C316 VTAIL.n174 VSUBS 0.013764f
C317 VTAIL.n175 VSUBS 0.030726f
C318 VTAIL.n176 VSUBS 0.030726f
C319 VTAIL.n177 VSUBS 0.013764f
C320 VTAIL.n178 VSUBS 0.012999f
C321 VTAIL.n179 VSUBS 0.024191f
C322 VTAIL.n180 VSUBS 0.024191f
C323 VTAIL.n181 VSUBS 0.012999f
C324 VTAIL.n182 VSUBS 0.013764f
C325 VTAIL.n183 VSUBS 0.030726f
C326 VTAIL.n184 VSUBS 0.030726f
C327 VTAIL.n185 VSUBS 0.013764f
C328 VTAIL.n186 VSUBS 0.012999f
C329 VTAIL.n187 VSUBS 0.024191f
C330 VTAIL.n188 VSUBS 0.024191f
C331 VTAIL.n189 VSUBS 0.012999f
C332 VTAIL.n190 VSUBS 0.013764f
C333 VTAIL.n191 VSUBS 0.030726f
C334 VTAIL.n192 VSUBS 0.030726f
C335 VTAIL.n193 VSUBS 0.013764f
C336 VTAIL.n194 VSUBS 0.012999f
C337 VTAIL.n195 VSUBS 0.024191f
C338 VTAIL.n196 VSUBS 0.062196f
C339 VTAIL.n197 VSUBS 0.012999f
C340 VTAIL.n198 VSUBS 0.013764f
C341 VTAIL.n199 VSUBS 0.068101f
C342 VTAIL.n200 VSUBS 0.045614f
C343 VTAIL.n201 VSUBS 0.324471f
C344 VTAIL.t9 VSUBS 0.345436f
C345 VTAIL.t7 VSUBS 0.345436f
C346 VTAIL.n202 VSUBS 2.75866f
C347 VTAIL.n203 VSUBS 1.0864f
C348 VTAIL.n204 VSUBS 0.013633f
C349 VTAIL.n205 VSUBS 0.030726f
C350 VTAIL.n206 VSUBS 0.013764f
C351 VTAIL.n207 VSUBS 0.024191f
C352 VTAIL.n208 VSUBS 0.012999f
C353 VTAIL.n209 VSUBS 0.030726f
C354 VTAIL.n210 VSUBS 0.013764f
C355 VTAIL.n211 VSUBS 0.024191f
C356 VTAIL.n212 VSUBS 0.012999f
C357 VTAIL.n213 VSUBS 0.030726f
C358 VTAIL.n214 VSUBS 0.013764f
C359 VTAIL.n215 VSUBS 0.024191f
C360 VTAIL.n216 VSUBS 0.012999f
C361 VTAIL.n217 VSUBS 0.030726f
C362 VTAIL.n218 VSUBS 0.013764f
C363 VTAIL.n219 VSUBS 0.024191f
C364 VTAIL.n220 VSUBS 0.012999f
C365 VTAIL.n221 VSUBS 0.030726f
C366 VTAIL.n222 VSUBS 0.013764f
C367 VTAIL.n223 VSUBS 0.024191f
C368 VTAIL.n224 VSUBS 0.012999f
C369 VTAIL.n225 VSUBS 0.030726f
C370 VTAIL.n226 VSUBS 0.013764f
C371 VTAIL.n227 VSUBS 0.024191f
C372 VTAIL.n228 VSUBS 0.012999f
C373 VTAIL.n229 VSUBS 0.030726f
C374 VTAIL.n230 VSUBS 0.013764f
C375 VTAIL.n231 VSUBS 0.024191f
C376 VTAIL.n232 VSUBS 0.012999f
C377 VTAIL.n233 VSUBS 0.030726f
C378 VTAIL.n234 VSUBS 0.013764f
C379 VTAIL.n235 VSUBS 0.256913f
C380 VTAIL.t13 VSUBS 0.066705f
C381 VTAIL.n236 VSUBS 0.023044f
C382 VTAIL.n237 VSUBS 0.023113f
C383 VTAIL.n238 VSUBS 0.012999f
C384 VTAIL.n239 VSUBS 1.83199f
C385 VTAIL.n240 VSUBS 0.024191f
C386 VTAIL.n241 VSUBS 0.012999f
C387 VTAIL.n242 VSUBS 0.013764f
C388 VTAIL.n243 VSUBS 0.030726f
C389 VTAIL.n244 VSUBS 0.030726f
C390 VTAIL.n245 VSUBS 0.013764f
C391 VTAIL.n246 VSUBS 0.012999f
C392 VTAIL.n247 VSUBS 0.024191f
C393 VTAIL.n248 VSUBS 0.024191f
C394 VTAIL.n249 VSUBS 0.012999f
C395 VTAIL.n250 VSUBS 0.013764f
C396 VTAIL.n251 VSUBS 0.030726f
C397 VTAIL.n252 VSUBS 0.030726f
C398 VTAIL.n253 VSUBS 0.030726f
C399 VTAIL.n254 VSUBS 0.013764f
C400 VTAIL.n255 VSUBS 0.012999f
C401 VTAIL.n256 VSUBS 0.024191f
C402 VTAIL.n257 VSUBS 0.024191f
C403 VTAIL.n258 VSUBS 0.012999f
C404 VTAIL.n259 VSUBS 0.013382f
C405 VTAIL.n260 VSUBS 0.013382f
C406 VTAIL.n261 VSUBS 0.030726f
C407 VTAIL.n262 VSUBS 0.030726f
C408 VTAIL.n263 VSUBS 0.013764f
C409 VTAIL.n264 VSUBS 0.012999f
C410 VTAIL.n265 VSUBS 0.024191f
C411 VTAIL.n266 VSUBS 0.024191f
C412 VTAIL.n267 VSUBS 0.012999f
C413 VTAIL.n268 VSUBS 0.013764f
C414 VTAIL.n269 VSUBS 0.030726f
C415 VTAIL.n270 VSUBS 0.030726f
C416 VTAIL.n271 VSUBS 0.013764f
C417 VTAIL.n272 VSUBS 0.012999f
C418 VTAIL.n273 VSUBS 0.024191f
C419 VTAIL.n274 VSUBS 0.024191f
C420 VTAIL.n275 VSUBS 0.012999f
C421 VTAIL.n276 VSUBS 0.013764f
C422 VTAIL.n277 VSUBS 0.030726f
C423 VTAIL.n278 VSUBS 0.030726f
C424 VTAIL.n279 VSUBS 0.013764f
C425 VTAIL.n280 VSUBS 0.012999f
C426 VTAIL.n281 VSUBS 0.024191f
C427 VTAIL.n282 VSUBS 0.024191f
C428 VTAIL.n283 VSUBS 0.012999f
C429 VTAIL.n284 VSUBS 0.013764f
C430 VTAIL.n285 VSUBS 0.030726f
C431 VTAIL.n286 VSUBS 0.030726f
C432 VTAIL.n287 VSUBS 0.013764f
C433 VTAIL.n288 VSUBS 0.012999f
C434 VTAIL.n289 VSUBS 0.024191f
C435 VTAIL.n290 VSUBS 0.024191f
C436 VTAIL.n291 VSUBS 0.012999f
C437 VTAIL.n292 VSUBS 0.013764f
C438 VTAIL.n293 VSUBS 0.030726f
C439 VTAIL.n294 VSUBS 0.030726f
C440 VTAIL.n295 VSUBS 0.013764f
C441 VTAIL.n296 VSUBS 0.012999f
C442 VTAIL.n297 VSUBS 0.024191f
C443 VTAIL.n298 VSUBS 0.062196f
C444 VTAIL.n299 VSUBS 0.012999f
C445 VTAIL.n300 VSUBS 0.013764f
C446 VTAIL.n301 VSUBS 0.068101f
C447 VTAIL.n302 VSUBS 0.045614f
C448 VTAIL.n303 VSUBS 2.09547f
C449 VTAIL.n304 VSUBS 0.013633f
C450 VTAIL.n305 VSUBS 0.030726f
C451 VTAIL.n306 VSUBS 0.013764f
C452 VTAIL.n307 VSUBS 0.024191f
C453 VTAIL.n308 VSUBS 0.012999f
C454 VTAIL.n309 VSUBS 0.030726f
C455 VTAIL.n310 VSUBS 0.013764f
C456 VTAIL.n311 VSUBS 0.024191f
C457 VTAIL.n312 VSUBS 0.012999f
C458 VTAIL.n313 VSUBS 0.030726f
C459 VTAIL.n314 VSUBS 0.013764f
C460 VTAIL.n315 VSUBS 0.024191f
C461 VTAIL.n316 VSUBS 0.012999f
C462 VTAIL.n317 VSUBS 0.030726f
C463 VTAIL.n318 VSUBS 0.013764f
C464 VTAIL.n319 VSUBS 0.024191f
C465 VTAIL.n320 VSUBS 0.012999f
C466 VTAIL.n321 VSUBS 0.030726f
C467 VTAIL.n322 VSUBS 0.013764f
C468 VTAIL.n323 VSUBS 0.024191f
C469 VTAIL.n324 VSUBS 0.012999f
C470 VTAIL.n325 VSUBS 0.030726f
C471 VTAIL.n326 VSUBS 0.013764f
C472 VTAIL.n327 VSUBS 0.024191f
C473 VTAIL.n328 VSUBS 0.012999f
C474 VTAIL.n329 VSUBS 0.030726f
C475 VTAIL.n330 VSUBS 0.030726f
C476 VTAIL.n331 VSUBS 0.013764f
C477 VTAIL.n332 VSUBS 0.024191f
C478 VTAIL.n333 VSUBS 0.012999f
C479 VTAIL.n334 VSUBS 0.030726f
C480 VTAIL.n335 VSUBS 0.013764f
C481 VTAIL.n336 VSUBS 0.256913f
C482 VTAIL.t1 VSUBS 0.066705f
C483 VTAIL.n337 VSUBS 0.023044f
C484 VTAIL.n338 VSUBS 0.023113f
C485 VTAIL.n339 VSUBS 0.012999f
C486 VTAIL.n340 VSUBS 1.83199f
C487 VTAIL.n341 VSUBS 0.024191f
C488 VTAIL.n342 VSUBS 0.012999f
C489 VTAIL.n343 VSUBS 0.013764f
C490 VTAIL.n344 VSUBS 0.030726f
C491 VTAIL.n345 VSUBS 0.030726f
C492 VTAIL.n346 VSUBS 0.013764f
C493 VTAIL.n347 VSUBS 0.012999f
C494 VTAIL.n348 VSUBS 0.024191f
C495 VTAIL.n349 VSUBS 0.024191f
C496 VTAIL.n350 VSUBS 0.012999f
C497 VTAIL.n351 VSUBS 0.013764f
C498 VTAIL.n352 VSUBS 0.030726f
C499 VTAIL.n353 VSUBS 0.030726f
C500 VTAIL.n354 VSUBS 0.013764f
C501 VTAIL.n355 VSUBS 0.012999f
C502 VTAIL.n356 VSUBS 0.024191f
C503 VTAIL.n357 VSUBS 0.024191f
C504 VTAIL.n358 VSUBS 0.012999f
C505 VTAIL.n359 VSUBS 0.013382f
C506 VTAIL.n360 VSUBS 0.013382f
C507 VTAIL.n361 VSUBS 0.030726f
C508 VTAIL.n362 VSUBS 0.030726f
C509 VTAIL.n363 VSUBS 0.013764f
C510 VTAIL.n364 VSUBS 0.012999f
C511 VTAIL.n365 VSUBS 0.024191f
C512 VTAIL.n366 VSUBS 0.024191f
C513 VTAIL.n367 VSUBS 0.012999f
C514 VTAIL.n368 VSUBS 0.013764f
C515 VTAIL.n369 VSUBS 0.030726f
C516 VTAIL.n370 VSUBS 0.030726f
C517 VTAIL.n371 VSUBS 0.013764f
C518 VTAIL.n372 VSUBS 0.012999f
C519 VTAIL.n373 VSUBS 0.024191f
C520 VTAIL.n374 VSUBS 0.024191f
C521 VTAIL.n375 VSUBS 0.012999f
C522 VTAIL.n376 VSUBS 0.013764f
C523 VTAIL.n377 VSUBS 0.030726f
C524 VTAIL.n378 VSUBS 0.030726f
C525 VTAIL.n379 VSUBS 0.013764f
C526 VTAIL.n380 VSUBS 0.012999f
C527 VTAIL.n381 VSUBS 0.024191f
C528 VTAIL.n382 VSUBS 0.024191f
C529 VTAIL.n383 VSUBS 0.012999f
C530 VTAIL.n384 VSUBS 0.013764f
C531 VTAIL.n385 VSUBS 0.030726f
C532 VTAIL.n386 VSUBS 0.030726f
C533 VTAIL.n387 VSUBS 0.013764f
C534 VTAIL.n388 VSUBS 0.012999f
C535 VTAIL.n389 VSUBS 0.024191f
C536 VTAIL.n390 VSUBS 0.024191f
C537 VTAIL.n391 VSUBS 0.012999f
C538 VTAIL.n392 VSUBS 0.013764f
C539 VTAIL.n393 VSUBS 0.030726f
C540 VTAIL.n394 VSUBS 0.030726f
C541 VTAIL.n395 VSUBS 0.013764f
C542 VTAIL.n396 VSUBS 0.012999f
C543 VTAIL.n397 VSUBS 0.024191f
C544 VTAIL.n398 VSUBS 0.062196f
C545 VTAIL.n399 VSUBS 0.012999f
C546 VTAIL.n400 VSUBS 0.013764f
C547 VTAIL.n401 VSUBS 0.068101f
C548 VTAIL.n402 VSUBS 0.045614f
C549 VTAIL.n403 VSUBS 2.09547f
C550 VTAIL.t3 VSUBS 0.345436f
C551 VTAIL.t0 VSUBS 0.345436f
C552 VTAIL.n404 VSUBS 2.75868f
C553 VTAIL.n405 VSUBS 1.08639f
C554 VTAIL.n406 VSUBS 0.013633f
C555 VTAIL.n407 VSUBS 0.030726f
C556 VTAIL.n408 VSUBS 0.013764f
C557 VTAIL.n409 VSUBS 0.024191f
C558 VTAIL.n410 VSUBS 0.012999f
C559 VTAIL.n411 VSUBS 0.030726f
C560 VTAIL.n412 VSUBS 0.013764f
C561 VTAIL.n413 VSUBS 0.024191f
C562 VTAIL.n414 VSUBS 0.012999f
C563 VTAIL.n415 VSUBS 0.030726f
C564 VTAIL.n416 VSUBS 0.013764f
C565 VTAIL.n417 VSUBS 0.024191f
C566 VTAIL.n418 VSUBS 0.012999f
C567 VTAIL.n419 VSUBS 0.030726f
C568 VTAIL.n420 VSUBS 0.013764f
C569 VTAIL.n421 VSUBS 0.024191f
C570 VTAIL.n422 VSUBS 0.012999f
C571 VTAIL.n423 VSUBS 0.030726f
C572 VTAIL.n424 VSUBS 0.013764f
C573 VTAIL.n425 VSUBS 0.024191f
C574 VTAIL.n426 VSUBS 0.012999f
C575 VTAIL.n427 VSUBS 0.030726f
C576 VTAIL.n428 VSUBS 0.013764f
C577 VTAIL.n429 VSUBS 0.024191f
C578 VTAIL.n430 VSUBS 0.012999f
C579 VTAIL.n431 VSUBS 0.030726f
C580 VTAIL.n432 VSUBS 0.030726f
C581 VTAIL.n433 VSUBS 0.013764f
C582 VTAIL.n434 VSUBS 0.024191f
C583 VTAIL.n435 VSUBS 0.012999f
C584 VTAIL.n436 VSUBS 0.030726f
C585 VTAIL.n437 VSUBS 0.013764f
C586 VTAIL.n438 VSUBS 0.256913f
C587 VTAIL.t6 VSUBS 0.066705f
C588 VTAIL.n439 VSUBS 0.023044f
C589 VTAIL.n440 VSUBS 0.023113f
C590 VTAIL.n441 VSUBS 0.012999f
C591 VTAIL.n442 VSUBS 1.83199f
C592 VTAIL.n443 VSUBS 0.024191f
C593 VTAIL.n444 VSUBS 0.012999f
C594 VTAIL.n445 VSUBS 0.013764f
C595 VTAIL.n446 VSUBS 0.030726f
C596 VTAIL.n447 VSUBS 0.030726f
C597 VTAIL.n448 VSUBS 0.013764f
C598 VTAIL.n449 VSUBS 0.012999f
C599 VTAIL.n450 VSUBS 0.024191f
C600 VTAIL.n451 VSUBS 0.024191f
C601 VTAIL.n452 VSUBS 0.012999f
C602 VTAIL.n453 VSUBS 0.013764f
C603 VTAIL.n454 VSUBS 0.030726f
C604 VTAIL.n455 VSUBS 0.030726f
C605 VTAIL.n456 VSUBS 0.013764f
C606 VTAIL.n457 VSUBS 0.012999f
C607 VTAIL.n458 VSUBS 0.024191f
C608 VTAIL.n459 VSUBS 0.024191f
C609 VTAIL.n460 VSUBS 0.012999f
C610 VTAIL.n461 VSUBS 0.013382f
C611 VTAIL.n462 VSUBS 0.013382f
C612 VTAIL.n463 VSUBS 0.030726f
C613 VTAIL.n464 VSUBS 0.030726f
C614 VTAIL.n465 VSUBS 0.013764f
C615 VTAIL.n466 VSUBS 0.012999f
C616 VTAIL.n467 VSUBS 0.024191f
C617 VTAIL.n468 VSUBS 0.024191f
C618 VTAIL.n469 VSUBS 0.012999f
C619 VTAIL.n470 VSUBS 0.013764f
C620 VTAIL.n471 VSUBS 0.030726f
C621 VTAIL.n472 VSUBS 0.030726f
C622 VTAIL.n473 VSUBS 0.013764f
C623 VTAIL.n474 VSUBS 0.012999f
C624 VTAIL.n475 VSUBS 0.024191f
C625 VTAIL.n476 VSUBS 0.024191f
C626 VTAIL.n477 VSUBS 0.012999f
C627 VTAIL.n478 VSUBS 0.013764f
C628 VTAIL.n479 VSUBS 0.030726f
C629 VTAIL.n480 VSUBS 0.030726f
C630 VTAIL.n481 VSUBS 0.013764f
C631 VTAIL.n482 VSUBS 0.012999f
C632 VTAIL.n483 VSUBS 0.024191f
C633 VTAIL.n484 VSUBS 0.024191f
C634 VTAIL.n485 VSUBS 0.012999f
C635 VTAIL.n486 VSUBS 0.013764f
C636 VTAIL.n487 VSUBS 0.030726f
C637 VTAIL.n488 VSUBS 0.030726f
C638 VTAIL.n489 VSUBS 0.013764f
C639 VTAIL.n490 VSUBS 0.012999f
C640 VTAIL.n491 VSUBS 0.024191f
C641 VTAIL.n492 VSUBS 0.024191f
C642 VTAIL.n493 VSUBS 0.012999f
C643 VTAIL.n494 VSUBS 0.013764f
C644 VTAIL.n495 VSUBS 0.030726f
C645 VTAIL.n496 VSUBS 0.030726f
C646 VTAIL.n497 VSUBS 0.013764f
C647 VTAIL.n498 VSUBS 0.012999f
C648 VTAIL.n499 VSUBS 0.024191f
C649 VTAIL.n500 VSUBS 0.062196f
C650 VTAIL.n501 VSUBS 0.012999f
C651 VTAIL.n502 VSUBS 0.013764f
C652 VTAIL.n503 VSUBS 0.068101f
C653 VTAIL.n504 VSUBS 0.045614f
C654 VTAIL.n505 VSUBS 0.324471f
C655 VTAIL.n506 VSUBS 0.013633f
C656 VTAIL.n507 VSUBS 0.030726f
C657 VTAIL.n508 VSUBS 0.013764f
C658 VTAIL.n509 VSUBS 0.024191f
C659 VTAIL.n510 VSUBS 0.012999f
C660 VTAIL.n511 VSUBS 0.030726f
C661 VTAIL.n512 VSUBS 0.013764f
C662 VTAIL.n513 VSUBS 0.024191f
C663 VTAIL.n514 VSUBS 0.012999f
C664 VTAIL.n515 VSUBS 0.030726f
C665 VTAIL.n516 VSUBS 0.013764f
C666 VTAIL.n517 VSUBS 0.024191f
C667 VTAIL.n518 VSUBS 0.012999f
C668 VTAIL.n519 VSUBS 0.030726f
C669 VTAIL.n520 VSUBS 0.013764f
C670 VTAIL.n521 VSUBS 0.024191f
C671 VTAIL.n522 VSUBS 0.012999f
C672 VTAIL.n523 VSUBS 0.030726f
C673 VTAIL.n524 VSUBS 0.013764f
C674 VTAIL.n525 VSUBS 0.024191f
C675 VTAIL.n526 VSUBS 0.012999f
C676 VTAIL.n527 VSUBS 0.030726f
C677 VTAIL.n528 VSUBS 0.013764f
C678 VTAIL.n529 VSUBS 0.024191f
C679 VTAIL.n530 VSUBS 0.012999f
C680 VTAIL.n531 VSUBS 0.030726f
C681 VTAIL.n532 VSUBS 0.030726f
C682 VTAIL.n533 VSUBS 0.013764f
C683 VTAIL.n534 VSUBS 0.024191f
C684 VTAIL.n535 VSUBS 0.012999f
C685 VTAIL.n536 VSUBS 0.030726f
C686 VTAIL.n537 VSUBS 0.013764f
C687 VTAIL.n538 VSUBS 0.256913f
C688 VTAIL.t12 VSUBS 0.066705f
C689 VTAIL.n539 VSUBS 0.023044f
C690 VTAIL.n540 VSUBS 0.023113f
C691 VTAIL.n541 VSUBS 0.012999f
C692 VTAIL.n542 VSUBS 1.83199f
C693 VTAIL.n543 VSUBS 0.024191f
C694 VTAIL.n544 VSUBS 0.012999f
C695 VTAIL.n545 VSUBS 0.013764f
C696 VTAIL.n546 VSUBS 0.030726f
C697 VTAIL.n547 VSUBS 0.030726f
C698 VTAIL.n548 VSUBS 0.013764f
C699 VTAIL.n549 VSUBS 0.012999f
C700 VTAIL.n550 VSUBS 0.024191f
C701 VTAIL.n551 VSUBS 0.024191f
C702 VTAIL.n552 VSUBS 0.012999f
C703 VTAIL.n553 VSUBS 0.013764f
C704 VTAIL.n554 VSUBS 0.030726f
C705 VTAIL.n555 VSUBS 0.030726f
C706 VTAIL.n556 VSUBS 0.013764f
C707 VTAIL.n557 VSUBS 0.012999f
C708 VTAIL.n558 VSUBS 0.024191f
C709 VTAIL.n559 VSUBS 0.024191f
C710 VTAIL.n560 VSUBS 0.012999f
C711 VTAIL.n561 VSUBS 0.013382f
C712 VTAIL.n562 VSUBS 0.013382f
C713 VTAIL.n563 VSUBS 0.030726f
C714 VTAIL.n564 VSUBS 0.030726f
C715 VTAIL.n565 VSUBS 0.013764f
C716 VTAIL.n566 VSUBS 0.012999f
C717 VTAIL.n567 VSUBS 0.024191f
C718 VTAIL.n568 VSUBS 0.024191f
C719 VTAIL.n569 VSUBS 0.012999f
C720 VTAIL.n570 VSUBS 0.013764f
C721 VTAIL.n571 VSUBS 0.030726f
C722 VTAIL.n572 VSUBS 0.030726f
C723 VTAIL.n573 VSUBS 0.013764f
C724 VTAIL.n574 VSUBS 0.012999f
C725 VTAIL.n575 VSUBS 0.024191f
C726 VTAIL.n576 VSUBS 0.024191f
C727 VTAIL.n577 VSUBS 0.012999f
C728 VTAIL.n578 VSUBS 0.013764f
C729 VTAIL.n579 VSUBS 0.030726f
C730 VTAIL.n580 VSUBS 0.030726f
C731 VTAIL.n581 VSUBS 0.013764f
C732 VTAIL.n582 VSUBS 0.012999f
C733 VTAIL.n583 VSUBS 0.024191f
C734 VTAIL.n584 VSUBS 0.024191f
C735 VTAIL.n585 VSUBS 0.012999f
C736 VTAIL.n586 VSUBS 0.013764f
C737 VTAIL.n587 VSUBS 0.030726f
C738 VTAIL.n588 VSUBS 0.030726f
C739 VTAIL.n589 VSUBS 0.013764f
C740 VTAIL.n590 VSUBS 0.012999f
C741 VTAIL.n591 VSUBS 0.024191f
C742 VTAIL.n592 VSUBS 0.024191f
C743 VTAIL.n593 VSUBS 0.012999f
C744 VTAIL.n594 VSUBS 0.013764f
C745 VTAIL.n595 VSUBS 0.030726f
C746 VTAIL.n596 VSUBS 0.030726f
C747 VTAIL.n597 VSUBS 0.013764f
C748 VTAIL.n598 VSUBS 0.012999f
C749 VTAIL.n599 VSUBS 0.024191f
C750 VTAIL.n600 VSUBS 0.062196f
C751 VTAIL.n601 VSUBS 0.012999f
C752 VTAIL.n602 VSUBS 0.013764f
C753 VTAIL.n603 VSUBS 0.068101f
C754 VTAIL.n604 VSUBS 0.045614f
C755 VTAIL.n605 VSUBS 0.324471f
C756 VTAIL.t14 VSUBS 0.345436f
C757 VTAIL.t11 VSUBS 0.345436f
C758 VTAIL.n606 VSUBS 2.75868f
C759 VTAIL.n607 VSUBS 1.08639f
C760 VTAIL.n608 VSUBS 0.013633f
C761 VTAIL.n609 VSUBS 0.030726f
C762 VTAIL.n610 VSUBS 0.013764f
C763 VTAIL.n611 VSUBS 0.024191f
C764 VTAIL.n612 VSUBS 0.012999f
C765 VTAIL.n613 VSUBS 0.030726f
C766 VTAIL.n614 VSUBS 0.013764f
C767 VTAIL.n615 VSUBS 0.024191f
C768 VTAIL.n616 VSUBS 0.012999f
C769 VTAIL.n617 VSUBS 0.030726f
C770 VTAIL.n618 VSUBS 0.013764f
C771 VTAIL.n619 VSUBS 0.024191f
C772 VTAIL.n620 VSUBS 0.012999f
C773 VTAIL.n621 VSUBS 0.030726f
C774 VTAIL.n622 VSUBS 0.013764f
C775 VTAIL.n623 VSUBS 0.024191f
C776 VTAIL.n624 VSUBS 0.012999f
C777 VTAIL.n625 VSUBS 0.030726f
C778 VTAIL.n626 VSUBS 0.013764f
C779 VTAIL.n627 VSUBS 0.024191f
C780 VTAIL.n628 VSUBS 0.012999f
C781 VTAIL.n629 VSUBS 0.030726f
C782 VTAIL.n630 VSUBS 0.013764f
C783 VTAIL.n631 VSUBS 0.024191f
C784 VTAIL.n632 VSUBS 0.012999f
C785 VTAIL.n633 VSUBS 0.030726f
C786 VTAIL.n634 VSUBS 0.030726f
C787 VTAIL.n635 VSUBS 0.013764f
C788 VTAIL.n636 VSUBS 0.024191f
C789 VTAIL.n637 VSUBS 0.012999f
C790 VTAIL.n638 VSUBS 0.030726f
C791 VTAIL.n639 VSUBS 0.013764f
C792 VTAIL.n640 VSUBS 0.256913f
C793 VTAIL.t10 VSUBS 0.066705f
C794 VTAIL.n641 VSUBS 0.023044f
C795 VTAIL.n642 VSUBS 0.023113f
C796 VTAIL.n643 VSUBS 0.012999f
C797 VTAIL.n644 VSUBS 1.83199f
C798 VTAIL.n645 VSUBS 0.024191f
C799 VTAIL.n646 VSUBS 0.012999f
C800 VTAIL.n647 VSUBS 0.013764f
C801 VTAIL.n648 VSUBS 0.030726f
C802 VTAIL.n649 VSUBS 0.030726f
C803 VTAIL.n650 VSUBS 0.013764f
C804 VTAIL.n651 VSUBS 0.012999f
C805 VTAIL.n652 VSUBS 0.024191f
C806 VTAIL.n653 VSUBS 0.024191f
C807 VTAIL.n654 VSUBS 0.012999f
C808 VTAIL.n655 VSUBS 0.013764f
C809 VTAIL.n656 VSUBS 0.030726f
C810 VTAIL.n657 VSUBS 0.030726f
C811 VTAIL.n658 VSUBS 0.013764f
C812 VTAIL.n659 VSUBS 0.012999f
C813 VTAIL.n660 VSUBS 0.024191f
C814 VTAIL.n661 VSUBS 0.024191f
C815 VTAIL.n662 VSUBS 0.012999f
C816 VTAIL.n663 VSUBS 0.013382f
C817 VTAIL.n664 VSUBS 0.013382f
C818 VTAIL.n665 VSUBS 0.030726f
C819 VTAIL.n666 VSUBS 0.030726f
C820 VTAIL.n667 VSUBS 0.013764f
C821 VTAIL.n668 VSUBS 0.012999f
C822 VTAIL.n669 VSUBS 0.024191f
C823 VTAIL.n670 VSUBS 0.024191f
C824 VTAIL.n671 VSUBS 0.012999f
C825 VTAIL.n672 VSUBS 0.013764f
C826 VTAIL.n673 VSUBS 0.030726f
C827 VTAIL.n674 VSUBS 0.030726f
C828 VTAIL.n675 VSUBS 0.013764f
C829 VTAIL.n676 VSUBS 0.012999f
C830 VTAIL.n677 VSUBS 0.024191f
C831 VTAIL.n678 VSUBS 0.024191f
C832 VTAIL.n679 VSUBS 0.012999f
C833 VTAIL.n680 VSUBS 0.013764f
C834 VTAIL.n681 VSUBS 0.030726f
C835 VTAIL.n682 VSUBS 0.030726f
C836 VTAIL.n683 VSUBS 0.013764f
C837 VTAIL.n684 VSUBS 0.012999f
C838 VTAIL.n685 VSUBS 0.024191f
C839 VTAIL.n686 VSUBS 0.024191f
C840 VTAIL.n687 VSUBS 0.012999f
C841 VTAIL.n688 VSUBS 0.013764f
C842 VTAIL.n689 VSUBS 0.030726f
C843 VTAIL.n690 VSUBS 0.030726f
C844 VTAIL.n691 VSUBS 0.013764f
C845 VTAIL.n692 VSUBS 0.012999f
C846 VTAIL.n693 VSUBS 0.024191f
C847 VTAIL.n694 VSUBS 0.024191f
C848 VTAIL.n695 VSUBS 0.012999f
C849 VTAIL.n696 VSUBS 0.013764f
C850 VTAIL.n697 VSUBS 0.030726f
C851 VTAIL.n698 VSUBS 0.030726f
C852 VTAIL.n699 VSUBS 0.013764f
C853 VTAIL.n700 VSUBS 0.012999f
C854 VTAIL.n701 VSUBS 0.024191f
C855 VTAIL.n702 VSUBS 0.062196f
C856 VTAIL.n703 VSUBS 0.012999f
C857 VTAIL.n704 VSUBS 0.013764f
C858 VTAIL.n705 VSUBS 0.068101f
C859 VTAIL.n706 VSUBS 0.045614f
C860 VTAIL.n707 VSUBS 2.09547f
C861 VTAIL.n708 VSUBS 0.013633f
C862 VTAIL.n709 VSUBS 0.030726f
C863 VTAIL.n710 VSUBS 0.013764f
C864 VTAIL.n711 VSUBS 0.024191f
C865 VTAIL.n712 VSUBS 0.012999f
C866 VTAIL.n713 VSUBS 0.030726f
C867 VTAIL.n714 VSUBS 0.013764f
C868 VTAIL.n715 VSUBS 0.024191f
C869 VTAIL.n716 VSUBS 0.012999f
C870 VTAIL.n717 VSUBS 0.030726f
C871 VTAIL.n718 VSUBS 0.013764f
C872 VTAIL.n719 VSUBS 0.024191f
C873 VTAIL.n720 VSUBS 0.012999f
C874 VTAIL.n721 VSUBS 0.030726f
C875 VTAIL.n722 VSUBS 0.013764f
C876 VTAIL.n723 VSUBS 0.024191f
C877 VTAIL.n724 VSUBS 0.012999f
C878 VTAIL.n725 VSUBS 0.030726f
C879 VTAIL.n726 VSUBS 0.013764f
C880 VTAIL.n727 VSUBS 0.024191f
C881 VTAIL.n728 VSUBS 0.012999f
C882 VTAIL.n729 VSUBS 0.030726f
C883 VTAIL.n730 VSUBS 0.013764f
C884 VTAIL.n731 VSUBS 0.024191f
C885 VTAIL.n732 VSUBS 0.012999f
C886 VTAIL.n733 VSUBS 0.030726f
C887 VTAIL.n734 VSUBS 0.013764f
C888 VTAIL.n735 VSUBS 0.024191f
C889 VTAIL.n736 VSUBS 0.012999f
C890 VTAIL.n737 VSUBS 0.030726f
C891 VTAIL.n738 VSUBS 0.013764f
C892 VTAIL.n739 VSUBS 0.256913f
C893 VTAIL.t15 VSUBS 0.066705f
C894 VTAIL.n740 VSUBS 0.023044f
C895 VTAIL.n741 VSUBS 0.023113f
C896 VTAIL.n742 VSUBS 0.012999f
C897 VTAIL.n743 VSUBS 1.83199f
C898 VTAIL.n744 VSUBS 0.024191f
C899 VTAIL.n745 VSUBS 0.012999f
C900 VTAIL.n746 VSUBS 0.013764f
C901 VTAIL.n747 VSUBS 0.030726f
C902 VTAIL.n748 VSUBS 0.030726f
C903 VTAIL.n749 VSUBS 0.013764f
C904 VTAIL.n750 VSUBS 0.012999f
C905 VTAIL.n751 VSUBS 0.024191f
C906 VTAIL.n752 VSUBS 0.024191f
C907 VTAIL.n753 VSUBS 0.012999f
C908 VTAIL.n754 VSUBS 0.013764f
C909 VTAIL.n755 VSUBS 0.030726f
C910 VTAIL.n756 VSUBS 0.030726f
C911 VTAIL.n757 VSUBS 0.030726f
C912 VTAIL.n758 VSUBS 0.013764f
C913 VTAIL.n759 VSUBS 0.012999f
C914 VTAIL.n760 VSUBS 0.024191f
C915 VTAIL.n761 VSUBS 0.024191f
C916 VTAIL.n762 VSUBS 0.012999f
C917 VTAIL.n763 VSUBS 0.013382f
C918 VTAIL.n764 VSUBS 0.013382f
C919 VTAIL.n765 VSUBS 0.030726f
C920 VTAIL.n766 VSUBS 0.030726f
C921 VTAIL.n767 VSUBS 0.013764f
C922 VTAIL.n768 VSUBS 0.012999f
C923 VTAIL.n769 VSUBS 0.024191f
C924 VTAIL.n770 VSUBS 0.024191f
C925 VTAIL.n771 VSUBS 0.012999f
C926 VTAIL.n772 VSUBS 0.013764f
C927 VTAIL.n773 VSUBS 0.030726f
C928 VTAIL.n774 VSUBS 0.030726f
C929 VTAIL.n775 VSUBS 0.013764f
C930 VTAIL.n776 VSUBS 0.012999f
C931 VTAIL.n777 VSUBS 0.024191f
C932 VTAIL.n778 VSUBS 0.024191f
C933 VTAIL.n779 VSUBS 0.012999f
C934 VTAIL.n780 VSUBS 0.013764f
C935 VTAIL.n781 VSUBS 0.030726f
C936 VTAIL.n782 VSUBS 0.030726f
C937 VTAIL.n783 VSUBS 0.013764f
C938 VTAIL.n784 VSUBS 0.012999f
C939 VTAIL.n785 VSUBS 0.024191f
C940 VTAIL.n786 VSUBS 0.024191f
C941 VTAIL.n787 VSUBS 0.012999f
C942 VTAIL.n788 VSUBS 0.013764f
C943 VTAIL.n789 VSUBS 0.030726f
C944 VTAIL.n790 VSUBS 0.030726f
C945 VTAIL.n791 VSUBS 0.013764f
C946 VTAIL.n792 VSUBS 0.012999f
C947 VTAIL.n793 VSUBS 0.024191f
C948 VTAIL.n794 VSUBS 0.024191f
C949 VTAIL.n795 VSUBS 0.012999f
C950 VTAIL.n796 VSUBS 0.013764f
C951 VTAIL.n797 VSUBS 0.030726f
C952 VTAIL.n798 VSUBS 0.030726f
C953 VTAIL.n799 VSUBS 0.013764f
C954 VTAIL.n800 VSUBS 0.012999f
C955 VTAIL.n801 VSUBS 0.024191f
C956 VTAIL.n802 VSUBS 0.062196f
C957 VTAIL.n803 VSUBS 0.012999f
C958 VTAIL.n804 VSUBS 0.013764f
C959 VTAIL.n805 VSUBS 0.068101f
C960 VTAIL.n806 VSUBS 0.045614f
C961 VTAIL.n807 VSUBS 2.09094f
C962 VP.t2 VSUBS 4.16204f
C963 VP.n0 VSUBS 1.52389f
C964 VP.n1 VSUBS 0.023194f
C965 VP.n2 VSUBS 0.037738f
C966 VP.n3 VSUBS 0.023194f
C967 VP.n4 VSUBS 0.033838f
C968 VP.n5 VSUBS 0.023194f
C969 VP.n6 VSUBS 0.03386f
C970 VP.n7 VSUBS 0.023194f
C971 VP.n8 VSUBS 0.031277f
C972 VP.n9 VSUBS 0.023194f
C973 VP.n10 VSUBS 0.029982f
C974 VP.n11 VSUBS 0.023194f
C975 VP.n12 VSUBS 0.028716f
C976 VP.t0 VSUBS 4.16204f
C977 VP.n13 VSUBS 1.52389f
C978 VP.n14 VSUBS 0.023194f
C979 VP.n15 VSUBS 0.037738f
C980 VP.n16 VSUBS 0.023194f
C981 VP.n17 VSUBS 0.033838f
C982 VP.n18 VSUBS 0.023194f
C983 VP.n19 VSUBS 0.03386f
C984 VP.n20 VSUBS 0.023194f
C985 VP.n21 VSUBS 0.031277f
C986 VP.t1 VSUBS 4.5082f
C987 VP.t6 VSUBS 4.16204f
C988 VP.n22 VSUBS 1.51411f
C989 VP.n23 VSUBS 1.44761f
C990 VP.n24 VSUBS 0.290527f
C991 VP.n25 VSUBS 0.023194f
C992 VP.n26 VSUBS 0.043229f
C993 VP.n27 VSUBS 0.043229f
C994 VP.n28 VSUBS 0.03386f
C995 VP.n29 VSUBS 0.023194f
C996 VP.n30 VSUBS 0.023194f
C997 VP.n31 VSUBS 0.023194f
C998 VP.n32 VSUBS 0.043229f
C999 VP.n33 VSUBS 0.043229f
C1000 VP.t7 VSUBS 4.16204f
C1001 VP.n34 VSUBS 1.43476f
C1002 VP.n35 VSUBS 0.031277f
C1003 VP.n36 VSUBS 0.023194f
C1004 VP.n37 VSUBS 0.023194f
C1005 VP.n38 VSUBS 0.023194f
C1006 VP.n39 VSUBS 0.043229f
C1007 VP.n40 VSUBS 0.043229f
C1008 VP.n41 VSUBS 0.029982f
C1009 VP.n42 VSUBS 0.023194f
C1010 VP.n43 VSUBS 0.023194f
C1011 VP.n44 VSUBS 0.023194f
C1012 VP.n45 VSUBS 0.043229f
C1013 VP.n46 VSUBS 0.043229f
C1014 VP.n47 VSUBS 0.028716f
C1015 VP.n48 VSUBS 0.037436f
C1016 VP.n49 VSUBS 1.71935f
C1017 VP.t5 VSUBS 4.16204f
C1018 VP.n50 VSUBS 1.52389f
C1019 VP.n51 VSUBS 1.73318f
C1020 VP.n52 VSUBS 0.037436f
C1021 VP.n53 VSUBS 0.023194f
C1022 VP.n54 VSUBS 0.043229f
C1023 VP.n55 VSUBS 0.043229f
C1024 VP.n56 VSUBS 0.037738f
C1025 VP.n57 VSUBS 0.023194f
C1026 VP.n58 VSUBS 0.023194f
C1027 VP.n59 VSUBS 0.023194f
C1028 VP.n60 VSUBS 0.043229f
C1029 VP.n61 VSUBS 0.043229f
C1030 VP.t4 VSUBS 4.16204f
C1031 VP.n62 VSUBS 1.43476f
C1032 VP.n63 VSUBS 0.033838f
C1033 VP.n64 VSUBS 0.023194f
C1034 VP.n65 VSUBS 0.023194f
C1035 VP.n66 VSUBS 0.023194f
C1036 VP.n67 VSUBS 0.043229f
C1037 VP.n68 VSUBS 0.043229f
C1038 VP.n69 VSUBS 0.03386f
C1039 VP.n70 VSUBS 0.023194f
C1040 VP.n71 VSUBS 0.023194f
C1041 VP.n72 VSUBS 0.023194f
C1042 VP.n73 VSUBS 0.043229f
C1043 VP.n74 VSUBS 0.043229f
C1044 VP.t3 VSUBS 4.16204f
C1045 VP.n75 VSUBS 1.43476f
C1046 VP.n76 VSUBS 0.031277f
C1047 VP.n77 VSUBS 0.023194f
C1048 VP.n78 VSUBS 0.023194f
C1049 VP.n79 VSUBS 0.023194f
C1050 VP.n80 VSUBS 0.043229f
C1051 VP.n81 VSUBS 0.043229f
C1052 VP.n82 VSUBS 0.029982f
C1053 VP.n83 VSUBS 0.023194f
C1054 VP.n84 VSUBS 0.023194f
C1055 VP.n85 VSUBS 0.023194f
C1056 VP.n86 VSUBS 0.043229f
C1057 VP.n87 VSUBS 0.043229f
C1058 VP.n88 VSUBS 0.028716f
C1059 VP.n89 VSUBS 0.037436f
C1060 VP.n90 VSUBS 0.065288f
C1061 B.n0 VSUBS 0.004689f
C1062 B.n1 VSUBS 0.004689f
C1063 B.n2 VSUBS 0.007415f
C1064 B.n3 VSUBS 0.007415f
C1065 B.n4 VSUBS 0.007415f
C1066 B.n5 VSUBS 0.007415f
C1067 B.n6 VSUBS 0.007415f
C1068 B.n7 VSUBS 0.007415f
C1069 B.n8 VSUBS 0.007415f
C1070 B.n9 VSUBS 0.007415f
C1071 B.n10 VSUBS 0.007415f
C1072 B.n11 VSUBS 0.007415f
C1073 B.n12 VSUBS 0.007415f
C1074 B.n13 VSUBS 0.007415f
C1075 B.n14 VSUBS 0.007415f
C1076 B.n15 VSUBS 0.007415f
C1077 B.n16 VSUBS 0.007415f
C1078 B.n17 VSUBS 0.007415f
C1079 B.n18 VSUBS 0.007415f
C1080 B.n19 VSUBS 0.007415f
C1081 B.n20 VSUBS 0.007415f
C1082 B.n21 VSUBS 0.007415f
C1083 B.n22 VSUBS 0.007415f
C1084 B.n23 VSUBS 0.007415f
C1085 B.n24 VSUBS 0.007415f
C1086 B.n25 VSUBS 0.007415f
C1087 B.n26 VSUBS 0.007415f
C1088 B.n27 VSUBS 0.007415f
C1089 B.n28 VSUBS 0.007415f
C1090 B.n29 VSUBS 0.007415f
C1091 B.n30 VSUBS 0.007415f
C1092 B.n31 VSUBS 0.007415f
C1093 B.n32 VSUBS 0.007415f
C1094 B.n33 VSUBS 0.007415f
C1095 B.n34 VSUBS 0.007415f
C1096 B.n35 VSUBS 0.01725f
C1097 B.n36 VSUBS 0.007415f
C1098 B.n37 VSUBS 0.007415f
C1099 B.n38 VSUBS 0.007415f
C1100 B.n39 VSUBS 0.007415f
C1101 B.n40 VSUBS 0.007415f
C1102 B.n41 VSUBS 0.007415f
C1103 B.n42 VSUBS 0.007415f
C1104 B.n43 VSUBS 0.007415f
C1105 B.n44 VSUBS 0.007415f
C1106 B.n45 VSUBS 0.007415f
C1107 B.n46 VSUBS 0.007415f
C1108 B.n47 VSUBS 0.007415f
C1109 B.n48 VSUBS 0.007415f
C1110 B.n49 VSUBS 0.007415f
C1111 B.n50 VSUBS 0.007415f
C1112 B.n51 VSUBS 0.007415f
C1113 B.n52 VSUBS 0.007415f
C1114 B.n53 VSUBS 0.007415f
C1115 B.n54 VSUBS 0.007415f
C1116 B.n55 VSUBS 0.007415f
C1117 B.n56 VSUBS 0.007415f
C1118 B.n57 VSUBS 0.007415f
C1119 B.n58 VSUBS 0.007415f
C1120 B.n59 VSUBS 0.007415f
C1121 B.n60 VSUBS 0.007415f
C1122 B.n61 VSUBS 0.007415f
C1123 B.n62 VSUBS 0.007415f
C1124 B.n63 VSUBS 0.007415f
C1125 B.n64 VSUBS 0.007415f
C1126 B.n65 VSUBS 0.007415f
C1127 B.t2 VSUBS 0.373481f
C1128 B.t1 VSUBS 0.4202f
C1129 B.t0 VSUBS 3.137f
C1130 B.n66 VSUBS 0.669523f
C1131 B.n67 VSUBS 0.353696f
C1132 B.n68 VSUBS 0.007415f
C1133 B.n69 VSUBS 0.007415f
C1134 B.n70 VSUBS 0.007415f
C1135 B.n71 VSUBS 0.007415f
C1136 B.t11 VSUBS 0.373485f
C1137 B.t10 VSUBS 0.420203f
C1138 B.t9 VSUBS 3.137f
C1139 B.n72 VSUBS 0.66952f
C1140 B.n73 VSUBS 0.353693f
C1141 B.n74 VSUBS 0.007415f
C1142 B.n75 VSUBS 0.007415f
C1143 B.n76 VSUBS 0.007415f
C1144 B.n77 VSUBS 0.007415f
C1145 B.n78 VSUBS 0.007415f
C1146 B.n79 VSUBS 0.007415f
C1147 B.n80 VSUBS 0.007415f
C1148 B.n81 VSUBS 0.007415f
C1149 B.n82 VSUBS 0.007415f
C1150 B.n83 VSUBS 0.007415f
C1151 B.n84 VSUBS 0.007415f
C1152 B.n85 VSUBS 0.007415f
C1153 B.n86 VSUBS 0.007415f
C1154 B.n87 VSUBS 0.007415f
C1155 B.n88 VSUBS 0.007415f
C1156 B.n89 VSUBS 0.007415f
C1157 B.n90 VSUBS 0.007415f
C1158 B.n91 VSUBS 0.007415f
C1159 B.n92 VSUBS 0.007415f
C1160 B.n93 VSUBS 0.007415f
C1161 B.n94 VSUBS 0.007415f
C1162 B.n95 VSUBS 0.007415f
C1163 B.n96 VSUBS 0.007415f
C1164 B.n97 VSUBS 0.007415f
C1165 B.n98 VSUBS 0.007415f
C1166 B.n99 VSUBS 0.007415f
C1167 B.n100 VSUBS 0.007415f
C1168 B.n101 VSUBS 0.007415f
C1169 B.n102 VSUBS 0.007415f
C1170 B.n103 VSUBS 0.01725f
C1171 B.n104 VSUBS 0.007415f
C1172 B.n105 VSUBS 0.007415f
C1173 B.n106 VSUBS 0.007415f
C1174 B.n107 VSUBS 0.007415f
C1175 B.n108 VSUBS 0.007415f
C1176 B.n109 VSUBS 0.007415f
C1177 B.n110 VSUBS 0.007415f
C1178 B.n111 VSUBS 0.007415f
C1179 B.n112 VSUBS 0.007415f
C1180 B.n113 VSUBS 0.007415f
C1181 B.n114 VSUBS 0.007415f
C1182 B.n115 VSUBS 0.007415f
C1183 B.n116 VSUBS 0.007415f
C1184 B.n117 VSUBS 0.007415f
C1185 B.n118 VSUBS 0.007415f
C1186 B.n119 VSUBS 0.007415f
C1187 B.n120 VSUBS 0.007415f
C1188 B.n121 VSUBS 0.007415f
C1189 B.n122 VSUBS 0.007415f
C1190 B.n123 VSUBS 0.007415f
C1191 B.n124 VSUBS 0.007415f
C1192 B.n125 VSUBS 0.007415f
C1193 B.n126 VSUBS 0.007415f
C1194 B.n127 VSUBS 0.007415f
C1195 B.n128 VSUBS 0.007415f
C1196 B.n129 VSUBS 0.007415f
C1197 B.n130 VSUBS 0.007415f
C1198 B.n131 VSUBS 0.007415f
C1199 B.n132 VSUBS 0.007415f
C1200 B.n133 VSUBS 0.007415f
C1201 B.n134 VSUBS 0.007415f
C1202 B.n135 VSUBS 0.007415f
C1203 B.n136 VSUBS 0.007415f
C1204 B.n137 VSUBS 0.007415f
C1205 B.n138 VSUBS 0.007415f
C1206 B.n139 VSUBS 0.007415f
C1207 B.n140 VSUBS 0.007415f
C1208 B.n141 VSUBS 0.007415f
C1209 B.n142 VSUBS 0.007415f
C1210 B.n143 VSUBS 0.007415f
C1211 B.n144 VSUBS 0.007415f
C1212 B.n145 VSUBS 0.007415f
C1213 B.n146 VSUBS 0.007415f
C1214 B.n147 VSUBS 0.007415f
C1215 B.n148 VSUBS 0.007415f
C1216 B.n149 VSUBS 0.007415f
C1217 B.n150 VSUBS 0.007415f
C1218 B.n151 VSUBS 0.007415f
C1219 B.n152 VSUBS 0.007415f
C1220 B.n153 VSUBS 0.007415f
C1221 B.n154 VSUBS 0.007415f
C1222 B.n155 VSUBS 0.007415f
C1223 B.n156 VSUBS 0.007415f
C1224 B.n157 VSUBS 0.007415f
C1225 B.n158 VSUBS 0.007415f
C1226 B.n159 VSUBS 0.007415f
C1227 B.n160 VSUBS 0.007415f
C1228 B.n161 VSUBS 0.007415f
C1229 B.n162 VSUBS 0.007415f
C1230 B.n163 VSUBS 0.007415f
C1231 B.n164 VSUBS 0.007415f
C1232 B.n165 VSUBS 0.007415f
C1233 B.n166 VSUBS 0.007415f
C1234 B.n167 VSUBS 0.007415f
C1235 B.n168 VSUBS 0.007415f
C1236 B.n169 VSUBS 0.007415f
C1237 B.n170 VSUBS 0.01725f
C1238 B.n171 VSUBS 0.007415f
C1239 B.n172 VSUBS 0.007415f
C1240 B.n173 VSUBS 0.007415f
C1241 B.n174 VSUBS 0.007415f
C1242 B.n175 VSUBS 0.007415f
C1243 B.n176 VSUBS 0.007415f
C1244 B.n177 VSUBS 0.007415f
C1245 B.n178 VSUBS 0.007415f
C1246 B.n179 VSUBS 0.007415f
C1247 B.n180 VSUBS 0.007415f
C1248 B.n181 VSUBS 0.007415f
C1249 B.n182 VSUBS 0.007415f
C1250 B.n183 VSUBS 0.007415f
C1251 B.n184 VSUBS 0.007415f
C1252 B.n185 VSUBS 0.007415f
C1253 B.n186 VSUBS 0.007415f
C1254 B.n187 VSUBS 0.007415f
C1255 B.n188 VSUBS 0.007415f
C1256 B.n189 VSUBS 0.007415f
C1257 B.n190 VSUBS 0.007415f
C1258 B.n191 VSUBS 0.007415f
C1259 B.n192 VSUBS 0.007415f
C1260 B.n193 VSUBS 0.007415f
C1261 B.n194 VSUBS 0.007415f
C1262 B.n195 VSUBS 0.007415f
C1263 B.n196 VSUBS 0.007415f
C1264 B.n197 VSUBS 0.007415f
C1265 B.n198 VSUBS 0.007415f
C1266 B.n199 VSUBS 0.007415f
C1267 B.t7 VSUBS 0.373485f
C1268 B.t8 VSUBS 0.420203f
C1269 B.t6 VSUBS 3.137f
C1270 B.n200 VSUBS 0.66952f
C1271 B.n201 VSUBS 0.353693f
C1272 B.n202 VSUBS 0.017179f
C1273 B.n203 VSUBS 0.007415f
C1274 B.n204 VSUBS 0.007415f
C1275 B.n205 VSUBS 0.007415f
C1276 B.n206 VSUBS 0.007415f
C1277 B.n207 VSUBS 0.007415f
C1278 B.t4 VSUBS 0.373481f
C1279 B.t5 VSUBS 0.4202f
C1280 B.t3 VSUBS 3.137f
C1281 B.n208 VSUBS 0.669523f
C1282 B.n209 VSUBS 0.353696f
C1283 B.n210 VSUBS 0.007415f
C1284 B.n211 VSUBS 0.007415f
C1285 B.n212 VSUBS 0.007415f
C1286 B.n213 VSUBS 0.007415f
C1287 B.n214 VSUBS 0.007415f
C1288 B.n215 VSUBS 0.007415f
C1289 B.n216 VSUBS 0.007415f
C1290 B.n217 VSUBS 0.007415f
C1291 B.n218 VSUBS 0.007415f
C1292 B.n219 VSUBS 0.007415f
C1293 B.n220 VSUBS 0.007415f
C1294 B.n221 VSUBS 0.007415f
C1295 B.n222 VSUBS 0.007415f
C1296 B.n223 VSUBS 0.007415f
C1297 B.n224 VSUBS 0.007415f
C1298 B.n225 VSUBS 0.007415f
C1299 B.n226 VSUBS 0.007415f
C1300 B.n227 VSUBS 0.007415f
C1301 B.n228 VSUBS 0.007415f
C1302 B.n229 VSUBS 0.007415f
C1303 B.n230 VSUBS 0.007415f
C1304 B.n231 VSUBS 0.007415f
C1305 B.n232 VSUBS 0.007415f
C1306 B.n233 VSUBS 0.007415f
C1307 B.n234 VSUBS 0.007415f
C1308 B.n235 VSUBS 0.007415f
C1309 B.n236 VSUBS 0.007415f
C1310 B.n237 VSUBS 0.007415f
C1311 B.n238 VSUBS 0.007415f
C1312 B.n239 VSUBS 0.015898f
C1313 B.n240 VSUBS 0.007415f
C1314 B.n241 VSUBS 0.007415f
C1315 B.n242 VSUBS 0.007415f
C1316 B.n243 VSUBS 0.007415f
C1317 B.n244 VSUBS 0.007415f
C1318 B.n245 VSUBS 0.007415f
C1319 B.n246 VSUBS 0.007415f
C1320 B.n247 VSUBS 0.007415f
C1321 B.n248 VSUBS 0.007415f
C1322 B.n249 VSUBS 0.007415f
C1323 B.n250 VSUBS 0.007415f
C1324 B.n251 VSUBS 0.007415f
C1325 B.n252 VSUBS 0.007415f
C1326 B.n253 VSUBS 0.007415f
C1327 B.n254 VSUBS 0.007415f
C1328 B.n255 VSUBS 0.007415f
C1329 B.n256 VSUBS 0.007415f
C1330 B.n257 VSUBS 0.007415f
C1331 B.n258 VSUBS 0.007415f
C1332 B.n259 VSUBS 0.007415f
C1333 B.n260 VSUBS 0.007415f
C1334 B.n261 VSUBS 0.007415f
C1335 B.n262 VSUBS 0.007415f
C1336 B.n263 VSUBS 0.007415f
C1337 B.n264 VSUBS 0.007415f
C1338 B.n265 VSUBS 0.007415f
C1339 B.n266 VSUBS 0.007415f
C1340 B.n267 VSUBS 0.007415f
C1341 B.n268 VSUBS 0.007415f
C1342 B.n269 VSUBS 0.007415f
C1343 B.n270 VSUBS 0.007415f
C1344 B.n271 VSUBS 0.007415f
C1345 B.n272 VSUBS 0.007415f
C1346 B.n273 VSUBS 0.007415f
C1347 B.n274 VSUBS 0.007415f
C1348 B.n275 VSUBS 0.007415f
C1349 B.n276 VSUBS 0.007415f
C1350 B.n277 VSUBS 0.007415f
C1351 B.n278 VSUBS 0.007415f
C1352 B.n279 VSUBS 0.007415f
C1353 B.n280 VSUBS 0.007415f
C1354 B.n281 VSUBS 0.007415f
C1355 B.n282 VSUBS 0.007415f
C1356 B.n283 VSUBS 0.007415f
C1357 B.n284 VSUBS 0.007415f
C1358 B.n285 VSUBS 0.007415f
C1359 B.n286 VSUBS 0.007415f
C1360 B.n287 VSUBS 0.007415f
C1361 B.n288 VSUBS 0.007415f
C1362 B.n289 VSUBS 0.007415f
C1363 B.n290 VSUBS 0.007415f
C1364 B.n291 VSUBS 0.007415f
C1365 B.n292 VSUBS 0.007415f
C1366 B.n293 VSUBS 0.007415f
C1367 B.n294 VSUBS 0.007415f
C1368 B.n295 VSUBS 0.007415f
C1369 B.n296 VSUBS 0.007415f
C1370 B.n297 VSUBS 0.007415f
C1371 B.n298 VSUBS 0.007415f
C1372 B.n299 VSUBS 0.007415f
C1373 B.n300 VSUBS 0.007415f
C1374 B.n301 VSUBS 0.007415f
C1375 B.n302 VSUBS 0.007415f
C1376 B.n303 VSUBS 0.007415f
C1377 B.n304 VSUBS 0.007415f
C1378 B.n305 VSUBS 0.007415f
C1379 B.n306 VSUBS 0.007415f
C1380 B.n307 VSUBS 0.007415f
C1381 B.n308 VSUBS 0.007415f
C1382 B.n309 VSUBS 0.007415f
C1383 B.n310 VSUBS 0.007415f
C1384 B.n311 VSUBS 0.007415f
C1385 B.n312 VSUBS 0.007415f
C1386 B.n313 VSUBS 0.007415f
C1387 B.n314 VSUBS 0.007415f
C1388 B.n315 VSUBS 0.007415f
C1389 B.n316 VSUBS 0.007415f
C1390 B.n317 VSUBS 0.007415f
C1391 B.n318 VSUBS 0.007415f
C1392 B.n319 VSUBS 0.007415f
C1393 B.n320 VSUBS 0.007415f
C1394 B.n321 VSUBS 0.007415f
C1395 B.n322 VSUBS 0.007415f
C1396 B.n323 VSUBS 0.007415f
C1397 B.n324 VSUBS 0.007415f
C1398 B.n325 VSUBS 0.007415f
C1399 B.n326 VSUBS 0.007415f
C1400 B.n327 VSUBS 0.007415f
C1401 B.n328 VSUBS 0.007415f
C1402 B.n329 VSUBS 0.007415f
C1403 B.n330 VSUBS 0.007415f
C1404 B.n331 VSUBS 0.007415f
C1405 B.n332 VSUBS 0.007415f
C1406 B.n333 VSUBS 0.007415f
C1407 B.n334 VSUBS 0.007415f
C1408 B.n335 VSUBS 0.007415f
C1409 B.n336 VSUBS 0.007415f
C1410 B.n337 VSUBS 0.007415f
C1411 B.n338 VSUBS 0.007415f
C1412 B.n339 VSUBS 0.007415f
C1413 B.n340 VSUBS 0.007415f
C1414 B.n341 VSUBS 0.007415f
C1415 B.n342 VSUBS 0.007415f
C1416 B.n343 VSUBS 0.007415f
C1417 B.n344 VSUBS 0.007415f
C1418 B.n345 VSUBS 0.007415f
C1419 B.n346 VSUBS 0.007415f
C1420 B.n347 VSUBS 0.007415f
C1421 B.n348 VSUBS 0.007415f
C1422 B.n349 VSUBS 0.007415f
C1423 B.n350 VSUBS 0.007415f
C1424 B.n351 VSUBS 0.007415f
C1425 B.n352 VSUBS 0.007415f
C1426 B.n353 VSUBS 0.007415f
C1427 B.n354 VSUBS 0.007415f
C1428 B.n355 VSUBS 0.007415f
C1429 B.n356 VSUBS 0.007415f
C1430 B.n357 VSUBS 0.007415f
C1431 B.n358 VSUBS 0.007415f
C1432 B.n359 VSUBS 0.007415f
C1433 B.n360 VSUBS 0.007415f
C1434 B.n361 VSUBS 0.007415f
C1435 B.n362 VSUBS 0.007415f
C1436 B.n363 VSUBS 0.007415f
C1437 B.n364 VSUBS 0.007415f
C1438 B.n365 VSUBS 0.007415f
C1439 B.n366 VSUBS 0.007415f
C1440 B.n367 VSUBS 0.007415f
C1441 B.n368 VSUBS 0.015898f
C1442 B.n369 VSUBS 0.01725f
C1443 B.n370 VSUBS 0.01725f
C1444 B.n371 VSUBS 0.007415f
C1445 B.n372 VSUBS 0.007415f
C1446 B.n373 VSUBS 0.007415f
C1447 B.n374 VSUBS 0.007415f
C1448 B.n375 VSUBS 0.007415f
C1449 B.n376 VSUBS 0.007415f
C1450 B.n377 VSUBS 0.007415f
C1451 B.n378 VSUBS 0.007415f
C1452 B.n379 VSUBS 0.007415f
C1453 B.n380 VSUBS 0.007415f
C1454 B.n381 VSUBS 0.007415f
C1455 B.n382 VSUBS 0.007415f
C1456 B.n383 VSUBS 0.007415f
C1457 B.n384 VSUBS 0.007415f
C1458 B.n385 VSUBS 0.007415f
C1459 B.n386 VSUBS 0.007415f
C1460 B.n387 VSUBS 0.007415f
C1461 B.n388 VSUBS 0.007415f
C1462 B.n389 VSUBS 0.007415f
C1463 B.n390 VSUBS 0.007415f
C1464 B.n391 VSUBS 0.007415f
C1465 B.n392 VSUBS 0.007415f
C1466 B.n393 VSUBS 0.007415f
C1467 B.n394 VSUBS 0.007415f
C1468 B.n395 VSUBS 0.007415f
C1469 B.n396 VSUBS 0.007415f
C1470 B.n397 VSUBS 0.007415f
C1471 B.n398 VSUBS 0.007415f
C1472 B.n399 VSUBS 0.007415f
C1473 B.n400 VSUBS 0.007415f
C1474 B.n401 VSUBS 0.007415f
C1475 B.n402 VSUBS 0.007415f
C1476 B.n403 VSUBS 0.007415f
C1477 B.n404 VSUBS 0.007415f
C1478 B.n405 VSUBS 0.007415f
C1479 B.n406 VSUBS 0.007415f
C1480 B.n407 VSUBS 0.007415f
C1481 B.n408 VSUBS 0.007415f
C1482 B.n409 VSUBS 0.007415f
C1483 B.n410 VSUBS 0.007415f
C1484 B.n411 VSUBS 0.007415f
C1485 B.n412 VSUBS 0.007415f
C1486 B.n413 VSUBS 0.007415f
C1487 B.n414 VSUBS 0.007415f
C1488 B.n415 VSUBS 0.007415f
C1489 B.n416 VSUBS 0.007415f
C1490 B.n417 VSUBS 0.007415f
C1491 B.n418 VSUBS 0.007415f
C1492 B.n419 VSUBS 0.007415f
C1493 B.n420 VSUBS 0.007415f
C1494 B.n421 VSUBS 0.007415f
C1495 B.n422 VSUBS 0.007415f
C1496 B.n423 VSUBS 0.007415f
C1497 B.n424 VSUBS 0.007415f
C1498 B.n425 VSUBS 0.007415f
C1499 B.n426 VSUBS 0.007415f
C1500 B.n427 VSUBS 0.007415f
C1501 B.n428 VSUBS 0.007415f
C1502 B.n429 VSUBS 0.007415f
C1503 B.n430 VSUBS 0.007415f
C1504 B.n431 VSUBS 0.007415f
C1505 B.n432 VSUBS 0.007415f
C1506 B.n433 VSUBS 0.007415f
C1507 B.n434 VSUBS 0.007415f
C1508 B.n435 VSUBS 0.007415f
C1509 B.n436 VSUBS 0.007415f
C1510 B.n437 VSUBS 0.007415f
C1511 B.n438 VSUBS 0.007415f
C1512 B.n439 VSUBS 0.007415f
C1513 B.n440 VSUBS 0.007415f
C1514 B.n441 VSUBS 0.007415f
C1515 B.n442 VSUBS 0.007415f
C1516 B.n443 VSUBS 0.007415f
C1517 B.n444 VSUBS 0.007415f
C1518 B.n445 VSUBS 0.007415f
C1519 B.n446 VSUBS 0.007415f
C1520 B.n447 VSUBS 0.007415f
C1521 B.n448 VSUBS 0.007415f
C1522 B.n449 VSUBS 0.007415f
C1523 B.n450 VSUBS 0.007415f
C1524 B.n451 VSUBS 0.007415f
C1525 B.n452 VSUBS 0.007415f
C1526 B.n453 VSUBS 0.007415f
C1527 B.n454 VSUBS 0.007415f
C1528 B.n455 VSUBS 0.007415f
C1529 B.n456 VSUBS 0.007415f
C1530 B.n457 VSUBS 0.007415f
C1531 B.n458 VSUBS 0.005125f
C1532 B.n459 VSUBS 0.017179f
C1533 B.n460 VSUBS 0.005997f
C1534 B.n461 VSUBS 0.007415f
C1535 B.n462 VSUBS 0.007415f
C1536 B.n463 VSUBS 0.007415f
C1537 B.n464 VSUBS 0.007415f
C1538 B.n465 VSUBS 0.007415f
C1539 B.n466 VSUBS 0.007415f
C1540 B.n467 VSUBS 0.007415f
C1541 B.n468 VSUBS 0.007415f
C1542 B.n469 VSUBS 0.007415f
C1543 B.n470 VSUBS 0.007415f
C1544 B.n471 VSUBS 0.007415f
C1545 B.n472 VSUBS 0.005997f
C1546 B.n473 VSUBS 0.007415f
C1547 B.n474 VSUBS 0.007415f
C1548 B.n475 VSUBS 0.005125f
C1549 B.n476 VSUBS 0.007415f
C1550 B.n477 VSUBS 0.007415f
C1551 B.n478 VSUBS 0.007415f
C1552 B.n479 VSUBS 0.007415f
C1553 B.n480 VSUBS 0.007415f
C1554 B.n481 VSUBS 0.007415f
C1555 B.n482 VSUBS 0.007415f
C1556 B.n483 VSUBS 0.007415f
C1557 B.n484 VSUBS 0.007415f
C1558 B.n485 VSUBS 0.007415f
C1559 B.n486 VSUBS 0.007415f
C1560 B.n487 VSUBS 0.007415f
C1561 B.n488 VSUBS 0.007415f
C1562 B.n489 VSUBS 0.007415f
C1563 B.n490 VSUBS 0.007415f
C1564 B.n491 VSUBS 0.007415f
C1565 B.n492 VSUBS 0.007415f
C1566 B.n493 VSUBS 0.007415f
C1567 B.n494 VSUBS 0.007415f
C1568 B.n495 VSUBS 0.007415f
C1569 B.n496 VSUBS 0.007415f
C1570 B.n497 VSUBS 0.007415f
C1571 B.n498 VSUBS 0.007415f
C1572 B.n499 VSUBS 0.007415f
C1573 B.n500 VSUBS 0.007415f
C1574 B.n501 VSUBS 0.007415f
C1575 B.n502 VSUBS 0.007415f
C1576 B.n503 VSUBS 0.007415f
C1577 B.n504 VSUBS 0.007415f
C1578 B.n505 VSUBS 0.007415f
C1579 B.n506 VSUBS 0.007415f
C1580 B.n507 VSUBS 0.007415f
C1581 B.n508 VSUBS 0.007415f
C1582 B.n509 VSUBS 0.007415f
C1583 B.n510 VSUBS 0.007415f
C1584 B.n511 VSUBS 0.007415f
C1585 B.n512 VSUBS 0.007415f
C1586 B.n513 VSUBS 0.007415f
C1587 B.n514 VSUBS 0.007415f
C1588 B.n515 VSUBS 0.007415f
C1589 B.n516 VSUBS 0.007415f
C1590 B.n517 VSUBS 0.007415f
C1591 B.n518 VSUBS 0.007415f
C1592 B.n519 VSUBS 0.007415f
C1593 B.n520 VSUBS 0.007415f
C1594 B.n521 VSUBS 0.007415f
C1595 B.n522 VSUBS 0.007415f
C1596 B.n523 VSUBS 0.007415f
C1597 B.n524 VSUBS 0.007415f
C1598 B.n525 VSUBS 0.007415f
C1599 B.n526 VSUBS 0.007415f
C1600 B.n527 VSUBS 0.007415f
C1601 B.n528 VSUBS 0.007415f
C1602 B.n529 VSUBS 0.007415f
C1603 B.n530 VSUBS 0.007415f
C1604 B.n531 VSUBS 0.007415f
C1605 B.n532 VSUBS 0.007415f
C1606 B.n533 VSUBS 0.007415f
C1607 B.n534 VSUBS 0.007415f
C1608 B.n535 VSUBS 0.007415f
C1609 B.n536 VSUBS 0.007415f
C1610 B.n537 VSUBS 0.007415f
C1611 B.n538 VSUBS 0.007415f
C1612 B.n539 VSUBS 0.007415f
C1613 B.n540 VSUBS 0.007415f
C1614 B.n541 VSUBS 0.007415f
C1615 B.n542 VSUBS 0.007415f
C1616 B.n543 VSUBS 0.007415f
C1617 B.n544 VSUBS 0.007415f
C1618 B.n545 VSUBS 0.007415f
C1619 B.n546 VSUBS 0.007415f
C1620 B.n547 VSUBS 0.007415f
C1621 B.n548 VSUBS 0.007415f
C1622 B.n549 VSUBS 0.007415f
C1623 B.n550 VSUBS 0.007415f
C1624 B.n551 VSUBS 0.007415f
C1625 B.n552 VSUBS 0.007415f
C1626 B.n553 VSUBS 0.007415f
C1627 B.n554 VSUBS 0.007415f
C1628 B.n555 VSUBS 0.007415f
C1629 B.n556 VSUBS 0.007415f
C1630 B.n557 VSUBS 0.007415f
C1631 B.n558 VSUBS 0.007415f
C1632 B.n559 VSUBS 0.007415f
C1633 B.n560 VSUBS 0.007415f
C1634 B.n561 VSUBS 0.007415f
C1635 B.n562 VSUBS 0.007415f
C1636 B.n563 VSUBS 0.01725f
C1637 B.n564 VSUBS 0.015898f
C1638 B.n565 VSUBS 0.015898f
C1639 B.n566 VSUBS 0.007415f
C1640 B.n567 VSUBS 0.007415f
C1641 B.n568 VSUBS 0.007415f
C1642 B.n569 VSUBS 0.007415f
C1643 B.n570 VSUBS 0.007415f
C1644 B.n571 VSUBS 0.007415f
C1645 B.n572 VSUBS 0.007415f
C1646 B.n573 VSUBS 0.007415f
C1647 B.n574 VSUBS 0.007415f
C1648 B.n575 VSUBS 0.007415f
C1649 B.n576 VSUBS 0.007415f
C1650 B.n577 VSUBS 0.007415f
C1651 B.n578 VSUBS 0.007415f
C1652 B.n579 VSUBS 0.007415f
C1653 B.n580 VSUBS 0.007415f
C1654 B.n581 VSUBS 0.007415f
C1655 B.n582 VSUBS 0.007415f
C1656 B.n583 VSUBS 0.007415f
C1657 B.n584 VSUBS 0.007415f
C1658 B.n585 VSUBS 0.007415f
C1659 B.n586 VSUBS 0.007415f
C1660 B.n587 VSUBS 0.007415f
C1661 B.n588 VSUBS 0.007415f
C1662 B.n589 VSUBS 0.007415f
C1663 B.n590 VSUBS 0.007415f
C1664 B.n591 VSUBS 0.007415f
C1665 B.n592 VSUBS 0.007415f
C1666 B.n593 VSUBS 0.007415f
C1667 B.n594 VSUBS 0.007415f
C1668 B.n595 VSUBS 0.007415f
C1669 B.n596 VSUBS 0.007415f
C1670 B.n597 VSUBS 0.007415f
C1671 B.n598 VSUBS 0.007415f
C1672 B.n599 VSUBS 0.007415f
C1673 B.n600 VSUBS 0.007415f
C1674 B.n601 VSUBS 0.007415f
C1675 B.n602 VSUBS 0.007415f
C1676 B.n603 VSUBS 0.007415f
C1677 B.n604 VSUBS 0.007415f
C1678 B.n605 VSUBS 0.007415f
C1679 B.n606 VSUBS 0.007415f
C1680 B.n607 VSUBS 0.007415f
C1681 B.n608 VSUBS 0.007415f
C1682 B.n609 VSUBS 0.007415f
C1683 B.n610 VSUBS 0.007415f
C1684 B.n611 VSUBS 0.007415f
C1685 B.n612 VSUBS 0.007415f
C1686 B.n613 VSUBS 0.007415f
C1687 B.n614 VSUBS 0.007415f
C1688 B.n615 VSUBS 0.007415f
C1689 B.n616 VSUBS 0.007415f
C1690 B.n617 VSUBS 0.007415f
C1691 B.n618 VSUBS 0.007415f
C1692 B.n619 VSUBS 0.007415f
C1693 B.n620 VSUBS 0.007415f
C1694 B.n621 VSUBS 0.007415f
C1695 B.n622 VSUBS 0.007415f
C1696 B.n623 VSUBS 0.007415f
C1697 B.n624 VSUBS 0.007415f
C1698 B.n625 VSUBS 0.007415f
C1699 B.n626 VSUBS 0.007415f
C1700 B.n627 VSUBS 0.007415f
C1701 B.n628 VSUBS 0.007415f
C1702 B.n629 VSUBS 0.007415f
C1703 B.n630 VSUBS 0.007415f
C1704 B.n631 VSUBS 0.007415f
C1705 B.n632 VSUBS 0.007415f
C1706 B.n633 VSUBS 0.007415f
C1707 B.n634 VSUBS 0.007415f
C1708 B.n635 VSUBS 0.007415f
C1709 B.n636 VSUBS 0.007415f
C1710 B.n637 VSUBS 0.007415f
C1711 B.n638 VSUBS 0.007415f
C1712 B.n639 VSUBS 0.007415f
C1713 B.n640 VSUBS 0.007415f
C1714 B.n641 VSUBS 0.007415f
C1715 B.n642 VSUBS 0.007415f
C1716 B.n643 VSUBS 0.007415f
C1717 B.n644 VSUBS 0.007415f
C1718 B.n645 VSUBS 0.007415f
C1719 B.n646 VSUBS 0.007415f
C1720 B.n647 VSUBS 0.007415f
C1721 B.n648 VSUBS 0.007415f
C1722 B.n649 VSUBS 0.007415f
C1723 B.n650 VSUBS 0.007415f
C1724 B.n651 VSUBS 0.007415f
C1725 B.n652 VSUBS 0.007415f
C1726 B.n653 VSUBS 0.007415f
C1727 B.n654 VSUBS 0.007415f
C1728 B.n655 VSUBS 0.007415f
C1729 B.n656 VSUBS 0.007415f
C1730 B.n657 VSUBS 0.007415f
C1731 B.n658 VSUBS 0.007415f
C1732 B.n659 VSUBS 0.007415f
C1733 B.n660 VSUBS 0.007415f
C1734 B.n661 VSUBS 0.007415f
C1735 B.n662 VSUBS 0.007415f
C1736 B.n663 VSUBS 0.007415f
C1737 B.n664 VSUBS 0.007415f
C1738 B.n665 VSUBS 0.007415f
C1739 B.n666 VSUBS 0.007415f
C1740 B.n667 VSUBS 0.007415f
C1741 B.n668 VSUBS 0.007415f
C1742 B.n669 VSUBS 0.007415f
C1743 B.n670 VSUBS 0.007415f
C1744 B.n671 VSUBS 0.007415f
C1745 B.n672 VSUBS 0.007415f
C1746 B.n673 VSUBS 0.007415f
C1747 B.n674 VSUBS 0.007415f
C1748 B.n675 VSUBS 0.007415f
C1749 B.n676 VSUBS 0.007415f
C1750 B.n677 VSUBS 0.007415f
C1751 B.n678 VSUBS 0.007415f
C1752 B.n679 VSUBS 0.007415f
C1753 B.n680 VSUBS 0.007415f
C1754 B.n681 VSUBS 0.007415f
C1755 B.n682 VSUBS 0.007415f
C1756 B.n683 VSUBS 0.007415f
C1757 B.n684 VSUBS 0.007415f
C1758 B.n685 VSUBS 0.007415f
C1759 B.n686 VSUBS 0.007415f
C1760 B.n687 VSUBS 0.007415f
C1761 B.n688 VSUBS 0.007415f
C1762 B.n689 VSUBS 0.007415f
C1763 B.n690 VSUBS 0.007415f
C1764 B.n691 VSUBS 0.007415f
C1765 B.n692 VSUBS 0.007415f
C1766 B.n693 VSUBS 0.007415f
C1767 B.n694 VSUBS 0.007415f
C1768 B.n695 VSUBS 0.007415f
C1769 B.n696 VSUBS 0.007415f
C1770 B.n697 VSUBS 0.007415f
C1771 B.n698 VSUBS 0.007415f
C1772 B.n699 VSUBS 0.007415f
C1773 B.n700 VSUBS 0.007415f
C1774 B.n701 VSUBS 0.007415f
C1775 B.n702 VSUBS 0.007415f
C1776 B.n703 VSUBS 0.007415f
C1777 B.n704 VSUBS 0.007415f
C1778 B.n705 VSUBS 0.007415f
C1779 B.n706 VSUBS 0.007415f
C1780 B.n707 VSUBS 0.007415f
C1781 B.n708 VSUBS 0.007415f
C1782 B.n709 VSUBS 0.007415f
C1783 B.n710 VSUBS 0.007415f
C1784 B.n711 VSUBS 0.007415f
C1785 B.n712 VSUBS 0.007415f
C1786 B.n713 VSUBS 0.007415f
C1787 B.n714 VSUBS 0.007415f
C1788 B.n715 VSUBS 0.007415f
C1789 B.n716 VSUBS 0.007415f
C1790 B.n717 VSUBS 0.007415f
C1791 B.n718 VSUBS 0.007415f
C1792 B.n719 VSUBS 0.007415f
C1793 B.n720 VSUBS 0.007415f
C1794 B.n721 VSUBS 0.007415f
C1795 B.n722 VSUBS 0.007415f
C1796 B.n723 VSUBS 0.007415f
C1797 B.n724 VSUBS 0.007415f
C1798 B.n725 VSUBS 0.007415f
C1799 B.n726 VSUBS 0.007415f
C1800 B.n727 VSUBS 0.007415f
C1801 B.n728 VSUBS 0.007415f
C1802 B.n729 VSUBS 0.007415f
C1803 B.n730 VSUBS 0.007415f
C1804 B.n731 VSUBS 0.007415f
C1805 B.n732 VSUBS 0.007415f
C1806 B.n733 VSUBS 0.007415f
C1807 B.n734 VSUBS 0.007415f
C1808 B.n735 VSUBS 0.007415f
C1809 B.n736 VSUBS 0.007415f
C1810 B.n737 VSUBS 0.007415f
C1811 B.n738 VSUBS 0.007415f
C1812 B.n739 VSUBS 0.007415f
C1813 B.n740 VSUBS 0.007415f
C1814 B.n741 VSUBS 0.007415f
C1815 B.n742 VSUBS 0.007415f
C1816 B.n743 VSUBS 0.007415f
C1817 B.n744 VSUBS 0.007415f
C1818 B.n745 VSUBS 0.007415f
C1819 B.n746 VSUBS 0.007415f
C1820 B.n747 VSUBS 0.007415f
C1821 B.n748 VSUBS 0.007415f
C1822 B.n749 VSUBS 0.007415f
C1823 B.n750 VSUBS 0.007415f
C1824 B.n751 VSUBS 0.007415f
C1825 B.n752 VSUBS 0.007415f
C1826 B.n753 VSUBS 0.007415f
C1827 B.n754 VSUBS 0.007415f
C1828 B.n755 VSUBS 0.007415f
C1829 B.n756 VSUBS 0.007415f
C1830 B.n757 VSUBS 0.007415f
C1831 B.n758 VSUBS 0.007415f
C1832 B.n759 VSUBS 0.007415f
C1833 B.n760 VSUBS 0.007415f
C1834 B.n761 VSUBS 0.007415f
C1835 B.n762 VSUBS 0.015898f
C1836 B.n763 VSUBS 0.016838f
C1837 B.n764 VSUBS 0.01631f
C1838 B.n765 VSUBS 0.007415f
C1839 B.n766 VSUBS 0.007415f
C1840 B.n767 VSUBS 0.007415f
C1841 B.n768 VSUBS 0.007415f
C1842 B.n769 VSUBS 0.007415f
C1843 B.n770 VSUBS 0.007415f
C1844 B.n771 VSUBS 0.007415f
C1845 B.n772 VSUBS 0.007415f
C1846 B.n773 VSUBS 0.007415f
C1847 B.n774 VSUBS 0.007415f
C1848 B.n775 VSUBS 0.007415f
C1849 B.n776 VSUBS 0.007415f
C1850 B.n777 VSUBS 0.007415f
C1851 B.n778 VSUBS 0.007415f
C1852 B.n779 VSUBS 0.007415f
C1853 B.n780 VSUBS 0.007415f
C1854 B.n781 VSUBS 0.007415f
C1855 B.n782 VSUBS 0.007415f
C1856 B.n783 VSUBS 0.007415f
C1857 B.n784 VSUBS 0.007415f
C1858 B.n785 VSUBS 0.007415f
C1859 B.n786 VSUBS 0.007415f
C1860 B.n787 VSUBS 0.007415f
C1861 B.n788 VSUBS 0.007415f
C1862 B.n789 VSUBS 0.007415f
C1863 B.n790 VSUBS 0.007415f
C1864 B.n791 VSUBS 0.007415f
C1865 B.n792 VSUBS 0.007415f
C1866 B.n793 VSUBS 0.007415f
C1867 B.n794 VSUBS 0.007415f
C1868 B.n795 VSUBS 0.007415f
C1869 B.n796 VSUBS 0.007415f
C1870 B.n797 VSUBS 0.007415f
C1871 B.n798 VSUBS 0.007415f
C1872 B.n799 VSUBS 0.007415f
C1873 B.n800 VSUBS 0.007415f
C1874 B.n801 VSUBS 0.007415f
C1875 B.n802 VSUBS 0.007415f
C1876 B.n803 VSUBS 0.007415f
C1877 B.n804 VSUBS 0.007415f
C1878 B.n805 VSUBS 0.007415f
C1879 B.n806 VSUBS 0.007415f
C1880 B.n807 VSUBS 0.007415f
C1881 B.n808 VSUBS 0.007415f
C1882 B.n809 VSUBS 0.007415f
C1883 B.n810 VSUBS 0.007415f
C1884 B.n811 VSUBS 0.007415f
C1885 B.n812 VSUBS 0.007415f
C1886 B.n813 VSUBS 0.007415f
C1887 B.n814 VSUBS 0.007415f
C1888 B.n815 VSUBS 0.007415f
C1889 B.n816 VSUBS 0.007415f
C1890 B.n817 VSUBS 0.007415f
C1891 B.n818 VSUBS 0.007415f
C1892 B.n819 VSUBS 0.007415f
C1893 B.n820 VSUBS 0.007415f
C1894 B.n821 VSUBS 0.007415f
C1895 B.n822 VSUBS 0.007415f
C1896 B.n823 VSUBS 0.007415f
C1897 B.n824 VSUBS 0.007415f
C1898 B.n825 VSUBS 0.007415f
C1899 B.n826 VSUBS 0.007415f
C1900 B.n827 VSUBS 0.007415f
C1901 B.n828 VSUBS 0.007415f
C1902 B.n829 VSUBS 0.007415f
C1903 B.n830 VSUBS 0.007415f
C1904 B.n831 VSUBS 0.007415f
C1905 B.n832 VSUBS 0.007415f
C1906 B.n833 VSUBS 0.007415f
C1907 B.n834 VSUBS 0.007415f
C1908 B.n835 VSUBS 0.007415f
C1909 B.n836 VSUBS 0.007415f
C1910 B.n837 VSUBS 0.007415f
C1911 B.n838 VSUBS 0.007415f
C1912 B.n839 VSUBS 0.007415f
C1913 B.n840 VSUBS 0.007415f
C1914 B.n841 VSUBS 0.007415f
C1915 B.n842 VSUBS 0.007415f
C1916 B.n843 VSUBS 0.007415f
C1917 B.n844 VSUBS 0.007415f
C1918 B.n845 VSUBS 0.007415f
C1919 B.n846 VSUBS 0.007415f
C1920 B.n847 VSUBS 0.007415f
C1921 B.n848 VSUBS 0.007415f
C1922 B.n849 VSUBS 0.007415f
C1923 B.n850 VSUBS 0.007415f
C1924 B.n851 VSUBS 0.007415f
C1925 B.n852 VSUBS 0.007415f
C1926 B.n853 VSUBS 0.005125f
C1927 B.n854 VSUBS 0.017179f
C1928 B.n855 VSUBS 0.005997f
C1929 B.n856 VSUBS 0.007415f
C1930 B.n857 VSUBS 0.007415f
C1931 B.n858 VSUBS 0.007415f
C1932 B.n859 VSUBS 0.007415f
C1933 B.n860 VSUBS 0.007415f
C1934 B.n861 VSUBS 0.007415f
C1935 B.n862 VSUBS 0.007415f
C1936 B.n863 VSUBS 0.007415f
C1937 B.n864 VSUBS 0.007415f
C1938 B.n865 VSUBS 0.007415f
C1939 B.n866 VSUBS 0.007415f
C1940 B.n867 VSUBS 0.005997f
C1941 B.n868 VSUBS 0.017179f
C1942 B.n869 VSUBS 0.005125f
C1943 B.n870 VSUBS 0.007415f
C1944 B.n871 VSUBS 0.007415f
C1945 B.n872 VSUBS 0.007415f
C1946 B.n873 VSUBS 0.007415f
C1947 B.n874 VSUBS 0.007415f
C1948 B.n875 VSUBS 0.007415f
C1949 B.n876 VSUBS 0.007415f
C1950 B.n877 VSUBS 0.007415f
C1951 B.n878 VSUBS 0.007415f
C1952 B.n879 VSUBS 0.007415f
C1953 B.n880 VSUBS 0.007415f
C1954 B.n881 VSUBS 0.007415f
C1955 B.n882 VSUBS 0.007415f
C1956 B.n883 VSUBS 0.007415f
C1957 B.n884 VSUBS 0.007415f
C1958 B.n885 VSUBS 0.007415f
C1959 B.n886 VSUBS 0.007415f
C1960 B.n887 VSUBS 0.007415f
C1961 B.n888 VSUBS 0.007415f
C1962 B.n889 VSUBS 0.007415f
C1963 B.n890 VSUBS 0.007415f
C1964 B.n891 VSUBS 0.007415f
C1965 B.n892 VSUBS 0.007415f
C1966 B.n893 VSUBS 0.007415f
C1967 B.n894 VSUBS 0.007415f
C1968 B.n895 VSUBS 0.007415f
C1969 B.n896 VSUBS 0.007415f
C1970 B.n897 VSUBS 0.007415f
C1971 B.n898 VSUBS 0.007415f
C1972 B.n899 VSUBS 0.007415f
C1973 B.n900 VSUBS 0.007415f
C1974 B.n901 VSUBS 0.007415f
C1975 B.n902 VSUBS 0.007415f
C1976 B.n903 VSUBS 0.007415f
C1977 B.n904 VSUBS 0.007415f
C1978 B.n905 VSUBS 0.007415f
C1979 B.n906 VSUBS 0.007415f
C1980 B.n907 VSUBS 0.007415f
C1981 B.n908 VSUBS 0.007415f
C1982 B.n909 VSUBS 0.007415f
C1983 B.n910 VSUBS 0.007415f
C1984 B.n911 VSUBS 0.007415f
C1985 B.n912 VSUBS 0.007415f
C1986 B.n913 VSUBS 0.007415f
C1987 B.n914 VSUBS 0.007415f
C1988 B.n915 VSUBS 0.007415f
C1989 B.n916 VSUBS 0.007415f
C1990 B.n917 VSUBS 0.007415f
C1991 B.n918 VSUBS 0.007415f
C1992 B.n919 VSUBS 0.007415f
C1993 B.n920 VSUBS 0.007415f
C1994 B.n921 VSUBS 0.007415f
C1995 B.n922 VSUBS 0.007415f
C1996 B.n923 VSUBS 0.007415f
C1997 B.n924 VSUBS 0.007415f
C1998 B.n925 VSUBS 0.007415f
C1999 B.n926 VSUBS 0.007415f
C2000 B.n927 VSUBS 0.007415f
C2001 B.n928 VSUBS 0.007415f
C2002 B.n929 VSUBS 0.007415f
C2003 B.n930 VSUBS 0.007415f
C2004 B.n931 VSUBS 0.007415f
C2005 B.n932 VSUBS 0.007415f
C2006 B.n933 VSUBS 0.007415f
C2007 B.n934 VSUBS 0.007415f
C2008 B.n935 VSUBS 0.007415f
C2009 B.n936 VSUBS 0.007415f
C2010 B.n937 VSUBS 0.007415f
C2011 B.n938 VSUBS 0.007415f
C2012 B.n939 VSUBS 0.007415f
C2013 B.n940 VSUBS 0.007415f
C2014 B.n941 VSUBS 0.007415f
C2015 B.n942 VSUBS 0.007415f
C2016 B.n943 VSUBS 0.007415f
C2017 B.n944 VSUBS 0.007415f
C2018 B.n945 VSUBS 0.007415f
C2019 B.n946 VSUBS 0.007415f
C2020 B.n947 VSUBS 0.007415f
C2021 B.n948 VSUBS 0.007415f
C2022 B.n949 VSUBS 0.007415f
C2023 B.n950 VSUBS 0.007415f
C2024 B.n951 VSUBS 0.007415f
C2025 B.n952 VSUBS 0.007415f
C2026 B.n953 VSUBS 0.007415f
C2027 B.n954 VSUBS 0.007415f
C2028 B.n955 VSUBS 0.007415f
C2029 B.n956 VSUBS 0.007415f
C2030 B.n957 VSUBS 0.007415f
C2031 B.n958 VSUBS 0.01725f
C2032 B.n959 VSUBS 0.015898f
C2033 B.n960 VSUBS 0.015898f
C2034 B.n961 VSUBS 0.007415f
C2035 B.n962 VSUBS 0.007415f
C2036 B.n963 VSUBS 0.007415f
C2037 B.n964 VSUBS 0.007415f
C2038 B.n965 VSUBS 0.007415f
C2039 B.n966 VSUBS 0.007415f
C2040 B.n967 VSUBS 0.007415f
C2041 B.n968 VSUBS 0.007415f
C2042 B.n969 VSUBS 0.007415f
C2043 B.n970 VSUBS 0.007415f
C2044 B.n971 VSUBS 0.007415f
C2045 B.n972 VSUBS 0.007415f
C2046 B.n973 VSUBS 0.007415f
C2047 B.n974 VSUBS 0.007415f
C2048 B.n975 VSUBS 0.007415f
C2049 B.n976 VSUBS 0.007415f
C2050 B.n977 VSUBS 0.007415f
C2051 B.n978 VSUBS 0.007415f
C2052 B.n979 VSUBS 0.007415f
C2053 B.n980 VSUBS 0.007415f
C2054 B.n981 VSUBS 0.007415f
C2055 B.n982 VSUBS 0.007415f
C2056 B.n983 VSUBS 0.007415f
C2057 B.n984 VSUBS 0.007415f
C2058 B.n985 VSUBS 0.007415f
C2059 B.n986 VSUBS 0.007415f
C2060 B.n987 VSUBS 0.007415f
C2061 B.n988 VSUBS 0.007415f
C2062 B.n989 VSUBS 0.007415f
C2063 B.n990 VSUBS 0.007415f
C2064 B.n991 VSUBS 0.007415f
C2065 B.n992 VSUBS 0.007415f
C2066 B.n993 VSUBS 0.007415f
C2067 B.n994 VSUBS 0.007415f
C2068 B.n995 VSUBS 0.007415f
C2069 B.n996 VSUBS 0.007415f
C2070 B.n997 VSUBS 0.007415f
C2071 B.n998 VSUBS 0.007415f
C2072 B.n999 VSUBS 0.007415f
C2073 B.n1000 VSUBS 0.007415f
C2074 B.n1001 VSUBS 0.007415f
C2075 B.n1002 VSUBS 0.007415f
C2076 B.n1003 VSUBS 0.007415f
C2077 B.n1004 VSUBS 0.007415f
C2078 B.n1005 VSUBS 0.007415f
C2079 B.n1006 VSUBS 0.007415f
C2080 B.n1007 VSUBS 0.007415f
C2081 B.n1008 VSUBS 0.007415f
C2082 B.n1009 VSUBS 0.007415f
C2083 B.n1010 VSUBS 0.007415f
C2084 B.n1011 VSUBS 0.007415f
C2085 B.n1012 VSUBS 0.007415f
C2086 B.n1013 VSUBS 0.007415f
C2087 B.n1014 VSUBS 0.007415f
C2088 B.n1015 VSUBS 0.007415f
C2089 B.n1016 VSUBS 0.007415f
C2090 B.n1017 VSUBS 0.007415f
C2091 B.n1018 VSUBS 0.007415f
C2092 B.n1019 VSUBS 0.007415f
C2093 B.n1020 VSUBS 0.007415f
C2094 B.n1021 VSUBS 0.007415f
C2095 B.n1022 VSUBS 0.007415f
C2096 B.n1023 VSUBS 0.007415f
C2097 B.n1024 VSUBS 0.007415f
C2098 B.n1025 VSUBS 0.007415f
C2099 B.n1026 VSUBS 0.007415f
C2100 B.n1027 VSUBS 0.007415f
C2101 B.n1028 VSUBS 0.007415f
C2102 B.n1029 VSUBS 0.007415f
C2103 B.n1030 VSUBS 0.007415f
C2104 B.n1031 VSUBS 0.007415f
C2105 B.n1032 VSUBS 0.007415f
C2106 B.n1033 VSUBS 0.007415f
C2107 B.n1034 VSUBS 0.007415f
C2108 B.n1035 VSUBS 0.007415f
C2109 B.n1036 VSUBS 0.007415f
C2110 B.n1037 VSUBS 0.007415f
C2111 B.n1038 VSUBS 0.007415f
C2112 B.n1039 VSUBS 0.007415f
C2113 B.n1040 VSUBS 0.007415f
C2114 B.n1041 VSUBS 0.007415f
C2115 B.n1042 VSUBS 0.007415f
C2116 B.n1043 VSUBS 0.007415f
C2117 B.n1044 VSUBS 0.007415f
C2118 B.n1045 VSUBS 0.007415f
C2119 B.n1046 VSUBS 0.007415f
C2120 B.n1047 VSUBS 0.007415f
C2121 B.n1048 VSUBS 0.007415f
C2122 B.n1049 VSUBS 0.007415f
C2123 B.n1050 VSUBS 0.007415f
C2124 B.n1051 VSUBS 0.007415f
C2125 B.n1052 VSUBS 0.007415f
C2126 B.n1053 VSUBS 0.007415f
C2127 B.n1054 VSUBS 0.007415f
C2128 B.n1055 VSUBS 0.007415f
C2129 B.n1056 VSUBS 0.007415f
C2130 B.n1057 VSUBS 0.007415f
C2131 B.n1058 VSUBS 0.007415f
C2132 B.n1059 VSUBS 0.016789f
.ends

