* NGSPICE file created from diff_pair_sample_1682.ext - technology: sky130A

.subckt diff_pair_sample_1682 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t12 B.t0 sky130_fd_pr__nfet_01v8 ad=2.34465 pd=14.54 as=2.34465 ps=14.54 w=14.21 l=2.97
X1 VDD2.t9 VN.t0 VTAIL.t9 B.t9 sky130_fd_pr__nfet_01v8 ad=2.34465 pd=14.54 as=5.5419 ps=29.2 w=14.21 l=2.97
X2 VTAIL.t3 VN.t1 VDD2.t8 B.t3 sky130_fd_pr__nfet_01v8 ad=2.34465 pd=14.54 as=2.34465 ps=14.54 w=14.21 l=2.97
X3 VTAIL.t19 VP.t1 VDD1.t8 B.t1 sky130_fd_pr__nfet_01v8 ad=2.34465 pd=14.54 as=2.34465 ps=14.54 w=14.21 l=2.97
X4 B.t23 B.t21 B.t22 B.t15 sky130_fd_pr__nfet_01v8 ad=5.5419 pd=29.2 as=0 ps=0 w=14.21 l=2.97
X5 VTAIL.t13 VP.t2 VDD1.t7 B.t5 sky130_fd_pr__nfet_01v8 ad=2.34465 pd=14.54 as=2.34465 ps=14.54 w=14.21 l=2.97
X6 VDD1.t6 VP.t3 VTAIL.t11 B.t8 sky130_fd_pr__nfet_01v8 ad=5.5419 pd=29.2 as=2.34465 ps=14.54 w=14.21 l=2.97
X7 VTAIL.t14 VP.t4 VDD1.t5 B.t6 sky130_fd_pr__nfet_01v8 ad=2.34465 pd=14.54 as=2.34465 ps=14.54 w=14.21 l=2.97
X8 VDD1.t4 VP.t5 VTAIL.t18 B.t9 sky130_fd_pr__nfet_01v8 ad=2.34465 pd=14.54 as=5.5419 ps=29.2 w=14.21 l=2.97
X9 VDD2.t7 VN.t2 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.34465 pd=14.54 as=2.34465 ps=14.54 w=14.21 l=2.97
X10 B.t20 B.t18 B.t19 B.t11 sky130_fd_pr__nfet_01v8 ad=5.5419 pd=29.2 as=0 ps=0 w=14.21 l=2.97
X11 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=5.5419 pd=29.2 as=0 ps=0 w=14.21 l=2.97
X12 VTAIL.t1 VN.t3 VDD2.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=2.34465 pd=14.54 as=2.34465 ps=14.54 w=14.21 l=2.97
X13 VDD2.t5 VN.t4 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=2.34465 pd=14.54 as=5.5419 ps=29.2 w=14.21 l=2.97
X14 VDD2.t4 VN.t5 VTAIL.t8 B.t8 sky130_fd_pr__nfet_01v8 ad=5.5419 pd=29.2 as=2.34465 ps=14.54 w=14.21 l=2.97
X15 VTAIL.t6 VN.t6 VDD2.t3 B.t6 sky130_fd_pr__nfet_01v8 ad=2.34465 pd=14.54 as=2.34465 ps=14.54 w=14.21 l=2.97
X16 VDD2.t2 VN.t7 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=5.5419 pd=29.2 as=2.34465 ps=14.54 w=14.21 l=2.97
X17 VDD1.t3 VP.t6 VTAIL.t10 B.t4 sky130_fd_pr__nfet_01v8 ad=5.5419 pd=29.2 as=2.34465 ps=14.54 w=14.21 l=2.97
X18 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=5.5419 pd=29.2 as=0 ps=0 w=14.21 l=2.97
X19 VTAIL.t15 VP.t7 VDD1.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=2.34465 pd=14.54 as=2.34465 ps=14.54 w=14.21 l=2.97
X20 VDD2.t1 VN.t8 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.34465 pd=14.54 as=2.34465 ps=14.54 w=14.21 l=2.97
X21 VDD1.t1 VP.t8 VTAIL.t17 B.t7 sky130_fd_pr__nfet_01v8 ad=2.34465 pd=14.54 as=5.5419 ps=29.2 w=14.21 l=2.97
X22 VDD1.t0 VP.t9 VTAIL.t16 B.t2 sky130_fd_pr__nfet_01v8 ad=2.34465 pd=14.54 as=2.34465 ps=14.54 w=14.21 l=2.97
X23 VTAIL.t5 VN.t9 VDD2.t0 B.t5 sky130_fd_pr__nfet_01v8 ad=2.34465 pd=14.54 as=2.34465 ps=14.54 w=14.21 l=2.97
R0 VP.n27 VP.n24 161.3
R1 VP.n29 VP.n28 161.3
R2 VP.n30 VP.n23 161.3
R3 VP.n32 VP.n31 161.3
R4 VP.n33 VP.n22 161.3
R5 VP.n35 VP.n34 161.3
R6 VP.n36 VP.n21 161.3
R7 VP.n39 VP.n38 161.3
R8 VP.n40 VP.n20 161.3
R9 VP.n42 VP.n41 161.3
R10 VP.n43 VP.n19 161.3
R11 VP.n45 VP.n44 161.3
R12 VP.n46 VP.n18 161.3
R13 VP.n48 VP.n47 161.3
R14 VP.n50 VP.n17 161.3
R15 VP.n52 VP.n51 161.3
R16 VP.n53 VP.n16 161.3
R17 VP.n55 VP.n54 161.3
R18 VP.n56 VP.n15 161.3
R19 VP.n58 VP.n57 161.3
R20 VP.n103 VP.n102 161.3
R21 VP.n101 VP.n1 161.3
R22 VP.n100 VP.n99 161.3
R23 VP.n98 VP.n2 161.3
R24 VP.n97 VP.n96 161.3
R25 VP.n95 VP.n3 161.3
R26 VP.n93 VP.n92 161.3
R27 VP.n91 VP.n4 161.3
R28 VP.n90 VP.n89 161.3
R29 VP.n88 VP.n5 161.3
R30 VP.n87 VP.n86 161.3
R31 VP.n85 VP.n6 161.3
R32 VP.n84 VP.n83 161.3
R33 VP.n81 VP.n7 161.3
R34 VP.n80 VP.n79 161.3
R35 VP.n78 VP.n8 161.3
R36 VP.n77 VP.n76 161.3
R37 VP.n75 VP.n9 161.3
R38 VP.n74 VP.n73 161.3
R39 VP.n72 VP.n10 161.3
R40 VP.n71 VP.n70 161.3
R41 VP.n68 VP.n11 161.3
R42 VP.n67 VP.n66 161.3
R43 VP.n65 VP.n12 161.3
R44 VP.n64 VP.n63 161.3
R45 VP.n62 VP.n13 161.3
R46 VP.n26 VP.t6 146.827
R47 VP.n61 VP.t3 115.308
R48 VP.n69 VP.t2 115.308
R49 VP.n82 VP.t0 115.308
R50 VP.n94 VP.t1 115.308
R51 VP.n0 VP.t8 115.308
R52 VP.n14 VP.t5 115.308
R53 VP.n49 VP.t7 115.308
R54 VP.n37 VP.t9 115.308
R55 VP.n25 VP.t4 115.308
R56 VP.n61 VP.n60 72.9405
R57 VP.n104 VP.n0 72.9405
R58 VP.n59 VP.n14 72.9405
R59 VP.n26 VP.n25 71.0033
R60 VP.n60 VP.n59 56.8705
R61 VP.n67 VP.n12 56.5193
R62 VP.n100 VP.n2 56.5193
R63 VP.n55 VP.n16 56.5193
R64 VP.n76 VP.n8 50.2061
R65 VP.n88 VP.n87 50.2061
R66 VP.n43 VP.n42 50.2061
R67 VP.n31 VP.n22 50.2061
R68 VP.n76 VP.n75 30.7807
R69 VP.n89 VP.n88 30.7807
R70 VP.n44 VP.n43 30.7807
R71 VP.n31 VP.n30 30.7807
R72 VP.n63 VP.n62 24.4675
R73 VP.n63 VP.n12 24.4675
R74 VP.n68 VP.n67 24.4675
R75 VP.n70 VP.n68 24.4675
R76 VP.n74 VP.n10 24.4675
R77 VP.n75 VP.n74 24.4675
R78 VP.n80 VP.n8 24.4675
R79 VP.n81 VP.n80 24.4675
R80 VP.n83 VP.n6 24.4675
R81 VP.n87 VP.n6 24.4675
R82 VP.n89 VP.n4 24.4675
R83 VP.n93 VP.n4 24.4675
R84 VP.n96 VP.n95 24.4675
R85 VP.n96 VP.n2 24.4675
R86 VP.n101 VP.n100 24.4675
R87 VP.n102 VP.n101 24.4675
R88 VP.n56 VP.n55 24.4675
R89 VP.n57 VP.n56 24.4675
R90 VP.n44 VP.n18 24.4675
R91 VP.n48 VP.n18 24.4675
R92 VP.n51 VP.n50 24.4675
R93 VP.n51 VP.n16 24.4675
R94 VP.n35 VP.n22 24.4675
R95 VP.n36 VP.n35 24.4675
R96 VP.n38 VP.n20 24.4675
R97 VP.n42 VP.n20 24.4675
R98 VP.n29 VP.n24 24.4675
R99 VP.n30 VP.n29 24.4675
R100 VP.n70 VP.n69 22.0208
R101 VP.n95 VP.n94 22.0208
R102 VP.n50 VP.n49 22.0208
R103 VP.n62 VP.n61 17.1274
R104 VP.n102 VP.n0 17.1274
R105 VP.n57 VP.n14 17.1274
R106 VP.n82 VP.n81 12.234
R107 VP.n83 VP.n82 12.234
R108 VP.n37 VP.n36 12.234
R109 VP.n38 VP.n37 12.234
R110 VP.n27 VP.n26 5.75991
R111 VP.n69 VP.n10 2.4472
R112 VP.n94 VP.n93 2.4472
R113 VP.n49 VP.n48 2.4472
R114 VP.n25 VP.n24 2.4472
R115 VP.n59 VP.n58 0.354971
R116 VP.n60 VP.n13 0.354971
R117 VP.n104 VP.n103 0.354971
R118 VP VP.n104 0.26696
R119 VP.n28 VP.n27 0.189894
R120 VP.n28 VP.n23 0.189894
R121 VP.n32 VP.n23 0.189894
R122 VP.n33 VP.n32 0.189894
R123 VP.n34 VP.n33 0.189894
R124 VP.n34 VP.n21 0.189894
R125 VP.n39 VP.n21 0.189894
R126 VP.n40 VP.n39 0.189894
R127 VP.n41 VP.n40 0.189894
R128 VP.n41 VP.n19 0.189894
R129 VP.n45 VP.n19 0.189894
R130 VP.n46 VP.n45 0.189894
R131 VP.n47 VP.n46 0.189894
R132 VP.n47 VP.n17 0.189894
R133 VP.n52 VP.n17 0.189894
R134 VP.n53 VP.n52 0.189894
R135 VP.n54 VP.n53 0.189894
R136 VP.n54 VP.n15 0.189894
R137 VP.n58 VP.n15 0.189894
R138 VP.n64 VP.n13 0.189894
R139 VP.n65 VP.n64 0.189894
R140 VP.n66 VP.n65 0.189894
R141 VP.n66 VP.n11 0.189894
R142 VP.n71 VP.n11 0.189894
R143 VP.n72 VP.n71 0.189894
R144 VP.n73 VP.n72 0.189894
R145 VP.n73 VP.n9 0.189894
R146 VP.n77 VP.n9 0.189894
R147 VP.n78 VP.n77 0.189894
R148 VP.n79 VP.n78 0.189894
R149 VP.n79 VP.n7 0.189894
R150 VP.n84 VP.n7 0.189894
R151 VP.n85 VP.n84 0.189894
R152 VP.n86 VP.n85 0.189894
R153 VP.n86 VP.n5 0.189894
R154 VP.n90 VP.n5 0.189894
R155 VP.n91 VP.n90 0.189894
R156 VP.n92 VP.n91 0.189894
R157 VP.n92 VP.n3 0.189894
R158 VP.n97 VP.n3 0.189894
R159 VP.n98 VP.n97 0.189894
R160 VP.n99 VP.n98 0.189894
R161 VP.n99 VP.n1 0.189894
R162 VP.n103 VP.n1 0.189894
R163 VTAIL.n320 VTAIL.n248 289.615
R164 VTAIL.n74 VTAIL.n2 289.615
R165 VTAIL.n242 VTAIL.n170 289.615
R166 VTAIL.n160 VTAIL.n88 289.615
R167 VTAIL.n272 VTAIL.n271 185
R168 VTAIL.n277 VTAIL.n276 185
R169 VTAIL.n279 VTAIL.n278 185
R170 VTAIL.n268 VTAIL.n267 185
R171 VTAIL.n285 VTAIL.n284 185
R172 VTAIL.n287 VTAIL.n286 185
R173 VTAIL.n264 VTAIL.n263 185
R174 VTAIL.n294 VTAIL.n293 185
R175 VTAIL.n295 VTAIL.n262 185
R176 VTAIL.n297 VTAIL.n296 185
R177 VTAIL.n260 VTAIL.n259 185
R178 VTAIL.n303 VTAIL.n302 185
R179 VTAIL.n305 VTAIL.n304 185
R180 VTAIL.n256 VTAIL.n255 185
R181 VTAIL.n311 VTAIL.n310 185
R182 VTAIL.n313 VTAIL.n312 185
R183 VTAIL.n252 VTAIL.n251 185
R184 VTAIL.n319 VTAIL.n318 185
R185 VTAIL.n321 VTAIL.n320 185
R186 VTAIL.n26 VTAIL.n25 185
R187 VTAIL.n31 VTAIL.n30 185
R188 VTAIL.n33 VTAIL.n32 185
R189 VTAIL.n22 VTAIL.n21 185
R190 VTAIL.n39 VTAIL.n38 185
R191 VTAIL.n41 VTAIL.n40 185
R192 VTAIL.n18 VTAIL.n17 185
R193 VTAIL.n48 VTAIL.n47 185
R194 VTAIL.n49 VTAIL.n16 185
R195 VTAIL.n51 VTAIL.n50 185
R196 VTAIL.n14 VTAIL.n13 185
R197 VTAIL.n57 VTAIL.n56 185
R198 VTAIL.n59 VTAIL.n58 185
R199 VTAIL.n10 VTAIL.n9 185
R200 VTAIL.n65 VTAIL.n64 185
R201 VTAIL.n67 VTAIL.n66 185
R202 VTAIL.n6 VTAIL.n5 185
R203 VTAIL.n73 VTAIL.n72 185
R204 VTAIL.n75 VTAIL.n74 185
R205 VTAIL.n243 VTAIL.n242 185
R206 VTAIL.n241 VTAIL.n240 185
R207 VTAIL.n174 VTAIL.n173 185
R208 VTAIL.n235 VTAIL.n234 185
R209 VTAIL.n233 VTAIL.n232 185
R210 VTAIL.n178 VTAIL.n177 185
R211 VTAIL.n227 VTAIL.n226 185
R212 VTAIL.n225 VTAIL.n224 185
R213 VTAIL.n182 VTAIL.n181 185
R214 VTAIL.n219 VTAIL.n218 185
R215 VTAIL.n217 VTAIL.n184 185
R216 VTAIL.n216 VTAIL.n215 185
R217 VTAIL.n187 VTAIL.n185 185
R218 VTAIL.n210 VTAIL.n209 185
R219 VTAIL.n208 VTAIL.n207 185
R220 VTAIL.n191 VTAIL.n190 185
R221 VTAIL.n202 VTAIL.n201 185
R222 VTAIL.n200 VTAIL.n199 185
R223 VTAIL.n195 VTAIL.n194 185
R224 VTAIL.n161 VTAIL.n160 185
R225 VTAIL.n159 VTAIL.n158 185
R226 VTAIL.n92 VTAIL.n91 185
R227 VTAIL.n153 VTAIL.n152 185
R228 VTAIL.n151 VTAIL.n150 185
R229 VTAIL.n96 VTAIL.n95 185
R230 VTAIL.n145 VTAIL.n144 185
R231 VTAIL.n143 VTAIL.n142 185
R232 VTAIL.n100 VTAIL.n99 185
R233 VTAIL.n137 VTAIL.n136 185
R234 VTAIL.n135 VTAIL.n102 185
R235 VTAIL.n134 VTAIL.n133 185
R236 VTAIL.n105 VTAIL.n103 185
R237 VTAIL.n128 VTAIL.n127 185
R238 VTAIL.n126 VTAIL.n125 185
R239 VTAIL.n109 VTAIL.n108 185
R240 VTAIL.n120 VTAIL.n119 185
R241 VTAIL.n118 VTAIL.n117 185
R242 VTAIL.n113 VTAIL.n112 185
R243 VTAIL.n273 VTAIL.t9 149.524
R244 VTAIL.n27 VTAIL.t17 149.524
R245 VTAIL.n196 VTAIL.t18 149.524
R246 VTAIL.n114 VTAIL.t7 149.524
R247 VTAIL.n277 VTAIL.n271 104.615
R248 VTAIL.n278 VTAIL.n277 104.615
R249 VTAIL.n278 VTAIL.n267 104.615
R250 VTAIL.n285 VTAIL.n267 104.615
R251 VTAIL.n286 VTAIL.n285 104.615
R252 VTAIL.n286 VTAIL.n263 104.615
R253 VTAIL.n294 VTAIL.n263 104.615
R254 VTAIL.n295 VTAIL.n294 104.615
R255 VTAIL.n296 VTAIL.n295 104.615
R256 VTAIL.n296 VTAIL.n259 104.615
R257 VTAIL.n303 VTAIL.n259 104.615
R258 VTAIL.n304 VTAIL.n303 104.615
R259 VTAIL.n304 VTAIL.n255 104.615
R260 VTAIL.n311 VTAIL.n255 104.615
R261 VTAIL.n312 VTAIL.n311 104.615
R262 VTAIL.n312 VTAIL.n251 104.615
R263 VTAIL.n319 VTAIL.n251 104.615
R264 VTAIL.n320 VTAIL.n319 104.615
R265 VTAIL.n31 VTAIL.n25 104.615
R266 VTAIL.n32 VTAIL.n31 104.615
R267 VTAIL.n32 VTAIL.n21 104.615
R268 VTAIL.n39 VTAIL.n21 104.615
R269 VTAIL.n40 VTAIL.n39 104.615
R270 VTAIL.n40 VTAIL.n17 104.615
R271 VTAIL.n48 VTAIL.n17 104.615
R272 VTAIL.n49 VTAIL.n48 104.615
R273 VTAIL.n50 VTAIL.n49 104.615
R274 VTAIL.n50 VTAIL.n13 104.615
R275 VTAIL.n57 VTAIL.n13 104.615
R276 VTAIL.n58 VTAIL.n57 104.615
R277 VTAIL.n58 VTAIL.n9 104.615
R278 VTAIL.n65 VTAIL.n9 104.615
R279 VTAIL.n66 VTAIL.n65 104.615
R280 VTAIL.n66 VTAIL.n5 104.615
R281 VTAIL.n73 VTAIL.n5 104.615
R282 VTAIL.n74 VTAIL.n73 104.615
R283 VTAIL.n242 VTAIL.n241 104.615
R284 VTAIL.n241 VTAIL.n173 104.615
R285 VTAIL.n234 VTAIL.n173 104.615
R286 VTAIL.n234 VTAIL.n233 104.615
R287 VTAIL.n233 VTAIL.n177 104.615
R288 VTAIL.n226 VTAIL.n177 104.615
R289 VTAIL.n226 VTAIL.n225 104.615
R290 VTAIL.n225 VTAIL.n181 104.615
R291 VTAIL.n218 VTAIL.n181 104.615
R292 VTAIL.n218 VTAIL.n217 104.615
R293 VTAIL.n217 VTAIL.n216 104.615
R294 VTAIL.n216 VTAIL.n185 104.615
R295 VTAIL.n209 VTAIL.n185 104.615
R296 VTAIL.n209 VTAIL.n208 104.615
R297 VTAIL.n208 VTAIL.n190 104.615
R298 VTAIL.n201 VTAIL.n190 104.615
R299 VTAIL.n201 VTAIL.n200 104.615
R300 VTAIL.n200 VTAIL.n194 104.615
R301 VTAIL.n160 VTAIL.n159 104.615
R302 VTAIL.n159 VTAIL.n91 104.615
R303 VTAIL.n152 VTAIL.n91 104.615
R304 VTAIL.n152 VTAIL.n151 104.615
R305 VTAIL.n151 VTAIL.n95 104.615
R306 VTAIL.n144 VTAIL.n95 104.615
R307 VTAIL.n144 VTAIL.n143 104.615
R308 VTAIL.n143 VTAIL.n99 104.615
R309 VTAIL.n136 VTAIL.n99 104.615
R310 VTAIL.n136 VTAIL.n135 104.615
R311 VTAIL.n135 VTAIL.n134 104.615
R312 VTAIL.n134 VTAIL.n103 104.615
R313 VTAIL.n127 VTAIL.n103 104.615
R314 VTAIL.n127 VTAIL.n126 104.615
R315 VTAIL.n126 VTAIL.n108 104.615
R316 VTAIL.n119 VTAIL.n108 104.615
R317 VTAIL.n119 VTAIL.n118 104.615
R318 VTAIL.n118 VTAIL.n112 104.615
R319 VTAIL.t9 VTAIL.n271 52.3082
R320 VTAIL.t17 VTAIL.n25 52.3082
R321 VTAIL.t18 VTAIL.n194 52.3082
R322 VTAIL.t7 VTAIL.n112 52.3082
R323 VTAIL.n327 VTAIL.n326 43.3918
R324 VTAIL.n1 VTAIL.n0 43.3918
R325 VTAIL.n81 VTAIL.n80 43.3918
R326 VTAIL.n83 VTAIL.n82 43.3918
R327 VTAIL.n169 VTAIL.n168 43.3918
R328 VTAIL.n167 VTAIL.n166 43.3918
R329 VTAIL.n87 VTAIL.n86 43.3918
R330 VTAIL.n85 VTAIL.n84 43.3918
R331 VTAIL.n325 VTAIL.n324 30.8278
R332 VTAIL.n79 VTAIL.n78 30.8278
R333 VTAIL.n247 VTAIL.n246 30.8278
R334 VTAIL.n165 VTAIL.n164 30.8278
R335 VTAIL.n85 VTAIL.n83 30.3065
R336 VTAIL.n325 VTAIL.n247 27.4617
R337 VTAIL.n297 VTAIL.n262 13.1884
R338 VTAIL.n51 VTAIL.n16 13.1884
R339 VTAIL.n219 VTAIL.n184 13.1884
R340 VTAIL.n137 VTAIL.n102 13.1884
R341 VTAIL.n293 VTAIL.n292 12.8005
R342 VTAIL.n298 VTAIL.n260 12.8005
R343 VTAIL.n47 VTAIL.n46 12.8005
R344 VTAIL.n52 VTAIL.n14 12.8005
R345 VTAIL.n220 VTAIL.n182 12.8005
R346 VTAIL.n215 VTAIL.n186 12.8005
R347 VTAIL.n138 VTAIL.n100 12.8005
R348 VTAIL.n133 VTAIL.n104 12.8005
R349 VTAIL.n291 VTAIL.n264 12.0247
R350 VTAIL.n302 VTAIL.n301 12.0247
R351 VTAIL.n45 VTAIL.n18 12.0247
R352 VTAIL.n56 VTAIL.n55 12.0247
R353 VTAIL.n224 VTAIL.n223 12.0247
R354 VTAIL.n214 VTAIL.n187 12.0247
R355 VTAIL.n142 VTAIL.n141 12.0247
R356 VTAIL.n132 VTAIL.n105 12.0247
R357 VTAIL.n288 VTAIL.n287 11.249
R358 VTAIL.n305 VTAIL.n258 11.249
R359 VTAIL.n42 VTAIL.n41 11.249
R360 VTAIL.n59 VTAIL.n12 11.249
R361 VTAIL.n227 VTAIL.n180 11.249
R362 VTAIL.n211 VTAIL.n210 11.249
R363 VTAIL.n145 VTAIL.n98 11.249
R364 VTAIL.n129 VTAIL.n128 11.249
R365 VTAIL.n284 VTAIL.n266 10.4732
R366 VTAIL.n306 VTAIL.n256 10.4732
R367 VTAIL.n38 VTAIL.n20 10.4732
R368 VTAIL.n60 VTAIL.n10 10.4732
R369 VTAIL.n228 VTAIL.n178 10.4732
R370 VTAIL.n207 VTAIL.n189 10.4732
R371 VTAIL.n146 VTAIL.n96 10.4732
R372 VTAIL.n125 VTAIL.n107 10.4732
R373 VTAIL.n273 VTAIL.n272 10.2747
R374 VTAIL.n27 VTAIL.n26 10.2747
R375 VTAIL.n196 VTAIL.n195 10.2747
R376 VTAIL.n114 VTAIL.n113 10.2747
R377 VTAIL.n283 VTAIL.n268 9.69747
R378 VTAIL.n310 VTAIL.n309 9.69747
R379 VTAIL.n37 VTAIL.n22 9.69747
R380 VTAIL.n64 VTAIL.n63 9.69747
R381 VTAIL.n232 VTAIL.n231 9.69747
R382 VTAIL.n206 VTAIL.n191 9.69747
R383 VTAIL.n150 VTAIL.n149 9.69747
R384 VTAIL.n124 VTAIL.n109 9.69747
R385 VTAIL.n324 VTAIL.n323 9.45567
R386 VTAIL.n78 VTAIL.n77 9.45567
R387 VTAIL.n246 VTAIL.n245 9.45567
R388 VTAIL.n164 VTAIL.n163 9.45567
R389 VTAIL.n250 VTAIL.n249 9.3005
R390 VTAIL.n323 VTAIL.n322 9.3005
R391 VTAIL.n315 VTAIL.n314 9.3005
R392 VTAIL.n254 VTAIL.n253 9.3005
R393 VTAIL.n309 VTAIL.n308 9.3005
R394 VTAIL.n307 VTAIL.n306 9.3005
R395 VTAIL.n258 VTAIL.n257 9.3005
R396 VTAIL.n301 VTAIL.n300 9.3005
R397 VTAIL.n299 VTAIL.n298 9.3005
R398 VTAIL.n275 VTAIL.n274 9.3005
R399 VTAIL.n270 VTAIL.n269 9.3005
R400 VTAIL.n281 VTAIL.n280 9.3005
R401 VTAIL.n283 VTAIL.n282 9.3005
R402 VTAIL.n266 VTAIL.n265 9.3005
R403 VTAIL.n289 VTAIL.n288 9.3005
R404 VTAIL.n291 VTAIL.n290 9.3005
R405 VTAIL.n292 VTAIL.n261 9.3005
R406 VTAIL.n317 VTAIL.n316 9.3005
R407 VTAIL.n4 VTAIL.n3 9.3005
R408 VTAIL.n77 VTAIL.n76 9.3005
R409 VTAIL.n69 VTAIL.n68 9.3005
R410 VTAIL.n8 VTAIL.n7 9.3005
R411 VTAIL.n63 VTAIL.n62 9.3005
R412 VTAIL.n61 VTAIL.n60 9.3005
R413 VTAIL.n12 VTAIL.n11 9.3005
R414 VTAIL.n55 VTAIL.n54 9.3005
R415 VTAIL.n53 VTAIL.n52 9.3005
R416 VTAIL.n29 VTAIL.n28 9.3005
R417 VTAIL.n24 VTAIL.n23 9.3005
R418 VTAIL.n35 VTAIL.n34 9.3005
R419 VTAIL.n37 VTAIL.n36 9.3005
R420 VTAIL.n20 VTAIL.n19 9.3005
R421 VTAIL.n43 VTAIL.n42 9.3005
R422 VTAIL.n45 VTAIL.n44 9.3005
R423 VTAIL.n46 VTAIL.n15 9.3005
R424 VTAIL.n71 VTAIL.n70 9.3005
R425 VTAIL.n172 VTAIL.n171 9.3005
R426 VTAIL.n239 VTAIL.n238 9.3005
R427 VTAIL.n237 VTAIL.n236 9.3005
R428 VTAIL.n176 VTAIL.n175 9.3005
R429 VTAIL.n231 VTAIL.n230 9.3005
R430 VTAIL.n229 VTAIL.n228 9.3005
R431 VTAIL.n180 VTAIL.n179 9.3005
R432 VTAIL.n223 VTAIL.n222 9.3005
R433 VTAIL.n221 VTAIL.n220 9.3005
R434 VTAIL.n186 VTAIL.n183 9.3005
R435 VTAIL.n214 VTAIL.n213 9.3005
R436 VTAIL.n212 VTAIL.n211 9.3005
R437 VTAIL.n189 VTAIL.n188 9.3005
R438 VTAIL.n206 VTAIL.n205 9.3005
R439 VTAIL.n204 VTAIL.n203 9.3005
R440 VTAIL.n193 VTAIL.n192 9.3005
R441 VTAIL.n198 VTAIL.n197 9.3005
R442 VTAIL.n245 VTAIL.n244 9.3005
R443 VTAIL.n116 VTAIL.n115 9.3005
R444 VTAIL.n111 VTAIL.n110 9.3005
R445 VTAIL.n122 VTAIL.n121 9.3005
R446 VTAIL.n124 VTAIL.n123 9.3005
R447 VTAIL.n107 VTAIL.n106 9.3005
R448 VTAIL.n130 VTAIL.n129 9.3005
R449 VTAIL.n132 VTAIL.n131 9.3005
R450 VTAIL.n104 VTAIL.n101 9.3005
R451 VTAIL.n163 VTAIL.n162 9.3005
R452 VTAIL.n90 VTAIL.n89 9.3005
R453 VTAIL.n157 VTAIL.n156 9.3005
R454 VTAIL.n155 VTAIL.n154 9.3005
R455 VTAIL.n94 VTAIL.n93 9.3005
R456 VTAIL.n149 VTAIL.n148 9.3005
R457 VTAIL.n147 VTAIL.n146 9.3005
R458 VTAIL.n98 VTAIL.n97 9.3005
R459 VTAIL.n141 VTAIL.n140 9.3005
R460 VTAIL.n139 VTAIL.n138 9.3005
R461 VTAIL.n280 VTAIL.n279 8.92171
R462 VTAIL.n313 VTAIL.n254 8.92171
R463 VTAIL.n34 VTAIL.n33 8.92171
R464 VTAIL.n67 VTAIL.n8 8.92171
R465 VTAIL.n235 VTAIL.n176 8.92171
R466 VTAIL.n203 VTAIL.n202 8.92171
R467 VTAIL.n153 VTAIL.n94 8.92171
R468 VTAIL.n121 VTAIL.n120 8.92171
R469 VTAIL.n276 VTAIL.n270 8.14595
R470 VTAIL.n314 VTAIL.n252 8.14595
R471 VTAIL.n324 VTAIL.n248 8.14595
R472 VTAIL.n30 VTAIL.n24 8.14595
R473 VTAIL.n68 VTAIL.n6 8.14595
R474 VTAIL.n78 VTAIL.n2 8.14595
R475 VTAIL.n246 VTAIL.n170 8.14595
R476 VTAIL.n236 VTAIL.n174 8.14595
R477 VTAIL.n199 VTAIL.n193 8.14595
R478 VTAIL.n164 VTAIL.n88 8.14595
R479 VTAIL.n154 VTAIL.n92 8.14595
R480 VTAIL.n117 VTAIL.n111 8.14595
R481 VTAIL.n275 VTAIL.n272 7.3702
R482 VTAIL.n318 VTAIL.n317 7.3702
R483 VTAIL.n322 VTAIL.n321 7.3702
R484 VTAIL.n29 VTAIL.n26 7.3702
R485 VTAIL.n72 VTAIL.n71 7.3702
R486 VTAIL.n76 VTAIL.n75 7.3702
R487 VTAIL.n244 VTAIL.n243 7.3702
R488 VTAIL.n240 VTAIL.n239 7.3702
R489 VTAIL.n198 VTAIL.n195 7.3702
R490 VTAIL.n162 VTAIL.n161 7.3702
R491 VTAIL.n158 VTAIL.n157 7.3702
R492 VTAIL.n116 VTAIL.n113 7.3702
R493 VTAIL.n318 VTAIL.n250 6.59444
R494 VTAIL.n321 VTAIL.n250 6.59444
R495 VTAIL.n72 VTAIL.n4 6.59444
R496 VTAIL.n75 VTAIL.n4 6.59444
R497 VTAIL.n243 VTAIL.n172 6.59444
R498 VTAIL.n240 VTAIL.n172 6.59444
R499 VTAIL.n161 VTAIL.n90 6.59444
R500 VTAIL.n158 VTAIL.n90 6.59444
R501 VTAIL.n276 VTAIL.n275 5.81868
R502 VTAIL.n317 VTAIL.n252 5.81868
R503 VTAIL.n322 VTAIL.n248 5.81868
R504 VTAIL.n30 VTAIL.n29 5.81868
R505 VTAIL.n71 VTAIL.n6 5.81868
R506 VTAIL.n76 VTAIL.n2 5.81868
R507 VTAIL.n244 VTAIL.n170 5.81868
R508 VTAIL.n239 VTAIL.n174 5.81868
R509 VTAIL.n199 VTAIL.n198 5.81868
R510 VTAIL.n162 VTAIL.n88 5.81868
R511 VTAIL.n157 VTAIL.n92 5.81868
R512 VTAIL.n117 VTAIL.n116 5.81868
R513 VTAIL.n279 VTAIL.n270 5.04292
R514 VTAIL.n314 VTAIL.n313 5.04292
R515 VTAIL.n33 VTAIL.n24 5.04292
R516 VTAIL.n68 VTAIL.n67 5.04292
R517 VTAIL.n236 VTAIL.n235 5.04292
R518 VTAIL.n202 VTAIL.n193 5.04292
R519 VTAIL.n154 VTAIL.n153 5.04292
R520 VTAIL.n120 VTAIL.n111 5.04292
R521 VTAIL.n280 VTAIL.n268 4.26717
R522 VTAIL.n310 VTAIL.n254 4.26717
R523 VTAIL.n34 VTAIL.n22 4.26717
R524 VTAIL.n64 VTAIL.n8 4.26717
R525 VTAIL.n232 VTAIL.n176 4.26717
R526 VTAIL.n203 VTAIL.n191 4.26717
R527 VTAIL.n150 VTAIL.n94 4.26717
R528 VTAIL.n121 VTAIL.n109 4.26717
R529 VTAIL.n284 VTAIL.n283 3.49141
R530 VTAIL.n309 VTAIL.n256 3.49141
R531 VTAIL.n38 VTAIL.n37 3.49141
R532 VTAIL.n63 VTAIL.n10 3.49141
R533 VTAIL.n231 VTAIL.n178 3.49141
R534 VTAIL.n207 VTAIL.n206 3.49141
R535 VTAIL.n149 VTAIL.n96 3.49141
R536 VTAIL.n125 VTAIL.n124 3.49141
R537 VTAIL.n87 VTAIL.n85 2.84533
R538 VTAIL.n165 VTAIL.n87 2.84533
R539 VTAIL.n169 VTAIL.n167 2.84533
R540 VTAIL.n247 VTAIL.n169 2.84533
R541 VTAIL.n83 VTAIL.n81 2.84533
R542 VTAIL.n81 VTAIL.n79 2.84533
R543 VTAIL.n327 VTAIL.n325 2.84533
R544 VTAIL.n274 VTAIL.n273 2.84303
R545 VTAIL.n28 VTAIL.n27 2.84303
R546 VTAIL.n115 VTAIL.n114 2.84303
R547 VTAIL.n197 VTAIL.n196 2.84303
R548 VTAIL.n287 VTAIL.n266 2.71565
R549 VTAIL.n306 VTAIL.n305 2.71565
R550 VTAIL.n41 VTAIL.n20 2.71565
R551 VTAIL.n60 VTAIL.n59 2.71565
R552 VTAIL.n228 VTAIL.n227 2.71565
R553 VTAIL.n210 VTAIL.n189 2.71565
R554 VTAIL.n146 VTAIL.n145 2.71565
R555 VTAIL.n128 VTAIL.n107 2.71565
R556 VTAIL VTAIL.n1 2.19231
R557 VTAIL.n288 VTAIL.n264 1.93989
R558 VTAIL.n302 VTAIL.n258 1.93989
R559 VTAIL.n42 VTAIL.n18 1.93989
R560 VTAIL.n56 VTAIL.n12 1.93989
R561 VTAIL.n224 VTAIL.n180 1.93989
R562 VTAIL.n211 VTAIL.n187 1.93989
R563 VTAIL.n142 VTAIL.n98 1.93989
R564 VTAIL.n129 VTAIL.n105 1.93989
R565 VTAIL.n167 VTAIL.n165 1.89274
R566 VTAIL.n79 VTAIL.n1 1.89274
R567 VTAIL.n326 VTAIL.t2 1.39388
R568 VTAIL.n326 VTAIL.t3 1.39388
R569 VTAIL.n0 VTAIL.t4 1.39388
R570 VTAIL.n0 VTAIL.t6 1.39388
R571 VTAIL.n80 VTAIL.t12 1.39388
R572 VTAIL.n80 VTAIL.t19 1.39388
R573 VTAIL.n82 VTAIL.t11 1.39388
R574 VTAIL.n82 VTAIL.t13 1.39388
R575 VTAIL.n168 VTAIL.t16 1.39388
R576 VTAIL.n168 VTAIL.t15 1.39388
R577 VTAIL.n166 VTAIL.t10 1.39388
R578 VTAIL.n166 VTAIL.t14 1.39388
R579 VTAIL.n86 VTAIL.t0 1.39388
R580 VTAIL.n86 VTAIL.t1 1.39388
R581 VTAIL.n84 VTAIL.t8 1.39388
R582 VTAIL.n84 VTAIL.t5 1.39388
R583 VTAIL.n293 VTAIL.n291 1.16414
R584 VTAIL.n301 VTAIL.n260 1.16414
R585 VTAIL.n47 VTAIL.n45 1.16414
R586 VTAIL.n55 VTAIL.n14 1.16414
R587 VTAIL.n223 VTAIL.n182 1.16414
R588 VTAIL.n215 VTAIL.n214 1.16414
R589 VTAIL.n141 VTAIL.n100 1.16414
R590 VTAIL.n133 VTAIL.n132 1.16414
R591 VTAIL VTAIL.n327 0.653517
R592 VTAIL.n292 VTAIL.n262 0.388379
R593 VTAIL.n298 VTAIL.n297 0.388379
R594 VTAIL.n46 VTAIL.n16 0.388379
R595 VTAIL.n52 VTAIL.n51 0.388379
R596 VTAIL.n220 VTAIL.n219 0.388379
R597 VTAIL.n186 VTAIL.n184 0.388379
R598 VTAIL.n138 VTAIL.n137 0.388379
R599 VTAIL.n104 VTAIL.n102 0.388379
R600 VTAIL.n274 VTAIL.n269 0.155672
R601 VTAIL.n281 VTAIL.n269 0.155672
R602 VTAIL.n282 VTAIL.n281 0.155672
R603 VTAIL.n282 VTAIL.n265 0.155672
R604 VTAIL.n289 VTAIL.n265 0.155672
R605 VTAIL.n290 VTAIL.n289 0.155672
R606 VTAIL.n290 VTAIL.n261 0.155672
R607 VTAIL.n299 VTAIL.n261 0.155672
R608 VTAIL.n300 VTAIL.n299 0.155672
R609 VTAIL.n300 VTAIL.n257 0.155672
R610 VTAIL.n307 VTAIL.n257 0.155672
R611 VTAIL.n308 VTAIL.n307 0.155672
R612 VTAIL.n308 VTAIL.n253 0.155672
R613 VTAIL.n315 VTAIL.n253 0.155672
R614 VTAIL.n316 VTAIL.n315 0.155672
R615 VTAIL.n316 VTAIL.n249 0.155672
R616 VTAIL.n323 VTAIL.n249 0.155672
R617 VTAIL.n28 VTAIL.n23 0.155672
R618 VTAIL.n35 VTAIL.n23 0.155672
R619 VTAIL.n36 VTAIL.n35 0.155672
R620 VTAIL.n36 VTAIL.n19 0.155672
R621 VTAIL.n43 VTAIL.n19 0.155672
R622 VTAIL.n44 VTAIL.n43 0.155672
R623 VTAIL.n44 VTAIL.n15 0.155672
R624 VTAIL.n53 VTAIL.n15 0.155672
R625 VTAIL.n54 VTAIL.n53 0.155672
R626 VTAIL.n54 VTAIL.n11 0.155672
R627 VTAIL.n61 VTAIL.n11 0.155672
R628 VTAIL.n62 VTAIL.n61 0.155672
R629 VTAIL.n62 VTAIL.n7 0.155672
R630 VTAIL.n69 VTAIL.n7 0.155672
R631 VTAIL.n70 VTAIL.n69 0.155672
R632 VTAIL.n70 VTAIL.n3 0.155672
R633 VTAIL.n77 VTAIL.n3 0.155672
R634 VTAIL.n245 VTAIL.n171 0.155672
R635 VTAIL.n238 VTAIL.n171 0.155672
R636 VTAIL.n238 VTAIL.n237 0.155672
R637 VTAIL.n237 VTAIL.n175 0.155672
R638 VTAIL.n230 VTAIL.n175 0.155672
R639 VTAIL.n230 VTAIL.n229 0.155672
R640 VTAIL.n229 VTAIL.n179 0.155672
R641 VTAIL.n222 VTAIL.n179 0.155672
R642 VTAIL.n222 VTAIL.n221 0.155672
R643 VTAIL.n221 VTAIL.n183 0.155672
R644 VTAIL.n213 VTAIL.n183 0.155672
R645 VTAIL.n213 VTAIL.n212 0.155672
R646 VTAIL.n212 VTAIL.n188 0.155672
R647 VTAIL.n205 VTAIL.n188 0.155672
R648 VTAIL.n205 VTAIL.n204 0.155672
R649 VTAIL.n204 VTAIL.n192 0.155672
R650 VTAIL.n197 VTAIL.n192 0.155672
R651 VTAIL.n163 VTAIL.n89 0.155672
R652 VTAIL.n156 VTAIL.n89 0.155672
R653 VTAIL.n156 VTAIL.n155 0.155672
R654 VTAIL.n155 VTAIL.n93 0.155672
R655 VTAIL.n148 VTAIL.n93 0.155672
R656 VTAIL.n148 VTAIL.n147 0.155672
R657 VTAIL.n147 VTAIL.n97 0.155672
R658 VTAIL.n140 VTAIL.n97 0.155672
R659 VTAIL.n140 VTAIL.n139 0.155672
R660 VTAIL.n139 VTAIL.n101 0.155672
R661 VTAIL.n131 VTAIL.n101 0.155672
R662 VTAIL.n131 VTAIL.n130 0.155672
R663 VTAIL.n130 VTAIL.n106 0.155672
R664 VTAIL.n123 VTAIL.n106 0.155672
R665 VTAIL.n123 VTAIL.n122 0.155672
R666 VTAIL.n122 VTAIL.n110 0.155672
R667 VTAIL.n115 VTAIL.n110 0.155672
R668 VDD1.n72 VDD1.n0 289.615
R669 VDD1.n151 VDD1.n79 289.615
R670 VDD1.n73 VDD1.n72 185
R671 VDD1.n71 VDD1.n70 185
R672 VDD1.n4 VDD1.n3 185
R673 VDD1.n65 VDD1.n64 185
R674 VDD1.n63 VDD1.n62 185
R675 VDD1.n8 VDD1.n7 185
R676 VDD1.n57 VDD1.n56 185
R677 VDD1.n55 VDD1.n54 185
R678 VDD1.n12 VDD1.n11 185
R679 VDD1.n49 VDD1.n48 185
R680 VDD1.n47 VDD1.n14 185
R681 VDD1.n46 VDD1.n45 185
R682 VDD1.n17 VDD1.n15 185
R683 VDD1.n40 VDD1.n39 185
R684 VDD1.n38 VDD1.n37 185
R685 VDD1.n21 VDD1.n20 185
R686 VDD1.n32 VDD1.n31 185
R687 VDD1.n30 VDD1.n29 185
R688 VDD1.n25 VDD1.n24 185
R689 VDD1.n103 VDD1.n102 185
R690 VDD1.n108 VDD1.n107 185
R691 VDD1.n110 VDD1.n109 185
R692 VDD1.n99 VDD1.n98 185
R693 VDD1.n116 VDD1.n115 185
R694 VDD1.n118 VDD1.n117 185
R695 VDD1.n95 VDD1.n94 185
R696 VDD1.n125 VDD1.n124 185
R697 VDD1.n126 VDD1.n93 185
R698 VDD1.n128 VDD1.n127 185
R699 VDD1.n91 VDD1.n90 185
R700 VDD1.n134 VDD1.n133 185
R701 VDD1.n136 VDD1.n135 185
R702 VDD1.n87 VDD1.n86 185
R703 VDD1.n142 VDD1.n141 185
R704 VDD1.n144 VDD1.n143 185
R705 VDD1.n83 VDD1.n82 185
R706 VDD1.n150 VDD1.n149 185
R707 VDD1.n152 VDD1.n151 185
R708 VDD1.n26 VDD1.t3 149.524
R709 VDD1.n104 VDD1.t6 149.524
R710 VDD1.n72 VDD1.n71 104.615
R711 VDD1.n71 VDD1.n3 104.615
R712 VDD1.n64 VDD1.n3 104.615
R713 VDD1.n64 VDD1.n63 104.615
R714 VDD1.n63 VDD1.n7 104.615
R715 VDD1.n56 VDD1.n7 104.615
R716 VDD1.n56 VDD1.n55 104.615
R717 VDD1.n55 VDD1.n11 104.615
R718 VDD1.n48 VDD1.n11 104.615
R719 VDD1.n48 VDD1.n47 104.615
R720 VDD1.n47 VDD1.n46 104.615
R721 VDD1.n46 VDD1.n15 104.615
R722 VDD1.n39 VDD1.n15 104.615
R723 VDD1.n39 VDD1.n38 104.615
R724 VDD1.n38 VDD1.n20 104.615
R725 VDD1.n31 VDD1.n20 104.615
R726 VDD1.n31 VDD1.n30 104.615
R727 VDD1.n30 VDD1.n24 104.615
R728 VDD1.n108 VDD1.n102 104.615
R729 VDD1.n109 VDD1.n108 104.615
R730 VDD1.n109 VDD1.n98 104.615
R731 VDD1.n116 VDD1.n98 104.615
R732 VDD1.n117 VDD1.n116 104.615
R733 VDD1.n117 VDD1.n94 104.615
R734 VDD1.n125 VDD1.n94 104.615
R735 VDD1.n126 VDD1.n125 104.615
R736 VDD1.n127 VDD1.n126 104.615
R737 VDD1.n127 VDD1.n90 104.615
R738 VDD1.n134 VDD1.n90 104.615
R739 VDD1.n135 VDD1.n134 104.615
R740 VDD1.n135 VDD1.n86 104.615
R741 VDD1.n142 VDD1.n86 104.615
R742 VDD1.n143 VDD1.n142 104.615
R743 VDD1.n143 VDD1.n82 104.615
R744 VDD1.n150 VDD1.n82 104.615
R745 VDD1.n151 VDD1.n150 104.615
R746 VDD1.n159 VDD1.n158 62.1489
R747 VDD1.n161 VDD1.n160 60.0706
R748 VDD1.n78 VDD1.n77 60.0706
R749 VDD1.n157 VDD1.n156 60.0706
R750 VDD1.t3 VDD1.n24 52.3082
R751 VDD1.t6 VDD1.n102 52.3082
R752 VDD1.n161 VDD1.n159 51.4837
R753 VDD1.n78 VDD1.n76 50.3514
R754 VDD1.n157 VDD1.n155 50.3514
R755 VDD1.n49 VDD1.n14 13.1884
R756 VDD1.n128 VDD1.n93 13.1884
R757 VDD1.n50 VDD1.n12 12.8005
R758 VDD1.n45 VDD1.n16 12.8005
R759 VDD1.n124 VDD1.n123 12.8005
R760 VDD1.n129 VDD1.n91 12.8005
R761 VDD1.n54 VDD1.n53 12.0247
R762 VDD1.n44 VDD1.n17 12.0247
R763 VDD1.n122 VDD1.n95 12.0247
R764 VDD1.n133 VDD1.n132 12.0247
R765 VDD1.n57 VDD1.n10 11.249
R766 VDD1.n41 VDD1.n40 11.249
R767 VDD1.n119 VDD1.n118 11.249
R768 VDD1.n136 VDD1.n89 11.249
R769 VDD1.n58 VDD1.n8 10.4732
R770 VDD1.n37 VDD1.n19 10.4732
R771 VDD1.n115 VDD1.n97 10.4732
R772 VDD1.n137 VDD1.n87 10.4732
R773 VDD1.n26 VDD1.n25 10.2747
R774 VDD1.n104 VDD1.n103 10.2747
R775 VDD1.n62 VDD1.n61 9.69747
R776 VDD1.n36 VDD1.n21 9.69747
R777 VDD1.n114 VDD1.n99 9.69747
R778 VDD1.n141 VDD1.n140 9.69747
R779 VDD1.n76 VDD1.n75 9.45567
R780 VDD1.n155 VDD1.n154 9.45567
R781 VDD1.n28 VDD1.n27 9.3005
R782 VDD1.n23 VDD1.n22 9.3005
R783 VDD1.n34 VDD1.n33 9.3005
R784 VDD1.n36 VDD1.n35 9.3005
R785 VDD1.n19 VDD1.n18 9.3005
R786 VDD1.n42 VDD1.n41 9.3005
R787 VDD1.n44 VDD1.n43 9.3005
R788 VDD1.n16 VDD1.n13 9.3005
R789 VDD1.n75 VDD1.n74 9.3005
R790 VDD1.n2 VDD1.n1 9.3005
R791 VDD1.n69 VDD1.n68 9.3005
R792 VDD1.n67 VDD1.n66 9.3005
R793 VDD1.n6 VDD1.n5 9.3005
R794 VDD1.n61 VDD1.n60 9.3005
R795 VDD1.n59 VDD1.n58 9.3005
R796 VDD1.n10 VDD1.n9 9.3005
R797 VDD1.n53 VDD1.n52 9.3005
R798 VDD1.n51 VDD1.n50 9.3005
R799 VDD1.n81 VDD1.n80 9.3005
R800 VDD1.n154 VDD1.n153 9.3005
R801 VDD1.n146 VDD1.n145 9.3005
R802 VDD1.n85 VDD1.n84 9.3005
R803 VDD1.n140 VDD1.n139 9.3005
R804 VDD1.n138 VDD1.n137 9.3005
R805 VDD1.n89 VDD1.n88 9.3005
R806 VDD1.n132 VDD1.n131 9.3005
R807 VDD1.n130 VDD1.n129 9.3005
R808 VDD1.n106 VDD1.n105 9.3005
R809 VDD1.n101 VDD1.n100 9.3005
R810 VDD1.n112 VDD1.n111 9.3005
R811 VDD1.n114 VDD1.n113 9.3005
R812 VDD1.n97 VDD1.n96 9.3005
R813 VDD1.n120 VDD1.n119 9.3005
R814 VDD1.n122 VDD1.n121 9.3005
R815 VDD1.n123 VDD1.n92 9.3005
R816 VDD1.n148 VDD1.n147 9.3005
R817 VDD1.n65 VDD1.n6 8.92171
R818 VDD1.n33 VDD1.n32 8.92171
R819 VDD1.n111 VDD1.n110 8.92171
R820 VDD1.n144 VDD1.n85 8.92171
R821 VDD1.n76 VDD1.n0 8.14595
R822 VDD1.n66 VDD1.n4 8.14595
R823 VDD1.n29 VDD1.n23 8.14595
R824 VDD1.n107 VDD1.n101 8.14595
R825 VDD1.n145 VDD1.n83 8.14595
R826 VDD1.n155 VDD1.n79 8.14595
R827 VDD1.n74 VDD1.n73 7.3702
R828 VDD1.n70 VDD1.n69 7.3702
R829 VDD1.n28 VDD1.n25 7.3702
R830 VDD1.n106 VDD1.n103 7.3702
R831 VDD1.n149 VDD1.n148 7.3702
R832 VDD1.n153 VDD1.n152 7.3702
R833 VDD1.n73 VDD1.n2 6.59444
R834 VDD1.n70 VDD1.n2 6.59444
R835 VDD1.n149 VDD1.n81 6.59444
R836 VDD1.n152 VDD1.n81 6.59444
R837 VDD1.n74 VDD1.n0 5.81868
R838 VDD1.n69 VDD1.n4 5.81868
R839 VDD1.n29 VDD1.n28 5.81868
R840 VDD1.n107 VDD1.n106 5.81868
R841 VDD1.n148 VDD1.n83 5.81868
R842 VDD1.n153 VDD1.n79 5.81868
R843 VDD1.n66 VDD1.n65 5.04292
R844 VDD1.n32 VDD1.n23 5.04292
R845 VDD1.n110 VDD1.n101 5.04292
R846 VDD1.n145 VDD1.n144 5.04292
R847 VDD1.n62 VDD1.n6 4.26717
R848 VDD1.n33 VDD1.n21 4.26717
R849 VDD1.n111 VDD1.n99 4.26717
R850 VDD1.n141 VDD1.n85 4.26717
R851 VDD1.n61 VDD1.n8 3.49141
R852 VDD1.n37 VDD1.n36 3.49141
R853 VDD1.n115 VDD1.n114 3.49141
R854 VDD1.n140 VDD1.n87 3.49141
R855 VDD1.n27 VDD1.n26 2.84303
R856 VDD1.n105 VDD1.n104 2.84303
R857 VDD1.n58 VDD1.n57 2.71565
R858 VDD1.n40 VDD1.n19 2.71565
R859 VDD1.n118 VDD1.n97 2.71565
R860 VDD1.n137 VDD1.n136 2.71565
R861 VDD1 VDD1.n161 2.07593
R862 VDD1.n54 VDD1.n10 1.93989
R863 VDD1.n41 VDD1.n17 1.93989
R864 VDD1.n119 VDD1.n95 1.93989
R865 VDD1.n133 VDD1.n89 1.93989
R866 VDD1.n160 VDD1.t2 1.39388
R867 VDD1.n160 VDD1.t4 1.39388
R868 VDD1.n77 VDD1.t5 1.39388
R869 VDD1.n77 VDD1.t0 1.39388
R870 VDD1.n158 VDD1.t8 1.39388
R871 VDD1.n158 VDD1.t1 1.39388
R872 VDD1.n156 VDD1.t7 1.39388
R873 VDD1.n156 VDD1.t9 1.39388
R874 VDD1.n53 VDD1.n12 1.16414
R875 VDD1.n45 VDD1.n44 1.16414
R876 VDD1.n124 VDD1.n122 1.16414
R877 VDD1.n132 VDD1.n91 1.16414
R878 VDD1 VDD1.n78 0.769897
R879 VDD1.n159 VDD1.n157 0.656361
R880 VDD1.n50 VDD1.n49 0.388379
R881 VDD1.n16 VDD1.n14 0.388379
R882 VDD1.n123 VDD1.n93 0.388379
R883 VDD1.n129 VDD1.n128 0.388379
R884 VDD1.n75 VDD1.n1 0.155672
R885 VDD1.n68 VDD1.n1 0.155672
R886 VDD1.n68 VDD1.n67 0.155672
R887 VDD1.n67 VDD1.n5 0.155672
R888 VDD1.n60 VDD1.n5 0.155672
R889 VDD1.n60 VDD1.n59 0.155672
R890 VDD1.n59 VDD1.n9 0.155672
R891 VDD1.n52 VDD1.n9 0.155672
R892 VDD1.n52 VDD1.n51 0.155672
R893 VDD1.n51 VDD1.n13 0.155672
R894 VDD1.n43 VDD1.n13 0.155672
R895 VDD1.n43 VDD1.n42 0.155672
R896 VDD1.n42 VDD1.n18 0.155672
R897 VDD1.n35 VDD1.n18 0.155672
R898 VDD1.n35 VDD1.n34 0.155672
R899 VDD1.n34 VDD1.n22 0.155672
R900 VDD1.n27 VDD1.n22 0.155672
R901 VDD1.n105 VDD1.n100 0.155672
R902 VDD1.n112 VDD1.n100 0.155672
R903 VDD1.n113 VDD1.n112 0.155672
R904 VDD1.n113 VDD1.n96 0.155672
R905 VDD1.n120 VDD1.n96 0.155672
R906 VDD1.n121 VDD1.n120 0.155672
R907 VDD1.n121 VDD1.n92 0.155672
R908 VDD1.n130 VDD1.n92 0.155672
R909 VDD1.n131 VDD1.n130 0.155672
R910 VDD1.n131 VDD1.n88 0.155672
R911 VDD1.n138 VDD1.n88 0.155672
R912 VDD1.n139 VDD1.n138 0.155672
R913 VDD1.n139 VDD1.n84 0.155672
R914 VDD1.n146 VDD1.n84 0.155672
R915 VDD1.n147 VDD1.n146 0.155672
R916 VDD1.n147 VDD1.n80 0.155672
R917 VDD1.n154 VDD1.n80 0.155672
R918 B.n864 B.n863 585
R919 B.n866 B.n179 585
R920 B.n869 B.n868 585
R921 B.n870 B.n178 585
R922 B.n872 B.n871 585
R923 B.n874 B.n177 585
R924 B.n877 B.n876 585
R925 B.n878 B.n176 585
R926 B.n880 B.n879 585
R927 B.n882 B.n175 585
R928 B.n885 B.n884 585
R929 B.n886 B.n174 585
R930 B.n888 B.n887 585
R931 B.n890 B.n173 585
R932 B.n893 B.n892 585
R933 B.n894 B.n172 585
R934 B.n896 B.n895 585
R935 B.n898 B.n171 585
R936 B.n901 B.n900 585
R937 B.n902 B.n170 585
R938 B.n904 B.n903 585
R939 B.n906 B.n169 585
R940 B.n909 B.n908 585
R941 B.n910 B.n168 585
R942 B.n912 B.n911 585
R943 B.n914 B.n167 585
R944 B.n917 B.n916 585
R945 B.n918 B.n166 585
R946 B.n920 B.n919 585
R947 B.n922 B.n165 585
R948 B.n925 B.n924 585
R949 B.n926 B.n164 585
R950 B.n928 B.n927 585
R951 B.n930 B.n163 585
R952 B.n933 B.n932 585
R953 B.n934 B.n162 585
R954 B.n936 B.n935 585
R955 B.n938 B.n161 585
R956 B.n941 B.n940 585
R957 B.n942 B.n160 585
R958 B.n944 B.n943 585
R959 B.n946 B.n159 585
R960 B.n949 B.n948 585
R961 B.n950 B.n158 585
R962 B.n952 B.n951 585
R963 B.n954 B.n157 585
R964 B.n956 B.n955 585
R965 B.n958 B.n957 585
R966 B.n961 B.n960 585
R967 B.n962 B.n152 585
R968 B.n964 B.n963 585
R969 B.n966 B.n151 585
R970 B.n969 B.n968 585
R971 B.n970 B.n150 585
R972 B.n972 B.n971 585
R973 B.n974 B.n149 585
R974 B.n977 B.n976 585
R975 B.n978 B.n146 585
R976 B.n981 B.n980 585
R977 B.n983 B.n145 585
R978 B.n986 B.n985 585
R979 B.n987 B.n144 585
R980 B.n989 B.n988 585
R981 B.n991 B.n143 585
R982 B.n994 B.n993 585
R983 B.n995 B.n142 585
R984 B.n997 B.n996 585
R985 B.n999 B.n141 585
R986 B.n1002 B.n1001 585
R987 B.n1003 B.n140 585
R988 B.n1005 B.n1004 585
R989 B.n1007 B.n139 585
R990 B.n1010 B.n1009 585
R991 B.n1011 B.n138 585
R992 B.n1013 B.n1012 585
R993 B.n1015 B.n137 585
R994 B.n1018 B.n1017 585
R995 B.n1019 B.n136 585
R996 B.n1021 B.n1020 585
R997 B.n1023 B.n135 585
R998 B.n1026 B.n1025 585
R999 B.n1027 B.n134 585
R1000 B.n1029 B.n1028 585
R1001 B.n1031 B.n133 585
R1002 B.n1034 B.n1033 585
R1003 B.n1035 B.n132 585
R1004 B.n1037 B.n1036 585
R1005 B.n1039 B.n131 585
R1006 B.n1042 B.n1041 585
R1007 B.n1043 B.n130 585
R1008 B.n1045 B.n1044 585
R1009 B.n1047 B.n129 585
R1010 B.n1050 B.n1049 585
R1011 B.n1051 B.n128 585
R1012 B.n1053 B.n1052 585
R1013 B.n1055 B.n127 585
R1014 B.n1058 B.n1057 585
R1015 B.n1059 B.n126 585
R1016 B.n1061 B.n1060 585
R1017 B.n1063 B.n125 585
R1018 B.n1066 B.n1065 585
R1019 B.n1067 B.n124 585
R1020 B.n1069 B.n1068 585
R1021 B.n1071 B.n123 585
R1022 B.n1074 B.n1073 585
R1023 B.n1075 B.n122 585
R1024 B.n862 B.n120 585
R1025 B.n1078 B.n120 585
R1026 B.n861 B.n119 585
R1027 B.n1079 B.n119 585
R1028 B.n860 B.n118 585
R1029 B.n1080 B.n118 585
R1030 B.n859 B.n858 585
R1031 B.n858 B.n114 585
R1032 B.n857 B.n113 585
R1033 B.n1086 B.n113 585
R1034 B.n856 B.n112 585
R1035 B.n1087 B.n112 585
R1036 B.n855 B.n111 585
R1037 B.n1088 B.n111 585
R1038 B.n854 B.n853 585
R1039 B.n853 B.n107 585
R1040 B.n852 B.n106 585
R1041 B.n1094 B.n106 585
R1042 B.n851 B.n105 585
R1043 B.n1095 B.n105 585
R1044 B.n850 B.n104 585
R1045 B.n1096 B.n104 585
R1046 B.n849 B.n848 585
R1047 B.n848 B.n100 585
R1048 B.n847 B.n99 585
R1049 B.n1102 B.n99 585
R1050 B.n846 B.n98 585
R1051 B.n1103 B.n98 585
R1052 B.n845 B.n97 585
R1053 B.n1104 B.n97 585
R1054 B.n844 B.n843 585
R1055 B.n843 B.n93 585
R1056 B.n842 B.n92 585
R1057 B.n1110 B.n92 585
R1058 B.n841 B.n91 585
R1059 B.n1111 B.n91 585
R1060 B.n840 B.n90 585
R1061 B.n1112 B.n90 585
R1062 B.n839 B.n838 585
R1063 B.n838 B.n86 585
R1064 B.n837 B.n85 585
R1065 B.n1118 B.n85 585
R1066 B.n836 B.n84 585
R1067 B.n1119 B.n84 585
R1068 B.n835 B.n83 585
R1069 B.n1120 B.n83 585
R1070 B.n834 B.n833 585
R1071 B.n833 B.n79 585
R1072 B.n832 B.n78 585
R1073 B.n1126 B.n78 585
R1074 B.n831 B.n77 585
R1075 B.n1127 B.n77 585
R1076 B.n830 B.n76 585
R1077 B.n1128 B.n76 585
R1078 B.n829 B.n828 585
R1079 B.n828 B.n72 585
R1080 B.n827 B.n71 585
R1081 B.n1134 B.n71 585
R1082 B.n826 B.n70 585
R1083 B.n1135 B.n70 585
R1084 B.n825 B.n69 585
R1085 B.n1136 B.n69 585
R1086 B.n824 B.n823 585
R1087 B.n823 B.n65 585
R1088 B.n822 B.n64 585
R1089 B.n1142 B.n64 585
R1090 B.n821 B.n63 585
R1091 B.n1143 B.n63 585
R1092 B.n820 B.n62 585
R1093 B.n1144 B.n62 585
R1094 B.n819 B.n818 585
R1095 B.n818 B.n58 585
R1096 B.n817 B.n57 585
R1097 B.n1150 B.n57 585
R1098 B.n816 B.n56 585
R1099 B.n1151 B.n56 585
R1100 B.n815 B.n55 585
R1101 B.n1152 B.n55 585
R1102 B.n814 B.n813 585
R1103 B.n813 B.n51 585
R1104 B.n812 B.n50 585
R1105 B.n1158 B.n50 585
R1106 B.n811 B.n49 585
R1107 B.n1159 B.n49 585
R1108 B.n810 B.n48 585
R1109 B.n1160 B.n48 585
R1110 B.n809 B.n808 585
R1111 B.n808 B.n44 585
R1112 B.n807 B.n43 585
R1113 B.n1166 B.n43 585
R1114 B.n806 B.n42 585
R1115 B.n1167 B.n42 585
R1116 B.n805 B.n41 585
R1117 B.n1168 B.n41 585
R1118 B.n804 B.n803 585
R1119 B.n803 B.n37 585
R1120 B.n802 B.n36 585
R1121 B.n1174 B.n36 585
R1122 B.n801 B.n35 585
R1123 B.n1175 B.n35 585
R1124 B.n800 B.n34 585
R1125 B.n1176 B.n34 585
R1126 B.n799 B.n798 585
R1127 B.n798 B.n30 585
R1128 B.n797 B.n29 585
R1129 B.n1182 B.n29 585
R1130 B.n796 B.n28 585
R1131 B.n1183 B.n28 585
R1132 B.n795 B.n27 585
R1133 B.n1184 B.n27 585
R1134 B.n794 B.n793 585
R1135 B.n793 B.n23 585
R1136 B.n792 B.n22 585
R1137 B.n1190 B.n22 585
R1138 B.n791 B.n21 585
R1139 B.n1191 B.n21 585
R1140 B.n790 B.n20 585
R1141 B.n1192 B.n20 585
R1142 B.n789 B.n788 585
R1143 B.n788 B.n16 585
R1144 B.n787 B.n15 585
R1145 B.n1198 B.n15 585
R1146 B.n786 B.n14 585
R1147 B.n1199 B.n14 585
R1148 B.n785 B.n13 585
R1149 B.n1200 B.n13 585
R1150 B.n784 B.n783 585
R1151 B.n783 B.n12 585
R1152 B.n782 B.n781 585
R1153 B.n782 B.n8 585
R1154 B.n780 B.n7 585
R1155 B.n1207 B.n7 585
R1156 B.n779 B.n6 585
R1157 B.n1208 B.n6 585
R1158 B.n778 B.n5 585
R1159 B.n1209 B.n5 585
R1160 B.n777 B.n776 585
R1161 B.n776 B.n4 585
R1162 B.n775 B.n180 585
R1163 B.n775 B.n774 585
R1164 B.n765 B.n181 585
R1165 B.n182 B.n181 585
R1166 B.n767 B.n766 585
R1167 B.n768 B.n767 585
R1168 B.n764 B.n187 585
R1169 B.n187 B.n186 585
R1170 B.n763 B.n762 585
R1171 B.n762 B.n761 585
R1172 B.n189 B.n188 585
R1173 B.n190 B.n189 585
R1174 B.n754 B.n753 585
R1175 B.n755 B.n754 585
R1176 B.n752 B.n195 585
R1177 B.n195 B.n194 585
R1178 B.n751 B.n750 585
R1179 B.n750 B.n749 585
R1180 B.n197 B.n196 585
R1181 B.n198 B.n197 585
R1182 B.n742 B.n741 585
R1183 B.n743 B.n742 585
R1184 B.n740 B.n203 585
R1185 B.n203 B.n202 585
R1186 B.n739 B.n738 585
R1187 B.n738 B.n737 585
R1188 B.n205 B.n204 585
R1189 B.n206 B.n205 585
R1190 B.n730 B.n729 585
R1191 B.n731 B.n730 585
R1192 B.n728 B.n211 585
R1193 B.n211 B.n210 585
R1194 B.n727 B.n726 585
R1195 B.n726 B.n725 585
R1196 B.n213 B.n212 585
R1197 B.n214 B.n213 585
R1198 B.n718 B.n717 585
R1199 B.n719 B.n718 585
R1200 B.n716 B.n219 585
R1201 B.n219 B.n218 585
R1202 B.n715 B.n714 585
R1203 B.n714 B.n713 585
R1204 B.n221 B.n220 585
R1205 B.n222 B.n221 585
R1206 B.n706 B.n705 585
R1207 B.n707 B.n706 585
R1208 B.n704 B.n227 585
R1209 B.n227 B.n226 585
R1210 B.n703 B.n702 585
R1211 B.n702 B.n701 585
R1212 B.n229 B.n228 585
R1213 B.n230 B.n229 585
R1214 B.n694 B.n693 585
R1215 B.n695 B.n694 585
R1216 B.n692 B.n235 585
R1217 B.n235 B.n234 585
R1218 B.n691 B.n690 585
R1219 B.n690 B.n689 585
R1220 B.n237 B.n236 585
R1221 B.n238 B.n237 585
R1222 B.n682 B.n681 585
R1223 B.n683 B.n682 585
R1224 B.n680 B.n243 585
R1225 B.n243 B.n242 585
R1226 B.n679 B.n678 585
R1227 B.n678 B.n677 585
R1228 B.n245 B.n244 585
R1229 B.n246 B.n245 585
R1230 B.n670 B.n669 585
R1231 B.n671 B.n670 585
R1232 B.n668 B.n251 585
R1233 B.n251 B.n250 585
R1234 B.n667 B.n666 585
R1235 B.n666 B.n665 585
R1236 B.n253 B.n252 585
R1237 B.n254 B.n253 585
R1238 B.n658 B.n657 585
R1239 B.n659 B.n658 585
R1240 B.n656 B.n259 585
R1241 B.n259 B.n258 585
R1242 B.n655 B.n654 585
R1243 B.n654 B.n653 585
R1244 B.n261 B.n260 585
R1245 B.n262 B.n261 585
R1246 B.n646 B.n645 585
R1247 B.n647 B.n646 585
R1248 B.n644 B.n266 585
R1249 B.n270 B.n266 585
R1250 B.n643 B.n642 585
R1251 B.n642 B.n641 585
R1252 B.n268 B.n267 585
R1253 B.n269 B.n268 585
R1254 B.n634 B.n633 585
R1255 B.n635 B.n634 585
R1256 B.n632 B.n275 585
R1257 B.n275 B.n274 585
R1258 B.n631 B.n630 585
R1259 B.n630 B.n629 585
R1260 B.n277 B.n276 585
R1261 B.n278 B.n277 585
R1262 B.n622 B.n621 585
R1263 B.n623 B.n622 585
R1264 B.n620 B.n283 585
R1265 B.n283 B.n282 585
R1266 B.n619 B.n618 585
R1267 B.n618 B.n617 585
R1268 B.n285 B.n284 585
R1269 B.n286 B.n285 585
R1270 B.n610 B.n609 585
R1271 B.n611 B.n610 585
R1272 B.n608 B.n291 585
R1273 B.n291 B.n290 585
R1274 B.n607 B.n606 585
R1275 B.n606 B.n605 585
R1276 B.n293 B.n292 585
R1277 B.n294 B.n293 585
R1278 B.n598 B.n597 585
R1279 B.n599 B.n598 585
R1280 B.n596 B.n299 585
R1281 B.n299 B.n298 585
R1282 B.n595 B.n594 585
R1283 B.n594 B.n593 585
R1284 B.n301 B.n300 585
R1285 B.n302 B.n301 585
R1286 B.n586 B.n585 585
R1287 B.n587 B.n586 585
R1288 B.n584 B.n307 585
R1289 B.n307 B.n306 585
R1290 B.n583 B.n582 585
R1291 B.n582 B.n581 585
R1292 B.n578 B.n311 585
R1293 B.n577 B.n576 585
R1294 B.n574 B.n312 585
R1295 B.n574 B.n310 585
R1296 B.n573 B.n572 585
R1297 B.n571 B.n570 585
R1298 B.n569 B.n314 585
R1299 B.n567 B.n566 585
R1300 B.n565 B.n315 585
R1301 B.n564 B.n563 585
R1302 B.n561 B.n316 585
R1303 B.n559 B.n558 585
R1304 B.n557 B.n317 585
R1305 B.n556 B.n555 585
R1306 B.n553 B.n318 585
R1307 B.n551 B.n550 585
R1308 B.n549 B.n319 585
R1309 B.n548 B.n547 585
R1310 B.n545 B.n320 585
R1311 B.n543 B.n542 585
R1312 B.n541 B.n321 585
R1313 B.n540 B.n539 585
R1314 B.n537 B.n322 585
R1315 B.n535 B.n534 585
R1316 B.n533 B.n323 585
R1317 B.n532 B.n531 585
R1318 B.n529 B.n324 585
R1319 B.n527 B.n526 585
R1320 B.n525 B.n325 585
R1321 B.n524 B.n523 585
R1322 B.n521 B.n326 585
R1323 B.n519 B.n518 585
R1324 B.n517 B.n327 585
R1325 B.n516 B.n515 585
R1326 B.n513 B.n328 585
R1327 B.n511 B.n510 585
R1328 B.n509 B.n329 585
R1329 B.n508 B.n507 585
R1330 B.n505 B.n330 585
R1331 B.n503 B.n502 585
R1332 B.n501 B.n331 585
R1333 B.n500 B.n499 585
R1334 B.n497 B.n332 585
R1335 B.n495 B.n494 585
R1336 B.n493 B.n333 585
R1337 B.n492 B.n491 585
R1338 B.n489 B.n334 585
R1339 B.n487 B.n486 585
R1340 B.n485 B.n335 585
R1341 B.n483 B.n482 585
R1342 B.n480 B.n338 585
R1343 B.n478 B.n477 585
R1344 B.n476 B.n339 585
R1345 B.n475 B.n474 585
R1346 B.n472 B.n340 585
R1347 B.n470 B.n469 585
R1348 B.n468 B.n341 585
R1349 B.n467 B.n466 585
R1350 B.n464 B.n342 585
R1351 B.n462 B.n461 585
R1352 B.n460 B.n343 585
R1353 B.n459 B.n458 585
R1354 B.n456 B.n347 585
R1355 B.n454 B.n453 585
R1356 B.n452 B.n348 585
R1357 B.n451 B.n450 585
R1358 B.n448 B.n349 585
R1359 B.n446 B.n445 585
R1360 B.n444 B.n350 585
R1361 B.n443 B.n442 585
R1362 B.n440 B.n351 585
R1363 B.n438 B.n437 585
R1364 B.n436 B.n352 585
R1365 B.n435 B.n434 585
R1366 B.n432 B.n353 585
R1367 B.n430 B.n429 585
R1368 B.n428 B.n354 585
R1369 B.n427 B.n426 585
R1370 B.n424 B.n355 585
R1371 B.n422 B.n421 585
R1372 B.n420 B.n356 585
R1373 B.n419 B.n418 585
R1374 B.n416 B.n357 585
R1375 B.n414 B.n413 585
R1376 B.n412 B.n358 585
R1377 B.n411 B.n410 585
R1378 B.n408 B.n359 585
R1379 B.n406 B.n405 585
R1380 B.n404 B.n360 585
R1381 B.n403 B.n402 585
R1382 B.n400 B.n361 585
R1383 B.n398 B.n397 585
R1384 B.n396 B.n362 585
R1385 B.n395 B.n394 585
R1386 B.n392 B.n363 585
R1387 B.n390 B.n389 585
R1388 B.n388 B.n364 585
R1389 B.n387 B.n386 585
R1390 B.n384 B.n365 585
R1391 B.n382 B.n381 585
R1392 B.n380 B.n366 585
R1393 B.n379 B.n378 585
R1394 B.n376 B.n367 585
R1395 B.n374 B.n373 585
R1396 B.n372 B.n368 585
R1397 B.n371 B.n370 585
R1398 B.n309 B.n308 585
R1399 B.n310 B.n309 585
R1400 B.n580 B.n579 585
R1401 B.n581 B.n580 585
R1402 B.n305 B.n304 585
R1403 B.n306 B.n305 585
R1404 B.n589 B.n588 585
R1405 B.n588 B.n587 585
R1406 B.n590 B.n303 585
R1407 B.n303 B.n302 585
R1408 B.n592 B.n591 585
R1409 B.n593 B.n592 585
R1410 B.n297 B.n296 585
R1411 B.n298 B.n297 585
R1412 B.n601 B.n600 585
R1413 B.n600 B.n599 585
R1414 B.n602 B.n295 585
R1415 B.n295 B.n294 585
R1416 B.n604 B.n603 585
R1417 B.n605 B.n604 585
R1418 B.n289 B.n288 585
R1419 B.n290 B.n289 585
R1420 B.n613 B.n612 585
R1421 B.n612 B.n611 585
R1422 B.n614 B.n287 585
R1423 B.n287 B.n286 585
R1424 B.n616 B.n615 585
R1425 B.n617 B.n616 585
R1426 B.n281 B.n280 585
R1427 B.n282 B.n281 585
R1428 B.n625 B.n624 585
R1429 B.n624 B.n623 585
R1430 B.n626 B.n279 585
R1431 B.n279 B.n278 585
R1432 B.n628 B.n627 585
R1433 B.n629 B.n628 585
R1434 B.n273 B.n272 585
R1435 B.n274 B.n273 585
R1436 B.n637 B.n636 585
R1437 B.n636 B.n635 585
R1438 B.n638 B.n271 585
R1439 B.n271 B.n269 585
R1440 B.n640 B.n639 585
R1441 B.n641 B.n640 585
R1442 B.n265 B.n264 585
R1443 B.n270 B.n265 585
R1444 B.n649 B.n648 585
R1445 B.n648 B.n647 585
R1446 B.n650 B.n263 585
R1447 B.n263 B.n262 585
R1448 B.n652 B.n651 585
R1449 B.n653 B.n652 585
R1450 B.n257 B.n256 585
R1451 B.n258 B.n257 585
R1452 B.n661 B.n660 585
R1453 B.n660 B.n659 585
R1454 B.n662 B.n255 585
R1455 B.n255 B.n254 585
R1456 B.n664 B.n663 585
R1457 B.n665 B.n664 585
R1458 B.n249 B.n248 585
R1459 B.n250 B.n249 585
R1460 B.n673 B.n672 585
R1461 B.n672 B.n671 585
R1462 B.n674 B.n247 585
R1463 B.n247 B.n246 585
R1464 B.n676 B.n675 585
R1465 B.n677 B.n676 585
R1466 B.n241 B.n240 585
R1467 B.n242 B.n241 585
R1468 B.n685 B.n684 585
R1469 B.n684 B.n683 585
R1470 B.n686 B.n239 585
R1471 B.n239 B.n238 585
R1472 B.n688 B.n687 585
R1473 B.n689 B.n688 585
R1474 B.n233 B.n232 585
R1475 B.n234 B.n233 585
R1476 B.n697 B.n696 585
R1477 B.n696 B.n695 585
R1478 B.n698 B.n231 585
R1479 B.n231 B.n230 585
R1480 B.n700 B.n699 585
R1481 B.n701 B.n700 585
R1482 B.n225 B.n224 585
R1483 B.n226 B.n225 585
R1484 B.n709 B.n708 585
R1485 B.n708 B.n707 585
R1486 B.n710 B.n223 585
R1487 B.n223 B.n222 585
R1488 B.n712 B.n711 585
R1489 B.n713 B.n712 585
R1490 B.n217 B.n216 585
R1491 B.n218 B.n217 585
R1492 B.n721 B.n720 585
R1493 B.n720 B.n719 585
R1494 B.n722 B.n215 585
R1495 B.n215 B.n214 585
R1496 B.n724 B.n723 585
R1497 B.n725 B.n724 585
R1498 B.n209 B.n208 585
R1499 B.n210 B.n209 585
R1500 B.n733 B.n732 585
R1501 B.n732 B.n731 585
R1502 B.n734 B.n207 585
R1503 B.n207 B.n206 585
R1504 B.n736 B.n735 585
R1505 B.n737 B.n736 585
R1506 B.n201 B.n200 585
R1507 B.n202 B.n201 585
R1508 B.n745 B.n744 585
R1509 B.n744 B.n743 585
R1510 B.n746 B.n199 585
R1511 B.n199 B.n198 585
R1512 B.n748 B.n747 585
R1513 B.n749 B.n748 585
R1514 B.n193 B.n192 585
R1515 B.n194 B.n193 585
R1516 B.n757 B.n756 585
R1517 B.n756 B.n755 585
R1518 B.n758 B.n191 585
R1519 B.n191 B.n190 585
R1520 B.n760 B.n759 585
R1521 B.n761 B.n760 585
R1522 B.n185 B.n184 585
R1523 B.n186 B.n185 585
R1524 B.n770 B.n769 585
R1525 B.n769 B.n768 585
R1526 B.n771 B.n183 585
R1527 B.n183 B.n182 585
R1528 B.n773 B.n772 585
R1529 B.n774 B.n773 585
R1530 B.n3 B.n0 585
R1531 B.n4 B.n3 585
R1532 B.n1206 B.n1 585
R1533 B.n1207 B.n1206 585
R1534 B.n1205 B.n1204 585
R1535 B.n1205 B.n8 585
R1536 B.n1203 B.n9 585
R1537 B.n12 B.n9 585
R1538 B.n1202 B.n1201 585
R1539 B.n1201 B.n1200 585
R1540 B.n11 B.n10 585
R1541 B.n1199 B.n11 585
R1542 B.n1197 B.n1196 585
R1543 B.n1198 B.n1197 585
R1544 B.n1195 B.n17 585
R1545 B.n17 B.n16 585
R1546 B.n1194 B.n1193 585
R1547 B.n1193 B.n1192 585
R1548 B.n19 B.n18 585
R1549 B.n1191 B.n19 585
R1550 B.n1189 B.n1188 585
R1551 B.n1190 B.n1189 585
R1552 B.n1187 B.n24 585
R1553 B.n24 B.n23 585
R1554 B.n1186 B.n1185 585
R1555 B.n1185 B.n1184 585
R1556 B.n26 B.n25 585
R1557 B.n1183 B.n26 585
R1558 B.n1181 B.n1180 585
R1559 B.n1182 B.n1181 585
R1560 B.n1179 B.n31 585
R1561 B.n31 B.n30 585
R1562 B.n1178 B.n1177 585
R1563 B.n1177 B.n1176 585
R1564 B.n33 B.n32 585
R1565 B.n1175 B.n33 585
R1566 B.n1173 B.n1172 585
R1567 B.n1174 B.n1173 585
R1568 B.n1171 B.n38 585
R1569 B.n38 B.n37 585
R1570 B.n1170 B.n1169 585
R1571 B.n1169 B.n1168 585
R1572 B.n40 B.n39 585
R1573 B.n1167 B.n40 585
R1574 B.n1165 B.n1164 585
R1575 B.n1166 B.n1165 585
R1576 B.n1163 B.n45 585
R1577 B.n45 B.n44 585
R1578 B.n1162 B.n1161 585
R1579 B.n1161 B.n1160 585
R1580 B.n47 B.n46 585
R1581 B.n1159 B.n47 585
R1582 B.n1157 B.n1156 585
R1583 B.n1158 B.n1157 585
R1584 B.n1155 B.n52 585
R1585 B.n52 B.n51 585
R1586 B.n1154 B.n1153 585
R1587 B.n1153 B.n1152 585
R1588 B.n54 B.n53 585
R1589 B.n1151 B.n54 585
R1590 B.n1149 B.n1148 585
R1591 B.n1150 B.n1149 585
R1592 B.n1147 B.n59 585
R1593 B.n59 B.n58 585
R1594 B.n1146 B.n1145 585
R1595 B.n1145 B.n1144 585
R1596 B.n61 B.n60 585
R1597 B.n1143 B.n61 585
R1598 B.n1141 B.n1140 585
R1599 B.n1142 B.n1141 585
R1600 B.n1139 B.n66 585
R1601 B.n66 B.n65 585
R1602 B.n1138 B.n1137 585
R1603 B.n1137 B.n1136 585
R1604 B.n68 B.n67 585
R1605 B.n1135 B.n68 585
R1606 B.n1133 B.n1132 585
R1607 B.n1134 B.n1133 585
R1608 B.n1131 B.n73 585
R1609 B.n73 B.n72 585
R1610 B.n1130 B.n1129 585
R1611 B.n1129 B.n1128 585
R1612 B.n75 B.n74 585
R1613 B.n1127 B.n75 585
R1614 B.n1125 B.n1124 585
R1615 B.n1126 B.n1125 585
R1616 B.n1123 B.n80 585
R1617 B.n80 B.n79 585
R1618 B.n1122 B.n1121 585
R1619 B.n1121 B.n1120 585
R1620 B.n82 B.n81 585
R1621 B.n1119 B.n82 585
R1622 B.n1117 B.n1116 585
R1623 B.n1118 B.n1117 585
R1624 B.n1115 B.n87 585
R1625 B.n87 B.n86 585
R1626 B.n1114 B.n1113 585
R1627 B.n1113 B.n1112 585
R1628 B.n89 B.n88 585
R1629 B.n1111 B.n89 585
R1630 B.n1109 B.n1108 585
R1631 B.n1110 B.n1109 585
R1632 B.n1107 B.n94 585
R1633 B.n94 B.n93 585
R1634 B.n1106 B.n1105 585
R1635 B.n1105 B.n1104 585
R1636 B.n96 B.n95 585
R1637 B.n1103 B.n96 585
R1638 B.n1101 B.n1100 585
R1639 B.n1102 B.n1101 585
R1640 B.n1099 B.n101 585
R1641 B.n101 B.n100 585
R1642 B.n1098 B.n1097 585
R1643 B.n1097 B.n1096 585
R1644 B.n103 B.n102 585
R1645 B.n1095 B.n103 585
R1646 B.n1093 B.n1092 585
R1647 B.n1094 B.n1093 585
R1648 B.n1091 B.n108 585
R1649 B.n108 B.n107 585
R1650 B.n1090 B.n1089 585
R1651 B.n1089 B.n1088 585
R1652 B.n110 B.n109 585
R1653 B.n1087 B.n110 585
R1654 B.n1085 B.n1084 585
R1655 B.n1086 B.n1085 585
R1656 B.n1083 B.n115 585
R1657 B.n115 B.n114 585
R1658 B.n1082 B.n1081 585
R1659 B.n1081 B.n1080 585
R1660 B.n117 B.n116 585
R1661 B.n1079 B.n117 585
R1662 B.n1077 B.n1076 585
R1663 B.n1078 B.n1077 585
R1664 B.n1210 B.n1209 585
R1665 B.n1208 B.n2 585
R1666 B.n1077 B.n122 458.866
R1667 B.n864 B.n120 458.866
R1668 B.n582 B.n309 458.866
R1669 B.n580 B.n311 458.866
R1670 B.n153 B.t22 384.442
R1671 B.n344 B.t20 384.442
R1672 B.n147 B.t16 384.442
R1673 B.n336 B.t13 384.442
R1674 B.n147 B.t14 323.851
R1675 B.n153 B.t21 323.851
R1676 B.n344 B.t18 323.851
R1677 B.n336 B.t10 323.851
R1678 B.n154 B.t23 320.442
R1679 B.n345 B.t19 320.442
R1680 B.n148 B.t17 320.442
R1681 B.n337 B.t12 320.442
R1682 B.n865 B.n121 256.663
R1683 B.n867 B.n121 256.663
R1684 B.n873 B.n121 256.663
R1685 B.n875 B.n121 256.663
R1686 B.n881 B.n121 256.663
R1687 B.n883 B.n121 256.663
R1688 B.n889 B.n121 256.663
R1689 B.n891 B.n121 256.663
R1690 B.n897 B.n121 256.663
R1691 B.n899 B.n121 256.663
R1692 B.n905 B.n121 256.663
R1693 B.n907 B.n121 256.663
R1694 B.n913 B.n121 256.663
R1695 B.n915 B.n121 256.663
R1696 B.n921 B.n121 256.663
R1697 B.n923 B.n121 256.663
R1698 B.n929 B.n121 256.663
R1699 B.n931 B.n121 256.663
R1700 B.n937 B.n121 256.663
R1701 B.n939 B.n121 256.663
R1702 B.n945 B.n121 256.663
R1703 B.n947 B.n121 256.663
R1704 B.n953 B.n121 256.663
R1705 B.n156 B.n121 256.663
R1706 B.n959 B.n121 256.663
R1707 B.n965 B.n121 256.663
R1708 B.n967 B.n121 256.663
R1709 B.n973 B.n121 256.663
R1710 B.n975 B.n121 256.663
R1711 B.n982 B.n121 256.663
R1712 B.n984 B.n121 256.663
R1713 B.n990 B.n121 256.663
R1714 B.n992 B.n121 256.663
R1715 B.n998 B.n121 256.663
R1716 B.n1000 B.n121 256.663
R1717 B.n1006 B.n121 256.663
R1718 B.n1008 B.n121 256.663
R1719 B.n1014 B.n121 256.663
R1720 B.n1016 B.n121 256.663
R1721 B.n1022 B.n121 256.663
R1722 B.n1024 B.n121 256.663
R1723 B.n1030 B.n121 256.663
R1724 B.n1032 B.n121 256.663
R1725 B.n1038 B.n121 256.663
R1726 B.n1040 B.n121 256.663
R1727 B.n1046 B.n121 256.663
R1728 B.n1048 B.n121 256.663
R1729 B.n1054 B.n121 256.663
R1730 B.n1056 B.n121 256.663
R1731 B.n1062 B.n121 256.663
R1732 B.n1064 B.n121 256.663
R1733 B.n1070 B.n121 256.663
R1734 B.n1072 B.n121 256.663
R1735 B.n575 B.n310 256.663
R1736 B.n313 B.n310 256.663
R1737 B.n568 B.n310 256.663
R1738 B.n562 B.n310 256.663
R1739 B.n560 B.n310 256.663
R1740 B.n554 B.n310 256.663
R1741 B.n552 B.n310 256.663
R1742 B.n546 B.n310 256.663
R1743 B.n544 B.n310 256.663
R1744 B.n538 B.n310 256.663
R1745 B.n536 B.n310 256.663
R1746 B.n530 B.n310 256.663
R1747 B.n528 B.n310 256.663
R1748 B.n522 B.n310 256.663
R1749 B.n520 B.n310 256.663
R1750 B.n514 B.n310 256.663
R1751 B.n512 B.n310 256.663
R1752 B.n506 B.n310 256.663
R1753 B.n504 B.n310 256.663
R1754 B.n498 B.n310 256.663
R1755 B.n496 B.n310 256.663
R1756 B.n490 B.n310 256.663
R1757 B.n488 B.n310 256.663
R1758 B.n481 B.n310 256.663
R1759 B.n479 B.n310 256.663
R1760 B.n473 B.n310 256.663
R1761 B.n471 B.n310 256.663
R1762 B.n465 B.n310 256.663
R1763 B.n463 B.n310 256.663
R1764 B.n457 B.n310 256.663
R1765 B.n455 B.n310 256.663
R1766 B.n449 B.n310 256.663
R1767 B.n447 B.n310 256.663
R1768 B.n441 B.n310 256.663
R1769 B.n439 B.n310 256.663
R1770 B.n433 B.n310 256.663
R1771 B.n431 B.n310 256.663
R1772 B.n425 B.n310 256.663
R1773 B.n423 B.n310 256.663
R1774 B.n417 B.n310 256.663
R1775 B.n415 B.n310 256.663
R1776 B.n409 B.n310 256.663
R1777 B.n407 B.n310 256.663
R1778 B.n401 B.n310 256.663
R1779 B.n399 B.n310 256.663
R1780 B.n393 B.n310 256.663
R1781 B.n391 B.n310 256.663
R1782 B.n385 B.n310 256.663
R1783 B.n383 B.n310 256.663
R1784 B.n377 B.n310 256.663
R1785 B.n375 B.n310 256.663
R1786 B.n369 B.n310 256.663
R1787 B.n1212 B.n1211 256.663
R1788 B.n1073 B.n1071 163.367
R1789 B.n1069 B.n124 163.367
R1790 B.n1065 B.n1063 163.367
R1791 B.n1061 B.n126 163.367
R1792 B.n1057 B.n1055 163.367
R1793 B.n1053 B.n128 163.367
R1794 B.n1049 B.n1047 163.367
R1795 B.n1045 B.n130 163.367
R1796 B.n1041 B.n1039 163.367
R1797 B.n1037 B.n132 163.367
R1798 B.n1033 B.n1031 163.367
R1799 B.n1029 B.n134 163.367
R1800 B.n1025 B.n1023 163.367
R1801 B.n1021 B.n136 163.367
R1802 B.n1017 B.n1015 163.367
R1803 B.n1013 B.n138 163.367
R1804 B.n1009 B.n1007 163.367
R1805 B.n1005 B.n140 163.367
R1806 B.n1001 B.n999 163.367
R1807 B.n997 B.n142 163.367
R1808 B.n993 B.n991 163.367
R1809 B.n989 B.n144 163.367
R1810 B.n985 B.n983 163.367
R1811 B.n981 B.n146 163.367
R1812 B.n976 B.n974 163.367
R1813 B.n972 B.n150 163.367
R1814 B.n968 B.n966 163.367
R1815 B.n964 B.n152 163.367
R1816 B.n960 B.n958 163.367
R1817 B.n955 B.n954 163.367
R1818 B.n952 B.n158 163.367
R1819 B.n948 B.n946 163.367
R1820 B.n944 B.n160 163.367
R1821 B.n940 B.n938 163.367
R1822 B.n936 B.n162 163.367
R1823 B.n932 B.n930 163.367
R1824 B.n928 B.n164 163.367
R1825 B.n924 B.n922 163.367
R1826 B.n920 B.n166 163.367
R1827 B.n916 B.n914 163.367
R1828 B.n912 B.n168 163.367
R1829 B.n908 B.n906 163.367
R1830 B.n904 B.n170 163.367
R1831 B.n900 B.n898 163.367
R1832 B.n896 B.n172 163.367
R1833 B.n892 B.n890 163.367
R1834 B.n888 B.n174 163.367
R1835 B.n884 B.n882 163.367
R1836 B.n880 B.n176 163.367
R1837 B.n876 B.n874 163.367
R1838 B.n872 B.n178 163.367
R1839 B.n868 B.n866 163.367
R1840 B.n582 B.n307 163.367
R1841 B.n586 B.n307 163.367
R1842 B.n586 B.n301 163.367
R1843 B.n594 B.n301 163.367
R1844 B.n594 B.n299 163.367
R1845 B.n598 B.n299 163.367
R1846 B.n598 B.n293 163.367
R1847 B.n606 B.n293 163.367
R1848 B.n606 B.n291 163.367
R1849 B.n610 B.n291 163.367
R1850 B.n610 B.n285 163.367
R1851 B.n618 B.n285 163.367
R1852 B.n618 B.n283 163.367
R1853 B.n622 B.n283 163.367
R1854 B.n622 B.n277 163.367
R1855 B.n630 B.n277 163.367
R1856 B.n630 B.n275 163.367
R1857 B.n634 B.n275 163.367
R1858 B.n634 B.n268 163.367
R1859 B.n642 B.n268 163.367
R1860 B.n642 B.n266 163.367
R1861 B.n646 B.n266 163.367
R1862 B.n646 B.n261 163.367
R1863 B.n654 B.n261 163.367
R1864 B.n654 B.n259 163.367
R1865 B.n658 B.n259 163.367
R1866 B.n658 B.n253 163.367
R1867 B.n666 B.n253 163.367
R1868 B.n666 B.n251 163.367
R1869 B.n670 B.n251 163.367
R1870 B.n670 B.n245 163.367
R1871 B.n678 B.n245 163.367
R1872 B.n678 B.n243 163.367
R1873 B.n682 B.n243 163.367
R1874 B.n682 B.n237 163.367
R1875 B.n690 B.n237 163.367
R1876 B.n690 B.n235 163.367
R1877 B.n694 B.n235 163.367
R1878 B.n694 B.n229 163.367
R1879 B.n702 B.n229 163.367
R1880 B.n702 B.n227 163.367
R1881 B.n706 B.n227 163.367
R1882 B.n706 B.n221 163.367
R1883 B.n714 B.n221 163.367
R1884 B.n714 B.n219 163.367
R1885 B.n718 B.n219 163.367
R1886 B.n718 B.n213 163.367
R1887 B.n726 B.n213 163.367
R1888 B.n726 B.n211 163.367
R1889 B.n730 B.n211 163.367
R1890 B.n730 B.n205 163.367
R1891 B.n738 B.n205 163.367
R1892 B.n738 B.n203 163.367
R1893 B.n742 B.n203 163.367
R1894 B.n742 B.n197 163.367
R1895 B.n750 B.n197 163.367
R1896 B.n750 B.n195 163.367
R1897 B.n754 B.n195 163.367
R1898 B.n754 B.n189 163.367
R1899 B.n762 B.n189 163.367
R1900 B.n762 B.n187 163.367
R1901 B.n767 B.n187 163.367
R1902 B.n767 B.n181 163.367
R1903 B.n775 B.n181 163.367
R1904 B.n776 B.n775 163.367
R1905 B.n776 B.n5 163.367
R1906 B.n6 B.n5 163.367
R1907 B.n7 B.n6 163.367
R1908 B.n782 B.n7 163.367
R1909 B.n783 B.n782 163.367
R1910 B.n783 B.n13 163.367
R1911 B.n14 B.n13 163.367
R1912 B.n15 B.n14 163.367
R1913 B.n788 B.n15 163.367
R1914 B.n788 B.n20 163.367
R1915 B.n21 B.n20 163.367
R1916 B.n22 B.n21 163.367
R1917 B.n793 B.n22 163.367
R1918 B.n793 B.n27 163.367
R1919 B.n28 B.n27 163.367
R1920 B.n29 B.n28 163.367
R1921 B.n798 B.n29 163.367
R1922 B.n798 B.n34 163.367
R1923 B.n35 B.n34 163.367
R1924 B.n36 B.n35 163.367
R1925 B.n803 B.n36 163.367
R1926 B.n803 B.n41 163.367
R1927 B.n42 B.n41 163.367
R1928 B.n43 B.n42 163.367
R1929 B.n808 B.n43 163.367
R1930 B.n808 B.n48 163.367
R1931 B.n49 B.n48 163.367
R1932 B.n50 B.n49 163.367
R1933 B.n813 B.n50 163.367
R1934 B.n813 B.n55 163.367
R1935 B.n56 B.n55 163.367
R1936 B.n57 B.n56 163.367
R1937 B.n818 B.n57 163.367
R1938 B.n818 B.n62 163.367
R1939 B.n63 B.n62 163.367
R1940 B.n64 B.n63 163.367
R1941 B.n823 B.n64 163.367
R1942 B.n823 B.n69 163.367
R1943 B.n70 B.n69 163.367
R1944 B.n71 B.n70 163.367
R1945 B.n828 B.n71 163.367
R1946 B.n828 B.n76 163.367
R1947 B.n77 B.n76 163.367
R1948 B.n78 B.n77 163.367
R1949 B.n833 B.n78 163.367
R1950 B.n833 B.n83 163.367
R1951 B.n84 B.n83 163.367
R1952 B.n85 B.n84 163.367
R1953 B.n838 B.n85 163.367
R1954 B.n838 B.n90 163.367
R1955 B.n91 B.n90 163.367
R1956 B.n92 B.n91 163.367
R1957 B.n843 B.n92 163.367
R1958 B.n843 B.n97 163.367
R1959 B.n98 B.n97 163.367
R1960 B.n99 B.n98 163.367
R1961 B.n848 B.n99 163.367
R1962 B.n848 B.n104 163.367
R1963 B.n105 B.n104 163.367
R1964 B.n106 B.n105 163.367
R1965 B.n853 B.n106 163.367
R1966 B.n853 B.n111 163.367
R1967 B.n112 B.n111 163.367
R1968 B.n113 B.n112 163.367
R1969 B.n858 B.n113 163.367
R1970 B.n858 B.n118 163.367
R1971 B.n119 B.n118 163.367
R1972 B.n120 B.n119 163.367
R1973 B.n576 B.n574 163.367
R1974 B.n574 B.n573 163.367
R1975 B.n570 B.n569 163.367
R1976 B.n567 B.n315 163.367
R1977 B.n563 B.n561 163.367
R1978 B.n559 B.n317 163.367
R1979 B.n555 B.n553 163.367
R1980 B.n551 B.n319 163.367
R1981 B.n547 B.n545 163.367
R1982 B.n543 B.n321 163.367
R1983 B.n539 B.n537 163.367
R1984 B.n535 B.n323 163.367
R1985 B.n531 B.n529 163.367
R1986 B.n527 B.n325 163.367
R1987 B.n523 B.n521 163.367
R1988 B.n519 B.n327 163.367
R1989 B.n515 B.n513 163.367
R1990 B.n511 B.n329 163.367
R1991 B.n507 B.n505 163.367
R1992 B.n503 B.n331 163.367
R1993 B.n499 B.n497 163.367
R1994 B.n495 B.n333 163.367
R1995 B.n491 B.n489 163.367
R1996 B.n487 B.n335 163.367
R1997 B.n482 B.n480 163.367
R1998 B.n478 B.n339 163.367
R1999 B.n474 B.n472 163.367
R2000 B.n470 B.n341 163.367
R2001 B.n466 B.n464 163.367
R2002 B.n462 B.n343 163.367
R2003 B.n458 B.n456 163.367
R2004 B.n454 B.n348 163.367
R2005 B.n450 B.n448 163.367
R2006 B.n446 B.n350 163.367
R2007 B.n442 B.n440 163.367
R2008 B.n438 B.n352 163.367
R2009 B.n434 B.n432 163.367
R2010 B.n430 B.n354 163.367
R2011 B.n426 B.n424 163.367
R2012 B.n422 B.n356 163.367
R2013 B.n418 B.n416 163.367
R2014 B.n414 B.n358 163.367
R2015 B.n410 B.n408 163.367
R2016 B.n406 B.n360 163.367
R2017 B.n402 B.n400 163.367
R2018 B.n398 B.n362 163.367
R2019 B.n394 B.n392 163.367
R2020 B.n390 B.n364 163.367
R2021 B.n386 B.n384 163.367
R2022 B.n382 B.n366 163.367
R2023 B.n378 B.n376 163.367
R2024 B.n374 B.n368 163.367
R2025 B.n370 B.n309 163.367
R2026 B.n580 B.n305 163.367
R2027 B.n588 B.n305 163.367
R2028 B.n588 B.n303 163.367
R2029 B.n592 B.n303 163.367
R2030 B.n592 B.n297 163.367
R2031 B.n600 B.n297 163.367
R2032 B.n600 B.n295 163.367
R2033 B.n604 B.n295 163.367
R2034 B.n604 B.n289 163.367
R2035 B.n612 B.n289 163.367
R2036 B.n612 B.n287 163.367
R2037 B.n616 B.n287 163.367
R2038 B.n616 B.n281 163.367
R2039 B.n624 B.n281 163.367
R2040 B.n624 B.n279 163.367
R2041 B.n628 B.n279 163.367
R2042 B.n628 B.n273 163.367
R2043 B.n636 B.n273 163.367
R2044 B.n636 B.n271 163.367
R2045 B.n640 B.n271 163.367
R2046 B.n640 B.n265 163.367
R2047 B.n648 B.n265 163.367
R2048 B.n648 B.n263 163.367
R2049 B.n652 B.n263 163.367
R2050 B.n652 B.n257 163.367
R2051 B.n660 B.n257 163.367
R2052 B.n660 B.n255 163.367
R2053 B.n664 B.n255 163.367
R2054 B.n664 B.n249 163.367
R2055 B.n672 B.n249 163.367
R2056 B.n672 B.n247 163.367
R2057 B.n676 B.n247 163.367
R2058 B.n676 B.n241 163.367
R2059 B.n684 B.n241 163.367
R2060 B.n684 B.n239 163.367
R2061 B.n688 B.n239 163.367
R2062 B.n688 B.n233 163.367
R2063 B.n696 B.n233 163.367
R2064 B.n696 B.n231 163.367
R2065 B.n700 B.n231 163.367
R2066 B.n700 B.n225 163.367
R2067 B.n708 B.n225 163.367
R2068 B.n708 B.n223 163.367
R2069 B.n712 B.n223 163.367
R2070 B.n712 B.n217 163.367
R2071 B.n720 B.n217 163.367
R2072 B.n720 B.n215 163.367
R2073 B.n724 B.n215 163.367
R2074 B.n724 B.n209 163.367
R2075 B.n732 B.n209 163.367
R2076 B.n732 B.n207 163.367
R2077 B.n736 B.n207 163.367
R2078 B.n736 B.n201 163.367
R2079 B.n744 B.n201 163.367
R2080 B.n744 B.n199 163.367
R2081 B.n748 B.n199 163.367
R2082 B.n748 B.n193 163.367
R2083 B.n756 B.n193 163.367
R2084 B.n756 B.n191 163.367
R2085 B.n760 B.n191 163.367
R2086 B.n760 B.n185 163.367
R2087 B.n769 B.n185 163.367
R2088 B.n769 B.n183 163.367
R2089 B.n773 B.n183 163.367
R2090 B.n773 B.n3 163.367
R2091 B.n1210 B.n3 163.367
R2092 B.n1206 B.n2 163.367
R2093 B.n1206 B.n1205 163.367
R2094 B.n1205 B.n9 163.367
R2095 B.n1201 B.n9 163.367
R2096 B.n1201 B.n11 163.367
R2097 B.n1197 B.n11 163.367
R2098 B.n1197 B.n17 163.367
R2099 B.n1193 B.n17 163.367
R2100 B.n1193 B.n19 163.367
R2101 B.n1189 B.n19 163.367
R2102 B.n1189 B.n24 163.367
R2103 B.n1185 B.n24 163.367
R2104 B.n1185 B.n26 163.367
R2105 B.n1181 B.n26 163.367
R2106 B.n1181 B.n31 163.367
R2107 B.n1177 B.n31 163.367
R2108 B.n1177 B.n33 163.367
R2109 B.n1173 B.n33 163.367
R2110 B.n1173 B.n38 163.367
R2111 B.n1169 B.n38 163.367
R2112 B.n1169 B.n40 163.367
R2113 B.n1165 B.n40 163.367
R2114 B.n1165 B.n45 163.367
R2115 B.n1161 B.n45 163.367
R2116 B.n1161 B.n47 163.367
R2117 B.n1157 B.n47 163.367
R2118 B.n1157 B.n52 163.367
R2119 B.n1153 B.n52 163.367
R2120 B.n1153 B.n54 163.367
R2121 B.n1149 B.n54 163.367
R2122 B.n1149 B.n59 163.367
R2123 B.n1145 B.n59 163.367
R2124 B.n1145 B.n61 163.367
R2125 B.n1141 B.n61 163.367
R2126 B.n1141 B.n66 163.367
R2127 B.n1137 B.n66 163.367
R2128 B.n1137 B.n68 163.367
R2129 B.n1133 B.n68 163.367
R2130 B.n1133 B.n73 163.367
R2131 B.n1129 B.n73 163.367
R2132 B.n1129 B.n75 163.367
R2133 B.n1125 B.n75 163.367
R2134 B.n1125 B.n80 163.367
R2135 B.n1121 B.n80 163.367
R2136 B.n1121 B.n82 163.367
R2137 B.n1117 B.n82 163.367
R2138 B.n1117 B.n87 163.367
R2139 B.n1113 B.n87 163.367
R2140 B.n1113 B.n89 163.367
R2141 B.n1109 B.n89 163.367
R2142 B.n1109 B.n94 163.367
R2143 B.n1105 B.n94 163.367
R2144 B.n1105 B.n96 163.367
R2145 B.n1101 B.n96 163.367
R2146 B.n1101 B.n101 163.367
R2147 B.n1097 B.n101 163.367
R2148 B.n1097 B.n103 163.367
R2149 B.n1093 B.n103 163.367
R2150 B.n1093 B.n108 163.367
R2151 B.n1089 B.n108 163.367
R2152 B.n1089 B.n110 163.367
R2153 B.n1085 B.n110 163.367
R2154 B.n1085 B.n115 163.367
R2155 B.n1081 B.n115 163.367
R2156 B.n1081 B.n117 163.367
R2157 B.n1077 B.n117 163.367
R2158 B.n1072 B.n122 71.676
R2159 B.n1071 B.n1070 71.676
R2160 B.n1064 B.n124 71.676
R2161 B.n1063 B.n1062 71.676
R2162 B.n1056 B.n126 71.676
R2163 B.n1055 B.n1054 71.676
R2164 B.n1048 B.n128 71.676
R2165 B.n1047 B.n1046 71.676
R2166 B.n1040 B.n130 71.676
R2167 B.n1039 B.n1038 71.676
R2168 B.n1032 B.n132 71.676
R2169 B.n1031 B.n1030 71.676
R2170 B.n1024 B.n134 71.676
R2171 B.n1023 B.n1022 71.676
R2172 B.n1016 B.n136 71.676
R2173 B.n1015 B.n1014 71.676
R2174 B.n1008 B.n138 71.676
R2175 B.n1007 B.n1006 71.676
R2176 B.n1000 B.n140 71.676
R2177 B.n999 B.n998 71.676
R2178 B.n992 B.n142 71.676
R2179 B.n991 B.n990 71.676
R2180 B.n984 B.n144 71.676
R2181 B.n983 B.n982 71.676
R2182 B.n975 B.n146 71.676
R2183 B.n974 B.n973 71.676
R2184 B.n967 B.n150 71.676
R2185 B.n966 B.n965 71.676
R2186 B.n959 B.n152 71.676
R2187 B.n958 B.n156 71.676
R2188 B.n954 B.n953 71.676
R2189 B.n947 B.n158 71.676
R2190 B.n946 B.n945 71.676
R2191 B.n939 B.n160 71.676
R2192 B.n938 B.n937 71.676
R2193 B.n931 B.n162 71.676
R2194 B.n930 B.n929 71.676
R2195 B.n923 B.n164 71.676
R2196 B.n922 B.n921 71.676
R2197 B.n915 B.n166 71.676
R2198 B.n914 B.n913 71.676
R2199 B.n907 B.n168 71.676
R2200 B.n906 B.n905 71.676
R2201 B.n899 B.n170 71.676
R2202 B.n898 B.n897 71.676
R2203 B.n891 B.n172 71.676
R2204 B.n890 B.n889 71.676
R2205 B.n883 B.n174 71.676
R2206 B.n882 B.n881 71.676
R2207 B.n875 B.n176 71.676
R2208 B.n874 B.n873 71.676
R2209 B.n867 B.n178 71.676
R2210 B.n866 B.n865 71.676
R2211 B.n865 B.n864 71.676
R2212 B.n868 B.n867 71.676
R2213 B.n873 B.n872 71.676
R2214 B.n876 B.n875 71.676
R2215 B.n881 B.n880 71.676
R2216 B.n884 B.n883 71.676
R2217 B.n889 B.n888 71.676
R2218 B.n892 B.n891 71.676
R2219 B.n897 B.n896 71.676
R2220 B.n900 B.n899 71.676
R2221 B.n905 B.n904 71.676
R2222 B.n908 B.n907 71.676
R2223 B.n913 B.n912 71.676
R2224 B.n916 B.n915 71.676
R2225 B.n921 B.n920 71.676
R2226 B.n924 B.n923 71.676
R2227 B.n929 B.n928 71.676
R2228 B.n932 B.n931 71.676
R2229 B.n937 B.n936 71.676
R2230 B.n940 B.n939 71.676
R2231 B.n945 B.n944 71.676
R2232 B.n948 B.n947 71.676
R2233 B.n953 B.n952 71.676
R2234 B.n955 B.n156 71.676
R2235 B.n960 B.n959 71.676
R2236 B.n965 B.n964 71.676
R2237 B.n968 B.n967 71.676
R2238 B.n973 B.n972 71.676
R2239 B.n976 B.n975 71.676
R2240 B.n982 B.n981 71.676
R2241 B.n985 B.n984 71.676
R2242 B.n990 B.n989 71.676
R2243 B.n993 B.n992 71.676
R2244 B.n998 B.n997 71.676
R2245 B.n1001 B.n1000 71.676
R2246 B.n1006 B.n1005 71.676
R2247 B.n1009 B.n1008 71.676
R2248 B.n1014 B.n1013 71.676
R2249 B.n1017 B.n1016 71.676
R2250 B.n1022 B.n1021 71.676
R2251 B.n1025 B.n1024 71.676
R2252 B.n1030 B.n1029 71.676
R2253 B.n1033 B.n1032 71.676
R2254 B.n1038 B.n1037 71.676
R2255 B.n1041 B.n1040 71.676
R2256 B.n1046 B.n1045 71.676
R2257 B.n1049 B.n1048 71.676
R2258 B.n1054 B.n1053 71.676
R2259 B.n1057 B.n1056 71.676
R2260 B.n1062 B.n1061 71.676
R2261 B.n1065 B.n1064 71.676
R2262 B.n1070 B.n1069 71.676
R2263 B.n1073 B.n1072 71.676
R2264 B.n575 B.n311 71.676
R2265 B.n573 B.n313 71.676
R2266 B.n569 B.n568 71.676
R2267 B.n562 B.n315 71.676
R2268 B.n561 B.n560 71.676
R2269 B.n554 B.n317 71.676
R2270 B.n553 B.n552 71.676
R2271 B.n546 B.n319 71.676
R2272 B.n545 B.n544 71.676
R2273 B.n538 B.n321 71.676
R2274 B.n537 B.n536 71.676
R2275 B.n530 B.n323 71.676
R2276 B.n529 B.n528 71.676
R2277 B.n522 B.n325 71.676
R2278 B.n521 B.n520 71.676
R2279 B.n514 B.n327 71.676
R2280 B.n513 B.n512 71.676
R2281 B.n506 B.n329 71.676
R2282 B.n505 B.n504 71.676
R2283 B.n498 B.n331 71.676
R2284 B.n497 B.n496 71.676
R2285 B.n490 B.n333 71.676
R2286 B.n489 B.n488 71.676
R2287 B.n481 B.n335 71.676
R2288 B.n480 B.n479 71.676
R2289 B.n473 B.n339 71.676
R2290 B.n472 B.n471 71.676
R2291 B.n465 B.n341 71.676
R2292 B.n464 B.n463 71.676
R2293 B.n457 B.n343 71.676
R2294 B.n456 B.n455 71.676
R2295 B.n449 B.n348 71.676
R2296 B.n448 B.n447 71.676
R2297 B.n441 B.n350 71.676
R2298 B.n440 B.n439 71.676
R2299 B.n433 B.n352 71.676
R2300 B.n432 B.n431 71.676
R2301 B.n425 B.n354 71.676
R2302 B.n424 B.n423 71.676
R2303 B.n417 B.n356 71.676
R2304 B.n416 B.n415 71.676
R2305 B.n409 B.n358 71.676
R2306 B.n408 B.n407 71.676
R2307 B.n401 B.n360 71.676
R2308 B.n400 B.n399 71.676
R2309 B.n393 B.n362 71.676
R2310 B.n392 B.n391 71.676
R2311 B.n385 B.n364 71.676
R2312 B.n384 B.n383 71.676
R2313 B.n377 B.n366 71.676
R2314 B.n376 B.n375 71.676
R2315 B.n369 B.n368 71.676
R2316 B.n576 B.n575 71.676
R2317 B.n570 B.n313 71.676
R2318 B.n568 B.n567 71.676
R2319 B.n563 B.n562 71.676
R2320 B.n560 B.n559 71.676
R2321 B.n555 B.n554 71.676
R2322 B.n552 B.n551 71.676
R2323 B.n547 B.n546 71.676
R2324 B.n544 B.n543 71.676
R2325 B.n539 B.n538 71.676
R2326 B.n536 B.n535 71.676
R2327 B.n531 B.n530 71.676
R2328 B.n528 B.n527 71.676
R2329 B.n523 B.n522 71.676
R2330 B.n520 B.n519 71.676
R2331 B.n515 B.n514 71.676
R2332 B.n512 B.n511 71.676
R2333 B.n507 B.n506 71.676
R2334 B.n504 B.n503 71.676
R2335 B.n499 B.n498 71.676
R2336 B.n496 B.n495 71.676
R2337 B.n491 B.n490 71.676
R2338 B.n488 B.n487 71.676
R2339 B.n482 B.n481 71.676
R2340 B.n479 B.n478 71.676
R2341 B.n474 B.n473 71.676
R2342 B.n471 B.n470 71.676
R2343 B.n466 B.n465 71.676
R2344 B.n463 B.n462 71.676
R2345 B.n458 B.n457 71.676
R2346 B.n455 B.n454 71.676
R2347 B.n450 B.n449 71.676
R2348 B.n447 B.n446 71.676
R2349 B.n442 B.n441 71.676
R2350 B.n439 B.n438 71.676
R2351 B.n434 B.n433 71.676
R2352 B.n431 B.n430 71.676
R2353 B.n426 B.n425 71.676
R2354 B.n423 B.n422 71.676
R2355 B.n418 B.n417 71.676
R2356 B.n415 B.n414 71.676
R2357 B.n410 B.n409 71.676
R2358 B.n407 B.n406 71.676
R2359 B.n402 B.n401 71.676
R2360 B.n399 B.n398 71.676
R2361 B.n394 B.n393 71.676
R2362 B.n391 B.n390 71.676
R2363 B.n386 B.n385 71.676
R2364 B.n383 B.n382 71.676
R2365 B.n378 B.n377 71.676
R2366 B.n375 B.n374 71.676
R2367 B.n370 B.n369 71.676
R2368 B.n1211 B.n1210 71.676
R2369 B.n1211 B.n2 71.676
R2370 B.n148 B.n147 64.0005
R2371 B.n154 B.n153 64.0005
R2372 B.n345 B.n344 64.0005
R2373 B.n337 B.n336 64.0005
R2374 B.n581 B.n310 63.7932
R2375 B.n1078 B.n121 63.7932
R2376 B.n979 B.n148 59.5399
R2377 B.n155 B.n154 59.5399
R2378 B.n346 B.n345 59.5399
R2379 B.n484 B.n337 59.5399
R2380 B.n581 B.n306 38.389
R2381 B.n587 B.n306 38.389
R2382 B.n587 B.n302 38.389
R2383 B.n593 B.n302 38.389
R2384 B.n593 B.n298 38.389
R2385 B.n599 B.n298 38.389
R2386 B.n599 B.n294 38.389
R2387 B.n605 B.n294 38.389
R2388 B.n611 B.n290 38.389
R2389 B.n611 B.n286 38.389
R2390 B.n617 B.n286 38.389
R2391 B.n617 B.n282 38.389
R2392 B.n623 B.n282 38.389
R2393 B.n623 B.n278 38.389
R2394 B.n629 B.n278 38.389
R2395 B.n629 B.n274 38.389
R2396 B.n635 B.n274 38.389
R2397 B.n635 B.n269 38.389
R2398 B.n641 B.n269 38.389
R2399 B.n641 B.n270 38.389
R2400 B.n647 B.n262 38.389
R2401 B.n653 B.n262 38.389
R2402 B.n653 B.n258 38.389
R2403 B.n659 B.n258 38.389
R2404 B.n659 B.n254 38.389
R2405 B.n665 B.n254 38.389
R2406 B.n665 B.n250 38.389
R2407 B.n671 B.n250 38.389
R2408 B.n677 B.n246 38.389
R2409 B.n677 B.n242 38.389
R2410 B.n683 B.n242 38.389
R2411 B.n683 B.n238 38.389
R2412 B.n689 B.n238 38.389
R2413 B.n689 B.n234 38.389
R2414 B.n695 B.n234 38.389
R2415 B.n695 B.n230 38.389
R2416 B.n701 B.n230 38.389
R2417 B.n707 B.n226 38.389
R2418 B.n707 B.n222 38.389
R2419 B.n713 B.n222 38.389
R2420 B.n713 B.n218 38.389
R2421 B.n719 B.n218 38.389
R2422 B.n719 B.n214 38.389
R2423 B.n725 B.n214 38.389
R2424 B.n725 B.n210 38.389
R2425 B.n731 B.n210 38.389
R2426 B.n737 B.n206 38.389
R2427 B.n737 B.n202 38.389
R2428 B.n743 B.n202 38.389
R2429 B.n743 B.n198 38.389
R2430 B.n749 B.n198 38.389
R2431 B.n749 B.n194 38.389
R2432 B.n755 B.n194 38.389
R2433 B.n755 B.n190 38.389
R2434 B.n761 B.n190 38.389
R2435 B.n768 B.n186 38.389
R2436 B.n768 B.n182 38.389
R2437 B.n774 B.n182 38.389
R2438 B.n774 B.n4 38.389
R2439 B.n1209 B.n4 38.389
R2440 B.n1209 B.n1208 38.389
R2441 B.n1208 B.n1207 38.389
R2442 B.n1207 B.n8 38.389
R2443 B.n12 B.n8 38.389
R2444 B.n1200 B.n12 38.389
R2445 B.n1200 B.n1199 38.389
R2446 B.n1198 B.n16 38.389
R2447 B.n1192 B.n16 38.389
R2448 B.n1192 B.n1191 38.389
R2449 B.n1191 B.n1190 38.389
R2450 B.n1190 B.n23 38.389
R2451 B.n1184 B.n23 38.389
R2452 B.n1184 B.n1183 38.389
R2453 B.n1183 B.n1182 38.389
R2454 B.n1182 B.n30 38.389
R2455 B.n1176 B.n1175 38.389
R2456 B.n1175 B.n1174 38.389
R2457 B.n1174 B.n37 38.389
R2458 B.n1168 B.n37 38.389
R2459 B.n1168 B.n1167 38.389
R2460 B.n1167 B.n1166 38.389
R2461 B.n1166 B.n44 38.389
R2462 B.n1160 B.n44 38.389
R2463 B.n1160 B.n1159 38.389
R2464 B.n1158 B.n51 38.389
R2465 B.n1152 B.n51 38.389
R2466 B.n1152 B.n1151 38.389
R2467 B.n1151 B.n1150 38.389
R2468 B.n1150 B.n58 38.389
R2469 B.n1144 B.n58 38.389
R2470 B.n1144 B.n1143 38.389
R2471 B.n1143 B.n1142 38.389
R2472 B.n1142 B.n65 38.389
R2473 B.n1136 B.n1135 38.389
R2474 B.n1135 B.n1134 38.389
R2475 B.n1134 B.n72 38.389
R2476 B.n1128 B.n72 38.389
R2477 B.n1128 B.n1127 38.389
R2478 B.n1127 B.n1126 38.389
R2479 B.n1126 B.n79 38.389
R2480 B.n1120 B.n79 38.389
R2481 B.n1119 B.n1118 38.389
R2482 B.n1118 B.n86 38.389
R2483 B.n1112 B.n86 38.389
R2484 B.n1112 B.n1111 38.389
R2485 B.n1111 B.n1110 38.389
R2486 B.n1110 B.n93 38.389
R2487 B.n1104 B.n93 38.389
R2488 B.n1104 B.n1103 38.389
R2489 B.n1103 B.n1102 38.389
R2490 B.n1102 B.n100 38.389
R2491 B.n1096 B.n100 38.389
R2492 B.n1096 B.n1095 38.389
R2493 B.n1094 B.n107 38.389
R2494 B.n1088 B.n107 38.389
R2495 B.n1088 B.n1087 38.389
R2496 B.n1087 B.n1086 38.389
R2497 B.n1086 B.n114 38.389
R2498 B.n1080 B.n114 38.389
R2499 B.n1080 B.n1079 38.389
R2500 B.n1079 B.n1078 38.389
R2501 B.t7 B.n186 36.6954
R2502 B.n1199 B.t4 36.6954
R2503 B.n671 B.t5 35.5663
R2504 B.n1136 B.t3 35.5663
R2505 B.n647 B.t8 29.921
R2506 B.n1120 B.t9 29.921
R2507 B.n579 B.n578 29.8151
R2508 B.n583 B.n308 29.8151
R2509 B.n863 B.n862 29.8151
R2510 B.n1076 B.n1075 29.8151
R2511 B.t11 B.n290 26.5337
R2512 B.n1095 B.t15 26.5337
R2513 B.t1 B.n206 25.4047
R2514 B.t6 B.n30 25.4047
R2515 B.n701 B.t0 24.2756
R2516 B.t2 B.n1158 24.2756
R2517 B B.n1212 18.0485
R2518 B.t0 B.n226 14.1139
R2519 B.n1159 B.t2 14.1139
R2520 B.n731 B.t1 12.9848
R2521 B.n1176 B.t6 12.9848
R2522 B.n605 B.t11 11.8558
R2523 B.t15 B.n1094 11.8558
R2524 B.n579 B.n304 10.6151
R2525 B.n589 B.n304 10.6151
R2526 B.n590 B.n589 10.6151
R2527 B.n591 B.n590 10.6151
R2528 B.n591 B.n296 10.6151
R2529 B.n601 B.n296 10.6151
R2530 B.n602 B.n601 10.6151
R2531 B.n603 B.n602 10.6151
R2532 B.n603 B.n288 10.6151
R2533 B.n613 B.n288 10.6151
R2534 B.n614 B.n613 10.6151
R2535 B.n615 B.n614 10.6151
R2536 B.n615 B.n280 10.6151
R2537 B.n625 B.n280 10.6151
R2538 B.n626 B.n625 10.6151
R2539 B.n627 B.n626 10.6151
R2540 B.n627 B.n272 10.6151
R2541 B.n637 B.n272 10.6151
R2542 B.n638 B.n637 10.6151
R2543 B.n639 B.n638 10.6151
R2544 B.n639 B.n264 10.6151
R2545 B.n649 B.n264 10.6151
R2546 B.n650 B.n649 10.6151
R2547 B.n651 B.n650 10.6151
R2548 B.n651 B.n256 10.6151
R2549 B.n661 B.n256 10.6151
R2550 B.n662 B.n661 10.6151
R2551 B.n663 B.n662 10.6151
R2552 B.n663 B.n248 10.6151
R2553 B.n673 B.n248 10.6151
R2554 B.n674 B.n673 10.6151
R2555 B.n675 B.n674 10.6151
R2556 B.n675 B.n240 10.6151
R2557 B.n685 B.n240 10.6151
R2558 B.n686 B.n685 10.6151
R2559 B.n687 B.n686 10.6151
R2560 B.n687 B.n232 10.6151
R2561 B.n697 B.n232 10.6151
R2562 B.n698 B.n697 10.6151
R2563 B.n699 B.n698 10.6151
R2564 B.n699 B.n224 10.6151
R2565 B.n709 B.n224 10.6151
R2566 B.n710 B.n709 10.6151
R2567 B.n711 B.n710 10.6151
R2568 B.n711 B.n216 10.6151
R2569 B.n721 B.n216 10.6151
R2570 B.n722 B.n721 10.6151
R2571 B.n723 B.n722 10.6151
R2572 B.n723 B.n208 10.6151
R2573 B.n733 B.n208 10.6151
R2574 B.n734 B.n733 10.6151
R2575 B.n735 B.n734 10.6151
R2576 B.n735 B.n200 10.6151
R2577 B.n745 B.n200 10.6151
R2578 B.n746 B.n745 10.6151
R2579 B.n747 B.n746 10.6151
R2580 B.n747 B.n192 10.6151
R2581 B.n757 B.n192 10.6151
R2582 B.n758 B.n757 10.6151
R2583 B.n759 B.n758 10.6151
R2584 B.n759 B.n184 10.6151
R2585 B.n770 B.n184 10.6151
R2586 B.n771 B.n770 10.6151
R2587 B.n772 B.n771 10.6151
R2588 B.n772 B.n0 10.6151
R2589 B.n578 B.n577 10.6151
R2590 B.n577 B.n312 10.6151
R2591 B.n572 B.n312 10.6151
R2592 B.n572 B.n571 10.6151
R2593 B.n571 B.n314 10.6151
R2594 B.n566 B.n314 10.6151
R2595 B.n566 B.n565 10.6151
R2596 B.n565 B.n564 10.6151
R2597 B.n564 B.n316 10.6151
R2598 B.n558 B.n316 10.6151
R2599 B.n558 B.n557 10.6151
R2600 B.n557 B.n556 10.6151
R2601 B.n556 B.n318 10.6151
R2602 B.n550 B.n318 10.6151
R2603 B.n550 B.n549 10.6151
R2604 B.n549 B.n548 10.6151
R2605 B.n548 B.n320 10.6151
R2606 B.n542 B.n320 10.6151
R2607 B.n542 B.n541 10.6151
R2608 B.n541 B.n540 10.6151
R2609 B.n540 B.n322 10.6151
R2610 B.n534 B.n322 10.6151
R2611 B.n534 B.n533 10.6151
R2612 B.n533 B.n532 10.6151
R2613 B.n532 B.n324 10.6151
R2614 B.n526 B.n324 10.6151
R2615 B.n526 B.n525 10.6151
R2616 B.n525 B.n524 10.6151
R2617 B.n524 B.n326 10.6151
R2618 B.n518 B.n326 10.6151
R2619 B.n518 B.n517 10.6151
R2620 B.n517 B.n516 10.6151
R2621 B.n516 B.n328 10.6151
R2622 B.n510 B.n328 10.6151
R2623 B.n510 B.n509 10.6151
R2624 B.n509 B.n508 10.6151
R2625 B.n508 B.n330 10.6151
R2626 B.n502 B.n330 10.6151
R2627 B.n502 B.n501 10.6151
R2628 B.n501 B.n500 10.6151
R2629 B.n500 B.n332 10.6151
R2630 B.n494 B.n332 10.6151
R2631 B.n494 B.n493 10.6151
R2632 B.n493 B.n492 10.6151
R2633 B.n492 B.n334 10.6151
R2634 B.n486 B.n334 10.6151
R2635 B.n486 B.n485 10.6151
R2636 B.n483 B.n338 10.6151
R2637 B.n477 B.n338 10.6151
R2638 B.n477 B.n476 10.6151
R2639 B.n476 B.n475 10.6151
R2640 B.n475 B.n340 10.6151
R2641 B.n469 B.n340 10.6151
R2642 B.n469 B.n468 10.6151
R2643 B.n468 B.n467 10.6151
R2644 B.n467 B.n342 10.6151
R2645 B.n461 B.n460 10.6151
R2646 B.n460 B.n459 10.6151
R2647 B.n459 B.n347 10.6151
R2648 B.n453 B.n347 10.6151
R2649 B.n453 B.n452 10.6151
R2650 B.n452 B.n451 10.6151
R2651 B.n451 B.n349 10.6151
R2652 B.n445 B.n349 10.6151
R2653 B.n445 B.n444 10.6151
R2654 B.n444 B.n443 10.6151
R2655 B.n443 B.n351 10.6151
R2656 B.n437 B.n351 10.6151
R2657 B.n437 B.n436 10.6151
R2658 B.n436 B.n435 10.6151
R2659 B.n435 B.n353 10.6151
R2660 B.n429 B.n353 10.6151
R2661 B.n429 B.n428 10.6151
R2662 B.n428 B.n427 10.6151
R2663 B.n427 B.n355 10.6151
R2664 B.n421 B.n355 10.6151
R2665 B.n421 B.n420 10.6151
R2666 B.n420 B.n419 10.6151
R2667 B.n419 B.n357 10.6151
R2668 B.n413 B.n357 10.6151
R2669 B.n413 B.n412 10.6151
R2670 B.n412 B.n411 10.6151
R2671 B.n411 B.n359 10.6151
R2672 B.n405 B.n359 10.6151
R2673 B.n405 B.n404 10.6151
R2674 B.n404 B.n403 10.6151
R2675 B.n403 B.n361 10.6151
R2676 B.n397 B.n361 10.6151
R2677 B.n397 B.n396 10.6151
R2678 B.n396 B.n395 10.6151
R2679 B.n395 B.n363 10.6151
R2680 B.n389 B.n363 10.6151
R2681 B.n389 B.n388 10.6151
R2682 B.n388 B.n387 10.6151
R2683 B.n387 B.n365 10.6151
R2684 B.n381 B.n365 10.6151
R2685 B.n381 B.n380 10.6151
R2686 B.n380 B.n379 10.6151
R2687 B.n379 B.n367 10.6151
R2688 B.n373 B.n367 10.6151
R2689 B.n373 B.n372 10.6151
R2690 B.n372 B.n371 10.6151
R2691 B.n371 B.n308 10.6151
R2692 B.n584 B.n583 10.6151
R2693 B.n585 B.n584 10.6151
R2694 B.n585 B.n300 10.6151
R2695 B.n595 B.n300 10.6151
R2696 B.n596 B.n595 10.6151
R2697 B.n597 B.n596 10.6151
R2698 B.n597 B.n292 10.6151
R2699 B.n607 B.n292 10.6151
R2700 B.n608 B.n607 10.6151
R2701 B.n609 B.n608 10.6151
R2702 B.n609 B.n284 10.6151
R2703 B.n619 B.n284 10.6151
R2704 B.n620 B.n619 10.6151
R2705 B.n621 B.n620 10.6151
R2706 B.n621 B.n276 10.6151
R2707 B.n631 B.n276 10.6151
R2708 B.n632 B.n631 10.6151
R2709 B.n633 B.n632 10.6151
R2710 B.n633 B.n267 10.6151
R2711 B.n643 B.n267 10.6151
R2712 B.n644 B.n643 10.6151
R2713 B.n645 B.n644 10.6151
R2714 B.n645 B.n260 10.6151
R2715 B.n655 B.n260 10.6151
R2716 B.n656 B.n655 10.6151
R2717 B.n657 B.n656 10.6151
R2718 B.n657 B.n252 10.6151
R2719 B.n667 B.n252 10.6151
R2720 B.n668 B.n667 10.6151
R2721 B.n669 B.n668 10.6151
R2722 B.n669 B.n244 10.6151
R2723 B.n679 B.n244 10.6151
R2724 B.n680 B.n679 10.6151
R2725 B.n681 B.n680 10.6151
R2726 B.n681 B.n236 10.6151
R2727 B.n691 B.n236 10.6151
R2728 B.n692 B.n691 10.6151
R2729 B.n693 B.n692 10.6151
R2730 B.n693 B.n228 10.6151
R2731 B.n703 B.n228 10.6151
R2732 B.n704 B.n703 10.6151
R2733 B.n705 B.n704 10.6151
R2734 B.n705 B.n220 10.6151
R2735 B.n715 B.n220 10.6151
R2736 B.n716 B.n715 10.6151
R2737 B.n717 B.n716 10.6151
R2738 B.n717 B.n212 10.6151
R2739 B.n727 B.n212 10.6151
R2740 B.n728 B.n727 10.6151
R2741 B.n729 B.n728 10.6151
R2742 B.n729 B.n204 10.6151
R2743 B.n739 B.n204 10.6151
R2744 B.n740 B.n739 10.6151
R2745 B.n741 B.n740 10.6151
R2746 B.n741 B.n196 10.6151
R2747 B.n751 B.n196 10.6151
R2748 B.n752 B.n751 10.6151
R2749 B.n753 B.n752 10.6151
R2750 B.n753 B.n188 10.6151
R2751 B.n763 B.n188 10.6151
R2752 B.n764 B.n763 10.6151
R2753 B.n766 B.n764 10.6151
R2754 B.n766 B.n765 10.6151
R2755 B.n765 B.n180 10.6151
R2756 B.n777 B.n180 10.6151
R2757 B.n778 B.n777 10.6151
R2758 B.n779 B.n778 10.6151
R2759 B.n780 B.n779 10.6151
R2760 B.n781 B.n780 10.6151
R2761 B.n784 B.n781 10.6151
R2762 B.n785 B.n784 10.6151
R2763 B.n786 B.n785 10.6151
R2764 B.n787 B.n786 10.6151
R2765 B.n789 B.n787 10.6151
R2766 B.n790 B.n789 10.6151
R2767 B.n791 B.n790 10.6151
R2768 B.n792 B.n791 10.6151
R2769 B.n794 B.n792 10.6151
R2770 B.n795 B.n794 10.6151
R2771 B.n796 B.n795 10.6151
R2772 B.n797 B.n796 10.6151
R2773 B.n799 B.n797 10.6151
R2774 B.n800 B.n799 10.6151
R2775 B.n801 B.n800 10.6151
R2776 B.n802 B.n801 10.6151
R2777 B.n804 B.n802 10.6151
R2778 B.n805 B.n804 10.6151
R2779 B.n806 B.n805 10.6151
R2780 B.n807 B.n806 10.6151
R2781 B.n809 B.n807 10.6151
R2782 B.n810 B.n809 10.6151
R2783 B.n811 B.n810 10.6151
R2784 B.n812 B.n811 10.6151
R2785 B.n814 B.n812 10.6151
R2786 B.n815 B.n814 10.6151
R2787 B.n816 B.n815 10.6151
R2788 B.n817 B.n816 10.6151
R2789 B.n819 B.n817 10.6151
R2790 B.n820 B.n819 10.6151
R2791 B.n821 B.n820 10.6151
R2792 B.n822 B.n821 10.6151
R2793 B.n824 B.n822 10.6151
R2794 B.n825 B.n824 10.6151
R2795 B.n826 B.n825 10.6151
R2796 B.n827 B.n826 10.6151
R2797 B.n829 B.n827 10.6151
R2798 B.n830 B.n829 10.6151
R2799 B.n831 B.n830 10.6151
R2800 B.n832 B.n831 10.6151
R2801 B.n834 B.n832 10.6151
R2802 B.n835 B.n834 10.6151
R2803 B.n836 B.n835 10.6151
R2804 B.n837 B.n836 10.6151
R2805 B.n839 B.n837 10.6151
R2806 B.n840 B.n839 10.6151
R2807 B.n841 B.n840 10.6151
R2808 B.n842 B.n841 10.6151
R2809 B.n844 B.n842 10.6151
R2810 B.n845 B.n844 10.6151
R2811 B.n846 B.n845 10.6151
R2812 B.n847 B.n846 10.6151
R2813 B.n849 B.n847 10.6151
R2814 B.n850 B.n849 10.6151
R2815 B.n851 B.n850 10.6151
R2816 B.n852 B.n851 10.6151
R2817 B.n854 B.n852 10.6151
R2818 B.n855 B.n854 10.6151
R2819 B.n856 B.n855 10.6151
R2820 B.n857 B.n856 10.6151
R2821 B.n859 B.n857 10.6151
R2822 B.n860 B.n859 10.6151
R2823 B.n861 B.n860 10.6151
R2824 B.n862 B.n861 10.6151
R2825 B.n1204 B.n1 10.6151
R2826 B.n1204 B.n1203 10.6151
R2827 B.n1203 B.n1202 10.6151
R2828 B.n1202 B.n10 10.6151
R2829 B.n1196 B.n10 10.6151
R2830 B.n1196 B.n1195 10.6151
R2831 B.n1195 B.n1194 10.6151
R2832 B.n1194 B.n18 10.6151
R2833 B.n1188 B.n18 10.6151
R2834 B.n1188 B.n1187 10.6151
R2835 B.n1187 B.n1186 10.6151
R2836 B.n1186 B.n25 10.6151
R2837 B.n1180 B.n25 10.6151
R2838 B.n1180 B.n1179 10.6151
R2839 B.n1179 B.n1178 10.6151
R2840 B.n1178 B.n32 10.6151
R2841 B.n1172 B.n32 10.6151
R2842 B.n1172 B.n1171 10.6151
R2843 B.n1171 B.n1170 10.6151
R2844 B.n1170 B.n39 10.6151
R2845 B.n1164 B.n39 10.6151
R2846 B.n1164 B.n1163 10.6151
R2847 B.n1163 B.n1162 10.6151
R2848 B.n1162 B.n46 10.6151
R2849 B.n1156 B.n46 10.6151
R2850 B.n1156 B.n1155 10.6151
R2851 B.n1155 B.n1154 10.6151
R2852 B.n1154 B.n53 10.6151
R2853 B.n1148 B.n53 10.6151
R2854 B.n1148 B.n1147 10.6151
R2855 B.n1147 B.n1146 10.6151
R2856 B.n1146 B.n60 10.6151
R2857 B.n1140 B.n60 10.6151
R2858 B.n1140 B.n1139 10.6151
R2859 B.n1139 B.n1138 10.6151
R2860 B.n1138 B.n67 10.6151
R2861 B.n1132 B.n67 10.6151
R2862 B.n1132 B.n1131 10.6151
R2863 B.n1131 B.n1130 10.6151
R2864 B.n1130 B.n74 10.6151
R2865 B.n1124 B.n74 10.6151
R2866 B.n1124 B.n1123 10.6151
R2867 B.n1123 B.n1122 10.6151
R2868 B.n1122 B.n81 10.6151
R2869 B.n1116 B.n81 10.6151
R2870 B.n1116 B.n1115 10.6151
R2871 B.n1115 B.n1114 10.6151
R2872 B.n1114 B.n88 10.6151
R2873 B.n1108 B.n88 10.6151
R2874 B.n1108 B.n1107 10.6151
R2875 B.n1107 B.n1106 10.6151
R2876 B.n1106 B.n95 10.6151
R2877 B.n1100 B.n95 10.6151
R2878 B.n1100 B.n1099 10.6151
R2879 B.n1099 B.n1098 10.6151
R2880 B.n1098 B.n102 10.6151
R2881 B.n1092 B.n102 10.6151
R2882 B.n1092 B.n1091 10.6151
R2883 B.n1091 B.n1090 10.6151
R2884 B.n1090 B.n109 10.6151
R2885 B.n1084 B.n109 10.6151
R2886 B.n1084 B.n1083 10.6151
R2887 B.n1083 B.n1082 10.6151
R2888 B.n1082 B.n116 10.6151
R2889 B.n1076 B.n116 10.6151
R2890 B.n1075 B.n1074 10.6151
R2891 B.n1074 B.n123 10.6151
R2892 B.n1068 B.n123 10.6151
R2893 B.n1068 B.n1067 10.6151
R2894 B.n1067 B.n1066 10.6151
R2895 B.n1066 B.n125 10.6151
R2896 B.n1060 B.n125 10.6151
R2897 B.n1060 B.n1059 10.6151
R2898 B.n1059 B.n1058 10.6151
R2899 B.n1058 B.n127 10.6151
R2900 B.n1052 B.n127 10.6151
R2901 B.n1052 B.n1051 10.6151
R2902 B.n1051 B.n1050 10.6151
R2903 B.n1050 B.n129 10.6151
R2904 B.n1044 B.n129 10.6151
R2905 B.n1044 B.n1043 10.6151
R2906 B.n1043 B.n1042 10.6151
R2907 B.n1042 B.n131 10.6151
R2908 B.n1036 B.n131 10.6151
R2909 B.n1036 B.n1035 10.6151
R2910 B.n1035 B.n1034 10.6151
R2911 B.n1034 B.n133 10.6151
R2912 B.n1028 B.n133 10.6151
R2913 B.n1028 B.n1027 10.6151
R2914 B.n1027 B.n1026 10.6151
R2915 B.n1026 B.n135 10.6151
R2916 B.n1020 B.n135 10.6151
R2917 B.n1020 B.n1019 10.6151
R2918 B.n1019 B.n1018 10.6151
R2919 B.n1018 B.n137 10.6151
R2920 B.n1012 B.n137 10.6151
R2921 B.n1012 B.n1011 10.6151
R2922 B.n1011 B.n1010 10.6151
R2923 B.n1010 B.n139 10.6151
R2924 B.n1004 B.n139 10.6151
R2925 B.n1004 B.n1003 10.6151
R2926 B.n1003 B.n1002 10.6151
R2927 B.n1002 B.n141 10.6151
R2928 B.n996 B.n141 10.6151
R2929 B.n996 B.n995 10.6151
R2930 B.n995 B.n994 10.6151
R2931 B.n994 B.n143 10.6151
R2932 B.n988 B.n143 10.6151
R2933 B.n988 B.n987 10.6151
R2934 B.n987 B.n986 10.6151
R2935 B.n986 B.n145 10.6151
R2936 B.n980 B.n145 10.6151
R2937 B.n978 B.n977 10.6151
R2938 B.n977 B.n149 10.6151
R2939 B.n971 B.n149 10.6151
R2940 B.n971 B.n970 10.6151
R2941 B.n970 B.n969 10.6151
R2942 B.n969 B.n151 10.6151
R2943 B.n963 B.n151 10.6151
R2944 B.n963 B.n962 10.6151
R2945 B.n962 B.n961 10.6151
R2946 B.n957 B.n956 10.6151
R2947 B.n956 B.n157 10.6151
R2948 B.n951 B.n157 10.6151
R2949 B.n951 B.n950 10.6151
R2950 B.n950 B.n949 10.6151
R2951 B.n949 B.n159 10.6151
R2952 B.n943 B.n159 10.6151
R2953 B.n943 B.n942 10.6151
R2954 B.n942 B.n941 10.6151
R2955 B.n941 B.n161 10.6151
R2956 B.n935 B.n161 10.6151
R2957 B.n935 B.n934 10.6151
R2958 B.n934 B.n933 10.6151
R2959 B.n933 B.n163 10.6151
R2960 B.n927 B.n163 10.6151
R2961 B.n927 B.n926 10.6151
R2962 B.n926 B.n925 10.6151
R2963 B.n925 B.n165 10.6151
R2964 B.n919 B.n165 10.6151
R2965 B.n919 B.n918 10.6151
R2966 B.n918 B.n917 10.6151
R2967 B.n917 B.n167 10.6151
R2968 B.n911 B.n167 10.6151
R2969 B.n911 B.n910 10.6151
R2970 B.n910 B.n909 10.6151
R2971 B.n909 B.n169 10.6151
R2972 B.n903 B.n169 10.6151
R2973 B.n903 B.n902 10.6151
R2974 B.n902 B.n901 10.6151
R2975 B.n901 B.n171 10.6151
R2976 B.n895 B.n171 10.6151
R2977 B.n895 B.n894 10.6151
R2978 B.n894 B.n893 10.6151
R2979 B.n893 B.n173 10.6151
R2980 B.n887 B.n173 10.6151
R2981 B.n887 B.n886 10.6151
R2982 B.n886 B.n885 10.6151
R2983 B.n885 B.n175 10.6151
R2984 B.n879 B.n175 10.6151
R2985 B.n879 B.n878 10.6151
R2986 B.n878 B.n877 10.6151
R2987 B.n877 B.n177 10.6151
R2988 B.n871 B.n177 10.6151
R2989 B.n871 B.n870 10.6151
R2990 B.n870 B.n869 10.6151
R2991 B.n869 B.n179 10.6151
R2992 B.n863 B.n179 10.6151
R2993 B.n485 B.n484 9.36635
R2994 B.n461 B.n346 9.36635
R2995 B.n980 B.n979 9.36635
R2996 B.n957 B.n155 9.36635
R2997 B.n270 B.t8 8.46855
R2998 B.t9 B.n1119 8.46855
R2999 B.n1212 B.n0 8.11757
R3000 B.n1212 B.n1 8.11757
R3001 B.t5 B.n246 2.82318
R3002 B.t3 B.n65 2.82318
R3003 B.n761 B.t7 1.69411
R3004 B.t4 B.n1198 1.69411
R3005 B.n484 B.n483 1.24928
R3006 B.n346 B.n342 1.24928
R3007 B.n979 B.n978 1.24928
R3008 B.n961 B.n155 1.24928
R3009 VN.n90 VN.n89 161.3
R3010 VN.n88 VN.n47 161.3
R3011 VN.n87 VN.n86 161.3
R3012 VN.n85 VN.n48 161.3
R3013 VN.n84 VN.n83 161.3
R3014 VN.n82 VN.n49 161.3
R3015 VN.n80 VN.n79 161.3
R3016 VN.n78 VN.n50 161.3
R3017 VN.n77 VN.n76 161.3
R3018 VN.n75 VN.n51 161.3
R3019 VN.n74 VN.n73 161.3
R3020 VN.n72 VN.n52 161.3
R3021 VN.n71 VN.n70 161.3
R3022 VN.n68 VN.n53 161.3
R3023 VN.n67 VN.n66 161.3
R3024 VN.n65 VN.n54 161.3
R3025 VN.n64 VN.n63 161.3
R3026 VN.n62 VN.n55 161.3
R3027 VN.n61 VN.n60 161.3
R3028 VN.n59 VN.n56 161.3
R3029 VN.n44 VN.n43 161.3
R3030 VN.n42 VN.n1 161.3
R3031 VN.n41 VN.n40 161.3
R3032 VN.n39 VN.n2 161.3
R3033 VN.n38 VN.n37 161.3
R3034 VN.n36 VN.n3 161.3
R3035 VN.n34 VN.n33 161.3
R3036 VN.n32 VN.n4 161.3
R3037 VN.n31 VN.n30 161.3
R3038 VN.n29 VN.n5 161.3
R3039 VN.n28 VN.n27 161.3
R3040 VN.n26 VN.n6 161.3
R3041 VN.n25 VN.n24 161.3
R3042 VN.n22 VN.n7 161.3
R3043 VN.n21 VN.n20 161.3
R3044 VN.n19 VN.n8 161.3
R3045 VN.n18 VN.n17 161.3
R3046 VN.n16 VN.n9 161.3
R3047 VN.n15 VN.n14 161.3
R3048 VN.n13 VN.n10 161.3
R3049 VN.n58 VN.t4 146.828
R3050 VN.n12 VN.t7 146.828
R3051 VN.n11 VN.t6 115.308
R3052 VN.n23 VN.t8 115.308
R3053 VN.n35 VN.t1 115.308
R3054 VN.n0 VN.t0 115.308
R3055 VN.n57 VN.t3 115.308
R3056 VN.n69 VN.t2 115.308
R3057 VN.n81 VN.t9 115.308
R3058 VN.n46 VN.t5 115.308
R3059 VN.n45 VN.n0 72.9405
R3060 VN.n91 VN.n46 72.9405
R3061 VN.n12 VN.n11 71.0033
R3062 VN.n58 VN.n57 71.0033
R3063 VN VN.n91 57.0359
R3064 VN.n41 VN.n2 56.5193
R3065 VN.n87 VN.n48 56.5193
R3066 VN.n17 VN.n8 50.2061
R3067 VN.n29 VN.n28 50.2061
R3068 VN.n63 VN.n54 50.2061
R3069 VN.n75 VN.n74 50.2061
R3070 VN.n17 VN.n16 30.7807
R3071 VN.n30 VN.n29 30.7807
R3072 VN.n63 VN.n62 30.7807
R3073 VN.n76 VN.n75 30.7807
R3074 VN.n15 VN.n10 24.4675
R3075 VN.n16 VN.n15 24.4675
R3076 VN.n21 VN.n8 24.4675
R3077 VN.n22 VN.n21 24.4675
R3078 VN.n24 VN.n6 24.4675
R3079 VN.n28 VN.n6 24.4675
R3080 VN.n30 VN.n4 24.4675
R3081 VN.n34 VN.n4 24.4675
R3082 VN.n37 VN.n36 24.4675
R3083 VN.n37 VN.n2 24.4675
R3084 VN.n42 VN.n41 24.4675
R3085 VN.n43 VN.n42 24.4675
R3086 VN.n62 VN.n61 24.4675
R3087 VN.n61 VN.n56 24.4675
R3088 VN.n74 VN.n52 24.4675
R3089 VN.n70 VN.n52 24.4675
R3090 VN.n68 VN.n67 24.4675
R3091 VN.n67 VN.n54 24.4675
R3092 VN.n83 VN.n48 24.4675
R3093 VN.n83 VN.n82 24.4675
R3094 VN.n80 VN.n50 24.4675
R3095 VN.n76 VN.n50 24.4675
R3096 VN.n89 VN.n88 24.4675
R3097 VN.n88 VN.n87 24.4675
R3098 VN.n36 VN.n35 22.0208
R3099 VN.n82 VN.n81 22.0208
R3100 VN.n43 VN.n0 17.1274
R3101 VN.n89 VN.n46 17.1274
R3102 VN.n23 VN.n22 12.234
R3103 VN.n24 VN.n23 12.234
R3104 VN.n70 VN.n69 12.234
R3105 VN.n69 VN.n68 12.234
R3106 VN.n59 VN.n58 5.75995
R3107 VN.n13 VN.n12 5.75995
R3108 VN.n11 VN.n10 2.4472
R3109 VN.n35 VN.n34 2.4472
R3110 VN.n57 VN.n56 2.4472
R3111 VN.n81 VN.n80 2.4472
R3112 VN.n91 VN.n90 0.354971
R3113 VN.n45 VN.n44 0.354971
R3114 VN VN.n45 0.26696
R3115 VN.n90 VN.n47 0.189894
R3116 VN.n86 VN.n47 0.189894
R3117 VN.n86 VN.n85 0.189894
R3118 VN.n85 VN.n84 0.189894
R3119 VN.n84 VN.n49 0.189894
R3120 VN.n79 VN.n49 0.189894
R3121 VN.n79 VN.n78 0.189894
R3122 VN.n78 VN.n77 0.189894
R3123 VN.n77 VN.n51 0.189894
R3124 VN.n73 VN.n51 0.189894
R3125 VN.n73 VN.n72 0.189894
R3126 VN.n72 VN.n71 0.189894
R3127 VN.n71 VN.n53 0.189894
R3128 VN.n66 VN.n53 0.189894
R3129 VN.n66 VN.n65 0.189894
R3130 VN.n65 VN.n64 0.189894
R3131 VN.n64 VN.n55 0.189894
R3132 VN.n60 VN.n55 0.189894
R3133 VN.n60 VN.n59 0.189894
R3134 VN.n14 VN.n13 0.189894
R3135 VN.n14 VN.n9 0.189894
R3136 VN.n18 VN.n9 0.189894
R3137 VN.n19 VN.n18 0.189894
R3138 VN.n20 VN.n19 0.189894
R3139 VN.n20 VN.n7 0.189894
R3140 VN.n25 VN.n7 0.189894
R3141 VN.n26 VN.n25 0.189894
R3142 VN.n27 VN.n26 0.189894
R3143 VN.n27 VN.n5 0.189894
R3144 VN.n31 VN.n5 0.189894
R3145 VN.n32 VN.n31 0.189894
R3146 VN.n33 VN.n32 0.189894
R3147 VN.n33 VN.n3 0.189894
R3148 VN.n38 VN.n3 0.189894
R3149 VN.n39 VN.n38 0.189894
R3150 VN.n40 VN.n39 0.189894
R3151 VN.n40 VN.n1 0.189894
R3152 VN.n44 VN.n1 0.189894
R3153 VDD2.n153 VDD2.n81 289.615
R3154 VDD2.n72 VDD2.n0 289.615
R3155 VDD2.n154 VDD2.n153 185
R3156 VDD2.n152 VDD2.n151 185
R3157 VDD2.n85 VDD2.n84 185
R3158 VDD2.n146 VDD2.n145 185
R3159 VDD2.n144 VDD2.n143 185
R3160 VDD2.n89 VDD2.n88 185
R3161 VDD2.n138 VDD2.n137 185
R3162 VDD2.n136 VDD2.n135 185
R3163 VDD2.n93 VDD2.n92 185
R3164 VDD2.n130 VDD2.n129 185
R3165 VDD2.n128 VDD2.n95 185
R3166 VDD2.n127 VDD2.n126 185
R3167 VDD2.n98 VDD2.n96 185
R3168 VDD2.n121 VDD2.n120 185
R3169 VDD2.n119 VDD2.n118 185
R3170 VDD2.n102 VDD2.n101 185
R3171 VDD2.n113 VDD2.n112 185
R3172 VDD2.n111 VDD2.n110 185
R3173 VDD2.n106 VDD2.n105 185
R3174 VDD2.n24 VDD2.n23 185
R3175 VDD2.n29 VDD2.n28 185
R3176 VDD2.n31 VDD2.n30 185
R3177 VDD2.n20 VDD2.n19 185
R3178 VDD2.n37 VDD2.n36 185
R3179 VDD2.n39 VDD2.n38 185
R3180 VDD2.n16 VDD2.n15 185
R3181 VDD2.n46 VDD2.n45 185
R3182 VDD2.n47 VDD2.n14 185
R3183 VDD2.n49 VDD2.n48 185
R3184 VDD2.n12 VDD2.n11 185
R3185 VDD2.n55 VDD2.n54 185
R3186 VDD2.n57 VDD2.n56 185
R3187 VDD2.n8 VDD2.n7 185
R3188 VDD2.n63 VDD2.n62 185
R3189 VDD2.n65 VDD2.n64 185
R3190 VDD2.n4 VDD2.n3 185
R3191 VDD2.n71 VDD2.n70 185
R3192 VDD2.n73 VDD2.n72 185
R3193 VDD2.n107 VDD2.t4 149.524
R3194 VDD2.n25 VDD2.t2 149.524
R3195 VDD2.n153 VDD2.n152 104.615
R3196 VDD2.n152 VDD2.n84 104.615
R3197 VDD2.n145 VDD2.n84 104.615
R3198 VDD2.n145 VDD2.n144 104.615
R3199 VDD2.n144 VDD2.n88 104.615
R3200 VDD2.n137 VDD2.n88 104.615
R3201 VDD2.n137 VDD2.n136 104.615
R3202 VDD2.n136 VDD2.n92 104.615
R3203 VDD2.n129 VDD2.n92 104.615
R3204 VDD2.n129 VDD2.n128 104.615
R3205 VDD2.n128 VDD2.n127 104.615
R3206 VDD2.n127 VDD2.n96 104.615
R3207 VDD2.n120 VDD2.n96 104.615
R3208 VDD2.n120 VDD2.n119 104.615
R3209 VDD2.n119 VDD2.n101 104.615
R3210 VDD2.n112 VDD2.n101 104.615
R3211 VDD2.n112 VDD2.n111 104.615
R3212 VDD2.n111 VDD2.n105 104.615
R3213 VDD2.n29 VDD2.n23 104.615
R3214 VDD2.n30 VDD2.n29 104.615
R3215 VDD2.n30 VDD2.n19 104.615
R3216 VDD2.n37 VDD2.n19 104.615
R3217 VDD2.n38 VDD2.n37 104.615
R3218 VDD2.n38 VDD2.n15 104.615
R3219 VDD2.n46 VDD2.n15 104.615
R3220 VDD2.n47 VDD2.n46 104.615
R3221 VDD2.n48 VDD2.n47 104.615
R3222 VDD2.n48 VDD2.n11 104.615
R3223 VDD2.n55 VDD2.n11 104.615
R3224 VDD2.n56 VDD2.n55 104.615
R3225 VDD2.n56 VDD2.n7 104.615
R3226 VDD2.n63 VDD2.n7 104.615
R3227 VDD2.n64 VDD2.n63 104.615
R3228 VDD2.n64 VDD2.n3 104.615
R3229 VDD2.n71 VDD2.n3 104.615
R3230 VDD2.n72 VDD2.n71 104.615
R3231 VDD2.n80 VDD2.n79 62.1489
R3232 VDD2 VDD2.n161 62.146
R3233 VDD2.n160 VDD2.n159 60.0706
R3234 VDD2.n78 VDD2.n77 60.0706
R3235 VDD2.t4 VDD2.n105 52.3082
R3236 VDD2.t2 VDD2.n23 52.3082
R3237 VDD2.n78 VDD2.n76 50.3514
R3238 VDD2.n158 VDD2.n80 49.4782
R3239 VDD2.n158 VDD2.n157 47.5066
R3240 VDD2.n130 VDD2.n95 13.1884
R3241 VDD2.n49 VDD2.n14 13.1884
R3242 VDD2.n131 VDD2.n93 12.8005
R3243 VDD2.n126 VDD2.n97 12.8005
R3244 VDD2.n45 VDD2.n44 12.8005
R3245 VDD2.n50 VDD2.n12 12.8005
R3246 VDD2.n135 VDD2.n134 12.0247
R3247 VDD2.n125 VDD2.n98 12.0247
R3248 VDD2.n43 VDD2.n16 12.0247
R3249 VDD2.n54 VDD2.n53 12.0247
R3250 VDD2.n138 VDD2.n91 11.249
R3251 VDD2.n122 VDD2.n121 11.249
R3252 VDD2.n40 VDD2.n39 11.249
R3253 VDD2.n57 VDD2.n10 11.249
R3254 VDD2.n139 VDD2.n89 10.4732
R3255 VDD2.n118 VDD2.n100 10.4732
R3256 VDD2.n36 VDD2.n18 10.4732
R3257 VDD2.n58 VDD2.n8 10.4732
R3258 VDD2.n107 VDD2.n106 10.2747
R3259 VDD2.n25 VDD2.n24 10.2747
R3260 VDD2.n143 VDD2.n142 9.69747
R3261 VDD2.n117 VDD2.n102 9.69747
R3262 VDD2.n35 VDD2.n20 9.69747
R3263 VDD2.n62 VDD2.n61 9.69747
R3264 VDD2.n157 VDD2.n156 9.45567
R3265 VDD2.n76 VDD2.n75 9.45567
R3266 VDD2.n109 VDD2.n108 9.3005
R3267 VDD2.n104 VDD2.n103 9.3005
R3268 VDD2.n115 VDD2.n114 9.3005
R3269 VDD2.n117 VDD2.n116 9.3005
R3270 VDD2.n100 VDD2.n99 9.3005
R3271 VDD2.n123 VDD2.n122 9.3005
R3272 VDD2.n125 VDD2.n124 9.3005
R3273 VDD2.n97 VDD2.n94 9.3005
R3274 VDD2.n156 VDD2.n155 9.3005
R3275 VDD2.n83 VDD2.n82 9.3005
R3276 VDD2.n150 VDD2.n149 9.3005
R3277 VDD2.n148 VDD2.n147 9.3005
R3278 VDD2.n87 VDD2.n86 9.3005
R3279 VDD2.n142 VDD2.n141 9.3005
R3280 VDD2.n140 VDD2.n139 9.3005
R3281 VDD2.n91 VDD2.n90 9.3005
R3282 VDD2.n134 VDD2.n133 9.3005
R3283 VDD2.n132 VDD2.n131 9.3005
R3284 VDD2.n2 VDD2.n1 9.3005
R3285 VDD2.n75 VDD2.n74 9.3005
R3286 VDD2.n67 VDD2.n66 9.3005
R3287 VDD2.n6 VDD2.n5 9.3005
R3288 VDD2.n61 VDD2.n60 9.3005
R3289 VDD2.n59 VDD2.n58 9.3005
R3290 VDD2.n10 VDD2.n9 9.3005
R3291 VDD2.n53 VDD2.n52 9.3005
R3292 VDD2.n51 VDD2.n50 9.3005
R3293 VDD2.n27 VDD2.n26 9.3005
R3294 VDD2.n22 VDD2.n21 9.3005
R3295 VDD2.n33 VDD2.n32 9.3005
R3296 VDD2.n35 VDD2.n34 9.3005
R3297 VDD2.n18 VDD2.n17 9.3005
R3298 VDD2.n41 VDD2.n40 9.3005
R3299 VDD2.n43 VDD2.n42 9.3005
R3300 VDD2.n44 VDD2.n13 9.3005
R3301 VDD2.n69 VDD2.n68 9.3005
R3302 VDD2.n146 VDD2.n87 8.92171
R3303 VDD2.n114 VDD2.n113 8.92171
R3304 VDD2.n32 VDD2.n31 8.92171
R3305 VDD2.n65 VDD2.n6 8.92171
R3306 VDD2.n157 VDD2.n81 8.14595
R3307 VDD2.n147 VDD2.n85 8.14595
R3308 VDD2.n110 VDD2.n104 8.14595
R3309 VDD2.n28 VDD2.n22 8.14595
R3310 VDD2.n66 VDD2.n4 8.14595
R3311 VDD2.n76 VDD2.n0 8.14595
R3312 VDD2.n155 VDD2.n154 7.3702
R3313 VDD2.n151 VDD2.n150 7.3702
R3314 VDD2.n109 VDD2.n106 7.3702
R3315 VDD2.n27 VDD2.n24 7.3702
R3316 VDD2.n70 VDD2.n69 7.3702
R3317 VDD2.n74 VDD2.n73 7.3702
R3318 VDD2.n154 VDD2.n83 6.59444
R3319 VDD2.n151 VDD2.n83 6.59444
R3320 VDD2.n70 VDD2.n2 6.59444
R3321 VDD2.n73 VDD2.n2 6.59444
R3322 VDD2.n155 VDD2.n81 5.81868
R3323 VDD2.n150 VDD2.n85 5.81868
R3324 VDD2.n110 VDD2.n109 5.81868
R3325 VDD2.n28 VDD2.n27 5.81868
R3326 VDD2.n69 VDD2.n4 5.81868
R3327 VDD2.n74 VDD2.n0 5.81868
R3328 VDD2.n147 VDD2.n146 5.04292
R3329 VDD2.n113 VDD2.n104 5.04292
R3330 VDD2.n31 VDD2.n22 5.04292
R3331 VDD2.n66 VDD2.n65 5.04292
R3332 VDD2.n143 VDD2.n87 4.26717
R3333 VDD2.n114 VDD2.n102 4.26717
R3334 VDD2.n32 VDD2.n20 4.26717
R3335 VDD2.n62 VDD2.n6 4.26717
R3336 VDD2.n142 VDD2.n89 3.49141
R3337 VDD2.n118 VDD2.n117 3.49141
R3338 VDD2.n36 VDD2.n35 3.49141
R3339 VDD2.n61 VDD2.n8 3.49141
R3340 VDD2.n160 VDD2.n158 2.84533
R3341 VDD2.n108 VDD2.n107 2.84303
R3342 VDD2.n26 VDD2.n25 2.84303
R3343 VDD2.n139 VDD2.n138 2.71565
R3344 VDD2.n121 VDD2.n100 2.71565
R3345 VDD2.n39 VDD2.n18 2.71565
R3346 VDD2.n58 VDD2.n57 2.71565
R3347 VDD2.n135 VDD2.n91 1.93989
R3348 VDD2.n122 VDD2.n98 1.93989
R3349 VDD2.n40 VDD2.n16 1.93989
R3350 VDD2.n54 VDD2.n10 1.93989
R3351 VDD2.n161 VDD2.t6 1.39388
R3352 VDD2.n161 VDD2.t5 1.39388
R3353 VDD2.n159 VDD2.t0 1.39388
R3354 VDD2.n159 VDD2.t7 1.39388
R3355 VDD2.n79 VDD2.t8 1.39388
R3356 VDD2.n79 VDD2.t9 1.39388
R3357 VDD2.n77 VDD2.t3 1.39388
R3358 VDD2.n77 VDD2.t1 1.39388
R3359 VDD2.n134 VDD2.n93 1.16414
R3360 VDD2.n126 VDD2.n125 1.16414
R3361 VDD2.n45 VDD2.n43 1.16414
R3362 VDD2.n53 VDD2.n12 1.16414
R3363 VDD2 VDD2.n160 0.769897
R3364 VDD2.n80 VDD2.n78 0.656361
R3365 VDD2.n131 VDD2.n130 0.388379
R3366 VDD2.n97 VDD2.n95 0.388379
R3367 VDD2.n44 VDD2.n14 0.388379
R3368 VDD2.n50 VDD2.n49 0.388379
R3369 VDD2.n156 VDD2.n82 0.155672
R3370 VDD2.n149 VDD2.n82 0.155672
R3371 VDD2.n149 VDD2.n148 0.155672
R3372 VDD2.n148 VDD2.n86 0.155672
R3373 VDD2.n141 VDD2.n86 0.155672
R3374 VDD2.n141 VDD2.n140 0.155672
R3375 VDD2.n140 VDD2.n90 0.155672
R3376 VDD2.n133 VDD2.n90 0.155672
R3377 VDD2.n133 VDD2.n132 0.155672
R3378 VDD2.n132 VDD2.n94 0.155672
R3379 VDD2.n124 VDD2.n94 0.155672
R3380 VDD2.n124 VDD2.n123 0.155672
R3381 VDD2.n123 VDD2.n99 0.155672
R3382 VDD2.n116 VDD2.n99 0.155672
R3383 VDD2.n116 VDD2.n115 0.155672
R3384 VDD2.n115 VDD2.n103 0.155672
R3385 VDD2.n108 VDD2.n103 0.155672
R3386 VDD2.n26 VDD2.n21 0.155672
R3387 VDD2.n33 VDD2.n21 0.155672
R3388 VDD2.n34 VDD2.n33 0.155672
R3389 VDD2.n34 VDD2.n17 0.155672
R3390 VDD2.n41 VDD2.n17 0.155672
R3391 VDD2.n42 VDD2.n41 0.155672
R3392 VDD2.n42 VDD2.n13 0.155672
R3393 VDD2.n51 VDD2.n13 0.155672
R3394 VDD2.n52 VDD2.n51 0.155672
R3395 VDD2.n52 VDD2.n9 0.155672
R3396 VDD2.n59 VDD2.n9 0.155672
R3397 VDD2.n60 VDD2.n59 0.155672
R3398 VDD2.n60 VDD2.n5 0.155672
R3399 VDD2.n67 VDD2.n5 0.155672
R3400 VDD2.n68 VDD2.n67 0.155672
R3401 VDD2.n68 VDD2.n1 0.155672
R3402 VDD2.n75 VDD2.n1 0.155672
C0 VP VDD1 13.3269f
C1 VP VN 9.35785f
C2 VP VDD2 0.630981f
C3 VDD1 VN 0.154248f
C4 VP VTAIL 13.5713f
C5 VDD1 VDD2 2.41587f
C6 VDD2 VN 12.8544f
C7 VDD1 VTAIL 11.4667f
C8 VN VTAIL 13.557f
C9 VDD2 VTAIL 11.52f
C10 VDD2 B 8.03546f
C11 VDD1 B 8.003937f
C12 VTAIL B 9.390512f
C13 VN B 20.095419f
C14 VP B 18.621319f
C15 VDD2.n0 B 0.034626f
C16 VDD2.n1 B 0.024057f
C17 VDD2.n2 B 0.012927f
C18 VDD2.n3 B 0.030555f
C19 VDD2.n4 B 0.013688f
C20 VDD2.n5 B 0.024057f
C21 VDD2.n6 B 0.012927f
C22 VDD2.n7 B 0.030555f
C23 VDD2.n8 B 0.013688f
C24 VDD2.n9 B 0.024057f
C25 VDD2.n10 B 0.012927f
C26 VDD2.n11 B 0.030555f
C27 VDD2.n12 B 0.013688f
C28 VDD2.n13 B 0.024057f
C29 VDD2.n14 B 0.013308f
C30 VDD2.n15 B 0.030555f
C31 VDD2.n16 B 0.013688f
C32 VDD2.n17 B 0.024057f
C33 VDD2.n18 B 0.012927f
C34 VDD2.n19 B 0.030555f
C35 VDD2.n20 B 0.013688f
C36 VDD2.n21 B 0.024057f
C37 VDD2.n22 B 0.012927f
C38 VDD2.n23 B 0.022917f
C39 VDD2.n24 B 0.0216f
C40 VDD2.t2 B 0.051892f
C41 VDD2.n25 B 0.193862f
C42 VDD2.n26 B 1.45013f
C43 VDD2.n27 B 0.012927f
C44 VDD2.n28 B 0.013688f
C45 VDD2.n29 B 0.030555f
C46 VDD2.n30 B 0.030555f
C47 VDD2.n31 B 0.013688f
C48 VDD2.n32 B 0.012927f
C49 VDD2.n33 B 0.024057f
C50 VDD2.n34 B 0.024057f
C51 VDD2.n35 B 0.012927f
C52 VDD2.n36 B 0.013688f
C53 VDD2.n37 B 0.030555f
C54 VDD2.n38 B 0.030555f
C55 VDD2.n39 B 0.013688f
C56 VDD2.n40 B 0.012927f
C57 VDD2.n41 B 0.024057f
C58 VDD2.n42 B 0.024057f
C59 VDD2.n43 B 0.012927f
C60 VDD2.n44 B 0.012927f
C61 VDD2.n45 B 0.013688f
C62 VDD2.n46 B 0.030555f
C63 VDD2.n47 B 0.030555f
C64 VDD2.n48 B 0.030555f
C65 VDD2.n49 B 0.013308f
C66 VDD2.n50 B 0.012927f
C67 VDD2.n51 B 0.024057f
C68 VDD2.n52 B 0.024057f
C69 VDD2.n53 B 0.012927f
C70 VDD2.n54 B 0.013688f
C71 VDD2.n55 B 0.030555f
C72 VDD2.n56 B 0.030555f
C73 VDD2.n57 B 0.013688f
C74 VDD2.n58 B 0.012927f
C75 VDD2.n59 B 0.024057f
C76 VDD2.n60 B 0.024057f
C77 VDD2.n61 B 0.012927f
C78 VDD2.n62 B 0.013688f
C79 VDD2.n63 B 0.030555f
C80 VDD2.n64 B 0.030555f
C81 VDD2.n65 B 0.013688f
C82 VDD2.n66 B 0.012927f
C83 VDD2.n67 B 0.024057f
C84 VDD2.n68 B 0.024057f
C85 VDD2.n69 B 0.012927f
C86 VDD2.n70 B 0.013688f
C87 VDD2.n71 B 0.030555f
C88 VDD2.n72 B 0.067583f
C89 VDD2.n73 B 0.013688f
C90 VDD2.n74 B 0.012927f
C91 VDD2.n75 B 0.053307f
C92 VDD2.n76 B 0.069523f
C93 VDD2.t3 B 0.270143f
C94 VDD2.t1 B 0.270143f
C95 VDD2.n77 B 2.42804f
C96 VDD2.n78 B 0.726378f
C97 VDD2.t8 B 0.270143f
C98 VDD2.t9 B 0.270143f
C99 VDD2.n79 B 2.44794f
C100 VDD2.n80 B 3.11872f
C101 VDD2.n81 B 0.034626f
C102 VDD2.n82 B 0.024057f
C103 VDD2.n83 B 0.012927f
C104 VDD2.n84 B 0.030555f
C105 VDD2.n85 B 0.013688f
C106 VDD2.n86 B 0.024057f
C107 VDD2.n87 B 0.012927f
C108 VDD2.n88 B 0.030555f
C109 VDD2.n89 B 0.013688f
C110 VDD2.n90 B 0.024057f
C111 VDD2.n91 B 0.012927f
C112 VDD2.n92 B 0.030555f
C113 VDD2.n93 B 0.013688f
C114 VDD2.n94 B 0.024057f
C115 VDD2.n95 B 0.013308f
C116 VDD2.n96 B 0.030555f
C117 VDD2.n97 B 0.012927f
C118 VDD2.n98 B 0.013688f
C119 VDD2.n99 B 0.024057f
C120 VDD2.n100 B 0.012927f
C121 VDD2.n101 B 0.030555f
C122 VDD2.n102 B 0.013688f
C123 VDD2.n103 B 0.024057f
C124 VDD2.n104 B 0.012927f
C125 VDD2.n105 B 0.022917f
C126 VDD2.n106 B 0.0216f
C127 VDD2.t4 B 0.051892f
C128 VDD2.n107 B 0.193862f
C129 VDD2.n108 B 1.45013f
C130 VDD2.n109 B 0.012927f
C131 VDD2.n110 B 0.013688f
C132 VDD2.n111 B 0.030555f
C133 VDD2.n112 B 0.030555f
C134 VDD2.n113 B 0.013688f
C135 VDD2.n114 B 0.012927f
C136 VDD2.n115 B 0.024057f
C137 VDD2.n116 B 0.024057f
C138 VDD2.n117 B 0.012927f
C139 VDD2.n118 B 0.013688f
C140 VDD2.n119 B 0.030555f
C141 VDD2.n120 B 0.030555f
C142 VDD2.n121 B 0.013688f
C143 VDD2.n122 B 0.012927f
C144 VDD2.n123 B 0.024057f
C145 VDD2.n124 B 0.024057f
C146 VDD2.n125 B 0.012927f
C147 VDD2.n126 B 0.013688f
C148 VDD2.n127 B 0.030555f
C149 VDD2.n128 B 0.030555f
C150 VDD2.n129 B 0.030555f
C151 VDD2.n130 B 0.013308f
C152 VDD2.n131 B 0.012927f
C153 VDD2.n132 B 0.024057f
C154 VDD2.n133 B 0.024057f
C155 VDD2.n134 B 0.012927f
C156 VDD2.n135 B 0.013688f
C157 VDD2.n136 B 0.030555f
C158 VDD2.n137 B 0.030555f
C159 VDD2.n138 B 0.013688f
C160 VDD2.n139 B 0.012927f
C161 VDD2.n140 B 0.024057f
C162 VDD2.n141 B 0.024057f
C163 VDD2.n142 B 0.012927f
C164 VDD2.n143 B 0.013688f
C165 VDD2.n144 B 0.030555f
C166 VDD2.n145 B 0.030555f
C167 VDD2.n146 B 0.013688f
C168 VDD2.n147 B 0.012927f
C169 VDD2.n148 B 0.024057f
C170 VDD2.n149 B 0.024057f
C171 VDD2.n150 B 0.012927f
C172 VDD2.n151 B 0.013688f
C173 VDD2.n152 B 0.030555f
C174 VDD2.n153 B 0.067583f
C175 VDD2.n154 B 0.013688f
C176 VDD2.n155 B 0.012927f
C177 VDD2.n156 B 0.053307f
C178 VDD2.n157 B 0.054521f
C179 VDD2.n158 B 3.08144f
C180 VDD2.t0 B 0.270143f
C181 VDD2.t7 B 0.270143f
C182 VDD2.n159 B 2.42804f
C183 VDD2.n160 B 0.483796f
C184 VDD2.t6 B 0.270143f
C185 VDD2.t5 B 0.270143f
C186 VDD2.n161 B 2.4479f
C187 VN.t0 B 2.23246f
C188 VN.n0 B 0.851852f
C189 VN.n1 B 0.019329f
C190 VN.n2 B 0.025523f
C191 VN.n3 B 0.019329f
C192 VN.t1 B 2.23246f
C193 VN.n4 B 0.036024f
C194 VN.n5 B 0.019329f
C195 VN.n6 B 0.036024f
C196 VN.n7 B 0.019329f
C197 VN.t8 B 2.23246f
C198 VN.n8 B 0.035475f
C199 VN.n9 B 0.019329f
C200 VN.n10 B 0.020017f
C201 VN.t6 B 2.23246f
C202 VN.n11 B 0.834204f
C203 VN.t7 B 2.42695f
C204 VN.n12 B 0.812215f
C205 VN.n13 B 0.209106f
C206 VN.n14 B 0.019329f
C207 VN.n15 B 0.036024f
C208 VN.n16 B 0.038722f
C209 VN.n17 B 0.018259f
C210 VN.n18 B 0.019329f
C211 VN.n19 B 0.019329f
C212 VN.n20 B 0.019329f
C213 VN.n21 B 0.036024f
C214 VN.n22 B 0.027131f
C215 VN.n23 B 0.779813f
C216 VN.n24 B 0.027131f
C217 VN.n25 B 0.019329f
C218 VN.n26 B 0.019329f
C219 VN.n27 B 0.019329f
C220 VN.n28 B 0.035475f
C221 VN.n29 B 0.018259f
C222 VN.n30 B 0.038722f
C223 VN.n31 B 0.019329f
C224 VN.n32 B 0.019329f
C225 VN.n33 B 0.019329f
C226 VN.n34 B 0.020017f
C227 VN.n35 B 0.779813f
C228 VN.n36 B 0.034245f
C229 VN.n37 B 0.036024f
C230 VN.n38 B 0.019329f
C231 VN.n39 B 0.019329f
C232 VN.n40 B 0.019329f
C233 VN.n41 B 0.030909f
C234 VN.n42 B 0.036024f
C235 VN.n43 B 0.030688f
C236 VN.n44 B 0.031196f
C237 VN.n45 B 0.042377f
C238 VN.t5 B 2.23246f
C239 VN.n46 B 0.851852f
C240 VN.n47 B 0.019329f
C241 VN.n48 B 0.025523f
C242 VN.n49 B 0.019329f
C243 VN.t9 B 2.23246f
C244 VN.n50 B 0.036024f
C245 VN.n51 B 0.019329f
C246 VN.n52 B 0.036024f
C247 VN.n53 B 0.019329f
C248 VN.t2 B 2.23246f
C249 VN.n54 B 0.035475f
C250 VN.n55 B 0.019329f
C251 VN.n56 B 0.020017f
C252 VN.t4 B 2.42695f
C253 VN.t3 B 2.23246f
C254 VN.n57 B 0.834204f
C255 VN.n58 B 0.812215f
C256 VN.n59 B 0.209106f
C257 VN.n60 B 0.019329f
C258 VN.n61 B 0.036024f
C259 VN.n62 B 0.038722f
C260 VN.n63 B 0.018259f
C261 VN.n64 B 0.019329f
C262 VN.n65 B 0.019329f
C263 VN.n66 B 0.019329f
C264 VN.n67 B 0.036024f
C265 VN.n68 B 0.027131f
C266 VN.n69 B 0.779813f
C267 VN.n70 B 0.027131f
C268 VN.n71 B 0.019329f
C269 VN.n72 B 0.019329f
C270 VN.n73 B 0.019329f
C271 VN.n74 B 0.035475f
C272 VN.n75 B 0.018259f
C273 VN.n76 B 0.038722f
C274 VN.n77 B 0.019329f
C275 VN.n78 B 0.019329f
C276 VN.n79 B 0.019329f
C277 VN.n80 B 0.020017f
C278 VN.n81 B 0.779813f
C279 VN.n82 B 0.034245f
C280 VN.n83 B 0.036024f
C281 VN.n84 B 0.019329f
C282 VN.n85 B 0.019329f
C283 VN.n86 B 0.019329f
C284 VN.n87 B 0.030909f
C285 VN.n88 B 0.036024f
C286 VN.n89 B 0.030688f
C287 VN.n90 B 0.031196f
C288 VN.n91 B 1.31828f
C289 VDD1.n0 B 0.035027f
C290 VDD1.n1 B 0.024336f
C291 VDD1.n2 B 0.013077f
C292 VDD1.n3 B 0.030909f
C293 VDD1.n4 B 0.013846f
C294 VDD1.n5 B 0.024336f
C295 VDD1.n6 B 0.013077f
C296 VDD1.n7 B 0.030909f
C297 VDD1.n8 B 0.013846f
C298 VDD1.n9 B 0.024336f
C299 VDD1.n10 B 0.013077f
C300 VDD1.n11 B 0.030909f
C301 VDD1.n12 B 0.013846f
C302 VDD1.n13 B 0.024336f
C303 VDD1.n14 B 0.013462f
C304 VDD1.n15 B 0.030909f
C305 VDD1.n16 B 0.013077f
C306 VDD1.n17 B 0.013846f
C307 VDD1.n18 B 0.024336f
C308 VDD1.n19 B 0.013077f
C309 VDD1.n20 B 0.030909f
C310 VDD1.n21 B 0.013846f
C311 VDD1.n22 B 0.024336f
C312 VDD1.n23 B 0.013077f
C313 VDD1.n24 B 0.023182f
C314 VDD1.n25 B 0.02185f
C315 VDD1.t3 B 0.052493f
C316 VDD1.n26 B 0.196105f
C317 VDD1.n27 B 1.46691f
C318 VDD1.n28 B 0.013077f
C319 VDD1.n29 B 0.013846f
C320 VDD1.n30 B 0.030909f
C321 VDD1.n31 B 0.030909f
C322 VDD1.n32 B 0.013846f
C323 VDD1.n33 B 0.013077f
C324 VDD1.n34 B 0.024336f
C325 VDD1.n35 B 0.024336f
C326 VDD1.n36 B 0.013077f
C327 VDD1.n37 B 0.013846f
C328 VDD1.n38 B 0.030909f
C329 VDD1.n39 B 0.030909f
C330 VDD1.n40 B 0.013846f
C331 VDD1.n41 B 0.013077f
C332 VDD1.n42 B 0.024336f
C333 VDD1.n43 B 0.024336f
C334 VDD1.n44 B 0.013077f
C335 VDD1.n45 B 0.013846f
C336 VDD1.n46 B 0.030909f
C337 VDD1.n47 B 0.030909f
C338 VDD1.n48 B 0.030909f
C339 VDD1.n49 B 0.013462f
C340 VDD1.n50 B 0.013077f
C341 VDD1.n51 B 0.024336f
C342 VDD1.n52 B 0.024336f
C343 VDD1.n53 B 0.013077f
C344 VDD1.n54 B 0.013846f
C345 VDD1.n55 B 0.030909f
C346 VDD1.n56 B 0.030909f
C347 VDD1.n57 B 0.013846f
C348 VDD1.n58 B 0.013077f
C349 VDD1.n59 B 0.024336f
C350 VDD1.n60 B 0.024336f
C351 VDD1.n61 B 0.013077f
C352 VDD1.n62 B 0.013846f
C353 VDD1.n63 B 0.030909f
C354 VDD1.n64 B 0.030909f
C355 VDD1.n65 B 0.013846f
C356 VDD1.n66 B 0.013077f
C357 VDD1.n67 B 0.024336f
C358 VDD1.n68 B 0.024336f
C359 VDD1.n69 B 0.013077f
C360 VDD1.n70 B 0.013846f
C361 VDD1.n71 B 0.030909f
C362 VDD1.n72 B 0.068365f
C363 VDD1.n73 B 0.013846f
C364 VDD1.n74 B 0.013077f
C365 VDD1.n75 B 0.053924f
C366 VDD1.n76 B 0.070328f
C367 VDD1.t5 B 0.273269f
C368 VDD1.t0 B 0.273269f
C369 VDD1.n77 B 2.45614f
C370 VDD1.n78 B 0.742823f
C371 VDD1.n79 B 0.035027f
C372 VDD1.n80 B 0.024336f
C373 VDD1.n81 B 0.013077f
C374 VDD1.n82 B 0.030909f
C375 VDD1.n83 B 0.013846f
C376 VDD1.n84 B 0.024336f
C377 VDD1.n85 B 0.013077f
C378 VDD1.n86 B 0.030909f
C379 VDD1.n87 B 0.013846f
C380 VDD1.n88 B 0.024336f
C381 VDD1.n89 B 0.013077f
C382 VDD1.n90 B 0.030909f
C383 VDD1.n91 B 0.013846f
C384 VDD1.n92 B 0.024336f
C385 VDD1.n93 B 0.013462f
C386 VDD1.n94 B 0.030909f
C387 VDD1.n95 B 0.013846f
C388 VDD1.n96 B 0.024336f
C389 VDD1.n97 B 0.013077f
C390 VDD1.n98 B 0.030909f
C391 VDD1.n99 B 0.013846f
C392 VDD1.n100 B 0.024336f
C393 VDD1.n101 B 0.013077f
C394 VDD1.n102 B 0.023182f
C395 VDD1.n103 B 0.02185f
C396 VDD1.t6 B 0.052493f
C397 VDD1.n104 B 0.196105f
C398 VDD1.n105 B 1.46691f
C399 VDD1.n106 B 0.013077f
C400 VDD1.n107 B 0.013846f
C401 VDD1.n108 B 0.030909f
C402 VDD1.n109 B 0.030909f
C403 VDD1.n110 B 0.013846f
C404 VDD1.n111 B 0.013077f
C405 VDD1.n112 B 0.024336f
C406 VDD1.n113 B 0.024336f
C407 VDD1.n114 B 0.013077f
C408 VDD1.n115 B 0.013846f
C409 VDD1.n116 B 0.030909f
C410 VDD1.n117 B 0.030909f
C411 VDD1.n118 B 0.013846f
C412 VDD1.n119 B 0.013077f
C413 VDD1.n120 B 0.024336f
C414 VDD1.n121 B 0.024336f
C415 VDD1.n122 B 0.013077f
C416 VDD1.n123 B 0.013077f
C417 VDD1.n124 B 0.013846f
C418 VDD1.n125 B 0.030909f
C419 VDD1.n126 B 0.030909f
C420 VDD1.n127 B 0.030909f
C421 VDD1.n128 B 0.013462f
C422 VDD1.n129 B 0.013077f
C423 VDD1.n130 B 0.024336f
C424 VDD1.n131 B 0.024336f
C425 VDD1.n132 B 0.013077f
C426 VDD1.n133 B 0.013846f
C427 VDD1.n134 B 0.030909f
C428 VDD1.n135 B 0.030909f
C429 VDD1.n136 B 0.013846f
C430 VDD1.n137 B 0.013077f
C431 VDD1.n138 B 0.024336f
C432 VDD1.n139 B 0.024336f
C433 VDD1.n140 B 0.013077f
C434 VDD1.n141 B 0.013846f
C435 VDD1.n142 B 0.030909f
C436 VDD1.n143 B 0.030909f
C437 VDD1.n144 B 0.013846f
C438 VDD1.n145 B 0.013077f
C439 VDD1.n146 B 0.024336f
C440 VDD1.n147 B 0.024336f
C441 VDD1.n148 B 0.013077f
C442 VDD1.n149 B 0.013846f
C443 VDD1.n150 B 0.030909f
C444 VDD1.n151 B 0.068365f
C445 VDD1.n152 B 0.013846f
C446 VDD1.n153 B 0.013077f
C447 VDD1.n154 B 0.053924f
C448 VDD1.n155 B 0.070328f
C449 VDD1.t7 B 0.273269f
C450 VDD1.t9 B 0.273269f
C451 VDD1.n156 B 2.45613f
C452 VDD1.n157 B 0.734783f
C453 VDD1.t8 B 0.273269f
C454 VDD1.t1 B 0.273269f
C455 VDD1.n158 B 2.47627f
C456 VDD1.n159 B 3.28781f
C457 VDD1.t2 B 0.273269f
C458 VDD1.t4 B 0.273269f
C459 VDD1.n160 B 2.45614f
C460 VDD1.n161 B 3.40698f
C461 VTAIL.t4 B 0.276755f
C462 VTAIL.t6 B 0.276755f
C463 VTAIL.n0 B 2.40908f
C464 VTAIL.n1 B 0.577835f
C465 VTAIL.n2 B 0.035474f
C466 VTAIL.n3 B 0.024646f
C467 VTAIL.n4 B 0.013244f
C468 VTAIL.n5 B 0.031303f
C469 VTAIL.n6 B 0.014023f
C470 VTAIL.n7 B 0.024646f
C471 VTAIL.n8 B 0.013244f
C472 VTAIL.n9 B 0.031303f
C473 VTAIL.n10 B 0.014023f
C474 VTAIL.n11 B 0.024646f
C475 VTAIL.n12 B 0.013244f
C476 VTAIL.n13 B 0.031303f
C477 VTAIL.n14 B 0.014023f
C478 VTAIL.n15 B 0.024646f
C479 VTAIL.n16 B 0.013633f
C480 VTAIL.n17 B 0.031303f
C481 VTAIL.n18 B 0.014023f
C482 VTAIL.n19 B 0.024646f
C483 VTAIL.n20 B 0.013244f
C484 VTAIL.n21 B 0.031303f
C485 VTAIL.n22 B 0.014023f
C486 VTAIL.n23 B 0.024646f
C487 VTAIL.n24 B 0.013244f
C488 VTAIL.n25 B 0.023478f
C489 VTAIL.n26 B 0.022129f
C490 VTAIL.t17 B 0.053162f
C491 VTAIL.n27 B 0.198606f
C492 VTAIL.n28 B 1.48562f
C493 VTAIL.n29 B 0.013244f
C494 VTAIL.n30 B 0.014023f
C495 VTAIL.n31 B 0.031303f
C496 VTAIL.n32 B 0.031303f
C497 VTAIL.n33 B 0.014023f
C498 VTAIL.n34 B 0.013244f
C499 VTAIL.n35 B 0.024646f
C500 VTAIL.n36 B 0.024646f
C501 VTAIL.n37 B 0.013244f
C502 VTAIL.n38 B 0.014023f
C503 VTAIL.n39 B 0.031303f
C504 VTAIL.n40 B 0.031303f
C505 VTAIL.n41 B 0.014023f
C506 VTAIL.n42 B 0.013244f
C507 VTAIL.n43 B 0.024646f
C508 VTAIL.n44 B 0.024646f
C509 VTAIL.n45 B 0.013244f
C510 VTAIL.n46 B 0.013244f
C511 VTAIL.n47 B 0.014023f
C512 VTAIL.n48 B 0.031303f
C513 VTAIL.n49 B 0.031303f
C514 VTAIL.n50 B 0.031303f
C515 VTAIL.n51 B 0.013633f
C516 VTAIL.n52 B 0.013244f
C517 VTAIL.n53 B 0.024646f
C518 VTAIL.n54 B 0.024646f
C519 VTAIL.n55 B 0.013244f
C520 VTAIL.n56 B 0.014023f
C521 VTAIL.n57 B 0.031303f
C522 VTAIL.n58 B 0.031303f
C523 VTAIL.n59 B 0.014023f
C524 VTAIL.n60 B 0.013244f
C525 VTAIL.n61 B 0.024646f
C526 VTAIL.n62 B 0.024646f
C527 VTAIL.n63 B 0.013244f
C528 VTAIL.n64 B 0.014023f
C529 VTAIL.n65 B 0.031303f
C530 VTAIL.n66 B 0.031303f
C531 VTAIL.n67 B 0.014023f
C532 VTAIL.n68 B 0.013244f
C533 VTAIL.n69 B 0.024646f
C534 VTAIL.n70 B 0.024646f
C535 VTAIL.n71 B 0.013244f
C536 VTAIL.n72 B 0.014023f
C537 VTAIL.n73 B 0.031303f
C538 VTAIL.n74 B 0.069237f
C539 VTAIL.n75 B 0.014023f
C540 VTAIL.n76 B 0.013244f
C541 VTAIL.n77 B 0.054611f
C542 VTAIL.n78 B 0.038818f
C543 VTAIL.n79 B 0.395915f
C544 VTAIL.t12 B 0.276755f
C545 VTAIL.t19 B 0.276755f
C546 VTAIL.n80 B 2.40908f
C547 VTAIL.n81 B 0.705344f
C548 VTAIL.t11 B 0.276755f
C549 VTAIL.t13 B 0.276755f
C550 VTAIL.n82 B 2.40908f
C551 VTAIL.n83 B 2.23889f
C552 VTAIL.t8 B 0.276755f
C553 VTAIL.t5 B 0.276755f
C554 VTAIL.n84 B 2.40908f
C555 VTAIL.n85 B 2.23888f
C556 VTAIL.t0 B 0.276755f
C557 VTAIL.t1 B 0.276755f
C558 VTAIL.n86 B 2.40908f
C559 VTAIL.n87 B 0.70534f
C560 VTAIL.n88 B 0.035474f
C561 VTAIL.n89 B 0.024646f
C562 VTAIL.n90 B 0.013244f
C563 VTAIL.n91 B 0.031303f
C564 VTAIL.n92 B 0.014023f
C565 VTAIL.n93 B 0.024646f
C566 VTAIL.n94 B 0.013244f
C567 VTAIL.n95 B 0.031303f
C568 VTAIL.n96 B 0.014023f
C569 VTAIL.n97 B 0.024646f
C570 VTAIL.n98 B 0.013244f
C571 VTAIL.n99 B 0.031303f
C572 VTAIL.n100 B 0.014023f
C573 VTAIL.n101 B 0.024646f
C574 VTAIL.n102 B 0.013633f
C575 VTAIL.n103 B 0.031303f
C576 VTAIL.n104 B 0.013244f
C577 VTAIL.n105 B 0.014023f
C578 VTAIL.n106 B 0.024646f
C579 VTAIL.n107 B 0.013244f
C580 VTAIL.n108 B 0.031303f
C581 VTAIL.n109 B 0.014023f
C582 VTAIL.n110 B 0.024646f
C583 VTAIL.n111 B 0.013244f
C584 VTAIL.n112 B 0.023478f
C585 VTAIL.n113 B 0.022129f
C586 VTAIL.t7 B 0.053162f
C587 VTAIL.n114 B 0.198606f
C588 VTAIL.n115 B 1.48562f
C589 VTAIL.n116 B 0.013244f
C590 VTAIL.n117 B 0.014023f
C591 VTAIL.n118 B 0.031303f
C592 VTAIL.n119 B 0.031303f
C593 VTAIL.n120 B 0.014023f
C594 VTAIL.n121 B 0.013244f
C595 VTAIL.n122 B 0.024646f
C596 VTAIL.n123 B 0.024646f
C597 VTAIL.n124 B 0.013244f
C598 VTAIL.n125 B 0.014023f
C599 VTAIL.n126 B 0.031303f
C600 VTAIL.n127 B 0.031303f
C601 VTAIL.n128 B 0.014023f
C602 VTAIL.n129 B 0.013244f
C603 VTAIL.n130 B 0.024646f
C604 VTAIL.n131 B 0.024646f
C605 VTAIL.n132 B 0.013244f
C606 VTAIL.n133 B 0.014023f
C607 VTAIL.n134 B 0.031303f
C608 VTAIL.n135 B 0.031303f
C609 VTAIL.n136 B 0.031303f
C610 VTAIL.n137 B 0.013633f
C611 VTAIL.n138 B 0.013244f
C612 VTAIL.n139 B 0.024646f
C613 VTAIL.n140 B 0.024646f
C614 VTAIL.n141 B 0.013244f
C615 VTAIL.n142 B 0.014023f
C616 VTAIL.n143 B 0.031303f
C617 VTAIL.n144 B 0.031303f
C618 VTAIL.n145 B 0.014023f
C619 VTAIL.n146 B 0.013244f
C620 VTAIL.n147 B 0.024646f
C621 VTAIL.n148 B 0.024646f
C622 VTAIL.n149 B 0.013244f
C623 VTAIL.n150 B 0.014023f
C624 VTAIL.n151 B 0.031303f
C625 VTAIL.n152 B 0.031303f
C626 VTAIL.n153 B 0.014023f
C627 VTAIL.n154 B 0.013244f
C628 VTAIL.n155 B 0.024646f
C629 VTAIL.n156 B 0.024646f
C630 VTAIL.n157 B 0.013244f
C631 VTAIL.n158 B 0.014023f
C632 VTAIL.n159 B 0.031303f
C633 VTAIL.n160 B 0.069237f
C634 VTAIL.n161 B 0.014023f
C635 VTAIL.n162 B 0.013244f
C636 VTAIL.n163 B 0.054611f
C637 VTAIL.n164 B 0.038818f
C638 VTAIL.n165 B 0.395915f
C639 VTAIL.t10 B 0.276755f
C640 VTAIL.t14 B 0.276755f
C641 VTAIL.n166 B 2.40908f
C642 VTAIL.n167 B 0.62969f
C643 VTAIL.t16 B 0.276755f
C644 VTAIL.t15 B 0.276755f
C645 VTAIL.n168 B 2.40908f
C646 VTAIL.n169 B 0.70534f
C647 VTAIL.n170 B 0.035474f
C648 VTAIL.n171 B 0.024646f
C649 VTAIL.n172 B 0.013244f
C650 VTAIL.n173 B 0.031303f
C651 VTAIL.n174 B 0.014023f
C652 VTAIL.n175 B 0.024646f
C653 VTAIL.n176 B 0.013244f
C654 VTAIL.n177 B 0.031303f
C655 VTAIL.n178 B 0.014023f
C656 VTAIL.n179 B 0.024646f
C657 VTAIL.n180 B 0.013244f
C658 VTAIL.n181 B 0.031303f
C659 VTAIL.n182 B 0.014023f
C660 VTAIL.n183 B 0.024646f
C661 VTAIL.n184 B 0.013633f
C662 VTAIL.n185 B 0.031303f
C663 VTAIL.n186 B 0.013244f
C664 VTAIL.n187 B 0.014023f
C665 VTAIL.n188 B 0.024646f
C666 VTAIL.n189 B 0.013244f
C667 VTAIL.n190 B 0.031303f
C668 VTAIL.n191 B 0.014023f
C669 VTAIL.n192 B 0.024646f
C670 VTAIL.n193 B 0.013244f
C671 VTAIL.n194 B 0.023478f
C672 VTAIL.n195 B 0.022129f
C673 VTAIL.t18 B 0.053162f
C674 VTAIL.n196 B 0.198606f
C675 VTAIL.n197 B 1.48562f
C676 VTAIL.n198 B 0.013244f
C677 VTAIL.n199 B 0.014023f
C678 VTAIL.n200 B 0.031303f
C679 VTAIL.n201 B 0.031303f
C680 VTAIL.n202 B 0.014023f
C681 VTAIL.n203 B 0.013244f
C682 VTAIL.n204 B 0.024646f
C683 VTAIL.n205 B 0.024646f
C684 VTAIL.n206 B 0.013244f
C685 VTAIL.n207 B 0.014023f
C686 VTAIL.n208 B 0.031303f
C687 VTAIL.n209 B 0.031303f
C688 VTAIL.n210 B 0.014023f
C689 VTAIL.n211 B 0.013244f
C690 VTAIL.n212 B 0.024646f
C691 VTAIL.n213 B 0.024646f
C692 VTAIL.n214 B 0.013244f
C693 VTAIL.n215 B 0.014023f
C694 VTAIL.n216 B 0.031303f
C695 VTAIL.n217 B 0.031303f
C696 VTAIL.n218 B 0.031303f
C697 VTAIL.n219 B 0.013633f
C698 VTAIL.n220 B 0.013244f
C699 VTAIL.n221 B 0.024646f
C700 VTAIL.n222 B 0.024646f
C701 VTAIL.n223 B 0.013244f
C702 VTAIL.n224 B 0.014023f
C703 VTAIL.n225 B 0.031303f
C704 VTAIL.n226 B 0.031303f
C705 VTAIL.n227 B 0.014023f
C706 VTAIL.n228 B 0.013244f
C707 VTAIL.n229 B 0.024646f
C708 VTAIL.n230 B 0.024646f
C709 VTAIL.n231 B 0.013244f
C710 VTAIL.n232 B 0.014023f
C711 VTAIL.n233 B 0.031303f
C712 VTAIL.n234 B 0.031303f
C713 VTAIL.n235 B 0.014023f
C714 VTAIL.n236 B 0.013244f
C715 VTAIL.n237 B 0.024646f
C716 VTAIL.n238 B 0.024646f
C717 VTAIL.n239 B 0.013244f
C718 VTAIL.n240 B 0.014023f
C719 VTAIL.n241 B 0.031303f
C720 VTAIL.n242 B 0.069237f
C721 VTAIL.n243 B 0.014023f
C722 VTAIL.n244 B 0.013244f
C723 VTAIL.n245 B 0.054611f
C724 VTAIL.n246 B 0.038818f
C725 VTAIL.n247 B 1.77919f
C726 VTAIL.n248 B 0.035474f
C727 VTAIL.n249 B 0.024646f
C728 VTAIL.n250 B 0.013244f
C729 VTAIL.n251 B 0.031303f
C730 VTAIL.n252 B 0.014023f
C731 VTAIL.n253 B 0.024646f
C732 VTAIL.n254 B 0.013244f
C733 VTAIL.n255 B 0.031303f
C734 VTAIL.n256 B 0.014023f
C735 VTAIL.n257 B 0.024646f
C736 VTAIL.n258 B 0.013244f
C737 VTAIL.n259 B 0.031303f
C738 VTAIL.n260 B 0.014023f
C739 VTAIL.n261 B 0.024646f
C740 VTAIL.n262 B 0.013633f
C741 VTAIL.n263 B 0.031303f
C742 VTAIL.n264 B 0.014023f
C743 VTAIL.n265 B 0.024646f
C744 VTAIL.n266 B 0.013244f
C745 VTAIL.n267 B 0.031303f
C746 VTAIL.n268 B 0.014023f
C747 VTAIL.n269 B 0.024646f
C748 VTAIL.n270 B 0.013244f
C749 VTAIL.n271 B 0.023478f
C750 VTAIL.n272 B 0.022129f
C751 VTAIL.t9 B 0.053162f
C752 VTAIL.n273 B 0.198606f
C753 VTAIL.n274 B 1.48562f
C754 VTAIL.n275 B 0.013244f
C755 VTAIL.n276 B 0.014023f
C756 VTAIL.n277 B 0.031303f
C757 VTAIL.n278 B 0.031303f
C758 VTAIL.n279 B 0.014023f
C759 VTAIL.n280 B 0.013244f
C760 VTAIL.n281 B 0.024646f
C761 VTAIL.n282 B 0.024646f
C762 VTAIL.n283 B 0.013244f
C763 VTAIL.n284 B 0.014023f
C764 VTAIL.n285 B 0.031303f
C765 VTAIL.n286 B 0.031303f
C766 VTAIL.n287 B 0.014023f
C767 VTAIL.n288 B 0.013244f
C768 VTAIL.n289 B 0.024646f
C769 VTAIL.n290 B 0.024646f
C770 VTAIL.n291 B 0.013244f
C771 VTAIL.n292 B 0.013244f
C772 VTAIL.n293 B 0.014023f
C773 VTAIL.n294 B 0.031303f
C774 VTAIL.n295 B 0.031303f
C775 VTAIL.n296 B 0.031303f
C776 VTAIL.n297 B 0.013633f
C777 VTAIL.n298 B 0.013244f
C778 VTAIL.n299 B 0.024646f
C779 VTAIL.n300 B 0.024646f
C780 VTAIL.n301 B 0.013244f
C781 VTAIL.n302 B 0.014023f
C782 VTAIL.n303 B 0.031303f
C783 VTAIL.n304 B 0.031303f
C784 VTAIL.n305 B 0.014023f
C785 VTAIL.n306 B 0.013244f
C786 VTAIL.n307 B 0.024646f
C787 VTAIL.n308 B 0.024646f
C788 VTAIL.n309 B 0.013244f
C789 VTAIL.n310 B 0.014023f
C790 VTAIL.n311 B 0.031303f
C791 VTAIL.n312 B 0.031303f
C792 VTAIL.n313 B 0.014023f
C793 VTAIL.n314 B 0.013244f
C794 VTAIL.n315 B 0.024646f
C795 VTAIL.n316 B 0.024646f
C796 VTAIL.n317 B 0.013244f
C797 VTAIL.n318 B 0.014023f
C798 VTAIL.n319 B 0.031303f
C799 VTAIL.n320 B 0.069237f
C800 VTAIL.n321 B 0.014023f
C801 VTAIL.n322 B 0.013244f
C802 VTAIL.n323 B 0.054611f
C803 VTAIL.n324 B 0.038818f
C804 VTAIL.n325 B 1.77919f
C805 VTAIL.t2 B 0.276755f
C806 VTAIL.t3 B 0.276755f
C807 VTAIL.n326 B 2.40908f
C808 VTAIL.n327 B 0.531281f
C809 VP.t8 B 2.25904f
C810 VP.n0 B 0.861996f
C811 VP.n1 B 0.019559f
C812 VP.n2 B 0.025827f
C813 VP.n3 B 0.019559f
C814 VP.t1 B 2.25904f
C815 VP.n4 B 0.036453f
C816 VP.n5 B 0.019559f
C817 VP.n6 B 0.036453f
C818 VP.n7 B 0.019559f
C819 VP.t0 B 2.25904f
C820 VP.n8 B 0.035897f
C821 VP.n9 B 0.019559f
C822 VP.n10 B 0.020256f
C823 VP.n11 B 0.019559f
C824 VP.n12 B 0.031277f
C825 VP.n13 B 0.031567f
C826 VP.t3 B 2.25904f
C827 VP.t5 B 2.25904f
C828 VP.n14 B 0.861996f
C829 VP.n15 B 0.019559f
C830 VP.n16 B 0.025827f
C831 VP.n17 B 0.019559f
C832 VP.t7 B 2.25904f
C833 VP.n18 B 0.036453f
C834 VP.n19 B 0.019559f
C835 VP.n20 B 0.036453f
C836 VP.n21 B 0.019559f
C837 VP.t9 B 2.25904f
C838 VP.n22 B 0.035897f
C839 VP.n23 B 0.019559f
C840 VP.n24 B 0.020256f
C841 VP.t6 B 2.45585f
C842 VP.t4 B 2.25904f
C843 VP.n25 B 0.844138f
C844 VP.n26 B 0.821887f
C845 VP.n27 B 0.211597f
C846 VP.n28 B 0.019559f
C847 VP.n29 B 0.036453f
C848 VP.n30 B 0.039183f
C849 VP.n31 B 0.018477f
C850 VP.n32 B 0.019559f
C851 VP.n33 B 0.019559f
C852 VP.n34 B 0.019559f
C853 VP.n35 B 0.036453f
C854 VP.n36 B 0.027454f
C855 VP.n37 B 0.789099f
C856 VP.n38 B 0.027454f
C857 VP.n39 B 0.019559f
C858 VP.n40 B 0.019559f
C859 VP.n41 B 0.019559f
C860 VP.n42 B 0.035897f
C861 VP.n43 B 0.018477f
C862 VP.n44 B 0.039183f
C863 VP.n45 B 0.019559f
C864 VP.n46 B 0.019559f
C865 VP.n47 B 0.019559f
C866 VP.n48 B 0.020256f
C867 VP.n49 B 0.789099f
C868 VP.n50 B 0.034653f
C869 VP.n51 B 0.036453f
C870 VP.n52 B 0.019559f
C871 VP.n53 B 0.019559f
C872 VP.n54 B 0.019559f
C873 VP.n55 B 0.031277f
C874 VP.n56 B 0.036453f
C875 VP.n57 B 0.031054f
C876 VP.n58 B 0.031567f
C877 VP.n59 B 1.3263f
C878 VP.n60 B 1.33867f
C879 VP.n61 B 0.861996f
C880 VP.n62 B 0.031054f
C881 VP.n63 B 0.036453f
C882 VP.n64 B 0.019559f
C883 VP.n65 B 0.019559f
C884 VP.n66 B 0.019559f
C885 VP.n67 B 0.025827f
C886 VP.n68 B 0.036453f
C887 VP.t2 B 2.25904f
C888 VP.n69 B 0.789099f
C889 VP.n70 B 0.034653f
C890 VP.n71 B 0.019559f
C891 VP.n72 B 0.019559f
C892 VP.n73 B 0.019559f
C893 VP.n74 B 0.036453f
C894 VP.n75 B 0.039183f
C895 VP.n76 B 0.018477f
C896 VP.n77 B 0.019559f
C897 VP.n78 B 0.019559f
C898 VP.n79 B 0.019559f
C899 VP.n80 B 0.036453f
C900 VP.n81 B 0.027454f
C901 VP.n82 B 0.789099f
C902 VP.n83 B 0.027454f
C903 VP.n84 B 0.019559f
C904 VP.n85 B 0.019559f
C905 VP.n86 B 0.019559f
C906 VP.n87 B 0.035897f
C907 VP.n88 B 0.018477f
C908 VP.n89 B 0.039183f
C909 VP.n90 B 0.019559f
C910 VP.n91 B 0.019559f
C911 VP.n92 B 0.019559f
C912 VP.n93 B 0.020256f
C913 VP.n94 B 0.789099f
C914 VP.n95 B 0.034653f
C915 VP.n96 B 0.036453f
C916 VP.n97 B 0.019559f
C917 VP.n98 B 0.019559f
C918 VP.n99 B 0.019559f
C919 VP.n100 B 0.031277f
C920 VP.n101 B 0.036453f
C921 VP.n102 B 0.031054f
C922 VP.n103 B 0.031567f
C923 VP.n104 B 0.042881f
.ends

