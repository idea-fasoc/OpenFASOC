* NGSPICE file created from diff_pair_sample_0486.ext - technology: sky130A

.subckt diff_pair_sample_0486 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t11 VP.t0 VDD1.t5 w_n3898_n1280# sky130_fd_pr__pfet_01v8 ad=0.2574 pd=1.89 as=0.2574 ps=1.89 w=1.56 l=3.33
X1 B.t11 B.t9 B.t10 w_n3898_n1280# sky130_fd_pr__pfet_01v8 ad=0.6084 pd=3.9 as=0 ps=0 w=1.56 l=3.33
X2 VDD1.t0 VP.t1 VTAIL.t10 w_n3898_n1280# sky130_fd_pr__pfet_01v8 ad=0.2574 pd=1.89 as=0.6084 ps=3.9 w=1.56 l=3.33
X3 VTAIL.t2 VN.t0 VDD2.t5 w_n3898_n1280# sky130_fd_pr__pfet_01v8 ad=0.2574 pd=1.89 as=0.2574 ps=1.89 w=1.56 l=3.33
X4 VDD2.t4 VN.t1 VTAIL.t4 w_n3898_n1280# sky130_fd_pr__pfet_01v8 ad=0.6084 pd=3.9 as=0.2574 ps=1.89 w=1.56 l=3.33
X5 VDD1.t2 VP.t2 VTAIL.t9 w_n3898_n1280# sky130_fd_pr__pfet_01v8 ad=0.6084 pd=3.9 as=0.2574 ps=1.89 w=1.56 l=3.33
X6 B.t8 B.t6 B.t7 w_n3898_n1280# sky130_fd_pr__pfet_01v8 ad=0.6084 pd=3.9 as=0 ps=0 w=1.56 l=3.33
X7 VDD2.t3 VN.t2 VTAIL.t5 w_n3898_n1280# sky130_fd_pr__pfet_01v8 ad=0.2574 pd=1.89 as=0.6084 ps=3.9 w=1.56 l=3.33
X8 B.t5 B.t3 B.t4 w_n3898_n1280# sky130_fd_pr__pfet_01v8 ad=0.6084 pd=3.9 as=0 ps=0 w=1.56 l=3.33
X9 VDD1.t1 VP.t3 VTAIL.t8 w_n3898_n1280# sky130_fd_pr__pfet_01v8 ad=0.6084 pd=3.9 as=0.2574 ps=1.89 w=1.56 l=3.33
X10 VTAIL.t7 VP.t4 VDD1.t3 w_n3898_n1280# sky130_fd_pr__pfet_01v8 ad=0.2574 pd=1.89 as=0.2574 ps=1.89 w=1.56 l=3.33
X11 VDD2.t2 VN.t3 VTAIL.t1 w_n3898_n1280# sky130_fd_pr__pfet_01v8 ad=0.2574 pd=1.89 as=0.6084 ps=3.9 w=1.56 l=3.33
X12 VDD2.t1 VN.t4 VTAIL.t3 w_n3898_n1280# sky130_fd_pr__pfet_01v8 ad=0.6084 pd=3.9 as=0.2574 ps=1.89 w=1.56 l=3.33
X13 VTAIL.t0 VN.t5 VDD2.t0 w_n3898_n1280# sky130_fd_pr__pfet_01v8 ad=0.2574 pd=1.89 as=0.2574 ps=1.89 w=1.56 l=3.33
X14 VDD1.t4 VP.t5 VTAIL.t6 w_n3898_n1280# sky130_fd_pr__pfet_01v8 ad=0.2574 pd=1.89 as=0.6084 ps=3.9 w=1.56 l=3.33
X15 B.t2 B.t0 B.t1 w_n3898_n1280# sky130_fd_pr__pfet_01v8 ad=0.6084 pd=3.9 as=0 ps=0 w=1.56 l=3.33
R0 VP.n16 VP.n15 161.3
R1 VP.n17 VP.n12 161.3
R2 VP.n19 VP.n18 161.3
R3 VP.n20 VP.n11 161.3
R4 VP.n22 VP.n21 161.3
R5 VP.n23 VP.n10 161.3
R6 VP.n25 VP.n24 161.3
R7 VP.n50 VP.n49 161.3
R8 VP.n48 VP.n1 161.3
R9 VP.n47 VP.n46 161.3
R10 VP.n45 VP.n2 161.3
R11 VP.n44 VP.n43 161.3
R12 VP.n42 VP.n3 161.3
R13 VP.n41 VP.n40 161.3
R14 VP.n39 VP.n4 161.3
R15 VP.n38 VP.n37 161.3
R16 VP.n36 VP.n5 161.3
R17 VP.n35 VP.n34 161.3
R18 VP.n33 VP.n6 161.3
R19 VP.n32 VP.n31 161.3
R20 VP.n30 VP.n7 161.3
R21 VP.n29 VP.n28 161.3
R22 VP.n27 VP.n8 82.1011
R23 VP.n51 VP.n0 82.1011
R24 VP.n26 VP.n9 82.1011
R25 VP.n35 VP.n6 56.4773
R26 VP.n43 VP.n2 56.4773
R27 VP.n18 VP.n11 56.4773
R28 VP.n14 VP.n13 49.9597
R29 VP.n14 VP.t2 44.2305
R30 VP.n27 VP.n26 43.6431
R31 VP.n30 VP.n29 24.3439
R32 VP.n31 VP.n30 24.3439
R33 VP.n31 VP.n6 24.3439
R34 VP.n36 VP.n35 24.3439
R35 VP.n37 VP.n36 24.3439
R36 VP.n37 VP.n4 24.3439
R37 VP.n41 VP.n4 24.3439
R38 VP.n42 VP.n41 24.3439
R39 VP.n43 VP.n42 24.3439
R40 VP.n47 VP.n2 24.3439
R41 VP.n48 VP.n47 24.3439
R42 VP.n49 VP.n48 24.3439
R43 VP.n22 VP.n11 24.3439
R44 VP.n23 VP.n22 24.3439
R45 VP.n24 VP.n23 24.3439
R46 VP.n16 VP.n13 24.3439
R47 VP.n17 VP.n16 24.3439
R48 VP.n18 VP.n17 24.3439
R49 VP.n4 VP.t0 11.2906
R50 VP.n8 VP.t3 11.2906
R51 VP.n0 VP.t1 11.2906
R52 VP.n13 VP.t4 11.2906
R53 VP.n9 VP.t5 11.2906
R54 VP.n29 VP.n8 7.7904
R55 VP.n49 VP.n0 7.7904
R56 VP.n24 VP.n9 7.7904
R57 VP.n15 VP.n14 3.24065
R58 VP.n26 VP.n25 0.355081
R59 VP.n28 VP.n27 0.355081
R60 VP.n51 VP.n50 0.355081
R61 VP VP.n51 0.26685
R62 VP.n15 VP.n12 0.189894
R63 VP.n19 VP.n12 0.189894
R64 VP.n20 VP.n19 0.189894
R65 VP.n21 VP.n20 0.189894
R66 VP.n21 VP.n10 0.189894
R67 VP.n25 VP.n10 0.189894
R68 VP.n28 VP.n7 0.189894
R69 VP.n32 VP.n7 0.189894
R70 VP.n33 VP.n32 0.189894
R71 VP.n34 VP.n33 0.189894
R72 VP.n34 VP.n5 0.189894
R73 VP.n38 VP.n5 0.189894
R74 VP.n39 VP.n38 0.189894
R75 VP.n40 VP.n39 0.189894
R76 VP.n40 VP.n3 0.189894
R77 VP.n44 VP.n3 0.189894
R78 VP.n45 VP.n44 0.189894
R79 VP.n46 VP.n45 0.189894
R80 VP.n46 VP.n1 0.189894
R81 VP.n50 VP.n1 0.189894
R82 VDD1 VDD1.t2 271.046
R83 VDD1.n1 VDD1.t1 270.932
R84 VDD1.n1 VDD1.n0 248.518
R85 VDD1.n3 VDD1.n2 247.785
R86 VDD1.n3 VDD1.n1 37.475
R87 VDD1.n2 VDD1.t3 20.837
R88 VDD1.n2 VDD1.t4 20.837
R89 VDD1.n0 VDD1.t5 20.837
R90 VDD1.n0 VDD1.t0 20.837
R91 VDD1 VDD1.n3 0.731103
R92 VTAIL.n10 VTAIL.t6 251.942
R93 VTAIL.n7 VTAIL.t5 251.942
R94 VTAIL.n11 VTAIL.t1 251.942
R95 VTAIL.n2 VTAIL.t10 251.942
R96 VTAIL.n1 VTAIL.n0 231.106
R97 VTAIL.n4 VTAIL.n3 231.106
R98 VTAIL.n9 VTAIL.n8 231.106
R99 VTAIL.n6 VTAIL.n5 231.106
R100 VTAIL.n0 VTAIL.t4 20.837
R101 VTAIL.n0 VTAIL.t2 20.837
R102 VTAIL.n3 VTAIL.t8 20.837
R103 VTAIL.n3 VTAIL.t11 20.837
R104 VTAIL.n8 VTAIL.t9 20.837
R105 VTAIL.n8 VTAIL.t7 20.837
R106 VTAIL.n5 VTAIL.t3 20.837
R107 VTAIL.n5 VTAIL.t0 20.837
R108 VTAIL.n6 VTAIL.n4 20.0221
R109 VTAIL.n11 VTAIL.n10 16.8669
R110 VTAIL.n7 VTAIL.n6 3.15567
R111 VTAIL.n10 VTAIL.n9 3.15567
R112 VTAIL.n4 VTAIL.n2 3.15567
R113 VTAIL VTAIL.n11 2.30869
R114 VTAIL.n9 VTAIL.n7 2.04791
R115 VTAIL.n2 VTAIL.n1 2.04791
R116 VTAIL VTAIL.n1 0.847483
R117 B.n422 B.n421 585
R118 B.n423 B.n46 585
R119 B.n425 B.n424 585
R120 B.n426 B.n45 585
R121 B.n428 B.n427 585
R122 B.n429 B.n44 585
R123 B.n431 B.n430 585
R124 B.n432 B.n43 585
R125 B.n434 B.n433 585
R126 B.n435 B.n42 585
R127 B.n437 B.n436 585
R128 B.n439 B.n39 585
R129 B.n441 B.n440 585
R130 B.n442 B.n38 585
R131 B.n444 B.n443 585
R132 B.n445 B.n37 585
R133 B.n447 B.n446 585
R134 B.n448 B.n36 585
R135 B.n450 B.n449 585
R136 B.n451 B.n33 585
R137 B.n454 B.n453 585
R138 B.n455 B.n32 585
R139 B.n457 B.n456 585
R140 B.n458 B.n31 585
R141 B.n460 B.n459 585
R142 B.n461 B.n30 585
R143 B.n463 B.n462 585
R144 B.n464 B.n29 585
R145 B.n466 B.n465 585
R146 B.n467 B.n28 585
R147 B.n469 B.n468 585
R148 B.n420 B.n47 585
R149 B.n419 B.n418 585
R150 B.n417 B.n48 585
R151 B.n416 B.n415 585
R152 B.n414 B.n49 585
R153 B.n413 B.n412 585
R154 B.n411 B.n50 585
R155 B.n410 B.n409 585
R156 B.n408 B.n51 585
R157 B.n407 B.n406 585
R158 B.n405 B.n52 585
R159 B.n404 B.n403 585
R160 B.n402 B.n53 585
R161 B.n401 B.n400 585
R162 B.n399 B.n54 585
R163 B.n398 B.n397 585
R164 B.n396 B.n55 585
R165 B.n395 B.n394 585
R166 B.n393 B.n56 585
R167 B.n392 B.n391 585
R168 B.n390 B.n57 585
R169 B.n389 B.n388 585
R170 B.n387 B.n58 585
R171 B.n386 B.n385 585
R172 B.n384 B.n59 585
R173 B.n383 B.n382 585
R174 B.n381 B.n60 585
R175 B.n380 B.n379 585
R176 B.n378 B.n61 585
R177 B.n377 B.n376 585
R178 B.n375 B.n62 585
R179 B.n374 B.n373 585
R180 B.n372 B.n63 585
R181 B.n371 B.n370 585
R182 B.n369 B.n64 585
R183 B.n368 B.n367 585
R184 B.n366 B.n65 585
R185 B.n365 B.n364 585
R186 B.n363 B.n66 585
R187 B.n362 B.n361 585
R188 B.n360 B.n67 585
R189 B.n359 B.n358 585
R190 B.n357 B.n68 585
R191 B.n356 B.n355 585
R192 B.n354 B.n69 585
R193 B.n353 B.n352 585
R194 B.n351 B.n70 585
R195 B.n350 B.n349 585
R196 B.n348 B.n71 585
R197 B.n347 B.n346 585
R198 B.n345 B.n72 585
R199 B.n344 B.n343 585
R200 B.n342 B.n73 585
R201 B.n341 B.n340 585
R202 B.n339 B.n74 585
R203 B.n338 B.n337 585
R204 B.n336 B.n75 585
R205 B.n335 B.n334 585
R206 B.n333 B.n76 585
R207 B.n332 B.n331 585
R208 B.n330 B.n77 585
R209 B.n329 B.n328 585
R210 B.n327 B.n78 585
R211 B.n326 B.n325 585
R212 B.n324 B.n79 585
R213 B.n323 B.n322 585
R214 B.n321 B.n80 585
R215 B.n320 B.n319 585
R216 B.n318 B.n81 585
R217 B.n317 B.n316 585
R218 B.n315 B.n82 585
R219 B.n314 B.n313 585
R220 B.n312 B.n83 585
R221 B.n311 B.n310 585
R222 B.n309 B.n84 585
R223 B.n308 B.n307 585
R224 B.n306 B.n85 585
R225 B.n305 B.n304 585
R226 B.n303 B.n86 585
R227 B.n302 B.n301 585
R228 B.n300 B.n87 585
R229 B.n299 B.n298 585
R230 B.n297 B.n88 585
R231 B.n296 B.n295 585
R232 B.n294 B.n89 585
R233 B.n293 B.n292 585
R234 B.n291 B.n90 585
R235 B.n290 B.n289 585
R236 B.n288 B.n91 585
R237 B.n287 B.n286 585
R238 B.n285 B.n92 585
R239 B.n284 B.n283 585
R240 B.n282 B.n93 585
R241 B.n281 B.n280 585
R242 B.n279 B.n94 585
R243 B.n278 B.n277 585
R244 B.n276 B.n95 585
R245 B.n275 B.n274 585
R246 B.n273 B.n96 585
R247 B.n272 B.n271 585
R248 B.n270 B.n97 585
R249 B.n269 B.n268 585
R250 B.n267 B.n98 585
R251 B.n219 B.n118 585
R252 B.n221 B.n220 585
R253 B.n222 B.n117 585
R254 B.n224 B.n223 585
R255 B.n225 B.n116 585
R256 B.n227 B.n226 585
R257 B.n228 B.n115 585
R258 B.n230 B.n229 585
R259 B.n231 B.n114 585
R260 B.n233 B.n232 585
R261 B.n234 B.n111 585
R262 B.n237 B.n236 585
R263 B.n238 B.n110 585
R264 B.n240 B.n239 585
R265 B.n241 B.n109 585
R266 B.n243 B.n242 585
R267 B.n244 B.n108 585
R268 B.n246 B.n245 585
R269 B.n247 B.n107 585
R270 B.n249 B.n248 585
R271 B.n251 B.n250 585
R272 B.n252 B.n103 585
R273 B.n254 B.n253 585
R274 B.n255 B.n102 585
R275 B.n257 B.n256 585
R276 B.n258 B.n101 585
R277 B.n260 B.n259 585
R278 B.n261 B.n100 585
R279 B.n263 B.n262 585
R280 B.n264 B.n99 585
R281 B.n266 B.n265 585
R282 B.n218 B.n217 585
R283 B.n216 B.n119 585
R284 B.n215 B.n214 585
R285 B.n213 B.n120 585
R286 B.n212 B.n211 585
R287 B.n210 B.n121 585
R288 B.n209 B.n208 585
R289 B.n207 B.n122 585
R290 B.n206 B.n205 585
R291 B.n204 B.n123 585
R292 B.n203 B.n202 585
R293 B.n201 B.n124 585
R294 B.n200 B.n199 585
R295 B.n198 B.n125 585
R296 B.n197 B.n196 585
R297 B.n195 B.n126 585
R298 B.n194 B.n193 585
R299 B.n192 B.n127 585
R300 B.n191 B.n190 585
R301 B.n189 B.n128 585
R302 B.n188 B.n187 585
R303 B.n186 B.n129 585
R304 B.n185 B.n184 585
R305 B.n183 B.n130 585
R306 B.n182 B.n181 585
R307 B.n180 B.n131 585
R308 B.n179 B.n178 585
R309 B.n177 B.n132 585
R310 B.n176 B.n175 585
R311 B.n174 B.n133 585
R312 B.n173 B.n172 585
R313 B.n171 B.n134 585
R314 B.n170 B.n169 585
R315 B.n168 B.n135 585
R316 B.n167 B.n166 585
R317 B.n165 B.n136 585
R318 B.n164 B.n163 585
R319 B.n162 B.n137 585
R320 B.n161 B.n160 585
R321 B.n159 B.n138 585
R322 B.n158 B.n157 585
R323 B.n156 B.n139 585
R324 B.n155 B.n154 585
R325 B.n153 B.n140 585
R326 B.n152 B.n151 585
R327 B.n150 B.n141 585
R328 B.n149 B.n148 585
R329 B.n147 B.n142 585
R330 B.n146 B.n145 585
R331 B.n144 B.n143 585
R332 B.n2 B.n0 585
R333 B.n545 B.n1 585
R334 B.n544 B.n543 585
R335 B.n542 B.n3 585
R336 B.n541 B.n540 585
R337 B.n539 B.n4 585
R338 B.n538 B.n537 585
R339 B.n536 B.n5 585
R340 B.n535 B.n534 585
R341 B.n533 B.n6 585
R342 B.n532 B.n531 585
R343 B.n530 B.n7 585
R344 B.n529 B.n528 585
R345 B.n527 B.n8 585
R346 B.n526 B.n525 585
R347 B.n524 B.n9 585
R348 B.n523 B.n522 585
R349 B.n521 B.n10 585
R350 B.n520 B.n519 585
R351 B.n518 B.n11 585
R352 B.n517 B.n516 585
R353 B.n515 B.n12 585
R354 B.n514 B.n513 585
R355 B.n512 B.n13 585
R356 B.n511 B.n510 585
R357 B.n509 B.n14 585
R358 B.n508 B.n507 585
R359 B.n506 B.n15 585
R360 B.n505 B.n504 585
R361 B.n503 B.n16 585
R362 B.n502 B.n501 585
R363 B.n500 B.n17 585
R364 B.n499 B.n498 585
R365 B.n497 B.n18 585
R366 B.n496 B.n495 585
R367 B.n494 B.n19 585
R368 B.n493 B.n492 585
R369 B.n491 B.n20 585
R370 B.n490 B.n489 585
R371 B.n488 B.n21 585
R372 B.n487 B.n486 585
R373 B.n485 B.n22 585
R374 B.n484 B.n483 585
R375 B.n482 B.n23 585
R376 B.n481 B.n480 585
R377 B.n479 B.n24 585
R378 B.n478 B.n477 585
R379 B.n476 B.n25 585
R380 B.n475 B.n474 585
R381 B.n473 B.n26 585
R382 B.n472 B.n471 585
R383 B.n470 B.n27 585
R384 B.n547 B.n546 585
R385 B.n219 B.n218 559.769
R386 B.n468 B.n27 559.769
R387 B.n267 B.n266 559.769
R388 B.n422 B.n47 559.769
R389 B.n104 B.t8 320.76
R390 B.n40 B.t10 320.76
R391 B.n112 B.t5 320.76
R392 B.n34 B.t1 320.76
R393 B.n105 B.t7 249.778
R394 B.n41 B.t11 249.778
R395 B.n113 B.t4 249.778
R396 B.n35 B.t2 249.778
R397 B.n104 B.t6 209.431
R398 B.n112 B.t3 209.431
R399 B.n34 B.t0 209.431
R400 B.n40 B.t9 209.431
R401 B.n218 B.n119 163.367
R402 B.n214 B.n119 163.367
R403 B.n214 B.n213 163.367
R404 B.n213 B.n212 163.367
R405 B.n212 B.n121 163.367
R406 B.n208 B.n121 163.367
R407 B.n208 B.n207 163.367
R408 B.n207 B.n206 163.367
R409 B.n206 B.n123 163.367
R410 B.n202 B.n123 163.367
R411 B.n202 B.n201 163.367
R412 B.n201 B.n200 163.367
R413 B.n200 B.n125 163.367
R414 B.n196 B.n125 163.367
R415 B.n196 B.n195 163.367
R416 B.n195 B.n194 163.367
R417 B.n194 B.n127 163.367
R418 B.n190 B.n127 163.367
R419 B.n190 B.n189 163.367
R420 B.n189 B.n188 163.367
R421 B.n188 B.n129 163.367
R422 B.n184 B.n129 163.367
R423 B.n184 B.n183 163.367
R424 B.n183 B.n182 163.367
R425 B.n182 B.n131 163.367
R426 B.n178 B.n131 163.367
R427 B.n178 B.n177 163.367
R428 B.n177 B.n176 163.367
R429 B.n176 B.n133 163.367
R430 B.n172 B.n133 163.367
R431 B.n172 B.n171 163.367
R432 B.n171 B.n170 163.367
R433 B.n170 B.n135 163.367
R434 B.n166 B.n135 163.367
R435 B.n166 B.n165 163.367
R436 B.n165 B.n164 163.367
R437 B.n164 B.n137 163.367
R438 B.n160 B.n137 163.367
R439 B.n160 B.n159 163.367
R440 B.n159 B.n158 163.367
R441 B.n158 B.n139 163.367
R442 B.n154 B.n139 163.367
R443 B.n154 B.n153 163.367
R444 B.n153 B.n152 163.367
R445 B.n152 B.n141 163.367
R446 B.n148 B.n141 163.367
R447 B.n148 B.n147 163.367
R448 B.n147 B.n146 163.367
R449 B.n146 B.n143 163.367
R450 B.n143 B.n2 163.367
R451 B.n546 B.n2 163.367
R452 B.n546 B.n545 163.367
R453 B.n545 B.n544 163.367
R454 B.n544 B.n3 163.367
R455 B.n540 B.n3 163.367
R456 B.n540 B.n539 163.367
R457 B.n539 B.n538 163.367
R458 B.n538 B.n5 163.367
R459 B.n534 B.n5 163.367
R460 B.n534 B.n533 163.367
R461 B.n533 B.n532 163.367
R462 B.n532 B.n7 163.367
R463 B.n528 B.n7 163.367
R464 B.n528 B.n527 163.367
R465 B.n527 B.n526 163.367
R466 B.n526 B.n9 163.367
R467 B.n522 B.n9 163.367
R468 B.n522 B.n521 163.367
R469 B.n521 B.n520 163.367
R470 B.n520 B.n11 163.367
R471 B.n516 B.n11 163.367
R472 B.n516 B.n515 163.367
R473 B.n515 B.n514 163.367
R474 B.n514 B.n13 163.367
R475 B.n510 B.n13 163.367
R476 B.n510 B.n509 163.367
R477 B.n509 B.n508 163.367
R478 B.n508 B.n15 163.367
R479 B.n504 B.n15 163.367
R480 B.n504 B.n503 163.367
R481 B.n503 B.n502 163.367
R482 B.n502 B.n17 163.367
R483 B.n498 B.n17 163.367
R484 B.n498 B.n497 163.367
R485 B.n497 B.n496 163.367
R486 B.n496 B.n19 163.367
R487 B.n492 B.n19 163.367
R488 B.n492 B.n491 163.367
R489 B.n491 B.n490 163.367
R490 B.n490 B.n21 163.367
R491 B.n486 B.n21 163.367
R492 B.n486 B.n485 163.367
R493 B.n485 B.n484 163.367
R494 B.n484 B.n23 163.367
R495 B.n480 B.n23 163.367
R496 B.n480 B.n479 163.367
R497 B.n479 B.n478 163.367
R498 B.n478 B.n25 163.367
R499 B.n474 B.n25 163.367
R500 B.n474 B.n473 163.367
R501 B.n473 B.n472 163.367
R502 B.n472 B.n27 163.367
R503 B.n220 B.n219 163.367
R504 B.n220 B.n117 163.367
R505 B.n224 B.n117 163.367
R506 B.n225 B.n224 163.367
R507 B.n226 B.n225 163.367
R508 B.n226 B.n115 163.367
R509 B.n230 B.n115 163.367
R510 B.n231 B.n230 163.367
R511 B.n232 B.n231 163.367
R512 B.n232 B.n111 163.367
R513 B.n237 B.n111 163.367
R514 B.n238 B.n237 163.367
R515 B.n239 B.n238 163.367
R516 B.n239 B.n109 163.367
R517 B.n243 B.n109 163.367
R518 B.n244 B.n243 163.367
R519 B.n245 B.n244 163.367
R520 B.n245 B.n107 163.367
R521 B.n249 B.n107 163.367
R522 B.n250 B.n249 163.367
R523 B.n250 B.n103 163.367
R524 B.n254 B.n103 163.367
R525 B.n255 B.n254 163.367
R526 B.n256 B.n255 163.367
R527 B.n256 B.n101 163.367
R528 B.n260 B.n101 163.367
R529 B.n261 B.n260 163.367
R530 B.n262 B.n261 163.367
R531 B.n262 B.n99 163.367
R532 B.n266 B.n99 163.367
R533 B.n268 B.n267 163.367
R534 B.n268 B.n97 163.367
R535 B.n272 B.n97 163.367
R536 B.n273 B.n272 163.367
R537 B.n274 B.n273 163.367
R538 B.n274 B.n95 163.367
R539 B.n278 B.n95 163.367
R540 B.n279 B.n278 163.367
R541 B.n280 B.n279 163.367
R542 B.n280 B.n93 163.367
R543 B.n284 B.n93 163.367
R544 B.n285 B.n284 163.367
R545 B.n286 B.n285 163.367
R546 B.n286 B.n91 163.367
R547 B.n290 B.n91 163.367
R548 B.n291 B.n290 163.367
R549 B.n292 B.n291 163.367
R550 B.n292 B.n89 163.367
R551 B.n296 B.n89 163.367
R552 B.n297 B.n296 163.367
R553 B.n298 B.n297 163.367
R554 B.n298 B.n87 163.367
R555 B.n302 B.n87 163.367
R556 B.n303 B.n302 163.367
R557 B.n304 B.n303 163.367
R558 B.n304 B.n85 163.367
R559 B.n308 B.n85 163.367
R560 B.n309 B.n308 163.367
R561 B.n310 B.n309 163.367
R562 B.n310 B.n83 163.367
R563 B.n314 B.n83 163.367
R564 B.n315 B.n314 163.367
R565 B.n316 B.n315 163.367
R566 B.n316 B.n81 163.367
R567 B.n320 B.n81 163.367
R568 B.n321 B.n320 163.367
R569 B.n322 B.n321 163.367
R570 B.n322 B.n79 163.367
R571 B.n326 B.n79 163.367
R572 B.n327 B.n326 163.367
R573 B.n328 B.n327 163.367
R574 B.n328 B.n77 163.367
R575 B.n332 B.n77 163.367
R576 B.n333 B.n332 163.367
R577 B.n334 B.n333 163.367
R578 B.n334 B.n75 163.367
R579 B.n338 B.n75 163.367
R580 B.n339 B.n338 163.367
R581 B.n340 B.n339 163.367
R582 B.n340 B.n73 163.367
R583 B.n344 B.n73 163.367
R584 B.n345 B.n344 163.367
R585 B.n346 B.n345 163.367
R586 B.n346 B.n71 163.367
R587 B.n350 B.n71 163.367
R588 B.n351 B.n350 163.367
R589 B.n352 B.n351 163.367
R590 B.n352 B.n69 163.367
R591 B.n356 B.n69 163.367
R592 B.n357 B.n356 163.367
R593 B.n358 B.n357 163.367
R594 B.n358 B.n67 163.367
R595 B.n362 B.n67 163.367
R596 B.n363 B.n362 163.367
R597 B.n364 B.n363 163.367
R598 B.n364 B.n65 163.367
R599 B.n368 B.n65 163.367
R600 B.n369 B.n368 163.367
R601 B.n370 B.n369 163.367
R602 B.n370 B.n63 163.367
R603 B.n374 B.n63 163.367
R604 B.n375 B.n374 163.367
R605 B.n376 B.n375 163.367
R606 B.n376 B.n61 163.367
R607 B.n380 B.n61 163.367
R608 B.n381 B.n380 163.367
R609 B.n382 B.n381 163.367
R610 B.n382 B.n59 163.367
R611 B.n386 B.n59 163.367
R612 B.n387 B.n386 163.367
R613 B.n388 B.n387 163.367
R614 B.n388 B.n57 163.367
R615 B.n392 B.n57 163.367
R616 B.n393 B.n392 163.367
R617 B.n394 B.n393 163.367
R618 B.n394 B.n55 163.367
R619 B.n398 B.n55 163.367
R620 B.n399 B.n398 163.367
R621 B.n400 B.n399 163.367
R622 B.n400 B.n53 163.367
R623 B.n404 B.n53 163.367
R624 B.n405 B.n404 163.367
R625 B.n406 B.n405 163.367
R626 B.n406 B.n51 163.367
R627 B.n410 B.n51 163.367
R628 B.n411 B.n410 163.367
R629 B.n412 B.n411 163.367
R630 B.n412 B.n49 163.367
R631 B.n416 B.n49 163.367
R632 B.n417 B.n416 163.367
R633 B.n418 B.n417 163.367
R634 B.n418 B.n47 163.367
R635 B.n468 B.n467 163.367
R636 B.n467 B.n466 163.367
R637 B.n466 B.n29 163.367
R638 B.n462 B.n29 163.367
R639 B.n462 B.n461 163.367
R640 B.n461 B.n460 163.367
R641 B.n460 B.n31 163.367
R642 B.n456 B.n31 163.367
R643 B.n456 B.n455 163.367
R644 B.n455 B.n454 163.367
R645 B.n454 B.n33 163.367
R646 B.n449 B.n33 163.367
R647 B.n449 B.n448 163.367
R648 B.n448 B.n447 163.367
R649 B.n447 B.n37 163.367
R650 B.n443 B.n37 163.367
R651 B.n443 B.n442 163.367
R652 B.n442 B.n441 163.367
R653 B.n441 B.n39 163.367
R654 B.n436 B.n39 163.367
R655 B.n436 B.n435 163.367
R656 B.n435 B.n434 163.367
R657 B.n434 B.n43 163.367
R658 B.n430 B.n43 163.367
R659 B.n430 B.n429 163.367
R660 B.n429 B.n428 163.367
R661 B.n428 B.n45 163.367
R662 B.n424 B.n45 163.367
R663 B.n424 B.n423 163.367
R664 B.n423 B.n422 163.367
R665 B.n105 B.n104 70.9823
R666 B.n113 B.n112 70.9823
R667 B.n35 B.n34 70.9823
R668 B.n41 B.n40 70.9823
R669 B.n106 B.n105 59.5399
R670 B.n235 B.n113 59.5399
R671 B.n452 B.n35 59.5399
R672 B.n438 B.n41 59.5399
R673 B.n470 B.n469 36.3712
R674 B.n421 B.n420 36.3712
R675 B.n265 B.n98 36.3712
R676 B.n217 B.n118 36.3712
R677 B B.n547 18.0485
R678 B.n469 B.n28 10.6151
R679 B.n465 B.n28 10.6151
R680 B.n465 B.n464 10.6151
R681 B.n464 B.n463 10.6151
R682 B.n463 B.n30 10.6151
R683 B.n459 B.n30 10.6151
R684 B.n459 B.n458 10.6151
R685 B.n458 B.n457 10.6151
R686 B.n457 B.n32 10.6151
R687 B.n453 B.n32 10.6151
R688 B.n451 B.n450 10.6151
R689 B.n450 B.n36 10.6151
R690 B.n446 B.n36 10.6151
R691 B.n446 B.n445 10.6151
R692 B.n445 B.n444 10.6151
R693 B.n444 B.n38 10.6151
R694 B.n440 B.n38 10.6151
R695 B.n440 B.n439 10.6151
R696 B.n437 B.n42 10.6151
R697 B.n433 B.n42 10.6151
R698 B.n433 B.n432 10.6151
R699 B.n432 B.n431 10.6151
R700 B.n431 B.n44 10.6151
R701 B.n427 B.n44 10.6151
R702 B.n427 B.n426 10.6151
R703 B.n426 B.n425 10.6151
R704 B.n425 B.n46 10.6151
R705 B.n421 B.n46 10.6151
R706 B.n269 B.n98 10.6151
R707 B.n270 B.n269 10.6151
R708 B.n271 B.n270 10.6151
R709 B.n271 B.n96 10.6151
R710 B.n275 B.n96 10.6151
R711 B.n276 B.n275 10.6151
R712 B.n277 B.n276 10.6151
R713 B.n277 B.n94 10.6151
R714 B.n281 B.n94 10.6151
R715 B.n282 B.n281 10.6151
R716 B.n283 B.n282 10.6151
R717 B.n283 B.n92 10.6151
R718 B.n287 B.n92 10.6151
R719 B.n288 B.n287 10.6151
R720 B.n289 B.n288 10.6151
R721 B.n289 B.n90 10.6151
R722 B.n293 B.n90 10.6151
R723 B.n294 B.n293 10.6151
R724 B.n295 B.n294 10.6151
R725 B.n295 B.n88 10.6151
R726 B.n299 B.n88 10.6151
R727 B.n300 B.n299 10.6151
R728 B.n301 B.n300 10.6151
R729 B.n301 B.n86 10.6151
R730 B.n305 B.n86 10.6151
R731 B.n306 B.n305 10.6151
R732 B.n307 B.n306 10.6151
R733 B.n307 B.n84 10.6151
R734 B.n311 B.n84 10.6151
R735 B.n312 B.n311 10.6151
R736 B.n313 B.n312 10.6151
R737 B.n313 B.n82 10.6151
R738 B.n317 B.n82 10.6151
R739 B.n318 B.n317 10.6151
R740 B.n319 B.n318 10.6151
R741 B.n319 B.n80 10.6151
R742 B.n323 B.n80 10.6151
R743 B.n324 B.n323 10.6151
R744 B.n325 B.n324 10.6151
R745 B.n325 B.n78 10.6151
R746 B.n329 B.n78 10.6151
R747 B.n330 B.n329 10.6151
R748 B.n331 B.n330 10.6151
R749 B.n331 B.n76 10.6151
R750 B.n335 B.n76 10.6151
R751 B.n336 B.n335 10.6151
R752 B.n337 B.n336 10.6151
R753 B.n337 B.n74 10.6151
R754 B.n341 B.n74 10.6151
R755 B.n342 B.n341 10.6151
R756 B.n343 B.n342 10.6151
R757 B.n343 B.n72 10.6151
R758 B.n347 B.n72 10.6151
R759 B.n348 B.n347 10.6151
R760 B.n349 B.n348 10.6151
R761 B.n349 B.n70 10.6151
R762 B.n353 B.n70 10.6151
R763 B.n354 B.n353 10.6151
R764 B.n355 B.n354 10.6151
R765 B.n355 B.n68 10.6151
R766 B.n359 B.n68 10.6151
R767 B.n360 B.n359 10.6151
R768 B.n361 B.n360 10.6151
R769 B.n361 B.n66 10.6151
R770 B.n365 B.n66 10.6151
R771 B.n366 B.n365 10.6151
R772 B.n367 B.n366 10.6151
R773 B.n367 B.n64 10.6151
R774 B.n371 B.n64 10.6151
R775 B.n372 B.n371 10.6151
R776 B.n373 B.n372 10.6151
R777 B.n373 B.n62 10.6151
R778 B.n377 B.n62 10.6151
R779 B.n378 B.n377 10.6151
R780 B.n379 B.n378 10.6151
R781 B.n379 B.n60 10.6151
R782 B.n383 B.n60 10.6151
R783 B.n384 B.n383 10.6151
R784 B.n385 B.n384 10.6151
R785 B.n385 B.n58 10.6151
R786 B.n389 B.n58 10.6151
R787 B.n390 B.n389 10.6151
R788 B.n391 B.n390 10.6151
R789 B.n391 B.n56 10.6151
R790 B.n395 B.n56 10.6151
R791 B.n396 B.n395 10.6151
R792 B.n397 B.n396 10.6151
R793 B.n397 B.n54 10.6151
R794 B.n401 B.n54 10.6151
R795 B.n402 B.n401 10.6151
R796 B.n403 B.n402 10.6151
R797 B.n403 B.n52 10.6151
R798 B.n407 B.n52 10.6151
R799 B.n408 B.n407 10.6151
R800 B.n409 B.n408 10.6151
R801 B.n409 B.n50 10.6151
R802 B.n413 B.n50 10.6151
R803 B.n414 B.n413 10.6151
R804 B.n415 B.n414 10.6151
R805 B.n415 B.n48 10.6151
R806 B.n419 B.n48 10.6151
R807 B.n420 B.n419 10.6151
R808 B.n221 B.n118 10.6151
R809 B.n222 B.n221 10.6151
R810 B.n223 B.n222 10.6151
R811 B.n223 B.n116 10.6151
R812 B.n227 B.n116 10.6151
R813 B.n228 B.n227 10.6151
R814 B.n229 B.n228 10.6151
R815 B.n229 B.n114 10.6151
R816 B.n233 B.n114 10.6151
R817 B.n234 B.n233 10.6151
R818 B.n236 B.n110 10.6151
R819 B.n240 B.n110 10.6151
R820 B.n241 B.n240 10.6151
R821 B.n242 B.n241 10.6151
R822 B.n242 B.n108 10.6151
R823 B.n246 B.n108 10.6151
R824 B.n247 B.n246 10.6151
R825 B.n248 B.n247 10.6151
R826 B.n252 B.n251 10.6151
R827 B.n253 B.n252 10.6151
R828 B.n253 B.n102 10.6151
R829 B.n257 B.n102 10.6151
R830 B.n258 B.n257 10.6151
R831 B.n259 B.n258 10.6151
R832 B.n259 B.n100 10.6151
R833 B.n263 B.n100 10.6151
R834 B.n264 B.n263 10.6151
R835 B.n265 B.n264 10.6151
R836 B.n217 B.n216 10.6151
R837 B.n216 B.n215 10.6151
R838 B.n215 B.n120 10.6151
R839 B.n211 B.n120 10.6151
R840 B.n211 B.n210 10.6151
R841 B.n210 B.n209 10.6151
R842 B.n209 B.n122 10.6151
R843 B.n205 B.n122 10.6151
R844 B.n205 B.n204 10.6151
R845 B.n204 B.n203 10.6151
R846 B.n203 B.n124 10.6151
R847 B.n199 B.n124 10.6151
R848 B.n199 B.n198 10.6151
R849 B.n198 B.n197 10.6151
R850 B.n197 B.n126 10.6151
R851 B.n193 B.n126 10.6151
R852 B.n193 B.n192 10.6151
R853 B.n192 B.n191 10.6151
R854 B.n191 B.n128 10.6151
R855 B.n187 B.n128 10.6151
R856 B.n187 B.n186 10.6151
R857 B.n186 B.n185 10.6151
R858 B.n185 B.n130 10.6151
R859 B.n181 B.n130 10.6151
R860 B.n181 B.n180 10.6151
R861 B.n180 B.n179 10.6151
R862 B.n179 B.n132 10.6151
R863 B.n175 B.n132 10.6151
R864 B.n175 B.n174 10.6151
R865 B.n174 B.n173 10.6151
R866 B.n173 B.n134 10.6151
R867 B.n169 B.n134 10.6151
R868 B.n169 B.n168 10.6151
R869 B.n168 B.n167 10.6151
R870 B.n167 B.n136 10.6151
R871 B.n163 B.n136 10.6151
R872 B.n163 B.n162 10.6151
R873 B.n162 B.n161 10.6151
R874 B.n161 B.n138 10.6151
R875 B.n157 B.n138 10.6151
R876 B.n157 B.n156 10.6151
R877 B.n156 B.n155 10.6151
R878 B.n155 B.n140 10.6151
R879 B.n151 B.n140 10.6151
R880 B.n151 B.n150 10.6151
R881 B.n150 B.n149 10.6151
R882 B.n149 B.n142 10.6151
R883 B.n145 B.n142 10.6151
R884 B.n145 B.n144 10.6151
R885 B.n144 B.n0 10.6151
R886 B.n543 B.n1 10.6151
R887 B.n543 B.n542 10.6151
R888 B.n542 B.n541 10.6151
R889 B.n541 B.n4 10.6151
R890 B.n537 B.n4 10.6151
R891 B.n537 B.n536 10.6151
R892 B.n536 B.n535 10.6151
R893 B.n535 B.n6 10.6151
R894 B.n531 B.n6 10.6151
R895 B.n531 B.n530 10.6151
R896 B.n530 B.n529 10.6151
R897 B.n529 B.n8 10.6151
R898 B.n525 B.n8 10.6151
R899 B.n525 B.n524 10.6151
R900 B.n524 B.n523 10.6151
R901 B.n523 B.n10 10.6151
R902 B.n519 B.n10 10.6151
R903 B.n519 B.n518 10.6151
R904 B.n518 B.n517 10.6151
R905 B.n517 B.n12 10.6151
R906 B.n513 B.n12 10.6151
R907 B.n513 B.n512 10.6151
R908 B.n512 B.n511 10.6151
R909 B.n511 B.n14 10.6151
R910 B.n507 B.n14 10.6151
R911 B.n507 B.n506 10.6151
R912 B.n506 B.n505 10.6151
R913 B.n505 B.n16 10.6151
R914 B.n501 B.n16 10.6151
R915 B.n501 B.n500 10.6151
R916 B.n500 B.n499 10.6151
R917 B.n499 B.n18 10.6151
R918 B.n495 B.n18 10.6151
R919 B.n495 B.n494 10.6151
R920 B.n494 B.n493 10.6151
R921 B.n493 B.n20 10.6151
R922 B.n489 B.n20 10.6151
R923 B.n489 B.n488 10.6151
R924 B.n488 B.n487 10.6151
R925 B.n487 B.n22 10.6151
R926 B.n483 B.n22 10.6151
R927 B.n483 B.n482 10.6151
R928 B.n482 B.n481 10.6151
R929 B.n481 B.n24 10.6151
R930 B.n477 B.n24 10.6151
R931 B.n477 B.n476 10.6151
R932 B.n476 B.n475 10.6151
R933 B.n475 B.n26 10.6151
R934 B.n471 B.n26 10.6151
R935 B.n471 B.n470 10.6151
R936 B.n452 B.n451 6.5566
R937 B.n439 B.n438 6.5566
R938 B.n236 B.n235 6.5566
R939 B.n248 B.n106 6.5566
R940 B.n453 B.n452 4.05904
R941 B.n438 B.n437 4.05904
R942 B.n235 B.n234 4.05904
R943 B.n251 B.n106 4.05904
R944 B.n547 B.n0 2.81026
R945 B.n547 B.n1 2.81026
R946 VN.n34 VN.n33 161.3
R947 VN.n32 VN.n19 161.3
R948 VN.n31 VN.n30 161.3
R949 VN.n29 VN.n20 161.3
R950 VN.n28 VN.n27 161.3
R951 VN.n26 VN.n21 161.3
R952 VN.n25 VN.n24 161.3
R953 VN.n16 VN.n15 161.3
R954 VN.n14 VN.n1 161.3
R955 VN.n13 VN.n12 161.3
R956 VN.n11 VN.n2 161.3
R957 VN.n10 VN.n9 161.3
R958 VN.n8 VN.n3 161.3
R959 VN.n7 VN.n6 161.3
R960 VN.n17 VN.n0 82.1011
R961 VN.n35 VN.n18 82.1011
R962 VN.n9 VN.n2 56.4773
R963 VN.n27 VN.n20 56.4773
R964 VN.n5 VN.n4 49.9597
R965 VN.n23 VN.n22 49.9597
R966 VN.n23 VN.t2 44.2307
R967 VN.n5 VN.t1 44.2307
R968 VN VN.n35 43.8085
R969 VN.n7 VN.n4 24.3439
R970 VN.n8 VN.n7 24.3439
R971 VN.n9 VN.n8 24.3439
R972 VN.n13 VN.n2 24.3439
R973 VN.n14 VN.n13 24.3439
R974 VN.n15 VN.n14 24.3439
R975 VN.n27 VN.n26 24.3439
R976 VN.n26 VN.n25 24.3439
R977 VN.n25 VN.n22 24.3439
R978 VN.n33 VN.n32 24.3439
R979 VN.n32 VN.n31 24.3439
R980 VN.n31 VN.n20 24.3439
R981 VN.n4 VN.t0 11.2906
R982 VN.n0 VN.t3 11.2906
R983 VN.n22 VN.t5 11.2906
R984 VN.n18 VN.t4 11.2906
R985 VN.n15 VN.n0 7.7904
R986 VN.n33 VN.n18 7.7904
R987 VN.n24 VN.n23 3.24066
R988 VN.n6 VN.n5 3.24066
R989 VN.n35 VN.n34 0.355081
R990 VN.n17 VN.n16 0.355081
R991 VN VN.n17 0.26685
R992 VN.n34 VN.n19 0.189894
R993 VN.n30 VN.n19 0.189894
R994 VN.n30 VN.n29 0.189894
R995 VN.n29 VN.n28 0.189894
R996 VN.n28 VN.n21 0.189894
R997 VN.n24 VN.n21 0.189894
R998 VN.n6 VN.n3 0.189894
R999 VN.n10 VN.n3 0.189894
R1000 VN.n11 VN.n10 0.189894
R1001 VN.n12 VN.n11 0.189894
R1002 VN.n12 VN.n1 0.189894
R1003 VN.n16 VN.n1 0.189894
R1004 VDD2.n1 VDD2.t4 270.932
R1005 VDD2.n2 VDD2.t1 268.62
R1006 VDD2.n1 VDD2.n0 248.518
R1007 VDD2 VDD2.n3 248.514
R1008 VDD2.n2 VDD2.n1 35.3144
R1009 VDD2.n3 VDD2.t0 20.837
R1010 VDD2.n3 VDD2.t3 20.837
R1011 VDD2.n0 VDD2.t5 20.837
R1012 VDD2.n0 VDD2.t2 20.837
R1013 VDD2 VDD2.n2 2.42507
C0 VDD1 B 1.44526f
C1 VP VTAIL 2.43622f
C2 VDD2 VP 0.527789f
C3 VP VN 5.72192f
C4 VP w_n3898_n1280# 7.90092f
C5 VDD2 VTAIL 4.53894f
C6 VN VTAIL 2.42209f
C7 w_n3898_n1280# VTAIL 1.55974f
C8 VDD1 VP 1.62682f
C9 VP B 2.0167f
C10 VDD2 VN 1.26093f
C11 VDD2 w_n3898_n1280# 1.85341f
C12 w_n3898_n1280# VN 7.40091f
C13 VDD1 VTAIL 4.48068f
C14 VTAIL B 1.38153f
C15 VDD2 VDD1 1.69145f
C16 VDD2 B 1.5374f
C17 VDD1 VN 0.158549f
C18 VN B 1.16916f
C19 VDD1 w_n3898_n1280# 1.74586f
C20 w_n3898_n1280# B 7.82988f
C21 VDD2 VSUBS 1.189525f
C22 VDD1 VSUBS 1.711094f
C23 VTAIL VSUBS 0.610042f
C24 VN VSUBS 6.66604f
C25 VP VSUBS 2.890996f
C26 B VSUBS 4.201984f
C27 w_n3898_n1280# VSUBS 63.942802f
C28 VDD2.t4 VSUBS 0.134702f
C29 VDD2.t5 VSUBS 0.021893f
C30 VDD2.t2 VSUBS 0.021893f
C31 VDD2.n0 VSUBS 0.082699f
C32 VDD2.n1 VSUBS 1.86885f
C33 VDD2.t1 VSUBS 0.131965f
C34 VDD2.n2 VSUBS 1.53062f
C35 VDD2.t0 VSUBS 0.021893f
C36 VDD2.t3 VSUBS 0.021893f
C37 VDD2.n3 VSUBS 0.082692f
C38 VN.t3 VSUBS 0.585071f
C39 VN.n0 VSUBS 0.478711f
C40 VN.n1 VSUBS 0.051109f
C41 VN.n2 VSUBS 0.06346f
C42 VN.n3 VSUBS 0.051109f
C43 VN.t0 VSUBS 0.585071f
C44 VN.n4 VSUBS 0.496744f
C45 VN.t1 VSUBS 1.08198f
C46 VN.n5 VSUBS 0.522857f
C47 VN.n6 VSUBS 0.623199f
C48 VN.n7 VSUBS 0.095732f
C49 VN.n8 VSUBS 0.095732f
C50 VN.n9 VSUBS 0.086409f
C51 VN.n10 VSUBS 0.051109f
C52 VN.n11 VSUBS 0.051109f
C53 VN.n12 VSUBS 0.051109f
C54 VN.n13 VSUBS 0.095732f
C55 VN.n14 VSUBS 0.095732f
C56 VN.n15 VSUBS 0.063591f
C57 VN.n16 VSUBS 0.082502f
C58 VN.n17 VSUBS 0.136851f
C59 VN.t4 VSUBS 0.585071f
C60 VN.n18 VSUBS 0.478711f
C61 VN.n19 VSUBS 0.051109f
C62 VN.n20 VSUBS 0.06346f
C63 VN.n21 VSUBS 0.051109f
C64 VN.t5 VSUBS 0.585071f
C65 VN.n22 VSUBS 0.496744f
C66 VN.t2 VSUBS 1.08198f
C67 VN.n23 VSUBS 0.522857f
C68 VN.n24 VSUBS 0.623199f
C69 VN.n25 VSUBS 0.095732f
C70 VN.n26 VSUBS 0.095732f
C71 VN.n27 VSUBS 0.086409f
C72 VN.n28 VSUBS 0.051109f
C73 VN.n29 VSUBS 0.051109f
C74 VN.n30 VSUBS 0.051109f
C75 VN.n31 VSUBS 0.095732f
C76 VN.n32 VSUBS 0.095732f
C77 VN.n33 VSUBS 0.063591f
C78 VN.n34 VSUBS 0.082502f
C79 VN.n35 VSUBS 2.40701f
C80 B.n0 VSUBS 0.007429f
C81 B.n1 VSUBS 0.007429f
C82 B.n2 VSUBS 0.011748f
C83 B.n3 VSUBS 0.011748f
C84 B.n4 VSUBS 0.011748f
C85 B.n5 VSUBS 0.011748f
C86 B.n6 VSUBS 0.011748f
C87 B.n7 VSUBS 0.011748f
C88 B.n8 VSUBS 0.011748f
C89 B.n9 VSUBS 0.011748f
C90 B.n10 VSUBS 0.011748f
C91 B.n11 VSUBS 0.011748f
C92 B.n12 VSUBS 0.011748f
C93 B.n13 VSUBS 0.011748f
C94 B.n14 VSUBS 0.011748f
C95 B.n15 VSUBS 0.011748f
C96 B.n16 VSUBS 0.011748f
C97 B.n17 VSUBS 0.011748f
C98 B.n18 VSUBS 0.011748f
C99 B.n19 VSUBS 0.011748f
C100 B.n20 VSUBS 0.011748f
C101 B.n21 VSUBS 0.011748f
C102 B.n22 VSUBS 0.011748f
C103 B.n23 VSUBS 0.011748f
C104 B.n24 VSUBS 0.011748f
C105 B.n25 VSUBS 0.011748f
C106 B.n26 VSUBS 0.011748f
C107 B.n27 VSUBS 0.028981f
C108 B.n28 VSUBS 0.011748f
C109 B.n29 VSUBS 0.011748f
C110 B.n30 VSUBS 0.011748f
C111 B.n31 VSUBS 0.011748f
C112 B.n32 VSUBS 0.011748f
C113 B.n33 VSUBS 0.011748f
C114 B.t2 VSUBS 0.05347f
C115 B.t1 VSUBS 0.070771f
C116 B.t0 VSUBS 0.438771f
C117 B.n34 VSUBS 0.119986f
C118 B.n35 VSUBS 0.094936f
C119 B.n36 VSUBS 0.011748f
C120 B.n37 VSUBS 0.011748f
C121 B.n38 VSUBS 0.011748f
C122 B.n39 VSUBS 0.011748f
C123 B.t11 VSUBS 0.05347f
C124 B.t10 VSUBS 0.070771f
C125 B.t9 VSUBS 0.438771f
C126 B.n40 VSUBS 0.119986f
C127 B.n41 VSUBS 0.094936f
C128 B.n42 VSUBS 0.011748f
C129 B.n43 VSUBS 0.011748f
C130 B.n44 VSUBS 0.011748f
C131 B.n45 VSUBS 0.011748f
C132 B.n46 VSUBS 0.011748f
C133 B.n47 VSUBS 0.028981f
C134 B.n48 VSUBS 0.011748f
C135 B.n49 VSUBS 0.011748f
C136 B.n50 VSUBS 0.011748f
C137 B.n51 VSUBS 0.011748f
C138 B.n52 VSUBS 0.011748f
C139 B.n53 VSUBS 0.011748f
C140 B.n54 VSUBS 0.011748f
C141 B.n55 VSUBS 0.011748f
C142 B.n56 VSUBS 0.011748f
C143 B.n57 VSUBS 0.011748f
C144 B.n58 VSUBS 0.011748f
C145 B.n59 VSUBS 0.011748f
C146 B.n60 VSUBS 0.011748f
C147 B.n61 VSUBS 0.011748f
C148 B.n62 VSUBS 0.011748f
C149 B.n63 VSUBS 0.011748f
C150 B.n64 VSUBS 0.011748f
C151 B.n65 VSUBS 0.011748f
C152 B.n66 VSUBS 0.011748f
C153 B.n67 VSUBS 0.011748f
C154 B.n68 VSUBS 0.011748f
C155 B.n69 VSUBS 0.011748f
C156 B.n70 VSUBS 0.011748f
C157 B.n71 VSUBS 0.011748f
C158 B.n72 VSUBS 0.011748f
C159 B.n73 VSUBS 0.011748f
C160 B.n74 VSUBS 0.011748f
C161 B.n75 VSUBS 0.011748f
C162 B.n76 VSUBS 0.011748f
C163 B.n77 VSUBS 0.011748f
C164 B.n78 VSUBS 0.011748f
C165 B.n79 VSUBS 0.011748f
C166 B.n80 VSUBS 0.011748f
C167 B.n81 VSUBS 0.011748f
C168 B.n82 VSUBS 0.011748f
C169 B.n83 VSUBS 0.011748f
C170 B.n84 VSUBS 0.011748f
C171 B.n85 VSUBS 0.011748f
C172 B.n86 VSUBS 0.011748f
C173 B.n87 VSUBS 0.011748f
C174 B.n88 VSUBS 0.011748f
C175 B.n89 VSUBS 0.011748f
C176 B.n90 VSUBS 0.011748f
C177 B.n91 VSUBS 0.011748f
C178 B.n92 VSUBS 0.011748f
C179 B.n93 VSUBS 0.011748f
C180 B.n94 VSUBS 0.011748f
C181 B.n95 VSUBS 0.011748f
C182 B.n96 VSUBS 0.011748f
C183 B.n97 VSUBS 0.011748f
C184 B.n98 VSUBS 0.028981f
C185 B.n99 VSUBS 0.011748f
C186 B.n100 VSUBS 0.011748f
C187 B.n101 VSUBS 0.011748f
C188 B.n102 VSUBS 0.011748f
C189 B.n103 VSUBS 0.011748f
C190 B.t7 VSUBS 0.05347f
C191 B.t8 VSUBS 0.070771f
C192 B.t6 VSUBS 0.438771f
C193 B.n104 VSUBS 0.119986f
C194 B.n105 VSUBS 0.094936f
C195 B.n106 VSUBS 0.02722f
C196 B.n107 VSUBS 0.011748f
C197 B.n108 VSUBS 0.011748f
C198 B.n109 VSUBS 0.011748f
C199 B.n110 VSUBS 0.011748f
C200 B.n111 VSUBS 0.011748f
C201 B.t4 VSUBS 0.05347f
C202 B.t5 VSUBS 0.070771f
C203 B.t3 VSUBS 0.438771f
C204 B.n112 VSUBS 0.119986f
C205 B.n113 VSUBS 0.094936f
C206 B.n114 VSUBS 0.011748f
C207 B.n115 VSUBS 0.011748f
C208 B.n116 VSUBS 0.011748f
C209 B.n117 VSUBS 0.011748f
C210 B.n118 VSUBS 0.030106f
C211 B.n119 VSUBS 0.011748f
C212 B.n120 VSUBS 0.011748f
C213 B.n121 VSUBS 0.011748f
C214 B.n122 VSUBS 0.011748f
C215 B.n123 VSUBS 0.011748f
C216 B.n124 VSUBS 0.011748f
C217 B.n125 VSUBS 0.011748f
C218 B.n126 VSUBS 0.011748f
C219 B.n127 VSUBS 0.011748f
C220 B.n128 VSUBS 0.011748f
C221 B.n129 VSUBS 0.011748f
C222 B.n130 VSUBS 0.011748f
C223 B.n131 VSUBS 0.011748f
C224 B.n132 VSUBS 0.011748f
C225 B.n133 VSUBS 0.011748f
C226 B.n134 VSUBS 0.011748f
C227 B.n135 VSUBS 0.011748f
C228 B.n136 VSUBS 0.011748f
C229 B.n137 VSUBS 0.011748f
C230 B.n138 VSUBS 0.011748f
C231 B.n139 VSUBS 0.011748f
C232 B.n140 VSUBS 0.011748f
C233 B.n141 VSUBS 0.011748f
C234 B.n142 VSUBS 0.011748f
C235 B.n143 VSUBS 0.011748f
C236 B.n144 VSUBS 0.011748f
C237 B.n145 VSUBS 0.011748f
C238 B.n146 VSUBS 0.011748f
C239 B.n147 VSUBS 0.011748f
C240 B.n148 VSUBS 0.011748f
C241 B.n149 VSUBS 0.011748f
C242 B.n150 VSUBS 0.011748f
C243 B.n151 VSUBS 0.011748f
C244 B.n152 VSUBS 0.011748f
C245 B.n153 VSUBS 0.011748f
C246 B.n154 VSUBS 0.011748f
C247 B.n155 VSUBS 0.011748f
C248 B.n156 VSUBS 0.011748f
C249 B.n157 VSUBS 0.011748f
C250 B.n158 VSUBS 0.011748f
C251 B.n159 VSUBS 0.011748f
C252 B.n160 VSUBS 0.011748f
C253 B.n161 VSUBS 0.011748f
C254 B.n162 VSUBS 0.011748f
C255 B.n163 VSUBS 0.011748f
C256 B.n164 VSUBS 0.011748f
C257 B.n165 VSUBS 0.011748f
C258 B.n166 VSUBS 0.011748f
C259 B.n167 VSUBS 0.011748f
C260 B.n168 VSUBS 0.011748f
C261 B.n169 VSUBS 0.011748f
C262 B.n170 VSUBS 0.011748f
C263 B.n171 VSUBS 0.011748f
C264 B.n172 VSUBS 0.011748f
C265 B.n173 VSUBS 0.011748f
C266 B.n174 VSUBS 0.011748f
C267 B.n175 VSUBS 0.011748f
C268 B.n176 VSUBS 0.011748f
C269 B.n177 VSUBS 0.011748f
C270 B.n178 VSUBS 0.011748f
C271 B.n179 VSUBS 0.011748f
C272 B.n180 VSUBS 0.011748f
C273 B.n181 VSUBS 0.011748f
C274 B.n182 VSUBS 0.011748f
C275 B.n183 VSUBS 0.011748f
C276 B.n184 VSUBS 0.011748f
C277 B.n185 VSUBS 0.011748f
C278 B.n186 VSUBS 0.011748f
C279 B.n187 VSUBS 0.011748f
C280 B.n188 VSUBS 0.011748f
C281 B.n189 VSUBS 0.011748f
C282 B.n190 VSUBS 0.011748f
C283 B.n191 VSUBS 0.011748f
C284 B.n192 VSUBS 0.011748f
C285 B.n193 VSUBS 0.011748f
C286 B.n194 VSUBS 0.011748f
C287 B.n195 VSUBS 0.011748f
C288 B.n196 VSUBS 0.011748f
C289 B.n197 VSUBS 0.011748f
C290 B.n198 VSUBS 0.011748f
C291 B.n199 VSUBS 0.011748f
C292 B.n200 VSUBS 0.011748f
C293 B.n201 VSUBS 0.011748f
C294 B.n202 VSUBS 0.011748f
C295 B.n203 VSUBS 0.011748f
C296 B.n204 VSUBS 0.011748f
C297 B.n205 VSUBS 0.011748f
C298 B.n206 VSUBS 0.011748f
C299 B.n207 VSUBS 0.011748f
C300 B.n208 VSUBS 0.011748f
C301 B.n209 VSUBS 0.011748f
C302 B.n210 VSUBS 0.011748f
C303 B.n211 VSUBS 0.011748f
C304 B.n212 VSUBS 0.011748f
C305 B.n213 VSUBS 0.011748f
C306 B.n214 VSUBS 0.011748f
C307 B.n215 VSUBS 0.011748f
C308 B.n216 VSUBS 0.011748f
C309 B.n217 VSUBS 0.028981f
C310 B.n218 VSUBS 0.028981f
C311 B.n219 VSUBS 0.030106f
C312 B.n220 VSUBS 0.011748f
C313 B.n221 VSUBS 0.011748f
C314 B.n222 VSUBS 0.011748f
C315 B.n223 VSUBS 0.011748f
C316 B.n224 VSUBS 0.011748f
C317 B.n225 VSUBS 0.011748f
C318 B.n226 VSUBS 0.011748f
C319 B.n227 VSUBS 0.011748f
C320 B.n228 VSUBS 0.011748f
C321 B.n229 VSUBS 0.011748f
C322 B.n230 VSUBS 0.011748f
C323 B.n231 VSUBS 0.011748f
C324 B.n232 VSUBS 0.011748f
C325 B.n233 VSUBS 0.011748f
C326 B.n234 VSUBS 0.00812f
C327 B.n235 VSUBS 0.02722f
C328 B.n236 VSUBS 0.009502f
C329 B.n237 VSUBS 0.011748f
C330 B.n238 VSUBS 0.011748f
C331 B.n239 VSUBS 0.011748f
C332 B.n240 VSUBS 0.011748f
C333 B.n241 VSUBS 0.011748f
C334 B.n242 VSUBS 0.011748f
C335 B.n243 VSUBS 0.011748f
C336 B.n244 VSUBS 0.011748f
C337 B.n245 VSUBS 0.011748f
C338 B.n246 VSUBS 0.011748f
C339 B.n247 VSUBS 0.011748f
C340 B.n248 VSUBS 0.009502f
C341 B.n249 VSUBS 0.011748f
C342 B.n250 VSUBS 0.011748f
C343 B.n251 VSUBS 0.00812f
C344 B.n252 VSUBS 0.011748f
C345 B.n253 VSUBS 0.011748f
C346 B.n254 VSUBS 0.011748f
C347 B.n255 VSUBS 0.011748f
C348 B.n256 VSUBS 0.011748f
C349 B.n257 VSUBS 0.011748f
C350 B.n258 VSUBS 0.011748f
C351 B.n259 VSUBS 0.011748f
C352 B.n260 VSUBS 0.011748f
C353 B.n261 VSUBS 0.011748f
C354 B.n262 VSUBS 0.011748f
C355 B.n263 VSUBS 0.011748f
C356 B.n264 VSUBS 0.011748f
C357 B.n265 VSUBS 0.030106f
C358 B.n266 VSUBS 0.030106f
C359 B.n267 VSUBS 0.028981f
C360 B.n268 VSUBS 0.011748f
C361 B.n269 VSUBS 0.011748f
C362 B.n270 VSUBS 0.011748f
C363 B.n271 VSUBS 0.011748f
C364 B.n272 VSUBS 0.011748f
C365 B.n273 VSUBS 0.011748f
C366 B.n274 VSUBS 0.011748f
C367 B.n275 VSUBS 0.011748f
C368 B.n276 VSUBS 0.011748f
C369 B.n277 VSUBS 0.011748f
C370 B.n278 VSUBS 0.011748f
C371 B.n279 VSUBS 0.011748f
C372 B.n280 VSUBS 0.011748f
C373 B.n281 VSUBS 0.011748f
C374 B.n282 VSUBS 0.011748f
C375 B.n283 VSUBS 0.011748f
C376 B.n284 VSUBS 0.011748f
C377 B.n285 VSUBS 0.011748f
C378 B.n286 VSUBS 0.011748f
C379 B.n287 VSUBS 0.011748f
C380 B.n288 VSUBS 0.011748f
C381 B.n289 VSUBS 0.011748f
C382 B.n290 VSUBS 0.011748f
C383 B.n291 VSUBS 0.011748f
C384 B.n292 VSUBS 0.011748f
C385 B.n293 VSUBS 0.011748f
C386 B.n294 VSUBS 0.011748f
C387 B.n295 VSUBS 0.011748f
C388 B.n296 VSUBS 0.011748f
C389 B.n297 VSUBS 0.011748f
C390 B.n298 VSUBS 0.011748f
C391 B.n299 VSUBS 0.011748f
C392 B.n300 VSUBS 0.011748f
C393 B.n301 VSUBS 0.011748f
C394 B.n302 VSUBS 0.011748f
C395 B.n303 VSUBS 0.011748f
C396 B.n304 VSUBS 0.011748f
C397 B.n305 VSUBS 0.011748f
C398 B.n306 VSUBS 0.011748f
C399 B.n307 VSUBS 0.011748f
C400 B.n308 VSUBS 0.011748f
C401 B.n309 VSUBS 0.011748f
C402 B.n310 VSUBS 0.011748f
C403 B.n311 VSUBS 0.011748f
C404 B.n312 VSUBS 0.011748f
C405 B.n313 VSUBS 0.011748f
C406 B.n314 VSUBS 0.011748f
C407 B.n315 VSUBS 0.011748f
C408 B.n316 VSUBS 0.011748f
C409 B.n317 VSUBS 0.011748f
C410 B.n318 VSUBS 0.011748f
C411 B.n319 VSUBS 0.011748f
C412 B.n320 VSUBS 0.011748f
C413 B.n321 VSUBS 0.011748f
C414 B.n322 VSUBS 0.011748f
C415 B.n323 VSUBS 0.011748f
C416 B.n324 VSUBS 0.011748f
C417 B.n325 VSUBS 0.011748f
C418 B.n326 VSUBS 0.011748f
C419 B.n327 VSUBS 0.011748f
C420 B.n328 VSUBS 0.011748f
C421 B.n329 VSUBS 0.011748f
C422 B.n330 VSUBS 0.011748f
C423 B.n331 VSUBS 0.011748f
C424 B.n332 VSUBS 0.011748f
C425 B.n333 VSUBS 0.011748f
C426 B.n334 VSUBS 0.011748f
C427 B.n335 VSUBS 0.011748f
C428 B.n336 VSUBS 0.011748f
C429 B.n337 VSUBS 0.011748f
C430 B.n338 VSUBS 0.011748f
C431 B.n339 VSUBS 0.011748f
C432 B.n340 VSUBS 0.011748f
C433 B.n341 VSUBS 0.011748f
C434 B.n342 VSUBS 0.011748f
C435 B.n343 VSUBS 0.011748f
C436 B.n344 VSUBS 0.011748f
C437 B.n345 VSUBS 0.011748f
C438 B.n346 VSUBS 0.011748f
C439 B.n347 VSUBS 0.011748f
C440 B.n348 VSUBS 0.011748f
C441 B.n349 VSUBS 0.011748f
C442 B.n350 VSUBS 0.011748f
C443 B.n351 VSUBS 0.011748f
C444 B.n352 VSUBS 0.011748f
C445 B.n353 VSUBS 0.011748f
C446 B.n354 VSUBS 0.011748f
C447 B.n355 VSUBS 0.011748f
C448 B.n356 VSUBS 0.011748f
C449 B.n357 VSUBS 0.011748f
C450 B.n358 VSUBS 0.011748f
C451 B.n359 VSUBS 0.011748f
C452 B.n360 VSUBS 0.011748f
C453 B.n361 VSUBS 0.011748f
C454 B.n362 VSUBS 0.011748f
C455 B.n363 VSUBS 0.011748f
C456 B.n364 VSUBS 0.011748f
C457 B.n365 VSUBS 0.011748f
C458 B.n366 VSUBS 0.011748f
C459 B.n367 VSUBS 0.011748f
C460 B.n368 VSUBS 0.011748f
C461 B.n369 VSUBS 0.011748f
C462 B.n370 VSUBS 0.011748f
C463 B.n371 VSUBS 0.011748f
C464 B.n372 VSUBS 0.011748f
C465 B.n373 VSUBS 0.011748f
C466 B.n374 VSUBS 0.011748f
C467 B.n375 VSUBS 0.011748f
C468 B.n376 VSUBS 0.011748f
C469 B.n377 VSUBS 0.011748f
C470 B.n378 VSUBS 0.011748f
C471 B.n379 VSUBS 0.011748f
C472 B.n380 VSUBS 0.011748f
C473 B.n381 VSUBS 0.011748f
C474 B.n382 VSUBS 0.011748f
C475 B.n383 VSUBS 0.011748f
C476 B.n384 VSUBS 0.011748f
C477 B.n385 VSUBS 0.011748f
C478 B.n386 VSUBS 0.011748f
C479 B.n387 VSUBS 0.011748f
C480 B.n388 VSUBS 0.011748f
C481 B.n389 VSUBS 0.011748f
C482 B.n390 VSUBS 0.011748f
C483 B.n391 VSUBS 0.011748f
C484 B.n392 VSUBS 0.011748f
C485 B.n393 VSUBS 0.011748f
C486 B.n394 VSUBS 0.011748f
C487 B.n395 VSUBS 0.011748f
C488 B.n396 VSUBS 0.011748f
C489 B.n397 VSUBS 0.011748f
C490 B.n398 VSUBS 0.011748f
C491 B.n399 VSUBS 0.011748f
C492 B.n400 VSUBS 0.011748f
C493 B.n401 VSUBS 0.011748f
C494 B.n402 VSUBS 0.011748f
C495 B.n403 VSUBS 0.011748f
C496 B.n404 VSUBS 0.011748f
C497 B.n405 VSUBS 0.011748f
C498 B.n406 VSUBS 0.011748f
C499 B.n407 VSUBS 0.011748f
C500 B.n408 VSUBS 0.011748f
C501 B.n409 VSUBS 0.011748f
C502 B.n410 VSUBS 0.011748f
C503 B.n411 VSUBS 0.011748f
C504 B.n412 VSUBS 0.011748f
C505 B.n413 VSUBS 0.011748f
C506 B.n414 VSUBS 0.011748f
C507 B.n415 VSUBS 0.011748f
C508 B.n416 VSUBS 0.011748f
C509 B.n417 VSUBS 0.011748f
C510 B.n418 VSUBS 0.011748f
C511 B.n419 VSUBS 0.011748f
C512 B.n420 VSUBS 0.030228f
C513 B.n421 VSUBS 0.02886f
C514 B.n422 VSUBS 0.030106f
C515 B.n423 VSUBS 0.011748f
C516 B.n424 VSUBS 0.011748f
C517 B.n425 VSUBS 0.011748f
C518 B.n426 VSUBS 0.011748f
C519 B.n427 VSUBS 0.011748f
C520 B.n428 VSUBS 0.011748f
C521 B.n429 VSUBS 0.011748f
C522 B.n430 VSUBS 0.011748f
C523 B.n431 VSUBS 0.011748f
C524 B.n432 VSUBS 0.011748f
C525 B.n433 VSUBS 0.011748f
C526 B.n434 VSUBS 0.011748f
C527 B.n435 VSUBS 0.011748f
C528 B.n436 VSUBS 0.011748f
C529 B.n437 VSUBS 0.00812f
C530 B.n438 VSUBS 0.02722f
C531 B.n439 VSUBS 0.009502f
C532 B.n440 VSUBS 0.011748f
C533 B.n441 VSUBS 0.011748f
C534 B.n442 VSUBS 0.011748f
C535 B.n443 VSUBS 0.011748f
C536 B.n444 VSUBS 0.011748f
C537 B.n445 VSUBS 0.011748f
C538 B.n446 VSUBS 0.011748f
C539 B.n447 VSUBS 0.011748f
C540 B.n448 VSUBS 0.011748f
C541 B.n449 VSUBS 0.011748f
C542 B.n450 VSUBS 0.011748f
C543 B.n451 VSUBS 0.009502f
C544 B.n452 VSUBS 0.02722f
C545 B.n453 VSUBS 0.00812f
C546 B.n454 VSUBS 0.011748f
C547 B.n455 VSUBS 0.011748f
C548 B.n456 VSUBS 0.011748f
C549 B.n457 VSUBS 0.011748f
C550 B.n458 VSUBS 0.011748f
C551 B.n459 VSUBS 0.011748f
C552 B.n460 VSUBS 0.011748f
C553 B.n461 VSUBS 0.011748f
C554 B.n462 VSUBS 0.011748f
C555 B.n463 VSUBS 0.011748f
C556 B.n464 VSUBS 0.011748f
C557 B.n465 VSUBS 0.011748f
C558 B.n466 VSUBS 0.011748f
C559 B.n467 VSUBS 0.011748f
C560 B.n468 VSUBS 0.030106f
C561 B.n469 VSUBS 0.030106f
C562 B.n470 VSUBS 0.028981f
C563 B.n471 VSUBS 0.011748f
C564 B.n472 VSUBS 0.011748f
C565 B.n473 VSUBS 0.011748f
C566 B.n474 VSUBS 0.011748f
C567 B.n475 VSUBS 0.011748f
C568 B.n476 VSUBS 0.011748f
C569 B.n477 VSUBS 0.011748f
C570 B.n478 VSUBS 0.011748f
C571 B.n479 VSUBS 0.011748f
C572 B.n480 VSUBS 0.011748f
C573 B.n481 VSUBS 0.011748f
C574 B.n482 VSUBS 0.011748f
C575 B.n483 VSUBS 0.011748f
C576 B.n484 VSUBS 0.011748f
C577 B.n485 VSUBS 0.011748f
C578 B.n486 VSUBS 0.011748f
C579 B.n487 VSUBS 0.011748f
C580 B.n488 VSUBS 0.011748f
C581 B.n489 VSUBS 0.011748f
C582 B.n490 VSUBS 0.011748f
C583 B.n491 VSUBS 0.011748f
C584 B.n492 VSUBS 0.011748f
C585 B.n493 VSUBS 0.011748f
C586 B.n494 VSUBS 0.011748f
C587 B.n495 VSUBS 0.011748f
C588 B.n496 VSUBS 0.011748f
C589 B.n497 VSUBS 0.011748f
C590 B.n498 VSUBS 0.011748f
C591 B.n499 VSUBS 0.011748f
C592 B.n500 VSUBS 0.011748f
C593 B.n501 VSUBS 0.011748f
C594 B.n502 VSUBS 0.011748f
C595 B.n503 VSUBS 0.011748f
C596 B.n504 VSUBS 0.011748f
C597 B.n505 VSUBS 0.011748f
C598 B.n506 VSUBS 0.011748f
C599 B.n507 VSUBS 0.011748f
C600 B.n508 VSUBS 0.011748f
C601 B.n509 VSUBS 0.011748f
C602 B.n510 VSUBS 0.011748f
C603 B.n511 VSUBS 0.011748f
C604 B.n512 VSUBS 0.011748f
C605 B.n513 VSUBS 0.011748f
C606 B.n514 VSUBS 0.011748f
C607 B.n515 VSUBS 0.011748f
C608 B.n516 VSUBS 0.011748f
C609 B.n517 VSUBS 0.011748f
C610 B.n518 VSUBS 0.011748f
C611 B.n519 VSUBS 0.011748f
C612 B.n520 VSUBS 0.011748f
C613 B.n521 VSUBS 0.011748f
C614 B.n522 VSUBS 0.011748f
C615 B.n523 VSUBS 0.011748f
C616 B.n524 VSUBS 0.011748f
C617 B.n525 VSUBS 0.011748f
C618 B.n526 VSUBS 0.011748f
C619 B.n527 VSUBS 0.011748f
C620 B.n528 VSUBS 0.011748f
C621 B.n529 VSUBS 0.011748f
C622 B.n530 VSUBS 0.011748f
C623 B.n531 VSUBS 0.011748f
C624 B.n532 VSUBS 0.011748f
C625 B.n533 VSUBS 0.011748f
C626 B.n534 VSUBS 0.011748f
C627 B.n535 VSUBS 0.011748f
C628 B.n536 VSUBS 0.011748f
C629 B.n537 VSUBS 0.011748f
C630 B.n538 VSUBS 0.011748f
C631 B.n539 VSUBS 0.011748f
C632 B.n540 VSUBS 0.011748f
C633 B.n541 VSUBS 0.011748f
C634 B.n542 VSUBS 0.011748f
C635 B.n543 VSUBS 0.011748f
C636 B.n544 VSUBS 0.011748f
C637 B.n545 VSUBS 0.011748f
C638 B.n546 VSUBS 0.011748f
C639 B.n547 VSUBS 0.026602f
C640 VTAIL.t4 VSUBS 0.046352f
C641 VTAIL.t2 VSUBS 0.046352f
C642 VTAIL.n0 VSUBS 0.146808f
C643 VTAIL.n1 VSUBS 0.689473f
C644 VTAIL.t10 VSUBS 0.254458f
C645 VTAIL.n2 VSUBS 0.987885f
C646 VTAIL.t8 VSUBS 0.046352f
C647 VTAIL.t11 VSUBS 0.046352f
C648 VTAIL.n3 VSUBS 0.146808f
C649 VTAIL.n4 VSUBS 2.15928f
C650 VTAIL.t3 VSUBS 0.046352f
C651 VTAIL.t0 VSUBS 0.046352f
C652 VTAIL.n5 VSUBS 0.146808f
C653 VTAIL.n6 VSUBS 2.15928f
C654 VTAIL.t5 VSUBS 0.254458f
C655 VTAIL.n7 VSUBS 0.987884f
C656 VTAIL.t9 VSUBS 0.046352f
C657 VTAIL.t7 VSUBS 0.046352f
C658 VTAIL.n8 VSUBS 0.146808f
C659 VTAIL.n9 VSUBS 0.969121f
C660 VTAIL.t6 VSUBS 0.254458f
C661 VTAIL.n10 VSUBS 1.79578f
C662 VTAIL.t1 VSUBS 0.254458f
C663 VTAIL.n11 VSUBS 1.69316f
C664 VDD1.t2 VSUBS 0.132954f
C665 VDD1.t1 VSUBS 0.132766f
C666 VDD1.t5 VSUBS 0.021579f
C667 VDD1.t0 VSUBS 0.021579f
C668 VDD1.n0 VSUBS 0.081511f
C669 VDD1.n1 VSUBS 1.93359f
C670 VDD1.t3 VSUBS 0.021579f
C671 VDD1.t4 VSUBS 0.021579f
C672 VDD1.n2 VSUBS 0.080341f
C673 VDD1.n3 VSUBS 1.55498f
C674 VP.t1 VSUBS 0.682601f
C675 VP.n0 VSUBS 0.558511f
C676 VP.n1 VSUBS 0.059629f
C677 VP.n2 VSUBS 0.074039f
C678 VP.n3 VSUBS 0.059629f
C679 VP.t0 VSUBS 0.682601f
C680 VP.n4 VSUBS 0.401053f
C681 VP.n5 VSUBS 0.059629f
C682 VP.n6 VSUBS 0.074039f
C683 VP.n7 VSUBS 0.059629f
C684 VP.t3 VSUBS 0.682601f
C685 VP.n8 VSUBS 0.558511f
C686 VP.t5 VSUBS 0.682601f
C687 VP.n9 VSUBS 0.558511f
C688 VP.n10 VSUBS 0.059629f
C689 VP.n11 VSUBS 0.074039f
C690 VP.n12 VSUBS 0.059629f
C691 VP.t4 VSUBS 0.682601f
C692 VP.n13 VSUBS 0.57955f
C693 VP.t2 VSUBS 1.26234f
C694 VP.n14 VSUBS 0.610017f
C695 VP.n15 VSUBS 0.727087f
C696 VP.n16 VSUBS 0.11169f
C697 VP.n17 VSUBS 0.11169f
C698 VP.n18 VSUBS 0.100813f
C699 VP.n19 VSUBS 0.059629f
C700 VP.n20 VSUBS 0.059629f
C701 VP.n21 VSUBS 0.059629f
C702 VP.n22 VSUBS 0.11169f
C703 VP.n23 VSUBS 0.11169f
C704 VP.n24 VSUBS 0.074191f
C705 VP.n25 VSUBS 0.096255f
C706 VP.n26 VSUBS 2.78261f
C707 VP.n27 VSUBS 2.83158f
C708 VP.n28 VSUBS 0.096255f
C709 VP.n29 VSUBS 0.074191f
C710 VP.n30 VSUBS 0.11169f
C711 VP.n31 VSUBS 0.11169f
C712 VP.n32 VSUBS 0.059629f
C713 VP.n33 VSUBS 0.059629f
C714 VP.n34 VSUBS 0.059629f
C715 VP.n35 VSUBS 0.100813f
C716 VP.n36 VSUBS 0.11169f
C717 VP.n37 VSUBS 0.11169f
C718 VP.n38 VSUBS 0.059629f
C719 VP.n39 VSUBS 0.059629f
C720 VP.n40 VSUBS 0.059629f
C721 VP.n41 VSUBS 0.11169f
C722 VP.n42 VSUBS 0.11169f
C723 VP.n43 VSUBS 0.100813f
C724 VP.n44 VSUBS 0.059629f
C725 VP.n45 VSUBS 0.059629f
C726 VP.n46 VSUBS 0.059629f
C727 VP.n47 VSUBS 0.11169f
C728 VP.n48 VSUBS 0.11169f
C729 VP.n49 VSUBS 0.074191f
C730 VP.n50 VSUBS 0.096255f
C731 VP.n51 VSUBS 0.159663f
.ends

