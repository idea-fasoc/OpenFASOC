* NGSPICE file created from diff_pair_sample_1314.ext - technology: sky130A

.subckt diff_pair_sample_1314 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t5 VP.t0 VTAIL.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=6.6105 pd=34.68 as=2.79675 ps=17.28 w=16.95 l=3.66
X1 B.t19 B.t17 B.t18 B.t11 sky130_fd_pr__nfet_01v8 ad=6.6105 pd=34.68 as=0 ps=0 w=16.95 l=3.66
X2 VTAIL.t7 VP.t1 VDD1.t4 B.t5 sky130_fd_pr__nfet_01v8 ad=2.79675 pd=17.28 as=2.79675 ps=17.28 w=16.95 l=3.66
X3 VDD1.t3 VP.t2 VTAIL.t6 B.t4 sky130_fd_pr__nfet_01v8 ad=2.79675 pd=17.28 as=6.6105 ps=34.68 w=16.95 l=3.66
X4 VTAIL.t10 VP.t3 VDD1.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=2.79675 pd=17.28 as=2.79675 ps=17.28 w=16.95 l=3.66
X5 VDD1.t1 VP.t4 VTAIL.t8 B.t2 sky130_fd_pr__nfet_01v8 ad=2.79675 pd=17.28 as=6.6105 ps=34.68 w=16.95 l=3.66
X6 VDD2.t5 VN.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=6.6105 pd=34.68 as=2.79675 ps=17.28 w=16.95 l=3.66
X7 VTAIL.t1 VN.t1 VDD2.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=2.79675 pd=17.28 as=2.79675 ps=17.28 w=16.95 l=3.66
X8 VDD2.t3 VN.t2 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.79675 pd=17.28 as=6.6105 ps=34.68 w=16.95 l=3.66
X9 VDD2.t2 VN.t3 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=6.6105 pd=34.68 as=2.79675 ps=17.28 w=16.95 l=3.66
X10 VDD2.t1 VN.t4 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=2.79675 pd=17.28 as=6.6105 ps=34.68 w=16.95 l=3.66
X11 B.t16 B.t14 B.t15 B.t7 sky130_fd_pr__nfet_01v8 ad=6.6105 pd=34.68 as=0 ps=0 w=16.95 l=3.66
X12 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=6.6105 pd=34.68 as=0 ps=0 w=16.95 l=3.66
X13 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=6.6105 pd=34.68 as=0 ps=0 w=16.95 l=3.66
X14 VTAIL.t5 VN.t5 VDD2.t0 B.t5 sky130_fd_pr__nfet_01v8 ad=2.79675 pd=17.28 as=2.79675 ps=17.28 w=16.95 l=3.66
X15 VDD1.t0 VP.t5 VTAIL.t9 B.t0 sky130_fd_pr__nfet_01v8 ad=6.6105 pd=34.68 as=2.79675 ps=17.28 w=16.95 l=3.66
R0 VP.n14 VP.n11 161.3
R1 VP.n16 VP.n15 161.3
R2 VP.n17 VP.n10 161.3
R3 VP.n19 VP.n18 161.3
R4 VP.n20 VP.n9 161.3
R5 VP.n22 VP.n21 161.3
R6 VP.n23 VP.n8 161.3
R7 VP.n49 VP.n0 161.3
R8 VP.n48 VP.n47 161.3
R9 VP.n46 VP.n1 161.3
R10 VP.n45 VP.n44 161.3
R11 VP.n43 VP.n2 161.3
R12 VP.n42 VP.n41 161.3
R13 VP.n40 VP.n3 161.3
R14 VP.n39 VP.n38 161.3
R15 VP.n37 VP.n4 161.3
R16 VP.n36 VP.n35 161.3
R17 VP.n34 VP.n5 161.3
R18 VP.n33 VP.n32 161.3
R19 VP.n31 VP.n6 161.3
R20 VP.n30 VP.n29 161.3
R21 VP.n28 VP.n7 161.3
R22 VP.n13 VP.t0 143.768
R23 VP.n38 VP.t1 111.612
R24 VP.n26 VP.t5 111.612
R25 VP.n50 VP.t2 111.612
R26 VP.n12 VP.t3 111.612
R27 VP.n24 VP.t4 111.612
R28 VP.n27 VP.n26 58.2041
R29 VP.n51 VP.n50 58.2041
R30 VP.n25 VP.n24 58.2041
R31 VP.n27 VP.n25 56.8032
R32 VP.n13 VP.n12 50.4706
R33 VP.n32 VP.n5 40.979
R34 VP.n44 VP.n43 40.979
R35 VP.n18 VP.n17 40.979
R36 VP.n32 VP.n31 40.0078
R37 VP.n44 VP.n1 40.0078
R38 VP.n18 VP.n9 40.0078
R39 VP.n30 VP.n7 24.4675
R40 VP.n31 VP.n30 24.4675
R41 VP.n36 VP.n5 24.4675
R42 VP.n37 VP.n36 24.4675
R43 VP.n38 VP.n37 24.4675
R44 VP.n38 VP.n3 24.4675
R45 VP.n42 VP.n3 24.4675
R46 VP.n43 VP.n42 24.4675
R47 VP.n48 VP.n1 24.4675
R48 VP.n49 VP.n48 24.4675
R49 VP.n22 VP.n9 24.4675
R50 VP.n23 VP.n22 24.4675
R51 VP.n12 VP.n11 24.4675
R52 VP.n16 VP.n11 24.4675
R53 VP.n17 VP.n16 24.4675
R54 VP.n26 VP.n7 23.9782
R55 VP.n50 VP.n49 23.9782
R56 VP.n24 VP.n23 23.9782
R57 VP.n14 VP.n13 2.54321
R58 VP.n25 VP.n8 0.417535
R59 VP.n28 VP.n27 0.417535
R60 VP.n51 VP.n0 0.417535
R61 VP VP.n51 0.394291
R62 VP.n15 VP.n14 0.189894
R63 VP.n15 VP.n10 0.189894
R64 VP.n19 VP.n10 0.189894
R65 VP.n20 VP.n19 0.189894
R66 VP.n21 VP.n20 0.189894
R67 VP.n21 VP.n8 0.189894
R68 VP.n29 VP.n28 0.189894
R69 VP.n29 VP.n6 0.189894
R70 VP.n33 VP.n6 0.189894
R71 VP.n34 VP.n33 0.189894
R72 VP.n35 VP.n34 0.189894
R73 VP.n35 VP.n4 0.189894
R74 VP.n39 VP.n4 0.189894
R75 VP.n40 VP.n39 0.189894
R76 VP.n41 VP.n40 0.189894
R77 VP.n41 VP.n2 0.189894
R78 VP.n45 VP.n2 0.189894
R79 VP.n46 VP.n45 0.189894
R80 VP.n47 VP.n46 0.189894
R81 VP.n47 VP.n0 0.189894
R82 VTAIL.n378 VTAIL.n290 289.615
R83 VTAIL.n90 VTAIL.n2 289.615
R84 VTAIL.n284 VTAIL.n196 289.615
R85 VTAIL.n188 VTAIL.n100 289.615
R86 VTAIL.n321 VTAIL.n320 185
R87 VTAIL.n318 VTAIL.n317 185
R88 VTAIL.n327 VTAIL.n326 185
R89 VTAIL.n329 VTAIL.n328 185
R90 VTAIL.n314 VTAIL.n313 185
R91 VTAIL.n335 VTAIL.n334 185
R92 VTAIL.n337 VTAIL.n336 185
R93 VTAIL.n310 VTAIL.n309 185
R94 VTAIL.n343 VTAIL.n342 185
R95 VTAIL.n345 VTAIL.n344 185
R96 VTAIL.n306 VTAIL.n305 185
R97 VTAIL.n351 VTAIL.n350 185
R98 VTAIL.n353 VTAIL.n352 185
R99 VTAIL.n302 VTAIL.n301 185
R100 VTAIL.n359 VTAIL.n358 185
R101 VTAIL.n362 VTAIL.n361 185
R102 VTAIL.n360 VTAIL.n298 185
R103 VTAIL.n367 VTAIL.n297 185
R104 VTAIL.n369 VTAIL.n368 185
R105 VTAIL.n371 VTAIL.n370 185
R106 VTAIL.n294 VTAIL.n293 185
R107 VTAIL.n377 VTAIL.n376 185
R108 VTAIL.n379 VTAIL.n378 185
R109 VTAIL.n33 VTAIL.n32 185
R110 VTAIL.n30 VTAIL.n29 185
R111 VTAIL.n39 VTAIL.n38 185
R112 VTAIL.n41 VTAIL.n40 185
R113 VTAIL.n26 VTAIL.n25 185
R114 VTAIL.n47 VTAIL.n46 185
R115 VTAIL.n49 VTAIL.n48 185
R116 VTAIL.n22 VTAIL.n21 185
R117 VTAIL.n55 VTAIL.n54 185
R118 VTAIL.n57 VTAIL.n56 185
R119 VTAIL.n18 VTAIL.n17 185
R120 VTAIL.n63 VTAIL.n62 185
R121 VTAIL.n65 VTAIL.n64 185
R122 VTAIL.n14 VTAIL.n13 185
R123 VTAIL.n71 VTAIL.n70 185
R124 VTAIL.n74 VTAIL.n73 185
R125 VTAIL.n72 VTAIL.n10 185
R126 VTAIL.n79 VTAIL.n9 185
R127 VTAIL.n81 VTAIL.n80 185
R128 VTAIL.n83 VTAIL.n82 185
R129 VTAIL.n6 VTAIL.n5 185
R130 VTAIL.n89 VTAIL.n88 185
R131 VTAIL.n91 VTAIL.n90 185
R132 VTAIL.n285 VTAIL.n284 185
R133 VTAIL.n283 VTAIL.n282 185
R134 VTAIL.n200 VTAIL.n199 185
R135 VTAIL.n277 VTAIL.n276 185
R136 VTAIL.n275 VTAIL.n274 185
R137 VTAIL.n273 VTAIL.n203 185
R138 VTAIL.n207 VTAIL.n204 185
R139 VTAIL.n268 VTAIL.n267 185
R140 VTAIL.n266 VTAIL.n265 185
R141 VTAIL.n209 VTAIL.n208 185
R142 VTAIL.n260 VTAIL.n259 185
R143 VTAIL.n258 VTAIL.n257 185
R144 VTAIL.n213 VTAIL.n212 185
R145 VTAIL.n252 VTAIL.n251 185
R146 VTAIL.n250 VTAIL.n249 185
R147 VTAIL.n217 VTAIL.n216 185
R148 VTAIL.n244 VTAIL.n243 185
R149 VTAIL.n242 VTAIL.n241 185
R150 VTAIL.n221 VTAIL.n220 185
R151 VTAIL.n236 VTAIL.n235 185
R152 VTAIL.n234 VTAIL.n233 185
R153 VTAIL.n225 VTAIL.n224 185
R154 VTAIL.n228 VTAIL.n227 185
R155 VTAIL.n189 VTAIL.n188 185
R156 VTAIL.n187 VTAIL.n186 185
R157 VTAIL.n104 VTAIL.n103 185
R158 VTAIL.n181 VTAIL.n180 185
R159 VTAIL.n179 VTAIL.n178 185
R160 VTAIL.n177 VTAIL.n107 185
R161 VTAIL.n111 VTAIL.n108 185
R162 VTAIL.n172 VTAIL.n171 185
R163 VTAIL.n170 VTAIL.n169 185
R164 VTAIL.n113 VTAIL.n112 185
R165 VTAIL.n164 VTAIL.n163 185
R166 VTAIL.n162 VTAIL.n161 185
R167 VTAIL.n117 VTAIL.n116 185
R168 VTAIL.n156 VTAIL.n155 185
R169 VTAIL.n154 VTAIL.n153 185
R170 VTAIL.n121 VTAIL.n120 185
R171 VTAIL.n148 VTAIL.n147 185
R172 VTAIL.n146 VTAIL.n145 185
R173 VTAIL.n125 VTAIL.n124 185
R174 VTAIL.n140 VTAIL.n139 185
R175 VTAIL.n138 VTAIL.n137 185
R176 VTAIL.n129 VTAIL.n128 185
R177 VTAIL.n132 VTAIL.n131 185
R178 VTAIL.t8 VTAIL.n226 147.659
R179 VTAIL.t4 VTAIL.n130 147.659
R180 VTAIL.t2 VTAIL.n319 147.659
R181 VTAIL.t6 VTAIL.n31 147.659
R182 VTAIL.n320 VTAIL.n317 104.615
R183 VTAIL.n327 VTAIL.n317 104.615
R184 VTAIL.n328 VTAIL.n327 104.615
R185 VTAIL.n328 VTAIL.n313 104.615
R186 VTAIL.n335 VTAIL.n313 104.615
R187 VTAIL.n336 VTAIL.n335 104.615
R188 VTAIL.n336 VTAIL.n309 104.615
R189 VTAIL.n343 VTAIL.n309 104.615
R190 VTAIL.n344 VTAIL.n343 104.615
R191 VTAIL.n344 VTAIL.n305 104.615
R192 VTAIL.n351 VTAIL.n305 104.615
R193 VTAIL.n352 VTAIL.n351 104.615
R194 VTAIL.n352 VTAIL.n301 104.615
R195 VTAIL.n359 VTAIL.n301 104.615
R196 VTAIL.n361 VTAIL.n359 104.615
R197 VTAIL.n361 VTAIL.n360 104.615
R198 VTAIL.n360 VTAIL.n297 104.615
R199 VTAIL.n369 VTAIL.n297 104.615
R200 VTAIL.n370 VTAIL.n369 104.615
R201 VTAIL.n370 VTAIL.n293 104.615
R202 VTAIL.n377 VTAIL.n293 104.615
R203 VTAIL.n378 VTAIL.n377 104.615
R204 VTAIL.n32 VTAIL.n29 104.615
R205 VTAIL.n39 VTAIL.n29 104.615
R206 VTAIL.n40 VTAIL.n39 104.615
R207 VTAIL.n40 VTAIL.n25 104.615
R208 VTAIL.n47 VTAIL.n25 104.615
R209 VTAIL.n48 VTAIL.n47 104.615
R210 VTAIL.n48 VTAIL.n21 104.615
R211 VTAIL.n55 VTAIL.n21 104.615
R212 VTAIL.n56 VTAIL.n55 104.615
R213 VTAIL.n56 VTAIL.n17 104.615
R214 VTAIL.n63 VTAIL.n17 104.615
R215 VTAIL.n64 VTAIL.n63 104.615
R216 VTAIL.n64 VTAIL.n13 104.615
R217 VTAIL.n71 VTAIL.n13 104.615
R218 VTAIL.n73 VTAIL.n71 104.615
R219 VTAIL.n73 VTAIL.n72 104.615
R220 VTAIL.n72 VTAIL.n9 104.615
R221 VTAIL.n81 VTAIL.n9 104.615
R222 VTAIL.n82 VTAIL.n81 104.615
R223 VTAIL.n82 VTAIL.n5 104.615
R224 VTAIL.n89 VTAIL.n5 104.615
R225 VTAIL.n90 VTAIL.n89 104.615
R226 VTAIL.n284 VTAIL.n283 104.615
R227 VTAIL.n283 VTAIL.n199 104.615
R228 VTAIL.n276 VTAIL.n199 104.615
R229 VTAIL.n276 VTAIL.n275 104.615
R230 VTAIL.n275 VTAIL.n203 104.615
R231 VTAIL.n207 VTAIL.n203 104.615
R232 VTAIL.n267 VTAIL.n207 104.615
R233 VTAIL.n267 VTAIL.n266 104.615
R234 VTAIL.n266 VTAIL.n208 104.615
R235 VTAIL.n259 VTAIL.n208 104.615
R236 VTAIL.n259 VTAIL.n258 104.615
R237 VTAIL.n258 VTAIL.n212 104.615
R238 VTAIL.n251 VTAIL.n212 104.615
R239 VTAIL.n251 VTAIL.n250 104.615
R240 VTAIL.n250 VTAIL.n216 104.615
R241 VTAIL.n243 VTAIL.n216 104.615
R242 VTAIL.n243 VTAIL.n242 104.615
R243 VTAIL.n242 VTAIL.n220 104.615
R244 VTAIL.n235 VTAIL.n220 104.615
R245 VTAIL.n235 VTAIL.n234 104.615
R246 VTAIL.n234 VTAIL.n224 104.615
R247 VTAIL.n227 VTAIL.n224 104.615
R248 VTAIL.n188 VTAIL.n187 104.615
R249 VTAIL.n187 VTAIL.n103 104.615
R250 VTAIL.n180 VTAIL.n103 104.615
R251 VTAIL.n180 VTAIL.n179 104.615
R252 VTAIL.n179 VTAIL.n107 104.615
R253 VTAIL.n111 VTAIL.n107 104.615
R254 VTAIL.n171 VTAIL.n111 104.615
R255 VTAIL.n171 VTAIL.n170 104.615
R256 VTAIL.n170 VTAIL.n112 104.615
R257 VTAIL.n163 VTAIL.n112 104.615
R258 VTAIL.n163 VTAIL.n162 104.615
R259 VTAIL.n162 VTAIL.n116 104.615
R260 VTAIL.n155 VTAIL.n116 104.615
R261 VTAIL.n155 VTAIL.n154 104.615
R262 VTAIL.n154 VTAIL.n120 104.615
R263 VTAIL.n147 VTAIL.n120 104.615
R264 VTAIL.n147 VTAIL.n146 104.615
R265 VTAIL.n146 VTAIL.n124 104.615
R266 VTAIL.n139 VTAIL.n124 104.615
R267 VTAIL.n139 VTAIL.n138 104.615
R268 VTAIL.n138 VTAIL.n128 104.615
R269 VTAIL.n131 VTAIL.n128 104.615
R270 VTAIL.n320 VTAIL.t2 52.3082
R271 VTAIL.n32 VTAIL.t6 52.3082
R272 VTAIL.n227 VTAIL.t8 52.3082
R273 VTAIL.n131 VTAIL.t4 52.3082
R274 VTAIL.n195 VTAIL.n194 46.9551
R275 VTAIL.n99 VTAIL.n98 46.9551
R276 VTAIL.n1 VTAIL.n0 46.9549
R277 VTAIL.n97 VTAIL.n96 46.9549
R278 VTAIL.n383 VTAIL.n382 35.0944
R279 VTAIL.n95 VTAIL.n94 35.0944
R280 VTAIL.n289 VTAIL.n288 35.0944
R281 VTAIL.n193 VTAIL.n192 35.0944
R282 VTAIL.n99 VTAIL.n97 33.8583
R283 VTAIL.n383 VTAIL.n289 30.4186
R284 VTAIL.n321 VTAIL.n319 15.6677
R285 VTAIL.n33 VTAIL.n31 15.6677
R286 VTAIL.n228 VTAIL.n226 15.6677
R287 VTAIL.n132 VTAIL.n130 15.6677
R288 VTAIL.n368 VTAIL.n367 13.1884
R289 VTAIL.n80 VTAIL.n79 13.1884
R290 VTAIL.n274 VTAIL.n273 13.1884
R291 VTAIL.n178 VTAIL.n177 13.1884
R292 VTAIL.n322 VTAIL.n318 12.8005
R293 VTAIL.n366 VTAIL.n298 12.8005
R294 VTAIL.n371 VTAIL.n296 12.8005
R295 VTAIL.n34 VTAIL.n30 12.8005
R296 VTAIL.n78 VTAIL.n10 12.8005
R297 VTAIL.n83 VTAIL.n8 12.8005
R298 VTAIL.n277 VTAIL.n202 12.8005
R299 VTAIL.n272 VTAIL.n204 12.8005
R300 VTAIL.n229 VTAIL.n225 12.8005
R301 VTAIL.n181 VTAIL.n106 12.8005
R302 VTAIL.n176 VTAIL.n108 12.8005
R303 VTAIL.n133 VTAIL.n129 12.8005
R304 VTAIL.n326 VTAIL.n325 12.0247
R305 VTAIL.n363 VTAIL.n362 12.0247
R306 VTAIL.n372 VTAIL.n294 12.0247
R307 VTAIL.n38 VTAIL.n37 12.0247
R308 VTAIL.n75 VTAIL.n74 12.0247
R309 VTAIL.n84 VTAIL.n6 12.0247
R310 VTAIL.n278 VTAIL.n200 12.0247
R311 VTAIL.n269 VTAIL.n268 12.0247
R312 VTAIL.n233 VTAIL.n232 12.0247
R313 VTAIL.n182 VTAIL.n104 12.0247
R314 VTAIL.n173 VTAIL.n172 12.0247
R315 VTAIL.n137 VTAIL.n136 12.0247
R316 VTAIL.n329 VTAIL.n316 11.249
R317 VTAIL.n358 VTAIL.n300 11.249
R318 VTAIL.n376 VTAIL.n375 11.249
R319 VTAIL.n41 VTAIL.n28 11.249
R320 VTAIL.n70 VTAIL.n12 11.249
R321 VTAIL.n88 VTAIL.n87 11.249
R322 VTAIL.n282 VTAIL.n281 11.249
R323 VTAIL.n265 VTAIL.n206 11.249
R324 VTAIL.n236 VTAIL.n223 11.249
R325 VTAIL.n186 VTAIL.n185 11.249
R326 VTAIL.n169 VTAIL.n110 11.249
R327 VTAIL.n140 VTAIL.n127 11.249
R328 VTAIL.n330 VTAIL.n314 10.4732
R329 VTAIL.n357 VTAIL.n302 10.4732
R330 VTAIL.n379 VTAIL.n292 10.4732
R331 VTAIL.n42 VTAIL.n26 10.4732
R332 VTAIL.n69 VTAIL.n14 10.4732
R333 VTAIL.n91 VTAIL.n4 10.4732
R334 VTAIL.n285 VTAIL.n198 10.4732
R335 VTAIL.n264 VTAIL.n209 10.4732
R336 VTAIL.n237 VTAIL.n221 10.4732
R337 VTAIL.n189 VTAIL.n102 10.4732
R338 VTAIL.n168 VTAIL.n113 10.4732
R339 VTAIL.n141 VTAIL.n125 10.4732
R340 VTAIL.n334 VTAIL.n333 9.69747
R341 VTAIL.n354 VTAIL.n353 9.69747
R342 VTAIL.n380 VTAIL.n290 9.69747
R343 VTAIL.n46 VTAIL.n45 9.69747
R344 VTAIL.n66 VTAIL.n65 9.69747
R345 VTAIL.n92 VTAIL.n2 9.69747
R346 VTAIL.n286 VTAIL.n196 9.69747
R347 VTAIL.n261 VTAIL.n260 9.69747
R348 VTAIL.n241 VTAIL.n240 9.69747
R349 VTAIL.n190 VTAIL.n100 9.69747
R350 VTAIL.n165 VTAIL.n164 9.69747
R351 VTAIL.n145 VTAIL.n144 9.69747
R352 VTAIL.n382 VTAIL.n381 9.45567
R353 VTAIL.n94 VTAIL.n93 9.45567
R354 VTAIL.n288 VTAIL.n287 9.45567
R355 VTAIL.n192 VTAIL.n191 9.45567
R356 VTAIL.n381 VTAIL.n380 9.3005
R357 VTAIL.n292 VTAIL.n291 9.3005
R358 VTAIL.n375 VTAIL.n374 9.3005
R359 VTAIL.n373 VTAIL.n372 9.3005
R360 VTAIL.n296 VTAIL.n295 9.3005
R361 VTAIL.n341 VTAIL.n340 9.3005
R362 VTAIL.n339 VTAIL.n338 9.3005
R363 VTAIL.n312 VTAIL.n311 9.3005
R364 VTAIL.n333 VTAIL.n332 9.3005
R365 VTAIL.n331 VTAIL.n330 9.3005
R366 VTAIL.n316 VTAIL.n315 9.3005
R367 VTAIL.n325 VTAIL.n324 9.3005
R368 VTAIL.n323 VTAIL.n322 9.3005
R369 VTAIL.n308 VTAIL.n307 9.3005
R370 VTAIL.n347 VTAIL.n346 9.3005
R371 VTAIL.n349 VTAIL.n348 9.3005
R372 VTAIL.n304 VTAIL.n303 9.3005
R373 VTAIL.n355 VTAIL.n354 9.3005
R374 VTAIL.n357 VTAIL.n356 9.3005
R375 VTAIL.n300 VTAIL.n299 9.3005
R376 VTAIL.n364 VTAIL.n363 9.3005
R377 VTAIL.n366 VTAIL.n365 9.3005
R378 VTAIL.n93 VTAIL.n92 9.3005
R379 VTAIL.n4 VTAIL.n3 9.3005
R380 VTAIL.n87 VTAIL.n86 9.3005
R381 VTAIL.n85 VTAIL.n84 9.3005
R382 VTAIL.n8 VTAIL.n7 9.3005
R383 VTAIL.n53 VTAIL.n52 9.3005
R384 VTAIL.n51 VTAIL.n50 9.3005
R385 VTAIL.n24 VTAIL.n23 9.3005
R386 VTAIL.n45 VTAIL.n44 9.3005
R387 VTAIL.n43 VTAIL.n42 9.3005
R388 VTAIL.n28 VTAIL.n27 9.3005
R389 VTAIL.n37 VTAIL.n36 9.3005
R390 VTAIL.n35 VTAIL.n34 9.3005
R391 VTAIL.n20 VTAIL.n19 9.3005
R392 VTAIL.n59 VTAIL.n58 9.3005
R393 VTAIL.n61 VTAIL.n60 9.3005
R394 VTAIL.n16 VTAIL.n15 9.3005
R395 VTAIL.n67 VTAIL.n66 9.3005
R396 VTAIL.n69 VTAIL.n68 9.3005
R397 VTAIL.n12 VTAIL.n11 9.3005
R398 VTAIL.n76 VTAIL.n75 9.3005
R399 VTAIL.n78 VTAIL.n77 9.3005
R400 VTAIL.n254 VTAIL.n253 9.3005
R401 VTAIL.n256 VTAIL.n255 9.3005
R402 VTAIL.n211 VTAIL.n210 9.3005
R403 VTAIL.n262 VTAIL.n261 9.3005
R404 VTAIL.n264 VTAIL.n263 9.3005
R405 VTAIL.n206 VTAIL.n205 9.3005
R406 VTAIL.n270 VTAIL.n269 9.3005
R407 VTAIL.n272 VTAIL.n271 9.3005
R408 VTAIL.n287 VTAIL.n286 9.3005
R409 VTAIL.n198 VTAIL.n197 9.3005
R410 VTAIL.n281 VTAIL.n280 9.3005
R411 VTAIL.n279 VTAIL.n278 9.3005
R412 VTAIL.n202 VTAIL.n201 9.3005
R413 VTAIL.n215 VTAIL.n214 9.3005
R414 VTAIL.n248 VTAIL.n247 9.3005
R415 VTAIL.n246 VTAIL.n245 9.3005
R416 VTAIL.n219 VTAIL.n218 9.3005
R417 VTAIL.n240 VTAIL.n239 9.3005
R418 VTAIL.n238 VTAIL.n237 9.3005
R419 VTAIL.n223 VTAIL.n222 9.3005
R420 VTAIL.n232 VTAIL.n231 9.3005
R421 VTAIL.n230 VTAIL.n229 9.3005
R422 VTAIL.n158 VTAIL.n157 9.3005
R423 VTAIL.n160 VTAIL.n159 9.3005
R424 VTAIL.n115 VTAIL.n114 9.3005
R425 VTAIL.n166 VTAIL.n165 9.3005
R426 VTAIL.n168 VTAIL.n167 9.3005
R427 VTAIL.n110 VTAIL.n109 9.3005
R428 VTAIL.n174 VTAIL.n173 9.3005
R429 VTAIL.n176 VTAIL.n175 9.3005
R430 VTAIL.n191 VTAIL.n190 9.3005
R431 VTAIL.n102 VTAIL.n101 9.3005
R432 VTAIL.n185 VTAIL.n184 9.3005
R433 VTAIL.n183 VTAIL.n182 9.3005
R434 VTAIL.n106 VTAIL.n105 9.3005
R435 VTAIL.n119 VTAIL.n118 9.3005
R436 VTAIL.n152 VTAIL.n151 9.3005
R437 VTAIL.n150 VTAIL.n149 9.3005
R438 VTAIL.n123 VTAIL.n122 9.3005
R439 VTAIL.n144 VTAIL.n143 9.3005
R440 VTAIL.n142 VTAIL.n141 9.3005
R441 VTAIL.n127 VTAIL.n126 9.3005
R442 VTAIL.n136 VTAIL.n135 9.3005
R443 VTAIL.n134 VTAIL.n133 9.3005
R444 VTAIL.n337 VTAIL.n312 8.92171
R445 VTAIL.n350 VTAIL.n304 8.92171
R446 VTAIL.n49 VTAIL.n24 8.92171
R447 VTAIL.n62 VTAIL.n16 8.92171
R448 VTAIL.n257 VTAIL.n211 8.92171
R449 VTAIL.n244 VTAIL.n219 8.92171
R450 VTAIL.n161 VTAIL.n115 8.92171
R451 VTAIL.n148 VTAIL.n123 8.92171
R452 VTAIL.n338 VTAIL.n310 8.14595
R453 VTAIL.n349 VTAIL.n306 8.14595
R454 VTAIL.n50 VTAIL.n22 8.14595
R455 VTAIL.n61 VTAIL.n18 8.14595
R456 VTAIL.n256 VTAIL.n213 8.14595
R457 VTAIL.n245 VTAIL.n217 8.14595
R458 VTAIL.n160 VTAIL.n117 8.14595
R459 VTAIL.n149 VTAIL.n121 8.14595
R460 VTAIL.n342 VTAIL.n341 7.3702
R461 VTAIL.n346 VTAIL.n345 7.3702
R462 VTAIL.n54 VTAIL.n53 7.3702
R463 VTAIL.n58 VTAIL.n57 7.3702
R464 VTAIL.n253 VTAIL.n252 7.3702
R465 VTAIL.n249 VTAIL.n248 7.3702
R466 VTAIL.n157 VTAIL.n156 7.3702
R467 VTAIL.n153 VTAIL.n152 7.3702
R468 VTAIL.n342 VTAIL.n308 6.59444
R469 VTAIL.n345 VTAIL.n308 6.59444
R470 VTAIL.n54 VTAIL.n20 6.59444
R471 VTAIL.n57 VTAIL.n20 6.59444
R472 VTAIL.n252 VTAIL.n215 6.59444
R473 VTAIL.n249 VTAIL.n215 6.59444
R474 VTAIL.n156 VTAIL.n119 6.59444
R475 VTAIL.n153 VTAIL.n119 6.59444
R476 VTAIL.n341 VTAIL.n310 5.81868
R477 VTAIL.n346 VTAIL.n306 5.81868
R478 VTAIL.n53 VTAIL.n22 5.81868
R479 VTAIL.n58 VTAIL.n18 5.81868
R480 VTAIL.n253 VTAIL.n213 5.81868
R481 VTAIL.n248 VTAIL.n217 5.81868
R482 VTAIL.n157 VTAIL.n117 5.81868
R483 VTAIL.n152 VTAIL.n121 5.81868
R484 VTAIL.n338 VTAIL.n337 5.04292
R485 VTAIL.n350 VTAIL.n349 5.04292
R486 VTAIL.n50 VTAIL.n49 5.04292
R487 VTAIL.n62 VTAIL.n61 5.04292
R488 VTAIL.n257 VTAIL.n256 5.04292
R489 VTAIL.n245 VTAIL.n244 5.04292
R490 VTAIL.n161 VTAIL.n160 5.04292
R491 VTAIL.n149 VTAIL.n148 5.04292
R492 VTAIL.n230 VTAIL.n226 4.38563
R493 VTAIL.n134 VTAIL.n130 4.38563
R494 VTAIL.n323 VTAIL.n319 4.38563
R495 VTAIL.n35 VTAIL.n31 4.38563
R496 VTAIL.n334 VTAIL.n312 4.26717
R497 VTAIL.n353 VTAIL.n304 4.26717
R498 VTAIL.n382 VTAIL.n290 4.26717
R499 VTAIL.n46 VTAIL.n24 4.26717
R500 VTAIL.n65 VTAIL.n16 4.26717
R501 VTAIL.n94 VTAIL.n2 4.26717
R502 VTAIL.n288 VTAIL.n196 4.26717
R503 VTAIL.n260 VTAIL.n211 4.26717
R504 VTAIL.n241 VTAIL.n219 4.26717
R505 VTAIL.n192 VTAIL.n100 4.26717
R506 VTAIL.n164 VTAIL.n115 4.26717
R507 VTAIL.n145 VTAIL.n123 4.26717
R508 VTAIL.n333 VTAIL.n314 3.49141
R509 VTAIL.n354 VTAIL.n302 3.49141
R510 VTAIL.n380 VTAIL.n379 3.49141
R511 VTAIL.n45 VTAIL.n26 3.49141
R512 VTAIL.n66 VTAIL.n14 3.49141
R513 VTAIL.n92 VTAIL.n91 3.49141
R514 VTAIL.n286 VTAIL.n285 3.49141
R515 VTAIL.n261 VTAIL.n209 3.49141
R516 VTAIL.n240 VTAIL.n221 3.49141
R517 VTAIL.n190 VTAIL.n189 3.49141
R518 VTAIL.n165 VTAIL.n113 3.49141
R519 VTAIL.n144 VTAIL.n125 3.49141
R520 VTAIL.n193 VTAIL.n99 3.44016
R521 VTAIL.n289 VTAIL.n195 3.44016
R522 VTAIL.n97 VTAIL.n95 3.44016
R523 VTAIL.n330 VTAIL.n329 2.71565
R524 VTAIL.n358 VTAIL.n357 2.71565
R525 VTAIL.n376 VTAIL.n292 2.71565
R526 VTAIL.n42 VTAIL.n41 2.71565
R527 VTAIL.n70 VTAIL.n69 2.71565
R528 VTAIL.n88 VTAIL.n4 2.71565
R529 VTAIL.n282 VTAIL.n198 2.71565
R530 VTAIL.n265 VTAIL.n264 2.71565
R531 VTAIL.n237 VTAIL.n236 2.71565
R532 VTAIL.n186 VTAIL.n102 2.71565
R533 VTAIL.n169 VTAIL.n168 2.71565
R534 VTAIL.n141 VTAIL.n140 2.71565
R535 VTAIL VTAIL.n383 2.52205
R536 VTAIL.n195 VTAIL.n193 2.19016
R537 VTAIL.n95 VTAIL.n1 2.19016
R538 VTAIL.n326 VTAIL.n316 1.93989
R539 VTAIL.n362 VTAIL.n300 1.93989
R540 VTAIL.n375 VTAIL.n294 1.93989
R541 VTAIL.n38 VTAIL.n28 1.93989
R542 VTAIL.n74 VTAIL.n12 1.93989
R543 VTAIL.n87 VTAIL.n6 1.93989
R544 VTAIL.n281 VTAIL.n200 1.93989
R545 VTAIL.n268 VTAIL.n206 1.93989
R546 VTAIL.n233 VTAIL.n223 1.93989
R547 VTAIL.n185 VTAIL.n104 1.93989
R548 VTAIL.n172 VTAIL.n110 1.93989
R549 VTAIL.n137 VTAIL.n127 1.93989
R550 VTAIL.n0 VTAIL.t3 1.16864
R551 VTAIL.n0 VTAIL.t1 1.16864
R552 VTAIL.n96 VTAIL.t9 1.16864
R553 VTAIL.n96 VTAIL.t7 1.16864
R554 VTAIL.n194 VTAIL.t11 1.16864
R555 VTAIL.n194 VTAIL.t10 1.16864
R556 VTAIL.n98 VTAIL.t0 1.16864
R557 VTAIL.n98 VTAIL.t5 1.16864
R558 VTAIL.n325 VTAIL.n318 1.16414
R559 VTAIL.n363 VTAIL.n298 1.16414
R560 VTAIL.n372 VTAIL.n371 1.16414
R561 VTAIL.n37 VTAIL.n30 1.16414
R562 VTAIL.n75 VTAIL.n10 1.16414
R563 VTAIL.n84 VTAIL.n83 1.16414
R564 VTAIL.n278 VTAIL.n277 1.16414
R565 VTAIL.n269 VTAIL.n204 1.16414
R566 VTAIL.n232 VTAIL.n225 1.16414
R567 VTAIL.n182 VTAIL.n181 1.16414
R568 VTAIL.n173 VTAIL.n108 1.16414
R569 VTAIL.n136 VTAIL.n129 1.16414
R570 VTAIL VTAIL.n1 0.918603
R571 VTAIL.n322 VTAIL.n321 0.388379
R572 VTAIL.n367 VTAIL.n366 0.388379
R573 VTAIL.n368 VTAIL.n296 0.388379
R574 VTAIL.n34 VTAIL.n33 0.388379
R575 VTAIL.n79 VTAIL.n78 0.388379
R576 VTAIL.n80 VTAIL.n8 0.388379
R577 VTAIL.n274 VTAIL.n202 0.388379
R578 VTAIL.n273 VTAIL.n272 0.388379
R579 VTAIL.n229 VTAIL.n228 0.388379
R580 VTAIL.n178 VTAIL.n106 0.388379
R581 VTAIL.n177 VTAIL.n176 0.388379
R582 VTAIL.n133 VTAIL.n132 0.388379
R583 VTAIL.n324 VTAIL.n323 0.155672
R584 VTAIL.n324 VTAIL.n315 0.155672
R585 VTAIL.n331 VTAIL.n315 0.155672
R586 VTAIL.n332 VTAIL.n331 0.155672
R587 VTAIL.n332 VTAIL.n311 0.155672
R588 VTAIL.n339 VTAIL.n311 0.155672
R589 VTAIL.n340 VTAIL.n339 0.155672
R590 VTAIL.n340 VTAIL.n307 0.155672
R591 VTAIL.n347 VTAIL.n307 0.155672
R592 VTAIL.n348 VTAIL.n347 0.155672
R593 VTAIL.n348 VTAIL.n303 0.155672
R594 VTAIL.n355 VTAIL.n303 0.155672
R595 VTAIL.n356 VTAIL.n355 0.155672
R596 VTAIL.n356 VTAIL.n299 0.155672
R597 VTAIL.n364 VTAIL.n299 0.155672
R598 VTAIL.n365 VTAIL.n364 0.155672
R599 VTAIL.n365 VTAIL.n295 0.155672
R600 VTAIL.n373 VTAIL.n295 0.155672
R601 VTAIL.n374 VTAIL.n373 0.155672
R602 VTAIL.n374 VTAIL.n291 0.155672
R603 VTAIL.n381 VTAIL.n291 0.155672
R604 VTAIL.n36 VTAIL.n35 0.155672
R605 VTAIL.n36 VTAIL.n27 0.155672
R606 VTAIL.n43 VTAIL.n27 0.155672
R607 VTAIL.n44 VTAIL.n43 0.155672
R608 VTAIL.n44 VTAIL.n23 0.155672
R609 VTAIL.n51 VTAIL.n23 0.155672
R610 VTAIL.n52 VTAIL.n51 0.155672
R611 VTAIL.n52 VTAIL.n19 0.155672
R612 VTAIL.n59 VTAIL.n19 0.155672
R613 VTAIL.n60 VTAIL.n59 0.155672
R614 VTAIL.n60 VTAIL.n15 0.155672
R615 VTAIL.n67 VTAIL.n15 0.155672
R616 VTAIL.n68 VTAIL.n67 0.155672
R617 VTAIL.n68 VTAIL.n11 0.155672
R618 VTAIL.n76 VTAIL.n11 0.155672
R619 VTAIL.n77 VTAIL.n76 0.155672
R620 VTAIL.n77 VTAIL.n7 0.155672
R621 VTAIL.n85 VTAIL.n7 0.155672
R622 VTAIL.n86 VTAIL.n85 0.155672
R623 VTAIL.n86 VTAIL.n3 0.155672
R624 VTAIL.n93 VTAIL.n3 0.155672
R625 VTAIL.n287 VTAIL.n197 0.155672
R626 VTAIL.n280 VTAIL.n197 0.155672
R627 VTAIL.n280 VTAIL.n279 0.155672
R628 VTAIL.n279 VTAIL.n201 0.155672
R629 VTAIL.n271 VTAIL.n201 0.155672
R630 VTAIL.n271 VTAIL.n270 0.155672
R631 VTAIL.n270 VTAIL.n205 0.155672
R632 VTAIL.n263 VTAIL.n205 0.155672
R633 VTAIL.n263 VTAIL.n262 0.155672
R634 VTAIL.n262 VTAIL.n210 0.155672
R635 VTAIL.n255 VTAIL.n210 0.155672
R636 VTAIL.n255 VTAIL.n254 0.155672
R637 VTAIL.n254 VTAIL.n214 0.155672
R638 VTAIL.n247 VTAIL.n214 0.155672
R639 VTAIL.n247 VTAIL.n246 0.155672
R640 VTAIL.n246 VTAIL.n218 0.155672
R641 VTAIL.n239 VTAIL.n218 0.155672
R642 VTAIL.n239 VTAIL.n238 0.155672
R643 VTAIL.n238 VTAIL.n222 0.155672
R644 VTAIL.n231 VTAIL.n222 0.155672
R645 VTAIL.n231 VTAIL.n230 0.155672
R646 VTAIL.n191 VTAIL.n101 0.155672
R647 VTAIL.n184 VTAIL.n101 0.155672
R648 VTAIL.n184 VTAIL.n183 0.155672
R649 VTAIL.n183 VTAIL.n105 0.155672
R650 VTAIL.n175 VTAIL.n105 0.155672
R651 VTAIL.n175 VTAIL.n174 0.155672
R652 VTAIL.n174 VTAIL.n109 0.155672
R653 VTAIL.n167 VTAIL.n109 0.155672
R654 VTAIL.n167 VTAIL.n166 0.155672
R655 VTAIL.n166 VTAIL.n114 0.155672
R656 VTAIL.n159 VTAIL.n114 0.155672
R657 VTAIL.n159 VTAIL.n158 0.155672
R658 VTAIL.n158 VTAIL.n118 0.155672
R659 VTAIL.n151 VTAIL.n118 0.155672
R660 VTAIL.n151 VTAIL.n150 0.155672
R661 VTAIL.n150 VTAIL.n122 0.155672
R662 VTAIL.n143 VTAIL.n122 0.155672
R663 VTAIL.n143 VTAIL.n142 0.155672
R664 VTAIL.n142 VTAIL.n126 0.155672
R665 VTAIL.n135 VTAIL.n126 0.155672
R666 VTAIL.n135 VTAIL.n134 0.155672
R667 VDD1.n88 VDD1.n0 289.615
R668 VDD1.n181 VDD1.n93 289.615
R669 VDD1.n89 VDD1.n88 185
R670 VDD1.n87 VDD1.n86 185
R671 VDD1.n4 VDD1.n3 185
R672 VDD1.n81 VDD1.n80 185
R673 VDD1.n79 VDD1.n78 185
R674 VDD1.n77 VDD1.n7 185
R675 VDD1.n11 VDD1.n8 185
R676 VDD1.n72 VDD1.n71 185
R677 VDD1.n70 VDD1.n69 185
R678 VDD1.n13 VDD1.n12 185
R679 VDD1.n64 VDD1.n63 185
R680 VDD1.n62 VDD1.n61 185
R681 VDD1.n17 VDD1.n16 185
R682 VDD1.n56 VDD1.n55 185
R683 VDD1.n54 VDD1.n53 185
R684 VDD1.n21 VDD1.n20 185
R685 VDD1.n48 VDD1.n47 185
R686 VDD1.n46 VDD1.n45 185
R687 VDD1.n25 VDD1.n24 185
R688 VDD1.n40 VDD1.n39 185
R689 VDD1.n38 VDD1.n37 185
R690 VDD1.n29 VDD1.n28 185
R691 VDD1.n32 VDD1.n31 185
R692 VDD1.n124 VDD1.n123 185
R693 VDD1.n121 VDD1.n120 185
R694 VDD1.n130 VDD1.n129 185
R695 VDD1.n132 VDD1.n131 185
R696 VDD1.n117 VDD1.n116 185
R697 VDD1.n138 VDD1.n137 185
R698 VDD1.n140 VDD1.n139 185
R699 VDD1.n113 VDD1.n112 185
R700 VDD1.n146 VDD1.n145 185
R701 VDD1.n148 VDD1.n147 185
R702 VDD1.n109 VDD1.n108 185
R703 VDD1.n154 VDD1.n153 185
R704 VDD1.n156 VDD1.n155 185
R705 VDD1.n105 VDD1.n104 185
R706 VDD1.n162 VDD1.n161 185
R707 VDD1.n165 VDD1.n164 185
R708 VDD1.n163 VDD1.n101 185
R709 VDD1.n170 VDD1.n100 185
R710 VDD1.n172 VDD1.n171 185
R711 VDD1.n174 VDD1.n173 185
R712 VDD1.n97 VDD1.n96 185
R713 VDD1.n180 VDD1.n179 185
R714 VDD1.n182 VDD1.n181 185
R715 VDD1.t5 VDD1.n30 147.659
R716 VDD1.t0 VDD1.n122 147.659
R717 VDD1.n88 VDD1.n87 104.615
R718 VDD1.n87 VDD1.n3 104.615
R719 VDD1.n80 VDD1.n3 104.615
R720 VDD1.n80 VDD1.n79 104.615
R721 VDD1.n79 VDD1.n7 104.615
R722 VDD1.n11 VDD1.n7 104.615
R723 VDD1.n71 VDD1.n11 104.615
R724 VDD1.n71 VDD1.n70 104.615
R725 VDD1.n70 VDD1.n12 104.615
R726 VDD1.n63 VDD1.n12 104.615
R727 VDD1.n63 VDD1.n62 104.615
R728 VDD1.n62 VDD1.n16 104.615
R729 VDD1.n55 VDD1.n16 104.615
R730 VDD1.n55 VDD1.n54 104.615
R731 VDD1.n54 VDD1.n20 104.615
R732 VDD1.n47 VDD1.n20 104.615
R733 VDD1.n47 VDD1.n46 104.615
R734 VDD1.n46 VDD1.n24 104.615
R735 VDD1.n39 VDD1.n24 104.615
R736 VDD1.n39 VDD1.n38 104.615
R737 VDD1.n38 VDD1.n28 104.615
R738 VDD1.n31 VDD1.n28 104.615
R739 VDD1.n123 VDD1.n120 104.615
R740 VDD1.n130 VDD1.n120 104.615
R741 VDD1.n131 VDD1.n130 104.615
R742 VDD1.n131 VDD1.n116 104.615
R743 VDD1.n138 VDD1.n116 104.615
R744 VDD1.n139 VDD1.n138 104.615
R745 VDD1.n139 VDD1.n112 104.615
R746 VDD1.n146 VDD1.n112 104.615
R747 VDD1.n147 VDD1.n146 104.615
R748 VDD1.n147 VDD1.n108 104.615
R749 VDD1.n154 VDD1.n108 104.615
R750 VDD1.n155 VDD1.n154 104.615
R751 VDD1.n155 VDD1.n104 104.615
R752 VDD1.n162 VDD1.n104 104.615
R753 VDD1.n164 VDD1.n162 104.615
R754 VDD1.n164 VDD1.n163 104.615
R755 VDD1.n163 VDD1.n100 104.615
R756 VDD1.n172 VDD1.n100 104.615
R757 VDD1.n173 VDD1.n172 104.615
R758 VDD1.n173 VDD1.n96 104.615
R759 VDD1.n180 VDD1.n96 104.615
R760 VDD1.n181 VDD1.n180 104.615
R761 VDD1.n187 VDD1.n186 64.4383
R762 VDD1.n189 VDD1.n188 63.6337
R763 VDD1 VDD1.n92 54.4112
R764 VDD1.n187 VDD1.n185 54.2976
R765 VDD1.n31 VDD1.t5 52.3082
R766 VDD1.n123 VDD1.t0 52.3082
R767 VDD1.n189 VDD1.n187 51.8091
R768 VDD1.n32 VDD1.n30 15.6677
R769 VDD1.n124 VDD1.n122 15.6677
R770 VDD1.n78 VDD1.n77 13.1884
R771 VDD1.n171 VDD1.n170 13.1884
R772 VDD1.n81 VDD1.n6 12.8005
R773 VDD1.n76 VDD1.n8 12.8005
R774 VDD1.n33 VDD1.n29 12.8005
R775 VDD1.n125 VDD1.n121 12.8005
R776 VDD1.n169 VDD1.n101 12.8005
R777 VDD1.n174 VDD1.n99 12.8005
R778 VDD1.n82 VDD1.n4 12.0247
R779 VDD1.n73 VDD1.n72 12.0247
R780 VDD1.n37 VDD1.n36 12.0247
R781 VDD1.n129 VDD1.n128 12.0247
R782 VDD1.n166 VDD1.n165 12.0247
R783 VDD1.n175 VDD1.n97 12.0247
R784 VDD1.n86 VDD1.n85 11.249
R785 VDD1.n69 VDD1.n10 11.249
R786 VDD1.n40 VDD1.n27 11.249
R787 VDD1.n132 VDD1.n119 11.249
R788 VDD1.n161 VDD1.n103 11.249
R789 VDD1.n179 VDD1.n178 11.249
R790 VDD1.n89 VDD1.n2 10.4732
R791 VDD1.n68 VDD1.n13 10.4732
R792 VDD1.n41 VDD1.n25 10.4732
R793 VDD1.n133 VDD1.n117 10.4732
R794 VDD1.n160 VDD1.n105 10.4732
R795 VDD1.n182 VDD1.n95 10.4732
R796 VDD1.n90 VDD1.n0 9.69747
R797 VDD1.n65 VDD1.n64 9.69747
R798 VDD1.n45 VDD1.n44 9.69747
R799 VDD1.n137 VDD1.n136 9.69747
R800 VDD1.n157 VDD1.n156 9.69747
R801 VDD1.n183 VDD1.n93 9.69747
R802 VDD1.n92 VDD1.n91 9.45567
R803 VDD1.n185 VDD1.n184 9.45567
R804 VDD1.n58 VDD1.n57 9.3005
R805 VDD1.n60 VDD1.n59 9.3005
R806 VDD1.n15 VDD1.n14 9.3005
R807 VDD1.n66 VDD1.n65 9.3005
R808 VDD1.n68 VDD1.n67 9.3005
R809 VDD1.n10 VDD1.n9 9.3005
R810 VDD1.n74 VDD1.n73 9.3005
R811 VDD1.n76 VDD1.n75 9.3005
R812 VDD1.n91 VDD1.n90 9.3005
R813 VDD1.n2 VDD1.n1 9.3005
R814 VDD1.n85 VDD1.n84 9.3005
R815 VDD1.n83 VDD1.n82 9.3005
R816 VDD1.n6 VDD1.n5 9.3005
R817 VDD1.n19 VDD1.n18 9.3005
R818 VDD1.n52 VDD1.n51 9.3005
R819 VDD1.n50 VDD1.n49 9.3005
R820 VDD1.n23 VDD1.n22 9.3005
R821 VDD1.n44 VDD1.n43 9.3005
R822 VDD1.n42 VDD1.n41 9.3005
R823 VDD1.n27 VDD1.n26 9.3005
R824 VDD1.n36 VDD1.n35 9.3005
R825 VDD1.n34 VDD1.n33 9.3005
R826 VDD1.n184 VDD1.n183 9.3005
R827 VDD1.n95 VDD1.n94 9.3005
R828 VDD1.n178 VDD1.n177 9.3005
R829 VDD1.n176 VDD1.n175 9.3005
R830 VDD1.n99 VDD1.n98 9.3005
R831 VDD1.n144 VDD1.n143 9.3005
R832 VDD1.n142 VDD1.n141 9.3005
R833 VDD1.n115 VDD1.n114 9.3005
R834 VDD1.n136 VDD1.n135 9.3005
R835 VDD1.n134 VDD1.n133 9.3005
R836 VDD1.n119 VDD1.n118 9.3005
R837 VDD1.n128 VDD1.n127 9.3005
R838 VDD1.n126 VDD1.n125 9.3005
R839 VDD1.n111 VDD1.n110 9.3005
R840 VDD1.n150 VDD1.n149 9.3005
R841 VDD1.n152 VDD1.n151 9.3005
R842 VDD1.n107 VDD1.n106 9.3005
R843 VDD1.n158 VDD1.n157 9.3005
R844 VDD1.n160 VDD1.n159 9.3005
R845 VDD1.n103 VDD1.n102 9.3005
R846 VDD1.n167 VDD1.n166 9.3005
R847 VDD1.n169 VDD1.n168 9.3005
R848 VDD1.n61 VDD1.n15 8.92171
R849 VDD1.n48 VDD1.n23 8.92171
R850 VDD1.n140 VDD1.n115 8.92171
R851 VDD1.n153 VDD1.n107 8.92171
R852 VDD1.n60 VDD1.n17 8.14595
R853 VDD1.n49 VDD1.n21 8.14595
R854 VDD1.n141 VDD1.n113 8.14595
R855 VDD1.n152 VDD1.n109 8.14595
R856 VDD1.n57 VDD1.n56 7.3702
R857 VDD1.n53 VDD1.n52 7.3702
R858 VDD1.n145 VDD1.n144 7.3702
R859 VDD1.n149 VDD1.n148 7.3702
R860 VDD1.n56 VDD1.n19 6.59444
R861 VDD1.n53 VDD1.n19 6.59444
R862 VDD1.n145 VDD1.n111 6.59444
R863 VDD1.n148 VDD1.n111 6.59444
R864 VDD1.n57 VDD1.n17 5.81868
R865 VDD1.n52 VDD1.n21 5.81868
R866 VDD1.n144 VDD1.n113 5.81868
R867 VDD1.n149 VDD1.n109 5.81868
R868 VDD1.n61 VDD1.n60 5.04292
R869 VDD1.n49 VDD1.n48 5.04292
R870 VDD1.n141 VDD1.n140 5.04292
R871 VDD1.n153 VDD1.n152 5.04292
R872 VDD1.n34 VDD1.n30 4.38563
R873 VDD1.n126 VDD1.n122 4.38563
R874 VDD1.n92 VDD1.n0 4.26717
R875 VDD1.n64 VDD1.n15 4.26717
R876 VDD1.n45 VDD1.n23 4.26717
R877 VDD1.n137 VDD1.n115 4.26717
R878 VDD1.n156 VDD1.n107 4.26717
R879 VDD1.n185 VDD1.n93 4.26717
R880 VDD1.n90 VDD1.n89 3.49141
R881 VDD1.n65 VDD1.n13 3.49141
R882 VDD1.n44 VDD1.n25 3.49141
R883 VDD1.n136 VDD1.n117 3.49141
R884 VDD1.n157 VDD1.n105 3.49141
R885 VDD1.n183 VDD1.n182 3.49141
R886 VDD1.n86 VDD1.n2 2.71565
R887 VDD1.n69 VDD1.n68 2.71565
R888 VDD1.n41 VDD1.n40 2.71565
R889 VDD1.n133 VDD1.n132 2.71565
R890 VDD1.n161 VDD1.n160 2.71565
R891 VDD1.n179 VDD1.n95 2.71565
R892 VDD1.n85 VDD1.n4 1.93989
R893 VDD1.n72 VDD1.n10 1.93989
R894 VDD1.n37 VDD1.n27 1.93989
R895 VDD1.n129 VDD1.n119 1.93989
R896 VDD1.n165 VDD1.n103 1.93989
R897 VDD1.n178 VDD1.n97 1.93989
R898 VDD1.n188 VDD1.t2 1.16864
R899 VDD1.n188 VDD1.t1 1.16864
R900 VDD1.n186 VDD1.t4 1.16864
R901 VDD1.n186 VDD1.t3 1.16864
R902 VDD1.n82 VDD1.n81 1.16414
R903 VDD1.n73 VDD1.n8 1.16414
R904 VDD1.n36 VDD1.n29 1.16414
R905 VDD1.n128 VDD1.n121 1.16414
R906 VDD1.n166 VDD1.n101 1.16414
R907 VDD1.n175 VDD1.n174 1.16414
R908 VDD1 VDD1.n189 0.802224
R909 VDD1.n78 VDD1.n6 0.388379
R910 VDD1.n77 VDD1.n76 0.388379
R911 VDD1.n33 VDD1.n32 0.388379
R912 VDD1.n125 VDD1.n124 0.388379
R913 VDD1.n170 VDD1.n169 0.388379
R914 VDD1.n171 VDD1.n99 0.388379
R915 VDD1.n91 VDD1.n1 0.155672
R916 VDD1.n84 VDD1.n1 0.155672
R917 VDD1.n84 VDD1.n83 0.155672
R918 VDD1.n83 VDD1.n5 0.155672
R919 VDD1.n75 VDD1.n5 0.155672
R920 VDD1.n75 VDD1.n74 0.155672
R921 VDD1.n74 VDD1.n9 0.155672
R922 VDD1.n67 VDD1.n9 0.155672
R923 VDD1.n67 VDD1.n66 0.155672
R924 VDD1.n66 VDD1.n14 0.155672
R925 VDD1.n59 VDD1.n14 0.155672
R926 VDD1.n59 VDD1.n58 0.155672
R927 VDD1.n58 VDD1.n18 0.155672
R928 VDD1.n51 VDD1.n18 0.155672
R929 VDD1.n51 VDD1.n50 0.155672
R930 VDD1.n50 VDD1.n22 0.155672
R931 VDD1.n43 VDD1.n22 0.155672
R932 VDD1.n43 VDD1.n42 0.155672
R933 VDD1.n42 VDD1.n26 0.155672
R934 VDD1.n35 VDD1.n26 0.155672
R935 VDD1.n35 VDD1.n34 0.155672
R936 VDD1.n127 VDD1.n126 0.155672
R937 VDD1.n127 VDD1.n118 0.155672
R938 VDD1.n134 VDD1.n118 0.155672
R939 VDD1.n135 VDD1.n134 0.155672
R940 VDD1.n135 VDD1.n114 0.155672
R941 VDD1.n142 VDD1.n114 0.155672
R942 VDD1.n143 VDD1.n142 0.155672
R943 VDD1.n143 VDD1.n110 0.155672
R944 VDD1.n150 VDD1.n110 0.155672
R945 VDD1.n151 VDD1.n150 0.155672
R946 VDD1.n151 VDD1.n106 0.155672
R947 VDD1.n158 VDD1.n106 0.155672
R948 VDD1.n159 VDD1.n158 0.155672
R949 VDD1.n159 VDD1.n102 0.155672
R950 VDD1.n167 VDD1.n102 0.155672
R951 VDD1.n168 VDD1.n167 0.155672
R952 VDD1.n168 VDD1.n98 0.155672
R953 VDD1.n176 VDD1.n98 0.155672
R954 VDD1.n177 VDD1.n176 0.155672
R955 VDD1.n177 VDD1.n94 0.155672
R956 VDD1.n184 VDD1.n94 0.155672
R957 B.n1060 B.n1059 585
R958 B.n406 B.n162 585
R959 B.n405 B.n404 585
R960 B.n403 B.n402 585
R961 B.n401 B.n400 585
R962 B.n399 B.n398 585
R963 B.n397 B.n396 585
R964 B.n395 B.n394 585
R965 B.n393 B.n392 585
R966 B.n391 B.n390 585
R967 B.n389 B.n388 585
R968 B.n387 B.n386 585
R969 B.n385 B.n384 585
R970 B.n383 B.n382 585
R971 B.n381 B.n380 585
R972 B.n379 B.n378 585
R973 B.n377 B.n376 585
R974 B.n375 B.n374 585
R975 B.n373 B.n372 585
R976 B.n371 B.n370 585
R977 B.n369 B.n368 585
R978 B.n367 B.n366 585
R979 B.n365 B.n364 585
R980 B.n363 B.n362 585
R981 B.n361 B.n360 585
R982 B.n359 B.n358 585
R983 B.n357 B.n356 585
R984 B.n355 B.n354 585
R985 B.n353 B.n352 585
R986 B.n351 B.n350 585
R987 B.n349 B.n348 585
R988 B.n347 B.n346 585
R989 B.n345 B.n344 585
R990 B.n343 B.n342 585
R991 B.n341 B.n340 585
R992 B.n339 B.n338 585
R993 B.n337 B.n336 585
R994 B.n335 B.n334 585
R995 B.n333 B.n332 585
R996 B.n331 B.n330 585
R997 B.n329 B.n328 585
R998 B.n327 B.n326 585
R999 B.n325 B.n324 585
R1000 B.n323 B.n322 585
R1001 B.n321 B.n320 585
R1002 B.n319 B.n318 585
R1003 B.n317 B.n316 585
R1004 B.n315 B.n314 585
R1005 B.n313 B.n312 585
R1006 B.n311 B.n310 585
R1007 B.n309 B.n308 585
R1008 B.n307 B.n306 585
R1009 B.n305 B.n304 585
R1010 B.n303 B.n302 585
R1011 B.n301 B.n300 585
R1012 B.n299 B.n298 585
R1013 B.n297 B.n296 585
R1014 B.n295 B.n294 585
R1015 B.n293 B.n292 585
R1016 B.n291 B.n290 585
R1017 B.n289 B.n288 585
R1018 B.n287 B.n286 585
R1019 B.n285 B.n284 585
R1020 B.n283 B.n282 585
R1021 B.n281 B.n280 585
R1022 B.n279 B.n278 585
R1023 B.n277 B.n276 585
R1024 B.n275 B.n274 585
R1025 B.n273 B.n272 585
R1026 B.n271 B.n270 585
R1027 B.n269 B.n268 585
R1028 B.n267 B.n266 585
R1029 B.n265 B.n264 585
R1030 B.n263 B.n262 585
R1031 B.n261 B.n260 585
R1032 B.n259 B.n258 585
R1033 B.n257 B.n256 585
R1034 B.n255 B.n254 585
R1035 B.n253 B.n252 585
R1036 B.n251 B.n250 585
R1037 B.n249 B.n248 585
R1038 B.n247 B.n246 585
R1039 B.n245 B.n244 585
R1040 B.n243 B.n242 585
R1041 B.n241 B.n240 585
R1042 B.n239 B.n238 585
R1043 B.n237 B.n236 585
R1044 B.n235 B.n234 585
R1045 B.n233 B.n232 585
R1046 B.n231 B.n230 585
R1047 B.n229 B.n228 585
R1048 B.n227 B.n226 585
R1049 B.n225 B.n224 585
R1050 B.n223 B.n222 585
R1051 B.n221 B.n220 585
R1052 B.n219 B.n218 585
R1053 B.n217 B.n216 585
R1054 B.n215 B.n214 585
R1055 B.n213 B.n212 585
R1056 B.n211 B.n210 585
R1057 B.n209 B.n208 585
R1058 B.n207 B.n206 585
R1059 B.n205 B.n204 585
R1060 B.n203 B.n202 585
R1061 B.n201 B.n200 585
R1062 B.n199 B.n198 585
R1063 B.n197 B.n196 585
R1064 B.n195 B.n194 585
R1065 B.n193 B.n192 585
R1066 B.n191 B.n190 585
R1067 B.n189 B.n188 585
R1068 B.n187 B.n186 585
R1069 B.n185 B.n184 585
R1070 B.n183 B.n182 585
R1071 B.n181 B.n180 585
R1072 B.n179 B.n178 585
R1073 B.n177 B.n176 585
R1074 B.n175 B.n174 585
R1075 B.n173 B.n172 585
R1076 B.n171 B.n170 585
R1077 B.n102 B.n101 585
R1078 B.n1065 B.n1064 585
R1079 B.n1058 B.n163 585
R1080 B.n163 B.n99 585
R1081 B.n1057 B.n98 585
R1082 B.n1069 B.n98 585
R1083 B.n1056 B.n97 585
R1084 B.n1070 B.n97 585
R1085 B.n1055 B.n96 585
R1086 B.n1071 B.n96 585
R1087 B.n1054 B.n1053 585
R1088 B.n1053 B.n92 585
R1089 B.n1052 B.n91 585
R1090 B.n1077 B.n91 585
R1091 B.n1051 B.n90 585
R1092 B.n1078 B.n90 585
R1093 B.n1050 B.n89 585
R1094 B.n1079 B.n89 585
R1095 B.n1049 B.n1048 585
R1096 B.n1048 B.n85 585
R1097 B.n1047 B.n84 585
R1098 B.n1085 B.n84 585
R1099 B.n1046 B.n83 585
R1100 B.n1086 B.n83 585
R1101 B.n1045 B.n82 585
R1102 B.n1087 B.n82 585
R1103 B.n1044 B.n1043 585
R1104 B.n1043 B.n78 585
R1105 B.n1042 B.n77 585
R1106 B.n1093 B.n77 585
R1107 B.n1041 B.n76 585
R1108 B.n1094 B.n76 585
R1109 B.n1040 B.n75 585
R1110 B.n1095 B.n75 585
R1111 B.n1039 B.n1038 585
R1112 B.n1038 B.n71 585
R1113 B.n1037 B.n70 585
R1114 B.n1101 B.n70 585
R1115 B.n1036 B.n69 585
R1116 B.n1102 B.n69 585
R1117 B.n1035 B.n68 585
R1118 B.n1103 B.n68 585
R1119 B.n1034 B.n1033 585
R1120 B.n1033 B.n64 585
R1121 B.n1032 B.n63 585
R1122 B.n1109 B.n63 585
R1123 B.n1031 B.n62 585
R1124 B.n1110 B.n62 585
R1125 B.n1030 B.n61 585
R1126 B.n1111 B.n61 585
R1127 B.n1029 B.n1028 585
R1128 B.n1028 B.n60 585
R1129 B.n1027 B.n56 585
R1130 B.n1117 B.n56 585
R1131 B.n1026 B.n55 585
R1132 B.n1118 B.n55 585
R1133 B.n1025 B.n54 585
R1134 B.n1119 B.n54 585
R1135 B.n1024 B.n1023 585
R1136 B.n1023 B.n50 585
R1137 B.n1022 B.n49 585
R1138 B.n1125 B.n49 585
R1139 B.n1021 B.n48 585
R1140 B.n1126 B.n48 585
R1141 B.n1020 B.n47 585
R1142 B.n1127 B.n47 585
R1143 B.n1019 B.n1018 585
R1144 B.n1018 B.n43 585
R1145 B.n1017 B.n42 585
R1146 B.n1133 B.n42 585
R1147 B.n1016 B.n41 585
R1148 B.n1134 B.n41 585
R1149 B.n1015 B.n40 585
R1150 B.n1135 B.n40 585
R1151 B.n1014 B.n1013 585
R1152 B.n1013 B.n36 585
R1153 B.n1012 B.n35 585
R1154 B.n1141 B.n35 585
R1155 B.n1011 B.n34 585
R1156 B.n1142 B.n34 585
R1157 B.n1010 B.n33 585
R1158 B.n1143 B.n33 585
R1159 B.n1009 B.n1008 585
R1160 B.n1008 B.n29 585
R1161 B.n1007 B.n28 585
R1162 B.n1149 B.n28 585
R1163 B.n1006 B.n27 585
R1164 B.n1150 B.n27 585
R1165 B.n1005 B.n26 585
R1166 B.n1151 B.n26 585
R1167 B.n1004 B.n1003 585
R1168 B.n1003 B.n22 585
R1169 B.n1002 B.n21 585
R1170 B.n1157 B.n21 585
R1171 B.n1001 B.n20 585
R1172 B.n1158 B.n20 585
R1173 B.n1000 B.n19 585
R1174 B.n1159 B.n19 585
R1175 B.n999 B.n998 585
R1176 B.n998 B.n15 585
R1177 B.n997 B.n14 585
R1178 B.n1165 B.n14 585
R1179 B.n996 B.n13 585
R1180 B.n1166 B.n13 585
R1181 B.n995 B.n12 585
R1182 B.n1167 B.n12 585
R1183 B.n994 B.n993 585
R1184 B.n993 B.n8 585
R1185 B.n992 B.n7 585
R1186 B.n1173 B.n7 585
R1187 B.n991 B.n6 585
R1188 B.n1174 B.n6 585
R1189 B.n990 B.n5 585
R1190 B.n1175 B.n5 585
R1191 B.n989 B.n988 585
R1192 B.n988 B.n4 585
R1193 B.n987 B.n407 585
R1194 B.n987 B.n986 585
R1195 B.n977 B.n408 585
R1196 B.n409 B.n408 585
R1197 B.n979 B.n978 585
R1198 B.n980 B.n979 585
R1199 B.n976 B.n414 585
R1200 B.n414 B.n413 585
R1201 B.n975 B.n974 585
R1202 B.n974 B.n973 585
R1203 B.n416 B.n415 585
R1204 B.n417 B.n416 585
R1205 B.n966 B.n965 585
R1206 B.n967 B.n966 585
R1207 B.n964 B.n422 585
R1208 B.n422 B.n421 585
R1209 B.n963 B.n962 585
R1210 B.n962 B.n961 585
R1211 B.n424 B.n423 585
R1212 B.n425 B.n424 585
R1213 B.n954 B.n953 585
R1214 B.n955 B.n954 585
R1215 B.n952 B.n430 585
R1216 B.n430 B.n429 585
R1217 B.n951 B.n950 585
R1218 B.n950 B.n949 585
R1219 B.n432 B.n431 585
R1220 B.n433 B.n432 585
R1221 B.n942 B.n941 585
R1222 B.n943 B.n942 585
R1223 B.n940 B.n438 585
R1224 B.n438 B.n437 585
R1225 B.n939 B.n938 585
R1226 B.n938 B.n937 585
R1227 B.n440 B.n439 585
R1228 B.n441 B.n440 585
R1229 B.n930 B.n929 585
R1230 B.n931 B.n930 585
R1231 B.n928 B.n446 585
R1232 B.n446 B.n445 585
R1233 B.n927 B.n926 585
R1234 B.n926 B.n925 585
R1235 B.n448 B.n447 585
R1236 B.n449 B.n448 585
R1237 B.n918 B.n917 585
R1238 B.n919 B.n918 585
R1239 B.n916 B.n454 585
R1240 B.n454 B.n453 585
R1241 B.n915 B.n914 585
R1242 B.n914 B.n913 585
R1243 B.n456 B.n455 585
R1244 B.n457 B.n456 585
R1245 B.n906 B.n905 585
R1246 B.n907 B.n906 585
R1247 B.n904 B.n462 585
R1248 B.n462 B.n461 585
R1249 B.n903 B.n902 585
R1250 B.n902 B.n901 585
R1251 B.n464 B.n463 585
R1252 B.n894 B.n464 585
R1253 B.n893 B.n892 585
R1254 B.n895 B.n893 585
R1255 B.n891 B.n469 585
R1256 B.n469 B.n468 585
R1257 B.n890 B.n889 585
R1258 B.n889 B.n888 585
R1259 B.n471 B.n470 585
R1260 B.n472 B.n471 585
R1261 B.n881 B.n880 585
R1262 B.n882 B.n881 585
R1263 B.n879 B.n477 585
R1264 B.n477 B.n476 585
R1265 B.n878 B.n877 585
R1266 B.n877 B.n876 585
R1267 B.n479 B.n478 585
R1268 B.n480 B.n479 585
R1269 B.n869 B.n868 585
R1270 B.n870 B.n869 585
R1271 B.n867 B.n485 585
R1272 B.n485 B.n484 585
R1273 B.n866 B.n865 585
R1274 B.n865 B.n864 585
R1275 B.n487 B.n486 585
R1276 B.n488 B.n487 585
R1277 B.n857 B.n856 585
R1278 B.n858 B.n857 585
R1279 B.n855 B.n493 585
R1280 B.n493 B.n492 585
R1281 B.n854 B.n853 585
R1282 B.n853 B.n852 585
R1283 B.n495 B.n494 585
R1284 B.n496 B.n495 585
R1285 B.n845 B.n844 585
R1286 B.n846 B.n845 585
R1287 B.n843 B.n501 585
R1288 B.n501 B.n500 585
R1289 B.n842 B.n841 585
R1290 B.n841 B.n840 585
R1291 B.n503 B.n502 585
R1292 B.n504 B.n503 585
R1293 B.n833 B.n832 585
R1294 B.n834 B.n833 585
R1295 B.n831 B.n509 585
R1296 B.n509 B.n508 585
R1297 B.n830 B.n829 585
R1298 B.n829 B.n828 585
R1299 B.n511 B.n510 585
R1300 B.n512 B.n511 585
R1301 B.n824 B.n823 585
R1302 B.n515 B.n514 585
R1303 B.n820 B.n819 585
R1304 B.n821 B.n820 585
R1305 B.n818 B.n576 585
R1306 B.n817 B.n816 585
R1307 B.n815 B.n814 585
R1308 B.n813 B.n812 585
R1309 B.n811 B.n810 585
R1310 B.n809 B.n808 585
R1311 B.n807 B.n806 585
R1312 B.n805 B.n804 585
R1313 B.n803 B.n802 585
R1314 B.n801 B.n800 585
R1315 B.n799 B.n798 585
R1316 B.n797 B.n796 585
R1317 B.n795 B.n794 585
R1318 B.n793 B.n792 585
R1319 B.n791 B.n790 585
R1320 B.n789 B.n788 585
R1321 B.n787 B.n786 585
R1322 B.n785 B.n784 585
R1323 B.n783 B.n782 585
R1324 B.n781 B.n780 585
R1325 B.n779 B.n778 585
R1326 B.n777 B.n776 585
R1327 B.n775 B.n774 585
R1328 B.n773 B.n772 585
R1329 B.n771 B.n770 585
R1330 B.n769 B.n768 585
R1331 B.n767 B.n766 585
R1332 B.n765 B.n764 585
R1333 B.n763 B.n762 585
R1334 B.n761 B.n760 585
R1335 B.n759 B.n758 585
R1336 B.n757 B.n756 585
R1337 B.n755 B.n754 585
R1338 B.n753 B.n752 585
R1339 B.n751 B.n750 585
R1340 B.n749 B.n748 585
R1341 B.n747 B.n746 585
R1342 B.n745 B.n744 585
R1343 B.n743 B.n742 585
R1344 B.n741 B.n740 585
R1345 B.n739 B.n738 585
R1346 B.n737 B.n736 585
R1347 B.n735 B.n734 585
R1348 B.n733 B.n732 585
R1349 B.n731 B.n730 585
R1350 B.n729 B.n728 585
R1351 B.n727 B.n726 585
R1352 B.n725 B.n724 585
R1353 B.n723 B.n722 585
R1354 B.n721 B.n720 585
R1355 B.n719 B.n718 585
R1356 B.n717 B.n716 585
R1357 B.n715 B.n714 585
R1358 B.n712 B.n711 585
R1359 B.n710 B.n709 585
R1360 B.n708 B.n707 585
R1361 B.n706 B.n705 585
R1362 B.n704 B.n703 585
R1363 B.n702 B.n701 585
R1364 B.n700 B.n699 585
R1365 B.n698 B.n697 585
R1366 B.n696 B.n695 585
R1367 B.n694 B.n693 585
R1368 B.n691 B.n690 585
R1369 B.n689 B.n688 585
R1370 B.n687 B.n686 585
R1371 B.n685 B.n684 585
R1372 B.n683 B.n682 585
R1373 B.n681 B.n680 585
R1374 B.n679 B.n678 585
R1375 B.n677 B.n676 585
R1376 B.n675 B.n674 585
R1377 B.n673 B.n672 585
R1378 B.n671 B.n670 585
R1379 B.n669 B.n668 585
R1380 B.n667 B.n666 585
R1381 B.n665 B.n664 585
R1382 B.n663 B.n662 585
R1383 B.n661 B.n660 585
R1384 B.n659 B.n658 585
R1385 B.n657 B.n656 585
R1386 B.n655 B.n654 585
R1387 B.n653 B.n652 585
R1388 B.n651 B.n650 585
R1389 B.n649 B.n648 585
R1390 B.n647 B.n646 585
R1391 B.n645 B.n644 585
R1392 B.n643 B.n642 585
R1393 B.n641 B.n640 585
R1394 B.n639 B.n638 585
R1395 B.n637 B.n636 585
R1396 B.n635 B.n634 585
R1397 B.n633 B.n632 585
R1398 B.n631 B.n630 585
R1399 B.n629 B.n628 585
R1400 B.n627 B.n626 585
R1401 B.n625 B.n624 585
R1402 B.n623 B.n622 585
R1403 B.n621 B.n620 585
R1404 B.n619 B.n618 585
R1405 B.n617 B.n616 585
R1406 B.n615 B.n614 585
R1407 B.n613 B.n612 585
R1408 B.n611 B.n610 585
R1409 B.n609 B.n608 585
R1410 B.n607 B.n606 585
R1411 B.n605 B.n604 585
R1412 B.n603 B.n602 585
R1413 B.n601 B.n600 585
R1414 B.n599 B.n598 585
R1415 B.n597 B.n596 585
R1416 B.n595 B.n594 585
R1417 B.n593 B.n592 585
R1418 B.n591 B.n590 585
R1419 B.n589 B.n588 585
R1420 B.n587 B.n586 585
R1421 B.n585 B.n584 585
R1422 B.n583 B.n582 585
R1423 B.n581 B.n575 585
R1424 B.n821 B.n575 585
R1425 B.n825 B.n513 585
R1426 B.n513 B.n512 585
R1427 B.n827 B.n826 585
R1428 B.n828 B.n827 585
R1429 B.n507 B.n506 585
R1430 B.n508 B.n507 585
R1431 B.n836 B.n835 585
R1432 B.n835 B.n834 585
R1433 B.n837 B.n505 585
R1434 B.n505 B.n504 585
R1435 B.n839 B.n838 585
R1436 B.n840 B.n839 585
R1437 B.n499 B.n498 585
R1438 B.n500 B.n499 585
R1439 B.n848 B.n847 585
R1440 B.n847 B.n846 585
R1441 B.n849 B.n497 585
R1442 B.n497 B.n496 585
R1443 B.n851 B.n850 585
R1444 B.n852 B.n851 585
R1445 B.n491 B.n490 585
R1446 B.n492 B.n491 585
R1447 B.n860 B.n859 585
R1448 B.n859 B.n858 585
R1449 B.n861 B.n489 585
R1450 B.n489 B.n488 585
R1451 B.n863 B.n862 585
R1452 B.n864 B.n863 585
R1453 B.n483 B.n482 585
R1454 B.n484 B.n483 585
R1455 B.n872 B.n871 585
R1456 B.n871 B.n870 585
R1457 B.n873 B.n481 585
R1458 B.n481 B.n480 585
R1459 B.n875 B.n874 585
R1460 B.n876 B.n875 585
R1461 B.n475 B.n474 585
R1462 B.n476 B.n475 585
R1463 B.n884 B.n883 585
R1464 B.n883 B.n882 585
R1465 B.n885 B.n473 585
R1466 B.n473 B.n472 585
R1467 B.n887 B.n886 585
R1468 B.n888 B.n887 585
R1469 B.n467 B.n466 585
R1470 B.n468 B.n467 585
R1471 B.n897 B.n896 585
R1472 B.n896 B.n895 585
R1473 B.n898 B.n465 585
R1474 B.n894 B.n465 585
R1475 B.n900 B.n899 585
R1476 B.n901 B.n900 585
R1477 B.n460 B.n459 585
R1478 B.n461 B.n460 585
R1479 B.n909 B.n908 585
R1480 B.n908 B.n907 585
R1481 B.n910 B.n458 585
R1482 B.n458 B.n457 585
R1483 B.n912 B.n911 585
R1484 B.n913 B.n912 585
R1485 B.n452 B.n451 585
R1486 B.n453 B.n452 585
R1487 B.n921 B.n920 585
R1488 B.n920 B.n919 585
R1489 B.n922 B.n450 585
R1490 B.n450 B.n449 585
R1491 B.n924 B.n923 585
R1492 B.n925 B.n924 585
R1493 B.n444 B.n443 585
R1494 B.n445 B.n444 585
R1495 B.n933 B.n932 585
R1496 B.n932 B.n931 585
R1497 B.n934 B.n442 585
R1498 B.n442 B.n441 585
R1499 B.n936 B.n935 585
R1500 B.n937 B.n936 585
R1501 B.n436 B.n435 585
R1502 B.n437 B.n436 585
R1503 B.n945 B.n944 585
R1504 B.n944 B.n943 585
R1505 B.n946 B.n434 585
R1506 B.n434 B.n433 585
R1507 B.n948 B.n947 585
R1508 B.n949 B.n948 585
R1509 B.n428 B.n427 585
R1510 B.n429 B.n428 585
R1511 B.n957 B.n956 585
R1512 B.n956 B.n955 585
R1513 B.n958 B.n426 585
R1514 B.n426 B.n425 585
R1515 B.n960 B.n959 585
R1516 B.n961 B.n960 585
R1517 B.n420 B.n419 585
R1518 B.n421 B.n420 585
R1519 B.n969 B.n968 585
R1520 B.n968 B.n967 585
R1521 B.n970 B.n418 585
R1522 B.n418 B.n417 585
R1523 B.n972 B.n971 585
R1524 B.n973 B.n972 585
R1525 B.n412 B.n411 585
R1526 B.n413 B.n412 585
R1527 B.n982 B.n981 585
R1528 B.n981 B.n980 585
R1529 B.n983 B.n410 585
R1530 B.n410 B.n409 585
R1531 B.n985 B.n984 585
R1532 B.n986 B.n985 585
R1533 B.n2 B.n0 585
R1534 B.n4 B.n2 585
R1535 B.n3 B.n1 585
R1536 B.n1174 B.n3 585
R1537 B.n1172 B.n1171 585
R1538 B.n1173 B.n1172 585
R1539 B.n1170 B.n9 585
R1540 B.n9 B.n8 585
R1541 B.n1169 B.n1168 585
R1542 B.n1168 B.n1167 585
R1543 B.n11 B.n10 585
R1544 B.n1166 B.n11 585
R1545 B.n1164 B.n1163 585
R1546 B.n1165 B.n1164 585
R1547 B.n1162 B.n16 585
R1548 B.n16 B.n15 585
R1549 B.n1161 B.n1160 585
R1550 B.n1160 B.n1159 585
R1551 B.n18 B.n17 585
R1552 B.n1158 B.n18 585
R1553 B.n1156 B.n1155 585
R1554 B.n1157 B.n1156 585
R1555 B.n1154 B.n23 585
R1556 B.n23 B.n22 585
R1557 B.n1153 B.n1152 585
R1558 B.n1152 B.n1151 585
R1559 B.n25 B.n24 585
R1560 B.n1150 B.n25 585
R1561 B.n1148 B.n1147 585
R1562 B.n1149 B.n1148 585
R1563 B.n1146 B.n30 585
R1564 B.n30 B.n29 585
R1565 B.n1145 B.n1144 585
R1566 B.n1144 B.n1143 585
R1567 B.n32 B.n31 585
R1568 B.n1142 B.n32 585
R1569 B.n1140 B.n1139 585
R1570 B.n1141 B.n1140 585
R1571 B.n1138 B.n37 585
R1572 B.n37 B.n36 585
R1573 B.n1137 B.n1136 585
R1574 B.n1136 B.n1135 585
R1575 B.n39 B.n38 585
R1576 B.n1134 B.n39 585
R1577 B.n1132 B.n1131 585
R1578 B.n1133 B.n1132 585
R1579 B.n1130 B.n44 585
R1580 B.n44 B.n43 585
R1581 B.n1129 B.n1128 585
R1582 B.n1128 B.n1127 585
R1583 B.n46 B.n45 585
R1584 B.n1126 B.n46 585
R1585 B.n1124 B.n1123 585
R1586 B.n1125 B.n1124 585
R1587 B.n1122 B.n51 585
R1588 B.n51 B.n50 585
R1589 B.n1121 B.n1120 585
R1590 B.n1120 B.n1119 585
R1591 B.n53 B.n52 585
R1592 B.n1118 B.n53 585
R1593 B.n1116 B.n1115 585
R1594 B.n1117 B.n1116 585
R1595 B.n1114 B.n57 585
R1596 B.n60 B.n57 585
R1597 B.n1113 B.n1112 585
R1598 B.n1112 B.n1111 585
R1599 B.n59 B.n58 585
R1600 B.n1110 B.n59 585
R1601 B.n1108 B.n1107 585
R1602 B.n1109 B.n1108 585
R1603 B.n1106 B.n65 585
R1604 B.n65 B.n64 585
R1605 B.n1105 B.n1104 585
R1606 B.n1104 B.n1103 585
R1607 B.n67 B.n66 585
R1608 B.n1102 B.n67 585
R1609 B.n1100 B.n1099 585
R1610 B.n1101 B.n1100 585
R1611 B.n1098 B.n72 585
R1612 B.n72 B.n71 585
R1613 B.n1097 B.n1096 585
R1614 B.n1096 B.n1095 585
R1615 B.n74 B.n73 585
R1616 B.n1094 B.n74 585
R1617 B.n1092 B.n1091 585
R1618 B.n1093 B.n1092 585
R1619 B.n1090 B.n79 585
R1620 B.n79 B.n78 585
R1621 B.n1089 B.n1088 585
R1622 B.n1088 B.n1087 585
R1623 B.n81 B.n80 585
R1624 B.n1086 B.n81 585
R1625 B.n1084 B.n1083 585
R1626 B.n1085 B.n1084 585
R1627 B.n1082 B.n86 585
R1628 B.n86 B.n85 585
R1629 B.n1081 B.n1080 585
R1630 B.n1080 B.n1079 585
R1631 B.n88 B.n87 585
R1632 B.n1078 B.n88 585
R1633 B.n1076 B.n1075 585
R1634 B.n1077 B.n1076 585
R1635 B.n1074 B.n93 585
R1636 B.n93 B.n92 585
R1637 B.n1073 B.n1072 585
R1638 B.n1072 B.n1071 585
R1639 B.n95 B.n94 585
R1640 B.n1070 B.n95 585
R1641 B.n1068 B.n1067 585
R1642 B.n1069 B.n1068 585
R1643 B.n1066 B.n100 585
R1644 B.n100 B.n99 585
R1645 B.n1177 B.n1176 585
R1646 B.n1176 B.n1175 585
R1647 B.n823 B.n513 502.111
R1648 B.n1064 B.n100 502.111
R1649 B.n575 B.n511 502.111
R1650 B.n1060 B.n163 502.111
R1651 B.n579 B.t16 445.062
R1652 B.n577 B.t9 445.062
R1653 B.n167 B.t12 445.062
R1654 B.n164 B.t18 445.062
R1655 B.n580 B.t15 367.68
R1656 B.n165 B.t19 367.68
R1657 B.n578 B.t8 367.68
R1658 B.n168 B.t13 367.68
R1659 B.n579 B.t14 320.842
R1660 B.n577 B.t6 320.842
R1661 B.n167 B.t10 320.842
R1662 B.n164 B.t17 320.842
R1663 B.n1062 B.n1061 256.663
R1664 B.n1062 B.n161 256.663
R1665 B.n1062 B.n160 256.663
R1666 B.n1062 B.n159 256.663
R1667 B.n1062 B.n158 256.663
R1668 B.n1062 B.n157 256.663
R1669 B.n1062 B.n156 256.663
R1670 B.n1062 B.n155 256.663
R1671 B.n1062 B.n154 256.663
R1672 B.n1062 B.n153 256.663
R1673 B.n1062 B.n152 256.663
R1674 B.n1062 B.n151 256.663
R1675 B.n1062 B.n150 256.663
R1676 B.n1062 B.n149 256.663
R1677 B.n1062 B.n148 256.663
R1678 B.n1062 B.n147 256.663
R1679 B.n1062 B.n146 256.663
R1680 B.n1062 B.n145 256.663
R1681 B.n1062 B.n144 256.663
R1682 B.n1062 B.n143 256.663
R1683 B.n1062 B.n142 256.663
R1684 B.n1062 B.n141 256.663
R1685 B.n1062 B.n140 256.663
R1686 B.n1062 B.n139 256.663
R1687 B.n1062 B.n138 256.663
R1688 B.n1062 B.n137 256.663
R1689 B.n1062 B.n136 256.663
R1690 B.n1062 B.n135 256.663
R1691 B.n1062 B.n134 256.663
R1692 B.n1062 B.n133 256.663
R1693 B.n1062 B.n132 256.663
R1694 B.n1062 B.n131 256.663
R1695 B.n1062 B.n130 256.663
R1696 B.n1062 B.n129 256.663
R1697 B.n1062 B.n128 256.663
R1698 B.n1062 B.n127 256.663
R1699 B.n1062 B.n126 256.663
R1700 B.n1062 B.n125 256.663
R1701 B.n1062 B.n124 256.663
R1702 B.n1062 B.n123 256.663
R1703 B.n1062 B.n122 256.663
R1704 B.n1062 B.n121 256.663
R1705 B.n1062 B.n120 256.663
R1706 B.n1062 B.n119 256.663
R1707 B.n1062 B.n118 256.663
R1708 B.n1062 B.n117 256.663
R1709 B.n1062 B.n116 256.663
R1710 B.n1062 B.n115 256.663
R1711 B.n1062 B.n114 256.663
R1712 B.n1062 B.n113 256.663
R1713 B.n1062 B.n112 256.663
R1714 B.n1062 B.n111 256.663
R1715 B.n1062 B.n110 256.663
R1716 B.n1062 B.n109 256.663
R1717 B.n1062 B.n108 256.663
R1718 B.n1062 B.n107 256.663
R1719 B.n1062 B.n106 256.663
R1720 B.n1062 B.n105 256.663
R1721 B.n1062 B.n104 256.663
R1722 B.n1062 B.n103 256.663
R1723 B.n1063 B.n1062 256.663
R1724 B.n822 B.n821 256.663
R1725 B.n821 B.n516 256.663
R1726 B.n821 B.n517 256.663
R1727 B.n821 B.n518 256.663
R1728 B.n821 B.n519 256.663
R1729 B.n821 B.n520 256.663
R1730 B.n821 B.n521 256.663
R1731 B.n821 B.n522 256.663
R1732 B.n821 B.n523 256.663
R1733 B.n821 B.n524 256.663
R1734 B.n821 B.n525 256.663
R1735 B.n821 B.n526 256.663
R1736 B.n821 B.n527 256.663
R1737 B.n821 B.n528 256.663
R1738 B.n821 B.n529 256.663
R1739 B.n821 B.n530 256.663
R1740 B.n821 B.n531 256.663
R1741 B.n821 B.n532 256.663
R1742 B.n821 B.n533 256.663
R1743 B.n821 B.n534 256.663
R1744 B.n821 B.n535 256.663
R1745 B.n821 B.n536 256.663
R1746 B.n821 B.n537 256.663
R1747 B.n821 B.n538 256.663
R1748 B.n821 B.n539 256.663
R1749 B.n821 B.n540 256.663
R1750 B.n821 B.n541 256.663
R1751 B.n821 B.n542 256.663
R1752 B.n821 B.n543 256.663
R1753 B.n821 B.n544 256.663
R1754 B.n821 B.n545 256.663
R1755 B.n821 B.n546 256.663
R1756 B.n821 B.n547 256.663
R1757 B.n821 B.n548 256.663
R1758 B.n821 B.n549 256.663
R1759 B.n821 B.n550 256.663
R1760 B.n821 B.n551 256.663
R1761 B.n821 B.n552 256.663
R1762 B.n821 B.n553 256.663
R1763 B.n821 B.n554 256.663
R1764 B.n821 B.n555 256.663
R1765 B.n821 B.n556 256.663
R1766 B.n821 B.n557 256.663
R1767 B.n821 B.n558 256.663
R1768 B.n821 B.n559 256.663
R1769 B.n821 B.n560 256.663
R1770 B.n821 B.n561 256.663
R1771 B.n821 B.n562 256.663
R1772 B.n821 B.n563 256.663
R1773 B.n821 B.n564 256.663
R1774 B.n821 B.n565 256.663
R1775 B.n821 B.n566 256.663
R1776 B.n821 B.n567 256.663
R1777 B.n821 B.n568 256.663
R1778 B.n821 B.n569 256.663
R1779 B.n821 B.n570 256.663
R1780 B.n821 B.n571 256.663
R1781 B.n821 B.n572 256.663
R1782 B.n821 B.n573 256.663
R1783 B.n821 B.n574 256.663
R1784 B.n827 B.n513 163.367
R1785 B.n827 B.n507 163.367
R1786 B.n835 B.n507 163.367
R1787 B.n835 B.n505 163.367
R1788 B.n839 B.n505 163.367
R1789 B.n839 B.n499 163.367
R1790 B.n847 B.n499 163.367
R1791 B.n847 B.n497 163.367
R1792 B.n851 B.n497 163.367
R1793 B.n851 B.n491 163.367
R1794 B.n859 B.n491 163.367
R1795 B.n859 B.n489 163.367
R1796 B.n863 B.n489 163.367
R1797 B.n863 B.n483 163.367
R1798 B.n871 B.n483 163.367
R1799 B.n871 B.n481 163.367
R1800 B.n875 B.n481 163.367
R1801 B.n875 B.n475 163.367
R1802 B.n883 B.n475 163.367
R1803 B.n883 B.n473 163.367
R1804 B.n887 B.n473 163.367
R1805 B.n887 B.n467 163.367
R1806 B.n896 B.n467 163.367
R1807 B.n896 B.n465 163.367
R1808 B.n900 B.n465 163.367
R1809 B.n900 B.n460 163.367
R1810 B.n908 B.n460 163.367
R1811 B.n908 B.n458 163.367
R1812 B.n912 B.n458 163.367
R1813 B.n912 B.n452 163.367
R1814 B.n920 B.n452 163.367
R1815 B.n920 B.n450 163.367
R1816 B.n924 B.n450 163.367
R1817 B.n924 B.n444 163.367
R1818 B.n932 B.n444 163.367
R1819 B.n932 B.n442 163.367
R1820 B.n936 B.n442 163.367
R1821 B.n936 B.n436 163.367
R1822 B.n944 B.n436 163.367
R1823 B.n944 B.n434 163.367
R1824 B.n948 B.n434 163.367
R1825 B.n948 B.n428 163.367
R1826 B.n956 B.n428 163.367
R1827 B.n956 B.n426 163.367
R1828 B.n960 B.n426 163.367
R1829 B.n960 B.n420 163.367
R1830 B.n968 B.n420 163.367
R1831 B.n968 B.n418 163.367
R1832 B.n972 B.n418 163.367
R1833 B.n972 B.n412 163.367
R1834 B.n981 B.n412 163.367
R1835 B.n981 B.n410 163.367
R1836 B.n985 B.n410 163.367
R1837 B.n985 B.n2 163.367
R1838 B.n1176 B.n2 163.367
R1839 B.n1176 B.n3 163.367
R1840 B.n1172 B.n3 163.367
R1841 B.n1172 B.n9 163.367
R1842 B.n1168 B.n9 163.367
R1843 B.n1168 B.n11 163.367
R1844 B.n1164 B.n11 163.367
R1845 B.n1164 B.n16 163.367
R1846 B.n1160 B.n16 163.367
R1847 B.n1160 B.n18 163.367
R1848 B.n1156 B.n18 163.367
R1849 B.n1156 B.n23 163.367
R1850 B.n1152 B.n23 163.367
R1851 B.n1152 B.n25 163.367
R1852 B.n1148 B.n25 163.367
R1853 B.n1148 B.n30 163.367
R1854 B.n1144 B.n30 163.367
R1855 B.n1144 B.n32 163.367
R1856 B.n1140 B.n32 163.367
R1857 B.n1140 B.n37 163.367
R1858 B.n1136 B.n37 163.367
R1859 B.n1136 B.n39 163.367
R1860 B.n1132 B.n39 163.367
R1861 B.n1132 B.n44 163.367
R1862 B.n1128 B.n44 163.367
R1863 B.n1128 B.n46 163.367
R1864 B.n1124 B.n46 163.367
R1865 B.n1124 B.n51 163.367
R1866 B.n1120 B.n51 163.367
R1867 B.n1120 B.n53 163.367
R1868 B.n1116 B.n53 163.367
R1869 B.n1116 B.n57 163.367
R1870 B.n1112 B.n57 163.367
R1871 B.n1112 B.n59 163.367
R1872 B.n1108 B.n59 163.367
R1873 B.n1108 B.n65 163.367
R1874 B.n1104 B.n65 163.367
R1875 B.n1104 B.n67 163.367
R1876 B.n1100 B.n67 163.367
R1877 B.n1100 B.n72 163.367
R1878 B.n1096 B.n72 163.367
R1879 B.n1096 B.n74 163.367
R1880 B.n1092 B.n74 163.367
R1881 B.n1092 B.n79 163.367
R1882 B.n1088 B.n79 163.367
R1883 B.n1088 B.n81 163.367
R1884 B.n1084 B.n81 163.367
R1885 B.n1084 B.n86 163.367
R1886 B.n1080 B.n86 163.367
R1887 B.n1080 B.n88 163.367
R1888 B.n1076 B.n88 163.367
R1889 B.n1076 B.n93 163.367
R1890 B.n1072 B.n93 163.367
R1891 B.n1072 B.n95 163.367
R1892 B.n1068 B.n95 163.367
R1893 B.n1068 B.n100 163.367
R1894 B.n820 B.n515 163.367
R1895 B.n820 B.n576 163.367
R1896 B.n816 B.n815 163.367
R1897 B.n812 B.n811 163.367
R1898 B.n808 B.n807 163.367
R1899 B.n804 B.n803 163.367
R1900 B.n800 B.n799 163.367
R1901 B.n796 B.n795 163.367
R1902 B.n792 B.n791 163.367
R1903 B.n788 B.n787 163.367
R1904 B.n784 B.n783 163.367
R1905 B.n780 B.n779 163.367
R1906 B.n776 B.n775 163.367
R1907 B.n772 B.n771 163.367
R1908 B.n768 B.n767 163.367
R1909 B.n764 B.n763 163.367
R1910 B.n760 B.n759 163.367
R1911 B.n756 B.n755 163.367
R1912 B.n752 B.n751 163.367
R1913 B.n748 B.n747 163.367
R1914 B.n744 B.n743 163.367
R1915 B.n740 B.n739 163.367
R1916 B.n736 B.n735 163.367
R1917 B.n732 B.n731 163.367
R1918 B.n728 B.n727 163.367
R1919 B.n724 B.n723 163.367
R1920 B.n720 B.n719 163.367
R1921 B.n716 B.n715 163.367
R1922 B.n711 B.n710 163.367
R1923 B.n707 B.n706 163.367
R1924 B.n703 B.n702 163.367
R1925 B.n699 B.n698 163.367
R1926 B.n695 B.n694 163.367
R1927 B.n690 B.n689 163.367
R1928 B.n686 B.n685 163.367
R1929 B.n682 B.n681 163.367
R1930 B.n678 B.n677 163.367
R1931 B.n674 B.n673 163.367
R1932 B.n670 B.n669 163.367
R1933 B.n666 B.n665 163.367
R1934 B.n662 B.n661 163.367
R1935 B.n658 B.n657 163.367
R1936 B.n654 B.n653 163.367
R1937 B.n650 B.n649 163.367
R1938 B.n646 B.n645 163.367
R1939 B.n642 B.n641 163.367
R1940 B.n638 B.n637 163.367
R1941 B.n634 B.n633 163.367
R1942 B.n630 B.n629 163.367
R1943 B.n626 B.n625 163.367
R1944 B.n622 B.n621 163.367
R1945 B.n618 B.n617 163.367
R1946 B.n614 B.n613 163.367
R1947 B.n610 B.n609 163.367
R1948 B.n606 B.n605 163.367
R1949 B.n602 B.n601 163.367
R1950 B.n598 B.n597 163.367
R1951 B.n594 B.n593 163.367
R1952 B.n590 B.n589 163.367
R1953 B.n586 B.n585 163.367
R1954 B.n582 B.n575 163.367
R1955 B.n829 B.n511 163.367
R1956 B.n829 B.n509 163.367
R1957 B.n833 B.n509 163.367
R1958 B.n833 B.n503 163.367
R1959 B.n841 B.n503 163.367
R1960 B.n841 B.n501 163.367
R1961 B.n845 B.n501 163.367
R1962 B.n845 B.n495 163.367
R1963 B.n853 B.n495 163.367
R1964 B.n853 B.n493 163.367
R1965 B.n857 B.n493 163.367
R1966 B.n857 B.n487 163.367
R1967 B.n865 B.n487 163.367
R1968 B.n865 B.n485 163.367
R1969 B.n869 B.n485 163.367
R1970 B.n869 B.n479 163.367
R1971 B.n877 B.n479 163.367
R1972 B.n877 B.n477 163.367
R1973 B.n881 B.n477 163.367
R1974 B.n881 B.n471 163.367
R1975 B.n889 B.n471 163.367
R1976 B.n889 B.n469 163.367
R1977 B.n893 B.n469 163.367
R1978 B.n893 B.n464 163.367
R1979 B.n902 B.n464 163.367
R1980 B.n902 B.n462 163.367
R1981 B.n906 B.n462 163.367
R1982 B.n906 B.n456 163.367
R1983 B.n914 B.n456 163.367
R1984 B.n914 B.n454 163.367
R1985 B.n918 B.n454 163.367
R1986 B.n918 B.n448 163.367
R1987 B.n926 B.n448 163.367
R1988 B.n926 B.n446 163.367
R1989 B.n930 B.n446 163.367
R1990 B.n930 B.n440 163.367
R1991 B.n938 B.n440 163.367
R1992 B.n938 B.n438 163.367
R1993 B.n942 B.n438 163.367
R1994 B.n942 B.n432 163.367
R1995 B.n950 B.n432 163.367
R1996 B.n950 B.n430 163.367
R1997 B.n954 B.n430 163.367
R1998 B.n954 B.n424 163.367
R1999 B.n962 B.n424 163.367
R2000 B.n962 B.n422 163.367
R2001 B.n966 B.n422 163.367
R2002 B.n966 B.n416 163.367
R2003 B.n974 B.n416 163.367
R2004 B.n974 B.n414 163.367
R2005 B.n979 B.n414 163.367
R2006 B.n979 B.n408 163.367
R2007 B.n987 B.n408 163.367
R2008 B.n988 B.n987 163.367
R2009 B.n988 B.n5 163.367
R2010 B.n6 B.n5 163.367
R2011 B.n7 B.n6 163.367
R2012 B.n993 B.n7 163.367
R2013 B.n993 B.n12 163.367
R2014 B.n13 B.n12 163.367
R2015 B.n14 B.n13 163.367
R2016 B.n998 B.n14 163.367
R2017 B.n998 B.n19 163.367
R2018 B.n20 B.n19 163.367
R2019 B.n21 B.n20 163.367
R2020 B.n1003 B.n21 163.367
R2021 B.n1003 B.n26 163.367
R2022 B.n27 B.n26 163.367
R2023 B.n28 B.n27 163.367
R2024 B.n1008 B.n28 163.367
R2025 B.n1008 B.n33 163.367
R2026 B.n34 B.n33 163.367
R2027 B.n35 B.n34 163.367
R2028 B.n1013 B.n35 163.367
R2029 B.n1013 B.n40 163.367
R2030 B.n41 B.n40 163.367
R2031 B.n42 B.n41 163.367
R2032 B.n1018 B.n42 163.367
R2033 B.n1018 B.n47 163.367
R2034 B.n48 B.n47 163.367
R2035 B.n49 B.n48 163.367
R2036 B.n1023 B.n49 163.367
R2037 B.n1023 B.n54 163.367
R2038 B.n55 B.n54 163.367
R2039 B.n56 B.n55 163.367
R2040 B.n1028 B.n56 163.367
R2041 B.n1028 B.n61 163.367
R2042 B.n62 B.n61 163.367
R2043 B.n63 B.n62 163.367
R2044 B.n1033 B.n63 163.367
R2045 B.n1033 B.n68 163.367
R2046 B.n69 B.n68 163.367
R2047 B.n70 B.n69 163.367
R2048 B.n1038 B.n70 163.367
R2049 B.n1038 B.n75 163.367
R2050 B.n76 B.n75 163.367
R2051 B.n77 B.n76 163.367
R2052 B.n1043 B.n77 163.367
R2053 B.n1043 B.n82 163.367
R2054 B.n83 B.n82 163.367
R2055 B.n84 B.n83 163.367
R2056 B.n1048 B.n84 163.367
R2057 B.n1048 B.n89 163.367
R2058 B.n90 B.n89 163.367
R2059 B.n91 B.n90 163.367
R2060 B.n1053 B.n91 163.367
R2061 B.n1053 B.n96 163.367
R2062 B.n97 B.n96 163.367
R2063 B.n98 B.n97 163.367
R2064 B.n163 B.n98 163.367
R2065 B.n170 B.n102 163.367
R2066 B.n174 B.n173 163.367
R2067 B.n178 B.n177 163.367
R2068 B.n182 B.n181 163.367
R2069 B.n186 B.n185 163.367
R2070 B.n190 B.n189 163.367
R2071 B.n194 B.n193 163.367
R2072 B.n198 B.n197 163.367
R2073 B.n202 B.n201 163.367
R2074 B.n206 B.n205 163.367
R2075 B.n210 B.n209 163.367
R2076 B.n214 B.n213 163.367
R2077 B.n218 B.n217 163.367
R2078 B.n222 B.n221 163.367
R2079 B.n226 B.n225 163.367
R2080 B.n230 B.n229 163.367
R2081 B.n234 B.n233 163.367
R2082 B.n238 B.n237 163.367
R2083 B.n242 B.n241 163.367
R2084 B.n246 B.n245 163.367
R2085 B.n250 B.n249 163.367
R2086 B.n254 B.n253 163.367
R2087 B.n258 B.n257 163.367
R2088 B.n262 B.n261 163.367
R2089 B.n266 B.n265 163.367
R2090 B.n270 B.n269 163.367
R2091 B.n274 B.n273 163.367
R2092 B.n278 B.n277 163.367
R2093 B.n282 B.n281 163.367
R2094 B.n286 B.n285 163.367
R2095 B.n290 B.n289 163.367
R2096 B.n294 B.n293 163.367
R2097 B.n298 B.n297 163.367
R2098 B.n302 B.n301 163.367
R2099 B.n306 B.n305 163.367
R2100 B.n310 B.n309 163.367
R2101 B.n314 B.n313 163.367
R2102 B.n318 B.n317 163.367
R2103 B.n322 B.n321 163.367
R2104 B.n326 B.n325 163.367
R2105 B.n330 B.n329 163.367
R2106 B.n334 B.n333 163.367
R2107 B.n338 B.n337 163.367
R2108 B.n342 B.n341 163.367
R2109 B.n346 B.n345 163.367
R2110 B.n350 B.n349 163.367
R2111 B.n354 B.n353 163.367
R2112 B.n358 B.n357 163.367
R2113 B.n362 B.n361 163.367
R2114 B.n366 B.n365 163.367
R2115 B.n370 B.n369 163.367
R2116 B.n374 B.n373 163.367
R2117 B.n378 B.n377 163.367
R2118 B.n382 B.n381 163.367
R2119 B.n386 B.n385 163.367
R2120 B.n390 B.n389 163.367
R2121 B.n394 B.n393 163.367
R2122 B.n398 B.n397 163.367
R2123 B.n402 B.n401 163.367
R2124 B.n404 B.n162 163.367
R2125 B.n580 B.n579 77.3823
R2126 B.n578 B.n577 77.3823
R2127 B.n168 B.n167 77.3823
R2128 B.n165 B.n164 77.3823
R2129 B.n823 B.n822 71.676
R2130 B.n576 B.n516 71.676
R2131 B.n815 B.n517 71.676
R2132 B.n811 B.n518 71.676
R2133 B.n807 B.n519 71.676
R2134 B.n803 B.n520 71.676
R2135 B.n799 B.n521 71.676
R2136 B.n795 B.n522 71.676
R2137 B.n791 B.n523 71.676
R2138 B.n787 B.n524 71.676
R2139 B.n783 B.n525 71.676
R2140 B.n779 B.n526 71.676
R2141 B.n775 B.n527 71.676
R2142 B.n771 B.n528 71.676
R2143 B.n767 B.n529 71.676
R2144 B.n763 B.n530 71.676
R2145 B.n759 B.n531 71.676
R2146 B.n755 B.n532 71.676
R2147 B.n751 B.n533 71.676
R2148 B.n747 B.n534 71.676
R2149 B.n743 B.n535 71.676
R2150 B.n739 B.n536 71.676
R2151 B.n735 B.n537 71.676
R2152 B.n731 B.n538 71.676
R2153 B.n727 B.n539 71.676
R2154 B.n723 B.n540 71.676
R2155 B.n719 B.n541 71.676
R2156 B.n715 B.n542 71.676
R2157 B.n710 B.n543 71.676
R2158 B.n706 B.n544 71.676
R2159 B.n702 B.n545 71.676
R2160 B.n698 B.n546 71.676
R2161 B.n694 B.n547 71.676
R2162 B.n689 B.n548 71.676
R2163 B.n685 B.n549 71.676
R2164 B.n681 B.n550 71.676
R2165 B.n677 B.n551 71.676
R2166 B.n673 B.n552 71.676
R2167 B.n669 B.n553 71.676
R2168 B.n665 B.n554 71.676
R2169 B.n661 B.n555 71.676
R2170 B.n657 B.n556 71.676
R2171 B.n653 B.n557 71.676
R2172 B.n649 B.n558 71.676
R2173 B.n645 B.n559 71.676
R2174 B.n641 B.n560 71.676
R2175 B.n637 B.n561 71.676
R2176 B.n633 B.n562 71.676
R2177 B.n629 B.n563 71.676
R2178 B.n625 B.n564 71.676
R2179 B.n621 B.n565 71.676
R2180 B.n617 B.n566 71.676
R2181 B.n613 B.n567 71.676
R2182 B.n609 B.n568 71.676
R2183 B.n605 B.n569 71.676
R2184 B.n601 B.n570 71.676
R2185 B.n597 B.n571 71.676
R2186 B.n593 B.n572 71.676
R2187 B.n589 B.n573 71.676
R2188 B.n585 B.n574 71.676
R2189 B.n1064 B.n1063 71.676
R2190 B.n170 B.n103 71.676
R2191 B.n174 B.n104 71.676
R2192 B.n178 B.n105 71.676
R2193 B.n182 B.n106 71.676
R2194 B.n186 B.n107 71.676
R2195 B.n190 B.n108 71.676
R2196 B.n194 B.n109 71.676
R2197 B.n198 B.n110 71.676
R2198 B.n202 B.n111 71.676
R2199 B.n206 B.n112 71.676
R2200 B.n210 B.n113 71.676
R2201 B.n214 B.n114 71.676
R2202 B.n218 B.n115 71.676
R2203 B.n222 B.n116 71.676
R2204 B.n226 B.n117 71.676
R2205 B.n230 B.n118 71.676
R2206 B.n234 B.n119 71.676
R2207 B.n238 B.n120 71.676
R2208 B.n242 B.n121 71.676
R2209 B.n246 B.n122 71.676
R2210 B.n250 B.n123 71.676
R2211 B.n254 B.n124 71.676
R2212 B.n258 B.n125 71.676
R2213 B.n262 B.n126 71.676
R2214 B.n266 B.n127 71.676
R2215 B.n270 B.n128 71.676
R2216 B.n274 B.n129 71.676
R2217 B.n278 B.n130 71.676
R2218 B.n282 B.n131 71.676
R2219 B.n286 B.n132 71.676
R2220 B.n290 B.n133 71.676
R2221 B.n294 B.n134 71.676
R2222 B.n298 B.n135 71.676
R2223 B.n302 B.n136 71.676
R2224 B.n306 B.n137 71.676
R2225 B.n310 B.n138 71.676
R2226 B.n314 B.n139 71.676
R2227 B.n318 B.n140 71.676
R2228 B.n322 B.n141 71.676
R2229 B.n326 B.n142 71.676
R2230 B.n330 B.n143 71.676
R2231 B.n334 B.n144 71.676
R2232 B.n338 B.n145 71.676
R2233 B.n342 B.n146 71.676
R2234 B.n346 B.n147 71.676
R2235 B.n350 B.n148 71.676
R2236 B.n354 B.n149 71.676
R2237 B.n358 B.n150 71.676
R2238 B.n362 B.n151 71.676
R2239 B.n366 B.n152 71.676
R2240 B.n370 B.n153 71.676
R2241 B.n374 B.n154 71.676
R2242 B.n378 B.n155 71.676
R2243 B.n382 B.n156 71.676
R2244 B.n386 B.n157 71.676
R2245 B.n390 B.n158 71.676
R2246 B.n394 B.n159 71.676
R2247 B.n398 B.n160 71.676
R2248 B.n402 B.n161 71.676
R2249 B.n1061 B.n162 71.676
R2250 B.n1061 B.n1060 71.676
R2251 B.n404 B.n161 71.676
R2252 B.n401 B.n160 71.676
R2253 B.n397 B.n159 71.676
R2254 B.n393 B.n158 71.676
R2255 B.n389 B.n157 71.676
R2256 B.n385 B.n156 71.676
R2257 B.n381 B.n155 71.676
R2258 B.n377 B.n154 71.676
R2259 B.n373 B.n153 71.676
R2260 B.n369 B.n152 71.676
R2261 B.n365 B.n151 71.676
R2262 B.n361 B.n150 71.676
R2263 B.n357 B.n149 71.676
R2264 B.n353 B.n148 71.676
R2265 B.n349 B.n147 71.676
R2266 B.n345 B.n146 71.676
R2267 B.n341 B.n145 71.676
R2268 B.n337 B.n144 71.676
R2269 B.n333 B.n143 71.676
R2270 B.n329 B.n142 71.676
R2271 B.n325 B.n141 71.676
R2272 B.n321 B.n140 71.676
R2273 B.n317 B.n139 71.676
R2274 B.n313 B.n138 71.676
R2275 B.n309 B.n137 71.676
R2276 B.n305 B.n136 71.676
R2277 B.n301 B.n135 71.676
R2278 B.n297 B.n134 71.676
R2279 B.n293 B.n133 71.676
R2280 B.n289 B.n132 71.676
R2281 B.n285 B.n131 71.676
R2282 B.n281 B.n130 71.676
R2283 B.n277 B.n129 71.676
R2284 B.n273 B.n128 71.676
R2285 B.n269 B.n127 71.676
R2286 B.n265 B.n126 71.676
R2287 B.n261 B.n125 71.676
R2288 B.n257 B.n124 71.676
R2289 B.n253 B.n123 71.676
R2290 B.n249 B.n122 71.676
R2291 B.n245 B.n121 71.676
R2292 B.n241 B.n120 71.676
R2293 B.n237 B.n119 71.676
R2294 B.n233 B.n118 71.676
R2295 B.n229 B.n117 71.676
R2296 B.n225 B.n116 71.676
R2297 B.n221 B.n115 71.676
R2298 B.n217 B.n114 71.676
R2299 B.n213 B.n113 71.676
R2300 B.n209 B.n112 71.676
R2301 B.n205 B.n111 71.676
R2302 B.n201 B.n110 71.676
R2303 B.n197 B.n109 71.676
R2304 B.n193 B.n108 71.676
R2305 B.n189 B.n107 71.676
R2306 B.n185 B.n106 71.676
R2307 B.n181 B.n105 71.676
R2308 B.n177 B.n104 71.676
R2309 B.n173 B.n103 71.676
R2310 B.n1063 B.n102 71.676
R2311 B.n822 B.n515 71.676
R2312 B.n816 B.n516 71.676
R2313 B.n812 B.n517 71.676
R2314 B.n808 B.n518 71.676
R2315 B.n804 B.n519 71.676
R2316 B.n800 B.n520 71.676
R2317 B.n796 B.n521 71.676
R2318 B.n792 B.n522 71.676
R2319 B.n788 B.n523 71.676
R2320 B.n784 B.n524 71.676
R2321 B.n780 B.n525 71.676
R2322 B.n776 B.n526 71.676
R2323 B.n772 B.n527 71.676
R2324 B.n768 B.n528 71.676
R2325 B.n764 B.n529 71.676
R2326 B.n760 B.n530 71.676
R2327 B.n756 B.n531 71.676
R2328 B.n752 B.n532 71.676
R2329 B.n748 B.n533 71.676
R2330 B.n744 B.n534 71.676
R2331 B.n740 B.n535 71.676
R2332 B.n736 B.n536 71.676
R2333 B.n732 B.n537 71.676
R2334 B.n728 B.n538 71.676
R2335 B.n724 B.n539 71.676
R2336 B.n720 B.n540 71.676
R2337 B.n716 B.n541 71.676
R2338 B.n711 B.n542 71.676
R2339 B.n707 B.n543 71.676
R2340 B.n703 B.n544 71.676
R2341 B.n699 B.n545 71.676
R2342 B.n695 B.n546 71.676
R2343 B.n690 B.n547 71.676
R2344 B.n686 B.n548 71.676
R2345 B.n682 B.n549 71.676
R2346 B.n678 B.n550 71.676
R2347 B.n674 B.n551 71.676
R2348 B.n670 B.n552 71.676
R2349 B.n666 B.n553 71.676
R2350 B.n662 B.n554 71.676
R2351 B.n658 B.n555 71.676
R2352 B.n654 B.n556 71.676
R2353 B.n650 B.n557 71.676
R2354 B.n646 B.n558 71.676
R2355 B.n642 B.n559 71.676
R2356 B.n638 B.n560 71.676
R2357 B.n634 B.n561 71.676
R2358 B.n630 B.n562 71.676
R2359 B.n626 B.n563 71.676
R2360 B.n622 B.n564 71.676
R2361 B.n618 B.n565 71.676
R2362 B.n614 B.n566 71.676
R2363 B.n610 B.n567 71.676
R2364 B.n606 B.n568 71.676
R2365 B.n602 B.n569 71.676
R2366 B.n598 B.n570 71.676
R2367 B.n594 B.n571 71.676
R2368 B.n590 B.n572 71.676
R2369 B.n586 B.n573 71.676
R2370 B.n582 B.n574 71.676
R2371 B.n821 B.n512 62.8576
R2372 B.n1062 B.n99 62.8576
R2373 B.n692 B.n580 59.5399
R2374 B.n713 B.n578 59.5399
R2375 B.n169 B.n168 59.5399
R2376 B.n166 B.n165 59.5399
R2377 B.n828 B.n512 33.6563
R2378 B.n828 B.n508 33.6563
R2379 B.n834 B.n508 33.6563
R2380 B.n834 B.n504 33.6563
R2381 B.n840 B.n504 33.6563
R2382 B.n840 B.n500 33.6563
R2383 B.n846 B.n500 33.6563
R2384 B.n846 B.n496 33.6563
R2385 B.n852 B.n496 33.6563
R2386 B.n858 B.n492 33.6563
R2387 B.n858 B.n488 33.6563
R2388 B.n864 B.n488 33.6563
R2389 B.n864 B.n484 33.6563
R2390 B.n870 B.n484 33.6563
R2391 B.n870 B.n480 33.6563
R2392 B.n876 B.n480 33.6563
R2393 B.n876 B.n476 33.6563
R2394 B.n882 B.n476 33.6563
R2395 B.n882 B.n472 33.6563
R2396 B.n888 B.n472 33.6563
R2397 B.n888 B.n468 33.6563
R2398 B.n895 B.n468 33.6563
R2399 B.n895 B.n894 33.6563
R2400 B.n901 B.n461 33.6563
R2401 B.n907 B.n461 33.6563
R2402 B.n907 B.n457 33.6563
R2403 B.n913 B.n457 33.6563
R2404 B.n913 B.n453 33.6563
R2405 B.n919 B.n453 33.6563
R2406 B.n919 B.n449 33.6563
R2407 B.n925 B.n449 33.6563
R2408 B.n925 B.n445 33.6563
R2409 B.n931 B.n445 33.6563
R2410 B.n937 B.n441 33.6563
R2411 B.n937 B.n437 33.6563
R2412 B.n943 B.n437 33.6563
R2413 B.n943 B.n433 33.6563
R2414 B.n949 B.n433 33.6563
R2415 B.n949 B.n429 33.6563
R2416 B.n955 B.n429 33.6563
R2417 B.n955 B.n425 33.6563
R2418 B.n961 B.n425 33.6563
R2419 B.n961 B.n421 33.6563
R2420 B.n967 B.n421 33.6563
R2421 B.n973 B.n417 33.6563
R2422 B.n973 B.n413 33.6563
R2423 B.n980 B.n413 33.6563
R2424 B.n980 B.n409 33.6563
R2425 B.n986 B.n409 33.6563
R2426 B.n986 B.n4 33.6563
R2427 B.n1175 B.n4 33.6563
R2428 B.n1175 B.n1174 33.6563
R2429 B.n1174 B.n1173 33.6563
R2430 B.n1173 B.n8 33.6563
R2431 B.n1167 B.n8 33.6563
R2432 B.n1167 B.n1166 33.6563
R2433 B.n1166 B.n1165 33.6563
R2434 B.n1165 B.n15 33.6563
R2435 B.n1159 B.n1158 33.6563
R2436 B.n1158 B.n1157 33.6563
R2437 B.n1157 B.n22 33.6563
R2438 B.n1151 B.n22 33.6563
R2439 B.n1151 B.n1150 33.6563
R2440 B.n1150 B.n1149 33.6563
R2441 B.n1149 B.n29 33.6563
R2442 B.n1143 B.n29 33.6563
R2443 B.n1143 B.n1142 33.6563
R2444 B.n1142 B.n1141 33.6563
R2445 B.n1141 B.n36 33.6563
R2446 B.n1135 B.n1134 33.6563
R2447 B.n1134 B.n1133 33.6563
R2448 B.n1133 B.n43 33.6563
R2449 B.n1127 B.n43 33.6563
R2450 B.n1127 B.n1126 33.6563
R2451 B.n1126 B.n1125 33.6563
R2452 B.n1125 B.n50 33.6563
R2453 B.n1119 B.n50 33.6563
R2454 B.n1119 B.n1118 33.6563
R2455 B.n1118 B.n1117 33.6563
R2456 B.n1111 B.n60 33.6563
R2457 B.n1111 B.n1110 33.6563
R2458 B.n1110 B.n1109 33.6563
R2459 B.n1109 B.n64 33.6563
R2460 B.n1103 B.n64 33.6563
R2461 B.n1103 B.n1102 33.6563
R2462 B.n1102 B.n1101 33.6563
R2463 B.n1101 B.n71 33.6563
R2464 B.n1095 B.n71 33.6563
R2465 B.n1095 B.n1094 33.6563
R2466 B.n1094 B.n1093 33.6563
R2467 B.n1093 B.n78 33.6563
R2468 B.n1087 B.n78 33.6563
R2469 B.n1087 B.n1086 33.6563
R2470 B.n1085 B.n85 33.6563
R2471 B.n1079 B.n85 33.6563
R2472 B.n1079 B.n1078 33.6563
R2473 B.n1078 B.n1077 33.6563
R2474 B.n1077 B.n92 33.6563
R2475 B.n1071 B.n92 33.6563
R2476 B.n1071 B.n1070 33.6563
R2477 B.n1070 B.n1069 33.6563
R2478 B.n1069 B.n99 33.6563
R2479 B.n1066 B.n1065 32.6249
R2480 B.n1059 B.n1058 32.6249
R2481 B.n581 B.n510 32.6249
R2482 B.n825 B.n824 32.6249
R2483 B.n901 B.t0 31.6765
R2484 B.n1117 B.t2 31.6765
R2485 B.t7 B.n492 29.6968
R2486 B.n1086 B.t11 29.6968
R2487 B.n931 B.t5 26.7272
R2488 B.n1135 B.t1 26.7272
R2489 B B.n1177 18.0485
R2490 B.n967 B.t4 17.8183
R2491 B.n1159 B.t3 17.8183
R2492 B.t4 B.n417 15.8385
R2493 B.t3 B.n15 15.8385
R2494 B.n1065 B.n101 10.6151
R2495 B.n171 B.n101 10.6151
R2496 B.n172 B.n171 10.6151
R2497 B.n175 B.n172 10.6151
R2498 B.n176 B.n175 10.6151
R2499 B.n179 B.n176 10.6151
R2500 B.n180 B.n179 10.6151
R2501 B.n183 B.n180 10.6151
R2502 B.n184 B.n183 10.6151
R2503 B.n187 B.n184 10.6151
R2504 B.n188 B.n187 10.6151
R2505 B.n191 B.n188 10.6151
R2506 B.n192 B.n191 10.6151
R2507 B.n195 B.n192 10.6151
R2508 B.n196 B.n195 10.6151
R2509 B.n199 B.n196 10.6151
R2510 B.n200 B.n199 10.6151
R2511 B.n203 B.n200 10.6151
R2512 B.n204 B.n203 10.6151
R2513 B.n207 B.n204 10.6151
R2514 B.n208 B.n207 10.6151
R2515 B.n211 B.n208 10.6151
R2516 B.n212 B.n211 10.6151
R2517 B.n215 B.n212 10.6151
R2518 B.n216 B.n215 10.6151
R2519 B.n219 B.n216 10.6151
R2520 B.n220 B.n219 10.6151
R2521 B.n223 B.n220 10.6151
R2522 B.n224 B.n223 10.6151
R2523 B.n227 B.n224 10.6151
R2524 B.n228 B.n227 10.6151
R2525 B.n231 B.n228 10.6151
R2526 B.n232 B.n231 10.6151
R2527 B.n235 B.n232 10.6151
R2528 B.n236 B.n235 10.6151
R2529 B.n239 B.n236 10.6151
R2530 B.n240 B.n239 10.6151
R2531 B.n243 B.n240 10.6151
R2532 B.n244 B.n243 10.6151
R2533 B.n247 B.n244 10.6151
R2534 B.n248 B.n247 10.6151
R2535 B.n251 B.n248 10.6151
R2536 B.n252 B.n251 10.6151
R2537 B.n255 B.n252 10.6151
R2538 B.n256 B.n255 10.6151
R2539 B.n259 B.n256 10.6151
R2540 B.n260 B.n259 10.6151
R2541 B.n263 B.n260 10.6151
R2542 B.n264 B.n263 10.6151
R2543 B.n267 B.n264 10.6151
R2544 B.n268 B.n267 10.6151
R2545 B.n271 B.n268 10.6151
R2546 B.n272 B.n271 10.6151
R2547 B.n275 B.n272 10.6151
R2548 B.n276 B.n275 10.6151
R2549 B.n280 B.n279 10.6151
R2550 B.n283 B.n280 10.6151
R2551 B.n284 B.n283 10.6151
R2552 B.n287 B.n284 10.6151
R2553 B.n288 B.n287 10.6151
R2554 B.n291 B.n288 10.6151
R2555 B.n292 B.n291 10.6151
R2556 B.n295 B.n292 10.6151
R2557 B.n296 B.n295 10.6151
R2558 B.n300 B.n299 10.6151
R2559 B.n303 B.n300 10.6151
R2560 B.n304 B.n303 10.6151
R2561 B.n307 B.n304 10.6151
R2562 B.n308 B.n307 10.6151
R2563 B.n311 B.n308 10.6151
R2564 B.n312 B.n311 10.6151
R2565 B.n315 B.n312 10.6151
R2566 B.n316 B.n315 10.6151
R2567 B.n319 B.n316 10.6151
R2568 B.n320 B.n319 10.6151
R2569 B.n323 B.n320 10.6151
R2570 B.n324 B.n323 10.6151
R2571 B.n327 B.n324 10.6151
R2572 B.n328 B.n327 10.6151
R2573 B.n331 B.n328 10.6151
R2574 B.n332 B.n331 10.6151
R2575 B.n335 B.n332 10.6151
R2576 B.n336 B.n335 10.6151
R2577 B.n339 B.n336 10.6151
R2578 B.n340 B.n339 10.6151
R2579 B.n343 B.n340 10.6151
R2580 B.n344 B.n343 10.6151
R2581 B.n347 B.n344 10.6151
R2582 B.n348 B.n347 10.6151
R2583 B.n351 B.n348 10.6151
R2584 B.n352 B.n351 10.6151
R2585 B.n355 B.n352 10.6151
R2586 B.n356 B.n355 10.6151
R2587 B.n359 B.n356 10.6151
R2588 B.n360 B.n359 10.6151
R2589 B.n363 B.n360 10.6151
R2590 B.n364 B.n363 10.6151
R2591 B.n367 B.n364 10.6151
R2592 B.n368 B.n367 10.6151
R2593 B.n371 B.n368 10.6151
R2594 B.n372 B.n371 10.6151
R2595 B.n375 B.n372 10.6151
R2596 B.n376 B.n375 10.6151
R2597 B.n379 B.n376 10.6151
R2598 B.n380 B.n379 10.6151
R2599 B.n383 B.n380 10.6151
R2600 B.n384 B.n383 10.6151
R2601 B.n387 B.n384 10.6151
R2602 B.n388 B.n387 10.6151
R2603 B.n391 B.n388 10.6151
R2604 B.n392 B.n391 10.6151
R2605 B.n395 B.n392 10.6151
R2606 B.n396 B.n395 10.6151
R2607 B.n399 B.n396 10.6151
R2608 B.n400 B.n399 10.6151
R2609 B.n403 B.n400 10.6151
R2610 B.n405 B.n403 10.6151
R2611 B.n406 B.n405 10.6151
R2612 B.n1059 B.n406 10.6151
R2613 B.n830 B.n510 10.6151
R2614 B.n831 B.n830 10.6151
R2615 B.n832 B.n831 10.6151
R2616 B.n832 B.n502 10.6151
R2617 B.n842 B.n502 10.6151
R2618 B.n843 B.n842 10.6151
R2619 B.n844 B.n843 10.6151
R2620 B.n844 B.n494 10.6151
R2621 B.n854 B.n494 10.6151
R2622 B.n855 B.n854 10.6151
R2623 B.n856 B.n855 10.6151
R2624 B.n856 B.n486 10.6151
R2625 B.n866 B.n486 10.6151
R2626 B.n867 B.n866 10.6151
R2627 B.n868 B.n867 10.6151
R2628 B.n868 B.n478 10.6151
R2629 B.n878 B.n478 10.6151
R2630 B.n879 B.n878 10.6151
R2631 B.n880 B.n879 10.6151
R2632 B.n880 B.n470 10.6151
R2633 B.n890 B.n470 10.6151
R2634 B.n891 B.n890 10.6151
R2635 B.n892 B.n891 10.6151
R2636 B.n892 B.n463 10.6151
R2637 B.n903 B.n463 10.6151
R2638 B.n904 B.n903 10.6151
R2639 B.n905 B.n904 10.6151
R2640 B.n905 B.n455 10.6151
R2641 B.n915 B.n455 10.6151
R2642 B.n916 B.n915 10.6151
R2643 B.n917 B.n916 10.6151
R2644 B.n917 B.n447 10.6151
R2645 B.n927 B.n447 10.6151
R2646 B.n928 B.n927 10.6151
R2647 B.n929 B.n928 10.6151
R2648 B.n929 B.n439 10.6151
R2649 B.n939 B.n439 10.6151
R2650 B.n940 B.n939 10.6151
R2651 B.n941 B.n940 10.6151
R2652 B.n941 B.n431 10.6151
R2653 B.n951 B.n431 10.6151
R2654 B.n952 B.n951 10.6151
R2655 B.n953 B.n952 10.6151
R2656 B.n953 B.n423 10.6151
R2657 B.n963 B.n423 10.6151
R2658 B.n964 B.n963 10.6151
R2659 B.n965 B.n964 10.6151
R2660 B.n965 B.n415 10.6151
R2661 B.n975 B.n415 10.6151
R2662 B.n976 B.n975 10.6151
R2663 B.n978 B.n976 10.6151
R2664 B.n978 B.n977 10.6151
R2665 B.n977 B.n407 10.6151
R2666 B.n989 B.n407 10.6151
R2667 B.n990 B.n989 10.6151
R2668 B.n991 B.n990 10.6151
R2669 B.n992 B.n991 10.6151
R2670 B.n994 B.n992 10.6151
R2671 B.n995 B.n994 10.6151
R2672 B.n996 B.n995 10.6151
R2673 B.n997 B.n996 10.6151
R2674 B.n999 B.n997 10.6151
R2675 B.n1000 B.n999 10.6151
R2676 B.n1001 B.n1000 10.6151
R2677 B.n1002 B.n1001 10.6151
R2678 B.n1004 B.n1002 10.6151
R2679 B.n1005 B.n1004 10.6151
R2680 B.n1006 B.n1005 10.6151
R2681 B.n1007 B.n1006 10.6151
R2682 B.n1009 B.n1007 10.6151
R2683 B.n1010 B.n1009 10.6151
R2684 B.n1011 B.n1010 10.6151
R2685 B.n1012 B.n1011 10.6151
R2686 B.n1014 B.n1012 10.6151
R2687 B.n1015 B.n1014 10.6151
R2688 B.n1016 B.n1015 10.6151
R2689 B.n1017 B.n1016 10.6151
R2690 B.n1019 B.n1017 10.6151
R2691 B.n1020 B.n1019 10.6151
R2692 B.n1021 B.n1020 10.6151
R2693 B.n1022 B.n1021 10.6151
R2694 B.n1024 B.n1022 10.6151
R2695 B.n1025 B.n1024 10.6151
R2696 B.n1026 B.n1025 10.6151
R2697 B.n1027 B.n1026 10.6151
R2698 B.n1029 B.n1027 10.6151
R2699 B.n1030 B.n1029 10.6151
R2700 B.n1031 B.n1030 10.6151
R2701 B.n1032 B.n1031 10.6151
R2702 B.n1034 B.n1032 10.6151
R2703 B.n1035 B.n1034 10.6151
R2704 B.n1036 B.n1035 10.6151
R2705 B.n1037 B.n1036 10.6151
R2706 B.n1039 B.n1037 10.6151
R2707 B.n1040 B.n1039 10.6151
R2708 B.n1041 B.n1040 10.6151
R2709 B.n1042 B.n1041 10.6151
R2710 B.n1044 B.n1042 10.6151
R2711 B.n1045 B.n1044 10.6151
R2712 B.n1046 B.n1045 10.6151
R2713 B.n1047 B.n1046 10.6151
R2714 B.n1049 B.n1047 10.6151
R2715 B.n1050 B.n1049 10.6151
R2716 B.n1051 B.n1050 10.6151
R2717 B.n1052 B.n1051 10.6151
R2718 B.n1054 B.n1052 10.6151
R2719 B.n1055 B.n1054 10.6151
R2720 B.n1056 B.n1055 10.6151
R2721 B.n1057 B.n1056 10.6151
R2722 B.n1058 B.n1057 10.6151
R2723 B.n824 B.n514 10.6151
R2724 B.n819 B.n514 10.6151
R2725 B.n819 B.n818 10.6151
R2726 B.n818 B.n817 10.6151
R2727 B.n817 B.n814 10.6151
R2728 B.n814 B.n813 10.6151
R2729 B.n813 B.n810 10.6151
R2730 B.n810 B.n809 10.6151
R2731 B.n809 B.n806 10.6151
R2732 B.n806 B.n805 10.6151
R2733 B.n805 B.n802 10.6151
R2734 B.n802 B.n801 10.6151
R2735 B.n801 B.n798 10.6151
R2736 B.n798 B.n797 10.6151
R2737 B.n797 B.n794 10.6151
R2738 B.n794 B.n793 10.6151
R2739 B.n793 B.n790 10.6151
R2740 B.n790 B.n789 10.6151
R2741 B.n789 B.n786 10.6151
R2742 B.n786 B.n785 10.6151
R2743 B.n785 B.n782 10.6151
R2744 B.n782 B.n781 10.6151
R2745 B.n781 B.n778 10.6151
R2746 B.n778 B.n777 10.6151
R2747 B.n777 B.n774 10.6151
R2748 B.n774 B.n773 10.6151
R2749 B.n773 B.n770 10.6151
R2750 B.n770 B.n769 10.6151
R2751 B.n769 B.n766 10.6151
R2752 B.n766 B.n765 10.6151
R2753 B.n765 B.n762 10.6151
R2754 B.n762 B.n761 10.6151
R2755 B.n761 B.n758 10.6151
R2756 B.n758 B.n757 10.6151
R2757 B.n757 B.n754 10.6151
R2758 B.n754 B.n753 10.6151
R2759 B.n753 B.n750 10.6151
R2760 B.n750 B.n749 10.6151
R2761 B.n749 B.n746 10.6151
R2762 B.n746 B.n745 10.6151
R2763 B.n745 B.n742 10.6151
R2764 B.n742 B.n741 10.6151
R2765 B.n741 B.n738 10.6151
R2766 B.n738 B.n737 10.6151
R2767 B.n737 B.n734 10.6151
R2768 B.n734 B.n733 10.6151
R2769 B.n733 B.n730 10.6151
R2770 B.n730 B.n729 10.6151
R2771 B.n729 B.n726 10.6151
R2772 B.n726 B.n725 10.6151
R2773 B.n725 B.n722 10.6151
R2774 B.n722 B.n721 10.6151
R2775 B.n721 B.n718 10.6151
R2776 B.n718 B.n717 10.6151
R2777 B.n717 B.n714 10.6151
R2778 B.n712 B.n709 10.6151
R2779 B.n709 B.n708 10.6151
R2780 B.n708 B.n705 10.6151
R2781 B.n705 B.n704 10.6151
R2782 B.n704 B.n701 10.6151
R2783 B.n701 B.n700 10.6151
R2784 B.n700 B.n697 10.6151
R2785 B.n697 B.n696 10.6151
R2786 B.n696 B.n693 10.6151
R2787 B.n691 B.n688 10.6151
R2788 B.n688 B.n687 10.6151
R2789 B.n687 B.n684 10.6151
R2790 B.n684 B.n683 10.6151
R2791 B.n683 B.n680 10.6151
R2792 B.n680 B.n679 10.6151
R2793 B.n679 B.n676 10.6151
R2794 B.n676 B.n675 10.6151
R2795 B.n675 B.n672 10.6151
R2796 B.n672 B.n671 10.6151
R2797 B.n671 B.n668 10.6151
R2798 B.n668 B.n667 10.6151
R2799 B.n667 B.n664 10.6151
R2800 B.n664 B.n663 10.6151
R2801 B.n663 B.n660 10.6151
R2802 B.n660 B.n659 10.6151
R2803 B.n659 B.n656 10.6151
R2804 B.n656 B.n655 10.6151
R2805 B.n655 B.n652 10.6151
R2806 B.n652 B.n651 10.6151
R2807 B.n651 B.n648 10.6151
R2808 B.n648 B.n647 10.6151
R2809 B.n647 B.n644 10.6151
R2810 B.n644 B.n643 10.6151
R2811 B.n643 B.n640 10.6151
R2812 B.n640 B.n639 10.6151
R2813 B.n639 B.n636 10.6151
R2814 B.n636 B.n635 10.6151
R2815 B.n635 B.n632 10.6151
R2816 B.n632 B.n631 10.6151
R2817 B.n631 B.n628 10.6151
R2818 B.n628 B.n627 10.6151
R2819 B.n627 B.n624 10.6151
R2820 B.n624 B.n623 10.6151
R2821 B.n623 B.n620 10.6151
R2822 B.n620 B.n619 10.6151
R2823 B.n619 B.n616 10.6151
R2824 B.n616 B.n615 10.6151
R2825 B.n615 B.n612 10.6151
R2826 B.n612 B.n611 10.6151
R2827 B.n611 B.n608 10.6151
R2828 B.n608 B.n607 10.6151
R2829 B.n607 B.n604 10.6151
R2830 B.n604 B.n603 10.6151
R2831 B.n603 B.n600 10.6151
R2832 B.n600 B.n599 10.6151
R2833 B.n599 B.n596 10.6151
R2834 B.n596 B.n595 10.6151
R2835 B.n595 B.n592 10.6151
R2836 B.n592 B.n591 10.6151
R2837 B.n591 B.n588 10.6151
R2838 B.n588 B.n587 10.6151
R2839 B.n587 B.n584 10.6151
R2840 B.n584 B.n583 10.6151
R2841 B.n583 B.n581 10.6151
R2842 B.n826 B.n825 10.6151
R2843 B.n826 B.n506 10.6151
R2844 B.n836 B.n506 10.6151
R2845 B.n837 B.n836 10.6151
R2846 B.n838 B.n837 10.6151
R2847 B.n838 B.n498 10.6151
R2848 B.n848 B.n498 10.6151
R2849 B.n849 B.n848 10.6151
R2850 B.n850 B.n849 10.6151
R2851 B.n850 B.n490 10.6151
R2852 B.n860 B.n490 10.6151
R2853 B.n861 B.n860 10.6151
R2854 B.n862 B.n861 10.6151
R2855 B.n862 B.n482 10.6151
R2856 B.n872 B.n482 10.6151
R2857 B.n873 B.n872 10.6151
R2858 B.n874 B.n873 10.6151
R2859 B.n874 B.n474 10.6151
R2860 B.n884 B.n474 10.6151
R2861 B.n885 B.n884 10.6151
R2862 B.n886 B.n885 10.6151
R2863 B.n886 B.n466 10.6151
R2864 B.n897 B.n466 10.6151
R2865 B.n898 B.n897 10.6151
R2866 B.n899 B.n898 10.6151
R2867 B.n899 B.n459 10.6151
R2868 B.n909 B.n459 10.6151
R2869 B.n910 B.n909 10.6151
R2870 B.n911 B.n910 10.6151
R2871 B.n911 B.n451 10.6151
R2872 B.n921 B.n451 10.6151
R2873 B.n922 B.n921 10.6151
R2874 B.n923 B.n922 10.6151
R2875 B.n923 B.n443 10.6151
R2876 B.n933 B.n443 10.6151
R2877 B.n934 B.n933 10.6151
R2878 B.n935 B.n934 10.6151
R2879 B.n935 B.n435 10.6151
R2880 B.n945 B.n435 10.6151
R2881 B.n946 B.n945 10.6151
R2882 B.n947 B.n946 10.6151
R2883 B.n947 B.n427 10.6151
R2884 B.n957 B.n427 10.6151
R2885 B.n958 B.n957 10.6151
R2886 B.n959 B.n958 10.6151
R2887 B.n959 B.n419 10.6151
R2888 B.n969 B.n419 10.6151
R2889 B.n970 B.n969 10.6151
R2890 B.n971 B.n970 10.6151
R2891 B.n971 B.n411 10.6151
R2892 B.n982 B.n411 10.6151
R2893 B.n983 B.n982 10.6151
R2894 B.n984 B.n983 10.6151
R2895 B.n984 B.n0 10.6151
R2896 B.n1171 B.n1 10.6151
R2897 B.n1171 B.n1170 10.6151
R2898 B.n1170 B.n1169 10.6151
R2899 B.n1169 B.n10 10.6151
R2900 B.n1163 B.n10 10.6151
R2901 B.n1163 B.n1162 10.6151
R2902 B.n1162 B.n1161 10.6151
R2903 B.n1161 B.n17 10.6151
R2904 B.n1155 B.n17 10.6151
R2905 B.n1155 B.n1154 10.6151
R2906 B.n1154 B.n1153 10.6151
R2907 B.n1153 B.n24 10.6151
R2908 B.n1147 B.n24 10.6151
R2909 B.n1147 B.n1146 10.6151
R2910 B.n1146 B.n1145 10.6151
R2911 B.n1145 B.n31 10.6151
R2912 B.n1139 B.n31 10.6151
R2913 B.n1139 B.n1138 10.6151
R2914 B.n1138 B.n1137 10.6151
R2915 B.n1137 B.n38 10.6151
R2916 B.n1131 B.n38 10.6151
R2917 B.n1131 B.n1130 10.6151
R2918 B.n1130 B.n1129 10.6151
R2919 B.n1129 B.n45 10.6151
R2920 B.n1123 B.n45 10.6151
R2921 B.n1123 B.n1122 10.6151
R2922 B.n1122 B.n1121 10.6151
R2923 B.n1121 B.n52 10.6151
R2924 B.n1115 B.n52 10.6151
R2925 B.n1115 B.n1114 10.6151
R2926 B.n1114 B.n1113 10.6151
R2927 B.n1113 B.n58 10.6151
R2928 B.n1107 B.n58 10.6151
R2929 B.n1107 B.n1106 10.6151
R2930 B.n1106 B.n1105 10.6151
R2931 B.n1105 B.n66 10.6151
R2932 B.n1099 B.n66 10.6151
R2933 B.n1099 B.n1098 10.6151
R2934 B.n1098 B.n1097 10.6151
R2935 B.n1097 B.n73 10.6151
R2936 B.n1091 B.n73 10.6151
R2937 B.n1091 B.n1090 10.6151
R2938 B.n1090 B.n1089 10.6151
R2939 B.n1089 B.n80 10.6151
R2940 B.n1083 B.n80 10.6151
R2941 B.n1083 B.n1082 10.6151
R2942 B.n1082 B.n1081 10.6151
R2943 B.n1081 B.n87 10.6151
R2944 B.n1075 B.n87 10.6151
R2945 B.n1075 B.n1074 10.6151
R2946 B.n1074 B.n1073 10.6151
R2947 B.n1073 B.n94 10.6151
R2948 B.n1067 B.n94 10.6151
R2949 B.n1067 B.n1066 10.6151
R2950 B.n276 B.n169 9.36635
R2951 B.n299 B.n166 9.36635
R2952 B.n714 B.n713 9.36635
R2953 B.n692 B.n691 9.36635
R2954 B.t5 B.n441 6.92963
R2955 B.t1 B.n36 6.92963
R2956 B.n852 B.t7 3.96001
R2957 B.t11 B.n1085 3.96001
R2958 B.n1177 B.n0 2.81026
R2959 B.n1177 B.n1 2.81026
R2960 B.n894 B.t0 1.98025
R2961 B.n60 B.t2 1.98025
R2962 B.n279 B.n169 1.24928
R2963 B.n296 B.n166 1.24928
R2964 B.n713 B.n712 1.24928
R2965 B.n693 B.n692 1.24928
R2966 VN.n33 VN.n18 161.3
R2967 VN.n32 VN.n31 161.3
R2968 VN.n30 VN.n19 161.3
R2969 VN.n29 VN.n28 161.3
R2970 VN.n27 VN.n20 161.3
R2971 VN.n26 VN.n25 161.3
R2972 VN.n24 VN.n21 161.3
R2973 VN.n15 VN.n0 161.3
R2974 VN.n14 VN.n13 161.3
R2975 VN.n12 VN.n1 161.3
R2976 VN.n11 VN.n10 161.3
R2977 VN.n9 VN.n2 161.3
R2978 VN.n8 VN.n7 161.3
R2979 VN.n6 VN.n3 161.3
R2980 VN.n5 VN.t3 143.768
R2981 VN.n23 VN.t4 143.768
R2982 VN.n4 VN.t1 111.612
R2983 VN.n16 VN.t2 111.612
R2984 VN.n22 VN.t5 111.612
R2985 VN.n34 VN.t0 111.612
R2986 VN.n17 VN.n16 58.2041
R2987 VN.n35 VN.n34 58.2041
R2988 VN VN.n35 56.8413
R2989 VN.n5 VN.n4 50.4706
R2990 VN.n23 VN.n22 50.4706
R2991 VN.n10 VN.n9 40.979
R2992 VN.n28 VN.n27 40.979
R2993 VN.n10 VN.n1 40.0078
R2994 VN.n28 VN.n19 40.0078
R2995 VN.n4 VN.n3 24.4675
R2996 VN.n8 VN.n3 24.4675
R2997 VN.n9 VN.n8 24.4675
R2998 VN.n14 VN.n1 24.4675
R2999 VN.n15 VN.n14 24.4675
R3000 VN.n27 VN.n26 24.4675
R3001 VN.n26 VN.n21 24.4675
R3002 VN.n22 VN.n21 24.4675
R3003 VN.n33 VN.n32 24.4675
R3004 VN.n32 VN.n19 24.4675
R3005 VN.n16 VN.n15 23.9782
R3006 VN.n34 VN.n33 23.9782
R3007 VN.n24 VN.n23 2.54324
R3008 VN.n6 VN.n5 2.54324
R3009 VN.n35 VN.n18 0.417535
R3010 VN.n17 VN.n0 0.417535
R3011 VN VN.n17 0.394291
R3012 VN.n31 VN.n18 0.189894
R3013 VN.n31 VN.n30 0.189894
R3014 VN.n30 VN.n29 0.189894
R3015 VN.n29 VN.n20 0.189894
R3016 VN.n25 VN.n20 0.189894
R3017 VN.n25 VN.n24 0.189894
R3018 VN.n7 VN.n6 0.189894
R3019 VN.n7 VN.n2 0.189894
R3020 VN.n11 VN.n2 0.189894
R3021 VN.n12 VN.n11 0.189894
R3022 VN.n13 VN.n12 0.189894
R3023 VN.n13 VN.n0 0.189894
R3024 VDD2.n183 VDD2.n95 289.615
R3025 VDD2.n88 VDD2.n0 289.615
R3026 VDD2.n184 VDD2.n183 185
R3027 VDD2.n182 VDD2.n181 185
R3028 VDD2.n99 VDD2.n98 185
R3029 VDD2.n176 VDD2.n175 185
R3030 VDD2.n174 VDD2.n173 185
R3031 VDD2.n172 VDD2.n102 185
R3032 VDD2.n106 VDD2.n103 185
R3033 VDD2.n167 VDD2.n166 185
R3034 VDD2.n165 VDD2.n164 185
R3035 VDD2.n108 VDD2.n107 185
R3036 VDD2.n159 VDD2.n158 185
R3037 VDD2.n157 VDD2.n156 185
R3038 VDD2.n112 VDD2.n111 185
R3039 VDD2.n151 VDD2.n150 185
R3040 VDD2.n149 VDD2.n148 185
R3041 VDD2.n116 VDD2.n115 185
R3042 VDD2.n143 VDD2.n142 185
R3043 VDD2.n141 VDD2.n140 185
R3044 VDD2.n120 VDD2.n119 185
R3045 VDD2.n135 VDD2.n134 185
R3046 VDD2.n133 VDD2.n132 185
R3047 VDD2.n124 VDD2.n123 185
R3048 VDD2.n127 VDD2.n126 185
R3049 VDD2.n31 VDD2.n30 185
R3050 VDD2.n28 VDD2.n27 185
R3051 VDD2.n37 VDD2.n36 185
R3052 VDD2.n39 VDD2.n38 185
R3053 VDD2.n24 VDD2.n23 185
R3054 VDD2.n45 VDD2.n44 185
R3055 VDD2.n47 VDD2.n46 185
R3056 VDD2.n20 VDD2.n19 185
R3057 VDD2.n53 VDD2.n52 185
R3058 VDD2.n55 VDD2.n54 185
R3059 VDD2.n16 VDD2.n15 185
R3060 VDD2.n61 VDD2.n60 185
R3061 VDD2.n63 VDD2.n62 185
R3062 VDD2.n12 VDD2.n11 185
R3063 VDD2.n69 VDD2.n68 185
R3064 VDD2.n72 VDD2.n71 185
R3065 VDD2.n70 VDD2.n8 185
R3066 VDD2.n77 VDD2.n7 185
R3067 VDD2.n79 VDD2.n78 185
R3068 VDD2.n81 VDD2.n80 185
R3069 VDD2.n4 VDD2.n3 185
R3070 VDD2.n87 VDD2.n86 185
R3071 VDD2.n89 VDD2.n88 185
R3072 VDD2.t5 VDD2.n125 147.659
R3073 VDD2.t2 VDD2.n29 147.659
R3074 VDD2.n183 VDD2.n182 104.615
R3075 VDD2.n182 VDD2.n98 104.615
R3076 VDD2.n175 VDD2.n98 104.615
R3077 VDD2.n175 VDD2.n174 104.615
R3078 VDD2.n174 VDD2.n102 104.615
R3079 VDD2.n106 VDD2.n102 104.615
R3080 VDD2.n166 VDD2.n106 104.615
R3081 VDD2.n166 VDD2.n165 104.615
R3082 VDD2.n165 VDD2.n107 104.615
R3083 VDD2.n158 VDD2.n107 104.615
R3084 VDD2.n158 VDD2.n157 104.615
R3085 VDD2.n157 VDD2.n111 104.615
R3086 VDD2.n150 VDD2.n111 104.615
R3087 VDD2.n150 VDD2.n149 104.615
R3088 VDD2.n149 VDD2.n115 104.615
R3089 VDD2.n142 VDD2.n115 104.615
R3090 VDD2.n142 VDD2.n141 104.615
R3091 VDD2.n141 VDD2.n119 104.615
R3092 VDD2.n134 VDD2.n119 104.615
R3093 VDD2.n134 VDD2.n133 104.615
R3094 VDD2.n133 VDD2.n123 104.615
R3095 VDD2.n126 VDD2.n123 104.615
R3096 VDD2.n30 VDD2.n27 104.615
R3097 VDD2.n37 VDD2.n27 104.615
R3098 VDD2.n38 VDD2.n37 104.615
R3099 VDD2.n38 VDD2.n23 104.615
R3100 VDD2.n45 VDD2.n23 104.615
R3101 VDD2.n46 VDD2.n45 104.615
R3102 VDD2.n46 VDD2.n19 104.615
R3103 VDD2.n53 VDD2.n19 104.615
R3104 VDD2.n54 VDD2.n53 104.615
R3105 VDD2.n54 VDD2.n15 104.615
R3106 VDD2.n61 VDD2.n15 104.615
R3107 VDD2.n62 VDD2.n61 104.615
R3108 VDD2.n62 VDD2.n11 104.615
R3109 VDD2.n69 VDD2.n11 104.615
R3110 VDD2.n71 VDD2.n69 104.615
R3111 VDD2.n71 VDD2.n70 104.615
R3112 VDD2.n70 VDD2.n7 104.615
R3113 VDD2.n79 VDD2.n7 104.615
R3114 VDD2.n80 VDD2.n79 104.615
R3115 VDD2.n80 VDD2.n3 104.615
R3116 VDD2.n87 VDD2.n3 104.615
R3117 VDD2.n88 VDD2.n87 104.615
R3118 VDD2.n94 VDD2.n93 64.4383
R3119 VDD2 VDD2.n189 64.4355
R3120 VDD2.n94 VDD2.n92 54.2976
R3121 VDD2.n126 VDD2.t5 52.3082
R3122 VDD2.n30 VDD2.t2 52.3082
R3123 VDD2.n188 VDD2.n187 51.7732
R3124 VDD2.n188 VDD2.n94 49.5062
R3125 VDD2.n127 VDD2.n125 15.6677
R3126 VDD2.n31 VDD2.n29 15.6677
R3127 VDD2.n173 VDD2.n172 13.1884
R3128 VDD2.n78 VDD2.n77 13.1884
R3129 VDD2.n176 VDD2.n101 12.8005
R3130 VDD2.n171 VDD2.n103 12.8005
R3131 VDD2.n128 VDD2.n124 12.8005
R3132 VDD2.n32 VDD2.n28 12.8005
R3133 VDD2.n76 VDD2.n8 12.8005
R3134 VDD2.n81 VDD2.n6 12.8005
R3135 VDD2.n177 VDD2.n99 12.0247
R3136 VDD2.n168 VDD2.n167 12.0247
R3137 VDD2.n132 VDD2.n131 12.0247
R3138 VDD2.n36 VDD2.n35 12.0247
R3139 VDD2.n73 VDD2.n72 12.0247
R3140 VDD2.n82 VDD2.n4 12.0247
R3141 VDD2.n181 VDD2.n180 11.249
R3142 VDD2.n164 VDD2.n105 11.249
R3143 VDD2.n135 VDD2.n122 11.249
R3144 VDD2.n39 VDD2.n26 11.249
R3145 VDD2.n68 VDD2.n10 11.249
R3146 VDD2.n86 VDD2.n85 11.249
R3147 VDD2.n184 VDD2.n97 10.4732
R3148 VDD2.n163 VDD2.n108 10.4732
R3149 VDD2.n136 VDD2.n120 10.4732
R3150 VDD2.n40 VDD2.n24 10.4732
R3151 VDD2.n67 VDD2.n12 10.4732
R3152 VDD2.n89 VDD2.n2 10.4732
R3153 VDD2.n185 VDD2.n95 9.69747
R3154 VDD2.n160 VDD2.n159 9.69747
R3155 VDD2.n140 VDD2.n139 9.69747
R3156 VDD2.n44 VDD2.n43 9.69747
R3157 VDD2.n64 VDD2.n63 9.69747
R3158 VDD2.n90 VDD2.n0 9.69747
R3159 VDD2.n187 VDD2.n186 9.45567
R3160 VDD2.n92 VDD2.n91 9.45567
R3161 VDD2.n153 VDD2.n152 9.3005
R3162 VDD2.n155 VDD2.n154 9.3005
R3163 VDD2.n110 VDD2.n109 9.3005
R3164 VDD2.n161 VDD2.n160 9.3005
R3165 VDD2.n163 VDD2.n162 9.3005
R3166 VDD2.n105 VDD2.n104 9.3005
R3167 VDD2.n169 VDD2.n168 9.3005
R3168 VDD2.n171 VDD2.n170 9.3005
R3169 VDD2.n186 VDD2.n185 9.3005
R3170 VDD2.n97 VDD2.n96 9.3005
R3171 VDD2.n180 VDD2.n179 9.3005
R3172 VDD2.n178 VDD2.n177 9.3005
R3173 VDD2.n101 VDD2.n100 9.3005
R3174 VDD2.n114 VDD2.n113 9.3005
R3175 VDD2.n147 VDD2.n146 9.3005
R3176 VDD2.n145 VDD2.n144 9.3005
R3177 VDD2.n118 VDD2.n117 9.3005
R3178 VDD2.n139 VDD2.n138 9.3005
R3179 VDD2.n137 VDD2.n136 9.3005
R3180 VDD2.n122 VDD2.n121 9.3005
R3181 VDD2.n131 VDD2.n130 9.3005
R3182 VDD2.n129 VDD2.n128 9.3005
R3183 VDD2.n91 VDD2.n90 9.3005
R3184 VDD2.n2 VDD2.n1 9.3005
R3185 VDD2.n85 VDD2.n84 9.3005
R3186 VDD2.n83 VDD2.n82 9.3005
R3187 VDD2.n6 VDD2.n5 9.3005
R3188 VDD2.n51 VDD2.n50 9.3005
R3189 VDD2.n49 VDD2.n48 9.3005
R3190 VDD2.n22 VDD2.n21 9.3005
R3191 VDD2.n43 VDD2.n42 9.3005
R3192 VDD2.n41 VDD2.n40 9.3005
R3193 VDD2.n26 VDD2.n25 9.3005
R3194 VDD2.n35 VDD2.n34 9.3005
R3195 VDD2.n33 VDD2.n32 9.3005
R3196 VDD2.n18 VDD2.n17 9.3005
R3197 VDD2.n57 VDD2.n56 9.3005
R3198 VDD2.n59 VDD2.n58 9.3005
R3199 VDD2.n14 VDD2.n13 9.3005
R3200 VDD2.n65 VDD2.n64 9.3005
R3201 VDD2.n67 VDD2.n66 9.3005
R3202 VDD2.n10 VDD2.n9 9.3005
R3203 VDD2.n74 VDD2.n73 9.3005
R3204 VDD2.n76 VDD2.n75 9.3005
R3205 VDD2.n156 VDD2.n110 8.92171
R3206 VDD2.n143 VDD2.n118 8.92171
R3207 VDD2.n47 VDD2.n22 8.92171
R3208 VDD2.n60 VDD2.n14 8.92171
R3209 VDD2.n155 VDD2.n112 8.14595
R3210 VDD2.n144 VDD2.n116 8.14595
R3211 VDD2.n48 VDD2.n20 8.14595
R3212 VDD2.n59 VDD2.n16 8.14595
R3213 VDD2.n152 VDD2.n151 7.3702
R3214 VDD2.n148 VDD2.n147 7.3702
R3215 VDD2.n52 VDD2.n51 7.3702
R3216 VDD2.n56 VDD2.n55 7.3702
R3217 VDD2.n151 VDD2.n114 6.59444
R3218 VDD2.n148 VDD2.n114 6.59444
R3219 VDD2.n52 VDD2.n18 6.59444
R3220 VDD2.n55 VDD2.n18 6.59444
R3221 VDD2.n152 VDD2.n112 5.81868
R3222 VDD2.n147 VDD2.n116 5.81868
R3223 VDD2.n51 VDD2.n20 5.81868
R3224 VDD2.n56 VDD2.n16 5.81868
R3225 VDD2.n156 VDD2.n155 5.04292
R3226 VDD2.n144 VDD2.n143 5.04292
R3227 VDD2.n48 VDD2.n47 5.04292
R3228 VDD2.n60 VDD2.n59 5.04292
R3229 VDD2.n129 VDD2.n125 4.38563
R3230 VDD2.n33 VDD2.n29 4.38563
R3231 VDD2.n187 VDD2.n95 4.26717
R3232 VDD2.n159 VDD2.n110 4.26717
R3233 VDD2.n140 VDD2.n118 4.26717
R3234 VDD2.n44 VDD2.n22 4.26717
R3235 VDD2.n63 VDD2.n14 4.26717
R3236 VDD2.n92 VDD2.n0 4.26717
R3237 VDD2.n185 VDD2.n184 3.49141
R3238 VDD2.n160 VDD2.n108 3.49141
R3239 VDD2.n139 VDD2.n120 3.49141
R3240 VDD2.n43 VDD2.n24 3.49141
R3241 VDD2.n64 VDD2.n12 3.49141
R3242 VDD2.n90 VDD2.n89 3.49141
R3243 VDD2.n181 VDD2.n97 2.71565
R3244 VDD2.n164 VDD2.n163 2.71565
R3245 VDD2.n136 VDD2.n135 2.71565
R3246 VDD2.n40 VDD2.n39 2.71565
R3247 VDD2.n68 VDD2.n67 2.71565
R3248 VDD2.n86 VDD2.n2 2.71565
R3249 VDD2 VDD2.n188 2.63843
R3250 VDD2.n180 VDD2.n99 1.93989
R3251 VDD2.n167 VDD2.n105 1.93989
R3252 VDD2.n132 VDD2.n122 1.93989
R3253 VDD2.n36 VDD2.n26 1.93989
R3254 VDD2.n72 VDD2.n10 1.93989
R3255 VDD2.n85 VDD2.n4 1.93989
R3256 VDD2.n189 VDD2.t0 1.16864
R3257 VDD2.n189 VDD2.t1 1.16864
R3258 VDD2.n93 VDD2.t4 1.16864
R3259 VDD2.n93 VDD2.t3 1.16864
R3260 VDD2.n177 VDD2.n176 1.16414
R3261 VDD2.n168 VDD2.n103 1.16414
R3262 VDD2.n131 VDD2.n124 1.16414
R3263 VDD2.n35 VDD2.n28 1.16414
R3264 VDD2.n73 VDD2.n8 1.16414
R3265 VDD2.n82 VDD2.n81 1.16414
R3266 VDD2.n173 VDD2.n101 0.388379
R3267 VDD2.n172 VDD2.n171 0.388379
R3268 VDD2.n128 VDD2.n127 0.388379
R3269 VDD2.n32 VDD2.n31 0.388379
R3270 VDD2.n77 VDD2.n76 0.388379
R3271 VDD2.n78 VDD2.n6 0.388379
R3272 VDD2.n186 VDD2.n96 0.155672
R3273 VDD2.n179 VDD2.n96 0.155672
R3274 VDD2.n179 VDD2.n178 0.155672
R3275 VDD2.n178 VDD2.n100 0.155672
R3276 VDD2.n170 VDD2.n100 0.155672
R3277 VDD2.n170 VDD2.n169 0.155672
R3278 VDD2.n169 VDD2.n104 0.155672
R3279 VDD2.n162 VDD2.n104 0.155672
R3280 VDD2.n162 VDD2.n161 0.155672
R3281 VDD2.n161 VDD2.n109 0.155672
R3282 VDD2.n154 VDD2.n109 0.155672
R3283 VDD2.n154 VDD2.n153 0.155672
R3284 VDD2.n153 VDD2.n113 0.155672
R3285 VDD2.n146 VDD2.n113 0.155672
R3286 VDD2.n146 VDD2.n145 0.155672
R3287 VDD2.n145 VDD2.n117 0.155672
R3288 VDD2.n138 VDD2.n117 0.155672
R3289 VDD2.n138 VDD2.n137 0.155672
R3290 VDD2.n137 VDD2.n121 0.155672
R3291 VDD2.n130 VDD2.n121 0.155672
R3292 VDD2.n130 VDD2.n129 0.155672
R3293 VDD2.n34 VDD2.n33 0.155672
R3294 VDD2.n34 VDD2.n25 0.155672
R3295 VDD2.n41 VDD2.n25 0.155672
R3296 VDD2.n42 VDD2.n41 0.155672
R3297 VDD2.n42 VDD2.n21 0.155672
R3298 VDD2.n49 VDD2.n21 0.155672
R3299 VDD2.n50 VDD2.n49 0.155672
R3300 VDD2.n50 VDD2.n17 0.155672
R3301 VDD2.n57 VDD2.n17 0.155672
R3302 VDD2.n58 VDD2.n57 0.155672
R3303 VDD2.n58 VDD2.n13 0.155672
R3304 VDD2.n65 VDD2.n13 0.155672
R3305 VDD2.n66 VDD2.n65 0.155672
R3306 VDD2.n66 VDD2.n9 0.155672
R3307 VDD2.n74 VDD2.n9 0.155672
R3308 VDD2.n75 VDD2.n74 0.155672
R3309 VDD2.n75 VDD2.n5 0.155672
R3310 VDD2.n83 VDD2.n5 0.155672
R3311 VDD2.n84 VDD2.n83 0.155672
R3312 VDD2.n84 VDD2.n1 0.155672
R3313 VDD2.n91 VDD2.n1 0.155672
C0 VDD1 VDD2 1.81963f
C1 VDD2 VP 0.54802f
C2 VDD2 VN 9.88356f
C3 VTAIL VDD1 9.68811f
C4 VTAIL VP 10.076599f
C5 VTAIL VN 10.062099f
C6 VDD1 VP 10.2762f
C7 VDD1 VN 0.151993f
C8 VP VN 8.878961f
C9 VTAIL VDD2 9.74613f
C10 VDD2 B 7.66148f
C11 VDD1 B 7.848125f
C12 VTAIL B 10.504504f
C13 VN B 16.423971f
C14 VP B 15.084857f
C15 VDD2.n0 B 0.030678f
C16 VDD2.n1 B 0.021116f
C17 VDD2.n2 B 0.011347f
C18 VDD2.n3 B 0.02682f
C19 VDD2.n4 B 0.012014f
C20 VDD2.n5 B 0.021116f
C21 VDD2.n6 B 0.011347f
C22 VDD2.n7 B 0.02682f
C23 VDD2.n8 B 0.012014f
C24 VDD2.n9 B 0.021116f
C25 VDD2.n10 B 0.011347f
C26 VDD2.n11 B 0.02682f
C27 VDD2.n12 B 0.012014f
C28 VDD2.n13 B 0.021116f
C29 VDD2.n14 B 0.011347f
C30 VDD2.n15 B 0.02682f
C31 VDD2.n16 B 0.012014f
C32 VDD2.n17 B 0.021116f
C33 VDD2.n18 B 0.011347f
C34 VDD2.n19 B 0.02682f
C35 VDD2.n20 B 0.012014f
C36 VDD2.n21 B 0.021116f
C37 VDD2.n22 B 0.011347f
C38 VDD2.n23 B 0.02682f
C39 VDD2.n24 B 0.012014f
C40 VDD2.n25 B 0.021116f
C41 VDD2.n26 B 0.011347f
C42 VDD2.n27 B 0.02682f
C43 VDD2.n28 B 0.012014f
C44 VDD2.n29 B 0.148047f
C45 VDD2.t2 B 0.044364f
C46 VDD2.n30 B 0.020115f
C47 VDD2.n31 B 0.015843f
C48 VDD2.n32 B 0.011347f
C49 VDD2.n33 B 1.56255f
C50 VDD2.n34 B 0.021116f
C51 VDD2.n35 B 0.011347f
C52 VDD2.n36 B 0.012014f
C53 VDD2.n37 B 0.02682f
C54 VDD2.n38 B 0.02682f
C55 VDD2.n39 B 0.012014f
C56 VDD2.n40 B 0.011347f
C57 VDD2.n41 B 0.021116f
C58 VDD2.n42 B 0.021116f
C59 VDD2.n43 B 0.011347f
C60 VDD2.n44 B 0.012014f
C61 VDD2.n45 B 0.02682f
C62 VDD2.n46 B 0.02682f
C63 VDD2.n47 B 0.012014f
C64 VDD2.n48 B 0.011347f
C65 VDD2.n49 B 0.021116f
C66 VDD2.n50 B 0.021116f
C67 VDD2.n51 B 0.011347f
C68 VDD2.n52 B 0.012014f
C69 VDD2.n53 B 0.02682f
C70 VDD2.n54 B 0.02682f
C71 VDD2.n55 B 0.012014f
C72 VDD2.n56 B 0.011347f
C73 VDD2.n57 B 0.021116f
C74 VDD2.n58 B 0.021116f
C75 VDD2.n59 B 0.011347f
C76 VDD2.n60 B 0.012014f
C77 VDD2.n61 B 0.02682f
C78 VDD2.n62 B 0.02682f
C79 VDD2.n63 B 0.012014f
C80 VDD2.n64 B 0.011347f
C81 VDD2.n65 B 0.021116f
C82 VDD2.n66 B 0.021116f
C83 VDD2.n67 B 0.011347f
C84 VDD2.n68 B 0.012014f
C85 VDD2.n69 B 0.02682f
C86 VDD2.n70 B 0.02682f
C87 VDD2.n71 B 0.02682f
C88 VDD2.n72 B 0.012014f
C89 VDD2.n73 B 0.011347f
C90 VDD2.n74 B 0.021116f
C91 VDD2.n75 B 0.021116f
C92 VDD2.n76 B 0.011347f
C93 VDD2.n77 B 0.011681f
C94 VDD2.n78 B 0.011681f
C95 VDD2.n79 B 0.02682f
C96 VDD2.n80 B 0.02682f
C97 VDD2.n81 B 0.012014f
C98 VDD2.n82 B 0.011347f
C99 VDD2.n83 B 0.021116f
C100 VDD2.n84 B 0.021116f
C101 VDD2.n85 B 0.011347f
C102 VDD2.n86 B 0.012014f
C103 VDD2.n87 B 0.02682f
C104 VDD2.n88 B 0.059824f
C105 VDD2.n89 B 0.012014f
C106 VDD2.n90 B 0.011347f
C107 VDD2.n91 B 0.053136f
C108 VDD2.n92 B 0.058333f
C109 VDD2.t4 B 0.282837f
C110 VDD2.t3 B 0.282837f
C111 VDD2.n93 B 2.5789f
C112 VDD2.n94 B 2.91107f
C113 VDD2.n95 B 0.030678f
C114 VDD2.n96 B 0.021116f
C115 VDD2.n97 B 0.011347f
C116 VDD2.n98 B 0.02682f
C117 VDD2.n99 B 0.012014f
C118 VDD2.n100 B 0.021116f
C119 VDD2.n101 B 0.011347f
C120 VDD2.n102 B 0.02682f
C121 VDD2.n103 B 0.012014f
C122 VDD2.n104 B 0.021116f
C123 VDD2.n105 B 0.011347f
C124 VDD2.n106 B 0.02682f
C125 VDD2.n107 B 0.02682f
C126 VDD2.n108 B 0.012014f
C127 VDD2.n109 B 0.021116f
C128 VDD2.n110 B 0.011347f
C129 VDD2.n111 B 0.02682f
C130 VDD2.n112 B 0.012014f
C131 VDD2.n113 B 0.021116f
C132 VDD2.n114 B 0.011347f
C133 VDD2.n115 B 0.02682f
C134 VDD2.n116 B 0.012014f
C135 VDD2.n117 B 0.021116f
C136 VDD2.n118 B 0.011347f
C137 VDD2.n119 B 0.02682f
C138 VDD2.n120 B 0.012014f
C139 VDD2.n121 B 0.021116f
C140 VDD2.n122 B 0.011347f
C141 VDD2.n123 B 0.02682f
C142 VDD2.n124 B 0.012014f
C143 VDD2.n125 B 0.148047f
C144 VDD2.t5 B 0.044364f
C145 VDD2.n126 B 0.020115f
C146 VDD2.n127 B 0.015843f
C147 VDD2.n128 B 0.011347f
C148 VDD2.n129 B 1.56255f
C149 VDD2.n130 B 0.021116f
C150 VDD2.n131 B 0.011347f
C151 VDD2.n132 B 0.012014f
C152 VDD2.n133 B 0.02682f
C153 VDD2.n134 B 0.02682f
C154 VDD2.n135 B 0.012014f
C155 VDD2.n136 B 0.011347f
C156 VDD2.n137 B 0.021116f
C157 VDD2.n138 B 0.021116f
C158 VDD2.n139 B 0.011347f
C159 VDD2.n140 B 0.012014f
C160 VDD2.n141 B 0.02682f
C161 VDD2.n142 B 0.02682f
C162 VDD2.n143 B 0.012014f
C163 VDD2.n144 B 0.011347f
C164 VDD2.n145 B 0.021116f
C165 VDD2.n146 B 0.021116f
C166 VDD2.n147 B 0.011347f
C167 VDD2.n148 B 0.012014f
C168 VDD2.n149 B 0.02682f
C169 VDD2.n150 B 0.02682f
C170 VDD2.n151 B 0.012014f
C171 VDD2.n152 B 0.011347f
C172 VDD2.n153 B 0.021116f
C173 VDD2.n154 B 0.021116f
C174 VDD2.n155 B 0.011347f
C175 VDD2.n156 B 0.012014f
C176 VDD2.n157 B 0.02682f
C177 VDD2.n158 B 0.02682f
C178 VDD2.n159 B 0.012014f
C179 VDD2.n160 B 0.011347f
C180 VDD2.n161 B 0.021116f
C181 VDD2.n162 B 0.021116f
C182 VDD2.n163 B 0.011347f
C183 VDD2.n164 B 0.012014f
C184 VDD2.n165 B 0.02682f
C185 VDD2.n166 B 0.02682f
C186 VDD2.n167 B 0.012014f
C187 VDD2.n168 B 0.011347f
C188 VDD2.n169 B 0.021116f
C189 VDD2.n170 B 0.021116f
C190 VDD2.n171 B 0.011347f
C191 VDD2.n172 B 0.011681f
C192 VDD2.n173 B 0.011681f
C193 VDD2.n174 B 0.02682f
C194 VDD2.n175 B 0.02682f
C195 VDD2.n176 B 0.012014f
C196 VDD2.n177 B 0.011347f
C197 VDD2.n178 B 0.021116f
C198 VDD2.n179 B 0.021116f
C199 VDD2.n180 B 0.011347f
C200 VDD2.n181 B 0.012014f
C201 VDD2.n182 B 0.02682f
C202 VDD2.n183 B 0.059824f
C203 VDD2.n184 B 0.012014f
C204 VDD2.n185 B 0.011347f
C205 VDD2.n186 B 0.053136f
C206 VDD2.n187 B 0.048332f
C207 VDD2.n188 B 2.72917f
C208 VDD2.t0 B 0.282837f
C209 VDD2.t1 B 0.282837f
C210 VDD2.n189 B 2.57887f
C211 VN.n0 B 0.033374f
C212 VN.t2 B 3.02406f
C213 VN.n1 B 0.035351f
C214 VN.n2 B 0.017743f
C215 VN.n3 B 0.033068f
C216 VN.t3 B 3.28858f
C217 VN.t1 B 3.02406f
C218 VN.n4 B 1.11691f
C219 VN.n5 B 1.06799f
C220 VN.n6 B 0.22631f
C221 VN.n7 B 0.017743f
C222 VN.n8 B 0.033068f
C223 VN.n9 B 0.035173f
C224 VN.n10 B 0.01435f
C225 VN.n11 B 0.017743f
C226 VN.n12 B 0.017743f
C227 VN.n13 B 0.017743f
C228 VN.n14 B 0.033068f
C229 VN.n15 B 0.032742f
C230 VN.n16 B 1.12237f
C231 VN.n17 B 0.050385f
C232 VN.n18 B 0.033374f
C233 VN.t0 B 3.02406f
C234 VN.n19 B 0.035351f
C235 VN.n20 B 0.017743f
C236 VN.n21 B 0.033068f
C237 VN.t4 B 3.28858f
C238 VN.t5 B 3.02406f
C239 VN.n22 B 1.11691f
C240 VN.n23 B 1.06799f
C241 VN.n24 B 0.22631f
C242 VN.n25 B 0.017743f
C243 VN.n26 B 0.033068f
C244 VN.n27 B 0.035173f
C245 VN.n28 B 0.01435f
C246 VN.n29 B 0.017743f
C247 VN.n30 B 0.017743f
C248 VN.n31 B 0.017743f
C249 VN.n32 B 0.033068f
C250 VN.n33 B 0.032742f
C251 VN.n34 B 1.12237f
C252 VN.n35 B 1.22694f
C253 VDD1.n0 B 0.03118f
C254 VDD1.n1 B 0.021462f
C255 VDD1.n2 B 0.011533f
C256 VDD1.n3 B 0.027259f
C257 VDD1.n4 B 0.012211f
C258 VDD1.n5 B 0.021462f
C259 VDD1.n6 B 0.011533f
C260 VDD1.n7 B 0.027259f
C261 VDD1.n8 B 0.012211f
C262 VDD1.n9 B 0.021462f
C263 VDD1.n10 B 0.011533f
C264 VDD1.n11 B 0.027259f
C265 VDD1.n12 B 0.027259f
C266 VDD1.n13 B 0.012211f
C267 VDD1.n14 B 0.021462f
C268 VDD1.n15 B 0.011533f
C269 VDD1.n16 B 0.027259f
C270 VDD1.n17 B 0.012211f
C271 VDD1.n18 B 0.021462f
C272 VDD1.n19 B 0.011533f
C273 VDD1.n20 B 0.027259f
C274 VDD1.n21 B 0.012211f
C275 VDD1.n22 B 0.021462f
C276 VDD1.n23 B 0.011533f
C277 VDD1.n24 B 0.027259f
C278 VDD1.n25 B 0.012211f
C279 VDD1.n26 B 0.021462f
C280 VDD1.n27 B 0.011533f
C281 VDD1.n28 B 0.027259f
C282 VDD1.n29 B 0.012211f
C283 VDD1.n30 B 0.15047f
C284 VDD1.t5 B 0.04509f
C285 VDD1.n31 B 0.020444f
C286 VDD1.n32 B 0.016103f
C287 VDD1.n33 B 0.011533f
C288 VDD1.n34 B 1.58812f
C289 VDD1.n35 B 0.021462f
C290 VDD1.n36 B 0.011533f
C291 VDD1.n37 B 0.012211f
C292 VDD1.n38 B 0.027259f
C293 VDD1.n39 B 0.027259f
C294 VDD1.n40 B 0.012211f
C295 VDD1.n41 B 0.011533f
C296 VDD1.n42 B 0.021462f
C297 VDD1.n43 B 0.021462f
C298 VDD1.n44 B 0.011533f
C299 VDD1.n45 B 0.012211f
C300 VDD1.n46 B 0.027259f
C301 VDD1.n47 B 0.027259f
C302 VDD1.n48 B 0.012211f
C303 VDD1.n49 B 0.011533f
C304 VDD1.n50 B 0.021462f
C305 VDD1.n51 B 0.021462f
C306 VDD1.n52 B 0.011533f
C307 VDD1.n53 B 0.012211f
C308 VDD1.n54 B 0.027259f
C309 VDD1.n55 B 0.027259f
C310 VDD1.n56 B 0.012211f
C311 VDD1.n57 B 0.011533f
C312 VDD1.n58 B 0.021462f
C313 VDD1.n59 B 0.021462f
C314 VDD1.n60 B 0.011533f
C315 VDD1.n61 B 0.012211f
C316 VDD1.n62 B 0.027259f
C317 VDD1.n63 B 0.027259f
C318 VDD1.n64 B 0.012211f
C319 VDD1.n65 B 0.011533f
C320 VDD1.n66 B 0.021462f
C321 VDD1.n67 B 0.021462f
C322 VDD1.n68 B 0.011533f
C323 VDD1.n69 B 0.012211f
C324 VDD1.n70 B 0.027259f
C325 VDD1.n71 B 0.027259f
C326 VDD1.n72 B 0.012211f
C327 VDD1.n73 B 0.011533f
C328 VDD1.n74 B 0.021462f
C329 VDD1.n75 B 0.021462f
C330 VDD1.n76 B 0.011533f
C331 VDD1.n77 B 0.011872f
C332 VDD1.n78 B 0.011872f
C333 VDD1.n79 B 0.027259f
C334 VDD1.n80 B 0.027259f
C335 VDD1.n81 B 0.012211f
C336 VDD1.n82 B 0.011533f
C337 VDD1.n83 B 0.021462f
C338 VDD1.n84 B 0.021462f
C339 VDD1.n85 B 0.011533f
C340 VDD1.n86 B 0.012211f
C341 VDD1.n87 B 0.027259f
C342 VDD1.n88 B 0.060803f
C343 VDD1.n89 B 0.012211f
C344 VDD1.n90 B 0.011533f
C345 VDD1.n91 B 0.054005f
C346 VDD1.n92 B 0.060093f
C347 VDD1.n93 B 0.03118f
C348 VDD1.n94 B 0.021462f
C349 VDD1.n95 B 0.011533f
C350 VDD1.n96 B 0.027259f
C351 VDD1.n97 B 0.012211f
C352 VDD1.n98 B 0.021462f
C353 VDD1.n99 B 0.011533f
C354 VDD1.n100 B 0.027259f
C355 VDD1.n101 B 0.012211f
C356 VDD1.n102 B 0.021462f
C357 VDD1.n103 B 0.011533f
C358 VDD1.n104 B 0.027259f
C359 VDD1.n105 B 0.012211f
C360 VDD1.n106 B 0.021462f
C361 VDD1.n107 B 0.011533f
C362 VDD1.n108 B 0.027259f
C363 VDD1.n109 B 0.012211f
C364 VDD1.n110 B 0.021462f
C365 VDD1.n111 B 0.011533f
C366 VDD1.n112 B 0.027259f
C367 VDD1.n113 B 0.012211f
C368 VDD1.n114 B 0.021462f
C369 VDD1.n115 B 0.011533f
C370 VDD1.n116 B 0.027259f
C371 VDD1.n117 B 0.012211f
C372 VDD1.n118 B 0.021462f
C373 VDD1.n119 B 0.011533f
C374 VDD1.n120 B 0.027259f
C375 VDD1.n121 B 0.012211f
C376 VDD1.n122 B 0.15047f
C377 VDD1.t0 B 0.04509f
C378 VDD1.n123 B 0.020444f
C379 VDD1.n124 B 0.016103f
C380 VDD1.n125 B 0.011533f
C381 VDD1.n126 B 1.58812f
C382 VDD1.n127 B 0.021462f
C383 VDD1.n128 B 0.011533f
C384 VDD1.n129 B 0.012211f
C385 VDD1.n130 B 0.027259f
C386 VDD1.n131 B 0.027259f
C387 VDD1.n132 B 0.012211f
C388 VDD1.n133 B 0.011533f
C389 VDD1.n134 B 0.021462f
C390 VDD1.n135 B 0.021462f
C391 VDD1.n136 B 0.011533f
C392 VDD1.n137 B 0.012211f
C393 VDD1.n138 B 0.027259f
C394 VDD1.n139 B 0.027259f
C395 VDD1.n140 B 0.012211f
C396 VDD1.n141 B 0.011533f
C397 VDD1.n142 B 0.021462f
C398 VDD1.n143 B 0.021462f
C399 VDD1.n144 B 0.011533f
C400 VDD1.n145 B 0.012211f
C401 VDD1.n146 B 0.027259f
C402 VDD1.n147 B 0.027259f
C403 VDD1.n148 B 0.012211f
C404 VDD1.n149 B 0.011533f
C405 VDD1.n150 B 0.021462f
C406 VDD1.n151 B 0.021462f
C407 VDD1.n152 B 0.011533f
C408 VDD1.n153 B 0.012211f
C409 VDD1.n154 B 0.027259f
C410 VDD1.n155 B 0.027259f
C411 VDD1.n156 B 0.012211f
C412 VDD1.n157 B 0.011533f
C413 VDD1.n158 B 0.021462f
C414 VDD1.n159 B 0.021462f
C415 VDD1.n160 B 0.011533f
C416 VDD1.n161 B 0.012211f
C417 VDD1.n162 B 0.027259f
C418 VDD1.n163 B 0.027259f
C419 VDD1.n164 B 0.027259f
C420 VDD1.n165 B 0.012211f
C421 VDD1.n166 B 0.011533f
C422 VDD1.n167 B 0.021462f
C423 VDD1.n168 B 0.021462f
C424 VDD1.n169 B 0.011533f
C425 VDD1.n170 B 0.011872f
C426 VDD1.n171 B 0.011872f
C427 VDD1.n172 B 0.027259f
C428 VDD1.n173 B 0.027259f
C429 VDD1.n174 B 0.012211f
C430 VDD1.n175 B 0.011533f
C431 VDD1.n176 B 0.021462f
C432 VDD1.n177 B 0.021462f
C433 VDD1.n178 B 0.011533f
C434 VDD1.n179 B 0.012211f
C435 VDD1.n180 B 0.027259f
C436 VDD1.n181 B 0.060803f
C437 VDD1.n182 B 0.012211f
C438 VDD1.n183 B 0.011533f
C439 VDD1.n184 B 0.054005f
C440 VDD1.n185 B 0.059287f
C441 VDD1.t4 B 0.287465f
C442 VDD1.t3 B 0.287465f
C443 VDD1.n186 B 2.6211f
C444 VDD1.n187 B 3.09301f
C445 VDD1.t2 B 0.287465f
C446 VDD1.t1 B 0.287465f
C447 VDD1.n188 B 2.61514f
C448 VDD1.n189 B 2.96923f
C449 VTAIL.t3 B 0.310474f
C450 VTAIL.t1 B 0.310474f
C451 VTAIL.n0 B 2.75898f
C452 VTAIL.n1 B 0.454823f
C453 VTAIL.n2 B 0.033675f
C454 VTAIL.n3 B 0.023179f
C455 VTAIL.n4 B 0.012456f
C456 VTAIL.n5 B 0.02944f
C457 VTAIL.n6 B 0.013188f
C458 VTAIL.n7 B 0.023179f
C459 VTAIL.n8 B 0.012456f
C460 VTAIL.n9 B 0.02944f
C461 VTAIL.n10 B 0.013188f
C462 VTAIL.n11 B 0.023179f
C463 VTAIL.n12 B 0.012456f
C464 VTAIL.n13 B 0.02944f
C465 VTAIL.n14 B 0.013188f
C466 VTAIL.n15 B 0.023179f
C467 VTAIL.n16 B 0.012456f
C468 VTAIL.n17 B 0.02944f
C469 VTAIL.n18 B 0.013188f
C470 VTAIL.n19 B 0.023179f
C471 VTAIL.n20 B 0.012456f
C472 VTAIL.n21 B 0.02944f
C473 VTAIL.n22 B 0.013188f
C474 VTAIL.n23 B 0.023179f
C475 VTAIL.n24 B 0.012456f
C476 VTAIL.n25 B 0.02944f
C477 VTAIL.n26 B 0.013188f
C478 VTAIL.n27 B 0.023179f
C479 VTAIL.n28 B 0.012456f
C480 VTAIL.n29 B 0.02944f
C481 VTAIL.n30 B 0.013188f
C482 VTAIL.n31 B 0.162514f
C483 VTAIL.t6 B 0.048699f
C484 VTAIL.n32 B 0.02208f
C485 VTAIL.n33 B 0.017391f
C486 VTAIL.n34 B 0.012456f
C487 VTAIL.n35 B 1.71524f
C488 VTAIL.n36 B 0.023179f
C489 VTAIL.n37 B 0.012456f
C490 VTAIL.n38 B 0.013188f
C491 VTAIL.n39 B 0.02944f
C492 VTAIL.n40 B 0.02944f
C493 VTAIL.n41 B 0.013188f
C494 VTAIL.n42 B 0.012456f
C495 VTAIL.n43 B 0.023179f
C496 VTAIL.n44 B 0.023179f
C497 VTAIL.n45 B 0.012456f
C498 VTAIL.n46 B 0.013188f
C499 VTAIL.n47 B 0.02944f
C500 VTAIL.n48 B 0.02944f
C501 VTAIL.n49 B 0.013188f
C502 VTAIL.n50 B 0.012456f
C503 VTAIL.n51 B 0.023179f
C504 VTAIL.n52 B 0.023179f
C505 VTAIL.n53 B 0.012456f
C506 VTAIL.n54 B 0.013188f
C507 VTAIL.n55 B 0.02944f
C508 VTAIL.n56 B 0.02944f
C509 VTAIL.n57 B 0.013188f
C510 VTAIL.n58 B 0.012456f
C511 VTAIL.n59 B 0.023179f
C512 VTAIL.n60 B 0.023179f
C513 VTAIL.n61 B 0.012456f
C514 VTAIL.n62 B 0.013188f
C515 VTAIL.n63 B 0.02944f
C516 VTAIL.n64 B 0.02944f
C517 VTAIL.n65 B 0.013188f
C518 VTAIL.n66 B 0.012456f
C519 VTAIL.n67 B 0.023179f
C520 VTAIL.n68 B 0.023179f
C521 VTAIL.n69 B 0.012456f
C522 VTAIL.n70 B 0.013188f
C523 VTAIL.n71 B 0.02944f
C524 VTAIL.n72 B 0.02944f
C525 VTAIL.n73 B 0.02944f
C526 VTAIL.n74 B 0.013188f
C527 VTAIL.n75 B 0.012456f
C528 VTAIL.n76 B 0.023179f
C529 VTAIL.n77 B 0.023179f
C530 VTAIL.n78 B 0.012456f
C531 VTAIL.n79 B 0.012822f
C532 VTAIL.n80 B 0.012822f
C533 VTAIL.n81 B 0.02944f
C534 VTAIL.n82 B 0.02944f
C535 VTAIL.n83 B 0.013188f
C536 VTAIL.n84 B 0.012456f
C537 VTAIL.n85 B 0.023179f
C538 VTAIL.n86 B 0.023179f
C539 VTAIL.n87 B 0.012456f
C540 VTAIL.n88 B 0.013188f
C541 VTAIL.n89 B 0.02944f
C542 VTAIL.n90 B 0.06567f
C543 VTAIL.n91 B 0.013188f
C544 VTAIL.n92 B 0.012456f
C545 VTAIL.n93 B 0.058328f
C546 VTAIL.n94 B 0.037084f
C547 VTAIL.n95 B 0.442932f
C548 VTAIL.t9 B 0.310474f
C549 VTAIL.t7 B 0.310474f
C550 VTAIL.n96 B 2.75898f
C551 VTAIL.n97 B 2.39965f
C552 VTAIL.t0 B 0.310474f
C553 VTAIL.t5 B 0.310474f
C554 VTAIL.n98 B 2.75899f
C555 VTAIL.n99 B 2.39964f
C556 VTAIL.n100 B 0.033675f
C557 VTAIL.n101 B 0.023179f
C558 VTAIL.n102 B 0.012456f
C559 VTAIL.n103 B 0.02944f
C560 VTAIL.n104 B 0.013188f
C561 VTAIL.n105 B 0.023179f
C562 VTAIL.n106 B 0.012456f
C563 VTAIL.n107 B 0.02944f
C564 VTAIL.n108 B 0.013188f
C565 VTAIL.n109 B 0.023179f
C566 VTAIL.n110 B 0.012456f
C567 VTAIL.n111 B 0.02944f
C568 VTAIL.n112 B 0.02944f
C569 VTAIL.n113 B 0.013188f
C570 VTAIL.n114 B 0.023179f
C571 VTAIL.n115 B 0.012456f
C572 VTAIL.n116 B 0.02944f
C573 VTAIL.n117 B 0.013188f
C574 VTAIL.n118 B 0.023179f
C575 VTAIL.n119 B 0.012456f
C576 VTAIL.n120 B 0.02944f
C577 VTAIL.n121 B 0.013188f
C578 VTAIL.n122 B 0.023179f
C579 VTAIL.n123 B 0.012456f
C580 VTAIL.n124 B 0.02944f
C581 VTAIL.n125 B 0.013188f
C582 VTAIL.n126 B 0.023179f
C583 VTAIL.n127 B 0.012456f
C584 VTAIL.n128 B 0.02944f
C585 VTAIL.n129 B 0.013188f
C586 VTAIL.n130 B 0.162514f
C587 VTAIL.t4 B 0.048699f
C588 VTAIL.n131 B 0.02208f
C589 VTAIL.n132 B 0.017391f
C590 VTAIL.n133 B 0.012456f
C591 VTAIL.n134 B 1.71524f
C592 VTAIL.n135 B 0.023179f
C593 VTAIL.n136 B 0.012456f
C594 VTAIL.n137 B 0.013188f
C595 VTAIL.n138 B 0.02944f
C596 VTAIL.n139 B 0.02944f
C597 VTAIL.n140 B 0.013188f
C598 VTAIL.n141 B 0.012456f
C599 VTAIL.n142 B 0.023179f
C600 VTAIL.n143 B 0.023179f
C601 VTAIL.n144 B 0.012456f
C602 VTAIL.n145 B 0.013188f
C603 VTAIL.n146 B 0.02944f
C604 VTAIL.n147 B 0.02944f
C605 VTAIL.n148 B 0.013188f
C606 VTAIL.n149 B 0.012456f
C607 VTAIL.n150 B 0.023179f
C608 VTAIL.n151 B 0.023179f
C609 VTAIL.n152 B 0.012456f
C610 VTAIL.n153 B 0.013188f
C611 VTAIL.n154 B 0.02944f
C612 VTAIL.n155 B 0.02944f
C613 VTAIL.n156 B 0.013188f
C614 VTAIL.n157 B 0.012456f
C615 VTAIL.n158 B 0.023179f
C616 VTAIL.n159 B 0.023179f
C617 VTAIL.n160 B 0.012456f
C618 VTAIL.n161 B 0.013188f
C619 VTAIL.n162 B 0.02944f
C620 VTAIL.n163 B 0.02944f
C621 VTAIL.n164 B 0.013188f
C622 VTAIL.n165 B 0.012456f
C623 VTAIL.n166 B 0.023179f
C624 VTAIL.n167 B 0.023179f
C625 VTAIL.n168 B 0.012456f
C626 VTAIL.n169 B 0.013188f
C627 VTAIL.n170 B 0.02944f
C628 VTAIL.n171 B 0.02944f
C629 VTAIL.n172 B 0.013188f
C630 VTAIL.n173 B 0.012456f
C631 VTAIL.n174 B 0.023179f
C632 VTAIL.n175 B 0.023179f
C633 VTAIL.n176 B 0.012456f
C634 VTAIL.n177 B 0.012822f
C635 VTAIL.n178 B 0.012822f
C636 VTAIL.n179 B 0.02944f
C637 VTAIL.n180 B 0.02944f
C638 VTAIL.n181 B 0.013188f
C639 VTAIL.n182 B 0.012456f
C640 VTAIL.n183 B 0.023179f
C641 VTAIL.n184 B 0.023179f
C642 VTAIL.n185 B 0.012456f
C643 VTAIL.n186 B 0.013188f
C644 VTAIL.n187 B 0.02944f
C645 VTAIL.n188 B 0.06567f
C646 VTAIL.n189 B 0.013188f
C647 VTAIL.n190 B 0.012456f
C648 VTAIL.n191 B 0.058328f
C649 VTAIL.n192 B 0.037084f
C650 VTAIL.n193 B 0.442932f
C651 VTAIL.t11 B 0.310474f
C652 VTAIL.t10 B 0.310474f
C653 VTAIL.n194 B 2.75899f
C654 VTAIL.n195 B 0.643144f
C655 VTAIL.n196 B 0.033675f
C656 VTAIL.n197 B 0.023179f
C657 VTAIL.n198 B 0.012456f
C658 VTAIL.n199 B 0.02944f
C659 VTAIL.n200 B 0.013188f
C660 VTAIL.n201 B 0.023179f
C661 VTAIL.n202 B 0.012456f
C662 VTAIL.n203 B 0.02944f
C663 VTAIL.n204 B 0.013188f
C664 VTAIL.n205 B 0.023179f
C665 VTAIL.n206 B 0.012456f
C666 VTAIL.n207 B 0.02944f
C667 VTAIL.n208 B 0.02944f
C668 VTAIL.n209 B 0.013188f
C669 VTAIL.n210 B 0.023179f
C670 VTAIL.n211 B 0.012456f
C671 VTAIL.n212 B 0.02944f
C672 VTAIL.n213 B 0.013188f
C673 VTAIL.n214 B 0.023179f
C674 VTAIL.n215 B 0.012456f
C675 VTAIL.n216 B 0.02944f
C676 VTAIL.n217 B 0.013188f
C677 VTAIL.n218 B 0.023179f
C678 VTAIL.n219 B 0.012456f
C679 VTAIL.n220 B 0.02944f
C680 VTAIL.n221 B 0.013188f
C681 VTAIL.n222 B 0.023179f
C682 VTAIL.n223 B 0.012456f
C683 VTAIL.n224 B 0.02944f
C684 VTAIL.n225 B 0.013188f
C685 VTAIL.n226 B 0.162514f
C686 VTAIL.t8 B 0.048699f
C687 VTAIL.n227 B 0.02208f
C688 VTAIL.n228 B 0.017391f
C689 VTAIL.n229 B 0.012456f
C690 VTAIL.n230 B 1.71524f
C691 VTAIL.n231 B 0.023179f
C692 VTAIL.n232 B 0.012456f
C693 VTAIL.n233 B 0.013188f
C694 VTAIL.n234 B 0.02944f
C695 VTAIL.n235 B 0.02944f
C696 VTAIL.n236 B 0.013188f
C697 VTAIL.n237 B 0.012456f
C698 VTAIL.n238 B 0.023179f
C699 VTAIL.n239 B 0.023179f
C700 VTAIL.n240 B 0.012456f
C701 VTAIL.n241 B 0.013188f
C702 VTAIL.n242 B 0.02944f
C703 VTAIL.n243 B 0.02944f
C704 VTAIL.n244 B 0.013188f
C705 VTAIL.n245 B 0.012456f
C706 VTAIL.n246 B 0.023179f
C707 VTAIL.n247 B 0.023179f
C708 VTAIL.n248 B 0.012456f
C709 VTAIL.n249 B 0.013188f
C710 VTAIL.n250 B 0.02944f
C711 VTAIL.n251 B 0.02944f
C712 VTAIL.n252 B 0.013188f
C713 VTAIL.n253 B 0.012456f
C714 VTAIL.n254 B 0.023179f
C715 VTAIL.n255 B 0.023179f
C716 VTAIL.n256 B 0.012456f
C717 VTAIL.n257 B 0.013188f
C718 VTAIL.n258 B 0.02944f
C719 VTAIL.n259 B 0.02944f
C720 VTAIL.n260 B 0.013188f
C721 VTAIL.n261 B 0.012456f
C722 VTAIL.n262 B 0.023179f
C723 VTAIL.n263 B 0.023179f
C724 VTAIL.n264 B 0.012456f
C725 VTAIL.n265 B 0.013188f
C726 VTAIL.n266 B 0.02944f
C727 VTAIL.n267 B 0.02944f
C728 VTAIL.n268 B 0.013188f
C729 VTAIL.n269 B 0.012456f
C730 VTAIL.n270 B 0.023179f
C731 VTAIL.n271 B 0.023179f
C732 VTAIL.n272 B 0.012456f
C733 VTAIL.n273 B 0.012822f
C734 VTAIL.n274 B 0.012822f
C735 VTAIL.n275 B 0.02944f
C736 VTAIL.n276 B 0.02944f
C737 VTAIL.n277 B 0.013188f
C738 VTAIL.n278 B 0.012456f
C739 VTAIL.n279 B 0.023179f
C740 VTAIL.n280 B 0.023179f
C741 VTAIL.n281 B 0.012456f
C742 VTAIL.n282 B 0.013188f
C743 VTAIL.n283 B 0.02944f
C744 VTAIL.n284 B 0.06567f
C745 VTAIL.n285 B 0.013188f
C746 VTAIL.n286 B 0.012456f
C747 VTAIL.n287 B 0.058328f
C748 VTAIL.n288 B 0.037084f
C749 VTAIL.n289 B 1.94252f
C750 VTAIL.n290 B 0.033675f
C751 VTAIL.n291 B 0.023179f
C752 VTAIL.n292 B 0.012456f
C753 VTAIL.n293 B 0.02944f
C754 VTAIL.n294 B 0.013188f
C755 VTAIL.n295 B 0.023179f
C756 VTAIL.n296 B 0.012456f
C757 VTAIL.n297 B 0.02944f
C758 VTAIL.n298 B 0.013188f
C759 VTAIL.n299 B 0.023179f
C760 VTAIL.n300 B 0.012456f
C761 VTAIL.n301 B 0.02944f
C762 VTAIL.n302 B 0.013188f
C763 VTAIL.n303 B 0.023179f
C764 VTAIL.n304 B 0.012456f
C765 VTAIL.n305 B 0.02944f
C766 VTAIL.n306 B 0.013188f
C767 VTAIL.n307 B 0.023179f
C768 VTAIL.n308 B 0.012456f
C769 VTAIL.n309 B 0.02944f
C770 VTAIL.n310 B 0.013188f
C771 VTAIL.n311 B 0.023179f
C772 VTAIL.n312 B 0.012456f
C773 VTAIL.n313 B 0.02944f
C774 VTAIL.n314 B 0.013188f
C775 VTAIL.n315 B 0.023179f
C776 VTAIL.n316 B 0.012456f
C777 VTAIL.n317 B 0.02944f
C778 VTAIL.n318 B 0.013188f
C779 VTAIL.n319 B 0.162514f
C780 VTAIL.t2 B 0.048699f
C781 VTAIL.n320 B 0.02208f
C782 VTAIL.n321 B 0.017391f
C783 VTAIL.n322 B 0.012456f
C784 VTAIL.n323 B 1.71524f
C785 VTAIL.n324 B 0.023179f
C786 VTAIL.n325 B 0.012456f
C787 VTAIL.n326 B 0.013188f
C788 VTAIL.n327 B 0.02944f
C789 VTAIL.n328 B 0.02944f
C790 VTAIL.n329 B 0.013188f
C791 VTAIL.n330 B 0.012456f
C792 VTAIL.n331 B 0.023179f
C793 VTAIL.n332 B 0.023179f
C794 VTAIL.n333 B 0.012456f
C795 VTAIL.n334 B 0.013188f
C796 VTAIL.n335 B 0.02944f
C797 VTAIL.n336 B 0.02944f
C798 VTAIL.n337 B 0.013188f
C799 VTAIL.n338 B 0.012456f
C800 VTAIL.n339 B 0.023179f
C801 VTAIL.n340 B 0.023179f
C802 VTAIL.n341 B 0.012456f
C803 VTAIL.n342 B 0.013188f
C804 VTAIL.n343 B 0.02944f
C805 VTAIL.n344 B 0.02944f
C806 VTAIL.n345 B 0.013188f
C807 VTAIL.n346 B 0.012456f
C808 VTAIL.n347 B 0.023179f
C809 VTAIL.n348 B 0.023179f
C810 VTAIL.n349 B 0.012456f
C811 VTAIL.n350 B 0.013188f
C812 VTAIL.n351 B 0.02944f
C813 VTAIL.n352 B 0.02944f
C814 VTAIL.n353 B 0.013188f
C815 VTAIL.n354 B 0.012456f
C816 VTAIL.n355 B 0.023179f
C817 VTAIL.n356 B 0.023179f
C818 VTAIL.n357 B 0.012456f
C819 VTAIL.n358 B 0.013188f
C820 VTAIL.n359 B 0.02944f
C821 VTAIL.n360 B 0.02944f
C822 VTAIL.n361 B 0.02944f
C823 VTAIL.n362 B 0.013188f
C824 VTAIL.n363 B 0.012456f
C825 VTAIL.n364 B 0.023179f
C826 VTAIL.n365 B 0.023179f
C827 VTAIL.n366 B 0.012456f
C828 VTAIL.n367 B 0.012822f
C829 VTAIL.n368 B 0.012822f
C830 VTAIL.n369 B 0.02944f
C831 VTAIL.n370 B 0.02944f
C832 VTAIL.n371 B 0.013188f
C833 VTAIL.n372 B 0.012456f
C834 VTAIL.n373 B 0.023179f
C835 VTAIL.n374 B 0.023179f
C836 VTAIL.n375 B 0.012456f
C837 VTAIL.n376 B 0.013188f
C838 VTAIL.n377 B 0.02944f
C839 VTAIL.n378 B 0.06567f
C840 VTAIL.n379 B 0.013188f
C841 VTAIL.n380 B 0.012456f
C842 VTAIL.n381 B 0.058328f
C843 VTAIL.n382 B 0.037084f
C844 VTAIL.n383 B 1.87395f
C845 VP.n0 B 0.033866f
C846 VP.t2 B 3.06857f
C847 VP.n1 B 0.035872f
C848 VP.n2 B 0.018004f
C849 VP.n3 B 0.033555f
C850 VP.n4 B 0.018004f
C851 VP.t1 B 3.06857f
C852 VP.n5 B 0.035691f
C853 VP.n6 B 0.018004f
C854 VP.n7 B 0.033224f
C855 VP.n8 B 0.033866f
C856 VP.t4 B 3.06857f
C857 VP.n9 B 0.035872f
C858 VP.n10 B 0.018004f
C859 VP.n11 B 0.033555f
C860 VP.t0 B 3.33698f
C861 VP.t3 B 3.06857f
C862 VP.n12 B 1.13335f
C863 VP.n13 B 1.08371f
C864 VP.n14 B 0.229641f
C865 VP.n15 B 0.018004f
C866 VP.n16 B 0.033555f
C867 VP.n17 B 0.035691f
C868 VP.n18 B 0.014561f
C869 VP.n19 B 0.018004f
C870 VP.n20 B 0.018004f
C871 VP.n21 B 0.018004f
C872 VP.n22 B 0.033555f
C873 VP.n23 B 0.033224f
C874 VP.n24 B 1.13889f
C875 VP.n25 B 1.2407f
C876 VP.t5 B 3.06857f
C877 VP.n26 B 1.13889f
C878 VP.n27 B 1.2521f
C879 VP.n28 B 0.033866f
C880 VP.n29 B 0.018004f
C881 VP.n30 B 0.033555f
C882 VP.n31 B 0.035872f
C883 VP.n32 B 0.014561f
C884 VP.n33 B 0.018004f
C885 VP.n34 B 0.018004f
C886 VP.n35 B 0.018004f
C887 VP.n36 B 0.033555f
C888 VP.n37 B 0.033555f
C889 VP.n38 B 1.07693f
C890 VP.n39 B 0.018004f
C891 VP.n40 B 0.018004f
C892 VP.n41 B 0.018004f
C893 VP.n42 B 0.033555f
C894 VP.n43 B 0.035691f
C895 VP.n44 B 0.014561f
C896 VP.n45 B 0.018004f
C897 VP.n46 B 0.018004f
C898 VP.n47 B 0.018004f
C899 VP.n48 B 0.033555f
C900 VP.n49 B 0.033224f
C901 VP.n50 B 1.13889f
C902 VP.n51 B 0.051126f
.ends

