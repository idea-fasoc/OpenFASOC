* NGSPICE file created from diff_pair_sample_0049.ext - technology: sky130A

.subckt diff_pair_sample_0049 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t1 VN.t0 VTAIL.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=4.953 pd=26.18 as=4.953 ps=26.18 w=12.7 l=1.61
X1 VDD1.t1 VP.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=4.953 pd=26.18 as=4.953 ps=26.18 w=12.7 l=1.61
X2 VDD1.t0 VP.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=4.953 pd=26.18 as=4.953 ps=26.18 w=12.7 l=1.61
X3 VDD2.t0 VN.t1 VTAIL.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=4.953 pd=26.18 as=4.953 ps=26.18 w=12.7 l=1.61
X4 B.t15 B.t13 B.t14 B.t10 sky130_fd_pr__nfet_01v8 ad=4.953 pd=26.18 as=0 ps=0 w=12.7 l=1.61
X5 B.t12 B.t9 B.t11 B.t10 sky130_fd_pr__nfet_01v8 ad=4.953 pd=26.18 as=0 ps=0 w=12.7 l=1.61
X6 B.t8 B.t6 B.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=4.953 pd=26.18 as=0 ps=0 w=12.7 l=1.61
X7 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=4.953 pd=26.18 as=0 ps=0 w=12.7 l=1.61
R0 VN VN.t1 337.955
R1 VN VN.t0 295.255
R2 VTAIL.n278 VTAIL.n277 289.615
R3 VTAIL.n68 VTAIL.n67 289.615
R4 VTAIL.n208 VTAIL.n207 289.615
R5 VTAIL.n138 VTAIL.n137 289.615
R6 VTAIL.n232 VTAIL.n231 185
R7 VTAIL.n237 VTAIL.n236 185
R8 VTAIL.n239 VTAIL.n238 185
R9 VTAIL.n228 VTAIL.n227 185
R10 VTAIL.n245 VTAIL.n244 185
R11 VTAIL.n247 VTAIL.n246 185
R12 VTAIL.n224 VTAIL.n223 185
R13 VTAIL.n253 VTAIL.n252 185
R14 VTAIL.n255 VTAIL.n254 185
R15 VTAIL.n220 VTAIL.n219 185
R16 VTAIL.n261 VTAIL.n260 185
R17 VTAIL.n263 VTAIL.n262 185
R18 VTAIL.n216 VTAIL.n215 185
R19 VTAIL.n269 VTAIL.n268 185
R20 VTAIL.n271 VTAIL.n270 185
R21 VTAIL.n212 VTAIL.n211 185
R22 VTAIL.n277 VTAIL.n276 185
R23 VTAIL.n22 VTAIL.n21 185
R24 VTAIL.n27 VTAIL.n26 185
R25 VTAIL.n29 VTAIL.n28 185
R26 VTAIL.n18 VTAIL.n17 185
R27 VTAIL.n35 VTAIL.n34 185
R28 VTAIL.n37 VTAIL.n36 185
R29 VTAIL.n14 VTAIL.n13 185
R30 VTAIL.n43 VTAIL.n42 185
R31 VTAIL.n45 VTAIL.n44 185
R32 VTAIL.n10 VTAIL.n9 185
R33 VTAIL.n51 VTAIL.n50 185
R34 VTAIL.n53 VTAIL.n52 185
R35 VTAIL.n6 VTAIL.n5 185
R36 VTAIL.n59 VTAIL.n58 185
R37 VTAIL.n61 VTAIL.n60 185
R38 VTAIL.n2 VTAIL.n1 185
R39 VTAIL.n67 VTAIL.n66 185
R40 VTAIL.n207 VTAIL.n206 185
R41 VTAIL.n142 VTAIL.n141 185
R42 VTAIL.n201 VTAIL.n200 185
R43 VTAIL.n199 VTAIL.n198 185
R44 VTAIL.n146 VTAIL.n145 185
R45 VTAIL.n193 VTAIL.n192 185
R46 VTAIL.n191 VTAIL.n190 185
R47 VTAIL.n150 VTAIL.n149 185
R48 VTAIL.n185 VTAIL.n184 185
R49 VTAIL.n183 VTAIL.n182 185
R50 VTAIL.n154 VTAIL.n153 185
R51 VTAIL.n177 VTAIL.n176 185
R52 VTAIL.n175 VTAIL.n174 185
R53 VTAIL.n158 VTAIL.n157 185
R54 VTAIL.n169 VTAIL.n168 185
R55 VTAIL.n167 VTAIL.n166 185
R56 VTAIL.n162 VTAIL.n161 185
R57 VTAIL.n137 VTAIL.n136 185
R58 VTAIL.n72 VTAIL.n71 185
R59 VTAIL.n131 VTAIL.n130 185
R60 VTAIL.n129 VTAIL.n128 185
R61 VTAIL.n76 VTAIL.n75 185
R62 VTAIL.n123 VTAIL.n122 185
R63 VTAIL.n121 VTAIL.n120 185
R64 VTAIL.n80 VTAIL.n79 185
R65 VTAIL.n115 VTAIL.n114 185
R66 VTAIL.n113 VTAIL.n112 185
R67 VTAIL.n84 VTAIL.n83 185
R68 VTAIL.n107 VTAIL.n106 185
R69 VTAIL.n105 VTAIL.n104 185
R70 VTAIL.n88 VTAIL.n87 185
R71 VTAIL.n99 VTAIL.n98 185
R72 VTAIL.n97 VTAIL.n96 185
R73 VTAIL.n92 VTAIL.n91 185
R74 VTAIL.n233 VTAIL.t2 147.659
R75 VTAIL.n23 VTAIL.t0 147.659
R76 VTAIL.n163 VTAIL.t1 147.659
R77 VTAIL.n93 VTAIL.t3 147.659
R78 VTAIL.n237 VTAIL.n231 104.615
R79 VTAIL.n238 VTAIL.n237 104.615
R80 VTAIL.n238 VTAIL.n227 104.615
R81 VTAIL.n245 VTAIL.n227 104.615
R82 VTAIL.n246 VTAIL.n245 104.615
R83 VTAIL.n246 VTAIL.n223 104.615
R84 VTAIL.n253 VTAIL.n223 104.615
R85 VTAIL.n254 VTAIL.n253 104.615
R86 VTAIL.n254 VTAIL.n219 104.615
R87 VTAIL.n261 VTAIL.n219 104.615
R88 VTAIL.n262 VTAIL.n261 104.615
R89 VTAIL.n262 VTAIL.n215 104.615
R90 VTAIL.n269 VTAIL.n215 104.615
R91 VTAIL.n270 VTAIL.n269 104.615
R92 VTAIL.n270 VTAIL.n211 104.615
R93 VTAIL.n277 VTAIL.n211 104.615
R94 VTAIL.n27 VTAIL.n21 104.615
R95 VTAIL.n28 VTAIL.n27 104.615
R96 VTAIL.n28 VTAIL.n17 104.615
R97 VTAIL.n35 VTAIL.n17 104.615
R98 VTAIL.n36 VTAIL.n35 104.615
R99 VTAIL.n36 VTAIL.n13 104.615
R100 VTAIL.n43 VTAIL.n13 104.615
R101 VTAIL.n44 VTAIL.n43 104.615
R102 VTAIL.n44 VTAIL.n9 104.615
R103 VTAIL.n51 VTAIL.n9 104.615
R104 VTAIL.n52 VTAIL.n51 104.615
R105 VTAIL.n52 VTAIL.n5 104.615
R106 VTAIL.n59 VTAIL.n5 104.615
R107 VTAIL.n60 VTAIL.n59 104.615
R108 VTAIL.n60 VTAIL.n1 104.615
R109 VTAIL.n67 VTAIL.n1 104.615
R110 VTAIL.n207 VTAIL.n141 104.615
R111 VTAIL.n200 VTAIL.n141 104.615
R112 VTAIL.n200 VTAIL.n199 104.615
R113 VTAIL.n199 VTAIL.n145 104.615
R114 VTAIL.n192 VTAIL.n145 104.615
R115 VTAIL.n192 VTAIL.n191 104.615
R116 VTAIL.n191 VTAIL.n149 104.615
R117 VTAIL.n184 VTAIL.n149 104.615
R118 VTAIL.n184 VTAIL.n183 104.615
R119 VTAIL.n183 VTAIL.n153 104.615
R120 VTAIL.n176 VTAIL.n153 104.615
R121 VTAIL.n176 VTAIL.n175 104.615
R122 VTAIL.n175 VTAIL.n157 104.615
R123 VTAIL.n168 VTAIL.n157 104.615
R124 VTAIL.n168 VTAIL.n167 104.615
R125 VTAIL.n167 VTAIL.n161 104.615
R126 VTAIL.n137 VTAIL.n71 104.615
R127 VTAIL.n130 VTAIL.n71 104.615
R128 VTAIL.n130 VTAIL.n129 104.615
R129 VTAIL.n129 VTAIL.n75 104.615
R130 VTAIL.n122 VTAIL.n75 104.615
R131 VTAIL.n122 VTAIL.n121 104.615
R132 VTAIL.n121 VTAIL.n79 104.615
R133 VTAIL.n114 VTAIL.n79 104.615
R134 VTAIL.n114 VTAIL.n113 104.615
R135 VTAIL.n113 VTAIL.n83 104.615
R136 VTAIL.n106 VTAIL.n83 104.615
R137 VTAIL.n106 VTAIL.n105 104.615
R138 VTAIL.n105 VTAIL.n87 104.615
R139 VTAIL.n98 VTAIL.n87 104.615
R140 VTAIL.n98 VTAIL.n97 104.615
R141 VTAIL.n97 VTAIL.n91 104.615
R142 VTAIL.t2 VTAIL.n231 52.3082
R143 VTAIL.t0 VTAIL.n21 52.3082
R144 VTAIL.t1 VTAIL.n161 52.3082
R145 VTAIL.t3 VTAIL.n91 52.3082
R146 VTAIL.n279 VTAIL.n278 36.0641
R147 VTAIL.n69 VTAIL.n68 36.0641
R148 VTAIL.n209 VTAIL.n208 36.0641
R149 VTAIL.n139 VTAIL.n138 36.0641
R150 VTAIL.n139 VTAIL.n69 26.66
R151 VTAIL.n279 VTAIL.n209 24.9876
R152 VTAIL.n233 VTAIL.n232 15.6677
R153 VTAIL.n23 VTAIL.n22 15.6677
R154 VTAIL.n163 VTAIL.n162 15.6677
R155 VTAIL.n93 VTAIL.n92 15.6677
R156 VTAIL.n236 VTAIL.n235 12.8005
R157 VTAIL.n276 VTAIL.n210 12.8005
R158 VTAIL.n26 VTAIL.n25 12.8005
R159 VTAIL.n66 VTAIL.n0 12.8005
R160 VTAIL.n206 VTAIL.n140 12.8005
R161 VTAIL.n166 VTAIL.n165 12.8005
R162 VTAIL.n136 VTAIL.n70 12.8005
R163 VTAIL.n96 VTAIL.n95 12.8005
R164 VTAIL.n239 VTAIL.n230 12.0247
R165 VTAIL.n275 VTAIL.n212 12.0247
R166 VTAIL.n29 VTAIL.n20 12.0247
R167 VTAIL.n65 VTAIL.n2 12.0247
R168 VTAIL.n205 VTAIL.n142 12.0247
R169 VTAIL.n169 VTAIL.n160 12.0247
R170 VTAIL.n135 VTAIL.n72 12.0247
R171 VTAIL.n99 VTAIL.n90 12.0247
R172 VTAIL.n240 VTAIL.n228 11.249
R173 VTAIL.n272 VTAIL.n271 11.249
R174 VTAIL.n30 VTAIL.n18 11.249
R175 VTAIL.n62 VTAIL.n61 11.249
R176 VTAIL.n202 VTAIL.n201 11.249
R177 VTAIL.n170 VTAIL.n158 11.249
R178 VTAIL.n132 VTAIL.n131 11.249
R179 VTAIL.n100 VTAIL.n88 11.249
R180 VTAIL.n244 VTAIL.n243 10.4732
R181 VTAIL.n268 VTAIL.n214 10.4732
R182 VTAIL.n34 VTAIL.n33 10.4732
R183 VTAIL.n58 VTAIL.n4 10.4732
R184 VTAIL.n198 VTAIL.n144 10.4732
R185 VTAIL.n174 VTAIL.n173 10.4732
R186 VTAIL.n128 VTAIL.n74 10.4732
R187 VTAIL.n104 VTAIL.n103 10.4732
R188 VTAIL.n247 VTAIL.n226 9.69747
R189 VTAIL.n267 VTAIL.n216 9.69747
R190 VTAIL.n37 VTAIL.n16 9.69747
R191 VTAIL.n57 VTAIL.n6 9.69747
R192 VTAIL.n197 VTAIL.n146 9.69747
R193 VTAIL.n177 VTAIL.n156 9.69747
R194 VTAIL.n127 VTAIL.n76 9.69747
R195 VTAIL.n107 VTAIL.n86 9.69747
R196 VTAIL.n274 VTAIL.n210 9.45567
R197 VTAIL.n64 VTAIL.n0 9.45567
R198 VTAIL.n204 VTAIL.n140 9.45567
R199 VTAIL.n134 VTAIL.n70 9.45567
R200 VTAIL.n257 VTAIL.n256 9.3005
R201 VTAIL.n259 VTAIL.n258 9.3005
R202 VTAIL.n218 VTAIL.n217 9.3005
R203 VTAIL.n265 VTAIL.n264 9.3005
R204 VTAIL.n267 VTAIL.n266 9.3005
R205 VTAIL.n214 VTAIL.n213 9.3005
R206 VTAIL.n273 VTAIL.n272 9.3005
R207 VTAIL.n275 VTAIL.n274 9.3005
R208 VTAIL.n251 VTAIL.n250 9.3005
R209 VTAIL.n249 VTAIL.n248 9.3005
R210 VTAIL.n226 VTAIL.n225 9.3005
R211 VTAIL.n243 VTAIL.n242 9.3005
R212 VTAIL.n241 VTAIL.n240 9.3005
R213 VTAIL.n230 VTAIL.n229 9.3005
R214 VTAIL.n235 VTAIL.n234 9.3005
R215 VTAIL.n222 VTAIL.n221 9.3005
R216 VTAIL.n47 VTAIL.n46 9.3005
R217 VTAIL.n49 VTAIL.n48 9.3005
R218 VTAIL.n8 VTAIL.n7 9.3005
R219 VTAIL.n55 VTAIL.n54 9.3005
R220 VTAIL.n57 VTAIL.n56 9.3005
R221 VTAIL.n4 VTAIL.n3 9.3005
R222 VTAIL.n63 VTAIL.n62 9.3005
R223 VTAIL.n65 VTAIL.n64 9.3005
R224 VTAIL.n41 VTAIL.n40 9.3005
R225 VTAIL.n39 VTAIL.n38 9.3005
R226 VTAIL.n16 VTAIL.n15 9.3005
R227 VTAIL.n33 VTAIL.n32 9.3005
R228 VTAIL.n31 VTAIL.n30 9.3005
R229 VTAIL.n20 VTAIL.n19 9.3005
R230 VTAIL.n25 VTAIL.n24 9.3005
R231 VTAIL.n12 VTAIL.n11 9.3005
R232 VTAIL.n205 VTAIL.n204 9.3005
R233 VTAIL.n203 VTAIL.n202 9.3005
R234 VTAIL.n144 VTAIL.n143 9.3005
R235 VTAIL.n197 VTAIL.n196 9.3005
R236 VTAIL.n195 VTAIL.n194 9.3005
R237 VTAIL.n148 VTAIL.n147 9.3005
R238 VTAIL.n189 VTAIL.n188 9.3005
R239 VTAIL.n187 VTAIL.n186 9.3005
R240 VTAIL.n152 VTAIL.n151 9.3005
R241 VTAIL.n181 VTAIL.n180 9.3005
R242 VTAIL.n179 VTAIL.n178 9.3005
R243 VTAIL.n156 VTAIL.n155 9.3005
R244 VTAIL.n173 VTAIL.n172 9.3005
R245 VTAIL.n171 VTAIL.n170 9.3005
R246 VTAIL.n160 VTAIL.n159 9.3005
R247 VTAIL.n165 VTAIL.n164 9.3005
R248 VTAIL.n119 VTAIL.n118 9.3005
R249 VTAIL.n78 VTAIL.n77 9.3005
R250 VTAIL.n125 VTAIL.n124 9.3005
R251 VTAIL.n127 VTAIL.n126 9.3005
R252 VTAIL.n74 VTAIL.n73 9.3005
R253 VTAIL.n133 VTAIL.n132 9.3005
R254 VTAIL.n135 VTAIL.n134 9.3005
R255 VTAIL.n117 VTAIL.n116 9.3005
R256 VTAIL.n82 VTAIL.n81 9.3005
R257 VTAIL.n111 VTAIL.n110 9.3005
R258 VTAIL.n109 VTAIL.n108 9.3005
R259 VTAIL.n86 VTAIL.n85 9.3005
R260 VTAIL.n103 VTAIL.n102 9.3005
R261 VTAIL.n101 VTAIL.n100 9.3005
R262 VTAIL.n90 VTAIL.n89 9.3005
R263 VTAIL.n95 VTAIL.n94 9.3005
R264 VTAIL.n248 VTAIL.n224 8.92171
R265 VTAIL.n264 VTAIL.n263 8.92171
R266 VTAIL.n38 VTAIL.n14 8.92171
R267 VTAIL.n54 VTAIL.n53 8.92171
R268 VTAIL.n194 VTAIL.n193 8.92171
R269 VTAIL.n178 VTAIL.n154 8.92171
R270 VTAIL.n124 VTAIL.n123 8.92171
R271 VTAIL.n108 VTAIL.n84 8.92171
R272 VTAIL.n252 VTAIL.n251 8.14595
R273 VTAIL.n260 VTAIL.n218 8.14595
R274 VTAIL.n42 VTAIL.n41 8.14595
R275 VTAIL.n50 VTAIL.n8 8.14595
R276 VTAIL.n190 VTAIL.n148 8.14595
R277 VTAIL.n182 VTAIL.n181 8.14595
R278 VTAIL.n120 VTAIL.n78 8.14595
R279 VTAIL.n112 VTAIL.n111 8.14595
R280 VTAIL.n255 VTAIL.n222 7.3702
R281 VTAIL.n259 VTAIL.n220 7.3702
R282 VTAIL.n45 VTAIL.n12 7.3702
R283 VTAIL.n49 VTAIL.n10 7.3702
R284 VTAIL.n189 VTAIL.n150 7.3702
R285 VTAIL.n185 VTAIL.n152 7.3702
R286 VTAIL.n119 VTAIL.n80 7.3702
R287 VTAIL.n115 VTAIL.n82 7.3702
R288 VTAIL.n256 VTAIL.n255 6.59444
R289 VTAIL.n256 VTAIL.n220 6.59444
R290 VTAIL.n46 VTAIL.n45 6.59444
R291 VTAIL.n46 VTAIL.n10 6.59444
R292 VTAIL.n186 VTAIL.n150 6.59444
R293 VTAIL.n186 VTAIL.n185 6.59444
R294 VTAIL.n116 VTAIL.n80 6.59444
R295 VTAIL.n116 VTAIL.n115 6.59444
R296 VTAIL.n252 VTAIL.n222 5.81868
R297 VTAIL.n260 VTAIL.n259 5.81868
R298 VTAIL.n42 VTAIL.n12 5.81868
R299 VTAIL.n50 VTAIL.n49 5.81868
R300 VTAIL.n190 VTAIL.n189 5.81868
R301 VTAIL.n182 VTAIL.n152 5.81868
R302 VTAIL.n120 VTAIL.n119 5.81868
R303 VTAIL.n112 VTAIL.n82 5.81868
R304 VTAIL.n251 VTAIL.n224 5.04292
R305 VTAIL.n263 VTAIL.n218 5.04292
R306 VTAIL.n41 VTAIL.n14 5.04292
R307 VTAIL.n53 VTAIL.n8 5.04292
R308 VTAIL.n193 VTAIL.n148 5.04292
R309 VTAIL.n181 VTAIL.n154 5.04292
R310 VTAIL.n123 VTAIL.n78 5.04292
R311 VTAIL.n111 VTAIL.n84 5.04292
R312 VTAIL.n234 VTAIL.n233 4.38563
R313 VTAIL.n24 VTAIL.n23 4.38563
R314 VTAIL.n164 VTAIL.n163 4.38563
R315 VTAIL.n94 VTAIL.n93 4.38563
R316 VTAIL.n248 VTAIL.n247 4.26717
R317 VTAIL.n264 VTAIL.n216 4.26717
R318 VTAIL.n38 VTAIL.n37 4.26717
R319 VTAIL.n54 VTAIL.n6 4.26717
R320 VTAIL.n194 VTAIL.n146 4.26717
R321 VTAIL.n178 VTAIL.n177 4.26717
R322 VTAIL.n124 VTAIL.n76 4.26717
R323 VTAIL.n108 VTAIL.n107 4.26717
R324 VTAIL.n244 VTAIL.n226 3.49141
R325 VTAIL.n268 VTAIL.n267 3.49141
R326 VTAIL.n34 VTAIL.n16 3.49141
R327 VTAIL.n58 VTAIL.n57 3.49141
R328 VTAIL.n198 VTAIL.n197 3.49141
R329 VTAIL.n174 VTAIL.n156 3.49141
R330 VTAIL.n128 VTAIL.n127 3.49141
R331 VTAIL.n104 VTAIL.n86 3.49141
R332 VTAIL.n243 VTAIL.n228 2.71565
R333 VTAIL.n271 VTAIL.n214 2.71565
R334 VTAIL.n33 VTAIL.n18 2.71565
R335 VTAIL.n61 VTAIL.n4 2.71565
R336 VTAIL.n201 VTAIL.n144 2.71565
R337 VTAIL.n173 VTAIL.n158 2.71565
R338 VTAIL.n131 VTAIL.n74 2.71565
R339 VTAIL.n103 VTAIL.n88 2.71565
R340 VTAIL.n240 VTAIL.n239 1.93989
R341 VTAIL.n272 VTAIL.n212 1.93989
R342 VTAIL.n30 VTAIL.n29 1.93989
R343 VTAIL.n62 VTAIL.n2 1.93989
R344 VTAIL.n202 VTAIL.n142 1.93989
R345 VTAIL.n170 VTAIL.n169 1.93989
R346 VTAIL.n132 VTAIL.n72 1.93989
R347 VTAIL.n100 VTAIL.n99 1.93989
R348 VTAIL.n209 VTAIL.n139 1.30653
R349 VTAIL.n236 VTAIL.n230 1.16414
R350 VTAIL.n276 VTAIL.n275 1.16414
R351 VTAIL.n26 VTAIL.n20 1.16414
R352 VTAIL.n66 VTAIL.n65 1.16414
R353 VTAIL.n206 VTAIL.n205 1.16414
R354 VTAIL.n166 VTAIL.n160 1.16414
R355 VTAIL.n136 VTAIL.n135 1.16414
R356 VTAIL.n96 VTAIL.n90 1.16414
R357 VTAIL VTAIL.n69 0.946621
R358 VTAIL.n235 VTAIL.n232 0.388379
R359 VTAIL.n278 VTAIL.n210 0.388379
R360 VTAIL.n25 VTAIL.n22 0.388379
R361 VTAIL.n68 VTAIL.n0 0.388379
R362 VTAIL.n208 VTAIL.n140 0.388379
R363 VTAIL.n165 VTAIL.n162 0.388379
R364 VTAIL.n138 VTAIL.n70 0.388379
R365 VTAIL.n95 VTAIL.n92 0.388379
R366 VTAIL VTAIL.n279 0.360414
R367 VTAIL.n234 VTAIL.n229 0.155672
R368 VTAIL.n241 VTAIL.n229 0.155672
R369 VTAIL.n242 VTAIL.n241 0.155672
R370 VTAIL.n242 VTAIL.n225 0.155672
R371 VTAIL.n249 VTAIL.n225 0.155672
R372 VTAIL.n250 VTAIL.n249 0.155672
R373 VTAIL.n250 VTAIL.n221 0.155672
R374 VTAIL.n257 VTAIL.n221 0.155672
R375 VTAIL.n258 VTAIL.n257 0.155672
R376 VTAIL.n258 VTAIL.n217 0.155672
R377 VTAIL.n265 VTAIL.n217 0.155672
R378 VTAIL.n266 VTAIL.n265 0.155672
R379 VTAIL.n266 VTAIL.n213 0.155672
R380 VTAIL.n273 VTAIL.n213 0.155672
R381 VTAIL.n274 VTAIL.n273 0.155672
R382 VTAIL.n24 VTAIL.n19 0.155672
R383 VTAIL.n31 VTAIL.n19 0.155672
R384 VTAIL.n32 VTAIL.n31 0.155672
R385 VTAIL.n32 VTAIL.n15 0.155672
R386 VTAIL.n39 VTAIL.n15 0.155672
R387 VTAIL.n40 VTAIL.n39 0.155672
R388 VTAIL.n40 VTAIL.n11 0.155672
R389 VTAIL.n47 VTAIL.n11 0.155672
R390 VTAIL.n48 VTAIL.n47 0.155672
R391 VTAIL.n48 VTAIL.n7 0.155672
R392 VTAIL.n55 VTAIL.n7 0.155672
R393 VTAIL.n56 VTAIL.n55 0.155672
R394 VTAIL.n56 VTAIL.n3 0.155672
R395 VTAIL.n63 VTAIL.n3 0.155672
R396 VTAIL.n64 VTAIL.n63 0.155672
R397 VTAIL.n204 VTAIL.n203 0.155672
R398 VTAIL.n203 VTAIL.n143 0.155672
R399 VTAIL.n196 VTAIL.n143 0.155672
R400 VTAIL.n196 VTAIL.n195 0.155672
R401 VTAIL.n195 VTAIL.n147 0.155672
R402 VTAIL.n188 VTAIL.n147 0.155672
R403 VTAIL.n188 VTAIL.n187 0.155672
R404 VTAIL.n187 VTAIL.n151 0.155672
R405 VTAIL.n180 VTAIL.n151 0.155672
R406 VTAIL.n180 VTAIL.n179 0.155672
R407 VTAIL.n179 VTAIL.n155 0.155672
R408 VTAIL.n172 VTAIL.n155 0.155672
R409 VTAIL.n172 VTAIL.n171 0.155672
R410 VTAIL.n171 VTAIL.n159 0.155672
R411 VTAIL.n164 VTAIL.n159 0.155672
R412 VTAIL.n134 VTAIL.n133 0.155672
R413 VTAIL.n133 VTAIL.n73 0.155672
R414 VTAIL.n126 VTAIL.n73 0.155672
R415 VTAIL.n126 VTAIL.n125 0.155672
R416 VTAIL.n125 VTAIL.n77 0.155672
R417 VTAIL.n118 VTAIL.n77 0.155672
R418 VTAIL.n118 VTAIL.n117 0.155672
R419 VTAIL.n117 VTAIL.n81 0.155672
R420 VTAIL.n110 VTAIL.n81 0.155672
R421 VTAIL.n110 VTAIL.n109 0.155672
R422 VTAIL.n109 VTAIL.n85 0.155672
R423 VTAIL.n102 VTAIL.n85 0.155672
R424 VTAIL.n102 VTAIL.n101 0.155672
R425 VTAIL.n101 VTAIL.n89 0.155672
R426 VTAIL.n94 VTAIL.n89 0.155672
R427 VDD2.n137 VDD2.n136 289.615
R428 VDD2.n68 VDD2.n67 289.615
R429 VDD2.n136 VDD2.n135 185
R430 VDD2.n71 VDD2.n70 185
R431 VDD2.n130 VDD2.n129 185
R432 VDD2.n128 VDD2.n127 185
R433 VDD2.n75 VDD2.n74 185
R434 VDD2.n122 VDD2.n121 185
R435 VDD2.n120 VDD2.n119 185
R436 VDD2.n79 VDD2.n78 185
R437 VDD2.n114 VDD2.n113 185
R438 VDD2.n112 VDD2.n111 185
R439 VDD2.n83 VDD2.n82 185
R440 VDD2.n106 VDD2.n105 185
R441 VDD2.n104 VDD2.n103 185
R442 VDD2.n87 VDD2.n86 185
R443 VDD2.n98 VDD2.n97 185
R444 VDD2.n96 VDD2.n95 185
R445 VDD2.n91 VDD2.n90 185
R446 VDD2.n22 VDD2.n21 185
R447 VDD2.n27 VDD2.n26 185
R448 VDD2.n29 VDD2.n28 185
R449 VDD2.n18 VDD2.n17 185
R450 VDD2.n35 VDD2.n34 185
R451 VDD2.n37 VDD2.n36 185
R452 VDD2.n14 VDD2.n13 185
R453 VDD2.n43 VDD2.n42 185
R454 VDD2.n45 VDD2.n44 185
R455 VDD2.n10 VDD2.n9 185
R456 VDD2.n51 VDD2.n50 185
R457 VDD2.n53 VDD2.n52 185
R458 VDD2.n6 VDD2.n5 185
R459 VDD2.n59 VDD2.n58 185
R460 VDD2.n61 VDD2.n60 185
R461 VDD2.n2 VDD2.n1 185
R462 VDD2.n67 VDD2.n66 185
R463 VDD2.n23 VDD2.t1 147.659
R464 VDD2.n92 VDD2.t0 147.659
R465 VDD2.n136 VDD2.n70 104.615
R466 VDD2.n129 VDD2.n70 104.615
R467 VDD2.n129 VDD2.n128 104.615
R468 VDD2.n128 VDD2.n74 104.615
R469 VDD2.n121 VDD2.n74 104.615
R470 VDD2.n121 VDD2.n120 104.615
R471 VDD2.n120 VDD2.n78 104.615
R472 VDD2.n113 VDD2.n78 104.615
R473 VDD2.n113 VDD2.n112 104.615
R474 VDD2.n112 VDD2.n82 104.615
R475 VDD2.n105 VDD2.n82 104.615
R476 VDD2.n105 VDD2.n104 104.615
R477 VDD2.n104 VDD2.n86 104.615
R478 VDD2.n97 VDD2.n86 104.615
R479 VDD2.n97 VDD2.n96 104.615
R480 VDD2.n96 VDD2.n90 104.615
R481 VDD2.n27 VDD2.n21 104.615
R482 VDD2.n28 VDD2.n27 104.615
R483 VDD2.n28 VDD2.n17 104.615
R484 VDD2.n35 VDD2.n17 104.615
R485 VDD2.n36 VDD2.n35 104.615
R486 VDD2.n36 VDD2.n13 104.615
R487 VDD2.n43 VDD2.n13 104.615
R488 VDD2.n44 VDD2.n43 104.615
R489 VDD2.n44 VDD2.n9 104.615
R490 VDD2.n51 VDD2.n9 104.615
R491 VDD2.n52 VDD2.n51 104.615
R492 VDD2.n52 VDD2.n5 104.615
R493 VDD2.n59 VDD2.n5 104.615
R494 VDD2.n60 VDD2.n59 104.615
R495 VDD2.n60 VDD2.n1 104.615
R496 VDD2.n67 VDD2.n1 104.615
R497 VDD2.n138 VDD2.n68 90.6955
R498 VDD2.n138 VDD2.n137 52.7429
R499 VDD2.t0 VDD2.n90 52.3082
R500 VDD2.t1 VDD2.n21 52.3082
R501 VDD2.n92 VDD2.n91 15.6677
R502 VDD2.n23 VDD2.n22 15.6677
R503 VDD2.n135 VDD2.n69 12.8005
R504 VDD2.n95 VDD2.n94 12.8005
R505 VDD2.n26 VDD2.n25 12.8005
R506 VDD2.n66 VDD2.n0 12.8005
R507 VDD2.n134 VDD2.n71 12.0247
R508 VDD2.n98 VDD2.n89 12.0247
R509 VDD2.n29 VDD2.n20 12.0247
R510 VDD2.n65 VDD2.n2 12.0247
R511 VDD2.n131 VDD2.n130 11.249
R512 VDD2.n99 VDD2.n87 11.249
R513 VDD2.n30 VDD2.n18 11.249
R514 VDD2.n62 VDD2.n61 11.249
R515 VDD2.n127 VDD2.n73 10.4732
R516 VDD2.n103 VDD2.n102 10.4732
R517 VDD2.n34 VDD2.n33 10.4732
R518 VDD2.n58 VDD2.n4 10.4732
R519 VDD2.n126 VDD2.n75 9.69747
R520 VDD2.n106 VDD2.n85 9.69747
R521 VDD2.n37 VDD2.n16 9.69747
R522 VDD2.n57 VDD2.n6 9.69747
R523 VDD2.n133 VDD2.n69 9.45567
R524 VDD2.n64 VDD2.n0 9.45567
R525 VDD2.n134 VDD2.n133 9.3005
R526 VDD2.n132 VDD2.n131 9.3005
R527 VDD2.n73 VDD2.n72 9.3005
R528 VDD2.n126 VDD2.n125 9.3005
R529 VDD2.n124 VDD2.n123 9.3005
R530 VDD2.n77 VDD2.n76 9.3005
R531 VDD2.n118 VDD2.n117 9.3005
R532 VDD2.n116 VDD2.n115 9.3005
R533 VDD2.n81 VDD2.n80 9.3005
R534 VDD2.n110 VDD2.n109 9.3005
R535 VDD2.n108 VDD2.n107 9.3005
R536 VDD2.n85 VDD2.n84 9.3005
R537 VDD2.n102 VDD2.n101 9.3005
R538 VDD2.n100 VDD2.n99 9.3005
R539 VDD2.n89 VDD2.n88 9.3005
R540 VDD2.n94 VDD2.n93 9.3005
R541 VDD2.n47 VDD2.n46 9.3005
R542 VDD2.n49 VDD2.n48 9.3005
R543 VDD2.n8 VDD2.n7 9.3005
R544 VDD2.n55 VDD2.n54 9.3005
R545 VDD2.n57 VDD2.n56 9.3005
R546 VDD2.n4 VDD2.n3 9.3005
R547 VDD2.n63 VDD2.n62 9.3005
R548 VDD2.n65 VDD2.n64 9.3005
R549 VDD2.n41 VDD2.n40 9.3005
R550 VDD2.n39 VDD2.n38 9.3005
R551 VDD2.n16 VDD2.n15 9.3005
R552 VDD2.n33 VDD2.n32 9.3005
R553 VDD2.n31 VDD2.n30 9.3005
R554 VDD2.n20 VDD2.n19 9.3005
R555 VDD2.n25 VDD2.n24 9.3005
R556 VDD2.n12 VDD2.n11 9.3005
R557 VDD2.n123 VDD2.n122 8.92171
R558 VDD2.n107 VDD2.n83 8.92171
R559 VDD2.n38 VDD2.n14 8.92171
R560 VDD2.n54 VDD2.n53 8.92171
R561 VDD2.n119 VDD2.n77 8.14595
R562 VDD2.n111 VDD2.n110 8.14595
R563 VDD2.n42 VDD2.n41 8.14595
R564 VDD2.n50 VDD2.n8 8.14595
R565 VDD2.n118 VDD2.n79 7.3702
R566 VDD2.n114 VDD2.n81 7.3702
R567 VDD2.n45 VDD2.n12 7.3702
R568 VDD2.n49 VDD2.n10 7.3702
R569 VDD2.n115 VDD2.n79 6.59444
R570 VDD2.n115 VDD2.n114 6.59444
R571 VDD2.n46 VDD2.n45 6.59444
R572 VDD2.n46 VDD2.n10 6.59444
R573 VDD2.n119 VDD2.n118 5.81868
R574 VDD2.n111 VDD2.n81 5.81868
R575 VDD2.n42 VDD2.n12 5.81868
R576 VDD2.n50 VDD2.n49 5.81868
R577 VDD2.n122 VDD2.n77 5.04292
R578 VDD2.n110 VDD2.n83 5.04292
R579 VDD2.n41 VDD2.n14 5.04292
R580 VDD2.n53 VDD2.n8 5.04292
R581 VDD2.n24 VDD2.n23 4.38563
R582 VDD2.n93 VDD2.n92 4.38563
R583 VDD2.n123 VDD2.n75 4.26717
R584 VDD2.n107 VDD2.n106 4.26717
R585 VDD2.n38 VDD2.n37 4.26717
R586 VDD2.n54 VDD2.n6 4.26717
R587 VDD2.n127 VDD2.n126 3.49141
R588 VDD2.n103 VDD2.n85 3.49141
R589 VDD2.n34 VDD2.n16 3.49141
R590 VDD2.n58 VDD2.n57 3.49141
R591 VDD2.n130 VDD2.n73 2.71565
R592 VDD2.n102 VDD2.n87 2.71565
R593 VDD2.n33 VDD2.n18 2.71565
R594 VDD2.n61 VDD2.n4 2.71565
R595 VDD2.n131 VDD2.n71 1.93989
R596 VDD2.n99 VDD2.n98 1.93989
R597 VDD2.n30 VDD2.n29 1.93989
R598 VDD2.n62 VDD2.n2 1.93989
R599 VDD2.n135 VDD2.n134 1.16414
R600 VDD2.n95 VDD2.n89 1.16414
R601 VDD2.n26 VDD2.n20 1.16414
R602 VDD2.n66 VDD2.n65 1.16414
R603 VDD2 VDD2.n138 0.476793
R604 VDD2.n137 VDD2.n69 0.388379
R605 VDD2.n94 VDD2.n91 0.388379
R606 VDD2.n25 VDD2.n22 0.388379
R607 VDD2.n68 VDD2.n0 0.388379
R608 VDD2.n133 VDD2.n132 0.155672
R609 VDD2.n132 VDD2.n72 0.155672
R610 VDD2.n125 VDD2.n72 0.155672
R611 VDD2.n125 VDD2.n124 0.155672
R612 VDD2.n124 VDD2.n76 0.155672
R613 VDD2.n117 VDD2.n76 0.155672
R614 VDD2.n117 VDD2.n116 0.155672
R615 VDD2.n116 VDD2.n80 0.155672
R616 VDD2.n109 VDD2.n80 0.155672
R617 VDD2.n109 VDD2.n108 0.155672
R618 VDD2.n108 VDD2.n84 0.155672
R619 VDD2.n101 VDD2.n84 0.155672
R620 VDD2.n101 VDD2.n100 0.155672
R621 VDD2.n100 VDD2.n88 0.155672
R622 VDD2.n93 VDD2.n88 0.155672
R623 VDD2.n24 VDD2.n19 0.155672
R624 VDD2.n31 VDD2.n19 0.155672
R625 VDD2.n32 VDD2.n31 0.155672
R626 VDD2.n32 VDD2.n15 0.155672
R627 VDD2.n39 VDD2.n15 0.155672
R628 VDD2.n40 VDD2.n39 0.155672
R629 VDD2.n40 VDD2.n11 0.155672
R630 VDD2.n47 VDD2.n11 0.155672
R631 VDD2.n48 VDD2.n47 0.155672
R632 VDD2.n48 VDD2.n7 0.155672
R633 VDD2.n55 VDD2.n7 0.155672
R634 VDD2.n56 VDD2.n55 0.155672
R635 VDD2.n56 VDD2.n3 0.155672
R636 VDD2.n63 VDD2.n3 0.155672
R637 VDD2.n64 VDD2.n63 0.155672
R638 B.n651 B.n650 585
R639 B.n652 B.n651 585
R640 B.n281 B.n87 585
R641 B.n280 B.n279 585
R642 B.n278 B.n277 585
R643 B.n276 B.n275 585
R644 B.n274 B.n273 585
R645 B.n272 B.n271 585
R646 B.n270 B.n269 585
R647 B.n268 B.n267 585
R648 B.n266 B.n265 585
R649 B.n264 B.n263 585
R650 B.n262 B.n261 585
R651 B.n260 B.n259 585
R652 B.n258 B.n257 585
R653 B.n256 B.n255 585
R654 B.n254 B.n253 585
R655 B.n252 B.n251 585
R656 B.n250 B.n249 585
R657 B.n248 B.n247 585
R658 B.n246 B.n245 585
R659 B.n244 B.n243 585
R660 B.n242 B.n241 585
R661 B.n240 B.n239 585
R662 B.n238 B.n237 585
R663 B.n236 B.n235 585
R664 B.n234 B.n233 585
R665 B.n232 B.n231 585
R666 B.n230 B.n229 585
R667 B.n228 B.n227 585
R668 B.n226 B.n225 585
R669 B.n224 B.n223 585
R670 B.n222 B.n221 585
R671 B.n220 B.n219 585
R672 B.n218 B.n217 585
R673 B.n216 B.n215 585
R674 B.n214 B.n213 585
R675 B.n212 B.n211 585
R676 B.n210 B.n209 585
R677 B.n208 B.n207 585
R678 B.n206 B.n205 585
R679 B.n204 B.n203 585
R680 B.n202 B.n201 585
R681 B.n200 B.n199 585
R682 B.n198 B.n197 585
R683 B.n195 B.n194 585
R684 B.n193 B.n192 585
R685 B.n191 B.n190 585
R686 B.n189 B.n188 585
R687 B.n187 B.n186 585
R688 B.n185 B.n184 585
R689 B.n183 B.n182 585
R690 B.n181 B.n180 585
R691 B.n179 B.n178 585
R692 B.n177 B.n176 585
R693 B.n175 B.n174 585
R694 B.n173 B.n172 585
R695 B.n171 B.n170 585
R696 B.n169 B.n168 585
R697 B.n167 B.n166 585
R698 B.n165 B.n164 585
R699 B.n163 B.n162 585
R700 B.n161 B.n160 585
R701 B.n159 B.n158 585
R702 B.n157 B.n156 585
R703 B.n155 B.n154 585
R704 B.n153 B.n152 585
R705 B.n151 B.n150 585
R706 B.n149 B.n148 585
R707 B.n147 B.n146 585
R708 B.n145 B.n144 585
R709 B.n143 B.n142 585
R710 B.n141 B.n140 585
R711 B.n139 B.n138 585
R712 B.n137 B.n136 585
R713 B.n135 B.n134 585
R714 B.n133 B.n132 585
R715 B.n131 B.n130 585
R716 B.n129 B.n128 585
R717 B.n127 B.n126 585
R718 B.n125 B.n124 585
R719 B.n123 B.n122 585
R720 B.n121 B.n120 585
R721 B.n119 B.n118 585
R722 B.n117 B.n116 585
R723 B.n115 B.n114 585
R724 B.n113 B.n112 585
R725 B.n111 B.n110 585
R726 B.n109 B.n108 585
R727 B.n107 B.n106 585
R728 B.n105 B.n104 585
R729 B.n103 B.n102 585
R730 B.n101 B.n100 585
R731 B.n99 B.n98 585
R732 B.n97 B.n96 585
R733 B.n95 B.n94 585
R734 B.n39 B.n38 585
R735 B.n655 B.n654 585
R736 B.n649 B.n88 585
R737 B.n88 B.n36 585
R738 B.n648 B.n35 585
R739 B.n659 B.n35 585
R740 B.n647 B.n34 585
R741 B.n660 B.n34 585
R742 B.n646 B.n33 585
R743 B.n661 B.n33 585
R744 B.n645 B.n644 585
R745 B.n644 B.n29 585
R746 B.n643 B.n28 585
R747 B.n667 B.n28 585
R748 B.n642 B.n27 585
R749 B.n668 B.n27 585
R750 B.n641 B.n26 585
R751 B.n669 B.n26 585
R752 B.n640 B.n639 585
R753 B.n639 B.n22 585
R754 B.n638 B.n21 585
R755 B.n675 B.n21 585
R756 B.n637 B.n20 585
R757 B.n676 B.n20 585
R758 B.n636 B.n19 585
R759 B.n677 B.n19 585
R760 B.n635 B.n634 585
R761 B.n634 B.n15 585
R762 B.n633 B.n14 585
R763 B.n683 B.n14 585
R764 B.n632 B.n13 585
R765 B.n684 B.n13 585
R766 B.n631 B.n12 585
R767 B.n685 B.n12 585
R768 B.n630 B.n629 585
R769 B.n629 B.n628 585
R770 B.n627 B.n626 585
R771 B.n627 B.n8 585
R772 B.n625 B.n7 585
R773 B.n692 B.n7 585
R774 B.n624 B.n6 585
R775 B.n693 B.n6 585
R776 B.n623 B.n5 585
R777 B.n694 B.n5 585
R778 B.n622 B.n621 585
R779 B.n621 B.n4 585
R780 B.n620 B.n282 585
R781 B.n620 B.n619 585
R782 B.n610 B.n283 585
R783 B.n284 B.n283 585
R784 B.n612 B.n611 585
R785 B.n613 B.n612 585
R786 B.n609 B.n289 585
R787 B.n289 B.n288 585
R788 B.n608 B.n607 585
R789 B.n607 B.n606 585
R790 B.n291 B.n290 585
R791 B.n292 B.n291 585
R792 B.n599 B.n598 585
R793 B.n600 B.n599 585
R794 B.n597 B.n297 585
R795 B.n297 B.n296 585
R796 B.n596 B.n595 585
R797 B.n595 B.n594 585
R798 B.n299 B.n298 585
R799 B.n300 B.n299 585
R800 B.n587 B.n586 585
R801 B.n588 B.n587 585
R802 B.n585 B.n304 585
R803 B.n308 B.n304 585
R804 B.n584 B.n583 585
R805 B.n583 B.n582 585
R806 B.n306 B.n305 585
R807 B.n307 B.n306 585
R808 B.n575 B.n574 585
R809 B.n576 B.n575 585
R810 B.n573 B.n313 585
R811 B.n313 B.n312 585
R812 B.n572 B.n571 585
R813 B.n571 B.n570 585
R814 B.n315 B.n314 585
R815 B.n316 B.n315 585
R816 B.n566 B.n565 585
R817 B.n319 B.n318 585
R818 B.n562 B.n561 585
R819 B.n563 B.n562 585
R820 B.n560 B.n367 585
R821 B.n559 B.n558 585
R822 B.n557 B.n556 585
R823 B.n555 B.n554 585
R824 B.n553 B.n552 585
R825 B.n551 B.n550 585
R826 B.n549 B.n548 585
R827 B.n547 B.n546 585
R828 B.n545 B.n544 585
R829 B.n543 B.n542 585
R830 B.n541 B.n540 585
R831 B.n539 B.n538 585
R832 B.n537 B.n536 585
R833 B.n535 B.n534 585
R834 B.n533 B.n532 585
R835 B.n531 B.n530 585
R836 B.n529 B.n528 585
R837 B.n527 B.n526 585
R838 B.n525 B.n524 585
R839 B.n523 B.n522 585
R840 B.n521 B.n520 585
R841 B.n519 B.n518 585
R842 B.n517 B.n516 585
R843 B.n515 B.n514 585
R844 B.n513 B.n512 585
R845 B.n511 B.n510 585
R846 B.n509 B.n508 585
R847 B.n507 B.n506 585
R848 B.n505 B.n504 585
R849 B.n503 B.n502 585
R850 B.n501 B.n500 585
R851 B.n499 B.n498 585
R852 B.n497 B.n496 585
R853 B.n495 B.n494 585
R854 B.n493 B.n492 585
R855 B.n491 B.n490 585
R856 B.n489 B.n488 585
R857 B.n487 B.n486 585
R858 B.n485 B.n484 585
R859 B.n483 B.n482 585
R860 B.n481 B.n480 585
R861 B.n478 B.n477 585
R862 B.n476 B.n475 585
R863 B.n474 B.n473 585
R864 B.n472 B.n471 585
R865 B.n470 B.n469 585
R866 B.n468 B.n467 585
R867 B.n466 B.n465 585
R868 B.n464 B.n463 585
R869 B.n462 B.n461 585
R870 B.n460 B.n459 585
R871 B.n458 B.n457 585
R872 B.n456 B.n455 585
R873 B.n454 B.n453 585
R874 B.n452 B.n451 585
R875 B.n450 B.n449 585
R876 B.n448 B.n447 585
R877 B.n446 B.n445 585
R878 B.n444 B.n443 585
R879 B.n442 B.n441 585
R880 B.n440 B.n439 585
R881 B.n438 B.n437 585
R882 B.n436 B.n435 585
R883 B.n434 B.n433 585
R884 B.n432 B.n431 585
R885 B.n430 B.n429 585
R886 B.n428 B.n427 585
R887 B.n426 B.n425 585
R888 B.n424 B.n423 585
R889 B.n422 B.n421 585
R890 B.n420 B.n419 585
R891 B.n418 B.n417 585
R892 B.n416 B.n415 585
R893 B.n414 B.n413 585
R894 B.n412 B.n411 585
R895 B.n410 B.n409 585
R896 B.n408 B.n407 585
R897 B.n406 B.n405 585
R898 B.n404 B.n403 585
R899 B.n402 B.n401 585
R900 B.n400 B.n399 585
R901 B.n398 B.n397 585
R902 B.n396 B.n395 585
R903 B.n394 B.n393 585
R904 B.n392 B.n391 585
R905 B.n390 B.n389 585
R906 B.n388 B.n387 585
R907 B.n386 B.n385 585
R908 B.n384 B.n383 585
R909 B.n382 B.n381 585
R910 B.n380 B.n379 585
R911 B.n378 B.n377 585
R912 B.n376 B.n375 585
R913 B.n374 B.n373 585
R914 B.n567 B.n317 585
R915 B.n317 B.n316 585
R916 B.n569 B.n568 585
R917 B.n570 B.n569 585
R918 B.n311 B.n310 585
R919 B.n312 B.n311 585
R920 B.n578 B.n577 585
R921 B.n577 B.n576 585
R922 B.n579 B.n309 585
R923 B.n309 B.n307 585
R924 B.n581 B.n580 585
R925 B.n582 B.n581 585
R926 B.n303 B.n302 585
R927 B.n308 B.n303 585
R928 B.n590 B.n589 585
R929 B.n589 B.n588 585
R930 B.n591 B.n301 585
R931 B.n301 B.n300 585
R932 B.n593 B.n592 585
R933 B.n594 B.n593 585
R934 B.n295 B.n294 585
R935 B.n296 B.n295 585
R936 B.n602 B.n601 585
R937 B.n601 B.n600 585
R938 B.n603 B.n293 585
R939 B.n293 B.n292 585
R940 B.n605 B.n604 585
R941 B.n606 B.n605 585
R942 B.n287 B.n286 585
R943 B.n288 B.n287 585
R944 B.n615 B.n614 585
R945 B.n614 B.n613 585
R946 B.n616 B.n285 585
R947 B.n285 B.n284 585
R948 B.n618 B.n617 585
R949 B.n619 B.n618 585
R950 B.n3 B.n0 585
R951 B.n4 B.n3 585
R952 B.n691 B.n1 585
R953 B.n692 B.n691 585
R954 B.n690 B.n689 585
R955 B.n690 B.n8 585
R956 B.n688 B.n9 585
R957 B.n628 B.n9 585
R958 B.n687 B.n686 585
R959 B.n686 B.n685 585
R960 B.n11 B.n10 585
R961 B.n684 B.n11 585
R962 B.n682 B.n681 585
R963 B.n683 B.n682 585
R964 B.n680 B.n16 585
R965 B.n16 B.n15 585
R966 B.n679 B.n678 585
R967 B.n678 B.n677 585
R968 B.n18 B.n17 585
R969 B.n676 B.n18 585
R970 B.n674 B.n673 585
R971 B.n675 B.n674 585
R972 B.n672 B.n23 585
R973 B.n23 B.n22 585
R974 B.n671 B.n670 585
R975 B.n670 B.n669 585
R976 B.n25 B.n24 585
R977 B.n668 B.n25 585
R978 B.n666 B.n665 585
R979 B.n667 B.n666 585
R980 B.n664 B.n30 585
R981 B.n30 B.n29 585
R982 B.n663 B.n662 585
R983 B.n662 B.n661 585
R984 B.n32 B.n31 585
R985 B.n660 B.n32 585
R986 B.n658 B.n657 585
R987 B.n659 B.n658 585
R988 B.n656 B.n37 585
R989 B.n37 B.n36 585
R990 B.n695 B.n694 585
R991 B.n693 B.n2 585
R992 B.n654 B.n37 497.305
R993 B.n651 B.n88 497.305
R994 B.n373 B.n315 497.305
R995 B.n565 B.n317 497.305
R996 B.n91 B.t13 395.933
R997 B.n89 B.t9 395.933
R998 B.n370 B.t6 395.933
R999 B.n368 B.t2 395.933
R1000 B.n89 B.t11 331.733
R1001 B.n370 B.t8 331.733
R1002 B.n91 B.t14 331.733
R1003 B.n368 B.t5 331.733
R1004 B.n90 B.t12 294.108
R1005 B.n371 B.t7 294.108
R1006 B.n92 B.t15 294.108
R1007 B.n369 B.t4 294.108
R1008 B.n652 B.n86 256.663
R1009 B.n652 B.n85 256.663
R1010 B.n652 B.n84 256.663
R1011 B.n652 B.n83 256.663
R1012 B.n652 B.n82 256.663
R1013 B.n652 B.n81 256.663
R1014 B.n652 B.n80 256.663
R1015 B.n652 B.n79 256.663
R1016 B.n652 B.n78 256.663
R1017 B.n652 B.n77 256.663
R1018 B.n652 B.n76 256.663
R1019 B.n652 B.n75 256.663
R1020 B.n652 B.n74 256.663
R1021 B.n652 B.n73 256.663
R1022 B.n652 B.n72 256.663
R1023 B.n652 B.n71 256.663
R1024 B.n652 B.n70 256.663
R1025 B.n652 B.n69 256.663
R1026 B.n652 B.n68 256.663
R1027 B.n652 B.n67 256.663
R1028 B.n652 B.n66 256.663
R1029 B.n652 B.n65 256.663
R1030 B.n652 B.n64 256.663
R1031 B.n652 B.n63 256.663
R1032 B.n652 B.n62 256.663
R1033 B.n652 B.n61 256.663
R1034 B.n652 B.n60 256.663
R1035 B.n652 B.n59 256.663
R1036 B.n652 B.n58 256.663
R1037 B.n652 B.n57 256.663
R1038 B.n652 B.n56 256.663
R1039 B.n652 B.n55 256.663
R1040 B.n652 B.n54 256.663
R1041 B.n652 B.n53 256.663
R1042 B.n652 B.n52 256.663
R1043 B.n652 B.n51 256.663
R1044 B.n652 B.n50 256.663
R1045 B.n652 B.n49 256.663
R1046 B.n652 B.n48 256.663
R1047 B.n652 B.n47 256.663
R1048 B.n652 B.n46 256.663
R1049 B.n652 B.n45 256.663
R1050 B.n652 B.n44 256.663
R1051 B.n652 B.n43 256.663
R1052 B.n652 B.n42 256.663
R1053 B.n652 B.n41 256.663
R1054 B.n652 B.n40 256.663
R1055 B.n653 B.n652 256.663
R1056 B.n564 B.n563 256.663
R1057 B.n563 B.n320 256.663
R1058 B.n563 B.n321 256.663
R1059 B.n563 B.n322 256.663
R1060 B.n563 B.n323 256.663
R1061 B.n563 B.n324 256.663
R1062 B.n563 B.n325 256.663
R1063 B.n563 B.n326 256.663
R1064 B.n563 B.n327 256.663
R1065 B.n563 B.n328 256.663
R1066 B.n563 B.n329 256.663
R1067 B.n563 B.n330 256.663
R1068 B.n563 B.n331 256.663
R1069 B.n563 B.n332 256.663
R1070 B.n563 B.n333 256.663
R1071 B.n563 B.n334 256.663
R1072 B.n563 B.n335 256.663
R1073 B.n563 B.n336 256.663
R1074 B.n563 B.n337 256.663
R1075 B.n563 B.n338 256.663
R1076 B.n563 B.n339 256.663
R1077 B.n563 B.n340 256.663
R1078 B.n563 B.n341 256.663
R1079 B.n563 B.n342 256.663
R1080 B.n563 B.n343 256.663
R1081 B.n563 B.n344 256.663
R1082 B.n563 B.n345 256.663
R1083 B.n563 B.n346 256.663
R1084 B.n563 B.n347 256.663
R1085 B.n563 B.n348 256.663
R1086 B.n563 B.n349 256.663
R1087 B.n563 B.n350 256.663
R1088 B.n563 B.n351 256.663
R1089 B.n563 B.n352 256.663
R1090 B.n563 B.n353 256.663
R1091 B.n563 B.n354 256.663
R1092 B.n563 B.n355 256.663
R1093 B.n563 B.n356 256.663
R1094 B.n563 B.n357 256.663
R1095 B.n563 B.n358 256.663
R1096 B.n563 B.n359 256.663
R1097 B.n563 B.n360 256.663
R1098 B.n563 B.n361 256.663
R1099 B.n563 B.n362 256.663
R1100 B.n563 B.n363 256.663
R1101 B.n563 B.n364 256.663
R1102 B.n563 B.n365 256.663
R1103 B.n563 B.n366 256.663
R1104 B.n697 B.n696 256.663
R1105 B.n94 B.n39 163.367
R1106 B.n98 B.n97 163.367
R1107 B.n102 B.n101 163.367
R1108 B.n106 B.n105 163.367
R1109 B.n110 B.n109 163.367
R1110 B.n114 B.n113 163.367
R1111 B.n118 B.n117 163.367
R1112 B.n122 B.n121 163.367
R1113 B.n126 B.n125 163.367
R1114 B.n130 B.n129 163.367
R1115 B.n134 B.n133 163.367
R1116 B.n138 B.n137 163.367
R1117 B.n142 B.n141 163.367
R1118 B.n146 B.n145 163.367
R1119 B.n150 B.n149 163.367
R1120 B.n154 B.n153 163.367
R1121 B.n158 B.n157 163.367
R1122 B.n162 B.n161 163.367
R1123 B.n166 B.n165 163.367
R1124 B.n170 B.n169 163.367
R1125 B.n174 B.n173 163.367
R1126 B.n178 B.n177 163.367
R1127 B.n182 B.n181 163.367
R1128 B.n186 B.n185 163.367
R1129 B.n190 B.n189 163.367
R1130 B.n194 B.n193 163.367
R1131 B.n199 B.n198 163.367
R1132 B.n203 B.n202 163.367
R1133 B.n207 B.n206 163.367
R1134 B.n211 B.n210 163.367
R1135 B.n215 B.n214 163.367
R1136 B.n219 B.n218 163.367
R1137 B.n223 B.n222 163.367
R1138 B.n227 B.n226 163.367
R1139 B.n231 B.n230 163.367
R1140 B.n235 B.n234 163.367
R1141 B.n239 B.n238 163.367
R1142 B.n243 B.n242 163.367
R1143 B.n247 B.n246 163.367
R1144 B.n251 B.n250 163.367
R1145 B.n255 B.n254 163.367
R1146 B.n259 B.n258 163.367
R1147 B.n263 B.n262 163.367
R1148 B.n267 B.n266 163.367
R1149 B.n271 B.n270 163.367
R1150 B.n275 B.n274 163.367
R1151 B.n279 B.n278 163.367
R1152 B.n651 B.n87 163.367
R1153 B.n571 B.n315 163.367
R1154 B.n571 B.n313 163.367
R1155 B.n575 B.n313 163.367
R1156 B.n575 B.n306 163.367
R1157 B.n583 B.n306 163.367
R1158 B.n583 B.n304 163.367
R1159 B.n587 B.n304 163.367
R1160 B.n587 B.n299 163.367
R1161 B.n595 B.n299 163.367
R1162 B.n595 B.n297 163.367
R1163 B.n599 B.n297 163.367
R1164 B.n599 B.n291 163.367
R1165 B.n607 B.n291 163.367
R1166 B.n607 B.n289 163.367
R1167 B.n612 B.n289 163.367
R1168 B.n612 B.n283 163.367
R1169 B.n620 B.n283 163.367
R1170 B.n621 B.n620 163.367
R1171 B.n621 B.n5 163.367
R1172 B.n6 B.n5 163.367
R1173 B.n7 B.n6 163.367
R1174 B.n627 B.n7 163.367
R1175 B.n629 B.n627 163.367
R1176 B.n629 B.n12 163.367
R1177 B.n13 B.n12 163.367
R1178 B.n14 B.n13 163.367
R1179 B.n634 B.n14 163.367
R1180 B.n634 B.n19 163.367
R1181 B.n20 B.n19 163.367
R1182 B.n21 B.n20 163.367
R1183 B.n639 B.n21 163.367
R1184 B.n639 B.n26 163.367
R1185 B.n27 B.n26 163.367
R1186 B.n28 B.n27 163.367
R1187 B.n644 B.n28 163.367
R1188 B.n644 B.n33 163.367
R1189 B.n34 B.n33 163.367
R1190 B.n35 B.n34 163.367
R1191 B.n88 B.n35 163.367
R1192 B.n562 B.n319 163.367
R1193 B.n562 B.n367 163.367
R1194 B.n558 B.n557 163.367
R1195 B.n554 B.n553 163.367
R1196 B.n550 B.n549 163.367
R1197 B.n546 B.n545 163.367
R1198 B.n542 B.n541 163.367
R1199 B.n538 B.n537 163.367
R1200 B.n534 B.n533 163.367
R1201 B.n530 B.n529 163.367
R1202 B.n526 B.n525 163.367
R1203 B.n522 B.n521 163.367
R1204 B.n518 B.n517 163.367
R1205 B.n514 B.n513 163.367
R1206 B.n510 B.n509 163.367
R1207 B.n506 B.n505 163.367
R1208 B.n502 B.n501 163.367
R1209 B.n498 B.n497 163.367
R1210 B.n494 B.n493 163.367
R1211 B.n490 B.n489 163.367
R1212 B.n486 B.n485 163.367
R1213 B.n482 B.n481 163.367
R1214 B.n477 B.n476 163.367
R1215 B.n473 B.n472 163.367
R1216 B.n469 B.n468 163.367
R1217 B.n465 B.n464 163.367
R1218 B.n461 B.n460 163.367
R1219 B.n457 B.n456 163.367
R1220 B.n453 B.n452 163.367
R1221 B.n449 B.n448 163.367
R1222 B.n445 B.n444 163.367
R1223 B.n441 B.n440 163.367
R1224 B.n437 B.n436 163.367
R1225 B.n433 B.n432 163.367
R1226 B.n429 B.n428 163.367
R1227 B.n425 B.n424 163.367
R1228 B.n421 B.n420 163.367
R1229 B.n417 B.n416 163.367
R1230 B.n413 B.n412 163.367
R1231 B.n409 B.n408 163.367
R1232 B.n405 B.n404 163.367
R1233 B.n401 B.n400 163.367
R1234 B.n397 B.n396 163.367
R1235 B.n393 B.n392 163.367
R1236 B.n389 B.n388 163.367
R1237 B.n385 B.n384 163.367
R1238 B.n381 B.n380 163.367
R1239 B.n377 B.n376 163.367
R1240 B.n569 B.n317 163.367
R1241 B.n569 B.n311 163.367
R1242 B.n577 B.n311 163.367
R1243 B.n577 B.n309 163.367
R1244 B.n581 B.n309 163.367
R1245 B.n581 B.n303 163.367
R1246 B.n589 B.n303 163.367
R1247 B.n589 B.n301 163.367
R1248 B.n593 B.n301 163.367
R1249 B.n593 B.n295 163.367
R1250 B.n601 B.n295 163.367
R1251 B.n601 B.n293 163.367
R1252 B.n605 B.n293 163.367
R1253 B.n605 B.n287 163.367
R1254 B.n614 B.n287 163.367
R1255 B.n614 B.n285 163.367
R1256 B.n618 B.n285 163.367
R1257 B.n618 B.n3 163.367
R1258 B.n695 B.n3 163.367
R1259 B.n691 B.n2 163.367
R1260 B.n691 B.n690 163.367
R1261 B.n690 B.n9 163.367
R1262 B.n686 B.n9 163.367
R1263 B.n686 B.n11 163.367
R1264 B.n682 B.n11 163.367
R1265 B.n682 B.n16 163.367
R1266 B.n678 B.n16 163.367
R1267 B.n678 B.n18 163.367
R1268 B.n674 B.n18 163.367
R1269 B.n674 B.n23 163.367
R1270 B.n670 B.n23 163.367
R1271 B.n670 B.n25 163.367
R1272 B.n666 B.n25 163.367
R1273 B.n666 B.n30 163.367
R1274 B.n662 B.n30 163.367
R1275 B.n662 B.n32 163.367
R1276 B.n658 B.n32 163.367
R1277 B.n658 B.n37 163.367
R1278 B.n563 B.n316 76.4956
R1279 B.n652 B.n36 76.4956
R1280 B.n654 B.n653 71.676
R1281 B.n94 B.n40 71.676
R1282 B.n98 B.n41 71.676
R1283 B.n102 B.n42 71.676
R1284 B.n106 B.n43 71.676
R1285 B.n110 B.n44 71.676
R1286 B.n114 B.n45 71.676
R1287 B.n118 B.n46 71.676
R1288 B.n122 B.n47 71.676
R1289 B.n126 B.n48 71.676
R1290 B.n130 B.n49 71.676
R1291 B.n134 B.n50 71.676
R1292 B.n138 B.n51 71.676
R1293 B.n142 B.n52 71.676
R1294 B.n146 B.n53 71.676
R1295 B.n150 B.n54 71.676
R1296 B.n154 B.n55 71.676
R1297 B.n158 B.n56 71.676
R1298 B.n162 B.n57 71.676
R1299 B.n166 B.n58 71.676
R1300 B.n170 B.n59 71.676
R1301 B.n174 B.n60 71.676
R1302 B.n178 B.n61 71.676
R1303 B.n182 B.n62 71.676
R1304 B.n186 B.n63 71.676
R1305 B.n190 B.n64 71.676
R1306 B.n194 B.n65 71.676
R1307 B.n199 B.n66 71.676
R1308 B.n203 B.n67 71.676
R1309 B.n207 B.n68 71.676
R1310 B.n211 B.n69 71.676
R1311 B.n215 B.n70 71.676
R1312 B.n219 B.n71 71.676
R1313 B.n223 B.n72 71.676
R1314 B.n227 B.n73 71.676
R1315 B.n231 B.n74 71.676
R1316 B.n235 B.n75 71.676
R1317 B.n239 B.n76 71.676
R1318 B.n243 B.n77 71.676
R1319 B.n247 B.n78 71.676
R1320 B.n251 B.n79 71.676
R1321 B.n255 B.n80 71.676
R1322 B.n259 B.n81 71.676
R1323 B.n263 B.n82 71.676
R1324 B.n267 B.n83 71.676
R1325 B.n271 B.n84 71.676
R1326 B.n275 B.n85 71.676
R1327 B.n279 B.n86 71.676
R1328 B.n87 B.n86 71.676
R1329 B.n278 B.n85 71.676
R1330 B.n274 B.n84 71.676
R1331 B.n270 B.n83 71.676
R1332 B.n266 B.n82 71.676
R1333 B.n262 B.n81 71.676
R1334 B.n258 B.n80 71.676
R1335 B.n254 B.n79 71.676
R1336 B.n250 B.n78 71.676
R1337 B.n246 B.n77 71.676
R1338 B.n242 B.n76 71.676
R1339 B.n238 B.n75 71.676
R1340 B.n234 B.n74 71.676
R1341 B.n230 B.n73 71.676
R1342 B.n226 B.n72 71.676
R1343 B.n222 B.n71 71.676
R1344 B.n218 B.n70 71.676
R1345 B.n214 B.n69 71.676
R1346 B.n210 B.n68 71.676
R1347 B.n206 B.n67 71.676
R1348 B.n202 B.n66 71.676
R1349 B.n198 B.n65 71.676
R1350 B.n193 B.n64 71.676
R1351 B.n189 B.n63 71.676
R1352 B.n185 B.n62 71.676
R1353 B.n181 B.n61 71.676
R1354 B.n177 B.n60 71.676
R1355 B.n173 B.n59 71.676
R1356 B.n169 B.n58 71.676
R1357 B.n165 B.n57 71.676
R1358 B.n161 B.n56 71.676
R1359 B.n157 B.n55 71.676
R1360 B.n153 B.n54 71.676
R1361 B.n149 B.n53 71.676
R1362 B.n145 B.n52 71.676
R1363 B.n141 B.n51 71.676
R1364 B.n137 B.n50 71.676
R1365 B.n133 B.n49 71.676
R1366 B.n129 B.n48 71.676
R1367 B.n125 B.n47 71.676
R1368 B.n121 B.n46 71.676
R1369 B.n117 B.n45 71.676
R1370 B.n113 B.n44 71.676
R1371 B.n109 B.n43 71.676
R1372 B.n105 B.n42 71.676
R1373 B.n101 B.n41 71.676
R1374 B.n97 B.n40 71.676
R1375 B.n653 B.n39 71.676
R1376 B.n565 B.n564 71.676
R1377 B.n367 B.n320 71.676
R1378 B.n557 B.n321 71.676
R1379 B.n553 B.n322 71.676
R1380 B.n549 B.n323 71.676
R1381 B.n545 B.n324 71.676
R1382 B.n541 B.n325 71.676
R1383 B.n537 B.n326 71.676
R1384 B.n533 B.n327 71.676
R1385 B.n529 B.n328 71.676
R1386 B.n525 B.n329 71.676
R1387 B.n521 B.n330 71.676
R1388 B.n517 B.n331 71.676
R1389 B.n513 B.n332 71.676
R1390 B.n509 B.n333 71.676
R1391 B.n505 B.n334 71.676
R1392 B.n501 B.n335 71.676
R1393 B.n497 B.n336 71.676
R1394 B.n493 B.n337 71.676
R1395 B.n489 B.n338 71.676
R1396 B.n485 B.n339 71.676
R1397 B.n481 B.n340 71.676
R1398 B.n476 B.n341 71.676
R1399 B.n472 B.n342 71.676
R1400 B.n468 B.n343 71.676
R1401 B.n464 B.n344 71.676
R1402 B.n460 B.n345 71.676
R1403 B.n456 B.n346 71.676
R1404 B.n452 B.n347 71.676
R1405 B.n448 B.n348 71.676
R1406 B.n444 B.n349 71.676
R1407 B.n440 B.n350 71.676
R1408 B.n436 B.n351 71.676
R1409 B.n432 B.n352 71.676
R1410 B.n428 B.n353 71.676
R1411 B.n424 B.n354 71.676
R1412 B.n420 B.n355 71.676
R1413 B.n416 B.n356 71.676
R1414 B.n412 B.n357 71.676
R1415 B.n408 B.n358 71.676
R1416 B.n404 B.n359 71.676
R1417 B.n400 B.n360 71.676
R1418 B.n396 B.n361 71.676
R1419 B.n392 B.n362 71.676
R1420 B.n388 B.n363 71.676
R1421 B.n384 B.n364 71.676
R1422 B.n380 B.n365 71.676
R1423 B.n376 B.n366 71.676
R1424 B.n564 B.n319 71.676
R1425 B.n558 B.n320 71.676
R1426 B.n554 B.n321 71.676
R1427 B.n550 B.n322 71.676
R1428 B.n546 B.n323 71.676
R1429 B.n542 B.n324 71.676
R1430 B.n538 B.n325 71.676
R1431 B.n534 B.n326 71.676
R1432 B.n530 B.n327 71.676
R1433 B.n526 B.n328 71.676
R1434 B.n522 B.n329 71.676
R1435 B.n518 B.n330 71.676
R1436 B.n514 B.n331 71.676
R1437 B.n510 B.n332 71.676
R1438 B.n506 B.n333 71.676
R1439 B.n502 B.n334 71.676
R1440 B.n498 B.n335 71.676
R1441 B.n494 B.n336 71.676
R1442 B.n490 B.n337 71.676
R1443 B.n486 B.n338 71.676
R1444 B.n482 B.n339 71.676
R1445 B.n477 B.n340 71.676
R1446 B.n473 B.n341 71.676
R1447 B.n469 B.n342 71.676
R1448 B.n465 B.n343 71.676
R1449 B.n461 B.n344 71.676
R1450 B.n457 B.n345 71.676
R1451 B.n453 B.n346 71.676
R1452 B.n449 B.n347 71.676
R1453 B.n445 B.n348 71.676
R1454 B.n441 B.n349 71.676
R1455 B.n437 B.n350 71.676
R1456 B.n433 B.n351 71.676
R1457 B.n429 B.n352 71.676
R1458 B.n425 B.n353 71.676
R1459 B.n421 B.n354 71.676
R1460 B.n417 B.n355 71.676
R1461 B.n413 B.n356 71.676
R1462 B.n409 B.n357 71.676
R1463 B.n405 B.n358 71.676
R1464 B.n401 B.n359 71.676
R1465 B.n397 B.n360 71.676
R1466 B.n393 B.n361 71.676
R1467 B.n389 B.n362 71.676
R1468 B.n385 B.n363 71.676
R1469 B.n381 B.n364 71.676
R1470 B.n377 B.n365 71.676
R1471 B.n373 B.n366 71.676
R1472 B.n696 B.n695 71.676
R1473 B.n696 B.n2 71.676
R1474 B.n93 B.n92 59.5399
R1475 B.n196 B.n90 59.5399
R1476 B.n372 B.n371 59.5399
R1477 B.n479 B.n369 59.5399
R1478 B.n570 B.n316 41.6138
R1479 B.n570 B.n312 41.6138
R1480 B.n576 B.n312 41.6138
R1481 B.n576 B.n307 41.6138
R1482 B.n582 B.n307 41.6138
R1483 B.n582 B.n308 41.6138
R1484 B.n588 B.n300 41.6138
R1485 B.n594 B.n300 41.6138
R1486 B.n594 B.n296 41.6138
R1487 B.n600 B.n296 41.6138
R1488 B.n600 B.n292 41.6138
R1489 B.n606 B.n292 41.6138
R1490 B.n606 B.n288 41.6138
R1491 B.n613 B.n288 41.6138
R1492 B.n619 B.n284 41.6138
R1493 B.n619 B.n4 41.6138
R1494 B.n694 B.n4 41.6138
R1495 B.n694 B.n693 41.6138
R1496 B.n693 B.n692 41.6138
R1497 B.n692 B.n8 41.6138
R1498 B.n628 B.n8 41.6138
R1499 B.n685 B.n684 41.6138
R1500 B.n684 B.n683 41.6138
R1501 B.n683 B.n15 41.6138
R1502 B.n677 B.n15 41.6138
R1503 B.n677 B.n676 41.6138
R1504 B.n676 B.n675 41.6138
R1505 B.n675 B.n22 41.6138
R1506 B.n669 B.n22 41.6138
R1507 B.n668 B.n667 41.6138
R1508 B.n667 B.n29 41.6138
R1509 B.n661 B.n29 41.6138
R1510 B.n661 B.n660 41.6138
R1511 B.n660 B.n659 41.6138
R1512 B.n659 B.n36 41.6138
R1513 B.t0 B.n284 39.778
R1514 B.n628 B.t1 39.778
R1515 B.n92 B.n91 37.6247
R1516 B.n90 B.n89 37.6247
R1517 B.n371 B.n370 37.6247
R1518 B.n369 B.n368 37.6247
R1519 B.n588 B.t3 36.1062
R1520 B.n669 B.t10 36.1062
R1521 B.n567 B.n566 32.3127
R1522 B.n374 B.n314 32.3127
R1523 B.n650 B.n649 32.3127
R1524 B.n656 B.n655 32.3127
R1525 B B.n697 18.0485
R1526 B.n568 B.n567 10.6151
R1527 B.n568 B.n310 10.6151
R1528 B.n578 B.n310 10.6151
R1529 B.n579 B.n578 10.6151
R1530 B.n580 B.n579 10.6151
R1531 B.n580 B.n302 10.6151
R1532 B.n590 B.n302 10.6151
R1533 B.n591 B.n590 10.6151
R1534 B.n592 B.n591 10.6151
R1535 B.n592 B.n294 10.6151
R1536 B.n602 B.n294 10.6151
R1537 B.n603 B.n602 10.6151
R1538 B.n604 B.n603 10.6151
R1539 B.n604 B.n286 10.6151
R1540 B.n615 B.n286 10.6151
R1541 B.n616 B.n615 10.6151
R1542 B.n617 B.n616 10.6151
R1543 B.n617 B.n0 10.6151
R1544 B.n566 B.n318 10.6151
R1545 B.n561 B.n318 10.6151
R1546 B.n561 B.n560 10.6151
R1547 B.n560 B.n559 10.6151
R1548 B.n559 B.n556 10.6151
R1549 B.n556 B.n555 10.6151
R1550 B.n555 B.n552 10.6151
R1551 B.n552 B.n551 10.6151
R1552 B.n551 B.n548 10.6151
R1553 B.n548 B.n547 10.6151
R1554 B.n547 B.n544 10.6151
R1555 B.n544 B.n543 10.6151
R1556 B.n543 B.n540 10.6151
R1557 B.n540 B.n539 10.6151
R1558 B.n539 B.n536 10.6151
R1559 B.n536 B.n535 10.6151
R1560 B.n535 B.n532 10.6151
R1561 B.n532 B.n531 10.6151
R1562 B.n531 B.n528 10.6151
R1563 B.n528 B.n527 10.6151
R1564 B.n527 B.n524 10.6151
R1565 B.n524 B.n523 10.6151
R1566 B.n523 B.n520 10.6151
R1567 B.n520 B.n519 10.6151
R1568 B.n519 B.n516 10.6151
R1569 B.n516 B.n515 10.6151
R1570 B.n515 B.n512 10.6151
R1571 B.n512 B.n511 10.6151
R1572 B.n511 B.n508 10.6151
R1573 B.n508 B.n507 10.6151
R1574 B.n507 B.n504 10.6151
R1575 B.n504 B.n503 10.6151
R1576 B.n503 B.n500 10.6151
R1577 B.n500 B.n499 10.6151
R1578 B.n499 B.n496 10.6151
R1579 B.n496 B.n495 10.6151
R1580 B.n495 B.n492 10.6151
R1581 B.n492 B.n491 10.6151
R1582 B.n491 B.n488 10.6151
R1583 B.n488 B.n487 10.6151
R1584 B.n487 B.n484 10.6151
R1585 B.n484 B.n483 10.6151
R1586 B.n483 B.n480 10.6151
R1587 B.n478 B.n475 10.6151
R1588 B.n475 B.n474 10.6151
R1589 B.n474 B.n471 10.6151
R1590 B.n471 B.n470 10.6151
R1591 B.n470 B.n467 10.6151
R1592 B.n467 B.n466 10.6151
R1593 B.n466 B.n463 10.6151
R1594 B.n463 B.n462 10.6151
R1595 B.n459 B.n458 10.6151
R1596 B.n458 B.n455 10.6151
R1597 B.n455 B.n454 10.6151
R1598 B.n454 B.n451 10.6151
R1599 B.n451 B.n450 10.6151
R1600 B.n450 B.n447 10.6151
R1601 B.n447 B.n446 10.6151
R1602 B.n446 B.n443 10.6151
R1603 B.n443 B.n442 10.6151
R1604 B.n442 B.n439 10.6151
R1605 B.n439 B.n438 10.6151
R1606 B.n438 B.n435 10.6151
R1607 B.n435 B.n434 10.6151
R1608 B.n434 B.n431 10.6151
R1609 B.n431 B.n430 10.6151
R1610 B.n430 B.n427 10.6151
R1611 B.n427 B.n426 10.6151
R1612 B.n426 B.n423 10.6151
R1613 B.n423 B.n422 10.6151
R1614 B.n422 B.n419 10.6151
R1615 B.n419 B.n418 10.6151
R1616 B.n418 B.n415 10.6151
R1617 B.n415 B.n414 10.6151
R1618 B.n414 B.n411 10.6151
R1619 B.n411 B.n410 10.6151
R1620 B.n410 B.n407 10.6151
R1621 B.n407 B.n406 10.6151
R1622 B.n406 B.n403 10.6151
R1623 B.n403 B.n402 10.6151
R1624 B.n402 B.n399 10.6151
R1625 B.n399 B.n398 10.6151
R1626 B.n398 B.n395 10.6151
R1627 B.n395 B.n394 10.6151
R1628 B.n394 B.n391 10.6151
R1629 B.n391 B.n390 10.6151
R1630 B.n390 B.n387 10.6151
R1631 B.n387 B.n386 10.6151
R1632 B.n386 B.n383 10.6151
R1633 B.n383 B.n382 10.6151
R1634 B.n382 B.n379 10.6151
R1635 B.n379 B.n378 10.6151
R1636 B.n378 B.n375 10.6151
R1637 B.n375 B.n374 10.6151
R1638 B.n572 B.n314 10.6151
R1639 B.n573 B.n572 10.6151
R1640 B.n574 B.n573 10.6151
R1641 B.n574 B.n305 10.6151
R1642 B.n584 B.n305 10.6151
R1643 B.n585 B.n584 10.6151
R1644 B.n586 B.n585 10.6151
R1645 B.n586 B.n298 10.6151
R1646 B.n596 B.n298 10.6151
R1647 B.n597 B.n596 10.6151
R1648 B.n598 B.n597 10.6151
R1649 B.n598 B.n290 10.6151
R1650 B.n608 B.n290 10.6151
R1651 B.n609 B.n608 10.6151
R1652 B.n611 B.n609 10.6151
R1653 B.n611 B.n610 10.6151
R1654 B.n610 B.n282 10.6151
R1655 B.n622 B.n282 10.6151
R1656 B.n623 B.n622 10.6151
R1657 B.n624 B.n623 10.6151
R1658 B.n625 B.n624 10.6151
R1659 B.n626 B.n625 10.6151
R1660 B.n630 B.n626 10.6151
R1661 B.n631 B.n630 10.6151
R1662 B.n632 B.n631 10.6151
R1663 B.n633 B.n632 10.6151
R1664 B.n635 B.n633 10.6151
R1665 B.n636 B.n635 10.6151
R1666 B.n637 B.n636 10.6151
R1667 B.n638 B.n637 10.6151
R1668 B.n640 B.n638 10.6151
R1669 B.n641 B.n640 10.6151
R1670 B.n642 B.n641 10.6151
R1671 B.n643 B.n642 10.6151
R1672 B.n645 B.n643 10.6151
R1673 B.n646 B.n645 10.6151
R1674 B.n647 B.n646 10.6151
R1675 B.n648 B.n647 10.6151
R1676 B.n649 B.n648 10.6151
R1677 B.n689 B.n1 10.6151
R1678 B.n689 B.n688 10.6151
R1679 B.n688 B.n687 10.6151
R1680 B.n687 B.n10 10.6151
R1681 B.n681 B.n10 10.6151
R1682 B.n681 B.n680 10.6151
R1683 B.n680 B.n679 10.6151
R1684 B.n679 B.n17 10.6151
R1685 B.n673 B.n17 10.6151
R1686 B.n673 B.n672 10.6151
R1687 B.n672 B.n671 10.6151
R1688 B.n671 B.n24 10.6151
R1689 B.n665 B.n24 10.6151
R1690 B.n665 B.n664 10.6151
R1691 B.n664 B.n663 10.6151
R1692 B.n663 B.n31 10.6151
R1693 B.n657 B.n31 10.6151
R1694 B.n657 B.n656 10.6151
R1695 B.n655 B.n38 10.6151
R1696 B.n95 B.n38 10.6151
R1697 B.n96 B.n95 10.6151
R1698 B.n99 B.n96 10.6151
R1699 B.n100 B.n99 10.6151
R1700 B.n103 B.n100 10.6151
R1701 B.n104 B.n103 10.6151
R1702 B.n107 B.n104 10.6151
R1703 B.n108 B.n107 10.6151
R1704 B.n111 B.n108 10.6151
R1705 B.n112 B.n111 10.6151
R1706 B.n115 B.n112 10.6151
R1707 B.n116 B.n115 10.6151
R1708 B.n119 B.n116 10.6151
R1709 B.n120 B.n119 10.6151
R1710 B.n123 B.n120 10.6151
R1711 B.n124 B.n123 10.6151
R1712 B.n127 B.n124 10.6151
R1713 B.n128 B.n127 10.6151
R1714 B.n131 B.n128 10.6151
R1715 B.n132 B.n131 10.6151
R1716 B.n135 B.n132 10.6151
R1717 B.n136 B.n135 10.6151
R1718 B.n139 B.n136 10.6151
R1719 B.n140 B.n139 10.6151
R1720 B.n143 B.n140 10.6151
R1721 B.n144 B.n143 10.6151
R1722 B.n147 B.n144 10.6151
R1723 B.n148 B.n147 10.6151
R1724 B.n151 B.n148 10.6151
R1725 B.n152 B.n151 10.6151
R1726 B.n155 B.n152 10.6151
R1727 B.n156 B.n155 10.6151
R1728 B.n159 B.n156 10.6151
R1729 B.n160 B.n159 10.6151
R1730 B.n163 B.n160 10.6151
R1731 B.n164 B.n163 10.6151
R1732 B.n167 B.n164 10.6151
R1733 B.n168 B.n167 10.6151
R1734 B.n171 B.n168 10.6151
R1735 B.n172 B.n171 10.6151
R1736 B.n175 B.n172 10.6151
R1737 B.n176 B.n175 10.6151
R1738 B.n180 B.n179 10.6151
R1739 B.n183 B.n180 10.6151
R1740 B.n184 B.n183 10.6151
R1741 B.n187 B.n184 10.6151
R1742 B.n188 B.n187 10.6151
R1743 B.n191 B.n188 10.6151
R1744 B.n192 B.n191 10.6151
R1745 B.n195 B.n192 10.6151
R1746 B.n200 B.n197 10.6151
R1747 B.n201 B.n200 10.6151
R1748 B.n204 B.n201 10.6151
R1749 B.n205 B.n204 10.6151
R1750 B.n208 B.n205 10.6151
R1751 B.n209 B.n208 10.6151
R1752 B.n212 B.n209 10.6151
R1753 B.n213 B.n212 10.6151
R1754 B.n216 B.n213 10.6151
R1755 B.n217 B.n216 10.6151
R1756 B.n220 B.n217 10.6151
R1757 B.n221 B.n220 10.6151
R1758 B.n224 B.n221 10.6151
R1759 B.n225 B.n224 10.6151
R1760 B.n228 B.n225 10.6151
R1761 B.n229 B.n228 10.6151
R1762 B.n232 B.n229 10.6151
R1763 B.n233 B.n232 10.6151
R1764 B.n236 B.n233 10.6151
R1765 B.n237 B.n236 10.6151
R1766 B.n240 B.n237 10.6151
R1767 B.n241 B.n240 10.6151
R1768 B.n244 B.n241 10.6151
R1769 B.n245 B.n244 10.6151
R1770 B.n248 B.n245 10.6151
R1771 B.n249 B.n248 10.6151
R1772 B.n252 B.n249 10.6151
R1773 B.n253 B.n252 10.6151
R1774 B.n256 B.n253 10.6151
R1775 B.n257 B.n256 10.6151
R1776 B.n260 B.n257 10.6151
R1777 B.n261 B.n260 10.6151
R1778 B.n264 B.n261 10.6151
R1779 B.n265 B.n264 10.6151
R1780 B.n268 B.n265 10.6151
R1781 B.n269 B.n268 10.6151
R1782 B.n272 B.n269 10.6151
R1783 B.n273 B.n272 10.6151
R1784 B.n276 B.n273 10.6151
R1785 B.n277 B.n276 10.6151
R1786 B.n280 B.n277 10.6151
R1787 B.n281 B.n280 10.6151
R1788 B.n650 B.n281 10.6151
R1789 B.n697 B.n0 8.11757
R1790 B.n697 B.n1 8.11757
R1791 B.n479 B.n478 6.5566
R1792 B.n462 B.n372 6.5566
R1793 B.n179 B.n93 6.5566
R1794 B.n196 B.n195 6.5566
R1795 B.n308 B.t3 5.50815
R1796 B.t10 B.n668 5.50815
R1797 B.n480 B.n479 4.05904
R1798 B.n459 B.n372 4.05904
R1799 B.n176 B.n93 4.05904
R1800 B.n197 B.n196 4.05904
R1801 B.n613 B.t0 1.83638
R1802 B.n685 B.t1 1.83638
R1803 VP.n0 VP.t1 337.671
R1804 VP.n0 VP.t0 295.108
R1805 VP VP.n0 0.146778
R1806 VDD1.n68 VDD1.n67 289.615
R1807 VDD1.n137 VDD1.n136 289.615
R1808 VDD1.n67 VDD1.n66 185
R1809 VDD1.n2 VDD1.n1 185
R1810 VDD1.n61 VDD1.n60 185
R1811 VDD1.n59 VDD1.n58 185
R1812 VDD1.n6 VDD1.n5 185
R1813 VDD1.n53 VDD1.n52 185
R1814 VDD1.n51 VDD1.n50 185
R1815 VDD1.n10 VDD1.n9 185
R1816 VDD1.n45 VDD1.n44 185
R1817 VDD1.n43 VDD1.n42 185
R1818 VDD1.n14 VDD1.n13 185
R1819 VDD1.n37 VDD1.n36 185
R1820 VDD1.n35 VDD1.n34 185
R1821 VDD1.n18 VDD1.n17 185
R1822 VDD1.n29 VDD1.n28 185
R1823 VDD1.n27 VDD1.n26 185
R1824 VDD1.n22 VDD1.n21 185
R1825 VDD1.n91 VDD1.n90 185
R1826 VDD1.n96 VDD1.n95 185
R1827 VDD1.n98 VDD1.n97 185
R1828 VDD1.n87 VDD1.n86 185
R1829 VDD1.n104 VDD1.n103 185
R1830 VDD1.n106 VDD1.n105 185
R1831 VDD1.n83 VDD1.n82 185
R1832 VDD1.n112 VDD1.n111 185
R1833 VDD1.n114 VDD1.n113 185
R1834 VDD1.n79 VDD1.n78 185
R1835 VDD1.n120 VDD1.n119 185
R1836 VDD1.n122 VDD1.n121 185
R1837 VDD1.n75 VDD1.n74 185
R1838 VDD1.n128 VDD1.n127 185
R1839 VDD1.n130 VDD1.n129 185
R1840 VDD1.n71 VDD1.n70 185
R1841 VDD1.n136 VDD1.n135 185
R1842 VDD1.n92 VDD1.t1 147.659
R1843 VDD1.n23 VDD1.t0 147.659
R1844 VDD1.n67 VDD1.n1 104.615
R1845 VDD1.n60 VDD1.n1 104.615
R1846 VDD1.n60 VDD1.n59 104.615
R1847 VDD1.n59 VDD1.n5 104.615
R1848 VDD1.n52 VDD1.n5 104.615
R1849 VDD1.n52 VDD1.n51 104.615
R1850 VDD1.n51 VDD1.n9 104.615
R1851 VDD1.n44 VDD1.n9 104.615
R1852 VDD1.n44 VDD1.n43 104.615
R1853 VDD1.n43 VDD1.n13 104.615
R1854 VDD1.n36 VDD1.n13 104.615
R1855 VDD1.n36 VDD1.n35 104.615
R1856 VDD1.n35 VDD1.n17 104.615
R1857 VDD1.n28 VDD1.n17 104.615
R1858 VDD1.n28 VDD1.n27 104.615
R1859 VDD1.n27 VDD1.n21 104.615
R1860 VDD1.n96 VDD1.n90 104.615
R1861 VDD1.n97 VDD1.n96 104.615
R1862 VDD1.n97 VDD1.n86 104.615
R1863 VDD1.n104 VDD1.n86 104.615
R1864 VDD1.n105 VDD1.n104 104.615
R1865 VDD1.n105 VDD1.n82 104.615
R1866 VDD1.n112 VDD1.n82 104.615
R1867 VDD1.n113 VDD1.n112 104.615
R1868 VDD1.n113 VDD1.n78 104.615
R1869 VDD1.n120 VDD1.n78 104.615
R1870 VDD1.n121 VDD1.n120 104.615
R1871 VDD1.n121 VDD1.n74 104.615
R1872 VDD1.n128 VDD1.n74 104.615
R1873 VDD1.n129 VDD1.n128 104.615
R1874 VDD1.n129 VDD1.n70 104.615
R1875 VDD1.n136 VDD1.n70 104.615
R1876 VDD1 VDD1.n137 91.6384
R1877 VDD1 VDD1.n68 53.2192
R1878 VDD1.t0 VDD1.n21 52.3082
R1879 VDD1.t1 VDD1.n90 52.3082
R1880 VDD1.n23 VDD1.n22 15.6677
R1881 VDD1.n92 VDD1.n91 15.6677
R1882 VDD1.n66 VDD1.n0 12.8005
R1883 VDD1.n26 VDD1.n25 12.8005
R1884 VDD1.n95 VDD1.n94 12.8005
R1885 VDD1.n135 VDD1.n69 12.8005
R1886 VDD1.n65 VDD1.n2 12.0247
R1887 VDD1.n29 VDD1.n20 12.0247
R1888 VDD1.n98 VDD1.n89 12.0247
R1889 VDD1.n134 VDD1.n71 12.0247
R1890 VDD1.n62 VDD1.n61 11.249
R1891 VDD1.n30 VDD1.n18 11.249
R1892 VDD1.n99 VDD1.n87 11.249
R1893 VDD1.n131 VDD1.n130 11.249
R1894 VDD1.n58 VDD1.n4 10.4732
R1895 VDD1.n34 VDD1.n33 10.4732
R1896 VDD1.n103 VDD1.n102 10.4732
R1897 VDD1.n127 VDD1.n73 10.4732
R1898 VDD1.n57 VDD1.n6 9.69747
R1899 VDD1.n37 VDD1.n16 9.69747
R1900 VDD1.n106 VDD1.n85 9.69747
R1901 VDD1.n126 VDD1.n75 9.69747
R1902 VDD1.n64 VDD1.n0 9.45567
R1903 VDD1.n133 VDD1.n69 9.45567
R1904 VDD1.n65 VDD1.n64 9.3005
R1905 VDD1.n63 VDD1.n62 9.3005
R1906 VDD1.n4 VDD1.n3 9.3005
R1907 VDD1.n57 VDD1.n56 9.3005
R1908 VDD1.n55 VDD1.n54 9.3005
R1909 VDD1.n8 VDD1.n7 9.3005
R1910 VDD1.n49 VDD1.n48 9.3005
R1911 VDD1.n47 VDD1.n46 9.3005
R1912 VDD1.n12 VDD1.n11 9.3005
R1913 VDD1.n41 VDD1.n40 9.3005
R1914 VDD1.n39 VDD1.n38 9.3005
R1915 VDD1.n16 VDD1.n15 9.3005
R1916 VDD1.n33 VDD1.n32 9.3005
R1917 VDD1.n31 VDD1.n30 9.3005
R1918 VDD1.n20 VDD1.n19 9.3005
R1919 VDD1.n25 VDD1.n24 9.3005
R1920 VDD1.n116 VDD1.n115 9.3005
R1921 VDD1.n118 VDD1.n117 9.3005
R1922 VDD1.n77 VDD1.n76 9.3005
R1923 VDD1.n124 VDD1.n123 9.3005
R1924 VDD1.n126 VDD1.n125 9.3005
R1925 VDD1.n73 VDD1.n72 9.3005
R1926 VDD1.n132 VDD1.n131 9.3005
R1927 VDD1.n134 VDD1.n133 9.3005
R1928 VDD1.n110 VDD1.n109 9.3005
R1929 VDD1.n108 VDD1.n107 9.3005
R1930 VDD1.n85 VDD1.n84 9.3005
R1931 VDD1.n102 VDD1.n101 9.3005
R1932 VDD1.n100 VDD1.n99 9.3005
R1933 VDD1.n89 VDD1.n88 9.3005
R1934 VDD1.n94 VDD1.n93 9.3005
R1935 VDD1.n81 VDD1.n80 9.3005
R1936 VDD1.n54 VDD1.n53 8.92171
R1937 VDD1.n38 VDD1.n14 8.92171
R1938 VDD1.n107 VDD1.n83 8.92171
R1939 VDD1.n123 VDD1.n122 8.92171
R1940 VDD1.n50 VDD1.n8 8.14595
R1941 VDD1.n42 VDD1.n41 8.14595
R1942 VDD1.n111 VDD1.n110 8.14595
R1943 VDD1.n119 VDD1.n77 8.14595
R1944 VDD1.n49 VDD1.n10 7.3702
R1945 VDD1.n45 VDD1.n12 7.3702
R1946 VDD1.n114 VDD1.n81 7.3702
R1947 VDD1.n118 VDD1.n79 7.3702
R1948 VDD1.n46 VDD1.n10 6.59444
R1949 VDD1.n46 VDD1.n45 6.59444
R1950 VDD1.n115 VDD1.n114 6.59444
R1951 VDD1.n115 VDD1.n79 6.59444
R1952 VDD1.n50 VDD1.n49 5.81868
R1953 VDD1.n42 VDD1.n12 5.81868
R1954 VDD1.n111 VDD1.n81 5.81868
R1955 VDD1.n119 VDD1.n118 5.81868
R1956 VDD1.n53 VDD1.n8 5.04292
R1957 VDD1.n41 VDD1.n14 5.04292
R1958 VDD1.n110 VDD1.n83 5.04292
R1959 VDD1.n122 VDD1.n77 5.04292
R1960 VDD1.n93 VDD1.n92 4.38563
R1961 VDD1.n24 VDD1.n23 4.38563
R1962 VDD1.n54 VDD1.n6 4.26717
R1963 VDD1.n38 VDD1.n37 4.26717
R1964 VDD1.n107 VDD1.n106 4.26717
R1965 VDD1.n123 VDD1.n75 4.26717
R1966 VDD1.n58 VDD1.n57 3.49141
R1967 VDD1.n34 VDD1.n16 3.49141
R1968 VDD1.n103 VDD1.n85 3.49141
R1969 VDD1.n127 VDD1.n126 3.49141
R1970 VDD1.n61 VDD1.n4 2.71565
R1971 VDD1.n33 VDD1.n18 2.71565
R1972 VDD1.n102 VDD1.n87 2.71565
R1973 VDD1.n130 VDD1.n73 2.71565
R1974 VDD1.n62 VDD1.n2 1.93989
R1975 VDD1.n30 VDD1.n29 1.93989
R1976 VDD1.n99 VDD1.n98 1.93989
R1977 VDD1.n131 VDD1.n71 1.93989
R1978 VDD1.n66 VDD1.n65 1.16414
R1979 VDD1.n26 VDD1.n20 1.16414
R1980 VDD1.n95 VDD1.n89 1.16414
R1981 VDD1.n135 VDD1.n134 1.16414
R1982 VDD1.n68 VDD1.n0 0.388379
R1983 VDD1.n25 VDD1.n22 0.388379
R1984 VDD1.n94 VDD1.n91 0.388379
R1985 VDD1.n137 VDD1.n69 0.388379
R1986 VDD1.n64 VDD1.n63 0.155672
R1987 VDD1.n63 VDD1.n3 0.155672
R1988 VDD1.n56 VDD1.n3 0.155672
R1989 VDD1.n56 VDD1.n55 0.155672
R1990 VDD1.n55 VDD1.n7 0.155672
R1991 VDD1.n48 VDD1.n7 0.155672
R1992 VDD1.n48 VDD1.n47 0.155672
R1993 VDD1.n47 VDD1.n11 0.155672
R1994 VDD1.n40 VDD1.n11 0.155672
R1995 VDD1.n40 VDD1.n39 0.155672
R1996 VDD1.n39 VDD1.n15 0.155672
R1997 VDD1.n32 VDD1.n15 0.155672
R1998 VDD1.n32 VDD1.n31 0.155672
R1999 VDD1.n31 VDD1.n19 0.155672
R2000 VDD1.n24 VDD1.n19 0.155672
R2001 VDD1.n93 VDD1.n88 0.155672
R2002 VDD1.n100 VDD1.n88 0.155672
R2003 VDD1.n101 VDD1.n100 0.155672
R2004 VDD1.n101 VDD1.n84 0.155672
R2005 VDD1.n108 VDD1.n84 0.155672
R2006 VDD1.n109 VDD1.n108 0.155672
R2007 VDD1.n109 VDD1.n80 0.155672
R2008 VDD1.n116 VDD1.n80 0.155672
R2009 VDD1.n117 VDD1.n116 0.155672
R2010 VDD1.n117 VDD1.n76 0.155672
R2011 VDD1.n124 VDD1.n76 0.155672
R2012 VDD1.n125 VDD1.n124 0.155672
R2013 VDD1.n125 VDD1.n72 0.155672
R2014 VDD1.n132 VDD1.n72 0.155672
R2015 VDD1.n133 VDD1.n132 0.155672
C0 VDD2 VDD1 0.558672f
C1 VTAIL VN 2.24357f
C2 VN VP 5.11387f
C3 VN VDD1 0.148002f
C4 VTAIL VP 2.25798f
C5 VN VDD2 2.67359f
C6 VTAIL VDD1 5.24891f
C7 VP VDD1 2.8142f
C8 VTAIL VDD2 5.29118f
C9 VP VDD2 0.291998f
C10 VDD2 B 4.20889f
C11 VDD1 B 6.805799f
C12 VTAIL B 7.1319f
C13 VN B 9.809731f
C14 VP B 5.196122f
C15 VDD1.n0 B 0.011325f
C16 VDD1.n1 B 0.025493f
C17 VDD1.n2 B 0.01142f
C18 VDD1.n3 B 0.020071f
C19 VDD1.n4 B 0.010785f
C20 VDD1.n5 B 0.025493f
C21 VDD1.n6 B 0.01142f
C22 VDD1.n7 B 0.020071f
C23 VDD1.n8 B 0.010785f
C24 VDD1.n9 B 0.025493f
C25 VDD1.n10 B 0.01142f
C26 VDD1.n11 B 0.020071f
C27 VDD1.n12 B 0.010785f
C28 VDD1.n13 B 0.025493f
C29 VDD1.n14 B 0.01142f
C30 VDD1.n15 B 0.020071f
C31 VDD1.n16 B 0.010785f
C32 VDD1.n17 B 0.025493f
C33 VDD1.n18 B 0.01142f
C34 VDD1.n19 B 0.020071f
C35 VDD1.n20 B 0.010785f
C36 VDD1.n21 B 0.019119f
C37 VDD1.n22 B 0.015059f
C38 VDD1.t0 B 0.041876f
C39 VDD1.n23 B 0.119333f
C40 VDD1.n24 B 1.09428f
C41 VDD1.n25 B 0.010785f
C42 VDD1.n26 B 0.01142f
C43 VDD1.n27 B 0.025493f
C44 VDD1.n28 B 0.025493f
C45 VDD1.n29 B 0.01142f
C46 VDD1.n30 B 0.010785f
C47 VDD1.n31 B 0.020071f
C48 VDD1.n32 B 0.020071f
C49 VDD1.n33 B 0.010785f
C50 VDD1.n34 B 0.01142f
C51 VDD1.n35 B 0.025493f
C52 VDD1.n36 B 0.025493f
C53 VDD1.n37 B 0.01142f
C54 VDD1.n38 B 0.010785f
C55 VDD1.n39 B 0.020071f
C56 VDD1.n40 B 0.020071f
C57 VDD1.n41 B 0.010785f
C58 VDD1.n42 B 0.01142f
C59 VDD1.n43 B 0.025493f
C60 VDD1.n44 B 0.025493f
C61 VDD1.n45 B 0.01142f
C62 VDD1.n46 B 0.010785f
C63 VDD1.n47 B 0.020071f
C64 VDD1.n48 B 0.020071f
C65 VDD1.n49 B 0.010785f
C66 VDD1.n50 B 0.01142f
C67 VDD1.n51 B 0.025493f
C68 VDD1.n52 B 0.025493f
C69 VDD1.n53 B 0.01142f
C70 VDD1.n54 B 0.010785f
C71 VDD1.n55 B 0.020071f
C72 VDD1.n56 B 0.020071f
C73 VDD1.n57 B 0.010785f
C74 VDD1.n58 B 0.01142f
C75 VDD1.n59 B 0.025493f
C76 VDD1.n60 B 0.025493f
C77 VDD1.n61 B 0.01142f
C78 VDD1.n62 B 0.010785f
C79 VDD1.n63 B 0.020071f
C80 VDD1.n64 B 0.052425f
C81 VDD1.n65 B 0.010785f
C82 VDD1.n66 B 0.01142f
C83 VDD1.n67 B 0.052792f
C84 VDD1.n68 B 0.059148f
C85 VDD1.n69 B 0.011325f
C86 VDD1.n70 B 0.025493f
C87 VDD1.n71 B 0.01142f
C88 VDD1.n72 B 0.020071f
C89 VDD1.n73 B 0.010785f
C90 VDD1.n74 B 0.025493f
C91 VDD1.n75 B 0.01142f
C92 VDD1.n76 B 0.020071f
C93 VDD1.n77 B 0.010785f
C94 VDD1.n78 B 0.025493f
C95 VDD1.n79 B 0.01142f
C96 VDD1.n80 B 0.020071f
C97 VDD1.n81 B 0.010785f
C98 VDD1.n82 B 0.025493f
C99 VDD1.n83 B 0.01142f
C100 VDD1.n84 B 0.020071f
C101 VDD1.n85 B 0.010785f
C102 VDD1.n86 B 0.025493f
C103 VDD1.n87 B 0.01142f
C104 VDD1.n88 B 0.020071f
C105 VDD1.n89 B 0.010785f
C106 VDD1.n90 B 0.019119f
C107 VDD1.n91 B 0.015059f
C108 VDD1.t1 B 0.041876f
C109 VDD1.n92 B 0.119333f
C110 VDD1.n93 B 1.09428f
C111 VDD1.n94 B 0.010785f
C112 VDD1.n95 B 0.01142f
C113 VDD1.n96 B 0.025493f
C114 VDD1.n97 B 0.025493f
C115 VDD1.n98 B 0.01142f
C116 VDD1.n99 B 0.010785f
C117 VDD1.n100 B 0.020071f
C118 VDD1.n101 B 0.020071f
C119 VDD1.n102 B 0.010785f
C120 VDD1.n103 B 0.01142f
C121 VDD1.n104 B 0.025493f
C122 VDD1.n105 B 0.025493f
C123 VDD1.n106 B 0.01142f
C124 VDD1.n107 B 0.010785f
C125 VDD1.n108 B 0.020071f
C126 VDD1.n109 B 0.020071f
C127 VDD1.n110 B 0.010785f
C128 VDD1.n111 B 0.01142f
C129 VDD1.n112 B 0.025493f
C130 VDD1.n113 B 0.025493f
C131 VDD1.n114 B 0.01142f
C132 VDD1.n115 B 0.010785f
C133 VDD1.n116 B 0.020071f
C134 VDD1.n117 B 0.020071f
C135 VDD1.n118 B 0.010785f
C136 VDD1.n119 B 0.01142f
C137 VDD1.n120 B 0.025493f
C138 VDD1.n121 B 0.025493f
C139 VDD1.n122 B 0.01142f
C140 VDD1.n123 B 0.010785f
C141 VDD1.n124 B 0.020071f
C142 VDD1.n125 B 0.020071f
C143 VDD1.n126 B 0.010785f
C144 VDD1.n127 B 0.01142f
C145 VDD1.n128 B 0.025493f
C146 VDD1.n129 B 0.025493f
C147 VDD1.n130 B 0.01142f
C148 VDD1.n131 B 0.010785f
C149 VDD1.n132 B 0.020071f
C150 VDD1.n133 B 0.052425f
C151 VDD1.n134 B 0.010785f
C152 VDD1.n135 B 0.01142f
C153 VDD1.n136 B 0.052792f
C154 VDD1.n137 B 0.583123f
C155 VP.t1 B 2.94641f
C156 VP.t0 B 2.63832f
C157 VP.n0 B 4.57001f
C158 VDD2.n0 B 0.011431f
C159 VDD2.n1 B 0.025731f
C160 VDD2.n2 B 0.011526f
C161 VDD2.n3 B 0.020259f
C162 VDD2.n4 B 0.010886f
C163 VDD2.n5 B 0.025731f
C164 VDD2.n6 B 0.011526f
C165 VDD2.n7 B 0.020259f
C166 VDD2.n8 B 0.010886f
C167 VDD2.n9 B 0.025731f
C168 VDD2.n10 B 0.011526f
C169 VDD2.n11 B 0.020259f
C170 VDD2.n12 B 0.010886f
C171 VDD2.n13 B 0.025731f
C172 VDD2.n14 B 0.011526f
C173 VDD2.n15 B 0.020259f
C174 VDD2.n16 B 0.010886f
C175 VDD2.n17 B 0.025731f
C176 VDD2.n18 B 0.011526f
C177 VDD2.n19 B 0.020259f
C178 VDD2.n20 B 0.010886f
C179 VDD2.n21 B 0.019298f
C180 VDD2.n22 B 0.0152f
C181 VDD2.t1 B 0.042268f
C182 VDD2.n23 B 0.12045f
C183 VDD2.n24 B 1.10452f
C184 VDD2.n25 B 0.010886f
C185 VDD2.n26 B 0.011526f
C186 VDD2.n27 B 0.025731f
C187 VDD2.n28 B 0.025731f
C188 VDD2.n29 B 0.011526f
C189 VDD2.n30 B 0.010886f
C190 VDD2.n31 B 0.020259f
C191 VDD2.n32 B 0.020259f
C192 VDD2.n33 B 0.010886f
C193 VDD2.n34 B 0.011526f
C194 VDD2.n35 B 0.025731f
C195 VDD2.n36 B 0.025731f
C196 VDD2.n37 B 0.011526f
C197 VDD2.n38 B 0.010886f
C198 VDD2.n39 B 0.020259f
C199 VDD2.n40 B 0.020259f
C200 VDD2.n41 B 0.010886f
C201 VDD2.n42 B 0.011526f
C202 VDD2.n43 B 0.025731f
C203 VDD2.n44 B 0.025731f
C204 VDD2.n45 B 0.011526f
C205 VDD2.n46 B 0.010886f
C206 VDD2.n47 B 0.020259f
C207 VDD2.n48 B 0.020259f
C208 VDD2.n49 B 0.010886f
C209 VDD2.n50 B 0.011526f
C210 VDD2.n51 B 0.025731f
C211 VDD2.n52 B 0.025731f
C212 VDD2.n53 B 0.011526f
C213 VDD2.n54 B 0.010886f
C214 VDD2.n55 B 0.020259f
C215 VDD2.n56 B 0.020259f
C216 VDD2.n57 B 0.010886f
C217 VDD2.n58 B 0.011526f
C218 VDD2.n59 B 0.025731f
C219 VDD2.n60 B 0.025731f
C220 VDD2.n61 B 0.011526f
C221 VDD2.n62 B 0.010886f
C222 VDD2.n63 B 0.020259f
C223 VDD2.n64 B 0.052916f
C224 VDD2.n65 B 0.010886f
C225 VDD2.n66 B 0.011526f
C226 VDD2.n67 B 0.053286f
C227 VDD2.n68 B 0.556437f
C228 VDD2.n69 B 0.011431f
C229 VDD2.n70 B 0.025731f
C230 VDD2.n71 B 0.011526f
C231 VDD2.n72 B 0.020259f
C232 VDD2.n73 B 0.010886f
C233 VDD2.n74 B 0.025731f
C234 VDD2.n75 B 0.011526f
C235 VDD2.n76 B 0.020259f
C236 VDD2.n77 B 0.010886f
C237 VDD2.n78 B 0.025731f
C238 VDD2.n79 B 0.011526f
C239 VDD2.n80 B 0.020259f
C240 VDD2.n81 B 0.010886f
C241 VDD2.n82 B 0.025731f
C242 VDD2.n83 B 0.011526f
C243 VDD2.n84 B 0.020259f
C244 VDD2.n85 B 0.010886f
C245 VDD2.n86 B 0.025731f
C246 VDD2.n87 B 0.011526f
C247 VDD2.n88 B 0.020259f
C248 VDD2.n89 B 0.010886f
C249 VDD2.n90 B 0.019298f
C250 VDD2.n91 B 0.0152f
C251 VDD2.t0 B 0.042268f
C252 VDD2.n92 B 0.12045f
C253 VDD2.n93 B 1.10452f
C254 VDD2.n94 B 0.010886f
C255 VDD2.n95 B 0.011526f
C256 VDD2.n96 B 0.025731f
C257 VDD2.n97 B 0.025731f
C258 VDD2.n98 B 0.011526f
C259 VDD2.n99 B 0.010886f
C260 VDD2.n100 B 0.020259f
C261 VDD2.n101 B 0.020259f
C262 VDD2.n102 B 0.010886f
C263 VDD2.n103 B 0.011526f
C264 VDD2.n104 B 0.025731f
C265 VDD2.n105 B 0.025731f
C266 VDD2.n106 B 0.011526f
C267 VDD2.n107 B 0.010886f
C268 VDD2.n108 B 0.020259f
C269 VDD2.n109 B 0.020259f
C270 VDD2.n110 B 0.010886f
C271 VDD2.n111 B 0.011526f
C272 VDD2.n112 B 0.025731f
C273 VDD2.n113 B 0.025731f
C274 VDD2.n114 B 0.011526f
C275 VDD2.n115 B 0.010886f
C276 VDD2.n116 B 0.020259f
C277 VDD2.n117 B 0.020259f
C278 VDD2.n118 B 0.010886f
C279 VDD2.n119 B 0.011526f
C280 VDD2.n120 B 0.025731f
C281 VDD2.n121 B 0.025731f
C282 VDD2.n122 B 0.011526f
C283 VDD2.n123 B 0.010886f
C284 VDD2.n124 B 0.020259f
C285 VDD2.n125 B 0.020259f
C286 VDD2.n126 B 0.010886f
C287 VDD2.n127 B 0.011526f
C288 VDD2.n128 B 0.025731f
C289 VDD2.n129 B 0.025731f
C290 VDD2.n130 B 0.011526f
C291 VDD2.n131 B 0.010886f
C292 VDD2.n132 B 0.020259f
C293 VDD2.n133 B 0.052916f
C294 VDD2.n134 B 0.010886f
C295 VDD2.n135 B 0.011526f
C296 VDD2.n136 B 0.053286f
C297 VDD2.n137 B 0.059046f
C298 VDD2.n138 B 2.40317f
C299 VTAIL.n0 B 0.011425f
C300 VTAIL.n1 B 0.025717f
C301 VTAIL.n2 B 0.011521f
C302 VTAIL.n3 B 0.020248f
C303 VTAIL.n4 B 0.01088f
C304 VTAIL.n5 B 0.025717f
C305 VTAIL.n6 B 0.011521f
C306 VTAIL.n7 B 0.020248f
C307 VTAIL.n8 B 0.01088f
C308 VTAIL.n9 B 0.025717f
C309 VTAIL.n10 B 0.011521f
C310 VTAIL.n11 B 0.020248f
C311 VTAIL.n12 B 0.01088f
C312 VTAIL.n13 B 0.025717f
C313 VTAIL.n14 B 0.011521f
C314 VTAIL.n15 B 0.020248f
C315 VTAIL.n16 B 0.01088f
C316 VTAIL.n17 B 0.025717f
C317 VTAIL.n18 B 0.011521f
C318 VTAIL.n19 B 0.020248f
C319 VTAIL.n20 B 0.01088f
C320 VTAIL.n21 B 0.019288f
C321 VTAIL.n22 B 0.015192f
C322 VTAIL.t0 B 0.042245f
C323 VTAIL.n23 B 0.120386f
C324 VTAIL.n24 B 1.10394f
C325 VTAIL.n25 B 0.01088f
C326 VTAIL.n26 B 0.011521f
C327 VTAIL.n27 B 0.025717f
C328 VTAIL.n28 B 0.025717f
C329 VTAIL.n29 B 0.011521f
C330 VTAIL.n30 B 0.01088f
C331 VTAIL.n31 B 0.020248f
C332 VTAIL.n32 B 0.020248f
C333 VTAIL.n33 B 0.01088f
C334 VTAIL.n34 B 0.011521f
C335 VTAIL.n35 B 0.025717f
C336 VTAIL.n36 B 0.025717f
C337 VTAIL.n37 B 0.011521f
C338 VTAIL.n38 B 0.01088f
C339 VTAIL.n39 B 0.020248f
C340 VTAIL.n40 B 0.020248f
C341 VTAIL.n41 B 0.01088f
C342 VTAIL.n42 B 0.011521f
C343 VTAIL.n43 B 0.025717f
C344 VTAIL.n44 B 0.025717f
C345 VTAIL.n45 B 0.011521f
C346 VTAIL.n46 B 0.01088f
C347 VTAIL.n47 B 0.020248f
C348 VTAIL.n48 B 0.020248f
C349 VTAIL.n49 B 0.01088f
C350 VTAIL.n50 B 0.011521f
C351 VTAIL.n51 B 0.025717f
C352 VTAIL.n52 B 0.025717f
C353 VTAIL.n53 B 0.011521f
C354 VTAIL.n54 B 0.01088f
C355 VTAIL.n55 B 0.020248f
C356 VTAIL.n56 B 0.020248f
C357 VTAIL.n57 B 0.01088f
C358 VTAIL.n58 B 0.011521f
C359 VTAIL.n59 B 0.025717f
C360 VTAIL.n60 B 0.025717f
C361 VTAIL.n61 B 0.011521f
C362 VTAIL.n62 B 0.01088f
C363 VTAIL.n63 B 0.020248f
C364 VTAIL.n64 B 0.052888f
C365 VTAIL.n65 B 0.01088f
C366 VTAIL.n66 B 0.011521f
C367 VTAIL.n67 B 0.053258f
C368 VTAIL.n68 B 0.045072f
C369 VTAIL.n69 B 1.28974f
C370 VTAIL.n70 B 0.011425f
C371 VTAIL.n71 B 0.025717f
C372 VTAIL.n72 B 0.011521f
C373 VTAIL.n73 B 0.020248f
C374 VTAIL.n74 B 0.01088f
C375 VTAIL.n75 B 0.025717f
C376 VTAIL.n76 B 0.011521f
C377 VTAIL.n77 B 0.020248f
C378 VTAIL.n78 B 0.01088f
C379 VTAIL.n79 B 0.025717f
C380 VTAIL.n80 B 0.011521f
C381 VTAIL.n81 B 0.020248f
C382 VTAIL.n82 B 0.01088f
C383 VTAIL.n83 B 0.025717f
C384 VTAIL.n84 B 0.011521f
C385 VTAIL.n85 B 0.020248f
C386 VTAIL.n86 B 0.01088f
C387 VTAIL.n87 B 0.025717f
C388 VTAIL.n88 B 0.011521f
C389 VTAIL.n89 B 0.020248f
C390 VTAIL.n90 B 0.01088f
C391 VTAIL.n91 B 0.019288f
C392 VTAIL.n92 B 0.015192f
C393 VTAIL.t3 B 0.042245f
C394 VTAIL.n93 B 0.120386f
C395 VTAIL.n94 B 1.10394f
C396 VTAIL.n95 B 0.01088f
C397 VTAIL.n96 B 0.011521f
C398 VTAIL.n97 B 0.025717f
C399 VTAIL.n98 B 0.025717f
C400 VTAIL.n99 B 0.011521f
C401 VTAIL.n100 B 0.01088f
C402 VTAIL.n101 B 0.020248f
C403 VTAIL.n102 B 0.020248f
C404 VTAIL.n103 B 0.01088f
C405 VTAIL.n104 B 0.011521f
C406 VTAIL.n105 B 0.025717f
C407 VTAIL.n106 B 0.025717f
C408 VTAIL.n107 B 0.011521f
C409 VTAIL.n108 B 0.01088f
C410 VTAIL.n109 B 0.020248f
C411 VTAIL.n110 B 0.020248f
C412 VTAIL.n111 B 0.01088f
C413 VTAIL.n112 B 0.011521f
C414 VTAIL.n113 B 0.025717f
C415 VTAIL.n114 B 0.025717f
C416 VTAIL.n115 B 0.011521f
C417 VTAIL.n116 B 0.01088f
C418 VTAIL.n117 B 0.020248f
C419 VTAIL.n118 B 0.020248f
C420 VTAIL.n119 B 0.01088f
C421 VTAIL.n120 B 0.011521f
C422 VTAIL.n121 B 0.025717f
C423 VTAIL.n122 B 0.025717f
C424 VTAIL.n123 B 0.011521f
C425 VTAIL.n124 B 0.01088f
C426 VTAIL.n125 B 0.020248f
C427 VTAIL.n126 B 0.020248f
C428 VTAIL.n127 B 0.01088f
C429 VTAIL.n128 B 0.011521f
C430 VTAIL.n129 B 0.025717f
C431 VTAIL.n130 B 0.025717f
C432 VTAIL.n131 B 0.011521f
C433 VTAIL.n132 B 0.01088f
C434 VTAIL.n133 B 0.020248f
C435 VTAIL.n134 B 0.052888f
C436 VTAIL.n135 B 0.01088f
C437 VTAIL.n136 B 0.011521f
C438 VTAIL.n137 B 0.053258f
C439 VTAIL.n138 B 0.045072f
C440 VTAIL.n139 B 1.31322f
C441 VTAIL.n140 B 0.011425f
C442 VTAIL.n141 B 0.025717f
C443 VTAIL.n142 B 0.011521f
C444 VTAIL.n143 B 0.020248f
C445 VTAIL.n144 B 0.01088f
C446 VTAIL.n145 B 0.025717f
C447 VTAIL.n146 B 0.011521f
C448 VTAIL.n147 B 0.020248f
C449 VTAIL.n148 B 0.01088f
C450 VTAIL.n149 B 0.025717f
C451 VTAIL.n150 B 0.011521f
C452 VTAIL.n151 B 0.020248f
C453 VTAIL.n152 B 0.01088f
C454 VTAIL.n153 B 0.025717f
C455 VTAIL.n154 B 0.011521f
C456 VTAIL.n155 B 0.020248f
C457 VTAIL.n156 B 0.01088f
C458 VTAIL.n157 B 0.025717f
C459 VTAIL.n158 B 0.011521f
C460 VTAIL.n159 B 0.020248f
C461 VTAIL.n160 B 0.01088f
C462 VTAIL.n161 B 0.019288f
C463 VTAIL.n162 B 0.015192f
C464 VTAIL.t1 B 0.042245f
C465 VTAIL.n163 B 0.120386f
C466 VTAIL.n164 B 1.10394f
C467 VTAIL.n165 B 0.01088f
C468 VTAIL.n166 B 0.011521f
C469 VTAIL.n167 B 0.025717f
C470 VTAIL.n168 B 0.025717f
C471 VTAIL.n169 B 0.011521f
C472 VTAIL.n170 B 0.01088f
C473 VTAIL.n171 B 0.020248f
C474 VTAIL.n172 B 0.020248f
C475 VTAIL.n173 B 0.01088f
C476 VTAIL.n174 B 0.011521f
C477 VTAIL.n175 B 0.025717f
C478 VTAIL.n176 B 0.025717f
C479 VTAIL.n177 B 0.011521f
C480 VTAIL.n178 B 0.01088f
C481 VTAIL.n179 B 0.020248f
C482 VTAIL.n180 B 0.020248f
C483 VTAIL.n181 B 0.01088f
C484 VTAIL.n182 B 0.011521f
C485 VTAIL.n183 B 0.025717f
C486 VTAIL.n184 B 0.025717f
C487 VTAIL.n185 B 0.011521f
C488 VTAIL.n186 B 0.01088f
C489 VTAIL.n187 B 0.020248f
C490 VTAIL.n188 B 0.020248f
C491 VTAIL.n189 B 0.01088f
C492 VTAIL.n190 B 0.011521f
C493 VTAIL.n191 B 0.025717f
C494 VTAIL.n192 B 0.025717f
C495 VTAIL.n193 B 0.011521f
C496 VTAIL.n194 B 0.01088f
C497 VTAIL.n195 B 0.020248f
C498 VTAIL.n196 B 0.020248f
C499 VTAIL.n197 B 0.01088f
C500 VTAIL.n198 B 0.011521f
C501 VTAIL.n199 B 0.025717f
C502 VTAIL.n200 B 0.025717f
C503 VTAIL.n201 B 0.011521f
C504 VTAIL.n202 B 0.01088f
C505 VTAIL.n203 B 0.020248f
C506 VTAIL.n204 B 0.052888f
C507 VTAIL.n205 B 0.01088f
C508 VTAIL.n206 B 0.011521f
C509 VTAIL.n207 B 0.053258f
C510 VTAIL.n208 B 0.045072f
C511 VTAIL.n209 B 1.2041f
C512 VTAIL.n210 B 0.011425f
C513 VTAIL.n211 B 0.025717f
C514 VTAIL.n212 B 0.011521f
C515 VTAIL.n213 B 0.020248f
C516 VTAIL.n214 B 0.01088f
C517 VTAIL.n215 B 0.025717f
C518 VTAIL.n216 B 0.011521f
C519 VTAIL.n217 B 0.020248f
C520 VTAIL.n218 B 0.01088f
C521 VTAIL.n219 B 0.025717f
C522 VTAIL.n220 B 0.011521f
C523 VTAIL.n221 B 0.020248f
C524 VTAIL.n222 B 0.01088f
C525 VTAIL.n223 B 0.025717f
C526 VTAIL.n224 B 0.011521f
C527 VTAIL.n225 B 0.020248f
C528 VTAIL.n226 B 0.01088f
C529 VTAIL.n227 B 0.025717f
C530 VTAIL.n228 B 0.011521f
C531 VTAIL.n229 B 0.020248f
C532 VTAIL.n230 B 0.01088f
C533 VTAIL.n231 B 0.019288f
C534 VTAIL.n232 B 0.015192f
C535 VTAIL.t2 B 0.042245f
C536 VTAIL.n233 B 0.120386f
C537 VTAIL.n234 B 1.10394f
C538 VTAIL.n235 B 0.01088f
C539 VTAIL.n236 B 0.011521f
C540 VTAIL.n237 B 0.025717f
C541 VTAIL.n238 B 0.025717f
C542 VTAIL.n239 B 0.011521f
C543 VTAIL.n240 B 0.01088f
C544 VTAIL.n241 B 0.020248f
C545 VTAIL.n242 B 0.020248f
C546 VTAIL.n243 B 0.01088f
C547 VTAIL.n244 B 0.011521f
C548 VTAIL.n245 B 0.025717f
C549 VTAIL.n246 B 0.025717f
C550 VTAIL.n247 B 0.011521f
C551 VTAIL.n248 B 0.01088f
C552 VTAIL.n249 B 0.020248f
C553 VTAIL.n250 B 0.020248f
C554 VTAIL.n251 B 0.01088f
C555 VTAIL.n252 B 0.011521f
C556 VTAIL.n253 B 0.025717f
C557 VTAIL.n254 B 0.025717f
C558 VTAIL.n255 B 0.011521f
C559 VTAIL.n256 B 0.01088f
C560 VTAIL.n257 B 0.020248f
C561 VTAIL.n258 B 0.020248f
C562 VTAIL.n259 B 0.01088f
C563 VTAIL.n260 B 0.011521f
C564 VTAIL.n261 B 0.025717f
C565 VTAIL.n262 B 0.025717f
C566 VTAIL.n263 B 0.011521f
C567 VTAIL.n264 B 0.01088f
C568 VTAIL.n265 B 0.020248f
C569 VTAIL.n266 B 0.020248f
C570 VTAIL.n267 B 0.01088f
C571 VTAIL.n268 B 0.011521f
C572 VTAIL.n269 B 0.025717f
C573 VTAIL.n270 B 0.025717f
C574 VTAIL.n271 B 0.011521f
C575 VTAIL.n272 B 0.01088f
C576 VTAIL.n273 B 0.020248f
C577 VTAIL.n274 B 0.052888f
C578 VTAIL.n275 B 0.01088f
C579 VTAIL.n276 B 0.011521f
C580 VTAIL.n277 B 0.053258f
C581 VTAIL.n278 B 0.045072f
C582 VTAIL.n279 B 1.14238f
C583 VN.t0 B 2.57243f
C584 VN.t1 B 2.87702f
.ends

