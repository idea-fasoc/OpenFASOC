* NGSPICE file created from diff_pair_sample_0906.ext - technology: sky130A

.subckt diff_pair_sample_0906 VTAIL VN VP B VDD2 VDD1
X0 B.t23 B.t21 B.t22 B.t18 sky130_fd_pr__nfet_01v8 ad=2.6793 pd=14.52 as=0 ps=0 w=6.87 l=1.16
X1 VDD1.t9 VP.t0 VTAIL.t10 B.t3 sky130_fd_pr__nfet_01v8 ad=1.13355 pd=7.2 as=1.13355 ps=7.2 w=6.87 l=1.16
X2 B.t20 B.t17 B.t19 B.t18 sky130_fd_pr__nfet_01v8 ad=2.6793 pd=14.52 as=0 ps=0 w=6.87 l=1.16
X3 VDD2.t9 VN.t0 VTAIL.t9 B.t7 sky130_fd_pr__nfet_01v8 ad=1.13355 pd=7.2 as=1.13355 ps=7.2 w=6.87 l=1.16
X4 VDD2.t8 VN.t1 VTAIL.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=1.13355 pd=7.2 as=1.13355 ps=7.2 w=6.87 l=1.16
X5 VTAIL.t12 VP.t1 VDD1.t8 B.t5 sky130_fd_pr__nfet_01v8 ad=1.13355 pd=7.2 as=1.13355 ps=7.2 w=6.87 l=1.16
X6 VDD2.t7 VN.t2 VTAIL.t8 B.t9 sky130_fd_pr__nfet_01v8 ad=2.6793 pd=14.52 as=1.13355 ps=7.2 w=6.87 l=1.16
X7 VTAIL.t0 VN.t3 VDD2.t6 B.t0 sky130_fd_pr__nfet_01v8 ad=1.13355 pd=7.2 as=1.13355 ps=7.2 w=6.87 l=1.16
X8 VDD1.t7 VP.t2 VTAIL.t19 B.t7 sky130_fd_pr__nfet_01v8 ad=1.13355 pd=7.2 as=1.13355 ps=7.2 w=6.87 l=1.16
X9 VDD1.t6 VP.t3 VTAIL.t16 B.t4 sky130_fd_pr__nfet_01v8 ad=1.13355 pd=7.2 as=2.6793 ps=14.52 w=6.87 l=1.16
X10 VTAIL.t3 VN.t4 VDD2.t5 B.t6 sky130_fd_pr__nfet_01v8 ad=1.13355 pd=7.2 as=1.13355 ps=7.2 w=6.87 l=1.16
X11 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=2.6793 pd=14.52 as=0 ps=0 w=6.87 l=1.16
X12 VDD1.t5 VP.t4 VTAIL.t18 B.t1 sky130_fd_pr__nfet_01v8 ad=1.13355 pd=7.2 as=2.6793 ps=14.52 w=6.87 l=1.16
X13 VDD1.t4 VP.t5 VTAIL.t17 B.t9 sky130_fd_pr__nfet_01v8 ad=2.6793 pd=14.52 as=1.13355 ps=7.2 w=6.87 l=1.16
X14 VTAIL.t11 VP.t6 VDD1.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=1.13355 pd=7.2 as=1.13355 ps=7.2 w=6.87 l=1.16
X15 VTAIL.t2 VN.t5 VDD2.t4 B.t5 sky130_fd_pr__nfet_01v8 ad=1.13355 pd=7.2 as=1.13355 ps=7.2 w=6.87 l=1.16
X16 VDD2.t3 VN.t6 VTAIL.t7 B.t1 sky130_fd_pr__nfet_01v8 ad=1.13355 pd=7.2 as=2.6793 ps=14.52 w=6.87 l=1.16
X17 VTAIL.t14 VP.t7 VDD1.t2 B.t6 sky130_fd_pr__nfet_01v8 ad=1.13355 pd=7.2 as=1.13355 ps=7.2 w=6.87 l=1.16
X18 VDD2.t2 VN.t7 VTAIL.t6 B.t8 sky130_fd_pr__nfet_01v8 ad=2.6793 pd=14.52 as=1.13355 ps=7.2 w=6.87 l=1.16
X19 VDD2.t1 VN.t8 VTAIL.t1 B.t4 sky130_fd_pr__nfet_01v8 ad=1.13355 pd=7.2 as=2.6793 ps=14.52 w=6.87 l=1.16
X20 VTAIL.t13 VP.t8 VDD1.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=1.13355 pd=7.2 as=1.13355 ps=7.2 w=6.87 l=1.16
X21 VDD1.t0 VP.t9 VTAIL.t15 B.t8 sky130_fd_pr__nfet_01v8 ad=2.6793 pd=14.52 as=1.13355 ps=7.2 w=6.87 l=1.16
X22 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=2.6793 pd=14.52 as=0 ps=0 w=6.87 l=1.16
X23 VTAIL.t5 VN.t9 VDD2.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=1.13355 pd=7.2 as=1.13355 ps=7.2 w=6.87 l=1.16
R0 B.n479 B.n478 585
R1 B.n479 B.n64 585
R2 B.n482 B.n481 585
R3 B.n483 B.n100 585
R4 B.n485 B.n484 585
R5 B.n487 B.n99 585
R6 B.n490 B.n489 585
R7 B.n491 B.n98 585
R8 B.n493 B.n492 585
R9 B.n495 B.n97 585
R10 B.n498 B.n497 585
R11 B.n499 B.n96 585
R12 B.n501 B.n500 585
R13 B.n503 B.n95 585
R14 B.n506 B.n505 585
R15 B.n507 B.n94 585
R16 B.n509 B.n508 585
R17 B.n511 B.n93 585
R18 B.n514 B.n513 585
R19 B.n515 B.n92 585
R20 B.n517 B.n516 585
R21 B.n519 B.n91 585
R22 B.n522 B.n521 585
R23 B.n523 B.n90 585
R24 B.n525 B.n524 585
R25 B.n527 B.n89 585
R26 B.n530 B.n529 585
R27 B.n531 B.n86 585
R28 B.n534 B.n533 585
R29 B.n536 B.n85 585
R30 B.n539 B.n538 585
R31 B.n540 B.n84 585
R32 B.n542 B.n541 585
R33 B.n544 B.n83 585
R34 B.n547 B.n546 585
R35 B.n548 B.n79 585
R36 B.n550 B.n549 585
R37 B.n552 B.n78 585
R38 B.n555 B.n554 585
R39 B.n556 B.n77 585
R40 B.n558 B.n557 585
R41 B.n560 B.n76 585
R42 B.n563 B.n562 585
R43 B.n564 B.n75 585
R44 B.n566 B.n565 585
R45 B.n568 B.n74 585
R46 B.n571 B.n570 585
R47 B.n572 B.n73 585
R48 B.n574 B.n573 585
R49 B.n576 B.n72 585
R50 B.n579 B.n578 585
R51 B.n580 B.n71 585
R52 B.n582 B.n581 585
R53 B.n584 B.n70 585
R54 B.n587 B.n586 585
R55 B.n588 B.n69 585
R56 B.n590 B.n589 585
R57 B.n592 B.n68 585
R58 B.n595 B.n594 585
R59 B.n596 B.n67 585
R60 B.n598 B.n597 585
R61 B.n600 B.n66 585
R62 B.n603 B.n602 585
R63 B.n604 B.n65 585
R64 B.n477 B.n63 585
R65 B.n607 B.n63 585
R66 B.n476 B.n62 585
R67 B.n608 B.n62 585
R68 B.n475 B.n61 585
R69 B.n609 B.n61 585
R70 B.n474 B.n473 585
R71 B.n473 B.n57 585
R72 B.n472 B.n56 585
R73 B.n615 B.n56 585
R74 B.n471 B.n55 585
R75 B.n616 B.n55 585
R76 B.n470 B.n54 585
R77 B.n617 B.n54 585
R78 B.n469 B.n468 585
R79 B.n468 B.n50 585
R80 B.n467 B.n49 585
R81 B.n623 B.n49 585
R82 B.n466 B.n48 585
R83 B.n624 B.n48 585
R84 B.n465 B.n47 585
R85 B.n625 B.n47 585
R86 B.n464 B.n463 585
R87 B.n463 B.n43 585
R88 B.n462 B.n42 585
R89 B.n631 B.n42 585
R90 B.n461 B.n41 585
R91 B.n632 B.n41 585
R92 B.n460 B.n40 585
R93 B.n633 B.n40 585
R94 B.n459 B.n458 585
R95 B.n458 B.n36 585
R96 B.n457 B.n35 585
R97 B.n639 B.n35 585
R98 B.n456 B.n34 585
R99 B.n640 B.n34 585
R100 B.n455 B.n33 585
R101 B.n641 B.n33 585
R102 B.n454 B.n453 585
R103 B.n453 B.n29 585
R104 B.n452 B.n28 585
R105 B.n647 B.n28 585
R106 B.n451 B.n27 585
R107 B.n648 B.n27 585
R108 B.n450 B.n26 585
R109 B.n649 B.n26 585
R110 B.n449 B.n448 585
R111 B.n448 B.n22 585
R112 B.n447 B.n21 585
R113 B.n655 B.n21 585
R114 B.n446 B.n20 585
R115 B.n656 B.n20 585
R116 B.n445 B.n19 585
R117 B.n657 B.n19 585
R118 B.n444 B.n443 585
R119 B.n443 B.n15 585
R120 B.n442 B.n14 585
R121 B.n663 B.n14 585
R122 B.n441 B.n13 585
R123 B.n664 B.n13 585
R124 B.n440 B.n12 585
R125 B.n665 B.n12 585
R126 B.n439 B.n438 585
R127 B.n438 B.n437 585
R128 B.n436 B.n435 585
R129 B.n436 B.n8 585
R130 B.n434 B.n7 585
R131 B.n672 B.n7 585
R132 B.n433 B.n6 585
R133 B.n673 B.n6 585
R134 B.n432 B.n5 585
R135 B.n674 B.n5 585
R136 B.n431 B.n430 585
R137 B.n430 B.n4 585
R138 B.n429 B.n101 585
R139 B.n429 B.n428 585
R140 B.n419 B.n102 585
R141 B.n103 B.n102 585
R142 B.n421 B.n420 585
R143 B.n422 B.n421 585
R144 B.n418 B.n108 585
R145 B.n108 B.n107 585
R146 B.n417 B.n416 585
R147 B.n416 B.n415 585
R148 B.n110 B.n109 585
R149 B.n111 B.n110 585
R150 B.n408 B.n407 585
R151 B.n409 B.n408 585
R152 B.n406 B.n116 585
R153 B.n116 B.n115 585
R154 B.n405 B.n404 585
R155 B.n404 B.n403 585
R156 B.n118 B.n117 585
R157 B.n119 B.n118 585
R158 B.n396 B.n395 585
R159 B.n397 B.n396 585
R160 B.n394 B.n123 585
R161 B.n127 B.n123 585
R162 B.n393 B.n392 585
R163 B.n392 B.n391 585
R164 B.n125 B.n124 585
R165 B.n126 B.n125 585
R166 B.n384 B.n383 585
R167 B.n385 B.n384 585
R168 B.n382 B.n131 585
R169 B.n135 B.n131 585
R170 B.n381 B.n380 585
R171 B.n380 B.n379 585
R172 B.n133 B.n132 585
R173 B.n134 B.n133 585
R174 B.n372 B.n371 585
R175 B.n373 B.n372 585
R176 B.n370 B.n139 585
R177 B.n143 B.n139 585
R178 B.n369 B.n368 585
R179 B.n368 B.n367 585
R180 B.n141 B.n140 585
R181 B.n142 B.n141 585
R182 B.n360 B.n359 585
R183 B.n361 B.n360 585
R184 B.n358 B.n148 585
R185 B.n148 B.n147 585
R186 B.n357 B.n356 585
R187 B.n356 B.n355 585
R188 B.n150 B.n149 585
R189 B.n151 B.n150 585
R190 B.n348 B.n347 585
R191 B.n349 B.n348 585
R192 B.n346 B.n155 585
R193 B.n159 B.n155 585
R194 B.n345 B.n344 585
R195 B.n344 B.n343 585
R196 B.n157 B.n156 585
R197 B.n158 B.n157 585
R198 B.n336 B.n335 585
R199 B.n337 B.n336 585
R200 B.n334 B.n164 585
R201 B.n164 B.n163 585
R202 B.n333 B.n332 585
R203 B.n332 B.n331 585
R204 B.n328 B.n168 585
R205 B.n327 B.n326 585
R206 B.n324 B.n169 585
R207 B.n324 B.n167 585
R208 B.n323 B.n322 585
R209 B.n321 B.n320 585
R210 B.n319 B.n171 585
R211 B.n317 B.n316 585
R212 B.n315 B.n172 585
R213 B.n314 B.n313 585
R214 B.n311 B.n173 585
R215 B.n309 B.n308 585
R216 B.n307 B.n174 585
R217 B.n306 B.n305 585
R218 B.n303 B.n175 585
R219 B.n301 B.n300 585
R220 B.n299 B.n176 585
R221 B.n298 B.n297 585
R222 B.n295 B.n177 585
R223 B.n293 B.n292 585
R224 B.n291 B.n178 585
R225 B.n290 B.n289 585
R226 B.n287 B.n179 585
R227 B.n285 B.n284 585
R228 B.n283 B.n180 585
R229 B.n282 B.n281 585
R230 B.n279 B.n181 585
R231 B.n277 B.n276 585
R232 B.n274 B.n182 585
R233 B.n273 B.n272 585
R234 B.n270 B.n185 585
R235 B.n268 B.n267 585
R236 B.n266 B.n186 585
R237 B.n265 B.n264 585
R238 B.n262 B.n187 585
R239 B.n260 B.n259 585
R240 B.n258 B.n188 585
R241 B.n256 B.n255 585
R242 B.n253 B.n191 585
R243 B.n251 B.n250 585
R244 B.n249 B.n192 585
R245 B.n248 B.n247 585
R246 B.n245 B.n193 585
R247 B.n243 B.n242 585
R248 B.n241 B.n194 585
R249 B.n240 B.n239 585
R250 B.n237 B.n195 585
R251 B.n235 B.n234 585
R252 B.n233 B.n196 585
R253 B.n232 B.n231 585
R254 B.n229 B.n197 585
R255 B.n227 B.n226 585
R256 B.n225 B.n198 585
R257 B.n224 B.n223 585
R258 B.n221 B.n199 585
R259 B.n219 B.n218 585
R260 B.n217 B.n200 585
R261 B.n216 B.n215 585
R262 B.n213 B.n201 585
R263 B.n211 B.n210 585
R264 B.n209 B.n202 585
R265 B.n208 B.n207 585
R266 B.n205 B.n203 585
R267 B.n166 B.n165 585
R268 B.n330 B.n329 585
R269 B.n331 B.n330 585
R270 B.n162 B.n161 585
R271 B.n163 B.n162 585
R272 B.n339 B.n338 585
R273 B.n338 B.n337 585
R274 B.n340 B.n160 585
R275 B.n160 B.n158 585
R276 B.n342 B.n341 585
R277 B.n343 B.n342 585
R278 B.n154 B.n153 585
R279 B.n159 B.n154 585
R280 B.n351 B.n350 585
R281 B.n350 B.n349 585
R282 B.n352 B.n152 585
R283 B.n152 B.n151 585
R284 B.n354 B.n353 585
R285 B.n355 B.n354 585
R286 B.n146 B.n145 585
R287 B.n147 B.n146 585
R288 B.n363 B.n362 585
R289 B.n362 B.n361 585
R290 B.n364 B.n144 585
R291 B.n144 B.n142 585
R292 B.n366 B.n365 585
R293 B.n367 B.n366 585
R294 B.n138 B.n137 585
R295 B.n143 B.n138 585
R296 B.n375 B.n374 585
R297 B.n374 B.n373 585
R298 B.n376 B.n136 585
R299 B.n136 B.n134 585
R300 B.n378 B.n377 585
R301 B.n379 B.n378 585
R302 B.n130 B.n129 585
R303 B.n135 B.n130 585
R304 B.n387 B.n386 585
R305 B.n386 B.n385 585
R306 B.n388 B.n128 585
R307 B.n128 B.n126 585
R308 B.n390 B.n389 585
R309 B.n391 B.n390 585
R310 B.n122 B.n121 585
R311 B.n127 B.n122 585
R312 B.n399 B.n398 585
R313 B.n398 B.n397 585
R314 B.n400 B.n120 585
R315 B.n120 B.n119 585
R316 B.n402 B.n401 585
R317 B.n403 B.n402 585
R318 B.n114 B.n113 585
R319 B.n115 B.n114 585
R320 B.n411 B.n410 585
R321 B.n410 B.n409 585
R322 B.n412 B.n112 585
R323 B.n112 B.n111 585
R324 B.n414 B.n413 585
R325 B.n415 B.n414 585
R326 B.n106 B.n105 585
R327 B.n107 B.n106 585
R328 B.n424 B.n423 585
R329 B.n423 B.n422 585
R330 B.n425 B.n104 585
R331 B.n104 B.n103 585
R332 B.n427 B.n426 585
R333 B.n428 B.n427 585
R334 B.n3 B.n0 585
R335 B.n4 B.n3 585
R336 B.n671 B.n1 585
R337 B.n672 B.n671 585
R338 B.n670 B.n669 585
R339 B.n670 B.n8 585
R340 B.n668 B.n9 585
R341 B.n437 B.n9 585
R342 B.n667 B.n666 585
R343 B.n666 B.n665 585
R344 B.n11 B.n10 585
R345 B.n664 B.n11 585
R346 B.n662 B.n661 585
R347 B.n663 B.n662 585
R348 B.n660 B.n16 585
R349 B.n16 B.n15 585
R350 B.n659 B.n658 585
R351 B.n658 B.n657 585
R352 B.n18 B.n17 585
R353 B.n656 B.n18 585
R354 B.n654 B.n653 585
R355 B.n655 B.n654 585
R356 B.n652 B.n23 585
R357 B.n23 B.n22 585
R358 B.n651 B.n650 585
R359 B.n650 B.n649 585
R360 B.n25 B.n24 585
R361 B.n648 B.n25 585
R362 B.n646 B.n645 585
R363 B.n647 B.n646 585
R364 B.n644 B.n30 585
R365 B.n30 B.n29 585
R366 B.n643 B.n642 585
R367 B.n642 B.n641 585
R368 B.n32 B.n31 585
R369 B.n640 B.n32 585
R370 B.n638 B.n637 585
R371 B.n639 B.n638 585
R372 B.n636 B.n37 585
R373 B.n37 B.n36 585
R374 B.n635 B.n634 585
R375 B.n634 B.n633 585
R376 B.n39 B.n38 585
R377 B.n632 B.n39 585
R378 B.n630 B.n629 585
R379 B.n631 B.n630 585
R380 B.n628 B.n44 585
R381 B.n44 B.n43 585
R382 B.n627 B.n626 585
R383 B.n626 B.n625 585
R384 B.n46 B.n45 585
R385 B.n624 B.n46 585
R386 B.n622 B.n621 585
R387 B.n623 B.n622 585
R388 B.n620 B.n51 585
R389 B.n51 B.n50 585
R390 B.n619 B.n618 585
R391 B.n618 B.n617 585
R392 B.n53 B.n52 585
R393 B.n616 B.n53 585
R394 B.n614 B.n613 585
R395 B.n615 B.n614 585
R396 B.n612 B.n58 585
R397 B.n58 B.n57 585
R398 B.n611 B.n610 585
R399 B.n610 B.n609 585
R400 B.n60 B.n59 585
R401 B.n608 B.n60 585
R402 B.n606 B.n605 585
R403 B.n607 B.n606 585
R404 B.n675 B.n674 585
R405 B.n673 B.n2 585
R406 B.n606 B.n65 454.062
R407 B.n479 B.n63 454.062
R408 B.n332 B.n166 454.062
R409 B.n330 B.n168 454.062
R410 B.n80 B.t14 346.632
R411 B.n87 B.t10 346.632
R412 B.n189 B.t17 346.632
R413 B.n183 B.t21 346.632
R414 B.n480 B.n64 256.663
R415 B.n486 B.n64 256.663
R416 B.n488 B.n64 256.663
R417 B.n494 B.n64 256.663
R418 B.n496 B.n64 256.663
R419 B.n502 B.n64 256.663
R420 B.n504 B.n64 256.663
R421 B.n510 B.n64 256.663
R422 B.n512 B.n64 256.663
R423 B.n518 B.n64 256.663
R424 B.n520 B.n64 256.663
R425 B.n526 B.n64 256.663
R426 B.n528 B.n64 256.663
R427 B.n535 B.n64 256.663
R428 B.n537 B.n64 256.663
R429 B.n543 B.n64 256.663
R430 B.n545 B.n64 256.663
R431 B.n551 B.n64 256.663
R432 B.n553 B.n64 256.663
R433 B.n559 B.n64 256.663
R434 B.n561 B.n64 256.663
R435 B.n567 B.n64 256.663
R436 B.n569 B.n64 256.663
R437 B.n575 B.n64 256.663
R438 B.n577 B.n64 256.663
R439 B.n583 B.n64 256.663
R440 B.n585 B.n64 256.663
R441 B.n591 B.n64 256.663
R442 B.n593 B.n64 256.663
R443 B.n599 B.n64 256.663
R444 B.n601 B.n64 256.663
R445 B.n325 B.n167 256.663
R446 B.n170 B.n167 256.663
R447 B.n318 B.n167 256.663
R448 B.n312 B.n167 256.663
R449 B.n310 B.n167 256.663
R450 B.n304 B.n167 256.663
R451 B.n302 B.n167 256.663
R452 B.n296 B.n167 256.663
R453 B.n294 B.n167 256.663
R454 B.n288 B.n167 256.663
R455 B.n286 B.n167 256.663
R456 B.n280 B.n167 256.663
R457 B.n278 B.n167 256.663
R458 B.n271 B.n167 256.663
R459 B.n269 B.n167 256.663
R460 B.n263 B.n167 256.663
R461 B.n261 B.n167 256.663
R462 B.n254 B.n167 256.663
R463 B.n252 B.n167 256.663
R464 B.n246 B.n167 256.663
R465 B.n244 B.n167 256.663
R466 B.n238 B.n167 256.663
R467 B.n236 B.n167 256.663
R468 B.n230 B.n167 256.663
R469 B.n228 B.n167 256.663
R470 B.n222 B.n167 256.663
R471 B.n220 B.n167 256.663
R472 B.n214 B.n167 256.663
R473 B.n212 B.n167 256.663
R474 B.n206 B.n167 256.663
R475 B.n204 B.n167 256.663
R476 B.n677 B.n676 256.663
R477 B.n602 B.n600 163.367
R478 B.n598 B.n67 163.367
R479 B.n594 B.n592 163.367
R480 B.n590 B.n69 163.367
R481 B.n586 B.n584 163.367
R482 B.n582 B.n71 163.367
R483 B.n578 B.n576 163.367
R484 B.n574 B.n73 163.367
R485 B.n570 B.n568 163.367
R486 B.n566 B.n75 163.367
R487 B.n562 B.n560 163.367
R488 B.n558 B.n77 163.367
R489 B.n554 B.n552 163.367
R490 B.n550 B.n79 163.367
R491 B.n546 B.n544 163.367
R492 B.n542 B.n84 163.367
R493 B.n538 B.n536 163.367
R494 B.n534 B.n86 163.367
R495 B.n529 B.n527 163.367
R496 B.n525 B.n90 163.367
R497 B.n521 B.n519 163.367
R498 B.n517 B.n92 163.367
R499 B.n513 B.n511 163.367
R500 B.n509 B.n94 163.367
R501 B.n505 B.n503 163.367
R502 B.n501 B.n96 163.367
R503 B.n497 B.n495 163.367
R504 B.n493 B.n98 163.367
R505 B.n489 B.n487 163.367
R506 B.n485 B.n100 163.367
R507 B.n481 B.n479 163.367
R508 B.n332 B.n164 163.367
R509 B.n336 B.n164 163.367
R510 B.n336 B.n157 163.367
R511 B.n344 B.n157 163.367
R512 B.n344 B.n155 163.367
R513 B.n348 B.n155 163.367
R514 B.n348 B.n150 163.367
R515 B.n356 B.n150 163.367
R516 B.n356 B.n148 163.367
R517 B.n360 B.n148 163.367
R518 B.n360 B.n141 163.367
R519 B.n368 B.n141 163.367
R520 B.n368 B.n139 163.367
R521 B.n372 B.n139 163.367
R522 B.n372 B.n133 163.367
R523 B.n380 B.n133 163.367
R524 B.n380 B.n131 163.367
R525 B.n384 B.n131 163.367
R526 B.n384 B.n125 163.367
R527 B.n392 B.n125 163.367
R528 B.n392 B.n123 163.367
R529 B.n396 B.n123 163.367
R530 B.n396 B.n118 163.367
R531 B.n404 B.n118 163.367
R532 B.n404 B.n116 163.367
R533 B.n408 B.n116 163.367
R534 B.n408 B.n110 163.367
R535 B.n416 B.n110 163.367
R536 B.n416 B.n108 163.367
R537 B.n421 B.n108 163.367
R538 B.n421 B.n102 163.367
R539 B.n429 B.n102 163.367
R540 B.n430 B.n429 163.367
R541 B.n430 B.n5 163.367
R542 B.n6 B.n5 163.367
R543 B.n7 B.n6 163.367
R544 B.n436 B.n7 163.367
R545 B.n438 B.n436 163.367
R546 B.n438 B.n12 163.367
R547 B.n13 B.n12 163.367
R548 B.n14 B.n13 163.367
R549 B.n443 B.n14 163.367
R550 B.n443 B.n19 163.367
R551 B.n20 B.n19 163.367
R552 B.n21 B.n20 163.367
R553 B.n448 B.n21 163.367
R554 B.n448 B.n26 163.367
R555 B.n27 B.n26 163.367
R556 B.n28 B.n27 163.367
R557 B.n453 B.n28 163.367
R558 B.n453 B.n33 163.367
R559 B.n34 B.n33 163.367
R560 B.n35 B.n34 163.367
R561 B.n458 B.n35 163.367
R562 B.n458 B.n40 163.367
R563 B.n41 B.n40 163.367
R564 B.n42 B.n41 163.367
R565 B.n463 B.n42 163.367
R566 B.n463 B.n47 163.367
R567 B.n48 B.n47 163.367
R568 B.n49 B.n48 163.367
R569 B.n468 B.n49 163.367
R570 B.n468 B.n54 163.367
R571 B.n55 B.n54 163.367
R572 B.n56 B.n55 163.367
R573 B.n473 B.n56 163.367
R574 B.n473 B.n61 163.367
R575 B.n62 B.n61 163.367
R576 B.n63 B.n62 163.367
R577 B.n326 B.n324 163.367
R578 B.n324 B.n323 163.367
R579 B.n320 B.n319 163.367
R580 B.n317 B.n172 163.367
R581 B.n313 B.n311 163.367
R582 B.n309 B.n174 163.367
R583 B.n305 B.n303 163.367
R584 B.n301 B.n176 163.367
R585 B.n297 B.n295 163.367
R586 B.n293 B.n178 163.367
R587 B.n289 B.n287 163.367
R588 B.n285 B.n180 163.367
R589 B.n281 B.n279 163.367
R590 B.n277 B.n182 163.367
R591 B.n272 B.n270 163.367
R592 B.n268 B.n186 163.367
R593 B.n264 B.n262 163.367
R594 B.n260 B.n188 163.367
R595 B.n255 B.n253 163.367
R596 B.n251 B.n192 163.367
R597 B.n247 B.n245 163.367
R598 B.n243 B.n194 163.367
R599 B.n239 B.n237 163.367
R600 B.n235 B.n196 163.367
R601 B.n231 B.n229 163.367
R602 B.n227 B.n198 163.367
R603 B.n223 B.n221 163.367
R604 B.n219 B.n200 163.367
R605 B.n215 B.n213 163.367
R606 B.n211 B.n202 163.367
R607 B.n207 B.n205 163.367
R608 B.n330 B.n162 163.367
R609 B.n338 B.n162 163.367
R610 B.n338 B.n160 163.367
R611 B.n342 B.n160 163.367
R612 B.n342 B.n154 163.367
R613 B.n350 B.n154 163.367
R614 B.n350 B.n152 163.367
R615 B.n354 B.n152 163.367
R616 B.n354 B.n146 163.367
R617 B.n362 B.n146 163.367
R618 B.n362 B.n144 163.367
R619 B.n366 B.n144 163.367
R620 B.n366 B.n138 163.367
R621 B.n374 B.n138 163.367
R622 B.n374 B.n136 163.367
R623 B.n378 B.n136 163.367
R624 B.n378 B.n130 163.367
R625 B.n386 B.n130 163.367
R626 B.n386 B.n128 163.367
R627 B.n390 B.n128 163.367
R628 B.n390 B.n122 163.367
R629 B.n398 B.n122 163.367
R630 B.n398 B.n120 163.367
R631 B.n402 B.n120 163.367
R632 B.n402 B.n114 163.367
R633 B.n410 B.n114 163.367
R634 B.n410 B.n112 163.367
R635 B.n414 B.n112 163.367
R636 B.n414 B.n106 163.367
R637 B.n423 B.n106 163.367
R638 B.n423 B.n104 163.367
R639 B.n427 B.n104 163.367
R640 B.n427 B.n3 163.367
R641 B.n675 B.n3 163.367
R642 B.n671 B.n2 163.367
R643 B.n671 B.n670 163.367
R644 B.n670 B.n9 163.367
R645 B.n666 B.n9 163.367
R646 B.n666 B.n11 163.367
R647 B.n662 B.n11 163.367
R648 B.n662 B.n16 163.367
R649 B.n658 B.n16 163.367
R650 B.n658 B.n18 163.367
R651 B.n654 B.n18 163.367
R652 B.n654 B.n23 163.367
R653 B.n650 B.n23 163.367
R654 B.n650 B.n25 163.367
R655 B.n646 B.n25 163.367
R656 B.n646 B.n30 163.367
R657 B.n642 B.n30 163.367
R658 B.n642 B.n32 163.367
R659 B.n638 B.n32 163.367
R660 B.n638 B.n37 163.367
R661 B.n634 B.n37 163.367
R662 B.n634 B.n39 163.367
R663 B.n630 B.n39 163.367
R664 B.n630 B.n44 163.367
R665 B.n626 B.n44 163.367
R666 B.n626 B.n46 163.367
R667 B.n622 B.n46 163.367
R668 B.n622 B.n51 163.367
R669 B.n618 B.n51 163.367
R670 B.n618 B.n53 163.367
R671 B.n614 B.n53 163.367
R672 B.n614 B.n58 163.367
R673 B.n610 B.n58 163.367
R674 B.n610 B.n60 163.367
R675 B.n606 B.n60 163.367
R676 B.n331 B.n167 105.971
R677 B.n607 B.n64 105.971
R678 B.n87 B.t12 99.2731
R679 B.n189 B.t20 99.2731
R680 B.n80 B.t15 99.2653
R681 B.n183 B.t23 99.2653
R682 B.n601 B.n65 71.676
R683 B.n600 B.n599 71.676
R684 B.n593 B.n67 71.676
R685 B.n592 B.n591 71.676
R686 B.n585 B.n69 71.676
R687 B.n584 B.n583 71.676
R688 B.n577 B.n71 71.676
R689 B.n576 B.n575 71.676
R690 B.n569 B.n73 71.676
R691 B.n568 B.n567 71.676
R692 B.n561 B.n75 71.676
R693 B.n560 B.n559 71.676
R694 B.n553 B.n77 71.676
R695 B.n552 B.n551 71.676
R696 B.n545 B.n79 71.676
R697 B.n544 B.n543 71.676
R698 B.n537 B.n84 71.676
R699 B.n536 B.n535 71.676
R700 B.n528 B.n86 71.676
R701 B.n527 B.n526 71.676
R702 B.n520 B.n90 71.676
R703 B.n519 B.n518 71.676
R704 B.n512 B.n92 71.676
R705 B.n511 B.n510 71.676
R706 B.n504 B.n94 71.676
R707 B.n503 B.n502 71.676
R708 B.n496 B.n96 71.676
R709 B.n495 B.n494 71.676
R710 B.n488 B.n98 71.676
R711 B.n487 B.n486 71.676
R712 B.n480 B.n100 71.676
R713 B.n481 B.n480 71.676
R714 B.n486 B.n485 71.676
R715 B.n489 B.n488 71.676
R716 B.n494 B.n493 71.676
R717 B.n497 B.n496 71.676
R718 B.n502 B.n501 71.676
R719 B.n505 B.n504 71.676
R720 B.n510 B.n509 71.676
R721 B.n513 B.n512 71.676
R722 B.n518 B.n517 71.676
R723 B.n521 B.n520 71.676
R724 B.n526 B.n525 71.676
R725 B.n529 B.n528 71.676
R726 B.n535 B.n534 71.676
R727 B.n538 B.n537 71.676
R728 B.n543 B.n542 71.676
R729 B.n546 B.n545 71.676
R730 B.n551 B.n550 71.676
R731 B.n554 B.n553 71.676
R732 B.n559 B.n558 71.676
R733 B.n562 B.n561 71.676
R734 B.n567 B.n566 71.676
R735 B.n570 B.n569 71.676
R736 B.n575 B.n574 71.676
R737 B.n578 B.n577 71.676
R738 B.n583 B.n582 71.676
R739 B.n586 B.n585 71.676
R740 B.n591 B.n590 71.676
R741 B.n594 B.n593 71.676
R742 B.n599 B.n598 71.676
R743 B.n602 B.n601 71.676
R744 B.n325 B.n168 71.676
R745 B.n323 B.n170 71.676
R746 B.n319 B.n318 71.676
R747 B.n312 B.n172 71.676
R748 B.n311 B.n310 71.676
R749 B.n304 B.n174 71.676
R750 B.n303 B.n302 71.676
R751 B.n296 B.n176 71.676
R752 B.n295 B.n294 71.676
R753 B.n288 B.n178 71.676
R754 B.n287 B.n286 71.676
R755 B.n280 B.n180 71.676
R756 B.n279 B.n278 71.676
R757 B.n271 B.n182 71.676
R758 B.n270 B.n269 71.676
R759 B.n263 B.n186 71.676
R760 B.n262 B.n261 71.676
R761 B.n254 B.n188 71.676
R762 B.n253 B.n252 71.676
R763 B.n246 B.n192 71.676
R764 B.n245 B.n244 71.676
R765 B.n238 B.n194 71.676
R766 B.n237 B.n236 71.676
R767 B.n230 B.n196 71.676
R768 B.n229 B.n228 71.676
R769 B.n222 B.n198 71.676
R770 B.n221 B.n220 71.676
R771 B.n214 B.n200 71.676
R772 B.n213 B.n212 71.676
R773 B.n206 B.n202 71.676
R774 B.n205 B.n204 71.676
R775 B.n326 B.n325 71.676
R776 B.n320 B.n170 71.676
R777 B.n318 B.n317 71.676
R778 B.n313 B.n312 71.676
R779 B.n310 B.n309 71.676
R780 B.n305 B.n304 71.676
R781 B.n302 B.n301 71.676
R782 B.n297 B.n296 71.676
R783 B.n294 B.n293 71.676
R784 B.n289 B.n288 71.676
R785 B.n286 B.n285 71.676
R786 B.n281 B.n280 71.676
R787 B.n278 B.n277 71.676
R788 B.n272 B.n271 71.676
R789 B.n269 B.n268 71.676
R790 B.n264 B.n263 71.676
R791 B.n261 B.n260 71.676
R792 B.n255 B.n254 71.676
R793 B.n252 B.n251 71.676
R794 B.n247 B.n246 71.676
R795 B.n244 B.n243 71.676
R796 B.n239 B.n238 71.676
R797 B.n236 B.n235 71.676
R798 B.n231 B.n230 71.676
R799 B.n228 B.n227 71.676
R800 B.n223 B.n222 71.676
R801 B.n220 B.n219 71.676
R802 B.n215 B.n214 71.676
R803 B.n212 B.n211 71.676
R804 B.n207 B.n206 71.676
R805 B.n204 B.n166 71.676
R806 B.n676 B.n675 71.676
R807 B.n676 B.n2 71.676
R808 B.n88 B.t13 70.3761
R809 B.n190 B.t19 70.3761
R810 B.n81 B.t16 70.3684
R811 B.n184 B.t22 70.3684
R812 B.n331 B.n163 61.5896
R813 B.n337 B.n163 61.5896
R814 B.n337 B.n158 61.5896
R815 B.n343 B.n158 61.5896
R816 B.n343 B.n159 61.5896
R817 B.n349 B.n151 61.5896
R818 B.n355 B.n151 61.5896
R819 B.n355 B.n147 61.5896
R820 B.n361 B.n147 61.5896
R821 B.n361 B.n142 61.5896
R822 B.n367 B.n142 61.5896
R823 B.n367 B.n143 61.5896
R824 B.n373 B.n134 61.5896
R825 B.n379 B.n134 61.5896
R826 B.n379 B.n135 61.5896
R827 B.n385 B.n126 61.5896
R828 B.n391 B.n126 61.5896
R829 B.n391 B.n127 61.5896
R830 B.n397 B.n119 61.5896
R831 B.n403 B.n119 61.5896
R832 B.n403 B.n115 61.5896
R833 B.n409 B.n115 61.5896
R834 B.n415 B.n111 61.5896
R835 B.n415 B.n107 61.5896
R836 B.n422 B.n107 61.5896
R837 B.n428 B.n103 61.5896
R838 B.n428 B.n4 61.5896
R839 B.n674 B.n4 61.5896
R840 B.n674 B.n673 61.5896
R841 B.n673 B.n672 61.5896
R842 B.n672 B.n8 61.5896
R843 B.n437 B.n8 61.5896
R844 B.n665 B.n664 61.5896
R845 B.n664 B.n663 61.5896
R846 B.n663 B.n15 61.5896
R847 B.n657 B.n656 61.5896
R848 B.n656 B.n655 61.5896
R849 B.n655 B.n22 61.5896
R850 B.n649 B.n22 61.5896
R851 B.n648 B.n647 61.5896
R852 B.n647 B.n29 61.5896
R853 B.n641 B.n29 61.5896
R854 B.n640 B.n639 61.5896
R855 B.n639 B.n36 61.5896
R856 B.n633 B.n36 61.5896
R857 B.n632 B.n631 61.5896
R858 B.n631 B.n43 61.5896
R859 B.n625 B.n43 61.5896
R860 B.n625 B.n624 61.5896
R861 B.n624 B.n623 61.5896
R862 B.n623 B.n50 61.5896
R863 B.n617 B.n50 61.5896
R864 B.n616 B.n615 61.5896
R865 B.n615 B.n57 61.5896
R866 B.n609 B.n57 61.5896
R867 B.n609 B.n608 61.5896
R868 B.n608 B.n607 61.5896
R869 B.n82 B.n81 59.5399
R870 B.n532 B.n88 59.5399
R871 B.n257 B.n190 59.5399
R872 B.n275 B.n184 59.5399
R873 B.n127 B.t7 57.9667
R874 B.t3 B.n648 57.9667
R875 B.n373 B.t8 50.721
R876 B.n633 B.t4 50.721
R877 B.n422 B.t1 43.4752
R878 B.n665 B.t9 43.4752
R879 B.t0 B.n111 41.6637
R880 B.t5 B.n15 41.6637
R881 B.n159 B.t18 36.2294
R882 B.t11 B.n616 36.2294
R883 B.n135 B.t2 34.418
R884 B.t6 B.n640 34.418
R885 B.n329 B.n328 29.5029
R886 B.n333 B.n165 29.5029
R887 B.n478 B.n477 29.5029
R888 B.n605 B.n604 29.5029
R889 B.n81 B.n80 28.8975
R890 B.n88 B.n87 28.8975
R891 B.n190 B.n189 28.8975
R892 B.n184 B.n183 28.8975
R893 B.n385 B.t2 27.1722
R894 B.n641 B.t6 27.1722
R895 B.n349 B.t18 25.3607
R896 B.n617 B.t11 25.3607
R897 B.n409 B.t0 19.9264
R898 B.n657 B.t5 19.9264
R899 B.t1 B.n103 18.115
R900 B.n437 B.t9 18.115
R901 B B.n677 18.0485
R902 B.n143 B.t8 10.8692
R903 B.t4 B.n632 10.8692
R904 B.n329 B.n161 10.6151
R905 B.n339 B.n161 10.6151
R906 B.n340 B.n339 10.6151
R907 B.n341 B.n340 10.6151
R908 B.n341 B.n153 10.6151
R909 B.n351 B.n153 10.6151
R910 B.n352 B.n351 10.6151
R911 B.n353 B.n352 10.6151
R912 B.n353 B.n145 10.6151
R913 B.n363 B.n145 10.6151
R914 B.n364 B.n363 10.6151
R915 B.n365 B.n364 10.6151
R916 B.n365 B.n137 10.6151
R917 B.n375 B.n137 10.6151
R918 B.n376 B.n375 10.6151
R919 B.n377 B.n376 10.6151
R920 B.n377 B.n129 10.6151
R921 B.n387 B.n129 10.6151
R922 B.n388 B.n387 10.6151
R923 B.n389 B.n388 10.6151
R924 B.n389 B.n121 10.6151
R925 B.n399 B.n121 10.6151
R926 B.n400 B.n399 10.6151
R927 B.n401 B.n400 10.6151
R928 B.n401 B.n113 10.6151
R929 B.n411 B.n113 10.6151
R930 B.n412 B.n411 10.6151
R931 B.n413 B.n412 10.6151
R932 B.n413 B.n105 10.6151
R933 B.n424 B.n105 10.6151
R934 B.n425 B.n424 10.6151
R935 B.n426 B.n425 10.6151
R936 B.n426 B.n0 10.6151
R937 B.n328 B.n327 10.6151
R938 B.n327 B.n169 10.6151
R939 B.n322 B.n169 10.6151
R940 B.n322 B.n321 10.6151
R941 B.n321 B.n171 10.6151
R942 B.n316 B.n171 10.6151
R943 B.n316 B.n315 10.6151
R944 B.n315 B.n314 10.6151
R945 B.n314 B.n173 10.6151
R946 B.n308 B.n173 10.6151
R947 B.n308 B.n307 10.6151
R948 B.n307 B.n306 10.6151
R949 B.n306 B.n175 10.6151
R950 B.n300 B.n175 10.6151
R951 B.n300 B.n299 10.6151
R952 B.n299 B.n298 10.6151
R953 B.n298 B.n177 10.6151
R954 B.n292 B.n177 10.6151
R955 B.n292 B.n291 10.6151
R956 B.n291 B.n290 10.6151
R957 B.n290 B.n179 10.6151
R958 B.n284 B.n179 10.6151
R959 B.n284 B.n283 10.6151
R960 B.n283 B.n282 10.6151
R961 B.n282 B.n181 10.6151
R962 B.n276 B.n181 10.6151
R963 B.n274 B.n273 10.6151
R964 B.n273 B.n185 10.6151
R965 B.n267 B.n185 10.6151
R966 B.n267 B.n266 10.6151
R967 B.n266 B.n265 10.6151
R968 B.n265 B.n187 10.6151
R969 B.n259 B.n187 10.6151
R970 B.n259 B.n258 10.6151
R971 B.n256 B.n191 10.6151
R972 B.n250 B.n191 10.6151
R973 B.n250 B.n249 10.6151
R974 B.n249 B.n248 10.6151
R975 B.n248 B.n193 10.6151
R976 B.n242 B.n193 10.6151
R977 B.n242 B.n241 10.6151
R978 B.n241 B.n240 10.6151
R979 B.n240 B.n195 10.6151
R980 B.n234 B.n195 10.6151
R981 B.n234 B.n233 10.6151
R982 B.n233 B.n232 10.6151
R983 B.n232 B.n197 10.6151
R984 B.n226 B.n197 10.6151
R985 B.n226 B.n225 10.6151
R986 B.n225 B.n224 10.6151
R987 B.n224 B.n199 10.6151
R988 B.n218 B.n199 10.6151
R989 B.n218 B.n217 10.6151
R990 B.n217 B.n216 10.6151
R991 B.n216 B.n201 10.6151
R992 B.n210 B.n201 10.6151
R993 B.n210 B.n209 10.6151
R994 B.n209 B.n208 10.6151
R995 B.n208 B.n203 10.6151
R996 B.n203 B.n165 10.6151
R997 B.n334 B.n333 10.6151
R998 B.n335 B.n334 10.6151
R999 B.n335 B.n156 10.6151
R1000 B.n345 B.n156 10.6151
R1001 B.n346 B.n345 10.6151
R1002 B.n347 B.n346 10.6151
R1003 B.n347 B.n149 10.6151
R1004 B.n357 B.n149 10.6151
R1005 B.n358 B.n357 10.6151
R1006 B.n359 B.n358 10.6151
R1007 B.n359 B.n140 10.6151
R1008 B.n369 B.n140 10.6151
R1009 B.n370 B.n369 10.6151
R1010 B.n371 B.n370 10.6151
R1011 B.n371 B.n132 10.6151
R1012 B.n381 B.n132 10.6151
R1013 B.n382 B.n381 10.6151
R1014 B.n383 B.n382 10.6151
R1015 B.n383 B.n124 10.6151
R1016 B.n393 B.n124 10.6151
R1017 B.n394 B.n393 10.6151
R1018 B.n395 B.n394 10.6151
R1019 B.n395 B.n117 10.6151
R1020 B.n405 B.n117 10.6151
R1021 B.n406 B.n405 10.6151
R1022 B.n407 B.n406 10.6151
R1023 B.n407 B.n109 10.6151
R1024 B.n417 B.n109 10.6151
R1025 B.n418 B.n417 10.6151
R1026 B.n420 B.n418 10.6151
R1027 B.n420 B.n419 10.6151
R1028 B.n419 B.n101 10.6151
R1029 B.n431 B.n101 10.6151
R1030 B.n432 B.n431 10.6151
R1031 B.n433 B.n432 10.6151
R1032 B.n434 B.n433 10.6151
R1033 B.n435 B.n434 10.6151
R1034 B.n439 B.n435 10.6151
R1035 B.n440 B.n439 10.6151
R1036 B.n441 B.n440 10.6151
R1037 B.n442 B.n441 10.6151
R1038 B.n444 B.n442 10.6151
R1039 B.n445 B.n444 10.6151
R1040 B.n446 B.n445 10.6151
R1041 B.n447 B.n446 10.6151
R1042 B.n449 B.n447 10.6151
R1043 B.n450 B.n449 10.6151
R1044 B.n451 B.n450 10.6151
R1045 B.n452 B.n451 10.6151
R1046 B.n454 B.n452 10.6151
R1047 B.n455 B.n454 10.6151
R1048 B.n456 B.n455 10.6151
R1049 B.n457 B.n456 10.6151
R1050 B.n459 B.n457 10.6151
R1051 B.n460 B.n459 10.6151
R1052 B.n461 B.n460 10.6151
R1053 B.n462 B.n461 10.6151
R1054 B.n464 B.n462 10.6151
R1055 B.n465 B.n464 10.6151
R1056 B.n466 B.n465 10.6151
R1057 B.n467 B.n466 10.6151
R1058 B.n469 B.n467 10.6151
R1059 B.n470 B.n469 10.6151
R1060 B.n471 B.n470 10.6151
R1061 B.n472 B.n471 10.6151
R1062 B.n474 B.n472 10.6151
R1063 B.n475 B.n474 10.6151
R1064 B.n476 B.n475 10.6151
R1065 B.n477 B.n476 10.6151
R1066 B.n669 B.n1 10.6151
R1067 B.n669 B.n668 10.6151
R1068 B.n668 B.n667 10.6151
R1069 B.n667 B.n10 10.6151
R1070 B.n661 B.n10 10.6151
R1071 B.n661 B.n660 10.6151
R1072 B.n660 B.n659 10.6151
R1073 B.n659 B.n17 10.6151
R1074 B.n653 B.n17 10.6151
R1075 B.n653 B.n652 10.6151
R1076 B.n652 B.n651 10.6151
R1077 B.n651 B.n24 10.6151
R1078 B.n645 B.n24 10.6151
R1079 B.n645 B.n644 10.6151
R1080 B.n644 B.n643 10.6151
R1081 B.n643 B.n31 10.6151
R1082 B.n637 B.n31 10.6151
R1083 B.n637 B.n636 10.6151
R1084 B.n636 B.n635 10.6151
R1085 B.n635 B.n38 10.6151
R1086 B.n629 B.n38 10.6151
R1087 B.n629 B.n628 10.6151
R1088 B.n628 B.n627 10.6151
R1089 B.n627 B.n45 10.6151
R1090 B.n621 B.n45 10.6151
R1091 B.n621 B.n620 10.6151
R1092 B.n620 B.n619 10.6151
R1093 B.n619 B.n52 10.6151
R1094 B.n613 B.n52 10.6151
R1095 B.n613 B.n612 10.6151
R1096 B.n612 B.n611 10.6151
R1097 B.n611 B.n59 10.6151
R1098 B.n605 B.n59 10.6151
R1099 B.n604 B.n603 10.6151
R1100 B.n603 B.n66 10.6151
R1101 B.n597 B.n66 10.6151
R1102 B.n597 B.n596 10.6151
R1103 B.n596 B.n595 10.6151
R1104 B.n595 B.n68 10.6151
R1105 B.n589 B.n68 10.6151
R1106 B.n589 B.n588 10.6151
R1107 B.n588 B.n587 10.6151
R1108 B.n587 B.n70 10.6151
R1109 B.n581 B.n70 10.6151
R1110 B.n581 B.n580 10.6151
R1111 B.n580 B.n579 10.6151
R1112 B.n579 B.n72 10.6151
R1113 B.n573 B.n72 10.6151
R1114 B.n573 B.n572 10.6151
R1115 B.n572 B.n571 10.6151
R1116 B.n571 B.n74 10.6151
R1117 B.n565 B.n74 10.6151
R1118 B.n565 B.n564 10.6151
R1119 B.n564 B.n563 10.6151
R1120 B.n563 B.n76 10.6151
R1121 B.n557 B.n76 10.6151
R1122 B.n557 B.n556 10.6151
R1123 B.n556 B.n555 10.6151
R1124 B.n555 B.n78 10.6151
R1125 B.n549 B.n548 10.6151
R1126 B.n548 B.n547 10.6151
R1127 B.n547 B.n83 10.6151
R1128 B.n541 B.n83 10.6151
R1129 B.n541 B.n540 10.6151
R1130 B.n540 B.n539 10.6151
R1131 B.n539 B.n85 10.6151
R1132 B.n533 B.n85 10.6151
R1133 B.n531 B.n530 10.6151
R1134 B.n530 B.n89 10.6151
R1135 B.n524 B.n89 10.6151
R1136 B.n524 B.n523 10.6151
R1137 B.n523 B.n522 10.6151
R1138 B.n522 B.n91 10.6151
R1139 B.n516 B.n91 10.6151
R1140 B.n516 B.n515 10.6151
R1141 B.n515 B.n514 10.6151
R1142 B.n514 B.n93 10.6151
R1143 B.n508 B.n93 10.6151
R1144 B.n508 B.n507 10.6151
R1145 B.n507 B.n506 10.6151
R1146 B.n506 B.n95 10.6151
R1147 B.n500 B.n95 10.6151
R1148 B.n500 B.n499 10.6151
R1149 B.n499 B.n498 10.6151
R1150 B.n498 B.n97 10.6151
R1151 B.n492 B.n97 10.6151
R1152 B.n492 B.n491 10.6151
R1153 B.n491 B.n490 10.6151
R1154 B.n490 B.n99 10.6151
R1155 B.n484 B.n99 10.6151
R1156 B.n484 B.n483 10.6151
R1157 B.n483 B.n482 10.6151
R1158 B.n482 B.n478 10.6151
R1159 B.n677 B.n0 8.11757
R1160 B.n677 B.n1 8.11757
R1161 B.n275 B.n274 6.5566
R1162 B.n258 B.n257 6.5566
R1163 B.n549 B.n82 6.5566
R1164 B.n533 B.n532 6.5566
R1165 B.n276 B.n275 4.05904
R1166 B.n257 B.n256 4.05904
R1167 B.n82 B.n78 4.05904
R1168 B.n532 B.n531 4.05904
R1169 B.n397 B.t7 3.62339
R1170 B.n649 B.t3 3.62339
R1171 VP.n32 VP.n7 174.512
R1172 VP.n54 VP.n53 174.512
R1173 VP.n31 VP.n30 174.512
R1174 VP.n14 VP.t5 172.143
R1175 VP.n16 VP.n15 161.3
R1176 VP.n17 VP.n12 161.3
R1177 VP.n19 VP.n18 161.3
R1178 VP.n21 VP.n20 161.3
R1179 VP.n22 VP.n10 161.3
R1180 VP.n25 VP.n24 161.3
R1181 VP.n26 VP.n9 161.3
R1182 VP.n28 VP.n27 161.3
R1183 VP.n29 VP.n8 161.3
R1184 VP.n52 VP.n0 161.3
R1185 VP.n51 VP.n50 161.3
R1186 VP.n49 VP.n1 161.3
R1187 VP.n48 VP.n47 161.3
R1188 VP.n45 VP.n2 161.3
R1189 VP.n44 VP.n43 161.3
R1190 VP.n42 VP.n41 161.3
R1191 VP.n40 VP.n4 161.3
R1192 VP.n39 VP.n38 161.3
R1193 VP.n37 VP.n36 161.3
R1194 VP.n35 VP.n6 161.3
R1195 VP.n34 VP.n33 161.3
R1196 VP.n7 VP.t9 142.731
R1197 VP.n5 VP.t6 142.731
R1198 VP.n3 VP.t2 142.731
R1199 VP.n46 VP.t8 142.731
R1200 VP.n53 VP.t4 142.731
R1201 VP.n30 VP.t3 142.731
R1202 VP.n23 VP.t7 142.731
R1203 VP.n11 VP.t0 142.731
R1204 VP.n13 VP.t1 142.731
R1205 VP.n14 VP.n13 52.0614
R1206 VP.n36 VP.n35 41.9503
R1207 VP.n51 VP.n1 41.9503
R1208 VP.n28 VP.n9 41.9503
R1209 VP.n32 VP.n31 41.2619
R1210 VP.n41 VP.n40 40.979
R1211 VP.n45 VP.n44 40.979
R1212 VP.n22 VP.n21 40.979
R1213 VP.n18 VP.n17 40.979
R1214 VP.n40 VP.n39 40.0078
R1215 VP.n47 VP.n45 40.0078
R1216 VP.n24 VP.n22 40.0078
R1217 VP.n17 VP.n16 40.0078
R1218 VP.n35 VP.n34 39.0365
R1219 VP.n52 VP.n51 39.0365
R1220 VP.n29 VP.n28 39.0365
R1221 VP.n15 VP.n14 27.217
R1222 VP.n36 VP.n5 12.7233
R1223 VP.n46 VP.n1 12.7233
R1224 VP.n23 VP.n9 12.7233
R1225 VP.n41 VP.n3 12.234
R1226 VP.n44 VP.n3 12.234
R1227 VP.n18 VP.n11 12.234
R1228 VP.n21 VP.n11 12.234
R1229 VP.n39 VP.n5 11.7447
R1230 VP.n47 VP.n46 11.7447
R1231 VP.n24 VP.n23 11.7447
R1232 VP.n16 VP.n13 11.7447
R1233 VP.n34 VP.n7 11.2553
R1234 VP.n53 VP.n52 11.2553
R1235 VP.n30 VP.n29 11.2553
R1236 VP.n15 VP.n12 0.189894
R1237 VP.n19 VP.n12 0.189894
R1238 VP.n20 VP.n19 0.189894
R1239 VP.n20 VP.n10 0.189894
R1240 VP.n25 VP.n10 0.189894
R1241 VP.n26 VP.n25 0.189894
R1242 VP.n27 VP.n26 0.189894
R1243 VP.n27 VP.n8 0.189894
R1244 VP.n31 VP.n8 0.189894
R1245 VP.n33 VP.n32 0.189894
R1246 VP.n33 VP.n6 0.189894
R1247 VP.n37 VP.n6 0.189894
R1248 VP.n38 VP.n37 0.189894
R1249 VP.n38 VP.n4 0.189894
R1250 VP.n42 VP.n4 0.189894
R1251 VP.n43 VP.n42 0.189894
R1252 VP.n43 VP.n2 0.189894
R1253 VP.n48 VP.n2 0.189894
R1254 VP.n49 VP.n48 0.189894
R1255 VP.n50 VP.n49 0.189894
R1256 VP.n50 VP.n0 0.189894
R1257 VP.n54 VP.n0 0.189894
R1258 VP VP.n54 0.0516364
R1259 VTAIL.n11 VTAIL.t7 54.1323
R1260 VTAIL.n17 VTAIL.t1 54.1322
R1261 VTAIL.n2 VTAIL.t18 54.1322
R1262 VTAIL.n16 VTAIL.t16 54.1322
R1263 VTAIL.n15 VTAIL.n14 51.2502
R1264 VTAIL.n13 VTAIL.n12 51.2502
R1265 VTAIL.n10 VTAIL.n9 51.2502
R1266 VTAIL.n8 VTAIL.n7 51.2502
R1267 VTAIL.n19 VTAIL.n18 51.2491
R1268 VTAIL.n1 VTAIL.n0 51.2491
R1269 VTAIL.n4 VTAIL.n3 51.2491
R1270 VTAIL.n6 VTAIL.n5 51.2491
R1271 VTAIL.n8 VTAIL.n6 20.8583
R1272 VTAIL.n17 VTAIL.n16 19.5738
R1273 VTAIL.n18 VTAIL.t4 2.8826
R1274 VTAIL.n18 VTAIL.t3 2.8826
R1275 VTAIL.n0 VTAIL.t8 2.8826
R1276 VTAIL.n0 VTAIL.t2 2.8826
R1277 VTAIL.n3 VTAIL.t19 2.8826
R1278 VTAIL.n3 VTAIL.t13 2.8826
R1279 VTAIL.n5 VTAIL.t15 2.8826
R1280 VTAIL.n5 VTAIL.t11 2.8826
R1281 VTAIL.n14 VTAIL.t10 2.8826
R1282 VTAIL.n14 VTAIL.t14 2.8826
R1283 VTAIL.n12 VTAIL.t17 2.8826
R1284 VTAIL.n12 VTAIL.t12 2.8826
R1285 VTAIL.n9 VTAIL.t9 2.8826
R1286 VTAIL.n9 VTAIL.t0 2.8826
R1287 VTAIL.n7 VTAIL.t6 2.8826
R1288 VTAIL.n7 VTAIL.t5 2.8826
R1289 VTAIL.n10 VTAIL.n8 1.28498
R1290 VTAIL.n11 VTAIL.n10 1.28498
R1291 VTAIL.n15 VTAIL.n13 1.28498
R1292 VTAIL.n16 VTAIL.n15 1.28498
R1293 VTAIL.n6 VTAIL.n4 1.28498
R1294 VTAIL.n4 VTAIL.n2 1.28498
R1295 VTAIL.n19 VTAIL.n17 1.28498
R1296 VTAIL.n13 VTAIL.n11 1.11257
R1297 VTAIL.n2 VTAIL.n1 1.11257
R1298 VTAIL VTAIL.n1 1.02205
R1299 VTAIL VTAIL.n19 0.263431
R1300 VDD1.n1 VDD1.t4 72.0956
R1301 VDD1.n3 VDD1.t0 72.0955
R1302 VDD1.n5 VDD1.n4 68.8359
R1303 VDD1.n1 VDD1.n0 67.929
R1304 VDD1.n7 VDD1.n6 67.9289
R1305 VDD1.n3 VDD1.n2 67.9279
R1306 VDD1.n7 VDD1.n5 36.9643
R1307 VDD1.n6 VDD1.t2 2.8826
R1308 VDD1.n6 VDD1.t6 2.8826
R1309 VDD1.n0 VDD1.t8 2.8826
R1310 VDD1.n0 VDD1.t9 2.8826
R1311 VDD1.n4 VDD1.t1 2.8826
R1312 VDD1.n4 VDD1.t5 2.8826
R1313 VDD1.n2 VDD1.t3 2.8826
R1314 VDD1.n2 VDD1.t7 2.8826
R1315 VDD1 VDD1.n7 0.905672
R1316 VDD1 VDD1.n1 0.37981
R1317 VDD1.n5 VDD1.n3 0.266275
R1318 VN.n23 VN.n22 174.512
R1319 VN.n47 VN.n46 174.512
R1320 VN.n6 VN.t2 172.143
R1321 VN.n31 VN.t6 172.143
R1322 VN.n45 VN.n24 161.3
R1323 VN.n44 VN.n43 161.3
R1324 VN.n42 VN.n25 161.3
R1325 VN.n41 VN.n40 161.3
R1326 VN.n39 VN.n26 161.3
R1327 VN.n38 VN.n37 161.3
R1328 VN.n36 VN.n35 161.3
R1329 VN.n34 VN.n29 161.3
R1330 VN.n33 VN.n32 161.3
R1331 VN.n21 VN.n0 161.3
R1332 VN.n20 VN.n19 161.3
R1333 VN.n18 VN.n1 161.3
R1334 VN.n17 VN.n16 161.3
R1335 VN.n14 VN.n2 161.3
R1336 VN.n13 VN.n12 161.3
R1337 VN.n11 VN.n10 161.3
R1338 VN.n9 VN.n4 161.3
R1339 VN.n8 VN.n7 161.3
R1340 VN.n5 VN.t5 142.731
R1341 VN.n3 VN.t1 142.731
R1342 VN.n15 VN.t4 142.731
R1343 VN.n22 VN.t8 142.731
R1344 VN.n30 VN.t3 142.731
R1345 VN.n28 VN.t0 142.731
R1346 VN.n27 VN.t9 142.731
R1347 VN.n46 VN.t7 142.731
R1348 VN.n6 VN.n5 52.0614
R1349 VN.n31 VN.n30 52.0614
R1350 VN.n20 VN.n1 41.9503
R1351 VN.n44 VN.n25 41.9503
R1352 VN VN.n47 41.6425
R1353 VN.n10 VN.n9 40.979
R1354 VN.n14 VN.n13 40.979
R1355 VN.n35 VN.n34 40.979
R1356 VN.n39 VN.n38 40.979
R1357 VN.n9 VN.n8 40.0078
R1358 VN.n16 VN.n14 40.0078
R1359 VN.n34 VN.n33 40.0078
R1360 VN.n40 VN.n39 40.0078
R1361 VN.n21 VN.n20 39.0365
R1362 VN.n45 VN.n44 39.0365
R1363 VN.n32 VN.n31 27.217
R1364 VN.n7 VN.n6 27.217
R1365 VN.n15 VN.n1 12.7233
R1366 VN.n27 VN.n25 12.7233
R1367 VN.n10 VN.n3 12.234
R1368 VN.n13 VN.n3 12.234
R1369 VN.n38 VN.n28 12.234
R1370 VN.n35 VN.n28 12.234
R1371 VN.n8 VN.n5 11.7447
R1372 VN.n16 VN.n15 11.7447
R1373 VN.n33 VN.n30 11.7447
R1374 VN.n40 VN.n27 11.7447
R1375 VN.n22 VN.n21 11.2553
R1376 VN.n46 VN.n45 11.2553
R1377 VN.n47 VN.n24 0.189894
R1378 VN.n43 VN.n24 0.189894
R1379 VN.n43 VN.n42 0.189894
R1380 VN.n42 VN.n41 0.189894
R1381 VN.n41 VN.n26 0.189894
R1382 VN.n37 VN.n26 0.189894
R1383 VN.n37 VN.n36 0.189894
R1384 VN.n36 VN.n29 0.189894
R1385 VN.n32 VN.n29 0.189894
R1386 VN.n7 VN.n4 0.189894
R1387 VN.n11 VN.n4 0.189894
R1388 VN.n12 VN.n11 0.189894
R1389 VN.n12 VN.n2 0.189894
R1390 VN.n17 VN.n2 0.189894
R1391 VN.n18 VN.n17 0.189894
R1392 VN.n19 VN.n18 0.189894
R1393 VN.n19 VN.n0 0.189894
R1394 VN.n23 VN.n0 0.189894
R1395 VN VN.n23 0.0516364
R1396 VDD2.n1 VDD2.t7 72.0955
R1397 VDD2.n4 VDD2.t2 70.8111
R1398 VDD2.n3 VDD2.n2 68.8359
R1399 VDD2 VDD2.n7 68.8341
R1400 VDD2.n6 VDD2.n5 67.929
R1401 VDD2.n1 VDD2.n0 67.9279
R1402 VDD2.n4 VDD2.n3 35.739
R1403 VDD2.n7 VDD2.t6 2.8826
R1404 VDD2.n7 VDD2.t3 2.8826
R1405 VDD2.n5 VDD2.t0 2.8826
R1406 VDD2.n5 VDD2.t9 2.8826
R1407 VDD2.n2 VDD2.t5 2.8826
R1408 VDD2.n2 VDD2.t1 2.8826
R1409 VDD2.n0 VDD2.t4 2.8826
R1410 VDD2.n0 VDD2.t8 2.8826
R1411 VDD2.n6 VDD2.n4 1.28498
R1412 VDD2 VDD2.n6 0.37981
R1413 VDD2.n3 VDD2.n1 0.266275
C0 VN VTAIL 5.38324f
C1 VDD2 VTAIL 8.05795f
C2 VP VN 5.32978f
C3 VP VDD2 0.398997f
C4 VN VDD1 0.149637f
C5 VDD2 VDD1 1.2503f
C6 VP VTAIL 5.39756f
C7 VDD2 VN 5.03992f
C8 VDD1 VTAIL 8.01694f
C9 VP VDD1 5.28647f
C10 VDD2 B 4.589587f
C11 VDD1 B 4.551146f
C12 VTAIL B 4.814776f
C13 VN B 10.84809f
C14 VP B 9.265246f
C15 VDD2.t7 B 1.36991f
C16 VDD2.t4 B 0.12565f
C17 VDD2.t8 B 0.12565f
C18 VDD2.n0 B 1.07374f
C19 VDD2.n1 B 0.630712f
C20 VDD2.t5 B 0.12565f
C21 VDD2.t1 B 0.12565f
C22 VDD2.n2 B 1.07842f
C23 VDD2.n3 B 1.69414f
C24 VDD2.t2 B 1.36389f
C25 VDD2.n4 B 1.98255f
C26 VDD2.t0 B 0.12565f
C27 VDD2.t9 B 0.12565f
C28 VDD2.n5 B 1.07375f
C29 VDD2.n6 B 0.304802f
C30 VDD2.t6 B 0.12565f
C31 VDD2.t3 B 0.12565f
C32 VDD2.n7 B 1.07839f
C33 VN.n0 B 0.035512f
C34 VN.t8 B 0.754613f
C35 VN.n1 B 0.054313f
C36 VN.n2 B 0.035512f
C37 VN.t1 B 0.754613f
C38 VN.n3 B 0.29704f
C39 VN.n4 B 0.035512f
C40 VN.t5 B 0.754613f
C41 VN.n5 B 0.347962f
C42 VN.t2 B 0.822677f
C43 VN.n6 B 0.370855f
C44 VN.n7 B 0.182923f
C45 VN.n8 B 0.053763f
C46 VN.n9 B 0.028721f
C47 VN.n10 B 0.05406f
C48 VN.n11 B 0.035512f
C49 VN.n12 B 0.035512f
C50 VN.n13 B 0.05406f
C51 VN.n14 B 0.028721f
C52 VN.t4 B 0.754613f
C53 VN.n15 B 0.29704f
C54 VN.n16 B 0.053763f
C55 VN.n17 B 0.035512f
C56 VN.n18 B 0.035512f
C57 VN.n19 B 0.035512f
C58 VN.n20 B 0.028812f
C59 VN.n21 B 0.053418f
C60 VN.n22 B 0.35157f
C61 VN.n23 B 0.031987f
C62 VN.n24 B 0.035512f
C63 VN.t7 B 0.754613f
C64 VN.n25 B 0.054313f
C65 VN.n26 B 0.035512f
C66 VN.t9 B 0.754613f
C67 VN.n27 B 0.29704f
C68 VN.t0 B 0.754613f
C69 VN.n28 B 0.29704f
C70 VN.n29 B 0.035512f
C71 VN.t3 B 0.754613f
C72 VN.n30 B 0.347962f
C73 VN.t6 B 0.822677f
C74 VN.n31 B 0.370855f
C75 VN.n32 B 0.182923f
C76 VN.n33 B 0.053763f
C77 VN.n34 B 0.028721f
C78 VN.n35 B 0.05406f
C79 VN.n36 B 0.035512f
C80 VN.n37 B 0.035512f
C81 VN.n38 B 0.05406f
C82 VN.n39 B 0.028721f
C83 VN.n40 B 0.053763f
C84 VN.n41 B 0.035512f
C85 VN.n42 B 0.035512f
C86 VN.n43 B 0.035512f
C87 VN.n44 B 0.028812f
C88 VN.n45 B 0.053418f
C89 VN.n46 B 0.35157f
C90 VN.n47 B 1.45067f
C91 VDD1.t4 B 1.38182f
C92 VDD1.t8 B 0.126741f
C93 VDD1.t9 B 0.126741f
C94 VDD1.n0 B 1.08307f
C95 VDD1.n1 B 0.64268f
C96 VDD1.t0 B 1.38181f
C97 VDD1.t3 B 0.126741f
C98 VDD1.t7 B 0.126741f
C99 VDD1.n2 B 1.08307f
C100 VDD1.n3 B 0.636189f
C101 VDD1.t1 B 0.126741f
C102 VDD1.t5 B 0.126741f
C103 VDD1.n4 B 1.08778f
C104 VDD1.n5 B 1.78854f
C105 VDD1.t2 B 0.126741f
C106 VDD1.t6 B 0.126741f
C107 VDD1.n6 B 1.08306f
C108 VDD1.n7 B 2.02142f
C109 VTAIL.t8 B 0.143702f
C110 VTAIL.t2 B 0.143702f
C111 VTAIL.n0 B 1.16238f
C112 VTAIL.n1 B 0.418321f
C113 VTAIL.t18 B 1.47919f
C114 VTAIL.n2 B 0.515855f
C115 VTAIL.t19 B 0.143702f
C116 VTAIL.t13 B 0.143702f
C117 VTAIL.n3 B 1.16238f
C118 VTAIL.n4 B 0.455452f
C119 VTAIL.t15 B 0.143702f
C120 VTAIL.t11 B 0.143702f
C121 VTAIL.n5 B 1.16238f
C122 VTAIL.n6 B 1.42971f
C123 VTAIL.t6 B 0.143702f
C124 VTAIL.t5 B 0.143702f
C125 VTAIL.n7 B 1.16239f
C126 VTAIL.n8 B 1.4297f
C127 VTAIL.t9 B 0.143702f
C128 VTAIL.t0 B 0.143702f
C129 VTAIL.n9 B 1.16239f
C130 VTAIL.n10 B 0.455444f
C131 VTAIL.t7 B 1.4792f
C132 VTAIL.n11 B 0.515842f
C133 VTAIL.t17 B 0.143702f
C134 VTAIL.t12 B 0.143702f
C135 VTAIL.n12 B 1.16239f
C136 VTAIL.n13 B 0.440738f
C137 VTAIL.t10 B 0.143702f
C138 VTAIL.t14 B 0.143702f
C139 VTAIL.n14 B 1.16239f
C140 VTAIL.n15 B 0.455444f
C141 VTAIL.t16 B 1.47919f
C142 VTAIL.n16 B 1.39526f
C143 VTAIL.t1 B 1.47919f
C144 VTAIL.n17 B 1.39526f
C145 VTAIL.t4 B 0.143702f
C146 VTAIL.t3 B 0.143702f
C147 VTAIL.n18 B 1.16238f
C148 VTAIL.n19 B 0.368322f
C149 VP.n0 B 0.036305f
C150 VP.t4 B 0.771485f
C151 VP.n1 B 0.055528f
C152 VP.n2 B 0.036305f
C153 VP.t2 B 0.771485f
C154 VP.n3 B 0.303682f
C155 VP.n4 B 0.036305f
C156 VP.t6 B 0.771485f
C157 VP.n5 B 0.303682f
C158 VP.n6 B 0.036305f
C159 VP.t9 B 0.771485f
C160 VP.n7 B 0.35943f
C161 VP.n8 B 0.036305f
C162 VP.t3 B 0.771485f
C163 VP.n9 B 0.055528f
C164 VP.n10 B 0.036305f
C165 VP.t0 B 0.771485f
C166 VP.n11 B 0.303682f
C167 VP.n12 B 0.036305f
C168 VP.t1 B 0.771485f
C169 VP.n13 B 0.355742f
C170 VP.t5 B 0.841072f
C171 VP.n14 B 0.379147f
C172 VP.n15 B 0.187013f
C173 VP.n16 B 0.054965f
C174 VP.n17 B 0.029363f
C175 VP.n18 B 0.055269f
C176 VP.n19 B 0.036305f
C177 VP.n20 B 0.036305f
C178 VP.n21 B 0.055269f
C179 VP.n22 B 0.029363f
C180 VP.t7 B 0.771485f
C181 VP.n23 B 0.303682f
C182 VP.n24 B 0.054965f
C183 VP.n25 B 0.036305f
C184 VP.n26 B 0.036305f
C185 VP.n27 B 0.036305f
C186 VP.n28 B 0.029456f
C187 VP.n29 B 0.054612f
C188 VP.n30 B 0.35943f
C189 VP.n31 B 1.45925f
C190 VP.n32 B 1.49088f
C191 VP.n33 B 0.036305f
C192 VP.n34 B 0.054612f
C193 VP.n35 B 0.029456f
C194 VP.n36 B 0.055528f
C195 VP.n37 B 0.036305f
C196 VP.n38 B 0.036305f
C197 VP.n39 B 0.054965f
C198 VP.n40 B 0.029363f
C199 VP.n41 B 0.055269f
C200 VP.n42 B 0.036305f
C201 VP.n43 B 0.036305f
C202 VP.n44 B 0.055269f
C203 VP.n45 B 0.029363f
C204 VP.t8 B 0.771485f
C205 VP.n46 B 0.303682f
C206 VP.n47 B 0.054965f
C207 VP.n48 B 0.036305f
C208 VP.n49 B 0.036305f
C209 VP.n50 B 0.036305f
C210 VP.n51 B 0.029456f
C211 VP.n52 B 0.054612f
C212 VP.n53 B 0.35943f
C213 VP.n54 B 0.032702f
.ends

