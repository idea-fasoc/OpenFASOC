* NGSPICE file created from diff_pair_sample_1146.ext - technology: sky130A

.subckt diff_pair_sample_1146 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t19 VP.t0 VDD1.t9 B.t9 sky130_fd_pr__nfet_01v8 ad=1.6533 pd=10.35 as=1.6533 ps=10.35 w=10.02 l=3.54
X1 VTAIL.t3 VN.t0 VDD2.t9 B.t3 sky130_fd_pr__nfet_01v8 ad=1.6533 pd=10.35 as=1.6533 ps=10.35 w=10.02 l=3.54
X2 B.t23 B.t21 B.t22 B.t15 sky130_fd_pr__nfet_01v8 ad=3.9078 pd=20.82 as=0 ps=0 w=10.02 l=3.54
X3 VTAIL.t18 VP.t1 VDD1.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=1.6533 pd=10.35 as=1.6533 ps=10.35 w=10.02 l=3.54
X4 VDD2.t8 VN.t1 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=3.9078 pd=20.82 as=1.6533 ps=10.35 w=10.02 l=3.54
X5 VDD1.t6 VP.t2 VTAIL.t17 B.t8 sky130_fd_pr__nfet_01v8 ad=1.6533 pd=10.35 as=3.9078 ps=20.82 w=10.02 l=3.54
X6 VTAIL.t4 VN.t2 VDD2.t7 B.t4 sky130_fd_pr__nfet_01v8 ad=1.6533 pd=10.35 as=1.6533 ps=10.35 w=10.02 l=3.54
X7 VTAIL.t16 VP.t3 VDD1.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=1.6533 pd=10.35 as=1.6533 ps=10.35 w=10.02 l=3.54
X8 VDD1.t0 VP.t4 VTAIL.t15 B.t1 sky130_fd_pr__nfet_01v8 ad=1.6533 pd=10.35 as=1.6533 ps=10.35 w=10.02 l=3.54
X9 VDD1.t3 VP.t5 VTAIL.t14 B.t5 sky130_fd_pr__nfet_01v8 ad=1.6533 pd=10.35 as=1.6533 ps=10.35 w=10.02 l=3.54
X10 VTAIL.t9 VN.t3 VDD2.t6 B.t9 sky130_fd_pr__nfet_01v8 ad=1.6533 pd=10.35 as=1.6533 ps=10.35 w=10.02 l=3.54
X11 B.t20 B.t18 B.t19 B.t11 sky130_fd_pr__nfet_01v8 ad=3.9078 pd=20.82 as=0 ps=0 w=10.02 l=3.54
X12 VDD1.t8 VP.t6 VTAIL.t13 B.t6 sky130_fd_pr__nfet_01v8 ad=1.6533 pd=10.35 as=3.9078 ps=20.82 w=10.02 l=3.54
X13 VDD2.t5 VN.t4 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.6533 pd=10.35 as=1.6533 ps=10.35 w=10.02 l=3.54
X14 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=3.9078 pd=20.82 as=0 ps=0 w=10.02 l=3.54
X15 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=3.9078 pd=20.82 as=0 ps=0 w=10.02 l=3.54
X16 VDD2.t4 VN.t5 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=1.6533 pd=10.35 as=3.9078 ps=20.82 w=10.02 l=3.54
X17 VDD2.t3 VN.t6 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=1.6533 pd=10.35 as=1.6533 ps=10.35 w=10.02 l=3.54
X18 VTAIL.t0 VN.t7 VDD2.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=1.6533 pd=10.35 as=1.6533 ps=10.35 w=10.02 l=3.54
X19 VDD1.t5 VP.t7 VTAIL.t12 B.t7 sky130_fd_pr__nfet_01v8 ad=3.9078 pd=20.82 as=1.6533 ps=10.35 w=10.02 l=3.54
X20 VDD2.t1 VN.t8 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=3.9078 pd=20.82 as=1.6533 ps=10.35 w=10.02 l=3.54
X21 VTAIL.t11 VP.t8 VDD1.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.6533 pd=10.35 as=1.6533 ps=10.35 w=10.02 l=3.54
X22 VDD1.t2 VP.t9 VTAIL.t10 B.t2 sky130_fd_pr__nfet_01v8 ad=3.9078 pd=20.82 as=1.6533 ps=10.35 w=10.02 l=3.54
X23 VDD2.t0 VN.t9 VTAIL.t8 B.t8 sky130_fd_pr__nfet_01v8 ad=1.6533 pd=10.35 as=3.9078 ps=20.82 w=10.02 l=3.54
R0 VP.n32 VP.n31 161.3
R1 VP.n33 VP.n28 161.3
R2 VP.n35 VP.n34 161.3
R3 VP.n36 VP.n27 161.3
R4 VP.n38 VP.n37 161.3
R5 VP.n39 VP.n26 161.3
R6 VP.n41 VP.n40 161.3
R7 VP.n42 VP.n25 161.3
R8 VP.n44 VP.n43 161.3
R9 VP.n45 VP.n24 161.3
R10 VP.n47 VP.n46 161.3
R11 VP.n48 VP.n23 161.3
R12 VP.n50 VP.n49 161.3
R13 VP.n51 VP.n22 161.3
R14 VP.n54 VP.n53 161.3
R15 VP.n55 VP.n21 161.3
R16 VP.n57 VP.n56 161.3
R17 VP.n58 VP.n20 161.3
R18 VP.n60 VP.n59 161.3
R19 VP.n61 VP.n19 161.3
R20 VP.n63 VP.n62 161.3
R21 VP.n64 VP.n18 161.3
R22 VP.n66 VP.n65 161.3
R23 VP.n117 VP.n116 161.3
R24 VP.n115 VP.n1 161.3
R25 VP.n114 VP.n113 161.3
R26 VP.n112 VP.n2 161.3
R27 VP.n111 VP.n110 161.3
R28 VP.n109 VP.n3 161.3
R29 VP.n108 VP.n107 161.3
R30 VP.n106 VP.n4 161.3
R31 VP.n105 VP.n104 161.3
R32 VP.n102 VP.n5 161.3
R33 VP.n101 VP.n100 161.3
R34 VP.n99 VP.n6 161.3
R35 VP.n98 VP.n97 161.3
R36 VP.n96 VP.n7 161.3
R37 VP.n95 VP.n94 161.3
R38 VP.n93 VP.n8 161.3
R39 VP.n92 VP.n91 161.3
R40 VP.n90 VP.n9 161.3
R41 VP.n89 VP.n88 161.3
R42 VP.n87 VP.n10 161.3
R43 VP.n86 VP.n85 161.3
R44 VP.n84 VP.n11 161.3
R45 VP.n83 VP.n82 161.3
R46 VP.n81 VP.n80 161.3
R47 VP.n79 VP.n13 161.3
R48 VP.n78 VP.n77 161.3
R49 VP.n76 VP.n14 161.3
R50 VP.n75 VP.n74 161.3
R51 VP.n73 VP.n15 161.3
R52 VP.n72 VP.n71 161.3
R53 VP.n70 VP.n16 161.3
R54 VP.n30 VP.t9 101.947
R55 VP.n69 VP.n68 78.4415
R56 VP.n118 VP.n0 78.4415
R57 VP.n67 VP.n17 78.4415
R58 VP.n8 VP.t4 68.2158
R59 VP.n68 VP.t7 68.2158
R60 VP.n12 VP.t0 68.2158
R61 VP.n103 VP.t3 68.2158
R62 VP.n0 VP.t6 68.2158
R63 VP.n25 VP.t5 68.2158
R64 VP.n17 VP.t2 68.2158
R65 VP.n52 VP.t1 68.2158
R66 VP.n29 VP.t8 68.2158
R67 VP.n69 VP.n67 56.8518
R68 VP.n30 VP.n29 56.6961
R69 VP.n74 VP.n14 56.5617
R70 VP.n110 VP.n2 56.5617
R71 VP.n59 VP.n19 56.5617
R72 VP.n89 VP.n10 46.874
R73 VP.n97 VP.n6 46.874
R74 VP.n46 VP.n23 46.874
R75 VP.n38 VP.n27 46.874
R76 VP.n85 VP.n10 34.28
R77 VP.n101 VP.n6 34.28
R78 VP.n50 VP.n23 34.28
R79 VP.n34 VP.n27 34.28
R80 VP.n72 VP.n16 24.5923
R81 VP.n73 VP.n72 24.5923
R82 VP.n74 VP.n73 24.5923
R83 VP.n78 VP.n14 24.5923
R84 VP.n79 VP.n78 24.5923
R85 VP.n80 VP.n79 24.5923
R86 VP.n84 VP.n83 24.5923
R87 VP.n85 VP.n84 24.5923
R88 VP.n90 VP.n89 24.5923
R89 VP.n91 VP.n90 24.5923
R90 VP.n91 VP.n8 24.5923
R91 VP.n95 VP.n8 24.5923
R92 VP.n96 VP.n95 24.5923
R93 VP.n97 VP.n96 24.5923
R94 VP.n102 VP.n101 24.5923
R95 VP.n104 VP.n102 24.5923
R96 VP.n108 VP.n4 24.5923
R97 VP.n109 VP.n108 24.5923
R98 VP.n110 VP.n109 24.5923
R99 VP.n114 VP.n2 24.5923
R100 VP.n115 VP.n114 24.5923
R101 VP.n116 VP.n115 24.5923
R102 VP.n63 VP.n19 24.5923
R103 VP.n64 VP.n63 24.5923
R104 VP.n65 VP.n64 24.5923
R105 VP.n51 VP.n50 24.5923
R106 VP.n53 VP.n51 24.5923
R107 VP.n57 VP.n21 24.5923
R108 VP.n58 VP.n57 24.5923
R109 VP.n59 VP.n58 24.5923
R110 VP.n39 VP.n38 24.5923
R111 VP.n40 VP.n39 24.5923
R112 VP.n40 VP.n25 24.5923
R113 VP.n44 VP.n25 24.5923
R114 VP.n45 VP.n44 24.5923
R115 VP.n46 VP.n45 24.5923
R116 VP.n33 VP.n32 24.5923
R117 VP.n34 VP.n33 24.5923
R118 VP.n83 VP.n12 18.1985
R119 VP.n104 VP.n103 18.1985
R120 VP.n53 VP.n52 18.1985
R121 VP.n32 VP.n29 18.1985
R122 VP.n68 VP.n16 11.8046
R123 VP.n116 VP.n0 11.8046
R124 VP.n65 VP.n17 11.8046
R125 VP.n80 VP.n12 6.39438
R126 VP.n103 VP.n4 6.39438
R127 VP.n52 VP.n21 6.39438
R128 VP.n31 VP.n30 3.08735
R129 VP.n67 VP.n66 0.354861
R130 VP.n70 VP.n69 0.354861
R131 VP.n118 VP.n117 0.354861
R132 VP VP.n118 0.267071
R133 VP.n31 VP.n28 0.189894
R134 VP.n35 VP.n28 0.189894
R135 VP.n36 VP.n35 0.189894
R136 VP.n37 VP.n36 0.189894
R137 VP.n37 VP.n26 0.189894
R138 VP.n41 VP.n26 0.189894
R139 VP.n42 VP.n41 0.189894
R140 VP.n43 VP.n42 0.189894
R141 VP.n43 VP.n24 0.189894
R142 VP.n47 VP.n24 0.189894
R143 VP.n48 VP.n47 0.189894
R144 VP.n49 VP.n48 0.189894
R145 VP.n49 VP.n22 0.189894
R146 VP.n54 VP.n22 0.189894
R147 VP.n55 VP.n54 0.189894
R148 VP.n56 VP.n55 0.189894
R149 VP.n56 VP.n20 0.189894
R150 VP.n60 VP.n20 0.189894
R151 VP.n61 VP.n60 0.189894
R152 VP.n62 VP.n61 0.189894
R153 VP.n62 VP.n18 0.189894
R154 VP.n66 VP.n18 0.189894
R155 VP.n71 VP.n70 0.189894
R156 VP.n71 VP.n15 0.189894
R157 VP.n75 VP.n15 0.189894
R158 VP.n76 VP.n75 0.189894
R159 VP.n77 VP.n76 0.189894
R160 VP.n77 VP.n13 0.189894
R161 VP.n81 VP.n13 0.189894
R162 VP.n82 VP.n81 0.189894
R163 VP.n82 VP.n11 0.189894
R164 VP.n86 VP.n11 0.189894
R165 VP.n87 VP.n86 0.189894
R166 VP.n88 VP.n87 0.189894
R167 VP.n88 VP.n9 0.189894
R168 VP.n92 VP.n9 0.189894
R169 VP.n93 VP.n92 0.189894
R170 VP.n94 VP.n93 0.189894
R171 VP.n94 VP.n7 0.189894
R172 VP.n98 VP.n7 0.189894
R173 VP.n99 VP.n98 0.189894
R174 VP.n100 VP.n99 0.189894
R175 VP.n100 VP.n5 0.189894
R176 VP.n105 VP.n5 0.189894
R177 VP.n106 VP.n105 0.189894
R178 VP.n107 VP.n106 0.189894
R179 VP.n107 VP.n3 0.189894
R180 VP.n111 VP.n3 0.189894
R181 VP.n112 VP.n111 0.189894
R182 VP.n113 VP.n112 0.189894
R183 VP.n113 VP.n1 0.189894
R184 VP.n117 VP.n1 0.189894
R185 VDD1.n48 VDD1.n0 289.615
R186 VDD1.n103 VDD1.n55 289.615
R187 VDD1.n49 VDD1.n48 185
R188 VDD1.n47 VDD1.n46 185
R189 VDD1.n4 VDD1.n3 185
R190 VDD1.n41 VDD1.n40 185
R191 VDD1.n39 VDD1.n6 185
R192 VDD1.n38 VDD1.n37 185
R193 VDD1.n9 VDD1.n7 185
R194 VDD1.n32 VDD1.n31 185
R195 VDD1.n30 VDD1.n29 185
R196 VDD1.n13 VDD1.n12 185
R197 VDD1.n24 VDD1.n23 185
R198 VDD1.n22 VDD1.n21 185
R199 VDD1.n17 VDD1.n16 185
R200 VDD1.n71 VDD1.n70 185
R201 VDD1.n76 VDD1.n75 185
R202 VDD1.n78 VDD1.n77 185
R203 VDD1.n67 VDD1.n66 185
R204 VDD1.n84 VDD1.n83 185
R205 VDD1.n86 VDD1.n85 185
R206 VDD1.n63 VDD1.n62 185
R207 VDD1.n93 VDD1.n92 185
R208 VDD1.n94 VDD1.n61 185
R209 VDD1.n96 VDD1.n95 185
R210 VDD1.n59 VDD1.n58 185
R211 VDD1.n102 VDD1.n101 185
R212 VDD1.n104 VDD1.n103 185
R213 VDD1.n18 VDD1.t2 149.524
R214 VDD1.n72 VDD1.t5 149.524
R215 VDD1.n48 VDD1.n47 104.615
R216 VDD1.n47 VDD1.n3 104.615
R217 VDD1.n40 VDD1.n3 104.615
R218 VDD1.n40 VDD1.n39 104.615
R219 VDD1.n39 VDD1.n38 104.615
R220 VDD1.n38 VDD1.n7 104.615
R221 VDD1.n31 VDD1.n7 104.615
R222 VDD1.n31 VDD1.n30 104.615
R223 VDD1.n30 VDD1.n12 104.615
R224 VDD1.n23 VDD1.n12 104.615
R225 VDD1.n23 VDD1.n22 104.615
R226 VDD1.n22 VDD1.n16 104.615
R227 VDD1.n76 VDD1.n70 104.615
R228 VDD1.n77 VDD1.n76 104.615
R229 VDD1.n77 VDD1.n66 104.615
R230 VDD1.n84 VDD1.n66 104.615
R231 VDD1.n85 VDD1.n84 104.615
R232 VDD1.n85 VDD1.n62 104.615
R233 VDD1.n93 VDD1.n62 104.615
R234 VDD1.n94 VDD1.n93 104.615
R235 VDD1.n95 VDD1.n94 104.615
R236 VDD1.n95 VDD1.n58 104.615
R237 VDD1.n102 VDD1.n58 104.615
R238 VDD1.n103 VDD1.n102 104.615
R239 VDD1.n111 VDD1.n110 66.2506
R240 VDD1.n54 VDD1.n53 63.804
R241 VDD1.n113 VDD1.n112 63.8038
R242 VDD1.n109 VDD1.n108 63.8038
R243 VDD1.n54 VDD1.n52 53.364
R244 VDD1.n109 VDD1.n107 53.364
R245 VDD1.t2 VDD1.n16 52.3082
R246 VDD1.t5 VDD1.n70 52.3082
R247 VDD1.n113 VDD1.n111 50.4513
R248 VDD1.n41 VDD1.n6 13.1884
R249 VDD1.n96 VDD1.n61 13.1884
R250 VDD1.n42 VDD1.n4 12.8005
R251 VDD1.n37 VDD1.n8 12.8005
R252 VDD1.n92 VDD1.n91 12.8005
R253 VDD1.n97 VDD1.n59 12.8005
R254 VDD1.n46 VDD1.n45 12.0247
R255 VDD1.n36 VDD1.n9 12.0247
R256 VDD1.n90 VDD1.n63 12.0247
R257 VDD1.n101 VDD1.n100 12.0247
R258 VDD1.n49 VDD1.n2 11.249
R259 VDD1.n33 VDD1.n32 11.249
R260 VDD1.n87 VDD1.n86 11.249
R261 VDD1.n104 VDD1.n57 11.249
R262 VDD1.n50 VDD1.n0 10.4732
R263 VDD1.n29 VDD1.n11 10.4732
R264 VDD1.n83 VDD1.n65 10.4732
R265 VDD1.n105 VDD1.n55 10.4732
R266 VDD1.n18 VDD1.n17 10.2747
R267 VDD1.n72 VDD1.n71 10.2747
R268 VDD1.n28 VDD1.n13 9.69747
R269 VDD1.n82 VDD1.n67 9.69747
R270 VDD1.n52 VDD1.n51 9.45567
R271 VDD1.n107 VDD1.n106 9.45567
R272 VDD1.n20 VDD1.n19 9.3005
R273 VDD1.n15 VDD1.n14 9.3005
R274 VDD1.n26 VDD1.n25 9.3005
R275 VDD1.n28 VDD1.n27 9.3005
R276 VDD1.n11 VDD1.n10 9.3005
R277 VDD1.n34 VDD1.n33 9.3005
R278 VDD1.n36 VDD1.n35 9.3005
R279 VDD1.n8 VDD1.n5 9.3005
R280 VDD1.n51 VDD1.n50 9.3005
R281 VDD1.n2 VDD1.n1 9.3005
R282 VDD1.n45 VDD1.n44 9.3005
R283 VDD1.n43 VDD1.n42 9.3005
R284 VDD1.n106 VDD1.n105 9.3005
R285 VDD1.n57 VDD1.n56 9.3005
R286 VDD1.n100 VDD1.n99 9.3005
R287 VDD1.n98 VDD1.n97 9.3005
R288 VDD1.n74 VDD1.n73 9.3005
R289 VDD1.n69 VDD1.n68 9.3005
R290 VDD1.n80 VDD1.n79 9.3005
R291 VDD1.n82 VDD1.n81 9.3005
R292 VDD1.n65 VDD1.n64 9.3005
R293 VDD1.n88 VDD1.n87 9.3005
R294 VDD1.n90 VDD1.n89 9.3005
R295 VDD1.n91 VDD1.n60 9.3005
R296 VDD1.n25 VDD1.n24 8.92171
R297 VDD1.n79 VDD1.n78 8.92171
R298 VDD1.n21 VDD1.n15 8.14595
R299 VDD1.n75 VDD1.n69 8.14595
R300 VDD1.n20 VDD1.n17 7.3702
R301 VDD1.n74 VDD1.n71 7.3702
R302 VDD1.n21 VDD1.n20 5.81868
R303 VDD1.n75 VDD1.n74 5.81868
R304 VDD1.n24 VDD1.n15 5.04292
R305 VDD1.n78 VDD1.n69 5.04292
R306 VDD1.n25 VDD1.n13 4.26717
R307 VDD1.n79 VDD1.n67 4.26717
R308 VDD1.n52 VDD1.n0 3.49141
R309 VDD1.n29 VDD1.n28 3.49141
R310 VDD1.n83 VDD1.n82 3.49141
R311 VDD1.n107 VDD1.n55 3.49141
R312 VDD1.n19 VDD1.n18 2.84303
R313 VDD1.n73 VDD1.n72 2.84303
R314 VDD1.n50 VDD1.n49 2.71565
R315 VDD1.n32 VDD1.n11 2.71565
R316 VDD1.n86 VDD1.n65 2.71565
R317 VDD1.n105 VDD1.n104 2.71565
R318 VDD1 VDD1.n113 2.44447
R319 VDD1.n112 VDD1.t7 1.97655
R320 VDD1.n112 VDD1.t6 1.97655
R321 VDD1.n53 VDD1.t4 1.97655
R322 VDD1.n53 VDD1.t3 1.97655
R323 VDD1.n110 VDD1.t1 1.97655
R324 VDD1.n110 VDD1.t8 1.97655
R325 VDD1.n108 VDD1.t9 1.97655
R326 VDD1.n108 VDD1.t0 1.97655
R327 VDD1.n46 VDD1.n2 1.93989
R328 VDD1.n33 VDD1.n9 1.93989
R329 VDD1.n87 VDD1.n63 1.93989
R330 VDD1.n101 VDD1.n57 1.93989
R331 VDD1.n45 VDD1.n4 1.16414
R332 VDD1.n37 VDD1.n36 1.16414
R333 VDD1.n92 VDD1.n90 1.16414
R334 VDD1.n100 VDD1.n59 1.16414
R335 VDD1 VDD1.n54 0.892741
R336 VDD1.n111 VDD1.n109 0.779206
R337 VDD1.n42 VDD1.n41 0.388379
R338 VDD1.n8 VDD1.n6 0.388379
R339 VDD1.n91 VDD1.n61 0.388379
R340 VDD1.n97 VDD1.n96 0.388379
R341 VDD1.n51 VDD1.n1 0.155672
R342 VDD1.n44 VDD1.n1 0.155672
R343 VDD1.n44 VDD1.n43 0.155672
R344 VDD1.n43 VDD1.n5 0.155672
R345 VDD1.n35 VDD1.n5 0.155672
R346 VDD1.n35 VDD1.n34 0.155672
R347 VDD1.n34 VDD1.n10 0.155672
R348 VDD1.n27 VDD1.n10 0.155672
R349 VDD1.n27 VDD1.n26 0.155672
R350 VDD1.n26 VDD1.n14 0.155672
R351 VDD1.n19 VDD1.n14 0.155672
R352 VDD1.n73 VDD1.n68 0.155672
R353 VDD1.n80 VDD1.n68 0.155672
R354 VDD1.n81 VDD1.n80 0.155672
R355 VDD1.n81 VDD1.n64 0.155672
R356 VDD1.n88 VDD1.n64 0.155672
R357 VDD1.n89 VDD1.n88 0.155672
R358 VDD1.n89 VDD1.n60 0.155672
R359 VDD1.n98 VDD1.n60 0.155672
R360 VDD1.n99 VDD1.n98 0.155672
R361 VDD1.n99 VDD1.n56 0.155672
R362 VDD1.n106 VDD1.n56 0.155672
R363 VTAIL.n224 VTAIL.n176 289.615
R364 VTAIL.n50 VTAIL.n2 289.615
R365 VTAIL.n170 VTAIL.n122 289.615
R366 VTAIL.n112 VTAIL.n64 289.615
R367 VTAIL.n192 VTAIL.n191 185
R368 VTAIL.n197 VTAIL.n196 185
R369 VTAIL.n199 VTAIL.n198 185
R370 VTAIL.n188 VTAIL.n187 185
R371 VTAIL.n205 VTAIL.n204 185
R372 VTAIL.n207 VTAIL.n206 185
R373 VTAIL.n184 VTAIL.n183 185
R374 VTAIL.n214 VTAIL.n213 185
R375 VTAIL.n215 VTAIL.n182 185
R376 VTAIL.n217 VTAIL.n216 185
R377 VTAIL.n180 VTAIL.n179 185
R378 VTAIL.n223 VTAIL.n222 185
R379 VTAIL.n225 VTAIL.n224 185
R380 VTAIL.n18 VTAIL.n17 185
R381 VTAIL.n23 VTAIL.n22 185
R382 VTAIL.n25 VTAIL.n24 185
R383 VTAIL.n14 VTAIL.n13 185
R384 VTAIL.n31 VTAIL.n30 185
R385 VTAIL.n33 VTAIL.n32 185
R386 VTAIL.n10 VTAIL.n9 185
R387 VTAIL.n40 VTAIL.n39 185
R388 VTAIL.n41 VTAIL.n8 185
R389 VTAIL.n43 VTAIL.n42 185
R390 VTAIL.n6 VTAIL.n5 185
R391 VTAIL.n49 VTAIL.n48 185
R392 VTAIL.n51 VTAIL.n50 185
R393 VTAIL.n171 VTAIL.n170 185
R394 VTAIL.n169 VTAIL.n168 185
R395 VTAIL.n126 VTAIL.n125 185
R396 VTAIL.n163 VTAIL.n162 185
R397 VTAIL.n161 VTAIL.n128 185
R398 VTAIL.n160 VTAIL.n159 185
R399 VTAIL.n131 VTAIL.n129 185
R400 VTAIL.n154 VTAIL.n153 185
R401 VTAIL.n152 VTAIL.n151 185
R402 VTAIL.n135 VTAIL.n134 185
R403 VTAIL.n146 VTAIL.n145 185
R404 VTAIL.n144 VTAIL.n143 185
R405 VTAIL.n139 VTAIL.n138 185
R406 VTAIL.n113 VTAIL.n112 185
R407 VTAIL.n111 VTAIL.n110 185
R408 VTAIL.n68 VTAIL.n67 185
R409 VTAIL.n105 VTAIL.n104 185
R410 VTAIL.n103 VTAIL.n70 185
R411 VTAIL.n102 VTAIL.n101 185
R412 VTAIL.n73 VTAIL.n71 185
R413 VTAIL.n96 VTAIL.n95 185
R414 VTAIL.n94 VTAIL.n93 185
R415 VTAIL.n77 VTAIL.n76 185
R416 VTAIL.n88 VTAIL.n87 185
R417 VTAIL.n86 VTAIL.n85 185
R418 VTAIL.n81 VTAIL.n80 185
R419 VTAIL.n193 VTAIL.t8 149.524
R420 VTAIL.n19 VTAIL.t13 149.524
R421 VTAIL.n140 VTAIL.t17 149.524
R422 VTAIL.n82 VTAIL.t6 149.524
R423 VTAIL.n197 VTAIL.n191 104.615
R424 VTAIL.n198 VTAIL.n197 104.615
R425 VTAIL.n198 VTAIL.n187 104.615
R426 VTAIL.n205 VTAIL.n187 104.615
R427 VTAIL.n206 VTAIL.n205 104.615
R428 VTAIL.n206 VTAIL.n183 104.615
R429 VTAIL.n214 VTAIL.n183 104.615
R430 VTAIL.n215 VTAIL.n214 104.615
R431 VTAIL.n216 VTAIL.n215 104.615
R432 VTAIL.n216 VTAIL.n179 104.615
R433 VTAIL.n223 VTAIL.n179 104.615
R434 VTAIL.n224 VTAIL.n223 104.615
R435 VTAIL.n23 VTAIL.n17 104.615
R436 VTAIL.n24 VTAIL.n23 104.615
R437 VTAIL.n24 VTAIL.n13 104.615
R438 VTAIL.n31 VTAIL.n13 104.615
R439 VTAIL.n32 VTAIL.n31 104.615
R440 VTAIL.n32 VTAIL.n9 104.615
R441 VTAIL.n40 VTAIL.n9 104.615
R442 VTAIL.n41 VTAIL.n40 104.615
R443 VTAIL.n42 VTAIL.n41 104.615
R444 VTAIL.n42 VTAIL.n5 104.615
R445 VTAIL.n49 VTAIL.n5 104.615
R446 VTAIL.n50 VTAIL.n49 104.615
R447 VTAIL.n170 VTAIL.n169 104.615
R448 VTAIL.n169 VTAIL.n125 104.615
R449 VTAIL.n162 VTAIL.n125 104.615
R450 VTAIL.n162 VTAIL.n161 104.615
R451 VTAIL.n161 VTAIL.n160 104.615
R452 VTAIL.n160 VTAIL.n129 104.615
R453 VTAIL.n153 VTAIL.n129 104.615
R454 VTAIL.n153 VTAIL.n152 104.615
R455 VTAIL.n152 VTAIL.n134 104.615
R456 VTAIL.n145 VTAIL.n134 104.615
R457 VTAIL.n145 VTAIL.n144 104.615
R458 VTAIL.n144 VTAIL.n138 104.615
R459 VTAIL.n112 VTAIL.n111 104.615
R460 VTAIL.n111 VTAIL.n67 104.615
R461 VTAIL.n104 VTAIL.n67 104.615
R462 VTAIL.n104 VTAIL.n103 104.615
R463 VTAIL.n103 VTAIL.n102 104.615
R464 VTAIL.n102 VTAIL.n71 104.615
R465 VTAIL.n95 VTAIL.n71 104.615
R466 VTAIL.n95 VTAIL.n94 104.615
R467 VTAIL.n94 VTAIL.n76 104.615
R468 VTAIL.n87 VTAIL.n76 104.615
R469 VTAIL.n87 VTAIL.n86 104.615
R470 VTAIL.n86 VTAIL.n80 104.615
R471 VTAIL.t8 VTAIL.n191 52.3082
R472 VTAIL.t13 VTAIL.n17 52.3082
R473 VTAIL.t17 VTAIL.n138 52.3082
R474 VTAIL.t6 VTAIL.n80 52.3082
R475 VTAIL.n121 VTAIL.n120 47.1252
R476 VTAIL.n119 VTAIL.n118 47.1252
R477 VTAIL.n63 VTAIL.n62 47.1252
R478 VTAIL.n61 VTAIL.n60 47.1252
R479 VTAIL.n231 VTAIL.n230 47.125
R480 VTAIL.n1 VTAIL.n0 47.125
R481 VTAIL.n57 VTAIL.n56 47.125
R482 VTAIL.n59 VTAIL.n58 47.125
R483 VTAIL.n229 VTAIL.n228 33.349
R484 VTAIL.n55 VTAIL.n54 33.349
R485 VTAIL.n175 VTAIL.n174 33.349
R486 VTAIL.n117 VTAIL.n116 33.349
R487 VTAIL.n61 VTAIL.n59 27.6772
R488 VTAIL.n229 VTAIL.n175 24.341
R489 VTAIL.n217 VTAIL.n182 13.1884
R490 VTAIL.n43 VTAIL.n8 13.1884
R491 VTAIL.n163 VTAIL.n128 13.1884
R492 VTAIL.n105 VTAIL.n70 13.1884
R493 VTAIL.n213 VTAIL.n212 12.8005
R494 VTAIL.n218 VTAIL.n180 12.8005
R495 VTAIL.n39 VTAIL.n38 12.8005
R496 VTAIL.n44 VTAIL.n6 12.8005
R497 VTAIL.n164 VTAIL.n126 12.8005
R498 VTAIL.n159 VTAIL.n130 12.8005
R499 VTAIL.n106 VTAIL.n68 12.8005
R500 VTAIL.n101 VTAIL.n72 12.8005
R501 VTAIL.n211 VTAIL.n184 12.0247
R502 VTAIL.n222 VTAIL.n221 12.0247
R503 VTAIL.n37 VTAIL.n10 12.0247
R504 VTAIL.n48 VTAIL.n47 12.0247
R505 VTAIL.n168 VTAIL.n167 12.0247
R506 VTAIL.n158 VTAIL.n131 12.0247
R507 VTAIL.n110 VTAIL.n109 12.0247
R508 VTAIL.n100 VTAIL.n73 12.0247
R509 VTAIL.n208 VTAIL.n207 11.249
R510 VTAIL.n225 VTAIL.n178 11.249
R511 VTAIL.n34 VTAIL.n33 11.249
R512 VTAIL.n51 VTAIL.n4 11.249
R513 VTAIL.n171 VTAIL.n124 11.249
R514 VTAIL.n155 VTAIL.n154 11.249
R515 VTAIL.n113 VTAIL.n66 11.249
R516 VTAIL.n97 VTAIL.n96 11.249
R517 VTAIL.n204 VTAIL.n186 10.4732
R518 VTAIL.n226 VTAIL.n176 10.4732
R519 VTAIL.n30 VTAIL.n12 10.4732
R520 VTAIL.n52 VTAIL.n2 10.4732
R521 VTAIL.n172 VTAIL.n122 10.4732
R522 VTAIL.n151 VTAIL.n133 10.4732
R523 VTAIL.n114 VTAIL.n64 10.4732
R524 VTAIL.n93 VTAIL.n75 10.4732
R525 VTAIL.n193 VTAIL.n192 10.2747
R526 VTAIL.n19 VTAIL.n18 10.2747
R527 VTAIL.n140 VTAIL.n139 10.2747
R528 VTAIL.n82 VTAIL.n81 10.2747
R529 VTAIL.n203 VTAIL.n188 9.69747
R530 VTAIL.n29 VTAIL.n14 9.69747
R531 VTAIL.n150 VTAIL.n135 9.69747
R532 VTAIL.n92 VTAIL.n77 9.69747
R533 VTAIL.n228 VTAIL.n227 9.45567
R534 VTAIL.n54 VTAIL.n53 9.45567
R535 VTAIL.n174 VTAIL.n173 9.45567
R536 VTAIL.n116 VTAIL.n115 9.45567
R537 VTAIL.n227 VTAIL.n226 9.3005
R538 VTAIL.n178 VTAIL.n177 9.3005
R539 VTAIL.n221 VTAIL.n220 9.3005
R540 VTAIL.n219 VTAIL.n218 9.3005
R541 VTAIL.n195 VTAIL.n194 9.3005
R542 VTAIL.n190 VTAIL.n189 9.3005
R543 VTAIL.n201 VTAIL.n200 9.3005
R544 VTAIL.n203 VTAIL.n202 9.3005
R545 VTAIL.n186 VTAIL.n185 9.3005
R546 VTAIL.n209 VTAIL.n208 9.3005
R547 VTAIL.n211 VTAIL.n210 9.3005
R548 VTAIL.n212 VTAIL.n181 9.3005
R549 VTAIL.n53 VTAIL.n52 9.3005
R550 VTAIL.n4 VTAIL.n3 9.3005
R551 VTAIL.n47 VTAIL.n46 9.3005
R552 VTAIL.n45 VTAIL.n44 9.3005
R553 VTAIL.n21 VTAIL.n20 9.3005
R554 VTAIL.n16 VTAIL.n15 9.3005
R555 VTAIL.n27 VTAIL.n26 9.3005
R556 VTAIL.n29 VTAIL.n28 9.3005
R557 VTAIL.n12 VTAIL.n11 9.3005
R558 VTAIL.n35 VTAIL.n34 9.3005
R559 VTAIL.n37 VTAIL.n36 9.3005
R560 VTAIL.n38 VTAIL.n7 9.3005
R561 VTAIL.n142 VTAIL.n141 9.3005
R562 VTAIL.n137 VTAIL.n136 9.3005
R563 VTAIL.n148 VTAIL.n147 9.3005
R564 VTAIL.n150 VTAIL.n149 9.3005
R565 VTAIL.n133 VTAIL.n132 9.3005
R566 VTAIL.n156 VTAIL.n155 9.3005
R567 VTAIL.n158 VTAIL.n157 9.3005
R568 VTAIL.n130 VTAIL.n127 9.3005
R569 VTAIL.n173 VTAIL.n172 9.3005
R570 VTAIL.n124 VTAIL.n123 9.3005
R571 VTAIL.n167 VTAIL.n166 9.3005
R572 VTAIL.n165 VTAIL.n164 9.3005
R573 VTAIL.n84 VTAIL.n83 9.3005
R574 VTAIL.n79 VTAIL.n78 9.3005
R575 VTAIL.n90 VTAIL.n89 9.3005
R576 VTAIL.n92 VTAIL.n91 9.3005
R577 VTAIL.n75 VTAIL.n74 9.3005
R578 VTAIL.n98 VTAIL.n97 9.3005
R579 VTAIL.n100 VTAIL.n99 9.3005
R580 VTAIL.n72 VTAIL.n69 9.3005
R581 VTAIL.n115 VTAIL.n114 9.3005
R582 VTAIL.n66 VTAIL.n65 9.3005
R583 VTAIL.n109 VTAIL.n108 9.3005
R584 VTAIL.n107 VTAIL.n106 9.3005
R585 VTAIL.n200 VTAIL.n199 8.92171
R586 VTAIL.n26 VTAIL.n25 8.92171
R587 VTAIL.n147 VTAIL.n146 8.92171
R588 VTAIL.n89 VTAIL.n88 8.92171
R589 VTAIL.n196 VTAIL.n190 8.14595
R590 VTAIL.n22 VTAIL.n16 8.14595
R591 VTAIL.n143 VTAIL.n137 8.14595
R592 VTAIL.n85 VTAIL.n79 8.14595
R593 VTAIL.n195 VTAIL.n192 7.3702
R594 VTAIL.n21 VTAIL.n18 7.3702
R595 VTAIL.n142 VTAIL.n139 7.3702
R596 VTAIL.n84 VTAIL.n81 7.3702
R597 VTAIL.n196 VTAIL.n195 5.81868
R598 VTAIL.n22 VTAIL.n21 5.81868
R599 VTAIL.n143 VTAIL.n142 5.81868
R600 VTAIL.n85 VTAIL.n84 5.81868
R601 VTAIL.n199 VTAIL.n190 5.04292
R602 VTAIL.n25 VTAIL.n16 5.04292
R603 VTAIL.n146 VTAIL.n137 5.04292
R604 VTAIL.n88 VTAIL.n79 5.04292
R605 VTAIL.n200 VTAIL.n188 4.26717
R606 VTAIL.n26 VTAIL.n14 4.26717
R607 VTAIL.n147 VTAIL.n135 4.26717
R608 VTAIL.n89 VTAIL.n77 4.26717
R609 VTAIL.n204 VTAIL.n203 3.49141
R610 VTAIL.n228 VTAIL.n176 3.49141
R611 VTAIL.n30 VTAIL.n29 3.49141
R612 VTAIL.n54 VTAIL.n2 3.49141
R613 VTAIL.n174 VTAIL.n122 3.49141
R614 VTAIL.n151 VTAIL.n150 3.49141
R615 VTAIL.n116 VTAIL.n64 3.49141
R616 VTAIL.n93 VTAIL.n92 3.49141
R617 VTAIL.n63 VTAIL.n61 3.33671
R618 VTAIL.n117 VTAIL.n63 3.33671
R619 VTAIL.n121 VTAIL.n119 3.33671
R620 VTAIL.n175 VTAIL.n121 3.33671
R621 VTAIL.n59 VTAIL.n57 3.33671
R622 VTAIL.n57 VTAIL.n55 3.33671
R623 VTAIL.n231 VTAIL.n229 3.33671
R624 VTAIL.n194 VTAIL.n193 2.84303
R625 VTAIL.n20 VTAIL.n19 2.84303
R626 VTAIL.n141 VTAIL.n140 2.84303
R627 VTAIL.n83 VTAIL.n82 2.84303
R628 VTAIL.n207 VTAIL.n186 2.71565
R629 VTAIL.n226 VTAIL.n225 2.71565
R630 VTAIL.n33 VTAIL.n12 2.71565
R631 VTAIL.n52 VTAIL.n51 2.71565
R632 VTAIL.n172 VTAIL.n171 2.71565
R633 VTAIL.n154 VTAIL.n133 2.71565
R634 VTAIL.n114 VTAIL.n113 2.71565
R635 VTAIL.n96 VTAIL.n75 2.71565
R636 VTAIL VTAIL.n1 2.56084
R637 VTAIL.n119 VTAIL.n117 2.13843
R638 VTAIL.n55 VTAIL.n1 2.13843
R639 VTAIL.n230 VTAIL.t5 1.97655
R640 VTAIL.n230 VTAIL.t3 1.97655
R641 VTAIL.n0 VTAIL.t2 1.97655
R642 VTAIL.n0 VTAIL.t4 1.97655
R643 VTAIL.n56 VTAIL.t15 1.97655
R644 VTAIL.n56 VTAIL.t16 1.97655
R645 VTAIL.n58 VTAIL.t12 1.97655
R646 VTAIL.n58 VTAIL.t19 1.97655
R647 VTAIL.n120 VTAIL.t14 1.97655
R648 VTAIL.n120 VTAIL.t18 1.97655
R649 VTAIL.n118 VTAIL.t10 1.97655
R650 VTAIL.n118 VTAIL.t11 1.97655
R651 VTAIL.n62 VTAIL.t1 1.97655
R652 VTAIL.n62 VTAIL.t0 1.97655
R653 VTAIL.n60 VTAIL.t7 1.97655
R654 VTAIL.n60 VTAIL.t9 1.97655
R655 VTAIL.n208 VTAIL.n184 1.93989
R656 VTAIL.n222 VTAIL.n178 1.93989
R657 VTAIL.n34 VTAIL.n10 1.93989
R658 VTAIL.n48 VTAIL.n4 1.93989
R659 VTAIL.n168 VTAIL.n124 1.93989
R660 VTAIL.n155 VTAIL.n131 1.93989
R661 VTAIL.n110 VTAIL.n66 1.93989
R662 VTAIL.n97 VTAIL.n73 1.93989
R663 VTAIL.n213 VTAIL.n211 1.16414
R664 VTAIL.n221 VTAIL.n180 1.16414
R665 VTAIL.n39 VTAIL.n37 1.16414
R666 VTAIL.n47 VTAIL.n6 1.16414
R667 VTAIL.n167 VTAIL.n126 1.16414
R668 VTAIL.n159 VTAIL.n158 1.16414
R669 VTAIL.n109 VTAIL.n68 1.16414
R670 VTAIL.n101 VTAIL.n100 1.16414
R671 VTAIL VTAIL.n231 0.776362
R672 VTAIL.n212 VTAIL.n182 0.388379
R673 VTAIL.n218 VTAIL.n217 0.388379
R674 VTAIL.n38 VTAIL.n8 0.388379
R675 VTAIL.n44 VTAIL.n43 0.388379
R676 VTAIL.n164 VTAIL.n163 0.388379
R677 VTAIL.n130 VTAIL.n128 0.388379
R678 VTAIL.n106 VTAIL.n105 0.388379
R679 VTAIL.n72 VTAIL.n70 0.388379
R680 VTAIL.n194 VTAIL.n189 0.155672
R681 VTAIL.n201 VTAIL.n189 0.155672
R682 VTAIL.n202 VTAIL.n201 0.155672
R683 VTAIL.n202 VTAIL.n185 0.155672
R684 VTAIL.n209 VTAIL.n185 0.155672
R685 VTAIL.n210 VTAIL.n209 0.155672
R686 VTAIL.n210 VTAIL.n181 0.155672
R687 VTAIL.n219 VTAIL.n181 0.155672
R688 VTAIL.n220 VTAIL.n219 0.155672
R689 VTAIL.n220 VTAIL.n177 0.155672
R690 VTAIL.n227 VTAIL.n177 0.155672
R691 VTAIL.n20 VTAIL.n15 0.155672
R692 VTAIL.n27 VTAIL.n15 0.155672
R693 VTAIL.n28 VTAIL.n27 0.155672
R694 VTAIL.n28 VTAIL.n11 0.155672
R695 VTAIL.n35 VTAIL.n11 0.155672
R696 VTAIL.n36 VTAIL.n35 0.155672
R697 VTAIL.n36 VTAIL.n7 0.155672
R698 VTAIL.n45 VTAIL.n7 0.155672
R699 VTAIL.n46 VTAIL.n45 0.155672
R700 VTAIL.n46 VTAIL.n3 0.155672
R701 VTAIL.n53 VTAIL.n3 0.155672
R702 VTAIL.n173 VTAIL.n123 0.155672
R703 VTAIL.n166 VTAIL.n123 0.155672
R704 VTAIL.n166 VTAIL.n165 0.155672
R705 VTAIL.n165 VTAIL.n127 0.155672
R706 VTAIL.n157 VTAIL.n127 0.155672
R707 VTAIL.n157 VTAIL.n156 0.155672
R708 VTAIL.n156 VTAIL.n132 0.155672
R709 VTAIL.n149 VTAIL.n132 0.155672
R710 VTAIL.n149 VTAIL.n148 0.155672
R711 VTAIL.n148 VTAIL.n136 0.155672
R712 VTAIL.n141 VTAIL.n136 0.155672
R713 VTAIL.n115 VTAIL.n65 0.155672
R714 VTAIL.n108 VTAIL.n65 0.155672
R715 VTAIL.n108 VTAIL.n107 0.155672
R716 VTAIL.n107 VTAIL.n69 0.155672
R717 VTAIL.n99 VTAIL.n69 0.155672
R718 VTAIL.n99 VTAIL.n98 0.155672
R719 VTAIL.n98 VTAIL.n74 0.155672
R720 VTAIL.n91 VTAIL.n74 0.155672
R721 VTAIL.n91 VTAIL.n90 0.155672
R722 VTAIL.n90 VTAIL.n78 0.155672
R723 VTAIL.n83 VTAIL.n78 0.155672
R724 B.n1029 B.n1028 585
R725 B.n1030 B.n1029 585
R726 B.n343 B.n180 585
R727 B.n342 B.n341 585
R728 B.n340 B.n339 585
R729 B.n338 B.n337 585
R730 B.n336 B.n335 585
R731 B.n334 B.n333 585
R732 B.n332 B.n331 585
R733 B.n330 B.n329 585
R734 B.n328 B.n327 585
R735 B.n326 B.n325 585
R736 B.n324 B.n323 585
R737 B.n322 B.n321 585
R738 B.n320 B.n319 585
R739 B.n318 B.n317 585
R740 B.n316 B.n315 585
R741 B.n314 B.n313 585
R742 B.n312 B.n311 585
R743 B.n310 B.n309 585
R744 B.n308 B.n307 585
R745 B.n306 B.n305 585
R746 B.n304 B.n303 585
R747 B.n302 B.n301 585
R748 B.n300 B.n299 585
R749 B.n298 B.n297 585
R750 B.n296 B.n295 585
R751 B.n294 B.n293 585
R752 B.n292 B.n291 585
R753 B.n290 B.n289 585
R754 B.n288 B.n287 585
R755 B.n286 B.n285 585
R756 B.n284 B.n283 585
R757 B.n282 B.n281 585
R758 B.n280 B.n279 585
R759 B.n278 B.n277 585
R760 B.n276 B.n275 585
R761 B.n273 B.n272 585
R762 B.n271 B.n270 585
R763 B.n269 B.n268 585
R764 B.n267 B.n266 585
R765 B.n265 B.n264 585
R766 B.n263 B.n262 585
R767 B.n261 B.n260 585
R768 B.n259 B.n258 585
R769 B.n257 B.n256 585
R770 B.n255 B.n254 585
R771 B.n253 B.n252 585
R772 B.n251 B.n250 585
R773 B.n249 B.n248 585
R774 B.n247 B.n246 585
R775 B.n245 B.n244 585
R776 B.n243 B.n242 585
R777 B.n241 B.n240 585
R778 B.n239 B.n238 585
R779 B.n237 B.n236 585
R780 B.n235 B.n234 585
R781 B.n233 B.n232 585
R782 B.n231 B.n230 585
R783 B.n229 B.n228 585
R784 B.n227 B.n226 585
R785 B.n225 B.n224 585
R786 B.n223 B.n222 585
R787 B.n221 B.n220 585
R788 B.n219 B.n218 585
R789 B.n217 B.n216 585
R790 B.n215 B.n214 585
R791 B.n213 B.n212 585
R792 B.n211 B.n210 585
R793 B.n209 B.n208 585
R794 B.n207 B.n206 585
R795 B.n205 B.n204 585
R796 B.n203 B.n202 585
R797 B.n201 B.n200 585
R798 B.n199 B.n198 585
R799 B.n197 B.n196 585
R800 B.n195 B.n194 585
R801 B.n193 B.n192 585
R802 B.n191 B.n190 585
R803 B.n189 B.n188 585
R804 B.n187 B.n186 585
R805 B.n138 B.n137 585
R806 B.n1027 B.n139 585
R807 B.n1031 B.n139 585
R808 B.n1026 B.n1025 585
R809 B.n1025 B.n135 585
R810 B.n1024 B.n134 585
R811 B.n1037 B.n134 585
R812 B.n1023 B.n133 585
R813 B.n1038 B.n133 585
R814 B.n1022 B.n132 585
R815 B.n1039 B.n132 585
R816 B.n1021 B.n1020 585
R817 B.n1020 B.n128 585
R818 B.n1019 B.n127 585
R819 B.n1045 B.n127 585
R820 B.n1018 B.n126 585
R821 B.n1046 B.n126 585
R822 B.n1017 B.n125 585
R823 B.n1047 B.n125 585
R824 B.n1016 B.n1015 585
R825 B.n1015 B.n124 585
R826 B.n1014 B.n120 585
R827 B.n1053 B.n120 585
R828 B.n1013 B.n119 585
R829 B.n1054 B.n119 585
R830 B.n1012 B.n118 585
R831 B.n1055 B.n118 585
R832 B.n1011 B.n1010 585
R833 B.n1010 B.n114 585
R834 B.n1009 B.n113 585
R835 B.n1061 B.n113 585
R836 B.n1008 B.n112 585
R837 B.n1062 B.n112 585
R838 B.n1007 B.n111 585
R839 B.n1063 B.n111 585
R840 B.n1006 B.n1005 585
R841 B.n1005 B.n107 585
R842 B.n1004 B.n106 585
R843 B.n1069 B.n106 585
R844 B.n1003 B.n105 585
R845 B.n1070 B.n105 585
R846 B.n1002 B.n104 585
R847 B.n1071 B.n104 585
R848 B.n1001 B.n1000 585
R849 B.n1000 B.n100 585
R850 B.n999 B.n99 585
R851 B.n1077 B.n99 585
R852 B.n998 B.n98 585
R853 B.n1078 B.n98 585
R854 B.n997 B.n97 585
R855 B.n1079 B.n97 585
R856 B.n996 B.n995 585
R857 B.n995 B.n93 585
R858 B.n994 B.n92 585
R859 B.n1085 B.n92 585
R860 B.n993 B.n91 585
R861 B.n1086 B.n91 585
R862 B.n992 B.n90 585
R863 B.n1087 B.n90 585
R864 B.n991 B.n990 585
R865 B.n990 B.n86 585
R866 B.n989 B.n85 585
R867 B.n1093 B.n85 585
R868 B.n988 B.n84 585
R869 B.n1094 B.n84 585
R870 B.n987 B.n83 585
R871 B.n1095 B.n83 585
R872 B.n986 B.n985 585
R873 B.n985 B.n79 585
R874 B.n984 B.n78 585
R875 B.n1101 B.n78 585
R876 B.n983 B.n77 585
R877 B.n1102 B.n77 585
R878 B.n982 B.n76 585
R879 B.n1103 B.n76 585
R880 B.n981 B.n980 585
R881 B.n980 B.n72 585
R882 B.n979 B.n71 585
R883 B.n1109 B.n71 585
R884 B.n978 B.n70 585
R885 B.n1110 B.n70 585
R886 B.n977 B.n69 585
R887 B.n1111 B.n69 585
R888 B.n976 B.n975 585
R889 B.n975 B.n65 585
R890 B.n974 B.n64 585
R891 B.n1117 B.n64 585
R892 B.n973 B.n63 585
R893 B.n1118 B.n63 585
R894 B.n972 B.n62 585
R895 B.n1119 B.n62 585
R896 B.n971 B.n970 585
R897 B.n970 B.n58 585
R898 B.n969 B.n57 585
R899 B.n1125 B.n57 585
R900 B.n968 B.n56 585
R901 B.n1126 B.n56 585
R902 B.n967 B.n55 585
R903 B.n1127 B.n55 585
R904 B.n966 B.n965 585
R905 B.n965 B.n51 585
R906 B.n964 B.n50 585
R907 B.n1133 B.n50 585
R908 B.n963 B.n49 585
R909 B.n1134 B.n49 585
R910 B.n962 B.n48 585
R911 B.n1135 B.n48 585
R912 B.n961 B.n960 585
R913 B.n960 B.n44 585
R914 B.n959 B.n43 585
R915 B.n1141 B.n43 585
R916 B.n958 B.n42 585
R917 B.n1142 B.n42 585
R918 B.n957 B.n41 585
R919 B.n1143 B.n41 585
R920 B.n956 B.n955 585
R921 B.n955 B.n40 585
R922 B.n954 B.n36 585
R923 B.n1149 B.n36 585
R924 B.n953 B.n35 585
R925 B.n1150 B.n35 585
R926 B.n952 B.n34 585
R927 B.n1151 B.n34 585
R928 B.n951 B.n950 585
R929 B.n950 B.n30 585
R930 B.n949 B.n29 585
R931 B.n1157 B.n29 585
R932 B.n948 B.n28 585
R933 B.n1158 B.n28 585
R934 B.n947 B.n27 585
R935 B.n1159 B.n27 585
R936 B.n946 B.n945 585
R937 B.n945 B.n23 585
R938 B.n944 B.n22 585
R939 B.n1165 B.n22 585
R940 B.n943 B.n21 585
R941 B.n1166 B.n21 585
R942 B.n942 B.n20 585
R943 B.n1167 B.n20 585
R944 B.n941 B.n940 585
R945 B.n940 B.n19 585
R946 B.n939 B.n15 585
R947 B.n1173 B.n15 585
R948 B.n938 B.n14 585
R949 B.n1174 B.n14 585
R950 B.n937 B.n13 585
R951 B.n1175 B.n13 585
R952 B.n936 B.n935 585
R953 B.n935 B.n12 585
R954 B.n934 B.n933 585
R955 B.n934 B.n8 585
R956 B.n932 B.n7 585
R957 B.n1182 B.n7 585
R958 B.n931 B.n6 585
R959 B.n1183 B.n6 585
R960 B.n930 B.n5 585
R961 B.n1184 B.n5 585
R962 B.n929 B.n928 585
R963 B.n928 B.n4 585
R964 B.n927 B.n344 585
R965 B.n927 B.n926 585
R966 B.n917 B.n345 585
R967 B.n346 B.n345 585
R968 B.n919 B.n918 585
R969 B.n920 B.n919 585
R970 B.n916 B.n351 585
R971 B.n351 B.n350 585
R972 B.n915 B.n914 585
R973 B.n914 B.n913 585
R974 B.n353 B.n352 585
R975 B.n906 B.n353 585
R976 B.n905 B.n904 585
R977 B.n907 B.n905 585
R978 B.n903 B.n358 585
R979 B.n358 B.n357 585
R980 B.n902 B.n901 585
R981 B.n901 B.n900 585
R982 B.n360 B.n359 585
R983 B.n361 B.n360 585
R984 B.n893 B.n892 585
R985 B.n894 B.n893 585
R986 B.n891 B.n366 585
R987 B.n366 B.n365 585
R988 B.n890 B.n889 585
R989 B.n889 B.n888 585
R990 B.n368 B.n367 585
R991 B.n369 B.n368 585
R992 B.n881 B.n880 585
R993 B.n882 B.n881 585
R994 B.n879 B.n374 585
R995 B.n374 B.n373 585
R996 B.n878 B.n877 585
R997 B.n877 B.n876 585
R998 B.n376 B.n375 585
R999 B.n869 B.n376 585
R1000 B.n868 B.n867 585
R1001 B.n870 B.n868 585
R1002 B.n866 B.n381 585
R1003 B.n381 B.n380 585
R1004 B.n865 B.n864 585
R1005 B.n864 B.n863 585
R1006 B.n383 B.n382 585
R1007 B.n384 B.n383 585
R1008 B.n856 B.n855 585
R1009 B.n857 B.n856 585
R1010 B.n854 B.n389 585
R1011 B.n389 B.n388 585
R1012 B.n853 B.n852 585
R1013 B.n852 B.n851 585
R1014 B.n391 B.n390 585
R1015 B.n392 B.n391 585
R1016 B.n844 B.n843 585
R1017 B.n845 B.n844 585
R1018 B.n842 B.n397 585
R1019 B.n397 B.n396 585
R1020 B.n841 B.n840 585
R1021 B.n840 B.n839 585
R1022 B.n399 B.n398 585
R1023 B.n400 B.n399 585
R1024 B.n832 B.n831 585
R1025 B.n833 B.n832 585
R1026 B.n830 B.n405 585
R1027 B.n405 B.n404 585
R1028 B.n829 B.n828 585
R1029 B.n828 B.n827 585
R1030 B.n407 B.n406 585
R1031 B.n408 B.n407 585
R1032 B.n820 B.n819 585
R1033 B.n821 B.n820 585
R1034 B.n818 B.n413 585
R1035 B.n413 B.n412 585
R1036 B.n817 B.n816 585
R1037 B.n816 B.n815 585
R1038 B.n415 B.n414 585
R1039 B.n416 B.n415 585
R1040 B.n808 B.n807 585
R1041 B.n809 B.n808 585
R1042 B.n806 B.n420 585
R1043 B.n424 B.n420 585
R1044 B.n805 B.n804 585
R1045 B.n804 B.n803 585
R1046 B.n422 B.n421 585
R1047 B.n423 B.n422 585
R1048 B.n796 B.n795 585
R1049 B.n797 B.n796 585
R1050 B.n794 B.n429 585
R1051 B.n429 B.n428 585
R1052 B.n793 B.n792 585
R1053 B.n792 B.n791 585
R1054 B.n431 B.n430 585
R1055 B.n432 B.n431 585
R1056 B.n784 B.n783 585
R1057 B.n785 B.n784 585
R1058 B.n782 B.n437 585
R1059 B.n437 B.n436 585
R1060 B.n781 B.n780 585
R1061 B.n780 B.n779 585
R1062 B.n439 B.n438 585
R1063 B.n440 B.n439 585
R1064 B.n772 B.n771 585
R1065 B.n773 B.n772 585
R1066 B.n770 B.n444 585
R1067 B.n448 B.n444 585
R1068 B.n769 B.n768 585
R1069 B.n768 B.n767 585
R1070 B.n446 B.n445 585
R1071 B.n447 B.n446 585
R1072 B.n760 B.n759 585
R1073 B.n761 B.n760 585
R1074 B.n758 B.n453 585
R1075 B.n453 B.n452 585
R1076 B.n757 B.n756 585
R1077 B.n756 B.n755 585
R1078 B.n455 B.n454 585
R1079 B.n456 B.n455 585
R1080 B.n748 B.n747 585
R1081 B.n749 B.n748 585
R1082 B.n746 B.n461 585
R1083 B.n461 B.n460 585
R1084 B.n745 B.n744 585
R1085 B.n744 B.n743 585
R1086 B.n463 B.n462 585
R1087 B.n464 B.n463 585
R1088 B.n736 B.n735 585
R1089 B.n737 B.n736 585
R1090 B.n734 B.n469 585
R1091 B.n469 B.n468 585
R1092 B.n733 B.n732 585
R1093 B.n732 B.n731 585
R1094 B.n471 B.n470 585
R1095 B.n724 B.n471 585
R1096 B.n723 B.n722 585
R1097 B.n725 B.n723 585
R1098 B.n721 B.n476 585
R1099 B.n476 B.n475 585
R1100 B.n720 B.n719 585
R1101 B.n719 B.n718 585
R1102 B.n478 B.n477 585
R1103 B.n479 B.n478 585
R1104 B.n711 B.n710 585
R1105 B.n712 B.n711 585
R1106 B.n709 B.n484 585
R1107 B.n484 B.n483 585
R1108 B.n708 B.n707 585
R1109 B.n707 B.n706 585
R1110 B.n486 B.n485 585
R1111 B.n487 B.n486 585
R1112 B.n699 B.n698 585
R1113 B.n700 B.n699 585
R1114 B.n490 B.n489 585
R1115 B.n538 B.n536 585
R1116 B.n539 B.n535 585
R1117 B.n539 B.n491 585
R1118 B.n542 B.n541 585
R1119 B.n543 B.n534 585
R1120 B.n545 B.n544 585
R1121 B.n547 B.n533 585
R1122 B.n550 B.n549 585
R1123 B.n551 B.n532 585
R1124 B.n553 B.n552 585
R1125 B.n555 B.n531 585
R1126 B.n558 B.n557 585
R1127 B.n559 B.n530 585
R1128 B.n561 B.n560 585
R1129 B.n563 B.n529 585
R1130 B.n566 B.n565 585
R1131 B.n567 B.n528 585
R1132 B.n569 B.n568 585
R1133 B.n571 B.n527 585
R1134 B.n574 B.n573 585
R1135 B.n575 B.n526 585
R1136 B.n577 B.n576 585
R1137 B.n579 B.n525 585
R1138 B.n582 B.n581 585
R1139 B.n583 B.n524 585
R1140 B.n585 B.n584 585
R1141 B.n587 B.n523 585
R1142 B.n590 B.n589 585
R1143 B.n591 B.n522 585
R1144 B.n593 B.n592 585
R1145 B.n595 B.n521 585
R1146 B.n598 B.n597 585
R1147 B.n599 B.n520 585
R1148 B.n601 B.n600 585
R1149 B.n603 B.n519 585
R1150 B.n606 B.n605 585
R1151 B.n608 B.n516 585
R1152 B.n610 B.n609 585
R1153 B.n612 B.n515 585
R1154 B.n615 B.n614 585
R1155 B.n616 B.n514 585
R1156 B.n618 B.n617 585
R1157 B.n620 B.n513 585
R1158 B.n623 B.n622 585
R1159 B.n624 B.n510 585
R1160 B.n627 B.n626 585
R1161 B.n629 B.n509 585
R1162 B.n632 B.n631 585
R1163 B.n633 B.n508 585
R1164 B.n635 B.n634 585
R1165 B.n637 B.n507 585
R1166 B.n640 B.n639 585
R1167 B.n641 B.n506 585
R1168 B.n643 B.n642 585
R1169 B.n645 B.n505 585
R1170 B.n648 B.n647 585
R1171 B.n649 B.n504 585
R1172 B.n651 B.n650 585
R1173 B.n653 B.n503 585
R1174 B.n656 B.n655 585
R1175 B.n657 B.n502 585
R1176 B.n659 B.n658 585
R1177 B.n661 B.n501 585
R1178 B.n664 B.n663 585
R1179 B.n665 B.n500 585
R1180 B.n667 B.n666 585
R1181 B.n669 B.n499 585
R1182 B.n672 B.n671 585
R1183 B.n673 B.n498 585
R1184 B.n675 B.n674 585
R1185 B.n677 B.n497 585
R1186 B.n680 B.n679 585
R1187 B.n681 B.n496 585
R1188 B.n683 B.n682 585
R1189 B.n685 B.n495 585
R1190 B.n688 B.n687 585
R1191 B.n689 B.n494 585
R1192 B.n691 B.n690 585
R1193 B.n693 B.n493 585
R1194 B.n696 B.n695 585
R1195 B.n697 B.n492 585
R1196 B.n702 B.n701 585
R1197 B.n701 B.n700 585
R1198 B.n703 B.n488 585
R1199 B.n488 B.n487 585
R1200 B.n705 B.n704 585
R1201 B.n706 B.n705 585
R1202 B.n482 B.n481 585
R1203 B.n483 B.n482 585
R1204 B.n714 B.n713 585
R1205 B.n713 B.n712 585
R1206 B.n715 B.n480 585
R1207 B.n480 B.n479 585
R1208 B.n717 B.n716 585
R1209 B.n718 B.n717 585
R1210 B.n474 B.n473 585
R1211 B.n475 B.n474 585
R1212 B.n727 B.n726 585
R1213 B.n726 B.n725 585
R1214 B.n728 B.n472 585
R1215 B.n724 B.n472 585
R1216 B.n730 B.n729 585
R1217 B.n731 B.n730 585
R1218 B.n467 B.n466 585
R1219 B.n468 B.n467 585
R1220 B.n739 B.n738 585
R1221 B.n738 B.n737 585
R1222 B.n740 B.n465 585
R1223 B.n465 B.n464 585
R1224 B.n742 B.n741 585
R1225 B.n743 B.n742 585
R1226 B.n459 B.n458 585
R1227 B.n460 B.n459 585
R1228 B.n751 B.n750 585
R1229 B.n750 B.n749 585
R1230 B.n752 B.n457 585
R1231 B.n457 B.n456 585
R1232 B.n754 B.n753 585
R1233 B.n755 B.n754 585
R1234 B.n451 B.n450 585
R1235 B.n452 B.n451 585
R1236 B.n763 B.n762 585
R1237 B.n762 B.n761 585
R1238 B.n764 B.n449 585
R1239 B.n449 B.n447 585
R1240 B.n766 B.n765 585
R1241 B.n767 B.n766 585
R1242 B.n443 B.n442 585
R1243 B.n448 B.n443 585
R1244 B.n775 B.n774 585
R1245 B.n774 B.n773 585
R1246 B.n776 B.n441 585
R1247 B.n441 B.n440 585
R1248 B.n778 B.n777 585
R1249 B.n779 B.n778 585
R1250 B.n435 B.n434 585
R1251 B.n436 B.n435 585
R1252 B.n787 B.n786 585
R1253 B.n786 B.n785 585
R1254 B.n788 B.n433 585
R1255 B.n433 B.n432 585
R1256 B.n790 B.n789 585
R1257 B.n791 B.n790 585
R1258 B.n427 B.n426 585
R1259 B.n428 B.n427 585
R1260 B.n799 B.n798 585
R1261 B.n798 B.n797 585
R1262 B.n800 B.n425 585
R1263 B.n425 B.n423 585
R1264 B.n802 B.n801 585
R1265 B.n803 B.n802 585
R1266 B.n419 B.n418 585
R1267 B.n424 B.n419 585
R1268 B.n811 B.n810 585
R1269 B.n810 B.n809 585
R1270 B.n812 B.n417 585
R1271 B.n417 B.n416 585
R1272 B.n814 B.n813 585
R1273 B.n815 B.n814 585
R1274 B.n411 B.n410 585
R1275 B.n412 B.n411 585
R1276 B.n823 B.n822 585
R1277 B.n822 B.n821 585
R1278 B.n824 B.n409 585
R1279 B.n409 B.n408 585
R1280 B.n826 B.n825 585
R1281 B.n827 B.n826 585
R1282 B.n403 B.n402 585
R1283 B.n404 B.n403 585
R1284 B.n835 B.n834 585
R1285 B.n834 B.n833 585
R1286 B.n836 B.n401 585
R1287 B.n401 B.n400 585
R1288 B.n838 B.n837 585
R1289 B.n839 B.n838 585
R1290 B.n395 B.n394 585
R1291 B.n396 B.n395 585
R1292 B.n847 B.n846 585
R1293 B.n846 B.n845 585
R1294 B.n848 B.n393 585
R1295 B.n393 B.n392 585
R1296 B.n850 B.n849 585
R1297 B.n851 B.n850 585
R1298 B.n387 B.n386 585
R1299 B.n388 B.n387 585
R1300 B.n859 B.n858 585
R1301 B.n858 B.n857 585
R1302 B.n860 B.n385 585
R1303 B.n385 B.n384 585
R1304 B.n862 B.n861 585
R1305 B.n863 B.n862 585
R1306 B.n379 B.n378 585
R1307 B.n380 B.n379 585
R1308 B.n872 B.n871 585
R1309 B.n871 B.n870 585
R1310 B.n873 B.n377 585
R1311 B.n869 B.n377 585
R1312 B.n875 B.n874 585
R1313 B.n876 B.n875 585
R1314 B.n372 B.n371 585
R1315 B.n373 B.n372 585
R1316 B.n884 B.n883 585
R1317 B.n883 B.n882 585
R1318 B.n885 B.n370 585
R1319 B.n370 B.n369 585
R1320 B.n887 B.n886 585
R1321 B.n888 B.n887 585
R1322 B.n364 B.n363 585
R1323 B.n365 B.n364 585
R1324 B.n896 B.n895 585
R1325 B.n895 B.n894 585
R1326 B.n897 B.n362 585
R1327 B.n362 B.n361 585
R1328 B.n899 B.n898 585
R1329 B.n900 B.n899 585
R1330 B.n356 B.n355 585
R1331 B.n357 B.n356 585
R1332 B.n909 B.n908 585
R1333 B.n908 B.n907 585
R1334 B.n910 B.n354 585
R1335 B.n906 B.n354 585
R1336 B.n912 B.n911 585
R1337 B.n913 B.n912 585
R1338 B.n349 B.n348 585
R1339 B.n350 B.n349 585
R1340 B.n922 B.n921 585
R1341 B.n921 B.n920 585
R1342 B.n923 B.n347 585
R1343 B.n347 B.n346 585
R1344 B.n925 B.n924 585
R1345 B.n926 B.n925 585
R1346 B.n3 B.n0 585
R1347 B.n4 B.n3 585
R1348 B.n1181 B.n1 585
R1349 B.n1182 B.n1181 585
R1350 B.n1180 B.n1179 585
R1351 B.n1180 B.n8 585
R1352 B.n1178 B.n9 585
R1353 B.n12 B.n9 585
R1354 B.n1177 B.n1176 585
R1355 B.n1176 B.n1175 585
R1356 B.n11 B.n10 585
R1357 B.n1174 B.n11 585
R1358 B.n1172 B.n1171 585
R1359 B.n1173 B.n1172 585
R1360 B.n1170 B.n16 585
R1361 B.n19 B.n16 585
R1362 B.n1169 B.n1168 585
R1363 B.n1168 B.n1167 585
R1364 B.n18 B.n17 585
R1365 B.n1166 B.n18 585
R1366 B.n1164 B.n1163 585
R1367 B.n1165 B.n1164 585
R1368 B.n1162 B.n24 585
R1369 B.n24 B.n23 585
R1370 B.n1161 B.n1160 585
R1371 B.n1160 B.n1159 585
R1372 B.n26 B.n25 585
R1373 B.n1158 B.n26 585
R1374 B.n1156 B.n1155 585
R1375 B.n1157 B.n1156 585
R1376 B.n1154 B.n31 585
R1377 B.n31 B.n30 585
R1378 B.n1153 B.n1152 585
R1379 B.n1152 B.n1151 585
R1380 B.n33 B.n32 585
R1381 B.n1150 B.n33 585
R1382 B.n1148 B.n1147 585
R1383 B.n1149 B.n1148 585
R1384 B.n1146 B.n37 585
R1385 B.n40 B.n37 585
R1386 B.n1145 B.n1144 585
R1387 B.n1144 B.n1143 585
R1388 B.n39 B.n38 585
R1389 B.n1142 B.n39 585
R1390 B.n1140 B.n1139 585
R1391 B.n1141 B.n1140 585
R1392 B.n1138 B.n45 585
R1393 B.n45 B.n44 585
R1394 B.n1137 B.n1136 585
R1395 B.n1136 B.n1135 585
R1396 B.n47 B.n46 585
R1397 B.n1134 B.n47 585
R1398 B.n1132 B.n1131 585
R1399 B.n1133 B.n1132 585
R1400 B.n1130 B.n52 585
R1401 B.n52 B.n51 585
R1402 B.n1129 B.n1128 585
R1403 B.n1128 B.n1127 585
R1404 B.n54 B.n53 585
R1405 B.n1126 B.n54 585
R1406 B.n1124 B.n1123 585
R1407 B.n1125 B.n1124 585
R1408 B.n1122 B.n59 585
R1409 B.n59 B.n58 585
R1410 B.n1121 B.n1120 585
R1411 B.n1120 B.n1119 585
R1412 B.n61 B.n60 585
R1413 B.n1118 B.n61 585
R1414 B.n1116 B.n1115 585
R1415 B.n1117 B.n1116 585
R1416 B.n1114 B.n66 585
R1417 B.n66 B.n65 585
R1418 B.n1113 B.n1112 585
R1419 B.n1112 B.n1111 585
R1420 B.n68 B.n67 585
R1421 B.n1110 B.n68 585
R1422 B.n1108 B.n1107 585
R1423 B.n1109 B.n1108 585
R1424 B.n1106 B.n73 585
R1425 B.n73 B.n72 585
R1426 B.n1105 B.n1104 585
R1427 B.n1104 B.n1103 585
R1428 B.n75 B.n74 585
R1429 B.n1102 B.n75 585
R1430 B.n1100 B.n1099 585
R1431 B.n1101 B.n1100 585
R1432 B.n1098 B.n80 585
R1433 B.n80 B.n79 585
R1434 B.n1097 B.n1096 585
R1435 B.n1096 B.n1095 585
R1436 B.n82 B.n81 585
R1437 B.n1094 B.n82 585
R1438 B.n1092 B.n1091 585
R1439 B.n1093 B.n1092 585
R1440 B.n1090 B.n87 585
R1441 B.n87 B.n86 585
R1442 B.n1089 B.n1088 585
R1443 B.n1088 B.n1087 585
R1444 B.n89 B.n88 585
R1445 B.n1086 B.n89 585
R1446 B.n1084 B.n1083 585
R1447 B.n1085 B.n1084 585
R1448 B.n1082 B.n94 585
R1449 B.n94 B.n93 585
R1450 B.n1081 B.n1080 585
R1451 B.n1080 B.n1079 585
R1452 B.n96 B.n95 585
R1453 B.n1078 B.n96 585
R1454 B.n1076 B.n1075 585
R1455 B.n1077 B.n1076 585
R1456 B.n1074 B.n101 585
R1457 B.n101 B.n100 585
R1458 B.n1073 B.n1072 585
R1459 B.n1072 B.n1071 585
R1460 B.n103 B.n102 585
R1461 B.n1070 B.n103 585
R1462 B.n1068 B.n1067 585
R1463 B.n1069 B.n1068 585
R1464 B.n1066 B.n108 585
R1465 B.n108 B.n107 585
R1466 B.n1065 B.n1064 585
R1467 B.n1064 B.n1063 585
R1468 B.n110 B.n109 585
R1469 B.n1062 B.n110 585
R1470 B.n1060 B.n1059 585
R1471 B.n1061 B.n1060 585
R1472 B.n1058 B.n115 585
R1473 B.n115 B.n114 585
R1474 B.n1057 B.n1056 585
R1475 B.n1056 B.n1055 585
R1476 B.n117 B.n116 585
R1477 B.n1054 B.n117 585
R1478 B.n1052 B.n1051 585
R1479 B.n1053 B.n1052 585
R1480 B.n1050 B.n121 585
R1481 B.n124 B.n121 585
R1482 B.n1049 B.n1048 585
R1483 B.n1048 B.n1047 585
R1484 B.n123 B.n122 585
R1485 B.n1046 B.n123 585
R1486 B.n1044 B.n1043 585
R1487 B.n1045 B.n1044 585
R1488 B.n1042 B.n129 585
R1489 B.n129 B.n128 585
R1490 B.n1041 B.n1040 585
R1491 B.n1040 B.n1039 585
R1492 B.n131 B.n130 585
R1493 B.n1038 B.n131 585
R1494 B.n1036 B.n1035 585
R1495 B.n1037 B.n1036 585
R1496 B.n1034 B.n136 585
R1497 B.n136 B.n135 585
R1498 B.n1033 B.n1032 585
R1499 B.n1032 B.n1031 585
R1500 B.n1185 B.n1184 585
R1501 B.n1183 B.n2 585
R1502 B.n1032 B.n138 497.305
R1503 B.n1029 B.n139 497.305
R1504 B.n699 B.n492 497.305
R1505 B.n701 B.n490 497.305
R1506 B.n181 B.t19 323.089
R1507 B.n511 B.t23 323.089
R1508 B.n183 B.t12 323.089
R1509 B.n517 B.t17 323.089
R1510 B.n183 B.t10 277.344
R1511 B.n181 B.t18 277.344
R1512 B.n511 B.t21 277.344
R1513 B.n517 B.t14 277.344
R1514 B.n1030 B.n179 256.663
R1515 B.n1030 B.n178 256.663
R1516 B.n1030 B.n177 256.663
R1517 B.n1030 B.n176 256.663
R1518 B.n1030 B.n175 256.663
R1519 B.n1030 B.n174 256.663
R1520 B.n1030 B.n173 256.663
R1521 B.n1030 B.n172 256.663
R1522 B.n1030 B.n171 256.663
R1523 B.n1030 B.n170 256.663
R1524 B.n1030 B.n169 256.663
R1525 B.n1030 B.n168 256.663
R1526 B.n1030 B.n167 256.663
R1527 B.n1030 B.n166 256.663
R1528 B.n1030 B.n165 256.663
R1529 B.n1030 B.n164 256.663
R1530 B.n1030 B.n163 256.663
R1531 B.n1030 B.n162 256.663
R1532 B.n1030 B.n161 256.663
R1533 B.n1030 B.n160 256.663
R1534 B.n1030 B.n159 256.663
R1535 B.n1030 B.n158 256.663
R1536 B.n1030 B.n157 256.663
R1537 B.n1030 B.n156 256.663
R1538 B.n1030 B.n155 256.663
R1539 B.n1030 B.n154 256.663
R1540 B.n1030 B.n153 256.663
R1541 B.n1030 B.n152 256.663
R1542 B.n1030 B.n151 256.663
R1543 B.n1030 B.n150 256.663
R1544 B.n1030 B.n149 256.663
R1545 B.n1030 B.n148 256.663
R1546 B.n1030 B.n147 256.663
R1547 B.n1030 B.n146 256.663
R1548 B.n1030 B.n145 256.663
R1549 B.n1030 B.n144 256.663
R1550 B.n1030 B.n143 256.663
R1551 B.n1030 B.n142 256.663
R1552 B.n1030 B.n141 256.663
R1553 B.n1030 B.n140 256.663
R1554 B.n537 B.n491 256.663
R1555 B.n540 B.n491 256.663
R1556 B.n546 B.n491 256.663
R1557 B.n548 B.n491 256.663
R1558 B.n554 B.n491 256.663
R1559 B.n556 B.n491 256.663
R1560 B.n562 B.n491 256.663
R1561 B.n564 B.n491 256.663
R1562 B.n570 B.n491 256.663
R1563 B.n572 B.n491 256.663
R1564 B.n578 B.n491 256.663
R1565 B.n580 B.n491 256.663
R1566 B.n586 B.n491 256.663
R1567 B.n588 B.n491 256.663
R1568 B.n594 B.n491 256.663
R1569 B.n596 B.n491 256.663
R1570 B.n602 B.n491 256.663
R1571 B.n604 B.n491 256.663
R1572 B.n611 B.n491 256.663
R1573 B.n613 B.n491 256.663
R1574 B.n619 B.n491 256.663
R1575 B.n621 B.n491 256.663
R1576 B.n628 B.n491 256.663
R1577 B.n630 B.n491 256.663
R1578 B.n636 B.n491 256.663
R1579 B.n638 B.n491 256.663
R1580 B.n644 B.n491 256.663
R1581 B.n646 B.n491 256.663
R1582 B.n652 B.n491 256.663
R1583 B.n654 B.n491 256.663
R1584 B.n660 B.n491 256.663
R1585 B.n662 B.n491 256.663
R1586 B.n668 B.n491 256.663
R1587 B.n670 B.n491 256.663
R1588 B.n676 B.n491 256.663
R1589 B.n678 B.n491 256.663
R1590 B.n684 B.n491 256.663
R1591 B.n686 B.n491 256.663
R1592 B.n692 B.n491 256.663
R1593 B.n694 B.n491 256.663
R1594 B.n1187 B.n1186 256.663
R1595 B.n182 B.t20 248.036
R1596 B.n512 B.t22 248.036
R1597 B.n184 B.t13 248.036
R1598 B.n518 B.t16 248.036
R1599 B.n188 B.n187 163.367
R1600 B.n192 B.n191 163.367
R1601 B.n196 B.n195 163.367
R1602 B.n200 B.n199 163.367
R1603 B.n204 B.n203 163.367
R1604 B.n208 B.n207 163.367
R1605 B.n212 B.n211 163.367
R1606 B.n216 B.n215 163.367
R1607 B.n220 B.n219 163.367
R1608 B.n224 B.n223 163.367
R1609 B.n228 B.n227 163.367
R1610 B.n232 B.n231 163.367
R1611 B.n236 B.n235 163.367
R1612 B.n240 B.n239 163.367
R1613 B.n244 B.n243 163.367
R1614 B.n248 B.n247 163.367
R1615 B.n252 B.n251 163.367
R1616 B.n256 B.n255 163.367
R1617 B.n260 B.n259 163.367
R1618 B.n264 B.n263 163.367
R1619 B.n268 B.n267 163.367
R1620 B.n272 B.n271 163.367
R1621 B.n277 B.n276 163.367
R1622 B.n281 B.n280 163.367
R1623 B.n285 B.n284 163.367
R1624 B.n289 B.n288 163.367
R1625 B.n293 B.n292 163.367
R1626 B.n297 B.n296 163.367
R1627 B.n301 B.n300 163.367
R1628 B.n305 B.n304 163.367
R1629 B.n309 B.n308 163.367
R1630 B.n313 B.n312 163.367
R1631 B.n317 B.n316 163.367
R1632 B.n321 B.n320 163.367
R1633 B.n325 B.n324 163.367
R1634 B.n329 B.n328 163.367
R1635 B.n333 B.n332 163.367
R1636 B.n337 B.n336 163.367
R1637 B.n341 B.n340 163.367
R1638 B.n1029 B.n180 163.367
R1639 B.n699 B.n486 163.367
R1640 B.n707 B.n486 163.367
R1641 B.n707 B.n484 163.367
R1642 B.n711 B.n484 163.367
R1643 B.n711 B.n478 163.367
R1644 B.n719 B.n478 163.367
R1645 B.n719 B.n476 163.367
R1646 B.n723 B.n476 163.367
R1647 B.n723 B.n471 163.367
R1648 B.n732 B.n471 163.367
R1649 B.n732 B.n469 163.367
R1650 B.n736 B.n469 163.367
R1651 B.n736 B.n463 163.367
R1652 B.n744 B.n463 163.367
R1653 B.n744 B.n461 163.367
R1654 B.n748 B.n461 163.367
R1655 B.n748 B.n455 163.367
R1656 B.n756 B.n455 163.367
R1657 B.n756 B.n453 163.367
R1658 B.n760 B.n453 163.367
R1659 B.n760 B.n446 163.367
R1660 B.n768 B.n446 163.367
R1661 B.n768 B.n444 163.367
R1662 B.n772 B.n444 163.367
R1663 B.n772 B.n439 163.367
R1664 B.n780 B.n439 163.367
R1665 B.n780 B.n437 163.367
R1666 B.n784 B.n437 163.367
R1667 B.n784 B.n431 163.367
R1668 B.n792 B.n431 163.367
R1669 B.n792 B.n429 163.367
R1670 B.n796 B.n429 163.367
R1671 B.n796 B.n422 163.367
R1672 B.n804 B.n422 163.367
R1673 B.n804 B.n420 163.367
R1674 B.n808 B.n420 163.367
R1675 B.n808 B.n415 163.367
R1676 B.n816 B.n415 163.367
R1677 B.n816 B.n413 163.367
R1678 B.n820 B.n413 163.367
R1679 B.n820 B.n407 163.367
R1680 B.n828 B.n407 163.367
R1681 B.n828 B.n405 163.367
R1682 B.n832 B.n405 163.367
R1683 B.n832 B.n399 163.367
R1684 B.n840 B.n399 163.367
R1685 B.n840 B.n397 163.367
R1686 B.n844 B.n397 163.367
R1687 B.n844 B.n391 163.367
R1688 B.n852 B.n391 163.367
R1689 B.n852 B.n389 163.367
R1690 B.n856 B.n389 163.367
R1691 B.n856 B.n383 163.367
R1692 B.n864 B.n383 163.367
R1693 B.n864 B.n381 163.367
R1694 B.n868 B.n381 163.367
R1695 B.n868 B.n376 163.367
R1696 B.n877 B.n376 163.367
R1697 B.n877 B.n374 163.367
R1698 B.n881 B.n374 163.367
R1699 B.n881 B.n368 163.367
R1700 B.n889 B.n368 163.367
R1701 B.n889 B.n366 163.367
R1702 B.n893 B.n366 163.367
R1703 B.n893 B.n360 163.367
R1704 B.n901 B.n360 163.367
R1705 B.n901 B.n358 163.367
R1706 B.n905 B.n358 163.367
R1707 B.n905 B.n353 163.367
R1708 B.n914 B.n353 163.367
R1709 B.n914 B.n351 163.367
R1710 B.n919 B.n351 163.367
R1711 B.n919 B.n345 163.367
R1712 B.n927 B.n345 163.367
R1713 B.n928 B.n927 163.367
R1714 B.n928 B.n5 163.367
R1715 B.n6 B.n5 163.367
R1716 B.n7 B.n6 163.367
R1717 B.n934 B.n7 163.367
R1718 B.n935 B.n934 163.367
R1719 B.n935 B.n13 163.367
R1720 B.n14 B.n13 163.367
R1721 B.n15 B.n14 163.367
R1722 B.n940 B.n15 163.367
R1723 B.n940 B.n20 163.367
R1724 B.n21 B.n20 163.367
R1725 B.n22 B.n21 163.367
R1726 B.n945 B.n22 163.367
R1727 B.n945 B.n27 163.367
R1728 B.n28 B.n27 163.367
R1729 B.n29 B.n28 163.367
R1730 B.n950 B.n29 163.367
R1731 B.n950 B.n34 163.367
R1732 B.n35 B.n34 163.367
R1733 B.n36 B.n35 163.367
R1734 B.n955 B.n36 163.367
R1735 B.n955 B.n41 163.367
R1736 B.n42 B.n41 163.367
R1737 B.n43 B.n42 163.367
R1738 B.n960 B.n43 163.367
R1739 B.n960 B.n48 163.367
R1740 B.n49 B.n48 163.367
R1741 B.n50 B.n49 163.367
R1742 B.n965 B.n50 163.367
R1743 B.n965 B.n55 163.367
R1744 B.n56 B.n55 163.367
R1745 B.n57 B.n56 163.367
R1746 B.n970 B.n57 163.367
R1747 B.n970 B.n62 163.367
R1748 B.n63 B.n62 163.367
R1749 B.n64 B.n63 163.367
R1750 B.n975 B.n64 163.367
R1751 B.n975 B.n69 163.367
R1752 B.n70 B.n69 163.367
R1753 B.n71 B.n70 163.367
R1754 B.n980 B.n71 163.367
R1755 B.n980 B.n76 163.367
R1756 B.n77 B.n76 163.367
R1757 B.n78 B.n77 163.367
R1758 B.n985 B.n78 163.367
R1759 B.n985 B.n83 163.367
R1760 B.n84 B.n83 163.367
R1761 B.n85 B.n84 163.367
R1762 B.n990 B.n85 163.367
R1763 B.n990 B.n90 163.367
R1764 B.n91 B.n90 163.367
R1765 B.n92 B.n91 163.367
R1766 B.n995 B.n92 163.367
R1767 B.n995 B.n97 163.367
R1768 B.n98 B.n97 163.367
R1769 B.n99 B.n98 163.367
R1770 B.n1000 B.n99 163.367
R1771 B.n1000 B.n104 163.367
R1772 B.n105 B.n104 163.367
R1773 B.n106 B.n105 163.367
R1774 B.n1005 B.n106 163.367
R1775 B.n1005 B.n111 163.367
R1776 B.n112 B.n111 163.367
R1777 B.n113 B.n112 163.367
R1778 B.n1010 B.n113 163.367
R1779 B.n1010 B.n118 163.367
R1780 B.n119 B.n118 163.367
R1781 B.n120 B.n119 163.367
R1782 B.n1015 B.n120 163.367
R1783 B.n1015 B.n125 163.367
R1784 B.n126 B.n125 163.367
R1785 B.n127 B.n126 163.367
R1786 B.n1020 B.n127 163.367
R1787 B.n1020 B.n132 163.367
R1788 B.n133 B.n132 163.367
R1789 B.n134 B.n133 163.367
R1790 B.n1025 B.n134 163.367
R1791 B.n1025 B.n139 163.367
R1792 B.n539 B.n538 163.367
R1793 B.n541 B.n539 163.367
R1794 B.n545 B.n534 163.367
R1795 B.n549 B.n547 163.367
R1796 B.n553 B.n532 163.367
R1797 B.n557 B.n555 163.367
R1798 B.n561 B.n530 163.367
R1799 B.n565 B.n563 163.367
R1800 B.n569 B.n528 163.367
R1801 B.n573 B.n571 163.367
R1802 B.n577 B.n526 163.367
R1803 B.n581 B.n579 163.367
R1804 B.n585 B.n524 163.367
R1805 B.n589 B.n587 163.367
R1806 B.n593 B.n522 163.367
R1807 B.n597 B.n595 163.367
R1808 B.n601 B.n520 163.367
R1809 B.n605 B.n603 163.367
R1810 B.n610 B.n516 163.367
R1811 B.n614 B.n612 163.367
R1812 B.n618 B.n514 163.367
R1813 B.n622 B.n620 163.367
R1814 B.n627 B.n510 163.367
R1815 B.n631 B.n629 163.367
R1816 B.n635 B.n508 163.367
R1817 B.n639 B.n637 163.367
R1818 B.n643 B.n506 163.367
R1819 B.n647 B.n645 163.367
R1820 B.n651 B.n504 163.367
R1821 B.n655 B.n653 163.367
R1822 B.n659 B.n502 163.367
R1823 B.n663 B.n661 163.367
R1824 B.n667 B.n500 163.367
R1825 B.n671 B.n669 163.367
R1826 B.n675 B.n498 163.367
R1827 B.n679 B.n677 163.367
R1828 B.n683 B.n496 163.367
R1829 B.n687 B.n685 163.367
R1830 B.n691 B.n494 163.367
R1831 B.n695 B.n693 163.367
R1832 B.n701 B.n488 163.367
R1833 B.n705 B.n488 163.367
R1834 B.n705 B.n482 163.367
R1835 B.n713 B.n482 163.367
R1836 B.n713 B.n480 163.367
R1837 B.n717 B.n480 163.367
R1838 B.n717 B.n474 163.367
R1839 B.n726 B.n474 163.367
R1840 B.n726 B.n472 163.367
R1841 B.n730 B.n472 163.367
R1842 B.n730 B.n467 163.367
R1843 B.n738 B.n467 163.367
R1844 B.n738 B.n465 163.367
R1845 B.n742 B.n465 163.367
R1846 B.n742 B.n459 163.367
R1847 B.n750 B.n459 163.367
R1848 B.n750 B.n457 163.367
R1849 B.n754 B.n457 163.367
R1850 B.n754 B.n451 163.367
R1851 B.n762 B.n451 163.367
R1852 B.n762 B.n449 163.367
R1853 B.n766 B.n449 163.367
R1854 B.n766 B.n443 163.367
R1855 B.n774 B.n443 163.367
R1856 B.n774 B.n441 163.367
R1857 B.n778 B.n441 163.367
R1858 B.n778 B.n435 163.367
R1859 B.n786 B.n435 163.367
R1860 B.n786 B.n433 163.367
R1861 B.n790 B.n433 163.367
R1862 B.n790 B.n427 163.367
R1863 B.n798 B.n427 163.367
R1864 B.n798 B.n425 163.367
R1865 B.n802 B.n425 163.367
R1866 B.n802 B.n419 163.367
R1867 B.n810 B.n419 163.367
R1868 B.n810 B.n417 163.367
R1869 B.n814 B.n417 163.367
R1870 B.n814 B.n411 163.367
R1871 B.n822 B.n411 163.367
R1872 B.n822 B.n409 163.367
R1873 B.n826 B.n409 163.367
R1874 B.n826 B.n403 163.367
R1875 B.n834 B.n403 163.367
R1876 B.n834 B.n401 163.367
R1877 B.n838 B.n401 163.367
R1878 B.n838 B.n395 163.367
R1879 B.n846 B.n395 163.367
R1880 B.n846 B.n393 163.367
R1881 B.n850 B.n393 163.367
R1882 B.n850 B.n387 163.367
R1883 B.n858 B.n387 163.367
R1884 B.n858 B.n385 163.367
R1885 B.n862 B.n385 163.367
R1886 B.n862 B.n379 163.367
R1887 B.n871 B.n379 163.367
R1888 B.n871 B.n377 163.367
R1889 B.n875 B.n377 163.367
R1890 B.n875 B.n372 163.367
R1891 B.n883 B.n372 163.367
R1892 B.n883 B.n370 163.367
R1893 B.n887 B.n370 163.367
R1894 B.n887 B.n364 163.367
R1895 B.n895 B.n364 163.367
R1896 B.n895 B.n362 163.367
R1897 B.n899 B.n362 163.367
R1898 B.n899 B.n356 163.367
R1899 B.n908 B.n356 163.367
R1900 B.n908 B.n354 163.367
R1901 B.n912 B.n354 163.367
R1902 B.n912 B.n349 163.367
R1903 B.n921 B.n349 163.367
R1904 B.n921 B.n347 163.367
R1905 B.n925 B.n347 163.367
R1906 B.n925 B.n3 163.367
R1907 B.n1185 B.n3 163.367
R1908 B.n1181 B.n2 163.367
R1909 B.n1181 B.n1180 163.367
R1910 B.n1180 B.n9 163.367
R1911 B.n1176 B.n9 163.367
R1912 B.n1176 B.n11 163.367
R1913 B.n1172 B.n11 163.367
R1914 B.n1172 B.n16 163.367
R1915 B.n1168 B.n16 163.367
R1916 B.n1168 B.n18 163.367
R1917 B.n1164 B.n18 163.367
R1918 B.n1164 B.n24 163.367
R1919 B.n1160 B.n24 163.367
R1920 B.n1160 B.n26 163.367
R1921 B.n1156 B.n26 163.367
R1922 B.n1156 B.n31 163.367
R1923 B.n1152 B.n31 163.367
R1924 B.n1152 B.n33 163.367
R1925 B.n1148 B.n33 163.367
R1926 B.n1148 B.n37 163.367
R1927 B.n1144 B.n37 163.367
R1928 B.n1144 B.n39 163.367
R1929 B.n1140 B.n39 163.367
R1930 B.n1140 B.n45 163.367
R1931 B.n1136 B.n45 163.367
R1932 B.n1136 B.n47 163.367
R1933 B.n1132 B.n47 163.367
R1934 B.n1132 B.n52 163.367
R1935 B.n1128 B.n52 163.367
R1936 B.n1128 B.n54 163.367
R1937 B.n1124 B.n54 163.367
R1938 B.n1124 B.n59 163.367
R1939 B.n1120 B.n59 163.367
R1940 B.n1120 B.n61 163.367
R1941 B.n1116 B.n61 163.367
R1942 B.n1116 B.n66 163.367
R1943 B.n1112 B.n66 163.367
R1944 B.n1112 B.n68 163.367
R1945 B.n1108 B.n68 163.367
R1946 B.n1108 B.n73 163.367
R1947 B.n1104 B.n73 163.367
R1948 B.n1104 B.n75 163.367
R1949 B.n1100 B.n75 163.367
R1950 B.n1100 B.n80 163.367
R1951 B.n1096 B.n80 163.367
R1952 B.n1096 B.n82 163.367
R1953 B.n1092 B.n82 163.367
R1954 B.n1092 B.n87 163.367
R1955 B.n1088 B.n87 163.367
R1956 B.n1088 B.n89 163.367
R1957 B.n1084 B.n89 163.367
R1958 B.n1084 B.n94 163.367
R1959 B.n1080 B.n94 163.367
R1960 B.n1080 B.n96 163.367
R1961 B.n1076 B.n96 163.367
R1962 B.n1076 B.n101 163.367
R1963 B.n1072 B.n101 163.367
R1964 B.n1072 B.n103 163.367
R1965 B.n1068 B.n103 163.367
R1966 B.n1068 B.n108 163.367
R1967 B.n1064 B.n108 163.367
R1968 B.n1064 B.n110 163.367
R1969 B.n1060 B.n110 163.367
R1970 B.n1060 B.n115 163.367
R1971 B.n1056 B.n115 163.367
R1972 B.n1056 B.n117 163.367
R1973 B.n1052 B.n117 163.367
R1974 B.n1052 B.n121 163.367
R1975 B.n1048 B.n121 163.367
R1976 B.n1048 B.n123 163.367
R1977 B.n1044 B.n123 163.367
R1978 B.n1044 B.n129 163.367
R1979 B.n1040 B.n129 163.367
R1980 B.n1040 B.n131 163.367
R1981 B.n1036 B.n131 163.367
R1982 B.n1036 B.n136 163.367
R1983 B.n1032 B.n136 163.367
R1984 B.n700 B.n491 84.1456
R1985 B.n1031 B.n1030 84.1456
R1986 B.n184 B.n183 75.0551
R1987 B.n182 B.n181 75.0551
R1988 B.n512 B.n511 75.0551
R1989 B.n518 B.n517 75.0551
R1990 B.n140 B.n138 71.676
R1991 B.n188 B.n141 71.676
R1992 B.n192 B.n142 71.676
R1993 B.n196 B.n143 71.676
R1994 B.n200 B.n144 71.676
R1995 B.n204 B.n145 71.676
R1996 B.n208 B.n146 71.676
R1997 B.n212 B.n147 71.676
R1998 B.n216 B.n148 71.676
R1999 B.n220 B.n149 71.676
R2000 B.n224 B.n150 71.676
R2001 B.n228 B.n151 71.676
R2002 B.n232 B.n152 71.676
R2003 B.n236 B.n153 71.676
R2004 B.n240 B.n154 71.676
R2005 B.n244 B.n155 71.676
R2006 B.n248 B.n156 71.676
R2007 B.n252 B.n157 71.676
R2008 B.n256 B.n158 71.676
R2009 B.n260 B.n159 71.676
R2010 B.n264 B.n160 71.676
R2011 B.n268 B.n161 71.676
R2012 B.n272 B.n162 71.676
R2013 B.n277 B.n163 71.676
R2014 B.n281 B.n164 71.676
R2015 B.n285 B.n165 71.676
R2016 B.n289 B.n166 71.676
R2017 B.n293 B.n167 71.676
R2018 B.n297 B.n168 71.676
R2019 B.n301 B.n169 71.676
R2020 B.n305 B.n170 71.676
R2021 B.n309 B.n171 71.676
R2022 B.n313 B.n172 71.676
R2023 B.n317 B.n173 71.676
R2024 B.n321 B.n174 71.676
R2025 B.n325 B.n175 71.676
R2026 B.n329 B.n176 71.676
R2027 B.n333 B.n177 71.676
R2028 B.n337 B.n178 71.676
R2029 B.n341 B.n179 71.676
R2030 B.n180 B.n179 71.676
R2031 B.n340 B.n178 71.676
R2032 B.n336 B.n177 71.676
R2033 B.n332 B.n176 71.676
R2034 B.n328 B.n175 71.676
R2035 B.n324 B.n174 71.676
R2036 B.n320 B.n173 71.676
R2037 B.n316 B.n172 71.676
R2038 B.n312 B.n171 71.676
R2039 B.n308 B.n170 71.676
R2040 B.n304 B.n169 71.676
R2041 B.n300 B.n168 71.676
R2042 B.n296 B.n167 71.676
R2043 B.n292 B.n166 71.676
R2044 B.n288 B.n165 71.676
R2045 B.n284 B.n164 71.676
R2046 B.n280 B.n163 71.676
R2047 B.n276 B.n162 71.676
R2048 B.n271 B.n161 71.676
R2049 B.n267 B.n160 71.676
R2050 B.n263 B.n159 71.676
R2051 B.n259 B.n158 71.676
R2052 B.n255 B.n157 71.676
R2053 B.n251 B.n156 71.676
R2054 B.n247 B.n155 71.676
R2055 B.n243 B.n154 71.676
R2056 B.n239 B.n153 71.676
R2057 B.n235 B.n152 71.676
R2058 B.n231 B.n151 71.676
R2059 B.n227 B.n150 71.676
R2060 B.n223 B.n149 71.676
R2061 B.n219 B.n148 71.676
R2062 B.n215 B.n147 71.676
R2063 B.n211 B.n146 71.676
R2064 B.n207 B.n145 71.676
R2065 B.n203 B.n144 71.676
R2066 B.n199 B.n143 71.676
R2067 B.n195 B.n142 71.676
R2068 B.n191 B.n141 71.676
R2069 B.n187 B.n140 71.676
R2070 B.n537 B.n490 71.676
R2071 B.n541 B.n540 71.676
R2072 B.n546 B.n545 71.676
R2073 B.n549 B.n548 71.676
R2074 B.n554 B.n553 71.676
R2075 B.n557 B.n556 71.676
R2076 B.n562 B.n561 71.676
R2077 B.n565 B.n564 71.676
R2078 B.n570 B.n569 71.676
R2079 B.n573 B.n572 71.676
R2080 B.n578 B.n577 71.676
R2081 B.n581 B.n580 71.676
R2082 B.n586 B.n585 71.676
R2083 B.n589 B.n588 71.676
R2084 B.n594 B.n593 71.676
R2085 B.n597 B.n596 71.676
R2086 B.n602 B.n601 71.676
R2087 B.n605 B.n604 71.676
R2088 B.n611 B.n610 71.676
R2089 B.n614 B.n613 71.676
R2090 B.n619 B.n618 71.676
R2091 B.n622 B.n621 71.676
R2092 B.n628 B.n627 71.676
R2093 B.n631 B.n630 71.676
R2094 B.n636 B.n635 71.676
R2095 B.n639 B.n638 71.676
R2096 B.n644 B.n643 71.676
R2097 B.n647 B.n646 71.676
R2098 B.n652 B.n651 71.676
R2099 B.n655 B.n654 71.676
R2100 B.n660 B.n659 71.676
R2101 B.n663 B.n662 71.676
R2102 B.n668 B.n667 71.676
R2103 B.n671 B.n670 71.676
R2104 B.n676 B.n675 71.676
R2105 B.n679 B.n678 71.676
R2106 B.n684 B.n683 71.676
R2107 B.n687 B.n686 71.676
R2108 B.n692 B.n691 71.676
R2109 B.n695 B.n694 71.676
R2110 B.n538 B.n537 71.676
R2111 B.n540 B.n534 71.676
R2112 B.n547 B.n546 71.676
R2113 B.n548 B.n532 71.676
R2114 B.n555 B.n554 71.676
R2115 B.n556 B.n530 71.676
R2116 B.n563 B.n562 71.676
R2117 B.n564 B.n528 71.676
R2118 B.n571 B.n570 71.676
R2119 B.n572 B.n526 71.676
R2120 B.n579 B.n578 71.676
R2121 B.n580 B.n524 71.676
R2122 B.n587 B.n586 71.676
R2123 B.n588 B.n522 71.676
R2124 B.n595 B.n594 71.676
R2125 B.n596 B.n520 71.676
R2126 B.n603 B.n602 71.676
R2127 B.n604 B.n516 71.676
R2128 B.n612 B.n611 71.676
R2129 B.n613 B.n514 71.676
R2130 B.n620 B.n619 71.676
R2131 B.n621 B.n510 71.676
R2132 B.n629 B.n628 71.676
R2133 B.n630 B.n508 71.676
R2134 B.n637 B.n636 71.676
R2135 B.n638 B.n506 71.676
R2136 B.n645 B.n644 71.676
R2137 B.n646 B.n504 71.676
R2138 B.n653 B.n652 71.676
R2139 B.n654 B.n502 71.676
R2140 B.n661 B.n660 71.676
R2141 B.n662 B.n500 71.676
R2142 B.n669 B.n668 71.676
R2143 B.n670 B.n498 71.676
R2144 B.n677 B.n676 71.676
R2145 B.n678 B.n496 71.676
R2146 B.n685 B.n684 71.676
R2147 B.n686 B.n494 71.676
R2148 B.n693 B.n692 71.676
R2149 B.n694 B.n492 71.676
R2150 B.n1186 B.n1185 71.676
R2151 B.n1186 B.n2 71.676
R2152 B.n185 B.n184 59.5399
R2153 B.n274 B.n182 59.5399
R2154 B.n625 B.n512 59.5399
R2155 B.n607 B.n518 59.5399
R2156 B.n700 B.n487 48.9054
R2157 B.n706 B.n487 48.9054
R2158 B.n706 B.n483 48.9054
R2159 B.n712 B.n483 48.9054
R2160 B.n712 B.n479 48.9054
R2161 B.n718 B.n479 48.9054
R2162 B.n718 B.n475 48.9054
R2163 B.n725 B.n475 48.9054
R2164 B.n725 B.n724 48.9054
R2165 B.n731 B.n468 48.9054
R2166 B.n737 B.n468 48.9054
R2167 B.n737 B.n464 48.9054
R2168 B.n743 B.n464 48.9054
R2169 B.n743 B.n460 48.9054
R2170 B.n749 B.n460 48.9054
R2171 B.n749 B.n456 48.9054
R2172 B.n755 B.n456 48.9054
R2173 B.n755 B.n452 48.9054
R2174 B.n761 B.n452 48.9054
R2175 B.n761 B.n447 48.9054
R2176 B.n767 B.n447 48.9054
R2177 B.n767 B.n448 48.9054
R2178 B.n773 B.n440 48.9054
R2179 B.n779 B.n440 48.9054
R2180 B.n779 B.n436 48.9054
R2181 B.n785 B.n436 48.9054
R2182 B.n785 B.n432 48.9054
R2183 B.n791 B.n432 48.9054
R2184 B.n791 B.n428 48.9054
R2185 B.n797 B.n428 48.9054
R2186 B.n797 B.n423 48.9054
R2187 B.n803 B.n423 48.9054
R2188 B.n803 B.n424 48.9054
R2189 B.n809 B.n416 48.9054
R2190 B.n815 B.n416 48.9054
R2191 B.n815 B.n412 48.9054
R2192 B.n821 B.n412 48.9054
R2193 B.n821 B.n408 48.9054
R2194 B.n827 B.n408 48.9054
R2195 B.n827 B.n404 48.9054
R2196 B.n833 B.n404 48.9054
R2197 B.n833 B.n400 48.9054
R2198 B.n839 B.n400 48.9054
R2199 B.n845 B.n396 48.9054
R2200 B.n845 B.n392 48.9054
R2201 B.n851 B.n392 48.9054
R2202 B.n851 B.n388 48.9054
R2203 B.n857 B.n388 48.9054
R2204 B.n857 B.n384 48.9054
R2205 B.n863 B.n384 48.9054
R2206 B.n863 B.n380 48.9054
R2207 B.n870 B.n380 48.9054
R2208 B.n870 B.n869 48.9054
R2209 B.n876 B.n373 48.9054
R2210 B.n882 B.n373 48.9054
R2211 B.n882 B.n369 48.9054
R2212 B.n888 B.n369 48.9054
R2213 B.n888 B.n365 48.9054
R2214 B.n894 B.n365 48.9054
R2215 B.n894 B.n361 48.9054
R2216 B.n900 B.n361 48.9054
R2217 B.n900 B.n357 48.9054
R2218 B.n907 B.n357 48.9054
R2219 B.n907 B.n906 48.9054
R2220 B.n913 B.n350 48.9054
R2221 B.n920 B.n350 48.9054
R2222 B.n920 B.n346 48.9054
R2223 B.n926 B.n346 48.9054
R2224 B.n926 B.n4 48.9054
R2225 B.n1184 B.n4 48.9054
R2226 B.n1184 B.n1183 48.9054
R2227 B.n1183 B.n1182 48.9054
R2228 B.n1182 B.n8 48.9054
R2229 B.n12 B.n8 48.9054
R2230 B.n1175 B.n12 48.9054
R2231 B.n1175 B.n1174 48.9054
R2232 B.n1174 B.n1173 48.9054
R2233 B.n1167 B.n19 48.9054
R2234 B.n1167 B.n1166 48.9054
R2235 B.n1166 B.n1165 48.9054
R2236 B.n1165 B.n23 48.9054
R2237 B.n1159 B.n23 48.9054
R2238 B.n1159 B.n1158 48.9054
R2239 B.n1158 B.n1157 48.9054
R2240 B.n1157 B.n30 48.9054
R2241 B.n1151 B.n30 48.9054
R2242 B.n1151 B.n1150 48.9054
R2243 B.n1150 B.n1149 48.9054
R2244 B.n1143 B.n40 48.9054
R2245 B.n1143 B.n1142 48.9054
R2246 B.n1142 B.n1141 48.9054
R2247 B.n1141 B.n44 48.9054
R2248 B.n1135 B.n44 48.9054
R2249 B.n1135 B.n1134 48.9054
R2250 B.n1134 B.n1133 48.9054
R2251 B.n1133 B.n51 48.9054
R2252 B.n1127 B.n51 48.9054
R2253 B.n1127 B.n1126 48.9054
R2254 B.n1125 B.n58 48.9054
R2255 B.n1119 B.n58 48.9054
R2256 B.n1119 B.n1118 48.9054
R2257 B.n1118 B.n1117 48.9054
R2258 B.n1117 B.n65 48.9054
R2259 B.n1111 B.n65 48.9054
R2260 B.n1111 B.n1110 48.9054
R2261 B.n1110 B.n1109 48.9054
R2262 B.n1109 B.n72 48.9054
R2263 B.n1103 B.n72 48.9054
R2264 B.n1102 B.n1101 48.9054
R2265 B.n1101 B.n79 48.9054
R2266 B.n1095 B.n79 48.9054
R2267 B.n1095 B.n1094 48.9054
R2268 B.n1094 B.n1093 48.9054
R2269 B.n1093 B.n86 48.9054
R2270 B.n1087 B.n86 48.9054
R2271 B.n1087 B.n1086 48.9054
R2272 B.n1086 B.n1085 48.9054
R2273 B.n1085 B.n93 48.9054
R2274 B.n1079 B.n93 48.9054
R2275 B.n1078 B.n1077 48.9054
R2276 B.n1077 B.n100 48.9054
R2277 B.n1071 B.n100 48.9054
R2278 B.n1071 B.n1070 48.9054
R2279 B.n1070 B.n1069 48.9054
R2280 B.n1069 B.n107 48.9054
R2281 B.n1063 B.n107 48.9054
R2282 B.n1063 B.n1062 48.9054
R2283 B.n1062 B.n1061 48.9054
R2284 B.n1061 B.n114 48.9054
R2285 B.n1055 B.n114 48.9054
R2286 B.n1055 B.n1054 48.9054
R2287 B.n1054 B.n1053 48.9054
R2288 B.n1047 B.n124 48.9054
R2289 B.n1047 B.n1046 48.9054
R2290 B.n1046 B.n1045 48.9054
R2291 B.n1045 B.n128 48.9054
R2292 B.n1039 B.n128 48.9054
R2293 B.n1039 B.n1038 48.9054
R2294 B.n1038 B.n1037 48.9054
R2295 B.n1037 B.n135 48.9054
R2296 B.n1031 B.n135 48.9054
R2297 B.n809 B.t9 46.0286
R2298 B.n1103 B.t3 46.0286
R2299 B.n731 B.t15 44.5902
R2300 B.n1053 B.t11 44.5902
R2301 B.n869 B.t0 40.2751
R2302 B.n40 B.t4 40.2751
R2303 B.n913 B.t6 38.8367
R2304 B.n1173 B.t2 38.8367
R2305 B.n448 B.t7 33.0832
R2306 B.t8 B.n1078 33.0832
R2307 B.n702 B.n489 32.3127
R2308 B.n698 B.n697 32.3127
R2309 B.n1028 B.n1027 32.3127
R2310 B.n1033 B.n137 32.3127
R2311 B.t1 B.n396 27.3297
R2312 B.n1126 B.t5 27.3297
R2313 B.n839 B.t1 21.5762
R2314 B.t5 B.n1125 21.5762
R2315 B B.n1187 18.0485
R2316 B.n773 B.t7 15.8227
R2317 B.n1079 B.t8 15.8227
R2318 B.n703 B.n702 10.6151
R2319 B.n704 B.n703 10.6151
R2320 B.n704 B.n481 10.6151
R2321 B.n714 B.n481 10.6151
R2322 B.n715 B.n714 10.6151
R2323 B.n716 B.n715 10.6151
R2324 B.n716 B.n473 10.6151
R2325 B.n727 B.n473 10.6151
R2326 B.n728 B.n727 10.6151
R2327 B.n729 B.n728 10.6151
R2328 B.n729 B.n466 10.6151
R2329 B.n739 B.n466 10.6151
R2330 B.n740 B.n739 10.6151
R2331 B.n741 B.n740 10.6151
R2332 B.n741 B.n458 10.6151
R2333 B.n751 B.n458 10.6151
R2334 B.n752 B.n751 10.6151
R2335 B.n753 B.n752 10.6151
R2336 B.n753 B.n450 10.6151
R2337 B.n763 B.n450 10.6151
R2338 B.n764 B.n763 10.6151
R2339 B.n765 B.n764 10.6151
R2340 B.n765 B.n442 10.6151
R2341 B.n775 B.n442 10.6151
R2342 B.n776 B.n775 10.6151
R2343 B.n777 B.n776 10.6151
R2344 B.n777 B.n434 10.6151
R2345 B.n787 B.n434 10.6151
R2346 B.n788 B.n787 10.6151
R2347 B.n789 B.n788 10.6151
R2348 B.n789 B.n426 10.6151
R2349 B.n799 B.n426 10.6151
R2350 B.n800 B.n799 10.6151
R2351 B.n801 B.n800 10.6151
R2352 B.n801 B.n418 10.6151
R2353 B.n811 B.n418 10.6151
R2354 B.n812 B.n811 10.6151
R2355 B.n813 B.n812 10.6151
R2356 B.n813 B.n410 10.6151
R2357 B.n823 B.n410 10.6151
R2358 B.n824 B.n823 10.6151
R2359 B.n825 B.n824 10.6151
R2360 B.n825 B.n402 10.6151
R2361 B.n835 B.n402 10.6151
R2362 B.n836 B.n835 10.6151
R2363 B.n837 B.n836 10.6151
R2364 B.n837 B.n394 10.6151
R2365 B.n847 B.n394 10.6151
R2366 B.n848 B.n847 10.6151
R2367 B.n849 B.n848 10.6151
R2368 B.n849 B.n386 10.6151
R2369 B.n859 B.n386 10.6151
R2370 B.n860 B.n859 10.6151
R2371 B.n861 B.n860 10.6151
R2372 B.n861 B.n378 10.6151
R2373 B.n872 B.n378 10.6151
R2374 B.n873 B.n872 10.6151
R2375 B.n874 B.n873 10.6151
R2376 B.n874 B.n371 10.6151
R2377 B.n884 B.n371 10.6151
R2378 B.n885 B.n884 10.6151
R2379 B.n886 B.n885 10.6151
R2380 B.n886 B.n363 10.6151
R2381 B.n896 B.n363 10.6151
R2382 B.n897 B.n896 10.6151
R2383 B.n898 B.n897 10.6151
R2384 B.n898 B.n355 10.6151
R2385 B.n909 B.n355 10.6151
R2386 B.n910 B.n909 10.6151
R2387 B.n911 B.n910 10.6151
R2388 B.n911 B.n348 10.6151
R2389 B.n922 B.n348 10.6151
R2390 B.n923 B.n922 10.6151
R2391 B.n924 B.n923 10.6151
R2392 B.n924 B.n0 10.6151
R2393 B.n536 B.n489 10.6151
R2394 B.n536 B.n535 10.6151
R2395 B.n542 B.n535 10.6151
R2396 B.n543 B.n542 10.6151
R2397 B.n544 B.n543 10.6151
R2398 B.n544 B.n533 10.6151
R2399 B.n550 B.n533 10.6151
R2400 B.n551 B.n550 10.6151
R2401 B.n552 B.n551 10.6151
R2402 B.n552 B.n531 10.6151
R2403 B.n558 B.n531 10.6151
R2404 B.n559 B.n558 10.6151
R2405 B.n560 B.n559 10.6151
R2406 B.n560 B.n529 10.6151
R2407 B.n566 B.n529 10.6151
R2408 B.n567 B.n566 10.6151
R2409 B.n568 B.n567 10.6151
R2410 B.n568 B.n527 10.6151
R2411 B.n574 B.n527 10.6151
R2412 B.n575 B.n574 10.6151
R2413 B.n576 B.n575 10.6151
R2414 B.n576 B.n525 10.6151
R2415 B.n582 B.n525 10.6151
R2416 B.n583 B.n582 10.6151
R2417 B.n584 B.n583 10.6151
R2418 B.n584 B.n523 10.6151
R2419 B.n590 B.n523 10.6151
R2420 B.n591 B.n590 10.6151
R2421 B.n592 B.n591 10.6151
R2422 B.n592 B.n521 10.6151
R2423 B.n598 B.n521 10.6151
R2424 B.n599 B.n598 10.6151
R2425 B.n600 B.n599 10.6151
R2426 B.n600 B.n519 10.6151
R2427 B.n606 B.n519 10.6151
R2428 B.n609 B.n608 10.6151
R2429 B.n609 B.n515 10.6151
R2430 B.n615 B.n515 10.6151
R2431 B.n616 B.n615 10.6151
R2432 B.n617 B.n616 10.6151
R2433 B.n617 B.n513 10.6151
R2434 B.n623 B.n513 10.6151
R2435 B.n624 B.n623 10.6151
R2436 B.n626 B.n509 10.6151
R2437 B.n632 B.n509 10.6151
R2438 B.n633 B.n632 10.6151
R2439 B.n634 B.n633 10.6151
R2440 B.n634 B.n507 10.6151
R2441 B.n640 B.n507 10.6151
R2442 B.n641 B.n640 10.6151
R2443 B.n642 B.n641 10.6151
R2444 B.n642 B.n505 10.6151
R2445 B.n648 B.n505 10.6151
R2446 B.n649 B.n648 10.6151
R2447 B.n650 B.n649 10.6151
R2448 B.n650 B.n503 10.6151
R2449 B.n656 B.n503 10.6151
R2450 B.n657 B.n656 10.6151
R2451 B.n658 B.n657 10.6151
R2452 B.n658 B.n501 10.6151
R2453 B.n664 B.n501 10.6151
R2454 B.n665 B.n664 10.6151
R2455 B.n666 B.n665 10.6151
R2456 B.n666 B.n499 10.6151
R2457 B.n672 B.n499 10.6151
R2458 B.n673 B.n672 10.6151
R2459 B.n674 B.n673 10.6151
R2460 B.n674 B.n497 10.6151
R2461 B.n680 B.n497 10.6151
R2462 B.n681 B.n680 10.6151
R2463 B.n682 B.n681 10.6151
R2464 B.n682 B.n495 10.6151
R2465 B.n688 B.n495 10.6151
R2466 B.n689 B.n688 10.6151
R2467 B.n690 B.n689 10.6151
R2468 B.n690 B.n493 10.6151
R2469 B.n696 B.n493 10.6151
R2470 B.n697 B.n696 10.6151
R2471 B.n698 B.n485 10.6151
R2472 B.n708 B.n485 10.6151
R2473 B.n709 B.n708 10.6151
R2474 B.n710 B.n709 10.6151
R2475 B.n710 B.n477 10.6151
R2476 B.n720 B.n477 10.6151
R2477 B.n721 B.n720 10.6151
R2478 B.n722 B.n721 10.6151
R2479 B.n722 B.n470 10.6151
R2480 B.n733 B.n470 10.6151
R2481 B.n734 B.n733 10.6151
R2482 B.n735 B.n734 10.6151
R2483 B.n735 B.n462 10.6151
R2484 B.n745 B.n462 10.6151
R2485 B.n746 B.n745 10.6151
R2486 B.n747 B.n746 10.6151
R2487 B.n747 B.n454 10.6151
R2488 B.n757 B.n454 10.6151
R2489 B.n758 B.n757 10.6151
R2490 B.n759 B.n758 10.6151
R2491 B.n759 B.n445 10.6151
R2492 B.n769 B.n445 10.6151
R2493 B.n770 B.n769 10.6151
R2494 B.n771 B.n770 10.6151
R2495 B.n771 B.n438 10.6151
R2496 B.n781 B.n438 10.6151
R2497 B.n782 B.n781 10.6151
R2498 B.n783 B.n782 10.6151
R2499 B.n783 B.n430 10.6151
R2500 B.n793 B.n430 10.6151
R2501 B.n794 B.n793 10.6151
R2502 B.n795 B.n794 10.6151
R2503 B.n795 B.n421 10.6151
R2504 B.n805 B.n421 10.6151
R2505 B.n806 B.n805 10.6151
R2506 B.n807 B.n806 10.6151
R2507 B.n807 B.n414 10.6151
R2508 B.n817 B.n414 10.6151
R2509 B.n818 B.n817 10.6151
R2510 B.n819 B.n818 10.6151
R2511 B.n819 B.n406 10.6151
R2512 B.n829 B.n406 10.6151
R2513 B.n830 B.n829 10.6151
R2514 B.n831 B.n830 10.6151
R2515 B.n831 B.n398 10.6151
R2516 B.n841 B.n398 10.6151
R2517 B.n842 B.n841 10.6151
R2518 B.n843 B.n842 10.6151
R2519 B.n843 B.n390 10.6151
R2520 B.n853 B.n390 10.6151
R2521 B.n854 B.n853 10.6151
R2522 B.n855 B.n854 10.6151
R2523 B.n855 B.n382 10.6151
R2524 B.n865 B.n382 10.6151
R2525 B.n866 B.n865 10.6151
R2526 B.n867 B.n866 10.6151
R2527 B.n867 B.n375 10.6151
R2528 B.n878 B.n375 10.6151
R2529 B.n879 B.n878 10.6151
R2530 B.n880 B.n879 10.6151
R2531 B.n880 B.n367 10.6151
R2532 B.n890 B.n367 10.6151
R2533 B.n891 B.n890 10.6151
R2534 B.n892 B.n891 10.6151
R2535 B.n892 B.n359 10.6151
R2536 B.n902 B.n359 10.6151
R2537 B.n903 B.n902 10.6151
R2538 B.n904 B.n903 10.6151
R2539 B.n904 B.n352 10.6151
R2540 B.n915 B.n352 10.6151
R2541 B.n916 B.n915 10.6151
R2542 B.n918 B.n916 10.6151
R2543 B.n918 B.n917 10.6151
R2544 B.n917 B.n344 10.6151
R2545 B.n929 B.n344 10.6151
R2546 B.n930 B.n929 10.6151
R2547 B.n931 B.n930 10.6151
R2548 B.n932 B.n931 10.6151
R2549 B.n933 B.n932 10.6151
R2550 B.n936 B.n933 10.6151
R2551 B.n937 B.n936 10.6151
R2552 B.n938 B.n937 10.6151
R2553 B.n939 B.n938 10.6151
R2554 B.n941 B.n939 10.6151
R2555 B.n942 B.n941 10.6151
R2556 B.n943 B.n942 10.6151
R2557 B.n944 B.n943 10.6151
R2558 B.n946 B.n944 10.6151
R2559 B.n947 B.n946 10.6151
R2560 B.n948 B.n947 10.6151
R2561 B.n949 B.n948 10.6151
R2562 B.n951 B.n949 10.6151
R2563 B.n952 B.n951 10.6151
R2564 B.n953 B.n952 10.6151
R2565 B.n954 B.n953 10.6151
R2566 B.n956 B.n954 10.6151
R2567 B.n957 B.n956 10.6151
R2568 B.n958 B.n957 10.6151
R2569 B.n959 B.n958 10.6151
R2570 B.n961 B.n959 10.6151
R2571 B.n962 B.n961 10.6151
R2572 B.n963 B.n962 10.6151
R2573 B.n964 B.n963 10.6151
R2574 B.n966 B.n964 10.6151
R2575 B.n967 B.n966 10.6151
R2576 B.n968 B.n967 10.6151
R2577 B.n969 B.n968 10.6151
R2578 B.n971 B.n969 10.6151
R2579 B.n972 B.n971 10.6151
R2580 B.n973 B.n972 10.6151
R2581 B.n974 B.n973 10.6151
R2582 B.n976 B.n974 10.6151
R2583 B.n977 B.n976 10.6151
R2584 B.n978 B.n977 10.6151
R2585 B.n979 B.n978 10.6151
R2586 B.n981 B.n979 10.6151
R2587 B.n982 B.n981 10.6151
R2588 B.n983 B.n982 10.6151
R2589 B.n984 B.n983 10.6151
R2590 B.n986 B.n984 10.6151
R2591 B.n987 B.n986 10.6151
R2592 B.n988 B.n987 10.6151
R2593 B.n989 B.n988 10.6151
R2594 B.n991 B.n989 10.6151
R2595 B.n992 B.n991 10.6151
R2596 B.n993 B.n992 10.6151
R2597 B.n994 B.n993 10.6151
R2598 B.n996 B.n994 10.6151
R2599 B.n997 B.n996 10.6151
R2600 B.n998 B.n997 10.6151
R2601 B.n999 B.n998 10.6151
R2602 B.n1001 B.n999 10.6151
R2603 B.n1002 B.n1001 10.6151
R2604 B.n1003 B.n1002 10.6151
R2605 B.n1004 B.n1003 10.6151
R2606 B.n1006 B.n1004 10.6151
R2607 B.n1007 B.n1006 10.6151
R2608 B.n1008 B.n1007 10.6151
R2609 B.n1009 B.n1008 10.6151
R2610 B.n1011 B.n1009 10.6151
R2611 B.n1012 B.n1011 10.6151
R2612 B.n1013 B.n1012 10.6151
R2613 B.n1014 B.n1013 10.6151
R2614 B.n1016 B.n1014 10.6151
R2615 B.n1017 B.n1016 10.6151
R2616 B.n1018 B.n1017 10.6151
R2617 B.n1019 B.n1018 10.6151
R2618 B.n1021 B.n1019 10.6151
R2619 B.n1022 B.n1021 10.6151
R2620 B.n1023 B.n1022 10.6151
R2621 B.n1024 B.n1023 10.6151
R2622 B.n1026 B.n1024 10.6151
R2623 B.n1027 B.n1026 10.6151
R2624 B.n1179 B.n1 10.6151
R2625 B.n1179 B.n1178 10.6151
R2626 B.n1178 B.n1177 10.6151
R2627 B.n1177 B.n10 10.6151
R2628 B.n1171 B.n10 10.6151
R2629 B.n1171 B.n1170 10.6151
R2630 B.n1170 B.n1169 10.6151
R2631 B.n1169 B.n17 10.6151
R2632 B.n1163 B.n17 10.6151
R2633 B.n1163 B.n1162 10.6151
R2634 B.n1162 B.n1161 10.6151
R2635 B.n1161 B.n25 10.6151
R2636 B.n1155 B.n25 10.6151
R2637 B.n1155 B.n1154 10.6151
R2638 B.n1154 B.n1153 10.6151
R2639 B.n1153 B.n32 10.6151
R2640 B.n1147 B.n32 10.6151
R2641 B.n1147 B.n1146 10.6151
R2642 B.n1146 B.n1145 10.6151
R2643 B.n1145 B.n38 10.6151
R2644 B.n1139 B.n38 10.6151
R2645 B.n1139 B.n1138 10.6151
R2646 B.n1138 B.n1137 10.6151
R2647 B.n1137 B.n46 10.6151
R2648 B.n1131 B.n46 10.6151
R2649 B.n1131 B.n1130 10.6151
R2650 B.n1130 B.n1129 10.6151
R2651 B.n1129 B.n53 10.6151
R2652 B.n1123 B.n53 10.6151
R2653 B.n1123 B.n1122 10.6151
R2654 B.n1122 B.n1121 10.6151
R2655 B.n1121 B.n60 10.6151
R2656 B.n1115 B.n60 10.6151
R2657 B.n1115 B.n1114 10.6151
R2658 B.n1114 B.n1113 10.6151
R2659 B.n1113 B.n67 10.6151
R2660 B.n1107 B.n67 10.6151
R2661 B.n1107 B.n1106 10.6151
R2662 B.n1106 B.n1105 10.6151
R2663 B.n1105 B.n74 10.6151
R2664 B.n1099 B.n74 10.6151
R2665 B.n1099 B.n1098 10.6151
R2666 B.n1098 B.n1097 10.6151
R2667 B.n1097 B.n81 10.6151
R2668 B.n1091 B.n81 10.6151
R2669 B.n1091 B.n1090 10.6151
R2670 B.n1090 B.n1089 10.6151
R2671 B.n1089 B.n88 10.6151
R2672 B.n1083 B.n88 10.6151
R2673 B.n1083 B.n1082 10.6151
R2674 B.n1082 B.n1081 10.6151
R2675 B.n1081 B.n95 10.6151
R2676 B.n1075 B.n95 10.6151
R2677 B.n1075 B.n1074 10.6151
R2678 B.n1074 B.n1073 10.6151
R2679 B.n1073 B.n102 10.6151
R2680 B.n1067 B.n102 10.6151
R2681 B.n1067 B.n1066 10.6151
R2682 B.n1066 B.n1065 10.6151
R2683 B.n1065 B.n109 10.6151
R2684 B.n1059 B.n109 10.6151
R2685 B.n1059 B.n1058 10.6151
R2686 B.n1058 B.n1057 10.6151
R2687 B.n1057 B.n116 10.6151
R2688 B.n1051 B.n116 10.6151
R2689 B.n1051 B.n1050 10.6151
R2690 B.n1050 B.n1049 10.6151
R2691 B.n1049 B.n122 10.6151
R2692 B.n1043 B.n122 10.6151
R2693 B.n1043 B.n1042 10.6151
R2694 B.n1042 B.n1041 10.6151
R2695 B.n1041 B.n130 10.6151
R2696 B.n1035 B.n130 10.6151
R2697 B.n1035 B.n1034 10.6151
R2698 B.n1034 B.n1033 10.6151
R2699 B.n186 B.n137 10.6151
R2700 B.n189 B.n186 10.6151
R2701 B.n190 B.n189 10.6151
R2702 B.n193 B.n190 10.6151
R2703 B.n194 B.n193 10.6151
R2704 B.n197 B.n194 10.6151
R2705 B.n198 B.n197 10.6151
R2706 B.n201 B.n198 10.6151
R2707 B.n202 B.n201 10.6151
R2708 B.n205 B.n202 10.6151
R2709 B.n206 B.n205 10.6151
R2710 B.n209 B.n206 10.6151
R2711 B.n210 B.n209 10.6151
R2712 B.n213 B.n210 10.6151
R2713 B.n214 B.n213 10.6151
R2714 B.n217 B.n214 10.6151
R2715 B.n218 B.n217 10.6151
R2716 B.n221 B.n218 10.6151
R2717 B.n222 B.n221 10.6151
R2718 B.n225 B.n222 10.6151
R2719 B.n226 B.n225 10.6151
R2720 B.n229 B.n226 10.6151
R2721 B.n230 B.n229 10.6151
R2722 B.n233 B.n230 10.6151
R2723 B.n234 B.n233 10.6151
R2724 B.n237 B.n234 10.6151
R2725 B.n238 B.n237 10.6151
R2726 B.n241 B.n238 10.6151
R2727 B.n242 B.n241 10.6151
R2728 B.n245 B.n242 10.6151
R2729 B.n246 B.n245 10.6151
R2730 B.n249 B.n246 10.6151
R2731 B.n250 B.n249 10.6151
R2732 B.n253 B.n250 10.6151
R2733 B.n254 B.n253 10.6151
R2734 B.n258 B.n257 10.6151
R2735 B.n261 B.n258 10.6151
R2736 B.n262 B.n261 10.6151
R2737 B.n265 B.n262 10.6151
R2738 B.n266 B.n265 10.6151
R2739 B.n269 B.n266 10.6151
R2740 B.n270 B.n269 10.6151
R2741 B.n273 B.n270 10.6151
R2742 B.n278 B.n275 10.6151
R2743 B.n279 B.n278 10.6151
R2744 B.n282 B.n279 10.6151
R2745 B.n283 B.n282 10.6151
R2746 B.n286 B.n283 10.6151
R2747 B.n287 B.n286 10.6151
R2748 B.n290 B.n287 10.6151
R2749 B.n291 B.n290 10.6151
R2750 B.n294 B.n291 10.6151
R2751 B.n295 B.n294 10.6151
R2752 B.n298 B.n295 10.6151
R2753 B.n299 B.n298 10.6151
R2754 B.n302 B.n299 10.6151
R2755 B.n303 B.n302 10.6151
R2756 B.n306 B.n303 10.6151
R2757 B.n307 B.n306 10.6151
R2758 B.n310 B.n307 10.6151
R2759 B.n311 B.n310 10.6151
R2760 B.n314 B.n311 10.6151
R2761 B.n315 B.n314 10.6151
R2762 B.n318 B.n315 10.6151
R2763 B.n319 B.n318 10.6151
R2764 B.n322 B.n319 10.6151
R2765 B.n323 B.n322 10.6151
R2766 B.n326 B.n323 10.6151
R2767 B.n327 B.n326 10.6151
R2768 B.n330 B.n327 10.6151
R2769 B.n331 B.n330 10.6151
R2770 B.n334 B.n331 10.6151
R2771 B.n335 B.n334 10.6151
R2772 B.n338 B.n335 10.6151
R2773 B.n339 B.n338 10.6151
R2774 B.n342 B.n339 10.6151
R2775 B.n343 B.n342 10.6151
R2776 B.n1028 B.n343 10.6151
R2777 B.n906 B.t6 10.0691
R2778 B.n19 B.t2 10.0691
R2779 B.n876 B.t0 8.63077
R2780 B.n1149 B.t4 8.63077
R2781 B.n1187 B.n0 8.11757
R2782 B.n1187 B.n1 8.11757
R2783 B.n608 B.n607 6.5566
R2784 B.n625 B.n624 6.5566
R2785 B.n257 B.n185 6.5566
R2786 B.n274 B.n273 6.5566
R2787 B.n724 B.t15 4.31564
R2788 B.n124 B.t11 4.31564
R2789 B.n607 B.n606 4.05904
R2790 B.n626 B.n625 4.05904
R2791 B.n254 B.n185 4.05904
R2792 B.n275 B.n274 4.05904
R2793 B.n424 B.t9 2.87726
R2794 B.t3 B.n1102 2.87726
R2795 VN.n100 VN.n99 161.3
R2796 VN.n98 VN.n52 161.3
R2797 VN.n97 VN.n96 161.3
R2798 VN.n95 VN.n53 161.3
R2799 VN.n94 VN.n93 161.3
R2800 VN.n92 VN.n54 161.3
R2801 VN.n91 VN.n90 161.3
R2802 VN.n89 VN.n55 161.3
R2803 VN.n88 VN.n87 161.3
R2804 VN.n86 VN.n56 161.3
R2805 VN.n85 VN.n84 161.3
R2806 VN.n83 VN.n58 161.3
R2807 VN.n82 VN.n81 161.3
R2808 VN.n80 VN.n59 161.3
R2809 VN.n79 VN.n78 161.3
R2810 VN.n77 VN.n60 161.3
R2811 VN.n76 VN.n75 161.3
R2812 VN.n74 VN.n61 161.3
R2813 VN.n73 VN.n72 161.3
R2814 VN.n71 VN.n62 161.3
R2815 VN.n70 VN.n69 161.3
R2816 VN.n68 VN.n63 161.3
R2817 VN.n67 VN.n66 161.3
R2818 VN.n49 VN.n48 161.3
R2819 VN.n47 VN.n1 161.3
R2820 VN.n46 VN.n45 161.3
R2821 VN.n44 VN.n2 161.3
R2822 VN.n43 VN.n42 161.3
R2823 VN.n41 VN.n3 161.3
R2824 VN.n40 VN.n39 161.3
R2825 VN.n38 VN.n4 161.3
R2826 VN.n37 VN.n36 161.3
R2827 VN.n34 VN.n5 161.3
R2828 VN.n33 VN.n32 161.3
R2829 VN.n31 VN.n6 161.3
R2830 VN.n30 VN.n29 161.3
R2831 VN.n28 VN.n7 161.3
R2832 VN.n27 VN.n26 161.3
R2833 VN.n25 VN.n8 161.3
R2834 VN.n24 VN.n23 161.3
R2835 VN.n22 VN.n9 161.3
R2836 VN.n21 VN.n20 161.3
R2837 VN.n19 VN.n10 161.3
R2838 VN.n18 VN.n17 161.3
R2839 VN.n16 VN.n11 161.3
R2840 VN.n15 VN.n14 161.3
R2841 VN.n65 VN.t5 101.947
R2842 VN.n13 VN.t8 101.947
R2843 VN.n50 VN.n0 78.4415
R2844 VN.n101 VN.n51 78.4415
R2845 VN.n8 VN.t6 68.2158
R2846 VN.n12 VN.t2 68.2158
R2847 VN.n35 VN.t0 68.2158
R2848 VN.n0 VN.t9 68.2158
R2849 VN.n60 VN.t4 68.2158
R2850 VN.n64 VN.t7 68.2158
R2851 VN.n57 VN.t3 68.2158
R2852 VN.n51 VN.t1 68.2158
R2853 VN VN.n101 57.0171
R2854 VN.n13 VN.n12 56.696
R2855 VN.n65 VN.n64 56.696
R2856 VN.n42 VN.n2 56.5617
R2857 VN.n93 VN.n53 56.5617
R2858 VN.n21 VN.n10 46.874
R2859 VN.n29 VN.n6 46.874
R2860 VN.n73 VN.n62 46.874
R2861 VN.n81 VN.n58 46.874
R2862 VN.n17 VN.n10 34.28
R2863 VN.n33 VN.n6 34.28
R2864 VN.n69 VN.n62 34.28
R2865 VN.n85 VN.n58 34.28
R2866 VN.n16 VN.n15 24.5923
R2867 VN.n17 VN.n16 24.5923
R2868 VN.n22 VN.n21 24.5923
R2869 VN.n23 VN.n22 24.5923
R2870 VN.n23 VN.n8 24.5923
R2871 VN.n27 VN.n8 24.5923
R2872 VN.n28 VN.n27 24.5923
R2873 VN.n29 VN.n28 24.5923
R2874 VN.n34 VN.n33 24.5923
R2875 VN.n36 VN.n34 24.5923
R2876 VN.n40 VN.n4 24.5923
R2877 VN.n41 VN.n40 24.5923
R2878 VN.n42 VN.n41 24.5923
R2879 VN.n46 VN.n2 24.5923
R2880 VN.n47 VN.n46 24.5923
R2881 VN.n48 VN.n47 24.5923
R2882 VN.n69 VN.n68 24.5923
R2883 VN.n68 VN.n67 24.5923
R2884 VN.n81 VN.n80 24.5923
R2885 VN.n80 VN.n79 24.5923
R2886 VN.n79 VN.n60 24.5923
R2887 VN.n75 VN.n60 24.5923
R2888 VN.n75 VN.n74 24.5923
R2889 VN.n74 VN.n73 24.5923
R2890 VN.n93 VN.n92 24.5923
R2891 VN.n92 VN.n91 24.5923
R2892 VN.n91 VN.n55 24.5923
R2893 VN.n87 VN.n86 24.5923
R2894 VN.n86 VN.n85 24.5923
R2895 VN.n99 VN.n98 24.5923
R2896 VN.n98 VN.n97 24.5923
R2897 VN.n97 VN.n53 24.5923
R2898 VN.n15 VN.n12 18.1985
R2899 VN.n36 VN.n35 18.1985
R2900 VN.n67 VN.n64 18.1985
R2901 VN.n87 VN.n57 18.1985
R2902 VN.n48 VN.n0 11.8046
R2903 VN.n99 VN.n51 11.8046
R2904 VN.n35 VN.n4 6.39438
R2905 VN.n57 VN.n55 6.39438
R2906 VN.n66 VN.n65 3.08737
R2907 VN.n14 VN.n13 3.08737
R2908 VN.n101 VN.n100 0.354861
R2909 VN.n50 VN.n49 0.354861
R2910 VN VN.n50 0.267071
R2911 VN.n100 VN.n52 0.189894
R2912 VN.n96 VN.n52 0.189894
R2913 VN.n96 VN.n95 0.189894
R2914 VN.n95 VN.n94 0.189894
R2915 VN.n94 VN.n54 0.189894
R2916 VN.n90 VN.n54 0.189894
R2917 VN.n90 VN.n89 0.189894
R2918 VN.n89 VN.n88 0.189894
R2919 VN.n88 VN.n56 0.189894
R2920 VN.n84 VN.n56 0.189894
R2921 VN.n84 VN.n83 0.189894
R2922 VN.n83 VN.n82 0.189894
R2923 VN.n82 VN.n59 0.189894
R2924 VN.n78 VN.n59 0.189894
R2925 VN.n78 VN.n77 0.189894
R2926 VN.n77 VN.n76 0.189894
R2927 VN.n76 VN.n61 0.189894
R2928 VN.n72 VN.n61 0.189894
R2929 VN.n72 VN.n71 0.189894
R2930 VN.n71 VN.n70 0.189894
R2931 VN.n70 VN.n63 0.189894
R2932 VN.n66 VN.n63 0.189894
R2933 VN.n14 VN.n11 0.189894
R2934 VN.n18 VN.n11 0.189894
R2935 VN.n19 VN.n18 0.189894
R2936 VN.n20 VN.n19 0.189894
R2937 VN.n20 VN.n9 0.189894
R2938 VN.n24 VN.n9 0.189894
R2939 VN.n25 VN.n24 0.189894
R2940 VN.n26 VN.n25 0.189894
R2941 VN.n26 VN.n7 0.189894
R2942 VN.n30 VN.n7 0.189894
R2943 VN.n31 VN.n30 0.189894
R2944 VN.n32 VN.n31 0.189894
R2945 VN.n32 VN.n5 0.189894
R2946 VN.n37 VN.n5 0.189894
R2947 VN.n38 VN.n37 0.189894
R2948 VN.n39 VN.n38 0.189894
R2949 VN.n39 VN.n3 0.189894
R2950 VN.n43 VN.n3 0.189894
R2951 VN.n44 VN.n43 0.189894
R2952 VN.n45 VN.n44 0.189894
R2953 VN.n45 VN.n1 0.189894
R2954 VN.n49 VN.n1 0.189894
R2955 VDD2.n105 VDD2.n57 289.615
R2956 VDD2.n48 VDD2.n0 289.615
R2957 VDD2.n106 VDD2.n105 185
R2958 VDD2.n104 VDD2.n103 185
R2959 VDD2.n61 VDD2.n60 185
R2960 VDD2.n98 VDD2.n97 185
R2961 VDD2.n96 VDD2.n63 185
R2962 VDD2.n95 VDD2.n94 185
R2963 VDD2.n66 VDD2.n64 185
R2964 VDD2.n89 VDD2.n88 185
R2965 VDD2.n87 VDD2.n86 185
R2966 VDD2.n70 VDD2.n69 185
R2967 VDD2.n81 VDD2.n80 185
R2968 VDD2.n79 VDD2.n78 185
R2969 VDD2.n74 VDD2.n73 185
R2970 VDD2.n16 VDD2.n15 185
R2971 VDD2.n21 VDD2.n20 185
R2972 VDD2.n23 VDD2.n22 185
R2973 VDD2.n12 VDD2.n11 185
R2974 VDD2.n29 VDD2.n28 185
R2975 VDD2.n31 VDD2.n30 185
R2976 VDD2.n8 VDD2.n7 185
R2977 VDD2.n38 VDD2.n37 185
R2978 VDD2.n39 VDD2.n6 185
R2979 VDD2.n41 VDD2.n40 185
R2980 VDD2.n4 VDD2.n3 185
R2981 VDD2.n47 VDD2.n46 185
R2982 VDD2.n49 VDD2.n48 185
R2983 VDD2.n75 VDD2.t8 149.524
R2984 VDD2.n17 VDD2.t1 149.524
R2985 VDD2.n105 VDD2.n104 104.615
R2986 VDD2.n104 VDD2.n60 104.615
R2987 VDD2.n97 VDD2.n60 104.615
R2988 VDD2.n97 VDD2.n96 104.615
R2989 VDD2.n96 VDD2.n95 104.615
R2990 VDD2.n95 VDD2.n64 104.615
R2991 VDD2.n88 VDD2.n64 104.615
R2992 VDD2.n88 VDD2.n87 104.615
R2993 VDD2.n87 VDD2.n69 104.615
R2994 VDD2.n80 VDD2.n69 104.615
R2995 VDD2.n80 VDD2.n79 104.615
R2996 VDD2.n79 VDD2.n73 104.615
R2997 VDD2.n21 VDD2.n15 104.615
R2998 VDD2.n22 VDD2.n21 104.615
R2999 VDD2.n22 VDD2.n11 104.615
R3000 VDD2.n29 VDD2.n11 104.615
R3001 VDD2.n30 VDD2.n29 104.615
R3002 VDD2.n30 VDD2.n7 104.615
R3003 VDD2.n38 VDD2.n7 104.615
R3004 VDD2.n39 VDD2.n38 104.615
R3005 VDD2.n40 VDD2.n39 104.615
R3006 VDD2.n40 VDD2.n3 104.615
R3007 VDD2.n47 VDD2.n3 104.615
R3008 VDD2.n48 VDD2.n47 104.615
R3009 VDD2.n56 VDD2.n55 66.2506
R3010 VDD2 VDD2.n113 66.2478
R3011 VDD2.n112 VDD2.n111 63.804
R3012 VDD2.n54 VDD2.n53 63.8038
R3013 VDD2.n54 VDD2.n52 53.364
R3014 VDD2.t8 VDD2.n73 52.3082
R3015 VDD2.t1 VDD2.n15 52.3082
R3016 VDD2.n110 VDD2.n109 50.0278
R3017 VDD2.n110 VDD2.n56 48.2002
R3018 VDD2.n98 VDD2.n63 13.1884
R3019 VDD2.n41 VDD2.n6 13.1884
R3020 VDD2.n99 VDD2.n61 12.8005
R3021 VDD2.n94 VDD2.n65 12.8005
R3022 VDD2.n37 VDD2.n36 12.8005
R3023 VDD2.n42 VDD2.n4 12.8005
R3024 VDD2.n103 VDD2.n102 12.0247
R3025 VDD2.n93 VDD2.n66 12.0247
R3026 VDD2.n35 VDD2.n8 12.0247
R3027 VDD2.n46 VDD2.n45 12.0247
R3028 VDD2.n106 VDD2.n59 11.249
R3029 VDD2.n90 VDD2.n89 11.249
R3030 VDD2.n32 VDD2.n31 11.249
R3031 VDD2.n49 VDD2.n2 11.249
R3032 VDD2.n107 VDD2.n57 10.4732
R3033 VDD2.n86 VDD2.n68 10.4732
R3034 VDD2.n28 VDD2.n10 10.4732
R3035 VDD2.n50 VDD2.n0 10.4732
R3036 VDD2.n75 VDD2.n74 10.2747
R3037 VDD2.n17 VDD2.n16 10.2747
R3038 VDD2.n85 VDD2.n70 9.69747
R3039 VDD2.n27 VDD2.n12 9.69747
R3040 VDD2.n109 VDD2.n108 9.45567
R3041 VDD2.n52 VDD2.n51 9.45567
R3042 VDD2.n77 VDD2.n76 9.3005
R3043 VDD2.n72 VDD2.n71 9.3005
R3044 VDD2.n83 VDD2.n82 9.3005
R3045 VDD2.n85 VDD2.n84 9.3005
R3046 VDD2.n68 VDD2.n67 9.3005
R3047 VDD2.n91 VDD2.n90 9.3005
R3048 VDD2.n93 VDD2.n92 9.3005
R3049 VDD2.n65 VDD2.n62 9.3005
R3050 VDD2.n108 VDD2.n107 9.3005
R3051 VDD2.n59 VDD2.n58 9.3005
R3052 VDD2.n102 VDD2.n101 9.3005
R3053 VDD2.n100 VDD2.n99 9.3005
R3054 VDD2.n51 VDD2.n50 9.3005
R3055 VDD2.n2 VDD2.n1 9.3005
R3056 VDD2.n45 VDD2.n44 9.3005
R3057 VDD2.n43 VDD2.n42 9.3005
R3058 VDD2.n19 VDD2.n18 9.3005
R3059 VDD2.n14 VDD2.n13 9.3005
R3060 VDD2.n25 VDD2.n24 9.3005
R3061 VDD2.n27 VDD2.n26 9.3005
R3062 VDD2.n10 VDD2.n9 9.3005
R3063 VDD2.n33 VDD2.n32 9.3005
R3064 VDD2.n35 VDD2.n34 9.3005
R3065 VDD2.n36 VDD2.n5 9.3005
R3066 VDD2.n82 VDD2.n81 8.92171
R3067 VDD2.n24 VDD2.n23 8.92171
R3068 VDD2.n78 VDD2.n72 8.14595
R3069 VDD2.n20 VDD2.n14 8.14595
R3070 VDD2.n77 VDD2.n74 7.3702
R3071 VDD2.n19 VDD2.n16 7.3702
R3072 VDD2.n78 VDD2.n77 5.81868
R3073 VDD2.n20 VDD2.n19 5.81868
R3074 VDD2.n81 VDD2.n72 5.04292
R3075 VDD2.n23 VDD2.n14 5.04292
R3076 VDD2.n82 VDD2.n70 4.26717
R3077 VDD2.n24 VDD2.n12 4.26717
R3078 VDD2.n109 VDD2.n57 3.49141
R3079 VDD2.n86 VDD2.n85 3.49141
R3080 VDD2.n28 VDD2.n27 3.49141
R3081 VDD2.n52 VDD2.n0 3.49141
R3082 VDD2.n112 VDD2.n110 3.33671
R3083 VDD2.n76 VDD2.n75 2.84303
R3084 VDD2.n18 VDD2.n17 2.84303
R3085 VDD2.n107 VDD2.n106 2.71565
R3086 VDD2.n89 VDD2.n68 2.71565
R3087 VDD2.n31 VDD2.n10 2.71565
R3088 VDD2.n50 VDD2.n49 2.71565
R3089 VDD2.n113 VDD2.t2 1.97655
R3090 VDD2.n113 VDD2.t4 1.97655
R3091 VDD2.n111 VDD2.t6 1.97655
R3092 VDD2.n111 VDD2.t5 1.97655
R3093 VDD2.n55 VDD2.t9 1.97655
R3094 VDD2.n55 VDD2.t0 1.97655
R3095 VDD2.n53 VDD2.t7 1.97655
R3096 VDD2.n53 VDD2.t3 1.97655
R3097 VDD2.n103 VDD2.n59 1.93989
R3098 VDD2.n90 VDD2.n66 1.93989
R3099 VDD2.n32 VDD2.n8 1.93989
R3100 VDD2.n46 VDD2.n2 1.93989
R3101 VDD2.n102 VDD2.n61 1.16414
R3102 VDD2.n94 VDD2.n93 1.16414
R3103 VDD2.n37 VDD2.n35 1.16414
R3104 VDD2.n45 VDD2.n4 1.16414
R3105 VDD2 VDD2.n112 0.892741
R3106 VDD2.n56 VDD2.n54 0.779206
R3107 VDD2.n99 VDD2.n98 0.388379
R3108 VDD2.n65 VDD2.n63 0.388379
R3109 VDD2.n36 VDD2.n6 0.388379
R3110 VDD2.n42 VDD2.n41 0.388379
R3111 VDD2.n108 VDD2.n58 0.155672
R3112 VDD2.n101 VDD2.n58 0.155672
R3113 VDD2.n101 VDD2.n100 0.155672
R3114 VDD2.n100 VDD2.n62 0.155672
R3115 VDD2.n92 VDD2.n62 0.155672
R3116 VDD2.n92 VDD2.n91 0.155672
R3117 VDD2.n91 VDD2.n67 0.155672
R3118 VDD2.n84 VDD2.n67 0.155672
R3119 VDD2.n84 VDD2.n83 0.155672
R3120 VDD2.n83 VDD2.n71 0.155672
R3121 VDD2.n76 VDD2.n71 0.155672
R3122 VDD2.n18 VDD2.n13 0.155672
R3123 VDD2.n25 VDD2.n13 0.155672
R3124 VDD2.n26 VDD2.n25 0.155672
R3125 VDD2.n26 VDD2.n9 0.155672
R3126 VDD2.n33 VDD2.n9 0.155672
R3127 VDD2.n34 VDD2.n33 0.155672
R3128 VDD2.n34 VDD2.n5 0.155672
R3129 VDD2.n43 VDD2.n5 0.155672
R3130 VDD2.n44 VDD2.n43 0.155672
R3131 VDD2.n44 VDD2.n1 0.155672
R3132 VDD2.n51 VDD2.n1 0.155672
C0 VN VDD1 0.155832f
C1 VN VTAIL 10.627201f
C2 VN VDD2 9.48831f
C3 VTAIL VDD1 10.038301f
C4 VDD1 VDD2 2.78652f
C5 VTAIL VDD2 10.096701f
C6 VN VP 9.40825f
C7 VP VDD1 10.032499f
C8 VTAIL VP 10.6414f
C9 VP VDD2 0.703721f
C10 VDD2 B 7.972547f
C11 VDD1 B 7.930423f
C12 VTAIL B 8.119215f
C13 VN B 22.471891f
C14 VP B 21.0623f
C15 VDD2.n0 B 0.034434f
C16 VDD2.n1 B 0.025225f
C17 VDD2.n2 B 0.013555f
C18 VDD2.n3 B 0.032038f
C19 VDD2.n4 B 0.014352f
C20 VDD2.n5 B 0.025225f
C21 VDD2.n6 B 0.013953f
C22 VDD2.n7 B 0.032038f
C23 VDD2.n8 B 0.014352f
C24 VDD2.n9 B 0.025225f
C25 VDD2.n10 B 0.013555f
C26 VDD2.n11 B 0.032038f
C27 VDD2.n12 B 0.014352f
C28 VDD2.n13 B 0.025225f
C29 VDD2.n14 B 0.013555f
C30 VDD2.n15 B 0.024029f
C31 VDD2.n16 B 0.022648f
C32 VDD2.t1 B 0.053843f
C33 VDD2.n17 B 0.162695f
C34 VDD2.n18 B 1.05038f
C35 VDD2.n19 B 0.013555f
C36 VDD2.n20 B 0.014352f
C37 VDD2.n21 B 0.032038f
C38 VDD2.n22 B 0.032038f
C39 VDD2.n23 B 0.014352f
C40 VDD2.n24 B 0.013555f
C41 VDD2.n25 B 0.025225f
C42 VDD2.n26 B 0.025225f
C43 VDD2.n27 B 0.013555f
C44 VDD2.n28 B 0.014352f
C45 VDD2.n29 B 0.032038f
C46 VDD2.n30 B 0.032038f
C47 VDD2.n31 B 0.014352f
C48 VDD2.n32 B 0.013555f
C49 VDD2.n33 B 0.025225f
C50 VDD2.n34 B 0.025225f
C51 VDD2.n35 B 0.013555f
C52 VDD2.n36 B 0.013555f
C53 VDD2.n37 B 0.014352f
C54 VDD2.n38 B 0.032038f
C55 VDD2.n39 B 0.032038f
C56 VDD2.n40 B 0.032038f
C57 VDD2.n41 B 0.013953f
C58 VDD2.n42 B 0.013555f
C59 VDD2.n43 B 0.025225f
C60 VDD2.n44 B 0.025225f
C61 VDD2.n45 B 0.013555f
C62 VDD2.n46 B 0.014352f
C63 VDD2.n47 B 0.032038f
C64 VDD2.n48 B 0.067551f
C65 VDD2.n49 B 0.014352f
C66 VDD2.n50 B 0.013555f
C67 VDD2.n51 B 0.060373f
C68 VDD2.n52 B 0.075139f
C69 VDD2.t7 B 0.19973f
C70 VDD2.t3 B 0.19973f
C71 VDD2.n53 B 1.75989f
C72 VDD2.n54 B 0.84082f
C73 VDD2.t9 B 0.19973f
C74 VDD2.t0 B 0.19973f
C75 VDD2.n55 B 1.7852f
C76 VDD2.n56 B 3.29877f
C77 VDD2.n57 B 0.034434f
C78 VDD2.n58 B 0.025225f
C79 VDD2.n59 B 0.013555f
C80 VDD2.n60 B 0.032038f
C81 VDD2.n61 B 0.014352f
C82 VDD2.n62 B 0.025225f
C83 VDD2.n63 B 0.013953f
C84 VDD2.n64 B 0.032038f
C85 VDD2.n65 B 0.013555f
C86 VDD2.n66 B 0.014352f
C87 VDD2.n67 B 0.025225f
C88 VDD2.n68 B 0.013555f
C89 VDD2.n69 B 0.032038f
C90 VDD2.n70 B 0.014352f
C91 VDD2.n71 B 0.025225f
C92 VDD2.n72 B 0.013555f
C93 VDD2.n73 B 0.024029f
C94 VDD2.n74 B 0.022648f
C95 VDD2.t8 B 0.053843f
C96 VDD2.n75 B 0.162695f
C97 VDD2.n76 B 1.05038f
C98 VDD2.n77 B 0.013555f
C99 VDD2.n78 B 0.014352f
C100 VDD2.n79 B 0.032038f
C101 VDD2.n80 B 0.032038f
C102 VDD2.n81 B 0.014352f
C103 VDD2.n82 B 0.013555f
C104 VDD2.n83 B 0.025225f
C105 VDD2.n84 B 0.025225f
C106 VDD2.n85 B 0.013555f
C107 VDD2.n86 B 0.014352f
C108 VDD2.n87 B 0.032038f
C109 VDD2.n88 B 0.032038f
C110 VDD2.n89 B 0.014352f
C111 VDD2.n90 B 0.013555f
C112 VDD2.n91 B 0.025225f
C113 VDD2.n92 B 0.025225f
C114 VDD2.n93 B 0.013555f
C115 VDD2.n94 B 0.014352f
C116 VDD2.n95 B 0.032038f
C117 VDD2.n96 B 0.032038f
C118 VDD2.n97 B 0.032038f
C119 VDD2.n98 B 0.013953f
C120 VDD2.n99 B 0.013555f
C121 VDD2.n100 B 0.025225f
C122 VDD2.n101 B 0.025225f
C123 VDD2.n102 B 0.013555f
C124 VDD2.n103 B 0.014352f
C125 VDD2.n104 B 0.032038f
C126 VDD2.n105 B 0.067551f
C127 VDD2.n106 B 0.014352f
C128 VDD2.n107 B 0.013555f
C129 VDD2.n108 B 0.060373f
C130 VDD2.n109 B 0.055076f
C131 VDD2.n110 B 3.13374f
C132 VDD2.t6 B 0.19973f
C133 VDD2.t5 B 0.19973f
C134 VDD2.n111 B 1.7599f
C135 VDD2.n112 B 0.548434f
C136 VDD2.t2 B 0.19973f
C137 VDD2.t4 B 0.19973f
C138 VDD2.n113 B 1.78515f
C139 VN.t9 B 1.73776f
C140 VN.n0 B 0.687683f
C141 VN.n1 B 0.018083f
C142 VN.n2 B 0.023535f
C143 VN.n3 B 0.018083f
C144 VN.n4 B 0.021283f
C145 VN.n5 B 0.018083f
C146 VN.n6 B 0.015603f
C147 VN.n7 B 0.018083f
C148 VN.t6 B 1.73776f
C149 VN.n8 B 0.632718f
C150 VN.n9 B 0.018083f
C151 VN.n10 B 0.015603f
C152 VN.n11 B 0.018083f
C153 VN.t2 B 1.73776f
C154 VN.n12 B 0.682164f
C155 VN.t8 B 1.98662f
C156 VN.n13 B 0.642494f
C157 VN.n14 B 0.223533f
C158 VN.n15 B 0.029229f
C159 VN.n16 B 0.033533f
C160 VN.n17 B 0.03634f
C161 VN.n18 B 0.018083f
C162 VN.n19 B 0.018083f
C163 VN.n20 B 0.018083f
C164 VN.n21 B 0.034163f
C165 VN.n22 B 0.033533f
C166 VN.n23 B 0.033533f
C167 VN.n24 B 0.018083f
C168 VN.n25 B 0.018083f
C169 VN.n26 B 0.018083f
C170 VN.n27 B 0.033533f
C171 VN.n28 B 0.033533f
C172 VN.n29 B 0.034163f
C173 VN.n30 B 0.018083f
C174 VN.n31 B 0.018083f
C175 VN.n32 B 0.018083f
C176 VN.n33 B 0.03634f
C177 VN.n34 B 0.033533f
C178 VN.t0 B 1.73776f
C179 VN.n35 B 0.61574f
C180 VN.n36 B 0.029229f
C181 VN.n37 B 0.018083f
C182 VN.n38 B 0.018083f
C183 VN.n39 B 0.018083f
C184 VN.n40 B 0.033533f
C185 VN.n41 B 0.033533f
C186 VN.n42 B 0.029038f
C187 VN.n43 B 0.018083f
C188 VN.n44 B 0.018083f
C189 VN.n45 B 0.018083f
C190 VN.n46 B 0.033533f
C191 VN.n47 B 0.033533f
C192 VN.n48 B 0.024925f
C193 VN.n49 B 0.029181f
C194 VN.n50 B 0.047676f
C195 VN.t1 B 1.73776f
C196 VN.n51 B 0.687683f
C197 VN.n52 B 0.018083f
C198 VN.n53 B 0.023535f
C199 VN.n54 B 0.018083f
C200 VN.n55 B 0.021283f
C201 VN.n56 B 0.018083f
C202 VN.t3 B 1.73776f
C203 VN.n57 B 0.61574f
C204 VN.n58 B 0.015603f
C205 VN.n59 B 0.018083f
C206 VN.t4 B 1.73776f
C207 VN.n60 B 0.632718f
C208 VN.n61 B 0.018083f
C209 VN.n62 B 0.015603f
C210 VN.n63 B 0.018083f
C211 VN.t7 B 1.73776f
C212 VN.n64 B 0.682164f
C213 VN.t5 B 1.98662f
C214 VN.n65 B 0.642494f
C215 VN.n66 B 0.223533f
C216 VN.n67 B 0.029229f
C217 VN.n68 B 0.033533f
C218 VN.n69 B 0.03634f
C219 VN.n70 B 0.018083f
C220 VN.n71 B 0.018083f
C221 VN.n72 B 0.018083f
C222 VN.n73 B 0.034163f
C223 VN.n74 B 0.033533f
C224 VN.n75 B 0.033533f
C225 VN.n76 B 0.018083f
C226 VN.n77 B 0.018083f
C227 VN.n78 B 0.018083f
C228 VN.n79 B 0.033533f
C229 VN.n80 B 0.033533f
C230 VN.n81 B 0.034163f
C231 VN.n82 B 0.018083f
C232 VN.n83 B 0.018083f
C233 VN.n84 B 0.018083f
C234 VN.n85 B 0.03634f
C235 VN.n86 B 0.033533f
C236 VN.n87 B 0.029229f
C237 VN.n88 B 0.018083f
C238 VN.n89 B 0.018083f
C239 VN.n90 B 0.018083f
C240 VN.n91 B 0.033533f
C241 VN.n92 B 0.033533f
C242 VN.n93 B 0.029038f
C243 VN.n94 B 0.018083f
C244 VN.n95 B 0.018083f
C245 VN.n96 B 0.018083f
C246 VN.n97 B 0.033533f
C247 VN.n98 B 0.033533f
C248 VN.n99 B 0.024925f
C249 VN.n100 B 0.029181f
C250 VN.n101 B 1.24295f
C251 VTAIL.t2 B 0.209476f
C252 VTAIL.t4 B 0.209476f
C253 VTAIL.n0 B 1.77154f
C254 VTAIL.n1 B 0.653517f
C255 VTAIL.n2 B 0.036114f
C256 VTAIL.n3 B 0.026455f
C257 VTAIL.n4 B 0.014216f
C258 VTAIL.n5 B 0.033601f
C259 VTAIL.n6 B 0.015052f
C260 VTAIL.n7 B 0.026455f
C261 VTAIL.n8 B 0.014634f
C262 VTAIL.n9 B 0.033601f
C263 VTAIL.n10 B 0.015052f
C264 VTAIL.n11 B 0.026455f
C265 VTAIL.n12 B 0.014216f
C266 VTAIL.n13 B 0.033601f
C267 VTAIL.n14 B 0.015052f
C268 VTAIL.n15 B 0.026455f
C269 VTAIL.n16 B 0.014216f
C270 VTAIL.n17 B 0.025201f
C271 VTAIL.n18 B 0.023754f
C272 VTAIL.t13 B 0.05647f
C273 VTAIL.n19 B 0.170633f
C274 VTAIL.n20 B 1.10163f
C275 VTAIL.n21 B 0.014216f
C276 VTAIL.n22 B 0.015052f
C277 VTAIL.n23 B 0.033601f
C278 VTAIL.n24 B 0.033601f
C279 VTAIL.n25 B 0.015052f
C280 VTAIL.n26 B 0.014216f
C281 VTAIL.n27 B 0.026455f
C282 VTAIL.n28 B 0.026455f
C283 VTAIL.n29 B 0.014216f
C284 VTAIL.n30 B 0.015052f
C285 VTAIL.n31 B 0.033601f
C286 VTAIL.n32 B 0.033601f
C287 VTAIL.n33 B 0.015052f
C288 VTAIL.n34 B 0.014216f
C289 VTAIL.n35 B 0.026455f
C290 VTAIL.n36 B 0.026455f
C291 VTAIL.n37 B 0.014216f
C292 VTAIL.n38 B 0.014216f
C293 VTAIL.n39 B 0.015052f
C294 VTAIL.n40 B 0.033601f
C295 VTAIL.n41 B 0.033601f
C296 VTAIL.n42 B 0.033601f
C297 VTAIL.n43 B 0.014634f
C298 VTAIL.n44 B 0.014216f
C299 VTAIL.n45 B 0.026455f
C300 VTAIL.n46 B 0.026455f
C301 VTAIL.n47 B 0.014216f
C302 VTAIL.n48 B 0.015052f
C303 VTAIL.n49 B 0.033601f
C304 VTAIL.n50 B 0.070847f
C305 VTAIL.n51 B 0.015052f
C306 VTAIL.n52 B 0.014216f
C307 VTAIL.n53 B 0.063319f
C308 VTAIL.n54 B 0.039513f
C309 VTAIL.n55 B 0.490463f
C310 VTAIL.t15 B 0.209476f
C311 VTAIL.t16 B 0.209476f
C312 VTAIL.n56 B 1.77154f
C313 VTAIL.n57 B 0.821803f
C314 VTAIL.t12 B 0.209476f
C315 VTAIL.t19 B 0.209476f
C316 VTAIL.n58 B 1.77154f
C317 VTAIL.n59 B 2.2019f
C318 VTAIL.t7 B 0.209476f
C319 VTAIL.t9 B 0.209476f
C320 VTAIL.n60 B 1.77156f
C321 VTAIL.n61 B 2.20189f
C322 VTAIL.t1 B 0.209476f
C323 VTAIL.t0 B 0.209476f
C324 VTAIL.n62 B 1.77156f
C325 VTAIL.n63 B 0.821792f
C326 VTAIL.n64 B 0.036114f
C327 VTAIL.n65 B 0.026455f
C328 VTAIL.n66 B 0.014216f
C329 VTAIL.n67 B 0.033601f
C330 VTAIL.n68 B 0.015052f
C331 VTAIL.n69 B 0.026455f
C332 VTAIL.n70 B 0.014634f
C333 VTAIL.n71 B 0.033601f
C334 VTAIL.n72 B 0.014216f
C335 VTAIL.n73 B 0.015052f
C336 VTAIL.n74 B 0.026455f
C337 VTAIL.n75 B 0.014216f
C338 VTAIL.n76 B 0.033601f
C339 VTAIL.n77 B 0.015052f
C340 VTAIL.n78 B 0.026455f
C341 VTAIL.n79 B 0.014216f
C342 VTAIL.n80 B 0.025201f
C343 VTAIL.n81 B 0.023754f
C344 VTAIL.t6 B 0.05647f
C345 VTAIL.n82 B 0.170633f
C346 VTAIL.n83 B 1.10163f
C347 VTAIL.n84 B 0.014216f
C348 VTAIL.n85 B 0.015052f
C349 VTAIL.n86 B 0.033601f
C350 VTAIL.n87 B 0.033601f
C351 VTAIL.n88 B 0.015052f
C352 VTAIL.n89 B 0.014216f
C353 VTAIL.n90 B 0.026455f
C354 VTAIL.n91 B 0.026455f
C355 VTAIL.n92 B 0.014216f
C356 VTAIL.n93 B 0.015052f
C357 VTAIL.n94 B 0.033601f
C358 VTAIL.n95 B 0.033601f
C359 VTAIL.n96 B 0.015052f
C360 VTAIL.n97 B 0.014216f
C361 VTAIL.n98 B 0.026455f
C362 VTAIL.n99 B 0.026455f
C363 VTAIL.n100 B 0.014216f
C364 VTAIL.n101 B 0.015052f
C365 VTAIL.n102 B 0.033601f
C366 VTAIL.n103 B 0.033601f
C367 VTAIL.n104 B 0.033601f
C368 VTAIL.n105 B 0.014634f
C369 VTAIL.n106 B 0.014216f
C370 VTAIL.n107 B 0.026455f
C371 VTAIL.n108 B 0.026455f
C372 VTAIL.n109 B 0.014216f
C373 VTAIL.n110 B 0.015052f
C374 VTAIL.n111 B 0.033601f
C375 VTAIL.n112 B 0.070847f
C376 VTAIL.n113 B 0.015052f
C377 VTAIL.n114 B 0.014216f
C378 VTAIL.n115 B 0.063319f
C379 VTAIL.n116 B 0.039513f
C380 VTAIL.n117 B 0.490463f
C381 VTAIL.t10 B 0.209476f
C382 VTAIL.t11 B 0.209476f
C383 VTAIL.n118 B 1.77156f
C384 VTAIL.n119 B 0.719645f
C385 VTAIL.t14 B 0.209476f
C386 VTAIL.t18 B 0.209476f
C387 VTAIL.n120 B 1.77156f
C388 VTAIL.n121 B 0.821792f
C389 VTAIL.n122 B 0.036114f
C390 VTAIL.n123 B 0.026455f
C391 VTAIL.n124 B 0.014216f
C392 VTAIL.n125 B 0.033601f
C393 VTAIL.n126 B 0.015052f
C394 VTAIL.n127 B 0.026455f
C395 VTAIL.n128 B 0.014634f
C396 VTAIL.n129 B 0.033601f
C397 VTAIL.n130 B 0.014216f
C398 VTAIL.n131 B 0.015052f
C399 VTAIL.n132 B 0.026455f
C400 VTAIL.n133 B 0.014216f
C401 VTAIL.n134 B 0.033601f
C402 VTAIL.n135 B 0.015052f
C403 VTAIL.n136 B 0.026455f
C404 VTAIL.n137 B 0.014216f
C405 VTAIL.n138 B 0.025201f
C406 VTAIL.n139 B 0.023754f
C407 VTAIL.t17 B 0.05647f
C408 VTAIL.n140 B 0.170633f
C409 VTAIL.n141 B 1.10163f
C410 VTAIL.n142 B 0.014216f
C411 VTAIL.n143 B 0.015052f
C412 VTAIL.n144 B 0.033601f
C413 VTAIL.n145 B 0.033601f
C414 VTAIL.n146 B 0.015052f
C415 VTAIL.n147 B 0.014216f
C416 VTAIL.n148 B 0.026455f
C417 VTAIL.n149 B 0.026455f
C418 VTAIL.n150 B 0.014216f
C419 VTAIL.n151 B 0.015052f
C420 VTAIL.n152 B 0.033601f
C421 VTAIL.n153 B 0.033601f
C422 VTAIL.n154 B 0.015052f
C423 VTAIL.n155 B 0.014216f
C424 VTAIL.n156 B 0.026455f
C425 VTAIL.n157 B 0.026455f
C426 VTAIL.n158 B 0.014216f
C427 VTAIL.n159 B 0.015052f
C428 VTAIL.n160 B 0.033601f
C429 VTAIL.n161 B 0.033601f
C430 VTAIL.n162 B 0.033601f
C431 VTAIL.n163 B 0.014634f
C432 VTAIL.n164 B 0.014216f
C433 VTAIL.n165 B 0.026455f
C434 VTAIL.n166 B 0.026455f
C435 VTAIL.n167 B 0.014216f
C436 VTAIL.n168 B 0.015052f
C437 VTAIL.n169 B 0.033601f
C438 VTAIL.n170 B 0.070847f
C439 VTAIL.n171 B 0.015052f
C440 VTAIL.n172 B 0.014216f
C441 VTAIL.n173 B 0.063319f
C442 VTAIL.n174 B 0.039513f
C443 VTAIL.n175 B 1.68832f
C444 VTAIL.n176 B 0.036114f
C445 VTAIL.n177 B 0.026455f
C446 VTAIL.n178 B 0.014216f
C447 VTAIL.n179 B 0.033601f
C448 VTAIL.n180 B 0.015052f
C449 VTAIL.n181 B 0.026455f
C450 VTAIL.n182 B 0.014634f
C451 VTAIL.n183 B 0.033601f
C452 VTAIL.n184 B 0.015052f
C453 VTAIL.n185 B 0.026455f
C454 VTAIL.n186 B 0.014216f
C455 VTAIL.n187 B 0.033601f
C456 VTAIL.n188 B 0.015052f
C457 VTAIL.n189 B 0.026455f
C458 VTAIL.n190 B 0.014216f
C459 VTAIL.n191 B 0.025201f
C460 VTAIL.n192 B 0.023754f
C461 VTAIL.t8 B 0.05647f
C462 VTAIL.n193 B 0.170633f
C463 VTAIL.n194 B 1.10163f
C464 VTAIL.n195 B 0.014216f
C465 VTAIL.n196 B 0.015052f
C466 VTAIL.n197 B 0.033601f
C467 VTAIL.n198 B 0.033601f
C468 VTAIL.n199 B 0.015052f
C469 VTAIL.n200 B 0.014216f
C470 VTAIL.n201 B 0.026455f
C471 VTAIL.n202 B 0.026455f
C472 VTAIL.n203 B 0.014216f
C473 VTAIL.n204 B 0.015052f
C474 VTAIL.n205 B 0.033601f
C475 VTAIL.n206 B 0.033601f
C476 VTAIL.n207 B 0.015052f
C477 VTAIL.n208 B 0.014216f
C478 VTAIL.n209 B 0.026455f
C479 VTAIL.n210 B 0.026455f
C480 VTAIL.n211 B 0.014216f
C481 VTAIL.n212 B 0.014216f
C482 VTAIL.n213 B 0.015052f
C483 VTAIL.n214 B 0.033601f
C484 VTAIL.n215 B 0.033601f
C485 VTAIL.n216 B 0.033601f
C486 VTAIL.n217 B 0.014634f
C487 VTAIL.n218 B 0.014216f
C488 VTAIL.n219 B 0.026455f
C489 VTAIL.n220 B 0.026455f
C490 VTAIL.n221 B 0.014216f
C491 VTAIL.n222 B 0.015052f
C492 VTAIL.n223 B 0.033601f
C493 VTAIL.n224 B 0.070847f
C494 VTAIL.n225 B 0.015052f
C495 VTAIL.n226 B 0.014216f
C496 VTAIL.n227 B 0.063319f
C497 VTAIL.n228 B 0.039513f
C498 VTAIL.n229 B 1.68832f
C499 VTAIL.t5 B 0.209476f
C500 VTAIL.t3 B 0.209476f
C501 VTAIL.n230 B 1.77154f
C502 VTAIL.n231 B 0.603546f
C503 VDD1.n0 B 0.034904f
C504 VDD1.n1 B 0.025569f
C505 VDD1.n2 B 0.01374f
C506 VDD1.n3 B 0.032475f
C507 VDD1.n4 B 0.014548f
C508 VDD1.n5 B 0.025569f
C509 VDD1.n6 B 0.014144f
C510 VDD1.n7 B 0.032475f
C511 VDD1.n8 B 0.01374f
C512 VDD1.n9 B 0.014548f
C513 VDD1.n10 B 0.025569f
C514 VDD1.n11 B 0.01374f
C515 VDD1.n12 B 0.032475f
C516 VDD1.n13 B 0.014548f
C517 VDD1.n14 B 0.025569f
C518 VDD1.n15 B 0.01374f
C519 VDD1.n16 B 0.024356f
C520 VDD1.n17 B 0.022957f
C521 VDD1.t2 B 0.054578f
C522 VDD1.n18 B 0.164914f
C523 VDD1.n19 B 1.06471f
C524 VDD1.n20 B 0.01374f
C525 VDD1.n21 B 0.014548f
C526 VDD1.n22 B 0.032475f
C527 VDD1.n23 B 0.032475f
C528 VDD1.n24 B 0.014548f
C529 VDD1.n25 B 0.01374f
C530 VDD1.n26 B 0.025569f
C531 VDD1.n27 B 0.025569f
C532 VDD1.n28 B 0.01374f
C533 VDD1.n29 B 0.014548f
C534 VDD1.n30 B 0.032475f
C535 VDD1.n31 B 0.032475f
C536 VDD1.n32 B 0.014548f
C537 VDD1.n33 B 0.01374f
C538 VDD1.n34 B 0.025569f
C539 VDD1.n35 B 0.025569f
C540 VDD1.n36 B 0.01374f
C541 VDD1.n37 B 0.014548f
C542 VDD1.n38 B 0.032475f
C543 VDD1.n39 B 0.032475f
C544 VDD1.n40 B 0.032475f
C545 VDD1.n41 B 0.014144f
C546 VDD1.n42 B 0.01374f
C547 VDD1.n43 B 0.025569f
C548 VDD1.n44 B 0.025569f
C549 VDD1.n45 B 0.01374f
C550 VDD1.n46 B 0.014548f
C551 VDD1.n47 B 0.032475f
C552 VDD1.n48 B 0.068473f
C553 VDD1.n49 B 0.014548f
C554 VDD1.n50 B 0.01374f
C555 VDD1.n51 B 0.061196f
C556 VDD1.n52 B 0.076164f
C557 VDD1.t4 B 0.202455f
C558 VDD1.t3 B 0.202455f
C559 VDD1.n53 B 1.78391f
C560 VDD1.n54 B 0.860875f
C561 VDD1.n55 B 0.034904f
C562 VDD1.n56 B 0.025569f
C563 VDD1.n57 B 0.01374f
C564 VDD1.n58 B 0.032475f
C565 VDD1.n59 B 0.014548f
C566 VDD1.n60 B 0.025569f
C567 VDD1.n61 B 0.014144f
C568 VDD1.n62 B 0.032475f
C569 VDD1.n63 B 0.014548f
C570 VDD1.n64 B 0.025569f
C571 VDD1.n65 B 0.01374f
C572 VDD1.n66 B 0.032475f
C573 VDD1.n67 B 0.014548f
C574 VDD1.n68 B 0.025569f
C575 VDD1.n69 B 0.01374f
C576 VDD1.n70 B 0.024356f
C577 VDD1.n71 B 0.022957f
C578 VDD1.t5 B 0.054578f
C579 VDD1.n72 B 0.164914f
C580 VDD1.n73 B 1.06471f
C581 VDD1.n74 B 0.01374f
C582 VDD1.n75 B 0.014548f
C583 VDD1.n76 B 0.032475f
C584 VDD1.n77 B 0.032475f
C585 VDD1.n78 B 0.014548f
C586 VDD1.n79 B 0.01374f
C587 VDD1.n80 B 0.025569f
C588 VDD1.n81 B 0.025569f
C589 VDD1.n82 B 0.01374f
C590 VDD1.n83 B 0.014548f
C591 VDD1.n84 B 0.032475f
C592 VDD1.n85 B 0.032475f
C593 VDD1.n86 B 0.014548f
C594 VDD1.n87 B 0.01374f
C595 VDD1.n88 B 0.025569f
C596 VDD1.n89 B 0.025569f
C597 VDD1.n90 B 0.01374f
C598 VDD1.n91 B 0.01374f
C599 VDD1.n92 B 0.014548f
C600 VDD1.n93 B 0.032475f
C601 VDD1.n94 B 0.032475f
C602 VDD1.n95 B 0.032475f
C603 VDD1.n96 B 0.014144f
C604 VDD1.n97 B 0.01374f
C605 VDD1.n98 B 0.025569f
C606 VDD1.n99 B 0.025569f
C607 VDD1.n100 B 0.01374f
C608 VDD1.n101 B 0.014548f
C609 VDD1.n102 B 0.032475f
C610 VDD1.n103 B 0.068473f
C611 VDD1.n104 B 0.014548f
C612 VDD1.n105 B 0.01374f
C613 VDD1.n106 B 0.061196f
C614 VDD1.n107 B 0.076164f
C615 VDD1.t9 B 0.202455f
C616 VDD1.t0 B 0.202455f
C617 VDD1.n108 B 1.7839f
C618 VDD1.n109 B 0.852289f
C619 VDD1.t1 B 0.202455f
C620 VDD1.t8 B 0.202455f
C621 VDD1.n110 B 1.80955f
C622 VDD1.n111 B 3.49642f
C623 VDD1.t7 B 0.202455f
C624 VDD1.t6 B 0.202455f
C625 VDD1.n112 B 1.7839f
C626 VDD1.n113 B 3.48705f
C627 VP.t6 B 1.76873f
C628 VP.n0 B 0.699942f
C629 VP.n1 B 0.018405f
C630 VP.n2 B 0.023954f
C631 VP.n3 B 0.018405f
C632 VP.n4 B 0.021662f
C633 VP.n5 B 0.018405f
C634 VP.n6 B 0.015881f
C635 VP.n7 B 0.018405f
C636 VP.t4 B 1.76873f
C637 VP.n8 B 0.643997f
C638 VP.n9 B 0.018405f
C639 VP.n10 B 0.015881f
C640 VP.n11 B 0.018405f
C641 VP.t0 B 1.76873f
C642 VP.n12 B 0.626716f
C643 VP.n13 B 0.018405f
C644 VP.n14 B 0.029556f
C645 VP.n15 B 0.018405f
C646 VP.n16 B 0.025369f
C647 VP.t2 B 1.76873f
C648 VP.n17 B 0.699942f
C649 VP.n18 B 0.018405f
C650 VP.n19 B 0.023954f
C651 VP.n20 B 0.018405f
C652 VP.n21 B 0.021662f
C653 VP.n22 B 0.018405f
C654 VP.n23 B 0.015881f
C655 VP.n24 B 0.018405f
C656 VP.t5 B 1.76873f
C657 VP.n25 B 0.643997f
C658 VP.n26 B 0.018405f
C659 VP.n27 B 0.015881f
C660 VP.n28 B 0.018405f
C661 VP.t8 B 1.76873f
C662 VP.n29 B 0.694325f
C663 VP.t9 B 2.02203f
C664 VP.n30 B 0.653948f
C665 VP.n31 B 0.227518f
C666 VP.n32 B 0.02975f
C667 VP.n33 B 0.034131f
C668 VP.n34 B 0.036988f
C669 VP.n35 B 0.018405f
C670 VP.n36 B 0.018405f
C671 VP.n37 B 0.018405f
C672 VP.n38 B 0.034772f
C673 VP.n39 B 0.034131f
C674 VP.n40 B 0.034131f
C675 VP.n41 B 0.018405f
C676 VP.n42 B 0.018405f
C677 VP.n43 B 0.018405f
C678 VP.n44 B 0.034131f
C679 VP.n45 B 0.034131f
C680 VP.n46 B 0.034772f
C681 VP.n47 B 0.018405f
C682 VP.n48 B 0.018405f
C683 VP.n49 B 0.018405f
C684 VP.n50 B 0.036988f
C685 VP.n51 B 0.034131f
C686 VP.t1 B 1.76873f
C687 VP.n52 B 0.626716f
C688 VP.n53 B 0.02975f
C689 VP.n54 B 0.018405f
C690 VP.n55 B 0.018405f
C691 VP.n56 B 0.018405f
C692 VP.n57 B 0.034131f
C693 VP.n58 B 0.034131f
C694 VP.n59 B 0.029556f
C695 VP.n60 B 0.018405f
C696 VP.n61 B 0.018405f
C697 VP.n62 B 0.018405f
C698 VP.n63 B 0.034131f
C699 VP.n64 B 0.034131f
C700 VP.n65 B 0.025369f
C701 VP.n66 B 0.029701f
C702 VP.n67 B 1.2579f
C703 VP.t7 B 1.76873f
C704 VP.n68 B 0.699942f
C705 VP.n69 B 1.26957f
C706 VP.n70 B 0.029701f
C707 VP.n71 B 0.018405f
C708 VP.n72 B 0.034131f
C709 VP.n73 B 0.034131f
C710 VP.n74 B 0.023954f
C711 VP.n75 B 0.018405f
C712 VP.n76 B 0.018405f
C713 VP.n77 B 0.018405f
C714 VP.n78 B 0.034131f
C715 VP.n79 B 0.034131f
C716 VP.n80 B 0.021662f
C717 VP.n81 B 0.018405f
C718 VP.n82 B 0.018405f
C719 VP.n83 B 0.02975f
C720 VP.n84 B 0.034131f
C721 VP.n85 B 0.036988f
C722 VP.n86 B 0.018405f
C723 VP.n87 B 0.018405f
C724 VP.n88 B 0.018405f
C725 VP.n89 B 0.034772f
C726 VP.n90 B 0.034131f
C727 VP.n91 B 0.034131f
C728 VP.n92 B 0.018405f
C729 VP.n93 B 0.018405f
C730 VP.n94 B 0.018405f
C731 VP.n95 B 0.034131f
C732 VP.n96 B 0.034131f
C733 VP.n97 B 0.034772f
C734 VP.n98 B 0.018405f
C735 VP.n99 B 0.018405f
C736 VP.n100 B 0.018405f
C737 VP.n101 B 0.036988f
C738 VP.n102 B 0.034131f
C739 VP.t3 B 1.76873f
C740 VP.n103 B 0.626716f
C741 VP.n104 B 0.02975f
C742 VP.n105 B 0.018405f
C743 VP.n106 B 0.018405f
C744 VP.n107 B 0.018405f
C745 VP.n108 B 0.034131f
C746 VP.n109 B 0.034131f
C747 VP.n110 B 0.029556f
C748 VP.n111 B 0.018405f
C749 VP.n112 B 0.018405f
C750 VP.n113 B 0.018405f
C751 VP.n114 B 0.034131f
C752 VP.n115 B 0.034131f
C753 VP.n116 B 0.025369f
C754 VP.n117 B 0.029701f
C755 VP.n118 B 0.048526f
.ends

