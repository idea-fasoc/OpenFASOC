* NGSPICE file created from diff_pair_sample_1388.ext - technology: sky130A

.subckt diff_pair_sample_1388 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t1 VP.t0 VTAIL.t3 w_n1190_n4430# sky130_fd_pr__pfet_01v8 ad=6.7431 pd=35.36 as=6.7431 ps=35.36 w=17.29 l=0.22
X1 B.t11 B.t9 B.t10 w_n1190_n4430# sky130_fd_pr__pfet_01v8 ad=6.7431 pd=35.36 as=0 ps=0 w=17.29 l=0.22
X2 VDD2.t1 VN.t0 VTAIL.t1 w_n1190_n4430# sky130_fd_pr__pfet_01v8 ad=6.7431 pd=35.36 as=6.7431 ps=35.36 w=17.29 l=0.22
X3 VDD1.t0 VP.t1 VTAIL.t2 w_n1190_n4430# sky130_fd_pr__pfet_01v8 ad=6.7431 pd=35.36 as=6.7431 ps=35.36 w=17.29 l=0.22
X4 B.t8 B.t6 B.t7 w_n1190_n4430# sky130_fd_pr__pfet_01v8 ad=6.7431 pd=35.36 as=0 ps=0 w=17.29 l=0.22
X5 B.t5 B.t3 B.t4 w_n1190_n4430# sky130_fd_pr__pfet_01v8 ad=6.7431 pd=35.36 as=0 ps=0 w=17.29 l=0.22
X6 B.t2 B.t0 B.t1 w_n1190_n4430# sky130_fd_pr__pfet_01v8 ad=6.7431 pd=35.36 as=0 ps=0 w=17.29 l=0.22
X7 VDD2.t0 VN.t1 VTAIL.t0 w_n1190_n4430# sky130_fd_pr__pfet_01v8 ad=6.7431 pd=35.36 as=6.7431 ps=35.36 w=17.29 l=0.22
R0 VP.n0 VP.t1 2265.31
R1 VP.n0 VP.t0 2222.95
R2 VP VP.n0 0.0516364
R3 VTAIL.n1 VTAIL.t0 56.9245
R4 VTAIL.n3 VTAIL.t1 56.9244
R5 VTAIL.n0 VTAIL.t3 56.9244
R6 VTAIL.n2 VTAIL.t2 56.9244
R7 VTAIL.n1 VTAIL.n0 28.2376
R8 VTAIL.n3 VTAIL.n2 27.7634
R9 VTAIL.n2 VTAIL.n1 0.707397
R10 VTAIL VTAIL.n0 0.647052
R11 VTAIL VTAIL.n3 0.0608448
R12 VDD1 VDD1.t1 113.776
R13 VDD1 VDD1.t0 73.7799
R14 B.n120 B.t6 2124.91
R15 B.n270 B.t9 2124.91
R16 B.n44 B.t0 2124.91
R17 B.n36 B.t3 2124.91
R18 B.n359 B.n86 585
R19 B.n358 B.n357 585
R20 B.n356 B.n87 585
R21 B.n355 B.n354 585
R22 B.n353 B.n88 585
R23 B.n352 B.n351 585
R24 B.n350 B.n89 585
R25 B.n349 B.n348 585
R26 B.n347 B.n90 585
R27 B.n346 B.n345 585
R28 B.n344 B.n91 585
R29 B.n343 B.n342 585
R30 B.n341 B.n92 585
R31 B.n340 B.n339 585
R32 B.n338 B.n93 585
R33 B.n337 B.n336 585
R34 B.n335 B.n94 585
R35 B.n334 B.n333 585
R36 B.n332 B.n95 585
R37 B.n331 B.n330 585
R38 B.n329 B.n96 585
R39 B.n328 B.n327 585
R40 B.n326 B.n97 585
R41 B.n325 B.n324 585
R42 B.n323 B.n98 585
R43 B.n322 B.n321 585
R44 B.n320 B.n99 585
R45 B.n319 B.n318 585
R46 B.n317 B.n100 585
R47 B.n316 B.n315 585
R48 B.n314 B.n101 585
R49 B.n313 B.n312 585
R50 B.n311 B.n102 585
R51 B.n310 B.n309 585
R52 B.n308 B.n103 585
R53 B.n307 B.n306 585
R54 B.n305 B.n104 585
R55 B.n304 B.n303 585
R56 B.n302 B.n105 585
R57 B.n301 B.n300 585
R58 B.n299 B.n106 585
R59 B.n298 B.n297 585
R60 B.n296 B.n107 585
R61 B.n295 B.n294 585
R62 B.n293 B.n108 585
R63 B.n292 B.n291 585
R64 B.n290 B.n109 585
R65 B.n289 B.n288 585
R66 B.n287 B.n110 585
R67 B.n286 B.n285 585
R68 B.n284 B.n111 585
R69 B.n283 B.n282 585
R70 B.n281 B.n112 585
R71 B.n280 B.n279 585
R72 B.n278 B.n113 585
R73 B.n277 B.n276 585
R74 B.n275 B.n114 585
R75 B.n274 B.n273 585
R76 B.n269 B.n115 585
R77 B.n268 B.n267 585
R78 B.n266 B.n116 585
R79 B.n265 B.n264 585
R80 B.n263 B.n117 585
R81 B.n262 B.n261 585
R82 B.n260 B.n118 585
R83 B.n259 B.n258 585
R84 B.n257 B.n119 585
R85 B.n255 B.n254 585
R86 B.n253 B.n122 585
R87 B.n252 B.n251 585
R88 B.n250 B.n123 585
R89 B.n249 B.n248 585
R90 B.n247 B.n124 585
R91 B.n246 B.n245 585
R92 B.n244 B.n125 585
R93 B.n243 B.n242 585
R94 B.n241 B.n126 585
R95 B.n240 B.n239 585
R96 B.n238 B.n127 585
R97 B.n237 B.n236 585
R98 B.n235 B.n128 585
R99 B.n234 B.n233 585
R100 B.n232 B.n129 585
R101 B.n231 B.n230 585
R102 B.n229 B.n130 585
R103 B.n228 B.n227 585
R104 B.n226 B.n131 585
R105 B.n225 B.n224 585
R106 B.n223 B.n132 585
R107 B.n222 B.n221 585
R108 B.n220 B.n133 585
R109 B.n219 B.n218 585
R110 B.n217 B.n134 585
R111 B.n216 B.n215 585
R112 B.n214 B.n135 585
R113 B.n213 B.n212 585
R114 B.n211 B.n136 585
R115 B.n210 B.n209 585
R116 B.n208 B.n137 585
R117 B.n207 B.n206 585
R118 B.n205 B.n138 585
R119 B.n204 B.n203 585
R120 B.n202 B.n139 585
R121 B.n201 B.n200 585
R122 B.n199 B.n140 585
R123 B.n198 B.n197 585
R124 B.n196 B.n141 585
R125 B.n195 B.n194 585
R126 B.n193 B.n142 585
R127 B.n192 B.n191 585
R128 B.n190 B.n143 585
R129 B.n189 B.n188 585
R130 B.n187 B.n144 585
R131 B.n186 B.n185 585
R132 B.n184 B.n145 585
R133 B.n183 B.n182 585
R134 B.n181 B.n146 585
R135 B.n180 B.n179 585
R136 B.n178 B.n147 585
R137 B.n177 B.n176 585
R138 B.n175 B.n148 585
R139 B.n174 B.n173 585
R140 B.n172 B.n149 585
R141 B.n171 B.n170 585
R142 B.n361 B.n360 585
R143 B.n362 B.n85 585
R144 B.n364 B.n363 585
R145 B.n365 B.n84 585
R146 B.n367 B.n366 585
R147 B.n368 B.n83 585
R148 B.n370 B.n369 585
R149 B.n371 B.n82 585
R150 B.n373 B.n372 585
R151 B.n374 B.n81 585
R152 B.n376 B.n375 585
R153 B.n377 B.n80 585
R154 B.n379 B.n378 585
R155 B.n380 B.n79 585
R156 B.n382 B.n381 585
R157 B.n383 B.n78 585
R158 B.n385 B.n384 585
R159 B.n386 B.n77 585
R160 B.n388 B.n387 585
R161 B.n389 B.n76 585
R162 B.n391 B.n390 585
R163 B.n392 B.n75 585
R164 B.n394 B.n393 585
R165 B.n395 B.n74 585
R166 B.n583 B.n582 585
R167 B.n581 B.n8 585
R168 B.n580 B.n579 585
R169 B.n578 B.n9 585
R170 B.n577 B.n576 585
R171 B.n575 B.n10 585
R172 B.n574 B.n573 585
R173 B.n572 B.n11 585
R174 B.n571 B.n570 585
R175 B.n569 B.n12 585
R176 B.n568 B.n567 585
R177 B.n566 B.n13 585
R178 B.n565 B.n564 585
R179 B.n563 B.n14 585
R180 B.n562 B.n561 585
R181 B.n560 B.n15 585
R182 B.n559 B.n558 585
R183 B.n557 B.n16 585
R184 B.n556 B.n555 585
R185 B.n554 B.n17 585
R186 B.n553 B.n552 585
R187 B.n551 B.n18 585
R188 B.n550 B.n549 585
R189 B.n548 B.n19 585
R190 B.n547 B.n546 585
R191 B.n545 B.n20 585
R192 B.n544 B.n543 585
R193 B.n542 B.n21 585
R194 B.n541 B.n540 585
R195 B.n539 B.n22 585
R196 B.n538 B.n537 585
R197 B.n536 B.n23 585
R198 B.n535 B.n534 585
R199 B.n533 B.n24 585
R200 B.n532 B.n531 585
R201 B.n530 B.n25 585
R202 B.n529 B.n528 585
R203 B.n527 B.n26 585
R204 B.n526 B.n525 585
R205 B.n524 B.n27 585
R206 B.n523 B.n522 585
R207 B.n521 B.n28 585
R208 B.n520 B.n519 585
R209 B.n518 B.n29 585
R210 B.n517 B.n516 585
R211 B.n515 B.n30 585
R212 B.n514 B.n513 585
R213 B.n512 B.n31 585
R214 B.n511 B.n510 585
R215 B.n509 B.n32 585
R216 B.n508 B.n507 585
R217 B.n506 B.n33 585
R218 B.n505 B.n504 585
R219 B.n503 B.n34 585
R220 B.n502 B.n501 585
R221 B.n500 B.n35 585
R222 B.n499 B.n498 585
R223 B.n497 B.n496 585
R224 B.n495 B.n39 585
R225 B.n494 B.n493 585
R226 B.n492 B.n40 585
R227 B.n491 B.n490 585
R228 B.n489 B.n41 585
R229 B.n488 B.n487 585
R230 B.n486 B.n42 585
R231 B.n485 B.n484 585
R232 B.n483 B.n43 585
R233 B.n481 B.n480 585
R234 B.n479 B.n46 585
R235 B.n478 B.n477 585
R236 B.n476 B.n47 585
R237 B.n475 B.n474 585
R238 B.n473 B.n48 585
R239 B.n472 B.n471 585
R240 B.n470 B.n49 585
R241 B.n469 B.n468 585
R242 B.n467 B.n50 585
R243 B.n466 B.n465 585
R244 B.n464 B.n51 585
R245 B.n463 B.n462 585
R246 B.n461 B.n52 585
R247 B.n460 B.n459 585
R248 B.n458 B.n53 585
R249 B.n457 B.n456 585
R250 B.n455 B.n54 585
R251 B.n454 B.n453 585
R252 B.n452 B.n55 585
R253 B.n451 B.n450 585
R254 B.n449 B.n56 585
R255 B.n448 B.n447 585
R256 B.n446 B.n57 585
R257 B.n445 B.n444 585
R258 B.n443 B.n58 585
R259 B.n442 B.n441 585
R260 B.n440 B.n59 585
R261 B.n439 B.n438 585
R262 B.n437 B.n60 585
R263 B.n436 B.n435 585
R264 B.n434 B.n61 585
R265 B.n433 B.n432 585
R266 B.n431 B.n62 585
R267 B.n430 B.n429 585
R268 B.n428 B.n63 585
R269 B.n427 B.n426 585
R270 B.n425 B.n64 585
R271 B.n424 B.n423 585
R272 B.n422 B.n65 585
R273 B.n421 B.n420 585
R274 B.n419 B.n66 585
R275 B.n418 B.n417 585
R276 B.n416 B.n67 585
R277 B.n415 B.n414 585
R278 B.n413 B.n68 585
R279 B.n412 B.n411 585
R280 B.n410 B.n69 585
R281 B.n409 B.n408 585
R282 B.n407 B.n70 585
R283 B.n406 B.n405 585
R284 B.n404 B.n71 585
R285 B.n403 B.n402 585
R286 B.n401 B.n72 585
R287 B.n400 B.n399 585
R288 B.n398 B.n73 585
R289 B.n397 B.n396 585
R290 B.n584 B.n7 585
R291 B.n586 B.n585 585
R292 B.n587 B.n6 585
R293 B.n589 B.n588 585
R294 B.n590 B.n5 585
R295 B.n592 B.n591 585
R296 B.n593 B.n4 585
R297 B.n595 B.n594 585
R298 B.n596 B.n3 585
R299 B.n598 B.n597 585
R300 B.n599 B.n0 585
R301 B.n2 B.n1 585
R302 B.n156 B.n155 585
R303 B.n157 B.n154 585
R304 B.n159 B.n158 585
R305 B.n160 B.n153 585
R306 B.n162 B.n161 585
R307 B.n163 B.n152 585
R308 B.n165 B.n164 585
R309 B.n166 B.n151 585
R310 B.n168 B.n167 585
R311 B.n169 B.n150 585
R312 B.n170 B.n169 478.086
R313 B.n360 B.n359 478.086
R314 B.n396 B.n395 478.086
R315 B.n582 B.n7 478.086
R316 B.n601 B.n600 256.663
R317 B.n600 B.n599 235.042
R318 B.n600 B.n2 235.042
R319 B.n170 B.n149 163.367
R320 B.n174 B.n149 163.367
R321 B.n175 B.n174 163.367
R322 B.n176 B.n175 163.367
R323 B.n176 B.n147 163.367
R324 B.n180 B.n147 163.367
R325 B.n181 B.n180 163.367
R326 B.n182 B.n181 163.367
R327 B.n182 B.n145 163.367
R328 B.n186 B.n145 163.367
R329 B.n187 B.n186 163.367
R330 B.n188 B.n187 163.367
R331 B.n188 B.n143 163.367
R332 B.n192 B.n143 163.367
R333 B.n193 B.n192 163.367
R334 B.n194 B.n193 163.367
R335 B.n194 B.n141 163.367
R336 B.n198 B.n141 163.367
R337 B.n199 B.n198 163.367
R338 B.n200 B.n199 163.367
R339 B.n200 B.n139 163.367
R340 B.n204 B.n139 163.367
R341 B.n205 B.n204 163.367
R342 B.n206 B.n205 163.367
R343 B.n206 B.n137 163.367
R344 B.n210 B.n137 163.367
R345 B.n211 B.n210 163.367
R346 B.n212 B.n211 163.367
R347 B.n212 B.n135 163.367
R348 B.n216 B.n135 163.367
R349 B.n217 B.n216 163.367
R350 B.n218 B.n217 163.367
R351 B.n218 B.n133 163.367
R352 B.n222 B.n133 163.367
R353 B.n223 B.n222 163.367
R354 B.n224 B.n223 163.367
R355 B.n224 B.n131 163.367
R356 B.n228 B.n131 163.367
R357 B.n229 B.n228 163.367
R358 B.n230 B.n229 163.367
R359 B.n230 B.n129 163.367
R360 B.n234 B.n129 163.367
R361 B.n235 B.n234 163.367
R362 B.n236 B.n235 163.367
R363 B.n236 B.n127 163.367
R364 B.n240 B.n127 163.367
R365 B.n241 B.n240 163.367
R366 B.n242 B.n241 163.367
R367 B.n242 B.n125 163.367
R368 B.n246 B.n125 163.367
R369 B.n247 B.n246 163.367
R370 B.n248 B.n247 163.367
R371 B.n248 B.n123 163.367
R372 B.n252 B.n123 163.367
R373 B.n253 B.n252 163.367
R374 B.n254 B.n253 163.367
R375 B.n254 B.n119 163.367
R376 B.n259 B.n119 163.367
R377 B.n260 B.n259 163.367
R378 B.n261 B.n260 163.367
R379 B.n261 B.n117 163.367
R380 B.n265 B.n117 163.367
R381 B.n266 B.n265 163.367
R382 B.n267 B.n266 163.367
R383 B.n267 B.n115 163.367
R384 B.n274 B.n115 163.367
R385 B.n275 B.n274 163.367
R386 B.n276 B.n275 163.367
R387 B.n276 B.n113 163.367
R388 B.n280 B.n113 163.367
R389 B.n281 B.n280 163.367
R390 B.n282 B.n281 163.367
R391 B.n282 B.n111 163.367
R392 B.n286 B.n111 163.367
R393 B.n287 B.n286 163.367
R394 B.n288 B.n287 163.367
R395 B.n288 B.n109 163.367
R396 B.n292 B.n109 163.367
R397 B.n293 B.n292 163.367
R398 B.n294 B.n293 163.367
R399 B.n294 B.n107 163.367
R400 B.n298 B.n107 163.367
R401 B.n299 B.n298 163.367
R402 B.n300 B.n299 163.367
R403 B.n300 B.n105 163.367
R404 B.n304 B.n105 163.367
R405 B.n305 B.n304 163.367
R406 B.n306 B.n305 163.367
R407 B.n306 B.n103 163.367
R408 B.n310 B.n103 163.367
R409 B.n311 B.n310 163.367
R410 B.n312 B.n311 163.367
R411 B.n312 B.n101 163.367
R412 B.n316 B.n101 163.367
R413 B.n317 B.n316 163.367
R414 B.n318 B.n317 163.367
R415 B.n318 B.n99 163.367
R416 B.n322 B.n99 163.367
R417 B.n323 B.n322 163.367
R418 B.n324 B.n323 163.367
R419 B.n324 B.n97 163.367
R420 B.n328 B.n97 163.367
R421 B.n329 B.n328 163.367
R422 B.n330 B.n329 163.367
R423 B.n330 B.n95 163.367
R424 B.n334 B.n95 163.367
R425 B.n335 B.n334 163.367
R426 B.n336 B.n335 163.367
R427 B.n336 B.n93 163.367
R428 B.n340 B.n93 163.367
R429 B.n341 B.n340 163.367
R430 B.n342 B.n341 163.367
R431 B.n342 B.n91 163.367
R432 B.n346 B.n91 163.367
R433 B.n347 B.n346 163.367
R434 B.n348 B.n347 163.367
R435 B.n348 B.n89 163.367
R436 B.n352 B.n89 163.367
R437 B.n353 B.n352 163.367
R438 B.n354 B.n353 163.367
R439 B.n354 B.n87 163.367
R440 B.n358 B.n87 163.367
R441 B.n359 B.n358 163.367
R442 B.n395 B.n394 163.367
R443 B.n394 B.n75 163.367
R444 B.n390 B.n75 163.367
R445 B.n390 B.n389 163.367
R446 B.n389 B.n388 163.367
R447 B.n388 B.n77 163.367
R448 B.n384 B.n77 163.367
R449 B.n384 B.n383 163.367
R450 B.n383 B.n382 163.367
R451 B.n382 B.n79 163.367
R452 B.n378 B.n79 163.367
R453 B.n378 B.n377 163.367
R454 B.n377 B.n376 163.367
R455 B.n376 B.n81 163.367
R456 B.n372 B.n81 163.367
R457 B.n372 B.n371 163.367
R458 B.n371 B.n370 163.367
R459 B.n370 B.n83 163.367
R460 B.n366 B.n83 163.367
R461 B.n366 B.n365 163.367
R462 B.n365 B.n364 163.367
R463 B.n364 B.n85 163.367
R464 B.n360 B.n85 163.367
R465 B.n582 B.n581 163.367
R466 B.n581 B.n580 163.367
R467 B.n580 B.n9 163.367
R468 B.n576 B.n9 163.367
R469 B.n576 B.n575 163.367
R470 B.n575 B.n574 163.367
R471 B.n574 B.n11 163.367
R472 B.n570 B.n11 163.367
R473 B.n570 B.n569 163.367
R474 B.n569 B.n568 163.367
R475 B.n568 B.n13 163.367
R476 B.n564 B.n13 163.367
R477 B.n564 B.n563 163.367
R478 B.n563 B.n562 163.367
R479 B.n562 B.n15 163.367
R480 B.n558 B.n15 163.367
R481 B.n558 B.n557 163.367
R482 B.n557 B.n556 163.367
R483 B.n556 B.n17 163.367
R484 B.n552 B.n17 163.367
R485 B.n552 B.n551 163.367
R486 B.n551 B.n550 163.367
R487 B.n550 B.n19 163.367
R488 B.n546 B.n19 163.367
R489 B.n546 B.n545 163.367
R490 B.n545 B.n544 163.367
R491 B.n544 B.n21 163.367
R492 B.n540 B.n21 163.367
R493 B.n540 B.n539 163.367
R494 B.n539 B.n538 163.367
R495 B.n538 B.n23 163.367
R496 B.n534 B.n23 163.367
R497 B.n534 B.n533 163.367
R498 B.n533 B.n532 163.367
R499 B.n532 B.n25 163.367
R500 B.n528 B.n25 163.367
R501 B.n528 B.n527 163.367
R502 B.n527 B.n526 163.367
R503 B.n526 B.n27 163.367
R504 B.n522 B.n27 163.367
R505 B.n522 B.n521 163.367
R506 B.n521 B.n520 163.367
R507 B.n520 B.n29 163.367
R508 B.n516 B.n29 163.367
R509 B.n516 B.n515 163.367
R510 B.n515 B.n514 163.367
R511 B.n514 B.n31 163.367
R512 B.n510 B.n31 163.367
R513 B.n510 B.n509 163.367
R514 B.n509 B.n508 163.367
R515 B.n508 B.n33 163.367
R516 B.n504 B.n33 163.367
R517 B.n504 B.n503 163.367
R518 B.n503 B.n502 163.367
R519 B.n502 B.n35 163.367
R520 B.n498 B.n35 163.367
R521 B.n498 B.n497 163.367
R522 B.n497 B.n39 163.367
R523 B.n493 B.n39 163.367
R524 B.n493 B.n492 163.367
R525 B.n492 B.n491 163.367
R526 B.n491 B.n41 163.367
R527 B.n487 B.n41 163.367
R528 B.n487 B.n486 163.367
R529 B.n486 B.n485 163.367
R530 B.n485 B.n43 163.367
R531 B.n480 B.n43 163.367
R532 B.n480 B.n479 163.367
R533 B.n479 B.n478 163.367
R534 B.n478 B.n47 163.367
R535 B.n474 B.n47 163.367
R536 B.n474 B.n473 163.367
R537 B.n473 B.n472 163.367
R538 B.n472 B.n49 163.367
R539 B.n468 B.n49 163.367
R540 B.n468 B.n467 163.367
R541 B.n467 B.n466 163.367
R542 B.n466 B.n51 163.367
R543 B.n462 B.n51 163.367
R544 B.n462 B.n461 163.367
R545 B.n461 B.n460 163.367
R546 B.n460 B.n53 163.367
R547 B.n456 B.n53 163.367
R548 B.n456 B.n455 163.367
R549 B.n455 B.n454 163.367
R550 B.n454 B.n55 163.367
R551 B.n450 B.n55 163.367
R552 B.n450 B.n449 163.367
R553 B.n449 B.n448 163.367
R554 B.n448 B.n57 163.367
R555 B.n444 B.n57 163.367
R556 B.n444 B.n443 163.367
R557 B.n443 B.n442 163.367
R558 B.n442 B.n59 163.367
R559 B.n438 B.n59 163.367
R560 B.n438 B.n437 163.367
R561 B.n437 B.n436 163.367
R562 B.n436 B.n61 163.367
R563 B.n432 B.n61 163.367
R564 B.n432 B.n431 163.367
R565 B.n431 B.n430 163.367
R566 B.n430 B.n63 163.367
R567 B.n426 B.n63 163.367
R568 B.n426 B.n425 163.367
R569 B.n425 B.n424 163.367
R570 B.n424 B.n65 163.367
R571 B.n420 B.n65 163.367
R572 B.n420 B.n419 163.367
R573 B.n419 B.n418 163.367
R574 B.n418 B.n67 163.367
R575 B.n414 B.n67 163.367
R576 B.n414 B.n413 163.367
R577 B.n413 B.n412 163.367
R578 B.n412 B.n69 163.367
R579 B.n408 B.n69 163.367
R580 B.n408 B.n407 163.367
R581 B.n407 B.n406 163.367
R582 B.n406 B.n71 163.367
R583 B.n402 B.n71 163.367
R584 B.n402 B.n401 163.367
R585 B.n401 B.n400 163.367
R586 B.n400 B.n73 163.367
R587 B.n396 B.n73 163.367
R588 B.n586 B.n7 163.367
R589 B.n587 B.n586 163.367
R590 B.n588 B.n587 163.367
R591 B.n588 B.n5 163.367
R592 B.n592 B.n5 163.367
R593 B.n593 B.n592 163.367
R594 B.n594 B.n593 163.367
R595 B.n594 B.n3 163.367
R596 B.n598 B.n3 163.367
R597 B.n599 B.n598 163.367
R598 B.n156 B.n2 163.367
R599 B.n157 B.n156 163.367
R600 B.n158 B.n157 163.367
R601 B.n158 B.n153 163.367
R602 B.n162 B.n153 163.367
R603 B.n163 B.n162 163.367
R604 B.n164 B.n163 163.367
R605 B.n164 B.n151 163.367
R606 B.n168 B.n151 163.367
R607 B.n169 B.n168 163.367
R608 B.n270 B.t10 122.567
R609 B.n44 B.t2 122.567
R610 B.n120 B.t7 122.546
R611 B.n36 B.t5 122.546
R612 B.n271 B.t11 111.901
R613 B.n45 B.t1 111.901
R614 B.n121 B.t8 111.879
R615 B.n37 B.t4 111.879
R616 B.n256 B.n121 59.5399
R617 B.n272 B.n271 59.5399
R618 B.n482 B.n45 59.5399
R619 B.n38 B.n37 59.5399
R620 B.n584 B.n583 31.0639
R621 B.n397 B.n74 31.0639
R622 B.n361 B.n86 31.0639
R623 B.n171 B.n150 31.0639
R624 B B.n601 18.0485
R625 B.n121 B.n120 10.6672
R626 B.n271 B.n270 10.6672
R627 B.n45 B.n44 10.6672
R628 B.n37 B.n36 10.6672
R629 B.n585 B.n584 10.6151
R630 B.n585 B.n6 10.6151
R631 B.n589 B.n6 10.6151
R632 B.n590 B.n589 10.6151
R633 B.n591 B.n590 10.6151
R634 B.n591 B.n4 10.6151
R635 B.n595 B.n4 10.6151
R636 B.n596 B.n595 10.6151
R637 B.n597 B.n596 10.6151
R638 B.n597 B.n0 10.6151
R639 B.n583 B.n8 10.6151
R640 B.n579 B.n8 10.6151
R641 B.n579 B.n578 10.6151
R642 B.n578 B.n577 10.6151
R643 B.n577 B.n10 10.6151
R644 B.n573 B.n10 10.6151
R645 B.n573 B.n572 10.6151
R646 B.n572 B.n571 10.6151
R647 B.n571 B.n12 10.6151
R648 B.n567 B.n12 10.6151
R649 B.n567 B.n566 10.6151
R650 B.n566 B.n565 10.6151
R651 B.n565 B.n14 10.6151
R652 B.n561 B.n14 10.6151
R653 B.n561 B.n560 10.6151
R654 B.n560 B.n559 10.6151
R655 B.n559 B.n16 10.6151
R656 B.n555 B.n16 10.6151
R657 B.n555 B.n554 10.6151
R658 B.n554 B.n553 10.6151
R659 B.n553 B.n18 10.6151
R660 B.n549 B.n18 10.6151
R661 B.n549 B.n548 10.6151
R662 B.n548 B.n547 10.6151
R663 B.n547 B.n20 10.6151
R664 B.n543 B.n20 10.6151
R665 B.n543 B.n542 10.6151
R666 B.n542 B.n541 10.6151
R667 B.n541 B.n22 10.6151
R668 B.n537 B.n22 10.6151
R669 B.n537 B.n536 10.6151
R670 B.n536 B.n535 10.6151
R671 B.n535 B.n24 10.6151
R672 B.n531 B.n24 10.6151
R673 B.n531 B.n530 10.6151
R674 B.n530 B.n529 10.6151
R675 B.n529 B.n26 10.6151
R676 B.n525 B.n26 10.6151
R677 B.n525 B.n524 10.6151
R678 B.n524 B.n523 10.6151
R679 B.n523 B.n28 10.6151
R680 B.n519 B.n28 10.6151
R681 B.n519 B.n518 10.6151
R682 B.n518 B.n517 10.6151
R683 B.n517 B.n30 10.6151
R684 B.n513 B.n30 10.6151
R685 B.n513 B.n512 10.6151
R686 B.n512 B.n511 10.6151
R687 B.n511 B.n32 10.6151
R688 B.n507 B.n32 10.6151
R689 B.n507 B.n506 10.6151
R690 B.n506 B.n505 10.6151
R691 B.n505 B.n34 10.6151
R692 B.n501 B.n34 10.6151
R693 B.n501 B.n500 10.6151
R694 B.n500 B.n499 10.6151
R695 B.n496 B.n495 10.6151
R696 B.n495 B.n494 10.6151
R697 B.n494 B.n40 10.6151
R698 B.n490 B.n40 10.6151
R699 B.n490 B.n489 10.6151
R700 B.n489 B.n488 10.6151
R701 B.n488 B.n42 10.6151
R702 B.n484 B.n42 10.6151
R703 B.n484 B.n483 10.6151
R704 B.n481 B.n46 10.6151
R705 B.n477 B.n46 10.6151
R706 B.n477 B.n476 10.6151
R707 B.n476 B.n475 10.6151
R708 B.n475 B.n48 10.6151
R709 B.n471 B.n48 10.6151
R710 B.n471 B.n470 10.6151
R711 B.n470 B.n469 10.6151
R712 B.n469 B.n50 10.6151
R713 B.n465 B.n50 10.6151
R714 B.n465 B.n464 10.6151
R715 B.n464 B.n463 10.6151
R716 B.n463 B.n52 10.6151
R717 B.n459 B.n52 10.6151
R718 B.n459 B.n458 10.6151
R719 B.n458 B.n457 10.6151
R720 B.n457 B.n54 10.6151
R721 B.n453 B.n54 10.6151
R722 B.n453 B.n452 10.6151
R723 B.n452 B.n451 10.6151
R724 B.n451 B.n56 10.6151
R725 B.n447 B.n56 10.6151
R726 B.n447 B.n446 10.6151
R727 B.n446 B.n445 10.6151
R728 B.n445 B.n58 10.6151
R729 B.n441 B.n58 10.6151
R730 B.n441 B.n440 10.6151
R731 B.n440 B.n439 10.6151
R732 B.n439 B.n60 10.6151
R733 B.n435 B.n60 10.6151
R734 B.n435 B.n434 10.6151
R735 B.n434 B.n433 10.6151
R736 B.n433 B.n62 10.6151
R737 B.n429 B.n62 10.6151
R738 B.n429 B.n428 10.6151
R739 B.n428 B.n427 10.6151
R740 B.n427 B.n64 10.6151
R741 B.n423 B.n64 10.6151
R742 B.n423 B.n422 10.6151
R743 B.n422 B.n421 10.6151
R744 B.n421 B.n66 10.6151
R745 B.n417 B.n66 10.6151
R746 B.n417 B.n416 10.6151
R747 B.n416 B.n415 10.6151
R748 B.n415 B.n68 10.6151
R749 B.n411 B.n68 10.6151
R750 B.n411 B.n410 10.6151
R751 B.n410 B.n409 10.6151
R752 B.n409 B.n70 10.6151
R753 B.n405 B.n70 10.6151
R754 B.n405 B.n404 10.6151
R755 B.n404 B.n403 10.6151
R756 B.n403 B.n72 10.6151
R757 B.n399 B.n72 10.6151
R758 B.n399 B.n398 10.6151
R759 B.n398 B.n397 10.6151
R760 B.n393 B.n74 10.6151
R761 B.n393 B.n392 10.6151
R762 B.n392 B.n391 10.6151
R763 B.n391 B.n76 10.6151
R764 B.n387 B.n76 10.6151
R765 B.n387 B.n386 10.6151
R766 B.n386 B.n385 10.6151
R767 B.n385 B.n78 10.6151
R768 B.n381 B.n78 10.6151
R769 B.n381 B.n380 10.6151
R770 B.n380 B.n379 10.6151
R771 B.n379 B.n80 10.6151
R772 B.n375 B.n80 10.6151
R773 B.n375 B.n374 10.6151
R774 B.n374 B.n373 10.6151
R775 B.n373 B.n82 10.6151
R776 B.n369 B.n82 10.6151
R777 B.n369 B.n368 10.6151
R778 B.n368 B.n367 10.6151
R779 B.n367 B.n84 10.6151
R780 B.n363 B.n84 10.6151
R781 B.n363 B.n362 10.6151
R782 B.n362 B.n361 10.6151
R783 B.n155 B.n1 10.6151
R784 B.n155 B.n154 10.6151
R785 B.n159 B.n154 10.6151
R786 B.n160 B.n159 10.6151
R787 B.n161 B.n160 10.6151
R788 B.n161 B.n152 10.6151
R789 B.n165 B.n152 10.6151
R790 B.n166 B.n165 10.6151
R791 B.n167 B.n166 10.6151
R792 B.n167 B.n150 10.6151
R793 B.n172 B.n171 10.6151
R794 B.n173 B.n172 10.6151
R795 B.n173 B.n148 10.6151
R796 B.n177 B.n148 10.6151
R797 B.n178 B.n177 10.6151
R798 B.n179 B.n178 10.6151
R799 B.n179 B.n146 10.6151
R800 B.n183 B.n146 10.6151
R801 B.n184 B.n183 10.6151
R802 B.n185 B.n184 10.6151
R803 B.n185 B.n144 10.6151
R804 B.n189 B.n144 10.6151
R805 B.n190 B.n189 10.6151
R806 B.n191 B.n190 10.6151
R807 B.n191 B.n142 10.6151
R808 B.n195 B.n142 10.6151
R809 B.n196 B.n195 10.6151
R810 B.n197 B.n196 10.6151
R811 B.n197 B.n140 10.6151
R812 B.n201 B.n140 10.6151
R813 B.n202 B.n201 10.6151
R814 B.n203 B.n202 10.6151
R815 B.n203 B.n138 10.6151
R816 B.n207 B.n138 10.6151
R817 B.n208 B.n207 10.6151
R818 B.n209 B.n208 10.6151
R819 B.n209 B.n136 10.6151
R820 B.n213 B.n136 10.6151
R821 B.n214 B.n213 10.6151
R822 B.n215 B.n214 10.6151
R823 B.n215 B.n134 10.6151
R824 B.n219 B.n134 10.6151
R825 B.n220 B.n219 10.6151
R826 B.n221 B.n220 10.6151
R827 B.n221 B.n132 10.6151
R828 B.n225 B.n132 10.6151
R829 B.n226 B.n225 10.6151
R830 B.n227 B.n226 10.6151
R831 B.n227 B.n130 10.6151
R832 B.n231 B.n130 10.6151
R833 B.n232 B.n231 10.6151
R834 B.n233 B.n232 10.6151
R835 B.n233 B.n128 10.6151
R836 B.n237 B.n128 10.6151
R837 B.n238 B.n237 10.6151
R838 B.n239 B.n238 10.6151
R839 B.n239 B.n126 10.6151
R840 B.n243 B.n126 10.6151
R841 B.n244 B.n243 10.6151
R842 B.n245 B.n244 10.6151
R843 B.n245 B.n124 10.6151
R844 B.n249 B.n124 10.6151
R845 B.n250 B.n249 10.6151
R846 B.n251 B.n250 10.6151
R847 B.n251 B.n122 10.6151
R848 B.n255 B.n122 10.6151
R849 B.n258 B.n257 10.6151
R850 B.n258 B.n118 10.6151
R851 B.n262 B.n118 10.6151
R852 B.n263 B.n262 10.6151
R853 B.n264 B.n263 10.6151
R854 B.n264 B.n116 10.6151
R855 B.n268 B.n116 10.6151
R856 B.n269 B.n268 10.6151
R857 B.n273 B.n269 10.6151
R858 B.n277 B.n114 10.6151
R859 B.n278 B.n277 10.6151
R860 B.n279 B.n278 10.6151
R861 B.n279 B.n112 10.6151
R862 B.n283 B.n112 10.6151
R863 B.n284 B.n283 10.6151
R864 B.n285 B.n284 10.6151
R865 B.n285 B.n110 10.6151
R866 B.n289 B.n110 10.6151
R867 B.n290 B.n289 10.6151
R868 B.n291 B.n290 10.6151
R869 B.n291 B.n108 10.6151
R870 B.n295 B.n108 10.6151
R871 B.n296 B.n295 10.6151
R872 B.n297 B.n296 10.6151
R873 B.n297 B.n106 10.6151
R874 B.n301 B.n106 10.6151
R875 B.n302 B.n301 10.6151
R876 B.n303 B.n302 10.6151
R877 B.n303 B.n104 10.6151
R878 B.n307 B.n104 10.6151
R879 B.n308 B.n307 10.6151
R880 B.n309 B.n308 10.6151
R881 B.n309 B.n102 10.6151
R882 B.n313 B.n102 10.6151
R883 B.n314 B.n313 10.6151
R884 B.n315 B.n314 10.6151
R885 B.n315 B.n100 10.6151
R886 B.n319 B.n100 10.6151
R887 B.n320 B.n319 10.6151
R888 B.n321 B.n320 10.6151
R889 B.n321 B.n98 10.6151
R890 B.n325 B.n98 10.6151
R891 B.n326 B.n325 10.6151
R892 B.n327 B.n326 10.6151
R893 B.n327 B.n96 10.6151
R894 B.n331 B.n96 10.6151
R895 B.n332 B.n331 10.6151
R896 B.n333 B.n332 10.6151
R897 B.n333 B.n94 10.6151
R898 B.n337 B.n94 10.6151
R899 B.n338 B.n337 10.6151
R900 B.n339 B.n338 10.6151
R901 B.n339 B.n92 10.6151
R902 B.n343 B.n92 10.6151
R903 B.n344 B.n343 10.6151
R904 B.n345 B.n344 10.6151
R905 B.n345 B.n90 10.6151
R906 B.n349 B.n90 10.6151
R907 B.n350 B.n349 10.6151
R908 B.n351 B.n350 10.6151
R909 B.n351 B.n88 10.6151
R910 B.n355 B.n88 10.6151
R911 B.n356 B.n355 10.6151
R912 B.n357 B.n356 10.6151
R913 B.n357 B.n86 10.6151
R914 B.n499 B.n38 8.74196
R915 B.n482 B.n481 8.74196
R916 B.n256 B.n255 8.74196
R917 B.n272 B.n114 8.74196
R918 B.n601 B.n0 8.11757
R919 B.n601 B.n1 8.11757
R920 B.n496 B.n38 1.87367
R921 B.n483 B.n482 1.87367
R922 B.n257 B.n256 1.87367
R923 B.n273 B.n272 1.87367
R924 VN VN.t1 2265.69
R925 VN VN.t0 2223
R926 VDD2.n0 VDD2.t1 113.133
R927 VDD2.n0 VDD2.t0 73.6032
R928 VDD2 VDD2.n0 0.177224
C0 B VTAIL 3.27292f
C1 VDD1 w_n1190_n4430# 1.92018f
C2 VDD1 VP 1.85571f
C3 w_n1190_n4430# VP 1.7333f
C4 VDD1 VN 0.148353f
C5 VDD2 VDD1 0.425142f
C6 w_n1190_n4430# VN 1.58685f
C7 VDD2 w_n1190_n4430# 1.92012f
C8 VN VP 5.3306f
C9 VDD2 VP 0.236096f
C10 B VDD1 1.69116f
C11 B w_n1190_n4430# 7.76918f
C12 B VP 0.937532f
C13 VDD2 VN 1.77544f
C14 VDD1 VTAIL 10.392799f
C15 B VN 0.706307f
C16 w_n1190_n4430# VTAIL 3.96176f
C17 B VDD2 1.7026f
C18 VTAIL VP 0.931162f
C19 VN VTAIL 0.91606f
C20 VDD2 VTAIL 10.4172f
C21 VDD2 VSUBS 0.893243f
C22 VDD1 VSUBS 4.570266f
C23 VTAIL VSUBS 0.210874f
C24 VN VSUBS 5.88097f
C25 VP VSUBS 1.172122f
C26 B VSUBS 2.593818f
C27 w_n1190_n4430# VSUBS 64.5028f
C28 VDD2.t1 VSUBS 3.73733f
C29 VDD2.t0 VSUBS 3.11012f
C30 VDD2.n0 VSUBS 3.52378f
C31 VN.t0 VSUBS 0.507075f
C32 VN.t1 VSUBS 0.547091f
C33 B.n0 VSUBS 0.006677f
C34 B.n1 VSUBS 0.006677f
C35 B.n2 VSUBS 0.009875f
C36 B.n3 VSUBS 0.007568f
C37 B.n4 VSUBS 0.007568f
C38 B.n5 VSUBS 0.007568f
C39 B.n6 VSUBS 0.007568f
C40 B.n7 VSUBS 0.016829f
C41 B.n8 VSUBS 0.007568f
C42 B.n9 VSUBS 0.007568f
C43 B.n10 VSUBS 0.007568f
C44 B.n11 VSUBS 0.007568f
C45 B.n12 VSUBS 0.007568f
C46 B.n13 VSUBS 0.007568f
C47 B.n14 VSUBS 0.007568f
C48 B.n15 VSUBS 0.007568f
C49 B.n16 VSUBS 0.007568f
C50 B.n17 VSUBS 0.007568f
C51 B.n18 VSUBS 0.007568f
C52 B.n19 VSUBS 0.007568f
C53 B.n20 VSUBS 0.007568f
C54 B.n21 VSUBS 0.007568f
C55 B.n22 VSUBS 0.007568f
C56 B.n23 VSUBS 0.007568f
C57 B.n24 VSUBS 0.007568f
C58 B.n25 VSUBS 0.007568f
C59 B.n26 VSUBS 0.007568f
C60 B.n27 VSUBS 0.007568f
C61 B.n28 VSUBS 0.007568f
C62 B.n29 VSUBS 0.007568f
C63 B.n30 VSUBS 0.007568f
C64 B.n31 VSUBS 0.007568f
C65 B.n32 VSUBS 0.007568f
C66 B.n33 VSUBS 0.007568f
C67 B.n34 VSUBS 0.007568f
C68 B.n35 VSUBS 0.007568f
C69 B.t4 VSUBS 0.629258f
C70 B.t5 VSUBS 0.634172f
C71 B.t3 VSUBS 0.158223f
C72 B.n36 VSUBS 0.110655f
C73 B.n37 VSUBS 0.067249f
C74 B.n38 VSUBS 0.017534f
C75 B.n39 VSUBS 0.007568f
C76 B.n40 VSUBS 0.007568f
C77 B.n41 VSUBS 0.007568f
C78 B.n42 VSUBS 0.007568f
C79 B.n43 VSUBS 0.007568f
C80 B.t1 VSUBS 0.629236f
C81 B.t2 VSUBS 0.634151f
C82 B.t0 VSUBS 0.158223f
C83 B.n44 VSUBS 0.110676f
C84 B.n45 VSUBS 0.06727f
C85 B.n46 VSUBS 0.007568f
C86 B.n47 VSUBS 0.007568f
C87 B.n48 VSUBS 0.007568f
C88 B.n49 VSUBS 0.007568f
C89 B.n50 VSUBS 0.007568f
C90 B.n51 VSUBS 0.007568f
C91 B.n52 VSUBS 0.007568f
C92 B.n53 VSUBS 0.007568f
C93 B.n54 VSUBS 0.007568f
C94 B.n55 VSUBS 0.007568f
C95 B.n56 VSUBS 0.007568f
C96 B.n57 VSUBS 0.007568f
C97 B.n58 VSUBS 0.007568f
C98 B.n59 VSUBS 0.007568f
C99 B.n60 VSUBS 0.007568f
C100 B.n61 VSUBS 0.007568f
C101 B.n62 VSUBS 0.007568f
C102 B.n63 VSUBS 0.007568f
C103 B.n64 VSUBS 0.007568f
C104 B.n65 VSUBS 0.007568f
C105 B.n66 VSUBS 0.007568f
C106 B.n67 VSUBS 0.007568f
C107 B.n68 VSUBS 0.007568f
C108 B.n69 VSUBS 0.007568f
C109 B.n70 VSUBS 0.007568f
C110 B.n71 VSUBS 0.007568f
C111 B.n72 VSUBS 0.007568f
C112 B.n73 VSUBS 0.007568f
C113 B.n74 VSUBS 0.016829f
C114 B.n75 VSUBS 0.007568f
C115 B.n76 VSUBS 0.007568f
C116 B.n77 VSUBS 0.007568f
C117 B.n78 VSUBS 0.007568f
C118 B.n79 VSUBS 0.007568f
C119 B.n80 VSUBS 0.007568f
C120 B.n81 VSUBS 0.007568f
C121 B.n82 VSUBS 0.007568f
C122 B.n83 VSUBS 0.007568f
C123 B.n84 VSUBS 0.007568f
C124 B.n85 VSUBS 0.007568f
C125 B.n86 VSUBS 0.016508f
C126 B.n87 VSUBS 0.007568f
C127 B.n88 VSUBS 0.007568f
C128 B.n89 VSUBS 0.007568f
C129 B.n90 VSUBS 0.007568f
C130 B.n91 VSUBS 0.007568f
C131 B.n92 VSUBS 0.007568f
C132 B.n93 VSUBS 0.007568f
C133 B.n94 VSUBS 0.007568f
C134 B.n95 VSUBS 0.007568f
C135 B.n96 VSUBS 0.007568f
C136 B.n97 VSUBS 0.007568f
C137 B.n98 VSUBS 0.007568f
C138 B.n99 VSUBS 0.007568f
C139 B.n100 VSUBS 0.007568f
C140 B.n101 VSUBS 0.007568f
C141 B.n102 VSUBS 0.007568f
C142 B.n103 VSUBS 0.007568f
C143 B.n104 VSUBS 0.007568f
C144 B.n105 VSUBS 0.007568f
C145 B.n106 VSUBS 0.007568f
C146 B.n107 VSUBS 0.007568f
C147 B.n108 VSUBS 0.007568f
C148 B.n109 VSUBS 0.007568f
C149 B.n110 VSUBS 0.007568f
C150 B.n111 VSUBS 0.007568f
C151 B.n112 VSUBS 0.007568f
C152 B.n113 VSUBS 0.007568f
C153 B.n114 VSUBS 0.0069f
C154 B.n115 VSUBS 0.007568f
C155 B.n116 VSUBS 0.007568f
C156 B.n117 VSUBS 0.007568f
C157 B.n118 VSUBS 0.007568f
C158 B.n119 VSUBS 0.007568f
C159 B.t8 VSUBS 0.629258f
C160 B.t7 VSUBS 0.634172f
C161 B.t6 VSUBS 0.158223f
C162 B.n120 VSUBS 0.110655f
C163 B.n121 VSUBS 0.067249f
C164 B.n122 VSUBS 0.007568f
C165 B.n123 VSUBS 0.007568f
C166 B.n124 VSUBS 0.007568f
C167 B.n125 VSUBS 0.007568f
C168 B.n126 VSUBS 0.007568f
C169 B.n127 VSUBS 0.007568f
C170 B.n128 VSUBS 0.007568f
C171 B.n129 VSUBS 0.007568f
C172 B.n130 VSUBS 0.007568f
C173 B.n131 VSUBS 0.007568f
C174 B.n132 VSUBS 0.007568f
C175 B.n133 VSUBS 0.007568f
C176 B.n134 VSUBS 0.007568f
C177 B.n135 VSUBS 0.007568f
C178 B.n136 VSUBS 0.007568f
C179 B.n137 VSUBS 0.007568f
C180 B.n138 VSUBS 0.007568f
C181 B.n139 VSUBS 0.007568f
C182 B.n140 VSUBS 0.007568f
C183 B.n141 VSUBS 0.007568f
C184 B.n142 VSUBS 0.007568f
C185 B.n143 VSUBS 0.007568f
C186 B.n144 VSUBS 0.007568f
C187 B.n145 VSUBS 0.007568f
C188 B.n146 VSUBS 0.007568f
C189 B.n147 VSUBS 0.007568f
C190 B.n148 VSUBS 0.007568f
C191 B.n149 VSUBS 0.007568f
C192 B.n150 VSUBS 0.016829f
C193 B.n151 VSUBS 0.007568f
C194 B.n152 VSUBS 0.007568f
C195 B.n153 VSUBS 0.007568f
C196 B.n154 VSUBS 0.007568f
C197 B.n155 VSUBS 0.007568f
C198 B.n156 VSUBS 0.007568f
C199 B.n157 VSUBS 0.007568f
C200 B.n158 VSUBS 0.007568f
C201 B.n159 VSUBS 0.007568f
C202 B.n160 VSUBS 0.007568f
C203 B.n161 VSUBS 0.007568f
C204 B.n162 VSUBS 0.007568f
C205 B.n163 VSUBS 0.007568f
C206 B.n164 VSUBS 0.007568f
C207 B.n165 VSUBS 0.007568f
C208 B.n166 VSUBS 0.007568f
C209 B.n167 VSUBS 0.007568f
C210 B.n168 VSUBS 0.007568f
C211 B.n169 VSUBS 0.016829f
C212 B.n170 VSUBS 0.017448f
C213 B.n171 VSUBS 0.017448f
C214 B.n172 VSUBS 0.007568f
C215 B.n173 VSUBS 0.007568f
C216 B.n174 VSUBS 0.007568f
C217 B.n175 VSUBS 0.007568f
C218 B.n176 VSUBS 0.007568f
C219 B.n177 VSUBS 0.007568f
C220 B.n178 VSUBS 0.007568f
C221 B.n179 VSUBS 0.007568f
C222 B.n180 VSUBS 0.007568f
C223 B.n181 VSUBS 0.007568f
C224 B.n182 VSUBS 0.007568f
C225 B.n183 VSUBS 0.007568f
C226 B.n184 VSUBS 0.007568f
C227 B.n185 VSUBS 0.007568f
C228 B.n186 VSUBS 0.007568f
C229 B.n187 VSUBS 0.007568f
C230 B.n188 VSUBS 0.007568f
C231 B.n189 VSUBS 0.007568f
C232 B.n190 VSUBS 0.007568f
C233 B.n191 VSUBS 0.007568f
C234 B.n192 VSUBS 0.007568f
C235 B.n193 VSUBS 0.007568f
C236 B.n194 VSUBS 0.007568f
C237 B.n195 VSUBS 0.007568f
C238 B.n196 VSUBS 0.007568f
C239 B.n197 VSUBS 0.007568f
C240 B.n198 VSUBS 0.007568f
C241 B.n199 VSUBS 0.007568f
C242 B.n200 VSUBS 0.007568f
C243 B.n201 VSUBS 0.007568f
C244 B.n202 VSUBS 0.007568f
C245 B.n203 VSUBS 0.007568f
C246 B.n204 VSUBS 0.007568f
C247 B.n205 VSUBS 0.007568f
C248 B.n206 VSUBS 0.007568f
C249 B.n207 VSUBS 0.007568f
C250 B.n208 VSUBS 0.007568f
C251 B.n209 VSUBS 0.007568f
C252 B.n210 VSUBS 0.007568f
C253 B.n211 VSUBS 0.007568f
C254 B.n212 VSUBS 0.007568f
C255 B.n213 VSUBS 0.007568f
C256 B.n214 VSUBS 0.007568f
C257 B.n215 VSUBS 0.007568f
C258 B.n216 VSUBS 0.007568f
C259 B.n217 VSUBS 0.007568f
C260 B.n218 VSUBS 0.007568f
C261 B.n219 VSUBS 0.007568f
C262 B.n220 VSUBS 0.007568f
C263 B.n221 VSUBS 0.007568f
C264 B.n222 VSUBS 0.007568f
C265 B.n223 VSUBS 0.007568f
C266 B.n224 VSUBS 0.007568f
C267 B.n225 VSUBS 0.007568f
C268 B.n226 VSUBS 0.007568f
C269 B.n227 VSUBS 0.007568f
C270 B.n228 VSUBS 0.007568f
C271 B.n229 VSUBS 0.007568f
C272 B.n230 VSUBS 0.007568f
C273 B.n231 VSUBS 0.007568f
C274 B.n232 VSUBS 0.007568f
C275 B.n233 VSUBS 0.007568f
C276 B.n234 VSUBS 0.007568f
C277 B.n235 VSUBS 0.007568f
C278 B.n236 VSUBS 0.007568f
C279 B.n237 VSUBS 0.007568f
C280 B.n238 VSUBS 0.007568f
C281 B.n239 VSUBS 0.007568f
C282 B.n240 VSUBS 0.007568f
C283 B.n241 VSUBS 0.007568f
C284 B.n242 VSUBS 0.007568f
C285 B.n243 VSUBS 0.007568f
C286 B.n244 VSUBS 0.007568f
C287 B.n245 VSUBS 0.007568f
C288 B.n246 VSUBS 0.007568f
C289 B.n247 VSUBS 0.007568f
C290 B.n248 VSUBS 0.007568f
C291 B.n249 VSUBS 0.007568f
C292 B.n250 VSUBS 0.007568f
C293 B.n251 VSUBS 0.007568f
C294 B.n252 VSUBS 0.007568f
C295 B.n253 VSUBS 0.007568f
C296 B.n254 VSUBS 0.007568f
C297 B.n255 VSUBS 0.0069f
C298 B.n256 VSUBS 0.017534f
C299 B.n257 VSUBS 0.004452f
C300 B.n258 VSUBS 0.007568f
C301 B.n259 VSUBS 0.007568f
C302 B.n260 VSUBS 0.007568f
C303 B.n261 VSUBS 0.007568f
C304 B.n262 VSUBS 0.007568f
C305 B.n263 VSUBS 0.007568f
C306 B.n264 VSUBS 0.007568f
C307 B.n265 VSUBS 0.007568f
C308 B.n266 VSUBS 0.007568f
C309 B.n267 VSUBS 0.007568f
C310 B.n268 VSUBS 0.007568f
C311 B.n269 VSUBS 0.007568f
C312 B.t11 VSUBS 0.629236f
C313 B.t10 VSUBS 0.634151f
C314 B.t9 VSUBS 0.158223f
C315 B.n270 VSUBS 0.110676f
C316 B.n271 VSUBS 0.06727f
C317 B.n272 VSUBS 0.017534f
C318 B.n273 VSUBS 0.004452f
C319 B.n274 VSUBS 0.007568f
C320 B.n275 VSUBS 0.007568f
C321 B.n276 VSUBS 0.007568f
C322 B.n277 VSUBS 0.007568f
C323 B.n278 VSUBS 0.007568f
C324 B.n279 VSUBS 0.007568f
C325 B.n280 VSUBS 0.007568f
C326 B.n281 VSUBS 0.007568f
C327 B.n282 VSUBS 0.007568f
C328 B.n283 VSUBS 0.007568f
C329 B.n284 VSUBS 0.007568f
C330 B.n285 VSUBS 0.007568f
C331 B.n286 VSUBS 0.007568f
C332 B.n287 VSUBS 0.007568f
C333 B.n288 VSUBS 0.007568f
C334 B.n289 VSUBS 0.007568f
C335 B.n290 VSUBS 0.007568f
C336 B.n291 VSUBS 0.007568f
C337 B.n292 VSUBS 0.007568f
C338 B.n293 VSUBS 0.007568f
C339 B.n294 VSUBS 0.007568f
C340 B.n295 VSUBS 0.007568f
C341 B.n296 VSUBS 0.007568f
C342 B.n297 VSUBS 0.007568f
C343 B.n298 VSUBS 0.007568f
C344 B.n299 VSUBS 0.007568f
C345 B.n300 VSUBS 0.007568f
C346 B.n301 VSUBS 0.007568f
C347 B.n302 VSUBS 0.007568f
C348 B.n303 VSUBS 0.007568f
C349 B.n304 VSUBS 0.007568f
C350 B.n305 VSUBS 0.007568f
C351 B.n306 VSUBS 0.007568f
C352 B.n307 VSUBS 0.007568f
C353 B.n308 VSUBS 0.007568f
C354 B.n309 VSUBS 0.007568f
C355 B.n310 VSUBS 0.007568f
C356 B.n311 VSUBS 0.007568f
C357 B.n312 VSUBS 0.007568f
C358 B.n313 VSUBS 0.007568f
C359 B.n314 VSUBS 0.007568f
C360 B.n315 VSUBS 0.007568f
C361 B.n316 VSUBS 0.007568f
C362 B.n317 VSUBS 0.007568f
C363 B.n318 VSUBS 0.007568f
C364 B.n319 VSUBS 0.007568f
C365 B.n320 VSUBS 0.007568f
C366 B.n321 VSUBS 0.007568f
C367 B.n322 VSUBS 0.007568f
C368 B.n323 VSUBS 0.007568f
C369 B.n324 VSUBS 0.007568f
C370 B.n325 VSUBS 0.007568f
C371 B.n326 VSUBS 0.007568f
C372 B.n327 VSUBS 0.007568f
C373 B.n328 VSUBS 0.007568f
C374 B.n329 VSUBS 0.007568f
C375 B.n330 VSUBS 0.007568f
C376 B.n331 VSUBS 0.007568f
C377 B.n332 VSUBS 0.007568f
C378 B.n333 VSUBS 0.007568f
C379 B.n334 VSUBS 0.007568f
C380 B.n335 VSUBS 0.007568f
C381 B.n336 VSUBS 0.007568f
C382 B.n337 VSUBS 0.007568f
C383 B.n338 VSUBS 0.007568f
C384 B.n339 VSUBS 0.007568f
C385 B.n340 VSUBS 0.007568f
C386 B.n341 VSUBS 0.007568f
C387 B.n342 VSUBS 0.007568f
C388 B.n343 VSUBS 0.007568f
C389 B.n344 VSUBS 0.007568f
C390 B.n345 VSUBS 0.007568f
C391 B.n346 VSUBS 0.007568f
C392 B.n347 VSUBS 0.007568f
C393 B.n348 VSUBS 0.007568f
C394 B.n349 VSUBS 0.007568f
C395 B.n350 VSUBS 0.007568f
C396 B.n351 VSUBS 0.007568f
C397 B.n352 VSUBS 0.007568f
C398 B.n353 VSUBS 0.007568f
C399 B.n354 VSUBS 0.007568f
C400 B.n355 VSUBS 0.007568f
C401 B.n356 VSUBS 0.007568f
C402 B.n357 VSUBS 0.007568f
C403 B.n358 VSUBS 0.007568f
C404 B.n359 VSUBS 0.017448f
C405 B.n360 VSUBS 0.016829f
C406 B.n361 VSUBS 0.017769f
C407 B.n362 VSUBS 0.007568f
C408 B.n363 VSUBS 0.007568f
C409 B.n364 VSUBS 0.007568f
C410 B.n365 VSUBS 0.007568f
C411 B.n366 VSUBS 0.007568f
C412 B.n367 VSUBS 0.007568f
C413 B.n368 VSUBS 0.007568f
C414 B.n369 VSUBS 0.007568f
C415 B.n370 VSUBS 0.007568f
C416 B.n371 VSUBS 0.007568f
C417 B.n372 VSUBS 0.007568f
C418 B.n373 VSUBS 0.007568f
C419 B.n374 VSUBS 0.007568f
C420 B.n375 VSUBS 0.007568f
C421 B.n376 VSUBS 0.007568f
C422 B.n377 VSUBS 0.007568f
C423 B.n378 VSUBS 0.007568f
C424 B.n379 VSUBS 0.007568f
C425 B.n380 VSUBS 0.007568f
C426 B.n381 VSUBS 0.007568f
C427 B.n382 VSUBS 0.007568f
C428 B.n383 VSUBS 0.007568f
C429 B.n384 VSUBS 0.007568f
C430 B.n385 VSUBS 0.007568f
C431 B.n386 VSUBS 0.007568f
C432 B.n387 VSUBS 0.007568f
C433 B.n388 VSUBS 0.007568f
C434 B.n389 VSUBS 0.007568f
C435 B.n390 VSUBS 0.007568f
C436 B.n391 VSUBS 0.007568f
C437 B.n392 VSUBS 0.007568f
C438 B.n393 VSUBS 0.007568f
C439 B.n394 VSUBS 0.007568f
C440 B.n395 VSUBS 0.016829f
C441 B.n396 VSUBS 0.017448f
C442 B.n397 VSUBS 0.017448f
C443 B.n398 VSUBS 0.007568f
C444 B.n399 VSUBS 0.007568f
C445 B.n400 VSUBS 0.007568f
C446 B.n401 VSUBS 0.007568f
C447 B.n402 VSUBS 0.007568f
C448 B.n403 VSUBS 0.007568f
C449 B.n404 VSUBS 0.007568f
C450 B.n405 VSUBS 0.007568f
C451 B.n406 VSUBS 0.007568f
C452 B.n407 VSUBS 0.007568f
C453 B.n408 VSUBS 0.007568f
C454 B.n409 VSUBS 0.007568f
C455 B.n410 VSUBS 0.007568f
C456 B.n411 VSUBS 0.007568f
C457 B.n412 VSUBS 0.007568f
C458 B.n413 VSUBS 0.007568f
C459 B.n414 VSUBS 0.007568f
C460 B.n415 VSUBS 0.007568f
C461 B.n416 VSUBS 0.007568f
C462 B.n417 VSUBS 0.007568f
C463 B.n418 VSUBS 0.007568f
C464 B.n419 VSUBS 0.007568f
C465 B.n420 VSUBS 0.007568f
C466 B.n421 VSUBS 0.007568f
C467 B.n422 VSUBS 0.007568f
C468 B.n423 VSUBS 0.007568f
C469 B.n424 VSUBS 0.007568f
C470 B.n425 VSUBS 0.007568f
C471 B.n426 VSUBS 0.007568f
C472 B.n427 VSUBS 0.007568f
C473 B.n428 VSUBS 0.007568f
C474 B.n429 VSUBS 0.007568f
C475 B.n430 VSUBS 0.007568f
C476 B.n431 VSUBS 0.007568f
C477 B.n432 VSUBS 0.007568f
C478 B.n433 VSUBS 0.007568f
C479 B.n434 VSUBS 0.007568f
C480 B.n435 VSUBS 0.007568f
C481 B.n436 VSUBS 0.007568f
C482 B.n437 VSUBS 0.007568f
C483 B.n438 VSUBS 0.007568f
C484 B.n439 VSUBS 0.007568f
C485 B.n440 VSUBS 0.007568f
C486 B.n441 VSUBS 0.007568f
C487 B.n442 VSUBS 0.007568f
C488 B.n443 VSUBS 0.007568f
C489 B.n444 VSUBS 0.007568f
C490 B.n445 VSUBS 0.007568f
C491 B.n446 VSUBS 0.007568f
C492 B.n447 VSUBS 0.007568f
C493 B.n448 VSUBS 0.007568f
C494 B.n449 VSUBS 0.007568f
C495 B.n450 VSUBS 0.007568f
C496 B.n451 VSUBS 0.007568f
C497 B.n452 VSUBS 0.007568f
C498 B.n453 VSUBS 0.007568f
C499 B.n454 VSUBS 0.007568f
C500 B.n455 VSUBS 0.007568f
C501 B.n456 VSUBS 0.007568f
C502 B.n457 VSUBS 0.007568f
C503 B.n458 VSUBS 0.007568f
C504 B.n459 VSUBS 0.007568f
C505 B.n460 VSUBS 0.007568f
C506 B.n461 VSUBS 0.007568f
C507 B.n462 VSUBS 0.007568f
C508 B.n463 VSUBS 0.007568f
C509 B.n464 VSUBS 0.007568f
C510 B.n465 VSUBS 0.007568f
C511 B.n466 VSUBS 0.007568f
C512 B.n467 VSUBS 0.007568f
C513 B.n468 VSUBS 0.007568f
C514 B.n469 VSUBS 0.007568f
C515 B.n470 VSUBS 0.007568f
C516 B.n471 VSUBS 0.007568f
C517 B.n472 VSUBS 0.007568f
C518 B.n473 VSUBS 0.007568f
C519 B.n474 VSUBS 0.007568f
C520 B.n475 VSUBS 0.007568f
C521 B.n476 VSUBS 0.007568f
C522 B.n477 VSUBS 0.007568f
C523 B.n478 VSUBS 0.007568f
C524 B.n479 VSUBS 0.007568f
C525 B.n480 VSUBS 0.007568f
C526 B.n481 VSUBS 0.0069f
C527 B.n482 VSUBS 0.017534f
C528 B.n483 VSUBS 0.004452f
C529 B.n484 VSUBS 0.007568f
C530 B.n485 VSUBS 0.007568f
C531 B.n486 VSUBS 0.007568f
C532 B.n487 VSUBS 0.007568f
C533 B.n488 VSUBS 0.007568f
C534 B.n489 VSUBS 0.007568f
C535 B.n490 VSUBS 0.007568f
C536 B.n491 VSUBS 0.007568f
C537 B.n492 VSUBS 0.007568f
C538 B.n493 VSUBS 0.007568f
C539 B.n494 VSUBS 0.007568f
C540 B.n495 VSUBS 0.007568f
C541 B.n496 VSUBS 0.004452f
C542 B.n497 VSUBS 0.007568f
C543 B.n498 VSUBS 0.007568f
C544 B.n499 VSUBS 0.0069f
C545 B.n500 VSUBS 0.007568f
C546 B.n501 VSUBS 0.007568f
C547 B.n502 VSUBS 0.007568f
C548 B.n503 VSUBS 0.007568f
C549 B.n504 VSUBS 0.007568f
C550 B.n505 VSUBS 0.007568f
C551 B.n506 VSUBS 0.007568f
C552 B.n507 VSUBS 0.007568f
C553 B.n508 VSUBS 0.007568f
C554 B.n509 VSUBS 0.007568f
C555 B.n510 VSUBS 0.007568f
C556 B.n511 VSUBS 0.007568f
C557 B.n512 VSUBS 0.007568f
C558 B.n513 VSUBS 0.007568f
C559 B.n514 VSUBS 0.007568f
C560 B.n515 VSUBS 0.007568f
C561 B.n516 VSUBS 0.007568f
C562 B.n517 VSUBS 0.007568f
C563 B.n518 VSUBS 0.007568f
C564 B.n519 VSUBS 0.007568f
C565 B.n520 VSUBS 0.007568f
C566 B.n521 VSUBS 0.007568f
C567 B.n522 VSUBS 0.007568f
C568 B.n523 VSUBS 0.007568f
C569 B.n524 VSUBS 0.007568f
C570 B.n525 VSUBS 0.007568f
C571 B.n526 VSUBS 0.007568f
C572 B.n527 VSUBS 0.007568f
C573 B.n528 VSUBS 0.007568f
C574 B.n529 VSUBS 0.007568f
C575 B.n530 VSUBS 0.007568f
C576 B.n531 VSUBS 0.007568f
C577 B.n532 VSUBS 0.007568f
C578 B.n533 VSUBS 0.007568f
C579 B.n534 VSUBS 0.007568f
C580 B.n535 VSUBS 0.007568f
C581 B.n536 VSUBS 0.007568f
C582 B.n537 VSUBS 0.007568f
C583 B.n538 VSUBS 0.007568f
C584 B.n539 VSUBS 0.007568f
C585 B.n540 VSUBS 0.007568f
C586 B.n541 VSUBS 0.007568f
C587 B.n542 VSUBS 0.007568f
C588 B.n543 VSUBS 0.007568f
C589 B.n544 VSUBS 0.007568f
C590 B.n545 VSUBS 0.007568f
C591 B.n546 VSUBS 0.007568f
C592 B.n547 VSUBS 0.007568f
C593 B.n548 VSUBS 0.007568f
C594 B.n549 VSUBS 0.007568f
C595 B.n550 VSUBS 0.007568f
C596 B.n551 VSUBS 0.007568f
C597 B.n552 VSUBS 0.007568f
C598 B.n553 VSUBS 0.007568f
C599 B.n554 VSUBS 0.007568f
C600 B.n555 VSUBS 0.007568f
C601 B.n556 VSUBS 0.007568f
C602 B.n557 VSUBS 0.007568f
C603 B.n558 VSUBS 0.007568f
C604 B.n559 VSUBS 0.007568f
C605 B.n560 VSUBS 0.007568f
C606 B.n561 VSUBS 0.007568f
C607 B.n562 VSUBS 0.007568f
C608 B.n563 VSUBS 0.007568f
C609 B.n564 VSUBS 0.007568f
C610 B.n565 VSUBS 0.007568f
C611 B.n566 VSUBS 0.007568f
C612 B.n567 VSUBS 0.007568f
C613 B.n568 VSUBS 0.007568f
C614 B.n569 VSUBS 0.007568f
C615 B.n570 VSUBS 0.007568f
C616 B.n571 VSUBS 0.007568f
C617 B.n572 VSUBS 0.007568f
C618 B.n573 VSUBS 0.007568f
C619 B.n574 VSUBS 0.007568f
C620 B.n575 VSUBS 0.007568f
C621 B.n576 VSUBS 0.007568f
C622 B.n577 VSUBS 0.007568f
C623 B.n578 VSUBS 0.007568f
C624 B.n579 VSUBS 0.007568f
C625 B.n580 VSUBS 0.007568f
C626 B.n581 VSUBS 0.007568f
C627 B.n582 VSUBS 0.017448f
C628 B.n583 VSUBS 0.017448f
C629 B.n584 VSUBS 0.016829f
C630 B.n585 VSUBS 0.007568f
C631 B.n586 VSUBS 0.007568f
C632 B.n587 VSUBS 0.007568f
C633 B.n588 VSUBS 0.007568f
C634 B.n589 VSUBS 0.007568f
C635 B.n590 VSUBS 0.007568f
C636 B.n591 VSUBS 0.007568f
C637 B.n592 VSUBS 0.007568f
C638 B.n593 VSUBS 0.007568f
C639 B.n594 VSUBS 0.007568f
C640 B.n595 VSUBS 0.007568f
C641 B.n596 VSUBS 0.007568f
C642 B.n597 VSUBS 0.007568f
C643 B.n598 VSUBS 0.007568f
C644 B.n599 VSUBS 0.009875f
C645 B.n600 VSUBS 0.01052f
C646 B.n601 VSUBS 0.02092f
C647 VDD1.t0 VSUBS 3.08813f
C648 VDD1.t1 VSUBS 3.73293f
C649 VTAIL.t3 VSUBS 4.20613f
C650 VTAIL.n0 VSUBS 2.83592f
C651 VTAIL.t0 VSUBS 4.20616f
C652 VTAIL.n1 VSUBS 2.8417f
C653 VTAIL.t2 VSUBS 4.20613f
C654 VTAIL.n2 VSUBS 2.796f
C655 VTAIL.t1 VSUBS 4.20613f
C656 VTAIL.n3 VSUBS 2.73364f
C657 VP.t1 VSUBS 0.552894f
C658 VP.t0 VSUBS 0.513304f
C659 VP.n0 VSUBS 4.22823f
.ends

