* NGSPICE file created from diff_pair_sample_1055.ext - technology: sky130A

.subckt diff_pair_sample_1055 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t1 VN.t0 VTAIL.t2 w_n2678_n4294# sky130_fd_pr__pfet_01v8 ad=6.4857 pd=34.04 as=6.4857 ps=34.04 w=16.63 l=3.94
X1 B.t11 B.t9 B.t10 w_n2678_n4294# sky130_fd_pr__pfet_01v8 ad=6.4857 pd=34.04 as=0 ps=0 w=16.63 l=3.94
X2 B.t8 B.t6 B.t7 w_n2678_n4294# sky130_fd_pr__pfet_01v8 ad=6.4857 pd=34.04 as=0 ps=0 w=16.63 l=3.94
X3 B.t5 B.t3 B.t4 w_n2678_n4294# sky130_fd_pr__pfet_01v8 ad=6.4857 pd=34.04 as=0 ps=0 w=16.63 l=3.94
X4 VDD2.t0 VN.t1 VTAIL.t3 w_n2678_n4294# sky130_fd_pr__pfet_01v8 ad=6.4857 pd=34.04 as=6.4857 ps=34.04 w=16.63 l=3.94
X5 VDD1.t1 VP.t0 VTAIL.t0 w_n2678_n4294# sky130_fd_pr__pfet_01v8 ad=6.4857 pd=34.04 as=6.4857 ps=34.04 w=16.63 l=3.94
X6 B.t2 B.t0 B.t1 w_n2678_n4294# sky130_fd_pr__pfet_01v8 ad=6.4857 pd=34.04 as=0 ps=0 w=16.63 l=3.94
X7 VDD1.t0 VP.t1 VTAIL.t1 w_n2678_n4294# sky130_fd_pr__pfet_01v8 ad=6.4857 pd=34.04 as=6.4857 ps=34.04 w=16.63 l=3.94
R0 VN VN.t1 188.29
R1 VN VN.t0 137.38
R2 VTAIL.n1 VTAIL.t3 58.5521
R3 VTAIL.n3 VTAIL.t2 58.5519
R4 VTAIL.n0 VTAIL.t0 58.5519
R5 VTAIL.n2 VTAIL.t1 58.5519
R6 VTAIL.n1 VTAIL.n0 34.0652
R7 VTAIL.n3 VTAIL.n2 30.3841
R8 VTAIL.n2 VTAIL.n1 2.31084
R9 VTAIL VTAIL.n0 1.44878
R10 VTAIL VTAIL.n3 0.862569
R11 VDD2.n0 VDD2.t1 120.588
R12 VDD2.n0 VDD2.t0 75.2307
R13 VDD2 VDD2.n0 0.978948
R14 B.n528 B.n527 585
R15 B.n529 B.n82 585
R16 B.n531 B.n530 585
R17 B.n532 B.n81 585
R18 B.n534 B.n533 585
R19 B.n535 B.n80 585
R20 B.n537 B.n536 585
R21 B.n538 B.n79 585
R22 B.n540 B.n539 585
R23 B.n541 B.n78 585
R24 B.n543 B.n542 585
R25 B.n544 B.n77 585
R26 B.n546 B.n545 585
R27 B.n547 B.n76 585
R28 B.n549 B.n548 585
R29 B.n550 B.n75 585
R30 B.n552 B.n551 585
R31 B.n553 B.n74 585
R32 B.n555 B.n554 585
R33 B.n556 B.n73 585
R34 B.n558 B.n557 585
R35 B.n559 B.n72 585
R36 B.n561 B.n560 585
R37 B.n562 B.n71 585
R38 B.n564 B.n563 585
R39 B.n565 B.n70 585
R40 B.n567 B.n566 585
R41 B.n568 B.n69 585
R42 B.n570 B.n569 585
R43 B.n571 B.n68 585
R44 B.n573 B.n572 585
R45 B.n574 B.n67 585
R46 B.n576 B.n575 585
R47 B.n577 B.n66 585
R48 B.n579 B.n578 585
R49 B.n580 B.n65 585
R50 B.n582 B.n581 585
R51 B.n583 B.n64 585
R52 B.n585 B.n584 585
R53 B.n586 B.n63 585
R54 B.n588 B.n587 585
R55 B.n589 B.n62 585
R56 B.n591 B.n590 585
R57 B.n592 B.n61 585
R58 B.n594 B.n593 585
R59 B.n595 B.n60 585
R60 B.n597 B.n596 585
R61 B.n598 B.n59 585
R62 B.n600 B.n599 585
R63 B.n601 B.n58 585
R64 B.n603 B.n602 585
R65 B.n604 B.n57 585
R66 B.n606 B.n605 585
R67 B.n607 B.n56 585
R68 B.n609 B.n608 585
R69 B.n611 B.n53 585
R70 B.n613 B.n612 585
R71 B.n614 B.n52 585
R72 B.n616 B.n615 585
R73 B.n617 B.n51 585
R74 B.n619 B.n618 585
R75 B.n620 B.n50 585
R76 B.n622 B.n621 585
R77 B.n623 B.n49 585
R78 B.n625 B.n624 585
R79 B.n627 B.n626 585
R80 B.n628 B.n45 585
R81 B.n630 B.n629 585
R82 B.n631 B.n44 585
R83 B.n633 B.n632 585
R84 B.n634 B.n43 585
R85 B.n636 B.n635 585
R86 B.n637 B.n42 585
R87 B.n639 B.n638 585
R88 B.n640 B.n41 585
R89 B.n642 B.n641 585
R90 B.n643 B.n40 585
R91 B.n645 B.n644 585
R92 B.n646 B.n39 585
R93 B.n648 B.n647 585
R94 B.n649 B.n38 585
R95 B.n651 B.n650 585
R96 B.n652 B.n37 585
R97 B.n654 B.n653 585
R98 B.n655 B.n36 585
R99 B.n657 B.n656 585
R100 B.n658 B.n35 585
R101 B.n660 B.n659 585
R102 B.n661 B.n34 585
R103 B.n663 B.n662 585
R104 B.n664 B.n33 585
R105 B.n666 B.n665 585
R106 B.n667 B.n32 585
R107 B.n669 B.n668 585
R108 B.n670 B.n31 585
R109 B.n672 B.n671 585
R110 B.n673 B.n30 585
R111 B.n675 B.n674 585
R112 B.n676 B.n29 585
R113 B.n678 B.n677 585
R114 B.n679 B.n28 585
R115 B.n681 B.n680 585
R116 B.n682 B.n27 585
R117 B.n684 B.n683 585
R118 B.n685 B.n26 585
R119 B.n687 B.n686 585
R120 B.n688 B.n25 585
R121 B.n690 B.n689 585
R122 B.n691 B.n24 585
R123 B.n693 B.n692 585
R124 B.n694 B.n23 585
R125 B.n696 B.n695 585
R126 B.n697 B.n22 585
R127 B.n699 B.n698 585
R128 B.n700 B.n21 585
R129 B.n702 B.n701 585
R130 B.n703 B.n20 585
R131 B.n705 B.n704 585
R132 B.n706 B.n19 585
R133 B.n708 B.n707 585
R134 B.n526 B.n83 585
R135 B.n525 B.n524 585
R136 B.n523 B.n84 585
R137 B.n522 B.n521 585
R138 B.n520 B.n85 585
R139 B.n519 B.n518 585
R140 B.n517 B.n86 585
R141 B.n516 B.n515 585
R142 B.n514 B.n87 585
R143 B.n513 B.n512 585
R144 B.n511 B.n88 585
R145 B.n510 B.n509 585
R146 B.n508 B.n89 585
R147 B.n507 B.n506 585
R148 B.n505 B.n90 585
R149 B.n504 B.n503 585
R150 B.n502 B.n91 585
R151 B.n501 B.n500 585
R152 B.n499 B.n92 585
R153 B.n498 B.n497 585
R154 B.n496 B.n93 585
R155 B.n495 B.n494 585
R156 B.n493 B.n94 585
R157 B.n492 B.n491 585
R158 B.n490 B.n95 585
R159 B.n489 B.n488 585
R160 B.n487 B.n96 585
R161 B.n486 B.n485 585
R162 B.n484 B.n97 585
R163 B.n483 B.n482 585
R164 B.n481 B.n98 585
R165 B.n480 B.n479 585
R166 B.n478 B.n99 585
R167 B.n477 B.n476 585
R168 B.n475 B.n100 585
R169 B.n474 B.n473 585
R170 B.n472 B.n101 585
R171 B.n471 B.n470 585
R172 B.n469 B.n102 585
R173 B.n468 B.n467 585
R174 B.n466 B.n103 585
R175 B.n465 B.n464 585
R176 B.n463 B.n104 585
R177 B.n462 B.n461 585
R178 B.n460 B.n105 585
R179 B.n459 B.n458 585
R180 B.n457 B.n106 585
R181 B.n456 B.n455 585
R182 B.n454 B.n107 585
R183 B.n453 B.n452 585
R184 B.n451 B.n108 585
R185 B.n450 B.n449 585
R186 B.n448 B.n109 585
R187 B.n447 B.n446 585
R188 B.n445 B.n110 585
R189 B.n444 B.n443 585
R190 B.n442 B.n111 585
R191 B.n441 B.n440 585
R192 B.n439 B.n112 585
R193 B.n438 B.n437 585
R194 B.n436 B.n113 585
R195 B.n435 B.n434 585
R196 B.n433 B.n114 585
R197 B.n432 B.n431 585
R198 B.n430 B.n115 585
R199 B.n429 B.n428 585
R200 B.n427 B.n116 585
R201 B.n246 B.n245 585
R202 B.n247 B.n180 585
R203 B.n249 B.n248 585
R204 B.n250 B.n179 585
R205 B.n252 B.n251 585
R206 B.n253 B.n178 585
R207 B.n255 B.n254 585
R208 B.n256 B.n177 585
R209 B.n258 B.n257 585
R210 B.n259 B.n176 585
R211 B.n261 B.n260 585
R212 B.n262 B.n175 585
R213 B.n264 B.n263 585
R214 B.n265 B.n174 585
R215 B.n267 B.n266 585
R216 B.n268 B.n173 585
R217 B.n270 B.n269 585
R218 B.n271 B.n172 585
R219 B.n273 B.n272 585
R220 B.n274 B.n171 585
R221 B.n276 B.n275 585
R222 B.n277 B.n170 585
R223 B.n279 B.n278 585
R224 B.n280 B.n169 585
R225 B.n282 B.n281 585
R226 B.n283 B.n168 585
R227 B.n285 B.n284 585
R228 B.n286 B.n167 585
R229 B.n288 B.n287 585
R230 B.n289 B.n166 585
R231 B.n291 B.n290 585
R232 B.n292 B.n165 585
R233 B.n294 B.n293 585
R234 B.n295 B.n164 585
R235 B.n297 B.n296 585
R236 B.n298 B.n163 585
R237 B.n300 B.n299 585
R238 B.n301 B.n162 585
R239 B.n303 B.n302 585
R240 B.n304 B.n161 585
R241 B.n306 B.n305 585
R242 B.n307 B.n160 585
R243 B.n309 B.n308 585
R244 B.n310 B.n159 585
R245 B.n312 B.n311 585
R246 B.n313 B.n158 585
R247 B.n315 B.n314 585
R248 B.n316 B.n157 585
R249 B.n318 B.n317 585
R250 B.n319 B.n156 585
R251 B.n321 B.n320 585
R252 B.n322 B.n155 585
R253 B.n324 B.n323 585
R254 B.n325 B.n154 585
R255 B.n327 B.n326 585
R256 B.n329 B.n151 585
R257 B.n331 B.n330 585
R258 B.n332 B.n150 585
R259 B.n334 B.n333 585
R260 B.n335 B.n149 585
R261 B.n337 B.n336 585
R262 B.n338 B.n148 585
R263 B.n340 B.n339 585
R264 B.n341 B.n147 585
R265 B.n343 B.n342 585
R266 B.n345 B.n344 585
R267 B.n346 B.n143 585
R268 B.n348 B.n347 585
R269 B.n349 B.n142 585
R270 B.n351 B.n350 585
R271 B.n352 B.n141 585
R272 B.n354 B.n353 585
R273 B.n355 B.n140 585
R274 B.n357 B.n356 585
R275 B.n358 B.n139 585
R276 B.n360 B.n359 585
R277 B.n361 B.n138 585
R278 B.n363 B.n362 585
R279 B.n364 B.n137 585
R280 B.n366 B.n365 585
R281 B.n367 B.n136 585
R282 B.n369 B.n368 585
R283 B.n370 B.n135 585
R284 B.n372 B.n371 585
R285 B.n373 B.n134 585
R286 B.n375 B.n374 585
R287 B.n376 B.n133 585
R288 B.n378 B.n377 585
R289 B.n379 B.n132 585
R290 B.n381 B.n380 585
R291 B.n382 B.n131 585
R292 B.n384 B.n383 585
R293 B.n385 B.n130 585
R294 B.n387 B.n386 585
R295 B.n388 B.n129 585
R296 B.n390 B.n389 585
R297 B.n391 B.n128 585
R298 B.n393 B.n392 585
R299 B.n394 B.n127 585
R300 B.n396 B.n395 585
R301 B.n397 B.n126 585
R302 B.n399 B.n398 585
R303 B.n400 B.n125 585
R304 B.n402 B.n401 585
R305 B.n403 B.n124 585
R306 B.n405 B.n404 585
R307 B.n406 B.n123 585
R308 B.n408 B.n407 585
R309 B.n409 B.n122 585
R310 B.n411 B.n410 585
R311 B.n412 B.n121 585
R312 B.n414 B.n413 585
R313 B.n415 B.n120 585
R314 B.n417 B.n416 585
R315 B.n418 B.n119 585
R316 B.n420 B.n419 585
R317 B.n421 B.n118 585
R318 B.n423 B.n422 585
R319 B.n424 B.n117 585
R320 B.n426 B.n425 585
R321 B.n244 B.n181 585
R322 B.n243 B.n242 585
R323 B.n241 B.n182 585
R324 B.n240 B.n239 585
R325 B.n238 B.n183 585
R326 B.n237 B.n236 585
R327 B.n235 B.n184 585
R328 B.n234 B.n233 585
R329 B.n232 B.n185 585
R330 B.n231 B.n230 585
R331 B.n229 B.n186 585
R332 B.n228 B.n227 585
R333 B.n226 B.n187 585
R334 B.n225 B.n224 585
R335 B.n223 B.n188 585
R336 B.n222 B.n221 585
R337 B.n220 B.n189 585
R338 B.n219 B.n218 585
R339 B.n217 B.n190 585
R340 B.n216 B.n215 585
R341 B.n214 B.n191 585
R342 B.n213 B.n212 585
R343 B.n211 B.n192 585
R344 B.n210 B.n209 585
R345 B.n208 B.n193 585
R346 B.n207 B.n206 585
R347 B.n205 B.n194 585
R348 B.n204 B.n203 585
R349 B.n202 B.n195 585
R350 B.n201 B.n200 585
R351 B.n199 B.n196 585
R352 B.n198 B.n197 585
R353 B.n2 B.n0 585
R354 B.n757 B.n1 585
R355 B.n756 B.n755 585
R356 B.n754 B.n3 585
R357 B.n753 B.n752 585
R358 B.n751 B.n4 585
R359 B.n750 B.n749 585
R360 B.n748 B.n5 585
R361 B.n747 B.n746 585
R362 B.n745 B.n6 585
R363 B.n744 B.n743 585
R364 B.n742 B.n7 585
R365 B.n741 B.n740 585
R366 B.n739 B.n8 585
R367 B.n738 B.n737 585
R368 B.n736 B.n9 585
R369 B.n735 B.n734 585
R370 B.n733 B.n10 585
R371 B.n732 B.n731 585
R372 B.n730 B.n11 585
R373 B.n729 B.n728 585
R374 B.n727 B.n12 585
R375 B.n726 B.n725 585
R376 B.n724 B.n13 585
R377 B.n723 B.n722 585
R378 B.n721 B.n14 585
R379 B.n720 B.n719 585
R380 B.n718 B.n15 585
R381 B.n717 B.n716 585
R382 B.n715 B.n16 585
R383 B.n714 B.n713 585
R384 B.n712 B.n17 585
R385 B.n711 B.n710 585
R386 B.n709 B.n18 585
R387 B.n759 B.n758 585
R388 B.n246 B.n181 540.549
R389 B.n709 B.n708 540.549
R390 B.n427 B.n426 540.549
R391 B.n528 B.n83 540.549
R392 B.n144 B.t3 311.171
R393 B.n152 B.t6 311.171
R394 B.n46 B.t9 311.171
R395 B.n54 B.t0 311.171
R396 B.n144 B.t5 195.174
R397 B.n54 B.t1 195.174
R398 B.n152 B.t8 195.154
R399 B.n46 B.t10 195.154
R400 B.n242 B.n181 163.367
R401 B.n242 B.n241 163.367
R402 B.n241 B.n240 163.367
R403 B.n240 B.n183 163.367
R404 B.n236 B.n183 163.367
R405 B.n236 B.n235 163.367
R406 B.n235 B.n234 163.367
R407 B.n234 B.n185 163.367
R408 B.n230 B.n185 163.367
R409 B.n230 B.n229 163.367
R410 B.n229 B.n228 163.367
R411 B.n228 B.n187 163.367
R412 B.n224 B.n187 163.367
R413 B.n224 B.n223 163.367
R414 B.n223 B.n222 163.367
R415 B.n222 B.n189 163.367
R416 B.n218 B.n189 163.367
R417 B.n218 B.n217 163.367
R418 B.n217 B.n216 163.367
R419 B.n216 B.n191 163.367
R420 B.n212 B.n191 163.367
R421 B.n212 B.n211 163.367
R422 B.n211 B.n210 163.367
R423 B.n210 B.n193 163.367
R424 B.n206 B.n193 163.367
R425 B.n206 B.n205 163.367
R426 B.n205 B.n204 163.367
R427 B.n204 B.n195 163.367
R428 B.n200 B.n195 163.367
R429 B.n200 B.n199 163.367
R430 B.n199 B.n198 163.367
R431 B.n198 B.n2 163.367
R432 B.n758 B.n2 163.367
R433 B.n758 B.n757 163.367
R434 B.n757 B.n756 163.367
R435 B.n756 B.n3 163.367
R436 B.n752 B.n3 163.367
R437 B.n752 B.n751 163.367
R438 B.n751 B.n750 163.367
R439 B.n750 B.n5 163.367
R440 B.n746 B.n5 163.367
R441 B.n746 B.n745 163.367
R442 B.n745 B.n744 163.367
R443 B.n744 B.n7 163.367
R444 B.n740 B.n7 163.367
R445 B.n740 B.n739 163.367
R446 B.n739 B.n738 163.367
R447 B.n738 B.n9 163.367
R448 B.n734 B.n9 163.367
R449 B.n734 B.n733 163.367
R450 B.n733 B.n732 163.367
R451 B.n732 B.n11 163.367
R452 B.n728 B.n11 163.367
R453 B.n728 B.n727 163.367
R454 B.n727 B.n726 163.367
R455 B.n726 B.n13 163.367
R456 B.n722 B.n13 163.367
R457 B.n722 B.n721 163.367
R458 B.n721 B.n720 163.367
R459 B.n720 B.n15 163.367
R460 B.n716 B.n15 163.367
R461 B.n716 B.n715 163.367
R462 B.n715 B.n714 163.367
R463 B.n714 B.n17 163.367
R464 B.n710 B.n17 163.367
R465 B.n710 B.n709 163.367
R466 B.n247 B.n246 163.367
R467 B.n248 B.n247 163.367
R468 B.n248 B.n179 163.367
R469 B.n252 B.n179 163.367
R470 B.n253 B.n252 163.367
R471 B.n254 B.n253 163.367
R472 B.n254 B.n177 163.367
R473 B.n258 B.n177 163.367
R474 B.n259 B.n258 163.367
R475 B.n260 B.n259 163.367
R476 B.n260 B.n175 163.367
R477 B.n264 B.n175 163.367
R478 B.n265 B.n264 163.367
R479 B.n266 B.n265 163.367
R480 B.n266 B.n173 163.367
R481 B.n270 B.n173 163.367
R482 B.n271 B.n270 163.367
R483 B.n272 B.n271 163.367
R484 B.n272 B.n171 163.367
R485 B.n276 B.n171 163.367
R486 B.n277 B.n276 163.367
R487 B.n278 B.n277 163.367
R488 B.n278 B.n169 163.367
R489 B.n282 B.n169 163.367
R490 B.n283 B.n282 163.367
R491 B.n284 B.n283 163.367
R492 B.n284 B.n167 163.367
R493 B.n288 B.n167 163.367
R494 B.n289 B.n288 163.367
R495 B.n290 B.n289 163.367
R496 B.n290 B.n165 163.367
R497 B.n294 B.n165 163.367
R498 B.n295 B.n294 163.367
R499 B.n296 B.n295 163.367
R500 B.n296 B.n163 163.367
R501 B.n300 B.n163 163.367
R502 B.n301 B.n300 163.367
R503 B.n302 B.n301 163.367
R504 B.n302 B.n161 163.367
R505 B.n306 B.n161 163.367
R506 B.n307 B.n306 163.367
R507 B.n308 B.n307 163.367
R508 B.n308 B.n159 163.367
R509 B.n312 B.n159 163.367
R510 B.n313 B.n312 163.367
R511 B.n314 B.n313 163.367
R512 B.n314 B.n157 163.367
R513 B.n318 B.n157 163.367
R514 B.n319 B.n318 163.367
R515 B.n320 B.n319 163.367
R516 B.n320 B.n155 163.367
R517 B.n324 B.n155 163.367
R518 B.n325 B.n324 163.367
R519 B.n326 B.n325 163.367
R520 B.n326 B.n151 163.367
R521 B.n331 B.n151 163.367
R522 B.n332 B.n331 163.367
R523 B.n333 B.n332 163.367
R524 B.n333 B.n149 163.367
R525 B.n337 B.n149 163.367
R526 B.n338 B.n337 163.367
R527 B.n339 B.n338 163.367
R528 B.n339 B.n147 163.367
R529 B.n343 B.n147 163.367
R530 B.n344 B.n343 163.367
R531 B.n344 B.n143 163.367
R532 B.n348 B.n143 163.367
R533 B.n349 B.n348 163.367
R534 B.n350 B.n349 163.367
R535 B.n350 B.n141 163.367
R536 B.n354 B.n141 163.367
R537 B.n355 B.n354 163.367
R538 B.n356 B.n355 163.367
R539 B.n356 B.n139 163.367
R540 B.n360 B.n139 163.367
R541 B.n361 B.n360 163.367
R542 B.n362 B.n361 163.367
R543 B.n362 B.n137 163.367
R544 B.n366 B.n137 163.367
R545 B.n367 B.n366 163.367
R546 B.n368 B.n367 163.367
R547 B.n368 B.n135 163.367
R548 B.n372 B.n135 163.367
R549 B.n373 B.n372 163.367
R550 B.n374 B.n373 163.367
R551 B.n374 B.n133 163.367
R552 B.n378 B.n133 163.367
R553 B.n379 B.n378 163.367
R554 B.n380 B.n379 163.367
R555 B.n380 B.n131 163.367
R556 B.n384 B.n131 163.367
R557 B.n385 B.n384 163.367
R558 B.n386 B.n385 163.367
R559 B.n386 B.n129 163.367
R560 B.n390 B.n129 163.367
R561 B.n391 B.n390 163.367
R562 B.n392 B.n391 163.367
R563 B.n392 B.n127 163.367
R564 B.n396 B.n127 163.367
R565 B.n397 B.n396 163.367
R566 B.n398 B.n397 163.367
R567 B.n398 B.n125 163.367
R568 B.n402 B.n125 163.367
R569 B.n403 B.n402 163.367
R570 B.n404 B.n403 163.367
R571 B.n404 B.n123 163.367
R572 B.n408 B.n123 163.367
R573 B.n409 B.n408 163.367
R574 B.n410 B.n409 163.367
R575 B.n410 B.n121 163.367
R576 B.n414 B.n121 163.367
R577 B.n415 B.n414 163.367
R578 B.n416 B.n415 163.367
R579 B.n416 B.n119 163.367
R580 B.n420 B.n119 163.367
R581 B.n421 B.n420 163.367
R582 B.n422 B.n421 163.367
R583 B.n422 B.n117 163.367
R584 B.n426 B.n117 163.367
R585 B.n428 B.n427 163.367
R586 B.n428 B.n115 163.367
R587 B.n432 B.n115 163.367
R588 B.n433 B.n432 163.367
R589 B.n434 B.n433 163.367
R590 B.n434 B.n113 163.367
R591 B.n438 B.n113 163.367
R592 B.n439 B.n438 163.367
R593 B.n440 B.n439 163.367
R594 B.n440 B.n111 163.367
R595 B.n444 B.n111 163.367
R596 B.n445 B.n444 163.367
R597 B.n446 B.n445 163.367
R598 B.n446 B.n109 163.367
R599 B.n450 B.n109 163.367
R600 B.n451 B.n450 163.367
R601 B.n452 B.n451 163.367
R602 B.n452 B.n107 163.367
R603 B.n456 B.n107 163.367
R604 B.n457 B.n456 163.367
R605 B.n458 B.n457 163.367
R606 B.n458 B.n105 163.367
R607 B.n462 B.n105 163.367
R608 B.n463 B.n462 163.367
R609 B.n464 B.n463 163.367
R610 B.n464 B.n103 163.367
R611 B.n468 B.n103 163.367
R612 B.n469 B.n468 163.367
R613 B.n470 B.n469 163.367
R614 B.n470 B.n101 163.367
R615 B.n474 B.n101 163.367
R616 B.n475 B.n474 163.367
R617 B.n476 B.n475 163.367
R618 B.n476 B.n99 163.367
R619 B.n480 B.n99 163.367
R620 B.n481 B.n480 163.367
R621 B.n482 B.n481 163.367
R622 B.n482 B.n97 163.367
R623 B.n486 B.n97 163.367
R624 B.n487 B.n486 163.367
R625 B.n488 B.n487 163.367
R626 B.n488 B.n95 163.367
R627 B.n492 B.n95 163.367
R628 B.n493 B.n492 163.367
R629 B.n494 B.n493 163.367
R630 B.n494 B.n93 163.367
R631 B.n498 B.n93 163.367
R632 B.n499 B.n498 163.367
R633 B.n500 B.n499 163.367
R634 B.n500 B.n91 163.367
R635 B.n504 B.n91 163.367
R636 B.n505 B.n504 163.367
R637 B.n506 B.n505 163.367
R638 B.n506 B.n89 163.367
R639 B.n510 B.n89 163.367
R640 B.n511 B.n510 163.367
R641 B.n512 B.n511 163.367
R642 B.n512 B.n87 163.367
R643 B.n516 B.n87 163.367
R644 B.n517 B.n516 163.367
R645 B.n518 B.n517 163.367
R646 B.n518 B.n85 163.367
R647 B.n522 B.n85 163.367
R648 B.n523 B.n522 163.367
R649 B.n524 B.n523 163.367
R650 B.n524 B.n83 163.367
R651 B.n708 B.n19 163.367
R652 B.n704 B.n19 163.367
R653 B.n704 B.n703 163.367
R654 B.n703 B.n702 163.367
R655 B.n702 B.n21 163.367
R656 B.n698 B.n21 163.367
R657 B.n698 B.n697 163.367
R658 B.n697 B.n696 163.367
R659 B.n696 B.n23 163.367
R660 B.n692 B.n23 163.367
R661 B.n692 B.n691 163.367
R662 B.n691 B.n690 163.367
R663 B.n690 B.n25 163.367
R664 B.n686 B.n25 163.367
R665 B.n686 B.n685 163.367
R666 B.n685 B.n684 163.367
R667 B.n684 B.n27 163.367
R668 B.n680 B.n27 163.367
R669 B.n680 B.n679 163.367
R670 B.n679 B.n678 163.367
R671 B.n678 B.n29 163.367
R672 B.n674 B.n29 163.367
R673 B.n674 B.n673 163.367
R674 B.n673 B.n672 163.367
R675 B.n672 B.n31 163.367
R676 B.n668 B.n31 163.367
R677 B.n668 B.n667 163.367
R678 B.n667 B.n666 163.367
R679 B.n666 B.n33 163.367
R680 B.n662 B.n33 163.367
R681 B.n662 B.n661 163.367
R682 B.n661 B.n660 163.367
R683 B.n660 B.n35 163.367
R684 B.n656 B.n35 163.367
R685 B.n656 B.n655 163.367
R686 B.n655 B.n654 163.367
R687 B.n654 B.n37 163.367
R688 B.n650 B.n37 163.367
R689 B.n650 B.n649 163.367
R690 B.n649 B.n648 163.367
R691 B.n648 B.n39 163.367
R692 B.n644 B.n39 163.367
R693 B.n644 B.n643 163.367
R694 B.n643 B.n642 163.367
R695 B.n642 B.n41 163.367
R696 B.n638 B.n41 163.367
R697 B.n638 B.n637 163.367
R698 B.n637 B.n636 163.367
R699 B.n636 B.n43 163.367
R700 B.n632 B.n43 163.367
R701 B.n632 B.n631 163.367
R702 B.n631 B.n630 163.367
R703 B.n630 B.n45 163.367
R704 B.n626 B.n45 163.367
R705 B.n626 B.n625 163.367
R706 B.n625 B.n49 163.367
R707 B.n621 B.n49 163.367
R708 B.n621 B.n620 163.367
R709 B.n620 B.n619 163.367
R710 B.n619 B.n51 163.367
R711 B.n615 B.n51 163.367
R712 B.n615 B.n614 163.367
R713 B.n614 B.n613 163.367
R714 B.n613 B.n53 163.367
R715 B.n608 B.n53 163.367
R716 B.n608 B.n607 163.367
R717 B.n607 B.n606 163.367
R718 B.n606 B.n57 163.367
R719 B.n602 B.n57 163.367
R720 B.n602 B.n601 163.367
R721 B.n601 B.n600 163.367
R722 B.n600 B.n59 163.367
R723 B.n596 B.n59 163.367
R724 B.n596 B.n595 163.367
R725 B.n595 B.n594 163.367
R726 B.n594 B.n61 163.367
R727 B.n590 B.n61 163.367
R728 B.n590 B.n589 163.367
R729 B.n589 B.n588 163.367
R730 B.n588 B.n63 163.367
R731 B.n584 B.n63 163.367
R732 B.n584 B.n583 163.367
R733 B.n583 B.n582 163.367
R734 B.n582 B.n65 163.367
R735 B.n578 B.n65 163.367
R736 B.n578 B.n577 163.367
R737 B.n577 B.n576 163.367
R738 B.n576 B.n67 163.367
R739 B.n572 B.n67 163.367
R740 B.n572 B.n571 163.367
R741 B.n571 B.n570 163.367
R742 B.n570 B.n69 163.367
R743 B.n566 B.n69 163.367
R744 B.n566 B.n565 163.367
R745 B.n565 B.n564 163.367
R746 B.n564 B.n71 163.367
R747 B.n560 B.n71 163.367
R748 B.n560 B.n559 163.367
R749 B.n559 B.n558 163.367
R750 B.n558 B.n73 163.367
R751 B.n554 B.n73 163.367
R752 B.n554 B.n553 163.367
R753 B.n553 B.n552 163.367
R754 B.n552 B.n75 163.367
R755 B.n548 B.n75 163.367
R756 B.n548 B.n547 163.367
R757 B.n547 B.n546 163.367
R758 B.n546 B.n77 163.367
R759 B.n542 B.n77 163.367
R760 B.n542 B.n541 163.367
R761 B.n541 B.n540 163.367
R762 B.n540 B.n79 163.367
R763 B.n536 B.n79 163.367
R764 B.n536 B.n535 163.367
R765 B.n535 B.n534 163.367
R766 B.n534 B.n81 163.367
R767 B.n530 B.n81 163.367
R768 B.n530 B.n529 163.367
R769 B.n529 B.n528 163.367
R770 B.n145 B.t4 112.362
R771 B.n55 B.t2 112.362
R772 B.n153 B.t7 112.341
R773 B.n47 B.t11 112.341
R774 B.n145 B.n144 82.8126
R775 B.n153 B.n152 82.8126
R776 B.n47 B.n46 82.8126
R777 B.n55 B.n54 82.8126
R778 B.n146 B.n145 59.5399
R779 B.n328 B.n153 59.5399
R780 B.n48 B.n47 59.5399
R781 B.n610 B.n55 59.5399
R782 B.n707 B.n18 35.1225
R783 B.n527 B.n526 35.1225
R784 B.n425 B.n116 35.1225
R785 B.n245 B.n244 35.1225
R786 B B.n759 18.0485
R787 B.n707 B.n706 10.6151
R788 B.n706 B.n705 10.6151
R789 B.n705 B.n20 10.6151
R790 B.n701 B.n20 10.6151
R791 B.n701 B.n700 10.6151
R792 B.n700 B.n699 10.6151
R793 B.n699 B.n22 10.6151
R794 B.n695 B.n22 10.6151
R795 B.n695 B.n694 10.6151
R796 B.n694 B.n693 10.6151
R797 B.n693 B.n24 10.6151
R798 B.n689 B.n24 10.6151
R799 B.n689 B.n688 10.6151
R800 B.n688 B.n687 10.6151
R801 B.n687 B.n26 10.6151
R802 B.n683 B.n26 10.6151
R803 B.n683 B.n682 10.6151
R804 B.n682 B.n681 10.6151
R805 B.n681 B.n28 10.6151
R806 B.n677 B.n28 10.6151
R807 B.n677 B.n676 10.6151
R808 B.n676 B.n675 10.6151
R809 B.n675 B.n30 10.6151
R810 B.n671 B.n30 10.6151
R811 B.n671 B.n670 10.6151
R812 B.n670 B.n669 10.6151
R813 B.n669 B.n32 10.6151
R814 B.n665 B.n32 10.6151
R815 B.n665 B.n664 10.6151
R816 B.n664 B.n663 10.6151
R817 B.n663 B.n34 10.6151
R818 B.n659 B.n34 10.6151
R819 B.n659 B.n658 10.6151
R820 B.n658 B.n657 10.6151
R821 B.n657 B.n36 10.6151
R822 B.n653 B.n36 10.6151
R823 B.n653 B.n652 10.6151
R824 B.n652 B.n651 10.6151
R825 B.n651 B.n38 10.6151
R826 B.n647 B.n38 10.6151
R827 B.n647 B.n646 10.6151
R828 B.n646 B.n645 10.6151
R829 B.n645 B.n40 10.6151
R830 B.n641 B.n40 10.6151
R831 B.n641 B.n640 10.6151
R832 B.n640 B.n639 10.6151
R833 B.n639 B.n42 10.6151
R834 B.n635 B.n42 10.6151
R835 B.n635 B.n634 10.6151
R836 B.n634 B.n633 10.6151
R837 B.n633 B.n44 10.6151
R838 B.n629 B.n44 10.6151
R839 B.n629 B.n628 10.6151
R840 B.n628 B.n627 10.6151
R841 B.n624 B.n623 10.6151
R842 B.n623 B.n622 10.6151
R843 B.n622 B.n50 10.6151
R844 B.n618 B.n50 10.6151
R845 B.n618 B.n617 10.6151
R846 B.n617 B.n616 10.6151
R847 B.n616 B.n52 10.6151
R848 B.n612 B.n52 10.6151
R849 B.n612 B.n611 10.6151
R850 B.n609 B.n56 10.6151
R851 B.n605 B.n56 10.6151
R852 B.n605 B.n604 10.6151
R853 B.n604 B.n603 10.6151
R854 B.n603 B.n58 10.6151
R855 B.n599 B.n58 10.6151
R856 B.n599 B.n598 10.6151
R857 B.n598 B.n597 10.6151
R858 B.n597 B.n60 10.6151
R859 B.n593 B.n60 10.6151
R860 B.n593 B.n592 10.6151
R861 B.n592 B.n591 10.6151
R862 B.n591 B.n62 10.6151
R863 B.n587 B.n62 10.6151
R864 B.n587 B.n586 10.6151
R865 B.n586 B.n585 10.6151
R866 B.n585 B.n64 10.6151
R867 B.n581 B.n64 10.6151
R868 B.n581 B.n580 10.6151
R869 B.n580 B.n579 10.6151
R870 B.n579 B.n66 10.6151
R871 B.n575 B.n66 10.6151
R872 B.n575 B.n574 10.6151
R873 B.n574 B.n573 10.6151
R874 B.n573 B.n68 10.6151
R875 B.n569 B.n68 10.6151
R876 B.n569 B.n568 10.6151
R877 B.n568 B.n567 10.6151
R878 B.n567 B.n70 10.6151
R879 B.n563 B.n70 10.6151
R880 B.n563 B.n562 10.6151
R881 B.n562 B.n561 10.6151
R882 B.n561 B.n72 10.6151
R883 B.n557 B.n72 10.6151
R884 B.n557 B.n556 10.6151
R885 B.n556 B.n555 10.6151
R886 B.n555 B.n74 10.6151
R887 B.n551 B.n74 10.6151
R888 B.n551 B.n550 10.6151
R889 B.n550 B.n549 10.6151
R890 B.n549 B.n76 10.6151
R891 B.n545 B.n76 10.6151
R892 B.n545 B.n544 10.6151
R893 B.n544 B.n543 10.6151
R894 B.n543 B.n78 10.6151
R895 B.n539 B.n78 10.6151
R896 B.n539 B.n538 10.6151
R897 B.n538 B.n537 10.6151
R898 B.n537 B.n80 10.6151
R899 B.n533 B.n80 10.6151
R900 B.n533 B.n532 10.6151
R901 B.n532 B.n531 10.6151
R902 B.n531 B.n82 10.6151
R903 B.n527 B.n82 10.6151
R904 B.n429 B.n116 10.6151
R905 B.n430 B.n429 10.6151
R906 B.n431 B.n430 10.6151
R907 B.n431 B.n114 10.6151
R908 B.n435 B.n114 10.6151
R909 B.n436 B.n435 10.6151
R910 B.n437 B.n436 10.6151
R911 B.n437 B.n112 10.6151
R912 B.n441 B.n112 10.6151
R913 B.n442 B.n441 10.6151
R914 B.n443 B.n442 10.6151
R915 B.n443 B.n110 10.6151
R916 B.n447 B.n110 10.6151
R917 B.n448 B.n447 10.6151
R918 B.n449 B.n448 10.6151
R919 B.n449 B.n108 10.6151
R920 B.n453 B.n108 10.6151
R921 B.n454 B.n453 10.6151
R922 B.n455 B.n454 10.6151
R923 B.n455 B.n106 10.6151
R924 B.n459 B.n106 10.6151
R925 B.n460 B.n459 10.6151
R926 B.n461 B.n460 10.6151
R927 B.n461 B.n104 10.6151
R928 B.n465 B.n104 10.6151
R929 B.n466 B.n465 10.6151
R930 B.n467 B.n466 10.6151
R931 B.n467 B.n102 10.6151
R932 B.n471 B.n102 10.6151
R933 B.n472 B.n471 10.6151
R934 B.n473 B.n472 10.6151
R935 B.n473 B.n100 10.6151
R936 B.n477 B.n100 10.6151
R937 B.n478 B.n477 10.6151
R938 B.n479 B.n478 10.6151
R939 B.n479 B.n98 10.6151
R940 B.n483 B.n98 10.6151
R941 B.n484 B.n483 10.6151
R942 B.n485 B.n484 10.6151
R943 B.n485 B.n96 10.6151
R944 B.n489 B.n96 10.6151
R945 B.n490 B.n489 10.6151
R946 B.n491 B.n490 10.6151
R947 B.n491 B.n94 10.6151
R948 B.n495 B.n94 10.6151
R949 B.n496 B.n495 10.6151
R950 B.n497 B.n496 10.6151
R951 B.n497 B.n92 10.6151
R952 B.n501 B.n92 10.6151
R953 B.n502 B.n501 10.6151
R954 B.n503 B.n502 10.6151
R955 B.n503 B.n90 10.6151
R956 B.n507 B.n90 10.6151
R957 B.n508 B.n507 10.6151
R958 B.n509 B.n508 10.6151
R959 B.n509 B.n88 10.6151
R960 B.n513 B.n88 10.6151
R961 B.n514 B.n513 10.6151
R962 B.n515 B.n514 10.6151
R963 B.n515 B.n86 10.6151
R964 B.n519 B.n86 10.6151
R965 B.n520 B.n519 10.6151
R966 B.n521 B.n520 10.6151
R967 B.n521 B.n84 10.6151
R968 B.n525 B.n84 10.6151
R969 B.n526 B.n525 10.6151
R970 B.n245 B.n180 10.6151
R971 B.n249 B.n180 10.6151
R972 B.n250 B.n249 10.6151
R973 B.n251 B.n250 10.6151
R974 B.n251 B.n178 10.6151
R975 B.n255 B.n178 10.6151
R976 B.n256 B.n255 10.6151
R977 B.n257 B.n256 10.6151
R978 B.n257 B.n176 10.6151
R979 B.n261 B.n176 10.6151
R980 B.n262 B.n261 10.6151
R981 B.n263 B.n262 10.6151
R982 B.n263 B.n174 10.6151
R983 B.n267 B.n174 10.6151
R984 B.n268 B.n267 10.6151
R985 B.n269 B.n268 10.6151
R986 B.n269 B.n172 10.6151
R987 B.n273 B.n172 10.6151
R988 B.n274 B.n273 10.6151
R989 B.n275 B.n274 10.6151
R990 B.n275 B.n170 10.6151
R991 B.n279 B.n170 10.6151
R992 B.n280 B.n279 10.6151
R993 B.n281 B.n280 10.6151
R994 B.n281 B.n168 10.6151
R995 B.n285 B.n168 10.6151
R996 B.n286 B.n285 10.6151
R997 B.n287 B.n286 10.6151
R998 B.n287 B.n166 10.6151
R999 B.n291 B.n166 10.6151
R1000 B.n292 B.n291 10.6151
R1001 B.n293 B.n292 10.6151
R1002 B.n293 B.n164 10.6151
R1003 B.n297 B.n164 10.6151
R1004 B.n298 B.n297 10.6151
R1005 B.n299 B.n298 10.6151
R1006 B.n299 B.n162 10.6151
R1007 B.n303 B.n162 10.6151
R1008 B.n304 B.n303 10.6151
R1009 B.n305 B.n304 10.6151
R1010 B.n305 B.n160 10.6151
R1011 B.n309 B.n160 10.6151
R1012 B.n310 B.n309 10.6151
R1013 B.n311 B.n310 10.6151
R1014 B.n311 B.n158 10.6151
R1015 B.n315 B.n158 10.6151
R1016 B.n316 B.n315 10.6151
R1017 B.n317 B.n316 10.6151
R1018 B.n317 B.n156 10.6151
R1019 B.n321 B.n156 10.6151
R1020 B.n322 B.n321 10.6151
R1021 B.n323 B.n322 10.6151
R1022 B.n323 B.n154 10.6151
R1023 B.n327 B.n154 10.6151
R1024 B.n330 B.n329 10.6151
R1025 B.n330 B.n150 10.6151
R1026 B.n334 B.n150 10.6151
R1027 B.n335 B.n334 10.6151
R1028 B.n336 B.n335 10.6151
R1029 B.n336 B.n148 10.6151
R1030 B.n340 B.n148 10.6151
R1031 B.n341 B.n340 10.6151
R1032 B.n342 B.n341 10.6151
R1033 B.n346 B.n345 10.6151
R1034 B.n347 B.n346 10.6151
R1035 B.n347 B.n142 10.6151
R1036 B.n351 B.n142 10.6151
R1037 B.n352 B.n351 10.6151
R1038 B.n353 B.n352 10.6151
R1039 B.n353 B.n140 10.6151
R1040 B.n357 B.n140 10.6151
R1041 B.n358 B.n357 10.6151
R1042 B.n359 B.n358 10.6151
R1043 B.n359 B.n138 10.6151
R1044 B.n363 B.n138 10.6151
R1045 B.n364 B.n363 10.6151
R1046 B.n365 B.n364 10.6151
R1047 B.n365 B.n136 10.6151
R1048 B.n369 B.n136 10.6151
R1049 B.n370 B.n369 10.6151
R1050 B.n371 B.n370 10.6151
R1051 B.n371 B.n134 10.6151
R1052 B.n375 B.n134 10.6151
R1053 B.n376 B.n375 10.6151
R1054 B.n377 B.n376 10.6151
R1055 B.n377 B.n132 10.6151
R1056 B.n381 B.n132 10.6151
R1057 B.n382 B.n381 10.6151
R1058 B.n383 B.n382 10.6151
R1059 B.n383 B.n130 10.6151
R1060 B.n387 B.n130 10.6151
R1061 B.n388 B.n387 10.6151
R1062 B.n389 B.n388 10.6151
R1063 B.n389 B.n128 10.6151
R1064 B.n393 B.n128 10.6151
R1065 B.n394 B.n393 10.6151
R1066 B.n395 B.n394 10.6151
R1067 B.n395 B.n126 10.6151
R1068 B.n399 B.n126 10.6151
R1069 B.n400 B.n399 10.6151
R1070 B.n401 B.n400 10.6151
R1071 B.n401 B.n124 10.6151
R1072 B.n405 B.n124 10.6151
R1073 B.n406 B.n405 10.6151
R1074 B.n407 B.n406 10.6151
R1075 B.n407 B.n122 10.6151
R1076 B.n411 B.n122 10.6151
R1077 B.n412 B.n411 10.6151
R1078 B.n413 B.n412 10.6151
R1079 B.n413 B.n120 10.6151
R1080 B.n417 B.n120 10.6151
R1081 B.n418 B.n417 10.6151
R1082 B.n419 B.n418 10.6151
R1083 B.n419 B.n118 10.6151
R1084 B.n423 B.n118 10.6151
R1085 B.n424 B.n423 10.6151
R1086 B.n425 B.n424 10.6151
R1087 B.n244 B.n243 10.6151
R1088 B.n243 B.n182 10.6151
R1089 B.n239 B.n182 10.6151
R1090 B.n239 B.n238 10.6151
R1091 B.n238 B.n237 10.6151
R1092 B.n237 B.n184 10.6151
R1093 B.n233 B.n184 10.6151
R1094 B.n233 B.n232 10.6151
R1095 B.n232 B.n231 10.6151
R1096 B.n231 B.n186 10.6151
R1097 B.n227 B.n186 10.6151
R1098 B.n227 B.n226 10.6151
R1099 B.n226 B.n225 10.6151
R1100 B.n225 B.n188 10.6151
R1101 B.n221 B.n188 10.6151
R1102 B.n221 B.n220 10.6151
R1103 B.n220 B.n219 10.6151
R1104 B.n219 B.n190 10.6151
R1105 B.n215 B.n190 10.6151
R1106 B.n215 B.n214 10.6151
R1107 B.n214 B.n213 10.6151
R1108 B.n213 B.n192 10.6151
R1109 B.n209 B.n192 10.6151
R1110 B.n209 B.n208 10.6151
R1111 B.n208 B.n207 10.6151
R1112 B.n207 B.n194 10.6151
R1113 B.n203 B.n194 10.6151
R1114 B.n203 B.n202 10.6151
R1115 B.n202 B.n201 10.6151
R1116 B.n201 B.n196 10.6151
R1117 B.n197 B.n196 10.6151
R1118 B.n197 B.n0 10.6151
R1119 B.n755 B.n1 10.6151
R1120 B.n755 B.n754 10.6151
R1121 B.n754 B.n753 10.6151
R1122 B.n753 B.n4 10.6151
R1123 B.n749 B.n4 10.6151
R1124 B.n749 B.n748 10.6151
R1125 B.n748 B.n747 10.6151
R1126 B.n747 B.n6 10.6151
R1127 B.n743 B.n6 10.6151
R1128 B.n743 B.n742 10.6151
R1129 B.n742 B.n741 10.6151
R1130 B.n741 B.n8 10.6151
R1131 B.n737 B.n8 10.6151
R1132 B.n737 B.n736 10.6151
R1133 B.n736 B.n735 10.6151
R1134 B.n735 B.n10 10.6151
R1135 B.n731 B.n10 10.6151
R1136 B.n731 B.n730 10.6151
R1137 B.n730 B.n729 10.6151
R1138 B.n729 B.n12 10.6151
R1139 B.n725 B.n12 10.6151
R1140 B.n725 B.n724 10.6151
R1141 B.n724 B.n723 10.6151
R1142 B.n723 B.n14 10.6151
R1143 B.n719 B.n14 10.6151
R1144 B.n719 B.n718 10.6151
R1145 B.n718 B.n717 10.6151
R1146 B.n717 B.n16 10.6151
R1147 B.n713 B.n16 10.6151
R1148 B.n713 B.n712 10.6151
R1149 B.n712 B.n711 10.6151
R1150 B.n711 B.n18 10.6151
R1151 B.n627 B.n48 9.36635
R1152 B.n610 B.n609 9.36635
R1153 B.n328 B.n327 9.36635
R1154 B.n345 B.n146 9.36635
R1155 B.n759 B.n0 2.81026
R1156 B.n759 B.n1 2.81026
R1157 B.n624 B.n48 1.24928
R1158 B.n611 B.n610 1.24928
R1159 B.n329 B.n328 1.24928
R1160 B.n342 B.n146 1.24928
R1161 VP.n0 VP.t1 188.476
R1162 VP.n0 VP.t0 136.76
R1163 VP VP.n0 0.621237
R1164 VDD1 VDD1.t1 122.034
R1165 VDD1 VDD1.t0 76.2091
C0 VP VDD2 0.388723f
C1 VN VDD1 0.148738f
C2 VN VDD2 3.96476f
C3 B w_n2678_n4294# 11.5547f
C4 VP w_n2678_n4294# 4.25452f
C5 VTAIL VDD1 6.49677f
C6 VTAIL VDD2 6.55672f
C7 VN w_n2678_n4294# 3.91051f
C8 VP B 1.90038f
C9 VDD1 VDD2 0.826086f
C10 VN B 1.32943f
C11 VP VN 6.94194f
C12 VTAIL w_n2678_n4294# 3.39999f
C13 VTAIL B 5.249741f
C14 VDD1 w_n2678_n4294# 2.24252f
C15 VTAIL VP 3.50422f
C16 VDD2 w_n2678_n4294# 2.28488f
C17 VTAIL VN 3.48904f
C18 VDD1 B 2.25583f
C19 B VDD2 2.29796f
C20 VP VDD1 4.20307f
C21 VDD2 VSUBS 1.240964f
C22 VDD1 VSUBS 7.181981f
C23 VTAIL VSUBS 1.320167f
C24 VN VSUBS 9.13893f
C25 VP VSUBS 2.243589f
C26 B VSUBS 5.283687f
C27 w_n2678_n4294# VSUBS 0.140788p
C28 VDD1.t0 VSUBS 4.09046f
C29 VDD1.t1 VSUBS 5.22857f
C30 VP.t1 VSUBS 6.8632f
C31 VP.t0 VSUBS 5.88886f
C32 VP.n0 VSUBS 6.01609f
C33 B.n0 VSUBS 0.003975f
C34 B.n1 VSUBS 0.003975f
C35 B.n2 VSUBS 0.006285f
C36 B.n3 VSUBS 0.006285f
C37 B.n4 VSUBS 0.006285f
C38 B.n5 VSUBS 0.006285f
C39 B.n6 VSUBS 0.006285f
C40 B.n7 VSUBS 0.006285f
C41 B.n8 VSUBS 0.006285f
C42 B.n9 VSUBS 0.006285f
C43 B.n10 VSUBS 0.006285f
C44 B.n11 VSUBS 0.006285f
C45 B.n12 VSUBS 0.006285f
C46 B.n13 VSUBS 0.006285f
C47 B.n14 VSUBS 0.006285f
C48 B.n15 VSUBS 0.006285f
C49 B.n16 VSUBS 0.006285f
C50 B.n17 VSUBS 0.006285f
C51 B.n18 VSUBS 0.01499f
C52 B.n19 VSUBS 0.006285f
C53 B.n20 VSUBS 0.006285f
C54 B.n21 VSUBS 0.006285f
C55 B.n22 VSUBS 0.006285f
C56 B.n23 VSUBS 0.006285f
C57 B.n24 VSUBS 0.006285f
C58 B.n25 VSUBS 0.006285f
C59 B.n26 VSUBS 0.006285f
C60 B.n27 VSUBS 0.006285f
C61 B.n28 VSUBS 0.006285f
C62 B.n29 VSUBS 0.006285f
C63 B.n30 VSUBS 0.006285f
C64 B.n31 VSUBS 0.006285f
C65 B.n32 VSUBS 0.006285f
C66 B.n33 VSUBS 0.006285f
C67 B.n34 VSUBS 0.006285f
C68 B.n35 VSUBS 0.006285f
C69 B.n36 VSUBS 0.006285f
C70 B.n37 VSUBS 0.006285f
C71 B.n38 VSUBS 0.006285f
C72 B.n39 VSUBS 0.006285f
C73 B.n40 VSUBS 0.006285f
C74 B.n41 VSUBS 0.006285f
C75 B.n42 VSUBS 0.006285f
C76 B.n43 VSUBS 0.006285f
C77 B.n44 VSUBS 0.006285f
C78 B.n45 VSUBS 0.006285f
C79 B.t11 VSUBS 0.501228f
C80 B.t10 VSUBS 0.526987f
C81 B.t9 VSUBS 2.70015f
C82 B.n46 VSUBS 0.325769f
C83 B.n47 VSUBS 0.069667f
C84 B.n48 VSUBS 0.014562f
C85 B.n49 VSUBS 0.006285f
C86 B.n50 VSUBS 0.006285f
C87 B.n51 VSUBS 0.006285f
C88 B.n52 VSUBS 0.006285f
C89 B.n53 VSUBS 0.006285f
C90 B.t2 VSUBS 0.501212f
C91 B.t1 VSUBS 0.526975f
C92 B.t0 VSUBS 2.70015f
C93 B.n54 VSUBS 0.325781f
C94 B.n55 VSUBS 0.069683f
C95 B.n56 VSUBS 0.006285f
C96 B.n57 VSUBS 0.006285f
C97 B.n58 VSUBS 0.006285f
C98 B.n59 VSUBS 0.006285f
C99 B.n60 VSUBS 0.006285f
C100 B.n61 VSUBS 0.006285f
C101 B.n62 VSUBS 0.006285f
C102 B.n63 VSUBS 0.006285f
C103 B.n64 VSUBS 0.006285f
C104 B.n65 VSUBS 0.006285f
C105 B.n66 VSUBS 0.006285f
C106 B.n67 VSUBS 0.006285f
C107 B.n68 VSUBS 0.006285f
C108 B.n69 VSUBS 0.006285f
C109 B.n70 VSUBS 0.006285f
C110 B.n71 VSUBS 0.006285f
C111 B.n72 VSUBS 0.006285f
C112 B.n73 VSUBS 0.006285f
C113 B.n74 VSUBS 0.006285f
C114 B.n75 VSUBS 0.006285f
C115 B.n76 VSUBS 0.006285f
C116 B.n77 VSUBS 0.006285f
C117 B.n78 VSUBS 0.006285f
C118 B.n79 VSUBS 0.006285f
C119 B.n80 VSUBS 0.006285f
C120 B.n81 VSUBS 0.006285f
C121 B.n82 VSUBS 0.006285f
C122 B.n83 VSUBS 0.01499f
C123 B.n84 VSUBS 0.006285f
C124 B.n85 VSUBS 0.006285f
C125 B.n86 VSUBS 0.006285f
C126 B.n87 VSUBS 0.006285f
C127 B.n88 VSUBS 0.006285f
C128 B.n89 VSUBS 0.006285f
C129 B.n90 VSUBS 0.006285f
C130 B.n91 VSUBS 0.006285f
C131 B.n92 VSUBS 0.006285f
C132 B.n93 VSUBS 0.006285f
C133 B.n94 VSUBS 0.006285f
C134 B.n95 VSUBS 0.006285f
C135 B.n96 VSUBS 0.006285f
C136 B.n97 VSUBS 0.006285f
C137 B.n98 VSUBS 0.006285f
C138 B.n99 VSUBS 0.006285f
C139 B.n100 VSUBS 0.006285f
C140 B.n101 VSUBS 0.006285f
C141 B.n102 VSUBS 0.006285f
C142 B.n103 VSUBS 0.006285f
C143 B.n104 VSUBS 0.006285f
C144 B.n105 VSUBS 0.006285f
C145 B.n106 VSUBS 0.006285f
C146 B.n107 VSUBS 0.006285f
C147 B.n108 VSUBS 0.006285f
C148 B.n109 VSUBS 0.006285f
C149 B.n110 VSUBS 0.006285f
C150 B.n111 VSUBS 0.006285f
C151 B.n112 VSUBS 0.006285f
C152 B.n113 VSUBS 0.006285f
C153 B.n114 VSUBS 0.006285f
C154 B.n115 VSUBS 0.006285f
C155 B.n116 VSUBS 0.01499f
C156 B.n117 VSUBS 0.006285f
C157 B.n118 VSUBS 0.006285f
C158 B.n119 VSUBS 0.006285f
C159 B.n120 VSUBS 0.006285f
C160 B.n121 VSUBS 0.006285f
C161 B.n122 VSUBS 0.006285f
C162 B.n123 VSUBS 0.006285f
C163 B.n124 VSUBS 0.006285f
C164 B.n125 VSUBS 0.006285f
C165 B.n126 VSUBS 0.006285f
C166 B.n127 VSUBS 0.006285f
C167 B.n128 VSUBS 0.006285f
C168 B.n129 VSUBS 0.006285f
C169 B.n130 VSUBS 0.006285f
C170 B.n131 VSUBS 0.006285f
C171 B.n132 VSUBS 0.006285f
C172 B.n133 VSUBS 0.006285f
C173 B.n134 VSUBS 0.006285f
C174 B.n135 VSUBS 0.006285f
C175 B.n136 VSUBS 0.006285f
C176 B.n137 VSUBS 0.006285f
C177 B.n138 VSUBS 0.006285f
C178 B.n139 VSUBS 0.006285f
C179 B.n140 VSUBS 0.006285f
C180 B.n141 VSUBS 0.006285f
C181 B.n142 VSUBS 0.006285f
C182 B.n143 VSUBS 0.006285f
C183 B.t4 VSUBS 0.501212f
C184 B.t5 VSUBS 0.526975f
C185 B.t3 VSUBS 2.70015f
C186 B.n144 VSUBS 0.325781f
C187 B.n145 VSUBS 0.069683f
C188 B.n146 VSUBS 0.014562f
C189 B.n147 VSUBS 0.006285f
C190 B.n148 VSUBS 0.006285f
C191 B.n149 VSUBS 0.006285f
C192 B.n150 VSUBS 0.006285f
C193 B.n151 VSUBS 0.006285f
C194 B.t7 VSUBS 0.501228f
C195 B.t8 VSUBS 0.526987f
C196 B.t6 VSUBS 2.70015f
C197 B.n152 VSUBS 0.325769f
C198 B.n153 VSUBS 0.069667f
C199 B.n154 VSUBS 0.006285f
C200 B.n155 VSUBS 0.006285f
C201 B.n156 VSUBS 0.006285f
C202 B.n157 VSUBS 0.006285f
C203 B.n158 VSUBS 0.006285f
C204 B.n159 VSUBS 0.006285f
C205 B.n160 VSUBS 0.006285f
C206 B.n161 VSUBS 0.006285f
C207 B.n162 VSUBS 0.006285f
C208 B.n163 VSUBS 0.006285f
C209 B.n164 VSUBS 0.006285f
C210 B.n165 VSUBS 0.006285f
C211 B.n166 VSUBS 0.006285f
C212 B.n167 VSUBS 0.006285f
C213 B.n168 VSUBS 0.006285f
C214 B.n169 VSUBS 0.006285f
C215 B.n170 VSUBS 0.006285f
C216 B.n171 VSUBS 0.006285f
C217 B.n172 VSUBS 0.006285f
C218 B.n173 VSUBS 0.006285f
C219 B.n174 VSUBS 0.006285f
C220 B.n175 VSUBS 0.006285f
C221 B.n176 VSUBS 0.006285f
C222 B.n177 VSUBS 0.006285f
C223 B.n178 VSUBS 0.006285f
C224 B.n179 VSUBS 0.006285f
C225 B.n180 VSUBS 0.006285f
C226 B.n181 VSUBS 0.01499f
C227 B.n182 VSUBS 0.006285f
C228 B.n183 VSUBS 0.006285f
C229 B.n184 VSUBS 0.006285f
C230 B.n185 VSUBS 0.006285f
C231 B.n186 VSUBS 0.006285f
C232 B.n187 VSUBS 0.006285f
C233 B.n188 VSUBS 0.006285f
C234 B.n189 VSUBS 0.006285f
C235 B.n190 VSUBS 0.006285f
C236 B.n191 VSUBS 0.006285f
C237 B.n192 VSUBS 0.006285f
C238 B.n193 VSUBS 0.006285f
C239 B.n194 VSUBS 0.006285f
C240 B.n195 VSUBS 0.006285f
C241 B.n196 VSUBS 0.006285f
C242 B.n197 VSUBS 0.006285f
C243 B.n198 VSUBS 0.006285f
C244 B.n199 VSUBS 0.006285f
C245 B.n200 VSUBS 0.006285f
C246 B.n201 VSUBS 0.006285f
C247 B.n202 VSUBS 0.006285f
C248 B.n203 VSUBS 0.006285f
C249 B.n204 VSUBS 0.006285f
C250 B.n205 VSUBS 0.006285f
C251 B.n206 VSUBS 0.006285f
C252 B.n207 VSUBS 0.006285f
C253 B.n208 VSUBS 0.006285f
C254 B.n209 VSUBS 0.006285f
C255 B.n210 VSUBS 0.006285f
C256 B.n211 VSUBS 0.006285f
C257 B.n212 VSUBS 0.006285f
C258 B.n213 VSUBS 0.006285f
C259 B.n214 VSUBS 0.006285f
C260 B.n215 VSUBS 0.006285f
C261 B.n216 VSUBS 0.006285f
C262 B.n217 VSUBS 0.006285f
C263 B.n218 VSUBS 0.006285f
C264 B.n219 VSUBS 0.006285f
C265 B.n220 VSUBS 0.006285f
C266 B.n221 VSUBS 0.006285f
C267 B.n222 VSUBS 0.006285f
C268 B.n223 VSUBS 0.006285f
C269 B.n224 VSUBS 0.006285f
C270 B.n225 VSUBS 0.006285f
C271 B.n226 VSUBS 0.006285f
C272 B.n227 VSUBS 0.006285f
C273 B.n228 VSUBS 0.006285f
C274 B.n229 VSUBS 0.006285f
C275 B.n230 VSUBS 0.006285f
C276 B.n231 VSUBS 0.006285f
C277 B.n232 VSUBS 0.006285f
C278 B.n233 VSUBS 0.006285f
C279 B.n234 VSUBS 0.006285f
C280 B.n235 VSUBS 0.006285f
C281 B.n236 VSUBS 0.006285f
C282 B.n237 VSUBS 0.006285f
C283 B.n238 VSUBS 0.006285f
C284 B.n239 VSUBS 0.006285f
C285 B.n240 VSUBS 0.006285f
C286 B.n241 VSUBS 0.006285f
C287 B.n242 VSUBS 0.006285f
C288 B.n243 VSUBS 0.006285f
C289 B.n244 VSUBS 0.01499f
C290 B.n245 VSUBS 0.015882f
C291 B.n246 VSUBS 0.015882f
C292 B.n247 VSUBS 0.006285f
C293 B.n248 VSUBS 0.006285f
C294 B.n249 VSUBS 0.006285f
C295 B.n250 VSUBS 0.006285f
C296 B.n251 VSUBS 0.006285f
C297 B.n252 VSUBS 0.006285f
C298 B.n253 VSUBS 0.006285f
C299 B.n254 VSUBS 0.006285f
C300 B.n255 VSUBS 0.006285f
C301 B.n256 VSUBS 0.006285f
C302 B.n257 VSUBS 0.006285f
C303 B.n258 VSUBS 0.006285f
C304 B.n259 VSUBS 0.006285f
C305 B.n260 VSUBS 0.006285f
C306 B.n261 VSUBS 0.006285f
C307 B.n262 VSUBS 0.006285f
C308 B.n263 VSUBS 0.006285f
C309 B.n264 VSUBS 0.006285f
C310 B.n265 VSUBS 0.006285f
C311 B.n266 VSUBS 0.006285f
C312 B.n267 VSUBS 0.006285f
C313 B.n268 VSUBS 0.006285f
C314 B.n269 VSUBS 0.006285f
C315 B.n270 VSUBS 0.006285f
C316 B.n271 VSUBS 0.006285f
C317 B.n272 VSUBS 0.006285f
C318 B.n273 VSUBS 0.006285f
C319 B.n274 VSUBS 0.006285f
C320 B.n275 VSUBS 0.006285f
C321 B.n276 VSUBS 0.006285f
C322 B.n277 VSUBS 0.006285f
C323 B.n278 VSUBS 0.006285f
C324 B.n279 VSUBS 0.006285f
C325 B.n280 VSUBS 0.006285f
C326 B.n281 VSUBS 0.006285f
C327 B.n282 VSUBS 0.006285f
C328 B.n283 VSUBS 0.006285f
C329 B.n284 VSUBS 0.006285f
C330 B.n285 VSUBS 0.006285f
C331 B.n286 VSUBS 0.006285f
C332 B.n287 VSUBS 0.006285f
C333 B.n288 VSUBS 0.006285f
C334 B.n289 VSUBS 0.006285f
C335 B.n290 VSUBS 0.006285f
C336 B.n291 VSUBS 0.006285f
C337 B.n292 VSUBS 0.006285f
C338 B.n293 VSUBS 0.006285f
C339 B.n294 VSUBS 0.006285f
C340 B.n295 VSUBS 0.006285f
C341 B.n296 VSUBS 0.006285f
C342 B.n297 VSUBS 0.006285f
C343 B.n298 VSUBS 0.006285f
C344 B.n299 VSUBS 0.006285f
C345 B.n300 VSUBS 0.006285f
C346 B.n301 VSUBS 0.006285f
C347 B.n302 VSUBS 0.006285f
C348 B.n303 VSUBS 0.006285f
C349 B.n304 VSUBS 0.006285f
C350 B.n305 VSUBS 0.006285f
C351 B.n306 VSUBS 0.006285f
C352 B.n307 VSUBS 0.006285f
C353 B.n308 VSUBS 0.006285f
C354 B.n309 VSUBS 0.006285f
C355 B.n310 VSUBS 0.006285f
C356 B.n311 VSUBS 0.006285f
C357 B.n312 VSUBS 0.006285f
C358 B.n313 VSUBS 0.006285f
C359 B.n314 VSUBS 0.006285f
C360 B.n315 VSUBS 0.006285f
C361 B.n316 VSUBS 0.006285f
C362 B.n317 VSUBS 0.006285f
C363 B.n318 VSUBS 0.006285f
C364 B.n319 VSUBS 0.006285f
C365 B.n320 VSUBS 0.006285f
C366 B.n321 VSUBS 0.006285f
C367 B.n322 VSUBS 0.006285f
C368 B.n323 VSUBS 0.006285f
C369 B.n324 VSUBS 0.006285f
C370 B.n325 VSUBS 0.006285f
C371 B.n326 VSUBS 0.006285f
C372 B.n327 VSUBS 0.005916f
C373 B.n328 VSUBS 0.014562f
C374 B.n329 VSUBS 0.003512f
C375 B.n330 VSUBS 0.006285f
C376 B.n331 VSUBS 0.006285f
C377 B.n332 VSUBS 0.006285f
C378 B.n333 VSUBS 0.006285f
C379 B.n334 VSUBS 0.006285f
C380 B.n335 VSUBS 0.006285f
C381 B.n336 VSUBS 0.006285f
C382 B.n337 VSUBS 0.006285f
C383 B.n338 VSUBS 0.006285f
C384 B.n339 VSUBS 0.006285f
C385 B.n340 VSUBS 0.006285f
C386 B.n341 VSUBS 0.006285f
C387 B.n342 VSUBS 0.003512f
C388 B.n343 VSUBS 0.006285f
C389 B.n344 VSUBS 0.006285f
C390 B.n345 VSUBS 0.005916f
C391 B.n346 VSUBS 0.006285f
C392 B.n347 VSUBS 0.006285f
C393 B.n348 VSUBS 0.006285f
C394 B.n349 VSUBS 0.006285f
C395 B.n350 VSUBS 0.006285f
C396 B.n351 VSUBS 0.006285f
C397 B.n352 VSUBS 0.006285f
C398 B.n353 VSUBS 0.006285f
C399 B.n354 VSUBS 0.006285f
C400 B.n355 VSUBS 0.006285f
C401 B.n356 VSUBS 0.006285f
C402 B.n357 VSUBS 0.006285f
C403 B.n358 VSUBS 0.006285f
C404 B.n359 VSUBS 0.006285f
C405 B.n360 VSUBS 0.006285f
C406 B.n361 VSUBS 0.006285f
C407 B.n362 VSUBS 0.006285f
C408 B.n363 VSUBS 0.006285f
C409 B.n364 VSUBS 0.006285f
C410 B.n365 VSUBS 0.006285f
C411 B.n366 VSUBS 0.006285f
C412 B.n367 VSUBS 0.006285f
C413 B.n368 VSUBS 0.006285f
C414 B.n369 VSUBS 0.006285f
C415 B.n370 VSUBS 0.006285f
C416 B.n371 VSUBS 0.006285f
C417 B.n372 VSUBS 0.006285f
C418 B.n373 VSUBS 0.006285f
C419 B.n374 VSUBS 0.006285f
C420 B.n375 VSUBS 0.006285f
C421 B.n376 VSUBS 0.006285f
C422 B.n377 VSUBS 0.006285f
C423 B.n378 VSUBS 0.006285f
C424 B.n379 VSUBS 0.006285f
C425 B.n380 VSUBS 0.006285f
C426 B.n381 VSUBS 0.006285f
C427 B.n382 VSUBS 0.006285f
C428 B.n383 VSUBS 0.006285f
C429 B.n384 VSUBS 0.006285f
C430 B.n385 VSUBS 0.006285f
C431 B.n386 VSUBS 0.006285f
C432 B.n387 VSUBS 0.006285f
C433 B.n388 VSUBS 0.006285f
C434 B.n389 VSUBS 0.006285f
C435 B.n390 VSUBS 0.006285f
C436 B.n391 VSUBS 0.006285f
C437 B.n392 VSUBS 0.006285f
C438 B.n393 VSUBS 0.006285f
C439 B.n394 VSUBS 0.006285f
C440 B.n395 VSUBS 0.006285f
C441 B.n396 VSUBS 0.006285f
C442 B.n397 VSUBS 0.006285f
C443 B.n398 VSUBS 0.006285f
C444 B.n399 VSUBS 0.006285f
C445 B.n400 VSUBS 0.006285f
C446 B.n401 VSUBS 0.006285f
C447 B.n402 VSUBS 0.006285f
C448 B.n403 VSUBS 0.006285f
C449 B.n404 VSUBS 0.006285f
C450 B.n405 VSUBS 0.006285f
C451 B.n406 VSUBS 0.006285f
C452 B.n407 VSUBS 0.006285f
C453 B.n408 VSUBS 0.006285f
C454 B.n409 VSUBS 0.006285f
C455 B.n410 VSUBS 0.006285f
C456 B.n411 VSUBS 0.006285f
C457 B.n412 VSUBS 0.006285f
C458 B.n413 VSUBS 0.006285f
C459 B.n414 VSUBS 0.006285f
C460 B.n415 VSUBS 0.006285f
C461 B.n416 VSUBS 0.006285f
C462 B.n417 VSUBS 0.006285f
C463 B.n418 VSUBS 0.006285f
C464 B.n419 VSUBS 0.006285f
C465 B.n420 VSUBS 0.006285f
C466 B.n421 VSUBS 0.006285f
C467 B.n422 VSUBS 0.006285f
C468 B.n423 VSUBS 0.006285f
C469 B.n424 VSUBS 0.006285f
C470 B.n425 VSUBS 0.015882f
C471 B.n426 VSUBS 0.015882f
C472 B.n427 VSUBS 0.01499f
C473 B.n428 VSUBS 0.006285f
C474 B.n429 VSUBS 0.006285f
C475 B.n430 VSUBS 0.006285f
C476 B.n431 VSUBS 0.006285f
C477 B.n432 VSUBS 0.006285f
C478 B.n433 VSUBS 0.006285f
C479 B.n434 VSUBS 0.006285f
C480 B.n435 VSUBS 0.006285f
C481 B.n436 VSUBS 0.006285f
C482 B.n437 VSUBS 0.006285f
C483 B.n438 VSUBS 0.006285f
C484 B.n439 VSUBS 0.006285f
C485 B.n440 VSUBS 0.006285f
C486 B.n441 VSUBS 0.006285f
C487 B.n442 VSUBS 0.006285f
C488 B.n443 VSUBS 0.006285f
C489 B.n444 VSUBS 0.006285f
C490 B.n445 VSUBS 0.006285f
C491 B.n446 VSUBS 0.006285f
C492 B.n447 VSUBS 0.006285f
C493 B.n448 VSUBS 0.006285f
C494 B.n449 VSUBS 0.006285f
C495 B.n450 VSUBS 0.006285f
C496 B.n451 VSUBS 0.006285f
C497 B.n452 VSUBS 0.006285f
C498 B.n453 VSUBS 0.006285f
C499 B.n454 VSUBS 0.006285f
C500 B.n455 VSUBS 0.006285f
C501 B.n456 VSUBS 0.006285f
C502 B.n457 VSUBS 0.006285f
C503 B.n458 VSUBS 0.006285f
C504 B.n459 VSUBS 0.006285f
C505 B.n460 VSUBS 0.006285f
C506 B.n461 VSUBS 0.006285f
C507 B.n462 VSUBS 0.006285f
C508 B.n463 VSUBS 0.006285f
C509 B.n464 VSUBS 0.006285f
C510 B.n465 VSUBS 0.006285f
C511 B.n466 VSUBS 0.006285f
C512 B.n467 VSUBS 0.006285f
C513 B.n468 VSUBS 0.006285f
C514 B.n469 VSUBS 0.006285f
C515 B.n470 VSUBS 0.006285f
C516 B.n471 VSUBS 0.006285f
C517 B.n472 VSUBS 0.006285f
C518 B.n473 VSUBS 0.006285f
C519 B.n474 VSUBS 0.006285f
C520 B.n475 VSUBS 0.006285f
C521 B.n476 VSUBS 0.006285f
C522 B.n477 VSUBS 0.006285f
C523 B.n478 VSUBS 0.006285f
C524 B.n479 VSUBS 0.006285f
C525 B.n480 VSUBS 0.006285f
C526 B.n481 VSUBS 0.006285f
C527 B.n482 VSUBS 0.006285f
C528 B.n483 VSUBS 0.006285f
C529 B.n484 VSUBS 0.006285f
C530 B.n485 VSUBS 0.006285f
C531 B.n486 VSUBS 0.006285f
C532 B.n487 VSUBS 0.006285f
C533 B.n488 VSUBS 0.006285f
C534 B.n489 VSUBS 0.006285f
C535 B.n490 VSUBS 0.006285f
C536 B.n491 VSUBS 0.006285f
C537 B.n492 VSUBS 0.006285f
C538 B.n493 VSUBS 0.006285f
C539 B.n494 VSUBS 0.006285f
C540 B.n495 VSUBS 0.006285f
C541 B.n496 VSUBS 0.006285f
C542 B.n497 VSUBS 0.006285f
C543 B.n498 VSUBS 0.006285f
C544 B.n499 VSUBS 0.006285f
C545 B.n500 VSUBS 0.006285f
C546 B.n501 VSUBS 0.006285f
C547 B.n502 VSUBS 0.006285f
C548 B.n503 VSUBS 0.006285f
C549 B.n504 VSUBS 0.006285f
C550 B.n505 VSUBS 0.006285f
C551 B.n506 VSUBS 0.006285f
C552 B.n507 VSUBS 0.006285f
C553 B.n508 VSUBS 0.006285f
C554 B.n509 VSUBS 0.006285f
C555 B.n510 VSUBS 0.006285f
C556 B.n511 VSUBS 0.006285f
C557 B.n512 VSUBS 0.006285f
C558 B.n513 VSUBS 0.006285f
C559 B.n514 VSUBS 0.006285f
C560 B.n515 VSUBS 0.006285f
C561 B.n516 VSUBS 0.006285f
C562 B.n517 VSUBS 0.006285f
C563 B.n518 VSUBS 0.006285f
C564 B.n519 VSUBS 0.006285f
C565 B.n520 VSUBS 0.006285f
C566 B.n521 VSUBS 0.006285f
C567 B.n522 VSUBS 0.006285f
C568 B.n523 VSUBS 0.006285f
C569 B.n524 VSUBS 0.006285f
C570 B.n525 VSUBS 0.006285f
C571 B.n526 VSUBS 0.01568f
C572 B.n527 VSUBS 0.015192f
C573 B.n528 VSUBS 0.015882f
C574 B.n529 VSUBS 0.006285f
C575 B.n530 VSUBS 0.006285f
C576 B.n531 VSUBS 0.006285f
C577 B.n532 VSUBS 0.006285f
C578 B.n533 VSUBS 0.006285f
C579 B.n534 VSUBS 0.006285f
C580 B.n535 VSUBS 0.006285f
C581 B.n536 VSUBS 0.006285f
C582 B.n537 VSUBS 0.006285f
C583 B.n538 VSUBS 0.006285f
C584 B.n539 VSUBS 0.006285f
C585 B.n540 VSUBS 0.006285f
C586 B.n541 VSUBS 0.006285f
C587 B.n542 VSUBS 0.006285f
C588 B.n543 VSUBS 0.006285f
C589 B.n544 VSUBS 0.006285f
C590 B.n545 VSUBS 0.006285f
C591 B.n546 VSUBS 0.006285f
C592 B.n547 VSUBS 0.006285f
C593 B.n548 VSUBS 0.006285f
C594 B.n549 VSUBS 0.006285f
C595 B.n550 VSUBS 0.006285f
C596 B.n551 VSUBS 0.006285f
C597 B.n552 VSUBS 0.006285f
C598 B.n553 VSUBS 0.006285f
C599 B.n554 VSUBS 0.006285f
C600 B.n555 VSUBS 0.006285f
C601 B.n556 VSUBS 0.006285f
C602 B.n557 VSUBS 0.006285f
C603 B.n558 VSUBS 0.006285f
C604 B.n559 VSUBS 0.006285f
C605 B.n560 VSUBS 0.006285f
C606 B.n561 VSUBS 0.006285f
C607 B.n562 VSUBS 0.006285f
C608 B.n563 VSUBS 0.006285f
C609 B.n564 VSUBS 0.006285f
C610 B.n565 VSUBS 0.006285f
C611 B.n566 VSUBS 0.006285f
C612 B.n567 VSUBS 0.006285f
C613 B.n568 VSUBS 0.006285f
C614 B.n569 VSUBS 0.006285f
C615 B.n570 VSUBS 0.006285f
C616 B.n571 VSUBS 0.006285f
C617 B.n572 VSUBS 0.006285f
C618 B.n573 VSUBS 0.006285f
C619 B.n574 VSUBS 0.006285f
C620 B.n575 VSUBS 0.006285f
C621 B.n576 VSUBS 0.006285f
C622 B.n577 VSUBS 0.006285f
C623 B.n578 VSUBS 0.006285f
C624 B.n579 VSUBS 0.006285f
C625 B.n580 VSUBS 0.006285f
C626 B.n581 VSUBS 0.006285f
C627 B.n582 VSUBS 0.006285f
C628 B.n583 VSUBS 0.006285f
C629 B.n584 VSUBS 0.006285f
C630 B.n585 VSUBS 0.006285f
C631 B.n586 VSUBS 0.006285f
C632 B.n587 VSUBS 0.006285f
C633 B.n588 VSUBS 0.006285f
C634 B.n589 VSUBS 0.006285f
C635 B.n590 VSUBS 0.006285f
C636 B.n591 VSUBS 0.006285f
C637 B.n592 VSUBS 0.006285f
C638 B.n593 VSUBS 0.006285f
C639 B.n594 VSUBS 0.006285f
C640 B.n595 VSUBS 0.006285f
C641 B.n596 VSUBS 0.006285f
C642 B.n597 VSUBS 0.006285f
C643 B.n598 VSUBS 0.006285f
C644 B.n599 VSUBS 0.006285f
C645 B.n600 VSUBS 0.006285f
C646 B.n601 VSUBS 0.006285f
C647 B.n602 VSUBS 0.006285f
C648 B.n603 VSUBS 0.006285f
C649 B.n604 VSUBS 0.006285f
C650 B.n605 VSUBS 0.006285f
C651 B.n606 VSUBS 0.006285f
C652 B.n607 VSUBS 0.006285f
C653 B.n608 VSUBS 0.006285f
C654 B.n609 VSUBS 0.005916f
C655 B.n610 VSUBS 0.014562f
C656 B.n611 VSUBS 0.003512f
C657 B.n612 VSUBS 0.006285f
C658 B.n613 VSUBS 0.006285f
C659 B.n614 VSUBS 0.006285f
C660 B.n615 VSUBS 0.006285f
C661 B.n616 VSUBS 0.006285f
C662 B.n617 VSUBS 0.006285f
C663 B.n618 VSUBS 0.006285f
C664 B.n619 VSUBS 0.006285f
C665 B.n620 VSUBS 0.006285f
C666 B.n621 VSUBS 0.006285f
C667 B.n622 VSUBS 0.006285f
C668 B.n623 VSUBS 0.006285f
C669 B.n624 VSUBS 0.003512f
C670 B.n625 VSUBS 0.006285f
C671 B.n626 VSUBS 0.006285f
C672 B.n627 VSUBS 0.005916f
C673 B.n628 VSUBS 0.006285f
C674 B.n629 VSUBS 0.006285f
C675 B.n630 VSUBS 0.006285f
C676 B.n631 VSUBS 0.006285f
C677 B.n632 VSUBS 0.006285f
C678 B.n633 VSUBS 0.006285f
C679 B.n634 VSUBS 0.006285f
C680 B.n635 VSUBS 0.006285f
C681 B.n636 VSUBS 0.006285f
C682 B.n637 VSUBS 0.006285f
C683 B.n638 VSUBS 0.006285f
C684 B.n639 VSUBS 0.006285f
C685 B.n640 VSUBS 0.006285f
C686 B.n641 VSUBS 0.006285f
C687 B.n642 VSUBS 0.006285f
C688 B.n643 VSUBS 0.006285f
C689 B.n644 VSUBS 0.006285f
C690 B.n645 VSUBS 0.006285f
C691 B.n646 VSUBS 0.006285f
C692 B.n647 VSUBS 0.006285f
C693 B.n648 VSUBS 0.006285f
C694 B.n649 VSUBS 0.006285f
C695 B.n650 VSUBS 0.006285f
C696 B.n651 VSUBS 0.006285f
C697 B.n652 VSUBS 0.006285f
C698 B.n653 VSUBS 0.006285f
C699 B.n654 VSUBS 0.006285f
C700 B.n655 VSUBS 0.006285f
C701 B.n656 VSUBS 0.006285f
C702 B.n657 VSUBS 0.006285f
C703 B.n658 VSUBS 0.006285f
C704 B.n659 VSUBS 0.006285f
C705 B.n660 VSUBS 0.006285f
C706 B.n661 VSUBS 0.006285f
C707 B.n662 VSUBS 0.006285f
C708 B.n663 VSUBS 0.006285f
C709 B.n664 VSUBS 0.006285f
C710 B.n665 VSUBS 0.006285f
C711 B.n666 VSUBS 0.006285f
C712 B.n667 VSUBS 0.006285f
C713 B.n668 VSUBS 0.006285f
C714 B.n669 VSUBS 0.006285f
C715 B.n670 VSUBS 0.006285f
C716 B.n671 VSUBS 0.006285f
C717 B.n672 VSUBS 0.006285f
C718 B.n673 VSUBS 0.006285f
C719 B.n674 VSUBS 0.006285f
C720 B.n675 VSUBS 0.006285f
C721 B.n676 VSUBS 0.006285f
C722 B.n677 VSUBS 0.006285f
C723 B.n678 VSUBS 0.006285f
C724 B.n679 VSUBS 0.006285f
C725 B.n680 VSUBS 0.006285f
C726 B.n681 VSUBS 0.006285f
C727 B.n682 VSUBS 0.006285f
C728 B.n683 VSUBS 0.006285f
C729 B.n684 VSUBS 0.006285f
C730 B.n685 VSUBS 0.006285f
C731 B.n686 VSUBS 0.006285f
C732 B.n687 VSUBS 0.006285f
C733 B.n688 VSUBS 0.006285f
C734 B.n689 VSUBS 0.006285f
C735 B.n690 VSUBS 0.006285f
C736 B.n691 VSUBS 0.006285f
C737 B.n692 VSUBS 0.006285f
C738 B.n693 VSUBS 0.006285f
C739 B.n694 VSUBS 0.006285f
C740 B.n695 VSUBS 0.006285f
C741 B.n696 VSUBS 0.006285f
C742 B.n697 VSUBS 0.006285f
C743 B.n698 VSUBS 0.006285f
C744 B.n699 VSUBS 0.006285f
C745 B.n700 VSUBS 0.006285f
C746 B.n701 VSUBS 0.006285f
C747 B.n702 VSUBS 0.006285f
C748 B.n703 VSUBS 0.006285f
C749 B.n704 VSUBS 0.006285f
C750 B.n705 VSUBS 0.006285f
C751 B.n706 VSUBS 0.006285f
C752 B.n707 VSUBS 0.015882f
C753 B.n708 VSUBS 0.015882f
C754 B.n709 VSUBS 0.01499f
C755 B.n710 VSUBS 0.006285f
C756 B.n711 VSUBS 0.006285f
C757 B.n712 VSUBS 0.006285f
C758 B.n713 VSUBS 0.006285f
C759 B.n714 VSUBS 0.006285f
C760 B.n715 VSUBS 0.006285f
C761 B.n716 VSUBS 0.006285f
C762 B.n717 VSUBS 0.006285f
C763 B.n718 VSUBS 0.006285f
C764 B.n719 VSUBS 0.006285f
C765 B.n720 VSUBS 0.006285f
C766 B.n721 VSUBS 0.006285f
C767 B.n722 VSUBS 0.006285f
C768 B.n723 VSUBS 0.006285f
C769 B.n724 VSUBS 0.006285f
C770 B.n725 VSUBS 0.006285f
C771 B.n726 VSUBS 0.006285f
C772 B.n727 VSUBS 0.006285f
C773 B.n728 VSUBS 0.006285f
C774 B.n729 VSUBS 0.006285f
C775 B.n730 VSUBS 0.006285f
C776 B.n731 VSUBS 0.006285f
C777 B.n732 VSUBS 0.006285f
C778 B.n733 VSUBS 0.006285f
C779 B.n734 VSUBS 0.006285f
C780 B.n735 VSUBS 0.006285f
C781 B.n736 VSUBS 0.006285f
C782 B.n737 VSUBS 0.006285f
C783 B.n738 VSUBS 0.006285f
C784 B.n739 VSUBS 0.006285f
C785 B.n740 VSUBS 0.006285f
C786 B.n741 VSUBS 0.006285f
C787 B.n742 VSUBS 0.006285f
C788 B.n743 VSUBS 0.006285f
C789 B.n744 VSUBS 0.006285f
C790 B.n745 VSUBS 0.006285f
C791 B.n746 VSUBS 0.006285f
C792 B.n747 VSUBS 0.006285f
C793 B.n748 VSUBS 0.006285f
C794 B.n749 VSUBS 0.006285f
C795 B.n750 VSUBS 0.006285f
C796 B.n751 VSUBS 0.006285f
C797 B.n752 VSUBS 0.006285f
C798 B.n753 VSUBS 0.006285f
C799 B.n754 VSUBS 0.006285f
C800 B.n755 VSUBS 0.006285f
C801 B.n756 VSUBS 0.006285f
C802 B.n757 VSUBS 0.006285f
C803 B.n758 VSUBS 0.006285f
C804 B.n759 VSUBS 0.014232f
C805 VDD2.t1 VSUBS 5.19819f
C806 VDD2.t0 VSUBS 4.10973f
C807 VDD2.n0 VSUBS 5.62671f
C808 VTAIL.t0 VSUBS 3.9145f
C809 VTAIL.n0 VSUBS 3.35205f
C810 VTAIL.t3 VSUBS 3.91451f
C811 VTAIL.n1 VSUBS 3.43271f
C812 VTAIL.t1 VSUBS 3.9145f
C813 VTAIL.n2 VSUBS 3.08828f
C814 VTAIL.t2 VSUBS 3.9145f
C815 VTAIL.n3 VSUBS 2.95277f
C816 VN.t0 VSUBS 5.69724f
C817 VN.t1 VSUBS 6.62805f
.ends

