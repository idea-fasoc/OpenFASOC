* NGSPICE file created from diff_pair_sample_0059.ext - technology: sky130A

.subckt diff_pair_sample_0059 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t1 VP.t0 VTAIL.t3 w_n2106_n1520# sky130_fd_pr__pfet_01v8 ad=1.0764 pd=6.3 as=1.0764 ps=6.3 w=2.76 l=2.51
X1 B.t11 B.t9 B.t10 w_n2106_n1520# sky130_fd_pr__pfet_01v8 ad=1.0764 pd=6.3 as=0 ps=0 w=2.76 l=2.51
X2 VDD1.t0 VP.t1 VTAIL.t2 w_n2106_n1520# sky130_fd_pr__pfet_01v8 ad=1.0764 pd=6.3 as=1.0764 ps=6.3 w=2.76 l=2.51
X3 VDD2.t1 VN.t0 VTAIL.t1 w_n2106_n1520# sky130_fd_pr__pfet_01v8 ad=1.0764 pd=6.3 as=1.0764 ps=6.3 w=2.76 l=2.51
X4 B.t8 B.t6 B.t7 w_n2106_n1520# sky130_fd_pr__pfet_01v8 ad=1.0764 pd=6.3 as=0 ps=0 w=2.76 l=2.51
X5 B.t5 B.t3 B.t4 w_n2106_n1520# sky130_fd_pr__pfet_01v8 ad=1.0764 pd=6.3 as=0 ps=0 w=2.76 l=2.51
X6 VDD2.t0 VN.t1 VTAIL.t0 w_n2106_n1520# sky130_fd_pr__pfet_01v8 ad=1.0764 pd=6.3 as=1.0764 ps=6.3 w=2.76 l=2.51
X7 B.t2 B.t0 B.t1 w_n2106_n1520# sky130_fd_pr__pfet_01v8 ad=1.0764 pd=6.3 as=0 ps=0 w=2.76 l=2.51
R0 VP.n0 VP.t0 113.133
R1 VP.n0 VP.t1 75.7159
R2 VP VP.n0 0.336784
R3 VTAIL.n1 VTAIL.t1 133.168
R4 VTAIL.n3 VTAIL.t0 133.168
R5 VTAIL.n0 VTAIL.t2 133.168
R6 VTAIL.n2 VTAIL.t3 133.168
R7 VTAIL.n1 VTAIL.n0 19.6427
R8 VTAIL.n3 VTAIL.n2 17.1945
R9 VTAIL.n2 VTAIL.n1 1.69447
R10 VTAIL VTAIL.n0 1.14059
R11 VTAIL VTAIL.n3 0.554379
R12 VDD1 VDD1.t0 181.919
R13 VDD1 VDD1.t1 150.518
R14 B.n271 B.n38 585
R15 B.n273 B.n272 585
R16 B.n274 B.n37 585
R17 B.n276 B.n275 585
R18 B.n277 B.n36 585
R19 B.n279 B.n278 585
R20 B.n280 B.n35 585
R21 B.n282 B.n281 585
R22 B.n283 B.n34 585
R23 B.n285 B.n284 585
R24 B.n286 B.n33 585
R25 B.n288 B.n287 585
R26 B.n289 B.n29 585
R27 B.n291 B.n290 585
R28 B.n292 B.n28 585
R29 B.n294 B.n293 585
R30 B.n295 B.n27 585
R31 B.n297 B.n296 585
R32 B.n298 B.n26 585
R33 B.n300 B.n299 585
R34 B.n301 B.n25 585
R35 B.n303 B.n302 585
R36 B.n304 B.n24 585
R37 B.n306 B.n305 585
R38 B.n308 B.n21 585
R39 B.n310 B.n309 585
R40 B.n311 B.n20 585
R41 B.n313 B.n312 585
R42 B.n314 B.n19 585
R43 B.n316 B.n315 585
R44 B.n317 B.n18 585
R45 B.n319 B.n318 585
R46 B.n320 B.n17 585
R47 B.n322 B.n321 585
R48 B.n323 B.n16 585
R49 B.n325 B.n324 585
R50 B.n326 B.n15 585
R51 B.n328 B.n327 585
R52 B.n270 B.n269 585
R53 B.n268 B.n39 585
R54 B.n267 B.n266 585
R55 B.n265 B.n40 585
R56 B.n264 B.n263 585
R57 B.n262 B.n41 585
R58 B.n261 B.n260 585
R59 B.n259 B.n42 585
R60 B.n258 B.n257 585
R61 B.n256 B.n43 585
R62 B.n255 B.n254 585
R63 B.n253 B.n44 585
R64 B.n252 B.n251 585
R65 B.n250 B.n45 585
R66 B.n249 B.n248 585
R67 B.n247 B.n46 585
R68 B.n246 B.n245 585
R69 B.n244 B.n47 585
R70 B.n243 B.n242 585
R71 B.n241 B.n48 585
R72 B.n240 B.n239 585
R73 B.n238 B.n49 585
R74 B.n237 B.n236 585
R75 B.n235 B.n50 585
R76 B.n234 B.n233 585
R77 B.n232 B.n51 585
R78 B.n231 B.n230 585
R79 B.n229 B.n52 585
R80 B.n228 B.n227 585
R81 B.n226 B.n53 585
R82 B.n225 B.n224 585
R83 B.n223 B.n54 585
R84 B.n222 B.n221 585
R85 B.n220 B.n55 585
R86 B.n219 B.n218 585
R87 B.n217 B.n56 585
R88 B.n216 B.n215 585
R89 B.n214 B.n57 585
R90 B.n213 B.n212 585
R91 B.n211 B.n58 585
R92 B.n210 B.n209 585
R93 B.n208 B.n59 585
R94 B.n207 B.n206 585
R95 B.n205 B.n60 585
R96 B.n204 B.n203 585
R97 B.n202 B.n61 585
R98 B.n201 B.n200 585
R99 B.n199 B.n62 585
R100 B.n198 B.n197 585
R101 B.n196 B.n63 585
R102 B.n195 B.n194 585
R103 B.n136 B.n87 585
R104 B.n138 B.n137 585
R105 B.n139 B.n86 585
R106 B.n141 B.n140 585
R107 B.n142 B.n85 585
R108 B.n144 B.n143 585
R109 B.n145 B.n84 585
R110 B.n147 B.n146 585
R111 B.n148 B.n83 585
R112 B.n150 B.n149 585
R113 B.n151 B.n82 585
R114 B.n153 B.n152 585
R115 B.n154 B.n81 585
R116 B.n156 B.n155 585
R117 B.n158 B.n78 585
R118 B.n160 B.n159 585
R119 B.n161 B.n77 585
R120 B.n163 B.n162 585
R121 B.n164 B.n76 585
R122 B.n166 B.n165 585
R123 B.n167 B.n75 585
R124 B.n169 B.n168 585
R125 B.n170 B.n74 585
R126 B.n172 B.n171 585
R127 B.n174 B.n173 585
R128 B.n175 B.n70 585
R129 B.n177 B.n176 585
R130 B.n178 B.n69 585
R131 B.n180 B.n179 585
R132 B.n181 B.n68 585
R133 B.n183 B.n182 585
R134 B.n184 B.n67 585
R135 B.n186 B.n185 585
R136 B.n187 B.n66 585
R137 B.n189 B.n188 585
R138 B.n190 B.n65 585
R139 B.n192 B.n191 585
R140 B.n193 B.n64 585
R141 B.n135 B.n134 585
R142 B.n133 B.n88 585
R143 B.n132 B.n131 585
R144 B.n130 B.n89 585
R145 B.n129 B.n128 585
R146 B.n127 B.n90 585
R147 B.n126 B.n125 585
R148 B.n124 B.n91 585
R149 B.n123 B.n122 585
R150 B.n121 B.n92 585
R151 B.n120 B.n119 585
R152 B.n118 B.n93 585
R153 B.n117 B.n116 585
R154 B.n115 B.n94 585
R155 B.n114 B.n113 585
R156 B.n112 B.n95 585
R157 B.n111 B.n110 585
R158 B.n109 B.n96 585
R159 B.n108 B.n107 585
R160 B.n106 B.n97 585
R161 B.n105 B.n104 585
R162 B.n103 B.n98 585
R163 B.n102 B.n101 585
R164 B.n100 B.n99 585
R165 B.n2 B.n0 585
R166 B.n365 B.n1 585
R167 B.n364 B.n363 585
R168 B.n362 B.n3 585
R169 B.n361 B.n360 585
R170 B.n359 B.n4 585
R171 B.n358 B.n357 585
R172 B.n356 B.n5 585
R173 B.n355 B.n354 585
R174 B.n353 B.n6 585
R175 B.n352 B.n351 585
R176 B.n350 B.n7 585
R177 B.n349 B.n348 585
R178 B.n347 B.n8 585
R179 B.n346 B.n345 585
R180 B.n344 B.n9 585
R181 B.n343 B.n342 585
R182 B.n341 B.n10 585
R183 B.n340 B.n339 585
R184 B.n338 B.n11 585
R185 B.n337 B.n336 585
R186 B.n335 B.n12 585
R187 B.n334 B.n333 585
R188 B.n332 B.n13 585
R189 B.n331 B.n330 585
R190 B.n329 B.n14 585
R191 B.n367 B.n366 585
R192 B.n136 B.n135 506.916
R193 B.n329 B.n328 506.916
R194 B.n195 B.n64 506.916
R195 B.n269 B.n38 506.916
R196 B.n71 B.t6 234.407
R197 B.n79 B.t3 234.407
R198 B.n22 B.t9 234.407
R199 B.n30 B.t0 234.407
R200 B.n71 B.t8 196.589
R201 B.n30 B.t1 196.589
R202 B.n79 B.t5 196.588
R203 B.n22 B.t10 196.588
R204 B.n135 B.n88 163.367
R205 B.n131 B.n88 163.367
R206 B.n131 B.n130 163.367
R207 B.n130 B.n129 163.367
R208 B.n129 B.n90 163.367
R209 B.n125 B.n90 163.367
R210 B.n125 B.n124 163.367
R211 B.n124 B.n123 163.367
R212 B.n123 B.n92 163.367
R213 B.n119 B.n92 163.367
R214 B.n119 B.n118 163.367
R215 B.n118 B.n117 163.367
R216 B.n117 B.n94 163.367
R217 B.n113 B.n94 163.367
R218 B.n113 B.n112 163.367
R219 B.n112 B.n111 163.367
R220 B.n111 B.n96 163.367
R221 B.n107 B.n96 163.367
R222 B.n107 B.n106 163.367
R223 B.n106 B.n105 163.367
R224 B.n105 B.n98 163.367
R225 B.n101 B.n98 163.367
R226 B.n101 B.n100 163.367
R227 B.n100 B.n2 163.367
R228 B.n366 B.n2 163.367
R229 B.n366 B.n365 163.367
R230 B.n365 B.n364 163.367
R231 B.n364 B.n3 163.367
R232 B.n360 B.n3 163.367
R233 B.n360 B.n359 163.367
R234 B.n359 B.n358 163.367
R235 B.n358 B.n5 163.367
R236 B.n354 B.n5 163.367
R237 B.n354 B.n353 163.367
R238 B.n353 B.n352 163.367
R239 B.n352 B.n7 163.367
R240 B.n348 B.n7 163.367
R241 B.n348 B.n347 163.367
R242 B.n347 B.n346 163.367
R243 B.n346 B.n9 163.367
R244 B.n342 B.n9 163.367
R245 B.n342 B.n341 163.367
R246 B.n341 B.n340 163.367
R247 B.n340 B.n11 163.367
R248 B.n336 B.n11 163.367
R249 B.n336 B.n335 163.367
R250 B.n335 B.n334 163.367
R251 B.n334 B.n13 163.367
R252 B.n330 B.n13 163.367
R253 B.n330 B.n329 163.367
R254 B.n137 B.n136 163.367
R255 B.n137 B.n86 163.367
R256 B.n141 B.n86 163.367
R257 B.n142 B.n141 163.367
R258 B.n143 B.n142 163.367
R259 B.n143 B.n84 163.367
R260 B.n147 B.n84 163.367
R261 B.n148 B.n147 163.367
R262 B.n149 B.n148 163.367
R263 B.n149 B.n82 163.367
R264 B.n153 B.n82 163.367
R265 B.n154 B.n153 163.367
R266 B.n155 B.n154 163.367
R267 B.n155 B.n78 163.367
R268 B.n160 B.n78 163.367
R269 B.n161 B.n160 163.367
R270 B.n162 B.n161 163.367
R271 B.n162 B.n76 163.367
R272 B.n166 B.n76 163.367
R273 B.n167 B.n166 163.367
R274 B.n168 B.n167 163.367
R275 B.n168 B.n74 163.367
R276 B.n172 B.n74 163.367
R277 B.n173 B.n172 163.367
R278 B.n173 B.n70 163.367
R279 B.n177 B.n70 163.367
R280 B.n178 B.n177 163.367
R281 B.n179 B.n178 163.367
R282 B.n179 B.n68 163.367
R283 B.n183 B.n68 163.367
R284 B.n184 B.n183 163.367
R285 B.n185 B.n184 163.367
R286 B.n185 B.n66 163.367
R287 B.n189 B.n66 163.367
R288 B.n190 B.n189 163.367
R289 B.n191 B.n190 163.367
R290 B.n191 B.n64 163.367
R291 B.n196 B.n195 163.367
R292 B.n197 B.n196 163.367
R293 B.n197 B.n62 163.367
R294 B.n201 B.n62 163.367
R295 B.n202 B.n201 163.367
R296 B.n203 B.n202 163.367
R297 B.n203 B.n60 163.367
R298 B.n207 B.n60 163.367
R299 B.n208 B.n207 163.367
R300 B.n209 B.n208 163.367
R301 B.n209 B.n58 163.367
R302 B.n213 B.n58 163.367
R303 B.n214 B.n213 163.367
R304 B.n215 B.n214 163.367
R305 B.n215 B.n56 163.367
R306 B.n219 B.n56 163.367
R307 B.n220 B.n219 163.367
R308 B.n221 B.n220 163.367
R309 B.n221 B.n54 163.367
R310 B.n225 B.n54 163.367
R311 B.n226 B.n225 163.367
R312 B.n227 B.n226 163.367
R313 B.n227 B.n52 163.367
R314 B.n231 B.n52 163.367
R315 B.n232 B.n231 163.367
R316 B.n233 B.n232 163.367
R317 B.n233 B.n50 163.367
R318 B.n237 B.n50 163.367
R319 B.n238 B.n237 163.367
R320 B.n239 B.n238 163.367
R321 B.n239 B.n48 163.367
R322 B.n243 B.n48 163.367
R323 B.n244 B.n243 163.367
R324 B.n245 B.n244 163.367
R325 B.n245 B.n46 163.367
R326 B.n249 B.n46 163.367
R327 B.n250 B.n249 163.367
R328 B.n251 B.n250 163.367
R329 B.n251 B.n44 163.367
R330 B.n255 B.n44 163.367
R331 B.n256 B.n255 163.367
R332 B.n257 B.n256 163.367
R333 B.n257 B.n42 163.367
R334 B.n261 B.n42 163.367
R335 B.n262 B.n261 163.367
R336 B.n263 B.n262 163.367
R337 B.n263 B.n40 163.367
R338 B.n267 B.n40 163.367
R339 B.n268 B.n267 163.367
R340 B.n269 B.n268 163.367
R341 B.n328 B.n15 163.367
R342 B.n324 B.n15 163.367
R343 B.n324 B.n323 163.367
R344 B.n323 B.n322 163.367
R345 B.n322 B.n17 163.367
R346 B.n318 B.n17 163.367
R347 B.n318 B.n317 163.367
R348 B.n317 B.n316 163.367
R349 B.n316 B.n19 163.367
R350 B.n312 B.n19 163.367
R351 B.n312 B.n311 163.367
R352 B.n311 B.n310 163.367
R353 B.n310 B.n21 163.367
R354 B.n305 B.n21 163.367
R355 B.n305 B.n304 163.367
R356 B.n304 B.n303 163.367
R357 B.n303 B.n25 163.367
R358 B.n299 B.n25 163.367
R359 B.n299 B.n298 163.367
R360 B.n298 B.n297 163.367
R361 B.n297 B.n27 163.367
R362 B.n293 B.n27 163.367
R363 B.n293 B.n292 163.367
R364 B.n292 B.n291 163.367
R365 B.n291 B.n29 163.367
R366 B.n287 B.n29 163.367
R367 B.n287 B.n286 163.367
R368 B.n286 B.n285 163.367
R369 B.n285 B.n34 163.367
R370 B.n281 B.n34 163.367
R371 B.n281 B.n280 163.367
R372 B.n280 B.n279 163.367
R373 B.n279 B.n36 163.367
R374 B.n275 B.n36 163.367
R375 B.n275 B.n274 163.367
R376 B.n274 B.n273 163.367
R377 B.n273 B.n38 163.367
R378 B.n72 B.t7 141.511
R379 B.n31 B.t2 141.511
R380 B.n80 B.t4 141.508
R381 B.n23 B.t11 141.508
R382 B.n73 B.n72 59.5399
R383 B.n157 B.n80 59.5399
R384 B.n307 B.n23 59.5399
R385 B.n32 B.n31 59.5399
R386 B.n72 B.n71 55.0793
R387 B.n80 B.n79 55.0793
R388 B.n23 B.n22 55.0793
R389 B.n31 B.n30 55.0793
R390 B.n327 B.n14 32.9371
R391 B.n271 B.n270 32.9371
R392 B.n194 B.n193 32.9371
R393 B.n134 B.n87 32.9371
R394 B B.n367 18.0485
R395 B.n327 B.n326 10.6151
R396 B.n326 B.n325 10.6151
R397 B.n325 B.n16 10.6151
R398 B.n321 B.n16 10.6151
R399 B.n321 B.n320 10.6151
R400 B.n320 B.n319 10.6151
R401 B.n319 B.n18 10.6151
R402 B.n315 B.n18 10.6151
R403 B.n315 B.n314 10.6151
R404 B.n314 B.n313 10.6151
R405 B.n313 B.n20 10.6151
R406 B.n309 B.n20 10.6151
R407 B.n309 B.n308 10.6151
R408 B.n306 B.n24 10.6151
R409 B.n302 B.n24 10.6151
R410 B.n302 B.n301 10.6151
R411 B.n301 B.n300 10.6151
R412 B.n300 B.n26 10.6151
R413 B.n296 B.n26 10.6151
R414 B.n296 B.n295 10.6151
R415 B.n295 B.n294 10.6151
R416 B.n294 B.n28 10.6151
R417 B.n290 B.n289 10.6151
R418 B.n289 B.n288 10.6151
R419 B.n288 B.n33 10.6151
R420 B.n284 B.n33 10.6151
R421 B.n284 B.n283 10.6151
R422 B.n283 B.n282 10.6151
R423 B.n282 B.n35 10.6151
R424 B.n278 B.n35 10.6151
R425 B.n278 B.n277 10.6151
R426 B.n277 B.n276 10.6151
R427 B.n276 B.n37 10.6151
R428 B.n272 B.n37 10.6151
R429 B.n272 B.n271 10.6151
R430 B.n194 B.n63 10.6151
R431 B.n198 B.n63 10.6151
R432 B.n199 B.n198 10.6151
R433 B.n200 B.n199 10.6151
R434 B.n200 B.n61 10.6151
R435 B.n204 B.n61 10.6151
R436 B.n205 B.n204 10.6151
R437 B.n206 B.n205 10.6151
R438 B.n206 B.n59 10.6151
R439 B.n210 B.n59 10.6151
R440 B.n211 B.n210 10.6151
R441 B.n212 B.n211 10.6151
R442 B.n212 B.n57 10.6151
R443 B.n216 B.n57 10.6151
R444 B.n217 B.n216 10.6151
R445 B.n218 B.n217 10.6151
R446 B.n218 B.n55 10.6151
R447 B.n222 B.n55 10.6151
R448 B.n223 B.n222 10.6151
R449 B.n224 B.n223 10.6151
R450 B.n224 B.n53 10.6151
R451 B.n228 B.n53 10.6151
R452 B.n229 B.n228 10.6151
R453 B.n230 B.n229 10.6151
R454 B.n230 B.n51 10.6151
R455 B.n234 B.n51 10.6151
R456 B.n235 B.n234 10.6151
R457 B.n236 B.n235 10.6151
R458 B.n236 B.n49 10.6151
R459 B.n240 B.n49 10.6151
R460 B.n241 B.n240 10.6151
R461 B.n242 B.n241 10.6151
R462 B.n242 B.n47 10.6151
R463 B.n246 B.n47 10.6151
R464 B.n247 B.n246 10.6151
R465 B.n248 B.n247 10.6151
R466 B.n248 B.n45 10.6151
R467 B.n252 B.n45 10.6151
R468 B.n253 B.n252 10.6151
R469 B.n254 B.n253 10.6151
R470 B.n254 B.n43 10.6151
R471 B.n258 B.n43 10.6151
R472 B.n259 B.n258 10.6151
R473 B.n260 B.n259 10.6151
R474 B.n260 B.n41 10.6151
R475 B.n264 B.n41 10.6151
R476 B.n265 B.n264 10.6151
R477 B.n266 B.n265 10.6151
R478 B.n266 B.n39 10.6151
R479 B.n270 B.n39 10.6151
R480 B.n138 B.n87 10.6151
R481 B.n139 B.n138 10.6151
R482 B.n140 B.n139 10.6151
R483 B.n140 B.n85 10.6151
R484 B.n144 B.n85 10.6151
R485 B.n145 B.n144 10.6151
R486 B.n146 B.n145 10.6151
R487 B.n146 B.n83 10.6151
R488 B.n150 B.n83 10.6151
R489 B.n151 B.n150 10.6151
R490 B.n152 B.n151 10.6151
R491 B.n152 B.n81 10.6151
R492 B.n156 B.n81 10.6151
R493 B.n159 B.n158 10.6151
R494 B.n159 B.n77 10.6151
R495 B.n163 B.n77 10.6151
R496 B.n164 B.n163 10.6151
R497 B.n165 B.n164 10.6151
R498 B.n165 B.n75 10.6151
R499 B.n169 B.n75 10.6151
R500 B.n170 B.n169 10.6151
R501 B.n171 B.n170 10.6151
R502 B.n175 B.n174 10.6151
R503 B.n176 B.n175 10.6151
R504 B.n176 B.n69 10.6151
R505 B.n180 B.n69 10.6151
R506 B.n181 B.n180 10.6151
R507 B.n182 B.n181 10.6151
R508 B.n182 B.n67 10.6151
R509 B.n186 B.n67 10.6151
R510 B.n187 B.n186 10.6151
R511 B.n188 B.n187 10.6151
R512 B.n188 B.n65 10.6151
R513 B.n192 B.n65 10.6151
R514 B.n193 B.n192 10.6151
R515 B.n134 B.n133 10.6151
R516 B.n133 B.n132 10.6151
R517 B.n132 B.n89 10.6151
R518 B.n128 B.n89 10.6151
R519 B.n128 B.n127 10.6151
R520 B.n127 B.n126 10.6151
R521 B.n126 B.n91 10.6151
R522 B.n122 B.n91 10.6151
R523 B.n122 B.n121 10.6151
R524 B.n121 B.n120 10.6151
R525 B.n120 B.n93 10.6151
R526 B.n116 B.n93 10.6151
R527 B.n116 B.n115 10.6151
R528 B.n115 B.n114 10.6151
R529 B.n114 B.n95 10.6151
R530 B.n110 B.n95 10.6151
R531 B.n110 B.n109 10.6151
R532 B.n109 B.n108 10.6151
R533 B.n108 B.n97 10.6151
R534 B.n104 B.n97 10.6151
R535 B.n104 B.n103 10.6151
R536 B.n103 B.n102 10.6151
R537 B.n102 B.n99 10.6151
R538 B.n99 B.n0 10.6151
R539 B.n363 B.n1 10.6151
R540 B.n363 B.n362 10.6151
R541 B.n362 B.n361 10.6151
R542 B.n361 B.n4 10.6151
R543 B.n357 B.n4 10.6151
R544 B.n357 B.n356 10.6151
R545 B.n356 B.n355 10.6151
R546 B.n355 B.n6 10.6151
R547 B.n351 B.n6 10.6151
R548 B.n351 B.n350 10.6151
R549 B.n350 B.n349 10.6151
R550 B.n349 B.n8 10.6151
R551 B.n345 B.n8 10.6151
R552 B.n345 B.n344 10.6151
R553 B.n344 B.n343 10.6151
R554 B.n343 B.n10 10.6151
R555 B.n339 B.n10 10.6151
R556 B.n339 B.n338 10.6151
R557 B.n338 B.n337 10.6151
R558 B.n337 B.n12 10.6151
R559 B.n333 B.n12 10.6151
R560 B.n333 B.n332 10.6151
R561 B.n332 B.n331 10.6151
R562 B.n331 B.n14 10.6151
R563 B.n308 B.n307 9.36635
R564 B.n290 B.n32 9.36635
R565 B.n157 B.n156 9.36635
R566 B.n174 B.n73 9.36635
R567 B.n367 B.n0 2.81026
R568 B.n367 B.n1 2.81026
R569 B.n307 B.n306 1.24928
R570 B.n32 B.n28 1.24928
R571 B.n158 B.n157 1.24928
R572 B.n171 B.n73 1.24928
R573 VN VN.t0 113.231
R574 VN VN.t1 76.0522
R575 VDD2.n0 VDD2.t0 180.782
R576 VDD2.n0 VDD2.t1 149.847
R577 VDD2 VDD2.n0 0.670759
C0 VDD1 VP 1.01126f
C1 VDD2 B 0.99319f
C2 VTAIL VN 1.04377f
C3 VP w_n2106_n1520# 2.96981f
C4 VDD2 VP 0.334774f
C5 VDD1 VN 0.153765f
C6 VP B 1.34725f
C7 VN w_n2106_n1520# 2.70449f
C8 VDD2 VN 0.831784f
C9 VDD1 VTAIL 2.59713f
C10 VTAIL w_n2106_n1520# 1.41625f
C11 VN B 0.907386f
C12 VDD2 VTAIL 2.64926f
C13 VDD1 w_n2106_n1520# 1.12394f
C14 VTAIL B 1.49798f
C15 VN VP 3.70385f
C16 VDD2 VDD1 0.662695f
C17 VTAIL VP 1.05792f
C18 VDD1 B 0.96368f
C19 VDD2 w_n2106_n1520# 1.14817f
C20 B w_n2106_n1520# 6.14045f
C21 VDD2 VSUBS 0.559242f
C22 VDD1 VSUBS 2.649555f
C23 VTAIL VSUBS 0.389329f
C24 VN VSUBS 5.2878f
C25 VP VSUBS 1.2044f
C26 B VSUBS 2.905889f
C27 w_n2106_n1520# VSUBS 40.612103f
C28 VDD2.t0 VSUBS 0.403652f
C29 VDD2.t1 VSUBS 0.261099f
C30 VDD2.n0 VSUBS 1.83472f
C31 VN.t1 VSUBS 1.19732f
C32 VN.t0 VSUBS 1.84762f
C33 B.n0 VSUBS 0.005191f
C34 B.n1 VSUBS 0.005191f
C35 B.n2 VSUBS 0.008209f
C36 B.n3 VSUBS 0.008209f
C37 B.n4 VSUBS 0.008209f
C38 B.n5 VSUBS 0.008209f
C39 B.n6 VSUBS 0.008209f
C40 B.n7 VSUBS 0.008209f
C41 B.n8 VSUBS 0.008209f
C42 B.n9 VSUBS 0.008209f
C43 B.n10 VSUBS 0.008209f
C44 B.n11 VSUBS 0.008209f
C45 B.n12 VSUBS 0.008209f
C46 B.n13 VSUBS 0.008209f
C47 B.n14 VSUBS 0.019186f
C48 B.n15 VSUBS 0.008209f
C49 B.n16 VSUBS 0.008209f
C50 B.n17 VSUBS 0.008209f
C51 B.n18 VSUBS 0.008209f
C52 B.n19 VSUBS 0.008209f
C53 B.n20 VSUBS 0.008209f
C54 B.n21 VSUBS 0.008209f
C55 B.t11 VSUBS 0.076302f
C56 B.t10 VSUBS 0.093835f
C57 B.t9 VSUBS 0.395784f
C58 B.n22 VSUBS 0.091204f
C59 B.n23 VSUBS 0.074285f
C60 B.n24 VSUBS 0.008209f
C61 B.n25 VSUBS 0.008209f
C62 B.n26 VSUBS 0.008209f
C63 B.n27 VSUBS 0.008209f
C64 B.n28 VSUBS 0.004587f
C65 B.n29 VSUBS 0.008209f
C66 B.t2 VSUBS 0.076302f
C67 B.t1 VSUBS 0.093835f
C68 B.t0 VSUBS 0.395784f
C69 B.n30 VSUBS 0.091204f
C70 B.n31 VSUBS 0.074285f
C71 B.n32 VSUBS 0.019019f
C72 B.n33 VSUBS 0.008209f
C73 B.n34 VSUBS 0.008209f
C74 B.n35 VSUBS 0.008209f
C75 B.n36 VSUBS 0.008209f
C76 B.n37 VSUBS 0.008209f
C77 B.n38 VSUBS 0.019444f
C78 B.n39 VSUBS 0.008209f
C79 B.n40 VSUBS 0.008209f
C80 B.n41 VSUBS 0.008209f
C81 B.n42 VSUBS 0.008209f
C82 B.n43 VSUBS 0.008209f
C83 B.n44 VSUBS 0.008209f
C84 B.n45 VSUBS 0.008209f
C85 B.n46 VSUBS 0.008209f
C86 B.n47 VSUBS 0.008209f
C87 B.n48 VSUBS 0.008209f
C88 B.n49 VSUBS 0.008209f
C89 B.n50 VSUBS 0.008209f
C90 B.n51 VSUBS 0.008209f
C91 B.n52 VSUBS 0.008209f
C92 B.n53 VSUBS 0.008209f
C93 B.n54 VSUBS 0.008209f
C94 B.n55 VSUBS 0.008209f
C95 B.n56 VSUBS 0.008209f
C96 B.n57 VSUBS 0.008209f
C97 B.n58 VSUBS 0.008209f
C98 B.n59 VSUBS 0.008209f
C99 B.n60 VSUBS 0.008209f
C100 B.n61 VSUBS 0.008209f
C101 B.n62 VSUBS 0.008209f
C102 B.n63 VSUBS 0.008209f
C103 B.n64 VSUBS 0.019444f
C104 B.n65 VSUBS 0.008209f
C105 B.n66 VSUBS 0.008209f
C106 B.n67 VSUBS 0.008209f
C107 B.n68 VSUBS 0.008209f
C108 B.n69 VSUBS 0.008209f
C109 B.n70 VSUBS 0.008209f
C110 B.t7 VSUBS 0.076302f
C111 B.t8 VSUBS 0.093835f
C112 B.t6 VSUBS 0.395784f
C113 B.n71 VSUBS 0.091204f
C114 B.n72 VSUBS 0.074285f
C115 B.n73 VSUBS 0.019019f
C116 B.n74 VSUBS 0.008209f
C117 B.n75 VSUBS 0.008209f
C118 B.n76 VSUBS 0.008209f
C119 B.n77 VSUBS 0.008209f
C120 B.n78 VSUBS 0.008209f
C121 B.t4 VSUBS 0.076302f
C122 B.t5 VSUBS 0.093835f
C123 B.t3 VSUBS 0.395784f
C124 B.n79 VSUBS 0.091204f
C125 B.n80 VSUBS 0.074285f
C126 B.n81 VSUBS 0.008209f
C127 B.n82 VSUBS 0.008209f
C128 B.n83 VSUBS 0.008209f
C129 B.n84 VSUBS 0.008209f
C130 B.n85 VSUBS 0.008209f
C131 B.n86 VSUBS 0.008209f
C132 B.n87 VSUBS 0.019444f
C133 B.n88 VSUBS 0.008209f
C134 B.n89 VSUBS 0.008209f
C135 B.n90 VSUBS 0.008209f
C136 B.n91 VSUBS 0.008209f
C137 B.n92 VSUBS 0.008209f
C138 B.n93 VSUBS 0.008209f
C139 B.n94 VSUBS 0.008209f
C140 B.n95 VSUBS 0.008209f
C141 B.n96 VSUBS 0.008209f
C142 B.n97 VSUBS 0.008209f
C143 B.n98 VSUBS 0.008209f
C144 B.n99 VSUBS 0.008209f
C145 B.n100 VSUBS 0.008209f
C146 B.n101 VSUBS 0.008209f
C147 B.n102 VSUBS 0.008209f
C148 B.n103 VSUBS 0.008209f
C149 B.n104 VSUBS 0.008209f
C150 B.n105 VSUBS 0.008209f
C151 B.n106 VSUBS 0.008209f
C152 B.n107 VSUBS 0.008209f
C153 B.n108 VSUBS 0.008209f
C154 B.n109 VSUBS 0.008209f
C155 B.n110 VSUBS 0.008209f
C156 B.n111 VSUBS 0.008209f
C157 B.n112 VSUBS 0.008209f
C158 B.n113 VSUBS 0.008209f
C159 B.n114 VSUBS 0.008209f
C160 B.n115 VSUBS 0.008209f
C161 B.n116 VSUBS 0.008209f
C162 B.n117 VSUBS 0.008209f
C163 B.n118 VSUBS 0.008209f
C164 B.n119 VSUBS 0.008209f
C165 B.n120 VSUBS 0.008209f
C166 B.n121 VSUBS 0.008209f
C167 B.n122 VSUBS 0.008209f
C168 B.n123 VSUBS 0.008209f
C169 B.n124 VSUBS 0.008209f
C170 B.n125 VSUBS 0.008209f
C171 B.n126 VSUBS 0.008209f
C172 B.n127 VSUBS 0.008209f
C173 B.n128 VSUBS 0.008209f
C174 B.n129 VSUBS 0.008209f
C175 B.n130 VSUBS 0.008209f
C176 B.n131 VSUBS 0.008209f
C177 B.n132 VSUBS 0.008209f
C178 B.n133 VSUBS 0.008209f
C179 B.n134 VSUBS 0.019186f
C180 B.n135 VSUBS 0.019186f
C181 B.n136 VSUBS 0.019444f
C182 B.n137 VSUBS 0.008209f
C183 B.n138 VSUBS 0.008209f
C184 B.n139 VSUBS 0.008209f
C185 B.n140 VSUBS 0.008209f
C186 B.n141 VSUBS 0.008209f
C187 B.n142 VSUBS 0.008209f
C188 B.n143 VSUBS 0.008209f
C189 B.n144 VSUBS 0.008209f
C190 B.n145 VSUBS 0.008209f
C191 B.n146 VSUBS 0.008209f
C192 B.n147 VSUBS 0.008209f
C193 B.n148 VSUBS 0.008209f
C194 B.n149 VSUBS 0.008209f
C195 B.n150 VSUBS 0.008209f
C196 B.n151 VSUBS 0.008209f
C197 B.n152 VSUBS 0.008209f
C198 B.n153 VSUBS 0.008209f
C199 B.n154 VSUBS 0.008209f
C200 B.n155 VSUBS 0.008209f
C201 B.n156 VSUBS 0.007726f
C202 B.n157 VSUBS 0.019019f
C203 B.n158 VSUBS 0.004587f
C204 B.n159 VSUBS 0.008209f
C205 B.n160 VSUBS 0.008209f
C206 B.n161 VSUBS 0.008209f
C207 B.n162 VSUBS 0.008209f
C208 B.n163 VSUBS 0.008209f
C209 B.n164 VSUBS 0.008209f
C210 B.n165 VSUBS 0.008209f
C211 B.n166 VSUBS 0.008209f
C212 B.n167 VSUBS 0.008209f
C213 B.n168 VSUBS 0.008209f
C214 B.n169 VSUBS 0.008209f
C215 B.n170 VSUBS 0.008209f
C216 B.n171 VSUBS 0.004587f
C217 B.n172 VSUBS 0.008209f
C218 B.n173 VSUBS 0.008209f
C219 B.n174 VSUBS 0.007726f
C220 B.n175 VSUBS 0.008209f
C221 B.n176 VSUBS 0.008209f
C222 B.n177 VSUBS 0.008209f
C223 B.n178 VSUBS 0.008209f
C224 B.n179 VSUBS 0.008209f
C225 B.n180 VSUBS 0.008209f
C226 B.n181 VSUBS 0.008209f
C227 B.n182 VSUBS 0.008209f
C228 B.n183 VSUBS 0.008209f
C229 B.n184 VSUBS 0.008209f
C230 B.n185 VSUBS 0.008209f
C231 B.n186 VSUBS 0.008209f
C232 B.n187 VSUBS 0.008209f
C233 B.n188 VSUBS 0.008209f
C234 B.n189 VSUBS 0.008209f
C235 B.n190 VSUBS 0.008209f
C236 B.n191 VSUBS 0.008209f
C237 B.n192 VSUBS 0.008209f
C238 B.n193 VSUBS 0.019444f
C239 B.n194 VSUBS 0.019186f
C240 B.n195 VSUBS 0.019186f
C241 B.n196 VSUBS 0.008209f
C242 B.n197 VSUBS 0.008209f
C243 B.n198 VSUBS 0.008209f
C244 B.n199 VSUBS 0.008209f
C245 B.n200 VSUBS 0.008209f
C246 B.n201 VSUBS 0.008209f
C247 B.n202 VSUBS 0.008209f
C248 B.n203 VSUBS 0.008209f
C249 B.n204 VSUBS 0.008209f
C250 B.n205 VSUBS 0.008209f
C251 B.n206 VSUBS 0.008209f
C252 B.n207 VSUBS 0.008209f
C253 B.n208 VSUBS 0.008209f
C254 B.n209 VSUBS 0.008209f
C255 B.n210 VSUBS 0.008209f
C256 B.n211 VSUBS 0.008209f
C257 B.n212 VSUBS 0.008209f
C258 B.n213 VSUBS 0.008209f
C259 B.n214 VSUBS 0.008209f
C260 B.n215 VSUBS 0.008209f
C261 B.n216 VSUBS 0.008209f
C262 B.n217 VSUBS 0.008209f
C263 B.n218 VSUBS 0.008209f
C264 B.n219 VSUBS 0.008209f
C265 B.n220 VSUBS 0.008209f
C266 B.n221 VSUBS 0.008209f
C267 B.n222 VSUBS 0.008209f
C268 B.n223 VSUBS 0.008209f
C269 B.n224 VSUBS 0.008209f
C270 B.n225 VSUBS 0.008209f
C271 B.n226 VSUBS 0.008209f
C272 B.n227 VSUBS 0.008209f
C273 B.n228 VSUBS 0.008209f
C274 B.n229 VSUBS 0.008209f
C275 B.n230 VSUBS 0.008209f
C276 B.n231 VSUBS 0.008209f
C277 B.n232 VSUBS 0.008209f
C278 B.n233 VSUBS 0.008209f
C279 B.n234 VSUBS 0.008209f
C280 B.n235 VSUBS 0.008209f
C281 B.n236 VSUBS 0.008209f
C282 B.n237 VSUBS 0.008209f
C283 B.n238 VSUBS 0.008209f
C284 B.n239 VSUBS 0.008209f
C285 B.n240 VSUBS 0.008209f
C286 B.n241 VSUBS 0.008209f
C287 B.n242 VSUBS 0.008209f
C288 B.n243 VSUBS 0.008209f
C289 B.n244 VSUBS 0.008209f
C290 B.n245 VSUBS 0.008209f
C291 B.n246 VSUBS 0.008209f
C292 B.n247 VSUBS 0.008209f
C293 B.n248 VSUBS 0.008209f
C294 B.n249 VSUBS 0.008209f
C295 B.n250 VSUBS 0.008209f
C296 B.n251 VSUBS 0.008209f
C297 B.n252 VSUBS 0.008209f
C298 B.n253 VSUBS 0.008209f
C299 B.n254 VSUBS 0.008209f
C300 B.n255 VSUBS 0.008209f
C301 B.n256 VSUBS 0.008209f
C302 B.n257 VSUBS 0.008209f
C303 B.n258 VSUBS 0.008209f
C304 B.n259 VSUBS 0.008209f
C305 B.n260 VSUBS 0.008209f
C306 B.n261 VSUBS 0.008209f
C307 B.n262 VSUBS 0.008209f
C308 B.n263 VSUBS 0.008209f
C309 B.n264 VSUBS 0.008209f
C310 B.n265 VSUBS 0.008209f
C311 B.n266 VSUBS 0.008209f
C312 B.n267 VSUBS 0.008209f
C313 B.n268 VSUBS 0.008209f
C314 B.n269 VSUBS 0.019186f
C315 B.n270 VSUBS 0.020147f
C316 B.n271 VSUBS 0.018482f
C317 B.n272 VSUBS 0.008209f
C318 B.n273 VSUBS 0.008209f
C319 B.n274 VSUBS 0.008209f
C320 B.n275 VSUBS 0.008209f
C321 B.n276 VSUBS 0.008209f
C322 B.n277 VSUBS 0.008209f
C323 B.n278 VSUBS 0.008209f
C324 B.n279 VSUBS 0.008209f
C325 B.n280 VSUBS 0.008209f
C326 B.n281 VSUBS 0.008209f
C327 B.n282 VSUBS 0.008209f
C328 B.n283 VSUBS 0.008209f
C329 B.n284 VSUBS 0.008209f
C330 B.n285 VSUBS 0.008209f
C331 B.n286 VSUBS 0.008209f
C332 B.n287 VSUBS 0.008209f
C333 B.n288 VSUBS 0.008209f
C334 B.n289 VSUBS 0.008209f
C335 B.n290 VSUBS 0.007726f
C336 B.n291 VSUBS 0.008209f
C337 B.n292 VSUBS 0.008209f
C338 B.n293 VSUBS 0.008209f
C339 B.n294 VSUBS 0.008209f
C340 B.n295 VSUBS 0.008209f
C341 B.n296 VSUBS 0.008209f
C342 B.n297 VSUBS 0.008209f
C343 B.n298 VSUBS 0.008209f
C344 B.n299 VSUBS 0.008209f
C345 B.n300 VSUBS 0.008209f
C346 B.n301 VSUBS 0.008209f
C347 B.n302 VSUBS 0.008209f
C348 B.n303 VSUBS 0.008209f
C349 B.n304 VSUBS 0.008209f
C350 B.n305 VSUBS 0.008209f
C351 B.n306 VSUBS 0.004587f
C352 B.n307 VSUBS 0.019019f
C353 B.n308 VSUBS 0.007726f
C354 B.n309 VSUBS 0.008209f
C355 B.n310 VSUBS 0.008209f
C356 B.n311 VSUBS 0.008209f
C357 B.n312 VSUBS 0.008209f
C358 B.n313 VSUBS 0.008209f
C359 B.n314 VSUBS 0.008209f
C360 B.n315 VSUBS 0.008209f
C361 B.n316 VSUBS 0.008209f
C362 B.n317 VSUBS 0.008209f
C363 B.n318 VSUBS 0.008209f
C364 B.n319 VSUBS 0.008209f
C365 B.n320 VSUBS 0.008209f
C366 B.n321 VSUBS 0.008209f
C367 B.n322 VSUBS 0.008209f
C368 B.n323 VSUBS 0.008209f
C369 B.n324 VSUBS 0.008209f
C370 B.n325 VSUBS 0.008209f
C371 B.n326 VSUBS 0.008209f
C372 B.n327 VSUBS 0.019444f
C373 B.n328 VSUBS 0.019444f
C374 B.n329 VSUBS 0.019186f
C375 B.n330 VSUBS 0.008209f
C376 B.n331 VSUBS 0.008209f
C377 B.n332 VSUBS 0.008209f
C378 B.n333 VSUBS 0.008209f
C379 B.n334 VSUBS 0.008209f
C380 B.n335 VSUBS 0.008209f
C381 B.n336 VSUBS 0.008209f
C382 B.n337 VSUBS 0.008209f
C383 B.n338 VSUBS 0.008209f
C384 B.n339 VSUBS 0.008209f
C385 B.n340 VSUBS 0.008209f
C386 B.n341 VSUBS 0.008209f
C387 B.n342 VSUBS 0.008209f
C388 B.n343 VSUBS 0.008209f
C389 B.n344 VSUBS 0.008209f
C390 B.n345 VSUBS 0.008209f
C391 B.n346 VSUBS 0.008209f
C392 B.n347 VSUBS 0.008209f
C393 B.n348 VSUBS 0.008209f
C394 B.n349 VSUBS 0.008209f
C395 B.n350 VSUBS 0.008209f
C396 B.n351 VSUBS 0.008209f
C397 B.n352 VSUBS 0.008209f
C398 B.n353 VSUBS 0.008209f
C399 B.n354 VSUBS 0.008209f
C400 B.n355 VSUBS 0.008209f
C401 B.n356 VSUBS 0.008209f
C402 B.n357 VSUBS 0.008209f
C403 B.n358 VSUBS 0.008209f
C404 B.n359 VSUBS 0.008209f
C405 B.n360 VSUBS 0.008209f
C406 B.n361 VSUBS 0.008209f
C407 B.n362 VSUBS 0.008209f
C408 B.n363 VSUBS 0.008209f
C409 B.n364 VSUBS 0.008209f
C410 B.n365 VSUBS 0.008209f
C411 B.n366 VSUBS 0.008209f
C412 B.n367 VSUBS 0.018587f
C413 VDD1.t1 VSUBS 0.25629f
C414 VDD1.t0 VSUBS 0.407494f
C415 VTAIL.t2 VSUBS 0.279496f
C416 VTAIL.n0 VSUBS 1.06277f
C417 VTAIL.t1 VSUBS 0.279497f
C418 VTAIL.n1 VSUBS 1.09769f
C419 VTAIL.t3 VSUBS 0.279496f
C420 VTAIL.n2 VSUBS 0.943311f
C421 VTAIL.t0 VSUBS 0.279496f
C422 VTAIL.n3 VSUBS 0.871419f
C423 VP.t0 VSUBS 1.94641f
C424 VP.t1 VSUBS 1.26423f
C425 VP.n0 VSUBS 3.37778f
.ends

