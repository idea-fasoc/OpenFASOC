* NGSPICE file created from diff_pair_sample_1305.ext - technology: sky130A

.subckt diff_pair_sample_1305 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t1 VN.t0 VTAIL.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=6.513 pd=34.18 as=6.513 ps=34.18 w=16.7 l=0.5
X1 B.t15 B.t13 B.t14 B.t10 sky130_fd_pr__nfet_01v8 ad=6.513 pd=34.18 as=0 ps=0 w=16.7 l=0.5
X2 B.t12 B.t9 B.t11 B.t10 sky130_fd_pr__nfet_01v8 ad=6.513 pd=34.18 as=0 ps=0 w=16.7 l=0.5
X3 VDD1.t1 VP.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=6.513 pd=34.18 as=6.513 ps=34.18 w=16.7 l=0.5
X4 B.t8 B.t6 B.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=6.513 pd=34.18 as=0 ps=0 w=16.7 l=0.5
X5 VDD2.t0 VN.t1 VTAIL.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=6.513 pd=34.18 as=6.513 ps=34.18 w=16.7 l=0.5
X6 VDD1.t0 VP.t1 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=6.513 pd=34.18 as=6.513 ps=34.18 w=16.7 l=0.5
X7 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=6.513 pd=34.18 as=0 ps=0 w=16.7 l=0.5
R0 VN VN.t0 1087.85
R1 VN VN.t1 1044.86
R2 VTAIL.n370 VTAIL.n282 289.615
R3 VTAIL.n88 VTAIL.n0 289.615
R4 VTAIL.n276 VTAIL.n188 289.615
R5 VTAIL.n182 VTAIL.n94 289.615
R6 VTAIL.n313 VTAIL.n312 185
R7 VTAIL.n310 VTAIL.n309 185
R8 VTAIL.n319 VTAIL.n318 185
R9 VTAIL.n321 VTAIL.n320 185
R10 VTAIL.n306 VTAIL.n305 185
R11 VTAIL.n327 VTAIL.n326 185
R12 VTAIL.n329 VTAIL.n328 185
R13 VTAIL.n302 VTAIL.n301 185
R14 VTAIL.n335 VTAIL.n334 185
R15 VTAIL.n337 VTAIL.n336 185
R16 VTAIL.n298 VTAIL.n297 185
R17 VTAIL.n343 VTAIL.n342 185
R18 VTAIL.n345 VTAIL.n344 185
R19 VTAIL.n294 VTAIL.n293 185
R20 VTAIL.n351 VTAIL.n350 185
R21 VTAIL.n354 VTAIL.n353 185
R22 VTAIL.n352 VTAIL.n290 185
R23 VTAIL.n359 VTAIL.n289 185
R24 VTAIL.n361 VTAIL.n360 185
R25 VTAIL.n363 VTAIL.n362 185
R26 VTAIL.n286 VTAIL.n285 185
R27 VTAIL.n369 VTAIL.n368 185
R28 VTAIL.n371 VTAIL.n370 185
R29 VTAIL.n31 VTAIL.n30 185
R30 VTAIL.n28 VTAIL.n27 185
R31 VTAIL.n37 VTAIL.n36 185
R32 VTAIL.n39 VTAIL.n38 185
R33 VTAIL.n24 VTAIL.n23 185
R34 VTAIL.n45 VTAIL.n44 185
R35 VTAIL.n47 VTAIL.n46 185
R36 VTAIL.n20 VTAIL.n19 185
R37 VTAIL.n53 VTAIL.n52 185
R38 VTAIL.n55 VTAIL.n54 185
R39 VTAIL.n16 VTAIL.n15 185
R40 VTAIL.n61 VTAIL.n60 185
R41 VTAIL.n63 VTAIL.n62 185
R42 VTAIL.n12 VTAIL.n11 185
R43 VTAIL.n69 VTAIL.n68 185
R44 VTAIL.n72 VTAIL.n71 185
R45 VTAIL.n70 VTAIL.n8 185
R46 VTAIL.n77 VTAIL.n7 185
R47 VTAIL.n79 VTAIL.n78 185
R48 VTAIL.n81 VTAIL.n80 185
R49 VTAIL.n4 VTAIL.n3 185
R50 VTAIL.n87 VTAIL.n86 185
R51 VTAIL.n89 VTAIL.n88 185
R52 VTAIL.n277 VTAIL.n276 185
R53 VTAIL.n275 VTAIL.n274 185
R54 VTAIL.n192 VTAIL.n191 185
R55 VTAIL.n269 VTAIL.n268 185
R56 VTAIL.n267 VTAIL.n266 185
R57 VTAIL.n265 VTAIL.n195 185
R58 VTAIL.n199 VTAIL.n196 185
R59 VTAIL.n260 VTAIL.n259 185
R60 VTAIL.n258 VTAIL.n257 185
R61 VTAIL.n201 VTAIL.n200 185
R62 VTAIL.n252 VTAIL.n251 185
R63 VTAIL.n250 VTAIL.n249 185
R64 VTAIL.n205 VTAIL.n204 185
R65 VTAIL.n244 VTAIL.n243 185
R66 VTAIL.n242 VTAIL.n241 185
R67 VTAIL.n209 VTAIL.n208 185
R68 VTAIL.n236 VTAIL.n235 185
R69 VTAIL.n234 VTAIL.n233 185
R70 VTAIL.n213 VTAIL.n212 185
R71 VTAIL.n228 VTAIL.n227 185
R72 VTAIL.n226 VTAIL.n225 185
R73 VTAIL.n217 VTAIL.n216 185
R74 VTAIL.n220 VTAIL.n219 185
R75 VTAIL.n183 VTAIL.n182 185
R76 VTAIL.n181 VTAIL.n180 185
R77 VTAIL.n98 VTAIL.n97 185
R78 VTAIL.n175 VTAIL.n174 185
R79 VTAIL.n173 VTAIL.n172 185
R80 VTAIL.n171 VTAIL.n101 185
R81 VTAIL.n105 VTAIL.n102 185
R82 VTAIL.n166 VTAIL.n165 185
R83 VTAIL.n164 VTAIL.n163 185
R84 VTAIL.n107 VTAIL.n106 185
R85 VTAIL.n158 VTAIL.n157 185
R86 VTAIL.n156 VTAIL.n155 185
R87 VTAIL.n111 VTAIL.n110 185
R88 VTAIL.n150 VTAIL.n149 185
R89 VTAIL.n148 VTAIL.n147 185
R90 VTAIL.n115 VTAIL.n114 185
R91 VTAIL.n142 VTAIL.n141 185
R92 VTAIL.n140 VTAIL.n139 185
R93 VTAIL.n119 VTAIL.n118 185
R94 VTAIL.n134 VTAIL.n133 185
R95 VTAIL.n132 VTAIL.n131 185
R96 VTAIL.n123 VTAIL.n122 185
R97 VTAIL.n126 VTAIL.n125 185
R98 VTAIL.t3 VTAIL.n218 147.659
R99 VTAIL.t1 VTAIL.n124 147.659
R100 VTAIL.t2 VTAIL.n311 147.659
R101 VTAIL.t0 VTAIL.n29 147.659
R102 VTAIL.n312 VTAIL.n309 104.615
R103 VTAIL.n319 VTAIL.n309 104.615
R104 VTAIL.n320 VTAIL.n319 104.615
R105 VTAIL.n320 VTAIL.n305 104.615
R106 VTAIL.n327 VTAIL.n305 104.615
R107 VTAIL.n328 VTAIL.n327 104.615
R108 VTAIL.n328 VTAIL.n301 104.615
R109 VTAIL.n335 VTAIL.n301 104.615
R110 VTAIL.n336 VTAIL.n335 104.615
R111 VTAIL.n336 VTAIL.n297 104.615
R112 VTAIL.n343 VTAIL.n297 104.615
R113 VTAIL.n344 VTAIL.n343 104.615
R114 VTAIL.n344 VTAIL.n293 104.615
R115 VTAIL.n351 VTAIL.n293 104.615
R116 VTAIL.n353 VTAIL.n351 104.615
R117 VTAIL.n353 VTAIL.n352 104.615
R118 VTAIL.n352 VTAIL.n289 104.615
R119 VTAIL.n361 VTAIL.n289 104.615
R120 VTAIL.n362 VTAIL.n361 104.615
R121 VTAIL.n362 VTAIL.n285 104.615
R122 VTAIL.n369 VTAIL.n285 104.615
R123 VTAIL.n370 VTAIL.n369 104.615
R124 VTAIL.n30 VTAIL.n27 104.615
R125 VTAIL.n37 VTAIL.n27 104.615
R126 VTAIL.n38 VTAIL.n37 104.615
R127 VTAIL.n38 VTAIL.n23 104.615
R128 VTAIL.n45 VTAIL.n23 104.615
R129 VTAIL.n46 VTAIL.n45 104.615
R130 VTAIL.n46 VTAIL.n19 104.615
R131 VTAIL.n53 VTAIL.n19 104.615
R132 VTAIL.n54 VTAIL.n53 104.615
R133 VTAIL.n54 VTAIL.n15 104.615
R134 VTAIL.n61 VTAIL.n15 104.615
R135 VTAIL.n62 VTAIL.n61 104.615
R136 VTAIL.n62 VTAIL.n11 104.615
R137 VTAIL.n69 VTAIL.n11 104.615
R138 VTAIL.n71 VTAIL.n69 104.615
R139 VTAIL.n71 VTAIL.n70 104.615
R140 VTAIL.n70 VTAIL.n7 104.615
R141 VTAIL.n79 VTAIL.n7 104.615
R142 VTAIL.n80 VTAIL.n79 104.615
R143 VTAIL.n80 VTAIL.n3 104.615
R144 VTAIL.n87 VTAIL.n3 104.615
R145 VTAIL.n88 VTAIL.n87 104.615
R146 VTAIL.n276 VTAIL.n275 104.615
R147 VTAIL.n275 VTAIL.n191 104.615
R148 VTAIL.n268 VTAIL.n191 104.615
R149 VTAIL.n268 VTAIL.n267 104.615
R150 VTAIL.n267 VTAIL.n195 104.615
R151 VTAIL.n199 VTAIL.n195 104.615
R152 VTAIL.n259 VTAIL.n199 104.615
R153 VTAIL.n259 VTAIL.n258 104.615
R154 VTAIL.n258 VTAIL.n200 104.615
R155 VTAIL.n251 VTAIL.n200 104.615
R156 VTAIL.n251 VTAIL.n250 104.615
R157 VTAIL.n250 VTAIL.n204 104.615
R158 VTAIL.n243 VTAIL.n204 104.615
R159 VTAIL.n243 VTAIL.n242 104.615
R160 VTAIL.n242 VTAIL.n208 104.615
R161 VTAIL.n235 VTAIL.n208 104.615
R162 VTAIL.n235 VTAIL.n234 104.615
R163 VTAIL.n234 VTAIL.n212 104.615
R164 VTAIL.n227 VTAIL.n212 104.615
R165 VTAIL.n227 VTAIL.n226 104.615
R166 VTAIL.n226 VTAIL.n216 104.615
R167 VTAIL.n219 VTAIL.n216 104.615
R168 VTAIL.n182 VTAIL.n181 104.615
R169 VTAIL.n181 VTAIL.n97 104.615
R170 VTAIL.n174 VTAIL.n97 104.615
R171 VTAIL.n174 VTAIL.n173 104.615
R172 VTAIL.n173 VTAIL.n101 104.615
R173 VTAIL.n105 VTAIL.n101 104.615
R174 VTAIL.n165 VTAIL.n105 104.615
R175 VTAIL.n165 VTAIL.n164 104.615
R176 VTAIL.n164 VTAIL.n106 104.615
R177 VTAIL.n157 VTAIL.n106 104.615
R178 VTAIL.n157 VTAIL.n156 104.615
R179 VTAIL.n156 VTAIL.n110 104.615
R180 VTAIL.n149 VTAIL.n110 104.615
R181 VTAIL.n149 VTAIL.n148 104.615
R182 VTAIL.n148 VTAIL.n114 104.615
R183 VTAIL.n141 VTAIL.n114 104.615
R184 VTAIL.n141 VTAIL.n140 104.615
R185 VTAIL.n140 VTAIL.n118 104.615
R186 VTAIL.n133 VTAIL.n118 104.615
R187 VTAIL.n133 VTAIL.n132 104.615
R188 VTAIL.n132 VTAIL.n122 104.615
R189 VTAIL.n125 VTAIL.n122 104.615
R190 VTAIL.n312 VTAIL.t2 52.3082
R191 VTAIL.n30 VTAIL.t0 52.3082
R192 VTAIL.n219 VTAIL.t3 52.3082
R193 VTAIL.n125 VTAIL.t1 52.3082
R194 VTAIL.n375 VTAIL.n374 30.246
R195 VTAIL.n93 VTAIL.n92 30.246
R196 VTAIL.n281 VTAIL.n280 30.246
R197 VTAIL.n187 VTAIL.n186 30.246
R198 VTAIL.n187 VTAIL.n93 28.2117
R199 VTAIL.n375 VTAIL.n281 27.4962
R200 VTAIL.n313 VTAIL.n311 15.6677
R201 VTAIL.n31 VTAIL.n29 15.6677
R202 VTAIL.n220 VTAIL.n218 15.6677
R203 VTAIL.n126 VTAIL.n124 15.6677
R204 VTAIL.n360 VTAIL.n359 13.1884
R205 VTAIL.n78 VTAIL.n77 13.1884
R206 VTAIL.n266 VTAIL.n265 13.1884
R207 VTAIL.n172 VTAIL.n171 13.1884
R208 VTAIL.n314 VTAIL.n310 12.8005
R209 VTAIL.n358 VTAIL.n290 12.8005
R210 VTAIL.n363 VTAIL.n288 12.8005
R211 VTAIL.n32 VTAIL.n28 12.8005
R212 VTAIL.n76 VTAIL.n8 12.8005
R213 VTAIL.n81 VTAIL.n6 12.8005
R214 VTAIL.n269 VTAIL.n194 12.8005
R215 VTAIL.n264 VTAIL.n196 12.8005
R216 VTAIL.n221 VTAIL.n217 12.8005
R217 VTAIL.n175 VTAIL.n100 12.8005
R218 VTAIL.n170 VTAIL.n102 12.8005
R219 VTAIL.n127 VTAIL.n123 12.8005
R220 VTAIL.n318 VTAIL.n317 12.0247
R221 VTAIL.n355 VTAIL.n354 12.0247
R222 VTAIL.n364 VTAIL.n286 12.0247
R223 VTAIL.n36 VTAIL.n35 12.0247
R224 VTAIL.n73 VTAIL.n72 12.0247
R225 VTAIL.n82 VTAIL.n4 12.0247
R226 VTAIL.n270 VTAIL.n192 12.0247
R227 VTAIL.n261 VTAIL.n260 12.0247
R228 VTAIL.n225 VTAIL.n224 12.0247
R229 VTAIL.n176 VTAIL.n98 12.0247
R230 VTAIL.n167 VTAIL.n166 12.0247
R231 VTAIL.n131 VTAIL.n130 12.0247
R232 VTAIL.n321 VTAIL.n308 11.249
R233 VTAIL.n350 VTAIL.n292 11.249
R234 VTAIL.n368 VTAIL.n367 11.249
R235 VTAIL.n39 VTAIL.n26 11.249
R236 VTAIL.n68 VTAIL.n10 11.249
R237 VTAIL.n86 VTAIL.n85 11.249
R238 VTAIL.n274 VTAIL.n273 11.249
R239 VTAIL.n257 VTAIL.n198 11.249
R240 VTAIL.n228 VTAIL.n215 11.249
R241 VTAIL.n180 VTAIL.n179 11.249
R242 VTAIL.n163 VTAIL.n104 11.249
R243 VTAIL.n134 VTAIL.n121 11.249
R244 VTAIL.n322 VTAIL.n306 10.4732
R245 VTAIL.n349 VTAIL.n294 10.4732
R246 VTAIL.n371 VTAIL.n284 10.4732
R247 VTAIL.n40 VTAIL.n24 10.4732
R248 VTAIL.n67 VTAIL.n12 10.4732
R249 VTAIL.n89 VTAIL.n2 10.4732
R250 VTAIL.n277 VTAIL.n190 10.4732
R251 VTAIL.n256 VTAIL.n201 10.4732
R252 VTAIL.n229 VTAIL.n213 10.4732
R253 VTAIL.n183 VTAIL.n96 10.4732
R254 VTAIL.n162 VTAIL.n107 10.4732
R255 VTAIL.n135 VTAIL.n119 10.4732
R256 VTAIL.n326 VTAIL.n325 9.69747
R257 VTAIL.n346 VTAIL.n345 9.69747
R258 VTAIL.n372 VTAIL.n282 9.69747
R259 VTAIL.n44 VTAIL.n43 9.69747
R260 VTAIL.n64 VTAIL.n63 9.69747
R261 VTAIL.n90 VTAIL.n0 9.69747
R262 VTAIL.n278 VTAIL.n188 9.69747
R263 VTAIL.n253 VTAIL.n252 9.69747
R264 VTAIL.n233 VTAIL.n232 9.69747
R265 VTAIL.n184 VTAIL.n94 9.69747
R266 VTAIL.n159 VTAIL.n158 9.69747
R267 VTAIL.n139 VTAIL.n138 9.69747
R268 VTAIL.n374 VTAIL.n373 9.45567
R269 VTAIL.n92 VTAIL.n91 9.45567
R270 VTAIL.n280 VTAIL.n279 9.45567
R271 VTAIL.n186 VTAIL.n185 9.45567
R272 VTAIL.n373 VTAIL.n372 9.3005
R273 VTAIL.n284 VTAIL.n283 9.3005
R274 VTAIL.n367 VTAIL.n366 9.3005
R275 VTAIL.n365 VTAIL.n364 9.3005
R276 VTAIL.n288 VTAIL.n287 9.3005
R277 VTAIL.n333 VTAIL.n332 9.3005
R278 VTAIL.n331 VTAIL.n330 9.3005
R279 VTAIL.n304 VTAIL.n303 9.3005
R280 VTAIL.n325 VTAIL.n324 9.3005
R281 VTAIL.n323 VTAIL.n322 9.3005
R282 VTAIL.n308 VTAIL.n307 9.3005
R283 VTAIL.n317 VTAIL.n316 9.3005
R284 VTAIL.n315 VTAIL.n314 9.3005
R285 VTAIL.n300 VTAIL.n299 9.3005
R286 VTAIL.n339 VTAIL.n338 9.3005
R287 VTAIL.n341 VTAIL.n340 9.3005
R288 VTAIL.n296 VTAIL.n295 9.3005
R289 VTAIL.n347 VTAIL.n346 9.3005
R290 VTAIL.n349 VTAIL.n348 9.3005
R291 VTAIL.n292 VTAIL.n291 9.3005
R292 VTAIL.n356 VTAIL.n355 9.3005
R293 VTAIL.n358 VTAIL.n357 9.3005
R294 VTAIL.n91 VTAIL.n90 9.3005
R295 VTAIL.n2 VTAIL.n1 9.3005
R296 VTAIL.n85 VTAIL.n84 9.3005
R297 VTAIL.n83 VTAIL.n82 9.3005
R298 VTAIL.n6 VTAIL.n5 9.3005
R299 VTAIL.n51 VTAIL.n50 9.3005
R300 VTAIL.n49 VTAIL.n48 9.3005
R301 VTAIL.n22 VTAIL.n21 9.3005
R302 VTAIL.n43 VTAIL.n42 9.3005
R303 VTAIL.n41 VTAIL.n40 9.3005
R304 VTAIL.n26 VTAIL.n25 9.3005
R305 VTAIL.n35 VTAIL.n34 9.3005
R306 VTAIL.n33 VTAIL.n32 9.3005
R307 VTAIL.n18 VTAIL.n17 9.3005
R308 VTAIL.n57 VTAIL.n56 9.3005
R309 VTAIL.n59 VTAIL.n58 9.3005
R310 VTAIL.n14 VTAIL.n13 9.3005
R311 VTAIL.n65 VTAIL.n64 9.3005
R312 VTAIL.n67 VTAIL.n66 9.3005
R313 VTAIL.n10 VTAIL.n9 9.3005
R314 VTAIL.n74 VTAIL.n73 9.3005
R315 VTAIL.n76 VTAIL.n75 9.3005
R316 VTAIL.n246 VTAIL.n245 9.3005
R317 VTAIL.n248 VTAIL.n247 9.3005
R318 VTAIL.n203 VTAIL.n202 9.3005
R319 VTAIL.n254 VTAIL.n253 9.3005
R320 VTAIL.n256 VTAIL.n255 9.3005
R321 VTAIL.n198 VTAIL.n197 9.3005
R322 VTAIL.n262 VTAIL.n261 9.3005
R323 VTAIL.n264 VTAIL.n263 9.3005
R324 VTAIL.n279 VTAIL.n278 9.3005
R325 VTAIL.n190 VTAIL.n189 9.3005
R326 VTAIL.n273 VTAIL.n272 9.3005
R327 VTAIL.n271 VTAIL.n270 9.3005
R328 VTAIL.n194 VTAIL.n193 9.3005
R329 VTAIL.n207 VTAIL.n206 9.3005
R330 VTAIL.n240 VTAIL.n239 9.3005
R331 VTAIL.n238 VTAIL.n237 9.3005
R332 VTAIL.n211 VTAIL.n210 9.3005
R333 VTAIL.n232 VTAIL.n231 9.3005
R334 VTAIL.n230 VTAIL.n229 9.3005
R335 VTAIL.n215 VTAIL.n214 9.3005
R336 VTAIL.n224 VTAIL.n223 9.3005
R337 VTAIL.n222 VTAIL.n221 9.3005
R338 VTAIL.n152 VTAIL.n151 9.3005
R339 VTAIL.n154 VTAIL.n153 9.3005
R340 VTAIL.n109 VTAIL.n108 9.3005
R341 VTAIL.n160 VTAIL.n159 9.3005
R342 VTAIL.n162 VTAIL.n161 9.3005
R343 VTAIL.n104 VTAIL.n103 9.3005
R344 VTAIL.n168 VTAIL.n167 9.3005
R345 VTAIL.n170 VTAIL.n169 9.3005
R346 VTAIL.n185 VTAIL.n184 9.3005
R347 VTAIL.n96 VTAIL.n95 9.3005
R348 VTAIL.n179 VTAIL.n178 9.3005
R349 VTAIL.n177 VTAIL.n176 9.3005
R350 VTAIL.n100 VTAIL.n99 9.3005
R351 VTAIL.n113 VTAIL.n112 9.3005
R352 VTAIL.n146 VTAIL.n145 9.3005
R353 VTAIL.n144 VTAIL.n143 9.3005
R354 VTAIL.n117 VTAIL.n116 9.3005
R355 VTAIL.n138 VTAIL.n137 9.3005
R356 VTAIL.n136 VTAIL.n135 9.3005
R357 VTAIL.n121 VTAIL.n120 9.3005
R358 VTAIL.n130 VTAIL.n129 9.3005
R359 VTAIL.n128 VTAIL.n127 9.3005
R360 VTAIL.n329 VTAIL.n304 8.92171
R361 VTAIL.n342 VTAIL.n296 8.92171
R362 VTAIL.n47 VTAIL.n22 8.92171
R363 VTAIL.n60 VTAIL.n14 8.92171
R364 VTAIL.n249 VTAIL.n203 8.92171
R365 VTAIL.n236 VTAIL.n211 8.92171
R366 VTAIL.n155 VTAIL.n109 8.92171
R367 VTAIL.n142 VTAIL.n117 8.92171
R368 VTAIL.n330 VTAIL.n302 8.14595
R369 VTAIL.n341 VTAIL.n298 8.14595
R370 VTAIL.n48 VTAIL.n20 8.14595
R371 VTAIL.n59 VTAIL.n16 8.14595
R372 VTAIL.n248 VTAIL.n205 8.14595
R373 VTAIL.n237 VTAIL.n209 8.14595
R374 VTAIL.n154 VTAIL.n111 8.14595
R375 VTAIL.n143 VTAIL.n115 8.14595
R376 VTAIL.n334 VTAIL.n333 7.3702
R377 VTAIL.n338 VTAIL.n337 7.3702
R378 VTAIL.n52 VTAIL.n51 7.3702
R379 VTAIL.n56 VTAIL.n55 7.3702
R380 VTAIL.n245 VTAIL.n244 7.3702
R381 VTAIL.n241 VTAIL.n240 7.3702
R382 VTAIL.n151 VTAIL.n150 7.3702
R383 VTAIL.n147 VTAIL.n146 7.3702
R384 VTAIL.n334 VTAIL.n300 6.59444
R385 VTAIL.n337 VTAIL.n300 6.59444
R386 VTAIL.n52 VTAIL.n18 6.59444
R387 VTAIL.n55 VTAIL.n18 6.59444
R388 VTAIL.n244 VTAIL.n207 6.59444
R389 VTAIL.n241 VTAIL.n207 6.59444
R390 VTAIL.n150 VTAIL.n113 6.59444
R391 VTAIL.n147 VTAIL.n113 6.59444
R392 VTAIL.n333 VTAIL.n302 5.81868
R393 VTAIL.n338 VTAIL.n298 5.81868
R394 VTAIL.n51 VTAIL.n20 5.81868
R395 VTAIL.n56 VTAIL.n16 5.81868
R396 VTAIL.n245 VTAIL.n205 5.81868
R397 VTAIL.n240 VTAIL.n209 5.81868
R398 VTAIL.n151 VTAIL.n111 5.81868
R399 VTAIL.n146 VTAIL.n115 5.81868
R400 VTAIL.n330 VTAIL.n329 5.04292
R401 VTAIL.n342 VTAIL.n341 5.04292
R402 VTAIL.n48 VTAIL.n47 5.04292
R403 VTAIL.n60 VTAIL.n59 5.04292
R404 VTAIL.n249 VTAIL.n248 5.04292
R405 VTAIL.n237 VTAIL.n236 5.04292
R406 VTAIL.n155 VTAIL.n154 5.04292
R407 VTAIL.n143 VTAIL.n142 5.04292
R408 VTAIL.n222 VTAIL.n218 4.38563
R409 VTAIL.n128 VTAIL.n124 4.38563
R410 VTAIL.n315 VTAIL.n311 4.38563
R411 VTAIL.n33 VTAIL.n29 4.38563
R412 VTAIL.n326 VTAIL.n304 4.26717
R413 VTAIL.n345 VTAIL.n296 4.26717
R414 VTAIL.n374 VTAIL.n282 4.26717
R415 VTAIL.n44 VTAIL.n22 4.26717
R416 VTAIL.n63 VTAIL.n14 4.26717
R417 VTAIL.n92 VTAIL.n0 4.26717
R418 VTAIL.n280 VTAIL.n188 4.26717
R419 VTAIL.n252 VTAIL.n203 4.26717
R420 VTAIL.n233 VTAIL.n211 4.26717
R421 VTAIL.n186 VTAIL.n94 4.26717
R422 VTAIL.n158 VTAIL.n109 4.26717
R423 VTAIL.n139 VTAIL.n117 4.26717
R424 VTAIL.n325 VTAIL.n306 3.49141
R425 VTAIL.n346 VTAIL.n294 3.49141
R426 VTAIL.n372 VTAIL.n371 3.49141
R427 VTAIL.n43 VTAIL.n24 3.49141
R428 VTAIL.n64 VTAIL.n12 3.49141
R429 VTAIL.n90 VTAIL.n89 3.49141
R430 VTAIL.n278 VTAIL.n277 3.49141
R431 VTAIL.n253 VTAIL.n201 3.49141
R432 VTAIL.n232 VTAIL.n213 3.49141
R433 VTAIL.n184 VTAIL.n183 3.49141
R434 VTAIL.n159 VTAIL.n107 3.49141
R435 VTAIL.n138 VTAIL.n119 3.49141
R436 VTAIL.n322 VTAIL.n321 2.71565
R437 VTAIL.n350 VTAIL.n349 2.71565
R438 VTAIL.n368 VTAIL.n284 2.71565
R439 VTAIL.n40 VTAIL.n39 2.71565
R440 VTAIL.n68 VTAIL.n67 2.71565
R441 VTAIL.n86 VTAIL.n2 2.71565
R442 VTAIL.n274 VTAIL.n190 2.71565
R443 VTAIL.n257 VTAIL.n256 2.71565
R444 VTAIL.n229 VTAIL.n228 2.71565
R445 VTAIL.n180 VTAIL.n96 2.71565
R446 VTAIL.n163 VTAIL.n162 2.71565
R447 VTAIL.n135 VTAIL.n134 2.71565
R448 VTAIL.n318 VTAIL.n308 1.93989
R449 VTAIL.n354 VTAIL.n292 1.93989
R450 VTAIL.n367 VTAIL.n286 1.93989
R451 VTAIL.n36 VTAIL.n26 1.93989
R452 VTAIL.n72 VTAIL.n10 1.93989
R453 VTAIL.n85 VTAIL.n4 1.93989
R454 VTAIL.n273 VTAIL.n192 1.93989
R455 VTAIL.n260 VTAIL.n198 1.93989
R456 VTAIL.n225 VTAIL.n215 1.93989
R457 VTAIL.n179 VTAIL.n98 1.93989
R458 VTAIL.n166 VTAIL.n104 1.93989
R459 VTAIL.n131 VTAIL.n121 1.93989
R460 VTAIL.n317 VTAIL.n310 1.16414
R461 VTAIL.n355 VTAIL.n290 1.16414
R462 VTAIL.n364 VTAIL.n363 1.16414
R463 VTAIL.n35 VTAIL.n28 1.16414
R464 VTAIL.n73 VTAIL.n8 1.16414
R465 VTAIL.n82 VTAIL.n81 1.16414
R466 VTAIL.n270 VTAIL.n269 1.16414
R467 VTAIL.n261 VTAIL.n196 1.16414
R468 VTAIL.n224 VTAIL.n217 1.16414
R469 VTAIL.n176 VTAIL.n175 1.16414
R470 VTAIL.n167 VTAIL.n102 1.16414
R471 VTAIL.n130 VTAIL.n123 1.16414
R472 VTAIL.n281 VTAIL.n187 0.828086
R473 VTAIL VTAIL.n93 0.707397
R474 VTAIL.n314 VTAIL.n313 0.388379
R475 VTAIL.n359 VTAIL.n358 0.388379
R476 VTAIL.n360 VTAIL.n288 0.388379
R477 VTAIL.n32 VTAIL.n31 0.388379
R478 VTAIL.n77 VTAIL.n76 0.388379
R479 VTAIL.n78 VTAIL.n6 0.388379
R480 VTAIL.n266 VTAIL.n194 0.388379
R481 VTAIL.n265 VTAIL.n264 0.388379
R482 VTAIL.n221 VTAIL.n220 0.388379
R483 VTAIL.n172 VTAIL.n100 0.388379
R484 VTAIL.n171 VTAIL.n170 0.388379
R485 VTAIL.n127 VTAIL.n126 0.388379
R486 VTAIL.n316 VTAIL.n315 0.155672
R487 VTAIL.n316 VTAIL.n307 0.155672
R488 VTAIL.n323 VTAIL.n307 0.155672
R489 VTAIL.n324 VTAIL.n323 0.155672
R490 VTAIL.n324 VTAIL.n303 0.155672
R491 VTAIL.n331 VTAIL.n303 0.155672
R492 VTAIL.n332 VTAIL.n331 0.155672
R493 VTAIL.n332 VTAIL.n299 0.155672
R494 VTAIL.n339 VTAIL.n299 0.155672
R495 VTAIL.n340 VTAIL.n339 0.155672
R496 VTAIL.n340 VTAIL.n295 0.155672
R497 VTAIL.n347 VTAIL.n295 0.155672
R498 VTAIL.n348 VTAIL.n347 0.155672
R499 VTAIL.n348 VTAIL.n291 0.155672
R500 VTAIL.n356 VTAIL.n291 0.155672
R501 VTAIL.n357 VTAIL.n356 0.155672
R502 VTAIL.n357 VTAIL.n287 0.155672
R503 VTAIL.n365 VTAIL.n287 0.155672
R504 VTAIL.n366 VTAIL.n365 0.155672
R505 VTAIL.n366 VTAIL.n283 0.155672
R506 VTAIL.n373 VTAIL.n283 0.155672
R507 VTAIL.n34 VTAIL.n33 0.155672
R508 VTAIL.n34 VTAIL.n25 0.155672
R509 VTAIL.n41 VTAIL.n25 0.155672
R510 VTAIL.n42 VTAIL.n41 0.155672
R511 VTAIL.n42 VTAIL.n21 0.155672
R512 VTAIL.n49 VTAIL.n21 0.155672
R513 VTAIL.n50 VTAIL.n49 0.155672
R514 VTAIL.n50 VTAIL.n17 0.155672
R515 VTAIL.n57 VTAIL.n17 0.155672
R516 VTAIL.n58 VTAIL.n57 0.155672
R517 VTAIL.n58 VTAIL.n13 0.155672
R518 VTAIL.n65 VTAIL.n13 0.155672
R519 VTAIL.n66 VTAIL.n65 0.155672
R520 VTAIL.n66 VTAIL.n9 0.155672
R521 VTAIL.n74 VTAIL.n9 0.155672
R522 VTAIL.n75 VTAIL.n74 0.155672
R523 VTAIL.n75 VTAIL.n5 0.155672
R524 VTAIL.n83 VTAIL.n5 0.155672
R525 VTAIL.n84 VTAIL.n83 0.155672
R526 VTAIL.n84 VTAIL.n1 0.155672
R527 VTAIL.n91 VTAIL.n1 0.155672
R528 VTAIL.n279 VTAIL.n189 0.155672
R529 VTAIL.n272 VTAIL.n189 0.155672
R530 VTAIL.n272 VTAIL.n271 0.155672
R531 VTAIL.n271 VTAIL.n193 0.155672
R532 VTAIL.n263 VTAIL.n193 0.155672
R533 VTAIL.n263 VTAIL.n262 0.155672
R534 VTAIL.n262 VTAIL.n197 0.155672
R535 VTAIL.n255 VTAIL.n197 0.155672
R536 VTAIL.n255 VTAIL.n254 0.155672
R537 VTAIL.n254 VTAIL.n202 0.155672
R538 VTAIL.n247 VTAIL.n202 0.155672
R539 VTAIL.n247 VTAIL.n246 0.155672
R540 VTAIL.n246 VTAIL.n206 0.155672
R541 VTAIL.n239 VTAIL.n206 0.155672
R542 VTAIL.n239 VTAIL.n238 0.155672
R543 VTAIL.n238 VTAIL.n210 0.155672
R544 VTAIL.n231 VTAIL.n210 0.155672
R545 VTAIL.n231 VTAIL.n230 0.155672
R546 VTAIL.n230 VTAIL.n214 0.155672
R547 VTAIL.n223 VTAIL.n214 0.155672
R548 VTAIL.n223 VTAIL.n222 0.155672
R549 VTAIL.n185 VTAIL.n95 0.155672
R550 VTAIL.n178 VTAIL.n95 0.155672
R551 VTAIL.n178 VTAIL.n177 0.155672
R552 VTAIL.n177 VTAIL.n99 0.155672
R553 VTAIL.n169 VTAIL.n99 0.155672
R554 VTAIL.n169 VTAIL.n168 0.155672
R555 VTAIL.n168 VTAIL.n103 0.155672
R556 VTAIL.n161 VTAIL.n103 0.155672
R557 VTAIL.n161 VTAIL.n160 0.155672
R558 VTAIL.n160 VTAIL.n108 0.155672
R559 VTAIL.n153 VTAIL.n108 0.155672
R560 VTAIL.n153 VTAIL.n152 0.155672
R561 VTAIL.n152 VTAIL.n112 0.155672
R562 VTAIL.n145 VTAIL.n112 0.155672
R563 VTAIL.n145 VTAIL.n144 0.155672
R564 VTAIL.n144 VTAIL.n116 0.155672
R565 VTAIL.n137 VTAIL.n116 0.155672
R566 VTAIL.n137 VTAIL.n136 0.155672
R567 VTAIL.n136 VTAIL.n120 0.155672
R568 VTAIL.n129 VTAIL.n120 0.155672
R569 VTAIL.n129 VTAIL.n128 0.155672
R570 VTAIL VTAIL.n375 0.12119
R571 VDD2.n181 VDD2.n93 289.615
R572 VDD2.n88 VDD2.n0 289.615
R573 VDD2.n182 VDD2.n181 185
R574 VDD2.n180 VDD2.n179 185
R575 VDD2.n97 VDD2.n96 185
R576 VDD2.n174 VDD2.n173 185
R577 VDD2.n172 VDD2.n171 185
R578 VDD2.n170 VDD2.n100 185
R579 VDD2.n104 VDD2.n101 185
R580 VDD2.n165 VDD2.n164 185
R581 VDD2.n163 VDD2.n162 185
R582 VDD2.n106 VDD2.n105 185
R583 VDD2.n157 VDD2.n156 185
R584 VDD2.n155 VDD2.n154 185
R585 VDD2.n110 VDD2.n109 185
R586 VDD2.n149 VDD2.n148 185
R587 VDD2.n147 VDD2.n146 185
R588 VDD2.n114 VDD2.n113 185
R589 VDD2.n141 VDD2.n140 185
R590 VDD2.n139 VDD2.n138 185
R591 VDD2.n118 VDD2.n117 185
R592 VDD2.n133 VDD2.n132 185
R593 VDD2.n131 VDD2.n130 185
R594 VDD2.n122 VDD2.n121 185
R595 VDD2.n125 VDD2.n124 185
R596 VDD2.n31 VDD2.n30 185
R597 VDD2.n28 VDD2.n27 185
R598 VDD2.n37 VDD2.n36 185
R599 VDD2.n39 VDD2.n38 185
R600 VDD2.n24 VDD2.n23 185
R601 VDD2.n45 VDD2.n44 185
R602 VDD2.n47 VDD2.n46 185
R603 VDD2.n20 VDD2.n19 185
R604 VDD2.n53 VDD2.n52 185
R605 VDD2.n55 VDD2.n54 185
R606 VDD2.n16 VDD2.n15 185
R607 VDD2.n61 VDD2.n60 185
R608 VDD2.n63 VDD2.n62 185
R609 VDD2.n12 VDD2.n11 185
R610 VDD2.n69 VDD2.n68 185
R611 VDD2.n72 VDD2.n71 185
R612 VDD2.n70 VDD2.n8 185
R613 VDD2.n77 VDD2.n7 185
R614 VDD2.n79 VDD2.n78 185
R615 VDD2.n81 VDD2.n80 185
R616 VDD2.n4 VDD2.n3 185
R617 VDD2.n87 VDD2.n86 185
R618 VDD2.n89 VDD2.n88 185
R619 VDD2.t1 VDD2.n123 147.659
R620 VDD2.t0 VDD2.n29 147.659
R621 VDD2.n181 VDD2.n180 104.615
R622 VDD2.n180 VDD2.n96 104.615
R623 VDD2.n173 VDD2.n96 104.615
R624 VDD2.n173 VDD2.n172 104.615
R625 VDD2.n172 VDD2.n100 104.615
R626 VDD2.n104 VDD2.n100 104.615
R627 VDD2.n164 VDD2.n104 104.615
R628 VDD2.n164 VDD2.n163 104.615
R629 VDD2.n163 VDD2.n105 104.615
R630 VDD2.n156 VDD2.n105 104.615
R631 VDD2.n156 VDD2.n155 104.615
R632 VDD2.n155 VDD2.n109 104.615
R633 VDD2.n148 VDD2.n109 104.615
R634 VDD2.n148 VDD2.n147 104.615
R635 VDD2.n147 VDD2.n113 104.615
R636 VDD2.n140 VDD2.n113 104.615
R637 VDD2.n140 VDD2.n139 104.615
R638 VDD2.n139 VDD2.n117 104.615
R639 VDD2.n132 VDD2.n117 104.615
R640 VDD2.n132 VDD2.n131 104.615
R641 VDD2.n131 VDD2.n121 104.615
R642 VDD2.n124 VDD2.n121 104.615
R643 VDD2.n30 VDD2.n27 104.615
R644 VDD2.n37 VDD2.n27 104.615
R645 VDD2.n38 VDD2.n37 104.615
R646 VDD2.n38 VDD2.n23 104.615
R647 VDD2.n45 VDD2.n23 104.615
R648 VDD2.n46 VDD2.n45 104.615
R649 VDD2.n46 VDD2.n19 104.615
R650 VDD2.n53 VDD2.n19 104.615
R651 VDD2.n54 VDD2.n53 104.615
R652 VDD2.n54 VDD2.n15 104.615
R653 VDD2.n61 VDD2.n15 104.615
R654 VDD2.n62 VDD2.n61 104.615
R655 VDD2.n62 VDD2.n11 104.615
R656 VDD2.n69 VDD2.n11 104.615
R657 VDD2.n71 VDD2.n69 104.615
R658 VDD2.n71 VDD2.n70 104.615
R659 VDD2.n70 VDD2.n7 104.615
R660 VDD2.n79 VDD2.n7 104.615
R661 VDD2.n80 VDD2.n79 104.615
R662 VDD2.n80 VDD2.n3 104.615
R663 VDD2.n87 VDD2.n3 104.615
R664 VDD2.n88 VDD2.n87 104.615
R665 VDD2.n186 VDD2.n92 86.429
R666 VDD2.n124 VDD2.t1 52.3082
R667 VDD2.n30 VDD2.t0 52.3082
R668 VDD2.n186 VDD2.n185 46.9247
R669 VDD2.n125 VDD2.n123 15.6677
R670 VDD2.n31 VDD2.n29 15.6677
R671 VDD2.n171 VDD2.n170 13.1884
R672 VDD2.n78 VDD2.n77 13.1884
R673 VDD2.n174 VDD2.n99 12.8005
R674 VDD2.n169 VDD2.n101 12.8005
R675 VDD2.n126 VDD2.n122 12.8005
R676 VDD2.n32 VDD2.n28 12.8005
R677 VDD2.n76 VDD2.n8 12.8005
R678 VDD2.n81 VDD2.n6 12.8005
R679 VDD2.n175 VDD2.n97 12.0247
R680 VDD2.n166 VDD2.n165 12.0247
R681 VDD2.n130 VDD2.n129 12.0247
R682 VDD2.n36 VDD2.n35 12.0247
R683 VDD2.n73 VDD2.n72 12.0247
R684 VDD2.n82 VDD2.n4 12.0247
R685 VDD2.n179 VDD2.n178 11.249
R686 VDD2.n162 VDD2.n103 11.249
R687 VDD2.n133 VDD2.n120 11.249
R688 VDD2.n39 VDD2.n26 11.249
R689 VDD2.n68 VDD2.n10 11.249
R690 VDD2.n86 VDD2.n85 11.249
R691 VDD2.n182 VDD2.n95 10.4732
R692 VDD2.n161 VDD2.n106 10.4732
R693 VDD2.n134 VDD2.n118 10.4732
R694 VDD2.n40 VDD2.n24 10.4732
R695 VDD2.n67 VDD2.n12 10.4732
R696 VDD2.n89 VDD2.n2 10.4732
R697 VDD2.n183 VDD2.n93 9.69747
R698 VDD2.n158 VDD2.n157 9.69747
R699 VDD2.n138 VDD2.n137 9.69747
R700 VDD2.n44 VDD2.n43 9.69747
R701 VDD2.n64 VDD2.n63 9.69747
R702 VDD2.n90 VDD2.n0 9.69747
R703 VDD2.n185 VDD2.n184 9.45567
R704 VDD2.n92 VDD2.n91 9.45567
R705 VDD2.n151 VDD2.n150 9.3005
R706 VDD2.n153 VDD2.n152 9.3005
R707 VDD2.n108 VDD2.n107 9.3005
R708 VDD2.n159 VDD2.n158 9.3005
R709 VDD2.n161 VDD2.n160 9.3005
R710 VDD2.n103 VDD2.n102 9.3005
R711 VDD2.n167 VDD2.n166 9.3005
R712 VDD2.n169 VDD2.n168 9.3005
R713 VDD2.n184 VDD2.n183 9.3005
R714 VDD2.n95 VDD2.n94 9.3005
R715 VDD2.n178 VDD2.n177 9.3005
R716 VDD2.n176 VDD2.n175 9.3005
R717 VDD2.n99 VDD2.n98 9.3005
R718 VDD2.n112 VDD2.n111 9.3005
R719 VDD2.n145 VDD2.n144 9.3005
R720 VDD2.n143 VDD2.n142 9.3005
R721 VDD2.n116 VDD2.n115 9.3005
R722 VDD2.n137 VDD2.n136 9.3005
R723 VDD2.n135 VDD2.n134 9.3005
R724 VDD2.n120 VDD2.n119 9.3005
R725 VDD2.n129 VDD2.n128 9.3005
R726 VDD2.n127 VDD2.n126 9.3005
R727 VDD2.n91 VDD2.n90 9.3005
R728 VDD2.n2 VDD2.n1 9.3005
R729 VDD2.n85 VDD2.n84 9.3005
R730 VDD2.n83 VDD2.n82 9.3005
R731 VDD2.n6 VDD2.n5 9.3005
R732 VDD2.n51 VDD2.n50 9.3005
R733 VDD2.n49 VDD2.n48 9.3005
R734 VDD2.n22 VDD2.n21 9.3005
R735 VDD2.n43 VDD2.n42 9.3005
R736 VDD2.n41 VDD2.n40 9.3005
R737 VDD2.n26 VDD2.n25 9.3005
R738 VDD2.n35 VDD2.n34 9.3005
R739 VDD2.n33 VDD2.n32 9.3005
R740 VDD2.n18 VDD2.n17 9.3005
R741 VDD2.n57 VDD2.n56 9.3005
R742 VDD2.n59 VDD2.n58 9.3005
R743 VDD2.n14 VDD2.n13 9.3005
R744 VDD2.n65 VDD2.n64 9.3005
R745 VDD2.n67 VDD2.n66 9.3005
R746 VDD2.n10 VDD2.n9 9.3005
R747 VDD2.n74 VDD2.n73 9.3005
R748 VDD2.n76 VDD2.n75 9.3005
R749 VDD2.n154 VDD2.n108 8.92171
R750 VDD2.n141 VDD2.n116 8.92171
R751 VDD2.n47 VDD2.n22 8.92171
R752 VDD2.n60 VDD2.n14 8.92171
R753 VDD2.n153 VDD2.n110 8.14595
R754 VDD2.n142 VDD2.n114 8.14595
R755 VDD2.n48 VDD2.n20 8.14595
R756 VDD2.n59 VDD2.n16 8.14595
R757 VDD2.n150 VDD2.n149 7.3702
R758 VDD2.n146 VDD2.n145 7.3702
R759 VDD2.n52 VDD2.n51 7.3702
R760 VDD2.n56 VDD2.n55 7.3702
R761 VDD2.n149 VDD2.n112 6.59444
R762 VDD2.n146 VDD2.n112 6.59444
R763 VDD2.n52 VDD2.n18 6.59444
R764 VDD2.n55 VDD2.n18 6.59444
R765 VDD2.n150 VDD2.n110 5.81868
R766 VDD2.n145 VDD2.n114 5.81868
R767 VDD2.n51 VDD2.n20 5.81868
R768 VDD2.n56 VDD2.n16 5.81868
R769 VDD2.n154 VDD2.n153 5.04292
R770 VDD2.n142 VDD2.n141 5.04292
R771 VDD2.n48 VDD2.n47 5.04292
R772 VDD2.n60 VDD2.n59 5.04292
R773 VDD2.n127 VDD2.n123 4.38563
R774 VDD2.n33 VDD2.n29 4.38563
R775 VDD2.n185 VDD2.n93 4.26717
R776 VDD2.n157 VDD2.n108 4.26717
R777 VDD2.n138 VDD2.n116 4.26717
R778 VDD2.n44 VDD2.n22 4.26717
R779 VDD2.n63 VDD2.n14 4.26717
R780 VDD2.n92 VDD2.n0 4.26717
R781 VDD2.n183 VDD2.n182 3.49141
R782 VDD2.n158 VDD2.n106 3.49141
R783 VDD2.n137 VDD2.n118 3.49141
R784 VDD2.n43 VDD2.n24 3.49141
R785 VDD2.n64 VDD2.n12 3.49141
R786 VDD2.n90 VDD2.n89 3.49141
R787 VDD2.n179 VDD2.n95 2.71565
R788 VDD2.n162 VDD2.n161 2.71565
R789 VDD2.n134 VDD2.n133 2.71565
R790 VDD2.n40 VDD2.n39 2.71565
R791 VDD2.n68 VDD2.n67 2.71565
R792 VDD2.n86 VDD2.n2 2.71565
R793 VDD2.n178 VDD2.n97 1.93989
R794 VDD2.n165 VDD2.n103 1.93989
R795 VDD2.n130 VDD2.n120 1.93989
R796 VDD2.n36 VDD2.n26 1.93989
R797 VDD2.n72 VDD2.n10 1.93989
R798 VDD2.n85 VDD2.n4 1.93989
R799 VDD2.n175 VDD2.n174 1.16414
R800 VDD2.n166 VDD2.n101 1.16414
R801 VDD2.n129 VDD2.n122 1.16414
R802 VDD2.n35 VDD2.n28 1.16414
R803 VDD2.n73 VDD2.n8 1.16414
R804 VDD2.n82 VDD2.n81 1.16414
R805 VDD2.n171 VDD2.n99 0.388379
R806 VDD2.n170 VDD2.n169 0.388379
R807 VDD2.n126 VDD2.n125 0.388379
R808 VDD2.n32 VDD2.n31 0.388379
R809 VDD2.n77 VDD2.n76 0.388379
R810 VDD2.n78 VDD2.n6 0.388379
R811 VDD2 VDD2.n186 0.237569
R812 VDD2.n184 VDD2.n94 0.155672
R813 VDD2.n177 VDD2.n94 0.155672
R814 VDD2.n177 VDD2.n176 0.155672
R815 VDD2.n176 VDD2.n98 0.155672
R816 VDD2.n168 VDD2.n98 0.155672
R817 VDD2.n168 VDD2.n167 0.155672
R818 VDD2.n167 VDD2.n102 0.155672
R819 VDD2.n160 VDD2.n102 0.155672
R820 VDD2.n160 VDD2.n159 0.155672
R821 VDD2.n159 VDD2.n107 0.155672
R822 VDD2.n152 VDD2.n107 0.155672
R823 VDD2.n152 VDD2.n151 0.155672
R824 VDD2.n151 VDD2.n111 0.155672
R825 VDD2.n144 VDD2.n111 0.155672
R826 VDD2.n144 VDD2.n143 0.155672
R827 VDD2.n143 VDD2.n115 0.155672
R828 VDD2.n136 VDD2.n115 0.155672
R829 VDD2.n136 VDD2.n135 0.155672
R830 VDD2.n135 VDD2.n119 0.155672
R831 VDD2.n128 VDD2.n119 0.155672
R832 VDD2.n128 VDD2.n127 0.155672
R833 VDD2.n34 VDD2.n33 0.155672
R834 VDD2.n34 VDD2.n25 0.155672
R835 VDD2.n41 VDD2.n25 0.155672
R836 VDD2.n42 VDD2.n41 0.155672
R837 VDD2.n42 VDD2.n21 0.155672
R838 VDD2.n49 VDD2.n21 0.155672
R839 VDD2.n50 VDD2.n49 0.155672
R840 VDD2.n50 VDD2.n17 0.155672
R841 VDD2.n57 VDD2.n17 0.155672
R842 VDD2.n58 VDD2.n57 0.155672
R843 VDD2.n58 VDD2.n13 0.155672
R844 VDD2.n65 VDD2.n13 0.155672
R845 VDD2.n66 VDD2.n65 0.155672
R846 VDD2.n66 VDD2.n9 0.155672
R847 VDD2.n74 VDD2.n9 0.155672
R848 VDD2.n75 VDD2.n74 0.155672
R849 VDD2.n75 VDD2.n5 0.155672
R850 VDD2.n83 VDD2.n5 0.155672
R851 VDD2.n84 VDD2.n83 0.155672
R852 VDD2.n84 VDD2.n1 0.155672
R853 VDD2.n91 VDD2.n1 0.155672
R854 B.n421 B.t9 1011.35
R855 B.n419 B.t13 1011.35
R856 B.n91 B.t2 1011.35
R857 B.n89 B.t6 1011.35
R858 B.n723 B.n722 585
R859 B.n724 B.n723 585
R860 B.n333 B.n88 585
R861 B.n332 B.n331 585
R862 B.n330 B.n329 585
R863 B.n328 B.n327 585
R864 B.n326 B.n325 585
R865 B.n324 B.n323 585
R866 B.n322 B.n321 585
R867 B.n320 B.n319 585
R868 B.n318 B.n317 585
R869 B.n316 B.n315 585
R870 B.n314 B.n313 585
R871 B.n312 B.n311 585
R872 B.n310 B.n309 585
R873 B.n308 B.n307 585
R874 B.n306 B.n305 585
R875 B.n304 B.n303 585
R876 B.n302 B.n301 585
R877 B.n300 B.n299 585
R878 B.n298 B.n297 585
R879 B.n296 B.n295 585
R880 B.n294 B.n293 585
R881 B.n292 B.n291 585
R882 B.n290 B.n289 585
R883 B.n288 B.n287 585
R884 B.n286 B.n285 585
R885 B.n284 B.n283 585
R886 B.n282 B.n281 585
R887 B.n280 B.n279 585
R888 B.n278 B.n277 585
R889 B.n276 B.n275 585
R890 B.n274 B.n273 585
R891 B.n272 B.n271 585
R892 B.n270 B.n269 585
R893 B.n268 B.n267 585
R894 B.n266 B.n265 585
R895 B.n264 B.n263 585
R896 B.n262 B.n261 585
R897 B.n260 B.n259 585
R898 B.n258 B.n257 585
R899 B.n256 B.n255 585
R900 B.n254 B.n253 585
R901 B.n252 B.n251 585
R902 B.n250 B.n249 585
R903 B.n248 B.n247 585
R904 B.n246 B.n245 585
R905 B.n244 B.n243 585
R906 B.n242 B.n241 585
R907 B.n240 B.n239 585
R908 B.n238 B.n237 585
R909 B.n236 B.n235 585
R910 B.n234 B.n233 585
R911 B.n232 B.n231 585
R912 B.n230 B.n229 585
R913 B.n228 B.n227 585
R914 B.n226 B.n225 585
R915 B.n223 B.n222 585
R916 B.n221 B.n220 585
R917 B.n219 B.n218 585
R918 B.n217 B.n216 585
R919 B.n215 B.n214 585
R920 B.n213 B.n212 585
R921 B.n211 B.n210 585
R922 B.n209 B.n208 585
R923 B.n207 B.n206 585
R924 B.n205 B.n204 585
R925 B.n203 B.n202 585
R926 B.n201 B.n200 585
R927 B.n199 B.n198 585
R928 B.n197 B.n196 585
R929 B.n195 B.n194 585
R930 B.n193 B.n192 585
R931 B.n191 B.n190 585
R932 B.n189 B.n188 585
R933 B.n187 B.n186 585
R934 B.n185 B.n184 585
R935 B.n183 B.n182 585
R936 B.n181 B.n180 585
R937 B.n179 B.n178 585
R938 B.n177 B.n176 585
R939 B.n175 B.n174 585
R940 B.n173 B.n172 585
R941 B.n171 B.n170 585
R942 B.n169 B.n168 585
R943 B.n167 B.n166 585
R944 B.n165 B.n164 585
R945 B.n163 B.n162 585
R946 B.n161 B.n160 585
R947 B.n159 B.n158 585
R948 B.n157 B.n156 585
R949 B.n155 B.n154 585
R950 B.n153 B.n152 585
R951 B.n151 B.n150 585
R952 B.n149 B.n148 585
R953 B.n147 B.n146 585
R954 B.n145 B.n144 585
R955 B.n143 B.n142 585
R956 B.n141 B.n140 585
R957 B.n139 B.n138 585
R958 B.n137 B.n136 585
R959 B.n135 B.n134 585
R960 B.n133 B.n132 585
R961 B.n131 B.n130 585
R962 B.n129 B.n128 585
R963 B.n127 B.n126 585
R964 B.n125 B.n124 585
R965 B.n123 B.n122 585
R966 B.n121 B.n120 585
R967 B.n119 B.n118 585
R968 B.n117 B.n116 585
R969 B.n115 B.n114 585
R970 B.n113 B.n112 585
R971 B.n111 B.n110 585
R972 B.n109 B.n108 585
R973 B.n107 B.n106 585
R974 B.n105 B.n104 585
R975 B.n103 B.n102 585
R976 B.n101 B.n100 585
R977 B.n99 B.n98 585
R978 B.n97 B.n96 585
R979 B.n95 B.n94 585
R980 B.n721 B.n27 585
R981 B.n725 B.n27 585
R982 B.n720 B.n26 585
R983 B.n726 B.n26 585
R984 B.n719 B.n718 585
R985 B.n718 B.n22 585
R986 B.n717 B.n21 585
R987 B.n732 B.n21 585
R988 B.n716 B.n20 585
R989 B.n733 B.n20 585
R990 B.n715 B.n19 585
R991 B.n734 B.n19 585
R992 B.n714 B.n713 585
R993 B.n713 B.n15 585
R994 B.n712 B.n14 585
R995 B.n740 B.n14 585
R996 B.n711 B.n13 585
R997 B.n741 B.n13 585
R998 B.n710 B.n12 585
R999 B.n742 B.n12 585
R1000 B.n709 B.n708 585
R1001 B.n708 B.n11 585
R1002 B.n707 B.n7 585
R1003 B.n748 B.n7 585
R1004 B.n706 B.n6 585
R1005 B.n749 B.n6 585
R1006 B.n705 B.n5 585
R1007 B.n750 B.n5 585
R1008 B.n704 B.n703 585
R1009 B.n703 B.n4 585
R1010 B.n702 B.n334 585
R1011 B.n702 B.n701 585
R1012 B.n691 B.n335 585
R1013 B.n694 B.n335 585
R1014 B.n693 B.n692 585
R1015 B.n695 B.n693 585
R1016 B.n690 B.n340 585
R1017 B.n340 B.n339 585
R1018 B.n689 B.n688 585
R1019 B.n688 B.n687 585
R1020 B.n342 B.n341 585
R1021 B.n343 B.n342 585
R1022 B.n680 B.n679 585
R1023 B.n681 B.n680 585
R1024 B.n678 B.n347 585
R1025 B.n351 B.n347 585
R1026 B.n677 B.n676 585
R1027 B.n676 B.n675 585
R1028 B.n349 B.n348 585
R1029 B.n350 B.n349 585
R1030 B.n668 B.n667 585
R1031 B.n669 B.n668 585
R1032 B.n666 B.n356 585
R1033 B.n356 B.n355 585
R1034 B.n660 B.n659 585
R1035 B.n658 B.n418 585
R1036 B.n657 B.n417 585
R1037 B.n662 B.n417 585
R1038 B.n656 B.n655 585
R1039 B.n654 B.n653 585
R1040 B.n652 B.n651 585
R1041 B.n650 B.n649 585
R1042 B.n648 B.n647 585
R1043 B.n646 B.n645 585
R1044 B.n644 B.n643 585
R1045 B.n642 B.n641 585
R1046 B.n640 B.n639 585
R1047 B.n638 B.n637 585
R1048 B.n636 B.n635 585
R1049 B.n634 B.n633 585
R1050 B.n632 B.n631 585
R1051 B.n630 B.n629 585
R1052 B.n628 B.n627 585
R1053 B.n626 B.n625 585
R1054 B.n624 B.n623 585
R1055 B.n622 B.n621 585
R1056 B.n620 B.n619 585
R1057 B.n618 B.n617 585
R1058 B.n616 B.n615 585
R1059 B.n614 B.n613 585
R1060 B.n612 B.n611 585
R1061 B.n610 B.n609 585
R1062 B.n608 B.n607 585
R1063 B.n606 B.n605 585
R1064 B.n604 B.n603 585
R1065 B.n602 B.n601 585
R1066 B.n600 B.n599 585
R1067 B.n598 B.n597 585
R1068 B.n596 B.n595 585
R1069 B.n594 B.n593 585
R1070 B.n592 B.n591 585
R1071 B.n590 B.n589 585
R1072 B.n588 B.n587 585
R1073 B.n586 B.n585 585
R1074 B.n584 B.n583 585
R1075 B.n582 B.n581 585
R1076 B.n580 B.n579 585
R1077 B.n578 B.n577 585
R1078 B.n576 B.n575 585
R1079 B.n574 B.n573 585
R1080 B.n572 B.n571 585
R1081 B.n570 B.n569 585
R1082 B.n568 B.n567 585
R1083 B.n566 B.n565 585
R1084 B.n564 B.n563 585
R1085 B.n562 B.n561 585
R1086 B.n560 B.n559 585
R1087 B.n558 B.n557 585
R1088 B.n556 B.n555 585
R1089 B.n554 B.n553 585
R1090 B.n552 B.n551 585
R1091 B.n549 B.n548 585
R1092 B.n547 B.n546 585
R1093 B.n545 B.n544 585
R1094 B.n543 B.n542 585
R1095 B.n541 B.n540 585
R1096 B.n539 B.n538 585
R1097 B.n537 B.n536 585
R1098 B.n535 B.n534 585
R1099 B.n533 B.n532 585
R1100 B.n531 B.n530 585
R1101 B.n529 B.n528 585
R1102 B.n527 B.n526 585
R1103 B.n525 B.n524 585
R1104 B.n523 B.n522 585
R1105 B.n521 B.n520 585
R1106 B.n519 B.n518 585
R1107 B.n517 B.n516 585
R1108 B.n515 B.n514 585
R1109 B.n513 B.n512 585
R1110 B.n511 B.n510 585
R1111 B.n509 B.n508 585
R1112 B.n507 B.n506 585
R1113 B.n505 B.n504 585
R1114 B.n503 B.n502 585
R1115 B.n501 B.n500 585
R1116 B.n499 B.n498 585
R1117 B.n497 B.n496 585
R1118 B.n495 B.n494 585
R1119 B.n493 B.n492 585
R1120 B.n491 B.n490 585
R1121 B.n489 B.n488 585
R1122 B.n487 B.n486 585
R1123 B.n485 B.n484 585
R1124 B.n483 B.n482 585
R1125 B.n481 B.n480 585
R1126 B.n479 B.n478 585
R1127 B.n477 B.n476 585
R1128 B.n475 B.n474 585
R1129 B.n473 B.n472 585
R1130 B.n471 B.n470 585
R1131 B.n469 B.n468 585
R1132 B.n467 B.n466 585
R1133 B.n465 B.n464 585
R1134 B.n463 B.n462 585
R1135 B.n461 B.n460 585
R1136 B.n459 B.n458 585
R1137 B.n457 B.n456 585
R1138 B.n455 B.n454 585
R1139 B.n453 B.n452 585
R1140 B.n451 B.n450 585
R1141 B.n449 B.n448 585
R1142 B.n447 B.n446 585
R1143 B.n445 B.n444 585
R1144 B.n443 B.n442 585
R1145 B.n441 B.n440 585
R1146 B.n439 B.n438 585
R1147 B.n437 B.n436 585
R1148 B.n435 B.n434 585
R1149 B.n433 B.n432 585
R1150 B.n431 B.n430 585
R1151 B.n429 B.n428 585
R1152 B.n427 B.n426 585
R1153 B.n425 B.n424 585
R1154 B.n358 B.n357 585
R1155 B.n665 B.n664 585
R1156 B.n354 B.n353 585
R1157 B.n355 B.n354 585
R1158 B.n671 B.n670 585
R1159 B.n670 B.n669 585
R1160 B.n672 B.n352 585
R1161 B.n352 B.n350 585
R1162 B.n674 B.n673 585
R1163 B.n675 B.n674 585
R1164 B.n346 B.n345 585
R1165 B.n351 B.n346 585
R1166 B.n683 B.n682 585
R1167 B.n682 B.n681 585
R1168 B.n684 B.n344 585
R1169 B.n344 B.n343 585
R1170 B.n686 B.n685 585
R1171 B.n687 B.n686 585
R1172 B.n338 B.n337 585
R1173 B.n339 B.n338 585
R1174 B.n697 B.n696 585
R1175 B.n696 B.n695 585
R1176 B.n698 B.n336 585
R1177 B.n694 B.n336 585
R1178 B.n700 B.n699 585
R1179 B.n701 B.n700 585
R1180 B.n2 B.n0 585
R1181 B.n4 B.n2 585
R1182 B.n3 B.n1 585
R1183 B.n749 B.n3 585
R1184 B.n747 B.n746 585
R1185 B.n748 B.n747 585
R1186 B.n745 B.n8 585
R1187 B.n11 B.n8 585
R1188 B.n744 B.n743 585
R1189 B.n743 B.n742 585
R1190 B.n10 B.n9 585
R1191 B.n741 B.n10 585
R1192 B.n739 B.n738 585
R1193 B.n740 B.n739 585
R1194 B.n737 B.n16 585
R1195 B.n16 B.n15 585
R1196 B.n736 B.n735 585
R1197 B.n735 B.n734 585
R1198 B.n18 B.n17 585
R1199 B.n733 B.n18 585
R1200 B.n731 B.n730 585
R1201 B.n732 B.n731 585
R1202 B.n729 B.n23 585
R1203 B.n23 B.n22 585
R1204 B.n728 B.n727 585
R1205 B.n727 B.n726 585
R1206 B.n25 B.n24 585
R1207 B.n725 B.n25 585
R1208 B.n752 B.n751 585
R1209 B.n751 B.n750 585
R1210 B.n660 B.n354 463.671
R1211 B.n94 B.n25 463.671
R1212 B.n664 B.n356 463.671
R1213 B.n723 B.n27 463.671
R1214 B.n421 B.t12 378.928
R1215 B.n89 B.t7 378.928
R1216 B.n419 B.t15 378.928
R1217 B.n91 B.t4 378.928
R1218 B.n422 B.t11 362.832
R1219 B.n90 B.t8 362.832
R1220 B.n420 B.t14 362.832
R1221 B.n92 B.t5 362.832
R1222 B.n724 B.n87 256.663
R1223 B.n724 B.n86 256.663
R1224 B.n724 B.n85 256.663
R1225 B.n724 B.n84 256.663
R1226 B.n724 B.n83 256.663
R1227 B.n724 B.n82 256.663
R1228 B.n724 B.n81 256.663
R1229 B.n724 B.n80 256.663
R1230 B.n724 B.n79 256.663
R1231 B.n724 B.n78 256.663
R1232 B.n724 B.n77 256.663
R1233 B.n724 B.n76 256.663
R1234 B.n724 B.n75 256.663
R1235 B.n724 B.n74 256.663
R1236 B.n724 B.n73 256.663
R1237 B.n724 B.n72 256.663
R1238 B.n724 B.n71 256.663
R1239 B.n724 B.n70 256.663
R1240 B.n724 B.n69 256.663
R1241 B.n724 B.n68 256.663
R1242 B.n724 B.n67 256.663
R1243 B.n724 B.n66 256.663
R1244 B.n724 B.n65 256.663
R1245 B.n724 B.n64 256.663
R1246 B.n724 B.n63 256.663
R1247 B.n724 B.n62 256.663
R1248 B.n724 B.n61 256.663
R1249 B.n724 B.n60 256.663
R1250 B.n724 B.n59 256.663
R1251 B.n724 B.n58 256.663
R1252 B.n724 B.n57 256.663
R1253 B.n724 B.n56 256.663
R1254 B.n724 B.n55 256.663
R1255 B.n724 B.n54 256.663
R1256 B.n724 B.n53 256.663
R1257 B.n724 B.n52 256.663
R1258 B.n724 B.n51 256.663
R1259 B.n724 B.n50 256.663
R1260 B.n724 B.n49 256.663
R1261 B.n724 B.n48 256.663
R1262 B.n724 B.n47 256.663
R1263 B.n724 B.n46 256.663
R1264 B.n724 B.n45 256.663
R1265 B.n724 B.n44 256.663
R1266 B.n724 B.n43 256.663
R1267 B.n724 B.n42 256.663
R1268 B.n724 B.n41 256.663
R1269 B.n724 B.n40 256.663
R1270 B.n724 B.n39 256.663
R1271 B.n724 B.n38 256.663
R1272 B.n724 B.n37 256.663
R1273 B.n724 B.n36 256.663
R1274 B.n724 B.n35 256.663
R1275 B.n724 B.n34 256.663
R1276 B.n724 B.n33 256.663
R1277 B.n724 B.n32 256.663
R1278 B.n724 B.n31 256.663
R1279 B.n724 B.n30 256.663
R1280 B.n724 B.n29 256.663
R1281 B.n724 B.n28 256.663
R1282 B.n662 B.n661 256.663
R1283 B.n662 B.n359 256.663
R1284 B.n662 B.n360 256.663
R1285 B.n662 B.n361 256.663
R1286 B.n662 B.n362 256.663
R1287 B.n662 B.n363 256.663
R1288 B.n662 B.n364 256.663
R1289 B.n662 B.n365 256.663
R1290 B.n662 B.n366 256.663
R1291 B.n662 B.n367 256.663
R1292 B.n662 B.n368 256.663
R1293 B.n662 B.n369 256.663
R1294 B.n662 B.n370 256.663
R1295 B.n662 B.n371 256.663
R1296 B.n662 B.n372 256.663
R1297 B.n662 B.n373 256.663
R1298 B.n662 B.n374 256.663
R1299 B.n662 B.n375 256.663
R1300 B.n662 B.n376 256.663
R1301 B.n662 B.n377 256.663
R1302 B.n662 B.n378 256.663
R1303 B.n662 B.n379 256.663
R1304 B.n662 B.n380 256.663
R1305 B.n662 B.n381 256.663
R1306 B.n662 B.n382 256.663
R1307 B.n662 B.n383 256.663
R1308 B.n662 B.n384 256.663
R1309 B.n662 B.n385 256.663
R1310 B.n662 B.n386 256.663
R1311 B.n662 B.n387 256.663
R1312 B.n662 B.n388 256.663
R1313 B.n662 B.n389 256.663
R1314 B.n662 B.n390 256.663
R1315 B.n662 B.n391 256.663
R1316 B.n662 B.n392 256.663
R1317 B.n662 B.n393 256.663
R1318 B.n662 B.n394 256.663
R1319 B.n662 B.n395 256.663
R1320 B.n662 B.n396 256.663
R1321 B.n662 B.n397 256.663
R1322 B.n662 B.n398 256.663
R1323 B.n662 B.n399 256.663
R1324 B.n662 B.n400 256.663
R1325 B.n662 B.n401 256.663
R1326 B.n662 B.n402 256.663
R1327 B.n662 B.n403 256.663
R1328 B.n662 B.n404 256.663
R1329 B.n662 B.n405 256.663
R1330 B.n662 B.n406 256.663
R1331 B.n662 B.n407 256.663
R1332 B.n662 B.n408 256.663
R1333 B.n662 B.n409 256.663
R1334 B.n662 B.n410 256.663
R1335 B.n662 B.n411 256.663
R1336 B.n662 B.n412 256.663
R1337 B.n662 B.n413 256.663
R1338 B.n662 B.n414 256.663
R1339 B.n662 B.n415 256.663
R1340 B.n662 B.n416 256.663
R1341 B.n663 B.n662 256.663
R1342 B.n670 B.n354 163.367
R1343 B.n670 B.n352 163.367
R1344 B.n674 B.n352 163.367
R1345 B.n674 B.n346 163.367
R1346 B.n682 B.n346 163.367
R1347 B.n682 B.n344 163.367
R1348 B.n686 B.n344 163.367
R1349 B.n686 B.n338 163.367
R1350 B.n696 B.n338 163.367
R1351 B.n696 B.n336 163.367
R1352 B.n700 B.n336 163.367
R1353 B.n700 B.n2 163.367
R1354 B.n751 B.n2 163.367
R1355 B.n751 B.n3 163.367
R1356 B.n747 B.n3 163.367
R1357 B.n747 B.n8 163.367
R1358 B.n743 B.n8 163.367
R1359 B.n743 B.n10 163.367
R1360 B.n739 B.n10 163.367
R1361 B.n739 B.n16 163.367
R1362 B.n735 B.n16 163.367
R1363 B.n735 B.n18 163.367
R1364 B.n731 B.n18 163.367
R1365 B.n731 B.n23 163.367
R1366 B.n727 B.n23 163.367
R1367 B.n727 B.n25 163.367
R1368 B.n418 B.n417 163.367
R1369 B.n655 B.n417 163.367
R1370 B.n653 B.n652 163.367
R1371 B.n649 B.n648 163.367
R1372 B.n645 B.n644 163.367
R1373 B.n641 B.n640 163.367
R1374 B.n637 B.n636 163.367
R1375 B.n633 B.n632 163.367
R1376 B.n629 B.n628 163.367
R1377 B.n625 B.n624 163.367
R1378 B.n621 B.n620 163.367
R1379 B.n617 B.n616 163.367
R1380 B.n613 B.n612 163.367
R1381 B.n609 B.n608 163.367
R1382 B.n605 B.n604 163.367
R1383 B.n601 B.n600 163.367
R1384 B.n597 B.n596 163.367
R1385 B.n593 B.n592 163.367
R1386 B.n589 B.n588 163.367
R1387 B.n585 B.n584 163.367
R1388 B.n581 B.n580 163.367
R1389 B.n577 B.n576 163.367
R1390 B.n573 B.n572 163.367
R1391 B.n569 B.n568 163.367
R1392 B.n565 B.n564 163.367
R1393 B.n561 B.n560 163.367
R1394 B.n557 B.n556 163.367
R1395 B.n553 B.n552 163.367
R1396 B.n548 B.n547 163.367
R1397 B.n544 B.n543 163.367
R1398 B.n540 B.n539 163.367
R1399 B.n536 B.n535 163.367
R1400 B.n532 B.n531 163.367
R1401 B.n528 B.n527 163.367
R1402 B.n524 B.n523 163.367
R1403 B.n520 B.n519 163.367
R1404 B.n516 B.n515 163.367
R1405 B.n512 B.n511 163.367
R1406 B.n508 B.n507 163.367
R1407 B.n504 B.n503 163.367
R1408 B.n500 B.n499 163.367
R1409 B.n496 B.n495 163.367
R1410 B.n492 B.n491 163.367
R1411 B.n488 B.n487 163.367
R1412 B.n484 B.n483 163.367
R1413 B.n480 B.n479 163.367
R1414 B.n476 B.n475 163.367
R1415 B.n472 B.n471 163.367
R1416 B.n468 B.n467 163.367
R1417 B.n464 B.n463 163.367
R1418 B.n460 B.n459 163.367
R1419 B.n456 B.n455 163.367
R1420 B.n452 B.n451 163.367
R1421 B.n448 B.n447 163.367
R1422 B.n444 B.n443 163.367
R1423 B.n440 B.n439 163.367
R1424 B.n436 B.n435 163.367
R1425 B.n432 B.n431 163.367
R1426 B.n428 B.n427 163.367
R1427 B.n424 B.n358 163.367
R1428 B.n668 B.n356 163.367
R1429 B.n668 B.n349 163.367
R1430 B.n676 B.n349 163.367
R1431 B.n676 B.n347 163.367
R1432 B.n680 B.n347 163.367
R1433 B.n680 B.n342 163.367
R1434 B.n688 B.n342 163.367
R1435 B.n688 B.n340 163.367
R1436 B.n693 B.n340 163.367
R1437 B.n693 B.n335 163.367
R1438 B.n702 B.n335 163.367
R1439 B.n703 B.n702 163.367
R1440 B.n703 B.n5 163.367
R1441 B.n6 B.n5 163.367
R1442 B.n7 B.n6 163.367
R1443 B.n708 B.n7 163.367
R1444 B.n708 B.n12 163.367
R1445 B.n13 B.n12 163.367
R1446 B.n14 B.n13 163.367
R1447 B.n713 B.n14 163.367
R1448 B.n713 B.n19 163.367
R1449 B.n20 B.n19 163.367
R1450 B.n21 B.n20 163.367
R1451 B.n718 B.n21 163.367
R1452 B.n718 B.n26 163.367
R1453 B.n27 B.n26 163.367
R1454 B.n98 B.n97 163.367
R1455 B.n102 B.n101 163.367
R1456 B.n106 B.n105 163.367
R1457 B.n110 B.n109 163.367
R1458 B.n114 B.n113 163.367
R1459 B.n118 B.n117 163.367
R1460 B.n122 B.n121 163.367
R1461 B.n126 B.n125 163.367
R1462 B.n130 B.n129 163.367
R1463 B.n134 B.n133 163.367
R1464 B.n138 B.n137 163.367
R1465 B.n142 B.n141 163.367
R1466 B.n146 B.n145 163.367
R1467 B.n150 B.n149 163.367
R1468 B.n154 B.n153 163.367
R1469 B.n158 B.n157 163.367
R1470 B.n162 B.n161 163.367
R1471 B.n166 B.n165 163.367
R1472 B.n170 B.n169 163.367
R1473 B.n174 B.n173 163.367
R1474 B.n178 B.n177 163.367
R1475 B.n182 B.n181 163.367
R1476 B.n186 B.n185 163.367
R1477 B.n190 B.n189 163.367
R1478 B.n194 B.n193 163.367
R1479 B.n198 B.n197 163.367
R1480 B.n202 B.n201 163.367
R1481 B.n206 B.n205 163.367
R1482 B.n210 B.n209 163.367
R1483 B.n214 B.n213 163.367
R1484 B.n218 B.n217 163.367
R1485 B.n222 B.n221 163.367
R1486 B.n227 B.n226 163.367
R1487 B.n231 B.n230 163.367
R1488 B.n235 B.n234 163.367
R1489 B.n239 B.n238 163.367
R1490 B.n243 B.n242 163.367
R1491 B.n247 B.n246 163.367
R1492 B.n251 B.n250 163.367
R1493 B.n255 B.n254 163.367
R1494 B.n259 B.n258 163.367
R1495 B.n263 B.n262 163.367
R1496 B.n267 B.n266 163.367
R1497 B.n271 B.n270 163.367
R1498 B.n275 B.n274 163.367
R1499 B.n279 B.n278 163.367
R1500 B.n283 B.n282 163.367
R1501 B.n287 B.n286 163.367
R1502 B.n291 B.n290 163.367
R1503 B.n295 B.n294 163.367
R1504 B.n299 B.n298 163.367
R1505 B.n303 B.n302 163.367
R1506 B.n307 B.n306 163.367
R1507 B.n311 B.n310 163.367
R1508 B.n315 B.n314 163.367
R1509 B.n319 B.n318 163.367
R1510 B.n323 B.n322 163.367
R1511 B.n327 B.n326 163.367
R1512 B.n331 B.n330 163.367
R1513 B.n723 B.n88 163.367
R1514 B.n661 B.n660 71.676
R1515 B.n655 B.n359 71.676
R1516 B.n652 B.n360 71.676
R1517 B.n648 B.n361 71.676
R1518 B.n644 B.n362 71.676
R1519 B.n640 B.n363 71.676
R1520 B.n636 B.n364 71.676
R1521 B.n632 B.n365 71.676
R1522 B.n628 B.n366 71.676
R1523 B.n624 B.n367 71.676
R1524 B.n620 B.n368 71.676
R1525 B.n616 B.n369 71.676
R1526 B.n612 B.n370 71.676
R1527 B.n608 B.n371 71.676
R1528 B.n604 B.n372 71.676
R1529 B.n600 B.n373 71.676
R1530 B.n596 B.n374 71.676
R1531 B.n592 B.n375 71.676
R1532 B.n588 B.n376 71.676
R1533 B.n584 B.n377 71.676
R1534 B.n580 B.n378 71.676
R1535 B.n576 B.n379 71.676
R1536 B.n572 B.n380 71.676
R1537 B.n568 B.n381 71.676
R1538 B.n564 B.n382 71.676
R1539 B.n560 B.n383 71.676
R1540 B.n556 B.n384 71.676
R1541 B.n552 B.n385 71.676
R1542 B.n547 B.n386 71.676
R1543 B.n543 B.n387 71.676
R1544 B.n539 B.n388 71.676
R1545 B.n535 B.n389 71.676
R1546 B.n531 B.n390 71.676
R1547 B.n527 B.n391 71.676
R1548 B.n523 B.n392 71.676
R1549 B.n519 B.n393 71.676
R1550 B.n515 B.n394 71.676
R1551 B.n511 B.n395 71.676
R1552 B.n507 B.n396 71.676
R1553 B.n503 B.n397 71.676
R1554 B.n499 B.n398 71.676
R1555 B.n495 B.n399 71.676
R1556 B.n491 B.n400 71.676
R1557 B.n487 B.n401 71.676
R1558 B.n483 B.n402 71.676
R1559 B.n479 B.n403 71.676
R1560 B.n475 B.n404 71.676
R1561 B.n471 B.n405 71.676
R1562 B.n467 B.n406 71.676
R1563 B.n463 B.n407 71.676
R1564 B.n459 B.n408 71.676
R1565 B.n455 B.n409 71.676
R1566 B.n451 B.n410 71.676
R1567 B.n447 B.n411 71.676
R1568 B.n443 B.n412 71.676
R1569 B.n439 B.n413 71.676
R1570 B.n435 B.n414 71.676
R1571 B.n431 B.n415 71.676
R1572 B.n427 B.n416 71.676
R1573 B.n663 B.n358 71.676
R1574 B.n94 B.n28 71.676
R1575 B.n98 B.n29 71.676
R1576 B.n102 B.n30 71.676
R1577 B.n106 B.n31 71.676
R1578 B.n110 B.n32 71.676
R1579 B.n114 B.n33 71.676
R1580 B.n118 B.n34 71.676
R1581 B.n122 B.n35 71.676
R1582 B.n126 B.n36 71.676
R1583 B.n130 B.n37 71.676
R1584 B.n134 B.n38 71.676
R1585 B.n138 B.n39 71.676
R1586 B.n142 B.n40 71.676
R1587 B.n146 B.n41 71.676
R1588 B.n150 B.n42 71.676
R1589 B.n154 B.n43 71.676
R1590 B.n158 B.n44 71.676
R1591 B.n162 B.n45 71.676
R1592 B.n166 B.n46 71.676
R1593 B.n170 B.n47 71.676
R1594 B.n174 B.n48 71.676
R1595 B.n178 B.n49 71.676
R1596 B.n182 B.n50 71.676
R1597 B.n186 B.n51 71.676
R1598 B.n190 B.n52 71.676
R1599 B.n194 B.n53 71.676
R1600 B.n198 B.n54 71.676
R1601 B.n202 B.n55 71.676
R1602 B.n206 B.n56 71.676
R1603 B.n210 B.n57 71.676
R1604 B.n214 B.n58 71.676
R1605 B.n218 B.n59 71.676
R1606 B.n222 B.n60 71.676
R1607 B.n227 B.n61 71.676
R1608 B.n231 B.n62 71.676
R1609 B.n235 B.n63 71.676
R1610 B.n239 B.n64 71.676
R1611 B.n243 B.n65 71.676
R1612 B.n247 B.n66 71.676
R1613 B.n251 B.n67 71.676
R1614 B.n255 B.n68 71.676
R1615 B.n259 B.n69 71.676
R1616 B.n263 B.n70 71.676
R1617 B.n267 B.n71 71.676
R1618 B.n271 B.n72 71.676
R1619 B.n275 B.n73 71.676
R1620 B.n279 B.n74 71.676
R1621 B.n283 B.n75 71.676
R1622 B.n287 B.n76 71.676
R1623 B.n291 B.n77 71.676
R1624 B.n295 B.n78 71.676
R1625 B.n299 B.n79 71.676
R1626 B.n303 B.n80 71.676
R1627 B.n307 B.n81 71.676
R1628 B.n311 B.n82 71.676
R1629 B.n315 B.n83 71.676
R1630 B.n319 B.n84 71.676
R1631 B.n323 B.n85 71.676
R1632 B.n327 B.n86 71.676
R1633 B.n331 B.n87 71.676
R1634 B.n88 B.n87 71.676
R1635 B.n330 B.n86 71.676
R1636 B.n326 B.n85 71.676
R1637 B.n322 B.n84 71.676
R1638 B.n318 B.n83 71.676
R1639 B.n314 B.n82 71.676
R1640 B.n310 B.n81 71.676
R1641 B.n306 B.n80 71.676
R1642 B.n302 B.n79 71.676
R1643 B.n298 B.n78 71.676
R1644 B.n294 B.n77 71.676
R1645 B.n290 B.n76 71.676
R1646 B.n286 B.n75 71.676
R1647 B.n282 B.n74 71.676
R1648 B.n278 B.n73 71.676
R1649 B.n274 B.n72 71.676
R1650 B.n270 B.n71 71.676
R1651 B.n266 B.n70 71.676
R1652 B.n262 B.n69 71.676
R1653 B.n258 B.n68 71.676
R1654 B.n254 B.n67 71.676
R1655 B.n250 B.n66 71.676
R1656 B.n246 B.n65 71.676
R1657 B.n242 B.n64 71.676
R1658 B.n238 B.n63 71.676
R1659 B.n234 B.n62 71.676
R1660 B.n230 B.n61 71.676
R1661 B.n226 B.n60 71.676
R1662 B.n221 B.n59 71.676
R1663 B.n217 B.n58 71.676
R1664 B.n213 B.n57 71.676
R1665 B.n209 B.n56 71.676
R1666 B.n205 B.n55 71.676
R1667 B.n201 B.n54 71.676
R1668 B.n197 B.n53 71.676
R1669 B.n193 B.n52 71.676
R1670 B.n189 B.n51 71.676
R1671 B.n185 B.n50 71.676
R1672 B.n181 B.n49 71.676
R1673 B.n177 B.n48 71.676
R1674 B.n173 B.n47 71.676
R1675 B.n169 B.n46 71.676
R1676 B.n165 B.n45 71.676
R1677 B.n161 B.n44 71.676
R1678 B.n157 B.n43 71.676
R1679 B.n153 B.n42 71.676
R1680 B.n149 B.n41 71.676
R1681 B.n145 B.n40 71.676
R1682 B.n141 B.n39 71.676
R1683 B.n137 B.n38 71.676
R1684 B.n133 B.n37 71.676
R1685 B.n129 B.n36 71.676
R1686 B.n125 B.n35 71.676
R1687 B.n121 B.n34 71.676
R1688 B.n117 B.n33 71.676
R1689 B.n113 B.n32 71.676
R1690 B.n109 B.n31 71.676
R1691 B.n105 B.n30 71.676
R1692 B.n101 B.n29 71.676
R1693 B.n97 B.n28 71.676
R1694 B.n661 B.n418 71.676
R1695 B.n653 B.n359 71.676
R1696 B.n649 B.n360 71.676
R1697 B.n645 B.n361 71.676
R1698 B.n641 B.n362 71.676
R1699 B.n637 B.n363 71.676
R1700 B.n633 B.n364 71.676
R1701 B.n629 B.n365 71.676
R1702 B.n625 B.n366 71.676
R1703 B.n621 B.n367 71.676
R1704 B.n617 B.n368 71.676
R1705 B.n613 B.n369 71.676
R1706 B.n609 B.n370 71.676
R1707 B.n605 B.n371 71.676
R1708 B.n601 B.n372 71.676
R1709 B.n597 B.n373 71.676
R1710 B.n593 B.n374 71.676
R1711 B.n589 B.n375 71.676
R1712 B.n585 B.n376 71.676
R1713 B.n581 B.n377 71.676
R1714 B.n577 B.n378 71.676
R1715 B.n573 B.n379 71.676
R1716 B.n569 B.n380 71.676
R1717 B.n565 B.n381 71.676
R1718 B.n561 B.n382 71.676
R1719 B.n557 B.n383 71.676
R1720 B.n553 B.n384 71.676
R1721 B.n548 B.n385 71.676
R1722 B.n544 B.n386 71.676
R1723 B.n540 B.n387 71.676
R1724 B.n536 B.n388 71.676
R1725 B.n532 B.n389 71.676
R1726 B.n528 B.n390 71.676
R1727 B.n524 B.n391 71.676
R1728 B.n520 B.n392 71.676
R1729 B.n516 B.n393 71.676
R1730 B.n512 B.n394 71.676
R1731 B.n508 B.n395 71.676
R1732 B.n504 B.n396 71.676
R1733 B.n500 B.n397 71.676
R1734 B.n496 B.n398 71.676
R1735 B.n492 B.n399 71.676
R1736 B.n488 B.n400 71.676
R1737 B.n484 B.n401 71.676
R1738 B.n480 B.n402 71.676
R1739 B.n476 B.n403 71.676
R1740 B.n472 B.n404 71.676
R1741 B.n468 B.n405 71.676
R1742 B.n464 B.n406 71.676
R1743 B.n460 B.n407 71.676
R1744 B.n456 B.n408 71.676
R1745 B.n452 B.n409 71.676
R1746 B.n448 B.n410 71.676
R1747 B.n444 B.n411 71.676
R1748 B.n440 B.n412 71.676
R1749 B.n436 B.n413 71.676
R1750 B.n432 B.n414 71.676
R1751 B.n428 B.n415 71.676
R1752 B.n424 B.n416 71.676
R1753 B.n664 B.n663 71.676
R1754 B.n662 B.n355 61.5145
R1755 B.n725 B.n724 61.5145
R1756 B.n423 B.n422 59.5399
R1757 B.n550 B.n420 59.5399
R1758 B.n93 B.n92 59.5399
R1759 B.n224 B.n90 59.5399
R1760 B.n669 B.n355 34.0082
R1761 B.n669 B.n350 34.0082
R1762 B.n675 B.n350 34.0082
R1763 B.n675 B.n351 34.0082
R1764 B.n681 B.n343 34.0082
R1765 B.n687 B.n343 34.0082
R1766 B.n687 B.n339 34.0082
R1767 B.n695 B.n339 34.0082
R1768 B.n695 B.n694 34.0082
R1769 B.n701 B.n4 34.0082
R1770 B.n750 B.n4 34.0082
R1771 B.n750 B.n749 34.0082
R1772 B.n749 B.n748 34.0082
R1773 B.n742 B.n11 34.0082
R1774 B.n742 B.n741 34.0082
R1775 B.n741 B.n740 34.0082
R1776 B.n740 B.n15 34.0082
R1777 B.n734 B.n15 34.0082
R1778 B.n733 B.n732 34.0082
R1779 B.n732 B.n22 34.0082
R1780 B.n726 B.n22 34.0082
R1781 B.n726 B.n725 34.0082
R1782 B.n722 B.n721 30.1273
R1783 B.n95 B.n24 30.1273
R1784 B.n666 B.n665 30.1273
R1785 B.n659 B.n353 30.1273
R1786 B.n701 B.t0 28.0069
R1787 B.n748 B.t1 28.0069
R1788 B B.n752 18.0485
R1789 B.n351 B.t10 18.0046
R1790 B.t3 B.n733 18.0046
R1791 B.n422 B.n421 16.0975
R1792 B.n420 B.n419 16.0975
R1793 B.n92 B.n91 16.0975
R1794 B.n90 B.n89 16.0975
R1795 B.n681 B.t10 16.0041
R1796 B.n734 B.t3 16.0041
R1797 B.n96 B.n95 10.6151
R1798 B.n99 B.n96 10.6151
R1799 B.n100 B.n99 10.6151
R1800 B.n103 B.n100 10.6151
R1801 B.n104 B.n103 10.6151
R1802 B.n107 B.n104 10.6151
R1803 B.n108 B.n107 10.6151
R1804 B.n111 B.n108 10.6151
R1805 B.n112 B.n111 10.6151
R1806 B.n115 B.n112 10.6151
R1807 B.n116 B.n115 10.6151
R1808 B.n119 B.n116 10.6151
R1809 B.n120 B.n119 10.6151
R1810 B.n123 B.n120 10.6151
R1811 B.n124 B.n123 10.6151
R1812 B.n127 B.n124 10.6151
R1813 B.n128 B.n127 10.6151
R1814 B.n131 B.n128 10.6151
R1815 B.n132 B.n131 10.6151
R1816 B.n135 B.n132 10.6151
R1817 B.n136 B.n135 10.6151
R1818 B.n139 B.n136 10.6151
R1819 B.n140 B.n139 10.6151
R1820 B.n143 B.n140 10.6151
R1821 B.n144 B.n143 10.6151
R1822 B.n147 B.n144 10.6151
R1823 B.n148 B.n147 10.6151
R1824 B.n151 B.n148 10.6151
R1825 B.n152 B.n151 10.6151
R1826 B.n155 B.n152 10.6151
R1827 B.n156 B.n155 10.6151
R1828 B.n159 B.n156 10.6151
R1829 B.n160 B.n159 10.6151
R1830 B.n163 B.n160 10.6151
R1831 B.n164 B.n163 10.6151
R1832 B.n167 B.n164 10.6151
R1833 B.n168 B.n167 10.6151
R1834 B.n171 B.n168 10.6151
R1835 B.n172 B.n171 10.6151
R1836 B.n175 B.n172 10.6151
R1837 B.n176 B.n175 10.6151
R1838 B.n179 B.n176 10.6151
R1839 B.n180 B.n179 10.6151
R1840 B.n183 B.n180 10.6151
R1841 B.n184 B.n183 10.6151
R1842 B.n187 B.n184 10.6151
R1843 B.n188 B.n187 10.6151
R1844 B.n191 B.n188 10.6151
R1845 B.n192 B.n191 10.6151
R1846 B.n195 B.n192 10.6151
R1847 B.n196 B.n195 10.6151
R1848 B.n199 B.n196 10.6151
R1849 B.n200 B.n199 10.6151
R1850 B.n203 B.n200 10.6151
R1851 B.n204 B.n203 10.6151
R1852 B.n208 B.n207 10.6151
R1853 B.n211 B.n208 10.6151
R1854 B.n212 B.n211 10.6151
R1855 B.n215 B.n212 10.6151
R1856 B.n216 B.n215 10.6151
R1857 B.n219 B.n216 10.6151
R1858 B.n220 B.n219 10.6151
R1859 B.n223 B.n220 10.6151
R1860 B.n228 B.n225 10.6151
R1861 B.n229 B.n228 10.6151
R1862 B.n232 B.n229 10.6151
R1863 B.n233 B.n232 10.6151
R1864 B.n236 B.n233 10.6151
R1865 B.n237 B.n236 10.6151
R1866 B.n240 B.n237 10.6151
R1867 B.n241 B.n240 10.6151
R1868 B.n244 B.n241 10.6151
R1869 B.n245 B.n244 10.6151
R1870 B.n248 B.n245 10.6151
R1871 B.n249 B.n248 10.6151
R1872 B.n252 B.n249 10.6151
R1873 B.n253 B.n252 10.6151
R1874 B.n256 B.n253 10.6151
R1875 B.n257 B.n256 10.6151
R1876 B.n260 B.n257 10.6151
R1877 B.n261 B.n260 10.6151
R1878 B.n264 B.n261 10.6151
R1879 B.n265 B.n264 10.6151
R1880 B.n268 B.n265 10.6151
R1881 B.n269 B.n268 10.6151
R1882 B.n272 B.n269 10.6151
R1883 B.n273 B.n272 10.6151
R1884 B.n276 B.n273 10.6151
R1885 B.n277 B.n276 10.6151
R1886 B.n280 B.n277 10.6151
R1887 B.n281 B.n280 10.6151
R1888 B.n284 B.n281 10.6151
R1889 B.n285 B.n284 10.6151
R1890 B.n288 B.n285 10.6151
R1891 B.n289 B.n288 10.6151
R1892 B.n292 B.n289 10.6151
R1893 B.n293 B.n292 10.6151
R1894 B.n296 B.n293 10.6151
R1895 B.n297 B.n296 10.6151
R1896 B.n300 B.n297 10.6151
R1897 B.n301 B.n300 10.6151
R1898 B.n304 B.n301 10.6151
R1899 B.n305 B.n304 10.6151
R1900 B.n308 B.n305 10.6151
R1901 B.n309 B.n308 10.6151
R1902 B.n312 B.n309 10.6151
R1903 B.n313 B.n312 10.6151
R1904 B.n316 B.n313 10.6151
R1905 B.n317 B.n316 10.6151
R1906 B.n320 B.n317 10.6151
R1907 B.n321 B.n320 10.6151
R1908 B.n324 B.n321 10.6151
R1909 B.n325 B.n324 10.6151
R1910 B.n328 B.n325 10.6151
R1911 B.n329 B.n328 10.6151
R1912 B.n332 B.n329 10.6151
R1913 B.n333 B.n332 10.6151
R1914 B.n722 B.n333 10.6151
R1915 B.n667 B.n666 10.6151
R1916 B.n667 B.n348 10.6151
R1917 B.n677 B.n348 10.6151
R1918 B.n678 B.n677 10.6151
R1919 B.n679 B.n678 10.6151
R1920 B.n679 B.n341 10.6151
R1921 B.n689 B.n341 10.6151
R1922 B.n690 B.n689 10.6151
R1923 B.n692 B.n690 10.6151
R1924 B.n692 B.n691 10.6151
R1925 B.n691 B.n334 10.6151
R1926 B.n704 B.n334 10.6151
R1927 B.n705 B.n704 10.6151
R1928 B.n706 B.n705 10.6151
R1929 B.n707 B.n706 10.6151
R1930 B.n709 B.n707 10.6151
R1931 B.n710 B.n709 10.6151
R1932 B.n711 B.n710 10.6151
R1933 B.n712 B.n711 10.6151
R1934 B.n714 B.n712 10.6151
R1935 B.n715 B.n714 10.6151
R1936 B.n716 B.n715 10.6151
R1937 B.n717 B.n716 10.6151
R1938 B.n719 B.n717 10.6151
R1939 B.n720 B.n719 10.6151
R1940 B.n721 B.n720 10.6151
R1941 B.n659 B.n658 10.6151
R1942 B.n658 B.n657 10.6151
R1943 B.n657 B.n656 10.6151
R1944 B.n656 B.n654 10.6151
R1945 B.n654 B.n651 10.6151
R1946 B.n651 B.n650 10.6151
R1947 B.n650 B.n647 10.6151
R1948 B.n647 B.n646 10.6151
R1949 B.n646 B.n643 10.6151
R1950 B.n643 B.n642 10.6151
R1951 B.n642 B.n639 10.6151
R1952 B.n639 B.n638 10.6151
R1953 B.n638 B.n635 10.6151
R1954 B.n635 B.n634 10.6151
R1955 B.n634 B.n631 10.6151
R1956 B.n631 B.n630 10.6151
R1957 B.n630 B.n627 10.6151
R1958 B.n627 B.n626 10.6151
R1959 B.n626 B.n623 10.6151
R1960 B.n623 B.n622 10.6151
R1961 B.n622 B.n619 10.6151
R1962 B.n619 B.n618 10.6151
R1963 B.n618 B.n615 10.6151
R1964 B.n615 B.n614 10.6151
R1965 B.n614 B.n611 10.6151
R1966 B.n611 B.n610 10.6151
R1967 B.n610 B.n607 10.6151
R1968 B.n607 B.n606 10.6151
R1969 B.n606 B.n603 10.6151
R1970 B.n603 B.n602 10.6151
R1971 B.n602 B.n599 10.6151
R1972 B.n599 B.n598 10.6151
R1973 B.n598 B.n595 10.6151
R1974 B.n595 B.n594 10.6151
R1975 B.n594 B.n591 10.6151
R1976 B.n591 B.n590 10.6151
R1977 B.n590 B.n587 10.6151
R1978 B.n587 B.n586 10.6151
R1979 B.n586 B.n583 10.6151
R1980 B.n583 B.n582 10.6151
R1981 B.n582 B.n579 10.6151
R1982 B.n579 B.n578 10.6151
R1983 B.n578 B.n575 10.6151
R1984 B.n575 B.n574 10.6151
R1985 B.n574 B.n571 10.6151
R1986 B.n571 B.n570 10.6151
R1987 B.n570 B.n567 10.6151
R1988 B.n567 B.n566 10.6151
R1989 B.n566 B.n563 10.6151
R1990 B.n563 B.n562 10.6151
R1991 B.n562 B.n559 10.6151
R1992 B.n559 B.n558 10.6151
R1993 B.n558 B.n555 10.6151
R1994 B.n555 B.n554 10.6151
R1995 B.n554 B.n551 10.6151
R1996 B.n549 B.n546 10.6151
R1997 B.n546 B.n545 10.6151
R1998 B.n545 B.n542 10.6151
R1999 B.n542 B.n541 10.6151
R2000 B.n541 B.n538 10.6151
R2001 B.n538 B.n537 10.6151
R2002 B.n537 B.n534 10.6151
R2003 B.n534 B.n533 10.6151
R2004 B.n530 B.n529 10.6151
R2005 B.n529 B.n526 10.6151
R2006 B.n526 B.n525 10.6151
R2007 B.n525 B.n522 10.6151
R2008 B.n522 B.n521 10.6151
R2009 B.n521 B.n518 10.6151
R2010 B.n518 B.n517 10.6151
R2011 B.n517 B.n514 10.6151
R2012 B.n514 B.n513 10.6151
R2013 B.n513 B.n510 10.6151
R2014 B.n510 B.n509 10.6151
R2015 B.n509 B.n506 10.6151
R2016 B.n506 B.n505 10.6151
R2017 B.n505 B.n502 10.6151
R2018 B.n502 B.n501 10.6151
R2019 B.n501 B.n498 10.6151
R2020 B.n498 B.n497 10.6151
R2021 B.n497 B.n494 10.6151
R2022 B.n494 B.n493 10.6151
R2023 B.n493 B.n490 10.6151
R2024 B.n490 B.n489 10.6151
R2025 B.n489 B.n486 10.6151
R2026 B.n486 B.n485 10.6151
R2027 B.n485 B.n482 10.6151
R2028 B.n482 B.n481 10.6151
R2029 B.n481 B.n478 10.6151
R2030 B.n478 B.n477 10.6151
R2031 B.n477 B.n474 10.6151
R2032 B.n474 B.n473 10.6151
R2033 B.n473 B.n470 10.6151
R2034 B.n470 B.n469 10.6151
R2035 B.n469 B.n466 10.6151
R2036 B.n466 B.n465 10.6151
R2037 B.n465 B.n462 10.6151
R2038 B.n462 B.n461 10.6151
R2039 B.n461 B.n458 10.6151
R2040 B.n458 B.n457 10.6151
R2041 B.n457 B.n454 10.6151
R2042 B.n454 B.n453 10.6151
R2043 B.n453 B.n450 10.6151
R2044 B.n450 B.n449 10.6151
R2045 B.n449 B.n446 10.6151
R2046 B.n446 B.n445 10.6151
R2047 B.n445 B.n442 10.6151
R2048 B.n442 B.n441 10.6151
R2049 B.n441 B.n438 10.6151
R2050 B.n438 B.n437 10.6151
R2051 B.n437 B.n434 10.6151
R2052 B.n434 B.n433 10.6151
R2053 B.n433 B.n430 10.6151
R2054 B.n430 B.n429 10.6151
R2055 B.n429 B.n426 10.6151
R2056 B.n426 B.n425 10.6151
R2057 B.n425 B.n357 10.6151
R2058 B.n665 B.n357 10.6151
R2059 B.n671 B.n353 10.6151
R2060 B.n672 B.n671 10.6151
R2061 B.n673 B.n672 10.6151
R2062 B.n673 B.n345 10.6151
R2063 B.n683 B.n345 10.6151
R2064 B.n684 B.n683 10.6151
R2065 B.n685 B.n684 10.6151
R2066 B.n685 B.n337 10.6151
R2067 B.n697 B.n337 10.6151
R2068 B.n698 B.n697 10.6151
R2069 B.n699 B.n698 10.6151
R2070 B.n699 B.n0 10.6151
R2071 B.n746 B.n1 10.6151
R2072 B.n746 B.n745 10.6151
R2073 B.n745 B.n744 10.6151
R2074 B.n744 B.n9 10.6151
R2075 B.n738 B.n9 10.6151
R2076 B.n738 B.n737 10.6151
R2077 B.n737 B.n736 10.6151
R2078 B.n736 B.n17 10.6151
R2079 B.n730 B.n17 10.6151
R2080 B.n730 B.n729 10.6151
R2081 B.n729 B.n728 10.6151
R2082 B.n728 B.n24 10.6151
R2083 B.n207 B.n93 7.18099
R2084 B.n224 B.n223 7.18099
R2085 B.n550 B.n549 7.18099
R2086 B.n533 B.n423 7.18099
R2087 B.n694 B.t0 6.00186
R2088 B.n11 B.t1 6.00186
R2089 B.n204 B.n93 3.43465
R2090 B.n225 B.n224 3.43465
R2091 B.n551 B.n550 3.43465
R2092 B.n530 B.n423 3.43465
R2093 B.n752 B.n0 2.81026
R2094 B.n752 B.n1 2.81026
R2095 VP.n0 VP.t1 1087.47
R2096 VP.n0 VP.t0 1044.81
R2097 VP VP.n0 0.0516364
R2098 VDD1.n88 VDD1.n0 289.615
R2099 VDD1.n181 VDD1.n93 289.615
R2100 VDD1.n89 VDD1.n88 185
R2101 VDD1.n87 VDD1.n86 185
R2102 VDD1.n4 VDD1.n3 185
R2103 VDD1.n81 VDD1.n80 185
R2104 VDD1.n79 VDD1.n78 185
R2105 VDD1.n77 VDD1.n7 185
R2106 VDD1.n11 VDD1.n8 185
R2107 VDD1.n72 VDD1.n71 185
R2108 VDD1.n70 VDD1.n69 185
R2109 VDD1.n13 VDD1.n12 185
R2110 VDD1.n64 VDD1.n63 185
R2111 VDD1.n62 VDD1.n61 185
R2112 VDD1.n17 VDD1.n16 185
R2113 VDD1.n56 VDD1.n55 185
R2114 VDD1.n54 VDD1.n53 185
R2115 VDD1.n21 VDD1.n20 185
R2116 VDD1.n48 VDD1.n47 185
R2117 VDD1.n46 VDD1.n45 185
R2118 VDD1.n25 VDD1.n24 185
R2119 VDD1.n40 VDD1.n39 185
R2120 VDD1.n38 VDD1.n37 185
R2121 VDD1.n29 VDD1.n28 185
R2122 VDD1.n32 VDD1.n31 185
R2123 VDD1.n124 VDD1.n123 185
R2124 VDD1.n121 VDD1.n120 185
R2125 VDD1.n130 VDD1.n129 185
R2126 VDD1.n132 VDD1.n131 185
R2127 VDD1.n117 VDD1.n116 185
R2128 VDD1.n138 VDD1.n137 185
R2129 VDD1.n140 VDD1.n139 185
R2130 VDD1.n113 VDD1.n112 185
R2131 VDD1.n146 VDD1.n145 185
R2132 VDD1.n148 VDD1.n147 185
R2133 VDD1.n109 VDD1.n108 185
R2134 VDD1.n154 VDD1.n153 185
R2135 VDD1.n156 VDD1.n155 185
R2136 VDD1.n105 VDD1.n104 185
R2137 VDD1.n162 VDD1.n161 185
R2138 VDD1.n165 VDD1.n164 185
R2139 VDD1.n163 VDD1.n101 185
R2140 VDD1.n170 VDD1.n100 185
R2141 VDD1.n172 VDD1.n171 185
R2142 VDD1.n174 VDD1.n173 185
R2143 VDD1.n97 VDD1.n96 185
R2144 VDD1.n180 VDD1.n179 185
R2145 VDD1.n182 VDD1.n181 185
R2146 VDD1.t0 VDD1.n30 147.659
R2147 VDD1.t1 VDD1.n122 147.659
R2148 VDD1.n88 VDD1.n87 104.615
R2149 VDD1.n87 VDD1.n3 104.615
R2150 VDD1.n80 VDD1.n3 104.615
R2151 VDD1.n80 VDD1.n79 104.615
R2152 VDD1.n79 VDD1.n7 104.615
R2153 VDD1.n11 VDD1.n7 104.615
R2154 VDD1.n71 VDD1.n11 104.615
R2155 VDD1.n71 VDD1.n70 104.615
R2156 VDD1.n70 VDD1.n12 104.615
R2157 VDD1.n63 VDD1.n12 104.615
R2158 VDD1.n63 VDD1.n62 104.615
R2159 VDD1.n62 VDD1.n16 104.615
R2160 VDD1.n55 VDD1.n16 104.615
R2161 VDD1.n55 VDD1.n54 104.615
R2162 VDD1.n54 VDD1.n20 104.615
R2163 VDD1.n47 VDD1.n20 104.615
R2164 VDD1.n47 VDD1.n46 104.615
R2165 VDD1.n46 VDD1.n24 104.615
R2166 VDD1.n39 VDD1.n24 104.615
R2167 VDD1.n39 VDD1.n38 104.615
R2168 VDD1.n38 VDD1.n28 104.615
R2169 VDD1.n31 VDD1.n28 104.615
R2170 VDD1.n123 VDD1.n120 104.615
R2171 VDD1.n130 VDD1.n120 104.615
R2172 VDD1.n131 VDD1.n130 104.615
R2173 VDD1.n131 VDD1.n116 104.615
R2174 VDD1.n138 VDD1.n116 104.615
R2175 VDD1.n139 VDD1.n138 104.615
R2176 VDD1.n139 VDD1.n112 104.615
R2177 VDD1.n146 VDD1.n112 104.615
R2178 VDD1.n147 VDD1.n146 104.615
R2179 VDD1.n147 VDD1.n108 104.615
R2180 VDD1.n154 VDD1.n108 104.615
R2181 VDD1.n155 VDD1.n154 104.615
R2182 VDD1.n155 VDD1.n104 104.615
R2183 VDD1.n162 VDD1.n104 104.615
R2184 VDD1.n164 VDD1.n162 104.615
R2185 VDD1.n164 VDD1.n163 104.615
R2186 VDD1.n163 VDD1.n100 104.615
R2187 VDD1.n172 VDD1.n100 104.615
R2188 VDD1.n173 VDD1.n172 104.615
R2189 VDD1.n173 VDD1.n96 104.615
R2190 VDD1.n180 VDD1.n96 104.615
R2191 VDD1.n181 VDD1.n180 104.615
R2192 VDD1 VDD1.n185 87.1327
R2193 VDD1.n31 VDD1.t0 52.3082
R2194 VDD1.n123 VDD1.t1 52.3082
R2195 VDD1 VDD1.n92 47.1618
R2196 VDD1.n32 VDD1.n30 15.6677
R2197 VDD1.n124 VDD1.n122 15.6677
R2198 VDD1.n78 VDD1.n77 13.1884
R2199 VDD1.n171 VDD1.n170 13.1884
R2200 VDD1.n81 VDD1.n6 12.8005
R2201 VDD1.n76 VDD1.n8 12.8005
R2202 VDD1.n33 VDD1.n29 12.8005
R2203 VDD1.n125 VDD1.n121 12.8005
R2204 VDD1.n169 VDD1.n101 12.8005
R2205 VDD1.n174 VDD1.n99 12.8005
R2206 VDD1.n82 VDD1.n4 12.0247
R2207 VDD1.n73 VDD1.n72 12.0247
R2208 VDD1.n37 VDD1.n36 12.0247
R2209 VDD1.n129 VDD1.n128 12.0247
R2210 VDD1.n166 VDD1.n165 12.0247
R2211 VDD1.n175 VDD1.n97 12.0247
R2212 VDD1.n86 VDD1.n85 11.249
R2213 VDD1.n69 VDD1.n10 11.249
R2214 VDD1.n40 VDD1.n27 11.249
R2215 VDD1.n132 VDD1.n119 11.249
R2216 VDD1.n161 VDD1.n103 11.249
R2217 VDD1.n179 VDD1.n178 11.249
R2218 VDD1.n89 VDD1.n2 10.4732
R2219 VDD1.n68 VDD1.n13 10.4732
R2220 VDD1.n41 VDD1.n25 10.4732
R2221 VDD1.n133 VDD1.n117 10.4732
R2222 VDD1.n160 VDD1.n105 10.4732
R2223 VDD1.n182 VDD1.n95 10.4732
R2224 VDD1.n90 VDD1.n0 9.69747
R2225 VDD1.n65 VDD1.n64 9.69747
R2226 VDD1.n45 VDD1.n44 9.69747
R2227 VDD1.n137 VDD1.n136 9.69747
R2228 VDD1.n157 VDD1.n156 9.69747
R2229 VDD1.n183 VDD1.n93 9.69747
R2230 VDD1.n92 VDD1.n91 9.45567
R2231 VDD1.n185 VDD1.n184 9.45567
R2232 VDD1.n58 VDD1.n57 9.3005
R2233 VDD1.n60 VDD1.n59 9.3005
R2234 VDD1.n15 VDD1.n14 9.3005
R2235 VDD1.n66 VDD1.n65 9.3005
R2236 VDD1.n68 VDD1.n67 9.3005
R2237 VDD1.n10 VDD1.n9 9.3005
R2238 VDD1.n74 VDD1.n73 9.3005
R2239 VDD1.n76 VDD1.n75 9.3005
R2240 VDD1.n91 VDD1.n90 9.3005
R2241 VDD1.n2 VDD1.n1 9.3005
R2242 VDD1.n85 VDD1.n84 9.3005
R2243 VDD1.n83 VDD1.n82 9.3005
R2244 VDD1.n6 VDD1.n5 9.3005
R2245 VDD1.n19 VDD1.n18 9.3005
R2246 VDD1.n52 VDD1.n51 9.3005
R2247 VDD1.n50 VDD1.n49 9.3005
R2248 VDD1.n23 VDD1.n22 9.3005
R2249 VDD1.n44 VDD1.n43 9.3005
R2250 VDD1.n42 VDD1.n41 9.3005
R2251 VDD1.n27 VDD1.n26 9.3005
R2252 VDD1.n36 VDD1.n35 9.3005
R2253 VDD1.n34 VDD1.n33 9.3005
R2254 VDD1.n184 VDD1.n183 9.3005
R2255 VDD1.n95 VDD1.n94 9.3005
R2256 VDD1.n178 VDD1.n177 9.3005
R2257 VDD1.n176 VDD1.n175 9.3005
R2258 VDD1.n99 VDD1.n98 9.3005
R2259 VDD1.n144 VDD1.n143 9.3005
R2260 VDD1.n142 VDD1.n141 9.3005
R2261 VDD1.n115 VDD1.n114 9.3005
R2262 VDD1.n136 VDD1.n135 9.3005
R2263 VDD1.n134 VDD1.n133 9.3005
R2264 VDD1.n119 VDD1.n118 9.3005
R2265 VDD1.n128 VDD1.n127 9.3005
R2266 VDD1.n126 VDD1.n125 9.3005
R2267 VDD1.n111 VDD1.n110 9.3005
R2268 VDD1.n150 VDD1.n149 9.3005
R2269 VDD1.n152 VDD1.n151 9.3005
R2270 VDD1.n107 VDD1.n106 9.3005
R2271 VDD1.n158 VDD1.n157 9.3005
R2272 VDD1.n160 VDD1.n159 9.3005
R2273 VDD1.n103 VDD1.n102 9.3005
R2274 VDD1.n167 VDD1.n166 9.3005
R2275 VDD1.n169 VDD1.n168 9.3005
R2276 VDD1.n61 VDD1.n15 8.92171
R2277 VDD1.n48 VDD1.n23 8.92171
R2278 VDD1.n140 VDD1.n115 8.92171
R2279 VDD1.n153 VDD1.n107 8.92171
R2280 VDD1.n60 VDD1.n17 8.14595
R2281 VDD1.n49 VDD1.n21 8.14595
R2282 VDD1.n141 VDD1.n113 8.14595
R2283 VDD1.n152 VDD1.n109 8.14595
R2284 VDD1.n57 VDD1.n56 7.3702
R2285 VDD1.n53 VDD1.n52 7.3702
R2286 VDD1.n145 VDD1.n144 7.3702
R2287 VDD1.n149 VDD1.n148 7.3702
R2288 VDD1.n56 VDD1.n19 6.59444
R2289 VDD1.n53 VDD1.n19 6.59444
R2290 VDD1.n145 VDD1.n111 6.59444
R2291 VDD1.n148 VDD1.n111 6.59444
R2292 VDD1.n57 VDD1.n17 5.81868
R2293 VDD1.n52 VDD1.n21 5.81868
R2294 VDD1.n144 VDD1.n113 5.81868
R2295 VDD1.n149 VDD1.n109 5.81868
R2296 VDD1.n61 VDD1.n60 5.04292
R2297 VDD1.n49 VDD1.n48 5.04292
R2298 VDD1.n141 VDD1.n140 5.04292
R2299 VDD1.n153 VDD1.n152 5.04292
R2300 VDD1.n34 VDD1.n30 4.38563
R2301 VDD1.n126 VDD1.n122 4.38563
R2302 VDD1.n92 VDD1.n0 4.26717
R2303 VDD1.n64 VDD1.n15 4.26717
R2304 VDD1.n45 VDD1.n23 4.26717
R2305 VDD1.n137 VDD1.n115 4.26717
R2306 VDD1.n156 VDD1.n107 4.26717
R2307 VDD1.n185 VDD1.n93 4.26717
R2308 VDD1.n90 VDD1.n89 3.49141
R2309 VDD1.n65 VDD1.n13 3.49141
R2310 VDD1.n44 VDD1.n25 3.49141
R2311 VDD1.n136 VDD1.n117 3.49141
R2312 VDD1.n157 VDD1.n105 3.49141
R2313 VDD1.n183 VDD1.n182 3.49141
R2314 VDD1.n86 VDD1.n2 2.71565
R2315 VDD1.n69 VDD1.n68 2.71565
R2316 VDD1.n41 VDD1.n40 2.71565
R2317 VDD1.n133 VDD1.n132 2.71565
R2318 VDD1.n161 VDD1.n160 2.71565
R2319 VDD1.n179 VDD1.n95 2.71565
R2320 VDD1.n85 VDD1.n4 1.93989
R2321 VDD1.n72 VDD1.n10 1.93989
R2322 VDD1.n37 VDD1.n27 1.93989
R2323 VDD1.n129 VDD1.n119 1.93989
R2324 VDD1.n165 VDD1.n103 1.93989
R2325 VDD1.n178 VDD1.n97 1.93989
R2326 VDD1.n82 VDD1.n81 1.16414
R2327 VDD1.n73 VDD1.n8 1.16414
R2328 VDD1.n36 VDD1.n29 1.16414
R2329 VDD1.n128 VDD1.n121 1.16414
R2330 VDD1.n166 VDD1.n101 1.16414
R2331 VDD1.n175 VDD1.n174 1.16414
R2332 VDD1.n78 VDD1.n6 0.388379
R2333 VDD1.n77 VDD1.n76 0.388379
R2334 VDD1.n33 VDD1.n32 0.388379
R2335 VDD1.n125 VDD1.n124 0.388379
R2336 VDD1.n170 VDD1.n169 0.388379
R2337 VDD1.n171 VDD1.n99 0.388379
R2338 VDD1.n91 VDD1.n1 0.155672
R2339 VDD1.n84 VDD1.n1 0.155672
R2340 VDD1.n84 VDD1.n83 0.155672
R2341 VDD1.n83 VDD1.n5 0.155672
R2342 VDD1.n75 VDD1.n5 0.155672
R2343 VDD1.n75 VDD1.n74 0.155672
R2344 VDD1.n74 VDD1.n9 0.155672
R2345 VDD1.n67 VDD1.n9 0.155672
R2346 VDD1.n67 VDD1.n66 0.155672
R2347 VDD1.n66 VDD1.n14 0.155672
R2348 VDD1.n59 VDD1.n14 0.155672
R2349 VDD1.n59 VDD1.n58 0.155672
R2350 VDD1.n58 VDD1.n18 0.155672
R2351 VDD1.n51 VDD1.n18 0.155672
R2352 VDD1.n51 VDD1.n50 0.155672
R2353 VDD1.n50 VDD1.n22 0.155672
R2354 VDD1.n43 VDD1.n22 0.155672
R2355 VDD1.n43 VDD1.n42 0.155672
R2356 VDD1.n42 VDD1.n26 0.155672
R2357 VDD1.n35 VDD1.n26 0.155672
R2358 VDD1.n35 VDD1.n34 0.155672
R2359 VDD1.n127 VDD1.n126 0.155672
R2360 VDD1.n127 VDD1.n118 0.155672
R2361 VDD1.n134 VDD1.n118 0.155672
R2362 VDD1.n135 VDD1.n134 0.155672
R2363 VDD1.n135 VDD1.n114 0.155672
R2364 VDD1.n142 VDD1.n114 0.155672
R2365 VDD1.n143 VDD1.n142 0.155672
R2366 VDD1.n143 VDD1.n110 0.155672
R2367 VDD1.n150 VDD1.n110 0.155672
R2368 VDD1.n151 VDD1.n150 0.155672
R2369 VDD1.n151 VDD1.n106 0.155672
R2370 VDD1.n158 VDD1.n106 0.155672
R2371 VDD1.n159 VDD1.n158 0.155672
R2372 VDD1.n159 VDD1.n102 0.155672
R2373 VDD1.n167 VDD1.n102 0.155672
R2374 VDD1.n168 VDD1.n167 0.155672
R2375 VDD1.n168 VDD1.n98 0.155672
R2376 VDD1.n176 VDD1.n98 0.155672
R2377 VDD1.n177 VDD1.n176 0.155672
R2378 VDD1.n177 VDD1.n94 0.155672
R2379 VDD1.n184 VDD1.n94 0.155672
C0 VDD1 VTAIL 8.040461f
C1 VN VTAIL 1.59051f
C2 VP VDD2 0.247813f
C3 VP VDD1 2.44127f
C4 VP VN 5.33965f
C5 VP VTAIL 1.60541f
C6 VDD1 VDD2 0.445151f
C7 VDD2 VN 2.34877f
C8 VDD2 VTAIL 8.069139f
C9 VDD1 VN 0.148831f
C10 VDD2 B 4.528234f
C11 VDD1 B 7.3743f
C12 VTAIL B 7.437111f
C13 VN B 9.187901f
C14 VP B 4.109175f
C15 VDD1.n0 B 0.027568f
C16 VDD1.n1 B 0.021468f
C17 VDD1.n2 B 0.011536f
C18 VDD1.n3 B 0.027267f
C19 VDD1.n4 B 0.012215f
C20 VDD1.n5 B 0.021468f
C21 VDD1.n6 B 0.011536f
C22 VDD1.n7 B 0.027267f
C23 VDD1.n8 B 0.012215f
C24 VDD1.n9 B 0.021468f
C25 VDD1.n10 B 0.011536f
C26 VDD1.n11 B 0.027267f
C27 VDD1.n12 B 0.027267f
C28 VDD1.n13 B 0.012215f
C29 VDD1.n14 B 0.021468f
C30 VDD1.n15 B 0.011536f
C31 VDD1.n16 B 0.027267f
C32 VDD1.n17 B 0.012215f
C33 VDD1.n18 B 0.021468f
C34 VDD1.n19 B 0.011536f
C35 VDD1.n20 B 0.027267f
C36 VDD1.n21 B 0.012215f
C37 VDD1.n22 B 0.021468f
C38 VDD1.n23 B 0.011536f
C39 VDD1.n24 B 0.027267f
C40 VDD1.n25 B 0.012215f
C41 VDD1.n26 B 0.021468f
C42 VDD1.n27 B 0.011536f
C43 VDD1.n28 B 0.027267f
C44 VDD1.n29 B 0.012215f
C45 VDD1.n30 B 0.149171f
C46 VDD1.t0 B 0.045085f
C47 VDD1.n31 B 0.02045f
C48 VDD1.n32 B 0.016107f
C49 VDD1.n33 B 0.011536f
C50 VDD1.n34 B 1.56401f
C51 VDD1.n35 B 0.021468f
C52 VDD1.n36 B 0.011536f
C53 VDD1.n37 B 0.012215f
C54 VDD1.n38 B 0.027267f
C55 VDD1.n39 B 0.027267f
C56 VDD1.n40 B 0.012215f
C57 VDD1.n41 B 0.011536f
C58 VDD1.n42 B 0.021468f
C59 VDD1.n43 B 0.021468f
C60 VDD1.n44 B 0.011536f
C61 VDD1.n45 B 0.012215f
C62 VDD1.n46 B 0.027267f
C63 VDD1.n47 B 0.027267f
C64 VDD1.n48 B 0.012215f
C65 VDD1.n49 B 0.011536f
C66 VDD1.n50 B 0.021468f
C67 VDD1.n51 B 0.021468f
C68 VDD1.n52 B 0.011536f
C69 VDD1.n53 B 0.012215f
C70 VDD1.n54 B 0.027267f
C71 VDD1.n55 B 0.027267f
C72 VDD1.n56 B 0.012215f
C73 VDD1.n57 B 0.011536f
C74 VDD1.n58 B 0.021468f
C75 VDD1.n59 B 0.021468f
C76 VDD1.n60 B 0.011536f
C77 VDD1.n61 B 0.012215f
C78 VDD1.n62 B 0.027267f
C79 VDD1.n63 B 0.027267f
C80 VDD1.n64 B 0.012215f
C81 VDD1.n65 B 0.011536f
C82 VDD1.n66 B 0.021468f
C83 VDD1.n67 B 0.021468f
C84 VDD1.n68 B 0.011536f
C85 VDD1.n69 B 0.012215f
C86 VDD1.n70 B 0.027267f
C87 VDD1.n71 B 0.027267f
C88 VDD1.n72 B 0.012215f
C89 VDD1.n73 B 0.011536f
C90 VDD1.n74 B 0.021468f
C91 VDD1.n75 B 0.021468f
C92 VDD1.n76 B 0.011536f
C93 VDD1.n77 B 0.011875f
C94 VDD1.n78 B 0.011875f
C95 VDD1.n79 B 0.027267f
C96 VDD1.n80 B 0.027267f
C97 VDD1.n81 B 0.012215f
C98 VDD1.n82 B 0.011536f
C99 VDD1.n83 B 0.021468f
C100 VDD1.n84 B 0.021468f
C101 VDD1.n85 B 0.011536f
C102 VDD1.n86 B 0.012215f
C103 VDD1.n87 B 0.027267f
C104 VDD1.n88 B 0.054418f
C105 VDD1.n89 B 0.012215f
C106 VDD1.n90 B 0.011536f
C107 VDD1.n91 B 0.04669f
C108 VDD1.n92 B 0.045013f
C109 VDD1.n93 B 0.027568f
C110 VDD1.n94 B 0.021468f
C111 VDD1.n95 B 0.011536f
C112 VDD1.n96 B 0.027267f
C113 VDD1.n97 B 0.012215f
C114 VDD1.n98 B 0.021468f
C115 VDD1.n99 B 0.011536f
C116 VDD1.n100 B 0.027267f
C117 VDD1.n101 B 0.012215f
C118 VDD1.n102 B 0.021468f
C119 VDD1.n103 B 0.011536f
C120 VDD1.n104 B 0.027267f
C121 VDD1.n105 B 0.012215f
C122 VDD1.n106 B 0.021468f
C123 VDD1.n107 B 0.011536f
C124 VDD1.n108 B 0.027267f
C125 VDD1.n109 B 0.012215f
C126 VDD1.n110 B 0.021468f
C127 VDD1.n111 B 0.011536f
C128 VDD1.n112 B 0.027267f
C129 VDD1.n113 B 0.012215f
C130 VDD1.n114 B 0.021468f
C131 VDD1.n115 B 0.011536f
C132 VDD1.n116 B 0.027267f
C133 VDD1.n117 B 0.012215f
C134 VDD1.n118 B 0.021468f
C135 VDD1.n119 B 0.011536f
C136 VDD1.n120 B 0.027267f
C137 VDD1.n121 B 0.012215f
C138 VDD1.n122 B 0.149171f
C139 VDD1.t1 B 0.045085f
C140 VDD1.n123 B 0.02045f
C141 VDD1.n124 B 0.016107f
C142 VDD1.n125 B 0.011536f
C143 VDD1.n126 B 1.56401f
C144 VDD1.n127 B 0.021468f
C145 VDD1.n128 B 0.011536f
C146 VDD1.n129 B 0.012215f
C147 VDD1.n130 B 0.027267f
C148 VDD1.n131 B 0.027267f
C149 VDD1.n132 B 0.012215f
C150 VDD1.n133 B 0.011536f
C151 VDD1.n134 B 0.021468f
C152 VDD1.n135 B 0.021468f
C153 VDD1.n136 B 0.011536f
C154 VDD1.n137 B 0.012215f
C155 VDD1.n138 B 0.027267f
C156 VDD1.n139 B 0.027267f
C157 VDD1.n140 B 0.012215f
C158 VDD1.n141 B 0.011536f
C159 VDD1.n142 B 0.021468f
C160 VDD1.n143 B 0.021468f
C161 VDD1.n144 B 0.011536f
C162 VDD1.n145 B 0.012215f
C163 VDD1.n146 B 0.027267f
C164 VDD1.n147 B 0.027267f
C165 VDD1.n148 B 0.012215f
C166 VDD1.n149 B 0.011536f
C167 VDD1.n150 B 0.021468f
C168 VDD1.n151 B 0.021468f
C169 VDD1.n152 B 0.011536f
C170 VDD1.n153 B 0.012215f
C171 VDD1.n154 B 0.027267f
C172 VDD1.n155 B 0.027267f
C173 VDD1.n156 B 0.012215f
C174 VDD1.n157 B 0.011536f
C175 VDD1.n158 B 0.021468f
C176 VDD1.n159 B 0.021468f
C177 VDD1.n160 B 0.011536f
C178 VDD1.n161 B 0.012215f
C179 VDD1.n162 B 0.027267f
C180 VDD1.n163 B 0.027267f
C181 VDD1.n164 B 0.027267f
C182 VDD1.n165 B 0.012215f
C183 VDD1.n166 B 0.011536f
C184 VDD1.n167 B 0.021468f
C185 VDD1.n168 B 0.021468f
C186 VDD1.n169 B 0.011536f
C187 VDD1.n170 B 0.011875f
C188 VDD1.n171 B 0.011875f
C189 VDD1.n172 B 0.027267f
C190 VDD1.n173 B 0.027267f
C191 VDD1.n174 B 0.012215f
C192 VDD1.n175 B 0.011536f
C193 VDD1.n176 B 0.021468f
C194 VDD1.n177 B 0.021468f
C195 VDD1.n178 B 0.011536f
C196 VDD1.n179 B 0.012215f
C197 VDD1.n180 B 0.027267f
C198 VDD1.n181 B 0.054418f
C199 VDD1.n182 B 0.012215f
C200 VDD1.n183 B 0.011536f
C201 VDD1.n184 B 0.04669f
C202 VDD1.n185 B 0.697019f
C203 VP.t1 B 1.3804f
C204 VP.t0 B 1.28045f
C205 VP.n0 B 5.02765f
C206 VDD2.n0 B 0.02778f
C207 VDD2.n1 B 0.021633f
C208 VDD2.n2 B 0.011625f
C209 VDD2.n3 B 0.027477f
C210 VDD2.n4 B 0.012309f
C211 VDD2.n5 B 0.021633f
C212 VDD2.n6 B 0.011625f
C213 VDD2.n7 B 0.027477f
C214 VDD2.n8 B 0.012309f
C215 VDD2.n9 B 0.021633f
C216 VDD2.n10 B 0.011625f
C217 VDD2.n11 B 0.027477f
C218 VDD2.n12 B 0.012309f
C219 VDD2.n13 B 0.021633f
C220 VDD2.n14 B 0.011625f
C221 VDD2.n15 B 0.027477f
C222 VDD2.n16 B 0.012309f
C223 VDD2.n17 B 0.021633f
C224 VDD2.n18 B 0.011625f
C225 VDD2.n19 B 0.027477f
C226 VDD2.n20 B 0.012309f
C227 VDD2.n21 B 0.021633f
C228 VDD2.n22 B 0.011625f
C229 VDD2.n23 B 0.027477f
C230 VDD2.n24 B 0.012309f
C231 VDD2.n25 B 0.021633f
C232 VDD2.n26 B 0.011625f
C233 VDD2.n27 B 0.027477f
C234 VDD2.n28 B 0.012309f
C235 VDD2.n29 B 0.150317f
C236 VDD2.t0 B 0.045432f
C237 VDD2.n30 B 0.020607f
C238 VDD2.n31 B 0.016231f
C239 VDD2.n32 B 0.011625f
C240 VDD2.n33 B 1.57603f
C241 VDD2.n34 B 0.021633f
C242 VDD2.n35 B 0.011625f
C243 VDD2.n36 B 0.012309f
C244 VDD2.n37 B 0.027477f
C245 VDD2.n38 B 0.027477f
C246 VDD2.n39 B 0.012309f
C247 VDD2.n40 B 0.011625f
C248 VDD2.n41 B 0.021633f
C249 VDD2.n42 B 0.021633f
C250 VDD2.n43 B 0.011625f
C251 VDD2.n44 B 0.012309f
C252 VDD2.n45 B 0.027477f
C253 VDD2.n46 B 0.027477f
C254 VDD2.n47 B 0.012309f
C255 VDD2.n48 B 0.011625f
C256 VDD2.n49 B 0.021633f
C257 VDD2.n50 B 0.021633f
C258 VDD2.n51 B 0.011625f
C259 VDD2.n52 B 0.012309f
C260 VDD2.n53 B 0.027477f
C261 VDD2.n54 B 0.027477f
C262 VDD2.n55 B 0.012309f
C263 VDD2.n56 B 0.011625f
C264 VDD2.n57 B 0.021633f
C265 VDD2.n58 B 0.021633f
C266 VDD2.n59 B 0.011625f
C267 VDD2.n60 B 0.012309f
C268 VDD2.n61 B 0.027477f
C269 VDD2.n62 B 0.027477f
C270 VDD2.n63 B 0.012309f
C271 VDD2.n64 B 0.011625f
C272 VDD2.n65 B 0.021633f
C273 VDD2.n66 B 0.021633f
C274 VDD2.n67 B 0.011625f
C275 VDD2.n68 B 0.012309f
C276 VDD2.n69 B 0.027477f
C277 VDD2.n70 B 0.027477f
C278 VDD2.n71 B 0.027477f
C279 VDD2.n72 B 0.012309f
C280 VDD2.n73 B 0.011625f
C281 VDD2.n74 B 0.021633f
C282 VDD2.n75 B 0.021633f
C283 VDD2.n76 B 0.011625f
C284 VDD2.n77 B 0.011967f
C285 VDD2.n78 B 0.011967f
C286 VDD2.n79 B 0.027477f
C287 VDD2.n80 B 0.027477f
C288 VDD2.n81 B 0.012309f
C289 VDD2.n82 B 0.011625f
C290 VDD2.n83 B 0.021633f
C291 VDD2.n84 B 0.021633f
C292 VDD2.n85 B 0.011625f
C293 VDD2.n86 B 0.012309f
C294 VDD2.n87 B 0.027477f
C295 VDD2.n88 B 0.054836f
C296 VDD2.n89 B 0.012309f
C297 VDD2.n90 B 0.011625f
C298 VDD2.n91 B 0.047049f
C299 VDD2.n92 B 0.672273f
C300 VDD2.n93 B 0.02778f
C301 VDD2.n94 B 0.021633f
C302 VDD2.n95 B 0.011625f
C303 VDD2.n96 B 0.027477f
C304 VDD2.n97 B 0.012309f
C305 VDD2.n98 B 0.021633f
C306 VDD2.n99 B 0.011625f
C307 VDD2.n100 B 0.027477f
C308 VDD2.n101 B 0.012309f
C309 VDD2.n102 B 0.021633f
C310 VDD2.n103 B 0.011625f
C311 VDD2.n104 B 0.027477f
C312 VDD2.n105 B 0.027477f
C313 VDD2.n106 B 0.012309f
C314 VDD2.n107 B 0.021633f
C315 VDD2.n108 B 0.011625f
C316 VDD2.n109 B 0.027477f
C317 VDD2.n110 B 0.012309f
C318 VDD2.n111 B 0.021633f
C319 VDD2.n112 B 0.011625f
C320 VDD2.n113 B 0.027477f
C321 VDD2.n114 B 0.012309f
C322 VDD2.n115 B 0.021633f
C323 VDD2.n116 B 0.011625f
C324 VDD2.n117 B 0.027477f
C325 VDD2.n118 B 0.012309f
C326 VDD2.n119 B 0.021633f
C327 VDD2.n120 B 0.011625f
C328 VDD2.n121 B 0.027477f
C329 VDD2.n122 B 0.012309f
C330 VDD2.n123 B 0.150317f
C331 VDD2.t1 B 0.045432f
C332 VDD2.n124 B 0.020607f
C333 VDD2.n125 B 0.016231f
C334 VDD2.n126 B 0.011625f
C335 VDD2.n127 B 1.57603f
C336 VDD2.n128 B 0.021633f
C337 VDD2.n129 B 0.011625f
C338 VDD2.n130 B 0.012309f
C339 VDD2.n131 B 0.027477f
C340 VDD2.n132 B 0.027477f
C341 VDD2.n133 B 0.012309f
C342 VDD2.n134 B 0.011625f
C343 VDD2.n135 B 0.021633f
C344 VDD2.n136 B 0.021633f
C345 VDD2.n137 B 0.011625f
C346 VDD2.n138 B 0.012309f
C347 VDD2.n139 B 0.027477f
C348 VDD2.n140 B 0.027477f
C349 VDD2.n141 B 0.012309f
C350 VDD2.n142 B 0.011625f
C351 VDD2.n143 B 0.021633f
C352 VDD2.n144 B 0.021633f
C353 VDD2.n145 B 0.011625f
C354 VDD2.n146 B 0.012309f
C355 VDD2.n147 B 0.027477f
C356 VDD2.n148 B 0.027477f
C357 VDD2.n149 B 0.012309f
C358 VDD2.n150 B 0.011625f
C359 VDD2.n151 B 0.021633f
C360 VDD2.n152 B 0.021633f
C361 VDD2.n153 B 0.011625f
C362 VDD2.n154 B 0.012309f
C363 VDD2.n155 B 0.027477f
C364 VDD2.n156 B 0.027477f
C365 VDD2.n157 B 0.012309f
C366 VDD2.n158 B 0.011625f
C367 VDD2.n159 B 0.021633f
C368 VDD2.n160 B 0.021633f
C369 VDD2.n161 B 0.011625f
C370 VDD2.n162 B 0.012309f
C371 VDD2.n163 B 0.027477f
C372 VDD2.n164 B 0.027477f
C373 VDD2.n165 B 0.012309f
C374 VDD2.n166 B 0.011625f
C375 VDD2.n167 B 0.021633f
C376 VDD2.n168 B 0.021633f
C377 VDD2.n169 B 0.011625f
C378 VDD2.n170 B 0.011967f
C379 VDD2.n171 B 0.011967f
C380 VDD2.n172 B 0.027477f
C381 VDD2.n173 B 0.027477f
C382 VDD2.n174 B 0.012309f
C383 VDD2.n175 B 0.011625f
C384 VDD2.n176 B 0.021633f
C385 VDD2.n177 B 0.021633f
C386 VDD2.n178 B 0.011625f
C387 VDD2.n179 B 0.012309f
C388 VDD2.n180 B 0.027477f
C389 VDD2.n181 B 0.054836f
C390 VDD2.n182 B 0.012309f
C391 VDD2.n183 B 0.011625f
C392 VDD2.n184 B 0.047049f
C393 VDD2.n185 B 0.045075f
C394 VDD2.n186 B 2.69299f
C395 VTAIL.n0 B 0.022581f
C396 VTAIL.n1 B 0.017584f
C397 VTAIL.n2 B 0.009449f
C398 VTAIL.n3 B 0.022334f
C399 VTAIL.n4 B 0.010005f
C400 VTAIL.n5 B 0.017584f
C401 VTAIL.n6 B 0.009449f
C402 VTAIL.n7 B 0.022334f
C403 VTAIL.n8 B 0.010005f
C404 VTAIL.n9 B 0.017584f
C405 VTAIL.n10 B 0.009449f
C406 VTAIL.n11 B 0.022334f
C407 VTAIL.n12 B 0.010005f
C408 VTAIL.n13 B 0.017584f
C409 VTAIL.n14 B 0.009449f
C410 VTAIL.n15 B 0.022334f
C411 VTAIL.n16 B 0.010005f
C412 VTAIL.n17 B 0.017584f
C413 VTAIL.n18 B 0.009449f
C414 VTAIL.n19 B 0.022334f
C415 VTAIL.n20 B 0.010005f
C416 VTAIL.n21 B 0.017584f
C417 VTAIL.n22 B 0.009449f
C418 VTAIL.n23 B 0.022334f
C419 VTAIL.n24 B 0.010005f
C420 VTAIL.n25 B 0.017584f
C421 VTAIL.n26 B 0.009449f
C422 VTAIL.n27 B 0.022334f
C423 VTAIL.n28 B 0.010005f
C424 VTAIL.n29 B 0.122182f
C425 VTAIL.t0 B 0.036928f
C426 VTAIL.n30 B 0.01675f
C427 VTAIL.n31 B 0.013193f
C428 VTAIL.n32 B 0.009449f
C429 VTAIL.n33 B 1.28105f
C430 VTAIL.n34 B 0.017584f
C431 VTAIL.n35 B 0.009449f
C432 VTAIL.n36 B 0.010005f
C433 VTAIL.n37 B 0.022334f
C434 VTAIL.n38 B 0.022334f
C435 VTAIL.n39 B 0.010005f
C436 VTAIL.n40 B 0.009449f
C437 VTAIL.n41 B 0.017584f
C438 VTAIL.n42 B 0.017584f
C439 VTAIL.n43 B 0.009449f
C440 VTAIL.n44 B 0.010005f
C441 VTAIL.n45 B 0.022334f
C442 VTAIL.n46 B 0.022334f
C443 VTAIL.n47 B 0.010005f
C444 VTAIL.n48 B 0.009449f
C445 VTAIL.n49 B 0.017584f
C446 VTAIL.n50 B 0.017584f
C447 VTAIL.n51 B 0.009449f
C448 VTAIL.n52 B 0.010005f
C449 VTAIL.n53 B 0.022334f
C450 VTAIL.n54 B 0.022334f
C451 VTAIL.n55 B 0.010005f
C452 VTAIL.n56 B 0.009449f
C453 VTAIL.n57 B 0.017584f
C454 VTAIL.n58 B 0.017584f
C455 VTAIL.n59 B 0.009449f
C456 VTAIL.n60 B 0.010005f
C457 VTAIL.n61 B 0.022334f
C458 VTAIL.n62 B 0.022334f
C459 VTAIL.n63 B 0.010005f
C460 VTAIL.n64 B 0.009449f
C461 VTAIL.n65 B 0.017584f
C462 VTAIL.n66 B 0.017584f
C463 VTAIL.n67 B 0.009449f
C464 VTAIL.n68 B 0.010005f
C465 VTAIL.n69 B 0.022334f
C466 VTAIL.n70 B 0.022334f
C467 VTAIL.n71 B 0.022334f
C468 VTAIL.n72 B 0.010005f
C469 VTAIL.n73 B 0.009449f
C470 VTAIL.n74 B 0.017584f
C471 VTAIL.n75 B 0.017584f
C472 VTAIL.n76 B 0.009449f
C473 VTAIL.n77 B 0.009727f
C474 VTAIL.n78 B 0.009727f
C475 VTAIL.n79 B 0.022334f
C476 VTAIL.n80 B 0.022334f
C477 VTAIL.n81 B 0.010005f
C478 VTAIL.n82 B 0.009449f
C479 VTAIL.n83 B 0.017584f
C480 VTAIL.n84 B 0.017584f
C481 VTAIL.n85 B 0.009449f
C482 VTAIL.n86 B 0.010005f
C483 VTAIL.n87 B 0.022334f
C484 VTAIL.n88 B 0.044573f
C485 VTAIL.n89 B 0.010005f
C486 VTAIL.n90 B 0.009449f
C487 VTAIL.n91 B 0.038243f
C488 VTAIL.n92 B 0.024476f
C489 VTAIL.n93 B 1.19034f
C490 VTAIL.n94 B 0.022581f
C491 VTAIL.n95 B 0.017584f
C492 VTAIL.n96 B 0.009449f
C493 VTAIL.n97 B 0.022334f
C494 VTAIL.n98 B 0.010005f
C495 VTAIL.n99 B 0.017584f
C496 VTAIL.n100 B 0.009449f
C497 VTAIL.n101 B 0.022334f
C498 VTAIL.n102 B 0.010005f
C499 VTAIL.n103 B 0.017584f
C500 VTAIL.n104 B 0.009449f
C501 VTAIL.n105 B 0.022334f
C502 VTAIL.n106 B 0.022334f
C503 VTAIL.n107 B 0.010005f
C504 VTAIL.n108 B 0.017584f
C505 VTAIL.n109 B 0.009449f
C506 VTAIL.n110 B 0.022334f
C507 VTAIL.n111 B 0.010005f
C508 VTAIL.n112 B 0.017584f
C509 VTAIL.n113 B 0.009449f
C510 VTAIL.n114 B 0.022334f
C511 VTAIL.n115 B 0.010005f
C512 VTAIL.n116 B 0.017584f
C513 VTAIL.n117 B 0.009449f
C514 VTAIL.n118 B 0.022334f
C515 VTAIL.n119 B 0.010005f
C516 VTAIL.n120 B 0.017584f
C517 VTAIL.n121 B 0.009449f
C518 VTAIL.n122 B 0.022334f
C519 VTAIL.n123 B 0.010005f
C520 VTAIL.n124 B 0.122182f
C521 VTAIL.t1 B 0.036928f
C522 VTAIL.n125 B 0.01675f
C523 VTAIL.n126 B 0.013193f
C524 VTAIL.n127 B 0.009449f
C525 VTAIL.n128 B 1.28105f
C526 VTAIL.n129 B 0.017584f
C527 VTAIL.n130 B 0.009449f
C528 VTAIL.n131 B 0.010005f
C529 VTAIL.n132 B 0.022334f
C530 VTAIL.n133 B 0.022334f
C531 VTAIL.n134 B 0.010005f
C532 VTAIL.n135 B 0.009449f
C533 VTAIL.n136 B 0.017584f
C534 VTAIL.n137 B 0.017584f
C535 VTAIL.n138 B 0.009449f
C536 VTAIL.n139 B 0.010005f
C537 VTAIL.n140 B 0.022334f
C538 VTAIL.n141 B 0.022334f
C539 VTAIL.n142 B 0.010005f
C540 VTAIL.n143 B 0.009449f
C541 VTAIL.n144 B 0.017584f
C542 VTAIL.n145 B 0.017584f
C543 VTAIL.n146 B 0.009449f
C544 VTAIL.n147 B 0.010005f
C545 VTAIL.n148 B 0.022334f
C546 VTAIL.n149 B 0.022334f
C547 VTAIL.n150 B 0.010005f
C548 VTAIL.n151 B 0.009449f
C549 VTAIL.n152 B 0.017584f
C550 VTAIL.n153 B 0.017584f
C551 VTAIL.n154 B 0.009449f
C552 VTAIL.n155 B 0.010005f
C553 VTAIL.n156 B 0.022334f
C554 VTAIL.n157 B 0.022334f
C555 VTAIL.n158 B 0.010005f
C556 VTAIL.n159 B 0.009449f
C557 VTAIL.n160 B 0.017584f
C558 VTAIL.n161 B 0.017584f
C559 VTAIL.n162 B 0.009449f
C560 VTAIL.n163 B 0.010005f
C561 VTAIL.n164 B 0.022334f
C562 VTAIL.n165 B 0.022334f
C563 VTAIL.n166 B 0.010005f
C564 VTAIL.n167 B 0.009449f
C565 VTAIL.n168 B 0.017584f
C566 VTAIL.n169 B 0.017584f
C567 VTAIL.n170 B 0.009449f
C568 VTAIL.n171 B 0.009727f
C569 VTAIL.n172 B 0.009727f
C570 VTAIL.n173 B 0.022334f
C571 VTAIL.n174 B 0.022334f
C572 VTAIL.n175 B 0.010005f
C573 VTAIL.n176 B 0.009449f
C574 VTAIL.n177 B 0.017584f
C575 VTAIL.n178 B 0.017584f
C576 VTAIL.n179 B 0.009449f
C577 VTAIL.n180 B 0.010005f
C578 VTAIL.n181 B 0.022334f
C579 VTAIL.n182 B 0.044573f
C580 VTAIL.n183 B 0.010005f
C581 VTAIL.n184 B 0.009449f
C582 VTAIL.n185 B 0.038243f
C583 VTAIL.n186 B 0.024476f
C584 VTAIL.n187 B 1.19718f
C585 VTAIL.n188 B 0.022581f
C586 VTAIL.n189 B 0.017584f
C587 VTAIL.n190 B 0.009449f
C588 VTAIL.n191 B 0.022334f
C589 VTAIL.n192 B 0.010005f
C590 VTAIL.n193 B 0.017584f
C591 VTAIL.n194 B 0.009449f
C592 VTAIL.n195 B 0.022334f
C593 VTAIL.n196 B 0.010005f
C594 VTAIL.n197 B 0.017584f
C595 VTAIL.n198 B 0.009449f
C596 VTAIL.n199 B 0.022334f
C597 VTAIL.n200 B 0.022334f
C598 VTAIL.n201 B 0.010005f
C599 VTAIL.n202 B 0.017584f
C600 VTAIL.n203 B 0.009449f
C601 VTAIL.n204 B 0.022334f
C602 VTAIL.n205 B 0.010005f
C603 VTAIL.n206 B 0.017584f
C604 VTAIL.n207 B 0.009449f
C605 VTAIL.n208 B 0.022334f
C606 VTAIL.n209 B 0.010005f
C607 VTAIL.n210 B 0.017584f
C608 VTAIL.n211 B 0.009449f
C609 VTAIL.n212 B 0.022334f
C610 VTAIL.n213 B 0.010005f
C611 VTAIL.n214 B 0.017584f
C612 VTAIL.n215 B 0.009449f
C613 VTAIL.n216 B 0.022334f
C614 VTAIL.n217 B 0.010005f
C615 VTAIL.n218 B 0.122182f
C616 VTAIL.t3 B 0.036928f
C617 VTAIL.n219 B 0.01675f
C618 VTAIL.n220 B 0.013193f
C619 VTAIL.n221 B 0.009449f
C620 VTAIL.n222 B 1.28105f
C621 VTAIL.n223 B 0.017584f
C622 VTAIL.n224 B 0.009449f
C623 VTAIL.n225 B 0.010005f
C624 VTAIL.n226 B 0.022334f
C625 VTAIL.n227 B 0.022334f
C626 VTAIL.n228 B 0.010005f
C627 VTAIL.n229 B 0.009449f
C628 VTAIL.n230 B 0.017584f
C629 VTAIL.n231 B 0.017584f
C630 VTAIL.n232 B 0.009449f
C631 VTAIL.n233 B 0.010005f
C632 VTAIL.n234 B 0.022334f
C633 VTAIL.n235 B 0.022334f
C634 VTAIL.n236 B 0.010005f
C635 VTAIL.n237 B 0.009449f
C636 VTAIL.n238 B 0.017584f
C637 VTAIL.n239 B 0.017584f
C638 VTAIL.n240 B 0.009449f
C639 VTAIL.n241 B 0.010005f
C640 VTAIL.n242 B 0.022334f
C641 VTAIL.n243 B 0.022334f
C642 VTAIL.n244 B 0.010005f
C643 VTAIL.n245 B 0.009449f
C644 VTAIL.n246 B 0.017584f
C645 VTAIL.n247 B 0.017584f
C646 VTAIL.n248 B 0.009449f
C647 VTAIL.n249 B 0.010005f
C648 VTAIL.n250 B 0.022334f
C649 VTAIL.n251 B 0.022334f
C650 VTAIL.n252 B 0.010005f
C651 VTAIL.n253 B 0.009449f
C652 VTAIL.n254 B 0.017584f
C653 VTAIL.n255 B 0.017584f
C654 VTAIL.n256 B 0.009449f
C655 VTAIL.n257 B 0.010005f
C656 VTAIL.n258 B 0.022334f
C657 VTAIL.n259 B 0.022334f
C658 VTAIL.n260 B 0.010005f
C659 VTAIL.n261 B 0.009449f
C660 VTAIL.n262 B 0.017584f
C661 VTAIL.n263 B 0.017584f
C662 VTAIL.n264 B 0.009449f
C663 VTAIL.n265 B 0.009727f
C664 VTAIL.n266 B 0.009727f
C665 VTAIL.n267 B 0.022334f
C666 VTAIL.n268 B 0.022334f
C667 VTAIL.n269 B 0.010005f
C668 VTAIL.n270 B 0.009449f
C669 VTAIL.n271 B 0.017584f
C670 VTAIL.n272 B 0.017584f
C671 VTAIL.n273 B 0.009449f
C672 VTAIL.n274 B 0.010005f
C673 VTAIL.n275 B 0.022334f
C674 VTAIL.n276 B 0.044573f
C675 VTAIL.n277 B 0.010005f
C676 VTAIL.n278 B 0.009449f
C677 VTAIL.n279 B 0.038243f
C678 VTAIL.n280 B 0.024476f
C679 VTAIL.n281 B 1.15664f
C680 VTAIL.n282 B 0.022581f
C681 VTAIL.n283 B 0.017584f
C682 VTAIL.n284 B 0.009449f
C683 VTAIL.n285 B 0.022334f
C684 VTAIL.n286 B 0.010005f
C685 VTAIL.n287 B 0.017584f
C686 VTAIL.n288 B 0.009449f
C687 VTAIL.n289 B 0.022334f
C688 VTAIL.n290 B 0.010005f
C689 VTAIL.n291 B 0.017584f
C690 VTAIL.n292 B 0.009449f
C691 VTAIL.n293 B 0.022334f
C692 VTAIL.n294 B 0.010005f
C693 VTAIL.n295 B 0.017584f
C694 VTAIL.n296 B 0.009449f
C695 VTAIL.n297 B 0.022334f
C696 VTAIL.n298 B 0.010005f
C697 VTAIL.n299 B 0.017584f
C698 VTAIL.n300 B 0.009449f
C699 VTAIL.n301 B 0.022334f
C700 VTAIL.n302 B 0.010005f
C701 VTAIL.n303 B 0.017584f
C702 VTAIL.n304 B 0.009449f
C703 VTAIL.n305 B 0.022334f
C704 VTAIL.n306 B 0.010005f
C705 VTAIL.n307 B 0.017584f
C706 VTAIL.n308 B 0.009449f
C707 VTAIL.n309 B 0.022334f
C708 VTAIL.n310 B 0.010005f
C709 VTAIL.n311 B 0.122182f
C710 VTAIL.t2 B 0.036928f
C711 VTAIL.n312 B 0.01675f
C712 VTAIL.n313 B 0.013193f
C713 VTAIL.n314 B 0.009449f
C714 VTAIL.n315 B 1.28105f
C715 VTAIL.n316 B 0.017584f
C716 VTAIL.n317 B 0.009449f
C717 VTAIL.n318 B 0.010005f
C718 VTAIL.n319 B 0.022334f
C719 VTAIL.n320 B 0.022334f
C720 VTAIL.n321 B 0.010005f
C721 VTAIL.n322 B 0.009449f
C722 VTAIL.n323 B 0.017584f
C723 VTAIL.n324 B 0.017584f
C724 VTAIL.n325 B 0.009449f
C725 VTAIL.n326 B 0.010005f
C726 VTAIL.n327 B 0.022334f
C727 VTAIL.n328 B 0.022334f
C728 VTAIL.n329 B 0.010005f
C729 VTAIL.n330 B 0.009449f
C730 VTAIL.n331 B 0.017584f
C731 VTAIL.n332 B 0.017584f
C732 VTAIL.n333 B 0.009449f
C733 VTAIL.n334 B 0.010005f
C734 VTAIL.n335 B 0.022334f
C735 VTAIL.n336 B 0.022334f
C736 VTAIL.n337 B 0.010005f
C737 VTAIL.n338 B 0.009449f
C738 VTAIL.n339 B 0.017584f
C739 VTAIL.n340 B 0.017584f
C740 VTAIL.n341 B 0.009449f
C741 VTAIL.n342 B 0.010005f
C742 VTAIL.n343 B 0.022334f
C743 VTAIL.n344 B 0.022334f
C744 VTAIL.n345 B 0.010005f
C745 VTAIL.n346 B 0.009449f
C746 VTAIL.n347 B 0.017584f
C747 VTAIL.n348 B 0.017584f
C748 VTAIL.n349 B 0.009449f
C749 VTAIL.n350 B 0.010005f
C750 VTAIL.n351 B 0.022334f
C751 VTAIL.n352 B 0.022334f
C752 VTAIL.n353 B 0.022334f
C753 VTAIL.n354 B 0.010005f
C754 VTAIL.n355 B 0.009449f
C755 VTAIL.n356 B 0.017584f
C756 VTAIL.n357 B 0.017584f
C757 VTAIL.n358 B 0.009449f
C758 VTAIL.n359 B 0.009727f
C759 VTAIL.n360 B 0.009727f
C760 VTAIL.n361 B 0.022334f
C761 VTAIL.n362 B 0.022334f
C762 VTAIL.n363 B 0.010005f
C763 VTAIL.n364 B 0.009449f
C764 VTAIL.n365 B 0.017584f
C765 VTAIL.n366 B 0.017584f
C766 VTAIL.n367 B 0.009449f
C767 VTAIL.n368 B 0.010005f
C768 VTAIL.n369 B 0.022334f
C769 VTAIL.n370 B 0.044573f
C770 VTAIL.n371 B 0.010005f
C771 VTAIL.n372 B 0.009449f
C772 VTAIL.n373 B 0.038243f
C773 VTAIL.n374 B 0.024476f
C774 VTAIL.n375 B 1.11659f
C775 VN.t1 B 1.25217f
C776 VN.t0 B 1.35202f
.ends

