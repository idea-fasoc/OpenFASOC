* NGSPICE file created from diff_pair_sample_1452.ext - technology: sky130A

.subckt diff_pair_sample_1452 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n3450_n4312# sky130_fd_pr__pfet_01v8 ad=6.5208 pd=34.22 as=0 ps=0 w=16.72 l=2.77
X1 VTAIL.t10 VP.t0 VDD1.t4 w_n3450_n4312# sky130_fd_pr__pfet_01v8 ad=2.7588 pd=17.05 as=2.7588 ps=17.05 w=16.72 l=2.77
X2 VTAIL.t9 VP.t1 VDD1.t3 w_n3450_n4312# sky130_fd_pr__pfet_01v8 ad=2.7588 pd=17.05 as=2.7588 ps=17.05 w=16.72 l=2.77
X3 VTAIL.t3 VN.t0 VDD2.t5 w_n3450_n4312# sky130_fd_pr__pfet_01v8 ad=2.7588 pd=17.05 as=2.7588 ps=17.05 w=16.72 l=2.77
X4 B.t8 B.t6 B.t7 w_n3450_n4312# sky130_fd_pr__pfet_01v8 ad=6.5208 pd=34.22 as=0 ps=0 w=16.72 l=2.77
X5 VDD1.t5 VP.t2 VTAIL.t8 w_n3450_n4312# sky130_fd_pr__pfet_01v8 ad=2.7588 pd=17.05 as=6.5208 ps=34.22 w=16.72 l=2.77
X6 VDD1.t1 VP.t3 VTAIL.t7 w_n3450_n4312# sky130_fd_pr__pfet_01v8 ad=6.5208 pd=34.22 as=2.7588 ps=17.05 w=16.72 l=2.77
X7 VDD2.t4 VN.t1 VTAIL.t1 w_n3450_n4312# sky130_fd_pr__pfet_01v8 ad=2.7588 pd=17.05 as=6.5208 ps=34.22 w=16.72 l=2.77
X8 VDD2.t3 VN.t2 VTAIL.t2 w_n3450_n4312# sky130_fd_pr__pfet_01v8 ad=6.5208 pd=34.22 as=2.7588 ps=17.05 w=16.72 l=2.77
X9 B.t5 B.t3 B.t4 w_n3450_n4312# sky130_fd_pr__pfet_01v8 ad=6.5208 pd=34.22 as=0 ps=0 w=16.72 l=2.77
X10 B.t2 B.t0 B.t1 w_n3450_n4312# sky130_fd_pr__pfet_01v8 ad=6.5208 pd=34.22 as=0 ps=0 w=16.72 l=2.77
X11 VDD2.t2 VN.t3 VTAIL.t11 w_n3450_n4312# sky130_fd_pr__pfet_01v8 ad=2.7588 pd=17.05 as=6.5208 ps=34.22 w=16.72 l=2.77
X12 VDD1.t2 VP.t4 VTAIL.t6 w_n3450_n4312# sky130_fd_pr__pfet_01v8 ad=2.7588 pd=17.05 as=6.5208 ps=34.22 w=16.72 l=2.77
X13 VTAIL.t4 VN.t4 VDD2.t1 w_n3450_n4312# sky130_fd_pr__pfet_01v8 ad=2.7588 pd=17.05 as=2.7588 ps=17.05 w=16.72 l=2.77
X14 VDD1.t0 VP.t5 VTAIL.t5 w_n3450_n4312# sky130_fd_pr__pfet_01v8 ad=6.5208 pd=34.22 as=2.7588 ps=17.05 w=16.72 l=2.77
X15 VDD2.t0 VN.t5 VTAIL.t0 w_n3450_n4312# sky130_fd_pr__pfet_01v8 ad=6.5208 pd=34.22 as=2.7588 ps=17.05 w=16.72 l=2.77
R0 B.n467 B.n134 585
R1 B.n466 B.n465 585
R2 B.n464 B.n135 585
R3 B.n463 B.n462 585
R4 B.n461 B.n136 585
R5 B.n460 B.n459 585
R6 B.n458 B.n137 585
R7 B.n457 B.n456 585
R8 B.n455 B.n138 585
R9 B.n454 B.n453 585
R10 B.n452 B.n139 585
R11 B.n451 B.n450 585
R12 B.n449 B.n140 585
R13 B.n448 B.n447 585
R14 B.n446 B.n141 585
R15 B.n445 B.n444 585
R16 B.n443 B.n142 585
R17 B.n442 B.n441 585
R18 B.n440 B.n143 585
R19 B.n439 B.n438 585
R20 B.n437 B.n144 585
R21 B.n436 B.n435 585
R22 B.n434 B.n145 585
R23 B.n433 B.n432 585
R24 B.n431 B.n146 585
R25 B.n430 B.n429 585
R26 B.n428 B.n147 585
R27 B.n427 B.n426 585
R28 B.n425 B.n148 585
R29 B.n424 B.n423 585
R30 B.n422 B.n149 585
R31 B.n421 B.n420 585
R32 B.n419 B.n150 585
R33 B.n418 B.n417 585
R34 B.n416 B.n151 585
R35 B.n415 B.n414 585
R36 B.n413 B.n152 585
R37 B.n412 B.n411 585
R38 B.n410 B.n153 585
R39 B.n409 B.n408 585
R40 B.n407 B.n154 585
R41 B.n406 B.n405 585
R42 B.n404 B.n155 585
R43 B.n403 B.n402 585
R44 B.n401 B.n156 585
R45 B.n400 B.n399 585
R46 B.n398 B.n157 585
R47 B.n397 B.n396 585
R48 B.n395 B.n158 585
R49 B.n394 B.n393 585
R50 B.n392 B.n159 585
R51 B.n391 B.n390 585
R52 B.n389 B.n160 585
R53 B.n388 B.n387 585
R54 B.n386 B.n161 585
R55 B.n385 B.n384 585
R56 B.n383 B.n382 585
R57 B.n381 B.n165 585
R58 B.n380 B.n379 585
R59 B.n378 B.n166 585
R60 B.n377 B.n376 585
R61 B.n375 B.n167 585
R62 B.n374 B.n373 585
R63 B.n372 B.n168 585
R64 B.n371 B.n370 585
R65 B.n368 B.n169 585
R66 B.n367 B.n366 585
R67 B.n365 B.n172 585
R68 B.n364 B.n363 585
R69 B.n362 B.n173 585
R70 B.n361 B.n360 585
R71 B.n359 B.n174 585
R72 B.n358 B.n357 585
R73 B.n356 B.n175 585
R74 B.n355 B.n354 585
R75 B.n353 B.n176 585
R76 B.n352 B.n351 585
R77 B.n350 B.n177 585
R78 B.n349 B.n348 585
R79 B.n347 B.n178 585
R80 B.n346 B.n345 585
R81 B.n344 B.n179 585
R82 B.n343 B.n342 585
R83 B.n341 B.n180 585
R84 B.n340 B.n339 585
R85 B.n338 B.n181 585
R86 B.n337 B.n336 585
R87 B.n335 B.n182 585
R88 B.n334 B.n333 585
R89 B.n332 B.n183 585
R90 B.n331 B.n330 585
R91 B.n329 B.n184 585
R92 B.n328 B.n327 585
R93 B.n326 B.n185 585
R94 B.n325 B.n324 585
R95 B.n323 B.n186 585
R96 B.n322 B.n321 585
R97 B.n320 B.n187 585
R98 B.n319 B.n318 585
R99 B.n317 B.n188 585
R100 B.n316 B.n315 585
R101 B.n314 B.n189 585
R102 B.n313 B.n312 585
R103 B.n311 B.n190 585
R104 B.n310 B.n309 585
R105 B.n308 B.n191 585
R106 B.n307 B.n306 585
R107 B.n305 B.n192 585
R108 B.n304 B.n303 585
R109 B.n302 B.n193 585
R110 B.n301 B.n300 585
R111 B.n299 B.n194 585
R112 B.n298 B.n297 585
R113 B.n296 B.n195 585
R114 B.n295 B.n294 585
R115 B.n293 B.n196 585
R116 B.n292 B.n291 585
R117 B.n290 B.n197 585
R118 B.n289 B.n288 585
R119 B.n287 B.n198 585
R120 B.n286 B.n285 585
R121 B.n469 B.n468 585
R122 B.n470 B.n133 585
R123 B.n472 B.n471 585
R124 B.n473 B.n132 585
R125 B.n475 B.n474 585
R126 B.n476 B.n131 585
R127 B.n478 B.n477 585
R128 B.n479 B.n130 585
R129 B.n481 B.n480 585
R130 B.n482 B.n129 585
R131 B.n484 B.n483 585
R132 B.n485 B.n128 585
R133 B.n487 B.n486 585
R134 B.n488 B.n127 585
R135 B.n490 B.n489 585
R136 B.n491 B.n126 585
R137 B.n493 B.n492 585
R138 B.n494 B.n125 585
R139 B.n496 B.n495 585
R140 B.n497 B.n124 585
R141 B.n499 B.n498 585
R142 B.n500 B.n123 585
R143 B.n502 B.n501 585
R144 B.n503 B.n122 585
R145 B.n505 B.n504 585
R146 B.n506 B.n121 585
R147 B.n508 B.n507 585
R148 B.n509 B.n120 585
R149 B.n511 B.n510 585
R150 B.n512 B.n119 585
R151 B.n514 B.n513 585
R152 B.n515 B.n118 585
R153 B.n517 B.n516 585
R154 B.n518 B.n117 585
R155 B.n520 B.n519 585
R156 B.n521 B.n116 585
R157 B.n523 B.n522 585
R158 B.n524 B.n115 585
R159 B.n526 B.n525 585
R160 B.n527 B.n114 585
R161 B.n529 B.n528 585
R162 B.n530 B.n113 585
R163 B.n532 B.n531 585
R164 B.n533 B.n112 585
R165 B.n535 B.n534 585
R166 B.n536 B.n111 585
R167 B.n538 B.n537 585
R168 B.n539 B.n110 585
R169 B.n541 B.n540 585
R170 B.n542 B.n109 585
R171 B.n544 B.n543 585
R172 B.n545 B.n108 585
R173 B.n547 B.n546 585
R174 B.n548 B.n107 585
R175 B.n550 B.n549 585
R176 B.n551 B.n106 585
R177 B.n553 B.n552 585
R178 B.n554 B.n105 585
R179 B.n556 B.n555 585
R180 B.n557 B.n104 585
R181 B.n559 B.n558 585
R182 B.n560 B.n103 585
R183 B.n562 B.n561 585
R184 B.n563 B.n102 585
R185 B.n565 B.n564 585
R186 B.n566 B.n101 585
R187 B.n568 B.n567 585
R188 B.n569 B.n100 585
R189 B.n571 B.n570 585
R190 B.n572 B.n99 585
R191 B.n574 B.n573 585
R192 B.n575 B.n98 585
R193 B.n577 B.n576 585
R194 B.n578 B.n97 585
R195 B.n580 B.n579 585
R196 B.n581 B.n96 585
R197 B.n583 B.n582 585
R198 B.n584 B.n95 585
R199 B.n586 B.n585 585
R200 B.n587 B.n94 585
R201 B.n589 B.n588 585
R202 B.n590 B.n93 585
R203 B.n592 B.n591 585
R204 B.n593 B.n92 585
R205 B.n595 B.n594 585
R206 B.n596 B.n91 585
R207 B.n598 B.n597 585
R208 B.n599 B.n90 585
R209 B.n601 B.n600 585
R210 B.n602 B.n89 585
R211 B.n785 B.n24 585
R212 B.n784 B.n783 585
R213 B.n782 B.n25 585
R214 B.n781 B.n780 585
R215 B.n779 B.n26 585
R216 B.n778 B.n777 585
R217 B.n776 B.n27 585
R218 B.n775 B.n774 585
R219 B.n773 B.n28 585
R220 B.n772 B.n771 585
R221 B.n770 B.n29 585
R222 B.n769 B.n768 585
R223 B.n767 B.n30 585
R224 B.n766 B.n765 585
R225 B.n764 B.n31 585
R226 B.n763 B.n762 585
R227 B.n761 B.n32 585
R228 B.n760 B.n759 585
R229 B.n758 B.n33 585
R230 B.n757 B.n756 585
R231 B.n755 B.n34 585
R232 B.n754 B.n753 585
R233 B.n752 B.n35 585
R234 B.n751 B.n750 585
R235 B.n749 B.n36 585
R236 B.n748 B.n747 585
R237 B.n746 B.n37 585
R238 B.n745 B.n744 585
R239 B.n743 B.n38 585
R240 B.n742 B.n741 585
R241 B.n740 B.n39 585
R242 B.n739 B.n738 585
R243 B.n737 B.n40 585
R244 B.n736 B.n735 585
R245 B.n734 B.n41 585
R246 B.n733 B.n732 585
R247 B.n731 B.n42 585
R248 B.n730 B.n729 585
R249 B.n728 B.n43 585
R250 B.n727 B.n726 585
R251 B.n725 B.n44 585
R252 B.n724 B.n723 585
R253 B.n722 B.n45 585
R254 B.n721 B.n720 585
R255 B.n719 B.n46 585
R256 B.n718 B.n717 585
R257 B.n716 B.n47 585
R258 B.n715 B.n714 585
R259 B.n713 B.n48 585
R260 B.n712 B.n711 585
R261 B.n710 B.n49 585
R262 B.n709 B.n708 585
R263 B.n707 B.n50 585
R264 B.n706 B.n705 585
R265 B.n704 B.n51 585
R266 B.n703 B.n702 585
R267 B.n701 B.n700 585
R268 B.n699 B.n55 585
R269 B.n698 B.n697 585
R270 B.n696 B.n56 585
R271 B.n695 B.n694 585
R272 B.n693 B.n57 585
R273 B.n692 B.n691 585
R274 B.n690 B.n58 585
R275 B.n689 B.n688 585
R276 B.n686 B.n59 585
R277 B.n685 B.n684 585
R278 B.n683 B.n62 585
R279 B.n682 B.n681 585
R280 B.n680 B.n63 585
R281 B.n679 B.n678 585
R282 B.n677 B.n64 585
R283 B.n676 B.n675 585
R284 B.n674 B.n65 585
R285 B.n673 B.n672 585
R286 B.n671 B.n66 585
R287 B.n670 B.n669 585
R288 B.n668 B.n67 585
R289 B.n667 B.n666 585
R290 B.n665 B.n68 585
R291 B.n664 B.n663 585
R292 B.n662 B.n69 585
R293 B.n661 B.n660 585
R294 B.n659 B.n70 585
R295 B.n658 B.n657 585
R296 B.n656 B.n71 585
R297 B.n655 B.n654 585
R298 B.n653 B.n72 585
R299 B.n652 B.n651 585
R300 B.n650 B.n73 585
R301 B.n649 B.n648 585
R302 B.n647 B.n74 585
R303 B.n646 B.n645 585
R304 B.n644 B.n75 585
R305 B.n643 B.n642 585
R306 B.n641 B.n76 585
R307 B.n640 B.n639 585
R308 B.n638 B.n77 585
R309 B.n637 B.n636 585
R310 B.n635 B.n78 585
R311 B.n634 B.n633 585
R312 B.n632 B.n79 585
R313 B.n631 B.n630 585
R314 B.n629 B.n80 585
R315 B.n628 B.n627 585
R316 B.n626 B.n81 585
R317 B.n625 B.n624 585
R318 B.n623 B.n82 585
R319 B.n622 B.n621 585
R320 B.n620 B.n83 585
R321 B.n619 B.n618 585
R322 B.n617 B.n84 585
R323 B.n616 B.n615 585
R324 B.n614 B.n85 585
R325 B.n613 B.n612 585
R326 B.n611 B.n86 585
R327 B.n610 B.n609 585
R328 B.n608 B.n87 585
R329 B.n607 B.n606 585
R330 B.n605 B.n88 585
R331 B.n604 B.n603 585
R332 B.n787 B.n786 585
R333 B.n788 B.n23 585
R334 B.n790 B.n789 585
R335 B.n791 B.n22 585
R336 B.n793 B.n792 585
R337 B.n794 B.n21 585
R338 B.n796 B.n795 585
R339 B.n797 B.n20 585
R340 B.n799 B.n798 585
R341 B.n800 B.n19 585
R342 B.n802 B.n801 585
R343 B.n803 B.n18 585
R344 B.n805 B.n804 585
R345 B.n806 B.n17 585
R346 B.n808 B.n807 585
R347 B.n809 B.n16 585
R348 B.n811 B.n810 585
R349 B.n812 B.n15 585
R350 B.n814 B.n813 585
R351 B.n815 B.n14 585
R352 B.n817 B.n816 585
R353 B.n818 B.n13 585
R354 B.n820 B.n819 585
R355 B.n821 B.n12 585
R356 B.n823 B.n822 585
R357 B.n824 B.n11 585
R358 B.n826 B.n825 585
R359 B.n827 B.n10 585
R360 B.n829 B.n828 585
R361 B.n830 B.n9 585
R362 B.n832 B.n831 585
R363 B.n833 B.n8 585
R364 B.n835 B.n834 585
R365 B.n836 B.n7 585
R366 B.n838 B.n837 585
R367 B.n839 B.n6 585
R368 B.n841 B.n840 585
R369 B.n842 B.n5 585
R370 B.n844 B.n843 585
R371 B.n845 B.n4 585
R372 B.n847 B.n846 585
R373 B.n848 B.n3 585
R374 B.n850 B.n849 585
R375 B.n851 B.n0 585
R376 B.n2 B.n1 585
R377 B.n221 B.n220 585
R378 B.n223 B.n222 585
R379 B.n224 B.n219 585
R380 B.n226 B.n225 585
R381 B.n227 B.n218 585
R382 B.n229 B.n228 585
R383 B.n230 B.n217 585
R384 B.n232 B.n231 585
R385 B.n233 B.n216 585
R386 B.n235 B.n234 585
R387 B.n236 B.n215 585
R388 B.n238 B.n237 585
R389 B.n239 B.n214 585
R390 B.n241 B.n240 585
R391 B.n242 B.n213 585
R392 B.n244 B.n243 585
R393 B.n245 B.n212 585
R394 B.n247 B.n246 585
R395 B.n248 B.n211 585
R396 B.n250 B.n249 585
R397 B.n251 B.n210 585
R398 B.n253 B.n252 585
R399 B.n254 B.n209 585
R400 B.n256 B.n255 585
R401 B.n257 B.n208 585
R402 B.n259 B.n258 585
R403 B.n260 B.n207 585
R404 B.n262 B.n261 585
R405 B.n263 B.n206 585
R406 B.n265 B.n264 585
R407 B.n266 B.n205 585
R408 B.n268 B.n267 585
R409 B.n269 B.n204 585
R410 B.n271 B.n270 585
R411 B.n272 B.n203 585
R412 B.n274 B.n273 585
R413 B.n275 B.n202 585
R414 B.n277 B.n276 585
R415 B.n278 B.n201 585
R416 B.n280 B.n279 585
R417 B.n281 B.n200 585
R418 B.n283 B.n282 585
R419 B.n284 B.n199 585
R420 B.n162 B.t4 520.611
R421 B.n60 B.t11 520.611
R422 B.n170 B.t1 520.611
R423 B.n52 B.t8 520.611
R424 B.n286 B.n199 478.086
R425 B.n468 B.n467 478.086
R426 B.n604 B.n89 478.086
R427 B.n786 B.n785 478.086
R428 B.n163 B.t5 460.49
R429 B.n61 B.t10 460.49
R430 B.n171 B.t2 460.49
R431 B.n53 B.t7 460.49
R432 B.n170 B.t0 353.76
R433 B.n162 B.t3 353.76
R434 B.n60 B.t9 353.76
R435 B.n52 B.t6 353.76
R436 B.n853 B.n852 256.663
R437 B.n852 B.n851 235.042
R438 B.n852 B.n2 235.042
R439 B.n287 B.n286 163.367
R440 B.n288 B.n287 163.367
R441 B.n288 B.n197 163.367
R442 B.n292 B.n197 163.367
R443 B.n293 B.n292 163.367
R444 B.n294 B.n293 163.367
R445 B.n294 B.n195 163.367
R446 B.n298 B.n195 163.367
R447 B.n299 B.n298 163.367
R448 B.n300 B.n299 163.367
R449 B.n300 B.n193 163.367
R450 B.n304 B.n193 163.367
R451 B.n305 B.n304 163.367
R452 B.n306 B.n305 163.367
R453 B.n306 B.n191 163.367
R454 B.n310 B.n191 163.367
R455 B.n311 B.n310 163.367
R456 B.n312 B.n311 163.367
R457 B.n312 B.n189 163.367
R458 B.n316 B.n189 163.367
R459 B.n317 B.n316 163.367
R460 B.n318 B.n317 163.367
R461 B.n318 B.n187 163.367
R462 B.n322 B.n187 163.367
R463 B.n323 B.n322 163.367
R464 B.n324 B.n323 163.367
R465 B.n324 B.n185 163.367
R466 B.n328 B.n185 163.367
R467 B.n329 B.n328 163.367
R468 B.n330 B.n329 163.367
R469 B.n330 B.n183 163.367
R470 B.n334 B.n183 163.367
R471 B.n335 B.n334 163.367
R472 B.n336 B.n335 163.367
R473 B.n336 B.n181 163.367
R474 B.n340 B.n181 163.367
R475 B.n341 B.n340 163.367
R476 B.n342 B.n341 163.367
R477 B.n342 B.n179 163.367
R478 B.n346 B.n179 163.367
R479 B.n347 B.n346 163.367
R480 B.n348 B.n347 163.367
R481 B.n348 B.n177 163.367
R482 B.n352 B.n177 163.367
R483 B.n353 B.n352 163.367
R484 B.n354 B.n353 163.367
R485 B.n354 B.n175 163.367
R486 B.n358 B.n175 163.367
R487 B.n359 B.n358 163.367
R488 B.n360 B.n359 163.367
R489 B.n360 B.n173 163.367
R490 B.n364 B.n173 163.367
R491 B.n365 B.n364 163.367
R492 B.n366 B.n365 163.367
R493 B.n366 B.n169 163.367
R494 B.n371 B.n169 163.367
R495 B.n372 B.n371 163.367
R496 B.n373 B.n372 163.367
R497 B.n373 B.n167 163.367
R498 B.n377 B.n167 163.367
R499 B.n378 B.n377 163.367
R500 B.n379 B.n378 163.367
R501 B.n379 B.n165 163.367
R502 B.n383 B.n165 163.367
R503 B.n384 B.n383 163.367
R504 B.n384 B.n161 163.367
R505 B.n388 B.n161 163.367
R506 B.n389 B.n388 163.367
R507 B.n390 B.n389 163.367
R508 B.n390 B.n159 163.367
R509 B.n394 B.n159 163.367
R510 B.n395 B.n394 163.367
R511 B.n396 B.n395 163.367
R512 B.n396 B.n157 163.367
R513 B.n400 B.n157 163.367
R514 B.n401 B.n400 163.367
R515 B.n402 B.n401 163.367
R516 B.n402 B.n155 163.367
R517 B.n406 B.n155 163.367
R518 B.n407 B.n406 163.367
R519 B.n408 B.n407 163.367
R520 B.n408 B.n153 163.367
R521 B.n412 B.n153 163.367
R522 B.n413 B.n412 163.367
R523 B.n414 B.n413 163.367
R524 B.n414 B.n151 163.367
R525 B.n418 B.n151 163.367
R526 B.n419 B.n418 163.367
R527 B.n420 B.n419 163.367
R528 B.n420 B.n149 163.367
R529 B.n424 B.n149 163.367
R530 B.n425 B.n424 163.367
R531 B.n426 B.n425 163.367
R532 B.n426 B.n147 163.367
R533 B.n430 B.n147 163.367
R534 B.n431 B.n430 163.367
R535 B.n432 B.n431 163.367
R536 B.n432 B.n145 163.367
R537 B.n436 B.n145 163.367
R538 B.n437 B.n436 163.367
R539 B.n438 B.n437 163.367
R540 B.n438 B.n143 163.367
R541 B.n442 B.n143 163.367
R542 B.n443 B.n442 163.367
R543 B.n444 B.n443 163.367
R544 B.n444 B.n141 163.367
R545 B.n448 B.n141 163.367
R546 B.n449 B.n448 163.367
R547 B.n450 B.n449 163.367
R548 B.n450 B.n139 163.367
R549 B.n454 B.n139 163.367
R550 B.n455 B.n454 163.367
R551 B.n456 B.n455 163.367
R552 B.n456 B.n137 163.367
R553 B.n460 B.n137 163.367
R554 B.n461 B.n460 163.367
R555 B.n462 B.n461 163.367
R556 B.n462 B.n135 163.367
R557 B.n466 B.n135 163.367
R558 B.n467 B.n466 163.367
R559 B.n600 B.n89 163.367
R560 B.n600 B.n599 163.367
R561 B.n599 B.n598 163.367
R562 B.n598 B.n91 163.367
R563 B.n594 B.n91 163.367
R564 B.n594 B.n593 163.367
R565 B.n593 B.n592 163.367
R566 B.n592 B.n93 163.367
R567 B.n588 B.n93 163.367
R568 B.n588 B.n587 163.367
R569 B.n587 B.n586 163.367
R570 B.n586 B.n95 163.367
R571 B.n582 B.n95 163.367
R572 B.n582 B.n581 163.367
R573 B.n581 B.n580 163.367
R574 B.n580 B.n97 163.367
R575 B.n576 B.n97 163.367
R576 B.n576 B.n575 163.367
R577 B.n575 B.n574 163.367
R578 B.n574 B.n99 163.367
R579 B.n570 B.n99 163.367
R580 B.n570 B.n569 163.367
R581 B.n569 B.n568 163.367
R582 B.n568 B.n101 163.367
R583 B.n564 B.n101 163.367
R584 B.n564 B.n563 163.367
R585 B.n563 B.n562 163.367
R586 B.n562 B.n103 163.367
R587 B.n558 B.n103 163.367
R588 B.n558 B.n557 163.367
R589 B.n557 B.n556 163.367
R590 B.n556 B.n105 163.367
R591 B.n552 B.n105 163.367
R592 B.n552 B.n551 163.367
R593 B.n551 B.n550 163.367
R594 B.n550 B.n107 163.367
R595 B.n546 B.n107 163.367
R596 B.n546 B.n545 163.367
R597 B.n545 B.n544 163.367
R598 B.n544 B.n109 163.367
R599 B.n540 B.n109 163.367
R600 B.n540 B.n539 163.367
R601 B.n539 B.n538 163.367
R602 B.n538 B.n111 163.367
R603 B.n534 B.n111 163.367
R604 B.n534 B.n533 163.367
R605 B.n533 B.n532 163.367
R606 B.n532 B.n113 163.367
R607 B.n528 B.n113 163.367
R608 B.n528 B.n527 163.367
R609 B.n527 B.n526 163.367
R610 B.n526 B.n115 163.367
R611 B.n522 B.n115 163.367
R612 B.n522 B.n521 163.367
R613 B.n521 B.n520 163.367
R614 B.n520 B.n117 163.367
R615 B.n516 B.n117 163.367
R616 B.n516 B.n515 163.367
R617 B.n515 B.n514 163.367
R618 B.n514 B.n119 163.367
R619 B.n510 B.n119 163.367
R620 B.n510 B.n509 163.367
R621 B.n509 B.n508 163.367
R622 B.n508 B.n121 163.367
R623 B.n504 B.n121 163.367
R624 B.n504 B.n503 163.367
R625 B.n503 B.n502 163.367
R626 B.n502 B.n123 163.367
R627 B.n498 B.n123 163.367
R628 B.n498 B.n497 163.367
R629 B.n497 B.n496 163.367
R630 B.n496 B.n125 163.367
R631 B.n492 B.n125 163.367
R632 B.n492 B.n491 163.367
R633 B.n491 B.n490 163.367
R634 B.n490 B.n127 163.367
R635 B.n486 B.n127 163.367
R636 B.n486 B.n485 163.367
R637 B.n485 B.n484 163.367
R638 B.n484 B.n129 163.367
R639 B.n480 B.n129 163.367
R640 B.n480 B.n479 163.367
R641 B.n479 B.n478 163.367
R642 B.n478 B.n131 163.367
R643 B.n474 B.n131 163.367
R644 B.n474 B.n473 163.367
R645 B.n473 B.n472 163.367
R646 B.n472 B.n133 163.367
R647 B.n468 B.n133 163.367
R648 B.n785 B.n784 163.367
R649 B.n784 B.n25 163.367
R650 B.n780 B.n25 163.367
R651 B.n780 B.n779 163.367
R652 B.n779 B.n778 163.367
R653 B.n778 B.n27 163.367
R654 B.n774 B.n27 163.367
R655 B.n774 B.n773 163.367
R656 B.n773 B.n772 163.367
R657 B.n772 B.n29 163.367
R658 B.n768 B.n29 163.367
R659 B.n768 B.n767 163.367
R660 B.n767 B.n766 163.367
R661 B.n766 B.n31 163.367
R662 B.n762 B.n31 163.367
R663 B.n762 B.n761 163.367
R664 B.n761 B.n760 163.367
R665 B.n760 B.n33 163.367
R666 B.n756 B.n33 163.367
R667 B.n756 B.n755 163.367
R668 B.n755 B.n754 163.367
R669 B.n754 B.n35 163.367
R670 B.n750 B.n35 163.367
R671 B.n750 B.n749 163.367
R672 B.n749 B.n748 163.367
R673 B.n748 B.n37 163.367
R674 B.n744 B.n37 163.367
R675 B.n744 B.n743 163.367
R676 B.n743 B.n742 163.367
R677 B.n742 B.n39 163.367
R678 B.n738 B.n39 163.367
R679 B.n738 B.n737 163.367
R680 B.n737 B.n736 163.367
R681 B.n736 B.n41 163.367
R682 B.n732 B.n41 163.367
R683 B.n732 B.n731 163.367
R684 B.n731 B.n730 163.367
R685 B.n730 B.n43 163.367
R686 B.n726 B.n43 163.367
R687 B.n726 B.n725 163.367
R688 B.n725 B.n724 163.367
R689 B.n724 B.n45 163.367
R690 B.n720 B.n45 163.367
R691 B.n720 B.n719 163.367
R692 B.n719 B.n718 163.367
R693 B.n718 B.n47 163.367
R694 B.n714 B.n47 163.367
R695 B.n714 B.n713 163.367
R696 B.n713 B.n712 163.367
R697 B.n712 B.n49 163.367
R698 B.n708 B.n49 163.367
R699 B.n708 B.n707 163.367
R700 B.n707 B.n706 163.367
R701 B.n706 B.n51 163.367
R702 B.n702 B.n51 163.367
R703 B.n702 B.n701 163.367
R704 B.n701 B.n55 163.367
R705 B.n697 B.n55 163.367
R706 B.n697 B.n696 163.367
R707 B.n696 B.n695 163.367
R708 B.n695 B.n57 163.367
R709 B.n691 B.n57 163.367
R710 B.n691 B.n690 163.367
R711 B.n690 B.n689 163.367
R712 B.n689 B.n59 163.367
R713 B.n684 B.n59 163.367
R714 B.n684 B.n683 163.367
R715 B.n683 B.n682 163.367
R716 B.n682 B.n63 163.367
R717 B.n678 B.n63 163.367
R718 B.n678 B.n677 163.367
R719 B.n677 B.n676 163.367
R720 B.n676 B.n65 163.367
R721 B.n672 B.n65 163.367
R722 B.n672 B.n671 163.367
R723 B.n671 B.n670 163.367
R724 B.n670 B.n67 163.367
R725 B.n666 B.n67 163.367
R726 B.n666 B.n665 163.367
R727 B.n665 B.n664 163.367
R728 B.n664 B.n69 163.367
R729 B.n660 B.n69 163.367
R730 B.n660 B.n659 163.367
R731 B.n659 B.n658 163.367
R732 B.n658 B.n71 163.367
R733 B.n654 B.n71 163.367
R734 B.n654 B.n653 163.367
R735 B.n653 B.n652 163.367
R736 B.n652 B.n73 163.367
R737 B.n648 B.n73 163.367
R738 B.n648 B.n647 163.367
R739 B.n647 B.n646 163.367
R740 B.n646 B.n75 163.367
R741 B.n642 B.n75 163.367
R742 B.n642 B.n641 163.367
R743 B.n641 B.n640 163.367
R744 B.n640 B.n77 163.367
R745 B.n636 B.n77 163.367
R746 B.n636 B.n635 163.367
R747 B.n635 B.n634 163.367
R748 B.n634 B.n79 163.367
R749 B.n630 B.n79 163.367
R750 B.n630 B.n629 163.367
R751 B.n629 B.n628 163.367
R752 B.n628 B.n81 163.367
R753 B.n624 B.n81 163.367
R754 B.n624 B.n623 163.367
R755 B.n623 B.n622 163.367
R756 B.n622 B.n83 163.367
R757 B.n618 B.n83 163.367
R758 B.n618 B.n617 163.367
R759 B.n617 B.n616 163.367
R760 B.n616 B.n85 163.367
R761 B.n612 B.n85 163.367
R762 B.n612 B.n611 163.367
R763 B.n611 B.n610 163.367
R764 B.n610 B.n87 163.367
R765 B.n606 B.n87 163.367
R766 B.n606 B.n605 163.367
R767 B.n605 B.n604 163.367
R768 B.n786 B.n23 163.367
R769 B.n790 B.n23 163.367
R770 B.n791 B.n790 163.367
R771 B.n792 B.n791 163.367
R772 B.n792 B.n21 163.367
R773 B.n796 B.n21 163.367
R774 B.n797 B.n796 163.367
R775 B.n798 B.n797 163.367
R776 B.n798 B.n19 163.367
R777 B.n802 B.n19 163.367
R778 B.n803 B.n802 163.367
R779 B.n804 B.n803 163.367
R780 B.n804 B.n17 163.367
R781 B.n808 B.n17 163.367
R782 B.n809 B.n808 163.367
R783 B.n810 B.n809 163.367
R784 B.n810 B.n15 163.367
R785 B.n814 B.n15 163.367
R786 B.n815 B.n814 163.367
R787 B.n816 B.n815 163.367
R788 B.n816 B.n13 163.367
R789 B.n820 B.n13 163.367
R790 B.n821 B.n820 163.367
R791 B.n822 B.n821 163.367
R792 B.n822 B.n11 163.367
R793 B.n826 B.n11 163.367
R794 B.n827 B.n826 163.367
R795 B.n828 B.n827 163.367
R796 B.n828 B.n9 163.367
R797 B.n832 B.n9 163.367
R798 B.n833 B.n832 163.367
R799 B.n834 B.n833 163.367
R800 B.n834 B.n7 163.367
R801 B.n838 B.n7 163.367
R802 B.n839 B.n838 163.367
R803 B.n840 B.n839 163.367
R804 B.n840 B.n5 163.367
R805 B.n844 B.n5 163.367
R806 B.n845 B.n844 163.367
R807 B.n846 B.n845 163.367
R808 B.n846 B.n3 163.367
R809 B.n850 B.n3 163.367
R810 B.n851 B.n850 163.367
R811 B.n221 B.n2 163.367
R812 B.n222 B.n221 163.367
R813 B.n222 B.n219 163.367
R814 B.n226 B.n219 163.367
R815 B.n227 B.n226 163.367
R816 B.n228 B.n227 163.367
R817 B.n228 B.n217 163.367
R818 B.n232 B.n217 163.367
R819 B.n233 B.n232 163.367
R820 B.n234 B.n233 163.367
R821 B.n234 B.n215 163.367
R822 B.n238 B.n215 163.367
R823 B.n239 B.n238 163.367
R824 B.n240 B.n239 163.367
R825 B.n240 B.n213 163.367
R826 B.n244 B.n213 163.367
R827 B.n245 B.n244 163.367
R828 B.n246 B.n245 163.367
R829 B.n246 B.n211 163.367
R830 B.n250 B.n211 163.367
R831 B.n251 B.n250 163.367
R832 B.n252 B.n251 163.367
R833 B.n252 B.n209 163.367
R834 B.n256 B.n209 163.367
R835 B.n257 B.n256 163.367
R836 B.n258 B.n257 163.367
R837 B.n258 B.n207 163.367
R838 B.n262 B.n207 163.367
R839 B.n263 B.n262 163.367
R840 B.n264 B.n263 163.367
R841 B.n264 B.n205 163.367
R842 B.n268 B.n205 163.367
R843 B.n269 B.n268 163.367
R844 B.n270 B.n269 163.367
R845 B.n270 B.n203 163.367
R846 B.n274 B.n203 163.367
R847 B.n275 B.n274 163.367
R848 B.n276 B.n275 163.367
R849 B.n276 B.n201 163.367
R850 B.n280 B.n201 163.367
R851 B.n281 B.n280 163.367
R852 B.n282 B.n281 163.367
R853 B.n282 B.n199 163.367
R854 B.n171 B.n170 60.1217
R855 B.n163 B.n162 60.1217
R856 B.n61 B.n60 60.1217
R857 B.n53 B.n52 60.1217
R858 B.n369 B.n171 59.5399
R859 B.n164 B.n163 59.5399
R860 B.n687 B.n61 59.5399
R861 B.n54 B.n53 59.5399
R862 B.n787 B.n24 31.0639
R863 B.n603 B.n602 31.0639
R864 B.n469 B.n134 31.0639
R865 B.n285 B.n284 31.0639
R866 B B.n853 18.0485
R867 B.n788 B.n787 10.6151
R868 B.n789 B.n788 10.6151
R869 B.n789 B.n22 10.6151
R870 B.n793 B.n22 10.6151
R871 B.n794 B.n793 10.6151
R872 B.n795 B.n794 10.6151
R873 B.n795 B.n20 10.6151
R874 B.n799 B.n20 10.6151
R875 B.n800 B.n799 10.6151
R876 B.n801 B.n800 10.6151
R877 B.n801 B.n18 10.6151
R878 B.n805 B.n18 10.6151
R879 B.n806 B.n805 10.6151
R880 B.n807 B.n806 10.6151
R881 B.n807 B.n16 10.6151
R882 B.n811 B.n16 10.6151
R883 B.n812 B.n811 10.6151
R884 B.n813 B.n812 10.6151
R885 B.n813 B.n14 10.6151
R886 B.n817 B.n14 10.6151
R887 B.n818 B.n817 10.6151
R888 B.n819 B.n818 10.6151
R889 B.n819 B.n12 10.6151
R890 B.n823 B.n12 10.6151
R891 B.n824 B.n823 10.6151
R892 B.n825 B.n824 10.6151
R893 B.n825 B.n10 10.6151
R894 B.n829 B.n10 10.6151
R895 B.n830 B.n829 10.6151
R896 B.n831 B.n830 10.6151
R897 B.n831 B.n8 10.6151
R898 B.n835 B.n8 10.6151
R899 B.n836 B.n835 10.6151
R900 B.n837 B.n836 10.6151
R901 B.n837 B.n6 10.6151
R902 B.n841 B.n6 10.6151
R903 B.n842 B.n841 10.6151
R904 B.n843 B.n842 10.6151
R905 B.n843 B.n4 10.6151
R906 B.n847 B.n4 10.6151
R907 B.n848 B.n847 10.6151
R908 B.n849 B.n848 10.6151
R909 B.n849 B.n0 10.6151
R910 B.n783 B.n24 10.6151
R911 B.n783 B.n782 10.6151
R912 B.n782 B.n781 10.6151
R913 B.n781 B.n26 10.6151
R914 B.n777 B.n26 10.6151
R915 B.n777 B.n776 10.6151
R916 B.n776 B.n775 10.6151
R917 B.n775 B.n28 10.6151
R918 B.n771 B.n28 10.6151
R919 B.n771 B.n770 10.6151
R920 B.n770 B.n769 10.6151
R921 B.n769 B.n30 10.6151
R922 B.n765 B.n30 10.6151
R923 B.n765 B.n764 10.6151
R924 B.n764 B.n763 10.6151
R925 B.n763 B.n32 10.6151
R926 B.n759 B.n32 10.6151
R927 B.n759 B.n758 10.6151
R928 B.n758 B.n757 10.6151
R929 B.n757 B.n34 10.6151
R930 B.n753 B.n34 10.6151
R931 B.n753 B.n752 10.6151
R932 B.n752 B.n751 10.6151
R933 B.n751 B.n36 10.6151
R934 B.n747 B.n36 10.6151
R935 B.n747 B.n746 10.6151
R936 B.n746 B.n745 10.6151
R937 B.n745 B.n38 10.6151
R938 B.n741 B.n38 10.6151
R939 B.n741 B.n740 10.6151
R940 B.n740 B.n739 10.6151
R941 B.n739 B.n40 10.6151
R942 B.n735 B.n40 10.6151
R943 B.n735 B.n734 10.6151
R944 B.n734 B.n733 10.6151
R945 B.n733 B.n42 10.6151
R946 B.n729 B.n42 10.6151
R947 B.n729 B.n728 10.6151
R948 B.n728 B.n727 10.6151
R949 B.n727 B.n44 10.6151
R950 B.n723 B.n44 10.6151
R951 B.n723 B.n722 10.6151
R952 B.n722 B.n721 10.6151
R953 B.n721 B.n46 10.6151
R954 B.n717 B.n46 10.6151
R955 B.n717 B.n716 10.6151
R956 B.n716 B.n715 10.6151
R957 B.n715 B.n48 10.6151
R958 B.n711 B.n48 10.6151
R959 B.n711 B.n710 10.6151
R960 B.n710 B.n709 10.6151
R961 B.n709 B.n50 10.6151
R962 B.n705 B.n50 10.6151
R963 B.n705 B.n704 10.6151
R964 B.n704 B.n703 10.6151
R965 B.n700 B.n699 10.6151
R966 B.n699 B.n698 10.6151
R967 B.n698 B.n56 10.6151
R968 B.n694 B.n56 10.6151
R969 B.n694 B.n693 10.6151
R970 B.n693 B.n692 10.6151
R971 B.n692 B.n58 10.6151
R972 B.n688 B.n58 10.6151
R973 B.n686 B.n685 10.6151
R974 B.n685 B.n62 10.6151
R975 B.n681 B.n62 10.6151
R976 B.n681 B.n680 10.6151
R977 B.n680 B.n679 10.6151
R978 B.n679 B.n64 10.6151
R979 B.n675 B.n64 10.6151
R980 B.n675 B.n674 10.6151
R981 B.n674 B.n673 10.6151
R982 B.n673 B.n66 10.6151
R983 B.n669 B.n66 10.6151
R984 B.n669 B.n668 10.6151
R985 B.n668 B.n667 10.6151
R986 B.n667 B.n68 10.6151
R987 B.n663 B.n68 10.6151
R988 B.n663 B.n662 10.6151
R989 B.n662 B.n661 10.6151
R990 B.n661 B.n70 10.6151
R991 B.n657 B.n70 10.6151
R992 B.n657 B.n656 10.6151
R993 B.n656 B.n655 10.6151
R994 B.n655 B.n72 10.6151
R995 B.n651 B.n72 10.6151
R996 B.n651 B.n650 10.6151
R997 B.n650 B.n649 10.6151
R998 B.n649 B.n74 10.6151
R999 B.n645 B.n74 10.6151
R1000 B.n645 B.n644 10.6151
R1001 B.n644 B.n643 10.6151
R1002 B.n643 B.n76 10.6151
R1003 B.n639 B.n76 10.6151
R1004 B.n639 B.n638 10.6151
R1005 B.n638 B.n637 10.6151
R1006 B.n637 B.n78 10.6151
R1007 B.n633 B.n78 10.6151
R1008 B.n633 B.n632 10.6151
R1009 B.n632 B.n631 10.6151
R1010 B.n631 B.n80 10.6151
R1011 B.n627 B.n80 10.6151
R1012 B.n627 B.n626 10.6151
R1013 B.n626 B.n625 10.6151
R1014 B.n625 B.n82 10.6151
R1015 B.n621 B.n82 10.6151
R1016 B.n621 B.n620 10.6151
R1017 B.n620 B.n619 10.6151
R1018 B.n619 B.n84 10.6151
R1019 B.n615 B.n84 10.6151
R1020 B.n615 B.n614 10.6151
R1021 B.n614 B.n613 10.6151
R1022 B.n613 B.n86 10.6151
R1023 B.n609 B.n86 10.6151
R1024 B.n609 B.n608 10.6151
R1025 B.n608 B.n607 10.6151
R1026 B.n607 B.n88 10.6151
R1027 B.n603 B.n88 10.6151
R1028 B.n602 B.n601 10.6151
R1029 B.n601 B.n90 10.6151
R1030 B.n597 B.n90 10.6151
R1031 B.n597 B.n596 10.6151
R1032 B.n596 B.n595 10.6151
R1033 B.n595 B.n92 10.6151
R1034 B.n591 B.n92 10.6151
R1035 B.n591 B.n590 10.6151
R1036 B.n590 B.n589 10.6151
R1037 B.n589 B.n94 10.6151
R1038 B.n585 B.n94 10.6151
R1039 B.n585 B.n584 10.6151
R1040 B.n584 B.n583 10.6151
R1041 B.n583 B.n96 10.6151
R1042 B.n579 B.n96 10.6151
R1043 B.n579 B.n578 10.6151
R1044 B.n578 B.n577 10.6151
R1045 B.n577 B.n98 10.6151
R1046 B.n573 B.n98 10.6151
R1047 B.n573 B.n572 10.6151
R1048 B.n572 B.n571 10.6151
R1049 B.n571 B.n100 10.6151
R1050 B.n567 B.n100 10.6151
R1051 B.n567 B.n566 10.6151
R1052 B.n566 B.n565 10.6151
R1053 B.n565 B.n102 10.6151
R1054 B.n561 B.n102 10.6151
R1055 B.n561 B.n560 10.6151
R1056 B.n560 B.n559 10.6151
R1057 B.n559 B.n104 10.6151
R1058 B.n555 B.n104 10.6151
R1059 B.n555 B.n554 10.6151
R1060 B.n554 B.n553 10.6151
R1061 B.n553 B.n106 10.6151
R1062 B.n549 B.n106 10.6151
R1063 B.n549 B.n548 10.6151
R1064 B.n548 B.n547 10.6151
R1065 B.n547 B.n108 10.6151
R1066 B.n543 B.n108 10.6151
R1067 B.n543 B.n542 10.6151
R1068 B.n542 B.n541 10.6151
R1069 B.n541 B.n110 10.6151
R1070 B.n537 B.n110 10.6151
R1071 B.n537 B.n536 10.6151
R1072 B.n536 B.n535 10.6151
R1073 B.n535 B.n112 10.6151
R1074 B.n531 B.n112 10.6151
R1075 B.n531 B.n530 10.6151
R1076 B.n530 B.n529 10.6151
R1077 B.n529 B.n114 10.6151
R1078 B.n525 B.n114 10.6151
R1079 B.n525 B.n524 10.6151
R1080 B.n524 B.n523 10.6151
R1081 B.n523 B.n116 10.6151
R1082 B.n519 B.n116 10.6151
R1083 B.n519 B.n518 10.6151
R1084 B.n518 B.n517 10.6151
R1085 B.n517 B.n118 10.6151
R1086 B.n513 B.n118 10.6151
R1087 B.n513 B.n512 10.6151
R1088 B.n512 B.n511 10.6151
R1089 B.n511 B.n120 10.6151
R1090 B.n507 B.n120 10.6151
R1091 B.n507 B.n506 10.6151
R1092 B.n506 B.n505 10.6151
R1093 B.n505 B.n122 10.6151
R1094 B.n501 B.n122 10.6151
R1095 B.n501 B.n500 10.6151
R1096 B.n500 B.n499 10.6151
R1097 B.n499 B.n124 10.6151
R1098 B.n495 B.n124 10.6151
R1099 B.n495 B.n494 10.6151
R1100 B.n494 B.n493 10.6151
R1101 B.n493 B.n126 10.6151
R1102 B.n489 B.n126 10.6151
R1103 B.n489 B.n488 10.6151
R1104 B.n488 B.n487 10.6151
R1105 B.n487 B.n128 10.6151
R1106 B.n483 B.n128 10.6151
R1107 B.n483 B.n482 10.6151
R1108 B.n482 B.n481 10.6151
R1109 B.n481 B.n130 10.6151
R1110 B.n477 B.n130 10.6151
R1111 B.n477 B.n476 10.6151
R1112 B.n476 B.n475 10.6151
R1113 B.n475 B.n132 10.6151
R1114 B.n471 B.n132 10.6151
R1115 B.n471 B.n470 10.6151
R1116 B.n470 B.n469 10.6151
R1117 B.n220 B.n1 10.6151
R1118 B.n223 B.n220 10.6151
R1119 B.n224 B.n223 10.6151
R1120 B.n225 B.n224 10.6151
R1121 B.n225 B.n218 10.6151
R1122 B.n229 B.n218 10.6151
R1123 B.n230 B.n229 10.6151
R1124 B.n231 B.n230 10.6151
R1125 B.n231 B.n216 10.6151
R1126 B.n235 B.n216 10.6151
R1127 B.n236 B.n235 10.6151
R1128 B.n237 B.n236 10.6151
R1129 B.n237 B.n214 10.6151
R1130 B.n241 B.n214 10.6151
R1131 B.n242 B.n241 10.6151
R1132 B.n243 B.n242 10.6151
R1133 B.n243 B.n212 10.6151
R1134 B.n247 B.n212 10.6151
R1135 B.n248 B.n247 10.6151
R1136 B.n249 B.n248 10.6151
R1137 B.n249 B.n210 10.6151
R1138 B.n253 B.n210 10.6151
R1139 B.n254 B.n253 10.6151
R1140 B.n255 B.n254 10.6151
R1141 B.n255 B.n208 10.6151
R1142 B.n259 B.n208 10.6151
R1143 B.n260 B.n259 10.6151
R1144 B.n261 B.n260 10.6151
R1145 B.n261 B.n206 10.6151
R1146 B.n265 B.n206 10.6151
R1147 B.n266 B.n265 10.6151
R1148 B.n267 B.n266 10.6151
R1149 B.n267 B.n204 10.6151
R1150 B.n271 B.n204 10.6151
R1151 B.n272 B.n271 10.6151
R1152 B.n273 B.n272 10.6151
R1153 B.n273 B.n202 10.6151
R1154 B.n277 B.n202 10.6151
R1155 B.n278 B.n277 10.6151
R1156 B.n279 B.n278 10.6151
R1157 B.n279 B.n200 10.6151
R1158 B.n283 B.n200 10.6151
R1159 B.n284 B.n283 10.6151
R1160 B.n285 B.n198 10.6151
R1161 B.n289 B.n198 10.6151
R1162 B.n290 B.n289 10.6151
R1163 B.n291 B.n290 10.6151
R1164 B.n291 B.n196 10.6151
R1165 B.n295 B.n196 10.6151
R1166 B.n296 B.n295 10.6151
R1167 B.n297 B.n296 10.6151
R1168 B.n297 B.n194 10.6151
R1169 B.n301 B.n194 10.6151
R1170 B.n302 B.n301 10.6151
R1171 B.n303 B.n302 10.6151
R1172 B.n303 B.n192 10.6151
R1173 B.n307 B.n192 10.6151
R1174 B.n308 B.n307 10.6151
R1175 B.n309 B.n308 10.6151
R1176 B.n309 B.n190 10.6151
R1177 B.n313 B.n190 10.6151
R1178 B.n314 B.n313 10.6151
R1179 B.n315 B.n314 10.6151
R1180 B.n315 B.n188 10.6151
R1181 B.n319 B.n188 10.6151
R1182 B.n320 B.n319 10.6151
R1183 B.n321 B.n320 10.6151
R1184 B.n321 B.n186 10.6151
R1185 B.n325 B.n186 10.6151
R1186 B.n326 B.n325 10.6151
R1187 B.n327 B.n326 10.6151
R1188 B.n327 B.n184 10.6151
R1189 B.n331 B.n184 10.6151
R1190 B.n332 B.n331 10.6151
R1191 B.n333 B.n332 10.6151
R1192 B.n333 B.n182 10.6151
R1193 B.n337 B.n182 10.6151
R1194 B.n338 B.n337 10.6151
R1195 B.n339 B.n338 10.6151
R1196 B.n339 B.n180 10.6151
R1197 B.n343 B.n180 10.6151
R1198 B.n344 B.n343 10.6151
R1199 B.n345 B.n344 10.6151
R1200 B.n345 B.n178 10.6151
R1201 B.n349 B.n178 10.6151
R1202 B.n350 B.n349 10.6151
R1203 B.n351 B.n350 10.6151
R1204 B.n351 B.n176 10.6151
R1205 B.n355 B.n176 10.6151
R1206 B.n356 B.n355 10.6151
R1207 B.n357 B.n356 10.6151
R1208 B.n357 B.n174 10.6151
R1209 B.n361 B.n174 10.6151
R1210 B.n362 B.n361 10.6151
R1211 B.n363 B.n362 10.6151
R1212 B.n363 B.n172 10.6151
R1213 B.n367 B.n172 10.6151
R1214 B.n368 B.n367 10.6151
R1215 B.n370 B.n168 10.6151
R1216 B.n374 B.n168 10.6151
R1217 B.n375 B.n374 10.6151
R1218 B.n376 B.n375 10.6151
R1219 B.n376 B.n166 10.6151
R1220 B.n380 B.n166 10.6151
R1221 B.n381 B.n380 10.6151
R1222 B.n382 B.n381 10.6151
R1223 B.n386 B.n385 10.6151
R1224 B.n387 B.n386 10.6151
R1225 B.n387 B.n160 10.6151
R1226 B.n391 B.n160 10.6151
R1227 B.n392 B.n391 10.6151
R1228 B.n393 B.n392 10.6151
R1229 B.n393 B.n158 10.6151
R1230 B.n397 B.n158 10.6151
R1231 B.n398 B.n397 10.6151
R1232 B.n399 B.n398 10.6151
R1233 B.n399 B.n156 10.6151
R1234 B.n403 B.n156 10.6151
R1235 B.n404 B.n403 10.6151
R1236 B.n405 B.n404 10.6151
R1237 B.n405 B.n154 10.6151
R1238 B.n409 B.n154 10.6151
R1239 B.n410 B.n409 10.6151
R1240 B.n411 B.n410 10.6151
R1241 B.n411 B.n152 10.6151
R1242 B.n415 B.n152 10.6151
R1243 B.n416 B.n415 10.6151
R1244 B.n417 B.n416 10.6151
R1245 B.n417 B.n150 10.6151
R1246 B.n421 B.n150 10.6151
R1247 B.n422 B.n421 10.6151
R1248 B.n423 B.n422 10.6151
R1249 B.n423 B.n148 10.6151
R1250 B.n427 B.n148 10.6151
R1251 B.n428 B.n427 10.6151
R1252 B.n429 B.n428 10.6151
R1253 B.n429 B.n146 10.6151
R1254 B.n433 B.n146 10.6151
R1255 B.n434 B.n433 10.6151
R1256 B.n435 B.n434 10.6151
R1257 B.n435 B.n144 10.6151
R1258 B.n439 B.n144 10.6151
R1259 B.n440 B.n439 10.6151
R1260 B.n441 B.n440 10.6151
R1261 B.n441 B.n142 10.6151
R1262 B.n445 B.n142 10.6151
R1263 B.n446 B.n445 10.6151
R1264 B.n447 B.n446 10.6151
R1265 B.n447 B.n140 10.6151
R1266 B.n451 B.n140 10.6151
R1267 B.n452 B.n451 10.6151
R1268 B.n453 B.n452 10.6151
R1269 B.n453 B.n138 10.6151
R1270 B.n457 B.n138 10.6151
R1271 B.n458 B.n457 10.6151
R1272 B.n459 B.n458 10.6151
R1273 B.n459 B.n136 10.6151
R1274 B.n463 B.n136 10.6151
R1275 B.n464 B.n463 10.6151
R1276 B.n465 B.n464 10.6151
R1277 B.n465 B.n134 10.6151
R1278 B.n853 B.n0 8.11757
R1279 B.n853 B.n1 8.11757
R1280 B.n700 B.n54 6.5566
R1281 B.n688 B.n687 6.5566
R1282 B.n370 B.n369 6.5566
R1283 B.n382 B.n164 6.5566
R1284 B.n703 B.n54 4.05904
R1285 B.n687 B.n686 4.05904
R1286 B.n369 B.n368 4.05904
R1287 B.n385 B.n164 4.05904
R1288 VP.n11 VP.t3 179.55
R1289 VP.n13 VP.n12 161.3
R1290 VP.n14 VP.n9 161.3
R1291 VP.n16 VP.n15 161.3
R1292 VP.n17 VP.n8 161.3
R1293 VP.n19 VP.n18 161.3
R1294 VP.n20 VP.n7 161.3
R1295 VP.n43 VP.n0 161.3
R1296 VP.n42 VP.n41 161.3
R1297 VP.n40 VP.n1 161.3
R1298 VP.n39 VP.n38 161.3
R1299 VP.n37 VP.n2 161.3
R1300 VP.n36 VP.n35 161.3
R1301 VP.n34 VP.n3 161.3
R1302 VP.n33 VP.n32 161.3
R1303 VP.n31 VP.n4 161.3
R1304 VP.n30 VP.n29 161.3
R1305 VP.n28 VP.n5 161.3
R1306 VP.n27 VP.n26 161.3
R1307 VP.n25 VP.n6 161.3
R1308 VP.n3 VP.t0 145.47
R1309 VP.n24 VP.t5 145.47
R1310 VP.n44 VP.t2 145.47
R1311 VP.n10 VP.t1 145.47
R1312 VP.n21 VP.t4 145.47
R1313 VP.n24 VP.n23 105.99
R1314 VP.n45 VP.n44 105.99
R1315 VP.n22 VP.n21 105.99
R1316 VP.n23 VP.n22 52.9012
R1317 VP.n11 VP.n10 49.0286
R1318 VP.n30 VP.n5 45.4209
R1319 VP.n38 VP.n1 45.4209
R1320 VP.n15 VP.n8 45.4209
R1321 VP.n31 VP.n30 35.7332
R1322 VP.n38 VP.n37 35.7332
R1323 VP.n15 VP.n14 35.7332
R1324 VP.n26 VP.n25 24.5923
R1325 VP.n26 VP.n5 24.5923
R1326 VP.n32 VP.n31 24.5923
R1327 VP.n32 VP.n3 24.5923
R1328 VP.n36 VP.n3 24.5923
R1329 VP.n37 VP.n36 24.5923
R1330 VP.n42 VP.n1 24.5923
R1331 VP.n43 VP.n42 24.5923
R1332 VP.n19 VP.n8 24.5923
R1333 VP.n20 VP.n19 24.5923
R1334 VP.n13 VP.n10 24.5923
R1335 VP.n14 VP.n13 24.5923
R1336 VP.n12 VP.n11 4.96469
R1337 VP.n25 VP.n24 4.91887
R1338 VP.n44 VP.n43 4.91887
R1339 VP.n21 VP.n20 4.91887
R1340 VP.n22 VP.n7 0.278335
R1341 VP.n23 VP.n6 0.278335
R1342 VP.n45 VP.n0 0.278335
R1343 VP.n12 VP.n9 0.189894
R1344 VP.n16 VP.n9 0.189894
R1345 VP.n17 VP.n16 0.189894
R1346 VP.n18 VP.n17 0.189894
R1347 VP.n18 VP.n7 0.189894
R1348 VP.n27 VP.n6 0.189894
R1349 VP.n28 VP.n27 0.189894
R1350 VP.n29 VP.n28 0.189894
R1351 VP.n29 VP.n4 0.189894
R1352 VP.n33 VP.n4 0.189894
R1353 VP.n34 VP.n33 0.189894
R1354 VP.n35 VP.n34 0.189894
R1355 VP.n35 VP.n2 0.189894
R1356 VP.n39 VP.n2 0.189894
R1357 VP.n40 VP.n39 0.189894
R1358 VP.n41 VP.n40 0.189894
R1359 VP.n41 VP.n0 0.189894
R1360 VP VP.n45 0.153485
R1361 VDD1.n88 VDD1.n0 756.745
R1362 VDD1.n181 VDD1.n93 756.745
R1363 VDD1.n89 VDD1.n88 585
R1364 VDD1.n87 VDD1.n86 585
R1365 VDD1.n4 VDD1.n3 585
R1366 VDD1.n81 VDD1.n80 585
R1367 VDD1.n79 VDD1.n78 585
R1368 VDD1.n77 VDD1.n7 585
R1369 VDD1.n11 VDD1.n8 585
R1370 VDD1.n72 VDD1.n71 585
R1371 VDD1.n70 VDD1.n69 585
R1372 VDD1.n13 VDD1.n12 585
R1373 VDD1.n64 VDD1.n63 585
R1374 VDD1.n62 VDD1.n61 585
R1375 VDD1.n17 VDD1.n16 585
R1376 VDD1.n56 VDD1.n55 585
R1377 VDD1.n54 VDD1.n53 585
R1378 VDD1.n21 VDD1.n20 585
R1379 VDD1.n48 VDD1.n47 585
R1380 VDD1.n46 VDD1.n45 585
R1381 VDD1.n25 VDD1.n24 585
R1382 VDD1.n40 VDD1.n39 585
R1383 VDD1.n38 VDD1.n37 585
R1384 VDD1.n29 VDD1.n28 585
R1385 VDD1.n32 VDD1.n31 585
R1386 VDD1.n124 VDD1.n123 585
R1387 VDD1.n121 VDD1.n120 585
R1388 VDD1.n130 VDD1.n129 585
R1389 VDD1.n132 VDD1.n131 585
R1390 VDD1.n117 VDD1.n116 585
R1391 VDD1.n138 VDD1.n137 585
R1392 VDD1.n140 VDD1.n139 585
R1393 VDD1.n113 VDD1.n112 585
R1394 VDD1.n146 VDD1.n145 585
R1395 VDD1.n148 VDD1.n147 585
R1396 VDD1.n109 VDD1.n108 585
R1397 VDD1.n154 VDD1.n153 585
R1398 VDD1.n156 VDD1.n155 585
R1399 VDD1.n105 VDD1.n104 585
R1400 VDD1.n162 VDD1.n161 585
R1401 VDD1.n165 VDD1.n164 585
R1402 VDD1.n163 VDD1.n101 585
R1403 VDD1.n170 VDD1.n100 585
R1404 VDD1.n172 VDD1.n171 585
R1405 VDD1.n174 VDD1.n173 585
R1406 VDD1.n97 VDD1.n96 585
R1407 VDD1.n180 VDD1.n179 585
R1408 VDD1.n182 VDD1.n181 585
R1409 VDD1.t1 VDD1.n30 327.466
R1410 VDD1.t0 VDD1.n122 327.466
R1411 VDD1.n88 VDD1.n87 171.744
R1412 VDD1.n87 VDD1.n3 171.744
R1413 VDD1.n80 VDD1.n3 171.744
R1414 VDD1.n80 VDD1.n79 171.744
R1415 VDD1.n79 VDD1.n7 171.744
R1416 VDD1.n11 VDD1.n7 171.744
R1417 VDD1.n71 VDD1.n11 171.744
R1418 VDD1.n71 VDD1.n70 171.744
R1419 VDD1.n70 VDD1.n12 171.744
R1420 VDD1.n63 VDD1.n12 171.744
R1421 VDD1.n63 VDD1.n62 171.744
R1422 VDD1.n62 VDD1.n16 171.744
R1423 VDD1.n55 VDD1.n16 171.744
R1424 VDD1.n55 VDD1.n54 171.744
R1425 VDD1.n54 VDD1.n20 171.744
R1426 VDD1.n47 VDD1.n20 171.744
R1427 VDD1.n47 VDD1.n46 171.744
R1428 VDD1.n46 VDD1.n24 171.744
R1429 VDD1.n39 VDD1.n24 171.744
R1430 VDD1.n39 VDD1.n38 171.744
R1431 VDD1.n38 VDD1.n28 171.744
R1432 VDD1.n31 VDD1.n28 171.744
R1433 VDD1.n123 VDD1.n120 171.744
R1434 VDD1.n130 VDD1.n120 171.744
R1435 VDD1.n131 VDD1.n130 171.744
R1436 VDD1.n131 VDD1.n116 171.744
R1437 VDD1.n138 VDD1.n116 171.744
R1438 VDD1.n139 VDD1.n138 171.744
R1439 VDD1.n139 VDD1.n112 171.744
R1440 VDD1.n146 VDD1.n112 171.744
R1441 VDD1.n147 VDD1.n146 171.744
R1442 VDD1.n147 VDD1.n108 171.744
R1443 VDD1.n154 VDD1.n108 171.744
R1444 VDD1.n155 VDD1.n154 171.744
R1445 VDD1.n155 VDD1.n104 171.744
R1446 VDD1.n162 VDD1.n104 171.744
R1447 VDD1.n164 VDD1.n162 171.744
R1448 VDD1.n164 VDD1.n163 171.744
R1449 VDD1.n163 VDD1.n100 171.744
R1450 VDD1.n172 VDD1.n100 171.744
R1451 VDD1.n173 VDD1.n172 171.744
R1452 VDD1.n173 VDD1.n96 171.744
R1453 VDD1.n180 VDD1.n96 171.744
R1454 VDD1.n181 VDD1.n180 171.744
R1455 VDD1.n31 VDD1.t1 85.8723
R1456 VDD1.n123 VDD1.t0 85.8723
R1457 VDD1.n187 VDD1.n186 68.4531
R1458 VDD1.n189 VDD1.n188 67.8403
R1459 VDD1 VDD1.n92 49.3751
R1460 VDD1.n187 VDD1.n185 49.2616
R1461 VDD1.n189 VDD1.n187 48.7337
R1462 VDD1.n32 VDD1.n30 16.3895
R1463 VDD1.n124 VDD1.n122 16.3895
R1464 VDD1.n78 VDD1.n77 13.1884
R1465 VDD1.n171 VDD1.n170 13.1884
R1466 VDD1.n81 VDD1.n6 12.8005
R1467 VDD1.n76 VDD1.n8 12.8005
R1468 VDD1.n33 VDD1.n29 12.8005
R1469 VDD1.n125 VDD1.n121 12.8005
R1470 VDD1.n169 VDD1.n101 12.8005
R1471 VDD1.n174 VDD1.n99 12.8005
R1472 VDD1.n82 VDD1.n4 12.0247
R1473 VDD1.n73 VDD1.n72 12.0247
R1474 VDD1.n37 VDD1.n36 12.0247
R1475 VDD1.n129 VDD1.n128 12.0247
R1476 VDD1.n166 VDD1.n165 12.0247
R1477 VDD1.n175 VDD1.n97 12.0247
R1478 VDD1.n86 VDD1.n85 11.249
R1479 VDD1.n69 VDD1.n10 11.249
R1480 VDD1.n40 VDD1.n27 11.249
R1481 VDD1.n132 VDD1.n119 11.249
R1482 VDD1.n161 VDD1.n103 11.249
R1483 VDD1.n179 VDD1.n178 11.249
R1484 VDD1.n89 VDD1.n2 10.4732
R1485 VDD1.n68 VDD1.n13 10.4732
R1486 VDD1.n41 VDD1.n25 10.4732
R1487 VDD1.n133 VDD1.n117 10.4732
R1488 VDD1.n160 VDD1.n105 10.4732
R1489 VDD1.n182 VDD1.n95 10.4732
R1490 VDD1.n90 VDD1.n0 9.69747
R1491 VDD1.n65 VDD1.n64 9.69747
R1492 VDD1.n45 VDD1.n44 9.69747
R1493 VDD1.n137 VDD1.n136 9.69747
R1494 VDD1.n157 VDD1.n156 9.69747
R1495 VDD1.n183 VDD1.n93 9.69747
R1496 VDD1.n92 VDD1.n91 9.45567
R1497 VDD1.n185 VDD1.n184 9.45567
R1498 VDD1.n58 VDD1.n57 9.3005
R1499 VDD1.n60 VDD1.n59 9.3005
R1500 VDD1.n15 VDD1.n14 9.3005
R1501 VDD1.n66 VDD1.n65 9.3005
R1502 VDD1.n68 VDD1.n67 9.3005
R1503 VDD1.n10 VDD1.n9 9.3005
R1504 VDD1.n74 VDD1.n73 9.3005
R1505 VDD1.n76 VDD1.n75 9.3005
R1506 VDD1.n91 VDD1.n90 9.3005
R1507 VDD1.n2 VDD1.n1 9.3005
R1508 VDD1.n85 VDD1.n84 9.3005
R1509 VDD1.n83 VDD1.n82 9.3005
R1510 VDD1.n6 VDD1.n5 9.3005
R1511 VDD1.n19 VDD1.n18 9.3005
R1512 VDD1.n52 VDD1.n51 9.3005
R1513 VDD1.n50 VDD1.n49 9.3005
R1514 VDD1.n23 VDD1.n22 9.3005
R1515 VDD1.n44 VDD1.n43 9.3005
R1516 VDD1.n42 VDD1.n41 9.3005
R1517 VDD1.n27 VDD1.n26 9.3005
R1518 VDD1.n36 VDD1.n35 9.3005
R1519 VDD1.n34 VDD1.n33 9.3005
R1520 VDD1.n184 VDD1.n183 9.3005
R1521 VDD1.n95 VDD1.n94 9.3005
R1522 VDD1.n178 VDD1.n177 9.3005
R1523 VDD1.n176 VDD1.n175 9.3005
R1524 VDD1.n99 VDD1.n98 9.3005
R1525 VDD1.n144 VDD1.n143 9.3005
R1526 VDD1.n142 VDD1.n141 9.3005
R1527 VDD1.n115 VDD1.n114 9.3005
R1528 VDD1.n136 VDD1.n135 9.3005
R1529 VDD1.n134 VDD1.n133 9.3005
R1530 VDD1.n119 VDD1.n118 9.3005
R1531 VDD1.n128 VDD1.n127 9.3005
R1532 VDD1.n126 VDD1.n125 9.3005
R1533 VDD1.n111 VDD1.n110 9.3005
R1534 VDD1.n150 VDD1.n149 9.3005
R1535 VDD1.n152 VDD1.n151 9.3005
R1536 VDD1.n107 VDD1.n106 9.3005
R1537 VDD1.n158 VDD1.n157 9.3005
R1538 VDD1.n160 VDD1.n159 9.3005
R1539 VDD1.n103 VDD1.n102 9.3005
R1540 VDD1.n167 VDD1.n166 9.3005
R1541 VDD1.n169 VDD1.n168 9.3005
R1542 VDD1.n61 VDD1.n15 8.92171
R1543 VDD1.n48 VDD1.n23 8.92171
R1544 VDD1.n140 VDD1.n115 8.92171
R1545 VDD1.n153 VDD1.n107 8.92171
R1546 VDD1.n60 VDD1.n17 8.14595
R1547 VDD1.n49 VDD1.n21 8.14595
R1548 VDD1.n141 VDD1.n113 8.14595
R1549 VDD1.n152 VDD1.n109 8.14595
R1550 VDD1.n57 VDD1.n56 7.3702
R1551 VDD1.n53 VDD1.n52 7.3702
R1552 VDD1.n145 VDD1.n144 7.3702
R1553 VDD1.n149 VDD1.n148 7.3702
R1554 VDD1.n56 VDD1.n19 6.59444
R1555 VDD1.n53 VDD1.n19 6.59444
R1556 VDD1.n145 VDD1.n111 6.59444
R1557 VDD1.n148 VDD1.n111 6.59444
R1558 VDD1.n57 VDD1.n17 5.81868
R1559 VDD1.n52 VDD1.n21 5.81868
R1560 VDD1.n144 VDD1.n113 5.81868
R1561 VDD1.n149 VDD1.n109 5.81868
R1562 VDD1.n61 VDD1.n60 5.04292
R1563 VDD1.n49 VDD1.n48 5.04292
R1564 VDD1.n141 VDD1.n140 5.04292
R1565 VDD1.n153 VDD1.n152 5.04292
R1566 VDD1.n92 VDD1.n0 4.26717
R1567 VDD1.n64 VDD1.n15 4.26717
R1568 VDD1.n45 VDD1.n23 4.26717
R1569 VDD1.n137 VDD1.n115 4.26717
R1570 VDD1.n156 VDD1.n107 4.26717
R1571 VDD1.n185 VDD1.n93 4.26717
R1572 VDD1.n34 VDD1.n30 3.70982
R1573 VDD1.n126 VDD1.n122 3.70982
R1574 VDD1.n90 VDD1.n89 3.49141
R1575 VDD1.n65 VDD1.n13 3.49141
R1576 VDD1.n44 VDD1.n25 3.49141
R1577 VDD1.n136 VDD1.n117 3.49141
R1578 VDD1.n157 VDD1.n105 3.49141
R1579 VDD1.n183 VDD1.n182 3.49141
R1580 VDD1.n86 VDD1.n2 2.71565
R1581 VDD1.n69 VDD1.n68 2.71565
R1582 VDD1.n41 VDD1.n40 2.71565
R1583 VDD1.n133 VDD1.n132 2.71565
R1584 VDD1.n161 VDD1.n160 2.71565
R1585 VDD1.n179 VDD1.n95 2.71565
R1586 VDD1.n188 VDD1.t3 1.94458
R1587 VDD1.n188 VDD1.t2 1.94458
R1588 VDD1.n186 VDD1.t4 1.94458
R1589 VDD1.n186 VDD1.t5 1.94458
R1590 VDD1.n85 VDD1.n4 1.93989
R1591 VDD1.n72 VDD1.n10 1.93989
R1592 VDD1.n37 VDD1.n27 1.93989
R1593 VDD1.n129 VDD1.n119 1.93989
R1594 VDD1.n165 VDD1.n103 1.93989
R1595 VDD1.n178 VDD1.n97 1.93989
R1596 VDD1.n82 VDD1.n81 1.16414
R1597 VDD1.n73 VDD1.n8 1.16414
R1598 VDD1.n36 VDD1.n29 1.16414
R1599 VDD1.n128 VDD1.n121 1.16414
R1600 VDD1.n166 VDD1.n101 1.16414
R1601 VDD1.n175 VDD1.n174 1.16414
R1602 VDD1 VDD1.n189 0.610414
R1603 VDD1.n78 VDD1.n6 0.388379
R1604 VDD1.n77 VDD1.n76 0.388379
R1605 VDD1.n33 VDD1.n32 0.388379
R1606 VDD1.n125 VDD1.n124 0.388379
R1607 VDD1.n170 VDD1.n169 0.388379
R1608 VDD1.n171 VDD1.n99 0.388379
R1609 VDD1.n91 VDD1.n1 0.155672
R1610 VDD1.n84 VDD1.n1 0.155672
R1611 VDD1.n84 VDD1.n83 0.155672
R1612 VDD1.n83 VDD1.n5 0.155672
R1613 VDD1.n75 VDD1.n5 0.155672
R1614 VDD1.n75 VDD1.n74 0.155672
R1615 VDD1.n74 VDD1.n9 0.155672
R1616 VDD1.n67 VDD1.n9 0.155672
R1617 VDD1.n67 VDD1.n66 0.155672
R1618 VDD1.n66 VDD1.n14 0.155672
R1619 VDD1.n59 VDD1.n14 0.155672
R1620 VDD1.n59 VDD1.n58 0.155672
R1621 VDD1.n58 VDD1.n18 0.155672
R1622 VDD1.n51 VDD1.n18 0.155672
R1623 VDD1.n51 VDD1.n50 0.155672
R1624 VDD1.n50 VDD1.n22 0.155672
R1625 VDD1.n43 VDD1.n22 0.155672
R1626 VDD1.n43 VDD1.n42 0.155672
R1627 VDD1.n42 VDD1.n26 0.155672
R1628 VDD1.n35 VDD1.n26 0.155672
R1629 VDD1.n35 VDD1.n34 0.155672
R1630 VDD1.n127 VDD1.n126 0.155672
R1631 VDD1.n127 VDD1.n118 0.155672
R1632 VDD1.n134 VDD1.n118 0.155672
R1633 VDD1.n135 VDD1.n134 0.155672
R1634 VDD1.n135 VDD1.n114 0.155672
R1635 VDD1.n142 VDD1.n114 0.155672
R1636 VDD1.n143 VDD1.n142 0.155672
R1637 VDD1.n143 VDD1.n110 0.155672
R1638 VDD1.n150 VDD1.n110 0.155672
R1639 VDD1.n151 VDD1.n150 0.155672
R1640 VDD1.n151 VDD1.n106 0.155672
R1641 VDD1.n158 VDD1.n106 0.155672
R1642 VDD1.n159 VDD1.n158 0.155672
R1643 VDD1.n159 VDD1.n102 0.155672
R1644 VDD1.n167 VDD1.n102 0.155672
R1645 VDD1.n168 VDD1.n167 0.155672
R1646 VDD1.n168 VDD1.n98 0.155672
R1647 VDD1.n176 VDD1.n98 0.155672
R1648 VDD1.n177 VDD1.n176 0.155672
R1649 VDD1.n177 VDD1.n94 0.155672
R1650 VDD1.n184 VDD1.n94 0.155672
R1651 VTAIL.n378 VTAIL.n290 756.745
R1652 VTAIL.n90 VTAIL.n2 756.745
R1653 VTAIL.n284 VTAIL.n196 756.745
R1654 VTAIL.n188 VTAIL.n100 756.745
R1655 VTAIL.n321 VTAIL.n320 585
R1656 VTAIL.n318 VTAIL.n317 585
R1657 VTAIL.n327 VTAIL.n326 585
R1658 VTAIL.n329 VTAIL.n328 585
R1659 VTAIL.n314 VTAIL.n313 585
R1660 VTAIL.n335 VTAIL.n334 585
R1661 VTAIL.n337 VTAIL.n336 585
R1662 VTAIL.n310 VTAIL.n309 585
R1663 VTAIL.n343 VTAIL.n342 585
R1664 VTAIL.n345 VTAIL.n344 585
R1665 VTAIL.n306 VTAIL.n305 585
R1666 VTAIL.n351 VTAIL.n350 585
R1667 VTAIL.n353 VTAIL.n352 585
R1668 VTAIL.n302 VTAIL.n301 585
R1669 VTAIL.n359 VTAIL.n358 585
R1670 VTAIL.n362 VTAIL.n361 585
R1671 VTAIL.n360 VTAIL.n298 585
R1672 VTAIL.n367 VTAIL.n297 585
R1673 VTAIL.n369 VTAIL.n368 585
R1674 VTAIL.n371 VTAIL.n370 585
R1675 VTAIL.n294 VTAIL.n293 585
R1676 VTAIL.n377 VTAIL.n376 585
R1677 VTAIL.n379 VTAIL.n378 585
R1678 VTAIL.n33 VTAIL.n32 585
R1679 VTAIL.n30 VTAIL.n29 585
R1680 VTAIL.n39 VTAIL.n38 585
R1681 VTAIL.n41 VTAIL.n40 585
R1682 VTAIL.n26 VTAIL.n25 585
R1683 VTAIL.n47 VTAIL.n46 585
R1684 VTAIL.n49 VTAIL.n48 585
R1685 VTAIL.n22 VTAIL.n21 585
R1686 VTAIL.n55 VTAIL.n54 585
R1687 VTAIL.n57 VTAIL.n56 585
R1688 VTAIL.n18 VTAIL.n17 585
R1689 VTAIL.n63 VTAIL.n62 585
R1690 VTAIL.n65 VTAIL.n64 585
R1691 VTAIL.n14 VTAIL.n13 585
R1692 VTAIL.n71 VTAIL.n70 585
R1693 VTAIL.n74 VTAIL.n73 585
R1694 VTAIL.n72 VTAIL.n10 585
R1695 VTAIL.n79 VTAIL.n9 585
R1696 VTAIL.n81 VTAIL.n80 585
R1697 VTAIL.n83 VTAIL.n82 585
R1698 VTAIL.n6 VTAIL.n5 585
R1699 VTAIL.n89 VTAIL.n88 585
R1700 VTAIL.n91 VTAIL.n90 585
R1701 VTAIL.n285 VTAIL.n284 585
R1702 VTAIL.n283 VTAIL.n282 585
R1703 VTAIL.n200 VTAIL.n199 585
R1704 VTAIL.n277 VTAIL.n276 585
R1705 VTAIL.n275 VTAIL.n274 585
R1706 VTAIL.n273 VTAIL.n203 585
R1707 VTAIL.n207 VTAIL.n204 585
R1708 VTAIL.n268 VTAIL.n267 585
R1709 VTAIL.n266 VTAIL.n265 585
R1710 VTAIL.n209 VTAIL.n208 585
R1711 VTAIL.n260 VTAIL.n259 585
R1712 VTAIL.n258 VTAIL.n257 585
R1713 VTAIL.n213 VTAIL.n212 585
R1714 VTAIL.n252 VTAIL.n251 585
R1715 VTAIL.n250 VTAIL.n249 585
R1716 VTAIL.n217 VTAIL.n216 585
R1717 VTAIL.n244 VTAIL.n243 585
R1718 VTAIL.n242 VTAIL.n241 585
R1719 VTAIL.n221 VTAIL.n220 585
R1720 VTAIL.n236 VTAIL.n235 585
R1721 VTAIL.n234 VTAIL.n233 585
R1722 VTAIL.n225 VTAIL.n224 585
R1723 VTAIL.n228 VTAIL.n227 585
R1724 VTAIL.n189 VTAIL.n188 585
R1725 VTAIL.n187 VTAIL.n186 585
R1726 VTAIL.n104 VTAIL.n103 585
R1727 VTAIL.n181 VTAIL.n180 585
R1728 VTAIL.n179 VTAIL.n178 585
R1729 VTAIL.n177 VTAIL.n107 585
R1730 VTAIL.n111 VTAIL.n108 585
R1731 VTAIL.n172 VTAIL.n171 585
R1732 VTAIL.n170 VTAIL.n169 585
R1733 VTAIL.n113 VTAIL.n112 585
R1734 VTAIL.n164 VTAIL.n163 585
R1735 VTAIL.n162 VTAIL.n161 585
R1736 VTAIL.n117 VTAIL.n116 585
R1737 VTAIL.n156 VTAIL.n155 585
R1738 VTAIL.n154 VTAIL.n153 585
R1739 VTAIL.n121 VTAIL.n120 585
R1740 VTAIL.n148 VTAIL.n147 585
R1741 VTAIL.n146 VTAIL.n145 585
R1742 VTAIL.n125 VTAIL.n124 585
R1743 VTAIL.n140 VTAIL.n139 585
R1744 VTAIL.n138 VTAIL.n137 585
R1745 VTAIL.n129 VTAIL.n128 585
R1746 VTAIL.n132 VTAIL.n131 585
R1747 VTAIL.t6 VTAIL.n226 327.466
R1748 VTAIL.t1 VTAIL.n130 327.466
R1749 VTAIL.t11 VTAIL.n319 327.466
R1750 VTAIL.t8 VTAIL.n31 327.466
R1751 VTAIL.n320 VTAIL.n317 171.744
R1752 VTAIL.n327 VTAIL.n317 171.744
R1753 VTAIL.n328 VTAIL.n327 171.744
R1754 VTAIL.n328 VTAIL.n313 171.744
R1755 VTAIL.n335 VTAIL.n313 171.744
R1756 VTAIL.n336 VTAIL.n335 171.744
R1757 VTAIL.n336 VTAIL.n309 171.744
R1758 VTAIL.n343 VTAIL.n309 171.744
R1759 VTAIL.n344 VTAIL.n343 171.744
R1760 VTAIL.n344 VTAIL.n305 171.744
R1761 VTAIL.n351 VTAIL.n305 171.744
R1762 VTAIL.n352 VTAIL.n351 171.744
R1763 VTAIL.n352 VTAIL.n301 171.744
R1764 VTAIL.n359 VTAIL.n301 171.744
R1765 VTAIL.n361 VTAIL.n359 171.744
R1766 VTAIL.n361 VTAIL.n360 171.744
R1767 VTAIL.n360 VTAIL.n297 171.744
R1768 VTAIL.n369 VTAIL.n297 171.744
R1769 VTAIL.n370 VTAIL.n369 171.744
R1770 VTAIL.n370 VTAIL.n293 171.744
R1771 VTAIL.n377 VTAIL.n293 171.744
R1772 VTAIL.n378 VTAIL.n377 171.744
R1773 VTAIL.n32 VTAIL.n29 171.744
R1774 VTAIL.n39 VTAIL.n29 171.744
R1775 VTAIL.n40 VTAIL.n39 171.744
R1776 VTAIL.n40 VTAIL.n25 171.744
R1777 VTAIL.n47 VTAIL.n25 171.744
R1778 VTAIL.n48 VTAIL.n47 171.744
R1779 VTAIL.n48 VTAIL.n21 171.744
R1780 VTAIL.n55 VTAIL.n21 171.744
R1781 VTAIL.n56 VTAIL.n55 171.744
R1782 VTAIL.n56 VTAIL.n17 171.744
R1783 VTAIL.n63 VTAIL.n17 171.744
R1784 VTAIL.n64 VTAIL.n63 171.744
R1785 VTAIL.n64 VTAIL.n13 171.744
R1786 VTAIL.n71 VTAIL.n13 171.744
R1787 VTAIL.n73 VTAIL.n71 171.744
R1788 VTAIL.n73 VTAIL.n72 171.744
R1789 VTAIL.n72 VTAIL.n9 171.744
R1790 VTAIL.n81 VTAIL.n9 171.744
R1791 VTAIL.n82 VTAIL.n81 171.744
R1792 VTAIL.n82 VTAIL.n5 171.744
R1793 VTAIL.n89 VTAIL.n5 171.744
R1794 VTAIL.n90 VTAIL.n89 171.744
R1795 VTAIL.n284 VTAIL.n283 171.744
R1796 VTAIL.n283 VTAIL.n199 171.744
R1797 VTAIL.n276 VTAIL.n199 171.744
R1798 VTAIL.n276 VTAIL.n275 171.744
R1799 VTAIL.n275 VTAIL.n203 171.744
R1800 VTAIL.n207 VTAIL.n203 171.744
R1801 VTAIL.n267 VTAIL.n207 171.744
R1802 VTAIL.n267 VTAIL.n266 171.744
R1803 VTAIL.n266 VTAIL.n208 171.744
R1804 VTAIL.n259 VTAIL.n208 171.744
R1805 VTAIL.n259 VTAIL.n258 171.744
R1806 VTAIL.n258 VTAIL.n212 171.744
R1807 VTAIL.n251 VTAIL.n212 171.744
R1808 VTAIL.n251 VTAIL.n250 171.744
R1809 VTAIL.n250 VTAIL.n216 171.744
R1810 VTAIL.n243 VTAIL.n216 171.744
R1811 VTAIL.n243 VTAIL.n242 171.744
R1812 VTAIL.n242 VTAIL.n220 171.744
R1813 VTAIL.n235 VTAIL.n220 171.744
R1814 VTAIL.n235 VTAIL.n234 171.744
R1815 VTAIL.n234 VTAIL.n224 171.744
R1816 VTAIL.n227 VTAIL.n224 171.744
R1817 VTAIL.n188 VTAIL.n187 171.744
R1818 VTAIL.n187 VTAIL.n103 171.744
R1819 VTAIL.n180 VTAIL.n103 171.744
R1820 VTAIL.n180 VTAIL.n179 171.744
R1821 VTAIL.n179 VTAIL.n107 171.744
R1822 VTAIL.n111 VTAIL.n107 171.744
R1823 VTAIL.n171 VTAIL.n111 171.744
R1824 VTAIL.n171 VTAIL.n170 171.744
R1825 VTAIL.n170 VTAIL.n112 171.744
R1826 VTAIL.n163 VTAIL.n112 171.744
R1827 VTAIL.n163 VTAIL.n162 171.744
R1828 VTAIL.n162 VTAIL.n116 171.744
R1829 VTAIL.n155 VTAIL.n116 171.744
R1830 VTAIL.n155 VTAIL.n154 171.744
R1831 VTAIL.n154 VTAIL.n120 171.744
R1832 VTAIL.n147 VTAIL.n120 171.744
R1833 VTAIL.n147 VTAIL.n146 171.744
R1834 VTAIL.n146 VTAIL.n124 171.744
R1835 VTAIL.n139 VTAIL.n124 171.744
R1836 VTAIL.n139 VTAIL.n138 171.744
R1837 VTAIL.n138 VTAIL.n128 171.744
R1838 VTAIL.n131 VTAIL.n128 171.744
R1839 VTAIL.n320 VTAIL.t11 85.8723
R1840 VTAIL.n32 VTAIL.t8 85.8723
R1841 VTAIL.n227 VTAIL.t6 85.8723
R1842 VTAIL.n131 VTAIL.t1 85.8723
R1843 VTAIL.n195 VTAIL.n194 51.1617
R1844 VTAIL.n99 VTAIL.n98 51.1617
R1845 VTAIL.n1 VTAIL.n0 51.1615
R1846 VTAIL.n97 VTAIL.n96 51.1615
R1847 VTAIL.n99 VTAIL.n97 32.1255
R1848 VTAIL.n383 VTAIL.n382 30.6338
R1849 VTAIL.n95 VTAIL.n94 30.6338
R1850 VTAIL.n289 VTAIL.n288 30.6338
R1851 VTAIL.n193 VTAIL.n192 30.6338
R1852 VTAIL.n383 VTAIL.n289 29.4531
R1853 VTAIL.n321 VTAIL.n319 16.3895
R1854 VTAIL.n33 VTAIL.n31 16.3895
R1855 VTAIL.n228 VTAIL.n226 16.3895
R1856 VTAIL.n132 VTAIL.n130 16.3895
R1857 VTAIL.n368 VTAIL.n367 13.1884
R1858 VTAIL.n80 VTAIL.n79 13.1884
R1859 VTAIL.n274 VTAIL.n273 13.1884
R1860 VTAIL.n178 VTAIL.n177 13.1884
R1861 VTAIL.n322 VTAIL.n318 12.8005
R1862 VTAIL.n366 VTAIL.n298 12.8005
R1863 VTAIL.n371 VTAIL.n296 12.8005
R1864 VTAIL.n34 VTAIL.n30 12.8005
R1865 VTAIL.n78 VTAIL.n10 12.8005
R1866 VTAIL.n83 VTAIL.n8 12.8005
R1867 VTAIL.n277 VTAIL.n202 12.8005
R1868 VTAIL.n272 VTAIL.n204 12.8005
R1869 VTAIL.n229 VTAIL.n225 12.8005
R1870 VTAIL.n181 VTAIL.n106 12.8005
R1871 VTAIL.n176 VTAIL.n108 12.8005
R1872 VTAIL.n133 VTAIL.n129 12.8005
R1873 VTAIL.n326 VTAIL.n325 12.0247
R1874 VTAIL.n363 VTAIL.n362 12.0247
R1875 VTAIL.n372 VTAIL.n294 12.0247
R1876 VTAIL.n38 VTAIL.n37 12.0247
R1877 VTAIL.n75 VTAIL.n74 12.0247
R1878 VTAIL.n84 VTAIL.n6 12.0247
R1879 VTAIL.n278 VTAIL.n200 12.0247
R1880 VTAIL.n269 VTAIL.n268 12.0247
R1881 VTAIL.n233 VTAIL.n232 12.0247
R1882 VTAIL.n182 VTAIL.n104 12.0247
R1883 VTAIL.n173 VTAIL.n172 12.0247
R1884 VTAIL.n137 VTAIL.n136 12.0247
R1885 VTAIL.n329 VTAIL.n316 11.249
R1886 VTAIL.n358 VTAIL.n300 11.249
R1887 VTAIL.n376 VTAIL.n375 11.249
R1888 VTAIL.n41 VTAIL.n28 11.249
R1889 VTAIL.n70 VTAIL.n12 11.249
R1890 VTAIL.n88 VTAIL.n87 11.249
R1891 VTAIL.n282 VTAIL.n281 11.249
R1892 VTAIL.n265 VTAIL.n206 11.249
R1893 VTAIL.n236 VTAIL.n223 11.249
R1894 VTAIL.n186 VTAIL.n185 11.249
R1895 VTAIL.n169 VTAIL.n110 11.249
R1896 VTAIL.n140 VTAIL.n127 11.249
R1897 VTAIL.n330 VTAIL.n314 10.4732
R1898 VTAIL.n357 VTAIL.n302 10.4732
R1899 VTAIL.n379 VTAIL.n292 10.4732
R1900 VTAIL.n42 VTAIL.n26 10.4732
R1901 VTAIL.n69 VTAIL.n14 10.4732
R1902 VTAIL.n91 VTAIL.n4 10.4732
R1903 VTAIL.n285 VTAIL.n198 10.4732
R1904 VTAIL.n264 VTAIL.n209 10.4732
R1905 VTAIL.n237 VTAIL.n221 10.4732
R1906 VTAIL.n189 VTAIL.n102 10.4732
R1907 VTAIL.n168 VTAIL.n113 10.4732
R1908 VTAIL.n141 VTAIL.n125 10.4732
R1909 VTAIL.n334 VTAIL.n333 9.69747
R1910 VTAIL.n354 VTAIL.n353 9.69747
R1911 VTAIL.n380 VTAIL.n290 9.69747
R1912 VTAIL.n46 VTAIL.n45 9.69747
R1913 VTAIL.n66 VTAIL.n65 9.69747
R1914 VTAIL.n92 VTAIL.n2 9.69747
R1915 VTAIL.n286 VTAIL.n196 9.69747
R1916 VTAIL.n261 VTAIL.n260 9.69747
R1917 VTAIL.n241 VTAIL.n240 9.69747
R1918 VTAIL.n190 VTAIL.n100 9.69747
R1919 VTAIL.n165 VTAIL.n164 9.69747
R1920 VTAIL.n145 VTAIL.n144 9.69747
R1921 VTAIL.n382 VTAIL.n381 9.45567
R1922 VTAIL.n94 VTAIL.n93 9.45567
R1923 VTAIL.n288 VTAIL.n287 9.45567
R1924 VTAIL.n192 VTAIL.n191 9.45567
R1925 VTAIL.n381 VTAIL.n380 9.3005
R1926 VTAIL.n292 VTAIL.n291 9.3005
R1927 VTAIL.n375 VTAIL.n374 9.3005
R1928 VTAIL.n373 VTAIL.n372 9.3005
R1929 VTAIL.n296 VTAIL.n295 9.3005
R1930 VTAIL.n341 VTAIL.n340 9.3005
R1931 VTAIL.n339 VTAIL.n338 9.3005
R1932 VTAIL.n312 VTAIL.n311 9.3005
R1933 VTAIL.n333 VTAIL.n332 9.3005
R1934 VTAIL.n331 VTAIL.n330 9.3005
R1935 VTAIL.n316 VTAIL.n315 9.3005
R1936 VTAIL.n325 VTAIL.n324 9.3005
R1937 VTAIL.n323 VTAIL.n322 9.3005
R1938 VTAIL.n308 VTAIL.n307 9.3005
R1939 VTAIL.n347 VTAIL.n346 9.3005
R1940 VTAIL.n349 VTAIL.n348 9.3005
R1941 VTAIL.n304 VTAIL.n303 9.3005
R1942 VTAIL.n355 VTAIL.n354 9.3005
R1943 VTAIL.n357 VTAIL.n356 9.3005
R1944 VTAIL.n300 VTAIL.n299 9.3005
R1945 VTAIL.n364 VTAIL.n363 9.3005
R1946 VTAIL.n366 VTAIL.n365 9.3005
R1947 VTAIL.n93 VTAIL.n92 9.3005
R1948 VTAIL.n4 VTAIL.n3 9.3005
R1949 VTAIL.n87 VTAIL.n86 9.3005
R1950 VTAIL.n85 VTAIL.n84 9.3005
R1951 VTAIL.n8 VTAIL.n7 9.3005
R1952 VTAIL.n53 VTAIL.n52 9.3005
R1953 VTAIL.n51 VTAIL.n50 9.3005
R1954 VTAIL.n24 VTAIL.n23 9.3005
R1955 VTAIL.n45 VTAIL.n44 9.3005
R1956 VTAIL.n43 VTAIL.n42 9.3005
R1957 VTAIL.n28 VTAIL.n27 9.3005
R1958 VTAIL.n37 VTAIL.n36 9.3005
R1959 VTAIL.n35 VTAIL.n34 9.3005
R1960 VTAIL.n20 VTAIL.n19 9.3005
R1961 VTAIL.n59 VTAIL.n58 9.3005
R1962 VTAIL.n61 VTAIL.n60 9.3005
R1963 VTAIL.n16 VTAIL.n15 9.3005
R1964 VTAIL.n67 VTAIL.n66 9.3005
R1965 VTAIL.n69 VTAIL.n68 9.3005
R1966 VTAIL.n12 VTAIL.n11 9.3005
R1967 VTAIL.n76 VTAIL.n75 9.3005
R1968 VTAIL.n78 VTAIL.n77 9.3005
R1969 VTAIL.n254 VTAIL.n253 9.3005
R1970 VTAIL.n256 VTAIL.n255 9.3005
R1971 VTAIL.n211 VTAIL.n210 9.3005
R1972 VTAIL.n262 VTAIL.n261 9.3005
R1973 VTAIL.n264 VTAIL.n263 9.3005
R1974 VTAIL.n206 VTAIL.n205 9.3005
R1975 VTAIL.n270 VTAIL.n269 9.3005
R1976 VTAIL.n272 VTAIL.n271 9.3005
R1977 VTAIL.n287 VTAIL.n286 9.3005
R1978 VTAIL.n198 VTAIL.n197 9.3005
R1979 VTAIL.n281 VTAIL.n280 9.3005
R1980 VTAIL.n279 VTAIL.n278 9.3005
R1981 VTAIL.n202 VTAIL.n201 9.3005
R1982 VTAIL.n215 VTAIL.n214 9.3005
R1983 VTAIL.n248 VTAIL.n247 9.3005
R1984 VTAIL.n246 VTAIL.n245 9.3005
R1985 VTAIL.n219 VTAIL.n218 9.3005
R1986 VTAIL.n240 VTAIL.n239 9.3005
R1987 VTAIL.n238 VTAIL.n237 9.3005
R1988 VTAIL.n223 VTAIL.n222 9.3005
R1989 VTAIL.n232 VTAIL.n231 9.3005
R1990 VTAIL.n230 VTAIL.n229 9.3005
R1991 VTAIL.n158 VTAIL.n157 9.3005
R1992 VTAIL.n160 VTAIL.n159 9.3005
R1993 VTAIL.n115 VTAIL.n114 9.3005
R1994 VTAIL.n166 VTAIL.n165 9.3005
R1995 VTAIL.n168 VTAIL.n167 9.3005
R1996 VTAIL.n110 VTAIL.n109 9.3005
R1997 VTAIL.n174 VTAIL.n173 9.3005
R1998 VTAIL.n176 VTAIL.n175 9.3005
R1999 VTAIL.n191 VTAIL.n190 9.3005
R2000 VTAIL.n102 VTAIL.n101 9.3005
R2001 VTAIL.n185 VTAIL.n184 9.3005
R2002 VTAIL.n183 VTAIL.n182 9.3005
R2003 VTAIL.n106 VTAIL.n105 9.3005
R2004 VTAIL.n119 VTAIL.n118 9.3005
R2005 VTAIL.n152 VTAIL.n151 9.3005
R2006 VTAIL.n150 VTAIL.n149 9.3005
R2007 VTAIL.n123 VTAIL.n122 9.3005
R2008 VTAIL.n144 VTAIL.n143 9.3005
R2009 VTAIL.n142 VTAIL.n141 9.3005
R2010 VTAIL.n127 VTAIL.n126 9.3005
R2011 VTAIL.n136 VTAIL.n135 9.3005
R2012 VTAIL.n134 VTAIL.n133 9.3005
R2013 VTAIL.n337 VTAIL.n312 8.92171
R2014 VTAIL.n350 VTAIL.n304 8.92171
R2015 VTAIL.n49 VTAIL.n24 8.92171
R2016 VTAIL.n62 VTAIL.n16 8.92171
R2017 VTAIL.n257 VTAIL.n211 8.92171
R2018 VTAIL.n244 VTAIL.n219 8.92171
R2019 VTAIL.n161 VTAIL.n115 8.92171
R2020 VTAIL.n148 VTAIL.n123 8.92171
R2021 VTAIL.n338 VTAIL.n310 8.14595
R2022 VTAIL.n349 VTAIL.n306 8.14595
R2023 VTAIL.n50 VTAIL.n22 8.14595
R2024 VTAIL.n61 VTAIL.n18 8.14595
R2025 VTAIL.n256 VTAIL.n213 8.14595
R2026 VTAIL.n245 VTAIL.n217 8.14595
R2027 VTAIL.n160 VTAIL.n117 8.14595
R2028 VTAIL.n149 VTAIL.n121 8.14595
R2029 VTAIL.n342 VTAIL.n341 7.3702
R2030 VTAIL.n346 VTAIL.n345 7.3702
R2031 VTAIL.n54 VTAIL.n53 7.3702
R2032 VTAIL.n58 VTAIL.n57 7.3702
R2033 VTAIL.n253 VTAIL.n252 7.3702
R2034 VTAIL.n249 VTAIL.n248 7.3702
R2035 VTAIL.n157 VTAIL.n156 7.3702
R2036 VTAIL.n153 VTAIL.n152 7.3702
R2037 VTAIL.n342 VTAIL.n308 6.59444
R2038 VTAIL.n345 VTAIL.n308 6.59444
R2039 VTAIL.n54 VTAIL.n20 6.59444
R2040 VTAIL.n57 VTAIL.n20 6.59444
R2041 VTAIL.n252 VTAIL.n215 6.59444
R2042 VTAIL.n249 VTAIL.n215 6.59444
R2043 VTAIL.n156 VTAIL.n119 6.59444
R2044 VTAIL.n153 VTAIL.n119 6.59444
R2045 VTAIL.n341 VTAIL.n310 5.81868
R2046 VTAIL.n346 VTAIL.n306 5.81868
R2047 VTAIL.n53 VTAIL.n22 5.81868
R2048 VTAIL.n58 VTAIL.n18 5.81868
R2049 VTAIL.n253 VTAIL.n213 5.81868
R2050 VTAIL.n248 VTAIL.n217 5.81868
R2051 VTAIL.n157 VTAIL.n117 5.81868
R2052 VTAIL.n152 VTAIL.n121 5.81868
R2053 VTAIL.n338 VTAIL.n337 5.04292
R2054 VTAIL.n350 VTAIL.n349 5.04292
R2055 VTAIL.n50 VTAIL.n49 5.04292
R2056 VTAIL.n62 VTAIL.n61 5.04292
R2057 VTAIL.n257 VTAIL.n256 5.04292
R2058 VTAIL.n245 VTAIL.n244 5.04292
R2059 VTAIL.n161 VTAIL.n160 5.04292
R2060 VTAIL.n149 VTAIL.n148 5.04292
R2061 VTAIL.n334 VTAIL.n312 4.26717
R2062 VTAIL.n353 VTAIL.n304 4.26717
R2063 VTAIL.n382 VTAIL.n290 4.26717
R2064 VTAIL.n46 VTAIL.n24 4.26717
R2065 VTAIL.n65 VTAIL.n16 4.26717
R2066 VTAIL.n94 VTAIL.n2 4.26717
R2067 VTAIL.n288 VTAIL.n196 4.26717
R2068 VTAIL.n260 VTAIL.n211 4.26717
R2069 VTAIL.n241 VTAIL.n219 4.26717
R2070 VTAIL.n192 VTAIL.n100 4.26717
R2071 VTAIL.n164 VTAIL.n115 4.26717
R2072 VTAIL.n145 VTAIL.n123 4.26717
R2073 VTAIL.n323 VTAIL.n319 3.70982
R2074 VTAIL.n35 VTAIL.n31 3.70982
R2075 VTAIL.n230 VTAIL.n226 3.70982
R2076 VTAIL.n134 VTAIL.n130 3.70982
R2077 VTAIL.n333 VTAIL.n314 3.49141
R2078 VTAIL.n354 VTAIL.n302 3.49141
R2079 VTAIL.n380 VTAIL.n379 3.49141
R2080 VTAIL.n45 VTAIL.n26 3.49141
R2081 VTAIL.n66 VTAIL.n14 3.49141
R2082 VTAIL.n92 VTAIL.n91 3.49141
R2083 VTAIL.n286 VTAIL.n285 3.49141
R2084 VTAIL.n261 VTAIL.n209 3.49141
R2085 VTAIL.n240 VTAIL.n221 3.49141
R2086 VTAIL.n190 VTAIL.n189 3.49141
R2087 VTAIL.n165 VTAIL.n113 3.49141
R2088 VTAIL.n144 VTAIL.n125 3.49141
R2089 VTAIL.n330 VTAIL.n329 2.71565
R2090 VTAIL.n358 VTAIL.n357 2.71565
R2091 VTAIL.n376 VTAIL.n292 2.71565
R2092 VTAIL.n42 VTAIL.n41 2.71565
R2093 VTAIL.n70 VTAIL.n69 2.71565
R2094 VTAIL.n88 VTAIL.n4 2.71565
R2095 VTAIL.n282 VTAIL.n198 2.71565
R2096 VTAIL.n265 VTAIL.n264 2.71565
R2097 VTAIL.n237 VTAIL.n236 2.71565
R2098 VTAIL.n186 VTAIL.n102 2.71565
R2099 VTAIL.n169 VTAIL.n168 2.71565
R2100 VTAIL.n141 VTAIL.n140 2.71565
R2101 VTAIL.n193 VTAIL.n99 2.67291
R2102 VTAIL.n289 VTAIL.n195 2.67291
R2103 VTAIL.n97 VTAIL.n95 2.67291
R2104 VTAIL VTAIL.n383 1.94662
R2105 VTAIL.n0 VTAIL.t2 1.94458
R2106 VTAIL.n0 VTAIL.t4 1.94458
R2107 VTAIL.n96 VTAIL.t5 1.94458
R2108 VTAIL.n96 VTAIL.t10 1.94458
R2109 VTAIL.n194 VTAIL.t7 1.94458
R2110 VTAIL.n194 VTAIL.t9 1.94458
R2111 VTAIL.n98 VTAIL.t0 1.94458
R2112 VTAIL.n98 VTAIL.t3 1.94458
R2113 VTAIL.n326 VTAIL.n316 1.93989
R2114 VTAIL.n362 VTAIL.n300 1.93989
R2115 VTAIL.n375 VTAIL.n294 1.93989
R2116 VTAIL.n38 VTAIL.n28 1.93989
R2117 VTAIL.n74 VTAIL.n12 1.93989
R2118 VTAIL.n87 VTAIL.n6 1.93989
R2119 VTAIL.n281 VTAIL.n200 1.93989
R2120 VTAIL.n268 VTAIL.n206 1.93989
R2121 VTAIL.n233 VTAIL.n223 1.93989
R2122 VTAIL.n185 VTAIL.n104 1.93989
R2123 VTAIL.n172 VTAIL.n110 1.93989
R2124 VTAIL.n137 VTAIL.n127 1.93989
R2125 VTAIL.n195 VTAIL.n193 1.80653
R2126 VTAIL.n95 VTAIL.n1 1.80653
R2127 VTAIL.n325 VTAIL.n318 1.16414
R2128 VTAIL.n363 VTAIL.n298 1.16414
R2129 VTAIL.n372 VTAIL.n371 1.16414
R2130 VTAIL.n37 VTAIL.n30 1.16414
R2131 VTAIL.n75 VTAIL.n10 1.16414
R2132 VTAIL.n84 VTAIL.n83 1.16414
R2133 VTAIL.n278 VTAIL.n277 1.16414
R2134 VTAIL.n269 VTAIL.n204 1.16414
R2135 VTAIL.n232 VTAIL.n225 1.16414
R2136 VTAIL.n182 VTAIL.n181 1.16414
R2137 VTAIL.n173 VTAIL.n108 1.16414
R2138 VTAIL.n136 VTAIL.n129 1.16414
R2139 VTAIL VTAIL.n1 0.726793
R2140 VTAIL.n322 VTAIL.n321 0.388379
R2141 VTAIL.n367 VTAIL.n366 0.388379
R2142 VTAIL.n368 VTAIL.n296 0.388379
R2143 VTAIL.n34 VTAIL.n33 0.388379
R2144 VTAIL.n79 VTAIL.n78 0.388379
R2145 VTAIL.n80 VTAIL.n8 0.388379
R2146 VTAIL.n274 VTAIL.n202 0.388379
R2147 VTAIL.n273 VTAIL.n272 0.388379
R2148 VTAIL.n229 VTAIL.n228 0.388379
R2149 VTAIL.n178 VTAIL.n106 0.388379
R2150 VTAIL.n177 VTAIL.n176 0.388379
R2151 VTAIL.n133 VTAIL.n132 0.388379
R2152 VTAIL.n324 VTAIL.n323 0.155672
R2153 VTAIL.n324 VTAIL.n315 0.155672
R2154 VTAIL.n331 VTAIL.n315 0.155672
R2155 VTAIL.n332 VTAIL.n331 0.155672
R2156 VTAIL.n332 VTAIL.n311 0.155672
R2157 VTAIL.n339 VTAIL.n311 0.155672
R2158 VTAIL.n340 VTAIL.n339 0.155672
R2159 VTAIL.n340 VTAIL.n307 0.155672
R2160 VTAIL.n347 VTAIL.n307 0.155672
R2161 VTAIL.n348 VTAIL.n347 0.155672
R2162 VTAIL.n348 VTAIL.n303 0.155672
R2163 VTAIL.n355 VTAIL.n303 0.155672
R2164 VTAIL.n356 VTAIL.n355 0.155672
R2165 VTAIL.n356 VTAIL.n299 0.155672
R2166 VTAIL.n364 VTAIL.n299 0.155672
R2167 VTAIL.n365 VTAIL.n364 0.155672
R2168 VTAIL.n365 VTAIL.n295 0.155672
R2169 VTAIL.n373 VTAIL.n295 0.155672
R2170 VTAIL.n374 VTAIL.n373 0.155672
R2171 VTAIL.n374 VTAIL.n291 0.155672
R2172 VTAIL.n381 VTAIL.n291 0.155672
R2173 VTAIL.n36 VTAIL.n35 0.155672
R2174 VTAIL.n36 VTAIL.n27 0.155672
R2175 VTAIL.n43 VTAIL.n27 0.155672
R2176 VTAIL.n44 VTAIL.n43 0.155672
R2177 VTAIL.n44 VTAIL.n23 0.155672
R2178 VTAIL.n51 VTAIL.n23 0.155672
R2179 VTAIL.n52 VTAIL.n51 0.155672
R2180 VTAIL.n52 VTAIL.n19 0.155672
R2181 VTAIL.n59 VTAIL.n19 0.155672
R2182 VTAIL.n60 VTAIL.n59 0.155672
R2183 VTAIL.n60 VTAIL.n15 0.155672
R2184 VTAIL.n67 VTAIL.n15 0.155672
R2185 VTAIL.n68 VTAIL.n67 0.155672
R2186 VTAIL.n68 VTAIL.n11 0.155672
R2187 VTAIL.n76 VTAIL.n11 0.155672
R2188 VTAIL.n77 VTAIL.n76 0.155672
R2189 VTAIL.n77 VTAIL.n7 0.155672
R2190 VTAIL.n85 VTAIL.n7 0.155672
R2191 VTAIL.n86 VTAIL.n85 0.155672
R2192 VTAIL.n86 VTAIL.n3 0.155672
R2193 VTAIL.n93 VTAIL.n3 0.155672
R2194 VTAIL.n287 VTAIL.n197 0.155672
R2195 VTAIL.n280 VTAIL.n197 0.155672
R2196 VTAIL.n280 VTAIL.n279 0.155672
R2197 VTAIL.n279 VTAIL.n201 0.155672
R2198 VTAIL.n271 VTAIL.n201 0.155672
R2199 VTAIL.n271 VTAIL.n270 0.155672
R2200 VTAIL.n270 VTAIL.n205 0.155672
R2201 VTAIL.n263 VTAIL.n205 0.155672
R2202 VTAIL.n263 VTAIL.n262 0.155672
R2203 VTAIL.n262 VTAIL.n210 0.155672
R2204 VTAIL.n255 VTAIL.n210 0.155672
R2205 VTAIL.n255 VTAIL.n254 0.155672
R2206 VTAIL.n254 VTAIL.n214 0.155672
R2207 VTAIL.n247 VTAIL.n214 0.155672
R2208 VTAIL.n247 VTAIL.n246 0.155672
R2209 VTAIL.n246 VTAIL.n218 0.155672
R2210 VTAIL.n239 VTAIL.n218 0.155672
R2211 VTAIL.n239 VTAIL.n238 0.155672
R2212 VTAIL.n238 VTAIL.n222 0.155672
R2213 VTAIL.n231 VTAIL.n222 0.155672
R2214 VTAIL.n231 VTAIL.n230 0.155672
R2215 VTAIL.n191 VTAIL.n101 0.155672
R2216 VTAIL.n184 VTAIL.n101 0.155672
R2217 VTAIL.n184 VTAIL.n183 0.155672
R2218 VTAIL.n183 VTAIL.n105 0.155672
R2219 VTAIL.n175 VTAIL.n105 0.155672
R2220 VTAIL.n175 VTAIL.n174 0.155672
R2221 VTAIL.n174 VTAIL.n109 0.155672
R2222 VTAIL.n167 VTAIL.n109 0.155672
R2223 VTAIL.n167 VTAIL.n166 0.155672
R2224 VTAIL.n166 VTAIL.n114 0.155672
R2225 VTAIL.n159 VTAIL.n114 0.155672
R2226 VTAIL.n159 VTAIL.n158 0.155672
R2227 VTAIL.n158 VTAIL.n118 0.155672
R2228 VTAIL.n151 VTAIL.n118 0.155672
R2229 VTAIL.n151 VTAIL.n150 0.155672
R2230 VTAIL.n150 VTAIL.n122 0.155672
R2231 VTAIL.n143 VTAIL.n122 0.155672
R2232 VTAIL.n143 VTAIL.n142 0.155672
R2233 VTAIL.n142 VTAIL.n126 0.155672
R2234 VTAIL.n135 VTAIL.n126 0.155672
R2235 VTAIL.n135 VTAIL.n134 0.155672
R2236 VN.n4 VN.t2 179.55
R2237 VN.n20 VN.t1 179.55
R2238 VN.n29 VN.n16 161.3
R2239 VN.n28 VN.n27 161.3
R2240 VN.n26 VN.n17 161.3
R2241 VN.n25 VN.n24 161.3
R2242 VN.n23 VN.n18 161.3
R2243 VN.n22 VN.n21 161.3
R2244 VN.n13 VN.n0 161.3
R2245 VN.n12 VN.n11 161.3
R2246 VN.n10 VN.n1 161.3
R2247 VN.n9 VN.n8 161.3
R2248 VN.n7 VN.n2 161.3
R2249 VN.n6 VN.n5 161.3
R2250 VN.n3 VN.t4 145.47
R2251 VN.n14 VN.t3 145.47
R2252 VN.n19 VN.t0 145.47
R2253 VN.n30 VN.t5 145.47
R2254 VN.n15 VN.n14 105.99
R2255 VN.n31 VN.n30 105.99
R2256 VN VN.n31 53.18
R2257 VN.n20 VN.n19 49.0286
R2258 VN.n4 VN.n3 49.0286
R2259 VN.n8 VN.n1 45.4209
R2260 VN.n24 VN.n17 45.4209
R2261 VN.n8 VN.n7 35.7332
R2262 VN.n24 VN.n23 35.7332
R2263 VN.n6 VN.n3 24.5923
R2264 VN.n7 VN.n6 24.5923
R2265 VN.n12 VN.n1 24.5923
R2266 VN.n13 VN.n12 24.5923
R2267 VN.n23 VN.n22 24.5923
R2268 VN.n22 VN.n19 24.5923
R2269 VN.n29 VN.n28 24.5923
R2270 VN.n28 VN.n17 24.5923
R2271 VN.n21 VN.n20 4.96469
R2272 VN.n5 VN.n4 4.96469
R2273 VN.n14 VN.n13 4.91887
R2274 VN.n30 VN.n29 4.91887
R2275 VN.n31 VN.n16 0.278335
R2276 VN.n15 VN.n0 0.278335
R2277 VN.n27 VN.n16 0.189894
R2278 VN.n27 VN.n26 0.189894
R2279 VN.n26 VN.n25 0.189894
R2280 VN.n25 VN.n18 0.189894
R2281 VN.n21 VN.n18 0.189894
R2282 VN.n5 VN.n2 0.189894
R2283 VN.n9 VN.n2 0.189894
R2284 VN.n10 VN.n9 0.189894
R2285 VN.n11 VN.n10 0.189894
R2286 VN.n11 VN.n0 0.189894
R2287 VN VN.n15 0.153485
R2288 VDD2.n183 VDD2.n95 756.745
R2289 VDD2.n88 VDD2.n0 756.745
R2290 VDD2.n184 VDD2.n183 585
R2291 VDD2.n182 VDD2.n181 585
R2292 VDD2.n99 VDD2.n98 585
R2293 VDD2.n176 VDD2.n175 585
R2294 VDD2.n174 VDD2.n173 585
R2295 VDD2.n172 VDD2.n102 585
R2296 VDD2.n106 VDD2.n103 585
R2297 VDD2.n167 VDD2.n166 585
R2298 VDD2.n165 VDD2.n164 585
R2299 VDD2.n108 VDD2.n107 585
R2300 VDD2.n159 VDD2.n158 585
R2301 VDD2.n157 VDD2.n156 585
R2302 VDD2.n112 VDD2.n111 585
R2303 VDD2.n151 VDD2.n150 585
R2304 VDD2.n149 VDD2.n148 585
R2305 VDD2.n116 VDD2.n115 585
R2306 VDD2.n143 VDD2.n142 585
R2307 VDD2.n141 VDD2.n140 585
R2308 VDD2.n120 VDD2.n119 585
R2309 VDD2.n135 VDD2.n134 585
R2310 VDD2.n133 VDD2.n132 585
R2311 VDD2.n124 VDD2.n123 585
R2312 VDD2.n127 VDD2.n126 585
R2313 VDD2.n31 VDD2.n30 585
R2314 VDD2.n28 VDD2.n27 585
R2315 VDD2.n37 VDD2.n36 585
R2316 VDD2.n39 VDD2.n38 585
R2317 VDD2.n24 VDD2.n23 585
R2318 VDD2.n45 VDD2.n44 585
R2319 VDD2.n47 VDD2.n46 585
R2320 VDD2.n20 VDD2.n19 585
R2321 VDD2.n53 VDD2.n52 585
R2322 VDD2.n55 VDD2.n54 585
R2323 VDD2.n16 VDD2.n15 585
R2324 VDD2.n61 VDD2.n60 585
R2325 VDD2.n63 VDD2.n62 585
R2326 VDD2.n12 VDD2.n11 585
R2327 VDD2.n69 VDD2.n68 585
R2328 VDD2.n72 VDD2.n71 585
R2329 VDD2.n70 VDD2.n8 585
R2330 VDD2.n77 VDD2.n7 585
R2331 VDD2.n79 VDD2.n78 585
R2332 VDD2.n81 VDD2.n80 585
R2333 VDD2.n4 VDD2.n3 585
R2334 VDD2.n87 VDD2.n86 585
R2335 VDD2.n89 VDD2.n88 585
R2336 VDD2.t0 VDD2.n125 327.466
R2337 VDD2.t3 VDD2.n29 327.466
R2338 VDD2.n183 VDD2.n182 171.744
R2339 VDD2.n182 VDD2.n98 171.744
R2340 VDD2.n175 VDD2.n98 171.744
R2341 VDD2.n175 VDD2.n174 171.744
R2342 VDD2.n174 VDD2.n102 171.744
R2343 VDD2.n106 VDD2.n102 171.744
R2344 VDD2.n166 VDD2.n106 171.744
R2345 VDD2.n166 VDD2.n165 171.744
R2346 VDD2.n165 VDD2.n107 171.744
R2347 VDD2.n158 VDD2.n107 171.744
R2348 VDD2.n158 VDD2.n157 171.744
R2349 VDD2.n157 VDD2.n111 171.744
R2350 VDD2.n150 VDD2.n111 171.744
R2351 VDD2.n150 VDD2.n149 171.744
R2352 VDD2.n149 VDD2.n115 171.744
R2353 VDD2.n142 VDD2.n115 171.744
R2354 VDD2.n142 VDD2.n141 171.744
R2355 VDD2.n141 VDD2.n119 171.744
R2356 VDD2.n134 VDD2.n119 171.744
R2357 VDD2.n134 VDD2.n133 171.744
R2358 VDD2.n133 VDD2.n123 171.744
R2359 VDD2.n126 VDD2.n123 171.744
R2360 VDD2.n30 VDD2.n27 171.744
R2361 VDD2.n37 VDD2.n27 171.744
R2362 VDD2.n38 VDD2.n37 171.744
R2363 VDD2.n38 VDD2.n23 171.744
R2364 VDD2.n45 VDD2.n23 171.744
R2365 VDD2.n46 VDD2.n45 171.744
R2366 VDD2.n46 VDD2.n19 171.744
R2367 VDD2.n53 VDD2.n19 171.744
R2368 VDD2.n54 VDD2.n53 171.744
R2369 VDD2.n54 VDD2.n15 171.744
R2370 VDD2.n61 VDD2.n15 171.744
R2371 VDD2.n62 VDD2.n61 171.744
R2372 VDD2.n62 VDD2.n11 171.744
R2373 VDD2.n69 VDD2.n11 171.744
R2374 VDD2.n71 VDD2.n69 171.744
R2375 VDD2.n71 VDD2.n70 171.744
R2376 VDD2.n70 VDD2.n7 171.744
R2377 VDD2.n79 VDD2.n7 171.744
R2378 VDD2.n80 VDD2.n79 171.744
R2379 VDD2.n80 VDD2.n3 171.744
R2380 VDD2.n87 VDD2.n3 171.744
R2381 VDD2.n88 VDD2.n87 171.744
R2382 VDD2.n126 VDD2.t0 85.8723
R2383 VDD2.n30 VDD2.t3 85.8723
R2384 VDD2.n94 VDD2.n93 68.4531
R2385 VDD2 VDD2.n189 68.4503
R2386 VDD2.n94 VDD2.n92 49.2616
R2387 VDD2.n188 VDD2.n187 47.3126
R2388 VDD2.n188 VDD2.n94 46.8144
R2389 VDD2.n127 VDD2.n125 16.3895
R2390 VDD2.n31 VDD2.n29 16.3895
R2391 VDD2.n173 VDD2.n172 13.1884
R2392 VDD2.n78 VDD2.n77 13.1884
R2393 VDD2.n176 VDD2.n101 12.8005
R2394 VDD2.n171 VDD2.n103 12.8005
R2395 VDD2.n128 VDD2.n124 12.8005
R2396 VDD2.n32 VDD2.n28 12.8005
R2397 VDD2.n76 VDD2.n8 12.8005
R2398 VDD2.n81 VDD2.n6 12.8005
R2399 VDD2.n177 VDD2.n99 12.0247
R2400 VDD2.n168 VDD2.n167 12.0247
R2401 VDD2.n132 VDD2.n131 12.0247
R2402 VDD2.n36 VDD2.n35 12.0247
R2403 VDD2.n73 VDD2.n72 12.0247
R2404 VDD2.n82 VDD2.n4 12.0247
R2405 VDD2.n181 VDD2.n180 11.249
R2406 VDD2.n164 VDD2.n105 11.249
R2407 VDD2.n135 VDD2.n122 11.249
R2408 VDD2.n39 VDD2.n26 11.249
R2409 VDD2.n68 VDD2.n10 11.249
R2410 VDD2.n86 VDD2.n85 11.249
R2411 VDD2.n184 VDD2.n97 10.4732
R2412 VDD2.n163 VDD2.n108 10.4732
R2413 VDD2.n136 VDD2.n120 10.4732
R2414 VDD2.n40 VDD2.n24 10.4732
R2415 VDD2.n67 VDD2.n12 10.4732
R2416 VDD2.n89 VDD2.n2 10.4732
R2417 VDD2.n185 VDD2.n95 9.69747
R2418 VDD2.n160 VDD2.n159 9.69747
R2419 VDD2.n140 VDD2.n139 9.69747
R2420 VDD2.n44 VDD2.n43 9.69747
R2421 VDD2.n64 VDD2.n63 9.69747
R2422 VDD2.n90 VDD2.n0 9.69747
R2423 VDD2.n187 VDD2.n186 9.45567
R2424 VDD2.n92 VDD2.n91 9.45567
R2425 VDD2.n153 VDD2.n152 9.3005
R2426 VDD2.n155 VDD2.n154 9.3005
R2427 VDD2.n110 VDD2.n109 9.3005
R2428 VDD2.n161 VDD2.n160 9.3005
R2429 VDD2.n163 VDD2.n162 9.3005
R2430 VDD2.n105 VDD2.n104 9.3005
R2431 VDD2.n169 VDD2.n168 9.3005
R2432 VDD2.n171 VDD2.n170 9.3005
R2433 VDD2.n186 VDD2.n185 9.3005
R2434 VDD2.n97 VDD2.n96 9.3005
R2435 VDD2.n180 VDD2.n179 9.3005
R2436 VDD2.n178 VDD2.n177 9.3005
R2437 VDD2.n101 VDD2.n100 9.3005
R2438 VDD2.n114 VDD2.n113 9.3005
R2439 VDD2.n147 VDD2.n146 9.3005
R2440 VDD2.n145 VDD2.n144 9.3005
R2441 VDD2.n118 VDD2.n117 9.3005
R2442 VDD2.n139 VDD2.n138 9.3005
R2443 VDD2.n137 VDD2.n136 9.3005
R2444 VDD2.n122 VDD2.n121 9.3005
R2445 VDD2.n131 VDD2.n130 9.3005
R2446 VDD2.n129 VDD2.n128 9.3005
R2447 VDD2.n91 VDD2.n90 9.3005
R2448 VDD2.n2 VDD2.n1 9.3005
R2449 VDD2.n85 VDD2.n84 9.3005
R2450 VDD2.n83 VDD2.n82 9.3005
R2451 VDD2.n6 VDD2.n5 9.3005
R2452 VDD2.n51 VDD2.n50 9.3005
R2453 VDD2.n49 VDD2.n48 9.3005
R2454 VDD2.n22 VDD2.n21 9.3005
R2455 VDD2.n43 VDD2.n42 9.3005
R2456 VDD2.n41 VDD2.n40 9.3005
R2457 VDD2.n26 VDD2.n25 9.3005
R2458 VDD2.n35 VDD2.n34 9.3005
R2459 VDD2.n33 VDD2.n32 9.3005
R2460 VDD2.n18 VDD2.n17 9.3005
R2461 VDD2.n57 VDD2.n56 9.3005
R2462 VDD2.n59 VDD2.n58 9.3005
R2463 VDD2.n14 VDD2.n13 9.3005
R2464 VDD2.n65 VDD2.n64 9.3005
R2465 VDD2.n67 VDD2.n66 9.3005
R2466 VDD2.n10 VDD2.n9 9.3005
R2467 VDD2.n74 VDD2.n73 9.3005
R2468 VDD2.n76 VDD2.n75 9.3005
R2469 VDD2.n156 VDD2.n110 8.92171
R2470 VDD2.n143 VDD2.n118 8.92171
R2471 VDD2.n47 VDD2.n22 8.92171
R2472 VDD2.n60 VDD2.n14 8.92171
R2473 VDD2.n155 VDD2.n112 8.14595
R2474 VDD2.n144 VDD2.n116 8.14595
R2475 VDD2.n48 VDD2.n20 8.14595
R2476 VDD2.n59 VDD2.n16 8.14595
R2477 VDD2.n152 VDD2.n151 7.3702
R2478 VDD2.n148 VDD2.n147 7.3702
R2479 VDD2.n52 VDD2.n51 7.3702
R2480 VDD2.n56 VDD2.n55 7.3702
R2481 VDD2.n151 VDD2.n114 6.59444
R2482 VDD2.n148 VDD2.n114 6.59444
R2483 VDD2.n52 VDD2.n18 6.59444
R2484 VDD2.n55 VDD2.n18 6.59444
R2485 VDD2.n152 VDD2.n112 5.81868
R2486 VDD2.n147 VDD2.n116 5.81868
R2487 VDD2.n51 VDD2.n20 5.81868
R2488 VDD2.n56 VDD2.n16 5.81868
R2489 VDD2.n156 VDD2.n155 5.04292
R2490 VDD2.n144 VDD2.n143 5.04292
R2491 VDD2.n48 VDD2.n47 5.04292
R2492 VDD2.n60 VDD2.n59 5.04292
R2493 VDD2.n187 VDD2.n95 4.26717
R2494 VDD2.n159 VDD2.n110 4.26717
R2495 VDD2.n140 VDD2.n118 4.26717
R2496 VDD2.n44 VDD2.n22 4.26717
R2497 VDD2.n63 VDD2.n14 4.26717
R2498 VDD2.n92 VDD2.n0 4.26717
R2499 VDD2.n129 VDD2.n125 3.70982
R2500 VDD2.n33 VDD2.n29 3.70982
R2501 VDD2.n185 VDD2.n184 3.49141
R2502 VDD2.n160 VDD2.n108 3.49141
R2503 VDD2.n139 VDD2.n120 3.49141
R2504 VDD2.n43 VDD2.n24 3.49141
R2505 VDD2.n64 VDD2.n12 3.49141
R2506 VDD2.n90 VDD2.n89 3.49141
R2507 VDD2.n181 VDD2.n97 2.71565
R2508 VDD2.n164 VDD2.n163 2.71565
R2509 VDD2.n136 VDD2.n135 2.71565
R2510 VDD2.n40 VDD2.n39 2.71565
R2511 VDD2.n68 VDD2.n67 2.71565
R2512 VDD2.n86 VDD2.n2 2.71565
R2513 VDD2 VDD2.n188 2.063
R2514 VDD2.n189 VDD2.t5 1.94458
R2515 VDD2.n189 VDD2.t4 1.94458
R2516 VDD2.n93 VDD2.t1 1.94458
R2517 VDD2.n93 VDD2.t2 1.94458
R2518 VDD2.n180 VDD2.n99 1.93989
R2519 VDD2.n167 VDD2.n105 1.93989
R2520 VDD2.n132 VDD2.n122 1.93989
R2521 VDD2.n36 VDD2.n26 1.93989
R2522 VDD2.n72 VDD2.n10 1.93989
R2523 VDD2.n85 VDD2.n4 1.93989
R2524 VDD2.n177 VDD2.n176 1.16414
R2525 VDD2.n168 VDD2.n103 1.16414
R2526 VDD2.n131 VDD2.n124 1.16414
R2527 VDD2.n35 VDD2.n28 1.16414
R2528 VDD2.n73 VDD2.n8 1.16414
R2529 VDD2.n82 VDD2.n81 1.16414
R2530 VDD2.n173 VDD2.n101 0.388379
R2531 VDD2.n172 VDD2.n171 0.388379
R2532 VDD2.n128 VDD2.n127 0.388379
R2533 VDD2.n32 VDD2.n31 0.388379
R2534 VDD2.n77 VDD2.n76 0.388379
R2535 VDD2.n78 VDD2.n6 0.388379
R2536 VDD2.n186 VDD2.n96 0.155672
R2537 VDD2.n179 VDD2.n96 0.155672
R2538 VDD2.n179 VDD2.n178 0.155672
R2539 VDD2.n178 VDD2.n100 0.155672
R2540 VDD2.n170 VDD2.n100 0.155672
R2541 VDD2.n170 VDD2.n169 0.155672
R2542 VDD2.n169 VDD2.n104 0.155672
R2543 VDD2.n162 VDD2.n104 0.155672
R2544 VDD2.n162 VDD2.n161 0.155672
R2545 VDD2.n161 VDD2.n109 0.155672
R2546 VDD2.n154 VDD2.n109 0.155672
R2547 VDD2.n154 VDD2.n153 0.155672
R2548 VDD2.n153 VDD2.n113 0.155672
R2549 VDD2.n146 VDD2.n113 0.155672
R2550 VDD2.n146 VDD2.n145 0.155672
R2551 VDD2.n145 VDD2.n117 0.155672
R2552 VDD2.n138 VDD2.n117 0.155672
R2553 VDD2.n138 VDD2.n137 0.155672
R2554 VDD2.n137 VDD2.n121 0.155672
R2555 VDD2.n130 VDD2.n121 0.155672
R2556 VDD2.n130 VDD2.n129 0.155672
R2557 VDD2.n34 VDD2.n33 0.155672
R2558 VDD2.n34 VDD2.n25 0.155672
R2559 VDD2.n41 VDD2.n25 0.155672
R2560 VDD2.n42 VDD2.n41 0.155672
R2561 VDD2.n42 VDD2.n21 0.155672
R2562 VDD2.n49 VDD2.n21 0.155672
R2563 VDD2.n50 VDD2.n49 0.155672
R2564 VDD2.n50 VDD2.n17 0.155672
R2565 VDD2.n57 VDD2.n17 0.155672
R2566 VDD2.n58 VDD2.n57 0.155672
R2567 VDD2.n58 VDD2.n13 0.155672
R2568 VDD2.n65 VDD2.n13 0.155672
R2569 VDD2.n66 VDD2.n65 0.155672
R2570 VDD2.n66 VDD2.n9 0.155672
R2571 VDD2.n74 VDD2.n9 0.155672
R2572 VDD2.n75 VDD2.n74 0.155672
R2573 VDD2.n75 VDD2.n5 0.155672
R2574 VDD2.n83 VDD2.n5 0.155672
R2575 VDD2.n84 VDD2.n83 0.155672
R2576 VDD2.n84 VDD2.n1 0.155672
R2577 VDD2.n91 VDD2.n1 0.155672
C0 VN VTAIL 9.315289f
C1 B VDD1 2.51202f
C2 w_n3450_n4312# VN 6.65814f
C3 B VDD2 2.59019f
C4 VDD1 VN 0.151177f
C5 VDD2 VN 9.33115f
C6 w_n3450_n4312# VTAIL 3.63843f
C7 B VP 2.0087f
C8 VDD1 VTAIL 9.43618f
C9 VP VN 7.96038f
C10 w_n3450_n4312# VDD1 2.65717f
C11 VDD2 VTAIL 9.4873f
C12 w_n3450_n4312# VDD2 2.74765f
C13 VP VTAIL 9.32963f
C14 B VN 1.26234f
C15 VDD1 VDD2 1.47287f
C16 w_n3450_n4312# VP 7.10465f
C17 VP VDD1 9.64933f
C18 B VTAIL 4.83208f
C19 VP VDD2 0.473295f
C20 w_n3450_n4312# B 11.234401f
C21 VDD2 VSUBS 2.09193f
C22 VDD1 VSUBS 2.014333f
C23 VTAIL VSUBS 1.389326f
C24 VN VSUBS 6.17375f
C25 VP VSUBS 3.233498f
C26 B VSUBS 5.205877f
C27 w_n3450_n4312# VSUBS 0.182119p
C28 VDD2.n0 VSUBS 0.027886f
C29 VDD2.n1 VSUBS 0.027158f
C30 VDD2.n2 VSUBS 0.014594f
C31 VDD2.n3 VSUBS 0.034494f
C32 VDD2.n4 VSUBS 0.015452f
C33 VDD2.n5 VSUBS 0.027158f
C34 VDD2.n6 VSUBS 0.014594f
C35 VDD2.n7 VSUBS 0.034494f
C36 VDD2.n8 VSUBS 0.015452f
C37 VDD2.n9 VSUBS 0.027158f
C38 VDD2.n10 VSUBS 0.014594f
C39 VDD2.n11 VSUBS 0.034494f
C40 VDD2.n12 VSUBS 0.015452f
C41 VDD2.n13 VSUBS 0.027158f
C42 VDD2.n14 VSUBS 0.014594f
C43 VDD2.n15 VSUBS 0.034494f
C44 VDD2.n16 VSUBS 0.015452f
C45 VDD2.n17 VSUBS 0.027158f
C46 VDD2.n18 VSUBS 0.014594f
C47 VDD2.n19 VSUBS 0.034494f
C48 VDD2.n20 VSUBS 0.015452f
C49 VDD2.n21 VSUBS 0.027158f
C50 VDD2.n22 VSUBS 0.014594f
C51 VDD2.n23 VSUBS 0.034494f
C52 VDD2.n24 VSUBS 0.015452f
C53 VDD2.n25 VSUBS 0.027158f
C54 VDD2.n26 VSUBS 0.014594f
C55 VDD2.n27 VSUBS 0.034494f
C56 VDD2.n28 VSUBS 0.015452f
C57 VDD2.n29 VSUBS 0.205221f
C58 VDD2.t3 VSUBS 0.073961f
C59 VDD2.n30 VSUBS 0.025871f
C60 VDD2.n31 VSUBS 0.021944f
C61 VDD2.n32 VSUBS 0.014594f
C62 VDD2.n33 VSUBS 1.94618f
C63 VDD2.n34 VSUBS 0.027158f
C64 VDD2.n35 VSUBS 0.014594f
C65 VDD2.n36 VSUBS 0.015452f
C66 VDD2.n37 VSUBS 0.034494f
C67 VDD2.n38 VSUBS 0.034494f
C68 VDD2.n39 VSUBS 0.015452f
C69 VDD2.n40 VSUBS 0.014594f
C70 VDD2.n41 VSUBS 0.027158f
C71 VDD2.n42 VSUBS 0.027158f
C72 VDD2.n43 VSUBS 0.014594f
C73 VDD2.n44 VSUBS 0.015452f
C74 VDD2.n45 VSUBS 0.034494f
C75 VDD2.n46 VSUBS 0.034494f
C76 VDD2.n47 VSUBS 0.015452f
C77 VDD2.n48 VSUBS 0.014594f
C78 VDD2.n49 VSUBS 0.027158f
C79 VDD2.n50 VSUBS 0.027158f
C80 VDD2.n51 VSUBS 0.014594f
C81 VDD2.n52 VSUBS 0.015452f
C82 VDD2.n53 VSUBS 0.034494f
C83 VDD2.n54 VSUBS 0.034494f
C84 VDD2.n55 VSUBS 0.015452f
C85 VDD2.n56 VSUBS 0.014594f
C86 VDD2.n57 VSUBS 0.027158f
C87 VDD2.n58 VSUBS 0.027158f
C88 VDD2.n59 VSUBS 0.014594f
C89 VDD2.n60 VSUBS 0.015452f
C90 VDD2.n61 VSUBS 0.034494f
C91 VDD2.n62 VSUBS 0.034494f
C92 VDD2.n63 VSUBS 0.015452f
C93 VDD2.n64 VSUBS 0.014594f
C94 VDD2.n65 VSUBS 0.027158f
C95 VDD2.n66 VSUBS 0.027158f
C96 VDD2.n67 VSUBS 0.014594f
C97 VDD2.n68 VSUBS 0.015452f
C98 VDD2.n69 VSUBS 0.034494f
C99 VDD2.n70 VSUBS 0.034494f
C100 VDD2.n71 VSUBS 0.034494f
C101 VDD2.n72 VSUBS 0.015452f
C102 VDD2.n73 VSUBS 0.014594f
C103 VDD2.n74 VSUBS 0.027158f
C104 VDD2.n75 VSUBS 0.027158f
C105 VDD2.n76 VSUBS 0.014594f
C106 VDD2.n77 VSUBS 0.015023f
C107 VDD2.n78 VSUBS 0.015023f
C108 VDD2.n79 VSUBS 0.034494f
C109 VDD2.n80 VSUBS 0.034494f
C110 VDD2.n81 VSUBS 0.015452f
C111 VDD2.n82 VSUBS 0.014594f
C112 VDD2.n83 VSUBS 0.027158f
C113 VDD2.n84 VSUBS 0.027158f
C114 VDD2.n85 VSUBS 0.014594f
C115 VDD2.n86 VSUBS 0.015452f
C116 VDD2.n87 VSUBS 0.034494f
C117 VDD2.n88 VSUBS 0.076846f
C118 VDD2.n89 VSUBS 0.015452f
C119 VDD2.n90 VSUBS 0.014594f
C120 VDD2.n91 VSUBS 0.059807f
C121 VDD2.n92 VSUBS 0.065796f
C122 VDD2.t1 VSUBS 0.358834f
C123 VDD2.t2 VSUBS 0.358834f
C124 VDD2.n93 VSUBS 2.95283f
C125 VDD2.n94 VSUBS 3.61913f
C126 VDD2.n95 VSUBS 0.027886f
C127 VDD2.n96 VSUBS 0.027158f
C128 VDD2.n97 VSUBS 0.014594f
C129 VDD2.n98 VSUBS 0.034494f
C130 VDD2.n99 VSUBS 0.015452f
C131 VDD2.n100 VSUBS 0.027158f
C132 VDD2.n101 VSUBS 0.014594f
C133 VDD2.n102 VSUBS 0.034494f
C134 VDD2.n103 VSUBS 0.015452f
C135 VDD2.n104 VSUBS 0.027158f
C136 VDD2.n105 VSUBS 0.014594f
C137 VDD2.n106 VSUBS 0.034494f
C138 VDD2.n107 VSUBS 0.034494f
C139 VDD2.n108 VSUBS 0.015452f
C140 VDD2.n109 VSUBS 0.027158f
C141 VDD2.n110 VSUBS 0.014594f
C142 VDD2.n111 VSUBS 0.034494f
C143 VDD2.n112 VSUBS 0.015452f
C144 VDD2.n113 VSUBS 0.027158f
C145 VDD2.n114 VSUBS 0.014594f
C146 VDD2.n115 VSUBS 0.034494f
C147 VDD2.n116 VSUBS 0.015452f
C148 VDD2.n117 VSUBS 0.027158f
C149 VDD2.n118 VSUBS 0.014594f
C150 VDD2.n119 VSUBS 0.034494f
C151 VDD2.n120 VSUBS 0.015452f
C152 VDD2.n121 VSUBS 0.027158f
C153 VDD2.n122 VSUBS 0.014594f
C154 VDD2.n123 VSUBS 0.034494f
C155 VDD2.n124 VSUBS 0.015452f
C156 VDD2.n125 VSUBS 0.205221f
C157 VDD2.t0 VSUBS 0.073961f
C158 VDD2.n126 VSUBS 0.025871f
C159 VDD2.n127 VSUBS 0.021944f
C160 VDD2.n128 VSUBS 0.014594f
C161 VDD2.n129 VSUBS 1.94618f
C162 VDD2.n130 VSUBS 0.027158f
C163 VDD2.n131 VSUBS 0.014594f
C164 VDD2.n132 VSUBS 0.015452f
C165 VDD2.n133 VSUBS 0.034494f
C166 VDD2.n134 VSUBS 0.034494f
C167 VDD2.n135 VSUBS 0.015452f
C168 VDD2.n136 VSUBS 0.014594f
C169 VDD2.n137 VSUBS 0.027158f
C170 VDD2.n138 VSUBS 0.027158f
C171 VDD2.n139 VSUBS 0.014594f
C172 VDD2.n140 VSUBS 0.015452f
C173 VDD2.n141 VSUBS 0.034494f
C174 VDD2.n142 VSUBS 0.034494f
C175 VDD2.n143 VSUBS 0.015452f
C176 VDD2.n144 VSUBS 0.014594f
C177 VDD2.n145 VSUBS 0.027158f
C178 VDD2.n146 VSUBS 0.027158f
C179 VDD2.n147 VSUBS 0.014594f
C180 VDD2.n148 VSUBS 0.015452f
C181 VDD2.n149 VSUBS 0.034494f
C182 VDD2.n150 VSUBS 0.034494f
C183 VDD2.n151 VSUBS 0.015452f
C184 VDD2.n152 VSUBS 0.014594f
C185 VDD2.n153 VSUBS 0.027158f
C186 VDD2.n154 VSUBS 0.027158f
C187 VDD2.n155 VSUBS 0.014594f
C188 VDD2.n156 VSUBS 0.015452f
C189 VDD2.n157 VSUBS 0.034494f
C190 VDD2.n158 VSUBS 0.034494f
C191 VDD2.n159 VSUBS 0.015452f
C192 VDD2.n160 VSUBS 0.014594f
C193 VDD2.n161 VSUBS 0.027158f
C194 VDD2.n162 VSUBS 0.027158f
C195 VDD2.n163 VSUBS 0.014594f
C196 VDD2.n164 VSUBS 0.015452f
C197 VDD2.n165 VSUBS 0.034494f
C198 VDD2.n166 VSUBS 0.034494f
C199 VDD2.n167 VSUBS 0.015452f
C200 VDD2.n168 VSUBS 0.014594f
C201 VDD2.n169 VSUBS 0.027158f
C202 VDD2.n170 VSUBS 0.027158f
C203 VDD2.n171 VSUBS 0.014594f
C204 VDD2.n172 VSUBS 0.015023f
C205 VDD2.n173 VSUBS 0.015023f
C206 VDD2.n174 VSUBS 0.034494f
C207 VDD2.n175 VSUBS 0.034494f
C208 VDD2.n176 VSUBS 0.015452f
C209 VDD2.n177 VSUBS 0.014594f
C210 VDD2.n178 VSUBS 0.027158f
C211 VDD2.n179 VSUBS 0.027158f
C212 VDD2.n180 VSUBS 0.014594f
C213 VDD2.n181 VSUBS 0.015452f
C214 VDD2.n182 VSUBS 0.034494f
C215 VDD2.n183 VSUBS 0.076846f
C216 VDD2.n184 VSUBS 0.015452f
C217 VDD2.n185 VSUBS 0.014594f
C218 VDD2.n186 VSUBS 0.059807f
C219 VDD2.n187 VSUBS 0.057033f
C220 VDD2.n188 VSUBS 3.22352f
C221 VDD2.t5 VSUBS 0.358834f
C222 VDD2.t4 VSUBS 0.358834f
C223 VDD2.n189 VSUBS 2.95278f
C224 VN.n0 VSUBS 0.035451f
C225 VN.t3 VSUBS 3.42071f
C226 VN.n1 VSUBS 0.051447f
C227 VN.n2 VSUBS 0.026891f
C228 VN.t4 VSUBS 3.42071f
C229 VN.n3 VSUBS 1.2833f
C230 VN.t2 VSUBS 3.67999f
C231 VN.n4 VSUBS 1.23004f
C232 VN.n5 VSUBS 0.281341f
C233 VN.n6 VSUBS 0.049867f
C234 VN.n7 VSUBS 0.054012f
C235 VN.n8 VSUBS 0.022588f
C236 VN.n9 VSUBS 0.026891f
C237 VN.n10 VSUBS 0.026891f
C238 VN.n11 VSUBS 0.026891f
C239 VN.n12 VSUBS 0.049867f
C240 VN.n13 VSUBS 0.030172f
C241 VN.n14 VSUBS 1.27624f
C242 VN.n15 VSUBS 0.048626f
C243 VN.n16 VSUBS 0.035451f
C244 VN.t5 VSUBS 3.42071f
C245 VN.n17 VSUBS 0.051447f
C246 VN.n18 VSUBS 0.026891f
C247 VN.t0 VSUBS 3.42071f
C248 VN.n19 VSUBS 1.2833f
C249 VN.t1 VSUBS 3.67999f
C250 VN.n20 VSUBS 1.23004f
C251 VN.n21 VSUBS 0.281341f
C252 VN.n22 VSUBS 0.049867f
C253 VN.n23 VSUBS 0.054012f
C254 VN.n24 VSUBS 0.022588f
C255 VN.n25 VSUBS 0.026891f
C256 VN.n26 VSUBS 0.026891f
C257 VN.n27 VSUBS 0.026891f
C258 VN.n28 VSUBS 0.049867f
C259 VN.n29 VSUBS 0.030172f
C260 VN.n30 VSUBS 1.27624f
C261 VN.n31 VSUBS 1.64296f
C262 VTAIL.t2 VSUBS 0.367768f
C263 VTAIL.t4 VSUBS 0.367768f
C264 VTAIL.n0 VSUBS 2.84058f
C265 VTAIL.n1 VSUBS 0.918901f
C266 VTAIL.n2 VSUBS 0.02858f
C267 VTAIL.n3 VSUBS 0.027834f
C268 VTAIL.n4 VSUBS 0.014957f
C269 VTAIL.n5 VSUBS 0.035353f
C270 VTAIL.n6 VSUBS 0.015837f
C271 VTAIL.n7 VSUBS 0.027834f
C272 VTAIL.n8 VSUBS 0.014957f
C273 VTAIL.n9 VSUBS 0.035353f
C274 VTAIL.n10 VSUBS 0.015837f
C275 VTAIL.n11 VSUBS 0.027834f
C276 VTAIL.n12 VSUBS 0.014957f
C277 VTAIL.n13 VSUBS 0.035353f
C278 VTAIL.n14 VSUBS 0.015837f
C279 VTAIL.n15 VSUBS 0.027834f
C280 VTAIL.n16 VSUBS 0.014957f
C281 VTAIL.n17 VSUBS 0.035353f
C282 VTAIL.n18 VSUBS 0.015837f
C283 VTAIL.n19 VSUBS 0.027834f
C284 VTAIL.n20 VSUBS 0.014957f
C285 VTAIL.n21 VSUBS 0.035353f
C286 VTAIL.n22 VSUBS 0.015837f
C287 VTAIL.n23 VSUBS 0.027834f
C288 VTAIL.n24 VSUBS 0.014957f
C289 VTAIL.n25 VSUBS 0.035353f
C290 VTAIL.n26 VSUBS 0.015837f
C291 VTAIL.n27 VSUBS 0.027834f
C292 VTAIL.n28 VSUBS 0.014957f
C293 VTAIL.n29 VSUBS 0.035353f
C294 VTAIL.n30 VSUBS 0.015837f
C295 VTAIL.n31 VSUBS 0.21033f
C296 VTAIL.t8 VSUBS 0.075803f
C297 VTAIL.n32 VSUBS 0.026515f
C298 VTAIL.n33 VSUBS 0.02249f
C299 VTAIL.n34 VSUBS 0.014957f
C300 VTAIL.n35 VSUBS 1.99463f
C301 VTAIL.n36 VSUBS 0.027834f
C302 VTAIL.n37 VSUBS 0.014957f
C303 VTAIL.n38 VSUBS 0.015837f
C304 VTAIL.n39 VSUBS 0.035353f
C305 VTAIL.n40 VSUBS 0.035353f
C306 VTAIL.n41 VSUBS 0.015837f
C307 VTAIL.n42 VSUBS 0.014957f
C308 VTAIL.n43 VSUBS 0.027834f
C309 VTAIL.n44 VSUBS 0.027834f
C310 VTAIL.n45 VSUBS 0.014957f
C311 VTAIL.n46 VSUBS 0.015837f
C312 VTAIL.n47 VSUBS 0.035353f
C313 VTAIL.n48 VSUBS 0.035353f
C314 VTAIL.n49 VSUBS 0.015837f
C315 VTAIL.n50 VSUBS 0.014957f
C316 VTAIL.n51 VSUBS 0.027834f
C317 VTAIL.n52 VSUBS 0.027834f
C318 VTAIL.n53 VSUBS 0.014957f
C319 VTAIL.n54 VSUBS 0.015837f
C320 VTAIL.n55 VSUBS 0.035353f
C321 VTAIL.n56 VSUBS 0.035353f
C322 VTAIL.n57 VSUBS 0.015837f
C323 VTAIL.n58 VSUBS 0.014957f
C324 VTAIL.n59 VSUBS 0.027834f
C325 VTAIL.n60 VSUBS 0.027834f
C326 VTAIL.n61 VSUBS 0.014957f
C327 VTAIL.n62 VSUBS 0.015837f
C328 VTAIL.n63 VSUBS 0.035353f
C329 VTAIL.n64 VSUBS 0.035353f
C330 VTAIL.n65 VSUBS 0.015837f
C331 VTAIL.n66 VSUBS 0.014957f
C332 VTAIL.n67 VSUBS 0.027834f
C333 VTAIL.n68 VSUBS 0.027834f
C334 VTAIL.n69 VSUBS 0.014957f
C335 VTAIL.n70 VSUBS 0.015837f
C336 VTAIL.n71 VSUBS 0.035353f
C337 VTAIL.n72 VSUBS 0.035353f
C338 VTAIL.n73 VSUBS 0.035353f
C339 VTAIL.n74 VSUBS 0.015837f
C340 VTAIL.n75 VSUBS 0.014957f
C341 VTAIL.n76 VSUBS 0.027834f
C342 VTAIL.n77 VSUBS 0.027834f
C343 VTAIL.n78 VSUBS 0.014957f
C344 VTAIL.n79 VSUBS 0.015397f
C345 VTAIL.n80 VSUBS 0.015397f
C346 VTAIL.n81 VSUBS 0.035353f
C347 VTAIL.n82 VSUBS 0.035353f
C348 VTAIL.n83 VSUBS 0.015837f
C349 VTAIL.n84 VSUBS 0.014957f
C350 VTAIL.n85 VSUBS 0.027834f
C351 VTAIL.n86 VSUBS 0.027834f
C352 VTAIL.n87 VSUBS 0.014957f
C353 VTAIL.n88 VSUBS 0.015837f
C354 VTAIL.n89 VSUBS 0.035353f
C355 VTAIL.n90 VSUBS 0.078759f
C356 VTAIL.n91 VSUBS 0.015837f
C357 VTAIL.n92 VSUBS 0.014957f
C358 VTAIL.n93 VSUBS 0.061296f
C359 VTAIL.n94 VSUBS 0.039209f
C360 VTAIL.n95 VSUBS 0.423726f
C361 VTAIL.t5 VSUBS 0.367768f
C362 VTAIL.t10 VSUBS 0.367768f
C363 VTAIL.n96 VSUBS 2.84058f
C364 VTAIL.n97 VSUBS 3.0817f
C365 VTAIL.t0 VSUBS 0.367768f
C366 VTAIL.t3 VSUBS 0.367768f
C367 VTAIL.n98 VSUBS 2.8406f
C368 VTAIL.n99 VSUBS 3.08168f
C369 VTAIL.n100 VSUBS 0.02858f
C370 VTAIL.n101 VSUBS 0.027834f
C371 VTAIL.n102 VSUBS 0.014957f
C372 VTAIL.n103 VSUBS 0.035353f
C373 VTAIL.n104 VSUBS 0.015837f
C374 VTAIL.n105 VSUBS 0.027834f
C375 VTAIL.n106 VSUBS 0.014957f
C376 VTAIL.n107 VSUBS 0.035353f
C377 VTAIL.n108 VSUBS 0.015837f
C378 VTAIL.n109 VSUBS 0.027834f
C379 VTAIL.n110 VSUBS 0.014957f
C380 VTAIL.n111 VSUBS 0.035353f
C381 VTAIL.n112 VSUBS 0.035353f
C382 VTAIL.n113 VSUBS 0.015837f
C383 VTAIL.n114 VSUBS 0.027834f
C384 VTAIL.n115 VSUBS 0.014957f
C385 VTAIL.n116 VSUBS 0.035353f
C386 VTAIL.n117 VSUBS 0.015837f
C387 VTAIL.n118 VSUBS 0.027834f
C388 VTAIL.n119 VSUBS 0.014957f
C389 VTAIL.n120 VSUBS 0.035353f
C390 VTAIL.n121 VSUBS 0.015837f
C391 VTAIL.n122 VSUBS 0.027834f
C392 VTAIL.n123 VSUBS 0.014957f
C393 VTAIL.n124 VSUBS 0.035353f
C394 VTAIL.n125 VSUBS 0.015837f
C395 VTAIL.n126 VSUBS 0.027834f
C396 VTAIL.n127 VSUBS 0.014957f
C397 VTAIL.n128 VSUBS 0.035353f
C398 VTAIL.n129 VSUBS 0.015837f
C399 VTAIL.n130 VSUBS 0.21033f
C400 VTAIL.t1 VSUBS 0.075803f
C401 VTAIL.n131 VSUBS 0.026515f
C402 VTAIL.n132 VSUBS 0.02249f
C403 VTAIL.n133 VSUBS 0.014957f
C404 VTAIL.n134 VSUBS 1.99463f
C405 VTAIL.n135 VSUBS 0.027834f
C406 VTAIL.n136 VSUBS 0.014957f
C407 VTAIL.n137 VSUBS 0.015837f
C408 VTAIL.n138 VSUBS 0.035353f
C409 VTAIL.n139 VSUBS 0.035353f
C410 VTAIL.n140 VSUBS 0.015837f
C411 VTAIL.n141 VSUBS 0.014957f
C412 VTAIL.n142 VSUBS 0.027834f
C413 VTAIL.n143 VSUBS 0.027834f
C414 VTAIL.n144 VSUBS 0.014957f
C415 VTAIL.n145 VSUBS 0.015837f
C416 VTAIL.n146 VSUBS 0.035353f
C417 VTAIL.n147 VSUBS 0.035353f
C418 VTAIL.n148 VSUBS 0.015837f
C419 VTAIL.n149 VSUBS 0.014957f
C420 VTAIL.n150 VSUBS 0.027834f
C421 VTAIL.n151 VSUBS 0.027834f
C422 VTAIL.n152 VSUBS 0.014957f
C423 VTAIL.n153 VSUBS 0.015837f
C424 VTAIL.n154 VSUBS 0.035353f
C425 VTAIL.n155 VSUBS 0.035353f
C426 VTAIL.n156 VSUBS 0.015837f
C427 VTAIL.n157 VSUBS 0.014957f
C428 VTAIL.n158 VSUBS 0.027834f
C429 VTAIL.n159 VSUBS 0.027834f
C430 VTAIL.n160 VSUBS 0.014957f
C431 VTAIL.n161 VSUBS 0.015837f
C432 VTAIL.n162 VSUBS 0.035353f
C433 VTAIL.n163 VSUBS 0.035353f
C434 VTAIL.n164 VSUBS 0.015837f
C435 VTAIL.n165 VSUBS 0.014957f
C436 VTAIL.n166 VSUBS 0.027834f
C437 VTAIL.n167 VSUBS 0.027834f
C438 VTAIL.n168 VSUBS 0.014957f
C439 VTAIL.n169 VSUBS 0.015837f
C440 VTAIL.n170 VSUBS 0.035353f
C441 VTAIL.n171 VSUBS 0.035353f
C442 VTAIL.n172 VSUBS 0.015837f
C443 VTAIL.n173 VSUBS 0.014957f
C444 VTAIL.n174 VSUBS 0.027834f
C445 VTAIL.n175 VSUBS 0.027834f
C446 VTAIL.n176 VSUBS 0.014957f
C447 VTAIL.n177 VSUBS 0.015397f
C448 VTAIL.n178 VSUBS 0.015397f
C449 VTAIL.n179 VSUBS 0.035353f
C450 VTAIL.n180 VSUBS 0.035353f
C451 VTAIL.n181 VSUBS 0.015837f
C452 VTAIL.n182 VSUBS 0.014957f
C453 VTAIL.n183 VSUBS 0.027834f
C454 VTAIL.n184 VSUBS 0.027834f
C455 VTAIL.n185 VSUBS 0.014957f
C456 VTAIL.n186 VSUBS 0.015837f
C457 VTAIL.n187 VSUBS 0.035353f
C458 VTAIL.n188 VSUBS 0.078759f
C459 VTAIL.n189 VSUBS 0.015837f
C460 VTAIL.n190 VSUBS 0.014957f
C461 VTAIL.n191 VSUBS 0.061296f
C462 VTAIL.n192 VSUBS 0.039209f
C463 VTAIL.n193 VSUBS 0.423726f
C464 VTAIL.t7 VSUBS 0.367768f
C465 VTAIL.t9 VSUBS 0.367768f
C466 VTAIL.n194 VSUBS 2.8406f
C467 VTAIL.n195 VSUBS 1.09343f
C468 VTAIL.n196 VSUBS 0.02858f
C469 VTAIL.n197 VSUBS 0.027834f
C470 VTAIL.n198 VSUBS 0.014957f
C471 VTAIL.n199 VSUBS 0.035353f
C472 VTAIL.n200 VSUBS 0.015837f
C473 VTAIL.n201 VSUBS 0.027834f
C474 VTAIL.n202 VSUBS 0.014957f
C475 VTAIL.n203 VSUBS 0.035353f
C476 VTAIL.n204 VSUBS 0.015837f
C477 VTAIL.n205 VSUBS 0.027834f
C478 VTAIL.n206 VSUBS 0.014957f
C479 VTAIL.n207 VSUBS 0.035353f
C480 VTAIL.n208 VSUBS 0.035353f
C481 VTAIL.n209 VSUBS 0.015837f
C482 VTAIL.n210 VSUBS 0.027834f
C483 VTAIL.n211 VSUBS 0.014957f
C484 VTAIL.n212 VSUBS 0.035353f
C485 VTAIL.n213 VSUBS 0.015837f
C486 VTAIL.n214 VSUBS 0.027834f
C487 VTAIL.n215 VSUBS 0.014957f
C488 VTAIL.n216 VSUBS 0.035353f
C489 VTAIL.n217 VSUBS 0.015837f
C490 VTAIL.n218 VSUBS 0.027834f
C491 VTAIL.n219 VSUBS 0.014957f
C492 VTAIL.n220 VSUBS 0.035353f
C493 VTAIL.n221 VSUBS 0.015837f
C494 VTAIL.n222 VSUBS 0.027834f
C495 VTAIL.n223 VSUBS 0.014957f
C496 VTAIL.n224 VSUBS 0.035353f
C497 VTAIL.n225 VSUBS 0.015837f
C498 VTAIL.n226 VSUBS 0.21033f
C499 VTAIL.t6 VSUBS 0.075803f
C500 VTAIL.n227 VSUBS 0.026515f
C501 VTAIL.n228 VSUBS 0.02249f
C502 VTAIL.n229 VSUBS 0.014957f
C503 VTAIL.n230 VSUBS 1.99463f
C504 VTAIL.n231 VSUBS 0.027834f
C505 VTAIL.n232 VSUBS 0.014957f
C506 VTAIL.n233 VSUBS 0.015837f
C507 VTAIL.n234 VSUBS 0.035353f
C508 VTAIL.n235 VSUBS 0.035353f
C509 VTAIL.n236 VSUBS 0.015837f
C510 VTAIL.n237 VSUBS 0.014957f
C511 VTAIL.n238 VSUBS 0.027834f
C512 VTAIL.n239 VSUBS 0.027834f
C513 VTAIL.n240 VSUBS 0.014957f
C514 VTAIL.n241 VSUBS 0.015837f
C515 VTAIL.n242 VSUBS 0.035353f
C516 VTAIL.n243 VSUBS 0.035353f
C517 VTAIL.n244 VSUBS 0.015837f
C518 VTAIL.n245 VSUBS 0.014957f
C519 VTAIL.n246 VSUBS 0.027834f
C520 VTAIL.n247 VSUBS 0.027834f
C521 VTAIL.n248 VSUBS 0.014957f
C522 VTAIL.n249 VSUBS 0.015837f
C523 VTAIL.n250 VSUBS 0.035353f
C524 VTAIL.n251 VSUBS 0.035353f
C525 VTAIL.n252 VSUBS 0.015837f
C526 VTAIL.n253 VSUBS 0.014957f
C527 VTAIL.n254 VSUBS 0.027834f
C528 VTAIL.n255 VSUBS 0.027834f
C529 VTAIL.n256 VSUBS 0.014957f
C530 VTAIL.n257 VSUBS 0.015837f
C531 VTAIL.n258 VSUBS 0.035353f
C532 VTAIL.n259 VSUBS 0.035353f
C533 VTAIL.n260 VSUBS 0.015837f
C534 VTAIL.n261 VSUBS 0.014957f
C535 VTAIL.n262 VSUBS 0.027834f
C536 VTAIL.n263 VSUBS 0.027834f
C537 VTAIL.n264 VSUBS 0.014957f
C538 VTAIL.n265 VSUBS 0.015837f
C539 VTAIL.n266 VSUBS 0.035353f
C540 VTAIL.n267 VSUBS 0.035353f
C541 VTAIL.n268 VSUBS 0.015837f
C542 VTAIL.n269 VSUBS 0.014957f
C543 VTAIL.n270 VSUBS 0.027834f
C544 VTAIL.n271 VSUBS 0.027834f
C545 VTAIL.n272 VSUBS 0.014957f
C546 VTAIL.n273 VSUBS 0.015397f
C547 VTAIL.n274 VSUBS 0.015397f
C548 VTAIL.n275 VSUBS 0.035353f
C549 VTAIL.n276 VSUBS 0.035353f
C550 VTAIL.n277 VSUBS 0.015837f
C551 VTAIL.n278 VSUBS 0.014957f
C552 VTAIL.n279 VSUBS 0.027834f
C553 VTAIL.n280 VSUBS 0.027834f
C554 VTAIL.n281 VSUBS 0.014957f
C555 VTAIL.n282 VSUBS 0.015837f
C556 VTAIL.n283 VSUBS 0.035353f
C557 VTAIL.n284 VSUBS 0.078759f
C558 VTAIL.n285 VSUBS 0.015837f
C559 VTAIL.n286 VSUBS 0.014957f
C560 VTAIL.n287 VSUBS 0.061296f
C561 VTAIL.n288 VSUBS 0.039209f
C562 VTAIL.n289 VSUBS 2.17229f
C563 VTAIL.n290 VSUBS 0.02858f
C564 VTAIL.n291 VSUBS 0.027834f
C565 VTAIL.n292 VSUBS 0.014957f
C566 VTAIL.n293 VSUBS 0.035353f
C567 VTAIL.n294 VSUBS 0.015837f
C568 VTAIL.n295 VSUBS 0.027834f
C569 VTAIL.n296 VSUBS 0.014957f
C570 VTAIL.n297 VSUBS 0.035353f
C571 VTAIL.n298 VSUBS 0.015837f
C572 VTAIL.n299 VSUBS 0.027834f
C573 VTAIL.n300 VSUBS 0.014957f
C574 VTAIL.n301 VSUBS 0.035353f
C575 VTAIL.n302 VSUBS 0.015837f
C576 VTAIL.n303 VSUBS 0.027834f
C577 VTAIL.n304 VSUBS 0.014957f
C578 VTAIL.n305 VSUBS 0.035353f
C579 VTAIL.n306 VSUBS 0.015837f
C580 VTAIL.n307 VSUBS 0.027834f
C581 VTAIL.n308 VSUBS 0.014957f
C582 VTAIL.n309 VSUBS 0.035353f
C583 VTAIL.n310 VSUBS 0.015837f
C584 VTAIL.n311 VSUBS 0.027834f
C585 VTAIL.n312 VSUBS 0.014957f
C586 VTAIL.n313 VSUBS 0.035353f
C587 VTAIL.n314 VSUBS 0.015837f
C588 VTAIL.n315 VSUBS 0.027834f
C589 VTAIL.n316 VSUBS 0.014957f
C590 VTAIL.n317 VSUBS 0.035353f
C591 VTAIL.n318 VSUBS 0.015837f
C592 VTAIL.n319 VSUBS 0.21033f
C593 VTAIL.t11 VSUBS 0.075803f
C594 VTAIL.n320 VSUBS 0.026515f
C595 VTAIL.n321 VSUBS 0.02249f
C596 VTAIL.n322 VSUBS 0.014957f
C597 VTAIL.n323 VSUBS 1.99463f
C598 VTAIL.n324 VSUBS 0.027834f
C599 VTAIL.n325 VSUBS 0.014957f
C600 VTAIL.n326 VSUBS 0.015837f
C601 VTAIL.n327 VSUBS 0.035353f
C602 VTAIL.n328 VSUBS 0.035353f
C603 VTAIL.n329 VSUBS 0.015837f
C604 VTAIL.n330 VSUBS 0.014957f
C605 VTAIL.n331 VSUBS 0.027834f
C606 VTAIL.n332 VSUBS 0.027834f
C607 VTAIL.n333 VSUBS 0.014957f
C608 VTAIL.n334 VSUBS 0.015837f
C609 VTAIL.n335 VSUBS 0.035353f
C610 VTAIL.n336 VSUBS 0.035353f
C611 VTAIL.n337 VSUBS 0.015837f
C612 VTAIL.n338 VSUBS 0.014957f
C613 VTAIL.n339 VSUBS 0.027834f
C614 VTAIL.n340 VSUBS 0.027834f
C615 VTAIL.n341 VSUBS 0.014957f
C616 VTAIL.n342 VSUBS 0.015837f
C617 VTAIL.n343 VSUBS 0.035353f
C618 VTAIL.n344 VSUBS 0.035353f
C619 VTAIL.n345 VSUBS 0.015837f
C620 VTAIL.n346 VSUBS 0.014957f
C621 VTAIL.n347 VSUBS 0.027834f
C622 VTAIL.n348 VSUBS 0.027834f
C623 VTAIL.n349 VSUBS 0.014957f
C624 VTAIL.n350 VSUBS 0.015837f
C625 VTAIL.n351 VSUBS 0.035353f
C626 VTAIL.n352 VSUBS 0.035353f
C627 VTAIL.n353 VSUBS 0.015837f
C628 VTAIL.n354 VSUBS 0.014957f
C629 VTAIL.n355 VSUBS 0.027834f
C630 VTAIL.n356 VSUBS 0.027834f
C631 VTAIL.n357 VSUBS 0.014957f
C632 VTAIL.n358 VSUBS 0.015837f
C633 VTAIL.n359 VSUBS 0.035353f
C634 VTAIL.n360 VSUBS 0.035353f
C635 VTAIL.n361 VSUBS 0.035353f
C636 VTAIL.n362 VSUBS 0.015837f
C637 VTAIL.n363 VSUBS 0.014957f
C638 VTAIL.n364 VSUBS 0.027834f
C639 VTAIL.n365 VSUBS 0.027834f
C640 VTAIL.n366 VSUBS 0.014957f
C641 VTAIL.n367 VSUBS 0.015397f
C642 VTAIL.n368 VSUBS 0.015397f
C643 VTAIL.n369 VSUBS 0.035353f
C644 VTAIL.n370 VSUBS 0.035353f
C645 VTAIL.n371 VSUBS 0.015837f
C646 VTAIL.n372 VSUBS 0.014957f
C647 VTAIL.n373 VSUBS 0.027834f
C648 VTAIL.n374 VSUBS 0.027834f
C649 VTAIL.n375 VSUBS 0.014957f
C650 VTAIL.n376 VSUBS 0.015837f
C651 VTAIL.n377 VSUBS 0.035353f
C652 VTAIL.n378 VSUBS 0.078759f
C653 VTAIL.n379 VSUBS 0.015837f
C654 VTAIL.n380 VSUBS 0.014957f
C655 VTAIL.n381 VSUBS 0.061296f
C656 VTAIL.n382 VSUBS 0.039209f
C657 VTAIL.n383 VSUBS 2.10715f
C658 VDD1.n0 VSUBS 0.027885f
C659 VDD1.n1 VSUBS 0.027158f
C660 VDD1.n2 VSUBS 0.014594f
C661 VDD1.n3 VSUBS 0.034494f
C662 VDD1.n4 VSUBS 0.015452f
C663 VDD1.n5 VSUBS 0.027158f
C664 VDD1.n6 VSUBS 0.014594f
C665 VDD1.n7 VSUBS 0.034494f
C666 VDD1.n8 VSUBS 0.015452f
C667 VDD1.n9 VSUBS 0.027158f
C668 VDD1.n10 VSUBS 0.014594f
C669 VDD1.n11 VSUBS 0.034494f
C670 VDD1.n12 VSUBS 0.034494f
C671 VDD1.n13 VSUBS 0.015452f
C672 VDD1.n14 VSUBS 0.027158f
C673 VDD1.n15 VSUBS 0.014594f
C674 VDD1.n16 VSUBS 0.034494f
C675 VDD1.n17 VSUBS 0.015452f
C676 VDD1.n18 VSUBS 0.027158f
C677 VDD1.n19 VSUBS 0.014594f
C678 VDD1.n20 VSUBS 0.034494f
C679 VDD1.n21 VSUBS 0.015452f
C680 VDD1.n22 VSUBS 0.027158f
C681 VDD1.n23 VSUBS 0.014594f
C682 VDD1.n24 VSUBS 0.034494f
C683 VDD1.n25 VSUBS 0.015452f
C684 VDD1.n26 VSUBS 0.027158f
C685 VDD1.n27 VSUBS 0.014594f
C686 VDD1.n28 VSUBS 0.034494f
C687 VDD1.n29 VSUBS 0.015452f
C688 VDD1.n30 VSUBS 0.205219f
C689 VDD1.t1 VSUBS 0.07396f
C690 VDD1.n31 VSUBS 0.02587f
C691 VDD1.n32 VSUBS 0.021943f
C692 VDD1.n33 VSUBS 0.014594f
C693 VDD1.n34 VSUBS 1.94616f
C694 VDD1.n35 VSUBS 0.027158f
C695 VDD1.n36 VSUBS 0.014594f
C696 VDD1.n37 VSUBS 0.015452f
C697 VDD1.n38 VSUBS 0.034494f
C698 VDD1.n39 VSUBS 0.034494f
C699 VDD1.n40 VSUBS 0.015452f
C700 VDD1.n41 VSUBS 0.014594f
C701 VDD1.n42 VSUBS 0.027158f
C702 VDD1.n43 VSUBS 0.027158f
C703 VDD1.n44 VSUBS 0.014594f
C704 VDD1.n45 VSUBS 0.015452f
C705 VDD1.n46 VSUBS 0.034494f
C706 VDD1.n47 VSUBS 0.034494f
C707 VDD1.n48 VSUBS 0.015452f
C708 VDD1.n49 VSUBS 0.014594f
C709 VDD1.n50 VSUBS 0.027158f
C710 VDD1.n51 VSUBS 0.027158f
C711 VDD1.n52 VSUBS 0.014594f
C712 VDD1.n53 VSUBS 0.015452f
C713 VDD1.n54 VSUBS 0.034494f
C714 VDD1.n55 VSUBS 0.034494f
C715 VDD1.n56 VSUBS 0.015452f
C716 VDD1.n57 VSUBS 0.014594f
C717 VDD1.n58 VSUBS 0.027158f
C718 VDD1.n59 VSUBS 0.027158f
C719 VDD1.n60 VSUBS 0.014594f
C720 VDD1.n61 VSUBS 0.015452f
C721 VDD1.n62 VSUBS 0.034494f
C722 VDD1.n63 VSUBS 0.034494f
C723 VDD1.n64 VSUBS 0.015452f
C724 VDD1.n65 VSUBS 0.014594f
C725 VDD1.n66 VSUBS 0.027158f
C726 VDD1.n67 VSUBS 0.027158f
C727 VDD1.n68 VSUBS 0.014594f
C728 VDD1.n69 VSUBS 0.015452f
C729 VDD1.n70 VSUBS 0.034494f
C730 VDD1.n71 VSUBS 0.034494f
C731 VDD1.n72 VSUBS 0.015452f
C732 VDD1.n73 VSUBS 0.014594f
C733 VDD1.n74 VSUBS 0.027158f
C734 VDD1.n75 VSUBS 0.027158f
C735 VDD1.n76 VSUBS 0.014594f
C736 VDD1.n77 VSUBS 0.015023f
C737 VDD1.n78 VSUBS 0.015023f
C738 VDD1.n79 VSUBS 0.034494f
C739 VDD1.n80 VSUBS 0.034494f
C740 VDD1.n81 VSUBS 0.015452f
C741 VDD1.n82 VSUBS 0.014594f
C742 VDD1.n83 VSUBS 0.027158f
C743 VDD1.n84 VSUBS 0.027158f
C744 VDD1.n85 VSUBS 0.014594f
C745 VDD1.n86 VSUBS 0.015452f
C746 VDD1.n87 VSUBS 0.034494f
C747 VDD1.n88 VSUBS 0.076845f
C748 VDD1.n89 VSUBS 0.015452f
C749 VDD1.n90 VSUBS 0.014594f
C750 VDD1.n91 VSUBS 0.059807f
C751 VDD1.n92 VSUBS 0.066686f
C752 VDD1.n93 VSUBS 0.027885f
C753 VDD1.n94 VSUBS 0.027158f
C754 VDD1.n95 VSUBS 0.014594f
C755 VDD1.n96 VSUBS 0.034494f
C756 VDD1.n97 VSUBS 0.015452f
C757 VDD1.n98 VSUBS 0.027158f
C758 VDD1.n99 VSUBS 0.014594f
C759 VDD1.n100 VSUBS 0.034494f
C760 VDD1.n101 VSUBS 0.015452f
C761 VDD1.n102 VSUBS 0.027158f
C762 VDD1.n103 VSUBS 0.014594f
C763 VDD1.n104 VSUBS 0.034494f
C764 VDD1.n105 VSUBS 0.015452f
C765 VDD1.n106 VSUBS 0.027158f
C766 VDD1.n107 VSUBS 0.014594f
C767 VDD1.n108 VSUBS 0.034494f
C768 VDD1.n109 VSUBS 0.015452f
C769 VDD1.n110 VSUBS 0.027158f
C770 VDD1.n111 VSUBS 0.014594f
C771 VDD1.n112 VSUBS 0.034494f
C772 VDD1.n113 VSUBS 0.015452f
C773 VDD1.n114 VSUBS 0.027158f
C774 VDD1.n115 VSUBS 0.014594f
C775 VDD1.n116 VSUBS 0.034494f
C776 VDD1.n117 VSUBS 0.015452f
C777 VDD1.n118 VSUBS 0.027158f
C778 VDD1.n119 VSUBS 0.014594f
C779 VDD1.n120 VSUBS 0.034494f
C780 VDD1.n121 VSUBS 0.015452f
C781 VDD1.n122 VSUBS 0.205219f
C782 VDD1.t0 VSUBS 0.07396f
C783 VDD1.n123 VSUBS 0.02587f
C784 VDD1.n124 VSUBS 0.021943f
C785 VDD1.n125 VSUBS 0.014594f
C786 VDD1.n126 VSUBS 1.94616f
C787 VDD1.n127 VSUBS 0.027158f
C788 VDD1.n128 VSUBS 0.014594f
C789 VDD1.n129 VSUBS 0.015452f
C790 VDD1.n130 VSUBS 0.034494f
C791 VDD1.n131 VSUBS 0.034494f
C792 VDD1.n132 VSUBS 0.015452f
C793 VDD1.n133 VSUBS 0.014594f
C794 VDD1.n134 VSUBS 0.027158f
C795 VDD1.n135 VSUBS 0.027158f
C796 VDD1.n136 VSUBS 0.014594f
C797 VDD1.n137 VSUBS 0.015452f
C798 VDD1.n138 VSUBS 0.034494f
C799 VDD1.n139 VSUBS 0.034494f
C800 VDD1.n140 VSUBS 0.015452f
C801 VDD1.n141 VSUBS 0.014594f
C802 VDD1.n142 VSUBS 0.027158f
C803 VDD1.n143 VSUBS 0.027158f
C804 VDD1.n144 VSUBS 0.014594f
C805 VDD1.n145 VSUBS 0.015452f
C806 VDD1.n146 VSUBS 0.034494f
C807 VDD1.n147 VSUBS 0.034494f
C808 VDD1.n148 VSUBS 0.015452f
C809 VDD1.n149 VSUBS 0.014594f
C810 VDD1.n150 VSUBS 0.027158f
C811 VDD1.n151 VSUBS 0.027158f
C812 VDD1.n152 VSUBS 0.014594f
C813 VDD1.n153 VSUBS 0.015452f
C814 VDD1.n154 VSUBS 0.034494f
C815 VDD1.n155 VSUBS 0.034494f
C816 VDD1.n156 VSUBS 0.015452f
C817 VDD1.n157 VSUBS 0.014594f
C818 VDD1.n158 VSUBS 0.027158f
C819 VDD1.n159 VSUBS 0.027158f
C820 VDD1.n160 VSUBS 0.014594f
C821 VDD1.n161 VSUBS 0.015452f
C822 VDD1.n162 VSUBS 0.034494f
C823 VDD1.n163 VSUBS 0.034494f
C824 VDD1.n164 VSUBS 0.034494f
C825 VDD1.n165 VSUBS 0.015452f
C826 VDD1.n166 VSUBS 0.014594f
C827 VDD1.n167 VSUBS 0.027158f
C828 VDD1.n168 VSUBS 0.027158f
C829 VDD1.n169 VSUBS 0.014594f
C830 VDD1.n170 VSUBS 0.015023f
C831 VDD1.n171 VSUBS 0.015023f
C832 VDD1.n172 VSUBS 0.034494f
C833 VDD1.n173 VSUBS 0.034494f
C834 VDD1.n174 VSUBS 0.015452f
C835 VDD1.n175 VSUBS 0.014594f
C836 VDD1.n176 VSUBS 0.027158f
C837 VDD1.n177 VSUBS 0.027158f
C838 VDD1.n178 VSUBS 0.014594f
C839 VDD1.n179 VSUBS 0.015452f
C840 VDD1.n180 VSUBS 0.034494f
C841 VDD1.n181 VSUBS 0.076845f
C842 VDD1.n182 VSUBS 0.015452f
C843 VDD1.n183 VSUBS 0.014594f
C844 VDD1.n184 VSUBS 0.059807f
C845 VDD1.n185 VSUBS 0.065795f
C846 VDD1.t4 VSUBS 0.35883f
C847 VDD1.t5 VSUBS 0.35883f
C848 VDD1.n186 VSUBS 2.95279f
C849 VDD1.n187 VSUBS 3.7624f
C850 VDD1.t3 VSUBS 0.35883f
C851 VDD1.t2 VSUBS 0.35883f
C852 VDD1.n188 VSUBS 2.94529f
C853 VDD1.n189 VSUBS 3.7857f
C854 VP.n0 VSUBS 0.038369f
C855 VP.t2 VSUBS 3.70227f
C856 VP.n1 VSUBS 0.055682f
C857 VP.n2 VSUBS 0.029104f
C858 VP.t0 VSUBS 3.70227f
C859 VP.n3 VSUBS 1.31317f
C860 VP.n4 VSUBS 0.029104f
C861 VP.n5 VSUBS 0.055682f
C862 VP.n6 VSUBS 0.038369f
C863 VP.t5 VSUBS 3.70227f
C864 VP.n7 VSUBS 0.038369f
C865 VP.t4 VSUBS 3.70227f
C866 VP.n8 VSUBS 0.055682f
C867 VP.n9 VSUBS 0.029104f
C868 VP.t1 VSUBS 3.70227f
C869 VP.n10 VSUBS 1.38893f
C870 VP.t3 VSUBS 3.98289f
C871 VP.n11 VSUBS 1.33128f
C872 VP.n12 VSUBS 0.304498f
C873 VP.n13 VSUBS 0.053971f
C874 VP.n14 VSUBS 0.058457f
C875 VP.n15 VSUBS 0.024448f
C876 VP.n16 VSUBS 0.029104f
C877 VP.n17 VSUBS 0.029104f
C878 VP.n18 VSUBS 0.029104f
C879 VP.n19 VSUBS 0.053971f
C880 VP.n20 VSUBS 0.032656f
C881 VP.n21 VSUBS 1.38129f
C882 VP.n22 VSUBS 1.76269f
C883 VP.n23 VSUBS 1.78252f
C884 VP.n24 VSUBS 1.38129f
C885 VP.n25 VSUBS 0.032656f
C886 VP.n26 VSUBS 0.053971f
C887 VP.n27 VSUBS 0.029104f
C888 VP.n28 VSUBS 0.029104f
C889 VP.n29 VSUBS 0.029104f
C890 VP.n30 VSUBS 0.024448f
C891 VP.n31 VSUBS 0.058457f
C892 VP.n32 VSUBS 0.053971f
C893 VP.n33 VSUBS 0.029104f
C894 VP.n34 VSUBS 0.029104f
C895 VP.n35 VSUBS 0.029104f
C896 VP.n36 VSUBS 0.053971f
C897 VP.n37 VSUBS 0.058457f
C898 VP.n38 VSUBS 0.024448f
C899 VP.n39 VSUBS 0.029104f
C900 VP.n40 VSUBS 0.029104f
C901 VP.n41 VSUBS 0.029104f
C902 VP.n42 VSUBS 0.053971f
C903 VP.n43 VSUBS 0.032656f
C904 VP.n44 VSUBS 1.38129f
C905 VP.n45 VSUBS 0.052628f
C906 B.n0 VSUBS 0.006935f
C907 B.n1 VSUBS 0.006935f
C908 B.n2 VSUBS 0.010256f
C909 B.n3 VSUBS 0.007859f
C910 B.n4 VSUBS 0.007859f
C911 B.n5 VSUBS 0.007859f
C912 B.n6 VSUBS 0.007859f
C913 B.n7 VSUBS 0.007859f
C914 B.n8 VSUBS 0.007859f
C915 B.n9 VSUBS 0.007859f
C916 B.n10 VSUBS 0.007859f
C917 B.n11 VSUBS 0.007859f
C918 B.n12 VSUBS 0.007859f
C919 B.n13 VSUBS 0.007859f
C920 B.n14 VSUBS 0.007859f
C921 B.n15 VSUBS 0.007859f
C922 B.n16 VSUBS 0.007859f
C923 B.n17 VSUBS 0.007859f
C924 B.n18 VSUBS 0.007859f
C925 B.n19 VSUBS 0.007859f
C926 B.n20 VSUBS 0.007859f
C927 B.n21 VSUBS 0.007859f
C928 B.n22 VSUBS 0.007859f
C929 B.n23 VSUBS 0.007859f
C930 B.n24 VSUBS 0.018502f
C931 B.n25 VSUBS 0.007859f
C932 B.n26 VSUBS 0.007859f
C933 B.n27 VSUBS 0.007859f
C934 B.n28 VSUBS 0.007859f
C935 B.n29 VSUBS 0.007859f
C936 B.n30 VSUBS 0.007859f
C937 B.n31 VSUBS 0.007859f
C938 B.n32 VSUBS 0.007859f
C939 B.n33 VSUBS 0.007859f
C940 B.n34 VSUBS 0.007859f
C941 B.n35 VSUBS 0.007859f
C942 B.n36 VSUBS 0.007859f
C943 B.n37 VSUBS 0.007859f
C944 B.n38 VSUBS 0.007859f
C945 B.n39 VSUBS 0.007859f
C946 B.n40 VSUBS 0.007859f
C947 B.n41 VSUBS 0.007859f
C948 B.n42 VSUBS 0.007859f
C949 B.n43 VSUBS 0.007859f
C950 B.n44 VSUBS 0.007859f
C951 B.n45 VSUBS 0.007859f
C952 B.n46 VSUBS 0.007859f
C953 B.n47 VSUBS 0.007859f
C954 B.n48 VSUBS 0.007859f
C955 B.n49 VSUBS 0.007859f
C956 B.n50 VSUBS 0.007859f
C957 B.n51 VSUBS 0.007859f
C958 B.t7 VSUBS 0.35944f
C959 B.t8 VSUBS 0.398869f
C960 B.t6 VSUBS 2.32891f
C961 B.n52 VSUBS 0.61926f
C962 B.n53 VSUBS 0.352633f
C963 B.n54 VSUBS 0.018209f
C964 B.n55 VSUBS 0.007859f
C965 B.n56 VSUBS 0.007859f
C966 B.n57 VSUBS 0.007859f
C967 B.n58 VSUBS 0.007859f
C968 B.n59 VSUBS 0.007859f
C969 B.t10 VSUBS 0.359444f
C970 B.t11 VSUBS 0.398872f
C971 B.t9 VSUBS 2.32891f
C972 B.n60 VSUBS 0.619257f
C973 B.n61 VSUBS 0.352629f
C974 B.n62 VSUBS 0.007859f
C975 B.n63 VSUBS 0.007859f
C976 B.n64 VSUBS 0.007859f
C977 B.n65 VSUBS 0.007859f
C978 B.n66 VSUBS 0.007859f
C979 B.n67 VSUBS 0.007859f
C980 B.n68 VSUBS 0.007859f
C981 B.n69 VSUBS 0.007859f
C982 B.n70 VSUBS 0.007859f
C983 B.n71 VSUBS 0.007859f
C984 B.n72 VSUBS 0.007859f
C985 B.n73 VSUBS 0.007859f
C986 B.n74 VSUBS 0.007859f
C987 B.n75 VSUBS 0.007859f
C988 B.n76 VSUBS 0.007859f
C989 B.n77 VSUBS 0.007859f
C990 B.n78 VSUBS 0.007859f
C991 B.n79 VSUBS 0.007859f
C992 B.n80 VSUBS 0.007859f
C993 B.n81 VSUBS 0.007859f
C994 B.n82 VSUBS 0.007859f
C995 B.n83 VSUBS 0.007859f
C996 B.n84 VSUBS 0.007859f
C997 B.n85 VSUBS 0.007859f
C998 B.n86 VSUBS 0.007859f
C999 B.n87 VSUBS 0.007859f
C1000 B.n88 VSUBS 0.007859f
C1001 B.n89 VSUBS 0.017097f
C1002 B.n90 VSUBS 0.007859f
C1003 B.n91 VSUBS 0.007859f
C1004 B.n92 VSUBS 0.007859f
C1005 B.n93 VSUBS 0.007859f
C1006 B.n94 VSUBS 0.007859f
C1007 B.n95 VSUBS 0.007859f
C1008 B.n96 VSUBS 0.007859f
C1009 B.n97 VSUBS 0.007859f
C1010 B.n98 VSUBS 0.007859f
C1011 B.n99 VSUBS 0.007859f
C1012 B.n100 VSUBS 0.007859f
C1013 B.n101 VSUBS 0.007859f
C1014 B.n102 VSUBS 0.007859f
C1015 B.n103 VSUBS 0.007859f
C1016 B.n104 VSUBS 0.007859f
C1017 B.n105 VSUBS 0.007859f
C1018 B.n106 VSUBS 0.007859f
C1019 B.n107 VSUBS 0.007859f
C1020 B.n108 VSUBS 0.007859f
C1021 B.n109 VSUBS 0.007859f
C1022 B.n110 VSUBS 0.007859f
C1023 B.n111 VSUBS 0.007859f
C1024 B.n112 VSUBS 0.007859f
C1025 B.n113 VSUBS 0.007859f
C1026 B.n114 VSUBS 0.007859f
C1027 B.n115 VSUBS 0.007859f
C1028 B.n116 VSUBS 0.007859f
C1029 B.n117 VSUBS 0.007859f
C1030 B.n118 VSUBS 0.007859f
C1031 B.n119 VSUBS 0.007859f
C1032 B.n120 VSUBS 0.007859f
C1033 B.n121 VSUBS 0.007859f
C1034 B.n122 VSUBS 0.007859f
C1035 B.n123 VSUBS 0.007859f
C1036 B.n124 VSUBS 0.007859f
C1037 B.n125 VSUBS 0.007859f
C1038 B.n126 VSUBS 0.007859f
C1039 B.n127 VSUBS 0.007859f
C1040 B.n128 VSUBS 0.007859f
C1041 B.n129 VSUBS 0.007859f
C1042 B.n130 VSUBS 0.007859f
C1043 B.n131 VSUBS 0.007859f
C1044 B.n132 VSUBS 0.007859f
C1045 B.n133 VSUBS 0.007859f
C1046 B.n134 VSUBS 0.017525f
C1047 B.n135 VSUBS 0.007859f
C1048 B.n136 VSUBS 0.007859f
C1049 B.n137 VSUBS 0.007859f
C1050 B.n138 VSUBS 0.007859f
C1051 B.n139 VSUBS 0.007859f
C1052 B.n140 VSUBS 0.007859f
C1053 B.n141 VSUBS 0.007859f
C1054 B.n142 VSUBS 0.007859f
C1055 B.n143 VSUBS 0.007859f
C1056 B.n144 VSUBS 0.007859f
C1057 B.n145 VSUBS 0.007859f
C1058 B.n146 VSUBS 0.007859f
C1059 B.n147 VSUBS 0.007859f
C1060 B.n148 VSUBS 0.007859f
C1061 B.n149 VSUBS 0.007859f
C1062 B.n150 VSUBS 0.007859f
C1063 B.n151 VSUBS 0.007859f
C1064 B.n152 VSUBS 0.007859f
C1065 B.n153 VSUBS 0.007859f
C1066 B.n154 VSUBS 0.007859f
C1067 B.n155 VSUBS 0.007859f
C1068 B.n156 VSUBS 0.007859f
C1069 B.n157 VSUBS 0.007859f
C1070 B.n158 VSUBS 0.007859f
C1071 B.n159 VSUBS 0.007859f
C1072 B.n160 VSUBS 0.007859f
C1073 B.n161 VSUBS 0.007859f
C1074 B.t5 VSUBS 0.359444f
C1075 B.t4 VSUBS 0.398872f
C1076 B.t3 VSUBS 2.32891f
C1077 B.n162 VSUBS 0.619257f
C1078 B.n163 VSUBS 0.352629f
C1079 B.n164 VSUBS 0.018209f
C1080 B.n165 VSUBS 0.007859f
C1081 B.n166 VSUBS 0.007859f
C1082 B.n167 VSUBS 0.007859f
C1083 B.n168 VSUBS 0.007859f
C1084 B.n169 VSUBS 0.007859f
C1085 B.t2 VSUBS 0.35944f
C1086 B.t1 VSUBS 0.398869f
C1087 B.t0 VSUBS 2.32891f
C1088 B.n170 VSUBS 0.61926f
C1089 B.n171 VSUBS 0.352633f
C1090 B.n172 VSUBS 0.007859f
C1091 B.n173 VSUBS 0.007859f
C1092 B.n174 VSUBS 0.007859f
C1093 B.n175 VSUBS 0.007859f
C1094 B.n176 VSUBS 0.007859f
C1095 B.n177 VSUBS 0.007859f
C1096 B.n178 VSUBS 0.007859f
C1097 B.n179 VSUBS 0.007859f
C1098 B.n180 VSUBS 0.007859f
C1099 B.n181 VSUBS 0.007859f
C1100 B.n182 VSUBS 0.007859f
C1101 B.n183 VSUBS 0.007859f
C1102 B.n184 VSUBS 0.007859f
C1103 B.n185 VSUBS 0.007859f
C1104 B.n186 VSUBS 0.007859f
C1105 B.n187 VSUBS 0.007859f
C1106 B.n188 VSUBS 0.007859f
C1107 B.n189 VSUBS 0.007859f
C1108 B.n190 VSUBS 0.007859f
C1109 B.n191 VSUBS 0.007859f
C1110 B.n192 VSUBS 0.007859f
C1111 B.n193 VSUBS 0.007859f
C1112 B.n194 VSUBS 0.007859f
C1113 B.n195 VSUBS 0.007859f
C1114 B.n196 VSUBS 0.007859f
C1115 B.n197 VSUBS 0.007859f
C1116 B.n198 VSUBS 0.007859f
C1117 B.n199 VSUBS 0.017097f
C1118 B.n200 VSUBS 0.007859f
C1119 B.n201 VSUBS 0.007859f
C1120 B.n202 VSUBS 0.007859f
C1121 B.n203 VSUBS 0.007859f
C1122 B.n204 VSUBS 0.007859f
C1123 B.n205 VSUBS 0.007859f
C1124 B.n206 VSUBS 0.007859f
C1125 B.n207 VSUBS 0.007859f
C1126 B.n208 VSUBS 0.007859f
C1127 B.n209 VSUBS 0.007859f
C1128 B.n210 VSUBS 0.007859f
C1129 B.n211 VSUBS 0.007859f
C1130 B.n212 VSUBS 0.007859f
C1131 B.n213 VSUBS 0.007859f
C1132 B.n214 VSUBS 0.007859f
C1133 B.n215 VSUBS 0.007859f
C1134 B.n216 VSUBS 0.007859f
C1135 B.n217 VSUBS 0.007859f
C1136 B.n218 VSUBS 0.007859f
C1137 B.n219 VSUBS 0.007859f
C1138 B.n220 VSUBS 0.007859f
C1139 B.n221 VSUBS 0.007859f
C1140 B.n222 VSUBS 0.007859f
C1141 B.n223 VSUBS 0.007859f
C1142 B.n224 VSUBS 0.007859f
C1143 B.n225 VSUBS 0.007859f
C1144 B.n226 VSUBS 0.007859f
C1145 B.n227 VSUBS 0.007859f
C1146 B.n228 VSUBS 0.007859f
C1147 B.n229 VSUBS 0.007859f
C1148 B.n230 VSUBS 0.007859f
C1149 B.n231 VSUBS 0.007859f
C1150 B.n232 VSUBS 0.007859f
C1151 B.n233 VSUBS 0.007859f
C1152 B.n234 VSUBS 0.007859f
C1153 B.n235 VSUBS 0.007859f
C1154 B.n236 VSUBS 0.007859f
C1155 B.n237 VSUBS 0.007859f
C1156 B.n238 VSUBS 0.007859f
C1157 B.n239 VSUBS 0.007859f
C1158 B.n240 VSUBS 0.007859f
C1159 B.n241 VSUBS 0.007859f
C1160 B.n242 VSUBS 0.007859f
C1161 B.n243 VSUBS 0.007859f
C1162 B.n244 VSUBS 0.007859f
C1163 B.n245 VSUBS 0.007859f
C1164 B.n246 VSUBS 0.007859f
C1165 B.n247 VSUBS 0.007859f
C1166 B.n248 VSUBS 0.007859f
C1167 B.n249 VSUBS 0.007859f
C1168 B.n250 VSUBS 0.007859f
C1169 B.n251 VSUBS 0.007859f
C1170 B.n252 VSUBS 0.007859f
C1171 B.n253 VSUBS 0.007859f
C1172 B.n254 VSUBS 0.007859f
C1173 B.n255 VSUBS 0.007859f
C1174 B.n256 VSUBS 0.007859f
C1175 B.n257 VSUBS 0.007859f
C1176 B.n258 VSUBS 0.007859f
C1177 B.n259 VSUBS 0.007859f
C1178 B.n260 VSUBS 0.007859f
C1179 B.n261 VSUBS 0.007859f
C1180 B.n262 VSUBS 0.007859f
C1181 B.n263 VSUBS 0.007859f
C1182 B.n264 VSUBS 0.007859f
C1183 B.n265 VSUBS 0.007859f
C1184 B.n266 VSUBS 0.007859f
C1185 B.n267 VSUBS 0.007859f
C1186 B.n268 VSUBS 0.007859f
C1187 B.n269 VSUBS 0.007859f
C1188 B.n270 VSUBS 0.007859f
C1189 B.n271 VSUBS 0.007859f
C1190 B.n272 VSUBS 0.007859f
C1191 B.n273 VSUBS 0.007859f
C1192 B.n274 VSUBS 0.007859f
C1193 B.n275 VSUBS 0.007859f
C1194 B.n276 VSUBS 0.007859f
C1195 B.n277 VSUBS 0.007859f
C1196 B.n278 VSUBS 0.007859f
C1197 B.n279 VSUBS 0.007859f
C1198 B.n280 VSUBS 0.007859f
C1199 B.n281 VSUBS 0.007859f
C1200 B.n282 VSUBS 0.007859f
C1201 B.n283 VSUBS 0.007859f
C1202 B.n284 VSUBS 0.017097f
C1203 B.n285 VSUBS 0.018502f
C1204 B.n286 VSUBS 0.018502f
C1205 B.n287 VSUBS 0.007859f
C1206 B.n288 VSUBS 0.007859f
C1207 B.n289 VSUBS 0.007859f
C1208 B.n290 VSUBS 0.007859f
C1209 B.n291 VSUBS 0.007859f
C1210 B.n292 VSUBS 0.007859f
C1211 B.n293 VSUBS 0.007859f
C1212 B.n294 VSUBS 0.007859f
C1213 B.n295 VSUBS 0.007859f
C1214 B.n296 VSUBS 0.007859f
C1215 B.n297 VSUBS 0.007859f
C1216 B.n298 VSUBS 0.007859f
C1217 B.n299 VSUBS 0.007859f
C1218 B.n300 VSUBS 0.007859f
C1219 B.n301 VSUBS 0.007859f
C1220 B.n302 VSUBS 0.007859f
C1221 B.n303 VSUBS 0.007859f
C1222 B.n304 VSUBS 0.007859f
C1223 B.n305 VSUBS 0.007859f
C1224 B.n306 VSUBS 0.007859f
C1225 B.n307 VSUBS 0.007859f
C1226 B.n308 VSUBS 0.007859f
C1227 B.n309 VSUBS 0.007859f
C1228 B.n310 VSUBS 0.007859f
C1229 B.n311 VSUBS 0.007859f
C1230 B.n312 VSUBS 0.007859f
C1231 B.n313 VSUBS 0.007859f
C1232 B.n314 VSUBS 0.007859f
C1233 B.n315 VSUBS 0.007859f
C1234 B.n316 VSUBS 0.007859f
C1235 B.n317 VSUBS 0.007859f
C1236 B.n318 VSUBS 0.007859f
C1237 B.n319 VSUBS 0.007859f
C1238 B.n320 VSUBS 0.007859f
C1239 B.n321 VSUBS 0.007859f
C1240 B.n322 VSUBS 0.007859f
C1241 B.n323 VSUBS 0.007859f
C1242 B.n324 VSUBS 0.007859f
C1243 B.n325 VSUBS 0.007859f
C1244 B.n326 VSUBS 0.007859f
C1245 B.n327 VSUBS 0.007859f
C1246 B.n328 VSUBS 0.007859f
C1247 B.n329 VSUBS 0.007859f
C1248 B.n330 VSUBS 0.007859f
C1249 B.n331 VSUBS 0.007859f
C1250 B.n332 VSUBS 0.007859f
C1251 B.n333 VSUBS 0.007859f
C1252 B.n334 VSUBS 0.007859f
C1253 B.n335 VSUBS 0.007859f
C1254 B.n336 VSUBS 0.007859f
C1255 B.n337 VSUBS 0.007859f
C1256 B.n338 VSUBS 0.007859f
C1257 B.n339 VSUBS 0.007859f
C1258 B.n340 VSUBS 0.007859f
C1259 B.n341 VSUBS 0.007859f
C1260 B.n342 VSUBS 0.007859f
C1261 B.n343 VSUBS 0.007859f
C1262 B.n344 VSUBS 0.007859f
C1263 B.n345 VSUBS 0.007859f
C1264 B.n346 VSUBS 0.007859f
C1265 B.n347 VSUBS 0.007859f
C1266 B.n348 VSUBS 0.007859f
C1267 B.n349 VSUBS 0.007859f
C1268 B.n350 VSUBS 0.007859f
C1269 B.n351 VSUBS 0.007859f
C1270 B.n352 VSUBS 0.007859f
C1271 B.n353 VSUBS 0.007859f
C1272 B.n354 VSUBS 0.007859f
C1273 B.n355 VSUBS 0.007859f
C1274 B.n356 VSUBS 0.007859f
C1275 B.n357 VSUBS 0.007859f
C1276 B.n358 VSUBS 0.007859f
C1277 B.n359 VSUBS 0.007859f
C1278 B.n360 VSUBS 0.007859f
C1279 B.n361 VSUBS 0.007859f
C1280 B.n362 VSUBS 0.007859f
C1281 B.n363 VSUBS 0.007859f
C1282 B.n364 VSUBS 0.007859f
C1283 B.n365 VSUBS 0.007859f
C1284 B.n366 VSUBS 0.007859f
C1285 B.n367 VSUBS 0.007859f
C1286 B.n368 VSUBS 0.005432f
C1287 B.n369 VSUBS 0.018209f
C1288 B.n370 VSUBS 0.006357f
C1289 B.n371 VSUBS 0.007859f
C1290 B.n372 VSUBS 0.007859f
C1291 B.n373 VSUBS 0.007859f
C1292 B.n374 VSUBS 0.007859f
C1293 B.n375 VSUBS 0.007859f
C1294 B.n376 VSUBS 0.007859f
C1295 B.n377 VSUBS 0.007859f
C1296 B.n378 VSUBS 0.007859f
C1297 B.n379 VSUBS 0.007859f
C1298 B.n380 VSUBS 0.007859f
C1299 B.n381 VSUBS 0.007859f
C1300 B.n382 VSUBS 0.006357f
C1301 B.n383 VSUBS 0.007859f
C1302 B.n384 VSUBS 0.007859f
C1303 B.n385 VSUBS 0.005432f
C1304 B.n386 VSUBS 0.007859f
C1305 B.n387 VSUBS 0.007859f
C1306 B.n388 VSUBS 0.007859f
C1307 B.n389 VSUBS 0.007859f
C1308 B.n390 VSUBS 0.007859f
C1309 B.n391 VSUBS 0.007859f
C1310 B.n392 VSUBS 0.007859f
C1311 B.n393 VSUBS 0.007859f
C1312 B.n394 VSUBS 0.007859f
C1313 B.n395 VSUBS 0.007859f
C1314 B.n396 VSUBS 0.007859f
C1315 B.n397 VSUBS 0.007859f
C1316 B.n398 VSUBS 0.007859f
C1317 B.n399 VSUBS 0.007859f
C1318 B.n400 VSUBS 0.007859f
C1319 B.n401 VSUBS 0.007859f
C1320 B.n402 VSUBS 0.007859f
C1321 B.n403 VSUBS 0.007859f
C1322 B.n404 VSUBS 0.007859f
C1323 B.n405 VSUBS 0.007859f
C1324 B.n406 VSUBS 0.007859f
C1325 B.n407 VSUBS 0.007859f
C1326 B.n408 VSUBS 0.007859f
C1327 B.n409 VSUBS 0.007859f
C1328 B.n410 VSUBS 0.007859f
C1329 B.n411 VSUBS 0.007859f
C1330 B.n412 VSUBS 0.007859f
C1331 B.n413 VSUBS 0.007859f
C1332 B.n414 VSUBS 0.007859f
C1333 B.n415 VSUBS 0.007859f
C1334 B.n416 VSUBS 0.007859f
C1335 B.n417 VSUBS 0.007859f
C1336 B.n418 VSUBS 0.007859f
C1337 B.n419 VSUBS 0.007859f
C1338 B.n420 VSUBS 0.007859f
C1339 B.n421 VSUBS 0.007859f
C1340 B.n422 VSUBS 0.007859f
C1341 B.n423 VSUBS 0.007859f
C1342 B.n424 VSUBS 0.007859f
C1343 B.n425 VSUBS 0.007859f
C1344 B.n426 VSUBS 0.007859f
C1345 B.n427 VSUBS 0.007859f
C1346 B.n428 VSUBS 0.007859f
C1347 B.n429 VSUBS 0.007859f
C1348 B.n430 VSUBS 0.007859f
C1349 B.n431 VSUBS 0.007859f
C1350 B.n432 VSUBS 0.007859f
C1351 B.n433 VSUBS 0.007859f
C1352 B.n434 VSUBS 0.007859f
C1353 B.n435 VSUBS 0.007859f
C1354 B.n436 VSUBS 0.007859f
C1355 B.n437 VSUBS 0.007859f
C1356 B.n438 VSUBS 0.007859f
C1357 B.n439 VSUBS 0.007859f
C1358 B.n440 VSUBS 0.007859f
C1359 B.n441 VSUBS 0.007859f
C1360 B.n442 VSUBS 0.007859f
C1361 B.n443 VSUBS 0.007859f
C1362 B.n444 VSUBS 0.007859f
C1363 B.n445 VSUBS 0.007859f
C1364 B.n446 VSUBS 0.007859f
C1365 B.n447 VSUBS 0.007859f
C1366 B.n448 VSUBS 0.007859f
C1367 B.n449 VSUBS 0.007859f
C1368 B.n450 VSUBS 0.007859f
C1369 B.n451 VSUBS 0.007859f
C1370 B.n452 VSUBS 0.007859f
C1371 B.n453 VSUBS 0.007859f
C1372 B.n454 VSUBS 0.007859f
C1373 B.n455 VSUBS 0.007859f
C1374 B.n456 VSUBS 0.007859f
C1375 B.n457 VSUBS 0.007859f
C1376 B.n458 VSUBS 0.007859f
C1377 B.n459 VSUBS 0.007859f
C1378 B.n460 VSUBS 0.007859f
C1379 B.n461 VSUBS 0.007859f
C1380 B.n462 VSUBS 0.007859f
C1381 B.n463 VSUBS 0.007859f
C1382 B.n464 VSUBS 0.007859f
C1383 B.n465 VSUBS 0.007859f
C1384 B.n466 VSUBS 0.007859f
C1385 B.n467 VSUBS 0.018502f
C1386 B.n468 VSUBS 0.017097f
C1387 B.n469 VSUBS 0.018073f
C1388 B.n470 VSUBS 0.007859f
C1389 B.n471 VSUBS 0.007859f
C1390 B.n472 VSUBS 0.007859f
C1391 B.n473 VSUBS 0.007859f
C1392 B.n474 VSUBS 0.007859f
C1393 B.n475 VSUBS 0.007859f
C1394 B.n476 VSUBS 0.007859f
C1395 B.n477 VSUBS 0.007859f
C1396 B.n478 VSUBS 0.007859f
C1397 B.n479 VSUBS 0.007859f
C1398 B.n480 VSUBS 0.007859f
C1399 B.n481 VSUBS 0.007859f
C1400 B.n482 VSUBS 0.007859f
C1401 B.n483 VSUBS 0.007859f
C1402 B.n484 VSUBS 0.007859f
C1403 B.n485 VSUBS 0.007859f
C1404 B.n486 VSUBS 0.007859f
C1405 B.n487 VSUBS 0.007859f
C1406 B.n488 VSUBS 0.007859f
C1407 B.n489 VSUBS 0.007859f
C1408 B.n490 VSUBS 0.007859f
C1409 B.n491 VSUBS 0.007859f
C1410 B.n492 VSUBS 0.007859f
C1411 B.n493 VSUBS 0.007859f
C1412 B.n494 VSUBS 0.007859f
C1413 B.n495 VSUBS 0.007859f
C1414 B.n496 VSUBS 0.007859f
C1415 B.n497 VSUBS 0.007859f
C1416 B.n498 VSUBS 0.007859f
C1417 B.n499 VSUBS 0.007859f
C1418 B.n500 VSUBS 0.007859f
C1419 B.n501 VSUBS 0.007859f
C1420 B.n502 VSUBS 0.007859f
C1421 B.n503 VSUBS 0.007859f
C1422 B.n504 VSUBS 0.007859f
C1423 B.n505 VSUBS 0.007859f
C1424 B.n506 VSUBS 0.007859f
C1425 B.n507 VSUBS 0.007859f
C1426 B.n508 VSUBS 0.007859f
C1427 B.n509 VSUBS 0.007859f
C1428 B.n510 VSUBS 0.007859f
C1429 B.n511 VSUBS 0.007859f
C1430 B.n512 VSUBS 0.007859f
C1431 B.n513 VSUBS 0.007859f
C1432 B.n514 VSUBS 0.007859f
C1433 B.n515 VSUBS 0.007859f
C1434 B.n516 VSUBS 0.007859f
C1435 B.n517 VSUBS 0.007859f
C1436 B.n518 VSUBS 0.007859f
C1437 B.n519 VSUBS 0.007859f
C1438 B.n520 VSUBS 0.007859f
C1439 B.n521 VSUBS 0.007859f
C1440 B.n522 VSUBS 0.007859f
C1441 B.n523 VSUBS 0.007859f
C1442 B.n524 VSUBS 0.007859f
C1443 B.n525 VSUBS 0.007859f
C1444 B.n526 VSUBS 0.007859f
C1445 B.n527 VSUBS 0.007859f
C1446 B.n528 VSUBS 0.007859f
C1447 B.n529 VSUBS 0.007859f
C1448 B.n530 VSUBS 0.007859f
C1449 B.n531 VSUBS 0.007859f
C1450 B.n532 VSUBS 0.007859f
C1451 B.n533 VSUBS 0.007859f
C1452 B.n534 VSUBS 0.007859f
C1453 B.n535 VSUBS 0.007859f
C1454 B.n536 VSUBS 0.007859f
C1455 B.n537 VSUBS 0.007859f
C1456 B.n538 VSUBS 0.007859f
C1457 B.n539 VSUBS 0.007859f
C1458 B.n540 VSUBS 0.007859f
C1459 B.n541 VSUBS 0.007859f
C1460 B.n542 VSUBS 0.007859f
C1461 B.n543 VSUBS 0.007859f
C1462 B.n544 VSUBS 0.007859f
C1463 B.n545 VSUBS 0.007859f
C1464 B.n546 VSUBS 0.007859f
C1465 B.n547 VSUBS 0.007859f
C1466 B.n548 VSUBS 0.007859f
C1467 B.n549 VSUBS 0.007859f
C1468 B.n550 VSUBS 0.007859f
C1469 B.n551 VSUBS 0.007859f
C1470 B.n552 VSUBS 0.007859f
C1471 B.n553 VSUBS 0.007859f
C1472 B.n554 VSUBS 0.007859f
C1473 B.n555 VSUBS 0.007859f
C1474 B.n556 VSUBS 0.007859f
C1475 B.n557 VSUBS 0.007859f
C1476 B.n558 VSUBS 0.007859f
C1477 B.n559 VSUBS 0.007859f
C1478 B.n560 VSUBS 0.007859f
C1479 B.n561 VSUBS 0.007859f
C1480 B.n562 VSUBS 0.007859f
C1481 B.n563 VSUBS 0.007859f
C1482 B.n564 VSUBS 0.007859f
C1483 B.n565 VSUBS 0.007859f
C1484 B.n566 VSUBS 0.007859f
C1485 B.n567 VSUBS 0.007859f
C1486 B.n568 VSUBS 0.007859f
C1487 B.n569 VSUBS 0.007859f
C1488 B.n570 VSUBS 0.007859f
C1489 B.n571 VSUBS 0.007859f
C1490 B.n572 VSUBS 0.007859f
C1491 B.n573 VSUBS 0.007859f
C1492 B.n574 VSUBS 0.007859f
C1493 B.n575 VSUBS 0.007859f
C1494 B.n576 VSUBS 0.007859f
C1495 B.n577 VSUBS 0.007859f
C1496 B.n578 VSUBS 0.007859f
C1497 B.n579 VSUBS 0.007859f
C1498 B.n580 VSUBS 0.007859f
C1499 B.n581 VSUBS 0.007859f
C1500 B.n582 VSUBS 0.007859f
C1501 B.n583 VSUBS 0.007859f
C1502 B.n584 VSUBS 0.007859f
C1503 B.n585 VSUBS 0.007859f
C1504 B.n586 VSUBS 0.007859f
C1505 B.n587 VSUBS 0.007859f
C1506 B.n588 VSUBS 0.007859f
C1507 B.n589 VSUBS 0.007859f
C1508 B.n590 VSUBS 0.007859f
C1509 B.n591 VSUBS 0.007859f
C1510 B.n592 VSUBS 0.007859f
C1511 B.n593 VSUBS 0.007859f
C1512 B.n594 VSUBS 0.007859f
C1513 B.n595 VSUBS 0.007859f
C1514 B.n596 VSUBS 0.007859f
C1515 B.n597 VSUBS 0.007859f
C1516 B.n598 VSUBS 0.007859f
C1517 B.n599 VSUBS 0.007859f
C1518 B.n600 VSUBS 0.007859f
C1519 B.n601 VSUBS 0.007859f
C1520 B.n602 VSUBS 0.017097f
C1521 B.n603 VSUBS 0.018502f
C1522 B.n604 VSUBS 0.018502f
C1523 B.n605 VSUBS 0.007859f
C1524 B.n606 VSUBS 0.007859f
C1525 B.n607 VSUBS 0.007859f
C1526 B.n608 VSUBS 0.007859f
C1527 B.n609 VSUBS 0.007859f
C1528 B.n610 VSUBS 0.007859f
C1529 B.n611 VSUBS 0.007859f
C1530 B.n612 VSUBS 0.007859f
C1531 B.n613 VSUBS 0.007859f
C1532 B.n614 VSUBS 0.007859f
C1533 B.n615 VSUBS 0.007859f
C1534 B.n616 VSUBS 0.007859f
C1535 B.n617 VSUBS 0.007859f
C1536 B.n618 VSUBS 0.007859f
C1537 B.n619 VSUBS 0.007859f
C1538 B.n620 VSUBS 0.007859f
C1539 B.n621 VSUBS 0.007859f
C1540 B.n622 VSUBS 0.007859f
C1541 B.n623 VSUBS 0.007859f
C1542 B.n624 VSUBS 0.007859f
C1543 B.n625 VSUBS 0.007859f
C1544 B.n626 VSUBS 0.007859f
C1545 B.n627 VSUBS 0.007859f
C1546 B.n628 VSUBS 0.007859f
C1547 B.n629 VSUBS 0.007859f
C1548 B.n630 VSUBS 0.007859f
C1549 B.n631 VSUBS 0.007859f
C1550 B.n632 VSUBS 0.007859f
C1551 B.n633 VSUBS 0.007859f
C1552 B.n634 VSUBS 0.007859f
C1553 B.n635 VSUBS 0.007859f
C1554 B.n636 VSUBS 0.007859f
C1555 B.n637 VSUBS 0.007859f
C1556 B.n638 VSUBS 0.007859f
C1557 B.n639 VSUBS 0.007859f
C1558 B.n640 VSUBS 0.007859f
C1559 B.n641 VSUBS 0.007859f
C1560 B.n642 VSUBS 0.007859f
C1561 B.n643 VSUBS 0.007859f
C1562 B.n644 VSUBS 0.007859f
C1563 B.n645 VSUBS 0.007859f
C1564 B.n646 VSUBS 0.007859f
C1565 B.n647 VSUBS 0.007859f
C1566 B.n648 VSUBS 0.007859f
C1567 B.n649 VSUBS 0.007859f
C1568 B.n650 VSUBS 0.007859f
C1569 B.n651 VSUBS 0.007859f
C1570 B.n652 VSUBS 0.007859f
C1571 B.n653 VSUBS 0.007859f
C1572 B.n654 VSUBS 0.007859f
C1573 B.n655 VSUBS 0.007859f
C1574 B.n656 VSUBS 0.007859f
C1575 B.n657 VSUBS 0.007859f
C1576 B.n658 VSUBS 0.007859f
C1577 B.n659 VSUBS 0.007859f
C1578 B.n660 VSUBS 0.007859f
C1579 B.n661 VSUBS 0.007859f
C1580 B.n662 VSUBS 0.007859f
C1581 B.n663 VSUBS 0.007859f
C1582 B.n664 VSUBS 0.007859f
C1583 B.n665 VSUBS 0.007859f
C1584 B.n666 VSUBS 0.007859f
C1585 B.n667 VSUBS 0.007859f
C1586 B.n668 VSUBS 0.007859f
C1587 B.n669 VSUBS 0.007859f
C1588 B.n670 VSUBS 0.007859f
C1589 B.n671 VSUBS 0.007859f
C1590 B.n672 VSUBS 0.007859f
C1591 B.n673 VSUBS 0.007859f
C1592 B.n674 VSUBS 0.007859f
C1593 B.n675 VSUBS 0.007859f
C1594 B.n676 VSUBS 0.007859f
C1595 B.n677 VSUBS 0.007859f
C1596 B.n678 VSUBS 0.007859f
C1597 B.n679 VSUBS 0.007859f
C1598 B.n680 VSUBS 0.007859f
C1599 B.n681 VSUBS 0.007859f
C1600 B.n682 VSUBS 0.007859f
C1601 B.n683 VSUBS 0.007859f
C1602 B.n684 VSUBS 0.007859f
C1603 B.n685 VSUBS 0.007859f
C1604 B.n686 VSUBS 0.005432f
C1605 B.n687 VSUBS 0.018209f
C1606 B.n688 VSUBS 0.006357f
C1607 B.n689 VSUBS 0.007859f
C1608 B.n690 VSUBS 0.007859f
C1609 B.n691 VSUBS 0.007859f
C1610 B.n692 VSUBS 0.007859f
C1611 B.n693 VSUBS 0.007859f
C1612 B.n694 VSUBS 0.007859f
C1613 B.n695 VSUBS 0.007859f
C1614 B.n696 VSUBS 0.007859f
C1615 B.n697 VSUBS 0.007859f
C1616 B.n698 VSUBS 0.007859f
C1617 B.n699 VSUBS 0.007859f
C1618 B.n700 VSUBS 0.006357f
C1619 B.n701 VSUBS 0.007859f
C1620 B.n702 VSUBS 0.007859f
C1621 B.n703 VSUBS 0.005432f
C1622 B.n704 VSUBS 0.007859f
C1623 B.n705 VSUBS 0.007859f
C1624 B.n706 VSUBS 0.007859f
C1625 B.n707 VSUBS 0.007859f
C1626 B.n708 VSUBS 0.007859f
C1627 B.n709 VSUBS 0.007859f
C1628 B.n710 VSUBS 0.007859f
C1629 B.n711 VSUBS 0.007859f
C1630 B.n712 VSUBS 0.007859f
C1631 B.n713 VSUBS 0.007859f
C1632 B.n714 VSUBS 0.007859f
C1633 B.n715 VSUBS 0.007859f
C1634 B.n716 VSUBS 0.007859f
C1635 B.n717 VSUBS 0.007859f
C1636 B.n718 VSUBS 0.007859f
C1637 B.n719 VSUBS 0.007859f
C1638 B.n720 VSUBS 0.007859f
C1639 B.n721 VSUBS 0.007859f
C1640 B.n722 VSUBS 0.007859f
C1641 B.n723 VSUBS 0.007859f
C1642 B.n724 VSUBS 0.007859f
C1643 B.n725 VSUBS 0.007859f
C1644 B.n726 VSUBS 0.007859f
C1645 B.n727 VSUBS 0.007859f
C1646 B.n728 VSUBS 0.007859f
C1647 B.n729 VSUBS 0.007859f
C1648 B.n730 VSUBS 0.007859f
C1649 B.n731 VSUBS 0.007859f
C1650 B.n732 VSUBS 0.007859f
C1651 B.n733 VSUBS 0.007859f
C1652 B.n734 VSUBS 0.007859f
C1653 B.n735 VSUBS 0.007859f
C1654 B.n736 VSUBS 0.007859f
C1655 B.n737 VSUBS 0.007859f
C1656 B.n738 VSUBS 0.007859f
C1657 B.n739 VSUBS 0.007859f
C1658 B.n740 VSUBS 0.007859f
C1659 B.n741 VSUBS 0.007859f
C1660 B.n742 VSUBS 0.007859f
C1661 B.n743 VSUBS 0.007859f
C1662 B.n744 VSUBS 0.007859f
C1663 B.n745 VSUBS 0.007859f
C1664 B.n746 VSUBS 0.007859f
C1665 B.n747 VSUBS 0.007859f
C1666 B.n748 VSUBS 0.007859f
C1667 B.n749 VSUBS 0.007859f
C1668 B.n750 VSUBS 0.007859f
C1669 B.n751 VSUBS 0.007859f
C1670 B.n752 VSUBS 0.007859f
C1671 B.n753 VSUBS 0.007859f
C1672 B.n754 VSUBS 0.007859f
C1673 B.n755 VSUBS 0.007859f
C1674 B.n756 VSUBS 0.007859f
C1675 B.n757 VSUBS 0.007859f
C1676 B.n758 VSUBS 0.007859f
C1677 B.n759 VSUBS 0.007859f
C1678 B.n760 VSUBS 0.007859f
C1679 B.n761 VSUBS 0.007859f
C1680 B.n762 VSUBS 0.007859f
C1681 B.n763 VSUBS 0.007859f
C1682 B.n764 VSUBS 0.007859f
C1683 B.n765 VSUBS 0.007859f
C1684 B.n766 VSUBS 0.007859f
C1685 B.n767 VSUBS 0.007859f
C1686 B.n768 VSUBS 0.007859f
C1687 B.n769 VSUBS 0.007859f
C1688 B.n770 VSUBS 0.007859f
C1689 B.n771 VSUBS 0.007859f
C1690 B.n772 VSUBS 0.007859f
C1691 B.n773 VSUBS 0.007859f
C1692 B.n774 VSUBS 0.007859f
C1693 B.n775 VSUBS 0.007859f
C1694 B.n776 VSUBS 0.007859f
C1695 B.n777 VSUBS 0.007859f
C1696 B.n778 VSUBS 0.007859f
C1697 B.n779 VSUBS 0.007859f
C1698 B.n780 VSUBS 0.007859f
C1699 B.n781 VSUBS 0.007859f
C1700 B.n782 VSUBS 0.007859f
C1701 B.n783 VSUBS 0.007859f
C1702 B.n784 VSUBS 0.007859f
C1703 B.n785 VSUBS 0.018502f
C1704 B.n786 VSUBS 0.017097f
C1705 B.n787 VSUBS 0.017097f
C1706 B.n788 VSUBS 0.007859f
C1707 B.n789 VSUBS 0.007859f
C1708 B.n790 VSUBS 0.007859f
C1709 B.n791 VSUBS 0.007859f
C1710 B.n792 VSUBS 0.007859f
C1711 B.n793 VSUBS 0.007859f
C1712 B.n794 VSUBS 0.007859f
C1713 B.n795 VSUBS 0.007859f
C1714 B.n796 VSUBS 0.007859f
C1715 B.n797 VSUBS 0.007859f
C1716 B.n798 VSUBS 0.007859f
C1717 B.n799 VSUBS 0.007859f
C1718 B.n800 VSUBS 0.007859f
C1719 B.n801 VSUBS 0.007859f
C1720 B.n802 VSUBS 0.007859f
C1721 B.n803 VSUBS 0.007859f
C1722 B.n804 VSUBS 0.007859f
C1723 B.n805 VSUBS 0.007859f
C1724 B.n806 VSUBS 0.007859f
C1725 B.n807 VSUBS 0.007859f
C1726 B.n808 VSUBS 0.007859f
C1727 B.n809 VSUBS 0.007859f
C1728 B.n810 VSUBS 0.007859f
C1729 B.n811 VSUBS 0.007859f
C1730 B.n812 VSUBS 0.007859f
C1731 B.n813 VSUBS 0.007859f
C1732 B.n814 VSUBS 0.007859f
C1733 B.n815 VSUBS 0.007859f
C1734 B.n816 VSUBS 0.007859f
C1735 B.n817 VSUBS 0.007859f
C1736 B.n818 VSUBS 0.007859f
C1737 B.n819 VSUBS 0.007859f
C1738 B.n820 VSUBS 0.007859f
C1739 B.n821 VSUBS 0.007859f
C1740 B.n822 VSUBS 0.007859f
C1741 B.n823 VSUBS 0.007859f
C1742 B.n824 VSUBS 0.007859f
C1743 B.n825 VSUBS 0.007859f
C1744 B.n826 VSUBS 0.007859f
C1745 B.n827 VSUBS 0.007859f
C1746 B.n828 VSUBS 0.007859f
C1747 B.n829 VSUBS 0.007859f
C1748 B.n830 VSUBS 0.007859f
C1749 B.n831 VSUBS 0.007859f
C1750 B.n832 VSUBS 0.007859f
C1751 B.n833 VSUBS 0.007859f
C1752 B.n834 VSUBS 0.007859f
C1753 B.n835 VSUBS 0.007859f
C1754 B.n836 VSUBS 0.007859f
C1755 B.n837 VSUBS 0.007859f
C1756 B.n838 VSUBS 0.007859f
C1757 B.n839 VSUBS 0.007859f
C1758 B.n840 VSUBS 0.007859f
C1759 B.n841 VSUBS 0.007859f
C1760 B.n842 VSUBS 0.007859f
C1761 B.n843 VSUBS 0.007859f
C1762 B.n844 VSUBS 0.007859f
C1763 B.n845 VSUBS 0.007859f
C1764 B.n846 VSUBS 0.007859f
C1765 B.n847 VSUBS 0.007859f
C1766 B.n848 VSUBS 0.007859f
C1767 B.n849 VSUBS 0.007859f
C1768 B.n850 VSUBS 0.007859f
C1769 B.n851 VSUBS 0.010256f
C1770 B.n852 VSUBS 0.010925f
C1771 B.n853 VSUBS 0.021726f
.ends

