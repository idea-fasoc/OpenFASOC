* NGSPICE file created from diff_pair_sample_0642.ext - technology: sky130A

.subckt diff_pair_sample_0642 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t12 VP.t0 VDD1.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=2.1483 pd=13.35 as=2.1483 ps=13.35 w=13.02 l=3.24
X1 VTAIL.t15 VN.t0 VDD2.t9 B.t21 sky130_fd_pr__nfet_01v8 ad=2.1483 pd=13.35 as=2.1483 ps=13.35 w=13.02 l=3.24
X2 VDD2.t8 VN.t1 VTAIL.t16 B.t22 sky130_fd_pr__nfet_01v8 ad=5.0778 pd=26.82 as=2.1483 ps=13.35 w=13.02 l=3.24
X3 B.t16 B.t14 B.t15 B.t4 sky130_fd_pr__nfet_01v8 ad=5.0778 pd=26.82 as=0 ps=0 w=13.02 l=3.24
X4 VDD1.t7 VP.t1 VTAIL.t11 B.t23 sky130_fd_pr__nfet_01v8 ad=2.1483 pd=13.35 as=2.1483 ps=13.35 w=13.02 l=3.24
X5 VDD1.t6 VP.t2 VTAIL.t10 B.t22 sky130_fd_pr__nfet_01v8 ad=5.0778 pd=26.82 as=2.1483 ps=13.35 w=13.02 l=3.24
X6 VDD1.t9 VP.t3 VTAIL.t9 B.t2 sky130_fd_pr__nfet_01v8 ad=2.1483 pd=13.35 as=5.0778 ps=26.82 w=13.02 l=3.24
X7 VDD2.t7 VN.t2 VTAIL.t19 B.t23 sky130_fd_pr__nfet_01v8 ad=2.1483 pd=13.35 as=2.1483 ps=13.35 w=13.02 l=3.24
X8 VDD2.t6 VN.t3 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.1483 pd=13.35 as=5.0778 ps=26.82 w=13.02 l=3.24
X9 VTAIL.t14 VN.t4 VDD2.t5 B.t17 sky130_fd_pr__nfet_01v8 ad=2.1483 pd=13.35 as=2.1483 ps=13.35 w=13.02 l=3.24
X10 VTAIL.t1 VN.t5 VDD2.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=2.1483 pd=13.35 as=2.1483 ps=13.35 w=13.02 l=3.24
X11 VTAIL.t8 VP.t4 VDD1.t8 B.t21 sky130_fd_pr__nfet_01v8 ad=2.1483 pd=13.35 as=2.1483 ps=13.35 w=13.02 l=3.24
X12 VDD2.t3 VN.t6 VTAIL.t13 B.t19 sky130_fd_pr__nfet_01v8 ad=2.1483 pd=13.35 as=5.0778 ps=26.82 w=13.02 l=3.24
X13 VTAIL.t7 VP.t5 VDD1.t3 B.t20 sky130_fd_pr__nfet_01v8 ad=2.1483 pd=13.35 as=2.1483 ps=13.35 w=13.02 l=3.24
X14 B.t13 B.t11 B.t12 B.t8 sky130_fd_pr__nfet_01v8 ad=5.0778 pd=26.82 as=0 ps=0 w=13.02 l=3.24
X15 VDD1.t2 VP.t6 VTAIL.t6 B.t19 sky130_fd_pr__nfet_01v8 ad=2.1483 pd=13.35 as=5.0778 ps=26.82 w=13.02 l=3.24
X16 VDD1.t5 VP.t7 VTAIL.t5 B.t18 sky130_fd_pr__nfet_01v8 ad=2.1483 pd=13.35 as=2.1483 ps=13.35 w=13.02 l=3.24
X17 B.t10 B.t7 B.t9 B.t8 sky130_fd_pr__nfet_01v8 ad=5.0778 pd=26.82 as=0 ps=0 w=13.02 l=3.24
X18 B.t6 B.t3 B.t5 B.t4 sky130_fd_pr__nfet_01v8 ad=5.0778 pd=26.82 as=0 ps=0 w=13.02 l=3.24
X19 VDD1.t4 VP.t8 VTAIL.t4 B.t0 sky130_fd_pr__nfet_01v8 ad=5.0778 pd=26.82 as=2.1483 ps=13.35 w=13.02 l=3.24
X20 VDD2.t2 VN.t7 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=5.0778 pd=26.82 as=2.1483 ps=13.35 w=13.02 l=3.24
X21 VDD2.t1 VN.t8 VTAIL.t18 B.t18 sky130_fd_pr__nfet_01v8 ad=2.1483 pd=13.35 as=2.1483 ps=13.35 w=13.02 l=3.24
X22 VTAIL.t3 VP.t9 VDD1.t1 B.t17 sky130_fd_pr__nfet_01v8 ad=2.1483 pd=13.35 as=2.1483 ps=13.35 w=13.02 l=3.24
X23 VTAIL.t17 VN.t9 VDD2.t0 B.t20 sky130_fd_pr__nfet_01v8 ad=2.1483 pd=13.35 as=2.1483 ps=13.35 w=13.02 l=3.24
R0 VP.n32 VP.n31 161.3
R1 VP.n33 VP.n28 161.3
R2 VP.n35 VP.n34 161.3
R3 VP.n36 VP.n27 161.3
R4 VP.n38 VP.n37 161.3
R5 VP.n39 VP.n26 161.3
R6 VP.n41 VP.n40 161.3
R7 VP.n43 VP.n42 161.3
R8 VP.n44 VP.n24 161.3
R9 VP.n46 VP.n45 161.3
R10 VP.n47 VP.n23 161.3
R11 VP.n49 VP.n48 161.3
R12 VP.n50 VP.n22 161.3
R13 VP.n52 VP.n51 161.3
R14 VP.n54 VP.n53 161.3
R15 VP.n55 VP.n20 161.3
R16 VP.n57 VP.n56 161.3
R17 VP.n58 VP.n19 161.3
R18 VP.n60 VP.n59 161.3
R19 VP.n61 VP.n18 161.3
R20 VP.n63 VP.n62 161.3
R21 VP.n109 VP.n108 161.3
R22 VP.n107 VP.n1 161.3
R23 VP.n106 VP.n105 161.3
R24 VP.n104 VP.n2 161.3
R25 VP.n103 VP.n102 161.3
R26 VP.n101 VP.n3 161.3
R27 VP.n100 VP.n99 161.3
R28 VP.n98 VP.n97 161.3
R29 VP.n96 VP.n5 161.3
R30 VP.n95 VP.n94 161.3
R31 VP.n93 VP.n6 161.3
R32 VP.n92 VP.n91 161.3
R33 VP.n90 VP.n7 161.3
R34 VP.n89 VP.n88 161.3
R35 VP.n87 VP.n86 161.3
R36 VP.n85 VP.n9 161.3
R37 VP.n84 VP.n83 161.3
R38 VP.n82 VP.n10 161.3
R39 VP.n81 VP.n80 161.3
R40 VP.n79 VP.n11 161.3
R41 VP.n78 VP.n77 161.3
R42 VP.n76 VP.n75 161.3
R43 VP.n74 VP.n13 161.3
R44 VP.n73 VP.n72 161.3
R45 VP.n71 VP.n14 161.3
R46 VP.n70 VP.n69 161.3
R47 VP.n68 VP.n15 161.3
R48 VP.n67 VP.n66 161.3
R49 VP.n30 VP.t2 130.256
R50 VP.n16 VP.t8 96.8468
R51 VP.n12 VP.t9 96.8468
R52 VP.n8 VP.t1 96.8468
R53 VP.n4 VP.t5 96.8468
R54 VP.n0 VP.t6 96.8468
R55 VP.n17 VP.t3 96.8468
R56 VP.n21 VP.t0 96.8468
R57 VP.n25 VP.t7 96.8468
R58 VP.n29 VP.t4 96.8468
R59 VP.n65 VP.n16 71.0639
R60 VP.n110 VP.n0 71.0639
R61 VP.n64 VP.n17 71.0639
R62 VP.n30 VP.n29 58.6193
R63 VP.n65 VP.n64 57.5336
R64 VP.n69 VP.n14 50.7491
R65 VP.n106 VP.n2 50.7491
R66 VP.n60 VP.n19 50.7491
R67 VP.n80 VP.n10 43.9677
R68 VP.n95 VP.n6 43.9677
R69 VP.n49 VP.n23 43.9677
R70 VP.n34 VP.n27 43.9677
R71 VP.n84 VP.n10 37.1863
R72 VP.n91 VP.n6 37.1863
R73 VP.n45 VP.n23 37.1863
R74 VP.n38 VP.n27 37.1863
R75 VP.n73 VP.n14 30.405
R76 VP.n102 VP.n2 30.405
R77 VP.n56 VP.n19 30.405
R78 VP.n68 VP.n67 24.5923
R79 VP.n69 VP.n68 24.5923
R80 VP.n74 VP.n73 24.5923
R81 VP.n75 VP.n74 24.5923
R82 VP.n79 VP.n78 24.5923
R83 VP.n80 VP.n79 24.5923
R84 VP.n85 VP.n84 24.5923
R85 VP.n86 VP.n85 24.5923
R86 VP.n90 VP.n89 24.5923
R87 VP.n91 VP.n90 24.5923
R88 VP.n96 VP.n95 24.5923
R89 VP.n97 VP.n96 24.5923
R90 VP.n101 VP.n100 24.5923
R91 VP.n102 VP.n101 24.5923
R92 VP.n107 VP.n106 24.5923
R93 VP.n108 VP.n107 24.5923
R94 VP.n61 VP.n60 24.5923
R95 VP.n62 VP.n61 24.5923
R96 VP.n50 VP.n49 24.5923
R97 VP.n51 VP.n50 24.5923
R98 VP.n55 VP.n54 24.5923
R99 VP.n56 VP.n55 24.5923
R100 VP.n39 VP.n38 24.5923
R101 VP.n40 VP.n39 24.5923
R102 VP.n44 VP.n43 24.5923
R103 VP.n45 VP.n44 24.5923
R104 VP.n33 VP.n32 24.5923
R105 VP.n34 VP.n33 24.5923
R106 VP.n67 VP.n16 19.1821
R107 VP.n108 VP.n0 19.1821
R108 VP.n62 VP.n17 19.1821
R109 VP.n78 VP.n12 15.7393
R110 VP.n97 VP.n4 15.7393
R111 VP.n51 VP.n21 15.7393
R112 VP.n32 VP.n29 15.7393
R113 VP.n86 VP.n8 12.2964
R114 VP.n89 VP.n8 12.2964
R115 VP.n40 VP.n25 12.2964
R116 VP.n43 VP.n25 12.2964
R117 VP.n75 VP.n12 8.85356
R118 VP.n100 VP.n4 8.85356
R119 VP.n54 VP.n21 8.85356
R120 VP.n31 VP.n30 3.93511
R121 VP.n64 VP.n63 0.354861
R122 VP.n66 VP.n65 0.354861
R123 VP.n110 VP.n109 0.354861
R124 VP VP.n110 0.267071
R125 VP.n31 VP.n28 0.189894
R126 VP.n35 VP.n28 0.189894
R127 VP.n36 VP.n35 0.189894
R128 VP.n37 VP.n36 0.189894
R129 VP.n37 VP.n26 0.189894
R130 VP.n41 VP.n26 0.189894
R131 VP.n42 VP.n41 0.189894
R132 VP.n42 VP.n24 0.189894
R133 VP.n46 VP.n24 0.189894
R134 VP.n47 VP.n46 0.189894
R135 VP.n48 VP.n47 0.189894
R136 VP.n48 VP.n22 0.189894
R137 VP.n52 VP.n22 0.189894
R138 VP.n53 VP.n52 0.189894
R139 VP.n53 VP.n20 0.189894
R140 VP.n57 VP.n20 0.189894
R141 VP.n58 VP.n57 0.189894
R142 VP.n59 VP.n58 0.189894
R143 VP.n59 VP.n18 0.189894
R144 VP.n63 VP.n18 0.189894
R145 VP.n66 VP.n15 0.189894
R146 VP.n70 VP.n15 0.189894
R147 VP.n71 VP.n70 0.189894
R148 VP.n72 VP.n71 0.189894
R149 VP.n72 VP.n13 0.189894
R150 VP.n76 VP.n13 0.189894
R151 VP.n77 VP.n76 0.189894
R152 VP.n77 VP.n11 0.189894
R153 VP.n81 VP.n11 0.189894
R154 VP.n82 VP.n81 0.189894
R155 VP.n83 VP.n82 0.189894
R156 VP.n83 VP.n9 0.189894
R157 VP.n87 VP.n9 0.189894
R158 VP.n88 VP.n87 0.189894
R159 VP.n88 VP.n7 0.189894
R160 VP.n92 VP.n7 0.189894
R161 VP.n93 VP.n92 0.189894
R162 VP.n94 VP.n93 0.189894
R163 VP.n94 VP.n5 0.189894
R164 VP.n98 VP.n5 0.189894
R165 VP.n99 VP.n98 0.189894
R166 VP.n99 VP.n3 0.189894
R167 VP.n103 VP.n3 0.189894
R168 VP.n104 VP.n103 0.189894
R169 VP.n105 VP.n104 0.189894
R170 VP.n105 VP.n1 0.189894
R171 VP.n109 VP.n1 0.189894
R172 VDD1.n1 VDD1.t6 69.2662
R173 VDD1.n3 VDD1.t4 69.265
R174 VDD1.n5 VDD1.n4 66.9195
R175 VDD1.n1 VDD1.n0 64.6679
R176 VDD1.n7 VDD1.n6 64.6667
R177 VDD1.n3 VDD1.n2 64.6667
R178 VDD1.n7 VDD1.n5 51.6798
R179 VDD1 VDD1.n7 2.2505
R180 VDD1.n6 VDD1.t0 1.52124
R181 VDD1.n6 VDD1.t9 1.52124
R182 VDD1.n0 VDD1.t8 1.52124
R183 VDD1.n0 VDD1.t5 1.52124
R184 VDD1.n4 VDD1.t3 1.52124
R185 VDD1.n4 VDD1.t2 1.52124
R186 VDD1.n2 VDD1.t1 1.52124
R187 VDD1.n2 VDD1.t7 1.52124
R188 VDD1 VDD1.n1 0.828086
R189 VDD1.n5 VDD1.n3 0.714551
R190 VTAIL.n11 VTAIL.t13 49.5098
R191 VTAIL.n17 VTAIL.t2 49.5087
R192 VTAIL.n2 VTAIL.t6 49.5087
R193 VTAIL.n16 VTAIL.t9 49.5087
R194 VTAIL.n15 VTAIL.n14 47.9891
R195 VTAIL.n13 VTAIL.n12 47.9891
R196 VTAIL.n10 VTAIL.n9 47.9891
R197 VTAIL.n8 VTAIL.n7 47.9891
R198 VTAIL.n19 VTAIL.n18 47.9879
R199 VTAIL.n1 VTAIL.n0 47.9879
R200 VTAIL.n4 VTAIL.n3 47.9879
R201 VTAIL.n6 VTAIL.n5 47.9879
R202 VTAIL.n8 VTAIL.n6 29.7462
R203 VTAIL.n17 VTAIL.n16 26.6686
R204 VTAIL.n10 VTAIL.n8 3.07809
R205 VTAIL.n11 VTAIL.n10 3.07809
R206 VTAIL.n15 VTAIL.n13 3.07809
R207 VTAIL.n16 VTAIL.n15 3.07809
R208 VTAIL.n6 VTAIL.n4 3.07809
R209 VTAIL.n4 VTAIL.n2 3.07809
R210 VTAIL.n19 VTAIL.n17 3.07809
R211 VTAIL VTAIL.n1 2.36688
R212 VTAIL.n13 VTAIL.n11 2.00912
R213 VTAIL.n2 VTAIL.n1 2.00912
R214 VTAIL.n18 VTAIL.t18 1.52124
R215 VTAIL.n18 VTAIL.t1 1.52124
R216 VTAIL.n0 VTAIL.t16 1.52124
R217 VTAIL.n0 VTAIL.t15 1.52124
R218 VTAIL.n3 VTAIL.t11 1.52124
R219 VTAIL.n3 VTAIL.t7 1.52124
R220 VTAIL.n5 VTAIL.t4 1.52124
R221 VTAIL.n5 VTAIL.t3 1.52124
R222 VTAIL.n14 VTAIL.t5 1.52124
R223 VTAIL.n14 VTAIL.t12 1.52124
R224 VTAIL.n12 VTAIL.t10 1.52124
R225 VTAIL.n12 VTAIL.t8 1.52124
R226 VTAIL.n9 VTAIL.t19 1.52124
R227 VTAIL.n9 VTAIL.t17 1.52124
R228 VTAIL.n7 VTAIL.t0 1.52124
R229 VTAIL.n7 VTAIL.t14 1.52124
R230 VTAIL VTAIL.n19 0.711707
R231 B.n1074 B.n1073 585
R232 B.n1075 B.n1074 585
R233 B.n377 B.n179 585
R234 B.n376 B.n375 585
R235 B.n374 B.n373 585
R236 B.n372 B.n371 585
R237 B.n370 B.n369 585
R238 B.n368 B.n367 585
R239 B.n366 B.n365 585
R240 B.n364 B.n363 585
R241 B.n362 B.n361 585
R242 B.n360 B.n359 585
R243 B.n358 B.n357 585
R244 B.n356 B.n355 585
R245 B.n354 B.n353 585
R246 B.n352 B.n351 585
R247 B.n350 B.n349 585
R248 B.n348 B.n347 585
R249 B.n346 B.n345 585
R250 B.n344 B.n343 585
R251 B.n342 B.n341 585
R252 B.n340 B.n339 585
R253 B.n338 B.n337 585
R254 B.n336 B.n335 585
R255 B.n334 B.n333 585
R256 B.n332 B.n331 585
R257 B.n330 B.n329 585
R258 B.n328 B.n327 585
R259 B.n326 B.n325 585
R260 B.n324 B.n323 585
R261 B.n322 B.n321 585
R262 B.n320 B.n319 585
R263 B.n318 B.n317 585
R264 B.n316 B.n315 585
R265 B.n314 B.n313 585
R266 B.n312 B.n311 585
R267 B.n310 B.n309 585
R268 B.n308 B.n307 585
R269 B.n306 B.n305 585
R270 B.n304 B.n303 585
R271 B.n302 B.n301 585
R272 B.n300 B.n299 585
R273 B.n298 B.n297 585
R274 B.n296 B.n295 585
R275 B.n294 B.n293 585
R276 B.n292 B.n291 585
R277 B.n290 B.n289 585
R278 B.n288 B.n287 585
R279 B.n286 B.n285 585
R280 B.n284 B.n283 585
R281 B.n282 B.n281 585
R282 B.n280 B.n279 585
R283 B.n278 B.n277 585
R284 B.n276 B.n275 585
R285 B.n274 B.n273 585
R286 B.n271 B.n270 585
R287 B.n269 B.n268 585
R288 B.n267 B.n266 585
R289 B.n265 B.n264 585
R290 B.n263 B.n262 585
R291 B.n261 B.n260 585
R292 B.n259 B.n258 585
R293 B.n257 B.n256 585
R294 B.n255 B.n254 585
R295 B.n253 B.n252 585
R296 B.n251 B.n250 585
R297 B.n249 B.n248 585
R298 B.n247 B.n246 585
R299 B.n245 B.n244 585
R300 B.n243 B.n242 585
R301 B.n241 B.n240 585
R302 B.n239 B.n238 585
R303 B.n237 B.n236 585
R304 B.n235 B.n234 585
R305 B.n233 B.n232 585
R306 B.n231 B.n230 585
R307 B.n229 B.n228 585
R308 B.n227 B.n226 585
R309 B.n225 B.n224 585
R310 B.n223 B.n222 585
R311 B.n221 B.n220 585
R312 B.n219 B.n218 585
R313 B.n217 B.n216 585
R314 B.n215 B.n214 585
R315 B.n213 B.n212 585
R316 B.n211 B.n210 585
R317 B.n209 B.n208 585
R318 B.n207 B.n206 585
R319 B.n205 B.n204 585
R320 B.n203 B.n202 585
R321 B.n201 B.n200 585
R322 B.n199 B.n198 585
R323 B.n197 B.n196 585
R324 B.n195 B.n194 585
R325 B.n193 B.n192 585
R326 B.n191 B.n190 585
R327 B.n189 B.n188 585
R328 B.n187 B.n186 585
R329 B.n130 B.n129 585
R330 B.n1078 B.n1077 585
R331 B.n1072 B.n180 585
R332 B.n180 B.n127 585
R333 B.n1071 B.n126 585
R334 B.n1082 B.n126 585
R335 B.n1070 B.n125 585
R336 B.n1083 B.n125 585
R337 B.n1069 B.n124 585
R338 B.n1084 B.n124 585
R339 B.n1068 B.n1067 585
R340 B.n1067 B.n120 585
R341 B.n1066 B.n119 585
R342 B.n1090 B.n119 585
R343 B.n1065 B.n118 585
R344 B.n1091 B.n118 585
R345 B.n1064 B.n117 585
R346 B.n1092 B.n117 585
R347 B.n1063 B.n1062 585
R348 B.n1062 B.n116 585
R349 B.n1061 B.n112 585
R350 B.n1098 B.n112 585
R351 B.n1060 B.n111 585
R352 B.n1099 B.n111 585
R353 B.n1059 B.n110 585
R354 B.n1100 B.n110 585
R355 B.n1058 B.n1057 585
R356 B.n1057 B.n106 585
R357 B.n1056 B.n105 585
R358 B.n1106 B.n105 585
R359 B.n1055 B.n104 585
R360 B.n1107 B.n104 585
R361 B.n1054 B.n103 585
R362 B.n1108 B.n103 585
R363 B.n1053 B.n1052 585
R364 B.n1052 B.n99 585
R365 B.n1051 B.n98 585
R366 B.n1114 B.n98 585
R367 B.n1050 B.n97 585
R368 B.n1115 B.n97 585
R369 B.n1049 B.n96 585
R370 B.n1116 B.n96 585
R371 B.n1048 B.n1047 585
R372 B.n1047 B.n92 585
R373 B.n1046 B.n91 585
R374 B.n1122 B.n91 585
R375 B.n1045 B.n90 585
R376 B.n1123 B.n90 585
R377 B.n1044 B.n89 585
R378 B.n1124 B.n89 585
R379 B.n1043 B.n1042 585
R380 B.n1042 B.n85 585
R381 B.n1041 B.n84 585
R382 B.n1130 B.n84 585
R383 B.n1040 B.n83 585
R384 B.n1131 B.n83 585
R385 B.n1039 B.n82 585
R386 B.n1132 B.n82 585
R387 B.n1038 B.n1037 585
R388 B.n1037 B.n78 585
R389 B.n1036 B.n77 585
R390 B.n1138 B.n77 585
R391 B.n1035 B.n76 585
R392 B.n1139 B.n76 585
R393 B.n1034 B.n75 585
R394 B.n1140 B.n75 585
R395 B.n1033 B.n1032 585
R396 B.n1032 B.n74 585
R397 B.n1031 B.n70 585
R398 B.n1146 B.n70 585
R399 B.n1030 B.n69 585
R400 B.n1147 B.n69 585
R401 B.n1029 B.n68 585
R402 B.n1148 B.n68 585
R403 B.n1028 B.n1027 585
R404 B.n1027 B.n64 585
R405 B.n1026 B.n63 585
R406 B.n1154 B.n63 585
R407 B.n1025 B.n62 585
R408 B.n1155 B.n62 585
R409 B.n1024 B.n61 585
R410 B.n1156 B.n61 585
R411 B.n1023 B.n1022 585
R412 B.n1022 B.n57 585
R413 B.n1021 B.n56 585
R414 B.n1162 B.n56 585
R415 B.n1020 B.n55 585
R416 B.n1163 B.n55 585
R417 B.n1019 B.n54 585
R418 B.n1164 B.n54 585
R419 B.n1018 B.n1017 585
R420 B.n1017 B.n50 585
R421 B.n1016 B.n49 585
R422 B.n1170 B.n49 585
R423 B.n1015 B.n48 585
R424 B.n1171 B.n48 585
R425 B.n1014 B.n47 585
R426 B.n1172 B.n47 585
R427 B.n1013 B.n1012 585
R428 B.n1012 B.n43 585
R429 B.n1011 B.n42 585
R430 B.n1178 B.n42 585
R431 B.n1010 B.n41 585
R432 B.n1179 B.n41 585
R433 B.n1009 B.n40 585
R434 B.n1180 B.n40 585
R435 B.n1008 B.n1007 585
R436 B.n1007 B.n36 585
R437 B.n1006 B.n35 585
R438 B.n1186 B.n35 585
R439 B.n1005 B.n34 585
R440 B.n1187 B.n34 585
R441 B.n1004 B.n33 585
R442 B.n1188 B.n33 585
R443 B.n1003 B.n1002 585
R444 B.n1002 B.n29 585
R445 B.n1001 B.n28 585
R446 B.n1194 B.n28 585
R447 B.n1000 B.n27 585
R448 B.n1195 B.n27 585
R449 B.n999 B.n26 585
R450 B.n1196 B.n26 585
R451 B.n998 B.n997 585
R452 B.n997 B.n22 585
R453 B.n996 B.n21 585
R454 B.n1202 B.n21 585
R455 B.n995 B.n20 585
R456 B.n1203 B.n20 585
R457 B.n994 B.n19 585
R458 B.n1204 B.n19 585
R459 B.n993 B.n992 585
R460 B.n992 B.n18 585
R461 B.n991 B.n14 585
R462 B.n1210 B.n14 585
R463 B.n990 B.n13 585
R464 B.n1211 B.n13 585
R465 B.n989 B.n12 585
R466 B.n1212 B.n12 585
R467 B.n988 B.n987 585
R468 B.n987 B.n8 585
R469 B.n986 B.n7 585
R470 B.n1218 B.n7 585
R471 B.n985 B.n6 585
R472 B.n1219 B.n6 585
R473 B.n984 B.n5 585
R474 B.n1220 B.n5 585
R475 B.n983 B.n982 585
R476 B.n982 B.n4 585
R477 B.n981 B.n378 585
R478 B.n981 B.n980 585
R479 B.n971 B.n379 585
R480 B.n380 B.n379 585
R481 B.n973 B.n972 585
R482 B.n974 B.n973 585
R483 B.n970 B.n385 585
R484 B.n385 B.n384 585
R485 B.n969 B.n968 585
R486 B.n968 B.n967 585
R487 B.n387 B.n386 585
R488 B.n960 B.n387 585
R489 B.n959 B.n958 585
R490 B.n961 B.n959 585
R491 B.n957 B.n392 585
R492 B.n392 B.n391 585
R493 B.n956 B.n955 585
R494 B.n955 B.n954 585
R495 B.n394 B.n393 585
R496 B.n395 B.n394 585
R497 B.n947 B.n946 585
R498 B.n948 B.n947 585
R499 B.n945 B.n400 585
R500 B.n400 B.n399 585
R501 B.n944 B.n943 585
R502 B.n943 B.n942 585
R503 B.n402 B.n401 585
R504 B.n403 B.n402 585
R505 B.n935 B.n934 585
R506 B.n936 B.n935 585
R507 B.n933 B.n408 585
R508 B.n408 B.n407 585
R509 B.n932 B.n931 585
R510 B.n931 B.n930 585
R511 B.n410 B.n409 585
R512 B.n411 B.n410 585
R513 B.n923 B.n922 585
R514 B.n924 B.n923 585
R515 B.n921 B.n416 585
R516 B.n416 B.n415 585
R517 B.n920 B.n919 585
R518 B.n919 B.n918 585
R519 B.n418 B.n417 585
R520 B.n419 B.n418 585
R521 B.n911 B.n910 585
R522 B.n912 B.n911 585
R523 B.n909 B.n424 585
R524 B.n424 B.n423 585
R525 B.n908 B.n907 585
R526 B.n907 B.n906 585
R527 B.n426 B.n425 585
R528 B.n427 B.n426 585
R529 B.n899 B.n898 585
R530 B.n900 B.n899 585
R531 B.n897 B.n432 585
R532 B.n432 B.n431 585
R533 B.n896 B.n895 585
R534 B.n895 B.n894 585
R535 B.n434 B.n433 585
R536 B.n435 B.n434 585
R537 B.n887 B.n886 585
R538 B.n888 B.n887 585
R539 B.n885 B.n440 585
R540 B.n440 B.n439 585
R541 B.n884 B.n883 585
R542 B.n883 B.n882 585
R543 B.n442 B.n441 585
R544 B.n443 B.n442 585
R545 B.n875 B.n874 585
R546 B.n876 B.n875 585
R547 B.n873 B.n448 585
R548 B.n448 B.n447 585
R549 B.n872 B.n871 585
R550 B.n871 B.n870 585
R551 B.n450 B.n449 585
R552 B.n863 B.n450 585
R553 B.n862 B.n861 585
R554 B.n864 B.n862 585
R555 B.n860 B.n455 585
R556 B.n455 B.n454 585
R557 B.n859 B.n858 585
R558 B.n858 B.n857 585
R559 B.n457 B.n456 585
R560 B.n458 B.n457 585
R561 B.n850 B.n849 585
R562 B.n851 B.n850 585
R563 B.n848 B.n463 585
R564 B.n463 B.n462 585
R565 B.n847 B.n846 585
R566 B.n846 B.n845 585
R567 B.n465 B.n464 585
R568 B.n466 B.n465 585
R569 B.n838 B.n837 585
R570 B.n839 B.n838 585
R571 B.n836 B.n470 585
R572 B.n474 B.n470 585
R573 B.n835 B.n834 585
R574 B.n834 B.n833 585
R575 B.n472 B.n471 585
R576 B.n473 B.n472 585
R577 B.n826 B.n825 585
R578 B.n827 B.n826 585
R579 B.n824 B.n479 585
R580 B.n479 B.n478 585
R581 B.n823 B.n822 585
R582 B.n822 B.n821 585
R583 B.n481 B.n480 585
R584 B.n482 B.n481 585
R585 B.n814 B.n813 585
R586 B.n815 B.n814 585
R587 B.n812 B.n487 585
R588 B.n487 B.n486 585
R589 B.n811 B.n810 585
R590 B.n810 B.n809 585
R591 B.n489 B.n488 585
R592 B.n490 B.n489 585
R593 B.n802 B.n801 585
R594 B.n803 B.n802 585
R595 B.n800 B.n495 585
R596 B.n495 B.n494 585
R597 B.n799 B.n798 585
R598 B.n798 B.n797 585
R599 B.n497 B.n496 585
R600 B.n790 B.n497 585
R601 B.n789 B.n788 585
R602 B.n791 B.n789 585
R603 B.n787 B.n502 585
R604 B.n502 B.n501 585
R605 B.n786 B.n785 585
R606 B.n785 B.n784 585
R607 B.n504 B.n503 585
R608 B.n505 B.n504 585
R609 B.n777 B.n776 585
R610 B.n778 B.n777 585
R611 B.n775 B.n510 585
R612 B.n510 B.n509 585
R613 B.n774 B.n773 585
R614 B.n773 B.n772 585
R615 B.n512 B.n511 585
R616 B.n513 B.n512 585
R617 B.n768 B.n767 585
R618 B.n516 B.n515 585
R619 B.n764 B.n763 585
R620 B.n765 B.n764 585
R621 B.n762 B.n565 585
R622 B.n761 B.n760 585
R623 B.n759 B.n758 585
R624 B.n757 B.n756 585
R625 B.n755 B.n754 585
R626 B.n753 B.n752 585
R627 B.n751 B.n750 585
R628 B.n749 B.n748 585
R629 B.n747 B.n746 585
R630 B.n745 B.n744 585
R631 B.n743 B.n742 585
R632 B.n741 B.n740 585
R633 B.n739 B.n738 585
R634 B.n737 B.n736 585
R635 B.n735 B.n734 585
R636 B.n733 B.n732 585
R637 B.n731 B.n730 585
R638 B.n729 B.n728 585
R639 B.n727 B.n726 585
R640 B.n725 B.n724 585
R641 B.n723 B.n722 585
R642 B.n721 B.n720 585
R643 B.n719 B.n718 585
R644 B.n717 B.n716 585
R645 B.n715 B.n714 585
R646 B.n713 B.n712 585
R647 B.n711 B.n710 585
R648 B.n709 B.n708 585
R649 B.n707 B.n706 585
R650 B.n705 B.n704 585
R651 B.n703 B.n702 585
R652 B.n701 B.n700 585
R653 B.n699 B.n698 585
R654 B.n697 B.n696 585
R655 B.n695 B.n694 585
R656 B.n693 B.n692 585
R657 B.n691 B.n690 585
R658 B.n689 B.n688 585
R659 B.n687 B.n686 585
R660 B.n685 B.n684 585
R661 B.n683 B.n682 585
R662 B.n681 B.n680 585
R663 B.n679 B.n678 585
R664 B.n677 B.n676 585
R665 B.n675 B.n674 585
R666 B.n673 B.n672 585
R667 B.n671 B.n670 585
R668 B.n669 B.n668 585
R669 B.n667 B.n666 585
R670 B.n665 B.n664 585
R671 B.n663 B.n662 585
R672 B.n660 B.n659 585
R673 B.n658 B.n657 585
R674 B.n656 B.n655 585
R675 B.n654 B.n653 585
R676 B.n652 B.n651 585
R677 B.n650 B.n649 585
R678 B.n648 B.n647 585
R679 B.n646 B.n645 585
R680 B.n644 B.n643 585
R681 B.n642 B.n641 585
R682 B.n640 B.n639 585
R683 B.n638 B.n637 585
R684 B.n636 B.n635 585
R685 B.n634 B.n633 585
R686 B.n632 B.n631 585
R687 B.n630 B.n629 585
R688 B.n628 B.n627 585
R689 B.n626 B.n625 585
R690 B.n624 B.n623 585
R691 B.n622 B.n621 585
R692 B.n620 B.n619 585
R693 B.n618 B.n617 585
R694 B.n616 B.n615 585
R695 B.n614 B.n613 585
R696 B.n612 B.n611 585
R697 B.n610 B.n609 585
R698 B.n608 B.n607 585
R699 B.n606 B.n605 585
R700 B.n604 B.n603 585
R701 B.n602 B.n601 585
R702 B.n600 B.n599 585
R703 B.n598 B.n597 585
R704 B.n596 B.n595 585
R705 B.n594 B.n593 585
R706 B.n592 B.n591 585
R707 B.n590 B.n589 585
R708 B.n588 B.n587 585
R709 B.n586 B.n585 585
R710 B.n584 B.n583 585
R711 B.n582 B.n581 585
R712 B.n580 B.n579 585
R713 B.n578 B.n577 585
R714 B.n576 B.n575 585
R715 B.n574 B.n573 585
R716 B.n572 B.n571 585
R717 B.n769 B.n514 585
R718 B.n514 B.n513 585
R719 B.n771 B.n770 585
R720 B.n772 B.n771 585
R721 B.n508 B.n507 585
R722 B.n509 B.n508 585
R723 B.n780 B.n779 585
R724 B.n779 B.n778 585
R725 B.n781 B.n506 585
R726 B.n506 B.n505 585
R727 B.n783 B.n782 585
R728 B.n784 B.n783 585
R729 B.n500 B.n499 585
R730 B.n501 B.n500 585
R731 B.n793 B.n792 585
R732 B.n792 B.n791 585
R733 B.n794 B.n498 585
R734 B.n790 B.n498 585
R735 B.n796 B.n795 585
R736 B.n797 B.n796 585
R737 B.n493 B.n492 585
R738 B.n494 B.n493 585
R739 B.n805 B.n804 585
R740 B.n804 B.n803 585
R741 B.n806 B.n491 585
R742 B.n491 B.n490 585
R743 B.n808 B.n807 585
R744 B.n809 B.n808 585
R745 B.n485 B.n484 585
R746 B.n486 B.n485 585
R747 B.n817 B.n816 585
R748 B.n816 B.n815 585
R749 B.n818 B.n483 585
R750 B.n483 B.n482 585
R751 B.n820 B.n819 585
R752 B.n821 B.n820 585
R753 B.n477 B.n476 585
R754 B.n478 B.n477 585
R755 B.n829 B.n828 585
R756 B.n828 B.n827 585
R757 B.n830 B.n475 585
R758 B.n475 B.n473 585
R759 B.n832 B.n831 585
R760 B.n833 B.n832 585
R761 B.n469 B.n468 585
R762 B.n474 B.n469 585
R763 B.n841 B.n840 585
R764 B.n840 B.n839 585
R765 B.n842 B.n467 585
R766 B.n467 B.n466 585
R767 B.n844 B.n843 585
R768 B.n845 B.n844 585
R769 B.n461 B.n460 585
R770 B.n462 B.n461 585
R771 B.n853 B.n852 585
R772 B.n852 B.n851 585
R773 B.n854 B.n459 585
R774 B.n459 B.n458 585
R775 B.n856 B.n855 585
R776 B.n857 B.n856 585
R777 B.n453 B.n452 585
R778 B.n454 B.n453 585
R779 B.n866 B.n865 585
R780 B.n865 B.n864 585
R781 B.n867 B.n451 585
R782 B.n863 B.n451 585
R783 B.n869 B.n868 585
R784 B.n870 B.n869 585
R785 B.n446 B.n445 585
R786 B.n447 B.n446 585
R787 B.n878 B.n877 585
R788 B.n877 B.n876 585
R789 B.n879 B.n444 585
R790 B.n444 B.n443 585
R791 B.n881 B.n880 585
R792 B.n882 B.n881 585
R793 B.n438 B.n437 585
R794 B.n439 B.n438 585
R795 B.n890 B.n889 585
R796 B.n889 B.n888 585
R797 B.n891 B.n436 585
R798 B.n436 B.n435 585
R799 B.n893 B.n892 585
R800 B.n894 B.n893 585
R801 B.n430 B.n429 585
R802 B.n431 B.n430 585
R803 B.n902 B.n901 585
R804 B.n901 B.n900 585
R805 B.n903 B.n428 585
R806 B.n428 B.n427 585
R807 B.n905 B.n904 585
R808 B.n906 B.n905 585
R809 B.n422 B.n421 585
R810 B.n423 B.n422 585
R811 B.n914 B.n913 585
R812 B.n913 B.n912 585
R813 B.n915 B.n420 585
R814 B.n420 B.n419 585
R815 B.n917 B.n916 585
R816 B.n918 B.n917 585
R817 B.n414 B.n413 585
R818 B.n415 B.n414 585
R819 B.n926 B.n925 585
R820 B.n925 B.n924 585
R821 B.n927 B.n412 585
R822 B.n412 B.n411 585
R823 B.n929 B.n928 585
R824 B.n930 B.n929 585
R825 B.n406 B.n405 585
R826 B.n407 B.n406 585
R827 B.n938 B.n937 585
R828 B.n937 B.n936 585
R829 B.n939 B.n404 585
R830 B.n404 B.n403 585
R831 B.n941 B.n940 585
R832 B.n942 B.n941 585
R833 B.n398 B.n397 585
R834 B.n399 B.n398 585
R835 B.n950 B.n949 585
R836 B.n949 B.n948 585
R837 B.n951 B.n396 585
R838 B.n396 B.n395 585
R839 B.n953 B.n952 585
R840 B.n954 B.n953 585
R841 B.n390 B.n389 585
R842 B.n391 B.n390 585
R843 B.n963 B.n962 585
R844 B.n962 B.n961 585
R845 B.n964 B.n388 585
R846 B.n960 B.n388 585
R847 B.n966 B.n965 585
R848 B.n967 B.n966 585
R849 B.n383 B.n382 585
R850 B.n384 B.n383 585
R851 B.n976 B.n975 585
R852 B.n975 B.n974 585
R853 B.n977 B.n381 585
R854 B.n381 B.n380 585
R855 B.n979 B.n978 585
R856 B.n980 B.n979 585
R857 B.n2 B.n0 585
R858 B.n4 B.n2 585
R859 B.n3 B.n1 585
R860 B.n1219 B.n3 585
R861 B.n1217 B.n1216 585
R862 B.n1218 B.n1217 585
R863 B.n1215 B.n9 585
R864 B.n9 B.n8 585
R865 B.n1214 B.n1213 585
R866 B.n1213 B.n1212 585
R867 B.n11 B.n10 585
R868 B.n1211 B.n11 585
R869 B.n1209 B.n1208 585
R870 B.n1210 B.n1209 585
R871 B.n1207 B.n15 585
R872 B.n18 B.n15 585
R873 B.n1206 B.n1205 585
R874 B.n1205 B.n1204 585
R875 B.n17 B.n16 585
R876 B.n1203 B.n17 585
R877 B.n1201 B.n1200 585
R878 B.n1202 B.n1201 585
R879 B.n1199 B.n23 585
R880 B.n23 B.n22 585
R881 B.n1198 B.n1197 585
R882 B.n1197 B.n1196 585
R883 B.n25 B.n24 585
R884 B.n1195 B.n25 585
R885 B.n1193 B.n1192 585
R886 B.n1194 B.n1193 585
R887 B.n1191 B.n30 585
R888 B.n30 B.n29 585
R889 B.n1190 B.n1189 585
R890 B.n1189 B.n1188 585
R891 B.n32 B.n31 585
R892 B.n1187 B.n32 585
R893 B.n1185 B.n1184 585
R894 B.n1186 B.n1185 585
R895 B.n1183 B.n37 585
R896 B.n37 B.n36 585
R897 B.n1182 B.n1181 585
R898 B.n1181 B.n1180 585
R899 B.n39 B.n38 585
R900 B.n1179 B.n39 585
R901 B.n1177 B.n1176 585
R902 B.n1178 B.n1177 585
R903 B.n1175 B.n44 585
R904 B.n44 B.n43 585
R905 B.n1174 B.n1173 585
R906 B.n1173 B.n1172 585
R907 B.n46 B.n45 585
R908 B.n1171 B.n46 585
R909 B.n1169 B.n1168 585
R910 B.n1170 B.n1169 585
R911 B.n1167 B.n51 585
R912 B.n51 B.n50 585
R913 B.n1166 B.n1165 585
R914 B.n1165 B.n1164 585
R915 B.n53 B.n52 585
R916 B.n1163 B.n53 585
R917 B.n1161 B.n1160 585
R918 B.n1162 B.n1161 585
R919 B.n1159 B.n58 585
R920 B.n58 B.n57 585
R921 B.n1158 B.n1157 585
R922 B.n1157 B.n1156 585
R923 B.n60 B.n59 585
R924 B.n1155 B.n60 585
R925 B.n1153 B.n1152 585
R926 B.n1154 B.n1153 585
R927 B.n1151 B.n65 585
R928 B.n65 B.n64 585
R929 B.n1150 B.n1149 585
R930 B.n1149 B.n1148 585
R931 B.n67 B.n66 585
R932 B.n1147 B.n67 585
R933 B.n1145 B.n1144 585
R934 B.n1146 B.n1145 585
R935 B.n1143 B.n71 585
R936 B.n74 B.n71 585
R937 B.n1142 B.n1141 585
R938 B.n1141 B.n1140 585
R939 B.n73 B.n72 585
R940 B.n1139 B.n73 585
R941 B.n1137 B.n1136 585
R942 B.n1138 B.n1137 585
R943 B.n1135 B.n79 585
R944 B.n79 B.n78 585
R945 B.n1134 B.n1133 585
R946 B.n1133 B.n1132 585
R947 B.n81 B.n80 585
R948 B.n1131 B.n81 585
R949 B.n1129 B.n1128 585
R950 B.n1130 B.n1129 585
R951 B.n1127 B.n86 585
R952 B.n86 B.n85 585
R953 B.n1126 B.n1125 585
R954 B.n1125 B.n1124 585
R955 B.n88 B.n87 585
R956 B.n1123 B.n88 585
R957 B.n1121 B.n1120 585
R958 B.n1122 B.n1121 585
R959 B.n1119 B.n93 585
R960 B.n93 B.n92 585
R961 B.n1118 B.n1117 585
R962 B.n1117 B.n1116 585
R963 B.n95 B.n94 585
R964 B.n1115 B.n95 585
R965 B.n1113 B.n1112 585
R966 B.n1114 B.n1113 585
R967 B.n1111 B.n100 585
R968 B.n100 B.n99 585
R969 B.n1110 B.n1109 585
R970 B.n1109 B.n1108 585
R971 B.n102 B.n101 585
R972 B.n1107 B.n102 585
R973 B.n1105 B.n1104 585
R974 B.n1106 B.n1105 585
R975 B.n1103 B.n107 585
R976 B.n107 B.n106 585
R977 B.n1102 B.n1101 585
R978 B.n1101 B.n1100 585
R979 B.n109 B.n108 585
R980 B.n1099 B.n109 585
R981 B.n1097 B.n1096 585
R982 B.n1098 B.n1097 585
R983 B.n1095 B.n113 585
R984 B.n116 B.n113 585
R985 B.n1094 B.n1093 585
R986 B.n1093 B.n1092 585
R987 B.n115 B.n114 585
R988 B.n1091 B.n115 585
R989 B.n1089 B.n1088 585
R990 B.n1090 B.n1089 585
R991 B.n1087 B.n121 585
R992 B.n121 B.n120 585
R993 B.n1086 B.n1085 585
R994 B.n1085 B.n1084 585
R995 B.n123 B.n122 585
R996 B.n1083 B.n123 585
R997 B.n1081 B.n1080 585
R998 B.n1082 B.n1081 585
R999 B.n1079 B.n128 585
R1000 B.n128 B.n127 585
R1001 B.n1222 B.n1221 585
R1002 B.n1221 B.n1220 585
R1003 B.n767 B.n514 502.111
R1004 B.n1077 B.n128 502.111
R1005 B.n571 B.n512 502.111
R1006 B.n1074 B.n180 502.111
R1007 B.n569 B.t11 305.69
R1008 B.n566 B.t7 305.69
R1009 B.n184 B.t3 305.69
R1010 B.n181 B.t14 305.69
R1011 B.n1075 B.n178 256.663
R1012 B.n1075 B.n177 256.663
R1013 B.n1075 B.n176 256.663
R1014 B.n1075 B.n175 256.663
R1015 B.n1075 B.n174 256.663
R1016 B.n1075 B.n173 256.663
R1017 B.n1075 B.n172 256.663
R1018 B.n1075 B.n171 256.663
R1019 B.n1075 B.n170 256.663
R1020 B.n1075 B.n169 256.663
R1021 B.n1075 B.n168 256.663
R1022 B.n1075 B.n167 256.663
R1023 B.n1075 B.n166 256.663
R1024 B.n1075 B.n165 256.663
R1025 B.n1075 B.n164 256.663
R1026 B.n1075 B.n163 256.663
R1027 B.n1075 B.n162 256.663
R1028 B.n1075 B.n161 256.663
R1029 B.n1075 B.n160 256.663
R1030 B.n1075 B.n159 256.663
R1031 B.n1075 B.n158 256.663
R1032 B.n1075 B.n157 256.663
R1033 B.n1075 B.n156 256.663
R1034 B.n1075 B.n155 256.663
R1035 B.n1075 B.n154 256.663
R1036 B.n1075 B.n153 256.663
R1037 B.n1075 B.n152 256.663
R1038 B.n1075 B.n151 256.663
R1039 B.n1075 B.n150 256.663
R1040 B.n1075 B.n149 256.663
R1041 B.n1075 B.n148 256.663
R1042 B.n1075 B.n147 256.663
R1043 B.n1075 B.n146 256.663
R1044 B.n1075 B.n145 256.663
R1045 B.n1075 B.n144 256.663
R1046 B.n1075 B.n143 256.663
R1047 B.n1075 B.n142 256.663
R1048 B.n1075 B.n141 256.663
R1049 B.n1075 B.n140 256.663
R1050 B.n1075 B.n139 256.663
R1051 B.n1075 B.n138 256.663
R1052 B.n1075 B.n137 256.663
R1053 B.n1075 B.n136 256.663
R1054 B.n1075 B.n135 256.663
R1055 B.n1075 B.n134 256.663
R1056 B.n1075 B.n133 256.663
R1057 B.n1075 B.n132 256.663
R1058 B.n1075 B.n131 256.663
R1059 B.n1076 B.n1075 256.663
R1060 B.n766 B.n765 256.663
R1061 B.n765 B.n517 256.663
R1062 B.n765 B.n518 256.663
R1063 B.n765 B.n519 256.663
R1064 B.n765 B.n520 256.663
R1065 B.n765 B.n521 256.663
R1066 B.n765 B.n522 256.663
R1067 B.n765 B.n523 256.663
R1068 B.n765 B.n524 256.663
R1069 B.n765 B.n525 256.663
R1070 B.n765 B.n526 256.663
R1071 B.n765 B.n527 256.663
R1072 B.n765 B.n528 256.663
R1073 B.n765 B.n529 256.663
R1074 B.n765 B.n530 256.663
R1075 B.n765 B.n531 256.663
R1076 B.n765 B.n532 256.663
R1077 B.n765 B.n533 256.663
R1078 B.n765 B.n534 256.663
R1079 B.n765 B.n535 256.663
R1080 B.n765 B.n536 256.663
R1081 B.n765 B.n537 256.663
R1082 B.n765 B.n538 256.663
R1083 B.n765 B.n539 256.663
R1084 B.n765 B.n540 256.663
R1085 B.n765 B.n541 256.663
R1086 B.n765 B.n542 256.663
R1087 B.n765 B.n543 256.663
R1088 B.n765 B.n544 256.663
R1089 B.n765 B.n545 256.663
R1090 B.n765 B.n546 256.663
R1091 B.n765 B.n547 256.663
R1092 B.n765 B.n548 256.663
R1093 B.n765 B.n549 256.663
R1094 B.n765 B.n550 256.663
R1095 B.n765 B.n551 256.663
R1096 B.n765 B.n552 256.663
R1097 B.n765 B.n553 256.663
R1098 B.n765 B.n554 256.663
R1099 B.n765 B.n555 256.663
R1100 B.n765 B.n556 256.663
R1101 B.n765 B.n557 256.663
R1102 B.n765 B.n558 256.663
R1103 B.n765 B.n559 256.663
R1104 B.n765 B.n560 256.663
R1105 B.n765 B.n561 256.663
R1106 B.n765 B.n562 256.663
R1107 B.n765 B.n563 256.663
R1108 B.n765 B.n564 256.663
R1109 B.n771 B.n514 163.367
R1110 B.n771 B.n508 163.367
R1111 B.n779 B.n508 163.367
R1112 B.n779 B.n506 163.367
R1113 B.n783 B.n506 163.367
R1114 B.n783 B.n500 163.367
R1115 B.n792 B.n500 163.367
R1116 B.n792 B.n498 163.367
R1117 B.n796 B.n498 163.367
R1118 B.n796 B.n493 163.367
R1119 B.n804 B.n493 163.367
R1120 B.n804 B.n491 163.367
R1121 B.n808 B.n491 163.367
R1122 B.n808 B.n485 163.367
R1123 B.n816 B.n485 163.367
R1124 B.n816 B.n483 163.367
R1125 B.n820 B.n483 163.367
R1126 B.n820 B.n477 163.367
R1127 B.n828 B.n477 163.367
R1128 B.n828 B.n475 163.367
R1129 B.n832 B.n475 163.367
R1130 B.n832 B.n469 163.367
R1131 B.n840 B.n469 163.367
R1132 B.n840 B.n467 163.367
R1133 B.n844 B.n467 163.367
R1134 B.n844 B.n461 163.367
R1135 B.n852 B.n461 163.367
R1136 B.n852 B.n459 163.367
R1137 B.n856 B.n459 163.367
R1138 B.n856 B.n453 163.367
R1139 B.n865 B.n453 163.367
R1140 B.n865 B.n451 163.367
R1141 B.n869 B.n451 163.367
R1142 B.n869 B.n446 163.367
R1143 B.n877 B.n446 163.367
R1144 B.n877 B.n444 163.367
R1145 B.n881 B.n444 163.367
R1146 B.n881 B.n438 163.367
R1147 B.n889 B.n438 163.367
R1148 B.n889 B.n436 163.367
R1149 B.n893 B.n436 163.367
R1150 B.n893 B.n430 163.367
R1151 B.n901 B.n430 163.367
R1152 B.n901 B.n428 163.367
R1153 B.n905 B.n428 163.367
R1154 B.n905 B.n422 163.367
R1155 B.n913 B.n422 163.367
R1156 B.n913 B.n420 163.367
R1157 B.n917 B.n420 163.367
R1158 B.n917 B.n414 163.367
R1159 B.n925 B.n414 163.367
R1160 B.n925 B.n412 163.367
R1161 B.n929 B.n412 163.367
R1162 B.n929 B.n406 163.367
R1163 B.n937 B.n406 163.367
R1164 B.n937 B.n404 163.367
R1165 B.n941 B.n404 163.367
R1166 B.n941 B.n398 163.367
R1167 B.n949 B.n398 163.367
R1168 B.n949 B.n396 163.367
R1169 B.n953 B.n396 163.367
R1170 B.n953 B.n390 163.367
R1171 B.n962 B.n390 163.367
R1172 B.n962 B.n388 163.367
R1173 B.n966 B.n388 163.367
R1174 B.n966 B.n383 163.367
R1175 B.n975 B.n383 163.367
R1176 B.n975 B.n381 163.367
R1177 B.n979 B.n381 163.367
R1178 B.n979 B.n2 163.367
R1179 B.n1221 B.n2 163.367
R1180 B.n1221 B.n3 163.367
R1181 B.n1217 B.n3 163.367
R1182 B.n1217 B.n9 163.367
R1183 B.n1213 B.n9 163.367
R1184 B.n1213 B.n11 163.367
R1185 B.n1209 B.n11 163.367
R1186 B.n1209 B.n15 163.367
R1187 B.n1205 B.n15 163.367
R1188 B.n1205 B.n17 163.367
R1189 B.n1201 B.n17 163.367
R1190 B.n1201 B.n23 163.367
R1191 B.n1197 B.n23 163.367
R1192 B.n1197 B.n25 163.367
R1193 B.n1193 B.n25 163.367
R1194 B.n1193 B.n30 163.367
R1195 B.n1189 B.n30 163.367
R1196 B.n1189 B.n32 163.367
R1197 B.n1185 B.n32 163.367
R1198 B.n1185 B.n37 163.367
R1199 B.n1181 B.n37 163.367
R1200 B.n1181 B.n39 163.367
R1201 B.n1177 B.n39 163.367
R1202 B.n1177 B.n44 163.367
R1203 B.n1173 B.n44 163.367
R1204 B.n1173 B.n46 163.367
R1205 B.n1169 B.n46 163.367
R1206 B.n1169 B.n51 163.367
R1207 B.n1165 B.n51 163.367
R1208 B.n1165 B.n53 163.367
R1209 B.n1161 B.n53 163.367
R1210 B.n1161 B.n58 163.367
R1211 B.n1157 B.n58 163.367
R1212 B.n1157 B.n60 163.367
R1213 B.n1153 B.n60 163.367
R1214 B.n1153 B.n65 163.367
R1215 B.n1149 B.n65 163.367
R1216 B.n1149 B.n67 163.367
R1217 B.n1145 B.n67 163.367
R1218 B.n1145 B.n71 163.367
R1219 B.n1141 B.n71 163.367
R1220 B.n1141 B.n73 163.367
R1221 B.n1137 B.n73 163.367
R1222 B.n1137 B.n79 163.367
R1223 B.n1133 B.n79 163.367
R1224 B.n1133 B.n81 163.367
R1225 B.n1129 B.n81 163.367
R1226 B.n1129 B.n86 163.367
R1227 B.n1125 B.n86 163.367
R1228 B.n1125 B.n88 163.367
R1229 B.n1121 B.n88 163.367
R1230 B.n1121 B.n93 163.367
R1231 B.n1117 B.n93 163.367
R1232 B.n1117 B.n95 163.367
R1233 B.n1113 B.n95 163.367
R1234 B.n1113 B.n100 163.367
R1235 B.n1109 B.n100 163.367
R1236 B.n1109 B.n102 163.367
R1237 B.n1105 B.n102 163.367
R1238 B.n1105 B.n107 163.367
R1239 B.n1101 B.n107 163.367
R1240 B.n1101 B.n109 163.367
R1241 B.n1097 B.n109 163.367
R1242 B.n1097 B.n113 163.367
R1243 B.n1093 B.n113 163.367
R1244 B.n1093 B.n115 163.367
R1245 B.n1089 B.n115 163.367
R1246 B.n1089 B.n121 163.367
R1247 B.n1085 B.n121 163.367
R1248 B.n1085 B.n123 163.367
R1249 B.n1081 B.n123 163.367
R1250 B.n1081 B.n128 163.367
R1251 B.n764 B.n516 163.367
R1252 B.n764 B.n565 163.367
R1253 B.n760 B.n759 163.367
R1254 B.n756 B.n755 163.367
R1255 B.n752 B.n751 163.367
R1256 B.n748 B.n747 163.367
R1257 B.n744 B.n743 163.367
R1258 B.n740 B.n739 163.367
R1259 B.n736 B.n735 163.367
R1260 B.n732 B.n731 163.367
R1261 B.n728 B.n727 163.367
R1262 B.n724 B.n723 163.367
R1263 B.n720 B.n719 163.367
R1264 B.n716 B.n715 163.367
R1265 B.n712 B.n711 163.367
R1266 B.n708 B.n707 163.367
R1267 B.n704 B.n703 163.367
R1268 B.n700 B.n699 163.367
R1269 B.n696 B.n695 163.367
R1270 B.n692 B.n691 163.367
R1271 B.n688 B.n687 163.367
R1272 B.n684 B.n683 163.367
R1273 B.n680 B.n679 163.367
R1274 B.n676 B.n675 163.367
R1275 B.n672 B.n671 163.367
R1276 B.n668 B.n667 163.367
R1277 B.n664 B.n663 163.367
R1278 B.n659 B.n658 163.367
R1279 B.n655 B.n654 163.367
R1280 B.n651 B.n650 163.367
R1281 B.n647 B.n646 163.367
R1282 B.n643 B.n642 163.367
R1283 B.n639 B.n638 163.367
R1284 B.n635 B.n634 163.367
R1285 B.n631 B.n630 163.367
R1286 B.n627 B.n626 163.367
R1287 B.n623 B.n622 163.367
R1288 B.n619 B.n618 163.367
R1289 B.n615 B.n614 163.367
R1290 B.n611 B.n610 163.367
R1291 B.n607 B.n606 163.367
R1292 B.n603 B.n602 163.367
R1293 B.n599 B.n598 163.367
R1294 B.n595 B.n594 163.367
R1295 B.n591 B.n590 163.367
R1296 B.n587 B.n586 163.367
R1297 B.n583 B.n582 163.367
R1298 B.n579 B.n578 163.367
R1299 B.n575 B.n574 163.367
R1300 B.n773 B.n512 163.367
R1301 B.n773 B.n510 163.367
R1302 B.n777 B.n510 163.367
R1303 B.n777 B.n504 163.367
R1304 B.n785 B.n504 163.367
R1305 B.n785 B.n502 163.367
R1306 B.n789 B.n502 163.367
R1307 B.n789 B.n497 163.367
R1308 B.n798 B.n497 163.367
R1309 B.n798 B.n495 163.367
R1310 B.n802 B.n495 163.367
R1311 B.n802 B.n489 163.367
R1312 B.n810 B.n489 163.367
R1313 B.n810 B.n487 163.367
R1314 B.n814 B.n487 163.367
R1315 B.n814 B.n481 163.367
R1316 B.n822 B.n481 163.367
R1317 B.n822 B.n479 163.367
R1318 B.n826 B.n479 163.367
R1319 B.n826 B.n472 163.367
R1320 B.n834 B.n472 163.367
R1321 B.n834 B.n470 163.367
R1322 B.n838 B.n470 163.367
R1323 B.n838 B.n465 163.367
R1324 B.n846 B.n465 163.367
R1325 B.n846 B.n463 163.367
R1326 B.n850 B.n463 163.367
R1327 B.n850 B.n457 163.367
R1328 B.n858 B.n457 163.367
R1329 B.n858 B.n455 163.367
R1330 B.n862 B.n455 163.367
R1331 B.n862 B.n450 163.367
R1332 B.n871 B.n450 163.367
R1333 B.n871 B.n448 163.367
R1334 B.n875 B.n448 163.367
R1335 B.n875 B.n442 163.367
R1336 B.n883 B.n442 163.367
R1337 B.n883 B.n440 163.367
R1338 B.n887 B.n440 163.367
R1339 B.n887 B.n434 163.367
R1340 B.n895 B.n434 163.367
R1341 B.n895 B.n432 163.367
R1342 B.n899 B.n432 163.367
R1343 B.n899 B.n426 163.367
R1344 B.n907 B.n426 163.367
R1345 B.n907 B.n424 163.367
R1346 B.n911 B.n424 163.367
R1347 B.n911 B.n418 163.367
R1348 B.n919 B.n418 163.367
R1349 B.n919 B.n416 163.367
R1350 B.n923 B.n416 163.367
R1351 B.n923 B.n410 163.367
R1352 B.n931 B.n410 163.367
R1353 B.n931 B.n408 163.367
R1354 B.n935 B.n408 163.367
R1355 B.n935 B.n402 163.367
R1356 B.n943 B.n402 163.367
R1357 B.n943 B.n400 163.367
R1358 B.n947 B.n400 163.367
R1359 B.n947 B.n394 163.367
R1360 B.n955 B.n394 163.367
R1361 B.n955 B.n392 163.367
R1362 B.n959 B.n392 163.367
R1363 B.n959 B.n387 163.367
R1364 B.n968 B.n387 163.367
R1365 B.n968 B.n385 163.367
R1366 B.n973 B.n385 163.367
R1367 B.n973 B.n379 163.367
R1368 B.n981 B.n379 163.367
R1369 B.n982 B.n981 163.367
R1370 B.n982 B.n5 163.367
R1371 B.n6 B.n5 163.367
R1372 B.n7 B.n6 163.367
R1373 B.n987 B.n7 163.367
R1374 B.n987 B.n12 163.367
R1375 B.n13 B.n12 163.367
R1376 B.n14 B.n13 163.367
R1377 B.n992 B.n14 163.367
R1378 B.n992 B.n19 163.367
R1379 B.n20 B.n19 163.367
R1380 B.n21 B.n20 163.367
R1381 B.n997 B.n21 163.367
R1382 B.n997 B.n26 163.367
R1383 B.n27 B.n26 163.367
R1384 B.n28 B.n27 163.367
R1385 B.n1002 B.n28 163.367
R1386 B.n1002 B.n33 163.367
R1387 B.n34 B.n33 163.367
R1388 B.n35 B.n34 163.367
R1389 B.n1007 B.n35 163.367
R1390 B.n1007 B.n40 163.367
R1391 B.n41 B.n40 163.367
R1392 B.n42 B.n41 163.367
R1393 B.n1012 B.n42 163.367
R1394 B.n1012 B.n47 163.367
R1395 B.n48 B.n47 163.367
R1396 B.n49 B.n48 163.367
R1397 B.n1017 B.n49 163.367
R1398 B.n1017 B.n54 163.367
R1399 B.n55 B.n54 163.367
R1400 B.n56 B.n55 163.367
R1401 B.n1022 B.n56 163.367
R1402 B.n1022 B.n61 163.367
R1403 B.n62 B.n61 163.367
R1404 B.n63 B.n62 163.367
R1405 B.n1027 B.n63 163.367
R1406 B.n1027 B.n68 163.367
R1407 B.n69 B.n68 163.367
R1408 B.n70 B.n69 163.367
R1409 B.n1032 B.n70 163.367
R1410 B.n1032 B.n75 163.367
R1411 B.n76 B.n75 163.367
R1412 B.n77 B.n76 163.367
R1413 B.n1037 B.n77 163.367
R1414 B.n1037 B.n82 163.367
R1415 B.n83 B.n82 163.367
R1416 B.n84 B.n83 163.367
R1417 B.n1042 B.n84 163.367
R1418 B.n1042 B.n89 163.367
R1419 B.n90 B.n89 163.367
R1420 B.n91 B.n90 163.367
R1421 B.n1047 B.n91 163.367
R1422 B.n1047 B.n96 163.367
R1423 B.n97 B.n96 163.367
R1424 B.n98 B.n97 163.367
R1425 B.n1052 B.n98 163.367
R1426 B.n1052 B.n103 163.367
R1427 B.n104 B.n103 163.367
R1428 B.n105 B.n104 163.367
R1429 B.n1057 B.n105 163.367
R1430 B.n1057 B.n110 163.367
R1431 B.n111 B.n110 163.367
R1432 B.n112 B.n111 163.367
R1433 B.n1062 B.n112 163.367
R1434 B.n1062 B.n117 163.367
R1435 B.n118 B.n117 163.367
R1436 B.n119 B.n118 163.367
R1437 B.n1067 B.n119 163.367
R1438 B.n1067 B.n124 163.367
R1439 B.n125 B.n124 163.367
R1440 B.n126 B.n125 163.367
R1441 B.n180 B.n126 163.367
R1442 B.n186 B.n130 163.367
R1443 B.n190 B.n189 163.367
R1444 B.n194 B.n193 163.367
R1445 B.n198 B.n197 163.367
R1446 B.n202 B.n201 163.367
R1447 B.n206 B.n205 163.367
R1448 B.n210 B.n209 163.367
R1449 B.n214 B.n213 163.367
R1450 B.n218 B.n217 163.367
R1451 B.n222 B.n221 163.367
R1452 B.n226 B.n225 163.367
R1453 B.n230 B.n229 163.367
R1454 B.n234 B.n233 163.367
R1455 B.n238 B.n237 163.367
R1456 B.n242 B.n241 163.367
R1457 B.n246 B.n245 163.367
R1458 B.n250 B.n249 163.367
R1459 B.n254 B.n253 163.367
R1460 B.n258 B.n257 163.367
R1461 B.n262 B.n261 163.367
R1462 B.n266 B.n265 163.367
R1463 B.n270 B.n269 163.367
R1464 B.n275 B.n274 163.367
R1465 B.n279 B.n278 163.367
R1466 B.n283 B.n282 163.367
R1467 B.n287 B.n286 163.367
R1468 B.n291 B.n290 163.367
R1469 B.n295 B.n294 163.367
R1470 B.n299 B.n298 163.367
R1471 B.n303 B.n302 163.367
R1472 B.n307 B.n306 163.367
R1473 B.n311 B.n310 163.367
R1474 B.n315 B.n314 163.367
R1475 B.n319 B.n318 163.367
R1476 B.n323 B.n322 163.367
R1477 B.n327 B.n326 163.367
R1478 B.n331 B.n330 163.367
R1479 B.n335 B.n334 163.367
R1480 B.n339 B.n338 163.367
R1481 B.n343 B.n342 163.367
R1482 B.n347 B.n346 163.367
R1483 B.n351 B.n350 163.367
R1484 B.n355 B.n354 163.367
R1485 B.n359 B.n358 163.367
R1486 B.n363 B.n362 163.367
R1487 B.n367 B.n366 163.367
R1488 B.n371 B.n370 163.367
R1489 B.n375 B.n374 163.367
R1490 B.n1074 B.n179 163.367
R1491 B.n569 B.t13 138.838
R1492 B.n181 B.t15 138.838
R1493 B.n566 B.t10 138.821
R1494 B.n184 B.t5 138.821
R1495 B.n765 B.n513 78.7652
R1496 B.n1075 B.n127 78.7652
R1497 B.n767 B.n766 71.676
R1498 B.n565 B.n517 71.676
R1499 B.n759 B.n518 71.676
R1500 B.n755 B.n519 71.676
R1501 B.n751 B.n520 71.676
R1502 B.n747 B.n521 71.676
R1503 B.n743 B.n522 71.676
R1504 B.n739 B.n523 71.676
R1505 B.n735 B.n524 71.676
R1506 B.n731 B.n525 71.676
R1507 B.n727 B.n526 71.676
R1508 B.n723 B.n527 71.676
R1509 B.n719 B.n528 71.676
R1510 B.n715 B.n529 71.676
R1511 B.n711 B.n530 71.676
R1512 B.n707 B.n531 71.676
R1513 B.n703 B.n532 71.676
R1514 B.n699 B.n533 71.676
R1515 B.n695 B.n534 71.676
R1516 B.n691 B.n535 71.676
R1517 B.n687 B.n536 71.676
R1518 B.n683 B.n537 71.676
R1519 B.n679 B.n538 71.676
R1520 B.n675 B.n539 71.676
R1521 B.n671 B.n540 71.676
R1522 B.n667 B.n541 71.676
R1523 B.n663 B.n542 71.676
R1524 B.n658 B.n543 71.676
R1525 B.n654 B.n544 71.676
R1526 B.n650 B.n545 71.676
R1527 B.n646 B.n546 71.676
R1528 B.n642 B.n547 71.676
R1529 B.n638 B.n548 71.676
R1530 B.n634 B.n549 71.676
R1531 B.n630 B.n550 71.676
R1532 B.n626 B.n551 71.676
R1533 B.n622 B.n552 71.676
R1534 B.n618 B.n553 71.676
R1535 B.n614 B.n554 71.676
R1536 B.n610 B.n555 71.676
R1537 B.n606 B.n556 71.676
R1538 B.n602 B.n557 71.676
R1539 B.n598 B.n558 71.676
R1540 B.n594 B.n559 71.676
R1541 B.n590 B.n560 71.676
R1542 B.n586 B.n561 71.676
R1543 B.n582 B.n562 71.676
R1544 B.n578 B.n563 71.676
R1545 B.n574 B.n564 71.676
R1546 B.n1077 B.n1076 71.676
R1547 B.n186 B.n131 71.676
R1548 B.n190 B.n132 71.676
R1549 B.n194 B.n133 71.676
R1550 B.n198 B.n134 71.676
R1551 B.n202 B.n135 71.676
R1552 B.n206 B.n136 71.676
R1553 B.n210 B.n137 71.676
R1554 B.n214 B.n138 71.676
R1555 B.n218 B.n139 71.676
R1556 B.n222 B.n140 71.676
R1557 B.n226 B.n141 71.676
R1558 B.n230 B.n142 71.676
R1559 B.n234 B.n143 71.676
R1560 B.n238 B.n144 71.676
R1561 B.n242 B.n145 71.676
R1562 B.n246 B.n146 71.676
R1563 B.n250 B.n147 71.676
R1564 B.n254 B.n148 71.676
R1565 B.n258 B.n149 71.676
R1566 B.n262 B.n150 71.676
R1567 B.n266 B.n151 71.676
R1568 B.n270 B.n152 71.676
R1569 B.n275 B.n153 71.676
R1570 B.n279 B.n154 71.676
R1571 B.n283 B.n155 71.676
R1572 B.n287 B.n156 71.676
R1573 B.n291 B.n157 71.676
R1574 B.n295 B.n158 71.676
R1575 B.n299 B.n159 71.676
R1576 B.n303 B.n160 71.676
R1577 B.n307 B.n161 71.676
R1578 B.n311 B.n162 71.676
R1579 B.n315 B.n163 71.676
R1580 B.n319 B.n164 71.676
R1581 B.n323 B.n165 71.676
R1582 B.n327 B.n166 71.676
R1583 B.n331 B.n167 71.676
R1584 B.n335 B.n168 71.676
R1585 B.n339 B.n169 71.676
R1586 B.n343 B.n170 71.676
R1587 B.n347 B.n171 71.676
R1588 B.n351 B.n172 71.676
R1589 B.n355 B.n173 71.676
R1590 B.n359 B.n174 71.676
R1591 B.n363 B.n175 71.676
R1592 B.n367 B.n176 71.676
R1593 B.n371 B.n177 71.676
R1594 B.n375 B.n178 71.676
R1595 B.n179 B.n178 71.676
R1596 B.n374 B.n177 71.676
R1597 B.n370 B.n176 71.676
R1598 B.n366 B.n175 71.676
R1599 B.n362 B.n174 71.676
R1600 B.n358 B.n173 71.676
R1601 B.n354 B.n172 71.676
R1602 B.n350 B.n171 71.676
R1603 B.n346 B.n170 71.676
R1604 B.n342 B.n169 71.676
R1605 B.n338 B.n168 71.676
R1606 B.n334 B.n167 71.676
R1607 B.n330 B.n166 71.676
R1608 B.n326 B.n165 71.676
R1609 B.n322 B.n164 71.676
R1610 B.n318 B.n163 71.676
R1611 B.n314 B.n162 71.676
R1612 B.n310 B.n161 71.676
R1613 B.n306 B.n160 71.676
R1614 B.n302 B.n159 71.676
R1615 B.n298 B.n158 71.676
R1616 B.n294 B.n157 71.676
R1617 B.n290 B.n156 71.676
R1618 B.n286 B.n155 71.676
R1619 B.n282 B.n154 71.676
R1620 B.n278 B.n153 71.676
R1621 B.n274 B.n152 71.676
R1622 B.n269 B.n151 71.676
R1623 B.n265 B.n150 71.676
R1624 B.n261 B.n149 71.676
R1625 B.n257 B.n148 71.676
R1626 B.n253 B.n147 71.676
R1627 B.n249 B.n146 71.676
R1628 B.n245 B.n145 71.676
R1629 B.n241 B.n144 71.676
R1630 B.n237 B.n143 71.676
R1631 B.n233 B.n142 71.676
R1632 B.n229 B.n141 71.676
R1633 B.n225 B.n140 71.676
R1634 B.n221 B.n139 71.676
R1635 B.n217 B.n138 71.676
R1636 B.n213 B.n137 71.676
R1637 B.n209 B.n136 71.676
R1638 B.n205 B.n135 71.676
R1639 B.n201 B.n134 71.676
R1640 B.n197 B.n133 71.676
R1641 B.n193 B.n132 71.676
R1642 B.n189 B.n131 71.676
R1643 B.n1076 B.n130 71.676
R1644 B.n766 B.n516 71.676
R1645 B.n760 B.n517 71.676
R1646 B.n756 B.n518 71.676
R1647 B.n752 B.n519 71.676
R1648 B.n748 B.n520 71.676
R1649 B.n744 B.n521 71.676
R1650 B.n740 B.n522 71.676
R1651 B.n736 B.n523 71.676
R1652 B.n732 B.n524 71.676
R1653 B.n728 B.n525 71.676
R1654 B.n724 B.n526 71.676
R1655 B.n720 B.n527 71.676
R1656 B.n716 B.n528 71.676
R1657 B.n712 B.n529 71.676
R1658 B.n708 B.n530 71.676
R1659 B.n704 B.n531 71.676
R1660 B.n700 B.n532 71.676
R1661 B.n696 B.n533 71.676
R1662 B.n692 B.n534 71.676
R1663 B.n688 B.n535 71.676
R1664 B.n684 B.n536 71.676
R1665 B.n680 B.n537 71.676
R1666 B.n676 B.n538 71.676
R1667 B.n672 B.n539 71.676
R1668 B.n668 B.n540 71.676
R1669 B.n664 B.n541 71.676
R1670 B.n659 B.n542 71.676
R1671 B.n655 B.n543 71.676
R1672 B.n651 B.n544 71.676
R1673 B.n647 B.n545 71.676
R1674 B.n643 B.n546 71.676
R1675 B.n639 B.n547 71.676
R1676 B.n635 B.n548 71.676
R1677 B.n631 B.n549 71.676
R1678 B.n627 B.n550 71.676
R1679 B.n623 B.n551 71.676
R1680 B.n619 B.n552 71.676
R1681 B.n615 B.n553 71.676
R1682 B.n611 B.n554 71.676
R1683 B.n607 B.n555 71.676
R1684 B.n603 B.n556 71.676
R1685 B.n599 B.n557 71.676
R1686 B.n595 B.n558 71.676
R1687 B.n591 B.n559 71.676
R1688 B.n587 B.n560 71.676
R1689 B.n583 B.n561 71.676
R1690 B.n579 B.n562 71.676
R1691 B.n575 B.n563 71.676
R1692 B.n571 B.n564 71.676
R1693 B.n570 B.t12 69.6015
R1694 B.n182 B.t16 69.6015
R1695 B.n567 B.t9 69.5848
R1696 B.n185 B.t6 69.5848
R1697 B.n570 B.n569 69.2369
R1698 B.n567 B.n566 69.2369
R1699 B.n185 B.n184 69.2369
R1700 B.n182 B.n181 69.2369
R1701 B.n661 B.n570 59.5399
R1702 B.n568 B.n567 59.5399
R1703 B.n272 B.n185 59.5399
R1704 B.n183 B.n182 59.5399
R1705 B.n772 B.n513 40.886
R1706 B.n772 B.n509 40.886
R1707 B.n778 B.n509 40.886
R1708 B.n778 B.n505 40.886
R1709 B.n784 B.n505 40.886
R1710 B.n784 B.n501 40.886
R1711 B.n791 B.n501 40.886
R1712 B.n791 B.n790 40.886
R1713 B.n797 B.n494 40.886
R1714 B.n803 B.n494 40.886
R1715 B.n803 B.n490 40.886
R1716 B.n809 B.n490 40.886
R1717 B.n809 B.n486 40.886
R1718 B.n815 B.n486 40.886
R1719 B.n815 B.n482 40.886
R1720 B.n821 B.n482 40.886
R1721 B.n821 B.n478 40.886
R1722 B.n827 B.n478 40.886
R1723 B.n827 B.n473 40.886
R1724 B.n833 B.n473 40.886
R1725 B.n833 B.n474 40.886
R1726 B.n839 B.n466 40.886
R1727 B.n845 B.n466 40.886
R1728 B.n845 B.n462 40.886
R1729 B.n851 B.n462 40.886
R1730 B.n851 B.n458 40.886
R1731 B.n857 B.n458 40.886
R1732 B.n857 B.n454 40.886
R1733 B.n864 B.n454 40.886
R1734 B.n864 B.n863 40.886
R1735 B.n870 B.n447 40.886
R1736 B.n876 B.n447 40.886
R1737 B.n876 B.n443 40.886
R1738 B.n882 B.n443 40.886
R1739 B.n882 B.n439 40.886
R1740 B.n888 B.n439 40.886
R1741 B.n888 B.n435 40.886
R1742 B.n894 B.n435 40.886
R1743 B.n894 B.n431 40.886
R1744 B.n900 B.n431 40.886
R1745 B.n906 B.n427 40.886
R1746 B.n906 B.n423 40.886
R1747 B.n912 B.n423 40.886
R1748 B.n912 B.n419 40.886
R1749 B.n918 B.n419 40.886
R1750 B.n918 B.n415 40.886
R1751 B.n924 B.n415 40.886
R1752 B.n924 B.n411 40.886
R1753 B.n930 B.n411 40.886
R1754 B.n936 B.n407 40.886
R1755 B.n936 B.n403 40.886
R1756 B.n942 B.n403 40.886
R1757 B.n942 B.n399 40.886
R1758 B.n948 B.n399 40.886
R1759 B.n948 B.n395 40.886
R1760 B.n954 B.n395 40.886
R1761 B.n954 B.n391 40.886
R1762 B.n961 B.n391 40.886
R1763 B.n961 B.n960 40.886
R1764 B.n967 B.n384 40.886
R1765 B.n974 B.n384 40.886
R1766 B.n974 B.n380 40.886
R1767 B.n980 B.n380 40.886
R1768 B.n980 B.n4 40.886
R1769 B.n1220 B.n4 40.886
R1770 B.n1220 B.n1219 40.886
R1771 B.n1219 B.n1218 40.886
R1772 B.n1218 B.n8 40.886
R1773 B.n1212 B.n8 40.886
R1774 B.n1212 B.n1211 40.886
R1775 B.n1211 B.n1210 40.886
R1776 B.n1204 B.n18 40.886
R1777 B.n1204 B.n1203 40.886
R1778 B.n1203 B.n1202 40.886
R1779 B.n1202 B.n22 40.886
R1780 B.n1196 B.n22 40.886
R1781 B.n1196 B.n1195 40.886
R1782 B.n1195 B.n1194 40.886
R1783 B.n1194 B.n29 40.886
R1784 B.n1188 B.n29 40.886
R1785 B.n1188 B.n1187 40.886
R1786 B.n1186 B.n36 40.886
R1787 B.n1180 B.n36 40.886
R1788 B.n1180 B.n1179 40.886
R1789 B.n1179 B.n1178 40.886
R1790 B.n1178 B.n43 40.886
R1791 B.n1172 B.n43 40.886
R1792 B.n1172 B.n1171 40.886
R1793 B.n1171 B.n1170 40.886
R1794 B.n1170 B.n50 40.886
R1795 B.n1164 B.n1163 40.886
R1796 B.n1163 B.n1162 40.886
R1797 B.n1162 B.n57 40.886
R1798 B.n1156 B.n57 40.886
R1799 B.n1156 B.n1155 40.886
R1800 B.n1155 B.n1154 40.886
R1801 B.n1154 B.n64 40.886
R1802 B.n1148 B.n64 40.886
R1803 B.n1148 B.n1147 40.886
R1804 B.n1147 B.n1146 40.886
R1805 B.n1140 B.n74 40.886
R1806 B.n1140 B.n1139 40.886
R1807 B.n1139 B.n1138 40.886
R1808 B.n1138 B.n78 40.886
R1809 B.n1132 B.n78 40.886
R1810 B.n1132 B.n1131 40.886
R1811 B.n1131 B.n1130 40.886
R1812 B.n1130 B.n85 40.886
R1813 B.n1124 B.n85 40.886
R1814 B.n1123 B.n1122 40.886
R1815 B.n1122 B.n92 40.886
R1816 B.n1116 B.n92 40.886
R1817 B.n1116 B.n1115 40.886
R1818 B.n1115 B.n1114 40.886
R1819 B.n1114 B.n99 40.886
R1820 B.n1108 B.n99 40.886
R1821 B.n1108 B.n1107 40.886
R1822 B.n1107 B.n1106 40.886
R1823 B.n1106 B.n106 40.886
R1824 B.n1100 B.n106 40.886
R1825 B.n1100 B.n1099 40.886
R1826 B.n1099 B.n1098 40.886
R1827 B.n1092 B.n116 40.886
R1828 B.n1092 B.n1091 40.886
R1829 B.n1091 B.n1090 40.886
R1830 B.n1090 B.n120 40.886
R1831 B.n1084 B.n120 40.886
R1832 B.n1084 B.n1083 40.886
R1833 B.n1083 B.n1082 40.886
R1834 B.n1082 B.n127 40.886
R1835 B.n839 B.t0 34.8734
R1836 B.t23 B.n427 34.8734
R1837 B.n967 B.t19 34.8734
R1838 B.n1210 B.t22 34.8734
R1839 B.t18 B.n50 34.8734
R1840 B.n1124 B.t2 34.8734
R1841 B.n1079 B.n1078 32.6249
R1842 B.n1073 B.n1072 32.6249
R1843 B.n572 B.n511 32.6249
R1844 B.n769 B.n768 32.6249
R1845 B.n863 B.t17 26.4558
R1846 B.n930 B.t20 26.4558
R1847 B.t21 B.n1186 26.4558
R1848 B.n74 B.t1 26.4558
R1849 B.n797 B.t8 22.8483
R1850 B.n1098 B.t4 22.8483
R1851 B B.n1222 18.0485
R1852 B.n790 B.t8 18.0382
R1853 B.n116 B.t4 18.0382
R1854 B.n870 B.t17 14.4307
R1855 B.t20 B.n407 14.4307
R1856 B.n1187 B.t21 14.4307
R1857 B.n1146 B.t1 14.4307
R1858 B.n1078 B.n129 10.6151
R1859 B.n187 B.n129 10.6151
R1860 B.n188 B.n187 10.6151
R1861 B.n191 B.n188 10.6151
R1862 B.n192 B.n191 10.6151
R1863 B.n195 B.n192 10.6151
R1864 B.n196 B.n195 10.6151
R1865 B.n199 B.n196 10.6151
R1866 B.n200 B.n199 10.6151
R1867 B.n203 B.n200 10.6151
R1868 B.n204 B.n203 10.6151
R1869 B.n207 B.n204 10.6151
R1870 B.n208 B.n207 10.6151
R1871 B.n211 B.n208 10.6151
R1872 B.n212 B.n211 10.6151
R1873 B.n215 B.n212 10.6151
R1874 B.n216 B.n215 10.6151
R1875 B.n219 B.n216 10.6151
R1876 B.n220 B.n219 10.6151
R1877 B.n223 B.n220 10.6151
R1878 B.n224 B.n223 10.6151
R1879 B.n227 B.n224 10.6151
R1880 B.n228 B.n227 10.6151
R1881 B.n231 B.n228 10.6151
R1882 B.n232 B.n231 10.6151
R1883 B.n235 B.n232 10.6151
R1884 B.n236 B.n235 10.6151
R1885 B.n239 B.n236 10.6151
R1886 B.n240 B.n239 10.6151
R1887 B.n243 B.n240 10.6151
R1888 B.n244 B.n243 10.6151
R1889 B.n247 B.n244 10.6151
R1890 B.n248 B.n247 10.6151
R1891 B.n251 B.n248 10.6151
R1892 B.n252 B.n251 10.6151
R1893 B.n255 B.n252 10.6151
R1894 B.n256 B.n255 10.6151
R1895 B.n259 B.n256 10.6151
R1896 B.n260 B.n259 10.6151
R1897 B.n263 B.n260 10.6151
R1898 B.n264 B.n263 10.6151
R1899 B.n267 B.n264 10.6151
R1900 B.n268 B.n267 10.6151
R1901 B.n271 B.n268 10.6151
R1902 B.n276 B.n273 10.6151
R1903 B.n277 B.n276 10.6151
R1904 B.n280 B.n277 10.6151
R1905 B.n281 B.n280 10.6151
R1906 B.n284 B.n281 10.6151
R1907 B.n285 B.n284 10.6151
R1908 B.n288 B.n285 10.6151
R1909 B.n289 B.n288 10.6151
R1910 B.n293 B.n292 10.6151
R1911 B.n296 B.n293 10.6151
R1912 B.n297 B.n296 10.6151
R1913 B.n300 B.n297 10.6151
R1914 B.n301 B.n300 10.6151
R1915 B.n304 B.n301 10.6151
R1916 B.n305 B.n304 10.6151
R1917 B.n308 B.n305 10.6151
R1918 B.n309 B.n308 10.6151
R1919 B.n312 B.n309 10.6151
R1920 B.n313 B.n312 10.6151
R1921 B.n316 B.n313 10.6151
R1922 B.n317 B.n316 10.6151
R1923 B.n320 B.n317 10.6151
R1924 B.n321 B.n320 10.6151
R1925 B.n324 B.n321 10.6151
R1926 B.n325 B.n324 10.6151
R1927 B.n328 B.n325 10.6151
R1928 B.n329 B.n328 10.6151
R1929 B.n332 B.n329 10.6151
R1930 B.n333 B.n332 10.6151
R1931 B.n336 B.n333 10.6151
R1932 B.n337 B.n336 10.6151
R1933 B.n340 B.n337 10.6151
R1934 B.n341 B.n340 10.6151
R1935 B.n344 B.n341 10.6151
R1936 B.n345 B.n344 10.6151
R1937 B.n348 B.n345 10.6151
R1938 B.n349 B.n348 10.6151
R1939 B.n352 B.n349 10.6151
R1940 B.n353 B.n352 10.6151
R1941 B.n356 B.n353 10.6151
R1942 B.n357 B.n356 10.6151
R1943 B.n360 B.n357 10.6151
R1944 B.n361 B.n360 10.6151
R1945 B.n364 B.n361 10.6151
R1946 B.n365 B.n364 10.6151
R1947 B.n368 B.n365 10.6151
R1948 B.n369 B.n368 10.6151
R1949 B.n372 B.n369 10.6151
R1950 B.n373 B.n372 10.6151
R1951 B.n376 B.n373 10.6151
R1952 B.n377 B.n376 10.6151
R1953 B.n1073 B.n377 10.6151
R1954 B.n774 B.n511 10.6151
R1955 B.n775 B.n774 10.6151
R1956 B.n776 B.n775 10.6151
R1957 B.n776 B.n503 10.6151
R1958 B.n786 B.n503 10.6151
R1959 B.n787 B.n786 10.6151
R1960 B.n788 B.n787 10.6151
R1961 B.n788 B.n496 10.6151
R1962 B.n799 B.n496 10.6151
R1963 B.n800 B.n799 10.6151
R1964 B.n801 B.n800 10.6151
R1965 B.n801 B.n488 10.6151
R1966 B.n811 B.n488 10.6151
R1967 B.n812 B.n811 10.6151
R1968 B.n813 B.n812 10.6151
R1969 B.n813 B.n480 10.6151
R1970 B.n823 B.n480 10.6151
R1971 B.n824 B.n823 10.6151
R1972 B.n825 B.n824 10.6151
R1973 B.n825 B.n471 10.6151
R1974 B.n835 B.n471 10.6151
R1975 B.n836 B.n835 10.6151
R1976 B.n837 B.n836 10.6151
R1977 B.n837 B.n464 10.6151
R1978 B.n847 B.n464 10.6151
R1979 B.n848 B.n847 10.6151
R1980 B.n849 B.n848 10.6151
R1981 B.n849 B.n456 10.6151
R1982 B.n859 B.n456 10.6151
R1983 B.n860 B.n859 10.6151
R1984 B.n861 B.n860 10.6151
R1985 B.n861 B.n449 10.6151
R1986 B.n872 B.n449 10.6151
R1987 B.n873 B.n872 10.6151
R1988 B.n874 B.n873 10.6151
R1989 B.n874 B.n441 10.6151
R1990 B.n884 B.n441 10.6151
R1991 B.n885 B.n884 10.6151
R1992 B.n886 B.n885 10.6151
R1993 B.n886 B.n433 10.6151
R1994 B.n896 B.n433 10.6151
R1995 B.n897 B.n896 10.6151
R1996 B.n898 B.n897 10.6151
R1997 B.n898 B.n425 10.6151
R1998 B.n908 B.n425 10.6151
R1999 B.n909 B.n908 10.6151
R2000 B.n910 B.n909 10.6151
R2001 B.n910 B.n417 10.6151
R2002 B.n920 B.n417 10.6151
R2003 B.n921 B.n920 10.6151
R2004 B.n922 B.n921 10.6151
R2005 B.n922 B.n409 10.6151
R2006 B.n932 B.n409 10.6151
R2007 B.n933 B.n932 10.6151
R2008 B.n934 B.n933 10.6151
R2009 B.n934 B.n401 10.6151
R2010 B.n944 B.n401 10.6151
R2011 B.n945 B.n944 10.6151
R2012 B.n946 B.n945 10.6151
R2013 B.n946 B.n393 10.6151
R2014 B.n956 B.n393 10.6151
R2015 B.n957 B.n956 10.6151
R2016 B.n958 B.n957 10.6151
R2017 B.n958 B.n386 10.6151
R2018 B.n969 B.n386 10.6151
R2019 B.n970 B.n969 10.6151
R2020 B.n972 B.n970 10.6151
R2021 B.n972 B.n971 10.6151
R2022 B.n971 B.n378 10.6151
R2023 B.n983 B.n378 10.6151
R2024 B.n984 B.n983 10.6151
R2025 B.n985 B.n984 10.6151
R2026 B.n986 B.n985 10.6151
R2027 B.n988 B.n986 10.6151
R2028 B.n989 B.n988 10.6151
R2029 B.n990 B.n989 10.6151
R2030 B.n991 B.n990 10.6151
R2031 B.n993 B.n991 10.6151
R2032 B.n994 B.n993 10.6151
R2033 B.n995 B.n994 10.6151
R2034 B.n996 B.n995 10.6151
R2035 B.n998 B.n996 10.6151
R2036 B.n999 B.n998 10.6151
R2037 B.n1000 B.n999 10.6151
R2038 B.n1001 B.n1000 10.6151
R2039 B.n1003 B.n1001 10.6151
R2040 B.n1004 B.n1003 10.6151
R2041 B.n1005 B.n1004 10.6151
R2042 B.n1006 B.n1005 10.6151
R2043 B.n1008 B.n1006 10.6151
R2044 B.n1009 B.n1008 10.6151
R2045 B.n1010 B.n1009 10.6151
R2046 B.n1011 B.n1010 10.6151
R2047 B.n1013 B.n1011 10.6151
R2048 B.n1014 B.n1013 10.6151
R2049 B.n1015 B.n1014 10.6151
R2050 B.n1016 B.n1015 10.6151
R2051 B.n1018 B.n1016 10.6151
R2052 B.n1019 B.n1018 10.6151
R2053 B.n1020 B.n1019 10.6151
R2054 B.n1021 B.n1020 10.6151
R2055 B.n1023 B.n1021 10.6151
R2056 B.n1024 B.n1023 10.6151
R2057 B.n1025 B.n1024 10.6151
R2058 B.n1026 B.n1025 10.6151
R2059 B.n1028 B.n1026 10.6151
R2060 B.n1029 B.n1028 10.6151
R2061 B.n1030 B.n1029 10.6151
R2062 B.n1031 B.n1030 10.6151
R2063 B.n1033 B.n1031 10.6151
R2064 B.n1034 B.n1033 10.6151
R2065 B.n1035 B.n1034 10.6151
R2066 B.n1036 B.n1035 10.6151
R2067 B.n1038 B.n1036 10.6151
R2068 B.n1039 B.n1038 10.6151
R2069 B.n1040 B.n1039 10.6151
R2070 B.n1041 B.n1040 10.6151
R2071 B.n1043 B.n1041 10.6151
R2072 B.n1044 B.n1043 10.6151
R2073 B.n1045 B.n1044 10.6151
R2074 B.n1046 B.n1045 10.6151
R2075 B.n1048 B.n1046 10.6151
R2076 B.n1049 B.n1048 10.6151
R2077 B.n1050 B.n1049 10.6151
R2078 B.n1051 B.n1050 10.6151
R2079 B.n1053 B.n1051 10.6151
R2080 B.n1054 B.n1053 10.6151
R2081 B.n1055 B.n1054 10.6151
R2082 B.n1056 B.n1055 10.6151
R2083 B.n1058 B.n1056 10.6151
R2084 B.n1059 B.n1058 10.6151
R2085 B.n1060 B.n1059 10.6151
R2086 B.n1061 B.n1060 10.6151
R2087 B.n1063 B.n1061 10.6151
R2088 B.n1064 B.n1063 10.6151
R2089 B.n1065 B.n1064 10.6151
R2090 B.n1066 B.n1065 10.6151
R2091 B.n1068 B.n1066 10.6151
R2092 B.n1069 B.n1068 10.6151
R2093 B.n1070 B.n1069 10.6151
R2094 B.n1071 B.n1070 10.6151
R2095 B.n1072 B.n1071 10.6151
R2096 B.n768 B.n515 10.6151
R2097 B.n763 B.n515 10.6151
R2098 B.n763 B.n762 10.6151
R2099 B.n762 B.n761 10.6151
R2100 B.n761 B.n758 10.6151
R2101 B.n758 B.n757 10.6151
R2102 B.n757 B.n754 10.6151
R2103 B.n754 B.n753 10.6151
R2104 B.n753 B.n750 10.6151
R2105 B.n750 B.n749 10.6151
R2106 B.n749 B.n746 10.6151
R2107 B.n746 B.n745 10.6151
R2108 B.n745 B.n742 10.6151
R2109 B.n742 B.n741 10.6151
R2110 B.n741 B.n738 10.6151
R2111 B.n738 B.n737 10.6151
R2112 B.n737 B.n734 10.6151
R2113 B.n734 B.n733 10.6151
R2114 B.n733 B.n730 10.6151
R2115 B.n730 B.n729 10.6151
R2116 B.n729 B.n726 10.6151
R2117 B.n726 B.n725 10.6151
R2118 B.n725 B.n722 10.6151
R2119 B.n722 B.n721 10.6151
R2120 B.n721 B.n718 10.6151
R2121 B.n718 B.n717 10.6151
R2122 B.n717 B.n714 10.6151
R2123 B.n714 B.n713 10.6151
R2124 B.n713 B.n710 10.6151
R2125 B.n710 B.n709 10.6151
R2126 B.n709 B.n706 10.6151
R2127 B.n706 B.n705 10.6151
R2128 B.n705 B.n702 10.6151
R2129 B.n702 B.n701 10.6151
R2130 B.n701 B.n698 10.6151
R2131 B.n698 B.n697 10.6151
R2132 B.n697 B.n694 10.6151
R2133 B.n694 B.n693 10.6151
R2134 B.n693 B.n690 10.6151
R2135 B.n690 B.n689 10.6151
R2136 B.n689 B.n686 10.6151
R2137 B.n686 B.n685 10.6151
R2138 B.n685 B.n682 10.6151
R2139 B.n682 B.n681 10.6151
R2140 B.n678 B.n677 10.6151
R2141 B.n677 B.n674 10.6151
R2142 B.n674 B.n673 10.6151
R2143 B.n673 B.n670 10.6151
R2144 B.n670 B.n669 10.6151
R2145 B.n669 B.n666 10.6151
R2146 B.n666 B.n665 10.6151
R2147 B.n665 B.n662 10.6151
R2148 B.n660 B.n657 10.6151
R2149 B.n657 B.n656 10.6151
R2150 B.n656 B.n653 10.6151
R2151 B.n653 B.n652 10.6151
R2152 B.n652 B.n649 10.6151
R2153 B.n649 B.n648 10.6151
R2154 B.n648 B.n645 10.6151
R2155 B.n645 B.n644 10.6151
R2156 B.n644 B.n641 10.6151
R2157 B.n641 B.n640 10.6151
R2158 B.n640 B.n637 10.6151
R2159 B.n637 B.n636 10.6151
R2160 B.n636 B.n633 10.6151
R2161 B.n633 B.n632 10.6151
R2162 B.n632 B.n629 10.6151
R2163 B.n629 B.n628 10.6151
R2164 B.n628 B.n625 10.6151
R2165 B.n625 B.n624 10.6151
R2166 B.n624 B.n621 10.6151
R2167 B.n621 B.n620 10.6151
R2168 B.n620 B.n617 10.6151
R2169 B.n617 B.n616 10.6151
R2170 B.n616 B.n613 10.6151
R2171 B.n613 B.n612 10.6151
R2172 B.n612 B.n609 10.6151
R2173 B.n609 B.n608 10.6151
R2174 B.n608 B.n605 10.6151
R2175 B.n605 B.n604 10.6151
R2176 B.n604 B.n601 10.6151
R2177 B.n601 B.n600 10.6151
R2178 B.n600 B.n597 10.6151
R2179 B.n597 B.n596 10.6151
R2180 B.n596 B.n593 10.6151
R2181 B.n593 B.n592 10.6151
R2182 B.n592 B.n589 10.6151
R2183 B.n589 B.n588 10.6151
R2184 B.n588 B.n585 10.6151
R2185 B.n585 B.n584 10.6151
R2186 B.n584 B.n581 10.6151
R2187 B.n581 B.n580 10.6151
R2188 B.n580 B.n577 10.6151
R2189 B.n577 B.n576 10.6151
R2190 B.n576 B.n573 10.6151
R2191 B.n573 B.n572 10.6151
R2192 B.n770 B.n769 10.6151
R2193 B.n770 B.n507 10.6151
R2194 B.n780 B.n507 10.6151
R2195 B.n781 B.n780 10.6151
R2196 B.n782 B.n781 10.6151
R2197 B.n782 B.n499 10.6151
R2198 B.n793 B.n499 10.6151
R2199 B.n794 B.n793 10.6151
R2200 B.n795 B.n794 10.6151
R2201 B.n795 B.n492 10.6151
R2202 B.n805 B.n492 10.6151
R2203 B.n806 B.n805 10.6151
R2204 B.n807 B.n806 10.6151
R2205 B.n807 B.n484 10.6151
R2206 B.n817 B.n484 10.6151
R2207 B.n818 B.n817 10.6151
R2208 B.n819 B.n818 10.6151
R2209 B.n819 B.n476 10.6151
R2210 B.n829 B.n476 10.6151
R2211 B.n830 B.n829 10.6151
R2212 B.n831 B.n830 10.6151
R2213 B.n831 B.n468 10.6151
R2214 B.n841 B.n468 10.6151
R2215 B.n842 B.n841 10.6151
R2216 B.n843 B.n842 10.6151
R2217 B.n843 B.n460 10.6151
R2218 B.n853 B.n460 10.6151
R2219 B.n854 B.n853 10.6151
R2220 B.n855 B.n854 10.6151
R2221 B.n855 B.n452 10.6151
R2222 B.n866 B.n452 10.6151
R2223 B.n867 B.n866 10.6151
R2224 B.n868 B.n867 10.6151
R2225 B.n868 B.n445 10.6151
R2226 B.n878 B.n445 10.6151
R2227 B.n879 B.n878 10.6151
R2228 B.n880 B.n879 10.6151
R2229 B.n880 B.n437 10.6151
R2230 B.n890 B.n437 10.6151
R2231 B.n891 B.n890 10.6151
R2232 B.n892 B.n891 10.6151
R2233 B.n892 B.n429 10.6151
R2234 B.n902 B.n429 10.6151
R2235 B.n903 B.n902 10.6151
R2236 B.n904 B.n903 10.6151
R2237 B.n904 B.n421 10.6151
R2238 B.n914 B.n421 10.6151
R2239 B.n915 B.n914 10.6151
R2240 B.n916 B.n915 10.6151
R2241 B.n916 B.n413 10.6151
R2242 B.n926 B.n413 10.6151
R2243 B.n927 B.n926 10.6151
R2244 B.n928 B.n927 10.6151
R2245 B.n928 B.n405 10.6151
R2246 B.n938 B.n405 10.6151
R2247 B.n939 B.n938 10.6151
R2248 B.n940 B.n939 10.6151
R2249 B.n940 B.n397 10.6151
R2250 B.n950 B.n397 10.6151
R2251 B.n951 B.n950 10.6151
R2252 B.n952 B.n951 10.6151
R2253 B.n952 B.n389 10.6151
R2254 B.n963 B.n389 10.6151
R2255 B.n964 B.n963 10.6151
R2256 B.n965 B.n964 10.6151
R2257 B.n965 B.n382 10.6151
R2258 B.n976 B.n382 10.6151
R2259 B.n977 B.n976 10.6151
R2260 B.n978 B.n977 10.6151
R2261 B.n978 B.n0 10.6151
R2262 B.n1216 B.n1 10.6151
R2263 B.n1216 B.n1215 10.6151
R2264 B.n1215 B.n1214 10.6151
R2265 B.n1214 B.n10 10.6151
R2266 B.n1208 B.n10 10.6151
R2267 B.n1208 B.n1207 10.6151
R2268 B.n1207 B.n1206 10.6151
R2269 B.n1206 B.n16 10.6151
R2270 B.n1200 B.n16 10.6151
R2271 B.n1200 B.n1199 10.6151
R2272 B.n1199 B.n1198 10.6151
R2273 B.n1198 B.n24 10.6151
R2274 B.n1192 B.n24 10.6151
R2275 B.n1192 B.n1191 10.6151
R2276 B.n1191 B.n1190 10.6151
R2277 B.n1190 B.n31 10.6151
R2278 B.n1184 B.n31 10.6151
R2279 B.n1184 B.n1183 10.6151
R2280 B.n1183 B.n1182 10.6151
R2281 B.n1182 B.n38 10.6151
R2282 B.n1176 B.n38 10.6151
R2283 B.n1176 B.n1175 10.6151
R2284 B.n1175 B.n1174 10.6151
R2285 B.n1174 B.n45 10.6151
R2286 B.n1168 B.n45 10.6151
R2287 B.n1168 B.n1167 10.6151
R2288 B.n1167 B.n1166 10.6151
R2289 B.n1166 B.n52 10.6151
R2290 B.n1160 B.n52 10.6151
R2291 B.n1160 B.n1159 10.6151
R2292 B.n1159 B.n1158 10.6151
R2293 B.n1158 B.n59 10.6151
R2294 B.n1152 B.n59 10.6151
R2295 B.n1152 B.n1151 10.6151
R2296 B.n1151 B.n1150 10.6151
R2297 B.n1150 B.n66 10.6151
R2298 B.n1144 B.n66 10.6151
R2299 B.n1144 B.n1143 10.6151
R2300 B.n1143 B.n1142 10.6151
R2301 B.n1142 B.n72 10.6151
R2302 B.n1136 B.n72 10.6151
R2303 B.n1136 B.n1135 10.6151
R2304 B.n1135 B.n1134 10.6151
R2305 B.n1134 B.n80 10.6151
R2306 B.n1128 B.n80 10.6151
R2307 B.n1128 B.n1127 10.6151
R2308 B.n1127 B.n1126 10.6151
R2309 B.n1126 B.n87 10.6151
R2310 B.n1120 B.n87 10.6151
R2311 B.n1120 B.n1119 10.6151
R2312 B.n1119 B.n1118 10.6151
R2313 B.n1118 B.n94 10.6151
R2314 B.n1112 B.n94 10.6151
R2315 B.n1112 B.n1111 10.6151
R2316 B.n1111 B.n1110 10.6151
R2317 B.n1110 B.n101 10.6151
R2318 B.n1104 B.n101 10.6151
R2319 B.n1104 B.n1103 10.6151
R2320 B.n1103 B.n1102 10.6151
R2321 B.n1102 B.n108 10.6151
R2322 B.n1096 B.n108 10.6151
R2323 B.n1096 B.n1095 10.6151
R2324 B.n1095 B.n1094 10.6151
R2325 B.n1094 B.n114 10.6151
R2326 B.n1088 B.n114 10.6151
R2327 B.n1088 B.n1087 10.6151
R2328 B.n1087 B.n1086 10.6151
R2329 B.n1086 B.n122 10.6151
R2330 B.n1080 B.n122 10.6151
R2331 B.n1080 B.n1079 10.6151
R2332 B.n273 B.n272 6.5566
R2333 B.n289 B.n183 6.5566
R2334 B.n678 B.n568 6.5566
R2335 B.n662 B.n661 6.5566
R2336 B.n474 B.t0 6.01307
R2337 B.n900 B.t23 6.01307
R2338 B.n960 B.t19 6.01307
R2339 B.n18 B.t22 6.01307
R2340 B.n1164 B.t18 6.01307
R2341 B.t2 B.n1123 6.01307
R2342 B.n272 B.n271 4.05904
R2343 B.n292 B.n183 4.05904
R2344 B.n681 B.n568 4.05904
R2345 B.n661 B.n660 4.05904
R2346 B.n1222 B.n0 2.81026
R2347 B.n1222 B.n1 2.81026
R2348 VN.n94 VN.n93 161.3
R2349 VN.n92 VN.n49 161.3
R2350 VN.n91 VN.n90 161.3
R2351 VN.n89 VN.n50 161.3
R2352 VN.n88 VN.n87 161.3
R2353 VN.n86 VN.n51 161.3
R2354 VN.n85 VN.n84 161.3
R2355 VN.n83 VN.n82 161.3
R2356 VN.n81 VN.n53 161.3
R2357 VN.n80 VN.n79 161.3
R2358 VN.n78 VN.n54 161.3
R2359 VN.n77 VN.n76 161.3
R2360 VN.n75 VN.n55 161.3
R2361 VN.n74 VN.n73 161.3
R2362 VN.n72 VN.n71 161.3
R2363 VN.n70 VN.n57 161.3
R2364 VN.n69 VN.n68 161.3
R2365 VN.n67 VN.n58 161.3
R2366 VN.n66 VN.n65 161.3
R2367 VN.n64 VN.n59 161.3
R2368 VN.n63 VN.n62 161.3
R2369 VN.n46 VN.n45 161.3
R2370 VN.n44 VN.n1 161.3
R2371 VN.n43 VN.n42 161.3
R2372 VN.n41 VN.n2 161.3
R2373 VN.n40 VN.n39 161.3
R2374 VN.n38 VN.n3 161.3
R2375 VN.n37 VN.n36 161.3
R2376 VN.n35 VN.n34 161.3
R2377 VN.n33 VN.n5 161.3
R2378 VN.n32 VN.n31 161.3
R2379 VN.n30 VN.n6 161.3
R2380 VN.n29 VN.n28 161.3
R2381 VN.n27 VN.n7 161.3
R2382 VN.n26 VN.n25 161.3
R2383 VN.n24 VN.n23 161.3
R2384 VN.n22 VN.n9 161.3
R2385 VN.n21 VN.n20 161.3
R2386 VN.n19 VN.n10 161.3
R2387 VN.n18 VN.n17 161.3
R2388 VN.n16 VN.n11 161.3
R2389 VN.n15 VN.n14 161.3
R2390 VN.n61 VN.t6 130.256
R2391 VN.n13 VN.t1 130.256
R2392 VN.n12 VN.t0 96.8468
R2393 VN.n8 VN.t8 96.8468
R2394 VN.n4 VN.t5 96.8468
R2395 VN.n0 VN.t3 96.8468
R2396 VN.n60 VN.t9 96.8468
R2397 VN.n56 VN.t2 96.8468
R2398 VN.n52 VN.t4 96.8468
R2399 VN.n48 VN.t7 96.8468
R2400 VN.n47 VN.n0 71.0639
R2401 VN.n95 VN.n48 71.0639
R2402 VN.n13 VN.n12 58.6193
R2403 VN.n61 VN.n60 58.6193
R2404 VN VN.n95 57.6989
R2405 VN.n43 VN.n2 50.7491
R2406 VN.n91 VN.n50 50.7491
R2407 VN.n17 VN.n10 43.9677
R2408 VN.n32 VN.n6 43.9677
R2409 VN.n65 VN.n58 43.9677
R2410 VN.n80 VN.n54 43.9677
R2411 VN.n21 VN.n10 37.1863
R2412 VN.n28 VN.n6 37.1863
R2413 VN.n69 VN.n58 37.1863
R2414 VN.n76 VN.n54 37.1863
R2415 VN.n39 VN.n2 30.405
R2416 VN.n87 VN.n50 30.405
R2417 VN.n16 VN.n15 24.5923
R2418 VN.n17 VN.n16 24.5923
R2419 VN.n22 VN.n21 24.5923
R2420 VN.n23 VN.n22 24.5923
R2421 VN.n27 VN.n26 24.5923
R2422 VN.n28 VN.n27 24.5923
R2423 VN.n33 VN.n32 24.5923
R2424 VN.n34 VN.n33 24.5923
R2425 VN.n38 VN.n37 24.5923
R2426 VN.n39 VN.n38 24.5923
R2427 VN.n44 VN.n43 24.5923
R2428 VN.n45 VN.n44 24.5923
R2429 VN.n65 VN.n64 24.5923
R2430 VN.n64 VN.n63 24.5923
R2431 VN.n76 VN.n75 24.5923
R2432 VN.n75 VN.n74 24.5923
R2433 VN.n71 VN.n70 24.5923
R2434 VN.n70 VN.n69 24.5923
R2435 VN.n87 VN.n86 24.5923
R2436 VN.n86 VN.n85 24.5923
R2437 VN.n82 VN.n81 24.5923
R2438 VN.n81 VN.n80 24.5923
R2439 VN.n93 VN.n92 24.5923
R2440 VN.n92 VN.n91 24.5923
R2441 VN.n45 VN.n0 19.1821
R2442 VN.n93 VN.n48 19.1821
R2443 VN.n15 VN.n12 15.7393
R2444 VN.n34 VN.n4 15.7393
R2445 VN.n63 VN.n60 15.7393
R2446 VN.n82 VN.n52 15.7393
R2447 VN.n23 VN.n8 12.2964
R2448 VN.n26 VN.n8 12.2964
R2449 VN.n74 VN.n56 12.2964
R2450 VN.n71 VN.n56 12.2964
R2451 VN.n37 VN.n4 8.85356
R2452 VN.n85 VN.n52 8.85356
R2453 VN.n14 VN.n13 3.93513
R2454 VN.n62 VN.n61 3.93513
R2455 VN.n95 VN.n94 0.354861
R2456 VN.n47 VN.n46 0.354861
R2457 VN VN.n47 0.267071
R2458 VN.n94 VN.n49 0.189894
R2459 VN.n90 VN.n49 0.189894
R2460 VN.n90 VN.n89 0.189894
R2461 VN.n89 VN.n88 0.189894
R2462 VN.n88 VN.n51 0.189894
R2463 VN.n84 VN.n51 0.189894
R2464 VN.n84 VN.n83 0.189894
R2465 VN.n83 VN.n53 0.189894
R2466 VN.n79 VN.n53 0.189894
R2467 VN.n79 VN.n78 0.189894
R2468 VN.n78 VN.n77 0.189894
R2469 VN.n77 VN.n55 0.189894
R2470 VN.n73 VN.n55 0.189894
R2471 VN.n73 VN.n72 0.189894
R2472 VN.n72 VN.n57 0.189894
R2473 VN.n68 VN.n57 0.189894
R2474 VN.n68 VN.n67 0.189894
R2475 VN.n67 VN.n66 0.189894
R2476 VN.n66 VN.n59 0.189894
R2477 VN.n62 VN.n59 0.189894
R2478 VN.n14 VN.n11 0.189894
R2479 VN.n18 VN.n11 0.189894
R2480 VN.n19 VN.n18 0.189894
R2481 VN.n20 VN.n19 0.189894
R2482 VN.n20 VN.n9 0.189894
R2483 VN.n24 VN.n9 0.189894
R2484 VN.n25 VN.n24 0.189894
R2485 VN.n25 VN.n7 0.189894
R2486 VN.n29 VN.n7 0.189894
R2487 VN.n30 VN.n29 0.189894
R2488 VN.n31 VN.n30 0.189894
R2489 VN.n31 VN.n5 0.189894
R2490 VN.n35 VN.n5 0.189894
R2491 VN.n36 VN.n35 0.189894
R2492 VN.n36 VN.n3 0.189894
R2493 VN.n40 VN.n3 0.189894
R2494 VN.n41 VN.n40 0.189894
R2495 VN.n42 VN.n41 0.189894
R2496 VN.n42 VN.n1 0.189894
R2497 VN.n46 VN.n1 0.189894
R2498 VDD2.n1 VDD2.t8 69.265
R2499 VDD2.n3 VDD2.n2 66.9195
R2500 VDD2 VDD2.n7 66.9167
R2501 VDD2.n4 VDD2.t2 66.1886
R2502 VDD2.n6 VDD2.n5 64.6679
R2503 VDD2.n1 VDD2.n0 64.6667
R2504 VDD2.n4 VDD2.n3 49.558
R2505 VDD2.n6 VDD2.n4 3.07809
R2506 VDD2.n7 VDD2.t0 1.52124
R2507 VDD2.n7 VDD2.t3 1.52124
R2508 VDD2.n5 VDD2.t5 1.52124
R2509 VDD2.n5 VDD2.t7 1.52124
R2510 VDD2.n2 VDD2.t4 1.52124
R2511 VDD2.n2 VDD2.t6 1.52124
R2512 VDD2.n0 VDD2.t9 1.52124
R2513 VDD2.n0 VDD2.t1 1.52124
R2514 VDD2 VDD2.n6 0.828086
R2515 VDD2.n3 VDD2.n1 0.714551
C0 VTAIL VP 12.8882f
C1 VN VDD1 0.154973f
C2 VN VDD2 12.004f
C3 VDD1 VP 12.510401f
C4 VTAIL VDD1 11.0688f
C5 VDD2 VP 0.66545f
C6 VTAIL VDD2 11.1244f
C7 VDD1 VDD2 2.59006f
C8 VN VP 9.52192f
C9 VN VTAIL 12.8739f
C10 VDD2 B 8.125386f
C11 VDD1 B 8.104184f
C12 VTAIL B 9.106122f
C13 VN B 21.26243f
C14 VP B 19.823484f
C15 VDD2.t8 B 2.89568f
C16 VDD2.t9 B 0.250475f
C17 VDD2.t1 B 0.250475f
C18 VDD2.n0 B 2.25174f
C19 VDD2.n1 B 0.975636f
C20 VDD2.t4 B 0.250475f
C21 VDD2.t6 B 0.250475f
C22 VDD2.n2 B 2.27267f
C23 VDD2.n3 B 3.20978f
C24 VDD2.t2 B 2.87319f
C25 VDD2.n4 B 3.35153f
C26 VDD2.t5 B 0.250475f
C27 VDD2.t7 B 0.250475f
C28 VDD2.n5 B 2.25175f
C29 VDD2.n6 B 0.499837f
C30 VDD2.t0 B 0.250475f
C31 VDD2.t3 B 0.250475f
C32 VDD2.n7 B 2.27263f
C33 VN.t3 B 2.11894f
C34 VN.n0 B 0.817823f
C35 VN.n1 B 0.018394f
C36 VN.n2 B 0.017615f
C37 VN.n3 B 0.018394f
C38 VN.t5 B 2.11894f
C39 VN.n4 B 0.74171f
C40 VN.n5 B 0.018394f
C41 VN.n6 B 0.015146f
C42 VN.n7 B 0.018394f
C43 VN.t8 B 2.11894f
C44 VN.n8 B 0.74171f
C45 VN.n9 B 0.018394f
C46 VN.n10 B 0.015146f
C47 VN.n11 B 0.018394f
C48 VN.t0 B 2.11894f
C49 VN.n12 B 0.804432f
C50 VN.t1 B 2.34326f
C51 VN.n13 B 0.766167f
C52 VN.n14 B 0.212996f
C53 VN.n15 B 0.028048f
C54 VN.n16 B 0.034111f
C55 VN.n17 B 0.035595f
C56 VN.n18 B 0.018394f
C57 VN.n19 B 0.018394f
C58 VN.n20 B 0.018394f
C59 VN.n21 B 0.036848f
C60 VN.n22 B 0.034111f
C61 VN.n23 B 0.025691f
C62 VN.n24 B 0.018394f
C63 VN.n25 B 0.018394f
C64 VN.n26 B 0.025691f
C65 VN.n27 B 0.034111f
C66 VN.n28 B 0.036848f
C67 VN.n29 B 0.018394f
C68 VN.n30 B 0.018394f
C69 VN.n31 B 0.018394f
C70 VN.n32 B 0.035595f
C71 VN.n33 B 0.034111f
C72 VN.n34 B 0.028048f
C73 VN.n35 B 0.018394f
C74 VN.n36 B 0.018394f
C75 VN.n37 B 0.023333f
C76 VN.n38 B 0.034111f
C77 VN.n39 B 0.036557f
C78 VN.n40 B 0.018394f
C79 VN.n41 B 0.018394f
C80 VN.n42 B 0.018394f
C81 VN.n43 B 0.033416f
C82 VN.n44 B 0.034111f
C83 VN.n45 B 0.030406f
C84 VN.n46 B 0.029683f
C85 VN.n47 B 0.040514f
C86 VN.t7 B 2.11894f
C87 VN.n48 B 0.817823f
C88 VN.n49 B 0.018394f
C89 VN.n50 B 0.017615f
C90 VN.n51 B 0.018394f
C91 VN.t4 B 2.11894f
C92 VN.n52 B 0.74171f
C93 VN.n53 B 0.018394f
C94 VN.n54 B 0.015146f
C95 VN.n55 B 0.018394f
C96 VN.t2 B 2.11894f
C97 VN.n56 B 0.74171f
C98 VN.n57 B 0.018394f
C99 VN.n58 B 0.015146f
C100 VN.n59 B 0.018394f
C101 VN.t9 B 2.11894f
C102 VN.n60 B 0.804432f
C103 VN.t6 B 2.34326f
C104 VN.n61 B 0.766167f
C105 VN.n62 B 0.212996f
C106 VN.n63 B 0.028048f
C107 VN.n64 B 0.034111f
C108 VN.n65 B 0.035595f
C109 VN.n66 B 0.018394f
C110 VN.n67 B 0.018394f
C111 VN.n68 B 0.018394f
C112 VN.n69 B 0.036848f
C113 VN.n70 B 0.034111f
C114 VN.n71 B 0.025691f
C115 VN.n72 B 0.018394f
C116 VN.n73 B 0.018394f
C117 VN.n74 B 0.025691f
C118 VN.n75 B 0.034111f
C119 VN.n76 B 0.036848f
C120 VN.n77 B 0.018394f
C121 VN.n78 B 0.018394f
C122 VN.n79 B 0.018394f
C123 VN.n80 B 0.035595f
C124 VN.n81 B 0.034111f
C125 VN.n82 B 0.028048f
C126 VN.n83 B 0.018394f
C127 VN.n84 B 0.018394f
C128 VN.n85 B 0.023333f
C129 VN.n86 B 0.034111f
C130 VN.n87 B 0.036557f
C131 VN.n88 B 0.018394f
C132 VN.n89 B 0.018394f
C133 VN.n90 B 0.018394f
C134 VN.n91 B 0.033416f
C135 VN.n92 B 0.034111f
C136 VN.n93 B 0.030406f
C137 VN.n94 B 0.029683f
C138 VN.n95 B 1.27683f
C139 VTAIL.t16 B 0.258711f
C140 VTAIL.t15 B 0.258711f
C141 VTAIL.n0 B 2.25798f
C142 VTAIL.n1 B 0.587973f
C143 VTAIL.t6 B 2.88046f
C144 VTAIL.n2 B 0.728683f
C145 VTAIL.t11 B 0.258711f
C146 VTAIL.t7 B 0.258711f
C147 VTAIL.n3 B 2.25798f
C148 VTAIL.n4 B 0.732207f
C149 VTAIL.t4 B 0.258711f
C150 VTAIL.t3 B 0.258711f
C151 VTAIL.n5 B 2.25798f
C152 VTAIL.n6 B 2.23253f
C153 VTAIL.t0 B 0.258711f
C154 VTAIL.t14 B 0.258711f
C155 VTAIL.n7 B 2.25799f
C156 VTAIL.n8 B 2.23252f
C157 VTAIL.t19 B 0.258711f
C158 VTAIL.t17 B 0.258711f
C159 VTAIL.n9 B 2.25799f
C160 VTAIL.n10 B 0.732196f
C161 VTAIL.t13 B 2.88048f
C162 VTAIL.n11 B 0.728667f
C163 VTAIL.t10 B 0.258711f
C164 VTAIL.t8 B 0.258711f
C165 VTAIL.n12 B 2.25799f
C166 VTAIL.n13 B 0.645586f
C167 VTAIL.t5 B 0.258711f
C168 VTAIL.t12 B 0.258711f
C169 VTAIL.n14 B 2.25799f
C170 VTAIL.n15 B 0.732196f
C171 VTAIL.t9 B 2.88046f
C172 VTAIL.n16 B 2.06626f
C173 VTAIL.t2 B 2.88046f
C174 VTAIL.n17 B 2.06626f
C175 VTAIL.t18 B 0.258711f
C176 VTAIL.t1 B 0.258711f
C177 VTAIL.n18 B 2.25798f
C178 VTAIL.n19 B 0.540477f
C179 VDD1.t6 B 2.94173f
C180 VDD1.t8 B 0.254458f
C181 VDD1.t5 B 0.254458f
C182 VDD1.n0 B 2.28755f
C183 VDD1.n1 B 0.999378f
C184 VDD1.t4 B 2.94172f
C185 VDD1.t1 B 0.254458f
C186 VDD1.t7 B 0.254458f
C187 VDD1.n2 B 2.28755f
C188 VDD1.n3 B 0.99115f
C189 VDD1.t3 B 0.254458f
C190 VDD1.t2 B 0.254458f
C191 VDD1.n4 B 2.30881f
C192 VDD1.n5 B 3.40257f
C193 VDD1.t0 B 0.254458f
C194 VDD1.t9 B 0.254458f
C195 VDD1.n6 B 2.28755f
C196 VDD1.n7 B 3.47108f
C197 VP.t6 B 2.15135f
C198 VP.n0 B 0.830334f
C199 VP.n1 B 0.018676f
C200 VP.n2 B 0.017885f
C201 VP.n3 B 0.018676f
C202 VP.t5 B 2.15135f
C203 VP.n4 B 0.753056f
C204 VP.n5 B 0.018676f
C205 VP.n6 B 0.015377f
C206 VP.n7 B 0.018676f
C207 VP.t1 B 2.15135f
C208 VP.n8 B 0.753056f
C209 VP.n9 B 0.018676f
C210 VP.n10 B 0.015377f
C211 VP.n11 B 0.018676f
C212 VP.t9 B 2.15135f
C213 VP.n12 B 0.753056f
C214 VP.n13 B 0.018676f
C215 VP.n14 B 0.017885f
C216 VP.n15 B 0.018676f
C217 VP.t8 B 2.15135f
C218 VP.n16 B 0.830334f
C219 VP.t3 B 2.15135f
C220 VP.n17 B 0.830334f
C221 VP.n18 B 0.018676f
C222 VP.n19 B 0.017885f
C223 VP.n20 B 0.018676f
C224 VP.t0 B 2.15135f
C225 VP.n21 B 0.753056f
C226 VP.n22 B 0.018676f
C227 VP.n23 B 0.015377f
C228 VP.n24 B 0.018676f
C229 VP.t7 B 2.15135f
C230 VP.n25 B 0.753056f
C231 VP.n26 B 0.018676f
C232 VP.n27 B 0.015377f
C233 VP.n28 B 0.018676f
C234 VP.t4 B 2.15135f
C235 VP.n29 B 0.816738f
C236 VP.t2 B 2.3791f
C237 VP.n30 B 0.777889f
C238 VP.n31 B 0.216255f
C239 VP.n32 B 0.028478f
C240 VP.n33 B 0.034633f
C241 VP.n34 B 0.036139f
C242 VP.n35 B 0.018676f
C243 VP.n36 B 0.018676f
C244 VP.n37 B 0.018676f
C245 VP.n38 B 0.037412f
C246 VP.n39 B 0.034633f
C247 VP.n40 B 0.026084f
C248 VP.n41 B 0.018676f
C249 VP.n42 B 0.018676f
C250 VP.n43 B 0.026084f
C251 VP.n44 B 0.034633f
C252 VP.n45 B 0.037412f
C253 VP.n46 B 0.018676f
C254 VP.n47 B 0.018676f
C255 VP.n48 B 0.018676f
C256 VP.n49 B 0.036139f
C257 VP.n50 B 0.034633f
C258 VP.n51 B 0.028478f
C259 VP.n52 B 0.018676f
C260 VP.n53 B 0.018676f
C261 VP.n54 B 0.02369f
C262 VP.n55 B 0.034633f
C263 VP.n56 B 0.037117f
C264 VP.n57 B 0.018676f
C265 VP.n58 B 0.018676f
C266 VP.n59 B 0.018676f
C267 VP.n60 B 0.033928f
C268 VP.n61 B 0.034633f
C269 VP.n62 B 0.030871f
C270 VP.n63 B 0.030138f
C271 VP.n64 B 1.28907f
C272 VP.n65 B 1.30077f
C273 VP.n66 B 0.030138f
C274 VP.n67 B 0.030871f
C275 VP.n68 B 0.034633f
C276 VP.n69 B 0.033928f
C277 VP.n70 B 0.018676f
C278 VP.n71 B 0.018676f
C279 VP.n72 B 0.018676f
C280 VP.n73 B 0.037117f
C281 VP.n74 B 0.034633f
C282 VP.n75 B 0.02369f
C283 VP.n76 B 0.018676f
C284 VP.n77 B 0.018676f
C285 VP.n78 B 0.028478f
C286 VP.n79 B 0.034633f
C287 VP.n80 B 0.036139f
C288 VP.n81 B 0.018676f
C289 VP.n82 B 0.018676f
C290 VP.n83 B 0.018676f
C291 VP.n84 B 0.037412f
C292 VP.n85 B 0.034633f
C293 VP.n86 B 0.026084f
C294 VP.n87 B 0.018676f
C295 VP.n88 B 0.018676f
C296 VP.n89 B 0.026084f
C297 VP.n90 B 0.034633f
C298 VP.n91 B 0.037412f
C299 VP.n92 B 0.018676f
C300 VP.n93 B 0.018676f
C301 VP.n94 B 0.018676f
C302 VP.n95 B 0.036139f
C303 VP.n96 B 0.034633f
C304 VP.n97 B 0.028478f
C305 VP.n98 B 0.018676f
C306 VP.n99 B 0.018676f
C307 VP.n100 B 0.02369f
C308 VP.n101 B 0.034633f
C309 VP.n102 B 0.037117f
C310 VP.n103 B 0.018676f
C311 VP.n104 B 0.018676f
C312 VP.n105 B 0.018676f
C313 VP.n106 B 0.033928f
C314 VP.n107 B 0.034633f
C315 VP.n108 B 0.030871f
C316 VP.n109 B 0.030138f
C317 VP.n110 B 0.041134f
.ends

