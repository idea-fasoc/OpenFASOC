* NGSPICE file created from diff_pair_sample_1183.ext - technology: sky130A

.subckt diff_pair_sample_1183 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t19 VN.t0 VDD2.t7 w_n2110_n2274# sky130_fd_pr__pfet_01v8 ad=1.07745 pd=6.86 as=1.07745 ps=6.86 w=6.53 l=0.62
X1 VDD2.t8 VN.t1 VTAIL.t18 w_n2110_n2274# sky130_fd_pr__pfet_01v8 ad=2.5467 pd=13.84 as=1.07745 ps=6.86 w=6.53 l=0.62
X2 VDD1.t9 VP.t0 VTAIL.t2 w_n2110_n2274# sky130_fd_pr__pfet_01v8 ad=1.07745 pd=6.86 as=2.5467 ps=13.84 w=6.53 l=0.62
X3 VTAIL.t7 VP.t1 VDD1.t8 w_n2110_n2274# sky130_fd_pr__pfet_01v8 ad=1.07745 pd=6.86 as=1.07745 ps=6.86 w=6.53 l=0.62
X4 B.t11 B.t9 B.t10 w_n2110_n2274# sky130_fd_pr__pfet_01v8 ad=2.5467 pd=13.84 as=0 ps=0 w=6.53 l=0.62
X5 VTAIL.t9 VP.t2 VDD1.t7 w_n2110_n2274# sky130_fd_pr__pfet_01v8 ad=1.07745 pd=6.86 as=1.07745 ps=6.86 w=6.53 l=0.62
X6 VDD1.t6 VP.t3 VTAIL.t6 w_n2110_n2274# sky130_fd_pr__pfet_01v8 ad=2.5467 pd=13.84 as=1.07745 ps=6.86 w=6.53 l=0.62
X7 VDD1.t5 VP.t4 VTAIL.t0 w_n2110_n2274# sky130_fd_pr__pfet_01v8 ad=1.07745 pd=6.86 as=1.07745 ps=6.86 w=6.53 l=0.62
X8 VTAIL.t8 VP.t5 VDD1.t4 w_n2110_n2274# sky130_fd_pr__pfet_01v8 ad=1.07745 pd=6.86 as=1.07745 ps=6.86 w=6.53 l=0.62
X9 B.t8 B.t6 B.t7 w_n2110_n2274# sky130_fd_pr__pfet_01v8 ad=2.5467 pd=13.84 as=0 ps=0 w=6.53 l=0.62
X10 VDD1.t3 VP.t6 VTAIL.t1 w_n2110_n2274# sky130_fd_pr__pfet_01v8 ad=2.5467 pd=13.84 as=1.07745 ps=6.86 w=6.53 l=0.62
X11 VDD2.t5 VN.t2 VTAIL.t17 w_n2110_n2274# sky130_fd_pr__pfet_01v8 ad=1.07745 pd=6.86 as=2.5467 ps=13.84 w=6.53 l=0.62
X12 VTAIL.t16 VN.t3 VDD2.t4 w_n2110_n2274# sky130_fd_pr__pfet_01v8 ad=1.07745 pd=6.86 as=1.07745 ps=6.86 w=6.53 l=0.62
X13 VDD1.t2 VP.t7 VTAIL.t4 w_n2110_n2274# sky130_fd_pr__pfet_01v8 ad=1.07745 pd=6.86 as=1.07745 ps=6.86 w=6.53 l=0.62
X14 VDD2.t3 VN.t4 VTAIL.t15 w_n2110_n2274# sky130_fd_pr__pfet_01v8 ad=2.5467 pd=13.84 as=1.07745 ps=6.86 w=6.53 l=0.62
X15 VTAIL.t14 VN.t5 VDD2.t9 w_n2110_n2274# sky130_fd_pr__pfet_01v8 ad=1.07745 pd=6.86 as=1.07745 ps=6.86 w=6.53 l=0.62
X16 VDD2.t6 VN.t6 VTAIL.t13 w_n2110_n2274# sky130_fd_pr__pfet_01v8 ad=1.07745 pd=6.86 as=1.07745 ps=6.86 w=6.53 l=0.62
X17 VDD2.t0 VN.t7 VTAIL.t12 w_n2110_n2274# sky130_fd_pr__pfet_01v8 ad=1.07745 pd=6.86 as=1.07745 ps=6.86 w=6.53 l=0.62
X18 VDD1.t1 VP.t8 VTAIL.t5 w_n2110_n2274# sky130_fd_pr__pfet_01v8 ad=1.07745 pd=6.86 as=2.5467 ps=13.84 w=6.53 l=0.62
X19 VTAIL.t11 VN.t8 VDD2.t1 w_n2110_n2274# sky130_fd_pr__pfet_01v8 ad=1.07745 pd=6.86 as=1.07745 ps=6.86 w=6.53 l=0.62
X20 B.t5 B.t3 B.t4 w_n2110_n2274# sky130_fd_pr__pfet_01v8 ad=2.5467 pd=13.84 as=0 ps=0 w=6.53 l=0.62
X21 VDD2.t2 VN.t9 VTAIL.t10 w_n2110_n2274# sky130_fd_pr__pfet_01v8 ad=1.07745 pd=6.86 as=2.5467 ps=13.84 w=6.53 l=0.62
X22 VTAIL.t3 VP.t9 VDD1.t0 w_n2110_n2274# sky130_fd_pr__pfet_01v8 ad=1.07745 pd=6.86 as=1.07745 ps=6.86 w=6.53 l=0.62
X23 B.t2 B.t0 B.t1 w_n2110_n2274# sky130_fd_pr__pfet_01v8 ad=2.5467 pd=13.84 as=0 ps=0 w=6.53 l=0.62
R0 VN.n2 VN.t4 344.397
R1 VN.n10 VN.t2 344.397
R2 VN.n1 VN.t5 317.577
R3 VN.n4 VN.t6 317.577
R4 VN.n5 VN.t8 317.577
R5 VN.n6 VN.t9 317.577
R6 VN.n9 VN.t0 317.577
R7 VN.n12 VN.t7 317.577
R8 VN.n13 VN.t3 317.577
R9 VN.n14 VN.t1 317.577
R10 VN.n7 VN.n6 161.3
R11 VN.n15 VN.n14 161.3
R12 VN.n13 VN.n8 80.6037
R13 VN.n12 VN.n11 80.6037
R14 VN.n5 VN.n0 80.6037
R15 VN.n4 VN.n3 80.6037
R16 VN.n4 VN.n1 48.2005
R17 VN.n5 VN.n4 48.2005
R18 VN.n6 VN.n5 48.2005
R19 VN.n12 VN.n9 48.2005
R20 VN.n13 VN.n12 48.2005
R21 VN.n14 VN.n13 48.2005
R22 VN.n11 VN.n10 45.2318
R23 VN.n3 VN.n2 45.2318
R24 VN VN.n15 38.635
R25 VN.n10 VN.n9 13.3799
R26 VN.n2 VN.n1 13.3799
R27 VN.n11 VN.n8 0.380177
R28 VN.n3 VN.n0 0.380177
R29 VN.n15 VN.n8 0.285035
R30 VN.n7 VN.n0 0.285035
R31 VN VN.n7 0.0516364
R32 VDD2.n69 VDD2.n68 756.745
R33 VDD2.n32 VDD2.n31 756.745
R34 VDD2.n68 VDD2.n67 585
R35 VDD2.n39 VDD2.n38 585
R36 VDD2.n62 VDD2.n61 585
R37 VDD2.n60 VDD2.n59 585
R38 VDD2.n43 VDD2.n42 585
R39 VDD2.n54 VDD2.n53 585
R40 VDD2.n52 VDD2.n51 585
R41 VDD2.n47 VDD2.n46 585
R42 VDD2.n10 VDD2.n9 585
R43 VDD2.n15 VDD2.n14 585
R44 VDD2.n17 VDD2.n16 585
R45 VDD2.n6 VDD2.n5 585
R46 VDD2.n23 VDD2.n22 585
R47 VDD2.n25 VDD2.n24 585
R48 VDD2.n2 VDD2.n1 585
R49 VDD2.n31 VDD2.n30 585
R50 VDD2.n48 VDD2.t8 329.084
R51 VDD2.n11 VDD2.t3 329.084
R52 VDD2.n68 VDD2.n38 171.744
R53 VDD2.n61 VDD2.n38 171.744
R54 VDD2.n61 VDD2.n60 171.744
R55 VDD2.n60 VDD2.n42 171.744
R56 VDD2.n53 VDD2.n42 171.744
R57 VDD2.n53 VDD2.n52 171.744
R58 VDD2.n52 VDD2.n46 171.744
R59 VDD2.n15 VDD2.n9 171.744
R60 VDD2.n16 VDD2.n15 171.744
R61 VDD2.n16 VDD2.n5 171.744
R62 VDD2.n23 VDD2.n5 171.744
R63 VDD2.n24 VDD2.n23 171.744
R64 VDD2.n24 VDD2.n1 171.744
R65 VDD2.n31 VDD2.n1 171.744
R66 VDD2.n36 VDD2.n35 91.7111
R67 VDD2 VDD2.n73 91.7081
R68 VDD2.n72 VDD2.n71 91.1532
R69 VDD2.n34 VDD2.n33 91.1522
R70 VDD2.t8 VDD2.n46 85.8723
R71 VDD2.t3 VDD2.n9 85.8723
R72 VDD2.n34 VDD2.n32 52.5922
R73 VDD2.n70 VDD2.n69 51.7732
R74 VDD2.n70 VDD2.n36 33.2347
R75 VDD2.n67 VDD2.n37 12.8005
R76 VDD2.n30 VDD2.n0 12.8005
R77 VDD2.n66 VDD2.n39 12.0247
R78 VDD2.n29 VDD2.n2 12.0247
R79 VDD2.n63 VDD2.n62 11.249
R80 VDD2.n26 VDD2.n25 11.249
R81 VDD2.n48 VDD2.n47 10.7233
R82 VDD2.n11 VDD2.n10 10.7233
R83 VDD2.n59 VDD2.n41 10.4732
R84 VDD2.n22 VDD2.n4 10.4732
R85 VDD2.n58 VDD2.n43 9.69747
R86 VDD2.n21 VDD2.n6 9.69747
R87 VDD2.n65 VDD2.n37 9.45567
R88 VDD2.n28 VDD2.n0 9.45567
R89 VDD2.n45 VDD2.n44 9.3005
R90 VDD2.n56 VDD2.n55 9.3005
R91 VDD2.n58 VDD2.n57 9.3005
R92 VDD2.n41 VDD2.n40 9.3005
R93 VDD2.n64 VDD2.n63 9.3005
R94 VDD2.n66 VDD2.n65 9.3005
R95 VDD2.n50 VDD2.n49 9.3005
R96 VDD2.n13 VDD2.n12 9.3005
R97 VDD2.n8 VDD2.n7 9.3005
R98 VDD2.n19 VDD2.n18 9.3005
R99 VDD2.n21 VDD2.n20 9.3005
R100 VDD2.n4 VDD2.n3 9.3005
R101 VDD2.n27 VDD2.n26 9.3005
R102 VDD2.n29 VDD2.n28 9.3005
R103 VDD2.n55 VDD2.n54 8.92171
R104 VDD2.n18 VDD2.n17 8.92171
R105 VDD2.n51 VDD2.n45 8.14595
R106 VDD2.n14 VDD2.n8 8.14595
R107 VDD2.n50 VDD2.n47 7.3702
R108 VDD2.n13 VDD2.n10 7.3702
R109 VDD2.n51 VDD2.n50 5.81868
R110 VDD2.n14 VDD2.n13 5.81868
R111 VDD2.n54 VDD2.n45 5.04292
R112 VDD2.n17 VDD2.n8 5.04292
R113 VDD2.n73 VDD2.t7 4.9783
R114 VDD2.n73 VDD2.t5 4.9783
R115 VDD2.n71 VDD2.t4 4.9783
R116 VDD2.n71 VDD2.t0 4.9783
R117 VDD2.n35 VDD2.t1 4.9783
R118 VDD2.n35 VDD2.t2 4.9783
R119 VDD2.n33 VDD2.t9 4.9783
R120 VDD2.n33 VDD2.t6 4.9783
R121 VDD2.n55 VDD2.n43 4.26717
R122 VDD2.n18 VDD2.n6 4.26717
R123 VDD2.n59 VDD2.n58 3.49141
R124 VDD2.n22 VDD2.n21 3.49141
R125 VDD2.n62 VDD2.n41 2.71565
R126 VDD2.n25 VDD2.n4 2.71565
R127 VDD2.n49 VDD2.n48 2.41347
R128 VDD2.n12 VDD2.n11 2.41347
R129 VDD2.n63 VDD2.n39 1.93989
R130 VDD2.n26 VDD2.n2 1.93989
R131 VDD2.n67 VDD2.n66 1.16414
R132 VDD2.n30 VDD2.n29 1.16414
R133 VDD2.n72 VDD2.n70 0.819465
R134 VDD2.n69 VDD2.n37 0.388379
R135 VDD2.n32 VDD2.n0 0.388379
R136 VDD2 VDD2.n72 0.263431
R137 VDD2.n65 VDD2.n64 0.155672
R138 VDD2.n64 VDD2.n40 0.155672
R139 VDD2.n57 VDD2.n40 0.155672
R140 VDD2.n57 VDD2.n56 0.155672
R141 VDD2.n56 VDD2.n44 0.155672
R142 VDD2.n49 VDD2.n44 0.155672
R143 VDD2.n12 VDD2.n7 0.155672
R144 VDD2.n19 VDD2.n7 0.155672
R145 VDD2.n20 VDD2.n19 0.155672
R146 VDD2.n20 VDD2.n3 0.155672
R147 VDD2.n27 VDD2.n3 0.155672
R148 VDD2.n28 VDD2.n27 0.155672
R149 VDD2.n36 VDD2.n34 0.149895
R150 VTAIL.n148 VTAIL.n147 756.745
R151 VTAIL.n34 VTAIL.n33 756.745
R152 VTAIL.n114 VTAIL.n113 756.745
R153 VTAIL.n76 VTAIL.n75 756.745
R154 VTAIL.n126 VTAIL.n125 585
R155 VTAIL.n131 VTAIL.n130 585
R156 VTAIL.n133 VTAIL.n132 585
R157 VTAIL.n122 VTAIL.n121 585
R158 VTAIL.n139 VTAIL.n138 585
R159 VTAIL.n141 VTAIL.n140 585
R160 VTAIL.n118 VTAIL.n117 585
R161 VTAIL.n147 VTAIL.n146 585
R162 VTAIL.n12 VTAIL.n11 585
R163 VTAIL.n17 VTAIL.n16 585
R164 VTAIL.n19 VTAIL.n18 585
R165 VTAIL.n8 VTAIL.n7 585
R166 VTAIL.n25 VTAIL.n24 585
R167 VTAIL.n27 VTAIL.n26 585
R168 VTAIL.n4 VTAIL.n3 585
R169 VTAIL.n33 VTAIL.n32 585
R170 VTAIL.n113 VTAIL.n112 585
R171 VTAIL.n84 VTAIL.n83 585
R172 VTAIL.n107 VTAIL.n106 585
R173 VTAIL.n105 VTAIL.n104 585
R174 VTAIL.n88 VTAIL.n87 585
R175 VTAIL.n99 VTAIL.n98 585
R176 VTAIL.n97 VTAIL.n96 585
R177 VTAIL.n92 VTAIL.n91 585
R178 VTAIL.n75 VTAIL.n74 585
R179 VTAIL.n46 VTAIL.n45 585
R180 VTAIL.n69 VTAIL.n68 585
R181 VTAIL.n67 VTAIL.n66 585
R182 VTAIL.n50 VTAIL.n49 585
R183 VTAIL.n61 VTAIL.n60 585
R184 VTAIL.n59 VTAIL.n58 585
R185 VTAIL.n54 VTAIL.n53 585
R186 VTAIL.n127 VTAIL.t10 329.084
R187 VTAIL.n13 VTAIL.t2 329.084
R188 VTAIL.n93 VTAIL.t5 329.084
R189 VTAIL.n55 VTAIL.t17 329.084
R190 VTAIL.n131 VTAIL.n125 171.744
R191 VTAIL.n132 VTAIL.n131 171.744
R192 VTAIL.n132 VTAIL.n121 171.744
R193 VTAIL.n139 VTAIL.n121 171.744
R194 VTAIL.n140 VTAIL.n139 171.744
R195 VTAIL.n140 VTAIL.n117 171.744
R196 VTAIL.n147 VTAIL.n117 171.744
R197 VTAIL.n17 VTAIL.n11 171.744
R198 VTAIL.n18 VTAIL.n17 171.744
R199 VTAIL.n18 VTAIL.n7 171.744
R200 VTAIL.n25 VTAIL.n7 171.744
R201 VTAIL.n26 VTAIL.n25 171.744
R202 VTAIL.n26 VTAIL.n3 171.744
R203 VTAIL.n33 VTAIL.n3 171.744
R204 VTAIL.n113 VTAIL.n83 171.744
R205 VTAIL.n106 VTAIL.n83 171.744
R206 VTAIL.n106 VTAIL.n105 171.744
R207 VTAIL.n105 VTAIL.n87 171.744
R208 VTAIL.n98 VTAIL.n87 171.744
R209 VTAIL.n98 VTAIL.n97 171.744
R210 VTAIL.n97 VTAIL.n91 171.744
R211 VTAIL.n75 VTAIL.n45 171.744
R212 VTAIL.n68 VTAIL.n45 171.744
R213 VTAIL.n68 VTAIL.n67 171.744
R214 VTAIL.n67 VTAIL.n49 171.744
R215 VTAIL.n60 VTAIL.n49 171.744
R216 VTAIL.n60 VTAIL.n59 171.744
R217 VTAIL.n59 VTAIL.n53 171.744
R218 VTAIL.t10 VTAIL.n125 85.8723
R219 VTAIL.t2 VTAIL.n11 85.8723
R220 VTAIL.t5 VTAIL.n91 85.8723
R221 VTAIL.t17 VTAIL.n53 85.8723
R222 VTAIL.n81 VTAIL.n80 74.4744
R223 VTAIL.n79 VTAIL.n78 74.4744
R224 VTAIL.n43 VTAIL.n42 74.4744
R225 VTAIL.n41 VTAIL.n40 74.4744
R226 VTAIL.n151 VTAIL.n150 74.4734
R227 VTAIL.n1 VTAIL.n0 74.4734
R228 VTAIL.n37 VTAIL.n36 74.4734
R229 VTAIL.n39 VTAIL.n38 74.4734
R230 VTAIL.n149 VTAIL.n148 35.0944
R231 VTAIL.n35 VTAIL.n34 35.0944
R232 VTAIL.n115 VTAIL.n114 35.0944
R233 VTAIL.n77 VTAIL.n76 35.0944
R234 VTAIL.n41 VTAIL.n39 19.6341
R235 VTAIL.n149 VTAIL.n115 18.8152
R236 VTAIL.n146 VTAIL.n116 12.8005
R237 VTAIL.n32 VTAIL.n2 12.8005
R238 VTAIL.n112 VTAIL.n82 12.8005
R239 VTAIL.n74 VTAIL.n44 12.8005
R240 VTAIL.n145 VTAIL.n118 12.0247
R241 VTAIL.n31 VTAIL.n4 12.0247
R242 VTAIL.n111 VTAIL.n84 12.0247
R243 VTAIL.n73 VTAIL.n46 12.0247
R244 VTAIL.n142 VTAIL.n141 11.249
R245 VTAIL.n28 VTAIL.n27 11.249
R246 VTAIL.n108 VTAIL.n107 11.249
R247 VTAIL.n70 VTAIL.n69 11.249
R248 VTAIL.n127 VTAIL.n126 10.7233
R249 VTAIL.n13 VTAIL.n12 10.7233
R250 VTAIL.n93 VTAIL.n92 10.7233
R251 VTAIL.n55 VTAIL.n54 10.7233
R252 VTAIL.n138 VTAIL.n120 10.4732
R253 VTAIL.n24 VTAIL.n6 10.4732
R254 VTAIL.n104 VTAIL.n86 10.4732
R255 VTAIL.n66 VTAIL.n48 10.4732
R256 VTAIL.n137 VTAIL.n122 9.69747
R257 VTAIL.n23 VTAIL.n8 9.69747
R258 VTAIL.n103 VTAIL.n88 9.69747
R259 VTAIL.n65 VTAIL.n50 9.69747
R260 VTAIL.n144 VTAIL.n116 9.45567
R261 VTAIL.n30 VTAIL.n2 9.45567
R262 VTAIL.n110 VTAIL.n82 9.45567
R263 VTAIL.n72 VTAIL.n44 9.45567
R264 VTAIL.n129 VTAIL.n128 9.3005
R265 VTAIL.n124 VTAIL.n123 9.3005
R266 VTAIL.n135 VTAIL.n134 9.3005
R267 VTAIL.n137 VTAIL.n136 9.3005
R268 VTAIL.n120 VTAIL.n119 9.3005
R269 VTAIL.n143 VTAIL.n142 9.3005
R270 VTAIL.n145 VTAIL.n144 9.3005
R271 VTAIL.n15 VTAIL.n14 9.3005
R272 VTAIL.n10 VTAIL.n9 9.3005
R273 VTAIL.n21 VTAIL.n20 9.3005
R274 VTAIL.n23 VTAIL.n22 9.3005
R275 VTAIL.n6 VTAIL.n5 9.3005
R276 VTAIL.n29 VTAIL.n28 9.3005
R277 VTAIL.n31 VTAIL.n30 9.3005
R278 VTAIL.n111 VTAIL.n110 9.3005
R279 VTAIL.n109 VTAIL.n108 9.3005
R280 VTAIL.n86 VTAIL.n85 9.3005
R281 VTAIL.n103 VTAIL.n102 9.3005
R282 VTAIL.n101 VTAIL.n100 9.3005
R283 VTAIL.n90 VTAIL.n89 9.3005
R284 VTAIL.n95 VTAIL.n94 9.3005
R285 VTAIL.n52 VTAIL.n51 9.3005
R286 VTAIL.n63 VTAIL.n62 9.3005
R287 VTAIL.n65 VTAIL.n64 9.3005
R288 VTAIL.n48 VTAIL.n47 9.3005
R289 VTAIL.n71 VTAIL.n70 9.3005
R290 VTAIL.n73 VTAIL.n72 9.3005
R291 VTAIL.n57 VTAIL.n56 9.3005
R292 VTAIL.n134 VTAIL.n133 8.92171
R293 VTAIL.n20 VTAIL.n19 8.92171
R294 VTAIL.n100 VTAIL.n99 8.92171
R295 VTAIL.n62 VTAIL.n61 8.92171
R296 VTAIL.n130 VTAIL.n124 8.14595
R297 VTAIL.n16 VTAIL.n10 8.14595
R298 VTAIL.n96 VTAIL.n90 8.14595
R299 VTAIL.n58 VTAIL.n52 8.14595
R300 VTAIL.n129 VTAIL.n126 7.3702
R301 VTAIL.n15 VTAIL.n12 7.3702
R302 VTAIL.n95 VTAIL.n92 7.3702
R303 VTAIL.n57 VTAIL.n54 7.3702
R304 VTAIL.n130 VTAIL.n129 5.81868
R305 VTAIL.n16 VTAIL.n15 5.81868
R306 VTAIL.n96 VTAIL.n95 5.81868
R307 VTAIL.n58 VTAIL.n57 5.81868
R308 VTAIL.n133 VTAIL.n124 5.04292
R309 VTAIL.n19 VTAIL.n10 5.04292
R310 VTAIL.n99 VTAIL.n90 5.04292
R311 VTAIL.n61 VTAIL.n52 5.04292
R312 VTAIL.n150 VTAIL.t13 4.9783
R313 VTAIL.n150 VTAIL.t11 4.9783
R314 VTAIL.n0 VTAIL.t15 4.9783
R315 VTAIL.n0 VTAIL.t14 4.9783
R316 VTAIL.n36 VTAIL.t0 4.9783
R317 VTAIL.n36 VTAIL.t7 4.9783
R318 VTAIL.n38 VTAIL.t1 4.9783
R319 VTAIL.n38 VTAIL.t8 4.9783
R320 VTAIL.n80 VTAIL.t4 4.9783
R321 VTAIL.n80 VTAIL.t9 4.9783
R322 VTAIL.n78 VTAIL.t6 4.9783
R323 VTAIL.n78 VTAIL.t3 4.9783
R324 VTAIL.n42 VTAIL.t12 4.9783
R325 VTAIL.n42 VTAIL.t19 4.9783
R326 VTAIL.n40 VTAIL.t18 4.9783
R327 VTAIL.n40 VTAIL.t16 4.9783
R328 VTAIL.n134 VTAIL.n122 4.26717
R329 VTAIL.n20 VTAIL.n8 4.26717
R330 VTAIL.n100 VTAIL.n88 4.26717
R331 VTAIL.n62 VTAIL.n50 4.26717
R332 VTAIL.n138 VTAIL.n137 3.49141
R333 VTAIL.n24 VTAIL.n23 3.49141
R334 VTAIL.n104 VTAIL.n103 3.49141
R335 VTAIL.n66 VTAIL.n65 3.49141
R336 VTAIL.n141 VTAIL.n120 2.71565
R337 VTAIL.n27 VTAIL.n6 2.71565
R338 VTAIL.n107 VTAIL.n86 2.71565
R339 VTAIL.n69 VTAIL.n48 2.71565
R340 VTAIL.n56 VTAIL.n55 2.41347
R341 VTAIL.n128 VTAIL.n127 2.41347
R342 VTAIL.n14 VTAIL.n13 2.41347
R343 VTAIL.n94 VTAIL.n93 2.41347
R344 VTAIL.n142 VTAIL.n118 1.93989
R345 VTAIL.n28 VTAIL.n4 1.93989
R346 VTAIL.n108 VTAIL.n84 1.93989
R347 VTAIL.n70 VTAIL.n46 1.93989
R348 VTAIL.n146 VTAIL.n145 1.16414
R349 VTAIL.n32 VTAIL.n31 1.16414
R350 VTAIL.n112 VTAIL.n111 1.16414
R351 VTAIL.n74 VTAIL.n73 1.16414
R352 VTAIL.n79 VTAIL.n77 0.87981
R353 VTAIL.n35 VTAIL.n1 0.87981
R354 VTAIL.n43 VTAIL.n41 0.819465
R355 VTAIL.n77 VTAIL.n43 0.819465
R356 VTAIL.n81 VTAIL.n79 0.819465
R357 VTAIL.n115 VTAIL.n81 0.819465
R358 VTAIL.n39 VTAIL.n37 0.819465
R359 VTAIL.n37 VTAIL.n35 0.819465
R360 VTAIL.n151 VTAIL.n149 0.819465
R361 VTAIL VTAIL.n1 0.672914
R362 VTAIL.n148 VTAIL.n116 0.388379
R363 VTAIL.n34 VTAIL.n2 0.388379
R364 VTAIL.n114 VTAIL.n82 0.388379
R365 VTAIL.n76 VTAIL.n44 0.388379
R366 VTAIL.n128 VTAIL.n123 0.155672
R367 VTAIL.n135 VTAIL.n123 0.155672
R368 VTAIL.n136 VTAIL.n135 0.155672
R369 VTAIL.n136 VTAIL.n119 0.155672
R370 VTAIL.n143 VTAIL.n119 0.155672
R371 VTAIL.n144 VTAIL.n143 0.155672
R372 VTAIL.n14 VTAIL.n9 0.155672
R373 VTAIL.n21 VTAIL.n9 0.155672
R374 VTAIL.n22 VTAIL.n21 0.155672
R375 VTAIL.n22 VTAIL.n5 0.155672
R376 VTAIL.n29 VTAIL.n5 0.155672
R377 VTAIL.n30 VTAIL.n29 0.155672
R378 VTAIL.n110 VTAIL.n109 0.155672
R379 VTAIL.n109 VTAIL.n85 0.155672
R380 VTAIL.n102 VTAIL.n85 0.155672
R381 VTAIL.n102 VTAIL.n101 0.155672
R382 VTAIL.n101 VTAIL.n89 0.155672
R383 VTAIL.n94 VTAIL.n89 0.155672
R384 VTAIL.n72 VTAIL.n71 0.155672
R385 VTAIL.n71 VTAIL.n47 0.155672
R386 VTAIL.n64 VTAIL.n47 0.155672
R387 VTAIL.n64 VTAIL.n63 0.155672
R388 VTAIL.n63 VTAIL.n51 0.155672
R389 VTAIL.n56 VTAIL.n51 0.155672
R390 VTAIL VTAIL.n151 0.147052
R391 VP.n4 VP.t3 344.397
R392 VP.n10 VP.t6 317.577
R393 VP.n1 VP.t5 317.577
R394 VP.n14 VP.t4 317.577
R395 VP.n15 VP.t1 317.577
R396 VP.n16 VP.t0 317.577
R397 VP.n8 VP.t8 317.577
R398 VP.n7 VP.t2 317.577
R399 VP.n6 VP.t7 317.577
R400 VP.n5 VP.t9 317.577
R401 VP.n17 VP.n16 161.3
R402 VP.n9 VP.n8 161.3
R403 VP.n11 VP.n10 161.3
R404 VP.n6 VP.n3 80.6037
R405 VP.n7 VP.n2 80.6037
R406 VP.n15 VP.n0 80.6037
R407 VP.n14 VP.n13 80.6037
R408 VP.n12 VP.n1 80.6037
R409 VP.n10 VP.n1 48.2005
R410 VP.n14 VP.n1 48.2005
R411 VP.n15 VP.n14 48.2005
R412 VP.n16 VP.n15 48.2005
R413 VP.n8 VP.n7 48.2005
R414 VP.n7 VP.n6 48.2005
R415 VP.n6 VP.n5 48.2005
R416 VP.n4 VP.n3 45.2318
R417 VP.n11 VP.n9 38.2543
R418 VP.n5 VP.n4 13.3799
R419 VP.n3 VP.n2 0.380177
R420 VP.n13 VP.n12 0.380177
R421 VP.n13 VP.n0 0.380177
R422 VP.n9 VP.n2 0.285035
R423 VP.n12 VP.n11 0.285035
R424 VP.n17 VP.n0 0.285035
R425 VP VP.n17 0.0516364
R426 VDD1.n32 VDD1.n31 756.745
R427 VDD1.n67 VDD1.n66 756.745
R428 VDD1.n31 VDD1.n30 585
R429 VDD1.n2 VDD1.n1 585
R430 VDD1.n25 VDD1.n24 585
R431 VDD1.n23 VDD1.n22 585
R432 VDD1.n6 VDD1.n5 585
R433 VDD1.n17 VDD1.n16 585
R434 VDD1.n15 VDD1.n14 585
R435 VDD1.n10 VDD1.n9 585
R436 VDD1.n45 VDD1.n44 585
R437 VDD1.n50 VDD1.n49 585
R438 VDD1.n52 VDD1.n51 585
R439 VDD1.n41 VDD1.n40 585
R440 VDD1.n58 VDD1.n57 585
R441 VDD1.n60 VDD1.n59 585
R442 VDD1.n37 VDD1.n36 585
R443 VDD1.n66 VDD1.n65 585
R444 VDD1.n11 VDD1.t6 329.084
R445 VDD1.n46 VDD1.t3 329.084
R446 VDD1.n31 VDD1.n1 171.744
R447 VDD1.n24 VDD1.n1 171.744
R448 VDD1.n24 VDD1.n23 171.744
R449 VDD1.n23 VDD1.n5 171.744
R450 VDD1.n16 VDD1.n5 171.744
R451 VDD1.n16 VDD1.n15 171.744
R452 VDD1.n15 VDD1.n9 171.744
R453 VDD1.n50 VDD1.n44 171.744
R454 VDD1.n51 VDD1.n50 171.744
R455 VDD1.n51 VDD1.n40 171.744
R456 VDD1.n58 VDD1.n40 171.744
R457 VDD1.n59 VDD1.n58 171.744
R458 VDD1.n59 VDD1.n36 171.744
R459 VDD1.n66 VDD1.n36 171.744
R460 VDD1.n71 VDD1.n70 91.7111
R461 VDD1.n34 VDD1.n33 91.1532
R462 VDD1.n69 VDD1.n68 91.1522
R463 VDD1.n73 VDD1.n72 91.1521
R464 VDD1.t6 VDD1.n9 85.8723
R465 VDD1.t3 VDD1.n44 85.8723
R466 VDD1.n34 VDD1.n32 52.5922
R467 VDD1.n69 VDD1.n67 52.5922
R468 VDD1.n73 VDD1.n71 34.2272
R469 VDD1.n30 VDD1.n0 12.8005
R470 VDD1.n65 VDD1.n35 12.8005
R471 VDD1.n29 VDD1.n2 12.0247
R472 VDD1.n64 VDD1.n37 12.0247
R473 VDD1.n26 VDD1.n25 11.249
R474 VDD1.n61 VDD1.n60 11.249
R475 VDD1.n11 VDD1.n10 10.7233
R476 VDD1.n46 VDD1.n45 10.7233
R477 VDD1.n22 VDD1.n4 10.4732
R478 VDD1.n57 VDD1.n39 10.4732
R479 VDD1.n21 VDD1.n6 9.69747
R480 VDD1.n56 VDD1.n41 9.69747
R481 VDD1.n28 VDD1.n0 9.45567
R482 VDD1.n63 VDD1.n35 9.45567
R483 VDD1.n8 VDD1.n7 9.3005
R484 VDD1.n19 VDD1.n18 9.3005
R485 VDD1.n21 VDD1.n20 9.3005
R486 VDD1.n4 VDD1.n3 9.3005
R487 VDD1.n27 VDD1.n26 9.3005
R488 VDD1.n29 VDD1.n28 9.3005
R489 VDD1.n13 VDD1.n12 9.3005
R490 VDD1.n48 VDD1.n47 9.3005
R491 VDD1.n43 VDD1.n42 9.3005
R492 VDD1.n54 VDD1.n53 9.3005
R493 VDD1.n56 VDD1.n55 9.3005
R494 VDD1.n39 VDD1.n38 9.3005
R495 VDD1.n62 VDD1.n61 9.3005
R496 VDD1.n64 VDD1.n63 9.3005
R497 VDD1.n18 VDD1.n17 8.92171
R498 VDD1.n53 VDD1.n52 8.92171
R499 VDD1.n14 VDD1.n8 8.14595
R500 VDD1.n49 VDD1.n43 8.14595
R501 VDD1.n13 VDD1.n10 7.3702
R502 VDD1.n48 VDD1.n45 7.3702
R503 VDD1.n14 VDD1.n13 5.81868
R504 VDD1.n49 VDD1.n48 5.81868
R505 VDD1.n17 VDD1.n8 5.04292
R506 VDD1.n52 VDD1.n43 5.04292
R507 VDD1.n72 VDD1.t7 4.9783
R508 VDD1.n72 VDD1.t1 4.9783
R509 VDD1.n33 VDD1.t0 4.9783
R510 VDD1.n33 VDD1.t2 4.9783
R511 VDD1.n70 VDD1.t8 4.9783
R512 VDD1.n70 VDD1.t9 4.9783
R513 VDD1.n68 VDD1.t4 4.9783
R514 VDD1.n68 VDD1.t5 4.9783
R515 VDD1.n18 VDD1.n6 4.26717
R516 VDD1.n53 VDD1.n41 4.26717
R517 VDD1.n22 VDD1.n21 3.49141
R518 VDD1.n57 VDD1.n56 3.49141
R519 VDD1.n25 VDD1.n4 2.71565
R520 VDD1.n60 VDD1.n39 2.71565
R521 VDD1.n12 VDD1.n11 2.41347
R522 VDD1.n47 VDD1.n46 2.41347
R523 VDD1.n26 VDD1.n2 1.93989
R524 VDD1.n61 VDD1.n37 1.93989
R525 VDD1.n30 VDD1.n29 1.16414
R526 VDD1.n65 VDD1.n64 1.16414
R527 VDD1 VDD1.n73 0.556535
R528 VDD1.n32 VDD1.n0 0.388379
R529 VDD1.n67 VDD1.n35 0.388379
R530 VDD1 VDD1.n34 0.263431
R531 VDD1.n28 VDD1.n27 0.155672
R532 VDD1.n27 VDD1.n3 0.155672
R533 VDD1.n20 VDD1.n3 0.155672
R534 VDD1.n20 VDD1.n19 0.155672
R535 VDD1.n19 VDD1.n7 0.155672
R536 VDD1.n12 VDD1.n7 0.155672
R537 VDD1.n47 VDD1.n42 0.155672
R538 VDD1.n54 VDD1.n42 0.155672
R539 VDD1.n55 VDD1.n54 0.155672
R540 VDD1.n55 VDD1.n38 0.155672
R541 VDD1.n62 VDD1.n38 0.155672
R542 VDD1.n63 VDD1.n62 0.155672
R543 VDD1.n71 VDD1.n69 0.149895
R544 B.n328 B.n49 585
R545 B.n330 B.n329 585
R546 B.n331 B.n48 585
R547 B.n333 B.n332 585
R548 B.n334 B.n47 585
R549 B.n336 B.n335 585
R550 B.n337 B.n46 585
R551 B.n339 B.n338 585
R552 B.n340 B.n45 585
R553 B.n342 B.n341 585
R554 B.n343 B.n44 585
R555 B.n345 B.n344 585
R556 B.n346 B.n43 585
R557 B.n348 B.n347 585
R558 B.n349 B.n42 585
R559 B.n351 B.n350 585
R560 B.n352 B.n41 585
R561 B.n354 B.n353 585
R562 B.n355 B.n40 585
R563 B.n357 B.n356 585
R564 B.n358 B.n39 585
R565 B.n360 B.n359 585
R566 B.n361 B.n38 585
R567 B.n363 B.n362 585
R568 B.n364 B.n37 585
R569 B.n366 B.n365 585
R570 B.n368 B.n367 585
R571 B.n369 B.n33 585
R572 B.n371 B.n370 585
R573 B.n372 B.n32 585
R574 B.n374 B.n373 585
R575 B.n375 B.n31 585
R576 B.n377 B.n376 585
R577 B.n378 B.n30 585
R578 B.n380 B.n379 585
R579 B.n382 B.n27 585
R580 B.n384 B.n383 585
R581 B.n385 B.n26 585
R582 B.n387 B.n386 585
R583 B.n388 B.n25 585
R584 B.n390 B.n389 585
R585 B.n391 B.n24 585
R586 B.n393 B.n392 585
R587 B.n394 B.n23 585
R588 B.n396 B.n395 585
R589 B.n397 B.n22 585
R590 B.n399 B.n398 585
R591 B.n400 B.n21 585
R592 B.n402 B.n401 585
R593 B.n403 B.n20 585
R594 B.n405 B.n404 585
R595 B.n406 B.n19 585
R596 B.n408 B.n407 585
R597 B.n409 B.n18 585
R598 B.n411 B.n410 585
R599 B.n412 B.n17 585
R600 B.n414 B.n413 585
R601 B.n415 B.n16 585
R602 B.n417 B.n416 585
R603 B.n418 B.n15 585
R604 B.n420 B.n419 585
R605 B.n327 B.n326 585
R606 B.n325 B.n50 585
R607 B.n324 B.n323 585
R608 B.n322 B.n51 585
R609 B.n321 B.n320 585
R610 B.n319 B.n52 585
R611 B.n318 B.n317 585
R612 B.n316 B.n53 585
R613 B.n315 B.n314 585
R614 B.n313 B.n54 585
R615 B.n312 B.n311 585
R616 B.n310 B.n55 585
R617 B.n309 B.n308 585
R618 B.n307 B.n56 585
R619 B.n306 B.n305 585
R620 B.n304 B.n57 585
R621 B.n303 B.n302 585
R622 B.n301 B.n58 585
R623 B.n300 B.n299 585
R624 B.n298 B.n59 585
R625 B.n297 B.n296 585
R626 B.n295 B.n60 585
R627 B.n294 B.n293 585
R628 B.n292 B.n61 585
R629 B.n291 B.n290 585
R630 B.n289 B.n62 585
R631 B.n288 B.n287 585
R632 B.n286 B.n63 585
R633 B.n285 B.n284 585
R634 B.n283 B.n64 585
R635 B.n282 B.n281 585
R636 B.n280 B.n65 585
R637 B.n279 B.n278 585
R638 B.n277 B.n66 585
R639 B.n276 B.n275 585
R640 B.n274 B.n67 585
R641 B.n273 B.n272 585
R642 B.n271 B.n68 585
R643 B.n270 B.n269 585
R644 B.n268 B.n69 585
R645 B.n267 B.n266 585
R646 B.n265 B.n70 585
R647 B.n264 B.n263 585
R648 B.n262 B.n71 585
R649 B.n261 B.n260 585
R650 B.n259 B.n72 585
R651 B.n258 B.n257 585
R652 B.n256 B.n73 585
R653 B.n255 B.n254 585
R654 B.n253 B.n74 585
R655 B.n252 B.n251 585
R656 B.n159 B.n158 585
R657 B.n160 B.n109 585
R658 B.n162 B.n161 585
R659 B.n163 B.n108 585
R660 B.n165 B.n164 585
R661 B.n166 B.n107 585
R662 B.n168 B.n167 585
R663 B.n169 B.n106 585
R664 B.n171 B.n170 585
R665 B.n172 B.n105 585
R666 B.n174 B.n173 585
R667 B.n175 B.n104 585
R668 B.n177 B.n176 585
R669 B.n178 B.n103 585
R670 B.n180 B.n179 585
R671 B.n181 B.n102 585
R672 B.n183 B.n182 585
R673 B.n184 B.n101 585
R674 B.n186 B.n185 585
R675 B.n187 B.n100 585
R676 B.n189 B.n188 585
R677 B.n190 B.n99 585
R678 B.n192 B.n191 585
R679 B.n193 B.n98 585
R680 B.n195 B.n194 585
R681 B.n196 B.n95 585
R682 B.n199 B.n198 585
R683 B.n200 B.n94 585
R684 B.n202 B.n201 585
R685 B.n203 B.n93 585
R686 B.n205 B.n204 585
R687 B.n206 B.n92 585
R688 B.n208 B.n207 585
R689 B.n209 B.n91 585
R690 B.n211 B.n210 585
R691 B.n213 B.n212 585
R692 B.n214 B.n87 585
R693 B.n216 B.n215 585
R694 B.n217 B.n86 585
R695 B.n219 B.n218 585
R696 B.n220 B.n85 585
R697 B.n222 B.n221 585
R698 B.n223 B.n84 585
R699 B.n225 B.n224 585
R700 B.n226 B.n83 585
R701 B.n228 B.n227 585
R702 B.n229 B.n82 585
R703 B.n231 B.n230 585
R704 B.n232 B.n81 585
R705 B.n234 B.n233 585
R706 B.n235 B.n80 585
R707 B.n237 B.n236 585
R708 B.n238 B.n79 585
R709 B.n240 B.n239 585
R710 B.n241 B.n78 585
R711 B.n243 B.n242 585
R712 B.n244 B.n77 585
R713 B.n246 B.n245 585
R714 B.n247 B.n76 585
R715 B.n249 B.n248 585
R716 B.n250 B.n75 585
R717 B.n157 B.n110 585
R718 B.n156 B.n155 585
R719 B.n154 B.n111 585
R720 B.n153 B.n152 585
R721 B.n151 B.n112 585
R722 B.n150 B.n149 585
R723 B.n148 B.n113 585
R724 B.n147 B.n146 585
R725 B.n145 B.n114 585
R726 B.n144 B.n143 585
R727 B.n142 B.n115 585
R728 B.n141 B.n140 585
R729 B.n139 B.n116 585
R730 B.n138 B.n137 585
R731 B.n136 B.n117 585
R732 B.n135 B.n134 585
R733 B.n133 B.n118 585
R734 B.n132 B.n131 585
R735 B.n130 B.n119 585
R736 B.n129 B.n128 585
R737 B.n127 B.n120 585
R738 B.n126 B.n125 585
R739 B.n124 B.n121 585
R740 B.n123 B.n122 585
R741 B.n2 B.n0 585
R742 B.n457 B.n1 585
R743 B.n456 B.n455 585
R744 B.n454 B.n3 585
R745 B.n453 B.n452 585
R746 B.n451 B.n4 585
R747 B.n450 B.n449 585
R748 B.n448 B.n5 585
R749 B.n447 B.n446 585
R750 B.n445 B.n6 585
R751 B.n444 B.n443 585
R752 B.n442 B.n7 585
R753 B.n441 B.n440 585
R754 B.n439 B.n8 585
R755 B.n438 B.n437 585
R756 B.n436 B.n9 585
R757 B.n435 B.n434 585
R758 B.n433 B.n10 585
R759 B.n432 B.n431 585
R760 B.n430 B.n11 585
R761 B.n429 B.n428 585
R762 B.n427 B.n12 585
R763 B.n426 B.n425 585
R764 B.n424 B.n13 585
R765 B.n423 B.n422 585
R766 B.n421 B.n14 585
R767 B.n459 B.n458 585
R768 B.n88 B.t9 457.904
R769 B.n96 B.t6 457.904
R770 B.n28 B.t0 457.904
R771 B.n34 B.t3 457.904
R772 B.n158 B.n157 449.257
R773 B.n421 B.n420 449.257
R774 B.n252 B.n75 449.257
R775 B.n326 B.n49 449.257
R776 B.n88 B.t11 295.702
R777 B.n34 B.t4 295.702
R778 B.n96 B.t8 295.702
R779 B.n28 B.t1 295.702
R780 B.n89 B.t10 277.277
R781 B.n35 B.t5 277.277
R782 B.n97 B.t7 277.277
R783 B.n29 B.t2 277.277
R784 B.n157 B.n156 163.367
R785 B.n156 B.n111 163.367
R786 B.n152 B.n111 163.367
R787 B.n152 B.n151 163.367
R788 B.n151 B.n150 163.367
R789 B.n150 B.n113 163.367
R790 B.n146 B.n113 163.367
R791 B.n146 B.n145 163.367
R792 B.n145 B.n144 163.367
R793 B.n144 B.n115 163.367
R794 B.n140 B.n115 163.367
R795 B.n140 B.n139 163.367
R796 B.n139 B.n138 163.367
R797 B.n138 B.n117 163.367
R798 B.n134 B.n117 163.367
R799 B.n134 B.n133 163.367
R800 B.n133 B.n132 163.367
R801 B.n132 B.n119 163.367
R802 B.n128 B.n119 163.367
R803 B.n128 B.n127 163.367
R804 B.n127 B.n126 163.367
R805 B.n126 B.n121 163.367
R806 B.n122 B.n121 163.367
R807 B.n122 B.n2 163.367
R808 B.n458 B.n2 163.367
R809 B.n458 B.n457 163.367
R810 B.n457 B.n456 163.367
R811 B.n456 B.n3 163.367
R812 B.n452 B.n3 163.367
R813 B.n452 B.n451 163.367
R814 B.n451 B.n450 163.367
R815 B.n450 B.n5 163.367
R816 B.n446 B.n5 163.367
R817 B.n446 B.n445 163.367
R818 B.n445 B.n444 163.367
R819 B.n444 B.n7 163.367
R820 B.n440 B.n7 163.367
R821 B.n440 B.n439 163.367
R822 B.n439 B.n438 163.367
R823 B.n438 B.n9 163.367
R824 B.n434 B.n9 163.367
R825 B.n434 B.n433 163.367
R826 B.n433 B.n432 163.367
R827 B.n432 B.n11 163.367
R828 B.n428 B.n11 163.367
R829 B.n428 B.n427 163.367
R830 B.n427 B.n426 163.367
R831 B.n426 B.n13 163.367
R832 B.n422 B.n13 163.367
R833 B.n422 B.n421 163.367
R834 B.n158 B.n109 163.367
R835 B.n162 B.n109 163.367
R836 B.n163 B.n162 163.367
R837 B.n164 B.n163 163.367
R838 B.n164 B.n107 163.367
R839 B.n168 B.n107 163.367
R840 B.n169 B.n168 163.367
R841 B.n170 B.n169 163.367
R842 B.n170 B.n105 163.367
R843 B.n174 B.n105 163.367
R844 B.n175 B.n174 163.367
R845 B.n176 B.n175 163.367
R846 B.n176 B.n103 163.367
R847 B.n180 B.n103 163.367
R848 B.n181 B.n180 163.367
R849 B.n182 B.n181 163.367
R850 B.n182 B.n101 163.367
R851 B.n186 B.n101 163.367
R852 B.n187 B.n186 163.367
R853 B.n188 B.n187 163.367
R854 B.n188 B.n99 163.367
R855 B.n192 B.n99 163.367
R856 B.n193 B.n192 163.367
R857 B.n194 B.n193 163.367
R858 B.n194 B.n95 163.367
R859 B.n199 B.n95 163.367
R860 B.n200 B.n199 163.367
R861 B.n201 B.n200 163.367
R862 B.n201 B.n93 163.367
R863 B.n205 B.n93 163.367
R864 B.n206 B.n205 163.367
R865 B.n207 B.n206 163.367
R866 B.n207 B.n91 163.367
R867 B.n211 B.n91 163.367
R868 B.n212 B.n211 163.367
R869 B.n212 B.n87 163.367
R870 B.n216 B.n87 163.367
R871 B.n217 B.n216 163.367
R872 B.n218 B.n217 163.367
R873 B.n218 B.n85 163.367
R874 B.n222 B.n85 163.367
R875 B.n223 B.n222 163.367
R876 B.n224 B.n223 163.367
R877 B.n224 B.n83 163.367
R878 B.n228 B.n83 163.367
R879 B.n229 B.n228 163.367
R880 B.n230 B.n229 163.367
R881 B.n230 B.n81 163.367
R882 B.n234 B.n81 163.367
R883 B.n235 B.n234 163.367
R884 B.n236 B.n235 163.367
R885 B.n236 B.n79 163.367
R886 B.n240 B.n79 163.367
R887 B.n241 B.n240 163.367
R888 B.n242 B.n241 163.367
R889 B.n242 B.n77 163.367
R890 B.n246 B.n77 163.367
R891 B.n247 B.n246 163.367
R892 B.n248 B.n247 163.367
R893 B.n248 B.n75 163.367
R894 B.n253 B.n252 163.367
R895 B.n254 B.n253 163.367
R896 B.n254 B.n73 163.367
R897 B.n258 B.n73 163.367
R898 B.n259 B.n258 163.367
R899 B.n260 B.n259 163.367
R900 B.n260 B.n71 163.367
R901 B.n264 B.n71 163.367
R902 B.n265 B.n264 163.367
R903 B.n266 B.n265 163.367
R904 B.n266 B.n69 163.367
R905 B.n270 B.n69 163.367
R906 B.n271 B.n270 163.367
R907 B.n272 B.n271 163.367
R908 B.n272 B.n67 163.367
R909 B.n276 B.n67 163.367
R910 B.n277 B.n276 163.367
R911 B.n278 B.n277 163.367
R912 B.n278 B.n65 163.367
R913 B.n282 B.n65 163.367
R914 B.n283 B.n282 163.367
R915 B.n284 B.n283 163.367
R916 B.n284 B.n63 163.367
R917 B.n288 B.n63 163.367
R918 B.n289 B.n288 163.367
R919 B.n290 B.n289 163.367
R920 B.n290 B.n61 163.367
R921 B.n294 B.n61 163.367
R922 B.n295 B.n294 163.367
R923 B.n296 B.n295 163.367
R924 B.n296 B.n59 163.367
R925 B.n300 B.n59 163.367
R926 B.n301 B.n300 163.367
R927 B.n302 B.n301 163.367
R928 B.n302 B.n57 163.367
R929 B.n306 B.n57 163.367
R930 B.n307 B.n306 163.367
R931 B.n308 B.n307 163.367
R932 B.n308 B.n55 163.367
R933 B.n312 B.n55 163.367
R934 B.n313 B.n312 163.367
R935 B.n314 B.n313 163.367
R936 B.n314 B.n53 163.367
R937 B.n318 B.n53 163.367
R938 B.n319 B.n318 163.367
R939 B.n320 B.n319 163.367
R940 B.n320 B.n51 163.367
R941 B.n324 B.n51 163.367
R942 B.n325 B.n324 163.367
R943 B.n326 B.n325 163.367
R944 B.n420 B.n15 163.367
R945 B.n416 B.n15 163.367
R946 B.n416 B.n415 163.367
R947 B.n415 B.n414 163.367
R948 B.n414 B.n17 163.367
R949 B.n410 B.n17 163.367
R950 B.n410 B.n409 163.367
R951 B.n409 B.n408 163.367
R952 B.n408 B.n19 163.367
R953 B.n404 B.n19 163.367
R954 B.n404 B.n403 163.367
R955 B.n403 B.n402 163.367
R956 B.n402 B.n21 163.367
R957 B.n398 B.n21 163.367
R958 B.n398 B.n397 163.367
R959 B.n397 B.n396 163.367
R960 B.n396 B.n23 163.367
R961 B.n392 B.n23 163.367
R962 B.n392 B.n391 163.367
R963 B.n391 B.n390 163.367
R964 B.n390 B.n25 163.367
R965 B.n386 B.n25 163.367
R966 B.n386 B.n385 163.367
R967 B.n385 B.n384 163.367
R968 B.n384 B.n27 163.367
R969 B.n379 B.n27 163.367
R970 B.n379 B.n378 163.367
R971 B.n378 B.n377 163.367
R972 B.n377 B.n31 163.367
R973 B.n373 B.n31 163.367
R974 B.n373 B.n372 163.367
R975 B.n372 B.n371 163.367
R976 B.n371 B.n33 163.367
R977 B.n367 B.n33 163.367
R978 B.n367 B.n366 163.367
R979 B.n366 B.n37 163.367
R980 B.n362 B.n37 163.367
R981 B.n362 B.n361 163.367
R982 B.n361 B.n360 163.367
R983 B.n360 B.n39 163.367
R984 B.n356 B.n39 163.367
R985 B.n356 B.n355 163.367
R986 B.n355 B.n354 163.367
R987 B.n354 B.n41 163.367
R988 B.n350 B.n41 163.367
R989 B.n350 B.n349 163.367
R990 B.n349 B.n348 163.367
R991 B.n348 B.n43 163.367
R992 B.n344 B.n43 163.367
R993 B.n344 B.n343 163.367
R994 B.n343 B.n342 163.367
R995 B.n342 B.n45 163.367
R996 B.n338 B.n45 163.367
R997 B.n338 B.n337 163.367
R998 B.n337 B.n336 163.367
R999 B.n336 B.n47 163.367
R1000 B.n332 B.n47 163.367
R1001 B.n332 B.n331 163.367
R1002 B.n331 B.n330 163.367
R1003 B.n330 B.n49 163.367
R1004 B.n90 B.n89 59.5399
R1005 B.n197 B.n97 59.5399
R1006 B.n381 B.n29 59.5399
R1007 B.n36 B.n35 59.5399
R1008 B.n419 B.n14 29.1907
R1009 B.n328 B.n327 29.1907
R1010 B.n251 B.n250 29.1907
R1011 B.n159 B.n110 29.1907
R1012 B.n89 B.n88 18.4247
R1013 B.n97 B.n96 18.4247
R1014 B.n29 B.n28 18.4247
R1015 B.n35 B.n34 18.4247
R1016 B B.n459 18.0485
R1017 B.n419 B.n418 10.6151
R1018 B.n418 B.n417 10.6151
R1019 B.n417 B.n16 10.6151
R1020 B.n413 B.n16 10.6151
R1021 B.n413 B.n412 10.6151
R1022 B.n412 B.n411 10.6151
R1023 B.n411 B.n18 10.6151
R1024 B.n407 B.n18 10.6151
R1025 B.n407 B.n406 10.6151
R1026 B.n406 B.n405 10.6151
R1027 B.n405 B.n20 10.6151
R1028 B.n401 B.n20 10.6151
R1029 B.n401 B.n400 10.6151
R1030 B.n400 B.n399 10.6151
R1031 B.n399 B.n22 10.6151
R1032 B.n395 B.n22 10.6151
R1033 B.n395 B.n394 10.6151
R1034 B.n394 B.n393 10.6151
R1035 B.n393 B.n24 10.6151
R1036 B.n389 B.n24 10.6151
R1037 B.n389 B.n388 10.6151
R1038 B.n388 B.n387 10.6151
R1039 B.n387 B.n26 10.6151
R1040 B.n383 B.n26 10.6151
R1041 B.n383 B.n382 10.6151
R1042 B.n380 B.n30 10.6151
R1043 B.n376 B.n30 10.6151
R1044 B.n376 B.n375 10.6151
R1045 B.n375 B.n374 10.6151
R1046 B.n374 B.n32 10.6151
R1047 B.n370 B.n32 10.6151
R1048 B.n370 B.n369 10.6151
R1049 B.n369 B.n368 10.6151
R1050 B.n365 B.n364 10.6151
R1051 B.n364 B.n363 10.6151
R1052 B.n363 B.n38 10.6151
R1053 B.n359 B.n38 10.6151
R1054 B.n359 B.n358 10.6151
R1055 B.n358 B.n357 10.6151
R1056 B.n357 B.n40 10.6151
R1057 B.n353 B.n40 10.6151
R1058 B.n353 B.n352 10.6151
R1059 B.n352 B.n351 10.6151
R1060 B.n351 B.n42 10.6151
R1061 B.n347 B.n42 10.6151
R1062 B.n347 B.n346 10.6151
R1063 B.n346 B.n345 10.6151
R1064 B.n345 B.n44 10.6151
R1065 B.n341 B.n44 10.6151
R1066 B.n341 B.n340 10.6151
R1067 B.n340 B.n339 10.6151
R1068 B.n339 B.n46 10.6151
R1069 B.n335 B.n46 10.6151
R1070 B.n335 B.n334 10.6151
R1071 B.n334 B.n333 10.6151
R1072 B.n333 B.n48 10.6151
R1073 B.n329 B.n48 10.6151
R1074 B.n329 B.n328 10.6151
R1075 B.n251 B.n74 10.6151
R1076 B.n255 B.n74 10.6151
R1077 B.n256 B.n255 10.6151
R1078 B.n257 B.n256 10.6151
R1079 B.n257 B.n72 10.6151
R1080 B.n261 B.n72 10.6151
R1081 B.n262 B.n261 10.6151
R1082 B.n263 B.n262 10.6151
R1083 B.n263 B.n70 10.6151
R1084 B.n267 B.n70 10.6151
R1085 B.n268 B.n267 10.6151
R1086 B.n269 B.n268 10.6151
R1087 B.n269 B.n68 10.6151
R1088 B.n273 B.n68 10.6151
R1089 B.n274 B.n273 10.6151
R1090 B.n275 B.n274 10.6151
R1091 B.n275 B.n66 10.6151
R1092 B.n279 B.n66 10.6151
R1093 B.n280 B.n279 10.6151
R1094 B.n281 B.n280 10.6151
R1095 B.n281 B.n64 10.6151
R1096 B.n285 B.n64 10.6151
R1097 B.n286 B.n285 10.6151
R1098 B.n287 B.n286 10.6151
R1099 B.n287 B.n62 10.6151
R1100 B.n291 B.n62 10.6151
R1101 B.n292 B.n291 10.6151
R1102 B.n293 B.n292 10.6151
R1103 B.n293 B.n60 10.6151
R1104 B.n297 B.n60 10.6151
R1105 B.n298 B.n297 10.6151
R1106 B.n299 B.n298 10.6151
R1107 B.n299 B.n58 10.6151
R1108 B.n303 B.n58 10.6151
R1109 B.n304 B.n303 10.6151
R1110 B.n305 B.n304 10.6151
R1111 B.n305 B.n56 10.6151
R1112 B.n309 B.n56 10.6151
R1113 B.n310 B.n309 10.6151
R1114 B.n311 B.n310 10.6151
R1115 B.n311 B.n54 10.6151
R1116 B.n315 B.n54 10.6151
R1117 B.n316 B.n315 10.6151
R1118 B.n317 B.n316 10.6151
R1119 B.n317 B.n52 10.6151
R1120 B.n321 B.n52 10.6151
R1121 B.n322 B.n321 10.6151
R1122 B.n323 B.n322 10.6151
R1123 B.n323 B.n50 10.6151
R1124 B.n327 B.n50 10.6151
R1125 B.n160 B.n159 10.6151
R1126 B.n161 B.n160 10.6151
R1127 B.n161 B.n108 10.6151
R1128 B.n165 B.n108 10.6151
R1129 B.n166 B.n165 10.6151
R1130 B.n167 B.n166 10.6151
R1131 B.n167 B.n106 10.6151
R1132 B.n171 B.n106 10.6151
R1133 B.n172 B.n171 10.6151
R1134 B.n173 B.n172 10.6151
R1135 B.n173 B.n104 10.6151
R1136 B.n177 B.n104 10.6151
R1137 B.n178 B.n177 10.6151
R1138 B.n179 B.n178 10.6151
R1139 B.n179 B.n102 10.6151
R1140 B.n183 B.n102 10.6151
R1141 B.n184 B.n183 10.6151
R1142 B.n185 B.n184 10.6151
R1143 B.n185 B.n100 10.6151
R1144 B.n189 B.n100 10.6151
R1145 B.n190 B.n189 10.6151
R1146 B.n191 B.n190 10.6151
R1147 B.n191 B.n98 10.6151
R1148 B.n195 B.n98 10.6151
R1149 B.n196 B.n195 10.6151
R1150 B.n198 B.n94 10.6151
R1151 B.n202 B.n94 10.6151
R1152 B.n203 B.n202 10.6151
R1153 B.n204 B.n203 10.6151
R1154 B.n204 B.n92 10.6151
R1155 B.n208 B.n92 10.6151
R1156 B.n209 B.n208 10.6151
R1157 B.n210 B.n209 10.6151
R1158 B.n214 B.n213 10.6151
R1159 B.n215 B.n214 10.6151
R1160 B.n215 B.n86 10.6151
R1161 B.n219 B.n86 10.6151
R1162 B.n220 B.n219 10.6151
R1163 B.n221 B.n220 10.6151
R1164 B.n221 B.n84 10.6151
R1165 B.n225 B.n84 10.6151
R1166 B.n226 B.n225 10.6151
R1167 B.n227 B.n226 10.6151
R1168 B.n227 B.n82 10.6151
R1169 B.n231 B.n82 10.6151
R1170 B.n232 B.n231 10.6151
R1171 B.n233 B.n232 10.6151
R1172 B.n233 B.n80 10.6151
R1173 B.n237 B.n80 10.6151
R1174 B.n238 B.n237 10.6151
R1175 B.n239 B.n238 10.6151
R1176 B.n239 B.n78 10.6151
R1177 B.n243 B.n78 10.6151
R1178 B.n244 B.n243 10.6151
R1179 B.n245 B.n244 10.6151
R1180 B.n245 B.n76 10.6151
R1181 B.n249 B.n76 10.6151
R1182 B.n250 B.n249 10.6151
R1183 B.n155 B.n110 10.6151
R1184 B.n155 B.n154 10.6151
R1185 B.n154 B.n153 10.6151
R1186 B.n153 B.n112 10.6151
R1187 B.n149 B.n112 10.6151
R1188 B.n149 B.n148 10.6151
R1189 B.n148 B.n147 10.6151
R1190 B.n147 B.n114 10.6151
R1191 B.n143 B.n114 10.6151
R1192 B.n143 B.n142 10.6151
R1193 B.n142 B.n141 10.6151
R1194 B.n141 B.n116 10.6151
R1195 B.n137 B.n116 10.6151
R1196 B.n137 B.n136 10.6151
R1197 B.n136 B.n135 10.6151
R1198 B.n135 B.n118 10.6151
R1199 B.n131 B.n118 10.6151
R1200 B.n131 B.n130 10.6151
R1201 B.n130 B.n129 10.6151
R1202 B.n129 B.n120 10.6151
R1203 B.n125 B.n120 10.6151
R1204 B.n125 B.n124 10.6151
R1205 B.n124 B.n123 10.6151
R1206 B.n123 B.n0 10.6151
R1207 B.n455 B.n1 10.6151
R1208 B.n455 B.n454 10.6151
R1209 B.n454 B.n453 10.6151
R1210 B.n453 B.n4 10.6151
R1211 B.n449 B.n4 10.6151
R1212 B.n449 B.n448 10.6151
R1213 B.n448 B.n447 10.6151
R1214 B.n447 B.n6 10.6151
R1215 B.n443 B.n6 10.6151
R1216 B.n443 B.n442 10.6151
R1217 B.n442 B.n441 10.6151
R1218 B.n441 B.n8 10.6151
R1219 B.n437 B.n8 10.6151
R1220 B.n437 B.n436 10.6151
R1221 B.n436 B.n435 10.6151
R1222 B.n435 B.n10 10.6151
R1223 B.n431 B.n10 10.6151
R1224 B.n431 B.n430 10.6151
R1225 B.n430 B.n429 10.6151
R1226 B.n429 B.n12 10.6151
R1227 B.n425 B.n12 10.6151
R1228 B.n425 B.n424 10.6151
R1229 B.n424 B.n423 10.6151
R1230 B.n423 B.n14 10.6151
R1231 B.n381 B.n380 6.5566
R1232 B.n368 B.n36 6.5566
R1233 B.n198 B.n197 6.5566
R1234 B.n210 B.n90 6.5566
R1235 B.n382 B.n381 4.05904
R1236 B.n365 B.n36 4.05904
R1237 B.n197 B.n196 4.05904
R1238 B.n213 B.n90 4.05904
R1239 B.n459 B.n0 2.81026
R1240 B.n459 B.n1 2.81026
C0 VP VDD2 0.330679f
C1 B VDD2 1.31418f
C2 VTAIL VDD2 9.30445f
C3 VDD2 VN 3.59792f
C4 VDD1 VP 3.7768f
C5 VDD1 B 1.27296f
C6 VDD1 VTAIL 9.267941f
C7 VDD1 VN 0.148961f
C8 VDD1 VDD2 0.921889f
C9 w_n2110_n2274# VP 4.06871f
C10 w_n2110_n2274# B 5.68856f
C11 w_n2110_n2274# VTAIL 2.16948f
C12 w_n2110_n2274# VN 3.80011f
C13 w_n2110_n2274# VDD2 1.64326f
C14 w_n2110_n2274# VDD1 1.60275f
C15 B VP 1.15334f
C16 VTAIL VP 3.68322f
C17 B VTAIL 1.71624f
C18 VP VN 4.46546f
C19 B VN 0.712591f
C20 VTAIL VN 3.66883f
C21 VDD2 VSUBS 1.144701f
C22 VDD1 VSUBS 0.951212f
C23 VTAIL VSUBS 0.441365f
C24 VN VSUBS 4.41441f
C25 VP VSUBS 1.44448f
C26 B VSUBS 2.44722f
C27 w_n2110_n2274# VSUBS 59.780502f
C28 B.n0 VSUBS 0.004061f
C29 B.n1 VSUBS 0.004061f
C30 B.n2 VSUBS 0.006422f
C31 B.n3 VSUBS 0.006422f
C32 B.n4 VSUBS 0.006422f
C33 B.n5 VSUBS 0.006422f
C34 B.n6 VSUBS 0.006422f
C35 B.n7 VSUBS 0.006422f
C36 B.n8 VSUBS 0.006422f
C37 B.n9 VSUBS 0.006422f
C38 B.n10 VSUBS 0.006422f
C39 B.n11 VSUBS 0.006422f
C40 B.n12 VSUBS 0.006422f
C41 B.n13 VSUBS 0.006422f
C42 B.n14 VSUBS 0.013532f
C43 B.n15 VSUBS 0.006422f
C44 B.n16 VSUBS 0.006422f
C45 B.n17 VSUBS 0.006422f
C46 B.n18 VSUBS 0.006422f
C47 B.n19 VSUBS 0.006422f
C48 B.n20 VSUBS 0.006422f
C49 B.n21 VSUBS 0.006422f
C50 B.n22 VSUBS 0.006422f
C51 B.n23 VSUBS 0.006422f
C52 B.n24 VSUBS 0.006422f
C53 B.n25 VSUBS 0.006422f
C54 B.n26 VSUBS 0.006422f
C55 B.n27 VSUBS 0.006422f
C56 B.t2 VSUBS 0.09048f
C57 B.t1 VSUBS 0.098957f
C58 B.t0 VSUBS 0.15829f
C59 B.n28 VSUBS 0.168028f
C60 B.n29 VSUBS 0.1452f
C61 B.n30 VSUBS 0.006422f
C62 B.n31 VSUBS 0.006422f
C63 B.n32 VSUBS 0.006422f
C64 B.n33 VSUBS 0.006422f
C65 B.t5 VSUBS 0.090482f
C66 B.t4 VSUBS 0.098958f
C67 B.t3 VSUBS 0.15829f
C68 B.n34 VSUBS 0.168026f
C69 B.n35 VSUBS 0.145198f
C70 B.n36 VSUBS 0.014879f
C71 B.n37 VSUBS 0.006422f
C72 B.n38 VSUBS 0.006422f
C73 B.n39 VSUBS 0.006422f
C74 B.n40 VSUBS 0.006422f
C75 B.n41 VSUBS 0.006422f
C76 B.n42 VSUBS 0.006422f
C77 B.n43 VSUBS 0.006422f
C78 B.n44 VSUBS 0.006422f
C79 B.n45 VSUBS 0.006422f
C80 B.n46 VSUBS 0.006422f
C81 B.n47 VSUBS 0.006422f
C82 B.n48 VSUBS 0.006422f
C83 B.n49 VSUBS 0.014423f
C84 B.n50 VSUBS 0.006422f
C85 B.n51 VSUBS 0.006422f
C86 B.n52 VSUBS 0.006422f
C87 B.n53 VSUBS 0.006422f
C88 B.n54 VSUBS 0.006422f
C89 B.n55 VSUBS 0.006422f
C90 B.n56 VSUBS 0.006422f
C91 B.n57 VSUBS 0.006422f
C92 B.n58 VSUBS 0.006422f
C93 B.n59 VSUBS 0.006422f
C94 B.n60 VSUBS 0.006422f
C95 B.n61 VSUBS 0.006422f
C96 B.n62 VSUBS 0.006422f
C97 B.n63 VSUBS 0.006422f
C98 B.n64 VSUBS 0.006422f
C99 B.n65 VSUBS 0.006422f
C100 B.n66 VSUBS 0.006422f
C101 B.n67 VSUBS 0.006422f
C102 B.n68 VSUBS 0.006422f
C103 B.n69 VSUBS 0.006422f
C104 B.n70 VSUBS 0.006422f
C105 B.n71 VSUBS 0.006422f
C106 B.n72 VSUBS 0.006422f
C107 B.n73 VSUBS 0.006422f
C108 B.n74 VSUBS 0.006422f
C109 B.n75 VSUBS 0.014423f
C110 B.n76 VSUBS 0.006422f
C111 B.n77 VSUBS 0.006422f
C112 B.n78 VSUBS 0.006422f
C113 B.n79 VSUBS 0.006422f
C114 B.n80 VSUBS 0.006422f
C115 B.n81 VSUBS 0.006422f
C116 B.n82 VSUBS 0.006422f
C117 B.n83 VSUBS 0.006422f
C118 B.n84 VSUBS 0.006422f
C119 B.n85 VSUBS 0.006422f
C120 B.n86 VSUBS 0.006422f
C121 B.n87 VSUBS 0.006422f
C122 B.t10 VSUBS 0.090482f
C123 B.t11 VSUBS 0.098958f
C124 B.t9 VSUBS 0.15829f
C125 B.n88 VSUBS 0.168026f
C126 B.n89 VSUBS 0.145198f
C127 B.n90 VSUBS 0.014879f
C128 B.n91 VSUBS 0.006422f
C129 B.n92 VSUBS 0.006422f
C130 B.n93 VSUBS 0.006422f
C131 B.n94 VSUBS 0.006422f
C132 B.n95 VSUBS 0.006422f
C133 B.t7 VSUBS 0.09048f
C134 B.t8 VSUBS 0.098957f
C135 B.t6 VSUBS 0.15829f
C136 B.n96 VSUBS 0.168028f
C137 B.n97 VSUBS 0.1452f
C138 B.n98 VSUBS 0.006422f
C139 B.n99 VSUBS 0.006422f
C140 B.n100 VSUBS 0.006422f
C141 B.n101 VSUBS 0.006422f
C142 B.n102 VSUBS 0.006422f
C143 B.n103 VSUBS 0.006422f
C144 B.n104 VSUBS 0.006422f
C145 B.n105 VSUBS 0.006422f
C146 B.n106 VSUBS 0.006422f
C147 B.n107 VSUBS 0.006422f
C148 B.n108 VSUBS 0.006422f
C149 B.n109 VSUBS 0.006422f
C150 B.n110 VSUBS 0.013532f
C151 B.n111 VSUBS 0.006422f
C152 B.n112 VSUBS 0.006422f
C153 B.n113 VSUBS 0.006422f
C154 B.n114 VSUBS 0.006422f
C155 B.n115 VSUBS 0.006422f
C156 B.n116 VSUBS 0.006422f
C157 B.n117 VSUBS 0.006422f
C158 B.n118 VSUBS 0.006422f
C159 B.n119 VSUBS 0.006422f
C160 B.n120 VSUBS 0.006422f
C161 B.n121 VSUBS 0.006422f
C162 B.n122 VSUBS 0.006422f
C163 B.n123 VSUBS 0.006422f
C164 B.n124 VSUBS 0.006422f
C165 B.n125 VSUBS 0.006422f
C166 B.n126 VSUBS 0.006422f
C167 B.n127 VSUBS 0.006422f
C168 B.n128 VSUBS 0.006422f
C169 B.n129 VSUBS 0.006422f
C170 B.n130 VSUBS 0.006422f
C171 B.n131 VSUBS 0.006422f
C172 B.n132 VSUBS 0.006422f
C173 B.n133 VSUBS 0.006422f
C174 B.n134 VSUBS 0.006422f
C175 B.n135 VSUBS 0.006422f
C176 B.n136 VSUBS 0.006422f
C177 B.n137 VSUBS 0.006422f
C178 B.n138 VSUBS 0.006422f
C179 B.n139 VSUBS 0.006422f
C180 B.n140 VSUBS 0.006422f
C181 B.n141 VSUBS 0.006422f
C182 B.n142 VSUBS 0.006422f
C183 B.n143 VSUBS 0.006422f
C184 B.n144 VSUBS 0.006422f
C185 B.n145 VSUBS 0.006422f
C186 B.n146 VSUBS 0.006422f
C187 B.n147 VSUBS 0.006422f
C188 B.n148 VSUBS 0.006422f
C189 B.n149 VSUBS 0.006422f
C190 B.n150 VSUBS 0.006422f
C191 B.n151 VSUBS 0.006422f
C192 B.n152 VSUBS 0.006422f
C193 B.n153 VSUBS 0.006422f
C194 B.n154 VSUBS 0.006422f
C195 B.n155 VSUBS 0.006422f
C196 B.n156 VSUBS 0.006422f
C197 B.n157 VSUBS 0.013532f
C198 B.n158 VSUBS 0.014423f
C199 B.n159 VSUBS 0.014423f
C200 B.n160 VSUBS 0.006422f
C201 B.n161 VSUBS 0.006422f
C202 B.n162 VSUBS 0.006422f
C203 B.n163 VSUBS 0.006422f
C204 B.n164 VSUBS 0.006422f
C205 B.n165 VSUBS 0.006422f
C206 B.n166 VSUBS 0.006422f
C207 B.n167 VSUBS 0.006422f
C208 B.n168 VSUBS 0.006422f
C209 B.n169 VSUBS 0.006422f
C210 B.n170 VSUBS 0.006422f
C211 B.n171 VSUBS 0.006422f
C212 B.n172 VSUBS 0.006422f
C213 B.n173 VSUBS 0.006422f
C214 B.n174 VSUBS 0.006422f
C215 B.n175 VSUBS 0.006422f
C216 B.n176 VSUBS 0.006422f
C217 B.n177 VSUBS 0.006422f
C218 B.n178 VSUBS 0.006422f
C219 B.n179 VSUBS 0.006422f
C220 B.n180 VSUBS 0.006422f
C221 B.n181 VSUBS 0.006422f
C222 B.n182 VSUBS 0.006422f
C223 B.n183 VSUBS 0.006422f
C224 B.n184 VSUBS 0.006422f
C225 B.n185 VSUBS 0.006422f
C226 B.n186 VSUBS 0.006422f
C227 B.n187 VSUBS 0.006422f
C228 B.n188 VSUBS 0.006422f
C229 B.n189 VSUBS 0.006422f
C230 B.n190 VSUBS 0.006422f
C231 B.n191 VSUBS 0.006422f
C232 B.n192 VSUBS 0.006422f
C233 B.n193 VSUBS 0.006422f
C234 B.n194 VSUBS 0.006422f
C235 B.n195 VSUBS 0.006422f
C236 B.n196 VSUBS 0.004439f
C237 B.n197 VSUBS 0.014879f
C238 B.n198 VSUBS 0.005194f
C239 B.n199 VSUBS 0.006422f
C240 B.n200 VSUBS 0.006422f
C241 B.n201 VSUBS 0.006422f
C242 B.n202 VSUBS 0.006422f
C243 B.n203 VSUBS 0.006422f
C244 B.n204 VSUBS 0.006422f
C245 B.n205 VSUBS 0.006422f
C246 B.n206 VSUBS 0.006422f
C247 B.n207 VSUBS 0.006422f
C248 B.n208 VSUBS 0.006422f
C249 B.n209 VSUBS 0.006422f
C250 B.n210 VSUBS 0.005194f
C251 B.n211 VSUBS 0.006422f
C252 B.n212 VSUBS 0.006422f
C253 B.n213 VSUBS 0.004439f
C254 B.n214 VSUBS 0.006422f
C255 B.n215 VSUBS 0.006422f
C256 B.n216 VSUBS 0.006422f
C257 B.n217 VSUBS 0.006422f
C258 B.n218 VSUBS 0.006422f
C259 B.n219 VSUBS 0.006422f
C260 B.n220 VSUBS 0.006422f
C261 B.n221 VSUBS 0.006422f
C262 B.n222 VSUBS 0.006422f
C263 B.n223 VSUBS 0.006422f
C264 B.n224 VSUBS 0.006422f
C265 B.n225 VSUBS 0.006422f
C266 B.n226 VSUBS 0.006422f
C267 B.n227 VSUBS 0.006422f
C268 B.n228 VSUBS 0.006422f
C269 B.n229 VSUBS 0.006422f
C270 B.n230 VSUBS 0.006422f
C271 B.n231 VSUBS 0.006422f
C272 B.n232 VSUBS 0.006422f
C273 B.n233 VSUBS 0.006422f
C274 B.n234 VSUBS 0.006422f
C275 B.n235 VSUBS 0.006422f
C276 B.n236 VSUBS 0.006422f
C277 B.n237 VSUBS 0.006422f
C278 B.n238 VSUBS 0.006422f
C279 B.n239 VSUBS 0.006422f
C280 B.n240 VSUBS 0.006422f
C281 B.n241 VSUBS 0.006422f
C282 B.n242 VSUBS 0.006422f
C283 B.n243 VSUBS 0.006422f
C284 B.n244 VSUBS 0.006422f
C285 B.n245 VSUBS 0.006422f
C286 B.n246 VSUBS 0.006422f
C287 B.n247 VSUBS 0.006422f
C288 B.n248 VSUBS 0.006422f
C289 B.n249 VSUBS 0.006422f
C290 B.n250 VSUBS 0.014423f
C291 B.n251 VSUBS 0.013532f
C292 B.n252 VSUBS 0.013532f
C293 B.n253 VSUBS 0.006422f
C294 B.n254 VSUBS 0.006422f
C295 B.n255 VSUBS 0.006422f
C296 B.n256 VSUBS 0.006422f
C297 B.n257 VSUBS 0.006422f
C298 B.n258 VSUBS 0.006422f
C299 B.n259 VSUBS 0.006422f
C300 B.n260 VSUBS 0.006422f
C301 B.n261 VSUBS 0.006422f
C302 B.n262 VSUBS 0.006422f
C303 B.n263 VSUBS 0.006422f
C304 B.n264 VSUBS 0.006422f
C305 B.n265 VSUBS 0.006422f
C306 B.n266 VSUBS 0.006422f
C307 B.n267 VSUBS 0.006422f
C308 B.n268 VSUBS 0.006422f
C309 B.n269 VSUBS 0.006422f
C310 B.n270 VSUBS 0.006422f
C311 B.n271 VSUBS 0.006422f
C312 B.n272 VSUBS 0.006422f
C313 B.n273 VSUBS 0.006422f
C314 B.n274 VSUBS 0.006422f
C315 B.n275 VSUBS 0.006422f
C316 B.n276 VSUBS 0.006422f
C317 B.n277 VSUBS 0.006422f
C318 B.n278 VSUBS 0.006422f
C319 B.n279 VSUBS 0.006422f
C320 B.n280 VSUBS 0.006422f
C321 B.n281 VSUBS 0.006422f
C322 B.n282 VSUBS 0.006422f
C323 B.n283 VSUBS 0.006422f
C324 B.n284 VSUBS 0.006422f
C325 B.n285 VSUBS 0.006422f
C326 B.n286 VSUBS 0.006422f
C327 B.n287 VSUBS 0.006422f
C328 B.n288 VSUBS 0.006422f
C329 B.n289 VSUBS 0.006422f
C330 B.n290 VSUBS 0.006422f
C331 B.n291 VSUBS 0.006422f
C332 B.n292 VSUBS 0.006422f
C333 B.n293 VSUBS 0.006422f
C334 B.n294 VSUBS 0.006422f
C335 B.n295 VSUBS 0.006422f
C336 B.n296 VSUBS 0.006422f
C337 B.n297 VSUBS 0.006422f
C338 B.n298 VSUBS 0.006422f
C339 B.n299 VSUBS 0.006422f
C340 B.n300 VSUBS 0.006422f
C341 B.n301 VSUBS 0.006422f
C342 B.n302 VSUBS 0.006422f
C343 B.n303 VSUBS 0.006422f
C344 B.n304 VSUBS 0.006422f
C345 B.n305 VSUBS 0.006422f
C346 B.n306 VSUBS 0.006422f
C347 B.n307 VSUBS 0.006422f
C348 B.n308 VSUBS 0.006422f
C349 B.n309 VSUBS 0.006422f
C350 B.n310 VSUBS 0.006422f
C351 B.n311 VSUBS 0.006422f
C352 B.n312 VSUBS 0.006422f
C353 B.n313 VSUBS 0.006422f
C354 B.n314 VSUBS 0.006422f
C355 B.n315 VSUBS 0.006422f
C356 B.n316 VSUBS 0.006422f
C357 B.n317 VSUBS 0.006422f
C358 B.n318 VSUBS 0.006422f
C359 B.n319 VSUBS 0.006422f
C360 B.n320 VSUBS 0.006422f
C361 B.n321 VSUBS 0.006422f
C362 B.n322 VSUBS 0.006422f
C363 B.n323 VSUBS 0.006422f
C364 B.n324 VSUBS 0.006422f
C365 B.n325 VSUBS 0.006422f
C366 B.n326 VSUBS 0.013532f
C367 B.n327 VSUBS 0.014381f
C368 B.n328 VSUBS 0.013574f
C369 B.n329 VSUBS 0.006422f
C370 B.n330 VSUBS 0.006422f
C371 B.n331 VSUBS 0.006422f
C372 B.n332 VSUBS 0.006422f
C373 B.n333 VSUBS 0.006422f
C374 B.n334 VSUBS 0.006422f
C375 B.n335 VSUBS 0.006422f
C376 B.n336 VSUBS 0.006422f
C377 B.n337 VSUBS 0.006422f
C378 B.n338 VSUBS 0.006422f
C379 B.n339 VSUBS 0.006422f
C380 B.n340 VSUBS 0.006422f
C381 B.n341 VSUBS 0.006422f
C382 B.n342 VSUBS 0.006422f
C383 B.n343 VSUBS 0.006422f
C384 B.n344 VSUBS 0.006422f
C385 B.n345 VSUBS 0.006422f
C386 B.n346 VSUBS 0.006422f
C387 B.n347 VSUBS 0.006422f
C388 B.n348 VSUBS 0.006422f
C389 B.n349 VSUBS 0.006422f
C390 B.n350 VSUBS 0.006422f
C391 B.n351 VSUBS 0.006422f
C392 B.n352 VSUBS 0.006422f
C393 B.n353 VSUBS 0.006422f
C394 B.n354 VSUBS 0.006422f
C395 B.n355 VSUBS 0.006422f
C396 B.n356 VSUBS 0.006422f
C397 B.n357 VSUBS 0.006422f
C398 B.n358 VSUBS 0.006422f
C399 B.n359 VSUBS 0.006422f
C400 B.n360 VSUBS 0.006422f
C401 B.n361 VSUBS 0.006422f
C402 B.n362 VSUBS 0.006422f
C403 B.n363 VSUBS 0.006422f
C404 B.n364 VSUBS 0.006422f
C405 B.n365 VSUBS 0.004439f
C406 B.n366 VSUBS 0.006422f
C407 B.n367 VSUBS 0.006422f
C408 B.n368 VSUBS 0.005194f
C409 B.n369 VSUBS 0.006422f
C410 B.n370 VSUBS 0.006422f
C411 B.n371 VSUBS 0.006422f
C412 B.n372 VSUBS 0.006422f
C413 B.n373 VSUBS 0.006422f
C414 B.n374 VSUBS 0.006422f
C415 B.n375 VSUBS 0.006422f
C416 B.n376 VSUBS 0.006422f
C417 B.n377 VSUBS 0.006422f
C418 B.n378 VSUBS 0.006422f
C419 B.n379 VSUBS 0.006422f
C420 B.n380 VSUBS 0.005194f
C421 B.n381 VSUBS 0.014879f
C422 B.n382 VSUBS 0.004439f
C423 B.n383 VSUBS 0.006422f
C424 B.n384 VSUBS 0.006422f
C425 B.n385 VSUBS 0.006422f
C426 B.n386 VSUBS 0.006422f
C427 B.n387 VSUBS 0.006422f
C428 B.n388 VSUBS 0.006422f
C429 B.n389 VSUBS 0.006422f
C430 B.n390 VSUBS 0.006422f
C431 B.n391 VSUBS 0.006422f
C432 B.n392 VSUBS 0.006422f
C433 B.n393 VSUBS 0.006422f
C434 B.n394 VSUBS 0.006422f
C435 B.n395 VSUBS 0.006422f
C436 B.n396 VSUBS 0.006422f
C437 B.n397 VSUBS 0.006422f
C438 B.n398 VSUBS 0.006422f
C439 B.n399 VSUBS 0.006422f
C440 B.n400 VSUBS 0.006422f
C441 B.n401 VSUBS 0.006422f
C442 B.n402 VSUBS 0.006422f
C443 B.n403 VSUBS 0.006422f
C444 B.n404 VSUBS 0.006422f
C445 B.n405 VSUBS 0.006422f
C446 B.n406 VSUBS 0.006422f
C447 B.n407 VSUBS 0.006422f
C448 B.n408 VSUBS 0.006422f
C449 B.n409 VSUBS 0.006422f
C450 B.n410 VSUBS 0.006422f
C451 B.n411 VSUBS 0.006422f
C452 B.n412 VSUBS 0.006422f
C453 B.n413 VSUBS 0.006422f
C454 B.n414 VSUBS 0.006422f
C455 B.n415 VSUBS 0.006422f
C456 B.n416 VSUBS 0.006422f
C457 B.n417 VSUBS 0.006422f
C458 B.n418 VSUBS 0.006422f
C459 B.n419 VSUBS 0.014423f
C460 B.n420 VSUBS 0.014423f
C461 B.n421 VSUBS 0.013532f
C462 B.n422 VSUBS 0.006422f
C463 B.n423 VSUBS 0.006422f
C464 B.n424 VSUBS 0.006422f
C465 B.n425 VSUBS 0.006422f
C466 B.n426 VSUBS 0.006422f
C467 B.n427 VSUBS 0.006422f
C468 B.n428 VSUBS 0.006422f
C469 B.n429 VSUBS 0.006422f
C470 B.n430 VSUBS 0.006422f
C471 B.n431 VSUBS 0.006422f
C472 B.n432 VSUBS 0.006422f
C473 B.n433 VSUBS 0.006422f
C474 B.n434 VSUBS 0.006422f
C475 B.n435 VSUBS 0.006422f
C476 B.n436 VSUBS 0.006422f
C477 B.n437 VSUBS 0.006422f
C478 B.n438 VSUBS 0.006422f
C479 B.n439 VSUBS 0.006422f
C480 B.n440 VSUBS 0.006422f
C481 B.n441 VSUBS 0.006422f
C482 B.n442 VSUBS 0.006422f
C483 B.n443 VSUBS 0.006422f
C484 B.n444 VSUBS 0.006422f
C485 B.n445 VSUBS 0.006422f
C486 B.n446 VSUBS 0.006422f
C487 B.n447 VSUBS 0.006422f
C488 B.n448 VSUBS 0.006422f
C489 B.n449 VSUBS 0.006422f
C490 B.n450 VSUBS 0.006422f
C491 B.n451 VSUBS 0.006422f
C492 B.n452 VSUBS 0.006422f
C493 B.n453 VSUBS 0.006422f
C494 B.n454 VSUBS 0.006422f
C495 B.n455 VSUBS 0.006422f
C496 B.n456 VSUBS 0.006422f
C497 B.n457 VSUBS 0.006422f
C498 B.n458 VSUBS 0.006422f
C499 B.n459 VSUBS 0.014542f
C500 VDD1.n0 VSUBS 0.014197f
C501 VDD1.n1 VSUBS 0.032021f
C502 VDD1.n2 VSUBS 0.014344f
C503 VDD1.n3 VSUBS 0.025212f
C504 VDD1.n4 VSUBS 0.013547f
C505 VDD1.n5 VSUBS 0.032021f
C506 VDD1.n6 VSUBS 0.014344f
C507 VDD1.n7 VSUBS 0.025212f
C508 VDD1.n8 VSUBS 0.013547f
C509 VDD1.n9 VSUBS 0.024016f
C510 VDD1.n10 VSUBS 0.024085f
C511 VDD1.t6 VSUBS 0.068849f
C512 VDD1.n11 VSUBS 0.136453f
C513 VDD1.n12 VSUBS 0.633901f
C514 VDD1.n13 VSUBS 0.013547f
C515 VDD1.n14 VSUBS 0.014344f
C516 VDD1.n15 VSUBS 0.032021f
C517 VDD1.n16 VSUBS 0.032021f
C518 VDD1.n17 VSUBS 0.014344f
C519 VDD1.n18 VSUBS 0.013547f
C520 VDD1.n19 VSUBS 0.025212f
C521 VDD1.n20 VSUBS 0.025212f
C522 VDD1.n21 VSUBS 0.013547f
C523 VDD1.n22 VSUBS 0.014344f
C524 VDD1.n23 VSUBS 0.032021f
C525 VDD1.n24 VSUBS 0.032021f
C526 VDD1.n25 VSUBS 0.014344f
C527 VDD1.n26 VSUBS 0.013547f
C528 VDD1.n27 VSUBS 0.025212f
C529 VDD1.n28 VSUBS 0.06413f
C530 VDD1.n29 VSUBS 0.013547f
C531 VDD1.n30 VSUBS 0.014344f
C532 VDD1.n31 VSUBS 0.071701f
C533 VDD1.n32 VSUBS 0.066571f
C534 VDD1.t0 VSUBS 0.130096f
C535 VDD1.t2 VSUBS 0.130096f
C536 VDD1.n33 VSUBS 0.900319f
C537 VDD1.n34 VSUBS 0.605805f
C538 VDD1.n35 VSUBS 0.014197f
C539 VDD1.n36 VSUBS 0.032021f
C540 VDD1.n37 VSUBS 0.014344f
C541 VDD1.n38 VSUBS 0.025212f
C542 VDD1.n39 VSUBS 0.013547f
C543 VDD1.n40 VSUBS 0.032021f
C544 VDD1.n41 VSUBS 0.014344f
C545 VDD1.n42 VSUBS 0.025212f
C546 VDD1.n43 VSUBS 0.013547f
C547 VDD1.n44 VSUBS 0.024016f
C548 VDD1.n45 VSUBS 0.024085f
C549 VDD1.t3 VSUBS 0.068849f
C550 VDD1.n46 VSUBS 0.136453f
C551 VDD1.n47 VSUBS 0.633902f
C552 VDD1.n48 VSUBS 0.013547f
C553 VDD1.n49 VSUBS 0.014344f
C554 VDD1.n50 VSUBS 0.032021f
C555 VDD1.n51 VSUBS 0.032021f
C556 VDD1.n52 VSUBS 0.014344f
C557 VDD1.n53 VSUBS 0.013547f
C558 VDD1.n54 VSUBS 0.025212f
C559 VDD1.n55 VSUBS 0.025212f
C560 VDD1.n56 VSUBS 0.013547f
C561 VDD1.n57 VSUBS 0.014344f
C562 VDD1.n58 VSUBS 0.032021f
C563 VDD1.n59 VSUBS 0.032021f
C564 VDD1.n60 VSUBS 0.014344f
C565 VDD1.n61 VSUBS 0.013547f
C566 VDD1.n62 VSUBS 0.025212f
C567 VDD1.n63 VSUBS 0.06413f
C568 VDD1.n64 VSUBS 0.013547f
C569 VDD1.n65 VSUBS 0.014344f
C570 VDD1.n66 VSUBS 0.071701f
C571 VDD1.n67 VSUBS 0.066571f
C572 VDD1.t4 VSUBS 0.130096f
C573 VDD1.t5 VSUBS 0.130096f
C574 VDD1.n68 VSUBS 0.900317f
C575 VDD1.n69 VSUBS 0.600496f
C576 VDD1.t8 VSUBS 0.130096f
C577 VDD1.t9 VSUBS 0.130096f
C578 VDD1.n70 VSUBS 0.903516f
C579 VDD1.n71 VSUBS 1.81513f
C580 VDD1.t7 VSUBS 0.130096f
C581 VDD1.t1 VSUBS 0.130096f
C582 VDD1.n72 VSUBS 0.900315f
C583 VDD1.n73 VSUBS 2.13214f
C584 VP.n0 VSUBS 0.104072f
C585 VP.t5 VSUBS 0.732088f
C586 VP.n1 VSUBS 0.347899f
C587 VP.n2 VSUBS 0.104072f
C588 VP.t8 VSUBS 0.732088f
C589 VP.t2 VSUBS 0.732088f
C590 VP.t7 VSUBS 0.732088f
C591 VP.n3 VSUBS 0.326707f
C592 VP.t9 VSUBS 0.732088f
C593 VP.t3 VSUBS 0.758091f
C594 VP.n4 VSUBS 0.3096f
C595 VP.n5 VSUBS 0.347899f
C596 VP.n6 VSUBS 0.347899f
C597 VP.n7 VSUBS 0.347899f
C598 VP.n8 VSUBS 0.333721f
C599 VP.n9 VSUBS 2.2164f
C600 VP.t6 VSUBS 0.732088f
C601 VP.n10 VSUBS 0.333721f
C602 VP.n11 VSUBS 2.27512f
C603 VP.n12 VSUBS 0.104072f
C604 VP.n13 VSUBS 0.124964f
C605 VP.t4 VSUBS 0.732088f
C606 VP.n14 VSUBS 0.347899f
C607 VP.t1 VSUBS 0.732088f
C608 VP.n15 VSUBS 0.347899f
C609 VP.t0 VSUBS 0.732088f
C610 VP.n16 VSUBS 0.333721f
C611 VP.n17 VSUBS 0.069314f
C612 VTAIL.t15 VSUBS 0.155043f
C613 VTAIL.t14 VSUBS 0.155043f
C614 VTAIL.n0 VSUBS 0.967022f
C615 VTAIL.n1 VSUBS 0.694083f
C616 VTAIL.n2 VSUBS 0.016919f
C617 VTAIL.n3 VSUBS 0.038162f
C618 VTAIL.n4 VSUBS 0.017095f
C619 VTAIL.n5 VSUBS 0.030046f
C620 VTAIL.n6 VSUBS 0.016145f
C621 VTAIL.n7 VSUBS 0.038162f
C622 VTAIL.n8 VSUBS 0.017095f
C623 VTAIL.n9 VSUBS 0.030046f
C624 VTAIL.n10 VSUBS 0.016145f
C625 VTAIL.n11 VSUBS 0.028621f
C626 VTAIL.n12 VSUBS 0.028703f
C627 VTAIL.t2 VSUBS 0.082051f
C628 VTAIL.n13 VSUBS 0.162619f
C629 VTAIL.n14 VSUBS 0.755458f
C630 VTAIL.n15 VSUBS 0.016145f
C631 VTAIL.n16 VSUBS 0.017095f
C632 VTAIL.n17 VSUBS 0.038162f
C633 VTAIL.n18 VSUBS 0.038162f
C634 VTAIL.n19 VSUBS 0.017095f
C635 VTAIL.n20 VSUBS 0.016145f
C636 VTAIL.n21 VSUBS 0.030046f
C637 VTAIL.n22 VSUBS 0.030046f
C638 VTAIL.n23 VSUBS 0.016145f
C639 VTAIL.n24 VSUBS 0.017095f
C640 VTAIL.n25 VSUBS 0.038162f
C641 VTAIL.n26 VSUBS 0.038162f
C642 VTAIL.n27 VSUBS 0.017095f
C643 VTAIL.n28 VSUBS 0.016145f
C644 VTAIL.n29 VSUBS 0.030046f
C645 VTAIL.n30 VSUBS 0.076428f
C646 VTAIL.n31 VSUBS 0.016145f
C647 VTAIL.n32 VSUBS 0.017095f
C648 VTAIL.n33 VSUBS 0.08545f
C649 VTAIL.n34 VSUBS 0.056444f
C650 VTAIL.n35 VSUBS 0.193562f
C651 VTAIL.t0 VSUBS 0.155043f
C652 VTAIL.t7 VSUBS 0.155043f
C653 VTAIL.n36 VSUBS 0.967022f
C654 VTAIL.n37 VSUBS 0.70243f
C655 VTAIL.t1 VSUBS 0.155043f
C656 VTAIL.t8 VSUBS 0.155043f
C657 VTAIL.n38 VSUBS 0.967022f
C658 VTAIL.n39 VSUBS 1.73486f
C659 VTAIL.t18 VSUBS 0.155043f
C660 VTAIL.t16 VSUBS 0.155043f
C661 VTAIL.n40 VSUBS 0.967026f
C662 VTAIL.n41 VSUBS 1.73485f
C663 VTAIL.t12 VSUBS 0.155043f
C664 VTAIL.t19 VSUBS 0.155043f
C665 VTAIL.n42 VSUBS 0.967026f
C666 VTAIL.n43 VSUBS 0.702426f
C667 VTAIL.n44 VSUBS 0.016919f
C668 VTAIL.n45 VSUBS 0.038162f
C669 VTAIL.n46 VSUBS 0.017095f
C670 VTAIL.n47 VSUBS 0.030046f
C671 VTAIL.n48 VSUBS 0.016145f
C672 VTAIL.n49 VSUBS 0.038162f
C673 VTAIL.n50 VSUBS 0.017095f
C674 VTAIL.n51 VSUBS 0.030046f
C675 VTAIL.n52 VSUBS 0.016145f
C676 VTAIL.n53 VSUBS 0.028621f
C677 VTAIL.n54 VSUBS 0.028703f
C678 VTAIL.t17 VSUBS 0.082051f
C679 VTAIL.n55 VSUBS 0.162619f
C680 VTAIL.n56 VSUBS 0.755458f
C681 VTAIL.n57 VSUBS 0.016145f
C682 VTAIL.n58 VSUBS 0.017095f
C683 VTAIL.n59 VSUBS 0.038162f
C684 VTAIL.n60 VSUBS 0.038162f
C685 VTAIL.n61 VSUBS 0.017095f
C686 VTAIL.n62 VSUBS 0.016145f
C687 VTAIL.n63 VSUBS 0.030046f
C688 VTAIL.n64 VSUBS 0.030046f
C689 VTAIL.n65 VSUBS 0.016145f
C690 VTAIL.n66 VSUBS 0.017095f
C691 VTAIL.n67 VSUBS 0.038162f
C692 VTAIL.n68 VSUBS 0.038162f
C693 VTAIL.n69 VSUBS 0.017095f
C694 VTAIL.n70 VSUBS 0.016145f
C695 VTAIL.n71 VSUBS 0.030046f
C696 VTAIL.n72 VSUBS 0.076428f
C697 VTAIL.n73 VSUBS 0.016145f
C698 VTAIL.n74 VSUBS 0.017095f
C699 VTAIL.n75 VSUBS 0.08545f
C700 VTAIL.n76 VSUBS 0.056444f
C701 VTAIL.n77 VSUBS 0.193562f
C702 VTAIL.t6 VSUBS 0.155043f
C703 VTAIL.t3 VSUBS 0.155043f
C704 VTAIL.n78 VSUBS 0.967026f
C705 VTAIL.n79 VSUBS 0.708268f
C706 VTAIL.t4 VSUBS 0.155043f
C707 VTAIL.t9 VSUBS 0.155043f
C708 VTAIL.n80 VSUBS 0.967026f
C709 VTAIL.n81 VSUBS 0.702426f
C710 VTAIL.n82 VSUBS 0.016919f
C711 VTAIL.n83 VSUBS 0.038162f
C712 VTAIL.n84 VSUBS 0.017095f
C713 VTAIL.n85 VSUBS 0.030046f
C714 VTAIL.n86 VSUBS 0.016145f
C715 VTAIL.n87 VSUBS 0.038162f
C716 VTAIL.n88 VSUBS 0.017095f
C717 VTAIL.n89 VSUBS 0.030046f
C718 VTAIL.n90 VSUBS 0.016145f
C719 VTAIL.n91 VSUBS 0.028621f
C720 VTAIL.n92 VSUBS 0.028703f
C721 VTAIL.t5 VSUBS 0.082051f
C722 VTAIL.n93 VSUBS 0.162619f
C723 VTAIL.n94 VSUBS 0.755458f
C724 VTAIL.n95 VSUBS 0.016145f
C725 VTAIL.n96 VSUBS 0.017095f
C726 VTAIL.n97 VSUBS 0.038162f
C727 VTAIL.n98 VSUBS 0.038162f
C728 VTAIL.n99 VSUBS 0.017095f
C729 VTAIL.n100 VSUBS 0.016145f
C730 VTAIL.n101 VSUBS 0.030046f
C731 VTAIL.n102 VSUBS 0.030046f
C732 VTAIL.n103 VSUBS 0.016145f
C733 VTAIL.n104 VSUBS 0.017095f
C734 VTAIL.n105 VSUBS 0.038162f
C735 VTAIL.n106 VSUBS 0.038162f
C736 VTAIL.n107 VSUBS 0.017095f
C737 VTAIL.n108 VSUBS 0.016145f
C738 VTAIL.n109 VSUBS 0.030046f
C739 VTAIL.n110 VSUBS 0.076428f
C740 VTAIL.n111 VSUBS 0.016145f
C741 VTAIL.n112 VSUBS 0.017095f
C742 VTAIL.n113 VSUBS 0.08545f
C743 VTAIL.n114 VSUBS 0.056444f
C744 VTAIL.n115 VSUBS 1.14086f
C745 VTAIL.n116 VSUBS 0.016919f
C746 VTAIL.n117 VSUBS 0.038162f
C747 VTAIL.n118 VSUBS 0.017095f
C748 VTAIL.n119 VSUBS 0.030046f
C749 VTAIL.n120 VSUBS 0.016145f
C750 VTAIL.n121 VSUBS 0.038162f
C751 VTAIL.n122 VSUBS 0.017095f
C752 VTAIL.n123 VSUBS 0.030046f
C753 VTAIL.n124 VSUBS 0.016145f
C754 VTAIL.n125 VSUBS 0.028621f
C755 VTAIL.n126 VSUBS 0.028703f
C756 VTAIL.t10 VSUBS 0.082051f
C757 VTAIL.n127 VSUBS 0.162619f
C758 VTAIL.n128 VSUBS 0.755458f
C759 VTAIL.n129 VSUBS 0.016145f
C760 VTAIL.n130 VSUBS 0.017095f
C761 VTAIL.n131 VSUBS 0.038162f
C762 VTAIL.n132 VSUBS 0.038162f
C763 VTAIL.n133 VSUBS 0.017095f
C764 VTAIL.n134 VSUBS 0.016145f
C765 VTAIL.n135 VSUBS 0.030046f
C766 VTAIL.n136 VSUBS 0.030046f
C767 VTAIL.n137 VSUBS 0.016145f
C768 VTAIL.n138 VSUBS 0.017095f
C769 VTAIL.n139 VSUBS 0.038162f
C770 VTAIL.n140 VSUBS 0.038162f
C771 VTAIL.n141 VSUBS 0.017095f
C772 VTAIL.n142 VSUBS 0.016145f
C773 VTAIL.n143 VSUBS 0.030046f
C774 VTAIL.n144 VSUBS 0.076428f
C775 VTAIL.n145 VSUBS 0.016145f
C776 VTAIL.n146 VSUBS 0.017095f
C777 VTAIL.n147 VSUBS 0.08545f
C778 VTAIL.n148 VSUBS 0.056444f
C779 VTAIL.n149 VSUBS 1.14086f
C780 VTAIL.t13 VSUBS 0.155043f
C781 VTAIL.t11 VSUBS 0.155043f
C782 VTAIL.n150 VSUBS 0.967022f
C783 VTAIL.n151 VSUBS 0.63733f
C784 VDD2.n0 VSUBS 0.01408f
C785 VDD2.n1 VSUBS 0.031758f
C786 VDD2.n2 VSUBS 0.014227f
C787 VDD2.n3 VSUBS 0.025004f
C788 VDD2.n4 VSUBS 0.013436f
C789 VDD2.n5 VSUBS 0.031758f
C790 VDD2.n6 VSUBS 0.014227f
C791 VDD2.n7 VSUBS 0.025004f
C792 VDD2.n8 VSUBS 0.013436f
C793 VDD2.n9 VSUBS 0.023819f
C794 VDD2.n10 VSUBS 0.023887f
C795 VDD2.t3 VSUBS 0.068283f
C796 VDD2.n11 VSUBS 0.135331f
C797 VDD2.n12 VSUBS 0.628693f
C798 VDD2.n13 VSUBS 0.013436f
C799 VDD2.n14 VSUBS 0.014227f
C800 VDD2.n15 VSUBS 0.031758f
C801 VDD2.n16 VSUBS 0.031758f
C802 VDD2.n17 VSUBS 0.014227f
C803 VDD2.n18 VSUBS 0.013436f
C804 VDD2.n19 VSUBS 0.025004f
C805 VDD2.n20 VSUBS 0.025004f
C806 VDD2.n21 VSUBS 0.013436f
C807 VDD2.n22 VSUBS 0.014227f
C808 VDD2.n23 VSUBS 0.031758f
C809 VDD2.n24 VSUBS 0.031758f
C810 VDD2.n25 VSUBS 0.014227f
C811 VDD2.n26 VSUBS 0.013436f
C812 VDD2.n27 VSUBS 0.025004f
C813 VDD2.n28 VSUBS 0.063603f
C814 VDD2.n29 VSUBS 0.013436f
C815 VDD2.n30 VSUBS 0.014227f
C816 VDD2.n31 VSUBS 0.071112f
C817 VDD2.n32 VSUBS 0.066024f
C818 VDD2.t9 VSUBS 0.129027f
C819 VDD2.t6 VSUBS 0.129027f
C820 VDD2.n33 VSUBS 0.892919f
C821 VDD2.n34 VSUBS 0.595561f
C822 VDD2.t1 VSUBS 0.129027f
C823 VDD2.t2 VSUBS 0.129027f
C824 VDD2.n35 VSUBS 0.896091f
C825 VDD2.n36 VSUBS 1.72708f
C826 VDD2.n37 VSUBS 0.01408f
C827 VDD2.n38 VSUBS 0.031758f
C828 VDD2.n39 VSUBS 0.014227f
C829 VDD2.n40 VSUBS 0.025004f
C830 VDD2.n41 VSUBS 0.013436f
C831 VDD2.n42 VSUBS 0.031758f
C832 VDD2.n43 VSUBS 0.014227f
C833 VDD2.n44 VSUBS 0.025004f
C834 VDD2.n45 VSUBS 0.013436f
C835 VDD2.n46 VSUBS 0.023819f
C836 VDD2.n47 VSUBS 0.023887f
C837 VDD2.t8 VSUBS 0.068283f
C838 VDD2.n48 VSUBS 0.135331f
C839 VDD2.n49 VSUBS 0.628693f
C840 VDD2.n50 VSUBS 0.013436f
C841 VDD2.n51 VSUBS 0.014227f
C842 VDD2.n52 VSUBS 0.031758f
C843 VDD2.n53 VSUBS 0.031758f
C844 VDD2.n54 VSUBS 0.014227f
C845 VDD2.n55 VSUBS 0.013436f
C846 VDD2.n56 VSUBS 0.025004f
C847 VDD2.n57 VSUBS 0.025004f
C848 VDD2.n58 VSUBS 0.013436f
C849 VDD2.n59 VSUBS 0.014227f
C850 VDD2.n60 VSUBS 0.031758f
C851 VDD2.n61 VSUBS 0.031758f
C852 VDD2.n62 VSUBS 0.014227f
C853 VDD2.n63 VSUBS 0.013436f
C854 VDD2.n64 VSUBS 0.025004f
C855 VDD2.n65 VSUBS 0.063603f
C856 VDD2.n66 VSUBS 0.013436f
C857 VDD2.n67 VSUBS 0.014227f
C858 VDD2.n68 VSUBS 0.071112f
C859 VDD2.n69 VSUBS 0.064201f
C860 VDD2.n70 VSUBS 1.69319f
C861 VDD2.t4 VSUBS 0.129027f
C862 VDD2.t0 VSUBS 0.129027f
C863 VDD2.n71 VSUBS 0.892921f
C864 VDD2.n72 VSUBS 0.485584f
C865 VDD2.t7 VSUBS 0.129027f
C866 VDD2.t5 VSUBS 0.129027f
C867 VDD2.n73 VSUBS 0.896065f
C868 VN.n0 VSUBS 0.100293f
C869 VN.t5 VSUBS 0.705503f
C870 VN.n1 VSUBS 0.335266f
C871 VN.t4 VSUBS 0.730562f
C872 VN.n2 VSUBS 0.298358f
C873 VN.n3 VSUBS 0.314844f
C874 VN.t6 VSUBS 0.705503f
C875 VN.n4 VSUBS 0.335266f
C876 VN.t8 VSUBS 0.705503f
C877 VN.n5 VSUBS 0.335266f
C878 VN.t9 VSUBS 0.705503f
C879 VN.n6 VSUBS 0.321602f
C880 VN.n7 VSUBS 0.066797f
C881 VN.n8 VSUBS 0.100293f
C882 VN.t0 VSUBS 0.705503f
C883 VN.n9 VSUBS 0.335266f
C884 VN.t7 VSUBS 0.705503f
C885 VN.t2 VSUBS 0.730562f
C886 VN.n10 VSUBS 0.298358f
C887 VN.n11 VSUBS 0.314844f
C888 VN.n12 VSUBS 0.335266f
C889 VN.t3 VSUBS 0.705503f
C890 VN.n13 VSUBS 0.335266f
C891 VN.t1 VSUBS 0.705503f
C892 VN.n14 VSUBS 0.321602f
C893 VN.n15 VSUBS 2.17569f
.ends

