* NGSPICE file created from diff_pair_sample_1142.ext - technology: sky130A

.subckt diff_pair_sample_1142 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t1 VN.t0 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=7.4217 pd=38.84 as=7.4217 ps=38.84 w=19.03 l=1.05
X1 VDD1.t1 VP.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=7.4217 pd=38.84 as=7.4217 ps=38.84 w=19.03 l=1.05
X2 VDD1.t0 VP.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=7.4217 pd=38.84 as=7.4217 ps=38.84 w=19.03 l=1.05
X3 B.t15 B.t13 B.t14 B.t3 sky130_fd_pr__nfet_01v8 ad=7.4217 pd=38.84 as=0 ps=0 w=19.03 l=1.05
X4 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=7.4217 pd=38.84 as=0 ps=0 w=19.03 l=1.05
X5 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=7.4217 pd=38.84 as=0 ps=0 w=19.03 l=1.05
X6 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=7.4217 pd=38.84 as=0 ps=0 w=19.03 l=1.05
X7 VDD2.t0 VN.t1 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=7.4217 pd=38.84 as=7.4217 ps=38.84 w=19.03 l=1.05
R0 VN VN.t0 681.994
R1 VN VN.t1 635.778
R2 VTAIL.n418 VTAIL.n318 289.615
R3 VTAIL.n100 VTAIL.n0 289.615
R4 VTAIL.n312 VTAIL.n212 289.615
R5 VTAIL.n206 VTAIL.n106 289.615
R6 VTAIL.n353 VTAIL.n352 185
R7 VTAIL.n350 VTAIL.n349 185
R8 VTAIL.n359 VTAIL.n358 185
R9 VTAIL.n361 VTAIL.n360 185
R10 VTAIL.n346 VTAIL.n345 185
R11 VTAIL.n367 VTAIL.n366 185
R12 VTAIL.n369 VTAIL.n368 185
R13 VTAIL.n342 VTAIL.n341 185
R14 VTAIL.n375 VTAIL.n374 185
R15 VTAIL.n377 VTAIL.n376 185
R16 VTAIL.n338 VTAIL.n337 185
R17 VTAIL.n383 VTAIL.n382 185
R18 VTAIL.n385 VTAIL.n384 185
R19 VTAIL.n334 VTAIL.n333 185
R20 VTAIL.n391 VTAIL.n390 185
R21 VTAIL.n394 VTAIL.n393 185
R22 VTAIL.n392 VTAIL.n330 185
R23 VTAIL.n399 VTAIL.n329 185
R24 VTAIL.n401 VTAIL.n400 185
R25 VTAIL.n403 VTAIL.n402 185
R26 VTAIL.n326 VTAIL.n325 185
R27 VTAIL.n409 VTAIL.n408 185
R28 VTAIL.n411 VTAIL.n410 185
R29 VTAIL.n322 VTAIL.n321 185
R30 VTAIL.n417 VTAIL.n416 185
R31 VTAIL.n419 VTAIL.n418 185
R32 VTAIL.n35 VTAIL.n34 185
R33 VTAIL.n32 VTAIL.n31 185
R34 VTAIL.n41 VTAIL.n40 185
R35 VTAIL.n43 VTAIL.n42 185
R36 VTAIL.n28 VTAIL.n27 185
R37 VTAIL.n49 VTAIL.n48 185
R38 VTAIL.n51 VTAIL.n50 185
R39 VTAIL.n24 VTAIL.n23 185
R40 VTAIL.n57 VTAIL.n56 185
R41 VTAIL.n59 VTAIL.n58 185
R42 VTAIL.n20 VTAIL.n19 185
R43 VTAIL.n65 VTAIL.n64 185
R44 VTAIL.n67 VTAIL.n66 185
R45 VTAIL.n16 VTAIL.n15 185
R46 VTAIL.n73 VTAIL.n72 185
R47 VTAIL.n76 VTAIL.n75 185
R48 VTAIL.n74 VTAIL.n12 185
R49 VTAIL.n81 VTAIL.n11 185
R50 VTAIL.n83 VTAIL.n82 185
R51 VTAIL.n85 VTAIL.n84 185
R52 VTAIL.n8 VTAIL.n7 185
R53 VTAIL.n91 VTAIL.n90 185
R54 VTAIL.n93 VTAIL.n92 185
R55 VTAIL.n4 VTAIL.n3 185
R56 VTAIL.n99 VTAIL.n98 185
R57 VTAIL.n101 VTAIL.n100 185
R58 VTAIL.n313 VTAIL.n312 185
R59 VTAIL.n311 VTAIL.n310 185
R60 VTAIL.n216 VTAIL.n215 185
R61 VTAIL.n305 VTAIL.n304 185
R62 VTAIL.n303 VTAIL.n302 185
R63 VTAIL.n220 VTAIL.n219 185
R64 VTAIL.n297 VTAIL.n296 185
R65 VTAIL.n295 VTAIL.n294 185
R66 VTAIL.n293 VTAIL.n223 185
R67 VTAIL.n227 VTAIL.n224 185
R68 VTAIL.n288 VTAIL.n287 185
R69 VTAIL.n286 VTAIL.n285 185
R70 VTAIL.n229 VTAIL.n228 185
R71 VTAIL.n280 VTAIL.n279 185
R72 VTAIL.n278 VTAIL.n277 185
R73 VTAIL.n233 VTAIL.n232 185
R74 VTAIL.n272 VTAIL.n271 185
R75 VTAIL.n270 VTAIL.n269 185
R76 VTAIL.n237 VTAIL.n236 185
R77 VTAIL.n264 VTAIL.n263 185
R78 VTAIL.n262 VTAIL.n261 185
R79 VTAIL.n241 VTAIL.n240 185
R80 VTAIL.n256 VTAIL.n255 185
R81 VTAIL.n254 VTAIL.n253 185
R82 VTAIL.n245 VTAIL.n244 185
R83 VTAIL.n248 VTAIL.n247 185
R84 VTAIL.n207 VTAIL.n206 185
R85 VTAIL.n205 VTAIL.n204 185
R86 VTAIL.n110 VTAIL.n109 185
R87 VTAIL.n199 VTAIL.n198 185
R88 VTAIL.n197 VTAIL.n196 185
R89 VTAIL.n114 VTAIL.n113 185
R90 VTAIL.n191 VTAIL.n190 185
R91 VTAIL.n189 VTAIL.n188 185
R92 VTAIL.n187 VTAIL.n117 185
R93 VTAIL.n121 VTAIL.n118 185
R94 VTAIL.n182 VTAIL.n181 185
R95 VTAIL.n180 VTAIL.n179 185
R96 VTAIL.n123 VTAIL.n122 185
R97 VTAIL.n174 VTAIL.n173 185
R98 VTAIL.n172 VTAIL.n171 185
R99 VTAIL.n127 VTAIL.n126 185
R100 VTAIL.n166 VTAIL.n165 185
R101 VTAIL.n164 VTAIL.n163 185
R102 VTAIL.n131 VTAIL.n130 185
R103 VTAIL.n158 VTAIL.n157 185
R104 VTAIL.n156 VTAIL.n155 185
R105 VTAIL.n135 VTAIL.n134 185
R106 VTAIL.n150 VTAIL.n149 185
R107 VTAIL.n148 VTAIL.n147 185
R108 VTAIL.n139 VTAIL.n138 185
R109 VTAIL.n142 VTAIL.n141 185
R110 VTAIL.t1 VTAIL.n246 147.659
R111 VTAIL.t2 VTAIL.n140 147.659
R112 VTAIL.t3 VTAIL.n351 147.659
R113 VTAIL.t0 VTAIL.n33 147.659
R114 VTAIL.n352 VTAIL.n349 104.615
R115 VTAIL.n359 VTAIL.n349 104.615
R116 VTAIL.n360 VTAIL.n359 104.615
R117 VTAIL.n360 VTAIL.n345 104.615
R118 VTAIL.n367 VTAIL.n345 104.615
R119 VTAIL.n368 VTAIL.n367 104.615
R120 VTAIL.n368 VTAIL.n341 104.615
R121 VTAIL.n375 VTAIL.n341 104.615
R122 VTAIL.n376 VTAIL.n375 104.615
R123 VTAIL.n376 VTAIL.n337 104.615
R124 VTAIL.n383 VTAIL.n337 104.615
R125 VTAIL.n384 VTAIL.n383 104.615
R126 VTAIL.n384 VTAIL.n333 104.615
R127 VTAIL.n391 VTAIL.n333 104.615
R128 VTAIL.n393 VTAIL.n391 104.615
R129 VTAIL.n393 VTAIL.n392 104.615
R130 VTAIL.n392 VTAIL.n329 104.615
R131 VTAIL.n401 VTAIL.n329 104.615
R132 VTAIL.n402 VTAIL.n401 104.615
R133 VTAIL.n402 VTAIL.n325 104.615
R134 VTAIL.n409 VTAIL.n325 104.615
R135 VTAIL.n410 VTAIL.n409 104.615
R136 VTAIL.n410 VTAIL.n321 104.615
R137 VTAIL.n417 VTAIL.n321 104.615
R138 VTAIL.n418 VTAIL.n417 104.615
R139 VTAIL.n34 VTAIL.n31 104.615
R140 VTAIL.n41 VTAIL.n31 104.615
R141 VTAIL.n42 VTAIL.n41 104.615
R142 VTAIL.n42 VTAIL.n27 104.615
R143 VTAIL.n49 VTAIL.n27 104.615
R144 VTAIL.n50 VTAIL.n49 104.615
R145 VTAIL.n50 VTAIL.n23 104.615
R146 VTAIL.n57 VTAIL.n23 104.615
R147 VTAIL.n58 VTAIL.n57 104.615
R148 VTAIL.n58 VTAIL.n19 104.615
R149 VTAIL.n65 VTAIL.n19 104.615
R150 VTAIL.n66 VTAIL.n65 104.615
R151 VTAIL.n66 VTAIL.n15 104.615
R152 VTAIL.n73 VTAIL.n15 104.615
R153 VTAIL.n75 VTAIL.n73 104.615
R154 VTAIL.n75 VTAIL.n74 104.615
R155 VTAIL.n74 VTAIL.n11 104.615
R156 VTAIL.n83 VTAIL.n11 104.615
R157 VTAIL.n84 VTAIL.n83 104.615
R158 VTAIL.n84 VTAIL.n7 104.615
R159 VTAIL.n91 VTAIL.n7 104.615
R160 VTAIL.n92 VTAIL.n91 104.615
R161 VTAIL.n92 VTAIL.n3 104.615
R162 VTAIL.n99 VTAIL.n3 104.615
R163 VTAIL.n100 VTAIL.n99 104.615
R164 VTAIL.n312 VTAIL.n311 104.615
R165 VTAIL.n311 VTAIL.n215 104.615
R166 VTAIL.n304 VTAIL.n215 104.615
R167 VTAIL.n304 VTAIL.n303 104.615
R168 VTAIL.n303 VTAIL.n219 104.615
R169 VTAIL.n296 VTAIL.n219 104.615
R170 VTAIL.n296 VTAIL.n295 104.615
R171 VTAIL.n295 VTAIL.n223 104.615
R172 VTAIL.n227 VTAIL.n223 104.615
R173 VTAIL.n287 VTAIL.n227 104.615
R174 VTAIL.n287 VTAIL.n286 104.615
R175 VTAIL.n286 VTAIL.n228 104.615
R176 VTAIL.n279 VTAIL.n228 104.615
R177 VTAIL.n279 VTAIL.n278 104.615
R178 VTAIL.n278 VTAIL.n232 104.615
R179 VTAIL.n271 VTAIL.n232 104.615
R180 VTAIL.n271 VTAIL.n270 104.615
R181 VTAIL.n270 VTAIL.n236 104.615
R182 VTAIL.n263 VTAIL.n236 104.615
R183 VTAIL.n263 VTAIL.n262 104.615
R184 VTAIL.n262 VTAIL.n240 104.615
R185 VTAIL.n255 VTAIL.n240 104.615
R186 VTAIL.n255 VTAIL.n254 104.615
R187 VTAIL.n254 VTAIL.n244 104.615
R188 VTAIL.n247 VTAIL.n244 104.615
R189 VTAIL.n206 VTAIL.n205 104.615
R190 VTAIL.n205 VTAIL.n109 104.615
R191 VTAIL.n198 VTAIL.n109 104.615
R192 VTAIL.n198 VTAIL.n197 104.615
R193 VTAIL.n197 VTAIL.n113 104.615
R194 VTAIL.n190 VTAIL.n113 104.615
R195 VTAIL.n190 VTAIL.n189 104.615
R196 VTAIL.n189 VTAIL.n117 104.615
R197 VTAIL.n121 VTAIL.n117 104.615
R198 VTAIL.n181 VTAIL.n121 104.615
R199 VTAIL.n181 VTAIL.n180 104.615
R200 VTAIL.n180 VTAIL.n122 104.615
R201 VTAIL.n173 VTAIL.n122 104.615
R202 VTAIL.n173 VTAIL.n172 104.615
R203 VTAIL.n172 VTAIL.n126 104.615
R204 VTAIL.n165 VTAIL.n126 104.615
R205 VTAIL.n165 VTAIL.n164 104.615
R206 VTAIL.n164 VTAIL.n130 104.615
R207 VTAIL.n157 VTAIL.n130 104.615
R208 VTAIL.n157 VTAIL.n156 104.615
R209 VTAIL.n156 VTAIL.n134 104.615
R210 VTAIL.n149 VTAIL.n134 104.615
R211 VTAIL.n149 VTAIL.n148 104.615
R212 VTAIL.n148 VTAIL.n138 104.615
R213 VTAIL.n141 VTAIL.n138 104.615
R214 VTAIL.n352 VTAIL.t3 52.3082
R215 VTAIL.n34 VTAIL.t0 52.3082
R216 VTAIL.n247 VTAIL.t1 52.3082
R217 VTAIL.n141 VTAIL.t2 52.3082
R218 VTAIL.n423 VTAIL.n422 33.5429
R219 VTAIL.n105 VTAIL.n104 33.5429
R220 VTAIL.n317 VTAIL.n316 33.5429
R221 VTAIL.n211 VTAIL.n210 33.5429
R222 VTAIL.n211 VTAIL.n105 31.1686
R223 VTAIL.n423 VTAIL.n317 29.9789
R224 VTAIL.n353 VTAIL.n351 15.6677
R225 VTAIL.n35 VTAIL.n33 15.6677
R226 VTAIL.n248 VTAIL.n246 15.6677
R227 VTAIL.n142 VTAIL.n140 15.6677
R228 VTAIL.n400 VTAIL.n399 13.1884
R229 VTAIL.n82 VTAIL.n81 13.1884
R230 VTAIL.n294 VTAIL.n293 13.1884
R231 VTAIL.n188 VTAIL.n187 13.1884
R232 VTAIL.n354 VTAIL.n350 12.8005
R233 VTAIL.n398 VTAIL.n330 12.8005
R234 VTAIL.n403 VTAIL.n328 12.8005
R235 VTAIL.n36 VTAIL.n32 12.8005
R236 VTAIL.n80 VTAIL.n12 12.8005
R237 VTAIL.n85 VTAIL.n10 12.8005
R238 VTAIL.n297 VTAIL.n222 12.8005
R239 VTAIL.n292 VTAIL.n224 12.8005
R240 VTAIL.n249 VTAIL.n245 12.8005
R241 VTAIL.n191 VTAIL.n116 12.8005
R242 VTAIL.n186 VTAIL.n118 12.8005
R243 VTAIL.n143 VTAIL.n139 12.8005
R244 VTAIL.n358 VTAIL.n357 12.0247
R245 VTAIL.n395 VTAIL.n394 12.0247
R246 VTAIL.n404 VTAIL.n326 12.0247
R247 VTAIL.n40 VTAIL.n39 12.0247
R248 VTAIL.n77 VTAIL.n76 12.0247
R249 VTAIL.n86 VTAIL.n8 12.0247
R250 VTAIL.n298 VTAIL.n220 12.0247
R251 VTAIL.n289 VTAIL.n288 12.0247
R252 VTAIL.n253 VTAIL.n252 12.0247
R253 VTAIL.n192 VTAIL.n114 12.0247
R254 VTAIL.n183 VTAIL.n182 12.0247
R255 VTAIL.n147 VTAIL.n146 12.0247
R256 VTAIL.n361 VTAIL.n348 11.249
R257 VTAIL.n390 VTAIL.n332 11.249
R258 VTAIL.n408 VTAIL.n407 11.249
R259 VTAIL.n43 VTAIL.n30 11.249
R260 VTAIL.n72 VTAIL.n14 11.249
R261 VTAIL.n90 VTAIL.n89 11.249
R262 VTAIL.n302 VTAIL.n301 11.249
R263 VTAIL.n285 VTAIL.n226 11.249
R264 VTAIL.n256 VTAIL.n243 11.249
R265 VTAIL.n196 VTAIL.n195 11.249
R266 VTAIL.n179 VTAIL.n120 11.249
R267 VTAIL.n150 VTAIL.n137 11.249
R268 VTAIL.n362 VTAIL.n346 10.4732
R269 VTAIL.n389 VTAIL.n334 10.4732
R270 VTAIL.n411 VTAIL.n324 10.4732
R271 VTAIL.n44 VTAIL.n28 10.4732
R272 VTAIL.n71 VTAIL.n16 10.4732
R273 VTAIL.n93 VTAIL.n6 10.4732
R274 VTAIL.n305 VTAIL.n218 10.4732
R275 VTAIL.n284 VTAIL.n229 10.4732
R276 VTAIL.n257 VTAIL.n241 10.4732
R277 VTAIL.n199 VTAIL.n112 10.4732
R278 VTAIL.n178 VTAIL.n123 10.4732
R279 VTAIL.n151 VTAIL.n135 10.4732
R280 VTAIL.n366 VTAIL.n365 9.69747
R281 VTAIL.n386 VTAIL.n385 9.69747
R282 VTAIL.n412 VTAIL.n322 9.69747
R283 VTAIL.n48 VTAIL.n47 9.69747
R284 VTAIL.n68 VTAIL.n67 9.69747
R285 VTAIL.n94 VTAIL.n4 9.69747
R286 VTAIL.n306 VTAIL.n216 9.69747
R287 VTAIL.n281 VTAIL.n280 9.69747
R288 VTAIL.n261 VTAIL.n260 9.69747
R289 VTAIL.n200 VTAIL.n110 9.69747
R290 VTAIL.n175 VTAIL.n174 9.69747
R291 VTAIL.n155 VTAIL.n154 9.69747
R292 VTAIL.n422 VTAIL.n421 9.45567
R293 VTAIL.n104 VTAIL.n103 9.45567
R294 VTAIL.n316 VTAIL.n315 9.45567
R295 VTAIL.n210 VTAIL.n209 9.45567
R296 VTAIL.n320 VTAIL.n319 9.3005
R297 VTAIL.n415 VTAIL.n414 9.3005
R298 VTAIL.n413 VTAIL.n412 9.3005
R299 VTAIL.n324 VTAIL.n323 9.3005
R300 VTAIL.n407 VTAIL.n406 9.3005
R301 VTAIL.n405 VTAIL.n404 9.3005
R302 VTAIL.n328 VTAIL.n327 9.3005
R303 VTAIL.n373 VTAIL.n372 9.3005
R304 VTAIL.n371 VTAIL.n370 9.3005
R305 VTAIL.n344 VTAIL.n343 9.3005
R306 VTAIL.n365 VTAIL.n364 9.3005
R307 VTAIL.n363 VTAIL.n362 9.3005
R308 VTAIL.n348 VTAIL.n347 9.3005
R309 VTAIL.n357 VTAIL.n356 9.3005
R310 VTAIL.n355 VTAIL.n354 9.3005
R311 VTAIL.n340 VTAIL.n339 9.3005
R312 VTAIL.n379 VTAIL.n378 9.3005
R313 VTAIL.n381 VTAIL.n380 9.3005
R314 VTAIL.n336 VTAIL.n335 9.3005
R315 VTAIL.n387 VTAIL.n386 9.3005
R316 VTAIL.n389 VTAIL.n388 9.3005
R317 VTAIL.n332 VTAIL.n331 9.3005
R318 VTAIL.n396 VTAIL.n395 9.3005
R319 VTAIL.n398 VTAIL.n397 9.3005
R320 VTAIL.n421 VTAIL.n420 9.3005
R321 VTAIL.n2 VTAIL.n1 9.3005
R322 VTAIL.n97 VTAIL.n96 9.3005
R323 VTAIL.n95 VTAIL.n94 9.3005
R324 VTAIL.n6 VTAIL.n5 9.3005
R325 VTAIL.n89 VTAIL.n88 9.3005
R326 VTAIL.n87 VTAIL.n86 9.3005
R327 VTAIL.n10 VTAIL.n9 9.3005
R328 VTAIL.n55 VTAIL.n54 9.3005
R329 VTAIL.n53 VTAIL.n52 9.3005
R330 VTAIL.n26 VTAIL.n25 9.3005
R331 VTAIL.n47 VTAIL.n46 9.3005
R332 VTAIL.n45 VTAIL.n44 9.3005
R333 VTAIL.n30 VTAIL.n29 9.3005
R334 VTAIL.n39 VTAIL.n38 9.3005
R335 VTAIL.n37 VTAIL.n36 9.3005
R336 VTAIL.n22 VTAIL.n21 9.3005
R337 VTAIL.n61 VTAIL.n60 9.3005
R338 VTAIL.n63 VTAIL.n62 9.3005
R339 VTAIL.n18 VTAIL.n17 9.3005
R340 VTAIL.n69 VTAIL.n68 9.3005
R341 VTAIL.n71 VTAIL.n70 9.3005
R342 VTAIL.n14 VTAIL.n13 9.3005
R343 VTAIL.n78 VTAIL.n77 9.3005
R344 VTAIL.n80 VTAIL.n79 9.3005
R345 VTAIL.n103 VTAIL.n102 9.3005
R346 VTAIL.n274 VTAIL.n273 9.3005
R347 VTAIL.n276 VTAIL.n275 9.3005
R348 VTAIL.n231 VTAIL.n230 9.3005
R349 VTAIL.n282 VTAIL.n281 9.3005
R350 VTAIL.n284 VTAIL.n283 9.3005
R351 VTAIL.n226 VTAIL.n225 9.3005
R352 VTAIL.n290 VTAIL.n289 9.3005
R353 VTAIL.n292 VTAIL.n291 9.3005
R354 VTAIL.n315 VTAIL.n314 9.3005
R355 VTAIL.n214 VTAIL.n213 9.3005
R356 VTAIL.n309 VTAIL.n308 9.3005
R357 VTAIL.n307 VTAIL.n306 9.3005
R358 VTAIL.n218 VTAIL.n217 9.3005
R359 VTAIL.n301 VTAIL.n300 9.3005
R360 VTAIL.n299 VTAIL.n298 9.3005
R361 VTAIL.n222 VTAIL.n221 9.3005
R362 VTAIL.n235 VTAIL.n234 9.3005
R363 VTAIL.n268 VTAIL.n267 9.3005
R364 VTAIL.n266 VTAIL.n265 9.3005
R365 VTAIL.n239 VTAIL.n238 9.3005
R366 VTAIL.n260 VTAIL.n259 9.3005
R367 VTAIL.n258 VTAIL.n257 9.3005
R368 VTAIL.n243 VTAIL.n242 9.3005
R369 VTAIL.n252 VTAIL.n251 9.3005
R370 VTAIL.n250 VTAIL.n249 9.3005
R371 VTAIL.n168 VTAIL.n167 9.3005
R372 VTAIL.n170 VTAIL.n169 9.3005
R373 VTAIL.n125 VTAIL.n124 9.3005
R374 VTAIL.n176 VTAIL.n175 9.3005
R375 VTAIL.n178 VTAIL.n177 9.3005
R376 VTAIL.n120 VTAIL.n119 9.3005
R377 VTAIL.n184 VTAIL.n183 9.3005
R378 VTAIL.n186 VTAIL.n185 9.3005
R379 VTAIL.n209 VTAIL.n208 9.3005
R380 VTAIL.n108 VTAIL.n107 9.3005
R381 VTAIL.n203 VTAIL.n202 9.3005
R382 VTAIL.n201 VTAIL.n200 9.3005
R383 VTAIL.n112 VTAIL.n111 9.3005
R384 VTAIL.n195 VTAIL.n194 9.3005
R385 VTAIL.n193 VTAIL.n192 9.3005
R386 VTAIL.n116 VTAIL.n115 9.3005
R387 VTAIL.n129 VTAIL.n128 9.3005
R388 VTAIL.n162 VTAIL.n161 9.3005
R389 VTAIL.n160 VTAIL.n159 9.3005
R390 VTAIL.n133 VTAIL.n132 9.3005
R391 VTAIL.n154 VTAIL.n153 9.3005
R392 VTAIL.n152 VTAIL.n151 9.3005
R393 VTAIL.n137 VTAIL.n136 9.3005
R394 VTAIL.n146 VTAIL.n145 9.3005
R395 VTAIL.n144 VTAIL.n143 9.3005
R396 VTAIL.n369 VTAIL.n344 8.92171
R397 VTAIL.n382 VTAIL.n336 8.92171
R398 VTAIL.n416 VTAIL.n415 8.92171
R399 VTAIL.n51 VTAIL.n26 8.92171
R400 VTAIL.n64 VTAIL.n18 8.92171
R401 VTAIL.n98 VTAIL.n97 8.92171
R402 VTAIL.n310 VTAIL.n309 8.92171
R403 VTAIL.n277 VTAIL.n231 8.92171
R404 VTAIL.n264 VTAIL.n239 8.92171
R405 VTAIL.n204 VTAIL.n203 8.92171
R406 VTAIL.n171 VTAIL.n125 8.92171
R407 VTAIL.n158 VTAIL.n133 8.92171
R408 VTAIL.n370 VTAIL.n342 8.14595
R409 VTAIL.n381 VTAIL.n338 8.14595
R410 VTAIL.n419 VTAIL.n320 8.14595
R411 VTAIL.n52 VTAIL.n24 8.14595
R412 VTAIL.n63 VTAIL.n20 8.14595
R413 VTAIL.n101 VTAIL.n2 8.14595
R414 VTAIL.n313 VTAIL.n214 8.14595
R415 VTAIL.n276 VTAIL.n233 8.14595
R416 VTAIL.n265 VTAIL.n237 8.14595
R417 VTAIL.n207 VTAIL.n108 8.14595
R418 VTAIL.n170 VTAIL.n127 8.14595
R419 VTAIL.n159 VTAIL.n131 8.14595
R420 VTAIL.n374 VTAIL.n373 7.3702
R421 VTAIL.n378 VTAIL.n377 7.3702
R422 VTAIL.n420 VTAIL.n318 7.3702
R423 VTAIL.n56 VTAIL.n55 7.3702
R424 VTAIL.n60 VTAIL.n59 7.3702
R425 VTAIL.n102 VTAIL.n0 7.3702
R426 VTAIL.n314 VTAIL.n212 7.3702
R427 VTAIL.n273 VTAIL.n272 7.3702
R428 VTAIL.n269 VTAIL.n268 7.3702
R429 VTAIL.n208 VTAIL.n106 7.3702
R430 VTAIL.n167 VTAIL.n166 7.3702
R431 VTAIL.n163 VTAIL.n162 7.3702
R432 VTAIL.n374 VTAIL.n340 6.59444
R433 VTAIL.n377 VTAIL.n340 6.59444
R434 VTAIL.n422 VTAIL.n318 6.59444
R435 VTAIL.n56 VTAIL.n22 6.59444
R436 VTAIL.n59 VTAIL.n22 6.59444
R437 VTAIL.n104 VTAIL.n0 6.59444
R438 VTAIL.n316 VTAIL.n212 6.59444
R439 VTAIL.n272 VTAIL.n235 6.59444
R440 VTAIL.n269 VTAIL.n235 6.59444
R441 VTAIL.n210 VTAIL.n106 6.59444
R442 VTAIL.n166 VTAIL.n129 6.59444
R443 VTAIL.n163 VTAIL.n129 6.59444
R444 VTAIL.n373 VTAIL.n342 5.81868
R445 VTAIL.n378 VTAIL.n338 5.81868
R446 VTAIL.n420 VTAIL.n419 5.81868
R447 VTAIL.n55 VTAIL.n24 5.81868
R448 VTAIL.n60 VTAIL.n20 5.81868
R449 VTAIL.n102 VTAIL.n101 5.81868
R450 VTAIL.n314 VTAIL.n313 5.81868
R451 VTAIL.n273 VTAIL.n233 5.81868
R452 VTAIL.n268 VTAIL.n237 5.81868
R453 VTAIL.n208 VTAIL.n207 5.81868
R454 VTAIL.n167 VTAIL.n127 5.81868
R455 VTAIL.n162 VTAIL.n131 5.81868
R456 VTAIL.n370 VTAIL.n369 5.04292
R457 VTAIL.n382 VTAIL.n381 5.04292
R458 VTAIL.n416 VTAIL.n320 5.04292
R459 VTAIL.n52 VTAIL.n51 5.04292
R460 VTAIL.n64 VTAIL.n63 5.04292
R461 VTAIL.n98 VTAIL.n2 5.04292
R462 VTAIL.n310 VTAIL.n214 5.04292
R463 VTAIL.n277 VTAIL.n276 5.04292
R464 VTAIL.n265 VTAIL.n264 5.04292
R465 VTAIL.n204 VTAIL.n108 5.04292
R466 VTAIL.n171 VTAIL.n170 5.04292
R467 VTAIL.n159 VTAIL.n158 5.04292
R468 VTAIL.n250 VTAIL.n246 4.38563
R469 VTAIL.n144 VTAIL.n140 4.38563
R470 VTAIL.n355 VTAIL.n351 4.38563
R471 VTAIL.n37 VTAIL.n33 4.38563
R472 VTAIL.n366 VTAIL.n344 4.26717
R473 VTAIL.n385 VTAIL.n336 4.26717
R474 VTAIL.n415 VTAIL.n322 4.26717
R475 VTAIL.n48 VTAIL.n26 4.26717
R476 VTAIL.n67 VTAIL.n18 4.26717
R477 VTAIL.n97 VTAIL.n4 4.26717
R478 VTAIL.n309 VTAIL.n216 4.26717
R479 VTAIL.n280 VTAIL.n231 4.26717
R480 VTAIL.n261 VTAIL.n239 4.26717
R481 VTAIL.n203 VTAIL.n110 4.26717
R482 VTAIL.n174 VTAIL.n125 4.26717
R483 VTAIL.n155 VTAIL.n133 4.26717
R484 VTAIL.n365 VTAIL.n346 3.49141
R485 VTAIL.n386 VTAIL.n334 3.49141
R486 VTAIL.n412 VTAIL.n411 3.49141
R487 VTAIL.n47 VTAIL.n28 3.49141
R488 VTAIL.n68 VTAIL.n16 3.49141
R489 VTAIL.n94 VTAIL.n93 3.49141
R490 VTAIL.n306 VTAIL.n305 3.49141
R491 VTAIL.n281 VTAIL.n229 3.49141
R492 VTAIL.n260 VTAIL.n241 3.49141
R493 VTAIL.n200 VTAIL.n199 3.49141
R494 VTAIL.n175 VTAIL.n123 3.49141
R495 VTAIL.n154 VTAIL.n135 3.49141
R496 VTAIL.n362 VTAIL.n361 2.71565
R497 VTAIL.n390 VTAIL.n389 2.71565
R498 VTAIL.n408 VTAIL.n324 2.71565
R499 VTAIL.n44 VTAIL.n43 2.71565
R500 VTAIL.n72 VTAIL.n71 2.71565
R501 VTAIL.n90 VTAIL.n6 2.71565
R502 VTAIL.n302 VTAIL.n218 2.71565
R503 VTAIL.n285 VTAIL.n284 2.71565
R504 VTAIL.n257 VTAIL.n256 2.71565
R505 VTAIL.n196 VTAIL.n112 2.71565
R506 VTAIL.n179 VTAIL.n178 2.71565
R507 VTAIL.n151 VTAIL.n150 2.71565
R508 VTAIL.n358 VTAIL.n348 1.93989
R509 VTAIL.n394 VTAIL.n332 1.93989
R510 VTAIL.n407 VTAIL.n326 1.93989
R511 VTAIL.n40 VTAIL.n30 1.93989
R512 VTAIL.n76 VTAIL.n14 1.93989
R513 VTAIL.n89 VTAIL.n8 1.93989
R514 VTAIL.n301 VTAIL.n220 1.93989
R515 VTAIL.n288 VTAIL.n226 1.93989
R516 VTAIL.n253 VTAIL.n243 1.93989
R517 VTAIL.n195 VTAIL.n114 1.93989
R518 VTAIL.n182 VTAIL.n120 1.93989
R519 VTAIL.n147 VTAIL.n137 1.93989
R520 VTAIL.n357 VTAIL.n350 1.16414
R521 VTAIL.n395 VTAIL.n330 1.16414
R522 VTAIL.n404 VTAIL.n403 1.16414
R523 VTAIL.n39 VTAIL.n32 1.16414
R524 VTAIL.n77 VTAIL.n12 1.16414
R525 VTAIL.n86 VTAIL.n85 1.16414
R526 VTAIL.n298 VTAIL.n297 1.16414
R527 VTAIL.n289 VTAIL.n224 1.16414
R528 VTAIL.n252 VTAIL.n245 1.16414
R529 VTAIL.n192 VTAIL.n191 1.16414
R530 VTAIL.n183 VTAIL.n118 1.16414
R531 VTAIL.n146 VTAIL.n139 1.16414
R532 VTAIL.n317 VTAIL.n211 1.06516
R533 VTAIL VTAIL.n105 0.825931
R534 VTAIL.n354 VTAIL.n353 0.388379
R535 VTAIL.n399 VTAIL.n398 0.388379
R536 VTAIL.n400 VTAIL.n328 0.388379
R537 VTAIL.n36 VTAIL.n35 0.388379
R538 VTAIL.n81 VTAIL.n80 0.388379
R539 VTAIL.n82 VTAIL.n10 0.388379
R540 VTAIL.n294 VTAIL.n222 0.388379
R541 VTAIL.n293 VTAIL.n292 0.388379
R542 VTAIL.n249 VTAIL.n248 0.388379
R543 VTAIL.n188 VTAIL.n116 0.388379
R544 VTAIL.n187 VTAIL.n186 0.388379
R545 VTAIL.n143 VTAIL.n142 0.388379
R546 VTAIL VTAIL.n423 0.239724
R547 VTAIL.n356 VTAIL.n355 0.155672
R548 VTAIL.n356 VTAIL.n347 0.155672
R549 VTAIL.n363 VTAIL.n347 0.155672
R550 VTAIL.n364 VTAIL.n363 0.155672
R551 VTAIL.n364 VTAIL.n343 0.155672
R552 VTAIL.n371 VTAIL.n343 0.155672
R553 VTAIL.n372 VTAIL.n371 0.155672
R554 VTAIL.n372 VTAIL.n339 0.155672
R555 VTAIL.n379 VTAIL.n339 0.155672
R556 VTAIL.n380 VTAIL.n379 0.155672
R557 VTAIL.n380 VTAIL.n335 0.155672
R558 VTAIL.n387 VTAIL.n335 0.155672
R559 VTAIL.n388 VTAIL.n387 0.155672
R560 VTAIL.n388 VTAIL.n331 0.155672
R561 VTAIL.n396 VTAIL.n331 0.155672
R562 VTAIL.n397 VTAIL.n396 0.155672
R563 VTAIL.n397 VTAIL.n327 0.155672
R564 VTAIL.n405 VTAIL.n327 0.155672
R565 VTAIL.n406 VTAIL.n405 0.155672
R566 VTAIL.n406 VTAIL.n323 0.155672
R567 VTAIL.n413 VTAIL.n323 0.155672
R568 VTAIL.n414 VTAIL.n413 0.155672
R569 VTAIL.n414 VTAIL.n319 0.155672
R570 VTAIL.n421 VTAIL.n319 0.155672
R571 VTAIL.n38 VTAIL.n37 0.155672
R572 VTAIL.n38 VTAIL.n29 0.155672
R573 VTAIL.n45 VTAIL.n29 0.155672
R574 VTAIL.n46 VTAIL.n45 0.155672
R575 VTAIL.n46 VTAIL.n25 0.155672
R576 VTAIL.n53 VTAIL.n25 0.155672
R577 VTAIL.n54 VTAIL.n53 0.155672
R578 VTAIL.n54 VTAIL.n21 0.155672
R579 VTAIL.n61 VTAIL.n21 0.155672
R580 VTAIL.n62 VTAIL.n61 0.155672
R581 VTAIL.n62 VTAIL.n17 0.155672
R582 VTAIL.n69 VTAIL.n17 0.155672
R583 VTAIL.n70 VTAIL.n69 0.155672
R584 VTAIL.n70 VTAIL.n13 0.155672
R585 VTAIL.n78 VTAIL.n13 0.155672
R586 VTAIL.n79 VTAIL.n78 0.155672
R587 VTAIL.n79 VTAIL.n9 0.155672
R588 VTAIL.n87 VTAIL.n9 0.155672
R589 VTAIL.n88 VTAIL.n87 0.155672
R590 VTAIL.n88 VTAIL.n5 0.155672
R591 VTAIL.n95 VTAIL.n5 0.155672
R592 VTAIL.n96 VTAIL.n95 0.155672
R593 VTAIL.n96 VTAIL.n1 0.155672
R594 VTAIL.n103 VTAIL.n1 0.155672
R595 VTAIL.n315 VTAIL.n213 0.155672
R596 VTAIL.n308 VTAIL.n213 0.155672
R597 VTAIL.n308 VTAIL.n307 0.155672
R598 VTAIL.n307 VTAIL.n217 0.155672
R599 VTAIL.n300 VTAIL.n217 0.155672
R600 VTAIL.n300 VTAIL.n299 0.155672
R601 VTAIL.n299 VTAIL.n221 0.155672
R602 VTAIL.n291 VTAIL.n221 0.155672
R603 VTAIL.n291 VTAIL.n290 0.155672
R604 VTAIL.n290 VTAIL.n225 0.155672
R605 VTAIL.n283 VTAIL.n225 0.155672
R606 VTAIL.n283 VTAIL.n282 0.155672
R607 VTAIL.n282 VTAIL.n230 0.155672
R608 VTAIL.n275 VTAIL.n230 0.155672
R609 VTAIL.n275 VTAIL.n274 0.155672
R610 VTAIL.n274 VTAIL.n234 0.155672
R611 VTAIL.n267 VTAIL.n234 0.155672
R612 VTAIL.n267 VTAIL.n266 0.155672
R613 VTAIL.n266 VTAIL.n238 0.155672
R614 VTAIL.n259 VTAIL.n238 0.155672
R615 VTAIL.n259 VTAIL.n258 0.155672
R616 VTAIL.n258 VTAIL.n242 0.155672
R617 VTAIL.n251 VTAIL.n242 0.155672
R618 VTAIL.n251 VTAIL.n250 0.155672
R619 VTAIL.n209 VTAIL.n107 0.155672
R620 VTAIL.n202 VTAIL.n107 0.155672
R621 VTAIL.n202 VTAIL.n201 0.155672
R622 VTAIL.n201 VTAIL.n111 0.155672
R623 VTAIL.n194 VTAIL.n111 0.155672
R624 VTAIL.n194 VTAIL.n193 0.155672
R625 VTAIL.n193 VTAIL.n115 0.155672
R626 VTAIL.n185 VTAIL.n115 0.155672
R627 VTAIL.n185 VTAIL.n184 0.155672
R628 VTAIL.n184 VTAIL.n119 0.155672
R629 VTAIL.n177 VTAIL.n119 0.155672
R630 VTAIL.n177 VTAIL.n176 0.155672
R631 VTAIL.n176 VTAIL.n124 0.155672
R632 VTAIL.n169 VTAIL.n124 0.155672
R633 VTAIL.n169 VTAIL.n168 0.155672
R634 VTAIL.n168 VTAIL.n128 0.155672
R635 VTAIL.n161 VTAIL.n128 0.155672
R636 VTAIL.n161 VTAIL.n160 0.155672
R637 VTAIL.n160 VTAIL.n132 0.155672
R638 VTAIL.n153 VTAIL.n132 0.155672
R639 VTAIL.n153 VTAIL.n152 0.155672
R640 VTAIL.n152 VTAIL.n136 0.155672
R641 VTAIL.n145 VTAIL.n136 0.155672
R642 VTAIL.n145 VTAIL.n144 0.155672
R643 VDD2.n205 VDD2.n105 289.615
R644 VDD2.n100 VDD2.n0 289.615
R645 VDD2.n206 VDD2.n205 185
R646 VDD2.n204 VDD2.n203 185
R647 VDD2.n109 VDD2.n108 185
R648 VDD2.n198 VDD2.n197 185
R649 VDD2.n196 VDD2.n195 185
R650 VDD2.n113 VDD2.n112 185
R651 VDD2.n190 VDD2.n189 185
R652 VDD2.n188 VDD2.n187 185
R653 VDD2.n186 VDD2.n116 185
R654 VDD2.n120 VDD2.n117 185
R655 VDD2.n181 VDD2.n180 185
R656 VDD2.n179 VDD2.n178 185
R657 VDD2.n122 VDD2.n121 185
R658 VDD2.n173 VDD2.n172 185
R659 VDD2.n171 VDD2.n170 185
R660 VDD2.n126 VDD2.n125 185
R661 VDD2.n165 VDD2.n164 185
R662 VDD2.n163 VDD2.n162 185
R663 VDD2.n130 VDD2.n129 185
R664 VDD2.n157 VDD2.n156 185
R665 VDD2.n155 VDD2.n154 185
R666 VDD2.n134 VDD2.n133 185
R667 VDD2.n149 VDD2.n148 185
R668 VDD2.n147 VDD2.n146 185
R669 VDD2.n138 VDD2.n137 185
R670 VDD2.n141 VDD2.n140 185
R671 VDD2.n35 VDD2.n34 185
R672 VDD2.n32 VDD2.n31 185
R673 VDD2.n41 VDD2.n40 185
R674 VDD2.n43 VDD2.n42 185
R675 VDD2.n28 VDD2.n27 185
R676 VDD2.n49 VDD2.n48 185
R677 VDD2.n51 VDD2.n50 185
R678 VDD2.n24 VDD2.n23 185
R679 VDD2.n57 VDD2.n56 185
R680 VDD2.n59 VDD2.n58 185
R681 VDD2.n20 VDD2.n19 185
R682 VDD2.n65 VDD2.n64 185
R683 VDD2.n67 VDD2.n66 185
R684 VDD2.n16 VDD2.n15 185
R685 VDD2.n73 VDD2.n72 185
R686 VDD2.n76 VDD2.n75 185
R687 VDD2.n74 VDD2.n12 185
R688 VDD2.n81 VDD2.n11 185
R689 VDD2.n83 VDD2.n82 185
R690 VDD2.n85 VDD2.n84 185
R691 VDD2.n8 VDD2.n7 185
R692 VDD2.n91 VDD2.n90 185
R693 VDD2.n93 VDD2.n92 185
R694 VDD2.n4 VDD2.n3 185
R695 VDD2.n99 VDD2.n98 185
R696 VDD2.n101 VDD2.n100 185
R697 VDD2.t1 VDD2.n139 147.659
R698 VDD2.t0 VDD2.n33 147.659
R699 VDD2.n205 VDD2.n204 104.615
R700 VDD2.n204 VDD2.n108 104.615
R701 VDD2.n197 VDD2.n108 104.615
R702 VDD2.n197 VDD2.n196 104.615
R703 VDD2.n196 VDD2.n112 104.615
R704 VDD2.n189 VDD2.n112 104.615
R705 VDD2.n189 VDD2.n188 104.615
R706 VDD2.n188 VDD2.n116 104.615
R707 VDD2.n120 VDD2.n116 104.615
R708 VDD2.n180 VDD2.n120 104.615
R709 VDD2.n180 VDD2.n179 104.615
R710 VDD2.n179 VDD2.n121 104.615
R711 VDD2.n172 VDD2.n121 104.615
R712 VDD2.n172 VDD2.n171 104.615
R713 VDD2.n171 VDD2.n125 104.615
R714 VDD2.n164 VDD2.n125 104.615
R715 VDD2.n164 VDD2.n163 104.615
R716 VDD2.n163 VDD2.n129 104.615
R717 VDD2.n156 VDD2.n129 104.615
R718 VDD2.n156 VDD2.n155 104.615
R719 VDD2.n155 VDD2.n133 104.615
R720 VDD2.n148 VDD2.n133 104.615
R721 VDD2.n148 VDD2.n147 104.615
R722 VDD2.n147 VDD2.n137 104.615
R723 VDD2.n140 VDD2.n137 104.615
R724 VDD2.n34 VDD2.n31 104.615
R725 VDD2.n41 VDD2.n31 104.615
R726 VDD2.n42 VDD2.n41 104.615
R727 VDD2.n42 VDD2.n27 104.615
R728 VDD2.n49 VDD2.n27 104.615
R729 VDD2.n50 VDD2.n49 104.615
R730 VDD2.n50 VDD2.n23 104.615
R731 VDD2.n57 VDD2.n23 104.615
R732 VDD2.n58 VDD2.n57 104.615
R733 VDD2.n58 VDD2.n19 104.615
R734 VDD2.n65 VDD2.n19 104.615
R735 VDD2.n66 VDD2.n65 104.615
R736 VDD2.n66 VDD2.n15 104.615
R737 VDD2.n73 VDD2.n15 104.615
R738 VDD2.n75 VDD2.n73 104.615
R739 VDD2.n75 VDD2.n74 104.615
R740 VDD2.n74 VDD2.n11 104.615
R741 VDD2.n83 VDD2.n11 104.615
R742 VDD2.n84 VDD2.n83 104.615
R743 VDD2.n84 VDD2.n7 104.615
R744 VDD2.n91 VDD2.n7 104.615
R745 VDD2.n92 VDD2.n91 104.615
R746 VDD2.n92 VDD2.n3 104.615
R747 VDD2.n99 VDD2.n3 104.615
R748 VDD2.n100 VDD2.n99 104.615
R749 VDD2.n210 VDD2.n104 92.6829
R750 VDD2.n140 VDD2.t1 52.3082
R751 VDD2.n34 VDD2.t0 52.3082
R752 VDD2.n210 VDD2.n209 50.2217
R753 VDD2.n141 VDD2.n139 15.6677
R754 VDD2.n35 VDD2.n33 15.6677
R755 VDD2.n187 VDD2.n186 13.1884
R756 VDD2.n82 VDD2.n81 13.1884
R757 VDD2.n190 VDD2.n115 12.8005
R758 VDD2.n185 VDD2.n117 12.8005
R759 VDD2.n142 VDD2.n138 12.8005
R760 VDD2.n36 VDD2.n32 12.8005
R761 VDD2.n80 VDD2.n12 12.8005
R762 VDD2.n85 VDD2.n10 12.8005
R763 VDD2.n191 VDD2.n113 12.0247
R764 VDD2.n182 VDD2.n181 12.0247
R765 VDD2.n146 VDD2.n145 12.0247
R766 VDD2.n40 VDD2.n39 12.0247
R767 VDD2.n77 VDD2.n76 12.0247
R768 VDD2.n86 VDD2.n8 12.0247
R769 VDD2.n195 VDD2.n194 11.249
R770 VDD2.n178 VDD2.n119 11.249
R771 VDD2.n149 VDD2.n136 11.249
R772 VDD2.n43 VDD2.n30 11.249
R773 VDD2.n72 VDD2.n14 11.249
R774 VDD2.n90 VDD2.n89 11.249
R775 VDD2.n198 VDD2.n111 10.4732
R776 VDD2.n177 VDD2.n122 10.4732
R777 VDD2.n150 VDD2.n134 10.4732
R778 VDD2.n44 VDD2.n28 10.4732
R779 VDD2.n71 VDD2.n16 10.4732
R780 VDD2.n93 VDD2.n6 10.4732
R781 VDD2.n199 VDD2.n109 9.69747
R782 VDD2.n174 VDD2.n173 9.69747
R783 VDD2.n154 VDD2.n153 9.69747
R784 VDD2.n48 VDD2.n47 9.69747
R785 VDD2.n68 VDD2.n67 9.69747
R786 VDD2.n94 VDD2.n4 9.69747
R787 VDD2.n209 VDD2.n208 9.45567
R788 VDD2.n104 VDD2.n103 9.45567
R789 VDD2.n167 VDD2.n166 9.3005
R790 VDD2.n169 VDD2.n168 9.3005
R791 VDD2.n124 VDD2.n123 9.3005
R792 VDD2.n175 VDD2.n174 9.3005
R793 VDD2.n177 VDD2.n176 9.3005
R794 VDD2.n119 VDD2.n118 9.3005
R795 VDD2.n183 VDD2.n182 9.3005
R796 VDD2.n185 VDD2.n184 9.3005
R797 VDD2.n208 VDD2.n207 9.3005
R798 VDD2.n107 VDD2.n106 9.3005
R799 VDD2.n202 VDD2.n201 9.3005
R800 VDD2.n200 VDD2.n199 9.3005
R801 VDD2.n111 VDD2.n110 9.3005
R802 VDD2.n194 VDD2.n193 9.3005
R803 VDD2.n192 VDD2.n191 9.3005
R804 VDD2.n115 VDD2.n114 9.3005
R805 VDD2.n128 VDD2.n127 9.3005
R806 VDD2.n161 VDD2.n160 9.3005
R807 VDD2.n159 VDD2.n158 9.3005
R808 VDD2.n132 VDD2.n131 9.3005
R809 VDD2.n153 VDD2.n152 9.3005
R810 VDD2.n151 VDD2.n150 9.3005
R811 VDD2.n136 VDD2.n135 9.3005
R812 VDD2.n145 VDD2.n144 9.3005
R813 VDD2.n143 VDD2.n142 9.3005
R814 VDD2.n2 VDD2.n1 9.3005
R815 VDD2.n97 VDD2.n96 9.3005
R816 VDD2.n95 VDD2.n94 9.3005
R817 VDD2.n6 VDD2.n5 9.3005
R818 VDD2.n89 VDD2.n88 9.3005
R819 VDD2.n87 VDD2.n86 9.3005
R820 VDD2.n10 VDD2.n9 9.3005
R821 VDD2.n55 VDD2.n54 9.3005
R822 VDD2.n53 VDD2.n52 9.3005
R823 VDD2.n26 VDD2.n25 9.3005
R824 VDD2.n47 VDD2.n46 9.3005
R825 VDD2.n45 VDD2.n44 9.3005
R826 VDD2.n30 VDD2.n29 9.3005
R827 VDD2.n39 VDD2.n38 9.3005
R828 VDD2.n37 VDD2.n36 9.3005
R829 VDD2.n22 VDD2.n21 9.3005
R830 VDD2.n61 VDD2.n60 9.3005
R831 VDD2.n63 VDD2.n62 9.3005
R832 VDD2.n18 VDD2.n17 9.3005
R833 VDD2.n69 VDD2.n68 9.3005
R834 VDD2.n71 VDD2.n70 9.3005
R835 VDD2.n14 VDD2.n13 9.3005
R836 VDD2.n78 VDD2.n77 9.3005
R837 VDD2.n80 VDD2.n79 9.3005
R838 VDD2.n103 VDD2.n102 9.3005
R839 VDD2.n203 VDD2.n202 8.92171
R840 VDD2.n170 VDD2.n124 8.92171
R841 VDD2.n157 VDD2.n132 8.92171
R842 VDD2.n51 VDD2.n26 8.92171
R843 VDD2.n64 VDD2.n18 8.92171
R844 VDD2.n98 VDD2.n97 8.92171
R845 VDD2.n206 VDD2.n107 8.14595
R846 VDD2.n169 VDD2.n126 8.14595
R847 VDD2.n158 VDD2.n130 8.14595
R848 VDD2.n52 VDD2.n24 8.14595
R849 VDD2.n63 VDD2.n20 8.14595
R850 VDD2.n101 VDD2.n2 8.14595
R851 VDD2.n207 VDD2.n105 7.3702
R852 VDD2.n166 VDD2.n165 7.3702
R853 VDD2.n162 VDD2.n161 7.3702
R854 VDD2.n56 VDD2.n55 7.3702
R855 VDD2.n60 VDD2.n59 7.3702
R856 VDD2.n102 VDD2.n0 7.3702
R857 VDD2.n209 VDD2.n105 6.59444
R858 VDD2.n165 VDD2.n128 6.59444
R859 VDD2.n162 VDD2.n128 6.59444
R860 VDD2.n56 VDD2.n22 6.59444
R861 VDD2.n59 VDD2.n22 6.59444
R862 VDD2.n104 VDD2.n0 6.59444
R863 VDD2.n207 VDD2.n206 5.81868
R864 VDD2.n166 VDD2.n126 5.81868
R865 VDD2.n161 VDD2.n130 5.81868
R866 VDD2.n55 VDD2.n24 5.81868
R867 VDD2.n60 VDD2.n20 5.81868
R868 VDD2.n102 VDD2.n101 5.81868
R869 VDD2.n203 VDD2.n107 5.04292
R870 VDD2.n170 VDD2.n169 5.04292
R871 VDD2.n158 VDD2.n157 5.04292
R872 VDD2.n52 VDD2.n51 5.04292
R873 VDD2.n64 VDD2.n63 5.04292
R874 VDD2.n98 VDD2.n2 5.04292
R875 VDD2.n143 VDD2.n139 4.38563
R876 VDD2.n37 VDD2.n33 4.38563
R877 VDD2.n202 VDD2.n109 4.26717
R878 VDD2.n173 VDD2.n124 4.26717
R879 VDD2.n154 VDD2.n132 4.26717
R880 VDD2.n48 VDD2.n26 4.26717
R881 VDD2.n67 VDD2.n18 4.26717
R882 VDD2.n97 VDD2.n4 4.26717
R883 VDD2.n199 VDD2.n198 3.49141
R884 VDD2.n174 VDD2.n122 3.49141
R885 VDD2.n153 VDD2.n134 3.49141
R886 VDD2.n47 VDD2.n28 3.49141
R887 VDD2.n68 VDD2.n16 3.49141
R888 VDD2.n94 VDD2.n93 3.49141
R889 VDD2.n195 VDD2.n111 2.71565
R890 VDD2.n178 VDD2.n177 2.71565
R891 VDD2.n150 VDD2.n149 2.71565
R892 VDD2.n44 VDD2.n43 2.71565
R893 VDD2.n72 VDD2.n71 2.71565
R894 VDD2.n90 VDD2.n6 2.71565
R895 VDD2.n194 VDD2.n113 1.93989
R896 VDD2.n181 VDD2.n119 1.93989
R897 VDD2.n146 VDD2.n136 1.93989
R898 VDD2.n40 VDD2.n30 1.93989
R899 VDD2.n76 VDD2.n14 1.93989
R900 VDD2.n89 VDD2.n8 1.93989
R901 VDD2.n191 VDD2.n190 1.16414
R902 VDD2.n182 VDD2.n117 1.16414
R903 VDD2.n145 VDD2.n138 1.16414
R904 VDD2.n39 VDD2.n32 1.16414
R905 VDD2.n77 VDD2.n12 1.16414
R906 VDD2.n86 VDD2.n85 1.16414
R907 VDD2.n187 VDD2.n115 0.388379
R908 VDD2.n186 VDD2.n185 0.388379
R909 VDD2.n142 VDD2.n141 0.388379
R910 VDD2.n36 VDD2.n35 0.388379
R911 VDD2.n81 VDD2.n80 0.388379
R912 VDD2.n82 VDD2.n10 0.388379
R913 VDD2 VDD2.n210 0.356103
R914 VDD2.n208 VDD2.n106 0.155672
R915 VDD2.n201 VDD2.n106 0.155672
R916 VDD2.n201 VDD2.n200 0.155672
R917 VDD2.n200 VDD2.n110 0.155672
R918 VDD2.n193 VDD2.n110 0.155672
R919 VDD2.n193 VDD2.n192 0.155672
R920 VDD2.n192 VDD2.n114 0.155672
R921 VDD2.n184 VDD2.n114 0.155672
R922 VDD2.n184 VDD2.n183 0.155672
R923 VDD2.n183 VDD2.n118 0.155672
R924 VDD2.n176 VDD2.n118 0.155672
R925 VDD2.n176 VDD2.n175 0.155672
R926 VDD2.n175 VDD2.n123 0.155672
R927 VDD2.n168 VDD2.n123 0.155672
R928 VDD2.n168 VDD2.n167 0.155672
R929 VDD2.n167 VDD2.n127 0.155672
R930 VDD2.n160 VDD2.n127 0.155672
R931 VDD2.n160 VDD2.n159 0.155672
R932 VDD2.n159 VDD2.n131 0.155672
R933 VDD2.n152 VDD2.n131 0.155672
R934 VDD2.n152 VDD2.n151 0.155672
R935 VDD2.n151 VDD2.n135 0.155672
R936 VDD2.n144 VDD2.n135 0.155672
R937 VDD2.n144 VDD2.n143 0.155672
R938 VDD2.n38 VDD2.n37 0.155672
R939 VDD2.n38 VDD2.n29 0.155672
R940 VDD2.n45 VDD2.n29 0.155672
R941 VDD2.n46 VDD2.n45 0.155672
R942 VDD2.n46 VDD2.n25 0.155672
R943 VDD2.n53 VDD2.n25 0.155672
R944 VDD2.n54 VDD2.n53 0.155672
R945 VDD2.n54 VDD2.n21 0.155672
R946 VDD2.n61 VDD2.n21 0.155672
R947 VDD2.n62 VDD2.n61 0.155672
R948 VDD2.n62 VDD2.n17 0.155672
R949 VDD2.n69 VDD2.n17 0.155672
R950 VDD2.n70 VDD2.n69 0.155672
R951 VDD2.n70 VDD2.n13 0.155672
R952 VDD2.n78 VDD2.n13 0.155672
R953 VDD2.n79 VDD2.n78 0.155672
R954 VDD2.n79 VDD2.n9 0.155672
R955 VDD2.n87 VDD2.n9 0.155672
R956 VDD2.n88 VDD2.n87 0.155672
R957 VDD2.n88 VDD2.n5 0.155672
R958 VDD2.n95 VDD2.n5 0.155672
R959 VDD2.n96 VDD2.n95 0.155672
R960 VDD2.n96 VDD2.n1 0.155672
R961 VDD2.n103 VDD2.n1 0.155672
R962 B.n432 B.t2 640.038
R963 B.n589 B.t13 640.038
R964 B.n104 B.t10 640.038
R965 B.n101 B.t6 640.038
R966 B.n810 B.n809 585
R967 B.n369 B.n100 585
R968 B.n368 B.n367 585
R969 B.n366 B.n365 585
R970 B.n364 B.n363 585
R971 B.n362 B.n361 585
R972 B.n360 B.n359 585
R973 B.n358 B.n357 585
R974 B.n356 B.n355 585
R975 B.n354 B.n353 585
R976 B.n352 B.n351 585
R977 B.n350 B.n349 585
R978 B.n348 B.n347 585
R979 B.n346 B.n345 585
R980 B.n344 B.n343 585
R981 B.n342 B.n341 585
R982 B.n340 B.n339 585
R983 B.n338 B.n337 585
R984 B.n336 B.n335 585
R985 B.n334 B.n333 585
R986 B.n332 B.n331 585
R987 B.n330 B.n329 585
R988 B.n328 B.n327 585
R989 B.n326 B.n325 585
R990 B.n324 B.n323 585
R991 B.n322 B.n321 585
R992 B.n320 B.n319 585
R993 B.n318 B.n317 585
R994 B.n316 B.n315 585
R995 B.n314 B.n313 585
R996 B.n312 B.n311 585
R997 B.n310 B.n309 585
R998 B.n308 B.n307 585
R999 B.n306 B.n305 585
R1000 B.n304 B.n303 585
R1001 B.n302 B.n301 585
R1002 B.n300 B.n299 585
R1003 B.n298 B.n297 585
R1004 B.n296 B.n295 585
R1005 B.n294 B.n293 585
R1006 B.n292 B.n291 585
R1007 B.n290 B.n289 585
R1008 B.n288 B.n287 585
R1009 B.n286 B.n285 585
R1010 B.n284 B.n283 585
R1011 B.n282 B.n281 585
R1012 B.n280 B.n279 585
R1013 B.n278 B.n277 585
R1014 B.n276 B.n275 585
R1015 B.n274 B.n273 585
R1016 B.n272 B.n271 585
R1017 B.n270 B.n269 585
R1018 B.n268 B.n267 585
R1019 B.n266 B.n265 585
R1020 B.n264 B.n263 585
R1021 B.n262 B.n261 585
R1022 B.n260 B.n259 585
R1023 B.n258 B.n257 585
R1024 B.n256 B.n255 585
R1025 B.n254 B.n253 585
R1026 B.n252 B.n251 585
R1027 B.n250 B.n249 585
R1028 B.n248 B.n247 585
R1029 B.n246 B.n245 585
R1030 B.n244 B.n243 585
R1031 B.n242 B.n241 585
R1032 B.n240 B.n239 585
R1033 B.n238 B.n237 585
R1034 B.n236 B.n235 585
R1035 B.n234 B.n233 585
R1036 B.n232 B.n231 585
R1037 B.n230 B.n229 585
R1038 B.n228 B.n227 585
R1039 B.n226 B.n225 585
R1040 B.n224 B.n223 585
R1041 B.n222 B.n221 585
R1042 B.n220 B.n219 585
R1043 B.n218 B.n217 585
R1044 B.n216 B.n215 585
R1045 B.n214 B.n213 585
R1046 B.n212 B.n211 585
R1047 B.n210 B.n209 585
R1048 B.n208 B.n207 585
R1049 B.n206 B.n205 585
R1050 B.n204 B.n203 585
R1051 B.n202 B.n201 585
R1052 B.n200 B.n199 585
R1053 B.n198 B.n197 585
R1054 B.n196 B.n195 585
R1055 B.n194 B.n193 585
R1056 B.n192 B.n191 585
R1057 B.n190 B.n189 585
R1058 B.n188 B.n187 585
R1059 B.n186 B.n185 585
R1060 B.n184 B.n183 585
R1061 B.n182 B.n181 585
R1062 B.n180 B.n179 585
R1063 B.n178 B.n177 585
R1064 B.n176 B.n175 585
R1065 B.n174 B.n173 585
R1066 B.n172 B.n171 585
R1067 B.n170 B.n169 585
R1068 B.n168 B.n167 585
R1069 B.n166 B.n165 585
R1070 B.n164 B.n163 585
R1071 B.n162 B.n161 585
R1072 B.n160 B.n159 585
R1073 B.n158 B.n157 585
R1074 B.n156 B.n155 585
R1075 B.n154 B.n153 585
R1076 B.n152 B.n151 585
R1077 B.n150 B.n149 585
R1078 B.n148 B.n147 585
R1079 B.n146 B.n145 585
R1080 B.n144 B.n143 585
R1081 B.n142 B.n141 585
R1082 B.n140 B.n139 585
R1083 B.n138 B.n137 585
R1084 B.n136 B.n135 585
R1085 B.n134 B.n133 585
R1086 B.n132 B.n131 585
R1087 B.n130 B.n129 585
R1088 B.n128 B.n127 585
R1089 B.n126 B.n125 585
R1090 B.n124 B.n123 585
R1091 B.n122 B.n121 585
R1092 B.n120 B.n119 585
R1093 B.n118 B.n117 585
R1094 B.n116 B.n115 585
R1095 B.n114 B.n113 585
R1096 B.n112 B.n111 585
R1097 B.n110 B.n109 585
R1098 B.n108 B.n107 585
R1099 B.n32 B.n31 585
R1100 B.n808 B.n33 585
R1101 B.n813 B.n33 585
R1102 B.n807 B.n806 585
R1103 B.n806 B.n29 585
R1104 B.n805 B.n28 585
R1105 B.n819 B.n28 585
R1106 B.n804 B.n27 585
R1107 B.n820 B.n27 585
R1108 B.n803 B.n26 585
R1109 B.n821 B.n26 585
R1110 B.n802 B.n801 585
R1111 B.n801 B.n25 585
R1112 B.n800 B.n21 585
R1113 B.n827 B.n21 585
R1114 B.n799 B.n20 585
R1115 B.n828 B.n20 585
R1116 B.n798 B.n19 585
R1117 B.n829 B.n19 585
R1118 B.n797 B.n796 585
R1119 B.n796 B.n15 585
R1120 B.n795 B.n14 585
R1121 B.n835 B.n14 585
R1122 B.n794 B.n13 585
R1123 B.n836 B.n13 585
R1124 B.n793 B.n12 585
R1125 B.n837 B.n12 585
R1126 B.n792 B.n791 585
R1127 B.n791 B.n8 585
R1128 B.n790 B.n7 585
R1129 B.n843 B.n7 585
R1130 B.n789 B.n6 585
R1131 B.n844 B.n6 585
R1132 B.n788 B.n5 585
R1133 B.n845 B.n5 585
R1134 B.n787 B.n786 585
R1135 B.n786 B.n4 585
R1136 B.n785 B.n370 585
R1137 B.n785 B.n784 585
R1138 B.n775 B.n371 585
R1139 B.n372 B.n371 585
R1140 B.n777 B.n776 585
R1141 B.n778 B.n777 585
R1142 B.n774 B.n377 585
R1143 B.n377 B.n376 585
R1144 B.n773 B.n772 585
R1145 B.n772 B.n771 585
R1146 B.n379 B.n378 585
R1147 B.n380 B.n379 585
R1148 B.n764 B.n763 585
R1149 B.n765 B.n764 585
R1150 B.n762 B.n385 585
R1151 B.n385 B.n384 585
R1152 B.n761 B.n760 585
R1153 B.n760 B.n759 585
R1154 B.n387 B.n386 585
R1155 B.n752 B.n387 585
R1156 B.n751 B.n750 585
R1157 B.n753 B.n751 585
R1158 B.n749 B.n392 585
R1159 B.n392 B.n391 585
R1160 B.n748 B.n747 585
R1161 B.n747 B.n746 585
R1162 B.n394 B.n393 585
R1163 B.n395 B.n394 585
R1164 B.n739 B.n738 585
R1165 B.n740 B.n739 585
R1166 B.n398 B.n397 585
R1167 B.n471 B.n469 585
R1168 B.n472 B.n468 585
R1169 B.n472 B.n399 585
R1170 B.n475 B.n474 585
R1171 B.n476 B.n467 585
R1172 B.n478 B.n477 585
R1173 B.n480 B.n466 585
R1174 B.n483 B.n482 585
R1175 B.n484 B.n465 585
R1176 B.n486 B.n485 585
R1177 B.n488 B.n464 585
R1178 B.n491 B.n490 585
R1179 B.n492 B.n463 585
R1180 B.n494 B.n493 585
R1181 B.n496 B.n462 585
R1182 B.n499 B.n498 585
R1183 B.n500 B.n461 585
R1184 B.n502 B.n501 585
R1185 B.n504 B.n460 585
R1186 B.n507 B.n506 585
R1187 B.n508 B.n459 585
R1188 B.n510 B.n509 585
R1189 B.n512 B.n458 585
R1190 B.n515 B.n514 585
R1191 B.n516 B.n457 585
R1192 B.n518 B.n517 585
R1193 B.n520 B.n456 585
R1194 B.n523 B.n522 585
R1195 B.n524 B.n455 585
R1196 B.n526 B.n525 585
R1197 B.n528 B.n454 585
R1198 B.n531 B.n530 585
R1199 B.n532 B.n453 585
R1200 B.n534 B.n533 585
R1201 B.n536 B.n452 585
R1202 B.n539 B.n538 585
R1203 B.n540 B.n451 585
R1204 B.n542 B.n541 585
R1205 B.n544 B.n450 585
R1206 B.n547 B.n546 585
R1207 B.n548 B.n449 585
R1208 B.n550 B.n549 585
R1209 B.n552 B.n448 585
R1210 B.n555 B.n554 585
R1211 B.n556 B.n447 585
R1212 B.n558 B.n557 585
R1213 B.n560 B.n446 585
R1214 B.n563 B.n562 585
R1215 B.n564 B.n445 585
R1216 B.n566 B.n565 585
R1217 B.n568 B.n444 585
R1218 B.n571 B.n570 585
R1219 B.n572 B.n443 585
R1220 B.n574 B.n573 585
R1221 B.n576 B.n442 585
R1222 B.n579 B.n578 585
R1223 B.n580 B.n441 585
R1224 B.n582 B.n581 585
R1225 B.n584 B.n440 585
R1226 B.n587 B.n586 585
R1227 B.n588 B.n439 585
R1228 B.n593 B.n592 585
R1229 B.n595 B.n438 585
R1230 B.n598 B.n597 585
R1231 B.n599 B.n437 585
R1232 B.n601 B.n600 585
R1233 B.n603 B.n436 585
R1234 B.n606 B.n605 585
R1235 B.n607 B.n435 585
R1236 B.n609 B.n608 585
R1237 B.n611 B.n434 585
R1238 B.n614 B.n613 585
R1239 B.n616 B.n431 585
R1240 B.n618 B.n617 585
R1241 B.n620 B.n430 585
R1242 B.n623 B.n622 585
R1243 B.n624 B.n429 585
R1244 B.n626 B.n625 585
R1245 B.n628 B.n428 585
R1246 B.n631 B.n630 585
R1247 B.n632 B.n427 585
R1248 B.n634 B.n633 585
R1249 B.n636 B.n426 585
R1250 B.n639 B.n638 585
R1251 B.n640 B.n425 585
R1252 B.n642 B.n641 585
R1253 B.n644 B.n424 585
R1254 B.n647 B.n646 585
R1255 B.n648 B.n423 585
R1256 B.n650 B.n649 585
R1257 B.n652 B.n422 585
R1258 B.n655 B.n654 585
R1259 B.n656 B.n421 585
R1260 B.n658 B.n657 585
R1261 B.n660 B.n420 585
R1262 B.n663 B.n662 585
R1263 B.n664 B.n419 585
R1264 B.n666 B.n665 585
R1265 B.n668 B.n418 585
R1266 B.n671 B.n670 585
R1267 B.n672 B.n417 585
R1268 B.n674 B.n673 585
R1269 B.n676 B.n416 585
R1270 B.n679 B.n678 585
R1271 B.n680 B.n415 585
R1272 B.n682 B.n681 585
R1273 B.n684 B.n414 585
R1274 B.n687 B.n686 585
R1275 B.n688 B.n413 585
R1276 B.n690 B.n689 585
R1277 B.n692 B.n412 585
R1278 B.n695 B.n694 585
R1279 B.n696 B.n411 585
R1280 B.n698 B.n697 585
R1281 B.n700 B.n410 585
R1282 B.n703 B.n702 585
R1283 B.n704 B.n409 585
R1284 B.n706 B.n705 585
R1285 B.n708 B.n408 585
R1286 B.n711 B.n710 585
R1287 B.n712 B.n407 585
R1288 B.n714 B.n713 585
R1289 B.n716 B.n406 585
R1290 B.n719 B.n718 585
R1291 B.n720 B.n405 585
R1292 B.n722 B.n721 585
R1293 B.n724 B.n404 585
R1294 B.n727 B.n726 585
R1295 B.n728 B.n403 585
R1296 B.n730 B.n729 585
R1297 B.n732 B.n402 585
R1298 B.n733 B.n401 585
R1299 B.n736 B.n735 585
R1300 B.n737 B.n400 585
R1301 B.n400 B.n399 585
R1302 B.n742 B.n741 585
R1303 B.n741 B.n740 585
R1304 B.n743 B.n396 585
R1305 B.n396 B.n395 585
R1306 B.n745 B.n744 585
R1307 B.n746 B.n745 585
R1308 B.n390 B.n389 585
R1309 B.n391 B.n390 585
R1310 B.n755 B.n754 585
R1311 B.n754 B.n753 585
R1312 B.n756 B.n388 585
R1313 B.n752 B.n388 585
R1314 B.n758 B.n757 585
R1315 B.n759 B.n758 585
R1316 B.n383 B.n382 585
R1317 B.n384 B.n383 585
R1318 B.n767 B.n766 585
R1319 B.n766 B.n765 585
R1320 B.n768 B.n381 585
R1321 B.n381 B.n380 585
R1322 B.n770 B.n769 585
R1323 B.n771 B.n770 585
R1324 B.n375 B.n374 585
R1325 B.n376 B.n375 585
R1326 B.n780 B.n779 585
R1327 B.n779 B.n778 585
R1328 B.n781 B.n373 585
R1329 B.n373 B.n372 585
R1330 B.n783 B.n782 585
R1331 B.n784 B.n783 585
R1332 B.n2 B.n0 585
R1333 B.n4 B.n2 585
R1334 B.n3 B.n1 585
R1335 B.n844 B.n3 585
R1336 B.n842 B.n841 585
R1337 B.n843 B.n842 585
R1338 B.n840 B.n9 585
R1339 B.n9 B.n8 585
R1340 B.n839 B.n838 585
R1341 B.n838 B.n837 585
R1342 B.n11 B.n10 585
R1343 B.n836 B.n11 585
R1344 B.n834 B.n833 585
R1345 B.n835 B.n834 585
R1346 B.n832 B.n16 585
R1347 B.n16 B.n15 585
R1348 B.n831 B.n830 585
R1349 B.n830 B.n829 585
R1350 B.n18 B.n17 585
R1351 B.n828 B.n18 585
R1352 B.n826 B.n825 585
R1353 B.n827 B.n826 585
R1354 B.n824 B.n22 585
R1355 B.n25 B.n22 585
R1356 B.n823 B.n822 585
R1357 B.n822 B.n821 585
R1358 B.n24 B.n23 585
R1359 B.n820 B.n24 585
R1360 B.n818 B.n817 585
R1361 B.n819 B.n818 585
R1362 B.n816 B.n30 585
R1363 B.n30 B.n29 585
R1364 B.n815 B.n814 585
R1365 B.n814 B.n813 585
R1366 B.n847 B.n846 585
R1367 B.n846 B.n845 585
R1368 B.n741 B.n398 559.769
R1369 B.n814 B.n32 559.769
R1370 B.n739 B.n400 559.769
R1371 B.n810 B.n33 559.769
R1372 B.n432 B.t5 430.356
R1373 B.n589 B.t15 430.356
R1374 B.n104 B.t11 430.356
R1375 B.n101 B.t8 430.356
R1376 B.n433 B.t4 403.592
R1377 B.n102 B.t9 403.592
R1378 B.n590 B.t14 403.592
R1379 B.n105 B.t12 403.592
R1380 B.n812 B.n811 256.663
R1381 B.n812 B.n99 256.663
R1382 B.n812 B.n98 256.663
R1383 B.n812 B.n97 256.663
R1384 B.n812 B.n96 256.663
R1385 B.n812 B.n95 256.663
R1386 B.n812 B.n94 256.663
R1387 B.n812 B.n93 256.663
R1388 B.n812 B.n92 256.663
R1389 B.n812 B.n91 256.663
R1390 B.n812 B.n90 256.663
R1391 B.n812 B.n89 256.663
R1392 B.n812 B.n88 256.663
R1393 B.n812 B.n87 256.663
R1394 B.n812 B.n86 256.663
R1395 B.n812 B.n85 256.663
R1396 B.n812 B.n84 256.663
R1397 B.n812 B.n83 256.663
R1398 B.n812 B.n82 256.663
R1399 B.n812 B.n81 256.663
R1400 B.n812 B.n80 256.663
R1401 B.n812 B.n79 256.663
R1402 B.n812 B.n78 256.663
R1403 B.n812 B.n77 256.663
R1404 B.n812 B.n76 256.663
R1405 B.n812 B.n75 256.663
R1406 B.n812 B.n74 256.663
R1407 B.n812 B.n73 256.663
R1408 B.n812 B.n72 256.663
R1409 B.n812 B.n71 256.663
R1410 B.n812 B.n70 256.663
R1411 B.n812 B.n69 256.663
R1412 B.n812 B.n68 256.663
R1413 B.n812 B.n67 256.663
R1414 B.n812 B.n66 256.663
R1415 B.n812 B.n65 256.663
R1416 B.n812 B.n64 256.663
R1417 B.n812 B.n63 256.663
R1418 B.n812 B.n62 256.663
R1419 B.n812 B.n61 256.663
R1420 B.n812 B.n60 256.663
R1421 B.n812 B.n59 256.663
R1422 B.n812 B.n58 256.663
R1423 B.n812 B.n57 256.663
R1424 B.n812 B.n56 256.663
R1425 B.n812 B.n55 256.663
R1426 B.n812 B.n54 256.663
R1427 B.n812 B.n53 256.663
R1428 B.n812 B.n52 256.663
R1429 B.n812 B.n51 256.663
R1430 B.n812 B.n50 256.663
R1431 B.n812 B.n49 256.663
R1432 B.n812 B.n48 256.663
R1433 B.n812 B.n47 256.663
R1434 B.n812 B.n46 256.663
R1435 B.n812 B.n45 256.663
R1436 B.n812 B.n44 256.663
R1437 B.n812 B.n43 256.663
R1438 B.n812 B.n42 256.663
R1439 B.n812 B.n41 256.663
R1440 B.n812 B.n40 256.663
R1441 B.n812 B.n39 256.663
R1442 B.n812 B.n38 256.663
R1443 B.n812 B.n37 256.663
R1444 B.n812 B.n36 256.663
R1445 B.n812 B.n35 256.663
R1446 B.n812 B.n34 256.663
R1447 B.n470 B.n399 256.663
R1448 B.n473 B.n399 256.663
R1449 B.n479 B.n399 256.663
R1450 B.n481 B.n399 256.663
R1451 B.n487 B.n399 256.663
R1452 B.n489 B.n399 256.663
R1453 B.n495 B.n399 256.663
R1454 B.n497 B.n399 256.663
R1455 B.n503 B.n399 256.663
R1456 B.n505 B.n399 256.663
R1457 B.n511 B.n399 256.663
R1458 B.n513 B.n399 256.663
R1459 B.n519 B.n399 256.663
R1460 B.n521 B.n399 256.663
R1461 B.n527 B.n399 256.663
R1462 B.n529 B.n399 256.663
R1463 B.n535 B.n399 256.663
R1464 B.n537 B.n399 256.663
R1465 B.n543 B.n399 256.663
R1466 B.n545 B.n399 256.663
R1467 B.n551 B.n399 256.663
R1468 B.n553 B.n399 256.663
R1469 B.n559 B.n399 256.663
R1470 B.n561 B.n399 256.663
R1471 B.n567 B.n399 256.663
R1472 B.n569 B.n399 256.663
R1473 B.n575 B.n399 256.663
R1474 B.n577 B.n399 256.663
R1475 B.n583 B.n399 256.663
R1476 B.n585 B.n399 256.663
R1477 B.n594 B.n399 256.663
R1478 B.n596 B.n399 256.663
R1479 B.n602 B.n399 256.663
R1480 B.n604 B.n399 256.663
R1481 B.n610 B.n399 256.663
R1482 B.n612 B.n399 256.663
R1483 B.n619 B.n399 256.663
R1484 B.n621 B.n399 256.663
R1485 B.n627 B.n399 256.663
R1486 B.n629 B.n399 256.663
R1487 B.n635 B.n399 256.663
R1488 B.n637 B.n399 256.663
R1489 B.n643 B.n399 256.663
R1490 B.n645 B.n399 256.663
R1491 B.n651 B.n399 256.663
R1492 B.n653 B.n399 256.663
R1493 B.n659 B.n399 256.663
R1494 B.n661 B.n399 256.663
R1495 B.n667 B.n399 256.663
R1496 B.n669 B.n399 256.663
R1497 B.n675 B.n399 256.663
R1498 B.n677 B.n399 256.663
R1499 B.n683 B.n399 256.663
R1500 B.n685 B.n399 256.663
R1501 B.n691 B.n399 256.663
R1502 B.n693 B.n399 256.663
R1503 B.n699 B.n399 256.663
R1504 B.n701 B.n399 256.663
R1505 B.n707 B.n399 256.663
R1506 B.n709 B.n399 256.663
R1507 B.n715 B.n399 256.663
R1508 B.n717 B.n399 256.663
R1509 B.n723 B.n399 256.663
R1510 B.n725 B.n399 256.663
R1511 B.n731 B.n399 256.663
R1512 B.n734 B.n399 256.663
R1513 B.n741 B.n396 163.367
R1514 B.n745 B.n396 163.367
R1515 B.n745 B.n390 163.367
R1516 B.n754 B.n390 163.367
R1517 B.n754 B.n388 163.367
R1518 B.n758 B.n388 163.367
R1519 B.n758 B.n383 163.367
R1520 B.n766 B.n383 163.367
R1521 B.n766 B.n381 163.367
R1522 B.n770 B.n381 163.367
R1523 B.n770 B.n375 163.367
R1524 B.n779 B.n375 163.367
R1525 B.n779 B.n373 163.367
R1526 B.n783 B.n373 163.367
R1527 B.n783 B.n2 163.367
R1528 B.n846 B.n2 163.367
R1529 B.n846 B.n3 163.367
R1530 B.n842 B.n3 163.367
R1531 B.n842 B.n9 163.367
R1532 B.n838 B.n9 163.367
R1533 B.n838 B.n11 163.367
R1534 B.n834 B.n11 163.367
R1535 B.n834 B.n16 163.367
R1536 B.n830 B.n16 163.367
R1537 B.n830 B.n18 163.367
R1538 B.n826 B.n18 163.367
R1539 B.n826 B.n22 163.367
R1540 B.n822 B.n22 163.367
R1541 B.n822 B.n24 163.367
R1542 B.n818 B.n24 163.367
R1543 B.n818 B.n30 163.367
R1544 B.n814 B.n30 163.367
R1545 B.n472 B.n471 163.367
R1546 B.n474 B.n472 163.367
R1547 B.n478 B.n467 163.367
R1548 B.n482 B.n480 163.367
R1549 B.n486 B.n465 163.367
R1550 B.n490 B.n488 163.367
R1551 B.n494 B.n463 163.367
R1552 B.n498 B.n496 163.367
R1553 B.n502 B.n461 163.367
R1554 B.n506 B.n504 163.367
R1555 B.n510 B.n459 163.367
R1556 B.n514 B.n512 163.367
R1557 B.n518 B.n457 163.367
R1558 B.n522 B.n520 163.367
R1559 B.n526 B.n455 163.367
R1560 B.n530 B.n528 163.367
R1561 B.n534 B.n453 163.367
R1562 B.n538 B.n536 163.367
R1563 B.n542 B.n451 163.367
R1564 B.n546 B.n544 163.367
R1565 B.n550 B.n449 163.367
R1566 B.n554 B.n552 163.367
R1567 B.n558 B.n447 163.367
R1568 B.n562 B.n560 163.367
R1569 B.n566 B.n445 163.367
R1570 B.n570 B.n568 163.367
R1571 B.n574 B.n443 163.367
R1572 B.n578 B.n576 163.367
R1573 B.n582 B.n441 163.367
R1574 B.n586 B.n584 163.367
R1575 B.n593 B.n439 163.367
R1576 B.n597 B.n595 163.367
R1577 B.n601 B.n437 163.367
R1578 B.n605 B.n603 163.367
R1579 B.n609 B.n435 163.367
R1580 B.n613 B.n611 163.367
R1581 B.n618 B.n431 163.367
R1582 B.n622 B.n620 163.367
R1583 B.n626 B.n429 163.367
R1584 B.n630 B.n628 163.367
R1585 B.n634 B.n427 163.367
R1586 B.n638 B.n636 163.367
R1587 B.n642 B.n425 163.367
R1588 B.n646 B.n644 163.367
R1589 B.n650 B.n423 163.367
R1590 B.n654 B.n652 163.367
R1591 B.n658 B.n421 163.367
R1592 B.n662 B.n660 163.367
R1593 B.n666 B.n419 163.367
R1594 B.n670 B.n668 163.367
R1595 B.n674 B.n417 163.367
R1596 B.n678 B.n676 163.367
R1597 B.n682 B.n415 163.367
R1598 B.n686 B.n684 163.367
R1599 B.n690 B.n413 163.367
R1600 B.n694 B.n692 163.367
R1601 B.n698 B.n411 163.367
R1602 B.n702 B.n700 163.367
R1603 B.n706 B.n409 163.367
R1604 B.n710 B.n708 163.367
R1605 B.n714 B.n407 163.367
R1606 B.n718 B.n716 163.367
R1607 B.n722 B.n405 163.367
R1608 B.n726 B.n724 163.367
R1609 B.n730 B.n403 163.367
R1610 B.n733 B.n732 163.367
R1611 B.n735 B.n400 163.367
R1612 B.n739 B.n394 163.367
R1613 B.n747 B.n394 163.367
R1614 B.n747 B.n392 163.367
R1615 B.n751 B.n392 163.367
R1616 B.n751 B.n387 163.367
R1617 B.n760 B.n387 163.367
R1618 B.n760 B.n385 163.367
R1619 B.n764 B.n385 163.367
R1620 B.n764 B.n379 163.367
R1621 B.n772 B.n379 163.367
R1622 B.n772 B.n377 163.367
R1623 B.n777 B.n377 163.367
R1624 B.n777 B.n371 163.367
R1625 B.n785 B.n371 163.367
R1626 B.n786 B.n785 163.367
R1627 B.n786 B.n5 163.367
R1628 B.n6 B.n5 163.367
R1629 B.n7 B.n6 163.367
R1630 B.n791 B.n7 163.367
R1631 B.n791 B.n12 163.367
R1632 B.n13 B.n12 163.367
R1633 B.n14 B.n13 163.367
R1634 B.n796 B.n14 163.367
R1635 B.n796 B.n19 163.367
R1636 B.n20 B.n19 163.367
R1637 B.n21 B.n20 163.367
R1638 B.n801 B.n21 163.367
R1639 B.n801 B.n26 163.367
R1640 B.n27 B.n26 163.367
R1641 B.n28 B.n27 163.367
R1642 B.n806 B.n28 163.367
R1643 B.n806 B.n33 163.367
R1644 B.n109 B.n108 163.367
R1645 B.n113 B.n112 163.367
R1646 B.n117 B.n116 163.367
R1647 B.n121 B.n120 163.367
R1648 B.n125 B.n124 163.367
R1649 B.n129 B.n128 163.367
R1650 B.n133 B.n132 163.367
R1651 B.n137 B.n136 163.367
R1652 B.n141 B.n140 163.367
R1653 B.n145 B.n144 163.367
R1654 B.n149 B.n148 163.367
R1655 B.n153 B.n152 163.367
R1656 B.n157 B.n156 163.367
R1657 B.n161 B.n160 163.367
R1658 B.n165 B.n164 163.367
R1659 B.n169 B.n168 163.367
R1660 B.n173 B.n172 163.367
R1661 B.n177 B.n176 163.367
R1662 B.n181 B.n180 163.367
R1663 B.n185 B.n184 163.367
R1664 B.n189 B.n188 163.367
R1665 B.n193 B.n192 163.367
R1666 B.n197 B.n196 163.367
R1667 B.n201 B.n200 163.367
R1668 B.n205 B.n204 163.367
R1669 B.n209 B.n208 163.367
R1670 B.n213 B.n212 163.367
R1671 B.n217 B.n216 163.367
R1672 B.n221 B.n220 163.367
R1673 B.n225 B.n224 163.367
R1674 B.n229 B.n228 163.367
R1675 B.n233 B.n232 163.367
R1676 B.n237 B.n236 163.367
R1677 B.n241 B.n240 163.367
R1678 B.n245 B.n244 163.367
R1679 B.n249 B.n248 163.367
R1680 B.n253 B.n252 163.367
R1681 B.n257 B.n256 163.367
R1682 B.n261 B.n260 163.367
R1683 B.n265 B.n264 163.367
R1684 B.n269 B.n268 163.367
R1685 B.n273 B.n272 163.367
R1686 B.n277 B.n276 163.367
R1687 B.n281 B.n280 163.367
R1688 B.n285 B.n284 163.367
R1689 B.n289 B.n288 163.367
R1690 B.n293 B.n292 163.367
R1691 B.n297 B.n296 163.367
R1692 B.n301 B.n300 163.367
R1693 B.n305 B.n304 163.367
R1694 B.n309 B.n308 163.367
R1695 B.n313 B.n312 163.367
R1696 B.n317 B.n316 163.367
R1697 B.n321 B.n320 163.367
R1698 B.n325 B.n324 163.367
R1699 B.n329 B.n328 163.367
R1700 B.n333 B.n332 163.367
R1701 B.n337 B.n336 163.367
R1702 B.n341 B.n340 163.367
R1703 B.n345 B.n344 163.367
R1704 B.n349 B.n348 163.367
R1705 B.n353 B.n352 163.367
R1706 B.n357 B.n356 163.367
R1707 B.n361 B.n360 163.367
R1708 B.n365 B.n364 163.367
R1709 B.n367 B.n100 163.367
R1710 B.n470 B.n398 71.676
R1711 B.n474 B.n473 71.676
R1712 B.n479 B.n478 71.676
R1713 B.n482 B.n481 71.676
R1714 B.n487 B.n486 71.676
R1715 B.n490 B.n489 71.676
R1716 B.n495 B.n494 71.676
R1717 B.n498 B.n497 71.676
R1718 B.n503 B.n502 71.676
R1719 B.n506 B.n505 71.676
R1720 B.n511 B.n510 71.676
R1721 B.n514 B.n513 71.676
R1722 B.n519 B.n518 71.676
R1723 B.n522 B.n521 71.676
R1724 B.n527 B.n526 71.676
R1725 B.n530 B.n529 71.676
R1726 B.n535 B.n534 71.676
R1727 B.n538 B.n537 71.676
R1728 B.n543 B.n542 71.676
R1729 B.n546 B.n545 71.676
R1730 B.n551 B.n550 71.676
R1731 B.n554 B.n553 71.676
R1732 B.n559 B.n558 71.676
R1733 B.n562 B.n561 71.676
R1734 B.n567 B.n566 71.676
R1735 B.n570 B.n569 71.676
R1736 B.n575 B.n574 71.676
R1737 B.n578 B.n577 71.676
R1738 B.n583 B.n582 71.676
R1739 B.n586 B.n585 71.676
R1740 B.n594 B.n593 71.676
R1741 B.n597 B.n596 71.676
R1742 B.n602 B.n601 71.676
R1743 B.n605 B.n604 71.676
R1744 B.n610 B.n609 71.676
R1745 B.n613 B.n612 71.676
R1746 B.n619 B.n618 71.676
R1747 B.n622 B.n621 71.676
R1748 B.n627 B.n626 71.676
R1749 B.n630 B.n629 71.676
R1750 B.n635 B.n634 71.676
R1751 B.n638 B.n637 71.676
R1752 B.n643 B.n642 71.676
R1753 B.n646 B.n645 71.676
R1754 B.n651 B.n650 71.676
R1755 B.n654 B.n653 71.676
R1756 B.n659 B.n658 71.676
R1757 B.n662 B.n661 71.676
R1758 B.n667 B.n666 71.676
R1759 B.n670 B.n669 71.676
R1760 B.n675 B.n674 71.676
R1761 B.n678 B.n677 71.676
R1762 B.n683 B.n682 71.676
R1763 B.n686 B.n685 71.676
R1764 B.n691 B.n690 71.676
R1765 B.n694 B.n693 71.676
R1766 B.n699 B.n698 71.676
R1767 B.n702 B.n701 71.676
R1768 B.n707 B.n706 71.676
R1769 B.n710 B.n709 71.676
R1770 B.n715 B.n714 71.676
R1771 B.n718 B.n717 71.676
R1772 B.n723 B.n722 71.676
R1773 B.n726 B.n725 71.676
R1774 B.n731 B.n730 71.676
R1775 B.n734 B.n733 71.676
R1776 B.n34 B.n32 71.676
R1777 B.n109 B.n35 71.676
R1778 B.n113 B.n36 71.676
R1779 B.n117 B.n37 71.676
R1780 B.n121 B.n38 71.676
R1781 B.n125 B.n39 71.676
R1782 B.n129 B.n40 71.676
R1783 B.n133 B.n41 71.676
R1784 B.n137 B.n42 71.676
R1785 B.n141 B.n43 71.676
R1786 B.n145 B.n44 71.676
R1787 B.n149 B.n45 71.676
R1788 B.n153 B.n46 71.676
R1789 B.n157 B.n47 71.676
R1790 B.n161 B.n48 71.676
R1791 B.n165 B.n49 71.676
R1792 B.n169 B.n50 71.676
R1793 B.n173 B.n51 71.676
R1794 B.n177 B.n52 71.676
R1795 B.n181 B.n53 71.676
R1796 B.n185 B.n54 71.676
R1797 B.n189 B.n55 71.676
R1798 B.n193 B.n56 71.676
R1799 B.n197 B.n57 71.676
R1800 B.n201 B.n58 71.676
R1801 B.n205 B.n59 71.676
R1802 B.n209 B.n60 71.676
R1803 B.n213 B.n61 71.676
R1804 B.n217 B.n62 71.676
R1805 B.n221 B.n63 71.676
R1806 B.n225 B.n64 71.676
R1807 B.n229 B.n65 71.676
R1808 B.n233 B.n66 71.676
R1809 B.n237 B.n67 71.676
R1810 B.n241 B.n68 71.676
R1811 B.n245 B.n69 71.676
R1812 B.n249 B.n70 71.676
R1813 B.n253 B.n71 71.676
R1814 B.n257 B.n72 71.676
R1815 B.n261 B.n73 71.676
R1816 B.n265 B.n74 71.676
R1817 B.n269 B.n75 71.676
R1818 B.n273 B.n76 71.676
R1819 B.n277 B.n77 71.676
R1820 B.n281 B.n78 71.676
R1821 B.n285 B.n79 71.676
R1822 B.n289 B.n80 71.676
R1823 B.n293 B.n81 71.676
R1824 B.n297 B.n82 71.676
R1825 B.n301 B.n83 71.676
R1826 B.n305 B.n84 71.676
R1827 B.n309 B.n85 71.676
R1828 B.n313 B.n86 71.676
R1829 B.n317 B.n87 71.676
R1830 B.n321 B.n88 71.676
R1831 B.n325 B.n89 71.676
R1832 B.n329 B.n90 71.676
R1833 B.n333 B.n91 71.676
R1834 B.n337 B.n92 71.676
R1835 B.n341 B.n93 71.676
R1836 B.n345 B.n94 71.676
R1837 B.n349 B.n95 71.676
R1838 B.n353 B.n96 71.676
R1839 B.n357 B.n97 71.676
R1840 B.n361 B.n98 71.676
R1841 B.n365 B.n99 71.676
R1842 B.n811 B.n100 71.676
R1843 B.n811 B.n810 71.676
R1844 B.n367 B.n99 71.676
R1845 B.n364 B.n98 71.676
R1846 B.n360 B.n97 71.676
R1847 B.n356 B.n96 71.676
R1848 B.n352 B.n95 71.676
R1849 B.n348 B.n94 71.676
R1850 B.n344 B.n93 71.676
R1851 B.n340 B.n92 71.676
R1852 B.n336 B.n91 71.676
R1853 B.n332 B.n90 71.676
R1854 B.n328 B.n89 71.676
R1855 B.n324 B.n88 71.676
R1856 B.n320 B.n87 71.676
R1857 B.n316 B.n86 71.676
R1858 B.n312 B.n85 71.676
R1859 B.n308 B.n84 71.676
R1860 B.n304 B.n83 71.676
R1861 B.n300 B.n82 71.676
R1862 B.n296 B.n81 71.676
R1863 B.n292 B.n80 71.676
R1864 B.n288 B.n79 71.676
R1865 B.n284 B.n78 71.676
R1866 B.n280 B.n77 71.676
R1867 B.n276 B.n76 71.676
R1868 B.n272 B.n75 71.676
R1869 B.n268 B.n74 71.676
R1870 B.n264 B.n73 71.676
R1871 B.n260 B.n72 71.676
R1872 B.n256 B.n71 71.676
R1873 B.n252 B.n70 71.676
R1874 B.n248 B.n69 71.676
R1875 B.n244 B.n68 71.676
R1876 B.n240 B.n67 71.676
R1877 B.n236 B.n66 71.676
R1878 B.n232 B.n65 71.676
R1879 B.n228 B.n64 71.676
R1880 B.n224 B.n63 71.676
R1881 B.n220 B.n62 71.676
R1882 B.n216 B.n61 71.676
R1883 B.n212 B.n60 71.676
R1884 B.n208 B.n59 71.676
R1885 B.n204 B.n58 71.676
R1886 B.n200 B.n57 71.676
R1887 B.n196 B.n56 71.676
R1888 B.n192 B.n55 71.676
R1889 B.n188 B.n54 71.676
R1890 B.n184 B.n53 71.676
R1891 B.n180 B.n52 71.676
R1892 B.n176 B.n51 71.676
R1893 B.n172 B.n50 71.676
R1894 B.n168 B.n49 71.676
R1895 B.n164 B.n48 71.676
R1896 B.n160 B.n47 71.676
R1897 B.n156 B.n46 71.676
R1898 B.n152 B.n45 71.676
R1899 B.n148 B.n44 71.676
R1900 B.n144 B.n43 71.676
R1901 B.n140 B.n42 71.676
R1902 B.n136 B.n41 71.676
R1903 B.n132 B.n40 71.676
R1904 B.n128 B.n39 71.676
R1905 B.n124 B.n38 71.676
R1906 B.n120 B.n37 71.676
R1907 B.n116 B.n36 71.676
R1908 B.n112 B.n35 71.676
R1909 B.n108 B.n34 71.676
R1910 B.n471 B.n470 71.676
R1911 B.n473 B.n467 71.676
R1912 B.n480 B.n479 71.676
R1913 B.n481 B.n465 71.676
R1914 B.n488 B.n487 71.676
R1915 B.n489 B.n463 71.676
R1916 B.n496 B.n495 71.676
R1917 B.n497 B.n461 71.676
R1918 B.n504 B.n503 71.676
R1919 B.n505 B.n459 71.676
R1920 B.n512 B.n511 71.676
R1921 B.n513 B.n457 71.676
R1922 B.n520 B.n519 71.676
R1923 B.n521 B.n455 71.676
R1924 B.n528 B.n527 71.676
R1925 B.n529 B.n453 71.676
R1926 B.n536 B.n535 71.676
R1927 B.n537 B.n451 71.676
R1928 B.n544 B.n543 71.676
R1929 B.n545 B.n449 71.676
R1930 B.n552 B.n551 71.676
R1931 B.n553 B.n447 71.676
R1932 B.n560 B.n559 71.676
R1933 B.n561 B.n445 71.676
R1934 B.n568 B.n567 71.676
R1935 B.n569 B.n443 71.676
R1936 B.n576 B.n575 71.676
R1937 B.n577 B.n441 71.676
R1938 B.n584 B.n583 71.676
R1939 B.n585 B.n439 71.676
R1940 B.n595 B.n594 71.676
R1941 B.n596 B.n437 71.676
R1942 B.n603 B.n602 71.676
R1943 B.n604 B.n435 71.676
R1944 B.n611 B.n610 71.676
R1945 B.n612 B.n431 71.676
R1946 B.n620 B.n619 71.676
R1947 B.n621 B.n429 71.676
R1948 B.n628 B.n627 71.676
R1949 B.n629 B.n427 71.676
R1950 B.n636 B.n635 71.676
R1951 B.n637 B.n425 71.676
R1952 B.n644 B.n643 71.676
R1953 B.n645 B.n423 71.676
R1954 B.n652 B.n651 71.676
R1955 B.n653 B.n421 71.676
R1956 B.n660 B.n659 71.676
R1957 B.n661 B.n419 71.676
R1958 B.n668 B.n667 71.676
R1959 B.n669 B.n417 71.676
R1960 B.n676 B.n675 71.676
R1961 B.n677 B.n415 71.676
R1962 B.n684 B.n683 71.676
R1963 B.n685 B.n413 71.676
R1964 B.n692 B.n691 71.676
R1965 B.n693 B.n411 71.676
R1966 B.n700 B.n699 71.676
R1967 B.n701 B.n409 71.676
R1968 B.n708 B.n707 71.676
R1969 B.n709 B.n407 71.676
R1970 B.n716 B.n715 71.676
R1971 B.n717 B.n405 71.676
R1972 B.n724 B.n723 71.676
R1973 B.n725 B.n403 71.676
R1974 B.n732 B.n731 71.676
R1975 B.n735 B.n734 71.676
R1976 B.n740 B.n399 62.8576
R1977 B.n813 B.n812 62.8576
R1978 B.n615 B.n433 59.5399
R1979 B.n591 B.n590 59.5399
R1980 B.n106 B.n105 59.5399
R1981 B.n103 B.n102 59.5399
R1982 B.n815 B.n31 36.3712
R1983 B.n809 B.n808 36.3712
R1984 B.n738 B.n737 36.3712
R1985 B.n742 B.n397 36.3712
R1986 B.n740 B.n395 30.7508
R1987 B.n746 B.n395 30.7508
R1988 B.n746 B.n391 30.7508
R1989 B.n753 B.n391 30.7508
R1990 B.n753 B.n752 30.7508
R1991 B.n759 B.n384 30.7508
R1992 B.n765 B.n384 30.7508
R1993 B.n765 B.n380 30.7508
R1994 B.n771 B.n380 30.7508
R1995 B.n771 B.n376 30.7508
R1996 B.n778 B.n376 30.7508
R1997 B.n784 B.n372 30.7508
R1998 B.n784 B.n4 30.7508
R1999 B.n845 B.n4 30.7508
R2000 B.n845 B.n844 30.7508
R2001 B.n844 B.n843 30.7508
R2002 B.n843 B.n8 30.7508
R2003 B.n837 B.n836 30.7508
R2004 B.n836 B.n835 30.7508
R2005 B.n835 B.n15 30.7508
R2006 B.n829 B.n15 30.7508
R2007 B.n829 B.n828 30.7508
R2008 B.n828 B.n827 30.7508
R2009 B.n821 B.n25 30.7508
R2010 B.n821 B.n820 30.7508
R2011 B.n820 B.n819 30.7508
R2012 B.n819 B.n29 30.7508
R2013 B.n813 B.n29 30.7508
R2014 B.n759 B.t3 27.5853
R2015 B.n827 B.t7 27.5853
R2016 B.n433 B.n432 26.7641
R2017 B.n590 B.n589 26.7641
R2018 B.n105 B.n104 26.7641
R2019 B.n102 B.n101 26.7641
R2020 B.t0 B.n372 19.4455
R2021 B.t1 B.n8 19.4455
R2022 B B.n847 18.0485
R2023 B.n778 B.t0 11.3057
R2024 B.n837 B.t1 11.3057
R2025 B.n107 B.n31 10.6151
R2026 B.n110 B.n107 10.6151
R2027 B.n111 B.n110 10.6151
R2028 B.n114 B.n111 10.6151
R2029 B.n115 B.n114 10.6151
R2030 B.n118 B.n115 10.6151
R2031 B.n119 B.n118 10.6151
R2032 B.n122 B.n119 10.6151
R2033 B.n123 B.n122 10.6151
R2034 B.n126 B.n123 10.6151
R2035 B.n127 B.n126 10.6151
R2036 B.n130 B.n127 10.6151
R2037 B.n131 B.n130 10.6151
R2038 B.n134 B.n131 10.6151
R2039 B.n135 B.n134 10.6151
R2040 B.n138 B.n135 10.6151
R2041 B.n139 B.n138 10.6151
R2042 B.n142 B.n139 10.6151
R2043 B.n143 B.n142 10.6151
R2044 B.n146 B.n143 10.6151
R2045 B.n147 B.n146 10.6151
R2046 B.n150 B.n147 10.6151
R2047 B.n151 B.n150 10.6151
R2048 B.n154 B.n151 10.6151
R2049 B.n155 B.n154 10.6151
R2050 B.n158 B.n155 10.6151
R2051 B.n159 B.n158 10.6151
R2052 B.n162 B.n159 10.6151
R2053 B.n163 B.n162 10.6151
R2054 B.n166 B.n163 10.6151
R2055 B.n167 B.n166 10.6151
R2056 B.n170 B.n167 10.6151
R2057 B.n171 B.n170 10.6151
R2058 B.n174 B.n171 10.6151
R2059 B.n175 B.n174 10.6151
R2060 B.n178 B.n175 10.6151
R2061 B.n179 B.n178 10.6151
R2062 B.n182 B.n179 10.6151
R2063 B.n183 B.n182 10.6151
R2064 B.n186 B.n183 10.6151
R2065 B.n187 B.n186 10.6151
R2066 B.n190 B.n187 10.6151
R2067 B.n191 B.n190 10.6151
R2068 B.n194 B.n191 10.6151
R2069 B.n195 B.n194 10.6151
R2070 B.n198 B.n195 10.6151
R2071 B.n199 B.n198 10.6151
R2072 B.n202 B.n199 10.6151
R2073 B.n203 B.n202 10.6151
R2074 B.n206 B.n203 10.6151
R2075 B.n207 B.n206 10.6151
R2076 B.n210 B.n207 10.6151
R2077 B.n211 B.n210 10.6151
R2078 B.n214 B.n211 10.6151
R2079 B.n215 B.n214 10.6151
R2080 B.n218 B.n215 10.6151
R2081 B.n219 B.n218 10.6151
R2082 B.n222 B.n219 10.6151
R2083 B.n223 B.n222 10.6151
R2084 B.n226 B.n223 10.6151
R2085 B.n227 B.n226 10.6151
R2086 B.n231 B.n230 10.6151
R2087 B.n234 B.n231 10.6151
R2088 B.n235 B.n234 10.6151
R2089 B.n238 B.n235 10.6151
R2090 B.n239 B.n238 10.6151
R2091 B.n242 B.n239 10.6151
R2092 B.n243 B.n242 10.6151
R2093 B.n246 B.n243 10.6151
R2094 B.n247 B.n246 10.6151
R2095 B.n251 B.n250 10.6151
R2096 B.n254 B.n251 10.6151
R2097 B.n255 B.n254 10.6151
R2098 B.n258 B.n255 10.6151
R2099 B.n259 B.n258 10.6151
R2100 B.n262 B.n259 10.6151
R2101 B.n263 B.n262 10.6151
R2102 B.n266 B.n263 10.6151
R2103 B.n267 B.n266 10.6151
R2104 B.n270 B.n267 10.6151
R2105 B.n271 B.n270 10.6151
R2106 B.n274 B.n271 10.6151
R2107 B.n275 B.n274 10.6151
R2108 B.n278 B.n275 10.6151
R2109 B.n279 B.n278 10.6151
R2110 B.n282 B.n279 10.6151
R2111 B.n283 B.n282 10.6151
R2112 B.n286 B.n283 10.6151
R2113 B.n287 B.n286 10.6151
R2114 B.n290 B.n287 10.6151
R2115 B.n291 B.n290 10.6151
R2116 B.n294 B.n291 10.6151
R2117 B.n295 B.n294 10.6151
R2118 B.n298 B.n295 10.6151
R2119 B.n299 B.n298 10.6151
R2120 B.n302 B.n299 10.6151
R2121 B.n303 B.n302 10.6151
R2122 B.n306 B.n303 10.6151
R2123 B.n307 B.n306 10.6151
R2124 B.n310 B.n307 10.6151
R2125 B.n311 B.n310 10.6151
R2126 B.n314 B.n311 10.6151
R2127 B.n315 B.n314 10.6151
R2128 B.n318 B.n315 10.6151
R2129 B.n319 B.n318 10.6151
R2130 B.n322 B.n319 10.6151
R2131 B.n323 B.n322 10.6151
R2132 B.n326 B.n323 10.6151
R2133 B.n327 B.n326 10.6151
R2134 B.n330 B.n327 10.6151
R2135 B.n331 B.n330 10.6151
R2136 B.n334 B.n331 10.6151
R2137 B.n335 B.n334 10.6151
R2138 B.n338 B.n335 10.6151
R2139 B.n339 B.n338 10.6151
R2140 B.n342 B.n339 10.6151
R2141 B.n343 B.n342 10.6151
R2142 B.n346 B.n343 10.6151
R2143 B.n347 B.n346 10.6151
R2144 B.n350 B.n347 10.6151
R2145 B.n351 B.n350 10.6151
R2146 B.n354 B.n351 10.6151
R2147 B.n355 B.n354 10.6151
R2148 B.n358 B.n355 10.6151
R2149 B.n359 B.n358 10.6151
R2150 B.n362 B.n359 10.6151
R2151 B.n363 B.n362 10.6151
R2152 B.n366 B.n363 10.6151
R2153 B.n368 B.n366 10.6151
R2154 B.n369 B.n368 10.6151
R2155 B.n809 B.n369 10.6151
R2156 B.n738 B.n393 10.6151
R2157 B.n748 B.n393 10.6151
R2158 B.n749 B.n748 10.6151
R2159 B.n750 B.n749 10.6151
R2160 B.n750 B.n386 10.6151
R2161 B.n761 B.n386 10.6151
R2162 B.n762 B.n761 10.6151
R2163 B.n763 B.n762 10.6151
R2164 B.n763 B.n378 10.6151
R2165 B.n773 B.n378 10.6151
R2166 B.n774 B.n773 10.6151
R2167 B.n776 B.n774 10.6151
R2168 B.n776 B.n775 10.6151
R2169 B.n775 B.n370 10.6151
R2170 B.n787 B.n370 10.6151
R2171 B.n788 B.n787 10.6151
R2172 B.n789 B.n788 10.6151
R2173 B.n790 B.n789 10.6151
R2174 B.n792 B.n790 10.6151
R2175 B.n793 B.n792 10.6151
R2176 B.n794 B.n793 10.6151
R2177 B.n795 B.n794 10.6151
R2178 B.n797 B.n795 10.6151
R2179 B.n798 B.n797 10.6151
R2180 B.n799 B.n798 10.6151
R2181 B.n800 B.n799 10.6151
R2182 B.n802 B.n800 10.6151
R2183 B.n803 B.n802 10.6151
R2184 B.n804 B.n803 10.6151
R2185 B.n805 B.n804 10.6151
R2186 B.n807 B.n805 10.6151
R2187 B.n808 B.n807 10.6151
R2188 B.n469 B.n397 10.6151
R2189 B.n469 B.n468 10.6151
R2190 B.n475 B.n468 10.6151
R2191 B.n476 B.n475 10.6151
R2192 B.n477 B.n476 10.6151
R2193 B.n477 B.n466 10.6151
R2194 B.n483 B.n466 10.6151
R2195 B.n484 B.n483 10.6151
R2196 B.n485 B.n484 10.6151
R2197 B.n485 B.n464 10.6151
R2198 B.n491 B.n464 10.6151
R2199 B.n492 B.n491 10.6151
R2200 B.n493 B.n492 10.6151
R2201 B.n493 B.n462 10.6151
R2202 B.n499 B.n462 10.6151
R2203 B.n500 B.n499 10.6151
R2204 B.n501 B.n500 10.6151
R2205 B.n501 B.n460 10.6151
R2206 B.n507 B.n460 10.6151
R2207 B.n508 B.n507 10.6151
R2208 B.n509 B.n508 10.6151
R2209 B.n509 B.n458 10.6151
R2210 B.n515 B.n458 10.6151
R2211 B.n516 B.n515 10.6151
R2212 B.n517 B.n516 10.6151
R2213 B.n517 B.n456 10.6151
R2214 B.n523 B.n456 10.6151
R2215 B.n524 B.n523 10.6151
R2216 B.n525 B.n524 10.6151
R2217 B.n525 B.n454 10.6151
R2218 B.n531 B.n454 10.6151
R2219 B.n532 B.n531 10.6151
R2220 B.n533 B.n532 10.6151
R2221 B.n533 B.n452 10.6151
R2222 B.n539 B.n452 10.6151
R2223 B.n540 B.n539 10.6151
R2224 B.n541 B.n540 10.6151
R2225 B.n541 B.n450 10.6151
R2226 B.n547 B.n450 10.6151
R2227 B.n548 B.n547 10.6151
R2228 B.n549 B.n548 10.6151
R2229 B.n549 B.n448 10.6151
R2230 B.n555 B.n448 10.6151
R2231 B.n556 B.n555 10.6151
R2232 B.n557 B.n556 10.6151
R2233 B.n557 B.n446 10.6151
R2234 B.n563 B.n446 10.6151
R2235 B.n564 B.n563 10.6151
R2236 B.n565 B.n564 10.6151
R2237 B.n565 B.n444 10.6151
R2238 B.n571 B.n444 10.6151
R2239 B.n572 B.n571 10.6151
R2240 B.n573 B.n572 10.6151
R2241 B.n573 B.n442 10.6151
R2242 B.n579 B.n442 10.6151
R2243 B.n580 B.n579 10.6151
R2244 B.n581 B.n580 10.6151
R2245 B.n581 B.n440 10.6151
R2246 B.n587 B.n440 10.6151
R2247 B.n588 B.n587 10.6151
R2248 B.n592 B.n588 10.6151
R2249 B.n598 B.n438 10.6151
R2250 B.n599 B.n598 10.6151
R2251 B.n600 B.n599 10.6151
R2252 B.n600 B.n436 10.6151
R2253 B.n606 B.n436 10.6151
R2254 B.n607 B.n606 10.6151
R2255 B.n608 B.n607 10.6151
R2256 B.n608 B.n434 10.6151
R2257 B.n614 B.n434 10.6151
R2258 B.n617 B.n616 10.6151
R2259 B.n617 B.n430 10.6151
R2260 B.n623 B.n430 10.6151
R2261 B.n624 B.n623 10.6151
R2262 B.n625 B.n624 10.6151
R2263 B.n625 B.n428 10.6151
R2264 B.n631 B.n428 10.6151
R2265 B.n632 B.n631 10.6151
R2266 B.n633 B.n632 10.6151
R2267 B.n633 B.n426 10.6151
R2268 B.n639 B.n426 10.6151
R2269 B.n640 B.n639 10.6151
R2270 B.n641 B.n640 10.6151
R2271 B.n641 B.n424 10.6151
R2272 B.n647 B.n424 10.6151
R2273 B.n648 B.n647 10.6151
R2274 B.n649 B.n648 10.6151
R2275 B.n649 B.n422 10.6151
R2276 B.n655 B.n422 10.6151
R2277 B.n656 B.n655 10.6151
R2278 B.n657 B.n656 10.6151
R2279 B.n657 B.n420 10.6151
R2280 B.n663 B.n420 10.6151
R2281 B.n664 B.n663 10.6151
R2282 B.n665 B.n664 10.6151
R2283 B.n665 B.n418 10.6151
R2284 B.n671 B.n418 10.6151
R2285 B.n672 B.n671 10.6151
R2286 B.n673 B.n672 10.6151
R2287 B.n673 B.n416 10.6151
R2288 B.n679 B.n416 10.6151
R2289 B.n680 B.n679 10.6151
R2290 B.n681 B.n680 10.6151
R2291 B.n681 B.n414 10.6151
R2292 B.n687 B.n414 10.6151
R2293 B.n688 B.n687 10.6151
R2294 B.n689 B.n688 10.6151
R2295 B.n689 B.n412 10.6151
R2296 B.n695 B.n412 10.6151
R2297 B.n696 B.n695 10.6151
R2298 B.n697 B.n696 10.6151
R2299 B.n697 B.n410 10.6151
R2300 B.n703 B.n410 10.6151
R2301 B.n704 B.n703 10.6151
R2302 B.n705 B.n704 10.6151
R2303 B.n705 B.n408 10.6151
R2304 B.n711 B.n408 10.6151
R2305 B.n712 B.n711 10.6151
R2306 B.n713 B.n712 10.6151
R2307 B.n713 B.n406 10.6151
R2308 B.n719 B.n406 10.6151
R2309 B.n720 B.n719 10.6151
R2310 B.n721 B.n720 10.6151
R2311 B.n721 B.n404 10.6151
R2312 B.n727 B.n404 10.6151
R2313 B.n728 B.n727 10.6151
R2314 B.n729 B.n728 10.6151
R2315 B.n729 B.n402 10.6151
R2316 B.n402 B.n401 10.6151
R2317 B.n736 B.n401 10.6151
R2318 B.n737 B.n736 10.6151
R2319 B.n743 B.n742 10.6151
R2320 B.n744 B.n743 10.6151
R2321 B.n744 B.n389 10.6151
R2322 B.n755 B.n389 10.6151
R2323 B.n756 B.n755 10.6151
R2324 B.n757 B.n756 10.6151
R2325 B.n757 B.n382 10.6151
R2326 B.n767 B.n382 10.6151
R2327 B.n768 B.n767 10.6151
R2328 B.n769 B.n768 10.6151
R2329 B.n769 B.n374 10.6151
R2330 B.n780 B.n374 10.6151
R2331 B.n781 B.n780 10.6151
R2332 B.n782 B.n781 10.6151
R2333 B.n782 B.n0 10.6151
R2334 B.n841 B.n1 10.6151
R2335 B.n841 B.n840 10.6151
R2336 B.n840 B.n839 10.6151
R2337 B.n839 B.n10 10.6151
R2338 B.n833 B.n10 10.6151
R2339 B.n833 B.n832 10.6151
R2340 B.n832 B.n831 10.6151
R2341 B.n831 B.n17 10.6151
R2342 B.n825 B.n17 10.6151
R2343 B.n825 B.n824 10.6151
R2344 B.n824 B.n823 10.6151
R2345 B.n823 B.n23 10.6151
R2346 B.n817 B.n23 10.6151
R2347 B.n817 B.n816 10.6151
R2348 B.n816 B.n815 10.6151
R2349 B.n227 B.n106 8.74196
R2350 B.n250 B.n103 8.74196
R2351 B.n592 B.n591 8.74196
R2352 B.n616 B.n615 8.74196
R2353 B.n752 B.t3 3.16597
R2354 B.n25 B.t7 3.16597
R2355 B.n847 B.n0 2.81026
R2356 B.n847 B.n1 2.81026
R2357 B.n230 B.n106 1.87367
R2358 B.n247 B.n103 1.87367
R2359 B.n591 B.n438 1.87367
R2360 B.n615 B.n614 1.87367
R2361 VP.n0 VP.t0 681.612
R2362 VP.n0 VP.t1 635.726
R2363 VP VP.n0 0.0516364
R2364 VDD1.n100 VDD1.n0 289.615
R2365 VDD1.n205 VDD1.n105 289.615
R2366 VDD1.n101 VDD1.n100 185
R2367 VDD1.n99 VDD1.n98 185
R2368 VDD1.n4 VDD1.n3 185
R2369 VDD1.n93 VDD1.n92 185
R2370 VDD1.n91 VDD1.n90 185
R2371 VDD1.n8 VDD1.n7 185
R2372 VDD1.n85 VDD1.n84 185
R2373 VDD1.n83 VDD1.n82 185
R2374 VDD1.n81 VDD1.n11 185
R2375 VDD1.n15 VDD1.n12 185
R2376 VDD1.n76 VDD1.n75 185
R2377 VDD1.n74 VDD1.n73 185
R2378 VDD1.n17 VDD1.n16 185
R2379 VDD1.n68 VDD1.n67 185
R2380 VDD1.n66 VDD1.n65 185
R2381 VDD1.n21 VDD1.n20 185
R2382 VDD1.n60 VDD1.n59 185
R2383 VDD1.n58 VDD1.n57 185
R2384 VDD1.n25 VDD1.n24 185
R2385 VDD1.n52 VDD1.n51 185
R2386 VDD1.n50 VDD1.n49 185
R2387 VDD1.n29 VDD1.n28 185
R2388 VDD1.n44 VDD1.n43 185
R2389 VDD1.n42 VDD1.n41 185
R2390 VDD1.n33 VDD1.n32 185
R2391 VDD1.n36 VDD1.n35 185
R2392 VDD1.n140 VDD1.n139 185
R2393 VDD1.n137 VDD1.n136 185
R2394 VDD1.n146 VDD1.n145 185
R2395 VDD1.n148 VDD1.n147 185
R2396 VDD1.n133 VDD1.n132 185
R2397 VDD1.n154 VDD1.n153 185
R2398 VDD1.n156 VDD1.n155 185
R2399 VDD1.n129 VDD1.n128 185
R2400 VDD1.n162 VDD1.n161 185
R2401 VDD1.n164 VDD1.n163 185
R2402 VDD1.n125 VDD1.n124 185
R2403 VDD1.n170 VDD1.n169 185
R2404 VDD1.n172 VDD1.n171 185
R2405 VDD1.n121 VDD1.n120 185
R2406 VDD1.n178 VDD1.n177 185
R2407 VDD1.n181 VDD1.n180 185
R2408 VDD1.n179 VDD1.n117 185
R2409 VDD1.n186 VDD1.n116 185
R2410 VDD1.n188 VDD1.n187 185
R2411 VDD1.n190 VDD1.n189 185
R2412 VDD1.n113 VDD1.n112 185
R2413 VDD1.n196 VDD1.n195 185
R2414 VDD1.n198 VDD1.n197 185
R2415 VDD1.n109 VDD1.n108 185
R2416 VDD1.n204 VDD1.n203 185
R2417 VDD1.n206 VDD1.n205 185
R2418 VDD1.t1 VDD1.n34 147.659
R2419 VDD1.t0 VDD1.n138 147.659
R2420 VDD1.n100 VDD1.n99 104.615
R2421 VDD1.n99 VDD1.n3 104.615
R2422 VDD1.n92 VDD1.n3 104.615
R2423 VDD1.n92 VDD1.n91 104.615
R2424 VDD1.n91 VDD1.n7 104.615
R2425 VDD1.n84 VDD1.n7 104.615
R2426 VDD1.n84 VDD1.n83 104.615
R2427 VDD1.n83 VDD1.n11 104.615
R2428 VDD1.n15 VDD1.n11 104.615
R2429 VDD1.n75 VDD1.n15 104.615
R2430 VDD1.n75 VDD1.n74 104.615
R2431 VDD1.n74 VDD1.n16 104.615
R2432 VDD1.n67 VDD1.n16 104.615
R2433 VDD1.n67 VDD1.n66 104.615
R2434 VDD1.n66 VDD1.n20 104.615
R2435 VDD1.n59 VDD1.n20 104.615
R2436 VDD1.n59 VDD1.n58 104.615
R2437 VDD1.n58 VDD1.n24 104.615
R2438 VDD1.n51 VDD1.n24 104.615
R2439 VDD1.n51 VDD1.n50 104.615
R2440 VDD1.n50 VDD1.n28 104.615
R2441 VDD1.n43 VDD1.n28 104.615
R2442 VDD1.n43 VDD1.n42 104.615
R2443 VDD1.n42 VDD1.n32 104.615
R2444 VDD1.n35 VDD1.n32 104.615
R2445 VDD1.n139 VDD1.n136 104.615
R2446 VDD1.n146 VDD1.n136 104.615
R2447 VDD1.n147 VDD1.n146 104.615
R2448 VDD1.n147 VDD1.n132 104.615
R2449 VDD1.n154 VDD1.n132 104.615
R2450 VDD1.n155 VDD1.n154 104.615
R2451 VDD1.n155 VDD1.n128 104.615
R2452 VDD1.n162 VDD1.n128 104.615
R2453 VDD1.n163 VDD1.n162 104.615
R2454 VDD1.n163 VDD1.n124 104.615
R2455 VDD1.n170 VDD1.n124 104.615
R2456 VDD1.n171 VDD1.n170 104.615
R2457 VDD1.n171 VDD1.n120 104.615
R2458 VDD1.n178 VDD1.n120 104.615
R2459 VDD1.n180 VDD1.n178 104.615
R2460 VDD1.n180 VDD1.n179 104.615
R2461 VDD1.n179 VDD1.n116 104.615
R2462 VDD1.n188 VDD1.n116 104.615
R2463 VDD1.n189 VDD1.n188 104.615
R2464 VDD1.n189 VDD1.n112 104.615
R2465 VDD1.n196 VDD1.n112 104.615
R2466 VDD1.n197 VDD1.n196 104.615
R2467 VDD1.n197 VDD1.n108 104.615
R2468 VDD1.n204 VDD1.n108 104.615
R2469 VDD1.n205 VDD1.n204 104.615
R2470 VDD1 VDD1.n209 93.5051
R2471 VDD1.n35 VDD1.t1 52.3082
R2472 VDD1.n139 VDD1.t0 52.3082
R2473 VDD1 VDD1.n104 50.5773
R2474 VDD1.n36 VDD1.n34 15.6677
R2475 VDD1.n140 VDD1.n138 15.6677
R2476 VDD1.n82 VDD1.n81 13.1884
R2477 VDD1.n187 VDD1.n186 13.1884
R2478 VDD1.n85 VDD1.n10 12.8005
R2479 VDD1.n80 VDD1.n12 12.8005
R2480 VDD1.n37 VDD1.n33 12.8005
R2481 VDD1.n141 VDD1.n137 12.8005
R2482 VDD1.n185 VDD1.n117 12.8005
R2483 VDD1.n190 VDD1.n115 12.8005
R2484 VDD1.n86 VDD1.n8 12.0247
R2485 VDD1.n77 VDD1.n76 12.0247
R2486 VDD1.n41 VDD1.n40 12.0247
R2487 VDD1.n145 VDD1.n144 12.0247
R2488 VDD1.n182 VDD1.n181 12.0247
R2489 VDD1.n191 VDD1.n113 12.0247
R2490 VDD1.n90 VDD1.n89 11.249
R2491 VDD1.n73 VDD1.n14 11.249
R2492 VDD1.n44 VDD1.n31 11.249
R2493 VDD1.n148 VDD1.n135 11.249
R2494 VDD1.n177 VDD1.n119 11.249
R2495 VDD1.n195 VDD1.n194 11.249
R2496 VDD1.n93 VDD1.n6 10.4732
R2497 VDD1.n72 VDD1.n17 10.4732
R2498 VDD1.n45 VDD1.n29 10.4732
R2499 VDD1.n149 VDD1.n133 10.4732
R2500 VDD1.n176 VDD1.n121 10.4732
R2501 VDD1.n198 VDD1.n111 10.4732
R2502 VDD1.n94 VDD1.n4 9.69747
R2503 VDD1.n69 VDD1.n68 9.69747
R2504 VDD1.n49 VDD1.n48 9.69747
R2505 VDD1.n153 VDD1.n152 9.69747
R2506 VDD1.n173 VDD1.n172 9.69747
R2507 VDD1.n199 VDD1.n109 9.69747
R2508 VDD1.n104 VDD1.n103 9.45567
R2509 VDD1.n209 VDD1.n208 9.45567
R2510 VDD1.n62 VDD1.n61 9.3005
R2511 VDD1.n64 VDD1.n63 9.3005
R2512 VDD1.n19 VDD1.n18 9.3005
R2513 VDD1.n70 VDD1.n69 9.3005
R2514 VDD1.n72 VDD1.n71 9.3005
R2515 VDD1.n14 VDD1.n13 9.3005
R2516 VDD1.n78 VDD1.n77 9.3005
R2517 VDD1.n80 VDD1.n79 9.3005
R2518 VDD1.n103 VDD1.n102 9.3005
R2519 VDD1.n2 VDD1.n1 9.3005
R2520 VDD1.n97 VDD1.n96 9.3005
R2521 VDD1.n95 VDD1.n94 9.3005
R2522 VDD1.n6 VDD1.n5 9.3005
R2523 VDD1.n89 VDD1.n88 9.3005
R2524 VDD1.n87 VDD1.n86 9.3005
R2525 VDD1.n10 VDD1.n9 9.3005
R2526 VDD1.n23 VDD1.n22 9.3005
R2527 VDD1.n56 VDD1.n55 9.3005
R2528 VDD1.n54 VDD1.n53 9.3005
R2529 VDD1.n27 VDD1.n26 9.3005
R2530 VDD1.n48 VDD1.n47 9.3005
R2531 VDD1.n46 VDD1.n45 9.3005
R2532 VDD1.n31 VDD1.n30 9.3005
R2533 VDD1.n40 VDD1.n39 9.3005
R2534 VDD1.n38 VDD1.n37 9.3005
R2535 VDD1.n107 VDD1.n106 9.3005
R2536 VDD1.n202 VDD1.n201 9.3005
R2537 VDD1.n200 VDD1.n199 9.3005
R2538 VDD1.n111 VDD1.n110 9.3005
R2539 VDD1.n194 VDD1.n193 9.3005
R2540 VDD1.n192 VDD1.n191 9.3005
R2541 VDD1.n115 VDD1.n114 9.3005
R2542 VDD1.n160 VDD1.n159 9.3005
R2543 VDD1.n158 VDD1.n157 9.3005
R2544 VDD1.n131 VDD1.n130 9.3005
R2545 VDD1.n152 VDD1.n151 9.3005
R2546 VDD1.n150 VDD1.n149 9.3005
R2547 VDD1.n135 VDD1.n134 9.3005
R2548 VDD1.n144 VDD1.n143 9.3005
R2549 VDD1.n142 VDD1.n141 9.3005
R2550 VDD1.n127 VDD1.n126 9.3005
R2551 VDD1.n166 VDD1.n165 9.3005
R2552 VDD1.n168 VDD1.n167 9.3005
R2553 VDD1.n123 VDD1.n122 9.3005
R2554 VDD1.n174 VDD1.n173 9.3005
R2555 VDD1.n176 VDD1.n175 9.3005
R2556 VDD1.n119 VDD1.n118 9.3005
R2557 VDD1.n183 VDD1.n182 9.3005
R2558 VDD1.n185 VDD1.n184 9.3005
R2559 VDD1.n208 VDD1.n207 9.3005
R2560 VDD1.n98 VDD1.n97 8.92171
R2561 VDD1.n65 VDD1.n19 8.92171
R2562 VDD1.n52 VDD1.n27 8.92171
R2563 VDD1.n156 VDD1.n131 8.92171
R2564 VDD1.n169 VDD1.n123 8.92171
R2565 VDD1.n203 VDD1.n202 8.92171
R2566 VDD1.n101 VDD1.n2 8.14595
R2567 VDD1.n64 VDD1.n21 8.14595
R2568 VDD1.n53 VDD1.n25 8.14595
R2569 VDD1.n157 VDD1.n129 8.14595
R2570 VDD1.n168 VDD1.n125 8.14595
R2571 VDD1.n206 VDD1.n107 8.14595
R2572 VDD1.n102 VDD1.n0 7.3702
R2573 VDD1.n61 VDD1.n60 7.3702
R2574 VDD1.n57 VDD1.n56 7.3702
R2575 VDD1.n161 VDD1.n160 7.3702
R2576 VDD1.n165 VDD1.n164 7.3702
R2577 VDD1.n207 VDD1.n105 7.3702
R2578 VDD1.n104 VDD1.n0 6.59444
R2579 VDD1.n60 VDD1.n23 6.59444
R2580 VDD1.n57 VDD1.n23 6.59444
R2581 VDD1.n161 VDD1.n127 6.59444
R2582 VDD1.n164 VDD1.n127 6.59444
R2583 VDD1.n209 VDD1.n105 6.59444
R2584 VDD1.n102 VDD1.n101 5.81868
R2585 VDD1.n61 VDD1.n21 5.81868
R2586 VDD1.n56 VDD1.n25 5.81868
R2587 VDD1.n160 VDD1.n129 5.81868
R2588 VDD1.n165 VDD1.n125 5.81868
R2589 VDD1.n207 VDD1.n206 5.81868
R2590 VDD1.n98 VDD1.n2 5.04292
R2591 VDD1.n65 VDD1.n64 5.04292
R2592 VDD1.n53 VDD1.n52 5.04292
R2593 VDD1.n157 VDD1.n156 5.04292
R2594 VDD1.n169 VDD1.n168 5.04292
R2595 VDD1.n203 VDD1.n107 5.04292
R2596 VDD1.n38 VDD1.n34 4.38563
R2597 VDD1.n142 VDD1.n138 4.38563
R2598 VDD1.n97 VDD1.n4 4.26717
R2599 VDD1.n68 VDD1.n19 4.26717
R2600 VDD1.n49 VDD1.n27 4.26717
R2601 VDD1.n153 VDD1.n131 4.26717
R2602 VDD1.n172 VDD1.n123 4.26717
R2603 VDD1.n202 VDD1.n109 4.26717
R2604 VDD1.n94 VDD1.n93 3.49141
R2605 VDD1.n69 VDD1.n17 3.49141
R2606 VDD1.n48 VDD1.n29 3.49141
R2607 VDD1.n152 VDD1.n133 3.49141
R2608 VDD1.n173 VDD1.n121 3.49141
R2609 VDD1.n199 VDD1.n198 3.49141
R2610 VDD1.n90 VDD1.n6 2.71565
R2611 VDD1.n73 VDD1.n72 2.71565
R2612 VDD1.n45 VDD1.n44 2.71565
R2613 VDD1.n149 VDD1.n148 2.71565
R2614 VDD1.n177 VDD1.n176 2.71565
R2615 VDD1.n195 VDD1.n111 2.71565
R2616 VDD1.n89 VDD1.n8 1.93989
R2617 VDD1.n76 VDD1.n14 1.93989
R2618 VDD1.n41 VDD1.n31 1.93989
R2619 VDD1.n145 VDD1.n135 1.93989
R2620 VDD1.n181 VDD1.n119 1.93989
R2621 VDD1.n194 VDD1.n113 1.93989
R2622 VDD1.n86 VDD1.n85 1.16414
R2623 VDD1.n77 VDD1.n12 1.16414
R2624 VDD1.n40 VDD1.n33 1.16414
R2625 VDD1.n144 VDD1.n137 1.16414
R2626 VDD1.n182 VDD1.n117 1.16414
R2627 VDD1.n191 VDD1.n190 1.16414
R2628 VDD1.n82 VDD1.n10 0.388379
R2629 VDD1.n81 VDD1.n80 0.388379
R2630 VDD1.n37 VDD1.n36 0.388379
R2631 VDD1.n141 VDD1.n140 0.388379
R2632 VDD1.n186 VDD1.n185 0.388379
R2633 VDD1.n187 VDD1.n115 0.388379
R2634 VDD1.n103 VDD1.n1 0.155672
R2635 VDD1.n96 VDD1.n1 0.155672
R2636 VDD1.n96 VDD1.n95 0.155672
R2637 VDD1.n95 VDD1.n5 0.155672
R2638 VDD1.n88 VDD1.n5 0.155672
R2639 VDD1.n88 VDD1.n87 0.155672
R2640 VDD1.n87 VDD1.n9 0.155672
R2641 VDD1.n79 VDD1.n9 0.155672
R2642 VDD1.n79 VDD1.n78 0.155672
R2643 VDD1.n78 VDD1.n13 0.155672
R2644 VDD1.n71 VDD1.n13 0.155672
R2645 VDD1.n71 VDD1.n70 0.155672
R2646 VDD1.n70 VDD1.n18 0.155672
R2647 VDD1.n63 VDD1.n18 0.155672
R2648 VDD1.n63 VDD1.n62 0.155672
R2649 VDD1.n62 VDD1.n22 0.155672
R2650 VDD1.n55 VDD1.n22 0.155672
R2651 VDD1.n55 VDD1.n54 0.155672
R2652 VDD1.n54 VDD1.n26 0.155672
R2653 VDD1.n47 VDD1.n26 0.155672
R2654 VDD1.n47 VDD1.n46 0.155672
R2655 VDD1.n46 VDD1.n30 0.155672
R2656 VDD1.n39 VDD1.n30 0.155672
R2657 VDD1.n39 VDD1.n38 0.155672
R2658 VDD1.n143 VDD1.n142 0.155672
R2659 VDD1.n143 VDD1.n134 0.155672
R2660 VDD1.n150 VDD1.n134 0.155672
R2661 VDD1.n151 VDD1.n150 0.155672
R2662 VDD1.n151 VDD1.n130 0.155672
R2663 VDD1.n158 VDD1.n130 0.155672
R2664 VDD1.n159 VDD1.n158 0.155672
R2665 VDD1.n159 VDD1.n126 0.155672
R2666 VDD1.n166 VDD1.n126 0.155672
R2667 VDD1.n167 VDD1.n166 0.155672
R2668 VDD1.n167 VDD1.n122 0.155672
R2669 VDD1.n174 VDD1.n122 0.155672
R2670 VDD1.n175 VDD1.n174 0.155672
R2671 VDD1.n175 VDD1.n118 0.155672
R2672 VDD1.n183 VDD1.n118 0.155672
R2673 VDD1.n184 VDD1.n183 0.155672
R2674 VDD1.n184 VDD1.n114 0.155672
R2675 VDD1.n192 VDD1.n114 0.155672
R2676 VDD1.n193 VDD1.n192 0.155672
R2677 VDD1.n193 VDD1.n110 0.155672
R2678 VDD1.n200 VDD1.n110 0.155672
R2679 VDD1.n201 VDD1.n200 0.155672
R2680 VDD1.n201 VDD1.n106 0.155672
R2681 VDD1.n208 VDD1.n106 0.155672
C0 VDD1 VDD2 0.498932f
C1 VDD2 VP 0.270487f
C2 VN VTAIL 2.70041f
C3 VDD1 VN 0.148748f
C4 VN VP 6.02164f
C5 VDD2 VN 3.4604f
C6 VDD1 VTAIL 7.55664f
C7 VTAIL VP 2.71516f
C8 VDD2 VTAIL 7.59081f
C9 VDD1 VP 3.5762f
C10 VDD2 B 5.149545f
C11 VDD1 B 8.178639f
C12 VTAIL B 9.271819f
C13 VN B 11.027189f
C14 VP B 4.930318f
C15 VDD1.n0 B 0.030171f
C16 VDD1.n1 B 0.020388f
C17 VDD1.n2 B 0.010956f
C18 VDD1.n3 B 0.025895f
C19 VDD1.n4 B 0.0116f
C20 VDD1.n5 B 0.020388f
C21 VDD1.n6 B 0.010956f
C22 VDD1.n7 B 0.025895f
C23 VDD1.n8 B 0.0116f
C24 VDD1.n9 B 0.020388f
C25 VDD1.n10 B 0.010956f
C26 VDD1.n11 B 0.025895f
C27 VDD1.n12 B 0.0116f
C28 VDD1.n13 B 0.020388f
C29 VDD1.n14 B 0.010956f
C30 VDD1.n15 B 0.025895f
C31 VDD1.n16 B 0.025895f
C32 VDD1.n17 B 0.0116f
C33 VDD1.n18 B 0.020388f
C34 VDD1.n19 B 0.010956f
C35 VDD1.n20 B 0.025895f
C36 VDD1.n21 B 0.0116f
C37 VDD1.n22 B 0.020388f
C38 VDD1.n23 B 0.010956f
C39 VDD1.n24 B 0.025895f
C40 VDD1.n25 B 0.0116f
C41 VDD1.n26 B 0.020388f
C42 VDD1.n27 B 0.010956f
C43 VDD1.n28 B 0.025895f
C44 VDD1.n29 B 0.0116f
C45 VDD1.n30 B 0.020388f
C46 VDD1.n31 B 0.010956f
C47 VDD1.n32 B 0.025895f
C48 VDD1.n33 B 0.0116f
C49 VDD1.n34 B 0.153576f
C50 VDD1.t1 B 0.04298f
C51 VDD1.n35 B 0.019421f
C52 VDD1.n36 B 0.015297f
C53 VDD1.n37 B 0.010956f
C54 VDD1.n38 B 1.70304f
C55 VDD1.n39 B 0.020388f
C56 VDD1.n40 B 0.010956f
C57 VDD1.n41 B 0.0116f
C58 VDD1.n42 B 0.025895f
C59 VDD1.n43 B 0.025895f
C60 VDD1.n44 B 0.0116f
C61 VDD1.n45 B 0.010956f
C62 VDD1.n46 B 0.020388f
C63 VDD1.n47 B 0.020388f
C64 VDD1.n48 B 0.010956f
C65 VDD1.n49 B 0.0116f
C66 VDD1.n50 B 0.025895f
C67 VDD1.n51 B 0.025895f
C68 VDD1.n52 B 0.0116f
C69 VDD1.n53 B 0.010956f
C70 VDD1.n54 B 0.020388f
C71 VDD1.n55 B 0.020388f
C72 VDD1.n56 B 0.010956f
C73 VDD1.n57 B 0.0116f
C74 VDD1.n58 B 0.025895f
C75 VDD1.n59 B 0.025895f
C76 VDD1.n60 B 0.0116f
C77 VDD1.n61 B 0.010956f
C78 VDD1.n62 B 0.020388f
C79 VDD1.n63 B 0.020388f
C80 VDD1.n64 B 0.010956f
C81 VDD1.n65 B 0.0116f
C82 VDD1.n66 B 0.025895f
C83 VDD1.n67 B 0.025895f
C84 VDD1.n68 B 0.0116f
C85 VDD1.n69 B 0.010956f
C86 VDD1.n70 B 0.020388f
C87 VDD1.n71 B 0.020388f
C88 VDD1.n72 B 0.010956f
C89 VDD1.n73 B 0.0116f
C90 VDD1.n74 B 0.025895f
C91 VDD1.n75 B 0.025895f
C92 VDD1.n76 B 0.0116f
C93 VDD1.n77 B 0.010956f
C94 VDD1.n78 B 0.020388f
C95 VDD1.n79 B 0.020388f
C96 VDD1.n80 B 0.010956f
C97 VDD1.n81 B 0.011278f
C98 VDD1.n82 B 0.011278f
C99 VDD1.n83 B 0.025895f
C100 VDD1.n84 B 0.025895f
C101 VDD1.n85 B 0.0116f
C102 VDD1.n86 B 0.010956f
C103 VDD1.n87 B 0.020388f
C104 VDD1.n88 B 0.020388f
C105 VDD1.n89 B 0.010956f
C106 VDD1.n90 B 0.0116f
C107 VDD1.n91 B 0.025895f
C108 VDD1.n92 B 0.025895f
C109 VDD1.n93 B 0.0116f
C110 VDD1.n94 B 0.010956f
C111 VDD1.n95 B 0.020388f
C112 VDD1.n96 B 0.020388f
C113 VDD1.n97 B 0.010956f
C114 VDD1.n98 B 0.0116f
C115 VDD1.n99 B 0.025895f
C116 VDD1.n100 B 0.058735f
C117 VDD1.n101 B 0.0116f
C118 VDD1.n102 B 0.010956f
C119 VDD1.n103 B 0.049076f
C120 VDD1.n104 B 0.047709f
C121 VDD1.n105 B 0.030171f
C122 VDD1.n106 B 0.020388f
C123 VDD1.n107 B 0.010956f
C124 VDD1.n108 B 0.025895f
C125 VDD1.n109 B 0.0116f
C126 VDD1.n110 B 0.020388f
C127 VDD1.n111 B 0.010956f
C128 VDD1.n112 B 0.025895f
C129 VDD1.n113 B 0.0116f
C130 VDD1.n114 B 0.020388f
C131 VDD1.n115 B 0.010956f
C132 VDD1.n116 B 0.025895f
C133 VDD1.n117 B 0.0116f
C134 VDD1.n118 B 0.020388f
C135 VDD1.n119 B 0.010956f
C136 VDD1.n120 B 0.025895f
C137 VDD1.n121 B 0.0116f
C138 VDD1.n122 B 0.020388f
C139 VDD1.n123 B 0.010956f
C140 VDD1.n124 B 0.025895f
C141 VDD1.n125 B 0.0116f
C142 VDD1.n126 B 0.020388f
C143 VDD1.n127 B 0.010956f
C144 VDD1.n128 B 0.025895f
C145 VDD1.n129 B 0.0116f
C146 VDD1.n130 B 0.020388f
C147 VDD1.n131 B 0.010956f
C148 VDD1.n132 B 0.025895f
C149 VDD1.n133 B 0.0116f
C150 VDD1.n134 B 0.020388f
C151 VDD1.n135 B 0.010956f
C152 VDD1.n136 B 0.025895f
C153 VDD1.n137 B 0.0116f
C154 VDD1.n138 B 0.153576f
C155 VDD1.t0 B 0.04298f
C156 VDD1.n139 B 0.019421f
C157 VDD1.n140 B 0.015297f
C158 VDD1.n141 B 0.010956f
C159 VDD1.n142 B 1.70304f
C160 VDD1.n143 B 0.020388f
C161 VDD1.n144 B 0.010956f
C162 VDD1.n145 B 0.0116f
C163 VDD1.n146 B 0.025895f
C164 VDD1.n147 B 0.025895f
C165 VDD1.n148 B 0.0116f
C166 VDD1.n149 B 0.010956f
C167 VDD1.n150 B 0.020388f
C168 VDD1.n151 B 0.020388f
C169 VDD1.n152 B 0.010956f
C170 VDD1.n153 B 0.0116f
C171 VDD1.n154 B 0.025895f
C172 VDD1.n155 B 0.025895f
C173 VDD1.n156 B 0.0116f
C174 VDD1.n157 B 0.010956f
C175 VDD1.n158 B 0.020388f
C176 VDD1.n159 B 0.020388f
C177 VDD1.n160 B 0.010956f
C178 VDD1.n161 B 0.0116f
C179 VDD1.n162 B 0.025895f
C180 VDD1.n163 B 0.025895f
C181 VDD1.n164 B 0.0116f
C182 VDD1.n165 B 0.010956f
C183 VDD1.n166 B 0.020388f
C184 VDD1.n167 B 0.020388f
C185 VDD1.n168 B 0.010956f
C186 VDD1.n169 B 0.0116f
C187 VDD1.n170 B 0.025895f
C188 VDD1.n171 B 0.025895f
C189 VDD1.n172 B 0.0116f
C190 VDD1.n173 B 0.010956f
C191 VDD1.n174 B 0.020388f
C192 VDD1.n175 B 0.020388f
C193 VDD1.n176 B 0.010956f
C194 VDD1.n177 B 0.0116f
C195 VDD1.n178 B 0.025895f
C196 VDD1.n179 B 0.025895f
C197 VDD1.n180 B 0.025895f
C198 VDD1.n181 B 0.0116f
C199 VDD1.n182 B 0.010956f
C200 VDD1.n183 B 0.020388f
C201 VDD1.n184 B 0.020388f
C202 VDD1.n185 B 0.010956f
C203 VDD1.n186 B 0.011278f
C204 VDD1.n187 B 0.011278f
C205 VDD1.n188 B 0.025895f
C206 VDD1.n189 B 0.025895f
C207 VDD1.n190 B 0.0116f
C208 VDD1.n191 B 0.010956f
C209 VDD1.n192 B 0.020388f
C210 VDD1.n193 B 0.020388f
C211 VDD1.n194 B 0.010956f
C212 VDD1.n195 B 0.0116f
C213 VDD1.n196 B 0.025895f
C214 VDD1.n197 B 0.025895f
C215 VDD1.n198 B 0.0116f
C216 VDD1.n199 B 0.010956f
C217 VDD1.n200 B 0.020388f
C218 VDD1.n201 B 0.020388f
C219 VDD1.n202 B 0.010956f
C220 VDD1.n203 B 0.0116f
C221 VDD1.n204 B 0.025895f
C222 VDD1.n205 B 0.058735f
C223 VDD1.n206 B 0.0116f
C224 VDD1.n207 B 0.010956f
C225 VDD1.n208 B 0.049076f
C226 VDD1.n209 B 0.750692f
C227 VP.t0 B 3.23376f
C228 VP.t1 B 3.02466f
C229 VP.n0 B 6.01404f
C230 VDD2.n0 B 0.030104f
C231 VDD2.n1 B 0.020343f
C232 VDD2.n2 B 0.010931f
C233 VDD2.n3 B 0.025838f
C234 VDD2.n4 B 0.011574f
C235 VDD2.n5 B 0.020343f
C236 VDD2.n6 B 0.010931f
C237 VDD2.n7 B 0.025838f
C238 VDD2.n8 B 0.011574f
C239 VDD2.n9 B 0.020343f
C240 VDD2.n10 B 0.010931f
C241 VDD2.n11 B 0.025838f
C242 VDD2.n12 B 0.011574f
C243 VDD2.n13 B 0.020343f
C244 VDD2.n14 B 0.010931f
C245 VDD2.n15 B 0.025838f
C246 VDD2.n16 B 0.011574f
C247 VDD2.n17 B 0.020343f
C248 VDD2.n18 B 0.010931f
C249 VDD2.n19 B 0.025838f
C250 VDD2.n20 B 0.011574f
C251 VDD2.n21 B 0.020343f
C252 VDD2.n22 B 0.010931f
C253 VDD2.n23 B 0.025838f
C254 VDD2.n24 B 0.011574f
C255 VDD2.n25 B 0.020343f
C256 VDD2.n26 B 0.010931f
C257 VDD2.n27 B 0.025838f
C258 VDD2.n28 B 0.011574f
C259 VDD2.n29 B 0.020343f
C260 VDD2.n30 B 0.010931f
C261 VDD2.n31 B 0.025838f
C262 VDD2.n32 B 0.011574f
C263 VDD2.n33 B 0.153235f
C264 VDD2.t0 B 0.042885f
C265 VDD2.n34 B 0.019378f
C266 VDD2.n35 B 0.015263f
C267 VDD2.n36 B 0.010931f
C268 VDD2.n37 B 1.69926f
C269 VDD2.n38 B 0.020343f
C270 VDD2.n39 B 0.010931f
C271 VDD2.n40 B 0.011574f
C272 VDD2.n41 B 0.025838f
C273 VDD2.n42 B 0.025838f
C274 VDD2.n43 B 0.011574f
C275 VDD2.n44 B 0.010931f
C276 VDD2.n45 B 0.020343f
C277 VDD2.n46 B 0.020343f
C278 VDD2.n47 B 0.010931f
C279 VDD2.n48 B 0.011574f
C280 VDD2.n49 B 0.025838f
C281 VDD2.n50 B 0.025838f
C282 VDD2.n51 B 0.011574f
C283 VDD2.n52 B 0.010931f
C284 VDD2.n53 B 0.020343f
C285 VDD2.n54 B 0.020343f
C286 VDD2.n55 B 0.010931f
C287 VDD2.n56 B 0.011574f
C288 VDD2.n57 B 0.025838f
C289 VDD2.n58 B 0.025838f
C290 VDD2.n59 B 0.011574f
C291 VDD2.n60 B 0.010931f
C292 VDD2.n61 B 0.020343f
C293 VDD2.n62 B 0.020343f
C294 VDD2.n63 B 0.010931f
C295 VDD2.n64 B 0.011574f
C296 VDD2.n65 B 0.025838f
C297 VDD2.n66 B 0.025838f
C298 VDD2.n67 B 0.011574f
C299 VDD2.n68 B 0.010931f
C300 VDD2.n69 B 0.020343f
C301 VDD2.n70 B 0.020343f
C302 VDD2.n71 B 0.010931f
C303 VDD2.n72 B 0.011574f
C304 VDD2.n73 B 0.025838f
C305 VDD2.n74 B 0.025838f
C306 VDD2.n75 B 0.025838f
C307 VDD2.n76 B 0.011574f
C308 VDD2.n77 B 0.010931f
C309 VDD2.n78 B 0.020343f
C310 VDD2.n79 B 0.020343f
C311 VDD2.n80 B 0.010931f
C312 VDD2.n81 B 0.011253f
C313 VDD2.n82 B 0.011253f
C314 VDD2.n83 B 0.025838f
C315 VDD2.n84 B 0.025838f
C316 VDD2.n85 B 0.011574f
C317 VDD2.n86 B 0.010931f
C318 VDD2.n87 B 0.020343f
C319 VDD2.n88 B 0.020343f
C320 VDD2.n89 B 0.010931f
C321 VDD2.n90 B 0.011574f
C322 VDD2.n91 B 0.025838f
C323 VDD2.n92 B 0.025838f
C324 VDD2.n93 B 0.011574f
C325 VDD2.n94 B 0.010931f
C326 VDD2.n95 B 0.020343f
C327 VDD2.n96 B 0.020343f
C328 VDD2.n97 B 0.010931f
C329 VDD2.n98 B 0.011574f
C330 VDD2.n99 B 0.025838f
C331 VDD2.n100 B 0.058604f
C332 VDD2.n101 B 0.011574f
C333 VDD2.n102 B 0.010931f
C334 VDD2.n103 B 0.048967f
C335 VDD2.n104 B 0.716816f
C336 VDD2.n105 B 0.030104f
C337 VDD2.n106 B 0.020343f
C338 VDD2.n107 B 0.010931f
C339 VDD2.n108 B 0.025838f
C340 VDD2.n109 B 0.011574f
C341 VDD2.n110 B 0.020343f
C342 VDD2.n111 B 0.010931f
C343 VDD2.n112 B 0.025838f
C344 VDD2.n113 B 0.011574f
C345 VDD2.n114 B 0.020343f
C346 VDD2.n115 B 0.010931f
C347 VDD2.n116 B 0.025838f
C348 VDD2.n117 B 0.011574f
C349 VDD2.n118 B 0.020343f
C350 VDD2.n119 B 0.010931f
C351 VDD2.n120 B 0.025838f
C352 VDD2.n121 B 0.025838f
C353 VDD2.n122 B 0.011574f
C354 VDD2.n123 B 0.020343f
C355 VDD2.n124 B 0.010931f
C356 VDD2.n125 B 0.025838f
C357 VDD2.n126 B 0.011574f
C358 VDD2.n127 B 0.020343f
C359 VDD2.n128 B 0.010931f
C360 VDD2.n129 B 0.025838f
C361 VDD2.n130 B 0.011574f
C362 VDD2.n131 B 0.020343f
C363 VDD2.n132 B 0.010931f
C364 VDD2.n133 B 0.025838f
C365 VDD2.n134 B 0.011574f
C366 VDD2.n135 B 0.020343f
C367 VDD2.n136 B 0.010931f
C368 VDD2.n137 B 0.025838f
C369 VDD2.n138 B 0.011574f
C370 VDD2.n139 B 0.153235f
C371 VDD2.t1 B 0.042885f
C372 VDD2.n140 B 0.019378f
C373 VDD2.n141 B 0.015263f
C374 VDD2.n142 B 0.010931f
C375 VDD2.n143 B 1.69926f
C376 VDD2.n144 B 0.020343f
C377 VDD2.n145 B 0.010931f
C378 VDD2.n146 B 0.011574f
C379 VDD2.n147 B 0.025838f
C380 VDD2.n148 B 0.025838f
C381 VDD2.n149 B 0.011574f
C382 VDD2.n150 B 0.010931f
C383 VDD2.n151 B 0.020343f
C384 VDD2.n152 B 0.020343f
C385 VDD2.n153 B 0.010931f
C386 VDD2.n154 B 0.011574f
C387 VDD2.n155 B 0.025838f
C388 VDD2.n156 B 0.025838f
C389 VDD2.n157 B 0.011574f
C390 VDD2.n158 B 0.010931f
C391 VDD2.n159 B 0.020343f
C392 VDD2.n160 B 0.020343f
C393 VDD2.n161 B 0.010931f
C394 VDD2.n162 B 0.011574f
C395 VDD2.n163 B 0.025838f
C396 VDD2.n164 B 0.025838f
C397 VDD2.n165 B 0.011574f
C398 VDD2.n166 B 0.010931f
C399 VDD2.n167 B 0.020343f
C400 VDD2.n168 B 0.020343f
C401 VDD2.n169 B 0.010931f
C402 VDD2.n170 B 0.011574f
C403 VDD2.n171 B 0.025838f
C404 VDD2.n172 B 0.025838f
C405 VDD2.n173 B 0.011574f
C406 VDD2.n174 B 0.010931f
C407 VDD2.n175 B 0.020343f
C408 VDD2.n176 B 0.020343f
C409 VDD2.n177 B 0.010931f
C410 VDD2.n178 B 0.011574f
C411 VDD2.n179 B 0.025838f
C412 VDD2.n180 B 0.025838f
C413 VDD2.n181 B 0.011574f
C414 VDD2.n182 B 0.010931f
C415 VDD2.n183 B 0.020343f
C416 VDD2.n184 B 0.020343f
C417 VDD2.n185 B 0.010931f
C418 VDD2.n186 B 0.011253f
C419 VDD2.n187 B 0.011253f
C420 VDD2.n188 B 0.025838f
C421 VDD2.n189 B 0.025838f
C422 VDD2.n190 B 0.011574f
C423 VDD2.n191 B 0.010931f
C424 VDD2.n192 B 0.020343f
C425 VDD2.n193 B 0.020343f
C426 VDD2.n194 B 0.010931f
C427 VDD2.n195 B 0.011574f
C428 VDD2.n196 B 0.025838f
C429 VDD2.n197 B 0.025838f
C430 VDD2.n198 B 0.011574f
C431 VDD2.n199 B 0.010931f
C432 VDD2.n200 B 0.020343f
C433 VDD2.n201 B 0.020343f
C434 VDD2.n202 B 0.010931f
C435 VDD2.n203 B 0.011574f
C436 VDD2.n204 B 0.025838f
C437 VDD2.n205 B 0.058604f
C438 VDD2.n206 B 0.011574f
C439 VDD2.n207 B 0.010931f
C440 VDD2.n208 B 0.048967f
C441 VDD2.n209 B 0.047156f
C442 VDD2.n210 B 2.83778f
C443 VTAIL.n0 B 0.029203f
C444 VTAIL.n1 B 0.019734f
C445 VTAIL.n2 B 0.010604f
C446 VTAIL.n3 B 0.025065f
C447 VTAIL.n4 B 0.011228f
C448 VTAIL.n5 B 0.019734f
C449 VTAIL.n6 B 0.010604f
C450 VTAIL.n7 B 0.025065f
C451 VTAIL.n8 B 0.011228f
C452 VTAIL.n9 B 0.019734f
C453 VTAIL.n10 B 0.010604f
C454 VTAIL.n11 B 0.025065f
C455 VTAIL.n12 B 0.011228f
C456 VTAIL.n13 B 0.019734f
C457 VTAIL.n14 B 0.010604f
C458 VTAIL.n15 B 0.025065f
C459 VTAIL.n16 B 0.011228f
C460 VTAIL.n17 B 0.019734f
C461 VTAIL.n18 B 0.010604f
C462 VTAIL.n19 B 0.025065f
C463 VTAIL.n20 B 0.011228f
C464 VTAIL.n21 B 0.019734f
C465 VTAIL.n22 B 0.010604f
C466 VTAIL.n23 B 0.025065f
C467 VTAIL.n24 B 0.011228f
C468 VTAIL.n25 B 0.019734f
C469 VTAIL.n26 B 0.010604f
C470 VTAIL.n27 B 0.025065f
C471 VTAIL.n28 B 0.011228f
C472 VTAIL.n29 B 0.019734f
C473 VTAIL.n30 B 0.010604f
C474 VTAIL.n31 B 0.025065f
C475 VTAIL.n32 B 0.011228f
C476 VTAIL.n33 B 0.14865f
C477 VTAIL.t0 B 0.041601f
C478 VTAIL.n34 B 0.018799f
C479 VTAIL.n35 B 0.014806f
C480 VTAIL.n36 B 0.010604f
C481 VTAIL.n37 B 1.64841f
C482 VTAIL.n38 B 0.019734f
C483 VTAIL.n39 B 0.010604f
C484 VTAIL.n40 B 0.011228f
C485 VTAIL.n41 B 0.025065f
C486 VTAIL.n42 B 0.025065f
C487 VTAIL.n43 B 0.011228f
C488 VTAIL.n44 B 0.010604f
C489 VTAIL.n45 B 0.019734f
C490 VTAIL.n46 B 0.019734f
C491 VTAIL.n47 B 0.010604f
C492 VTAIL.n48 B 0.011228f
C493 VTAIL.n49 B 0.025065f
C494 VTAIL.n50 B 0.025065f
C495 VTAIL.n51 B 0.011228f
C496 VTAIL.n52 B 0.010604f
C497 VTAIL.n53 B 0.019734f
C498 VTAIL.n54 B 0.019734f
C499 VTAIL.n55 B 0.010604f
C500 VTAIL.n56 B 0.011228f
C501 VTAIL.n57 B 0.025065f
C502 VTAIL.n58 B 0.025065f
C503 VTAIL.n59 B 0.011228f
C504 VTAIL.n60 B 0.010604f
C505 VTAIL.n61 B 0.019734f
C506 VTAIL.n62 B 0.019734f
C507 VTAIL.n63 B 0.010604f
C508 VTAIL.n64 B 0.011228f
C509 VTAIL.n65 B 0.025065f
C510 VTAIL.n66 B 0.025065f
C511 VTAIL.n67 B 0.011228f
C512 VTAIL.n68 B 0.010604f
C513 VTAIL.n69 B 0.019734f
C514 VTAIL.n70 B 0.019734f
C515 VTAIL.n71 B 0.010604f
C516 VTAIL.n72 B 0.011228f
C517 VTAIL.n73 B 0.025065f
C518 VTAIL.n74 B 0.025065f
C519 VTAIL.n75 B 0.025065f
C520 VTAIL.n76 B 0.011228f
C521 VTAIL.n77 B 0.010604f
C522 VTAIL.n78 B 0.019734f
C523 VTAIL.n79 B 0.019734f
C524 VTAIL.n80 B 0.010604f
C525 VTAIL.n81 B 0.010916f
C526 VTAIL.n82 B 0.010916f
C527 VTAIL.n83 B 0.025065f
C528 VTAIL.n84 B 0.025065f
C529 VTAIL.n85 B 0.011228f
C530 VTAIL.n86 B 0.010604f
C531 VTAIL.n87 B 0.019734f
C532 VTAIL.n88 B 0.019734f
C533 VTAIL.n89 B 0.010604f
C534 VTAIL.n90 B 0.011228f
C535 VTAIL.n91 B 0.025065f
C536 VTAIL.n92 B 0.025065f
C537 VTAIL.n93 B 0.011228f
C538 VTAIL.n94 B 0.010604f
C539 VTAIL.n95 B 0.019734f
C540 VTAIL.n96 B 0.019734f
C541 VTAIL.n97 B 0.010604f
C542 VTAIL.n98 B 0.011228f
C543 VTAIL.n99 B 0.025065f
C544 VTAIL.n100 B 0.056851f
C545 VTAIL.n101 B 0.011228f
C546 VTAIL.n102 B 0.010604f
C547 VTAIL.n103 B 0.047502f
C548 VTAIL.n104 B 0.032133f
C549 VTAIL.n105 B 1.53403f
C550 VTAIL.n106 B 0.029203f
C551 VTAIL.n107 B 0.019734f
C552 VTAIL.n108 B 0.010604f
C553 VTAIL.n109 B 0.025065f
C554 VTAIL.n110 B 0.011228f
C555 VTAIL.n111 B 0.019734f
C556 VTAIL.n112 B 0.010604f
C557 VTAIL.n113 B 0.025065f
C558 VTAIL.n114 B 0.011228f
C559 VTAIL.n115 B 0.019734f
C560 VTAIL.n116 B 0.010604f
C561 VTAIL.n117 B 0.025065f
C562 VTAIL.n118 B 0.011228f
C563 VTAIL.n119 B 0.019734f
C564 VTAIL.n120 B 0.010604f
C565 VTAIL.n121 B 0.025065f
C566 VTAIL.n122 B 0.025065f
C567 VTAIL.n123 B 0.011228f
C568 VTAIL.n124 B 0.019734f
C569 VTAIL.n125 B 0.010604f
C570 VTAIL.n126 B 0.025065f
C571 VTAIL.n127 B 0.011228f
C572 VTAIL.n128 B 0.019734f
C573 VTAIL.n129 B 0.010604f
C574 VTAIL.n130 B 0.025065f
C575 VTAIL.n131 B 0.011228f
C576 VTAIL.n132 B 0.019734f
C577 VTAIL.n133 B 0.010604f
C578 VTAIL.n134 B 0.025065f
C579 VTAIL.n135 B 0.011228f
C580 VTAIL.n136 B 0.019734f
C581 VTAIL.n137 B 0.010604f
C582 VTAIL.n138 B 0.025065f
C583 VTAIL.n139 B 0.011228f
C584 VTAIL.n140 B 0.14865f
C585 VTAIL.t2 B 0.041601f
C586 VTAIL.n141 B 0.018799f
C587 VTAIL.n142 B 0.014806f
C588 VTAIL.n143 B 0.010604f
C589 VTAIL.n144 B 1.64841f
C590 VTAIL.n145 B 0.019734f
C591 VTAIL.n146 B 0.010604f
C592 VTAIL.n147 B 0.011228f
C593 VTAIL.n148 B 0.025065f
C594 VTAIL.n149 B 0.025065f
C595 VTAIL.n150 B 0.011228f
C596 VTAIL.n151 B 0.010604f
C597 VTAIL.n152 B 0.019734f
C598 VTAIL.n153 B 0.019734f
C599 VTAIL.n154 B 0.010604f
C600 VTAIL.n155 B 0.011228f
C601 VTAIL.n156 B 0.025065f
C602 VTAIL.n157 B 0.025065f
C603 VTAIL.n158 B 0.011228f
C604 VTAIL.n159 B 0.010604f
C605 VTAIL.n160 B 0.019734f
C606 VTAIL.n161 B 0.019734f
C607 VTAIL.n162 B 0.010604f
C608 VTAIL.n163 B 0.011228f
C609 VTAIL.n164 B 0.025065f
C610 VTAIL.n165 B 0.025065f
C611 VTAIL.n166 B 0.011228f
C612 VTAIL.n167 B 0.010604f
C613 VTAIL.n168 B 0.019734f
C614 VTAIL.n169 B 0.019734f
C615 VTAIL.n170 B 0.010604f
C616 VTAIL.n171 B 0.011228f
C617 VTAIL.n172 B 0.025065f
C618 VTAIL.n173 B 0.025065f
C619 VTAIL.n174 B 0.011228f
C620 VTAIL.n175 B 0.010604f
C621 VTAIL.n176 B 0.019734f
C622 VTAIL.n177 B 0.019734f
C623 VTAIL.n178 B 0.010604f
C624 VTAIL.n179 B 0.011228f
C625 VTAIL.n180 B 0.025065f
C626 VTAIL.n181 B 0.025065f
C627 VTAIL.n182 B 0.011228f
C628 VTAIL.n183 B 0.010604f
C629 VTAIL.n184 B 0.019734f
C630 VTAIL.n185 B 0.019734f
C631 VTAIL.n186 B 0.010604f
C632 VTAIL.n187 B 0.010916f
C633 VTAIL.n188 B 0.010916f
C634 VTAIL.n189 B 0.025065f
C635 VTAIL.n190 B 0.025065f
C636 VTAIL.n191 B 0.011228f
C637 VTAIL.n192 B 0.010604f
C638 VTAIL.n193 B 0.019734f
C639 VTAIL.n194 B 0.019734f
C640 VTAIL.n195 B 0.010604f
C641 VTAIL.n196 B 0.011228f
C642 VTAIL.n197 B 0.025065f
C643 VTAIL.n198 B 0.025065f
C644 VTAIL.n199 B 0.011228f
C645 VTAIL.n200 B 0.010604f
C646 VTAIL.n201 B 0.019734f
C647 VTAIL.n202 B 0.019734f
C648 VTAIL.n203 B 0.010604f
C649 VTAIL.n204 B 0.011228f
C650 VTAIL.n205 B 0.025065f
C651 VTAIL.n206 B 0.056851f
C652 VTAIL.n207 B 0.011228f
C653 VTAIL.n208 B 0.010604f
C654 VTAIL.n209 B 0.047502f
C655 VTAIL.n210 B 0.032133f
C656 VTAIL.n211 B 1.54925f
C657 VTAIL.n212 B 0.029203f
C658 VTAIL.n213 B 0.019734f
C659 VTAIL.n214 B 0.010604f
C660 VTAIL.n215 B 0.025065f
C661 VTAIL.n216 B 0.011228f
C662 VTAIL.n217 B 0.019734f
C663 VTAIL.n218 B 0.010604f
C664 VTAIL.n219 B 0.025065f
C665 VTAIL.n220 B 0.011228f
C666 VTAIL.n221 B 0.019734f
C667 VTAIL.n222 B 0.010604f
C668 VTAIL.n223 B 0.025065f
C669 VTAIL.n224 B 0.011228f
C670 VTAIL.n225 B 0.019734f
C671 VTAIL.n226 B 0.010604f
C672 VTAIL.n227 B 0.025065f
C673 VTAIL.n228 B 0.025065f
C674 VTAIL.n229 B 0.011228f
C675 VTAIL.n230 B 0.019734f
C676 VTAIL.n231 B 0.010604f
C677 VTAIL.n232 B 0.025065f
C678 VTAIL.n233 B 0.011228f
C679 VTAIL.n234 B 0.019734f
C680 VTAIL.n235 B 0.010604f
C681 VTAIL.n236 B 0.025065f
C682 VTAIL.n237 B 0.011228f
C683 VTAIL.n238 B 0.019734f
C684 VTAIL.n239 B 0.010604f
C685 VTAIL.n240 B 0.025065f
C686 VTAIL.n241 B 0.011228f
C687 VTAIL.n242 B 0.019734f
C688 VTAIL.n243 B 0.010604f
C689 VTAIL.n244 B 0.025065f
C690 VTAIL.n245 B 0.011228f
C691 VTAIL.n246 B 0.14865f
C692 VTAIL.t1 B 0.041601f
C693 VTAIL.n247 B 0.018799f
C694 VTAIL.n248 B 0.014806f
C695 VTAIL.n249 B 0.010604f
C696 VTAIL.n250 B 1.64841f
C697 VTAIL.n251 B 0.019734f
C698 VTAIL.n252 B 0.010604f
C699 VTAIL.n253 B 0.011228f
C700 VTAIL.n254 B 0.025065f
C701 VTAIL.n255 B 0.025065f
C702 VTAIL.n256 B 0.011228f
C703 VTAIL.n257 B 0.010604f
C704 VTAIL.n258 B 0.019734f
C705 VTAIL.n259 B 0.019734f
C706 VTAIL.n260 B 0.010604f
C707 VTAIL.n261 B 0.011228f
C708 VTAIL.n262 B 0.025065f
C709 VTAIL.n263 B 0.025065f
C710 VTAIL.n264 B 0.011228f
C711 VTAIL.n265 B 0.010604f
C712 VTAIL.n266 B 0.019734f
C713 VTAIL.n267 B 0.019734f
C714 VTAIL.n268 B 0.010604f
C715 VTAIL.n269 B 0.011228f
C716 VTAIL.n270 B 0.025065f
C717 VTAIL.n271 B 0.025065f
C718 VTAIL.n272 B 0.011228f
C719 VTAIL.n273 B 0.010604f
C720 VTAIL.n274 B 0.019734f
C721 VTAIL.n275 B 0.019734f
C722 VTAIL.n276 B 0.010604f
C723 VTAIL.n277 B 0.011228f
C724 VTAIL.n278 B 0.025065f
C725 VTAIL.n279 B 0.025065f
C726 VTAIL.n280 B 0.011228f
C727 VTAIL.n281 B 0.010604f
C728 VTAIL.n282 B 0.019734f
C729 VTAIL.n283 B 0.019734f
C730 VTAIL.n284 B 0.010604f
C731 VTAIL.n285 B 0.011228f
C732 VTAIL.n286 B 0.025065f
C733 VTAIL.n287 B 0.025065f
C734 VTAIL.n288 B 0.011228f
C735 VTAIL.n289 B 0.010604f
C736 VTAIL.n290 B 0.019734f
C737 VTAIL.n291 B 0.019734f
C738 VTAIL.n292 B 0.010604f
C739 VTAIL.n293 B 0.010916f
C740 VTAIL.n294 B 0.010916f
C741 VTAIL.n295 B 0.025065f
C742 VTAIL.n296 B 0.025065f
C743 VTAIL.n297 B 0.011228f
C744 VTAIL.n298 B 0.010604f
C745 VTAIL.n299 B 0.019734f
C746 VTAIL.n300 B 0.019734f
C747 VTAIL.n301 B 0.010604f
C748 VTAIL.n302 B 0.011228f
C749 VTAIL.n303 B 0.025065f
C750 VTAIL.n304 B 0.025065f
C751 VTAIL.n305 B 0.011228f
C752 VTAIL.n306 B 0.010604f
C753 VTAIL.n307 B 0.019734f
C754 VTAIL.n308 B 0.019734f
C755 VTAIL.n309 B 0.010604f
C756 VTAIL.n310 B 0.011228f
C757 VTAIL.n311 B 0.025065f
C758 VTAIL.n312 B 0.056851f
C759 VTAIL.n313 B 0.011228f
C760 VTAIL.n314 B 0.010604f
C761 VTAIL.n315 B 0.047502f
C762 VTAIL.n316 B 0.032133f
C763 VTAIL.n317 B 1.4736f
C764 VTAIL.n318 B 0.029203f
C765 VTAIL.n319 B 0.019734f
C766 VTAIL.n320 B 0.010604f
C767 VTAIL.n321 B 0.025065f
C768 VTAIL.n322 B 0.011228f
C769 VTAIL.n323 B 0.019734f
C770 VTAIL.n324 B 0.010604f
C771 VTAIL.n325 B 0.025065f
C772 VTAIL.n326 B 0.011228f
C773 VTAIL.n327 B 0.019734f
C774 VTAIL.n328 B 0.010604f
C775 VTAIL.n329 B 0.025065f
C776 VTAIL.n330 B 0.011228f
C777 VTAIL.n331 B 0.019734f
C778 VTAIL.n332 B 0.010604f
C779 VTAIL.n333 B 0.025065f
C780 VTAIL.n334 B 0.011228f
C781 VTAIL.n335 B 0.019734f
C782 VTAIL.n336 B 0.010604f
C783 VTAIL.n337 B 0.025065f
C784 VTAIL.n338 B 0.011228f
C785 VTAIL.n339 B 0.019734f
C786 VTAIL.n340 B 0.010604f
C787 VTAIL.n341 B 0.025065f
C788 VTAIL.n342 B 0.011228f
C789 VTAIL.n343 B 0.019734f
C790 VTAIL.n344 B 0.010604f
C791 VTAIL.n345 B 0.025065f
C792 VTAIL.n346 B 0.011228f
C793 VTAIL.n347 B 0.019734f
C794 VTAIL.n348 B 0.010604f
C795 VTAIL.n349 B 0.025065f
C796 VTAIL.n350 B 0.011228f
C797 VTAIL.n351 B 0.14865f
C798 VTAIL.t3 B 0.041601f
C799 VTAIL.n352 B 0.018799f
C800 VTAIL.n353 B 0.014806f
C801 VTAIL.n354 B 0.010604f
C802 VTAIL.n355 B 1.64841f
C803 VTAIL.n356 B 0.019734f
C804 VTAIL.n357 B 0.010604f
C805 VTAIL.n358 B 0.011228f
C806 VTAIL.n359 B 0.025065f
C807 VTAIL.n360 B 0.025065f
C808 VTAIL.n361 B 0.011228f
C809 VTAIL.n362 B 0.010604f
C810 VTAIL.n363 B 0.019734f
C811 VTAIL.n364 B 0.019734f
C812 VTAIL.n365 B 0.010604f
C813 VTAIL.n366 B 0.011228f
C814 VTAIL.n367 B 0.025065f
C815 VTAIL.n368 B 0.025065f
C816 VTAIL.n369 B 0.011228f
C817 VTAIL.n370 B 0.010604f
C818 VTAIL.n371 B 0.019734f
C819 VTAIL.n372 B 0.019734f
C820 VTAIL.n373 B 0.010604f
C821 VTAIL.n374 B 0.011228f
C822 VTAIL.n375 B 0.025065f
C823 VTAIL.n376 B 0.025065f
C824 VTAIL.n377 B 0.011228f
C825 VTAIL.n378 B 0.010604f
C826 VTAIL.n379 B 0.019734f
C827 VTAIL.n380 B 0.019734f
C828 VTAIL.n381 B 0.010604f
C829 VTAIL.n382 B 0.011228f
C830 VTAIL.n383 B 0.025065f
C831 VTAIL.n384 B 0.025065f
C832 VTAIL.n385 B 0.011228f
C833 VTAIL.n386 B 0.010604f
C834 VTAIL.n387 B 0.019734f
C835 VTAIL.n388 B 0.019734f
C836 VTAIL.n389 B 0.010604f
C837 VTAIL.n390 B 0.011228f
C838 VTAIL.n391 B 0.025065f
C839 VTAIL.n392 B 0.025065f
C840 VTAIL.n393 B 0.025065f
C841 VTAIL.n394 B 0.011228f
C842 VTAIL.n395 B 0.010604f
C843 VTAIL.n396 B 0.019734f
C844 VTAIL.n397 B 0.019734f
C845 VTAIL.n398 B 0.010604f
C846 VTAIL.n399 B 0.010916f
C847 VTAIL.n400 B 0.010916f
C848 VTAIL.n401 B 0.025065f
C849 VTAIL.n402 B 0.025065f
C850 VTAIL.n403 B 0.011228f
C851 VTAIL.n404 B 0.010604f
C852 VTAIL.n405 B 0.019734f
C853 VTAIL.n406 B 0.019734f
C854 VTAIL.n407 B 0.010604f
C855 VTAIL.n408 B 0.011228f
C856 VTAIL.n409 B 0.025065f
C857 VTAIL.n410 B 0.025065f
C858 VTAIL.n411 B 0.011228f
C859 VTAIL.n412 B 0.010604f
C860 VTAIL.n413 B 0.019734f
C861 VTAIL.n414 B 0.019734f
C862 VTAIL.n415 B 0.010604f
C863 VTAIL.n416 B 0.011228f
C864 VTAIL.n417 B 0.025065f
C865 VTAIL.n418 B 0.056851f
C866 VTAIL.n419 B 0.011228f
C867 VTAIL.n420 B 0.010604f
C868 VTAIL.n421 B 0.047502f
C869 VTAIL.n422 B 0.032133f
C870 VTAIL.n423 B 1.42111f
C871 VN.t1 B 2.98348f
C872 VN.t0 B 3.19339f
.ends

