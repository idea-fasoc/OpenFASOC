* NGSPICE file created from diff_pair_sample_0738.ext - technology: sky130A

.subckt diff_pair_sample_0738 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VN.t0 VDD2.t3 w_n3290_n1504# sky130_fd_pr__pfet_01v8 ad=1.0452 pd=6.14 as=0.4422 ps=3.01 w=2.68 l=1.99
X1 VDD1.t7 VP.t0 VTAIL.t5 w_n3290_n1504# sky130_fd_pr__pfet_01v8 ad=0.4422 pd=3.01 as=1.0452 ps=6.14 w=2.68 l=1.99
X2 VDD2.t2 VN.t1 VTAIL.t14 w_n3290_n1504# sky130_fd_pr__pfet_01v8 ad=0.4422 pd=3.01 as=0.4422 ps=3.01 w=2.68 l=1.99
X3 VDD2.t1 VN.t2 VTAIL.t13 w_n3290_n1504# sky130_fd_pr__pfet_01v8 ad=0.4422 pd=3.01 as=1.0452 ps=6.14 w=2.68 l=1.99
X4 B.t11 B.t9 B.t10 w_n3290_n1504# sky130_fd_pr__pfet_01v8 ad=1.0452 pd=6.14 as=0 ps=0 w=2.68 l=1.99
X5 B.t8 B.t6 B.t7 w_n3290_n1504# sky130_fd_pr__pfet_01v8 ad=1.0452 pd=6.14 as=0 ps=0 w=2.68 l=1.99
X6 VTAIL.t12 VN.t3 VDD2.t5 w_n3290_n1504# sky130_fd_pr__pfet_01v8 ad=0.4422 pd=3.01 as=0.4422 ps=3.01 w=2.68 l=1.99
X7 VTAIL.t3 VP.t1 VDD1.t6 w_n3290_n1504# sky130_fd_pr__pfet_01v8 ad=0.4422 pd=3.01 as=0.4422 ps=3.01 w=2.68 l=1.99
X8 VDD1.t5 VP.t2 VTAIL.t4 w_n3290_n1504# sky130_fd_pr__pfet_01v8 ad=0.4422 pd=3.01 as=1.0452 ps=6.14 w=2.68 l=1.99
X9 B.t5 B.t3 B.t4 w_n3290_n1504# sky130_fd_pr__pfet_01v8 ad=1.0452 pd=6.14 as=0 ps=0 w=2.68 l=1.99
X10 VTAIL.t11 VN.t4 VDD2.t4 w_n3290_n1504# sky130_fd_pr__pfet_01v8 ad=0.4422 pd=3.01 as=0.4422 ps=3.01 w=2.68 l=1.99
X11 B.t2 B.t0 B.t1 w_n3290_n1504# sky130_fd_pr__pfet_01v8 ad=1.0452 pd=6.14 as=0 ps=0 w=2.68 l=1.99
X12 VDD2.t6 VN.t5 VTAIL.t10 w_n3290_n1504# sky130_fd_pr__pfet_01v8 ad=0.4422 pd=3.01 as=0.4422 ps=3.01 w=2.68 l=1.99
X13 VDD2.t0 VN.t6 VTAIL.t9 w_n3290_n1504# sky130_fd_pr__pfet_01v8 ad=0.4422 pd=3.01 as=1.0452 ps=6.14 w=2.68 l=1.99
X14 VTAIL.t1 VP.t3 VDD1.t4 w_n3290_n1504# sky130_fd_pr__pfet_01v8 ad=1.0452 pd=6.14 as=0.4422 ps=3.01 w=2.68 l=1.99
X15 VTAIL.t0 VP.t4 VDD1.t3 w_n3290_n1504# sky130_fd_pr__pfet_01v8 ad=0.4422 pd=3.01 as=0.4422 ps=3.01 w=2.68 l=1.99
X16 VDD1.t2 VP.t5 VTAIL.t6 w_n3290_n1504# sky130_fd_pr__pfet_01v8 ad=0.4422 pd=3.01 as=0.4422 ps=3.01 w=2.68 l=1.99
X17 VTAIL.t8 VN.t7 VDD2.t7 w_n3290_n1504# sky130_fd_pr__pfet_01v8 ad=1.0452 pd=6.14 as=0.4422 ps=3.01 w=2.68 l=1.99
X18 VTAIL.t7 VP.t6 VDD1.t1 w_n3290_n1504# sky130_fd_pr__pfet_01v8 ad=1.0452 pd=6.14 as=0.4422 ps=3.01 w=2.68 l=1.99
X19 VDD1.t0 VP.t7 VTAIL.t2 w_n3290_n1504# sky130_fd_pr__pfet_01v8 ad=0.4422 pd=3.01 as=0.4422 ps=3.01 w=2.68 l=1.99
R0 VN.n43 VN.n23 161.3
R1 VN.n42 VN.n41 161.3
R2 VN.n40 VN.n24 161.3
R3 VN.n39 VN.n38 161.3
R4 VN.n36 VN.n25 161.3
R5 VN.n35 VN.n34 161.3
R6 VN.n33 VN.n26 161.3
R7 VN.n32 VN.n31 161.3
R8 VN.n30 VN.n27 161.3
R9 VN.n20 VN.n0 161.3
R10 VN.n19 VN.n18 161.3
R11 VN.n17 VN.n1 161.3
R12 VN.n16 VN.n15 161.3
R13 VN.n13 VN.n2 161.3
R14 VN.n12 VN.n11 161.3
R15 VN.n10 VN.n3 161.3
R16 VN.n9 VN.n8 161.3
R17 VN.n7 VN.n4 161.3
R18 VN.n22 VN.n21 87.2365
R19 VN.n45 VN.n44 87.2365
R20 VN.n5 VN.t0 63.3496
R21 VN.n28 VN.t2 63.3496
R22 VN.n6 VN.n5 62.2957
R23 VN.n29 VN.n28 62.2957
R24 VN.n19 VN.n1 56.4773
R25 VN.n42 VN.n24 56.4773
R26 VN VN.n45 41.339
R27 VN.n8 VN.n3 40.4106
R28 VN.n12 VN.n3 40.4106
R29 VN.n31 VN.n26 40.4106
R30 VN.n35 VN.n26 40.4106
R31 VN.n6 VN.t1 32.4568
R32 VN.n14 VN.t3 32.4568
R33 VN.n21 VN.t6 32.4568
R34 VN.n29 VN.t4 32.4568
R35 VN.n37 VN.t5 32.4568
R36 VN.n44 VN.t7 32.4568
R37 VN.n8 VN.n7 24.3439
R38 VN.n13 VN.n12 24.3439
R39 VN.n15 VN.n1 24.3439
R40 VN.n20 VN.n19 24.3439
R41 VN.n31 VN.n30 24.3439
R42 VN.n38 VN.n24 24.3439
R43 VN.n36 VN.n35 24.3439
R44 VN.n43 VN.n42 24.3439
R45 VN.n21 VN.n20 23.3702
R46 VN.n44 VN.n43 23.3702
R47 VN.n15 VN.n14 16.554
R48 VN.n38 VN.n37 16.554
R49 VN.n28 VN.n27 12.8355
R50 VN.n5 VN.n4 12.8355
R51 VN.n7 VN.n6 7.7904
R52 VN.n14 VN.n13 7.7904
R53 VN.n30 VN.n29 7.7904
R54 VN.n37 VN.n36 7.7904
R55 VN.n45 VN.n23 0.278398
R56 VN.n22 VN.n0 0.278398
R57 VN.n41 VN.n23 0.189894
R58 VN.n41 VN.n40 0.189894
R59 VN.n40 VN.n39 0.189894
R60 VN.n39 VN.n25 0.189894
R61 VN.n34 VN.n25 0.189894
R62 VN.n34 VN.n33 0.189894
R63 VN.n33 VN.n32 0.189894
R64 VN.n32 VN.n27 0.189894
R65 VN.n9 VN.n4 0.189894
R66 VN.n10 VN.n9 0.189894
R67 VN.n11 VN.n10 0.189894
R68 VN.n11 VN.n2 0.189894
R69 VN.n16 VN.n2 0.189894
R70 VN.n17 VN.n16 0.189894
R71 VN.n18 VN.n17 0.189894
R72 VN.n18 VN.n0 0.189894
R73 VN VN.n22 0.153422
R74 VDD2.n2 VDD2.n1 152.523
R75 VDD2.n2 VDD2.n0 152.523
R76 VDD2 VDD2.n5 152.519
R77 VDD2.n4 VDD2.n3 151.577
R78 VDD2.n4 VDD2.n2 35.0256
R79 VDD2.n5 VDD2.t4 12.1292
R80 VDD2.n5 VDD2.t1 12.1292
R81 VDD2.n3 VDD2.t7 12.1292
R82 VDD2.n3 VDD2.t6 12.1292
R83 VDD2.n1 VDD2.t5 12.1292
R84 VDD2.n1 VDD2.t0 12.1292
R85 VDD2.n0 VDD2.t3 12.1292
R86 VDD2.n0 VDD2.t2 12.1292
R87 VDD2 VDD2.n4 1.05869
R88 VTAIL.n98 VTAIL.n92 756.745
R89 VTAIL.n8 VTAIL.n2 756.745
R90 VTAIL.n20 VTAIL.n14 756.745
R91 VTAIL.n34 VTAIL.n28 756.745
R92 VTAIL.n86 VTAIL.n80 756.745
R93 VTAIL.n72 VTAIL.n66 756.745
R94 VTAIL.n60 VTAIL.n54 756.745
R95 VTAIL.n46 VTAIL.n40 756.745
R96 VTAIL.n97 VTAIL.n96 585
R97 VTAIL.n99 VTAIL.n98 585
R98 VTAIL.n7 VTAIL.n6 585
R99 VTAIL.n9 VTAIL.n8 585
R100 VTAIL.n19 VTAIL.n18 585
R101 VTAIL.n21 VTAIL.n20 585
R102 VTAIL.n33 VTAIL.n32 585
R103 VTAIL.n35 VTAIL.n34 585
R104 VTAIL.n87 VTAIL.n86 585
R105 VTAIL.n85 VTAIL.n84 585
R106 VTAIL.n73 VTAIL.n72 585
R107 VTAIL.n71 VTAIL.n70 585
R108 VTAIL.n61 VTAIL.n60 585
R109 VTAIL.n59 VTAIL.n58 585
R110 VTAIL.n47 VTAIL.n46 585
R111 VTAIL.n45 VTAIL.n44 585
R112 VTAIL.n95 VTAIL.t9 357.269
R113 VTAIL.n5 VTAIL.t15 357.269
R114 VTAIL.n17 VTAIL.t4 357.269
R115 VTAIL.n31 VTAIL.t7 357.269
R116 VTAIL.n83 VTAIL.t5 357.269
R117 VTAIL.n69 VTAIL.t1 357.269
R118 VTAIL.n57 VTAIL.t13 357.269
R119 VTAIL.n43 VTAIL.t8 357.269
R120 VTAIL.n98 VTAIL.n97 171.744
R121 VTAIL.n8 VTAIL.n7 171.744
R122 VTAIL.n20 VTAIL.n19 171.744
R123 VTAIL.n34 VTAIL.n33 171.744
R124 VTAIL.n86 VTAIL.n85 171.744
R125 VTAIL.n72 VTAIL.n71 171.744
R126 VTAIL.n60 VTAIL.n59 171.744
R127 VTAIL.n46 VTAIL.n45 171.744
R128 VTAIL.n1 VTAIL.n0 134.899
R129 VTAIL.n27 VTAIL.n26 134.899
R130 VTAIL.n79 VTAIL.n78 134.899
R131 VTAIL.n53 VTAIL.n52 134.899
R132 VTAIL.n97 VTAIL.t9 85.8723
R133 VTAIL.n7 VTAIL.t15 85.8723
R134 VTAIL.n19 VTAIL.t4 85.8723
R135 VTAIL.n33 VTAIL.t7 85.8723
R136 VTAIL.n85 VTAIL.t5 85.8723
R137 VTAIL.n71 VTAIL.t1 85.8723
R138 VTAIL.n59 VTAIL.t13 85.8723
R139 VTAIL.n45 VTAIL.t8 85.8723
R140 VTAIL.n103 VTAIL.n102 30.6338
R141 VTAIL.n13 VTAIL.n12 30.6338
R142 VTAIL.n25 VTAIL.n24 30.6338
R143 VTAIL.n39 VTAIL.n38 30.6338
R144 VTAIL.n91 VTAIL.n90 30.6338
R145 VTAIL.n77 VTAIL.n76 30.6338
R146 VTAIL.n65 VTAIL.n64 30.6338
R147 VTAIL.n51 VTAIL.n50 30.6338
R148 VTAIL.n103 VTAIL.n91 16.6772
R149 VTAIL.n51 VTAIL.n39 16.6772
R150 VTAIL.n0 VTAIL.t14 12.1292
R151 VTAIL.n0 VTAIL.t12 12.1292
R152 VTAIL.n26 VTAIL.t2 12.1292
R153 VTAIL.n26 VTAIL.t3 12.1292
R154 VTAIL.n78 VTAIL.t6 12.1292
R155 VTAIL.n78 VTAIL.t0 12.1292
R156 VTAIL.n52 VTAIL.t10 12.1292
R157 VTAIL.n52 VTAIL.t11 12.1292
R158 VTAIL.n96 VTAIL.n95 10.3978
R159 VTAIL.n6 VTAIL.n5 10.3978
R160 VTAIL.n18 VTAIL.n17 10.3978
R161 VTAIL.n32 VTAIL.n31 10.3978
R162 VTAIL.n84 VTAIL.n83 10.3978
R163 VTAIL.n70 VTAIL.n69 10.3978
R164 VTAIL.n58 VTAIL.n57 10.3978
R165 VTAIL.n44 VTAIL.n43 10.3978
R166 VTAIL.n102 VTAIL.n101 9.45567
R167 VTAIL.n12 VTAIL.n11 9.45567
R168 VTAIL.n24 VTAIL.n23 9.45567
R169 VTAIL.n38 VTAIL.n37 9.45567
R170 VTAIL.n90 VTAIL.n89 9.45567
R171 VTAIL.n76 VTAIL.n75 9.45567
R172 VTAIL.n64 VTAIL.n63 9.45567
R173 VTAIL.n50 VTAIL.n49 9.45567
R174 VTAIL.n94 VTAIL.n93 9.3005
R175 VTAIL.n101 VTAIL.n100 9.3005
R176 VTAIL.n4 VTAIL.n3 9.3005
R177 VTAIL.n11 VTAIL.n10 9.3005
R178 VTAIL.n16 VTAIL.n15 9.3005
R179 VTAIL.n23 VTAIL.n22 9.3005
R180 VTAIL.n30 VTAIL.n29 9.3005
R181 VTAIL.n37 VTAIL.n36 9.3005
R182 VTAIL.n82 VTAIL.n81 9.3005
R183 VTAIL.n89 VTAIL.n88 9.3005
R184 VTAIL.n75 VTAIL.n74 9.3005
R185 VTAIL.n68 VTAIL.n67 9.3005
R186 VTAIL.n63 VTAIL.n62 9.3005
R187 VTAIL.n56 VTAIL.n55 9.3005
R188 VTAIL.n49 VTAIL.n48 9.3005
R189 VTAIL.n42 VTAIL.n41 9.3005
R190 VTAIL.n102 VTAIL.n92 8.92171
R191 VTAIL.n12 VTAIL.n2 8.92171
R192 VTAIL.n24 VTAIL.n14 8.92171
R193 VTAIL.n38 VTAIL.n28 8.92171
R194 VTAIL.n90 VTAIL.n80 8.92171
R195 VTAIL.n76 VTAIL.n66 8.92171
R196 VTAIL.n64 VTAIL.n54 8.92171
R197 VTAIL.n50 VTAIL.n40 8.92171
R198 VTAIL.n100 VTAIL.n99 8.14595
R199 VTAIL.n10 VTAIL.n9 8.14595
R200 VTAIL.n22 VTAIL.n21 8.14595
R201 VTAIL.n36 VTAIL.n35 8.14595
R202 VTAIL.n88 VTAIL.n87 8.14595
R203 VTAIL.n74 VTAIL.n73 8.14595
R204 VTAIL.n62 VTAIL.n61 8.14595
R205 VTAIL.n48 VTAIL.n47 8.14595
R206 VTAIL.n96 VTAIL.n94 7.3702
R207 VTAIL.n6 VTAIL.n4 7.3702
R208 VTAIL.n18 VTAIL.n16 7.3702
R209 VTAIL.n32 VTAIL.n30 7.3702
R210 VTAIL.n84 VTAIL.n82 7.3702
R211 VTAIL.n70 VTAIL.n68 7.3702
R212 VTAIL.n58 VTAIL.n56 7.3702
R213 VTAIL.n44 VTAIL.n42 7.3702
R214 VTAIL.n99 VTAIL.n94 5.81868
R215 VTAIL.n9 VTAIL.n4 5.81868
R216 VTAIL.n21 VTAIL.n16 5.81868
R217 VTAIL.n35 VTAIL.n30 5.81868
R218 VTAIL.n87 VTAIL.n82 5.81868
R219 VTAIL.n73 VTAIL.n68 5.81868
R220 VTAIL.n61 VTAIL.n56 5.81868
R221 VTAIL.n47 VTAIL.n42 5.81868
R222 VTAIL.n100 VTAIL.n92 5.04292
R223 VTAIL.n10 VTAIL.n2 5.04292
R224 VTAIL.n22 VTAIL.n14 5.04292
R225 VTAIL.n36 VTAIL.n28 5.04292
R226 VTAIL.n88 VTAIL.n80 5.04292
R227 VTAIL.n74 VTAIL.n66 5.04292
R228 VTAIL.n62 VTAIL.n54 5.04292
R229 VTAIL.n48 VTAIL.n40 5.04292
R230 VTAIL.n95 VTAIL.n93 2.74506
R231 VTAIL.n5 VTAIL.n3 2.74506
R232 VTAIL.n17 VTAIL.n15 2.74506
R233 VTAIL.n31 VTAIL.n29 2.74506
R234 VTAIL.n83 VTAIL.n81 2.74506
R235 VTAIL.n69 VTAIL.n67 2.74506
R236 VTAIL.n57 VTAIL.n55 2.74506
R237 VTAIL.n43 VTAIL.n41 2.74506
R238 VTAIL.n53 VTAIL.n51 2.0005
R239 VTAIL.n65 VTAIL.n53 2.0005
R240 VTAIL.n79 VTAIL.n77 2.0005
R241 VTAIL.n91 VTAIL.n79 2.0005
R242 VTAIL.n39 VTAIL.n27 2.0005
R243 VTAIL.n27 VTAIL.n25 2.0005
R244 VTAIL.n13 VTAIL.n1 2.0005
R245 VTAIL VTAIL.n103 1.94231
R246 VTAIL.n77 VTAIL.n65 0.470328
R247 VTAIL.n25 VTAIL.n13 0.470328
R248 VTAIL.n101 VTAIL.n93 0.155672
R249 VTAIL.n11 VTAIL.n3 0.155672
R250 VTAIL.n23 VTAIL.n15 0.155672
R251 VTAIL.n37 VTAIL.n29 0.155672
R252 VTAIL.n89 VTAIL.n81 0.155672
R253 VTAIL.n75 VTAIL.n67 0.155672
R254 VTAIL.n63 VTAIL.n55 0.155672
R255 VTAIL.n49 VTAIL.n41 0.155672
R256 VTAIL VTAIL.n1 0.0586897
R257 VP.n14 VP.n11 161.3
R258 VP.n16 VP.n15 161.3
R259 VP.n17 VP.n10 161.3
R260 VP.n19 VP.n18 161.3
R261 VP.n20 VP.n9 161.3
R262 VP.n23 VP.n22 161.3
R263 VP.n24 VP.n8 161.3
R264 VP.n26 VP.n25 161.3
R265 VP.n27 VP.n7 161.3
R266 VP.n52 VP.n0 161.3
R267 VP.n51 VP.n50 161.3
R268 VP.n49 VP.n1 161.3
R269 VP.n48 VP.n47 161.3
R270 VP.n45 VP.n2 161.3
R271 VP.n44 VP.n43 161.3
R272 VP.n42 VP.n3 161.3
R273 VP.n41 VP.n40 161.3
R274 VP.n39 VP.n4 161.3
R275 VP.n37 VP.n36 161.3
R276 VP.n35 VP.n5 161.3
R277 VP.n34 VP.n33 161.3
R278 VP.n32 VP.n6 161.3
R279 VP.n31 VP.n30 87.2365
R280 VP.n54 VP.n53 87.2365
R281 VP.n29 VP.n28 87.2365
R282 VP.n12 VP.t3 63.3496
R283 VP.n13 VP.n12 62.2957
R284 VP.n33 VP.n5 56.4773
R285 VP.n51 VP.n1 56.4773
R286 VP.n26 VP.n8 56.4773
R287 VP.n30 VP.n29 41.0601
R288 VP.n40 VP.n3 40.4106
R289 VP.n44 VP.n3 40.4106
R290 VP.n19 VP.n10 40.4106
R291 VP.n15 VP.n10 40.4106
R292 VP.n31 VP.t6 32.4568
R293 VP.n38 VP.t7 32.4568
R294 VP.n46 VP.t1 32.4568
R295 VP.n53 VP.t2 32.4568
R296 VP.n28 VP.t0 32.4568
R297 VP.n21 VP.t4 32.4568
R298 VP.n13 VP.t5 32.4568
R299 VP.n33 VP.n32 24.3439
R300 VP.n37 VP.n5 24.3439
R301 VP.n40 VP.n39 24.3439
R302 VP.n45 VP.n44 24.3439
R303 VP.n47 VP.n1 24.3439
R304 VP.n52 VP.n51 24.3439
R305 VP.n27 VP.n26 24.3439
R306 VP.n20 VP.n19 24.3439
R307 VP.n22 VP.n8 24.3439
R308 VP.n15 VP.n14 24.3439
R309 VP.n32 VP.n31 23.3702
R310 VP.n53 VP.n52 23.3702
R311 VP.n28 VP.n27 23.3702
R312 VP.n38 VP.n37 16.554
R313 VP.n47 VP.n46 16.554
R314 VP.n22 VP.n21 16.554
R315 VP.n12 VP.n11 12.8355
R316 VP.n39 VP.n38 7.7904
R317 VP.n46 VP.n45 7.7904
R318 VP.n21 VP.n20 7.7904
R319 VP.n14 VP.n13 7.7904
R320 VP.n29 VP.n7 0.278398
R321 VP.n30 VP.n6 0.278398
R322 VP.n54 VP.n0 0.278398
R323 VP.n16 VP.n11 0.189894
R324 VP.n17 VP.n16 0.189894
R325 VP.n18 VP.n17 0.189894
R326 VP.n18 VP.n9 0.189894
R327 VP.n23 VP.n9 0.189894
R328 VP.n24 VP.n23 0.189894
R329 VP.n25 VP.n24 0.189894
R330 VP.n25 VP.n7 0.189894
R331 VP.n34 VP.n6 0.189894
R332 VP.n35 VP.n34 0.189894
R333 VP.n36 VP.n35 0.189894
R334 VP.n36 VP.n4 0.189894
R335 VP.n41 VP.n4 0.189894
R336 VP.n42 VP.n41 0.189894
R337 VP.n43 VP.n42 0.189894
R338 VP.n43 VP.n2 0.189894
R339 VP.n48 VP.n2 0.189894
R340 VP.n49 VP.n48 0.189894
R341 VP.n50 VP.n49 0.189894
R342 VP.n50 VP.n0 0.189894
R343 VP VP.n54 0.153422
R344 VDD1 VDD1.n0 152.636
R345 VDD1.n3 VDD1.n2 152.523
R346 VDD1.n3 VDD1.n1 152.523
R347 VDD1.n5 VDD1.n4 151.577
R348 VDD1.n5 VDD1.n3 35.6087
R349 VDD1.n4 VDD1.t3 12.1292
R350 VDD1.n4 VDD1.t7 12.1292
R351 VDD1.n0 VDD1.t4 12.1292
R352 VDD1.n0 VDD1.t2 12.1292
R353 VDD1.n2 VDD1.t6 12.1292
R354 VDD1.n2 VDD1.t5 12.1292
R355 VDD1.n1 VDD1.t1 12.1292
R356 VDD1.n1 VDD1.t0 12.1292
R357 VDD1 VDD1.n5 0.94231
R358 B.n381 B.n46 585
R359 B.n383 B.n382 585
R360 B.n384 B.n45 585
R361 B.n386 B.n385 585
R362 B.n387 B.n44 585
R363 B.n389 B.n388 585
R364 B.n390 B.n43 585
R365 B.n392 B.n391 585
R366 B.n393 B.n42 585
R367 B.n395 B.n394 585
R368 B.n396 B.n41 585
R369 B.n398 B.n397 585
R370 B.n399 B.n40 585
R371 B.n401 B.n400 585
R372 B.n403 B.n37 585
R373 B.n405 B.n404 585
R374 B.n406 B.n36 585
R375 B.n408 B.n407 585
R376 B.n409 B.n35 585
R377 B.n411 B.n410 585
R378 B.n412 B.n34 585
R379 B.n414 B.n413 585
R380 B.n415 B.n33 585
R381 B.n417 B.n416 585
R382 B.n419 B.n418 585
R383 B.n420 B.n29 585
R384 B.n422 B.n421 585
R385 B.n423 B.n28 585
R386 B.n425 B.n424 585
R387 B.n426 B.n27 585
R388 B.n428 B.n427 585
R389 B.n429 B.n26 585
R390 B.n431 B.n430 585
R391 B.n432 B.n25 585
R392 B.n434 B.n433 585
R393 B.n435 B.n24 585
R394 B.n437 B.n436 585
R395 B.n438 B.n23 585
R396 B.n380 B.n379 585
R397 B.n378 B.n47 585
R398 B.n377 B.n376 585
R399 B.n375 B.n48 585
R400 B.n374 B.n373 585
R401 B.n372 B.n49 585
R402 B.n371 B.n370 585
R403 B.n369 B.n50 585
R404 B.n368 B.n367 585
R405 B.n366 B.n51 585
R406 B.n365 B.n364 585
R407 B.n363 B.n52 585
R408 B.n362 B.n361 585
R409 B.n360 B.n53 585
R410 B.n359 B.n358 585
R411 B.n357 B.n54 585
R412 B.n356 B.n355 585
R413 B.n354 B.n55 585
R414 B.n353 B.n352 585
R415 B.n351 B.n56 585
R416 B.n350 B.n349 585
R417 B.n348 B.n57 585
R418 B.n347 B.n346 585
R419 B.n345 B.n58 585
R420 B.n344 B.n343 585
R421 B.n342 B.n59 585
R422 B.n341 B.n340 585
R423 B.n339 B.n60 585
R424 B.n338 B.n337 585
R425 B.n336 B.n61 585
R426 B.n335 B.n334 585
R427 B.n333 B.n62 585
R428 B.n332 B.n331 585
R429 B.n330 B.n63 585
R430 B.n329 B.n328 585
R431 B.n327 B.n64 585
R432 B.n326 B.n325 585
R433 B.n324 B.n65 585
R434 B.n323 B.n322 585
R435 B.n321 B.n66 585
R436 B.n320 B.n319 585
R437 B.n318 B.n67 585
R438 B.n317 B.n316 585
R439 B.n315 B.n68 585
R440 B.n314 B.n313 585
R441 B.n312 B.n69 585
R442 B.n311 B.n310 585
R443 B.n309 B.n70 585
R444 B.n308 B.n307 585
R445 B.n306 B.n71 585
R446 B.n305 B.n304 585
R447 B.n303 B.n72 585
R448 B.n302 B.n301 585
R449 B.n300 B.n73 585
R450 B.n299 B.n298 585
R451 B.n297 B.n74 585
R452 B.n296 B.n295 585
R453 B.n294 B.n75 585
R454 B.n293 B.n292 585
R455 B.n291 B.n76 585
R456 B.n290 B.n289 585
R457 B.n288 B.n77 585
R458 B.n287 B.n286 585
R459 B.n285 B.n78 585
R460 B.n284 B.n283 585
R461 B.n282 B.n79 585
R462 B.n281 B.n280 585
R463 B.n279 B.n80 585
R464 B.n278 B.n277 585
R465 B.n276 B.n81 585
R466 B.n275 B.n274 585
R467 B.n273 B.n82 585
R468 B.n272 B.n271 585
R469 B.n270 B.n83 585
R470 B.n269 B.n268 585
R471 B.n267 B.n84 585
R472 B.n266 B.n265 585
R473 B.n264 B.n85 585
R474 B.n263 B.n262 585
R475 B.n261 B.n86 585
R476 B.n260 B.n259 585
R477 B.n258 B.n87 585
R478 B.n257 B.n256 585
R479 B.n255 B.n88 585
R480 B.n254 B.n253 585
R481 B.n195 B.n112 585
R482 B.n197 B.n196 585
R483 B.n198 B.n111 585
R484 B.n200 B.n199 585
R485 B.n201 B.n110 585
R486 B.n203 B.n202 585
R487 B.n204 B.n109 585
R488 B.n206 B.n205 585
R489 B.n207 B.n108 585
R490 B.n209 B.n208 585
R491 B.n210 B.n107 585
R492 B.n212 B.n211 585
R493 B.n213 B.n106 585
R494 B.n215 B.n214 585
R495 B.n217 B.n103 585
R496 B.n219 B.n218 585
R497 B.n220 B.n102 585
R498 B.n222 B.n221 585
R499 B.n223 B.n101 585
R500 B.n225 B.n224 585
R501 B.n226 B.n100 585
R502 B.n228 B.n227 585
R503 B.n229 B.n99 585
R504 B.n231 B.n230 585
R505 B.n233 B.n232 585
R506 B.n234 B.n95 585
R507 B.n236 B.n235 585
R508 B.n237 B.n94 585
R509 B.n239 B.n238 585
R510 B.n240 B.n93 585
R511 B.n242 B.n241 585
R512 B.n243 B.n92 585
R513 B.n245 B.n244 585
R514 B.n246 B.n91 585
R515 B.n248 B.n247 585
R516 B.n249 B.n90 585
R517 B.n251 B.n250 585
R518 B.n252 B.n89 585
R519 B.n194 B.n193 585
R520 B.n192 B.n113 585
R521 B.n191 B.n190 585
R522 B.n189 B.n114 585
R523 B.n188 B.n187 585
R524 B.n186 B.n115 585
R525 B.n185 B.n184 585
R526 B.n183 B.n116 585
R527 B.n182 B.n181 585
R528 B.n180 B.n117 585
R529 B.n179 B.n178 585
R530 B.n177 B.n118 585
R531 B.n176 B.n175 585
R532 B.n174 B.n119 585
R533 B.n173 B.n172 585
R534 B.n171 B.n120 585
R535 B.n170 B.n169 585
R536 B.n168 B.n121 585
R537 B.n167 B.n166 585
R538 B.n165 B.n122 585
R539 B.n164 B.n163 585
R540 B.n162 B.n123 585
R541 B.n161 B.n160 585
R542 B.n159 B.n124 585
R543 B.n158 B.n157 585
R544 B.n156 B.n125 585
R545 B.n155 B.n154 585
R546 B.n153 B.n126 585
R547 B.n152 B.n151 585
R548 B.n150 B.n127 585
R549 B.n149 B.n148 585
R550 B.n147 B.n128 585
R551 B.n146 B.n145 585
R552 B.n144 B.n129 585
R553 B.n143 B.n142 585
R554 B.n141 B.n130 585
R555 B.n140 B.n139 585
R556 B.n138 B.n131 585
R557 B.n137 B.n136 585
R558 B.n135 B.n132 585
R559 B.n134 B.n133 585
R560 B.n2 B.n0 585
R561 B.n501 B.n1 585
R562 B.n500 B.n499 585
R563 B.n498 B.n3 585
R564 B.n497 B.n496 585
R565 B.n495 B.n4 585
R566 B.n494 B.n493 585
R567 B.n492 B.n5 585
R568 B.n491 B.n490 585
R569 B.n489 B.n6 585
R570 B.n488 B.n487 585
R571 B.n486 B.n7 585
R572 B.n485 B.n484 585
R573 B.n483 B.n8 585
R574 B.n482 B.n481 585
R575 B.n480 B.n9 585
R576 B.n479 B.n478 585
R577 B.n477 B.n10 585
R578 B.n476 B.n475 585
R579 B.n474 B.n11 585
R580 B.n473 B.n472 585
R581 B.n471 B.n12 585
R582 B.n470 B.n469 585
R583 B.n468 B.n13 585
R584 B.n467 B.n466 585
R585 B.n465 B.n14 585
R586 B.n464 B.n463 585
R587 B.n462 B.n15 585
R588 B.n461 B.n460 585
R589 B.n459 B.n16 585
R590 B.n458 B.n457 585
R591 B.n456 B.n17 585
R592 B.n455 B.n454 585
R593 B.n453 B.n18 585
R594 B.n452 B.n451 585
R595 B.n450 B.n19 585
R596 B.n449 B.n448 585
R597 B.n447 B.n20 585
R598 B.n446 B.n445 585
R599 B.n444 B.n21 585
R600 B.n443 B.n442 585
R601 B.n441 B.n22 585
R602 B.n440 B.n439 585
R603 B.n503 B.n502 585
R604 B.n195 B.n194 535.745
R605 B.n440 B.n23 535.745
R606 B.n254 B.n89 535.745
R607 B.n381 B.n380 535.745
R608 B.n96 B.t2 272.736
R609 B.n38 B.t7 272.736
R610 B.n104 B.t11 272.736
R611 B.n30 B.t4 272.736
R612 B.n96 B.t0 239.351
R613 B.n104 B.t9 239.351
R614 B.n30 B.t3 239.351
R615 B.n38 B.t6 239.351
R616 B.n97 B.t1 227.743
R617 B.n39 B.t8 227.743
R618 B.n105 B.t10 227.743
R619 B.n31 B.t5 227.743
R620 B.n194 B.n113 163.367
R621 B.n190 B.n113 163.367
R622 B.n190 B.n189 163.367
R623 B.n189 B.n188 163.367
R624 B.n188 B.n115 163.367
R625 B.n184 B.n115 163.367
R626 B.n184 B.n183 163.367
R627 B.n183 B.n182 163.367
R628 B.n182 B.n117 163.367
R629 B.n178 B.n117 163.367
R630 B.n178 B.n177 163.367
R631 B.n177 B.n176 163.367
R632 B.n176 B.n119 163.367
R633 B.n172 B.n119 163.367
R634 B.n172 B.n171 163.367
R635 B.n171 B.n170 163.367
R636 B.n170 B.n121 163.367
R637 B.n166 B.n121 163.367
R638 B.n166 B.n165 163.367
R639 B.n165 B.n164 163.367
R640 B.n164 B.n123 163.367
R641 B.n160 B.n123 163.367
R642 B.n160 B.n159 163.367
R643 B.n159 B.n158 163.367
R644 B.n158 B.n125 163.367
R645 B.n154 B.n125 163.367
R646 B.n154 B.n153 163.367
R647 B.n153 B.n152 163.367
R648 B.n152 B.n127 163.367
R649 B.n148 B.n127 163.367
R650 B.n148 B.n147 163.367
R651 B.n147 B.n146 163.367
R652 B.n146 B.n129 163.367
R653 B.n142 B.n129 163.367
R654 B.n142 B.n141 163.367
R655 B.n141 B.n140 163.367
R656 B.n140 B.n131 163.367
R657 B.n136 B.n131 163.367
R658 B.n136 B.n135 163.367
R659 B.n135 B.n134 163.367
R660 B.n134 B.n2 163.367
R661 B.n502 B.n2 163.367
R662 B.n502 B.n501 163.367
R663 B.n501 B.n500 163.367
R664 B.n500 B.n3 163.367
R665 B.n496 B.n3 163.367
R666 B.n496 B.n495 163.367
R667 B.n495 B.n494 163.367
R668 B.n494 B.n5 163.367
R669 B.n490 B.n5 163.367
R670 B.n490 B.n489 163.367
R671 B.n489 B.n488 163.367
R672 B.n488 B.n7 163.367
R673 B.n484 B.n7 163.367
R674 B.n484 B.n483 163.367
R675 B.n483 B.n482 163.367
R676 B.n482 B.n9 163.367
R677 B.n478 B.n9 163.367
R678 B.n478 B.n477 163.367
R679 B.n477 B.n476 163.367
R680 B.n476 B.n11 163.367
R681 B.n472 B.n11 163.367
R682 B.n472 B.n471 163.367
R683 B.n471 B.n470 163.367
R684 B.n470 B.n13 163.367
R685 B.n466 B.n13 163.367
R686 B.n466 B.n465 163.367
R687 B.n465 B.n464 163.367
R688 B.n464 B.n15 163.367
R689 B.n460 B.n15 163.367
R690 B.n460 B.n459 163.367
R691 B.n459 B.n458 163.367
R692 B.n458 B.n17 163.367
R693 B.n454 B.n17 163.367
R694 B.n454 B.n453 163.367
R695 B.n453 B.n452 163.367
R696 B.n452 B.n19 163.367
R697 B.n448 B.n19 163.367
R698 B.n448 B.n447 163.367
R699 B.n447 B.n446 163.367
R700 B.n446 B.n21 163.367
R701 B.n442 B.n21 163.367
R702 B.n442 B.n441 163.367
R703 B.n441 B.n440 163.367
R704 B.n196 B.n195 163.367
R705 B.n196 B.n111 163.367
R706 B.n200 B.n111 163.367
R707 B.n201 B.n200 163.367
R708 B.n202 B.n201 163.367
R709 B.n202 B.n109 163.367
R710 B.n206 B.n109 163.367
R711 B.n207 B.n206 163.367
R712 B.n208 B.n207 163.367
R713 B.n208 B.n107 163.367
R714 B.n212 B.n107 163.367
R715 B.n213 B.n212 163.367
R716 B.n214 B.n213 163.367
R717 B.n214 B.n103 163.367
R718 B.n219 B.n103 163.367
R719 B.n220 B.n219 163.367
R720 B.n221 B.n220 163.367
R721 B.n221 B.n101 163.367
R722 B.n225 B.n101 163.367
R723 B.n226 B.n225 163.367
R724 B.n227 B.n226 163.367
R725 B.n227 B.n99 163.367
R726 B.n231 B.n99 163.367
R727 B.n232 B.n231 163.367
R728 B.n232 B.n95 163.367
R729 B.n236 B.n95 163.367
R730 B.n237 B.n236 163.367
R731 B.n238 B.n237 163.367
R732 B.n238 B.n93 163.367
R733 B.n242 B.n93 163.367
R734 B.n243 B.n242 163.367
R735 B.n244 B.n243 163.367
R736 B.n244 B.n91 163.367
R737 B.n248 B.n91 163.367
R738 B.n249 B.n248 163.367
R739 B.n250 B.n249 163.367
R740 B.n250 B.n89 163.367
R741 B.n255 B.n254 163.367
R742 B.n256 B.n255 163.367
R743 B.n256 B.n87 163.367
R744 B.n260 B.n87 163.367
R745 B.n261 B.n260 163.367
R746 B.n262 B.n261 163.367
R747 B.n262 B.n85 163.367
R748 B.n266 B.n85 163.367
R749 B.n267 B.n266 163.367
R750 B.n268 B.n267 163.367
R751 B.n268 B.n83 163.367
R752 B.n272 B.n83 163.367
R753 B.n273 B.n272 163.367
R754 B.n274 B.n273 163.367
R755 B.n274 B.n81 163.367
R756 B.n278 B.n81 163.367
R757 B.n279 B.n278 163.367
R758 B.n280 B.n279 163.367
R759 B.n280 B.n79 163.367
R760 B.n284 B.n79 163.367
R761 B.n285 B.n284 163.367
R762 B.n286 B.n285 163.367
R763 B.n286 B.n77 163.367
R764 B.n290 B.n77 163.367
R765 B.n291 B.n290 163.367
R766 B.n292 B.n291 163.367
R767 B.n292 B.n75 163.367
R768 B.n296 B.n75 163.367
R769 B.n297 B.n296 163.367
R770 B.n298 B.n297 163.367
R771 B.n298 B.n73 163.367
R772 B.n302 B.n73 163.367
R773 B.n303 B.n302 163.367
R774 B.n304 B.n303 163.367
R775 B.n304 B.n71 163.367
R776 B.n308 B.n71 163.367
R777 B.n309 B.n308 163.367
R778 B.n310 B.n309 163.367
R779 B.n310 B.n69 163.367
R780 B.n314 B.n69 163.367
R781 B.n315 B.n314 163.367
R782 B.n316 B.n315 163.367
R783 B.n316 B.n67 163.367
R784 B.n320 B.n67 163.367
R785 B.n321 B.n320 163.367
R786 B.n322 B.n321 163.367
R787 B.n322 B.n65 163.367
R788 B.n326 B.n65 163.367
R789 B.n327 B.n326 163.367
R790 B.n328 B.n327 163.367
R791 B.n328 B.n63 163.367
R792 B.n332 B.n63 163.367
R793 B.n333 B.n332 163.367
R794 B.n334 B.n333 163.367
R795 B.n334 B.n61 163.367
R796 B.n338 B.n61 163.367
R797 B.n339 B.n338 163.367
R798 B.n340 B.n339 163.367
R799 B.n340 B.n59 163.367
R800 B.n344 B.n59 163.367
R801 B.n345 B.n344 163.367
R802 B.n346 B.n345 163.367
R803 B.n346 B.n57 163.367
R804 B.n350 B.n57 163.367
R805 B.n351 B.n350 163.367
R806 B.n352 B.n351 163.367
R807 B.n352 B.n55 163.367
R808 B.n356 B.n55 163.367
R809 B.n357 B.n356 163.367
R810 B.n358 B.n357 163.367
R811 B.n358 B.n53 163.367
R812 B.n362 B.n53 163.367
R813 B.n363 B.n362 163.367
R814 B.n364 B.n363 163.367
R815 B.n364 B.n51 163.367
R816 B.n368 B.n51 163.367
R817 B.n369 B.n368 163.367
R818 B.n370 B.n369 163.367
R819 B.n370 B.n49 163.367
R820 B.n374 B.n49 163.367
R821 B.n375 B.n374 163.367
R822 B.n376 B.n375 163.367
R823 B.n376 B.n47 163.367
R824 B.n380 B.n47 163.367
R825 B.n436 B.n23 163.367
R826 B.n436 B.n435 163.367
R827 B.n435 B.n434 163.367
R828 B.n434 B.n25 163.367
R829 B.n430 B.n25 163.367
R830 B.n430 B.n429 163.367
R831 B.n429 B.n428 163.367
R832 B.n428 B.n27 163.367
R833 B.n424 B.n27 163.367
R834 B.n424 B.n423 163.367
R835 B.n423 B.n422 163.367
R836 B.n422 B.n29 163.367
R837 B.n418 B.n29 163.367
R838 B.n418 B.n417 163.367
R839 B.n417 B.n33 163.367
R840 B.n413 B.n33 163.367
R841 B.n413 B.n412 163.367
R842 B.n412 B.n411 163.367
R843 B.n411 B.n35 163.367
R844 B.n407 B.n35 163.367
R845 B.n407 B.n406 163.367
R846 B.n406 B.n405 163.367
R847 B.n405 B.n37 163.367
R848 B.n400 B.n37 163.367
R849 B.n400 B.n399 163.367
R850 B.n399 B.n398 163.367
R851 B.n398 B.n41 163.367
R852 B.n394 B.n41 163.367
R853 B.n394 B.n393 163.367
R854 B.n393 B.n392 163.367
R855 B.n392 B.n43 163.367
R856 B.n388 B.n43 163.367
R857 B.n388 B.n387 163.367
R858 B.n387 B.n386 163.367
R859 B.n386 B.n45 163.367
R860 B.n382 B.n45 163.367
R861 B.n382 B.n381 163.367
R862 B.n98 B.n97 59.5399
R863 B.n216 B.n105 59.5399
R864 B.n32 B.n31 59.5399
R865 B.n402 B.n39 59.5399
R866 B.n97 B.n96 44.9944
R867 B.n105 B.n104 44.9944
R868 B.n31 B.n30 44.9944
R869 B.n39 B.n38 44.9944
R870 B.n439 B.n438 34.8103
R871 B.n379 B.n46 34.8103
R872 B.n253 B.n252 34.8103
R873 B.n193 B.n112 34.8103
R874 B B.n503 18.0485
R875 B.n438 B.n437 10.6151
R876 B.n437 B.n24 10.6151
R877 B.n433 B.n24 10.6151
R878 B.n433 B.n432 10.6151
R879 B.n432 B.n431 10.6151
R880 B.n431 B.n26 10.6151
R881 B.n427 B.n26 10.6151
R882 B.n427 B.n426 10.6151
R883 B.n426 B.n425 10.6151
R884 B.n425 B.n28 10.6151
R885 B.n421 B.n28 10.6151
R886 B.n421 B.n420 10.6151
R887 B.n420 B.n419 10.6151
R888 B.n416 B.n415 10.6151
R889 B.n415 B.n414 10.6151
R890 B.n414 B.n34 10.6151
R891 B.n410 B.n34 10.6151
R892 B.n410 B.n409 10.6151
R893 B.n409 B.n408 10.6151
R894 B.n408 B.n36 10.6151
R895 B.n404 B.n36 10.6151
R896 B.n404 B.n403 10.6151
R897 B.n401 B.n40 10.6151
R898 B.n397 B.n40 10.6151
R899 B.n397 B.n396 10.6151
R900 B.n396 B.n395 10.6151
R901 B.n395 B.n42 10.6151
R902 B.n391 B.n42 10.6151
R903 B.n391 B.n390 10.6151
R904 B.n390 B.n389 10.6151
R905 B.n389 B.n44 10.6151
R906 B.n385 B.n44 10.6151
R907 B.n385 B.n384 10.6151
R908 B.n384 B.n383 10.6151
R909 B.n383 B.n46 10.6151
R910 B.n253 B.n88 10.6151
R911 B.n257 B.n88 10.6151
R912 B.n258 B.n257 10.6151
R913 B.n259 B.n258 10.6151
R914 B.n259 B.n86 10.6151
R915 B.n263 B.n86 10.6151
R916 B.n264 B.n263 10.6151
R917 B.n265 B.n264 10.6151
R918 B.n265 B.n84 10.6151
R919 B.n269 B.n84 10.6151
R920 B.n270 B.n269 10.6151
R921 B.n271 B.n270 10.6151
R922 B.n271 B.n82 10.6151
R923 B.n275 B.n82 10.6151
R924 B.n276 B.n275 10.6151
R925 B.n277 B.n276 10.6151
R926 B.n277 B.n80 10.6151
R927 B.n281 B.n80 10.6151
R928 B.n282 B.n281 10.6151
R929 B.n283 B.n282 10.6151
R930 B.n283 B.n78 10.6151
R931 B.n287 B.n78 10.6151
R932 B.n288 B.n287 10.6151
R933 B.n289 B.n288 10.6151
R934 B.n289 B.n76 10.6151
R935 B.n293 B.n76 10.6151
R936 B.n294 B.n293 10.6151
R937 B.n295 B.n294 10.6151
R938 B.n295 B.n74 10.6151
R939 B.n299 B.n74 10.6151
R940 B.n300 B.n299 10.6151
R941 B.n301 B.n300 10.6151
R942 B.n301 B.n72 10.6151
R943 B.n305 B.n72 10.6151
R944 B.n306 B.n305 10.6151
R945 B.n307 B.n306 10.6151
R946 B.n307 B.n70 10.6151
R947 B.n311 B.n70 10.6151
R948 B.n312 B.n311 10.6151
R949 B.n313 B.n312 10.6151
R950 B.n313 B.n68 10.6151
R951 B.n317 B.n68 10.6151
R952 B.n318 B.n317 10.6151
R953 B.n319 B.n318 10.6151
R954 B.n319 B.n66 10.6151
R955 B.n323 B.n66 10.6151
R956 B.n324 B.n323 10.6151
R957 B.n325 B.n324 10.6151
R958 B.n325 B.n64 10.6151
R959 B.n329 B.n64 10.6151
R960 B.n330 B.n329 10.6151
R961 B.n331 B.n330 10.6151
R962 B.n331 B.n62 10.6151
R963 B.n335 B.n62 10.6151
R964 B.n336 B.n335 10.6151
R965 B.n337 B.n336 10.6151
R966 B.n337 B.n60 10.6151
R967 B.n341 B.n60 10.6151
R968 B.n342 B.n341 10.6151
R969 B.n343 B.n342 10.6151
R970 B.n343 B.n58 10.6151
R971 B.n347 B.n58 10.6151
R972 B.n348 B.n347 10.6151
R973 B.n349 B.n348 10.6151
R974 B.n349 B.n56 10.6151
R975 B.n353 B.n56 10.6151
R976 B.n354 B.n353 10.6151
R977 B.n355 B.n354 10.6151
R978 B.n355 B.n54 10.6151
R979 B.n359 B.n54 10.6151
R980 B.n360 B.n359 10.6151
R981 B.n361 B.n360 10.6151
R982 B.n361 B.n52 10.6151
R983 B.n365 B.n52 10.6151
R984 B.n366 B.n365 10.6151
R985 B.n367 B.n366 10.6151
R986 B.n367 B.n50 10.6151
R987 B.n371 B.n50 10.6151
R988 B.n372 B.n371 10.6151
R989 B.n373 B.n372 10.6151
R990 B.n373 B.n48 10.6151
R991 B.n377 B.n48 10.6151
R992 B.n378 B.n377 10.6151
R993 B.n379 B.n378 10.6151
R994 B.n197 B.n112 10.6151
R995 B.n198 B.n197 10.6151
R996 B.n199 B.n198 10.6151
R997 B.n199 B.n110 10.6151
R998 B.n203 B.n110 10.6151
R999 B.n204 B.n203 10.6151
R1000 B.n205 B.n204 10.6151
R1001 B.n205 B.n108 10.6151
R1002 B.n209 B.n108 10.6151
R1003 B.n210 B.n209 10.6151
R1004 B.n211 B.n210 10.6151
R1005 B.n211 B.n106 10.6151
R1006 B.n215 B.n106 10.6151
R1007 B.n218 B.n217 10.6151
R1008 B.n218 B.n102 10.6151
R1009 B.n222 B.n102 10.6151
R1010 B.n223 B.n222 10.6151
R1011 B.n224 B.n223 10.6151
R1012 B.n224 B.n100 10.6151
R1013 B.n228 B.n100 10.6151
R1014 B.n229 B.n228 10.6151
R1015 B.n230 B.n229 10.6151
R1016 B.n234 B.n233 10.6151
R1017 B.n235 B.n234 10.6151
R1018 B.n235 B.n94 10.6151
R1019 B.n239 B.n94 10.6151
R1020 B.n240 B.n239 10.6151
R1021 B.n241 B.n240 10.6151
R1022 B.n241 B.n92 10.6151
R1023 B.n245 B.n92 10.6151
R1024 B.n246 B.n245 10.6151
R1025 B.n247 B.n246 10.6151
R1026 B.n247 B.n90 10.6151
R1027 B.n251 B.n90 10.6151
R1028 B.n252 B.n251 10.6151
R1029 B.n193 B.n192 10.6151
R1030 B.n192 B.n191 10.6151
R1031 B.n191 B.n114 10.6151
R1032 B.n187 B.n114 10.6151
R1033 B.n187 B.n186 10.6151
R1034 B.n186 B.n185 10.6151
R1035 B.n185 B.n116 10.6151
R1036 B.n181 B.n116 10.6151
R1037 B.n181 B.n180 10.6151
R1038 B.n180 B.n179 10.6151
R1039 B.n179 B.n118 10.6151
R1040 B.n175 B.n118 10.6151
R1041 B.n175 B.n174 10.6151
R1042 B.n174 B.n173 10.6151
R1043 B.n173 B.n120 10.6151
R1044 B.n169 B.n120 10.6151
R1045 B.n169 B.n168 10.6151
R1046 B.n168 B.n167 10.6151
R1047 B.n167 B.n122 10.6151
R1048 B.n163 B.n122 10.6151
R1049 B.n163 B.n162 10.6151
R1050 B.n162 B.n161 10.6151
R1051 B.n161 B.n124 10.6151
R1052 B.n157 B.n124 10.6151
R1053 B.n157 B.n156 10.6151
R1054 B.n156 B.n155 10.6151
R1055 B.n155 B.n126 10.6151
R1056 B.n151 B.n126 10.6151
R1057 B.n151 B.n150 10.6151
R1058 B.n150 B.n149 10.6151
R1059 B.n149 B.n128 10.6151
R1060 B.n145 B.n128 10.6151
R1061 B.n145 B.n144 10.6151
R1062 B.n144 B.n143 10.6151
R1063 B.n143 B.n130 10.6151
R1064 B.n139 B.n130 10.6151
R1065 B.n139 B.n138 10.6151
R1066 B.n138 B.n137 10.6151
R1067 B.n137 B.n132 10.6151
R1068 B.n133 B.n132 10.6151
R1069 B.n133 B.n0 10.6151
R1070 B.n499 B.n1 10.6151
R1071 B.n499 B.n498 10.6151
R1072 B.n498 B.n497 10.6151
R1073 B.n497 B.n4 10.6151
R1074 B.n493 B.n4 10.6151
R1075 B.n493 B.n492 10.6151
R1076 B.n492 B.n491 10.6151
R1077 B.n491 B.n6 10.6151
R1078 B.n487 B.n6 10.6151
R1079 B.n487 B.n486 10.6151
R1080 B.n486 B.n485 10.6151
R1081 B.n485 B.n8 10.6151
R1082 B.n481 B.n8 10.6151
R1083 B.n481 B.n480 10.6151
R1084 B.n480 B.n479 10.6151
R1085 B.n479 B.n10 10.6151
R1086 B.n475 B.n10 10.6151
R1087 B.n475 B.n474 10.6151
R1088 B.n474 B.n473 10.6151
R1089 B.n473 B.n12 10.6151
R1090 B.n469 B.n12 10.6151
R1091 B.n469 B.n468 10.6151
R1092 B.n468 B.n467 10.6151
R1093 B.n467 B.n14 10.6151
R1094 B.n463 B.n14 10.6151
R1095 B.n463 B.n462 10.6151
R1096 B.n462 B.n461 10.6151
R1097 B.n461 B.n16 10.6151
R1098 B.n457 B.n16 10.6151
R1099 B.n457 B.n456 10.6151
R1100 B.n456 B.n455 10.6151
R1101 B.n455 B.n18 10.6151
R1102 B.n451 B.n18 10.6151
R1103 B.n451 B.n450 10.6151
R1104 B.n450 B.n449 10.6151
R1105 B.n449 B.n20 10.6151
R1106 B.n445 B.n20 10.6151
R1107 B.n445 B.n444 10.6151
R1108 B.n444 B.n443 10.6151
R1109 B.n443 B.n22 10.6151
R1110 B.n439 B.n22 10.6151
R1111 B.n419 B.n32 9.36635
R1112 B.n402 B.n401 9.36635
R1113 B.n216 B.n215 9.36635
R1114 B.n233 B.n98 9.36635
R1115 B.n503 B.n0 2.81026
R1116 B.n503 B.n1 2.81026
R1117 B.n416 B.n32 1.24928
R1118 B.n403 B.n402 1.24928
R1119 B.n217 B.n216 1.24928
R1120 B.n230 B.n98 1.24928
C0 VDD1 B 1.21235f
C1 B VN 0.976121f
C2 VDD1 VP 2.46808f
C3 VP VN 5.20186f
C4 VDD1 VTAIL 4.46275f
C5 VTAIL VN 2.96624f
C6 VDD1 VN 0.155572f
C7 B w_n3290_n1504# 6.59161f
C8 w_n3290_n1504# VP 6.7798f
C9 w_n3290_n1504# VTAIL 1.98672f
C10 VDD1 w_n3290_n1504# 1.50447f
C11 w_n3290_n1504# VN 6.35737f
C12 VDD2 B 1.28938f
C13 VDD2 VP 0.460508f
C14 VDD2 VTAIL 4.51307f
C15 VDD1 VDD2 1.46057f
C16 VDD2 VN 2.16518f
C17 VDD2 w_n3290_n1504# 1.593f
C18 B VP 1.68532f
C19 B VTAIL 1.69209f
C20 VTAIL VP 2.98034f
C21 VDD2 VSUBS 1.255716f
C22 VDD1 VSUBS 1.809571f
C23 VTAIL VSUBS 0.498273f
C24 VN VSUBS 5.82023f
C25 VP VSUBS 2.428663f
C26 B VSUBS 3.329546f
C27 w_n3290_n1504# VSUBS 62.8127f
C28 B.n0 VSUBS 0.005049f
C29 B.n1 VSUBS 0.005049f
C30 B.n2 VSUBS 0.007985f
C31 B.n3 VSUBS 0.007985f
C32 B.n4 VSUBS 0.007985f
C33 B.n5 VSUBS 0.007985f
C34 B.n6 VSUBS 0.007985f
C35 B.n7 VSUBS 0.007985f
C36 B.n8 VSUBS 0.007985f
C37 B.n9 VSUBS 0.007985f
C38 B.n10 VSUBS 0.007985f
C39 B.n11 VSUBS 0.007985f
C40 B.n12 VSUBS 0.007985f
C41 B.n13 VSUBS 0.007985f
C42 B.n14 VSUBS 0.007985f
C43 B.n15 VSUBS 0.007985f
C44 B.n16 VSUBS 0.007985f
C45 B.n17 VSUBS 0.007985f
C46 B.n18 VSUBS 0.007985f
C47 B.n19 VSUBS 0.007985f
C48 B.n20 VSUBS 0.007985f
C49 B.n21 VSUBS 0.007985f
C50 B.n22 VSUBS 0.007985f
C51 B.n23 VSUBS 0.020087f
C52 B.n24 VSUBS 0.007985f
C53 B.n25 VSUBS 0.007985f
C54 B.n26 VSUBS 0.007985f
C55 B.n27 VSUBS 0.007985f
C56 B.n28 VSUBS 0.007985f
C57 B.n29 VSUBS 0.007985f
C58 B.t5 VSUBS 0.047693f
C59 B.t4 VSUBS 0.061162f
C60 B.t3 VSUBS 0.294804f
C61 B.n30 VSUBS 0.10703f
C62 B.n31 VSUBS 0.093034f
C63 B.n32 VSUBS 0.0185f
C64 B.n33 VSUBS 0.007985f
C65 B.n34 VSUBS 0.007985f
C66 B.n35 VSUBS 0.007985f
C67 B.n36 VSUBS 0.007985f
C68 B.n37 VSUBS 0.007985f
C69 B.t8 VSUBS 0.047694f
C70 B.t7 VSUBS 0.061163f
C71 B.t6 VSUBS 0.294804f
C72 B.n38 VSUBS 0.10703f
C73 B.n39 VSUBS 0.093034f
C74 B.n40 VSUBS 0.007985f
C75 B.n41 VSUBS 0.007985f
C76 B.n42 VSUBS 0.007985f
C77 B.n43 VSUBS 0.007985f
C78 B.n44 VSUBS 0.007985f
C79 B.n45 VSUBS 0.007985f
C80 B.n46 VSUBS 0.019201f
C81 B.n47 VSUBS 0.007985f
C82 B.n48 VSUBS 0.007985f
C83 B.n49 VSUBS 0.007985f
C84 B.n50 VSUBS 0.007985f
C85 B.n51 VSUBS 0.007985f
C86 B.n52 VSUBS 0.007985f
C87 B.n53 VSUBS 0.007985f
C88 B.n54 VSUBS 0.007985f
C89 B.n55 VSUBS 0.007985f
C90 B.n56 VSUBS 0.007985f
C91 B.n57 VSUBS 0.007985f
C92 B.n58 VSUBS 0.007985f
C93 B.n59 VSUBS 0.007985f
C94 B.n60 VSUBS 0.007985f
C95 B.n61 VSUBS 0.007985f
C96 B.n62 VSUBS 0.007985f
C97 B.n63 VSUBS 0.007985f
C98 B.n64 VSUBS 0.007985f
C99 B.n65 VSUBS 0.007985f
C100 B.n66 VSUBS 0.007985f
C101 B.n67 VSUBS 0.007985f
C102 B.n68 VSUBS 0.007985f
C103 B.n69 VSUBS 0.007985f
C104 B.n70 VSUBS 0.007985f
C105 B.n71 VSUBS 0.007985f
C106 B.n72 VSUBS 0.007985f
C107 B.n73 VSUBS 0.007985f
C108 B.n74 VSUBS 0.007985f
C109 B.n75 VSUBS 0.007985f
C110 B.n76 VSUBS 0.007985f
C111 B.n77 VSUBS 0.007985f
C112 B.n78 VSUBS 0.007985f
C113 B.n79 VSUBS 0.007985f
C114 B.n80 VSUBS 0.007985f
C115 B.n81 VSUBS 0.007985f
C116 B.n82 VSUBS 0.007985f
C117 B.n83 VSUBS 0.007985f
C118 B.n84 VSUBS 0.007985f
C119 B.n85 VSUBS 0.007985f
C120 B.n86 VSUBS 0.007985f
C121 B.n87 VSUBS 0.007985f
C122 B.n88 VSUBS 0.007985f
C123 B.n89 VSUBS 0.020087f
C124 B.n90 VSUBS 0.007985f
C125 B.n91 VSUBS 0.007985f
C126 B.n92 VSUBS 0.007985f
C127 B.n93 VSUBS 0.007985f
C128 B.n94 VSUBS 0.007985f
C129 B.n95 VSUBS 0.007985f
C130 B.t1 VSUBS 0.047694f
C131 B.t2 VSUBS 0.061163f
C132 B.t0 VSUBS 0.294804f
C133 B.n96 VSUBS 0.10703f
C134 B.n97 VSUBS 0.093034f
C135 B.n98 VSUBS 0.0185f
C136 B.n99 VSUBS 0.007985f
C137 B.n100 VSUBS 0.007985f
C138 B.n101 VSUBS 0.007985f
C139 B.n102 VSUBS 0.007985f
C140 B.n103 VSUBS 0.007985f
C141 B.t10 VSUBS 0.047693f
C142 B.t11 VSUBS 0.061162f
C143 B.t9 VSUBS 0.294804f
C144 B.n104 VSUBS 0.10703f
C145 B.n105 VSUBS 0.093034f
C146 B.n106 VSUBS 0.007985f
C147 B.n107 VSUBS 0.007985f
C148 B.n108 VSUBS 0.007985f
C149 B.n109 VSUBS 0.007985f
C150 B.n110 VSUBS 0.007985f
C151 B.n111 VSUBS 0.007985f
C152 B.n112 VSUBS 0.020086f
C153 B.n113 VSUBS 0.007985f
C154 B.n114 VSUBS 0.007985f
C155 B.n115 VSUBS 0.007985f
C156 B.n116 VSUBS 0.007985f
C157 B.n117 VSUBS 0.007985f
C158 B.n118 VSUBS 0.007985f
C159 B.n119 VSUBS 0.007985f
C160 B.n120 VSUBS 0.007985f
C161 B.n121 VSUBS 0.007985f
C162 B.n122 VSUBS 0.007985f
C163 B.n123 VSUBS 0.007985f
C164 B.n124 VSUBS 0.007985f
C165 B.n125 VSUBS 0.007985f
C166 B.n126 VSUBS 0.007985f
C167 B.n127 VSUBS 0.007985f
C168 B.n128 VSUBS 0.007985f
C169 B.n129 VSUBS 0.007985f
C170 B.n130 VSUBS 0.007985f
C171 B.n131 VSUBS 0.007985f
C172 B.n132 VSUBS 0.007985f
C173 B.n133 VSUBS 0.007985f
C174 B.n134 VSUBS 0.007985f
C175 B.n135 VSUBS 0.007985f
C176 B.n136 VSUBS 0.007985f
C177 B.n137 VSUBS 0.007985f
C178 B.n138 VSUBS 0.007985f
C179 B.n139 VSUBS 0.007985f
C180 B.n140 VSUBS 0.007985f
C181 B.n141 VSUBS 0.007985f
C182 B.n142 VSUBS 0.007985f
C183 B.n143 VSUBS 0.007985f
C184 B.n144 VSUBS 0.007985f
C185 B.n145 VSUBS 0.007985f
C186 B.n146 VSUBS 0.007985f
C187 B.n147 VSUBS 0.007985f
C188 B.n148 VSUBS 0.007985f
C189 B.n149 VSUBS 0.007985f
C190 B.n150 VSUBS 0.007985f
C191 B.n151 VSUBS 0.007985f
C192 B.n152 VSUBS 0.007985f
C193 B.n153 VSUBS 0.007985f
C194 B.n154 VSUBS 0.007985f
C195 B.n155 VSUBS 0.007985f
C196 B.n156 VSUBS 0.007985f
C197 B.n157 VSUBS 0.007985f
C198 B.n158 VSUBS 0.007985f
C199 B.n159 VSUBS 0.007985f
C200 B.n160 VSUBS 0.007985f
C201 B.n161 VSUBS 0.007985f
C202 B.n162 VSUBS 0.007985f
C203 B.n163 VSUBS 0.007985f
C204 B.n164 VSUBS 0.007985f
C205 B.n165 VSUBS 0.007985f
C206 B.n166 VSUBS 0.007985f
C207 B.n167 VSUBS 0.007985f
C208 B.n168 VSUBS 0.007985f
C209 B.n169 VSUBS 0.007985f
C210 B.n170 VSUBS 0.007985f
C211 B.n171 VSUBS 0.007985f
C212 B.n172 VSUBS 0.007985f
C213 B.n173 VSUBS 0.007985f
C214 B.n174 VSUBS 0.007985f
C215 B.n175 VSUBS 0.007985f
C216 B.n176 VSUBS 0.007985f
C217 B.n177 VSUBS 0.007985f
C218 B.n178 VSUBS 0.007985f
C219 B.n179 VSUBS 0.007985f
C220 B.n180 VSUBS 0.007985f
C221 B.n181 VSUBS 0.007985f
C222 B.n182 VSUBS 0.007985f
C223 B.n183 VSUBS 0.007985f
C224 B.n184 VSUBS 0.007985f
C225 B.n185 VSUBS 0.007985f
C226 B.n186 VSUBS 0.007985f
C227 B.n187 VSUBS 0.007985f
C228 B.n188 VSUBS 0.007985f
C229 B.n189 VSUBS 0.007985f
C230 B.n190 VSUBS 0.007985f
C231 B.n191 VSUBS 0.007985f
C232 B.n192 VSUBS 0.007985f
C233 B.n193 VSUBS 0.018899f
C234 B.n194 VSUBS 0.018899f
C235 B.n195 VSUBS 0.020087f
C236 B.n196 VSUBS 0.007985f
C237 B.n197 VSUBS 0.007985f
C238 B.n198 VSUBS 0.007985f
C239 B.n199 VSUBS 0.007985f
C240 B.n200 VSUBS 0.007985f
C241 B.n201 VSUBS 0.007985f
C242 B.n202 VSUBS 0.007985f
C243 B.n203 VSUBS 0.007985f
C244 B.n204 VSUBS 0.007985f
C245 B.n205 VSUBS 0.007985f
C246 B.n206 VSUBS 0.007985f
C247 B.n207 VSUBS 0.007985f
C248 B.n208 VSUBS 0.007985f
C249 B.n209 VSUBS 0.007985f
C250 B.n210 VSUBS 0.007985f
C251 B.n211 VSUBS 0.007985f
C252 B.n212 VSUBS 0.007985f
C253 B.n213 VSUBS 0.007985f
C254 B.n214 VSUBS 0.007985f
C255 B.n215 VSUBS 0.007515f
C256 B.n216 VSUBS 0.0185f
C257 B.n217 VSUBS 0.004462f
C258 B.n218 VSUBS 0.007985f
C259 B.n219 VSUBS 0.007985f
C260 B.n220 VSUBS 0.007985f
C261 B.n221 VSUBS 0.007985f
C262 B.n222 VSUBS 0.007985f
C263 B.n223 VSUBS 0.007985f
C264 B.n224 VSUBS 0.007985f
C265 B.n225 VSUBS 0.007985f
C266 B.n226 VSUBS 0.007985f
C267 B.n227 VSUBS 0.007985f
C268 B.n228 VSUBS 0.007985f
C269 B.n229 VSUBS 0.007985f
C270 B.n230 VSUBS 0.004462f
C271 B.n231 VSUBS 0.007985f
C272 B.n232 VSUBS 0.007985f
C273 B.n233 VSUBS 0.007515f
C274 B.n234 VSUBS 0.007985f
C275 B.n235 VSUBS 0.007985f
C276 B.n236 VSUBS 0.007985f
C277 B.n237 VSUBS 0.007985f
C278 B.n238 VSUBS 0.007985f
C279 B.n239 VSUBS 0.007985f
C280 B.n240 VSUBS 0.007985f
C281 B.n241 VSUBS 0.007985f
C282 B.n242 VSUBS 0.007985f
C283 B.n243 VSUBS 0.007985f
C284 B.n244 VSUBS 0.007985f
C285 B.n245 VSUBS 0.007985f
C286 B.n246 VSUBS 0.007985f
C287 B.n247 VSUBS 0.007985f
C288 B.n248 VSUBS 0.007985f
C289 B.n249 VSUBS 0.007985f
C290 B.n250 VSUBS 0.007985f
C291 B.n251 VSUBS 0.007985f
C292 B.n252 VSUBS 0.020086f
C293 B.n253 VSUBS 0.018899f
C294 B.n254 VSUBS 0.018899f
C295 B.n255 VSUBS 0.007985f
C296 B.n256 VSUBS 0.007985f
C297 B.n257 VSUBS 0.007985f
C298 B.n258 VSUBS 0.007985f
C299 B.n259 VSUBS 0.007985f
C300 B.n260 VSUBS 0.007985f
C301 B.n261 VSUBS 0.007985f
C302 B.n262 VSUBS 0.007985f
C303 B.n263 VSUBS 0.007985f
C304 B.n264 VSUBS 0.007985f
C305 B.n265 VSUBS 0.007985f
C306 B.n266 VSUBS 0.007985f
C307 B.n267 VSUBS 0.007985f
C308 B.n268 VSUBS 0.007985f
C309 B.n269 VSUBS 0.007985f
C310 B.n270 VSUBS 0.007985f
C311 B.n271 VSUBS 0.007985f
C312 B.n272 VSUBS 0.007985f
C313 B.n273 VSUBS 0.007985f
C314 B.n274 VSUBS 0.007985f
C315 B.n275 VSUBS 0.007985f
C316 B.n276 VSUBS 0.007985f
C317 B.n277 VSUBS 0.007985f
C318 B.n278 VSUBS 0.007985f
C319 B.n279 VSUBS 0.007985f
C320 B.n280 VSUBS 0.007985f
C321 B.n281 VSUBS 0.007985f
C322 B.n282 VSUBS 0.007985f
C323 B.n283 VSUBS 0.007985f
C324 B.n284 VSUBS 0.007985f
C325 B.n285 VSUBS 0.007985f
C326 B.n286 VSUBS 0.007985f
C327 B.n287 VSUBS 0.007985f
C328 B.n288 VSUBS 0.007985f
C329 B.n289 VSUBS 0.007985f
C330 B.n290 VSUBS 0.007985f
C331 B.n291 VSUBS 0.007985f
C332 B.n292 VSUBS 0.007985f
C333 B.n293 VSUBS 0.007985f
C334 B.n294 VSUBS 0.007985f
C335 B.n295 VSUBS 0.007985f
C336 B.n296 VSUBS 0.007985f
C337 B.n297 VSUBS 0.007985f
C338 B.n298 VSUBS 0.007985f
C339 B.n299 VSUBS 0.007985f
C340 B.n300 VSUBS 0.007985f
C341 B.n301 VSUBS 0.007985f
C342 B.n302 VSUBS 0.007985f
C343 B.n303 VSUBS 0.007985f
C344 B.n304 VSUBS 0.007985f
C345 B.n305 VSUBS 0.007985f
C346 B.n306 VSUBS 0.007985f
C347 B.n307 VSUBS 0.007985f
C348 B.n308 VSUBS 0.007985f
C349 B.n309 VSUBS 0.007985f
C350 B.n310 VSUBS 0.007985f
C351 B.n311 VSUBS 0.007985f
C352 B.n312 VSUBS 0.007985f
C353 B.n313 VSUBS 0.007985f
C354 B.n314 VSUBS 0.007985f
C355 B.n315 VSUBS 0.007985f
C356 B.n316 VSUBS 0.007985f
C357 B.n317 VSUBS 0.007985f
C358 B.n318 VSUBS 0.007985f
C359 B.n319 VSUBS 0.007985f
C360 B.n320 VSUBS 0.007985f
C361 B.n321 VSUBS 0.007985f
C362 B.n322 VSUBS 0.007985f
C363 B.n323 VSUBS 0.007985f
C364 B.n324 VSUBS 0.007985f
C365 B.n325 VSUBS 0.007985f
C366 B.n326 VSUBS 0.007985f
C367 B.n327 VSUBS 0.007985f
C368 B.n328 VSUBS 0.007985f
C369 B.n329 VSUBS 0.007985f
C370 B.n330 VSUBS 0.007985f
C371 B.n331 VSUBS 0.007985f
C372 B.n332 VSUBS 0.007985f
C373 B.n333 VSUBS 0.007985f
C374 B.n334 VSUBS 0.007985f
C375 B.n335 VSUBS 0.007985f
C376 B.n336 VSUBS 0.007985f
C377 B.n337 VSUBS 0.007985f
C378 B.n338 VSUBS 0.007985f
C379 B.n339 VSUBS 0.007985f
C380 B.n340 VSUBS 0.007985f
C381 B.n341 VSUBS 0.007985f
C382 B.n342 VSUBS 0.007985f
C383 B.n343 VSUBS 0.007985f
C384 B.n344 VSUBS 0.007985f
C385 B.n345 VSUBS 0.007985f
C386 B.n346 VSUBS 0.007985f
C387 B.n347 VSUBS 0.007985f
C388 B.n348 VSUBS 0.007985f
C389 B.n349 VSUBS 0.007985f
C390 B.n350 VSUBS 0.007985f
C391 B.n351 VSUBS 0.007985f
C392 B.n352 VSUBS 0.007985f
C393 B.n353 VSUBS 0.007985f
C394 B.n354 VSUBS 0.007985f
C395 B.n355 VSUBS 0.007985f
C396 B.n356 VSUBS 0.007985f
C397 B.n357 VSUBS 0.007985f
C398 B.n358 VSUBS 0.007985f
C399 B.n359 VSUBS 0.007985f
C400 B.n360 VSUBS 0.007985f
C401 B.n361 VSUBS 0.007985f
C402 B.n362 VSUBS 0.007985f
C403 B.n363 VSUBS 0.007985f
C404 B.n364 VSUBS 0.007985f
C405 B.n365 VSUBS 0.007985f
C406 B.n366 VSUBS 0.007985f
C407 B.n367 VSUBS 0.007985f
C408 B.n368 VSUBS 0.007985f
C409 B.n369 VSUBS 0.007985f
C410 B.n370 VSUBS 0.007985f
C411 B.n371 VSUBS 0.007985f
C412 B.n372 VSUBS 0.007985f
C413 B.n373 VSUBS 0.007985f
C414 B.n374 VSUBS 0.007985f
C415 B.n375 VSUBS 0.007985f
C416 B.n376 VSUBS 0.007985f
C417 B.n377 VSUBS 0.007985f
C418 B.n378 VSUBS 0.007985f
C419 B.n379 VSUBS 0.019784f
C420 B.n380 VSUBS 0.018899f
C421 B.n381 VSUBS 0.020087f
C422 B.n382 VSUBS 0.007985f
C423 B.n383 VSUBS 0.007985f
C424 B.n384 VSUBS 0.007985f
C425 B.n385 VSUBS 0.007985f
C426 B.n386 VSUBS 0.007985f
C427 B.n387 VSUBS 0.007985f
C428 B.n388 VSUBS 0.007985f
C429 B.n389 VSUBS 0.007985f
C430 B.n390 VSUBS 0.007985f
C431 B.n391 VSUBS 0.007985f
C432 B.n392 VSUBS 0.007985f
C433 B.n393 VSUBS 0.007985f
C434 B.n394 VSUBS 0.007985f
C435 B.n395 VSUBS 0.007985f
C436 B.n396 VSUBS 0.007985f
C437 B.n397 VSUBS 0.007985f
C438 B.n398 VSUBS 0.007985f
C439 B.n399 VSUBS 0.007985f
C440 B.n400 VSUBS 0.007985f
C441 B.n401 VSUBS 0.007515f
C442 B.n402 VSUBS 0.0185f
C443 B.n403 VSUBS 0.004462f
C444 B.n404 VSUBS 0.007985f
C445 B.n405 VSUBS 0.007985f
C446 B.n406 VSUBS 0.007985f
C447 B.n407 VSUBS 0.007985f
C448 B.n408 VSUBS 0.007985f
C449 B.n409 VSUBS 0.007985f
C450 B.n410 VSUBS 0.007985f
C451 B.n411 VSUBS 0.007985f
C452 B.n412 VSUBS 0.007985f
C453 B.n413 VSUBS 0.007985f
C454 B.n414 VSUBS 0.007985f
C455 B.n415 VSUBS 0.007985f
C456 B.n416 VSUBS 0.004462f
C457 B.n417 VSUBS 0.007985f
C458 B.n418 VSUBS 0.007985f
C459 B.n419 VSUBS 0.007515f
C460 B.n420 VSUBS 0.007985f
C461 B.n421 VSUBS 0.007985f
C462 B.n422 VSUBS 0.007985f
C463 B.n423 VSUBS 0.007985f
C464 B.n424 VSUBS 0.007985f
C465 B.n425 VSUBS 0.007985f
C466 B.n426 VSUBS 0.007985f
C467 B.n427 VSUBS 0.007985f
C468 B.n428 VSUBS 0.007985f
C469 B.n429 VSUBS 0.007985f
C470 B.n430 VSUBS 0.007985f
C471 B.n431 VSUBS 0.007985f
C472 B.n432 VSUBS 0.007985f
C473 B.n433 VSUBS 0.007985f
C474 B.n434 VSUBS 0.007985f
C475 B.n435 VSUBS 0.007985f
C476 B.n436 VSUBS 0.007985f
C477 B.n437 VSUBS 0.007985f
C478 B.n438 VSUBS 0.020086f
C479 B.n439 VSUBS 0.018899f
C480 B.n440 VSUBS 0.018899f
C481 B.n441 VSUBS 0.007985f
C482 B.n442 VSUBS 0.007985f
C483 B.n443 VSUBS 0.007985f
C484 B.n444 VSUBS 0.007985f
C485 B.n445 VSUBS 0.007985f
C486 B.n446 VSUBS 0.007985f
C487 B.n447 VSUBS 0.007985f
C488 B.n448 VSUBS 0.007985f
C489 B.n449 VSUBS 0.007985f
C490 B.n450 VSUBS 0.007985f
C491 B.n451 VSUBS 0.007985f
C492 B.n452 VSUBS 0.007985f
C493 B.n453 VSUBS 0.007985f
C494 B.n454 VSUBS 0.007985f
C495 B.n455 VSUBS 0.007985f
C496 B.n456 VSUBS 0.007985f
C497 B.n457 VSUBS 0.007985f
C498 B.n458 VSUBS 0.007985f
C499 B.n459 VSUBS 0.007985f
C500 B.n460 VSUBS 0.007985f
C501 B.n461 VSUBS 0.007985f
C502 B.n462 VSUBS 0.007985f
C503 B.n463 VSUBS 0.007985f
C504 B.n464 VSUBS 0.007985f
C505 B.n465 VSUBS 0.007985f
C506 B.n466 VSUBS 0.007985f
C507 B.n467 VSUBS 0.007985f
C508 B.n468 VSUBS 0.007985f
C509 B.n469 VSUBS 0.007985f
C510 B.n470 VSUBS 0.007985f
C511 B.n471 VSUBS 0.007985f
C512 B.n472 VSUBS 0.007985f
C513 B.n473 VSUBS 0.007985f
C514 B.n474 VSUBS 0.007985f
C515 B.n475 VSUBS 0.007985f
C516 B.n476 VSUBS 0.007985f
C517 B.n477 VSUBS 0.007985f
C518 B.n478 VSUBS 0.007985f
C519 B.n479 VSUBS 0.007985f
C520 B.n480 VSUBS 0.007985f
C521 B.n481 VSUBS 0.007985f
C522 B.n482 VSUBS 0.007985f
C523 B.n483 VSUBS 0.007985f
C524 B.n484 VSUBS 0.007985f
C525 B.n485 VSUBS 0.007985f
C526 B.n486 VSUBS 0.007985f
C527 B.n487 VSUBS 0.007985f
C528 B.n488 VSUBS 0.007985f
C529 B.n489 VSUBS 0.007985f
C530 B.n490 VSUBS 0.007985f
C531 B.n491 VSUBS 0.007985f
C532 B.n492 VSUBS 0.007985f
C533 B.n493 VSUBS 0.007985f
C534 B.n494 VSUBS 0.007985f
C535 B.n495 VSUBS 0.007985f
C536 B.n496 VSUBS 0.007985f
C537 B.n497 VSUBS 0.007985f
C538 B.n498 VSUBS 0.007985f
C539 B.n499 VSUBS 0.007985f
C540 B.n500 VSUBS 0.007985f
C541 B.n501 VSUBS 0.007985f
C542 B.n502 VSUBS 0.007985f
C543 B.n503 VSUBS 0.018081f
C544 VDD1.t4 VSUBS 0.053269f
C545 VDD1.t2 VSUBS 0.053269f
C546 VDD1.n0 VSUBS 0.259061f
C547 VDD1.t1 VSUBS 0.053269f
C548 VDD1.t0 VSUBS 0.053269f
C549 VDD1.n1 VSUBS 0.258583f
C550 VDD1.t6 VSUBS 0.053269f
C551 VDD1.t5 VSUBS 0.053269f
C552 VDD1.n2 VSUBS 0.258583f
C553 VDD1.n3 VSUBS 2.65186f
C554 VDD1.t3 VSUBS 0.053269f
C555 VDD1.t7 VSUBS 0.053269f
C556 VDD1.n4 VSUBS 0.255084f
C557 VDD1.n5 VSUBS 2.15879f
C558 VP.n0 VSUBS 0.072347f
C559 VP.t2 VSUBS 0.718111f
C560 VP.n1 VSUBS 0.09123f
C561 VP.n2 VSUBS 0.054871f
C562 VP.t1 VSUBS 0.718111f
C563 VP.n3 VSUBS 0.044403f
C564 VP.n4 VSUBS 0.054871f
C565 VP.t7 VSUBS 0.718111f
C566 VP.n5 VSUBS 0.09123f
C567 VP.n6 VSUBS 0.072347f
C568 VP.t6 VSUBS 0.718111f
C569 VP.n7 VSUBS 0.072347f
C570 VP.t0 VSUBS 0.718111f
C571 VP.n8 VSUBS 0.09123f
C572 VP.n9 VSUBS 0.054871f
C573 VP.t4 VSUBS 0.718111f
C574 VP.n10 VSUBS 0.044403f
C575 VP.n11 VSUBS 0.409987f
C576 VP.t5 VSUBS 0.718111f
C577 VP.t3 VSUBS 1.01103f
C578 VP.n12 VSUBS 0.447874f
C579 VP.n13 VSUBS 0.447483f
C580 VP.n14 VSUBS 0.068272f
C581 VP.n15 VSUBS 0.109639f
C582 VP.n16 VSUBS 0.054871f
C583 VP.n17 VSUBS 0.054871f
C584 VP.n18 VSUBS 0.054871f
C585 VP.n19 VSUBS 0.109639f
C586 VP.n20 VSUBS 0.068272f
C587 VP.n21 VSUBS 0.324118f
C588 VP.n22 VSUBS 0.08654f
C589 VP.n23 VSUBS 0.054871f
C590 VP.n24 VSUBS 0.054871f
C591 VP.n25 VSUBS 0.054871f
C592 VP.n26 VSUBS 0.069672f
C593 VP.n27 VSUBS 0.100749f
C594 VP.n28 VSUBS 0.505122f
C595 VP.n29 VSUBS 2.22124f
C596 VP.n30 VSUBS 2.26914f
C597 VP.n31 VSUBS 0.505122f
C598 VP.n32 VSUBS 0.100749f
C599 VP.n33 VSUBS 0.069672f
C600 VP.n34 VSUBS 0.054871f
C601 VP.n35 VSUBS 0.054871f
C602 VP.n36 VSUBS 0.054871f
C603 VP.n37 VSUBS 0.08654f
C604 VP.n38 VSUBS 0.324118f
C605 VP.n39 VSUBS 0.068272f
C606 VP.n40 VSUBS 0.109639f
C607 VP.n41 VSUBS 0.054871f
C608 VP.n42 VSUBS 0.054871f
C609 VP.n43 VSUBS 0.054871f
C610 VP.n44 VSUBS 0.109639f
C611 VP.n45 VSUBS 0.068272f
C612 VP.n46 VSUBS 0.324118f
C613 VP.n47 VSUBS 0.08654f
C614 VP.n48 VSUBS 0.054871f
C615 VP.n49 VSUBS 0.054871f
C616 VP.n50 VSUBS 0.054871f
C617 VP.n51 VSUBS 0.069672f
C618 VP.n52 VSUBS 0.100749f
C619 VP.n53 VSUBS 0.505122f
C620 VP.n54 VSUBS 0.060168f
C621 VTAIL.t14 VSUBS 0.05902f
C622 VTAIL.t12 VSUBS 0.05902f
C623 VTAIL.n0 VSUBS 0.240018f
C624 VTAIL.n1 VSUBS 0.539418f
C625 VTAIL.n2 VSUBS 0.03145f
C626 VTAIL.n3 VSUBS 0.227327f
C627 VTAIL.n4 VSUBS 0.014975f
C628 VTAIL.t15 VSUBS 0.082975f
C629 VTAIL.n5 VSUBS 0.099864f
C630 VTAIL.n6 VSUBS 0.025101f
C631 VTAIL.n7 VSUBS 0.026547f
C632 VTAIL.n8 VSUBS 0.088512f
C633 VTAIL.n9 VSUBS 0.015856f
C634 VTAIL.n10 VSUBS 0.014975f
C635 VTAIL.n11 VSUBS 0.06137f
C636 VTAIL.n12 VSUBS 0.044541f
C637 VTAIL.n13 VSUBS 0.243869f
C638 VTAIL.n14 VSUBS 0.03145f
C639 VTAIL.n15 VSUBS 0.227327f
C640 VTAIL.n16 VSUBS 0.014975f
C641 VTAIL.t4 VSUBS 0.082975f
C642 VTAIL.n17 VSUBS 0.099864f
C643 VTAIL.n18 VSUBS 0.025101f
C644 VTAIL.n19 VSUBS 0.026547f
C645 VTAIL.n20 VSUBS 0.088512f
C646 VTAIL.n21 VSUBS 0.015856f
C647 VTAIL.n22 VSUBS 0.014975f
C648 VTAIL.n23 VSUBS 0.06137f
C649 VTAIL.n24 VSUBS 0.044541f
C650 VTAIL.n25 VSUBS 0.243869f
C651 VTAIL.t2 VSUBS 0.05902f
C652 VTAIL.t3 VSUBS 0.05902f
C653 VTAIL.n26 VSUBS 0.240018f
C654 VTAIL.n27 VSUBS 0.713788f
C655 VTAIL.n28 VSUBS 0.03145f
C656 VTAIL.n29 VSUBS 0.227327f
C657 VTAIL.n30 VSUBS 0.014975f
C658 VTAIL.t7 VSUBS 0.082975f
C659 VTAIL.n31 VSUBS 0.099864f
C660 VTAIL.n32 VSUBS 0.025101f
C661 VTAIL.n33 VSUBS 0.026547f
C662 VTAIL.n34 VSUBS 0.088512f
C663 VTAIL.n35 VSUBS 0.015856f
C664 VTAIL.n36 VSUBS 0.014975f
C665 VTAIL.n37 VSUBS 0.06137f
C666 VTAIL.n38 VSUBS 0.044541f
C667 VTAIL.n39 VSUBS 0.967296f
C668 VTAIL.n40 VSUBS 0.03145f
C669 VTAIL.n41 VSUBS 0.227327f
C670 VTAIL.n42 VSUBS 0.014975f
C671 VTAIL.t8 VSUBS 0.082975f
C672 VTAIL.n43 VSUBS 0.099864f
C673 VTAIL.n44 VSUBS 0.025101f
C674 VTAIL.n45 VSUBS 0.026547f
C675 VTAIL.n46 VSUBS 0.088512f
C676 VTAIL.n47 VSUBS 0.015856f
C677 VTAIL.n48 VSUBS 0.014975f
C678 VTAIL.n49 VSUBS 0.06137f
C679 VTAIL.n50 VSUBS 0.044541f
C680 VTAIL.n51 VSUBS 0.967296f
C681 VTAIL.t10 VSUBS 0.05902f
C682 VTAIL.t11 VSUBS 0.05902f
C683 VTAIL.n52 VSUBS 0.240019f
C684 VTAIL.n53 VSUBS 0.713787f
C685 VTAIL.n54 VSUBS 0.03145f
C686 VTAIL.n55 VSUBS 0.227327f
C687 VTAIL.n56 VSUBS 0.014975f
C688 VTAIL.t13 VSUBS 0.082975f
C689 VTAIL.n57 VSUBS 0.099864f
C690 VTAIL.n58 VSUBS 0.025101f
C691 VTAIL.n59 VSUBS 0.026547f
C692 VTAIL.n60 VSUBS 0.088512f
C693 VTAIL.n61 VSUBS 0.015856f
C694 VTAIL.n62 VSUBS 0.014975f
C695 VTAIL.n63 VSUBS 0.06137f
C696 VTAIL.n64 VSUBS 0.044541f
C697 VTAIL.n65 VSUBS 0.243869f
C698 VTAIL.n66 VSUBS 0.03145f
C699 VTAIL.n67 VSUBS 0.227327f
C700 VTAIL.n68 VSUBS 0.014975f
C701 VTAIL.t1 VSUBS 0.082975f
C702 VTAIL.n69 VSUBS 0.099864f
C703 VTAIL.n70 VSUBS 0.025101f
C704 VTAIL.n71 VSUBS 0.026547f
C705 VTAIL.n72 VSUBS 0.088512f
C706 VTAIL.n73 VSUBS 0.015856f
C707 VTAIL.n74 VSUBS 0.014975f
C708 VTAIL.n75 VSUBS 0.06137f
C709 VTAIL.n76 VSUBS 0.044541f
C710 VTAIL.n77 VSUBS 0.243869f
C711 VTAIL.t6 VSUBS 0.05902f
C712 VTAIL.t0 VSUBS 0.05902f
C713 VTAIL.n78 VSUBS 0.240019f
C714 VTAIL.n79 VSUBS 0.713787f
C715 VTAIL.n80 VSUBS 0.03145f
C716 VTAIL.n81 VSUBS 0.227327f
C717 VTAIL.n82 VSUBS 0.014975f
C718 VTAIL.t5 VSUBS 0.082975f
C719 VTAIL.n83 VSUBS 0.099864f
C720 VTAIL.n84 VSUBS 0.025101f
C721 VTAIL.n85 VSUBS 0.026547f
C722 VTAIL.n86 VSUBS 0.088512f
C723 VTAIL.n87 VSUBS 0.015856f
C724 VTAIL.n88 VSUBS 0.014975f
C725 VTAIL.n89 VSUBS 0.06137f
C726 VTAIL.n90 VSUBS 0.044541f
C727 VTAIL.n91 VSUBS 0.967296f
C728 VTAIL.n92 VSUBS 0.03145f
C729 VTAIL.n93 VSUBS 0.227327f
C730 VTAIL.n94 VSUBS 0.014975f
C731 VTAIL.t9 VSUBS 0.082975f
C732 VTAIL.n95 VSUBS 0.099864f
C733 VTAIL.n96 VSUBS 0.025101f
C734 VTAIL.n97 VSUBS 0.026547f
C735 VTAIL.n98 VSUBS 0.088512f
C736 VTAIL.n99 VSUBS 0.015856f
C737 VTAIL.n100 VSUBS 0.014975f
C738 VTAIL.n101 VSUBS 0.06137f
C739 VTAIL.n102 VSUBS 0.044541f
C740 VTAIL.n103 VSUBS 0.962071f
C741 VDD2.t3 VSUBS 0.051672f
C742 VDD2.t2 VSUBS 0.051672f
C743 VDD2.n0 VSUBS 0.25083f
C744 VDD2.t5 VSUBS 0.051672f
C745 VDD2.t0 VSUBS 0.051672f
C746 VDD2.n1 VSUBS 0.25083f
C747 VDD2.n2 VSUBS 2.52096f
C748 VDD2.t7 VSUBS 0.051672f
C749 VDD2.t6 VSUBS 0.051672f
C750 VDD2.n3 VSUBS 0.247435f
C751 VDD2.n4 VSUBS 2.06448f
C752 VDD2.t4 VSUBS 0.051672f
C753 VDD2.t1 VSUBS 0.051672f
C754 VDD2.n5 VSUBS 0.250816f
C755 VN.n0 VSUBS 0.069148f
C756 VN.t6 VSUBS 0.686361f
C757 VN.n1 VSUBS 0.087197f
C758 VN.n2 VSUBS 0.052445f
C759 VN.t3 VSUBS 0.686361f
C760 VN.n3 VSUBS 0.04244f
C761 VN.n4 VSUBS 0.39186f
C762 VN.t1 VSUBS 0.686361f
C763 VN.t0 VSUBS 0.966331f
C764 VN.n5 VSUBS 0.428073f
C765 VN.n6 VSUBS 0.427698f
C766 VN.n7 VSUBS 0.065253f
C767 VN.n8 VSUBS 0.104792f
C768 VN.n9 VSUBS 0.052445f
C769 VN.n10 VSUBS 0.052445f
C770 VN.n11 VSUBS 0.052445f
C771 VN.n12 VSUBS 0.104792f
C772 VN.n13 VSUBS 0.065253f
C773 VN.n14 VSUBS 0.309788f
C774 VN.n15 VSUBS 0.082714f
C775 VN.n16 VSUBS 0.052445f
C776 VN.n17 VSUBS 0.052445f
C777 VN.n18 VSUBS 0.052445f
C778 VN.n19 VSUBS 0.066592f
C779 VN.n20 VSUBS 0.096295f
C780 VN.n21 VSUBS 0.482789f
C781 VN.n22 VSUBS 0.057508f
C782 VN.n23 VSUBS 0.069148f
C783 VN.t7 VSUBS 0.686361f
C784 VN.n24 VSUBS 0.087197f
C785 VN.n25 VSUBS 0.052445f
C786 VN.t5 VSUBS 0.686361f
C787 VN.n26 VSUBS 0.04244f
C788 VN.n27 VSUBS 0.39186f
C789 VN.t4 VSUBS 0.686361f
C790 VN.t2 VSUBS 0.966331f
C791 VN.n28 VSUBS 0.428073f
C792 VN.n29 VSUBS 0.427698f
C793 VN.n30 VSUBS 0.065253f
C794 VN.n31 VSUBS 0.104792f
C795 VN.n32 VSUBS 0.052445f
C796 VN.n33 VSUBS 0.052445f
C797 VN.n34 VSUBS 0.052445f
C798 VN.n35 VSUBS 0.104792f
C799 VN.n36 VSUBS 0.065253f
C800 VN.n37 VSUBS 0.309788f
C801 VN.n38 VSUBS 0.082714f
C802 VN.n39 VSUBS 0.052445f
C803 VN.n40 VSUBS 0.052445f
C804 VN.n41 VSUBS 0.052445f
C805 VN.n42 VSUBS 0.066592f
C806 VN.n43 VSUBS 0.096295f
C807 VN.n44 VSUBS 0.482789f
C808 VN.n45 VSUBS 2.15218f
.ends

