* NGSPICE file created from diff_pair_sample_0509.ext - technology: sky130A

.subckt diff_pair_sample_0509 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VP.t0 VDD1.t2 B.t7 sky130_fd_pr__nfet_01v8 ad=2.27205 pd=14.1 as=2.27205 ps=14.1 w=13.77 l=1.82
X1 VTAIL.t14 VP.t1 VDD1.t4 B.t0 sky130_fd_pr__nfet_01v8 ad=5.3703 pd=28.32 as=2.27205 ps=14.1 w=13.77 l=1.82
X2 VDD2.t7 VN.t0 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.27205 pd=14.1 as=2.27205 ps=14.1 w=13.77 l=1.82
X3 VDD1.t6 VP.t2 VTAIL.t13 B.t1 sky130_fd_pr__nfet_01v8 ad=2.27205 pd=14.1 as=5.3703 ps=28.32 w=13.77 l=1.82
X4 VDD1.t0 VP.t3 VTAIL.t12 B.t2 sky130_fd_pr__nfet_01v8 ad=2.27205 pd=14.1 as=2.27205 ps=14.1 w=13.77 l=1.82
X5 VTAIL.t5 VN.t1 VDD2.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=5.3703 pd=28.32 as=2.27205 ps=14.1 w=13.77 l=1.82
X6 VDD2.t5 VN.t2 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.27205 pd=14.1 as=5.3703 ps=28.32 w=13.77 l=1.82
X7 B.t21 B.t19 B.t20 B.t9 sky130_fd_pr__nfet_01v8 ad=5.3703 pd=28.32 as=0 ps=0 w=13.77 l=1.82
X8 VTAIL.t7 VN.t3 VDD2.t4 B.t7 sky130_fd_pr__nfet_01v8 ad=2.27205 pd=14.1 as=2.27205 ps=14.1 w=13.77 l=1.82
X9 B.t18 B.t16 B.t17 B.t13 sky130_fd_pr__nfet_01v8 ad=5.3703 pd=28.32 as=0 ps=0 w=13.77 l=1.82
X10 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=5.3703 pd=28.32 as=0 ps=0 w=13.77 l=1.82
X11 VDD2.t3 VN.t4 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.27205 pd=14.1 as=2.27205 ps=14.1 w=13.77 l=1.82
X12 VTAIL.t0 VN.t5 VDD2.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=5.3703 pd=28.32 as=2.27205 ps=14.1 w=13.77 l=1.82
X13 VDD2.t1 VN.t6 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=2.27205 pd=14.1 as=5.3703 ps=28.32 w=13.77 l=1.82
X14 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=5.3703 pd=28.32 as=0 ps=0 w=13.77 l=1.82
X15 VTAIL.t6 VN.t7 VDD2.t0 B.t6 sky130_fd_pr__nfet_01v8 ad=2.27205 pd=14.1 as=2.27205 ps=14.1 w=13.77 l=1.82
X16 VTAIL.t11 VP.t4 VDD1.t7 B.t5 sky130_fd_pr__nfet_01v8 ad=5.3703 pd=28.32 as=2.27205 ps=14.1 w=13.77 l=1.82
X17 VTAIL.t10 VP.t5 VDD1.t1 B.t6 sky130_fd_pr__nfet_01v8 ad=2.27205 pd=14.1 as=2.27205 ps=14.1 w=13.77 l=1.82
X18 VDD1.t3 VP.t6 VTAIL.t9 B.t3 sky130_fd_pr__nfet_01v8 ad=2.27205 pd=14.1 as=2.27205 ps=14.1 w=13.77 l=1.82
X19 VDD1.t5 VP.t7 VTAIL.t8 B.t4 sky130_fd_pr__nfet_01v8 ad=2.27205 pd=14.1 as=5.3703 ps=28.32 w=13.77 l=1.82
R0 VP.n10 VP.t1 213.773
R1 VP.n28 VP.t4 182.339
R2 VP.n35 VP.t6 182.339
R3 VP.n42 VP.t5 182.339
R4 VP.n49 VP.t7 182.339
R5 VP.n25 VP.t2 182.339
R6 VP.n18 VP.t0 182.339
R7 VP.n11 VP.t3 182.339
R8 VP.n13 VP.n12 161.3
R9 VP.n14 VP.n9 161.3
R10 VP.n16 VP.n15 161.3
R11 VP.n17 VP.n8 161.3
R12 VP.n20 VP.n19 161.3
R13 VP.n21 VP.n7 161.3
R14 VP.n23 VP.n22 161.3
R15 VP.n24 VP.n6 161.3
R16 VP.n48 VP.n0 161.3
R17 VP.n47 VP.n46 161.3
R18 VP.n45 VP.n1 161.3
R19 VP.n44 VP.n43 161.3
R20 VP.n41 VP.n2 161.3
R21 VP.n40 VP.n39 161.3
R22 VP.n38 VP.n3 161.3
R23 VP.n37 VP.n36 161.3
R24 VP.n34 VP.n4 161.3
R25 VP.n33 VP.n32 161.3
R26 VP.n31 VP.n5 161.3
R27 VP.n30 VP.n29 161.3
R28 VP.n28 VP.n27 87.5128
R29 VP.n50 VP.n49 87.5128
R30 VP.n26 VP.n25 87.5128
R31 VP.n40 VP.n3 56.5193
R32 VP.n16 VP.n9 56.5193
R33 VP.n11 VP.n10 53.8955
R34 VP.n33 VP.n5 50.2061
R35 VP.n47 VP.n1 50.2061
R36 VP.n23 VP.n7 50.2061
R37 VP.n27 VP.n26 48.6208
R38 VP.n29 VP.n5 30.7807
R39 VP.n48 VP.n47 30.7807
R40 VP.n24 VP.n23 30.7807
R41 VP.n34 VP.n33 24.4675
R42 VP.n36 VP.n3 24.4675
R43 VP.n41 VP.n40 24.4675
R44 VP.n43 VP.n1 24.4675
R45 VP.n17 VP.n16 24.4675
R46 VP.n19 VP.n7 24.4675
R47 VP.n12 VP.n9 24.4675
R48 VP.n29 VP.n28 23.2442
R49 VP.n49 VP.n48 23.2442
R50 VP.n25 VP.n24 23.2442
R51 VP.n36 VP.n35 15.9041
R52 VP.n42 VP.n41 15.9041
R53 VP.n18 VP.n17 15.9041
R54 VP.n12 VP.n11 15.9041
R55 VP.n13 VP.n10 12.7761
R56 VP.n35 VP.n34 8.56395
R57 VP.n43 VP.n42 8.56395
R58 VP.n19 VP.n18 8.56395
R59 VP.n26 VP.n6 0.278367
R60 VP.n30 VP.n27 0.278367
R61 VP.n50 VP.n0 0.278367
R62 VP.n14 VP.n13 0.189894
R63 VP.n15 VP.n14 0.189894
R64 VP.n15 VP.n8 0.189894
R65 VP.n20 VP.n8 0.189894
R66 VP.n21 VP.n20 0.189894
R67 VP.n22 VP.n21 0.189894
R68 VP.n22 VP.n6 0.189894
R69 VP.n31 VP.n30 0.189894
R70 VP.n32 VP.n31 0.189894
R71 VP.n32 VP.n4 0.189894
R72 VP.n37 VP.n4 0.189894
R73 VP.n38 VP.n37 0.189894
R74 VP.n39 VP.n38 0.189894
R75 VP.n39 VP.n2 0.189894
R76 VP.n44 VP.n2 0.189894
R77 VP.n45 VP.n44 0.189894
R78 VP.n46 VP.n45 0.189894
R79 VP.n46 VP.n0 0.189894
R80 VP VP.n50 0.153454
R81 VDD1 VDD1.n0 66.1248
R82 VDD1.n3 VDD1.n2 66.011
R83 VDD1.n3 VDD1.n1 66.011
R84 VDD1.n5 VDD1.n4 65.1397
R85 VDD1.n5 VDD1.n3 44.5095
R86 VDD1.n4 VDD1.t2 1.43841
R87 VDD1.n4 VDD1.t6 1.43841
R88 VDD1.n0 VDD1.t4 1.43841
R89 VDD1.n0 VDD1.t0 1.43841
R90 VDD1.n2 VDD1.t1 1.43841
R91 VDD1.n2 VDD1.t5 1.43841
R92 VDD1.n1 VDD1.t7 1.43841
R93 VDD1.n1 VDD1.t3 1.43841
R94 VDD1 VDD1.n5 0.869035
R95 VTAIL.n11 VTAIL.t14 49.899
R96 VTAIL.n10 VTAIL.t4 49.899
R97 VTAIL.n7 VTAIL.t5 49.899
R98 VTAIL.n15 VTAIL.t1 49.8988
R99 VTAIL.n2 VTAIL.t0 49.8988
R100 VTAIL.n3 VTAIL.t8 49.8988
R101 VTAIL.n6 VTAIL.t11 49.8988
R102 VTAIL.n14 VTAIL.t13 49.8988
R103 VTAIL.n13 VTAIL.n12 48.4611
R104 VTAIL.n9 VTAIL.n8 48.4611
R105 VTAIL.n1 VTAIL.n0 48.4609
R106 VTAIL.n5 VTAIL.n4 48.4609
R107 VTAIL.n15 VTAIL.n14 26.091
R108 VTAIL.n7 VTAIL.n6 26.091
R109 VTAIL.n9 VTAIL.n7 1.85395
R110 VTAIL.n10 VTAIL.n9 1.85395
R111 VTAIL.n13 VTAIL.n11 1.85395
R112 VTAIL.n14 VTAIL.n13 1.85395
R113 VTAIL.n6 VTAIL.n5 1.85395
R114 VTAIL.n5 VTAIL.n3 1.85395
R115 VTAIL.n2 VTAIL.n1 1.85395
R116 VTAIL VTAIL.n15 1.79576
R117 VTAIL.n0 VTAIL.t2 1.43841
R118 VTAIL.n0 VTAIL.t7 1.43841
R119 VTAIL.n4 VTAIL.t9 1.43841
R120 VTAIL.n4 VTAIL.t10 1.43841
R121 VTAIL.n12 VTAIL.t12 1.43841
R122 VTAIL.n12 VTAIL.t15 1.43841
R123 VTAIL.n8 VTAIL.t3 1.43841
R124 VTAIL.n8 VTAIL.t6 1.43841
R125 VTAIL.n11 VTAIL.n10 0.470328
R126 VTAIL.n3 VTAIL.n2 0.470328
R127 VTAIL VTAIL.n1 0.0586897
R128 B.n841 B.n840 585
R129 B.n842 B.n841 585
R130 B.n332 B.n126 585
R131 B.n331 B.n330 585
R132 B.n329 B.n328 585
R133 B.n327 B.n326 585
R134 B.n325 B.n324 585
R135 B.n323 B.n322 585
R136 B.n321 B.n320 585
R137 B.n319 B.n318 585
R138 B.n317 B.n316 585
R139 B.n315 B.n314 585
R140 B.n313 B.n312 585
R141 B.n311 B.n310 585
R142 B.n309 B.n308 585
R143 B.n307 B.n306 585
R144 B.n305 B.n304 585
R145 B.n303 B.n302 585
R146 B.n301 B.n300 585
R147 B.n299 B.n298 585
R148 B.n297 B.n296 585
R149 B.n295 B.n294 585
R150 B.n293 B.n292 585
R151 B.n291 B.n290 585
R152 B.n289 B.n288 585
R153 B.n287 B.n286 585
R154 B.n285 B.n284 585
R155 B.n283 B.n282 585
R156 B.n281 B.n280 585
R157 B.n279 B.n278 585
R158 B.n277 B.n276 585
R159 B.n275 B.n274 585
R160 B.n273 B.n272 585
R161 B.n271 B.n270 585
R162 B.n269 B.n268 585
R163 B.n267 B.n266 585
R164 B.n265 B.n264 585
R165 B.n263 B.n262 585
R166 B.n261 B.n260 585
R167 B.n259 B.n258 585
R168 B.n257 B.n256 585
R169 B.n255 B.n254 585
R170 B.n253 B.n252 585
R171 B.n251 B.n250 585
R172 B.n249 B.n248 585
R173 B.n247 B.n246 585
R174 B.n245 B.n244 585
R175 B.n243 B.n242 585
R176 B.n241 B.n240 585
R177 B.n239 B.n238 585
R178 B.n237 B.n236 585
R179 B.n235 B.n234 585
R180 B.n233 B.n232 585
R181 B.n231 B.n230 585
R182 B.n229 B.n228 585
R183 B.n227 B.n226 585
R184 B.n225 B.n224 585
R185 B.n222 B.n221 585
R186 B.n220 B.n219 585
R187 B.n218 B.n217 585
R188 B.n216 B.n215 585
R189 B.n214 B.n213 585
R190 B.n212 B.n211 585
R191 B.n210 B.n209 585
R192 B.n208 B.n207 585
R193 B.n206 B.n205 585
R194 B.n204 B.n203 585
R195 B.n202 B.n201 585
R196 B.n200 B.n199 585
R197 B.n198 B.n197 585
R198 B.n196 B.n195 585
R199 B.n194 B.n193 585
R200 B.n192 B.n191 585
R201 B.n190 B.n189 585
R202 B.n188 B.n187 585
R203 B.n186 B.n185 585
R204 B.n184 B.n183 585
R205 B.n182 B.n181 585
R206 B.n180 B.n179 585
R207 B.n178 B.n177 585
R208 B.n176 B.n175 585
R209 B.n174 B.n173 585
R210 B.n172 B.n171 585
R211 B.n170 B.n169 585
R212 B.n168 B.n167 585
R213 B.n166 B.n165 585
R214 B.n164 B.n163 585
R215 B.n162 B.n161 585
R216 B.n160 B.n159 585
R217 B.n158 B.n157 585
R218 B.n156 B.n155 585
R219 B.n154 B.n153 585
R220 B.n152 B.n151 585
R221 B.n150 B.n149 585
R222 B.n148 B.n147 585
R223 B.n146 B.n145 585
R224 B.n144 B.n143 585
R225 B.n142 B.n141 585
R226 B.n140 B.n139 585
R227 B.n138 B.n137 585
R228 B.n136 B.n135 585
R229 B.n134 B.n133 585
R230 B.n75 B.n74 585
R231 B.n845 B.n844 585
R232 B.n839 B.n127 585
R233 B.n127 B.n72 585
R234 B.n838 B.n71 585
R235 B.n849 B.n71 585
R236 B.n837 B.n70 585
R237 B.n850 B.n70 585
R238 B.n836 B.n69 585
R239 B.n851 B.n69 585
R240 B.n835 B.n834 585
R241 B.n834 B.n65 585
R242 B.n833 B.n64 585
R243 B.n857 B.n64 585
R244 B.n832 B.n63 585
R245 B.n858 B.n63 585
R246 B.n831 B.n62 585
R247 B.n859 B.n62 585
R248 B.n830 B.n829 585
R249 B.n829 B.n58 585
R250 B.n828 B.n57 585
R251 B.n865 B.n57 585
R252 B.n827 B.n56 585
R253 B.n866 B.n56 585
R254 B.n826 B.n55 585
R255 B.n867 B.n55 585
R256 B.n825 B.n824 585
R257 B.n824 B.n51 585
R258 B.n823 B.n50 585
R259 B.n873 B.n50 585
R260 B.n822 B.n49 585
R261 B.n874 B.n49 585
R262 B.n821 B.n48 585
R263 B.n875 B.n48 585
R264 B.n820 B.n819 585
R265 B.n819 B.n44 585
R266 B.n818 B.n43 585
R267 B.n881 B.n43 585
R268 B.n817 B.n42 585
R269 B.n882 B.n42 585
R270 B.n816 B.n41 585
R271 B.n883 B.n41 585
R272 B.n815 B.n814 585
R273 B.n814 B.n37 585
R274 B.n813 B.n36 585
R275 B.n889 B.n36 585
R276 B.n812 B.n35 585
R277 B.n890 B.n35 585
R278 B.n811 B.n34 585
R279 B.n891 B.n34 585
R280 B.n810 B.n809 585
R281 B.n809 B.n30 585
R282 B.n808 B.n29 585
R283 B.n897 B.n29 585
R284 B.n807 B.n28 585
R285 B.n898 B.n28 585
R286 B.n806 B.n27 585
R287 B.n899 B.n27 585
R288 B.n805 B.n804 585
R289 B.n804 B.n26 585
R290 B.n803 B.n22 585
R291 B.n905 B.n22 585
R292 B.n802 B.n21 585
R293 B.n906 B.n21 585
R294 B.n801 B.n20 585
R295 B.n907 B.n20 585
R296 B.n800 B.n799 585
R297 B.n799 B.n16 585
R298 B.n798 B.n15 585
R299 B.n913 B.n15 585
R300 B.n797 B.n14 585
R301 B.n914 B.n14 585
R302 B.n796 B.n13 585
R303 B.n915 B.n13 585
R304 B.n795 B.n794 585
R305 B.n794 B.n12 585
R306 B.n793 B.n792 585
R307 B.n793 B.n8 585
R308 B.n791 B.n7 585
R309 B.n922 B.n7 585
R310 B.n790 B.n6 585
R311 B.n923 B.n6 585
R312 B.n789 B.n5 585
R313 B.n924 B.n5 585
R314 B.n788 B.n787 585
R315 B.n787 B.n4 585
R316 B.n786 B.n333 585
R317 B.n786 B.n785 585
R318 B.n776 B.n334 585
R319 B.n335 B.n334 585
R320 B.n778 B.n777 585
R321 B.n779 B.n778 585
R322 B.n775 B.n339 585
R323 B.n343 B.n339 585
R324 B.n774 B.n773 585
R325 B.n773 B.n772 585
R326 B.n341 B.n340 585
R327 B.n342 B.n341 585
R328 B.n765 B.n764 585
R329 B.n766 B.n765 585
R330 B.n763 B.n348 585
R331 B.n348 B.n347 585
R332 B.n762 B.n761 585
R333 B.n761 B.n760 585
R334 B.n350 B.n349 585
R335 B.n753 B.n350 585
R336 B.n752 B.n751 585
R337 B.n754 B.n752 585
R338 B.n750 B.n355 585
R339 B.n355 B.n354 585
R340 B.n749 B.n748 585
R341 B.n748 B.n747 585
R342 B.n357 B.n356 585
R343 B.n358 B.n357 585
R344 B.n740 B.n739 585
R345 B.n741 B.n740 585
R346 B.n738 B.n362 585
R347 B.n366 B.n362 585
R348 B.n737 B.n736 585
R349 B.n736 B.n735 585
R350 B.n364 B.n363 585
R351 B.n365 B.n364 585
R352 B.n728 B.n727 585
R353 B.n729 B.n728 585
R354 B.n726 B.n371 585
R355 B.n371 B.n370 585
R356 B.n725 B.n724 585
R357 B.n724 B.n723 585
R358 B.n373 B.n372 585
R359 B.n374 B.n373 585
R360 B.n716 B.n715 585
R361 B.n717 B.n716 585
R362 B.n714 B.n379 585
R363 B.n379 B.n378 585
R364 B.n713 B.n712 585
R365 B.n712 B.n711 585
R366 B.n381 B.n380 585
R367 B.n382 B.n381 585
R368 B.n704 B.n703 585
R369 B.n705 B.n704 585
R370 B.n702 B.n387 585
R371 B.n387 B.n386 585
R372 B.n701 B.n700 585
R373 B.n700 B.n699 585
R374 B.n389 B.n388 585
R375 B.n390 B.n389 585
R376 B.n692 B.n691 585
R377 B.n693 B.n692 585
R378 B.n690 B.n394 585
R379 B.n398 B.n394 585
R380 B.n689 B.n688 585
R381 B.n688 B.n687 585
R382 B.n396 B.n395 585
R383 B.n397 B.n396 585
R384 B.n680 B.n679 585
R385 B.n681 B.n680 585
R386 B.n678 B.n403 585
R387 B.n403 B.n402 585
R388 B.n677 B.n676 585
R389 B.n676 B.n675 585
R390 B.n405 B.n404 585
R391 B.n406 B.n405 585
R392 B.n671 B.n670 585
R393 B.n409 B.n408 585
R394 B.n667 B.n666 585
R395 B.n668 B.n667 585
R396 B.n665 B.n460 585
R397 B.n664 B.n663 585
R398 B.n662 B.n661 585
R399 B.n660 B.n659 585
R400 B.n658 B.n657 585
R401 B.n656 B.n655 585
R402 B.n654 B.n653 585
R403 B.n652 B.n651 585
R404 B.n650 B.n649 585
R405 B.n648 B.n647 585
R406 B.n646 B.n645 585
R407 B.n644 B.n643 585
R408 B.n642 B.n641 585
R409 B.n640 B.n639 585
R410 B.n638 B.n637 585
R411 B.n636 B.n635 585
R412 B.n634 B.n633 585
R413 B.n632 B.n631 585
R414 B.n630 B.n629 585
R415 B.n628 B.n627 585
R416 B.n626 B.n625 585
R417 B.n624 B.n623 585
R418 B.n622 B.n621 585
R419 B.n620 B.n619 585
R420 B.n618 B.n617 585
R421 B.n616 B.n615 585
R422 B.n614 B.n613 585
R423 B.n612 B.n611 585
R424 B.n610 B.n609 585
R425 B.n608 B.n607 585
R426 B.n606 B.n605 585
R427 B.n604 B.n603 585
R428 B.n602 B.n601 585
R429 B.n600 B.n599 585
R430 B.n598 B.n597 585
R431 B.n596 B.n595 585
R432 B.n594 B.n593 585
R433 B.n592 B.n591 585
R434 B.n590 B.n589 585
R435 B.n588 B.n587 585
R436 B.n586 B.n585 585
R437 B.n584 B.n583 585
R438 B.n582 B.n581 585
R439 B.n580 B.n579 585
R440 B.n578 B.n577 585
R441 B.n576 B.n575 585
R442 B.n574 B.n573 585
R443 B.n572 B.n571 585
R444 B.n570 B.n569 585
R445 B.n568 B.n567 585
R446 B.n566 B.n565 585
R447 B.n564 B.n563 585
R448 B.n562 B.n561 585
R449 B.n559 B.n558 585
R450 B.n557 B.n556 585
R451 B.n555 B.n554 585
R452 B.n553 B.n552 585
R453 B.n551 B.n550 585
R454 B.n549 B.n548 585
R455 B.n547 B.n546 585
R456 B.n545 B.n544 585
R457 B.n543 B.n542 585
R458 B.n541 B.n540 585
R459 B.n539 B.n538 585
R460 B.n537 B.n536 585
R461 B.n535 B.n534 585
R462 B.n533 B.n532 585
R463 B.n531 B.n530 585
R464 B.n529 B.n528 585
R465 B.n527 B.n526 585
R466 B.n525 B.n524 585
R467 B.n523 B.n522 585
R468 B.n521 B.n520 585
R469 B.n519 B.n518 585
R470 B.n517 B.n516 585
R471 B.n515 B.n514 585
R472 B.n513 B.n512 585
R473 B.n511 B.n510 585
R474 B.n509 B.n508 585
R475 B.n507 B.n506 585
R476 B.n505 B.n504 585
R477 B.n503 B.n502 585
R478 B.n501 B.n500 585
R479 B.n499 B.n498 585
R480 B.n497 B.n496 585
R481 B.n495 B.n494 585
R482 B.n493 B.n492 585
R483 B.n491 B.n490 585
R484 B.n489 B.n488 585
R485 B.n487 B.n486 585
R486 B.n485 B.n484 585
R487 B.n483 B.n482 585
R488 B.n481 B.n480 585
R489 B.n479 B.n478 585
R490 B.n477 B.n476 585
R491 B.n475 B.n474 585
R492 B.n473 B.n472 585
R493 B.n471 B.n470 585
R494 B.n469 B.n468 585
R495 B.n467 B.n466 585
R496 B.n672 B.n407 585
R497 B.n407 B.n406 585
R498 B.n674 B.n673 585
R499 B.n675 B.n674 585
R500 B.n401 B.n400 585
R501 B.n402 B.n401 585
R502 B.n683 B.n682 585
R503 B.n682 B.n681 585
R504 B.n684 B.n399 585
R505 B.n399 B.n397 585
R506 B.n686 B.n685 585
R507 B.n687 B.n686 585
R508 B.n393 B.n392 585
R509 B.n398 B.n393 585
R510 B.n695 B.n694 585
R511 B.n694 B.n693 585
R512 B.n696 B.n391 585
R513 B.n391 B.n390 585
R514 B.n698 B.n697 585
R515 B.n699 B.n698 585
R516 B.n385 B.n384 585
R517 B.n386 B.n385 585
R518 B.n707 B.n706 585
R519 B.n706 B.n705 585
R520 B.n708 B.n383 585
R521 B.n383 B.n382 585
R522 B.n710 B.n709 585
R523 B.n711 B.n710 585
R524 B.n377 B.n376 585
R525 B.n378 B.n377 585
R526 B.n719 B.n718 585
R527 B.n718 B.n717 585
R528 B.n720 B.n375 585
R529 B.n375 B.n374 585
R530 B.n722 B.n721 585
R531 B.n723 B.n722 585
R532 B.n369 B.n368 585
R533 B.n370 B.n369 585
R534 B.n731 B.n730 585
R535 B.n730 B.n729 585
R536 B.n732 B.n367 585
R537 B.n367 B.n365 585
R538 B.n734 B.n733 585
R539 B.n735 B.n734 585
R540 B.n361 B.n360 585
R541 B.n366 B.n361 585
R542 B.n743 B.n742 585
R543 B.n742 B.n741 585
R544 B.n744 B.n359 585
R545 B.n359 B.n358 585
R546 B.n746 B.n745 585
R547 B.n747 B.n746 585
R548 B.n353 B.n352 585
R549 B.n354 B.n353 585
R550 B.n756 B.n755 585
R551 B.n755 B.n754 585
R552 B.n757 B.n351 585
R553 B.n753 B.n351 585
R554 B.n759 B.n758 585
R555 B.n760 B.n759 585
R556 B.n346 B.n345 585
R557 B.n347 B.n346 585
R558 B.n768 B.n767 585
R559 B.n767 B.n766 585
R560 B.n769 B.n344 585
R561 B.n344 B.n342 585
R562 B.n771 B.n770 585
R563 B.n772 B.n771 585
R564 B.n338 B.n337 585
R565 B.n343 B.n338 585
R566 B.n781 B.n780 585
R567 B.n780 B.n779 585
R568 B.n782 B.n336 585
R569 B.n336 B.n335 585
R570 B.n784 B.n783 585
R571 B.n785 B.n784 585
R572 B.n3 B.n0 585
R573 B.n4 B.n3 585
R574 B.n921 B.n1 585
R575 B.n922 B.n921 585
R576 B.n920 B.n919 585
R577 B.n920 B.n8 585
R578 B.n918 B.n9 585
R579 B.n12 B.n9 585
R580 B.n917 B.n916 585
R581 B.n916 B.n915 585
R582 B.n11 B.n10 585
R583 B.n914 B.n11 585
R584 B.n912 B.n911 585
R585 B.n913 B.n912 585
R586 B.n910 B.n17 585
R587 B.n17 B.n16 585
R588 B.n909 B.n908 585
R589 B.n908 B.n907 585
R590 B.n19 B.n18 585
R591 B.n906 B.n19 585
R592 B.n904 B.n903 585
R593 B.n905 B.n904 585
R594 B.n902 B.n23 585
R595 B.n26 B.n23 585
R596 B.n901 B.n900 585
R597 B.n900 B.n899 585
R598 B.n25 B.n24 585
R599 B.n898 B.n25 585
R600 B.n896 B.n895 585
R601 B.n897 B.n896 585
R602 B.n894 B.n31 585
R603 B.n31 B.n30 585
R604 B.n893 B.n892 585
R605 B.n892 B.n891 585
R606 B.n33 B.n32 585
R607 B.n890 B.n33 585
R608 B.n888 B.n887 585
R609 B.n889 B.n888 585
R610 B.n886 B.n38 585
R611 B.n38 B.n37 585
R612 B.n885 B.n884 585
R613 B.n884 B.n883 585
R614 B.n40 B.n39 585
R615 B.n882 B.n40 585
R616 B.n880 B.n879 585
R617 B.n881 B.n880 585
R618 B.n878 B.n45 585
R619 B.n45 B.n44 585
R620 B.n877 B.n876 585
R621 B.n876 B.n875 585
R622 B.n47 B.n46 585
R623 B.n874 B.n47 585
R624 B.n872 B.n871 585
R625 B.n873 B.n872 585
R626 B.n870 B.n52 585
R627 B.n52 B.n51 585
R628 B.n869 B.n868 585
R629 B.n868 B.n867 585
R630 B.n54 B.n53 585
R631 B.n866 B.n54 585
R632 B.n864 B.n863 585
R633 B.n865 B.n864 585
R634 B.n862 B.n59 585
R635 B.n59 B.n58 585
R636 B.n861 B.n860 585
R637 B.n860 B.n859 585
R638 B.n61 B.n60 585
R639 B.n858 B.n61 585
R640 B.n856 B.n855 585
R641 B.n857 B.n856 585
R642 B.n854 B.n66 585
R643 B.n66 B.n65 585
R644 B.n853 B.n852 585
R645 B.n852 B.n851 585
R646 B.n68 B.n67 585
R647 B.n850 B.n68 585
R648 B.n848 B.n847 585
R649 B.n849 B.n848 585
R650 B.n846 B.n73 585
R651 B.n73 B.n72 585
R652 B.n925 B.n924 585
R653 B.n923 B.n2 585
R654 B.n844 B.n73 554.963
R655 B.n841 B.n127 554.963
R656 B.n466 B.n405 554.963
R657 B.n670 B.n407 554.963
R658 B.n131 B.t8 388.8
R659 B.n128 B.t19 388.8
R660 B.n464 B.t12 388.8
R661 B.n461 B.t16 388.8
R662 B.n842 B.n125 256.663
R663 B.n842 B.n124 256.663
R664 B.n842 B.n123 256.663
R665 B.n842 B.n122 256.663
R666 B.n842 B.n121 256.663
R667 B.n842 B.n120 256.663
R668 B.n842 B.n119 256.663
R669 B.n842 B.n118 256.663
R670 B.n842 B.n117 256.663
R671 B.n842 B.n116 256.663
R672 B.n842 B.n115 256.663
R673 B.n842 B.n114 256.663
R674 B.n842 B.n113 256.663
R675 B.n842 B.n112 256.663
R676 B.n842 B.n111 256.663
R677 B.n842 B.n110 256.663
R678 B.n842 B.n109 256.663
R679 B.n842 B.n108 256.663
R680 B.n842 B.n107 256.663
R681 B.n842 B.n106 256.663
R682 B.n842 B.n105 256.663
R683 B.n842 B.n104 256.663
R684 B.n842 B.n103 256.663
R685 B.n842 B.n102 256.663
R686 B.n842 B.n101 256.663
R687 B.n842 B.n100 256.663
R688 B.n842 B.n99 256.663
R689 B.n842 B.n98 256.663
R690 B.n842 B.n97 256.663
R691 B.n842 B.n96 256.663
R692 B.n842 B.n95 256.663
R693 B.n842 B.n94 256.663
R694 B.n842 B.n93 256.663
R695 B.n842 B.n92 256.663
R696 B.n842 B.n91 256.663
R697 B.n842 B.n90 256.663
R698 B.n842 B.n89 256.663
R699 B.n842 B.n88 256.663
R700 B.n842 B.n87 256.663
R701 B.n842 B.n86 256.663
R702 B.n842 B.n85 256.663
R703 B.n842 B.n84 256.663
R704 B.n842 B.n83 256.663
R705 B.n842 B.n82 256.663
R706 B.n842 B.n81 256.663
R707 B.n842 B.n80 256.663
R708 B.n842 B.n79 256.663
R709 B.n842 B.n78 256.663
R710 B.n842 B.n77 256.663
R711 B.n842 B.n76 256.663
R712 B.n843 B.n842 256.663
R713 B.n669 B.n668 256.663
R714 B.n668 B.n410 256.663
R715 B.n668 B.n411 256.663
R716 B.n668 B.n412 256.663
R717 B.n668 B.n413 256.663
R718 B.n668 B.n414 256.663
R719 B.n668 B.n415 256.663
R720 B.n668 B.n416 256.663
R721 B.n668 B.n417 256.663
R722 B.n668 B.n418 256.663
R723 B.n668 B.n419 256.663
R724 B.n668 B.n420 256.663
R725 B.n668 B.n421 256.663
R726 B.n668 B.n422 256.663
R727 B.n668 B.n423 256.663
R728 B.n668 B.n424 256.663
R729 B.n668 B.n425 256.663
R730 B.n668 B.n426 256.663
R731 B.n668 B.n427 256.663
R732 B.n668 B.n428 256.663
R733 B.n668 B.n429 256.663
R734 B.n668 B.n430 256.663
R735 B.n668 B.n431 256.663
R736 B.n668 B.n432 256.663
R737 B.n668 B.n433 256.663
R738 B.n668 B.n434 256.663
R739 B.n668 B.n435 256.663
R740 B.n668 B.n436 256.663
R741 B.n668 B.n437 256.663
R742 B.n668 B.n438 256.663
R743 B.n668 B.n439 256.663
R744 B.n668 B.n440 256.663
R745 B.n668 B.n441 256.663
R746 B.n668 B.n442 256.663
R747 B.n668 B.n443 256.663
R748 B.n668 B.n444 256.663
R749 B.n668 B.n445 256.663
R750 B.n668 B.n446 256.663
R751 B.n668 B.n447 256.663
R752 B.n668 B.n448 256.663
R753 B.n668 B.n449 256.663
R754 B.n668 B.n450 256.663
R755 B.n668 B.n451 256.663
R756 B.n668 B.n452 256.663
R757 B.n668 B.n453 256.663
R758 B.n668 B.n454 256.663
R759 B.n668 B.n455 256.663
R760 B.n668 B.n456 256.663
R761 B.n668 B.n457 256.663
R762 B.n668 B.n458 256.663
R763 B.n668 B.n459 256.663
R764 B.n927 B.n926 256.663
R765 B.n133 B.n75 163.367
R766 B.n137 B.n136 163.367
R767 B.n141 B.n140 163.367
R768 B.n145 B.n144 163.367
R769 B.n149 B.n148 163.367
R770 B.n153 B.n152 163.367
R771 B.n157 B.n156 163.367
R772 B.n161 B.n160 163.367
R773 B.n165 B.n164 163.367
R774 B.n169 B.n168 163.367
R775 B.n173 B.n172 163.367
R776 B.n177 B.n176 163.367
R777 B.n181 B.n180 163.367
R778 B.n185 B.n184 163.367
R779 B.n189 B.n188 163.367
R780 B.n193 B.n192 163.367
R781 B.n197 B.n196 163.367
R782 B.n201 B.n200 163.367
R783 B.n205 B.n204 163.367
R784 B.n209 B.n208 163.367
R785 B.n213 B.n212 163.367
R786 B.n217 B.n216 163.367
R787 B.n221 B.n220 163.367
R788 B.n226 B.n225 163.367
R789 B.n230 B.n229 163.367
R790 B.n234 B.n233 163.367
R791 B.n238 B.n237 163.367
R792 B.n242 B.n241 163.367
R793 B.n246 B.n245 163.367
R794 B.n250 B.n249 163.367
R795 B.n254 B.n253 163.367
R796 B.n258 B.n257 163.367
R797 B.n262 B.n261 163.367
R798 B.n266 B.n265 163.367
R799 B.n270 B.n269 163.367
R800 B.n274 B.n273 163.367
R801 B.n278 B.n277 163.367
R802 B.n282 B.n281 163.367
R803 B.n286 B.n285 163.367
R804 B.n290 B.n289 163.367
R805 B.n294 B.n293 163.367
R806 B.n298 B.n297 163.367
R807 B.n302 B.n301 163.367
R808 B.n306 B.n305 163.367
R809 B.n310 B.n309 163.367
R810 B.n314 B.n313 163.367
R811 B.n318 B.n317 163.367
R812 B.n322 B.n321 163.367
R813 B.n326 B.n325 163.367
R814 B.n330 B.n329 163.367
R815 B.n841 B.n126 163.367
R816 B.n676 B.n405 163.367
R817 B.n676 B.n403 163.367
R818 B.n680 B.n403 163.367
R819 B.n680 B.n396 163.367
R820 B.n688 B.n396 163.367
R821 B.n688 B.n394 163.367
R822 B.n692 B.n394 163.367
R823 B.n692 B.n389 163.367
R824 B.n700 B.n389 163.367
R825 B.n700 B.n387 163.367
R826 B.n704 B.n387 163.367
R827 B.n704 B.n381 163.367
R828 B.n712 B.n381 163.367
R829 B.n712 B.n379 163.367
R830 B.n716 B.n379 163.367
R831 B.n716 B.n373 163.367
R832 B.n724 B.n373 163.367
R833 B.n724 B.n371 163.367
R834 B.n728 B.n371 163.367
R835 B.n728 B.n364 163.367
R836 B.n736 B.n364 163.367
R837 B.n736 B.n362 163.367
R838 B.n740 B.n362 163.367
R839 B.n740 B.n357 163.367
R840 B.n748 B.n357 163.367
R841 B.n748 B.n355 163.367
R842 B.n752 B.n355 163.367
R843 B.n752 B.n350 163.367
R844 B.n761 B.n350 163.367
R845 B.n761 B.n348 163.367
R846 B.n765 B.n348 163.367
R847 B.n765 B.n341 163.367
R848 B.n773 B.n341 163.367
R849 B.n773 B.n339 163.367
R850 B.n778 B.n339 163.367
R851 B.n778 B.n334 163.367
R852 B.n786 B.n334 163.367
R853 B.n787 B.n786 163.367
R854 B.n787 B.n5 163.367
R855 B.n6 B.n5 163.367
R856 B.n7 B.n6 163.367
R857 B.n793 B.n7 163.367
R858 B.n794 B.n793 163.367
R859 B.n794 B.n13 163.367
R860 B.n14 B.n13 163.367
R861 B.n15 B.n14 163.367
R862 B.n799 B.n15 163.367
R863 B.n799 B.n20 163.367
R864 B.n21 B.n20 163.367
R865 B.n22 B.n21 163.367
R866 B.n804 B.n22 163.367
R867 B.n804 B.n27 163.367
R868 B.n28 B.n27 163.367
R869 B.n29 B.n28 163.367
R870 B.n809 B.n29 163.367
R871 B.n809 B.n34 163.367
R872 B.n35 B.n34 163.367
R873 B.n36 B.n35 163.367
R874 B.n814 B.n36 163.367
R875 B.n814 B.n41 163.367
R876 B.n42 B.n41 163.367
R877 B.n43 B.n42 163.367
R878 B.n819 B.n43 163.367
R879 B.n819 B.n48 163.367
R880 B.n49 B.n48 163.367
R881 B.n50 B.n49 163.367
R882 B.n824 B.n50 163.367
R883 B.n824 B.n55 163.367
R884 B.n56 B.n55 163.367
R885 B.n57 B.n56 163.367
R886 B.n829 B.n57 163.367
R887 B.n829 B.n62 163.367
R888 B.n63 B.n62 163.367
R889 B.n64 B.n63 163.367
R890 B.n834 B.n64 163.367
R891 B.n834 B.n69 163.367
R892 B.n70 B.n69 163.367
R893 B.n71 B.n70 163.367
R894 B.n127 B.n71 163.367
R895 B.n667 B.n409 163.367
R896 B.n667 B.n460 163.367
R897 B.n663 B.n662 163.367
R898 B.n659 B.n658 163.367
R899 B.n655 B.n654 163.367
R900 B.n651 B.n650 163.367
R901 B.n647 B.n646 163.367
R902 B.n643 B.n642 163.367
R903 B.n639 B.n638 163.367
R904 B.n635 B.n634 163.367
R905 B.n631 B.n630 163.367
R906 B.n627 B.n626 163.367
R907 B.n623 B.n622 163.367
R908 B.n619 B.n618 163.367
R909 B.n615 B.n614 163.367
R910 B.n611 B.n610 163.367
R911 B.n607 B.n606 163.367
R912 B.n603 B.n602 163.367
R913 B.n599 B.n598 163.367
R914 B.n595 B.n594 163.367
R915 B.n591 B.n590 163.367
R916 B.n587 B.n586 163.367
R917 B.n583 B.n582 163.367
R918 B.n579 B.n578 163.367
R919 B.n575 B.n574 163.367
R920 B.n571 B.n570 163.367
R921 B.n567 B.n566 163.367
R922 B.n563 B.n562 163.367
R923 B.n558 B.n557 163.367
R924 B.n554 B.n553 163.367
R925 B.n550 B.n549 163.367
R926 B.n546 B.n545 163.367
R927 B.n542 B.n541 163.367
R928 B.n538 B.n537 163.367
R929 B.n534 B.n533 163.367
R930 B.n530 B.n529 163.367
R931 B.n526 B.n525 163.367
R932 B.n522 B.n521 163.367
R933 B.n518 B.n517 163.367
R934 B.n514 B.n513 163.367
R935 B.n510 B.n509 163.367
R936 B.n506 B.n505 163.367
R937 B.n502 B.n501 163.367
R938 B.n498 B.n497 163.367
R939 B.n494 B.n493 163.367
R940 B.n490 B.n489 163.367
R941 B.n486 B.n485 163.367
R942 B.n482 B.n481 163.367
R943 B.n478 B.n477 163.367
R944 B.n474 B.n473 163.367
R945 B.n470 B.n469 163.367
R946 B.n674 B.n407 163.367
R947 B.n674 B.n401 163.367
R948 B.n682 B.n401 163.367
R949 B.n682 B.n399 163.367
R950 B.n686 B.n399 163.367
R951 B.n686 B.n393 163.367
R952 B.n694 B.n393 163.367
R953 B.n694 B.n391 163.367
R954 B.n698 B.n391 163.367
R955 B.n698 B.n385 163.367
R956 B.n706 B.n385 163.367
R957 B.n706 B.n383 163.367
R958 B.n710 B.n383 163.367
R959 B.n710 B.n377 163.367
R960 B.n718 B.n377 163.367
R961 B.n718 B.n375 163.367
R962 B.n722 B.n375 163.367
R963 B.n722 B.n369 163.367
R964 B.n730 B.n369 163.367
R965 B.n730 B.n367 163.367
R966 B.n734 B.n367 163.367
R967 B.n734 B.n361 163.367
R968 B.n742 B.n361 163.367
R969 B.n742 B.n359 163.367
R970 B.n746 B.n359 163.367
R971 B.n746 B.n353 163.367
R972 B.n755 B.n353 163.367
R973 B.n755 B.n351 163.367
R974 B.n759 B.n351 163.367
R975 B.n759 B.n346 163.367
R976 B.n767 B.n346 163.367
R977 B.n767 B.n344 163.367
R978 B.n771 B.n344 163.367
R979 B.n771 B.n338 163.367
R980 B.n780 B.n338 163.367
R981 B.n780 B.n336 163.367
R982 B.n784 B.n336 163.367
R983 B.n784 B.n3 163.367
R984 B.n925 B.n3 163.367
R985 B.n921 B.n2 163.367
R986 B.n921 B.n920 163.367
R987 B.n920 B.n9 163.367
R988 B.n916 B.n9 163.367
R989 B.n916 B.n11 163.367
R990 B.n912 B.n11 163.367
R991 B.n912 B.n17 163.367
R992 B.n908 B.n17 163.367
R993 B.n908 B.n19 163.367
R994 B.n904 B.n19 163.367
R995 B.n904 B.n23 163.367
R996 B.n900 B.n23 163.367
R997 B.n900 B.n25 163.367
R998 B.n896 B.n25 163.367
R999 B.n896 B.n31 163.367
R1000 B.n892 B.n31 163.367
R1001 B.n892 B.n33 163.367
R1002 B.n888 B.n33 163.367
R1003 B.n888 B.n38 163.367
R1004 B.n884 B.n38 163.367
R1005 B.n884 B.n40 163.367
R1006 B.n880 B.n40 163.367
R1007 B.n880 B.n45 163.367
R1008 B.n876 B.n45 163.367
R1009 B.n876 B.n47 163.367
R1010 B.n872 B.n47 163.367
R1011 B.n872 B.n52 163.367
R1012 B.n868 B.n52 163.367
R1013 B.n868 B.n54 163.367
R1014 B.n864 B.n54 163.367
R1015 B.n864 B.n59 163.367
R1016 B.n860 B.n59 163.367
R1017 B.n860 B.n61 163.367
R1018 B.n856 B.n61 163.367
R1019 B.n856 B.n66 163.367
R1020 B.n852 B.n66 163.367
R1021 B.n852 B.n68 163.367
R1022 B.n848 B.n68 163.367
R1023 B.n848 B.n73 163.367
R1024 B.n128 B.t20 112.575
R1025 B.n464 B.t15 112.575
R1026 B.n131 B.t10 112.556
R1027 B.n461 B.t18 112.556
R1028 B.n668 B.n406 80.284
R1029 B.n842 B.n72 80.284
R1030 B.n844 B.n843 71.676
R1031 B.n133 B.n76 71.676
R1032 B.n137 B.n77 71.676
R1033 B.n141 B.n78 71.676
R1034 B.n145 B.n79 71.676
R1035 B.n149 B.n80 71.676
R1036 B.n153 B.n81 71.676
R1037 B.n157 B.n82 71.676
R1038 B.n161 B.n83 71.676
R1039 B.n165 B.n84 71.676
R1040 B.n169 B.n85 71.676
R1041 B.n173 B.n86 71.676
R1042 B.n177 B.n87 71.676
R1043 B.n181 B.n88 71.676
R1044 B.n185 B.n89 71.676
R1045 B.n189 B.n90 71.676
R1046 B.n193 B.n91 71.676
R1047 B.n197 B.n92 71.676
R1048 B.n201 B.n93 71.676
R1049 B.n205 B.n94 71.676
R1050 B.n209 B.n95 71.676
R1051 B.n213 B.n96 71.676
R1052 B.n217 B.n97 71.676
R1053 B.n221 B.n98 71.676
R1054 B.n226 B.n99 71.676
R1055 B.n230 B.n100 71.676
R1056 B.n234 B.n101 71.676
R1057 B.n238 B.n102 71.676
R1058 B.n242 B.n103 71.676
R1059 B.n246 B.n104 71.676
R1060 B.n250 B.n105 71.676
R1061 B.n254 B.n106 71.676
R1062 B.n258 B.n107 71.676
R1063 B.n262 B.n108 71.676
R1064 B.n266 B.n109 71.676
R1065 B.n270 B.n110 71.676
R1066 B.n274 B.n111 71.676
R1067 B.n278 B.n112 71.676
R1068 B.n282 B.n113 71.676
R1069 B.n286 B.n114 71.676
R1070 B.n290 B.n115 71.676
R1071 B.n294 B.n116 71.676
R1072 B.n298 B.n117 71.676
R1073 B.n302 B.n118 71.676
R1074 B.n306 B.n119 71.676
R1075 B.n310 B.n120 71.676
R1076 B.n314 B.n121 71.676
R1077 B.n318 B.n122 71.676
R1078 B.n322 B.n123 71.676
R1079 B.n326 B.n124 71.676
R1080 B.n330 B.n125 71.676
R1081 B.n126 B.n125 71.676
R1082 B.n329 B.n124 71.676
R1083 B.n325 B.n123 71.676
R1084 B.n321 B.n122 71.676
R1085 B.n317 B.n121 71.676
R1086 B.n313 B.n120 71.676
R1087 B.n309 B.n119 71.676
R1088 B.n305 B.n118 71.676
R1089 B.n301 B.n117 71.676
R1090 B.n297 B.n116 71.676
R1091 B.n293 B.n115 71.676
R1092 B.n289 B.n114 71.676
R1093 B.n285 B.n113 71.676
R1094 B.n281 B.n112 71.676
R1095 B.n277 B.n111 71.676
R1096 B.n273 B.n110 71.676
R1097 B.n269 B.n109 71.676
R1098 B.n265 B.n108 71.676
R1099 B.n261 B.n107 71.676
R1100 B.n257 B.n106 71.676
R1101 B.n253 B.n105 71.676
R1102 B.n249 B.n104 71.676
R1103 B.n245 B.n103 71.676
R1104 B.n241 B.n102 71.676
R1105 B.n237 B.n101 71.676
R1106 B.n233 B.n100 71.676
R1107 B.n229 B.n99 71.676
R1108 B.n225 B.n98 71.676
R1109 B.n220 B.n97 71.676
R1110 B.n216 B.n96 71.676
R1111 B.n212 B.n95 71.676
R1112 B.n208 B.n94 71.676
R1113 B.n204 B.n93 71.676
R1114 B.n200 B.n92 71.676
R1115 B.n196 B.n91 71.676
R1116 B.n192 B.n90 71.676
R1117 B.n188 B.n89 71.676
R1118 B.n184 B.n88 71.676
R1119 B.n180 B.n87 71.676
R1120 B.n176 B.n86 71.676
R1121 B.n172 B.n85 71.676
R1122 B.n168 B.n84 71.676
R1123 B.n164 B.n83 71.676
R1124 B.n160 B.n82 71.676
R1125 B.n156 B.n81 71.676
R1126 B.n152 B.n80 71.676
R1127 B.n148 B.n79 71.676
R1128 B.n144 B.n78 71.676
R1129 B.n140 B.n77 71.676
R1130 B.n136 B.n76 71.676
R1131 B.n843 B.n75 71.676
R1132 B.n670 B.n669 71.676
R1133 B.n460 B.n410 71.676
R1134 B.n662 B.n411 71.676
R1135 B.n658 B.n412 71.676
R1136 B.n654 B.n413 71.676
R1137 B.n650 B.n414 71.676
R1138 B.n646 B.n415 71.676
R1139 B.n642 B.n416 71.676
R1140 B.n638 B.n417 71.676
R1141 B.n634 B.n418 71.676
R1142 B.n630 B.n419 71.676
R1143 B.n626 B.n420 71.676
R1144 B.n622 B.n421 71.676
R1145 B.n618 B.n422 71.676
R1146 B.n614 B.n423 71.676
R1147 B.n610 B.n424 71.676
R1148 B.n606 B.n425 71.676
R1149 B.n602 B.n426 71.676
R1150 B.n598 B.n427 71.676
R1151 B.n594 B.n428 71.676
R1152 B.n590 B.n429 71.676
R1153 B.n586 B.n430 71.676
R1154 B.n582 B.n431 71.676
R1155 B.n578 B.n432 71.676
R1156 B.n574 B.n433 71.676
R1157 B.n570 B.n434 71.676
R1158 B.n566 B.n435 71.676
R1159 B.n562 B.n436 71.676
R1160 B.n557 B.n437 71.676
R1161 B.n553 B.n438 71.676
R1162 B.n549 B.n439 71.676
R1163 B.n545 B.n440 71.676
R1164 B.n541 B.n441 71.676
R1165 B.n537 B.n442 71.676
R1166 B.n533 B.n443 71.676
R1167 B.n529 B.n444 71.676
R1168 B.n525 B.n445 71.676
R1169 B.n521 B.n446 71.676
R1170 B.n517 B.n447 71.676
R1171 B.n513 B.n448 71.676
R1172 B.n509 B.n449 71.676
R1173 B.n505 B.n450 71.676
R1174 B.n501 B.n451 71.676
R1175 B.n497 B.n452 71.676
R1176 B.n493 B.n453 71.676
R1177 B.n489 B.n454 71.676
R1178 B.n485 B.n455 71.676
R1179 B.n481 B.n456 71.676
R1180 B.n477 B.n457 71.676
R1181 B.n473 B.n458 71.676
R1182 B.n469 B.n459 71.676
R1183 B.n669 B.n409 71.676
R1184 B.n663 B.n410 71.676
R1185 B.n659 B.n411 71.676
R1186 B.n655 B.n412 71.676
R1187 B.n651 B.n413 71.676
R1188 B.n647 B.n414 71.676
R1189 B.n643 B.n415 71.676
R1190 B.n639 B.n416 71.676
R1191 B.n635 B.n417 71.676
R1192 B.n631 B.n418 71.676
R1193 B.n627 B.n419 71.676
R1194 B.n623 B.n420 71.676
R1195 B.n619 B.n421 71.676
R1196 B.n615 B.n422 71.676
R1197 B.n611 B.n423 71.676
R1198 B.n607 B.n424 71.676
R1199 B.n603 B.n425 71.676
R1200 B.n599 B.n426 71.676
R1201 B.n595 B.n427 71.676
R1202 B.n591 B.n428 71.676
R1203 B.n587 B.n429 71.676
R1204 B.n583 B.n430 71.676
R1205 B.n579 B.n431 71.676
R1206 B.n575 B.n432 71.676
R1207 B.n571 B.n433 71.676
R1208 B.n567 B.n434 71.676
R1209 B.n563 B.n435 71.676
R1210 B.n558 B.n436 71.676
R1211 B.n554 B.n437 71.676
R1212 B.n550 B.n438 71.676
R1213 B.n546 B.n439 71.676
R1214 B.n542 B.n440 71.676
R1215 B.n538 B.n441 71.676
R1216 B.n534 B.n442 71.676
R1217 B.n530 B.n443 71.676
R1218 B.n526 B.n444 71.676
R1219 B.n522 B.n445 71.676
R1220 B.n518 B.n446 71.676
R1221 B.n514 B.n447 71.676
R1222 B.n510 B.n448 71.676
R1223 B.n506 B.n449 71.676
R1224 B.n502 B.n450 71.676
R1225 B.n498 B.n451 71.676
R1226 B.n494 B.n452 71.676
R1227 B.n490 B.n453 71.676
R1228 B.n486 B.n454 71.676
R1229 B.n482 B.n455 71.676
R1230 B.n478 B.n456 71.676
R1231 B.n474 B.n457 71.676
R1232 B.n470 B.n458 71.676
R1233 B.n466 B.n459 71.676
R1234 B.n926 B.n925 71.676
R1235 B.n926 B.n2 71.676
R1236 B.n129 B.t21 70.8773
R1237 B.n465 B.t14 70.8773
R1238 B.n132 B.t11 70.8595
R1239 B.n462 B.t17 70.8595
R1240 B.n223 B.n132 59.5399
R1241 B.n130 B.n129 59.5399
R1242 B.n560 B.n465 59.5399
R1243 B.n463 B.n462 59.5399
R1244 B.n132 B.n131 41.6975
R1245 B.n129 B.n128 41.6975
R1246 B.n465 B.n464 41.6975
R1247 B.n462 B.n461 41.6975
R1248 B.n675 B.n406 39.2759
R1249 B.n675 B.n402 39.2759
R1250 B.n681 B.n402 39.2759
R1251 B.n681 B.n397 39.2759
R1252 B.n687 B.n397 39.2759
R1253 B.n687 B.n398 39.2759
R1254 B.n693 B.n390 39.2759
R1255 B.n699 B.n390 39.2759
R1256 B.n699 B.n386 39.2759
R1257 B.n705 B.n386 39.2759
R1258 B.n705 B.n382 39.2759
R1259 B.n711 B.n382 39.2759
R1260 B.n711 B.n378 39.2759
R1261 B.n717 B.n378 39.2759
R1262 B.n723 B.n374 39.2759
R1263 B.n723 B.n370 39.2759
R1264 B.n729 B.n370 39.2759
R1265 B.n729 B.n365 39.2759
R1266 B.n735 B.n365 39.2759
R1267 B.n735 B.n366 39.2759
R1268 B.n741 B.n358 39.2759
R1269 B.n747 B.n358 39.2759
R1270 B.n747 B.n354 39.2759
R1271 B.n754 B.n354 39.2759
R1272 B.n754 B.n753 39.2759
R1273 B.n760 B.n347 39.2759
R1274 B.n766 B.n347 39.2759
R1275 B.n766 B.n342 39.2759
R1276 B.n772 B.n342 39.2759
R1277 B.n772 B.n343 39.2759
R1278 B.n779 B.n335 39.2759
R1279 B.n785 B.n335 39.2759
R1280 B.n785 B.n4 39.2759
R1281 B.n924 B.n4 39.2759
R1282 B.n924 B.n923 39.2759
R1283 B.n923 B.n922 39.2759
R1284 B.n922 B.n8 39.2759
R1285 B.n12 B.n8 39.2759
R1286 B.n915 B.n12 39.2759
R1287 B.n914 B.n913 39.2759
R1288 B.n913 B.n16 39.2759
R1289 B.n907 B.n16 39.2759
R1290 B.n907 B.n906 39.2759
R1291 B.n906 B.n905 39.2759
R1292 B.n899 B.n26 39.2759
R1293 B.n899 B.n898 39.2759
R1294 B.n898 B.n897 39.2759
R1295 B.n897 B.n30 39.2759
R1296 B.n891 B.n30 39.2759
R1297 B.n890 B.n889 39.2759
R1298 B.n889 B.n37 39.2759
R1299 B.n883 B.n37 39.2759
R1300 B.n883 B.n882 39.2759
R1301 B.n882 B.n881 39.2759
R1302 B.n881 B.n44 39.2759
R1303 B.n875 B.n874 39.2759
R1304 B.n874 B.n873 39.2759
R1305 B.n873 B.n51 39.2759
R1306 B.n867 B.n51 39.2759
R1307 B.n867 B.n866 39.2759
R1308 B.n866 B.n865 39.2759
R1309 B.n865 B.n58 39.2759
R1310 B.n859 B.n58 39.2759
R1311 B.n858 B.n857 39.2759
R1312 B.n857 B.n65 39.2759
R1313 B.n851 B.n65 39.2759
R1314 B.n851 B.n850 39.2759
R1315 B.n850 B.n849 39.2759
R1316 B.n849 B.n72 39.2759
R1317 B.n840 B.n839 36.059
R1318 B.n672 B.n671 36.059
R1319 B.n467 B.n404 36.059
R1320 B.n846 B.n845 36.059
R1321 B.n741 B.t3 35.8104
R1322 B.n891 B.t7 35.8104
R1323 B.n693 B.t13 30.0346
R1324 B.n717 B.t5 30.0346
R1325 B.n875 B.t1 30.0346
R1326 B.n859 B.t9 30.0346
R1327 B.n343 B.t4 28.8795
R1328 B.t0 B.n914 28.8795
R1329 B.n760 B.t6 23.1037
R1330 B.n905 B.t2 23.1037
R1331 B B.n927 18.0485
R1332 B.n753 B.t6 16.1727
R1333 B.n26 B.t2 16.1727
R1334 B.n673 B.n672 10.6151
R1335 B.n673 B.n400 10.6151
R1336 B.n683 B.n400 10.6151
R1337 B.n684 B.n683 10.6151
R1338 B.n685 B.n684 10.6151
R1339 B.n685 B.n392 10.6151
R1340 B.n695 B.n392 10.6151
R1341 B.n696 B.n695 10.6151
R1342 B.n697 B.n696 10.6151
R1343 B.n697 B.n384 10.6151
R1344 B.n707 B.n384 10.6151
R1345 B.n708 B.n707 10.6151
R1346 B.n709 B.n708 10.6151
R1347 B.n709 B.n376 10.6151
R1348 B.n719 B.n376 10.6151
R1349 B.n720 B.n719 10.6151
R1350 B.n721 B.n720 10.6151
R1351 B.n721 B.n368 10.6151
R1352 B.n731 B.n368 10.6151
R1353 B.n732 B.n731 10.6151
R1354 B.n733 B.n732 10.6151
R1355 B.n733 B.n360 10.6151
R1356 B.n743 B.n360 10.6151
R1357 B.n744 B.n743 10.6151
R1358 B.n745 B.n744 10.6151
R1359 B.n745 B.n352 10.6151
R1360 B.n756 B.n352 10.6151
R1361 B.n757 B.n756 10.6151
R1362 B.n758 B.n757 10.6151
R1363 B.n758 B.n345 10.6151
R1364 B.n768 B.n345 10.6151
R1365 B.n769 B.n768 10.6151
R1366 B.n770 B.n769 10.6151
R1367 B.n770 B.n337 10.6151
R1368 B.n781 B.n337 10.6151
R1369 B.n782 B.n781 10.6151
R1370 B.n783 B.n782 10.6151
R1371 B.n783 B.n0 10.6151
R1372 B.n671 B.n408 10.6151
R1373 B.n666 B.n408 10.6151
R1374 B.n666 B.n665 10.6151
R1375 B.n665 B.n664 10.6151
R1376 B.n664 B.n661 10.6151
R1377 B.n661 B.n660 10.6151
R1378 B.n660 B.n657 10.6151
R1379 B.n657 B.n656 10.6151
R1380 B.n656 B.n653 10.6151
R1381 B.n653 B.n652 10.6151
R1382 B.n652 B.n649 10.6151
R1383 B.n649 B.n648 10.6151
R1384 B.n648 B.n645 10.6151
R1385 B.n645 B.n644 10.6151
R1386 B.n644 B.n641 10.6151
R1387 B.n641 B.n640 10.6151
R1388 B.n640 B.n637 10.6151
R1389 B.n637 B.n636 10.6151
R1390 B.n636 B.n633 10.6151
R1391 B.n633 B.n632 10.6151
R1392 B.n632 B.n629 10.6151
R1393 B.n629 B.n628 10.6151
R1394 B.n628 B.n625 10.6151
R1395 B.n625 B.n624 10.6151
R1396 B.n624 B.n621 10.6151
R1397 B.n621 B.n620 10.6151
R1398 B.n620 B.n617 10.6151
R1399 B.n617 B.n616 10.6151
R1400 B.n616 B.n613 10.6151
R1401 B.n613 B.n612 10.6151
R1402 B.n612 B.n609 10.6151
R1403 B.n609 B.n608 10.6151
R1404 B.n608 B.n605 10.6151
R1405 B.n605 B.n604 10.6151
R1406 B.n604 B.n601 10.6151
R1407 B.n601 B.n600 10.6151
R1408 B.n600 B.n597 10.6151
R1409 B.n597 B.n596 10.6151
R1410 B.n596 B.n593 10.6151
R1411 B.n593 B.n592 10.6151
R1412 B.n592 B.n589 10.6151
R1413 B.n589 B.n588 10.6151
R1414 B.n588 B.n585 10.6151
R1415 B.n585 B.n584 10.6151
R1416 B.n584 B.n581 10.6151
R1417 B.n581 B.n580 10.6151
R1418 B.n577 B.n576 10.6151
R1419 B.n576 B.n573 10.6151
R1420 B.n573 B.n572 10.6151
R1421 B.n572 B.n569 10.6151
R1422 B.n569 B.n568 10.6151
R1423 B.n568 B.n565 10.6151
R1424 B.n565 B.n564 10.6151
R1425 B.n564 B.n561 10.6151
R1426 B.n559 B.n556 10.6151
R1427 B.n556 B.n555 10.6151
R1428 B.n555 B.n552 10.6151
R1429 B.n552 B.n551 10.6151
R1430 B.n551 B.n548 10.6151
R1431 B.n548 B.n547 10.6151
R1432 B.n547 B.n544 10.6151
R1433 B.n544 B.n543 10.6151
R1434 B.n543 B.n540 10.6151
R1435 B.n540 B.n539 10.6151
R1436 B.n539 B.n536 10.6151
R1437 B.n536 B.n535 10.6151
R1438 B.n535 B.n532 10.6151
R1439 B.n532 B.n531 10.6151
R1440 B.n531 B.n528 10.6151
R1441 B.n528 B.n527 10.6151
R1442 B.n527 B.n524 10.6151
R1443 B.n524 B.n523 10.6151
R1444 B.n523 B.n520 10.6151
R1445 B.n520 B.n519 10.6151
R1446 B.n519 B.n516 10.6151
R1447 B.n516 B.n515 10.6151
R1448 B.n515 B.n512 10.6151
R1449 B.n512 B.n511 10.6151
R1450 B.n511 B.n508 10.6151
R1451 B.n508 B.n507 10.6151
R1452 B.n507 B.n504 10.6151
R1453 B.n504 B.n503 10.6151
R1454 B.n503 B.n500 10.6151
R1455 B.n500 B.n499 10.6151
R1456 B.n499 B.n496 10.6151
R1457 B.n496 B.n495 10.6151
R1458 B.n495 B.n492 10.6151
R1459 B.n492 B.n491 10.6151
R1460 B.n491 B.n488 10.6151
R1461 B.n488 B.n487 10.6151
R1462 B.n487 B.n484 10.6151
R1463 B.n484 B.n483 10.6151
R1464 B.n483 B.n480 10.6151
R1465 B.n480 B.n479 10.6151
R1466 B.n479 B.n476 10.6151
R1467 B.n476 B.n475 10.6151
R1468 B.n475 B.n472 10.6151
R1469 B.n472 B.n471 10.6151
R1470 B.n471 B.n468 10.6151
R1471 B.n468 B.n467 10.6151
R1472 B.n677 B.n404 10.6151
R1473 B.n678 B.n677 10.6151
R1474 B.n679 B.n678 10.6151
R1475 B.n679 B.n395 10.6151
R1476 B.n689 B.n395 10.6151
R1477 B.n690 B.n689 10.6151
R1478 B.n691 B.n690 10.6151
R1479 B.n691 B.n388 10.6151
R1480 B.n701 B.n388 10.6151
R1481 B.n702 B.n701 10.6151
R1482 B.n703 B.n702 10.6151
R1483 B.n703 B.n380 10.6151
R1484 B.n713 B.n380 10.6151
R1485 B.n714 B.n713 10.6151
R1486 B.n715 B.n714 10.6151
R1487 B.n715 B.n372 10.6151
R1488 B.n725 B.n372 10.6151
R1489 B.n726 B.n725 10.6151
R1490 B.n727 B.n726 10.6151
R1491 B.n727 B.n363 10.6151
R1492 B.n737 B.n363 10.6151
R1493 B.n738 B.n737 10.6151
R1494 B.n739 B.n738 10.6151
R1495 B.n739 B.n356 10.6151
R1496 B.n749 B.n356 10.6151
R1497 B.n750 B.n749 10.6151
R1498 B.n751 B.n750 10.6151
R1499 B.n751 B.n349 10.6151
R1500 B.n762 B.n349 10.6151
R1501 B.n763 B.n762 10.6151
R1502 B.n764 B.n763 10.6151
R1503 B.n764 B.n340 10.6151
R1504 B.n774 B.n340 10.6151
R1505 B.n775 B.n774 10.6151
R1506 B.n777 B.n775 10.6151
R1507 B.n777 B.n776 10.6151
R1508 B.n776 B.n333 10.6151
R1509 B.n788 B.n333 10.6151
R1510 B.n789 B.n788 10.6151
R1511 B.n790 B.n789 10.6151
R1512 B.n791 B.n790 10.6151
R1513 B.n792 B.n791 10.6151
R1514 B.n795 B.n792 10.6151
R1515 B.n796 B.n795 10.6151
R1516 B.n797 B.n796 10.6151
R1517 B.n798 B.n797 10.6151
R1518 B.n800 B.n798 10.6151
R1519 B.n801 B.n800 10.6151
R1520 B.n802 B.n801 10.6151
R1521 B.n803 B.n802 10.6151
R1522 B.n805 B.n803 10.6151
R1523 B.n806 B.n805 10.6151
R1524 B.n807 B.n806 10.6151
R1525 B.n808 B.n807 10.6151
R1526 B.n810 B.n808 10.6151
R1527 B.n811 B.n810 10.6151
R1528 B.n812 B.n811 10.6151
R1529 B.n813 B.n812 10.6151
R1530 B.n815 B.n813 10.6151
R1531 B.n816 B.n815 10.6151
R1532 B.n817 B.n816 10.6151
R1533 B.n818 B.n817 10.6151
R1534 B.n820 B.n818 10.6151
R1535 B.n821 B.n820 10.6151
R1536 B.n822 B.n821 10.6151
R1537 B.n823 B.n822 10.6151
R1538 B.n825 B.n823 10.6151
R1539 B.n826 B.n825 10.6151
R1540 B.n827 B.n826 10.6151
R1541 B.n828 B.n827 10.6151
R1542 B.n830 B.n828 10.6151
R1543 B.n831 B.n830 10.6151
R1544 B.n832 B.n831 10.6151
R1545 B.n833 B.n832 10.6151
R1546 B.n835 B.n833 10.6151
R1547 B.n836 B.n835 10.6151
R1548 B.n837 B.n836 10.6151
R1549 B.n838 B.n837 10.6151
R1550 B.n839 B.n838 10.6151
R1551 B.n919 B.n1 10.6151
R1552 B.n919 B.n918 10.6151
R1553 B.n918 B.n917 10.6151
R1554 B.n917 B.n10 10.6151
R1555 B.n911 B.n10 10.6151
R1556 B.n911 B.n910 10.6151
R1557 B.n910 B.n909 10.6151
R1558 B.n909 B.n18 10.6151
R1559 B.n903 B.n18 10.6151
R1560 B.n903 B.n902 10.6151
R1561 B.n902 B.n901 10.6151
R1562 B.n901 B.n24 10.6151
R1563 B.n895 B.n24 10.6151
R1564 B.n895 B.n894 10.6151
R1565 B.n894 B.n893 10.6151
R1566 B.n893 B.n32 10.6151
R1567 B.n887 B.n32 10.6151
R1568 B.n887 B.n886 10.6151
R1569 B.n886 B.n885 10.6151
R1570 B.n885 B.n39 10.6151
R1571 B.n879 B.n39 10.6151
R1572 B.n879 B.n878 10.6151
R1573 B.n878 B.n877 10.6151
R1574 B.n877 B.n46 10.6151
R1575 B.n871 B.n46 10.6151
R1576 B.n871 B.n870 10.6151
R1577 B.n870 B.n869 10.6151
R1578 B.n869 B.n53 10.6151
R1579 B.n863 B.n53 10.6151
R1580 B.n863 B.n862 10.6151
R1581 B.n862 B.n861 10.6151
R1582 B.n861 B.n60 10.6151
R1583 B.n855 B.n60 10.6151
R1584 B.n855 B.n854 10.6151
R1585 B.n854 B.n853 10.6151
R1586 B.n853 B.n67 10.6151
R1587 B.n847 B.n67 10.6151
R1588 B.n847 B.n846 10.6151
R1589 B.n845 B.n74 10.6151
R1590 B.n134 B.n74 10.6151
R1591 B.n135 B.n134 10.6151
R1592 B.n138 B.n135 10.6151
R1593 B.n139 B.n138 10.6151
R1594 B.n142 B.n139 10.6151
R1595 B.n143 B.n142 10.6151
R1596 B.n146 B.n143 10.6151
R1597 B.n147 B.n146 10.6151
R1598 B.n150 B.n147 10.6151
R1599 B.n151 B.n150 10.6151
R1600 B.n154 B.n151 10.6151
R1601 B.n155 B.n154 10.6151
R1602 B.n158 B.n155 10.6151
R1603 B.n159 B.n158 10.6151
R1604 B.n162 B.n159 10.6151
R1605 B.n163 B.n162 10.6151
R1606 B.n166 B.n163 10.6151
R1607 B.n167 B.n166 10.6151
R1608 B.n170 B.n167 10.6151
R1609 B.n171 B.n170 10.6151
R1610 B.n174 B.n171 10.6151
R1611 B.n175 B.n174 10.6151
R1612 B.n178 B.n175 10.6151
R1613 B.n179 B.n178 10.6151
R1614 B.n182 B.n179 10.6151
R1615 B.n183 B.n182 10.6151
R1616 B.n186 B.n183 10.6151
R1617 B.n187 B.n186 10.6151
R1618 B.n190 B.n187 10.6151
R1619 B.n191 B.n190 10.6151
R1620 B.n194 B.n191 10.6151
R1621 B.n195 B.n194 10.6151
R1622 B.n198 B.n195 10.6151
R1623 B.n199 B.n198 10.6151
R1624 B.n202 B.n199 10.6151
R1625 B.n203 B.n202 10.6151
R1626 B.n206 B.n203 10.6151
R1627 B.n207 B.n206 10.6151
R1628 B.n210 B.n207 10.6151
R1629 B.n211 B.n210 10.6151
R1630 B.n214 B.n211 10.6151
R1631 B.n215 B.n214 10.6151
R1632 B.n218 B.n215 10.6151
R1633 B.n219 B.n218 10.6151
R1634 B.n222 B.n219 10.6151
R1635 B.n227 B.n224 10.6151
R1636 B.n228 B.n227 10.6151
R1637 B.n231 B.n228 10.6151
R1638 B.n232 B.n231 10.6151
R1639 B.n235 B.n232 10.6151
R1640 B.n236 B.n235 10.6151
R1641 B.n239 B.n236 10.6151
R1642 B.n240 B.n239 10.6151
R1643 B.n244 B.n243 10.6151
R1644 B.n247 B.n244 10.6151
R1645 B.n248 B.n247 10.6151
R1646 B.n251 B.n248 10.6151
R1647 B.n252 B.n251 10.6151
R1648 B.n255 B.n252 10.6151
R1649 B.n256 B.n255 10.6151
R1650 B.n259 B.n256 10.6151
R1651 B.n260 B.n259 10.6151
R1652 B.n263 B.n260 10.6151
R1653 B.n264 B.n263 10.6151
R1654 B.n267 B.n264 10.6151
R1655 B.n268 B.n267 10.6151
R1656 B.n271 B.n268 10.6151
R1657 B.n272 B.n271 10.6151
R1658 B.n275 B.n272 10.6151
R1659 B.n276 B.n275 10.6151
R1660 B.n279 B.n276 10.6151
R1661 B.n280 B.n279 10.6151
R1662 B.n283 B.n280 10.6151
R1663 B.n284 B.n283 10.6151
R1664 B.n287 B.n284 10.6151
R1665 B.n288 B.n287 10.6151
R1666 B.n291 B.n288 10.6151
R1667 B.n292 B.n291 10.6151
R1668 B.n295 B.n292 10.6151
R1669 B.n296 B.n295 10.6151
R1670 B.n299 B.n296 10.6151
R1671 B.n300 B.n299 10.6151
R1672 B.n303 B.n300 10.6151
R1673 B.n304 B.n303 10.6151
R1674 B.n307 B.n304 10.6151
R1675 B.n308 B.n307 10.6151
R1676 B.n311 B.n308 10.6151
R1677 B.n312 B.n311 10.6151
R1678 B.n315 B.n312 10.6151
R1679 B.n316 B.n315 10.6151
R1680 B.n319 B.n316 10.6151
R1681 B.n320 B.n319 10.6151
R1682 B.n323 B.n320 10.6151
R1683 B.n324 B.n323 10.6151
R1684 B.n327 B.n324 10.6151
R1685 B.n328 B.n327 10.6151
R1686 B.n331 B.n328 10.6151
R1687 B.n332 B.n331 10.6151
R1688 B.n840 B.n332 10.6151
R1689 B.n779 B.t4 10.3969
R1690 B.n915 B.t0 10.3969
R1691 B.n398 B.t13 9.24177
R1692 B.t5 B.n374 9.24177
R1693 B.t1 B.n44 9.24177
R1694 B.t9 B.n858 9.24177
R1695 B.n927 B.n0 8.11757
R1696 B.n927 B.n1 8.11757
R1697 B.n577 B.n463 6.5566
R1698 B.n561 B.n560 6.5566
R1699 B.n224 B.n223 6.5566
R1700 B.n240 B.n130 6.5566
R1701 B.n580 B.n463 4.05904
R1702 B.n560 B.n559 4.05904
R1703 B.n223 B.n222 4.05904
R1704 B.n243 B.n130 4.05904
R1705 B.n366 B.t3 3.46598
R1706 B.t7 B.n890 3.46598
R1707 VN.n4 VN.t5 213.773
R1708 VN.n25 VN.t6 213.773
R1709 VN.n5 VN.t4 182.339
R1710 VN.n12 VN.t3 182.339
R1711 VN.n19 VN.t2 182.339
R1712 VN.n26 VN.t7 182.339
R1713 VN.n33 VN.t0 182.339
R1714 VN.n40 VN.t1 182.339
R1715 VN.n39 VN.n21 161.3
R1716 VN.n38 VN.n37 161.3
R1717 VN.n36 VN.n22 161.3
R1718 VN.n35 VN.n34 161.3
R1719 VN.n32 VN.n23 161.3
R1720 VN.n31 VN.n30 161.3
R1721 VN.n29 VN.n24 161.3
R1722 VN.n28 VN.n27 161.3
R1723 VN.n18 VN.n0 161.3
R1724 VN.n17 VN.n16 161.3
R1725 VN.n15 VN.n1 161.3
R1726 VN.n14 VN.n13 161.3
R1727 VN.n11 VN.n2 161.3
R1728 VN.n10 VN.n9 161.3
R1729 VN.n8 VN.n3 161.3
R1730 VN.n7 VN.n6 161.3
R1731 VN.n20 VN.n19 87.5128
R1732 VN.n41 VN.n40 87.5128
R1733 VN.n10 VN.n3 56.5193
R1734 VN.n31 VN.n24 56.5193
R1735 VN.n5 VN.n4 53.8955
R1736 VN.n26 VN.n25 53.8955
R1737 VN.n17 VN.n1 50.2061
R1738 VN.n38 VN.n22 50.2061
R1739 VN VN.n41 48.8997
R1740 VN.n18 VN.n17 30.7807
R1741 VN.n39 VN.n38 30.7807
R1742 VN.n6 VN.n3 24.4675
R1743 VN.n11 VN.n10 24.4675
R1744 VN.n13 VN.n1 24.4675
R1745 VN.n27 VN.n24 24.4675
R1746 VN.n34 VN.n22 24.4675
R1747 VN.n32 VN.n31 24.4675
R1748 VN.n19 VN.n18 23.2442
R1749 VN.n40 VN.n39 23.2442
R1750 VN.n6 VN.n5 15.9041
R1751 VN.n12 VN.n11 15.9041
R1752 VN.n27 VN.n26 15.9041
R1753 VN.n33 VN.n32 15.9041
R1754 VN.n28 VN.n25 12.7761
R1755 VN.n7 VN.n4 12.7761
R1756 VN.n13 VN.n12 8.56395
R1757 VN.n34 VN.n33 8.56395
R1758 VN.n41 VN.n21 0.278367
R1759 VN.n20 VN.n0 0.278367
R1760 VN.n37 VN.n21 0.189894
R1761 VN.n37 VN.n36 0.189894
R1762 VN.n36 VN.n35 0.189894
R1763 VN.n35 VN.n23 0.189894
R1764 VN.n30 VN.n23 0.189894
R1765 VN.n30 VN.n29 0.189894
R1766 VN.n29 VN.n28 0.189894
R1767 VN.n8 VN.n7 0.189894
R1768 VN.n9 VN.n8 0.189894
R1769 VN.n9 VN.n2 0.189894
R1770 VN.n14 VN.n2 0.189894
R1771 VN.n15 VN.n14 0.189894
R1772 VN.n16 VN.n15 0.189894
R1773 VN.n16 VN.n0 0.189894
R1774 VN VN.n20 0.153454
R1775 VDD2.n2 VDD2.n1 66.011
R1776 VDD2.n2 VDD2.n0 66.011
R1777 VDD2 VDD2.n5 66.0082
R1778 VDD2.n4 VDD2.n3 65.1399
R1779 VDD2.n4 VDD2.n2 43.9265
R1780 VDD2.n5 VDD2.t0 1.43841
R1781 VDD2.n5 VDD2.t1 1.43841
R1782 VDD2.n3 VDD2.t6 1.43841
R1783 VDD2.n3 VDD2.t7 1.43841
R1784 VDD2.n1 VDD2.t4 1.43841
R1785 VDD2.n1 VDD2.t5 1.43841
R1786 VDD2.n0 VDD2.t2 1.43841
R1787 VDD2.n0 VDD2.t3 1.43841
R1788 VDD2 VDD2.n4 0.985414
C0 VDD1 VTAIL 8.91512f
C1 VDD1 VP 9.409019f
C2 VTAIL VN 9.19303f
C3 VP VN 7.03866f
C4 VDD1 VDD2 1.3704f
C5 VDD2 VN 9.12367f
C6 VTAIL VP 9.20714f
C7 VTAIL VDD2 8.96431f
C8 VP VDD2 0.436502f
C9 VDD1 VN 0.150149f
C10 VDD2 B 4.729352f
C11 VDD1 B 5.080945f
C12 VTAIL B 10.973066f
C13 VN B 12.734929f
C14 VP B 11.160074f
C15 VDD2.t2 B 0.268946f
C16 VDD2.t3 B 0.268946f
C17 VDD2.n0 B 2.43064f
C18 VDD2.t4 B 0.268946f
C19 VDD2.t5 B 0.268946f
C20 VDD2.n1 B 2.43064f
C21 VDD2.n2 B 2.88955f
C22 VDD2.t6 B 0.268946f
C23 VDD2.t7 B 0.268946f
C24 VDD2.n3 B 2.42503f
C25 VDD2.n4 B 2.77627f
C26 VDD2.t0 B 0.268946f
C27 VDD2.t1 B 0.268946f
C28 VDD2.n5 B 2.4306f
C29 VN.n0 B 0.035929f
C30 VN.t2 B 1.86767f
C31 VN.n1 B 0.050017f
C32 VN.n2 B 0.027252f
C33 VN.t3 B 1.86767f
C34 VN.n3 B 0.039783f
C35 VN.t5 B 1.98394f
C36 VN.n4 B 0.732531f
C37 VN.t4 B 1.86767f
C38 VN.n5 B 0.727889f
C39 VN.n6 B 0.042013f
C40 VN.n7 B 0.199652f
C41 VN.n8 B 0.027252f
C42 VN.n9 B 0.027252f
C43 VN.n10 B 0.039783f
C44 VN.n11 B 0.042013f
C45 VN.n12 B 0.663074f
C46 VN.n13 B 0.03449f
C47 VN.n14 B 0.027252f
C48 VN.n15 B 0.027252f
C49 VN.n16 B 0.027252f
C50 VN.n17 B 0.025744f
C51 VN.n18 B 0.05334f
C52 VN.n19 B 0.744742f
C53 VN.n20 B 0.029626f
C54 VN.n21 B 0.035929f
C55 VN.t1 B 1.86767f
C56 VN.n22 B 0.050017f
C57 VN.n23 B 0.027252f
C58 VN.t0 B 1.86767f
C59 VN.n24 B 0.039783f
C60 VN.t6 B 1.98394f
C61 VN.n25 B 0.732531f
C62 VN.t7 B 1.86767f
C63 VN.n26 B 0.727889f
C64 VN.n27 B 0.042013f
C65 VN.n28 B 0.199652f
C66 VN.n29 B 0.027252f
C67 VN.n30 B 0.027252f
C68 VN.n31 B 0.039783f
C69 VN.n32 B 0.042013f
C70 VN.n33 B 0.663074f
C71 VN.n34 B 0.03449f
C72 VN.n35 B 0.027252f
C73 VN.n36 B 0.027252f
C74 VN.n37 B 0.027252f
C75 VN.n38 B 0.025744f
C76 VN.n39 B 0.05334f
C77 VN.n40 B 0.744742f
C78 VN.n41 B 1.45403f
C79 VTAIL.t2 B 0.206374f
C80 VTAIL.t7 B 0.206374f
C81 VTAIL.n0 B 1.81007f
C82 VTAIL.n1 B 0.292915f
C83 VTAIL.t0 B 2.31047f
C84 VTAIL.n2 B 0.380503f
C85 VTAIL.t8 B 2.31047f
C86 VTAIL.n3 B 0.380503f
C87 VTAIL.t9 B 0.206374f
C88 VTAIL.t10 B 0.206374f
C89 VTAIL.n4 B 1.81007f
C90 VTAIL.n5 B 0.402625f
C91 VTAIL.t11 B 2.31047f
C92 VTAIL.n6 B 1.44812f
C93 VTAIL.t5 B 2.31047f
C94 VTAIL.n7 B 1.44812f
C95 VTAIL.t3 B 0.206374f
C96 VTAIL.t6 B 0.206374f
C97 VTAIL.n8 B 1.81007f
C98 VTAIL.n9 B 0.402623f
C99 VTAIL.t4 B 2.31047f
C100 VTAIL.n10 B 0.380501f
C101 VTAIL.t14 B 2.31047f
C102 VTAIL.n11 B 0.380501f
C103 VTAIL.t12 B 0.206374f
C104 VTAIL.t15 B 0.206374f
C105 VTAIL.n12 B 1.81007f
C106 VTAIL.n13 B 0.402623f
C107 VTAIL.t13 B 2.31047f
C108 VTAIL.n14 B 1.44812f
C109 VTAIL.t1 B 2.31047f
C110 VTAIL.n15 B 1.44456f
C111 VDD1.t4 B 0.270553f
C112 VDD1.t0 B 0.270553f
C113 VDD1.n0 B 2.44601f
C114 VDD1.t7 B 0.270553f
C115 VDD1.t3 B 0.270553f
C116 VDD1.n1 B 2.44516f
C117 VDD1.t1 B 0.270553f
C118 VDD1.t5 B 0.270553f
C119 VDD1.n2 B 2.44516f
C120 VDD1.n3 B 2.959f
C121 VDD1.t2 B 0.270553f
C122 VDD1.t6 B 0.270553f
C123 VDD1.n4 B 2.43952f
C124 VDD1.n5 B 2.8232f
C125 VP.n0 B 0.03641f
C126 VP.t7 B 1.89268f
C127 VP.n1 B 0.050687f
C128 VP.n2 B 0.027617f
C129 VP.t5 B 1.89268f
C130 VP.n3 B 0.040316f
C131 VP.n4 B 0.027617f
C132 VP.t6 B 1.89268f
C133 VP.n5 B 0.026089f
C134 VP.n6 B 0.03641f
C135 VP.t2 B 1.89268f
C136 VP.n7 B 0.050687f
C137 VP.n8 B 0.027617f
C138 VP.t0 B 1.89268f
C139 VP.n9 B 0.040316f
C140 VP.t1 B 2.01051f
C141 VP.n10 B 0.742341f
C142 VP.t3 B 1.89268f
C143 VP.n11 B 0.737637f
C144 VP.n12 B 0.042576f
C145 VP.n13 B 0.202326f
C146 VP.n14 B 0.027617f
C147 VP.n15 B 0.027617f
C148 VP.n16 B 0.040316f
C149 VP.n17 B 0.042576f
C150 VP.n18 B 0.671954f
C151 VP.n19 B 0.034952f
C152 VP.n20 B 0.027617f
C153 VP.n21 B 0.027617f
C154 VP.n22 B 0.027617f
C155 VP.n23 B 0.026089f
C156 VP.n24 B 0.054054f
C157 VP.n25 B 0.754716f
C158 VP.n26 B 1.45859f
C159 VP.n27 B 1.47901f
C160 VP.t4 B 1.89268f
C161 VP.n28 B 0.754716f
C162 VP.n29 B 0.054054f
C163 VP.n30 B 0.03641f
C164 VP.n31 B 0.027617f
C165 VP.n32 B 0.027617f
C166 VP.n33 B 0.050687f
C167 VP.n34 B 0.034952f
C168 VP.n35 B 0.671954f
C169 VP.n36 B 0.042576f
C170 VP.n37 B 0.027617f
C171 VP.n38 B 0.027617f
C172 VP.n39 B 0.027617f
C173 VP.n40 B 0.040316f
C174 VP.n41 B 0.042576f
C175 VP.n42 B 0.671954f
C176 VP.n43 B 0.034952f
C177 VP.n44 B 0.027617f
C178 VP.n45 B 0.027617f
C179 VP.n46 B 0.027617f
C180 VP.n47 B 0.026089f
C181 VP.n48 B 0.054054f
C182 VP.n49 B 0.754716f
C183 VP.n50 B 0.030023f
.ends

