* NGSPICE file created from diff_pair_sample_0654.ext - technology: sky130A

.subckt diff_pair_sample_0654 VTAIL VN VP B VDD2 VDD1
X0 B.t17 B.t15 B.t16 B.t9 sky130_fd_pr__nfet_01v8 ad=3.8961 pd=20.76 as=0 ps=0 w=9.99 l=1.29
X1 VDD2.t3 VN.t0 VTAIL.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=1.64835 pd=10.32 as=3.8961 ps=20.76 w=9.99 l=1.29
X2 VTAIL.t3 VP.t0 VDD1.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=3.8961 pd=20.76 as=1.64835 ps=10.32 w=9.99 l=1.29
X3 B.t14 B.t12 B.t13 B.t5 sky130_fd_pr__nfet_01v8 ad=3.8961 pd=20.76 as=0 ps=0 w=9.99 l=1.29
X4 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=3.8961 pd=20.76 as=0 ps=0 w=9.99 l=1.29
X5 VDD1.t2 VP.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.64835 pd=10.32 as=3.8961 ps=20.76 w=9.99 l=1.29
X6 VTAIL.t1 VP.t2 VDD1.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=3.8961 pd=20.76 as=1.64835 ps=10.32 w=9.99 l=1.29
X7 VDD1.t0 VP.t3 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.64835 pd=10.32 as=3.8961 ps=20.76 w=9.99 l=1.29
X8 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=3.8961 pd=20.76 as=0 ps=0 w=9.99 l=1.29
X9 VDD2.t2 VN.t1 VTAIL.t7 B.t0 sky130_fd_pr__nfet_01v8 ad=1.64835 pd=10.32 as=3.8961 ps=20.76 w=9.99 l=1.29
X10 VTAIL.t4 VN.t2 VDD2.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=3.8961 pd=20.76 as=1.64835 ps=10.32 w=9.99 l=1.29
X11 VTAIL.t5 VN.t3 VDD2.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=3.8961 pd=20.76 as=1.64835 ps=10.32 w=9.99 l=1.29
R0 B.n436 B.n88 585
R1 B.n88 B.n43 585
R2 B.n438 B.n437 585
R3 B.n440 B.n87 585
R4 B.n443 B.n442 585
R5 B.n444 B.n86 585
R6 B.n446 B.n445 585
R7 B.n448 B.n85 585
R8 B.n451 B.n450 585
R9 B.n452 B.n84 585
R10 B.n454 B.n453 585
R11 B.n456 B.n83 585
R12 B.n459 B.n458 585
R13 B.n460 B.n82 585
R14 B.n462 B.n461 585
R15 B.n464 B.n81 585
R16 B.n467 B.n466 585
R17 B.n468 B.n80 585
R18 B.n470 B.n469 585
R19 B.n472 B.n79 585
R20 B.n475 B.n474 585
R21 B.n476 B.n78 585
R22 B.n478 B.n477 585
R23 B.n480 B.n77 585
R24 B.n483 B.n482 585
R25 B.n484 B.n76 585
R26 B.n486 B.n485 585
R27 B.n488 B.n75 585
R28 B.n491 B.n490 585
R29 B.n492 B.n74 585
R30 B.n494 B.n493 585
R31 B.n496 B.n73 585
R32 B.n499 B.n498 585
R33 B.n500 B.n72 585
R34 B.n502 B.n501 585
R35 B.n504 B.n71 585
R36 B.n507 B.n506 585
R37 B.n509 B.n68 585
R38 B.n511 B.n510 585
R39 B.n513 B.n67 585
R40 B.n516 B.n515 585
R41 B.n517 B.n66 585
R42 B.n519 B.n518 585
R43 B.n521 B.n65 585
R44 B.n524 B.n523 585
R45 B.n525 B.n62 585
R46 B.n528 B.n527 585
R47 B.n530 B.n61 585
R48 B.n533 B.n532 585
R49 B.n534 B.n60 585
R50 B.n536 B.n535 585
R51 B.n538 B.n59 585
R52 B.n541 B.n540 585
R53 B.n542 B.n58 585
R54 B.n544 B.n543 585
R55 B.n546 B.n57 585
R56 B.n549 B.n548 585
R57 B.n550 B.n56 585
R58 B.n552 B.n551 585
R59 B.n554 B.n55 585
R60 B.n557 B.n556 585
R61 B.n558 B.n54 585
R62 B.n560 B.n559 585
R63 B.n562 B.n53 585
R64 B.n565 B.n564 585
R65 B.n566 B.n52 585
R66 B.n568 B.n567 585
R67 B.n570 B.n51 585
R68 B.n573 B.n572 585
R69 B.n574 B.n50 585
R70 B.n576 B.n575 585
R71 B.n578 B.n49 585
R72 B.n581 B.n580 585
R73 B.n582 B.n48 585
R74 B.n584 B.n583 585
R75 B.n586 B.n47 585
R76 B.n589 B.n588 585
R77 B.n590 B.n46 585
R78 B.n592 B.n591 585
R79 B.n594 B.n45 585
R80 B.n597 B.n596 585
R81 B.n598 B.n44 585
R82 B.n435 B.n42 585
R83 B.n601 B.n42 585
R84 B.n434 B.n41 585
R85 B.n602 B.n41 585
R86 B.n433 B.n40 585
R87 B.n603 B.n40 585
R88 B.n432 B.n431 585
R89 B.n431 B.n36 585
R90 B.n430 B.n35 585
R91 B.n609 B.n35 585
R92 B.n429 B.n34 585
R93 B.n610 B.n34 585
R94 B.n428 B.n33 585
R95 B.n611 B.n33 585
R96 B.n427 B.n426 585
R97 B.n426 B.n29 585
R98 B.n425 B.n28 585
R99 B.n617 B.n28 585
R100 B.n424 B.n27 585
R101 B.n618 B.n27 585
R102 B.n423 B.n26 585
R103 B.n619 B.n26 585
R104 B.n422 B.n421 585
R105 B.n421 B.n22 585
R106 B.n420 B.n21 585
R107 B.n625 B.n21 585
R108 B.n419 B.n20 585
R109 B.n626 B.n20 585
R110 B.n418 B.n19 585
R111 B.n627 B.n19 585
R112 B.n417 B.n416 585
R113 B.n416 B.n15 585
R114 B.n415 B.n14 585
R115 B.n633 B.n14 585
R116 B.n414 B.n13 585
R117 B.n634 B.n13 585
R118 B.n413 B.n12 585
R119 B.n635 B.n12 585
R120 B.n412 B.n411 585
R121 B.n411 B.n410 585
R122 B.n409 B.n408 585
R123 B.n409 B.n8 585
R124 B.n407 B.n7 585
R125 B.n642 B.n7 585
R126 B.n406 B.n6 585
R127 B.n643 B.n6 585
R128 B.n405 B.n5 585
R129 B.n644 B.n5 585
R130 B.n404 B.n403 585
R131 B.n403 B.n4 585
R132 B.n402 B.n89 585
R133 B.n402 B.n401 585
R134 B.n392 B.n90 585
R135 B.n91 B.n90 585
R136 B.n394 B.n393 585
R137 B.n395 B.n394 585
R138 B.n391 B.n96 585
R139 B.n96 B.n95 585
R140 B.n390 B.n389 585
R141 B.n389 B.n388 585
R142 B.n98 B.n97 585
R143 B.n99 B.n98 585
R144 B.n381 B.n380 585
R145 B.n382 B.n381 585
R146 B.n379 B.n103 585
R147 B.n107 B.n103 585
R148 B.n378 B.n377 585
R149 B.n377 B.n376 585
R150 B.n105 B.n104 585
R151 B.n106 B.n105 585
R152 B.n369 B.n368 585
R153 B.n370 B.n369 585
R154 B.n367 B.n112 585
R155 B.n112 B.n111 585
R156 B.n366 B.n365 585
R157 B.n365 B.n364 585
R158 B.n114 B.n113 585
R159 B.n115 B.n114 585
R160 B.n357 B.n356 585
R161 B.n358 B.n357 585
R162 B.n355 B.n119 585
R163 B.n123 B.n119 585
R164 B.n354 B.n353 585
R165 B.n353 B.n352 585
R166 B.n121 B.n120 585
R167 B.n122 B.n121 585
R168 B.n345 B.n344 585
R169 B.n346 B.n345 585
R170 B.n343 B.n128 585
R171 B.n128 B.n127 585
R172 B.n342 B.n341 585
R173 B.n341 B.n340 585
R174 B.n337 B.n132 585
R175 B.n336 B.n335 585
R176 B.n333 B.n133 585
R177 B.n333 B.n131 585
R178 B.n332 B.n331 585
R179 B.n330 B.n329 585
R180 B.n328 B.n135 585
R181 B.n326 B.n325 585
R182 B.n324 B.n136 585
R183 B.n323 B.n322 585
R184 B.n320 B.n137 585
R185 B.n318 B.n317 585
R186 B.n316 B.n138 585
R187 B.n315 B.n314 585
R188 B.n312 B.n139 585
R189 B.n310 B.n309 585
R190 B.n308 B.n140 585
R191 B.n307 B.n306 585
R192 B.n304 B.n141 585
R193 B.n302 B.n301 585
R194 B.n300 B.n142 585
R195 B.n299 B.n298 585
R196 B.n296 B.n143 585
R197 B.n294 B.n293 585
R198 B.n292 B.n144 585
R199 B.n291 B.n290 585
R200 B.n288 B.n145 585
R201 B.n286 B.n285 585
R202 B.n284 B.n146 585
R203 B.n283 B.n282 585
R204 B.n280 B.n147 585
R205 B.n278 B.n277 585
R206 B.n276 B.n148 585
R207 B.n275 B.n274 585
R208 B.n272 B.n149 585
R209 B.n270 B.n269 585
R210 B.n268 B.n150 585
R211 B.n266 B.n265 585
R212 B.n263 B.n153 585
R213 B.n261 B.n260 585
R214 B.n259 B.n154 585
R215 B.n258 B.n257 585
R216 B.n255 B.n155 585
R217 B.n253 B.n252 585
R218 B.n251 B.n156 585
R219 B.n250 B.n249 585
R220 B.n247 B.n246 585
R221 B.n245 B.n244 585
R222 B.n243 B.n161 585
R223 B.n241 B.n240 585
R224 B.n239 B.n162 585
R225 B.n238 B.n237 585
R226 B.n235 B.n163 585
R227 B.n233 B.n232 585
R228 B.n231 B.n164 585
R229 B.n230 B.n229 585
R230 B.n227 B.n165 585
R231 B.n225 B.n224 585
R232 B.n223 B.n166 585
R233 B.n222 B.n221 585
R234 B.n219 B.n167 585
R235 B.n217 B.n216 585
R236 B.n215 B.n168 585
R237 B.n214 B.n213 585
R238 B.n211 B.n169 585
R239 B.n209 B.n208 585
R240 B.n207 B.n170 585
R241 B.n206 B.n205 585
R242 B.n203 B.n171 585
R243 B.n201 B.n200 585
R244 B.n199 B.n172 585
R245 B.n198 B.n197 585
R246 B.n195 B.n173 585
R247 B.n193 B.n192 585
R248 B.n191 B.n174 585
R249 B.n190 B.n189 585
R250 B.n187 B.n175 585
R251 B.n185 B.n184 585
R252 B.n183 B.n176 585
R253 B.n182 B.n181 585
R254 B.n179 B.n177 585
R255 B.n130 B.n129 585
R256 B.n339 B.n338 585
R257 B.n340 B.n339 585
R258 B.n126 B.n125 585
R259 B.n127 B.n126 585
R260 B.n348 B.n347 585
R261 B.n347 B.n346 585
R262 B.n349 B.n124 585
R263 B.n124 B.n122 585
R264 B.n351 B.n350 585
R265 B.n352 B.n351 585
R266 B.n118 B.n117 585
R267 B.n123 B.n118 585
R268 B.n360 B.n359 585
R269 B.n359 B.n358 585
R270 B.n361 B.n116 585
R271 B.n116 B.n115 585
R272 B.n363 B.n362 585
R273 B.n364 B.n363 585
R274 B.n110 B.n109 585
R275 B.n111 B.n110 585
R276 B.n372 B.n371 585
R277 B.n371 B.n370 585
R278 B.n373 B.n108 585
R279 B.n108 B.n106 585
R280 B.n375 B.n374 585
R281 B.n376 B.n375 585
R282 B.n102 B.n101 585
R283 B.n107 B.n102 585
R284 B.n384 B.n383 585
R285 B.n383 B.n382 585
R286 B.n385 B.n100 585
R287 B.n100 B.n99 585
R288 B.n387 B.n386 585
R289 B.n388 B.n387 585
R290 B.n94 B.n93 585
R291 B.n95 B.n94 585
R292 B.n397 B.n396 585
R293 B.n396 B.n395 585
R294 B.n398 B.n92 585
R295 B.n92 B.n91 585
R296 B.n400 B.n399 585
R297 B.n401 B.n400 585
R298 B.n3 B.n0 585
R299 B.n4 B.n3 585
R300 B.n641 B.n1 585
R301 B.n642 B.n641 585
R302 B.n640 B.n639 585
R303 B.n640 B.n8 585
R304 B.n638 B.n9 585
R305 B.n410 B.n9 585
R306 B.n637 B.n636 585
R307 B.n636 B.n635 585
R308 B.n11 B.n10 585
R309 B.n634 B.n11 585
R310 B.n632 B.n631 585
R311 B.n633 B.n632 585
R312 B.n630 B.n16 585
R313 B.n16 B.n15 585
R314 B.n629 B.n628 585
R315 B.n628 B.n627 585
R316 B.n18 B.n17 585
R317 B.n626 B.n18 585
R318 B.n624 B.n623 585
R319 B.n625 B.n624 585
R320 B.n622 B.n23 585
R321 B.n23 B.n22 585
R322 B.n621 B.n620 585
R323 B.n620 B.n619 585
R324 B.n25 B.n24 585
R325 B.n618 B.n25 585
R326 B.n616 B.n615 585
R327 B.n617 B.n616 585
R328 B.n614 B.n30 585
R329 B.n30 B.n29 585
R330 B.n613 B.n612 585
R331 B.n612 B.n611 585
R332 B.n32 B.n31 585
R333 B.n610 B.n32 585
R334 B.n608 B.n607 585
R335 B.n609 B.n608 585
R336 B.n606 B.n37 585
R337 B.n37 B.n36 585
R338 B.n605 B.n604 585
R339 B.n604 B.n603 585
R340 B.n39 B.n38 585
R341 B.n602 B.n39 585
R342 B.n600 B.n599 585
R343 B.n601 B.n600 585
R344 B.n645 B.n644 585
R345 B.n643 B.n2 585
R346 B.n600 B.n44 482.89
R347 B.n88 B.n42 482.89
R348 B.n341 B.n130 482.89
R349 B.n339 B.n132 482.89
R350 B.n63 B.t8 391.197
R351 B.n69 B.t15 391.197
R352 B.n157 B.t4 391.197
R353 B.n151 B.t12 391.197
R354 B.n69 B.t16 278.872
R355 B.n157 B.t7 278.872
R356 B.n63 B.t10 278.872
R357 B.n151 B.t14 278.872
R358 B.n439 B.n43 256.663
R359 B.n441 B.n43 256.663
R360 B.n447 B.n43 256.663
R361 B.n449 B.n43 256.663
R362 B.n455 B.n43 256.663
R363 B.n457 B.n43 256.663
R364 B.n463 B.n43 256.663
R365 B.n465 B.n43 256.663
R366 B.n471 B.n43 256.663
R367 B.n473 B.n43 256.663
R368 B.n479 B.n43 256.663
R369 B.n481 B.n43 256.663
R370 B.n487 B.n43 256.663
R371 B.n489 B.n43 256.663
R372 B.n495 B.n43 256.663
R373 B.n497 B.n43 256.663
R374 B.n503 B.n43 256.663
R375 B.n505 B.n43 256.663
R376 B.n512 B.n43 256.663
R377 B.n514 B.n43 256.663
R378 B.n520 B.n43 256.663
R379 B.n522 B.n43 256.663
R380 B.n529 B.n43 256.663
R381 B.n531 B.n43 256.663
R382 B.n537 B.n43 256.663
R383 B.n539 B.n43 256.663
R384 B.n545 B.n43 256.663
R385 B.n547 B.n43 256.663
R386 B.n553 B.n43 256.663
R387 B.n555 B.n43 256.663
R388 B.n561 B.n43 256.663
R389 B.n563 B.n43 256.663
R390 B.n569 B.n43 256.663
R391 B.n571 B.n43 256.663
R392 B.n577 B.n43 256.663
R393 B.n579 B.n43 256.663
R394 B.n585 B.n43 256.663
R395 B.n587 B.n43 256.663
R396 B.n593 B.n43 256.663
R397 B.n595 B.n43 256.663
R398 B.n334 B.n131 256.663
R399 B.n134 B.n131 256.663
R400 B.n327 B.n131 256.663
R401 B.n321 B.n131 256.663
R402 B.n319 B.n131 256.663
R403 B.n313 B.n131 256.663
R404 B.n311 B.n131 256.663
R405 B.n305 B.n131 256.663
R406 B.n303 B.n131 256.663
R407 B.n297 B.n131 256.663
R408 B.n295 B.n131 256.663
R409 B.n289 B.n131 256.663
R410 B.n287 B.n131 256.663
R411 B.n281 B.n131 256.663
R412 B.n279 B.n131 256.663
R413 B.n273 B.n131 256.663
R414 B.n271 B.n131 256.663
R415 B.n264 B.n131 256.663
R416 B.n262 B.n131 256.663
R417 B.n256 B.n131 256.663
R418 B.n254 B.n131 256.663
R419 B.n248 B.n131 256.663
R420 B.n160 B.n131 256.663
R421 B.n242 B.n131 256.663
R422 B.n236 B.n131 256.663
R423 B.n234 B.n131 256.663
R424 B.n228 B.n131 256.663
R425 B.n226 B.n131 256.663
R426 B.n220 B.n131 256.663
R427 B.n218 B.n131 256.663
R428 B.n212 B.n131 256.663
R429 B.n210 B.n131 256.663
R430 B.n204 B.n131 256.663
R431 B.n202 B.n131 256.663
R432 B.n196 B.n131 256.663
R433 B.n194 B.n131 256.663
R434 B.n188 B.n131 256.663
R435 B.n186 B.n131 256.663
R436 B.n180 B.n131 256.663
R437 B.n178 B.n131 256.663
R438 B.n647 B.n646 256.663
R439 B.n70 B.t17 247.453
R440 B.n158 B.t6 247.453
R441 B.n64 B.t11 247.453
R442 B.n152 B.t13 247.453
R443 B.n596 B.n594 163.367
R444 B.n592 B.n46 163.367
R445 B.n588 B.n586 163.367
R446 B.n584 B.n48 163.367
R447 B.n580 B.n578 163.367
R448 B.n576 B.n50 163.367
R449 B.n572 B.n570 163.367
R450 B.n568 B.n52 163.367
R451 B.n564 B.n562 163.367
R452 B.n560 B.n54 163.367
R453 B.n556 B.n554 163.367
R454 B.n552 B.n56 163.367
R455 B.n548 B.n546 163.367
R456 B.n544 B.n58 163.367
R457 B.n540 B.n538 163.367
R458 B.n536 B.n60 163.367
R459 B.n532 B.n530 163.367
R460 B.n528 B.n62 163.367
R461 B.n523 B.n521 163.367
R462 B.n519 B.n66 163.367
R463 B.n515 B.n513 163.367
R464 B.n511 B.n68 163.367
R465 B.n506 B.n504 163.367
R466 B.n502 B.n72 163.367
R467 B.n498 B.n496 163.367
R468 B.n494 B.n74 163.367
R469 B.n490 B.n488 163.367
R470 B.n486 B.n76 163.367
R471 B.n482 B.n480 163.367
R472 B.n478 B.n78 163.367
R473 B.n474 B.n472 163.367
R474 B.n470 B.n80 163.367
R475 B.n466 B.n464 163.367
R476 B.n462 B.n82 163.367
R477 B.n458 B.n456 163.367
R478 B.n454 B.n84 163.367
R479 B.n450 B.n448 163.367
R480 B.n446 B.n86 163.367
R481 B.n442 B.n440 163.367
R482 B.n438 B.n88 163.367
R483 B.n341 B.n128 163.367
R484 B.n345 B.n128 163.367
R485 B.n345 B.n121 163.367
R486 B.n353 B.n121 163.367
R487 B.n353 B.n119 163.367
R488 B.n357 B.n119 163.367
R489 B.n357 B.n114 163.367
R490 B.n365 B.n114 163.367
R491 B.n365 B.n112 163.367
R492 B.n369 B.n112 163.367
R493 B.n369 B.n105 163.367
R494 B.n377 B.n105 163.367
R495 B.n377 B.n103 163.367
R496 B.n381 B.n103 163.367
R497 B.n381 B.n98 163.367
R498 B.n389 B.n98 163.367
R499 B.n389 B.n96 163.367
R500 B.n394 B.n96 163.367
R501 B.n394 B.n90 163.367
R502 B.n402 B.n90 163.367
R503 B.n403 B.n402 163.367
R504 B.n403 B.n5 163.367
R505 B.n6 B.n5 163.367
R506 B.n7 B.n6 163.367
R507 B.n409 B.n7 163.367
R508 B.n411 B.n409 163.367
R509 B.n411 B.n12 163.367
R510 B.n13 B.n12 163.367
R511 B.n14 B.n13 163.367
R512 B.n416 B.n14 163.367
R513 B.n416 B.n19 163.367
R514 B.n20 B.n19 163.367
R515 B.n21 B.n20 163.367
R516 B.n421 B.n21 163.367
R517 B.n421 B.n26 163.367
R518 B.n27 B.n26 163.367
R519 B.n28 B.n27 163.367
R520 B.n426 B.n28 163.367
R521 B.n426 B.n33 163.367
R522 B.n34 B.n33 163.367
R523 B.n35 B.n34 163.367
R524 B.n431 B.n35 163.367
R525 B.n431 B.n40 163.367
R526 B.n41 B.n40 163.367
R527 B.n42 B.n41 163.367
R528 B.n335 B.n333 163.367
R529 B.n333 B.n332 163.367
R530 B.n329 B.n328 163.367
R531 B.n326 B.n136 163.367
R532 B.n322 B.n320 163.367
R533 B.n318 B.n138 163.367
R534 B.n314 B.n312 163.367
R535 B.n310 B.n140 163.367
R536 B.n306 B.n304 163.367
R537 B.n302 B.n142 163.367
R538 B.n298 B.n296 163.367
R539 B.n294 B.n144 163.367
R540 B.n290 B.n288 163.367
R541 B.n286 B.n146 163.367
R542 B.n282 B.n280 163.367
R543 B.n278 B.n148 163.367
R544 B.n274 B.n272 163.367
R545 B.n270 B.n150 163.367
R546 B.n265 B.n263 163.367
R547 B.n261 B.n154 163.367
R548 B.n257 B.n255 163.367
R549 B.n253 B.n156 163.367
R550 B.n249 B.n247 163.367
R551 B.n244 B.n243 163.367
R552 B.n241 B.n162 163.367
R553 B.n237 B.n235 163.367
R554 B.n233 B.n164 163.367
R555 B.n229 B.n227 163.367
R556 B.n225 B.n166 163.367
R557 B.n221 B.n219 163.367
R558 B.n217 B.n168 163.367
R559 B.n213 B.n211 163.367
R560 B.n209 B.n170 163.367
R561 B.n205 B.n203 163.367
R562 B.n201 B.n172 163.367
R563 B.n197 B.n195 163.367
R564 B.n193 B.n174 163.367
R565 B.n189 B.n187 163.367
R566 B.n185 B.n176 163.367
R567 B.n181 B.n179 163.367
R568 B.n339 B.n126 163.367
R569 B.n347 B.n126 163.367
R570 B.n347 B.n124 163.367
R571 B.n351 B.n124 163.367
R572 B.n351 B.n118 163.367
R573 B.n359 B.n118 163.367
R574 B.n359 B.n116 163.367
R575 B.n363 B.n116 163.367
R576 B.n363 B.n110 163.367
R577 B.n371 B.n110 163.367
R578 B.n371 B.n108 163.367
R579 B.n375 B.n108 163.367
R580 B.n375 B.n102 163.367
R581 B.n383 B.n102 163.367
R582 B.n383 B.n100 163.367
R583 B.n387 B.n100 163.367
R584 B.n387 B.n94 163.367
R585 B.n396 B.n94 163.367
R586 B.n396 B.n92 163.367
R587 B.n400 B.n92 163.367
R588 B.n400 B.n3 163.367
R589 B.n645 B.n3 163.367
R590 B.n641 B.n2 163.367
R591 B.n641 B.n640 163.367
R592 B.n640 B.n9 163.367
R593 B.n636 B.n9 163.367
R594 B.n636 B.n11 163.367
R595 B.n632 B.n11 163.367
R596 B.n632 B.n16 163.367
R597 B.n628 B.n16 163.367
R598 B.n628 B.n18 163.367
R599 B.n624 B.n18 163.367
R600 B.n624 B.n23 163.367
R601 B.n620 B.n23 163.367
R602 B.n620 B.n25 163.367
R603 B.n616 B.n25 163.367
R604 B.n616 B.n30 163.367
R605 B.n612 B.n30 163.367
R606 B.n612 B.n32 163.367
R607 B.n608 B.n32 163.367
R608 B.n608 B.n37 163.367
R609 B.n604 B.n37 163.367
R610 B.n604 B.n39 163.367
R611 B.n600 B.n39 163.367
R612 B.n340 B.n131 84.311
R613 B.n601 B.n43 84.311
R614 B.n595 B.n44 71.676
R615 B.n594 B.n593 71.676
R616 B.n587 B.n46 71.676
R617 B.n586 B.n585 71.676
R618 B.n579 B.n48 71.676
R619 B.n578 B.n577 71.676
R620 B.n571 B.n50 71.676
R621 B.n570 B.n569 71.676
R622 B.n563 B.n52 71.676
R623 B.n562 B.n561 71.676
R624 B.n555 B.n54 71.676
R625 B.n554 B.n553 71.676
R626 B.n547 B.n56 71.676
R627 B.n546 B.n545 71.676
R628 B.n539 B.n58 71.676
R629 B.n538 B.n537 71.676
R630 B.n531 B.n60 71.676
R631 B.n530 B.n529 71.676
R632 B.n522 B.n62 71.676
R633 B.n521 B.n520 71.676
R634 B.n514 B.n66 71.676
R635 B.n513 B.n512 71.676
R636 B.n505 B.n68 71.676
R637 B.n504 B.n503 71.676
R638 B.n497 B.n72 71.676
R639 B.n496 B.n495 71.676
R640 B.n489 B.n74 71.676
R641 B.n488 B.n487 71.676
R642 B.n481 B.n76 71.676
R643 B.n480 B.n479 71.676
R644 B.n473 B.n78 71.676
R645 B.n472 B.n471 71.676
R646 B.n465 B.n80 71.676
R647 B.n464 B.n463 71.676
R648 B.n457 B.n82 71.676
R649 B.n456 B.n455 71.676
R650 B.n449 B.n84 71.676
R651 B.n448 B.n447 71.676
R652 B.n441 B.n86 71.676
R653 B.n440 B.n439 71.676
R654 B.n439 B.n438 71.676
R655 B.n442 B.n441 71.676
R656 B.n447 B.n446 71.676
R657 B.n450 B.n449 71.676
R658 B.n455 B.n454 71.676
R659 B.n458 B.n457 71.676
R660 B.n463 B.n462 71.676
R661 B.n466 B.n465 71.676
R662 B.n471 B.n470 71.676
R663 B.n474 B.n473 71.676
R664 B.n479 B.n478 71.676
R665 B.n482 B.n481 71.676
R666 B.n487 B.n486 71.676
R667 B.n490 B.n489 71.676
R668 B.n495 B.n494 71.676
R669 B.n498 B.n497 71.676
R670 B.n503 B.n502 71.676
R671 B.n506 B.n505 71.676
R672 B.n512 B.n511 71.676
R673 B.n515 B.n514 71.676
R674 B.n520 B.n519 71.676
R675 B.n523 B.n522 71.676
R676 B.n529 B.n528 71.676
R677 B.n532 B.n531 71.676
R678 B.n537 B.n536 71.676
R679 B.n540 B.n539 71.676
R680 B.n545 B.n544 71.676
R681 B.n548 B.n547 71.676
R682 B.n553 B.n552 71.676
R683 B.n556 B.n555 71.676
R684 B.n561 B.n560 71.676
R685 B.n564 B.n563 71.676
R686 B.n569 B.n568 71.676
R687 B.n572 B.n571 71.676
R688 B.n577 B.n576 71.676
R689 B.n580 B.n579 71.676
R690 B.n585 B.n584 71.676
R691 B.n588 B.n587 71.676
R692 B.n593 B.n592 71.676
R693 B.n596 B.n595 71.676
R694 B.n334 B.n132 71.676
R695 B.n332 B.n134 71.676
R696 B.n328 B.n327 71.676
R697 B.n321 B.n136 71.676
R698 B.n320 B.n319 71.676
R699 B.n313 B.n138 71.676
R700 B.n312 B.n311 71.676
R701 B.n305 B.n140 71.676
R702 B.n304 B.n303 71.676
R703 B.n297 B.n142 71.676
R704 B.n296 B.n295 71.676
R705 B.n289 B.n144 71.676
R706 B.n288 B.n287 71.676
R707 B.n281 B.n146 71.676
R708 B.n280 B.n279 71.676
R709 B.n273 B.n148 71.676
R710 B.n272 B.n271 71.676
R711 B.n264 B.n150 71.676
R712 B.n263 B.n262 71.676
R713 B.n256 B.n154 71.676
R714 B.n255 B.n254 71.676
R715 B.n248 B.n156 71.676
R716 B.n247 B.n160 71.676
R717 B.n243 B.n242 71.676
R718 B.n236 B.n162 71.676
R719 B.n235 B.n234 71.676
R720 B.n228 B.n164 71.676
R721 B.n227 B.n226 71.676
R722 B.n220 B.n166 71.676
R723 B.n219 B.n218 71.676
R724 B.n212 B.n168 71.676
R725 B.n211 B.n210 71.676
R726 B.n204 B.n170 71.676
R727 B.n203 B.n202 71.676
R728 B.n196 B.n172 71.676
R729 B.n195 B.n194 71.676
R730 B.n188 B.n174 71.676
R731 B.n187 B.n186 71.676
R732 B.n180 B.n176 71.676
R733 B.n179 B.n178 71.676
R734 B.n335 B.n334 71.676
R735 B.n329 B.n134 71.676
R736 B.n327 B.n326 71.676
R737 B.n322 B.n321 71.676
R738 B.n319 B.n318 71.676
R739 B.n314 B.n313 71.676
R740 B.n311 B.n310 71.676
R741 B.n306 B.n305 71.676
R742 B.n303 B.n302 71.676
R743 B.n298 B.n297 71.676
R744 B.n295 B.n294 71.676
R745 B.n290 B.n289 71.676
R746 B.n287 B.n286 71.676
R747 B.n282 B.n281 71.676
R748 B.n279 B.n278 71.676
R749 B.n274 B.n273 71.676
R750 B.n271 B.n270 71.676
R751 B.n265 B.n264 71.676
R752 B.n262 B.n261 71.676
R753 B.n257 B.n256 71.676
R754 B.n254 B.n253 71.676
R755 B.n249 B.n248 71.676
R756 B.n244 B.n160 71.676
R757 B.n242 B.n241 71.676
R758 B.n237 B.n236 71.676
R759 B.n234 B.n233 71.676
R760 B.n229 B.n228 71.676
R761 B.n226 B.n225 71.676
R762 B.n221 B.n220 71.676
R763 B.n218 B.n217 71.676
R764 B.n213 B.n212 71.676
R765 B.n210 B.n209 71.676
R766 B.n205 B.n204 71.676
R767 B.n202 B.n201 71.676
R768 B.n197 B.n196 71.676
R769 B.n194 B.n193 71.676
R770 B.n189 B.n188 71.676
R771 B.n186 B.n185 71.676
R772 B.n181 B.n180 71.676
R773 B.n178 B.n130 71.676
R774 B.n646 B.n645 71.676
R775 B.n646 B.n2 71.676
R776 B.n526 B.n64 59.5399
R777 B.n508 B.n70 59.5399
R778 B.n159 B.n158 59.5399
R779 B.n267 B.n152 59.5399
R780 B.n340 B.n127 49.0015
R781 B.n346 B.n127 49.0015
R782 B.n346 B.n122 49.0015
R783 B.n352 B.n122 49.0015
R784 B.n352 B.n123 49.0015
R785 B.n358 B.n115 49.0015
R786 B.n364 B.n115 49.0015
R787 B.n364 B.n111 49.0015
R788 B.n370 B.n111 49.0015
R789 B.n370 B.n106 49.0015
R790 B.n376 B.n106 49.0015
R791 B.n376 B.n107 49.0015
R792 B.n382 B.n99 49.0015
R793 B.n388 B.n99 49.0015
R794 B.n388 B.n95 49.0015
R795 B.n395 B.n95 49.0015
R796 B.n401 B.n91 49.0015
R797 B.n401 B.n4 49.0015
R798 B.n644 B.n4 49.0015
R799 B.n644 B.n643 49.0015
R800 B.n643 B.n642 49.0015
R801 B.n642 B.n8 49.0015
R802 B.n410 B.n8 49.0015
R803 B.n635 B.n634 49.0015
R804 B.n634 B.n633 49.0015
R805 B.n633 B.n15 49.0015
R806 B.n627 B.n15 49.0015
R807 B.n626 B.n625 49.0015
R808 B.n625 B.n22 49.0015
R809 B.n619 B.n22 49.0015
R810 B.n619 B.n618 49.0015
R811 B.n618 B.n617 49.0015
R812 B.n617 B.n29 49.0015
R813 B.n611 B.n29 49.0015
R814 B.n610 B.n609 49.0015
R815 B.n609 B.n36 49.0015
R816 B.n603 B.n36 49.0015
R817 B.n603 B.n602 49.0015
R818 B.n602 B.n601 49.0015
R819 B.n123 B.t5 38.1924
R820 B.t9 B.n610 38.1924
R821 B.n107 B.t1 36.7512
R822 B.t2 B.n626 36.7512
R823 B.n64 B.n63 31.4187
R824 B.n70 B.n69 31.4187
R825 B.n158 B.n157 31.4187
R826 B.n152 B.n151 31.4187
R827 B.n338 B.n337 31.3761
R828 B.n342 B.n129 31.3761
R829 B.n436 B.n435 31.3761
R830 B.n599 B.n598 31.3761
R831 B.n395 B.t0 25.2216
R832 B.n635 B.t3 25.2216
R833 B.t0 B.n91 23.7804
R834 B.n410 B.t3 23.7804
R835 B B.n647 18.0485
R836 B.n382 B.t1 12.2507
R837 B.n627 B.t2 12.2507
R838 B.n358 B.t5 10.8095
R839 B.n611 B.t9 10.8095
R840 B.n338 B.n125 10.6151
R841 B.n348 B.n125 10.6151
R842 B.n349 B.n348 10.6151
R843 B.n350 B.n349 10.6151
R844 B.n350 B.n117 10.6151
R845 B.n360 B.n117 10.6151
R846 B.n361 B.n360 10.6151
R847 B.n362 B.n361 10.6151
R848 B.n362 B.n109 10.6151
R849 B.n372 B.n109 10.6151
R850 B.n373 B.n372 10.6151
R851 B.n374 B.n373 10.6151
R852 B.n374 B.n101 10.6151
R853 B.n384 B.n101 10.6151
R854 B.n385 B.n384 10.6151
R855 B.n386 B.n385 10.6151
R856 B.n386 B.n93 10.6151
R857 B.n397 B.n93 10.6151
R858 B.n398 B.n397 10.6151
R859 B.n399 B.n398 10.6151
R860 B.n399 B.n0 10.6151
R861 B.n337 B.n336 10.6151
R862 B.n336 B.n133 10.6151
R863 B.n331 B.n133 10.6151
R864 B.n331 B.n330 10.6151
R865 B.n330 B.n135 10.6151
R866 B.n325 B.n135 10.6151
R867 B.n325 B.n324 10.6151
R868 B.n324 B.n323 10.6151
R869 B.n323 B.n137 10.6151
R870 B.n317 B.n137 10.6151
R871 B.n317 B.n316 10.6151
R872 B.n316 B.n315 10.6151
R873 B.n315 B.n139 10.6151
R874 B.n309 B.n139 10.6151
R875 B.n309 B.n308 10.6151
R876 B.n308 B.n307 10.6151
R877 B.n307 B.n141 10.6151
R878 B.n301 B.n141 10.6151
R879 B.n301 B.n300 10.6151
R880 B.n300 B.n299 10.6151
R881 B.n299 B.n143 10.6151
R882 B.n293 B.n143 10.6151
R883 B.n293 B.n292 10.6151
R884 B.n292 B.n291 10.6151
R885 B.n291 B.n145 10.6151
R886 B.n285 B.n145 10.6151
R887 B.n285 B.n284 10.6151
R888 B.n284 B.n283 10.6151
R889 B.n283 B.n147 10.6151
R890 B.n277 B.n147 10.6151
R891 B.n277 B.n276 10.6151
R892 B.n276 B.n275 10.6151
R893 B.n275 B.n149 10.6151
R894 B.n269 B.n149 10.6151
R895 B.n269 B.n268 10.6151
R896 B.n266 B.n153 10.6151
R897 B.n260 B.n153 10.6151
R898 B.n260 B.n259 10.6151
R899 B.n259 B.n258 10.6151
R900 B.n258 B.n155 10.6151
R901 B.n252 B.n155 10.6151
R902 B.n252 B.n251 10.6151
R903 B.n251 B.n250 10.6151
R904 B.n246 B.n245 10.6151
R905 B.n245 B.n161 10.6151
R906 B.n240 B.n161 10.6151
R907 B.n240 B.n239 10.6151
R908 B.n239 B.n238 10.6151
R909 B.n238 B.n163 10.6151
R910 B.n232 B.n163 10.6151
R911 B.n232 B.n231 10.6151
R912 B.n231 B.n230 10.6151
R913 B.n230 B.n165 10.6151
R914 B.n224 B.n165 10.6151
R915 B.n224 B.n223 10.6151
R916 B.n223 B.n222 10.6151
R917 B.n222 B.n167 10.6151
R918 B.n216 B.n167 10.6151
R919 B.n216 B.n215 10.6151
R920 B.n215 B.n214 10.6151
R921 B.n214 B.n169 10.6151
R922 B.n208 B.n169 10.6151
R923 B.n208 B.n207 10.6151
R924 B.n207 B.n206 10.6151
R925 B.n206 B.n171 10.6151
R926 B.n200 B.n171 10.6151
R927 B.n200 B.n199 10.6151
R928 B.n199 B.n198 10.6151
R929 B.n198 B.n173 10.6151
R930 B.n192 B.n173 10.6151
R931 B.n192 B.n191 10.6151
R932 B.n191 B.n190 10.6151
R933 B.n190 B.n175 10.6151
R934 B.n184 B.n175 10.6151
R935 B.n184 B.n183 10.6151
R936 B.n183 B.n182 10.6151
R937 B.n182 B.n177 10.6151
R938 B.n177 B.n129 10.6151
R939 B.n343 B.n342 10.6151
R940 B.n344 B.n343 10.6151
R941 B.n344 B.n120 10.6151
R942 B.n354 B.n120 10.6151
R943 B.n355 B.n354 10.6151
R944 B.n356 B.n355 10.6151
R945 B.n356 B.n113 10.6151
R946 B.n366 B.n113 10.6151
R947 B.n367 B.n366 10.6151
R948 B.n368 B.n367 10.6151
R949 B.n368 B.n104 10.6151
R950 B.n378 B.n104 10.6151
R951 B.n379 B.n378 10.6151
R952 B.n380 B.n379 10.6151
R953 B.n380 B.n97 10.6151
R954 B.n390 B.n97 10.6151
R955 B.n391 B.n390 10.6151
R956 B.n393 B.n391 10.6151
R957 B.n393 B.n392 10.6151
R958 B.n392 B.n89 10.6151
R959 B.n404 B.n89 10.6151
R960 B.n405 B.n404 10.6151
R961 B.n406 B.n405 10.6151
R962 B.n407 B.n406 10.6151
R963 B.n408 B.n407 10.6151
R964 B.n412 B.n408 10.6151
R965 B.n413 B.n412 10.6151
R966 B.n414 B.n413 10.6151
R967 B.n415 B.n414 10.6151
R968 B.n417 B.n415 10.6151
R969 B.n418 B.n417 10.6151
R970 B.n419 B.n418 10.6151
R971 B.n420 B.n419 10.6151
R972 B.n422 B.n420 10.6151
R973 B.n423 B.n422 10.6151
R974 B.n424 B.n423 10.6151
R975 B.n425 B.n424 10.6151
R976 B.n427 B.n425 10.6151
R977 B.n428 B.n427 10.6151
R978 B.n429 B.n428 10.6151
R979 B.n430 B.n429 10.6151
R980 B.n432 B.n430 10.6151
R981 B.n433 B.n432 10.6151
R982 B.n434 B.n433 10.6151
R983 B.n435 B.n434 10.6151
R984 B.n639 B.n1 10.6151
R985 B.n639 B.n638 10.6151
R986 B.n638 B.n637 10.6151
R987 B.n637 B.n10 10.6151
R988 B.n631 B.n10 10.6151
R989 B.n631 B.n630 10.6151
R990 B.n630 B.n629 10.6151
R991 B.n629 B.n17 10.6151
R992 B.n623 B.n17 10.6151
R993 B.n623 B.n622 10.6151
R994 B.n622 B.n621 10.6151
R995 B.n621 B.n24 10.6151
R996 B.n615 B.n24 10.6151
R997 B.n615 B.n614 10.6151
R998 B.n614 B.n613 10.6151
R999 B.n613 B.n31 10.6151
R1000 B.n607 B.n31 10.6151
R1001 B.n607 B.n606 10.6151
R1002 B.n606 B.n605 10.6151
R1003 B.n605 B.n38 10.6151
R1004 B.n599 B.n38 10.6151
R1005 B.n598 B.n597 10.6151
R1006 B.n597 B.n45 10.6151
R1007 B.n591 B.n45 10.6151
R1008 B.n591 B.n590 10.6151
R1009 B.n590 B.n589 10.6151
R1010 B.n589 B.n47 10.6151
R1011 B.n583 B.n47 10.6151
R1012 B.n583 B.n582 10.6151
R1013 B.n582 B.n581 10.6151
R1014 B.n581 B.n49 10.6151
R1015 B.n575 B.n49 10.6151
R1016 B.n575 B.n574 10.6151
R1017 B.n574 B.n573 10.6151
R1018 B.n573 B.n51 10.6151
R1019 B.n567 B.n51 10.6151
R1020 B.n567 B.n566 10.6151
R1021 B.n566 B.n565 10.6151
R1022 B.n565 B.n53 10.6151
R1023 B.n559 B.n53 10.6151
R1024 B.n559 B.n558 10.6151
R1025 B.n558 B.n557 10.6151
R1026 B.n557 B.n55 10.6151
R1027 B.n551 B.n55 10.6151
R1028 B.n551 B.n550 10.6151
R1029 B.n550 B.n549 10.6151
R1030 B.n549 B.n57 10.6151
R1031 B.n543 B.n57 10.6151
R1032 B.n543 B.n542 10.6151
R1033 B.n542 B.n541 10.6151
R1034 B.n541 B.n59 10.6151
R1035 B.n535 B.n59 10.6151
R1036 B.n535 B.n534 10.6151
R1037 B.n534 B.n533 10.6151
R1038 B.n533 B.n61 10.6151
R1039 B.n527 B.n61 10.6151
R1040 B.n525 B.n524 10.6151
R1041 B.n524 B.n65 10.6151
R1042 B.n518 B.n65 10.6151
R1043 B.n518 B.n517 10.6151
R1044 B.n517 B.n516 10.6151
R1045 B.n516 B.n67 10.6151
R1046 B.n510 B.n67 10.6151
R1047 B.n510 B.n509 10.6151
R1048 B.n507 B.n71 10.6151
R1049 B.n501 B.n71 10.6151
R1050 B.n501 B.n500 10.6151
R1051 B.n500 B.n499 10.6151
R1052 B.n499 B.n73 10.6151
R1053 B.n493 B.n73 10.6151
R1054 B.n493 B.n492 10.6151
R1055 B.n492 B.n491 10.6151
R1056 B.n491 B.n75 10.6151
R1057 B.n485 B.n75 10.6151
R1058 B.n485 B.n484 10.6151
R1059 B.n484 B.n483 10.6151
R1060 B.n483 B.n77 10.6151
R1061 B.n477 B.n77 10.6151
R1062 B.n477 B.n476 10.6151
R1063 B.n476 B.n475 10.6151
R1064 B.n475 B.n79 10.6151
R1065 B.n469 B.n79 10.6151
R1066 B.n469 B.n468 10.6151
R1067 B.n468 B.n467 10.6151
R1068 B.n467 B.n81 10.6151
R1069 B.n461 B.n81 10.6151
R1070 B.n461 B.n460 10.6151
R1071 B.n460 B.n459 10.6151
R1072 B.n459 B.n83 10.6151
R1073 B.n453 B.n83 10.6151
R1074 B.n453 B.n452 10.6151
R1075 B.n452 B.n451 10.6151
R1076 B.n451 B.n85 10.6151
R1077 B.n445 B.n85 10.6151
R1078 B.n445 B.n444 10.6151
R1079 B.n444 B.n443 10.6151
R1080 B.n443 B.n87 10.6151
R1081 B.n437 B.n87 10.6151
R1082 B.n437 B.n436 10.6151
R1083 B.n647 B.n0 8.11757
R1084 B.n647 B.n1 8.11757
R1085 B.n267 B.n266 6.5566
R1086 B.n250 B.n159 6.5566
R1087 B.n526 B.n525 6.5566
R1088 B.n509 B.n508 6.5566
R1089 B.n268 B.n267 4.05904
R1090 B.n246 B.n159 4.05904
R1091 B.n527 B.n526 4.05904
R1092 B.n508 B.n507 4.05904
R1093 VN.n0 VN.t3 223.963
R1094 VN.n1 VN.t1 223.963
R1095 VN.n0 VN.t0 223.738
R1096 VN.n1 VN.t2 223.738
R1097 VN VN.n1 59.1186
R1098 VN VN.n0 18.0466
R1099 VTAIL.n426 VTAIL.n378 289.615
R1100 VTAIL.n48 VTAIL.n0 289.615
R1101 VTAIL.n102 VTAIL.n54 289.615
R1102 VTAIL.n156 VTAIL.n108 289.615
R1103 VTAIL.n372 VTAIL.n324 289.615
R1104 VTAIL.n318 VTAIL.n270 289.615
R1105 VTAIL.n264 VTAIL.n216 289.615
R1106 VTAIL.n210 VTAIL.n162 289.615
R1107 VTAIL.n394 VTAIL.n393 185
R1108 VTAIL.n399 VTAIL.n398 185
R1109 VTAIL.n401 VTAIL.n400 185
R1110 VTAIL.n390 VTAIL.n389 185
R1111 VTAIL.n407 VTAIL.n406 185
R1112 VTAIL.n409 VTAIL.n408 185
R1113 VTAIL.n386 VTAIL.n385 185
R1114 VTAIL.n416 VTAIL.n415 185
R1115 VTAIL.n417 VTAIL.n384 185
R1116 VTAIL.n419 VTAIL.n418 185
R1117 VTAIL.n382 VTAIL.n381 185
R1118 VTAIL.n425 VTAIL.n424 185
R1119 VTAIL.n427 VTAIL.n426 185
R1120 VTAIL.n16 VTAIL.n15 185
R1121 VTAIL.n21 VTAIL.n20 185
R1122 VTAIL.n23 VTAIL.n22 185
R1123 VTAIL.n12 VTAIL.n11 185
R1124 VTAIL.n29 VTAIL.n28 185
R1125 VTAIL.n31 VTAIL.n30 185
R1126 VTAIL.n8 VTAIL.n7 185
R1127 VTAIL.n38 VTAIL.n37 185
R1128 VTAIL.n39 VTAIL.n6 185
R1129 VTAIL.n41 VTAIL.n40 185
R1130 VTAIL.n4 VTAIL.n3 185
R1131 VTAIL.n47 VTAIL.n46 185
R1132 VTAIL.n49 VTAIL.n48 185
R1133 VTAIL.n70 VTAIL.n69 185
R1134 VTAIL.n75 VTAIL.n74 185
R1135 VTAIL.n77 VTAIL.n76 185
R1136 VTAIL.n66 VTAIL.n65 185
R1137 VTAIL.n83 VTAIL.n82 185
R1138 VTAIL.n85 VTAIL.n84 185
R1139 VTAIL.n62 VTAIL.n61 185
R1140 VTAIL.n92 VTAIL.n91 185
R1141 VTAIL.n93 VTAIL.n60 185
R1142 VTAIL.n95 VTAIL.n94 185
R1143 VTAIL.n58 VTAIL.n57 185
R1144 VTAIL.n101 VTAIL.n100 185
R1145 VTAIL.n103 VTAIL.n102 185
R1146 VTAIL.n124 VTAIL.n123 185
R1147 VTAIL.n129 VTAIL.n128 185
R1148 VTAIL.n131 VTAIL.n130 185
R1149 VTAIL.n120 VTAIL.n119 185
R1150 VTAIL.n137 VTAIL.n136 185
R1151 VTAIL.n139 VTAIL.n138 185
R1152 VTAIL.n116 VTAIL.n115 185
R1153 VTAIL.n146 VTAIL.n145 185
R1154 VTAIL.n147 VTAIL.n114 185
R1155 VTAIL.n149 VTAIL.n148 185
R1156 VTAIL.n112 VTAIL.n111 185
R1157 VTAIL.n155 VTAIL.n154 185
R1158 VTAIL.n157 VTAIL.n156 185
R1159 VTAIL.n373 VTAIL.n372 185
R1160 VTAIL.n371 VTAIL.n370 185
R1161 VTAIL.n328 VTAIL.n327 185
R1162 VTAIL.n365 VTAIL.n364 185
R1163 VTAIL.n363 VTAIL.n330 185
R1164 VTAIL.n362 VTAIL.n361 185
R1165 VTAIL.n333 VTAIL.n331 185
R1166 VTAIL.n356 VTAIL.n355 185
R1167 VTAIL.n354 VTAIL.n353 185
R1168 VTAIL.n337 VTAIL.n336 185
R1169 VTAIL.n348 VTAIL.n347 185
R1170 VTAIL.n346 VTAIL.n345 185
R1171 VTAIL.n341 VTAIL.n340 185
R1172 VTAIL.n319 VTAIL.n318 185
R1173 VTAIL.n317 VTAIL.n316 185
R1174 VTAIL.n274 VTAIL.n273 185
R1175 VTAIL.n311 VTAIL.n310 185
R1176 VTAIL.n309 VTAIL.n276 185
R1177 VTAIL.n308 VTAIL.n307 185
R1178 VTAIL.n279 VTAIL.n277 185
R1179 VTAIL.n302 VTAIL.n301 185
R1180 VTAIL.n300 VTAIL.n299 185
R1181 VTAIL.n283 VTAIL.n282 185
R1182 VTAIL.n294 VTAIL.n293 185
R1183 VTAIL.n292 VTAIL.n291 185
R1184 VTAIL.n287 VTAIL.n286 185
R1185 VTAIL.n265 VTAIL.n264 185
R1186 VTAIL.n263 VTAIL.n262 185
R1187 VTAIL.n220 VTAIL.n219 185
R1188 VTAIL.n257 VTAIL.n256 185
R1189 VTAIL.n255 VTAIL.n222 185
R1190 VTAIL.n254 VTAIL.n253 185
R1191 VTAIL.n225 VTAIL.n223 185
R1192 VTAIL.n248 VTAIL.n247 185
R1193 VTAIL.n246 VTAIL.n245 185
R1194 VTAIL.n229 VTAIL.n228 185
R1195 VTAIL.n240 VTAIL.n239 185
R1196 VTAIL.n238 VTAIL.n237 185
R1197 VTAIL.n233 VTAIL.n232 185
R1198 VTAIL.n211 VTAIL.n210 185
R1199 VTAIL.n209 VTAIL.n208 185
R1200 VTAIL.n166 VTAIL.n165 185
R1201 VTAIL.n203 VTAIL.n202 185
R1202 VTAIL.n201 VTAIL.n168 185
R1203 VTAIL.n200 VTAIL.n199 185
R1204 VTAIL.n171 VTAIL.n169 185
R1205 VTAIL.n194 VTAIL.n193 185
R1206 VTAIL.n192 VTAIL.n191 185
R1207 VTAIL.n175 VTAIL.n174 185
R1208 VTAIL.n186 VTAIL.n185 185
R1209 VTAIL.n184 VTAIL.n183 185
R1210 VTAIL.n179 VTAIL.n178 185
R1211 VTAIL.n395 VTAIL.t6 149.524
R1212 VTAIL.n17 VTAIL.t5 149.524
R1213 VTAIL.n71 VTAIL.t0 149.524
R1214 VTAIL.n125 VTAIL.t1 149.524
R1215 VTAIL.n342 VTAIL.t2 149.524
R1216 VTAIL.n288 VTAIL.t3 149.524
R1217 VTAIL.n234 VTAIL.t7 149.524
R1218 VTAIL.n180 VTAIL.t4 149.524
R1219 VTAIL.n399 VTAIL.n393 104.615
R1220 VTAIL.n400 VTAIL.n399 104.615
R1221 VTAIL.n400 VTAIL.n389 104.615
R1222 VTAIL.n407 VTAIL.n389 104.615
R1223 VTAIL.n408 VTAIL.n407 104.615
R1224 VTAIL.n408 VTAIL.n385 104.615
R1225 VTAIL.n416 VTAIL.n385 104.615
R1226 VTAIL.n417 VTAIL.n416 104.615
R1227 VTAIL.n418 VTAIL.n417 104.615
R1228 VTAIL.n418 VTAIL.n381 104.615
R1229 VTAIL.n425 VTAIL.n381 104.615
R1230 VTAIL.n426 VTAIL.n425 104.615
R1231 VTAIL.n21 VTAIL.n15 104.615
R1232 VTAIL.n22 VTAIL.n21 104.615
R1233 VTAIL.n22 VTAIL.n11 104.615
R1234 VTAIL.n29 VTAIL.n11 104.615
R1235 VTAIL.n30 VTAIL.n29 104.615
R1236 VTAIL.n30 VTAIL.n7 104.615
R1237 VTAIL.n38 VTAIL.n7 104.615
R1238 VTAIL.n39 VTAIL.n38 104.615
R1239 VTAIL.n40 VTAIL.n39 104.615
R1240 VTAIL.n40 VTAIL.n3 104.615
R1241 VTAIL.n47 VTAIL.n3 104.615
R1242 VTAIL.n48 VTAIL.n47 104.615
R1243 VTAIL.n75 VTAIL.n69 104.615
R1244 VTAIL.n76 VTAIL.n75 104.615
R1245 VTAIL.n76 VTAIL.n65 104.615
R1246 VTAIL.n83 VTAIL.n65 104.615
R1247 VTAIL.n84 VTAIL.n83 104.615
R1248 VTAIL.n84 VTAIL.n61 104.615
R1249 VTAIL.n92 VTAIL.n61 104.615
R1250 VTAIL.n93 VTAIL.n92 104.615
R1251 VTAIL.n94 VTAIL.n93 104.615
R1252 VTAIL.n94 VTAIL.n57 104.615
R1253 VTAIL.n101 VTAIL.n57 104.615
R1254 VTAIL.n102 VTAIL.n101 104.615
R1255 VTAIL.n129 VTAIL.n123 104.615
R1256 VTAIL.n130 VTAIL.n129 104.615
R1257 VTAIL.n130 VTAIL.n119 104.615
R1258 VTAIL.n137 VTAIL.n119 104.615
R1259 VTAIL.n138 VTAIL.n137 104.615
R1260 VTAIL.n138 VTAIL.n115 104.615
R1261 VTAIL.n146 VTAIL.n115 104.615
R1262 VTAIL.n147 VTAIL.n146 104.615
R1263 VTAIL.n148 VTAIL.n147 104.615
R1264 VTAIL.n148 VTAIL.n111 104.615
R1265 VTAIL.n155 VTAIL.n111 104.615
R1266 VTAIL.n156 VTAIL.n155 104.615
R1267 VTAIL.n372 VTAIL.n371 104.615
R1268 VTAIL.n371 VTAIL.n327 104.615
R1269 VTAIL.n364 VTAIL.n327 104.615
R1270 VTAIL.n364 VTAIL.n363 104.615
R1271 VTAIL.n363 VTAIL.n362 104.615
R1272 VTAIL.n362 VTAIL.n331 104.615
R1273 VTAIL.n355 VTAIL.n331 104.615
R1274 VTAIL.n355 VTAIL.n354 104.615
R1275 VTAIL.n354 VTAIL.n336 104.615
R1276 VTAIL.n347 VTAIL.n336 104.615
R1277 VTAIL.n347 VTAIL.n346 104.615
R1278 VTAIL.n346 VTAIL.n340 104.615
R1279 VTAIL.n318 VTAIL.n317 104.615
R1280 VTAIL.n317 VTAIL.n273 104.615
R1281 VTAIL.n310 VTAIL.n273 104.615
R1282 VTAIL.n310 VTAIL.n309 104.615
R1283 VTAIL.n309 VTAIL.n308 104.615
R1284 VTAIL.n308 VTAIL.n277 104.615
R1285 VTAIL.n301 VTAIL.n277 104.615
R1286 VTAIL.n301 VTAIL.n300 104.615
R1287 VTAIL.n300 VTAIL.n282 104.615
R1288 VTAIL.n293 VTAIL.n282 104.615
R1289 VTAIL.n293 VTAIL.n292 104.615
R1290 VTAIL.n292 VTAIL.n286 104.615
R1291 VTAIL.n264 VTAIL.n263 104.615
R1292 VTAIL.n263 VTAIL.n219 104.615
R1293 VTAIL.n256 VTAIL.n219 104.615
R1294 VTAIL.n256 VTAIL.n255 104.615
R1295 VTAIL.n255 VTAIL.n254 104.615
R1296 VTAIL.n254 VTAIL.n223 104.615
R1297 VTAIL.n247 VTAIL.n223 104.615
R1298 VTAIL.n247 VTAIL.n246 104.615
R1299 VTAIL.n246 VTAIL.n228 104.615
R1300 VTAIL.n239 VTAIL.n228 104.615
R1301 VTAIL.n239 VTAIL.n238 104.615
R1302 VTAIL.n238 VTAIL.n232 104.615
R1303 VTAIL.n210 VTAIL.n209 104.615
R1304 VTAIL.n209 VTAIL.n165 104.615
R1305 VTAIL.n202 VTAIL.n165 104.615
R1306 VTAIL.n202 VTAIL.n201 104.615
R1307 VTAIL.n201 VTAIL.n200 104.615
R1308 VTAIL.n200 VTAIL.n169 104.615
R1309 VTAIL.n193 VTAIL.n169 104.615
R1310 VTAIL.n193 VTAIL.n192 104.615
R1311 VTAIL.n192 VTAIL.n174 104.615
R1312 VTAIL.n185 VTAIL.n174 104.615
R1313 VTAIL.n185 VTAIL.n184 104.615
R1314 VTAIL.n184 VTAIL.n178 104.615
R1315 VTAIL.t6 VTAIL.n393 52.3082
R1316 VTAIL.t5 VTAIL.n15 52.3082
R1317 VTAIL.t0 VTAIL.n69 52.3082
R1318 VTAIL.t1 VTAIL.n123 52.3082
R1319 VTAIL.t2 VTAIL.n340 52.3082
R1320 VTAIL.t3 VTAIL.n286 52.3082
R1321 VTAIL.t7 VTAIL.n232 52.3082
R1322 VTAIL.t4 VTAIL.n178 52.3082
R1323 VTAIL.n431 VTAIL.n430 32.7672
R1324 VTAIL.n53 VTAIL.n52 32.7672
R1325 VTAIL.n107 VTAIL.n106 32.7672
R1326 VTAIL.n161 VTAIL.n160 32.7672
R1327 VTAIL.n377 VTAIL.n376 32.7672
R1328 VTAIL.n323 VTAIL.n322 32.7672
R1329 VTAIL.n269 VTAIL.n268 32.7672
R1330 VTAIL.n215 VTAIL.n214 32.7672
R1331 VTAIL.n431 VTAIL.n377 22.3755
R1332 VTAIL.n215 VTAIL.n161 22.3755
R1333 VTAIL.n419 VTAIL.n384 13.1884
R1334 VTAIL.n41 VTAIL.n6 13.1884
R1335 VTAIL.n95 VTAIL.n60 13.1884
R1336 VTAIL.n149 VTAIL.n114 13.1884
R1337 VTAIL.n365 VTAIL.n330 13.1884
R1338 VTAIL.n311 VTAIL.n276 13.1884
R1339 VTAIL.n257 VTAIL.n222 13.1884
R1340 VTAIL.n203 VTAIL.n168 13.1884
R1341 VTAIL.n415 VTAIL.n414 12.8005
R1342 VTAIL.n420 VTAIL.n382 12.8005
R1343 VTAIL.n37 VTAIL.n36 12.8005
R1344 VTAIL.n42 VTAIL.n4 12.8005
R1345 VTAIL.n91 VTAIL.n90 12.8005
R1346 VTAIL.n96 VTAIL.n58 12.8005
R1347 VTAIL.n145 VTAIL.n144 12.8005
R1348 VTAIL.n150 VTAIL.n112 12.8005
R1349 VTAIL.n366 VTAIL.n328 12.8005
R1350 VTAIL.n361 VTAIL.n332 12.8005
R1351 VTAIL.n312 VTAIL.n274 12.8005
R1352 VTAIL.n307 VTAIL.n278 12.8005
R1353 VTAIL.n258 VTAIL.n220 12.8005
R1354 VTAIL.n253 VTAIL.n224 12.8005
R1355 VTAIL.n204 VTAIL.n166 12.8005
R1356 VTAIL.n199 VTAIL.n170 12.8005
R1357 VTAIL.n413 VTAIL.n386 12.0247
R1358 VTAIL.n424 VTAIL.n423 12.0247
R1359 VTAIL.n35 VTAIL.n8 12.0247
R1360 VTAIL.n46 VTAIL.n45 12.0247
R1361 VTAIL.n89 VTAIL.n62 12.0247
R1362 VTAIL.n100 VTAIL.n99 12.0247
R1363 VTAIL.n143 VTAIL.n116 12.0247
R1364 VTAIL.n154 VTAIL.n153 12.0247
R1365 VTAIL.n370 VTAIL.n369 12.0247
R1366 VTAIL.n360 VTAIL.n333 12.0247
R1367 VTAIL.n316 VTAIL.n315 12.0247
R1368 VTAIL.n306 VTAIL.n279 12.0247
R1369 VTAIL.n262 VTAIL.n261 12.0247
R1370 VTAIL.n252 VTAIL.n225 12.0247
R1371 VTAIL.n208 VTAIL.n207 12.0247
R1372 VTAIL.n198 VTAIL.n171 12.0247
R1373 VTAIL.n410 VTAIL.n409 11.249
R1374 VTAIL.n427 VTAIL.n380 11.249
R1375 VTAIL.n32 VTAIL.n31 11.249
R1376 VTAIL.n49 VTAIL.n2 11.249
R1377 VTAIL.n86 VTAIL.n85 11.249
R1378 VTAIL.n103 VTAIL.n56 11.249
R1379 VTAIL.n140 VTAIL.n139 11.249
R1380 VTAIL.n157 VTAIL.n110 11.249
R1381 VTAIL.n373 VTAIL.n326 11.249
R1382 VTAIL.n357 VTAIL.n356 11.249
R1383 VTAIL.n319 VTAIL.n272 11.249
R1384 VTAIL.n303 VTAIL.n302 11.249
R1385 VTAIL.n265 VTAIL.n218 11.249
R1386 VTAIL.n249 VTAIL.n248 11.249
R1387 VTAIL.n211 VTAIL.n164 11.249
R1388 VTAIL.n195 VTAIL.n194 11.249
R1389 VTAIL.n406 VTAIL.n388 10.4732
R1390 VTAIL.n428 VTAIL.n378 10.4732
R1391 VTAIL.n28 VTAIL.n10 10.4732
R1392 VTAIL.n50 VTAIL.n0 10.4732
R1393 VTAIL.n82 VTAIL.n64 10.4732
R1394 VTAIL.n104 VTAIL.n54 10.4732
R1395 VTAIL.n136 VTAIL.n118 10.4732
R1396 VTAIL.n158 VTAIL.n108 10.4732
R1397 VTAIL.n374 VTAIL.n324 10.4732
R1398 VTAIL.n353 VTAIL.n335 10.4732
R1399 VTAIL.n320 VTAIL.n270 10.4732
R1400 VTAIL.n299 VTAIL.n281 10.4732
R1401 VTAIL.n266 VTAIL.n216 10.4732
R1402 VTAIL.n245 VTAIL.n227 10.4732
R1403 VTAIL.n212 VTAIL.n162 10.4732
R1404 VTAIL.n191 VTAIL.n173 10.4732
R1405 VTAIL.n395 VTAIL.n394 10.2747
R1406 VTAIL.n17 VTAIL.n16 10.2747
R1407 VTAIL.n71 VTAIL.n70 10.2747
R1408 VTAIL.n125 VTAIL.n124 10.2747
R1409 VTAIL.n342 VTAIL.n341 10.2747
R1410 VTAIL.n288 VTAIL.n287 10.2747
R1411 VTAIL.n234 VTAIL.n233 10.2747
R1412 VTAIL.n180 VTAIL.n179 10.2747
R1413 VTAIL.n405 VTAIL.n390 9.69747
R1414 VTAIL.n27 VTAIL.n12 9.69747
R1415 VTAIL.n81 VTAIL.n66 9.69747
R1416 VTAIL.n135 VTAIL.n120 9.69747
R1417 VTAIL.n352 VTAIL.n337 9.69747
R1418 VTAIL.n298 VTAIL.n283 9.69747
R1419 VTAIL.n244 VTAIL.n229 9.69747
R1420 VTAIL.n190 VTAIL.n175 9.69747
R1421 VTAIL.n430 VTAIL.n429 9.45567
R1422 VTAIL.n52 VTAIL.n51 9.45567
R1423 VTAIL.n106 VTAIL.n105 9.45567
R1424 VTAIL.n160 VTAIL.n159 9.45567
R1425 VTAIL.n376 VTAIL.n375 9.45567
R1426 VTAIL.n322 VTAIL.n321 9.45567
R1427 VTAIL.n268 VTAIL.n267 9.45567
R1428 VTAIL.n214 VTAIL.n213 9.45567
R1429 VTAIL.n429 VTAIL.n428 9.3005
R1430 VTAIL.n380 VTAIL.n379 9.3005
R1431 VTAIL.n423 VTAIL.n422 9.3005
R1432 VTAIL.n421 VTAIL.n420 9.3005
R1433 VTAIL.n397 VTAIL.n396 9.3005
R1434 VTAIL.n392 VTAIL.n391 9.3005
R1435 VTAIL.n403 VTAIL.n402 9.3005
R1436 VTAIL.n405 VTAIL.n404 9.3005
R1437 VTAIL.n388 VTAIL.n387 9.3005
R1438 VTAIL.n411 VTAIL.n410 9.3005
R1439 VTAIL.n413 VTAIL.n412 9.3005
R1440 VTAIL.n414 VTAIL.n383 9.3005
R1441 VTAIL.n51 VTAIL.n50 9.3005
R1442 VTAIL.n2 VTAIL.n1 9.3005
R1443 VTAIL.n45 VTAIL.n44 9.3005
R1444 VTAIL.n43 VTAIL.n42 9.3005
R1445 VTAIL.n19 VTAIL.n18 9.3005
R1446 VTAIL.n14 VTAIL.n13 9.3005
R1447 VTAIL.n25 VTAIL.n24 9.3005
R1448 VTAIL.n27 VTAIL.n26 9.3005
R1449 VTAIL.n10 VTAIL.n9 9.3005
R1450 VTAIL.n33 VTAIL.n32 9.3005
R1451 VTAIL.n35 VTAIL.n34 9.3005
R1452 VTAIL.n36 VTAIL.n5 9.3005
R1453 VTAIL.n105 VTAIL.n104 9.3005
R1454 VTAIL.n56 VTAIL.n55 9.3005
R1455 VTAIL.n99 VTAIL.n98 9.3005
R1456 VTAIL.n97 VTAIL.n96 9.3005
R1457 VTAIL.n73 VTAIL.n72 9.3005
R1458 VTAIL.n68 VTAIL.n67 9.3005
R1459 VTAIL.n79 VTAIL.n78 9.3005
R1460 VTAIL.n81 VTAIL.n80 9.3005
R1461 VTAIL.n64 VTAIL.n63 9.3005
R1462 VTAIL.n87 VTAIL.n86 9.3005
R1463 VTAIL.n89 VTAIL.n88 9.3005
R1464 VTAIL.n90 VTAIL.n59 9.3005
R1465 VTAIL.n159 VTAIL.n158 9.3005
R1466 VTAIL.n110 VTAIL.n109 9.3005
R1467 VTAIL.n153 VTAIL.n152 9.3005
R1468 VTAIL.n151 VTAIL.n150 9.3005
R1469 VTAIL.n127 VTAIL.n126 9.3005
R1470 VTAIL.n122 VTAIL.n121 9.3005
R1471 VTAIL.n133 VTAIL.n132 9.3005
R1472 VTAIL.n135 VTAIL.n134 9.3005
R1473 VTAIL.n118 VTAIL.n117 9.3005
R1474 VTAIL.n141 VTAIL.n140 9.3005
R1475 VTAIL.n143 VTAIL.n142 9.3005
R1476 VTAIL.n144 VTAIL.n113 9.3005
R1477 VTAIL.n344 VTAIL.n343 9.3005
R1478 VTAIL.n339 VTAIL.n338 9.3005
R1479 VTAIL.n350 VTAIL.n349 9.3005
R1480 VTAIL.n352 VTAIL.n351 9.3005
R1481 VTAIL.n335 VTAIL.n334 9.3005
R1482 VTAIL.n358 VTAIL.n357 9.3005
R1483 VTAIL.n360 VTAIL.n359 9.3005
R1484 VTAIL.n332 VTAIL.n329 9.3005
R1485 VTAIL.n375 VTAIL.n374 9.3005
R1486 VTAIL.n326 VTAIL.n325 9.3005
R1487 VTAIL.n369 VTAIL.n368 9.3005
R1488 VTAIL.n367 VTAIL.n366 9.3005
R1489 VTAIL.n290 VTAIL.n289 9.3005
R1490 VTAIL.n285 VTAIL.n284 9.3005
R1491 VTAIL.n296 VTAIL.n295 9.3005
R1492 VTAIL.n298 VTAIL.n297 9.3005
R1493 VTAIL.n281 VTAIL.n280 9.3005
R1494 VTAIL.n304 VTAIL.n303 9.3005
R1495 VTAIL.n306 VTAIL.n305 9.3005
R1496 VTAIL.n278 VTAIL.n275 9.3005
R1497 VTAIL.n321 VTAIL.n320 9.3005
R1498 VTAIL.n272 VTAIL.n271 9.3005
R1499 VTAIL.n315 VTAIL.n314 9.3005
R1500 VTAIL.n313 VTAIL.n312 9.3005
R1501 VTAIL.n236 VTAIL.n235 9.3005
R1502 VTAIL.n231 VTAIL.n230 9.3005
R1503 VTAIL.n242 VTAIL.n241 9.3005
R1504 VTAIL.n244 VTAIL.n243 9.3005
R1505 VTAIL.n227 VTAIL.n226 9.3005
R1506 VTAIL.n250 VTAIL.n249 9.3005
R1507 VTAIL.n252 VTAIL.n251 9.3005
R1508 VTAIL.n224 VTAIL.n221 9.3005
R1509 VTAIL.n267 VTAIL.n266 9.3005
R1510 VTAIL.n218 VTAIL.n217 9.3005
R1511 VTAIL.n261 VTAIL.n260 9.3005
R1512 VTAIL.n259 VTAIL.n258 9.3005
R1513 VTAIL.n182 VTAIL.n181 9.3005
R1514 VTAIL.n177 VTAIL.n176 9.3005
R1515 VTAIL.n188 VTAIL.n187 9.3005
R1516 VTAIL.n190 VTAIL.n189 9.3005
R1517 VTAIL.n173 VTAIL.n172 9.3005
R1518 VTAIL.n196 VTAIL.n195 9.3005
R1519 VTAIL.n198 VTAIL.n197 9.3005
R1520 VTAIL.n170 VTAIL.n167 9.3005
R1521 VTAIL.n213 VTAIL.n212 9.3005
R1522 VTAIL.n164 VTAIL.n163 9.3005
R1523 VTAIL.n207 VTAIL.n206 9.3005
R1524 VTAIL.n205 VTAIL.n204 9.3005
R1525 VTAIL.n402 VTAIL.n401 8.92171
R1526 VTAIL.n24 VTAIL.n23 8.92171
R1527 VTAIL.n78 VTAIL.n77 8.92171
R1528 VTAIL.n132 VTAIL.n131 8.92171
R1529 VTAIL.n349 VTAIL.n348 8.92171
R1530 VTAIL.n295 VTAIL.n294 8.92171
R1531 VTAIL.n241 VTAIL.n240 8.92171
R1532 VTAIL.n187 VTAIL.n186 8.92171
R1533 VTAIL.n398 VTAIL.n392 8.14595
R1534 VTAIL.n20 VTAIL.n14 8.14595
R1535 VTAIL.n74 VTAIL.n68 8.14595
R1536 VTAIL.n128 VTAIL.n122 8.14595
R1537 VTAIL.n345 VTAIL.n339 8.14595
R1538 VTAIL.n291 VTAIL.n285 8.14595
R1539 VTAIL.n237 VTAIL.n231 8.14595
R1540 VTAIL.n183 VTAIL.n177 8.14595
R1541 VTAIL.n397 VTAIL.n394 7.3702
R1542 VTAIL.n19 VTAIL.n16 7.3702
R1543 VTAIL.n73 VTAIL.n70 7.3702
R1544 VTAIL.n127 VTAIL.n124 7.3702
R1545 VTAIL.n344 VTAIL.n341 7.3702
R1546 VTAIL.n290 VTAIL.n287 7.3702
R1547 VTAIL.n236 VTAIL.n233 7.3702
R1548 VTAIL.n182 VTAIL.n179 7.3702
R1549 VTAIL.n398 VTAIL.n397 5.81868
R1550 VTAIL.n20 VTAIL.n19 5.81868
R1551 VTAIL.n74 VTAIL.n73 5.81868
R1552 VTAIL.n128 VTAIL.n127 5.81868
R1553 VTAIL.n345 VTAIL.n344 5.81868
R1554 VTAIL.n291 VTAIL.n290 5.81868
R1555 VTAIL.n237 VTAIL.n236 5.81868
R1556 VTAIL.n183 VTAIL.n182 5.81868
R1557 VTAIL.n401 VTAIL.n392 5.04292
R1558 VTAIL.n23 VTAIL.n14 5.04292
R1559 VTAIL.n77 VTAIL.n68 5.04292
R1560 VTAIL.n131 VTAIL.n122 5.04292
R1561 VTAIL.n348 VTAIL.n339 5.04292
R1562 VTAIL.n294 VTAIL.n285 5.04292
R1563 VTAIL.n240 VTAIL.n231 5.04292
R1564 VTAIL.n186 VTAIL.n177 5.04292
R1565 VTAIL.n402 VTAIL.n390 4.26717
R1566 VTAIL.n24 VTAIL.n12 4.26717
R1567 VTAIL.n78 VTAIL.n66 4.26717
R1568 VTAIL.n132 VTAIL.n120 4.26717
R1569 VTAIL.n349 VTAIL.n337 4.26717
R1570 VTAIL.n295 VTAIL.n283 4.26717
R1571 VTAIL.n241 VTAIL.n229 4.26717
R1572 VTAIL.n187 VTAIL.n175 4.26717
R1573 VTAIL.n406 VTAIL.n405 3.49141
R1574 VTAIL.n430 VTAIL.n378 3.49141
R1575 VTAIL.n28 VTAIL.n27 3.49141
R1576 VTAIL.n52 VTAIL.n0 3.49141
R1577 VTAIL.n82 VTAIL.n81 3.49141
R1578 VTAIL.n106 VTAIL.n54 3.49141
R1579 VTAIL.n136 VTAIL.n135 3.49141
R1580 VTAIL.n160 VTAIL.n108 3.49141
R1581 VTAIL.n376 VTAIL.n324 3.49141
R1582 VTAIL.n353 VTAIL.n352 3.49141
R1583 VTAIL.n322 VTAIL.n270 3.49141
R1584 VTAIL.n299 VTAIL.n298 3.49141
R1585 VTAIL.n268 VTAIL.n216 3.49141
R1586 VTAIL.n245 VTAIL.n244 3.49141
R1587 VTAIL.n214 VTAIL.n162 3.49141
R1588 VTAIL.n191 VTAIL.n190 3.49141
R1589 VTAIL.n396 VTAIL.n395 2.84303
R1590 VTAIL.n18 VTAIL.n17 2.84303
R1591 VTAIL.n72 VTAIL.n71 2.84303
R1592 VTAIL.n126 VTAIL.n125 2.84303
R1593 VTAIL.n343 VTAIL.n342 2.84303
R1594 VTAIL.n289 VTAIL.n288 2.84303
R1595 VTAIL.n235 VTAIL.n234 2.84303
R1596 VTAIL.n181 VTAIL.n180 2.84303
R1597 VTAIL.n409 VTAIL.n388 2.71565
R1598 VTAIL.n428 VTAIL.n427 2.71565
R1599 VTAIL.n31 VTAIL.n10 2.71565
R1600 VTAIL.n50 VTAIL.n49 2.71565
R1601 VTAIL.n85 VTAIL.n64 2.71565
R1602 VTAIL.n104 VTAIL.n103 2.71565
R1603 VTAIL.n139 VTAIL.n118 2.71565
R1604 VTAIL.n158 VTAIL.n157 2.71565
R1605 VTAIL.n374 VTAIL.n373 2.71565
R1606 VTAIL.n356 VTAIL.n335 2.71565
R1607 VTAIL.n320 VTAIL.n319 2.71565
R1608 VTAIL.n302 VTAIL.n281 2.71565
R1609 VTAIL.n266 VTAIL.n265 2.71565
R1610 VTAIL.n248 VTAIL.n227 2.71565
R1611 VTAIL.n212 VTAIL.n211 2.71565
R1612 VTAIL.n194 VTAIL.n173 2.71565
R1613 VTAIL.n410 VTAIL.n386 1.93989
R1614 VTAIL.n424 VTAIL.n380 1.93989
R1615 VTAIL.n32 VTAIL.n8 1.93989
R1616 VTAIL.n46 VTAIL.n2 1.93989
R1617 VTAIL.n86 VTAIL.n62 1.93989
R1618 VTAIL.n100 VTAIL.n56 1.93989
R1619 VTAIL.n140 VTAIL.n116 1.93989
R1620 VTAIL.n154 VTAIL.n110 1.93989
R1621 VTAIL.n370 VTAIL.n326 1.93989
R1622 VTAIL.n357 VTAIL.n333 1.93989
R1623 VTAIL.n316 VTAIL.n272 1.93989
R1624 VTAIL.n303 VTAIL.n279 1.93989
R1625 VTAIL.n262 VTAIL.n218 1.93989
R1626 VTAIL.n249 VTAIL.n225 1.93989
R1627 VTAIL.n208 VTAIL.n164 1.93989
R1628 VTAIL.n195 VTAIL.n171 1.93989
R1629 VTAIL.n269 VTAIL.n215 1.39705
R1630 VTAIL.n377 VTAIL.n323 1.39705
R1631 VTAIL.n161 VTAIL.n107 1.39705
R1632 VTAIL.n415 VTAIL.n413 1.16414
R1633 VTAIL.n423 VTAIL.n382 1.16414
R1634 VTAIL.n37 VTAIL.n35 1.16414
R1635 VTAIL.n45 VTAIL.n4 1.16414
R1636 VTAIL.n91 VTAIL.n89 1.16414
R1637 VTAIL.n99 VTAIL.n58 1.16414
R1638 VTAIL.n145 VTAIL.n143 1.16414
R1639 VTAIL.n153 VTAIL.n112 1.16414
R1640 VTAIL.n369 VTAIL.n328 1.16414
R1641 VTAIL.n361 VTAIL.n360 1.16414
R1642 VTAIL.n315 VTAIL.n274 1.16414
R1643 VTAIL.n307 VTAIL.n306 1.16414
R1644 VTAIL.n261 VTAIL.n220 1.16414
R1645 VTAIL.n253 VTAIL.n252 1.16414
R1646 VTAIL.n207 VTAIL.n166 1.16414
R1647 VTAIL.n199 VTAIL.n198 1.16414
R1648 VTAIL VTAIL.n53 0.756965
R1649 VTAIL VTAIL.n431 0.640586
R1650 VTAIL.n323 VTAIL.n269 0.470328
R1651 VTAIL.n107 VTAIL.n53 0.470328
R1652 VTAIL.n414 VTAIL.n384 0.388379
R1653 VTAIL.n420 VTAIL.n419 0.388379
R1654 VTAIL.n36 VTAIL.n6 0.388379
R1655 VTAIL.n42 VTAIL.n41 0.388379
R1656 VTAIL.n90 VTAIL.n60 0.388379
R1657 VTAIL.n96 VTAIL.n95 0.388379
R1658 VTAIL.n144 VTAIL.n114 0.388379
R1659 VTAIL.n150 VTAIL.n149 0.388379
R1660 VTAIL.n366 VTAIL.n365 0.388379
R1661 VTAIL.n332 VTAIL.n330 0.388379
R1662 VTAIL.n312 VTAIL.n311 0.388379
R1663 VTAIL.n278 VTAIL.n276 0.388379
R1664 VTAIL.n258 VTAIL.n257 0.388379
R1665 VTAIL.n224 VTAIL.n222 0.388379
R1666 VTAIL.n204 VTAIL.n203 0.388379
R1667 VTAIL.n170 VTAIL.n168 0.388379
R1668 VTAIL.n396 VTAIL.n391 0.155672
R1669 VTAIL.n403 VTAIL.n391 0.155672
R1670 VTAIL.n404 VTAIL.n403 0.155672
R1671 VTAIL.n404 VTAIL.n387 0.155672
R1672 VTAIL.n411 VTAIL.n387 0.155672
R1673 VTAIL.n412 VTAIL.n411 0.155672
R1674 VTAIL.n412 VTAIL.n383 0.155672
R1675 VTAIL.n421 VTAIL.n383 0.155672
R1676 VTAIL.n422 VTAIL.n421 0.155672
R1677 VTAIL.n422 VTAIL.n379 0.155672
R1678 VTAIL.n429 VTAIL.n379 0.155672
R1679 VTAIL.n18 VTAIL.n13 0.155672
R1680 VTAIL.n25 VTAIL.n13 0.155672
R1681 VTAIL.n26 VTAIL.n25 0.155672
R1682 VTAIL.n26 VTAIL.n9 0.155672
R1683 VTAIL.n33 VTAIL.n9 0.155672
R1684 VTAIL.n34 VTAIL.n33 0.155672
R1685 VTAIL.n34 VTAIL.n5 0.155672
R1686 VTAIL.n43 VTAIL.n5 0.155672
R1687 VTAIL.n44 VTAIL.n43 0.155672
R1688 VTAIL.n44 VTAIL.n1 0.155672
R1689 VTAIL.n51 VTAIL.n1 0.155672
R1690 VTAIL.n72 VTAIL.n67 0.155672
R1691 VTAIL.n79 VTAIL.n67 0.155672
R1692 VTAIL.n80 VTAIL.n79 0.155672
R1693 VTAIL.n80 VTAIL.n63 0.155672
R1694 VTAIL.n87 VTAIL.n63 0.155672
R1695 VTAIL.n88 VTAIL.n87 0.155672
R1696 VTAIL.n88 VTAIL.n59 0.155672
R1697 VTAIL.n97 VTAIL.n59 0.155672
R1698 VTAIL.n98 VTAIL.n97 0.155672
R1699 VTAIL.n98 VTAIL.n55 0.155672
R1700 VTAIL.n105 VTAIL.n55 0.155672
R1701 VTAIL.n126 VTAIL.n121 0.155672
R1702 VTAIL.n133 VTAIL.n121 0.155672
R1703 VTAIL.n134 VTAIL.n133 0.155672
R1704 VTAIL.n134 VTAIL.n117 0.155672
R1705 VTAIL.n141 VTAIL.n117 0.155672
R1706 VTAIL.n142 VTAIL.n141 0.155672
R1707 VTAIL.n142 VTAIL.n113 0.155672
R1708 VTAIL.n151 VTAIL.n113 0.155672
R1709 VTAIL.n152 VTAIL.n151 0.155672
R1710 VTAIL.n152 VTAIL.n109 0.155672
R1711 VTAIL.n159 VTAIL.n109 0.155672
R1712 VTAIL.n375 VTAIL.n325 0.155672
R1713 VTAIL.n368 VTAIL.n325 0.155672
R1714 VTAIL.n368 VTAIL.n367 0.155672
R1715 VTAIL.n367 VTAIL.n329 0.155672
R1716 VTAIL.n359 VTAIL.n329 0.155672
R1717 VTAIL.n359 VTAIL.n358 0.155672
R1718 VTAIL.n358 VTAIL.n334 0.155672
R1719 VTAIL.n351 VTAIL.n334 0.155672
R1720 VTAIL.n351 VTAIL.n350 0.155672
R1721 VTAIL.n350 VTAIL.n338 0.155672
R1722 VTAIL.n343 VTAIL.n338 0.155672
R1723 VTAIL.n321 VTAIL.n271 0.155672
R1724 VTAIL.n314 VTAIL.n271 0.155672
R1725 VTAIL.n314 VTAIL.n313 0.155672
R1726 VTAIL.n313 VTAIL.n275 0.155672
R1727 VTAIL.n305 VTAIL.n275 0.155672
R1728 VTAIL.n305 VTAIL.n304 0.155672
R1729 VTAIL.n304 VTAIL.n280 0.155672
R1730 VTAIL.n297 VTAIL.n280 0.155672
R1731 VTAIL.n297 VTAIL.n296 0.155672
R1732 VTAIL.n296 VTAIL.n284 0.155672
R1733 VTAIL.n289 VTAIL.n284 0.155672
R1734 VTAIL.n267 VTAIL.n217 0.155672
R1735 VTAIL.n260 VTAIL.n217 0.155672
R1736 VTAIL.n260 VTAIL.n259 0.155672
R1737 VTAIL.n259 VTAIL.n221 0.155672
R1738 VTAIL.n251 VTAIL.n221 0.155672
R1739 VTAIL.n251 VTAIL.n250 0.155672
R1740 VTAIL.n250 VTAIL.n226 0.155672
R1741 VTAIL.n243 VTAIL.n226 0.155672
R1742 VTAIL.n243 VTAIL.n242 0.155672
R1743 VTAIL.n242 VTAIL.n230 0.155672
R1744 VTAIL.n235 VTAIL.n230 0.155672
R1745 VTAIL.n213 VTAIL.n163 0.155672
R1746 VTAIL.n206 VTAIL.n163 0.155672
R1747 VTAIL.n206 VTAIL.n205 0.155672
R1748 VTAIL.n205 VTAIL.n167 0.155672
R1749 VTAIL.n197 VTAIL.n167 0.155672
R1750 VTAIL.n197 VTAIL.n196 0.155672
R1751 VTAIL.n196 VTAIL.n172 0.155672
R1752 VTAIL.n189 VTAIL.n172 0.155672
R1753 VTAIL.n189 VTAIL.n188 0.155672
R1754 VTAIL.n188 VTAIL.n176 0.155672
R1755 VTAIL.n181 VTAIL.n176 0.155672
R1756 VDD2.n2 VDD2.n0 99.7385
R1757 VDD2.n2 VDD2.n1 63.222
R1758 VDD2.n1 VDD2.t1 1.98248
R1759 VDD2.n1 VDD2.t2 1.98248
R1760 VDD2.n0 VDD2.t0 1.98248
R1761 VDD2.n0 VDD2.t3 1.98248
R1762 VDD2 VDD2.n2 0.0586897
R1763 VP.n2 VP.t0 223.963
R1764 VP.n2 VP.t3 223.738
R1765 VP.n3 VP.t2 186.636
R1766 VP.n9 VP.t1 186.636
R1767 VP.n4 VP.n3 170.597
R1768 VP.n10 VP.n9 170.597
R1769 VP.n8 VP.n0 161.3
R1770 VP.n7 VP.n6 161.3
R1771 VP.n5 VP.n1 161.3
R1772 VP.n4 VP.n2 58.7379
R1773 VP.n7 VP.n1 40.4934
R1774 VP.n8 VP.n7 40.4934
R1775 VP.n3 VP.n1 15.17
R1776 VP.n9 VP.n8 15.17
R1777 VP.n5 VP.n4 0.189894
R1778 VP.n6 VP.n5 0.189894
R1779 VP.n6 VP.n0 0.189894
R1780 VP.n10 VP.n0 0.189894
R1781 VP VP.n10 0.0516364
R1782 VDD1 VDD1.n1 100.263
R1783 VDD1 VDD1.n0 63.2802
R1784 VDD1.n0 VDD1.t3 1.98248
R1785 VDD1.n0 VDD1.t0 1.98248
R1786 VDD1.n1 VDD1.t1 1.98248
R1787 VDD1.n1 VDD1.t2 1.98248
C0 VP VN 4.87429f
C1 VP VDD1 3.54546f
C2 VDD1 VN 0.14763f
C3 VP VDD2 0.310762f
C4 VDD2 VN 3.38273f
C5 VP VTAIL 3.1826f
C6 VN VTAIL 3.1685f
C7 VDD2 VDD1 0.706218f
C8 VDD1 VTAIL 5.03376f
C9 VDD2 VTAIL 5.07919f
C10 VDD2 B 2.873437f
C11 VDD1 B 6.33964f
C12 VTAIL B 8.071807f
C13 VN B 8.37735f
C14 VP B 6.007477f
C15 VDD1.t3 B 0.210848f
C16 VDD1.t0 B 0.210848f
C17 VDD1.n0 B 1.85726f
C18 VDD1.t1 B 0.210848f
C19 VDD1.t2 B 0.210848f
C20 VDD1.n1 B 2.41081f
C21 VP.n0 B 0.039234f
C22 VP.t1 B 1.36969f
C23 VP.n1 B 0.064259f
C24 VP.t0 B 1.47694f
C25 VP.t3 B 1.47627f
C26 VP.n2 B 2.30491f
C27 VP.t2 B 1.36969f
C28 VP.n3 B 0.58439f
C29 VP.n4 B 2.10223f
C30 VP.n5 B 0.039234f
C31 VP.n6 B 0.039234f
C32 VP.n7 B 0.031717f
C33 VP.n8 B 0.064259f
C34 VP.n9 B 0.58439f
C35 VP.n10 B 0.034784f
C36 VDD2.t0 B 0.213324f
C37 VDD2.t3 B 0.213324f
C38 VDD2.n0 B 2.41406f
C39 VDD2.t1 B 0.213324f
C40 VDD2.t2 B 0.213324f
C41 VDD2.n1 B 1.87873f
C42 VDD2.n2 B 3.22649f
C43 VTAIL.n0 B 0.022013f
C44 VTAIL.n1 B 0.016368f
C45 VTAIL.n2 B 0.008796f
C46 VTAIL.n3 B 0.02079f
C47 VTAIL.n4 B 0.009313f
C48 VTAIL.n5 B 0.016368f
C49 VTAIL.n6 B 0.009054f
C50 VTAIL.n7 B 0.02079f
C51 VTAIL.n8 B 0.009313f
C52 VTAIL.n9 B 0.016368f
C53 VTAIL.n10 B 0.008796f
C54 VTAIL.n11 B 0.02079f
C55 VTAIL.n12 B 0.009313f
C56 VTAIL.n13 B 0.016368f
C57 VTAIL.n14 B 0.008796f
C58 VTAIL.n15 B 0.015592f
C59 VTAIL.n16 B 0.014697f
C60 VTAIL.t5 B 0.034936f
C61 VTAIL.n17 B 0.105385f
C62 VTAIL.n18 B 0.679413f
C63 VTAIL.n19 B 0.008796f
C64 VTAIL.n20 B 0.009313f
C65 VTAIL.n21 B 0.02079f
C66 VTAIL.n22 B 0.02079f
C67 VTAIL.n23 B 0.009313f
C68 VTAIL.n24 B 0.008796f
C69 VTAIL.n25 B 0.016368f
C70 VTAIL.n26 B 0.016368f
C71 VTAIL.n27 B 0.008796f
C72 VTAIL.n28 B 0.009313f
C73 VTAIL.n29 B 0.02079f
C74 VTAIL.n30 B 0.02079f
C75 VTAIL.n31 B 0.009313f
C76 VTAIL.n32 B 0.008796f
C77 VTAIL.n33 B 0.016368f
C78 VTAIL.n34 B 0.016368f
C79 VTAIL.n35 B 0.008796f
C80 VTAIL.n36 B 0.008796f
C81 VTAIL.n37 B 0.009313f
C82 VTAIL.n38 B 0.02079f
C83 VTAIL.n39 B 0.02079f
C84 VTAIL.n40 B 0.02079f
C85 VTAIL.n41 B 0.009054f
C86 VTAIL.n42 B 0.008796f
C87 VTAIL.n43 B 0.016368f
C88 VTAIL.n44 B 0.016368f
C89 VTAIL.n45 B 0.008796f
C90 VTAIL.n46 B 0.009313f
C91 VTAIL.n47 B 0.02079f
C92 VTAIL.n48 B 0.043248f
C93 VTAIL.n49 B 0.009313f
C94 VTAIL.n50 B 0.008796f
C95 VTAIL.n51 B 0.038505f
C96 VTAIL.n52 B 0.024039f
C97 VTAIL.n53 B 0.079036f
C98 VTAIL.n54 B 0.022013f
C99 VTAIL.n55 B 0.016368f
C100 VTAIL.n56 B 0.008796f
C101 VTAIL.n57 B 0.02079f
C102 VTAIL.n58 B 0.009313f
C103 VTAIL.n59 B 0.016368f
C104 VTAIL.n60 B 0.009054f
C105 VTAIL.n61 B 0.02079f
C106 VTAIL.n62 B 0.009313f
C107 VTAIL.n63 B 0.016368f
C108 VTAIL.n64 B 0.008796f
C109 VTAIL.n65 B 0.02079f
C110 VTAIL.n66 B 0.009313f
C111 VTAIL.n67 B 0.016368f
C112 VTAIL.n68 B 0.008796f
C113 VTAIL.n69 B 0.015592f
C114 VTAIL.n70 B 0.014697f
C115 VTAIL.t0 B 0.034936f
C116 VTAIL.n71 B 0.105385f
C117 VTAIL.n72 B 0.679413f
C118 VTAIL.n73 B 0.008796f
C119 VTAIL.n74 B 0.009313f
C120 VTAIL.n75 B 0.02079f
C121 VTAIL.n76 B 0.02079f
C122 VTAIL.n77 B 0.009313f
C123 VTAIL.n78 B 0.008796f
C124 VTAIL.n79 B 0.016368f
C125 VTAIL.n80 B 0.016368f
C126 VTAIL.n81 B 0.008796f
C127 VTAIL.n82 B 0.009313f
C128 VTAIL.n83 B 0.02079f
C129 VTAIL.n84 B 0.02079f
C130 VTAIL.n85 B 0.009313f
C131 VTAIL.n86 B 0.008796f
C132 VTAIL.n87 B 0.016368f
C133 VTAIL.n88 B 0.016368f
C134 VTAIL.n89 B 0.008796f
C135 VTAIL.n90 B 0.008796f
C136 VTAIL.n91 B 0.009313f
C137 VTAIL.n92 B 0.02079f
C138 VTAIL.n93 B 0.02079f
C139 VTAIL.n94 B 0.02079f
C140 VTAIL.n95 B 0.009054f
C141 VTAIL.n96 B 0.008796f
C142 VTAIL.n97 B 0.016368f
C143 VTAIL.n98 B 0.016368f
C144 VTAIL.n99 B 0.008796f
C145 VTAIL.n100 B 0.009313f
C146 VTAIL.n101 B 0.02079f
C147 VTAIL.n102 B 0.043248f
C148 VTAIL.n103 B 0.009313f
C149 VTAIL.n104 B 0.008796f
C150 VTAIL.n105 B 0.038505f
C151 VTAIL.n106 B 0.024039f
C152 VTAIL.n107 B 0.112796f
C153 VTAIL.n108 B 0.022013f
C154 VTAIL.n109 B 0.016368f
C155 VTAIL.n110 B 0.008796f
C156 VTAIL.n111 B 0.02079f
C157 VTAIL.n112 B 0.009313f
C158 VTAIL.n113 B 0.016368f
C159 VTAIL.n114 B 0.009054f
C160 VTAIL.n115 B 0.02079f
C161 VTAIL.n116 B 0.009313f
C162 VTAIL.n117 B 0.016368f
C163 VTAIL.n118 B 0.008796f
C164 VTAIL.n119 B 0.02079f
C165 VTAIL.n120 B 0.009313f
C166 VTAIL.n121 B 0.016368f
C167 VTAIL.n122 B 0.008796f
C168 VTAIL.n123 B 0.015592f
C169 VTAIL.n124 B 0.014697f
C170 VTAIL.t1 B 0.034936f
C171 VTAIL.n125 B 0.105385f
C172 VTAIL.n126 B 0.679413f
C173 VTAIL.n127 B 0.008796f
C174 VTAIL.n128 B 0.009313f
C175 VTAIL.n129 B 0.02079f
C176 VTAIL.n130 B 0.02079f
C177 VTAIL.n131 B 0.009313f
C178 VTAIL.n132 B 0.008796f
C179 VTAIL.n133 B 0.016368f
C180 VTAIL.n134 B 0.016368f
C181 VTAIL.n135 B 0.008796f
C182 VTAIL.n136 B 0.009313f
C183 VTAIL.n137 B 0.02079f
C184 VTAIL.n138 B 0.02079f
C185 VTAIL.n139 B 0.009313f
C186 VTAIL.n140 B 0.008796f
C187 VTAIL.n141 B 0.016368f
C188 VTAIL.n142 B 0.016368f
C189 VTAIL.n143 B 0.008796f
C190 VTAIL.n144 B 0.008796f
C191 VTAIL.n145 B 0.009313f
C192 VTAIL.n146 B 0.02079f
C193 VTAIL.n147 B 0.02079f
C194 VTAIL.n148 B 0.02079f
C195 VTAIL.n149 B 0.009054f
C196 VTAIL.n150 B 0.008796f
C197 VTAIL.n151 B 0.016368f
C198 VTAIL.n152 B 0.016368f
C199 VTAIL.n153 B 0.008796f
C200 VTAIL.n154 B 0.009313f
C201 VTAIL.n155 B 0.02079f
C202 VTAIL.n156 B 0.043248f
C203 VTAIL.n157 B 0.009313f
C204 VTAIL.n158 B 0.008796f
C205 VTAIL.n159 B 0.038505f
C206 VTAIL.n160 B 0.024039f
C207 VTAIL.n161 B 0.838237f
C208 VTAIL.n162 B 0.022013f
C209 VTAIL.n163 B 0.016368f
C210 VTAIL.n164 B 0.008796f
C211 VTAIL.n165 B 0.02079f
C212 VTAIL.n166 B 0.009313f
C213 VTAIL.n167 B 0.016368f
C214 VTAIL.n168 B 0.009054f
C215 VTAIL.n169 B 0.02079f
C216 VTAIL.n170 B 0.008796f
C217 VTAIL.n171 B 0.009313f
C218 VTAIL.n172 B 0.016368f
C219 VTAIL.n173 B 0.008796f
C220 VTAIL.n174 B 0.02079f
C221 VTAIL.n175 B 0.009313f
C222 VTAIL.n176 B 0.016368f
C223 VTAIL.n177 B 0.008796f
C224 VTAIL.n178 B 0.015592f
C225 VTAIL.n179 B 0.014697f
C226 VTAIL.t4 B 0.034936f
C227 VTAIL.n180 B 0.105385f
C228 VTAIL.n181 B 0.679413f
C229 VTAIL.n182 B 0.008796f
C230 VTAIL.n183 B 0.009313f
C231 VTAIL.n184 B 0.02079f
C232 VTAIL.n185 B 0.02079f
C233 VTAIL.n186 B 0.009313f
C234 VTAIL.n187 B 0.008796f
C235 VTAIL.n188 B 0.016368f
C236 VTAIL.n189 B 0.016368f
C237 VTAIL.n190 B 0.008796f
C238 VTAIL.n191 B 0.009313f
C239 VTAIL.n192 B 0.02079f
C240 VTAIL.n193 B 0.02079f
C241 VTAIL.n194 B 0.009313f
C242 VTAIL.n195 B 0.008796f
C243 VTAIL.n196 B 0.016368f
C244 VTAIL.n197 B 0.016368f
C245 VTAIL.n198 B 0.008796f
C246 VTAIL.n199 B 0.009313f
C247 VTAIL.n200 B 0.02079f
C248 VTAIL.n201 B 0.02079f
C249 VTAIL.n202 B 0.02079f
C250 VTAIL.n203 B 0.009054f
C251 VTAIL.n204 B 0.008796f
C252 VTAIL.n205 B 0.016368f
C253 VTAIL.n206 B 0.016368f
C254 VTAIL.n207 B 0.008796f
C255 VTAIL.n208 B 0.009313f
C256 VTAIL.n209 B 0.02079f
C257 VTAIL.n210 B 0.043248f
C258 VTAIL.n211 B 0.009313f
C259 VTAIL.n212 B 0.008796f
C260 VTAIL.n213 B 0.038505f
C261 VTAIL.n214 B 0.024039f
C262 VTAIL.n215 B 0.838237f
C263 VTAIL.n216 B 0.022013f
C264 VTAIL.n217 B 0.016368f
C265 VTAIL.n218 B 0.008796f
C266 VTAIL.n219 B 0.02079f
C267 VTAIL.n220 B 0.009313f
C268 VTAIL.n221 B 0.016368f
C269 VTAIL.n222 B 0.009054f
C270 VTAIL.n223 B 0.02079f
C271 VTAIL.n224 B 0.008796f
C272 VTAIL.n225 B 0.009313f
C273 VTAIL.n226 B 0.016368f
C274 VTAIL.n227 B 0.008796f
C275 VTAIL.n228 B 0.02079f
C276 VTAIL.n229 B 0.009313f
C277 VTAIL.n230 B 0.016368f
C278 VTAIL.n231 B 0.008796f
C279 VTAIL.n232 B 0.015592f
C280 VTAIL.n233 B 0.014697f
C281 VTAIL.t7 B 0.034936f
C282 VTAIL.n234 B 0.105385f
C283 VTAIL.n235 B 0.679413f
C284 VTAIL.n236 B 0.008796f
C285 VTAIL.n237 B 0.009313f
C286 VTAIL.n238 B 0.02079f
C287 VTAIL.n239 B 0.02079f
C288 VTAIL.n240 B 0.009313f
C289 VTAIL.n241 B 0.008796f
C290 VTAIL.n242 B 0.016368f
C291 VTAIL.n243 B 0.016368f
C292 VTAIL.n244 B 0.008796f
C293 VTAIL.n245 B 0.009313f
C294 VTAIL.n246 B 0.02079f
C295 VTAIL.n247 B 0.02079f
C296 VTAIL.n248 B 0.009313f
C297 VTAIL.n249 B 0.008796f
C298 VTAIL.n250 B 0.016368f
C299 VTAIL.n251 B 0.016368f
C300 VTAIL.n252 B 0.008796f
C301 VTAIL.n253 B 0.009313f
C302 VTAIL.n254 B 0.02079f
C303 VTAIL.n255 B 0.02079f
C304 VTAIL.n256 B 0.02079f
C305 VTAIL.n257 B 0.009054f
C306 VTAIL.n258 B 0.008796f
C307 VTAIL.n259 B 0.016368f
C308 VTAIL.n260 B 0.016368f
C309 VTAIL.n261 B 0.008796f
C310 VTAIL.n262 B 0.009313f
C311 VTAIL.n263 B 0.02079f
C312 VTAIL.n264 B 0.043248f
C313 VTAIL.n265 B 0.009313f
C314 VTAIL.n266 B 0.008796f
C315 VTAIL.n267 B 0.038505f
C316 VTAIL.n268 B 0.024039f
C317 VTAIL.n269 B 0.112796f
C318 VTAIL.n270 B 0.022013f
C319 VTAIL.n271 B 0.016368f
C320 VTAIL.n272 B 0.008796f
C321 VTAIL.n273 B 0.02079f
C322 VTAIL.n274 B 0.009313f
C323 VTAIL.n275 B 0.016368f
C324 VTAIL.n276 B 0.009054f
C325 VTAIL.n277 B 0.02079f
C326 VTAIL.n278 B 0.008796f
C327 VTAIL.n279 B 0.009313f
C328 VTAIL.n280 B 0.016368f
C329 VTAIL.n281 B 0.008796f
C330 VTAIL.n282 B 0.02079f
C331 VTAIL.n283 B 0.009313f
C332 VTAIL.n284 B 0.016368f
C333 VTAIL.n285 B 0.008796f
C334 VTAIL.n286 B 0.015592f
C335 VTAIL.n287 B 0.014697f
C336 VTAIL.t3 B 0.034936f
C337 VTAIL.n288 B 0.105385f
C338 VTAIL.n289 B 0.679413f
C339 VTAIL.n290 B 0.008796f
C340 VTAIL.n291 B 0.009313f
C341 VTAIL.n292 B 0.02079f
C342 VTAIL.n293 B 0.02079f
C343 VTAIL.n294 B 0.009313f
C344 VTAIL.n295 B 0.008796f
C345 VTAIL.n296 B 0.016368f
C346 VTAIL.n297 B 0.016368f
C347 VTAIL.n298 B 0.008796f
C348 VTAIL.n299 B 0.009313f
C349 VTAIL.n300 B 0.02079f
C350 VTAIL.n301 B 0.02079f
C351 VTAIL.n302 B 0.009313f
C352 VTAIL.n303 B 0.008796f
C353 VTAIL.n304 B 0.016368f
C354 VTAIL.n305 B 0.016368f
C355 VTAIL.n306 B 0.008796f
C356 VTAIL.n307 B 0.009313f
C357 VTAIL.n308 B 0.02079f
C358 VTAIL.n309 B 0.02079f
C359 VTAIL.n310 B 0.02079f
C360 VTAIL.n311 B 0.009054f
C361 VTAIL.n312 B 0.008796f
C362 VTAIL.n313 B 0.016368f
C363 VTAIL.n314 B 0.016368f
C364 VTAIL.n315 B 0.008796f
C365 VTAIL.n316 B 0.009313f
C366 VTAIL.n317 B 0.02079f
C367 VTAIL.n318 B 0.043248f
C368 VTAIL.n319 B 0.009313f
C369 VTAIL.n320 B 0.008796f
C370 VTAIL.n321 B 0.038505f
C371 VTAIL.n322 B 0.024039f
C372 VTAIL.n323 B 0.112796f
C373 VTAIL.n324 B 0.022013f
C374 VTAIL.n325 B 0.016368f
C375 VTAIL.n326 B 0.008796f
C376 VTAIL.n327 B 0.02079f
C377 VTAIL.n328 B 0.009313f
C378 VTAIL.n329 B 0.016368f
C379 VTAIL.n330 B 0.009054f
C380 VTAIL.n331 B 0.02079f
C381 VTAIL.n332 B 0.008796f
C382 VTAIL.n333 B 0.009313f
C383 VTAIL.n334 B 0.016368f
C384 VTAIL.n335 B 0.008796f
C385 VTAIL.n336 B 0.02079f
C386 VTAIL.n337 B 0.009313f
C387 VTAIL.n338 B 0.016368f
C388 VTAIL.n339 B 0.008796f
C389 VTAIL.n340 B 0.015592f
C390 VTAIL.n341 B 0.014697f
C391 VTAIL.t2 B 0.034936f
C392 VTAIL.n342 B 0.105385f
C393 VTAIL.n343 B 0.679413f
C394 VTAIL.n344 B 0.008796f
C395 VTAIL.n345 B 0.009313f
C396 VTAIL.n346 B 0.02079f
C397 VTAIL.n347 B 0.02079f
C398 VTAIL.n348 B 0.009313f
C399 VTAIL.n349 B 0.008796f
C400 VTAIL.n350 B 0.016368f
C401 VTAIL.n351 B 0.016368f
C402 VTAIL.n352 B 0.008796f
C403 VTAIL.n353 B 0.009313f
C404 VTAIL.n354 B 0.02079f
C405 VTAIL.n355 B 0.02079f
C406 VTAIL.n356 B 0.009313f
C407 VTAIL.n357 B 0.008796f
C408 VTAIL.n358 B 0.016368f
C409 VTAIL.n359 B 0.016368f
C410 VTAIL.n360 B 0.008796f
C411 VTAIL.n361 B 0.009313f
C412 VTAIL.n362 B 0.02079f
C413 VTAIL.n363 B 0.02079f
C414 VTAIL.n364 B 0.02079f
C415 VTAIL.n365 B 0.009054f
C416 VTAIL.n366 B 0.008796f
C417 VTAIL.n367 B 0.016368f
C418 VTAIL.n368 B 0.016368f
C419 VTAIL.n369 B 0.008796f
C420 VTAIL.n370 B 0.009313f
C421 VTAIL.n371 B 0.02079f
C422 VTAIL.n372 B 0.043248f
C423 VTAIL.n373 B 0.009313f
C424 VTAIL.n374 B 0.008796f
C425 VTAIL.n375 B 0.038505f
C426 VTAIL.n376 B 0.024039f
C427 VTAIL.n377 B 0.838237f
C428 VTAIL.n378 B 0.022013f
C429 VTAIL.n379 B 0.016368f
C430 VTAIL.n380 B 0.008796f
C431 VTAIL.n381 B 0.02079f
C432 VTAIL.n382 B 0.009313f
C433 VTAIL.n383 B 0.016368f
C434 VTAIL.n384 B 0.009054f
C435 VTAIL.n385 B 0.02079f
C436 VTAIL.n386 B 0.009313f
C437 VTAIL.n387 B 0.016368f
C438 VTAIL.n388 B 0.008796f
C439 VTAIL.n389 B 0.02079f
C440 VTAIL.n390 B 0.009313f
C441 VTAIL.n391 B 0.016368f
C442 VTAIL.n392 B 0.008796f
C443 VTAIL.n393 B 0.015592f
C444 VTAIL.n394 B 0.014697f
C445 VTAIL.t6 B 0.034936f
C446 VTAIL.n395 B 0.105385f
C447 VTAIL.n396 B 0.679413f
C448 VTAIL.n397 B 0.008796f
C449 VTAIL.n398 B 0.009313f
C450 VTAIL.n399 B 0.02079f
C451 VTAIL.n400 B 0.02079f
C452 VTAIL.n401 B 0.009313f
C453 VTAIL.n402 B 0.008796f
C454 VTAIL.n403 B 0.016368f
C455 VTAIL.n404 B 0.016368f
C456 VTAIL.n405 B 0.008796f
C457 VTAIL.n406 B 0.009313f
C458 VTAIL.n407 B 0.02079f
C459 VTAIL.n408 B 0.02079f
C460 VTAIL.n409 B 0.009313f
C461 VTAIL.n410 B 0.008796f
C462 VTAIL.n411 B 0.016368f
C463 VTAIL.n412 B 0.016368f
C464 VTAIL.n413 B 0.008796f
C465 VTAIL.n414 B 0.008796f
C466 VTAIL.n415 B 0.009313f
C467 VTAIL.n416 B 0.02079f
C468 VTAIL.n417 B 0.02079f
C469 VTAIL.n418 B 0.02079f
C470 VTAIL.n419 B 0.009054f
C471 VTAIL.n420 B 0.008796f
C472 VTAIL.n421 B 0.016368f
C473 VTAIL.n422 B 0.016368f
C474 VTAIL.n423 B 0.008796f
C475 VTAIL.n424 B 0.009313f
C476 VTAIL.n425 B 0.02079f
C477 VTAIL.n426 B 0.043248f
C478 VTAIL.n427 B 0.009313f
C479 VTAIL.n428 B 0.008796f
C480 VTAIL.n429 B 0.038505f
C481 VTAIL.n430 B 0.024039f
C482 VTAIL.n431 B 0.79834f
C483 VN.t3 B 1.45728f
C484 VN.t0 B 1.45662f
C485 VN.n0 B 1.10294f
C486 VN.t1 B 1.45728f
C487 VN.t2 B 1.45662f
C488 VN.n1 B 2.29528f
.ends

