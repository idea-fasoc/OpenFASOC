* NGSPICE file created from diff_pair_sample_1686.ext - technology: sky130A

.subckt diff_pair_sample_1686 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t11 VP.t0 VDD1.t4 B.t5 sky130_fd_pr__nfet_01v8 ad=2.2605 pd=14.03 as=2.2605 ps=14.03 w=13.7 l=0.72
X1 VDD2.t5 VN.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.2605 pd=14.03 as=5.343 ps=28.18 w=13.7 l=0.72
X2 B.t19 B.t17 B.t18 B.t11 sky130_fd_pr__nfet_01v8 ad=5.343 pd=28.18 as=0 ps=0 w=13.7 l=0.72
X3 VTAIL.t10 VP.t1 VDD1.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=2.2605 pd=14.03 as=2.2605 ps=14.03 w=13.7 l=0.72
X4 VTAIL.t5 VN.t1 VDD2.t4 B.t5 sky130_fd_pr__nfet_01v8 ad=2.2605 pd=14.03 as=2.2605 ps=14.03 w=13.7 l=0.72
X5 B.t16 B.t14 B.t15 B.t7 sky130_fd_pr__nfet_01v8 ad=5.343 pd=28.18 as=0 ps=0 w=13.7 l=0.72
X6 VDD1.t2 VP.t2 VTAIL.t9 B.t0 sky130_fd_pr__nfet_01v8 ad=2.2605 pd=14.03 as=5.343 ps=28.18 w=13.7 l=0.72
X7 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=5.343 pd=28.18 as=0 ps=0 w=13.7 l=0.72
X8 VDD1.t5 VP.t3 VTAIL.t8 B.t3 sky130_fd_pr__nfet_01v8 ad=2.2605 pd=14.03 as=5.343 ps=28.18 w=13.7 l=0.72
X9 VDD2.t3 VN.t2 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=5.343 pd=28.18 as=2.2605 ps=14.03 w=13.7 l=0.72
X10 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=5.343 pd=28.18 as=0 ps=0 w=13.7 l=0.72
X11 VDD2.t2 VN.t3 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.2605 pd=14.03 as=5.343 ps=28.18 w=13.7 l=0.72
X12 VDD1.t0 VP.t4 VTAIL.t7 B.t2 sky130_fd_pr__nfet_01v8 ad=5.343 pd=28.18 as=2.2605 ps=14.03 w=13.7 l=0.72
X13 VTAIL.t1 VN.t4 VDD2.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.2605 pd=14.03 as=2.2605 ps=14.03 w=13.7 l=0.72
X14 VDD1.t1 VP.t5 VTAIL.t6 B.t4 sky130_fd_pr__nfet_01v8 ad=5.343 pd=28.18 as=2.2605 ps=14.03 w=13.7 l=0.72
X15 VDD2.t0 VN.t5 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=5.343 pd=28.18 as=2.2605 ps=14.03 w=13.7 l=0.72
R0 VP.n3 VP.t5 535.115
R1 VP.n8 VP.t4 513.13
R2 VP.n12 VP.t1 513.13
R3 VP.n14 VP.t3 513.13
R4 VP.n6 VP.t2 513.13
R5 VP.n4 VP.t0 513.13
R6 VP.n15 VP.n14 161.3
R7 VP.n5 VP.n2 161.3
R8 VP.n7 VP.n6 161.3
R9 VP.n13 VP.n0 161.3
R10 VP.n12 VP.n11 161.3
R11 VP.n10 VP.n1 161.3
R12 VP.n9 VP.n8 161.3
R13 VP.n3 VP.n2 44.859
R14 VP.n9 VP.n7 42.5876
R15 VP.n8 VP.n1 27.752
R16 VP.n14 VP.n13 27.752
R17 VP.n6 VP.n5 27.752
R18 VP.n12 VP.n1 20.449
R19 VP.n13 VP.n12 20.449
R20 VP.n5 VP.n4 20.449
R21 VP.n4 VP.n3 19.9186
R22 VP.n7 VP.n2 0.189894
R23 VP.n10 VP.n9 0.189894
R24 VP.n11 VP.n10 0.189894
R25 VP.n11 VP.n0 0.189894
R26 VP.n15 VP.n0 0.189894
R27 VP VP.n15 0.0516364
R28 VDD1 VDD1.t1 65.9646
R29 VDD1.n1 VDD1.t0 65.8509
R30 VDD1.n1 VDD1.n0 63.953
R31 VDD1.n3 VDD1.n2 63.7821
R32 VDD1.n3 VDD1.n1 39.503
R33 VDD1.n2 VDD1.t4 1.44576
R34 VDD1.n2 VDD1.t2 1.44576
R35 VDD1.n0 VDD1.t3 1.44576
R36 VDD1.n0 VDD1.t5 1.44576
R37 VDD1 VDD1.n3 0.168603
R38 VTAIL.n7 VTAIL.t3 48.5487
R39 VTAIL.n11 VTAIL.t0 48.5485
R40 VTAIL.n2 VTAIL.t8 48.5485
R41 VTAIL.n10 VTAIL.t9 48.5485
R42 VTAIL.n9 VTAIL.n8 47.1035
R43 VTAIL.n6 VTAIL.n5 47.1035
R44 VTAIL.n1 VTAIL.n0 47.1033
R45 VTAIL.n4 VTAIL.n3 47.1033
R46 VTAIL.n6 VTAIL.n4 25.9876
R47 VTAIL.n11 VTAIL.n10 25.0824
R48 VTAIL.n0 VTAIL.t4 1.44576
R49 VTAIL.n0 VTAIL.t5 1.44576
R50 VTAIL.n3 VTAIL.t7 1.44576
R51 VTAIL.n3 VTAIL.t10 1.44576
R52 VTAIL.n8 VTAIL.t6 1.44576
R53 VTAIL.n8 VTAIL.t11 1.44576
R54 VTAIL.n5 VTAIL.t2 1.44576
R55 VTAIL.n5 VTAIL.t1 1.44576
R56 VTAIL.n9 VTAIL.n7 0.922914
R57 VTAIL.n2 VTAIL.n1 0.922914
R58 VTAIL.n7 VTAIL.n6 0.905672
R59 VTAIL.n10 VTAIL.n9 0.905672
R60 VTAIL.n4 VTAIL.n2 0.905672
R61 VTAIL VTAIL.n11 0.62119
R62 VTAIL VTAIL.n1 0.284983
R63 B.n97 B.t17 661.295
R64 B.n94 B.t10 661.295
R65 B.n501 B.t14 661.295
R66 B.n368 B.t6 661.295
R67 B.n691 B.n690 585
R68 B.n692 B.n691 585
R69 B.n300 B.n93 585
R70 B.n299 B.n298 585
R71 B.n297 B.n296 585
R72 B.n295 B.n294 585
R73 B.n293 B.n292 585
R74 B.n291 B.n290 585
R75 B.n289 B.n288 585
R76 B.n287 B.n286 585
R77 B.n285 B.n284 585
R78 B.n283 B.n282 585
R79 B.n281 B.n280 585
R80 B.n279 B.n278 585
R81 B.n277 B.n276 585
R82 B.n275 B.n274 585
R83 B.n273 B.n272 585
R84 B.n271 B.n270 585
R85 B.n269 B.n268 585
R86 B.n267 B.n266 585
R87 B.n265 B.n264 585
R88 B.n263 B.n262 585
R89 B.n261 B.n260 585
R90 B.n259 B.n258 585
R91 B.n257 B.n256 585
R92 B.n255 B.n254 585
R93 B.n253 B.n252 585
R94 B.n251 B.n250 585
R95 B.n249 B.n248 585
R96 B.n247 B.n246 585
R97 B.n245 B.n244 585
R98 B.n243 B.n242 585
R99 B.n241 B.n240 585
R100 B.n239 B.n238 585
R101 B.n237 B.n236 585
R102 B.n235 B.n234 585
R103 B.n233 B.n232 585
R104 B.n231 B.n230 585
R105 B.n229 B.n228 585
R106 B.n227 B.n226 585
R107 B.n225 B.n224 585
R108 B.n223 B.n222 585
R109 B.n221 B.n220 585
R110 B.n219 B.n218 585
R111 B.n217 B.n216 585
R112 B.n215 B.n214 585
R113 B.n213 B.n212 585
R114 B.n211 B.n210 585
R115 B.n209 B.n208 585
R116 B.n207 B.n206 585
R117 B.n205 B.n204 585
R118 B.n203 B.n202 585
R119 B.n201 B.n200 585
R120 B.n199 B.n198 585
R121 B.n197 B.n196 585
R122 B.n195 B.n194 585
R123 B.n193 B.n192 585
R124 B.n190 B.n189 585
R125 B.n188 B.n187 585
R126 B.n186 B.n185 585
R127 B.n184 B.n183 585
R128 B.n182 B.n181 585
R129 B.n180 B.n179 585
R130 B.n178 B.n177 585
R131 B.n176 B.n175 585
R132 B.n174 B.n173 585
R133 B.n172 B.n171 585
R134 B.n170 B.n169 585
R135 B.n168 B.n167 585
R136 B.n166 B.n165 585
R137 B.n164 B.n163 585
R138 B.n162 B.n161 585
R139 B.n160 B.n159 585
R140 B.n158 B.n157 585
R141 B.n156 B.n155 585
R142 B.n154 B.n153 585
R143 B.n152 B.n151 585
R144 B.n150 B.n149 585
R145 B.n148 B.n147 585
R146 B.n146 B.n145 585
R147 B.n144 B.n143 585
R148 B.n142 B.n141 585
R149 B.n140 B.n139 585
R150 B.n138 B.n137 585
R151 B.n136 B.n135 585
R152 B.n134 B.n133 585
R153 B.n132 B.n131 585
R154 B.n130 B.n129 585
R155 B.n128 B.n127 585
R156 B.n126 B.n125 585
R157 B.n124 B.n123 585
R158 B.n122 B.n121 585
R159 B.n120 B.n119 585
R160 B.n118 B.n117 585
R161 B.n116 B.n115 585
R162 B.n114 B.n113 585
R163 B.n112 B.n111 585
R164 B.n110 B.n109 585
R165 B.n108 B.n107 585
R166 B.n106 B.n105 585
R167 B.n104 B.n103 585
R168 B.n102 B.n101 585
R169 B.n100 B.n99 585
R170 B.n40 B.n39 585
R171 B.n689 B.n41 585
R172 B.n693 B.n41 585
R173 B.n688 B.n687 585
R174 B.n687 B.n37 585
R175 B.n686 B.n36 585
R176 B.n699 B.n36 585
R177 B.n685 B.n35 585
R178 B.n700 B.n35 585
R179 B.n684 B.n34 585
R180 B.n701 B.n34 585
R181 B.n683 B.n682 585
R182 B.n682 B.n30 585
R183 B.n681 B.n29 585
R184 B.n707 B.n29 585
R185 B.n680 B.n28 585
R186 B.n708 B.n28 585
R187 B.n679 B.n27 585
R188 B.n709 B.n27 585
R189 B.n678 B.n677 585
R190 B.n677 B.n23 585
R191 B.n676 B.n22 585
R192 B.n715 B.n22 585
R193 B.n675 B.n21 585
R194 B.n716 B.n21 585
R195 B.n674 B.n20 585
R196 B.n717 B.n20 585
R197 B.n673 B.n672 585
R198 B.n672 B.n16 585
R199 B.n671 B.n15 585
R200 B.n723 B.n15 585
R201 B.n670 B.n14 585
R202 B.n724 B.n14 585
R203 B.n669 B.n13 585
R204 B.n725 B.n13 585
R205 B.n668 B.n667 585
R206 B.n667 B.n12 585
R207 B.n666 B.n665 585
R208 B.n666 B.n8 585
R209 B.n664 B.n7 585
R210 B.n732 B.n7 585
R211 B.n663 B.n6 585
R212 B.n733 B.n6 585
R213 B.n662 B.n5 585
R214 B.n734 B.n5 585
R215 B.n661 B.n660 585
R216 B.n660 B.n4 585
R217 B.n659 B.n301 585
R218 B.n659 B.n658 585
R219 B.n648 B.n302 585
R220 B.n651 B.n302 585
R221 B.n650 B.n649 585
R222 B.n652 B.n650 585
R223 B.n647 B.n307 585
R224 B.n307 B.n306 585
R225 B.n646 B.n645 585
R226 B.n645 B.n644 585
R227 B.n309 B.n308 585
R228 B.n310 B.n309 585
R229 B.n637 B.n636 585
R230 B.n638 B.n637 585
R231 B.n635 B.n314 585
R232 B.n318 B.n314 585
R233 B.n634 B.n633 585
R234 B.n633 B.n632 585
R235 B.n316 B.n315 585
R236 B.n317 B.n316 585
R237 B.n625 B.n624 585
R238 B.n626 B.n625 585
R239 B.n623 B.n323 585
R240 B.n323 B.n322 585
R241 B.n622 B.n621 585
R242 B.n621 B.n620 585
R243 B.n325 B.n324 585
R244 B.n326 B.n325 585
R245 B.n613 B.n612 585
R246 B.n614 B.n613 585
R247 B.n611 B.n331 585
R248 B.n331 B.n330 585
R249 B.n610 B.n609 585
R250 B.n609 B.n608 585
R251 B.n333 B.n332 585
R252 B.n334 B.n333 585
R253 B.n601 B.n600 585
R254 B.n602 B.n601 585
R255 B.n337 B.n336 585
R256 B.n394 B.n393 585
R257 B.n395 B.n391 585
R258 B.n391 B.n338 585
R259 B.n397 B.n396 585
R260 B.n399 B.n390 585
R261 B.n402 B.n401 585
R262 B.n403 B.n389 585
R263 B.n405 B.n404 585
R264 B.n407 B.n388 585
R265 B.n410 B.n409 585
R266 B.n411 B.n387 585
R267 B.n413 B.n412 585
R268 B.n415 B.n386 585
R269 B.n418 B.n417 585
R270 B.n419 B.n385 585
R271 B.n421 B.n420 585
R272 B.n423 B.n384 585
R273 B.n426 B.n425 585
R274 B.n427 B.n383 585
R275 B.n429 B.n428 585
R276 B.n431 B.n382 585
R277 B.n434 B.n433 585
R278 B.n435 B.n381 585
R279 B.n437 B.n436 585
R280 B.n439 B.n380 585
R281 B.n442 B.n441 585
R282 B.n443 B.n379 585
R283 B.n445 B.n444 585
R284 B.n447 B.n378 585
R285 B.n450 B.n449 585
R286 B.n451 B.n377 585
R287 B.n453 B.n452 585
R288 B.n455 B.n376 585
R289 B.n458 B.n457 585
R290 B.n459 B.n375 585
R291 B.n461 B.n460 585
R292 B.n463 B.n374 585
R293 B.n466 B.n465 585
R294 B.n467 B.n373 585
R295 B.n469 B.n468 585
R296 B.n471 B.n372 585
R297 B.n474 B.n473 585
R298 B.n475 B.n371 585
R299 B.n477 B.n476 585
R300 B.n479 B.n370 585
R301 B.n482 B.n481 585
R302 B.n483 B.n367 585
R303 B.n486 B.n485 585
R304 B.n488 B.n366 585
R305 B.n491 B.n490 585
R306 B.n492 B.n365 585
R307 B.n494 B.n493 585
R308 B.n496 B.n364 585
R309 B.n499 B.n498 585
R310 B.n500 B.n363 585
R311 B.n505 B.n504 585
R312 B.n507 B.n362 585
R313 B.n510 B.n509 585
R314 B.n511 B.n361 585
R315 B.n513 B.n512 585
R316 B.n515 B.n360 585
R317 B.n518 B.n517 585
R318 B.n519 B.n359 585
R319 B.n521 B.n520 585
R320 B.n523 B.n358 585
R321 B.n526 B.n525 585
R322 B.n527 B.n357 585
R323 B.n529 B.n528 585
R324 B.n531 B.n356 585
R325 B.n534 B.n533 585
R326 B.n535 B.n355 585
R327 B.n537 B.n536 585
R328 B.n539 B.n354 585
R329 B.n542 B.n541 585
R330 B.n543 B.n353 585
R331 B.n545 B.n544 585
R332 B.n547 B.n352 585
R333 B.n550 B.n549 585
R334 B.n551 B.n351 585
R335 B.n553 B.n552 585
R336 B.n555 B.n350 585
R337 B.n558 B.n557 585
R338 B.n559 B.n349 585
R339 B.n561 B.n560 585
R340 B.n563 B.n348 585
R341 B.n566 B.n565 585
R342 B.n567 B.n347 585
R343 B.n569 B.n568 585
R344 B.n571 B.n346 585
R345 B.n574 B.n573 585
R346 B.n575 B.n345 585
R347 B.n577 B.n576 585
R348 B.n579 B.n344 585
R349 B.n582 B.n581 585
R350 B.n583 B.n343 585
R351 B.n585 B.n584 585
R352 B.n587 B.n342 585
R353 B.n590 B.n589 585
R354 B.n591 B.n341 585
R355 B.n593 B.n592 585
R356 B.n595 B.n340 585
R357 B.n598 B.n597 585
R358 B.n599 B.n339 585
R359 B.n604 B.n603 585
R360 B.n603 B.n602 585
R361 B.n605 B.n335 585
R362 B.n335 B.n334 585
R363 B.n607 B.n606 585
R364 B.n608 B.n607 585
R365 B.n329 B.n328 585
R366 B.n330 B.n329 585
R367 B.n616 B.n615 585
R368 B.n615 B.n614 585
R369 B.n617 B.n327 585
R370 B.n327 B.n326 585
R371 B.n619 B.n618 585
R372 B.n620 B.n619 585
R373 B.n321 B.n320 585
R374 B.n322 B.n321 585
R375 B.n628 B.n627 585
R376 B.n627 B.n626 585
R377 B.n629 B.n319 585
R378 B.n319 B.n317 585
R379 B.n631 B.n630 585
R380 B.n632 B.n631 585
R381 B.n313 B.n312 585
R382 B.n318 B.n313 585
R383 B.n640 B.n639 585
R384 B.n639 B.n638 585
R385 B.n641 B.n311 585
R386 B.n311 B.n310 585
R387 B.n643 B.n642 585
R388 B.n644 B.n643 585
R389 B.n305 B.n304 585
R390 B.n306 B.n305 585
R391 B.n654 B.n653 585
R392 B.n653 B.n652 585
R393 B.n655 B.n303 585
R394 B.n651 B.n303 585
R395 B.n657 B.n656 585
R396 B.n658 B.n657 585
R397 B.n3 B.n0 585
R398 B.n4 B.n3 585
R399 B.n731 B.n1 585
R400 B.n732 B.n731 585
R401 B.n730 B.n729 585
R402 B.n730 B.n8 585
R403 B.n728 B.n9 585
R404 B.n12 B.n9 585
R405 B.n727 B.n726 585
R406 B.n726 B.n725 585
R407 B.n11 B.n10 585
R408 B.n724 B.n11 585
R409 B.n722 B.n721 585
R410 B.n723 B.n722 585
R411 B.n720 B.n17 585
R412 B.n17 B.n16 585
R413 B.n719 B.n718 585
R414 B.n718 B.n717 585
R415 B.n19 B.n18 585
R416 B.n716 B.n19 585
R417 B.n714 B.n713 585
R418 B.n715 B.n714 585
R419 B.n712 B.n24 585
R420 B.n24 B.n23 585
R421 B.n711 B.n710 585
R422 B.n710 B.n709 585
R423 B.n26 B.n25 585
R424 B.n708 B.n26 585
R425 B.n706 B.n705 585
R426 B.n707 B.n706 585
R427 B.n704 B.n31 585
R428 B.n31 B.n30 585
R429 B.n703 B.n702 585
R430 B.n702 B.n701 585
R431 B.n33 B.n32 585
R432 B.n700 B.n33 585
R433 B.n698 B.n697 585
R434 B.n699 B.n698 585
R435 B.n696 B.n38 585
R436 B.n38 B.n37 585
R437 B.n695 B.n694 585
R438 B.n694 B.n693 585
R439 B.n735 B.n734 585
R440 B.n733 B.n2 585
R441 B.n694 B.n40 478.086
R442 B.n691 B.n41 478.086
R443 B.n601 B.n339 478.086
R444 B.n603 B.n337 478.086
R445 B.n692 B.n92 256.663
R446 B.n692 B.n91 256.663
R447 B.n692 B.n90 256.663
R448 B.n692 B.n89 256.663
R449 B.n692 B.n88 256.663
R450 B.n692 B.n87 256.663
R451 B.n692 B.n86 256.663
R452 B.n692 B.n85 256.663
R453 B.n692 B.n84 256.663
R454 B.n692 B.n83 256.663
R455 B.n692 B.n82 256.663
R456 B.n692 B.n81 256.663
R457 B.n692 B.n80 256.663
R458 B.n692 B.n79 256.663
R459 B.n692 B.n78 256.663
R460 B.n692 B.n77 256.663
R461 B.n692 B.n76 256.663
R462 B.n692 B.n75 256.663
R463 B.n692 B.n74 256.663
R464 B.n692 B.n73 256.663
R465 B.n692 B.n72 256.663
R466 B.n692 B.n71 256.663
R467 B.n692 B.n70 256.663
R468 B.n692 B.n69 256.663
R469 B.n692 B.n68 256.663
R470 B.n692 B.n67 256.663
R471 B.n692 B.n66 256.663
R472 B.n692 B.n65 256.663
R473 B.n692 B.n64 256.663
R474 B.n692 B.n63 256.663
R475 B.n692 B.n62 256.663
R476 B.n692 B.n61 256.663
R477 B.n692 B.n60 256.663
R478 B.n692 B.n59 256.663
R479 B.n692 B.n58 256.663
R480 B.n692 B.n57 256.663
R481 B.n692 B.n56 256.663
R482 B.n692 B.n55 256.663
R483 B.n692 B.n54 256.663
R484 B.n692 B.n53 256.663
R485 B.n692 B.n52 256.663
R486 B.n692 B.n51 256.663
R487 B.n692 B.n50 256.663
R488 B.n692 B.n49 256.663
R489 B.n692 B.n48 256.663
R490 B.n692 B.n47 256.663
R491 B.n692 B.n46 256.663
R492 B.n692 B.n45 256.663
R493 B.n692 B.n44 256.663
R494 B.n692 B.n43 256.663
R495 B.n692 B.n42 256.663
R496 B.n392 B.n338 256.663
R497 B.n398 B.n338 256.663
R498 B.n400 B.n338 256.663
R499 B.n406 B.n338 256.663
R500 B.n408 B.n338 256.663
R501 B.n414 B.n338 256.663
R502 B.n416 B.n338 256.663
R503 B.n422 B.n338 256.663
R504 B.n424 B.n338 256.663
R505 B.n430 B.n338 256.663
R506 B.n432 B.n338 256.663
R507 B.n438 B.n338 256.663
R508 B.n440 B.n338 256.663
R509 B.n446 B.n338 256.663
R510 B.n448 B.n338 256.663
R511 B.n454 B.n338 256.663
R512 B.n456 B.n338 256.663
R513 B.n462 B.n338 256.663
R514 B.n464 B.n338 256.663
R515 B.n470 B.n338 256.663
R516 B.n472 B.n338 256.663
R517 B.n478 B.n338 256.663
R518 B.n480 B.n338 256.663
R519 B.n487 B.n338 256.663
R520 B.n489 B.n338 256.663
R521 B.n495 B.n338 256.663
R522 B.n497 B.n338 256.663
R523 B.n506 B.n338 256.663
R524 B.n508 B.n338 256.663
R525 B.n514 B.n338 256.663
R526 B.n516 B.n338 256.663
R527 B.n522 B.n338 256.663
R528 B.n524 B.n338 256.663
R529 B.n530 B.n338 256.663
R530 B.n532 B.n338 256.663
R531 B.n538 B.n338 256.663
R532 B.n540 B.n338 256.663
R533 B.n546 B.n338 256.663
R534 B.n548 B.n338 256.663
R535 B.n554 B.n338 256.663
R536 B.n556 B.n338 256.663
R537 B.n562 B.n338 256.663
R538 B.n564 B.n338 256.663
R539 B.n570 B.n338 256.663
R540 B.n572 B.n338 256.663
R541 B.n578 B.n338 256.663
R542 B.n580 B.n338 256.663
R543 B.n586 B.n338 256.663
R544 B.n588 B.n338 256.663
R545 B.n594 B.n338 256.663
R546 B.n596 B.n338 256.663
R547 B.n737 B.n736 256.663
R548 B.n101 B.n100 163.367
R549 B.n105 B.n104 163.367
R550 B.n109 B.n108 163.367
R551 B.n113 B.n112 163.367
R552 B.n117 B.n116 163.367
R553 B.n121 B.n120 163.367
R554 B.n125 B.n124 163.367
R555 B.n129 B.n128 163.367
R556 B.n133 B.n132 163.367
R557 B.n137 B.n136 163.367
R558 B.n141 B.n140 163.367
R559 B.n145 B.n144 163.367
R560 B.n149 B.n148 163.367
R561 B.n153 B.n152 163.367
R562 B.n157 B.n156 163.367
R563 B.n161 B.n160 163.367
R564 B.n165 B.n164 163.367
R565 B.n169 B.n168 163.367
R566 B.n173 B.n172 163.367
R567 B.n177 B.n176 163.367
R568 B.n181 B.n180 163.367
R569 B.n185 B.n184 163.367
R570 B.n189 B.n188 163.367
R571 B.n194 B.n193 163.367
R572 B.n198 B.n197 163.367
R573 B.n202 B.n201 163.367
R574 B.n206 B.n205 163.367
R575 B.n210 B.n209 163.367
R576 B.n214 B.n213 163.367
R577 B.n218 B.n217 163.367
R578 B.n222 B.n221 163.367
R579 B.n226 B.n225 163.367
R580 B.n230 B.n229 163.367
R581 B.n234 B.n233 163.367
R582 B.n238 B.n237 163.367
R583 B.n242 B.n241 163.367
R584 B.n246 B.n245 163.367
R585 B.n250 B.n249 163.367
R586 B.n254 B.n253 163.367
R587 B.n258 B.n257 163.367
R588 B.n262 B.n261 163.367
R589 B.n266 B.n265 163.367
R590 B.n270 B.n269 163.367
R591 B.n274 B.n273 163.367
R592 B.n278 B.n277 163.367
R593 B.n282 B.n281 163.367
R594 B.n286 B.n285 163.367
R595 B.n290 B.n289 163.367
R596 B.n294 B.n293 163.367
R597 B.n298 B.n297 163.367
R598 B.n691 B.n93 163.367
R599 B.n601 B.n333 163.367
R600 B.n609 B.n333 163.367
R601 B.n609 B.n331 163.367
R602 B.n613 B.n331 163.367
R603 B.n613 B.n325 163.367
R604 B.n621 B.n325 163.367
R605 B.n621 B.n323 163.367
R606 B.n625 B.n323 163.367
R607 B.n625 B.n316 163.367
R608 B.n633 B.n316 163.367
R609 B.n633 B.n314 163.367
R610 B.n637 B.n314 163.367
R611 B.n637 B.n309 163.367
R612 B.n645 B.n309 163.367
R613 B.n645 B.n307 163.367
R614 B.n650 B.n307 163.367
R615 B.n650 B.n302 163.367
R616 B.n659 B.n302 163.367
R617 B.n660 B.n659 163.367
R618 B.n660 B.n5 163.367
R619 B.n6 B.n5 163.367
R620 B.n7 B.n6 163.367
R621 B.n666 B.n7 163.367
R622 B.n667 B.n666 163.367
R623 B.n667 B.n13 163.367
R624 B.n14 B.n13 163.367
R625 B.n15 B.n14 163.367
R626 B.n672 B.n15 163.367
R627 B.n672 B.n20 163.367
R628 B.n21 B.n20 163.367
R629 B.n22 B.n21 163.367
R630 B.n677 B.n22 163.367
R631 B.n677 B.n27 163.367
R632 B.n28 B.n27 163.367
R633 B.n29 B.n28 163.367
R634 B.n682 B.n29 163.367
R635 B.n682 B.n34 163.367
R636 B.n35 B.n34 163.367
R637 B.n36 B.n35 163.367
R638 B.n687 B.n36 163.367
R639 B.n687 B.n41 163.367
R640 B.n393 B.n391 163.367
R641 B.n397 B.n391 163.367
R642 B.n401 B.n399 163.367
R643 B.n405 B.n389 163.367
R644 B.n409 B.n407 163.367
R645 B.n413 B.n387 163.367
R646 B.n417 B.n415 163.367
R647 B.n421 B.n385 163.367
R648 B.n425 B.n423 163.367
R649 B.n429 B.n383 163.367
R650 B.n433 B.n431 163.367
R651 B.n437 B.n381 163.367
R652 B.n441 B.n439 163.367
R653 B.n445 B.n379 163.367
R654 B.n449 B.n447 163.367
R655 B.n453 B.n377 163.367
R656 B.n457 B.n455 163.367
R657 B.n461 B.n375 163.367
R658 B.n465 B.n463 163.367
R659 B.n469 B.n373 163.367
R660 B.n473 B.n471 163.367
R661 B.n477 B.n371 163.367
R662 B.n481 B.n479 163.367
R663 B.n486 B.n367 163.367
R664 B.n490 B.n488 163.367
R665 B.n494 B.n365 163.367
R666 B.n498 B.n496 163.367
R667 B.n505 B.n363 163.367
R668 B.n509 B.n507 163.367
R669 B.n513 B.n361 163.367
R670 B.n517 B.n515 163.367
R671 B.n521 B.n359 163.367
R672 B.n525 B.n523 163.367
R673 B.n529 B.n357 163.367
R674 B.n533 B.n531 163.367
R675 B.n537 B.n355 163.367
R676 B.n541 B.n539 163.367
R677 B.n545 B.n353 163.367
R678 B.n549 B.n547 163.367
R679 B.n553 B.n351 163.367
R680 B.n557 B.n555 163.367
R681 B.n561 B.n349 163.367
R682 B.n565 B.n563 163.367
R683 B.n569 B.n347 163.367
R684 B.n573 B.n571 163.367
R685 B.n577 B.n345 163.367
R686 B.n581 B.n579 163.367
R687 B.n585 B.n343 163.367
R688 B.n589 B.n587 163.367
R689 B.n593 B.n341 163.367
R690 B.n597 B.n595 163.367
R691 B.n603 B.n335 163.367
R692 B.n607 B.n335 163.367
R693 B.n607 B.n329 163.367
R694 B.n615 B.n329 163.367
R695 B.n615 B.n327 163.367
R696 B.n619 B.n327 163.367
R697 B.n619 B.n321 163.367
R698 B.n627 B.n321 163.367
R699 B.n627 B.n319 163.367
R700 B.n631 B.n319 163.367
R701 B.n631 B.n313 163.367
R702 B.n639 B.n313 163.367
R703 B.n639 B.n311 163.367
R704 B.n643 B.n311 163.367
R705 B.n643 B.n305 163.367
R706 B.n653 B.n305 163.367
R707 B.n653 B.n303 163.367
R708 B.n657 B.n303 163.367
R709 B.n657 B.n3 163.367
R710 B.n735 B.n3 163.367
R711 B.n731 B.n2 163.367
R712 B.n731 B.n730 163.367
R713 B.n730 B.n9 163.367
R714 B.n726 B.n9 163.367
R715 B.n726 B.n11 163.367
R716 B.n722 B.n11 163.367
R717 B.n722 B.n17 163.367
R718 B.n718 B.n17 163.367
R719 B.n718 B.n19 163.367
R720 B.n714 B.n19 163.367
R721 B.n714 B.n24 163.367
R722 B.n710 B.n24 163.367
R723 B.n710 B.n26 163.367
R724 B.n706 B.n26 163.367
R725 B.n706 B.n31 163.367
R726 B.n702 B.n31 163.367
R727 B.n702 B.n33 163.367
R728 B.n698 B.n33 163.367
R729 B.n698 B.n38 163.367
R730 B.n694 B.n38 163.367
R731 B.n94 B.t12 89.8907
R732 B.n501 B.t16 89.8907
R733 B.n97 B.t18 89.8729
R734 B.n368 B.t9 89.8729
R735 B.n42 B.n40 71.676
R736 B.n101 B.n43 71.676
R737 B.n105 B.n44 71.676
R738 B.n109 B.n45 71.676
R739 B.n113 B.n46 71.676
R740 B.n117 B.n47 71.676
R741 B.n121 B.n48 71.676
R742 B.n125 B.n49 71.676
R743 B.n129 B.n50 71.676
R744 B.n133 B.n51 71.676
R745 B.n137 B.n52 71.676
R746 B.n141 B.n53 71.676
R747 B.n145 B.n54 71.676
R748 B.n149 B.n55 71.676
R749 B.n153 B.n56 71.676
R750 B.n157 B.n57 71.676
R751 B.n161 B.n58 71.676
R752 B.n165 B.n59 71.676
R753 B.n169 B.n60 71.676
R754 B.n173 B.n61 71.676
R755 B.n177 B.n62 71.676
R756 B.n181 B.n63 71.676
R757 B.n185 B.n64 71.676
R758 B.n189 B.n65 71.676
R759 B.n194 B.n66 71.676
R760 B.n198 B.n67 71.676
R761 B.n202 B.n68 71.676
R762 B.n206 B.n69 71.676
R763 B.n210 B.n70 71.676
R764 B.n214 B.n71 71.676
R765 B.n218 B.n72 71.676
R766 B.n222 B.n73 71.676
R767 B.n226 B.n74 71.676
R768 B.n230 B.n75 71.676
R769 B.n234 B.n76 71.676
R770 B.n238 B.n77 71.676
R771 B.n242 B.n78 71.676
R772 B.n246 B.n79 71.676
R773 B.n250 B.n80 71.676
R774 B.n254 B.n81 71.676
R775 B.n258 B.n82 71.676
R776 B.n262 B.n83 71.676
R777 B.n266 B.n84 71.676
R778 B.n270 B.n85 71.676
R779 B.n274 B.n86 71.676
R780 B.n278 B.n87 71.676
R781 B.n282 B.n88 71.676
R782 B.n286 B.n89 71.676
R783 B.n290 B.n90 71.676
R784 B.n294 B.n91 71.676
R785 B.n298 B.n92 71.676
R786 B.n93 B.n92 71.676
R787 B.n297 B.n91 71.676
R788 B.n293 B.n90 71.676
R789 B.n289 B.n89 71.676
R790 B.n285 B.n88 71.676
R791 B.n281 B.n87 71.676
R792 B.n277 B.n86 71.676
R793 B.n273 B.n85 71.676
R794 B.n269 B.n84 71.676
R795 B.n265 B.n83 71.676
R796 B.n261 B.n82 71.676
R797 B.n257 B.n81 71.676
R798 B.n253 B.n80 71.676
R799 B.n249 B.n79 71.676
R800 B.n245 B.n78 71.676
R801 B.n241 B.n77 71.676
R802 B.n237 B.n76 71.676
R803 B.n233 B.n75 71.676
R804 B.n229 B.n74 71.676
R805 B.n225 B.n73 71.676
R806 B.n221 B.n72 71.676
R807 B.n217 B.n71 71.676
R808 B.n213 B.n70 71.676
R809 B.n209 B.n69 71.676
R810 B.n205 B.n68 71.676
R811 B.n201 B.n67 71.676
R812 B.n197 B.n66 71.676
R813 B.n193 B.n65 71.676
R814 B.n188 B.n64 71.676
R815 B.n184 B.n63 71.676
R816 B.n180 B.n62 71.676
R817 B.n176 B.n61 71.676
R818 B.n172 B.n60 71.676
R819 B.n168 B.n59 71.676
R820 B.n164 B.n58 71.676
R821 B.n160 B.n57 71.676
R822 B.n156 B.n56 71.676
R823 B.n152 B.n55 71.676
R824 B.n148 B.n54 71.676
R825 B.n144 B.n53 71.676
R826 B.n140 B.n52 71.676
R827 B.n136 B.n51 71.676
R828 B.n132 B.n50 71.676
R829 B.n128 B.n49 71.676
R830 B.n124 B.n48 71.676
R831 B.n120 B.n47 71.676
R832 B.n116 B.n46 71.676
R833 B.n112 B.n45 71.676
R834 B.n108 B.n44 71.676
R835 B.n104 B.n43 71.676
R836 B.n100 B.n42 71.676
R837 B.n392 B.n337 71.676
R838 B.n398 B.n397 71.676
R839 B.n401 B.n400 71.676
R840 B.n406 B.n405 71.676
R841 B.n409 B.n408 71.676
R842 B.n414 B.n413 71.676
R843 B.n417 B.n416 71.676
R844 B.n422 B.n421 71.676
R845 B.n425 B.n424 71.676
R846 B.n430 B.n429 71.676
R847 B.n433 B.n432 71.676
R848 B.n438 B.n437 71.676
R849 B.n441 B.n440 71.676
R850 B.n446 B.n445 71.676
R851 B.n449 B.n448 71.676
R852 B.n454 B.n453 71.676
R853 B.n457 B.n456 71.676
R854 B.n462 B.n461 71.676
R855 B.n465 B.n464 71.676
R856 B.n470 B.n469 71.676
R857 B.n473 B.n472 71.676
R858 B.n478 B.n477 71.676
R859 B.n481 B.n480 71.676
R860 B.n487 B.n486 71.676
R861 B.n490 B.n489 71.676
R862 B.n495 B.n494 71.676
R863 B.n498 B.n497 71.676
R864 B.n506 B.n505 71.676
R865 B.n509 B.n508 71.676
R866 B.n514 B.n513 71.676
R867 B.n517 B.n516 71.676
R868 B.n522 B.n521 71.676
R869 B.n525 B.n524 71.676
R870 B.n530 B.n529 71.676
R871 B.n533 B.n532 71.676
R872 B.n538 B.n537 71.676
R873 B.n541 B.n540 71.676
R874 B.n546 B.n545 71.676
R875 B.n549 B.n548 71.676
R876 B.n554 B.n553 71.676
R877 B.n557 B.n556 71.676
R878 B.n562 B.n561 71.676
R879 B.n565 B.n564 71.676
R880 B.n570 B.n569 71.676
R881 B.n573 B.n572 71.676
R882 B.n578 B.n577 71.676
R883 B.n581 B.n580 71.676
R884 B.n586 B.n585 71.676
R885 B.n589 B.n588 71.676
R886 B.n594 B.n593 71.676
R887 B.n597 B.n596 71.676
R888 B.n393 B.n392 71.676
R889 B.n399 B.n398 71.676
R890 B.n400 B.n389 71.676
R891 B.n407 B.n406 71.676
R892 B.n408 B.n387 71.676
R893 B.n415 B.n414 71.676
R894 B.n416 B.n385 71.676
R895 B.n423 B.n422 71.676
R896 B.n424 B.n383 71.676
R897 B.n431 B.n430 71.676
R898 B.n432 B.n381 71.676
R899 B.n439 B.n438 71.676
R900 B.n440 B.n379 71.676
R901 B.n447 B.n446 71.676
R902 B.n448 B.n377 71.676
R903 B.n455 B.n454 71.676
R904 B.n456 B.n375 71.676
R905 B.n463 B.n462 71.676
R906 B.n464 B.n373 71.676
R907 B.n471 B.n470 71.676
R908 B.n472 B.n371 71.676
R909 B.n479 B.n478 71.676
R910 B.n480 B.n367 71.676
R911 B.n488 B.n487 71.676
R912 B.n489 B.n365 71.676
R913 B.n496 B.n495 71.676
R914 B.n497 B.n363 71.676
R915 B.n507 B.n506 71.676
R916 B.n508 B.n361 71.676
R917 B.n515 B.n514 71.676
R918 B.n516 B.n359 71.676
R919 B.n523 B.n522 71.676
R920 B.n524 B.n357 71.676
R921 B.n531 B.n530 71.676
R922 B.n532 B.n355 71.676
R923 B.n539 B.n538 71.676
R924 B.n540 B.n353 71.676
R925 B.n547 B.n546 71.676
R926 B.n548 B.n351 71.676
R927 B.n555 B.n554 71.676
R928 B.n556 B.n349 71.676
R929 B.n563 B.n562 71.676
R930 B.n564 B.n347 71.676
R931 B.n571 B.n570 71.676
R932 B.n572 B.n345 71.676
R933 B.n579 B.n578 71.676
R934 B.n580 B.n343 71.676
R935 B.n587 B.n586 71.676
R936 B.n588 B.n341 71.676
R937 B.n595 B.n594 71.676
R938 B.n596 B.n339 71.676
R939 B.n736 B.n735 71.676
R940 B.n736 B.n2 71.676
R941 B.n602 B.n338 70.1454
R942 B.n693 B.n692 70.1454
R943 B.n95 B.t13 69.5271
R944 B.n502 B.t15 69.5271
R945 B.n98 B.t19 69.5093
R946 B.n369 B.t8 69.5093
R947 B.n191 B.n98 59.5399
R948 B.n96 B.n95 59.5399
R949 B.n503 B.n502 59.5399
R950 B.n484 B.n369 59.5399
R951 B.n602 B.n334 39.4208
R952 B.n608 B.n334 39.4208
R953 B.n608 B.n330 39.4208
R954 B.n614 B.n330 39.4208
R955 B.n620 B.n326 39.4208
R956 B.n620 B.n322 39.4208
R957 B.n626 B.n322 39.4208
R958 B.n626 B.n317 39.4208
R959 B.n632 B.n317 39.4208
R960 B.n632 B.n318 39.4208
R961 B.n638 B.n310 39.4208
R962 B.n644 B.n310 39.4208
R963 B.n652 B.n306 39.4208
R964 B.n652 B.n651 39.4208
R965 B.n658 B.n4 39.4208
R966 B.n734 B.n4 39.4208
R967 B.n734 B.n733 39.4208
R968 B.n733 B.n732 39.4208
R969 B.n732 B.n8 39.4208
R970 B.n725 B.n12 39.4208
R971 B.n725 B.n724 39.4208
R972 B.n723 B.n16 39.4208
R973 B.n717 B.n16 39.4208
R974 B.n716 B.n715 39.4208
R975 B.n715 B.n23 39.4208
R976 B.n709 B.n23 39.4208
R977 B.n709 B.n708 39.4208
R978 B.n708 B.n707 39.4208
R979 B.n707 B.n30 39.4208
R980 B.n701 B.n700 39.4208
R981 B.n700 B.n699 39.4208
R982 B.n699 B.n37 39.4208
R983 B.n693 B.n37 39.4208
R984 B.n614 B.t7 34.7831
R985 B.n701 B.t11 34.7831
R986 B.n638 B.t2 32.4643
R987 B.n717 B.t0 32.4643
R988 B.n604 B.n336 31.0639
R989 B.n600 B.n599 31.0639
R990 B.n690 B.n689 31.0639
R991 B.n695 B.n39 31.0639
R992 B.t1 B.n306 28.986
R993 B.n724 B.t5 28.986
R994 B.n658 B.t3 25.5077
R995 B.t4 B.n8 25.5077
R996 B.n98 B.n97 20.3641
R997 B.n95 B.n94 20.3641
R998 B.n502 B.n501 20.3641
R999 B.n369 B.n368 20.3641
R1000 B B.n737 18.0485
R1001 B.n651 B.t3 13.9135
R1002 B.n12 B.t4 13.9135
R1003 B.n605 B.n604 10.6151
R1004 B.n606 B.n605 10.6151
R1005 B.n606 B.n328 10.6151
R1006 B.n616 B.n328 10.6151
R1007 B.n617 B.n616 10.6151
R1008 B.n618 B.n617 10.6151
R1009 B.n618 B.n320 10.6151
R1010 B.n628 B.n320 10.6151
R1011 B.n629 B.n628 10.6151
R1012 B.n630 B.n629 10.6151
R1013 B.n630 B.n312 10.6151
R1014 B.n640 B.n312 10.6151
R1015 B.n641 B.n640 10.6151
R1016 B.n642 B.n641 10.6151
R1017 B.n642 B.n304 10.6151
R1018 B.n654 B.n304 10.6151
R1019 B.n655 B.n654 10.6151
R1020 B.n656 B.n655 10.6151
R1021 B.n656 B.n0 10.6151
R1022 B.n394 B.n336 10.6151
R1023 B.n395 B.n394 10.6151
R1024 B.n396 B.n395 10.6151
R1025 B.n396 B.n390 10.6151
R1026 B.n402 B.n390 10.6151
R1027 B.n403 B.n402 10.6151
R1028 B.n404 B.n403 10.6151
R1029 B.n404 B.n388 10.6151
R1030 B.n410 B.n388 10.6151
R1031 B.n411 B.n410 10.6151
R1032 B.n412 B.n411 10.6151
R1033 B.n412 B.n386 10.6151
R1034 B.n418 B.n386 10.6151
R1035 B.n419 B.n418 10.6151
R1036 B.n420 B.n419 10.6151
R1037 B.n420 B.n384 10.6151
R1038 B.n426 B.n384 10.6151
R1039 B.n427 B.n426 10.6151
R1040 B.n428 B.n427 10.6151
R1041 B.n428 B.n382 10.6151
R1042 B.n434 B.n382 10.6151
R1043 B.n435 B.n434 10.6151
R1044 B.n436 B.n435 10.6151
R1045 B.n436 B.n380 10.6151
R1046 B.n442 B.n380 10.6151
R1047 B.n443 B.n442 10.6151
R1048 B.n444 B.n443 10.6151
R1049 B.n444 B.n378 10.6151
R1050 B.n450 B.n378 10.6151
R1051 B.n451 B.n450 10.6151
R1052 B.n452 B.n451 10.6151
R1053 B.n452 B.n376 10.6151
R1054 B.n458 B.n376 10.6151
R1055 B.n459 B.n458 10.6151
R1056 B.n460 B.n459 10.6151
R1057 B.n460 B.n374 10.6151
R1058 B.n466 B.n374 10.6151
R1059 B.n467 B.n466 10.6151
R1060 B.n468 B.n467 10.6151
R1061 B.n468 B.n372 10.6151
R1062 B.n474 B.n372 10.6151
R1063 B.n475 B.n474 10.6151
R1064 B.n476 B.n475 10.6151
R1065 B.n476 B.n370 10.6151
R1066 B.n482 B.n370 10.6151
R1067 B.n483 B.n482 10.6151
R1068 B.n485 B.n366 10.6151
R1069 B.n491 B.n366 10.6151
R1070 B.n492 B.n491 10.6151
R1071 B.n493 B.n492 10.6151
R1072 B.n493 B.n364 10.6151
R1073 B.n499 B.n364 10.6151
R1074 B.n500 B.n499 10.6151
R1075 B.n504 B.n500 10.6151
R1076 B.n510 B.n362 10.6151
R1077 B.n511 B.n510 10.6151
R1078 B.n512 B.n511 10.6151
R1079 B.n512 B.n360 10.6151
R1080 B.n518 B.n360 10.6151
R1081 B.n519 B.n518 10.6151
R1082 B.n520 B.n519 10.6151
R1083 B.n520 B.n358 10.6151
R1084 B.n526 B.n358 10.6151
R1085 B.n527 B.n526 10.6151
R1086 B.n528 B.n527 10.6151
R1087 B.n528 B.n356 10.6151
R1088 B.n534 B.n356 10.6151
R1089 B.n535 B.n534 10.6151
R1090 B.n536 B.n535 10.6151
R1091 B.n536 B.n354 10.6151
R1092 B.n542 B.n354 10.6151
R1093 B.n543 B.n542 10.6151
R1094 B.n544 B.n543 10.6151
R1095 B.n544 B.n352 10.6151
R1096 B.n550 B.n352 10.6151
R1097 B.n551 B.n550 10.6151
R1098 B.n552 B.n551 10.6151
R1099 B.n552 B.n350 10.6151
R1100 B.n558 B.n350 10.6151
R1101 B.n559 B.n558 10.6151
R1102 B.n560 B.n559 10.6151
R1103 B.n560 B.n348 10.6151
R1104 B.n566 B.n348 10.6151
R1105 B.n567 B.n566 10.6151
R1106 B.n568 B.n567 10.6151
R1107 B.n568 B.n346 10.6151
R1108 B.n574 B.n346 10.6151
R1109 B.n575 B.n574 10.6151
R1110 B.n576 B.n575 10.6151
R1111 B.n576 B.n344 10.6151
R1112 B.n582 B.n344 10.6151
R1113 B.n583 B.n582 10.6151
R1114 B.n584 B.n583 10.6151
R1115 B.n584 B.n342 10.6151
R1116 B.n590 B.n342 10.6151
R1117 B.n591 B.n590 10.6151
R1118 B.n592 B.n591 10.6151
R1119 B.n592 B.n340 10.6151
R1120 B.n598 B.n340 10.6151
R1121 B.n599 B.n598 10.6151
R1122 B.n600 B.n332 10.6151
R1123 B.n610 B.n332 10.6151
R1124 B.n611 B.n610 10.6151
R1125 B.n612 B.n611 10.6151
R1126 B.n612 B.n324 10.6151
R1127 B.n622 B.n324 10.6151
R1128 B.n623 B.n622 10.6151
R1129 B.n624 B.n623 10.6151
R1130 B.n624 B.n315 10.6151
R1131 B.n634 B.n315 10.6151
R1132 B.n635 B.n634 10.6151
R1133 B.n636 B.n635 10.6151
R1134 B.n636 B.n308 10.6151
R1135 B.n646 B.n308 10.6151
R1136 B.n647 B.n646 10.6151
R1137 B.n649 B.n647 10.6151
R1138 B.n649 B.n648 10.6151
R1139 B.n648 B.n301 10.6151
R1140 B.n661 B.n301 10.6151
R1141 B.n662 B.n661 10.6151
R1142 B.n663 B.n662 10.6151
R1143 B.n664 B.n663 10.6151
R1144 B.n665 B.n664 10.6151
R1145 B.n668 B.n665 10.6151
R1146 B.n669 B.n668 10.6151
R1147 B.n670 B.n669 10.6151
R1148 B.n671 B.n670 10.6151
R1149 B.n673 B.n671 10.6151
R1150 B.n674 B.n673 10.6151
R1151 B.n675 B.n674 10.6151
R1152 B.n676 B.n675 10.6151
R1153 B.n678 B.n676 10.6151
R1154 B.n679 B.n678 10.6151
R1155 B.n680 B.n679 10.6151
R1156 B.n681 B.n680 10.6151
R1157 B.n683 B.n681 10.6151
R1158 B.n684 B.n683 10.6151
R1159 B.n685 B.n684 10.6151
R1160 B.n686 B.n685 10.6151
R1161 B.n688 B.n686 10.6151
R1162 B.n689 B.n688 10.6151
R1163 B.n729 B.n1 10.6151
R1164 B.n729 B.n728 10.6151
R1165 B.n728 B.n727 10.6151
R1166 B.n727 B.n10 10.6151
R1167 B.n721 B.n10 10.6151
R1168 B.n721 B.n720 10.6151
R1169 B.n720 B.n719 10.6151
R1170 B.n719 B.n18 10.6151
R1171 B.n713 B.n18 10.6151
R1172 B.n713 B.n712 10.6151
R1173 B.n712 B.n711 10.6151
R1174 B.n711 B.n25 10.6151
R1175 B.n705 B.n25 10.6151
R1176 B.n705 B.n704 10.6151
R1177 B.n704 B.n703 10.6151
R1178 B.n703 B.n32 10.6151
R1179 B.n697 B.n32 10.6151
R1180 B.n697 B.n696 10.6151
R1181 B.n696 B.n695 10.6151
R1182 B.n99 B.n39 10.6151
R1183 B.n102 B.n99 10.6151
R1184 B.n103 B.n102 10.6151
R1185 B.n106 B.n103 10.6151
R1186 B.n107 B.n106 10.6151
R1187 B.n110 B.n107 10.6151
R1188 B.n111 B.n110 10.6151
R1189 B.n114 B.n111 10.6151
R1190 B.n115 B.n114 10.6151
R1191 B.n118 B.n115 10.6151
R1192 B.n119 B.n118 10.6151
R1193 B.n122 B.n119 10.6151
R1194 B.n123 B.n122 10.6151
R1195 B.n126 B.n123 10.6151
R1196 B.n127 B.n126 10.6151
R1197 B.n130 B.n127 10.6151
R1198 B.n131 B.n130 10.6151
R1199 B.n134 B.n131 10.6151
R1200 B.n135 B.n134 10.6151
R1201 B.n138 B.n135 10.6151
R1202 B.n139 B.n138 10.6151
R1203 B.n142 B.n139 10.6151
R1204 B.n143 B.n142 10.6151
R1205 B.n146 B.n143 10.6151
R1206 B.n147 B.n146 10.6151
R1207 B.n150 B.n147 10.6151
R1208 B.n151 B.n150 10.6151
R1209 B.n154 B.n151 10.6151
R1210 B.n155 B.n154 10.6151
R1211 B.n158 B.n155 10.6151
R1212 B.n159 B.n158 10.6151
R1213 B.n162 B.n159 10.6151
R1214 B.n163 B.n162 10.6151
R1215 B.n166 B.n163 10.6151
R1216 B.n167 B.n166 10.6151
R1217 B.n170 B.n167 10.6151
R1218 B.n171 B.n170 10.6151
R1219 B.n174 B.n171 10.6151
R1220 B.n175 B.n174 10.6151
R1221 B.n178 B.n175 10.6151
R1222 B.n179 B.n178 10.6151
R1223 B.n182 B.n179 10.6151
R1224 B.n183 B.n182 10.6151
R1225 B.n186 B.n183 10.6151
R1226 B.n187 B.n186 10.6151
R1227 B.n190 B.n187 10.6151
R1228 B.n195 B.n192 10.6151
R1229 B.n196 B.n195 10.6151
R1230 B.n199 B.n196 10.6151
R1231 B.n200 B.n199 10.6151
R1232 B.n203 B.n200 10.6151
R1233 B.n204 B.n203 10.6151
R1234 B.n207 B.n204 10.6151
R1235 B.n208 B.n207 10.6151
R1236 B.n212 B.n211 10.6151
R1237 B.n215 B.n212 10.6151
R1238 B.n216 B.n215 10.6151
R1239 B.n219 B.n216 10.6151
R1240 B.n220 B.n219 10.6151
R1241 B.n223 B.n220 10.6151
R1242 B.n224 B.n223 10.6151
R1243 B.n227 B.n224 10.6151
R1244 B.n228 B.n227 10.6151
R1245 B.n231 B.n228 10.6151
R1246 B.n232 B.n231 10.6151
R1247 B.n235 B.n232 10.6151
R1248 B.n236 B.n235 10.6151
R1249 B.n239 B.n236 10.6151
R1250 B.n240 B.n239 10.6151
R1251 B.n243 B.n240 10.6151
R1252 B.n244 B.n243 10.6151
R1253 B.n247 B.n244 10.6151
R1254 B.n248 B.n247 10.6151
R1255 B.n251 B.n248 10.6151
R1256 B.n252 B.n251 10.6151
R1257 B.n255 B.n252 10.6151
R1258 B.n256 B.n255 10.6151
R1259 B.n259 B.n256 10.6151
R1260 B.n260 B.n259 10.6151
R1261 B.n263 B.n260 10.6151
R1262 B.n264 B.n263 10.6151
R1263 B.n267 B.n264 10.6151
R1264 B.n268 B.n267 10.6151
R1265 B.n271 B.n268 10.6151
R1266 B.n272 B.n271 10.6151
R1267 B.n275 B.n272 10.6151
R1268 B.n276 B.n275 10.6151
R1269 B.n279 B.n276 10.6151
R1270 B.n280 B.n279 10.6151
R1271 B.n283 B.n280 10.6151
R1272 B.n284 B.n283 10.6151
R1273 B.n287 B.n284 10.6151
R1274 B.n288 B.n287 10.6151
R1275 B.n291 B.n288 10.6151
R1276 B.n292 B.n291 10.6151
R1277 B.n295 B.n292 10.6151
R1278 B.n296 B.n295 10.6151
R1279 B.n299 B.n296 10.6151
R1280 B.n300 B.n299 10.6151
R1281 B.n690 B.n300 10.6151
R1282 B.n644 B.t1 10.4353
R1283 B.t5 B.n723 10.4353
R1284 B.n737 B.n0 8.11757
R1285 B.n737 B.n1 8.11757
R1286 B.n318 B.t2 6.95702
R1287 B.t0 B.n716 6.95702
R1288 B.n485 B.n484 6.5566
R1289 B.n504 B.n503 6.5566
R1290 B.n192 B.n191 6.5566
R1291 B.n208 B.n96 6.5566
R1292 B.t7 B.n326 4.63818
R1293 B.t11 B.n30 4.63818
R1294 B.n484 B.n483 4.05904
R1295 B.n503 B.n362 4.05904
R1296 B.n191 B.n190 4.05904
R1297 B.n211 B.n96 4.05904
R1298 VN.n1 VN.t2 535.115
R1299 VN.n7 VN.t3 535.115
R1300 VN.n2 VN.t1 513.13
R1301 VN.n4 VN.t0 513.13
R1302 VN.n8 VN.t4 513.13
R1303 VN.n10 VN.t5 513.13
R1304 VN.n5 VN.n4 161.3
R1305 VN.n11 VN.n10 161.3
R1306 VN.n9 VN.n6 161.3
R1307 VN.n3 VN.n0 161.3
R1308 VN.n7 VN.n6 44.859
R1309 VN.n1 VN.n0 44.859
R1310 VN VN.n11 42.9683
R1311 VN.n4 VN.n3 27.752
R1312 VN.n10 VN.n9 27.752
R1313 VN.n3 VN.n2 20.449
R1314 VN.n9 VN.n8 20.449
R1315 VN.n2 VN.n1 19.9186
R1316 VN.n8 VN.n7 19.9186
R1317 VN.n11 VN.n6 0.189894
R1318 VN.n5 VN.n0 0.189894
R1319 VN VN.n5 0.0516364
R1320 VDD2.n1 VDD2.t3 65.8509
R1321 VDD2.n2 VDD2.t0 65.2275
R1322 VDD2.n1 VDD2.n0 63.953
R1323 VDD2 VDD2.n3 63.9502
R1324 VDD2.n2 VDD2.n1 38.4674
R1325 VDD2.n3 VDD2.t1 1.44576
R1326 VDD2.n3 VDD2.t2 1.44576
R1327 VDD2.n0 VDD2.t4 1.44576
R1328 VDD2.n0 VDD2.t5 1.44576
R1329 VDD2 VDD2.n2 0.737569
C0 VDD2 VDD1 0.717139f
C1 VTAIL VP 4.6157f
C2 VTAIL VN 4.601029f
C3 VDD1 VP 5.12305f
C4 VDD2 VP 0.299704f
C5 VDD1 VN 0.148303f
C6 VDD2 VN 4.97673f
C7 VDD1 VTAIL 10.9559f
C8 VDD2 VTAIL 10.989201f
C9 VN VP 5.41249f
C10 VDD2 B 4.805881f
C11 VDD1 B 5.039551f
C12 VTAIL B 7.029971f
C13 VN B 7.989849f
C14 VP B 5.940913f
C15 VDD2.t3 B 2.90639f
C16 VDD2.t4 B 0.252493f
C17 VDD2.t5 B 0.252493f
C18 VDD2.n0 B 2.27572f
C19 VDD2.n1 B 2.03775f
C20 VDD2.t0 B 2.90352f
C21 VDD2.n2 B 2.24673f
C22 VDD2.t1 B 0.252493f
C23 VDD2.t2 B 0.252493f
C24 VDD2.n3 B 2.2757f
C25 VN.n0 B 0.189904f
C26 VN.t2 B 1.29657f
C27 VN.n1 B 0.48218f
C28 VN.t1 B 1.2761f
C29 VN.n2 B 0.501857f
C30 VN.n3 B 0.010317f
C31 VN.t0 B 1.2761f
C32 VN.n4 B 0.495367f
C33 VN.n5 B 0.035234f
C34 VN.n6 B 0.189904f
C35 VN.t3 B 1.29657f
C36 VN.n7 B 0.48218f
C37 VN.t4 B 1.2761f
C38 VN.n8 B 0.501857f
C39 VN.n9 B 0.010317f
C40 VN.t5 B 1.2761f
C41 VN.n10 B 0.495367f
C42 VN.n11 B 1.95021f
C43 VTAIL.t4 B 0.260313f
C44 VTAIL.t5 B 0.260313f
C45 VTAIL.n0 B 2.27883f
C46 VTAIL.n1 B 0.3201f
C47 VTAIL.t8 B 2.90755f
C48 VTAIL.n2 B 0.449415f
C49 VTAIL.t7 B 0.260313f
C50 VTAIL.t10 B 0.260313f
C51 VTAIL.n3 B 2.27883f
C52 VTAIL.n4 B 1.67865f
C53 VTAIL.t2 B 0.260313f
C54 VTAIL.t1 B 0.260313f
C55 VTAIL.n5 B 2.27883f
C56 VTAIL.n6 B 1.67864f
C57 VTAIL.t3 B 2.90755f
C58 VTAIL.n7 B 0.449412f
C59 VTAIL.t6 B 0.260313f
C60 VTAIL.t11 B 0.260313f
C61 VTAIL.n8 B 2.27883f
C62 VTAIL.n9 B 0.368187f
C63 VTAIL.t9 B 2.90755f
C64 VTAIL.n10 B 1.68974f
C65 VTAIL.t0 B 2.90755f
C66 VTAIL.n11 B 1.6677f
C67 VDD1.t1 B 2.9095f
C68 VDD1.t0 B 2.9089f
C69 VDD1.t3 B 0.25271f
C70 VDD1.t5 B 0.25271f
C71 VDD1.n0 B 2.27768f
C72 VDD1.n1 B 2.11244f
C73 VDD1.t4 B 0.25271f
C74 VDD1.t2 B 0.25271f
C75 VDD1.n2 B 2.27693f
C76 VDD1.n3 B 2.22711f
C77 VP.n0 B 0.045965f
C78 VP.n1 B 0.01043f
C79 VP.n2 B 0.191988f
C80 VP.t2 B 1.29011f
C81 VP.t0 B 1.29011f
C82 VP.t5 B 1.3108f
C83 VP.n3 B 0.487472f
C84 VP.n4 B 0.507364f
C85 VP.n5 B 0.01043f
C86 VP.n6 B 0.500804f
C87 VP.n7 B 1.94147f
C88 VP.t4 B 1.29011f
C89 VP.n8 B 0.500804f
C90 VP.n9 B 1.98038f
C91 VP.n10 B 0.045965f
C92 VP.n11 B 0.045965f
C93 VP.t1 B 1.29011f
C94 VP.n12 B 0.503354f
C95 VP.n13 B 0.01043f
C96 VP.t3 B 1.29011f
C97 VP.n14 B 0.500804f
C98 VP.n15 B 0.035621f
.ends

