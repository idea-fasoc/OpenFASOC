* NGSPICE file created from diff_pair_sample_0975.ext - technology: sky130A

.subckt diff_pair_sample_0975 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t9 VN.t0 VTAIL.t17 B.t4 sky130_fd_pr__nfet_01v8 ad=1.482 pd=8.38 as=0.627 ps=4.13 w=3.8 l=3.44
X1 VTAIL.t10 VN.t1 VDD2.t8 B.t8 sky130_fd_pr__nfet_01v8 ad=0.627 pd=4.13 as=0.627 ps=4.13 w=3.8 l=3.44
X2 VDD1.t9 VP.t0 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=1.482 pd=8.38 as=0.627 ps=4.13 w=3.8 l=3.44
X3 VTAIL.t16 VN.t2 VDD2.t7 B.t0 sky130_fd_pr__nfet_01v8 ad=0.627 pd=4.13 as=0.627 ps=4.13 w=3.8 l=3.44
X4 B.t23 B.t21 B.t22 B.t18 sky130_fd_pr__nfet_01v8 ad=1.482 pd=8.38 as=0 ps=0 w=3.8 l=3.44
X5 VDD2.t6 VN.t3 VTAIL.t14 B.t7 sky130_fd_pr__nfet_01v8 ad=0.627 pd=4.13 as=1.482 ps=8.38 w=3.8 l=3.44
X6 VDD1.t8 VP.t1 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=0.627 pd=4.13 as=1.482 ps=8.38 w=3.8 l=3.44
X7 VTAIL.t0 VP.t2 VDD1.t7 B.t0 sky130_fd_pr__nfet_01v8 ad=0.627 pd=4.13 as=0.627 ps=4.13 w=3.8 l=3.44
X8 B.t20 B.t17 B.t19 B.t18 sky130_fd_pr__nfet_01v8 ad=1.482 pd=8.38 as=0 ps=0 w=3.8 l=3.44
X9 VDD2.t5 VN.t4 VTAIL.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=0.627 pd=4.13 as=0.627 ps=4.13 w=3.8 l=3.44
X10 VDD2.t4 VN.t5 VTAIL.t15 B.t6 sky130_fd_pr__nfet_01v8 ad=0.627 pd=4.13 as=0.627 ps=4.13 w=3.8 l=3.44
X11 VDD2.t3 VN.t6 VTAIL.t18 B.t1 sky130_fd_pr__nfet_01v8 ad=0.627 pd=4.13 as=1.482 ps=8.38 w=3.8 l=3.44
X12 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=1.482 pd=8.38 as=0 ps=0 w=3.8 l=3.44
X13 VDD2.t2 VN.t7 VTAIL.t19 B.t5 sky130_fd_pr__nfet_01v8 ad=1.482 pd=8.38 as=0.627 ps=4.13 w=3.8 l=3.44
X14 VDD1.t6 VP.t3 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=0.627 pd=4.13 as=0.627 ps=4.13 w=3.8 l=3.44
X15 VDD1.t5 VP.t4 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.482 pd=8.38 as=0.627 ps=4.13 w=3.8 l=3.44
X16 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=1.482 pd=8.38 as=0 ps=0 w=3.8 l=3.44
X17 VDD1.t4 VP.t5 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.627 pd=4.13 as=0.627 ps=4.13 w=3.8 l=3.44
X18 VTAIL.t2 VP.t6 VDD1.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=0.627 pd=4.13 as=0.627 ps=4.13 w=3.8 l=3.44
X19 VTAIL.t13 VN.t8 VDD2.t1 B.t9 sky130_fd_pr__nfet_01v8 ad=0.627 pd=4.13 as=0.627 ps=4.13 w=3.8 l=3.44
X20 VTAIL.t9 VP.t7 VDD1.t2 B.t9 sky130_fd_pr__nfet_01v8 ad=0.627 pd=4.13 as=0.627 ps=4.13 w=3.8 l=3.44
X21 VTAIL.t8 VP.t8 VDD1.t1 B.t8 sky130_fd_pr__nfet_01v8 ad=0.627 pd=4.13 as=0.627 ps=4.13 w=3.8 l=3.44
X22 VTAIL.t12 VN.t9 VDD2.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=0.627 pd=4.13 as=0.627 ps=4.13 w=3.8 l=3.44
X23 VDD1.t0 VP.t9 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.627 pd=4.13 as=1.482 ps=8.38 w=3.8 l=3.44
R0 VN.n102 VN.n101 161.3
R1 VN.n100 VN.n53 161.3
R2 VN.n99 VN.n98 161.3
R3 VN.n97 VN.n54 161.3
R4 VN.n96 VN.n95 161.3
R5 VN.n94 VN.n55 161.3
R6 VN.n93 VN.n92 161.3
R7 VN.n91 VN.n90 161.3
R8 VN.n89 VN.n57 161.3
R9 VN.n88 VN.n87 161.3
R10 VN.n86 VN.n58 161.3
R11 VN.n85 VN.n84 161.3
R12 VN.n83 VN.n59 161.3
R13 VN.n82 VN.n81 161.3
R14 VN.n80 VN.n60 161.3
R15 VN.n79 VN.n78 161.3
R16 VN.n77 VN.n61 161.3
R17 VN.n76 VN.n75 161.3
R18 VN.n74 VN.n63 161.3
R19 VN.n73 VN.n72 161.3
R20 VN.n71 VN.n64 161.3
R21 VN.n70 VN.n69 161.3
R22 VN.n68 VN.n65 161.3
R23 VN.n50 VN.n49 161.3
R24 VN.n48 VN.n1 161.3
R25 VN.n47 VN.n46 161.3
R26 VN.n45 VN.n2 161.3
R27 VN.n44 VN.n43 161.3
R28 VN.n42 VN.n3 161.3
R29 VN.n41 VN.n40 161.3
R30 VN.n39 VN.n38 161.3
R31 VN.n37 VN.n5 161.3
R32 VN.n36 VN.n35 161.3
R33 VN.n34 VN.n6 161.3
R34 VN.n33 VN.n32 161.3
R35 VN.n31 VN.n7 161.3
R36 VN.n30 VN.n29 161.3
R37 VN.n28 VN.n8 161.3
R38 VN.n27 VN.n26 161.3
R39 VN.n24 VN.n9 161.3
R40 VN.n23 VN.n22 161.3
R41 VN.n21 VN.n10 161.3
R42 VN.n20 VN.n19 161.3
R43 VN.n18 VN.n11 161.3
R44 VN.n17 VN.n16 161.3
R45 VN.n15 VN.n12 161.3
R46 VN.n51 VN.n0 75.9823
R47 VN.n103 VN.n52 75.9823
R48 VN.n14 VN.n13 73.9636
R49 VN.n67 VN.n66 73.9636
R50 VN.n67 VN.t6 59.4414
R51 VN.n14 VN.t7 59.4414
R52 VN.n19 VN.n10 53.6554
R53 VN.n32 VN.n6 53.6554
R54 VN.n72 VN.n63 53.6554
R55 VN.n84 VN.n58 53.6554
R56 VN VN.n103 51.7746
R57 VN.n43 VN.n2 49.7803
R58 VN.n95 VN.n54 49.7803
R59 VN.n47 VN.n2 31.3737
R60 VN.n99 VN.n54 31.3737
R61 VN.n23 VN.n10 27.4986
R62 VN.n32 VN.n31 27.4986
R63 VN.n76 VN.n63 27.4986
R64 VN.n84 VN.n83 27.4986
R65 VN.n13 VN.t2 26.6226
R66 VN.n25 VN.t4 26.6226
R67 VN.n4 VN.t1 26.6226
R68 VN.n0 VN.t3 26.6226
R69 VN.n66 VN.t9 26.6226
R70 VN.n62 VN.t5 26.6226
R71 VN.n56 VN.t8 26.6226
R72 VN.n52 VN.t0 26.6226
R73 VN.n17 VN.n12 24.5923
R74 VN.n18 VN.n17 24.5923
R75 VN.n19 VN.n18 24.5923
R76 VN.n24 VN.n23 24.5923
R77 VN.n26 VN.n24 24.5923
R78 VN.n30 VN.n8 24.5923
R79 VN.n31 VN.n30 24.5923
R80 VN.n36 VN.n6 24.5923
R81 VN.n37 VN.n36 24.5923
R82 VN.n38 VN.n37 24.5923
R83 VN.n42 VN.n41 24.5923
R84 VN.n43 VN.n42 24.5923
R85 VN.n48 VN.n47 24.5923
R86 VN.n49 VN.n48 24.5923
R87 VN.n72 VN.n71 24.5923
R88 VN.n71 VN.n70 24.5923
R89 VN.n70 VN.n65 24.5923
R90 VN.n83 VN.n82 24.5923
R91 VN.n82 VN.n60 24.5923
R92 VN.n78 VN.n77 24.5923
R93 VN.n77 VN.n76 24.5923
R94 VN.n95 VN.n94 24.5923
R95 VN.n94 VN.n93 24.5923
R96 VN.n90 VN.n89 24.5923
R97 VN.n89 VN.n88 24.5923
R98 VN.n88 VN.n58 24.5923
R99 VN.n101 VN.n100 24.5923
R100 VN.n100 VN.n99 24.5923
R101 VN.n41 VN.n4 23.6087
R102 VN.n93 VN.n56 23.6087
R103 VN.n49 VN.n0 14.2638
R104 VN.n101 VN.n52 14.2638
R105 VN.n26 VN.n25 12.2964
R106 VN.n25 VN.n8 12.2964
R107 VN.n62 VN.n60 12.2964
R108 VN.n78 VN.n62 12.2964
R109 VN.n68 VN.n67 4.18336
R110 VN.n15 VN.n14 4.18336
R111 VN.n13 VN.n12 0.984173
R112 VN.n38 VN.n4 0.984173
R113 VN.n66 VN.n65 0.984173
R114 VN.n90 VN.n56 0.984173
R115 VN.n103 VN.n102 0.354861
R116 VN.n51 VN.n50 0.354861
R117 VN VN.n51 0.267071
R118 VN.n102 VN.n53 0.189894
R119 VN.n98 VN.n53 0.189894
R120 VN.n98 VN.n97 0.189894
R121 VN.n97 VN.n96 0.189894
R122 VN.n96 VN.n55 0.189894
R123 VN.n92 VN.n55 0.189894
R124 VN.n92 VN.n91 0.189894
R125 VN.n91 VN.n57 0.189894
R126 VN.n87 VN.n57 0.189894
R127 VN.n87 VN.n86 0.189894
R128 VN.n86 VN.n85 0.189894
R129 VN.n85 VN.n59 0.189894
R130 VN.n81 VN.n59 0.189894
R131 VN.n81 VN.n80 0.189894
R132 VN.n80 VN.n79 0.189894
R133 VN.n79 VN.n61 0.189894
R134 VN.n75 VN.n61 0.189894
R135 VN.n75 VN.n74 0.189894
R136 VN.n74 VN.n73 0.189894
R137 VN.n73 VN.n64 0.189894
R138 VN.n69 VN.n64 0.189894
R139 VN.n69 VN.n68 0.189894
R140 VN.n16 VN.n15 0.189894
R141 VN.n16 VN.n11 0.189894
R142 VN.n20 VN.n11 0.189894
R143 VN.n21 VN.n20 0.189894
R144 VN.n22 VN.n21 0.189894
R145 VN.n22 VN.n9 0.189894
R146 VN.n27 VN.n9 0.189894
R147 VN.n28 VN.n27 0.189894
R148 VN.n29 VN.n28 0.189894
R149 VN.n29 VN.n7 0.189894
R150 VN.n33 VN.n7 0.189894
R151 VN.n34 VN.n33 0.189894
R152 VN.n35 VN.n34 0.189894
R153 VN.n35 VN.n5 0.189894
R154 VN.n39 VN.n5 0.189894
R155 VN.n40 VN.n39 0.189894
R156 VN.n40 VN.n3 0.189894
R157 VN.n44 VN.n3 0.189894
R158 VN.n45 VN.n44 0.189894
R159 VN.n46 VN.n45 0.189894
R160 VN.n46 VN.n1 0.189894
R161 VN.n50 VN.n1 0.189894
R162 VTAIL.n88 VTAIL.n74 289.615
R163 VTAIL.n16 VTAIL.n2 289.615
R164 VTAIL.n68 VTAIL.n54 289.615
R165 VTAIL.n44 VTAIL.n30 289.615
R166 VTAIL.n81 VTAIL.n80 185
R167 VTAIL.n78 VTAIL.n77 185
R168 VTAIL.n87 VTAIL.n86 185
R169 VTAIL.n89 VTAIL.n88 185
R170 VTAIL.n9 VTAIL.n8 185
R171 VTAIL.n6 VTAIL.n5 185
R172 VTAIL.n15 VTAIL.n14 185
R173 VTAIL.n17 VTAIL.n16 185
R174 VTAIL.n69 VTAIL.n68 185
R175 VTAIL.n67 VTAIL.n66 185
R176 VTAIL.n58 VTAIL.n57 185
R177 VTAIL.n61 VTAIL.n60 185
R178 VTAIL.n45 VTAIL.n44 185
R179 VTAIL.n43 VTAIL.n42 185
R180 VTAIL.n34 VTAIL.n33 185
R181 VTAIL.n37 VTAIL.n36 185
R182 VTAIL.t14 VTAIL.n79 147.888
R183 VTAIL.t1 VTAIL.n7 147.888
R184 VTAIL.t7 VTAIL.n59 147.888
R185 VTAIL.t18 VTAIL.n35 147.888
R186 VTAIL.n80 VTAIL.n77 104.615
R187 VTAIL.n87 VTAIL.n77 104.615
R188 VTAIL.n88 VTAIL.n87 104.615
R189 VTAIL.n8 VTAIL.n5 104.615
R190 VTAIL.n15 VTAIL.n5 104.615
R191 VTAIL.n16 VTAIL.n15 104.615
R192 VTAIL.n68 VTAIL.n67 104.615
R193 VTAIL.n67 VTAIL.n57 104.615
R194 VTAIL.n60 VTAIL.n57 104.615
R195 VTAIL.n44 VTAIL.n43 104.615
R196 VTAIL.n43 VTAIL.n33 104.615
R197 VTAIL.n36 VTAIL.n33 104.615
R198 VTAIL.n53 VTAIL.n52 56.0096
R199 VTAIL.n51 VTAIL.n50 56.0096
R200 VTAIL.n29 VTAIL.n28 56.0096
R201 VTAIL.n27 VTAIL.n26 56.0096
R202 VTAIL.n95 VTAIL.n94 56.0094
R203 VTAIL.n1 VTAIL.n0 56.0094
R204 VTAIL.n23 VTAIL.n22 56.0094
R205 VTAIL.n25 VTAIL.n24 56.0094
R206 VTAIL.n80 VTAIL.t14 52.3082
R207 VTAIL.n8 VTAIL.t1 52.3082
R208 VTAIL.n60 VTAIL.t7 52.3082
R209 VTAIL.n36 VTAIL.t18 52.3082
R210 VTAIL.n93 VTAIL.n92 31.4096
R211 VTAIL.n21 VTAIL.n20 31.4096
R212 VTAIL.n73 VTAIL.n72 31.4096
R213 VTAIL.n49 VTAIL.n48 31.4096
R214 VTAIL.n27 VTAIL.n25 22.1427
R215 VTAIL.n93 VTAIL.n73 18.8927
R216 VTAIL.n81 VTAIL.n79 15.6496
R217 VTAIL.n9 VTAIL.n7 15.6496
R218 VTAIL.n61 VTAIL.n59 15.6496
R219 VTAIL.n37 VTAIL.n35 15.6496
R220 VTAIL.n82 VTAIL.n78 12.8005
R221 VTAIL.n10 VTAIL.n6 12.8005
R222 VTAIL.n62 VTAIL.n58 12.8005
R223 VTAIL.n38 VTAIL.n34 12.8005
R224 VTAIL.n86 VTAIL.n85 12.0247
R225 VTAIL.n14 VTAIL.n13 12.0247
R226 VTAIL.n66 VTAIL.n65 12.0247
R227 VTAIL.n42 VTAIL.n41 12.0247
R228 VTAIL.n89 VTAIL.n76 11.249
R229 VTAIL.n17 VTAIL.n4 11.249
R230 VTAIL.n69 VTAIL.n56 11.249
R231 VTAIL.n45 VTAIL.n32 11.249
R232 VTAIL.n90 VTAIL.n74 10.4732
R233 VTAIL.n18 VTAIL.n2 10.4732
R234 VTAIL.n70 VTAIL.n54 10.4732
R235 VTAIL.n46 VTAIL.n30 10.4732
R236 VTAIL.n92 VTAIL.n91 9.45567
R237 VTAIL.n20 VTAIL.n19 9.45567
R238 VTAIL.n72 VTAIL.n71 9.45567
R239 VTAIL.n48 VTAIL.n47 9.45567
R240 VTAIL.n91 VTAIL.n90 9.3005
R241 VTAIL.n76 VTAIL.n75 9.3005
R242 VTAIL.n85 VTAIL.n84 9.3005
R243 VTAIL.n83 VTAIL.n82 9.3005
R244 VTAIL.n19 VTAIL.n18 9.3005
R245 VTAIL.n4 VTAIL.n3 9.3005
R246 VTAIL.n13 VTAIL.n12 9.3005
R247 VTAIL.n11 VTAIL.n10 9.3005
R248 VTAIL.n71 VTAIL.n70 9.3005
R249 VTAIL.n56 VTAIL.n55 9.3005
R250 VTAIL.n65 VTAIL.n64 9.3005
R251 VTAIL.n63 VTAIL.n62 9.3005
R252 VTAIL.n47 VTAIL.n46 9.3005
R253 VTAIL.n32 VTAIL.n31 9.3005
R254 VTAIL.n41 VTAIL.n40 9.3005
R255 VTAIL.n39 VTAIL.n38 9.3005
R256 VTAIL.n94 VTAIL.t11 5.21103
R257 VTAIL.n94 VTAIL.t10 5.21103
R258 VTAIL.n0 VTAIL.t19 5.21103
R259 VTAIL.n0 VTAIL.t16 5.21103
R260 VTAIL.n22 VTAIL.t6 5.21103
R261 VTAIL.n22 VTAIL.t2 5.21103
R262 VTAIL.n24 VTAIL.t4 5.21103
R263 VTAIL.n24 VTAIL.t9 5.21103
R264 VTAIL.n52 VTAIL.t3 5.21103
R265 VTAIL.n52 VTAIL.t8 5.21103
R266 VTAIL.n50 VTAIL.t5 5.21103
R267 VTAIL.n50 VTAIL.t0 5.21103
R268 VTAIL.n28 VTAIL.t15 5.21103
R269 VTAIL.n28 VTAIL.t12 5.21103
R270 VTAIL.n26 VTAIL.t17 5.21103
R271 VTAIL.n26 VTAIL.t13 5.21103
R272 VTAIL.n83 VTAIL.n79 4.40546
R273 VTAIL.n11 VTAIL.n7 4.40546
R274 VTAIL.n63 VTAIL.n59 4.40546
R275 VTAIL.n39 VTAIL.n35 4.40546
R276 VTAIL.n92 VTAIL.n74 3.49141
R277 VTAIL.n20 VTAIL.n2 3.49141
R278 VTAIL.n72 VTAIL.n54 3.49141
R279 VTAIL.n48 VTAIL.n30 3.49141
R280 VTAIL.n29 VTAIL.n27 3.2505
R281 VTAIL.n49 VTAIL.n29 3.2505
R282 VTAIL.n53 VTAIL.n51 3.2505
R283 VTAIL.n73 VTAIL.n53 3.2505
R284 VTAIL.n25 VTAIL.n23 3.2505
R285 VTAIL.n23 VTAIL.n21 3.2505
R286 VTAIL.n95 VTAIL.n93 3.2505
R287 VTAIL.n90 VTAIL.n89 2.71565
R288 VTAIL.n18 VTAIL.n17 2.71565
R289 VTAIL.n70 VTAIL.n69 2.71565
R290 VTAIL.n46 VTAIL.n45 2.71565
R291 VTAIL VTAIL.n1 2.49619
R292 VTAIL.n51 VTAIL.n49 2.09533
R293 VTAIL.n21 VTAIL.n1 2.09533
R294 VTAIL.n86 VTAIL.n76 1.93989
R295 VTAIL.n14 VTAIL.n4 1.93989
R296 VTAIL.n66 VTAIL.n56 1.93989
R297 VTAIL.n42 VTAIL.n32 1.93989
R298 VTAIL.n85 VTAIL.n78 1.16414
R299 VTAIL.n13 VTAIL.n6 1.16414
R300 VTAIL.n65 VTAIL.n58 1.16414
R301 VTAIL.n41 VTAIL.n34 1.16414
R302 VTAIL VTAIL.n95 0.75481
R303 VTAIL.n82 VTAIL.n81 0.388379
R304 VTAIL.n10 VTAIL.n9 0.388379
R305 VTAIL.n62 VTAIL.n61 0.388379
R306 VTAIL.n38 VTAIL.n37 0.388379
R307 VTAIL.n84 VTAIL.n83 0.155672
R308 VTAIL.n84 VTAIL.n75 0.155672
R309 VTAIL.n91 VTAIL.n75 0.155672
R310 VTAIL.n12 VTAIL.n11 0.155672
R311 VTAIL.n12 VTAIL.n3 0.155672
R312 VTAIL.n19 VTAIL.n3 0.155672
R313 VTAIL.n71 VTAIL.n55 0.155672
R314 VTAIL.n64 VTAIL.n55 0.155672
R315 VTAIL.n64 VTAIL.n63 0.155672
R316 VTAIL.n47 VTAIL.n31 0.155672
R317 VTAIL.n40 VTAIL.n31 0.155672
R318 VTAIL.n40 VTAIL.n39 0.155672
R319 VDD2.n37 VDD2.n23 289.615
R320 VDD2.n14 VDD2.n0 289.615
R321 VDD2.n38 VDD2.n37 185
R322 VDD2.n36 VDD2.n35 185
R323 VDD2.n27 VDD2.n26 185
R324 VDD2.n30 VDD2.n29 185
R325 VDD2.n7 VDD2.n6 185
R326 VDD2.n4 VDD2.n3 185
R327 VDD2.n13 VDD2.n12 185
R328 VDD2.n15 VDD2.n14 185
R329 VDD2.t9 VDD2.n28 147.888
R330 VDD2.t2 VDD2.n5 147.888
R331 VDD2.n37 VDD2.n36 104.615
R332 VDD2.n36 VDD2.n26 104.615
R333 VDD2.n29 VDD2.n26 104.615
R334 VDD2.n6 VDD2.n3 104.615
R335 VDD2.n13 VDD2.n3 104.615
R336 VDD2.n14 VDD2.n13 104.615
R337 VDD2.n22 VDD2.n21 75.0704
R338 VDD2 VDD2.n45 75.0675
R339 VDD2.n44 VDD2.n43 72.6883
R340 VDD2.n20 VDD2.n19 72.6882
R341 VDD2.n29 VDD2.t9 52.3082
R342 VDD2.n6 VDD2.t2 52.3082
R343 VDD2.n20 VDD2.n18 51.3384
R344 VDD2.n42 VDD2.n41 48.0884
R345 VDD2.n42 VDD2.n22 42.4287
R346 VDD2.n30 VDD2.n28 15.6496
R347 VDD2.n7 VDD2.n5 15.6496
R348 VDD2.n31 VDD2.n27 12.8005
R349 VDD2.n8 VDD2.n4 12.8005
R350 VDD2.n35 VDD2.n34 12.0247
R351 VDD2.n12 VDD2.n11 12.0247
R352 VDD2.n38 VDD2.n25 11.249
R353 VDD2.n15 VDD2.n2 11.249
R354 VDD2.n39 VDD2.n23 10.4732
R355 VDD2.n16 VDD2.n0 10.4732
R356 VDD2.n41 VDD2.n40 9.45567
R357 VDD2.n18 VDD2.n17 9.45567
R358 VDD2.n40 VDD2.n39 9.3005
R359 VDD2.n25 VDD2.n24 9.3005
R360 VDD2.n34 VDD2.n33 9.3005
R361 VDD2.n32 VDD2.n31 9.3005
R362 VDD2.n17 VDD2.n16 9.3005
R363 VDD2.n2 VDD2.n1 9.3005
R364 VDD2.n11 VDD2.n10 9.3005
R365 VDD2.n9 VDD2.n8 9.3005
R366 VDD2.n45 VDD2.t0 5.21103
R367 VDD2.n45 VDD2.t3 5.21103
R368 VDD2.n43 VDD2.t1 5.21103
R369 VDD2.n43 VDD2.t4 5.21103
R370 VDD2.n21 VDD2.t8 5.21103
R371 VDD2.n21 VDD2.t6 5.21103
R372 VDD2.n19 VDD2.t7 5.21103
R373 VDD2.n19 VDD2.t5 5.21103
R374 VDD2.n32 VDD2.n28 4.40546
R375 VDD2.n9 VDD2.n5 4.40546
R376 VDD2.n41 VDD2.n23 3.49141
R377 VDD2.n18 VDD2.n0 3.49141
R378 VDD2.n44 VDD2.n42 3.2505
R379 VDD2.n39 VDD2.n38 2.71565
R380 VDD2.n16 VDD2.n15 2.71565
R381 VDD2.n35 VDD2.n25 1.93989
R382 VDD2.n12 VDD2.n2 1.93989
R383 VDD2.n34 VDD2.n27 1.16414
R384 VDD2.n11 VDD2.n4 1.16414
R385 VDD2 VDD2.n44 0.87119
R386 VDD2.n22 VDD2.n20 0.757654
R387 VDD2.n31 VDD2.n30 0.388379
R388 VDD2.n8 VDD2.n7 0.388379
R389 VDD2.n40 VDD2.n24 0.155672
R390 VDD2.n33 VDD2.n24 0.155672
R391 VDD2.n33 VDD2.n32 0.155672
R392 VDD2.n10 VDD2.n9 0.155672
R393 VDD2.n10 VDD2.n1 0.155672
R394 VDD2.n17 VDD2.n1 0.155672
R395 B.n743 B.n742 585
R396 B.n743 B.n134 585
R397 B.n746 B.n745 585
R398 B.n747 B.n161 585
R399 B.n749 B.n748 585
R400 B.n751 B.n160 585
R401 B.n754 B.n753 585
R402 B.n755 B.n159 585
R403 B.n757 B.n756 585
R404 B.n759 B.n158 585
R405 B.n762 B.n761 585
R406 B.n763 B.n157 585
R407 B.n765 B.n764 585
R408 B.n767 B.n156 585
R409 B.n770 B.n769 585
R410 B.n771 B.n155 585
R411 B.n773 B.n772 585
R412 B.n775 B.n154 585
R413 B.n778 B.n777 585
R414 B.n780 B.n151 585
R415 B.n782 B.n781 585
R416 B.n784 B.n150 585
R417 B.n787 B.n786 585
R418 B.n788 B.n149 585
R419 B.n790 B.n789 585
R420 B.n792 B.n148 585
R421 B.n794 B.n793 585
R422 B.n796 B.n795 585
R423 B.n799 B.n798 585
R424 B.n800 B.n143 585
R425 B.n802 B.n801 585
R426 B.n804 B.n142 585
R427 B.n807 B.n806 585
R428 B.n808 B.n141 585
R429 B.n810 B.n809 585
R430 B.n812 B.n140 585
R431 B.n815 B.n814 585
R432 B.n816 B.n139 585
R433 B.n818 B.n817 585
R434 B.n820 B.n138 585
R435 B.n823 B.n822 585
R436 B.n824 B.n137 585
R437 B.n826 B.n825 585
R438 B.n828 B.n136 585
R439 B.n831 B.n830 585
R440 B.n832 B.n135 585
R441 B.n741 B.n133 585
R442 B.n835 B.n133 585
R443 B.n740 B.n132 585
R444 B.n836 B.n132 585
R445 B.n739 B.n131 585
R446 B.n837 B.n131 585
R447 B.n738 B.n737 585
R448 B.n737 B.n127 585
R449 B.n736 B.n126 585
R450 B.n843 B.n126 585
R451 B.n735 B.n125 585
R452 B.n844 B.n125 585
R453 B.n734 B.n124 585
R454 B.n845 B.n124 585
R455 B.n733 B.n732 585
R456 B.n732 B.n120 585
R457 B.n731 B.n119 585
R458 B.n851 B.n119 585
R459 B.n730 B.n118 585
R460 B.n852 B.n118 585
R461 B.n729 B.n117 585
R462 B.n853 B.n117 585
R463 B.n728 B.n727 585
R464 B.n727 B.n113 585
R465 B.n726 B.n112 585
R466 B.n859 B.n112 585
R467 B.n725 B.n111 585
R468 B.n860 B.n111 585
R469 B.n724 B.n110 585
R470 B.n861 B.n110 585
R471 B.n723 B.n722 585
R472 B.n722 B.n106 585
R473 B.n721 B.n105 585
R474 B.n867 B.n105 585
R475 B.n720 B.n104 585
R476 B.n868 B.n104 585
R477 B.n719 B.n103 585
R478 B.n869 B.n103 585
R479 B.n718 B.n717 585
R480 B.n717 B.n99 585
R481 B.n716 B.n98 585
R482 B.n875 B.n98 585
R483 B.n715 B.n97 585
R484 B.n876 B.n97 585
R485 B.n714 B.n96 585
R486 B.n877 B.n96 585
R487 B.n713 B.n712 585
R488 B.n712 B.t7 585
R489 B.n711 B.n92 585
R490 B.n883 B.n92 585
R491 B.n710 B.n91 585
R492 B.n884 B.n91 585
R493 B.n709 B.n90 585
R494 B.n885 B.n90 585
R495 B.n708 B.n707 585
R496 B.n707 B.n86 585
R497 B.n706 B.n85 585
R498 B.n891 B.n85 585
R499 B.n705 B.n84 585
R500 B.n892 B.n84 585
R501 B.n704 B.n83 585
R502 B.n893 B.n83 585
R503 B.n703 B.n702 585
R504 B.n702 B.n79 585
R505 B.n701 B.n78 585
R506 B.n899 B.n78 585
R507 B.n700 B.n77 585
R508 B.n900 B.n77 585
R509 B.n699 B.n76 585
R510 B.n901 B.n76 585
R511 B.n698 B.n697 585
R512 B.n697 B.n72 585
R513 B.n696 B.n71 585
R514 B.n907 B.n71 585
R515 B.n695 B.n70 585
R516 B.n908 B.n70 585
R517 B.n694 B.n69 585
R518 B.n909 B.n69 585
R519 B.n693 B.n692 585
R520 B.n692 B.n65 585
R521 B.n691 B.n64 585
R522 B.n915 B.n64 585
R523 B.n690 B.n63 585
R524 B.n916 B.n63 585
R525 B.n689 B.n62 585
R526 B.n917 B.n62 585
R527 B.n688 B.n687 585
R528 B.n687 B.n58 585
R529 B.n686 B.n57 585
R530 B.n923 B.n57 585
R531 B.n685 B.n56 585
R532 B.n924 B.n56 585
R533 B.n684 B.n55 585
R534 B.n925 B.n55 585
R535 B.n683 B.n682 585
R536 B.n682 B.n51 585
R537 B.n681 B.n50 585
R538 B.n931 B.n50 585
R539 B.n680 B.n49 585
R540 B.n932 B.n49 585
R541 B.n679 B.n48 585
R542 B.n933 B.n48 585
R543 B.n678 B.n677 585
R544 B.n677 B.n44 585
R545 B.n676 B.n43 585
R546 B.n939 B.n43 585
R547 B.n675 B.n42 585
R548 B.n940 B.n42 585
R549 B.n674 B.n41 585
R550 B.n941 B.n41 585
R551 B.n673 B.n672 585
R552 B.n672 B.n37 585
R553 B.n671 B.n36 585
R554 B.n947 B.n36 585
R555 B.n670 B.n35 585
R556 B.n948 B.n35 585
R557 B.n669 B.n34 585
R558 B.n949 B.n34 585
R559 B.n668 B.n667 585
R560 B.n667 B.n30 585
R561 B.n666 B.n29 585
R562 B.n955 B.n29 585
R563 B.n665 B.n28 585
R564 B.n956 B.n28 585
R565 B.n664 B.n27 585
R566 B.n957 B.n27 585
R567 B.n663 B.n662 585
R568 B.n662 B.n23 585
R569 B.n661 B.n22 585
R570 B.n963 B.n22 585
R571 B.n660 B.n21 585
R572 B.n964 B.n21 585
R573 B.n659 B.n20 585
R574 B.n965 B.n20 585
R575 B.n658 B.n657 585
R576 B.n657 B.n19 585
R577 B.n656 B.n15 585
R578 B.n971 B.n15 585
R579 B.n655 B.n14 585
R580 B.n972 B.n14 585
R581 B.n654 B.n13 585
R582 B.n973 B.n13 585
R583 B.n653 B.n652 585
R584 B.n652 B.n12 585
R585 B.n651 B.n650 585
R586 B.n651 B.n8 585
R587 B.n649 B.n7 585
R588 B.n980 B.n7 585
R589 B.n648 B.n6 585
R590 B.n981 B.n6 585
R591 B.n647 B.n5 585
R592 B.n982 B.n5 585
R593 B.n646 B.n645 585
R594 B.n645 B.n4 585
R595 B.n644 B.n162 585
R596 B.n644 B.n643 585
R597 B.n634 B.n163 585
R598 B.n164 B.n163 585
R599 B.n636 B.n635 585
R600 B.n637 B.n636 585
R601 B.n633 B.n169 585
R602 B.n169 B.n168 585
R603 B.n632 B.n631 585
R604 B.n631 B.n630 585
R605 B.n171 B.n170 585
R606 B.n623 B.n171 585
R607 B.n622 B.n621 585
R608 B.n624 B.n622 585
R609 B.n620 B.n176 585
R610 B.n176 B.n175 585
R611 B.n619 B.n618 585
R612 B.n618 B.n617 585
R613 B.n178 B.n177 585
R614 B.n179 B.n178 585
R615 B.n610 B.n609 585
R616 B.n611 B.n610 585
R617 B.n608 B.n184 585
R618 B.n184 B.n183 585
R619 B.n607 B.n606 585
R620 B.n606 B.n605 585
R621 B.n186 B.n185 585
R622 B.n187 B.n186 585
R623 B.n598 B.n597 585
R624 B.n599 B.n598 585
R625 B.n596 B.n192 585
R626 B.n192 B.n191 585
R627 B.n595 B.n594 585
R628 B.n594 B.n593 585
R629 B.n194 B.n193 585
R630 B.n195 B.n194 585
R631 B.n586 B.n585 585
R632 B.n587 B.n586 585
R633 B.n584 B.n200 585
R634 B.n200 B.n199 585
R635 B.n583 B.n582 585
R636 B.n582 B.n581 585
R637 B.n202 B.n201 585
R638 B.n203 B.n202 585
R639 B.n574 B.n573 585
R640 B.n575 B.n574 585
R641 B.n572 B.n208 585
R642 B.n208 B.n207 585
R643 B.n571 B.n570 585
R644 B.n570 B.n569 585
R645 B.n210 B.n209 585
R646 B.n211 B.n210 585
R647 B.n562 B.n561 585
R648 B.n563 B.n562 585
R649 B.n560 B.n215 585
R650 B.n219 B.n215 585
R651 B.n559 B.n558 585
R652 B.n558 B.n557 585
R653 B.n217 B.n216 585
R654 B.n218 B.n217 585
R655 B.n550 B.n549 585
R656 B.n551 B.n550 585
R657 B.n548 B.n224 585
R658 B.n224 B.n223 585
R659 B.n547 B.n546 585
R660 B.n546 B.n545 585
R661 B.n226 B.n225 585
R662 B.n227 B.n226 585
R663 B.n538 B.n537 585
R664 B.n539 B.n538 585
R665 B.n536 B.n232 585
R666 B.n232 B.n231 585
R667 B.n535 B.n534 585
R668 B.n534 B.n533 585
R669 B.n234 B.n233 585
R670 B.n235 B.n234 585
R671 B.n526 B.n525 585
R672 B.n527 B.n526 585
R673 B.n524 B.n240 585
R674 B.n240 B.n239 585
R675 B.n523 B.n522 585
R676 B.n522 B.n521 585
R677 B.n242 B.n241 585
R678 B.n243 B.n242 585
R679 B.n514 B.n513 585
R680 B.n515 B.n514 585
R681 B.n512 B.n248 585
R682 B.n248 B.n247 585
R683 B.n511 B.n510 585
R684 B.n510 B.n509 585
R685 B.n250 B.n249 585
R686 B.n251 B.n250 585
R687 B.n502 B.n501 585
R688 B.n503 B.n502 585
R689 B.n500 B.n256 585
R690 B.n256 B.n255 585
R691 B.n499 B.n498 585
R692 B.n498 B.n497 585
R693 B.n258 B.n257 585
R694 B.t4 B.n258 585
R695 B.n490 B.n489 585
R696 B.n491 B.n490 585
R697 B.n488 B.n263 585
R698 B.n263 B.n262 585
R699 B.n487 B.n486 585
R700 B.n486 B.n485 585
R701 B.n265 B.n264 585
R702 B.n266 B.n265 585
R703 B.n478 B.n477 585
R704 B.n479 B.n478 585
R705 B.n476 B.n271 585
R706 B.n271 B.n270 585
R707 B.n475 B.n474 585
R708 B.n474 B.n473 585
R709 B.n273 B.n272 585
R710 B.n274 B.n273 585
R711 B.n466 B.n465 585
R712 B.n467 B.n466 585
R713 B.n464 B.n279 585
R714 B.n279 B.n278 585
R715 B.n463 B.n462 585
R716 B.n462 B.n461 585
R717 B.n281 B.n280 585
R718 B.n282 B.n281 585
R719 B.n454 B.n453 585
R720 B.n455 B.n454 585
R721 B.n452 B.n287 585
R722 B.n287 B.n286 585
R723 B.n451 B.n450 585
R724 B.n450 B.n449 585
R725 B.n289 B.n288 585
R726 B.n290 B.n289 585
R727 B.n442 B.n441 585
R728 B.n443 B.n442 585
R729 B.n440 B.n295 585
R730 B.n295 B.n294 585
R731 B.n439 B.n438 585
R732 B.n438 B.n437 585
R733 B.n297 B.n296 585
R734 B.n298 B.n297 585
R735 B.n430 B.n429 585
R736 B.n431 B.n430 585
R737 B.n428 B.n303 585
R738 B.n303 B.n302 585
R739 B.n427 B.n426 585
R740 B.n426 B.n425 585
R741 B.n422 B.n307 585
R742 B.n421 B.n420 585
R743 B.n418 B.n308 585
R744 B.n418 B.n306 585
R745 B.n417 B.n416 585
R746 B.n415 B.n414 585
R747 B.n413 B.n310 585
R748 B.n411 B.n410 585
R749 B.n409 B.n311 585
R750 B.n408 B.n407 585
R751 B.n405 B.n312 585
R752 B.n403 B.n402 585
R753 B.n401 B.n313 585
R754 B.n400 B.n399 585
R755 B.n397 B.n314 585
R756 B.n395 B.n394 585
R757 B.n393 B.n315 585
R758 B.n392 B.n391 585
R759 B.n389 B.n316 585
R760 B.n387 B.n386 585
R761 B.n385 B.n317 585
R762 B.n384 B.n383 585
R763 B.n381 B.n321 585
R764 B.n379 B.n378 585
R765 B.n377 B.n322 585
R766 B.n376 B.n375 585
R767 B.n373 B.n323 585
R768 B.n371 B.n370 585
R769 B.n368 B.n324 585
R770 B.n367 B.n366 585
R771 B.n364 B.n327 585
R772 B.n362 B.n361 585
R773 B.n360 B.n328 585
R774 B.n359 B.n358 585
R775 B.n356 B.n329 585
R776 B.n354 B.n353 585
R777 B.n352 B.n330 585
R778 B.n351 B.n350 585
R779 B.n348 B.n331 585
R780 B.n346 B.n345 585
R781 B.n344 B.n332 585
R782 B.n343 B.n342 585
R783 B.n340 B.n333 585
R784 B.n338 B.n337 585
R785 B.n336 B.n335 585
R786 B.n305 B.n304 585
R787 B.n424 B.n423 585
R788 B.n425 B.n424 585
R789 B.n301 B.n300 585
R790 B.n302 B.n301 585
R791 B.n433 B.n432 585
R792 B.n432 B.n431 585
R793 B.n434 B.n299 585
R794 B.n299 B.n298 585
R795 B.n436 B.n435 585
R796 B.n437 B.n436 585
R797 B.n293 B.n292 585
R798 B.n294 B.n293 585
R799 B.n445 B.n444 585
R800 B.n444 B.n443 585
R801 B.n446 B.n291 585
R802 B.n291 B.n290 585
R803 B.n448 B.n447 585
R804 B.n449 B.n448 585
R805 B.n285 B.n284 585
R806 B.n286 B.n285 585
R807 B.n457 B.n456 585
R808 B.n456 B.n455 585
R809 B.n458 B.n283 585
R810 B.n283 B.n282 585
R811 B.n460 B.n459 585
R812 B.n461 B.n460 585
R813 B.n277 B.n276 585
R814 B.n278 B.n277 585
R815 B.n469 B.n468 585
R816 B.n468 B.n467 585
R817 B.n470 B.n275 585
R818 B.n275 B.n274 585
R819 B.n472 B.n471 585
R820 B.n473 B.n472 585
R821 B.n269 B.n268 585
R822 B.n270 B.n269 585
R823 B.n481 B.n480 585
R824 B.n480 B.n479 585
R825 B.n482 B.n267 585
R826 B.n267 B.n266 585
R827 B.n484 B.n483 585
R828 B.n485 B.n484 585
R829 B.n261 B.n260 585
R830 B.n262 B.n261 585
R831 B.n493 B.n492 585
R832 B.n492 B.n491 585
R833 B.n494 B.n259 585
R834 B.n259 B.t4 585
R835 B.n496 B.n495 585
R836 B.n497 B.n496 585
R837 B.n254 B.n253 585
R838 B.n255 B.n254 585
R839 B.n505 B.n504 585
R840 B.n504 B.n503 585
R841 B.n506 B.n252 585
R842 B.n252 B.n251 585
R843 B.n508 B.n507 585
R844 B.n509 B.n508 585
R845 B.n246 B.n245 585
R846 B.n247 B.n246 585
R847 B.n517 B.n516 585
R848 B.n516 B.n515 585
R849 B.n518 B.n244 585
R850 B.n244 B.n243 585
R851 B.n520 B.n519 585
R852 B.n521 B.n520 585
R853 B.n238 B.n237 585
R854 B.n239 B.n238 585
R855 B.n529 B.n528 585
R856 B.n528 B.n527 585
R857 B.n530 B.n236 585
R858 B.n236 B.n235 585
R859 B.n532 B.n531 585
R860 B.n533 B.n532 585
R861 B.n230 B.n229 585
R862 B.n231 B.n230 585
R863 B.n541 B.n540 585
R864 B.n540 B.n539 585
R865 B.n542 B.n228 585
R866 B.n228 B.n227 585
R867 B.n544 B.n543 585
R868 B.n545 B.n544 585
R869 B.n222 B.n221 585
R870 B.n223 B.n222 585
R871 B.n553 B.n552 585
R872 B.n552 B.n551 585
R873 B.n554 B.n220 585
R874 B.n220 B.n218 585
R875 B.n556 B.n555 585
R876 B.n557 B.n556 585
R877 B.n214 B.n213 585
R878 B.n219 B.n214 585
R879 B.n565 B.n564 585
R880 B.n564 B.n563 585
R881 B.n566 B.n212 585
R882 B.n212 B.n211 585
R883 B.n568 B.n567 585
R884 B.n569 B.n568 585
R885 B.n206 B.n205 585
R886 B.n207 B.n206 585
R887 B.n577 B.n576 585
R888 B.n576 B.n575 585
R889 B.n578 B.n204 585
R890 B.n204 B.n203 585
R891 B.n580 B.n579 585
R892 B.n581 B.n580 585
R893 B.n198 B.n197 585
R894 B.n199 B.n198 585
R895 B.n589 B.n588 585
R896 B.n588 B.n587 585
R897 B.n590 B.n196 585
R898 B.n196 B.n195 585
R899 B.n592 B.n591 585
R900 B.n593 B.n592 585
R901 B.n190 B.n189 585
R902 B.n191 B.n190 585
R903 B.n601 B.n600 585
R904 B.n600 B.n599 585
R905 B.n602 B.n188 585
R906 B.n188 B.n187 585
R907 B.n604 B.n603 585
R908 B.n605 B.n604 585
R909 B.n182 B.n181 585
R910 B.n183 B.n182 585
R911 B.n613 B.n612 585
R912 B.n612 B.n611 585
R913 B.n614 B.n180 585
R914 B.n180 B.n179 585
R915 B.n616 B.n615 585
R916 B.n617 B.n616 585
R917 B.n174 B.n173 585
R918 B.n175 B.n174 585
R919 B.n626 B.n625 585
R920 B.n625 B.n624 585
R921 B.n627 B.n172 585
R922 B.n623 B.n172 585
R923 B.n629 B.n628 585
R924 B.n630 B.n629 585
R925 B.n167 B.n166 585
R926 B.n168 B.n167 585
R927 B.n639 B.n638 585
R928 B.n638 B.n637 585
R929 B.n640 B.n165 585
R930 B.n165 B.n164 585
R931 B.n642 B.n641 585
R932 B.n643 B.n642 585
R933 B.n3 B.n0 585
R934 B.n4 B.n3 585
R935 B.n979 B.n1 585
R936 B.n980 B.n979 585
R937 B.n978 B.n977 585
R938 B.n978 B.n8 585
R939 B.n976 B.n9 585
R940 B.n12 B.n9 585
R941 B.n975 B.n974 585
R942 B.n974 B.n973 585
R943 B.n11 B.n10 585
R944 B.n972 B.n11 585
R945 B.n970 B.n969 585
R946 B.n971 B.n970 585
R947 B.n968 B.n16 585
R948 B.n19 B.n16 585
R949 B.n967 B.n966 585
R950 B.n966 B.n965 585
R951 B.n18 B.n17 585
R952 B.n964 B.n18 585
R953 B.n962 B.n961 585
R954 B.n963 B.n962 585
R955 B.n960 B.n24 585
R956 B.n24 B.n23 585
R957 B.n959 B.n958 585
R958 B.n958 B.n957 585
R959 B.n26 B.n25 585
R960 B.n956 B.n26 585
R961 B.n954 B.n953 585
R962 B.n955 B.n954 585
R963 B.n952 B.n31 585
R964 B.n31 B.n30 585
R965 B.n951 B.n950 585
R966 B.n950 B.n949 585
R967 B.n33 B.n32 585
R968 B.n948 B.n33 585
R969 B.n946 B.n945 585
R970 B.n947 B.n946 585
R971 B.n944 B.n38 585
R972 B.n38 B.n37 585
R973 B.n943 B.n942 585
R974 B.n942 B.n941 585
R975 B.n40 B.n39 585
R976 B.n940 B.n40 585
R977 B.n938 B.n937 585
R978 B.n939 B.n938 585
R979 B.n936 B.n45 585
R980 B.n45 B.n44 585
R981 B.n935 B.n934 585
R982 B.n934 B.n933 585
R983 B.n47 B.n46 585
R984 B.n932 B.n47 585
R985 B.n930 B.n929 585
R986 B.n931 B.n930 585
R987 B.n928 B.n52 585
R988 B.n52 B.n51 585
R989 B.n927 B.n926 585
R990 B.n926 B.n925 585
R991 B.n54 B.n53 585
R992 B.n924 B.n54 585
R993 B.n922 B.n921 585
R994 B.n923 B.n922 585
R995 B.n920 B.n59 585
R996 B.n59 B.n58 585
R997 B.n919 B.n918 585
R998 B.n918 B.n917 585
R999 B.n61 B.n60 585
R1000 B.n916 B.n61 585
R1001 B.n914 B.n913 585
R1002 B.n915 B.n914 585
R1003 B.n912 B.n66 585
R1004 B.n66 B.n65 585
R1005 B.n911 B.n910 585
R1006 B.n910 B.n909 585
R1007 B.n68 B.n67 585
R1008 B.n908 B.n68 585
R1009 B.n906 B.n905 585
R1010 B.n907 B.n906 585
R1011 B.n904 B.n73 585
R1012 B.n73 B.n72 585
R1013 B.n903 B.n902 585
R1014 B.n902 B.n901 585
R1015 B.n75 B.n74 585
R1016 B.n900 B.n75 585
R1017 B.n898 B.n897 585
R1018 B.n899 B.n898 585
R1019 B.n896 B.n80 585
R1020 B.n80 B.n79 585
R1021 B.n895 B.n894 585
R1022 B.n894 B.n893 585
R1023 B.n82 B.n81 585
R1024 B.n892 B.n82 585
R1025 B.n890 B.n889 585
R1026 B.n891 B.n890 585
R1027 B.n888 B.n87 585
R1028 B.n87 B.n86 585
R1029 B.n887 B.n886 585
R1030 B.n886 B.n885 585
R1031 B.n89 B.n88 585
R1032 B.n884 B.n89 585
R1033 B.n882 B.n881 585
R1034 B.n883 B.n882 585
R1035 B.n880 B.n93 585
R1036 B.n93 B.t7 585
R1037 B.n879 B.n878 585
R1038 B.n878 B.n877 585
R1039 B.n95 B.n94 585
R1040 B.n876 B.n95 585
R1041 B.n874 B.n873 585
R1042 B.n875 B.n874 585
R1043 B.n872 B.n100 585
R1044 B.n100 B.n99 585
R1045 B.n871 B.n870 585
R1046 B.n870 B.n869 585
R1047 B.n102 B.n101 585
R1048 B.n868 B.n102 585
R1049 B.n866 B.n865 585
R1050 B.n867 B.n866 585
R1051 B.n864 B.n107 585
R1052 B.n107 B.n106 585
R1053 B.n863 B.n862 585
R1054 B.n862 B.n861 585
R1055 B.n109 B.n108 585
R1056 B.n860 B.n109 585
R1057 B.n858 B.n857 585
R1058 B.n859 B.n858 585
R1059 B.n856 B.n114 585
R1060 B.n114 B.n113 585
R1061 B.n855 B.n854 585
R1062 B.n854 B.n853 585
R1063 B.n116 B.n115 585
R1064 B.n852 B.n116 585
R1065 B.n850 B.n849 585
R1066 B.n851 B.n850 585
R1067 B.n848 B.n121 585
R1068 B.n121 B.n120 585
R1069 B.n847 B.n846 585
R1070 B.n846 B.n845 585
R1071 B.n123 B.n122 585
R1072 B.n844 B.n123 585
R1073 B.n842 B.n841 585
R1074 B.n843 B.n842 585
R1075 B.n840 B.n128 585
R1076 B.n128 B.n127 585
R1077 B.n839 B.n838 585
R1078 B.n838 B.n837 585
R1079 B.n130 B.n129 585
R1080 B.n836 B.n130 585
R1081 B.n834 B.n833 585
R1082 B.n835 B.n834 585
R1083 B.n983 B.n982 585
R1084 B.n981 B.n2 585
R1085 B.n834 B.n135 487.695
R1086 B.n743 B.n133 487.695
R1087 B.n426 B.n305 487.695
R1088 B.n424 B.n307 487.695
R1089 B.n744 B.n134 256.663
R1090 B.n750 B.n134 256.663
R1091 B.n752 B.n134 256.663
R1092 B.n758 B.n134 256.663
R1093 B.n760 B.n134 256.663
R1094 B.n766 B.n134 256.663
R1095 B.n768 B.n134 256.663
R1096 B.n774 B.n134 256.663
R1097 B.n776 B.n134 256.663
R1098 B.n783 B.n134 256.663
R1099 B.n785 B.n134 256.663
R1100 B.n791 B.n134 256.663
R1101 B.n147 B.n134 256.663
R1102 B.n797 B.n134 256.663
R1103 B.n803 B.n134 256.663
R1104 B.n805 B.n134 256.663
R1105 B.n811 B.n134 256.663
R1106 B.n813 B.n134 256.663
R1107 B.n819 B.n134 256.663
R1108 B.n821 B.n134 256.663
R1109 B.n827 B.n134 256.663
R1110 B.n829 B.n134 256.663
R1111 B.n419 B.n306 256.663
R1112 B.n309 B.n306 256.663
R1113 B.n412 B.n306 256.663
R1114 B.n406 B.n306 256.663
R1115 B.n404 B.n306 256.663
R1116 B.n398 B.n306 256.663
R1117 B.n396 B.n306 256.663
R1118 B.n390 B.n306 256.663
R1119 B.n388 B.n306 256.663
R1120 B.n382 B.n306 256.663
R1121 B.n380 B.n306 256.663
R1122 B.n374 B.n306 256.663
R1123 B.n372 B.n306 256.663
R1124 B.n365 B.n306 256.663
R1125 B.n363 B.n306 256.663
R1126 B.n357 B.n306 256.663
R1127 B.n355 B.n306 256.663
R1128 B.n349 B.n306 256.663
R1129 B.n347 B.n306 256.663
R1130 B.n341 B.n306 256.663
R1131 B.n339 B.n306 256.663
R1132 B.n334 B.n306 256.663
R1133 B.n985 B.n984 256.663
R1134 B.n144 B.t21 235.661
R1135 B.n152 B.t17 235.661
R1136 B.n325 B.t14 235.661
R1137 B.n318 B.t10 235.661
R1138 B.n152 B.t19 214.496
R1139 B.n325 B.t16 214.496
R1140 B.n144 B.t22 214.496
R1141 B.n318 B.t13 214.496
R1142 B.n830 B.n828 163.367
R1143 B.n826 B.n137 163.367
R1144 B.n822 B.n820 163.367
R1145 B.n818 B.n139 163.367
R1146 B.n814 B.n812 163.367
R1147 B.n810 B.n141 163.367
R1148 B.n806 B.n804 163.367
R1149 B.n802 B.n143 163.367
R1150 B.n798 B.n796 163.367
R1151 B.n793 B.n792 163.367
R1152 B.n790 B.n149 163.367
R1153 B.n786 B.n784 163.367
R1154 B.n782 B.n151 163.367
R1155 B.n777 B.n775 163.367
R1156 B.n773 B.n155 163.367
R1157 B.n769 B.n767 163.367
R1158 B.n765 B.n157 163.367
R1159 B.n761 B.n759 163.367
R1160 B.n757 B.n159 163.367
R1161 B.n753 B.n751 163.367
R1162 B.n749 B.n161 163.367
R1163 B.n745 B.n743 163.367
R1164 B.n426 B.n303 163.367
R1165 B.n430 B.n303 163.367
R1166 B.n430 B.n297 163.367
R1167 B.n438 B.n297 163.367
R1168 B.n438 B.n295 163.367
R1169 B.n442 B.n295 163.367
R1170 B.n442 B.n289 163.367
R1171 B.n450 B.n289 163.367
R1172 B.n450 B.n287 163.367
R1173 B.n454 B.n287 163.367
R1174 B.n454 B.n281 163.367
R1175 B.n462 B.n281 163.367
R1176 B.n462 B.n279 163.367
R1177 B.n466 B.n279 163.367
R1178 B.n466 B.n273 163.367
R1179 B.n474 B.n273 163.367
R1180 B.n474 B.n271 163.367
R1181 B.n478 B.n271 163.367
R1182 B.n478 B.n265 163.367
R1183 B.n486 B.n265 163.367
R1184 B.n486 B.n263 163.367
R1185 B.n490 B.n263 163.367
R1186 B.n490 B.n258 163.367
R1187 B.n498 B.n258 163.367
R1188 B.n498 B.n256 163.367
R1189 B.n502 B.n256 163.367
R1190 B.n502 B.n250 163.367
R1191 B.n510 B.n250 163.367
R1192 B.n510 B.n248 163.367
R1193 B.n514 B.n248 163.367
R1194 B.n514 B.n242 163.367
R1195 B.n522 B.n242 163.367
R1196 B.n522 B.n240 163.367
R1197 B.n526 B.n240 163.367
R1198 B.n526 B.n234 163.367
R1199 B.n534 B.n234 163.367
R1200 B.n534 B.n232 163.367
R1201 B.n538 B.n232 163.367
R1202 B.n538 B.n226 163.367
R1203 B.n546 B.n226 163.367
R1204 B.n546 B.n224 163.367
R1205 B.n550 B.n224 163.367
R1206 B.n550 B.n217 163.367
R1207 B.n558 B.n217 163.367
R1208 B.n558 B.n215 163.367
R1209 B.n562 B.n215 163.367
R1210 B.n562 B.n210 163.367
R1211 B.n570 B.n210 163.367
R1212 B.n570 B.n208 163.367
R1213 B.n574 B.n208 163.367
R1214 B.n574 B.n202 163.367
R1215 B.n582 B.n202 163.367
R1216 B.n582 B.n200 163.367
R1217 B.n586 B.n200 163.367
R1218 B.n586 B.n194 163.367
R1219 B.n594 B.n194 163.367
R1220 B.n594 B.n192 163.367
R1221 B.n598 B.n192 163.367
R1222 B.n598 B.n186 163.367
R1223 B.n606 B.n186 163.367
R1224 B.n606 B.n184 163.367
R1225 B.n610 B.n184 163.367
R1226 B.n610 B.n178 163.367
R1227 B.n618 B.n178 163.367
R1228 B.n618 B.n176 163.367
R1229 B.n622 B.n176 163.367
R1230 B.n622 B.n171 163.367
R1231 B.n631 B.n171 163.367
R1232 B.n631 B.n169 163.367
R1233 B.n636 B.n169 163.367
R1234 B.n636 B.n163 163.367
R1235 B.n644 B.n163 163.367
R1236 B.n645 B.n644 163.367
R1237 B.n645 B.n5 163.367
R1238 B.n6 B.n5 163.367
R1239 B.n7 B.n6 163.367
R1240 B.n651 B.n7 163.367
R1241 B.n652 B.n651 163.367
R1242 B.n652 B.n13 163.367
R1243 B.n14 B.n13 163.367
R1244 B.n15 B.n14 163.367
R1245 B.n657 B.n15 163.367
R1246 B.n657 B.n20 163.367
R1247 B.n21 B.n20 163.367
R1248 B.n22 B.n21 163.367
R1249 B.n662 B.n22 163.367
R1250 B.n662 B.n27 163.367
R1251 B.n28 B.n27 163.367
R1252 B.n29 B.n28 163.367
R1253 B.n667 B.n29 163.367
R1254 B.n667 B.n34 163.367
R1255 B.n35 B.n34 163.367
R1256 B.n36 B.n35 163.367
R1257 B.n672 B.n36 163.367
R1258 B.n672 B.n41 163.367
R1259 B.n42 B.n41 163.367
R1260 B.n43 B.n42 163.367
R1261 B.n677 B.n43 163.367
R1262 B.n677 B.n48 163.367
R1263 B.n49 B.n48 163.367
R1264 B.n50 B.n49 163.367
R1265 B.n682 B.n50 163.367
R1266 B.n682 B.n55 163.367
R1267 B.n56 B.n55 163.367
R1268 B.n57 B.n56 163.367
R1269 B.n687 B.n57 163.367
R1270 B.n687 B.n62 163.367
R1271 B.n63 B.n62 163.367
R1272 B.n64 B.n63 163.367
R1273 B.n692 B.n64 163.367
R1274 B.n692 B.n69 163.367
R1275 B.n70 B.n69 163.367
R1276 B.n71 B.n70 163.367
R1277 B.n697 B.n71 163.367
R1278 B.n697 B.n76 163.367
R1279 B.n77 B.n76 163.367
R1280 B.n78 B.n77 163.367
R1281 B.n702 B.n78 163.367
R1282 B.n702 B.n83 163.367
R1283 B.n84 B.n83 163.367
R1284 B.n85 B.n84 163.367
R1285 B.n707 B.n85 163.367
R1286 B.n707 B.n90 163.367
R1287 B.n91 B.n90 163.367
R1288 B.n92 B.n91 163.367
R1289 B.n712 B.n92 163.367
R1290 B.n712 B.n96 163.367
R1291 B.n97 B.n96 163.367
R1292 B.n98 B.n97 163.367
R1293 B.n717 B.n98 163.367
R1294 B.n717 B.n103 163.367
R1295 B.n104 B.n103 163.367
R1296 B.n105 B.n104 163.367
R1297 B.n722 B.n105 163.367
R1298 B.n722 B.n110 163.367
R1299 B.n111 B.n110 163.367
R1300 B.n112 B.n111 163.367
R1301 B.n727 B.n112 163.367
R1302 B.n727 B.n117 163.367
R1303 B.n118 B.n117 163.367
R1304 B.n119 B.n118 163.367
R1305 B.n732 B.n119 163.367
R1306 B.n732 B.n124 163.367
R1307 B.n125 B.n124 163.367
R1308 B.n126 B.n125 163.367
R1309 B.n737 B.n126 163.367
R1310 B.n737 B.n131 163.367
R1311 B.n132 B.n131 163.367
R1312 B.n133 B.n132 163.367
R1313 B.n420 B.n418 163.367
R1314 B.n418 B.n417 163.367
R1315 B.n414 B.n413 163.367
R1316 B.n411 B.n311 163.367
R1317 B.n407 B.n405 163.367
R1318 B.n403 B.n313 163.367
R1319 B.n399 B.n397 163.367
R1320 B.n395 B.n315 163.367
R1321 B.n391 B.n389 163.367
R1322 B.n387 B.n317 163.367
R1323 B.n383 B.n381 163.367
R1324 B.n379 B.n322 163.367
R1325 B.n375 B.n373 163.367
R1326 B.n371 B.n324 163.367
R1327 B.n366 B.n364 163.367
R1328 B.n362 B.n328 163.367
R1329 B.n358 B.n356 163.367
R1330 B.n354 B.n330 163.367
R1331 B.n350 B.n348 163.367
R1332 B.n346 B.n332 163.367
R1333 B.n342 B.n340 163.367
R1334 B.n338 B.n335 163.367
R1335 B.n424 B.n301 163.367
R1336 B.n432 B.n301 163.367
R1337 B.n432 B.n299 163.367
R1338 B.n436 B.n299 163.367
R1339 B.n436 B.n293 163.367
R1340 B.n444 B.n293 163.367
R1341 B.n444 B.n291 163.367
R1342 B.n448 B.n291 163.367
R1343 B.n448 B.n285 163.367
R1344 B.n456 B.n285 163.367
R1345 B.n456 B.n283 163.367
R1346 B.n460 B.n283 163.367
R1347 B.n460 B.n277 163.367
R1348 B.n468 B.n277 163.367
R1349 B.n468 B.n275 163.367
R1350 B.n472 B.n275 163.367
R1351 B.n472 B.n269 163.367
R1352 B.n480 B.n269 163.367
R1353 B.n480 B.n267 163.367
R1354 B.n484 B.n267 163.367
R1355 B.n484 B.n261 163.367
R1356 B.n492 B.n261 163.367
R1357 B.n492 B.n259 163.367
R1358 B.n496 B.n259 163.367
R1359 B.n496 B.n254 163.367
R1360 B.n504 B.n254 163.367
R1361 B.n504 B.n252 163.367
R1362 B.n508 B.n252 163.367
R1363 B.n508 B.n246 163.367
R1364 B.n516 B.n246 163.367
R1365 B.n516 B.n244 163.367
R1366 B.n520 B.n244 163.367
R1367 B.n520 B.n238 163.367
R1368 B.n528 B.n238 163.367
R1369 B.n528 B.n236 163.367
R1370 B.n532 B.n236 163.367
R1371 B.n532 B.n230 163.367
R1372 B.n540 B.n230 163.367
R1373 B.n540 B.n228 163.367
R1374 B.n544 B.n228 163.367
R1375 B.n544 B.n222 163.367
R1376 B.n552 B.n222 163.367
R1377 B.n552 B.n220 163.367
R1378 B.n556 B.n220 163.367
R1379 B.n556 B.n214 163.367
R1380 B.n564 B.n214 163.367
R1381 B.n564 B.n212 163.367
R1382 B.n568 B.n212 163.367
R1383 B.n568 B.n206 163.367
R1384 B.n576 B.n206 163.367
R1385 B.n576 B.n204 163.367
R1386 B.n580 B.n204 163.367
R1387 B.n580 B.n198 163.367
R1388 B.n588 B.n198 163.367
R1389 B.n588 B.n196 163.367
R1390 B.n592 B.n196 163.367
R1391 B.n592 B.n190 163.367
R1392 B.n600 B.n190 163.367
R1393 B.n600 B.n188 163.367
R1394 B.n604 B.n188 163.367
R1395 B.n604 B.n182 163.367
R1396 B.n612 B.n182 163.367
R1397 B.n612 B.n180 163.367
R1398 B.n616 B.n180 163.367
R1399 B.n616 B.n174 163.367
R1400 B.n625 B.n174 163.367
R1401 B.n625 B.n172 163.367
R1402 B.n629 B.n172 163.367
R1403 B.n629 B.n167 163.367
R1404 B.n638 B.n167 163.367
R1405 B.n638 B.n165 163.367
R1406 B.n642 B.n165 163.367
R1407 B.n642 B.n3 163.367
R1408 B.n983 B.n3 163.367
R1409 B.n979 B.n2 163.367
R1410 B.n979 B.n978 163.367
R1411 B.n978 B.n9 163.367
R1412 B.n974 B.n9 163.367
R1413 B.n974 B.n11 163.367
R1414 B.n970 B.n11 163.367
R1415 B.n970 B.n16 163.367
R1416 B.n966 B.n16 163.367
R1417 B.n966 B.n18 163.367
R1418 B.n962 B.n18 163.367
R1419 B.n962 B.n24 163.367
R1420 B.n958 B.n24 163.367
R1421 B.n958 B.n26 163.367
R1422 B.n954 B.n26 163.367
R1423 B.n954 B.n31 163.367
R1424 B.n950 B.n31 163.367
R1425 B.n950 B.n33 163.367
R1426 B.n946 B.n33 163.367
R1427 B.n946 B.n38 163.367
R1428 B.n942 B.n38 163.367
R1429 B.n942 B.n40 163.367
R1430 B.n938 B.n40 163.367
R1431 B.n938 B.n45 163.367
R1432 B.n934 B.n45 163.367
R1433 B.n934 B.n47 163.367
R1434 B.n930 B.n47 163.367
R1435 B.n930 B.n52 163.367
R1436 B.n926 B.n52 163.367
R1437 B.n926 B.n54 163.367
R1438 B.n922 B.n54 163.367
R1439 B.n922 B.n59 163.367
R1440 B.n918 B.n59 163.367
R1441 B.n918 B.n61 163.367
R1442 B.n914 B.n61 163.367
R1443 B.n914 B.n66 163.367
R1444 B.n910 B.n66 163.367
R1445 B.n910 B.n68 163.367
R1446 B.n906 B.n68 163.367
R1447 B.n906 B.n73 163.367
R1448 B.n902 B.n73 163.367
R1449 B.n902 B.n75 163.367
R1450 B.n898 B.n75 163.367
R1451 B.n898 B.n80 163.367
R1452 B.n894 B.n80 163.367
R1453 B.n894 B.n82 163.367
R1454 B.n890 B.n82 163.367
R1455 B.n890 B.n87 163.367
R1456 B.n886 B.n87 163.367
R1457 B.n886 B.n89 163.367
R1458 B.n882 B.n89 163.367
R1459 B.n882 B.n93 163.367
R1460 B.n878 B.n93 163.367
R1461 B.n878 B.n95 163.367
R1462 B.n874 B.n95 163.367
R1463 B.n874 B.n100 163.367
R1464 B.n870 B.n100 163.367
R1465 B.n870 B.n102 163.367
R1466 B.n866 B.n102 163.367
R1467 B.n866 B.n107 163.367
R1468 B.n862 B.n107 163.367
R1469 B.n862 B.n109 163.367
R1470 B.n858 B.n109 163.367
R1471 B.n858 B.n114 163.367
R1472 B.n854 B.n114 163.367
R1473 B.n854 B.n116 163.367
R1474 B.n850 B.n116 163.367
R1475 B.n850 B.n121 163.367
R1476 B.n846 B.n121 163.367
R1477 B.n846 B.n123 163.367
R1478 B.n842 B.n123 163.367
R1479 B.n842 B.n128 163.367
R1480 B.n838 B.n128 163.367
R1481 B.n838 B.n130 163.367
R1482 B.n834 B.n130 163.367
R1483 B.n425 B.n306 161.213
R1484 B.n835 B.n134 161.213
R1485 B.n153 B.t20 141.381
R1486 B.n326 B.t15 141.381
R1487 B.n145 B.t23 141.381
R1488 B.n319 B.t12 141.381
R1489 B.n425 B.n302 82.4247
R1490 B.n431 B.n302 82.4247
R1491 B.n431 B.n298 82.4247
R1492 B.n437 B.n298 82.4247
R1493 B.n437 B.n294 82.4247
R1494 B.n443 B.n294 82.4247
R1495 B.n443 B.n290 82.4247
R1496 B.n449 B.n290 82.4247
R1497 B.n455 B.n286 82.4247
R1498 B.n455 B.n282 82.4247
R1499 B.n461 B.n282 82.4247
R1500 B.n461 B.n278 82.4247
R1501 B.n467 B.n278 82.4247
R1502 B.n467 B.n274 82.4247
R1503 B.n473 B.n274 82.4247
R1504 B.n473 B.n270 82.4247
R1505 B.n479 B.n270 82.4247
R1506 B.n479 B.n266 82.4247
R1507 B.n485 B.n266 82.4247
R1508 B.n485 B.n262 82.4247
R1509 B.n491 B.n262 82.4247
R1510 B.n491 B.t4 82.4247
R1511 B.n497 B.t4 82.4247
R1512 B.n497 B.n255 82.4247
R1513 B.n503 B.n255 82.4247
R1514 B.n503 B.n251 82.4247
R1515 B.n509 B.n251 82.4247
R1516 B.n509 B.n247 82.4247
R1517 B.n515 B.n247 82.4247
R1518 B.n515 B.n243 82.4247
R1519 B.n521 B.n243 82.4247
R1520 B.n521 B.n239 82.4247
R1521 B.n527 B.n239 82.4247
R1522 B.n533 B.n235 82.4247
R1523 B.n533 B.n231 82.4247
R1524 B.n539 B.n231 82.4247
R1525 B.n539 B.n227 82.4247
R1526 B.n545 B.n227 82.4247
R1527 B.n545 B.n223 82.4247
R1528 B.n551 B.n223 82.4247
R1529 B.n551 B.n218 82.4247
R1530 B.n557 B.n218 82.4247
R1531 B.n557 B.n219 82.4247
R1532 B.n563 B.n211 82.4247
R1533 B.n569 B.n211 82.4247
R1534 B.n569 B.n207 82.4247
R1535 B.n575 B.n207 82.4247
R1536 B.n575 B.n203 82.4247
R1537 B.n581 B.n203 82.4247
R1538 B.n581 B.n199 82.4247
R1539 B.n587 B.n199 82.4247
R1540 B.n587 B.n195 82.4247
R1541 B.n593 B.n195 82.4247
R1542 B.n599 B.n191 82.4247
R1543 B.n599 B.n187 82.4247
R1544 B.n605 B.n187 82.4247
R1545 B.n605 B.n183 82.4247
R1546 B.n611 B.n183 82.4247
R1547 B.n611 B.n179 82.4247
R1548 B.n617 B.n179 82.4247
R1549 B.n617 B.n175 82.4247
R1550 B.n624 B.n175 82.4247
R1551 B.n624 B.n623 82.4247
R1552 B.n630 B.n168 82.4247
R1553 B.n637 B.n168 82.4247
R1554 B.n637 B.n164 82.4247
R1555 B.n643 B.n164 82.4247
R1556 B.n643 B.n4 82.4247
R1557 B.n982 B.n4 82.4247
R1558 B.n982 B.n981 82.4247
R1559 B.n981 B.n980 82.4247
R1560 B.n980 B.n8 82.4247
R1561 B.n12 B.n8 82.4247
R1562 B.n973 B.n12 82.4247
R1563 B.n973 B.n972 82.4247
R1564 B.n972 B.n971 82.4247
R1565 B.n965 B.n19 82.4247
R1566 B.n965 B.n964 82.4247
R1567 B.n964 B.n963 82.4247
R1568 B.n963 B.n23 82.4247
R1569 B.n957 B.n23 82.4247
R1570 B.n957 B.n956 82.4247
R1571 B.n956 B.n955 82.4247
R1572 B.n955 B.n30 82.4247
R1573 B.n949 B.n30 82.4247
R1574 B.n949 B.n948 82.4247
R1575 B.n947 B.n37 82.4247
R1576 B.n941 B.n37 82.4247
R1577 B.n941 B.n940 82.4247
R1578 B.n940 B.n939 82.4247
R1579 B.n939 B.n44 82.4247
R1580 B.n933 B.n44 82.4247
R1581 B.n933 B.n932 82.4247
R1582 B.n932 B.n931 82.4247
R1583 B.n931 B.n51 82.4247
R1584 B.n925 B.n51 82.4247
R1585 B.n924 B.n923 82.4247
R1586 B.n923 B.n58 82.4247
R1587 B.n917 B.n58 82.4247
R1588 B.n917 B.n916 82.4247
R1589 B.n916 B.n915 82.4247
R1590 B.n915 B.n65 82.4247
R1591 B.n909 B.n65 82.4247
R1592 B.n909 B.n908 82.4247
R1593 B.n908 B.n907 82.4247
R1594 B.n907 B.n72 82.4247
R1595 B.n901 B.n900 82.4247
R1596 B.n900 B.n899 82.4247
R1597 B.n899 B.n79 82.4247
R1598 B.n893 B.n79 82.4247
R1599 B.n893 B.n892 82.4247
R1600 B.n892 B.n891 82.4247
R1601 B.n891 B.n86 82.4247
R1602 B.n885 B.n86 82.4247
R1603 B.n885 B.n884 82.4247
R1604 B.n884 B.n883 82.4247
R1605 B.n883 B.t7 82.4247
R1606 B.n877 B.t7 82.4247
R1607 B.n877 B.n876 82.4247
R1608 B.n876 B.n875 82.4247
R1609 B.n875 B.n99 82.4247
R1610 B.n869 B.n99 82.4247
R1611 B.n869 B.n868 82.4247
R1612 B.n868 B.n867 82.4247
R1613 B.n867 B.n106 82.4247
R1614 B.n861 B.n106 82.4247
R1615 B.n861 B.n860 82.4247
R1616 B.n860 B.n859 82.4247
R1617 B.n859 B.n113 82.4247
R1618 B.n853 B.n113 82.4247
R1619 B.n853 B.n852 82.4247
R1620 B.n851 B.n120 82.4247
R1621 B.n845 B.n120 82.4247
R1622 B.n845 B.n844 82.4247
R1623 B.n844 B.n843 82.4247
R1624 B.n843 B.n127 82.4247
R1625 B.n837 B.n127 82.4247
R1626 B.n837 B.n836 82.4247
R1627 B.n836 B.n835 82.4247
R1628 B.t9 B.n235 75.152
R1629 B.t8 B.n72 75.152
R1630 B.n145 B.n144 73.1157
R1631 B.n153 B.n152 73.1157
R1632 B.n326 B.n325 73.1157
R1633 B.n319 B.n318 73.1157
R1634 B.n829 B.n135 71.676
R1635 B.n828 B.n827 71.676
R1636 B.n821 B.n137 71.676
R1637 B.n820 B.n819 71.676
R1638 B.n813 B.n139 71.676
R1639 B.n812 B.n811 71.676
R1640 B.n805 B.n141 71.676
R1641 B.n804 B.n803 71.676
R1642 B.n797 B.n143 71.676
R1643 B.n796 B.n147 71.676
R1644 B.n792 B.n791 71.676
R1645 B.n785 B.n149 71.676
R1646 B.n784 B.n783 71.676
R1647 B.n776 B.n151 71.676
R1648 B.n775 B.n774 71.676
R1649 B.n768 B.n155 71.676
R1650 B.n767 B.n766 71.676
R1651 B.n760 B.n157 71.676
R1652 B.n759 B.n758 71.676
R1653 B.n752 B.n159 71.676
R1654 B.n751 B.n750 71.676
R1655 B.n744 B.n161 71.676
R1656 B.n745 B.n744 71.676
R1657 B.n750 B.n749 71.676
R1658 B.n753 B.n752 71.676
R1659 B.n758 B.n757 71.676
R1660 B.n761 B.n760 71.676
R1661 B.n766 B.n765 71.676
R1662 B.n769 B.n768 71.676
R1663 B.n774 B.n773 71.676
R1664 B.n777 B.n776 71.676
R1665 B.n783 B.n782 71.676
R1666 B.n786 B.n785 71.676
R1667 B.n791 B.n790 71.676
R1668 B.n793 B.n147 71.676
R1669 B.n798 B.n797 71.676
R1670 B.n803 B.n802 71.676
R1671 B.n806 B.n805 71.676
R1672 B.n811 B.n810 71.676
R1673 B.n814 B.n813 71.676
R1674 B.n819 B.n818 71.676
R1675 B.n822 B.n821 71.676
R1676 B.n827 B.n826 71.676
R1677 B.n830 B.n829 71.676
R1678 B.n419 B.n307 71.676
R1679 B.n417 B.n309 71.676
R1680 B.n413 B.n412 71.676
R1681 B.n406 B.n311 71.676
R1682 B.n405 B.n404 71.676
R1683 B.n398 B.n313 71.676
R1684 B.n397 B.n396 71.676
R1685 B.n390 B.n315 71.676
R1686 B.n389 B.n388 71.676
R1687 B.n382 B.n317 71.676
R1688 B.n381 B.n380 71.676
R1689 B.n374 B.n322 71.676
R1690 B.n373 B.n372 71.676
R1691 B.n365 B.n324 71.676
R1692 B.n364 B.n363 71.676
R1693 B.n357 B.n328 71.676
R1694 B.n356 B.n355 71.676
R1695 B.n349 B.n330 71.676
R1696 B.n348 B.n347 71.676
R1697 B.n341 B.n332 71.676
R1698 B.n340 B.n339 71.676
R1699 B.n335 B.n334 71.676
R1700 B.n420 B.n419 71.676
R1701 B.n414 B.n309 71.676
R1702 B.n412 B.n411 71.676
R1703 B.n407 B.n406 71.676
R1704 B.n404 B.n403 71.676
R1705 B.n399 B.n398 71.676
R1706 B.n396 B.n395 71.676
R1707 B.n391 B.n390 71.676
R1708 B.n388 B.n387 71.676
R1709 B.n383 B.n382 71.676
R1710 B.n380 B.n379 71.676
R1711 B.n375 B.n374 71.676
R1712 B.n372 B.n371 71.676
R1713 B.n366 B.n365 71.676
R1714 B.n363 B.n362 71.676
R1715 B.n358 B.n357 71.676
R1716 B.n355 B.n354 71.676
R1717 B.n350 B.n349 71.676
R1718 B.n347 B.n346 71.676
R1719 B.n342 B.n341 71.676
R1720 B.n339 B.n338 71.676
R1721 B.n334 B.n305 71.676
R1722 B.n984 B.n983 71.676
R1723 B.n984 B.n2 71.676
R1724 B.n563 B.t6 67.8793
R1725 B.n925 B.t3 67.8793
R1726 B.t2 B.n191 60.6066
R1727 B.n948 B.t0 60.6066
R1728 B.n146 B.n145 59.5399
R1729 B.n779 B.n153 59.5399
R1730 B.n369 B.n326 59.5399
R1731 B.n320 B.n319 59.5399
R1732 B.n449 B.t11 58.1823
R1733 B.t18 B.n851 58.1823
R1734 B.n630 B.t1 53.3338
R1735 B.n971 B.t5 53.3338
R1736 B.n423 B.n422 31.6883
R1737 B.n427 B.n304 31.6883
R1738 B.n742 B.n741 31.6883
R1739 B.n833 B.n832 31.6883
R1740 B.n623 B.t1 29.0914
R1741 B.n19 B.t5 29.0914
R1742 B.t11 B.n286 24.2429
R1743 B.n852 B.t18 24.2429
R1744 B.n593 B.t2 21.8187
R1745 B.t0 B.n947 21.8187
R1746 B B.n985 18.0485
R1747 B.n219 B.t6 14.546
R1748 B.t3 B.n924 14.546
R1749 B.n423 B.n300 10.6151
R1750 B.n433 B.n300 10.6151
R1751 B.n434 B.n433 10.6151
R1752 B.n435 B.n434 10.6151
R1753 B.n435 B.n292 10.6151
R1754 B.n445 B.n292 10.6151
R1755 B.n446 B.n445 10.6151
R1756 B.n447 B.n446 10.6151
R1757 B.n447 B.n284 10.6151
R1758 B.n457 B.n284 10.6151
R1759 B.n458 B.n457 10.6151
R1760 B.n459 B.n458 10.6151
R1761 B.n459 B.n276 10.6151
R1762 B.n469 B.n276 10.6151
R1763 B.n470 B.n469 10.6151
R1764 B.n471 B.n470 10.6151
R1765 B.n471 B.n268 10.6151
R1766 B.n481 B.n268 10.6151
R1767 B.n482 B.n481 10.6151
R1768 B.n483 B.n482 10.6151
R1769 B.n483 B.n260 10.6151
R1770 B.n493 B.n260 10.6151
R1771 B.n494 B.n493 10.6151
R1772 B.n495 B.n494 10.6151
R1773 B.n495 B.n253 10.6151
R1774 B.n505 B.n253 10.6151
R1775 B.n506 B.n505 10.6151
R1776 B.n507 B.n506 10.6151
R1777 B.n507 B.n245 10.6151
R1778 B.n517 B.n245 10.6151
R1779 B.n518 B.n517 10.6151
R1780 B.n519 B.n518 10.6151
R1781 B.n519 B.n237 10.6151
R1782 B.n529 B.n237 10.6151
R1783 B.n530 B.n529 10.6151
R1784 B.n531 B.n530 10.6151
R1785 B.n531 B.n229 10.6151
R1786 B.n541 B.n229 10.6151
R1787 B.n542 B.n541 10.6151
R1788 B.n543 B.n542 10.6151
R1789 B.n543 B.n221 10.6151
R1790 B.n553 B.n221 10.6151
R1791 B.n554 B.n553 10.6151
R1792 B.n555 B.n554 10.6151
R1793 B.n555 B.n213 10.6151
R1794 B.n565 B.n213 10.6151
R1795 B.n566 B.n565 10.6151
R1796 B.n567 B.n566 10.6151
R1797 B.n567 B.n205 10.6151
R1798 B.n577 B.n205 10.6151
R1799 B.n578 B.n577 10.6151
R1800 B.n579 B.n578 10.6151
R1801 B.n579 B.n197 10.6151
R1802 B.n589 B.n197 10.6151
R1803 B.n590 B.n589 10.6151
R1804 B.n591 B.n590 10.6151
R1805 B.n591 B.n189 10.6151
R1806 B.n601 B.n189 10.6151
R1807 B.n602 B.n601 10.6151
R1808 B.n603 B.n602 10.6151
R1809 B.n603 B.n181 10.6151
R1810 B.n613 B.n181 10.6151
R1811 B.n614 B.n613 10.6151
R1812 B.n615 B.n614 10.6151
R1813 B.n615 B.n173 10.6151
R1814 B.n626 B.n173 10.6151
R1815 B.n627 B.n626 10.6151
R1816 B.n628 B.n627 10.6151
R1817 B.n628 B.n166 10.6151
R1818 B.n639 B.n166 10.6151
R1819 B.n640 B.n639 10.6151
R1820 B.n641 B.n640 10.6151
R1821 B.n641 B.n0 10.6151
R1822 B.n422 B.n421 10.6151
R1823 B.n421 B.n308 10.6151
R1824 B.n416 B.n308 10.6151
R1825 B.n416 B.n415 10.6151
R1826 B.n415 B.n310 10.6151
R1827 B.n410 B.n310 10.6151
R1828 B.n410 B.n409 10.6151
R1829 B.n409 B.n408 10.6151
R1830 B.n408 B.n312 10.6151
R1831 B.n402 B.n312 10.6151
R1832 B.n402 B.n401 10.6151
R1833 B.n401 B.n400 10.6151
R1834 B.n400 B.n314 10.6151
R1835 B.n394 B.n314 10.6151
R1836 B.n394 B.n393 10.6151
R1837 B.n393 B.n392 10.6151
R1838 B.n392 B.n316 10.6151
R1839 B.n386 B.n385 10.6151
R1840 B.n385 B.n384 10.6151
R1841 B.n384 B.n321 10.6151
R1842 B.n378 B.n321 10.6151
R1843 B.n378 B.n377 10.6151
R1844 B.n377 B.n376 10.6151
R1845 B.n376 B.n323 10.6151
R1846 B.n370 B.n323 10.6151
R1847 B.n368 B.n367 10.6151
R1848 B.n367 B.n327 10.6151
R1849 B.n361 B.n327 10.6151
R1850 B.n361 B.n360 10.6151
R1851 B.n360 B.n359 10.6151
R1852 B.n359 B.n329 10.6151
R1853 B.n353 B.n329 10.6151
R1854 B.n353 B.n352 10.6151
R1855 B.n352 B.n351 10.6151
R1856 B.n351 B.n331 10.6151
R1857 B.n345 B.n331 10.6151
R1858 B.n345 B.n344 10.6151
R1859 B.n344 B.n343 10.6151
R1860 B.n343 B.n333 10.6151
R1861 B.n337 B.n333 10.6151
R1862 B.n337 B.n336 10.6151
R1863 B.n336 B.n304 10.6151
R1864 B.n428 B.n427 10.6151
R1865 B.n429 B.n428 10.6151
R1866 B.n429 B.n296 10.6151
R1867 B.n439 B.n296 10.6151
R1868 B.n440 B.n439 10.6151
R1869 B.n441 B.n440 10.6151
R1870 B.n441 B.n288 10.6151
R1871 B.n451 B.n288 10.6151
R1872 B.n452 B.n451 10.6151
R1873 B.n453 B.n452 10.6151
R1874 B.n453 B.n280 10.6151
R1875 B.n463 B.n280 10.6151
R1876 B.n464 B.n463 10.6151
R1877 B.n465 B.n464 10.6151
R1878 B.n465 B.n272 10.6151
R1879 B.n475 B.n272 10.6151
R1880 B.n476 B.n475 10.6151
R1881 B.n477 B.n476 10.6151
R1882 B.n477 B.n264 10.6151
R1883 B.n487 B.n264 10.6151
R1884 B.n488 B.n487 10.6151
R1885 B.n489 B.n488 10.6151
R1886 B.n489 B.n257 10.6151
R1887 B.n499 B.n257 10.6151
R1888 B.n500 B.n499 10.6151
R1889 B.n501 B.n500 10.6151
R1890 B.n501 B.n249 10.6151
R1891 B.n511 B.n249 10.6151
R1892 B.n512 B.n511 10.6151
R1893 B.n513 B.n512 10.6151
R1894 B.n513 B.n241 10.6151
R1895 B.n523 B.n241 10.6151
R1896 B.n524 B.n523 10.6151
R1897 B.n525 B.n524 10.6151
R1898 B.n525 B.n233 10.6151
R1899 B.n535 B.n233 10.6151
R1900 B.n536 B.n535 10.6151
R1901 B.n537 B.n536 10.6151
R1902 B.n537 B.n225 10.6151
R1903 B.n547 B.n225 10.6151
R1904 B.n548 B.n547 10.6151
R1905 B.n549 B.n548 10.6151
R1906 B.n549 B.n216 10.6151
R1907 B.n559 B.n216 10.6151
R1908 B.n560 B.n559 10.6151
R1909 B.n561 B.n560 10.6151
R1910 B.n561 B.n209 10.6151
R1911 B.n571 B.n209 10.6151
R1912 B.n572 B.n571 10.6151
R1913 B.n573 B.n572 10.6151
R1914 B.n573 B.n201 10.6151
R1915 B.n583 B.n201 10.6151
R1916 B.n584 B.n583 10.6151
R1917 B.n585 B.n584 10.6151
R1918 B.n585 B.n193 10.6151
R1919 B.n595 B.n193 10.6151
R1920 B.n596 B.n595 10.6151
R1921 B.n597 B.n596 10.6151
R1922 B.n597 B.n185 10.6151
R1923 B.n607 B.n185 10.6151
R1924 B.n608 B.n607 10.6151
R1925 B.n609 B.n608 10.6151
R1926 B.n609 B.n177 10.6151
R1927 B.n619 B.n177 10.6151
R1928 B.n620 B.n619 10.6151
R1929 B.n621 B.n620 10.6151
R1930 B.n621 B.n170 10.6151
R1931 B.n632 B.n170 10.6151
R1932 B.n633 B.n632 10.6151
R1933 B.n635 B.n633 10.6151
R1934 B.n635 B.n634 10.6151
R1935 B.n634 B.n162 10.6151
R1936 B.n646 B.n162 10.6151
R1937 B.n647 B.n646 10.6151
R1938 B.n648 B.n647 10.6151
R1939 B.n649 B.n648 10.6151
R1940 B.n650 B.n649 10.6151
R1941 B.n653 B.n650 10.6151
R1942 B.n654 B.n653 10.6151
R1943 B.n655 B.n654 10.6151
R1944 B.n656 B.n655 10.6151
R1945 B.n658 B.n656 10.6151
R1946 B.n659 B.n658 10.6151
R1947 B.n660 B.n659 10.6151
R1948 B.n661 B.n660 10.6151
R1949 B.n663 B.n661 10.6151
R1950 B.n664 B.n663 10.6151
R1951 B.n665 B.n664 10.6151
R1952 B.n666 B.n665 10.6151
R1953 B.n668 B.n666 10.6151
R1954 B.n669 B.n668 10.6151
R1955 B.n670 B.n669 10.6151
R1956 B.n671 B.n670 10.6151
R1957 B.n673 B.n671 10.6151
R1958 B.n674 B.n673 10.6151
R1959 B.n675 B.n674 10.6151
R1960 B.n676 B.n675 10.6151
R1961 B.n678 B.n676 10.6151
R1962 B.n679 B.n678 10.6151
R1963 B.n680 B.n679 10.6151
R1964 B.n681 B.n680 10.6151
R1965 B.n683 B.n681 10.6151
R1966 B.n684 B.n683 10.6151
R1967 B.n685 B.n684 10.6151
R1968 B.n686 B.n685 10.6151
R1969 B.n688 B.n686 10.6151
R1970 B.n689 B.n688 10.6151
R1971 B.n690 B.n689 10.6151
R1972 B.n691 B.n690 10.6151
R1973 B.n693 B.n691 10.6151
R1974 B.n694 B.n693 10.6151
R1975 B.n695 B.n694 10.6151
R1976 B.n696 B.n695 10.6151
R1977 B.n698 B.n696 10.6151
R1978 B.n699 B.n698 10.6151
R1979 B.n700 B.n699 10.6151
R1980 B.n701 B.n700 10.6151
R1981 B.n703 B.n701 10.6151
R1982 B.n704 B.n703 10.6151
R1983 B.n705 B.n704 10.6151
R1984 B.n706 B.n705 10.6151
R1985 B.n708 B.n706 10.6151
R1986 B.n709 B.n708 10.6151
R1987 B.n710 B.n709 10.6151
R1988 B.n711 B.n710 10.6151
R1989 B.n713 B.n711 10.6151
R1990 B.n714 B.n713 10.6151
R1991 B.n715 B.n714 10.6151
R1992 B.n716 B.n715 10.6151
R1993 B.n718 B.n716 10.6151
R1994 B.n719 B.n718 10.6151
R1995 B.n720 B.n719 10.6151
R1996 B.n721 B.n720 10.6151
R1997 B.n723 B.n721 10.6151
R1998 B.n724 B.n723 10.6151
R1999 B.n725 B.n724 10.6151
R2000 B.n726 B.n725 10.6151
R2001 B.n728 B.n726 10.6151
R2002 B.n729 B.n728 10.6151
R2003 B.n730 B.n729 10.6151
R2004 B.n731 B.n730 10.6151
R2005 B.n733 B.n731 10.6151
R2006 B.n734 B.n733 10.6151
R2007 B.n735 B.n734 10.6151
R2008 B.n736 B.n735 10.6151
R2009 B.n738 B.n736 10.6151
R2010 B.n739 B.n738 10.6151
R2011 B.n740 B.n739 10.6151
R2012 B.n741 B.n740 10.6151
R2013 B.n977 B.n1 10.6151
R2014 B.n977 B.n976 10.6151
R2015 B.n976 B.n975 10.6151
R2016 B.n975 B.n10 10.6151
R2017 B.n969 B.n10 10.6151
R2018 B.n969 B.n968 10.6151
R2019 B.n968 B.n967 10.6151
R2020 B.n967 B.n17 10.6151
R2021 B.n961 B.n17 10.6151
R2022 B.n961 B.n960 10.6151
R2023 B.n960 B.n959 10.6151
R2024 B.n959 B.n25 10.6151
R2025 B.n953 B.n25 10.6151
R2026 B.n953 B.n952 10.6151
R2027 B.n952 B.n951 10.6151
R2028 B.n951 B.n32 10.6151
R2029 B.n945 B.n32 10.6151
R2030 B.n945 B.n944 10.6151
R2031 B.n944 B.n943 10.6151
R2032 B.n943 B.n39 10.6151
R2033 B.n937 B.n39 10.6151
R2034 B.n937 B.n936 10.6151
R2035 B.n936 B.n935 10.6151
R2036 B.n935 B.n46 10.6151
R2037 B.n929 B.n46 10.6151
R2038 B.n929 B.n928 10.6151
R2039 B.n928 B.n927 10.6151
R2040 B.n927 B.n53 10.6151
R2041 B.n921 B.n53 10.6151
R2042 B.n921 B.n920 10.6151
R2043 B.n920 B.n919 10.6151
R2044 B.n919 B.n60 10.6151
R2045 B.n913 B.n60 10.6151
R2046 B.n913 B.n912 10.6151
R2047 B.n912 B.n911 10.6151
R2048 B.n911 B.n67 10.6151
R2049 B.n905 B.n67 10.6151
R2050 B.n905 B.n904 10.6151
R2051 B.n904 B.n903 10.6151
R2052 B.n903 B.n74 10.6151
R2053 B.n897 B.n74 10.6151
R2054 B.n897 B.n896 10.6151
R2055 B.n896 B.n895 10.6151
R2056 B.n895 B.n81 10.6151
R2057 B.n889 B.n81 10.6151
R2058 B.n889 B.n888 10.6151
R2059 B.n888 B.n887 10.6151
R2060 B.n887 B.n88 10.6151
R2061 B.n881 B.n88 10.6151
R2062 B.n881 B.n880 10.6151
R2063 B.n880 B.n879 10.6151
R2064 B.n879 B.n94 10.6151
R2065 B.n873 B.n94 10.6151
R2066 B.n873 B.n872 10.6151
R2067 B.n872 B.n871 10.6151
R2068 B.n871 B.n101 10.6151
R2069 B.n865 B.n101 10.6151
R2070 B.n865 B.n864 10.6151
R2071 B.n864 B.n863 10.6151
R2072 B.n863 B.n108 10.6151
R2073 B.n857 B.n108 10.6151
R2074 B.n857 B.n856 10.6151
R2075 B.n856 B.n855 10.6151
R2076 B.n855 B.n115 10.6151
R2077 B.n849 B.n115 10.6151
R2078 B.n849 B.n848 10.6151
R2079 B.n848 B.n847 10.6151
R2080 B.n847 B.n122 10.6151
R2081 B.n841 B.n122 10.6151
R2082 B.n841 B.n840 10.6151
R2083 B.n840 B.n839 10.6151
R2084 B.n839 B.n129 10.6151
R2085 B.n833 B.n129 10.6151
R2086 B.n832 B.n831 10.6151
R2087 B.n831 B.n136 10.6151
R2088 B.n825 B.n136 10.6151
R2089 B.n825 B.n824 10.6151
R2090 B.n824 B.n823 10.6151
R2091 B.n823 B.n138 10.6151
R2092 B.n817 B.n138 10.6151
R2093 B.n817 B.n816 10.6151
R2094 B.n816 B.n815 10.6151
R2095 B.n815 B.n140 10.6151
R2096 B.n809 B.n140 10.6151
R2097 B.n809 B.n808 10.6151
R2098 B.n808 B.n807 10.6151
R2099 B.n807 B.n142 10.6151
R2100 B.n801 B.n142 10.6151
R2101 B.n801 B.n800 10.6151
R2102 B.n800 B.n799 10.6151
R2103 B.n795 B.n794 10.6151
R2104 B.n794 B.n148 10.6151
R2105 B.n789 B.n148 10.6151
R2106 B.n789 B.n788 10.6151
R2107 B.n788 B.n787 10.6151
R2108 B.n787 B.n150 10.6151
R2109 B.n781 B.n150 10.6151
R2110 B.n781 B.n780 10.6151
R2111 B.n778 B.n154 10.6151
R2112 B.n772 B.n154 10.6151
R2113 B.n772 B.n771 10.6151
R2114 B.n771 B.n770 10.6151
R2115 B.n770 B.n156 10.6151
R2116 B.n764 B.n156 10.6151
R2117 B.n764 B.n763 10.6151
R2118 B.n763 B.n762 10.6151
R2119 B.n762 B.n158 10.6151
R2120 B.n756 B.n158 10.6151
R2121 B.n756 B.n755 10.6151
R2122 B.n755 B.n754 10.6151
R2123 B.n754 B.n160 10.6151
R2124 B.n748 B.n160 10.6151
R2125 B.n748 B.n747 10.6151
R2126 B.n747 B.n746 10.6151
R2127 B.n746 B.n742 10.6151
R2128 B.n985 B.n0 8.11757
R2129 B.n985 B.n1 8.11757
R2130 B.n527 B.t9 7.27323
R2131 B.n901 B.t8 7.27323
R2132 B.n386 B.n320 6.5566
R2133 B.n370 B.n369 6.5566
R2134 B.n795 B.n146 6.5566
R2135 B.n780 B.n779 6.5566
R2136 B.n320 B.n316 4.05904
R2137 B.n369 B.n368 4.05904
R2138 B.n799 B.n146 4.05904
R2139 B.n779 B.n778 4.05904
R2140 VP.n32 VP.n29 161.3
R2141 VP.n34 VP.n33 161.3
R2142 VP.n35 VP.n28 161.3
R2143 VP.n37 VP.n36 161.3
R2144 VP.n38 VP.n27 161.3
R2145 VP.n40 VP.n39 161.3
R2146 VP.n41 VP.n26 161.3
R2147 VP.n44 VP.n43 161.3
R2148 VP.n45 VP.n25 161.3
R2149 VP.n47 VP.n46 161.3
R2150 VP.n48 VP.n24 161.3
R2151 VP.n50 VP.n49 161.3
R2152 VP.n51 VP.n23 161.3
R2153 VP.n53 VP.n52 161.3
R2154 VP.n54 VP.n22 161.3
R2155 VP.n56 VP.n55 161.3
R2156 VP.n58 VP.n57 161.3
R2157 VP.n59 VP.n20 161.3
R2158 VP.n61 VP.n60 161.3
R2159 VP.n62 VP.n19 161.3
R2160 VP.n64 VP.n63 161.3
R2161 VP.n65 VP.n18 161.3
R2162 VP.n67 VP.n66 161.3
R2163 VP.n117 VP.n116 161.3
R2164 VP.n115 VP.n1 161.3
R2165 VP.n114 VP.n113 161.3
R2166 VP.n112 VP.n2 161.3
R2167 VP.n111 VP.n110 161.3
R2168 VP.n109 VP.n3 161.3
R2169 VP.n108 VP.n107 161.3
R2170 VP.n106 VP.n105 161.3
R2171 VP.n104 VP.n5 161.3
R2172 VP.n103 VP.n102 161.3
R2173 VP.n101 VP.n6 161.3
R2174 VP.n100 VP.n99 161.3
R2175 VP.n98 VP.n7 161.3
R2176 VP.n97 VP.n96 161.3
R2177 VP.n95 VP.n8 161.3
R2178 VP.n94 VP.n93 161.3
R2179 VP.n91 VP.n9 161.3
R2180 VP.n90 VP.n89 161.3
R2181 VP.n88 VP.n10 161.3
R2182 VP.n87 VP.n86 161.3
R2183 VP.n85 VP.n11 161.3
R2184 VP.n84 VP.n83 161.3
R2185 VP.n82 VP.n12 161.3
R2186 VP.n81 VP.n80 161.3
R2187 VP.n78 VP.n13 161.3
R2188 VP.n77 VP.n76 161.3
R2189 VP.n75 VP.n14 161.3
R2190 VP.n74 VP.n73 161.3
R2191 VP.n72 VP.n15 161.3
R2192 VP.n71 VP.n70 161.3
R2193 VP.n69 VP.n16 75.9823
R2194 VP.n118 VP.n0 75.9823
R2195 VP.n68 VP.n17 75.9823
R2196 VP.n31 VP.n30 73.9636
R2197 VP.n31 VP.t0 59.4412
R2198 VP.n86 VP.n10 53.6554
R2199 VP.n99 VP.n6 53.6554
R2200 VP.n49 VP.n23 53.6554
R2201 VP.n36 VP.n27 53.6554
R2202 VP.n69 VP.n68 51.6094
R2203 VP.n77 VP.n14 49.7803
R2204 VP.n110 VP.n2 49.7803
R2205 VP.n60 VP.n19 49.7803
R2206 VP.n73 VP.n14 31.3737
R2207 VP.n114 VP.n2 31.3737
R2208 VP.n64 VP.n19 31.3737
R2209 VP.n90 VP.n10 27.4986
R2210 VP.n99 VP.n98 27.4986
R2211 VP.n49 VP.n48 27.4986
R2212 VP.n40 VP.n27 27.4986
R2213 VP.n16 VP.t4 26.6226
R2214 VP.n79 VP.t7 26.6226
R2215 VP.n92 VP.t3 26.6226
R2216 VP.n4 VP.t6 26.6226
R2217 VP.n0 VP.t9 26.6226
R2218 VP.n17 VP.t1 26.6226
R2219 VP.n21 VP.t8 26.6226
R2220 VP.n42 VP.t5 26.6226
R2221 VP.n30 VP.t2 26.6226
R2222 VP.n72 VP.n71 24.5923
R2223 VP.n73 VP.n72 24.5923
R2224 VP.n78 VP.n77 24.5923
R2225 VP.n80 VP.n78 24.5923
R2226 VP.n84 VP.n12 24.5923
R2227 VP.n85 VP.n84 24.5923
R2228 VP.n86 VP.n85 24.5923
R2229 VP.n91 VP.n90 24.5923
R2230 VP.n93 VP.n91 24.5923
R2231 VP.n97 VP.n8 24.5923
R2232 VP.n98 VP.n97 24.5923
R2233 VP.n103 VP.n6 24.5923
R2234 VP.n104 VP.n103 24.5923
R2235 VP.n105 VP.n104 24.5923
R2236 VP.n109 VP.n108 24.5923
R2237 VP.n110 VP.n109 24.5923
R2238 VP.n115 VP.n114 24.5923
R2239 VP.n116 VP.n115 24.5923
R2240 VP.n65 VP.n64 24.5923
R2241 VP.n66 VP.n65 24.5923
R2242 VP.n53 VP.n23 24.5923
R2243 VP.n54 VP.n53 24.5923
R2244 VP.n55 VP.n54 24.5923
R2245 VP.n59 VP.n58 24.5923
R2246 VP.n60 VP.n59 24.5923
R2247 VP.n41 VP.n40 24.5923
R2248 VP.n43 VP.n41 24.5923
R2249 VP.n47 VP.n25 24.5923
R2250 VP.n48 VP.n47 24.5923
R2251 VP.n34 VP.n29 24.5923
R2252 VP.n35 VP.n34 24.5923
R2253 VP.n36 VP.n35 24.5923
R2254 VP.n80 VP.n79 23.6087
R2255 VP.n108 VP.n4 23.6087
R2256 VP.n58 VP.n21 23.6087
R2257 VP.n71 VP.n16 14.2638
R2258 VP.n116 VP.n0 14.2638
R2259 VP.n66 VP.n17 14.2638
R2260 VP.n93 VP.n92 12.2964
R2261 VP.n92 VP.n8 12.2964
R2262 VP.n43 VP.n42 12.2964
R2263 VP.n42 VP.n25 12.2964
R2264 VP.n32 VP.n31 4.18334
R2265 VP.n79 VP.n12 0.984173
R2266 VP.n105 VP.n4 0.984173
R2267 VP.n55 VP.n21 0.984173
R2268 VP.n30 VP.n29 0.984173
R2269 VP.n68 VP.n67 0.354861
R2270 VP.n70 VP.n69 0.354861
R2271 VP.n118 VP.n117 0.354861
R2272 VP VP.n118 0.267071
R2273 VP.n33 VP.n32 0.189894
R2274 VP.n33 VP.n28 0.189894
R2275 VP.n37 VP.n28 0.189894
R2276 VP.n38 VP.n37 0.189894
R2277 VP.n39 VP.n38 0.189894
R2278 VP.n39 VP.n26 0.189894
R2279 VP.n44 VP.n26 0.189894
R2280 VP.n45 VP.n44 0.189894
R2281 VP.n46 VP.n45 0.189894
R2282 VP.n46 VP.n24 0.189894
R2283 VP.n50 VP.n24 0.189894
R2284 VP.n51 VP.n50 0.189894
R2285 VP.n52 VP.n51 0.189894
R2286 VP.n52 VP.n22 0.189894
R2287 VP.n56 VP.n22 0.189894
R2288 VP.n57 VP.n56 0.189894
R2289 VP.n57 VP.n20 0.189894
R2290 VP.n61 VP.n20 0.189894
R2291 VP.n62 VP.n61 0.189894
R2292 VP.n63 VP.n62 0.189894
R2293 VP.n63 VP.n18 0.189894
R2294 VP.n67 VP.n18 0.189894
R2295 VP.n70 VP.n15 0.189894
R2296 VP.n74 VP.n15 0.189894
R2297 VP.n75 VP.n74 0.189894
R2298 VP.n76 VP.n75 0.189894
R2299 VP.n76 VP.n13 0.189894
R2300 VP.n81 VP.n13 0.189894
R2301 VP.n82 VP.n81 0.189894
R2302 VP.n83 VP.n82 0.189894
R2303 VP.n83 VP.n11 0.189894
R2304 VP.n87 VP.n11 0.189894
R2305 VP.n88 VP.n87 0.189894
R2306 VP.n89 VP.n88 0.189894
R2307 VP.n89 VP.n9 0.189894
R2308 VP.n94 VP.n9 0.189894
R2309 VP.n95 VP.n94 0.189894
R2310 VP.n96 VP.n95 0.189894
R2311 VP.n96 VP.n7 0.189894
R2312 VP.n100 VP.n7 0.189894
R2313 VP.n101 VP.n100 0.189894
R2314 VP.n102 VP.n101 0.189894
R2315 VP.n102 VP.n5 0.189894
R2316 VP.n106 VP.n5 0.189894
R2317 VP.n107 VP.n106 0.189894
R2318 VP.n107 VP.n3 0.189894
R2319 VP.n111 VP.n3 0.189894
R2320 VP.n112 VP.n111 0.189894
R2321 VP.n113 VP.n112 0.189894
R2322 VP.n113 VP.n1 0.189894
R2323 VP.n117 VP.n1 0.189894
R2324 VDD1.n14 VDD1.n0 289.615
R2325 VDD1.n35 VDD1.n21 289.615
R2326 VDD1.n15 VDD1.n14 185
R2327 VDD1.n13 VDD1.n12 185
R2328 VDD1.n4 VDD1.n3 185
R2329 VDD1.n7 VDD1.n6 185
R2330 VDD1.n28 VDD1.n27 185
R2331 VDD1.n25 VDD1.n24 185
R2332 VDD1.n34 VDD1.n33 185
R2333 VDD1.n36 VDD1.n35 185
R2334 VDD1.t9 VDD1.n5 147.888
R2335 VDD1.t5 VDD1.n26 147.888
R2336 VDD1.n14 VDD1.n13 104.615
R2337 VDD1.n13 VDD1.n3 104.615
R2338 VDD1.n6 VDD1.n3 104.615
R2339 VDD1.n27 VDD1.n24 104.615
R2340 VDD1.n34 VDD1.n24 104.615
R2341 VDD1.n35 VDD1.n34 104.615
R2342 VDD1.n43 VDD1.n42 75.0704
R2343 VDD1.n20 VDD1.n19 72.6883
R2344 VDD1.n45 VDD1.n44 72.6882
R2345 VDD1.n41 VDD1.n40 72.6882
R2346 VDD1.n6 VDD1.t9 52.3082
R2347 VDD1.n27 VDD1.t5 52.3082
R2348 VDD1.n20 VDD1.n18 51.3384
R2349 VDD1.n41 VDD1.n39 51.3384
R2350 VDD1.n45 VDD1.n43 44.6367
R2351 VDD1.n7 VDD1.n5 15.6496
R2352 VDD1.n28 VDD1.n26 15.6496
R2353 VDD1.n8 VDD1.n4 12.8005
R2354 VDD1.n29 VDD1.n25 12.8005
R2355 VDD1.n12 VDD1.n11 12.0247
R2356 VDD1.n33 VDD1.n32 12.0247
R2357 VDD1.n15 VDD1.n2 11.249
R2358 VDD1.n36 VDD1.n23 11.249
R2359 VDD1.n16 VDD1.n0 10.4732
R2360 VDD1.n37 VDD1.n21 10.4732
R2361 VDD1.n18 VDD1.n17 9.45567
R2362 VDD1.n39 VDD1.n38 9.45567
R2363 VDD1.n17 VDD1.n16 9.3005
R2364 VDD1.n2 VDD1.n1 9.3005
R2365 VDD1.n11 VDD1.n10 9.3005
R2366 VDD1.n9 VDD1.n8 9.3005
R2367 VDD1.n38 VDD1.n37 9.3005
R2368 VDD1.n23 VDD1.n22 9.3005
R2369 VDD1.n32 VDD1.n31 9.3005
R2370 VDD1.n30 VDD1.n29 9.3005
R2371 VDD1.n44 VDD1.t1 5.21103
R2372 VDD1.n44 VDD1.t8 5.21103
R2373 VDD1.n19 VDD1.t7 5.21103
R2374 VDD1.n19 VDD1.t4 5.21103
R2375 VDD1.n42 VDD1.t3 5.21103
R2376 VDD1.n42 VDD1.t0 5.21103
R2377 VDD1.n40 VDD1.t2 5.21103
R2378 VDD1.n40 VDD1.t6 5.21103
R2379 VDD1.n9 VDD1.n5 4.40546
R2380 VDD1.n30 VDD1.n26 4.40546
R2381 VDD1.n18 VDD1.n0 3.49141
R2382 VDD1.n39 VDD1.n21 3.49141
R2383 VDD1.n16 VDD1.n15 2.71565
R2384 VDD1.n37 VDD1.n36 2.71565
R2385 VDD1 VDD1.n45 2.37981
R2386 VDD1.n12 VDD1.n2 1.93989
R2387 VDD1.n33 VDD1.n23 1.93989
R2388 VDD1.n11 VDD1.n4 1.16414
R2389 VDD1.n32 VDD1.n25 1.16414
R2390 VDD1 VDD1.n20 0.87119
R2391 VDD1.n43 VDD1.n41 0.757654
R2392 VDD1.n8 VDD1.n7 0.388379
R2393 VDD1.n29 VDD1.n28 0.388379
R2394 VDD1.n17 VDD1.n1 0.155672
R2395 VDD1.n10 VDD1.n1 0.155672
R2396 VDD1.n10 VDD1.n9 0.155672
R2397 VDD1.n31 VDD1.n30 0.155672
R2398 VDD1.n31 VDD1.n22 0.155672
R2399 VDD1.n38 VDD1.n22 0.155672
C0 VP VDD2 0.695822f
C1 VN VDD2 3.92291f
C2 VTAIL VDD2 7.506431f
C3 VDD1 VP 4.45481f
C4 VN VDD1 0.160043f
C5 VDD1 VTAIL 7.4477f
C6 VDD1 VDD2 2.72073f
C7 VN VP 8.11497f
C8 VTAIL VP 5.63609f
C9 VN VTAIL 5.62195f
C10 VDD2 B 6.84079f
C11 VDD1 B 6.735372f
C12 VTAIL B 4.943583f
C13 VN B 21.3671f
C14 VP B 19.83666f
C15 VDD1.n0 B 0.037516f
C16 VDD1.n1 B 0.028911f
C17 VDD1.n2 B 0.015535f
C18 VDD1.n3 B 0.03672f
C19 VDD1.n4 B 0.016449f
C20 VDD1.n5 B 0.109176f
C21 VDD1.t9 B 0.060506f
C22 VDD1.n6 B 0.02754f
C23 VDD1.n7 B 0.021612f
C24 VDD1.n8 B 0.015535f
C25 VDD1.n9 B 0.394209f
C26 VDD1.n10 B 0.028911f
C27 VDD1.n11 B 0.015535f
C28 VDD1.n12 B 0.016449f
C29 VDD1.n13 B 0.03672f
C30 VDD1.n14 B 0.073974f
C31 VDD1.n15 B 0.016449f
C32 VDD1.n16 B 0.015535f
C33 VDD1.n17 B 0.065247f
C34 VDD1.n18 B 0.083384f
C35 VDD1.t7 B 0.086816f
C36 VDD1.t4 B 0.086816f
C37 VDD1.n19 B 0.677035f
C38 VDD1.n20 B 0.941365f
C39 VDD1.n21 B 0.037516f
C40 VDD1.n22 B 0.028911f
C41 VDD1.n23 B 0.015535f
C42 VDD1.n24 B 0.03672f
C43 VDD1.n25 B 0.016449f
C44 VDD1.n26 B 0.109176f
C45 VDD1.t5 B 0.060506f
C46 VDD1.n27 B 0.02754f
C47 VDD1.n28 B 0.021612f
C48 VDD1.n29 B 0.015535f
C49 VDD1.n30 B 0.394209f
C50 VDD1.n31 B 0.028911f
C51 VDD1.n32 B 0.015535f
C52 VDD1.n33 B 0.016449f
C53 VDD1.n34 B 0.03672f
C54 VDD1.n35 B 0.073974f
C55 VDD1.n36 B 0.016449f
C56 VDD1.n37 B 0.015535f
C57 VDD1.n38 B 0.065247f
C58 VDD1.n39 B 0.083384f
C59 VDD1.t2 B 0.086816f
C60 VDD1.t6 B 0.086816f
C61 VDD1.n40 B 0.677032f
C62 VDD1.n41 B 0.931677f
C63 VDD1.t3 B 0.086816f
C64 VDD1.t0 B 0.086816f
C65 VDD1.n42 B 0.701124f
C66 VDD1.n43 B 3.43768f
C67 VDD1.t1 B 0.086816f
C68 VDD1.t8 B 0.086816f
C69 VDD1.n44 B 0.677032f
C70 VDD1.n45 B 3.32793f
C71 VP.t9 B 0.788747f
C72 VP.n0 B 0.404871f
C73 VP.n1 B 0.023601f
C74 VP.n2 B 0.021924f
C75 VP.n3 B 0.023601f
C76 VP.t6 B 0.788747f
C77 VP.n4 B 0.309802f
C78 VP.n5 B 0.023601f
C79 VP.n6 B 0.041425f
C80 VP.n7 B 0.023601f
C81 VP.n8 B 0.032963f
C82 VP.n9 B 0.023601f
C83 VP.n10 B 0.02518f
C84 VP.n11 B 0.023601f
C85 VP.n12 B 0.023024f
C86 VP.n13 B 0.023601f
C87 VP.n14 B 0.021924f
C88 VP.n15 B 0.023601f
C89 VP.t4 B 0.788747f
C90 VP.n16 B 0.404871f
C91 VP.t1 B 0.788747f
C92 VP.n17 B 0.404871f
C93 VP.n18 B 0.023601f
C94 VP.n19 B 0.021924f
C95 VP.n20 B 0.023601f
C96 VP.t8 B 0.788747f
C97 VP.n21 B 0.309802f
C98 VP.n22 B 0.023601f
C99 VP.n23 B 0.041425f
C100 VP.n24 B 0.023601f
C101 VP.n25 B 0.032963f
C102 VP.n26 B 0.023601f
C103 VP.n27 B 0.02518f
C104 VP.n28 B 0.023601f
C105 VP.n29 B 0.023024f
C106 VP.t0 B 1.05429f
C107 VP.t2 B 0.788747f
C108 VP.n30 B 0.381304f
C109 VP.n31 B 0.377042f
C110 VP.n32 B 0.28163f
C111 VP.n33 B 0.023601f
C112 VP.n34 B 0.043765f
C113 VP.n35 B 0.043765f
C114 VP.n36 B 0.041425f
C115 VP.n37 B 0.023601f
C116 VP.n38 B 0.023601f
C117 VP.n39 B 0.023601f
C118 VP.n40 B 0.045775f
C119 VP.n41 B 0.043765f
C120 VP.t5 B 0.788747f
C121 VP.n42 B 0.309802f
C122 VP.n43 B 0.032963f
C123 VP.n44 B 0.023601f
C124 VP.n45 B 0.023601f
C125 VP.n46 B 0.023601f
C126 VP.n47 B 0.043765f
C127 VP.n48 B 0.045775f
C128 VP.n49 B 0.02518f
C129 VP.n50 B 0.023601f
C130 VP.n51 B 0.023601f
C131 VP.n52 B 0.023601f
C132 VP.n53 B 0.043765f
C133 VP.n54 B 0.043765f
C134 VP.n55 B 0.023024f
C135 VP.n56 B 0.023601f
C136 VP.n57 B 0.023601f
C137 VP.n58 B 0.042901f
C138 VP.n59 B 0.043765f
C139 VP.n60 B 0.043328f
C140 VP.n61 B 0.023601f
C141 VP.n62 B 0.023601f
C142 VP.n63 B 0.023601f
C143 VP.n64 B 0.047128f
C144 VP.n65 B 0.043765f
C145 VP.n66 B 0.034691f
C146 VP.n67 B 0.038085f
C147 VP.n68 B 1.4075f
C148 VP.n69 B 1.42398f
C149 VP.n70 B 0.038085f
C150 VP.n71 B 0.034691f
C151 VP.n72 B 0.043765f
C152 VP.n73 B 0.047128f
C153 VP.n74 B 0.023601f
C154 VP.n75 B 0.023601f
C155 VP.n76 B 0.023601f
C156 VP.n77 B 0.043328f
C157 VP.n78 B 0.043765f
C158 VP.t7 B 0.788747f
C159 VP.n79 B 0.309802f
C160 VP.n80 B 0.042901f
C161 VP.n81 B 0.023601f
C162 VP.n82 B 0.023601f
C163 VP.n83 B 0.023601f
C164 VP.n84 B 0.043765f
C165 VP.n85 B 0.043765f
C166 VP.n86 B 0.041425f
C167 VP.n87 B 0.023601f
C168 VP.n88 B 0.023601f
C169 VP.n89 B 0.023601f
C170 VP.n90 B 0.045775f
C171 VP.n91 B 0.043765f
C172 VP.t3 B 0.788747f
C173 VP.n92 B 0.309802f
C174 VP.n93 B 0.032963f
C175 VP.n94 B 0.023601f
C176 VP.n95 B 0.023601f
C177 VP.n96 B 0.023601f
C178 VP.n97 B 0.043765f
C179 VP.n98 B 0.045775f
C180 VP.n99 B 0.02518f
C181 VP.n100 B 0.023601f
C182 VP.n101 B 0.023601f
C183 VP.n102 B 0.023601f
C184 VP.n103 B 0.043765f
C185 VP.n104 B 0.043765f
C186 VP.n105 B 0.023024f
C187 VP.n106 B 0.023601f
C188 VP.n107 B 0.023601f
C189 VP.n108 B 0.042901f
C190 VP.n109 B 0.043765f
C191 VP.n110 B 0.043328f
C192 VP.n111 B 0.023601f
C193 VP.n112 B 0.023601f
C194 VP.n113 B 0.023601f
C195 VP.n114 B 0.047128f
C196 VP.n115 B 0.043765f
C197 VP.n116 B 0.034691f
C198 VP.n117 B 0.038085f
C199 VP.n118 B 0.058891f
C200 VDD2.n0 B 0.036498f
C201 VDD2.n1 B 0.028127f
C202 VDD2.n2 B 0.015114f
C203 VDD2.n3 B 0.035724f
C204 VDD2.n4 B 0.016003f
C205 VDD2.n5 B 0.106214f
C206 VDD2.t2 B 0.058864f
C207 VDD2.n6 B 0.026793f
C208 VDD2.n7 B 0.021026f
C209 VDD2.n8 B 0.015114f
C210 VDD2.n9 B 0.383513f
C211 VDD2.n10 B 0.028127f
C212 VDD2.n11 B 0.015114f
C213 VDD2.n12 B 0.016003f
C214 VDD2.n13 B 0.035724f
C215 VDD2.n14 B 0.071967f
C216 VDD2.n15 B 0.016003f
C217 VDD2.n16 B 0.015114f
C218 VDD2.n17 B 0.063476f
C219 VDD2.n18 B 0.081122f
C220 VDD2.t7 B 0.084461f
C221 VDD2.t5 B 0.084461f
C222 VDD2.n19 B 0.658663f
C223 VDD2.n20 B 0.906399f
C224 VDD2.t8 B 0.084461f
C225 VDD2.t6 B 0.084461f
C226 VDD2.n21 B 0.682101f
C227 VDD2.n22 B 3.18666f
C228 VDD2.n23 B 0.036498f
C229 VDD2.n24 B 0.028127f
C230 VDD2.n25 B 0.015114f
C231 VDD2.n26 B 0.035724f
C232 VDD2.n27 B 0.016003f
C233 VDD2.n28 B 0.106214f
C234 VDD2.t9 B 0.058864f
C235 VDD2.n29 B 0.026793f
C236 VDD2.n30 B 0.021026f
C237 VDD2.n31 B 0.015114f
C238 VDD2.n32 B 0.383513f
C239 VDD2.n33 B 0.028127f
C240 VDD2.n34 B 0.015114f
C241 VDD2.n35 B 0.016003f
C242 VDD2.n36 B 0.035724f
C243 VDD2.n37 B 0.071967f
C244 VDD2.n38 B 0.016003f
C245 VDD2.n39 B 0.015114f
C246 VDD2.n40 B 0.063476f
C247 VDD2.n41 B 0.059102f
C248 VDD2.n42 B 2.90126f
C249 VDD2.t1 B 0.084461f
C250 VDD2.t4 B 0.084461f
C251 VDD2.n43 B 0.658667f
C252 VDD2.n44 B 0.590016f
C253 VDD2.t0 B 0.084461f
C254 VDD2.t3 B 0.084461f
C255 VDD2.n45 B 0.682057f
C256 VTAIL.t19 B 0.098977f
C257 VTAIL.t16 B 0.098977f
C258 VTAIL.n0 B 0.698167f
C259 VTAIL.n1 B 0.770233f
C260 VTAIL.n2 B 0.042771f
C261 VTAIL.n3 B 0.032961f
C262 VTAIL.n4 B 0.017712f
C263 VTAIL.n5 B 0.041864f
C264 VTAIL.n6 B 0.018754f
C265 VTAIL.n7 B 0.12447f
C266 VTAIL.t1 B 0.068981f
C267 VTAIL.n8 B 0.031398f
C268 VTAIL.n9 B 0.02464f
C269 VTAIL.n10 B 0.017712f
C270 VTAIL.n11 B 0.44943f
C271 VTAIL.n12 B 0.032961f
C272 VTAIL.n13 B 0.017712f
C273 VTAIL.n14 B 0.018754f
C274 VTAIL.n15 B 0.041864f
C275 VTAIL.n16 B 0.084336f
C276 VTAIL.n17 B 0.018754f
C277 VTAIL.n18 B 0.017712f
C278 VTAIL.n19 B 0.074386f
C279 VTAIL.n20 B 0.046487f
C280 VTAIL.n21 B 0.594794f
C281 VTAIL.t6 B 0.098977f
C282 VTAIL.t2 B 0.098977f
C283 VTAIL.n22 B 0.698167f
C284 VTAIL.n23 B 0.973033f
C285 VTAIL.t4 B 0.098977f
C286 VTAIL.t9 B 0.098977f
C287 VTAIL.n24 B 0.698167f
C288 VTAIL.n25 B 2.11386f
C289 VTAIL.t17 B 0.098977f
C290 VTAIL.t13 B 0.098977f
C291 VTAIL.n26 B 0.698172f
C292 VTAIL.n27 B 2.11386f
C293 VTAIL.t15 B 0.098977f
C294 VTAIL.t12 B 0.098977f
C295 VTAIL.n28 B 0.698172f
C296 VTAIL.n29 B 0.973028f
C297 VTAIL.n30 B 0.042771f
C298 VTAIL.n31 B 0.032961f
C299 VTAIL.n32 B 0.017712f
C300 VTAIL.n33 B 0.041864f
C301 VTAIL.n34 B 0.018754f
C302 VTAIL.n35 B 0.12447f
C303 VTAIL.t18 B 0.068981f
C304 VTAIL.n36 B 0.031398f
C305 VTAIL.n37 B 0.02464f
C306 VTAIL.n38 B 0.017712f
C307 VTAIL.n39 B 0.44943f
C308 VTAIL.n40 B 0.032961f
C309 VTAIL.n41 B 0.017712f
C310 VTAIL.n42 B 0.018754f
C311 VTAIL.n43 B 0.041864f
C312 VTAIL.n44 B 0.084336f
C313 VTAIL.n45 B 0.018754f
C314 VTAIL.n46 B 0.017712f
C315 VTAIL.n47 B 0.074386f
C316 VTAIL.n48 B 0.046487f
C317 VTAIL.n49 B 0.594794f
C318 VTAIL.t5 B 0.098977f
C319 VTAIL.t0 B 0.098977f
C320 VTAIL.n50 B 0.698172f
C321 VTAIL.n51 B 0.850341f
C322 VTAIL.t3 B 0.098977f
C323 VTAIL.t8 B 0.098977f
C324 VTAIL.n52 B 0.698172f
C325 VTAIL.n53 B 0.973028f
C326 VTAIL.n54 B 0.042771f
C327 VTAIL.n55 B 0.032961f
C328 VTAIL.n56 B 0.017712f
C329 VTAIL.n57 B 0.041864f
C330 VTAIL.n58 B 0.018754f
C331 VTAIL.n59 B 0.12447f
C332 VTAIL.t7 B 0.068981f
C333 VTAIL.n60 B 0.031398f
C334 VTAIL.n61 B 0.02464f
C335 VTAIL.n62 B 0.017712f
C336 VTAIL.n63 B 0.44943f
C337 VTAIL.n64 B 0.032961f
C338 VTAIL.n65 B 0.017712f
C339 VTAIL.n66 B 0.018754f
C340 VTAIL.n67 B 0.041864f
C341 VTAIL.n68 B 0.084336f
C342 VTAIL.n69 B 0.018754f
C343 VTAIL.n70 B 0.017712f
C344 VTAIL.n71 B 0.074386f
C345 VTAIL.n72 B 0.046487f
C346 VTAIL.n73 B 1.51314f
C347 VTAIL.n74 B 0.042771f
C348 VTAIL.n75 B 0.032961f
C349 VTAIL.n76 B 0.017712f
C350 VTAIL.n77 B 0.041864f
C351 VTAIL.n78 B 0.018754f
C352 VTAIL.n79 B 0.12447f
C353 VTAIL.t14 B 0.068981f
C354 VTAIL.n80 B 0.031398f
C355 VTAIL.n81 B 0.02464f
C356 VTAIL.n82 B 0.017712f
C357 VTAIL.n83 B 0.44943f
C358 VTAIL.n84 B 0.032961f
C359 VTAIL.n85 B 0.017712f
C360 VTAIL.n86 B 0.018754f
C361 VTAIL.n87 B 0.041864f
C362 VTAIL.n88 B 0.084336f
C363 VTAIL.n89 B 0.018754f
C364 VTAIL.n90 B 0.017712f
C365 VTAIL.n91 B 0.074386f
C366 VTAIL.n92 B 0.046487f
C367 VTAIL.n93 B 1.51314f
C368 VTAIL.t11 B 0.098977f
C369 VTAIL.t10 B 0.098977f
C370 VTAIL.n94 B 0.698167f
C371 VTAIL.n95 B 0.707973f
C372 VN.t3 B 0.761357f
C373 VN.n0 B 0.390811f
C374 VN.n1 B 0.022781f
C375 VN.n2 B 0.021163f
C376 VN.n3 B 0.022781f
C377 VN.t1 B 0.761357f
C378 VN.n4 B 0.299044f
C379 VN.n5 B 0.022781f
C380 VN.n6 B 0.039986f
C381 VN.n7 B 0.022781f
C382 VN.n8 B 0.031818f
C383 VN.n9 B 0.022781f
C384 VN.n10 B 0.024306f
C385 VN.n11 B 0.022781f
C386 VN.n12 B 0.022224f
C387 VN.t2 B 0.761357f
C388 VN.n13 B 0.368063f
C389 VN.t7 B 1.01768f
C390 VN.n14 B 0.363949f
C391 VN.n15 B 0.271849f
C392 VN.n16 B 0.022781f
C393 VN.n17 B 0.042246f
C394 VN.n18 B 0.042246f
C395 VN.n19 B 0.039986f
C396 VN.n20 B 0.022781f
C397 VN.n21 B 0.022781f
C398 VN.n22 B 0.022781f
C399 VN.n23 B 0.044185f
C400 VN.n24 B 0.042246f
C401 VN.t4 B 0.761357f
C402 VN.n25 B 0.299044f
C403 VN.n26 B 0.031818f
C404 VN.n27 B 0.022781f
C405 VN.n28 B 0.022781f
C406 VN.n29 B 0.022781f
C407 VN.n30 B 0.042246f
C408 VN.n31 B 0.044185f
C409 VN.n32 B 0.024306f
C410 VN.n33 B 0.022781f
C411 VN.n34 B 0.022781f
C412 VN.n35 B 0.022781f
C413 VN.n36 B 0.042246f
C414 VN.n37 B 0.042246f
C415 VN.n38 B 0.022224f
C416 VN.n39 B 0.022781f
C417 VN.n40 B 0.022781f
C418 VN.n41 B 0.041411f
C419 VN.n42 B 0.042246f
C420 VN.n43 B 0.041824f
C421 VN.n44 B 0.022781f
C422 VN.n45 B 0.022781f
C423 VN.n46 B 0.022781f
C424 VN.n47 B 0.045491f
C425 VN.n48 B 0.042246f
C426 VN.n49 B 0.033486f
C427 VN.n50 B 0.036763f
C428 VN.n51 B 0.056846f
C429 VN.t0 B 0.761357f
C430 VN.n52 B 0.390811f
C431 VN.n53 B 0.022781f
C432 VN.n54 B 0.021163f
C433 VN.n55 B 0.022781f
C434 VN.t8 B 0.761357f
C435 VN.n56 B 0.299044f
C436 VN.n57 B 0.022781f
C437 VN.n58 B 0.039986f
C438 VN.n59 B 0.022781f
C439 VN.n60 B 0.031818f
C440 VN.n61 B 0.022781f
C441 VN.t5 B 0.761357f
C442 VN.n62 B 0.299044f
C443 VN.n63 B 0.024306f
C444 VN.n64 B 0.022781f
C445 VN.n65 B 0.022224f
C446 VN.t6 B 1.01768f
C447 VN.t9 B 0.761357f
C448 VN.n66 B 0.368063f
C449 VN.n67 B 0.363949f
C450 VN.n68 B 0.271849f
C451 VN.n69 B 0.022781f
C452 VN.n70 B 0.042246f
C453 VN.n71 B 0.042246f
C454 VN.n72 B 0.039986f
C455 VN.n73 B 0.022781f
C456 VN.n74 B 0.022781f
C457 VN.n75 B 0.022781f
C458 VN.n76 B 0.044185f
C459 VN.n77 B 0.042246f
C460 VN.n78 B 0.031818f
C461 VN.n79 B 0.022781f
C462 VN.n80 B 0.022781f
C463 VN.n81 B 0.022781f
C464 VN.n82 B 0.042246f
C465 VN.n83 B 0.044185f
C466 VN.n84 B 0.024306f
C467 VN.n85 B 0.022781f
C468 VN.n86 B 0.022781f
C469 VN.n87 B 0.022781f
C470 VN.n88 B 0.042246f
C471 VN.n89 B 0.042246f
C472 VN.n90 B 0.022224f
C473 VN.n91 B 0.022781f
C474 VN.n92 B 0.022781f
C475 VN.n93 B 0.041411f
C476 VN.n94 B 0.042246f
C477 VN.n95 B 0.041824f
C478 VN.n96 B 0.022781f
C479 VN.n97 B 0.022781f
C480 VN.n98 B 0.022781f
C481 VN.n99 B 0.045491f
C482 VN.n100 B 0.042246f
C483 VN.n101 B 0.033486f
C484 VN.n102 B 0.036763f
C485 VN.n103 B 1.36783f
.ends

