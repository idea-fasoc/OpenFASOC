* NGSPICE file created from diff_pair_sample_1368.ext - technology: sky130A

.subckt diff_pair_sample_1368 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n2752_n1790# sky130_fd_pr__pfet_01v8 ad=1.6029 pd=9 as=0 ps=0 w=4.11 l=2.64
X1 B.t8 B.t6 B.t7 w_n2752_n1790# sky130_fd_pr__pfet_01v8 ad=1.6029 pd=9 as=0 ps=0 w=4.11 l=2.64
X2 VTAIL.t7 VN.t0 VDD2.t3 w_n2752_n1790# sky130_fd_pr__pfet_01v8 ad=1.6029 pd=9 as=0.67815 ps=4.44 w=4.11 l=2.64
X3 B.t5 B.t3 B.t4 w_n2752_n1790# sky130_fd_pr__pfet_01v8 ad=1.6029 pd=9 as=0 ps=0 w=4.11 l=2.64
X4 VDD1.t3 VP.t0 VTAIL.t2 w_n2752_n1790# sky130_fd_pr__pfet_01v8 ad=0.67815 pd=4.44 as=1.6029 ps=9 w=4.11 l=2.64
X5 VDD2.t1 VN.t1 VTAIL.t6 w_n2752_n1790# sky130_fd_pr__pfet_01v8 ad=0.67815 pd=4.44 as=1.6029 ps=9 w=4.11 l=2.64
X6 VDD2.t0 VN.t2 VTAIL.t5 w_n2752_n1790# sky130_fd_pr__pfet_01v8 ad=0.67815 pd=4.44 as=1.6029 ps=9 w=4.11 l=2.64
X7 VTAIL.t4 VN.t3 VDD2.t2 w_n2752_n1790# sky130_fd_pr__pfet_01v8 ad=1.6029 pd=9 as=0.67815 ps=4.44 w=4.11 l=2.64
X8 VTAIL.t0 VP.t1 VDD1.t2 w_n2752_n1790# sky130_fd_pr__pfet_01v8 ad=1.6029 pd=9 as=0.67815 ps=4.44 w=4.11 l=2.64
X9 VDD1.t1 VP.t2 VTAIL.t1 w_n2752_n1790# sky130_fd_pr__pfet_01v8 ad=0.67815 pd=4.44 as=1.6029 ps=9 w=4.11 l=2.64
X10 B.t2 B.t0 B.t1 w_n2752_n1790# sky130_fd_pr__pfet_01v8 ad=1.6029 pd=9 as=0 ps=0 w=4.11 l=2.64
X11 VTAIL.t3 VP.t3 VDD1.t0 w_n2752_n1790# sky130_fd_pr__pfet_01v8 ad=1.6029 pd=9 as=0.67815 ps=4.44 w=4.11 l=2.64
R0 B.n245 B.n244 585
R1 B.n243 B.n82 585
R2 B.n242 B.n241 585
R3 B.n240 B.n83 585
R4 B.n239 B.n238 585
R5 B.n237 B.n84 585
R6 B.n236 B.n235 585
R7 B.n234 B.n85 585
R8 B.n233 B.n232 585
R9 B.n231 B.n86 585
R10 B.n230 B.n229 585
R11 B.n228 B.n87 585
R12 B.n227 B.n226 585
R13 B.n225 B.n88 585
R14 B.n224 B.n223 585
R15 B.n222 B.n89 585
R16 B.n221 B.n220 585
R17 B.n219 B.n90 585
R18 B.n218 B.n217 585
R19 B.n213 B.n91 585
R20 B.n212 B.n211 585
R21 B.n210 B.n92 585
R22 B.n209 B.n208 585
R23 B.n207 B.n93 585
R24 B.n206 B.n205 585
R25 B.n204 B.n94 585
R26 B.n203 B.n202 585
R27 B.n201 B.n95 585
R28 B.n199 B.n198 585
R29 B.n197 B.n98 585
R30 B.n196 B.n195 585
R31 B.n194 B.n99 585
R32 B.n193 B.n192 585
R33 B.n191 B.n100 585
R34 B.n190 B.n189 585
R35 B.n188 B.n101 585
R36 B.n187 B.n186 585
R37 B.n185 B.n102 585
R38 B.n184 B.n183 585
R39 B.n182 B.n103 585
R40 B.n181 B.n180 585
R41 B.n179 B.n104 585
R42 B.n178 B.n177 585
R43 B.n176 B.n105 585
R44 B.n175 B.n174 585
R45 B.n173 B.n106 585
R46 B.n246 B.n81 585
R47 B.n248 B.n247 585
R48 B.n249 B.n80 585
R49 B.n251 B.n250 585
R50 B.n252 B.n79 585
R51 B.n254 B.n253 585
R52 B.n255 B.n78 585
R53 B.n257 B.n256 585
R54 B.n258 B.n77 585
R55 B.n260 B.n259 585
R56 B.n261 B.n76 585
R57 B.n263 B.n262 585
R58 B.n264 B.n75 585
R59 B.n266 B.n265 585
R60 B.n267 B.n74 585
R61 B.n269 B.n268 585
R62 B.n270 B.n73 585
R63 B.n272 B.n271 585
R64 B.n273 B.n72 585
R65 B.n275 B.n274 585
R66 B.n276 B.n71 585
R67 B.n278 B.n277 585
R68 B.n279 B.n70 585
R69 B.n281 B.n280 585
R70 B.n282 B.n69 585
R71 B.n284 B.n283 585
R72 B.n285 B.n68 585
R73 B.n287 B.n286 585
R74 B.n288 B.n67 585
R75 B.n290 B.n289 585
R76 B.n291 B.n66 585
R77 B.n293 B.n292 585
R78 B.n294 B.n65 585
R79 B.n296 B.n295 585
R80 B.n297 B.n64 585
R81 B.n299 B.n298 585
R82 B.n300 B.n63 585
R83 B.n302 B.n301 585
R84 B.n303 B.n62 585
R85 B.n305 B.n304 585
R86 B.n306 B.n61 585
R87 B.n308 B.n307 585
R88 B.n309 B.n60 585
R89 B.n311 B.n310 585
R90 B.n312 B.n59 585
R91 B.n314 B.n313 585
R92 B.n315 B.n58 585
R93 B.n317 B.n316 585
R94 B.n318 B.n57 585
R95 B.n320 B.n319 585
R96 B.n321 B.n56 585
R97 B.n323 B.n322 585
R98 B.n324 B.n55 585
R99 B.n326 B.n325 585
R100 B.n327 B.n54 585
R101 B.n329 B.n328 585
R102 B.n330 B.n53 585
R103 B.n332 B.n331 585
R104 B.n333 B.n52 585
R105 B.n335 B.n334 585
R106 B.n336 B.n51 585
R107 B.n338 B.n337 585
R108 B.n339 B.n50 585
R109 B.n341 B.n340 585
R110 B.n342 B.n49 585
R111 B.n344 B.n343 585
R112 B.n345 B.n48 585
R113 B.n347 B.n346 585
R114 B.n348 B.n47 585
R115 B.n350 B.n349 585
R116 B.n420 B.n19 585
R117 B.n419 B.n418 585
R118 B.n417 B.n20 585
R119 B.n416 B.n415 585
R120 B.n414 B.n21 585
R121 B.n413 B.n412 585
R122 B.n411 B.n22 585
R123 B.n410 B.n409 585
R124 B.n408 B.n23 585
R125 B.n407 B.n406 585
R126 B.n405 B.n24 585
R127 B.n404 B.n403 585
R128 B.n402 B.n25 585
R129 B.n401 B.n400 585
R130 B.n399 B.n26 585
R131 B.n398 B.n397 585
R132 B.n396 B.n27 585
R133 B.n395 B.n394 585
R134 B.n393 B.n392 585
R135 B.n391 B.n31 585
R136 B.n390 B.n389 585
R137 B.n388 B.n32 585
R138 B.n387 B.n386 585
R139 B.n385 B.n33 585
R140 B.n384 B.n383 585
R141 B.n382 B.n34 585
R142 B.n381 B.n380 585
R143 B.n379 B.n35 585
R144 B.n377 B.n376 585
R145 B.n375 B.n38 585
R146 B.n374 B.n373 585
R147 B.n372 B.n39 585
R148 B.n371 B.n370 585
R149 B.n369 B.n40 585
R150 B.n368 B.n367 585
R151 B.n366 B.n41 585
R152 B.n365 B.n364 585
R153 B.n363 B.n42 585
R154 B.n362 B.n361 585
R155 B.n360 B.n43 585
R156 B.n359 B.n358 585
R157 B.n357 B.n44 585
R158 B.n356 B.n355 585
R159 B.n354 B.n45 585
R160 B.n353 B.n352 585
R161 B.n351 B.n46 585
R162 B.n422 B.n421 585
R163 B.n423 B.n18 585
R164 B.n425 B.n424 585
R165 B.n426 B.n17 585
R166 B.n428 B.n427 585
R167 B.n429 B.n16 585
R168 B.n431 B.n430 585
R169 B.n432 B.n15 585
R170 B.n434 B.n433 585
R171 B.n435 B.n14 585
R172 B.n437 B.n436 585
R173 B.n438 B.n13 585
R174 B.n440 B.n439 585
R175 B.n441 B.n12 585
R176 B.n443 B.n442 585
R177 B.n444 B.n11 585
R178 B.n446 B.n445 585
R179 B.n447 B.n10 585
R180 B.n449 B.n448 585
R181 B.n450 B.n9 585
R182 B.n452 B.n451 585
R183 B.n453 B.n8 585
R184 B.n455 B.n454 585
R185 B.n456 B.n7 585
R186 B.n458 B.n457 585
R187 B.n459 B.n6 585
R188 B.n461 B.n460 585
R189 B.n462 B.n5 585
R190 B.n464 B.n463 585
R191 B.n465 B.n4 585
R192 B.n467 B.n466 585
R193 B.n468 B.n3 585
R194 B.n470 B.n469 585
R195 B.n471 B.n0 585
R196 B.n2 B.n1 585
R197 B.n124 B.n123 585
R198 B.n125 B.n122 585
R199 B.n127 B.n126 585
R200 B.n128 B.n121 585
R201 B.n130 B.n129 585
R202 B.n131 B.n120 585
R203 B.n133 B.n132 585
R204 B.n134 B.n119 585
R205 B.n136 B.n135 585
R206 B.n137 B.n118 585
R207 B.n139 B.n138 585
R208 B.n140 B.n117 585
R209 B.n142 B.n141 585
R210 B.n143 B.n116 585
R211 B.n145 B.n144 585
R212 B.n146 B.n115 585
R213 B.n148 B.n147 585
R214 B.n149 B.n114 585
R215 B.n151 B.n150 585
R216 B.n152 B.n113 585
R217 B.n154 B.n153 585
R218 B.n155 B.n112 585
R219 B.n157 B.n156 585
R220 B.n158 B.n111 585
R221 B.n160 B.n159 585
R222 B.n161 B.n110 585
R223 B.n163 B.n162 585
R224 B.n164 B.n109 585
R225 B.n166 B.n165 585
R226 B.n167 B.n108 585
R227 B.n169 B.n168 585
R228 B.n170 B.n107 585
R229 B.n172 B.n171 585
R230 B.n173 B.n172 502.111
R231 B.n244 B.n81 502.111
R232 B.n351 B.n350 502.111
R233 B.n422 B.n19 502.111
R234 B.n473 B.n472 256.663
R235 B.n96 B.t6 245.625
R236 B.n214 B.t0 245.625
R237 B.n36 B.t9 245.625
R238 B.n28 B.t3 245.625
R239 B.n472 B.n471 235.042
R240 B.n472 B.n2 235.042
R241 B.n214 B.t1 177.214
R242 B.n36 B.t11 177.214
R243 B.n96 B.t7 177.212
R244 B.n28 B.t5 177.212
R245 B.n174 B.n173 163.367
R246 B.n174 B.n105 163.367
R247 B.n178 B.n105 163.367
R248 B.n179 B.n178 163.367
R249 B.n180 B.n179 163.367
R250 B.n180 B.n103 163.367
R251 B.n184 B.n103 163.367
R252 B.n185 B.n184 163.367
R253 B.n186 B.n185 163.367
R254 B.n186 B.n101 163.367
R255 B.n190 B.n101 163.367
R256 B.n191 B.n190 163.367
R257 B.n192 B.n191 163.367
R258 B.n192 B.n99 163.367
R259 B.n196 B.n99 163.367
R260 B.n197 B.n196 163.367
R261 B.n198 B.n197 163.367
R262 B.n198 B.n95 163.367
R263 B.n203 B.n95 163.367
R264 B.n204 B.n203 163.367
R265 B.n205 B.n204 163.367
R266 B.n205 B.n93 163.367
R267 B.n209 B.n93 163.367
R268 B.n210 B.n209 163.367
R269 B.n211 B.n210 163.367
R270 B.n211 B.n91 163.367
R271 B.n218 B.n91 163.367
R272 B.n219 B.n218 163.367
R273 B.n220 B.n219 163.367
R274 B.n220 B.n89 163.367
R275 B.n224 B.n89 163.367
R276 B.n225 B.n224 163.367
R277 B.n226 B.n225 163.367
R278 B.n226 B.n87 163.367
R279 B.n230 B.n87 163.367
R280 B.n231 B.n230 163.367
R281 B.n232 B.n231 163.367
R282 B.n232 B.n85 163.367
R283 B.n236 B.n85 163.367
R284 B.n237 B.n236 163.367
R285 B.n238 B.n237 163.367
R286 B.n238 B.n83 163.367
R287 B.n242 B.n83 163.367
R288 B.n243 B.n242 163.367
R289 B.n244 B.n243 163.367
R290 B.n350 B.n47 163.367
R291 B.n346 B.n47 163.367
R292 B.n346 B.n345 163.367
R293 B.n345 B.n344 163.367
R294 B.n344 B.n49 163.367
R295 B.n340 B.n49 163.367
R296 B.n340 B.n339 163.367
R297 B.n339 B.n338 163.367
R298 B.n338 B.n51 163.367
R299 B.n334 B.n51 163.367
R300 B.n334 B.n333 163.367
R301 B.n333 B.n332 163.367
R302 B.n332 B.n53 163.367
R303 B.n328 B.n53 163.367
R304 B.n328 B.n327 163.367
R305 B.n327 B.n326 163.367
R306 B.n326 B.n55 163.367
R307 B.n322 B.n55 163.367
R308 B.n322 B.n321 163.367
R309 B.n321 B.n320 163.367
R310 B.n320 B.n57 163.367
R311 B.n316 B.n57 163.367
R312 B.n316 B.n315 163.367
R313 B.n315 B.n314 163.367
R314 B.n314 B.n59 163.367
R315 B.n310 B.n59 163.367
R316 B.n310 B.n309 163.367
R317 B.n309 B.n308 163.367
R318 B.n308 B.n61 163.367
R319 B.n304 B.n61 163.367
R320 B.n304 B.n303 163.367
R321 B.n303 B.n302 163.367
R322 B.n302 B.n63 163.367
R323 B.n298 B.n63 163.367
R324 B.n298 B.n297 163.367
R325 B.n297 B.n296 163.367
R326 B.n296 B.n65 163.367
R327 B.n292 B.n65 163.367
R328 B.n292 B.n291 163.367
R329 B.n291 B.n290 163.367
R330 B.n290 B.n67 163.367
R331 B.n286 B.n67 163.367
R332 B.n286 B.n285 163.367
R333 B.n285 B.n284 163.367
R334 B.n284 B.n69 163.367
R335 B.n280 B.n69 163.367
R336 B.n280 B.n279 163.367
R337 B.n279 B.n278 163.367
R338 B.n278 B.n71 163.367
R339 B.n274 B.n71 163.367
R340 B.n274 B.n273 163.367
R341 B.n273 B.n272 163.367
R342 B.n272 B.n73 163.367
R343 B.n268 B.n73 163.367
R344 B.n268 B.n267 163.367
R345 B.n267 B.n266 163.367
R346 B.n266 B.n75 163.367
R347 B.n262 B.n75 163.367
R348 B.n262 B.n261 163.367
R349 B.n261 B.n260 163.367
R350 B.n260 B.n77 163.367
R351 B.n256 B.n77 163.367
R352 B.n256 B.n255 163.367
R353 B.n255 B.n254 163.367
R354 B.n254 B.n79 163.367
R355 B.n250 B.n79 163.367
R356 B.n250 B.n249 163.367
R357 B.n249 B.n248 163.367
R358 B.n248 B.n81 163.367
R359 B.n418 B.n19 163.367
R360 B.n418 B.n417 163.367
R361 B.n417 B.n416 163.367
R362 B.n416 B.n21 163.367
R363 B.n412 B.n21 163.367
R364 B.n412 B.n411 163.367
R365 B.n411 B.n410 163.367
R366 B.n410 B.n23 163.367
R367 B.n406 B.n23 163.367
R368 B.n406 B.n405 163.367
R369 B.n405 B.n404 163.367
R370 B.n404 B.n25 163.367
R371 B.n400 B.n25 163.367
R372 B.n400 B.n399 163.367
R373 B.n399 B.n398 163.367
R374 B.n398 B.n27 163.367
R375 B.n394 B.n27 163.367
R376 B.n394 B.n393 163.367
R377 B.n393 B.n31 163.367
R378 B.n389 B.n31 163.367
R379 B.n389 B.n388 163.367
R380 B.n388 B.n387 163.367
R381 B.n387 B.n33 163.367
R382 B.n383 B.n33 163.367
R383 B.n383 B.n382 163.367
R384 B.n382 B.n381 163.367
R385 B.n381 B.n35 163.367
R386 B.n376 B.n35 163.367
R387 B.n376 B.n375 163.367
R388 B.n375 B.n374 163.367
R389 B.n374 B.n39 163.367
R390 B.n370 B.n39 163.367
R391 B.n370 B.n369 163.367
R392 B.n369 B.n368 163.367
R393 B.n368 B.n41 163.367
R394 B.n364 B.n41 163.367
R395 B.n364 B.n363 163.367
R396 B.n363 B.n362 163.367
R397 B.n362 B.n43 163.367
R398 B.n358 B.n43 163.367
R399 B.n358 B.n357 163.367
R400 B.n357 B.n356 163.367
R401 B.n356 B.n45 163.367
R402 B.n352 B.n45 163.367
R403 B.n352 B.n351 163.367
R404 B.n423 B.n422 163.367
R405 B.n424 B.n423 163.367
R406 B.n424 B.n17 163.367
R407 B.n428 B.n17 163.367
R408 B.n429 B.n428 163.367
R409 B.n430 B.n429 163.367
R410 B.n430 B.n15 163.367
R411 B.n434 B.n15 163.367
R412 B.n435 B.n434 163.367
R413 B.n436 B.n435 163.367
R414 B.n436 B.n13 163.367
R415 B.n440 B.n13 163.367
R416 B.n441 B.n440 163.367
R417 B.n442 B.n441 163.367
R418 B.n442 B.n11 163.367
R419 B.n446 B.n11 163.367
R420 B.n447 B.n446 163.367
R421 B.n448 B.n447 163.367
R422 B.n448 B.n9 163.367
R423 B.n452 B.n9 163.367
R424 B.n453 B.n452 163.367
R425 B.n454 B.n453 163.367
R426 B.n454 B.n7 163.367
R427 B.n458 B.n7 163.367
R428 B.n459 B.n458 163.367
R429 B.n460 B.n459 163.367
R430 B.n460 B.n5 163.367
R431 B.n464 B.n5 163.367
R432 B.n465 B.n464 163.367
R433 B.n466 B.n465 163.367
R434 B.n466 B.n3 163.367
R435 B.n470 B.n3 163.367
R436 B.n471 B.n470 163.367
R437 B.n124 B.n2 163.367
R438 B.n125 B.n124 163.367
R439 B.n126 B.n125 163.367
R440 B.n126 B.n121 163.367
R441 B.n130 B.n121 163.367
R442 B.n131 B.n130 163.367
R443 B.n132 B.n131 163.367
R444 B.n132 B.n119 163.367
R445 B.n136 B.n119 163.367
R446 B.n137 B.n136 163.367
R447 B.n138 B.n137 163.367
R448 B.n138 B.n117 163.367
R449 B.n142 B.n117 163.367
R450 B.n143 B.n142 163.367
R451 B.n144 B.n143 163.367
R452 B.n144 B.n115 163.367
R453 B.n148 B.n115 163.367
R454 B.n149 B.n148 163.367
R455 B.n150 B.n149 163.367
R456 B.n150 B.n113 163.367
R457 B.n154 B.n113 163.367
R458 B.n155 B.n154 163.367
R459 B.n156 B.n155 163.367
R460 B.n156 B.n111 163.367
R461 B.n160 B.n111 163.367
R462 B.n161 B.n160 163.367
R463 B.n162 B.n161 163.367
R464 B.n162 B.n109 163.367
R465 B.n166 B.n109 163.367
R466 B.n167 B.n166 163.367
R467 B.n168 B.n167 163.367
R468 B.n168 B.n107 163.367
R469 B.n172 B.n107 163.367
R470 B.n215 B.t2 119.615
R471 B.n37 B.t10 119.615
R472 B.n97 B.t8 119.612
R473 B.n29 B.t4 119.612
R474 B.n200 B.n97 59.5399
R475 B.n216 B.n215 59.5399
R476 B.n378 B.n37 59.5399
R477 B.n30 B.n29 59.5399
R478 B.n97 B.n96 57.6005
R479 B.n215 B.n214 57.6005
R480 B.n37 B.n36 57.6005
R481 B.n29 B.n28 57.6005
R482 B.n421 B.n420 32.6249
R483 B.n349 B.n46 32.6249
R484 B.n246 B.n245 32.6249
R485 B.n171 B.n106 32.6249
R486 B B.n473 18.0485
R487 B.n421 B.n18 10.6151
R488 B.n425 B.n18 10.6151
R489 B.n426 B.n425 10.6151
R490 B.n427 B.n426 10.6151
R491 B.n427 B.n16 10.6151
R492 B.n431 B.n16 10.6151
R493 B.n432 B.n431 10.6151
R494 B.n433 B.n432 10.6151
R495 B.n433 B.n14 10.6151
R496 B.n437 B.n14 10.6151
R497 B.n438 B.n437 10.6151
R498 B.n439 B.n438 10.6151
R499 B.n439 B.n12 10.6151
R500 B.n443 B.n12 10.6151
R501 B.n444 B.n443 10.6151
R502 B.n445 B.n444 10.6151
R503 B.n445 B.n10 10.6151
R504 B.n449 B.n10 10.6151
R505 B.n450 B.n449 10.6151
R506 B.n451 B.n450 10.6151
R507 B.n451 B.n8 10.6151
R508 B.n455 B.n8 10.6151
R509 B.n456 B.n455 10.6151
R510 B.n457 B.n456 10.6151
R511 B.n457 B.n6 10.6151
R512 B.n461 B.n6 10.6151
R513 B.n462 B.n461 10.6151
R514 B.n463 B.n462 10.6151
R515 B.n463 B.n4 10.6151
R516 B.n467 B.n4 10.6151
R517 B.n468 B.n467 10.6151
R518 B.n469 B.n468 10.6151
R519 B.n469 B.n0 10.6151
R520 B.n420 B.n419 10.6151
R521 B.n419 B.n20 10.6151
R522 B.n415 B.n20 10.6151
R523 B.n415 B.n414 10.6151
R524 B.n414 B.n413 10.6151
R525 B.n413 B.n22 10.6151
R526 B.n409 B.n22 10.6151
R527 B.n409 B.n408 10.6151
R528 B.n408 B.n407 10.6151
R529 B.n407 B.n24 10.6151
R530 B.n403 B.n24 10.6151
R531 B.n403 B.n402 10.6151
R532 B.n402 B.n401 10.6151
R533 B.n401 B.n26 10.6151
R534 B.n397 B.n26 10.6151
R535 B.n397 B.n396 10.6151
R536 B.n396 B.n395 10.6151
R537 B.n392 B.n391 10.6151
R538 B.n391 B.n390 10.6151
R539 B.n390 B.n32 10.6151
R540 B.n386 B.n32 10.6151
R541 B.n386 B.n385 10.6151
R542 B.n385 B.n384 10.6151
R543 B.n384 B.n34 10.6151
R544 B.n380 B.n34 10.6151
R545 B.n380 B.n379 10.6151
R546 B.n377 B.n38 10.6151
R547 B.n373 B.n38 10.6151
R548 B.n373 B.n372 10.6151
R549 B.n372 B.n371 10.6151
R550 B.n371 B.n40 10.6151
R551 B.n367 B.n40 10.6151
R552 B.n367 B.n366 10.6151
R553 B.n366 B.n365 10.6151
R554 B.n365 B.n42 10.6151
R555 B.n361 B.n42 10.6151
R556 B.n361 B.n360 10.6151
R557 B.n360 B.n359 10.6151
R558 B.n359 B.n44 10.6151
R559 B.n355 B.n44 10.6151
R560 B.n355 B.n354 10.6151
R561 B.n354 B.n353 10.6151
R562 B.n353 B.n46 10.6151
R563 B.n349 B.n348 10.6151
R564 B.n348 B.n347 10.6151
R565 B.n347 B.n48 10.6151
R566 B.n343 B.n48 10.6151
R567 B.n343 B.n342 10.6151
R568 B.n342 B.n341 10.6151
R569 B.n341 B.n50 10.6151
R570 B.n337 B.n50 10.6151
R571 B.n337 B.n336 10.6151
R572 B.n336 B.n335 10.6151
R573 B.n335 B.n52 10.6151
R574 B.n331 B.n52 10.6151
R575 B.n331 B.n330 10.6151
R576 B.n330 B.n329 10.6151
R577 B.n329 B.n54 10.6151
R578 B.n325 B.n54 10.6151
R579 B.n325 B.n324 10.6151
R580 B.n324 B.n323 10.6151
R581 B.n323 B.n56 10.6151
R582 B.n319 B.n56 10.6151
R583 B.n319 B.n318 10.6151
R584 B.n318 B.n317 10.6151
R585 B.n317 B.n58 10.6151
R586 B.n313 B.n58 10.6151
R587 B.n313 B.n312 10.6151
R588 B.n312 B.n311 10.6151
R589 B.n311 B.n60 10.6151
R590 B.n307 B.n60 10.6151
R591 B.n307 B.n306 10.6151
R592 B.n306 B.n305 10.6151
R593 B.n305 B.n62 10.6151
R594 B.n301 B.n62 10.6151
R595 B.n301 B.n300 10.6151
R596 B.n300 B.n299 10.6151
R597 B.n299 B.n64 10.6151
R598 B.n295 B.n64 10.6151
R599 B.n295 B.n294 10.6151
R600 B.n294 B.n293 10.6151
R601 B.n293 B.n66 10.6151
R602 B.n289 B.n66 10.6151
R603 B.n289 B.n288 10.6151
R604 B.n288 B.n287 10.6151
R605 B.n287 B.n68 10.6151
R606 B.n283 B.n68 10.6151
R607 B.n283 B.n282 10.6151
R608 B.n282 B.n281 10.6151
R609 B.n281 B.n70 10.6151
R610 B.n277 B.n70 10.6151
R611 B.n277 B.n276 10.6151
R612 B.n276 B.n275 10.6151
R613 B.n275 B.n72 10.6151
R614 B.n271 B.n72 10.6151
R615 B.n271 B.n270 10.6151
R616 B.n270 B.n269 10.6151
R617 B.n269 B.n74 10.6151
R618 B.n265 B.n74 10.6151
R619 B.n265 B.n264 10.6151
R620 B.n264 B.n263 10.6151
R621 B.n263 B.n76 10.6151
R622 B.n259 B.n76 10.6151
R623 B.n259 B.n258 10.6151
R624 B.n258 B.n257 10.6151
R625 B.n257 B.n78 10.6151
R626 B.n253 B.n78 10.6151
R627 B.n253 B.n252 10.6151
R628 B.n252 B.n251 10.6151
R629 B.n251 B.n80 10.6151
R630 B.n247 B.n80 10.6151
R631 B.n247 B.n246 10.6151
R632 B.n123 B.n1 10.6151
R633 B.n123 B.n122 10.6151
R634 B.n127 B.n122 10.6151
R635 B.n128 B.n127 10.6151
R636 B.n129 B.n128 10.6151
R637 B.n129 B.n120 10.6151
R638 B.n133 B.n120 10.6151
R639 B.n134 B.n133 10.6151
R640 B.n135 B.n134 10.6151
R641 B.n135 B.n118 10.6151
R642 B.n139 B.n118 10.6151
R643 B.n140 B.n139 10.6151
R644 B.n141 B.n140 10.6151
R645 B.n141 B.n116 10.6151
R646 B.n145 B.n116 10.6151
R647 B.n146 B.n145 10.6151
R648 B.n147 B.n146 10.6151
R649 B.n147 B.n114 10.6151
R650 B.n151 B.n114 10.6151
R651 B.n152 B.n151 10.6151
R652 B.n153 B.n152 10.6151
R653 B.n153 B.n112 10.6151
R654 B.n157 B.n112 10.6151
R655 B.n158 B.n157 10.6151
R656 B.n159 B.n158 10.6151
R657 B.n159 B.n110 10.6151
R658 B.n163 B.n110 10.6151
R659 B.n164 B.n163 10.6151
R660 B.n165 B.n164 10.6151
R661 B.n165 B.n108 10.6151
R662 B.n169 B.n108 10.6151
R663 B.n170 B.n169 10.6151
R664 B.n171 B.n170 10.6151
R665 B.n175 B.n106 10.6151
R666 B.n176 B.n175 10.6151
R667 B.n177 B.n176 10.6151
R668 B.n177 B.n104 10.6151
R669 B.n181 B.n104 10.6151
R670 B.n182 B.n181 10.6151
R671 B.n183 B.n182 10.6151
R672 B.n183 B.n102 10.6151
R673 B.n187 B.n102 10.6151
R674 B.n188 B.n187 10.6151
R675 B.n189 B.n188 10.6151
R676 B.n189 B.n100 10.6151
R677 B.n193 B.n100 10.6151
R678 B.n194 B.n193 10.6151
R679 B.n195 B.n194 10.6151
R680 B.n195 B.n98 10.6151
R681 B.n199 B.n98 10.6151
R682 B.n202 B.n201 10.6151
R683 B.n202 B.n94 10.6151
R684 B.n206 B.n94 10.6151
R685 B.n207 B.n206 10.6151
R686 B.n208 B.n207 10.6151
R687 B.n208 B.n92 10.6151
R688 B.n212 B.n92 10.6151
R689 B.n213 B.n212 10.6151
R690 B.n217 B.n213 10.6151
R691 B.n221 B.n90 10.6151
R692 B.n222 B.n221 10.6151
R693 B.n223 B.n222 10.6151
R694 B.n223 B.n88 10.6151
R695 B.n227 B.n88 10.6151
R696 B.n228 B.n227 10.6151
R697 B.n229 B.n228 10.6151
R698 B.n229 B.n86 10.6151
R699 B.n233 B.n86 10.6151
R700 B.n234 B.n233 10.6151
R701 B.n235 B.n234 10.6151
R702 B.n235 B.n84 10.6151
R703 B.n239 B.n84 10.6151
R704 B.n240 B.n239 10.6151
R705 B.n241 B.n240 10.6151
R706 B.n241 B.n82 10.6151
R707 B.n245 B.n82 10.6151
R708 B.n395 B.n30 9.36635
R709 B.n378 B.n377 9.36635
R710 B.n200 B.n199 9.36635
R711 B.n216 B.n90 9.36635
R712 B.n473 B.n0 8.11757
R713 B.n473 B.n1 8.11757
R714 B.n392 B.n30 1.24928
R715 B.n379 B.n378 1.24928
R716 B.n201 B.n200 1.24928
R717 B.n217 B.n216 1.24928
R718 VN.n0 VN.t0 73.996
R719 VN.n1 VN.t1 73.996
R720 VN.n0 VN.t2 73.2135
R721 VN.n1 VN.t3 73.2135
R722 VN VN.n1 45.038
R723 VN VN.n0 4.25389
R724 VDD2.n2 VDD2.n0 141.579
R725 VDD2.n2 VDD2.n1 106.641
R726 VDD2.n1 VDD2.t2 7.90926
R727 VDD2.n1 VDD2.t1 7.90926
R728 VDD2.n0 VDD2.t3 7.90926
R729 VDD2.n0 VDD2.t0 7.90926
R730 VDD2 VDD2.n2 0.0586897
R731 VTAIL.n5 VTAIL.t0 97.8712
R732 VTAIL.n4 VTAIL.t6 97.8712
R733 VTAIL.n3 VTAIL.t4 97.8712
R734 VTAIL.n7 VTAIL.t5 97.8709
R735 VTAIL.n0 VTAIL.t7 97.8709
R736 VTAIL.n1 VTAIL.t2 97.8709
R737 VTAIL.n2 VTAIL.t3 97.8709
R738 VTAIL.n6 VTAIL.t1 97.8709
R739 VTAIL.n7 VTAIL.n6 18.4703
R740 VTAIL.n3 VTAIL.n2 18.4703
R741 VTAIL.n4 VTAIL.n3 2.56084
R742 VTAIL.n6 VTAIL.n5 2.56084
R743 VTAIL.n2 VTAIL.n1 2.56084
R744 VTAIL VTAIL.n0 1.33886
R745 VTAIL VTAIL.n7 1.22248
R746 VTAIL.n5 VTAIL.n4 0.470328
R747 VTAIL.n1 VTAIL.n0 0.470328
R748 VP.n14 VP.n0 161.3
R749 VP.n13 VP.n12 161.3
R750 VP.n11 VP.n1 161.3
R751 VP.n10 VP.n9 161.3
R752 VP.n8 VP.n2 161.3
R753 VP.n7 VP.n6 161.3
R754 VP.n5 VP.n3 99.257
R755 VP.n16 VP.n15 99.257
R756 VP.n4 VP.t1 73.996
R757 VP.n4 VP.t2 73.2135
R758 VP.n9 VP.n1 56.5193
R759 VP.n5 VP.n4 44.7591
R760 VP.n3 VP.t3 37.5198
R761 VP.n15 VP.t0 37.5198
R762 VP.n8 VP.n7 24.4675
R763 VP.n9 VP.n8 24.4675
R764 VP.n13 VP.n1 24.4675
R765 VP.n14 VP.n13 24.4675
R766 VP.n7 VP.n3 11.5
R767 VP.n15 VP.n14 11.5
R768 VP.n6 VP.n5 0.278367
R769 VP.n16 VP.n0 0.278367
R770 VP.n6 VP.n2 0.189894
R771 VP.n10 VP.n2 0.189894
R772 VP.n11 VP.n10 0.189894
R773 VP.n12 VP.n11 0.189894
R774 VP.n12 VP.n0 0.189894
R775 VP VP.n16 0.153454
R776 VDD1 VDD1.n1 142.105
R777 VDD1 VDD1.n0 106.7
R778 VDD1.n0 VDD1.t2 7.90926
R779 VDD1.n0 VDD1.t1 7.90926
R780 VDD1.n1 VDD1.t0 7.90926
R781 VDD1.n1 VDD1.t3 7.90926
C0 w_n2752_n1790# VDD1 1.25058f
C1 w_n2752_n1790# VP 4.86252f
C2 VN B 1.02737f
C3 VTAIL B 2.33335f
C4 VTAIL VN 2.25168f
C5 B VDD1 1.05512f
C6 VP B 1.61463f
C7 w_n2752_n1790# VDD2 1.30722f
C8 VN VDD1 0.153368f
C9 VTAIL VDD1 3.54817f
C10 VP VN 4.76116f
C11 VTAIL VP 2.26579f
C12 VP VDD1 2.08742f
C13 VDD2 B 1.10807f
C14 VDD2 VN 1.84041f
C15 w_n2752_n1790# B 7.09952f
C16 VTAIL VDD2 3.60264f
C17 w_n2752_n1790# VN 4.50938f
C18 w_n2752_n1790# VTAIL 2.1877f
C19 VDD2 VDD1 1.03068f
C20 VP VDD2 0.401619f
C21 VDD2 VSUBS 0.692142f
C22 VDD1 VSUBS 4.702996f
C23 VTAIL VSUBS 0.632764f
C24 VN VSUBS 5.07759f
C25 VP VSUBS 1.851754f
C26 B VSUBS 3.453346f
C27 w_n2752_n1790# VSUBS 61.986f
C28 VDD1.t2 VSUBS 0.092174f
C29 VDD1.t1 VSUBS 0.092174f
C30 VDD1.n0 VSUBS 0.543506f
C31 VDD1.t0 VSUBS 0.092174f
C32 VDD1.t3 VSUBS 0.092174f
C33 VDD1.n1 VSUBS 0.90616f
C34 VP.n0 VSUBS 0.064192f
C35 VP.t0 VSUBS 1.36046f
C36 VP.n1 VSUBS 0.071077f
C37 VP.n2 VSUBS 0.048689f
C38 VP.t3 VSUBS 1.36046f
C39 VP.n3 VSUBS 0.708647f
C40 VP.t2 VSUBS 1.77568f
C41 VP.t1 VSUBS 1.78442f
C42 VP.n4 VSUBS 3.24872f
C43 VP.n5 VSUBS 2.22726f
C44 VP.n6 VSUBS 0.064192f
C45 VP.n7 VSUBS 0.066998f
C46 VP.n8 VSUBS 0.090744f
C47 VP.n9 VSUBS 0.071077f
C48 VP.n10 VSUBS 0.048689f
C49 VP.n11 VSUBS 0.048689f
C50 VP.n12 VSUBS 0.048689f
C51 VP.n13 VSUBS 0.090744f
C52 VP.n14 VSUBS 0.066998f
C53 VP.n15 VSUBS 0.708646f
C54 VP.n16 VSUBS 0.077802f
C55 VTAIL.t7 VSUBS 0.717491f
C56 VTAIL.n0 VSUBS 0.705115f
C57 VTAIL.t2 VSUBS 0.717491f
C58 VTAIL.n1 VSUBS 0.824874f
C59 VTAIL.t3 VSUBS 0.717491f
C60 VTAIL.n2 VSUBS 1.79014f
C61 VTAIL.t4 VSUBS 0.717494f
C62 VTAIL.n3 VSUBS 1.79014f
C63 VTAIL.t6 VSUBS 0.717494f
C64 VTAIL.n4 VSUBS 0.824872f
C65 VTAIL.t0 VSUBS 0.717494f
C66 VTAIL.n5 VSUBS 0.824872f
C67 VTAIL.t1 VSUBS 0.717492f
C68 VTAIL.n6 VSUBS 1.79014f
C69 VTAIL.t5 VSUBS 0.717491f
C70 VTAIL.n7 VSUBS 1.65898f
C71 VDD2.t3 VSUBS 0.060385f
C72 VDD2.t0 VSUBS 0.060385f
C73 VDD2.n0 VSUBS 0.581729f
C74 VDD2.t2 VSUBS 0.060385f
C75 VDD2.t1 VSUBS 0.060385f
C76 VDD2.n1 VSUBS 0.355827f
C77 VDD2.n2 VSUBS 2.26352f
C78 VN.t0 VSUBS 1.46094f
C79 VN.t2 VSUBS 1.45378f
C80 VN.n0 VSUBS 0.891577f
C81 VN.t1 VSUBS 1.46094f
C82 VN.t3 VSUBS 1.45378f
C83 VN.n1 VSUBS 2.68108f
C84 B.n0 VSUBS 0.008128f
C85 B.n1 VSUBS 0.008128f
C86 B.n2 VSUBS 0.012021f
C87 B.n3 VSUBS 0.009212f
C88 B.n4 VSUBS 0.009212f
C89 B.n5 VSUBS 0.009212f
C90 B.n6 VSUBS 0.009212f
C91 B.n7 VSUBS 0.009212f
C92 B.n8 VSUBS 0.009212f
C93 B.n9 VSUBS 0.009212f
C94 B.n10 VSUBS 0.009212f
C95 B.n11 VSUBS 0.009212f
C96 B.n12 VSUBS 0.009212f
C97 B.n13 VSUBS 0.009212f
C98 B.n14 VSUBS 0.009212f
C99 B.n15 VSUBS 0.009212f
C100 B.n16 VSUBS 0.009212f
C101 B.n17 VSUBS 0.009212f
C102 B.n18 VSUBS 0.009212f
C103 B.n19 VSUBS 0.021712f
C104 B.n20 VSUBS 0.009212f
C105 B.n21 VSUBS 0.009212f
C106 B.n22 VSUBS 0.009212f
C107 B.n23 VSUBS 0.009212f
C108 B.n24 VSUBS 0.009212f
C109 B.n25 VSUBS 0.009212f
C110 B.n26 VSUBS 0.009212f
C111 B.n27 VSUBS 0.009212f
C112 B.t4 VSUBS 0.143449f
C113 B.t5 VSUBS 0.168586f
C114 B.t3 VSUBS 0.686719f
C115 B.n28 VSUBS 0.122054f
C116 B.n29 VSUBS 0.090475f
C117 B.n30 VSUBS 0.021342f
C118 B.n31 VSUBS 0.009212f
C119 B.n32 VSUBS 0.009212f
C120 B.n33 VSUBS 0.009212f
C121 B.n34 VSUBS 0.009212f
C122 B.n35 VSUBS 0.009212f
C123 B.t10 VSUBS 0.143449f
C124 B.t11 VSUBS 0.168586f
C125 B.t9 VSUBS 0.686719f
C126 B.n36 VSUBS 0.122055f
C127 B.n37 VSUBS 0.090475f
C128 B.n38 VSUBS 0.009212f
C129 B.n39 VSUBS 0.009212f
C130 B.n40 VSUBS 0.009212f
C131 B.n41 VSUBS 0.009212f
C132 B.n42 VSUBS 0.009212f
C133 B.n43 VSUBS 0.009212f
C134 B.n44 VSUBS 0.009212f
C135 B.n45 VSUBS 0.009212f
C136 B.n46 VSUBS 0.021712f
C137 B.n47 VSUBS 0.009212f
C138 B.n48 VSUBS 0.009212f
C139 B.n49 VSUBS 0.009212f
C140 B.n50 VSUBS 0.009212f
C141 B.n51 VSUBS 0.009212f
C142 B.n52 VSUBS 0.009212f
C143 B.n53 VSUBS 0.009212f
C144 B.n54 VSUBS 0.009212f
C145 B.n55 VSUBS 0.009212f
C146 B.n56 VSUBS 0.009212f
C147 B.n57 VSUBS 0.009212f
C148 B.n58 VSUBS 0.009212f
C149 B.n59 VSUBS 0.009212f
C150 B.n60 VSUBS 0.009212f
C151 B.n61 VSUBS 0.009212f
C152 B.n62 VSUBS 0.009212f
C153 B.n63 VSUBS 0.009212f
C154 B.n64 VSUBS 0.009212f
C155 B.n65 VSUBS 0.009212f
C156 B.n66 VSUBS 0.009212f
C157 B.n67 VSUBS 0.009212f
C158 B.n68 VSUBS 0.009212f
C159 B.n69 VSUBS 0.009212f
C160 B.n70 VSUBS 0.009212f
C161 B.n71 VSUBS 0.009212f
C162 B.n72 VSUBS 0.009212f
C163 B.n73 VSUBS 0.009212f
C164 B.n74 VSUBS 0.009212f
C165 B.n75 VSUBS 0.009212f
C166 B.n76 VSUBS 0.009212f
C167 B.n77 VSUBS 0.009212f
C168 B.n78 VSUBS 0.009212f
C169 B.n79 VSUBS 0.009212f
C170 B.n80 VSUBS 0.009212f
C171 B.n81 VSUBS 0.021366f
C172 B.n82 VSUBS 0.009212f
C173 B.n83 VSUBS 0.009212f
C174 B.n84 VSUBS 0.009212f
C175 B.n85 VSUBS 0.009212f
C176 B.n86 VSUBS 0.009212f
C177 B.n87 VSUBS 0.009212f
C178 B.n88 VSUBS 0.009212f
C179 B.n89 VSUBS 0.009212f
C180 B.n90 VSUBS 0.00867f
C181 B.n91 VSUBS 0.009212f
C182 B.n92 VSUBS 0.009212f
C183 B.n93 VSUBS 0.009212f
C184 B.n94 VSUBS 0.009212f
C185 B.n95 VSUBS 0.009212f
C186 B.t8 VSUBS 0.143449f
C187 B.t7 VSUBS 0.168586f
C188 B.t6 VSUBS 0.686719f
C189 B.n96 VSUBS 0.122054f
C190 B.n97 VSUBS 0.090475f
C191 B.n98 VSUBS 0.009212f
C192 B.n99 VSUBS 0.009212f
C193 B.n100 VSUBS 0.009212f
C194 B.n101 VSUBS 0.009212f
C195 B.n102 VSUBS 0.009212f
C196 B.n103 VSUBS 0.009212f
C197 B.n104 VSUBS 0.009212f
C198 B.n105 VSUBS 0.009212f
C199 B.n106 VSUBS 0.021712f
C200 B.n107 VSUBS 0.009212f
C201 B.n108 VSUBS 0.009212f
C202 B.n109 VSUBS 0.009212f
C203 B.n110 VSUBS 0.009212f
C204 B.n111 VSUBS 0.009212f
C205 B.n112 VSUBS 0.009212f
C206 B.n113 VSUBS 0.009212f
C207 B.n114 VSUBS 0.009212f
C208 B.n115 VSUBS 0.009212f
C209 B.n116 VSUBS 0.009212f
C210 B.n117 VSUBS 0.009212f
C211 B.n118 VSUBS 0.009212f
C212 B.n119 VSUBS 0.009212f
C213 B.n120 VSUBS 0.009212f
C214 B.n121 VSUBS 0.009212f
C215 B.n122 VSUBS 0.009212f
C216 B.n123 VSUBS 0.009212f
C217 B.n124 VSUBS 0.009212f
C218 B.n125 VSUBS 0.009212f
C219 B.n126 VSUBS 0.009212f
C220 B.n127 VSUBS 0.009212f
C221 B.n128 VSUBS 0.009212f
C222 B.n129 VSUBS 0.009212f
C223 B.n130 VSUBS 0.009212f
C224 B.n131 VSUBS 0.009212f
C225 B.n132 VSUBS 0.009212f
C226 B.n133 VSUBS 0.009212f
C227 B.n134 VSUBS 0.009212f
C228 B.n135 VSUBS 0.009212f
C229 B.n136 VSUBS 0.009212f
C230 B.n137 VSUBS 0.009212f
C231 B.n138 VSUBS 0.009212f
C232 B.n139 VSUBS 0.009212f
C233 B.n140 VSUBS 0.009212f
C234 B.n141 VSUBS 0.009212f
C235 B.n142 VSUBS 0.009212f
C236 B.n143 VSUBS 0.009212f
C237 B.n144 VSUBS 0.009212f
C238 B.n145 VSUBS 0.009212f
C239 B.n146 VSUBS 0.009212f
C240 B.n147 VSUBS 0.009212f
C241 B.n148 VSUBS 0.009212f
C242 B.n149 VSUBS 0.009212f
C243 B.n150 VSUBS 0.009212f
C244 B.n151 VSUBS 0.009212f
C245 B.n152 VSUBS 0.009212f
C246 B.n153 VSUBS 0.009212f
C247 B.n154 VSUBS 0.009212f
C248 B.n155 VSUBS 0.009212f
C249 B.n156 VSUBS 0.009212f
C250 B.n157 VSUBS 0.009212f
C251 B.n158 VSUBS 0.009212f
C252 B.n159 VSUBS 0.009212f
C253 B.n160 VSUBS 0.009212f
C254 B.n161 VSUBS 0.009212f
C255 B.n162 VSUBS 0.009212f
C256 B.n163 VSUBS 0.009212f
C257 B.n164 VSUBS 0.009212f
C258 B.n165 VSUBS 0.009212f
C259 B.n166 VSUBS 0.009212f
C260 B.n167 VSUBS 0.009212f
C261 B.n168 VSUBS 0.009212f
C262 B.n169 VSUBS 0.009212f
C263 B.n170 VSUBS 0.009212f
C264 B.n171 VSUBS 0.021366f
C265 B.n172 VSUBS 0.021366f
C266 B.n173 VSUBS 0.021712f
C267 B.n174 VSUBS 0.009212f
C268 B.n175 VSUBS 0.009212f
C269 B.n176 VSUBS 0.009212f
C270 B.n177 VSUBS 0.009212f
C271 B.n178 VSUBS 0.009212f
C272 B.n179 VSUBS 0.009212f
C273 B.n180 VSUBS 0.009212f
C274 B.n181 VSUBS 0.009212f
C275 B.n182 VSUBS 0.009212f
C276 B.n183 VSUBS 0.009212f
C277 B.n184 VSUBS 0.009212f
C278 B.n185 VSUBS 0.009212f
C279 B.n186 VSUBS 0.009212f
C280 B.n187 VSUBS 0.009212f
C281 B.n188 VSUBS 0.009212f
C282 B.n189 VSUBS 0.009212f
C283 B.n190 VSUBS 0.009212f
C284 B.n191 VSUBS 0.009212f
C285 B.n192 VSUBS 0.009212f
C286 B.n193 VSUBS 0.009212f
C287 B.n194 VSUBS 0.009212f
C288 B.n195 VSUBS 0.009212f
C289 B.n196 VSUBS 0.009212f
C290 B.n197 VSUBS 0.009212f
C291 B.n198 VSUBS 0.009212f
C292 B.n199 VSUBS 0.00867f
C293 B.n200 VSUBS 0.021342f
C294 B.n201 VSUBS 0.005148f
C295 B.n202 VSUBS 0.009212f
C296 B.n203 VSUBS 0.009212f
C297 B.n204 VSUBS 0.009212f
C298 B.n205 VSUBS 0.009212f
C299 B.n206 VSUBS 0.009212f
C300 B.n207 VSUBS 0.009212f
C301 B.n208 VSUBS 0.009212f
C302 B.n209 VSUBS 0.009212f
C303 B.n210 VSUBS 0.009212f
C304 B.n211 VSUBS 0.009212f
C305 B.n212 VSUBS 0.009212f
C306 B.n213 VSUBS 0.009212f
C307 B.t2 VSUBS 0.143449f
C308 B.t1 VSUBS 0.168586f
C309 B.t0 VSUBS 0.686719f
C310 B.n214 VSUBS 0.122055f
C311 B.n215 VSUBS 0.090475f
C312 B.n216 VSUBS 0.021342f
C313 B.n217 VSUBS 0.005148f
C314 B.n218 VSUBS 0.009212f
C315 B.n219 VSUBS 0.009212f
C316 B.n220 VSUBS 0.009212f
C317 B.n221 VSUBS 0.009212f
C318 B.n222 VSUBS 0.009212f
C319 B.n223 VSUBS 0.009212f
C320 B.n224 VSUBS 0.009212f
C321 B.n225 VSUBS 0.009212f
C322 B.n226 VSUBS 0.009212f
C323 B.n227 VSUBS 0.009212f
C324 B.n228 VSUBS 0.009212f
C325 B.n229 VSUBS 0.009212f
C326 B.n230 VSUBS 0.009212f
C327 B.n231 VSUBS 0.009212f
C328 B.n232 VSUBS 0.009212f
C329 B.n233 VSUBS 0.009212f
C330 B.n234 VSUBS 0.009212f
C331 B.n235 VSUBS 0.009212f
C332 B.n236 VSUBS 0.009212f
C333 B.n237 VSUBS 0.009212f
C334 B.n238 VSUBS 0.009212f
C335 B.n239 VSUBS 0.009212f
C336 B.n240 VSUBS 0.009212f
C337 B.n241 VSUBS 0.009212f
C338 B.n242 VSUBS 0.009212f
C339 B.n243 VSUBS 0.009212f
C340 B.n244 VSUBS 0.021712f
C341 B.n245 VSUBS 0.020622f
C342 B.n246 VSUBS 0.022456f
C343 B.n247 VSUBS 0.009212f
C344 B.n248 VSUBS 0.009212f
C345 B.n249 VSUBS 0.009212f
C346 B.n250 VSUBS 0.009212f
C347 B.n251 VSUBS 0.009212f
C348 B.n252 VSUBS 0.009212f
C349 B.n253 VSUBS 0.009212f
C350 B.n254 VSUBS 0.009212f
C351 B.n255 VSUBS 0.009212f
C352 B.n256 VSUBS 0.009212f
C353 B.n257 VSUBS 0.009212f
C354 B.n258 VSUBS 0.009212f
C355 B.n259 VSUBS 0.009212f
C356 B.n260 VSUBS 0.009212f
C357 B.n261 VSUBS 0.009212f
C358 B.n262 VSUBS 0.009212f
C359 B.n263 VSUBS 0.009212f
C360 B.n264 VSUBS 0.009212f
C361 B.n265 VSUBS 0.009212f
C362 B.n266 VSUBS 0.009212f
C363 B.n267 VSUBS 0.009212f
C364 B.n268 VSUBS 0.009212f
C365 B.n269 VSUBS 0.009212f
C366 B.n270 VSUBS 0.009212f
C367 B.n271 VSUBS 0.009212f
C368 B.n272 VSUBS 0.009212f
C369 B.n273 VSUBS 0.009212f
C370 B.n274 VSUBS 0.009212f
C371 B.n275 VSUBS 0.009212f
C372 B.n276 VSUBS 0.009212f
C373 B.n277 VSUBS 0.009212f
C374 B.n278 VSUBS 0.009212f
C375 B.n279 VSUBS 0.009212f
C376 B.n280 VSUBS 0.009212f
C377 B.n281 VSUBS 0.009212f
C378 B.n282 VSUBS 0.009212f
C379 B.n283 VSUBS 0.009212f
C380 B.n284 VSUBS 0.009212f
C381 B.n285 VSUBS 0.009212f
C382 B.n286 VSUBS 0.009212f
C383 B.n287 VSUBS 0.009212f
C384 B.n288 VSUBS 0.009212f
C385 B.n289 VSUBS 0.009212f
C386 B.n290 VSUBS 0.009212f
C387 B.n291 VSUBS 0.009212f
C388 B.n292 VSUBS 0.009212f
C389 B.n293 VSUBS 0.009212f
C390 B.n294 VSUBS 0.009212f
C391 B.n295 VSUBS 0.009212f
C392 B.n296 VSUBS 0.009212f
C393 B.n297 VSUBS 0.009212f
C394 B.n298 VSUBS 0.009212f
C395 B.n299 VSUBS 0.009212f
C396 B.n300 VSUBS 0.009212f
C397 B.n301 VSUBS 0.009212f
C398 B.n302 VSUBS 0.009212f
C399 B.n303 VSUBS 0.009212f
C400 B.n304 VSUBS 0.009212f
C401 B.n305 VSUBS 0.009212f
C402 B.n306 VSUBS 0.009212f
C403 B.n307 VSUBS 0.009212f
C404 B.n308 VSUBS 0.009212f
C405 B.n309 VSUBS 0.009212f
C406 B.n310 VSUBS 0.009212f
C407 B.n311 VSUBS 0.009212f
C408 B.n312 VSUBS 0.009212f
C409 B.n313 VSUBS 0.009212f
C410 B.n314 VSUBS 0.009212f
C411 B.n315 VSUBS 0.009212f
C412 B.n316 VSUBS 0.009212f
C413 B.n317 VSUBS 0.009212f
C414 B.n318 VSUBS 0.009212f
C415 B.n319 VSUBS 0.009212f
C416 B.n320 VSUBS 0.009212f
C417 B.n321 VSUBS 0.009212f
C418 B.n322 VSUBS 0.009212f
C419 B.n323 VSUBS 0.009212f
C420 B.n324 VSUBS 0.009212f
C421 B.n325 VSUBS 0.009212f
C422 B.n326 VSUBS 0.009212f
C423 B.n327 VSUBS 0.009212f
C424 B.n328 VSUBS 0.009212f
C425 B.n329 VSUBS 0.009212f
C426 B.n330 VSUBS 0.009212f
C427 B.n331 VSUBS 0.009212f
C428 B.n332 VSUBS 0.009212f
C429 B.n333 VSUBS 0.009212f
C430 B.n334 VSUBS 0.009212f
C431 B.n335 VSUBS 0.009212f
C432 B.n336 VSUBS 0.009212f
C433 B.n337 VSUBS 0.009212f
C434 B.n338 VSUBS 0.009212f
C435 B.n339 VSUBS 0.009212f
C436 B.n340 VSUBS 0.009212f
C437 B.n341 VSUBS 0.009212f
C438 B.n342 VSUBS 0.009212f
C439 B.n343 VSUBS 0.009212f
C440 B.n344 VSUBS 0.009212f
C441 B.n345 VSUBS 0.009212f
C442 B.n346 VSUBS 0.009212f
C443 B.n347 VSUBS 0.009212f
C444 B.n348 VSUBS 0.009212f
C445 B.n349 VSUBS 0.021366f
C446 B.n350 VSUBS 0.021366f
C447 B.n351 VSUBS 0.021712f
C448 B.n352 VSUBS 0.009212f
C449 B.n353 VSUBS 0.009212f
C450 B.n354 VSUBS 0.009212f
C451 B.n355 VSUBS 0.009212f
C452 B.n356 VSUBS 0.009212f
C453 B.n357 VSUBS 0.009212f
C454 B.n358 VSUBS 0.009212f
C455 B.n359 VSUBS 0.009212f
C456 B.n360 VSUBS 0.009212f
C457 B.n361 VSUBS 0.009212f
C458 B.n362 VSUBS 0.009212f
C459 B.n363 VSUBS 0.009212f
C460 B.n364 VSUBS 0.009212f
C461 B.n365 VSUBS 0.009212f
C462 B.n366 VSUBS 0.009212f
C463 B.n367 VSUBS 0.009212f
C464 B.n368 VSUBS 0.009212f
C465 B.n369 VSUBS 0.009212f
C466 B.n370 VSUBS 0.009212f
C467 B.n371 VSUBS 0.009212f
C468 B.n372 VSUBS 0.009212f
C469 B.n373 VSUBS 0.009212f
C470 B.n374 VSUBS 0.009212f
C471 B.n375 VSUBS 0.009212f
C472 B.n376 VSUBS 0.009212f
C473 B.n377 VSUBS 0.00867f
C474 B.n378 VSUBS 0.021342f
C475 B.n379 VSUBS 0.005148f
C476 B.n380 VSUBS 0.009212f
C477 B.n381 VSUBS 0.009212f
C478 B.n382 VSUBS 0.009212f
C479 B.n383 VSUBS 0.009212f
C480 B.n384 VSUBS 0.009212f
C481 B.n385 VSUBS 0.009212f
C482 B.n386 VSUBS 0.009212f
C483 B.n387 VSUBS 0.009212f
C484 B.n388 VSUBS 0.009212f
C485 B.n389 VSUBS 0.009212f
C486 B.n390 VSUBS 0.009212f
C487 B.n391 VSUBS 0.009212f
C488 B.n392 VSUBS 0.005148f
C489 B.n393 VSUBS 0.009212f
C490 B.n394 VSUBS 0.009212f
C491 B.n395 VSUBS 0.00867f
C492 B.n396 VSUBS 0.009212f
C493 B.n397 VSUBS 0.009212f
C494 B.n398 VSUBS 0.009212f
C495 B.n399 VSUBS 0.009212f
C496 B.n400 VSUBS 0.009212f
C497 B.n401 VSUBS 0.009212f
C498 B.n402 VSUBS 0.009212f
C499 B.n403 VSUBS 0.009212f
C500 B.n404 VSUBS 0.009212f
C501 B.n405 VSUBS 0.009212f
C502 B.n406 VSUBS 0.009212f
C503 B.n407 VSUBS 0.009212f
C504 B.n408 VSUBS 0.009212f
C505 B.n409 VSUBS 0.009212f
C506 B.n410 VSUBS 0.009212f
C507 B.n411 VSUBS 0.009212f
C508 B.n412 VSUBS 0.009212f
C509 B.n413 VSUBS 0.009212f
C510 B.n414 VSUBS 0.009212f
C511 B.n415 VSUBS 0.009212f
C512 B.n416 VSUBS 0.009212f
C513 B.n417 VSUBS 0.009212f
C514 B.n418 VSUBS 0.009212f
C515 B.n419 VSUBS 0.009212f
C516 B.n420 VSUBS 0.021712f
C517 B.n421 VSUBS 0.021366f
C518 B.n422 VSUBS 0.021366f
C519 B.n423 VSUBS 0.009212f
C520 B.n424 VSUBS 0.009212f
C521 B.n425 VSUBS 0.009212f
C522 B.n426 VSUBS 0.009212f
C523 B.n427 VSUBS 0.009212f
C524 B.n428 VSUBS 0.009212f
C525 B.n429 VSUBS 0.009212f
C526 B.n430 VSUBS 0.009212f
C527 B.n431 VSUBS 0.009212f
C528 B.n432 VSUBS 0.009212f
C529 B.n433 VSUBS 0.009212f
C530 B.n434 VSUBS 0.009212f
C531 B.n435 VSUBS 0.009212f
C532 B.n436 VSUBS 0.009212f
C533 B.n437 VSUBS 0.009212f
C534 B.n438 VSUBS 0.009212f
C535 B.n439 VSUBS 0.009212f
C536 B.n440 VSUBS 0.009212f
C537 B.n441 VSUBS 0.009212f
C538 B.n442 VSUBS 0.009212f
C539 B.n443 VSUBS 0.009212f
C540 B.n444 VSUBS 0.009212f
C541 B.n445 VSUBS 0.009212f
C542 B.n446 VSUBS 0.009212f
C543 B.n447 VSUBS 0.009212f
C544 B.n448 VSUBS 0.009212f
C545 B.n449 VSUBS 0.009212f
C546 B.n450 VSUBS 0.009212f
C547 B.n451 VSUBS 0.009212f
C548 B.n452 VSUBS 0.009212f
C549 B.n453 VSUBS 0.009212f
C550 B.n454 VSUBS 0.009212f
C551 B.n455 VSUBS 0.009212f
C552 B.n456 VSUBS 0.009212f
C553 B.n457 VSUBS 0.009212f
C554 B.n458 VSUBS 0.009212f
C555 B.n459 VSUBS 0.009212f
C556 B.n460 VSUBS 0.009212f
C557 B.n461 VSUBS 0.009212f
C558 B.n462 VSUBS 0.009212f
C559 B.n463 VSUBS 0.009212f
C560 B.n464 VSUBS 0.009212f
C561 B.n465 VSUBS 0.009212f
C562 B.n466 VSUBS 0.009212f
C563 B.n467 VSUBS 0.009212f
C564 B.n468 VSUBS 0.009212f
C565 B.n469 VSUBS 0.009212f
C566 B.n470 VSUBS 0.009212f
C567 B.n471 VSUBS 0.012021f
C568 B.n472 VSUBS 0.012805f
C569 B.n473 VSUBS 0.025464f
.ends

