* NGSPICE file created from diff_pair_sample_1330.ext - technology: sky130A

.subckt diff_pair_sample_1330 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t5 VN.t0 VTAIL.t11 B.t0 sky130_fd_pr__nfet_01v8 ad=1.2285 pd=7.08 as=0.51975 ps=3.48 w=3.15 l=2.44
X1 VDD1.t5 VP.t0 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.51975 pd=3.48 as=1.2285 ps=7.08 w=3.15 l=2.44
X2 B.t19 B.t17 B.t18 B.t11 sky130_fd_pr__nfet_01v8 ad=1.2285 pd=7.08 as=0 ps=0 w=3.15 l=2.44
X3 VTAIL.t3 VP.t1 VDD1.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=0.51975 pd=3.48 as=0.51975 ps=3.48 w=3.15 l=2.44
X4 VDD1.t3 VP.t2 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.2285 pd=7.08 as=0.51975 ps=3.48 w=3.15 l=2.44
X5 B.t16 B.t14 B.t15 B.t7 sky130_fd_pr__nfet_01v8 ad=1.2285 pd=7.08 as=0 ps=0 w=3.15 l=2.44
X6 VDD2.t4 VN.t1 VTAIL.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=0.51975 pd=3.48 as=1.2285 ps=7.08 w=3.15 l=2.44
X7 VTAIL.t7 VN.t2 VDD2.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.51975 pd=3.48 as=0.51975 ps=3.48 w=3.15 l=2.44
X8 VDD2.t2 VN.t3 VTAIL.t10 B.t2 sky130_fd_pr__nfet_01v8 ad=0.51975 pd=3.48 as=1.2285 ps=7.08 w=3.15 l=2.44
X9 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=1.2285 pd=7.08 as=0 ps=0 w=3.15 l=2.44
X10 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=1.2285 pd=7.08 as=0 ps=0 w=3.15 l=2.44
X11 VTAIL.t5 VP.t3 VDD1.t2 B.t5 sky130_fd_pr__nfet_01v8 ad=0.51975 pd=3.48 as=0.51975 ps=3.48 w=3.15 l=2.44
X12 VDD2.t1 VN.t4 VTAIL.t9 B.t4 sky130_fd_pr__nfet_01v8 ad=1.2285 pd=7.08 as=0.51975 ps=3.48 w=3.15 l=2.44
X13 VDD1.t1 VP.t4 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.2285 pd=7.08 as=0.51975 ps=3.48 w=3.15 l=2.44
X14 VDD1.t0 VP.t5 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.51975 pd=3.48 as=1.2285 ps=7.08 w=3.15 l=2.44
X15 VTAIL.t8 VN.t5 VDD2.t0 B.t5 sky130_fd_pr__nfet_01v8 ad=0.51975 pd=3.48 as=0.51975 ps=3.48 w=3.15 l=2.44
R0 VN.n25 VN.n14 161.3
R1 VN.n24 VN.n23 161.3
R2 VN.n22 VN.n15 161.3
R3 VN.n21 VN.n20 161.3
R4 VN.n19 VN.n16 161.3
R5 VN.n11 VN.n0 161.3
R6 VN.n10 VN.n9 161.3
R7 VN.n8 VN.n1 161.3
R8 VN.n7 VN.n6 161.3
R9 VN.n5 VN.n2 161.3
R10 VN.n13 VN.n12 97.5443
R11 VN.n27 VN.n26 97.5443
R12 VN.n3 VN.t0 65.7772
R13 VN.n17 VN.t3 65.7772
R14 VN.n6 VN.n1 51.663
R15 VN.n20 VN.n15 51.663
R16 VN.n4 VN.n3 48.034
R17 VN.n18 VN.n17 48.034
R18 VN VN.n27 41.6535
R19 VN.n4 VN.t5 31.1132
R20 VN.n12 VN.t1 31.1132
R21 VN.n18 VN.t2 31.1132
R22 VN.n26 VN.t4 31.1132
R23 VN.n10 VN.n1 29.3238
R24 VN.n24 VN.n15 29.3238
R25 VN.n5 VN.n4 24.4675
R26 VN.n6 VN.n5 24.4675
R27 VN.n11 VN.n10 24.4675
R28 VN.n20 VN.n19 24.4675
R29 VN.n19 VN.n18 24.4675
R30 VN.n25 VN.n24 24.4675
R31 VN.n12 VN.n11 13.2127
R32 VN.n26 VN.n25 13.2127
R33 VN.n17 VN.n16 6.62503
R34 VN.n3 VN.n2 6.62503
R35 VN.n27 VN.n14 0.278367
R36 VN.n13 VN.n0 0.278367
R37 VN.n23 VN.n14 0.189894
R38 VN.n23 VN.n22 0.189894
R39 VN.n22 VN.n21 0.189894
R40 VN.n21 VN.n16 0.189894
R41 VN.n7 VN.n2 0.189894
R42 VN.n8 VN.n7 0.189894
R43 VN.n9 VN.n8 0.189894
R44 VN.n9 VN.n0 0.189894
R45 VN VN.n13 0.153454
R46 VTAIL.n66 VTAIL.n56 289.615
R47 VTAIL.n12 VTAIL.n2 289.615
R48 VTAIL.n50 VTAIL.n40 289.615
R49 VTAIL.n32 VTAIL.n22 289.615
R50 VTAIL.n60 VTAIL.n59 185
R51 VTAIL.n65 VTAIL.n64 185
R52 VTAIL.n67 VTAIL.n66 185
R53 VTAIL.n6 VTAIL.n5 185
R54 VTAIL.n11 VTAIL.n10 185
R55 VTAIL.n13 VTAIL.n12 185
R56 VTAIL.n51 VTAIL.n50 185
R57 VTAIL.n49 VTAIL.n48 185
R58 VTAIL.n44 VTAIL.n43 185
R59 VTAIL.n33 VTAIL.n32 185
R60 VTAIL.n31 VTAIL.n30 185
R61 VTAIL.n26 VTAIL.n25 185
R62 VTAIL.n61 VTAIL.t6 148.606
R63 VTAIL.n7 VTAIL.t2 148.606
R64 VTAIL.n45 VTAIL.t1 148.606
R65 VTAIL.n27 VTAIL.t10 148.606
R66 VTAIL.n65 VTAIL.n59 104.615
R67 VTAIL.n66 VTAIL.n65 104.615
R68 VTAIL.n11 VTAIL.n5 104.615
R69 VTAIL.n12 VTAIL.n11 104.615
R70 VTAIL.n50 VTAIL.n49 104.615
R71 VTAIL.n49 VTAIL.n43 104.615
R72 VTAIL.n32 VTAIL.n31 104.615
R73 VTAIL.n31 VTAIL.n25 104.615
R74 VTAIL.n39 VTAIL.n38 61.6522
R75 VTAIL.n21 VTAIL.n20 61.6522
R76 VTAIL.n1 VTAIL.n0 61.6521
R77 VTAIL.n19 VTAIL.n18 61.6521
R78 VTAIL.t6 VTAIL.n59 52.3082
R79 VTAIL.t2 VTAIL.n5 52.3082
R80 VTAIL.t1 VTAIL.n43 52.3082
R81 VTAIL.t10 VTAIL.n25 52.3082
R82 VTAIL.n71 VTAIL.n70 32.7672
R83 VTAIL.n17 VTAIL.n16 32.7672
R84 VTAIL.n55 VTAIL.n54 32.7672
R85 VTAIL.n37 VTAIL.n36 32.7672
R86 VTAIL.n21 VTAIL.n19 19.8583
R87 VTAIL.n71 VTAIL.n55 17.4703
R88 VTAIL.n61 VTAIL.n60 15.5966
R89 VTAIL.n7 VTAIL.n6 15.5966
R90 VTAIL.n45 VTAIL.n44 15.5966
R91 VTAIL.n27 VTAIL.n26 15.5966
R92 VTAIL.n64 VTAIL.n63 12.8005
R93 VTAIL.n10 VTAIL.n9 12.8005
R94 VTAIL.n48 VTAIL.n47 12.8005
R95 VTAIL.n30 VTAIL.n29 12.8005
R96 VTAIL.n67 VTAIL.n58 12.0247
R97 VTAIL.n13 VTAIL.n4 12.0247
R98 VTAIL.n51 VTAIL.n42 12.0247
R99 VTAIL.n33 VTAIL.n24 12.0247
R100 VTAIL.n68 VTAIL.n56 11.249
R101 VTAIL.n14 VTAIL.n2 11.249
R102 VTAIL.n52 VTAIL.n40 11.249
R103 VTAIL.n34 VTAIL.n22 11.249
R104 VTAIL.n70 VTAIL.n69 9.45567
R105 VTAIL.n16 VTAIL.n15 9.45567
R106 VTAIL.n54 VTAIL.n53 9.45567
R107 VTAIL.n36 VTAIL.n35 9.45567
R108 VTAIL.n69 VTAIL.n68 9.3005
R109 VTAIL.n58 VTAIL.n57 9.3005
R110 VTAIL.n63 VTAIL.n62 9.3005
R111 VTAIL.n15 VTAIL.n14 9.3005
R112 VTAIL.n4 VTAIL.n3 9.3005
R113 VTAIL.n9 VTAIL.n8 9.3005
R114 VTAIL.n53 VTAIL.n52 9.3005
R115 VTAIL.n42 VTAIL.n41 9.3005
R116 VTAIL.n47 VTAIL.n46 9.3005
R117 VTAIL.n35 VTAIL.n34 9.3005
R118 VTAIL.n24 VTAIL.n23 9.3005
R119 VTAIL.n29 VTAIL.n28 9.3005
R120 VTAIL.n0 VTAIL.t11 6.28621
R121 VTAIL.n0 VTAIL.t8 6.28621
R122 VTAIL.n18 VTAIL.t4 6.28621
R123 VTAIL.n18 VTAIL.t3 6.28621
R124 VTAIL.n38 VTAIL.t0 6.28621
R125 VTAIL.n38 VTAIL.t5 6.28621
R126 VTAIL.n20 VTAIL.t9 6.28621
R127 VTAIL.n20 VTAIL.t7 6.28621
R128 VTAIL.n62 VTAIL.n61 4.46457
R129 VTAIL.n8 VTAIL.n7 4.46457
R130 VTAIL.n46 VTAIL.n45 4.46457
R131 VTAIL.n28 VTAIL.n27 4.46457
R132 VTAIL.n70 VTAIL.n56 2.71565
R133 VTAIL.n16 VTAIL.n2 2.71565
R134 VTAIL.n54 VTAIL.n40 2.71565
R135 VTAIL.n36 VTAIL.n22 2.71565
R136 VTAIL.n37 VTAIL.n21 2.38843
R137 VTAIL.n55 VTAIL.n39 2.38843
R138 VTAIL.n19 VTAIL.n17 2.38843
R139 VTAIL.n68 VTAIL.n67 1.93989
R140 VTAIL.n14 VTAIL.n13 1.93989
R141 VTAIL.n52 VTAIL.n51 1.93989
R142 VTAIL.n34 VTAIL.n33 1.93989
R143 VTAIL VTAIL.n71 1.73326
R144 VTAIL.n39 VTAIL.n37 1.66429
R145 VTAIL.n17 VTAIL.n1 1.66429
R146 VTAIL.n64 VTAIL.n58 1.16414
R147 VTAIL.n10 VTAIL.n4 1.16414
R148 VTAIL.n48 VTAIL.n42 1.16414
R149 VTAIL.n30 VTAIL.n24 1.16414
R150 VTAIL VTAIL.n1 0.655672
R151 VTAIL.n63 VTAIL.n60 0.388379
R152 VTAIL.n9 VTAIL.n6 0.388379
R153 VTAIL.n47 VTAIL.n44 0.388379
R154 VTAIL.n29 VTAIL.n26 0.388379
R155 VTAIL.n62 VTAIL.n57 0.155672
R156 VTAIL.n69 VTAIL.n57 0.155672
R157 VTAIL.n8 VTAIL.n3 0.155672
R158 VTAIL.n15 VTAIL.n3 0.155672
R159 VTAIL.n53 VTAIL.n41 0.155672
R160 VTAIL.n46 VTAIL.n41 0.155672
R161 VTAIL.n35 VTAIL.n23 0.155672
R162 VTAIL.n28 VTAIL.n23 0.155672
R163 VDD2.n27 VDD2.n17 289.615
R164 VDD2.n10 VDD2.n0 289.615
R165 VDD2.n28 VDD2.n27 185
R166 VDD2.n26 VDD2.n25 185
R167 VDD2.n21 VDD2.n20 185
R168 VDD2.n4 VDD2.n3 185
R169 VDD2.n9 VDD2.n8 185
R170 VDD2.n11 VDD2.n10 185
R171 VDD2.n22 VDD2.t1 148.606
R172 VDD2.n5 VDD2.t5 148.606
R173 VDD2.n27 VDD2.n26 104.615
R174 VDD2.n26 VDD2.n20 104.615
R175 VDD2.n9 VDD2.n3 104.615
R176 VDD2.n10 VDD2.n9 104.615
R177 VDD2.n16 VDD2.n15 78.8725
R178 VDD2 VDD2.n33 78.8697
R179 VDD2.t1 VDD2.n20 52.3082
R180 VDD2.t5 VDD2.n3 52.3082
R181 VDD2.n16 VDD2.n14 51.1816
R182 VDD2.n32 VDD2.n31 49.446
R183 VDD2.n32 VDD2.n16 34.1916
R184 VDD2.n22 VDD2.n21 15.5966
R185 VDD2.n5 VDD2.n4 15.5966
R186 VDD2.n25 VDD2.n24 12.8005
R187 VDD2.n8 VDD2.n7 12.8005
R188 VDD2.n28 VDD2.n19 12.0247
R189 VDD2.n11 VDD2.n2 12.0247
R190 VDD2.n29 VDD2.n17 11.249
R191 VDD2.n12 VDD2.n0 11.249
R192 VDD2.n31 VDD2.n30 9.45567
R193 VDD2.n14 VDD2.n13 9.45567
R194 VDD2.n30 VDD2.n29 9.3005
R195 VDD2.n19 VDD2.n18 9.3005
R196 VDD2.n24 VDD2.n23 9.3005
R197 VDD2.n13 VDD2.n12 9.3005
R198 VDD2.n2 VDD2.n1 9.3005
R199 VDD2.n7 VDD2.n6 9.3005
R200 VDD2.n33 VDD2.t3 6.28621
R201 VDD2.n33 VDD2.t2 6.28621
R202 VDD2.n15 VDD2.t0 6.28621
R203 VDD2.n15 VDD2.t4 6.28621
R204 VDD2.n23 VDD2.n22 4.46457
R205 VDD2.n6 VDD2.n5 4.46457
R206 VDD2.n31 VDD2.n17 2.71565
R207 VDD2.n14 VDD2.n0 2.71565
R208 VDD2.n29 VDD2.n28 1.93989
R209 VDD2.n12 VDD2.n11 1.93989
R210 VDD2 VDD2.n32 1.84964
R211 VDD2.n25 VDD2.n19 1.16414
R212 VDD2.n8 VDD2.n2 1.16414
R213 VDD2.n24 VDD2.n21 0.388379
R214 VDD2.n7 VDD2.n4 0.388379
R215 VDD2.n30 VDD2.n18 0.155672
R216 VDD2.n23 VDD2.n18 0.155672
R217 VDD2.n6 VDD2.n1 0.155672
R218 VDD2.n13 VDD2.n1 0.155672
R219 B.n541 B.n540 585
R220 B.n542 B.n541 585
R221 B.n180 B.n97 585
R222 B.n179 B.n178 585
R223 B.n177 B.n176 585
R224 B.n175 B.n174 585
R225 B.n173 B.n172 585
R226 B.n171 B.n170 585
R227 B.n169 B.n168 585
R228 B.n167 B.n166 585
R229 B.n165 B.n164 585
R230 B.n163 B.n162 585
R231 B.n161 B.n160 585
R232 B.n159 B.n158 585
R233 B.n157 B.n156 585
R234 B.n155 B.n154 585
R235 B.n153 B.n152 585
R236 B.n150 B.n149 585
R237 B.n148 B.n147 585
R238 B.n146 B.n145 585
R239 B.n144 B.n143 585
R240 B.n142 B.n141 585
R241 B.n140 B.n139 585
R242 B.n138 B.n137 585
R243 B.n136 B.n135 585
R244 B.n134 B.n133 585
R245 B.n132 B.n131 585
R246 B.n130 B.n129 585
R247 B.n128 B.n127 585
R248 B.n126 B.n125 585
R249 B.n124 B.n123 585
R250 B.n122 B.n121 585
R251 B.n120 B.n119 585
R252 B.n118 B.n117 585
R253 B.n116 B.n115 585
R254 B.n114 B.n113 585
R255 B.n112 B.n111 585
R256 B.n110 B.n109 585
R257 B.n108 B.n107 585
R258 B.n106 B.n105 585
R259 B.n104 B.n103 585
R260 B.n75 B.n74 585
R261 B.n539 B.n76 585
R262 B.n543 B.n76 585
R263 B.n538 B.n537 585
R264 B.n537 B.n72 585
R265 B.n536 B.n71 585
R266 B.n549 B.n71 585
R267 B.n535 B.n70 585
R268 B.n550 B.n70 585
R269 B.n534 B.n69 585
R270 B.n551 B.n69 585
R271 B.n533 B.n532 585
R272 B.n532 B.n65 585
R273 B.n531 B.n64 585
R274 B.n557 B.n64 585
R275 B.n530 B.n63 585
R276 B.n558 B.n63 585
R277 B.n529 B.n62 585
R278 B.n559 B.n62 585
R279 B.n528 B.n527 585
R280 B.n527 B.n58 585
R281 B.n526 B.n57 585
R282 B.n565 B.n57 585
R283 B.n525 B.n56 585
R284 B.n566 B.n56 585
R285 B.n524 B.n55 585
R286 B.n567 B.n55 585
R287 B.n523 B.n522 585
R288 B.n522 B.n51 585
R289 B.n521 B.n50 585
R290 B.n573 B.n50 585
R291 B.n520 B.n49 585
R292 B.n574 B.n49 585
R293 B.n519 B.n48 585
R294 B.n575 B.n48 585
R295 B.n518 B.n517 585
R296 B.n517 B.n44 585
R297 B.n516 B.n43 585
R298 B.n581 B.n43 585
R299 B.n515 B.n42 585
R300 B.n582 B.n42 585
R301 B.n514 B.n41 585
R302 B.n583 B.n41 585
R303 B.n513 B.n512 585
R304 B.n512 B.n37 585
R305 B.n511 B.n36 585
R306 B.n589 B.n36 585
R307 B.n510 B.n35 585
R308 B.n590 B.n35 585
R309 B.n509 B.n34 585
R310 B.n591 B.n34 585
R311 B.n508 B.n507 585
R312 B.n507 B.n30 585
R313 B.n506 B.n29 585
R314 B.n597 B.n29 585
R315 B.n505 B.n28 585
R316 B.n598 B.n28 585
R317 B.n504 B.n27 585
R318 B.n599 B.n27 585
R319 B.n503 B.n502 585
R320 B.n502 B.n23 585
R321 B.n501 B.n22 585
R322 B.n605 B.n22 585
R323 B.n500 B.n21 585
R324 B.n606 B.n21 585
R325 B.n499 B.n20 585
R326 B.n607 B.n20 585
R327 B.n498 B.n497 585
R328 B.n497 B.n16 585
R329 B.n496 B.n15 585
R330 B.n613 B.n15 585
R331 B.n495 B.n14 585
R332 B.n614 B.n14 585
R333 B.n494 B.n13 585
R334 B.n615 B.n13 585
R335 B.n493 B.n492 585
R336 B.n492 B.n12 585
R337 B.n491 B.n490 585
R338 B.n491 B.n8 585
R339 B.n489 B.n7 585
R340 B.n622 B.n7 585
R341 B.n488 B.n6 585
R342 B.n623 B.n6 585
R343 B.n487 B.n5 585
R344 B.n624 B.n5 585
R345 B.n486 B.n485 585
R346 B.n485 B.n4 585
R347 B.n484 B.n181 585
R348 B.n484 B.n483 585
R349 B.n474 B.n182 585
R350 B.n183 B.n182 585
R351 B.n476 B.n475 585
R352 B.n477 B.n476 585
R353 B.n473 B.n188 585
R354 B.n188 B.n187 585
R355 B.n472 B.n471 585
R356 B.n471 B.n470 585
R357 B.n190 B.n189 585
R358 B.n191 B.n190 585
R359 B.n463 B.n462 585
R360 B.n464 B.n463 585
R361 B.n461 B.n196 585
R362 B.n196 B.n195 585
R363 B.n460 B.n459 585
R364 B.n459 B.n458 585
R365 B.n198 B.n197 585
R366 B.n199 B.n198 585
R367 B.n451 B.n450 585
R368 B.n452 B.n451 585
R369 B.n449 B.n204 585
R370 B.n204 B.n203 585
R371 B.n448 B.n447 585
R372 B.n447 B.n446 585
R373 B.n206 B.n205 585
R374 B.n207 B.n206 585
R375 B.n439 B.n438 585
R376 B.n440 B.n439 585
R377 B.n437 B.n212 585
R378 B.n212 B.n211 585
R379 B.n436 B.n435 585
R380 B.n435 B.n434 585
R381 B.n214 B.n213 585
R382 B.n215 B.n214 585
R383 B.n427 B.n426 585
R384 B.n428 B.n427 585
R385 B.n425 B.n220 585
R386 B.n220 B.n219 585
R387 B.n424 B.n423 585
R388 B.n423 B.n422 585
R389 B.n222 B.n221 585
R390 B.n223 B.n222 585
R391 B.n415 B.n414 585
R392 B.n416 B.n415 585
R393 B.n413 B.n228 585
R394 B.n228 B.n227 585
R395 B.n412 B.n411 585
R396 B.n411 B.n410 585
R397 B.n230 B.n229 585
R398 B.n231 B.n230 585
R399 B.n403 B.n402 585
R400 B.n404 B.n403 585
R401 B.n401 B.n236 585
R402 B.n236 B.n235 585
R403 B.n400 B.n399 585
R404 B.n399 B.n398 585
R405 B.n238 B.n237 585
R406 B.n239 B.n238 585
R407 B.n391 B.n390 585
R408 B.n392 B.n391 585
R409 B.n389 B.n243 585
R410 B.n247 B.n243 585
R411 B.n388 B.n387 585
R412 B.n387 B.n386 585
R413 B.n245 B.n244 585
R414 B.n246 B.n245 585
R415 B.n379 B.n378 585
R416 B.n380 B.n379 585
R417 B.n377 B.n252 585
R418 B.n252 B.n251 585
R419 B.n376 B.n375 585
R420 B.n375 B.n374 585
R421 B.n254 B.n253 585
R422 B.n255 B.n254 585
R423 B.n367 B.n366 585
R424 B.n368 B.n367 585
R425 B.n258 B.n257 585
R426 B.n286 B.n284 585
R427 B.n287 B.n283 585
R428 B.n287 B.n259 585
R429 B.n290 B.n289 585
R430 B.n291 B.n282 585
R431 B.n293 B.n292 585
R432 B.n295 B.n281 585
R433 B.n298 B.n297 585
R434 B.n299 B.n280 585
R435 B.n301 B.n300 585
R436 B.n303 B.n279 585
R437 B.n306 B.n305 585
R438 B.n307 B.n278 585
R439 B.n309 B.n308 585
R440 B.n311 B.n277 585
R441 B.n314 B.n313 585
R442 B.n316 B.n274 585
R443 B.n318 B.n317 585
R444 B.n320 B.n273 585
R445 B.n323 B.n322 585
R446 B.n324 B.n272 585
R447 B.n326 B.n325 585
R448 B.n328 B.n271 585
R449 B.n331 B.n330 585
R450 B.n332 B.n268 585
R451 B.n335 B.n334 585
R452 B.n337 B.n267 585
R453 B.n340 B.n339 585
R454 B.n341 B.n266 585
R455 B.n343 B.n342 585
R456 B.n345 B.n265 585
R457 B.n348 B.n347 585
R458 B.n349 B.n264 585
R459 B.n351 B.n350 585
R460 B.n353 B.n263 585
R461 B.n356 B.n355 585
R462 B.n357 B.n262 585
R463 B.n359 B.n358 585
R464 B.n361 B.n261 585
R465 B.n364 B.n363 585
R466 B.n365 B.n260 585
R467 B.n370 B.n369 585
R468 B.n369 B.n368 585
R469 B.n371 B.n256 585
R470 B.n256 B.n255 585
R471 B.n373 B.n372 585
R472 B.n374 B.n373 585
R473 B.n250 B.n249 585
R474 B.n251 B.n250 585
R475 B.n382 B.n381 585
R476 B.n381 B.n380 585
R477 B.n383 B.n248 585
R478 B.n248 B.n246 585
R479 B.n385 B.n384 585
R480 B.n386 B.n385 585
R481 B.n242 B.n241 585
R482 B.n247 B.n242 585
R483 B.n394 B.n393 585
R484 B.n393 B.n392 585
R485 B.n395 B.n240 585
R486 B.n240 B.n239 585
R487 B.n397 B.n396 585
R488 B.n398 B.n397 585
R489 B.n234 B.n233 585
R490 B.n235 B.n234 585
R491 B.n406 B.n405 585
R492 B.n405 B.n404 585
R493 B.n407 B.n232 585
R494 B.n232 B.n231 585
R495 B.n409 B.n408 585
R496 B.n410 B.n409 585
R497 B.n226 B.n225 585
R498 B.n227 B.n226 585
R499 B.n418 B.n417 585
R500 B.n417 B.n416 585
R501 B.n419 B.n224 585
R502 B.n224 B.n223 585
R503 B.n421 B.n420 585
R504 B.n422 B.n421 585
R505 B.n218 B.n217 585
R506 B.n219 B.n218 585
R507 B.n430 B.n429 585
R508 B.n429 B.n428 585
R509 B.n431 B.n216 585
R510 B.n216 B.n215 585
R511 B.n433 B.n432 585
R512 B.n434 B.n433 585
R513 B.n210 B.n209 585
R514 B.n211 B.n210 585
R515 B.n442 B.n441 585
R516 B.n441 B.n440 585
R517 B.n443 B.n208 585
R518 B.n208 B.n207 585
R519 B.n445 B.n444 585
R520 B.n446 B.n445 585
R521 B.n202 B.n201 585
R522 B.n203 B.n202 585
R523 B.n454 B.n453 585
R524 B.n453 B.n452 585
R525 B.n455 B.n200 585
R526 B.n200 B.n199 585
R527 B.n457 B.n456 585
R528 B.n458 B.n457 585
R529 B.n194 B.n193 585
R530 B.n195 B.n194 585
R531 B.n466 B.n465 585
R532 B.n465 B.n464 585
R533 B.n467 B.n192 585
R534 B.n192 B.n191 585
R535 B.n469 B.n468 585
R536 B.n470 B.n469 585
R537 B.n186 B.n185 585
R538 B.n187 B.n186 585
R539 B.n479 B.n478 585
R540 B.n478 B.n477 585
R541 B.n480 B.n184 585
R542 B.n184 B.n183 585
R543 B.n482 B.n481 585
R544 B.n483 B.n482 585
R545 B.n3 B.n0 585
R546 B.n4 B.n3 585
R547 B.n621 B.n1 585
R548 B.n622 B.n621 585
R549 B.n620 B.n619 585
R550 B.n620 B.n8 585
R551 B.n618 B.n9 585
R552 B.n12 B.n9 585
R553 B.n617 B.n616 585
R554 B.n616 B.n615 585
R555 B.n11 B.n10 585
R556 B.n614 B.n11 585
R557 B.n612 B.n611 585
R558 B.n613 B.n612 585
R559 B.n610 B.n17 585
R560 B.n17 B.n16 585
R561 B.n609 B.n608 585
R562 B.n608 B.n607 585
R563 B.n19 B.n18 585
R564 B.n606 B.n19 585
R565 B.n604 B.n603 585
R566 B.n605 B.n604 585
R567 B.n602 B.n24 585
R568 B.n24 B.n23 585
R569 B.n601 B.n600 585
R570 B.n600 B.n599 585
R571 B.n26 B.n25 585
R572 B.n598 B.n26 585
R573 B.n596 B.n595 585
R574 B.n597 B.n596 585
R575 B.n594 B.n31 585
R576 B.n31 B.n30 585
R577 B.n593 B.n592 585
R578 B.n592 B.n591 585
R579 B.n33 B.n32 585
R580 B.n590 B.n33 585
R581 B.n588 B.n587 585
R582 B.n589 B.n588 585
R583 B.n586 B.n38 585
R584 B.n38 B.n37 585
R585 B.n585 B.n584 585
R586 B.n584 B.n583 585
R587 B.n40 B.n39 585
R588 B.n582 B.n40 585
R589 B.n580 B.n579 585
R590 B.n581 B.n580 585
R591 B.n578 B.n45 585
R592 B.n45 B.n44 585
R593 B.n577 B.n576 585
R594 B.n576 B.n575 585
R595 B.n47 B.n46 585
R596 B.n574 B.n47 585
R597 B.n572 B.n571 585
R598 B.n573 B.n572 585
R599 B.n570 B.n52 585
R600 B.n52 B.n51 585
R601 B.n569 B.n568 585
R602 B.n568 B.n567 585
R603 B.n54 B.n53 585
R604 B.n566 B.n54 585
R605 B.n564 B.n563 585
R606 B.n565 B.n564 585
R607 B.n562 B.n59 585
R608 B.n59 B.n58 585
R609 B.n561 B.n560 585
R610 B.n560 B.n559 585
R611 B.n61 B.n60 585
R612 B.n558 B.n61 585
R613 B.n556 B.n555 585
R614 B.n557 B.n556 585
R615 B.n554 B.n66 585
R616 B.n66 B.n65 585
R617 B.n553 B.n552 585
R618 B.n552 B.n551 585
R619 B.n68 B.n67 585
R620 B.n550 B.n68 585
R621 B.n548 B.n547 585
R622 B.n549 B.n548 585
R623 B.n546 B.n73 585
R624 B.n73 B.n72 585
R625 B.n545 B.n544 585
R626 B.n544 B.n543 585
R627 B.n625 B.n624 585
R628 B.n623 B.n2 585
R629 B.n544 B.n75 511.721
R630 B.n541 B.n76 511.721
R631 B.n367 B.n260 511.721
R632 B.n369 B.n258 511.721
R633 B.n542 B.n96 256.663
R634 B.n542 B.n95 256.663
R635 B.n542 B.n94 256.663
R636 B.n542 B.n93 256.663
R637 B.n542 B.n92 256.663
R638 B.n542 B.n91 256.663
R639 B.n542 B.n90 256.663
R640 B.n542 B.n89 256.663
R641 B.n542 B.n88 256.663
R642 B.n542 B.n87 256.663
R643 B.n542 B.n86 256.663
R644 B.n542 B.n85 256.663
R645 B.n542 B.n84 256.663
R646 B.n542 B.n83 256.663
R647 B.n542 B.n82 256.663
R648 B.n542 B.n81 256.663
R649 B.n542 B.n80 256.663
R650 B.n542 B.n79 256.663
R651 B.n542 B.n78 256.663
R652 B.n542 B.n77 256.663
R653 B.n285 B.n259 256.663
R654 B.n288 B.n259 256.663
R655 B.n294 B.n259 256.663
R656 B.n296 B.n259 256.663
R657 B.n302 B.n259 256.663
R658 B.n304 B.n259 256.663
R659 B.n310 B.n259 256.663
R660 B.n312 B.n259 256.663
R661 B.n319 B.n259 256.663
R662 B.n321 B.n259 256.663
R663 B.n327 B.n259 256.663
R664 B.n329 B.n259 256.663
R665 B.n336 B.n259 256.663
R666 B.n338 B.n259 256.663
R667 B.n344 B.n259 256.663
R668 B.n346 B.n259 256.663
R669 B.n352 B.n259 256.663
R670 B.n354 B.n259 256.663
R671 B.n360 B.n259 256.663
R672 B.n362 B.n259 256.663
R673 B.n627 B.n626 256.663
R674 B.n100 B.t14 238.905
R675 B.n98 B.t6 238.905
R676 B.n269 B.t10 238.905
R677 B.n275 B.t17 238.905
R678 B.n98 B.t8 184.93
R679 B.n269 B.t13 184.93
R680 B.n100 B.t15 184.93
R681 B.n275 B.t19 184.93
R682 B.n368 B.n259 178.873
R683 B.n543 B.n542 178.873
R684 B.n105 B.n104 163.367
R685 B.n109 B.n108 163.367
R686 B.n113 B.n112 163.367
R687 B.n117 B.n116 163.367
R688 B.n121 B.n120 163.367
R689 B.n125 B.n124 163.367
R690 B.n129 B.n128 163.367
R691 B.n133 B.n132 163.367
R692 B.n137 B.n136 163.367
R693 B.n141 B.n140 163.367
R694 B.n145 B.n144 163.367
R695 B.n149 B.n148 163.367
R696 B.n154 B.n153 163.367
R697 B.n158 B.n157 163.367
R698 B.n162 B.n161 163.367
R699 B.n166 B.n165 163.367
R700 B.n170 B.n169 163.367
R701 B.n174 B.n173 163.367
R702 B.n178 B.n177 163.367
R703 B.n541 B.n97 163.367
R704 B.n367 B.n254 163.367
R705 B.n375 B.n254 163.367
R706 B.n375 B.n252 163.367
R707 B.n379 B.n252 163.367
R708 B.n379 B.n245 163.367
R709 B.n387 B.n245 163.367
R710 B.n387 B.n243 163.367
R711 B.n391 B.n243 163.367
R712 B.n391 B.n238 163.367
R713 B.n399 B.n238 163.367
R714 B.n399 B.n236 163.367
R715 B.n403 B.n236 163.367
R716 B.n403 B.n230 163.367
R717 B.n411 B.n230 163.367
R718 B.n411 B.n228 163.367
R719 B.n415 B.n228 163.367
R720 B.n415 B.n222 163.367
R721 B.n423 B.n222 163.367
R722 B.n423 B.n220 163.367
R723 B.n427 B.n220 163.367
R724 B.n427 B.n214 163.367
R725 B.n435 B.n214 163.367
R726 B.n435 B.n212 163.367
R727 B.n439 B.n212 163.367
R728 B.n439 B.n206 163.367
R729 B.n447 B.n206 163.367
R730 B.n447 B.n204 163.367
R731 B.n451 B.n204 163.367
R732 B.n451 B.n198 163.367
R733 B.n459 B.n198 163.367
R734 B.n459 B.n196 163.367
R735 B.n463 B.n196 163.367
R736 B.n463 B.n190 163.367
R737 B.n471 B.n190 163.367
R738 B.n471 B.n188 163.367
R739 B.n476 B.n188 163.367
R740 B.n476 B.n182 163.367
R741 B.n484 B.n182 163.367
R742 B.n485 B.n484 163.367
R743 B.n485 B.n5 163.367
R744 B.n6 B.n5 163.367
R745 B.n7 B.n6 163.367
R746 B.n491 B.n7 163.367
R747 B.n492 B.n491 163.367
R748 B.n492 B.n13 163.367
R749 B.n14 B.n13 163.367
R750 B.n15 B.n14 163.367
R751 B.n497 B.n15 163.367
R752 B.n497 B.n20 163.367
R753 B.n21 B.n20 163.367
R754 B.n22 B.n21 163.367
R755 B.n502 B.n22 163.367
R756 B.n502 B.n27 163.367
R757 B.n28 B.n27 163.367
R758 B.n29 B.n28 163.367
R759 B.n507 B.n29 163.367
R760 B.n507 B.n34 163.367
R761 B.n35 B.n34 163.367
R762 B.n36 B.n35 163.367
R763 B.n512 B.n36 163.367
R764 B.n512 B.n41 163.367
R765 B.n42 B.n41 163.367
R766 B.n43 B.n42 163.367
R767 B.n517 B.n43 163.367
R768 B.n517 B.n48 163.367
R769 B.n49 B.n48 163.367
R770 B.n50 B.n49 163.367
R771 B.n522 B.n50 163.367
R772 B.n522 B.n55 163.367
R773 B.n56 B.n55 163.367
R774 B.n57 B.n56 163.367
R775 B.n527 B.n57 163.367
R776 B.n527 B.n62 163.367
R777 B.n63 B.n62 163.367
R778 B.n64 B.n63 163.367
R779 B.n532 B.n64 163.367
R780 B.n532 B.n69 163.367
R781 B.n70 B.n69 163.367
R782 B.n71 B.n70 163.367
R783 B.n537 B.n71 163.367
R784 B.n537 B.n76 163.367
R785 B.n287 B.n286 163.367
R786 B.n289 B.n287 163.367
R787 B.n293 B.n282 163.367
R788 B.n297 B.n295 163.367
R789 B.n301 B.n280 163.367
R790 B.n305 B.n303 163.367
R791 B.n309 B.n278 163.367
R792 B.n313 B.n311 163.367
R793 B.n318 B.n274 163.367
R794 B.n322 B.n320 163.367
R795 B.n326 B.n272 163.367
R796 B.n330 B.n328 163.367
R797 B.n335 B.n268 163.367
R798 B.n339 B.n337 163.367
R799 B.n343 B.n266 163.367
R800 B.n347 B.n345 163.367
R801 B.n351 B.n264 163.367
R802 B.n355 B.n353 163.367
R803 B.n359 B.n262 163.367
R804 B.n363 B.n361 163.367
R805 B.n369 B.n256 163.367
R806 B.n373 B.n256 163.367
R807 B.n373 B.n250 163.367
R808 B.n381 B.n250 163.367
R809 B.n381 B.n248 163.367
R810 B.n385 B.n248 163.367
R811 B.n385 B.n242 163.367
R812 B.n393 B.n242 163.367
R813 B.n393 B.n240 163.367
R814 B.n397 B.n240 163.367
R815 B.n397 B.n234 163.367
R816 B.n405 B.n234 163.367
R817 B.n405 B.n232 163.367
R818 B.n409 B.n232 163.367
R819 B.n409 B.n226 163.367
R820 B.n417 B.n226 163.367
R821 B.n417 B.n224 163.367
R822 B.n421 B.n224 163.367
R823 B.n421 B.n218 163.367
R824 B.n429 B.n218 163.367
R825 B.n429 B.n216 163.367
R826 B.n433 B.n216 163.367
R827 B.n433 B.n210 163.367
R828 B.n441 B.n210 163.367
R829 B.n441 B.n208 163.367
R830 B.n445 B.n208 163.367
R831 B.n445 B.n202 163.367
R832 B.n453 B.n202 163.367
R833 B.n453 B.n200 163.367
R834 B.n457 B.n200 163.367
R835 B.n457 B.n194 163.367
R836 B.n465 B.n194 163.367
R837 B.n465 B.n192 163.367
R838 B.n469 B.n192 163.367
R839 B.n469 B.n186 163.367
R840 B.n478 B.n186 163.367
R841 B.n478 B.n184 163.367
R842 B.n482 B.n184 163.367
R843 B.n482 B.n3 163.367
R844 B.n625 B.n3 163.367
R845 B.n621 B.n2 163.367
R846 B.n621 B.n620 163.367
R847 B.n620 B.n9 163.367
R848 B.n616 B.n9 163.367
R849 B.n616 B.n11 163.367
R850 B.n612 B.n11 163.367
R851 B.n612 B.n17 163.367
R852 B.n608 B.n17 163.367
R853 B.n608 B.n19 163.367
R854 B.n604 B.n19 163.367
R855 B.n604 B.n24 163.367
R856 B.n600 B.n24 163.367
R857 B.n600 B.n26 163.367
R858 B.n596 B.n26 163.367
R859 B.n596 B.n31 163.367
R860 B.n592 B.n31 163.367
R861 B.n592 B.n33 163.367
R862 B.n588 B.n33 163.367
R863 B.n588 B.n38 163.367
R864 B.n584 B.n38 163.367
R865 B.n584 B.n40 163.367
R866 B.n580 B.n40 163.367
R867 B.n580 B.n45 163.367
R868 B.n576 B.n45 163.367
R869 B.n576 B.n47 163.367
R870 B.n572 B.n47 163.367
R871 B.n572 B.n52 163.367
R872 B.n568 B.n52 163.367
R873 B.n568 B.n54 163.367
R874 B.n564 B.n54 163.367
R875 B.n564 B.n59 163.367
R876 B.n560 B.n59 163.367
R877 B.n560 B.n61 163.367
R878 B.n556 B.n61 163.367
R879 B.n556 B.n66 163.367
R880 B.n552 B.n66 163.367
R881 B.n552 B.n68 163.367
R882 B.n548 B.n68 163.367
R883 B.n548 B.n73 163.367
R884 B.n544 B.n73 163.367
R885 B.n99 B.t9 131.209
R886 B.n270 B.t12 131.209
R887 B.n101 B.t16 131.209
R888 B.n276 B.t18 131.209
R889 B.n368 B.n255 88.7839
R890 B.n374 B.n255 88.7839
R891 B.n374 B.n251 88.7839
R892 B.n380 B.n251 88.7839
R893 B.n380 B.n246 88.7839
R894 B.n386 B.n246 88.7839
R895 B.n386 B.n247 88.7839
R896 B.n392 B.n239 88.7839
R897 B.n398 B.n239 88.7839
R898 B.n398 B.n235 88.7839
R899 B.n404 B.n235 88.7839
R900 B.n404 B.n231 88.7839
R901 B.n410 B.n231 88.7839
R902 B.n410 B.n227 88.7839
R903 B.n416 B.n227 88.7839
R904 B.n416 B.n223 88.7839
R905 B.n422 B.n223 88.7839
R906 B.n428 B.n219 88.7839
R907 B.n428 B.n215 88.7839
R908 B.n434 B.n215 88.7839
R909 B.n434 B.n211 88.7839
R910 B.n440 B.n211 88.7839
R911 B.n440 B.n207 88.7839
R912 B.n446 B.n207 88.7839
R913 B.n452 B.n203 88.7839
R914 B.n452 B.n199 88.7839
R915 B.n458 B.n199 88.7839
R916 B.n458 B.n195 88.7839
R917 B.n464 B.n195 88.7839
R918 B.n464 B.n191 88.7839
R919 B.n470 B.n191 88.7839
R920 B.n477 B.n187 88.7839
R921 B.n477 B.n183 88.7839
R922 B.n483 B.n183 88.7839
R923 B.n483 B.n4 88.7839
R924 B.n624 B.n4 88.7839
R925 B.n624 B.n623 88.7839
R926 B.n623 B.n622 88.7839
R927 B.n622 B.n8 88.7839
R928 B.n12 B.n8 88.7839
R929 B.n615 B.n12 88.7839
R930 B.n615 B.n614 88.7839
R931 B.n613 B.n16 88.7839
R932 B.n607 B.n16 88.7839
R933 B.n607 B.n606 88.7839
R934 B.n606 B.n605 88.7839
R935 B.n605 B.n23 88.7839
R936 B.n599 B.n23 88.7839
R937 B.n599 B.n598 88.7839
R938 B.n597 B.n30 88.7839
R939 B.n591 B.n30 88.7839
R940 B.n591 B.n590 88.7839
R941 B.n590 B.n589 88.7839
R942 B.n589 B.n37 88.7839
R943 B.n583 B.n37 88.7839
R944 B.n583 B.n582 88.7839
R945 B.n581 B.n44 88.7839
R946 B.n575 B.n44 88.7839
R947 B.n575 B.n574 88.7839
R948 B.n574 B.n573 88.7839
R949 B.n573 B.n51 88.7839
R950 B.n567 B.n51 88.7839
R951 B.n567 B.n566 88.7839
R952 B.n566 B.n565 88.7839
R953 B.n565 B.n58 88.7839
R954 B.n559 B.n58 88.7839
R955 B.n558 B.n557 88.7839
R956 B.n557 B.n65 88.7839
R957 B.n551 B.n65 88.7839
R958 B.n551 B.n550 88.7839
R959 B.n550 B.n549 88.7839
R960 B.n549 B.n72 88.7839
R961 B.n543 B.n72 88.7839
R962 B.n392 B.t11 73.1162
R963 B.n470 B.t2 73.1162
R964 B.t0 B.n613 73.1162
R965 B.n559 B.t7 73.1162
R966 B.n77 B.n75 71.676
R967 B.n105 B.n78 71.676
R968 B.n109 B.n79 71.676
R969 B.n113 B.n80 71.676
R970 B.n117 B.n81 71.676
R971 B.n121 B.n82 71.676
R972 B.n125 B.n83 71.676
R973 B.n129 B.n84 71.676
R974 B.n133 B.n85 71.676
R975 B.n137 B.n86 71.676
R976 B.n141 B.n87 71.676
R977 B.n145 B.n88 71.676
R978 B.n149 B.n89 71.676
R979 B.n154 B.n90 71.676
R980 B.n158 B.n91 71.676
R981 B.n162 B.n92 71.676
R982 B.n166 B.n93 71.676
R983 B.n170 B.n94 71.676
R984 B.n174 B.n95 71.676
R985 B.n178 B.n96 71.676
R986 B.n97 B.n96 71.676
R987 B.n177 B.n95 71.676
R988 B.n173 B.n94 71.676
R989 B.n169 B.n93 71.676
R990 B.n165 B.n92 71.676
R991 B.n161 B.n91 71.676
R992 B.n157 B.n90 71.676
R993 B.n153 B.n89 71.676
R994 B.n148 B.n88 71.676
R995 B.n144 B.n87 71.676
R996 B.n140 B.n86 71.676
R997 B.n136 B.n85 71.676
R998 B.n132 B.n84 71.676
R999 B.n128 B.n83 71.676
R1000 B.n124 B.n82 71.676
R1001 B.n120 B.n81 71.676
R1002 B.n116 B.n80 71.676
R1003 B.n112 B.n79 71.676
R1004 B.n108 B.n78 71.676
R1005 B.n104 B.n77 71.676
R1006 B.n285 B.n258 71.676
R1007 B.n289 B.n288 71.676
R1008 B.n294 B.n293 71.676
R1009 B.n297 B.n296 71.676
R1010 B.n302 B.n301 71.676
R1011 B.n305 B.n304 71.676
R1012 B.n310 B.n309 71.676
R1013 B.n313 B.n312 71.676
R1014 B.n319 B.n318 71.676
R1015 B.n322 B.n321 71.676
R1016 B.n327 B.n326 71.676
R1017 B.n330 B.n329 71.676
R1018 B.n336 B.n335 71.676
R1019 B.n339 B.n338 71.676
R1020 B.n344 B.n343 71.676
R1021 B.n347 B.n346 71.676
R1022 B.n352 B.n351 71.676
R1023 B.n355 B.n354 71.676
R1024 B.n360 B.n359 71.676
R1025 B.n363 B.n362 71.676
R1026 B.n286 B.n285 71.676
R1027 B.n288 B.n282 71.676
R1028 B.n295 B.n294 71.676
R1029 B.n296 B.n280 71.676
R1030 B.n303 B.n302 71.676
R1031 B.n304 B.n278 71.676
R1032 B.n311 B.n310 71.676
R1033 B.n312 B.n274 71.676
R1034 B.n320 B.n319 71.676
R1035 B.n321 B.n272 71.676
R1036 B.n328 B.n327 71.676
R1037 B.n329 B.n268 71.676
R1038 B.n337 B.n336 71.676
R1039 B.n338 B.n266 71.676
R1040 B.n345 B.n344 71.676
R1041 B.n346 B.n264 71.676
R1042 B.n353 B.n352 71.676
R1043 B.n354 B.n262 71.676
R1044 B.n361 B.n360 71.676
R1045 B.n362 B.n260 71.676
R1046 B.n626 B.n625 71.676
R1047 B.n626 B.n2 71.676
R1048 B.n446 B.t3 60.0598
R1049 B.t5 B.n597 60.0598
R1050 B.n102 B.n101 59.5399
R1051 B.n151 B.n99 59.5399
R1052 B.n333 B.n270 59.5399
R1053 B.n315 B.n276 59.5399
R1054 B.n101 B.n100 53.7217
R1055 B.n99 B.n98 53.7217
R1056 B.n270 B.n269 53.7217
R1057 B.n276 B.n275 53.7217
R1058 B.n422 B.t4 47.0035
R1059 B.t1 B.n581 47.0035
R1060 B.t4 B.n219 41.7809
R1061 B.n582 B.t1 41.7809
R1062 B.n370 B.n257 33.2493
R1063 B.n366 B.n365 33.2493
R1064 B.n540 B.n539 33.2493
R1065 B.n545 B.n74 33.2493
R1066 B.t3 B.n203 28.7245
R1067 B.n598 B.t5 28.7245
R1068 B B.n627 18.0485
R1069 B.n247 B.t11 15.6682
R1070 B.t2 B.n187 15.6682
R1071 B.n614 B.t0 15.6682
R1072 B.t7 B.n558 15.6682
R1073 B.n371 B.n370 10.6151
R1074 B.n372 B.n371 10.6151
R1075 B.n372 B.n249 10.6151
R1076 B.n382 B.n249 10.6151
R1077 B.n383 B.n382 10.6151
R1078 B.n384 B.n383 10.6151
R1079 B.n384 B.n241 10.6151
R1080 B.n394 B.n241 10.6151
R1081 B.n395 B.n394 10.6151
R1082 B.n396 B.n395 10.6151
R1083 B.n396 B.n233 10.6151
R1084 B.n406 B.n233 10.6151
R1085 B.n407 B.n406 10.6151
R1086 B.n408 B.n407 10.6151
R1087 B.n408 B.n225 10.6151
R1088 B.n418 B.n225 10.6151
R1089 B.n419 B.n418 10.6151
R1090 B.n420 B.n419 10.6151
R1091 B.n420 B.n217 10.6151
R1092 B.n430 B.n217 10.6151
R1093 B.n431 B.n430 10.6151
R1094 B.n432 B.n431 10.6151
R1095 B.n432 B.n209 10.6151
R1096 B.n442 B.n209 10.6151
R1097 B.n443 B.n442 10.6151
R1098 B.n444 B.n443 10.6151
R1099 B.n444 B.n201 10.6151
R1100 B.n454 B.n201 10.6151
R1101 B.n455 B.n454 10.6151
R1102 B.n456 B.n455 10.6151
R1103 B.n456 B.n193 10.6151
R1104 B.n466 B.n193 10.6151
R1105 B.n467 B.n466 10.6151
R1106 B.n468 B.n467 10.6151
R1107 B.n468 B.n185 10.6151
R1108 B.n479 B.n185 10.6151
R1109 B.n480 B.n479 10.6151
R1110 B.n481 B.n480 10.6151
R1111 B.n481 B.n0 10.6151
R1112 B.n284 B.n257 10.6151
R1113 B.n284 B.n283 10.6151
R1114 B.n290 B.n283 10.6151
R1115 B.n291 B.n290 10.6151
R1116 B.n292 B.n291 10.6151
R1117 B.n292 B.n281 10.6151
R1118 B.n298 B.n281 10.6151
R1119 B.n299 B.n298 10.6151
R1120 B.n300 B.n299 10.6151
R1121 B.n300 B.n279 10.6151
R1122 B.n306 B.n279 10.6151
R1123 B.n307 B.n306 10.6151
R1124 B.n308 B.n307 10.6151
R1125 B.n308 B.n277 10.6151
R1126 B.n314 B.n277 10.6151
R1127 B.n317 B.n316 10.6151
R1128 B.n317 B.n273 10.6151
R1129 B.n323 B.n273 10.6151
R1130 B.n324 B.n323 10.6151
R1131 B.n325 B.n324 10.6151
R1132 B.n325 B.n271 10.6151
R1133 B.n331 B.n271 10.6151
R1134 B.n332 B.n331 10.6151
R1135 B.n334 B.n267 10.6151
R1136 B.n340 B.n267 10.6151
R1137 B.n341 B.n340 10.6151
R1138 B.n342 B.n341 10.6151
R1139 B.n342 B.n265 10.6151
R1140 B.n348 B.n265 10.6151
R1141 B.n349 B.n348 10.6151
R1142 B.n350 B.n349 10.6151
R1143 B.n350 B.n263 10.6151
R1144 B.n356 B.n263 10.6151
R1145 B.n357 B.n356 10.6151
R1146 B.n358 B.n357 10.6151
R1147 B.n358 B.n261 10.6151
R1148 B.n364 B.n261 10.6151
R1149 B.n365 B.n364 10.6151
R1150 B.n366 B.n253 10.6151
R1151 B.n376 B.n253 10.6151
R1152 B.n377 B.n376 10.6151
R1153 B.n378 B.n377 10.6151
R1154 B.n378 B.n244 10.6151
R1155 B.n388 B.n244 10.6151
R1156 B.n389 B.n388 10.6151
R1157 B.n390 B.n389 10.6151
R1158 B.n390 B.n237 10.6151
R1159 B.n400 B.n237 10.6151
R1160 B.n401 B.n400 10.6151
R1161 B.n402 B.n401 10.6151
R1162 B.n402 B.n229 10.6151
R1163 B.n412 B.n229 10.6151
R1164 B.n413 B.n412 10.6151
R1165 B.n414 B.n413 10.6151
R1166 B.n414 B.n221 10.6151
R1167 B.n424 B.n221 10.6151
R1168 B.n425 B.n424 10.6151
R1169 B.n426 B.n425 10.6151
R1170 B.n426 B.n213 10.6151
R1171 B.n436 B.n213 10.6151
R1172 B.n437 B.n436 10.6151
R1173 B.n438 B.n437 10.6151
R1174 B.n438 B.n205 10.6151
R1175 B.n448 B.n205 10.6151
R1176 B.n449 B.n448 10.6151
R1177 B.n450 B.n449 10.6151
R1178 B.n450 B.n197 10.6151
R1179 B.n460 B.n197 10.6151
R1180 B.n461 B.n460 10.6151
R1181 B.n462 B.n461 10.6151
R1182 B.n462 B.n189 10.6151
R1183 B.n472 B.n189 10.6151
R1184 B.n473 B.n472 10.6151
R1185 B.n475 B.n473 10.6151
R1186 B.n475 B.n474 10.6151
R1187 B.n474 B.n181 10.6151
R1188 B.n486 B.n181 10.6151
R1189 B.n487 B.n486 10.6151
R1190 B.n488 B.n487 10.6151
R1191 B.n489 B.n488 10.6151
R1192 B.n490 B.n489 10.6151
R1193 B.n493 B.n490 10.6151
R1194 B.n494 B.n493 10.6151
R1195 B.n495 B.n494 10.6151
R1196 B.n496 B.n495 10.6151
R1197 B.n498 B.n496 10.6151
R1198 B.n499 B.n498 10.6151
R1199 B.n500 B.n499 10.6151
R1200 B.n501 B.n500 10.6151
R1201 B.n503 B.n501 10.6151
R1202 B.n504 B.n503 10.6151
R1203 B.n505 B.n504 10.6151
R1204 B.n506 B.n505 10.6151
R1205 B.n508 B.n506 10.6151
R1206 B.n509 B.n508 10.6151
R1207 B.n510 B.n509 10.6151
R1208 B.n511 B.n510 10.6151
R1209 B.n513 B.n511 10.6151
R1210 B.n514 B.n513 10.6151
R1211 B.n515 B.n514 10.6151
R1212 B.n516 B.n515 10.6151
R1213 B.n518 B.n516 10.6151
R1214 B.n519 B.n518 10.6151
R1215 B.n520 B.n519 10.6151
R1216 B.n521 B.n520 10.6151
R1217 B.n523 B.n521 10.6151
R1218 B.n524 B.n523 10.6151
R1219 B.n525 B.n524 10.6151
R1220 B.n526 B.n525 10.6151
R1221 B.n528 B.n526 10.6151
R1222 B.n529 B.n528 10.6151
R1223 B.n530 B.n529 10.6151
R1224 B.n531 B.n530 10.6151
R1225 B.n533 B.n531 10.6151
R1226 B.n534 B.n533 10.6151
R1227 B.n535 B.n534 10.6151
R1228 B.n536 B.n535 10.6151
R1229 B.n538 B.n536 10.6151
R1230 B.n539 B.n538 10.6151
R1231 B.n619 B.n1 10.6151
R1232 B.n619 B.n618 10.6151
R1233 B.n618 B.n617 10.6151
R1234 B.n617 B.n10 10.6151
R1235 B.n611 B.n10 10.6151
R1236 B.n611 B.n610 10.6151
R1237 B.n610 B.n609 10.6151
R1238 B.n609 B.n18 10.6151
R1239 B.n603 B.n18 10.6151
R1240 B.n603 B.n602 10.6151
R1241 B.n602 B.n601 10.6151
R1242 B.n601 B.n25 10.6151
R1243 B.n595 B.n25 10.6151
R1244 B.n595 B.n594 10.6151
R1245 B.n594 B.n593 10.6151
R1246 B.n593 B.n32 10.6151
R1247 B.n587 B.n32 10.6151
R1248 B.n587 B.n586 10.6151
R1249 B.n586 B.n585 10.6151
R1250 B.n585 B.n39 10.6151
R1251 B.n579 B.n39 10.6151
R1252 B.n579 B.n578 10.6151
R1253 B.n578 B.n577 10.6151
R1254 B.n577 B.n46 10.6151
R1255 B.n571 B.n46 10.6151
R1256 B.n571 B.n570 10.6151
R1257 B.n570 B.n569 10.6151
R1258 B.n569 B.n53 10.6151
R1259 B.n563 B.n53 10.6151
R1260 B.n563 B.n562 10.6151
R1261 B.n562 B.n561 10.6151
R1262 B.n561 B.n60 10.6151
R1263 B.n555 B.n60 10.6151
R1264 B.n555 B.n554 10.6151
R1265 B.n554 B.n553 10.6151
R1266 B.n553 B.n67 10.6151
R1267 B.n547 B.n67 10.6151
R1268 B.n547 B.n546 10.6151
R1269 B.n546 B.n545 10.6151
R1270 B.n103 B.n74 10.6151
R1271 B.n106 B.n103 10.6151
R1272 B.n107 B.n106 10.6151
R1273 B.n110 B.n107 10.6151
R1274 B.n111 B.n110 10.6151
R1275 B.n114 B.n111 10.6151
R1276 B.n115 B.n114 10.6151
R1277 B.n118 B.n115 10.6151
R1278 B.n119 B.n118 10.6151
R1279 B.n122 B.n119 10.6151
R1280 B.n123 B.n122 10.6151
R1281 B.n126 B.n123 10.6151
R1282 B.n127 B.n126 10.6151
R1283 B.n130 B.n127 10.6151
R1284 B.n131 B.n130 10.6151
R1285 B.n135 B.n134 10.6151
R1286 B.n138 B.n135 10.6151
R1287 B.n139 B.n138 10.6151
R1288 B.n142 B.n139 10.6151
R1289 B.n143 B.n142 10.6151
R1290 B.n146 B.n143 10.6151
R1291 B.n147 B.n146 10.6151
R1292 B.n150 B.n147 10.6151
R1293 B.n155 B.n152 10.6151
R1294 B.n156 B.n155 10.6151
R1295 B.n159 B.n156 10.6151
R1296 B.n160 B.n159 10.6151
R1297 B.n163 B.n160 10.6151
R1298 B.n164 B.n163 10.6151
R1299 B.n167 B.n164 10.6151
R1300 B.n168 B.n167 10.6151
R1301 B.n171 B.n168 10.6151
R1302 B.n172 B.n171 10.6151
R1303 B.n175 B.n172 10.6151
R1304 B.n176 B.n175 10.6151
R1305 B.n179 B.n176 10.6151
R1306 B.n180 B.n179 10.6151
R1307 B.n540 B.n180 10.6151
R1308 B.n627 B.n0 8.11757
R1309 B.n627 B.n1 8.11757
R1310 B.n316 B.n315 6.5566
R1311 B.n333 B.n332 6.5566
R1312 B.n134 B.n102 6.5566
R1313 B.n151 B.n150 6.5566
R1314 B.n315 B.n314 4.05904
R1315 B.n334 B.n333 4.05904
R1316 B.n131 B.n102 4.05904
R1317 B.n152 B.n151 4.05904
R1318 VP.n11 VP.n8 161.3
R1319 VP.n13 VP.n12 161.3
R1320 VP.n14 VP.n7 161.3
R1321 VP.n16 VP.n15 161.3
R1322 VP.n17 VP.n6 161.3
R1323 VP.n37 VP.n0 161.3
R1324 VP.n36 VP.n35 161.3
R1325 VP.n34 VP.n1 161.3
R1326 VP.n33 VP.n32 161.3
R1327 VP.n31 VP.n2 161.3
R1328 VP.n30 VP.n29 161.3
R1329 VP.n28 VP.n3 161.3
R1330 VP.n27 VP.n26 161.3
R1331 VP.n25 VP.n4 161.3
R1332 VP.n24 VP.n23 161.3
R1333 VP.n22 VP.n5 161.3
R1334 VP.n21 VP.n20 97.5443
R1335 VP.n39 VP.n38 97.5443
R1336 VP.n19 VP.n18 97.5443
R1337 VP.n9 VP.t4 65.7772
R1338 VP.n26 VP.n25 51.663
R1339 VP.n32 VP.n1 51.663
R1340 VP.n12 VP.n7 51.663
R1341 VP.n10 VP.n9 48.034
R1342 VP.n21 VP.n19 41.3746
R1343 VP.n30 VP.t1 31.1132
R1344 VP.n20 VP.t2 31.1132
R1345 VP.n38 VP.t0 31.1132
R1346 VP.n10 VP.t3 31.1132
R1347 VP.n18 VP.t5 31.1132
R1348 VP.n25 VP.n24 29.3238
R1349 VP.n36 VP.n1 29.3238
R1350 VP.n16 VP.n7 29.3238
R1351 VP.n24 VP.n5 24.4675
R1352 VP.n26 VP.n3 24.4675
R1353 VP.n30 VP.n3 24.4675
R1354 VP.n31 VP.n30 24.4675
R1355 VP.n32 VP.n31 24.4675
R1356 VP.n37 VP.n36 24.4675
R1357 VP.n17 VP.n16 24.4675
R1358 VP.n11 VP.n10 24.4675
R1359 VP.n12 VP.n11 24.4675
R1360 VP.n20 VP.n5 13.2127
R1361 VP.n38 VP.n37 13.2127
R1362 VP.n18 VP.n17 13.2127
R1363 VP.n9 VP.n8 6.62503
R1364 VP.n19 VP.n6 0.278367
R1365 VP.n22 VP.n21 0.278367
R1366 VP.n39 VP.n0 0.278367
R1367 VP.n13 VP.n8 0.189894
R1368 VP.n14 VP.n13 0.189894
R1369 VP.n15 VP.n14 0.189894
R1370 VP.n15 VP.n6 0.189894
R1371 VP.n23 VP.n22 0.189894
R1372 VP.n23 VP.n4 0.189894
R1373 VP.n27 VP.n4 0.189894
R1374 VP.n28 VP.n27 0.189894
R1375 VP.n29 VP.n28 0.189894
R1376 VP.n29 VP.n2 0.189894
R1377 VP.n33 VP.n2 0.189894
R1378 VP.n34 VP.n33 0.189894
R1379 VP.n35 VP.n34 0.189894
R1380 VP.n35 VP.n0 0.189894
R1381 VP VP.n39 0.153454
R1382 VDD1.n10 VDD1.n0 289.615
R1383 VDD1.n25 VDD1.n15 289.615
R1384 VDD1.n11 VDD1.n10 185
R1385 VDD1.n9 VDD1.n8 185
R1386 VDD1.n4 VDD1.n3 185
R1387 VDD1.n19 VDD1.n18 185
R1388 VDD1.n24 VDD1.n23 185
R1389 VDD1.n26 VDD1.n25 185
R1390 VDD1.n5 VDD1.t1 148.606
R1391 VDD1.n20 VDD1.t3 148.606
R1392 VDD1.n10 VDD1.n9 104.615
R1393 VDD1.n9 VDD1.n3 104.615
R1394 VDD1.n24 VDD1.n18 104.615
R1395 VDD1.n25 VDD1.n24 104.615
R1396 VDD1.n31 VDD1.n30 78.8725
R1397 VDD1.n33 VDD1.n32 78.3309
R1398 VDD1.t1 VDD1.n3 52.3082
R1399 VDD1.t3 VDD1.n18 52.3082
R1400 VDD1 VDD1.n14 51.2951
R1401 VDD1.n31 VDD1.n29 51.1816
R1402 VDD1.n33 VDD1.n31 35.9686
R1403 VDD1.n5 VDD1.n4 15.5966
R1404 VDD1.n20 VDD1.n19 15.5966
R1405 VDD1.n8 VDD1.n7 12.8005
R1406 VDD1.n23 VDD1.n22 12.8005
R1407 VDD1.n11 VDD1.n2 12.0247
R1408 VDD1.n26 VDD1.n17 12.0247
R1409 VDD1.n12 VDD1.n0 11.249
R1410 VDD1.n27 VDD1.n15 11.249
R1411 VDD1.n14 VDD1.n13 9.45567
R1412 VDD1.n29 VDD1.n28 9.45567
R1413 VDD1.n13 VDD1.n12 9.3005
R1414 VDD1.n2 VDD1.n1 9.3005
R1415 VDD1.n7 VDD1.n6 9.3005
R1416 VDD1.n28 VDD1.n27 9.3005
R1417 VDD1.n17 VDD1.n16 9.3005
R1418 VDD1.n22 VDD1.n21 9.3005
R1419 VDD1.n32 VDD1.t2 6.28621
R1420 VDD1.n32 VDD1.t0 6.28621
R1421 VDD1.n30 VDD1.t4 6.28621
R1422 VDD1.n30 VDD1.t5 6.28621
R1423 VDD1.n6 VDD1.n5 4.46457
R1424 VDD1.n21 VDD1.n20 4.46457
R1425 VDD1.n14 VDD1.n0 2.71565
R1426 VDD1.n29 VDD1.n15 2.71565
R1427 VDD1.n12 VDD1.n11 1.93989
R1428 VDD1.n27 VDD1.n26 1.93989
R1429 VDD1.n8 VDD1.n2 1.16414
R1430 VDD1.n23 VDD1.n17 1.16414
R1431 VDD1 VDD1.n33 0.539293
R1432 VDD1.n7 VDD1.n4 0.388379
R1433 VDD1.n22 VDD1.n19 0.388379
R1434 VDD1.n13 VDD1.n1 0.155672
R1435 VDD1.n6 VDD1.n1 0.155672
R1436 VDD1.n21 VDD1.n16 0.155672
R1437 VDD1.n28 VDD1.n16 0.155672
C0 VDD2 VP 0.449655f
C1 VN VP 5.13781f
C2 VDD1 VP 2.31886f
C3 VDD2 VN 2.02708f
C4 VDD2 VDD1 1.34346f
C5 VDD1 VN 0.155494f
C6 VTAIL VP 2.73851f
C7 VDD2 VTAIL 4.47049f
C8 VTAIL VN 2.72436f
C9 VDD1 VTAIL 4.41872f
C10 VDD2 B 4.280426f
C11 VDD1 B 4.407257f
C12 VTAIL B 3.843351f
C13 VN B 11.60429f
C14 VP B 10.22261f
C15 VDD1.n0 B 0.029961f
C16 VDD1.n1 B 0.022734f
C17 VDD1.n2 B 0.012217f
C18 VDD1.n3 B 0.021657f
C19 VDD1.n4 B 0.016838f
C20 VDD1.t1 B 0.048414f
C21 VDD1.n5 B 0.083252f
C22 VDD1.n6 B 0.240432f
C23 VDD1.n7 B 0.012217f
C24 VDD1.n8 B 0.012935f
C25 VDD1.n9 B 0.028875f
C26 VDD1.n10 B 0.058984f
C27 VDD1.n11 B 0.012935f
C28 VDD1.n12 B 0.012217f
C29 VDD1.n13 B 0.053481f
C30 VDD1.n14 B 0.054841f
C31 VDD1.n15 B 0.029961f
C32 VDD1.n16 B 0.022734f
C33 VDD1.n17 B 0.012217f
C34 VDD1.n18 B 0.021657f
C35 VDD1.n19 B 0.016838f
C36 VDD1.t3 B 0.048414f
C37 VDD1.n20 B 0.083252f
C38 VDD1.n21 B 0.240432f
C39 VDD1.n22 B 0.012217f
C40 VDD1.n23 B 0.012935f
C41 VDD1.n24 B 0.028875f
C42 VDD1.n25 B 0.058984f
C43 VDD1.n26 B 0.012935f
C44 VDD1.n27 B 0.012217f
C45 VDD1.n28 B 0.053481f
C46 VDD1.n29 B 0.054185f
C47 VDD1.t4 B 0.056591f
C48 VDD1.t5 B 0.056591f
C49 VDD1.n30 B 0.427929f
C50 VDD1.n31 B 1.97742f
C51 VDD1.t2 B 0.056591f
C52 VDD1.t0 B 0.056591f
C53 VDD1.n32 B 0.425211f
C54 VDD1.n33 B 1.85153f
C55 VP.n0 B 0.041078f
C56 VP.t0 B 0.600106f
C57 VP.n1 B 0.030917f
C58 VP.n2 B 0.031157f
C59 VP.t1 B 0.600106f
C60 VP.n3 B 0.05807f
C61 VP.n4 B 0.031157f
C62 VP.n5 B 0.044882f
C63 VP.n6 B 0.041078f
C64 VP.t5 B 0.600106f
C65 VP.n7 B 0.030917f
C66 VP.n8 B 0.296096f
C67 VP.t3 B 0.600106f
C68 VP.t4 B 0.83215f
C69 VP.n9 B 0.320012f
C70 VP.n10 B 0.355818f
C71 VP.n11 B 0.05807f
C72 VP.n12 B 0.056259f
C73 VP.n13 B 0.031157f
C74 VP.n14 B 0.031157f
C75 VP.n15 B 0.031157f
C76 VP.n16 B 0.061868f
C77 VP.n17 B 0.044882f
C78 VP.n18 B 0.355796f
C79 VP.n19 B 1.28984f
C80 VP.t2 B 0.600106f
C81 VP.n20 B 0.355796f
C82 VP.n21 B 1.31691f
C83 VP.n22 B 0.041078f
C84 VP.n23 B 0.031157f
C85 VP.n24 B 0.061868f
C86 VP.n25 B 0.030917f
C87 VP.n26 B 0.056259f
C88 VP.n27 B 0.031157f
C89 VP.n28 B 0.031157f
C90 VP.n29 B 0.031157f
C91 VP.n30 B 0.281778f
C92 VP.n31 B 0.05807f
C93 VP.n32 B 0.056259f
C94 VP.n33 B 0.031157f
C95 VP.n34 B 0.031157f
C96 VP.n35 B 0.031157f
C97 VP.n36 B 0.061868f
C98 VP.n37 B 0.044882f
C99 VP.n38 B 0.355796f
C100 VP.n39 B 0.046567f
C101 VDD2.n0 B 0.029436f
C102 VDD2.n1 B 0.022336f
C103 VDD2.n2 B 0.012002f
C104 VDD2.n3 B 0.021277f
C105 VDD2.n4 B 0.016542f
C106 VDD2.t5 B 0.047565f
C107 VDD2.n5 B 0.081792f
C108 VDD2.n6 B 0.236215f
C109 VDD2.n7 B 0.012002f
C110 VDD2.n8 B 0.012708f
C111 VDD2.n9 B 0.028369f
C112 VDD2.n10 B 0.05795f
C113 VDD2.n11 B 0.012708f
C114 VDD2.n12 B 0.012002f
C115 VDD2.n13 B 0.052543f
C116 VDD2.n14 B 0.053234f
C117 VDD2.t0 B 0.055599f
C118 VDD2.t4 B 0.055599f
C119 VDD2.n15 B 0.420424f
C120 VDD2.n16 B 1.84341f
C121 VDD2.n17 B 0.029436f
C122 VDD2.n18 B 0.022336f
C123 VDD2.n19 B 0.012002f
C124 VDD2.n20 B 0.021277f
C125 VDD2.n21 B 0.016542f
C126 VDD2.t1 B 0.047565f
C127 VDD2.n22 B 0.081792f
C128 VDD2.n23 B 0.236215f
C129 VDD2.n24 B 0.012002f
C130 VDD2.n25 B 0.012708f
C131 VDD2.n26 B 0.028369f
C132 VDD2.n27 B 0.05795f
C133 VDD2.n28 B 0.012708f
C134 VDD2.n29 B 0.012002f
C135 VDD2.n30 B 0.052543f
C136 VDD2.n31 B 0.047512f
C137 VDD2.n32 B 1.62477f
C138 VDD2.t3 B 0.055599f
C139 VDD2.t2 B 0.055599f
C140 VDD2.n33 B 0.420403f
C141 VTAIL.t11 B 0.076627f
C142 VTAIL.t8 B 0.076627f
C143 VTAIL.n0 B 0.51466f
C144 VTAIL.n1 B 0.480964f
C145 VTAIL.n2 B 0.040569f
C146 VTAIL.n3 B 0.030783f
C147 VTAIL.n4 B 0.016542f
C148 VTAIL.n5 B 0.029324f
C149 VTAIL.n6 B 0.022799f
C150 VTAIL.t2 B 0.065554f
C151 VTAIL.n7 B 0.112726f
C152 VTAIL.n8 B 0.325555f
C153 VTAIL.n9 B 0.016542f
C154 VTAIL.n10 B 0.017515f
C155 VTAIL.n11 B 0.039098f
C156 VTAIL.n12 B 0.079867f
C157 VTAIL.n13 B 0.017515f
C158 VTAIL.n14 B 0.016542f
C159 VTAIL.n15 B 0.072416f
C160 VTAIL.n16 B 0.044236f
C161 VTAIL.n17 B 0.428898f
C162 VTAIL.t4 B 0.076627f
C163 VTAIL.t3 B 0.076627f
C164 VTAIL.n18 B 0.51466f
C165 VTAIL.n19 B 1.64904f
C166 VTAIL.t9 B 0.076627f
C167 VTAIL.t7 B 0.076627f
C168 VTAIL.n20 B 0.514663f
C169 VTAIL.n21 B 1.64903f
C170 VTAIL.n22 B 0.040569f
C171 VTAIL.n23 B 0.030783f
C172 VTAIL.n24 B 0.016542f
C173 VTAIL.n25 B 0.029324f
C174 VTAIL.n26 B 0.022799f
C175 VTAIL.t10 B 0.065554f
C176 VTAIL.n27 B 0.112726f
C177 VTAIL.n28 B 0.325555f
C178 VTAIL.n29 B 0.016542f
C179 VTAIL.n30 B 0.017515f
C180 VTAIL.n31 B 0.039098f
C181 VTAIL.n32 B 0.079867f
C182 VTAIL.n33 B 0.017515f
C183 VTAIL.n34 B 0.016542f
C184 VTAIL.n35 B 0.072416f
C185 VTAIL.n36 B 0.044236f
C186 VTAIL.n37 B 0.428898f
C187 VTAIL.t0 B 0.076627f
C188 VTAIL.t5 B 0.076627f
C189 VTAIL.n38 B 0.514663f
C190 VTAIL.n39 B 0.652834f
C191 VTAIL.n40 B 0.040569f
C192 VTAIL.n41 B 0.030783f
C193 VTAIL.n42 B 0.016542f
C194 VTAIL.n43 B 0.029324f
C195 VTAIL.n44 B 0.022799f
C196 VTAIL.t1 B 0.065554f
C197 VTAIL.n45 B 0.112726f
C198 VTAIL.n46 B 0.325555f
C199 VTAIL.n47 B 0.016542f
C200 VTAIL.n48 B 0.017515f
C201 VTAIL.n49 B 0.039098f
C202 VTAIL.n50 B 0.079867f
C203 VTAIL.n51 B 0.017515f
C204 VTAIL.n52 B 0.016542f
C205 VTAIL.n53 B 0.072416f
C206 VTAIL.n54 B 0.044236f
C207 VTAIL.n55 B 1.18824f
C208 VTAIL.n56 B 0.040569f
C209 VTAIL.n57 B 0.030783f
C210 VTAIL.n58 B 0.016542f
C211 VTAIL.n59 B 0.029324f
C212 VTAIL.n60 B 0.022799f
C213 VTAIL.t6 B 0.065554f
C214 VTAIL.n61 B 0.112726f
C215 VTAIL.n62 B 0.325555f
C216 VTAIL.n63 B 0.016542f
C217 VTAIL.n64 B 0.017515f
C218 VTAIL.n65 B 0.039098f
C219 VTAIL.n66 B 0.079867f
C220 VTAIL.n67 B 0.017515f
C221 VTAIL.n68 B 0.016542f
C222 VTAIL.n69 B 0.072416f
C223 VTAIL.n70 B 0.044236f
C224 VTAIL.n71 B 1.12325f
C225 VN.n0 B 0.039686f
C226 VN.t1 B 0.579767f
C227 VN.n1 B 0.029869f
C228 VN.n2 B 0.28606f
C229 VN.t5 B 0.579767f
C230 VN.t0 B 0.803946f
C231 VN.n3 B 0.309166f
C232 VN.n4 B 0.343758f
C233 VN.n5 B 0.056102f
C234 VN.n6 B 0.054352f
C235 VN.n7 B 0.030101f
C236 VN.n8 B 0.030101f
C237 VN.n9 B 0.030101f
C238 VN.n10 B 0.059771f
C239 VN.n11 B 0.043361f
C240 VN.n12 B 0.343737f
C241 VN.n13 B 0.044989f
C242 VN.n14 B 0.039686f
C243 VN.t4 B 0.579767f
C244 VN.n15 B 0.029869f
C245 VN.n16 B 0.28606f
C246 VN.t2 B 0.579767f
C247 VN.t3 B 0.803946f
C248 VN.n17 B 0.309166f
C249 VN.n18 B 0.343758f
C250 VN.n19 B 0.056102f
C251 VN.n20 B 0.054352f
C252 VN.n21 B 0.030101f
C253 VN.n22 B 0.030101f
C254 VN.n23 B 0.030101f
C255 VN.n24 B 0.059771f
C256 VN.n25 B 0.043361f
C257 VN.n26 B 0.343737f
C258 VN.n27 B 1.26283f
.ends

