* NGSPICE file created from diff_pair_sample_0243.ext - technology: sky130A

.subckt diff_pair_sample_0243 VTAIL VN VP B VDD2 VDD1
X0 B.t15 B.t13 B.t14 B.t10 sky130_fd_pr__nfet_01v8 ad=2.7027 pd=14.64 as=0 ps=0 w=6.93 l=2.91
X1 B.t12 B.t9 B.t11 B.t10 sky130_fd_pr__nfet_01v8 ad=2.7027 pd=14.64 as=0 ps=0 w=6.93 l=2.91
X2 B.t8 B.t6 B.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=2.7027 pd=14.64 as=0 ps=0 w=6.93 l=2.91
X3 VDD2.t1 VN.t0 VTAIL.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=2.7027 pd=14.64 as=2.7027 ps=14.64 w=6.93 l=2.91
X4 VDD1.t1 VP.t0 VTAIL.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=2.7027 pd=14.64 as=2.7027 ps=14.64 w=6.93 l=2.91
X5 VDD2.t0 VN.t1 VTAIL.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=2.7027 pd=14.64 as=2.7027 ps=14.64 w=6.93 l=2.91
X6 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=2.7027 pd=14.64 as=0 ps=0 w=6.93 l=2.91
X7 VDD1.t0 VP.t1 VTAIL.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=2.7027 pd=14.64 as=2.7027 ps=14.64 w=6.93 l=2.91
R0 B.n542 B.n541 585
R1 B.n543 B.n542 585
R2 B.n210 B.n84 585
R3 B.n209 B.n208 585
R4 B.n207 B.n206 585
R5 B.n205 B.n204 585
R6 B.n203 B.n202 585
R7 B.n201 B.n200 585
R8 B.n199 B.n198 585
R9 B.n197 B.n196 585
R10 B.n195 B.n194 585
R11 B.n193 B.n192 585
R12 B.n191 B.n190 585
R13 B.n189 B.n188 585
R14 B.n187 B.n186 585
R15 B.n185 B.n184 585
R16 B.n183 B.n182 585
R17 B.n181 B.n180 585
R18 B.n179 B.n178 585
R19 B.n177 B.n176 585
R20 B.n175 B.n174 585
R21 B.n173 B.n172 585
R22 B.n171 B.n170 585
R23 B.n169 B.n168 585
R24 B.n167 B.n166 585
R25 B.n165 B.n164 585
R26 B.n163 B.n162 585
R27 B.n161 B.n160 585
R28 B.n159 B.n158 585
R29 B.n157 B.n156 585
R30 B.n155 B.n154 585
R31 B.n153 B.n152 585
R32 B.n151 B.n150 585
R33 B.n149 B.n148 585
R34 B.n147 B.n146 585
R35 B.n145 B.n144 585
R36 B.n143 B.n142 585
R37 B.n140 B.n139 585
R38 B.n138 B.n137 585
R39 B.n136 B.n135 585
R40 B.n134 B.n133 585
R41 B.n132 B.n131 585
R42 B.n130 B.n129 585
R43 B.n128 B.n127 585
R44 B.n126 B.n125 585
R45 B.n124 B.n123 585
R46 B.n122 B.n121 585
R47 B.n120 B.n119 585
R48 B.n118 B.n117 585
R49 B.n116 B.n115 585
R50 B.n114 B.n113 585
R51 B.n112 B.n111 585
R52 B.n110 B.n109 585
R53 B.n108 B.n107 585
R54 B.n106 B.n105 585
R55 B.n104 B.n103 585
R56 B.n102 B.n101 585
R57 B.n100 B.n99 585
R58 B.n98 B.n97 585
R59 B.n96 B.n95 585
R60 B.n94 B.n93 585
R61 B.n92 B.n91 585
R62 B.n53 B.n52 585
R63 B.n546 B.n545 585
R64 B.n540 B.n85 585
R65 B.n85 B.n50 585
R66 B.n539 B.n49 585
R67 B.n550 B.n49 585
R68 B.n538 B.n48 585
R69 B.n551 B.n48 585
R70 B.n537 B.n47 585
R71 B.n552 B.n47 585
R72 B.n536 B.n535 585
R73 B.n535 B.n43 585
R74 B.n534 B.n42 585
R75 B.n558 B.n42 585
R76 B.n533 B.n41 585
R77 B.n559 B.n41 585
R78 B.n532 B.n40 585
R79 B.n560 B.n40 585
R80 B.n531 B.n530 585
R81 B.n530 B.n36 585
R82 B.n529 B.n35 585
R83 B.n566 B.n35 585
R84 B.n528 B.n34 585
R85 B.n567 B.n34 585
R86 B.n527 B.n33 585
R87 B.n568 B.n33 585
R88 B.n526 B.n525 585
R89 B.n525 B.n29 585
R90 B.n524 B.n28 585
R91 B.n574 B.n28 585
R92 B.n523 B.n27 585
R93 B.n575 B.n27 585
R94 B.n522 B.n26 585
R95 B.n576 B.n26 585
R96 B.n521 B.n520 585
R97 B.n520 B.n22 585
R98 B.n519 B.n21 585
R99 B.n582 B.n21 585
R100 B.n518 B.n20 585
R101 B.n583 B.n20 585
R102 B.n517 B.n19 585
R103 B.n584 B.n19 585
R104 B.n516 B.n515 585
R105 B.n515 B.n18 585
R106 B.n514 B.n14 585
R107 B.n590 B.n14 585
R108 B.n513 B.n13 585
R109 B.n591 B.n13 585
R110 B.n512 B.n12 585
R111 B.n592 B.n12 585
R112 B.n511 B.n510 585
R113 B.n510 B.n8 585
R114 B.n509 B.n7 585
R115 B.n598 B.n7 585
R116 B.n508 B.n6 585
R117 B.n599 B.n6 585
R118 B.n507 B.n5 585
R119 B.n600 B.n5 585
R120 B.n506 B.n505 585
R121 B.n505 B.n4 585
R122 B.n504 B.n211 585
R123 B.n504 B.n503 585
R124 B.n494 B.n212 585
R125 B.n213 B.n212 585
R126 B.n496 B.n495 585
R127 B.n497 B.n496 585
R128 B.n493 B.n218 585
R129 B.n218 B.n217 585
R130 B.n492 B.n491 585
R131 B.n491 B.n490 585
R132 B.n220 B.n219 585
R133 B.n483 B.n220 585
R134 B.n482 B.n481 585
R135 B.n484 B.n482 585
R136 B.n480 B.n225 585
R137 B.n225 B.n224 585
R138 B.n479 B.n478 585
R139 B.n478 B.n477 585
R140 B.n227 B.n226 585
R141 B.n228 B.n227 585
R142 B.n470 B.n469 585
R143 B.n471 B.n470 585
R144 B.n468 B.n233 585
R145 B.n233 B.n232 585
R146 B.n467 B.n466 585
R147 B.n466 B.n465 585
R148 B.n235 B.n234 585
R149 B.n236 B.n235 585
R150 B.n458 B.n457 585
R151 B.n459 B.n458 585
R152 B.n456 B.n241 585
R153 B.n241 B.n240 585
R154 B.n455 B.n454 585
R155 B.n454 B.n453 585
R156 B.n243 B.n242 585
R157 B.n244 B.n243 585
R158 B.n446 B.n445 585
R159 B.n447 B.n446 585
R160 B.n444 B.n249 585
R161 B.n249 B.n248 585
R162 B.n443 B.n442 585
R163 B.n442 B.n441 585
R164 B.n251 B.n250 585
R165 B.n252 B.n251 585
R166 B.n434 B.n433 585
R167 B.n435 B.n434 585
R168 B.n432 B.n257 585
R169 B.n257 B.n256 585
R170 B.n431 B.n430 585
R171 B.n430 B.n429 585
R172 B.n259 B.n258 585
R173 B.n260 B.n259 585
R174 B.n425 B.n424 585
R175 B.n263 B.n262 585
R176 B.n421 B.n420 585
R177 B.n422 B.n421 585
R178 B.n419 B.n294 585
R179 B.n418 B.n417 585
R180 B.n416 B.n415 585
R181 B.n414 B.n413 585
R182 B.n412 B.n411 585
R183 B.n410 B.n409 585
R184 B.n408 B.n407 585
R185 B.n406 B.n405 585
R186 B.n404 B.n403 585
R187 B.n402 B.n401 585
R188 B.n400 B.n399 585
R189 B.n398 B.n397 585
R190 B.n396 B.n395 585
R191 B.n394 B.n393 585
R192 B.n392 B.n391 585
R193 B.n390 B.n389 585
R194 B.n388 B.n387 585
R195 B.n386 B.n385 585
R196 B.n384 B.n383 585
R197 B.n382 B.n381 585
R198 B.n380 B.n379 585
R199 B.n378 B.n377 585
R200 B.n376 B.n375 585
R201 B.n374 B.n373 585
R202 B.n372 B.n371 585
R203 B.n370 B.n369 585
R204 B.n368 B.n367 585
R205 B.n366 B.n365 585
R206 B.n364 B.n363 585
R207 B.n362 B.n361 585
R208 B.n360 B.n359 585
R209 B.n358 B.n357 585
R210 B.n356 B.n355 585
R211 B.n353 B.n352 585
R212 B.n351 B.n350 585
R213 B.n349 B.n348 585
R214 B.n347 B.n346 585
R215 B.n345 B.n344 585
R216 B.n343 B.n342 585
R217 B.n341 B.n340 585
R218 B.n339 B.n338 585
R219 B.n337 B.n336 585
R220 B.n335 B.n334 585
R221 B.n333 B.n332 585
R222 B.n331 B.n330 585
R223 B.n329 B.n328 585
R224 B.n327 B.n326 585
R225 B.n325 B.n324 585
R226 B.n323 B.n322 585
R227 B.n321 B.n320 585
R228 B.n319 B.n318 585
R229 B.n317 B.n316 585
R230 B.n315 B.n314 585
R231 B.n313 B.n312 585
R232 B.n311 B.n310 585
R233 B.n309 B.n308 585
R234 B.n307 B.n306 585
R235 B.n305 B.n304 585
R236 B.n303 B.n302 585
R237 B.n301 B.n300 585
R238 B.n426 B.n261 585
R239 B.n261 B.n260 585
R240 B.n428 B.n427 585
R241 B.n429 B.n428 585
R242 B.n255 B.n254 585
R243 B.n256 B.n255 585
R244 B.n437 B.n436 585
R245 B.n436 B.n435 585
R246 B.n438 B.n253 585
R247 B.n253 B.n252 585
R248 B.n440 B.n439 585
R249 B.n441 B.n440 585
R250 B.n247 B.n246 585
R251 B.n248 B.n247 585
R252 B.n449 B.n448 585
R253 B.n448 B.n447 585
R254 B.n450 B.n245 585
R255 B.n245 B.n244 585
R256 B.n452 B.n451 585
R257 B.n453 B.n452 585
R258 B.n239 B.n238 585
R259 B.n240 B.n239 585
R260 B.n461 B.n460 585
R261 B.n460 B.n459 585
R262 B.n462 B.n237 585
R263 B.n237 B.n236 585
R264 B.n464 B.n463 585
R265 B.n465 B.n464 585
R266 B.n231 B.n230 585
R267 B.n232 B.n231 585
R268 B.n473 B.n472 585
R269 B.n472 B.n471 585
R270 B.n474 B.n229 585
R271 B.n229 B.n228 585
R272 B.n476 B.n475 585
R273 B.n477 B.n476 585
R274 B.n223 B.n222 585
R275 B.n224 B.n223 585
R276 B.n486 B.n485 585
R277 B.n485 B.n484 585
R278 B.n487 B.n221 585
R279 B.n483 B.n221 585
R280 B.n489 B.n488 585
R281 B.n490 B.n489 585
R282 B.n216 B.n215 585
R283 B.n217 B.n216 585
R284 B.n499 B.n498 585
R285 B.n498 B.n497 585
R286 B.n500 B.n214 585
R287 B.n214 B.n213 585
R288 B.n502 B.n501 585
R289 B.n503 B.n502 585
R290 B.n2 B.n0 585
R291 B.n4 B.n2 585
R292 B.n3 B.n1 585
R293 B.n599 B.n3 585
R294 B.n597 B.n596 585
R295 B.n598 B.n597 585
R296 B.n595 B.n9 585
R297 B.n9 B.n8 585
R298 B.n594 B.n593 585
R299 B.n593 B.n592 585
R300 B.n11 B.n10 585
R301 B.n591 B.n11 585
R302 B.n589 B.n588 585
R303 B.n590 B.n589 585
R304 B.n587 B.n15 585
R305 B.n18 B.n15 585
R306 B.n586 B.n585 585
R307 B.n585 B.n584 585
R308 B.n17 B.n16 585
R309 B.n583 B.n17 585
R310 B.n581 B.n580 585
R311 B.n582 B.n581 585
R312 B.n579 B.n23 585
R313 B.n23 B.n22 585
R314 B.n578 B.n577 585
R315 B.n577 B.n576 585
R316 B.n25 B.n24 585
R317 B.n575 B.n25 585
R318 B.n573 B.n572 585
R319 B.n574 B.n573 585
R320 B.n571 B.n30 585
R321 B.n30 B.n29 585
R322 B.n570 B.n569 585
R323 B.n569 B.n568 585
R324 B.n32 B.n31 585
R325 B.n567 B.n32 585
R326 B.n565 B.n564 585
R327 B.n566 B.n565 585
R328 B.n563 B.n37 585
R329 B.n37 B.n36 585
R330 B.n562 B.n561 585
R331 B.n561 B.n560 585
R332 B.n39 B.n38 585
R333 B.n559 B.n39 585
R334 B.n557 B.n556 585
R335 B.n558 B.n557 585
R336 B.n555 B.n44 585
R337 B.n44 B.n43 585
R338 B.n554 B.n553 585
R339 B.n553 B.n552 585
R340 B.n46 B.n45 585
R341 B.n551 B.n46 585
R342 B.n549 B.n548 585
R343 B.n550 B.n549 585
R344 B.n547 B.n51 585
R345 B.n51 B.n50 585
R346 B.n602 B.n601 585
R347 B.n601 B.n600 585
R348 B.n424 B.n261 526.135
R349 B.n545 B.n51 526.135
R350 B.n300 B.n259 526.135
R351 B.n542 B.n85 526.135
R352 B.n298 B.t13 265.865
R353 B.n295 B.t9 265.865
R354 B.n89 B.t2 265.865
R355 B.n86 B.t6 265.865
R356 B.n543 B.n83 256.663
R357 B.n543 B.n82 256.663
R358 B.n543 B.n81 256.663
R359 B.n543 B.n80 256.663
R360 B.n543 B.n79 256.663
R361 B.n543 B.n78 256.663
R362 B.n543 B.n77 256.663
R363 B.n543 B.n76 256.663
R364 B.n543 B.n75 256.663
R365 B.n543 B.n74 256.663
R366 B.n543 B.n73 256.663
R367 B.n543 B.n72 256.663
R368 B.n543 B.n71 256.663
R369 B.n543 B.n70 256.663
R370 B.n543 B.n69 256.663
R371 B.n543 B.n68 256.663
R372 B.n543 B.n67 256.663
R373 B.n543 B.n66 256.663
R374 B.n543 B.n65 256.663
R375 B.n543 B.n64 256.663
R376 B.n543 B.n63 256.663
R377 B.n543 B.n62 256.663
R378 B.n543 B.n61 256.663
R379 B.n543 B.n60 256.663
R380 B.n543 B.n59 256.663
R381 B.n543 B.n58 256.663
R382 B.n543 B.n57 256.663
R383 B.n543 B.n56 256.663
R384 B.n543 B.n55 256.663
R385 B.n543 B.n54 256.663
R386 B.n544 B.n543 256.663
R387 B.n423 B.n422 256.663
R388 B.n422 B.n264 256.663
R389 B.n422 B.n265 256.663
R390 B.n422 B.n266 256.663
R391 B.n422 B.n267 256.663
R392 B.n422 B.n268 256.663
R393 B.n422 B.n269 256.663
R394 B.n422 B.n270 256.663
R395 B.n422 B.n271 256.663
R396 B.n422 B.n272 256.663
R397 B.n422 B.n273 256.663
R398 B.n422 B.n274 256.663
R399 B.n422 B.n275 256.663
R400 B.n422 B.n276 256.663
R401 B.n422 B.n277 256.663
R402 B.n422 B.n278 256.663
R403 B.n422 B.n279 256.663
R404 B.n422 B.n280 256.663
R405 B.n422 B.n281 256.663
R406 B.n422 B.n282 256.663
R407 B.n422 B.n283 256.663
R408 B.n422 B.n284 256.663
R409 B.n422 B.n285 256.663
R410 B.n422 B.n286 256.663
R411 B.n422 B.n287 256.663
R412 B.n422 B.n288 256.663
R413 B.n422 B.n289 256.663
R414 B.n422 B.n290 256.663
R415 B.n422 B.n291 256.663
R416 B.n422 B.n292 256.663
R417 B.n422 B.n293 256.663
R418 B.n428 B.n261 163.367
R419 B.n428 B.n255 163.367
R420 B.n436 B.n255 163.367
R421 B.n436 B.n253 163.367
R422 B.n440 B.n253 163.367
R423 B.n440 B.n247 163.367
R424 B.n448 B.n247 163.367
R425 B.n448 B.n245 163.367
R426 B.n452 B.n245 163.367
R427 B.n452 B.n239 163.367
R428 B.n460 B.n239 163.367
R429 B.n460 B.n237 163.367
R430 B.n464 B.n237 163.367
R431 B.n464 B.n231 163.367
R432 B.n472 B.n231 163.367
R433 B.n472 B.n229 163.367
R434 B.n476 B.n229 163.367
R435 B.n476 B.n223 163.367
R436 B.n485 B.n223 163.367
R437 B.n485 B.n221 163.367
R438 B.n489 B.n221 163.367
R439 B.n489 B.n216 163.367
R440 B.n498 B.n216 163.367
R441 B.n498 B.n214 163.367
R442 B.n502 B.n214 163.367
R443 B.n502 B.n2 163.367
R444 B.n601 B.n2 163.367
R445 B.n601 B.n3 163.367
R446 B.n597 B.n3 163.367
R447 B.n597 B.n9 163.367
R448 B.n593 B.n9 163.367
R449 B.n593 B.n11 163.367
R450 B.n589 B.n11 163.367
R451 B.n589 B.n15 163.367
R452 B.n585 B.n15 163.367
R453 B.n585 B.n17 163.367
R454 B.n581 B.n17 163.367
R455 B.n581 B.n23 163.367
R456 B.n577 B.n23 163.367
R457 B.n577 B.n25 163.367
R458 B.n573 B.n25 163.367
R459 B.n573 B.n30 163.367
R460 B.n569 B.n30 163.367
R461 B.n569 B.n32 163.367
R462 B.n565 B.n32 163.367
R463 B.n565 B.n37 163.367
R464 B.n561 B.n37 163.367
R465 B.n561 B.n39 163.367
R466 B.n557 B.n39 163.367
R467 B.n557 B.n44 163.367
R468 B.n553 B.n44 163.367
R469 B.n553 B.n46 163.367
R470 B.n549 B.n46 163.367
R471 B.n549 B.n51 163.367
R472 B.n421 B.n263 163.367
R473 B.n421 B.n294 163.367
R474 B.n417 B.n416 163.367
R475 B.n413 B.n412 163.367
R476 B.n409 B.n408 163.367
R477 B.n405 B.n404 163.367
R478 B.n401 B.n400 163.367
R479 B.n397 B.n396 163.367
R480 B.n393 B.n392 163.367
R481 B.n389 B.n388 163.367
R482 B.n385 B.n384 163.367
R483 B.n381 B.n380 163.367
R484 B.n377 B.n376 163.367
R485 B.n373 B.n372 163.367
R486 B.n369 B.n368 163.367
R487 B.n365 B.n364 163.367
R488 B.n361 B.n360 163.367
R489 B.n357 B.n356 163.367
R490 B.n352 B.n351 163.367
R491 B.n348 B.n347 163.367
R492 B.n344 B.n343 163.367
R493 B.n340 B.n339 163.367
R494 B.n336 B.n335 163.367
R495 B.n332 B.n331 163.367
R496 B.n328 B.n327 163.367
R497 B.n324 B.n323 163.367
R498 B.n320 B.n319 163.367
R499 B.n316 B.n315 163.367
R500 B.n312 B.n311 163.367
R501 B.n308 B.n307 163.367
R502 B.n304 B.n303 163.367
R503 B.n430 B.n259 163.367
R504 B.n430 B.n257 163.367
R505 B.n434 B.n257 163.367
R506 B.n434 B.n251 163.367
R507 B.n442 B.n251 163.367
R508 B.n442 B.n249 163.367
R509 B.n446 B.n249 163.367
R510 B.n446 B.n243 163.367
R511 B.n454 B.n243 163.367
R512 B.n454 B.n241 163.367
R513 B.n458 B.n241 163.367
R514 B.n458 B.n235 163.367
R515 B.n466 B.n235 163.367
R516 B.n466 B.n233 163.367
R517 B.n470 B.n233 163.367
R518 B.n470 B.n227 163.367
R519 B.n478 B.n227 163.367
R520 B.n478 B.n225 163.367
R521 B.n482 B.n225 163.367
R522 B.n482 B.n220 163.367
R523 B.n491 B.n220 163.367
R524 B.n491 B.n218 163.367
R525 B.n496 B.n218 163.367
R526 B.n496 B.n212 163.367
R527 B.n504 B.n212 163.367
R528 B.n505 B.n504 163.367
R529 B.n505 B.n5 163.367
R530 B.n6 B.n5 163.367
R531 B.n7 B.n6 163.367
R532 B.n510 B.n7 163.367
R533 B.n510 B.n12 163.367
R534 B.n13 B.n12 163.367
R535 B.n14 B.n13 163.367
R536 B.n515 B.n14 163.367
R537 B.n515 B.n19 163.367
R538 B.n20 B.n19 163.367
R539 B.n21 B.n20 163.367
R540 B.n520 B.n21 163.367
R541 B.n520 B.n26 163.367
R542 B.n27 B.n26 163.367
R543 B.n28 B.n27 163.367
R544 B.n525 B.n28 163.367
R545 B.n525 B.n33 163.367
R546 B.n34 B.n33 163.367
R547 B.n35 B.n34 163.367
R548 B.n530 B.n35 163.367
R549 B.n530 B.n40 163.367
R550 B.n41 B.n40 163.367
R551 B.n42 B.n41 163.367
R552 B.n535 B.n42 163.367
R553 B.n535 B.n47 163.367
R554 B.n48 B.n47 163.367
R555 B.n49 B.n48 163.367
R556 B.n85 B.n49 163.367
R557 B.n91 B.n53 163.367
R558 B.n95 B.n94 163.367
R559 B.n99 B.n98 163.367
R560 B.n103 B.n102 163.367
R561 B.n107 B.n106 163.367
R562 B.n111 B.n110 163.367
R563 B.n115 B.n114 163.367
R564 B.n119 B.n118 163.367
R565 B.n123 B.n122 163.367
R566 B.n127 B.n126 163.367
R567 B.n131 B.n130 163.367
R568 B.n135 B.n134 163.367
R569 B.n139 B.n138 163.367
R570 B.n144 B.n143 163.367
R571 B.n148 B.n147 163.367
R572 B.n152 B.n151 163.367
R573 B.n156 B.n155 163.367
R574 B.n160 B.n159 163.367
R575 B.n164 B.n163 163.367
R576 B.n168 B.n167 163.367
R577 B.n172 B.n171 163.367
R578 B.n176 B.n175 163.367
R579 B.n180 B.n179 163.367
R580 B.n184 B.n183 163.367
R581 B.n188 B.n187 163.367
R582 B.n192 B.n191 163.367
R583 B.n196 B.n195 163.367
R584 B.n200 B.n199 163.367
R585 B.n204 B.n203 163.367
R586 B.n208 B.n207 163.367
R587 B.n542 B.n84 163.367
R588 B.n298 B.t15 134.351
R589 B.n86 B.t7 134.351
R590 B.n295 B.t12 134.344
R591 B.n89 B.t4 134.344
R592 B.n422 B.n260 121.671
R593 B.n543 B.n50 121.671
R594 B.n424 B.n423 71.676
R595 B.n294 B.n264 71.676
R596 B.n416 B.n265 71.676
R597 B.n412 B.n266 71.676
R598 B.n408 B.n267 71.676
R599 B.n404 B.n268 71.676
R600 B.n400 B.n269 71.676
R601 B.n396 B.n270 71.676
R602 B.n392 B.n271 71.676
R603 B.n388 B.n272 71.676
R604 B.n384 B.n273 71.676
R605 B.n380 B.n274 71.676
R606 B.n376 B.n275 71.676
R607 B.n372 B.n276 71.676
R608 B.n368 B.n277 71.676
R609 B.n364 B.n278 71.676
R610 B.n360 B.n279 71.676
R611 B.n356 B.n280 71.676
R612 B.n351 B.n281 71.676
R613 B.n347 B.n282 71.676
R614 B.n343 B.n283 71.676
R615 B.n339 B.n284 71.676
R616 B.n335 B.n285 71.676
R617 B.n331 B.n286 71.676
R618 B.n327 B.n287 71.676
R619 B.n323 B.n288 71.676
R620 B.n319 B.n289 71.676
R621 B.n315 B.n290 71.676
R622 B.n311 B.n291 71.676
R623 B.n307 B.n292 71.676
R624 B.n303 B.n293 71.676
R625 B.n545 B.n544 71.676
R626 B.n91 B.n54 71.676
R627 B.n95 B.n55 71.676
R628 B.n99 B.n56 71.676
R629 B.n103 B.n57 71.676
R630 B.n107 B.n58 71.676
R631 B.n111 B.n59 71.676
R632 B.n115 B.n60 71.676
R633 B.n119 B.n61 71.676
R634 B.n123 B.n62 71.676
R635 B.n127 B.n63 71.676
R636 B.n131 B.n64 71.676
R637 B.n135 B.n65 71.676
R638 B.n139 B.n66 71.676
R639 B.n144 B.n67 71.676
R640 B.n148 B.n68 71.676
R641 B.n152 B.n69 71.676
R642 B.n156 B.n70 71.676
R643 B.n160 B.n71 71.676
R644 B.n164 B.n72 71.676
R645 B.n168 B.n73 71.676
R646 B.n172 B.n74 71.676
R647 B.n176 B.n75 71.676
R648 B.n180 B.n76 71.676
R649 B.n184 B.n77 71.676
R650 B.n188 B.n78 71.676
R651 B.n192 B.n79 71.676
R652 B.n196 B.n80 71.676
R653 B.n200 B.n81 71.676
R654 B.n204 B.n82 71.676
R655 B.n208 B.n83 71.676
R656 B.n84 B.n83 71.676
R657 B.n207 B.n82 71.676
R658 B.n203 B.n81 71.676
R659 B.n199 B.n80 71.676
R660 B.n195 B.n79 71.676
R661 B.n191 B.n78 71.676
R662 B.n187 B.n77 71.676
R663 B.n183 B.n76 71.676
R664 B.n179 B.n75 71.676
R665 B.n175 B.n74 71.676
R666 B.n171 B.n73 71.676
R667 B.n167 B.n72 71.676
R668 B.n163 B.n71 71.676
R669 B.n159 B.n70 71.676
R670 B.n155 B.n69 71.676
R671 B.n151 B.n68 71.676
R672 B.n147 B.n67 71.676
R673 B.n143 B.n66 71.676
R674 B.n138 B.n65 71.676
R675 B.n134 B.n64 71.676
R676 B.n130 B.n63 71.676
R677 B.n126 B.n62 71.676
R678 B.n122 B.n61 71.676
R679 B.n118 B.n60 71.676
R680 B.n114 B.n59 71.676
R681 B.n110 B.n58 71.676
R682 B.n106 B.n57 71.676
R683 B.n102 B.n56 71.676
R684 B.n98 B.n55 71.676
R685 B.n94 B.n54 71.676
R686 B.n544 B.n53 71.676
R687 B.n423 B.n263 71.676
R688 B.n417 B.n264 71.676
R689 B.n413 B.n265 71.676
R690 B.n409 B.n266 71.676
R691 B.n405 B.n267 71.676
R692 B.n401 B.n268 71.676
R693 B.n397 B.n269 71.676
R694 B.n393 B.n270 71.676
R695 B.n389 B.n271 71.676
R696 B.n385 B.n272 71.676
R697 B.n381 B.n273 71.676
R698 B.n377 B.n274 71.676
R699 B.n373 B.n275 71.676
R700 B.n369 B.n276 71.676
R701 B.n365 B.n277 71.676
R702 B.n361 B.n278 71.676
R703 B.n357 B.n279 71.676
R704 B.n352 B.n280 71.676
R705 B.n348 B.n281 71.676
R706 B.n344 B.n282 71.676
R707 B.n340 B.n283 71.676
R708 B.n336 B.n284 71.676
R709 B.n332 B.n285 71.676
R710 B.n328 B.n286 71.676
R711 B.n324 B.n287 71.676
R712 B.n320 B.n288 71.676
R713 B.n316 B.n289 71.676
R714 B.n312 B.n290 71.676
R715 B.n308 B.n291 71.676
R716 B.n304 B.n292 71.676
R717 B.n300 B.n293 71.676
R718 B.n299 B.t14 71.5148
R719 B.n87 B.t8 71.5148
R720 B.n296 B.t11 71.507
R721 B.n90 B.t5 71.507
R722 B.n299 B.n298 62.8369
R723 B.n296 B.n295 62.8369
R724 B.n90 B.n89 62.8369
R725 B.n87 B.n86 62.8369
R726 B.n429 B.n260 61.2869
R727 B.n429 B.n256 61.2869
R728 B.n435 B.n256 61.2869
R729 B.n435 B.n252 61.2869
R730 B.n441 B.n252 61.2869
R731 B.n441 B.n248 61.2869
R732 B.n447 B.n248 61.2869
R733 B.n453 B.n244 61.2869
R734 B.n453 B.n240 61.2869
R735 B.n459 B.n240 61.2869
R736 B.n459 B.n236 61.2869
R737 B.n465 B.n236 61.2869
R738 B.n465 B.n232 61.2869
R739 B.n471 B.n232 61.2869
R740 B.n471 B.n228 61.2869
R741 B.n477 B.n228 61.2869
R742 B.n477 B.n224 61.2869
R743 B.n484 B.n224 61.2869
R744 B.n484 B.n483 61.2869
R745 B.n490 B.n217 61.2869
R746 B.n497 B.n217 61.2869
R747 B.n497 B.n213 61.2869
R748 B.n503 B.n213 61.2869
R749 B.n503 B.n4 61.2869
R750 B.n600 B.n4 61.2869
R751 B.n600 B.n599 61.2869
R752 B.n599 B.n598 61.2869
R753 B.n598 B.n8 61.2869
R754 B.n592 B.n8 61.2869
R755 B.n592 B.n591 61.2869
R756 B.n591 B.n590 61.2869
R757 B.n584 B.n18 61.2869
R758 B.n584 B.n583 61.2869
R759 B.n583 B.n582 61.2869
R760 B.n582 B.n22 61.2869
R761 B.n576 B.n22 61.2869
R762 B.n576 B.n575 61.2869
R763 B.n575 B.n574 61.2869
R764 B.n574 B.n29 61.2869
R765 B.n568 B.n29 61.2869
R766 B.n568 B.n567 61.2869
R767 B.n567 B.n566 61.2869
R768 B.n566 B.n36 61.2869
R769 B.n560 B.n559 61.2869
R770 B.n559 B.n558 61.2869
R771 B.n558 B.n43 61.2869
R772 B.n552 B.n43 61.2869
R773 B.n552 B.n551 61.2869
R774 B.n551 B.n550 61.2869
R775 B.n550 B.n50 61.2869
R776 B.n354 B.n299 59.5399
R777 B.n297 B.n296 59.5399
R778 B.n141 B.n90 59.5399
R779 B.n88 B.n87 59.5399
R780 B.n447 B.t10 54.978
R781 B.n560 B.t3 54.978
R782 B.n483 B.t0 38.7551
R783 B.n18 B.t1 38.7551
R784 B.n547 B.n546 34.1859
R785 B.n541 B.n540 34.1859
R786 B.n301 B.n258 34.1859
R787 B.n426 B.n425 34.1859
R788 B.n490 B.t0 22.5322
R789 B.n590 B.t1 22.5322
R790 B B.n602 18.0485
R791 B.n546 B.n52 10.6151
R792 B.n92 B.n52 10.6151
R793 B.n93 B.n92 10.6151
R794 B.n96 B.n93 10.6151
R795 B.n97 B.n96 10.6151
R796 B.n100 B.n97 10.6151
R797 B.n101 B.n100 10.6151
R798 B.n104 B.n101 10.6151
R799 B.n105 B.n104 10.6151
R800 B.n108 B.n105 10.6151
R801 B.n109 B.n108 10.6151
R802 B.n112 B.n109 10.6151
R803 B.n113 B.n112 10.6151
R804 B.n116 B.n113 10.6151
R805 B.n117 B.n116 10.6151
R806 B.n120 B.n117 10.6151
R807 B.n121 B.n120 10.6151
R808 B.n124 B.n121 10.6151
R809 B.n125 B.n124 10.6151
R810 B.n128 B.n125 10.6151
R811 B.n129 B.n128 10.6151
R812 B.n132 B.n129 10.6151
R813 B.n133 B.n132 10.6151
R814 B.n136 B.n133 10.6151
R815 B.n137 B.n136 10.6151
R816 B.n140 B.n137 10.6151
R817 B.n145 B.n142 10.6151
R818 B.n146 B.n145 10.6151
R819 B.n149 B.n146 10.6151
R820 B.n150 B.n149 10.6151
R821 B.n153 B.n150 10.6151
R822 B.n154 B.n153 10.6151
R823 B.n157 B.n154 10.6151
R824 B.n158 B.n157 10.6151
R825 B.n162 B.n161 10.6151
R826 B.n165 B.n162 10.6151
R827 B.n166 B.n165 10.6151
R828 B.n169 B.n166 10.6151
R829 B.n170 B.n169 10.6151
R830 B.n173 B.n170 10.6151
R831 B.n174 B.n173 10.6151
R832 B.n177 B.n174 10.6151
R833 B.n178 B.n177 10.6151
R834 B.n181 B.n178 10.6151
R835 B.n182 B.n181 10.6151
R836 B.n185 B.n182 10.6151
R837 B.n186 B.n185 10.6151
R838 B.n189 B.n186 10.6151
R839 B.n190 B.n189 10.6151
R840 B.n193 B.n190 10.6151
R841 B.n194 B.n193 10.6151
R842 B.n197 B.n194 10.6151
R843 B.n198 B.n197 10.6151
R844 B.n201 B.n198 10.6151
R845 B.n202 B.n201 10.6151
R846 B.n205 B.n202 10.6151
R847 B.n206 B.n205 10.6151
R848 B.n209 B.n206 10.6151
R849 B.n210 B.n209 10.6151
R850 B.n541 B.n210 10.6151
R851 B.n431 B.n258 10.6151
R852 B.n432 B.n431 10.6151
R853 B.n433 B.n432 10.6151
R854 B.n433 B.n250 10.6151
R855 B.n443 B.n250 10.6151
R856 B.n444 B.n443 10.6151
R857 B.n445 B.n444 10.6151
R858 B.n445 B.n242 10.6151
R859 B.n455 B.n242 10.6151
R860 B.n456 B.n455 10.6151
R861 B.n457 B.n456 10.6151
R862 B.n457 B.n234 10.6151
R863 B.n467 B.n234 10.6151
R864 B.n468 B.n467 10.6151
R865 B.n469 B.n468 10.6151
R866 B.n469 B.n226 10.6151
R867 B.n479 B.n226 10.6151
R868 B.n480 B.n479 10.6151
R869 B.n481 B.n480 10.6151
R870 B.n481 B.n219 10.6151
R871 B.n492 B.n219 10.6151
R872 B.n493 B.n492 10.6151
R873 B.n495 B.n493 10.6151
R874 B.n495 B.n494 10.6151
R875 B.n494 B.n211 10.6151
R876 B.n506 B.n211 10.6151
R877 B.n507 B.n506 10.6151
R878 B.n508 B.n507 10.6151
R879 B.n509 B.n508 10.6151
R880 B.n511 B.n509 10.6151
R881 B.n512 B.n511 10.6151
R882 B.n513 B.n512 10.6151
R883 B.n514 B.n513 10.6151
R884 B.n516 B.n514 10.6151
R885 B.n517 B.n516 10.6151
R886 B.n518 B.n517 10.6151
R887 B.n519 B.n518 10.6151
R888 B.n521 B.n519 10.6151
R889 B.n522 B.n521 10.6151
R890 B.n523 B.n522 10.6151
R891 B.n524 B.n523 10.6151
R892 B.n526 B.n524 10.6151
R893 B.n527 B.n526 10.6151
R894 B.n528 B.n527 10.6151
R895 B.n529 B.n528 10.6151
R896 B.n531 B.n529 10.6151
R897 B.n532 B.n531 10.6151
R898 B.n533 B.n532 10.6151
R899 B.n534 B.n533 10.6151
R900 B.n536 B.n534 10.6151
R901 B.n537 B.n536 10.6151
R902 B.n538 B.n537 10.6151
R903 B.n539 B.n538 10.6151
R904 B.n540 B.n539 10.6151
R905 B.n425 B.n262 10.6151
R906 B.n420 B.n262 10.6151
R907 B.n420 B.n419 10.6151
R908 B.n419 B.n418 10.6151
R909 B.n418 B.n415 10.6151
R910 B.n415 B.n414 10.6151
R911 B.n414 B.n411 10.6151
R912 B.n411 B.n410 10.6151
R913 B.n410 B.n407 10.6151
R914 B.n407 B.n406 10.6151
R915 B.n406 B.n403 10.6151
R916 B.n403 B.n402 10.6151
R917 B.n402 B.n399 10.6151
R918 B.n399 B.n398 10.6151
R919 B.n398 B.n395 10.6151
R920 B.n395 B.n394 10.6151
R921 B.n394 B.n391 10.6151
R922 B.n391 B.n390 10.6151
R923 B.n390 B.n387 10.6151
R924 B.n387 B.n386 10.6151
R925 B.n386 B.n383 10.6151
R926 B.n383 B.n382 10.6151
R927 B.n382 B.n379 10.6151
R928 B.n379 B.n378 10.6151
R929 B.n378 B.n375 10.6151
R930 B.n375 B.n374 10.6151
R931 B.n371 B.n370 10.6151
R932 B.n370 B.n367 10.6151
R933 B.n367 B.n366 10.6151
R934 B.n366 B.n363 10.6151
R935 B.n363 B.n362 10.6151
R936 B.n362 B.n359 10.6151
R937 B.n359 B.n358 10.6151
R938 B.n358 B.n355 10.6151
R939 B.n353 B.n350 10.6151
R940 B.n350 B.n349 10.6151
R941 B.n349 B.n346 10.6151
R942 B.n346 B.n345 10.6151
R943 B.n345 B.n342 10.6151
R944 B.n342 B.n341 10.6151
R945 B.n341 B.n338 10.6151
R946 B.n338 B.n337 10.6151
R947 B.n337 B.n334 10.6151
R948 B.n334 B.n333 10.6151
R949 B.n333 B.n330 10.6151
R950 B.n330 B.n329 10.6151
R951 B.n329 B.n326 10.6151
R952 B.n326 B.n325 10.6151
R953 B.n325 B.n322 10.6151
R954 B.n322 B.n321 10.6151
R955 B.n321 B.n318 10.6151
R956 B.n318 B.n317 10.6151
R957 B.n317 B.n314 10.6151
R958 B.n314 B.n313 10.6151
R959 B.n313 B.n310 10.6151
R960 B.n310 B.n309 10.6151
R961 B.n309 B.n306 10.6151
R962 B.n306 B.n305 10.6151
R963 B.n305 B.n302 10.6151
R964 B.n302 B.n301 10.6151
R965 B.n427 B.n426 10.6151
R966 B.n427 B.n254 10.6151
R967 B.n437 B.n254 10.6151
R968 B.n438 B.n437 10.6151
R969 B.n439 B.n438 10.6151
R970 B.n439 B.n246 10.6151
R971 B.n449 B.n246 10.6151
R972 B.n450 B.n449 10.6151
R973 B.n451 B.n450 10.6151
R974 B.n451 B.n238 10.6151
R975 B.n461 B.n238 10.6151
R976 B.n462 B.n461 10.6151
R977 B.n463 B.n462 10.6151
R978 B.n463 B.n230 10.6151
R979 B.n473 B.n230 10.6151
R980 B.n474 B.n473 10.6151
R981 B.n475 B.n474 10.6151
R982 B.n475 B.n222 10.6151
R983 B.n486 B.n222 10.6151
R984 B.n487 B.n486 10.6151
R985 B.n488 B.n487 10.6151
R986 B.n488 B.n215 10.6151
R987 B.n499 B.n215 10.6151
R988 B.n500 B.n499 10.6151
R989 B.n501 B.n500 10.6151
R990 B.n501 B.n0 10.6151
R991 B.n596 B.n1 10.6151
R992 B.n596 B.n595 10.6151
R993 B.n595 B.n594 10.6151
R994 B.n594 B.n10 10.6151
R995 B.n588 B.n10 10.6151
R996 B.n588 B.n587 10.6151
R997 B.n587 B.n586 10.6151
R998 B.n586 B.n16 10.6151
R999 B.n580 B.n16 10.6151
R1000 B.n580 B.n579 10.6151
R1001 B.n579 B.n578 10.6151
R1002 B.n578 B.n24 10.6151
R1003 B.n572 B.n24 10.6151
R1004 B.n572 B.n571 10.6151
R1005 B.n571 B.n570 10.6151
R1006 B.n570 B.n31 10.6151
R1007 B.n564 B.n31 10.6151
R1008 B.n564 B.n563 10.6151
R1009 B.n563 B.n562 10.6151
R1010 B.n562 B.n38 10.6151
R1011 B.n556 B.n38 10.6151
R1012 B.n556 B.n555 10.6151
R1013 B.n555 B.n554 10.6151
R1014 B.n554 B.n45 10.6151
R1015 B.n548 B.n45 10.6151
R1016 B.n548 B.n547 10.6151
R1017 B.n142 B.n141 6.5566
R1018 B.n158 B.n88 6.5566
R1019 B.n371 B.n297 6.5566
R1020 B.n355 B.n354 6.5566
R1021 B.t10 B.n244 6.30939
R1022 B.t3 B.n36 6.30939
R1023 B.n141 B.n140 4.05904
R1024 B.n161 B.n88 4.05904
R1025 B.n374 B.n297 4.05904
R1026 B.n354 B.n353 4.05904
R1027 B.n602 B.n0 2.81026
R1028 B.n602 B.n1 2.81026
R1029 VN VN.t1 140.129
R1030 VN VN.t0 98.9203
R1031 VTAIL.n1 VTAIL.t3 55.271
R1032 VTAIL.n3 VTAIL.t2 55.2709
R1033 VTAIL.n0 VTAIL.t1 55.2709
R1034 VTAIL.n2 VTAIL.t0 55.2709
R1035 VTAIL.n1 VTAIL.n0 23.9272
R1036 VTAIL.n3 VTAIL.n2 21.1341
R1037 VTAIL.n2 VTAIL.n1 1.86688
R1038 VTAIL VTAIL.n0 1.22679
R1039 VTAIL VTAIL.n3 0.640586
R1040 VDD2.n0 VDD2.t1 107.169
R1041 VDD2.n0 VDD2.t0 71.9497
R1042 VDD2 VDD2.n0 0.756965
R1043 VP.n0 VP.t0 140.126
R1044 VP.n0 VP.t1 98.489
R1045 VP VP.n0 0.431811
R1046 VDD1 VDD1.t0 108.392
R1047 VDD1 VDD1.t1 72.7061
C0 VP VDD1 1.9334f
C1 VDD1 VTAIL 3.80228f
C2 VN VP 4.66216f
C3 VN VTAIL 1.74842f
C4 VN VDD1 0.148264f
C5 VP VDD2 0.345712f
C6 VDD2 VTAIL 3.85633f
C7 VDD1 VDD2 0.711635f
C8 VN VDD2 1.73753f
C9 VP VTAIL 1.76262f
C10 VDD2 B 3.588531f
C11 VDD1 B 5.5343f
C12 VTAIL B 5.215442f
C13 VN B 8.35279f
C14 VP B 6.307882f
C15 VDD1.t1 B 0.836503f
C16 VDD1.t0 B 1.12806f
C17 VP.t1 B 1.19944f
C18 VP.t0 B 1.53896f
C19 VP.n0 B 1.90843f
C20 VDD2.t1 B 1.1505f
C21 VDD2.t0 B 0.868419f
C22 VDD2.n0 B 1.77951f
C23 VTAIL.t1 B 0.903318f
C24 VTAIL.n0 B 1.0606f
C25 VTAIL.t3 B 0.903326f
C26 VTAIL.n1 B 1.09352f
C27 VTAIL.t0 B 0.903318f
C28 VTAIL.n2 B 0.94984f
C29 VTAIL.t2 B 0.903318f
C30 VTAIL.n3 B 0.886756f
C31 VN.t0 B 1.19454f
C32 VN.t1 B 1.53198f
.ends

