* NGSPICE file created from diff_pair_sample_0672.ext - technology: sky130A

.subckt diff_pair_sample_0672 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t7 VP.t0 VDD1.t0 w_n2476_n3408# sky130_fd_pr__pfet_01v8 ad=4.758 pd=25.18 as=2.013 ps=12.53 w=12.2 l=2.18
X1 VDD1.t3 VP.t1 VTAIL.t6 w_n2476_n3408# sky130_fd_pr__pfet_01v8 ad=2.013 pd=12.53 as=4.758 ps=25.18 w=12.2 l=2.18
X2 VDD1.t1 VP.t2 VTAIL.t5 w_n2476_n3408# sky130_fd_pr__pfet_01v8 ad=2.013 pd=12.53 as=4.758 ps=25.18 w=12.2 l=2.18
X3 VTAIL.t1 VN.t0 VDD2.t3 w_n2476_n3408# sky130_fd_pr__pfet_01v8 ad=4.758 pd=25.18 as=2.013 ps=12.53 w=12.2 l=2.18
X4 VTAIL.t4 VP.t3 VDD1.t2 w_n2476_n3408# sky130_fd_pr__pfet_01v8 ad=4.758 pd=25.18 as=2.013 ps=12.53 w=12.2 l=2.18
X5 VDD2.t2 VN.t1 VTAIL.t2 w_n2476_n3408# sky130_fd_pr__pfet_01v8 ad=2.013 pd=12.53 as=4.758 ps=25.18 w=12.2 l=2.18
X6 B.t11 B.t9 B.t10 w_n2476_n3408# sky130_fd_pr__pfet_01v8 ad=4.758 pd=25.18 as=0 ps=0 w=12.2 l=2.18
X7 VDD2.t1 VN.t2 VTAIL.t3 w_n2476_n3408# sky130_fd_pr__pfet_01v8 ad=2.013 pd=12.53 as=4.758 ps=25.18 w=12.2 l=2.18
X8 B.t8 B.t6 B.t7 w_n2476_n3408# sky130_fd_pr__pfet_01v8 ad=4.758 pd=25.18 as=0 ps=0 w=12.2 l=2.18
X9 VTAIL.t0 VN.t3 VDD2.t0 w_n2476_n3408# sky130_fd_pr__pfet_01v8 ad=4.758 pd=25.18 as=2.013 ps=12.53 w=12.2 l=2.18
X10 B.t5 B.t3 B.t4 w_n2476_n3408# sky130_fd_pr__pfet_01v8 ad=4.758 pd=25.18 as=0 ps=0 w=12.2 l=2.18
X11 B.t2 B.t0 B.t1 w_n2476_n3408# sky130_fd_pr__pfet_01v8 ad=4.758 pd=25.18 as=0 ps=0 w=12.2 l=2.18
R0 VP.n3 VP.t3 170.489
R1 VP.n3 VP.t1 169.856
R2 VP.n12 VP.n0 161.3
R3 VP.n11 VP.n10 161.3
R4 VP.n9 VP.n1 161.3
R5 VP.n8 VP.n7 161.3
R6 VP.n6 VP.n2 161.3
R7 VP.n5 VP.t0 134.873
R8 VP.n13 VP.t2 134.873
R9 VP.n5 VP.n4 98.3664
R10 VP.n14 VP.n13 98.3664
R11 VP.n4 VP.n3 50.9621
R12 VP.n7 VP.n1 40.577
R13 VP.n11 VP.n1 40.577
R14 VP.n7 VP.n6 24.5923
R15 VP.n12 VP.n11 24.5923
R16 VP.n6 VP.n5 12.5423
R17 VP.n13 VP.n12 12.5423
R18 VP.n4 VP.n2 0.278335
R19 VP.n14 VP.n0 0.278335
R20 VP.n8 VP.n2 0.189894
R21 VP.n9 VP.n8 0.189894
R22 VP.n10 VP.n9 0.189894
R23 VP.n10 VP.n0 0.189894
R24 VP VP.n14 0.153485
R25 VDD1 VDD1.n1 116.638
R26 VDD1 VDD1.n0 75.4487
R27 VDD1.n0 VDD1.t2 2.66484
R28 VDD1.n0 VDD1.t3 2.66484
R29 VDD1.n1 VDD1.t0 2.66484
R30 VDD1.n1 VDD1.t1 2.66484
R31 VTAIL.n522 VTAIL.n462 756.745
R32 VTAIL.n60 VTAIL.n0 756.745
R33 VTAIL.n126 VTAIL.n66 756.745
R34 VTAIL.n192 VTAIL.n132 756.745
R35 VTAIL.n456 VTAIL.n396 756.745
R36 VTAIL.n390 VTAIL.n330 756.745
R37 VTAIL.n324 VTAIL.n264 756.745
R38 VTAIL.n258 VTAIL.n198 756.745
R39 VTAIL.n482 VTAIL.n481 585
R40 VTAIL.n487 VTAIL.n486 585
R41 VTAIL.n489 VTAIL.n488 585
R42 VTAIL.n478 VTAIL.n477 585
R43 VTAIL.n495 VTAIL.n494 585
R44 VTAIL.n497 VTAIL.n496 585
R45 VTAIL.n474 VTAIL.n473 585
R46 VTAIL.n504 VTAIL.n503 585
R47 VTAIL.n505 VTAIL.n472 585
R48 VTAIL.n507 VTAIL.n506 585
R49 VTAIL.n470 VTAIL.n469 585
R50 VTAIL.n513 VTAIL.n512 585
R51 VTAIL.n515 VTAIL.n514 585
R52 VTAIL.n466 VTAIL.n465 585
R53 VTAIL.n521 VTAIL.n520 585
R54 VTAIL.n523 VTAIL.n522 585
R55 VTAIL.n20 VTAIL.n19 585
R56 VTAIL.n25 VTAIL.n24 585
R57 VTAIL.n27 VTAIL.n26 585
R58 VTAIL.n16 VTAIL.n15 585
R59 VTAIL.n33 VTAIL.n32 585
R60 VTAIL.n35 VTAIL.n34 585
R61 VTAIL.n12 VTAIL.n11 585
R62 VTAIL.n42 VTAIL.n41 585
R63 VTAIL.n43 VTAIL.n10 585
R64 VTAIL.n45 VTAIL.n44 585
R65 VTAIL.n8 VTAIL.n7 585
R66 VTAIL.n51 VTAIL.n50 585
R67 VTAIL.n53 VTAIL.n52 585
R68 VTAIL.n4 VTAIL.n3 585
R69 VTAIL.n59 VTAIL.n58 585
R70 VTAIL.n61 VTAIL.n60 585
R71 VTAIL.n86 VTAIL.n85 585
R72 VTAIL.n91 VTAIL.n90 585
R73 VTAIL.n93 VTAIL.n92 585
R74 VTAIL.n82 VTAIL.n81 585
R75 VTAIL.n99 VTAIL.n98 585
R76 VTAIL.n101 VTAIL.n100 585
R77 VTAIL.n78 VTAIL.n77 585
R78 VTAIL.n108 VTAIL.n107 585
R79 VTAIL.n109 VTAIL.n76 585
R80 VTAIL.n111 VTAIL.n110 585
R81 VTAIL.n74 VTAIL.n73 585
R82 VTAIL.n117 VTAIL.n116 585
R83 VTAIL.n119 VTAIL.n118 585
R84 VTAIL.n70 VTAIL.n69 585
R85 VTAIL.n125 VTAIL.n124 585
R86 VTAIL.n127 VTAIL.n126 585
R87 VTAIL.n152 VTAIL.n151 585
R88 VTAIL.n157 VTAIL.n156 585
R89 VTAIL.n159 VTAIL.n158 585
R90 VTAIL.n148 VTAIL.n147 585
R91 VTAIL.n165 VTAIL.n164 585
R92 VTAIL.n167 VTAIL.n166 585
R93 VTAIL.n144 VTAIL.n143 585
R94 VTAIL.n174 VTAIL.n173 585
R95 VTAIL.n175 VTAIL.n142 585
R96 VTAIL.n177 VTAIL.n176 585
R97 VTAIL.n140 VTAIL.n139 585
R98 VTAIL.n183 VTAIL.n182 585
R99 VTAIL.n185 VTAIL.n184 585
R100 VTAIL.n136 VTAIL.n135 585
R101 VTAIL.n191 VTAIL.n190 585
R102 VTAIL.n193 VTAIL.n192 585
R103 VTAIL.n457 VTAIL.n456 585
R104 VTAIL.n455 VTAIL.n454 585
R105 VTAIL.n400 VTAIL.n399 585
R106 VTAIL.n449 VTAIL.n448 585
R107 VTAIL.n447 VTAIL.n446 585
R108 VTAIL.n404 VTAIL.n403 585
R109 VTAIL.n441 VTAIL.n440 585
R110 VTAIL.n439 VTAIL.n406 585
R111 VTAIL.n438 VTAIL.n437 585
R112 VTAIL.n409 VTAIL.n407 585
R113 VTAIL.n432 VTAIL.n431 585
R114 VTAIL.n430 VTAIL.n429 585
R115 VTAIL.n413 VTAIL.n412 585
R116 VTAIL.n424 VTAIL.n423 585
R117 VTAIL.n422 VTAIL.n421 585
R118 VTAIL.n417 VTAIL.n416 585
R119 VTAIL.n391 VTAIL.n390 585
R120 VTAIL.n389 VTAIL.n388 585
R121 VTAIL.n334 VTAIL.n333 585
R122 VTAIL.n383 VTAIL.n382 585
R123 VTAIL.n381 VTAIL.n380 585
R124 VTAIL.n338 VTAIL.n337 585
R125 VTAIL.n375 VTAIL.n374 585
R126 VTAIL.n373 VTAIL.n340 585
R127 VTAIL.n372 VTAIL.n371 585
R128 VTAIL.n343 VTAIL.n341 585
R129 VTAIL.n366 VTAIL.n365 585
R130 VTAIL.n364 VTAIL.n363 585
R131 VTAIL.n347 VTAIL.n346 585
R132 VTAIL.n358 VTAIL.n357 585
R133 VTAIL.n356 VTAIL.n355 585
R134 VTAIL.n351 VTAIL.n350 585
R135 VTAIL.n325 VTAIL.n324 585
R136 VTAIL.n323 VTAIL.n322 585
R137 VTAIL.n268 VTAIL.n267 585
R138 VTAIL.n317 VTAIL.n316 585
R139 VTAIL.n315 VTAIL.n314 585
R140 VTAIL.n272 VTAIL.n271 585
R141 VTAIL.n309 VTAIL.n308 585
R142 VTAIL.n307 VTAIL.n274 585
R143 VTAIL.n306 VTAIL.n305 585
R144 VTAIL.n277 VTAIL.n275 585
R145 VTAIL.n300 VTAIL.n299 585
R146 VTAIL.n298 VTAIL.n297 585
R147 VTAIL.n281 VTAIL.n280 585
R148 VTAIL.n292 VTAIL.n291 585
R149 VTAIL.n290 VTAIL.n289 585
R150 VTAIL.n285 VTAIL.n284 585
R151 VTAIL.n259 VTAIL.n258 585
R152 VTAIL.n257 VTAIL.n256 585
R153 VTAIL.n202 VTAIL.n201 585
R154 VTAIL.n251 VTAIL.n250 585
R155 VTAIL.n249 VTAIL.n248 585
R156 VTAIL.n206 VTAIL.n205 585
R157 VTAIL.n243 VTAIL.n242 585
R158 VTAIL.n241 VTAIL.n208 585
R159 VTAIL.n240 VTAIL.n239 585
R160 VTAIL.n211 VTAIL.n209 585
R161 VTAIL.n234 VTAIL.n233 585
R162 VTAIL.n232 VTAIL.n231 585
R163 VTAIL.n215 VTAIL.n214 585
R164 VTAIL.n226 VTAIL.n225 585
R165 VTAIL.n224 VTAIL.n223 585
R166 VTAIL.n219 VTAIL.n218 585
R167 VTAIL.n483 VTAIL.t3 329.036
R168 VTAIL.n21 VTAIL.t0 329.036
R169 VTAIL.n87 VTAIL.t5 329.036
R170 VTAIL.n153 VTAIL.t7 329.036
R171 VTAIL.n418 VTAIL.t6 329.036
R172 VTAIL.n352 VTAIL.t4 329.036
R173 VTAIL.n286 VTAIL.t2 329.036
R174 VTAIL.n220 VTAIL.t1 329.036
R175 VTAIL.n487 VTAIL.n481 171.744
R176 VTAIL.n488 VTAIL.n487 171.744
R177 VTAIL.n488 VTAIL.n477 171.744
R178 VTAIL.n495 VTAIL.n477 171.744
R179 VTAIL.n496 VTAIL.n495 171.744
R180 VTAIL.n496 VTAIL.n473 171.744
R181 VTAIL.n504 VTAIL.n473 171.744
R182 VTAIL.n505 VTAIL.n504 171.744
R183 VTAIL.n506 VTAIL.n505 171.744
R184 VTAIL.n506 VTAIL.n469 171.744
R185 VTAIL.n513 VTAIL.n469 171.744
R186 VTAIL.n514 VTAIL.n513 171.744
R187 VTAIL.n514 VTAIL.n465 171.744
R188 VTAIL.n521 VTAIL.n465 171.744
R189 VTAIL.n522 VTAIL.n521 171.744
R190 VTAIL.n25 VTAIL.n19 171.744
R191 VTAIL.n26 VTAIL.n25 171.744
R192 VTAIL.n26 VTAIL.n15 171.744
R193 VTAIL.n33 VTAIL.n15 171.744
R194 VTAIL.n34 VTAIL.n33 171.744
R195 VTAIL.n34 VTAIL.n11 171.744
R196 VTAIL.n42 VTAIL.n11 171.744
R197 VTAIL.n43 VTAIL.n42 171.744
R198 VTAIL.n44 VTAIL.n43 171.744
R199 VTAIL.n44 VTAIL.n7 171.744
R200 VTAIL.n51 VTAIL.n7 171.744
R201 VTAIL.n52 VTAIL.n51 171.744
R202 VTAIL.n52 VTAIL.n3 171.744
R203 VTAIL.n59 VTAIL.n3 171.744
R204 VTAIL.n60 VTAIL.n59 171.744
R205 VTAIL.n91 VTAIL.n85 171.744
R206 VTAIL.n92 VTAIL.n91 171.744
R207 VTAIL.n92 VTAIL.n81 171.744
R208 VTAIL.n99 VTAIL.n81 171.744
R209 VTAIL.n100 VTAIL.n99 171.744
R210 VTAIL.n100 VTAIL.n77 171.744
R211 VTAIL.n108 VTAIL.n77 171.744
R212 VTAIL.n109 VTAIL.n108 171.744
R213 VTAIL.n110 VTAIL.n109 171.744
R214 VTAIL.n110 VTAIL.n73 171.744
R215 VTAIL.n117 VTAIL.n73 171.744
R216 VTAIL.n118 VTAIL.n117 171.744
R217 VTAIL.n118 VTAIL.n69 171.744
R218 VTAIL.n125 VTAIL.n69 171.744
R219 VTAIL.n126 VTAIL.n125 171.744
R220 VTAIL.n157 VTAIL.n151 171.744
R221 VTAIL.n158 VTAIL.n157 171.744
R222 VTAIL.n158 VTAIL.n147 171.744
R223 VTAIL.n165 VTAIL.n147 171.744
R224 VTAIL.n166 VTAIL.n165 171.744
R225 VTAIL.n166 VTAIL.n143 171.744
R226 VTAIL.n174 VTAIL.n143 171.744
R227 VTAIL.n175 VTAIL.n174 171.744
R228 VTAIL.n176 VTAIL.n175 171.744
R229 VTAIL.n176 VTAIL.n139 171.744
R230 VTAIL.n183 VTAIL.n139 171.744
R231 VTAIL.n184 VTAIL.n183 171.744
R232 VTAIL.n184 VTAIL.n135 171.744
R233 VTAIL.n191 VTAIL.n135 171.744
R234 VTAIL.n192 VTAIL.n191 171.744
R235 VTAIL.n456 VTAIL.n455 171.744
R236 VTAIL.n455 VTAIL.n399 171.744
R237 VTAIL.n448 VTAIL.n399 171.744
R238 VTAIL.n448 VTAIL.n447 171.744
R239 VTAIL.n447 VTAIL.n403 171.744
R240 VTAIL.n440 VTAIL.n403 171.744
R241 VTAIL.n440 VTAIL.n439 171.744
R242 VTAIL.n439 VTAIL.n438 171.744
R243 VTAIL.n438 VTAIL.n407 171.744
R244 VTAIL.n431 VTAIL.n407 171.744
R245 VTAIL.n431 VTAIL.n430 171.744
R246 VTAIL.n430 VTAIL.n412 171.744
R247 VTAIL.n423 VTAIL.n412 171.744
R248 VTAIL.n423 VTAIL.n422 171.744
R249 VTAIL.n422 VTAIL.n416 171.744
R250 VTAIL.n390 VTAIL.n389 171.744
R251 VTAIL.n389 VTAIL.n333 171.744
R252 VTAIL.n382 VTAIL.n333 171.744
R253 VTAIL.n382 VTAIL.n381 171.744
R254 VTAIL.n381 VTAIL.n337 171.744
R255 VTAIL.n374 VTAIL.n337 171.744
R256 VTAIL.n374 VTAIL.n373 171.744
R257 VTAIL.n373 VTAIL.n372 171.744
R258 VTAIL.n372 VTAIL.n341 171.744
R259 VTAIL.n365 VTAIL.n341 171.744
R260 VTAIL.n365 VTAIL.n364 171.744
R261 VTAIL.n364 VTAIL.n346 171.744
R262 VTAIL.n357 VTAIL.n346 171.744
R263 VTAIL.n357 VTAIL.n356 171.744
R264 VTAIL.n356 VTAIL.n350 171.744
R265 VTAIL.n324 VTAIL.n323 171.744
R266 VTAIL.n323 VTAIL.n267 171.744
R267 VTAIL.n316 VTAIL.n267 171.744
R268 VTAIL.n316 VTAIL.n315 171.744
R269 VTAIL.n315 VTAIL.n271 171.744
R270 VTAIL.n308 VTAIL.n271 171.744
R271 VTAIL.n308 VTAIL.n307 171.744
R272 VTAIL.n307 VTAIL.n306 171.744
R273 VTAIL.n306 VTAIL.n275 171.744
R274 VTAIL.n299 VTAIL.n275 171.744
R275 VTAIL.n299 VTAIL.n298 171.744
R276 VTAIL.n298 VTAIL.n280 171.744
R277 VTAIL.n291 VTAIL.n280 171.744
R278 VTAIL.n291 VTAIL.n290 171.744
R279 VTAIL.n290 VTAIL.n284 171.744
R280 VTAIL.n258 VTAIL.n257 171.744
R281 VTAIL.n257 VTAIL.n201 171.744
R282 VTAIL.n250 VTAIL.n201 171.744
R283 VTAIL.n250 VTAIL.n249 171.744
R284 VTAIL.n249 VTAIL.n205 171.744
R285 VTAIL.n242 VTAIL.n205 171.744
R286 VTAIL.n242 VTAIL.n241 171.744
R287 VTAIL.n241 VTAIL.n240 171.744
R288 VTAIL.n240 VTAIL.n209 171.744
R289 VTAIL.n233 VTAIL.n209 171.744
R290 VTAIL.n233 VTAIL.n232 171.744
R291 VTAIL.n232 VTAIL.n214 171.744
R292 VTAIL.n225 VTAIL.n214 171.744
R293 VTAIL.n225 VTAIL.n224 171.744
R294 VTAIL.n224 VTAIL.n218 171.744
R295 VTAIL.t3 VTAIL.n481 85.8723
R296 VTAIL.t0 VTAIL.n19 85.8723
R297 VTAIL.t5 VTAIL.n85 85.8723
R298 VTAIL.t7 VTAIL.n151 85.8723
R299 VTAIL.t6 VTAIL.n416 85.8723
R300 VTAIL.t4 VTAIL.n350 85.8723
R301 VTAIL.t2 VTAIL.n284 85.8723
R302 VTAIL.t1 VTAIL.n218 85.8723
R303 VTAIL.n527 VTAIL.n526 33.7369
R304 VTAIL.n65 VTAIL.n64 33.7369
R305 VTAIL.n131 VTAIL.n130 33.7369
R306 VTAIL.n197 VTAIL.n196 33.7369
R307 VTAIL.n461 VTAIL.n460 33.7369
R308 VTAIL.n395 VTAIL.n394 33.7369
R309 VTAIL.n329 VTAIL.n328 33.7369
R310 VTAIL.n263 VTAIL.n262 33.7369
R311 VTAIL.n527 VTAIL.n461 25.0479
R312 VTAIL.n263 VTAIL.n197 25.0479
R313 VTAIL.n507 VTAIL.n472 13.1884
R314 VTAIL.n45 VTAIL.n10 13.1884
R315 VTAIL.n111 VTAIL.n76 13.1884
R316 VTAIL.n177 VTAIL.n142 13.1884
R317 VTAIL.n441 VTAIL.n406 13.1884
R318 VTAIL.n375 VTAIL.n340 13.1884
R319 VTAIL.n309 VTAIL.n274 13.1884
R320 VTAIL.n243 VTAIL.n208 13.1884
R321 VTAIL.n503 VTAIL.n502 12.8005
R322 VTAIL.n508 VTAIL.n470 12.8005
R323 VTAIL.n41 VTAIL.n40 12.8005
R324 VTAIL.n46 VTAIL.n8 12.8005
R325 VTAIL.n107 VTAIL.n106 12.8005
R326 VTAIL.n112 VTAIL.n74 12.8005
R327 VTAIL.n173 VTAIL.n172 12.8005
R328 VTAIL.n178 VTAIL.n140 12.8005
R329 VTAIL.n442 VTAIL.n404 12.8005
R330 VTAIL.n437 VTAIL.n408 12.8005
R331 VTAIL.n376 VTAIL.n338 12.8005
R332 VTAIL.n371 VTAIL.n342 12.8005
R333 VTAIL.n310 VTAIL.n272 12.8005
R334 VTAIL.n305 VTAIL.n276 12.8005
R335 VTAIL.n244 VTAIL.n206 12.8005
R336 VTAIL.n239 VTAIL.n210 12.8005
R337 VTAIL.n501 VTAIL.n474 12.0247
R338 VTAIL.n512 VTAIL.n511 12.0247
R339 VTAIL.n39 VTAIL.n12 12.0247
R340 VTAIL.n50 VTAIL.n49 12.0247
R341 VTAIL.n105 VTAIL.n78 12.0247
R342 VTAIL.n116 VTAIL.n115 12.0247
R343 VTAIL.n171 VTAIL.n144 12.0247
R344 VTAIL.n182 VTAIL.n181 12.0247
R345 VTAIL.n446 VTAIL.n445 12.0247
R346 VTAIL.n436 VTAIL.n409 12.0247
R347 VTAIL.n380 VTAIL.n379 12.0247
R348 VTAIL.n370 VTAIL.n343 12.0247
R349 VTAIL.n314 VTAIL.n313 12.0247
R350 VTAIL.n304 VTAIL.n277 12.0247
R351 VTAIL.n248 VTAIL.n247 12.0247
R352 VTAIL.n238 VTAIL.n211 12.0247
R353 VTAIL.n498 VTAIL.n497 11.249
R354 VTAIL.n515 VTAIL.n468 11.249
R355 VTAIL.n36 VTAIL.n35 11.249
R356 VTAIL.n53 VTAIL.n6 11.249
R357 VTAIL.n102 VTAIL.n101 11.249
R358 VTAIL.n119 VTAIL.n72 11.249
R359 VTAIL.n168 VTAIL.n167 11.249
R360 VTAIL.n185 VTAIL.n138 11.249
R361 VTAIL.n449 VTAIL.n402 11.249
R362 VTAIL.n433 VTAIL.n432 11.249
R363 VTAIL.n383 VTAIL.n336 11.249
R364 VTAIL.n367 VTAIL.n366 11.249
R365 VTAIL.n317 VTAIL.n270 11.249
R366 VTAIL.n301 VTAIL.n300 11.249
R367 VTAIL.n251 VTAIL.n204 11.249
R368 VTAIL.n235 VTAIL.n234 11.249
R369 VTAIL.n483 VTAIL.n482 10.7239
R370 VTAIL.n21 VTAIL.n20 10.7239
R371 VTAIL.n87 VTAIL.n86 10.7239
R372 VTAIL.n153 VTAIL.n152 10.7239
R373 VTAIL.n418 VTAIL.n417 10.7239
R374 VTAIL.n352 VTAIL.n351 10.7239
R375 VTAIL.n286 VTAIL.n285 10.7239
R376 VTAIL.n220 VTAIL.n219 10.7239
R377 VTAIL.n494 VTAIL.n476 10.4732
R378 VTAIL.n516 VTAIL.n466 10.4732
R379 VTAIL.n32 VTAIL.n14 10.4732
R380 VTAIL.n54 VTAIL.n4 10.4732
R381 VTAIL.n98 VTAIL.n80 10.4732
R382 VTAIL.n120 VTAIL.n70 10.4732
R383 VTAIL.n164 VTAIL.n146 10.4732
R384 VTAIL.n186 VTAIL.n136 10.4732
R385 VTAIL.n450 VTAIL.n400 10.4732
R386 VTAIL.n429 VTAIL.n411 10.4732
R387 VTAIL.n384 VTAIL.n334 10.4732
R388 VTAIL.n363 VTAIL.n345 10.4732
R389 VTAIL.n318 VTAIL.n268 10.4732
R390 VTAIL.n297 VTAIL.n279 10.4732
R391 VTAIL.n252 VTAIL.n202 10.4732
R392 VTAIL.n231 VTAIL.n213 10.4732
R393 VTAIL.n493 VTAIL.n478 9.69747
R394 VTAIL.n520 VTAIL.n519 9.69747
R395 VTAIL.n31 VTAIL.n16 9.69747
R396 VTAIL.n58 VTAIL.n57 9.69747
R397 VTAIL.n97 VTAIL.n82 9.69747
R398 VTAIL.n124 VTAIL.n123 9.69747
R399 VTAIL.n163 VTAIL.n148 9.69747
R400 VTAIL.n190 VTAIL.n189 9.69747
R401 VTAIL.n454 VTAIL.n453 9.69747
R402 VTAIL.n428 VTAIL.n413 9.69747
R403 VTAIL.n388 VTAIL.n387 9.69747
R404 VTAIL.n362 VTAIL.n347 9.69747
R405 VTAIL.n322 VTAIL.n321 9.69747
R406 VTAIL.n296 VTAIL.n281 9.69747
R407 VTAIL.n256 VTAIL.n255 9.69747
R408 VTAIL.n230 VTAIL.n215 9.69747
R409 VTAIL.n526 VTAIL.n525 9.45567
R410 VTAIL.n64 VTAIL.n63 9.45567
R411 VTAIL.n130 VTAIL.n129 9.45567
R412 VTAIL.n196 VTAIL.n195 9.45567
R413 VTAIL.n460 VTAIL.n459 9.45567
R414 VTAIL.n394 VTAIL.n393 9.45567
R415 VTAIL.n328 VTAIL.n327 9.45567
R416 VTAIL.n262 VTAIL.n261 9.45567
R417 VTAIL.n525 VTAIL.n524 9.3005
R418 VTAIL.n464 VTAIL.n463 9.3005
R419 VTAIL.n519 VTAIL.n518 9.3005
R420 VTAIL.n517 VTAIL.n516 9.3005
R421 VTAIL.n468 VTAIL.n467 9.3005
R422 VTAIL.n511 VTAIL.n510 9.3005
R423 VTAIL.n509 VTAIL.n508 9.3005
R424 VTAIL.n485 VTAIL.n484 9.3005
R425 VTAIL.n480 VTAIL.n479 9.3005
R426 VTAIL.n491 VTAIL.n490 9.3005
R427 VTAIL.n493 VTAIL.n492 9.3005
R428 VTAIL.n476 VTAIL.n475 9.3005
R429 VTAIL.n499 VTAIL.n498 9.3005
R430 VTAIL.n501 VTAIL.n500 9.3005
R431 VTAIL.n502 VTAIL.n471 9.3005
R432 VTAIL.n63 VTAIL.n62 9.3005
R433 VTAIL.n2 VTAIL.n1 9.3005
R434 VTAIL.n57 VTAIL.n56 9.3005
R435 VTAIL.n55 VTAIL.n54 9.3005
R436 VTAIL.n6 VTAIL.n5 9.3005
R437 VTAIL.n49 VTAIL.n48 9.3005
R438 VTAIL.n47 VTAIL.n46 9.3005
R439 VTAIL.n23 VTAIL.n22 9.3005
R440 VTAIL.n18 VTAIL.n17 9.3005
R441 VTAIL.n29 VTAIL.n28 9.3005
R442 VTAIL.n31 VTAIL.n30 9.3005
R443 VTAIL.n14 VTAIL.n13 9.3005
R444 VTAIL.n37 VTAIL.n36 9.3005
R445 VTAIL.n39 VTAIL.n38 9.3005
R446 VTAIL.n40 VTAIL.n9 9.3005
R447 VTAIL.n129 VTAIL.n128 9.3005
R448 VTAIL.n68 VTAIL.n67 9.3005
R449 VTAIL.n123 VTAIL.n122 9.3005
R450 VTAIL.n121 VTAIL.n120 9.3005
R451 VTAIL.n72 VTAIL.n71 9.3005
R452 VTAIL.n115 VTAIL.n114 9.3005
R453 VTAIL.n113 VTAIL.n112 9.3005
R454 VTAIL.n89 VTAIL.n88 9.3005
R455 VTAIL.n84 VTAIL.n83 9.3005
R456 VTAIL.n95 VTAIL.n94 9.3005
R457 VTAIL.n97 VTAIL.n96 9.3005
R458 VTAIL.n80 VTAIL.n79 9.3005
R459 VTAIL.n103 VTAIL.n102 9.3005
R460 VTAIL.n105 VTAIL.n104 9.3005
R461 VTAIL.n106 VTAIL.n75 9.3005
R462 VTAIL.n195 VTAIL.n194 9.3005
R463 VTAIL.n134 VTAIL.n133 9.3005
R464 VTAIL.n189 VTAIL.n188 9.3005
R465 VTAIL.n187 VTAIL.n186 9.3005
R466 VTAIL.n138 VTAIL.n137 9.3005
R467 VTAIL.n181 VTAIL.n180 9.3005
R468 VTAIL.n179 VTAIL.n178 9.3005
R469 VTAIL.n155 VTAIL.n154 9.3005
R470 VTAIL.n150 VTAIL.n149 9.3005
R471 VTAIL.n161 VTAIL.n160 9.3005
R472 VTAIL.n163 VTAIL.n162 9.3005
R473 VTAIL.n146 VTAIL.n145 9.3005
R474 VTAIL.n169 VTAIL.n168 9.3005
R475 VTAIL.n171 VTAIL.n170 9.3005
R476 VTAIL.n172 VTAIL.n141 9.3005
R477 VTAIL.n420 VTAIL.n419 9.3005
R478 VTAIL.n415 VTAIL.n414 9.3005
R479 VTAIL.n426 VTAIL.n425 9.3005
R480 VTAIL.n428 VTAIL.n427 9.3005
R481 VTAIL.n411 VTAIL.n410 9.3005
R482 VTAIL.n434 VTAIL.n433 9.3005
R483 VTAIL.n436 VTAIL.n435 9.3005
R484 VTAIL.n408 VTAIL.n405 9.3005
R485 VTAIL.n459 VTAIL.n458 9.3005
R486 VTAIL.n398 VTAIL.n397 9.3005
R487 VTAIL.n453 VTAIL.n452 9.3005
R488 VTAIL.n451 VTAIL.n450 9.3005
R489 VTAIL.n402 VTAIL.n401 9.3005
R490 VTAIL.n445 VTAIL.n444 9.3005
R491 VTAIL.n443 VTAIL.n442 9.3005
R492 VTAIL.n354 VTAIL.n353 9.3005
R493 VTAIL.n349 VTAIL.n348 9.3005
R494 VTAIL.n360 VTAIL.n359 9.3005
R495 VTAIL.n362 VTAIL.n361 9.3005
R496 VTAIL.n345 VTAIL.n344 9.3005
R497 VTAIL.n368 VTAIL.n367 9.3005
R498 VTAIL.n370 VTAIL.n369 9.3005
R499 VTAIL.n342 VTAIL.n339 9.3005
R500 VTAIL.n393 VTAIL.n392 9.3005
R501 VTAIL.n332 VTAIL.n331 9.3005
R502 VTAIL.n387 VTAIL.n386 9.3005
R503 VTAIL.n385 VTAIL.n384 9.3005
R504 VTAIL.n336 VTAIL.n335 9.3005
R505 VTAIL.n379 VTAIL.n378 9.3005
R506 VTAIL.n377 VTAIL.n376 9.3005
R507 VTAIL.n288 VTAIL.n287 9.3005
R508 VTAIL.n283 VTAIL.n282 9.3005
R509 VTAIL.n294 VTAIL.n293 9.3005
R510 VTAIL.n296 VTAIL.n295 9.3005
R511 VTAIL.n279 VTAIL.n278 9.3005
R512 VTAIL.n302 VTAIL.n301 9.3005
R513 VTAIL.n304 VTAIL.n303 9.3005
R514 VTAIL.n276 VTAIL.n273 9.3005
R515 VTAIL.n327 VTAIL.n326 9.3005
R516 VTAIL.n266 VTAIL.n265 9.3005
R517 VTAIL.n321 VTAIL.n320 9.3005
R518 VTAIL.n319 VTAIL.n318 9.3005
R519 VTAIL.n270 VTAIL.n269 9.3005
R520 VTAIL.n313 VTAIL.n312 9.3005
R521 VTAIL.n311 VTAIL.n310 9.3005
R522 VTAIL.n222 VTAIL.n221 9.3005
R523 VTAIL.n217 VTAIL.n216 9.3005
R524 VTAIL.n228 VTAIL.n227 9.3005
R525 VTAIL.n230 VTAIL.n229 9.3005
R526 VTAIL.n213 VTAIL.n212 9.3005
R527 VTAIL.n236 VTAIL.n235 9.3005
R528 VTAIL.n238 VTAIL.n237 9.3005
R529 VTAIL.n210 VTAIL.n207 9.3005
R530 VTAIL.n261 VTAIL.n260 9.3005
R531 VTAIL.n200 VTAIL.n199 9.3005
R532 VTAIL.n255 VTAIL.n254 9.3005
R533 VTAIL.n253 VTAIL.n252 9.3005
R534 VTAIL.n204 VTAIL.n203 9.3005
R535 VTAIL.n247 VTAIL.n246 9.3005
R536 VTAIL.n245 VTAIL.n244 9.3005
R537 VTAIL.n490 VTAIL.n489 8.92171
R538 VTAIL.n523 VTAIL.n464 8.92171
R539 VTAIL.n28 VTAIL.n27 8.92171
R540 VTAIL.n61 VTAIL.n2 8.92171
R541 VTAIL.n94 VTAIL.n93 8.92171
R542 VTAIL.n127 VTAIL.n68 8.92171
R543 VTAIL.n160 VTAIL.n159 8.92171
R544 VTAIL.n193 VTAIL.n134 8.92171
R545 VTAIL.n457 VTAIL.n398 8.92171
R546 VTAIL.n425 VTAIL.n424 8.92171
R547 VTAIL.n391 VTAIL.n332 8.92171
R548 VTAIL.n359 VTAIL.n358 8.92171
R549 VTAIL.n325 VTAIL.n266 8.92171
R550 VTAIL.n293 VTAIL.n292 8.92171
R551 VTAIL.n259 VTAIL.n200 8.92171
R552 VTAIL.n227 VTAIL.n226 8.92171
R553 VTAIL.n486 VTAIL.n480 8.14595
R554 VTAIL.n524 VTAIL.n462 8.14595
R555 VTAIL.n24 VTAIL.n18 8.14595
R556 VTAIL.n62 VTAIL.n0 8.14595
R557 VTAIL.n90 VTAIL.n84 8.14595
R558 VTAIL.n128 VTAIL.n66 8.14595
R559 VTAIL.n156 VTAIL.n150 8.14595
R560 VTAIL.n194 VTAIL.n132 8.14595
R561 VTAIL.n458 VTAIL.n396 8.14595
R562 VTAIL.n421 VTAIL.n415 8.14595
R563 VTAIL.n392 VTAIL.n330 8.14595
R564 VTAIL.n355 VTAIL.n349 8.14595
R565 VTAIL.n326 VTAIL.n264 8.14595
R566 VTAIL.n289 VTAIL.n283 8.14595
R567 VTAIL.n260 VTAIL.n198 8.14595
R568 VTAIL.n223 VTAIL.n217 8.14595
R569 VTAIL.n485 VTAIL.n482 7.3702
R570 VTAIL.n23 VTAIL.n20 7.3702
R571 VTAIL.n89 VTAIL.n86 7.3702
R572 VTAIL.n155 VTAIL.n152 7.3702
R573 VTAIL.n420 VTAIL.n417 7.3702
R574 VTAIL.n354 VTAIL.n351 7.3702
R575 VTAIL.n288 VTAIL.n285 7.3702
R576 VTAIL.n222 VTAIL.n219 7.3702
R577 VTAIL.n486 VTAIL.n485 5.81868
R578 VTAIL.n526 VTAIL.n462 5.81868
R579 VTAIL.n24 VTAIL.n23 5.81868
R580 VTAIL.n64 VTAIL.n0 5.81868
R581 VTAIL.n90 VTAIL.n89 5.81868
R582 VTAIL.n130 VTAIL.n66 5.81868
R583 VTAIL.n156 VTAIL.n155 5.81868
R584 VTAIL.n196 VTAIL.n132 5.81868
R585 VTAIL.n460 VTAIL.n396 5.81868
R586 VTAIL.n421 VTAIL.n420 5.81868
R587 VTAIL.n394 VTAIL.n330 5.81868
R588 VTAIL.n355 VTAIL.n354 5.81868
R589 VTAIL.n328 VTAIL.n264 5.81868
R590 VTAIL.n289 VTAIL.n288 5.81868
R591 VTAIL.n262 VTAIL.n198 5.81868
R592 VTAIL.n223 VTAIL.n222 5.81868
R593 VTAIL.n489 VTAIL.n480 5.04292
R594 VTAIL.n524 VTAIL.n523 5.04292
R595 VTAIL.n27 VTAIL.n18 5.04292
R596 VTAIL.n62 VTAIL.n61 5.04292
R597 VTAIL.n93 VTAIL.n84 5.04292
R598 VTAIL.n128 VTAIL.n127 5.04292
R599 VTAIL.n159 VTAIL.n150 5.04292
R600 VTAIL.n194 VTAIL.n193 5.04292
R601 VTAIL.n458 VTAIL.n457 5.04292
R602 VTAIL.n424 VTAIL.n415 5.04292
R603 VTAIL.n392 VTAIL.n391 5.04292
R604 VTAIL.n358 VTAIL.n349 5.04292
R605 VTAIL.n326 VTAIL.n325 5.04292
R606 VTAIL.n292 VTAIL.n283 5.04292
R607 VTAIL.n260 VTAIL.n259 5.04292
R608 VTAIL.n226 VTAIL.n217 5.04292
R609 VTAIL.n490 VTAIL.n478 4.26717
R610 VTAIL.n520 VTAIL.n464 4.26717
R611 VTAIL.n28 VTAIL.n16 4.26717
R612 VTAIL.n58 VTAIL.n2 4.26717
R613 VTAIL.n94 VTAIL.n82 4.26717
R614 VTAIL.n124 VTAIL.n68 4.26717
R615 VTAIL.n160 VTAIL.n148 4.26717
R616 VTAIL.n190 VTAIL.n134 4.26717
R617 VTAIL.n454 VTAIL.n398 4.26717
R618 VTAIL.n425 VTAIL.n413 4.26717
R619 VTAIL.n388 VTAIL.n332 4.26717
R620 VTAIL.n359 VTAIL.n347 4.26717
R621 VTAIL.n322 VTAIL.n266 4.26717
R622 VTAIL.n293 VTAIL.n281 4.26717
R623 VTAIL.n256 VTAIL.n200 4.26717
R624 VTAIL.n227 VTAIL.n215 4.26717
R625 VTAIL.n494 VTAIL.n493 3.49141
R626 VTAIL.n519 VTAIL.n466 3.49141
R627 VTAIL.n32 VTAIL.n31 3.49141
R628 VTAIL.n57 VTAIL.n4 3.49141
R629 VTAIL.n98 VTAIL.n97 3.49141
R630 VTAIL.n123 VTAIL.n70 3.49141
R631 VTAIL.n164 VTAIL.n163 3.49141
R632 VTAIL.n189 VTAIL.n136 3.49141
R633 VTAIL.n453 VTAIL.n400 3.49141
R634 VTAIL.n429 VTAIL.n428 3.49141
R635 VTAIL.n387 VTAIL.n334 3.49141
R636 VTAIL.n363 VTAIL.n362 3.49141
R637 VTAIL.n321 VTAIL.n268 3.49141
R638 VTAIL.n297 VTAIL.n296 3.49141
R639 VTAIL.n255 VTAIL.n202 3.49141
R640 VTAIL.n231 VTAIL.n230 3.49141
R641 VTAIL.n497 VTAIL.n476 2.71565
R642 VTAIL.n516 VTAIL.n515 2.71565
R643 VTAIL.n35 VTAIL.n14 2.71565
R644 VTAIL.n54 VTAIL.n53 2.71565
R645 VTAIL.n101 VTAIL.n80 2.71565
R646 VTAIL.n120 VTAIL.n119 2.71565
R647 VTAIL.n167 VTAIL.n146 2.71565
R648 VTAIL.n186 VTAIL.n185 2.71565
R649 VTAIL.n450 VTAIL.n449 2.71565
R650 VTAIL.n432 VTAIL.n411 2.71565
R651 VTAIL.n384 VTAIL.n383 2.71565
R652 VTAIL.n366 VTAIL.n345 2.71565
R653 VTAIL.n318 VTAIL.n317 2.71565
R654 VTAIL.n300 VTAIL.n279 2.71565
R655 VTAIL.n252 VTAIL.n251 2.71565
R656 VTAIL.n234 VTAIL.n213 2.71565
R657 VTAIL.n419 VTAIL.n418 2.41282
R658 VTAIL.n353 VTAIL.n352 2.41282
R659 VTAIL.n287 VTAIL.n286 2.41282
R660 VTAIL.n221 VTAIL.n220 2.41282
R661 VTAIL.n484 VTAIL.n483 2.41282
R662 VTAIL.n22 VTAIL.n21 2.41282
R663 VTAIL.n88 VTAIL.n87 2.41282
R664 VTAIL.n154 VTAIL.n153 2.41282
R665 VTAIL.n329 VTAIL.n263 2.16429
R666 VTAIL.n461 VTAIL.n395 2.16429
R667 VTAIL.n197 VTAIL.n131 2.16429
R668 VTAIL.n498 VTAIL.n474 1.93989
R669 VTAIL.n512 VTAIL.n468 1.93989
R670 VTAIL.n36 VTAIL.n12 1.93989
R671 VTAIL.n50 VTAIL.n6 1.93989
R672 VTAIL.n102 VTAIL.n78 1.93989
R673 VTAIL.n116 VTAIL.n72 1.93989
R674 VTAIL.n168 VTAIL.n144 1.93989
R675 VTAIL.n182 VTAIL.n138 1.93989
R676 VTAIL.n446 VTAIL.n402 1.93989
R677 VTAIL.n433 VTAIL.n409 1.93989
R678 VTAIL.n380 VTAIL.n336 1.93989
R679 VTAIL.n367 VTAIL.n343 1.93989
R680 VTAIL.n314 VTAIL.n270 1.93989
R681 VTAIL.n301 VTAIL.n277 1.93989
R682 VTAIL.n248 VTAIL.n204 1.93989
R683 VTAIL.n235 VTAIL.n211 1.93989
R684 VTAIL.n503 VTAIL.n501 1.16414
R685 VTAIL.n511 VTAIL.n470 1.16414
R686 VTAIL.n41 VTAIL.n39 1.16414
R687 VTAIL.n49 VTAIL.n8 1.16414
R688 VTAIL.n107 VTAIL.n105 1.16414
R689 VTAIL.n115 VTAIL.n74 1.16414
R690 VTAIL.n173 VTAIL.n171 1.16414
R691 VTAIL.n181 VTAIL.n140 1.16414
R692 VTAIL.n445 VTAIL.n404 1.16414
R693 VTAIL.n437 VTAIL.n436 1.16414
R694 VTAIL.n379 VTAIL.n338 1.16414
R695 VTAIL.n371 VTAIL.n370 1.16414
R696 VTAIL.n313 VTAIL.n272 1.16414
R697 VTAIL.n305 VTAIL.n304 1.16414
R698 VTAIL.n247 VTAIL.n206 1.16414
R699 VTAIL.n239 VTAIL.n238 1.16414
R700 VTAIL VTAIL.n65 1.14059
R701 VTAIL VTAIL.n527 1.02421
R702 VTAIL.n395 VTAIL.n329 0.470328
R703 VTAIL.n131 VTAIL.n65 0.470328
R704 VTAIL.n502 VTAIL.n472 0.388379
R705 VTAIL.n508 VTAIL.n507 0.388379
R706 VTAIL.n40 VTAIL.n10 0.388379
R707 VTAIL.n46 VTAIL.n45 0.388379
R708 VTAIL.n106 VTAIL.n76 0.388379
R709 VTAIL.n112 VTAIL.n111 0.388379
R710 VTAIL.n172 VTAIL.n142 0.388379
R711 VTAIL.n178 VTAIL.n177 0.388379
R712 VTAIL.n442 VTAIL.n441 0.388379
R713 VTAIL.n408 VTAIL.n406 0.388379
R714 VTAIL.n376 VTAIL.n375 0.388379
R715 VTAIL.n342 VTAIL.n340 0.388379
R716 VTAIL.n310 VTAIL.n309 0.388379
R717 VTAIL.n276 VTAIL.n274 0.388379
R718 VTAIL.n244 VTAIL.n243 0.388379
R719 VTAIL.n210 VTAIL.n208 0.388379
R720 VTAIL.n484 VTAIL.n479 0.155672
R721 VTAIL.n491 VTAIL.n479 0.155672
R722 VTAIL.n492 VTAIL.n491 0.155672
R723 VTAIL.n492 VTAIL.n475 0.155672
R724 VTAIL.n499 VTAIL.n475 0.155672
R725 VTAIL.n500 VTAIL.n499 0.155672
R726 VTAIL.n500 VTAIL.n471 0.155672
R727 VTAIL.n509 VTAIL.n471 0.155672
R728 VTAIL.n510 VTAIL.n509 0.155672
R729 VTAIL.n510 VTAIL.n467 0.155672
R730 VTAIL.n517 VTAIL.n467 0.155672
R731 VTAIL.n518 VTAIL.n517 0.155672
R732 VTAIL.n518 VTAIL.n463 0.155672
R733 VTAIL.n525 VTAIL.n463 0.155672
R734 VTAIL.n22 VTAIL.n17 0.155672
R735 VTAIL.n29 VTAIL.n17 0.155672
R736 VTAIL.n30 VTAIL.n29 0.155672
R737 VTAIL.n30 VTAIL.n13 0.155672
R738 VTAIL.n37 VTAIL.n13 0.155672
R739 VTAIL.n38 VTAIL.n37 0.155672
R740 VTAIL.n38 VTAIL.n9 0.155672
R741 VTAIL.n47 VTAIL.n9 0.155672
R742 VTAIL.n48 VTAIL.n47 0.155672
R743 VTAIL.n48 VTAIL.n5 0.155672
R744 VTAIL.n55 VTAIL.n5 0.155672
R745 VTAIL.n56 VTAIL.n55 0.155672
R746 VTAIL.n56 VTAIL.n1 0.155672
R747 VTAIL.n63 VTAIL.n1 0.155672
R748 VTAIL.n88 VTAIL.n83 0.155672
R749 VTAIL.n95 VTAIL.n83 0.155672
R750 VTAIL.n96 VTAIL.n95 0.155672
R751 VTAIL.n96 VTAIL.n79 0.155672
R752 VTAIL.n103 VTAIL.n79 0.155672
R753 VTAIL.n104 VTAIL.n103 0.155672
R754 VTAIL.n104 VTAIL.n75 0.155672
R755 VTAIL.n113 VTAIL.n75 0.155672
R756 VTAIL.n114 VTAIL.n113 0.155672
R757 VTAIL.n114 VTAIL.n71 0.155672
R758 VTAIL.n121 VTAIL.n71 0.155672
R759 VTAIL.n122 VTAIL.n121 0.155672
R760 VTAIL.n122 VTAIL.n67 0.155672
R761 VTAIL.n129 VTAIL.n67 0.155672
R762 VTAIL.n154 VTAIL.n149 0.155672
R763 VTAIL.n161 VTAIL.n149 0.155672
R764 VTAIL.n162 VTAIL.n161 0.155672
R765 VTAIL.n162 VTAIL.n145 0.155672
R766 VTAIL.n169 VTAIL.n145 0.155672
R767 VTAIL.n170 VTAIL.n169 0.155672
R768 VTAIL.n170 VTAIL.n141 0.155672
R769 VTAIL.n179 VTAIL.n141 0.155672
R770 VTAIL.n180 VTAIL.n179 0.155672
R771 VTAIL.n180 VTAIL.n137 0.155672
R772 VTAIL.n187 VTAIL.n137 0.155672
R773 VTAIL.n188 VTAIL.n187 0.155672
R774 VTAIL.n188 VTAIL.n133 0.155672
R775 VTAIL.n195 VTAIL.n133 0.155672
R776 VTAIL.n459 VTAIL.n397 0.155672
R777 VTAIL.n452 VTAIL.n397 0.155672
R778 VTAIL.n452 VTAIL.n451 0.155672
R779 VTAIL.n451 VTAIL.n401 0.155672
R780 VTAIL.n444 VTAIL.n401 0.155672
R781 VTAIL.n444 VTAIL.n443 0.155672
R782 VTAIL.n443 VTAIL.n405 0.155672
R783 VTAIL.n435 VTAIL.n405 0.155672
R784 VTAIL.n435 VTAIL.n434 0.155672
R785 VTAIL.n434 VTAIL.n410 0.155672
R786 VTAIL.n427 VTAIL.n410 0.155672
R787 VTAIL.n427 VTAIL.n426 0.155672
R788 VTAIL.n426 VTAIL.n414 0.155672
R789 VTAIL.n419 VTAIL.n414 0.155672
R790 VTAIL.n393 VTAIL.n331 0.155672
R791 VTAIL.n386 VTAIL.n331 0.155672
R792 VTAIL.n386 VTAIL.n385 0.155672
R793 VTAIL.n385 VTAIL.n335 0.155672
R794 VTAIL.n378 VTAIL.n335 0.155672
R795 VTAIL.n378 VTAIL.n377 0.155672
R796 VTAIL.n377 VTAIL.n339 0.155672
R797 VTAIL.n369 VTAIL.n339 0.155672
R798 VTAIL.n369 VTAIL.n368 0.155672
R799 VTAIL.n368 VTAIL.n344 0.155672
R800 VTAIL.n361 VTAIL.n344 0.155672
R801 VTAIL.n361 VTAIL.n360 0.155672
R802 VTAIL.n360 VTAIL.n348 0.155672
R803 VTAIL.n353 VTAIL.n348 0.155672
R804 VTAIL.n327 VTAIL.n265 0.155672
R805 VTAIL.n320 VTAIL.n265 0.155672
R806 VTAIL.n320 VTAIL.n319 0.155672
R807 VTAIL.n319 VTAIL.n269 0.155672
R808 VTAIL.n312 VTAIL.n269 0.155672
R809 VTAIL.n312 VTAIL.n311 0.155672
R810 VTAIL.n311 VTAIL.n273 0.155672
R811 VTAIL.n303 VTAIL.n273 0.155672
R812 VTAIL.n303 VTAIL.n302 0.155672
R813 VTAIL.n302 VTAIL.n278 0.155672
R814 VTAIL.n295 VTAIL.n278 0.155672
R815 VTAIL.n295 VTAIL.n294 0.155672
R816 VTAIL.n294 VTAIL.n282 0.155672
R817 VTAIL.n287 VTAIL.n282 0.155672
R818 VTAIL.n261 VTAIL.n199 0.155672
R819 VTAIL.n254 VTAIL.n199 0.155672
R820 VTAIL.n254 VTAIL.n253 0.155672
R821 VTAIL.n253 VTAIL.n203 0.155672
R822 VTAIL.n246 VTAIL.n203 0.155672
R823 VTAIL.n246 VTAIL.n245 0.155672
R824 VTAIL.n245 VTAIL.n207 0.155672
R825 VTAIL.n237 VTAIL.n207 0.155672
R826 VTAIL.n237 VTAIL.n236 0.155672
R827 VTAIL.n236 VTAIL.n212 0.155672
R828 VTAIL.n229 VTAIL.n212 0.155672
R829 VTAIL.n229 VTAIL.n228 0.155672
R830 VTAIL.n228 VTAIL.n216 0.155672
R831 VTAIL.n221 VTAIL.n216 0.155672
R832 VN.n0 VN.t3 170.489
R833 VN.n1 VN.t1 170.489
R834 VN.n0 VN.t2 169.856
R835 VN.n1 VN.t0 169.856
R836 VN VN.n1 51.2409
R837 VN VN.n0 5.88109
R838 VDD2.n2 VDD2.n0 116.114
R839 VDD2.n2 VDD2.n1 75.3905
R840 VDD2.n1 VDD2.t3 2.66484
R841 VDD2.n1 VDD2.t2 2.66484
R842 VDD2.n0 VDD2.t0 2.66484
R843 VDD2.n0 VDD2.t1 2.66484
R844 VDD2 VDD2.n2 0.0586897
R845 B.n443 B.n68 585
R846 B.n445 B.n444 585
R847 B.n446 B.n67 585
R848 B.n448 B.n447 585
R849 B.n449 B.n66 585
R850 B.n451 B.n450 585
R851 B.n452 B.n65 585
R852 B.n454 B.n453 585
R853 B.n455 B.n64 585
R854 B.n457 B.n456 585
R855 B.n458 B.n63 585
R856 B.n460 B.n459 585
R857 B.n461 B.n62 585
R858 B.n463 B.n462 585
R859 B.n464 B.n61 585
R860 B.n466 B.n465 585
R861 B.n467 B.n60 585
R862 B.n469 B.n468 585
R863 B.n470 B.n59 585
R864 B.n472 B.n471 585
R865 B.n473 B.n58 585
R866 B.n475 B.n474 585
R867 B.n476 B.n57 585
R868 B.n478 B.n477 585
R869 B.n479 B.n56 585
R870 B.n481 B.n480 585
R871 B.n482 B.n55 585
R872 B.n484 B.n483 585
R873 B.n485 B.n54 585
R874 B.n487 B.n486 585
R875 B.n488 B.n53 585
R876 B.n490 B.n489 585
R877 B.n491 B.n52 585
R878 B.n493 B.n492 585
R879 B.n494 B.n51 585
R880 B.n496 B.n495 585
R881 B.n497 B.n50 585
R882 B.n499 B.n498 585
R883 B.n500 B.n49 585
R884 B.n502 B.n501 585
R885 B.n503 B.n48 585
R886 B.n505 B.n504 585
R887 B.n507 B.n45 585
R888 B.n509 B.n508 585
R889 B.n510 B.n44 585
R890 B.n512 B.n511 585
R891 B.n513 B.n43 585
R892 B.n515 B.n514 585
R893 B.n516 B.n42 585
R894 B.n518 B.n517 585
R895 B.n519 B.n41 585
R896 B.n521 B.n520 585
R897 B.n523 B.n522 585
R898 B.n524 B.n37 585
R899 B.n526 B.n525 585
R900 B.n527 B.n36 585
R901 B.n529 B.n528 585
R902 B.n530 B.n35 585
R903 B.n532 B.n531 585
R904 B.n533 B.n34 585
R905 B.n535 B.n534 585
R906 B.n536 B.n33 585
R907 B.n538 B.n537 585
R908 B.n539 B.n32 585
R909 B.n541 B.n540 585
R910 B.n542 B.n31 585
R911 B.n544 B.n543 585
R912 B.n545 B.n30 585
R913 B.n547 B.n546 585
R914 B.n548 B.n29 585
R915 B.n550 B.n549 585
R916 B.n551 B.n28 585
R917 B.n553 B.n552 585
R918 B.n554 B.n27 585
R919 B.n556 B.n555 585
R920 B.n557 B.n26 585
R921 B.n559 B.n558 585
R922 B.n560 B.n25 585
R923 B.n562 B.n561 585
R924 B.n563 B.n24 585
R925 B.n565 B.n564 585
R926 B.n566 B.n23 585
R927 B.n568 B.n567 585
R928 B.n569 B.n22 585
R929 B.n571 B.n570 585
R930 B.n572 B.n21 585
R931 B.n574 B.n573 585
R932 B.n575 B.n20 585
R933 B.n577 B.n576 585
R934 B.n578 B.n19 585
R935 B.n580 B.n579 585
R936 B.n581 B.n18 585
R937 B.n583 B.n582 585
R938 B.n584 B.n17 585
R939 B.n442 B.n441 585
R940 B.n440 B.n69 585
R941 B.n439 B.n438 585
R942 B.n437 B.n70 585
R943 B.n436 B.n435 585
R944 B.n434 B.n71 585
R945 B.n433 B.n432 585
R946 B.n431 B.n72 585
R947 B.n430 B.n429 585
R948 B.n428 B.n73 585
R949 B.n427 B.n426 585
R950 B.n425 B.n74 585
R951 B.n424 B.n423 585
R952 B.n422 B.n75 585
R953 B.n421 B.n420 585
R954 B.n419 B.n76 585
R955 B.n418 B.n417 585
R956 B.n416 B.n77 585
R957 B.n415 B.n414 585
R958 B.n413 B.n78 585
R959 B.n412 B.n411 585
R960 B.n410 B.n79 585
R961 B.n409 B.n408 585
R962 B.n407 B.n80 585
R963 B.n406 B.n405 585
R964 B.n404 B.n81 585
R965 B.n403 B.n402 585
R966 B.n401 B.n82 585
R967 B.n400 B.n399 585
R968 B.n398 B.n83 585
R969 B.n397 B.n396 585
R970 B.n395 B.n84 585
R971 B.n394 B.n393 585
R972 B.n392 B.n85 585
R973 B.n391 B.n390 585
R974 B.n389 B.n86 585
R975 B.n388 B.n387 585
R976 B.n386 B.n87 585
R977 B.n385 B.n384 585
R978 B.n383 B.n88 585
R979 B.n382 B.n381 585
R980 B.n380 B.n89 585
R981 B.n379 B.n378 585
R982 B.n377 B.n90 585
R983 B.n376 B.n375 585
R984 B.n374 B.n91 585
R985 B.n373 B.n372 585
R986 B.n371 B.n92 585
R987 B.n370 B.n369 585
R988 B.n368 B.n93 585
R989 B.n367 B.n366 585
R990 B.n365 B.n94 585
R991 B.n364 B.n363 585
R992 B.n362 B.n95 585
R993 B.n361 B.n360 585
R994 B.n359 B.n96 585
R995 B.n358 B.n357 585
R996 B.n356 B.n97 585
R997 B.n355 B.n354 585
R998 B.n353 B.n98 585
R999 B.n352 B.n351 585
R1000 B.n209 B.n150 585
R1001 B.n211 B.n210 585
R1002 B.n212 B.n149 585
R1003 B.n214 B.n213 585
R1004 B.n215 B.n148 585
R1005 B.n217 B.n216 585
R1006 B.n218 B.n147 585
R1007 B.n220 B.n219 585
R1008 B.n221 B.n146 585
R1009 B.n223 B.n222 585
R1010 B.n224 B.n145 585
R1011 B.n226 B.n225 585
R1012 B.n227 B.n144 585
R1013 B.n229 B.n228 585
R1014 B.n230 B.n143 585
R1015 B.n232 B.n231 585
R1016 B.n233 B.n142 585
R1017 B.n235 B.n234 585
R1018 B.n236 B.n141 585
R1019 B.n238 B.n237 585
R1020 B.n239 B.n140 585
R1021 B.n241 B.n240 585
R1022 B.n242 B.n139 585
R1023 B.n244 B.n243 585
R1024 B.n245 B.n138 585
R1025 B.n247 B.n246 585
R1026 B.n248 B.n137 585
R1027 B.n250 B.n249 585
R1028 B.n251 B.n136 585
R1029 B.n253 B.n252 585
R1030 B.n254 B.n135 585
R1031 B.n256 B.n255 585
R1032 B.n257 B.n134 585
R1033 B.n259 B.n258 585
R1034 B.n260 B.n133 585
R1035 B.n262 B.n261 585
R1036 B.n263 B.n132 585
R1037 B.n265 B.n264 585
R1038 B.n266 B.n131 585
R1039 B.n268 B.n267 585
R1040 B.n269 B.n130 585
R1041 B.n271 B.n270 585
R1042 B.n273 B.n127 585
R1043 B.n275 B.n274 585
R1044 B.n276 B.n126 585
R1045 B.n278 B.n277 585
R1046 B.n279 B.n125 585
R1047 B.n281 B.n280 585
R1048 B.n282 B.n124 585
R1049 B.n284 B.n283 585
R1050 B.n285 B.n123 585
R1051 B.n287 B.n286 585
R1052 B.n289 B.n288 585
R1053 B.n290 B.n119 585
R1054 B.n292 B.n291 585
R1055 B.n293 B.n118 585
R1056 B.n295 B.n294 585
R1057 B.n296 B.n117 585
R1058 B.n298 B.n297 585
R1059 B.n299 B.n116 585
R1060 B.n301 B.n300 585
R1061 B.n302 B.n115 585
R1062 B.n304 B.n303 585
R1063 B.n305 B.n114 585
R1064 B.n307 B.n306 585
R1065 B.n308 B.n113 585
R1066 B.n310 B.n309 585
R1067 B.n311 B.n112 585
R1068 B.n313 B.n312 585
R1069 B.n314 B.n111 585
R1070 B.n316 B.n315 585
R1071 B.n317 B.n110 585
R1072 B.n319 B.n318 585
R1073 B.n320 B.n109 585
R1074 B.n322 B.n321 585
R1075 B.n323 B.n108 585
R1076 B.n325 B.n324 585
R1077 B.n326 B.n107 585
R1078 B.n328 B.n327 585
R1079 B.n329 B.n106 585
R1080 B.n331 B.n330 585
R1081 B.n332 B.n105 585
R1082 B.n334 B.n333 585
R1083 B.n335 B.n104 585
R1084 B.n337 B.n336 585
R1085 B.n338 B.n103 585
R1086 B.n340 B.n339 585
R1087 B.n341 B.n102 585
R1088 B.n343 B.n342 585
R1089 B.n344 B.n101 585
R1090 B.n346 B.n345 585
R1091 B.n347 B.n100 585
R1092 B.n349 B.n348 585
R1093 B.n350 B.n99 585
R1094 B.n208 B.n207 585
R1095 B.n206 B.n151 585
R1096 B.n205 B.n204 585
R1097 B.n203 B.n152 585
R1098 B.n202 B.n201 585
R1099 B.n200 B.n153 585
R1100 B.n199 B.n198 585
R1101 B.n197 B.n154 585
R1102 B.n196 B.n195 585
R1103 B.n194 B.n155 585
R1104 B.n193 B.n192 585
R1105 B.n191 B.n156 585
R1106 B.n190 B.n189 585
R1107 B.n188 B.n157 585
R1108 B.n187 B.n186 585
R1109 B.n185 B.n158 585
R1110 B.n184 B.n183 585
R1111 B.n182 B.n159 585
R1112 B.n181 B.n180 585
R1113 B.n179 B.n160 585
R1114 B.n178 B.n177 585
R1115 B.n176 B.n161 585
R1116 B.n175 B.n174 585
R1117 B.n173 B.n162 585
R1118 B.n172 B.n171 585
R1119 B.n170 B.n163 585
R1120 B.n169 B.n168 585
R1121 B.n167 B.n164 585
R1122 B.n166 B.n165 585
R1123 B.n2 B.n0 585
R1124 B.n629 B.n1 585
R1125 B.n628 B.n627 585
R1126 B.n626 B.n3 585
R1127 B.n625 B.n624 585
R1128 B.n623 B.n4 585
R1129 B.n622 B.n621 585
R1130 B.n620 B.n5 585
R1131 B.n619 B.n618 585
R1132 B.n617 B.n6 585
R1133 B.n616 B.n615 585
R1134 B.n614 B.n7 585
R1135 B.n613 B.n612 585
R1136 B.n611 B.n8 585
R1137 B.n610 B.n609 585
R1138 B.n608 B.n9 585
R1139 B.n607 B.n606 585
R1140 B.n605 B.n10 585
R1141 B.n604 B.n603 585
R1142 B.n602 B.n11 585
R1143 B.n601 B.n600 585
R1144 B.n599 B.n12 585
R1145 B.n598 B.n597 585
R1146 B.n596 B.n13 585
R1147 B.n595 B.n594 585
R1148 B.n593 B.n14 585
R1149 B.n592 B.n591 585
R1150 B.n590 B.n15 585
R1151 B.n589 B.n588 585
R1152 B.n587 B.n16 585
R1153 B.n586 B.n585 585
R1154 B.n631 B.n630 585
R1155 B.n209 B.n208 540.549
R1156 B.n586 B.n17 540.549
R1157 B.n352 B.n99 540.549
R1158 B.n443 B.n442 540.549
R1159 B.n120 B.t2 428.087
R1160 B.n46 B.t10 428.087
R1161 B.n128 B.t5 428.087
R1162 B.n38 B.t7 428.087
R1163 B.n121 B.t1 379.409
R1164 B.n47 B.t11 379.409
R1165 B.n129 B.t4 379.409
R1166 B.n39 B.t8 379.409
R1167 B.n120 B.t0 342.183
R1168 B.n128 B.t3 342.183
R1169 B.n38 B.t6 342.183
R1170 B.n46 B.t9 342.183
R1171 B.n208 B.n151 163.367
R1172 B.n204 B.n151 163.367
R1173 B.n204 B.n203 163.367
R1174 B.n203 B.n202 163.367
R1175 B.n202 B.n153 163.367
R1176 B.n198 B.n153 163.367
R1177 B.n198 B.n197 163.367
R1178 B.n197 B.n196 163.367
R1179 B.n196 B.n155 163.367
R1180 B.n192 B.n155 163.367
R1181 B.n192 B.n191 163.367
R1182 B.n191 B.n190 163.367
R1183 B.n190 B.n157 163.367
R1184 B.n186 B.n157 163.367
R1185 B.n186 B.n185 163.367
R1186 B.n185 B.n184 163.367
R1187 B.n184 B.n159 163.367
R1188 B.n180 B.n159 163.367
R1189 B.n180 B.n179 163.367
R1190 B.n179 B.n178 163.367
R1191 B.n178 B.n161 163.367
R1192 B.n174 B.n161 163.367
R1193 B.n174 B.n173 163.367
R1194 B.n173 B.n172 163.367
R1195 B.n172 B.n163 163.367
R1196 B.n168 B.n163 163.367
R1197 B.n168 B.n167 163.367
R1198 B.n167 B.n166 163.367
R1199 B.n166 B.n2 163.367
R1200 B.n630 B.n2 163.367
R1201 B.n630 B.n629 163.367
R1202 B.n629 B.n628 163.367
R1203 B.n628 B.n3 163.367
R1204 B.n624 B.n3 163.367
R1205 B.n624 B.n623 163.367
R1206 B.n623 B.n622 163.367
R1207 B.n622 B.n5 163.367
R1208 B.n618 B.n5 163.367
R1209 B.n618 B.n617 163.367
R1210 B.n617 B.n616 163.367
R1211 B.n616 B.n7 163.367
R1212 B.n612 B.n7 163.367
R1213 B.n612 B.n611 163.367
R1214 B.n611 B.n610 163.367
R1215 B.n610 B.n9 163.367
R1216 B.n606 B.n9 163.367
R1217 B.n606 B.n605 163.367
R1218 B.n605 B.n604 163.367
R1219 B.n604 B.n11 163.367
R1220 B.n600 B.n11 163.367
R1221 B.n600 B.n599 163.367
R1222 B.n599 B.n598 163.367
R1223 B.n598 B.n13 163.367
R1224 B.n594 B.n13 163.367
R1225 B.n594 B.n593 163.367
R1226 B.n593 B.n592 163.367
R1227 B.n592 B.n15 163.367
R1228 B.n588 B.n15 163.367
R1229 B.n588 B.n587 163.367
R1230 B.n587 B.n586 163.367
R1231 B.n210 B.n209 163.367
R1232 B.n210 B.n149 163.367
R1233 B.n214 B.n149 163.367
R1234 B.n215 B.n214 163.367
R1235 B.n216 B.n215 163.367
R1236 B.n216 B.n147 163.367
R1237 B.n220 B.n147 163.367
R1238 B.n221 B.n220 163.367
R1239 B.n222 B.n221 163.367
R1240 B.n222 B.n145 163.367
R1241 B.n226 B.n145 163.367
R1242 B.n227 B.n226 163.367
R1243 B.n228 B.n227 163.367
R1244 B.n228 B.n143 163.367
R1245 B.n232 B.n143 163.367
R1246 B.n233 B.n232 163.367
R1247 B.n234 B.n233 163.367
R1248 B.n234 B.n141 163.367
R1249 B.n238 B.n141 163.367
R1250 B.n239 B.n238 163.367
R1251 B.n240 B.n239 163.367
R1252 B.n240 B.n139 163.367
R1253 B.n244 B.n139 163.367
R1254 B.n245 B.n244 163.367
R1255 B.n246 B.n245 163.367
R1256 B.n246 B.n137 163.367
R1257 B.n250 B.n137 163.367
R1258 B.n251 B.n250 163.367
R1259 B.n252 B.n251 163.367
R1260 B.n252 B.n135 163.367
R1261 B.n256 B.n135 163.367
R1262 B.n257 B.n256 163.367
R1263 B.n258 B.n257 163.367
R1264 B.n258 B.n133 163.367
R1265 B.n262 B.n133 163.367
R1266 B.n263 B.n262 163.367
R1267 B.n264 B.n263 163.367
R1268 B.n264 B.n131 163.367
R1269 B.n268 B.n131 163.367
R1270 B.n269 B.n268 163.367
R1271 B.n270 B.n269 163.367
R1272 B.n270 B.n127 163.367
R1273 B.n275 B.n127 163.367
R1274 B.n276 B.n275 163.367
R1275 B.n277 B.n276 163.367
R1276 B.n277 B.n125 163.367
R1277 B.n281 B.n125 163.367
R1278 B.n282 B.n281 163.367
R1279 B.n283 B.n282 163.367
R1280 B.n283 B.n123 163.367
R1281 B.n287 B.n123 163.367
R1282 B.n288 B.n287 163.367
R1283 B.n288 B.n119 163.367
R1284 B.n292 B.n119 163.367
R1285 B.n293 B.n292 163.367
R1286 B.n294 B.n293 163.367
R1287 B.n294 B.n117 163.367
R1288 B.n298 B.n117 163.367
R1289 B.n299 B.n298 163.367
R1290 B.n300 B.n299 163.367
R1291 B.n300 B.n115 163.367
R1292 B.n304 B.n115 163.367
R1293 B.n305 B.n304 163.367
R1294 B.n306 B.n305 163.367
R1295 B.n306 B.n113 163.367
R1296 B.n310 B.n113 163.367
R1297 B.n311 B.n310 163.367
R1298 B.n312 B.n311 163.367
R1299 B.n312 B.n111 163.367
R1300 B.n316 B.n111 163.367
R1301 B.n317 B.n316 163.367
R1302 B.n318 B.n317 163.367
R1303 B.n318 B.n109 163.367
R1304 B.n322 B.n109 163.367
R1305 B.n323 B.n322 163.367
R1306 B.n324 B.n323 163.367
R1307 B.n324 B.n107 163.367
R1308 B.n328 B.n107 163.367
R1309 B.n329 B.n328 163.367
R1310 B.n330 B.n329 163.367
R1311 B.n330 B.n105 163.367
R1312 B.n334 B.n105 163.367
R1313 B.n335 B.n334 163.367
R1314 B.n336 B.n335 163.367
R1315 B.n336 B.n103 163.367
R1316 B.n340 B.n103 163.367
R1317 B.n341 B.n340 163.367
R1318 B.n342 B.n341 163.367
R1319 B.n342 B.n101 163.367
R1320 B.n346 B.n101 163.367
R1321 B.n347 B.n346 163.367
R1322 B.n348 B.n347 163.367
R1323 B.n348 B.n99 163.367
R1324 B.n353 B.n352 163.367
R1325 B.n354 B.n353 163.367
R1326 B.n354 B.n97 163.367
R1327 B.n358 B.n97 163.367
R1328 B.n359 B.n358 163.367
R1329 B.n360 B.n359 163.367
R1330 B.n360 B.n95 163.367
R1331 B.n364 B.n95 163.367
R1332 B.n365 B.n364 163.367
R1333 B.n366 B.n365 163.367
R1334 B.n366 B.n93 163.367
R1335 B.n370 B.n93 163.367
R1336 B.n371 B.n370 163.367
R1337 B.n372 B.n371 163.367
R1338 B.n372 B.n91 163.367
R1339 B.n376 B.n91 163.367
R1340 B.n377 B.n376 163.367
R1341 B.n378 B.n377 163.367
R1342 B.n378 B.n89 163.367
R1343 B.n382 B.n89 163.367
R1344 B.n383 B.n382 163.367
R1345 B.n384 B.n383 163.367
R1346 B.n384 B.n87 163.367
R1347 B.n388 B.n87 163.367
R1348 B.n389 B.n388 163.367
R1349 B.n390 B.n389 163.367
R1350 B.n390 B.n85 163.367
R1351 B.n394 B.n85 163.367
R1352 B.n395 B.n394 163.367
R1353 B.n396 B.n395 163.367
R1354 B.n396 B.n83 163.367
R1355 B.n400 B.n83 163.367
R1356 B.n401 B.n400 163.367
R1357 B.n402 B.n401 163.367
R1358 B.n402 B.n81 163.367
R1359 B.n406 B.n81 163.367
R1360 B.n407 B.n406 163.367
R1361 B.n408 B.n407 163.367
R1362 B.n408 B.n79 163.367
R1363 B.n412 B.n79 163.367
R1364 B.n413 B.n412 163.367
R1365 B.n414 B.n413 163.367
R1366 B.n414 B.n77 163.367
R1367 B.n418 B.n77 163.367
R1368 B.n419 B.n418 163.367
R1369 B.n420 B.n419 163.367
R1370 B.n420 B.n75 163.367
R1371 B.n424 B.n75 163.367
R1372 B.n425 B.n424 163.367
R1373 B.n426 B.n425 163.367
R1374 B.n426 B.n73 163.367
R1375 B.n430 B.n73 163.367
R1376 B.n431 B.n430 163.367
R1377 B.n432 B.n431 163.367
R1378 B.n432 B.n71 163.367
R1379 B.n436 B.n71 163.367
R1380 B.n437 B.n436 163.367
R1381 B.n438 B.n437 163.367
R1382 B.n438 B.n69 163.367
R1383 B.n442 B.n69 163.367
R1384 B.n582 B.n17 163.367
R1385 B.n582 B.n581 163.367
R1386 B.n581 B.n580 163.367
R1387 B.n580 B.n19 163.367
R1388 B.n576 B.n19 163.367
R1389 B.n576 B.n575 163.367
R1390 B.n575 B.n574 163.367
R1391 B.n574 B.n21 163.367
R1392 B.n570 B.n21 163.367
R1393 B.n570 B.n569 163.367
R1394 B.n569 B.n568 163.367
R1395 B.n568 B.n23 163.367
R1396 B.n564 B.n23 163.367
R1397 B.n564 B.n563 163.367
R1398 B.n563 B.n562 163.367
R1399 B.n562 B.n25 163.367
R1400 B.n558 B.n25 163.367
R1401 B.n558 B.n557 163.367
R1402 B.n557 B.n556 163.367
R1403 B.n556 B.n27 163.367
R1404 B.n552 B.n27 163.367
R1405 B.n552 B.n551 163.367
R1406 B.n551 B.n550 163.367
R1407 B.n550 B.n29 163.367
R1408 B.n546 B.n29 163.367
R1409 B.n546 B.n545 163.367
R1410 B.n545 B.n544 163.367
R1411 B.n544 B.n31 163.367
R1412 B.n540 B.n31 163.367
R1413 B.n540 B.n539 163.367
R1414 B.n539 B.n538 163.367
R1415 B.n538 B.n33 163.367
R1416 B.n534 B.n33 163.367
R1417 B.n534 B.n533 163.367
R1418 B.n533 B.n532 163.367
R1419 B.n532 B.n35 163.367
R1420 B.n528 B.n35 163.367
R1421 B.n528 B.n527 163.367
R1422 B.n527 B.n526 163.367
R1423 B.n526 B.n37 163.367
R1424 B.n522 B.n37 163.367
R1425 B.n522 B.n521 163.367
R1426 B.n521 B.n41 163.367
R1427 B.n517 B.n41 163.367
R1428 B.n517 B.n516 163.367
R1429 B.n516 B.n515 163.367
R1430 B.n515 B.n43 163.367
R1431 B.n511 B.n43 163.367
R1432 B.n511 B.n510 163.367
R1433 B.n510 B.n509 163.367
R1434 B.n509 B.n45 163.367
R1435 B.n504 B.n45 163.367
R1436 B.n504 B.n503 163.367
R1437 B.n503 B.n502 163.367
R1438 B.n502 B.n49 163.367
R1439 B.n498 B.n49 163.367
R1440 B.n498 B.n497 163.367
R1441 B.n497 B.n496 163.367
R1442 B.n496 B.n51 163.367
R1443 B.n492 B.n51 163.367
R1444 B.n492 B.n491 163.367
R1445 B.n491 B.n490 163.367
R1446 B.n490 B.n53 163.367
R1447 B.n486 B.n53 163.367
R1448 B.n486 B.n485 163.367
R1449 B.n485 B.n484 163.367
R1450 B.n484 B.n55 163.367
R1451 B.n480 B.n55 163.367
R1452 B.n480 B.n479 163.367
R1453 B.n479 B.n478 163.367
R1454 B.n478 B.n57 163.367
R1455 B.n474 B.n57 163.367
R1456 B.n474 B.n473 163.367
R1457 B.n473 B.n472 163.367
R1458 B.n472 B.n59 163.367
R1459 B.n468 B.n59 163.367
R1460 B.n468 B.n467 163.367
R1461 B.n467 B.n466 163.367
R1462 B.n466 B.n61 163.367
R1463 B.n462 B.n61 163.367
R1464 B.n462 B.n461 163.367
R1465 B.n461 B.n460 163.367
R1466 B.n460 B.n63 163.367
R1467 B.n456 B.n63 163.367
R1468 B.n456 B.n455 163.367
R1469 B.n455 B.n454 163.367
R1470 B.n454 B.n65 163.367
R1471 B.n450 B.n65 163.367
R1472 B.n450 B.n449 163.367
R1473 B.n449 B.n448 163.367
R1474 B.n448 B.n67 163.367
R1475 B.n444 B.n67 163.367
R1476 B.n444 B.n443 163.367
R1477 B.n122 B.n121 59.5399
R1478 B.n272 B.n129 59.5399
R1479 B.n40 B.n39 59.5399
R1480 B.n506 B.n47 59.5399
R1481 B.n121 B.n120 48.6793
R1482 B.n129 B.n128 48.6793
R1483 B.n39 B.n38 48.6793
R1484 B.n47 B.n46 48.6793
R1485 B.n585 B.n584 35.1225
R1486 B.n441 B.n68 35.1225
R1487 B.n351 B.n350 35.1225
R1488 B.n207 B.n150 35.1225
R1489 B B.n631 18.0485
R1490 B.n584 B.n583 10.6151
R1491 B.n583 B.n18 10.6151
R1492 B.n579 B.n18 10.6151
R1493 B.n579 B.n578 10.6151
R1494 B.n578 B.n577 10.6151
R1495 B.n577 B.n20 10.6151
R1496 B.n573 B.n20 10.6151
R1497 B.n573 B.n572 10.6151
R1498 B.n572 B.n571 10.6151
R1499 B.n571 B.n22 10.6151
R1500 B.n567 B.n22 10.6151
R1501 B.n567 B.n566 10.6151
R1502 B.n566 B.n565 10.6151
R1503 B.n565 B.n24 10.6151
R1504 B.n561 B.n24 10.6151
R1505 B.n561 B.n560 10.6151
R1506 B.n560 B.n559 10.6151
R1507 B.n559 B.n26 10.6151
R1508 B.n555 B.n26 10.6151
R1509 B.n555 B.n554 10.6151
R1510 B.n554 B.n553 10.6151
R1511 B.n553 B.n28 10.6151
R1512 B.n549 B.n28 10.6151
R1513 B.n549 B.n548 10.6151
R1514 B.n548 B.n547 10.6151
R1515 B.n547 B.n30 10.6151
R1516 B.n543 B.n30 10.6151
R1517 B.n543 B.n542 10.6151
R1518 B.n542 B.n541 10.6151
R1519 B.n541 B.n32 10.6151
R1520 B.n537 B.n32 10.6151
R1521 B.n537 B.n536 10.6151
R1522 B.n536 B.n535 10.6151
R1523 B.n535 B.n34 10.6151
R1524 B.n531 B.n34 10.6151
R1525 B.n531 B.n530 10.6151
R1526 B.n530 B.n529 10.6151
R1527 B.n529 B.n36 10.6151
R1528 B.n525 B.n36 10.6151
R1529 B.n525 B.n524 10.6151
R1530 B.n524 B.n523 10.6151
R1531 B.n520 B.n519 10.6151
R1532 B.n519 B.n518 10.6151
R1533 B.n518 B.n42 10.6151
R1534 B.n514 B.n42 10.6151
R1535 B.n514 B.n513 10.6151
R1536 B.n513 B.n512 10.6151
R1537 B.n512 B.n44 10.6151
R1538 B.n508 B.n44 10.6151
R1539 B.n508 B.n507 10.6151
R1540 B.n505 B.n48 10.6151
R1541 B.n501 B.n48 10.6151
R1542 B.n501 B.n500 10.6151
R1543 B.n500 B.n499 10.6151
R1544 B.n499 B.n50 10.6151
R1545 B.n495 B.n50 10.6151
R1546 B.n495 B.n494 10.6151
R1547 B.n494 B.n493 10.6151
R1548 B.n493 B.n52 10.6151
R1549 B.n489 B.n52 10.6151
R1550 B.n489 B.n488 10.6151
R1551 B.n488 B.n487 10.6151
R1552 B.n487 B.n54 10.6151
R1553 B.n483 B.n54 10.6151
R1554 B.n483 B.n482 10.6151
R1555 B.n482 B.n481 10.6151
R1556 B.n481 B.n56 10.6151
R1557 B.n477 B.n56 10.6151
R1558 B.n477 B.n476 10.6151
R1559 B.n476 B.n475 10.6151
R1560 B.n475 B.n58 10.6151
R1561 B.n471 B.n58 10.6151
R1562 B.n471 B.n470 10.6151
R1563 B.n470 B.n469 10.6151
R1564 B.n469 B.n60 10.6151
R1565 B.n465 B.n60 10.6151
R1566 B.n465 B.n464 10.6151
R1567 B.n464 B.n463 10.6151
R1568 B.n463 B.n62 10.6151
R1569 B.n459 B.n62 10.6151
R1570 B.n459 B.n458 10.6151
R1571 B.n458 B.n457 10.6151
R1572 B.n457 B.n64 10.6151
R1573 B.n453 B.n64 10.6151
R1574 B.n453 B.n452 10.6151
R1575 B.n452 B.n451 10.6151
R1576 B.n451 B.n66 10.6151
R1577 B.n447 B.n66 10.6151
R1578 B.n447 B.n446 10.6151
R1579 B.n446 B.n445 10.6151
R1580 B.n445 B.n68 10.6151
R1581 B.n351 B.n98 10.6151
R1582 B.n355 B.n98 10.6151
R1583 B.n356 B.n355 10.6151
R1584 B.n357 B.n356 10.6151
R1585 B.n357 B.n96 10.6151
R1586 B.n361 B.n96 10.6151
R1587 B.n362 B.n361 10.6151
R1588 B.n363 B.n362 10.6151
R1589 B.n363 B.n94 10.6151
R1590 B.n367 B.n94 10.6151
R1591 B.n368 B.n367 10.6151
R1592 B.n369 B.n368 10.6151
R1593 B.n369 B.n92 10.6151
R1594 B.n373 B.n92 10.6151
R1595 B.n374 B.n373 10.6151
R1596 B.n375 B.n374 10.6151
R1597 B.n375 B.n90 10.6151
R1598 B.n379 B.n90 10.6151
R1599 B.n380 B.n379 10.6151
R1600 B.n381 B.n380 10.6151
R1601 B.n381 B.n88 10.6151
R1602 B.n385 B.n88 10.6151
R1603 B.n386 B.n385 10.6151
R1604 B.n387 B.n386 10.6151
R1605 B.n387 B.n86 10.6151
R1606 B.n391 B.n86 10.6151
R1607 B.n392 B.n391 10.6151
R1608 B.n393 B.n392 10.6151
R1609 B.n393 B.n84 10.6151
R1610 B.n397 B.n84 10.6151
R1611 B.n398 B.n397 10.6151
R1612 B.n399 B.n398 10.6151
R1613 B.n399 B.n82 10.6151
R1614 B.n403 B.n82 10.6151
R1615 B.n404 B.n403 10.6151
R1616 B.n405 B.n404 10.6151
R1617 B.n405 B.n80 10.6151
R1618 B.n409 B.n80 10.6151
R1619 B.n410 B.n409 10.6151
R1620 B.n411 B.n410 10.6151
R1621 B.n411 B.n78 10.6151
R1622 B.n415 B.n78 10.6151
R1623 B.n416 B.n415 10.6151
R1624 B.n417 B.n416 10.6151
R1625 B.n417 B.n76 10.6151
R1626 B.n421 B.n76 10.6151
R1627 B.n422 B.n421 10.6151
R1628 B.n423 B.n422 10.6151
R1629 B.n423 B.n74 10.6151
R1630 B.n427 B.n74 10.6151
R1631 B.n428 B.n427 10.6151
R1632 B.n429 B.n428 10.6151
R1633 B.n429 B.n72 10.6151
R1634 B.n433 B.n72 10.6151
R1635 B.n434 B.n433 10.6151
R1636 B.n435 B.n434 10.6151
R1637 B.n435 B.n70 10.6151
R1638 B.n439 B.n70 10.6151
R1639 B.n440 B.n439 10.6151
R1640 B.n441 B.n440 10.6151
R1641 B.n211 B.n150 10.6151
R1642 B.n212 B.n211 10.6151
R1643 B.n213 B.n212 10.6151
R1644 B.n213 B.n148 10.6151
R1645 B.n217 B.n148 10.6151
R1646 B.n218 B.n217 10.6151
R1647 B.n219 B.n218 10.6151
R1648 B.n219 B.n146 10.6151
R1649 B.n223 B.n146 10.6151
R1650 B.n224 B.n223 10.6151
R1651 B.n225 B.n224 10.6151
R1652 B.n225 B.n144 10.6151
R1653 B.n229 B.n144 10.6151
R1654 B.n230 B.n229 10.6151
R1655 B.n231 B.n230 10.6151
R1656 B.n231 B.n142 10.6151
R1657 B.n235 B.n142 10.6151
R1658 B.n236 B.n235 10.6151
R1659 B.n237 B.n236 10.6151
R1660 B.n237 B.n140 10.6151
R1661 B.n241 B.n140 10.6151
R1662 B.n242 B.n241 10.6151
R1663 B.n243 B.n242 10.6151
R1664 B.n243 B.n138 10.6151
R1665 B.n247 B.n138 10.6151
R1666 B.n248 B.n247 10.6151
R1667 B.n249 B.n248 10.6151
R1668 B.n249 B.n136 10.6151
R1669 B.n253 B.n136 10.6151
R1670 B.n254 B.n253 10.6151
R1671 B.n255 B.n254 10.6151
R1672 B.n255 B.n134 10.6151
R1673 B.n259 B.n134 10.6151
R1674 B.n260 B.n259 10.6151
R1675 B.n261 B.n260 10.6151
R1676 B.n261 B.n132 10.6151
R1677 B.n265 B.n132 10.6151
R1678 B.n266 B.n265 10.6151
R1679 B.n267 B.n266 10.6151
R1680 B.n267 B.n130 10.6151
R1681 B.n271 B.n130 10.6151
R1682 B.n274 B.n273 10.6151
R1683 B.n274 B.n126 10.6151
R1684 B.n278 B.n126 10.6151
R1685 B.n279 B.n278 10.6151
R1686 B.n280 B.n279 10.6151
R1687 B.n280 B.n124 10.6151
R1688 B.n284 B.n124 10.6151
R1689 B.n285 B.n284 10.6151
R1690 B.n286 B.n285 10.6151
R1691 B.n290 B.n289 10.6151
R1692 B.n291 B.n290 10.6151
R1693 B.n291 B.n118 10.6151
R1694 B.n295 B.n118 10.6151
R1695 B.n296 B.n295 10.6151
R1696 B.n297 B.n296 10.6151
R1697 B.n297 B.n116 10.6151
R1698 B.n301 B.n116 10.6151
R1699 B.n302 B.n301 10.6151
R1700 B.n303 B.n302 10.6151
R1701 B.n303 B.n114 10.6151
R1702 B.n307 B.n114 10.6151
R1703 B.n308 B.n307 10.6151
R1704 B.n309 B.n308 10.6151
R1705 B.n309 B.n112 10.6151
R1706 B.n313 B.n112 10.6151
R1707 B.n314 B.n313 10.6151
R1708 B.n315 B.n314 10.6151
R1709 B.n315 B.n110 10.6151
R1710 B.n319 B.n110 10.6151
R1711 B.n320 B.n319 10.6151
R1712 B.n321 B.n320 10.6151
R1713 B.n321 B.n108 10.6151
R1714 B.n325 B.n108 10.6151
R1715 B.n326 B.n325 10.6151
R1716 B.n327 B.n326 10.6151
R1717 B.n327 B.n106 10.6151
R1718 B.n331 B.n106 10.6151
R1719 B.n332 B.n331 10.6151
R1720 B.n333 B.n332 10.6151
R1721 B.n333 B.n104 10.6151
R1722 B.n337 B.n104 10.6151
R1723 B.n338 B.n337 10.6151
R1724 B.n339 B.n338 10.6151
R1725 B.n339 B.n102 10.6151
R1726 B.n343 B.n102 10.6151
R1727 B.n344 B.n343 10.6151
R1728 B.n345 B.n344 10.6151
R1729 B.n345 B.n100 10.6151
R1730 B.n349 B.n100 10.6151
R1731 B.n350 B.n349 10.6151
R1732 B.n207 B.n206 10.6151
R1733 B.n206 B.n205 10.6151
R1734 B.n205 B.n152 10.6151
R1735 B.n201 B.n152 10.6151
R1736 B.n201 B.n200 10.6151
R1737 B.n200 B.n199 10.6151
R1738 B.n199 B.n154 10.6151
R1739 B.n195 B.n154 10.6151
R1740 B.n195 B.n194 10.6151
R1741 B.n194 B.n193 10.6151
R1742 B.n193 B.n156 10.6151
R1743 B.n189 B.n156 10.6151
R1744 B.n189 B.n188 10.6151
R1745 B.n188 B.n187 10.6151
R1746 B.n187 B.n158 10.6151
R1747 B.n183 B.n158 10.6151
R1748 B.n183 B.n182 10.6151
R1749 B.n182 B.n181 10.6151
R1750 B.n181 B.n160 10.6151
R1751 B.n177 B.n160 10.6151
R1752 B.n177 B.n176 10.6151
R1753 B.n176 B.n175 10.6151
R1754 B.n175 B.n162 10.6151
R1755 B.n171 B.n162 10.6151
R1756 B.n171 B.n170 10.6151
R1757 B.n170 B.n169 10.6151
R1758 B.n169 B.n164 10.6151
R1759 B.n165 B.n164 10.6151
R1760 B.n165 B.n0 10.6151
R1761 B.n627 B.n1 10.6151
R1762 B.n627 B.n626 10.6151
R1763 B.n626 B.n625 10.6151
R1764 B.n625 B.n4 10.6151
R1765 B.n621 B.n4 10.6151
R1766 B.n621 B.n620 10.6151
R1767 B.n620 B.n619 10.6151
R1768 B.n619 B.n6 10.6151
R1769 B.n615 B.n6 10.6151
R1770 B.n615 B.n614 10.6151
R1771 B.n614 B.n613 10.6151
R1772 B.n613 B.n8 10.6151
R1773 B.n609 B.n8 10.6151
R1774 B.n609 B.n608 10.6151
R1775 B.n608 B.n607 10.6151
R1776 B.n607 B.n10 10.6151
R1777 B.n603 B.n10 10.6151
R1778 B.n603 B.n602 10.6151
R1779 B.n602 B.n601 10.6151
R1780 B.n601 B.n12 10.6151
R1781 B.n597 B.n12 10.6151
R1782 B.n597 B.n596 10.6151
R1783 B.n596 B.n595 10.6151
R1784 B.n595 B.n14 10.6151
R1785 B.n591 B.n14 10.6151
R1786 B.n591 B.n590 10.6151
R1787 B.n590 B.n589 10.6151
R1788 B.n589 B.n16 10.6151
R1789 B.n585 B.n16 10.6151
R1790 B.n523 B.n40 9.36635
R1791 B.n506 B.n505 9.36635
R1792 B.n272 B.n271 9.36635
R1793 B.n289 B.n122 9.36635
R1794 B.n631 B.n0 2.81026
R1795 B.n631 B.n1 2.81026
R1796 B.n520 B.n40 1.24928
R1797 B.n507 B.n506 1.24928
R1798 B.n273 B.n272 1.24928
R1799 B.n286 B.n122 1.24928
C0 w_n2476_n3408# VDD1 1.37424f
C1 B VN 1.03478f
C2 B VTAIL 4.81166f
C3 w_n2476_n3408# VN 4.12686f
C4 w_n2476_n3408# VTAIL 4.01724f
C5 B VP 1.55926f
C6 w_n2476_n3408# VP 4.4441f
C7 VDD1 VDD2 0.926826f
C8 w_n2476_n3408# B 8.78556f
C9 VDD2 VN 4.6658f
C10 VTAIL VDD2 5.47458f
C11 VP VDD2 0.367742f
C12 VDD1 VN 0.148782f
C13 VTAIL VDD1 5.42318f
C14 VTAIL VN 4.50526f
C15 B VDD2 1.23954f
C16 VDD1 VP 4.88412f
C17 w_n2476_n3408# VDD2 1.42096f
C18 VP VN 5.92533f
C19 VTAIL VP 4.51936f
C20 B VDD1 1.19429f
C21 VDD2 VSUBS 0.878507f
C22 VDD1 VSUBS 5.51967f
C23 VTAIL VSUBS 1.171549f
C24 VN VSUBS 5.27352f
C25 VP VSUBS 2.071434f
C26 B VSUBS 3.925962f
C27 w_n2476_n3408# VSUBS 0.103843p
C28 B.n0 VSUBS 0.004388f
C29 B.n1 VSUBS 0.004388f
C30 B.n2 VSUBS 0.006939f
C31 B.n3 VSUBS 0.006939f
C32 B.n4 VSUBS 0.006939f
C33 B.n5 VSUBS 0.006939f
C34 B.n6 VSUBS 0.006939f
C35 B.n7 VSUBS 0.006939f
C36 B.n8 VSUBS 0.006939f
C37 B.n9 VSUBS 0.006939f
C38 B.n10 VSUBS 0.006939f
C39 B.n11 VSUBS 0.006939f
C40 B.n12 VSUBS 0.006939f
C41 B.n13 VSUBS 0.006939f
C42 B.n14 VSUBS 0.006939f
C43 B.n15 VSUBS 0.006939f
C44 B.n16 VSUBS 0.006939f
C45 B.n17 VSUBS 0.01757f
C46 B.n18 VSUBS 0.006939f
C47 B.n19 VSUBS 0.006939f
C48 B.n20 VSUBS 0.006939f
C49 B.n21 VSUBS 0.006939f
C50 B.n22 VSUBS 0.006939f
C51 B.n23 VSUBS 0.006939f
C52 B.n24 VSUBS 0.006939f
C53 B.n25 VSUBS 0.006939f
C54 B.n26 VSUBS 0.006939f
C55 B.n27 VSUBS 0.006939f
C56 B.n28 VSUBS 0.006939f
C57 B.n29 VSUBS 0.006939f
C58 B.n30 VSUBS 0.006939f
C59 B.n31 VSUBS 0.006939f
C60 B.n32 VSUBS 0.006939f
C61 B.n33 VSUBS 0.006939f
C62 B.n34 VSUBS 0.006939f
C63 B.n35 VSUBS 0.006939f
C64 B.n36 VSUBS 0.006939f
C65 B.n37 VSUBS 0.006939f
C66 B.t8 VSUBS 0.213792f
C67 B.t7 VSUBS 0.241146f
C68 B.t6 VSUBS 1.18477f
C69 B.n38 VSUBS 0.378251f
C70 B.n39 VSUBS 0.250444f
C71 B.n40 VSUBS 0.016076f
C72 B.n41 VSUBS 0.006939f
C73 B.n42 VSUBS 0.006939f
C74 B.n43 VSUBS 0.006939f
C75 B.n44 VSUBS 0.006939f
C76 B.n45 VSUBS 0.006939f
C77 B.t11 VSUBS 0.213795f
C78 B.t10 VSUBS 0.241148f
C79 B.t9 VSUBS 1.18477f
C80 B.n46 VSUBS 0.378248f
C81 B.n47 VSUBS 0.250441f
C82 B.n48 VSUBS 0.006939f
C83 B.n49 VSUBS 0.006939f
C84 B.n50 VSUBS 0.006939f
C85 B.n51 VSUBS 0.006939f
C86 B.n52 VSUBS 0.006939f
C87 B.n53 VSUBS 0.006939f
C88 B.n54 VSUBS 0.006939f
C89 B.n55 VSUBS 0.006939f
C90 B.n56 VSUBS 0.006939f
C91 B.n57 VSUBS 0.006939f
C92 B.n58 VSUBS 0.006939f
C93 B.n59 VSUBS 0.006939f
C94 B.n60 VSUBS 0.006939f
C95 B.n61 VSUBS 0.006939f
C96 B.n62 VSUBS 0.006939f
C97 B.n63 VSUBS 0.006939f
C98 B.n64 VSUBS 0.006939f
C99 B.n65 VSUBS 0.006939f
C100 B.n66 VSUBS 0.006939f
C101 B.n67 VSUBS 0.006939f
C102 B.n68 VSUBS 0.016808f
C103 B.n69 VSUBS 0.006939f
C104 B.n70 VSUBS 0.006939f
C105 B.n71 VSUBS 0.006939f
C106 B.n72 VSUBS 0.006939f
C107 B.n73 VSUBS 0.006939f
C108 B.n74 VSUBS 0.006939f
C109 B.n75 VSUBS 0.006939f
C110 B.n76 VSUBS 0.006939f
C111 B.n77 VSUBS 0.006939f
C112 B.n78 VSUBS 0.006939f
C113 B.n79 VSUBS 0.006939f
C114 B.n80 VSUBS 0.006939f
C115 B.n81 VSUBS 0.006939f
C116 B.n82 VSUBS 0.006939f
C117 B.n83 VSUBS 0.006939f
C118 B.n84 VSUBS 0.006939f
C119 B.n85 VSUBS 0.006939f
C120 B.n86 VSUBS 0.006939f
C121 B.n87 VSUBS 0.006939f
C122 B.n88 VSUBS 0.006939f
C123 B.n89 VSUBS 0.006939f
C124 B.n90 VSUBS 0.006939f
C125 B.n91 VSUBS 0.006939f
C126 B.n92 VSUBS 0.006939f
C127 B.n93 VSUBS 0.006939f
C128 B.n94 VSUBS 0.006939f
C129 B.n95 VSUBS 0.006939f
C130 B.n96 VSUBS 0.006939f
C131 B.n97 VSUBS 0.006939f
C132 B.n98 VSUBS 0.006939f
C133 B.n99 VSUBS 0.01757f
C134 B.n100 VSUBS 0.006939f
C135 B.n101 VSUBS 0.006939f
C136 B.n102 VSUBS 0.006939f
C137 B.n103 VSUBS 0.006939f
C138 B.n104 VSUBS 0.006939f
C139 B.n105 VSUBS 0.006939f
C140 B.n106 VSUBS 0.006939f
C141 B.n107 VSUBS 0.006939f
C142 B.n108 VSUBS 0.006939f
C143 B.n109 VSUBS 0.006939f
C144 B.n110 VSUBS 0.006939f
C145 B.n111 VSUBS 0.006939f
C146 B.n112 VSUBS 0.006939f
C147 B.n113 VSUBS 0.006939f
C148 B.n114 VSUBS 0.006939f
C149 B.n115 VSUBS 0.006939f
C150 B.n116 VSUBS 0.006939f
C151 B.n117 VSUBS 0.006939f
C152 B.n118 VSUBS 0.006939f
C153 B.n119 VSUBS 0.006939f
C154 B.t1 VSUBS 0.213795f
C155 B.t2 VSUBS 0.241148f
C156 B.t0 VSUBS 1.18477f
C157 B.n120 VSUBS 0.378248f
C158 B.n121 VSUBS 0.250441f
C159 B.n122 VSUBS 0.016076f
C160 B.n123 VSUBS 0.006939f
C161 B.n124 VSUBS 0.006939f
C162 B.n125 VSUBS 0.006939f
C163 B.n126 VSUBS 0.006939f
C164 B.n127 VSUBS 0.006939f
C165 B.t4 VSUBS 0.213792f
C166 B.t5 VSUBS 0.241146f
C167 B.t3 VSUBS 1.18477f
C168 B.n128 VSUBS 0.378251f
C169 B.n129 VSUBS 0.250444f
C170 B.n130 VSUBS 0.006939f
C171 B.n131 VSUBS 0.006939f
C172 B.n132 VSUBS 0.006939f
C173 B.n133 VSUBS 0.006939f
C174 B.n134 VSUBS 0.006939f
C175 B.n135 VSUBS 0.006939f
C176 B.n136 VSUBS 0.006939f
C177 B.n137 VSUBS 0.006939f
C178 B.n138 VSUBS 0.006939f
C179 B.n139 VSUBS 0.006939f
C180 B.n140 VSUBS 0.006939f
C181 B.n141 VSUBS 0.006939f
C182 B.n142 VSUBS 0.006939f
C183 B.n143 VSUBS 0.006939f
C184 B.n144 VSUBS 0.006939f
C185 B.n145 VSUBS 0.006939f
C186 B.n146 VSUBS 0.006939f
C187 B.n147 VSUBS 0.006939f
C188 B.n148 VSUBS 0.006939f
C189 B.n149 VSUBS 0.006939f
C190 B.n150 VSUBS 0.01757f
C191 B.n151 VSUBS 0.006939f
C192 B.n152 VSUBS 0.006939f
C193 B.n153 VSUBS 0.006939f
C194 B.n154 VSUBS 0.006939f
C195 B.n155 VSUBS 0.006939f
C196 B.n156 VSUBS 0.006939f
C197 B.n157 VSUBS 0.006939f
C198 B.n158 VSUBS 0.006939f
C199 B.n159 VSUBS 0.006939f
C200 B.n160 VSUBS 0.006939f
C201 B.n161 VSUBS 0.006939f
C202 B.n162 VSUBS 0.006939f
C203 B.n163 VSUBS 0.006939f
C204 B.n164 VSUBS 0.006939f
C205 B.n165 VSUBS 0.006939f
C206 B.n166 VSUBS 0.006939f
C207 B.n167 VSUBS 0.006939f
C208 B.n168 VSUBS 0.006939f
C209 B.n169 VSUBS 0.006939f
C210 B.n170 VSUBS 0.006939f
C211 B.n171 VSUBS 0.006939f
C212 B.n172 VSUBS 0.006939f
C213 B.n173 VSUBS 0.006939f
C214 B.n174 VSUBS 0.006939f
C215 B.n175 VSUBS 0.006939f
C216 B.n176 VSUBS 0.006939f
C217 B.n177 VSUBS 0.006939f
C218 B.n178 VSUBS 0.006939f
C219 B.n179 VSUBS 0.006939f
C220 B.n180 VSUBS 0.006939f
C221 B.n181 VSUBS 0.006939f
C222 B.n182 VSUBS 0.006939f
C223 B.n183 VSUBS 0.006939f
C224 B.n184 VSUBS 0.006939f
C225 B.n185 VSUBS 0.006939f
C226 B.n186 VSUBS 0.006939f
C227 B.n187 VSUBS 0.006939f
C228 B.n188 VSUBS 0.006939f
C229 B.n189 VSUBS 0.006939f
C230 B.n190 VSUBS 0.006939f
C231 B.n191 VSUBS 0.006939f
C232 B.n192 VSUBS 0.006939f
C233 B.n193 VSUBS 0.006939f
C234 B.n194 VSUBS 0.006939f
C235 B.n195 VSUBS 0.006939f
C236 B.n196 VSUBS 0.006939f
C237 B.n197 VSUBS 0.006939f
C238 B.n198 VSUBS 0.006939f
C239 B.n199 VSUBS 0.006939f
C240 B.n200 VSUBS 0.006939f
C241 B.n201 VSUBS 0.006939f
C242 B.n202 VSUBS 0.006939f
C243 B.n203 VSUBS 0.006939f
C244 B.n204 VSUBS 0.006939f
C245 B.n205 VSUBS 0.006939f
C246 B.n206 VSUBS 0.006939f
C247 B.n207 VSUBS 0.01651f
C248 B.n208 VSUBS 0.01651f
C249 B.n209 VSUBS 0.01757f
C250 B.n210 VSUBS 0.006939f
C251 B.n211 VSUBS 0.006939f
C252 B.n212 VSUBS 0.006939f
C253 B.n213 VSUBS 0.006939f
C254 B.n214 VSUBS 0.006939f
C255 B.n215 VSUBS 0.006939f
C256 B.n216 VSUBS 0.006939f
C257 B.n217 VSUBS 0.006939f
C258 B.n218 VSUBS 0.006939f
C259 B.n219 VSUBS 0.006939f
C260 B.n220 VSUBS 0.006939f
C261 B.n221 VSUBS 0.006939f
C262 B.n222 VSUBS 0.006939f
C263 B.n223 VSUBS 0.006939f
C264 B.n224 VSUBS 0.006939f
C265 B.n225 VSUBS 0.006939f
C266 B.n226 VSUBS 0.006939f
C267 B.n227 VSUBS 0.006939f
C268 B.n228 VSUBS 0.006939f
C269 B.n229 VSUBS 0.006939f
C270 B.n230 VSUBS 0.006939f
C271 B.n231 VSUBS 0.006939f
C272 B.n232 VSUBS 0.006939f
C273 B.n233 VSUBS 0.006939f
C274 B.n234 VSUBS 0.006939f
C275 B.n235 VSUBS 0.006939f
C276 B.n236 VSUBS 0.006939f
C277 B.n237 VSUBS 0.006939f
C278 B.n238 VSUBS 0.006939f
C279 B.n239 VSUBS 0.006939f
C280 B.n240 VSUBS 0.006939f
C281 B.n241 VSUBS 0.006939f
C282 B.n242 VSUBS 0.006939f
C283 B.n243 VSUBS 0.006939f
C284 B.n244 VSUBS 0.006939f
C285 B.n245 VSUBS 0.006939f
C286 B.n246 VSUBS 0.006939f
C287 B.n247 VSUBS 0.006939f
C288 B.n248 VSUBS 0.006939f
C289 B.n249 VSUBS 0.006939f
C290 B.n250 VSUBS 0.006939f
C291 B.n251 VSUBS 0.006939f
C292 B.n252 VSUBS 0.006939f
C293 B.n253 VSUBS 0.006939f
C294 B.n254 VSUBS 0.006939f
C295 B.n255 VSUBS 0.006939f
C296 B.n256 VSUBS 0.006939f
C297 B.n257 VSUBS 0.006939f
C298 B.n258 VSUBS 0.006939f
C299 B.n259 VSUBS 0.006939f
C300 B.n260 VSUBS 0.006939f
C301 B.n261 VSUBS 0.006939f
C302 B.n262 VSUBS 0.006939f
C303 B.n263 VSUBS 0.006939f
C304 B.n264 VSUBS 0.006939f
C305 B.n265 VSUBS 0.006939f
C306 B.n266 VSUBS 0.006939f
C307 B.n267 VSUBS 0.006939f
C308 B.n268 VSUBS 0.006939f
C309 B.n269 VSUBS 0.006939f
C310 B.n270 VSUBS 0.006939f
C311 B.n271 VSUBS 0.00653f
C312 B.n272 VSUBS 0.016076f
C313 B.n273 VSUBS 0.003877f
C314 B.n274 VSUBS 0.006939f
C315 B.n275 VSUBS 0.006939f
C316 B.n276 VSUBS 0.006939f
C317 B.n277 VSUBS 0.006939f
C318 B.n278 VSUBS 0.006939f
C319 B.n279 VSUBS 0.006939f
C320 B.n280 VSUBS 0.006939f
C321 B.n281 VSUBS 0.006939f
C322 B.n282 VSUBS 0.006939f
C323 B.n283 VSUBS 0.006939f
C324 B.n284 VSUBS 0.006939f
C325 B.n285 VSUBS 0.006939f
C326 B.n286 VSUBS 0.003877f
C327 B.n287 VSUBS 0.006939f
C328 B.n288 VSUBS 0.006939f
C329 B.n289 VSUBS 0.00653f
C330 B.n290 VSUBS 0.006939f
C331 B.n291 VSUBS 0.006939f
C332 B.n292 VSUBS 0.006939f
C333 B.n293 VSUBS 0.006939f
C334 B.n294 VSUBS 0.006939f
C335 B.n295 VSUBS 0.006939f
C336 B.n296 VSUBS 0.006939f
C337 B.n297 VSUBS 0.006939f
C338 B.n298 VSUBS 0.006939f
C339 B.n299 VSUBS 0.006939f
C340 B.n300 VSUBS 0.006939f
C341 B.n301 VSUBS 0.006939f
C342 B.n302 VSUBS 0.006939f
C343 B.n303 VSUBS 0.006939f
C344 B.n304 VSUBS 0.006939f
C345 B.n305 VSUBS 0.006939f
C346 B.n306 VSUBS 0.006939f
C347 B.n307 VSUBS 0.006939f
C348 B.n308 VSUBS 0.006939f
C349 B.n309 VSUBS 0.006939f
C350 B.n310 VSUBS 0.006939f
C351 B.n311 VSUBS 0.006939f
C352 B.n312 VSUBS 0.006939f
C353 B.n313 VSUBS 0.006939f
C354 B.n314 VSUBS 0.006939f
C355 B.n315 VSUBS 0.006939f
C356 B.n316 VSUBS 0.006939f
C357 B.n317 VSUBS 0.006939f
C358 B.n318 VSUBS 0.006939f
C359 B.n319 VSUBS 0.006939f
C360 B.n320 VSUBS 0.006939f
C361 B.n321 VSUBS 0.006939f
C362 B.n322 VSUBS 0.006939f
C363 B.n323 VSUBS 0.006939f
C364 B.n324 VSUBS 0.006939f
C365 B.n325 VSUBS 0.006939f
C366 B.n326 VSUBS 0.006939f
C367 B.n327 VSUBS 0.006939f
C368 B.n328 VSUBS 0.006939f
C369 B.n329 VSUBS 0.006939f
C370 B.n330 VSUBS 0.006939f
C371 B.n331 VSUBS 0.006939f
C372 B.n332 VSUBS 0.006939f
C373 B.n333 VSUBS 0.006939f
C374 B.n334 VSUBS 0.006939f
C375 B.n335 VSUBS 0.006939f
C376 B.n336 VSUBS 0.006939f
C377 B.n337 VSUBS 0.006939f
C378 B.n338 VSUBS 0.006939f
C379 B.n339 VSUBS 0.006939f
C380 B.n340 VSUBS 0.006939f
C381 B.n341 VSUBS 0.006939f
C382 B.n342 VSUBS 0.006939f
C383 B.n343 VSUBS 0.006939f
C384 B.n344 VSUBS 0.006939f
C385 B.n345 VSUBS 0.006939f
C386 B.n346 VSUBS 0.006939f
C387 B.n347 VSUBS 0.006939f
C388 B.n348 VSUBS 0.006939f
C389 B.n349 VSUBS 0.006939f
C390 B.n350 VSUBS 0.01757f
C391 B.n351 VSUBS 0.01651f
C392 B.n352 VSUBS 0.01651f
C393 B.n353 VSUBS 0.006939f
C394 B.n354 VSUBS 0.006939f
C395 B.n355 VSUBS 0.006939f
C396 B.n356 VSUBS 0.006939f
C397 B.n357 VSUBS 0.006939f
C398 B.n358 VSUBS 0.006939f
C399 B.n359 VSUBS 0.006939f
C400 B.n360 VSUBS 0.006939f
C401 B.n361 VSUBS 0.006939f
C402 B.n362 VSUBS 0.006939f
C403 B.n363 VSUBS 0.006939f
C404 B.n364 VSUBS 0.006939f
C405 B.n365 VSUBS 0.006939f
C406 B.n366 VSUBS 0.006939f
C407 B.n367 VSUBS 0.006939f
C408 B.n368 VSUBS 0.006939f
C409 B.n369 VSUBS 0.006939f
C410 B.n370 VSUBS 0.006939f
C411 B.n371 VSUBS 0.006939f
C412 B.n372 VSUBS 0.006939f
C413 B.n373 VSUBS 0.006939f
C414 B.n374 VSUBS 0.006939f
C415 B.n375 VSUBS 0.006939f
C416 B.n376 VSUBS 0.006939f
C417 B.n377 VSUBS 0.006939f
C418 B.n378 VSUBS 0.006939f
C419 B.n379 VSUBS 0.006939f
C420 B.n380 VSUBS 0.006939f
C421 B.n381 VSUBS 0.006939f
C422 B.n382 VSUBS 0.006939f
C423 B.n383 VSUBS 0.006939f
C424 B.n384 VSUBS 0.006939f
C425 B.n385 VSUBS 0.006939f
C426 B.n386 VSUBS 0.006939f
C427 B.n387 VSUBS 0.006939f
C428 B.n388 VSUBS 0.006939f
C429 B.n389 VSUBS 0.006939f
C430 B.n390 VSUBS 0.006939f
C431 B.n391 VSUBS 0.006939f
C432 B.n392 VSUBS 0.006939f
C433 B.n393 VSUBS 0.006939f
C434 B.n394 VSUBS 0.006939f
C435 B.n395 VSUBS 0.006939f
C436 B.n396 VSUBS 0.006939f
C437 B.n397 VSUBS 0.006939f
C438 B.n398 VSUBS 0.006939f
C439 B.n399 VSUBS 0.006939f
C440 B.n400 VSUBS 0.006939f
C441 B.n401 VSUBS 0.006939f
C442 B.n402 VSUBS 0.006939f
C443 B.n403 VSUBS 0.006939f
C444 B.n404 VSUBS 0.006939f
C445 B.n405 VSUBS 0.006939f
C446 B.n406 VSUBS 0.006939f
C447 B.n407 VSUBS 0.006939f
C448 B.n408 VSUBS 0.006939f
C449 B.n409 VSUBS 0.006939f
C450 B.n410 VSUBS 0.006939f
C451 B.n411 VSUBS 0.006939f
C452 B.n412 VSUBS 0.006939f
C453 B.n413 VSUBS 0.006939f
C454 B.n414 VSUBS 0.006939f
C455 B.n415 VSUBS 0.006939f
C456 B.n416 VSUBS 0.006939f
C457 B.n417 VSUBS 0.006939f
C458 B.n418 VSUBS 0.006939f
C459 B.n419 VSUBS 0.006939f
C460 B.n420 VSUBS 0.006939f
C461 B.n421 VSUBS 0.006939f
C462 B.n422 VSUBS 0.006939f
C463 B.n423 VSUBS 0.006939f
C464 B.n424 VSUBS 0.006939f
C465 B.n425 VSUBS 0.006939f
C466 B.n426 VSUBS 0.006939f
C467 B.n427 VSUBS 0.006939f
C468 B.n428 VSUBS 0.006939f
C469 B.n429 VSUBS 0.006939f
C470 B.n430 VSUBS 0.006939f
C471 B.n431 VSUBS 0.006939f
C472 B.n432 VSUBS 0.006939f
C473 B.n433 VSUBS 0.006939f
C474 B.n434 VSUBS 0.006939f
C475 B.n435 VSUBS 0.006939f
C476 B.n436 VSUBS 0.006939f
C477 B.n437 VSUBS 0.006939f
C478 B.n438 VSUBS 0.006939f
C479 B.n439 VSUBS 0.006939f
C480 B.n440 VSUBS 0.006939f
C481 B.n441 VSUBS 0.017273f
C482 B.n442 VSUBS 0.01651f
C483 B.n443 VSUBS 0.01757f
C484 B.n444 VSUBS 0.006939f
C485 B.n445 VSUBS 0.006939f
C486 B.n446 VSUBS 0.006939f
C487 B.n447 VSUBS 0.006939f
C488 B.n448 VSUBS 0.006939f
C489 B.n449 VSUBS 0.006939f
C490 B.n450 VSUBS 0.006939f
C491 B.n451 VSUBS 0.006939f
C492 B.n452 VSUBS 0.006939f
C493 B.n453 VSUBS 0.006939f
C494 B.n454 VSUBS 0.006939f
C495 B.n455 VSUBS 0.006939f
C496 B.n456 VSUBS 0.006939f
C497 B.n457 VSUBS 0.006939f
C498 B.n458 VSUBS 0.006939f
C499 B.n459 VSUBS 0.006939f
C500 B.n460 VSUBS 0.006939f
C501 B.n461 VSUBS 0.006939f
C502 B.n462 VSUBS 0.006939f
C503 B.n463 VSUBS 0.006939f
C504 B.n464 VSUBS 0.006939f
C505 B.n465 VSUBS 0.006939f
C506 B.n466 VSUBS 0.006939f
C507 B.n467 VSUBS 0.006939f
C508 B.n468 VSUBS 0.006939f
C509 B.n469 VSUBS 0.006939f
C510 B.n470 VSUBS 0.006939f
C511 B.n471 VSUBS 0.006939f
C512 B.n472 VSUBS 0.006939f
C513 B.n473 VSUBS 0.006939f
C514 B.n474 VSUBS 0.006939f
C515 B.n475 VSUBS 0.006939f
C516 B.n476 VSUBS 0.006939f
C517 B.n477 VSUBS 0.006939f
C518 B.n478 VSUBS 0.006939f
C519 B.n479 VSUBS 0.006939f
C520 B.n480 VSUBS 0.006939f
C521 B.n481 VSUBS 0.006939f
C522 B.n482 VSUBS 0.006939f
C523 B.n483 VSUBS 0.006939f
C524 B.n484 VSUBS 0.006939f
C525 B.n485 VSUBS 0.006939f
C526 B.n486 VSUBS 0.006939f
C527 B.n487 VSUBS 0.006939f
C528 B.n488 VSUBS 0.006939f
C529 B.n489 VSUBS 0.006939f
C530 B.n490 VSUBS 0.006939f
C531 B.n491 VSUBS 0.006939f
C532 B.n492 VSUBS 0.006939f
C533 B.n493 VSUBS 0.006939f
C534 B.n494 VSUBS 0.006939f
C535 B.n495 VSUBS 0.006939f
C536 B.n496 VSUBS 0.006939f
C537 B.n497 VSUBS 0.006939f
C538 B.n498 VSUBS 0.006939f
C539 B.n499 VSUBS 0.006939f
C540 B.n500 VSUBS 0.006939f
C541 B.n501 VSUBS 0.006939f
C542 B.n502 VSUBS 0.006939f
C543 B.n503 VSUBS 0.006939f
C544 B.n504 VSUBS 0.006939f
C545 B.n505 VSUBS 0.00653f
C546 B.n506 VSUBS 0.016076f
C547 B.n507 VSUBS 0.003877f
C548 B.n508 VSUBS 0.006939f
C549 B.n509 VSUBS 0.006939f
C550 B.n510 VSUBS 0.006939f
C551 B.n511 VSUBS 0.006939f
C552 B.n512 VSUBS 0.006939f
C553 B.n513 VSUBS 0.006939f
C554 B.n514 VSUBS 0.006939f
C555 B.n515 VSUBS 0.006939f
C556 B.n516 VSUBS 0.006939f
C557 B.n517 VSUBS 0.006939f
C558 B.n518 VSUBS 0.006939f
C559 B.n519 VSUBS 0.006939f
C560 B.n520 VSUBS 0.003877f
C561 B.n521 VSUBS 0.006939f
C562 B.n522 VSUBS 0.006939f
C563 B.n523 VSUBS 0.00653f
C564 B.n524 VSUBS 0.006939f
C565 B.n525 VSUBS 0.006939f
C566 B.n526 VSUBS 0.006939f
C567 B.n527 VSUBS 0.006939f
C568 B.n528 VSUBS 0.006939f
C569 B.n529 VSUBS 0.006939f
C570 B.n530 VSUBS 0.006939f
C571 B.n531 VSUBS 0.006939f
C572 B.n532 VSUBS 0.006939f
C573 B.n533 VSUBS 0.006939f
C574 B.n534 VSUBS 0.006939f
C575 B.n535 VSUBS 0.006939f
C576 B.n536 VSUBS 0.006939f
C577 B.n537 VSUBS 0.006939f
C578 B.n538 VSUBS 0.006939f
C579 B.n539 VSUBS 0.006939f
C580 B.n540 VSUBS 0.006939f
C581 B.n541 VSUBS 0.006939f
C582 B.n542 VSUBS 0.006939f
C583 B.n543 VSUBS 0.006939f
C584 B.n544 VSUBS 0.006939f
C585 B.n545 VSUBS 0.006939f
C586 B.n546 VSUBS 0.006939f
C587 B.n547 VSUBS 0.006939f
C588 B.n548 VSUBS 0.006939f
C589 B.n549 VSUBS 0.006939f
C590 B.n550 VSUBS 0.006939f
C591 B.n551 VSUBS 0.006939f
C592 B.n552 VSUBS 0.006939f
C593 B.n553 VSUBS 0.006939f
C594 B.n554 VSUBS 0.006939f
C595 B.n555 VSUBS 0.006939f
C596 B.n556 VSUBS 0.006939f
C597 B.n557 VSUBS 0.006939f
C598 B.n558 VSUBS 0.006939f
C599 B.n559 VSUBS 0.006939f
C600 B.n560 VSUBS 0.006939f
C601 B.n561 VSUBS 0.006939f
C602 B.n562 VSUBS 0.006939f
C603 B.n563 VSUBS 0.006939f
C604 B.n564 VSUBS 0.006939f
C605 B.n565 VSUBS 0.006939f
C606 B.n566 VSUBS 0.006939f
C607 B.n567 VSUBS 0.006939f
C608 B.n568 VSUBS 0.006939f
C609 B.n569 VSUBS 0.006939f
C610 B.n570 VSUBS 0.006939f
C611 B.n571 VSUBS 0.006939f
C612 B.n572 VSUBS 0.006939f
C613 B.n573 VSUBS 0.006939f
C614 B.n574 VSUBS 0.006939f
C615 B.n575 VSUBS 0.006939f
C616 B.n576 VSUBS 0.006939f
C617 B.n577 VSUBS 0.006939f
C618 B.n578 VSUBS 0.006939f
C619 B.n579 VSUBS 0.006939f
C620 B.n580 VSUBS 0.006939f
C621 B.n581 VSUBS 0.006939f
C622 B.n582 VSUBS 0.006939f
C623 B.n583 VSUBS 0.006939f
C624 B.n584 VSUBS 0.01757f
C625 B.n585 VSUBS 0.01651f
C626 B.n586 VSUBS 0.01651f
C627 B.n587 VSUBS 0.006939f
C628 B.n588 VSUBS 0.006939f
C629 B.n589 VSUBS 0.006939f
C630 B.n590 VSUBS 0.006939f
C631 B.n591 VSUBS 0.006939f
C632 B.n592 VSUBS 0.006939f
C633 B.n593 VSUBS 0.006939f
C634 B.n594 VSUBS 0.006939f
C635 B.n595 VSUBS 0.006939f
C636 B.n596 VSUBS 0.006939f
C637 B.n597 VSUBS 0.006939f
C638 B.n598 VSUBS 0.006939f
C639 B.n599 VSUBS 0.006939f
C640 B.n600 VSUBS 0.006939f
C641 B.n601 VSUBS 0.006939f
C642 B.n602 VSUBS 0.006939f
C643 B.n603 VSUBS 0.006939f
C644 B.n604 VSUBS 0.006939f
C645 B.n605 VSUBS 0.006939f
C646 B.n606 VSUBS 0.006939f
C647 B.n607 VSUBS 0.006939f
C648 B.n608 VSUBS 0.006939f
C649 B.n609 VSUBS 0.006939f
C650 B.n610 VSUBS 0.006939f
C651 B.n611 VSUBS 0.006939f
C652 B.n612 VSUBS 0.006939f
C653 B.n613 VSUBS 0.006939f
C654 B.n614 VSUBS 0.006939f
C655 B.n615 VSUBS 0.006939f
C656 B.n616 VSUBS 0.006939f
C657 B.n617 VSUBS 0.006939f
C658 B.n618 VSUBS 0.006939f
C659 B.n619 VSUBS 0.006939f
C660 B.n620 VSUBS 0.006939f
C661 B.n621 VSUBS 0.006939f
C662 B.n622 VSUBS 0.006939f
C663 B.n623 VSUBS 0.006939f
C664 B.n624 VSUBS 0.006939f
C665 B.n625 VSUBS 0.006939f
C666 B.n626 VSUBS 0.006939f
C667 B.n627 VSUBS 0.006939f
C668 B.n628 VSUBS 0.006939f
C669 B.n629 VSUBS 0.006939f
C670 B.n630 VSUBS 0.006939f
C671 B.n631 VSUBS 0.015711f
C672 VDD2.t0 VSUBS 0.259178f
C673 VDD2.t1 VSUBS 0.259178f
C674 VDD2.n0 VSUBS 2.71425f
C675 VDD2.t3 VSUBS 0.259178f
C676 VDD2.t2 VSUBS 0.259178f
C677 VDD2.n1 VSUBS 2.03342f
C678 VDD2.n2 VSUBS 4.22239f
C679 VN.t3 VSUBS 2.84478f
C680 VN.t2 VSUBS 2.84059f
C681 VN.n0 VSUBS 1.89163f
C682 VN.t1 VSUBS 2.84478f
C683 VN.t0 VSUBS 2.84059f
C684 VN.n1 VSUBS 3.6698f
C685 VTAIL.n0 VSUBS 0.026261f
C686 VTAIL.n1 VSUBS 0.023271f
C687 VTAIL.n2 VSUBS 0.012505f
C688 VTAIL.n3 VSUBS 0.029556f
C689 VTAIL.n4 VSUBS 0.01324f
C690 VTAIL.n5 VSUBS 0.023271f
C691 VTAIL.n6 VSUBS 0.012505f
C692 VTAIL.n7 VSUBS 0.029556f
C693 VTAIL.n8 VSUBS 0.01324f
C694 VTAIL.n9 VSUBS 0.023271f
C695 VTAIL.n10 VSUBS 0.012872f
C696 VTAIL.n11 VSUBS 0.029556f
C697 VTAIL.n12 VSUBS 0.01324f
C698 VTAIL.n13 VSUBS 0.023271f
C699 VTAIL.n14 VSUBS 0.012505f
C700 VTAIL.n15 VSUBS 0.029556f
C701 VTAIL.n16 VSUBS 0.01324f
C702 VTAIL.n17 VSUBS 0.023271f
C703 VTAIL.n18 VSUBS 0.012505f
C704 VTAIL.n19 VSUBS 0.022167f
C705 VTAIL.n20 VSUBS 0.022234f
C706 VTAIL.t0 VSUBS 0.063708f
C707 VTAIL.n21 VSUBS 0.185376f
C708 VTAIL.n22 VSUBS 1.16375f
C709 VTAIL.n23 VSUBS 0.012505f
C710 VTAIL.n24 VSUBS 0.01324f
C711 VTAIL.n25 VSUBS 0.029556f
C712 VTAIL.n26 VSUBS 0.029556f
C713 VTAIL.n27 VSUBS 0.01324f
C714 VTAIL.n28 VSUBS 0.012505f
C715 VTAIL.n29 VSUBS 0.023271f
C716 VTAIL.n30 VSUBS 0.023271f
C717 VTAIL.n31 VSUBS 0.012505f
C718 VTAIL.n32 VSUBS 0.01324f
C719 VTAIL.n33 VSUBS 0.029556f
C720 VTAIL.n34 VSUBS 0.029556f
C721 VTAIL.n35 VSUBS 0.01324f
C722 VTAIL.n36 VSUBS 0.012505f
C723 VTAIL.n37 VSUBS 0.023271f
C724 VTAIL.n38 VSUBS 0.023271f
C725 VTAIL.n39 VSUBS 0.012505f
C726 VTAIL.n40 VSUBS 0.012505f
C727 VTAIL.n41 VSUBS 0.01324f
C728 VTAIL.n42 VSUBS 0.029556f
C729 VTAIL.n43 VSUBS 0.029556f
C730 VTAIL.n44 VSUBS 0.029556f
C731 VTAIL.n45 VSUBS 0.012872f
C732 VTAIL.n46 VSUBS 0.012505f
C733 VTAIL.n47 VSUBS 0.023271f
C734 VTAIL.n48 VSUBS 0.023271f
C735 VTAIL.n49 VSUBS 0.012505f
C736 VTAIL.n50 VSUBS 0.01324f
C737 VTAIL.n51 VSUBS 0.029556f
C738 VTAIL.n52 VSUBS 0.029556f
C739 VTAIL.n53 VSUBS 0.01324f
C740 VTAIL.n54 VSUBS 0.012505f
C741 VTAIL.n55 VSUBS 0.023271f
C742 VTAIL.n56 VSUBS 0.023271f
C743 VTAIL.n57 VSUBS 0.012505f
C744 VTAIL.n58 VSUBS 0.01324f
C745 VTAIL.n59 VSUBS 0.029556f
C746 VTAIL.n60 VSUBS 0.07391f
C747 VTAIL.n61 VSUBS 0.01324f
C748 VTAIL.n62 VSUBS 0.012505f
C749 VTAIL.n63 VSUBS 0.056332f
C750 VTAIL.n64 VSUBS 0.03735f
C751 VTAIL.n65 VSUBS 0.142029f
C752 VTAIL.n66 VSUBS 0.026261f
C753 VTAIL.n67 VSUBS 0.023271f
C754 VTAIL.n68 VSUBS 0.012505f
C755 VTAIL.n69 VSUBS 0.029556f
C756 VTAIL.n70 VSUBS 0.01324f
C757 VTAIL.n71 VSUBS 0.023271f
C758 VTAIL.n72 VSUBS 0.012505f
C759 VTAIL.n73 VSUBS 0.029556f
C760 VTAIL.n74 VSUBS 0.01324f
C761 VTAIL.n75 VSUBS 0.023271f
C762 VTAIL.n76 VSUBS 0.012872f
C763 VTAIL.n77 VSUBS 0.029556f
C764 VTAIL.n78 VSUBS 0.01324f
C765 VTAIL.n79 VSUBS 0.023271f
C766 VTAIL.n80 VSUBS 0.012505f
C767 VTAIL.n81 VSUBS 0.029556f
C768 VTAIL.n82 VSUBS 0.01324f
C769 VTAIL.n83 VSUBS 0.023271f
C770 VTAIL.n84 VSUBS 0.012505f
C771 VTAIL.n85 VSUBS 0.022167f
C772 VTAIL.n86 VSUBS 0.022234f
C773 VTAIL.t5 VSUBS 0.063708f
C774 VTAIL.n87 VSUBS 0.185376f
C775 VTAIL.n88 VSUBS 1.16375f
C776 VTAIL.n89 VSUBS 0.012505f
C777 VTAIL.n90 VSUBS 0.01324f
C778 VTAIL.n91 VSUBS 0.029556f
C779 VTAIL.n92 VSUBS 0.029556f
C780 VTAIL.n93 VSUBS 0.01324f
C781 VTAIL.n94 VSUBS 0.012505f
C782 VTAIL.n95 VSUBS 0.023271f
C783 VTAIL.n96 VSUBS 0.023271f
C784 VTAIL.n97 VSUBS 0.012505f
C785 VTAIL.n98 VSUBS 0.01324f
C786 VTAIL.n99 VSUBS 0.029556f
C787 VTAIL.n100 VSUBS 0.029556f
C788 VTAIL.n101 VSUBS 0.01324f
C789 VTAIL.n102 VSUBS 0.012505f
C790 VTAIL.n103 VSUBS 0.023271f
C791 VTAIL.n104 VSUBS 0.023271f
C792 VTAIL.n105 VSUBS 0.012505f
C793 VTAIL.n106 VSUBS 0.012505f
C794 VTAIL.n107 VSUBS 0.01324f
C795 VTAIL.n108 VSUBS 0.029556f
C796 VTAIL.n109 VSUBS 0.029556f
C797 VTAIL.n110 VSUBS 0.029556f
C798 VTAIL.n111 VSUBS 0.012872f
C799 VTAIL.n112 VSUBS 0.012505f
C800 VTAIL.n113 VSUBS 0.023271f
C801 VTAIL.n114 VSUBS 0.023271f
C802 VTAIL.n115 VSUBS 0.012505f
C803 VTAIL.n116 VSUBS 0.01324f
C804 VTAIL.n117 VSUBS 0.029556f
C805 VTAIL.n118 VSUBS 0.029556f
C806 VTAIL.n119 VSUBS 0.01324f
C807 VTAIL.n120 VSUBS 0.012505f
C808 VTAIL.n121 VSUBS 0.023271f
C809 VTAIL.n122 VSUBS 0.023271f
C810 VTAIL.n123 VSUBS 0.012505f
C811 VTAIL.n124 VSUBS 0.01324f
C812 VTAIL.n125 VSUBS 0.029556f
C813 VTAIL.n126 VSUBS 0.07391f
C814 VTAIL.n127 VSUBS 0.01324f
C815 VTAIL.n128 VSUBS 0.012505f
C816 VTAIL.n129 VSUBS 0.056332f
C817 VTAIL.n130 VSUBS 0.03735f
C818 VTAIL.n131 VSUBS 0.21879f
C819 VTAIL.n132 VSUBS 0.026261f
C820 VTAIL.n133 VSUBS 0.023271f
C821 VTAIL.n134 VSUBS 0.012505f
C822 VTAIL.n135 VSUBS 0.029556f
C823 VTAIL.n136 VSUBS 0.01324f
C824 VTAIL.n137 VSUBS 0.023271f
C825 VTAIL.n138 VSUBS 0.012505f
C826 VTAIL.n139 VSUBS 0.029556f
C827 VTAIL.n140 VSUBS 0.01324f
C828 VTAIL.n141 VSUBS 0.023271f
C829 VTAIL.n142 VSUBS 0.012872f
C830 VTAIL.n143 VSUBS 0.029556f
C831 VTAIL.n144 VSUBS 0.01324f
C832 VTAIL.n145 VSUBS 0.023271f
C833 VTAIL.n146 VSUBS 0.012505f
C834 VTAIL.n147 VSUBS 0.029556f
C835 VTAIL.n148 VSUBS 0.01324f
C836 VTAIL.n149 VSUBS 0.023271f
C837 VTAIL.n150 VSUBS 0.012505f
C838 VTAIL.n151 VSUBS 0.022167f
C839 VTAIL.n152 VSUBS 0.022234f
C840 VTAIL.t7 VSUBS 0.063708f
C841 VTAIL.n153 VSUBS 0.185376f
C842 VTAIL.n154 VSUBS 1.16375f
C843 VTAIL.n155 VSUBS 0.012505f
C844 VTAIL.n156 VSUBS 0.01324f
C845 VTAIL.n157 VSUBS 0.029556f
C846 VTAIL.n158 VSUBS 0.029556f
C847 VTAIL.n159 VSUBS 0.01324f
C848 VTAIL.n160 VSUBS 0.012505f
C849 VTAIL.n161 VSUBS 0.023271f
C850 VTAIL.n162 VSUBS 0.023271f
C851 VTAIL.n163 VSUBS 0.012505f
C852 VTAIL.n164 VSUBS 0.01324f
C853 VTAIL.n165 VSUBS 0.029556f
C854 VTAIL.n166 VSUBS 0.029556f
C855 VTAIL.n167 VSUBS 0.01324f
C856 VTAIL.n168 VSUBS 0.012505f
C857 VTAIL.n169 VSUBS 0.023271f
C858 VTAIL.n170 VSUBS 0.023271f
C859 VTAIL.n171 VSUBS 0.012505f
C860 VTAIL.n172 VSUBS 0.012505f
C861 VTAIL.n173 VSUBS 0.01324f
C862 VTAIL.n174 VSUBS 0.029556f
C863 VTAIL.n175 VSUBS 0.029556f
C864 VTAIL.n176 VSUBS 0.029556f
C865 VTAIL.n177 VSUBS 0.012872f
C866 VTAIL.n178 VSUBS 0.012505f
C867 VTAIL.n179 VSUBS 0.023271f
C868 VTAIL.n180 VSUBS 0.023271f
C869 VTAIL.n181 VSUBS 0.012505f
C870 VTAIL.n182 VSUBS 0.01324f
C871 VTAIL.n183 VSUBS 0.029556f
C872 VTAIL.n184 VSUBS 0.029556f
C873 VTAIL.n185 VSUBS 0.01324f
C874 VTAIL.n186 VSUBS 0.012505f
C875 VTAIL.n187 VSUBS 0.023271f
C876 VTAIL.n188 VSUBS 0.023271f
C877 VTAIL.n189 VSUBS 0.012505f
C878 VTAIL.n190 VSUBS 0.01324f
C879 VTAIL.n191 VSUBS 0.029556f
C880 VTAIL.n192 VSUBS 0.07391f
C881 VTAIL.n193 VSUBS 0.01324f
C882 VTAIL.n194 VSUBS 0.012505f
C883 VTAIL.n195 VSUBS 0.056332f
C884 VTAIL.n196 VSUBS 0.03735f
C885 VTAIL.n197 VSUBS 1.45053f
C886 VTAIL.n198 VSUBS 0.026261f
C887 VTAIL.n199 VSUBS 0.023271f
C888 VTAIL.n200 VSUBS 0.012505f
C889 VTAIL.n201 VSUBS 0.029556f
C890 VTAIL.n202 VSUBS 0.01324f
C891 VTAIL.n203 VSUBS 0.023271f
C892 VTAIL.n204 VSUBS 0.012505f
C893 VTAIL.n205 VSUBS 0.029556f
C894 VTAIL.n206 VSUBS 0.01324f
C895 VTAIL.n207 VSUBS 0.023271f
C896 VTAIL.n208 VSUBS 0.012872f
C897 VTAIL.n209 VSUBS 0.029556f
C898 VTAIL.n210 VSUBS 0.012505f
C899 VTAIL.n211 VSUBS 0.01324f
C900 VTAIL.n212 VSUBS 0.023271f
C901 VTAIL.n213 VSUBS 0.012505f
C902 VTAIL.n214 VSUBS 0.029556f
C903 VTAIL.n215 VSUBS 0.01324f
C904 VTAIL.n216 VSUBS 0.023271f
C905 VTAIL.n217 VSUBS 0.012505f
C906 VTAIL.n218 VSUBS 0.022167f
C907 VTAIL.n219 VSUBS 0.022234f
C908 VTAIL.t1 VSUBS 0.063708f
C909 VTAIL.n220 VSUBS 0.185376f
C910 VTAIL.n221 VSUBS 1.16375f
C911 VTAIL.n222 VSUBS 0.012505f
C912 VTAIL.n223 VSUBS 0.01324f
C913 VTAIL.n224 VSUBS 0.029556f
C914 VTAIL.n225 VSUBS 0.029556f
C915 VTAIL.n226 VSUBS 0.01324f
C916 VTAIL.n227 VSUBS 0.012505f
C917 VTAIL.n228 VSUBS 0.023271f
C918 VTAIL.n229 VSUBS 0.023271f
C919 VTAIL.n230 VSUBS 0.012505f
C920 VTAIL.n231 VSUBS 0.01324f
C921 VTAIL.n232 VSUBS 0.029556f
C922 VTAIL.n233 VSUBS 0.029556f
C923 VTAIL.n234 VSUBS 0.01324f
C924 VTAIL.n235 VSUBS 0.012505f
C925 VTAIL.n236 VSUBS 0.023271f
C926 VTAIL.n237 VSUBS 0.023271f
C927 VTAIL.n238 VSUBS 0.012505f
C928 VTAIL.n239 VSUBS 0.01324f
C929 VTAIL.n240 VSUBS 0.029556f
C930 VTAIL.n241 VSUBS 0.029556f
C931 VTAIL.n242 VSUBS 0.029556f
C932 VTAIL.n243 VSUBS 0.012872f
C933 VTAIL.n244 VSUBS 0.012505f
C934 VTAIL.n245 VSUBS 0.023271f
C935 VTAIL.n246 VSUBS 0.023271f
C936 VTAIL.n247 VSUBS 0.012505f
C937 VTAIL.n248 VSUBS 0.01324f
C938 VTAIL.n249 VSUBS 0.029556f
C939 VTAIL.n250 VSUBS 0.029556f
C940 VTAIL.n251 VSUBS 0.01324f
C941 VTAIL.n252 VSUBS 0.012505f
C942 VTAIL.n253 VSUBS 0.023271f
C943 VTAIL.n254 VSUBS 0.023271f
C944 VTAIL.n255 VSUBS 0.012505f
C945 VTAIL.n256 VSUBS 0.01324f
C946 VTAIL.n257 VSUBS 0.029556f
C947 VTAIL.n258 VSUBS 0.07391f
C948 VTAIL.n259 VSUBS 0.01324f
C949 VTAIL.n260 VSUBS 0.012505f
C950 VTAIL.n261 VSUBS 0.056332f
C951 VTAIL.n262 VSUBS 0.03735f
C952 VTAIL.n263 VSUBS 1.45053f
C953 VTAIL.n264 VSUBS 0.026261f
C954 VTAIL.n265 VSUBS 0.023271f
C955 VTAIL.n266 VSUBS 0.012505f
C956 VTAIL.n267 VSUBS 0.029556f
C957 VTAIL.n268 VSUBS 0.01324f
C958 VTAIL.n269 VSUBS 0.023271f
C959 VTAIL.n270 VSUBS 0.012505f
C960 VTAIL.n271 VSUBS 0.029556f
C961 VTAIL.n272 VSUBS 0.01324f
C962 VTAIL.n273 VSUBS 0.023271f
C963 VTAIL.n274 VSUBS 0.012872f
C964 VTAIL.n275 VSUBS 0.029556f
C965 VTAIL.n276 VSUBS 0.012505f
C966 VTAIL.n277 VSUBS 0.01324f
C967 VTAIL.n278 VSUBS 0.023271f
C968 VTAIL.n279 VSUBS 0.012505f
C969 VTAIL.n280 VSUBS 0.029556f
C970 VTAIL.n281 VSUBS 0.01324f
C971 VTAIL.n282 VSUBS 0.023271f
C972 VTAIL.n283 VSUBS 0.012505f
C973 VTAIL.n284 VSUBS 0.022167f
C974 VTAIL.n285 VSUBS 0.022234f
C975 VTAIL.t2 VSUBS 0.063708f
C976 VTAIL.n286 VSUBS 0.185376f
C977 VTAIL.n287 VSUBS 1.16375f
C978 VTAIL.n288 VSUBS 0.012505f
C979 VTAIL.n289 VSUBS 0.01324f
C980 VTAIL.n290 VSUBS 0.029556f
C981 VTAIL.n291 VSUBS 0.029556f
C982 VTAIL.n292 VSUBS 0.01324f
C983 VTAIL.n293 VSUBS 0.012505f
C984 VTAIL.n294 VSUBS 0.023271f
C985 VTAIL.n295 VSUBS 0.023271f
C986 VTAIL.n296 VSUBS 0.012505f
C987 VTAIL.n297 VSUBS 0.01324f
C988 VTAIL.n298 VSUBS 0.029556f
C989 VTAIL.n299 VSUBS 0.029556f
C990 VTAIL.n300 VSUBS 0.01324f
C991 VTAIL.n301 VSUBS 0.012505f
C992 VTAIL.n302 VSUBS 0.023271f
C993 VTAIL.n303 VSUBS 0.023271f
C994 VTAIL.n304 VSUBS 0.012505f
C995 VTAIL.n305 VSUBS 0.01324f
C996 VTAIL.n306 VSUBS 0.029556f
C997 VTAIL.n307 VSUBS 0.029556f
C998 VTAIL.n308 VSUBS 0.029556f
C999 VTAIL.n309 VSUBS 0.012872f
C1000 VTAIL.n310 VSUBS 0.012505f
C1001 VTAIL.n311 VSUBS 0.023271f
C1002 VTAIL.n312 VSUBS 0.023271f
C1003 VTAIL.n313 VSUBS 0.012505f
C1004 VTAIL.n314 VSUBS 0.01324f
C1005 VTAIL.n315 VSUBS 0.029556f
C1006 VTAIL.n316 VSUBS 0.029556f
C1007 VTAIL.n317 VSUBS 0.01324f
C1008 VTAIL.n318 VSUBS 0.012505f
C1009 VTAIL.n319 VSUBS 0.023271f
C1010 VTAIL.n320 VSUBS 0.023271f
C1011 VTAIL.n321 VSUBS 0.012505f
C1012 VTAIL.n322 VSUBS 0.01324f
C1013 VTAIL.n323 VSUBS 0.029556f
C1014 VTAIL.n324 VSUBS 0.07391f
C1015 VTAIL.n325 VSUBS 0.01324f
C1016 VTAIL.n326 VSUBS 0.012505f
C1017 VTAIL.n327 VSUBS 0.056332f
C1018 VTAIL.n328 VSUBS 0.03735f
C1019 VTAIL.n329 VSUBS 0.21879f
C1020 VTAIL.n330 VSUBS 0.026261f
C1021 VTAIL.n331 VSUBS 0.023271f
C1022 VTAIL.n332 VSUBS 0.012505f
C1023 VTAIL.n333 VSUBS 0.029556f
C1024 VTAIL.n334 VSUBS 0.01324f
C1025 VTAIL.n335 VSUBS 0.023271f
C1026 VTAIL.n336 VSUBS 0.012505f
C1027 VTAIL.n337 VSUBS 0.029556f
C1028 VTAIL.n338 VSUBS 0.01324f
C1029 VTAIL.n339 VSUBS 0.023271f
C1030 VTAIL.n340 VSUBS 0.012872f
C1031 VTAIL.n341 VSUBS 0.029556f
C1032 VTAIL.n342 VSUBS 0.012505f
C1033 VTAIL.n343 VSUBS 0.01324f
C1034 VTAIL.n344 VSUBS 0.023271f
C1035 VTAIL.n345 VSUBS 0.012505f
C1036 VTAIL.n346 VSUBS 0.029556f
C1037 VTAIL.n347 VSUBS 0.01324f
C1038 VTAIL.n348 VSUBS 0.023271f
C1039 VTAIL.n349 VSUBS 0.012505f
C1040 VTAIL.n350 VSUBS 0.022167f
C1041 VTAIL.n351 VSUBS 0.022234f
C1042 VTAIL.t4 VSUBS 0.063708f
C1043 VTAIL.n352 VSUBS 0.185376f
C1044 VTAIL.n353 VSUBS 1.16375f
C1045 VTAIL.n354 VSUBS 0.012505f
C1046 VTAIL.n355 VSUBS 0.01324f
C1047 VTAIL.n356 VSUBS 0.029556f
C1048 VTAIL.n357 VSUBS 0.029556f
C1049 VTAIL.n358 VSUBS 0.01324f
C1050 VTAIL.n359 VSUBS 0.012505f
C1051 VTAIL.n360 VSUBS 0.023271f
C1052 VTAIL.n361 VSUBS 0.023271f
C1053 VTAIL.n362 VSUBS 0.012505f
C1054 VTAIL.n363 VSUBS 0.01324f
C1055 VTAIL.n364 VSUBS 0.029556f
C1056 VTAIL.n365 VSUBS 0.029556f
C1057 VTAIL.n366 VSUBS 0.01324f
C1058 VTAIL.n367 VSUBS 0.012505f
C1059 VTAIL.n368 VSUBS 0.023271f
C1060 VTAIL.n369 VSUBS 0.023271f
C1061 VTAIL.n370 VSUBS 0.012505f
C1062 VTAIL.n371 VSUBS 0.01324f
C1063 VTAIL.n372 VSUBS 0.029556f
C1064 VTAIL.n373 VSUBS 0.029556f
C1065 VTAIL.n374 VSUBS 0.029556f
C1066 VTAIL.n375 VSUBS 0.012872f
C1067 VTAIL.n376 VSUBS 0.012505f
C1068 VTAIL.n377 VSUBS 0.023271f
C1069 VTAIL.n378 VSUBS 0.023271f
C1070 VTAIL.n379 VSUBS 0.012505f
C1071 VTAIL.n380 VSUBS 0.01324f
C1072 VTAIL.n381 VSUBS 0.029556f
C1073 VTAIL.n382 VSUBS 0.029556f
C1074 VTAIL.n383 VSUBS 0.01324f
C1075 VTAIL.n384 VSUBS 0.012505f
C1076 VTAIL.n385 VSUBS 0.023271f
C1077 VTAIL.n386 VSUBS 0.023271f
C1078 VTAIL.n387 VSUBS 0.012505f
C1079 VTAIL.n388 VSUBS 0.01324f
C1080 VTAIL.n389 VSUBS 0.029556f
C1081 VTAIL.n390 VSUBS 0.07391f
C1082 VTAIL.n391 VSUBS 0.01324f
C1083 VTAIL.n392 VSUBS 0.012505f
C1084 VTAIL.n393 VSUBS 0.056332f
C1085 VTAIL.n394 VSUBS 0.03735f
C1086 VTAIL.n395 VSUBS 0.21879f
C1087 VTAIL.n396 VSUBS 0.026261f
C1088 VTAIL.n397 VSUBS 0.023271f
C1089 VTAIL.n398 VSUBS 0.012505f
C1090 VTAIL.n399 VSUBS 0.029556f
C1091 VTAIL.n400 VSUBS 0.01324f
C1092 VTAIL.n401 VSUBS 0.023271f
C1093 VTAIL.n402 VSUBS 0.012505f
C1094 VTAIL.n403 VSUBS 0.029556f
C1095 VTAIL.n404 VSUBS 0.01324f
C1096 VTAIL.n405 VSUBS 0.023271f
C1097 VTAIL.n406 VSUBS 0.012872f
C1098 VTAIL.n407 VSUBS 0.029556f
C1099 VTAIL.n408 VSUBS 0.012505f
C1100 VTAIL.n409 VSUBS 0.01324f
C1101 VTAIL.n410 VSUBS 0.023271f
C1102 VTAIL.n411 VSUBS 0.012505f
C1103 VTAIL.n412 VSUBS 0.029556f
C1104 VTAIL.n413 VSUBS 0.01324f
C1105 VTAIL.n414 VSUBS 0.023271f
C1106 VTAIL.n415 VSUBS 0.012505f
C1107 VTAIL.n416 VSUBS 0.022167f
C1108 VTAIL.n417 VSUBS 0.022234f
C1109 VTAIL.t6 VSUBS 0.063708f
C1110 VTAIL.n418 VSUBS 0.185376f
C1111 VTAIL.n419 VSUBS 1.16375f
C1112 VTAIL.n420 VSUBS 0.012505f
C1113 VTAIL.n421 VSUBS 0.01324f
C1114 VTAIL.n422 VSUBS 0.029556f
C1115 VTAIL.n423 VSUBS 0.029556f
C1116 VTAIL.n424 VSUBS 0.01324f
C1117 VTAIL.n425 VSUBS 0.012505f
C1118 VTAIL.n426 VSUBS 0.023271f
C1119 VTAIL.n427 VSUBS 0.023271f
C1120 VTAIL.n428 VSUBS 0.012505f
C1121 VTAIL.n429 VSUBS 0.01324f
C1122 VTAIL.n430 VSUBS 0.029556f
C1123 VTAIL.n431 VSUBS 0.029556f
C1124 VTAIL.n432 VSUBS 0.01324f
C1125 VTAIL.n433 VSUBS 0.012505f
C1126 VTAIL.n434 VSUBS 0.023271f
C1127 VTAIL.n435 VSUBS 0.023271f
C1128 VTAIL.n436 VSUBS 0.012505f
C1129 VTAIL.n437 VSUBS 0.01324f
C1130 VTAIL.n438 VSUBS 0.029556f
C1131 VTAIL.n439 VSUBS 0.029556f
C1132 VTAIL.n440 VSUBS 0.029556f
C1133 VTAIL.n441 VSUBS 0.012872f
C1134 VTAIL.n442 VSUBS 0.012505f
C1135 VTAIL.n443 VSUBS 0.023271f
C1136 VTAIL.n444 VSUBS 0.023271f
C1137 VTAIL.n445 VSUBS 0.012505f
C1138 VTAIL.n446 VSUBS 0.01324f
C1139 VTAIL.n447 VSUBS 0.029556f
C1140 VTAIL.n448 VSUBS 0.029556f
C1141 VTAIL.n449 VSUBS 0.01324f
C1142 VTAIL.n450 VSUBS 0.012505f
C1143 VTAIL.n451 VSUBS 0.023271f
C1144 VTAIL.n452 VSUBS 0.023271f
C1145 VTAIL.n453 VSUBS 0.012505f
C1146 VTAIL.n454 VSUBS 0.01324f
C1147 VTAIL.n455 VSUBS 0.029556f
C1148 VTAIL.n456 VSUBS 0.07391f
C1149 VTAIL.n457 VSUBS 0.01324f
C1150 VTAIL.n458 VSUBS 0.012505f
C1151 VTAIL.n459 VSUBS 0.056332f
C1152 VTAIL.n460 VSUBS 0.03735f
C1153 VTAIL.n461 VSUBS 1.45053f
C1154 VTAIL.n462 VSUBS 0.026261f
C1155 VTAIL.n463 VSUBS 0.023271f
C1156 VTAIL.n464 VSUBS 0.012505f
C1157 VTAIL.n465 VSUBS 0.029556f
C1158 VTAIL.n466 VSUBS 0.01324f
C1159 VTAIL.n467 VSUBS 0.023271f
C1160 VTAIL.n468 VSUBS 0.012505f
C1161 VTAIL.n469 VSUBS 0.029556f
C1162 VTAIL.n470 VSUBS 0.01324f
C1163 VTAIL.n471 VSUBS 0.023271f
C1164 VTAIL.n472 VSUBS 0.012872f
C1165 VTAIL.n473 VSUBS 0.029556f
C1166 VTAIL.n474 VSUBS 0.01324f
C1167 VTAIL.n475 VSUBS 0.023271f
C1168 VTAIL.n476 VSUBS 0.012505f
C1169 VTAIL.n477 VSUBS 0.029556f
C1170 VTAIL.n478 VSUBS 0.01324f
C1171 VTAIL.n479 VSUBS 0.023271f
C1172 VTAIL.n480 VSUBS 0.012505f
C1173 VTAIL.n481 VSUBS 0.022167f
C1174 VTAIL.n482 VSUBS 0.022234f
C1175 VTAIL.t3 VSUBS 0.063708f
C1176 VTAIL.n483 VSUBS 0.185376f
C1177 VTAIL.n484 VSUBS 1.16375f
C1178 VTAIL.n485 VSUBS 0.012505f
C1179 VTAIL.n486 VSUBS 0.01324f
C1180 VTAIL.n487 VSUBS 0.029556f
C1181 VTAIL.n488 VSUBS 0.029556f
C1182 VTAIL.n489 VSUBS 0.01324f
C1183 VTAIL.n490 VSUBS 0.012505f
C1184 VTAIL.n491 VSUBS 0.023271f
C1185 VTAIL.n492 VSUBS 0.023271f
C1186 VTAIL.n493 VSUBS 0.012505f
C1187 VTAIL.n494 VSUBS 0.01324f
C1188 VTAIL.n495 VSUBS 0.029556f
C1189 VTAIL.n496 VSUBS 0.029556f
C1190 VTAIL.n497 VSUBS 0.01324f
C1191 VTAIL.n498 VSUBS 0.012505f
C1192 VTAIL.n499 VSUBS 0.023271f
C1193 VTAIL.n500 VSUBS 0.023271f
C1194 VTAIL.n501 VSUBS 0.012505f
C1195 VTAIL.n502 VSUBS 0.012505f
C1196 VTAIL.n503 VSUBS 0.01324f
C1197 VTAIL.n504 VSUBS 0.029556f
C1198 VTAIL.n505 VSUBS 0.029556f
C1199 VTAIL.n506 VSUBS 0.029556f
C1200 VTAIL.n507 VSUBS 0.012872f
C1201 VTAIL.n508 VSUBS 0.012505f
C1202 VTAIL.n509 VSUBS 0.023271f
C1203 VTAIL.n510 VSUBS 0.023271f
C1204 VTAIL.n511 VSUBS 0.012505f
C1205 VTAIL.n512 VSUBS 0.01324f
C1206 VTAIL.n513 VSUBS 0.029556f
C1207 VTAIL.n514 VSUBS 0.029556f
C1208 VTAIL.n515 VSUBS 0.01324f
C1209 VTAIL.n516 VSUBS 0.012505f
C1210 VTAIL.n517 VSUBS 0.023271f
C1211 VTAIL.n518 VSUBS 0.023271f
C1212 VTAIL.n519 VSUBS 0.012505f
C1213 VTAIL.n520 VSUBS 0.01324f
C1214 VTAIL.n521 VSUBS 0.029556f
C1215 VTAIL.n522 VSUBS 0.07391f
C1216 VTAIL.n523 VSUBS 0.01324f
C1217 VTAIL.n524 VSUBS 0.012505f
C1218 VTAIL.n525 VSUBS 0.056332f
C1219 VTAIL.n526 VSUBS 0.03735f
C1220 VTAIL.n527 VSUBS 1.36504f
C1221 VDD1.t2 VSUBS 0.259196f
C1222 VDD1.t3 VSUBS 0.259196f
C1223 VDD1.n0 VSUBS 2.03411f
C1224 VDD1.t0 VSUBS 0.259196f
C1225 VDD1.t1 VSUBS 0.259196f
C1226 VDD1.n1 VSUBS 2.73909f
C1227 VP.n0 VSUBS 0.048813f
C1228 VP.t2 VSUBS 2.68436f
C1229 VP.n1 VSUBS 0.029905f
C1230 VP.n2 VSUBS 0.048813f
C1231 VP.t0 VSUBS 2.68436f
C1232 VP.t1 VSUBS 2.92227f
C1233 VP.t3 VSUBS 2.92657f
C1234 VP.n3 VSUBS 3.75609f
C1235 VP.n4 VSUBS 2.02291f
C1236 VP.n5 VSUBS 1.06099f
C1237 VP.n6 VSUBS 0.052053f
C1238 VP.n7 VSUBS 0.073203f
C1239 VP.n8 VSUBS 0.037027f
C1240 VP.n9 VSUBS 0.037027f
C1241 VP.n10 VSUBS 0.037027f
C1242 VP.n11 VSUBS 0.073203f
C1243 VP.n12 VSUBS 0.052053f
C1244 VP.n13 VSUBS 1.06099f
C1245 VP.n14 VSUBS 0.053398f
.ends

