* NGSPICE file created from diff_pair_sample_0295.ext - technology: sky130A

.subckt diff_pair_sample_0295 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n1910_n3148# sky130_fd_pr__pfet_01v8 ad=4.251 pd=22.58 as=0 ps=0 w=10.9 l=2.02
X1 B.t8 B.t6 B.t7 w_n1910_n3148# sky130_fd_pr__pfet_01v8 ad=4.251 pd=22.58 as=0 ps=0 w=10.9 l=2.02
X2 VDD2.t1 VN.t0 VTAIL.t3 w_n1910_n3148# sky130_fd_pr__pfet_01v8 ad=4.251 pd=22.58 as=4.251 ps=22.58 w=10.9 l=2.02
X3 B.t5 B.t3 B.t4 w_n1910_n3148# sky130_fd_pr__pfet_01v8 ad=4.251 pd=22.58 as=0 ps=0 w=10.9 l=2.02
X4 VDD2.t0 VN.t1 VTAIL.t2 w_n1910_n3148# sky130_fd_pr__pfet_01v8 ad=4.251 pd=22.58 as=4.251 ps=22.58 w=10.9 l=2.02
X5 VDD1.t1 VP.t0 VTAIL.t0 w_n1910_n3148# sky130_fd_pr__pfet_01v8 ad=4.251 pd=22.58 as=4.251 ps=22.58 w=10.9 l=2.02
X6 B.t2 B.t0 B.t1 w_n1910_n3148# sky130_fd_pr__pfet_01v8 ad=4.251 pd=22.58 as=0 ps=0 w=10.9 l=2.02
X7 VDD1.t0 VP.t1 VTAIL.t1 w_n1910_n3148# sky130_fd_pr__pfet_01v8 ad=4.251 pd=22.58 as=4.251 ps=22.58 w=10.9 l=2.02
R0 B.n371 B.n60 585
R1 B.n373 B.n372 585
R2 B.n374 B.n59 585
R3 B.n376 B.n375 585
R4 B.n377 B.n58 585
R5 B.n379 B.n378 585
R6 B.n380 B.n57 585
R7 B.n382 B.n381 585
R8 B.n383 B.n56 585
R9 B.n385 B.n384 585
R10 B.n386 B.n55 585
R11 B.n388 B.n387 585
R12 B.n389 B.n54 585
R13 B.n391 B.n390 585
R14 B.n392 B.n53 585
R15 B.n394 B.n393 585
R16 B.n395 B.n52 585
R17 B.n397 B.n396 585
R18 B.n398 B.n51 585
R19 B.n400 B.n399 585
R20 B.n401 B.n50 585
R21 B.n403 B.n402 585
R22 B.n404 B.n49 585
R23 B.n406 B.n405 585
R24 B.n407 B.n48 585
R25 B.n409 B.n408 585
R26 B.n410 B.n47 585
R27 B.n412 B.n411 585
R28 B.n413 B.n46 585
R29 B.n415 B.n414 585
R30 B.n416 B.n45 585
R31 B.n418 B.n417 585
R32 B.n419 B.n44 585
R33 B.n421 B.n420 585
R34 B.n422 B.n43 585
R35 B.n424 B.n423 585
R36 B.n425 B.n42 585
R37 B.n427 B.n426 585
R38 B.n429 B.n39 585
R39 B.n431 B.n430 585
R40 B.n432 B.n38 585
R41 B.n434 B.n433 585
R42 B.n435 B.n37 585
R43 B.n437 B.n436 585
R44 B.n438 B.n36 585
R45 B.n440 B.n439 585
R46 B.n441 B.n35 585
R47 B.n443 B.n442 585
R48 B.n445 B.n444 585
R49 B.n446 B.n31 585
R50 B.n448 B.n447 585
R51 B.n449 B.n30 585
R52 B.n451 B.n450 585
R53 B.n452 B.n29 585
R54 B.n454 B.n453 585
R55 B.n455 B.n28 585
R56 B.n457 B.n456 585
R57 B.n458 B.n27 585
R58 B.n460 B.n459 585
R59 B.n461 B.n26 585
R60 B.n463 B.n462 585
R61 B.n464 B.n25 585
R62 B.n466 B.n465 585
R63 B.n467 B.n24 585
R64 B.n469 B.n468 585
R65 B.n470 B.n23 585
R66 B.n472 B.n471 585
R67 B.n473 B.n22 585
R68 B.n475 B.n474 585
R69 B.n476 B.n21 585
R70 B.n478 B.n477 585
R71 B.n479 B.n20 585
R72 B.n481 B.n480 585
R73 B.n482 B.n19 585
R74 B.n484 B.n483 585
R75 B.n485 B.n18 585
R76 B.n487 B.n486 585
R77 B.n488 B.n17 585
R78 B.n490 B.n489 585
R79 B.n491 B.n16 585
R80 B.n493 B.n492 585
R81 B.n494 B.n15 585
R82 B.n496 B.n495 585
R83 B.n497 B.n14 585
R84 B.n499 B.n498 585
R85 B.n500 B.n13 585
R86 B.n370 B.n369 585
R87 B.n368 B.n61 585
R88 B.n367 B.n366 585
R89 B.n365 B.n62 585
R90 B.n364 B.n363 585
R91 B.n362 B.n63 585
R92 B.n361 B.n360 585
R93 B.n359 B.n64 585
R94 B.n358 B.n357 585
R95 B.n356 B.n65 585
R96 B.n355 B.n354 585
R97 B.n353 B.n66 585
R98 B.n352 B.n351 585
R99 B.n350 B.n67 585
R100 B.n349 B.n348 585
R101 B.n347 B.n68 585
R102 B.n346 B.n345 585
R103 B.n344 B.n69 585
R104 B.n343 B.n342 585
R105 B.n341 B.n70 585
R106 B.n340 B.n339 585
R107 B.n338 B.n71 585
R108 B.n337 B.n336 585
R109 B.n335 B.n72 585
R110 B.n334 B.n333 585
R111 B.n332 B.n73 585
R112 B.n331 B.n330 585
R113 B.n329 B.n74 585
R114 B.n328 B.n327 585
R115 B.n326 B.n75 585
R116 B.n325 B.n324 585
R117 B.n323 B.n76 585
R118 B.n322 B.n321 585
R119 B.n320 B.n77 585
R120 B.n319 B.n318 585
R121 B.n317 B.n78 585
R122 B.n316 B.n315 585
R123 B.n314 B.n79 585
R124 B.n313 B.n312 585
R125 B.n311 B.n80 585
R126 B.n310 B.n309 585
R127 B.n308 B.n81 585
R128 B.n307 B.n306 585
R129 B.n305 B.n82 585
R130 B.n304 B.n303 585
R131 B.n173 B.n130 585
R132 B.n175 B.n174 585
R133 B.n176 B.n129 585
R134 B.n178 B.n177 585
R135 B.n179 B.n128 585
R136 B.n181 B.n180 585
R137 B.n182 B.n127 585
R138 B.n184 B.n183 585
R139 B.n185 B.n126 585
R140 B.n187 B.n186 585
R141 B.n188 B.n125 585
R142 B.n190 B.n189 585
R143 B.n191 B.n124 585
R144 B.n193 B.n192 585
R145 B.n194 B.n123 585
R146 B.n196 B.n195 585
R147 B.n197 B.n122 585
R148 B.n199 B.n198 585
R149 B.n200 B.n121 585
R150 B.n202 B.n201 585
R151 B.n203 B.n120 585
R152 B.n205 B.n204 585
R153 B.n206 B.n119 585
R154 B.n208 B.n207 585
R155 B.n209 B.n118 585
R156 B.n211 B.n210 585
R157 B.n212 B.n117 585
R158 B.n214 B.n213 585
R159 B.n215 B.n116 585
R160 B.n217 B.n216 585
R161 B.n218 B.n115 585
R162 B.n220 B.n219 585
R163 B.n221 B.n114 585
R164 B.n223 B.n222 585
R165 B.n224 B.n113 585
R166 B.n226 B.n225 585
R167 B.n227 B.n112 585
R168 B.n229 B.n228 585
R169 B.n231 B.n109 585
R170 B.n233 B.n232 585
R171 B.n234 B.n108 585
R172 B.n236 B.n235 585
R173 B.n237 B.n107 585
R174 B.n239 B.n238 585
R175 B.n240 B.n106 585
R176 B.n242 B.n241 585
R177 B.n243 B.n105 585
R178 B.n245 B.n244 585
R179 B.n247 B.n246 585
R180 B.n248 B.n101 585
R181 B.n250 B.n249 585
R182 B.n251 B.n100 585
R183 B.n253 B.n252 585
R184 B.n254 B.n99 585
R185 B.n256 B.n255 585
R186 B.n257 B.n98 585
R187 B.n259 B.n258 585
R188 B.n260 B.n97 585
R189 B.n262 B.n261 585
R190 B.n263 B.n96 585
R191 B.n265 B.n264 585
R192 B.n266 B.n95 585
R193 B.n268 B.n267 585
R194 B.n269 B.n94 585
R195 B.n271 B.n270 585
R196 B.n272 B.n93 585
R197 B.n274 B.n273 585
R198 B.n275 B.n92 585
R199 B.n277 B.n276 585
R200 B.n278 B.n91 585
R201 B.n280 B.n279 585
R202 B.n281 B.n90 585
R203 B.n283 B.n282 585
R204 B.n284 B.n89 585
R205 B.n286 B.n285 585
R206 B.n287 B.n88 585
R207 B.n289 B.n288 585
R208 B.n290 B.n87 585
R209 B.n292 B.n291 585
R210 B.n293 B.n86 585
R211 B.n295 B.n294 585
R212 B.n296 B.n85 585
R213 B.n298 B.n297 585
R214 B.n299 B.n84 585
R215 B.n301 B.n300 585
R216 B.n302 B.n83 585
R217 B.n172 B.n171 585
R218 B.n170 B.n131 585
R219 B.n169 B.n168 585
R220 B.n167 B.n132 585
R221 B.n166 B.n165 585
R222 B.n164 B.n133 585
R223 B.n163 B.n162 585
R224 B.n161 B.n134 585
R225 B.n160 B.n159 585
R226 B.n158 B.n135 585
R227 B.n157 B.n156 585
R228 B.n155 B.n136 585
R229 B.n154 B.n153 585
R230 B.n152 B.n137 585
R231 B.n151 B.n150 585
R232 B.n149 B.n138 585
R233 B.n148 B.n147 585
R234 B.n146 B.n139 585
R235 B.n145 B.n144 585
R236 B.n143 B.n140 585
R237 B.n142 B.n141 585
R238 B.n2 B.n0 585
R239 B.n533 B.n1 585
R240 B.n532 B.n531 585
R241 B.n530 B.n3 585
R242 B.n529 B.n528 585
R243 B.n527 B.n4 585
R244 B.n526 B.n525 585
R245 B.n524 B.n5 585
R246 B.n523 B.n522 585
R247 B.n521 B.n6 585
R248 B.n520 B.n519 585
R249 B.n518 B.n7 585
R250 B.n517 B.n516 585
R251 B.n515 B.n8 585
R252 B.n514 B.n513 585
R253 B.n512 B.n9 585
R254 B.n511 B.n510 585
R255 B.n509 B.n10 585
R256 B.n508 B.n507 585
R257 B.n506 B.n11 585
R258 B.n505 B.n504 585
R259 B.n503 B.n12 585
R260 B.n502 B.n501 585
R261 B.n535 B.n534 585
R262 B.n173 B.n172 516.524
R263 B.n502 B.n13 516.524
R264 B.n304 B.n83 516.524
R265 B.n371 B.n370 516.524
R266 B.n102 B.t9 337.009
R267 B.n110 B.t6 337.009
R268 B.n32 B.t3 337.009
R269 B.n40 B.t0 337.009
R270 B.n172 B.n131 163.367
R271 B.n168 B.n131 163.367
R272 B.n168 B.n167 163.367
R273 B.n167 B.n166 163.367
R274 B.n166 B.n133 163.367
R275 B.n162 B.n133 163.367
R276 B.n162 B.n161 163.367
R277 B.n161 B.n160 163.367
R278 B.n160 B.n135 163.367
R279 B.n156 B.n135 163.367
R280 B.n156 B.n155 163.367
R281 B.n155 B.n154 163.367
R282 B.n154 B.n137 163.367
R283 B.n150 B.n137 163.367
R284 B.n150 B.n149 163.367
R285 B.n149 B.n148 163.367
R286 B.n148 B.n139 163.367
R287 B.n144 B.n139 163.367
R288 B.n144 B.n143 163.367
R289 B.n143 B.n142 163.367
R290 B.n142 B.n2 163.367
R291 B.n534 B.n2 163.367
R292 B.n534 B.n533 163.367
R293 B.n533 B.n532 163.367
R294 B.n532 B.n3 163.367
R295 B.n528 B.n3 163.367
R296 B.n528 B.n527 163.367
R297 B.n527 B.n526 163.367
R298 B.n526 B.n5 163.367
R299 B.n522 B.n5 163.367
R300 B.n522 B.n521 163.367
R301 B.n521 B.n520 163.367
R302 B.n520 B.n7 163.367
R303 B.n516 B.n7 163.367
R304 B.n516 B.n515 163.367
R305 B.n515 B.n514 163.367
R306 B.n514 B.n9 163.367
R307 B.n510 B.n9 163.367
R308 B.n510 B.n509 163.367
R309 B.n509 B.n508 163.367
R310 B.n508 B.n11 163.367
R311 B.n504 B.n11 163.367
R312 B.n504 B.n503 163.367
R313 B.n503 B.n502 163.367
R314 B.n174 B.n173 163.367
R315 B.n174 B.n129 163.367
R316 B.n178 B.n129 163.367
R317 B.n179 B.n178 163.367
R318 B.n180 B.n179 163.367
R319 B.n180 B.n127 163.367
R320 B.n184 B.n127 163.367
R321 B.n185 B.n184 163.367
R322 B.n186 B.n185 163.367
R323 B.n186 B.n125 163.367
R324 B.n190 B.n125 163.367
R325 B.n191 B.n190 163.367
R326 B.n192 B.n191 163.367
R327 B.n192 B.n123 163.367
R328 B.n196 B.n123 163.367
R329 B.n197 B.n196 163.367
R330 B.n198 B.n197 163.367
R331 B.n198 B.n121 163.367
R332 B.n202 B.n121 163.367
R333 B.n203 B.n202 163.367
R334 B.n204 B.n203 163.367
R335 B.n204 B.n119 163.367
R336 B.n208 B.n119 163.367
R337 B.n209 B.n208 163.367
R338 B.n210 B.n209 163.367
R339 B.n210 B.n117 163.367
R340 B.n214 B.n117 163.367
R341 B.n215 B.n214 163.367
R342 B.n216 B.n215 163.367
R343 B.n216 B.n115 163.367
R344 B.n220 B.n115 163.367
R345 B.n221 B.n220 163.367
R346 B.n222 B.n221 163.367
R347 B.n222 B.n113 163.367
R348 B.n226 B.n113 163.367
R349 B.n227 B.n226 163.367
R350 B.n228 B.n227 163.367
R351 B.n228 B.n109 163.367
R352 B.n233 B.n109 163.367
R353 B.n234 B.n233 163.367
R354 B.n235 B.n234 163.367
R355 B.n235 B.n107 163.367
R356 B.n239 B.n107 163.367
R357 B.n240 B.n239 163.367
R358 B.n241 B.n240 163.367
R359 B.n241 B.n105 163.367
R360 B.n245 B.n105 163.367
R361 B.n246 B.n245 163.367
R362 B.n246 B.n101 163.367
R363 B.n250 B.n101 163.367
R364 B.n251 B.n250 163.367
R365 B.n252 B.n251 163.367
R366 B.n252 B.n99 163.367
R367 B.n256 B.n99 163.367
R368 B.n257 B.n256 163.367
R369 B.n258 B.n257 163.367
R370 B.n258 B.n97 163.367
R371 B.n262 B.n97 163.367
R372 B.n263 B.n262 163.367
R373 B.n264 B.n263 163.367
R374 B.n264 B.n95 163.367
R375 B.n268 B.n95 163.367
R376 B.n269 B.n268 163.367
R377 B.n270 B.n269 163.367
R378 B.n270 B.n93 163.367
R379 B.n274 B.n93 163.367
R380 B.n275 B.n274 163.367
R381 B.n276 B.n275 163.367
R382 B.n276 B.n91 163.367
R383 B.n280 B.n91 163.367
R384 B.n281 B.n280 163.367
R385 B.n282 B.n281 163.367
R386 B.n282 B.n89 163.367
R387 B.n286 B.n89 163.367
R388 B.n287 B.n286 163.367
R389 B.n288 B.n287 163.367
R390 B.n288 B.n87 163.367
R391 B.n292 B.n87 163.367
R392 B.n293 B.n292 163.367
R393 B.n294 B.n293 163.367
R394 B.n294 B.n85 163.367
R395 B.n298 B.n85 163.367
R396 B.n299 B.n298 163.367
R397 B.n300 B.n299 163.367
R398 B.n300 B.n83 163.367
R399 B.n305 B.n304 163.367
R400 B.n306 B.n305 163.367
R401 B.n306 B.n81 163.367
R402 B.n310 B.n81 163.367
R403 B.n311 B.n310 163.367
R404 B.n312 B.n311 163.367
R405 B.n312 B.n79 163.367
R406 B.n316 B.n79 163.367
R407 B.n317 B.n316 163.367
R408 B.n318 B.n317 163.367
R409 B.n318 B.n77 163.367
R410 B.n322 B.n77 163.367
R411 B.n323 B.n322 163.367
R412 B.n324 B.n323 163.367
R413 B.n324 B.n75 163.367
R414 B.n328 B.n75 163.367
R415 B.n329 B.n328 163.367
R416 B.n330 B.n329 163.367
R417 B.n330 B.n73 163.367
R418 B.n334 B.n73 163.367
R419 B.n335 B.n334 163.367
R420 B.n336 B.n335 163.367
R421 B.n336 B.n71 163.367
R422 B.n340 B.n71 163.367
R423 B.n341 B.n340 163.367
R424 B.n342 B.n341 163.367
R425 B.n342 B.n69 163.367
R426 B.n346 B.n69 163.367
R427 B.n347 B.n346 163.367
R428 B.n348 B.n347 163.367
R429 B.n348 B.n67 163.367
R430 B.n352 B.n67 163.367
R431 B.n353 B.n352 163.367
R432 B.n354 B.n353 163.367
R433 B.n354 B.n65 163.367
R434 B.n358 B.n65 163.367
R435 B.n359 B.n358 163.367
R436 B.n360 B.n359 163.367
R437 B.n360 B.n63 163.367
R438 B.n364 B.n63 163.367
R439 B.n365 B.n364 163.367
R440 B.n366 B.n365 163.367
R441 B.n366 B.n61 163.367
R442 B.n370 B.n61 163.367
R443 B.n498 B.n13 163.367
R444 B.n498 B.n497 163.367
R445 B.n497 B.n496 163.367
R446 B.n496 B.n15 163.367
R447 B.n492 B.n15 163.367
R448 B.n492 B.n491 163.367
R449 B.n491 B.n490 163.367
R450 B.n490 B.n17 163.367
R451 B.n486 B.n17 163.367
R452 B.n486 B.n485 163.367
R453 B.n485 B.n484 163.367
R454 B.n484 B.n19 163.367
R455 B.n480 B.n19 163.367
R456 B.n480 B.n479 163.367
R457 B.n479 B.n478 163.367
R458 B.n478 B.n21 163.367
R459 B.n474 B.n21 163.367
R460 B.n474 B.n473 163.367
R461 B.n473 B.n472 163.367
R462 B.n472 B.n23 163.367
R463 B.n468 B.n23 163.367
R464 B.n468 B.n467 163.367
R465 B.n467 B.n466 163.367
R466 B.n466 B.n25 163.367
R467 B.n462 B.n25 163.367
R468 B.n462 B.n461 163.367
R469 B.n461 B.n460 163.367
R470 B.n460 B.n27 163.367
R471 B.n456 B.n27 163.367
R472 B.n456 B.n455 163.367
R473 B.n455 B.n454 163.367
R474 B.n454 B.n29 163.367
R475 B.n450 B.n29 163.367
R476 B.n450 B.n449 163.367
R477 B.n449 B.n448 163.367
R478 B.n448 B.n31 163.367
R479 B.n444 B.n31 163.367
R480 B.n444 B.n443 163.367
R481 B.n443 B.n35 163.367
R482 B.n439 B.n35 163.367
R483 B.n439 B.n438 163.367
R484 B.n438 B.n437 163.367
R485 B.n437 B.n37 163.367
R486 B.n433 B.n37 163.367
R487 B.n433 B.n432 163.367
R488 B.n432 B.n431 163.367
R489 B.n431 B.n39 163.367
R490 B.n426 B.n39 163.367
R491 B.n426 B.n425 163.367
R492 B.n425 B.n424 163.367
R493 B.n424 B.n43 163.367
R494 B.n420 B.n43 163.367
R495 B.n420 B.n419 163.367
R496 B.n419 B.n418 163.367
R497 B.n418 B.n45 163.367
R498 B.n414 B.n45 163.367
R499 B.n414 B.n413 163.367
R500 B.n413 B.n412 163.367
R501 B.n412 B.n47 163.367
R502 B.n408 B.n47 163.367
R503 B.n408 B.n407 163.367
R504 B.n407 B.n406 163.367
R505 B.n406 B.n49 163.367
R506 B.n402 B.n49 163.367
R507 B.n402 B.n401 163.367
R508 B.n401 B.n400 163.367
R509 B.n400 B.n51 163.367
R510 B.n396 B.n51 163.367
R511 B.n396 B.n395 163.367
R512 B.n395 B.n394 163.367
R513 B.n394 B.n53 163.367
R514 B.n390 B.n53 163.367
R515 B.n390 B.n389 163.367
R516 B.n389 B.n388 163.367
R517 B.n388 B.n55 163.367
R518 B.n384 B.n55 163.367
R519 B.n384 B.n383 163.367
R520 B.n383 B.n382 163.367
R521 B.n382 B.n57 163.367
R522 B.n378 B.n57 163.367
R523 B.n378 B.n377 163.367
R524 B.n377 B.n376 163.367
R525 B.n376 B.n59 163.367
R526 B.n372 B.n59 163.367
R527 B.n372 B.n371 163.367
R528 B.n102 B.t11 153.35
R529 B.n40 B.t1 153.35
R530 B.n110 B.t8 153.337
R531 B.n32 B.t4 153.337
R532 B.n103 B.t10 107.775
R533 B.n41 B.t2 107.775
R534 B.n111 B.t7 107.761
R535 B.n33 B.t5 107.761
R536 B.n104 B.n103 59.5399
R537 B.n230 B.n111 59.5399
R538 B.n34 B.n33 59.5399
R539 B.n428 B.n41 59.5399
R540 B.n103 B.n102 45.5763
R541 B.n111 B.n110 45.5763
R542 B.n33 B.n32 45.5763
R543 B.n41 B.n40 45.5763
R544 B.n501 B.n500 33.5615
R545 B.n369 B.n60 33.5615
R546 B.n303 B.n302 33.5615
R547 B.n171 B.n130 33.5615
R548 B B.n535 18.0485
R549 B.n500 B.n499 10.6151
R550 B.n499 B.n14 10.6151
R551 B.n495 B.n14 10.6151
R552 B.n495 B.n494 10.6151
R553 B.n494 B.n493 10.6151
R554 B.n493 B.n16 10.6151
R555 B.n489 B.n16 10.6151
R556 B.n489 B.n488 10.6151
R557 B.n488 B.n487 10.6151
R558 B.n487 B.n18 10.6151
R559 B.n483 B.n18 10.6151
R560 B.n483 B.n482 10.6151
R561 B.n482 B.n481 10.6151
R562 B.n481 B.n20 10.6151
R563 B.n477 B.n20 10.6151
R564 B.n477 B.n476 10.6151
R565 B.n476 B.n475 10.6151
R566 B.n475 B.n22 10.6151
R567 B.n471 B.n22 10.6151
R568 B.n471 B.n470 10.6151
R569 B.n470 B.n469 10.6151
R570 B.n469 B.n24 10.6151
R571 B.n465 B.n24 10.6151
R572 B.n465 B.n464 10.6151
R573 B.n464 B.n463 10.6151
R574 B.n463 B.n26 10.6151
R575 B.n459 B.n26 10.6151
R576 B.n459 B.n458 10.6151
R577 B.n458 B.n457 10.6151
R578 B.n457 B.n28 10.6151
R579 B.n453 B.n28 10.6151
R580 B.n453 B.n452 10.6151
R581 B.n452 B.n451 10.6151
R582 B.n451 B.n30 10.6151
R583 B.n447 B.n30 10.6151
R584 B.n447 B.n446 10.6151
R585 B.n446 B.n445 10.6151
R586 B.n442 B.n441 10.6151
R587 B.n441 B.n440 10.6151
R588 B.n440 B.n36 10.6151
R589 B.n436 B.n36 10.6151
R590 B.n436 B.n435 10.6151
R591 B.n435 B.n434 10.6151
R592 B.n434 B.n38 10.6151
R593 B.n430 B.n38 10.6151
R594 B.n430 B.n429 10.6151
R595 B.n427 B.n42 10.6151
R596 B.n423 B.n42 10.6151
R597 B.n423 B.n422 10.6151
R598 B.n422 B.n421 10.6151
R599 B.n421 B.n44 10.6151
R600 B.n417 B.n44 10.6151
R601 B.n417 B.n416 10.6151
R602 B.n416 B.n415 10.6151
R603 B.n415 B.n46 10.6151
R604 B.n411 B.n46 10.6151
R605 B.n411 B.n410 10.6151
R606 B.n410 B.n409 10.6151
R607 B.n409 B.n48 10.6151
R608 B.n405 B.n48 10.6151
R609 B.n405 B.n404 10.6151
R610 B.n404 B.n403 10.6151
R611 B.n403 B.n50 10.6151
R612 B.n399 B.n50 10.6151
R613 B.n399 B.n398 10.6151
R614 B.n398 B.n397 10.6151
R615 B.n397 B.n52 10.6151
R616 B.n393 B.n52 10.6151
R617 B.n393 B.n392 10.6151
R618 B.n392 B.n391 10.6151
R619 B.n391 B.n54 10.6151
R620 B.n387 B.n54 10.6151
R621 B.n387 B.n386 10.6151
R622 B.n386 B.n385 10.6151
R623 B.n385 B.n56 10.6151
R624 B.n381 B.n56 10.6151
R625 B.n381 B.n380 10.6151
R626 B.n380 B.n379 10.6151
R627 B.n379 B.n58 10.6151
R628 B.n375 B.n58 10.6151
R629 B.n375 B.n374 10.6151
R630 B.n374 B.n373 10.6151
R631 B.n373 B.n60 10.6151
R632 B.n303 B.n82 10.6151
R633 B.n307 B.n82 10.6151
R634 B.n308 B.n307 10.6151
R635 B.n309 B.n308 10.6151
R636 B.n309 B.n80 10.6151
R637 B.n313 B.n80 10.6151
R638 B.n314 B.n313 10.6151
R639 B.n315 B.n314 10.6151
R640 B.n315 B.n78 10.6151
R641 B.n319 B.n78 10.6151
R642 B.n320 B.n319 10.6151
R643 B.n321 B.n320 10.6151
R644 B.n321 B.n76 10.6151
R645 B.n325 B.n76 10.6151
R646 B.n326 B.n325 10.6151
R647 B.n327 B.n326 10.6151
R648 B.n327 B.n74 10.6151
R649 B.n331 B.n74 10.6151
R650 B.n332 B.n331 10.6151
R651 B.n333 B.n332 10.6151
R652 B.n333 B.n72 10.6151
R653 B.n337 B.n72 10.6151
R654 B.n338 B.n337 10.6151
R655 B.n339 B.n338 10.6151
R656 B.n339 B.n70 10.6151
R657 B.n343 B.n70 10.6151
R658 B.n344 B.n343 10.6151
R659 B.n345 B.n344 10.6151
R660 B.n345 B.n68 10.6151
R661 B.n349 B.n68 10.6151
R662 B.n350 B.n349 10.6151
R663 B.n351 B.n350 10.6151
R664 B.n351 B.n66 10.6151
R665 B.n355 B.n66 10.6151
R666 B.n356 B.n355 10.6151
R667 B.n357 B.n356 10.6151
R668 B.n357 B.n64 10.6151
R669 B.n361 B.n64 10.6151
R670 B.n362 B.n361 10.6151
R671 B.n363 B.n362 10.6151
R672 B.n363 B.n62 10.6151
R673 B.n367 B.n62 10.6151
R674 B.n368 B.n367 10.6151
R675 B.n369 B.n368 10.6151
R676 B.n175 B.n130 10.6151
R677 B.n176 B.n175 10.6151
R678 B.n177 B.n176 10.6151
R679 B.n177 B.n128 10.6151
R680 B.n181 B.n128 10.6151
R681 B.n182 B.n181 10.6151
R682 B.n183 B.n182 10.6151
R683 B.n183 B.n126 10.6151
R684 B.n187 B.n126 10.6151
R685 B.n188 B.n187 10.6151
R686 B.n189 B.n188 10.6151
R687 B.n189 B.n124 10.6151
R688 B.n193 B.n124 10.6151
R689 B.n194 B.n193 10.6151
R690 B.n195 B.n194 10.6151
R691 B.n195 B.n122 10.6151
R692 B.n199 B.n122 10.6151
R693 B.n200 B.n199 10.6151
R694 B.n201 B.n200 10.6151
R695 B.n201 B.n120 10.6151
R696 B.n205 B.n120 10.6151
R697 B.n206 B.n205 10.6151
R698 B.n207 B.n206 10.6151
R699 B.n207 B.n118 10.6151
R700 B.n211 B.n118 10.6151
R701 B.n212 B.n211 10.6151
R702 B.n213 B.n212 10.6151
R703 B.n213 B.n116 10.6151
R704 B.n217 B.n116 10.6151
R705 B.n218 B.n217 10.6151
R706 B.n219 B.n218 10.6151
R707 B.n219 B.n114 10.6151
R708 B.n223 B.n114 10.6151
R709 B.n224 B.n223 10.6151
R710 B.n225 B.n224 10.6151
R711 B.n225 B.n112 10.6151
R712 B.n229 B.n112 10.6151
R713 B.n232 B.n231 10.6151
R714 B.n232 B.n108 10.6151
R715 B.n236 B.n108 10.6151
R716 B.n237 B.n236 10.6151
R717 B.n238 B.n237 10.6151
R718 B.n238 B.n106 10.6151
R719 B.n242 B.n106 10.6151
R720 B.n243 B.n242 10.6151
R721 B.n244 B.n243 10.6151
R722 B.n248 B.n247 10.6151
R723 B.n249 B.n248 10.6151
R724 B.n249 B.n100 10.6151
R725 B.n253 B.n100 10.6151
R726 B.n254 B.n253 10.6151
R727 B.n255 B.n254 10.6151
R728 B.n255 B.n98 10.6151
R729 B.n259 B.n98 10.6151
R730 B.n260 B.n259 10.6151
R731 B.n261 B.n260 10.6151
R732 B.n261 B.n96 10.6151
R733 B.n265 B.n96 10.6151
R734 B.n266 B.n265 10.6151
R735 B.n267 B.n266 10.6151
R736 B.n267 B.n94 10.6151
R737 B.n271 B.n94 10.6151
R738 B.n272 B.n271 10.6151
R739 B.n273 B.n272 10.6151
R740 B.n273 B.n92 10.6151
R741 B.n277 B.n92 10.6151
R742 B.n278 B.n277 10.6151
R743 B.n279 B.n278 10.6151
R744 B.n279 B.n90 10.6151
R745 B.n283 B.n90 10.6151
R746 B.n284 B.n283 10.6151
R747 B.n285 B.n284 10.6151
R748 B.n285 B.n88 10.6151
R749 B.n289 B.n88 10.6151
R750 B.n290 B.n289 10.6151
R751 B.n291 B.n290 10.6151
R752 B.n291 B.n86 10.6151
R753 B.n295 B.n86 10.6151
R754 B.n296 B.n295 10.6151
R755 B.n297 B.n296 10.6151
R756 B.n297 B.n84 10.6151
R757 B.n301 B.n84 10.6151
R758 B.n302 B.n301 10.6151
R759 B.n171 B.n170 10.6151
R760 B.n170 B.n169 10.6151
R761 B.n169 B.n132 10.6151
R762 B.n165 B.n132 10.6151
R763 B.n165 B.n164 10.6151
R764 B.n164 B.n163 10.6151
R765 B.n163 B.n134 10.6151
R766 B.n159 B.n134 10.6151
R767 B.n159 B.n158 10.6151
R768 B.n158 B.n157 10.6151
R769 B.n157 B.n136 10.6151
R770 B.n153 B.n136 10.6151
R771 B.n153 B.n152 10.6151
R772 B.n152 B.n151 10.6151
R773 B.n151 B.n138 10.6151
R774 B.n147 B.n138 10.6151
R775 B.n147 B.n146 10.6151
R776 B.n146 B.n145 10.6151
R777 B.n145 B.n140 10.6151
R778 B.n141 B.n140 10.6151
R779 B.n141 B.n0 10.6151
R780 B.n531 B.n1 10.6151
R781 B.n531 B.n530 10.6151
R782 B.n530 B.n529 10.6151
R783 B.n529 B.n4 10.6151
R784 B.n525 B.n4 10.6151
R785 B.n525 B.n524 10.6151
R786 B.n524 B.n523 10.6151
R787 B.n523 B.n6 10.6151
R788 B.n519 B.n6 10.6151
R789 B.n519 B.n518 10.6151
R790 B.n518 B.n517 10.6151
R791 B.n517 B.n8 10.6151
R792 B.n513 B.n8 10.6151
R793 B.n513 B.n512 10.6151
R794 B.n512 B.n511 10.6151
R795 B.n511 B.n10 10.6151
R796 B.n507 B.n10 10.6151
R797 B.n507 B.n506 10.6151
R798 B.n506 B.n505 10.6151
R799 B.n505 B.n12 10.6151
R800 B.n501 B.n12 10.6151
R801 B.n445 B.n34 9.36635
R802 B.n428 B.n427 9.36635
R803 B.n230 B.n229 9.36635
R804 B.n247 B.n104 9.36635
R805 B.n535 B.n0 2.81026
R806 B.n535 B.n1 2.81026
R807 B.n442 B.n34 1.24928
R808 B.n429 B.n428 1.24928
R809 B.n231 B.n230 1.24928
R810 B.n244 B.n104 1.24928
R811 VN VN.t0 231.357
R812 VN VN.t1 189.123
R813 VTAIL.n1 VTAIL.t3 65.3354
R814 VTAIL.n3 VTAIL.t2 65.3344
R815 VTAIL.n0 VTAIL.t1 65.3344
R816 VTAIL.n2 VTAIL.t0 65.3342
R817 VTAIL.n1 VTAIL.n0 25.8152
R818 VTAIL.n3 VTAIL.n2 23.7893
R819 VTAIL.n2 VTAIL.n1 1.48326
R820 VTAIL VTAIL.n0 1.03498
R821 VTAIL VTAIL.n3 0.448776
R822 VDD2.n0 VDD2.t0 119.121
R823 VDD2.n0 VDD2.t1 82.013
R824 VDD2 VDD2.n0 0.565155
R825 VP.n0 VP.t0 231.166
R826 VP.n0 VP.t1 188.881
R827 VP VP.n0 0.241678
R828 VDD1 VDD1.t0 120.153
R829 VDD1 VDD1.t1 82.5776
C0 VTAIL w_n1910_n3148# 2.61467f
C1 B VN 0.935703f
C2 VTAIL VDD2 4.76036f
C3 VTAIL VDD1 4.71405f
C4 VP VTAIL 2.12386f
C5 VDD2 w_n1910_n3148# 1.658f
C6 VDD1 w_n1910_n3148# 1.63906f
C7 VP w_n1910_n3148# 2.8068f
C8 VDD2 VDD1 0.605524f
C9 VP VDD2 0.308307f
C10 VP VDD1 2.59905f
C11 VTAIL VN 2.10953f
C12 VN w_n1910_n3148# 2.56476f
C13 VTAIL B 3.17435f
C14 B w_n1910_n3148# 7.874411f
C15 VN VDD2 2.44092f
C16 VN VDD1 0.147522f
C17 VP VN 4.98004f
C18 B VDD2 1.5651f
C19 B VDD1 1.54016f
C20 VP B 1.33131f
C21 VDD2 VSUBS 0.807239f
C22 VDD1 VSUBS 4.165875f
C23 VTAIL VSUBS 0.893161f
C24 VN VSUBS 7.470251f
C25 VP VSUBS 1.474222f
C26 B VSUBS 3.368532f
C27 w_n1910_n3148# VSUBS 74.1462f
C28 VDD1.t1 VSUBS 1.78405f
C29 VDD1.t0 VSUBS 2.28417f
C30 VP.t0 VSUBS 3.78759f
C31 VP.t1 VSUBS 3.24081f
C32 VP.n0 VSUBS 5.39098f
C33 VDD2.t0 VSUBS 2.24752f
C34 VDD2.t1 VSUBS 1.77477f
C35 VDD2.n0 VSUBS 3.0741f
C36 VTAIL.t1 VSUBS 2.43305f
C37 VTAIL.n0 VSUBS 2.49568f
C38 VTAIL.t3 VSUBS 2.43306f
C39 VTAIL.n1 VSUBS 2.53834f
C40 VTAIL.t0 VSUBS 2.43304f
C41 VTAIL.n2 VSUBS 2.34556f
C42 VTAIL.t2 VSUBS 2.43305f
C43 VTAIL.n3 VSUBS 2.24711f
C44 VN.t1 VSUBS 3.12172f
C45 VN.t0 VSUBS 3.65275f
C46 B.n0 VSUBS 0.004187f
C47 B.n1 VSUBS 0.004187f
C48 B.n2 VSUBS 0.006622f
C49 B.n3 VSUBS 0.006622f
C50 B.n4 VSUBS 0.006622f
C51 B.n5 VSUBS 0.006622f
C52 B.n6 VSUBS 0.006622f
C53 B.n7 VSUBS 0.006622f
C54 B.n8 VSUBS 0.006622f
C55 B.n9 VSUBS 0.006622f
C56 B.n10 VSUBS 0.006622f
C57 B.n11 VSUBS 0.006622f
C58 B.n12 VSUBS 0.006622f
C59 B.n13 VSUBS 0.015989f
C60 B.n14 VSUBS 0.006622f
C61 B.n15 VSUBS 0.006622f
C62 B.n16 VSUBS 0.006622f
C63 B.n17 VSUBS 0.006622f
C64 B.n18 VSUBS 0.006622f
C65 B.n19 VSUBS 0.006622f
C66 B.n20 VSUBS 0.006622f
C67 B.n21 VSUBS 0.006622f
C68 B.n22 VSUBS 0.006622f
C69 B.n23 VSUBS 0.006622f
C70 B.n24 VSUBS 0.006622f
C71 B.n25 VSUBS 0.006622f
C72 B.n26 VSUBS 0.006622f
C73 B.n27 VSUBS 0.006622f
C74 B.n28 VSUBS 0.006622f
C75 B.n29 VSUBS 0.006622f
C76 B.n30 VSUBS 0.006622f
C77 B.n31 VSUBS 0.006622f
C78 B.t5 VSUBS 0.332377f
C79 B.t4 VSUBS 0.349061f
C80 B.t3 VSUBS 0.937812f
C81 B.n32 VSUBS 0.171117f
C82 B.n33 VSUBS 0.065574f
C83 B.n34 VSUBS 0.015342f
C84 B.n35 VSUBS 0.006622f
C85 B.n36 VSUBS 0.006622f
C86 B.n37 VSUBS 0.006622f
C87 B.n38 VSUBS 0.006622f
C88 B.n39 VSUBS 0.006622f
C89 B.t2 VSUBS 0.332372f
C90 B.t1 VSUBS 0.349055f
C91 B.t0 VSUBS 0.937812f
C92 B.n40 VSUBS 0.171122f
C93 B.n41 VSUBS 0.06558f
C94 B.n42 VSUBS 0.006622f
C95 B.n43 VSUBS 0.006622f
C96 B.n44 VSUBS 0.006622f
C97 B.n45 VSUBS 0.006622f
C98 B.n46 VSUBS 0.006622f
C99 B.n47 VSUBS 0.006622f
C100 B.n48 VSUBS 0.006622f
C101 B.n49 VSUBS 0.006622f
C102 B.n50 VSUBS 0.006622f
C103 B.n51 VSUBS 0.006622f
C104 B.n52 VSUBS 0.006622f
C105 B.n53 VSUBS 0.006622f
C106 B.n54 VSUBS 0.006622f
C107 B.n55 VSUBS 0.006622f
C108 B.n56 VSUBS 0.006622f
C109 B.n57 VSUBS 0.006622f
C110 B.n58 VSUBS 0.006622f
C111 B.n59 VSUBS 0.006622f
C112 B.n60 VSUBS 0.015228f
C113 B.n61 VSUBS 0.006622f
C114 B.n62 VSUBS 0.006622f
C115 B.n63 VSUBS 0.006622f
C116 B.n64 VSUBS 0.006622f
C117 B.n65 VSUBS 0.006622f
C118 B.n66 VSUBS 0.006622f
C119 B.n67 VSUBS 0.006622f
C120 B.n68 VSUBS 0.006622f
C121 B.n69 VSUBS 0.006622f
C122 B.n70 VSUBS 0.006622f
C123 B.n71 VSUBS 0.006622f
C124 B.n72 VSUBS 0.006622f
C125 B.n73 VSUBS 0.006622f
C126 B.n74 VSUBS 0.006622f
C127 B.n75 VSUBS 0.006622f
C128 B.n76 VSUBS 0.006622f
C129 B.n77 VSUBS 0.006622f
C130 B.n78 VSUBS 0.006622f
C131 B.n79 VSUBS 0.006622f
C132 B.n80 VSUBS 0.006622f
C133 B.n81 VSUBS 0.006622f
C134 B.n82 VSUBS 0.006622f
C135 B.n83 VSUBS 0.015989f
C136 B.n84 VSUBS 0.006622f
C137 B.n85 VSUBS 0.006622f
C138 B.n86 VSUBS 0.006622f
C139 B.n87 VSUBS 0.006622f
C140 B.n88 VSUBS 0.006622f
C141 B.n89 VSUBS 0.006622f
C142 B.n90 VSUBS 0.006622f
C143 B.n91 VSUBS 0.006622f
C144 B.n92 VSUBS 0.006622f
C145 B.n93 VSUBS 0.006622f
C146 B.n94 VSUBS 0.006622f
C147 B.n95 VSUBS 0.006622f
C148 B.n96 VSUBS 0.006622f
C149 B.n97 VSUBS 0.006622f
C150 B.n98 VSUBS 0.006622f
C151 B.n99 VSUBS 0.006622f
C152 B.n100 VSUBS 0.006622f
C153 B.n101 VSUBS 0.006622f
C154 B.t10 VSUBS 0.332372f
C155 B.t11 VSUBS 0.349055f
C156 B.t9 VSUBS 0.937812f
C157 B.n102 VSUBS 0.171122f
C158 B.n103 VSUBS 0.06558f
C159 B.n104 VSUBS 0.015342f
C160 B.n105 VSUBS 0.006622f
C161 B.n106 VSUBS 0.006622f
C162 B.n107 VSUBS 0.006622f
C163 B.n108 VSUBS 0.006622f
C164 B.n109 VSUBS 0.006622f
C165 B.t7 VSUBS 0.332377f
C166 B.t8 VSUBS 0.349061f
C167 B.t6 VSUBS 0.937812f
C168 B.n110 VSUBS 0.171117f
C169 B.n111 VSUBS 0.065574f
C170 B.n112 VSUBS 0.006622f
C171 B.n113 VSUBS 0.006622f
C172 B.n114 VSUBS 0.006622f
C173 B.n115 VSUBS 0.006622f
C174 B.n116 VSUBS 0.006622f
C175 B.n117 VSUBS 0.006622f
C176 B.n118 VSUBS 0.006622f
C177 B.n119 VSUBS 0.006622f
C178 B.n120 VSUBS 0.006622f
C179 B.n121 VSUBS 0.006622f
C180 B.n122 VSUBS 0.006622f
C181 B.n123 VSUBS 0.006622f
C182 B.n124 VSUBS 0.006622f
C183 B.n125 VSUBS 0.006622f
C184 B.n126 VSUBS 0.006622f
C185 B.n127 VSUBS 0.006622f
C186 B.n128 VSUBS 0.006622f
C187 B.n129 VSUBS 0.006622f
C188 B.n130 VSUBS 0.015989f
C189 B.n131 VSUBS 0.006622f
C190 B.n132 VSUBS 0.006622f
C191 B.n133 VSUBS 0.006622f
C192 B.n134 VSUBS 0.006622f
C193 B.n135 VSUBS 0.006622f
C194 B.n136 VSUBS 0.006622f
C195 B.n137 VSUBS 0.006622f
C196 B.n138 VSUBS 0.006622f
C197 B.n139 VSUBS 0.006622f
C198 B.n140 VSUBS 0.006622f
C199 B.n141 VSUBS 0.006622f
C200 B.n142 VSUBS 0.006622f
C201 B.n143 VSUBS 0.006622f
C202 B.n144 VSUBS 0.006622f
C203 B.n145 VSUBS 0.006622f
C204 B.n146 VSUBS 0.006622f
C205 B.n147 VSUBS 0.006622f
C206 B.n148 VSUBS 0.006622f
C207 B.n149 VSUBS 0.006622f
C208 B.n150 VSUBS 0.006622f
C209 B.n151 VSUBS 0.006622f
C210 B.n152 VSUBS 0.006622f
C211 B.n153 VSUBS 0.006622f
C212 B.n154 VSUBS 0.006622f
C213 B.n155 VSUBS 0.006622f
C214 B.n156 VSUBS 0.006622f
C215 B.n157 VSUBS 0.006622f
C216 B.n158 VSUBS 0.006622f
C217 B.n159 VSUBS 0.006622f
C218 B.n160 VSUBS 0.006622f
C219 B.n161 VSUBS 0.006622f
C220 B.n162 VSUBS 0.006622f
C221 B.n163 VSUBS 0.006622f
C222 B.n164 VSUBS 0.006622f
C223 B.n165 VSUBS 0.006622f
C224 B.n166 VSUBS 0.006622f
C225 B.n167 VSUBS 0.006622f
C226 B.n168 VSUBS 0.006622f
C227 B.n169 VSUBS 0.006622f
C228 B.n170 VSUBS 0.006622f
C229 B.n171 VSUBS 0.015562f
C230 B.n172 VSUBS 0.015562f
C231 B.n173 VSUBS 0.015989f
C232 B.n174 VSUBS 0.006622f
C233 B.n175 VSUBS 0.006622f
C234 B.n176 VSUBS 0.006622f
C235 B.n177 VSUBS 0.006622f
C236 B.n178 VSUBS 0.006622f
C237 B.n179 VSUBS 0.006622f
C238 B.n180 VSUBS 0.006622f
C239 B.n181 VSUBS 0.006622f
C240 B.n182 VSUBS 0.006622f
C241 B.n183 VSUBS 0.006622f
C242 B.n184 VSUBS 0.006622f
C243 B.n185 VSUBS 0.006622f
C244 B.n186 VSUBS 0.006622f
C245 B.n187 VSUBS 0.006622f
C246 B.n188 VSUBS 0.006622f
C247 B.n189 VSUBS 0.006622f
C248 B.n190 VSUBS 0.006622f
C249 B.n191 VSUBS 0.006622f
C250 B.n192 VSUBS 0.006622f
C251 B.n193 VSUBS 0.006622f
C252 B.n194 VSUBS 0.006622f
C253 B.n195 VSUBS 0.006622f
C254 B.n196 VSUBS 0.006622f
C255 B.n197 VSUBS 0.006622f
C256 B.n198 VSUBS 0.006622f
C257 B.n199 VSUBS 0.006622f
C258 B.n200 VSUBS 0.006622f
C259 B.n201 VSUBS 0.006622f
C260 B.n202 VSUBS 0.006622f
C261 B.n203 VSUBS 0.006622f
C262 B.n204 VSUBS 0.006622f
C263 B.n205 VSUBS 0.006622f
C264 B.n206 VSUBS 0.006622f
C265 B.n207 VSUBS 0.006622f
C266 B.n208 VSUBS 0.006622f
C267 B.n209 VSUBS 0.006622f
C268 B.n210 VSUBS 0.006622f
C269 B.n211 VSUBS 0.006622f
C270 B.n212 VSUBS 0.006622f
C271 B.n213 VSUBS 0.006622f
C272 B.n214 VSUBS 0.006622f
C273 B.n215 VSUBS 0.006622f
C274 B.n216 VSUBS 0.006622f
C275 B.n217 VSUBS 0.006622f
C276 B.n218 VSUBS 0.006622f
C277 B.n219 VSUBS 0.006622f
C278 B.n220 VSUBS 0.006622f
C279 B.n221 VSUBS 0.006622f
C280 B.n222 VSUBS 0.006622f
C281 B.n223 VSUBS 0.006622f
C282 B.n224 VSUBS 0.006622f
C283 B.n225 VSUBS 0.006622f
C284 B.n226 VSUBS 0.006622f
C285 B.n227 VSUBS 0.006622f
C286 B.n228 VSUBS 0.006622f
C287 B.n229 VSUBS 0.006232f
C288 B.n230 VSUBS 0.015342f
C289 B.n231 VSUBS 0.0037f
C290 B.n232 VSUBS 0.006622f
C291 B.n233 VSUBS 0.006622f
C292 B.n234 VSUBS 0.006622f
C293 B.n235 VSUBS 0.006622f
C294 B.n236 VSUBS 0.006622f
C295 B.n237 VSUBS 0.006622f
C296 B.n238 VSUBS 0.006622f
C297 B.n239 VSUBS 0.006622f
C298 B.n240 VSUBS 0.006622f
C299 B.n241 VSUBS 0.006622f
C300 B.n242 VSUBS 0.006622f
C301 B.n243 VSUBS 0.006622f
C302 B.n244 VSUBS 0.0037f
C303 B.n245 VSUBS 0.006622f
C304 B.n246 VSUBS 0.006622f
C305 B.n247 VSUBS 0.006232f
C306 B.n248 VSUBS 0.006622f
C307 B.n249 VSUBS 0.006622f
C308 B.n250 VSUBS 0.006622f
C309 B.n251 VSUBS 0.006622f
C310 B.n252 VSUBS 0.006622f
C311 B.n253 VSUBS 0.006622f
C312 B.n254 VSUBS 0.006622f
C313 B.n255 VSUBS 0.006622f
C314 B.n256 VSUBS 0.006622f
C315 B.n257 VSUBS 0.006622f
C316 B.n258 VSUBS 0.006622f
C317 B.n259 VSUBS 0.006622f
C318 B.n260 VSUBS 0.006622f
C319 B.n261 VSUBS 0.006622f
C320 B.n262 VSUBS 0.006622f
C321 B.n263 VSUBS 0.006622f
C322 B.n264 VSUBS 0.006622f
C323 B.n265 VSUBS 0.006622f
C324 B.n266 VSUBS 0.006622f
C325 B.n267 VSUBS 0.006622f
C326 B.n268 VSUBS 0.006622f
C327 B.n269 VSUBS 0.006622f
C328 B.n270 VSUBS 0.006622f
C329 B.n271 VSUBS 0.006622f
C330 B.n272 VSUBS 0.006622f
C331 B.n273 VSUBS 0.006622f
C332 B.n274 VSUBS 0.006622f
C333 B.n275 VSUBS 0.006622f
C334 B.n276 VSUBS 0.006622f
C335 B.n277 VSUBS 0.006622f
C336 B.n278 VSUBS 0.006622f
C337 B.n279 VSUBS 0.006622f
C338 B.n280 VSUBS 0.006622f
C339 B.n281 VSUBS 0.006622f
C340 B.n282 VSUBS 0.006622f
C341 B.n283 VSUBS 0.006622f
C342 B.n284 VSUBS 0.006622f
C343 B.n285 VSUBS 0.006622f
C344 B.n286 VSUBS 0.006622f
C345 B.n287 VSUBS 0.006622f
C346 B.n288 VSUBS 0.006622f
C347 B.n289 VSUBS 0.006622f
C348 B.n290 VSUBS 0.006622f
C349 B.n291 VSUBS 0.006622f
C350 B.n292 VSUBS 0.006622f
C351 B.n293 VSUBS 0.006622f
C352 B.n294 VSUBS 0.006622f
C353 B.n295 VSUBS 0.006622f
C354 B.n296 VSUBS 0.006622f
C355 B.n297 VSUBS 0.006622f
C356 B.n298 VSUBS 0.006622f
C357 B.n299 VSUBS 0.006622f
C358 B.n300 VSUBS 0.006622f
C359 B.n301 VSUBS 0.006622f
C360 B.n302 VSUBS 0.015989f
C361 B.n303 VSUBS 0.015562f
C362 B.n304 VSUBS 0.015562f
C363 B.n305 VSUBS 0.006622f
C364 B.n306 VSUBS 0.006622f
C365 B.n307 VSUBS 0.006622f
C366 B.n308 VSUBS 0.006622f
C367 B.n309 VSUBS 0.006622f
C368 B.n310 VSUBS 0.006622f
C369 B.n311 VSUBS 0.006622f
C370 B.n312 VSUBS 0.006622f
C371 B.n313 VSUBS 0.006622f
C372 B.n314 VSUBS 0.006622f
C373 B.n315 VSUBS 0.006622f
C374 B.n316 VSUBS 0.006622f
C375 B.n317 VSUBS 0.006622f
C376 B.n318 VSUBS 0.006622f
C377 B.n319 VSUBS 0.006622f
C378 B.n320 VSUBS 0.006622f
C379 B.n321 VSUBS 0.006622f
C380 B.n322 VSUBS 0.006622f
C381 B.n323 VSUBS 0.006622f
C382 B.n324 VSUBS 0.006622f
C383 B.n325 VSUBS 0.006622f
C384 B.n326 VSUBS 0.006622f
C385 B.n327 VSUBS 0.006622f
C386 B.n328 VSUBS 0.006622f
C387 B.n329 VSUBS 0.006622f
C388 B.n330 VSUBS 0.006622f
C389 B.n331 VSUBS 0.006622f
C390 B.n332 VSUBS 0.006622f
C391 B.n333 VSUBS 0.006622f
C392 B.n334 VSUBS 0.006622f
C393 B.n335 VSUBS 0.006622f
C394 B.n336 VSUBS 0.006622f
C395 B.n337 VSUBS 0.006622f
C396 B.n338 VSUBS 0.006622f
C397 B.n339 VSUBS 0.006622f
C398 B.n340 VSUBS 0.006622f
C399 B.n341 VSUBS 0.006622f
C400 B.n342 VSUBS 0.006622f
C401 B.n343 VSUBS 0.006622f
C402 B.n344 VSUBS 0.006622f
C403 B.n345 VSUBS 0.006622f
C404 B.n346 VSUBS 0.006622f
C405 B.n347 VSUBS 0.006622f
C406 B.n348 VSUBS 0.006622f
C407 B.n349 VSUBS 0.006622f
C408 B.n350 VSUBS 0.006622f
C409 B.n351 VSUBS 0.006622f
C410 B.n352 VSUBS 0.006622f
C411 B.n353 VSUBS 0.006622f
C412 B.n354 VSUBS 0.006622f
C413 B.n355 VSUBS 0.006622f
C414 B.n356 VSUBS 0.006622f
C415 B.n357 VSUBS 0.006622f
C416 B.n358 VSUBS 0.006622f
C417 B.n359 VSUBS 0.006622f
C418 B.n360 VSUBS 0.006622f
C419 B.n361 VSUBS 0.006622f
C420 B.n362 VSUBS 0.006622f
C421 B.n363 VSUBS 0.006622f
C422 B.n364 VSUBS 0.006622f
C423 B.n365 VSUBS 0.006622f
C424 B.n366 VSUBS 0.006622f
C425 B.n367 VSUBS 0.006622f
C426 B.n368 VSUBS 0.006622f
C427 B.n369 VSUBS 0.016323f
C428 B.n370 VSUBS 0.015562f
C429 B.n371 VSUBS 0.015989f
C430 B.n372 VSUBS 0.006622f
C431 B.n373 VSUBS 0.006622f
C432 B.n374 VSUBS 0.006622f
C433 B.n375 VSUBS 0.006622f
C434 B.n376 VSUBS 0.006622f
C435 B.n377 VSUBS 0.006622f
C436 B.n378 VSUBS 0.006622f
C437 B.n379 VSUBS 0.006622f
C438 B.n380 VSUBS 0.006622f
C439 B.n381 VSUBS 0.006622f
C440 B.n382 VSUBS 0.006622f
C441 B.n383 VSUBS 0.006622f
C442 B.n384 VSUBS 0.006622f
C443 B.n385 VSUBS 0.006622f
C444 B.n386 VSUBS 0.006622f
C445 B.n387 VSUBS 0.006622f
C446 B.n388 VSUBS 0.006622f
C447 B.n389 VSUBS 0.006622f
C448 B.n390 VSUBS 0.006622f
C449 B.n391 VSUBS 0.006622f
C450 B.n392 VSUBS 0.006622f
C451 B.n393 VSUBS 0.006622f
C452 B.n394 VSUBS 0.006622f
C453 B.n395 VSUBS 0.006622f
C454 B.n396 VSUBS 0.006622f
C455 B.n397 VSUBS 0.006622f
C456 B.n398 VSUBS 0.006622f
C457 B.n399 VSUBS 0.006622f
C458 B.n400 VSUBS 0.006622f
C459 B.n401 VSUBS 0.006622f
C460 B.n402 VSUBS 0.006622f
C461 B.n403 VSUBS 0.006622f
C462 B.n404 VSUBS 0.006622f
C463 B.n405 VSUBS 0.006622f
C464 B.n406 VSUBS 0.006622f
C465 B.n407 VSUBS 0.006622f
C466 B.n408 VSUBS 0.006622f
C467 B.n409 VSUBS 0.006622f
C468 B.n410 VSUBS 0.006622f
C469 B.n411 VSUBS 0.006622f
C470 B.n412 VSUBS 0.006622f
C471 B.n413 VSUBS 0.006622f
C472 B.n414 VSUBS 0.006622f
C473 B.n415 VSUBS 0.006622f
C474 B.n416 VSUBS 0.006622f
C475 B.n417 VSUBS 0.006622f
C476 B.n418 VSUBS 0.006622f
C477 B.n419 VSUBS 0.006622f
C478 B.n420 VSUBS 0.006622f
C479 B.n421 VSUBS 0.006622f
C480 B.n422 VSUBS 0.006622f
C481 B.n423 VSUBS 0.006622f
C482 B.n424 VSUBS 0.006622f
C483 B.n425 VSUBS 0.006622f
C484 B.n426 VSUBS 0.006622f
C485 B.n427 VSUBS 0.006232f
C486 B.n428 VSUBS 0.015342f
C487 B.n429 VSUBS 0.0037f
C488 B.n430 VSUBS 0.006622f
C489 B.n431 VSUBS 0.006622f
C490 B.n432 VSUBS 0.006622f
C491 B.n433 VSUBS 0.006622f
C492 B.n434 VSUBS 0.006622f
C493 B.n435 VSUBS 0.006622f
C494 B.n436 VSUBS 0.006622f
C495 B.n437 VSUBS 0.006622f
C496 B.n438 VSUBS 0.006622f
C497 B.n439 VSUBS 0.006622f
C498 B.n440 VSUBS 0.006622f
C499 B.n441 VSUBS 0.006622f
C500 B.n442 VSUBS 0.0037f
C501 B.n443 VSUBS 0.006622f
C502 B.n444 VSUBS 0.006622f
C503 B.n445 VSUBS 0.006232f
C504 B.n446 VSUBS 0.006622f
C505 B.n447 VSUBS 0.006622f
C506 B.n448 VSUBS 0.006622f
C507 B.n449 VSUBS 0.006622f
C508 B.n450 VSUBS 0.006622f
C509 B.n451 VSUBS 0.006622f
C510 B.n452 VSUBS 0.006622f
C511 B.n453 VSUBS 0.006622f
C512 B.n454 VSUBS 0.006622f
C513 B.n455 VSUBS 0.006622f
C514 B.n456 VSUBS 0.006622f
C515 B.n457 VSUBS 0.006622f
C516 B.n458 VSUBS 0.006622f
C517 B.n459 VSUBS 0.006622f
C518 B.n460 VSUBS 0.006622f
C519 B.n461 VSUBS 0.006622f
C520 B.n462 VSUBS 0.006622f
C521 B.n463 VSUBS 0.006622f
C522 B.n464 VSUBS 0.006622f
C523 B.n465 VSUBS 0.006622f
C524 B.n466 VSUBS 0.006622f
C525 B.n467 VSUBS 0.006622f
C526 B.n468 VSUBS 0.006622f
C527 B.n469 VSUBS 0.006622f
C528 B.n470 VSUBS 0.006622f
C529 B.n471 VSUBS 0.006622f
C530 B.n472 VSUBS 0.006622f
C531 B.n473 VSUBS 0.006622f
C532 B.n474 VSUBS 0.006622f
C533 B.n475 VSUBS 0.006622f
C534 B.n476 VSUBS 0.006622f
C535 B.n477 VSUBS 0.006622f
C536 B.n478 VSUBS 0.006622f
C537 B.n479 VSUBS 0.006622f
C538 B.n480 VSUBS 0.006622f
C539 B.n481 VSUBS 0.006622f
C540 B.n482 VSUBS 0.006622f
C541 B.n483 VSUBS 0.006622f
C542 B.n484 VSUBS 0.006622f
C543 B.n485 VSUBS 0.006622f
C544 B.n486 VSUBS 0.006622f
C545 B.n487 VSUBS 0.006622f
C546 B.n488 VSUBS 0.006622f
C547 B.n489 VSUBS 0.006622f
C548 B.n490 VSUBS 0.006622f
C549 B.n491 VSUBS 0.006622f
C550 B.n492 VSUBS 0.006622f
C551 B.n493 VSUBS 0.006622f
C552 B.n494 VSUBS 0.006622f
C553 B.n495 VSUBS 0.006622f
C554 B.n496 VSUBS 0.006622f
C555 B.n497 VSUBS 0.006622f
C556 B.n498 VSUBS 0.006622f
C557 B.n499 VSUBS 0.006622f
C558 B.n500 VSUBS 0.015989f
C559 B.n501 VSUBS 0.015562f
C560 B.n502 VSUBS 0.015562f
C561 B.n503 VSUBS 0.006622f
C562 B.n504 VSUBS 0.006622f
C563 B.n505 VSUBS 0.006622f
C564 B.n506 VSUBS 0.006622f
C565 B.n507 VSUBS 0.006622f
C566 B.n508 VSUBS 0.006622f
C567 B.n509 VSUBS 0.006622f
C568 B.n510 VSUBS 0.006622f
C569 B.n511 VSUBS 0.006622f
C570 B.n512 VSUBS 0.006622f
C571 B.n513 VSUBS 0.006622f
C572 B.n514 VSUBS 0.006622f
C573 B.n515 VSUBS 0.006622f
C574 B.n516 VSUBS 0.006622f
C575 B.n517 VSUBS 0.006622f
C576 B.n518 VSUBS 0.006622f
C577 B.n519 VSUBS 0.006622f
C578 B.n520 VSUBS 0.006622f
C579 B.n521 VSUBS 0.006622f
C580 B.n522 VSUBS 0.006622f
C581 B.n523 VSUBS 0.006622f
C582 B.n524 VSUBS 0.006622f
C583 B.n525 VSUBS 0.006622f
C584 B.n526 VSUBS 0.006622f
C585 B.n527 VSUBS 0.006622f
C586 B.n528 VSUBS 0.006622f
C587 B.n529 VSUBS 0.006622f
C588 B.n530 VSUBS 0.006622f
C589 B.n531 VSUBS 0.006622f
C590 B.n532 VSUBS 0.006622f
C591 B.n533 VSUBS 0.006622f
C592 B.n534 VSUBS 0.006622f
C593 B.n535 VSUBS 0.014994f
.ends

