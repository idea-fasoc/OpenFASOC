* NGSPICE file created from diff_pair_sample_1563.ext - technology: sky130A

.subckt diff_pair_sample_1563 VTAIL VN VP B VDD2 VDD1
X0 B.t15 B.t13 B.t14 B.t3 sky130_fd_pr__nfet_01v8 ad=6.4623 pd=33.92 as=0 ps=0 w=16.57 l=1.71
X1 VDD1.t1 VP.t0 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=6.4623 pd=33.92 as=6.4623 ps=33.92 w=16.57 l=1.71
X2 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=6.4623 pd=33.92 as=0 ps=0 w=16.57 l=1.71
X3 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=6.4623 pd=33.92 as=0 ps=0 w=16.57 l=1.71
X4 VDD2.t1 VN.t0 VTAIL.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=6.4623 pd=33.92 as=6.4623 ps=33.92 w=16.57 l=1.71
X5 VDD2.t0 VN.t1 VTAIL.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=6.4623 pd=33.92 as=6.4623 ps=33.92 w=16.57 l=1.71
X6 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=6.4623 pd=33.92 as=0 ps=0 w=16.57 l=1.71
X7 VDD1.t0 VP.t1 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=6.4623 pd=33.92 as=6.4623 ps=33.92 w=16.57 l=1.71
R0 B.n772 B.n771 585
R1 B.n341 B.n100 585
R2 B.n340 B.n339 585
R3 B.n338 B.n337 585
R4 B.n336 B.n335 585
R5 B.n334 B.n333 585
R6 B.n332 B.n331 585
R7 B.n330 B.n329 585
R8 B.n328 B.n327 585
R9 B.n326 B.n325 585
R10 B.n324 B.n323 585
R11 B.n322 B.n321 585
R12 B.n320 B.n319 585
R13 B.n318 B.n317 585
R14 B.n316 B.n315 585
R15 B.n314 B.n313 585
R16 B.n312 B.n311 585
R17 B.n310 B.n309 585
R18 B.n308 B.n307 585
R19 B.n306 B.n305 585
R20 B.n304 B.n303 585
R21 B.n302 B.n301 585
R22 B.n300 B.n299 585
R23 B.n298 B.n297 585
R24 B.n296 B.n295 585
R25 B.n294 B.n293 585
R26 B.n292 B.n291 585
R27 B.n290 B.n289 585
R28 B.n288 B.n287 585
R29 B.n286 B.n285 585
R30 B.n284 B.n283 585
R31 B.n282 B.n281 585
R32 B.n280 B.n279 585
R33 B.n278 B.n277 585
R34 B.n276 B.n275 585
R35 B.n274 B.n273 585
R36 B.n272 B.n271 585
R37 B.n270 B.n269 585
R38 B.n268 B.n267 585
R39 B.n266 B.n265 585
R40 B.n264 B.n263 585
R41 B.n262 B.n261 585
R42 B.n260 B.n259 585
R43 B.n258 B.n257 585
R44 B.n256 B.n255 585
R45 B.n254 B.n253 585
R46 B.n252 B.n251 585
R47 B.n250 B.n249 585
R48 B.n248 B.n247 585
R49 B.n246 B.n245 585
R50 B.n244 B.n243 585
R51 B.n242 B.n241 585
R52 B.n240 B.n239 585
R53 B.n238 B.n237 585
R54 B.n236 B.n235 585
R55 B.n233 B.n232 585
R56 B.n231 B.n230 585
R57 B.n229 B.n228 585
R58 B.n227 B.n226 585
R59 B.n225 B.n224 585
R60 B.n223 B.n222 585
R61 B.n221 B.n220 585
R62 B.n219 B.n218 585
R63 B.n217 B.n216 585
R64 B.n215 B.n214 585
R65 B.n212 B.n211 585
R66 B.n210 B.n209 585
R67 B.n208 B.n207 585
R68 B.n206 B.n205 585
R69 B.n204 B.n203 585
R70 B.n202 B.n201 585
R71 B.n200 B.n199 585
R72 B.n198 B.n197 585
R73 B.n196 B.n195 585
R74 B.n194 B.n193 585
R75 B.n192 B.n191 585
R76 B.n190 B.n189 585
R77 B.n188 B.n187 585
R78 B.n186 B.n185 585
R79 B.n184 B.n183 585
R80 B.n182 B.n181 585
R81 B.n180 B.n179 585
R82 B.n178 B.n177 585
R83 B.n176 B.n175 585
R84 B.n174 B.n173 585
R85 B.n172 B.n171 585
R86 B.n170 B.n169 585
R87 B.n168 B.n167 585
R88 B.n166 B.n165 585
R89 B.n164 B.n163 585
R90 B.n162 B.n161 585
R91 B.n160 B.n159 585
R92 B.n158 B.n157 585
R93 B.n156 B.n155 585
R94 B.n154 B.n153 585
R95 B.n152 B.n151 585
R96 B.n150 B.n149 585
R97 B.n148 B.n147 585
R98 B.n146 B.n145 585
R99 B.n144 B.n143 585
R100 B.n142 B.n141 585
R101 B.n140 B.n139 585
R102 B.n138 B.n137 585
R103 B.n136 B.n135 585
R104 B.n134 B.n133 585
R105 B.n132 B.n131 585
R106 B.n130 B.n129 585
R107 B.n128 B.n127 585
R108 B.n126 B.n125 585
R109 B.n124 B.n123 585
R110 B.n122 B.n121 585
R111 B.n120 B.n119 585
R112 B.n118 B.n117 585
R113 B.n116 B.n115 585
R114 B.n114 B.n113 585
R115 B.n112 B.n111 585
R116 B.n110 B.n109 585
R117 B.n108 B.n107 585
R118 B.n106 B.n105 585
R119 B.n39 B.n38 585
R120 B.n770 B.n40 585
R121 B.n775 B.n40 585
R122 B.n769 B.n768 585
R123 B.n768 B.n36 585
R124 B.n767 B.n35 585
R125 B.n781 B.n35 585
R126 B.n766 B.n34 585
R127 B.n782 B.n34 585
R128 B.n765 B.n33 585
R129 B.n783 B.n33 585
R130 B.n764 B.n763 585
R131 B.n763 B.n29 585
R132 B.n762 B.n28 585
R133 B.n789 B.n28 585
R134 B.n761 B.n27 585
R135 B.n790 B.n27 585
R136 B.n760 B.n26 585
R137 B.n791 B.n26 585
R138 B.n759 B.n758 585
R139 B.n758 B.n22 585
R140 B.n757 B.n21 585
R141 B.n797 B.n21 585
R142 B.n756 B.n20 585
R143 B.n798 B.n20 585
R144 B.n755 B.n19 585
R145 B.n799 B.n19 585
R146 B.n754 B.n753 585
R147 B.n753 B.n15 585
R148 B.n752 B.n14 585
R149 B.n805 B.n14 585
R150 B.n751 B.n13 585
R151 B.n806 B.n13 585
R152 B.n750 B.n12 585
R153 B.n807 B.n12 585
R154 B.n749 B.n748 585
R155 B.n748 B.n8 585
R156 B.n747 B.n7 585
R157 B.n813 B.n7 585
R158 B.n746 B.n6 585
R159 B.n814 B.n6 585
R160 B.n745 B.n5 585
R161 B.n815 B.n5 585
R162 B.n744 B.n743 585
R163 B.n743 B.n4 585
R164 B.n742 B.n342 585
R165 B.n742 B.n741 585
R166 B.n732 B.n343 585
R167 B.n344 B.n343 585
R168 B.n734 B.n733 585
R169 B.n735 B.n734 585
R170 B.n731 B.n348 585
R171 B.n352 B.n348 585
R172 B.n730 B.n729 585
R173 B.n729 B.n728 585
R174 B.n350 B.n349 585
R175 B.n351 B.n350 585
R176 B.n721 B.n720 585
R177 B.n722 B.n721 585
R178 B.n719 B.n357 585
R179 B.n357 B.n356 585
R180 B.n718 B.n717 585
R181 B.n717 B.n716 585
R182 B.n359 B.n358 585
R183 B.n360 B.n359 585
R184 B.n709 B.n708 585
R185 B.n710 B.n709 585
R186 B.n707 B.n365 585
R187 B.n365 B.n364 585
R188 B.n706 B.n705 585
R189 B.n705 B.n704 585
R190 B.n367 B.n366 585
R191 B.n368 B.n367 585
R192 B.n697 B.n696 585
R193 B.n698 B.n697 585
R194 B.n695 B.n373 585
R195 B.n373 B.n372 585
R196 B.n694 B.n693 585
R197 B.n693 B.n692 585
R198 B.n375 B.n374 585
R199 B.n376 B.n375 585
R200 B.n685 B.n684 585
R201 B.n686 B.n685 585
R202 B.n379 B.n378 585
R203 B.n448 B.n447 585
R204 B.n449 B.n445 585
R205 B.n445 B.n380 585
R206 B.n451 B.n450 585
R207 B.n453 B.n444 585
R208 B.n456 B.n455 585
R209 B.n457 B.n443 585
R210 B.n459 B.n458 585
R211 B.n461 B.n442 585
R212 B.n464 B.n463 585
R213 B.n465 B.n441 585
R214 B.n467 B.n466 585
R215 B.n469 B.n440 585
R216 B.n472 B.n471 585
R217 B.n473 B.n439 585
R218 B.n475 B.n474 585
R219 B.n477 B.n438 585
R220 B.n480 B.n479 585
R221 B.n481 B.n437 585
R222 B.n483 B.n482 585
R223 B.n485 B.n436 585
R224 B.n488 B.n487 585
R225 B.n489 B.n435 585
R226 B.n491 B.n490 585
R227 B.n493 B.n434 585
R228 B.n496 B.n495 585
R229 B.n497 B.n433 585
R230 B.n499 B.n498 585
R231 B.n501 B.n432 585
R232 B.n504 B.n503 585
R233 B.n505 B.n431 585
R234 B.n507 B.n506 585
R235 B.n509 B.n430 585
R236 B.n512 B.n511 585
R237 B.n513 B.n429 585
R238 B.n515 B.n514 585
R239 B.n517 B.n428 585
R240 B.n520 B.n519 585
R241 B.n521 B.n427 585
R242 B.n523 B.n522 585
R243 B.n525 B.n426 585
R244 B.n528 B.n527 585
R245 B.n529 B.n425 585
R246 B.n531 B.n530 585
R247 B.n533 B.n424 585
R248 B.n536 B.n535 585
R249 B.n537 B.n423 585
R250 B.n539 B.n538 585
R251 B.n541 B.n422 585
R252 B.n544 B.n543 585
R253 B.n545 B.n421 585
R254 B.n547 B.n546 585
R255 B.n549 B.n420 585
R256 B.n552 B.n551 585
R257 B.n553 B.n417 585
R258 B.n556 B.n555 585
R259 B.n558 B.n416 585
R260 B.n561 B.n560 585
R261 B.n562 B.n415 585
R262 B.n564 B.n563 585
R263 B.n566 B.n414 585
R264 B.n569 B.n568 585
R265 B.n570 B.n413 585
R266 B.n572 B.n571 585
R267 B.n574 B.n412 585
R268 B.n577 B.n576 585
R269 B.n578 B.n408 585
R270 B.n580 B.n579 585
R271 B.n582 B.n407 585
R272 B.n585 B.n584 585
R273 B.n586 B.n406 585
R274 B.n588 B.n587 585
R275 B.n590 B.n405 585
R276 B.n593 B.n592 585
R277 B.n594 B.n404 585
R278 B.n596 B.n595 585
R279 B.n598 B.n403 585
R280 B.n601 B.n600 585
R281 B.n602 B.n402 585
R282 B.n604 B.n603 585
R283 B.n606 B.n401 585
R284 B.n609 B.n608 585
R285 B.n610 B.n400 585
R286 B.n612 B.n611 585
R287 B.n614 B.n399 585
R288 B.n617 B.n616 585
R289 B.n618 B.n398 585
R290 B.n620 B.n619 585
R291 B.n622 B.n397 585
R292 B.n625 B.n624 585
R293 B.n626 B.n396 585
R294 B.n628 B.n627 585
R295 B.n630 B.n395 585
R296 B.n633 B.n632 585
R297 B.n634 B.n394 585
R298 B.n636 B.n635 585
R299 B.n638 B.n393 585
R300 B.n641 B.n640 585
R301 B.n642 B.n392 585
R302 B.n644 B.n643 585
R303 B.n646 B.n391 585
R304 B.n649 B.n648 585
R305 B.n650 B.n390 585
R306 B.n652 B.n651 585
R307 B.n654 B.n389 585
R308 B.n657 B.n656 585
R309 B.n658 B.n388 585
R310 B.n660 B.n659 585
R311 B.n662 B.n387 585
R312 B.n665 B.n664 585
R313 B.n666 B.n386 585
R314 B.n668 B.n667 585
R315 B.n670 B.n385 585
R316 B.n673 B.n672 585
R317 B.n674 B.n384 585
R318 B.n676 B.n675 585
R319 B.n678 B.n383 585
R320 B.n679 B.n382 585
R321 B.n682 B.n681 585
R322 B.n683 B.n381 585
R323 B.n381 B.n380 585
R324 B.n688 B.n687 585
R325 B.n687 B.n686 585
R326 B.n689 B.n377 585
R327 B.n377 B.n376 585
R328 B.n691 B.n690 585
R329 B.n692 B.n691 585
R330 B.n371 B.n370 585
R331 B.n372 B.n371 585
R332 B.n700 B.n699 585
R333 B.n699 B.n698 585
R334 B.n701 B.n369 585
R335 B.n369 B.n368 585
R336 B.n703 B.n702 585
R337 B.n704 B.n703 585
R338 B.n363 B.n362 585
R339 B.n364 B.n363 585
R340 B.n712 B.n711 585
R341 B.n711 B.n710 585
R342 B.n713 B.n361 585
R343 B.n361 B.n360 585
R344 B.n715 B.n714 585
R345 B.n716 B.n715 585
R346 B.n355 B.n354 585
R347 B.n356 B.n355 585
R348 B.n724 B.n723 585
R349 B.n723 B.n722 585
R350 B.n725 B.n353 585
R351 B.n353 B.n351 585
R352 B.n727 B.n726 585
R353 B.n728 B.n727 585
R354 B.n347 B.n346 585
R355 B.n352 B.n347 585
R356 B.n737 B.n736 585
R357 B.n736 B.n735 585
R358 B.n738 B.n345 585
R359 B.n345 B.n344 585
R360 B.n740 B.n739 585
R361 B.n741 B.n740 585
R362 B.n2 B.n0 585
R363 B.n4 B.n2 585
R364 B.n3 B.n1 585
R365 B.n814 B.n3 585
R366 B.n812 B.n811 585
R367 B.n813 B.n812 585
R368 B.n810 B.n9 585
R369 B.n9 B.n8 585
R370 B.n809 B.n808 585
R371 B.n808 B.n807 585
R372 B.n11 B.n10 585
R373 B.n806 B.n11 585
R374 B.n804 B.n803 585
R375 B.n805 B.n804 585
R376 B.n802 B.n16 585
R377 B.n16 B.n15 585
R378 B.n801 B.n800 585
R379 B.n800 B.n799 585
R380 B.n18 B.n17 585
R381 B.n798 B.n18 585
R382 B.n796 B.n795 585
R383 B.n797 B.n796 585
R384 B.n794 B.n23 585
R385 B.n23 B.n22 585
R386 B.n793 B.n792 585
R387 B.n792 B.n791 585
R388 B.n25 B.n24 585
R389 B.n790 B.n25 585
R390 B.n788 B.n787 585
R391 B.n789 B.n788 585
R392 B.n786 B.n30 585
R393 B.n30 B.n29 585
R394 B.n785 B.n784 585
R395 B.n784 B.n783 585
R396 B.n32 B.n31 585
R397 B.n782 B.n32 585
R398 B.n780 B.n779 585
R399 B.n781 B.n780 585
R400 B.n778 B.n37 585
R401 B.n37 B.n36 585
R402 B.n777 B.n776 585
R403 B.n776 B.n775 585
R404 B.n817 B.n816 585
R405 B.n816 B.n815 585
R406 B.n687 B.n379 492.5
R407 B.n776 B.n39 492.5
R408 B.n685 B.n381 492.5
R409 B.n772 B.n40 492.5
R410 B.n409 B.t6 439.675
R411 B.n418 B.t10 439.675
R412 B.n103 B.t2 439.675
R413 B.n101 B.t13 439.675
R414 B.n774 B.n773 256.663
R415 B.n774 B.n99 256.663
R416 B.n774 B.n98 256.663
R417 B.n774 B.n97 256.663
R418 B.n774 B.n96 256.663
R419 B.n774 B.n95 256.663
R420 B.n774 B.n94 256.663
R421 B.n774 B.n93 256.663
R422 B.n774 B.n92 256.663
R423 B.n774 B.n91 256.663
R424 B.n774 B.n90 256.663
R425 B.n774 B.n89 256.663
R426 B.n774 B.n88 256.663
R427 B.n774 B.n87 256.663
R428 B.n774 B.n86 256.663
R429 B.n774 B.n85 256.663
R430 B.n774 B.n84 256.663
R431 B.n774 B.n83 256.663
R432 B.n774 B.n82 256.663
R433 B.n774 B.n81 256.663
R434 B.n774 B.n80 256.663
R435 B.n774 B.n79 256.663
R436 B.n774 B.n78 256.663
R437 B.n774 B.n77 256.663
R438 B.n774 B.n76 256.663
R439 B.n774 B.n75 256.663
R440 B.n774 B.n74 256.663
R441 B.n774 B.n73 256.663
R442 B.n774 B.n72 256.663
R443 B.n774 B.n71 256.663
R444 B.n774 B.n70 256.663
R445 B.n774 B.n69 256.663
R446 B.n774 B.n68 256.663
R447 B.n774 B.n67 256.663
R448 B.n774 B.n66 256.663
R449 B.n774 B.n65 256.663
R450 B.n774 B.n64 256.663
R451 B.n774 B.n63 256.663
R452 B.n774 B.n62 256.663
R453 B.n774 B.n61 256.663
R454 B.n774 B.n60 256.663
R455 B.n774 B.n59 256.663
R456 B.n774 B.n58 256.663
R457 B.n774 B.n57 256.663
R458 B.n774 B.n56 256.663
R459 B.n774 B.n55 256.663
R460 B.n774 B.n54 256.663
R461 B.n774 B.n53 256.663
R462 B.n774 B.n52 256.663
R463 B.n774 B.n51 256.663
R464 B.n774 B.n50 256.663
R465 B.n774 B.n49 256.663
R466 B.n774 B.n48 256.663
R467 B.n774 B.n47 256.663
R468 B.n774 B.n46 256.663
R469 B.n774 B.n45 256.663
R470 B.n774 B.n44 256.663
R471 B.n774 B.n43 256.663
R472 B.n774 B.n42 256.663
R473 B.n774 B.n41 256.663
R474 B.n446 B.n380 256.663
R475 B.n452 B.n380 256.663
R476 B.n454 B.n380 256.663
R477 B.n460 B.n380 256.663
R478 B.n462 B.n380 256.663
R479 B.n468 B.n380 256.663
R480 B.n470 B.n380 256.663
R481 B.n476 B.n380 256.663
R482 B.n478 B.n380 256.663
R483 B.n484 B.n380 256.663
R484 B.n486 B.n380 256.663
R485 B.n492 B.n380 256.663
R486 B.n494 B.n380 256.663
R487 B.n500 B.n380 256.663
R488 B.n502 B.n380 256.663
R489 B.n508 B.n380 256.663
R490 B.n510 B.n380 256.663
R491 B.n516 B.n380 256.663
R492 B.n518 B.n380 256.663
R493 B.n524 B.n380 256.663
R494 B.n526 B.n380 256.663
R495 B.n532 B.n380 256.663
R496 B.n534 B.n380 256.663
R497 B.n540 B.n380 256.663
R498 B.n542 B.n380 256.663
R499 B.n548 B.n380 256.663
R500 B.n550 B.n380 256.663
R501 B.n557 B.n380 256.663
R502 B.n559 B.n380 256.663
R503 B.n565 B.n380 256.663
R504 B.n567 B.n380 256.663
R505 B.n573 B.n380 256.663
R506 B.n575 B.n380 256.663
R507 B.n581 B.n380 256.663
R508 B.n583 B.n380 256.663
R509 B.n589 B.n380 256.663
R510 B.n591 B.n380 256.663
R511 B.n597 B.n380 256.663
R512 B.n599 B.n380 256.663
R513 B.n605 B.n380 256.663
R514 B.n607 B.n380 256.663
R515 B.n613 B.n380 256.663
R516 B.n615 B.n380 256.663
R517 B.n621 B.n380 256.663
R518 B.n623 B.n380 256.663
R519 B.n629 B.n380 256.663
R520 B.n631 B.n380 256.663
R521 B.n637 B.n380 256.663
R522 B.n639 B.n380 256.663
R523 B.n645 B.n380 256.663
R524 B.n647 B.n380 256.663
R525 B.n653 B.n380 256.663
R526 B.n655 B.n380 256.663
R527 B.n661 B.n380 256.663
R528 B.n663 B.n380 256.663
R529 B.n669 B.n380 256.663
R530 B.n671 B.n380 256.663
R531 B.n677 B.n380 256.663
R532 B.n680 B.n380 256.663
R533 B.n687 B.n377 163.367
R534 B.n691 B.n377 163.367
R535 B.n691 B.n371 163.367
R536 B.n699 B.n371 163.367
R537 B.n699 B.n369 163.367
R538 B.n703 B.n369 163.367
R539 B.n703 B.n363 163.367
R540 B.n711 B.n363 163.367
R541 B.n711 B.n361 163.367
R542 B.n715 B.n361 163.367
R543 B.n715 B.n355 163.367
R544 B.n723 B.n355 163.367
R545 B.n723 B.n353 163.367
R546 B.n727 B.n353 163.367
R547 B.n727 B.n347 163.367
R548 B.n736 B.n347 163.367
R549 B.n736 B.n345 163.367
R550 B.n740 B.n345 163.367
R551 B.n740 B.n2 163.367
R552 B.n816 B.n2 163.367
R553 B.n816 B.n3 163.367
R554 B.n812 B.n3 163.367
R555 B.n812 B.n9 163.367
R556 B.n808 B.n9 163.367
R557 B.n808 B.n11 163.367
R558 B.n804 B.n11 163.367
R559 B.n804 B.n16 163.367
R560 B.n800 B.n16 163.367
R561 B.n800 B.n18 163.367
R562 B.n796 B.n18 163.367
R563 B.n796 B.n23 163.367
R564 B.n792 B.n23 163.367
R565 B.n792 B.n25 163.367
R566 B.n788 B.n25 163.367
R567 B.n788 B.n30 163.367
R568 B.n784 B.n30 163.367
R569 B.n784 B.n32 163.367
R570 B.n780 B.n32 163.367
R571 B.n780 B.n37 163.367
R572 B.n776 B.n37 163.367
R573 B.n447 B.n445 163.367
R574 B.n451 B.n445 163.367
R575 B.n455 B.n453 163.367
R576 B.n459 B.n443 163.367
R577 B.n463 B.n461 163.367
R578 B.n467 B.n441 163.367
R579 B.n471 B.n469 163.367
R580 B.n475 B.n439 163.367
R581 B.n479 B.n477 163.367
R582 B.n483 B.n437 163.367
R583 B.n487 B.n485 163.367
R584 B.n491 B.n435 163.367
R585 B.n495 B.n493 163.367
R586 B.n499 B.n433 163.367
R587 B.n503 B.n501 163.367
R588 B.n507 B.n431 163.367
R589 B.n511 B.n509 163.367
R590 B.n515 B.n429 163.367
R591 B.n519 B.n517 163.367
R592 B.n523 B.n427 163.367
R593 B.n527 B.n525 163.367
R594 B.n531 B.n425 163.367
R595 B.n535 B.n533 163.367
R596 B.n539 B.n423 163.367
R597 B.n543 B.n541 163.367
R598 B.n547 B.n421 163.367
R599 B.n551 B.n549 163.367
R600 B.n556 B.n417 163.367
R601 B.n560 B.n558 163.367
R602 B.n564 B.n415 163.367
R603 B.n568 B.n566 163.367
R604 B.n572 B.n413 163.367
R605 B.n576 B.n574 163.367
R606 B.n580 B.n408 163.367
R607 B.n584 B.n582 163.367
R608 B.n588 B.n406 163.367
R609 B.n592 B.n590 163.367
R610 B.n596 B.n404 163.367
R611 B.n600 B.n598 163.367
R612 B.n604 B.n402 163.367
R613 B.n608 B.n606 163.367
R614 B.n612 B.n400 163.367
R615 B.n616 B.n614 163.367
R616 B.n620 B.n398 163.367
R617 B.n624 B.n622 163.367
R618 B.n628 B.n396 163.367
R619 B.n632 B.n630 163.367
R620 B.n636 B.n394 163.367
R621 B.n640 B.n638 163.367
R622 B.n644 B.n392 163.367
R623 B.n648 B.n646 163.367
R624 B.n652 B.n390 163.367
R625 B.n656 B.n654 163.367
R626 B.n660 B.n388 163.367
R627 B.n664 B.n662 163.367
R628 B.n668 B.n386 163.367
R629 B.n672 B.n670 163.367
R630 B.n676 B.n384 163.367
R631 B.n679 B.n678 163.367
R632 B.n681 B.n381 163.367
R633 B.n685 B.n375 163.367
R634 B.n693 B.n375 163.367
R635 B.n693 B.n373 163.367
R636 B.n697 B.n373 163.367
R637 B.n697 B.n367 163.367
R638 B.n705 B.n367 163.367
R639 B.n705 B.n365 163.367
R640 B.n709 B.n365 163.367
R641 B.n709 B.n359 163.367
R642 B.n717 B.n359 163.367
R643 B.n717 B.n357 163.367
R644 B.n721 B.n357 163.367
R645 B.n721 B.n350 163.367
R646 B.n729 B.n350 163.367
R647 B.n729 B.n348 163.367
R648 B.n734 B.n348 163.367
R649 B.n734 B.n343 163.367
R650 B.n742 B.n343 163.367
R651 B.n743 B.n742 163.367
R652 B.n743 B.n5 163.367
R653 B.n6 B.n5 163.367
R654 B.n7 B.n6 163.367
R655 B.n748 B.n7 163.367
R656 B.n748 B.n12 163.367
R657 B.n13 B.n12 163.367
R658 B.n14 B.n13 163.367
R659 B.n753 B.n14 163.367
R660 B.n753 B.n19 163.367
R661 B.n20 B.n19 163.367
R662 B.n21 B.n20 163.367
R663 B.n758 B.n21 163.367
R664 B.n758 B.n26 163.367
R665 B.n27 B.n26 163.367
R666 B.n28 B.n27 163.367
R667 B.n763 B.n28 163.367
R668 B.n763 B.n33 163.367
R669 B.n34 B.n33 163.367
R670 B.n35 B.n34 163.367
R671 B.n768 B.n35 163.367
R672 B.n768 B.n40 163.367
R673 B.n107 B.n106 163.367
R674 B.n111 B.n110 163.367
R675 B.n115 B.n114 163.367
R676 B.n119 B.n118 163.367
R677 B.n123 B.n122 163.367
R678 B.n127 B.n126 163.367
R679 B.n131 B.n130 163.367
R680 B.n135 B.n134 163.367
R681 B.n139 B.n138 163.367
R682 B.n143 B.n142 163.367
R683 B.n147 B.n146 163.367
R684 B.n151 B.n150 163.367
R685 B.n155 B.n154 163.367
R686 B.n159 B.n158 163.367
R687 B.n163 B.n162 163.367
R688 B.n167 B.n166 163.367
R689 B.n171 B.n170 163.367
R690 B.n175 B.n174 163.367
R691 B.n179 B.n178 163.367
R692 B.n183 B.n182 163.367
R693 B.n187 B.n186 163.367
R694 B.n191 B.n190 163.367
R695 B.n195 B.n194 163.367
R696 B.n199 B.n198 163.367
R697 B.n203 B.n202 163.367
R698 B.n207 B.n206 163.367
R699 B.n211 B.n210 163.367
R700 B.n216 B.n215 163.367
R701 B.n220 B.n219 163.367
R702 B.n224 B.n223 163.367
R703 B.n228 B.n227 163.367
R704 B.n232 B.n231 163.367
R705 B.n237 B.n236 163.367
R706 B.n241 B.n240 163.367
R707 B.n245 B.n244 163.367
R708 B.n249 B.n248 163.367
R709 B.n253 B.n252 163.367
R710 B.n257 B.n256 163.367
R711 B.n261 B.n260 163.367
R712 B.n265 B.n264 163.367
R713 B.n269 B.n268 163.367
R714 B.n273 B.n272 163.367
R715 B.n277 B.n276 163.367
R716 B.n281 B.n280 163.367
R717 B.n285 B.n284 163.367
R718 B.n289 B.n288 163.367
R719 B.n293 B.n292 163.367
R720 B.n297 B.n296 163.367
R721 B.n301 B.n300 163.367
R722 B.n305 B.n304 163.367
R723 B.n309 B.n308 163.367
R724 B.n313 B.n312 163.367
R725 B.n317 B.n316 163.367
R726 B.n321 B.n320 163.367
R727 B.n325 B.n324 163.367
R728 B.n329 B.n328 163.367
R729 B.n333 B.n332 163.367
R730 B.n337 B.n336 163.367
R731 B.n339 B.n100 163.367
R732 B.n409 B.t9 111.754
R733 B.n101 B.t14 111.754
R734 B.n418 B.t12 111.731
R735 B.n103 B.t4 111.731
R736 B.n410 B.t8 72.1898
R737 B.n102 B.t15 72.1898
R738 B.n419 B.t11 72.1681
R739 B.n104 B.t5 72.1681
R740 B.n446 B.n379 71.676
R741 B.n452 B.n451 71.676
R742 B.n455 B.n454 71.676
R743 B.n460 B.n459 71.676
R744 B.n463 B.n462 71.676
R745 B.n468 B.n467 71.676
R746 B.n471 B.n470 71.676
R747 B.n476 B.n475 71.676
R748 B.n479 B.n478 71.676
R749 B.n484 B.n483 71.676
R750 B.n487 B.n486 71.676
R751 B.n492 B.n491 71.676
R752 B.n495 B.n494 71.676
R753 B.n500 B.n499 71.676
R754 B.n503 B.n502 71.676
R755 B.n508 B.n507 71.676
R756 B.n511 B.n510 71.676
R757 B.n516 B.n515 71.676
R758 B.n519 B.n518 71.676
R759 B.n524 B.n523 71.676
R760 B.n527 B.n526 71.676
R761 B.n532 B.n531 71.676
R762 B.n535 B.n534 71.676
R763 B.n540 B.n539 71.676
R764 B.n543 B.n542 71.676
R765 B.n548 B.n547 71.676
R766 B.n551 B.n550 71.676
R767 B.n557 B.n556 71.676
R768 B.n560 B.n559 71.676
R769 B.n565 B.n564 71.676
R770 B.n568 B.n567 71.676
R771 B.n573 B.n572 71.676
R772 B.n576 B.n575 71.676
R773 B.n581 B.n580 71.676
R774 B.n584 B.n583 71.676
R775 B.n589 B.n588 71.676
R776 B.n592 B.n591 71.676
R777 B.n597 B.n596 71.676
R778 B.n600 B.n599 71.676
R779 B.n605 B.n604 71.676
R780 B.n608 B.n607 71.676
R781 B.n613 B.n612 71.676
R782 B.n616 B.n615 71.676
R783 B.n621 B.n620 71.676
R784 B.n624 B.n623 71.676
R785 B.n629 B.n628 71.676
R786 B.n632 B.n631 71.676
R787 B.n637 B.n636 71.676
R788 B.n640 B.n639 71.676
R789 B.n645 B.n644 71.676
R790 B.n648 B.n647 71.676
R791 B.n653 B.n652 71.676
R792 B.n656 B.n655 71.676
R793 B.n661 B.n660 71.676
R794 B.n664 B.n663 71.676
R795 B.n669 B.n668 71.676
R796 B.n672 B.n671 71.676
R797 B.n677 B.n676 71.676
R798 B.n680 B.n679 71.676
R799 B.n41 B.n39 71.676
R800 B.n107 B.n42 71.676
R801 B.n111 B.n43 71.676
R802 B.n115 B.n44 71.676
R803 B.n119 B.n45 71.676
R804 B.n123 B.n46 71.676
R805 B.n127 B.n47 71.676
R806 B.n131 B.n48 71.676
R807 B.n135 B.n49 71.676
R808 B.n139 B.n50 71.676
R809 B.n143 B.n51 71.676
R810 B.n147 B.n52 71.676
R811 B.n151 B.n53 71.676
R812 B.n155 B.n54 71.676
R813 B.n159 B.n55 71.676
R814 B.n163 B.n56 71.676
R815 B.n167 B.n57 71.676
R816 B.n171 B.n58 71.676
R817 B.n175 B.n59 71.676
R818 B.n179 B.n60 71.676
R819 B.n183 B.n61 71.676
R820 B.n187 B.n62 71.676
R821 B.n191 B.n63 71.676
R822 B.n195 B.n64 71.676
R823 B.n199 B.n65 71.676
R824 B.n203 B.n66 71.676
R825 B.n207 B.n67 71.676
R826 B.n211 B.n68 71.676
R827 B.n216 B.n69 71.676
R828 B.n220 B.n70 71.676
R829 B.n224 B.n71 71.676
R830 B.n228 B.n72 71.676
R831 B.n232 B.n73 71.676
R832 B.n237 B.n74 71.676
R833 B.n241 B.n75 71.676
R834 B.n245 B.n76 71.676
R835 B.n249 B.n77 71.676
R836 B.n253 B.n78 71.676
R837 B.n257 B.n79 71.676
R838 B.n261 B.n80 71.676
R839 B.n265 B.n81 71.676
R840 B.n269 B.n82 71.676
R841 B.n273 B.n83 71.676
R842 B.n277 B.n84 71.676
R843 B.n281 B.n85 71.676
R844 B.n285 B.n86 71.676
R845 B.n289 B.n87 71.676
R846 B.n293 B.n88 71.676
R847 B.n297 B.n89 71.676
R848 B.n301 B.n90 71.676
R849 B.n305 B.n91 71.676
R850 B.n309 B.n92 71.676
R851 B.n313 B.n93 71.676
R852 B.n317 B.n94 71.676
R853 B.n321 B.n95 71.676
R854 B.n325 B.n96 71.676
R855 B.n329 B.n97 71.676
R856 B.n333 B.n98 71.676
R857 B.n337 B.n99 71.676
R858 B.n773 B.n100 71.676
R859 B.n773 B.n772 71.676
R860 B.n339 B.n99 71.676
R861 B.n336 B.n98 71.676
R862 B.n332 B.n97 71.676
R863 B.n328 B.n96 71.676
R864 B.n324 B.n95 71.676
R865 B.n320 B.n94 71.676
R866 B.n316 B.n93 71.676
R867 B.n312 B.n92 71.676
R868 B.n308 B.n91 71.676
R869 B.n304 B.n90 71.676
R870 B.n300 B.n89 71.676
R871 B.n296 B.n88 71.676
R872 B.n292 B.n87 71.676
R873 B.n288 B.n86 71.676
R874 B.n284 B.n85 71.676
R875 B.n280 B.n84 71.676
R876 B.n276 B.n83 71.676
R877 B.n272 B.n82 71.676
R878 B.n268 B.n81 71.676
R879 B.n264 B.n80 71.676
R880 B.n260 B.n79 71.676
R881 B.n256 B.n78 71.676
R882 B.n252 B.n77 71.676
R883 B.n248 B.n76 71.676
R884 B.n244 B.n75 71.676
R885 B.n240 B.n74 71.676
R886 B.n236 B.n73 71.676
R887 B.n231 B.n72 71.676
R888 B.n227 B.n71 71.676
R889 B.n223 B.n70 71.676
R890 B.n219 B.n69 71.676
R891 B.n215 B.n68 71.676
R892 B.n210 B.n67 71.676
R893 B.n206 B.n66 71.676
R894 B.n202 B.n65 71.676
R895 B.n198 B.n64 71.676
R896 B.n194 B.n63 71.676
R897 B.n190 B.n62 71.676
R898 B.n186 B.n61 71.676
R899 B.n182 B.n60 71.676
R900 B.n178 B.n59 71.676
R901 B.n174 B.n58 71.676
R902 B.n170 B.n57 71.676
R903 B.n166 B.n56 71.676
R904 B.n162 B.n55 71.676
R905 B.n158 B.n54 71.676
R906 B.n154 B.n53 71.676
R907 B.n150 B.n52 71.676
R908 B.n146 B.n51 71.676
R909 B.n142 B.n50 71.676
R910 B.n138 B.n49 71.676
R911 B.n134 B.n48 71.676
R912 B.n130 B.n47 71.676
R913 B.n126 B.n46 71.676
R914 B.n122 B.n45 71.676
R915 B.n118 B.n44 71.676
R916 B.n114 B.n43 71.676
R917 B.n110 B.n42 71.676
R918 B.n106 B.n41 71.676
R919 B.n447 B.n446 71.676
R920 B.n453 B.n452 71.676
R921 B.n454 B.n443 71.676
R922 B.n461 B.n460 71.676
R923 B.n462 B.n441 71.676
R924 B.n469 B.n468 71.676
R925 B.n470 B.n439 71.676
R926 B.n477 B.n476 71.676
R927 B.n478 B.n437 71.676
R928 B.n485 B.n484 71.676
R929 B.n486 B.n435 71.676
R930 B.n493 B.n492 71.676
R931 B.n494 B.n433 71.676
R932 B.n501 B.n500 71.676
R933 B.n502 B.n431 71.676
R934 B.n509 B.n508 71.676
R935 B.n510 B.n429 71.676
R936 B.n517 B.n516 71.676
R937 B.n518 B.n427 71.676
R938 B.n525 B.n524 71.676
R939 B.n526 B.n425 71.676
R940 B.n533 B.n532 71.676
R941 B.n534 B.n423 71.676
R942 B.n541 B.n540 71.676
R943 B.n542 B.n421 71.676
R944 B.n549 B.n548 71.676
R945 B.n550 B.n417 71.676
R946 B.n558 B.n557 71.676
R947 B.n559 B.n415 71.676
R948 B.n566 B.n565 71.676
R949 B.n567 B.n413 71.676
R950 B.n574 B.n573 71.676
R951 B.n575 B.n408 71.676
R952 B.n582 B.n581 71.676
R953 B.n583 B.n406 71.676
R954 B.n590 B.n589 71.676
R955 B.n591 B.n404 71.676
R956 B.n598 B.n597 71.676
R957 B.n599 B.n402 71.676
R958 B.n606 B.n605 71.676
R959 B.n607 B.n400 71.676
R960 B.n614 B.n613 71.676
R961 B.n615 B.n398 71.676
R962 B.n622 B.n621 71.676
R963 B.n623 B.n396 71.676
R964 B.n630 B.n629 71.676
R965 B.n631 B.n394 71.676
R966 B.n638 B.n637 71.676
R967 B.n639 B.n392 71.676
R968 B.n646 B.n645 71.676
R969 B.n647 B.n390 71.676
R970 B.n654 B.n653 71.676
R971 B.n655 B.n388 71.676
R972 B.n662 B.n661 71.676
R973 B.n663 B.n386 71.676
R974 B.n670 B.n669 71.676
R975 B.n671 B.n384 71.676
R976 B.n678 B.n677 71.676
R977 B.n681 B.n680 71.676
R978 B.n686 B.n380 65.9653
R979 B.n775 B.n774 65.9653
R980 B.n411 B.n410 59.5399
R981 B.n554 B.n419 59.5399
R982 B.n213 B.n104 59.5399
R983 B.n234 B.n102 59.5399
R984 B.n410 B.n409 39.5641
R985 B.n419 B.n418 39.5641
R986 B.n104 B.n103 39.5641
R987 B.n102 B.n101 39.5641
R988 B.n686 B.n376 34.2417
R989 B.n692 B.n376 34.2417
R990 B.n692 B.n372 34.2417
R991 B.n698 B.n372 34.2417
R992 B.n698 B.n368 34.2417
R993 B.n704 B.n368 34.2417
R994 B.n710 B.n364 34.2417
R995 B.n710 B.n360 34.2417
R996 B.n716 B.n360 34.2417
R997 B.n716 B.n356 34.2417
R998 B.n722 B.n356 34.2417
R999 B.n722 B.n351 34.2417
R1000 B.n728 B.n351 34.2417
R1001 B.n728 B.n352 34.2417
R1002 B.n735 B.n344 34.2417
R1003 B.n741 B.n344 34.2417
R1004 B.n741 B.n4 34.2417
R1005 B.n815 B.n4 34.2417
R1006 B.n815 B.n814 34.2417
R1007 B.n814 B.n813 34.2417
R1008 B.n813 B.n8 34.2417
R1009 B.n807 B.n8 34.2417
R1010 B.n806 B.n805 34.2417
R1011 B.n805 B.n15 34.2417
R1012 B.n799 B.n15 34.2417
R1013 B.n799 B.n798 34.2417
R1014 B.n798 B.n797 34.2417
R1015 B.n797 B.n22 34.2417
R1016 B.n791 B.n22 34.2417
R1017 B.n791 B.n790 34.2417
R1018 B.n789 B.n29 34.2417
R1019 B.n783 B.n29 34.2417
R1020 B.n783 B.n782 34.2417
R1021 B.n782 B.n781 34.2417
R1022 B.n781 B.n36 34.2417
R1023 B.n775 B.n36 34.2417
R1024 B.n777 B.n38 32.0005
R1025 B.n771 B.n770 32.0005
R1026 B.n684 B.n683 32.0005
R1027 B.n688 B.n378 32.0005
R1028 B.t7 B.n364 27.6956
R1029 B.n790 B.t3 27.6956
R1030 B.n735 B.t0 20.646
R1031 B.n807 B.t1 20.646
R1032 B B.n817 18.0485
R1033 B.n352 B.t0 13.5963
R1034 B.t1 B.n806 13.5963
R1035 B.n105 B.n38 10.6151
R1036 B.n108 B.n105 10.6151
R1037 B.n109 B.n108 10.6151
R1038 B.n112 B.n109 10.6151
R1039 B.n113 B.n112 10.6151
R1040 B.n116 B.n113 10.6151
R1041 B.n117 B.n116 10.6151
R1042 B.n120 B.n117 10.6151
R1043 B.n121 B.n120 10.6151
R1044 B.n124 B.n121 10.6151
R1045 B.n125 B.n124 10.6151
R1046 B.n128 B.n125 10.6151
R1047 B.n129 B.n128 10.6151
R1048 B.n132 B.n129 10.6151
R1049 B.n133 B.n132 10.6151
R1050 B.n136 B.n133 10.6151
R1051 B.n137 B.n136 10.6151
R1052 B.n140 B.n137 10.6151
R1053 B.n141 B.n140 10.6151
R1054 B.n144 B.n141 10.6151
R1055 B.n145 B.n144 10.6151
R1056 B.n148 B.n145 10.6151
R1057 B.n149 B.n148 10.6151
R1058 B.n152 B.n149 10.6151
R1059 B.n153 B.n152 10.6151
R1060 B.n156 B.n153 10.6151
R1061 B.n157 B.n156 10.6151
R1062 B.n160 B.n157 10.6151
R1063 B.n161 B.n160 10.6151
R1064 B.n164 B.n161 10.6151
R1065 B.n165 B.n164 10.6151
R1066 B.n168 B.n165 10.6151
R1067 B.n169 B.n168 10.6151
R1068 B.n172 B.n169 10.6151
R1069 B.n173 B.n172 10.6151
R1070 B.n176 B.n173 10.6151
R1071 B.n177 B.n176 10.6151
R1072 B.n180 B.n177 10.6151
R1073 B.n181 B.n180 10.6151
R1074 B.n184 B.n181 10.6151
R1075 B.n185 B.n184 10.6151
R1076 B.n188 B.n185 10.6151
R1077 B.n189 B.n188 10.6151
R1078 B.n192 B.n189 10.6151
R1079 B.n193 B.n192 10.6151
R1080 B.n196 B.n193 10.6151
R1081 B.n197 B.n196 10.6151
R1082 B.n200 B.n197 10.6151
R1083 B.n201 B.n200 10.6151
R1084 B.n204 B.n201 10.6151
R1085 B.n205 B.n204 10.6151
R1086 B.n208 B.n205 10.6151
R1087 B.n209 B.n208 10.6151
R1088 B.n212 B.n209 10.6151
R1089 B.n217 B.n214 10.6151
R1090 B.n218 B.n217 10.6151
R1091 B.n221 B.n218 10.6151
R1092 B.n222 B.n221 10.6151
R1093 B.n225 B.n222 10.6151
R1094 B.n226 B.n225 10.6151
R1095 B.n229 B.n226 10.6151
R1096 B.n230 B.n229 10.6151
R1097 B.n233 B.n230 10.6151
R1098 B.n238 B.n235 10.6151
R1099 B.n239 B.n238 10.6151
R1100 B.n242 B.n239 10.6151
R1101 B.n243 B.n242 10.6151
R1102 B.n246 B.n243 10.6151
R1103 B.n247 B.n246 10.6151
R1104 B.n250 B.n247 10.6151
R1105 B.n251 B.n250 10.6151
R1106 B.n254 B.n251 10.6151
R1107 B.n255 B.n254 10.6151
R1108 B.n258 B.n255 10.6151
R1109 B.n259 B.n258 10.6151
R1110 B.n262 B.n259 10.6151
R1111 B.n263 B.n262 10.6151
R1112 B.n266 B.n263 10.6151
R1113 B.n267 B.n266 10.6151
R1114 B.n270 B.n267 10.6151
R1115 B.n271 B.n270 10.6151
R1116 B.n274 B.n271 10.6151
R1117 B.n275 B.n274 10.6151
R1118 B.n278 B.n275 10.6151
R1119 B.n279 B.n278 10.6151
R1120 B.n282 B.n279 10.6151
R1121 B.n283 B.n282 10.6151
R1122 B.n286 B.n283 10.6151
R1123 B.n287 B.n286 10.6151
R1124 B.n290 B.n287 10.6151
R1125 B.n291 B.n290 10.6151
R1126 B.n294 B.n291 10.6151
R1127 B.n295 B.n294 10.6151
R1128 B.n298 B.n295 10.6151
R1129 B.n299 B.n298 10.6151
R1130 B.n302 B.n299 10.6151
R1131 B.n303 B.n302 10.6151
R1132 B.n306 B.n303 10.6151
R1133 B.n307 B.n306 10.6151
R1134 B.n310 B.n307 10.6151
R1135 B.n311 B.n310 10.6151
R1136 B.n314 B.n311 10.6151
R1137 B.n315 B.n314 10.6151
R1138 B.n318 B.n315 10.6151
R1139 B.n319 B.n318 10.6151
R1140 B.n322 B.n319 10.6151
R1141 B.n323 B.n322 10.6151
R1142 B.n326 B.n323 10.6151
R1143 B.n327 B.n326 10.6151
R1144 B.n330 B.n327 10.6151
R1145 B.n331 B.n330 10.6151
R1146 B.n334 B.n331 10.6151
R1147 B.n335 B.n334 10.6151
R1148 B.n338 B.n335 10.6151
R1149 B.n340 B.n338 10.6151
R1150 B.n341 B.n340 10.6151
R1151 B.n771 B.n341 10.6151
R1152 B.n684 B.n374 10.6151
R1153 B.n694 B.n374 10.6151
R1154 B.n695 B.n694 10.6151
R1155 B.n696 B.n695 10.6151
R1156 B.n696 B.n366 10.6151
R1157 B.n706 B.n366 10.6151
R1158 B.n707 B.n706 10.6151
R1159 B.n708 B.n707 10.6151
R1160 B.n708 B.n358 10.6151
R1161 B.n718 B.n358 10.6151
R1162 B.n719 B.n718 10.6151
R1163 B.n720 B.n719 10.6151
R1164 B.n720 B.n349 10.6151
R1165 B.n730 B.n349 10.6151
R1166 B.n731 B.n730 10.6151
R1167 B.n733 B.n731 10.6151
R1168 B.n733 B.n732 10.6151
R1169 B.n732 B.n342 10.6151
R1170 B.n744 B.n342 10.6151
R1171 B.n745 B.n744 10.6151
R1172 B.n746 B.n745 10.6151
R1173 B.n747 B.n746 10.6151
R1174 B.n749 B.n747 10.6151
R1175 B.n750 B.n749 10.6151
R1176 B.n751 B.n750 10.6151
R1177 B.n752 B.n751 10.6151
R1178 B.n754 B.n752 10.6151
R1179 B.n755 B.n754 10.6151
R1180 B.n756 B.n755 10.6151
R1181 B.n757 B.n756 10.6151
R1182 B.n759 B.n757 10.6151
R1183 B.n760 B.n759 10.6151
R1184 B.n761 B.n760 10.6151
R1185 B.n762 B.n761 10.6151
R1186 B.n764 B.n762 10.6151
R1187 B.n765 B.n764 10.6151
R1188 B.n766 B.n765 10.6151
R1189 B.n767 B.n766 10.6151
R1190 B.n769 B.n767 10.6151
R1191 B.n770 B.n769 10.6151
R1192 B.n448 B.n378 10.6151
R1193 B.n449 B.n448 10.6151
R1194 B.n450 B.n449 10.6151
R1195 B.n450 B.n444 10.6151
R1196 B.n456 B.n444 10.6151
R1197 B.n457 B.n456 10.6151
R1198 B.n458 B.n457 10.6151
R1199 B.n458 B.n442 10.6151
R1200 B.n464 B.n442 10.6151
R1201 B.n465 B.n464 10.6151
R1202 B.n466 B.n465 10.6151
R1203 B.n466 B.n440 10.6151
R1204 B.n472 B.n440 10.6151
R1205 B.n473 B.n472 10.6151
R1206 B.n474 B.n473 10.6151
R1207 B.n474 B.n438 10.6151
R1208 B.n480 B.n438 10.6151
R1209 B.n481 B.n480 10.6151
R1210 B.n482 B.n481 10.6151
R1211 B.n482 B.n436 10.6151
R1212 B.n488 B.n436 10.6151
R1213 B.n489 B.n488 10.6151
R1214 B.n490 B.n489 10.6151
R1215 B.n490 B.n434 10.6151
R1216 B.n496 B.n434 10.6151
R1217 B.n497 B.n496 10.6151
R1218 B.n498 B.n497 10.6151
R1219 B.n498 B.n432 10.6151
R1220 B.n504 B.n432 10.6151
R1221 B.n505 B.n504 10.6151
R1222 B.n506 B.n505 10.6151
R1223 B.n506 B.n430 10.6151
R1224 B.n512 B.n430 10.6151
R1225 B.n513 B.n512 10.6151
R1226 B.n514 B.n513 10.6151
R1227 B.n514 B.n428 10.6151
R1228 B.n520 B.n428 10.6151
R1229 B.n521 B.n520 10.6151
R1230 B.n522 B.n521 10.6151
R1231 B.n522 B.n426 10.6151
R1232 B.n528 B.n426 10.6151
R1233 B.n529 B.n528 10.6151
R1234 B.n530 B.n529 10.6151
R1235 B.n530 B.n424 10.6151
R1236 B.n536 B.n424 10.6151
R1237 B.n537 B.n536 10.6151
R1238 B.n538 B.n537 10.6151
R1239 B.n538 B.n422 10.6151
R1240 B.n544 B.n422 10.6151
R1241 B.n545 B.n544 10.6151
R1242 B.n546 B.n545 10.6151
R1243 B.n546 B.n420 10.6151
R1244 B.n552 B.n420 10.6151
R1245 B.n553 B.n552 10.6151
R1246 B.n555 B.n416 10.6151
R1247 B.n561 B.n416 10.6151
R1248 B.n562 B.n561 10.6151
R1249 B.n563 B.n562 10.6151
R1250 B.n563 B.n414 10.6151
R1251 B.n569 B.n414 10.6151
R1252 B.n570 B.n569 10.6151
R1253 B.n571 B.n570 10.6151
R1254 B.n571 B.n412 10.6151
R1255 B.n578 B.n577 10.6151
R1256 B.n579 B.n578 10.6151
R1257 B.n579 B.n407 10.6151
R1258 B.n585 B.n407 10.6151
R1259 B.n586 B.n585 10.6151
R1260 B.n587 B.n586 10.6151
R1261 B.n587 B.n405 10.6151
R1262 B.n593 B.n405 10.6151
R1263 B.n594 B.n593 10.6151
R1264 B.n595 B.n594 10.6151
R1265 B.n595 B.n403 10.6151
R1266 B.n601 B.n403 10.6151
R1267 B.n602 B.n601 10.6151
R1268 B.n603 B.n602 10.6151
R1269 B.n603 B.n401 10.6151
R1270 B.n609 B.n401 10.6151
R1271 B.n610 B.n609 10.6151
R1272 B.n611 B.n610 10.6151
R1273 B.n611 B.n399 10.6151
R1274 B.n617 B.n399 10.6151
R1275 B.n618 B.n617 10.6151
R1276 B.n619 B.n618 10.6151
R1277 B.n619 B.n397 10.6151
R1278 B.n625 B.n397 10.6151
R1279 B.n626 B.n625 10.6151
R1280 B.n627 B.n626 10.6151
R1281 B.n627 B.n395 10.6151
R1282 B.n633 B.n395 10.6151
R1283 B.n634 B.n633 10.6151
R1284 B.n635 B.n634 10.6151
R1285 B.n635 B.n393 10.6151
R1286 B.n641 B.n393 10.6151
R1287 B.n642 B.n641 10.6151
R1288 B.n643 B.n642 10.6151
R1289 B.n643 B.n391 10.6151
R1290 B.n649 B.n391 10.6151
R1291 B.n650 B.n649 10.6151
R1292 B.n651 B.n650 10.6151
R1293 B.n651 B.n389 10.6151
R1294 B.n657 B.n389 10.6151
R1295 B.n658 B.n657 10.6151
R1296 B.n659 B.n658 10.6151
R1297 B.n659 B.n387 10.6151
R1298 B.n665 B.n387 10.6151
R1299 B.n666 B.n665 10.6151
R1300 B.n667 B.n666 10.6151
R1301 B.n667 B.n385 10.6151
R1302 B.n673 B.n385 10.6151
R1303 B.n674 B.n673 10.6151
R1304 B.n675 B.n674 10.6151
R1305 B.n675 B.n383 10.6151
R1306 B.n383 B.n382 10.6151
R1307 B.n682 B.n382 10.6151
R1308 B.n683 B.n682 10.6151
R1309 B.n689 B.n688 10.6151
R1310 B.n690 B.n689 10.6151
R1311 B.n690 B.n370 10.6151
R1312 B.n700 B.n370 10.6151
R1313 B.n701 B.n700 10.6151
R1314 B.n702 B.n701 10.6151
R1315 B.n702 B.n362 10.6151
R1316 B.n712 B.n362 10.6151
R1317 B.n713 B.n712 10.6151
R1318 B.n714 B.n713 10.6151
R1319 B.n714 B.n354 10.6151
R1320 B.n724 B.n354 10.6151
R1321 B.n725 B.n724 10.6151
R1322 B.n726 B.n725 10.6151
R1323 B.n726 B.n346 10.6151
R1324 B.n737 B.n346 10.6151
R1325 B.n738 B.n737 10.6151
R1326 B.n739 B.n738 10.6151
R1327 B.n739 B.n0 10.6151
R1328 B.n811 B.n1 10.6151
R1329 B.n811 B.n810 10.6151
R1330 B.n810 B.n809 10.6151
R1331 B.n809 B.n10 10.6151
R1332 B.n803 B.n10 10.6151
R1333 B.n803 B.n802 10.6151
R1334 B.n802 B.n801 10.6151
R1335 B.n801 B.n17 10.6151
R1336 B.n795 B.n17 10.6151
R1337 B.n795 B.n794 10.6151
R1338 B.n794 B.n793 10.6151
R1339 B.n793 B.n24 10.6151
R1340 B.n787 B.n24 10.6151
R1341 B.n787 B.n786 10.6151
R1342 B.n786 B.n785 10.6151
R1343 B.n785 B.n31 10.6151
R1344 B.n779 B.n31 10.6151
R1345 B.n779 B.n778 10.6151
R1346 B.n778 B.n777 10.6151
R1347 B.n213 B.n212 9.36635
R1348 B.n235 B.n234 9.36635
R1349 B.n554 B.n553 9.36635
R1350 B.n577 B.n411 9.36635
R1351 B.n704 B.t7 6.54662
R1352 B.t3 B.n789 6.54662
R1353 B.n817 B.n0 2.81026
R1354 B.n817 B.n1 2.81026
R1355 B.n214 B.n213 1.24928
R1356 B.n234 B.n233 1.24928
R1357 B.n555 B.n554 1.24928
R1358 B.n412 B.n411 1.24928
R1359 VP.n0 VP.t1 338.149
R1360 VP.n0 VP.t0 292.392
R1361 VP VP.n0 0.241678
R1362 VTAIL.n1 VTAIL.t1 47.787
R1363 VTAIL.n3 VTAIL.t0 47.7868
R1364 VTAIL.n0 VTAIL.t2 47.7868
R1365 VTAIL.n2 VTAIL.t3 47.7868
R1366 VTAIL.n1 VTAIL.n0 30.1686
R1367 VTAIL.n3 VTAIL.n2 28.41
R1368 VTAIL.n2 VTAIL.n1 1.34964
R1369 VTAIL VTAIL.n0 0.968172
R1370 VTAIL VTAIL.n3 0.381966
R1371 VDD1 VDD1.t1 106.891
R1372 VDD1 VDD1.t0 64.9634
R1373 VN VN.t0 338.341
R1374 VN VN.t1 292.632
R1375 VDD2.n0 VDD2.t0 105.927
R1376 VDD2.n0 VDD2.t1 64.4655
R1377 VDD2 VDD2.n0 0.498345
C0 VTAIL VP 2.88275f
C1 VDD1 VDD2 0.570668f
C2 VDD1 VN 0.147714f
C3 VDD1 VTAIL 6.3462f
C4 VDD2 VN 3.46192f
C5 VDD1 VP 3.60626f
C6 VDD2 VTAIL 6.38806f
C7 VTAIL VN 2.86826f
C8 VDD2 VP 0.296251f
C9 VN VP 5.88671f
C10 VDD2 B 4.940475f
C11 VDD1 B 8.21898f
C12 VTAIL B 8.714002f
C13 VN B 11.11537f
C14 VP B 5.609659f
C15 VDD2.t0 B 3.66873f
C16 VDD2.t1 B 3.0569f
C17 VDD2.n0 B 3.08461f
C18 VN.t1 B 3.22745f
C19 VN.t0 B 3.62024f
C20 VDD1.t0 B 3.0361f
C21 VDD1.t1 B 3.67363f
C22 VTAIL.t2 B 2.93352f
C23 VTAIL.n0 B 1.72319f
C24 VTAIL.t1 B 2.93352f
C25 VTAIL.n1 B 1.74749f
C26 VTAIL.t3 B 2.93352f
C27 VTAIL.n2 B 1.63547f
C28 VTAIL.t0 B 2.93352f
C29 VTAIL.n3 B 1.57382f
C30 VP.t1 B 3.66191f
C31 VP.t0 B 3.26708f
C32 VP.n0 B 5.41483f
.ends

