* NGSPICE file created from diff_pair_sample_0799.ext - technology: sky130A

.subckt diff_pair_sample_0799 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n2650_n1878# sky130_fd_pr__pfet_01v8 ad=1.7745 pd=9.88 as=0 ps=0 w=4.55 l=1.35
X1 B.t8 B.t6 B.t7 w_n2650_n1878# sky130_fd_pr__pfet_01v8 ad=1.7745 pd=9.88 as=0 ps=0 w=4.55 l=1.35
X2 VDD2.t7 VN.t0 VTAIL.t13 w_n2650_n1878# sky130_fd_pr__pfet_01v8 ad=0.75075 pd=4.88 as=1.7745 ps=9.88 w=4.55 l=1.35
X3 VTAIL.t6 VP.t0 VDD1.t7 w_n2650_n1878# sky130_fd_pr__pfet_01v8 ad=1.7745 pd=9.88 as=0.75075 ps=4.88 w=4.55 l=1.35
X4 VDD1.t6 VP.t1 VTAIL.t5 w_n2650_n1878# sky130_fd_pr__pfet_01v8 ad=0.75075 pd=4.88 as=0.75075 ps=4.88 w=4.55 l=1.35
X5 VDD2.t6 VN.t1 VTAIL.t11 w_n2650_n1878# sky130_fd_pr__pfet_01v8 ad=0.75075 pd=4.88 as=1.7745 ps=9.88 w=4.55 l=1.35
X6 B.t5 B.t3 B.t4 w_n2650_n1878# sky130_fd_pr__pfet_01v8 ad=1.7745 pd=9.88 as=0 ps=0 w=4.55 l=1.35
X7 B.t2 B.t0 B.t1 w_n2650_n1878# sky130_fd_pr__pfet_01v8 ad=1.7745 pd=9.88 as=0 ps=0 w=4.55 l=1.35
X8 VDD2.t5 VN.t2 VTAIL.t9 w_n2650_n1878# sky130_fd_pr__pfet_01v8 ad=0.75075 pd=4.88 as=0.75075 ps=4.88 w=4.55 l=1.35
X9 VTAIL.t15 VN.t3 VDD2.t4 w_n2650_n1878# sky130_fd_pr__pfet_01v8 ad=1.7745 pd=9.88 as=0.75075 ps=4.88 w=4.55 l=1.35
X10 VDD1.t5 VP.t2 VTAIL.t2 w_n2650_n1878# sky130_fd_pr__pfet_01v8 ad=0.75075 pd=4.88 as=1.7745 ps=9.88 w=4.55 l=1.35
X11 VTAIL.t8 VN.t4 VDD2.t3 w_n2650_n1878# sky130_fd_pr__pfet_01v8 ad=0.75075 pd=4.88 as=0.75075 ps=4.88 w=4.55 l=1.35
X12 VDD1.t4 VP.t3 VTAIL.t4 w_n2650_n1878# sky130_fd_pr__pfet_01v8 ad=0.75075 pd=4.88 as=0.75075 ps=4.88 w=4.55 l=1.35
X13 VDD2.t2 VN.t5 VTAIL.t14 w_n2650_n1878# sky130_fd_pr__pfet_01v8 ad=0.75075 pd=4.88 as=0.75075 ps=4.88 w=4.55 l=1.35
X14 VDD1.t3 VP.t4 VTAIL.t3 w_n2650_n1878# sky130_fd_pr__pfet_01v8 ad=0.75075 pd=4.88 as=1.7745 ps=9.88 w=4.55 l=1.35
X15 VTAIL.t12 VN.t6 VDD2.t1 w_n2650_n1878# sky130_fd_pr__pfet_01v8 ad=0.75075 pd=4.88 as=0.75075 ps=4.88 w=4.55 l=1.35
X16 VTAIL.t7 VP.t5 VDD1.t2 w_n2650_n1878# sky130_fd_pr__pfet_01v8 ad=0.75075 pd=4.88 as=0.75075 ps=4.88 w=4.55 l=1.35
X17 VTAIL.t10 VN.t7 VDD2.t0 w_n2650_n1878# sky130_fd_pr__pfet_01v8 ad=1.7745 pd=9.88 as=0.75075 ps=4.88 w=4.55 l=1.35
X18 VTAIL.t1 VP.t6 VDD1.t1 w_n2650_n1878# sky130_fd_pr__pfet_01v8 ad=0.75075 pd=4.88 as=0.75075 ps=4.88 w=4.55 l=1.35
X19 VTAIL.t0 VP.t7 VDD1.t0 w_n2650_n1878# sky130_fd_pr__pfet_01v8 ad=1.7745 pd=9.88 as=0.75075 ps=4.88 w=4.55 l=1.35
R0 B.n351 B.n350 585
R1 B.n352 B.n47 585
R2 B.n354 B.n353 585
R3 B.n355 B.n46 585
R4 B.n357 B.n356 585
R5 B.n358 B.n45 585
R6 B.n360 B.n359 585
R7 B.n361 B.n44 585
R8 B.n363 B.n362 585
R9 B.n364 B.n43 585
R10 B.n366 B.n365 585
R11 B.n367 B.n42 585
R12 B.n369 B.n368 585
R13 B.n370 B.n41 585
R14 B.n372 B.n371 585
R15 B.n373 B.n40 585
R16 B.n375 B.n374 585
R17 B.n376 B.n39 585
R18 B.n378 B.n377 585
R19 B.n379 B.n36 585
R20 B.n382 B.n381 585
R21 B.n383 B.n35 585
R22 B.n385 B.n384 585
R23 B.n386 B.n34 585
R24 B.n388 B.n387 585
R25 B.n389 B.n33 585
R26 B.n391 B.n390 585
R27 B.n392 B.n29 585
R28 B.n394 B.n393 585
R29 B.n395 B.n28 585
R30 B.n397 B.n396 585
R31 B.n398 B.n27 585
R32 B.n400 B.n399 585
R33 B.n401 B.n26 585
R34 B.n403 B.n402 585
R35 B.n404 B.n25 585
R36 B.n406 B.n405 585
R37 B.n407 B.n24 585
R38 B.n409 B.n408 585
R39 B.n410 B.n23 585
R40 B.n412 B.n411 585
R41 B.n413 B.n22 585
R42 B.n415 B.n414 585
R43 B.n416 B.n21 585
R44 B.n418 B.n417 585
R45 B.n419 B.n20 585
R46 B.n421 B.n420 585
R47 B.n422 B.n19 585
R48 B.n424 B.n423 585
R49 B.n349 B.n48 585
R50 B.n348 B.n347 585
R51 B.n346 B.n49 585
R52 B.n345 B.n344 585
R53 B.n343 B.n50 585
R54 B.n342 B.n341 585
R55 B.n340 B.n51 585
R56 B.n339 B.n338 585
R57 B.n337 B.n52 585
R58 B.n336 B.n335 585
R59 B.n334 B.n53 585
R60 B.n333 B.n332 585
R61 B.n331 B.n54 585
R62 B.n330 B.n329 585
R63 B.n328 B.n55 585
R64 B.n327 B.n326 585
R65 B.n325 B.n56 585
R66 B.n324 B.n323 585
R67 B.n322 B.n57 585
R68 B.n321 B.n320 585
R69 B.n319 B.n58 585
R70 B.n318 B.n317 585
R71 B.n316 B.n59 585
R72 B.n315 B.n314 585
R73 B.n313 B.n60 585
R74 B.n312 B.n311 585
R75 B.n310 B.n61 585
R76 B.n309 B.n308 585
R77 B.n307 B.n62 585
R78 B.n306 B.n305 585
R79 B.n304 B.n63 585
R80 B.n303 B.n302 585
R81 B.n301 B.n64 585
R82 B.n300 B.n299 585
R83 B.n298 B.n65 585
R84 B.n297 B.n296 585
R85 B.n295 B.n66 585
R86 B.n294 B.n293 585
R87 B.n292 B.n67 585
R88 B.n291 B.n290 585
R89 B.n289 B.n68 585
R90 B.n288 B.n287 585
R91 B.n286 B.n69 585
R92 B.n285 B.n284 585
R93 B.n283 B.n70 585
R94 B.n282 B.n281 585
R95 B.n280 B.n71 585
R96 B.n279 B.n278 585
R97 B.n277 B.n72 585
R98 B.n276 B.n275 585
R99 B.n274 B.n73 585
R100 B.n273 B.n272 585
R101 B.n271 B.n74 585
R102 B.n270 B.n269 585
R103 B.n268 B.n75 585
R104 B.n267 B.n266 585
R105 B.n265 B.n76 585
R106 B.n264 B.n263 585
R107 B.n262 B.n77 585
R108 B.n261 B.n260 585
R109 B.n259 B.n78 585
R110 B.n258 B.n257 585
R111 B.n256 B.n79 585
R112 B.n255 B.n254 585
R113 B.n253 B.n80 585
R114 B.n252 B.n251 585
R115 B.n250 B.n81 585
R116 B.n173 B.n172 585
R117 B.n174 B.n107 585
R118 B.n176 B.n175 585
R119 B.n177 B.n106 585
R120 B.n179 B.n178 585
R121 B.n180 B.n105 585
R122 B.n182 B.n181 585
R123 B.n183 B.n104 585
R124 B.n185 B.n184 585
R125 B.n186 B.n103 585
R126 B.n188 B.n187 585
R127 B.n189 B.n102 585
R128 B.n191 B.n190 585
R129 B.n192 B.n101 585
R130 B.n194 B.n193 585
R131 B.n195 B.n100 585
R132 B.n197 B.n196 585
R133 B.n198 B.n99 585
R134 B.n200 B.n199 585
R135 B.n201 B.n96 585
R136 B.n204 B.n203 585
R137 B.n205 B.n95 585
R138 B.n207 B.n206 585
R139 B.n208 B.n94 585
R140 B.n210 B.n209 585
R141 B.n211 B.n93 585
R142 B.n213 B.n212 585
R143 B.n214 B.n92 585
R144 B.n219 B.n218 585
R145 B.n220 B.n91 585
R146 B.n222 B.n221 585
R147 B.n223 B.n90 585
R148 B.n225 B.n224 585
R149 B.n226 B.n89 585
R150 B.n228 B.n227 585
R151 B.n229 B.n88 585
R152 B.n231 B.n230 585
R153 B.n232 B.n87 585
R154 B.n234 B.n233 585
R155 B.n235 B.n86 585
R156 B.n237 B.n236 585
R157 B.n238 B.n85 585
R158 B.n240 B.n239 585
R159 B.n241 B.n84 585
R160 B.n243 B.n242 585
R161 B.n244 B.n83 585
R162 B.n246 B.n245 585
R163 B.n247 B.n82 585
R164 B.n249 B.n248 585
R165 B.n171 B.n108 585
R166 B.n170 B.n169 585
R167 B.n168 B.n109 585
R168 B.n167 B.n166 585
R169 B.n165 B.n110 585
R170 B.n164 B.n163 585
R171 B.n162 B.n111 585
R172 B.n161 B.n160 585
R173 B.n159 B.n112 585
R174 B.n158 B.n157 585
R175 B.n156 B.n113 585
R176 B.n155 B.n154 585
R177 B.n153 B.n114 585
R178 B.n152 B.n151 585
R179 B.n150 B.n115 585
R180 B.n149 B.n148 585
R181 B.n147 B.n116 585
R182 B.n146 B.n145 585
R183 B.n144 B.n117 585
R184 B.n143 B.n142 585
R185 B.n141 B.n118 585
R186 B.n140 B.n139 585
R187 B.n138 B.n119 585
R188 B.n137 B.n136 585
R189 B.n135 B.n120 585
R190 B.n134 B.n133 585
R191 B.n132 B.n121 585
R192 B.n131 B.n130 585
R193 B.n129 B.n122 585
R194 B.n128 B.n127 585
R195 B.n126 B.n123 585
R196 B.n125 B.n124 585
R197 B.n2 B.n0 585
R198 B.n473 B.n1 585
R199 B.n472 B.n471 585
R200 B.n470 B.n3 585
R201 B.n469 B.n468 585
R202 B.n467 B.n4 585
R203 B.n466 B.n465 585
R204 B.n464 B.n5 585
R205 B.n463 B.n462 585
R206 B.n461 B.n6 585
R207 B.n460 B.n459 585
R208 B.n458 B.n7 585
R209 B.n457 B.n456 585
R210 B.n455 B.n8 585
R211 B.n454 B.n453 585
R212 B.n452 B.n9 585
R213 B.n451 B.n450 585
R214 B.n449 B.n10 585
R215 B.n448 B.n447 585
R216 B.n446 B.n11 585
R217 B.n445 B.n444 585
R218 B.n443 B.n12 585
R219 B.n442 B.n441 585
R220 B.n440 B.n13 585
R221 B.n439 B.n438 585
R222 B.n437 B.n14 585
R223 B.n436 B.n435 585
R224 B.n434 B.n15 585
R225 B.n433 B.n432 585
R226 B.n431 B.n16 585
R227 B.n430 B.n429 585
R228 B.n428 B.n17 585
R229 B.n427 B.n426 585
R230 B.n425 B.n18 585
R231 B.n475 B.n474 585
R232 B.n173 B.n108 468.476
R233 B.n425 B.n424 468.476
R234 B.n250 B.n249 468.476
R235 B.n351 B.n48 468.476
R236 B.n215 B.t3 286.06
R237 B.n97 B.t6 286.06
R238 B.n30 B.t0 286.06
R239 B.n37 B.t9 286.06
R240 B.n215 B.t5 275.957
R241 B.n37 B.t10 275.957
R242 B.n97 B.t8 275.957
R243 B.n30 B.t1 275.957
R244 B.n216 B.t4 243.375
R245 B.n38 B.t11 243.375
R246 B.n98 B.t7 243.375
R247 B.n31 B.t2 243.375
R248 B.n169 B.n108 163.367
R249 B.n169 B.n168 163.367
R250 B.n168 B.n167 163.367
R251 B.n167 B.n110 163.367
R252 B.n163 B.n110 163.367
R253 B.n163 B.n162 163.367
R254 B.n162 B.n161 163.367
R255 B.n161 B.n112 163.367
R256 B.n157 B.n112 163.367
R257 B.n157 B.n156 163.367
R258 B.n156 B.n155 163.367
R259 B.n155 B.n114 163.367
R260 B.n151 B.n114 163.367
R261 B.n151 B.n150 163.367
R262 B.n150 B.n149 163.367
R263 B.n149 B.n116 163.367
R264 B.n145 B.n116 163.367
R265 B.n145 B.n144 163.367
R266 B.n144 B.n143 163.367
R267 B.n143 B.n118 163.367
R268 B.n139 B.n118 163.367
R269 B.n139 B.n138 163.367
R270 B.n138 B.n137 163.367
R271 B.n137 B.n120 163.367
R272 B.n133 B.n120 163.367
R273 B.n133 B.n132 163.367
R274 B.n132 B.n131 163.367
R275 B.n131 B.n122 163.367
R276 B.n127 B.n122 163.367
R277 B.n127 B.n126 163.367
R278 B.n126 B.n125 163.367
R279 B.n125 B.n2 163.367
R280 B.n474 B.n2 163.367
R281 B.n474 B.n473 163.367
R282 B.n473 B.n472 163.367
R283 B.n472 B.n3 163.367
R284 B.n468 B.n3 163.367
R285 B.n468 B.n467 163.367
R286 B.n467 B.n466 163.367
R287 B.n466 B.n5 163.367
R288 B.n462 B.n5 163.367
R289 B.n462 B.n461 163.367
R290 B.n461 B.n460 163.367
R291 B.n460 B.n7 163.367
R292 B.n456 B.n7 163.367
R293 B.n456 B.n455 163.367
R294 B.n455 B.n454 163.367
R295 B.n454 B.n9 163.367
R296 B.n450 B.n9 163.367
R297 B.n450 B.n449 163.367
R298 B.n449 B.n448 163.367
R299 B.n448 B.n11 163.367
R300 B.n444 B.n11 163.367
R301 B.n444 B.n443 163.367
R302 B.n443 B.n442 163.367
R303 B.n442 B.n13 163.367
R304 B.n438 B.n13 163.367
R305 B.n438 B.n437 163.367
R306 B.n437 B.n436 163.367
R307 B.n436 B.n15 163.367
R308 B.n432 B.n15 163.367
R309 B.n432 B.n431 163.367
R310 B.n431 B.n430 163.367
R311 B.n430 B.n17 163.367
R312 B.n426 B.n17 163.367
R313 B.n426 B.n425 163.367
R314 B.n174 B.n173 163.367
R315 B.n175 B.n174 163.367
R316 B.n175 B.n106 163.367
R317 B.n179 B.n106 163.367
R318 B.n180 B.n179 163.367
R319 B.n181 B.n180 163.367
R320 B.n181 B.n104 163.367
R321 B.n185 B.n104 163.367
R322 B.n186 B.n185 163.367
R323 B.n187 B.n186 163.367
R324 B.n187 B.n102 163.367
R325 B.n191 B.n102 163.367
R326 B.n192 B.n191 163.367
R327 B.n193 B.n192 163.367
R328 B.n193 B.n100 163.367
R329 B.n197 B.n100 163.367
R330 B.n198 B.n197 163.367
R331 B.n199 B.n198 163.367
R332 B.n199 B.n96 163.367
R333 B.n204 B.n96 163.367
R334 B.n205 B.n204 163.367
R335 B.n206 B.n205 163.367
R336 B.n206 B.n94 163.367
R337 B.n210 B.n94 163.367
R338 B.n211 B.n210 163.367
R339 B.n212 B.n211 163.367
R340 B.n212 B.n92 163.367
R341 B.n219 B.n92 163.367
R342 B.n220 B.n219 163.367
R343 B.n221 B.n220 163.367
R344 B.n221 B.n90 163.367
R345 B.n225 B.n90 163.367
R346 B.n226 B.n225 163.367
R347 B.n227 B.n226 163.367
R348 B.n227 B.n88 163.367
R349 B.n231 B.n88 163.367
R350 B.n232 B.n231 163.367
R351 B.n233 B.n232 163.367
R352 B.n233 B.n86 163.367
R353 B.n237 B.n86 163.367
R354 B.n238 B.n237 163.367
R355 B.n239 B.n238 163.367
R356 B.n239 B.n84 163.367
R357 B.n243 B.n84 163.367
R358 B.n244 B.n243 163.367
R359 B.n245 B.n244 163.367
R360 B.n245 B.n82 163.367
R361 B.n249 B.n82 163.367
R362 B.n251 B.n250 163.367
R363 B.n251 B.n80 163.367
R364 B.n255 B.n80 163.367
R365 B.n256 B.n255 163.367
R366 B.n257 B.n256 163.367
R367 B.n257 B.n78 163.367
R368 B.n261 B.n78 163.367
R369 B.n262 B.n261 163.367
R370 B.n263 B.n262 163.367
R371 B.n263 B.n76 163.367
R372 B.n267 B.n76 163.367
R373 B.n268 B.n267 163.367
R374 B.n269 B.n268 163.367
R375 B.n269 B.n74 163.367
R376 B.n273 B.n74 163.367
R377 B.n274 B.n273 163.367
R378 B.n275 B.n274 163.367
R379 B.n275 B.n72 163.367
R380 B.n279 B.n72 163.367
R381 B.n280 B.n279 163.367
R382 B.n281 B.n280 163.367
R383 B.n281 B.n70 163.367
R384 B.n285 B.n70 163.367
R385 B.n286 B.n285 163.367
R386 B.n287 B.n286 163.367
R387 B.n287 B.n68 163.367
R388 B.n291 B.n68 163.367
R389 B.n292 B.n291 163.367
R390 B.n293 B.n292 163.367
R391 B.n293 B.n66 163.367
R392 B.n297 B.n66 163.367
R393 B.n298 B.n297 163.367
R394 B.n299 B.n298 163.367
R395 B.n299 B.n64 163.367
R396 B.n303 B.n64 163.367
R397 B.n304 B.n303 163.367
R398 B.n305 B.n304 163.367
R399 B.n305 B.n62 163.367
R400 B.n309 B.n62 163.367
R401 B.n310 B.n309 163.367
R402 B.n311 B.n310 163.367
R403 B.n311 B.n60 163.367
R404 B.n315 B.n60 163.367
R405 B.n316 B.n315 163.367
R406 B.n317 B.n316 163.367
R407 B.n317 B.n58 163.367
R408 B.n321 B.n58 163.367
R409 B.n322 B.n321 163.367
R410 B.n323 B.n322 163.367
R411 B.n323 B.n56 163.367
R412 B.n327 B.n56 163.367
R413 B.n328 B.n327 163.367
R414 B.n329 B.n328 163.367
R415 B.n329 B.n54 163.367
R416 B.n333 B.n54 163.367
R417 B.n334 B.n333 163.367
R418 B.n335 B.n334 163.367
R419 B.n335 B.n52 163.367
R420 B.n339 B.n52 163.367
R421 B.n340 B.n339 163.367
R422 B.n341 B.n340 163.367
R423 B.n341 B.n50 163.367
R424 B.n345 B.n50 163.367
R425 B.n346 B.n345 163.367
R426 B.n347 B.n346 163.367
R427 B.n347 B.n48 163.367
R428 B.n424 B.n19 163.367
R429 B.n420 B.n19 163.367
R430 B.n420 B.n419 163.367
R431 B.n419 B.n418 163.367
R432 B.n418 B.n21 163.367
R433 B.n414 B.n21 163.367
R434 B.n414 B.n413 163.367
R435 B.n413 B.n412 163.367
R436 B.n412 B.n23 163.367
R437 B.n408 B.n23 163.367
R438 B.n408 B.n407 163.367
R439 B.n407 B.n406 163.367
R440 B.n406 B.n25 163.367
R441 B.n402 B.n25 163.367
R442 B.n402 B.n401 163.367
R443 B.n401 B.n400 163.367
R444 B.n400 B.n27 163.367
R445 B.n396 B.n27 163.367
R446 B.n396 B.n395 163.367
R447 B.n395 B.n394 163.367
R448 B.n394 B.n29 163.367
R449 B.n390 B.n29 163.367
R450 B.n390 B.n389 163.367
R451 B.n389 B.n388 163.367
R452 B.n388 B.n34 163.367
R453 B.n384 B.n34 163.367
R454 B.n384 B.n383 163.367
R455 B.n383 B.n382 163.367
R456 B.n382 B.n36 163.367
R457 B.n377 B.n36 163.367
R458 B.n377 B.n376 163.367
R459 B.n376 B.n375 163.367
R460 B.n375 B.n40 163.367
R461 B.n371 B.n40 163.367
R462 B.n371 B.n370 163.367
R463 B.n370 B.n369 163.367
R464 B.n369 B.n42 163.367
R465 B.n365 B.n42 163.367
R466 B.n365 B.n364 163.367
R467 B.n364 B.n363 163.367
R468 B.n363 B.n44 163.367
R469 B.n359 B.n44 163.367
R470 B.n359 B.n358 163.367
R471 B.n358 B.n357 163.367
R472 B.n357 B.n46 163.367
R473 B.n353 B.n46 163.367
R474 B.n353 B.n352 163.367
R475 B.n352 B.n351 163.367
R476 B.n217 B.n216 59.5399
R477 B.n202 B.n98 59.5399
R478 B.n32 B.n31 59.5399
R479 B.n380 B.n38 59.5399
R480 B.n216 B.n215 32.5823
R481 B.n98 B.n97 32.5823
R482 B.n31 B.n30 32.5823
R483 B.n38 B.n37 32.5823
R484 B.n423 B.n18 30.4395
R485 B.n248 B.n81 30.4395
R486 B.n172 B.n171 30.4395
R487 B.n350 B.n349 30.4395
R488 B B.n475 18.0485
R489 B.n423 B.n422 10.6151
R490 B.n422 B.n421 10.6151
R491 B.n421 B.n20 10.6151
R492 B.n417 B.n20 10.6151
R493 B.n417 B.n416 10.6151
R494 B.n416 B.n415 10.6151
R495 B.n415 B.n22 10.6151
R496 B.n411 B.n22 10.6151
R497 B.n411 B.n410 10.6151
R498 B.n410 B.n409 10.6151
R499 B.n409 B.n24 10.6151
R500 B.n405 B.n24 10.6151
R501 B.n405 B.n404 10.6151
R502 B.n404 B.n403 10.6151
R503 B.n403 B.n26 10.6151
R504 B.n399 B.n26 10.6151
R505 B.n399 B.n398 10.6151
R506 B.n398 B.n397 10.6151
R507 B.n397 B.n28 10.6151
R508 B.n393 B.n392 10.6151
R509 B.n392 B.n391 10.6151
R510 B.n391 B.n33 10.6151
R511 B.n387 B.n33 10.6151
R512 B.n387 B.n386 10.6151
R513 B.n386 B.n385 10.6151
R514 B.n385 B.n35 10.6151
R515 B.n381 B.n35 10.6151
R516 B.n379 B.n378 10.6151
R517 B.n378 B.n39 10.6151
R518 B.n374 B.n39 10.6151
R519 B.n374 B.n373 10.6151
R520 B.n373 B.n372 10.6151
R521 B.n372 B.n41 10.6151
R522 B.n368 B.n41 10.6151
R523 B.n368 B.n367 10.6151
R524 B.n367 B.n366 10.6151
R525 B.n366 B.n43 10.6151
R526 B.n362 B.n43 10.6151
R527 B.n362 B.n361 10.6151
R528 B.n361 B.n360 10.6151
R529 B.n360 B.n45 10.6151
R530 B.n356 B.n45 10.6151
R531 B.n356 B.n355 10.6151
R532 B.n355 B.n354 10.6151
R533 B.n354 B.n47 10.6151
R534 B.n350 B.n47 10.6151
R535 B.n252 B.n81 10.6151
R536 B.n253 B.n252 10.6151
R537 B.n254 B.n253 10.6151
R538 B.n254 B.n79 10.6151
R539 B.n258 B.n79 10.6151
R540 B.n259 B.n258 10.6151
R541 B.n260 B.n259 10.6151
R542 B.n260 B.n77 10.6151
R543 B.n264 B.n77 10.6151
R544 B.n265 B.n264 10.6151
R545 B.n266 B.n265 10.6151
R546 B.n266 B.n75 10.6151
R547 B.n270 B.n75 10.6151
R548 B.n271 B.n270 10.6151
R549 B.n272 B.n271 10.6151
R550 B.n272 B.n73 10.6151
R551 B.n276 B.n73 10.6151
R552 B.n277 B.n276 10.6151
R553 B.n278 B.n277 10.6151
R554 B.n278 B.n71 10.6151
R555 B.n282 B.n71 10.6151
R556 B.n283 B.n282 10.6151
R557 B.n284 B.n283 10.6151
R558 B.n284 B.n69 10.6151
R559 B.n288 B.n69 10.6151
R560 B.n289 B.n288 10.6151
R561 B.n290 B.n289 10.6151
R562 B.n290 B.n67 10.6151
R563 B.n294 B.n67 10.6151
R564 B.n295 B.n294 10.6151
R565 B.n296 B.n295 10.6151
R566 B.n296 B.n65 10.6151
R567 B.n300 B.n65 10.6151
R568 B.n301 B.n300 10.6151
R569 B.n302 B.n301 10.6151
R570 B.n302 B.n63 10.6151
R571 B.n306 B.n63 10.6151
R572 B.n307 B.n306 10.6151
R573 B.n308 B.n307 10.6151
R574 B.n308 B.n61 10.6151
R575 B.n312 B.n61 10.6151
R576 B.n313 B.n312 10.6151
R577 B.n314 B.n313 10.6151
R578 B.n314 B.n59 10.6151
R579 B.n318 B.n59 10.6151
R580 B.n319 B.n318 10.6151
R581 B.n320 B.n319 10.6151
R582 B.n320 B.n57 10.6151
R583 B.n324 B.n57 10.6151
R584 B.n325 B.n324 10.6151
R585 B.n326 B.n325 10.6151
R586 B.n326 B.n55 10.6151
R587 B.n330 B.n55 10.6151
R588 B.n331 B.n330 10.6151
R589 B.n332 B.n331 10.6151
R590 B.n332 B.n53 10.6151
R591 B.n336 B.n53 10.6151
R592 B.n337 B.n336 10.6151
R593 B.n338 B.n337 10.6151
R594 B.n338 B.n51 10.6151
R595 B.n342 B.n51 10.6151
R596 B.n343 B.n342 10.6151
R597 B.n344 B.n343 10.6151
R598 B.n344 B.n49 10.6151
R599 B.n348 B.n49 10.6151
R600 B.n349 B.n348 10.6151
R601 B.n172 B.n107 10.6151
R602 B.n176 B.n107 10.6151
R603 B.n177 B.n176 10.6151
R604 B.n178 B.n177 10.6151
R605 B.n178 B.n105 10.6151
R606 B.n182 B.n105 10.6151
R607 B.n183 B.n182 10.6151
R608 B.n184 B.n183 10.6151
R609 B.n184 B.n103 10.6151
R610 B.n188 B.n103 10.6151
R611 B.n189 B.n188 10.6151
R612 B.n190 B.n189 10.6151
R613 B.n190 B.n101 10.6151
R614 B.n194 B.n101 10.6151
R615 B.n195 B.n194 10.6151
R616 B.n196 B.n195 10.6151
R617 B.n196 B.n99 10.6151
R618 B.n200 B.n99 10.6151
R619 B.n201 B.n200 10.6151
R620 B.n203 B.n95 10.6151
R621 B.n207 B.n95 10.6151
R622 B.n208 B.n207 10.6151
R623 B.n209 B.n208 10.6151
R624 B.n209 B.n93 10.6151
R625 B.n213 B.n93 10.6151
R626 B.n214 B.n213 10.6151
R627 B.n218 B.n214 10.6151
R628 B.n222 B.n91 10.6151
R629 B.n223 B.n222 10.6151
R630 B.n224 B.n223 10.6151
R631 B.n224 B.n89 10.6151
R632 B.n228 B.n89 10.6151
R633 B.n229 B.n228 10.6151
R634 B.n230 B.n229 10.6151
R635 B.n230 B.n87 10.6151
R636 B.n234 B.n87 10.6151
R637 B.n235 B.n234 10.6151
R638 B.n236 B.n235 10.6151
R639 B.n236 B.n85 10.6151
R640 B.n240 B.n85 10.6151
R641 B.n241 B.n240 10.6151
R642 B.n242 B.n241 10.6151
R643 B.n242 B.n83 10.6151
R644 B.n246 B.n83 10.6151
R645 B.n247 B.n246 10.6151
R646 B.n248 B.n247 10.6151
R647 B.n171 B.n170 10.6151
R648 B.n170 B.n109 10.6151
R649 B.n166 B.n109 10.6151
R650 B.n166 B.n165 10.6151
R651 B.n165 B.n164 10.6151
R652 B.n164 B.n111 10.6151
R653 B.n160 B.n111 10.6151
R654 B.n160 B.n159 10.6151
R655 B.n159 B.n158 10.6151
R656 B.n158 B.n113 10.6151
R657 B.n154 B.n113 10.6151
R658 B.n154 B.n153 10.6151
R659 B.n153 B.n152 10.6151
R660 B.n152 B.n115 10.6151
R661 B.n148 B.n115 10.6151
R662 B.n148 B.n147 10.6151
R663 B.n147 B.n146 10.6151
R664 B.n146 B.n117 10.6151
R665 B.n142 B.n117 10.6151
R666 B.n142 B.n141 10.6151
R667 B.n141 B.n140 10.6151
R668 B.n140 B.n119 10.6151
R669 B.n136 B.n119 10.6151
R670 B.n136 B.n135 10.6151
R671 B.n135 B.n134 10.6151
R672 B.n134 B.n121 10.6151
R673 B.n130 B.n121 10.6151
R674 B.n130 B.n129 10.6151
R675 B.n129 B.n128 10.6151
R676 B.n128 B.n123 10.6151
R677 B.n124 B.n123 10.6151
R678 B.n124 B.n0 10.6151
R679 B.n471 B.n1 10.6151
R680 B.n471 B.n470 10.6151
R681 B.n470 B.n469 10.6151
R682 B.n469 B.n4 10.6151
R683 B.n465 B.n4 10.6151
R684 B.n465 B.n464 10.6151
R685 B.n464 B.n463 10.6151
R686 B.n463 B.n6 10.6151
R687 B.n459 B.n6 10.6151
R688 B.n459 B.n458 10.6151
R689 B.n458 B.n457 10.6151
R690 B.n457 B.n8 10.6151
R691 B.n453 B.n8 10.6151
R692 B.n453 B.n452 10.6151
R693 B.n452 B.n451 10.6151
R694 B.n451 B.n10 10.6151
R695 B.n447 B.n10 10.6151
R696 B.n447 B.n446 10.6151
R697 B.n446 B.n445 10.6151
R698 B.n445 B.n12 10.6151
R699 B.n441 B.n12 10.6151
R700 B.n441 B.n440 10.6151
R701 B.n440 B.n439 10.6151
R702 B.n439 B.n14 10.6151
R703 B.n435 B.n14 10.6151
R704 B.n435 B.n434 10.6151
R705 B.n434 B.n433 10.6151
R706 B.n433 B.n16 10.6151
R707 B.n429 B.n16 10.6151
R708 B.n429 B.n428 10.6151
R709 B.n428 B.n427 10.6151
R710 B.n427 B.n18 10.6151
R711 B.n393 B.n32 6.5566
R712 B.n381 B.n380 6.5566
R713 B.n203 B.n202 6.5566
R714 B.n218 B.n217 6.5566
R715 B.n32 B.n28 4.05904
R716 B.n380 B.n379 4.05904
R717 B.n202 B.n201 4.05904
R718 B.n217 B.n91 4.05904
R719 B.n475 B.n0 2.81026
R720 B.n475 B.n1 2.81026
R721 VN.n18 VN.n17 172.555
R722 VN.n37 VN.n36 172.555
R723 VN.n35 VN.n19 161.3
R724 VN.n34 VN.n33 161.3
R725 VN.n32 VN.n20 161.3
R726 VN.n31 VN.n30 161.3
R727 VN.n29 VN.n21 161.3
R728 VN.n28 VN.n27 161.3
R729 VN.n26 VN.n23 161.3
R730 VN.n16 VN.n0 161.3
R731 VN.n15 VN.n14 161.3
R732 VN.n13 VN.n1 161.3
R733 VN.n12 VN.n11 161.3
R734 VN.n9 VN.n2 161.3
R735 VN.n8 VN.n7 161.3
R736 VN.n6 VN.n3 161.3
R737 VN.n5 VN.t3 110.861
R738 VN.n25 VN.t1 110.861
R739 VN.n4 VN.t5 81.2264
R740 VN.n10 VN.t4 81.2264
R741 VN.n17 VN.t0 81.2264
R742 VN.n24 VN.t6 81.2264
R743 VN.n22 VN.t2 81.2264
R744 VN.n36 VN.t7 81.2264
R745 VN.n5 VN.n4 60.7907
R746 VN.n25 VN.n24 60.7907
R747 VN.n9 VN.n8 56.5193
R748 VN.n29 VN.n28 56.5193
R749 VN.n15 VN.n1 47.2923
R750 VN.n34 VN.n20 47.2923
R751 VN VN.n37 39.7221
R752 VN.n16 VN.n15 33.6945
R753 VN.n35 VN.n34 33.6945
R754 VN.n26 VN.n25 27.0659
R755 VN.n6 VN.n5 27.0659
R756 VN.n8 VN.n3 24.4675
R757 VN.n11 VN.n9 24.4675
R758 VN.n28 VN.n23 24.4675
R759 VN.n30 VN.n29 24.4675
R760 VN.n10 VN.n1 20.0634
R761 VN.n22 VN.n20 20.0634
R762 VN.n17 VN.n16 13.2127
R763 VN.n36 VN.n35 13.2127
R764 VN.n4 VN.n3 4.40456
R765 VN.n11 VN.n10 4.40456
R766 VN.n24 VN.n23 4.40456
R767 VN.n30 VN.n22 4.40456
R768 VN.n37 VN.n19 0.189894
R769 VN.n33 VN.n19 0.189894
R770 VN.n33 VN.n32 0.189894
R771 VN.n32 VN.n31 0.189894
R772 VN.n31 VN.n21 0.189894
R773 VN.n27 VN.n21 0.189894
R774 VN.n27 VN.n26 0.189894
R775 VN.n7 VN.n6 0.189894
R776 VN.n7 VN.n2 0.189894
R777 VN.n12 VN.n2 0.189894
R778 VN.n13 VN.n12 0.189894
R779 VN.n14 VN.n13 0.189894
R780 VN.n14 VN.n0 0.189894
R781 VN.n18 VN.n0 0.189894
R782 VN VN.n18 0.0516364
R783 VTAIL.n194 VTAIL.n176 756.745
R784 VTAIL.n20 VTAIL.n2 756.745
R785 VTAIL.n44 VTAIL.n26 756.745
R786 VTAIL.n70 VTAIL.n52 756.745
R787 VTAIL.n170 VTAIL.n152 756.745
R788 VTAIL.n144 VTAIL.n126 756.745
R789 VTAIL.n120 VTAIL.n102 756.745
R790 VTAIL.n94 VTAIL.n76 756.745
R791 VTAIL.n185 VTAIL.n184 585
R792 VTAIL.n187 VTAIL.n186 585
R793 VTAIL.n180 VTAIL.n179 585
R794 VTAIL.n193 VTAIL.n192 585
R795 VTAIL.n195 VTAIL.n194 585
R796 VTAIL.n11 VTAIL.n10 585
R797 VTAIL.n13 VTAIL.n12 585
R798 VTAIL.n6 VTAIL.n5 585
R799 VTAIL.n19 VTAIL.n18 585
R800 VTAIL.n21 VTAIL.n20 585
R801 VTAIL.n35 VTAIL.n34 585
R802 VTAIL.n37 VTAIL.n36 585
R803 VTAIL.n30 VTAIL.n29 585
R804 VTAIL.n43 VTAIL.n42 585
R805 VTAIL.n45 VTAIL.n44 585
R806 VTAIL.n61 VTAIL.n60 585
R807 VTAIL.n63 VTAIL.n62 585
R808 VTAIL.n56 VTAIL.n55 585
R809 VTAIL.n69 VTAIL.n68 585
R810 VTAIL.n71 VTAIL.n70 585
R811 VTAIL.n171 VTAIL.n170 585
R812 VTAIL.n169 VTAIL.n168 585
R813 VTAIL.n156 VTAIL.n155 585
R814 VTAIL.n163 VTAIL.n162 585
R815 VTAIL.n161 VTAIL.n160 585
R816 VTAIL.n145 VTAIL.n144 585
R817 VTAIL.n143 VTAIL.n142 585
R818 VTAIL.n130 VTAIL.n129 585
R819 VTAIL.n137 VTAIL.n136 585
R820 VTAIL.n135 VTAIL.n134 585
R821 VTAIL.n121 VTAIL.n120 585
R822 VTAIL.n119 VTAIL.n118 585
R823 VTAIL.n106 VTAIL.n105 585
R824 VTAIL.n113 VTAIL.n112 585
R825 VTAIL.n111 VTAIL.n110 585
R826 VTAIL.n95 VTAIL.n94 585
R827 VTAIL.n93 VTAIL.n92 585
R828 VTAIL.n80 VTAIL.n79 585
R829 VTAIL.n87 VTAIL.n86 585
R830 VTAIL.n85 VTAIL.n84 585
R831 VTAIL.n183 VTAIL.t13 328.587
R832 VTAIL.n9 VTAIL.t15 328.587
R833 VTAIL.n33 VTAIL.t3 328.587
R834 VTAIL.n59 VTAIL.t0 328.587
R835 VTAIL.n159 VTAIL.t2 328.587
R836 VTAIL.n133 VTAIL.t6 328.587
R837 VTAIL.n109 VTAIL.t11 328.587
R838 VTAIL.n83 VTAIL.t10 328.587
R839 VTAIL.n186 VTAIL.n185 171.744
R840 VTAIL.n186 VTAIL.n179 171.744
R841 VTAIL.n193 VTAIL.n179 171.744
R842 VTAIL.n194 VTAIL.n193 171.744
R843 VTAIL.n12 VTAIL.n11 171.744
R844 VTAIL.n12 VTAIL.n5 171.744
R845 VTAIL.n19 VTAIL.n5 171.744
R846 VTAIL.n20 VTAIL.n19 171.744
R847 VTAIL.n36 VTAIL.n35 171.744
R848 VTAIL.n36 VTAIL.n29 171.744
R849 VTAIL.n43 VTAIL.n29 171.744
R850 VTAIL.n44 VTAIL.n43 171.744
R851 VTAIL.n62 VTAIL.n61 171.744
R852 VTAIL.n62 VTAIL.n55 171.744
R853 VTAIL.n69 VTAIL.n55 171.744
R854 VTAIL.n70 VTAIL.n69 171.744
R855 VTAIL.n170 VTAIL.n169 171.744
R856 VTAIL.n169 VTAIL.n155 171.744
R857 VTAIL.n162 VTAIL.n155 171.744
R858 VTAIL.n162 VTAIL.n161 171.744
R859 VTAIL.n144 VTAIL.n143 171.744
R860 VTAIL.n143 VTAIL.n129 171.744
R861 VTAIL.n136 VTAIL.n129 171.744
R862 VTAIL.n136 VTAIL.n135 171.744
R863 VTAIL.n120 VTAIL.n119 171.744
R864 VTAIL.n119 VTAIL.n105 171.744
R865 VTAIL.n112 VTAIL.n105 171.744
R866 VTAIL.n112 VTAIL.n111 171.744
R867 VTAIL.n94 VTAIL.n93 171.744
R868 VTAIL.n93 VTAIL.n79 171.744
R869 VTAIL.n86 VTAIL.n79 171.744
R870 VTAIL.n86 VTAIL.n85 171.744
R871 VTAIL.n151 VTAIL.n150 87.2071
R872 VTAIL.n101 VTAIL.n100 87.2071
R873 VTAIL.n1 VTAIL.n0 87.2069
R874 VTAIL.n51 VTAIL.n50 87.2069
R875 VTAIL.n185 VTAIL.t13 85.8723
R876 VTAIL.n11 VTAIL.t15 85.8723
R877 VTAIL.n35 VTAIL.t3 85.8723
R878 VTAIL.n61 VTAIL.t0 85.8723
R879 VTAIL.n161 VTAIL.t2 85.8723
R880 VTAIL.n135 VTAIL.t6 85.8723
R881 VTAIL.n111 VTAIL.t11 85.8723
R882 VTAIL.n85 VTAIL.t10 85.8723
R883 VTAIL.n199 VTAIL.n198 31.9914
R884 VTAIL.n25 VTAIL.n24 31.9914
R885 VTAIL.n49 VTAIL.n48 31.9914
R886 VTAIL.n75 VTAIL.n74 31.9914
R887 VTAIL.n175 VTAIL.n174 31.9914
R888 VTAIL.n149 VTAIL.n148 31.9914
R889 VTAIL.n125 VTAIL.n124 31.9914
R890 VTAIL.n99 VTAIL.n98 31.9914
R891 VTAIL.n199 VTAIL.n175 17.7376
R892 VTAIL.n99 VTAIL.n75 17.7376
R893 VTAIL.n184 VTAIL.n183 16.3651
R894 VTAIL.n10 VTAIL.n9 16.3651
R895 VTAIL.n34 VTAIL.n33 16.3651
R896 VTAIL.n60 VTAIL.n59 16.3651
R897 VTAIL.n160 VTAIL.n159 16.3651
R898 VTAIL.n134 VTAIL.n133 16.3651
R899 VTAIL.n110 VTAIL.n109 16.3651
R900 VTAIL.n84 VTAIL.n83 16.3651
R901 VTAIL.n187 VTAIL.n182 12.8005
R902 VTAIL.n13 VTAIL.n8 12.8005
R903 VTAIL.n37 VTAIL.n32 12.8005
R904 VTAIL.n63 VTAIL.n58 12.8005
R905 VTAIL.n163 VTAIL.n158 12.8005
R906 VTAIL.n137 VTAIL.n132 12.8005
R907 VTAIL.n113 VTAIL.n108 12.8005
R908 VTAIL.n87 VTAIL.n82 12.8005
R909 VTAIL.n188 VTAIL.n180 12.0247
R910 VTAIL.n14 VTAIL.n6 12.0247
R911 VTAIL.n38 VTAIL.n30 12.0247
R912 VTAIL.n64 VTAIL.n56 12.0247
R913 VTAIL.n164 VTAIL.n156 12.0247
R914 VTAIL.n138 VTAIL.n130 12.0247
R915 VTAIL.n114 VTAIL.n106 12.0247
R916 VTAIL.n88 VTAIL.n80 12.0247
R917 VTAIL.n192 VTAIL.n191 11.249
R918 VTAIL.n18 VTAIL.n17 11.249
R919 VTAIL.n42 VTAIL.n41 11.249
R920 VTAIL.n68 VTAIL.n67 11.249
R921 VTAIL.n168 VTAIL.n167 11.249
R922 VTAIL.n142 VTAIL.n141 11.249
R923 VTAIL.n118 VTAIL.n117 11.249
R924 VTAIL.n92 VTAIL.n91 11.249
R925 VTAIL.n195 VTAIL.n178 10.4732
R926 VTAIL.n21 VTAIL.n4 10.4732
R927 VTAIL.n45 VTAIL.n28 10.4732
R928 VTAIL.n71 VTAIL.n54 10.4732
R929 VTAIL.n171 VTAIL.n154 10.4732
R930 VTAIL.n145 VTAIL.n128 10.4732
R931 VTAIL.n121 VTAIL.n104 10.4732
R932 VTAIL.n95 VTAIL.n78 10.4732
R933 VTAIL.n196 VTAIL.n176 9.69747
R934 VTAIL.n22 VTAIL.n2 9.69747
R935 VTAIL.n46 VTAIL.n26 9.69747
R936 VTAIL.n72 VTAIL.n52 9.69747
R937 VTAIL.n172 VTAIL.n152 9.69747
R938 VTAIL.n146 VTAIL.n126 9.69747
R939 VTAIL.n122 VTAIL.n102 9.69747
R940 VTAIL.n96 VTAIL.n76 9.69747
R941 VTAIL.n198 VTAIL.n197 9.45567
R942 VTAIL.n24 VTAIL.n23 9.45567
R943 VTAIL.n48 VTAIL.n47 9.45567
R944 VTAIL.n74 VTAIL.n73 9.45567
R945 VTAIL.n174 VTAIL.n173 9.45567
R946 VTAIL.n148 VTAIL.n147 9.45567
R947 VTAIL.n124 VTAIL.n123 9.45567
R948 VTAIL.n98 VTAIL.n97 9.45567
R949 VTAIL.n197 VTAIL.n196 9.3005
R950 VTAIL.n178 VTAIL.n177 9.3005
R951 VTAIL.n191 VTAIL.n190 9.3005
R952 VTAIL.n189 VTAIL.n188 9.3005
R953 VTAIL.n182 VTAIL.n181 9.3005
R954 VTAIL.n23 VTAIL.n22 9.3005
R955 VTAIL.n4 VTAIL.n3 9.3005
R956 VTAIL.n17 VTAIL.n16 9.3005
R957 VTAIL.n15 VTAIL.n14 9.3005
R958 VTAIL.n8 VTAIL.n7 9.3005
R959 VTAIL.n47 VTAIL.n46 9.3005
R960 VTAIL.n28 VTAIL.n27 9.3005
R961 VTAIL.n41 VTAIL.n40 9.3005
R962 VTAIL.n39 VTAIL.n38 9.3005
R963 VTAIL.n32 VTAIL.n31 9.3005
R964 VTAIL.n73 VTAIL.n72 9.3005
R965 VTAIL.n54 VTAIL.n53 9.3005
R966 VTAIL.n67 VTAIL.n66 9.3005
R967 VTAIL.n65 VTAIL.n64 9.3005
R968 VTAIL.n58 VTAIL.n57 9.3005
R969 VTAIL.n173 VTAIL.n172 9.3005
R970 VTAIL.n154 VTAIL.n153 9.3005
R971 VTAIL.n167 VTAIL.n166 9.3005
R972 VTAIL.n165 VTAIL.n164 9.3005
R973 VTAIL.n158 VTAIL.n157 9.3005
R974 VTAIL.n147 VTAIL.n146 9.3005
R975 VTAIL.n128 VTAIL.n127 9.3005
R976 VTAIL.n141 VTAIL.n140 9.3005
R977 VTAIL.n139 VTAIL.n138 9.3005
R978 VTAIL.n132 VTAIL.n131 9.3005
R979 VTAIL.n123 VTAIL.n122 9.3005
R980 VTAIL.n104 VTAIL.n103 9.3005
R981 VTAIL.n117 VTAIL.n116 9.3005
R982 VTAIL.n115 VTAIL.n114 9.3005
R983 VTAIL.n108 VTAIL.n107 9.3005
R984 VTAIL.n97 VTAIL.n96 9.3005
R985 VTAIL.n78 VTAIL.n77 9.3005
R986 VTAIL.n91 VTAIL.n90 9.3005
R987 VTAIL.n89 VTAIL.n88 9.3005
R988 VTAIL.n82 VTAIL.n81 9.3005
R989 VTAIL.n0 VTAIL.t14 7.14446
R990 VTAIL.n0 VTAIL.t8 7.14446
R991 VTAIL.n50 VTAIL.t5 7.14446
R992 VTAIL.n50 VTAIL.t1 7.14446
R993 VTAIL.n150 VTAIL.t4 7.14446
R994 VTAIL.n150 VTAIL.t7 7.14446
R995 VTAIL.n100 VTAIL.t9 7.14446
R996 VTAIL.n100 VTAIL.t12 7.14446
R997 VTAIL.n198 VTAIL.n176 4.26717
R998 VTAIL.n24 VTAIL.n2 4.26717
R999 VTAIL.n48 VTAIL.n26 4.26717
R1000 VTAIL.n74 VTAIL.n52 4.26717
R1001 VTAIL.n174 VTAIL.n152 4.26717
R1002 VTAIL.n148 VTAIL.n126 4.26717
R1003 VTAIL.n124 VTAIL.n102 4.26717
R1004 VTAIL.n98 VTAIL.n76 4.26717
R1005 VTAIL.n183 VTAIL.n181 3.73474
R1006 VTAIL.n9 VTAIL.n7 3.73474
R1007 VTAIL.n33 VTAIL.n31 3.73474
R1008 VTAIL.n59 VTAIL.n57 3.73474
R1009 VTAIL.n159 VTAIL.n157 3.73474
R1010 VTAIL.n133 VTAIL.n131 3.73474
R1011 VTAIL.n109 VTAIL.n107 3.73474
R1012 VTAIL.n83 VTAIL.n81 3.73474
R1013 VTAIL.n196 VTAIL.n195 3.49141
R1014 VTAIL.n22 VTAIL.n21 3.49141
R1015 VTAIL.n46 VTAIL.n45 3.49141
R1016 VTAIL.n72 VTAIL.n71 3.49141
R1017 VTAIL.n172 VTAIL.n171 3.49141
R1018 VTAIL.n146 VTAIL.n145 3.49141
R1019 VTAIL.n122 VTAIL.n121 3.49141
R1020 VTAIL.n96 VTAIL.n95 3.49141
R1021 VTAIL.n192 VTAIL.n178 2.71565
R1022 VTAIL.n18 VTAIL.n4 2.71565
R1023 VTAIL.n42 VTAIL.n28 2.71565
R1024 VTAIL.n68 VTAIL.n54 2.71565
R1025 VTAIL.n168 VTAIL.n154 2.71565
R1026 VTAIL.n142 VTAIL.n128 2.71565
R1027 VTAIL.n118 VTAIL.n104 2.71565
R1028 VTAIL.n92 VTAIL.n78 2.71565
R1029 VTAIL.n191 VTAIL.n180 1.93989
R1030 VTAIL.n17 VTAIL.n6 1.93989
R1031 VTAIL.n41 VTAIL.n30 1.93989
R1032 VTAIL.n67 VTAIL.n56 1.93989
R1033 VTAIL.n167 VTAIL.n156 1.93989
R1034 VTAIL.n141 VTAIL.n130 1.93989
R1035 VTAIL.n117 VTAIL.n106 1.93989
R1036 VTAIL.n91 VTAIL.n80 1.93989
R1037 VTAIL.n101 VTAIL.n99 1.44878
R1038 VTAIL.n125 VTAIL.n101 1.44878
R1039 VTAIL.n151 VTAIL.n149 1.44878
R1040 VTAIL.n175 VTAIL.n151 1.44878
R1041 VTAIL.n75 VTAIL.n51 1.44878
R1042 VTAIL.n51 VTAIL.n49 1.44878
R1043 VTAIL.n25 VTAIL.n1 1.44878
R1044 VTAIL VTAIL.n199 1.39059
R1045 VTAIL.n188 VTAIL.n187 1.16414
R1046 VTAIL.n14 VTAIL.n13 1.16414
R1047 VTAIL.n38 VTAIL.n37 1.16414
R1048 VTAIL.n64 VTAIL.n63 1.16414
R1049 VTAIL.n164 VTAIL.n163 1.16414
R1050 VTAIL.n138 VTAIL.n137 1.16414
R1051 VTAIL.n114 VTAIL.n113 1.16414
R1052 VTAIL.n88 VTAIL.n87 1.16414
R1053 VTAIL.n149 VTAIL.n125 0.470328
R1054 VTAIL.n49 VTAIL.n25 0.470328
R1055 VTAIL.n184 VTAIL.n182 0.388379
R1056 VTAIL.n10 VTAIL.n8 0.388379
R1057 VTAIL.n34 VTAIL.n32 0.388379
R1058 VTAIL.n60 VTAIL.n58 0.388379
R1059 VTAIL.n160 VTAIL.n158 0.388379
R1060 VTAIL.n134 VTAIL.n132 0.388379
R1061 VTAIL.n110 VTAIL.n108 0.388379
R1062 VTAIL.n84 VTAIL.n82 0.388379
R1063 VTAIL.n189 VTAIL.n181 0.155672
R1064 VTAIL.n190 VTAIL.n189 0.155672
R1065 VTAIL.n190 VTAIL.n177 0.155672
R1066 VTAIL.n197 VTAIL.n177 0.155672
R1067 VTAIL.n15 VTAIL.n7 0.155672
R1068 VTAIL.n16 VTAIL.n15 0.155672
R1069 VTAIL.n16 VTAIL.n3 0.155672
R1070 VTAIL.n23 VTAIL.n3 0.155672
R1071 VTAIL.n39 VTAIL.n31 0.155672
R1072 VTAIL.n40 VTAIL.n39 0.155672
R1073 VTAIL.n40 VTAIL.n27 0.155672
R1074 VTAIL.n47 VTAIL.n27 0.155672
R1075 VTAIL.n65 VTAIL.n57 0.155672
R1076 VTAIL.n66 VTAIL.n65 0.155672
R1077 VTAIL.n66 VTAIL.n53 0.155672
R1078 VTAIL.n73 VTAIL.n53 0.155672
R1079 VTAIL.n173 VTAIL.n153 0.155672
R1080 VTAIL.n166 VTAIL.n153 0.155672
R1081 VTAIL.n166 VTAIL.n165 0.155672
R1082 VTAIL.n165 VTAIL.n157 0.155672
R1083 VTAIL.n147 VTAIL.n127 0.155672
R1084 VTAIL.n140 VTAIL.n127 0.155672
R1085 VTAIL.n140 VTAIL.n139 0.155672
R1086 VTAIL.n139 VTAIL.n131 0.155672
R1087 VTAIL.n123 VTAIL.n103 0.155672
R1088 VTAIL.n116 VTAIL.n103 0.155672
R1089 VTAIL.n116 VTAIL.n115 0.155672
R1090 VTAIL.n115 VTAIL.n107 0.155672
R1091 VTAIL.n97 VTAIL.n77 0.155672
R1092 VTAIL.n90 VTAIL.n77 0.155672
R1093 VTAIL.n90 VTAIL.n89 0.155672
R1094 VTAIL.n89 VTAIL.n81 0.155672
R1095 VTAIL VTAIL.n1 0.0586897
R1096 VDD2.n2 VDD2.n1 104.555
R1097 VDD2.n2 VDD2.n0 104.555
R1098 VDD2 VDD2.n5 104.552
R1099 VDD2.n4 VDD2.n3 103.885
R1100 VDD2.n4 VDD2.n2 34.1549
R1101 VDD2.n5 VDD2.t1 7.14446
R1102 VDD2.n5 VDD2.t6 7.14446
R1103 VDD2.n3 VDD2.t0 7.14446
R1104 VDD2.n3 VDD2.t5 7.14446
R1105 VDD2.n1 VDD2.t3 7.14446
R1106 VDD2.n1 VDD2.t7 7.14446
R1107 VDD2.n0 VDD2.t4 7.14446
R1108 VDD2.n0 VDD2.t2 7.14446
R1109 VDD2 VDD2.n4 0.782828
R1110 VP.n25 VP.n5 172.555
R1111 VP.n44 VP.n43 172.555
R1112 VP.n24 VP.n23 172.555
R1113 VP.n12 VP.n9 161.3
R1114 VP.n14 VP.n13 161.3
R1115 VP.n15 VP.n8 161.3
R1116 VP.n18 VP.n17 161.3
R1117 VP.n19 VP.n7 161.3
R1118 VP.n21 VP.n20 161.3
R1119 VP.n22 VP.n6 161.3
R1120 VP.n42 VP.n0 161.3
R1121 VP.n41 VP.n40 161.3
R1122 VP.n39 VP.n1 161.3
R1123 VP.n38 VP.n37 161.3
R1124 VP.n35 VP.n2 161.3
R1125 VP.n34 VP.n33 161.3
R1126 VP.n32 VP.n3 161.3
R1127 VP.n31 VP.n30 161.3
R1128 VP.n28 VP.n4 161.3
R1129 VP.n27 VP.n26 161.3
R1130 VP.n11 VP.t0 110.861
R1131 VP.n5 VP.t7 81.2264
R1132 VP.n29 VP.t1 81.2264
R1133 VP.n36 VP.t6 81.2264
R1134 VP.n43 VP.t4 81.2264
R1135 VP.n23 VP.t2 81.2264
R1136 VP.n16 VP.t5 81.2264
R1137 VP.n10 VP.t3 81.2264
R1138 VP.n11 VP.n10 60.7907
R1139 VP.n35 VP.n34 56.5193
R1140 VP.n15 VP.n14 56.5193
R1141 VP.n30 VP.n28 47.2923
R1142 VP.n41 VP.n1 47.2923
R1143 VP.n21 VP.n7 47.2923
R1144 VP.n25 VP.n24 39.3414
R1145 VP.n28 VP.n27 33.6945
R1146 VP.n42 VP.n41 33.6945
R1147 VP.n22 VP.n21 33.6945
R1148 VP.n12 VP.n11 27.0659
R1149 VP.n34 VP.n3 24.4675
R1150 VP.n37 VP.n35 24.4675
R1151 VP.n17 VP.n15 24.4675
R1152 VP.n14 VP.n9 24.4675
R1153 VP.n30 VP.n29 20.0634
R1154 VP.n36 VP.n1 20.0634
R1155 VP.n16 VP.n7 20.0634
R1156 VP.n27 VP.n5 13.2127
R1157 VP.n43 VP.n42 13.2127
R1158 VP.n23 VP.n22 13.2127
R1159 VP.n29 VP.n3 4.40456
R1160 VP.n37 VP.n36 4.40456
R1161 VP.n17 VP.n16 4.40456
R1162 VP.n10 VP.n9 4.40456
R1163 VP.n13 VP.n12 0.189894
R1164 VP.n13 VP.n8 0.189894
R1165 VP.n18 VP.n8 0.189894
R1166 VP.n19 VP.n18 0.189894
R1167 VP.n20 VP.n19 0.189894
R1168 VP.n20 VP.n6 0.189894
R1169 VP.n24 VP.n6 0.189894
R1170 VP.n26 VP.n25 0.189894
R1171 VP.n26 VP.n4 0.189894
R1172 VP.n31 VP.n4 0.189894
R1173 VP.n32 VP.n31 0.189894
R1174 VP.n33 VP.n32 0.189894
R1175 VP.n33 VP.n2 0.189894
R1176 VP.n38 VP.n2 0.189894
R1177 VP.n39 VP.n38 0.189894
R1178 VP.n40 VP.n39 0.189894
R1179 VP.n40 VP.n0 0.189894
R1180 VP.n44 VP.n0 0.189894
R1181 VP VP.n44 0.0516364
R1182 VDD1 VDD1.n0 104.668
R1183 VDD1.n3 VDD1.n2 104.555
R1184 VDD1.n3 VDD1.n1 104.555
R1185 VDD1.n5 VDD1.n4 103.885
R1186 VDD1.n5 VDD1.n3 34.738
R1187 VDD1.n4 VDD1.t2 7.14446
R1188 VDD1.n4 VDD1.t5 7.14446
R1189 VDD1.n0 VDD1.t7 7.14446
R1190 VDD1.n0 VDD1.t4 7.14446
R1191 VDD1.n2 VDD1.t1 7.14446
R1192 VDD1.n2 VDD1.t3 7.14446
R1193 VDD1.n1 VDD1.t0 7.14446
R1194 VDD1.n1 VDD1.t6 7.14446
R1195 VDD1 VDD1.n5 0.666448
C0 w_n2650_n1878# VP 5.24626f
C1 w_n2650_n1878# B 6.11756f
C2 B VP 1.42385f
C3 VN VTAIL 3.43048f
C4 VN VDD1 0.153184f
C5 VDD2 VN 3.03316f
C6 w_n2650_n1878# VN 4.9061f
C7 VDD1 VTAIL 5.01186f
C8 VP VN 4.75937f
C9 B VN 0.860088f
C10 VDD2 VTAIL 5.05789f
C11 VDD2 VDD1 1.15064f
C12 w_n2650_n1878# VTAIL 2.37382f
C13 w_n2650_n1878# VDD1 1.33431f
C14 VP VTAIL 3.44459f
C15 VP VDD1 3.26954f
C16 B VTAIL 2.08724f
C17 B VDD1 1.06781f
C18 w_n2650_n1878# VDD2 1.3962f
C19 VDD2 VP 0.39076f
C20 VDD2 B 1.1247f
C21 VDD2 VSUBS 1.169622f
C22 VDD1 VSUBS 1.597455f
C23 VTAIL VSUBS 0.534176f
C24 VN VSUBS 4.81913f
C25 VP VSUBS 1.856105f
C26 B VSUBS 2.829213f
C27 w_n2650_n1878# VSUBS 62.487003f
C28 VDD1.t7 VSUBS 0.090899f
C29 VDD1.t4 VSUBS 0.090899f
C30 VDD1.n0 VSUBS 0.558452f
C31 VDD1.t0 VSUBS 0.090899f
C32 VDD1.t6 VSUBS 0.090899f
C33 VDD1.n1 VSUBS 0.557785f
C34 VDD1.t1 VSUBS 0.090899f
C35 VDD1.t3 VSUBS 0.090899f
C36 VDD1.n2 VSUBS 0.557785f
C37 VDD1.n3 VSUBS 2.51505f
C38 VDD1.t2 VSUBS 0.090899f
C39 VDD1.t5 VSUBS 0.090899f
C40 VDD1.n4 VSUBS 0.554212f
C41 VDD1.n5 VSUBS 2.14885f
C42 VP.n0 VSUBS 0.053266f
C43 VP.t4 VSUBS 0.849762f
C44 VP.n1 VSUBS 0.091868f
C45 VP.n2 VSUBS 0.053266f
C46 VP.n3 VSUBS 0.059085f
C47 VP.n4 VSUBS 0.053266f
C48 VP.t7 VSUBS 0.849762f
C49 VP.n5 VSUBS 0.458454f
C50 VP.n6 VSUBS 0.053266f
C51 VP.t2 VSUBS 0.849762f
C52 VP.n7 VSUBS 0.091868f
C53 VP.n8 VSUBS 0.053266f
C54 VP.n9 VSUBS 0.059085f
C55 VP.t0 VSUBS 0.991674f
C56 VP.t3 VSUBS 0.849762f
C57 VP.n10 VSUBS 0.429206f
C58 VP.n11 VSUBS 0.468156f
C59 VP.n12 VSUBS 0.283646f
C60 VP.n13 VSUBS 0.053266f
C61 VP.n14 VSUBS 0.077759f
C62 VP.n15 VSUBS 0.077759f
C63 VP.t5 VSUBS 0.849762f
C64 VP.n16 VSUBS 0.354658f
C65 VP.n17 VSUBS 0.059085f
C66 VP.n18 VSUBS 0.053266f
C67 VP.n19 VSUBS 0.053266f
C68 VP.n20 VSUBS 0.053266f
C69 VP.n21 VSUBS 0.04651f
C70 VP.n22 VSUBS 0.085047f
C71 VP.n23 VSUBS 0.458454f
C72 VP.n24 VSUBS 1.97387f
C73 VP.n25 VSUBS 2.02254f
C74 VP.n26 VSUBS 0.053266f
C75 VP.n27 VSUBS 0.085047f
C76 VP.n28 VSUBS 0.04651f
C77 VP.t1 VSUBS 0.849762f
C78 VP.n29 VSUBS 0.354658f
C79 VP.n30 VSUBS 0.091868f
C80 VP.n31 VSUBS 0.053266f
C81 VP.n32 VSUBS 0.053266f
C82 VP.n33 VSUBS 0.053266f
C83 VP.n34 VSUBS 0.077759f
C84 VP.n35 VSUBS 0.077759f
C85 VP.t6 VSUBS 0.849762f
C86 VP.n36 VSUBS 0.354658f
C87 VP.n37 VSUBS 0.059085f
C88 VP.n38 VSUBS 0.053266f
C89 VP.n39 VSUBS 0.053266f
C90 VP.n40 VSUBS 0.053266f
C91 VP.n41 VSUBS 0.04651f
C92 VP.n42 VSUBS 0.085047f
C93 VP.n43 VSUBS 0.458454f
C94 VP.n44 VSUBS 0.048522f
C95 VDD2.t4 VSUBS 0.089718f
C96 VDD2.t2 VSUBS 0.089718f
C97 VDD2.n0 VSUBS 0.550538f
C98 VDD2.t3 VSUBS 0.089718f
C99 VDD2.t7 VSUBS 0.089718f
C100 VDD2.n1 VSUBS 0.550538f
C101 VDD2.n2 VSUBS 2.42938f
C102 VDD2.t0 VSUBS 0.089718f
C103 VDD2.t5 VSUBS 0.089718f
C104 VDD2.n3 VSUBS 0.547014f
C105 VDD2.n4 VSUBS 2.09112f
C106 VDD2.t1 VSUBS 0.089718f
C107 VDD2.t6 VSUBS 0.089718f
C108 VDD2.n5 VSUBS 0.550516f
C109 VTAIL.t14 VSUBS 0.104507f
C110 VTAIL.t8 VSUBS 0.104507f
C111 VTAIL.n0 VSUBS 0.55577f
C112 VTAIL.n1 VSUBS 0.614174f
C113 VTAIL.n2 VSUBS 0.030707f
C114 VTAIL.n3 VSUBS 0.029066f
C115 VTAIL.n4 VSUBS 0.015619f
C116 VTAIL.n5 VSUBS 0.036917f
C117 VTAIL.n6 VSUBS 0.016537f
C118 VTAIL.n7 VSUBS 0.47378f
C119 VTAIL.n8 VSUBS 0.015619f
C120 VTAIL.t15 VSUBS 0.080118f
C121 VTAIL.n9 VSUBS 0.116798f
C122 VTAIL.n10 VSUBS 0.023387f
C123 VTAIL.n11 VSUBS 0.027688f
C124 VTAIL.n12 VSUBS 0.036917f
C125 VTAIL.n13 VSUBS 0.016537f
C126 VTAIL.n14 VSUBS 0.015619f
C127 VTAIL.n15 VSUBS 0.029066f
C128 VTAIL.n16 VSUBS 0.029066f
C129 VTAIL.n17 VSUBS 0.015619f
C130 VTAIL.n18 VSUBS 0.016537f
C131 VTAIL.n19 VSUBS 0.036917f
C132 VTAIL.n20 VSUBS 0.08518f
C133 VTAIL.n21 VSUBS 0.016537f
C134 VTAIL.n22 VSUBS 0.015619f
C135 VTAIL.n23 VSUBS 0.066787f
C136 VTAIL.n24 VSUBS 0.042638f
C137 VTAIL.n25 VSUBS 0.204242f
C138 VTAIL.n26 VSUBS 0.030707f
C139 VTAIL.n27 VSUBS 0.029066f
C140 VTAIL.n28 VSUBS 0.015619f
C141 VTAIL.n29 VSUBS 0.036917f
C142 VTAIL.n30 VSUBS 0.016537f
C143 VTAIL.n31 VSUBS 0.47378f
C144 VTAIL.n32 VSUBS 0.015619f
C145 VTAIL.t3 VSUBS 0.080118f
C146 VTAIL.n33 VSUBS 0.116798f
C147 VTAIL.n34 VSUBS 0.023387f
C148 VTAIL.n35 VSUBS 0.027688f
C149 VTAIL.n36 VSUBS 0.036917f
C150 VTAIL.n37 VSUBS 0.016537f
C151 VTAIL.n38 VSUBS 0.015619f
C152 VTAIL.n39 VSUBS 0.029066f
C153 VTAIL.n40 VSUBS 0.029066f
C154 VTAIL.n41 VSUBS 0.015619f
C155 VTAIL.n42 VSUBS 0.016537f
C156 VTAIL.n43 VSUBS 0.036917f
C157 VTAIL.n44 VSUBS 0.08518f
C158 VTAIL.n45 VSUBS 0.016537f
C159 VTAIL.n46 VSUBS 0.015619f
C160 VTAIL.n47 VSUBS 0.066787f
C161 VTAIL.n48 VSUBS 0.042638f
C162 VTAIL.n49 VSUBS 0.204242f
C163 VTAIL.t5 VSUBS 0.104507f
C164 VTAIL.t1 VSUBS 0.104507f
C165 VTAIL.n50 VSUBS 0.55577f
C166 VTAIL.n51 VSUBS 0.744364f
C167 VTAIL.n52 VSUBS 0.030707f
C168 VTAIL.n53 VSUBS 0.029066f
C169 VTAIL.n54 VSUBS 0.015619f
C170 VTAIL.n55 VSUBS 0.036917f
C171 VTAIL.n56 VSUBS 0.016537f
C172 VTAIL.n57 VSUBS 0.47378f
C173 VTAIL.n58 VSUBS 0.015619f
C174 VTAIL.t0 VSUBS 0.080118f
C175 VTAIL.n59 VSUBS 0.116798f
C176 VTAIL.n60 VSUBS 0.023387f
C177 VTAIL.n61 VSUBS 0.027688f
C178 VTAIL.n62 VSUBS 0.036917f
C179 VTAIL.n63 VSUBS 0.016537f
C180 VTAIL.n64 VSUBS 0.015619f
C181 VTAIL.n65 VSUBS 0.029066f
C182 VTAIL.n66 VSUBS 0.029066f
C183 VTAIL.n67 VSUBS 0.015619f
C184 VTAIL.n68 VSUBS 0.016537f
C185 VTAIL.n69 VSUBS 0.036917f
C186 VTAIL.n70 VSUBS 0.08518f
C187 VTAIL.n71 VSUBS 0.016537f
C188 VTAIL.n72 VSUBS 0.015619f
C189 VTAIL.n73 VSUBS 0.066787f
C190 VTAIL.n74 VSUBS 0.042638f
C191 VTAIL.n75 VSUBS 1.05806f
C192 VTAIL.n76 VSUBS 0.030707f
C193 VTAIL.n77 VSUBS 0.029066f
C194 VTAIL.n78 VSUBS 0.015619f
C195 VTAIL.n79 VSUBS 0.036917f
C196 VTAIL.n80 VSUBS 0.016537f
C197 VTAIL.n81 VSUBS 0.473779f
C198 VTAIL.n82 VSUBS 0.015619f
C199 VTAIL.t10 VSUBS 0.080118f
C200 VTAIL.n83 VSUBS 0.116798f
C201 VTAIL.n84 VSUBS 0.023387f
C202 VTAIL.n85 VSUBS 0.027688f
C203 VTAIL.n86 VSUBS 0.036917f
C204 VTAIL.n87 VSUBS 0.016537f
C205 VTAIL.n88 VSUBS 0.015619f
C206 VTAIL.n89 VSUBS 0.029066f
C207 VTAIL.n90 VSUBS 0.029066f
C208 VTAIL.n91 VSUBS 0.015619f
C209 VTAIL.n92 VSUBS 0.016537f
C210 VTAIL.n93 VSUBS 0.036917f
C211 VTAIL.n94 VSUBS 0.08518f
C212 VTAIL.n95 VSUBS 0.016537f
C213 VTAIL.n96 VSUBS 0.015619f
C214 VTAIL.n97 VSUBS 0.066787f
C215 VTAIL.n98 VSUBS 0.042638f
C216 VTAIL.n99 VSUBS 1.05806f
C217 VTAIL.t9 VSUBS 0.104507f
C218 VTAIL.t12 VSUBS 0.104507f
C219 VTAIL.n100 VSUBS 0.555774f
C220 VTAIL.n101 VSUBS 0.74436f
C221 VTAIL.n102 VSUBS 0.030707f
C222 VTAIL.n103 VSUBS 0.029066f
C223 VTAIL.n104 VSUBS 0.015619f
C224 VTAIL.n105 VSUBS 0.036917f
C225 VTAIL.n106 VSUBS 0.016537f
C226 VTAIL.n107 VSUBS 0.473779f
C227 VTAIL.n108 VSUBS 0.015619f
C228 VTAIL.t11 VSUBS 0.080118f
C229 VTAIL.n109 VSUBS 0.116798f
C230 VTAIL.n110 VSUBS 0.023387f
C231 VTAIL.n111 VSUBS 0.027688f
C232 VTAIL.n112 VSUBS 0.036917f
C233 VTAIL.n113 VSUBS 0.016537f
C234 VTAIL.n114 VSUBS 0.015619f
C235 VTAIL.n115 VSUBS 0.029066f
C236 VTAIL.n116 VSUBS 0.029066f
C237 VTAIL.n117 VSUBS 0.015619f
C238 VTAIL.n118 VSUBS 0.016537f
C239 VTAIL.n119 VSUBS 0.036917f
C240 VTAIL.n120 VSUBS 0.08518f
C241 VTAIL.n121 VSUBS 0.016537f
C242 VTAIL.n122 VSUBS 0.015619f
C243 VTAIL.n123 VSUBS 0.066787f
C244 VTAIL.n124 VSUBS 0.042638f
C245 VTAIL.n125 VSUBS 0.204242f
C246 VTAIL.n126 VSUBS 0.030707f
C247 VTAIL.n127 VSUBS 0.029066f
C248 VTAIL.n128 VSUBS 0.015619f
C249 VTAIL.n129 VSUBS 0.036917f
C250 VTAIL.n130 VSUBS 0.016537f
C251 VTAIL.n131 VSUBS 0.473779f
C252 VTAIL.n132 VSUBS 0.015619f
C253 VTAIL.t6 VSUBS 0.080118f
C254 VTAIL.n133 VSUBS 0.116798f
C255 VTAIL.n134 VSUBS 0.023387f
C256 VTAIL.n135 VSUBS 0.027688f
C257 VTAIL.n136 VSUBS 0.036917f
C258 VTAIL.n137 VSUBS 0.016537f
C259 VTAIL.n138 VSUBS 0.015619f
C260 VTAIL.n139 VSUBS 0.029066f
C261 VTAIL.n140 VSUBS 0.029066f
C262 VTAIL.n141 VSUBS 0.015619f
C263 VTAIL.n142 VSUBS 0.016537f
C264 VTAIL.n143 VSUBS 0.036917f
C265 VTAIL.n144 VSUBS 0.08518f
C266 VTAIL.n145 VSUBS 0.016537f
C267 VTAIL.n146 VSUBS 0.015619f
C268 VTAIL.n147 VSUBS 0.066787f
C269 VTAIL.n148 VSUBS 0.042638f
C270 VTAIL.n149 VSUBS 0.204242f
C271 VTAIL.t4 VSUBS 0.104507f
C272 VTAIL.t7 VSUBS 0.104507f
C273 VTAIL.n150 VSUBS 0.555774f
C274 VTAIL.n151 VSUBS 0.74436f
C275 VTAIL.n152 VSUBS 0.030707f
C276 VTAIL.n153 VSUBS 0.029066f
C277 VTAIL.n154 VSUBS 0.015619f
C278 VTAIL.n155 VSUBS 0.036917f
C279 VTAIL.n156 VSUBS 0.016537f
C280 VTAIL.n157 VSUBS 0.473779f
C281 VTAIL.n158 VSUBS 0.015619f
C282 VTAIL.t2 VSUBS 0.080118f
C283 VTAIL.n159 VSUBS 0.116798f
C284 VTAIL.n160 VSUBS 0.023387f
C285 VTAIL.n161 VSUBS 0.027688f
C286 VTAIL.n162 VSUBS 0.036917f
C287 VTAIL.n163 VSUBS 0.016537f
C288 VTAIL.n164 VSUBS 0.015619f
C289 VTAIL.n165 VSUBS 0.029066f
C290 VTAIL.n166 VSUBS 0.029066f
C291 VTAIL.n167 VSUBS 0.015619f
C292 VTAIL.n168 VSUBS 0.016537f
C293 VTAIL.n169 VSUBS 0.036917f
C294 VTAIL.n170 VSUBS 0.08518f
C295 VTAIL.n171 VSUBS 0.016537f
C296 VTAIL.n172 VSUBS 0.015619f
C297 VTAIL.n173 VSUBS 0.066787f
C298 VTAIL.n174 VSUBS 0.042638f
C299 VTAIL.n175 VSUBS 1.05806f
C300 VTAIL.n176 VSUBS 0.030707f
C301 VTAIL.n177 VSUBS 0.029066f
C302 VTAIL.n178 VSUBS 0.015619f
C303 VTAIL.n179 VSUBS 0.036917f
C304 VTAIL.n180 VSUBS 0.016537f
C305 VTAIL.n181 VSUBS 0.47378f
C306 VTAIL.n182 VSUBS 0.015619f
C307 VTAIL.t13 VSUBS 0.080118f
C308 VTAIL.n183 VSUBS 0.116798f
C309 VTAIL.n184 VSUBS 0.023387f
C310 VTAIL.n185 VSUBS 0.027688f
C311 VTAIL.n186 VSUBS 0.036917f
C312 VTAIL.n187 VSUBS 0.016537f
C313 VTAIL.n188 VSUBS 0.015619f
C314 VTAIL.n189 VSUBS 0.029066f
C315 VTAIL.n190 VSUBS 0.029066f
C316 VTAIL.n191 VSUBS 0.015619f
C317 VTAIL.n192 VSUBS 0.016537f
C318 VTAIL.n193 VSUBS 0.036917f
C319 VTAIL.n194 VSUBS 0.08518f
C320 VTAIL.n195 VSUBS 0.016537f
C321 VTAIL.n196 VSUBS 0.015619f
C322 VTAIL.n197 VSUBS 0.066787f
C323 VTAIL.n198 VSUBS 0.042638f
C324 VTAIL.n199 VSUBS 1.05261f
C325 VN.n0 VSUBS 0.051123f
C326 VN.t0 VSUBS 0.815574f
C327 VN.n1 VSUBS 0.088172f
C328 VN.n2 VSUBS 0.051123f
C329 VN.n3 VSUBS 0.056708f
C330 VN.t3 VSUBS 0.951778f
C331 VN.t5 VSUBS 0.815574f
C332 VN.n4 VSUBS 0.411938f
C333 VN.n5 VSUBS 0.449321f
C334 VN.n6 VSUBS 0.272234f
C335 VN.n7 VSUBS 0.051123f
C336 VN.n8 VSUBS 0.074631f
C337 VN.n9 VSUBS 0.074631f
C338 VN.t4 VSUBS 0.815574f
C339 VN.n10 VSUBS 0.34039f
C340 VN.n11 VSUBS 0.056708f
C341 VN.n12 VSUBS 0.051123f
C342 VN.n13 VSUBS 0.051123f
C343 VN.n14 VSUBS 0.051123f
C344 VN.n15 VSUBS 0.044639f
C345 VN.n16 VSUBS 0.081626f
C346 VN.n17 VSUBS 0.44001f
C347 VN.n18 VSUBS 0.04657f
C348 VN.n19 VSUBS 0.051123f
C349 VN.t7 VSUBS 0.815574f
C350 VN.n20 VSUBS 0.088172f
C351 VN.n21 VSUBS 0.051123f
C352 VN.t2 VSUBS 0.815574f
C353 VN.n22 VSUBS 0.34039f
C354 VN.n23 VSUBS 0.056708f
C355 VN.t1 VSUBS 0.951778f
C356 VN.t6 VSUBS 0.815574f
C357 VN.n24 VSUBS 0.411938f
C358 VN.n25 VSUBS 0.449321f
C359 VN.n26 VSUBS 0.272234f
C360 VN.n27 VSUBS 0.051123f
C361 VN.n28 VSUBS 0.074631f
C362 VN.n29 VSUBS 0.074631f
C363 VN.n30 VSUBS 0.056708f
C364 VN.n31 VSUBS 0.051123f
C365 VN.n32 VSUBS 0.051123f
C366 VN.n33 VSUBS 0.051123f
C367 VN.n34 VSUBS 0.044639f
C368 VN.n35 VSUBS 0.081626f
C369 VN.n36 VSUBS 0.44001f
C370 VN.n37 VSUBS 1.92816f
C371 B.n0 VSUBS 0.005828f
C372 B.n1 VSUBS 0.005828f
C373 B.n2 VSUBS 0.009217f
C374 B.n3 VSUBS 0.009217f
C375 B.n4 VSUBS 0.009217f
C376 B.n5 VSUBS 0.009217f
C377 B.n6 VSUBS 0.009217f
C378 B.n7 VSUBS 0.009217f
C379 B.n8 VSUBS 0.009217f
C380 B.n9 VSUBS 0.009217f
C381 B.n10 VSUBS 0.009217f
C382 B.n11 VSUBS 0.009217f
C383 B.n12 VSUBS 0.009217f
C384 B.n13 VSUBS 0.009217f
C385 B.n14 VSUBS 0.009217f
C386 B.n15 VSUBS 0.009217f
C387 B.n16 VSUBS 0.009217f
C388 B.n17 VSUBS 0.009217f
C389 B.n18 VSUBS 0.020217f
C390 B.n19 VSUBS 0.009217f
C391 B.n20 VSUBS 0.009217f
C392 B.n21 VSUBS 0.009217f
C393 B.n22 VSUBS 0.009217f
C394 B.n23 VSUBS 0.009217f
C395 B.n24 VSUBS 0.009217f
C396 B.n25 VSUBS 0.009217f
C397 B.n26 VSUBS 0.009217f
C398 B.n27 VSUBS 0.009217f
C399 B.n28 VSUBS 0.00637f
C400 B.n29 VSUBS 0.009217f
C401 B.t2 VSUBS 0.086428f
C402 B.t1 VSUBS 0.103948f
C403 B.t0 VSUBS 0.374546f
C404 B.n30 VSUBS 0.187978f
C405 B.n31 VSUBS 0.161537f
C406 B.n32 VSUBS 0.021354f
C407 B.n33 VSUBS 0.009217f
C408 B.n34 VSUBS 0.009217f
C409 B.n35 VSUBS 0.009217f
C410 B.n36 VSUBS 0.009217f
C411 B.t11 VSUBS 0.086429f
C412 B.t10 VSUBS 0.10395f
C413 B.t9 VSUBS 0.374546f
C414 B.n37 VSUBS 0.187977f
C415 B.n38 VSUBS 0.161535f
C416 B.n39 VSUBS 0.009217f
C417 B.n40 VSUBS 0.009217f
C418 B.n41 VSUBS 0.009217f
C419 B.n42 VSUBS 0.009217f
C420 B.n43 VSUBS 0.009217f
C421 B.n44 VSUBS 0.009217f
C422 B.n45 VSUBS 0.009217f
C423 B.n46 VSUBS 0.009217f
C424 B.n47 VSUBS 0.009217f
C425 B.n48 VSUBS 0.020217f
C426 B.n49 VSUBS 0.009217f
C427 B.n50 VSUBS 0.009217f
C428 B.n51 VSUBS 0.009217f
C429 B.n52 VSUBS 0.009217f
C430 B.n53 VSUBS 0.009217f
C431 B.n54 VSUBS 0.009217f
C432 B.n55 VSUBS 0.009217f
C433 B.n56 VSUBS 0.009217f
C434 B.n57 VSUBS 0.009217f
C435 B.n58 VSUBS 0.009217f
C436 B.n59 VSUBS 0.009217f
C437 B.n60 VSUBS 0.009217f
C438 B.n61 VSUBS 0.009217f
C439 B.n62 VSUBS 0.009217f
C440 B.n63 VSUBS 0.009217f
C441 B.n64 VSUBS 0.009217f
C442 B.n65 VSUBS 0.009217f
C443 B.n66 VSUBS 0.009217f
C444 B.n67 VSUBS 0.009217f
C445 B.n68 VSUBS 0.009217f
C446 B.n69 VSUBS 0.009217f
C447 B.n70 VSUBS 0.009217f
C448 B.n71 VSUBS 0.009217f
C449 B.n72 VSUBS 0.009217f
C450 B.n73 VSUBS 0.009217f
C451 B.n74 VSUBS 0.009217f
C452 B.n75 VSUBS 0.009217f
C453 B.n76 VSUBS 0.009217f
C454 B.n77 VSUBS 0.009217f
C455 B.n78 VSUBS 0.009217f
C456 B.n79 VSUBS 0.009217f
C457 B.n80 VSUBS 0.009217f
C458 B.n81 VSUBS 0.020217f
C459 B.n82 VSUBS 0.009217f
C460 B.n83 VSUBS 0.009217f
C461 B.n84 VSUBS 0.009217f
C462 B.n85 VSUBS 0.009217f
C463 B.n86 VSUBS 0.009217f
C464 B.n87 VSUBS 0.009217f
C465 B.n88 VSUBS 0.009217f
C466 B.n89 VSUBS 0.009217f
C467 B.n90 VSUBS 0.009217f
C468 B.n91 VSUBS 0.00637f
C469 B.n92 VSUBS 0.009217f
C470 B.n93 VSUBS 0.009217f
C471 B.n94 VSUBS 0.009217f
C472 B.n95 VSUBS 0.009217f
C473 B.n96 VSUBS 0.009217f
C474 B.t7 VSUBS 0.086428f
C475 B.t8 VSUBS 0.103948f
C476 B.t6 VSUBS 0.374546f
C477 B.n97 VSUBS 0.187978f
C478 B.n98 VSUBS 0.161537f
C479 B.n99 VSUBS 0.009217f
C480 B.n100 VSUBS 0.009217f
C481 B.n101 VSUBS 0.009217f
C482 B.n102 VSUBS 0.009217f
C483 B.n103 VSUBS 0.009217f
C484 B.n104 VSUBS 0.009217f
C485 B.n105 VSUBS 0.009217f
C486 B.n106 VSUBS 0.009217f
C487 B.n107 VSUBS 0.009217f
C488 B.n108 VSUBS 0.020217f
C489 B.n109 VSUBS 0.009217f
C490 B.n110 VSUBS 0.009217f
C491 B.n111 VSUBS 0.009217f
C492 B.n112 VSUBS 0.009217f
C493 B.n113 VSUBS 0.009217f
C494 B.n114 VSUBS 0.009217f
C495 B.n115 VSUBS 0.009217f
C496 B.n116 VSUBS 0.009217f
C497 B.n117 VSUBS 0.009217f
C498 B.n118 VSUBS 0.009217f
C499 B.n119 VSUBS 0.009217f
C500 B.n120 VSUBS 0.009217f
C501 B.n121 VSUBS 0.009217f
C502 B.n122 VSUBS 0.009217f
C503 B.n123 VSUBS 0.009217f
C504 B.n124 VSUBS 0.009217f
C505 B.n125 VSUBS 0.009217f
C506 B.n126 VSUBS 0.009217f
C507 B.n127 VSUBS 0.009217f
C508 B.n128 VSUBS 0.009217f
C509 B.n129 VSUBS 0.009217f
C510 B.n130 VSUBS 0.009217f
C511 B.n131 VSUBS 0.009217f
C512 B.n132 VSUBS 0.009217f
C513 B.n133 VSUBS 0.009217f
C514 B.n134 VSUBS 0.009217f
C515 B.n135 VSUBS 0.009217f
C516 B.n136 VSUBS 0.009217f
C517 B.n137 VSUBS 0.009217f
C518 B.n138 VSUBS 0.009217f
C519 B.n139 VSUBS 0.009217f
C520 B.n140 VSUBS 0.009217f
C521 B.n141 VSUBS 0.009217f
C522 B.n142 VSUBS 0.009217f
C523 B.n143 VSUBS 0.009217f
C524 B.n144 VSUBS 0.009217f
C525 B.n145 VSUBS 0.009217f
C526 B.n146 VSUBS 0.009217f
C527 B.n147 VSUBS 0.009217f
C528 B.n148 VSUBS 0.009217f
C529 B.n149 VSUBS 0.009217f
C530 B.n150 VSUBS 0.009217f
C531 B.n151 VSUBS 0.009217f
C532 B.n152 VSUBS 0.009217f
C533 B.n153 VSUBS 0.009217f
C534 B.n154 VSUBS 0.009217f
C535 B.n155 VSUBS 0.009217f
C536 B.n156 VSUBS 0.009217f
C537 B.n157 VSUBS 0.009217f
C538 B.n158 VSUBS 0.009217f
C539 B.n159 VSUBS 0.009217f
C540 B.n160 VSUBS 0.009217f
C541 B.n161 VSUBS 0.009217f
C542 B.n162 VSUBS 0.009217f
C543 B.n163 VSUBS 0.009217f
C544 B.n164 VSUBS 0.009217f
C545 B.n165 VSUBS 0.009217f
C546 B.n166 VSUBS 0.009217f
C547 B.n167 VSUBS 0.009217f
C548 B.n168 VSUBS 0.009217f
C549 B.n169 VSUBS 0.009217f
C550 B.n170 VSUBS 0.009217f
C551 B.n171 VSUBS 0.020217f
C552 B.n172 VSUBS 0.020987f
C553 B.n173 VSUBS 0.020987f
C554 B.n174 VSUBS 0.009217f
C555 B.n175 VSUBS 0.009217f
C556 B.n176 VSUBS 0.009217f
C557 B.n177 VSUBS 0.009217f
C558 B.n178 VSUBS 0.009217f
C559 B.n179 VSUBS 0.009217f
C560 B.n180 VSUBS 0.009217f
C561 B.n181 VSUBS 0.009217f
C562 B.n182 VSUBS 0.009217f
C563 B.n183 VSUBS 0.009217f
C564 B.n184 VSUBS 0.009217f
C565 B.n185 VSUBS 0.009217f
C566 B.n186 VSUBS 0.009217f
C567 B.n187 VSUBS 0.009217f
C568 B.n188 VSUBS 0.009217f
C569 B.n189 VSUBS 0.009217f
C570 B.n190 VSUBS 0.009217f
C571 B.n191 VSUBS 0.009217f
C572 B.n192 VSUBS 0.009217f
C573 B.n193 VSUBS 0.009217f
C574 B.n194 VSUBS 0.009217f
C575 B.n195 VSUBS 0.009217f
C576 B.n196 VSUBS 0.009217f
C577 B.n197 VSUBS 0.009217f
C578 B.n198 VSUBS 0.009217f
C579 B.n199 VSUBS 0.009217f
C580 B.n200 VSUBS 0.009217f
C581 B.n201 VSUBS 0.00637f
C582 B.n202 VSUBS 0.021354f
C583 B.n203 VSUBS 0.007455f
C584 B.n204 VSUBS 0.009217f
C585 B.n205 VSUBS 0.009217f
C586 B.n206 VSUBS 0.009217f
C587 B.n207 VSUBS 0.009217f
C588 B.n208 VSUBS 0.009217f
C589 B.n209 VSUBS 0.009217f
C590 B.n210 VSUBS 0.009217f
C591 B.n211 VSUBS 0.009217f
C592 B.n212 VSUBS 0.009217f
C593 B.n213 VSUBS 0.009217f
C594 B.n214 VSUBS 0.009217f
C595 B.t4 VSUBS 0.086429f
C596 B.t5 VSUBS 0.10395f
C597 B.t3 VSUBS 0.374546f
C598 B.n215 VSUBS 0.187977f
C599 B.n216 VSUBS 0.161535f
C600 B.n217 VSUBS 0.021354f
C601 B.n218 VSUBS 0.007455f
C602 B.n219 VSUBS 0.009217f
C603 B.n220 VSUBS 0.009217f
C604 B.n221 VSUBS 0.009217f
C605 B.n222 VSUBS 0.009217f
C606 B.n223 VSUBS 0.009217f
C607 B.n224 VSUBS 0.009217f
C608 B.n225 VSUBS 0.009217f
C609 B.n226 VSUBS 0.009217f
C610 B.n227 VSUBS 0.009217f
C611 B.n228 VSUBS 0.009217f
C612 B.n229 VSUBS 0.009217f
C613 B.n230 VSUBS 0.009217f
C614 B.n231 VSUBS 0.009217f
C615 B.n232 VSUBS 0.009217f
C616 B.n233 VSUBS 0.009217f
C617 B.n234 VSUBS 0.009217f
C618 B.n235 VSUBS 0.009217f
C619 B.n236 VSUBS 0.009217f
C620 B.n237 VSUBS 0.009217f
C621 B.n238 VSUBS 0.009217f
C622 B.n239 VSUBS 0.009217f
C623 B.n240 VSUBS 0.009217f
C624 B.n241 VSUBS 0.009217f
C625 B.n242 VSUBS 0.009217f
C626 B.n243 VSUBS 0.009217f
C627 B.n244 VSUBS 0.009217f
C628 B.n245 VSUBS 0.009217f
C629 B.n246 VSUBS 0.009217f
C630 B.n247 VSUBS 0.009217f
C631 B.n248 VSUBS 0.020987f
C632 B.n249 VSUBS 0.020987f
C633 B.n250 VSUBS 0.020217f
C634 B.n251 VSUBS 0.009217f
C635 B.n252 VSUBS 0.009217f
C636 B.n253 VSUBS 0.009217f
C637 B.n254 VSUBS 0.009217f
C638 B.n255 VSUBS 0.009217f
C639 B.n256 VSUBS 0.009217f
C640 B.n257 VSUBS 0.009217f
C641 B.n258 VSUBS 0.009217f
C642 B.n259 VSUBS 0.009217f
C643 B.n260 VSUBS 0.009217f
C644 B.n261 VSUBS 0.009217f
C645 B.n262 VSUBS 0.009217f
C646 B.n263 VSUBS 0.009217f
C647 B.n264 VSUBS 0.009217f
C648 B.n265 VSUBS 0.009217f
C649 B.n266 VSUBS 0.009217f
C650 B.n267 VSUBS 0.009217f
C651 B.n268 VSUBS 0.009217f
C652 B.n269 VSUBS 0.009217f
C653 B.n270 VSUBS 0.009217f
C654 B.n271 VSUBS 0.009217f
C655 B.n272 VSUBS 0.009217f
C656 B.n273 VSUBS 0.009217f
C657 B.n274 VSUBS 0.009217f
C658 B.n275 VSUBS 0.009217f
C659 B.n276 VSUBS 0.009217f
C660 B.n277 VSUBS 0.009217f
C661 B.n278 VSUBS 0.009217f
C662 B.n279 VSUBS 0.009217f
C663 B.n280 VSUBS 0.009217f
C664 B.n281 VSUBS 0.009217f
C665 B.n282 VSUBS 0.009217f
C666 B.n283 VSUBS 0.009217f
C667 B.n284 VSUBS 0.009217f
C668 B.n285 VSUBS 0.009217f
C669 B.n286 VSUBS 0.009217f
C670 B.n287 VSUBS 0.009217f
C671 B.n288 VSUBS 0.009217f
C672 B.n289 VSUBS 0.009217f
C673 B.n290 VSUBS 0.009217f
C674 B.n291 VSUBS 0.009217f
C675 B.n292 VSUBS 0.009217f
C676 B.n293 VSUBS 0.009217f
C677 B.n294 VSUBS 0.009217f
C678 B.n295 VSUBS 0.009217f
C679 B.n296 VSUBS 0.009217f
C680 B.n297 VSUBS 0.009217f
C681 B.n298 VSUBS 0.009217f
C682 B.n299 VSUBS 0.009217f
C683 B.n300 VSUBS 0.009217f
C684 B.n301 VSUBS 0.009217f
C685 B.n302 VSUBS 0.009217f
C686 B.n303 VSUBS 0.009217f
C687 B.n304 VSUBS 0.009217f
C688 B.n305 VSUBS 0.009217f
C689 B.n306 VSUBS 0.009217f
C690 B.n307 VSUBS 0.009217f
C691 B.n308 VSUBS 0.009217f
C692 B.n309 VSUBS 0.009217f
C693 B.n310 VSUBS 0.009217f
C694 B.n311 VSUBS 0.009217f
C695 B.n312 VSUBS 0.009217f
C696 B.n313 VSUBS 0.009217f
C697 B.n314 VSUBS 0.009217f
C698 B.n315 VSUBS 0.009217f
C699 B.n316 VSUBS 0.009217f
C700 B.n317 VSUBS 0.009217f
C701 B.n318 VSUBS 0.009217f
C702 B.n319 VSUBS 0.009217f
C703 B.n320 VSUBS 0.009217f
C704 B.n321 VSUBS 0.009217f
C705 B.n322 VSUBS 0.009217f
C706 B.n323 VSUBS 0.009217f
C707 B.n324 VSUBS 0.009217f
C708 B.n325 VSUBS 0.009217f
C709 B.n326 VSUBS 0.009217f
C710 B.n327 VSUBS 0.009217f
C711 B.n328 VSUBS 0.009217f
C712 B.n329 VSUBS 0.009217f
C713 B.n330 VSUBS 0.009217f
C714 B.n331 VSUBS 0.009217f
C715 B.n332 VSUBS 0.009217f
C716 B.n333 VSUBS 0.009217f
C717 B.n334 VSUBS 0.009217f
C718 B.n335 VSUBS 0.009217f
C719 B.n336 VSUBS 0.009217f
C720 B.n337 VSUBS 0.009217f
C721 B.n338 VSUBS 0.009217f
C722 B.n339 VSUBS 0.009217f
C723 B.n340 VSUBS 0.009217f
C724 B.n341 VSUBS 0.009217f
C725 B.n342 VSUBS 0.009217f
C726 B.n343 VSUBS 0.009217f
C727 B.n344 VSUBS 0.009217f
C728 B.n345 VSUBS 0.009217f
C729 B.n346 VSUBS 0.009217f
C730 B.n347 VSUBS 0.009217f
C731 B.n348 VSUBS 0.009217f
C732 B.n349 VSUBS 0.021386f
C733 B.n350 VSUBS 0.019818f
C734 B.n351 VSUBS 0.020987f
C735 B.n352 VSUBS 0.009217f
C736 B.n353 VSUBS 0.009217f
C737 B.n354 VSUBS 0.009217f
C738 B.n355 VSUBS 0.009217f
C739 B.n356 VSUBS 0.009217f
C740 B.n357 VSUBS 0.009217f
C741 B.n358 VSUBS 0.009217f
C742 B.n359 VSUBS 0.009217f
C743 B.n360 VSUBS 0.009217f
C744 B.n361 VSUBS 0.009217f
C745 B.n362 VSUBS 0.009217f
C746 B.n363 VSUBS 0.009217f
C747 B.n364 VSUBS 0.009217f
C748 B.n365 VSUBS 0.009217f
C749 B.n366 VSUBS 0.009217f
C750 B.n367 VSUBS 0.009217f
C751 B.n368 VSUBS 0.009217f
C752 B.n369 VSUBS 0.009217f
C753 B.n370 VSUBS 0.009217f
C754 B.n371 VSUBS 0.009217f
C755 B.n372 VSUBS 0.009217f
C756 B.n373 VSUBS 0.009217f
C757 B.n374 VSUBS 0.009217f
C758 B.n375 VSUBS 0.009217f
C759 B.n376 VSUBS 0.009217f
C760 B.n377 VSUBS 0.009217f
C761 B.n378 VSUBS 0.009217f
C762 B.n379 VSUBS 0.00637f
C763 B.n380 VSUBS 0.021354f
C764 B.n381 VSUBS 0.007455f
C765 B.n382 VSUBS 0.009217f
C766 B.n383 VSUBS 0.009217f
C767 B.n384 VSUBS 0.009217f
C768 B.n385 VSUBS 0.009217f
C769 B.n386 VSUBS 0.009217f
C770 B.n387 VSUBS 0.009217f
C771 B.n388 VSUBS 0.009217f
C772 B.n389 VSUBS 0.009217f
C773 B.n390 VSUBS 0.009217f
C774 B.n391 VSUBS 0.009217f
C775 B.n392 VSUBS 0.009217f
C776 B.n393 VSUBS 0.007455f
C777 B.n394 VSUBS 0.009217f
C778 B.n395 VSUBS 0.009217f
C779 B.n396 VSUBS 0.009217f
C780 B.n397 VSUBS 0.009217f
C781 B.n398 VSUBS 0.009217f
C782 B.n399 VSUBS 0.009217f
C783 B.n400 VSUBS 0.009217f
C784 B.n401 VSUBS 0.009217f
C785 B.n402 VSUBS 0.009217f
C786 B.n403 VSUBS 0.009217f
C787 B.n404 VSUBS 0.009217f
C788 B.n405 VSUBS 0.009217f
C789 B.n406 VSUBS 0.009217f
C790 B.n407 VSUBS 0.009217f
C791 B.n408 VSUBS 0.009217f
C792 B.n409 VSUBS 0.009217f
C793 B.n410 VSUBS 0.009217f
C794 B.n411 VSUBS 0.009217f
C795 B.n412 VSUBS 0.009217f
C796 B.n413 VSUBS 0.009217f
C797 B.n414 VSUBS 0.009217f
C798 B.n415 VSUBS 0.009217f
C799 B.n416 VSUBS 0.009217f
C800 B.n417 VSUBS 0.009217f
C801 B.n418 VSUBS 0.009217f
C802 B.n419 VSUBS 0.009217f
C803 B.n420 VSUBS 0.009217f
C804 B.n421 VSUBS 0.009217f
C805 B.n422 VSUBS 0.009217f
C806 B.n423 VSUBS 0.020987f
C807 B.n424 VSUBS 0.020987f
C808 B.n425 VSUBS 0.020217f
C809 B.n426 VSUBS 0.009217f
C810 B.n427 VSUBS 0.009217f
C811 B.n428 VSUBS 0.009217f
C812 B.n429 VSUBS 0.009217f
C813 B.n430 VSUBS 0.009217f
C814 B.n431 VSUBS 0.009217f
C815 B.n432 VSUBS 0.009217f
C816 B.n433 VSUBS 0.009217f
C817 B.n434 VSUBS 0.009217f
C818 B.n435 VSUBS 0.009217f
C819 B.n436 VSUBS 0.009217f
C820 B.n437 VSUBS 0.009217f
C821 B.n438 VSUBS 0.009217f
C822 B.n439 VSUBS 0.009217f
C823 B.n440 VSUBS 0.009217f
C824 B.n441 VSUBS 0.009217f
C825 B.n442 VSUBS 0.009217f
C826 B.n443 VSUBS 0.009217f
C827 B.n444 VSUBS 0.009217f
C828 B.n445 VSUBS 0.009217f
C829 B.n446 VSUBS 0.009217f
C830 B.n447 VSUBS 0.009217f
C831 B.n448 VSUBS 0.009217f
C832 B.n449 VSUBS 0.009217f
C833 B.n450 VSUBS 0.009217f
C834 B.n451 VSUBS 0.009217f
C835 B.n452 VSUBS 0.009217f
C836 B.n453 VSUBS 0.009217f
C837 B.n454 VSUBS 0.009217f
C838 B.n455 VSUBS 0.009217f
C839 B.n456 VSUBS 0.009217f
C840 B.n457 VSUBS 0.009217f
C841 B.n458 VSUBS 0.009217f
C842 B.n459 VSUBS 0.009217f
C843 B.n460 VSUBS 0.009217f
C844 B.n461 VSUBS 0.009217f
C845 B.n462 VSUBS 0.009217f
C846 B.n463 VSUBS 0.009217f
C847 B.n464 VSUBS 0.009217f
C848 B.n465 VSUBS 0.009217f
C849 B.n466 VSUBS 0.009217f
C850 B.n467 VSUBS 0.009217f
C851 B.n468 VSUBS 0.009217f
C852 B.n469 VSUBS 0.009217f
C853 B.n470 VSUBS 0.009217f
C854 B.n471 VSUBS 0.009217f
C855 B.n472 VSUBS 0.009217f
C856 B.n473 VSUBS 0.009217f
C857 B.n474 VSUBS 0.009217f
C858 B.n475 VSUBS 0.02087f
.ends

