* NGSPICE file created from diff_pair_sample_0735.ext - technology: sky130A

.subckt diff_pair_sample_0735 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t11 VP.t0 VDD1.t4 B.t0 sky130_fd_pr__nfet_01v8 ad=0.7194 pd=4.69 as=0.7194 ps=4.69 w=4.36 l=2.88
X1 VDD2.t5 VN.t0 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=1.7004 pd=9.5 as=0.7194 ps=4.69 w=4.36 l=2.88
X2 VDD1.t2 VP.t1 VTAIL.t10 B.t4 sky130_fd_pr__nfet_01v8 ad=0.7194 pd=4.69 as=1.7004 ps=9.5 w=4.36 l=2.88
X3 VTAIL.t2 VN.t1 VDD2.t4 B.t2 sky130_fd_pr__nfet_01v8 ad=0.7194 pd=4.69 as=0.7194 ps=4.69 w=4.36 l=2.88
X4 B.t19 B.t17 B.t18 B.t14 sky130_fd_pr__nfet_01v8 ad=1.7004 pd=9.5 as=0 ps=0 w=4.36 l=2.88
X5 VDD2.t3 VN.t2 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.7194 pd=4.69 as=1.7004 ps=9.5 w=4.36 l=2.88
X6 VDD1.t0 VP.t2 VTAIL.t9 B.t1 sky130_fd_pr__nfet_01v8 ad=0.7194 pd=4.69 as=1.7004 ps=9.5 w=4.36 l=2.88
X7 VDD1.t3 VP.t3 VTAIL.t8 B.t3 sky130_fd_pr__nfet_01v8 ad=1.7004 pd=9.5 as=0.7194 ps=4.69 w=4.36 l=2.88
X8 VTAIL.t0 VN.t3 VDD2.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=0.7194 pd=4.69 as=0.7194 ps=4.69 w=4.36 l=2.88
X9 B.t16 B.t13 B.t15 B.t14 sky130_fd_pr__nfet_01v8 ad=1.7004 pd=9.5 as=0 ps=0 w=4.36 l=2.88
X10 VDD2.t1 VN.t4 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=0.7194 pd=4.69 as=1.7004 ps=9.5 w=4.36 l=2.88
X11 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=1.7004 pd=9.5 as=0 ps=0 w=4.36 l=2.88
X12 VDD2.t0 VN.t5 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.7004 pd=9.5 as=0.7194 ps=4.69 w=4.36 l=2.88
X13 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=1.7004 pd=9.5 as=0 ps=0 w=4.36 l=2.88
X14 VTAIL.t7 VP.t4 VDD1.t5 B.t2 sky130_fd_pr__nfet_01v8 ad=0.7194 pd=4.69 as=0.7194 ps=4.69 w=4.36 l=2.88
X15 VDD1.t1 VP.t5 VTAIL.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=1.7004 pd=9.5 as=0.7194 ps=4.69 w=4.36 l=2.88
R0 VP.n13 VP.n10 161.3
R1 VP.n15 VP.n14 161.3
R2 VP.n16 VP.n9 161.3
R3 VP.n18 VP.n17 161.3
R4 VP.n19 VP.n8 161.3
R5 VP.n21 VP.n20 161.3
R6 VP.n43 VP.n42 161.3
R7 VP.n41 VP.n1 161.3
R8 VP.n40 VP.n39 161.3
R9 VP.n38 VP.n2 161.3
R10 VP.n37 VP.n36 161.3
R11 VP.n35 VP.n3 161.3
R12 VP.n33 VP.n32 161.3
R13 VP.n31 VP.n4 161.3
R14 VP.n30 VP.n29 161.3
R15 VP.n28 VP.n5 161.3
R16 VP.n27 VP.n26 161.3
R17 VP.n25 VP.n6 161.3
R18 VP.n11 VP.t3 68.3832
R19 VP.n24 VP.n23 67.6211
R20 VP.n44 VP.n0 67.6211
R21 VP.n22 VP.n7 67.6211
R22 VP.n12 VP.n11 61.7085
R23 VP.n29 VP.n28 54.6242
R24 VP.n40 VP.n2 54.6242
R25 VP.n18 VP.n9 54.6242
R26 VP.n24 VP.n22 44.117
R27 VP.n23 VP.t5 36.4852
R28 VP.n34 VP.t4 36.4852
R29 VP.n0 VP.t1 36.4852
R30 VP.n7 VP.t2 36.4852
R31 VP.n12 VP.t0 36.4852
R32 VP.n28 VP.n27 26.5299
R33 VP.n41 VP.n40 26.5299
R34 VP.n19 VP.n18 26.5299
R35 VP.n27 VP.n6 24.5923
R36 VP.n29 VP.n4 24.5923
R37 VP.n33 VP.n4 24.5923
R38 VP.n36 VP.n35 24.5923
R39 VP.n36 VP.n2 24.5923
R40 VP.n42 VP.n41 24.5923
R41 VP.n20 VP.n19 24.5923
R42 VP.n14 VP.n13 24.5923
R43 VP.n14 VP.n9 24.5923
R44 VP.n23 VP.n6 22.625
R45 VP.n42 VP.n0 22.625
R46 VP.n20 VP.n7 22.625
R47 VP.n34 VP.n33 12.2964
R48 VP.n35 VP.n34 12.2964
R49 VP.n13 VP.n12 12.2964
R50 VP.n11 VP.n10 5.34744
R51 VP.n22 VP.n21 0.354861
R52 VP.n25 VP.n24 0.354861
R53 VP.n44 VP.n43 0.354861
R54 VP VP.n44 0.267071
R55 VP.n15 VP.n10 0.189894
R56 VP.n16 VP.n15 0.189894
R57 VP.n17 VP.n16 0.189894
R58 VP.n17 VP.n8 0.189894
R59 VP.n21 VP.n8 0.189894
R60 VP.n26 VP.n25 0.189894
R61 VP.n26 VP.n5 0.189894
R62 VP.n30 VP.n5 0.189894
R63 VP.n31 VP.n30 0.189894
R64 VP.n32 VP.n31 0.189894
R65 VP.n32 VP.n3 0.189894
R66 VP.n37 VP.n3 0.189894
R67 VP.n38 VP.n37 0.189894
R68 VP.n39 VP.n38 0.189894
R69 VP.n39 VP.n1 0.189894
R70 VP.n43 VP.n1 0.189894
R71 VDD1 VDD1.t3 81.6964
R72 VDD1.n1 VDD1.t1 81.5826
R73 VDD1.n1 VDD1.n0 75.6577
R74 VDD1.n3 VDD1.n2 75.0213
R75 VDD1.n3 VDD1.n1 38.4341
R76 VDD1.n2 VDD1.t4 4.54178
R77 VDD1.n2 VDD1.t0 4.54178
R78 VDD1.n0 VDD1.t5 4.54178
R79 VDD1.n0 VDD1.t2 4.54178
R80 VDD1 VDD1.n3 0.634121
R81 VTAIL.n7 VTAIL.t4 62.884
R82 VTAIL.n10 VTAIL.t9 62.8837
R83 VTAIL.n11 VTAIL.t1 62.8837
R84 VTAIL.n2 VTAIL.t10 62.8837
R85 VTAIL.n9 VTAIL.n8 58.3427
R86 VTAIL.n6 VTAIL.n5 58.3427
R87 VTAIL.n1 VTAIL.n0 58.3425
R88 VTAIL.n4 VTAIL.n3 58.3425
R89 VTAIL.n6 VTAIL.n4 21.66
R90 VTAIL.n11 VTAIL.n10 18.8927
R91 VTAIL.n0 VTAIL.t3 4.54178
R92 VTAIL.n0 VTAIL.t0 4.54178
R93 VTAIL.n3 VTAIL.t6 4.54178
R94 VTAIL.n3 VTAIL.t7 4.54178
R95 VTAIL.n8 VTAIL.t8 4.54178
R96 VTAIL.n8 VTAIL.t11 4.54178
R97 VTAIL.n5 VTAIL.t5 4.54178
R98 VTAIL.n5 VTAIL.t2 4.54178
R99 VTAIL.n7 VTAIL.n6 2.76774
R100 VTAIL.n10 VTAIL.n9 2.76774
R101 VTAIL.n4 VTAIL.n2 2.76774
R102 VTAIL VTAIL.n11 2.01774
R103 VTAIL.n9 VTAIL.n7 1.85395
R104 VTAIL.n2 VTAIL.n1 1.85395
R105 VTAIL VTAIL.n1 0.7505
R106 B.n527 B.n526 585
R107 B.n529 B.n114 585
R108 B.n532 B.n531 585
R109 B.n533 B.n113 585
R110 B.n535 B.n534 585
R111 B.n537 B.n112 585
R112 B.n540 B.n539 585
R113 B.n541 B.n111 585
R114 B.n543 B.n542 585
R115 B.n545 B.n110 585
R116 B.n548 B.n547 585
R117 B.n549 B.n109 585
R118 B.n551 B.n550 585
R119 B.n553 B.n108 585
R120 B.n556 B.n555 585
R121 B.n557 B.n107 585
R122 B.n559 B.n558 585
R123 B.n561 B.n106 585
R124 B.n564 B.n563 585
R125 B.n566 B.n103 585
R126 B.n568 B.n567 585
R127 B.n570 B.n102 585
R128 B.n573 B.n572 585
R129 B.n574 B.n101 585
R130 B.n576 B.n575 585
R131 B.n578 B.n100 585
R132 B.n581 B.n580 585
R133 B.n582 B.n96 585
R134 B.n584 B.n583 585
R135 B.n586 B.n95 585
R136 B.n589 B.n588 585
R137 B.n590 B.n94 585
R138 B.n592 B.n591 585
R139 B.n594 B.n93 585
R140 B.n597 B.n596 585
R141 B.n598 B.n92 585
R142 B.n600 B.n599 585
R143 B.n602 B.n91 585
R144 B.n605 B.n604 585
R145 B.n606 B.n90 585
R146 B.n608 B.n607 585
R147 B.n610 B.n89 585
R148 B.n613 B.n612 585
R149 B.n614 B.n88 585
R150 B.n616 B.n615 585
R151 B.n618 B.n87 585
R152 B.n621 B.n620 585
R153 B.n622 B.n86 585
R154 B.n525 B.n84 585
R155 B.n625 B.n84 585
R156 B.n524 B.n83 585
R157 B.n626 B.n83 585
R158 B.n523 B.n82 585
R159 B.n627 B.n82 585
R160 B.n522 B.n521 585
R161 B.n521 B.n78 585
R162 B.n520 B.n77 585
R163 B.n633 B.n77 585
R164 B.n519 B.n76 585
R165 B.n634 B.n76 585
R166 B.n518 B.n75 585
R167 B.n635 B.n75 585
R168 B.n517 B.n516 585
R169 B.n516 B.n71 585
R170 B.n515 B.n70 585
R171 B.n641 B.n70 585
R172 B.n514 B.n69 585
R173 B.n642 B.n69 585
R174 B.n513 B.n68 585
R175 B.n643 B.n68 585
R176 B.n512 B.n511 585
R177 B.n511 B.n64 585
R178 B.n510 B.n63 585
R179 B.n649 B.n63 585
R180 B.n509 B.n62 585
R181 B.n650 B.n62 585
R182 B.n508 B.n61 585
R183 B.n651 B.n61 585
R184 B.n507 B.n506 585
R185 B.n506 B.n57 585
R186 B.n505 B.n56 585
R187 B.n657 B.n56 585
R188 B.n504 B.n55 585
R189 B.n658 B.n55 585
R190 B.n503 B.n54 585
R191 B.n659 B.n54 585
R192 B.n502 B.n501 585
R193 B.n501 B.n50 585
R194 B.n500 B.n49 585
R195 B.n665 B.n49 585
R196 B.n499 B.n48 585
R197 B.n666 B.n48 585
R198 B.n498 B.n47 585
R199 B.n667 B.n47 585
R200 B.n497 B.n496 585
R201 B.n496 B.n43 585
R202 B.n495 B.n42 585
R203 B.n673 B.n42 585
R204 B.n494 B.n41 585
R205 B.n674 B.n41 585
R206 B.n493 B.n40 585
R207 B.n675 B.n40 585
R208 B.n492 B.n491 585
R209 B.n491 B.n36 585
R210 B.n490 B.n35 585
R211 B.n681 B.n35 585
R212 B.n489 B.n34 585
R213 B.n682 B.n34 585
R214 B.n488 B.n33 585
R215 B.n683 B.n33 585
R216 B.n487 B.n486 585
R217 B.n486 B.n29 585
R218 B.n485 B.n28 585
R219 B.n689 B.n28 585
R220 B.n484 B.n27 585
R221 B.n690 B.n27 585
R222 B.n483 B.n26 585
R223 B.n691 B.n26 585
R224 B.n482 B.n481 585
R225 B.n481 B.n22 585
R226 B.n480 B.n21 585
R227 B.n697 B.n21 585
R228 B.n479 B.n20 585
R229 B.n698 B.n20 585
R230 B.n478 B.n19 585
R231 B.n699 B.n19 585
R232 B.n477 B.n476 585
R233 B.n476 B.n18 585
R234 B.n475 B.n14 585
R235 B.n705 B.n14 585
R236 B.n474 B.n13 585
R237 B.n706 B.n13 585
R238 B.n473 B.n12 585
R239 B.n707 B.n12 585
R240 B.n472 B.n471 585
R241 B.n471 B.n8 585
R242 B.n470 B.n7 585
R243 B.n713 B.n7 585
R244 B.n469 B.n6 585
R245 B.n714 B.n6 585
R246 B.n468 B.n5 585
R247 B.n715 B.n5 585
R248 B.n467 B.n466 585
R249 B.n466 B.n4 585
R250 B.n465 B.n115 585
R251 B.n465 B.n464 585
R252 B.n455 B.n116 585
R253 B.n117 B.n116 585
R254 B.n457 B.n456 585
R255 B.n458 B.n457 585
R256 B.n454 B.n122 585
R257 B.n122 B.n121 585
R258 B.n453 B.n452 585
R259 B.n452 B.n451 585
R260 B.n124 B.n123 585
R261 B.n444 B.n124 585
R262 B.n443 B.n442 585
R263 B.n445 B.n443 585
R264 B.n441 B.n129 585
R265 B.n129 B.n128 585
R266 B.n440 B.n439 585
R267 B.n439 B.n438 585
R268 B.n131 B.n130 585
R269 B.n132 B.n131 585
R270 B.n431 B.n430 585
R271 B.n432 B.n431 585
R272 B.n429 B.n137 585
R273 B.n137 B.n136 585
R274 B.n428 B.n427 585
R275 B.n427 B.n426 585
R276 B.n139 B.n138 585
R277 B.n140 B.n139 585
R278 B.n419 B.n418 585
R279 B.n420 B.n419 585
R280 B.n417 B.n145 585
R281 B.n145 B.n144 585
R282 B.n416 B.n415 585
R283 B.n415 B.n414 585
R284 B.n147 B.n146 585
R285 B.n148 B.n147 585
R286 B.n407 B.n406 585
R287 B.n408 B.n407 585
R288 B.n405 B.n153 585
R289 B.n153 B.n152 585
R290 B.n404 B.n403 585
R291 B.n403 B.n402 585
R292 B.n155 B.n154 585
R293 B.n156 B.n155 585
R294 B.n395 B.n394 585
R295 B.n396 B.n395 585
R296 B.n393 B.n161 585
R297 B.n161 B.n160 585
R298 B.n392 B.n391 585
R299 B.n391 B.n390 585
R300 B.n163 B.n162 585
R301 B.n164 B.n163 585
R302 B.n383 B.n382 585
R303 B.n384 B.n383 585
R304 B.n381 B.n169 585
R305 B.n169 B.n168 585
R306 B.n380 B.n379 585
R307 B.n379 B.n378 585
R308 B.n171 B.n170 585
R309 B.n172 B.n171 585
R310 B.n371 B.n370 585
R311 B.n372 B.n371 585
R312 B.n369 B.n177 585
R313 B.n177 B.n176 585
R314 B.n368 B.n367 585
R315 B.n367 B.n366 585
R316 B.n179 B.n178 585
R317 B.n180 B.n179 585
R318 B.n359 B.n358 585
R319 B.n360 B.n359 585
R320 B.n357 B.n185 585
R321 B.n185 B.n184 585
R322 B.n356 B.n355 585
R323 B.n355 B.n354 585
R324 B.n187 B.n186 585
R325 B.n188 B.n187 585
R326 B.n347 B.n346 585
R327 B.n348 B.n347 585
R328 B.n345 B.n193 585
R329 B.n193 B.n192 585
R330 B.n344 B.n343 585
R331 B.n343 B.n342 585
R332 B.n195 B.n194 585
R333 B.n196 B.n195 585
R334 B.n335 B.n334 585
R335 B.n336 B.n335 585
R336 B.n333 B.n201 585
R337 B.n201 B.n200 585
R338 B.n332 B.n331 585
R339 B.n331 B.n330 585
R340 B.n327 B.n205 585
R341 B.n326 B.n325 585
R342 B.n323 B.n206 585
R343 B.n323 B.n204 585
R344 B.n322 B.n321 585
R345 B.n320 B.n319 585
R346 B.n318 B.n208 585
R347 B.n316 B.n315 585
R348 B.n314 B.n209 585
R349 B.n313 B.n312 585
R350 B.n310 B.n210 585
R351 B.n308 B.n307 585
R352 B.n306 B.n211 585
R353 B.n305 B.n304 585
R354 B.n302 B.n212 585
R355 B.n300 B.n299 585
R356 B.n298 B.n213 585
R357 B.n297 B.n296 585
R358 B.n294 B.n214 585
R359 B.n292 B.n291 585
R360 B.n289 B.n215 585
R361 B.n288 B.n287 585
R362 B.n285 B.n218 585
R363 B.n283 B.n282 585
R364 B.n281 B.n219 585
R365 B.n280 B.n279 585
R366 B.n277 B.n220 585
R367 B.n275 B.n274 585
R368 B.n273 B.n221 585
R369 B.n272 B.n271 585
R370 B.n269 B.n268 585
R371 B.n267 B.n266 585
R372 B.n265 B.n226 585
R373 B.n263 B.n262 585
R374 B.n261 B.n227 585
R375 B.n260 B.n259 585
R376 B.n257 B.n228 585
R377 B.n255 B.n254 585
R378 B.n253 B.n229 585
R379 B.n252 B.n251 585
R380 B.n249 B.n230 585
R381 B.n247 B.n246 585
R382 B.n245 B.n231 585
R383 B.n244 B.n243 585
R384 B.n241 B.n232 585
R385 B.n239 B.n238 585
R386 B.n237 B.n233 585
R387 B.n236 B.n235 585
R388 B.n203 B.n202 585
R389 B.n204 B.n203 585
R390 B.n329 B.n328 585
R391 B.n330 B.n329 585
R392 B.n199 B.n198 585
R393 B.n200 B.n199 585
R394 B.n338 B.n337 585
R395 B.n337 B.n336 585
R396 B.n339 B.n197 585
R397 B.n197 B.n196 585
R398 B.n341 B.n340 585
R399 B.n342 B.n341 585
R400 B.n191 B.n190 585
R401 B.n192 B.n191 585
R402 B.n350 B.n349 585
R403 B.n349 B.n348 585
R404 B.n351 B.n189 585
R405 B.n189 B.n188 585
R406 B.n353 B.n352 585
R407 B.n354 B.n353 585
R408 B.n183 B.n182 585
R409 B.n184 B.n183 585
R410 B.n362 B.n361 585
R411 B.n361 B.n360 585
R412 B.n363 B.n181 585
R413 B.n181 B.n180 585
R414 B.n365 B.n364 585
R415 B.n366 B.n365 585
R416 B.n175 B.n174 585
R417 B.n176 B.n175 585
R418 B.n374 B.n373 585
R419 B.n373 B.n372 585
R420 B.n375 B.n173 585
R421 B.n173 B.n172 585
R422 B.n377 B.n376 585
R423 B.n378 B.n377 585
R424 B.n167 B.n166 585
R425 B.n168 B.n167 585
R426 B.n386 B.n385 585
R427 B.n385 B.n384 585
R428 B.n387 B.n165 585
R429 B.n165 B.n164 585
R430 B.n389 B.n388 585
R431 B.n390 B.n389 585
R432 B.n159 B.n158 585
R433 B.n160 B.n159 585
R434 B.n398 B.n397 585
R435 B.n397 B.n396 585
R436 B.n399 B.n157 585
R437 B.n157 B.n156 585
R438 B.n401 B.n400 585
R439 B.n402 B.n401 585
R440 B.n151 B.n150 585
R441 B.n152 B.n151 585
R442 B.n410 B.n409 585
R443 B.n409 B.n408 585
R444 B.n411 B.n149 585
R445 B.n149 B.n148 585
R446 B.n413 B.n412 585
R447 B.n414 B.n413 585
R448 B.n143 B.n142 585
R449 B.n144 B.n143 585
R450 B.n422 B.n421 585
R451 B.n421 B.n420 585
R452 B.n423 B.n141 585
R453 B.n141 B.n140 585
R454 B.n425 B.n424 585
R455 B.n426 B.n425 585
R456 B.n135 B.n134 585
R457 B.n136 B.n135 585
R458 B.n434 B.n433 585
R459 B.n433 B.n432 585
R460 B.n435 B.n133 585
R461 B.n133 B.n132 585
R462 B.n437 B.n436 585
R463 B.n438 B.n437 585
R464 B.n127 B.n126 585
R465 B.n128 B.n127 585
R466 B.n447 B.n446 585
R467 B.n446 B.n445 585
R468 B.n448 B.n125 585
R469 B.n444 B.n125 585
R470 B.n450 B.n449 585
R471 B.n451 B.n450 585
R472 B.n120 B.n119 585
R473 B.n121 B.n120 585
R474 B.n460 B.n459 585
R475 B.n459 B.n458 585
R476 B.n461 B.n118 585
R477 B.n118 B.n117 585
R478 B.n463 B.n462 585
R479 B.n464 B.n463 585
R480 B.n2 B.n0 585
R481 B.n4 B.n2 585
R482 B.n3 B.n1 585
R483 B.n714 B.n3 585
R484 B.n712 B.n711 585
R485 B.n713 B.n712 585
R486 B.n710 B.n9 585
R487 B.n9 B.n8 585
R488 B.n709 B.n708 585
R489 B.n708 B.n707 585
R490 B.n11 B.n10 585
R491 B.n706 B.n11 585
R492 B.n704 B.n703 585
R493 B.n705 B.n704 585
R494 B.n702 B.n15 585
R495 B.n18 B.n15 585
R496 B.n701 B.n700 585
R497 B.n700 B.n699 585
R498 B.n17 B.n16 585
R499 B.n698 B.n17 585
R500 B.n696 B.n695 585
R501 B.n697 B.n696 585
R502 B.n694 B.n23 585
R503 B.n23 B.n22 585
R504 B.n693 B.n692 585
R505 B.n692 B.n691 585
R506 B.n25 B.n24 585
R507 B.n690 B.n25 585
R508 B.n688 B.n687 585
R509 B.n689 B.n688 585
R510 B.n686 B.n30 585
R511 B.n30 B.n29 585
R512 B.n685 B.n684 585
R513 B.n684 B.n683 585
R514 B.n32 B.n31 585
R515 B.n682 B.n32 585
R516 B.n680 B.n679 585
R517 B.n681 B.n680 585
R518 B.n678 B.n37 585
R519 B.n37 B.n36 585
R520 B.n677 B.n676 585
R521 B.n676 B.n675 585
R522 B.n39 B.n38 585
R523 B.n674 B.n39 585
R524 B.n672 B.n671 585
R525 B.n673 B.n672 585
R526 B.n670 B.n44 585
R527 B.n44 B.n43 585
R528 B.n669 B.n668 585
R529 B.n668 B.n667 585
R530 B.n46 B.n45 585
R531 B.n666 B.n46 585
R532 B.n664 B.n663 585
R533 B.n665 B.n664 585
R534 B.n662 B.n51 585
R535 B.n51 B.n50 585
R536 B.n661 B.n660 585
R537 B.n660 B.n659 585
R538 B.n53 B.n52 585
R539 B.n658 B.n53 585
R540 B.n656 B.n655 585
R541 B.n657 B.n656 585
R542 B.n654 B.n58 585
R543 B.n58 B.n57 585
R544 B.n653 B.n652 585
R545 B.n652 B.n651 585
R546 B.n60 B.n59 585
R547 B.n650 B.n60 585
R548 B.n648 B.n647 585
R549 B.n649 B.n648 585
R550 B.n646 B.n65 585
R551 B.n65 B.n64 585
R552 B.n645 B.n644 585
R553 B.n644 B.n643 585
R554 B.n67 B.n66 585
R555 B.n642 B.n67 585
R556 B.n640 B.n639 585
R557 B.n641 B.n640 585
R558 B.n638 B.n72 585
R559 B.n72 B.n71 585
R560 B.n637 B.n636 585
R561 B.n636 B.n635 585
R562 B.n74 B.n73 585
R563 B.n634 B.n74 585
R564 B.n632 B.n631 585
R565 B.n633 B.n632 585
R566 B.n630 B.n79 585
R567 B.n79 B.n78 585
R568 B.n629 B.n628 585
R569 B.n628 B.n627 585
R570 B.n81 B.n80 585
R571 B.n626 B.n81 585
R572 B.n624 B.n623 585
R573 B.n625 B.n624 585
R574 B.n717 B.n716 585
R575 B.n716 B.n715 585
R576 B.n329 B.n205 468.476
R577 B.n624 B.n86 468.476
R578 B.n331 B.n203 468.476
R579 B.n527 B.n84 468.476
R580 B.n528 B.n85 256.663
R581 B.n530 B.n85 256.663
R582 B.n536 B.n85 256.663
R583 B.n538 B.n85 256.663
R584 B.n544 B.n85 256.663
R585 B.n546 B.n85 256.663
R586 B.n552 B.n85 256.663
R587 B.n554 B.n85 256.663
R588 B.n560 B.n85 256.663
R589 B.n562 B.n85 256.663
R590 B.n569 B.n85 256.663
R591 B.n571 B.n85 256.663
R592 B.n577 B.n85 256.663
R593 B.n579 B.n85 256.663
R594 B.n585 B.n85 256.663
R595 B.n587 B.n85 256.663
R596 B.n593 B.n85 256.663
R597 B.n595 B.n85 256.663
R598 B.n601 B.n85 256.663
R599 B.n603 B.n85 256.663
R600 B.n609 B.n85 256.663
R601 B.n611 B.n85 256.663
R602 B.n617 B.n85 256.663
R603 B.n619 B.n85 256.663
R604 B.n324 B.n204 256.663
R605 B.n207 B.n204 256.663
R606 B.n317 B.n204 256.663
R607 B.n311 B.n204 256.663
R608 B.n309 B.n204 256.663
R609 B.n303 B.n204 256.663
R610 B.n301 B.n204 256.663
R611 B.n295 B.n204 256.663
R612 B.n293 B.n204 256.663
R613 B.n286 B.n204 256.663
R614 B.n284 B.n204 256.663
R615 B.n278 B.n204 256.663
R616 B.n276 B.n204 256.663
R617 B.n270 B.n204 256.663
R618 B.n225 B.n204 256.663
R619 B.n264 B.n204 256.663
R620 B.n258 B.n204 256.663
R621 B.n256 B.n204 256.663
R622 B.n250 B.n204 256.663
R623 B.n248 B.n204 256.663
R624 B.n242 B.n204 256.663
R625 B.n240 B.n204 256.663
R626 B.n234 B.n204 256.663
R627 B.n222 B.t10 244.918
R628 B.n216 B.t6 244.918
R629 B.n97 B.t13 244.918
R630 B.n104 B.t17 244.918
R631 B.n329 B.n199 163.367
R632 B.n337 B.n199 163.367
R633 B.n337 B.n197 163.367
R634 B.n341 B.n197 163.367
R635 B.n341 B.n191 163.367
R636 B.n349 B.n191 163.367
R637 B.n349 B.n189 163.367
R638 B.n353 B.n189 163.367
R639 B.n353 B.n183 163.367
R640 B.n361 B.n183 163.367
R641 B.n361 B.n181 163.367
R642 B.n365 B.n181 163.367
R643 B.n365 B.n175 163.367
R644 B.n373 B.n175 163.367
R645 B.n373 B.n173 163.367
R646 B.n377 B.n173 163.367
R647 B.n377 B.n167 163.367
R648 B.n385 B.n167 163.367
R649 B.n385 B.n165 163.367
R650 B.n389 B.n165 163.367
R651 B.n389 B.n159 163.367
R652 B.n397 B.n159 163.367
R653 B.n397 B.n157 163.367
R654 B.n401 B.n157 163.367
R655 B.n401 B.n151 163.367
R656 B.n409 B.n151 163.367
R657 B.n409 B.n149 163.367
R658 B.n413 B.n149 163.367
R659 B.n413 B.n143 163.367
R660 B.n421 B.n143 163.367
R661 B.n421 B.n141 163.367
R662 B.n425 B.n141 163.367
R663 B.n425 B.n135 163.367
R664 B.n433 B.n135 163.367
R665 B.n433 B.n133 163.367
R666 B.n437 B.n133 163.367
R667 B.n437 B.n127 163.367
R668 B.n446 B.n127 163.367
R669 B.n446 B.n125 163.367
R670 B.n450 B.n125 163.367
R671 B.n450 B.n120 163.367
R672 B.n459 B.n120 163.367
R673 B.n459 B.n118 163.367
R674 B.n463 B.n118 163.367
R675 B.n463 B.n2 163.367
R676 B.n716 B.n2 163.367
R677 B.n716 B.n3 163.367
R678 B.n712 B.n3 163.367
R679 B.n712 B.n9 163.367
R680 B.n708 B.n9 163.367
R681 B.n708 B.n11 163.367
R682 B.n704 B.n11 163.367
R683 B.n704 B.n15 163.367
R684 B.n700 B.n15 163.367
R685 B.n700 B.n17 163.367
R686 B.n696 B.n17 163.367
R687 B.n696 B.n23 163.367
R688 B.n692 B.n23 163.367
R689 B.n692 B.n25 163.367
R690 B.n688 B.n25 163.367
R691 B.n688 B.n30 163.367
R692 B.n684 B.n30 163.367
R693 B.n684 B.n32 163.367
R694 B.n680 B.n32 163.367
R695 B.n680 B.n37 163.367
R696 B.n676 B.n37 163.367
R697 B.n676 B.n39 163.367
R698 B.n672 B.n39 163.367
R699 B.n672 B.n44 163.367
R700 B.n668 B.n44 163.367
R701 B.n668 B.n46 163.367
R702 B.n664 B.n46 163.367
R703 B.n664 B.n51 163.367
R704 B.n660 B.n51 163.367
R705 B.n660 B.n53 163.367
R706 B.n656 B.n53 163.367
R707 B.n656 B.n58 163.367
R708 B.n652 B.n58 163.367
R709 B.n652 B.n60 163.367
R710 B.n648 B.n60 163.367
R711 B.n648 B.n65 163.367
R712 B.n644 B.n65 163.367
R713 B.n644 B.n67 163.367
R714 B.n640 B.n67 163.367
R715 B.n640 B.n72 163.367
R716 B.n636 B.n72 163.367
R717 B.n636 B.n74 163.367
R718 B.n632 B.n74 163.367
R719 B.n632 B.n79 163.367
R720 B.n628 B.n79 163.367
R721 B.n628 B.n81 163.367
R722 B.n624 B.n81 163.367
R723 B.n325 B.n323 163.367
R724 B.n323 B.n322 163.367
R725 B.n319 B.n318 163.367
R726 B.n316 B.n209 163.367
R727 B.n312 B.n310 163.367
R728 B.n308 B.n211 163.367
R729 B.n304 B.n302 163.367
R730 B.n300 B.n213 163.367
R731 B.n296 B.n294 163.367
R732 B.n292 B.n215 163.367
R733 B.n287 B.n285 163.367
R734 B.n283 B.n219 163.367
R735 B.n279 B.n277 163.367
R736 B.n275 B.n221 163.367
R737 B.n271 B.n269 163.367
R738 B.n266 B.n265 163.367
R739 B.n263 B.n227 163.367
R740 B.n259 B.n257 163.367
R741 B.n255 B.n229 163.367
R742 B.n251 B.n249 163.367
R743 B.n247 B.n231 163.367
R744 B.n243 B.n241 163.367
R745 B.n239 B.n233 163.367
R746 B.n235 B.n203 163.367
R747 B.n331 B.n201 163.367
R748 B.n335 B.n201 163.367
R749 B.n335 B.n195 163.367
R750 B.n343 B.n195 163.367
R751 B.n343 B.n193 163.367
R752 B.n347 B.n193 163.367
R753 B.n347 B.n187 163.367
R754 B.n355 B.n187 163.367
R755 B.n355 B.n185 163.367
R756 B.n359 B.n185 163.367
R757 B.n359 B.n179 163.367
R758 B.n367 B.n179 163.367
R759 B.n367 B.n177 163.367
R760 B.n371 B.n177 163.367
R761 B.n371 B.n171 163.367
R762 B.n379 B.n171 163.367
R763 B.n379 B.n169 163.367
R764 B.n383 B.n169 163.367
R765 B.n383 B.n163 163.367
R766 B.n391 B.n163 163.367
R767 B.n391 B.n161 163.367
R768 B.n395 B.n161 163.367
R769 B.n395 B.n155 163.367
R770 B.n403 B.n155 163.367
R771 B.n403 B.n153 163.367
R772 B.n407 B.n153 163.367
R773 B.n407 B.n147 163.367
R774 B.n415 B.n147 163.367
R775 B.n415 B.n145 163.367
R776 B.n419 B.n145 163.367
R777 B.n419 B.n139 163.367
R778 B.n427 B.n139 163.367
R779 B.n427 B.n137 163.367
R780 B.n431 B.n137 163.367
R781 B.n431 B.n131 163.367
R782 B.n439 B.n131 163.367
R783 B.n439 B.n129 163.367
R784 B.n443 B.n129 163.367
R785 B.n443 B.n124 163.367
R786 B.n452 B.n124 163.367
R787 B.n452 B.n122 163.367
R788 B.n457 B.n122 163.367
R789 B.n457 B.n116 163.367
R790 B.n465 B.n116 163.367
R791 B.n466 B.n465 163.367
R792 B.n466 B.n5 163.367
R793 B.n6 B.n5 163.367
R794 B.n7 B.n6 163.367
R795 B.n471 B.n7 163.367
R796 B.n471 B.n12 163.367
R797 B.n13 B.n12 163.367
R798 B.n14 B.n13 163.367
R799 B.n476 B.n14 163.367
R800 B.n476 B.n19 163.367
R801 B.n20 B.n19 163.367
R802 B.n21 B.n20 163.367
R803 B.n481 B.n21 163.367
R804 B.n481 B.n26 163.367
R805 B.n27 B.n26 163.367
R806 B.n28 B.n27 163.367
R807 B.n486 B.n28 163.367
R808 B.n486 B.n33 163.367
R809 B.n34 B.n33 163.367
R810 B.n35 B.n34 163.367
R811 B.n491 B.n35 163.367
R812 B.n491 B.n40 163.367
R813 B.n41 B.n40 163.367
R814 B.n42 B.n41 163.367
R815 B.n496 B.n42 163.367
R816 B.n496 B.n47 163.367
R817 B.n48 B.n47 163.367
R818 B.n49 B.n48 163.367
R819 B.n501 B.n49 163.367
R820 B.n501 B.n54 163.367
R821 B.n55 B.n54 163.367
R822 B.n56 B.n55 163.367
R823 B.n506 B.n56 163.367
R824 B.n506 B.n61 163.367
R825 B.n62 B.n61 163.367
R826 B.n63 B.n62 163.367
R827 B.n511 B.n63 163.367
R828 B.n511 B.n68 163.367
R829 B.n69 B.n68 163.367
R830 B.n70 B.n69 163.367
R831 B.n516 B.n70 163.367
R832 B.n516 B.n75 163.367
R833 B.n76 B.n75 163.367
R834 B.n77 B.n76 163.367
R835 B.n521 B.n77 163.367
R836 B.n521 B.n82 163.367
R837 B.n83 B.n82 163.367
R838 B.n84 B.n83 163.367
R839 B.n620 B.n618 163.367
R840 B.n616 B.n88 163.367
R841 B.n612 B.n610 163.367
R842 B.n608 B.n90 163.367
R843 B.n604 B.n602 163.367
R844 B.n600 B.n92 163.367
R845 B.n596 B.n594 163.367
R846 B.n592 B.n94 163.367
R847 B.n588 B.n586 163.367
R848 B.n584 B.n96 163.367
R849 B.n580 B.n578 163.367
R850 B.n576 B.n101 163.367
R851 B.n572 B.n570 163.367
R852 B.n568 B.n103 163.367
R853 B.n563 B.n561 163.367
R854 B.n559 B.n107 163.367
R855 B.n555 B.n553 163.367
R856 B.n551 B.n109 163.367
R857 B.n547 B.n545 163.367
R858 B.n543 B.n111 163.367
R859 B.n539 B.n537 163.367
R860 B.n535 B.n113 163.367
R861 B.n531 B.n529 163.367
R862 B.n222 B.t12 138.641
R863 B.n104 B.t18 138.641
R864 B.n216 B.t9 138.637
R865 B.n97 B.t15 138.637
R866 B.n330 B.n204 131.292
R867 B.n625 B.n85 131.292
R868 B.n330 B.n200 77.6341
R869 B.n336 B.n200 77.6341
R870 B.n336 B.n196 77.6341
R871 B.n342 B.n196 77.6341
R872 B.n342 B.n192 77.6341
R873 B.n348 B.n192 77.6341
R874 B.n348 B.n188 77.6341
R875 B.n354 B.n188 77.6341
R876 B.n360 B.n184 77.6341
R877 B.n360 B.n180 77.6341
R878 B.n366 B.n180 77.6341
R879 B.n366 B.n176 77.6341
R880 B.n372 B.n176 77.6341
R881 B.n372 B.n172 77.6341
R882 B.n378 B.n172 77.6341
R883 B.n378 B.n168 77.6341
R884 B.n384 B.n168 77.6341
R885 B.n384 B.n164 77.6341
R886 B.n390 B.n164 77.6341
R887 B.n396 B.n160 77.6341
R888 B.n396 B.n156 77.6341
R889 B.n402 B.n156 77.6341
R890 B.n402 B.n152 77.6341
R891 B.n408 B.n152 77.6341
R892 B.n408 B.n148 77.6341
R893 B.n414 B.n148 77.6341
R894 B.n414 B.n144 77.6341
R895 B.n420 B.n144 77.6341
R896 B.n426 B.n140 77.6341
R897 B.n426 B.n136 77.6341
R898 B.n432 B.n136 77.6341
R899 B.n432 B.n132 77.6341
R900 B.n438 B.n132 77.6341
R901 B.n438 B.n128 77.6341
R902 B.n445 B.n128 77.6341
R903 B.n445 B.n444 77.6341
R904 B.n451 B.n121 77.6341
R905 B.n458 B.n121 77.6341
R906 B.n458 B.n117 77.6341
R907 B.n464 B.n117 77.6341
R908 B.n464 B.n4 77.6341
R909 B.n715 B.n4 77.6341
R910 B.n715 B.n714 77.6341
R911 B.n714 B.n713 77.6341
R912 B.n713 B.n8 77.6341
R913 B.n707 B.n8 77.6341
R914 B.n707 B.n706 77.6341
R915 B.n706 B.n705 77.6341
R916 B.n699 B.n18 77.6341
R917 B.n699 B.n698 77.6341
R918 B.n698 B.n697 77.6341
R919 B.n697 B.n22 77.6341
R920 B.n691 B.n22 77.6341
R921 B.n691 B.n690 77.6341
R922 B.n690 B.n689 77.6341
R923 B.n689 B.n29 77.6341
R924 B.n683 B.n682 77.6341
R925 B.n682 B.n681 77.6341
R926 B.n681 B.n36 77.6341
R927 B.n675 B.n36 77.6341
R928 B.n675 B.n674 77.6341
R929 B.n674 B.n673 77.6341
R930 B.n673 B.n43 77.6341
R931 B.n667 B.n43 77.6341
R932 B.n667 B.n666 77.6341
R933 B.n665 B.n50 77.6341
R934 B.n659 B.n50 77.6341
R935 B.n659 B.n658 77.6341
R936 B.n658 B.n657 77.6341
R937 B.n657 B.n57 77.6341
R938 B.n651 B.n57 77.6341
R939 B.n651 B.n650 77.6341
R940 B.n650 B.n649 77.6341
R941 B.n649 B.n64 77.6341
R942 B.n643 B.n64 77.6341
R943 B.n643 B.n642 77.6341
R944 B.n641 B.n71 77.6341
R945 B.n635 B.n71 77.6341
R946 B.n635 B.n634 77.6341
R947 B.n634 B.n633 77.6341
R948 B.n633 B.n78 77.6341
R949 B.n627 B.n78 77.6341
R950 B.n627 B.n626 77.6341
R951 B.n626 B.n625 77.6341
R952 B.n223 B.t11 76.3861
R953 B.n105 B.t19 76.3861
R954 B.n217 B.t8 76.3822
R955 B.n98 B.t16 76.3822
R956 B.n324 B.n205 71.676
R957 B.n322 B.n207 71.676
R958 B.n318 B.n317 71.676
R959 B.n311 B.n209 71.676
R960 B.n310 B.n309 71.676
R961 B.n303 B.n211 71.676
R962 B.n302 B.n301 71.676
R963 B.n295 B.n213 71.676
R964 B.n294 B.n293 71.676
R965 B.n286 B.n215 71.676
R966 B.n285 B.n284 71.676
R967 B.n278 B.n219 71.676
R968 B.n277 B.n276 71.676
R969 B.n270 B.n221 71.676
R970 B.n269 B.n225 71.676
R971 B.n265 B.n264 71.676
R972 B.n258 B.n227 71.676
R973 B.n257 B.n256 71.676
R974 B.n250 B.n229 71.676
R975 B.n249 B.n248 71.676
R976 B.n242 B.n231 71.676
R977 B.n241 B.n240 71.676
R978 B.n234 B.n233 71.676
R979 B.n619 B.n86 71.676
R980 B.n618 B.n617 71.676
R981 B.n611 B.n88 71.676
R982 B.n610 B.n609 71.676
R983 B.n603 B.n90 71.676
R984 B.n602 B.n601 71.676
R985 B.n595 B.n92 71.676
R986 B.n594 B.n593 71.676
R987 B.n587 B.n94 71.676
R988 B.n586 B.n585 71.676
R989 B.n579 B.n96 71.676
R990 B.n578 B.n577 71.676
R991 B.n571 B.n101 71.676
R992 B.n570 B.n569 71.676
R993 B.n562 B.n103 71.676
R994 B.n561 B.n560 71.676
R995 B.n554 B.n107 71.676
R996 B.n553 B.n552 71.676
R997 B.n546 B.n109 71.676
R998 B.n545 B.n544 71.676
R999 B.n538 B.n111 71.676
R1000 B.n537 B.n536 71.676
R1001 B.n530 B.n113 71.676
R1002 B.n529 B.n528 71.676
R1003 B.n528 B.n527 71.676
R1004 B.n531 B.n530 71.676
R1005 B.n536 B.n535 71.676
R1006 B.n539 B.n538 71.676
R1007 B.n544 B.n543 71.676
R1008 B.n547 B.n546 71.676
R1009 B.n552 B.n551 71.676
R1010 B.n555 B.n554 71.676
R1011 B.n560 B.n559 71.676
R1012 B.n563 B.n562 71.676
R1013 B.n569 B.n568 71.676
R1014 B.n572 B.n571 71.676
R1015 B.n577 B.n576 71.676
R1016 B.n580 B.n579 71.676
R1017 B.n585 B.n584 71.676
R1018 B.n588 B.n587 71.676
R1019 B.n593 B.n592 71.676
R1020 B.n596 B.n595 71.676
R1021 B.n601 B.n600 71.676
R1022 B.n604 B.n603 71.676
R1023 B.n609 B.n608 71.676
R1024 B.n612 B.n611 71.676
R1025 B.n617 B.n616 71.676
R1026 B.n620 B.n619 71.676
R1027 B.n325 B.n324 71.676
R1028 B.n319 B.n207 71.676
R1029 B.n317 B.n316 71.676
R1030 B.n312 B.n311 71.676
R1031 B.n309 B.n308 71.676
R1032 B.n304 B.n303 71.676
R1033 B.n301 B.n300 71.676
R1034 B.n296 B.n295 71.676
R1035 B.n293 B.n292 71.676
R1036 B.n287 B.n286 71.676
R1037 B.n284 B.n283 71.676
R1038 B.n279 B.n278 71.676
R1039 B.n276 B.n275 71.676
R1040 B.n271 B.n270 71.676
R1041 B.n266 B.n225 71.676
R1042 B.n264 B.n263 71.676
R1043 B.n259 B.n258 71.676
R1044 B.n256 B.n255 71.676
R1045 B.n251 B.n250 71.676
R1046 B.n248 B.n247 71.676
R1047 B.n243 B.n242 71.676
R1048 B.n240 B.n239 71.676
R1049 B.n235 B.n234 71.676
R1050 B.t7 B.n184 66.2174
R1051 B.n642 B.t14 66.2174
R1052 B.n223 B.n222 62.255
R1053 B.n217 B.n216 62.255
R1054 B.n98 B.n97 62.255
R1055 B.n105 B.n104 62.255
R1056 B.n390 B.t5 61.6507
R1057 B.t1 B.n665 61.6507
R1058 B.n224 B.n223 59.5399
R1059 B.n290 B.n217 59.5399
R1060 B.n99 B.n98 59.5399
R1061 B.n565 B.n105 59.5399
R1062 B.t2 B.n140 59.3674
R1063 B.t0 B.n29 59.3674
R1064 B.n444 B.t4 52.5174
R1065 B.n18 B.t3 52.5174
R1066 B.n623 B.n622 30.4395
R1067 B.n526 B.n525 30.4395
R1068 B.n332 B.n202 30.4395
R1069 B.n328 B.n327 30.4395
R1070 B.n451 B.t4 25.1173
R1071 B.n705 B.t3 25.1173
R1072 B.n420 B.t2 18.2672
R1073 B.n683 B.t0 18.2672
R1074 B B.n717 18.0485
R1075 B.t5 B.n160 15.9839
R1076 B.n666 B.t1 15.9839
R1077 B.n354 B.t7 11.4172
R1078 B.t14 B.n641 11.4172
R1079 B.n622 B.n621 10.6151
R1080 B.n621 B.n87 10.6151
R1081 B.n615 B.n87 10.6151
R1082 B.n615 B.n614 10.6151
R1083 B.n614 B.n613 10.6151
R1084 B.n613 B.n89 10.6151
R1085 B.n607 B.n89 10.6151
R1086 B.n607 B.n606 10.6151
R1087 B.n606 B.n605 10.6151
R1088 B.n605 B.n91 10.6151
R1089 B.n599 B.n91 10.6151
R1090 B.n599 B.n598 10.6151
R1091 B.n598 B.n597 10.6151
R1092 B.n597 B.n93 10.6151
R1093 B.n591 B.n93 10.6151
R1094 B.n591 B.n590 10.6151
R1095 B.n590 B.n589 10.6151
R1096 B.n589 B.n95 10.6151
R1097 B.n583 B.n582 10.6151
R1098 B.n582 B.n581 10.6151
R1099 B.n581 B.n100 10.6151
R1100 B.n575 B.n100 10.6151
R1101 B.n575 B.n574 10.6151
R1102 B.n574 B.n573 10.6151
R1103 B.n573 B.n102 10.6151
R1104 B.n567 B.n102 10.6151
R1105 B.n567 B.n566 10.6151
R1106 B.n564 B.n106 10.6151
R1107 B.n558 B.n106 10.6151
R1108 B.n558 B.n557 10.6151
R1109 B.n557 B.n556 10.6151
R1110 B.n556 B.n108 10.6151
R1111 B.n550 B.n108 10.6151
R1112 B.n550 B.n549 10.6151
R1113 B.n549 B.n548 10.6151
R1114 B.n548 B.n110 10.6151
R1115 B.n542 B.n110 10.6151
R1116 B.n542 B.n541 10.6151
R1117 B.n541 B.n540 10.6151
R1118 B.n540 B.n112 10.6151
R1119 B.n534 B.n112 10.6151
R1120 B.n534 B.n533 10.6151
R1121 B.n533 B.n532 10.6151
R1122 B.n532 B.n114 10.6151
R1123 B.n526 B.n114 10.6151
R1124 B.n333 B.n332 10.6151
R1125 B.n334 B.n333 10.6151
R1126 B.n334 B.n194 10.6151
R1127 B.n344 B.n194 10.6151
R1128 B.n345 B.n344 10.6151
R1129 B.n346 B.n345 10.6151
R1130 B.n346 B.n186 10.6151
R1131 B.n356 B.n186 10.6151
R1132 B.n357 B.n356 10.6151
R1133 B.n358 B.n357 10.6151
R1134 B.n358 B.n178 10.6151
R1135 B.n368 B.n178 10.6151
R1136 B.n369 B.n368 10.6151
R1137 B.n370 B.n369 10.6151
R1138 B.n370 B.n170 10.6151
R1139 B.n380 B.n170 10.6151
R1140 B.n381 B.n380 10.6151
R1141 B.n382 B.n381 10.6151
R1142 B.n382 B.n162 10.6151
R1143 B.n392 B.n162 10.6151
R1144 B.n393 B.n392 10.6151
R1145 B.n394 B.n393 10.6151
R1146 B.n394 B.n154 10.6151
R1147 B.n404 B.n154 10.6151
R1148 B.n405 B.n404 10.6151
R1149 B.n406 B.n405 10.6151
R1150 B.n406 B.n146 10.6151
R1151 B.n416 B.n146 10.6151
R1152 B.n417 B.n416 10.6151
R1153 B.n418 B.n417 10.6151
R1154 B.n418 B.n138 10.6151
R1155 B.n428 B.n138 10.6151
R1156 B.n429 B.n428 10.6151
R1157 B.n430 B.n429 10.6151
R1158 B.n430 B.n130 10.6151
R1159 B.n440 B.n130 10.6151
R1160 B.n441 B.n440 10.6151
R1161 B.n442 B.n441 10.6151
R1162 B.n442 B.n123 10.6151
R1163 B.n453 B.n123 10.6151
R1164 B.n454 B.n453 10.6151
R1165 B.n456 B.n454 10.6151
R1166 B.n456 B.n455 10.6151
R1167 B.n455 B.n115 10.6151
R1168 B.n467 B.n115 10.6151
R1169 B.n468 B.n467 10.6151
R1170 B.n469 B.n468 10.6151
R1171 B.n470 B.n469 10.6151
R1172 B.n472 B.n470 10.6151
R1173 B.n473 B.n472 10.6151
R1174 B.n474 B.n473 10.6151
R1175 B.n475 B.n474 10.6151
R1176 B.n477 B.n475 10.6151
R1177 B.n478 B.n477 10.6151
R1178 B.n479 B.n478 10.6151
R1179 B.n480 B.n479 10.6151
R1180 B.n482 B.n480 10.6151
R1181 B.n483 B.n482 10.6151
R1182 B.n484 B.n483 10.6151
R1183 B.n485 B.n484 10.6151
R1184 B.n487 B.n485 10.6151
R1185 B.n488 B.n487 10.6151
R1186 B.n489 B.n488 10.6151
R1187 B.n490 B.n489 10.6151
R1188 B.n492 B.n490 10.6151
R1189 B.n493 B.n492 10.6151
R1190 B.n494 B.n493 10.6151
R1191 B.n495 B.n494 10.6151
R1192 B.n497 B.n495 10.6151
R1193 B.n498 B.n497 10.6151
R1194 B.n499 B.n498 10.6151
R1195 B.n500 B.n499 10.6151
R1196 B.n502 B.n500 10.6151
R1197 B.n503 B.n502 10.6151
R1198 B.n504 B.n503 10.6151
R1199 B.n505 B.n504 10.6151
R1200 B.n507 B.n505 10.6151
R1201 B.n508 B.n507 10.6151
R1202 B.n509 B.n508 10.6151
R1203 B.n510 B.n509 10.6151
R1204 B.n512 B.n510 10.6151
R1205 B.n513 B.n512 10.6151
R1206 B.n514 B.n513 10.6151
R1207 B.n515 B.n514 10.6151
R1208 B.n517 B.n515 10.6151
R1209 B.n518 B.n517 10.6151
R1210 B.n519 B.n518 10.6151
R1211 B.n520 B.n519 10.6151
R1212 B.n522 B.n520 10.6151
R1213 B.n523 B.n522 10.6151
R1214 B.n524 B.n523 10.6151
R1215 B.n525 B.n524 10.6151
R1216 B.n327 B.n326 10.6151
R1217 B.n326 B.n206 10.6151
R1218 B.n321 B.n206 10.6151
R1219 B.n321 B.n320 10.6151
R1220 B.n320 B.n208 10.6151
R1221 B.n315 B.n208 10.6151
R1222 B.n315 B.n314 10.6151
R1223 B.n314 B.n313 10.6151
R1224 B.n313 B.n210 10.6151
R1225 B.n307 B.n210 10.6151
R1226 B.n307 B.n306 10.6151
R1227 B.n306 B.n305 10.6151
R1228 B.n305 B.n212 10.6151
R1229 B.n299 B.n212 10.6151
R1230 B.n299 B.n298 10.6151
R1231 B.n298 B.n297 10.6151
R1232 B.n297 B.n214 10.6151
R1233 B.n291 B.n214 10.6151
R1234 B.n289 B.n288 10.6151
R1235 B.n288 B.n218 10.6151
R1236 B.n282 B.n218 10.6151
R1237 B.n282 B.n281 10.6151
R1238 B.n281 B.n280 10.6151
R1239 B.n280 B.n220 10.6151
R1240 B.n274 B.n220 10.6151
R1241 B.n274 B.n273 10.6151
R1242 B.n273 B.n272 10.6151
R1243 B.n268 B.n267 10.6151
R1244 B.n267 B.n226 10.6151
R1245 B.n262 B.n226 10.6151
R1246 B.n262 B.n261 10.6151
R1247 B.n261 B.n260 10.6151
R1248 B.n260 B.n228 10.6151
R1249 B.n254 B.n228 10.6151
R1250 B.n254 B.n253 10.6151
R1251 B.n253 B.n252 10.6151
R1252 B.n252 B.n230 10.6151
R1253 B.n246 B.n230 10.6151
R1254 B.n246 B.n245 10.6151
R1255 B.n245 B.n244 10.6151
R1256 B.n244 B.n232 10.6151
R1257 B.n238 B.n232 10.6151
R1258 B.n238 B.n237 10.6151
R1259 B.n237 B.n236 10.6151
R1260 B.n236 B.n202 10.6151
R1261 B.n328 B.n198 10.6151
R1262 B.n338 B.n198 10.6151
R1263 B.n339 B.n338 10.6151
R1264 B.n340 B.n339 10.6151
R1265 B.n340 B.n190 10.6151
R1266 B.n350 B.n190 10.6151
R1267 B.n351 B.n350 10.6151
R1268 B.n352 B.n351 10.6151
R1269 B.n352 B.n182 10.6151
R1270 B.n362 B.n182 10.6151
R1271 B.n363 B.n362 10.6151
R1272 B.n364 B.n363 10.6151
R1273 B.n364 B.n174 10.6151
R1274 B.n374 B.n174 10.6151
R1275 B.n375 B.n374 10.6151
R1276 B.n376 B.n375 10.6151
R1277 B.n376 B.n166 10.6151
R1278 B.n386 B.n166 10.6151
R1279 B.n387 B.n386 10.6151
R1280 B.n388 B.n387 10.6151
R1281 B.n388 B.n158 10.6151
R1282 B.n398 B.n158 10.6151
R1283 B.n399 B.n398 10.6151
R1284 B.n400 B.n399 10.6151
R1285 B.n400 B.n150 10.6151
R1286 B.n410 B.n150 10.6151
R1287 B.n411 B.n410 10.6151
R1288 B.n412 B.n411 10.6151
R1289 B.n412 B.n142 10.6151
R1290 B.n422 B.n142 10.6151
R1291 B.n423 B.n422 10.6151
R1292 B.n424 B.n423 10.6151
R1293 B.n424 B.n134 10.6151
R1294 B.n434 B.n134 10.6151
R1295 B.n435 B.n434 10.6151
R1296 B.n436 B.n435 10.6151
R1297 B.n436 B.n126 10.6151
R1298 B.n447 B.n126 10.6151
R1299 B.n448 B.n447 10.6151
R1300 B.n449 B.n448 10.6151
R1301 B.n449 B.n119 10.6151
R1302 B.n460 B.n119 10.6151
R1303 B.n461 B.n460 10.6151
R1304 B.n462 B.n461 10.6151
R1305 B.n462 B.n0 10.6151
R1306 B.n711 B.n1 10.6151
R1307 B.n711 B.n710 10.6151
R1308 B.n710 B.n709 10.6151
R1309 B.n709 B.n10 10.6151
R1310 B.n703 B.n10 10.6151
R1311 B.n703 B.n702 10.6151
R1312 B.n702 B.n701 10.6151
R1313 B.n701 B.n16 10.6151
R1314 B.n695 B.n16 10.6151
R1315 B.n695 B.n694 10.6151
R1316 B.n694 B.n693 10.6151
R1317 B.n693 B.n24 10.6151
R1318 B.n687 B.n24 10.6151
R1319 B.n687 B.n686 10.6151
R1320 B.n686 B.n685 10.6151
R1321 B.n685 B.n31 10.6151
R1322 B.n679 B.n31 10.6151
R1323 B.n679 B.n678 10.6151
R1324 B.n678 B.n677 10.6151
R1325 B.n677 B.n38 10.6151
R1326 B.n671 B.n38 10.6151
R1327 B.n671 B.n670 10.6151
R1328 B.n670 B.n669 10.6151
R1329 B.n669 B.n45 10.6151
R1330 B.n663 B.n45 10.6151
R1331 B.n663 B.n662 10.6151
R1332 B.n662 B.n661 10.6151
R1333 B.n661 B.n52 10.6151
R1334 B.n655 B.n52 10.6151
R1335 B.n655 B.n654 10.6151
R1336 B.n654 B.n653 10.6151
R1337 B.n653 B.n59 10.6151
R1338 B.n647 B.n59 10.6151
R1339 B.n647 B.n646 10.6151
R1340 B.n646 B.n645 10.6151
R1341 B.n645 B.n66 10.6151
R1342 B.n639 B.n66 10.6151
R1343 B.n639 B.n638 10.6151
R1344 B.n638 B.n637 10.6151
R1345 B.n637 B.n73 10.6151
R1346 B.n631 B.n73 10.6151
R1347 B.n631 B.n630 10.6151
R1348 B.n630 B.n629 10.6151
R1349 B.n629 B.n80 10.6151
R1350 B.n623 B.n80 10.6151
R1351 B.n99 B.n95 9.36635
R1352 B.n565 B.n564 9.36635
R1353 B.n291 B.n290 9.36635
R1354 B.n268 B.n224 9.36635
R1355 B.n717 B.n0 2.81026
R1356 B.n717 B.n1 2.81026
R1357 B.n583 B.n99 1.24928
R1358 B.n566 B.n565 1.24928
R1359 B.n290 B.n289 1.24928
R1360 B.n272 B.n224 1.24928
R1361 VN.n30 VN.n29 161.3
R1362 VN.n28 VN.n17 161.3
R1363 VN.n27 VN.n26 161.3
R1364 VN.n25 VN.n18 161.3
R1365 VN.n24 VN.n23 161.3
R1366 VN.n22 VN.n19 161.3
R1367 VN.n14 VN.n13 161.3
R1368 VN.n12 VN.n1 161.3
R1369 VN.n11 VN.n10 161.3
R1370 VN.n9 VN.n2 161.3
R1371 VN.n8 VN.n7 161.3
R1372 VN.n6 VN.n3 161.3
R1373 VN.n20 VN.t4 68.3835
R1374 VN.n4 VN.t5 68.3835
R1375 VN.n15 VN.n0 67.6211
R1376 VN.n31 VN.n16 67.6211
R1377 VN.n5 VN.n4 61.7085
R1378 VN.n21 VN.n20 61.7085
R1379 VN.n11 VN.n2 54.6242
R1380 VN.n27 VN.n18 54.6242
R1381 VN VN.n31 44.2822
R1382 VN.n5 VN.t3 36.4852
R1383 VN.n0 VN.t2 36.4852
R1384 VN.n21 VN.t1 36.4852
R1385 VN.n16 VN.t0 36.4852
R1386 VN.n12 VN.n11 26.5299
R1387 VN.n28 VN.n27 26.5299
R1388 VN.n7 VN.n6 24.5923
R1389 VN.n7 VN.n2 24.5923
R1390 VN.n13 VN.n12 24.5923
R1391 VN.n23 VN.n18 24.5923
R1392 VN.n23 VN.n22 24.5923
R1393 VN.n29 VN.n28 24.5923
R1394 VN.n13 VN.n0 22.625
R1395 VN.n29 VN.n16 22.625
R1396 VN.n6 VN.n5 12.2964
R1397 VN.n22 VN.n21 12.2964
R1398 VN.n4 VN.n3 5.34748
R1399 VN.n20 VN.n19 5.34748
R1400 VN.n31 VN.n30 0.354861
R1401 VN.n15 VN.n14 0.354861
R1402 VN VN.n15 0.267071
R1403 VN.n30 VN.n17 0.189894
R1404 VN.n26 VN.n17 0.189894
R1405 VN.n26 VN.n25 0.189894
R1406 VN.n25 VN.n24 0.189894
R1407 VN.n24 VN.n19 0.189894
R1408 VN.n8 VN.n3 0.189894
R1409 VN.n9 VN.n8 0.189894
R1410 VN.n10 VN.n9 0.189894
R1411 VN.n10 VN.n1 0.189894
R1412 VN.n14 VN.n1 0.189894
R1413 VDD2.n1 VDD2.t0 81.5826
R1414 VDD2.n2 VDD2.t5 79.5627
R1415 VDD2.n1 VDD2.n0 75.6577
R1416 VDD2 VDD2.n3 75.6549
R1417 VDD2.n2 VDD2.n1 36.4674
R1418 VDD2.n3 VDD2.t4 4.54178
R1419 VDD2.n3 VDD2.t1 4.54178
R1420 VDD2.n0 VDD2.t2 4.54178
R1421 VDD2.n0 VDD2.t3 4.54178
R1422 VDD2 VDD2.n2 2.13412
C0 VDD2 VN 2.73813f
C1 VDD1 VP 3.06649f
C2 VP VTAIL 3.50767f
C3 VDD1 VTAIL 5.12468f
C4 VP VN 5.78651f
C5 VDD1 VN 0.15558f
C6 VTAIL VN 3.4935f
C7 VDD2 VP 0.486448f
C8 VDD1 VDD2 1.51564f
C9 VDD2 VTAIL 5.17928f
C10 VDD2 B 4.83805f
C11 VDD1 B 5.169194f
C12 VTAIL B 4.568295f
C13 VN B 12.996921f
C14 VP B 11.643878f
C15 VDD2.t0 B 0.779376f
C16 VDD2.t2 B 0.075935f
C17 VDD2.t3 B 0.075935f
C18 VDD2.n0 B 0.608771f
C19 VDD2.n1 B 2.23377f
C20 VDD2.t5 B 0.770265f
C21 VDD2.n2 B 1.97855f
C22 VDD2.t4 B 0.075935f
C23 VDD2.t1 B 0.075935f
C24 VDD2.n3 B 0.608746f
C25 VN.t2 B 0.855626f
C26 VN.n0 B 0.437175f
C27 VN.n1 B 0.026327f
C28 VN.n2 B 0.045641f
C29 VN.n3 B 0.279774f
C30 VN.t3 B 0.855626f
C31 VN.t5 B 1.09187f
C32 VN.n4 B 0.400227f
C33 VN.n5 B 0.414337f
C34 VN.n6 B 0.036771f
C35 VN.n7 B 0.048821f
C36 VN.n8 B 0.026327f
C37 VN.n9 B 0.026327f
C38 VN.n10 B 0.026327f
C39 VN.n11 B 0.029281f
C40 VN.n12 B 0.050441f
C41 VN.n13 B 0.046893f
C42 VN.n14 B 0.042485f
C43 VN.n15 B 0.050694f
C44 VN.t0 B 0.855626f
C45 VN.n16 B 0.437175f
C46 VN.n17 B 0.026327f
C47 VN.n18 B 0.045641f
C48 VN.n19 B 0.279774f
C49 VN.t1 B 0.855626f
C50 VN.t4 B 1.09187f
C51 VN.n20 B 0.400227f
C52 VN.n21 B 0.414337f
C53 VN.n22 B 0.036771f
C54 VN.n23 B 0.048821f
C55 VN.n24 B 0.026327f
C56 VN.n25 B 0.026327f
C57 VN.n26 B 0.026327f
C58 VN.n27 B 0.029281f
C59 VN.n28 B 0.050441f
C60 VN.n29 B 0.046893f
C61 VN.n30 B 0.042485f
C62 VN.n31 B 1.24173f
C63 VTAIL.t3 B 0.101301f
C64 VTAIL.t0 B 0.101301f
C65 VTAIL.n0 B 0.742822f
C66 VTAIL.n1 B 0.502566f
C67 VTAIL.t10 B 0.952815f
C68 VTAIL.n2 B 0.759958f
C69 VTAIL.t6 B 0.101301f
C70 VTAIL.t7 B 0.101301f
C71 VTAIL.n3 B 0.742822f
C72 VTAIL.n4 B 1.79789f
C73 VTAIL.t5 B 0.101301f
C74 VTAIL.t2 B 0.101301f
C75 VTAIL.n5 B 0.742826f
C76 VTAIL.n6 B 1.79788f
C77 VTAIL.t4 B 0.952819f
C78 VTAIL.n7 B 0.759954f
C79 VTAIL.t8 B 0.101301f
C80 VTAIL.t11 B 0.101301f
C81 VTAIL.n8 B 0.742826f
C82 VTAIL.n9 B 0.693673f
C83 VTAIL.t9 B 0.952815f
C84 VTAIL.n10 B 1.602f
C85 VTAIL.t1 B 0.952815f
C86 VTAIL.n11 B 1.53095f
C87 VDD1.t3 B 0.801446f
C88 VDD1.t1 B 0.800722f
C89 VDD1.t5 B 0.078015f
C90 VDD1.t2 B 0.078015f
C91 VDD1.n0 B 0.625444f
C92 VDD1.n1 B 2.40687f
C93 VDD1.t4 B 0.078015f
C94 VDD1.t0 B 0.078015f
C95 VDD1.n2 B 0.621772f
C96 VDD1.n3 B 2.05373f
C97 VP.t1 B 0.886882f
C98 VP.n0 B 0.453146f
C99 VP.n1 B 0.027289f
C100 VP.n2 B 0.047308f
C101 VP.n3 B 0.027289f
C102 VP.t4 B 0.886882f
C103 VP.n4 B 0.050605f
C104 VP.n5 B 0.027289f
C105 VP.n6 B 0.048606f
C106 VP.t2 B 0.886882f
C107 VP.n7 B 0.453146f
C108 VP.n8 B 0.027289f
C109 VP.n9 B 0.047308f
C110 VP.n10 B 0.289995f
C111 VP.t0 B 0.886882f
C112 VP.t3 B 1.13175f
C113 VP.n11 B 0.414848f
C114 VP.n12 B 0.429473f
C115 VP.n13 B 0.038114f
C116 VP.n14 B 0.050605f
C117 VP.n15 B 0.027289f
C118 VP.n16 B 0.027289f
C119 VP.n17 B 0.027289f
C120 VP.n18 B 0.03035f
C121 VP.n19 B 0.052283f
C122 VP.n20 B 0.048606f
C123 VP.n21 B 0.044037f
C124 VP.n22 B 1.27541f
C125 VP.t5 B 0.886882f
C126 VP.n23 B 0.453146f
C127 VP.n24 B 1.29771f
C128 VP.n25 B 0.044037f
C129 VP.n26 B 0.027289f
C130 VP.n27 B 0.052283f
C131 VP.n28 B 0.03035f
C132 VP.n29 B 0.047308f
C133 VP.n30 B 0.027289f
C134 VP.n31 B 0.027289f
C135 VP.n32 B 0.027289f
C136 VP.n33 B 0.038114f
C137 VP.n34 B 0.345082f
C138 VP.n35 B 0.038114f
C139 VP.n36 B 0.050605f
C140 VP.n37 B 0.027289f
C141 VP.n38 B 0.027289f
C142 VP.n39 B 0.027289f
C143 VP.n40 B 0.03035f
C144 VP.n41 B 0.052283f
C145 VP.n42 B 0.048606f
C146 VP.n43 B 0.044037f
C147 VP.n44 B 0.052546f
.ends

