* NGSPICE file created from diff_pair_sample_0093.ext - technology: sky130A

.subckt diff_pair_sample_0093 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t9 w_n4522_n1170# sky130_fd_pr__pfet_01v8 ad=0.16665 pd=1.34 as=0.3939 ps=2.8 w=1.01 l=2.63
X1 B.t11 B.t9 B.t10 w_n4522_n1170# sky130_fd_pr__pfet_01v8 ad=0.3939 pd=2.8 as=0 ps=0 w=1.01 l=2.63
X2 VDD1.t8 VP.t1 VTAIL.t8 w_n4522_n1170# sky130_fd_pr__pfet_01v8 ad=0.16665 pd=1.34 as=0.3939 ps=2.8 w=1.01 l=2.63
X3 VTAIL.t5 VP.t2 VDD1.t7 w_n4522_n1170# sky130_fd_pr__pfet_01v8 ad=0.16665 pd=1.34 as=0.16665 ps=1.34 w=1.01 l=2.63
X4 VDD2.t9 VN.t0 VTAIL.t19 w_n4522_n1170# sky130_fd_pr__pfet_01v8 ad=0.16665 pd=1.34 as=0.16665 ps=1.34 w=1.01 l=2.63
X5 VDD2.t8 VN.t1 VTAIL.t17 w_n4522_n1170# sky130_fd_pr__pfet_01v8 ad=0.16665 pd=1.34 as=0.3939 ps=2.8 w=1.01 l=2.63
X6 VTAIL.t14 VN.t2 VDD2.t7 w_n4522_n1170# sky130_fd_pr__pfet_01v8 ad=0.16665 pd=1.34 as=0.16665 ps=1.34 w=1.01 l=2.63
X7 VTAIL.t3 VN.t3 VDD2.t6 w_n4522_n1170# sky130_fd_pr__pfet_01v8 ad=0.16665 pd=1.34 as=0.16665 ps=1.34 w=1.01 l=2.63
X8 VTAIL.t12 VP.t3 VDD1.t6 w_n4522_n1170# sky130_fd_pr__pfet_01v8 ad=0.16665 pd=1.34 as=0.16665 ps=1.34 w=1.01 l=2.63
X9 B.t8 B.t6 B.t7 w_n4522_n1170# sky130_fd_pr__pfet_01v8 ad=0.3939 pd=2.8 as=0 ps=0 w=1.01 l=2.63
X10 VDD1.t5 VP.t4 VTAIL.t6 w_n4522_n1170# sky130_fd_pr__pfet_01v8 ad=0.3939 pd=2.8 as=0.16665 ps=1.34 w=1.01 l=2.63
X11 VDD2.t5 VN.t4 VTAIL.t2 w_n4522_n1170# sky130_fd_pr__pfet_01v8 ad=0.16665 pd=1.34 as=0.3939 ps=2.8 w=1.01 l=2.63
X12 VTAIL.t7 VP.t5 VDD1.t4 w_n4522_n1170# sky130_fd_pr__pfet_01v8 ad=0.16665 pd=1.34 as=0.16665 ps=1.34 w=1.01 l=2.63
X13 VTAIL.t18 VN.t5 VDD2.t4 w_n4522_n1170# sky130_fd_pr__pfet_01v8 ad=0.16665 pd=1.34 as=0.16665 ps=1.34 w=1.01 l=2.63
X14 VDD2.t3 VN.t6 VTAIL.t16 w_n4522_n1170# sky130_fd_pr__pfet_01v8 ad=0.3939 pd=2.8 as=0.16665 ps=1.34 w=1.01 l=2.63
X15 B.t5 B.t3 B.t4 w_n4522_n1170# sky130_fd_pr__pfet_01v8 ad=0.3939 pd=2.8 as=0 ps=0 w=1.01 l=2.63
X16 VDD1.t3 VP.t6 VTAIL.t10 w_n4522_n1170# sky130_fd_pr__pfet_01v8 ad=0.16665 pd=1.34 as=0.16665 ps=1.34 w=1.01 l=2.63
X17 VDD2.t2 VN.t7 VTAIL.t15 w_n4522_n1170# sky130_fd_pr__pfet_01v8 ad=0.16665 pd=1.34 as=0.16665 ps=1.34 w=1.01 l=2.63
X18 VDD2.t1 VN.t8 VTAIL.t0 w_n4522_n1170# sky130_fd_pr__pfet_01v8 ad=0.3939 pd=2.8 as=0.16665 ps=1.34 w=1.01 l=2.63
X19 VDD1.t2 VP.t7 VTAIL.t13 w_n4522_n1170# sky130_fd_pr__pfet_01v8 ad=0.16665 pd=1.34 as=0.16665 ps=1.34 w=1.01 l=2.63
X20 B.t2 B.t0 B.t1 w_n4522_n1170# sky130_fd_pr__pfet_01v8 ad=0.3939 pd=2.8 as=0 ps=0 w=1.01 l=2.63
X21 VDD1.t1 VP.t8 VTAIL.t11 w_n4522_n1170# sky130_fd_pr__pfet_01v8 ad=0.3939 pd=2.8 as=0.16665 ps=1.34 w=1.01 l=2.63
X22 VTAIL.t1 VN.t9 VDD2.t0 w_n4522_n1170# sky130_fd_pr__pfet_01v8 ad=0.16665 pd=1.34 as=0.16665 ps=1.34 w=1.01 l=2.63
X23 VTAIL.t4 VP.t9 VDD1.t0 w_n4522_n1170# sky130_fd_pr__pfet_01v8 ad=0.16665 pd=1.34 as=0.16665 ps=1.34 w=1.01 l=2.63
R0 VP.n25 VP.n22 161.3
R1 VP.n27 VP.n26 161.3
R2 VP.n28 VP.n21 161.3
R3 VP.n30 VP.n29 161.3
R4 VP.n31 VP.n20 161.3
R5 VP.n33 VP.n32 161.3
R6 VP.n35 VP.n19 161.3
R7 VP.n37 VP.n36 161.3
R8 VP.n38 VP.n18 161.3
R9 VP.n40 VP.n39 161.3
R10 VP.n41 VP.n17 161.3
R11 VP.n43 VP.n42 161.3
R12 VP.n45 VP.n44 161.3
R13 VP.n46 VP.n15 161.3
R14 VP.n48 VP.n47 161.3
R15 VP.n49 VP.n14 161.3
R16 VP.n51 VP.n50 161.3
R17 VP.n52 VP.n13 161.3
R18 VP.n94 VP.n0 161.3
R19 VP.n93 VP.n92 161.3
R20 VP.n91 VP.n1 161.3
R21 VP.n90 VP.n89 161.3
R22 VP.n88 VP.n2 161.3
R23 VP.n87 VP.n86 161.3
R24 VP.n85 VP.n84 161.3
R25 VP.n83 VP.n4 161.3
R26 VP.n82 VP.n81 161.3
R27 VP.n80 VP.n5 161.3
R28 VP.n79 VP.n78 161.3
R29 VP.n77 VP.n6 161.3
R30 VP.n75 VP.n74 161.3
R31 VP.n73 VP.n7 161.3
R32 VP.n72 VP.n71 161.3
R33 VP.n70 VP.n8 161.3
R34 VP.n69 VP.n68 161.3
R35 VP.n67 VP.n9 161.3
R36 VP.n66 VP.n65 161.3
R37 VP.n63 VP.n10 161.3
R38 VP.n62 VP.n61 161.3
R39 VP.n60 VP.n11 161.3
R40 VP.n59 VP.n58 161.3
R41 VP.n57 VP.n12 161.3
R42 VP.n56 VP.n55 102.438
R43 VP.n96 VP.n95 102.438
R44 VP.n54 VP.n53 102.438
R45 VP.n24 VP.n23 62.0711
R46 VP.n62 VP.n11 56.5193
R47 VP.n71 VP.n70 56.5193
R48 VP.n82 VP.n5 56.5193
R49 VP.n89 VP.n1 56.5193
R50 VP.n47 VP.n14 56.5193
R51 VP.n40 VP.n18 56.5193
R52 VP.n29 VP.n28 56.5193
R53 VP.n55 VP.n54 44.9541
R54 VP.n24 VP.t4 42.3725
R55 VP.n58 VP.n57 24.4675
R56 VP.n58 VP.n11 24.4675
R57 VP.n63 VP.n62 24.4675
R58 VP.n65 VP.n63 24.4675
R59 VP.n69 VP.n9 24.4675
R60 VP.n70 VP.n69 24.4675
R61 VP.n71 VP.n7 24.4675
R62 VP.n75 VP.n7 24.4675
R63 VP.n78 VP.n77 24.4675
R64 VP.n78 VP.n5 24.4675
R65 VP.n83 VP.n82 24.4675
R66 VP.n84 VP.n83 24.4675
R67 VP.n88 VP.n87 24.4675
R68 VP.n89 VP.n88 24.4675
R69 VP.n93 VP.n1 24.4675
R70 VP.n94 VP.n93 24.4675
R71 VP.n51 VP.n14 24.4675
R72 VP.n52 VP.n51 24.4675
R73 VP.n41 VP.n40 24.4675
R74 VP.n42 VP.n41 24.4675
R75 VP.n46 VP.n45 24.4675
R76 VP.n47 VP.n46 24.4675
R77 VP.n29 VP.n20 24.4675
R78 VP.n33 VP.n20 24.4675
R79 VP.n36 VP.n35 24.4675
R80 VP.n36 VP.n18 24.4675
R81 VP.n27 VP.n22 24.4675
R82 VP.n28 VP.n27 24.4675
R83 VP.n65 VP.n64 14.1914
R84 VP.n87 VP.n3 14.1914
R85 VP.n45 VP.n16 14.1914
R86 VP.n76 VP.n75 12.234
R87 VP.n77 VP.n76 12.234
R88 VP.n34 VP.n33 12.234
R89 VP.n35 VP.n34 12.234
R90 VP.n64 VP.n9 10.2766
R91 VP.n84 VP.n3 10.2766
R92 VP.n42 VP.n16 10.2766
R93 VP.n23 VP.n22 10.2766
R94 VP.n56 VP.t8 9.25563
R95 VP.n64 VP.t9 9.25563
R96 VP.n76 VP.t6 9.25563
R97 VP.n3 VP.t3 9.25563
R98 VP.n95 VP.t0 9.25563
R99 VP.n53 VP.t1 9.25563
R100 VP.n16 VP.t5 9.25563
R101 VP.n34 VP.t7 9.25563
R102 VP.n23 VP.t2 9.25563
R103 VP.n57 VP.n56 8.31928
R104 VP.n95 VP.n94 8.31928
R105 VP.n53 VP.n52 8.31928
R106 VP.n25 VP.n24 6.95571
R107 VP.n54 VP.n13 0.278367
R108 VP.n55 VP.n12 0.278367
R109 VP.n96 VP.n0 0.278367
R110 VP.n26 VP.n25 0.189894
R111 VP.n26 VP.n21 0.189894
R112 VP.n30 VP.n21 0.189894
R113 VP.n31 VP.n30 0.189894
R114 VP.n32 VP.n31 0.189894
R115 VP.n32 VP.n19 0.189894
R116 VP.n37 VP.n19 0.189894
R117 VP.n38 VP.n37 0.189894
R118 VP.n39 VP.n38 0.189894
R119 VP.n39 VP.n17 0.189894
R120 VP.n43 VP.n17 0.189894
R121 VP.n44 VP.n43 0.189894
R122 VP.n44 VP.n15 0.189894
R123 VP.n48 VP.n15 0.189894
R124 VP.n49 VP.n48 0.189894
R125 VP.n50 VP.n49 0.189894
R126 VP.n50 VP.n13 0.189894
R127 VP.n59 VP.n12 0.189894
R128 VP.n60 VP.n59 0.189894
R129 VP.n61 VP.n60 0.189894
R130 VP.n61 VP.n10 0.189894
R131 VP.n66 VP.n10 0.189894
R132 VP.n67 VP.n66 0.189894
R133 VP.n68 VP.n67 0.189894
R134 VP.n68 VP.n8 0.189894
R135 VP.n72 VP.n8 0.189894
R136 VP.n73 VP.n72 0.189894
R137 VP.n74 VP.n73 0.189894
R138 VP.n74 VP.n6 0.189894
R139 VP.n79 VP.n6 0.189894
R140 VP.n80 VP.n79 0.189894
R141 VP.n81 VP.n80 0.189894
R142 VP.n81 VP.n4 0.189894
R143 VP.n85 VP.n4 0.189894
R144 VP.n86 VP.n85 0.189894
R145 VP.n86 VP.n2 0.189894
R146 VP.n90 VP.n2 0.189894
R147 VP.n91 VP.n90 0.189894
R148 VP.n92 VP.n91 0.189894
R149 VP.n92 VP.n0 0.189894
R150 VP VP.n96 0.153454
R151 VTAIL.n16 VTAIL.t8 655.832
R152 VTAIL.n11 VTAIL.t2 655.832
R153 VTAIL.n17 VTAIL.t17 655.831
R154 VTAIL.n2 VTAIL.t9 655.831
R155 VTAIL.n15 VTAIL.n14 623.649
R156 VTAIL.n13 VTAIL.n12 623.649
R157 VTAIL.n10 VTAIL.n9 623.649
R158 VTAIL.n8 VTAIL.n7 623.649
R159 VTAIL.n19 VTAIL.n18 623.646
R160 VTAIL.n1 VTAIL.n0 623.646
R161 VTAIL.n4 VTAIL.n3 623.646
R162 VTAIL.n6 VTAIL.n5 623.646
R163 VTAIL.n18 VTAIL.t15 32.1837
R164 VTAIL.n18 VTAIL.t18 32.1837
R165 VTAIL.n0 VTAIL.t0 32.1837
R166 VTAIL.n0 VTAIL.t14 32.1837
R167 VTAIL.n3 VTAIL.t10 32.1837
R168 VTAIL.n3 VTAIL.t12 32.1837
R169 VTAIL.n5 VTAIL.t11 32.1837
R170 VTAIL.n5 VTAIL.t4 32.1837
R171 VTAIL.n14 VTAIL.t13 32.1837
R172 VTAIL.n14 VTAIL.t7 32.1837
R173 VTAIL.n12 VTAIL.t6 32.1837
R174 VTAIL.n12 VTAIL.t5 32.1837
R175 VTAIL.n9 VTAIL.t19 32.1837
R176 VTAIL.n9 VTAIL.t3 32.1837
R177 VTAIL.n7 VTAIL.t16 32.1837
R178 VTAIL.n7 VTAIL.t1 32.1837
R179 VTAIL.n8 VTAIL.n6 18.341
R180 VTAIL.n17 VTAIL.n16 15.7893
R181 VTAIL.n10 VTAIL.n8 2.55222
R182 VTAIL.n11 VTAIL.n10 2.55222
R183 VTAIL.n15 VTAIL.n13 2.55222
R184 VTAIL.n16 VTAIL.n15 2.55222
R185 VTAIL.n6 VTAIL.n4 2.55222
R186 VTAIL.n4 VTAIL.n2 2.55222
R187 VTAIL.n19 VTAIL.n17 2.55222
R188 VTAIL VTAIL.n1 1.97248
R189 VTAIL.n13 VTAIL.n11 1.74619
R190 VTAIL.n2 VTAIL.n1 1.74619
R191 VTAIL VTAIL.n19 0.580241
R192 VDD1.n1 VDD1.t5 675.062
R193 VDD1.n3 VDD1.t1 675.061
R194 VDD1.n5 VDD1.n4 642.184
R195 VDD1.n7 VDD1.n6 640.327
R196 VDD1.n1 VDD1.n0 640.327
R197 VDD1.n3 VDD1.n2 640.326
R198 VDD1.n7 VDD1.n5 38.5656
R199 VDD1.n6 VDD1.t4 32.1837
R200 VDD1.n6 VDD1.t8 32.1837
R201 VDD1.n0 VDD1.t7 32.1837
R202 VDD1.n0 VDD1.t2 32.1837
R203 VDD1.n4 VDD1.t6 32.1837
R204 VDD1.n4 VDD1.t9 32.1837
R205 VDD1.n2 VDD1.t0 32.1837
R206 VDD1.n2 VDD1.t3 32.1837
R207 VDD1 VDD1.n7 1.8561
R208 VDD1 VDD1.n1 0.696621
R209 VDD1.n5 VDD1.n3 0.583085
R210 B.n258 B.t7 703.875
R211 B.n117 B.t1 703.875
R212 B.n45 B.t11 703.875
R213 B.n38 B.t5 703.875
R214 B.n259 B.t8 646.468
R215 B.n118 B.t2 646.468
R216 B.n46 B.t10 646.468
R217 B.n39 B.t4 646.468
R218 B.n291 B.n112 585
R219 B.n290 B.n289 585
R220 B.n288 B.n113 585
R221 B.n287 B.n286 585
R222 B.n285 B.n114 585
R223 B.n284 B.n283 585
R224 B.n282 B.n115 585
R225 B.n281 B.n280 585
R226 B.n279 B.n116 585
R227 B.n277 B.n276 585
R228 B.n275 B.n119 585
R229 B.n274 B.n273 585
R230 B.n272 B.n120 585
R231 B.n271 B.n270 585
R232 B.n269 B.n121 585
R233 B.n268 B.n267 585
R234 B.n266 B.n122 585
R235 B.n265 B.n264 585
R236 B.n263 B.n123 585
R237 B.n262 B.n261 585
R238 B.n257 B.n124 585
R239 B.n256 B.n255 585
R240 B.n254 B.n125 585
R241 B.n253 B.n252 585
R242 B.n251 B.n126 585
R243 B.n250 B.n249 585
R244 B.n248 B.n127 585
R245 B.n247 B.n246 585
R246 B.n293 B.n292 585
R247 B.n294 B.n111 585
R248 B.n296 B.n295 585
R249 B.n297 B.n110 585
R250 B.n299 B.n298 585
R251 B.n300 B.n109 585
R252 B.n302 B.n301 585
R253 B.n303 B.n108 585
R254 B.n305 B.n304 585
R255 B.n306 B.n107 585
R256 B.n308 B.n307 585
R257 B.n309 B.n106 585
R258 B.n311 B.n310 585
R259 B.n312 B.n105 585
R260 B.n314 B.n313 585
R261 B.n315 B.n104 585
R262 B.n317 B.n316 585
R263 B.n318 B.n103 585
R264 B.n320 B.n319 585
R265 B.n321 B.n102 585
R266 B.n323 B.n322 585
R267 B.n324 B.n101 585
R268 B.n326 B.n325 585
R269 B.n327 B.n100 585
R270 B.n329 B.n328 585
R271 B.n330 B.n99 585
R272 B.n332 B.n331 585
R273 B.n333 B.n98 585
R274 B.n335 B.n334 585
R275 B.n336 B.n97 585
R276 B.n338 B.n337 585
R277 B.n339 B.n96 585
R278 B.n341 B.n340 585
R279 B.n342 B.n95 585
R280 B.n344 B.n343 585
R281 B.n345 B.n94 585
R282 B.n347 B.n346 585
R283 B.n348 B.n93 585
R284 B.n350 B.n349 585
R285 B.n351 B.n92 585
R286 B.n353 B.n352 585
R287 B.n354 B.n91 585
R288 B.n356 B.n355 585
R289 B.n357 B.n90 585
R290 B.n359 B.n358 585
R291 B.n360 B.n89 585
R292 B.n362 B.n361 585
R293 B.n363 B.n88 585
R294 B.n365 B.n364 585
R295 B.n366 B.n87 585
R296 B.n368 B.n367 585
R297 B.n369 B.n86 585
R298 B.n371 B.n370 585
R299 B.n372 B.n85 585
R300 B.n374 B.n373 585
R301 B.n375 B.n84 585
R302 B.n377 B.n376 585
R303 B.n378 B.n83 585
R304 B.n380 B.n379 585
R305 B.n381 B.n82 585
R306 B.n383 B.n382 585
R307 B.n384 B.n81 585
R308 B.n386 B.n385 585
R309 B.n387 B.n80 585
R310 B.n389 B.n388 585
R311 B.n390 B.n79 585
R312 B.n392 B.n391 585
R313 B.n393 B.n78 585
R314 B.n395 B.n394 585
R315 B.n396 B.n77 585
R316 B.n398 B.n397 585
R317 B.n399 B.n76 585
R318 B.n401 B.n400 585
R319 B.n402 B.n75 585
R320 B.n404 B.n403 585
R321 B.n405 B.n74 585
R322 B.n407 B.n406 585
R323 B.n408 B.n73 585
R324 B.n410 B.n409 585
R325 B.n411 B.n72 585
R326 B.n413 B.n412 585
R327 B.n414 B.n71 585
R328 B.n416 B.n415 585
R329 B.n417 B.n70 585
R330 B.n419 B.n418 585
R331 B.n420 B.n69 585
R332 B.n422 B.n421 585
R333 B.n423 B.n68 585
R334 B.n425 B.n424 585
R335 B.n426 B.n67 585
R336 B.n428 B.n427 585
R337 B.n429 B.n66 585
R338 B.n431 B.n430 585
R339 B.n432 B.n65 585
R340 B.n434 B.n433 585
R341 B.n435 B.n64 585
R342 B.n437 B.n436 585
R343 B.n438 B.n63 585
R344 B.n440 B.n439 585
R345 B.n441 B.n62 585
R346 B.n443 B.n442 585
R347 B.n444 B.n61 585
R348 B.n446 B.n445 585
R349 B.n447 B.n60 585
R350 B.n449 B.n448 585
R351 B.n450 B.n59 585
R352 B.n452 B.n451 585
R353 B.n453 B.n58 585
R354 B.n455 B.n454 585
R355 B.n456 B.n57 585
R356 B.n458 B.n457 585
R357 B.n459 B.n56 585
R358 B.n461 B.n460 585
R359 B.n462 B.n55 585
R360 B.n464 B.n463 585
R361 B.n465 B.n54 585
R362 B.n467 B.n466 585
R363 B.n468 B.n53 585
R364 B.n470 B.n469 585
R365 B.n471 B.n52 585
R366 B.n473 B.n472 585
R367 B.n474 B.n51 585
R368 B.n517 B.n32 585
R369 B.n516 B.n515 585
R370 B.n514 B.n33 585
R371 B.n513 B.n512 585
R372 B.n511 B.n34 585
R373 B.n510 B.n509 585
R374 B.n508 B.n35 585
R375 B.n507 B.n506 585
R376 B.n505 B.n36 585
R377 B.n504 B.n503 585
R378 B.n502 B.n37 585
R379 B.n501 B.n500 585
R380 B.n499 B.n41 585
R381 B.n498 B.n497 585
R382 B.n496 B.n42 585
R383 B.n495 B.n494 585
R384 B.n493 B.n43 585
R385 B.n492 B.n491 585
R386 B.n490 B.n44 585
R387 B.n488 B.n487 585
R388 B.n486 B.n47 585
R389 B.n485 B.n484 585
R390 B.n483 B.n48 585
R391 B.n482 B.n481 585
R392 B.n480 B.n49 585
R393 B.n479 B.n478 585
R394 B.n477 B.n50 585
R395 B.n476 B.n475 585
R396 B.n519 B.n518 585
R397 B.n520 B.n31 585
R398 B.n522 B.n521 585
R399 B.n523 B.n30 585
R400 B.n525 B.n524 585
R401 B.n526 B.n29 585
R402 B.n528 B.n527 585
R403 B.n529 B.n28 585
R404 B.n531 B.n530 585
R405 B.n532 B.n27 585
R406 B.n534 B.n533 585
R407 B.n535 B.n26 585
R408 B.n537 B.n536 585
R409 B.n538 B.n25 585
R410 B.n540 B.n539 585
R411 B.n541 B.n24 585
R412 B.n543 B.n542 585
R413 B.n544 B.n23 585
R414 B.n546 B.n545 585
R415 B.n547 B.n22 585
R416 B.n549 B.n548 585
R417 B.n550 B.n21 585
R418 B.n552 B.n551 585
R419 B.n553 B.n20 585
R420 B.n555 B.n554 585
R421 B.n556 B.n19 585
R422 B.n558 B.n557 585
R423 B.n559 B.n18 585
R424 B.n561 B.n560 585
R425 B.n562 B.n17 585
R426 B.n564 B.n563 585
R427 B.n565 B.n16 585
R428 B.n567 B.n566 585
R429 B.n568 B.n15 585
R430 B.n570 B.n569 585
R431 B.n571 B.n14 585
R432 B.n573 B.n572 585
R433 B.n574 B.n13 585
R434 B.n576 B.n575 585
R435 B.n577 B.n12 585
R436 B.n579 B.n578 585
R437 B.n580 B.n11 585
R438 B.n582 B.n581 585
R439 B.n583 B.n10 585
R440 B.n585 B.n584 585
R441 B.n586 B.n9 585
R442 B.n588 B.n587 585
R443 B.n589 B.n8 585
R444 B.n591 B.n590 585
R445 B.n592 B.n7 585
R446 B.n594 B.n593 585
R447 B.n595 B.n6 585
R448 B.n597 B.n596 585
R449 B.n598 B.n5 585
R450 B.n600 B.n599 585
R451 B.n601 B.n4 585
R452 B.n603 B.n602 585
R453 B.n604 B.n3 585
R454 B.n606 B.n605 585
R455 B.n607 B.n0 585
R456 B.n2 B.n1 585
R457 B.n158 B.n157 585
R458 B.n160 B.n159 585
R459 B.n161 B.n156 585
R460 B.n163 B.n162 585
R461 B.n164 B.n155 585
R462 B.n166 B.n165 585
R463 B.n167 B.n154 585
R464 B.n169 B.n168 585
R465 B.n170 B.n153 585
R466 B.n172 B.n171 585
R467 B.n173 B.n152 585
R468 B.n175 B.n174 585
R469 B.n176 B.n151 585
R470 B.n178 B.n177 585
R471 B.n179 B.n150 585
R472 B.n181 B.n180 585
R473 B.n182 B.n149 585
R474 B.n184 B.n183 585
R475 B.n185 B.n148 585
R476 B.n187 B.n186 585
R477 B.n188 B.n147 585
R478 B.n190 B.n189 585
R479 B.n191 B.n146 585
R480 B.n193 B.n192 585
R481 B.n194 B.n145 585
R482 B.n196 B.n195 585
R483 B.n197 B.n144 585
R484 B.n199 B.n198 585
R485 B.n200 B.n143 585
R486 B.n202 B.n201 585
R487 B.n203 B.n142 585
R488 B.n205 B.n204 585
R489 B.n206 B.n141 585
R490 B.n208 B.n207 585
R491 B.n209 B.n140 585
R492 B.n211 B.n210 585
R493 B.n212 B.n139 585
R494 B.n214 B.n213 585
R495 B.n215 B.n138 585
R496 B.n217 B.n216 585
R497 B.n218 B.n137 585
R498 B.n220 B.n219 585
R499 B.n221 B.n136 585
R500 B.n223 B.n222 585
R501 B.n224 B.n135 585
R502 B.n226 B.n225 585
R503 B.n227 B.n134 585
R504 B.n229 B.n228 585
R505 B.n230 B.n133 585
R506 B.n232 B.n231 585
R507 B.n233 B.n132 585
R508 B.n235 B.n234 585
R509 B.n236 B.n131 585
R510 B.n238 B.n237 585
R511 B.n239 B.n130 585
R512 B.n241 B.n240 585
R513 B.n242 B.n129 585
R514 B.n244 B.n243 585
R515 B.n245 B.n128 585
R516 B.n247 B.n128 487.695
R517 B.n293 B.n112 487.695
R518 B.n475 B.n474 487.695
R519 B.n518 B.n517 487.695
R520 B.n609 B.n608 256.663
R521 B.n608 B.n607 235.042
R522 B.n608 B.n2 235.042
R523 B.n258 B.t6 208.966
R524 B.n117 B.t0 208.966
R525 B.n45 B.t9 208.966
R526 B.n38 B.t3 208.966
R527 B.n248 B.n247 163.367
R528 B.n249 B.n248 163.367
R529 B.n249 B.n126 163.367
R530 B.n253 B.n126 163.367
R531 B.n254 B.n253 163.367
R532 B.n255 B.n254 163.367
R533 B.n255 B.n124 163.367
R534 B.n262 B.n124 163.367
R535 B.n263 B.n262 163.367
R536 B.n264 B.n263 163.367
R537 B.n264 B.n122 163.367
R538 B.n268 B.n122 163.367
R539 B.n269 B.n268 163.367
R540 B.n270 B.n269 163.367
R541 B.n270 B.n120 163.367
R542 B.n274 B.n120 163.367
R543 B.n275 B.n274 163.367
R544 B.n276 B.n275 163.367
R545 B.n276 B.n116 163.367
R546 B.n281 B.n116 163.367
R547 B.n282 B.n281 163.367
R548 B.n283 B.n282 163.367
R549 B.n283 B.n114 163.367
R550 B.n287 B.n114 163.367
R551 B.n288 B.n287 163.367
R552 B.n289 B.n288 163.367
R553 B.n289 B.n112 163.367
R554 B.n474 B.n473 163.367
R555 B.n473 B.n52 163.367
R556 B.n469 B.n52 163.367
R557 B.n469 B.n468 163.367
R558 B.n468 B.n467 163.367
R559 B.n467 B.n54 163.367
R560 B.n463 B.n54 163.367
R561 B.n463 B.n462 163.367
R562 B.n462 B.n461 163.367
R563 B.n461 B.n56 163.367
R564 B.n457 B.n56 163.367
R565 B.n457 B.n456 163.367
R566 B.n456 B.n455 163.367
R567 B.n455 B.n58 163.367
R568 B.n451 B.n58 163.367
R569 B.n451 B.n450 163.367
R570 B.n450 B.n449 163.367
R571 B.n449 B.n60 163.367
R572 B.n445 B.n60 163.367
R573 B.n445 B.n444 163.367
R574 B.n444 B.n443 163.367
R575 B.n443 B.n62 163.367
R576 B.n439 B.n62 163.367
R577 B.n439 B.n438 163.367
R578 B.n438 B.n437 163.367
R579 B.n437 B.n64 163.367
R580 B.n433 B.n64 163.367
R581 B.n433 B.n432 163.367
R582 B.n432 B.n431 163.367
R583 B.n431 B.n66 163.367
R584 B.n427 B.n66 163.367
R585 B.n427 B.n426 163.367
R586 B.n426 B.n425 163.367
R587 B.n425 B.n68 163.367
R588 B.n421 B.n68 163.367
R589 B.n421 B.n420 163.367
R590 B.n420 B.n419 163.367
R591 B.n419 B.n70 163.367
R592 B.n415 B.n70 163.367
R593 B.n415 B.n414 163.367
R594 B.n414 B.n413 163.367
R595 B.n413 B.n72 163.367
R596 B.n409 B.n72 163.367
R597 B.n409 B.n408 163.367
R598 B.n408 B.n407 163.367
R599 B.n407 B.n74 163.367
R600 B.n403 B.n74 163.367
R601 B.n403 B.n402 163.367
R602 B.n402 B.n401 163.367
R603 B.n401 B.n76 163.367
R604 B.n397 B.n76 163.367
R605 B.n397 B.n396 163.367
R606 B.n396 B.n395 163.367
R607 B.n395 B.n78 163.367
R608 B.n391 B.n78 163.367
R609 B.n391 B.n390 163.367
R610 B.n390 B.n389 163.367
R611 B.n389 B.n80 163.367
R612 B.n385 B.n80 163.367
R613 B.n385 B.n384 163.367
R614 B.n384 B.n383 163.367
R615 B.n383 B.n82 163.367
R616 B.n379 B.n82 163.367
R617 B.n379 B.n378 163.367
R618 B.n378 B.n377 163.367
R619 B.n377 B.n84 163.367
R620 B.n373 B.n84 163.367
R621 B.n373 B.n372 163.367
R622 B.n372 B.n371 163.367
R623 B.n371 B.n86 163.367
R624 B.n367 B.n86 163.367
R625 B.n367 B.n366 163.367
R626 B.n366 B.n365 163.367
R627 B.n365 B.n88 163.367
R628 B.n361 B.n88 163.367
R629 B.n361 B.n360 163.367
R630 B.n360 B.n359 163.367
R631 B.n359 B.n90 163.367
R632 B.n355 B.n90 163.367
R633 B.n355 B.n354 163.367
R634 B.n354 B.n353 163.367
R635 B.n353 B.n92 163.367
R636 B.n349 B.n92 163.367
R637 B.n349 B.n348 163.367
R638 B.n348 B.n347 163.367
R639 B.n347 B.n94 163.367
R640 B.n343 B.n94 163.367
R641 B.n343 B.n342 163.367
R642 B.n342 B.n341 163.367
R643 B.n341 B.n96 163.367
R644 B.n337 B.n96 163.367
R645 B.n337 B.n336 163.367
R646 B.n336 B.n335 163.367
R647 B.n335 B.n98 163.367
R648 B.n331 B.n98 163.367
R649 B.n331 B.n330 163.367
R650 B.n330 B.n329 163.367
R651 B.n329 B.n100 163.367
R652 B.n325 B.n100 163.367
R653 B.n325 B.n324 163.367
R654 B.n324 B.n323 163.367
R655 B.n323 B.n102 163.367
R656 B.n319 B.n102 163.367
R657 B.n319 B.n318 163.367
R658 B.n318 B.n317 163.367
R659 B.n317 B.n104 163.367
R660 B.n313 B.n104 163.367
R661 B.n313 B.n312 163.367
R662 B.n312 B.n311 163.367
R663 B.n311 B.n106 163.367
R664 B.n307 B.n106 163.367
R665 B.n307 B.n306 163.367
R666 B.n306 B.n305 163.367
R667 B.n305 B.n108 163.367
R668 B.n301 B.n108 163.367
R669 B.n301 B.n300 163.367
R670 B.n300 B.n299 163.367
R671 B.n299 B.n110 163.367
R672 B.n295 B.n110 163.367
R673 B.n295 B.n294 163.367
R674 B.n294 B.n293 163.367
R675 B.n517 B.n516 163.367
R676 B.n516 B.n33 163.367
R677 B.n512 B.n33 163.367
R678 B.n512 B.n511 163.367
R679 B.n511 B.n510 163.367
R680 B.n510 B.n35 163.367
R681 B.n506 B.n35 163.367
R682 B.n506 B.n505 163.367
R683 B.n505 B.n504 163.367
R684 B.n504 B.n37 163.367
R685 B.n500 B.n37 163.367
R686 B.n500 B.n499 163.367
R687 B.n499 B.n498 163.367
R688 B.n498 B.n42 163.367
R689 B.n494 B.n42 163.367
R690 B.n494 B.n493 163.367
R691 B.n493 B.n492 163.367
R692 B.n492 B.n44 163.367
R693 B.n487 B.n44 163.367
R694 B.n487 B.n486 163.367
R695 B.n486 B.n485 163.367
R696 B.n485 B.n48 163.367
R697 B.n481 B.n48 163.367
R698 B.n481 B.n480 163.367
R699 B.n480 B.n479 163.367
R700 B.n479 B.n50 163.367
R701 B.n475 B.n50 163.367
R702 B.n518 B.n31 163.367
R703 B.n522 B.n31 163.367
R704 B.n523 B.n522 163.367
R705 B.n524 B.n523 163.367
R706 B.n524 B.n29 163.367
R707 B.n528 B.n29 163.367
R708 B.n529 B.n528 163.367
R709 B.n530 B.n529 163.367
R710 B.n530 B.n27 163.367
R711 B.n534 B.n27 163.367
R712 B.n535 B.n534 163.367
R713 B.n536 B.n535 163.367
R714 B.n536 B.n25 163.367
R715 B.n540 B.n25 163.367
R716 B.n541 B.n540 163.367
R717 B.n542 B.n541 163.367
R718 B.n542 B.n23 163.367
R719 B.n546 B.n23 163.367
R720 B.n547 B.n546 163.367
R721 B.n548 B.n547 163.367
R722 B.n548 B.n21 163.367
R723 B.n552 B.n21 163.367
R724 B.n553 B.n552 163.367
R725 B.n554 B.n553 163.367
R726 B.n554 B.n19 163.367
R727 B.n558 B.n19 163.367
R728 B.n559 B.n558 163.367
R729 B.n560 B.n559 163.367
R730 B.n560 B.n17 163.367
R731 B.n564 B.n17 163.367
R732 B.n565 B.n564 163.367
R733 B.n566 B.n565 163.367
R734 B.n566 B.n15 163.367
R735 B.n570 B.n15 163.367
R736 B.n571 B.n570 163.367
R737 B.n572 B.n571 163.367
R738 B.n572 B.n13 163.367
R739 B.n576 B.n13 163.367
R740 B.n577 B.n576 163.367
R741 B.n578 B.n577 163.367
R742 B.n578 B.n11 163.367
R743 B.n582 B.n11 163.367
R744 B.n583 B.n582 163.367
R745 B.n584 B.n583 163.367
R746 B.n584 B.n9 163.367
R747 B.n588 B.n9 163.367
R748 B.n589 B.n588 163.367
R749 B.n590 B.n589 163.367
R750 B.n590 B.n7 163.367
R751 B.n594 B.n7 163.367
R752 B.n595 B.n594 163.367
R753 B.n596 B.n595 163.367
R754 B.n596 B.n5 163.367
R755 B.n600 B.n5 163.367
R756 B.n601 B.n600 163.367
R757 B.n602 B.n601 163.367
R758 B.n602 B.n3 163.367
R759 B.n606 B.n3 163.367
R760 B.n607 B.n606 163.367
R761 B.n158 B.n2 163.367
R762 B.n159 B.n158 163.367
R763 B.n159 B.n156 163.367
R764 B.n163 B.n156 163.367
R765 B.n164 B.n163 163.367
R766 B.n165 B.n164 163.367
R767 B.n165 B.n154 163.367
R768 B.n169 B.n154 163.367
R769 B.n170 B.n169 163.367
R770 B.n171 B.n170 163.367
R771 B.n171 B.n152 163.367
R772 B.n175 B.n152 163.367
R773 B.n176 B.n175 163.367
R774 B.n177 B.n176 163.367
R775 B.n177 B.n150 163.367
R776 B.n181 B.n150 163.367
R777 B.n182 B.n181 163.367
R778 B.n183 B.n182 163.367
R779 B.n183 B.n148 163.367
R780 B.n187 B.n148 163.367
R781 B.n188 B.n187 163.367
R782 B.n189 B.n188 163.367
R783 B.n189 B.n146 163.367
R784 B.n193 B.n146 163.367
R785 B.n194 B.n193 163.367
R786 B.n195 B.n194 163.367
R787 B.n195 B.n144 163.367
R788 B.n199 B.n144 163.367
R789 B.n200 B.n199 163.367
R790 B.n201 B.n200 163.367
R791 B.n201 B.n142 163.367
R792 B.n205 B.n142 163.367
R793 B.n206 B.n205 163.367
R794 B.n207 B.n206 163.367
R795 B.n207 B.n140 163.367
R796 B.n211 B.n140 163.367
R797 B.n212 B.n211 163.367
R798 B.n213 B.n212 163.367
R799 B.n213 B.n138 163.367
R800 B.n217 B.n138 163.367
R801 B.n218 B.n217 163.367
R802 B.n219 B.n218 163.367
R803 B.n219 B.n136 163.367
R804 B.n223 B.n136 163.367
R805 B.n224 B.n223 163.367
R806 B.n225 B.n224 163.367
R807 B.n225 B.n134 163.367
R808 B.n229 B.n134 163.367
R809 B.n230 B.n229 163.367
R810 B.n231 B.n230 163.367
R811 B.n231 B.n132 163.367
R812 B.n235 B.n132 163.367
R813 B.n236 B.n235 163.367
R814 B.n237 B.n236 163.367
R815 B.n237 B.n130 163.367
R816 B.n241 B.n130 163.367
R817 B.n242 B.n241 163.367
R818 B.n243 B.n242 163.367
R819 B.n243 B.n128 163.367
R820 B.n260 B.n259 59.5399
R821 B.n278 B.n118 59.5399
R822 B.n489 B.n46 59.5399
R823 B.n40 B.n39 59.5399
R824 B.n259 B.n258 57.4066
R825 B.n118 B.n117 57.4066
R826 B.n46 B.n45 57.4066
R827 B.n39 B.n38 57.4066
R828 B.n519 B.n32 31.6883
R829 B.n476 B.n51 31.6883
R830 B.n292 B.n291 31.6883
R831 B.n246 B.n245 31.6883
R832 B B.n609 18.0485
R833 B.n520 B.n519 10.6151
R834 B.n521 B.n520 10.6151
R835 B.n521 B.n30 10.6151
R836 B.n525 B.n30 10.6151
R837 B.n526 B.n525 10.6151
R838 B.n527 B.n526 10.6151
R839 B.n527 B.n28 10.6151
R840 B.n531 B.n28 10.6151
R841 B.n532 B.n531 10.6151
R842 B.n533 B.n532 10.6151
R843 B.n533 B.n26 10.6151
R844 B.n537 B.n26 10.6151
R845 B.n538 B.n537 10.6151
R846 B.n539 B.n538 10.6151
R847 B.n539 B.n24 10.6151
R848 B.n543 B.n24 10.6151
R849 B.n544 B.n543 10.6151
R850 B.n545 B.n544 10.6151
R851 B.n545 B.n22 10.6151
R852 B.n549 B.n22 10.6151
R853 B.n550 B.n549 10.6151
R854 B.n551 B.n550 10.6151
R855 B.n551 B.n20 10.6151
R856 B.n555 B.n20 10.6151
R857 B.n556 B.n555 10.6151
R858 B.n557 B.n556 10.6151
R859 B.n557 B.n18 10.6151
R860 B.n561 B.n18 10.6151
R861 B.n562 B.n561 10.6151
R862 B.n563 B.n562 10.6151
R863 B.n563 B.n16 10.6151
R864 B.n567 B.n16 10.6151
R865 B.n568 B.n567 10.6151
R866 B.n569 B.n568 10.6151
R867 B.n569 B.n14 10.6151
R868 B.n573 B.n14 10.6151
R869 B.n574 B.n573 10.6151
R870 B.n575 B.n574 10.6151
R871 B.n575 B.n12 10.6151
R872 B.n579 B.n12 10.6151
R873 B.n580 B.n579 10.6151
R874 B.n581 B.n580 10.6151
R875 B.n581 B.n10 10.6151
R876 B.n585 B.n10 10.6151
R877 B.n586 B.n585 10.6151
R878 B.n587 B.n586 10.6151
R879 B.n587 B.n8 10.6151
R880 B.n591 B.n8 10.6151
R881 B.n592 B.n591 10.6151
R882 B.n593 B.n592 10.6151
R883 B.n593 B.n6 10.6151
R884 B.n597 B.n6 10.6151
R885 B.n598 B.n597 10.6151
R886 B.n599 B.n598 10.6151
R887 B.n599 B.n4 10.6151
R888 B.n603 B.n4 10.6151
R889 B.n604 B.n603 10.6151
R890 B.n605 B.n604 10.6151
R891 B.n605 B.n0 10.6151
R892 B.n515 B.n32 10.6151
R893 B.n515 B.n514 10.6151
R894 B.n514 B.n513 10.6151
R895 B.n513 B.n34 10.6151
R896 B.n509 B.n34 10.6151
R897 B.n509 B.n508 10.6151
R898 B.n508 B.n507 10.6151
R899 B.n507 B.n36 10.6151
R900 B.n503 B.n502 10.6151
R901 B.n502 B.n501 10.6151
R902 B.n501 B.n41 10.6151
R903 B.n497 B.n41 10.6151
R904 B.n497 B.n496 10.6151
R905 B.n496 B.n495 10.6151
R906 B.n495 B.n43 10.6151
R907 B.n491 B.n43 10.6151
R908 B.n491 B.n490 10.6151
R909 B.n488 B.n47 10.6151
R910 B.n484 B.n47 10.6151
R911 B.n484 B.n483 10.6151
R912 B.n483 B.n482 10.6151
R913 B.n482 B.n49 10.6151
R914 B.n478 B.n49 10.6151
R915 B.n478 B.n477 10.6151
R916 B.n477 B.n476 10.6151
R917 B.n472 B.n51 10.6151
R918 B.n472 B.n471 10.6151
R919 B.n471 B.n470 10.6151
R920 B.n470 B.n53 10.6151
R921 B.n466 B.n53 10.6151
R922 B.n466 B.n465 10.6151
R923 B.n465 B.n464 10.6151
R924 B.n464 B.n55 10.6151
R925 B.n460 B.n55 10.6151
R926 B.n460 B.n459 10.6151
R927 B.n459 B.n458 10.6151
R928 B.n458 B.n57 10.6151
R929 B.n454 B.n57 10.6151
R930 B.n454 B.n453 10.6151
R931 B.n453 B.n452 10.6151
R932 B.n452 B.n59 10.6151
R933 B.n448 B.n59 10.6151
R934 B.n448 B.n447 10.6151
R935 B.n447 B.n446 10.6151
R936 B.n446 B.n61 10.6151
R937 B.n442 B.n61 10.6151
R938 B.n442 B.n441 10.6151
R939 B.n441 B.n440 10.6151
R940 B.n440 B.n63 10.6151
R941 B.n436 B.n63 10.6151
R942 B.n436 B.n435 10.6151
R943 B.n435 B.n434 10.6151
R944 B.n434 B.n65 10.6151
R945 B.n430 B.n65 10.6151
R946 B.n430 B.n429 10.6151
R947 B.n429 B.n428 10.6151
R948 B.n428 B.n67 10.6151
R949 B.n424 B.n67 10.6151
R950 B.n424 B.n423 10.6151
R951 B.n423 B.n422 10.6151
R952 B.n422 B.n69 10.6151
R953 B.n418 B.n69 10.6151
R954 B.n418 B.n417 10.6151
R955 B.n417 B.n416 10.6151
R956 B.n416 B.n71 10.6151
R957 B.n412 B.n71 10.6151
R958 B.n412 B.n411 10.6151
R959 B.n411 B.n410 10.6151
R960 B.n410 B.n73 10.6151
R961 B.n406 B.n73 10.6151
R962 B.n406 B.n405 10.6151
R963 B.n405 B.n404 10.6151
R964 B.n404 B.n75 10.6151
R965 B.n400 B.n75 10.6151
R966 B.n400 B.n399 10.6151
R967 B.n399 B.n398 10.6151
R968 B.n398 B.n77 10.6151
R969 B.n394 B.n77 10.6151
R970 B.n394 B.n393 10.6151
R971 B.n393 B.n392 10.6151
R972 B.n392 B.n79 10.6151
R973 B.n388 B.n79 10.6151
R974 B.n388 B.n387 10.6151
R975 B.n387 B.n386 10.6151
R976 B.n386 B.n81 10.6151
R977 B.n382 B.n81 10.6151
R978 B.n382 B.n381 10.6151
R979 B.n381 B.n380 10.6151
R980 B.n380 B.n83 10.6151
R981 B.n376 B.n83 10.6151
R982 B.n376 B.n375 10.6151
R983 B.n375 B.n374 10.6151
R984 B.n374 B.n85 10.6151
R985 B.n370 B.n85 10.6151
R986 B.n370 B.n369 10.6151
R987 B.n369 B.n368 10.6151
R988 B.n368 B.n87 10.6151
R989 B.n364 B.n87 10.6151
R990 B.n364 B.n363 10.6151
R991 B.n363 B.n362 10.6151
R992 B.n362 B.n89 10.6151
R993 B.n358 B.n89 10.6151
R994 B.n358 B.n357 10.6151
R995 B.n357 B.n356 10.6151
R996 B.n356 B.n91 10.6151
R997 B.n352 B.n91 10.6151
R998 B.n352 B.n351 10.6151
R999 B.n351 B.n350 10.6151
R1000 B.n350 B.n93 10.6151
R1001 B.n346 B.n93 10.6151
R1002 B.n346 B.n345 10.6151
R1003 B.n345 B.n344 10.6151
R1004 B.n344 B.n95 10.6151
R1005 B.n340 B.n95 10.6151
R1006 B.n340 B.n339 10.6151
R1007 B.n339 B.n338 10.6151
R1008 B.n338 B.n97 10.6151
R1009 B.n334 B.n97 10.6151
R1010 B.n334 B.n333 10.6151
R1011 B.n333 B.n332 10.6151
R1012 B.n332 B.n99 10.6151
R1013 B.n328 B.n99 10.6151
R1014 B.n328 B.n327 10.6151
R1015 B.n327 B.n326 10.6151
R1016 B.n326 B.n101 10.6151
R1017 B.n322 B.n101 10.6151
R1018 B.n322 B.n321 10.6151
R1019 B.n321 B.n320 10.6151
R1020 B.n320 B.n103 10.6151
R1021 B.n316 B.n103 10.6151
R1022 B.n316 B.n315 10.6151
R1023 B.n315 B.n314 10.6151
R1024 B.n314 B.n105 10.6151
R1025 B.n310 B.n105 10.6151
R1026 B.n310 B.n309 10.6151
R1027 B.n309 B.n308 10.6151
R1028 B.n308 B.n107 10.6151
R1029 B.n304 B.n107 10.6151
R1030 B.n304 B.n303 10.6151
R1031 B.n303 B.n302 10.6151
R1032 B.n302 B.n109 10.6151
R1033 B.n298 B.n109 10.6151
R1034 B.n298 B.n297 10.6151
R1035 B.n297 B.n296 10.6151
R1036 B.n296 B.n111 10.6151
R1037 B.n292 B.n111 10.6151
R1038 B.n157 B.n1 10.6151
R1039 B.n160 B.n157 10.6151
R1040 B.n161 B.n160 10.6151
R1041 B.n162 B.n161 10.6151
R1042 B.n162 B.n155 10.6151
R1043 B.n166 B.n155 10.6151
R1044 B.n167 B.n166 10.6151
R1045 B.n168 B.n167 10.6151
R1046 B.n168 B.n153 10.6151
R1047 B.n172 B.n153 10.6151
R1048 B.n173 B.n172 10.6151
R1049 B.n174 B.n173 10.6151
R1050 B.n174 B.n151 10.6151
R1051 B.n178 B.n151 10.6151
R1052 B.n179 B.n178 10.6151
R1053 B.n180 B.n179 10.6151
R1054 B.n180 B.n149 10.6151
R1055 B.n184 B.n149 10.6151
R1056 B.n185 B.n184 10.6151
R1057 B.n186 B.n185 10.6151
R1058 B.n186 B.n147 10.6151
R1059 B.n190 B.n147 10.6151
R1060 B.n191 B.n190 10.6151
R1061 B.n192 B.n191 10.6151
R1062 B.n192 B.n145 10.6151
R1063 B.n196 B.n145 10.6151
R1064 B.n197 B.n196 10.6151
R1065 B.n198 B.n197 10.6151
R1066 B.n198 B.n143 10.6151
R1067 B.n202 B.n143 10.6151
R1068 B.n203 B.n202 10.6151
R1069 B.n204 B.n203 10.6151
R1070 B.n204 B.n141 10.6151
R1071 B.n208 B.n141 10.6151
R1072 B.n209 B.n208 10.6151
R1073 B.n210 B.n209 10.6151
R1074 B.n210 B.n139 10.6151
R1075 B.n214 B.n139 10.6151
R1076 B.n215 B.n214 10.6151
R1077 B.n216 B.n215 10.6151
R1078 B.n216 B.n137 10.6151
R1079 B.n220 B.n137 10.6151
R1080 B.n221 B.n220 10.6151
R1081 B.n222 B.n221 10.6151
R1082 B.n222 B.n135 10.6151
R1083 B.n226 B.n135 10.6151
R1084 B.n227 B.n226 10.6151
R1085 B.n228 B.n227 10.6151
R1086 B.n228 B.n133 10.6151
R1087 B.n232 B.n133 10.6151
R1088 B.n233 B.n232 10.6151
R1089 B.n234 B.n233 10.6151
R1090 B.n234 B.n131 10.6151
R1091 B.n238 B.n131 10.6151
R1092 B.n239 B.n238 10.6151
R1093 B.n240 B.n239 10.6151
R1094 B.n240 B.n129 10.6151
R1095 B.n244 B.n129 10.6151
R1096 B.n245 B.n244 10.6151
R1097 B.n246 B.n127 10.6151
R1098 B.n250 B.n127 10.6151
R1099 B.n251 B.n250 10.6151
R1100 B.n252 B.n251 10.6151
R1101 B.n252 B.n125 10.6151
R1102 B.n256 B.n125 10.6151
R1103 B.n257 B.n256 10.6151
R1104 B.n261 B.n257 10.6151
R1105 B.n265 B.n123 10.6151
R1106 B.n266 B.n265 10.6151
R1107 B.n267 B.n266 10.6151
R1108 B.n267 B.n121 10.6151
R1109 B.n271 B.n121 10.6151
R1110 B.n272 B.n271 10.6151
R1111 B.n273 B.n272 10.6151
R1112 B.n273 B.n119 10.6151
R1113 B.n277 B.n119 10.6151
R1114 B.n280 B.n279 10.6151
R1115 B.n280 B.n115 10.6151
R1116 B.n284 B.n115 10.6151
R1117 B.n285 B.n284 10.6151
R1118 B.n286 B.n285 10.6151
R1119 B.n286 B.n113 10.6151
R1120 B.n290 B.n113 10.6151
R1121 B.n291 B.n290 10.6151
R1122 B.n40 B.n36 9.36635
R1123 B.n489 B.n488 9.36635
R1124 B.n261 B.n260 9.36635
R1125 B.n279 B.n278 9.36635
R1126 B.n609 B.n0 8.11757
R1127 B.n609 B.n1 8.11757
R1128 B.n503 B.n40 1.24928
R1129 B.n490 B.n489 1.24928
R1130 B.n260 B.n123 1.24928
R1131 B.n278 B.n277 1.24928
R1132 VN.n81 VN.n42 161.3
R1133 VN.n80 VN.n79 161.3
R1134 VN.n78 VN.n43 161.3
R1135 VN.n77 VN.n76 161.3
R1136 VN.n75 VN.n44 161.3
R1137 VN.n74 VN.n73 161.3
R1138 VN.n72 VN.n71 161.3
R1139 VN.n70 VN.n46 161.3
R1140 VN.n69 VN.n68 161.3
R1141 VN.n67 VN.n47 161.3
R1142 VN.n66 VN.n65 161.3
R1143 VN.n64 VN.n48 161.3
R1144 VN.n62 VN.n61 161.3
R1145 VN.n60 VN.n49 161.3
R1146 VN.n59 VN.n58 161.3
R1147 VN.n57 VN.n50 161.3
R1148 VN.n56 VN.n55 161.3
R1149 VN.n54 VN.n51 161.3
R1150 VN.n39 VN.n0 161.3
R1151 VN.n38 VN.n37 161.3
R1152 VN.n36 VN.n1 161.3
R1153 VN.n35 VN.n34 161.3
R1154 VN.n33 VN.n2 161.3
R1155 VN.n32 VN.n31 161.3
R1156 VN.n30 VN.n29 161.3
R1157 VN.n28 VN.n4 161.3
R1158 VN.n27 VN.n26 161.3
R1159 VN.n25 VN.n5 161.3
R1160 VN.n24 VN.n23 161.3
R1161 VN.n22 VN.n6 161.3
R1162 VN.n20 VN.n19 161.3
R1163 VN.n18 VN.n7 161.3
R1164 VN.n17 VN.n16 161.3
R1165 VN.n15 VN.n8 161.3
R1166 VN.n14 VN.n13 161.3
R1167 VN.n12 VN.n9 161.3
R1168 VN.n41 VN.n40 102.438
R1169 VN.n83 VN.n82 102.438
R1170 VN.n11 VN.n10 62.0711
R1171 VN.n53 VN.n52 62.0711
R1172 VN.n16 VN.n15 56.5193
R1173 VN.n27 VN.n5 56.5193
R1174 VN.n34 VN.n1 56.5193
R1175 VN.n58 VN.n57 56.5193
R1176 VN.n69 VN.n47 56.5193
R1177 VN.n76 VN.n43 56.5193
R1178 VN VN.n83 45.233
R1179 VN.n11 VN.t8 42.3725
R1180 VN.n53 VN.t4 42.3725
R1181 VN.n14 VN.n9 24.4675
R1182 VN.n15 VN.n14 24.4675
R1183 VN.n16 VN.n7 24.4675
R1184 VN.n20 VN.n7 24.4675
R1185 VN.n23 VN.n22 24.4675
R1186 VN.n23 VN.n5 24.4675
R1187 VN.n28 VN.n27 24.4675
R1188 VN.n29 VN.n28 24.4675
R1189 VN.n33 VN.n32 24.4675
R1190 VN.n34 VN.n33 24.4675
R1191 VN.n38 VN.n1 24.4675
R1192 VN.n39 VN.n38 24.4675
R1193 VN.n57 VN.n56 24.4675
R1194 VN.n56 VN.n51 24.4675
R1195 VN.n65 VN.n47 24.4675
R1196 VN.n65 VN.n64 24.4675
R1197 VN.n62 VN.n49 24.4675
R1198 VN.n58 VN.n49 24.4675
R1199 VN.n76 VN.n75 24.4675
R1200 VN.n75 VN.n74 24.4675
R1201 VN.n71 VN.n70 24.4675
R1202 VN.n70 VN.n69 24.4675
R1203 VN.n81 VN.n80 24.4675
R1204 VN.n80 VN.n43 24.4675
R1205 VN.n32 VN.n3 14.1914
R1206 VN.n74 VN.n45 14.1914
R1207 VN.n21 VN.n20 12.234
R1208 VN.n22 VN.n21 12.234
R1209 VN.n64 VN.n63 12.234
R1210 VN.n63 VN.n62 12.234
R1211 VN.n10 VN.n9 10.2766
R1212 VN.n29 VN.n3 10.2766
R1213 VN.n52 VN.n51 10.2766
R1214 VN.n71 VN.n45 10.2766
R1215 VN.n10 VN.t2 9.25563
R1216 VN.n21 VN.t7 9.25563
R1217 VN.n3 VN.t5 9.25563
R1218 VN.n40 VN.t1 9.25563
R1219 VN.n52 VN.t3 9.25563
R1220 VN.n63 VN.t0 9.25563
R1221 VN.n45 VN.t9 9.25563
R1222 VN.n82 VN.t6 9.25563
R1223 VN.n40 VN.n39 8.31928
R1224 VN.n82 VN.n81 8.31928
R1225 VN.n54 VN.n53 6.95571
R1226 VN.n12 VN.n11 6.95571
R1227 VN.n83 VN.n42 0.278367
R1228 VN.n41 VN.n0 0.278367
R1229 VN.n79 VN.n42 0.189894
R1230 VN.n79 VN.n78 0.189894
R1231 VN.n78 VN.n77 0.189894
R1232 VN.n77 VN.n44 0.189894
R1233 VN.n73 VN.n44 0.189894
R1234 VN.n73 VN.n72 0.189894
R1235 VN.n72 VN.n46 0.189894
R1236 VN.n68 VN.n46 0.189894
R1237 VN.n68 VN.n67 0.189894
R1238 VN.n67 VN.n66 0.189894
R1239 VN.n66 VN.n48 0.189894
R1240 VN.n61 VN.n48 0.189894
R1241 VN.n61 VN.n60 0.189894
R1242 VN.n60 VN.n59 0.189894
R1243 VN.n59 VN.n50 0.189894
R1244 VN.n55 VN.n50 0.189894
R1245 VN.n55 VN.n54 0.189894
R1246 VN.n13 VN.n12 0.189894
R1247 VN.n13 VN.n8 0.189894
R1248 VN.n17 VN.n8 0.189894
R1249 VN.n18 VN.n17 0.189894
R1250 VN.n19 VN.n18 0.189894
R1251 VN.n19 VN.n6 0.189894
R1252 VN.n24 VN.n6 0.189894
R1253 VN.n25 VN.n24 0.189894
R1254 VN.n26 VN.n25 0.189894
R1255 VN.n26 VN.n4 0.189894
R1256 VN.n30 VN.n4 0.189894
R1257 VN.n31 VN.n30 0.189894
R1258 VN.n31 VN.n2 0.189894
R1259 VN.n35 VN.n2 0.189894
R1260 VN.n36 VN.n35 0.189894
R1261 VN.n37 VN.n36 0.189894
R1262 VN.n37 VN.n0 0.189894
R1263 VN VN.n41 0.153454
R1264 VDD2.n1 VDD2.t1 675.061
R1265 VDD2.n4 VDD2.t3 672.51
R1266 VDD2.n3 VDD2.n2 642.184
R1267 VDD2 VDD2.n7 642.183
R1268 VDD2.n6 VDD2.n5 640.327
R1269 VDD2.n1 VDD2.n0 640.326
R1270 VDD2.n4 VDD2.n3 36.7067
R1271 VDD2.n7 VDD2.t6 32.1837
R1272 VDD2.n7 VDD2.t5 32.1837
R1273 VDD2.n5 VDD2.t0 32.1837
R1274 VDD2.n5 VDD2.t9 32.1837
R1275 VDD2.n2 VDD2.t4 32.1837
R1276 VDD2.n2 VDD2.t8 32.1837
R1277 VDD2.n0 VDD2.t7 32.1837
R1278 VDD2.n0 VDD2.t2 32.1837
R1279 VDD2.n6 VDD2.n4 2.55222
R1280 VDD2 VDD2.n6 0.696621
R1281 VDD2.n3 VDD2.n1 0.583085
C0 VN VDD1 0.161519f
C1 VTAIL VP 2.9833f
C2 B w_n4522_n1170# 7.60509f
C3 VN VTAIL 2.96918f
C4 VDD1 VTAIL 5.35501f
C5 VDD2 VP 0.596787f
C6 VN VDD2 1.37811f
C7 VDD1 VDD2 2.19384f
C8 VTAIL VDD2 5.40871f
C9 w_n4522_n1170# VP 10.100201f
C10 B VP 2.13235f
C11 VN w_n4522_n1170# 9.51905f
C12 VDD1 w_n4522_n1170# 2.03044f
C13 VN B 1.14326f
C14 VDD1 B 1.62187f
C15 VTAIL w_n4522_n1170# 1.61288f
C16 VTAIL B 1.11336f
C17 VDD2 w_n4522_n1170# 2.17448f
C18 B VDD2 1.74158f
C19 VN VP 6.41625f
C20 VDD1 VP 1.80865f
C21 VDD2 VSUBS 1.686894f
C22 VDD1 VSUBS 1.66871f
C23 VTAIL VSUBS 0.564526f
C24 VN VSUBS 8.05424f
C25 VP VSUBS 3.588434f
C26 B VSUBS 4.191217f
C27 w_n4522_n1170# VSUBS 68.20979f
C28 VDD2.t1 VSUBS 0.144816f
C29 VDD2.t7 VSUBS 0.027311f
C30 VDD2.t2 VSUBS 0.027311f
C31 VDD2.n0 VSUBS 0.073959f
C32 VDD2.n1 VSUBS 1.19166f
C33 VDD2.t4 VSUBS 0.027311f
C34 VDD2.t8 VSUBS 0.027311f
C35 VDD2.n2 VSUBS 0.076198f
C36 VDD2.n3 VSUBS 3.10833f
C37 VDD2.t3 VSUBS 0.142646f
C38 VDD2.n4 VSUBS 3.01084f
C39 VDD2.t0 VSUBS 0.027311f
C40 VDD2.t9 VSUBS 0.027311f
C41 VDD2.n5 VSUBS 0.073959f
C42 VDD2.n6 VSUBS 0.631082f
C43 VDD2.t6 VSUBS 0.027311f
C44 VDD2.t5 VSUBS 0.027311f
C45 VDD2.n7 VSUBS 0.076192f
C46 VN.n0 VSUBS 0.076811f
C47 VN.t1 VSUBS 0.290568f
C48 VN.n1 VSUBS 0.094791f
C49 VN.n2 VSUBS 0.058261f
C50 VN.t5 VSUBS 0.290568f
C51 VN.n3 VSUBS 0.198177f
C52 VN.n4 VSUBS 0.058261f
C53 VN.n5 VSUBS 0.081803f
C54 VN.n6 VSUBS 0.058261f
C55 VN.t7 VSUBS 0.290568f
C56 VN.n7 VSUBS 0.108583f
C57 VN.n8 VSUBS 0.058261f
C58 VN.n9 VSUBS 0.077491f
C59 VN.t8 VSUBS 0.728712f
C60 VN.t2 VSUBS 0.290568f
C61 VN.n10 VSUBS 0.362952f
C62 VN.n11 VSUBS 0.36747f
C63 VN.n12 VSUBS 0.564886f
C64 VN.n13 VSUBS 0.058261f
C65 VN.n14 VSUBS 0.108583f
C66 VN.n15 VSUBS 0.088297f
C67 VN.n16 VSUBS 0.081803f
C68 VN.n17 VSUBS 0.058261f
C69 VN.n18 VSUBS 0.058261f
C70 VN.n19 VSUBS 0.058261f
C71 VN.n20 VSUBS 0.081779f
C72 VN.n21 VSUBS 0.198177f
C73 VN.n22 VSUBS 0.081779f
C74 VN.n23 VSUBS 0.108583f
C75 VN.n24 VSUBS 0.058261f
C76 VN.n25 VSUBS 0.058261f
C77 VN.n26 VSUBS 0.058261f
C78 VN.n27 VSUBS 0.088297f
C79 VN.n28 VSUBS 0.108583f
C80 VN.n29 VSUBS 0.077491f
C81 VN.n30 VSUBS 0.058261f
C82 VN.n31 VSUBS 0.058261f
C83 VN.n32 VSUBS 0.086068f
C84 VN.n33 VSUBS 0.108583f
C85 VN.n34 VSUBS 0.075309f
C86 VN.n35 VSUBS 0.058261f
C87 VN.n36 VSUBS 0.058261f
C88 VN.n37 VSUBS 0.058261f
C89 VN.n38 VSUBS 0.108583f
C90 VN.n39 VSUBS 0.073202f
C91 VN.n40 VSUBS 0.390566f
C92 VN.n41 VSUBS 0.09781f
C93 VN.n42 VSUBS 0.076811f
C94 VN.t6 VSUBS 0.290568f
C95 VN.n43 VSUBS 0.094791f
C96 VN.n44 VSUBS 0.058261f
C97 VN.t9 VSUBS 0.290568f
C98 VN.n45 VSUBS 0.198177f
C99 VN.n46 VSUBS 0.058261f
C100 VN.n47 VSUBS 0.081803f
C101 VN.n48 VSUBS 0.058261f
C102 VN.t0 VSUBS 0.290568f
C103 VN.n49 VSUBS 0.108583f
C104 VN.n50 VSUBS 0.058261f
C105 VN.n51 VSUBS 0.077491f
C106 VN.t4 VSUBS 0.728712f
C107 VN.t3 VSUBS 0.290568f
C108 VN.n52 VSUBS 0.362952f
C109 VN.n53 VSUBS 0.36747f
C110 VN.n54 VSUBS 0.564886f
C111 VN.n55 VSUBS 0.058261f
C112 VN.n56 VSUBS 0.108583f
C113 VN.n57 VSUBS 0.088297f
C114 VN.n58 VSUBS 0.081803f
C115 VN.n59 VSUBS 0.058261f
C116 VN.n60 VSUBS 0.058261f
C117 VN.n61 VSUBS 0.058261f
C118 VN.n62 VSUBS 0.081779f
C119 VN.n63 VSUBS 0.198177f
C120 VN.n64 VSUBS 0.081779f
C121 VN.n65 VSUBS 0.108583f
C122 VN.n66 VSUBS 0.058261f
C123 VN.n67 VSUBS 0.058261f
C124 VN.n68 VSUBS 0.058261f
C125 VN.n69 VSUBS 0.088297f
C126 VN.n70 VSUBS 0.108583f
C127 VN.n71 VSUBS 0.077491f
C128 VN.n72 VSUBS 0.058261f
C129 VN.n73 VSUBS 0.058261f
C130 VN.n74 VSUBS 0.086068f
C131 VN.n75 VSUBS 0.108583f
C132 VN.n76 VSUBS 0.075309f
C133 VN.n77 VSUBS 0.058261f
C134 VN.n78 VSUBS 0.058261f
C135 VN.n79 VSUBS 0.058261f
C136 VN.n80 VSUBS 0.108583f
C137 VN.n81 VSUBS 0.073202f
C138 VN.n82 VSUBS 0.390566f
C139 VN.n83 VSUBS 2.79581f
C140 B.n0 VSUBS 0.010801f
C141 B.n1 VSUBS 0.010801f
C142 B.n2 VSUBS 0.015973f
C143 B.n3 VSUBS 0.012241f
C144 B.n4 VSUBS 0.012241f
C145 B.n5 VSUBS 0.012241f
C146 B.n6 VSUBS 0.012241f
C147 B.n7 VSUBS 0.012241f
C148 B.n8 VSUBS 0.012241f
C149 B.n9 VSUBS 0.012241f
C150 B.n10 VSUBS 0.012241f
C151 B.n11 VSUBS 0.012241f
C152 B.n12 VSUBS 0.012241f
C153 B.n13 VSUBS 0.012241f
C154 B.n14 VSUBS 0.012241f
C155 B.n15 VSUBS 0.012241f
C156 B.n16 VSUBS 0.012241f
C157 B.n17 VSUBS 0.012241f
C158 B.n18 VSUBS 0.012241f
C159 B.n19 VSUBS 0.012241f
C160 B.n20 VSUBS 0.012241f
C161 B.n21 VSUBS 0.012241f
C162 B.n22 VSUBS 0.012241f
C163 B.n23 VSUBS 0.012241f
C164 B.n24 VSUBS 0.012241f
C165 B.n25 VSUBS 0.012241f
C166 B.n26 VSUBS 0.012241f
C167 B.n27 VSUBS 0.012241f
C168 B.n28 VSUBS 0.012241f
C169 B.n29 VSUBS 0.012241f
C170 B.n30 VSUBS 0.012241f
C171 B.n31 VSUBS 0.012241f
C172 B.n32 VSUBS 0.0285f
C173 B.n33 VSUBS 0.012241f
C174 B.n34 VSUBS 0.012241f
C175 B.n35 VSUBS 0.012241f
C176 B.n36 VSUBS 0.011521f
C177 B.n37 VSUBS 0.012241f
C178 B.t4 VSUBS 0.034389f
C179 B.t5 VSUBS 0.039522f
C180 B.t3 VSUBS 0.23559f
C181 B.n38 VSUBS 0.107911f
C182 B.n39 VSUBS 0.080394f
C183 B.n40 VSUBS 0.02836f
C184 B.n41 VSUBS 0.012241f
C185 B.n42 VSUBS 0.012241f
C186 B.n43 VSUBS 0.012241f
C187 B.n44 VSUBS 0.012241f
C188 B.t10 VSUBS 0.034389f
C189 B.t11 VSUBS 0.039522f
C190 B.t9 VSUBS 0.23559f
C191 B.n45 VSUBS 0.107911f
C192 B.n46 VSUBS 0.080394f
C193 B.n47 VSUBS 0.012241f
C194 B.n48 VSUBS 0.012241f
C195 B.n49 VSUBS 0.012241f
C196 B.n50 VSUBS 0.012241f
C197 B.n51 VSUBS 0.027664f
C198 B.n52 VSUBS 0.012241f
C199 B.n53 VSUBS 0.012241f
C200 B.n54 VSUBS 0.012241f
C201 B.n55 VSUBS 0.012241f
C202 B.n56 VSUBS 0.012241f
C203 B.n57 VSUBS 0.012241f
C204 B.n58 VSUBS 0.012241f
C205 B.n59 VSUBS 0.012241f
C206 B.n60 VSUBS 0.012241f
C207 B.n61 VSUBS 0.012241f
C208 B.n62 VSUBS 0.012241f
C209 B.n63 VSUBS 0.012241f
C210 B.n64 VSUBS 0.012241f
C211 B.n65 VSUBS 0.012241f
C212 B.n66 VSUBS 0.012241f
C213 B.n67 VSUBS 0.012241f
C214 B.n68 VSUBS 0.012241f
C215 B.n69 VSUBS 0.012241f
C216 B.n70 VSUBS 0.012241f
C217 B.n71 VSUBS 0.012241f
C218 B.n72 VSUBS 0.012241f
C219 B.n73 VSUBS 0.012241f
C220 B.n74 VSUBS 0.012241f
C221 B.n75 VSUBS 0.012241f
C222 B.n76 VSUBS 0.012241f
C223 B.n77 VSUBS 0.012241f
C224 B.n78 VSUBS 0.012241f
C225 B.n79 VSUBS 0.012241f
C226 B.n80 VSUBS 0.012241f
C227 B.n81 VSUBS 0.012241f
C228 B.n82 VSUBS 0.012241f
C229 B.n83 VSUBS 0.012241f
C230 B.n84 VSUBS 0.012241f
C231 B.n85 VSUBS 0.012241f
C232 B.n86 VSUBS 0.012241f
C233 B.n87 VSUBS 0.012241f
C234 B.n88 VSUBS 0.012241f
C235 B.n89 VSUBS 0.012241f
C236 B.n90 VSUBS 0.012241f
C237 B.n91 VSUBS 0.012241f
C238 B.n92 VSUBS 0.012241f
C239 B.n93 VSUBS 0.012241f
C240 B.n94 VSUBS 0.012241f
C241 B.n95 VSUBS 0.012241f
C242 B.n96 VSUBS 0.012241f
C243 B.n97 VSUBS 0.012241f
C244 B.n98 VSUBS 0.012241f
C245 B.n99 VSUBS 0.012241f
C246 B.n100 VSUBS 0.012241f
C247 B.n101 VSUBS 0.012241f
C248 B.n102 VSUBS 0.012241f
C249 B.n103 VSUBS 0.012241f
C250 B.n104 VSUBS 0.012241f
C251 B.n105 VSUBS 0.012241f
C252 B.n106 VSUBS 0.012241f
C253 B.n107 VSUBS 0.012241f
C254 B.n108 VSUBS 0.012241f
C255 B.n109 VSUBS 0.012241f
C256 B.n110 VSUBS 0.012241f
C257 B.n111 VSUBS 0.012241f
C258 B.n112 VSUBS 0.0285f
C259 B.n113 VSUBS 0.012241f
C260 B.n114 VSUBS 0.012241f
C261 B.n115 VSUBS 0.012241f
C262 B.n116 VSUBS 0.012241f
C263 B.t2 VSUBS 0.034389f
C264 B.t1 VSUBS 0.039522f
C265 B.t0 VSUBS 0.23559f
C266 B.n117 VSUBS 0.107911f
C267 B.n118 VSUBS 0.080394f
C268 B.n119 VSUBS 0.012241f
C269 B.n120 VSUBS 0.012241f
C270 B.n121 VSUBS 0.012241f
C271 B.n122 VSUBS 0.012241f
C272 B.n123 VSUBS 0.00684f
C273 B.n124 VSUBS 0.012241f
C274 B.n125 VSUBS 0.012241f
C275 B.n126 VSUBS 0.012241f
C276 B.n127 VSUBS 0.012241f
C277 B.n128 VSUBS 0.027664f
C278 B.n129 VSUBS 0.012241f
C279 B.n130 VSUBS 0.012241f
C280 B.n131 VSUBS 0.012241f
C281 B.n132 VSUBS 0.012241f
C282 B.n133 VSUBS 0.012241f
C283 B.n134 VSUBS 0.012241f
C284 B.n135 VSUBS 0.012241f
C285 B.n136 VSUBS 0.012241f
C286 B.n137 VSUBS 0.012241f
C287 B.n138 VSUBS 0.012241f
C288 B.n139 VSUBS 0.012241f
C289 B.n140 VSUBS 0.012241f
C290 B.n141 VSUBS 0.012241f
C291 B.n142 VSUBS 0.012241f
C292 B.n143 VSUBS 0.012241f
C293 B.n144 VSUBS 0.012241f
C294 B.n145 VSUBS 0.012241f
C295 B.n146 VSUBS 0.012241f
C296 B.n147 VSUBS 0.012241f
C297 B.n148 VSUBS 0.012241f
C298 B.n149 VSUBS 0.012241f
C299 B.n150 VSUBS 0.012241f
C300 B.n151 VSUBS 0.012241f
C301 B.n152 VSUBS 0.012241f
C302 B.n153 VSUBS 0.012241f
C303 B.n154 VSUBS 0.012241f
C304 B.n155 VSUBS 0.012241f
C305 B.n156 VSUBS 0.012241f
C306 B.n157 VSUBS 0.012241f
C307 B.n158 VSUBS 0.012241f
C308 B.n159 VSUBS 0.012241f
C309 B.n160 VSUBS 0.012241f
C310 B.n161 VSUBS 0.012241f
C311 B.n162 VSUBS 0.012241f
C312 B.n163 VSUBS 0.012241f
C313 B.n164 VSUBS 0.012241f
C314 B.n165 VSUBS 0.012241f
C315 B.n166 VSUBS 0.012241f
C316 B.n167 VSUBS 0.012241f
C317 B.n168 VSUBS 0.012241f
C318 B.n169 VSUBS 0.012241f
C319 B.n170 VSUBS 0.012241f
C320 B.n171 VSUBS 0.012241f
C321 B.n172 VSUBS 0.012241f
C322 B.n173 VSUBS 0.012241f
C323 B.n174 VSUBS 0.012241f
C324 B.n175 VSUBS 0.012241f
C325 B.n176 VSUBS 0.012241f
C326 B.n177 VSUBS 0.012241f
C327 B.n178 VSUBS 0.012241f
C328 B.n179 VSUBS 0.012241f
C329 B.n180 VSUBS 0.012241f
C330 B.n181 VSUBS 0.012241f
C331 B.n182 VSUBS 0.012241f
C332 B.n183 VSUBS 0.012241f
C333 B.n184 VSUBS 0.012241f
C334 B.n185 VSUBS 0.012241f
C335 B.n186 VSUBS 0.012241f
C336 B.n187 VSUBS 0.012241f
C337 B.n188 VSUBS 0.012241f
C338 B.n189 VSUBS 0.012241f
C339 B.n190 VSUBS 0.012241f
C340 B.n191 VSUBS 0.012241f
C341 B.n192 VSUBS 0.012241f
C342 B.n193 VSUBS 0.012241f
C343 B.n194 VSUBS 0.012241f
C344 B.n195 VSUBS 0.012241f
C345 B.n196 VSUBS 0.012241f
C346 B.n197 VSUBS 0.012241f
C347 B.n198 VSUBS 0.012241f
C348 B.n199 VSUBS 0.012241f
C349 B.n200 VSUBS 0.012241f
C350 B.n201 VSUBS 0.012241f
C351 B.n202 VSUBS 0.012241f
C352 B.n203 VSUBS 0.012241f
C353 B.n204 VSUBS 0.012241f
C354 B.n205 VSUBS 0.012241f
C355 B.n206 VSUBS 0.012241f
C356 B.n207 VSUBS 0.012241f
C357 B.n208 VSUBS 0.012241f
C358 B.n209 VSUBS 0.012241f
C359 B.n210 VSUBS 0.012241f
C360 B.n211 VSUBS 0.012241f
C361 B.n212 VSUBS 0.012241f
C362 B.n213 VSUBS 0.012241f
C363 B.n214 VSUBS 0.012241f
C364 B.n215 VSUBS 0.012241f
C365 B.n216 VSUBS 0.012241f
C366 B.n217 VSUBS 0.012241f
C367 B.n218 VSUBS 0.012241f
C368 B.n219 VSUBS 0.012241f
C369 B.n220 VSUBS 0.012241f
C370 B.n221 VSUBS 0.012241f
C371 B.n222 VSUBS 0.012241f
C372 B.n223 VSUBS 0.012241f
C373 B.n224 VSUBS 0.012241f
C374 B.n225 VSUBS 0.012241f
C375 B.n226 VSUBS 0.012241f
C376 B.n227 VSUBS 0.012241f
C377 B.n228 VSUBS 0.012241f
C378 B.n229 VSUBS 0.012241f
C379 B.n230 VSUBS 0.012241f
C380 B.n231 VSUBS 0.012241f
C381 B.n232 VSUBS 0.012241f
C382 B.n233 VSUBS 0.012241f
C383 B.n234 VSUBS 0.012241f
C384 B.n235 VSUBS 0.012241f
C385 B.n236 VSUBS 0.012241f
C386 B.n237 VSUBS 0.012241f
C387 B.n238 VSUBS 0.012241f
C388 B.n239 VSUBS 0.012241f
C389 B.n240 VSUBS 0.012241f
C390 B.n241 VSUBS 0.012241f
C391 B.n242 VSUBS 0.012241f
C392 B.n243 VSUBS 0.012241f
C393 B.n244 VSUBS 0.012241f
C394 B.n245 VSUBS 0.027664f
C395 B.n246 VSUBS 0.0285f
C396 B.n247 VSUBS 0.0285f
C397 B.n248 VSUBS 0.012241f
C398 B.n249 VSUBS 0.012241f
C399 B.n250 VSUBS 0.012241f
C400 B.n251 VSUBS 0.012241f
C401 B.n252 VSUBS 0.012241f
C402 B.n253 VSUBS 0.012241f
C403 B.n254 VSUBS 0.012241f
C404 B.n255 VSUBS 0.012241f
C405 B.n256 VSUBS 0.012241f
C406 B.n257 VSUBS 0.012241f
C407 B.t8 VSUBS 0.034389f
C408 B.t7 VSUBS 0.039522f
C409 B.t6 VSUBS 0.23559f
C410 B.n258 VSUBS 0.107911f
C411 B.n259 VSUBS 0.080394f
C412 B.n260 VSUBS 0.02836f
C413 B.n261 VSUBS 0.011521f
C414 B.n262 VSUBS 0.012241f
C415 B.n263 VSUBS 0.012241f
C416 B.n264 VSUBS 0.012241f
C417 B.n265 VSUBS 0.012241f
C418 B.n266 VSUBS 0.012241f
C419 B.n267 VSUBS 0.012241f
C420 B.n268 VSUBS 0.012241f
C421 B.n269 VSUBS 0.012241f
C422 B.n270 VSUBS 0.012241f
C423 B.n271 VSUBS 0.012241f
C424 B.n272 VSUBS 0.012241f
C425 B.n273 VSUBS 0.012241f
C426 B.n274 VSUBS 0.012241f
C427 B.n275 VSUBS 0.012241f
C428 B.n276 VSUBS 0.012241f
C429 B.n277 VSUBS 0.00684f
C430 B.n278 VSUBS 0.02836f
C431 B.n279 VSUBS 0.011521f
C432 B.n280 VSUBS 0.012241f
C433 B.n281 VSUBS 0.012241f
C434 B.n282 VSUBS 0.012241f
C435 B.n283 VSUBS 0.012241f
C436 B.n284 VSUBS 0.012241f
C437 B.n285 VSUBS 0.012241f
C438 B.n286 VSUBS 0.012241f
C439 B.n287 VSUBS 0.012241f
C440 B.n288 VSUBS 0.012241f
C441 B.n289 VSUBS 0.012241f
C442 B.n290 VSUBS 0.012241f
C443 B.n291 VSUBS 0.027009f
C444 B.n292 VSUBS 0.029154f
C445 B.n293 VSUBS 0.027664f
C446 B.n294 VSUBS 0.012241f
C447 B.n295 VSUBS 0.012241f
C448 B.n296 VSUBS 0.012241f
C449 B.n297 VSUBS 0.012241f
C450 B.n298 VSUBS 0.012241f
C451 B.n299 VSUBS 0.012241f
C452 B.n300 VSUBS 0.012241f
C453 B.n301 VSUBS 0.012241f
C454 B.n302 VSUBS 0.012241f
C455 B.n303 VSUBS 0.012241f
C456 B.n304 VSUBS 0.012241f
C457 B.n305 VSUBS 0.012241f
C458 B.n306 VSUBS 0.012241f
C459 B.n307 VSUBS 0.012241f
C460 B.n308 VSUBS 0.012241f
C461 B.n309 VSUBS 0.012241f
C462 B.n310 VSUBS 0.012241f
C463 B.n311 VSUBS 0.012241f
C464 B.n312 VSUBS 0.012241f
C465 B.n313 VSUBS 0.012241f
C466 B.n314 VSUBS 0.012241f
C467 B.n315 VSUBS 0.012241f
C468 B.n316 VSUBS 0.012241f
C469 B.n317 VSUBS 0.012241f
C470 B.n318 VSUBS 0.012241f
C471 B.n319 VSUBS 0.012241f
C472 B.n320 VSUBS 0.012241f
C473 B.n321 VSUBS 0.012241f
C474 B.n322 VSUBS 0.012241f
C475 B.n323 VSUBS 0.012241f
C476 B.n324 VSUBS 0.012241f
C477 B.n325 VSUBS 0.012241f
C478 B.n326 VSUBS 0.012241f
C479 B.n327 VSUBS 0.012241f
C480 B.n328 VSUBS 0.012241f
C481 B.n329 VSUBS 0.012241f
C482 B.n330 VSUBS 0.012241f
C483 B.n331 VSUBS 0.012241f
C484 B.n332 VSUBS 0.012241f
C485 B.n333 VSUBS 0.012241f
C486 B.n334 VSUBS 0.012241f
C487 B.n335 VSUBS 0.012241f
C488 B.n336 VSUBS 0.012241f
C489 B.n337 VSUBS 0.012241f
C490 B.n338 VSUBS 0.012241f
C491 B.n339 VSUBS 0.012241f
C492 B.n340 VSUBS 0.012241f
C493 B.n341 VSUBS 0.012241f
C494 B.n342 VSUBS 0.012241f
C495 B.n343 VSUBS 0.012241f
C496 B.n344 VSUBS 0.012241f
C497 B.n345 VSUBS 0.012241f
C498 B.n346 VSUBS 0.012241f
C499 B.n347 VSUBS 0.012241f
C500 B.n348 VSUBS 0.012241f
C501 B.n349 VSUBS 0.012241f
C502 B.n350 VSUBS 0.012241f
C503 B.n351 VSUBS 0.012241f
C504 B.n352 VSUBS 0.012241f
C505 B.n353 VSUBS 0.012241f
C506 B.n354 VSUBS 0.012241f
C507 B.n355 VSUBS 0.012241f
C508 B.n356 VSUBS 0.012241f
C509 B.n357 VSUBS 0.012241f
C510 B.n358 VSUBS 0.012241f
C511 B.n359 VSUBS 0.012241f
C512 B.n360 VSUBS 0.012241f
C513 B.n361 VSUBS 0.012241f
C514 B.n362 VSUBS 0.012241f
C515 B.n363 VSUBS 0.012241f
C516 B.n364 VSUBS 0.012241f
C517 B.n365 VSUBS 0.012241f
C518 B.n366 VSUBS 0.012241f
C519 B.n367 VSUBS 0.012241f
C520 B.n368 VSUBS 0.012241f
C521 B.n369 VSUBS 0.012241f
C522 B.n370 VSUBS 0.012241f
C523 B.n371 VSUBS 0.012241f
C524 B.n372 VSUBS 0.012241f
C525 B.n373 VSUBS 0.012241f
C526 B.n374 VSUBS 0.012241f
C527 B.n375 VSUBS 0.012241f
C528 B.n376 VSUBS 0.012241f
C529 B.n377 VSUBS 0.012241f
C530 B.n378 VSUBS 0.012241f
C531 B.n379 VSUBS 0.012241f
C532 B.n380 VSUBS 0.012241f
C533 B.n381 VSUBS 0.012241f
C534 B.n382 VSUBS 0.012241f
C535 B.n383 VSUBS 0.012241f
C536 B.n384 VSUBS 0.012241f
C537 B.n385 VSUBS 0.012241f
C538 B.n386 VSUBS 0.012241f
C539 B.n387 VSUBS 0.012241f
C540 B.n388 VSUBS 0.012241f
C541 B.n389 VSUBS 0.012241f
C542 B.n390 VSUBS 0.012241f
C543 B.n391 VSUBS 0.012241f
C544 B.n392 VSUBS 0.012241f
C545 B.n393 VSUBS 0.012241f
C546 B.n394 VSUBS 0.012241f
C547 B.n395 VSUBS 0.012241f
C548 B.n396 VSUBS 0.012241f
C549 B.n397 VSUBS 0.012241f
C550 B.n398 VSUBS 0.012241f
C551 B.n399 VSUBS 0.012241f
C552 B.n400 VSUBS 0.012241f
C553 B.n401 VSUBS 0.012241f
C554 B.n402 VSUBS 0.012241f
C555 B.n403 VSUBS 0.012241f
C556 B.n404 VSUBS 0.012241f
C557 B.n405 VSUBS 0.012241f
C558 B.n406 VSUBS 0.012241f
C559 B.n407 VSUBS 0.012241f
C560 B.n408 VSUBS 0.012241f
C561 B.n409 VSUBS 0.012241f
C562 B.n410 VSUBS 0.012241f
C563 B.n411 VSUBS 0.012241f
C564 B.n412 VSUBS 0.012241f
C565 B.n413 VSUBS 0.012241f
C566 B.n414 VSUBS 0.012241f
C567 B.n415 VSUBS 0.012241f
C568 B.n416 VSUBS 0.012241f
C569 B.n417 VSUBS 0.012241f
C570 B.n418 VSUBS 0.012241f
C571 B.n419 VSUBS 0.012241f
C572 B.n420 VSUBS 0.012241f
C573 B.n421 VSUBS 0.012241f
C574 B.n422 VSUBS 0.012241f
C575 B.n423 VSUBS 0.012241f
C576 B.n424 VSUBS 0.012241f
C577 B.n425 VSUBS 0.012241f
C578 B.n426 VSUBS 0.012241f
C579 B.n427 VSUBS 0.012241f
C580 B.n428 VSUBS 0.012241f
C581 B.n429 VSUBS 0.012241f
C582 B.n430 VSUBS 0.012241f
C583 B.n431 VSUBS 0.012241f
C584 B.n432 VSUBS 0.012241f
C585 B.n433 VSUBS 0.012241f
C586 B.n434 VSUBS 0.012241f
C587 B.n435 VSUBS 0.012241f
C588 B.n436 VSUBS 0.012241f
C589 B.n437 VSUBS 0.012241f
C590 B.n438 VSUBS 0.012241f
C591 B.n439 VSUBS 0.012241f
C592 B.n440 VSUBS 0.012241f
C593 B.n441 VSUBS 0.012241f
C594 B.n442 VSUBS 0.012241f
C595 B.n443 VSUBS 0.012241f
C596 B.n444 VSUBS 0.012241f
C597 B.n445 VSUBS 0.012241f
C598 B.n446 VSUBS 0.012241f
C599 B.n447 VSUBS 0.012241f
C600 B.n448 VSUBS 0.012241f
C601 B.n449 VSUBS 0.012241f
C602 B.n450 VSUBS 0.012241f
C603 B.n451 VSUBS 0.012241f
C604 B.n452 VSUBS 0.012241f
C605 B.n453 VSUBS 0.012241f
C606 B.n454 VSUBS 0.012241f
C607 B.n455 VSUBS 0.012241f
C608 B.n456 VSUBS 0.012241f
C609 B.n457 VSUBS 0.012241f
C610 B.n458 VSUBS 0.012241f
C611 B.n459 VSUBS 0.012241f
C612 B.n460 VSUBS 0.012241f
C613 B.n461 VSUBS 0.012241f
C614 B.n462 VSUBS 0.012241f
C615 B.n463 VSUBS 0.012241f
C616 B.n464 VSUBS 0.012241f
C617 B.n465 VSUBS 0.012241f
C618 B.n466 VSUBS 0.012241f
C619 B.n467 VSUBS 0.012241f
C620 B.n468 VSUBS 0.012241f
C621 B.n469 VSUBS 0.012241f
C622 B.n470 VSUBS 0.012241f
C623 B.n471 VSUBS 0.012241f
C624 B.n472 VSUBS 0.012241f
C625 B.n473 VSUBS 0.012241f
C626 B.n474 VSUBS 0.027664f
C627 B.n475 VSUBS 0.0285f
C628 B.n476 VSUBS 0.0285f
C629 B.n477 VSUBS 0.012241f
C630 B.n478 VSUBS 0.012241f
C631 B.n479 VSUBS 0.012241f
C632 B.n480 VSUBS 0.012241f
C633 B.n481 VSUBS 0.012241f
C634 B.n482 VSUBS 0.012241f
C635 B.n483 VSUBS 0.012241f
C636 B.n484 VSUBS 0.012241f
C637 B.n485 VSUBS 0.012241f
C638 B.n486 VSUBS 0.012241f
C639 B.n487 VSUBS 0.012241f
C640 B.n488 VSUBS 0.011521f
C641 B.n489 VSUBS 0.02836f
C642 B.n490 VSUBS 0.00684f
C643 B.n491 VSUBS 0.012241f
C644 B.n492 VSUBS 0.012241f
C645 B.n493 VSUBS 0.012241f
C646 B.n494 VSUBS 0.012241f
C647 B.n495 VSUBS 0.012241f
C648 B.n496 VSUBS 0.012241f
C649 B.n497 VSUBS 0.012241f
C650 B.n498 VSUBS 0.012241f
C651 B.n499 VSUBS 0.012241f
C652 B.n500 VSUBS 0.012241f
C653 B.n501 VSUBS 0.012241f
C654 B.n502 VSUBS 0.012241f
C655 B.n503 VSUBS 0.00684f
C656 B.n504 VSUBS 0.012241f
C657 B.n505 VSUBS 0.012241f
C658 B.n506 VSUBS 0.012241f
C659 B.n507 VSUBS 0.012241f
C660 B.n508 VSUBS 0.012241f
C661 B.n509 VSUBS 0.012241f
C662 B.n510 VSUBS 0.012241f
C663 B.n511 VSUBS 0.012241f
C664 B.n512 VSUBS 0.012241f
C665 B.n513 VSUBS 0.012241f
C666 B.n514 VSUBS 0.012241f
C667 B.n515 VSUBS 0.012241f
C668 B.n516 VSUBS 0.012241f
C669 B.n517 VSUBS 0.0285f
C670 B.n518 VSUBS 0.027664f
C671 B.n519 VSUBS 0.027664f
C672 B.n520 VSUBS 0.012241f
C673 B.n521 VSUBS 0.012241f
C674 B.n522 VSUBS 0.012241f
C675 B.n523 VSUBS 0.012241f
C676 B.n524 VSUBS 0.012241f
C677 B.n525 VSUBS 0.012241f
C678 B.n526 VSUBS 0.012241f
C679 B.n527 VSUBS 0.012241f
C680 B.n528 VSUBS 0.012241f
C681 B.n529 VSUBS 0.012241f
C682 B.n530 VSUBS 0.012241f
C683 B.n531 VSUBS 0.012241f
C684 B.n532 VSUBS 0.012241f
C685 B.n533 VSUBS 0.012241f
C686 B.n534 VSUBS 0.012241f
C687 B.n535 VSUBS 0.012241f
C688 B.n536 VSUBS 0.012241f
C689 B.n537 VSUBS 0.012241f
C690 B.n538 VSUBS 0.012241f
C691 B.n539 VSUBS 0.012241f
C692 B.n540 VSUBS 0.012241f
C693 B.n541 VSUBS 0.012241f
C694 B.n542 VSUBS 0.012241f
C695 B.n543 VSUBS 0.012241f
C696 B.n544 VSUBS 0.012241f
C697 B.n545 VSUBS 0.012241f
C698 B.n546 VSUBS 0.012241f
C699 B.n547 VSUBS 0.012241f
C700 B.n548 VSUBS 0.012241f
C701 B.n549 VSUBS 0.012241f
C702 B.n550 VSUBS 0.012241f
C703 B.n551 VSUBS 0.012241f
C704 B.n552 VSUBS 0.012241f
C705 B.n553 VSUBS 0.012241f
C706 B.n554 VSUBS 0.012241f
C707 B.n555 VSUBS 0.012241f
C708 B.n556 VSUBS 0.012241f
C709 B.n557 VSUBS 0.012241f
C710 B.n558 VSUBS 0.012241f
C711 B.n559 VSUBS 0.012241f
C712 B.n560 VSUBS 0.012241f
C713 B.n561 VSUBS 0.012241f
C714 B.n562 VSUBS 0.012241f
C715 B.n563 VSUBS 0.012241f
C716 B.n564 VSUBS 0.012241f
C717 B.n565 VSUBS 0.012241f
C718 B.n566 VSUBS 0.012241f
C719 B.n567 VSUBS 0.012241f
C720 B.n568 VSUBS 0.012241f
C721 B.n569 VSUBS 0.012241f
C722 B.n570 VSUBS 0.012241f
C723 B.n571 VSUBS 0.012241f
C724 B.n572 VSUBS 0.012241f
C725 B.n573 VSUBS 0.012241f
C726 B.n574 VSUBS 0.012241f
C727 B.n575 VSUBS 0.012241f
C728 B.n576 VSUBS 0.012241f
C729 B.n577 VSUBS 0.012241f
C730 B.n578 VSUBS 0.012241f
C731 B.n579 VSUBS 0.012241f
C732 B.n580 VSUBS 0.012241f
C733 B.n581 VSUBS 0.012241f
C734 B.n582 VSUBS 0.012241f
C735 B.n583 VSUBS 0.012241f
C736 B.n584 VSUBS 0.012241f
C737 B.n585 VSUBS 0.012241f
C738 B.n586 VSUBS 0.012241f
C739 B.n587 VSUBS 0.012241f
C740 B.n588 VSUBS 0.012241f
C741 B.n589 VSUBS 0.012241f
C742 B.n590 VSUBS 0.012241f
C743 B.n591 VSUBS 0.012241f
C744 B.n592 VSUBS 0.012241f
C745 B.n593 VSUBS 0.012241f
C746 B.n594 VSUBS 0.012241f
C747 B.n595 VSUBS 0.012241f
C748 B.n596 VSUBS 0.012241f
C749 B.n597 VSUBS 0.012241f
C750 B.n598 VSUBS 0.012241f
C751 B.n599 VSUBS 0.012241f
C752 B.n600 VSUBS 0.012241f
C753 B.n601 VSUBS 0.012241f
C754 B.n602 VSUBS 0.012241f
C755 B.n603 VSUBS 0.012241f
C756 B.n604 VSUBS 0.012241f
C757 B.n605 VSUBS 0.012241f
C758 B.n606 VSUBS 0.012241f
C759 B.n607 VSUBS 0.015973f
C760 B.n608 VSUBS 0.017016f
C761 B.n609 VSUBS 0.033838f
C762 VDD1.t5 VSUBS 0.140054f
C763 VDD1.t7 VSUBS 0.026413f
C764 VDD1.t2 VSUBS 0.026413f
C765 VDD1.n0 VSUBS 0.071527f
C766 VDD1.n1 VSUBS 1.16327f
C767 VDD1.t1 VSUBS 0.140054f
C768 VDD1.t0 VSUBS 0.026413f
C769 VDD1.t3 VSUBS 0.026413f
C770 VDD1.n2 VSUBS 0.071527f
C771 VDD1.n3 VSUBS 1.15248f
C772 VDD1.t6 VSUBS 0.026413f
C773 VDD1.t9 VSUBS 0.026413f
C774 VDD1.n4 VSUBS 0.073692f
C775 VDD1.n5 VSUBS 3.15884f
C776 VDD1.t4 VSUBS 0.026413f
C777 VDD1.t8 VSUBS 0.026413f
C778 VDD1.n6 VSUBS 0.071527f
C779 VDD1.n7 VSUBS 3.07362f
C780 VTAIL.t0 VSUBS 0.033879f
C781 VTAIL.t14 VSUBS 0.033879f
C782 VTAIL.n0 VSUBS 0.082906f
C783 VTAIL.n1 VSUBS 0.798263f
C784 VTAIL.t9 VSUBS 0.168363f
C785 VTAIL.n2 VSUBS 0.884498f
C786 VTAIL.t10 VSUBS 0.033879f
C787 VTAIL.t12 VSUBS 0.033879f
C788 VTAIL.n3 VSUBS 0.082906f
C789 VTAIL.n4 VSUBS 0.987805f
C790 VTAIL.t11 VSUBS 0.033879f
C791 VTAIL.t4 VSUBS 0.033879f
C792 VTAIL.n5 VSUBS 0.082906f
C793 VTAIL.n6 VSUBS 2.03251f
C794 VTAIL.t16 VSUBS 0.033879f
C795 VTAIL.t1 VSUBS 0.033879f
C796 VTAIL.n7 VSUBS 0.082906f
C797 VTAIL.n8 VSUBS 2.03251f
C798 VTAIL.t19 VSUBS 0.033879f
C799 VTAIL.t3 VSUBS 0.033879f
C800 VTAIL.n9 VSUBS 0.082906f
C801 VTAIL.n10 VSUBS 0.987804f
C802 VTAIL.t2 VSUBS 0.168363f
C803 VTAIL.n11 VSUBS 0.884498f
C804 VTAIL.t6 VSUBS 0.033879f
C805 VTAIL.t5 VSUBS 0.033879f
C806 VTAIL.n12 VSUBS 0.082906f
C807 VTAIL.n13 VSUBS 0.877558f
C808 VTAIL.t13 VSUBS 0.033879f
C809 VTAIL.t7 VSUBS 0.033879f
C810 VTAIL.n14 VSUBS 0.082906f
C811 VTAIL.n15 VSUBS 0.987804f
C812 VTAIL.t8 VSUBS 0.168363f
C813 VTAIL.n16 VSUBS 1.69044f
C814 VTAIL.t17 VSUBS 0.168363f
C815 VTAIL.n17 VSUBS 1.69044f
C816 VTAIL.t15 VSUBS 0.033879f
C817 VTAIL.t18 VSUBS 0.033879f
C818 VTAIL.n18 VSUBS 0.082906f
C819 VTAIL.n19 VSUBS 0.718084f
C820 VP.n0 VSUBS 0.088166f
C821 VP.t0 VSUBS 0.333523f
C822 VP.n1 VSUBS 0.108804f
C823 VP.n2 VSUBS 0.066873f
C824 VP.t3 VSUBS 0.333523f
C825 VP.n3 VSUBS 0.227473f
C826 VP.n4 VSUBS 0.066873f
C827 VP.n5 VSUBS 0.093896f
C828 VP.n6 VSUBS 0.066873f
C829 VP.t6 VSUBS 0.333523f
C830 VP.n7 VSUBS 0.124636f
C831 VP.n8 VSUBS 0.066873f
C832 VP.n9 VSUBS 0.088946f
C833 VP.n10 VSUBS 0.066873f
C834 VP.n11 VSUBS 0.108804f
C835 VP.n12 VSUBS 0.088166f
C836 VP.t8 VSUBS 0.333523f
C837 VP.n13 VSUBS 0.088166f
C838 VP.t1 VSUBS 0.333523f
C839 VP.n14 VSUBS 0.108804f
C840 VP.n15 VSUBS 0.066873f
C841 VP.t5 VSUBS 0.333523f
C842 VP.n16 VSUBS 0.227473f
C843 VP.n17 VSUBS 0.066873f
C844 VP.n18 VSUBS 0.093896f
C845 VP.n19 VSUBS 0.066873f
C846 VP.t7 VSUBS 0.333523f
C847 VP.n20 VSUBS 0.124636f
C848 VP.n21 VSUBS 0.066873f
C849 VP.n22 VSUBS 0.088946f
C850 VP.t4 VSUBS 0.836439f
C851 VP.t2 VSUBS 0.333523f
C852 VP.n23 VSUBS 0.416607f
C853 VP.n24 VSUBS 0.421794f
C854 VP.n25 VSUBS 0.648394f
C855 VP.n26 VSUBS 0.066873f
C856 VP.n27 VSUBS 0.124636f
C857 VP.n28 VSUBS 0.10135f
C858 VP.n29 VSUBS 0.093896f
C859 VP.n30 VSUBS 0.066873f
C860 VP.n31 VSUBS 0.066873f
C861 VP.n32 VSUBS 0.066873f
C862 VP.n33 VSUBS 0.093869f
C863 VP.n34 VSUBS 0.227473f
C864 VP.n35 VSUBS 0.093869f
C865 VP.n36 VSUBS 0.124636f
C866 VP.n37 VSUBS 0.066873f
C867 VP.n38 VSUBS 0.066873f
C868 VP.n39 VSUBS 0.066873f
C869 VP.n40 VSUBS 0.10135f
C870 VP.n41 VSUBS 0.124636f
C871 VP.n42 VSUBS 0.088946f
C872 VP.n43 VSUBS 0.066873f
C873 VP.n44 VSUBS 0.066873f
C874 VP.n45 VSUBS 0.098791f
C875 VP.n46 VSUBS 0.124636f
C876 VP.n47 VSUBS 0.086442f
C877 VP.n48 VSUBS 0.066873f
C878 VP.n49 VSUBS 0.066873f
C879 VP.n50 VSUBS 0.066873f
C880 VP.n51 VSUBS 0.124636f
C881 VP.n52 VSUBS 0.084024f
C882 VP.n53 VSUBS 0.448304f
C883 VP.n54 VSUBS 3.17254f
C884 VP.n55 VSUBS 3.22602f
C885 VP.n56 VSUBS 0.448304f
C886 VP.n57 VSUBS 0.084024f
C887 VP.n58 VSUBS 0.124636f
C888 VP.n59 VSUBS 0.066873f
C889 VP.n60 VSUBS 0.066873f
C890 VP.n61 VSUBS 0.066873f
C891 VP.n62 VSUBS 0.086442f
C892 VP.n63 VSUBS 0.124636f
C893 VP.t9 VSUBS 0.333523f
C894 VP.n64 VSUBS 0.227473f
C895 VP.n65 VSUBS 0.098791f
C896 VP.n66 VSUBS 0.066873f
C897 VP.n67 VSUBS 0.066873f
C898 VP.n68 VSUBS 0.066873f
C899 VP.n69 VSUBS 0.124636f
C900 VP.n70 VSUBS 0.10135f
C901 VP.n71 VSUBS 0.093896f
C902 VP.n72 VSUBS 0.066873f
C903 VP.n73 VSUBS 0.066873f
C904 VP.n74 VSUBS 0.066873f
C905 VP.n75 VSUBS 0.093869f
C906 VP.n76 VSUBS 0.227473f
C907 VP.n77 VSUBS 0.093869f
C908 VP.n78 VSUBS 0.124636f
C909 VP.n79 VSUBS 0.066873f
C910 VP.n80 VSUBS 0.066873f
C911 VP.n81 VSUBS 0.066873f
C912 VP.n82 VSUBS 0.10135f
C913 VP.n83 VSUBS 0.124636f
C914 VP.n84 VSUBS 0.088946f
C915 VP.n85 VSUBS 0.066873f
C916 VP.n86 VSUBS 0.066873f
C917 VP.n87 VSUBS 0.098791f
C918 VP.n88 VSUBS 0.124636f
C919 VP.n89 VSUBS 0.086442f
C920 VP.n90 VSUBS 0.066873f
C921 VP.n91 VSUBS 0.066873f
C922 VP.n92 VSUBS 0.066873f
C923 VP.n93 VSUBS 0.124636f
C924 VP.n94 VSUBS 0.084024f
C925 VP.n95 VSUBS 0.448304f
C926 VP.n96 VSUBS 0.112269f
.ends

