* NGSPICE file created from diff_pair_sample_0643.ext - technology: sky130A

.subckt diff_pair_sample_0643 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t7 VN.t0 VTAIL.t14 B.t6 sky130_fd_pr__nfet_01v8 ad=0.9306 pd=5.97 as=0.9306 ps=5.97 w=5.64 l=0.51
X1 B.t21 B.t19 B.t20 B.t9 sky130_fd_pr__nfet_01v8 ad=2.1996 pd=12.06 as=0 ps=0 w=5.64 l=0.51
X2 VTAIL.t3 VP.t0 VDD1.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=0.9306 pd=5.97 as=0.9306 ps=5.97 w=5.64 l=0.51
X3 VDD1.t6 VP.t1 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=0.9306 pd=5.97 as=0.9306 ps=5.97 w=5.64 l=0.51
X4 B.t18 B.t16 B.t17 B.t13 sky130_fd_pr__nfet_01v8 ad=2.1996 pd=12.06 as=0 ps=0 w=5.64 l=0.51
X5 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=2.1996 pd=12.06 as=0 ps=0 w=5.64 l=0.51
X6 VTAIL.t4 VP.t2 VDD1.t5 B.t4 sky130_fd_pr__nfet_01v8 ad=2.1996 pd=12.06 as=0.9306 ps=5.97 w=5.64 l=0.51
X7 VDD1.t4 VP.t3 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=0.9306 pd=5.97 as=0.9306 ps=5.97 w=5.64 l=0.51
X8 VTAIL.t11 VN.t1 VDD2.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=0.9306 pd=5.97 as=0.9306 ps=5.97 w=5.64 l=0.51
X9 VTAIL.t1 VP.t4 VDD1.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=2.1996 pd=12.06 as=0.9306 ps=5.97 w=5.64 l=0.51
X10 VTAIL.t10 VN.t2 VDD2.t5 B.t1 sky130_fd_pr__nfet_01v8 ad=2.1996 pd=12.06 as=0.9306 ps=5.97 w=5.64 l=0.51
X11 VDD2.t4 VN.t3 VTAIL.t13 B.t0 sky130_fd_pr__nfet_01v8 ad=0.9306 pd=5.97 as=2.1996 ps=12.06 w=5.64 l=0.51
X12 VDD2.t3 VN.t4 VTAIL.t12 B.t5 sky130_fd_pr__nfet_01v8 ad=0.9306 pd=5.97 as=0.9306 ps=5.97 w=5.64 l=0.51
X13 VDD1.t2 VP.t5 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.9306 pd=5.97 as=2.1996 ps=12.06 w=5.64 l=0.51
X14 VTAIL.t9 VN.t5 VDD2.t2 B.t7 sky130_fd_pr__nfet_01v8 ad=0.9306 pd=5.97 as=0.9306 ps=5.97 w=5.64 l=0.51
X15 VTAIL.t15 VN.t6 VDD2.t1 B.t4 sky130_fd_pr__nfet_01v8 ad=2.1996 pd=12.06 as=0.9306 ps=5.97 w=5.64 l=0.51
X16 VDD2.t0 VN.t7 VTAIL.t8 B.t2 sky130_fd_pr__nfet_01v8 ad=0.9306 pd=5.97 as=2.1996 ps=12.06 w=5.64 l=0.51
X17 VTAIL.t7 VP.t6 VDD1.t1 B.t7 sky130_fd_pr__nfet_01v8 ad=0.9306 pd=5.97 as=0.9306 ps=5.97 w=5.64 l=0.51
X18 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=2.1996 pd=12.06 as=0 ps=0 w=5.64 l=0.51
X19 VDD1.t0 VP.t7 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.9306 pd=5.97 as=2.1996 ps=12.06 w=5.64 l=0.51
R0 VN.n2 VN.t2 364.978
R1 VN.n10 VN.t3 364.978
R2 VN.n6 VN.t7 344.274
R3 VN.n14 VN.t6 344.274
R4 VN.n1 VN.t4 343.543
R5 VN.n5 VN.t5 343.543
R6 VN.n9 VN.t1 343.543
R7 VN.n13 VN.t0 343.543
R8 VN.n7 VN.n6 161.3
R9 VN.n15 VN.n14 161.3
R10 VN.n13 VN.n8 161.3
R11 VN.n12 VN.n11 161.3
R12 VN.n5 VN.n0 161.3
R13 VN.n4 VN.n3 161.3
R14 VN.n11 VN.n10 70.5418
R15 VN.n3 VN.n2 70.5418
R16 VN.n6 VN.n5 47.4702
R17 VN.n14 VN.n13 47.4702
R18 VN VN.n15 36.7827
R19 VN.n4 VN.n1 24.1005
R20 VN.n5 VN.n4 24.1005
R21 VN.n13 VN.n12 24.1005
R22 VN.n12 VN.n9 24.1005
R23 VN.n10 VN.n9 20.6807
R24 VN.n2 VN.n1 20.6807
R25 VN.n15 VN.n8 0.189894
R26 VN.n11 VN.n8 0.189894
R27 VN.n3 VN.n0 0.189894
R28 VN.n7 VN.n0 0.189894
R29 VN VN.n7 0.0516364
R30 VTAIL.n11 VTAIL.t1 54.7019
R31 VTAIL.n10 VTAIL.t13 54.7019
R32 VTAIL.n7 VTAIL.t15 54.7019
R33 VTAIL.n15 VTAIL.t8 54.7017
R34 VTAIL.n2 VTAIL.t10 54.7017
R35 VTAIL.n3 VTAIL.t0 54.7017
R36 VTAIL.n6 VTAIL.t4 54.7017
R37 VTAIL.n14 VTAIL.t2 54.7017
R38 VTAIL.n13 VTAIL.n12 51.1912
R39 VTAIL.n9 VTAIL.n8 51.1912
R40 VTAIL.n1 VTAIL.n0 51.191
R41 VTAIL.n5 VTAIL.n4 51.191
R42 VTAIL.n15 VTAIL.n14 17.9531
R43 VTAIL.n7 VTAIL.n6 17.9531
R44 VTAIL.n0 VTAIL.t12 3.51114
R45 VTAIL.n0 VTAIL.t9 3.51114
R46 VTAIL.n4 VTAIL.t6 3.51114
R47 VTAIL.n4 VTAIL.t3 3.51114
R48 VTAIL.n12 VTAIL.t5 3.51114
R49 VTAIL.n12 VTAIL.t7 3.51114
R50 VTAIL.n8 VTAIL.t14 3.51114
R51 VTAIL.n8 VTAIL.t11 3.51114
R52 VTAIL.n9 VTAIL.n7 0.724638
R53 VTAIL.n10 VTAIL.n9 0.724638
R54 VTAIL.n13 VTAIL.n11 0.724638
R55 VTAIL.n14 VTAIL.n13 0.724638
R56 VTAIL.n6 VTAIL.n5 0.724638
R57 VTAIL.n5 VTAIL.n3 0.724638
R58 VTAIL.n2 VTAIL.n1 0.724638
R59 VTAIL VTAIL.n15 0.666448
R60 VTAIL.n11 VTAIL.n10 0.470328
R61 VTAIL.n3 VTAIL.n2 0.470328
R62 VTAIL VTAIL.n1 0.0586897
R63 VDD2.n2 VDD2.n1 68.1765
R64 VDD2.n2 VDD2.n0 68.1765
R65 VDD2 VDD2.n5 68.1737
R66 VDD2.n4 VDD2.n3 67.87
R67 VDD2.n4 VDD2.n2 31.836
R68 VDD2.n5 VDD2.t6 3.51114
R69 VDD2.n5 VDD2.t4 3.51114
R70 VDD2.n3 VDD2.t1 3.51114
R71 VDD2.n3 VDD2.t7 3.51114
R72 VDD2.n1 VDD2.t2 3.51114
R73 VDD2.n1 VDD2.t0 3.51114
R74 VDD2.n0 VDD2.t5 3.51114
R75 VDD2.n0 VDD2.t3 3.51114
R76 VDD2 VDD2.n4 0.420759
R77 B.n451 B.n450 585
R78 B.n452 B.n451 585
R79 B.n180 B.n69 585
R80 B.n179 B.n178 585
R81 B.n177 B.n176 585
R82 B.n175 B.n174 585
R83 B.n173 B.n172 585
R84 B.n171 B.n170 585
R85 B.n169 B.n168 585
R86 B.n167 B.n166 585
R87 B.n165 B.n164 585
R88 B.n163 B.n162 585
R89 B.n161 B.n160 585
R90 B.n159 B.n158 585
R91 B.n157 B.n156 585
R92 B.n155 B.n154 585
R93 B.n153 B.n152 585
R94 B.n151 B.n150 585
R95 B.n149 B.n148 585
R96 B.n147 B.n146 585
R97 B.n145 B.n144 585
R98 B.n143 B.n142 585
R99 B.n141 B.n140 585
R100 B.n139 B.n138 585
R101 B.n137 B.n136 585
R102 B.n135 B.n134 585
R103 B.n133 B.n132 585
R104 B.n131 B.n130 585
R105 B.n129 B.n128 585
R106 B.n127 B.n126 585
R107 B.n125 B.n124 585
R108 B.n123 B.n122 585
R109 B.n121 B.n120 585
R110 B.n118 B.n117 585
R111 B.n116 B.n115 585
R112 B.n114 B.n113 585
R113 B.n112 B.n111 585
R114 B.n110 B.n109 585
R115 B.n108 B.n107 585
R116 B.n106 B.n105 585
R117 B.n104 B.n103 585
R118 B.n102 B.n101 585
R119 B.n100 B.n99 585
R120 B.n98 B.n97 585
R121 B.n96 B.n95 585
R122 B.n94 B.n93 585
R123 B.n92 B.n91 585
R124 B.n90 B.n89 585
R125 B.n88 B.n87 585
R126 B.n86 B.n85 585
R127 B.n84 B.n83 585
R128 B.n82 B.n81 585
R129 B.n80 B.n79 585
R130 B.n78 B.n77 585
R131 B.n76 B.n75 585
R132 B.n40 B.n39 585
R133 B.n449 B.n41 585
R134 B.n453 B.n41 585
R135 B.n448 B.n447 585
R136 B.n447 B.n37 585
R137 B.n446 B.n36 585
R138 B.n459 B.n36 585
R139 B.n445 B.n35 585
R140 B.n460 B.n35 585
R141 B.n444 B.n34 585
R142 B.n461 B.n34 585
R143 B.n443 B.n442 585
R144 B.n442 B.n30 585
R145 B.n441 B.n29 585
R146 B.n467 B.n29 585
R147 B.n440 B.n28 585
R148 B.n468 B.n28 585
R149 B.n439 B.n27 585
R150 B.n469 B.n27 585
R151 B.n438 B.n437 585
R152 B.n437 B.n23 585
R153 B.n436 B.n22 585
R154 B.n475 B.n22 585
R155 B.n435 B.n21 585
R156 B.n476 B.n21 585
R157 B.n434 B.n20 585
R158 B.n477 B.n20 585
R159 B.n433 B.n432 585
R160 B.n432 B.n16 585
R161 B.n431 B.n15 585
R162 B.n483 B.n15 585
R163 B.n430 B.n14 585
R164 B.n484 B.n14 585
R165 B.n429 B.n13 585
R166 B.n485 B.n13 585
R167 B.n428 B.n427 585
R168 B.n427 B.n12 585
R169 B.n426 B.n425 585
R170 B.n426 B.n8 585
R171 B.n424 B.n7 585
R172 B.n492 B.n7 585
R173 B.n423 B.n6 585
R174 B.n493 B.n6 585
R175 B.n422 B.n5 585
R176 B.n494 B.n5 585
R177 B.n421 B.n420 585
R178 B.n420 B.n4 585
R179 B.n419 B.n181 585
R180 B.n419 B.n418 585
R181 B.n408 B.n182 585
R182 B.n411 B.n182 585
R183 B.n410 B.n409 585
R184 B.n412 B.n410 585
R185 B.n407 B.n186 585
R186 B.n190 B.n186 585
R187 B.n406 B.n405 585
R188 B.n405 B.n404 585
R189 B.n188 B.n187 585
R190 B.n189 B.n188 585
R191 B.n397 B.n396 585
R192 B.n398 B.n397 585
R193 B.n395 B.n195 585
R194 B.n195 B.n194 585
R195 B.n394 B.n393 585
R196 B.n393 B.n392 585
R197 B.n197 B.n196 585
R198 B.n198 B.n197 585
R199 B.n385 B.n384 585
R200 B.n386 B.n385 585
R201 B.n383 B.n203 585
R202 B.n203 B.n202 585
R203 B.n382 B.n381 585
R204 B.n381 B.n380 585
R205 B.n205 B.n204 585
R206 B.n206 B.n205 585
R207 B.n373 B.n372 585
R208 B.n374 B.n373 585
R209 B.n371 B.n211 585
R210 B.n211 B.n210 585
R211 B.n370 B.n369 585
R212 B.n369 B.n368 585
R213 B.n213 B.n212 585
R214 B.n214 B.n213 585
R215 B.n361 B.n360 585
R216 B.n362 B.n361 585
R217 B.n217 B.n216 585
R218 B.n250 B.n249 585
R219 B.n251 B.n247 585
R220 B.n247 B.n218 585
R221 B.n253 B.n252 585
R222 B.n255 B.n246 585
R223 B.n258 B.n257 585
R224 B.n259 B.n245 585
R225 B.n261 B.n260 585
R226 B.n263 B.n244 585
R227 B.n266 B.n265 585
R228 B.n267 B.n243 585
R229 B.n269 B.n268 585
R230 B.n271 B.n242 585
R231 B.n274 B.n273 585
R232 B.n275 B.n241 585
R233 B.n277 B.n276 585
R234 B.n279 B.n240 585
R235 B.n282 B.n281 585
R236 B.n283 B.n239 585
R237 B.n285 B.n284 585
R238 B.n287 B.n238 585
R239 B.n290 B.n289 585
R240 B.n291 B.n235 585
R241 B.n294 B.n293 585
R242 B.n296 B.n234 585
R243 B.n299 B.n298 585
R244 B.n300 B.n233 585
R245 B.n302 B.n301 585
R246 B.n304 B.n232 585
R247 B.n307 B.n306 585
R248 B.n308 B.n231 585
R249 B.n313 B.n312 585
R250 B.n315 B.n230 585
R251 B.n318 B.n317 585
R252 B.n319 B.n229 585
R253 B.n321 B.n320 585
R254 B.n323 B.n228 585
R255 B.n326 B.n325 585
R256 B.n327 B.n227 585
R257 B.n329 B.n328 585
R258 B.n331 B.n226 585
R259 B.n334 B.n333 585
R260 B.n335 B.n225 585
R261 B.n337 B.n336 585
R262 B.n339 B.n224 585
R263 B.n342 B.n341 585
R264 B.n343 B.n223 585
R265 B.n345 B.n344 585
R266 B.n347 B.n222 585
R267 B.n350 B.n349 585
R268 B.n351 B.n221 585
R269 B.n353 B.n352 585
R270 B.n355 B.n220 585
R271 B.n358 B.n357 585
R272 B.n359 B.n219 585
R273 B.n364 B.n363 585
R274 B.n363 B.n362 585
R275 B.n365 B.n215 585
R276 B.n215 B.n214 585
R277 B.n367 B.n366 585
R278 B.n368 B.n367 585
R279 B.n209 B.n208 585
R280 B.n210 B.n209 585
R281 B.n376 B.n375 585
R282 B.n375 B.n374 585
R283 B.n377 B.n207 585
R284 B.n207 B.n206 585
R285 B.n379 B.n378 585
R286 B.n380 B.n379 585
R287 B.n201 B.n200 585
R288 B.n202 B.n201 585
R289 B.n388 B.n387 585
R290 B.n387 B.n386 585
R291 B.n389 B.n199 585
R292 B.n199 B.n198 585
R293 B.n391 B.n390 585
R294 B.n392 B.n391 585
R295 B.n193 B.n192 585
R296 B.n194 B.n193 585
R297 B.n400 B.n399 585
R298 B.n399 B.n398 585
R299 B.n401 B.n191 585
R300 B.n191 B.n189 585
R301 B.n403 B.n402 585
R302 B.n404 B.n403 585
R303 B.n185 B.n184 585
R304 B.n190 B.n185 585
R305 B.n414 B.n413 585
R306 B.n413 B.n412 585
R307 B.n415 B.n183 585
R308 B.n411 B.n183 585
R309 B.n417 B.n416 585
R310 B.n418 B.n417 585
R311 B.n3 B.n0 585
R312 B.n4 B.n3 585
R313 B.n491 B.n1 585
R314 B.n492 B.n491 585
R315 B.n490 B.n489 585
R316 B.n490 B.n8 585
R317 B.n488 B.n9 585
R318 B.n12 B.n9 585
R319 B.n487 B.n486 585
R320 B.n486 B.n485 585
R321 B.n11 B.n10 585
R322 B.n484 B.n11 585
R323 B.n482 B.n481 585
R324 B.n483 B.n482 585
R325 B.n480 B.n17 585
R326 B.n17 B.n16 585
R327 B.n479 B.n478 585
R328 B.n478 B.n477 585
R329 B.n19 B.n18 585
R330 B.n476 B.n19 585
R331 B.n474 B.n473 585
R332 B.n475 B.n474 585
R333 B.n472 B.n24 585
R334 B.n24 B.n23 585
R335 B.n471 B.n470 585
R336 B.n470 B.n469 585
R337 B.n26 B.n25 585
R338 B.n468 B.n26 585
R339 B.n466 B.n465 585
R340 B.n467 B.n466 585
R341 B.n464 B.n31 585
R342 B.n31 B.n30 585
R343 B.n463 B.n462 585
R344 B.n462 B.n461 585
R345 B.n33 B.n32 585
R346 B.n460 B.n33 585
R347 B.n458 B.n457 585
R348 B.n459 B.n458 585
R349 B.n456 B.n38 585
R350 B.n38 B.n37 585
R351 B.n455 B.n454 585
R352 B.n454 B.n453 585
R353 B.n495 B.n494 585
R354 B.n493 B.n2 585
R355 B.n454 B.n40 526.135
R356 B.n451 B.n41 526.135
R357 B.n361 B.n219 526.135
R358 B.n363 B.n217 526.135
R359 B.n73 B.t19 472.69
R360 B.n70 B.t8 472.69
R361 B.n309 B.t16 472.69
R362 B.n236 B.t12 472.69
R363 B.n452 B.n68 256.663
R364 B.n452 B.n67 256.663
R365 B.n452 B.n66 256.663
R366 B.n452 B.n65 256.663
R367 B.n452 B.n64 256.663
R368 B.n452 B.n63 256.663
R369 B.n452 B.n62 256.663
R370 B.n452 B.n61 256.663
R371 B.n452 B.n60 256.663
R372 B.n452 B.n59 256.663
R373 B.n452 B.n58 256.663
R374 B.n452 B.n57 256.663
R375 B.n452 B.n56 256.663
R376 B.n452 B.n55 256.663
R377 B.n452 B.n54 256.663
R378 B.n452 B.n53 256.663
R379 B.n452 B.n52 256.663
R380 B.n452 B.n51 256.663
R381 B.n452 B.n50 256.663
R382 B.n452 B.n49 256.663
R383 B.n452 B.n48 256.663
R384 B.n452 B.n47 256.663
R385 B.n452 B.n46 256.663
R386 B.n452 B.n45 256.663
R387 B.n452 B.n44 256.663
R388 B.n452 B.n43 256.663
R389 B.n452 B.n42 256.663
R390 B.n248 B.n218 256.663
R391 B.n254 B.n218 256.663
R392 B.n256 B.n218 256.663
R393 B.n262 B.n218 256.663
R394 B.n264 B.n218 256.663
R395 B.n270 B.n218 256.663
R396 B.n272 B.n218 256.663
R397 B.n278 B.n218 256.663
R398 B.n280 B.n218 256.663
R399 B.n286 B.n218 256.663
R400 B.n288 B.n218 256.663
R401 B.n295 B.n218 256.663
R402 B.n297 B.n218 256.663
R403 B.n303 B.n218 256.663
R404 B.n305 B.n218 256.663
R405 B.n314 B.n218 256.663
R406 B.n316 B.n218 256.663
R407 B.n322 B.n218 256.663
R408 B.n324 B.n218 256.663
R409 B.n330 B.n218 256.663
R410 B.n332 B.n218 256.663
R411 B.n338 B.n218 256.663
R412 B.n340 B.n218 256.663
R413 B.n346 B.n218 256.663
R414 B.n348 B.n218 256.663
R415 B.n354 B.n218 256.663
R416 B.n356 B.n218 256.663
R417 B.n497 B.n496 256.663
R418 B.n77 B.n76 163.367
R419 B.n81 B.n80 163.367
R420 B.n85 B.n84 163.367
R421 B.n89 B.n88 163.367
R422 B.n93 B.n92 163.367
R423 B.n97 B.n96 163.367
R424 B.n101 B.n100 163.367
R425 B.n105 B.n104 163.367
R426 B.n109 B.n108 163.367
R427 B.n113 B.n112 163.367
R428 B.n117 B.n116 163.367
R429 B.n122 B.n121 163.367
R430 B.n126 B.n125 163.367
R431 B.n130 B.n129 163.367
R432 B.n134 B.n133 163.367
R433 B.n138 B.n137 163.367
R434 B.n142 B.n141 163.367
R435 B.n146 B.n145 163.367
R436 B.n150 B.n149 163.367
R437 B.n154 B.n153 163.367
R438 B.n158 B.n157 163.367
R439 B.n162 B.n161 163.367
R440 B.n166 B.n165 163.367
R441 B.n170 B.n169 163.367
R442 B.n174 B.n173 163.367
R443 B.n178 B.n177 163.367
R444 B.n451 B.n69 163.367
R445 B.n361 B.n213 163.367
R446 B.n369 B.n213 163.367
R447 B.n369 B.n211 163.367
R448 B.n373 B.n211 163.367
R449 B.n373 B.n205 163.367
R450 B.n381 B.n205 163.367
R451 B.n381 B.n203 163.367
R452 B.n385 B.n203 163.367
R453 B.n385 B.n197 163.367
R454 B.n393 B.n197 163.367
R455 B.n393 B.n195 163.367
R456 B.n397 B.n195 163.367
R457 B.n397 B.n188 163.367
R458 B.n405 B.n188 163.367
R459 B.n405 B.n186 163.367
R460 B.n410 B.n186 163.367
R461 B.n410 B.n182 163.367
R462 B.n419 B.n182 163.367
R463 B.n420 B.n419 163.367
R464 B.n420 B.n5 163.367
R465 B.n6 B.n5 163.367
R466 B.n7 B.n6 163.367
R467 B.n426 B.n7 163.367
R468 B.n427 B.n426 163.367
R469 B.n427 B.n13 163.367
R470 B.n14 B.n13 163.367
R471 B.n15 B.n14 163.367
R472 B.n432 B.n15 163.367
R473 B.n432 B.n20 163.367
R474 B.n21 B.n20 163.367
R475 B.n22 B.n21 163.367
R476 B.n437 B.n22 163.367
R477 B.n437 B.n27 163.367
R478 B.n28 B.n27 163.367
R479 B.n29 B.n28 163.367
R480 B.n442 B.n29 163.367
R481 B.n442 B.n34 163.367
R482 B.n35 B.n34 163.367
R483 B.n36 B.n35 163.367
R484 B.n447 B.n36 163.367
R485 B.n447 B.n41 163.367
R486 B.n249 B.n247 163.367
R487 B.n253 B.n247 163.367
R488 B.n257 B.n255 163.367
R489 B.n261 B.n245 163.367
R490 B.n265 B.n263 163.367
R491 B.n269 B.n243 163.367
R492 B.n273 B.n271 163.367
R493 B.n277 B.n241 163.367
R494 B.n281 B.n279 163.367
R495 B.n285 B.n239 163.367
R496 B.n289 B.n287 163.367
R497 B.n294 B.n235 163.367
R498 B.n298 B.n296 163.367
R499 B.n302 B.n233 163.367
R500 B.n306 B.n304 163.367
R501 B.n313 B.n231 163.367
R502 B.n317 B.n315 163.367
R503 B.n321 B.n229 163.367
R504 B.n325 B.n323 163.367
R505 B.n329 B.n227 163.367
R506 B.n333 B.n331 163.367
R507 B.n337 B.n225 163.367
R508 B.n341 B.n339 163.367
R509 B.n345 B.n223 163.367
R510 B.n349 B.n347 163.367
R511 B.n353 B.n221 163.367
R512 B.n357 B.n355 163.367
R513 B.n363 B.n215 163.367
R514 B.n367 B.n215 163.367
R515 B.n367 B.n209 163.367
R516 B.n375 B.n209 163.367
R517 B.n375 B.n207 163.367
R518 B.n379 B.n207 163.367
R519 B.n379 B.n201 163.367
R520 B.n387 B.n201 163.367
R521 B.n387 B.n199 163.367
R522 B.n391 B.n199 163.367
R523 B.n391 B.n193 163.367
R524 B.n399 B.n193 163.367
R525 B.n399 B.n191 163.367
R526 B.n403 B.n191 163.367
R527 B.n403 B.n185 163.367
R528 B.n413 B.n185 163.367
R529 B.n413 B.n183 163.367
R530 B.n417 B.n183 163.367
R531 B.n417 B.n3 163.367
R532 B.n495 B.n3 163.367
R533 B.n491 B.n2 163.367
R534 B.n491 B.n490 163.367
R535 B.n490 B.n9 163.367
R536 B.n486 B.n9 163.367
R537 B.n486 B.n11 163.367
R538 B.n482 B.n11 163.367
R539 B.n482 B.n17 163.367
R540 B.n478 B.n17 163.367
R541 B.n478 B.n19 163.367
R542 B.n474 B.n19 163.367
R543 B.n474 B.n24 163.367
R544 B.n470 B.n24 163.367
R545 B.n470 B.n26 163.367
R546 B.n466 B.n26 163.367
R547 B.n466 B.n31 163.367
R548 B.n462 B.n31 163.367
R549 B.n462 B.n33 163.367
R550 B.n458 B.n33 163.367
R551 B.n458 B.n38 163.367
R552 B.n454 B.n38 163.367
R553 B.n362 B.n218 121.942
R554 B.n453 B.n452 121.942
R555 B.n70 B.t10 89.8447
R556 B.n309 B.t18 89.8447
R557 B.n73 B.t20 89.8389
R558 B.n236 B.t15 89.8389
R559 B.n71 B.t11 73.5538
R560 B.n310 B.t17 73.5538
R561 B.n74 B.t21 73.548
R562 B.n237 B.t14 73.548
R563 B.n42 B.n40 71.676
R564 B.n77 B.n43 71.676
R565 B.n81 B.n44 71.676
R566 B.n85 B.n45 71.676
R567 B.n89 B.n46 71.676
R568 B.n93 B.n47 71.676
R569 B.n97 B.n48 71.676
R570 B.n101 B.n49 71.676
R571 B.n105 B.n50 71.676
R572 B.n109 B.n51 71.676
R573 B.n113 B.n52 71.676
R574 B.n117 B.n53 71.676
R575 B.n122 B.n54 71.676
R576 B.n126 B.n55 71.676
R577 B.n130 B.n56 71.676
R578 B.n134 B.n57 71.676
R579 B.n138 B.n58 71.676
R580 B.n142 B.n59 71.676
R581 B.n146 B.n60 71.676
R582 B.n150 B.n61 71.676
R583 B.n154 B.n62 71.676
R584 B.n158 B.n63 71.676
R585 B.n162 B.n64 71.676
R586 B.n166 B.n65 71.676
R587 B.n170 B.n66 71.676
R588 B.n174 B.n67 71.676
R589 B.n178 B.n68 71.676
R590 B.n69 B.n68 71.676
R591 B.n177 B.n67 71.676
R592 B.n173 B.n66 71.676
R593 B.n169 B.n65 71.676
R594 B.n165 B.n64 71.676
R595 B.n161 B.n63 71.676
R596 B.n157 B.n62 71.676
R597 B.n153 B.n61 71.676
R598 B.n149 B.n60 71.676
R599 B.n145 B.n59 71.676
R600 B.n141 B.n58 71.676
R601 B.n137 B.n57 71.676
R602 B.n133 B.n56 71.676
R603 B.n129 B.n55 71.676
R604 B.n125 B.n54 71.676
R605 B.n121 B.n53 71.676
R606 B.n116 B.n52 71.676
R607 B.n112 B.n51 71.676
R608 B.n108 B.n50 71.676
R609 B.n104 B.n49 71.676
R610 B.n100 B.n48 71.676
R611 B.n96 B.n47 71.676
R612 B.n92 B.n46 71.676
R613 B.n88 B.n45 71.676
R614 B.n84 B.n44 71.676
R615 B.n80 B.n43 71.676
R616 B.n76 B.n42 71.676
R617 B.n248 B.n217 71.676
R618 B.n254 B.n253 71.676
R619 B.n257 B.n256 71.676
R620 B.n262 B.n261 71.676
R621 B.n265 B.n264 71.676
R622 B.n270 B.n269 71.676
R623 B.n273 B.n272 71.676
R624 B.n278 B.n277 71.676
R625 B.n281 B.n280 71.676
R626 B.n286 B.n285 71.676
R627 B.n289 B.n288 71.676
R628 B.n295 B.n294 71.676
R629 B.n298 B.n297 71.676
R630 B.n303 B.n302 71.676
R631 B.n306 B.n305 71.676
R632 B.n314 B.n313 71.676
R633 B.n317 B.n316 71.676
R634 B.n322 B.n321 71.676
R635 B.n325 B.n324 71.676
R636 B.n330 B.n329 71.676
R637 B.n333 B.n332 71.676
R638 B.n338 B.n337 71.676
R639 B.n341 B.n340 71.676
R640 B.n346 B.n345 71.676
R641 B.n349 B.n348 71.676
R642 B.n354 B.n353 71.676
R643 B.n357 B.n356 71.676
R644 B.n249 B.n248 71.676
R645 B.n255 B.n254 71.676
R646 B.n256 B.n245 71.676
R647 B.n263 B.n262 71.676
R648 B.n264 B.n243 71.676
R649 B.n271 B.n270 71.676
R650 B.n272 B.n241 71.676
R651 B.n279 B.n278 71.676
R652 B.n280 B.n239 71.676
R653 B.n287 B.n286 71.676
R654 B.n288 B.n235 71.676
R655 B.n296 B.n295 71.676
R656 B.n297 B.n233 71.676
R657 B.n304 B.n303 71.676
R658 B.n305 B.n231 71.676
R659 B.n315 B.n314 71.676
R660 B.n316 B.n229 71.676
R661 B.n323 B.n322 71.676
R662 B.n324 B.n227 71.676
R663 B.n331 B.n330 71.676
R664 B.n332 B.n225 71.676
R665 B.n339 B.n338 71.676
R666 B.n340 B.n223 71.676
R667 B.n347 B.n346 71.676
R668 B.n348 B.n221 71.676
R669 B.n355 B.n354 71.676
R670 B.n356 B.n219 71.676
R671 B.n496 B.n495 71.676
R672 B.n496 B.n2 71.676
R673 B.n362 B.n214 68.53
R674 B.n368 B.n214 68.53
R675 B.n368 B.n210 68.53
R676 B.n374 B.n210 68.53
R677 B.n380 B.n206 68.53
R678 B.n380 B.n202 68.53
R679 B.n386 B.n202 68.53
R680 B.n386 B.n198 68.53
R681 B.n392 B.n198 68.53
R682 B.n398 B.n194 68.53
R683 B.n404 B.n189 68.53
R684 B.n404 B.n190 68.53
R685 B.n412 B.n411 68.53
R686 B.n418 B.n4 68.53
R687 B.n494 B.n4 68.53
R688 B.n494 B.n493 68.53
R689 B.n493 B.n492 68.53
R690 B.n492 B.n8 68.53
R691 B.n485 B.n12 68.53
R692 B.n484 B.n483 68.53
R693 B.n483 B.n16 68.53
R694 B.n477 B.n476 68.53
R695 B.n475 B.n23 68.53
R696 B.n469 B.n23 68.53
R697 B.n469 B.n468 68.53
R698 B.n468 B.n467 68.53
R699 B.n467 B.n30 68.53
R700 B.n461 B.n460 68.53
R701 B.n460 B.n459 68.53
R702 B.n459 B.n37 68.53
R703 B.n453 B.n37 68.53
R704 B.n119 B.n74 59.5399
R705 B.n72 B.n71 59.5399
R706 B.n311 B.n310 59.5399
R707 B.n292 B.n237 59.5399
R708 B.n412 B.t3 55.4288
R709 B.n485 B.t5 55.4288
R710 B.t4 B.n194 51.3977
R711 B.n476 B.t2 51.3977
R712 B.n398 B.t6 49.3821
R713 B.n477 B.t7 49.3821
R714 B.n411 B.t0 45.3509
R715 B.n12 B.t1 45.3509
R716 B.n374 B.t13 39.3042
R717 B.n461 B.t9 39.3042
R718 B.n364 B.n216 34.1859
R719 B.n360 B.n359 34.1859
R720 B.n450 B.n449 34.1859
R721 B.n455 B.n39 34.1859
R722 B.t13 B.n206 29.2263
R723 B.t9 B.n30 29.2263
R724 B.n418 B.t0 23.1796
R725 B.t1 B.n8 23.1796
R726 B.t6 B.n189 19.1485
R727 B.t7 B.n16 19.1485
R728 B B.n497 18.0485
R729 B.n392 B.t4 17.1329
R730 B.t2 B.n475 17.1329
R731 B.n74 B.n73 16.2914
R732 B.n71 B.n70 16.2914
R733 B.n310 B.n309 16.2914
R734 B.n237 B.n236 16.2914
R735 B.n190 B.t3 13.1017
R736 B.t5 B.n484 13.1017
R737 B.n365 B.n364 10.6151
R738 B.n366 B.n365 10.6151
R739 B.n366 B.n208 10.6151
R740 B.n376 B.n208 10.6151
R741 B.n377 B.n376 10.6151
R742 B.n378 B.n377 10.6151
R743 B.n378 B.n200 10.6151
R744 B.n388 B.n200 10.6151
R745 B.n389 B.n388 10.6151
R746 B.n390 B.n389 10.6151
R747 B.n390 B.n192 10.6151
R748 B.n400 B.n192 10.6151
R749 B.n401 B.n400 10.6151
R750 B.n402 B.n401 10.6151
R751 B.n402 B.n184 10.6151
R752 B.n414 B.n184 10.6151
R753 B.n415 B.n414 10.6151
R754 B.n416 B.n415 10.6151
R755 B.n416 B.n0 10.6151
R756 B.n250 B.n216 10.6151
R757 B.n251 B.n250 10.6151
R758 B.n252 B.n251 10.6151
R759 B.n252 B.n246 10.6151
R760 B.n258 B.n246 10.6151
R761 B.n259 B.n258 10.6151
R762 B.n260 B.n259 10.6151
R763 B.n260 B.n244 10.6151
R764 B.n266 B.n244 10.6151
R765 B.n267 B.n266 10.6151
R766 B.n268 B.n267 10.6151
R767 B.n268 B.n242 10.6151
R768 B.n274 B.n242 10.6151
R769 B.n275 B.n274 10.6151
R770 B.n276 B.n275 10.6151
R771 B.n276 B.n240 10.6151
R772 B.n282 B.n240 10.6151
R773 B.n283 B.n282 10.6151
R774 B.n284 B.n283 10.6151
R775 B.n284 B.n238 10.6151
R776 B.n290 B.n238 10.6151
R777 B.n291 B.n290 10.6151
R778 B.n293 B.n234 10.6151
R779 B.n299 B.n234 10.6151
R780 B.n300 B.n299 10.6151
R781 B.n301 B.n300 10.6151
R782 B.n301 B.n232 10.6151
R783 B.n307 B.n232 10.6151
R784 B.n308 B.n307 10.6151
R785 B.n312 B.n308 10.6151
R786 B.n318 B.n230 10.6151
R787 B.n319 B.n318 10.6151
R788 B.n320 B.n319 10.6151
R789 B.n320 B.n228 10.6151
R790 B.n326 B.n228 10.6151
R791 B.n327 B.n326 10.6151
R792 B.n328 B.n327 10.6151
R793 B.n328 B.n226 10.6151
R794 B.n334 B.n226 10.6151
R795 B.n335 B.n334 10.6151
R796 B.n336 B.n335 10.6151
R797 B.n336 B.n224 10.6151
R798 B.n342 B.n224 10.6151
R799 B.n343 B.n342 10.6151
R800 B.n344 B.n343 10.6151
R801 B.n344 B.n222 10.6151
R802 B.n350 B.n222 10.6151
R803 B.n351 B.n350 10.6151
R804 B.n352 B.n351 10.6151
R805 B.n352 B.n220 10.6151
R806 B.n358 B.n220 10.6151
R807 B.n359 B.n358 10.6151
R808 B.n360 B.n212 10.6151
R809 B.n370 B.n212 10.6151
R810 B.n371 B.n370 10.6151
R811 B.n372 B.n371 10.6151
R812 B.n372 B.n204 10.6151
R813 B.n382 B.n204 10.6151
R814 B.n383 B.n382 10.6151
R815 B.n384 B.n383 10.6151
R816 B.n384 B.n196 10.6151
R817 B.n394 B.n196 10.6151
R818 B.n395 B.n394 10.6151
R819 B.n396 B.n395 10.6151
R820 B.n396 B.n187 10.6151
R821 B.n406 B.n187 10.6151
R822 B.n407 B.n406 10.6151
R823 B.n409 B.n407 10.6151
R824 B.n409 B.n408 10.6151
R825 B.n408 B.n181 10.6151
R826 B.n421 B.n181 10.6151
R827 B.n422 B.n421 10.6151
R828 B.n423 B.n422 10.6151
R829 B.n424 B.n423 10.6151
R830 B.n425 B.n424 10.6151
R831 B.n428 B.n425 10.6151
R832 B.n429 B.n428 10.6151
R833 B.n430 B.n429 10.6151
R834 B.n431 B.n430 10.6151
R835 B.n433 B.n431 10.6151
R836 B.n434 B.n433 10.6151
R837 B.n435 B.n434 10.6151
R838 B.n436 B.n435 10.6151
R839 B.n438 B.n436 10.6151
R840 B.n439 B.n438 10.6151
R841 B.n440 B.n439 10.6151
R842 B.n441 B.n440 10.6151
R843 B.n443 B.n441 10.6151
R844 B.n444 B.n443 10.6151
R845 B.n445 B.n444 10.6151
R846 B.n446 B.n445 10.6151
R847 B.n448 B.n446 10.6151
R848 B.n449 B.n448 10.6151
R849 B.n489 B.n1 10.6151
R850 B.n489 B.n488 10.6151
R851 B.n488 B.n487 10.6151
R852 B.n487 B.n10 10.6151
R853 B.n481 B.n10 10.6151
R854 B.n481 B.n480 10.6151
R855 B.n480 B.n479 10.6151
R856 B.n479 B.n18 10.6151
R857 B.n473 B.n18 10.6151
R858 B.n473 B.n472 10.6151
R859 B.n472 B.n471 10.6151
R860 B.n471 B.n25 10.6151
R861 B.n465 B.n25 10.6151
R862 B.n465 B.n464 10.6151
R863 B.n464 B.n463 10.6151
R864 B.n463 B.n32 10.6151
R865 B.n457 B.n32 10.6151
R866 B.n457 B.n456 10.6151
R867 B.n456 B.n455 10.6151
R868 B.n75 B.n39 10.6151
R869 B.n78 B.n75 10.6151
R870 B.n79 B.n78 10.6151
R871 B.n82 B.n79 10.6151
R872 B.n83 B.n82 10.6151
R873 B.n86 B.n83 10.6151
R874 B.n87 B.n86 10.6151
R875 B.n90 B.n87 10.6151
R876 B.n91 B.n90 10.6151
R877 B.n94 B.n91 10.6151
R878 B.n95 B.n94 10.6151
R879 B.n98 B.n95 10.6151
R880 B.n99 B.n98 10.6151
R881 B.n102 B.n99 10.6151
R882 B.n103 B.n102 10.6151
R883 B.n106 B.n103 10.6151
R884 B.n107 B.n106 10.6151
R885 B.n110 B.n107 10.6151
R886 B.n111 B.n110 10.6151
R887 B.n114 B.n111 10.6151
R888 B.n115 B.n114 10.6151
R889 B.n118 B.n115 10.6151
R890 B.n123 B.n120 10.6151
R891 B.n124 B.n123 10.6151
R892 B.n127 B.n124 10.6151
R893 B.n128 B.n127 10.6151
R894 B.n131 B.n128 10.6151
R895 B.n132 B.n131 10.6151
R896 B.n135 B.n132 10.6151
R897 B.n136 B.n135 10.6151
R898 B.n140 B.n139 10.6151
R899 B.n143 B.n140 10.6151
R900 B.n144 B.n143 10.6151
R901 B.n147 B.n144 10.6151
R902 B.n148 B.n147 10.6151
R903 B.n151 B.n148 10.6151
R904 B.n152 B.n151 10.6151
R905 B.n155 B.n152 10.6151
R906 B.n156 B.n155 10.6151
R907 B.n159 B.n156 10.6151
R908 B.n160 B.n159 10.6151
R909 B.n163 B.n160 10.6151
R910 B.n164 B.n163 10.6151
R911 B.n167 B.n164 10.6151
R912 B.n168 B.n167 10.6151
R913 B.n171 B.n168 10.6151
R914 B.n172 B.n171 10.6151
R915 B.n175 B.n172 10.6151
R916 B.n176 B.n175 10.6151
R917 B.n179 B.n176 10.6151
R918 B.n180 B.n179 10.6151
R919 B.n450 B.n180 10.6151
R920 B.n497 B.n0 8.11757
R921 B.n497 B.n1 8.11757
R922 B.n293 B.n292 6.5566
R923 B.n312 B.n311 6.5566
R924 B.n120 B.n119 6.5566
R925 B.n136 B.n72 6.5566
R926 B.n292 B.n291 4.05904
R927 B.n311 B.n230 4.05904
R928 B.n119 B.n118 4.05904
R929 B.n139 B.n72 4.05904
R930 VP.n4 VP.t4 364.978
R931 VP.n16 VP.t7 344.274
R932 VP.n10 VP.t2 344.274
R933 VP.n8 VP.t5 344.274
R934 VP.n1 VP.t1 343.543
R935 VP.n15 VP.t0 343.543
R936 VP.n7 VP.t6 343.543
R937 VP.n3 VP.t3 343.543
R938 VP.n17 VP.n16 161.3
R939 VP.n6 VP.n5 161.3
R940 VP.n7 VP.n2 161.3
R941 VP.n9 VP.n8 161.3
R942 VP.n15 VP.n0 161.3
R943 VP.n14 VP.n13 161.3
R944 VP.n12 VP.n1 161.3
R945 VP.n11 VP.n10 161.3
R946 VP.n5 VP.n4 70.5418
R947 VP.n10 VP.n1 47.4702
R948 VP.n16 VP.n15 47.4702
R949 VP.n8 VP.n7 47.4702
R950 VP.n11 VP.n9 36.402
R951 VP.n14 VP.n1 24.1005
R952 VP.n15 VP.n14 24.1005
R953 VP.n6 VP.n3 24.1005
R954 VP.n7 VP.n6 24.1005
R955 VP.n4 VP.n3 20.6807
R956 VP.n5 VP.n2 0.189894
R957 VP.n9 VP.n2 0.189894
R958 VP.n12 VP.n11 0.189894
R959 VP.n13 VP.n12 0.189894
R960 VP.n13 VP.n0 0.189894
R961 VP.n17 VP.n0 0.189894
R962 VP VP.n17 0.0516364
R963 VDD1 VDD1.n0 68.2903
R964 VDD1.n3 VDD1.n2 68.1765
R965 VDD1.n3 VDD1.n1 68.1765
R966 VDD1.n5 VDD1.n4 67.8699
R967 VDD1.n5 VDD1.n3 32.419
R968 VDD1.n4 VDD1.t1 3.51114
R969 VDD1.n4 VDD1.t2 3.51114
R970 VDD1.n0 VDD1.t3 3.51114
R971 VDD1.n0 VDD1.t4 3.51114
R972 VDD1.n2 VDD1.t7 3.51114
R973 VDD1.n2 VDD1.t0 3.51114
R974 VDD1.n1 VDD1.t5 3.51114
R975 VDD1.n1 VDD1.t6 3.51114
R976 VDD1 VDD1.n5 0.304379
C0 VTAIL VP 2.37626f
C1 VDD1 VDD2 0.733039f
C2 VTAIL VDD2 7.09602f
C3 VTAIL VDD1 7.05561f
C4 VN VP 3.92296f
C5 VN VDD2 2.36877f
C6 VN VDD1 0.148283f
C7 VN VTAIL 2.36215f
C8 VP VDD2 0.297607f
C9 VP VDD1 2.51776f
C10 VDD2 B 2.812014f
C11 VDD1 B 3.026811f
C12 VTAIL B 5.068369f
C13 VN B 7.10894f
C14 VP B 5.383237f
C15 VDD1.t3 B 0.127073f
C16 VDD1.t4 B 0.127073f
C17 VDD1.n0 B 1.05381f
C18 VDD1.t5 B 0.127073f
C19 VDD1.t6 B 0.127073f
C20 VDD1.n1 B 1.05319f
C21 VDD1.t7 B 0.127073f
C22 VDD1.t0 B 0.127073f
C23 VDD1.n2 B 1.05319f
C24 VDD1.n3 B 1.97056f
C25 VDD1.t1 B 0.127073f
C26 VDD1.t2 B 0.127073f
C27 VDD1.n4 B 1.05167f
C28 VDD1.n5 B 1.98999f
C29 VP.n0 B 0.050683f
C30 VP.t1 B 0.423766f
C31 VP.n1 B 0.20798f
C32 VP.n2 B 0.050683f
C33 VP.t6 B 0.423766f
C34 VP.t3 B 0.423766f
C35 VP.n3 B 0.20798f
C36 VP.t4 B 0.435678f
C37 VP.n4 B 0.19162f
C38 VP.n5 B 0.168214f
C39 VP.n6 B 0.011501f
C40 VP.n7 B 0.20798f
C41 VP.t5 B 0.424173f
C42 VP.n8 B 0.20273f
C43 VP.n9 B 1.62681f
C44 VP.t2 B 0.424173f
C45 VP.n10 B 0.20273f
C46 VP.n11 B 1.67701f
C47 VP.n12 B 0.050683f
C48 VP.n13 B 0.050683f
C49 VP.n14 B 0.011501f
C50 VP.t0 B 0.423766f
C51 VP.n15 B 0.20798f
C52 VP.t7 B 0.424173f
C53 VP.n16 B 0.20273f
C54 VP.n17 B 0.039277f
C55 VDD2.t5 B 0.127144f
C56 VDD2.t3 B 0.127144f
C57 VDD2.n0 B 1.05378f
C58 VDD2.t2 B 0.127144f
C59 VDD2.t0 B 0.127144f
C60 VDD2.n1 B 1.05378f
C61 VDD2.n2 B 1.91032f
C62 VDD2.t1 B 0.127144f
C63 VDD2.t7 B 0.127144f
C64 VDD2.n3 B 1.05226f
C65 VDD2.n4 B 1.95776f
C66 VDD2.t6 B 0.127144f
C67 VDD2.t4 B 0.127144f
C68 VDD2.n5 B 1.05375f
C69 VTAIL.t12 B 0.102552f
C70 VTAIL.t9 B 0.102552f
C71 VTAIL.n0 B 0.789676f
C72 VTAIL.n1 B 0.271395f
C73 VTAIL.t10 B 1.00731f
C74 VTAIL.n2 B 0.363963f
C75 VTAIL.t0 B 1.00731f
C76 VTAIL.n3 B 0.363963f
C77 VTAIL.t6 B 0.102552f
C78 VTAIL.t3 B 0.102552f
C79 VTAIL.n4 B 0.789676f
C80 VTAIL.n5 B 0.32077f
C81 VTAIL.t4 B 1.00731f
C82 VTAIL.n6 B 1.05586f
C83 VTAIL.t15 B 1.00732f
C84 VTAIL.n7 B 1.05586f
C85 VTAIL.t14 B 0.102552f
C86 VTAIL.t11 B 0.102552f
C87 VTAIL.n8 B 0.78968f
C88 VTAIL.n9 B 0.320766f
C89 VTAIL.t13 B 1.00732f
C90 VTAIL.n10 B 0.363959f
C91 VTAIL.t1 B 1.00732f
C92 VTAIL.n11 B 0.363959f
C93 VTAIL.t5 B 0.102552f
C94 VTAIL.t7 B 0.102552f
C95 VTAIL.n12 B 0.78968f
C96 VTAIL.n13 B 0.320766f
C97 VTAIL.t2 B 1.00731f
C98 VTAIL.n14 B 1.05586f
C99 VTAIL.t8 B 1.00731f
C100 VTAIL.n15 B 1.05155f
C101 VN.n0 B 0.049704f
C102 VN.t4 B 0.415586f
C103 VN.n1 B 0.203965f
C104 VN.t2 B 0.427268f
C105 VN.n2 B 0.187922f
C106 VN.n3 B 0.164967f
C107 VN.n4 B 0.011279f
C108 VN.t5 B 0.415586f
C109 VN.n5 B 0.203965f
C110 VN.t7 B 0.415985f
C111 VN.n6 B 0.198817f
C112 VN.n7 B 0.038519f
C113 VN.n8 B 0.049704f
C114 VN.t6 B 0.415985f
C115 VN.t1 B 0.415586f
C116 VN.n9 B 0.203965f
C117 VN.t3 B 0.427268f
C118 VN.n10 B 0.187922f
C119 VN.n11 B 0.164967f
C120 VN.n12 B 0.011279f
C121 VN.t0 B 0.415586f
C122 VN.n13 B 0.203965f
C123 VN.n14 B 0.198817f
C124 VN.n15 B 1.62835f
.ends

