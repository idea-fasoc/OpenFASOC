* NGSPICE file created from diff_pair_sample_0342.ext - technology: sky130A

.subckt diff_pair_sample_0342 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t19 VN.t0 VDD2.t6 B.t22 sky130_fd_pr__nfet_01v8 ad=0.2739 pd=1.99 as=0.2739 ps=1.99 w=1.66 l=2.85
X1 VDD1.t9 VP.t0 VTAIL.t6 B.t20 sky130_fd_pr__nfet_01v8 ad=0.2739 pd=1.99 as=0.6474 ps=4.1 w=1.66 l=2.85
X2 VTAIL.t18 VN.t1 VDD2.t9 B.t3 sky130_fd_pr__nfet_01v8 ad=0.2739 pd=1.99 as=0.2739 ps=1.99 w=1.66 l=2.85
X3 B.t17 B.t15 B.t16 B.t12 sky130_fd_pr__nfet_01v8 ad=0.6474 pd=4.1 as=0 ps=0 w=1.66 l=2.85
X4 VTAIL.t17 VN.t2 VDD2.t5 B.t18 sky130_fd_pr__nfet_01v8 ad=0.2739 pd=1.99 as=0.2739 ps=1.99 w=1.66 l=2.85
X5 VDD2.t2 VN.t3 VTAIL.t16 B.t21 sky130_fd_pr__nfet_01v8 ad=0.6474 pd=4.1 as=0.2739 ps=1.99 w=1.66 l=2.85
X6 VDD1.t8 VP.t1 VTAIL.t9 B.t23 sky130_fd_pr__nfet_01v8 ad=0.2739 pd=1.99 as=0.2739 ps=1.99 w=1.66 l=2.85
X7 B.t14 B.t11 B.t13 B.t12 sky130_fd_pr__nfet_01v8 ad=0.6474 pd=4.1 as=0 ps=0 w=1.66 l=2.85
X8 VDD1.t7 VP.t2 VTAIL.t7 B.t21 sky130_fd_pr__nfet_01v8 ad=0.6474 pd=4.1 as=0.2739 ps=1.99 w=1.66 l=2.85
X9 VTAIL.t15 VN.t4 VDD2.t0 B.t19 sky130_fd_pr__nfet_01v8 ad=0.2739 pd=1.99 as=0.2739 ps=1.99 w=1.66 l=2.85
X10 VDD2.t1 VN.t5 VTAIL.t14 B.t2 sky130_fd_pr__nfet_01v8 ad=0.2739 pd=1.99 as=0.6474 ps=4.1 w=1.66 l=2.85
X11 VTAIL.t4 VP.t3 VDD1.t6 B.t18 sky130_fd_pr__nfet_01v8 ad=0.2739 pd=1.99 as=0.2739 ps=1.99 w=1.66 l=2.85
X12 B.t10 B.t8 B.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=0.6474 pd=4.1 as=0 ps=0 w=1.66 l=2.85
X13 VDD2.t8 VN.t6 VTAIL.t13 B.t1 sky130_fd_pr__nfet_01v8 ad=0.6474 pd=4.1 as=0.2739 ps=1.99 w=1.66 l=2.85
X14 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=0.6474 pd=4.1 as=0 ps=0 w=1.66 l=2.85
X15 VDD1.t5 VP.t4 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.2739 pd=1.99 as=0.6474 ps=4.1 w=1.66 l=2.85
X16 VDD1.t4 VP.t5 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.6474 pd=4.1 as=0.2739 ps=1.99 w=1.66 l=2.85
X17 VDD2.t3 VN.t7 VTAIL.t12 B.t20 sky130_fd_pr__nfet_01v8 ad=0.2739 pd=1.99 as=0.6474 ps=4.1 w=1.66 l=2.85
X18 VTAIL.t3 VP.t6 VDD1.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.2739 pd=1.99 as=0.2739 ps=1.99 w=1.66 l=2.85
X19 VDD2.t4 VN.t8 VTAIL.t11 B.t23 sky130_fd_pr__nfet_01v8 ad=0.2739 pd=1.99 as=0.2739 ps=1.99 w=1.66 l=2.85
X20 VTAIL.t8 VP.t7 VDD1.t2 B.t22 sky130_fd_pr__nfet_01v8 ad=0.2739 pd=1.99 as=0.2739 ps=1.99 w=1.66 l=2.85
X21 VTAIL.t5 VP.t8 VDD1.t1 B.t19 sky130_fd_pr__nfet_01v8 ad=0.2739 pd=1.99 as=0.2739 ps=1.99 w=1.66 l=2.85
X22 VDD2.t7 VN.t9 VTAIL.t10 B.t0 sky130_fd_pr__nfet_01v8 ad=0.2739 pd=1.99 as=0.2739 ps=1.99 w=1.66 l=2.85
X23 VDD1.t0 VP.t9 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.2739 pd=1.99 as=0.2739 ps=1.99 w=1.66 l=2.85
R0 VN.n85 VN.n44 161.3
R1 VN.n84 VN.n83 161.3
R2 VN.n82 VN.n45 161.3
R3 VN.n81 VN.n80 161.3
R4 VN.n79 VN.n46 161.3
R5 VN.n78 VN.n77 161.3
R6 VN.n76 VN.n47 161.3
R7 VN.n75 VN.n74 161.3
R8 VN.n73 VN.n48 161.3
R9 VN.n72 VN.n71 161.3
R10 VN.n70 VN.n50 161.3
R11 VN.n69 VN.n68 161.3
R12 VN.n67 VN.n51 161.3
R13 VN.n65 VN.n64 161.3
R14 VN.n63 VN.n52 161.3
R15 VN.n62 VN.n61 161.3
R16 VN.n60 VN.n53 161.3
R17 VN.n59 VN.n58 161.3
R18 VN.n57 VN.n54 161.3
R19 VN.n41 VN.n0 161.3
R20 VN.n40 VN.n39 161.3
R21 VN.n38 VN.n1 161.3
R22 VN.n37 VN.n36 161.3
R23 VN.n35 VN.n2 161.3
R24 VN.n34 VN.n33 161.3
R25 VN.n32 VN.n3 161.3
R26 VN.n31 VN.n30 161.3
R27 VN.n28 VN.n4 161.3
R28 VN.n27 VN.n26 161.3
R29 VN.n25 VN.n5 161.3
R30 VN.n24 VN.n23 161.3
R31 VN.n22 VN.n6 161.3
R32 VN.n20 VN.n19 161.3
R33 VN.n18 VN.n7 161.3
R34 VN.n17 VN.n16 161.3
R35 VN.n15 VN.n8 161.3
R36 VN.n14 VN.n13 161.3
R37 VN.n12 VN.n9 161.3
R38 VN.n43 VN.n42 105.499
R39 VN.n87 VN.n86 105.499
R40 VN.n16 VN.n15 56.0773
R41 VN.n27 VN.n5 56.0773
R42 VN.n61 VN.n60 56.0773
R43 VN.n72 VN.n50 56.0773
R44 VN.n11 VN.n10 52.6217
R45 VN.n56 VN.n55 52.6217
R46 VN.n11 VN.t3 48.2268
R47 VN.n56 VN.t5 48.2268
R48 VN VN.n87 46.93
R49 VN.n36 VN.n1 42.5146
R50 VN.n80 VN.n45 42.5146
R51 VN.n36 VN.n35 38.6395
R52 VN.n80 VN.n79 38.6395
R53 VN.n15 VN.n14 25.0767
R54 VN.n28 VN.n27 25.0767
R55 VN.n60 VN.n59 25.0767
R56 VN.n73 VN.n72 25.0767
R57 VN.n14 VN.n9 24.5923
R58 VN.n16 VN.n7 24.5923
R59 VN.n20 VN.n7 24.5923
R60 VN.n23 VN.n22 24.5923
R61 VN.n23 VN.n5 24.5923
R62 VN.n30 VN.n28 24.5923
R63 VN.n34 VN.n3 24.5923
R64 VN.n35 VN.n34 24.5923
R65 VN.n40 VN.n1 24.5923
R66 VN.n41 VN.n40 24.5923
R67 VN.n59 VN.n54 24.5923
R68 VN.n68 VN.n50 24.5923
R69 VN.n68 VN.n67 24.5923
R70 VN.n65 VN.n52 24.5923
R71 VN.n61 VN.n52 24.5923
R72 VN.n79 VN.n78 24.5923
R73 VN.n78 VN.n47 24.5923
R74 VN.n74 VN.n73 24.5923
R75 VN.n85 VN.n84 24.5923
R76 VN.n84 VN.n45 24.5923
R77 VN.n10 VN.n9 21.1495
R78 VN.n30 VN.n29 21.1495
R79 VN.n55 VN.n54 21.1495
R80 VN.n74 VN.n49 21.1495
R81 VN.n10 VN.t4 14.0377
R82 VN.n21 VN.t8 14.0377
R83 VN.n29 VN.t0 14.0377
R84 VN.n42 VN.t7 14.0377
R85 VN.n55 VN.t1 14.0377
R86 VN.n66 VN.t9 14.0377
R87 VN.n49 VN.t2 14.0377
R88 VN.n86 VN.t6 14.0377
R89 VN.n21 VN.n20 12.2964
R90 VN.n22 VN.n21 12.2964
R91 VN.n67 VN.n66 12.2964
R92 VN.n66 VN.n65 12.2964
R93 VN.n42 VN.n41 5.4107
R94 VN.n86 VN.n85 5.4107
R95 VN.n57 VN.n56 4.94439
R96 VN.n12 VN.n11 4.94439
R97 VN.n29 VN.n3 3.44336
R98 VN.n49 VN.n47 3.44336
R99 VN.n87 VN.n44 0.278335
R100 VN.n43 VN.n0 0.278335
R101 VN.n83 VN.n44 0.189894
R102 VN.n83 VN.n82 0.189894
R103 VN.n82 VN.n81 0.189894
R104 VN.n81 VN.n46 0.189894
R105 VN.n77 VN.n46 0.189894
R106 VN.n77 VN.n76 0.189894
R107 VN.n76 VN.n75 0.189894
R108 VN.n75 VN.n48 0.189894
R109 VN.n71 VN.n48 0.189894
R110 VN.n71 VN.n70 0.189894
R111 VN.n70 VN.n69 0.189894
R112 VN.n69 VN.n51 0.189894
R113 VN.n64 VN.n51 0.189894
R114 VN.n64 VN.n63 0.189894
R115 VN.n63 VN.n62 0.189894
R116 VN.n62 VN.n53 0.189894
R117 VN.n58 VN.n53 0.189894
R118 VN.n58 VN.n57 0.189894
R119 VN.n13 VN.n12 0.189894
R120 VN.n13 VN.n8 0.189894
R121 VN.n17 VN.n8 0.189894
R122 VN.n18 VN.n17 0.189894
R123 VN.n19 VN.n18 0.189894
R124 VN.n19 VN.n6 0.189894
R125 VN.n24 VN.n6 0.189894
R126 VN.n25 VN.n24 0.189894
R127 VN.n26 VN.n25 0.189894
R128 VN.n26 VN.n4 0.189894
R129 VN.n31 VN.n4 0.189894
R130 VN.n32 VN.n31 0.189894
R131 VN.n33 VN.n32 0.189894
R132 VN.n33 VN.n2 0.189894
R133 VN.n37 VN.n2 0.189894
R134 VN.n38 VN.n37 0.189894
R135 VN.n39 VN.n38 0.189894
R136 VN.n39 VN.n0 0.189894
R137 VN VN.n43 0.153485
R138 VDD2.n1 VDD2.t2 131.034
R139 VDD2.n4 VDD2.t8 128.292
R140 VDD2.n3 VDD2.n2 118.365
R141 VDD2 VDD2.n7 118.362
R142 VDD2.n1 VDD2.n0 116.365
R143 VDD2.n6 VDD2.n5 116.365
R144 VDD2.n4 VDD2.n3 38.1679
R145 VDD2.n7 VDD2.t9 11.9282
R146 VDD2.n7 VDD2.t1 11.9282
R147 VDD2.n5 VDD2.t5 11.9282
R148 VDD2.n5 VDD2.t7 11.9282
R149 VDD2.n2 VDD2.t6 11.9282
R150 VDD2.n2 VDD2.t3 11.9282
R151 VDD2.n0 VDD2.t0 11.9282
R152 VDD2.n0 VDD2.t4 11.9282
R153 VDD2.n6 VDD2.n4 2.74188
R154 VDD2 VDD2.n6 0.744035
R155 VDD2.n3 VDD2.n1 0.630499
R156 VTAIL.n17 VTAIL.t12 111.614
R157 VTAIL.n2 VTAIL.t2 111.614
R158 VTAIL.n16 VTAIL.t6 111.614
R159 VTAIL.n11 VTAIL.t14 111.614
R160 VTAIL.n19 VTAIL.n18 99.6854
R161 VTAIL.n1 VTAIL.n0 99.6854
R162 VTAIL.n4 VTAIL.n3 99.6854
R163 VTAIL.n6 VTAIL.n5 99.6854
R164 VTAIL.n15 VTAIL.n14 99.6854
R165 VTAIL.n13 VTAIL.n12 99.6854
R166 VTAIL.n10 VTAIL.n9 99.6854
R167 VTAIL.n8 VTAIL.n7 99.6854
R168 VTAIL.n8 VTAIL.n6 19.2807
R169 VTAIL.n17 VTAIL.n16 16.5393
R170 VTAIL.n18 VTAIL.t11 11.9282
R171 VTAIL.n18 VTAIL.t19 11.9282
R172 VTAIL.n0 VTAIL.t16 11.9282
R173 VTAIL.n0 VTAIL.t15 11.9282
R174 VTAIL.n3 VTAIL.t0 11.9282
R175 VTAIL.n3 VTAIL.t3 11.9282
R176 VTAIL.n5 VTAIL.t1 11.9282
R177 VTAIL.n5 VTAIL.t4 11.9282
R178 VTAIL.n14 VTAIL.t9 11.9282
R179 VTAIL.n14 VTAIL.t8 11.9282
R180 VTAIL.n12 VTAIL.t7 11.9282
R181 VTAIL.n12 VTAIL.t5 11.9282
R182 VTAIL.n9 VTAIL.t10 11.9282
R183 VTAIL.n9 VTAIL.t18 11.9282
R184 VTAIL.n7 VTAIL.t13 11.9282
R185 VTAIL.n7 VTAIL.t17 11.9282
R186 VTAIL.n10 VTAIL.n8 2.74188
R187 VTAIL.n11 VTAIL.n10 2.74188
R188 VTAIL.n15 VTAIL.n13 2.74188
R189 VTAIL.n16 VTAIL.n15 2.74188
R190 VTAIL.n6 VTAIL.n4 2.74188
R191 VTAIL.n4 VTAIL.n2 2.74188
R192 VTAIL.n19 VTAIL.n17 2.74188
R193 VTAIL VTAIL.n1 2.11472
R194 VTAIL.n13 VTAIL.n11 1.84102
R195 VTAIL.n2 VTAIL.n1 1.84102
R196 VTAIL VTAIL.n19 0.627655
R197 B.n684 B.n683 585
R198 B.n198 B.n133 585
R199 B.n197 B.n196 585
R200 B.n195 B.n194 585
R201 B.n193 B.n192 585
R202 B.n191 B.n190 585
R203 B.n189 B.n188 585
R204 B.n187 B.n186 585
R205 B.n185 B.n184 585
R206 B.n183 B.n182 585
R207 B.n181 B.n180 585
R208 B.n178 B.n177 585
R209 B.n176 B.n175 585
R210 B.n174 B.n173 585
R211 B.n172 B.n171 585
R212 B.n170 B.n169 585
R213 B.n168 B.n167 585
R214 B.n166 B.n165 585
R215 B.n164 B.n163 585
R216 B.n162 B.n161 585
R217 B.n160 B.n159 585
R218 B.n157 B.n156 585
R219 B.n155 B.n154 585
R220 B.n153 B.n152 585
R221 B.n151 B.n150 585
R222 B.n149 B.n148 585
R223 B.n147 B.n146 585
R224 B.n145 B.n144 585
R225 B.n143 B.n142 585
R226 B.n141 B.n140 585
R227 B.n139 B.n138 585
R228 B.n116 B.n115 585
R229 B.n682 B.n117 585
R230 B.n687 B.n117 585
R231 B.n681 B.n680 585
R232 B.n680 B.n113 585
R233 B.n679 B.n112 585
R234 B.n693 B.n112 585
R235 B.n678 B.n111 585
R236 B.n694 B.n111 585
R237 B.n677 B.n110 585
R238 B.n695 B.n110 585
R239 B.n676 B.n675 585
R240 B.n675 B.n106 585
R241 B.n674 B.n105 585
R242 B.n701 B.n105 585
R243 B.n673 B.n104 585
R244 B.n702 B.n104 585
R245 B.n672 B.n103 585
R246 B.n703 B.n103 585
R247 B.n671 B.n670 585
R248 B.n670 B.n99 585
R249 B.n669 B.n98 585
R250 B.n709 B.n98 585
R251 B.n668 B.n97 585
R252 B.n710 B.n97 585
R253 B.n667 B.n96 585
R254 B.n711 B.n96 585
R255 B.n666 B.n665 585
R256 B.n665 B.n92 585
R257 B.n664 B.n91 585
R258 B.n717 B.n91 585
R259 B.n663 B.n90 585
R260 B.n718 B.n90 585
R261 B.n662 B.n89 585
R262 B.n719 B.n89 585
R263 B.n661 B.n660 585
R264 B.n660 B.n85 585
R265 B.n659 B.n84 585
R266 B.n725 B.n84 585
R267 B.n658 B.n83 585
R268 B.n726 B.n83 585
R269 B.n657 B.n82 585
R270 B.n727 B.n82 585
R271 B.n656 B.n655 585
R272 B.n655 B.n78 585
R273 B.n654 B.n77 585
R274 B.n733 B.n77 585
R275 B.n653 B.n76 585
R276 B.n734 B.n76 585
R277 B.n652 B.n75 585
R278 B.n735 B.n75 585
R279 B.n651 B.n650 585
R280 B.n650 B.n71 585
R281 B.n649 B.n70 585
R282 B.n741 B.n70 585
R283 B.n648 B.n69 585
R284 B.n742 B.n69 585
R285 B.n647 B.n68 585
R286 B.n743 B.n68 585
R287 B.n646 B.n645 585
R288 B.n645 B.n67 585
R289 B.n644 B.n63 585
R290 B.n749 B.n63 585
R291 B.n643 B.n62 585
R292 B.n750 B.n62 585
R293 B.n642 B.n61 585
R294 B.n751 B.n61 585
R295 B.n641 B.n640 585
R296 B.n640 B.n57 585
R297 B.n639 B.n56 585
R298 B.n757 B.n56 585
R299 B.n638 B.n55 585
R300 B.n758 B.n55 585
R301 B.n637 B.n54 585
R302 B.n759 B.n54 585
R303 B.n636 B.n635 585
R304 B.n635 B.n50 585
R305 B.n634 B.n49 585
R306 B.n765 B.n49 585
R307 B.n633 B.n48 585
R308 B.n766 B.n48 585
R309 B.n632 B.n47 585
R310 B.n767 B.n47 585
R311 B.n631 B.n630 585
R312 B.n630 B.n43 585
R313 B.n629 B.n42 585
R314 B.n773 B.n42 585
R315 B.n628 B.n41 585
R316 B.n774 B.n41 585
R317 B.n627 B.n40 585
R318 B.n775 B.n40 585
R319 B.n626 B.n625 585
R320 B.n625 B.n36 585
R321 B.n624 B.n35 585
R322 B.n781 B.n35 585
R323 B.n623 B.n34 585
R324 B.n782 B.n34 585
R325 B.n622 B.n33 585
R326 B.n783 B.n33 585
R327 B.n621 B.n620 585
R328 B.n620 B.n29 585
R329 B.n619 B.n28 585
R330 B.n789 B.n28 585
R331 B.n618 B.n27 585
R332 B.n790 B.n27 585
R333 B.n617 B.n26 585
R334 B.n791 B.n26 585
R335 B.n616 B.n615 585
R336 B.n615 B.n22 585
R337 B.n614 B.n21 585
R338 B.n797 B.n21 585
R339 B.n613 B.n20 585
R340 B.n798 B.n20 585
R341 B.n612 B.n19 585
R342 B.n799 B.n19 585
R343 B.n611 B.n610 585
R344 B.n610 B.n18 585
R345 B.n609 B.n14 585
R346 B.n805 B.n14 585
R347 B.n608 B.n13 585
R348 B.n806 B.n13 585
R349 B.n607 B.n12 585
R350 B.n807 B.n12 585
R351 B.n606 B.n605 585
R352 B.n605 B.n8 585
R353 B.n604 B.n7 585
R354 B.n813 B.n7 585
R355 B.n603 B.n6 585
R356 B.n814 B.n6 585
R357 B.n602 B.n5 585
R358 B.n815 B.n5 585
R359 B.n601 B.n600 585
R360 B.n600 B.n4 585
R361 B.n599 B.n199 585
R362 B.n599 B.n598 585
R363 B.n589 B.n200 585
R364 B.n201 B.n200 585
R365 B.n591 B.n590 585
R366 B.n592 B.n591 585
R367 B.n588 B.n206 585
R368 B.n206 B.n205 585
R369 B.n587 B.n586 585
R370 B.n586 B.n585 585
R371 B.n208 B.n207 585
R372 B.n578 B.n208 585
R373 B.n577 B.n576 585
R374 B.n579 B.n577 585
R375 B.n575 B.n213 585
R376 B.n213 B.n212 585
R377 B.n574 B.n573 585
R378 B.n573 B.n572 585
R379 B.n215 B.n214 585
R380 B.n216 B.n215 585
R381 B.n565 B.n564 585
R382 B.n566 B.n565 585
R383 B.n563 B.n221 585
R384 B.n221 B.n220 585
R385 B.n562 B.n561 585
R386 B.n561 B.n560 585
R387 B.n223 B.n222 585
R388 B.n224 B.n223 585
R389 B.n553 B.n552 585
R390 B.n554 B.n553 585
R391 B.n551 B.n229 585
R392 B.n229 B.n228 585
R393 B.n550 B.n549 585
R394 B.n549 B.n548 585
R395 B.n231 B.n230 585
R396 B.n232 B.n231 585
R397 B.n541 B.n540 585
R398 B.n542 B.n541 585
R399 B.n539 B.n237 585
R400 B.n237 B.n236 585
R401 B.n538 B.n537 585
R402 B.n537 B.n536 585
R403 B.n239 B.n238 585
R404 B.n240 B.n239 585
R405 B.n529 B.n528 585
R406 B.n530 B.n529 585
R407 B.n527 B.n244 585
R408 B.n248 B.n244 585
R409 B.n526 B.n525 585
R410 B.n525 B.n524 585
R411 B.n246 B.n245 585
R412 B.n247 B.n246 585
R413 B.n517 B.n516 585
R414 B.n518 B.n517 585
R415 B.n515 B.n253 585
R416 B.n253 B.n252 585
R417 B.n514 B.n513 585
R418 B.n513 B.n512 585
R419 B.n255 B.n254 585
R420 B.n256 B.n255 585
R421 B.n505 B.n504 585
R422 B.n506 B.n505 585
R423 B.n503 B.n261 585
R424 B.n261 B.n260 585
R425 B.n502 B.n501 585
R426 B.n501 B.n500 585
R427 B.n263 B.n262 585
R428 B.n493 B.n263 585
R429 B.n492 B.n491 585
R430 B.n494 B.n492 585
R431 B.n490 B.n268 585
R432 B.n268 B.n267 585
R433 B.n489 B.n488 585
R434 B.n488 B.n487 585
R435 B.n270 B.n269 585
R436 B.n271 B.n270 585
R437 B.n480 B.n479 585
R438 B.n481 B.n480 585
R439 B.n478 B.n276 585
R440 B.n276 B.n275 585
R441 B.n477 B.n476 585
R442 B.n476 B.n475 585
R443 B.n278 B.n277 585
R444 B.n279 B.n278 585
R445 B.n468 B.n467 585
R446 B.n469 B.n468 585
R447 B.n466 B.n284 585
R448 B.n284 B.n283 585
R449 B.n465 B.n464 585
R450 B.n464 B.n463 585
R451 B.n286 B.n285 585
R452 B.n287 B.n286 585
R453 B.n456 B.n455 585
R454 B.n457 B.n456 585
R455 B.n454 B.n292 585
R456 B.n292 B.n291 585
R457 B.n453 B.n452 585
R458 B.n452 B.n451 585
R459 B.n294 B.n293 585
R460 B.n295 B.n294 585
R461 B.n444 B.n443 585
R462 B.n445 B.n444 585
R463 B.n442 B.n300 585
R464 B.n300 B.n299 585
R465 B.n441 B.n440 585
R466 B.n440 B.n439 585
R467 B.n302 B.n301 585
R468 B.n303 B.n302 585
R469 B.n432 B.n431 585
R470 B.n433 B.n432 585
R471 B.n430 B.n307 585
R472 B.n311 B.n307 585
R473 B.n429 B.n428 585
R474 B.n428 B.n427 585
R475 B.n309 B.n308 585
R476 B.n310 B.n309 585
R477 B.n420 B.n419 585
R478 B.n421 B.n420 585
R479 B.n418 B.n316 585
R480 B.n316 B.n315 585
R481 B.n417 B.n416 585
R482 B.n416 B.n415 585
R483 B.n318 B.n317 585
R484 B.n319 B.n318 585
R485 B.n408 B.n407 585
R486 B.n409 B.n408 585
R487 B.n322 B.n321 585
R488 B.n347 B.n346 585
R489 B.n348 B.n344 585
R490 B.n344 B.n323 585
R491 B.n350 B.n349 585
R492 B.n352 B.n343 585
R493 B.n355 B.n354 585
R494 B.n356 B.n342 585
R495 B.n358 B.n357 585
R496 B.n360 B.n341 585
R497 B.n363 B.n362 585
R498 B.n364 B.n338 585
R499 B.n367 B.n366 585
R500 B.n369 B.n337 585
R501 B.n372 B.n371 585
R502 B.n373 B.n336 585
R503 B.n375 B.n374 585
R504 B.n377 B.n335 585
R505 B.n380 B.n379 585
R506 B.n381 B.n334 585
R507 B.n383 B.n382 585
R508 B.n385 B.n333 585
R509 B.n388 B.n387 585
R510 B.n389 B.n329 585
R511 B.n391 B.n390 585
R512 B.n393 B.n328 585
R513 B.n396 B.n395 585
R514 B.n397 B.n327 585
R515 B.n399 B.n398 585
R516 B.n401 B.n326 585
R517 B.n402 B.n325 585
R518 B.n405 B.n404 585
R519 B.n406 B.n324 585
R520 B.n324 B.n323 585
R521 B.n411 B.n410 585
R522 B.n410 B.n409 585
R523 B.n412 B.n320 585
R524 B.n320 B.n319 585
R525 B.n414 B.n413 585
R526 B.n415 B.n414 585
R527 B.n314 B.n313 585
R528 B.n315 B.n314 585
R529 B.n423 B.n422 585
R530 B.n422 B.n421 585
R531 B.n424 B.n312 585
R532 B.n312 B.n310 585
R533 B.n426 B.n425 585
R534 B.n427 B.n426 585
R535 B.n306 B.n305 585
R536 B.n311 B.n306 585
R537 B.n435 B.n434 585
R538 B.n434 B.n433 585
R539 B.n436 B.n304 585
R540 B.n304 B.n303 585
R541 B.n438 B.n437 585
R542 B.n439 B.n438 585
R543 B.n298 B.n297 585
R544 B.n299 B.n298 585
R545 B.n447 B.n446 585
R546 B.n446 B.n445 585
R547 B.n448 B.n296 585
R548 B.n296 B.n295 585
R549 B.n450 B.n449 585
R550 B.n451 B.n450 585
R551 B.n290 B.n289 585
R552 B.n291 B.n290 585
R553 B.n459 B.n458 585
R554 B.n458 B.n457 585
R555 B.n460 B.n288 585
R556 B.n288 B.n287 585
R557 B.n462 B.n461 585
R558 B.n463 B.n462 585
R559 B.n282 B.n281 585
R560 B.n283 B.n282 585
R561 B.n471 B.n470 585
R562 B.n470 B.n469 585
R563 B.n472 B.n280 585
R564 B.n280 B.n279 585
R565 B.n474 B.n473 585
R566 B.n475 B.n474 585
R567 B.n274 B.n273 585
R568 B.n275 B.n274 585
R569 B.n483 B.n482 585
R570 B.n482 B.n481 585
R571 B.n484 B.n272 585
R572 B.n272 B.n271 585
R573 B.n486 B.n485 585
R574 B.n487 B.n486 585
R575 B.n266 B.n265 585
R576 B.n267 B.n266 585
R577 B.n496 B.n495 585
R578 B.n495 B.n494 585
R579 B.n497 B.n264 585
R580 B.n493 B.n264 585
R581 B.n499 B.n498 585
R582 B.n500 B.n499 585
R583 B.n259 B.n258 585
R584 B.n260 B.n259 585
R585 B.n508 B.n507 585
R586 B.n507 B.n506 585
R587 B.n509 B.n257 585
R588 B.n257 B.n256 585
R589 B.n511 B.n510 585
R590 B.n512 B.n511 585
R591 B.n251 B.n250 585
R592 B.n252 B.n251 585
R593 B.n520 B.n519 585
R594 B.n519 B.n518 585
R595 B.n521 B.n249 585
R596 B.n249 B.n247 585
R597 B.n523 B.n522 585
R598 B.n524 B.n523 585
R599 B.n243 B.n242 585
R600 B.n248 B.n243 585
R601 B.n532 B.n531 585
R602 B.n531 B.n530 585
R603 B.n533 B.n241 585
R604 B.n241 B.n240 585
R605 B.n535 B.n534 585
R606 B.n536 B.n535 585
R607 B.n235 B.n234 585
R608 B.n236 B.n235 585
R609 B.n544 B.n543 585
R610 B.n543 B.n542 585
R611 B.n545 B.n233 585
R612 B.n233 B.n232 585
R613 B.n547 B.n546 585
R614 B.n548 B.n547 585
R615 B.n227 B.n226 585
R616 B.n228 B.n227 585
R617 B.n556 B.n555 585
R618 B.n555 B.n554 585
R619 B.n557 B.n225 585
R620 B.n225 B.n224 585
R621 B.n559 B.n558 585
R622 B.n560 B.n559 585
R623 B.n219 B.n218 585
R624 B.n220 B.n219 585
R625 B.n568 B.n567 585
R626 B.n567 B.n566 585
R627 B.n569 B.n217 585
R628 B.n217 B.n216 585
R629 B.n571 B.n570 585
R630 B.n572 B.n571 585
R631 B.n211 B.n210 585
R632 B.n212 B.n211 585
R633 B.n581 B.n580 585
R634 B.n580 B.n579 585
R635 B.n582 B.n209 585
R636 B.n578 B.n209 585
R637 B.n584 B.n583 585
R638 B.n585 B.n584 585
R639 B.n204 B.n203 585
R640 B.n205 B.n204 585
R641 B.n594 B.n593 585
R642 B.n593 B.n592 585
R643 B.n595 B.n202 585
R644 B.n202 B.n201 585
R645 B.n597 B.n596 585
R646 B.n598 B.n597 585
R647 B.n2 B.n0 585
R648 B.n4 B.n2 585
R649 B.n3 B.n1 585
R650 B.n814 B.n3 585
R651 B.n812 B.n811 585
R652 B.n813 B.n812 585
R653 B.n810 B.n9 585
R654 B.n9 B.n8 585
R655 B.n809 B.n808 585
R656 B.n808 B.n807 585
R657 B.n11 B.n10 585
R658 B.n806 B.n11 585
R659 B.n804 B.n803 585
R660 B.n805 B.n804 585
R661 B.n802 B.n15 585
R662 B.n18 B.n15 585
R663 B.n801 B.n800 585
R664 B.n800 B.n799 585
R665 B.n17 B.n16 585
R666 B.n798 B.n17 585
R667 B.n796 B.n795 585
R668 B.n797 B.n796 585
R669 B.n794 B.n23 585
R670 B.n23 B.n22 585
R671 B.n793 B.n792 585
R672 B.n792 B.n791 585
R673 B.n25 B.n24 585
R674 B.n790 B.n25 585
R675 B.n788 B.n787 585
R676 B.n789 B.n788 585
R677 B.n786 B.n30 585
R678 B.n30 B.n29 585
R679 B.n785 B.n784 585
R680 B.n784 B.n783 585
R681 B.n32 B.n31 585
R682 B.n782 B.n32 585
R683 B.n780 B.n779 585
R684 B.n781 B.n780 585
R685 B.n778 B.n37 585
R686 B.n37 B.n36 585
R687 B.n777 B.n776 585
R688 B.n776 B.n775 585
R689 B.n39 B.n38 585
R690 B.n774 B.n39 585
R691 B.n772 B.n771 585
R692 B.n773 B.n772 585
R693 B.n770 B.n44 585
R694 B.n44 B.n43 585
R695 B.n769 B.n768 585
R696 B.n768 B.n767 585
R697 B.n46 B.n45 585
R698 B.n766 B.n46 585
R699 B.n764 B.n763 585
R700 B.n765 B.n764 585
R701 B.n762 B.n51 585
R702 B.n51 B.n50 585
R703 B.n761 B.n760 585
R704 B.n760 B.n759 585
R705 B.n53 B.n52 585
R706 B.n758 B.n53 585
R707 B.n756 B.n755 585
R708 B.n757 B.n756 585
R709 B.n754 B.n58 585
R710 B.n58 B.n57 585
R711 B.n753 B.n752 585
R712 B.n752 B.n751 585
R713 B.n60 B.n59 585
R714 B.n750 B.n60 585
R715 B.n748 B.n747 585
R716 B.n749 B.n748 585
R717 B.n746 B.n64 585
R718 B.n67 B.n64 585
R719 B.n745 B.n744 585
R720 B.n744 B.n743 585
R721 B.n66 B.n65 585
R722 B.n742 B.n66 585
R723 B.n740 B.n739 585
R724 B.n741 B.n740 585
R725 B.n738 B.n72 585
R726 B.n72 B.n71 585
R727 B.n737 B.n736 585
R728 B.n736 B.n735 585
R729 B.n74 B.n73 585
R730 B.n734 B.n74 585
R731 B.n732 B.n731 585
R732 B.n733 B.n732 585
R733 B.n730 B.n79 585
R734 B.n79 B.n78 585
R735 B.n729 B.n728 585
R736 B.n728 B.n727 585
R737 B.n81 B.n80 585
R738 B.n726 B.n81 585
R739 B.n724 B.n723 585
R740 B.n725 B.n724 585
R741 B.n722 B.n86 585
R742 B.n86 B.n85 585
R743 B.n721 B.n720 585
R744 B.n720 B.n719 585
R745 B.n88 B.n87 585
R746 B.n718 B.n88 585
R747 B.n716 B.n715 585
R748 B.n717 B.n716 585
R749 B.n714 B.n93 585
R750 B.n93 B.n92 585
R751 B.n713 B.n712 585
R752 B.n712 B.n711 585
R753 B.n95 B.n94 585
R754 B.n710 B.n95 585
R755 B.n708 B.n707 585
R756 B.n709 B.n708 585
R757 B.n706 B.n100 585
R758 B.n100 B.n99 585
R759 B.n705 B.n704 585
R760 B.n704 B.n703 585
R761 B.n102 B.n101 585
R762 B.n702 B.n102 585
R763 B.n700 B.n699 585
R764 B.n701 B.n700 585
R765 B.n698 B.n107 585
R766 B.n107 B.n106 585
R767 B.n697 B.n696 585
R768 B.n696 B.n695 585
R769 B.n109 B.n108 585
R770 B.n694 B.n109 585
R771 B.n692 B.n691 585
R772 B.n693 B.n692 585
R773 B.n690 B.n114 585
R774 B.n114 B.n113 585
R775 B.n689 B.n688 585
R776 B.n688 B.n687 585
R777 B.n817 B.n816 585
R778 B.n816 B.n815 585
R779 B.n410 B.n322 535.745
R780 B.n688 B.n116 535.745
R781 B.n408 B.n324 535.745
R782 B.n684 B.n117 535.745
R783 B.n686 B.n685 256.663
R784 B.n686 B.n132 256.663
R785 B.n686 B.n131 256.663
R786 B.n686 B.n130 256.663
R787 B.n686 B.n129 256.663
R788 B.n686 B.n128 256.663
R789 B.n686 B.n127 256.663
R790 B.n686 B.n126 256.663
R791 B.n686 B.n125 256.663
R792 B.n686 B.n124 256.663
R793 B.n686 B.n123 256.663
R794 B.n686 B.n122 256.663
R795 B.n686 B.n121 256.663
R796 B.n686 B.n120 256.663
R797 B.n686 B.n119 256.663
R798 B.n686 B.n118 256.663
R799 B.n345 B.n323 256.663
R800 B.n351 B.n323 256.663
R801 B.n353 B.n323 256.663
R802 B.n359 B.n323 256.663
R803 B.n361 B.n323 256.663
R804 B.n368 B.n323 256.663
R805 B.n370 B.n323 256.663
R806 B.n376 B.n323 256.663
R807 B.n378 B.n323 256.663
R808 B.n384 B.n323 256.663
R809 B.n386 B.n323 256.663
R810 B.n392 B.n323 256.663
R811 B.n394 B.n323 256.663
R812 B.n400 B.n323 256.663
R813 B.n403 B.n323 256.663
R814 B.n330 B.t8 222.433
R815 B.n339 B.t4 222.433
R816 B.n136 B.t15 222.433
R817 B.n134 B.t11 222.433
R818 B.n409 B.n323 220.476
R819 B.n687 B.n686 220.476
R820 B.n330 B.t10 170.843
R821 B.n134 B.t13 170.843
R822 B.n339 B.t7 170.843
R823 B.n136 B.t16 170.843
R824 B.n410 B.n320 163.367
R825 B.n414 B.n320 163.367
R826 B.n414 B.n314 163.367
R827 B.n422 B.n314 163.367
R828 B.n422 B.n312 163.367
R829 B.n426 B.n312 163.367
R830 B.n426 B.n306 163.367
R831 B.n434 B.n306 163.367
R832 B.n434 B.n304 163.367
R833 B.n438 B.n304 163.367
R834 B.n438 B.n298 163.367
R835 B.n446 B.n298 163.367
R836 B.n446 B.n296 163.367
R837 B.n450 B.n296 163.367
R838 B.n450 B.n290 163.367
R839 B.n458 B.n290 163.367
R840 B.n458 B.n288 163.367
R841 B.n462 B.n288 163.367
R842 B.n462 B.n282 163.367
R843 B.n470 B.n282 163.367
R844 B.n470 B.n280 163.367
R845 B.n474 B.n280 163.367
R846 B.n474 B.n274 163.367
R847 B.n482 B.n274 163.367
R848 B.n482 B.n272 163.367
R849 B.n486 B.n272 163.367
R850 B.n486 B.n266 163.367
R851 B.n495 B.n266 163.367
R852 B.n495 B.n264 163.367
R853 B.n499 B.n264 163.367
R854 B.n499 B.n259 163.367
R855 B.n507 B.n259 163.367
R856 B.n507 B.n257 163.367
R857 B.n511 B.n257 163.367
R858 B.n511 B.n251 163.367
R859 B.n519 B.n251 163.367
R860 B.n519 B.n249 163.367
R861 B.n523 B.n249 163.367
R862 B.n523 B.n243 163.367
R863 B.n531 B.n243 163.367
R864 B.n531 B.n241 163.367
R865 B.n535 B.n241 163.367
R866 B.n535 B.n235 163.367
R867 B.n543 B.n235 163.367
R868 B.n543 B.n233 163.367
R869 B.n547 B.n233 163.367
R870 B.n547 B.n227 163.367
R871 B.n555 B.n227 163.367
R872 B.n555 B.n225 163.367
R873 B.n559 B.n225 163.367
R874 B.n559 B.n219 163.367
R875 B.n567 B.n219 163.367
R876 B.n567 B.n217 163.367
R877 B.n571 B.n217 163.367
R878 B.n571 B.n211 163.367
R879 B.n580 B.n211 163.367
R880 B.n580 B.n209 163.367
R881 B.n584 B.n209 163.367
R882 B.n584 B.n204 163.367
R883 B.n593 B.n204 163.367
R884 B.n593 B.n202 163.367
R885 B.n597 B.n202 163.367
R886 B.n597 B.n2 163.367
R887 B.n816 B.n2 163.367
R888 B.n816 B.n3 163.367
R889 B.n812 B.n3 163.367
R890 B.n812 B.n9 163.367
R891 B.n808 B.n9 163.367
R892 B.n808 B.n11 163.367
R893 B.n804 B.n11 163.367
R894 B.n804 B.n15 163.367
R895 B.n800 B.n15 163.367
R896 B.n800 B.n17 163.367
R897 B.n796 B.n17 163.367
R898 B.n796 B.n23 163.367
R899 B.n792 B.n23 163.367
R900 B.n792 B.n25 163.367
R901 B.n788 B.n25 163.367
R902 B.n788 B.n30 163.367
R903 B.n784 B.n30 163.367
R904 B.n784 B.n32 163.367
R905 B.n780 B.n32 163.367
R906 B.n780 B.n37 163.367
R907 B.n776 B.n37 163.367
R908 B.n776 B.n39 163.367
R909 B.n772 B.n39 163.367
R910 B.n772 B.n44 163.367
R911 B.n768 B.n44 163.367
R912 B.n768 B.n46 163.367
R913 B.n764 B.n46 163.367
R914 B.n764 B.n51 163.367
R915 B.n760 B.n51 163.367
R916 B.n760 B.n53 163.367
R917 B.n756 B.n53 163.367
R918 B.n756 B.n58 163.367
R919 B.n752 B.n58 163.367
R920 B.n752 B.n60 163.367
R921 B.n748 B.n60 163.367
R922 B.n748 B.n64 163.367
R923 B.n744 B.n64 163.367
R924 B.n744 B.n66 163.367
R925 B.n740 B.n66 163.367
R926 B.n740 B.n72 163.367
R927 B.n736 B.n72 163.367
R928 B.n736 B.n74 163.367
R929 B.n732 B.n74 163.367
R930 B.n732 B.n79 163.367
R931 B.n728 B.n79 163.367
R932 B.n728 B.n81 163.367
R933 B.n724 B.n81 163.367
R934 B.n724 B.n86 163.367
R935 B.n720 B.n86 163.367
R936 B.n720 B.n88 163.367
R937 B.n716 B.n88 163.367
R938 B.n716 B.n93 163.367
R939 B.n712 B.n93 163.367
R940 B.n712 B.n95 163.367
R941 B.n708 B.n95 163.367
R942 B.n708 B.n100 163.367
R943 B.n704 B.n100 163.367
R944 B.n704 B.n102 163.367
R945 B.n700 B.n102 163.367
R946 B.n700 B.n107 163.367
R947 B.n696 B.n107 163.367
R948 B.n696 B.n109 163.367
R949 B.n692 B.n109 163.367
R950 B.n692 B.n114 163.367
R951 B.n688 B.n114 163.367
R952 B.n346 B.n344 163.367
R953 B.n350 B.n344 163.367
R954 B.n354 B.n352 163.367
R955 B.n358 B.n342 163.367
R956 B.n362 B.n360 163.367
R957 B.n367 B.n338 163.367
R958 B.n371 B.n369 163.367
R959 B.n375 B.n336 163.367
R960 B.n379 B.n377 163.367
R961 B.n383 B.n334 163.367
R962 B.n387 B.n385 163.367
R963 B.n391 B.n329 163.367
R964 B.n395 B.n393 163.367
R965 B.n399 B.n327 163.367
R966 B.n402 B.n401 163.367
R967 B.n404 B.n324 163.367
R968 B.n408 B.n318 163.367
R969 B.n416 B.n318 163.367
R970 B.n416 B.n316 163.367
R971 B.n420 B.n316 163.367
R972 B.n420 B.n309 163.367
R973 B.n428 B.n309 163.367
R974 B.n428 B.n307 163.367
R975 B.n432 B.n307 163.367
R976 B.n432 B.n302 163.367
R977 B.n440 B.n302 163.367
R978 B.n440 B.n300 163.367
R979 B.n444 B.n300 163.367
R980 B.n444 B.n294 163.367
R981 B.n452 B.n294 163.367
R982 B.n452 B.n292 163.367
R983 B.n456 B.n292 163.367
R984 B.n456 B.n286 163.367
R985 B.n464 B.n286 163.367
R986 B.n464 B.n284 163.367
R987 B.n468 B.n284 163.367
R988 B.n468 B.n278 163.367
R989 B.n476 B.n278 163.367
R990 B.n476 B.n276 163.367
R991 B.n480 B.n276 163.367
R992 B.n480 B.n270 163.367
R993 B.n488 B.n270 163.367
R994 B.n488 B.n268 163.367
R995 B.n492 B.n268 163.367
R996 B.n492 B.n263 163.367
R997 B.n501 B.n263 163.367
R998 B.n501 B.n261 163.367
R999 B.n505 B.n261 163.367
R1000 B.n505 B.n255 163.367
R1001 B.n513 B.n255 163.367
R1002 B.n513 B.n253 163.367
R1003 B.n517 B.n253 163.367
R1004 B.n517 B.n246 163.367
R1005 B.n525 B.n246 163.367
R1006 B.n525 B.n244 163.367
R1007 B.n529 B.n244 163.367
R1008 B.n529 B.n239 163.367
R1009 B.n537 B.n239 163.367
R1010 B.n537 B.n237 163.367
R1011 B.n541 B.n237 163.367
R1012 B.n541 B.n231 163.367
R1013 B.n549 B.n231 163.367
R1014 B.n549 B.n229 163.367
R1015 B.n553 B.n229 163.367
R1016 B.n553 B.n223 163.367
R1017 B.n561 B.n223 163.367
R1018 B.n561 B.n221 163.367
R1019 B.n565 B.n221 163.367
R1020 B.n565 B.n215 163.367
R1021 B.n573 B.n215 163.367
R1022 B.n573 B.n213 163.367
R1023 B.n577 B.n213 163.367
R1024 B.n577 B.n208 163.367
R1025 B.n586 B.n208 163.367
R1026 B.n586 B.n206 163.367
R1027 B.n591 B.n206 163.367
R1028 B.n591 B.n200 163.367
R1029 B.n599 B.n200 163.367
R1030 B.n600 B.n599 163.367
R1031 B.n600 B.n5 163.367
R1032 B.n6 B.n5 163.367
R1033 B.n7 B.n6 163.367
R1034 B.n605 B.n7 163.367
R1035 B.n605 B.n12 163.367
R1036 B.n13 B.n12 163.367
R1037 B.n14 B.n13 163.367
R1038 B.n610 B.n14 163.367
R1039 B.n610 B.n19 163.367
R1040 B.n20 B.n19 163.367
R1041 B.n21 B.n20 163.367
R1042 B.n615 B.n21 163.367
R1043 B.n615 B.n26 163.367
R1044 B.n27 B.n26 163.367
R1045 B.n28 B.n27 163.367
R1046 B.n620 B.n28 163.367
R1047 B.n620 B.n33 163.367
R1048 B.n34 B.n33 163.367
R1049 B.n35 B.n34 163.367
R1050 B.n625 B.n35 163.367
R1051 B.n625 B.n40 163.367
R1052 B.n41 B.n40 163.367
R1053 B.n42 B.n41 163.367
R1054 B.n630 B.n42 163.367
R1055 B.n630 B.n47 163.367
R1056 B.n48 B.n47 163.367
R1057 B.n49 B.n48 163.367
R1058 B.n635 B.n49 163.367
R1059 B.n635 B.n54 163.367
R1060 B.n55 B.n54 163.367
R1061 B.n56 B.n55 163.367
R1062 B.n640 B.n56 163.367
R1063 B.n640 B.n61 163.367
R1064 B.n62 B.n61 163.367
R1065 B.n63 B.n62 163.367
R1066 B.n645 B.n63 163.367
R1067 B.n645 B.n68 163.367
R1068 B.n69 B.n68 163.367
R1069 B.n70 B.n69 163.367
R1070 B.n650 B.n70 163.367
R1071 B.n650 B.n75 163.367
R1072 B.n76 B.n75 163.367
R1073 B.n77 B.n76 163.367
R1074 B.n655 B.n77 163.367
R1075 B.n655 B.n82 163.367
R1076 B.n83 B.n82 163.367
R1077 B.n84 B.n83 163.367
R1078 B.n660 B.n84 163.367
R1079 B.n660 B.n89 163.367
R1080 B.n90 B.n89 163.367
R1081 B.n91 B.n90 163.367
R1082 B.n665 B.n91 163.367
R1083 B.n665 B.n96 163.367
R1084 B.n97 B.n96 163.367
R1085 B.n98 B.n97 163.367
R1086 B.n670 B.n98 163.367
R1087 B.n670 B.n103 163.367
R1088 B.n104 B.n103 163.367
R1089 B.n105 B.n104 163.367
R1090 B.n675 B.n105 163.367
R1091 B.n675 B.n110 163.367
R1092 B.n111 B.n110 163.367
R1093 B.n112 B.n111 163.367
R1094 B.n680 B.n112 163.367
R1095 B.n680 B.n117 163.367
R1096 B.n140 B.n139 163.367
R1097 B.n144 B.n143 163.367
R1098 B.n148 B.n147 163.367
R1099 B.n152 B.n151 163.367
R1100 B.n156 B.n155 163.367
R1101 B.n161 B.n160 163.367
R1102 B.n165 B.n164 163.367
R1103 B.n169 B.n168 163.367
R1104 B.n173 B.n172 163.367
R1105 B.n177 B.n176 163.367
R1106 B.n182 B.n181 163.367
R1107 B.n186 B.n185 163.367
R1108 B.n190 B.n189 163.367
R1109 B.n194 B.n193 163.367
R1110 B.n196 B.n133 163.367
R1111 B.n331 B.t9 109.171
R1112 B.n135 B.t14 109.171
R1113 B.n340 B.t6 109.169
R1114 B.n137 B.t17 109.169
R1115 B.n409 B.n319 107.859
R1116 B.n415 B.n319 107.859
R1117 B.n415 B.n315 107.859
R1118 B.n421 B.n315 107.859
R1119 B.n421 B.n310 107.859
R1120 B.n427 B.n310 107.859
R1121 B.n427 B.n311 107.859
R1122 B.n433 B.n303 107.859
R1123 B.n439 B.n303 107.859
R1124 B.n439 B.n299 107.859
R1125 B.n445 B.n299 107.859
R1126 B.n445 B.n295 107.859
R1127 B.n451 B.n295 107.859
R1128 B.n451 B.n291 107.859
R1129 B.n457 B.n291 107.859
R1130 B.n457 B.n287 107.859
R1131 B.n463 B.n287 107.859
R1132 B.n463 B.n283 107.859
R1133 B.n469 B.n283 107.859
R1134 B.n475 B.n279 107.859
R1135 B.n475 B.n275 107.859
R1136 B.n481 B.n275 107.859
R1137 B.n481 B.n271 107.859
R1138 B.n487 B.n271 107.859
R1139 B.n487 B.n267 107.859
R1140 B.n494 B.n267 107.859
R1141 B.n494 B.n493 107.859
R1142 B.n500 B.n260 107.859
R1143 B.n506 B.n260 107.859
R1144 B.n506 B.n256 107.859
R1145 B.n512 B.n256 107.859
R1146 B.n512 B.n252 107.859
R1147 B.n518 B.n252 107.859
R1148 B.n518 B.n247 107.859
R1149 B.n524 B.n247 107.859
R1150 B.n524 B.n248 107.859
R1151 B.n530 B.n240 107.859
R1152 B.n536 B.n240 107.859
R1153 B.n536 B.n236 107.859
R1154 B.n542 B.n236 107.859
R1155 B.n542 B.n232 107.859
R1156 B.n548 B.n232 107.859
R1157 B.n548 B.n228 107.859
R1158 B.n554 B.n228 107.859
R1159 B.n560 B.n224 107.859
R1160 B.n560 B.n220 107.859
R1161 B.n566 B.n220 107.859
R1162 B.n566 B.n216 107.859
R1163 B.n572 B.n216 107.859
R1164 B.n572 B.n212 107.859
R1165 B.n579 B.n212 107.859
R1166 B.n579 B.n578 107.859
R1167 B.n585 B.n205 107.859
R1168 B.n592 B.n205 107.859
R1169 B.n592 B.n201 107.859
R1170 B.n598 B.n201 107.859
R1171 B.n598 B.n4 107.859
R1172 B.n815 B.n4 107.859
R1173 B.n815 B.n814 107.859
R1174 B.n814 B.n813 107.859
R1175 B.n813 B.n8 107.859
R1176 B.n807 B.n8 107.859
R1177 B.n807 B.n806 107.859
R1178 B.n806 B.n805 107.859
R1179 B.n799 B.n18 107.859
R1180 B.n799 B.n798 107.859
R1181 B.n798 B.n797 107.859
R1182 B.n797 B.n22 107.859
R1183 B.n791 B.n22 107.859
R1184 B.n791 B.n790 107.859
R1185 B.n790 B.n789 107.859
R1186 B.n789 B.n29 107.859
R1187 B.n783 B.n782 107.859
R1188 B.n782 B.n781 107.859
R1189 B.n781 B.n36 107.859
R1190 B.n775 B.n36 107.859
R1191 B.n775 B.n774 107.859
R1192 B.n774 B.n773 107.859
R1193 B.n773 B.n43 107.859
R1194 B.n767 B.n43 107.859
R1195 B.n766 B.n765 107.859
R1196 B.n765 B.n50 107.859
R1197 B.n759 B.n50 107.859
R1198 B.n759 B.n758 107.859
R1199 B.n758 B.n757 107.859
R1200 B.n757 B.n57 107.859
R1201 B.n751 B.n57 107.859
R1202 B.n751 B.n750 107.859
R1203 B.n750 B.n749 107.859
R1204 B.n743 B.n67 107.859
R1205 B.n743 B.n742 107.859
R1206 B.n742 B.n741 107.859
R1207 B.n741 B.n71 107.859
R1208 B.n735 B.n71 107.859
R1209 B.n735 B.n734 107.859
R1210 B.n734 B.n733 107.859
R1211 B.n733 B.n78 107.859
R1212 B.n727 B.n726 107.859
R1213 B.n726 B.n725 107.859
R1214 B.n725 B.n85 107.859
R1215 B.n719 B.n85 107.859
R1216 B.n719 B.n718 107.859
R1217 B.n718 B.n717 107.859
R1218 B.n717 B.n92 107.859
R1219 B.n711 B.n92 107.859
R1220 B.n711 B.n710 107.859
R1221 B.n710 B.n709 107.859
R1222 B.n709 B.n99 107.859
R1223 B.n703 B.n99 107.859
R1224 B.n702 B.n701 107.859
R1225 B.n701 B.n106 107.859
R1226 B.n695 B.n106 107.859
R1227 B.n695 B.n694 107.859
R1228 B.n694 B.n693 107.859
R1229 B.n693 B.n113 107.859
R1230 B.n687 B.n113 107.859
R1231 B.n530 B.t0 106.273
R1232 B.n767 B.t23 106.273
R1233 B.n311 B.t5 80.8945
R1234 B.t12 B.n702 80.8945
R1235 B.n578 B.t2 77.7222
R1236 B.n18 B.t21 77.7222
R1237 B.t1 B.n279 74.5499
R1238 B.t20 B.n78 74.5499
R1239 B.n345 B.n322 71.676
R1240 B.n351 B.n350 71.676
R1241 B.n354 B.n353 71.676
R1242 B.n359 B.n358 71.676
R1243 B.n362 B.n361 71.676
R1244 B.n368 B.n367 71.676
R1245 B.n371 B.n370 71.676
R1246 B.n376 B.n375 71.676
R1247 B.n379 B.n378 71.676
R1248 B.n384 B.n383 71.676
R1249 B.n387 B.n386 71.676
R1250 B.n392 B.n391 71.676
R1251 B.n395 B.n394 71.676
R1252 B.n400 B.n399 71.676
R1253 B.n403 B.n402 71.676
R1254 B.n118 B.n116 71.676
R1255 B.n140 B.n119 71.676
R1256 B.n144 B.n120 71.676
R1257 B.n148 B.n121 71.676
R1258 B.n152 B.n122 71.676
R1259 B.n156 B.n123 71.676
R1260 B.n161 B.n124 71.676
R1261 B.n165 B.n125 71.676
R1262 B.n169 B.n126 71.676
R1263 B.n173 B.n127 71.676
R1264 B.n177 B.n128 71.676
R1265 B.n182 B.n129 71.676
R1266 B.n186 B.n130 71.676
R1267 B.n190 B.n131 71.676
R1268 B.n194 B.n132 71.676
R1269 B.n685 B.n133 71.676
R1270 B.n685 B.n684 71.676
R1271 B.n196 B.n132 71.676
R1272 B.n193 B.n131 71.676
R1273 B.n189 B.n130 71.676
R1274 B.n185 B.n129 71.676
R1275 B.n181 B.n128 71.676
R1276 B.n176 B.n127 71.676
R1277 B.n172 B.n126 71.676
R1278 B.n168 B.n125 71.676
R1279 B.n164 B.n124 71.676
R1280 B.n160 B.n123 71.676
R1281 B.n155 B.n122 71.676
R1282 B.n151 B.n121 71.676
R1283 B.n147 B.n120 71.676
R1284 B.n143 B.n119 71.676
R1285 B.n139 B.n118 71.676
R1286 B.n346 B.n345 71.676
R1287 B.n352 B.n351 71.676
R1288 B.n353 B.n342 71.676
R1289 B.n360 B.n359 71.676
R1290 B.n361 B.n338 71.676
R1291 B.n369 B.n368 71.676
R1292 B.n370 B.n336 71.676
R1293 B.n377 B.n376 71.676
R1294 B.n378 B.n334 71.676
R1295 B.n385 B.n384 71.676
R1296 B.n386 B.n329 71.676
R1297 B.n393 B.n392 71.676
R1298 B.n394 B.n327 71.676
R1299 B.n401 B.n400 71.676
R1300 B.n404 B.n403 71.676
R1301 B.n493 B.t18 71.3776
R1302 B.n67 B.t22 71.3776
R1303 B.t3 B.n224 68.2053
R1304 B.t19 B.n29 68.2053
R1305 B.n331 B.n330 61.6732
R1306 B.n340 B.n339 61.6732
R1307 B.n137 B.n136 61.6732
R1308 B.n135 B.n134 61.6732
R1309 B.n332 B.n331 59.5399
R1310 B.n365 B.n340 59.5399
R1311 B.n158 B.n137 59.5399
R1312 B.n179 B.n135 59.5399
R1313 B.n554 B.t3 39.6544
R1314 B.n783 B.t19 39.6544
R1315 B.n500 B.t18 36.4821
R1316 B.n749 B.t22 36.4821
R1317 B.n689 B.n115 34.8103
R1318 B.n683 B.n682 34.8103
R1319 B.n407 B.n406 34.8103
R1320 B.n411 B.n321 34.8103
R1321 B.n469 B.t1 33.3098
R1322 B.n727 B.t20 33.3098
R1323 B.n585 B.t2 30.1375
R1324 B.n805 B.t21 30.1375
R1325 B.n433 B.t5 26.9652
R1326 B.n703 B.t12 26.9652
R1327 B B.n817 18.0485
R1328 B.n138 B.n115 10.6151
R1329 B.n141 B.n138 10.6151
R1330 B.n142 B.n141 10.6151
R1331 B.n145 B.n142 10.6151
R1332 B.n146 B.n145 10.6151
R1333 B.n149 B.n146 10.6151
R1334 B.n150 B.n149 10.6151
R1335 B.n153 B.n150 10.6151
R1336 B.n154 B.n153 10.6151
R1337 B.n157 B.n154 10.6151
R1338 B.n162 B.n159 10.6151
R1339 B.n163 B.n162 10.6151
R1340 B.n166 B.n163 10.6151
R1341 B.n167 B.n166 10.6151
R1342 B.n170 B.n167 10.6151
R1343 B.n171 B.n170 10.6151
R1344 B.n174 B.n171 10.6151
R1345 B.n175 B.n174 10.6151
R1346 B.n178 B.n175 10.6151
R1347 B.n183 B.n180 10.6151
R1348 B.n184 B.n183 10.6151
R1349 B.n187 B.n184 10.6151
R1350 B.n188 B.n187 10.6151
R1351 B.n191 B.n188 10.6151
R1352 B.n192 B.n191 10.6151
R1353 B.n195 B.n192 10.6151
R1354 B.n197 B.n195 10.6151
R1355 B.n198 B.n197 10.6151
R1356 B.n683 B.n198 10.6151
R1357 B.n407 B.n317 10.6151
R1358 B.n417 B.n317 10.6151
R1359 B.n418 B.n417 10.6151
R1360 B.n419 B.n418 10.6151
R1361 B.n419 B.n308 10.6151
R1362 B.n429 B.n308 10.6151
R1363 B.n430 B.n429 10.6151
R1364 B.n431 B.n430 10.6151
R1365 B.n431 B.n301 10.6151
R1366 B.n441 B.n301 10.6151
R1367 B.n442 B.n441 10.6151
R1368 B.n443 B.n442 10.6151
R1369 B.n443 B.n293 10.6151
R1370 B.n453 B.n293 10.6151
R1371 B.n454 B.n453 10.6151
R1372 B.n455 B.n454 10.6151
R1373 B.n455 B.n285 10.6151
R1374 B.n465 B.n285 10.6151
R1375 B.n466 B.n465 10.6151
R1376 B.n467 B.n466 10.6151
R1377 B.n467 B.n277 10.6151
R1378 B.n477 B.n277 10.6151
R1379 B.n478 B.n477 10.6151
R1380 B.n479 B.n478 10.6151
R1381 B.n479 B.n269 10.6151
R1382 B.n489 B.n269 10.6151
R1383 B.n490 B.n489 10.6151
R1384 B.n491 B.n490 10.6151
R1385 B.n491 B.n262 10.6151
R1386 B.n502 B.n262 10.6151
R1387 B.n503 B.n502 10.6151
R1388 B.n504 B.n503 10.6151
R1389 B.n504 B.n254 10.6151
R1390 B.n514 B.n254 10.6151
R1391 B.n515 B.n514 10.6151
R1392 B.n516 B.n515 10.6151
R1393 B.n516 B.n245 10.6151
R1394 B.n526 B.n245 10.6151
R1395 B.n527 B.n526 10.6151
R1396 B.n528 B.n527 10.6151
R1397 B.n528 B.n238 10.6151
R1398 B.n538 B.n238 10.6151
R1399 B.n539 B.n538 10.6151
R1400 B.n540 B.n539 10.6151
R1401 B.n540 B.n230 10.6151
R1402 B.n550 B.n230 10.6151
R1403 B.n551 B.n550 10.6151
R1404 B.n552 B.n551 10.6151
R1405 B.n552 B.n222 10.6151
R1406 B.n562 B.n222 10.6151
R1407 B.n563 B.n562 10.6151
R1408 B.n564 B.n563 10.6151
R1409 B.n564 B.n214 10.6151
R1410 B.n574 B.n214 10.6151
R1411 B.n575 B.n574 10.6151
R1412 B.n576 B.n575 10.6151
R1413 B.n576 B.n207 10.6151
R1414 B.n587 B.n207 10.6151
R1415 B.n588 B.n587 10.6151
R1416 B.n590 B.n588 10.6151
R1417 B.n590 B.n589 10.6151
R1418 B.n589 B.n199 10.6151
R1419 B.n601 B.n199 10.6151
R1420 B.n602 B.n601 10.6151
R1421 B.n603 B.n602 10.6151
R1422 B.n604 B.n603 10.6151
R1423 B.n606 B.n604 10.6151
R1424 B.n607 B.n606 10.6151
R1425 B.n608 B.n607 10.6151
R1426 B.n609 B.n608 10.6151
R1427 B.n611 B.n609 10.6151
R1428 B.n612 B.n611 10.6151
R1429 B.n613 B.n612 10.6151
R1430 B.n614 B.n613 10.6151
R1431 B.n616 B.n614 10.6151
R1432 B.n617 B.n616 10.6151
R1433 B.n618 B.n617 10.6151
R1434 B.n619 B.n618 10.6151
R1435 B.n621 B.n619 10.6151
R1436 B.n622 B.n621 10.6151
R1437 B.n623 B.n622 10.6151
R1438 B.n624 B.n623 10.6151
R1439 B.n626 B.n624 10.6151
R1440 B.n627 B.n626 10.6151
R1441 B.n628 B.n627 10.6151
R1442 B.n629 B.n628 10.6151
R1443 B.n631 B.n629 10.6151
R1444 B.n632 B.n631 10.6151
R1445 B.n633 B.n632 10.6151
R1446 B.n634 B.n633 10.6151
R1447 B.n636 B.n634 10.6151
R1448 B.n637 B.n636 10.6151
R1449 B.n638 B.n637 10.6151
R1450 B.n639 B.n638 10.6151
R1451 B.n641 B.n639 10.6151
R1452 B.n642 B.n641 10.6151
R1453 B.n643 B.n642 10.6151
R1454 B.n644 B.n643 10.6151
R1455 B.n646 B.n644 10.6151
R1456 B.n647 B.n646 10.6151
R1457 B.n648 B.n647 10.6151
R1458 B.n649 B.n648 10.6151
R1459 B.n651 B.n649 10.6151
R1460 B.n652 B.n651 10.6151
R1461 B.n653 B.n652 10.6151
R1462 B.n654 B.n653 10.6151
R1463 B.n656 B.n654 10.6151
R1464 B.n657 B.n656 10.6151
R1465 B.n658 B.n657 10.6151
R1466 B.n659 B.n658 10.6151
R1467 B.n661 B.n659 10.6151
R1468 B.n662 B.n661 10.6151
R1469 B.n663 B.n662 10.6151
R1470 B.n664 B.n663 10.6151
R1471 B.n666 B.n664 10.6151
R1472 B.n667 B.n666 10.6151
R1473 B.n668 B.n667 10.6151
R1474 B.n669 B.n668 10.6151
R1475 B.n671 B.n669 10.6151
R1476 B.n672 B.n671 10.6151
R1477 B.n673 B.n672 10.6151
R1478 B.n674 B.n673 10.6151
R1479 B.n676 B.n674 10.6151
R1480 B.n677 B.n676 10.6151
R1481 B.n678 B.n677 10.6151
R1482 B.n679 B.n678 10.6151
R1483 B.n681 B.n679 10.6151
R1484 B.n682 B.n681 10.6151
R1485 B.n347 B.n321 10.6151
R1486 B.n348 B.n347 10.6151
R1487 B.n349 B.n348 10.6151
R1488 B.n349 B.n343 10.6151
R1489 B.n355 B.n343 10.6151
R1490 B.n356 B.n355 10.6151
R1491 B.n357 B.n356 10.6151
R1492 B.n357 B.n341 10.6151
R1493 B.n363 B.n341 10.6151
R1494 B.n364 B.n363 10.6151
R1495 B.n366 B.n337 10.6151
R1496 B.n372 B.n337 10.6151
R1497 B.n373 B.n372 10.6151
R1498 B.n374 B.n373 10.6151
R1499 B.n374 B.n335 10.6151
R1500 B.n380 B.n335 10.6151
R1501 B.n381 B.n380 10.6151
R1502 B.n382 B.n381 10.6151
R1503 B.n382 B.n333 10.6151
R1504 B.n389 B.n388 10.6151
R1505 B.n390 B.n389 10.6151
R1506 B.n390 B.n328 10.6151
R1507 B.n396 B.n328 10.6151
R1508 B.n397 B.n396 10.6151
R1509 B.n398 B.n397 10.6151
R1510 B.n398 B.n326 10.6151
R1511 B.n326 B.n325 10.6151
R1512 B.n405 B.n325 10.6151
R1513 B.n406 B.n405 10.6151
R1514 B.n412 B.n411 10.6151
R1515 B.n413 B.n412 10.6151
R1516 B.n413 B.n313 10.6151
R1517 B.n423 B.n313 10.6151
R1518 B.n424 B.n423 10.6151
R1519 B.n425 B.n424 10.6151
R1520 B.n425 B.n305 10.6151
R1521 B.n435 B.n305 10.6151
R1522 B.n436 B.n435 10.6151
R1523 B.n437 B.n436 10.6151
R1524 B.n437 B.n297 10.6151
R1525 B.n447 B.n297 10.6151
R1526 B.n448 B.n447 10.6151
R1527 B.n449 B.n448 10.6151
R1528 B.n449 B.n289 10.6151
R1529 B.n459 B.n289 10.6151
R1530 B.n460 B.n459 10.6151
R1531 B.n461 B.n460 10.6151
R1532 B.n461 B.n281 10.6151
R1533 B.n471 B.n281 10.6151
R1534 B.n472 B.n471 10.6151
R1535 B.n473 B.n472 10.6151
R1536 B.n473 B.n273 10.6151
R1537 B.n483 B.n273 10.6151
R1538 B.n484 B.n483 10.6151
R1539 B.n485 B.n484 10.6151
R1540 B.n485 B.n265 10.6151
R1541 B.n496 B.n265 10.6151
R1542 B.n497 B.n496 10.6151
R1543 B.n498 B.n497 10.6151
R1544 B.n498 B.n258 10.6151
R1545 B.n508 B.n258 10.6151
R1546 B.n509 B.n508 10.6151
R1547 B.n510 B.n509 10.6151
R1548 B.n510 B.n250 10.6151
R1549 B.n520 B.n250 10.6151
R1550 B.n521 B.n520 10.6151
R1551 B.n522 B.n521 10.6151
R1552 B.n522 B.n242 10.6151
R1553 B.n532 B.n242 10.6151
R1554 B.n533 B.n532 10.6151
R1555 B.n534 B.n533 10.6151
R1556 B.n534 B.n234 10.6151
R1557 B.n544 B.n234 10.6151
R1558 B.n545 B.n544 10.6151
R1559 B.n546 B.n545 10.6151
R1560 B.n546 B.n226 10.6151
R1561 B.n556 B.n226 10.6151
R1562 B.n557 B.n556 10.6151
R1563 B.n558 B.n557 10.6151
R1564 B.n558 B.n218 10.6151
R1565 B.n568 B.n218 10.6151
R1566 B.n569 B.n568 10.6151
R1567 B.n570 B.n569 10.6151
R1568 B.n570 B.n210 10.6151
R1569 B.n581 B.n210 10.6151
R1570 B.n582 B.n581 10.6151
R1571 B.n583 B.n582 10.6151
R1572 B.n583 B.n203 10.6151
R1573 B.n594 B.n203 10.6151
R1574 B.n595 B.n594 10.6151
R1575 B.n596 B.n595 10.6151
R1576 B.n596 B.n0 10.6151
R1577 B.n811 B.n1 10.6151
R1578 B.n811 B.n810 10.6151
R1579 B.n810 B.n809 10.6151
R1580 B.n809 B.n10 10.6151
R1581 B.n803 B.n10 10.6151
R1582 B.n803 B.n802 10.6151
R1583 B.n802 B.n801 10.6151
R1584 B.n801 B.n16 10.6151
R1585 B.n795 B.n16 10.6151
R1586 B.n795 B.n794 10.6151
R1587 B.n794 B.n793 10.6151
R1588 B.n793 B.n24 10.6151
R1589 B.n787 B.n24 10.6151
R1590 B.n787 B.n786 10.6151
R1591 B.n786 B.n785 10.6151
R1592 B.n785 B.n31 10.6151
R1593 B.n779 B.n31 10.6151
R1594 B.n779 B.n778 10.6151
R1595 B.n778 B.n777 10.6151
R1596 B.n777 B.n38 10.6151
R1597 B.n771 B.n38 10.6151
R1598 B.n771 B.n770 10.6151
R1599 B.n770 B.n769 10.6151
R1600 B.n769 B.n45 10.6151
R1601 B.n763 B.n45 10.6151
R1602 B.n763 B.n762 10.6151
R1603 B.n762 B.n761 10.6151
R1604 B.n761 B.n52 10.6151
R1605 B.n755 B.n52 10.6151
R1606 B.n755 B.n754 10.6151
R1607 B.n754 B.n753 10.6151
R1608 B.n753 B.n59 10.6151
R1609 B.n747 B.n59 10.6151
R1610 B.n747 B.n746 10.6151
R1611 B.n746 B.n745 10.6151
R1612 B.n745 B.n65 10.6151
R1613 B.n739 B.n65 10.6151
R1614 B.n739 B.n738 10.6151
R1615 B.n738 B.n737 10.6151
R1616 B.n737 B.n73 10.6151
R1617 B.n731 B.n73 10.6151
R1618 B.n731 B.n730 10.6151
R1619 B.n730 B.n729 10.6151
R1620 B.n729 B.n80 10.6151
R1621 B.n723 B.n80 10.6151
R1622 B.n723 B.n722 10.6151
R1623 B.n722 B.n721 10.6151
R1624 B.n721 B.n87 10.6151
R1625 B.n715 B.n87 10.6151
R1626 B.n715 B.n714 10.6151
R1627 B.n714 B.n713 10.6151
R1628 B.n713 B.n94 10.6151
R1629 B.n707 B.n94 10.6151
R1630 B.n707 B.n706 10.6151
R1631 B.n706 B.n705 10.6151
R1632 B.n705 B.n101 10.6151
R1633 B.n699 B.n101 10.6151
R1634 B.n699 B.n698 10.6151
R1635 B.n698 B.n697 10.6151
R1636 B.n697 B.n108 10.6151
R1637 B.n691 B.n108 10.6151
R1638 B.n691 B.n690 10.6151
R1639 B.n690 B.n689 10.6151
R1640 B.n158 B.n157 9.36635
R1641 B.n180 B.n179 9.36635
R1642 B.n365 B.n364 9.36635
R1643 B.n388 B.n332 9.36635
R1644 B.n817 B.n0 2.81026
R1645 B.n817 B.n1 2.81026
R1646 B.n248 B.t0 1.58666
R1647 B.t23 B.n766 1.58666
R1648 B.n159 B.n158 1.24928
R1649 B.n179 B.n178 1.24928
R1650 B.n366 B.n365 1.24928
R1651 B.n333 B.n332 1.24928
R1652 VP.n26 VP.n23 161.3
R1653 VP.n28 VP.n27 161.3
R1654 VP.n29 VP.n22 161.3
R1655 VP.n31 VP.n30 161.3
R1656 VP.n32 VP.n21 161.3
R1657 VP.n34 VP.n33 161.3
R1658 VP.n36 VP.n20 161.3
R1659 VP.n38 VP.n37 161.3
R1660 VP.n39 VP.n19 161.3
R1661 VP.n41 VP.n40 161.3
R1662 VP.n42 VP.n18 161.3
R1663 VP.n45 VP.n44 161.3
R1664 VP.n46 VP.n17 161.3
R1665 VP.n48 VP.n47 161.3
R1666 VP.n49 VP.n16 161.3
R1667 VP.n51 VP.n50 161.3
R1668 VP.n52 VP.n15 161.3
R1669 VP.n54 VP.n53 161.3
R1670 VP.n55 VP.n14 161.3
R1671 VP.n100 VP.n0 161.3
R1672 VP.n99 VP.n98 161.3
R1673 VP.n97 VP.n1 161.3
R1674 VP.n96 VP.n95 161.3
R1675 VP.n94 VP.n2 161.3
R1676 VP.n93 VP.n92 161.3
R1677 VP.n91 VP.n3 161.3
R1678 VP.n90 VP.n89 161.3
R1679 VP.n87 VP.n4 161.3
R1680 VP.n86 VP.n85 161.3
R1681 VP.n84 VP.n5 161.3
R1682 VP.n83 VP.n82 161.3
R1683 VP.n81 VP.n6 161.3
R1684 VP.n79 VP.n78 161.3
R1685 VP.n77 VP.n7 161.3
R1686 VP.n76 VP.n75 161.3
R1687 VP.n74 VP.n8 161.3
R1688 VP.n73 VP.n72 161.3
R1689 VP.n71 VP.n9 161.3
R1690 VP.n70 VP.n69 161.3
R1691 VP.n67 VP.n10 161.3
R1692 VP.n66 VP.n65 161.3
R1693 VP.n64 VP.n11 161.3
R1694 VP.n63 VP.n62 161.3
R1695 VP.n61 VP.n12 161.3
R1696 VP.n60 VP.n59 161.3
R1697 VP.n58 VP.n13 105.499
R1698 VP.n102 VP.n101 105.499
R1699 VP.n57 VP.n56 105.499
R1700 VP.n75 VP.n74 56.0773
R1701 VP.n86 VP.n5 56.0773
R1702 VP.n41 VP.n19 56.0773
R1703 VP.n30 VP.n29 56.0773
R1704 VP.n25 VP.n24 52.6217
R1705 VP.n25 VP.t2 48.2268
R1706 VP.n58 VP.n57 46.6512
R1707 VP.n62 VP.n11 42.5146
R1708 VP.n95 VP.n1 42.5146
R1709 VP.n50 VP.n15 42.5146
R1710 VP.n66 VP.n11 38.6395
R1711 VP.n95 VP.n94 38.6395
R1712 VP.n50 VP.n49 38.6395
R1713 VP.n74 VP.n73 25.0767
R1714 VP.n87 VP.n86 25.0767
R1715 VP.n42 VP.n41 25.0767
R1716 VP.n29 VP.n28 25.0767
R1717 VP.n61 VP.n60 24.5923
R1718 VP.n62 VP.n61 24.5923
R1719 VP.n67 VP.n66 24.5923
R1720 VP.n69 VP.n67 24.5923
R1721 VP.n73 VP.n9 24.5923
R1722 VP.n75 VP.n7 24.5923
R1723 VP.n79 VP.n7 24.5923
R1724 VP.n82 VP.n81 24.5923
R1725 VP.n82 VP.n5 24.5923
R1726 VP.n89 VP.n87 24.5923
R1727 VP.n93 VP.n3 24.5923
R1728 VP.n94 VP.n93 24.5923
R1729 VP.n99 VP.n1 24.5923
R1730 VP.n100 VP.n99 24.5923
R1731 VP.n54 VP.n15 24.5923
R1732 VP.n55 VP.n54 24.5923
R1733 VP.n44 VP.n42 24.5923
R1734 VP.n48 VP.n17 24.5923
R1735 VP.n49 VP.n48 24.5923
R1736 VP.n30 VP.n21 24.5923
R1737 VP.n34 VP.n21 24.5923
R1738 VP.n37 VP.n36 24.5923
R1739 VP.n37 VP.n19 24.5923
R1740 VP.n28 VP.n23 24.5923
R1741 VP.n68 VP.n9 21.1495
R1742 VP.n89 VP.n88 21.1495
R1743 VP.n44 VP.n43 21.1495
R1744 VP.n24 VP.n23 21.1495
R1745 VP.n13 VP.t5 14.0377
R1746 VP.n68 VP.t3 14.0377
R1747 VP.n80 VP.t9 14.0377
R1748 VP.n88 VP.t6 14.0377
R1749 VP.n101 VP.t4 14.0377
R1750 VP.n56 VP.t0 14.0377
R1751 VP.n43 VP.t7 14.0377
R1752 VP.n35 VP.t1 14.0377
R1753 VP.n24 VP.t8 14.0377
R1754 VP.n80 VP.n79 12.2964
R1755 VP.n81 VP.n80 12.2964
R1756 VP.n35 VP.n34 12.2964
R1757 VP.n36 VP.n35 12.2964
R1758 VP.n60 VP.n13 5.4107
R1759 VP.n101 VP.n100 5.4107
R1760 VP.n56 VP.n55 5.4107
R1761 VP.n26 VP.n25 4.94439
R1762 VP.n69 VP.n68 3.44336
R1763 VP.n88 VP.n3 3.44336
R1764 VP.n43 VP.n17 3.44336
R1765 VP.n57 VP.n14 0.278335
R1766 VP.n59 VP.n58 0.278335
R1767 VP.n102 VP.n0 0.278335
R1768 VP.n27 VP.n26 0.189894
R1769 VP.n27 VP.n22 0.189894
R1770 VP.n31 VP.n22 0.189894
R1771 VP.n32 VP.n31 0.189894
R1772 VP.n33 VP.n32 0.189894
R1773 VP.n33 VP.n20 0.189894
R1774 VP.n38 VP.n20 0.189894
R1775 VP.n39 VP.n38 0.189894
R1776 VP.n40 VP.n39 0.189894
R1777 VP.n40 VP.n18 0.189894
R1778 VP.n45 VP.n18 0.189894
R1779 VP.n46 VP.n45 0.189894
R1780 VP.n47 VP.n46 0.189894
R1781 VP.n47 VP.n16 0.189894
R1782 VP.n51 VP.n16 0.189894
R1783 VP.n52 VP.n51 0.189894
R1784 VP.n53 VP.n52 0.189894
R1785 VP.n53 VP.n14 0.189894
R1786 VP.n59 VP.n12 0.189894
R1787 VP.n63 VP.n12 0.189894
R1788 VP.n64 VP.n63 0.189894
R1789 VP.n65 VP.n64 0.189894
R1790 VP.n65 VP.n10 0.189894
R1791 VP.n70 VP.n10 0.189894
R1792 VP.n71 VP.n70 0.189894
R1793 VP.n72 VP.n71 0.189894
R1794 VP.n72 VP.n8 0.189894
R1795 VP.n76 VP.n8 0.189894
R1796 VP.n77 VP.n76 0.189894
R1797 VP.n78 VP.n77 0.189894
R1798 VP.n78 VP.n6 0.189894
R1799 VP.n83 VP.n6 0.189894
R1800 VP.n84 VP.n83 0.189894
R1801 VP.n85 VP.n84 0.189894
R1802 VP.n85 VP.n4 0.189894
R1803 VP.n90 VP.n4 0.189894
R1804 VP.n91 VP.n90 0.189894
R1805 VP.n92 VP.n91 0.189894
R1806 VP.n92 VP.n2 0.189894
R1807 VP.n96 VP.n2 0.189894
R1808 VP.n97 VP.n96 0.189894
R1809 VP.n98 VP.n97 0.189894
R1810 VP.n98 VP.n0 0.189894
R1811 VP VP.n102 0.153485
R1812 VDD1.n1 VDD1.t7 131.034
R1813 VDD1.n3 VDD1.t4 131.034
R1814 VDD1.n5 VDD1.n4 118.365
R1815 VDD1.n3 VDD1.n2 116.365
R1816 VDD1.n7 VDD1.n6 116.365
R1817 VDD1.n1 VDD1.n0 116.365
R1818 VDD1.n7 VDD1.n5 40.1216
R1819 VDD1.n6 VDD1.t2 11.9282
R1820 VDD1.n6 VDD1.t9 11.9282
R1821 VDD1.n0 VDD1.t1 11.9282
R1822 VDD1.n0 VDD1.t8 11.9282
R1823 VDD1.n4 VDD1.t3 11.9282
R1824 VDD1.n4 VDD1.t5 11.9282
R1825 VDD1.n2 VDD1.t6 11.9282
R1826 VDD1.n2 VDD1.t0 11.9282
R1827 VDD1 VDD1.n7 1.99834
R1828 VDD1 VDD1.n1 0.744035
R1829 VDD1.n5 VDD1.n3 0.630499
C0 VN VDD2 1.96238f
C1 VDD1 VTAIL 5.9012f
C2 VP VDD1 2.42051f
C3 VDD2 VTAIL 5.95626f
C4 VP VDD2 0.6235f
C5 VN VTAIL 3.56337f
C6 VP VN 6.851009f
C7 VDD2 VDD1 2.33525f
C8 VN VDD1 0.16112f
C9 VP VTAIL 3.5775f
C10 VDD2 B 5.651857f
C11 VDD1 B 5.6762f
C12 VTAIL B 3.690101f
C13 VN B 18.303299f
C14 VP B 16.858114f
C15 VDD1.t7 B 0.328222f
C16 VDD1.t1 B 0.040675f
C17 VDD1.t8 B 0.040675f
C18 VDD1.n0 B 0.23416f
C19 VDD1.n1 B 1.11499f
C20 VDD1.t4 B 0.328222f
C21 VDD1.t6 B 0.040675f
C22 VDD1.t0 B 0.040675f
C23 VDD1.n2 B 0.23416f
C24 VDD1.n3 B 1.10479f
C25 VDD1.t3 B 0.040675f
C26 VDD1.t5 B 0.040675f
C27 VDD1.n4 B 0.246303f
C28 VDD1.n5 B 3.13127f
C29 VDD1.t2 B 0.040675f
C30 VDD1.t9 B 0.040675f
C31 VDD1.n6 B 0.23416f
C32 VDD1.n7 B 3.04443f
C33 VP.n0 B 0.040903f
C34 VP.t4 B 0.328761f
C35 VP.n1 B 0.060649f
C36 VP.n2 B 0.031026f
C37 VP.n3 B 0.033108f
C38 VP.n4 B 0.031026f
C39 VP.n5 B 0.052751f
C40 VP.n6 B 0.031026f
C41 VP.t9 B 0.328761f
C42 VP.n7 B 0.057536f
C43 VP.n8 B 0.031026f
C44 VP.n9 B 0.053559f
C45 VP.n10 B 0.031026f
C46 VP.n11 B 0.025218f
C47 VP.n12 B 0.031026f
C48 VP.t5 B 0.328761f
C49 VP.n13 B 0.271322f
C50 VP.n14 B 0.040903f
C51 VP.t0 B 0.328761f
C52 VP.n15 B 0.060649f
C53 VP.n16 B 0.031026f
C54 VP.n17 B 0.033108f
C55 VP.n18 B 0.031026f
C56 VP.n19 B 0.052751f
C57 VP.n20 B 0.031026f
C58 VP.t1 B 0.328761f
C59 VP.n21 B 0.057536f
C60 VP.n22 B 0.031026f
C61 VP.n23 B 0.053559f
C62 VP.t2 B 0.594533f
C63 VP.t8 B 0.328761f
C64 VP.n24 B 0.271728f
C65 VP.n25 B 0.260015f
C66 VP.n26 B 0.327206f
C67 VP.n27 B 0.031026f
C68 VP.n28 B 0.058073f
C69 VP.n29 B 0.036915f
C70 VP.n30 B 0.052751f
C71 VP.n31 B 0.031026f
C72 VP.n32 B 0.031026f
C73 VP.n33 B 0.031026f
C74 VP.n34 B 0.043334f
C75 VP.n35 B 0.165525f
C76 VP.n36 B 0.043334f
C77 VP.n37 B 0.057536f
C78 VP.n38 B 0.031026f
C79 VP.n39 B 0.031026f
C80 VP.n40 B 0.031026f
C81 VP.n41 B 0.036915f
C82 VP.n42 B 0.058073f
C83 VP.t7 B 0.328761f
C84 VP.n43 B 0.165525f
C85 VP.n44 B 0.053559f
C86 VP.n45 B 0.031026f
C87 VP.n46 B 0.031026f
C88 VP.n47 B 0.031026f
C89 VP.n48 B 0.057536f
C90 VP.n49 B 0.061873f
C91 VP.n50 B 0.025218f
C92 VP.n51 B 0.031026f
C93 VP.n52 B 0.031026f
C94 VP.n53 B 0.031026f
C95 VP.n54 B 0.057536f
C96 VP.n55 B 0.035381f
C97 VP.n56 B 0.271322f
C98 VP.n57 B 1.56312f
C99 VP.n58 B 1.5871f
C100 VP.n59 B 0.040903f
C101 VP.n60 B 0.035381f
C102 VP.n61 B 0.057536f
C103 VP.n62 B 0.060649f
C104 VP.n63 B 0.031026f
C105 VP.n64 B 0.031026f
C106 VP.n65 B 0.031026f
C107 VP.n66 B 0.061873f
C108 VP.n67 B 0.057536f
C109 VP.t3 B 0.328761f
C110 VP.n68 B 0.165525f
C111 VP.n69 B 0.033108f
C112 VP.n70 B 0.031026f
C113 VP.n71 B 0.031026f
C114 VP.n72 B 0.031026f
C115 VP.n73 B 0.058073f
C116 VP.n74 B 0.036915f
C117 VP.n75 B 0.052751f
C118 VP.n76 B 0.031026f
C119 VP.n77 B 0.031026f
C120 VP.n78 B 0.031026f
C121 VP.n79 B 0.043334f
C122 VP.n80 B 0.165525f
C123 VP.n81 B 0.043334f
C124 VP.n82 B 0.057536f
C125 VP.n83 B 0.031026f
C126 VP.n84 B 0.031026f
C127 VP.n85 B 0.031026f
C128 VP.n86 B 0.036915f
C129 VP.n87 B 0.058073f
C130 VP.t6 B 0.328761f
C131 VP.n88 B 0.165525f
C132 VP.n89 B 0.053559f
C133 VP.n90 B 0.031026f
C134 VP.n91 B 0.031026f
C135 VP.n92 B 0.031026f
C136 VP.n93 B 0.057536f
C137 VP.n94 B 0.061873f
C138 VP.n95 B 0.025218f
C139 VP.n96 B 0.031026f
C140 VP.n97 B 0.031026f
C141 VP.n98 B 0.031026f
C142 VP.n99 B 0.057536f
C143 VP.n100 B 0.035381f
C144 VP.n101 B 0.271322f
C145 VP.n102 B 0.056674f
C146 VTAIL.t16 B 0.051118f
C147 VTAIL.t15 B 0.051118f
C148 VTAIL.n0 B 0.246785f
C149 VTAIL.n1 B 0.78238f
C150 VTAIL.t2 B 0.350389f
C151 VTAIL.n2 B 0.896938f
C152 VTAIL.t0 B 0.051118f
C153 VTAIL.t3 B 0.051118f
C154 VTAIL.n3 B 0.246785f
C155 VTAIL.n4 B 0.974246f
C156 VTAIL.t1 B 0.051118f
C157 VTAIL.t4 B 0.051118f
C158 VTAIL.n5 B 0.246785f
C159 VTAIL.n6 B 2.0275f
C160 VTAIL.t13 B 0.051118f
C161 VTAIL.t17 B 0.051118f
C162 VTAIL.n7 B 0.246786f
C163 VTAIL.n8 B 2.02749f
C164 VTAIL.t10 B 0.051118f
C165 VTAIL.t18 B 0.051118f
C166 VTAIL.n9 B 0.246786f
C167 VTAIL.n10 B 0.974245f
C168 VTAIL.t14 B 0.35039f
C169 VTAIL.n11 B 0.896937f
C170 VTAIL.t7 B 0.051118f
C171 VTAIL.t5 B 0.051118f
C172 VTAIL.n12 B 0.246786f
C173 VTAIL.n13 B 0.861128f
C174 VTAIL.t9 B 0.051118f
C175 VTAIL.t8 B 0.051118f
C176 VTAIL.n14 B 0.246786f
C177 VTAIL.n15 B 0.974245f
C178 VTAIL.t6 B 0.35039f
C179 VTAIL.n16 B 1.71908f
C180 VTAIL.t12 B 0.350389f
C181 VTAIL.n17 B 1.71908f
C182 VTAIL.t11 B 0.051118f
C183 VTAIL.t19 B 0.051118f
C184 VTAIL.n18 B 0.246785f
C185 VTAIL.n19 B 0.708773f
C186 VDD2.t2 B 0.259811f
C187 VDD2.t0 B 0.032197f
C188 VDD2.t4 B 0.032197f
C189 VDD2.n0 B 0.185354f
C190 VDD2.n1 B 0.874516f
C191 VDD2.t6 B 0.032197f
C192 VDD2.t3 B 0.032197f
C193 VDD2.n2 B 0.194966f
C194 VDD2.n3 B 2.35898f
C195 VDD2.t8 B 0.250762f
C196 VDD2.n4 B 2.30327f
C197 VDD2.t5 B 0.032197f
C198 VDD2.t7 B 0.032197f
C199 VDD2.n5 B 0.185355f
C200 VDD2.n6 B 0.459078f
C201 VDD2.t9 B 0.032197f
C202 VDD2.t1 B 0.032197f
C203 VDD2.n7 B 0.194945f
C204 VN.n0 B 0.033181f
C205 VN.t7 B 0.266694f
C206 VN.n1 B 0.049199f
C207 VN.n2 B 0.025169f
C208 VN.n3 B 0.026858f
C209 VN.n4 B 0.025169f
C210 VN.n5 B 0.042792f
C211 VN.n6 B 0.025169f
C212 VN.t8 B 0.266694f
C213 VN.n7 B 0.046674f
C214 VN.n8 B 0.025169f
C215 VN.n9 B 0.043448f
C216 VN.t3 B 0.482292f
C217 VN.t4 B 0.266694f
C218 VN.n10 B 0.220429f
C219 VN.n11 B 0.210927f
C220 VN.n12 B 0.265433f
C221 VN.n13 B 0.025169f
C222 VN.n14 B 0.04711f
C223 VN.n15 B 0.029945f
C224 VN.n16 B 0.042792f
C225 VN.n17 B 0.025169f
C226 VN.n18 B 0.025169f
C227 VN.n19 B 0.025169f
C228 VN.n20 B 0.035153f
C229 VN.n21 B 0.134276f
C230 VN.n22 B 0.035153f
C231 VN.n23 B 0.046674f
C232 VN.n24 B 0.025169f
C233 VN.n25 B 0.025169f
C234 VN.n26 B 0.025169f
C235 VN.n27 B 0.029945f
C236 VN.n28 B 0.04711f
C237 VN.t0 B 0.266694f
C238 VN.n29 B 0.134276f
C239 VN.n30 B 0.043448f
C240 VN.n31 B 0.025169f
C241 VN.n32 B 0.025169f
C242 VN.n33 B 0.025169f
C243 VN.n34 B 0.046674f
C244 VN.n35 B 0.050192f
C245 VN.n36 B 0.020457f
C246 VN.n37 B 0.025169f
C247 VN.n38 B 0.025169f
C248 VN.n39 B 0.025169f
C249 VN.n40 B 0.046674f
C250 VN.n41 B 0.028701f
C251 VN.n42 B 0.2201f
C252 VN.n43 B 0.045975f
C253 VN.n44 B 0.033181f
C254 VN.t6 B 0.266694f
C255 VN.n45 B 0.049199f
C256 VN.n46 B 0.025169f
C257 VN.n47 B 0.026858f
C258 VN.n48 B 0.025169f
C259 VN.t2 B 0.266694f
C260 VN.n49 B 0.134276f
C261 VN.n50 B 0.042792f
C262 VN.n51 B 0.025169f
C263 VN.t9 B 0.266694f
C264 VN.n52 B 0.046674f
C265 VN.n53 B 0.025169f
C266 VN.n54 B 0.043448f
C267 VN.t5 B 0.482292f
C268 VN.t1 B 0.266694f
C269 VN.n55 B 0.220429f
C270 VN.n56 B 0.210927f
C271 VN.n57 B 0.265433f
C272 VN.n58 B 0.025169f
C273 VN.n59 B 0.04711f
C274 VN.n60 B 0.029945f
C275 VN.n61 B 0.042792f
C276 VN.n62 B 0.025169f
C277 VN.n63 B 0.025169f
C278 VN.n64 B 0.025169f
C279 VN.n65 B 0.035153f
C280 VN.n66 B 0.134276f
C281 VN.n67 B 0.035153f
C282 VN.n68 B 0.046674f
C283 VN.n69 B 0.025169f
C284 VN.n70 B 0.025169f
C285 VN.n71 B 0.025169f
C286 VN.n72 B 0.029945f
C287 VN.n73 B 0.04711f
C288 VN.n74 B 0.043448f
C289 VN.n75 B 0.025169f
C290 VN.n76 B 0.025169f
C291 VN.n77 B 0.025169f
C292 VN.n78 B 0.046674f
C293 VN.n79 B 0.050192f
C294 VN.n80 B 0.020457f
C295 VN.n81 B 0.025169f
C296 VN.n82 B 0.025169f
C297 VN.n83 B 0.025169f
C298 VN.n84 B 0.046674f
C299 VN.n85 B 0.028701f
C300 VN.n86 B 0.2201f
C301 VN.n87 B 1.2817f
.ends

