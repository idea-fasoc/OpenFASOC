* NGSPICE file created from diff_pair_sample_0838.ext - technology: sky130A

.subckt diff_pair_sample_0838 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t7 VN.t0 VTAIL.t8 B.t4 sky130_fd_pr__nfet_01v8 ad=0.68475 pd=4.48 as=0.68475 ps=4.48 w=4.15 l=2.95
X1 VTAIL.t3 VP.t0 VDD1.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=0.68475 pd=4.48 as=0.68475 ps=4.48 w=4.15 l=2.95
X2 B.t21 B.t19 B.t20 B.t9 sky130_fd_pr__nfet_01v8 ad=1.6185 pd=9.08 as=0 ps=0 w=4.15 l=2.95
X3 B.t18 B.t16 B.t17 B.t13 sky130_fd_pr__nfet_01v8 ad=1.6185 pd=9.08 as=0 ps=0 w=4.15 l=2.95
X4 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=1.6185 pd=9.08 as=0 ps=0 w=4.15 l=2.95
X5 VDD1.t6 VP.t1 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=0.68475 pd=4.48 as=0.68475 ps=4.48 w=4.15 l=2.95
X6 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=1.6185 pd=9.08 as=0 ps=0 w=4.15 l=2.95
X7 VTAIL.t10 VN.t1 VDD2.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=0.68475 pd=4.48 as=0.68475 ps=4.48 w=4.15 l=2.95
X8 VTAIL.t11 VN.t2 VDD2.t5 B.t1 sky130_fd_pr__nfet_01v8 ad=1.6185 pd=9.08 as=0.68475 ps=4.48 w=4.15 l=2.95
X9 VDD1.t5 VP.t2 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=0.68475 pd=4.48 as=1.6185 ps=9.08 w=4.15 l=2.95
X10 VDD2.t4 VN.t3 VTAIL.t12 B.t5 sky130_fd_pr__nfet_01v8 ad=0.68475 pd=4.48 as=1.6185 ps=9.08 w=4.15 l=2.95
X11 VTAIL.t9 VN.t4 VDD2.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.68475 pd=4.48 as=0.68475 ps=4.48 w=4.15 l=2.95
X12 VTAIL.t0 VP.t3 VDD1.t4 B.t0 sky130_fd_pr__nfet_01v8 ad=1.6185 pd=9.08 as=0.68475 ps=4.48 w=4.15 l=2.95
X13 VDD1.t3 VP.t4 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.68475 pd=4.48 as=1.6185 ps=9.08 w=4.15 l=2.95
X14 VTAIL.t6 VP.t5 VDD1.t2 B.t6 sky130_fd_pr__nfet_01v8 ad=0.68475 pd=4.48 as=0.68475 ps=4.48 w=4.15 l=2.95
X15 VDD2.t2 VN.t5 VTAIL.t13 B.t2 sky130_fd_pr__nfet_01v8 ad=0.68475 pd=4.48 as=1.6185 ps=9.08 w=4.15 l=2.95
X16 VDD1.t1 VP.t6 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=0.68475 pd=4.48 as=0.68475 ps=4.48 w=4.15 l=2.95
X17 VTAIL.t14 VN.t6 VDD2.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=1.6185 pd=9.08 as=0.68475 ps=4.48 w=4.15 l=2.95
X18 VDD2.t0 VN.t7 VTAIL.t15 B.t7 sky130_fd_pr__nfet_01v8 ad=0.68475 pd=4.48 as=0.68475 ps=4.48 w=4.15 l=2.95
X19 VTAIL.t1 VP.t7 VDD1.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=1.6185 pd=9.08 as=0.68475 ps=4.48 w=4.15 l=2.95
R0 VN.n60 VN.n59 161.3
R1 VN.n58 VN.n32 161.3
R2 VN.n57 VN.n56 161.3
R3 VN.n55 VN.n33 161.3
R4 VN.n54 VN.n53 161.3
R5 VN.n52 VN.n34 161.3
R6 VN.n50 VN.n49 161.3
R7 VN.n48 VN.n35 161.3
R8 VN.n47 VN.n46 161.3
R9 VN.n45 VN.n36 161.3
R10 VN.n44 VN.n43 161.3
R11 VN.n42 VN.n37 161.3
R12 VN.n41 VN.n40 161.3
R13 VN.n29 VN.n28 161.3
R14 VN.n27 VN.n1 161.3
R15 VN.n26 VN.n25 161.3
R16 VN.n24 VN.n2 161.3
R17 VN.n23 VN.n22 161.3
R18 VN.n21 VN.n3 161.3
R19 VN.n19 VN.n18 161.3
R20 VN.n17 VN.n4 161.3
R21 VN.n16 VN.n15 161.3
R22 VN.n14 VN.n5 161.3
R23 VN.n13 VN.n12 161.3
R24 VN.n11 VN.n6 161.3
R25 VN.n10 VN.n9 161.3
R26 VN.n30 VN.n0 69.5151
R27 VN.n61 VN.n31 69.5151
R28 VN.n39 VN.n38 66.8451
R29 VN.n8 VN.n7 66.8451
R30 VN.n38 VN.t3 65.6241
R31 VN.n7 VN.t2 65.6241
R32 VN.n26 VN.n2 56.5193
R33 VN.n57 VN.n33 56.5193
R34 VN VN.n61 46.8692
R35 VN.n14 VN.n13 40.4934
R36 VN.n15 VN.n14 40.4934
R37 VN.n45 VN.n44 40.4934
R38 VN.n46 VN.n45 40.4934
R39 VN.n8 VN.t0 33.9039
R40 VN.n20 VN.t1 33.9039
R41 VN.n0 VN.t5 33.9039
R42 VN.n39 VN.t4 33.9039
R43 VN.n51 VN.t7 33.9039
R44 VN.n31 VN.t6 33.9039
R45 VN.n9 VN.n6 24.4675
R46 VN.n13 VN.n6 24.4675
R47 VN.n15 VN.n4 24.4675
R48 VN.n19 VN.n4 24.4675
R49 VN.n22 VN.n21 24.4675
R50 VN.n22 VN.n2 24.4675
R51 VN.n27 VN.n26 24.4675
R52 VN.n28 VN.n27 24.4675
R53 VN.n44 VN.n37 24.4675
R54 VN.n40 VN.n37 24.4675
R55 VN.n53 VN.n33 24.4675
R56 VN.n53 VN.n52 24.4675
R57 VN.n50 VN.n35 24.4675
R58 VN.n46 VN.n35 24.4675
R59 VN.n59 VN.n58 24.4675
R60 VN.n58 VN.n57 24.4675
R61 VN.n28 VN.n0 20.5528
R62 VN.n59 VN.n31 20.5528
R63 VN.n21 VN.n20 17.6167
R64 VN.n52 VN.n51 17.6167
R65 VN.n9 VN.n8 6.85126
R66 VN.n20 VN.n19 6.85126
R67 VN.n40 VN.n39 6.85126
R68 VN.n51 VN.n50 6.85126
R69 VN.n41 VN.n38 5.51404
R70 VN.n10 VN.n7 5.51404
R71 VN.n61 VN.n60 0.354971
R72 VN.n30 VN.n29 0.354971
R73 VN VN.n30 0.26696
R74 VN.n60 VN.n32 0.189894
R75 VN.n56 VN.n32 0.189894
R76 VN.n56 VN.n55 0.189894
R77 VN.n55 VN.n54 0.189894
R78 VN.n54 VN.n34 0.189894
R79 VN.n49 VN.n34 0.189894
R80 VN.n49 VN.n48 0.189894
R81 VN.n48 VN.n47 0.189894
R82 VN.n47 VN.n36 0.189894
R83 VN.n43 VN.n36 0.189894
R84 VN.n43 VN.n42 0.189894
R85 VN.n42 VN.n41 0.189894
R86 VN.n11 VN.n10 0.189894
R87 VN.n12 VN.n11 0.189894
R88 VN.n12 VN.n5 0.189894
R89 VN.n16 VN.n5 0.189894
R90 VN.n17 VN.n16 0.189894
R91 VN.n18 VN.n17 0.189894
R92 VN.n18 VN.n3 0.189894
R93 VN.n23 VN.n3 0.189894
R94 VN.n24 VN.n23 0.189894
R95 VN.n25 VN.n24 0.189894
R96 VN.n25 VN.n1 0.189894
R97 VN.n29 VN.n1 0.189894
R98 VTAIL.n11 VTAIL.t1 59.041
R99 VTAIL.n10 VTAIL.t12 59.041
R100 VTAIL.n7 VTAIL.t14 59.041
R101 VTAIL.n15 VTAIL.t13 59.0408
R102 VTAIL.n2 VTAIL.t11 59.0408
R103 VTAIL.n3 VTAIL.t5 59.0408
R104 VTAIL.n6 VTAIL.t0 59.0408
R105 VTAIL.n14 VTAIL.t2 59.0408
R106 VTAIL.n13 VTAIL.n12 54.27
R107 VTAIL.n9 VTAIL.n8 54.27
R108 VTAIL.n1 VTAIL.n0 54.2697
R109 VTAIL.n5 VTAIL.n4 54.2697
R110 VTAIL.n15 VTAIL.n14 18.7721
R111 VTAIL.n7 VTAIL.n6 18.7721
R112 VTAIL.n0 VTAIL.t8 4.77158
R113 VTAIL.n0 VTAIL.t10 4.77158
R114 VTAIL.n4 VTAIL.t7 4.77158
R115 VTAIL.n4 VTAIL.t3 4.77158
R116 VTAIL.n12 VTAIL.t4 4.77158
R117 VTAIL.n12 VTAIL.t6 4.77158
R118 VTAIL.n8 VTAIL.t15 4.77158
R119 VTAIL.n8 VTAIL.t9 4.77158
R120 VTAIL.n9 VTAIL.n7 2.82809
R121 VTAIL.n10 VTAIL.n9 2.82809
R122 VTAIL.n13 VTAIL.n11 2.82809
R123 VTAIL.n14 VTAIL.n13 2.82809
R124 VTAIL.n6 VTAIL.n5 2.82809
R125 VTAIL.n5 VTAIL.n3 2.82809
R126 VTAIL.n2 VTAIL.n1 2.82809
R127 VTAIL VTAIL.n15 2.7699
R128 VTAIL.n11 VTAIL.n10 0.470328
R129 VTAIL.n3 VTAIL.n2 0.470328
R130 VTAIL VTAIL.n1 0.0586897
R131 VDD2.n2 VDD2.n1 72.307
R132 VDD2.n2 VDD2.n0 72.307
R133 VDD2 VDD2.n5 72.3042
R134 VDD2.n4 VDD2.n3 70.9487
R135 VDD2.n4 VDD2.n2 40.017
R136 VDD2.n5 VDD2.t3 4.77158
R137 VDD2.n5 VDD2.t4 4.77158
R138 VDD2.n3 VDD2.t1 4.77158
R139 VDD2.n3 VDD2.t0 4.77158
R140 VDD2.n1 VDD2.t6 4.77158
R141 VDD2.n1 VDD2.t2 4.77158
R142 VDD2.n0 VDD2.t5 4.77158
R143 VDD2.n0 VDD2.t7 4.77158
R144 VDD2 VDD2.n4 1.47248
R145 B.n699 B.n698 585
R146 B.n700 B.n699 585
R147 B.n223 B.n128 585
R148 B.n222 B.n221 585
R149 B.n220 B.n219 585
R150 B.n218 B.n217 585
R151 B.n216 B.n215 585
R152 B.n214 B.n213 585
R153 B.n212 B.n211 585
R154 B.n210 B.n209 585
R155 B.n208 B.n207 585
R156 B.n206 B.n205 585
R157 B.n204 B.n203 585
R158 B.n202 B.n201 585
R159 B.n200 B.n199 585
R160 B.n198 B.n197 585
R161 B.n196 B.n195 585
R162 B.n194 B.n193 585
R163 B.n192 B.n191 585
R164 B.n190 B.n189 585
R165 B.n188 B.n187 585
R166 B.n186 B.n185 585
R167 B.n184 B.n183 585
R168 B.n182 B.n181 585
R169 B.n180 B.n179 585
R170 B.n178 B.n177 585
R171 B.n176 B.n175 585
R172 B.n174 B.n173 585
R173 B.n172 B.n171 585
R174 B.n169 B.n168 585
R175 B.n167 B.n166 585
R176 B.n165 B.n164 585
R177 B.n163 B.n162 585
R178 B.n161 B.n160 585
R179 B.n159 B.n158 585
R180 B.n157 B.n156 585
R181 B.n155 B.n154 585
R182 B.n153 B.n152 585
R183 B.n151 B.n150 585
R184 B.n149 B.n148 585
R185 B.n147 B.n146 585
R186 B.n145 B.n144 585
R187 B.n143 B.n142 585
R188 B.n141 B.n140 585
R189 B.n139 B.n138 585
R190 B.n137 B.n136 585
R191 B.n135 B.n134 585
R192 B.n103 B.n102 585
R193 B.n697 B.n104 585
R194 B.n701 B.n104 585
R195 B.n696 B.n695 585
R196 B.n695 B.n100 585
R197 B.n694 B.n99 585
R198 B.n707 B.n99 585
R199 B.n693 B.n98 585
R200 B.n708 B.n98 585
R201 B.n692 B.n97 585
R202 B.n709 B.n97 585
R203 B.n691 B.n690 585
R204 B.n690 B.n93 585
R205 B.n689 B.n92 585
R206 B.n715 B.n92 585
R207 B.n688 B.n91 585
R208 B.n716 B.n91 585
R209 B.n687 B.n90 585
R210 B.n717 B.n90 585
R211 B.n686 B.n685 585
R212 B.n685 B.n86 585
R213 B.n684 B.n85 585
R214 B.n723 B.n85 585
R215 B.n683 B.n84 585
R216 B.n724 B.n84 585
R217 B.n682 B.n83 585
R218 B.n725 B.n83 585
R219 B.n681 B.n680 585
R220 B.n680 B.n79 585
R221 B.n679 B.n78 585
R222 B.n731 B.n78 585
R223 B.n678 B.n77 585
R224 B.n732 B.n77 585
R225 B.n677 B.n76 585
R226 B.n733 B.n76 585
R227 B.n676 B.n675 585
R228 B.n675 B.n72 585
R229 B.n674 B.n71 585
R230 B.n739 B.n71 585
R231 B.n673 B.n70 585
R232 B.n740 B.n70 585
R233 B.n672 B.n69 585
R234 B.n741 B.n69 585
R235 B.n671 B.n670 585
R236 B.n670 B.n68 585
R237 B.n669 B.n64 585
R238 B.n747 B.n64 585
R239 B.n668 B.n63 585
R240 B.n748 B.n63 585
R241 B.n667 B.n62 585
R242 B.n749 B.n62 585
R243 B.n666 B.n665 585
R244 B.n665 B.n58 585
R245 B.n664 B.n57 585
R246 B.n755 B.n57 585
R247 B.n663 B.n56 585
R248 B.n756 B.n56 585
R249 B.n662 B.n55 585
R250 B.n757 B.n55 585
R251 B.n661 B.n660 585
R252 B.n660 B.n51 585
R253 B.n659 B.n50 585
R254 B.n763 B.n50 585
R255 B.n658 B.n49 585
R256 B.n764 B.n49 585
R257 B.n657 B.n48 585
R258 B.n765 B.n48 585
R259 B.n656 B.n655 585
R260 B.n655 B.n44 585
R261 B.n654 B.n43 585
R262 B.n771 B.n43 585
R263 B.n653 B.n42 585
R264 B.n772 B.n42 585
R265 B.n652 B.n41 585
R266 B.n773 B.n41 585
R267 B.n651 B.n650 585
R268 B.n650 B.n37 585
R269 B.n649 B.n36 585
R270 B.n779 B.n36 585
R271 B.n648 B.n35 585
R272 B.n780 B.n35 585
R273 B.n647 B.n34 585
R274 B.n781 B.n34 585
R275 B.n646 B.n645 585
R276 B.n645 B.n30 585
R277 B.n644 B.n29 585
R278 B.n787 B.n29 585
R279 B.n643 B.n28 585
R280 B.n788 B.n28 585
R281 B.n642 B.n27 585
R282 B.n789 B.n27 585
R283 B.n641 B.n640 585
R284 B.n640 B.n23 585
R285 B.n639 B.n22 585
R286 B.n795 B.n22 585
R287 B.n638 B.n21 585
R288 B.n796 B.n21 585
R289 B.n637 B.n20 585
R290 B.n797 B.n20 585
R291 B.n636 B.n635 585
R292 B.n635 B.n16 585
R293 B.n634 B.n15 585
R294 B.n803 B.n15 585
R295 B.n633 B.n14 585
R296 B.n804 B.n14 585
R297 B.n632 B.n13 585
R298 B.n805 B.n13 585
R299 B.n631 B.n630 585
R300 B.n630 B.n12 585
R301 B.n629 B.n628 585
R302 B.n629 B.n8 585
R303 B.n627 B.n7 585
R304 B.n812 B.n7 585
R305 B.n626 B.n6 585
R306 B.n813 B.n6 585
R307 B.n625 B.n5 585
R308 B.n814 B.n5 585
R309 B.n624 B.n623 585
R310 B.n623 B.n4 585
R311 B.n622 B.n224 585
R312 B.n622 B.n621 585
R313 B.n612 B.n225 585
R314 B.n226 B.n225 585
R315 B.n614 B.n613 585
R316 B.n615 B.n614 585
R317 B.n611 B.n231 585
R318 B.n231 B.n230 585
R319 B.n610 B.n609 585
R320 B.n609 B.n608 585
R321 B.n233 B.n232 585
R322 B.n234 B.n233 585
R323 B.n601 B.n600 585
R324 B.n602 B.n601 585
R325 B.n599 B.n239 585
R326 B.n239 B.n238 585
R327 B.n598 B.n597 585
R328 B.n597 B.n596 585
R329 B.n241 B.n240 585
R330 B.n242 B.n241 585
R331 B.n589 B.n588 585
R332 B.n590 B.n589 585
R333 B.n587 B.n247 585
R334 B.n247 B.n246 585
R335 B.n586 B.n585 585
R336 B.n585 B.n584 585
R337 B.n249 B.n248 585
R338 B.n250 B.n249 585
R339 B.n577 B.n576 585
R340 B.n578 B.n577 585
R341 B.n575 B.n255 585
R342 B.n255 B.n254 585
R343 B.n574 B.n573 585
R344 B.n573 B.n572 585
R345 B.n257 B.n256 585
R346 B.n258 B.n257 585
R347 B.n565 B.n564 585
R348 B.n566 B.n565 585
R349 B.n563 B.n263 585
R350 B.n263 B.n262 585
R351 B.n562 B.n561 585
R352 B.n561 B.n560 585
R353 B.n265 B.n264 585
R354 B.n266 B.n265 585
R355 B.n553 B.n552 585
R356 B.n554 B.n553 585
R357 B.n551 B.n271 585
R358 B.n271 B.n270 585
R359 B.n550 B.n549 585
R360 B.n549 B.n548 585
R361 B.n273 B.n272 585
R362 B.n274 B.n273 585
R363 B.n541 B.n540 585
R364 B.n542 B.n541 585
R365 B.n539 B.n279 585
R366 B.n279 B.n278 585
R367 B.n538 B.n537 585
R368 B.n537 B.n536 585
R369 B.n281 B.n280 585
R370 B.n282 B.n281 585
R371 B.n529 B.n528 585
R372 B.n530 B.n529 585
R373 B.n527 B.n287 585
R374 B.n287 B.n286 585
R375 B.n526 B.n525 585
R376 B.n525 B.n524 585
R377 B.n289 B.n288 585
R378 B.n517 B.n289 585
R379 B.n516 B.n515 585
R380 B.n518 B.n516 585
R381 B.n514 B.n294 585
R382 B.n294 B.n293 585
R383 B.n513 B.n512 585
R384 B.n512 B.n511 585
R385 B.n296 B.n295 585
R386 B.n297 B.n296 585
R387 B.n504 B.n503 585
R388 B.n505 B.n504 585
R389 B.n502 B.n302 585
R390 B.n302 B.n301 585
R391 B.n501 B.n500 585
R392 B.n500 B.n499 585
R393 B.n304 B.n303 585
R394 B.n305 B.n304 585
R395 B.n492 B.n491 585
R396 B.n493 B.n492 585
R397 B.n490 B.n310 585
R398 B.n310 B.n309 585
R399 B.n489 B.n488 585
R400 B.n488 B.n487 585
R401 B.n312 B.n311 585
R402 B.n313 B.n312 585
R403 B.n480 B.n479 585
R404 B.n481 B.n480 585
R405 B.n478 B.n318 585
R406 B.n318 B.n317 585
R407 B.n477 B.n476 585
R408 B.n476 B.n475 585
R409 B.n320 B.n319 585
R410 B.n321 B.n320 585
R411 B.n468 B.n467 585
R412 B.n469 B.n468 585
R413 B.n466 B.n326 585
R414 B.n326 B.n325 585
R415 B.n465 B.n464 585
R416 B.n464 B.n463 585
R417 B.n328 B.n327 585
R418 B.n329 B.n328 585
R419 B.n456 B.n455 585
R420 B.n457 B.n456 585
R421 B.n332 B.n331 585
R422 B.n361 B.n360 585
R423 B.n362 B.n358 585
R424 B.n358 B.n333 585
R425 B.n364 B.n363 585
R426 B.n366 B.n357 585
R427 B.n369 B.n368 585
R428 B.n370 B.n356 585
R429 B.n372 B.n371 585
R430 B.n374 B.n355 585
R431 B.n377 B.n376 585
R432 B.n378 B.n354 585
R433 B.n380 B.n379 585
R434 B.n382 B.n353 585
R435 B.n385 B.n384 585
R436 B.n386 B.n352 585
R437 B.n388 B.n387 585
R438 B.n390 B.n351 585
R439 B.n393 B.n392 585
R440 B.n394 B.n348 585
R441 B.n397 B.n396 585
R442 B.n399 B.n347 585
R443 B.n402 B.n401 585
R444 B.n403 B.n346 585
R445 B.n405 B.n404 585
R446 B.n407 B.n345 585
R447 B.n410 B.n409 585
R448 B.n411 B.n344 585
R449 B.n416 B.n415 585
R450 B.n418 B.n343 585
R451 B.n421 B.n420 585
R452 B.n422 B.n342 585
R453 B.n424 B.n423 585
R454 B.n426 B.n341 585
R455 B.n429 B.n428 585
R456 B.n430 B.n340 585
R457 B.n432 B.n431 585
R458 B.n434 B.n339 585
R459 B.n437 B.n436 585
R460 B.n438 B.n338 585
R461 B.n440 B.n439 585
R462 B.n442 B.n337 585
R463 B.n445 B.n444 585
R464 B.n446 B.n336 585
R465 B.n448 B.n447 585
R466 B.n450 B.n335 585
R467 B.n453 B.n452 585
R468 B.n454 B.n334 585
R469 B.n459 B.n458 585
R470 B.n458 B.n457 585
R471 B.n460 B.n330 585
R472 B.n330 B.n329 585
R473 B.n462 B.n461 585
R474 B.n463 B.n462 585
R475 B.n324 B.n323 585
R476 B.n325 B.n324 585
R477 B.n471 B.n470 585
R478 B.n470 B.n469 585
R479 B.n472 B.n322 585
R480 B.n322 B.n321 585
R481 B.n474 B.n473 585
R482 B.n475 B.n474 585
R483 B.n316 B.n315 585
R484 B.n317 B.n316 585
R485 B.n483 B.n482 585
R486 B.n482 B.n481 585
R487 B.n484 B.n314 585
R488 B.n314 B.n313 585
R489 B.n486 B.n485 585
R490 B.n487 B.n486 585
R491 B.n308 B.n307 585
R492 B.n309 B.n308 585
R493 B.n495 B.n494 585
R494 B.n494 B.n493 585
R495 B.n496 B.n306 585
R496 B.n306 B.n305 585
R497 B.n498 B.n497 585
R498 B.n499 B.n498 585
R499 B.n300 B.n299 585
R500 B.n301 B.n300 585
R501 B.n507 B.n506 585
R502 B.n506 B.n505 585
R503 B.n508 B.n298 585
R504 B.n298 B.n297 585
R505 B.n510 B.n509 585
R506 B.n511 B.n510 585
R507 B.n292 B.n291 585
R508 B.n293 B.n292 585
R509 B.n520 B.n519 585
R510 B.n519 B.n518 585
R511 B.n521 B.n290 585
R512 B.n517 B.n290 585
R513 B.n523 B.n522 585
R514 B.n524 B.n523 585
R515 B.n285 B.n284 585
R516 B.n286 B.n285 585
R517 B.n532 B.n531 585
R518 B.n531 B.n530 585
R519 B.n533 B.n283 585
R520 B.n283 B.n282 585
R521 B.n535 B.n534 585
R522 B.n536 B.n535 585
R523 B.n277 B.n276 585
R524 B.n278 B.n277 585
R525 B.n544 B.n543 585
R526 B.n543 B.n542 585
R527 B.n545 B.n275 585
R528 B.n275 B.n274 585
R529 B.n547 B.n546 585
R530 B.n548 B.n547 585
R531 B.n269 B.n268 585
R532 B.n270 B.n269 585
R533 B.n556 B.n555 585
R534 B.n555 B.n554 585
R535 B.n557 B.n267 585
R536 B.n267 B.n266 585
R537 B.n559 B.n558 585
R538 B.n560 B.n559 585
R539 B.n261 B.n260 585
R540 B.n262 B.n261 585
R541 B.n568 B.n567 585
R542 B.n567 B.n566 585
R543 B.n569 B.n259 585
R544 B.n259 B.n258 585
R545 B.n571 B.n570 585
R546 B.n572 B.n571 585
R547 B.n253 B.n252 585
R548 B.n254 B.n253 585
R549 B.n580 B.n579 585
R550 B.n579 B.n578 585
R551 B.n581 B.n251 585
R552 B.n251 B.n250 585
R553 B.n583 B.n582 585
R554 B.n584 B.n583 585
R555 B.n245 B.n244 585
R556 B.n246 B.n245 585
R557 B.n592 B.n591 585
R558 B.n591 B.n590 585
R559 B.n593 B.n243 585
R560 B.n243 B.n242 585
R561 B.n595 B.n594 585
R562 B.n596 B.n595 585
R563 B.n237 B.n236 585
R564 B.n238 B.n237 585
R565 B.n604 B.n603 585
R566 B.n603 B.n602 585
R567 B.n605 B.n235 585
R568 B.n235 B.n234 585
R569 B.n607 B.n606 585
R570 B.n608 B.n607 585
R571 B.n229 B.n228 585
R572 B.n230 B.n229 585
R573 B.n617 B.n616 585
R574 B.n616 B.n615 585
R575 B.n618 B.n227 585
R576 B.n227 B.n226 585
R577 B.n620 B.n619 585
R578 B.n621 B.n620 585
R579 B.n3 B.n0 585
R580 B.n4 B.n3 585
R581 B.n811 B.n1 585
R582 B.n812 B.n811 585
R583 B.n810 B.n809 585
R584 B.n810 B.n8 585
R585 B.n808 B.n9 585
R586 B.n12 B.n9 585
R587 B.n807 B.n806 585
R588 B.n806 B.n805 585
R589 B.n11 B.n10 585
R590 B.n804 B.n11 585
R591 B.n802 B.n801 585
R592 B.n803 B.n802 585
R593 B.n800 B.n17 585
R594 B.n17 B.n16 585
R595 B.n799 B.n798 585
R596 B.n798 B.n797 585
R597 B.n19 B.n18 585
R598 B.n796 B.n19 585
R599 B.n794 B.n793 585
R600 B.n795 B.n794 585
R601 B.n792 B.n24 585
R602 B.n24 B.n23 585
R603 B.n791 B.n790 585
R604 B.n790 B.n789 585
R605 B.n26 B.n25 585
R606 B.n788 B.n26 585
R607 B.n786 B.n785 585
R608 B.n787 B.n786 585
R609 B.n784 B.n31 585
R610 B.n31 B.n30 585
R611 B.n783 B.n782 585
R612 B.n782 B.n781 585
R613 B.n33 B.n32 585
R614 B.n780 B.n33 585
R615 B.n778 B.n777 585
R616 B.n779 B.n778 585
R617 B.n776 B.n38 585
R618 B.n38 B.n37 585
R619 B.n775 B.n774 585
R620 B.n774 B.n773 585
R621 B.n40 B.n39 585
R622 B.n772 B.n40 585
R623 B.n770 B.n769 585
R624 B.n771 B.n770 585
R625 B.n768 B.n45 585
R626 B.n45 B.n44 585
R627 B.n767 B.n766 585
R628 B.n766 B.n765 585
R629 B.n47 B.n46 585
R630 B.n764 B.n47 585
R631 B.n762 B.n761 585
R632 B.n763 B.n762 585
R633 B.n760 B.n52 585
R634 B.n52 B.n51 585
R635 B.n759 B.n758 585
R636 B.n758 B.n757 585
R637 B.n54 B.n53 585
R638 B.n756 B.n54 585
R639 B.n754 B.n753 585
R640 B.n755 B.n754 585
R641 B.n752 B.n59 585
R642 B.n59 B.n58 585
R643 B.n751 B.n750 585
R644 B.n750 B.n749 585
R645 B.n61 B.n60 585
R646 B.n748 B.n61 585
R647 B.n746 B.n745 585
R648 B.n747 B.n746 585
R649 B.n744 B.n65 585
R650 B.n68 B.n65 585
R651 B.n743 B.n742 585
R652 B.n742 B.n741 585
R653 B.n67 B.n66 585
R654 B.n740 B.n67 585
R655 B.n738 B.n737 585
R656 B.n739 B.n738 585
R657 B.n736 B.n73 585
R658 B.n73 B.n72 585
R659 B.n735 B.n734 585
R660 B.n734 B.n733 585
R661 B.n75 B.n74 585
R662 B.n732 B.n75 585
R663 B.n730 B.n729 585
R664 B.n731 B.n730 585
R665 B.n728 B.n80 585
R666 B.n80 B.n79 585
R667 B.n727 B.n726 585
R668 B.n726 B.n725 585
R669 B.n82 B.n81 585
R670 B.n724 B.n82 585
R671 B.n722 B.n721 585
R672 B.n723 B.n722 585
R673 B.n720 B.n87 585
R674 B.n87 B.n86 585
R675 B.n719 B.n718 585
R676 B.n718 B.n717 585
R677 B.n89 B.n88 585
R678 B.n716 B.n89 585
R679 B.n714 B.n713 585
R680 B.n715 B.n714 585
R681 B.n712 B.n94 585
R682 B.n94 B.n93 585
R683 B.n711 B.n710 585
R684 B.n710 B.n709 585
R685 B.n96 B.n95 585
R686 B.n708 B.n96 585
R687 B.n706 B.n705 585
R688 B.n707 B.n706 585
R689 B.n704 B.n101 585
R690 B.n101 B.n100 585
R691 B.n703 B.n702 585
R692 B.n702 B.n701 585
R693 B.n815 B.n814 585
R694 B.n813 B.n2 585
R695 B.n702 B.n103 444.452
R696 B.n699 B.n104 444.452
R697 B.n456 B.n334 444.452
R698 B.n458 B.n332 444.452
R699 B.n700 B.n127 256.663
R700 B.n700 B.n126 256.663
R701 B.n700 B.n125 256.663
R702 B.n700 B.n124 256.663
R703 B.n700 B.n123 256.663
R704 B.n700 B.n122 256.663
R705 B.n700 B.n121 256.663
R706 B.n700 B.n120 256.663
R707 B.n700 B.n119 256.663
R708 B.n700 B.n118 256.663
R709 B.n700 B.n117 256.663
R710 B.n700 B.n116 256.663
R711 B.n700 B.n115 256.663
R712 B.n700 B.n114 256.663
R713 B.n700 B.n113 256.663
R714 B.n700 B.n112 256.663
R715 B.n700 B.n111 256.663
R716 B.n700 B.n110 256.663
R717 B.n700 B.n109 256.663
R718 B.n700 B.n108 256.663
R719 B.n700 B.n107 256.663
R720 B.n700 B.n106 256.663
R721 B.n700 B.n105 256.663
R722 B.n359 B.n333 256.663
R723 B.n365 B.n333 256.663
R724 B.n367 B.n333 256.663
R725 B.n373 B.n333 256.663
R726 B.n375 B.n333 256.663
R727 B.n381 B.n333 256.663
R728 B.n383 B.n333 256.663
R729 B.n389 B.n333 256.663
R730 B.n391 B.n333 256.663
R731 B.n398 B.n333 256.663
R732 B.n400 B.n333 256.663
R733 B.n406 B.n333 256.663
R734 B.n408 B.n333 256.663
R735 B.n417 B.n333 256.663
R736 B.n419 B.n333 256.663
R737 B.n425 B.n333 256.663
R738 B.n427 B.n333 256.663
R739 B.n433 B.n333 256.663
R740 B.n435 B.n333 256.663
R741 B.n441 B.n333 256.663
R742 B.n443 B.n333 256.663
R743 B.n449 B.n333 256.663
R744 B.n451 B.n333 256.663
R745 B.n817 B.n816 256.663
R746 B.n132 B.t12 242.423
R747 B.n129 B.t16 242.423
R748 B.n412 B.t19 242.423
R749 B.n349 B.t8 242.423
R750 B.n136 B.n135 163.367
R751 B.n140 B.n139 163.367
R752 B.n144 B.n143 163.367
R753 B.n148 B.n147 163.367
R754 B.n152 B.n151 163.367
R755 B.n156 B.n155 163.367
R756 B.n160 B.n159 163.367
R757 B.n164 B.n163 163.367
R758 B.n168 B.n167 163.367
R759 B.n173 B.n172 163.367
R760 B.n177 B.n176 163.367
R761 B.n181 B.n180 163.367
R762 B.n185 B.n184 163.367
R763 B.n189 B.n188 163.367
R764 B.n193 B.n192 163.367
R765 B.n197 B.n196 163.367
R766 B.n201 B.n200 163.367
R767 B.n205 B.n204 163.367
R768 B.n209 B.n208 163.367
R769 B.n213 B.n212 163.367
R770 B.n217 B.n216 163.367
R771 B.n221 B.n220 163.367
R772 B.n699 B.n128 163.367
R773 B.n456 B.n328 163.367
R774 B.n464 B.n328 163.367
R775 B.n464 B.n326 163.367
R776 B.n468 B.n326 163.367
R777 B.n468 B.n320 163.367
R778 B.n476 B.n320 163.367
R779 B.n476 B.n318 163.367
R780 B.n480 B.n318 163.367
R781 B.n480 B.n312 163.367
R782 B.n488 B.n312 163.367
R783 B.n488 B.n310 163.367
R784 B.n492 B.n310 163.367
R785 B.n492 B.n304 163.367
R786 B.n500 B.n304 163.367
R787 B.n500 B.n302 163.367
R788 B.n504 B.n302 163.367
R789 B.n504 B.n296 163.367
R790 B.n512 B.n296 163.367
R791 B.n512 B.n294 163.367
R792 B.n516 B.n294 163.367
R793 B.n516 B.n289 163.367
R794 B.n525 B.n289 163.367
R795 B.n525 B.n287 163.367
R796 B.n529 B.n287 163.367
R797 B.n529 B.n281 163.367
R798 B.n537 B.n281 163.367
R799 B.n537 B.n279 163.367
R800 B.n541 B.n279 163.367
R801 B.n541 B.n273 163.367
R802 B.n549 B.n273 163.367
R803 B.n549 B.n271 163.367
R804 B.n553 B.n271 163.367
R805 B.n553 B.n265 163.367
R806 B.n561 B.n265 163.367
R807 B.n561 B.n263 163.367
R808 B.n565 B.n263 163.367
R809 B.n565 B.n257 163.367
R810 B.n573 B.n257 163.367
R811 B.n573 B.n255 163.367
R812 B.n577 B.n255 163.367
R813 B.n577 B.n249 163.367
R814 B.n585 B.n249 163.367
R815 B.n585 B.n247 163.367
R816 B.n589 B.n247 163.367
R817 B.n589 B.n241 163.367
R818 B.n597 B.n241 163.367
R819 B.n597 B.n239 163.367
R820 B.n601 B.n239 163.367
R821 B.n601 B.n233 163.367
R822 B.n609 B.n233 163.367
R823 B.n609 B.n231 163.367
R824 B.n614 B.n231 163.367
R825 B.n614 B.n225 163.367
R826 B.n622 B.n225 163.367
R827 B.n623 B.n622 163.367
R828 B.n623 B.n5 163.367
R829 B.n6 B.n5 163.367
R830 B.n7 B.n6 163.367
R831 B.n629 B.n7 163.367
R832 B.n630 B.n629 163.367
R833 B.n630 B.n13 163.367
R834 B.n14 B.n13 163.367
R835 B.n15 B.n14 163.367
R836 B.n635 B.n15 163.367
R837 B.n635 B.n20 163.367
R838 B.n21 B.n20 163.367
R839 B.n22 B.n21 163.367
R840 B.n640 B.n22 163.367
R841 B.n640 B.n27 163.367
R842 B.n28 B.n27 163.367
R843 B.n29 B.n28 163.367
R844 B.n645 B.n29 163.367
R845 B.n645 B.n34 163.367
R846 B.n35 B.n34 163.367
R847 B.n36 B.n35 163.367
R848 B.n650 B.n36 163.367
R849 B.n650 B.n41 163.367
R850 B.n42 B.n41 163.367
R851 B.n43 B.n42 163.367
R852 B.n655 B.n43 163.367
R853 B.n655 B.n48 163.367
R854 B.n49 B.n48 163.367
R855 B.n50 B.n49 163.367
R856 B.n660 B.n50 163.367
R857 B.n660 B.n55 163.367
R858 B.n56 B.n55 163.367
R859 B.n57 B.n56 163.367
R860 B.n665 B.n57 163.367
R861 B.n665 B.n62 163.367
R862 B.n63 B.n62 163.367
R863 B.n64 B.n63 163.367
R864 B.n670 B.n64 163.367
R865 B.n670 B.n69 163.367
R866 B.n70 B.n69 163.367
R867 B.n71 B.n70 163.367
R868 B.n675 B.n71 163.367
R869 B.n675 B.n76 163.367
R870 B.n77 B.n76 163.367
R871 B.n78 B.n77 163.367
R872 B.n680 B.n78 163.367
R873 B.n680 B.n83 163.367
R874 B.n84 B.n83 163.367
R875 B.n85 B.n84 163.367
R876 B.n685 B.n85 163.367
R877 B.n685 B.n90 163.367
R878 B.n91 B.n90 163.367
R879 B.n92 B.n91 163.367
R880 B.n690 B.n92 163.367
R881 B.n690 B.n97 163.367
R882 B.n98 B.n97 163.367
R883 B.n99 B.n98 163.367
R884 B.n695 B.n99 163.367
R885 B.n695 B.n104 163.367
R886 B.n360 B.n358 163.367
R887 B.n364 B.n358 163.367
R888 B.n368 B.n366 163.367
R889 B.n372 B.n356 163.367
R890 B.n376 B.n374 163.367
R891 B.n380 B.n354 163.367
R892 B.n384 B.n382 163.367
R893 B.n388 B.n352 163.367
R894 B.n392 B.n390 163.367
R895 B.n397 B.n348 163.367
R896 B.n401 B.n399 163.367
R897 B.n405 B.n346 163.367
R898 B.n409 B.n407 163.367
R899 B.n416 B.n344 163.367
R900 B.n420 B.n418 163.367
R901 B.n424 B.n342 163.367
R902 B.n428 B.n426 163.367
R903 B.n432 B.n340 163.367
R904 B.n436 B.n434 163.367
R905 B.n440 B.n338 163.367
R906 B.n444 B.n442 163.367
R907 B.n448 B.n336 163.367
R908 B.n452 B.n450 163.367
R909 B.n458 B.n330 163.367
R910 B.n462 B.n330 163.367
R911 B.n462 B.n324 163.367
R912 B.n470 B.n324 163.367
R913 B.n470 B.n322 163.367
R914 B.n474 B.n322 163.367
R915 B.n474 B.n316 163.367
R916 B.n482 B.n316 163.367
R917 B.n482 B.n314 163.367
R918 B.n486 B.n314 163.367
R919 B.n486 B.n308 163.367
R920 B.n494 B.n308 163.367
R921 B.n494 B.n306 163.367
R922 B.n498 B.n306 163.367
R923 B.n498 B.n300 163.367
R924 B.n506 B.n300 163.367
R925 B.n506 B.n298 163.367
R926 B.n510 B.n298 163.367
R927 B.n510 B.n292 163.367
R928 B.n519 B.n292 163.367
R929 B.n519 B.n290 163.367
R930 B.n523 B.n290 163.367
R931 B.n523 B.n285 163.367
R932 B.n531 B.n285 163.367
R933 B.n531 B.n283 163.367
R934 B.n535 B.n283 163.367
R935 B.n535 B.n277 163.367
R936 B.n543 B.n277 163.367
R937 B.n543 B.n275 163.367
R938 B.n547 B.n275 163.367
R939 B.n547 B.n269 163.367
R940 B.n555 B.n269 163.367
R941 B.n555 B.n267 163.367
R942 B.n559 B.n267 163.367
R943 B.n559 B.n261 163.367
R944 B.n567 B.n261 163.367
R945 B.n567 B.n259 163.367
R946 B.n571 B.n259 163.367
R947 B.n571 B.n253 163.367
R948 B.n579 B.n253 163.367
R949 B.n579 B.n251 163.367
R950 B.n583 B.n251 163.367
R951 B.n583 B.n245 163.367
R952 B.n591 B.n245 163.367
R953 B.n591 B.n243 163.367
R954 B.n595 B.n243 163.367
R955 B.n595 B.n237 163.367
R956 B.n603 B.n237 163.367
R957 B.n603 B.n235 163.367
R958 B.n607 B.n235 163.367
R959 B.n607 B.n229 163.367
R960 B.n616 B.n229 163.367
R961 B.n616 B.n227 163.367
R962 B.n620 B.n227 163.367
R963 B.n620 B.n3 163.367
R964 B.n815 B.n3 163.367
R965 B.n811 B.n2 163.367
R966 B.n811 B.n810 163.367
R967 B.n810 B.n9 163.367
R968 B.n806 B.n9 163.367
R969 B.n806 B.n11 163.367
R970 B.n802 B.n11 163.367
R971 B.n802 B.n17 163.367
R972 B.n798 B.n17 163.367
R973 B.n798 B.n19 163.367
R974 B.n794 B.n19 163.367
R975 B.n794 B.n24 163.367
R976 B.n790 B.n24 163.367
R977 B.n790 B.n26 163.367
R978 B.n786 B.n26 163.367
R979 B.n786 B.n31 163.367
R980 B.n782 B.n31 163.367
R981 B.n782 B.n33 163.367
R982 B.n778 B.n33 163.367
R983 B.n778 B.n38 163.367
R984 B.n774 B.n38 163.367
R985 B.n774 B.n40 163.367
R986 B.n770 B.n40 163.367
R987 B.n770 B.n45 163.367
R988 B.n766 B.n45 163.367
R989 B.n766 B.n47 163.367
R990 B.n762 B.n47 163.367
R991 B.n762 B.n52 163.367
R992 B.n758 B.n52 163.367
R993 B.n758 B.n54 163.367
R994 B.n754 B.n54 163.367
R995 B.n754 B.n59 163.367
R996 B.n750 B.n59 163.367
R997 B.n750 B.n61 163.367
R998 B.n746 B.n61 163.367
R999 B.n746 B.n65 163.367
R1000 B.n742 B.n65 163.367
R1001 B.n742 B.n67 163.367
R1002 B.n738 B.n67 163.367
R1003 B.n738 B.n73 163.367
R1004 B.n734 B.n73 163.367
R1005 B.n734 B.n75 163.367
R1006 B.n730 B.n75 163.367
R1007 B.n730 B.n80 163.367
R1008 B.n726 B.n80 163.367
R1009 B.n726 B.n82 163.367
R1010 B.n722 B.n82 163.367
R1011 B.n722 B.n87 163.367
R1012 B.n718 B.n87 163.367
R1013 B.n718 B.n89 163.367
R1014 B.n714 B.n89 163.367
R1015 B.n714 B.n94 163.367
R1016 B.n710 B.n94 163.367
R1017 B.n710 B.n96 163.367
R1018 B.n706 B.n96 163.367
R1019 B.n706 B.n101 163.367
R1020 B.n702 B.n101 163.367
R1021 B.n129 B.t17 136.155
R1022 B.n412 B.t21 136.155
R1023 B.n132 B.t14 136.151
R1024 B.n349 B.t11 136.151
R1025 B.n457 B.n333 131.883
R1026 B.n701 B.n700 131.883
R1027 B.n457 B.n329 79.3639
R1028 B.n463 B.n329 79.3639
R1029 B.n463 B.n325 79.3639
R1030 B.n469 B.n325 79.3639
R1031 B.n469 B.n321 79.3639
R1032 B.n475 B.n321 79.3639
R1033 B.n475 B.n317 79.3639
R1034 B.n481 B.n317 79.3639
R1035 B.n487 B.n313 79.3639
R1036 B.n487 B.n309 79.3639
R1037 B.n493 B.n309 79.3639
R1038 B.n493 B.n305 79.3639
R1039 B.n499 B.n305 79.3639
R1040 B.n499 B.n301 79.3639
R1041 B.n505 B.n301 79.3639
R1042 B.n505 B.n297 79.3639
R1043 B.n511 B.n297 79.3639
R1044 B.n511 B.n293 79.3639
R1045 B.n518 B.n293 79.3639
R1046 B.n518 B.n517 79.3639
R1047 B.n524 B.n286 79.3639
R1048 B.n530 B.n286 79.3639
R1049 B.n530 B.n282 79.3639
R1050 B.n536 B.n282 79.3639
R1051 B.n536 B.n278 79.3639
R1052 B.n542 B.n278 79.3639
R1053 B.n542 B.n274 79.3639
R1054 B.n548 B.n274 79.3639
R1055 B.n554 B.n270 79.3639
R1056 B.n554 B.n266 79.3639
R1057 B.n560 B.n266 79.3639
R1058 B.n560 B.n262 79.3639
R1059 B.n566 B.n262 79.3639
R1060 B.n566 B.n258 79.3639
R1061 B.n572 B.n258 79.3639
R1062 B.n572 B.n254 79.3639
R1063 B.n578 B.n254 79.3639
R1064 B.n584 B.n250 79.3639
R1065 B.n584 B.n246 79.3639
R1066 B.n590 B.n246 79.3639
R1067 B.n590 B.n242 79.3639
R1068 B.n596 B.n242 79.3639
R1069 B.n596 B.n238 79.3639
R1070 B.n602 B.n238 79.3639
R1071 B.n602 B.n234 79.3639
R1072 B.n608 B.n234 79.3639
R1073 B.n615 B.n230 79.3639
R1074 B.n615 B.n226 79.3639
R1075 B.n621 B.n226 79.3639
R1076 B.n621 B.n4 79.3639
R1077 B.n814 B.n4 79.3639
R1078 B.n814 B.n813 79.3639
R1079 B.n813 B.n812 79.3639
R1080 B.n812 B.n8 79.3639
R1081 B.n12 B.n8 79.3639
R1082 B.n805 B.n12 79.3639
R1083 B.n805 B.n804 79.3639
R1084 B.n803 B.n16 79.3639
R1085 B.n797 B.n16 79.3639
R1086 B.n797 B.n796 79.3639
R1087 B.n796 B.n795 79.3639
R1088 B.n795 B.n23 79.3639
R1089 B.n789 B.n23 79.3639
R1090 B.n789 B.n788 79.3639
R1091 B.n788 B.n787 79.3639
R1092 B.n787 B.n30 79.3639
R1093 B.n781 B.n780 79.3639
R1094 B.n780 B.n779 79.3639
R1095 B.n779 B.n37 79.3639
R1096 B.n773 B.n37 79.3639
R1097 B.n773 B.n772 79.3639
R1098 B.n772 B.n771 79.3639
R1099 B.n771 B.n44 79.3639
R1100 B.n765 B.n44 79.3639
R1101 B.n765 B.n764 79.3639
R1102 B.n763 B.n51 79.3639
R1103 B.n757 B.n51 79.3639
R1104 B.n757 B.n756 79.3639
R1105 B.n756 B.n755 79.3639
R1106 B.n755 B.n58 79.3639
R1107 B.n749 B.n58 79.3639
R1108 B.n749 B.n748 79.3639
R1109 B.n748 B.n747 79.3639
R1110 B.n741 B.n68 79.3639
R1111 B.n741 B.n740 79.3639
R1112 B.n740 B.n739 79.3639
R1113 B.n739 B.n72 79.3639
R1114 B.n733 B.n72 79.3639
R1115 B.n733 B.n732 79.3639
R1116 B.n732 B.n731 79.3639
R1117 B.n731 B.n79 79.3639
R1118 B.n725 B.n79 79.3639
R1119 B.n725 B.n724 79.3639
R1120 B.n724 B.n723 79.3639
R1121 B.n723 B.n86 79.3639
R1122 B.n717 B.n716 79.3639
R1123 B.n716 B.n715 79.3639
R1124 B.n715 B.n93 79.3639
R1125 B.n709 B.n93 79.3639
R1126 B.n709 B.n708 79.3639
R1127 B.n708 B.n707 79.3639
R1128 B.n707 B.n100 79.3639
R1129 B.n701 B.n100 79.3639
R1130 B.t5 B.n230 73.5284
R1131 B.n804 B.t1 73.5284
R1132 B.n130 B.t18 72.5432
R1133 B.n413 B.t20 72.5432
R1134 B.n133 B.t15 72.5393
R1135 B.n350 B.t10 72.5393
R1136 B.n105 B.n103 71.676
R1137 B.n136 B.n106 71.676
R1138 B.n140 B.n107 71.676
R1139 B.n144 B.n108 71.676
R1140 B.n148 B.n109 71.676
R1141 B.n152 B.n110 71.676
R1142 B.n156 B.n111 71.676
R1143 B.n160 B.n112 71.676
R1144 B.n164 B.n113 71.676
R1145 B.n168 B.n114 71.676
R1146 B.n173 B.n115 71.676
R1147 B.n177 B.n116 71.676
R1148 B.n181 B.n117 71.676
R1149 B.n185 B.n118 71.676
R1150 B.n189 B.n119 71.676
R1151 B.n193 B.n120 71.676
R1152 B.n197 B.n121 71.676
R1153 B.n201 B.n122 71.676
R1154 B.n205 B.n123 71.676
R1155 B.n209 B.n124 71.676
R1156 B.n213 B.n125 71.676
R1157 B.n217 B.n126 71.676
R1158 B.n221 B.n127 71.676
R1159 B.n128 B.n127 71.676
R1160 B.n220 B.n126 71.676
R1161 B.n216 B.n125 71.676
R1162 B.n212 B.n124 71.676
R1163 B.n208 B.n123 71.676
R1164 B.n204 B.n122 71.676
R1165 B.n200 B.n121 71.676
R1166 B.n196 B.n120 71.676
R1167 B.n192 B.n119 71.676
R1168 B.n188 B.n118 71.676
R1169 B.n184 B.n117 71.676
R1170 B.n180 B.n116 71.676
R1171 B.n176 B.n115 71.676
R1172 B.n172 B.n114 71.676
R1173 B.n167 B.n113 71.676
R1174 B.n163 B.n112 71.676
R1175 B.n159 B.n111 71.676
R1176 B.n155 B.n110 71.676
R1177 B.n151 B.n109 71.676
R1178 B.n147 B.n108 71.676
R1179 B.n143 B.n107 71.676
R1180 B.n139 B.n106 71.676
R1181 B.n135 B.n105 71.676
R1182 B.n359 B.n332 71.676
R1183 B.n365 B.n364 71.676
R1184 B.n368 B.n367 71.676
R1185 B.n373 B.n372 71.676
R1186 B.n376 B.n375 71.676
R1187 B.n381 B.n380 71.676
R1188 B.n384 B.n383 71.676
R1189 B.n389 B.n388 71.676
R1190 B.n392 B.n391 71.676
R1191 B.n398 B.n397 71.676
R1192 B.n401 B.n400 71.676
R1193 B.n406 B.n405 71.676
R1194 B.n409 B.n408 71.676
R1195 B.n417 B.n416 71.676
R1196 B.n420 B.n419 71.676
R1197 B.n425 B.n424 71.676
R1198 B.n428 B.n427 71.676
R1199 B.n433 B.n432 71.676
R1200 B.n436 B.n435 71.676
R1201 B.n441 B.n440 71.676
R1202 B.n444 B.n443 71.676
R1203 B.n449 B.n448 71.676
R1204 B.n452 B.n451 71.676
R1205 B.n360 B.n359 71.676
R1206 B.n366 B.n365 71.676
R1207 B.n367 B.n356 71.676
R1208 B.n374 B.n373 71.676
R1209 B.n375 B.n354 71.676
R1210 B.n382 B.n381 71.676
R1211 B.n383 B.n352 71.676
R1212 B.n390 B.n389 71.676
R1213 B.n391 B.n348 71.676
R1214 B.n399 B.n398 71.676
R1215 B.n400 B.n346 71.676
R1216 B.n407 B.n406 71.676
R1217 B.n408 B.n344 71.676
R1218 B.n418 B.n417 71.676
R1219 B.n419 B.n342 71.676
R1220 B.n426 B.n425 71.676
R1221 B.n427 B.n340 71.676
R1222 B.n434 B.n433 71.676
R1223 B.n435 B.n338 71.676
R1224 B.n442 B.n441 71.676
R1225 B.n443 B.n336 71.676
R1226 B.n450 B.n449 71.676
R1227 B.n451 B.n334 71.676
R1228 B.n816 B.n815 71.676
R1229 B.n816 B.n2 71.676
R1230 B.n524 B.t0 68.8599
R1231 B.n747 B.t2 68.8599
R1232 B.n133 B.n132 63.6126
R1233 B.n130 B.n129 63.6126
R1234 B.n413 B.n412 63.6126
R1235 B.n350 B.n349 63.6126
R1236 B.n548 B.t7 61.8573
R1237 B.t6 B.n763 61.8573
R1238 B.n170 B.n133 59.5399
R1239 B.n131 B.n130 59.5399
R1240 B.n414 B.n413 59.5399
R1241 B.n395 B.n350 59.5399
R1242 B.t9 B.n313 57.1888
R1243 B.t13 B.n86 57.1888
R1244 B.t3 B.n250 45.5177
R1245 B.t4 B.n30 45.5177
R1246 B.n578 B.t3 33.8467
R1247 B.n781 B.t4 33.8467
R1248 B.n459 B.n331 28.8785
R1249 B.n455 B.n454 28.8785
R1250 B.n698 B.n697 28.8785
R1251 B.n703 B.n102 28.8785
R1252 B.n481 B.t9 22.1756
R1253 B.n717 B.t13 22.1756
R1254 B B.n817 18.0485
R1255 B.t7 B.n270 17.5071
R1256 B.n764 B.t6 17.5071
R1257 B.n460 B.n459 10.6151
R1258 B.n461 B.n460 10.6151
R1259 B.n461 B.n323 10.6151
R1260 B.n471 B.n323 10.6151
R1261 B.n472 B.n471 10.6151
R1262 B.n473 B.n472 10.6151
R1263 B.n473 B.n315 10.6151
R1264 B.n483 B.n315 10.6151
R1265 B.n484 B.n483 10.6151
R1266 B.n485 B.n484 10.6151
R1267 B.n485 B.n307 10.6151
R1268 B.n495 B.n307 10.6151
R1269 B.n496 B.n495 10.6151
R1270 B.n497 B.n496 10.6151
R1271 B.n497 B.n299 10.6151
R1272 B.n507 B.n299 10.6151
R1273 B.n508 B.n507 10.6151
R1274 B.n509 B.n508 10.6151
R1275 B.n509 B.n291 10.6151
R1276 B.n520 B.n291 10.6151
R1277 B.n521 B.n520 10.6151
R1278 B.n522 B.n521 10.6151
R1279 B.n522 B.n284 10.6151
R1280 B.n532 B.n284 10.6151
R1281 B.n533 B.n532 10.6151
R1282 B.n534 B.n533 10.6151
R1283 B.n534 B.n276 10.6151
R1284 B.n544 B.n276 10.6151
R1285 B.n545 B.n544 10.6151
R1286 B.n546 B.n545 10.6151
R1287 B.n546 B.n268 10.6151
R1288 B.n556 B.n268 10.6151
R1289 B.n557 B.n556 10.6151
R1290 B.n558 B.n557 10.6151
R1291 B.n558 B.n260 10.6151
R1292 B.n568 B.n260 10.6151
R1293 B.n569 B.n568 10.6151
R1294 B.n570 B.n569 10.6151
R1295 B.n570 B.n252 10.6151
R1296 B.n580 B.n252 10.6151
R1297 B.n581 B.n580 10.6151
R1298 B.n582 B.n581 10.6151
R1299 B.n582 B.n244 10.6151
R1300 B.n592 B.n244 10.6151
R1301 B.n593 B.n592 10.6151
R1302 B.n594 B.n593 10.6151
R1303 B.n594 B.n236 10.6151
R1304 B.n604 B.n236 10.6151
R1305 B.n605 B.n604 10.6151
R1306 B.n606 B.n605 10.6151
R1307 B.n606 B.n228 10.6151
R1308 B.n617 B.n228 10.6151
R1309 B.n618 B.n617 10.6151
R1310 B.n619 B.n618 10.6151
R1311 B.n619 B.n0 10.6151
R1312 B.n361 B.n331 10.6151
R1313 B.n362 B.n361 10.6151
R1314 B.n363 B.n362 10.6151
R1315 B.n363 B.n357 10.6151
R1316 B.n369 B.n357 10.6151
R1317 B.n370 B.n369 10.6151
R1318 B.n371 B.n370 10.6151
R1319 B.n371 B.n355 10.6151
R1320 B.n377 B.n355 10.6151
R1321 B.n378 B.n377 10.6151
R1322 B.n379 B.n378 10.6151
R1323 B.n379 B.n353 10.6151
R1324 B.n385 B.n353 10.6151
R1325 B.n386 B.n385 10.6151
R1326 B.n387 B.n386 10.6151
R1327 B.n387 B.n351 10.6151
R1328 B.n393 B.n351 10.6151
R1329 B.n394 B.n393 10.6151
R1330 B.n396 B.n347 10.6151
R1331 B.n402 B.n347 10.6151
R1332 B.n403 B.n402 10.6151
R1333 B.n404 B.n403 10.6151
R1334 B.n404 B.n345 10.6151
R1335 B.n410 B.n345 10.6151
R1336 B.n411 B.n410 10.6151
R1337 B.n415 B.n411 10.6151
R1338 B.n421 B.n343 10.6151
R1339 B.n422 B.n421 10.6151
R1340 B.n423 B.n422 10.6151
R1341 B.n423 B.n341 10.6151
R1342 B.n429 B.n341 10.6151
R1343 B.n430 B.n429 10.6151
R1344 B.n431 B.n430 10.6151
R1345 B.n431 B.n339 10.6151
R1346 B.n437 B.n339 10.6151
R1347 B.n438 B.n437 10.6151
R1348 B.n439 B.n438 10.6151
R1349 B.n439 B.n337 10.6151
R1350 B.n445 B.n337 10.6151
R1351 B.n446 B.n445 10.6151
R1352 B.n447 B.n446 10.6151
R1353 B.n447 B.n335 10.6151
R1354 B.n453 B.n335 10.6151
R1355 B.n454 B.n453 10.6151
R1356 B.n455 B.n327 10.6151
R1357 B.n465 B.n327 10.6151
R1358 B.n466 B.n465 10.6151
R1359 B.n467 B.n466 10.6151
R1360 B.n467 B.n319 10.6151
R1361 B.n477 B.n319 10.6151
R1362 B.n478 B.n477 10.6151
R1363 B.n479 B.n478 10.6151
R1364 B.n479 B.n311 10.6151
R1365 B.n489 B.n311 10.6151
R1366 B.n490 B.n489 10.6151
R1367 B.n491 B.n490 10.6151
R1368 B.n491 B.n303 10.6151
R1369 B.n501 B.n303 10.6151
R1370 B.n502 B.n501 10.6151
R1371 B.n503 B.n502 10.6151
R1372 B.n503 B.n295 10.6151
R1373 B.n513 B.n295 10.6151
R1374 B.n514 B.n513 10.6151
R1375 B.n515 B.n514 10.6151
R1376 B.n515 B.n288 10.6151
R1377 B.n526 B.n288 10.6151
R1378 B.n527 B.n526 10.6151
R1379 B.n528 B.n527 10.6151
R1380 B.n528 B.n280 10.6151
R1381 B.n538 B.n280 10.6151
R1382 B.n539 B.n538 10.6151
R1383 B.n540 B.n539 10.6151
R1384 B.n540 B.n272 10.6151
R1385 B.n550 B.n272 10.6151
R1386 B.n551 B.n550 10.6151
R1387 B.n552 B.n551 10.6151
R1388 B.n552 B.n264 10.6151
R1389 B.n562 B.n264 10.6151
R1390 B.n563 B.n562 10.6151
R1391 B.n564 B.n563 10.6151
R1392 B.n564 B.n256 10.6151
R1393 B.n574 B.n256 10.6151
R1394 B.n575 B.n574 10.6151
R1395 B.n576 B.n575 10.6151
R1396 B.n576 B.n248 10.6151
R1397 B.n586 B.n248 10.6151
R1398 B.n587 B.n586 10.6151
R1399 B.n588 B.n587 10.6151
R1400 B.n588 B.n240 10.6151
R1401 B.n598 B.n240 10.6151
R1402 B.n599 B.n598 10.6151
R1403 B.n600 B.n599 10.6151
R1404 B.n600 B.n232 10.6151
R1405 B.n610 B.n232 10.6151
R1406 B.n611 B.n610 10.6151
R1407 B.n613 B.n611 10.6151
R1408 B.n613 B.n612 10.6151
R1409 B.n612 B.n224 10.6151
R1410 B.n624 B.n224 10.6151
R1411 B.n625 B.n624 10.6151
R1412 B.n626 B.n625 10.6151
R1413 B.n627 B.n626 10.6151
R1414 B.n628 B.n627 10.6151
R1415 B.n631 B.n628 10.6151
R1416 B.n632 B.n631 10.6151
R1417 B.n633 B.n632 10.6151
R1418 B.n634 B.n633 10.6151
R1419 B.n636 B.n634 10.6151
R1420 B.n637 B.n636 10.6151
R1421 B.n638 B.n637 10.6151
R1422 B.n639 B.n638 10.6151
R1423 B.n641 B.n639 10.6151
R1424 B.n642 B.n641 10.6151
R1425 B.n643 B.n642 10.6151
R1426 B.n644 B.n643 10.6151
R1427 B.n646 B.n644 10.6151
R1428 B.n647 B.n646 10.6151
R1429 B.n648 B.n647 10.6151
R1430 B.n649 B.n648 10.6151
R1431 B.n651 B.n649 10.6151
R1432 B.n652 B.n651 10.6151
R1433 B.n653 B.n652 10.6151
R1434 B.n654 B.n653 10.6151
R1435 B.n656 B.n654 10.6151
R1436 B.n657 B.n656 10.6151
R1437 B.n658 B.n657 10.6151
R1438 B.n659 B.n658 10.6151
R1439 B.n661 B.n659 10.6151
R1440 B.n662 B.n661 10.6151
R1441 B.n663 B.n662 10.6151
R1442 B.n664 B.n663 10.6151
R1443 B.n666 B.n664 10.6151
R1444 B.n667 B.n666 10.6151
R1445 B.n668 B.n667 10.6151
R1446 B.n669 B.n668 10.6151
R1447 B.n671 B.n669 10.6151
R1448 B.n672 B.n671 10.6151
R1449 B.n673 B.n672 10.6151
R1450 B.n674 B.n673 10.6151
R1451 B.n676 B.n674 10.6151
R1452 B.n677 B.n676 10.6151
R1453 B.n678 B.n677 10.6151
R1454 B.n679 B.n678 10.6151
R1455 B.n681 B.n679 10.6151
R1456 B.n682 B.n681 10.6151
R1457 B.n683 B.n682 10.6151
R1458 B.n684 B.n683 10.6151
R1459 B.n686 B.n684 10.6151
R1460 B.n687 B.n686 10.6151
R1461 B.n688 B.n687 10.6151
R1462 B.n689 B.n688 10.6151
R1463 B.n691 B.n689 10.6151
R1464 B.n692 B.n691 10.6151
R1465 B.n693 B.n692 10.6151
R1466 B.n694 B.n693 10.6151
R1467 B.n696 B.n694 10.6151
R1468 B.n697 B.n696 10.6151
R1469 B.n809 B.n1 10.6151
R1470 B.n809 B.n808 10.6151
R1471 B.n808 B.n807 10.6151
R1472 B.n807 B.n10 10.6151
R1473 B.n801 B.n10 10.6151
R1474 B.n801 B.n800 10.6151
R1475 B.n800 B.n799 10.6151
R1476 B.n799 B.n18 10.6151
R1477 B.n793 B.n18 10.6151
R1478 B.n793 B.n792 10.6151
R1479 B.n792 B.n791 10.6151
R1480 B.n791 B.n25 10.6151
R1481 B.n785 B.n25 10.6151
R1482 B.n785 B.n784 10.6151
R1483 B.n784 B.n783 10.6151
R1484 B.n783 B.n32 10.6151
R1485 B.n777 B.n32 10.6151
R1486 B.n777 B.n776 10.6151
R1487 B.n776 B.n775 10.6151
R1488 B.n775 B.n39 10.6151
R1489 B.n769 B.n39 10.6151
R1490 B.n769 B.n768 10.6151
R1491 B.n768 B.n767 10.6151
R1492 B.n767 B.n46 10.6151
R1493 B.n761 B.n46 10.6151
R1494 B.n761 B.n760 10.6151
R1495 B.n760 B.n759 10.6151
R1496 B.n759 B.n53 10.6151
R1497 B.n753 B.n53 10.6151
R1498 B.n753 B.n752 10.6151
R1499 B.n752 B.n751 10.6151
R1500 B.n751 B.n60 10.6151
R1501 B.n745 B.n60 10.6151
R1502 B.n745 B.n744 10.6151
R1503 B.n744 B.n743 10.6151
R1504 B.n743 B.n66 10.6151
R1505 B.n737 B.n66 10.6151
R1506 B.n737 B.n736 10.6151
R1507 B.n736 B.n735 10.6151
R1508 B.n735 B.n74 10.6151
R1509 B.n729 B.n74 10.6151
R1510 B.n729 B.n728 10.6151
R1511 B.n728 B.n727 10.6151
R1512 B.n727 B.n81 10.6151
R1513 B.n721 B.n81 10.6151
R1514 B.n721 B.n720 10.6151
R1515 B.n720 B.n719 10.6151
R1516 B.n719 B.n88 10.6151
R1517 B.n713 B.n88 10.6151
R1518 B.n713 B.n712 10.6151
R1519 B.n712 B.n711 10.6151
R1520 B.n711 B.n95 10.6151
R1521 B.n705 B.n95 10.6151
R1522 B.n705 B.n704 10.6151
R1523 B.n704 B.n703 10.6151
R1524 B.n134 B.n102 10.6151
R1525 B.n137 B.n134 10.6151
R1526 B.n138 B.n137 10.6151
R1527 B.n141 B.n138 10.6151
R1528 B.n142 B.n141 10.6151
R1529 B.n145 B.n142 10.6151
R1530 B.n146 B.n145 10.6151
R1531 B.n149 B.n146 10.6151
R1532 B.n150 B.n149 10.6151
R1533 B.n153 B.n150 10.6151
R1534 B.n154 B.n153 10.6151
R1535 B.n157 B.n154 10.6151
R1536 B.n158 B.n157 10.6151
R1537 B.n161 B.n158 10.6151
R1538 B.n162 B.n161 10.6151
R1539 B.n165 B.n162 10.6151
R1540 B.n166 B.n165 10.6151
R1541 B.n169 B.n166 10.6151
R1542 B.n174 B.n171 10.6151
R1543 B.n175 B.n174 10.6151
R1544 B.n178 B.n175 10.6151
R1545 B.n179 B.n178 10.6151
R1546 B.n182 B.n179 10.6151
R1547 B.n183 B.n182 10.6151
R1548 B.n186 B.n183 10.6151
R1549 B.n187 B.n186 10.6151
R1550 B.n191 B.n190 10.6151
R1551 B.n194 B.n191 10.6151
R1552 B.n195 B.n194 10.6151
R1553 B.n198 B.n195 10.6151
R1554 B.n199 B.n198 10.6151
R1555 B.n202 B.n199 10.6151
R1556 B.n203 B.n202 10.6151
R1557 B.n206 B.n203 10.6151
R1558 B.n207 B.n206 10.6151
R1559 B.n210 B.n207 10.6151
R1560 B.n211 B.n210 10.6151
R1561 B.n214 B.n211 10.6151
R1562 B.n215 B.n214 10.6151
R1563 B.n218 B.n215 10.6151
R1564 B.n219 B.n218 10.6151
R1565 B.n222 B.n219 10.6151
R1566 B.n223 B.n222 10.6151
R1567 B.n698 B.n223 10.6151
R1568 B.n517 B.t0 10.5045
R1569 B.n68 B.t2 10.5045
R1570 B.n817 B.n0 8.11757
R1571 B.n817 B.n1 8.11757
R1572 B.n396 B.n395 6.5566
R1573 B.n415 B.n414 6.5566
R1574 B.n171 B.n170 6.5566
R1575 B.n187 B.n131 6.5566
R1576 B.n608 B.t5 5.83604
R1577 B.t1 B.n803 5.83604
R1578 B.n395 B.n394 4.05904
R1579 B.n414 B.n343 4.05904
R1580 B.n170 B.n169 4.05904
R1581 B.n190 B.n131 4.05904
R1582 VP.n21 VP.n20 161.3
R1583 VP.n22 VP.n17 161.3
R1584 VP.n24 VP.n23 161.3
R1585 VP.n25 VP.n16 161.3
R1586 VP.n27 VP.n26 161.3
R1587 VP.n28 VP.n15 161.3
R1588 VP.n30 VP.n29 161.3
R1589 VP.n32 VP.n14 161.3
R1590 VP.n34 VP.n33 161.3
R1591 VP.n35 VP.n13 161.3
R1592 VP.n37 VP.n36 161.3
R1593 VP.n38 VP.n12 161.3
R1594 VP.n40 VP.n39 161.3
R1595 VP.n73 VP.n72 161.3
R1596 VP.n71 VP.n1 161.3
R1597 VP.n70 VP.n69 161.3
R1598 VP.n68 VP.n2 161.3
R1599 VP.n67 VP.n66 161.3
R1600 VP.n65 VP.n3 161.3
R1601 VP.n63 VP.n62 161.3
R1602 VP.n61 VP.n4 161.3
R1603 VP.n60 VP.n59 161.3
R1604 VP.n58 VP.n5 161.3
R1605 VP.n57 VP.n56 161.3
R1606 VP.n55 VP.n6 161.3
R1607 VP.n54 VP.n53 161.3
R1608 VP.n51 VP.n7 161.3
R1609 VP.n50 VP.n49 161.3
R1610 VP.n48 VP.n8 161.3
R1611 VP.n47 VP.n46 161.3
R1612 VP.n45 VP.n9 161.3
R1613 VP.n44 VP.n43 161.3
R1614 VP.n42 VP.n10 69.5151
R1615 VP.n74 VP.n0 69.5151
R1616 VP.n41 VP.n11 69.5151
R1617 VP.n19 VP.n18 66.8452
R1618 VP.n18 VP.t7 65.6239
R1619 VP.n46 VP.n8 56.5193
R1620 VP.n70 VP.n2 56.5193
R1621 VP.n37 VP.n13 56.5193
R1622 VP.n42 VP.n41 46.7039
R1623 VP.n58 VP.n57 40.4934
R1624 VP.n59 VP.n58 40.4934
R1625 VP.n26 VP.n25 40.4934
R1626 VP.n25 VP.n24 40.4934
R1627 VP.n10 VP.t3 33.9039
R1628 VP.n52 VP.t1 33.9039
R1629 VP.n64 VP.t0 33.9039
R1630 VP.n0 VP.t2 33.9039
R1631 VP.n11 VP.t4 33.9039
R1632 VP.n31 VP.t5 33.9039
R1633 VP.n19 VP.t6 33.9039
R1634 VP.n45 VP.n44 24.4675
R1635 VP.n46 VP.n45 24.4675
R1636 VP.n50 VP.n8 24.4675
R1637 VP.n51 VP.n50 24.4675
R1638 VP.n53 VP.n6 24.4675
R1639 VP.n57 VP.n6 24.4675
R1640 VP.n59 VP.n4 24.4675
R1641 VP.n63 VP.n4 24.4675
R1642 VP.n66 VP.n65 24.4675
R1643 VP.n66 VP.n2 24.4675
R1644 VP.n71 VP.n70 24.4675
R1645 VP.n72 VP.n71 24.4675
R1646 VP.n38 VP.n37 24.4675
R1647 VP.n39 VP.n38 24.4675
R1648 VP.n26 VP.n15 24.4675
R1649 VP.n30 VP.n15 24.4675
R1650 VP.n33 VP.n32 24.4675
R1651 VP.n33 VP.n13 24.4675
R1652 VP.n20 VP.n17 24.4675
R1653 VP.n24 VP.n17 24.4675
R1654 VP.n44 VP.n10 20.5528
R1655 VP.n72 VP.n0 20.5528
R1656 VP.n39 VP.n11 20.5528
R1657 VP.n52 VP.n51 17.6167
R1658 VP.n65 VP.n64 17.6167
R1659 VP.n32 VP.n31 17.6167
R1660 VP.n53 VP.n52 6.85126
R1661 VP.n64 VP.n63 6.85126
R1662 VP.n31 VP.n30 6.85126
R1663 VP.n20 VP.n19 6.85126
R1664 VP.n21 VP.n18 5.514
R1665 VP.n41 VP.n40 0.354971
R1666 VP.n43 VP.n42 0.354971
R1667 VP.n74 VP.n73 0.354971
R1668 VP VP.n74 0.26696
R1669 VP.n22 VP.n21 0.189894
R1670 VP.n23 VP.n22 0.189894
R1671 VP.n23 VP.n16 0.189894
R1672 VP.n27 VP.n16 0.189894
R1673 VP.n28 VP.n27 0.189894
R1674 VP.n29 VP.n28 0.189894
R1675 VP.n29 VP.n14 0.189894
R1676 VP.n34 VP.n14 0.189894
R1677 VP.n35 VP.n34 0.189894
R1678 VP.n36 VP.n35 0.189894
R1679 VP.n36 VP.n12 0.189894
R1680 VP.n40 VP.n12 0.189894
R1681 VP.n43 VP.n9 0.189894
R1682 VP.n47 VP.n9 0.189894
R1683 VP.n48 VP.n47 0.189894
R1684 VP.n49 VP.n48 0.189894
R1685 VP.n49 VP.n7 0.189894
R1686 VP.n54 VP.n7 0.189894
R1687 VP.n55 VP.n54 0.189894
R1688 VP.n56 VP.n55 0.189894
R1689 VP.n56 VP.n5 0.189894
R1690 VP.n60 VP.n5 0.189894
R1691 VP.n61 VP.n60 0.189894
R1692 VP.n62 VP.n61 0.189894
R1693 VP.n62 VP.n3 0.189894
R1694 VP.n67 VP.n3 0.189894
R1695 VP.n68 VP.n67 0.189894
R1696 VP.n69 VP.n68 0.189894
R1697 VP.n69 VP.n1 0.189894
R1698 VP.n73 VP.n1 0.189894
R1699 VDD1 VDD1.n0 72.4207
R1700 VDD1.n3 VDD1.n2 72.307
R1701 VDD1.n3 VDD1.n1 72.307
R1702 VDD1.n5 VDD1.n4 70.9486
R1703 VDD1.n5 VDD1.n3 40.6
R1704 VDD1.n4 VDD1.t2 4.77158
R1705 VDD1.n4 VDD1.t3 4.77158
R1706 VDD1.n0 VDD1.t0 4.77158
R1707 VDD1.n0 VDD1.t1 4.77158
R1708 VDD1.n2 VDD1.t7 4.77158
R1709 VDD1.n2 VDD1.t5 4.77158
R1710 VDD1.n1 VDD1.t4 4.77158
R1711 VDD1.n1 VDD1.t6 4.77158
R1712 VDD1 VDD1.n5 1.3561
C0 VP VDD1 3.77862f
C1 VDD2 VN 3.37578f
C2 VDD1 VTAIL 5.70579f
C3 VP VN 6.64513f
C4 VDD2 VP 0.561849f
C5 VTAIL VN 4.48093f
C6 VDD2 VTAIL 5.76255f
C7 VP VTAIL 4.49504f
C8 VDD1 VN 0.15669f
C9 VDD2 VDD1 1.96053f
C10 VDD2 B 5.058959f
C11 VDD1 B 5.540306f
C12 VTAIL B 5.566135f
C13 VN B 16.11706f
C14 VP B 14.697908f
C15 VDD1.t0 B 0.081421f
C16 VDD1.t1 B 0.081421f
C17 VDD1.n0 B 0.655647f
C18 VDD1.t4 B 0.081421f
C19 VDD1.t6 B 0.081421f
C20 VDD1.n1 B 0.65464f
C21 VDD1.t7 B 0.081421f
C22 VDD1.t5 B 0.081421f
C23 VDD1.n2 B 0.65464f
C24 VDD1.n3 B 3.00933f
C25 VDD1.t2 B 0.081421f
C26 VDD1.t3 B 0.081421f
C27 VDD1.n4 B 0.644519f
C28 VDD1.n5 B 2.46742f
C29 VP.t2 B 0.810497f
C30 VP.n0 B 0.418347f
C31 VP.n1 B 0.025687f
C32 VP.n2 B 0.039645f
C33 VP.n3 B 0.025687f
C34 VP.t0 B 0.810497f
C35 VP.n4 B 0.047873f
C36 VP.n5 B 0.025687f
C37 VP.n6 B 0.047873f
C38 VP.n7 B 0.025687f
C39 VP.t1 B 0.810497f
C40 VP.n8 B 0.039645f
C41 VP.n9 B 0.025687f
C42 VP.t3 B 0.810497f
C43 VP.n10 B 0.418347f
C44 VP.t4 B 0.810497f
C45 VP.n11 B 0.418347f
C46 VP.n12 B 0.025687f
C47 VP.n13 B 0.039645f
C48 VP.n14 B 0.025687f
C49 VP.t5 B 0.810497f
C50 VP.n15 B 0.047873f
C51 VP.n16 B 0.025687f
C52 VP.n17 B 0.047873f
C53 VP.t7 B 1.04631f
C54 VP.n18 B 0.384628f
C55 VP.t6 B 0.810497f
C56 VP.n19 B 0.393284f
C57 VP.n20 B 0.030856f
C58 VP.n21 B 0.276088f
C59 VP.n22 B 0.025687f
C60 VP.n23 B 0.025687f
C61 VP.n24 B 0.051052f
C62 VP.n25 B 0.020765f
C63 VP.n26 B 0.051052f
C64 VP.n27 B 0.025687f
C65 VP.n28 B 0.025687f
C66 VP.n29 B 0.025687f
C67 VP.n30 B 0.030856f
C68 VP.n31 B 0.317396f
C69 VP.n32 B 0.041255f
C70 VP.n33 B 0.047873f
C71 VP.n34 B 0.025687f
C72 VP.n35 B 0.025687f
C73 VP.n36 B 0.025687f
C74 VP.n37 B 0.03535f
C75 VP.n38 B 0.047873f
C76 VP.n39 B 0.044092f
C77 VP.n40 B 0.041457f
C78 VP.n41 B 1.31215f
C79 VP.n42 B 1.33192f
C80 VP.n43 B 0.041457f
C81 VP.n44 B 0.044092f
C82 VP.n45 B 0.047873f
C83 VP.n46 B 0.03535f
C84 VP.n47 B 0.025687f
C85 VP.n48 B 0.025687f
C86 VP.n49 B 0.025687f
C87 VP.n50 B 0.047873f
C88 VP.n51 B 0.041255f
C89 VP.n52 B 0.317396f
C90 VP.n53 B 0.030856f
C91 VP.n54 B 0.025687f
C92 VP.n55 B 0.025687f
C93 VP.n56 B 0.025687f
C94 VP.n57 B 0.051052f
C95 VP.n58 B 0.020765f
C96 VP.n59 B 0.051052f
C97 VP.n60 B 0.025687f
C98 VP.n61 B 0.025687f
C99 VP.n62 B 0.025687f
C100 VP.n63 B 0.030856f
C101 VP.n64 B 0.317396f
C102 VP.n65 B 0.041255f
C103 VP.n66 B 0.047873f
C104 VP.n67 B 0.025687f
C105 VP.n68 B 0.025687f
C106 VP.n69 B 0.025687f
C107 VP.n70 B 0.03535f
C108 VP.n71 B 0.047873f
C109 VP.n72 B 0.044092f
C110 VP.n73 B 0.041457f
C111 VP.n74 B 0.052396f
C112 VDD2.t5 B 0.079619f
C113 VDD2.t7 B 0.079619f
C114 VDD2.n0 B 0.640147f
C115 VDD2.t6 B 0.079619f
C116 VDD2.t2 B 0.079619f
C117 VDD2.n1 B 0.640147f
C118 VDD2.n2 B 2.89213f
C119 VDD2.t1 B 0.079619f
C120 VDD2.t0 B 0.079619f
C121 VDD2.n3 B 0.630252f
C122 VDD2.n4 B 2.3828f
C123 VDD2.t3 B 0.079619f
C124 VDD2.t4 B 0.079619f
C125 VDD2.n5 B 0.640114f
C126 VTAIL.t8 B 0.086726f
C127 VTAIL.t10 B 0.086726f
C128 VTAIL.n0 B 0.62475f
C129 VTAIL.n1 B 0.477708f
C130 VTAIL.t11 B 0.798682f
C131 VTAIL.n2 B 0.575376f
C132 VTAIL.t5 B 0.798682f
C133 VTAIL.n3 B 0.575376f
C134 VTAIL.t7 B 0.086726f
C135 VTAIL.t3 B 0.086726f
C136 VTAIL.n4 B 0.62475f
C137 VTAIL.n5 B 0.713694f
C138 VTAIL.t0 B 0.798682f
C139 VTAIL.n6 B 1.44036f
C140 VTAIL.t14 B 0.798686f
C141 VTAIL.n7 B 1.44036f
C142 VTAIL.t15 B 0.086726f
C143 VTAIL.t9 B 0.086726f
C144 VTAIL.n8 B 0.624753f
C145 VTAIL.n9 B 0.71369f
C146 VTAIL.t12 B 0.798686f
C147 VTAIL.n10 B 0.575372f
C148 VTAIL.t1 B 0.798686f
C149 VTAIL.n11 B 0.575372f
C150 VTAIL.t4 B 0.086726f
C151 VTAIL.t6 B 0.086726f
C152 VTAIL.n12 B 0.624753f
C153 VTAIL.n13 B 0.71369f
C154 VTAIL.t2 B 0.798682f
C155 VTAIL.n14 B 1.44036f
C156 VTAIL.t13 B 0.798682f
C157 VTAIL.n15 B 1.43541f
C158 VN.t5 B 0.786832f
C159 VN.n0 B 0.406132f
C160 VN.n1 B 0.024937f
C161 VN.n2 B 0.038487f
C162 VN.n3 B 0.024937f
C163 VN.t1 B 0.786832f
C164 VN.n4 B 0.046475f
C165 VN.n5 B 0.024937f
C166 VN.n6 B 0.046475f
C167 VN.t2 B 1.01576f
C168 VN.n7 B 0.373397f
C169 VN.t0 B 0.786832f
C170 VN.n8 B 0.3818f
C171 VN.n9 B 0.029955f
C172 VN.n10 B 0.268026f
C173 VN.n11 B 0.024937f
C174 VN.n12 B 0.024937f
C175 VN.n13 B 0.049561f
C176 VN.n14 B 0.020159f
C177 VN.n15 B 0.049561f
C178 VN.n16 B 0.024937f
C179 VN.n17 B 0.024937f
C180 VN.n18 B 0.024937f
C181 VN.n19 B 0.029955f
C182 VN.n20 B 0.308129f
C183 VN.n21 B 0.040051f
C184 VN.n22 B 0.046475f
C185 VN.n23 B 0.024937f
C186 VN.n24 B 0.024937f
C187 VN.n25 B 0.024937f
C188 VN.n26 B 0.034318f
C189 VN.n27 B 0.046475f
C190 VN.n28 B 0.042804f
C191 VN.n29 B 0.040247f
C192 VN.n30 B 0.050866f
C193 VN.t6 B 0.786832f
C194 VN.n31 B 0.406132f
C195 VN.n32 B 0.024937f
C196 VN.n33 B 0.038487f
C197 VN.n34 B 0.024937f
C198 VN.t7 B 0.786832f
C199 VN.n35 B 0.046475f
C200 VN.n36 B 0.024937f
C201 VN.n37 B 0.046475f
C202 VN.t3 B 1.01576f
C203 VN.n38 B 0.373397f
C204 VN.t4 B 0.786832f
C205 VN.n39 B 0.3818f
C206 VN.n40 B 0.029955f
C207 VN.n41 B 0.268027f
C208 VN.n42 B 0.024937f
C209 VN.n43 B 0.024937f
C210 VN.n44 B 0.049561f
C211 VN.n45 B 0.020159f
C212 VN.n46 B 0.049561f
C213 VN.n47 B 0.024937f
C214 VN.n48 B 0.024937f
C215 VN.n49 B 0.024937f
C216 VN.n50 B 0.029955f
C217 VN.n51 B 0.308129f
C218 VN.n52 B 0.040051f
C219 VN.n53 B 0.046475f
C220 VN.n54 B 0.024937f
C221 VN.n55 B 0.024937f
C222 VN.n56 B 0.024937f
C223 VN.n57 B 0.034318f
C224 VN.n58 B 0.046475f
C225 VN.n59 B 0.042804f
C226 VN.n60 B 0.040247f
C227 VN.n61 B 1.28429f
.ends

