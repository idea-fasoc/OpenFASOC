* NGSPICE file created from diff_pair_sample_0404.ext - technology: sky130A

.subckt diff_pair_sample_0404 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t1 VN.t0 VTAIL.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=3.0888 pd=16.62 as=3.0888 ps=16.62 w=7.92 l=0.23
X1 B.t15 B.t13 B.t14 B.t3 sky130_fd_pr__nfet_01v8 ad=3.0888 pd=16.62 as=0 ps=0 w=7.92 l=0.23
X2 VDD2.t0 VN.t1 VTAIL.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=3.0888 pd=16.62 as=3.0888 ps=16.62 w=7.92 l=0.23
X3 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=3.0888 pd=16.62 as=0 ps=0 w=7.92 l=0.23
X4 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=3.0888 pd=16.62 as=0 ps=0 w=7.92 l=0.23
X5 VDD1.t1 VP.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=3.0888 pd=16.62 as=3.0888 ps=16.62 w=7.92 l=0.23
X6 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=3.0888 pd=16.62 as=0 ps=0 w=7.92 l=0.23
X7 VDD1.t0 VP.t1 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=3.0888 pd=16.62 as=3.0888 ps=16.62 w=7.92 l=0.23
R0 VN VN.t0 1187.17
R1 VN VN.t1 1151.55
R2 VTAIL.n162 VTAIL.n126 289.615
R3 VTAIL.n36 VTAIL.n0 289.615
R4 VTAIL.n120 VTAIL.n84 289.615
R5 VTAIL.n78 VTAIL.n42 289.615
R6 VTAIL.n138 VTAIL.n137 185
R7 VTAIL.n143 VTAIL.n142 185
R8 VTAIL.n145 VTAIL.n144 185
R9 VTAIL.n134 VTAIL.n133 185
R10 VTAIL.n151 VTAIL.n150 185
R11 VTAIL.n153 VTAIL.n152 185
R12 VTAIL.n130 VTAIL.n129 185
R13 VTAIL.n160 VTAIL.n159 185
R14 VTAIL.n161 VTAIL.n128 185
R15 VTAIL.n163 VTAIL.n162 185
R16 VTAIL.n12 VTAIL.n11 185
R17 VTAIL.n17 VTAIL.n16 185
R18 VTAIL.n19 VTAIL.n18 185
R19 VTAIL.n8 VTAIL.n7 185
R20 VTAIL.n25 VTAIL.n24 185
R21 VTAIL.n27 VTAIL.n26 185
R22 VTAIL.n4 VTAIL.n3 185
R23 VTAIL.n34 VTAIL.n33 185
R24 VTAIL.n35 VTAIL.n2 185
R25 VTAIL.n37 VTAIL.n36 185
R26 VTAIL.n121 VTAIL.n120 185
R27 VTAIL.n119 VTAIL.n86 185
R28 VTAIL.n118 VTAIL.n117 185
R29 VTAIL.n89 VTAIL.n87 185
R30 VTAIL.n112 VTAIL.n111 185
R31 VTAIL.n110 VTAIL.n109 185
R32 VTAIL.n93 VTAIL.n92 185
R33 VTAIL.n104 VTAIL.n103 185
R34 VTAIL.n102 VTAIL.n101 185
R35 VTAIL.n97 VTAIL.n96 185
R36 VTAIL.n79 VTAIL.n78 185
R37 VTAIL.n77 VTAIL.n44 185
R38 VTAIL.n76 VTAIL.n75 185
R39 VTAIL.n47 VTAIL.n45 185
R40 VTAIL.n70 VTAIL.n69 185
R41 VTAIL.n68 VTAIL.n67 185
R42 VTAIL.n51 VTAIL.n50 185
R43 VTAIL.n62 VTAIL.n61 185
R44 VTAIL.n60 VTAIL.n59 185
R45 VTAIL.n55 VTAIL.n54 185
R46 VTAIL.n139 VTAIL.t2 149.524
R47 VTAIL.n13 VTAIL.t0 149.524
R48 VTAIL.n98 VTAIL.t3 149.524
R49 VTAIL.n56 VTAIL.t1 149.524
R50 VTAIL.n143 VTAIL.n137 104.615
R51 VTAIL.n144 VTAIL.n143 104.615
R52 VTAIL.n144 VTAIL.n133 104.615
R53 VTAIL.n151 VTAIL.n133 104.615
R54 VTAIL.n152 VTAIL.n151 104.615
R55 VTAIL.n152 VTAIL.n129 104.615
R56 VTAIL.n160 VTAIL.n129 104.615
R57 VTAIL.n161 VTAIL.n160 104.615
R58 VTAIL.n162 VTAIL.n161 104.615
R59 VTAIL.n17 VTAIL.n11 104.615
R60 VTAIL.n18 VTAIL.n17 104.615
R61 VTAIL.n18 VTAIL.n7 104.615
R62 VTAIL.n25 VTAIL.n7 104.615
R63 VTAIL.n26 VTAIL.n25 104.615
R64 VTAIL.n26 VTAIL.n3 104.615
R65 VTAIL.n34 VTAIL.n3 104.615
R66 VTAIL.n35 VTAIL.n34 104.615
R67 VTAIL.n36 VTAIL.n35 104.615
R68 VTAIL.n120 VTAIL.n119 104.615
R69 VTAIL.n119 VTAIL.n118 104.615
R70 VTAIL.n118 VTAIL.n87 104.615
R71 VTAIL.n111 VTAIL.n87 104.615
R72 VTAIL.n111 VTAIL.n110 104.615
R73 VTAIL.n110 VTAIL.n92 104.615
R74 VTAIL.n103 VTAIL.n92 104.615
R75 VTAIL.n103 VTAIL.n102 104.615
R76 VTAIL.n102 VTAIL.n96 104.615
R77 VTAIL.n78 VTAIL.n77 104.615
R78 VTAIL.n77 VTAIL.n76 104.615
R79 VTAIL.n76 VTAIL.n45 104.615
R80 VTAIL.n69 VTAIL.n45 104.615
R81 VTAIL.n69 VTAIL.n68 104.615
R82 VTAIL.n68 VTAIL.n50 104.615
R83 VTAIL.n61 VTAIL.n50 104.615
R84 VTAIL.n61 VTAIL.n60 104.615
R85 VTAIL.n60 VTAIL.n54 104.615
R86 VTAIL.t2 VTAIL.n137 52.3082
R87 VTAIL.t0 VTAIL.n11 52.3082
R88 VTAIL.t3 VTAIL.n96 52.3082
R89 VTAIL.t1 VTAIL.n54 52.3082
R90 VTAIL.n167 VTAIL.n166 34.5126
R91 VTAIL.n41 VTAIL.n40 34.5126
R92 VTAIL.n125 VTAIL.n124 34.5126
R93 VTAIL.n83 VTAIL.n82 34.5126
R94 VTAIL.n83 VTAIL.n41 20.1772
R95 VTAIL.n167 VTAIL.n125 19.6945
R96 VTAIL.n163 VTAIL.n128 13.1884
R97 VTAIL.n37 VTAIL.n2 13.1884
R98 VTAIL.n121 VTAIL.n86 13.1884
R99 VTAIL.n79 VTAIL.n44 13.1884
R100 VTAIL.n159 VTAIL.n158 12.8005
R101 VTAIL.n164 VTAIL.n126 12.8005
R102 VTAIL.n33 VTAIL.n32 12.8005
R103 VTAIL.n38 VTAIL.n0 12.8005
R104 VTAIL.n122 VTAIL.n84 12.8005
R105 VTAIL.n117 VTAIL.n88 12.8005
R106 VTAIL.n80 VTAIL.n42 12.8005
R107 VTAIL.n75 VTAIL.n46 12.8005
R108 VTAIL.n157 VTAIL.n130 12.0247
R109 VTAIL.n31 VTAIL.n4 12.0247
R110 VTAIL.n116 VTAIL.n89 12.0247
R111 VTAIL.n74 VTAIL.n47 12.0247
R112 VTAIL.n154 VTAIL.n153 11.249
R113 VTAIL.n28 VTAIL.n27 11.249
R114 VTAIL.n113 VTAIL.n112 11.249
R115 VTAIL.n71 VTAIL.n70 11.249
R116 VTAIL.n150 VTAIL.n132 10.4732
R117 VTAIL.n24 VTAIL.n6 10.4732
R118 VTAIL.n109 VTAIL.n91 10.4732
R119 VTAIL.n67 VTAIL.n49 10.4732
R120 VTAIL.n139 VTAIL.n138 10.2747
R121 VTAIL.n13 VTAIL.n12 10.2747
R122 VTAIL.n98 VTAIL.n97 10.2747
R123 VTAIL.n56 VTAIL.n55 10.2747
R124 VTAIL.n149 VTAIL.n134 9.69747
R125 VTAIL.n23 VTAIL.n8 9.69747
R126 VTAIL.n108 VTAIL.n93 9.69747
R127 VTAIL.n66 VTAIL.n51 9.69747
R128 VTAIL.n166 VTAIL.n165 9.45567
R129 VTAIL.n40 VTAIL.n39 9.45567
R130 VTAIL.n124 VTAIL.n123 9.45567
R131 VTAIL.n82 VTAIL.n81 9.45567
R132 VTAIL.n165 VTAIL.n164 9.3005
R133 VTAIL.n141 VTAIL.n140 9.3005
R134 VTAIL.n136 VTAIL.n135 9.3005
R135 VTAIL.n147 VTAIL.n146 9.3005
R136 VTAIL.n149 VTAIL.n148 9.3005
R137 VTAIL.n132 VTAIL.n131 9.3005
R138 VTAIL.n155 VTAIL.n154 9.3005
R139 VTAIL.n157 VTAIL.n156 9.3005
R140 VTAIL.n158 VTAIL.n127 9.3005
R141 VTAIL.n39 VTAIL.n38 9.3005
R142 VTAIL.n15 VTAIL.n14 9.3005
R143 VTAIL.n10 VTAIL.n9 9.3005
R144 VTAIL.n21 VTAIL.n20 9.3005
R145 VTAIL.n23 VTAIL.n22 9.3005
R146 VTAIL.n6 VTAIL.n5 9.3005
R147 VTAIL.n29 VTAIL.n28 9.3005
R148 VTAIL.n31 VTAIL.n30 9.3005
R149 VTAIL.n32 VTAIL.n1 9.3005
R150 VTAIL.n100 VTAIL.n99 9.3005
R151 VTAIL.n95 VTAIL.n94 9.3005
R152 VTAIL.n106 VTAIL.n105 9.3005
R153 VTAIL.n108 VTAIL.n107 9.3005
R154 VTAIL.n91 VTAIL.n90 9.3005
R155 VTAIL.n114 VTAIL.n113 9.3005
R156 VTAIL.n116 VTAIL.n115 9.3005
R157 VTAIL.n88 VTAIL.n85 9.3005
R158 VTAIL.n123 VTAIL.n122 9.3005
R159 VTAIL.n58 VTAIL.n57 9.3005
R160 VTAIL.n53 VTAIL.n52 9.3005
R161 VTAIL.n64 VTAIL.n63 9.3005
R162 VTAIL.n66 VTAIL.n65 9.3005
R163 VTAIL.n49 VTAIL.n48 9.3005
R164 VTAIL.n72 VTAIL.n71 9.3005
R165 VTAIL.n74 VTAIL.n73 9.3005
R166 VTAIL.n46 VTAIL.n43 9.3005
R167 VTAIL.n81 VTAIL.n80 9.3005
R168 VTAIL.n146 VTAIL.n145 8.92171
R169 VTAIL.n20 VTAIL.n19 8.92171
R170 VTAIL.n105 VTAIL.n104 8.92171
R171 VTAIL.n63 VTAIL.n62 8.92171
R172 VTAIL.n142 VTAIL.n136 8.14595
R173 VTAIL.n16 VTAIL.n10 8.14595
R174 VTAIL.n101 VTAIL.n95 8.14595
R175 VTAIL.n59 VTAIL.n53 8.14595
R176 VTAIL.n141 VTAIL.n138 7.3702
R177 VTAIL.n15 VTAIL.n12 7.3702
R178 VTAIL.n100 VTAIL.n97 7.3702
R179 VTAIL.n58 VTAIL.n55 7.3702
R180 VTAIL.n142 VTAIL.n141 5.81868
R181 VTAIL.n16 VTAIL.n15 5.81868
R182 VTAIL.n101 VTAIL.n100 5.81868
R183 VTAIL.n59 VTAIL.n58 5.81868
R184 VTAIL.n145 VTAIL.n136 5.04292
R185 VTAIL.n19 VTAIL.n10 5.04292
R186 VTAIL.n104 VTAIL.n95 5.04292
R187 VTAIL.n62 VTAIL.n53 5.04292
R188 VTAIL.n146 VTAIL.n134 4.26717
R189 VTAIL.n20 VTAIL.n8 4.26717
R190 VTAIL.n105 VTAIL.n93 4.26717
R191 VTAIL.n63 VTAIL.n51 4.26717
R192 VTAIL.n150 VTAIL.n149 3.49141
R193 VTAIL.n24 VTAIL.n23 3.49141
R194 VTAIL.n109 VTAIL.n108 3.49141
R195 VTAIL.n67 VTAIL.n66 3.49141
R196 VTAIL.n140 VTAIL.n139 2.84304
R197 VTAIL.n14 VTAIL.n13 2.84304
R198 VTAIL.n99 VTAIL.n98 2.84304
R199 VTAIL.n57 VTAIL.n56 2.84304
R200 VTAIL.n153 VTAIL.n132 2.71565
R201 VTAIL.n27 VTAIL.n6 2.71565
R202 VTAIL.n112 VTAIL.n91 2.71565
R203 VTAIL.n70 VTAIL.n49 2.71565
R204 VTAIL.n154 VTAIL.n130 1.93989
R205 VTAIL.n28 VTAIL.n4 1.93989
R206 VTAIL.n113 VTAIL.n89 1.93989
R207 VTAIL.n71 VTAIL.n47 1.93989
R208 VTAIL.n159 VTAIL.n157 1.16414
R209 VTAIL.n166 VTAIL.n126 1.16414
R210 VTAIL.n33 VTAIL.n31 1.16414
R211 VTAIL.n40 VTAIL.n0 1.16414
R212 VTAIL.n124 VTAIL.n84 1.16414
R213 VTAIL.n117 VTAIL.n116 1.16414
R214 VTAIL.n82 VTAIL.n42 1.16414
R215 VTAIL.n75 VTAIL.n74 1.16414
R216 VTAIL.n125 VTAIL.n83 0.711707
R217 VTAIL VTAIL.n41 0.649207
R218 VTAIL.n158 VTAIL.n128 0.388379
R219 VTAIL.n164 VTAIL.n163 0.388379
R220 VTAIL.n32 VTAIL.n2 0.388379
R221 VTAIL.n38 VTAIL.n37 0.388379
R222 VTAIL.n122 VTAIL.n121 0.388379
R223 VTAIL.n88 VTAIL.n86 0.388379
R224 VTAIL.n80 VTAIL.n79 0.388379
R225 VTAIL.n46 VTAIL.n44 0.388379
R226 VTAIL.n140 VTAIL.n135 0.155672
R227 VTAIL.n147 VTAIL.n135 0.155672
R228 VTAIL.n148 VTAIL.n147 0.155672
R229 VTAIL.n148 VTAIL.n131 0.155672
R230 VTAIL.n155 VTAIL.n131 0.155672
R231 VTAIL.n156 VTAIL.n155 0.155672
R232 VTAIL.n156 VTAIL.n127 0.155672
R233 VTAIL.n165 VTAIL.n127 0.155672
R234 VTAIL.n14 VTAIL.n9 0.155672
R235 VTAIL.n21 VTAIL.n9 0.155672
R236 VTAIL.n22 VTAIL.n21 0.155672
R237 VTAIL.n22 VTAIL.n5 0.155672
R238 VTAIL.n29 VTAIL.n5 0.155672
R239 VTAIL.n30 VTAIL.n29 0.155672
R240 VTAIL.n30 VTAIL.n1 0.155672
R241 VTAIL.n39 VTAIL.n1 0.155672
R242 VTAIL.n123 VTAIL.n85 0.155672
R243 VTAIL.n115 VTAIL.n85 0.155672
R244 VTAIL.n115 VTAIL.n114 0.155672
R245 VTAIL.n114 VTAIL.n90 0.155672
R246 VTAIL.n107 VTAIL.n90 0.155672
R247 VTAIL.n107 VTAIL.n106 0.155672
R248 VTAIL.n106 VTAIL.n94 0.155672
R249 VTAIL.n99 VTAIL.n94 0.155672
R250 VTAIL.n81 VTAIL.n43 0.155672
R251 VTAIL.n73 VTAIL.n43 0.155672
R252 VTAIL.n73 VTAIL.n72 0.155672
R253 VTAIL.n72 VTAIL.n48 0.155672
R254 VTAIL.n65 VTAIL.n48 0.155672
R255 VTAIL.n65 VTAIL.n64 0.155672
R256 VTAIL.n64 VTAIL.n52 0.155672
R257 VTAIL.n57 VTAIL.n52 0.155672
R258 VTAIL VTAIL.n167 0.063
R259 VDD2.n77 VDD2.n41 289.615
R260 VDD2.n36 VDD2.n0 289.615
R261 VDD2.n78 VDD2.n77 185
R262 VDD2.n76 VDD2.n43 185
R263 VDD2.n75 VDD2.n74 185
R264 VDD2.n46 VDD2.n44 185
R265 VDD2.n69 VDD2.n68 185
R266 VDD2.n67 VDD2.n66 185
R267 VDD2.n50 VDD2.n49 185
R268 VDD2.n61 VDD2.n60 185
R269 VDD2.n59 VDD2.n58 185
R270 VDD2.n54 VDD2.n53 185
R271 VDD2.n12 VDD2.n11 185
R272 VDD2.n17 VDD2.n16 185
R273 VDD2.n19 VDD2.n18 185
R274 VDD2.n8 VDD2.n7 185
R275 VDD2.n25 VDD2.n24 185
R276 VDD2.n27 VDD2.n26 185
R277 VDD2.n4 VDD2.n3 185
R278 VDD2.n34 VDD2.n33 185
R279 VDD2.n35 VDD2.n2 185
R280 VDD2.n37 VDD2.n36 185
R281 VDD2.n55 VDD2.t1 149.524
R282 VDD2.n13 VDD2.t0 149.524
R283 VDD2.n77 VDD2.n76 104.615
R284 VDD2.n76 VDD2.n75 104.615
R285 VDD2.n75 VDD2.n44 104.615
R286 VDD2.n68 VDD2.n44 104.615
R287 VDD2.n68 VDD2.n67 104.615
R288 VDD2.n67 VDD2.n49 104.615
R289 VDD2.n60 VDD2.n49 104.615
R290 VDD2.n60 VDD2.n59 104.615
R291 VDD2.n59 VDD2.n53 104.615
R292 VDD2.n17 VDD2.n11 104.615
R293 VDD2.n18 VDD2.n17 104.615
R294 VDD2.n18 VDD2.n7 104.615
R295 VDD2.n25 VDD2.n7 104.615
R296 VDD2.n26 VDD2.n25 104.615
R297 VDD2.n26 VDD2.n3 104.615
R298 VDD2.n34 VDD2.n3 104.615
R299 VDD2.n35 VDD2.n34 104.615
R300 VDD2.n36 VDD2.n35 104.615
R301 VDD2.n82 VDD2.n40 82.6612
R302 VDD2.t1 VDD2.n53 52.3082
R303 VDD2.t0 VDD2.n11 52.3082
R304 VDD2.n82 VDD2.n81 51.1914
R305 VDD2.n78 VDD2.n43 13.1884
R306 VDD2.n37 VDD2.n2 13.1884
R307 VDD2.n79 VDD2.n41 12.8005
R308 VDD2.n74 VDD2.n45 12.8005
R309 VDD2.n33 VDD2.n32 12.8005
R310 VDD2.n38 VDD2.n0 12.8005
R311 VDD2.n73 VDD2.n46 12.0247
R312 VDD2.n31 VDD2.n4 12.0247
R313 VDD2.n70 VDD2.n69 11.249
R314 VDD2.n28 VDD2.n27 11.249
R315 VDD2.n66 VDD2.n48 10.4732
R316 VDD2.n24 VDD2.n6 10.4732
R317 VDD2.n55 VDD2.n54 10.2747
R318 VDD2.n13 VDD2.n12 10.2747
R319 VDD2.n65 VDD2.n50 9.69747
R320 VDD2.n23 VDD2.n8 9.69747
R321 VDD2.n81 VDD2.n80 9.45567
R322 VDD2.n40 VDD2.n39 9.45567
R323 VDD2.n57 VDD2.n56 9.3005
R324 VDD2.n52 VDD2.n51 9.3005
R325 VDD2.n63 VDD2.n62 9.3005
R326 VDD2.n65 VDD2.n64 9.3005
R327 VDD2.n48 VDD2.n47 9.3005
R328 VDD2.n71 VDD2.n70 9.3005
R329 VDD2.n73 VDD2.n72 9.3005
R330 VDD2.n45 VDD2.n42 9.3005
R331 VDD2.n80 VDD2.n79 9.3005
R332 VDD2.n39 VDD2.n38 9.3005
R333 VDD2.n15 VDD2.n14 9.3005
R334 VDD2.n10 VDD2.n9 9.3005
R335 VDD2.n21 VDD2.n20 9.3005
R336 VDD2.n23 VDD2.n22 9.3005
R337 VDD2.n6 VDD2.n5 9.3005
R338 VDD2.n29 VDD2.n28 9.3005
R339 VDD2.n31 VDD2.n30 9.3005
R340 VDD2.n32 VDD2.n1 9.3005
R341 VDD2.n62 VDD2.n61 8.92171
R342 VDD2.n20 VDD2.n19 8.92171
R343 VDD2.n58 VDD2.n52 8.14595
R344 VDD2.n16 VDD2.n10 8.14595
R345 VDD2.n57 VDD2.n54 7.3702
R346 VDD2.n15 VDD2.n12 7.3702
R347 VDD2.n58 VDD2.n57 5.81868
R348 VDD2.n16 VDD2.n15 5.81868
R349 VDD2.n61 VDD2.n52 5.04292
R350 VDD2.n19 VDD2.n10 5.04292
R351 VDD2.n62 VDD2.n50 4.26717
R352 VDD2.n20 VDD2.n8 4.26717
R353 VDD2.n66 VDD2.n65 3.49141
R354 VDD2.n24 VDD2.n23 3.49141
R355 VDD2.n56 VDD2.n55 2.84304
R356 VDD2.n14 VDD2.n13 2.84304
R357 VDD2.n69 VDD2.n48 2.71565
R358 VDD2.n27 VDD2.n6 2.71565
R359 VDD2.n70 VDD2.n46 1.93989
R360 VDD2.n28 VDD2.n4 1.93989
R361 VDD2.n81 VDD2.n41 1.16414
R362 VDD2.n74 VDD2.n73 1.16414
R363 VDD2.n33 VDD2.n31 1.16414
R364 VDD2.n40 VDD2.n0 1.16414
R365 VDD2.n79 VDD2.n78 0.388379
R366 VDD2.n45 VDD2.n43 0.388379
R367 VDD2.n32 VDD2.n2 0.388379
R368 VDD2.n38 VDD2.n37 0.388379
R369 VDD2 VDD2.n82 0.179379
R370 VDD2.n80 VDD2.n42 0.155672
R371 VDD2.n72 VDD2.n42 0.155672
R372 VDD2.n72 VDD2.n71 0.155672
R373 VDD2.n71 VDD2.n47 0.155672
R374 VDD2.n64 VDD2.n47 0.155672
R375 VDD2.n64 VDD2.n63 0.155672
R376 VDD2.n63 VDD2.n51 0.155672
R377 VDD2.n56 VDD2.n51 0.155672
R378 VDD2.n14 VDD2.n9 0.155672
R379 VDD2.n21 VDD2.n9 0.155672
R380 VDD2.n22 VDD2.n21 0.155672
R381 VDD2.n22 VDD2.n5 0.155672
R382 VDD2.n29 VDD2.n5 0.155672
R383 VDD2.n30 VDD2.n29 0.155672
R384 VDD2.n30 VDD2.n1 0.155672
R385 VDD2.n39 VDD2.n1 0.155672
R386 B.n64 B.t10 1058.37
R387 B.n62 B.t6 1058.37
R388 B.n260 B.t2 1058.37
R389 B.n258 B.t13 1058.37
R390 B.n450 B.n449 585
R391 B.n451 B.n450 585
R392 B.n202 B.n61 585
R393 B.n201 B.n200 585
R394 B.n199 B.n198 585
R395 B.n197 B.n196 585
R396 B.n195 B.n194 585
R397 B.n193 B.n192 585
R398 B.n191 B.n190 585
R399 B.n189 B.n188 585
R400 B.n187 B.n186 585
R401 B.n185 B.n184 585
R402 B.n183 B.n182 585
R403 B.n181 B.n180 585
R404 B.n179 B.n178 585
R405 B.n177 B.n176 585
R406 B.n175 B.n174 585
R407 B.n173 B.n172 585
R408 B.n171 B.n170 585
R409 B.n169 B.n168 585
R410 B.n167 B.n166 585
R411 B.n165 B.n164 585
R412 B.n163 B.n162 585
R413 B.n161 B.n160 585
R414 B.n159 B.n158 585
R415 B.n157 B.n156 585
R416 B.n155 B.n154 585
R417 B.n153 B.n152 585
R418 B.n151 B.n150 585
R419 B.n149 B.n148 585
R420 B.n147 B.n146 585
R421 B.n144 B.n143 585
R422 B.n142 B.n141 585
R423 B.n140 B.n139 585
R424 B.n138 B.n137 585
R425 B.n136 B.n135 585
R426 B.n134 B.n133 585
R427 B.n132 B.n131 585
R428 B.n130 B.n129 585
R429 B.n128 B.n127 585
R430 B.n126 B.n125 585
R431 B.n124 B.n123 585
R432 B.n122 B.n121 585
R433 B.n120 B.n119 585
R434 B.n118 B.n117 585
R435 B.n116 B.n115 585
R436 B.n114 B.n113 585
R437 B.n112 B.n111 585
R438 B.n110 B.n109 585
R439 B.n108 B.n107 585
R440 B.n106 B.n105 585
R441 B.n104 B.n103 585
R442 B.n102 B.n101 585
R443 B.n100 B.n99 585
R444 B.n98 B.n97 585
R445 B.n96 B.n95 585
R446 B.n94 B.n93 585
R447 B.n92 B.n91 585
R448 B.n90 B.n89 585
R449 B.n88 B.n87 585
R450 B.n86 B.n85 585
R451 B.n84 B.n83 585
R452 B.n82 B.n81 585
R453 B.n80 B.n79 585
R454 B.n78 B.n77 585
R455 B.n76 B.n75 585
R456 B.n74 B.n73 585
R457 B.n72 B.n71 585
R458 B.n70 B.n69 585
R459 B.n68 B.n67 585
R460 B.n448 B.n26 585
R461 B.n452 B.n26 585
R462 B.n447 B.n25 585
R463 B.n453 B.n25 585
R464 B.n446 B.n445 585
R465 B.n445 B.n21 585
R466 B.n444 B.n20 585
R467 B.n459 B.n20 585
R468 B.n443 B.n19 585
R469 B.n460 B.n19 585
R470 B.n442 B.n18 585
R471 B.n461 B.n18 585
R472 B.n441 B.n440 585
R473 B.n440 B.n13 585
R474 B.n439 B.n12 585
R475 B.n467 B.n12 585
R476 B.n438 B.n11 585
R477 B.n468 B.n11 585
R478 B.n437 B.n10 585
R479 B.n469 B.n10 585
R480 B.n436 B.n7 585
R481 B.n472 B.n7 585
R482 B.n435 B.n6 585
R483 B.n473 B.n6 585
R484 B.n434 B.n5 585
R485 B.n474 B.n5 585
R486 B.n433 B.n432 585
R487 B.n432 B.n4 585
R488 B.n431 B.n203 585
R489 B.n431 B.n430 585
R490 B.n421 B.n204 585
R491 B.n205 B.n204 585
R492 B.n423 B.n422 585
R493 B.n424 B.n423 585
R494 B.n420 B.n210 585
R495 B.n210 B.n209 585
R496 B.n419 B.n418 585
R497 B.n418 B.n417 585
R498 B.n212 B.n211 585
R499 B.n410 B.n212 585
R500 B.n409 B.n408 585
R501 B.n411 B.n409 585
R502 B.n407 B.n217 585
R503 B.n217 B.n216 585
R504 B.n406 B.n405 585
R505 B.n405 B.n404 585
R506 B.n219 B.n218 585
R507 B.n220 B.n219 585
R508 B.n400 B.n399 585
R509 B.n223 B.n222 585
R510 B.n396 B.n395 585
R511 B.n397 B.n396 585
R512 B.n394 B.n257 585
R513 B.n393 B.n392 585
R514 B.n391 B.n390 585
R515 B.n389 B.n388 585
R516 B.n387 B.n386 585
R517 B.n385 B.n384 585
R518 B.n383 B.n382 585
R519 B.n381 B.n380 585
R520 B.n379 B.n378 585
R521 B.n377 B.n376 585
R522 B.n375 B.n374 585
R523 B.n373 B.n372 585
R524 B.n371 B.n370 585
R525 B.n369 B.n368 585
R526 B.n367 B.n366 585
R527 B.n365 B.n364 585
R528 B.n363 B.n362 585
R529 B.n361 B.n360 585
R530 B.n359 B.n358 585
R531 B.n357 B.n356 585
R532 B.n355 B.n354 585
R533 B.n353 B.n352 585
R534 B.n351 B.n350 585
R535 B.n349 B.n348 585
R536 B.n347 B.n346 585
R537 B.n345 B.n344 585
R538 B.n343 B.n342 585
R539 B.n340 B.n339 585
R540 B.n338 B.n337 585
R541 B.n336 B.n335 585
R542 B.n334 B.n333 585
R543 B.n332 B.n331 585
R544 B.n330 B.n329 585
R545 B.n328 B.n327 585
R546 B.n326 B.n325 585
R547 B.n324 B.n323 585
R548 B.n322 B.n321 585
R549 B.n320 B.n319 585
R550 B.n318 B.n317 585
R551 B.n316 B.n315 585
R552 B.n314 B.n313 585
R553 B.n312 B.n311 585
R554 B.n310 B.n309 585
R555 B.n308 B.n307 585
R556 B.n306 B.n305 585
R557 B.n304 B.n303 585
R558 B.n302 B.n301 585
R559 B.n300 B.n299 585
R560 B.n298 B.n297 585
R561 B.n296 B.n295 585
R562 B.n294 B.n293 585
R563 B.n292 B.n291 585
R564 B.n290 B.n289 585
R565 B.n288 B.n287 585
R566 B.n286 B.n285 585
R567 B.n284 B.n283 585
R568 B.n282 B.n281 585
R569 B.n280 B.n279 585
R570 B.n278 B.n277 585
R571 B.n276 B.n275 585
R572 B.n274 B.n273 585
R573 B.n272 B.n271 585
R574 B.n270 B.n269 585
R575 B.n268 B.n267 585
R576 B.n266 B.n265 585
R577 B.n264 B.n263 585
R578 B.n401 B.n221 585
R579 B.n221 B.n220 585
R580 B.n403 B.n402 585
R581 B.n404 B.n403 585
R582 B.n215 B.n214 585
R583 B.n216 B.n215 585
R584 B.n413 B.n412 585
R585 B.n412 B.n411 585
R586 B.n414 B.n213 585
R587 B.n410 B.n213 585
R588 B.n416 B.n415 585
R589 B.n417 B.n416 585
R590 B.n208 B.n207 585
R591 B.n209 B.n208 585
R592 B.n426 B.n425 585
R593 B.n425 B.n424 585
R594 B.n427 B.n206 585
R595 B.n206 B.n205 585
R596 B.n429 B.n428 585
R597 B.n430 B.n429 585
R598 B.n3 B.n0 585
R599 B.n4 B.n3 585
R600 B.n471 B.n1 585
R601 B.n472 B.n471 585
R602 B.n470 B.n9 585
R603 B.n470 B.n469 585
R604 B.n15 B.n8 585
R605 B.n468 B.n8 585
R606 B.n466 B.n465 585
R607 B.n467 B.n466 585
R608 B.n464 B.n14 585
R609 B.n14 B.n13 585
R610 B.n463 B.n462 585
R611 B.n462 B.n461 585
R612 B.n17 B.n16 585
R613 B.n460 B.n17 585
R614 B.n458 B.n457 585
R615 B.n459 B.n458 585
R616 B.n456 B.n22 585
R617 B.n22 B.n21 585
R618 B.n455 B.n454 585
R619 B.n454 B.n453 585
R620 B.n24 B.n23 585
R621 B.n452 B.n24 585
R622 B.n475 B.n474 585
R623 B.n473 B.n2 585
R624 B.n67 B.n24 478.086
R625 B.n450 B.n26 478.086
R626 B.n263 B.n219 478.086
R627 B.n399 B.n221 478.086
R628 B.n451 B.n60 256.663
R629 B.n451 B.n59 256.663
R630 B.n451 B.n58 256.663
R631 B.n451 B.n57 256.663
R632 B.n451 B.n56 256.663
R633 B.n451 B.n55 256.663
R634 B.n451 B.n54 256.663
R635 B.n451 B.n53 256.663
R636 B.n451 B.n52 256.663
R637 B.n451 B.n51 256.663
R638 B.n451 B.n50 256.663
R639 B.n451 B.n49 256.663
R640 B.n451 B.n48 256.663
R641 B.n451 B.n47 256.663
R642 B.n451 B.n46 256.663
R643 B.n451 B.n45 256.663
R644 B.n451 B.n44 256.663
R645 B.n451 B.n43 256.663
R646 B.n451 B.n42 256.663
R647 B.n451 B.n41 256.663
R648 B.n451 B.n40 256.663
R649 B.n451 B.n39 256.663
R650 B.n451 B.n38 256.663
R651 B.n451 B.n37 256.663
R652 B.n451 B.n36 256.663
R653 B.n451 B.n35 256.663
R654 B.n451 B.n34 256.663
R655 B.n451 B.n33 256.663
R656 B.n451 B.n32 256.663
R657 B.n451 B.n31 256.663
R658 B.n451 B.n30 256.663
R659 B.n451 B.n29 256.663
R660 B.n451 B.n28 256.663
R661 B.n451 B.n27 256.663
R662 B.n398 B.n397 256.663
R663 B.n397 B.n224 256.663
R664 B.n397 B.n225 256.663
R665 B.n397 B.n226 256.663
R666 B.n397 B.n227 256.663
R667 B.n397 B.n228 256.663
R668 B.n397 B.n229 256.663
R669 B.n397 B.n230 256.663
R670 B.n397 B.n231 256.663
R671 B.n397 B.n232 256.663
R672 B.n397 B.n233 256.663
R673 B.n397 B.n234 256.663
R674 B.n397 B.n235 256.663
R675 B.n397 B.n236 256.663
R676 B.n397 B.n237 256.663
R677 B.n397 B.n238 256.663
R678 B.n397 B.n239 256.663
R679 B.n397 B.n240 256.663
R680 B.n397 B.n241 256.663
R681 B.n397 B.n242 256.663
R682 B.n397 B.n243 256.663
R683 B.n397 B.n244 256.663
R684 B.n397 B.n245 256.663
R685 B.n397 B.n246 256.663
R686 B.n397 B.n247 256.663
R687 B.n397 B.n248 256.663
R688 B.n397 B.n249 256.663
R689 B.n397 B.n250 256.663
R690 B.n397 B.n251 256.663
R691 B.n397 B.n252 256.663
R692 B.n397 B.n253 256.663
R693 B.n397 B.n254 256.663
R694 B.n397 B.n255 256.663
R695 B.n397 B.n256 256.663
R696 B.n477 B.n476 256.663
R697 B.n62 B.t8 222.601
R698 B.n260 B.t5 222.601
R699 B.n64 B.t11 222.601
R700 B.n258 B.t15 222.601
R701 B.n63 B.t9 211.739
R702 B.n261 B.t4 211.739
R703 B.n65 B.t12 211.739
R704 B.n259 B.t14 211.739
R705 B.n71 B.n70 163.367
R706 B.n75 B.n74 163.367
R707 B.n79 B.n78 163.367
R708 B.n83 B.n82 163.367
R709 B.n87 B.n86 163.367
R710 B.n91 B.n90 163.367
R711 B.n95 B.n94 163.367
R712 B.n99 B.n98 163.367
R713 B.n103 B.n102 163.367
R714 B.n107 B.n106 163.367
R715 B.n111 B.n110 163.367
R716 B.n115 B.n114 163.367
R717 B.n119 B.n118 163.367
R718 B.n123 B.n122 163.367
R719 B.n127 B.n126 163.367
R720 B.n131 B.n130 163.367
R721 B.n135 B.n134 163.367
R722 B.n139 B.n138 163.367
R723 B.n143 B.n142 163.367
R724 B.n148 B.n147 163.367
R725 B.n152 B.n151 163.367
R726 B.n156 B.n155 163.367
R727 B.n160 B.n159 163.367
R728 B.n164 B.n163 163.367
R729 B.n168 B.n167 163.367
R730 B.n172 B.n171 163.367
R731 B.n176 B.n175 163.367
R732 B.n180 B.n179 163.367
R733 B.n184 B.n183 163.367
R734 B.n188 B.n187 163.367
R735 B.n192 B.n191 163.367
R736 B.n196 B.n195 163.367
R737 B.n200 B.n199 163.367
R738 B.n450 B.n61 163.367
R739 B.n405 B.n219 163.367
R740 B.n405 B.n217 163.367
R741 B.n409 B.n217 163.367
R742 B.n409 B.n212 163.367
R743 B.n418 B.n212 163.367
R744 B.n418 B.n210 163.367
R745 B.n423 B.n210 163.367
R746 B.n423 B.n204 163.367
R747 B.n431 B.n204 163.367
R748 B.n432 B.n431 163.367
R749 B.n432 B.n5 163.367
R750 B.n6 B.n5 163.367
R751 B.n7 B.n6 163.367
R752 B.n10 B.n7 163.367
R753 B.n11 B.n10 163.367
R754 B.n12 B.n11 163.367
R755 B.n440 B.n12 163.367
R756 B.n440 B.n18 163.367
R757 B.n19 B.n18 163.367
R758 B.n20 B.n19 163.367
R759 B.n445 B.n20 163.367
R760 B.n445 B.n25 163.367
R761 B.n26 B.n25 163.367
R762 B.n396 B.n223 163.367
R763 B.n396 B.n257 163.367
R764 B.n392 B.n391 163.367
R765 B.n388 B.n387 163.367
R766 B.n384 B.n383 163.367
R767 B.n380 B.n379 163.367
R768 B.n376 B.n375 163.367
R769 B.n372 B.n371 163.367
R770 B.n368 B.n367 163.367
R771 B.n364 B.n363 163.367
R772 B.n360 B.n359 163.367
R773 B.n356 B.n355 163.367
R774 B.n352 B.n351 163.367
R775 B.n348 B.n347 163.367
R776 B.n344 B.n343 163.367
R777 B.n339 B.n338 163.367
R778 B.n335 B.n334 163.367
R779 B.n331 B.n330 163.367
R780 B.n327 B.n326 163.367
R781 B.n323 B.n322 163.367
R782 B.n319 B.n318 163.367
R783 B.n315 B.n314 163.367
R784 B.n311 B.n310 163.367
R785 B.n307 B.n306 163.367
R786 B.n303 B.n302 163.367
R787 B.n299 B.n298 163.367
R788 B.n295 B.n294 163.367
R789 B.n291 B.n290 163.367
R790 B.n287 B.n286 163.367
R791 B.n283 B.n282 163.367
R792 B.n279 B.n278 163.367
R793 B.n275 B.n274 163.367
R794 B.n271 B.n270 163.367
R795 B.n267 B.n266 163.367
R796 B.n403 B.n221 163.367
R797 B.n403 B.n215 163.367
R798 B.n412 B.n215 163.367
R799 B.n412 B.n213 163.367
R800 B.n416 B.n213 163.367
R801 B.n416 B.n208 163.367
R802 B.n425 B.n208 163.367
R803 B.n425 B.n206 163.367
R804 B.n429 B.n206 163.367
R805 B.n429 B.n3 163.367
R806 B.n475 B.n3 163.367
R807 B.n471 B.n2 163.367
R808 B.n471 B.n470 163.367
R809 B.n470 B.n8 163.367
R810 B.n466 B.n8 163.367
R811 B.n466 B.n14 163.367
R812 B.n462 B.n14 163.367
R813 B.n462 B.n17 163.367
R814 B.n458 B.n17 163.367
R815 B.n458 B.n22 163.367
R816 B.n454 B.n22 163.367
R817 B.n454 B.n24 163.367
R818 B.n397 B.n220 97.3898
R819 B.n452 B.n451 97.3898
R820 B.n67 B.n27 71.676
R821 B.n71 B.n28 71.676
R822 B.n75 B.n29 71.676
R823 B.n79 B.n30 71.676
R824 B.n83 B.n31 71.676
R825 B.n87 B.n32 71.676
R826 B.n91 B.n33 71.676
R827 B.n95 B.n34 71.676
R828 B.n99 B.n35 71.676
R829 B.n103 B.n36 71.676
R830 B.n107 B.n37 71.676
R831 B.n111 B.n38 71.676
R832 B.n115 B.n39 71.676
R833 B.n119 B.n40 71.676
R834 B.n123 B.n41 71.676
R835 B.n127 B.n42 71.676
R836 B.n131 B.n43 71.676
R837 B.n135 B.n44 71.676
R838 B.n139 B.n45 71.676
R839 B.n143 B.n46 71.676
R840 B.n148 B.n47 71.676
R841 B.n152 B.n48 71.676
R842 B.n156 B.n49 71.676
R843 B.n160 B.n50 71.676
R844 B.n164 B.n51 71.676
R845 B.n168 B.n52 71.676
R846 B.n172 B.n53 71.676
R847 B.n176 B.n54 71.676
R848 B.n180 B.n55 71.676
R849 B.n184 B.n56 71.676
R850 B.n188 B.n57 71.676
R851 B.n192 B.n58 71.676
R852 B.n196 B.n59 71.676
R853 B.n200 B.n60 71.676
R854 B.n61 B.n60 71.676
R855 B.n199 B.n59 71.676
R856 B.n195 B.n58 71.676
R857 B.n191 B.n57 71.676
R858 B.n187 B.n56 71.676
R859 B.n183 B.n55 71.676
R860 B.n179 B.n54 71.676
R861 B.n175 B.n53 71.676
R862 B.n171 B.n52 71.676
R863 B.n167 B.n51 71.676
R864 B.n163 B.n50 71.676
R865 B.n159 B.n49 71.676
R866 B.n155 B.n48 71.676
R867 B.n151 B.n47 71.676
R868 B.n147 B.n46 71.676
R869 B.n142 B.n45 71.676
R870 B.n138 B.n44 71.676
R871 B.n134 B.n43 71.676
R872 B.n130 B.n42 71.676
R873 B.n126 B.n41 71.676
R874 B.n122 B.n40 71.676
R875 B.n118 B.n39 71.676
R876 B.n114 B.n38 71.676
R877 B.n110 B.n37 71.676
R878 B.n106 B.n36 71.676
R879 B.n102 B.n35 71.676
R880 B.n98 B.n34 71.676
R881 B.n94 B.n33 71.676
R882 B.n90 B.n32 71.676
R883 B.n86 B.n31 71.676
R884 B.n82 B.n30 71.676
R885 B.n78 B.n29 71.676
R886 B.n74 B.n28 71.676
R887 B.n70 B.n27 71.676
R888 B.n399 B.n398 71.676
R889 B.n257 B.n224 71.676
R890 B.n391 B.n225 71.676
R891 B.n387 B.n226 71.676
R892 B.n383 B.n227 71.676
R893 B.n379 B.n228 71.676
R894 B.n375 B.n229 71.676
R895 B.n371 B.n230 71.676
R896 B.n367 B.n231 71.676
R897 B.n363 B.n232 71.676
R898 B.n359 B.n233 71.676
R899 B.n355 B.n234 71.676
R900 B.n351 B.n235 71.676
R901 B.n347 B.n236 71.676
R902 B.n343 B.n237 71.676
R903 B.n338 B.n238 71.676
R904 B.n334 B.n239 71.676
R905 B.n330 B.n240 71.676
R906 B.n326 B.n241 71.676
R907 B.n322 B.n242 71.676
R908 B.n318 B.n243 71.676
R909 B.n314 B.n244 71.676
R910 B.n310 B.n245 71.676
R911 B.n306 B.n246 71.676
R912 B.n302 B.n247 71.676
R913 B.n298 B.n248 71.676
R914 B.n294 B.n249 71.676
R915 B.n290 B.n250 71.676
R916 B.n286 B.n251 71.676
R917 B.n282 B.n252 71.676
R918 B.n278 B.n253 71.676
R919 B.n274 B.n254 71.676
R920 B.n270 B.n255 71.676
R921 B.n266 B.n256 71.676
R922 B.n398 B.n223 71.676
R923 B.n392 B.n224 71.676
R924 B.n388 B.n225 71.676
R925 B.n384 B.n226 71.676
R926 B.n380 B.n227 71.676
R927 B.n376 B.n228 71.676
R928 B.n372 B.n229 71.676
R929 B.n368 B.n230 71.676
R930 B.n364 B.n231 71.676
R931 B.n360 B.n232 71.676
R932 B.n356 B.n233 71.676
R933 B.n352 B.n234 71.676
R934 B.n348 B.n235 71.676
R935 B.n344 B.n236 71.676
R936 B.n339 B.n237 71.676
R937 B.n335 B.n238 71.676
R938 B.n331 B.n239 71.676
R939 B.n327 B.n240 71.676
R940 B.n323 B.n241 71.676
R941 B.n319 B.n242 71.676
R942 B.n315 B.n243 71.676
R943 B.n311 B.n244 71.676
R944 B.n307 B.n245 71.676
R945 B.n303 B.n246 71.676
R946 B.n299 B.n247 71.676
R947 B.n295 B.n248 71.676
R948 B.n291 B.n249 71.676
R949 B.n287 B.n250 71.676
R950 B.n283 B.n251 71.676
R951 B.n279 B.n252 71.676
R952 B.n275 B.n253 71.676
R953 B.n271 B.n254 71.676
R954 B.n267 B.n255 71.676
R955 B.n263 B.n256 71.676
R956 B.n476 B.n475 71.676
R957 B.n476 B.n2 71.676
R958 B.n66 B.n65 59.5399
R959 B.n145 B.n63 59.5399
R960 B.n262 B.n261 59.5399
R961 B.n341 B.n259 59.5399
R962 B.n404 B.n220 56.6028
R963 B.n404 B.n216 56.6028
R964 B.n411 B.n216 56.6028
R965 B.n411 B.n410 56.6028
R966 B.n417 B.n209 56.6028
R967 B.n424 B.n209 56.6028
R968 B.n424 B.n205 56.6028
R969 B.n430 B.n205 56.6028
R970 B.n474 B.n4 56.6028
R971 B.n474 B.n473 56.6028
R972 B.n473 B.n472 56.6028
R973 B.n469 B.n468 56.6028
R974 B.n468 B.n467 56.6028
R975 B.n467 B.n13 56.6028
R976 B.n461 B.n13 56.6028
R977 B.n460 B.n459 56.6028
R978 B.n459 B.n21 56.6028
R979 B.n453 B.n21 56.6028
R980 B.n453 B.n452 56.6028
R981 B.t0 B.n4 52.4409
R982 B.n472 B.t1 52.4409
R983 B.n417 B.t3 44.117
R984 B.n461 B.t7 44.117
R985 B.n401 B.n400 31.0639
R986 B.n264 B.n218 31.0639
R987 B.n449 B.n448 31.0639
R988 B.n68 B.n23 31.0639
R989 B B.n477 18.0485
R990 B.n410 B.t3 12.4863
R991 B.t7 B.n460 12.4863
R992 B.n65 B.n64 10.8611
R993 B.n63 B.n62 10.8611
R994 B.n261 B.n260 10.8611
R995 B.n259 B.n258 10.8611
R996 B.n402 B.n401 10.6151
R997 B.n402 B.n214 10.6151
R998 B.n413 B.n214 10.6151
R999 B.n414 B.n413 10.6151
R1000 B.n415 B.n414 10.6151
R1001 B.n415 B.n207 10.6151
R1002 B.n426 B.n207 10.6151
R1003 B.n427 B.n426 10.6151
R1004 B.n428 B.n427 10.6151
R1005 B.n428 B.n0 10.6151
R1006 B.n400 B.n222 10.6151
R1007 B.n395 B.n222 10.6151
R1008 B.n395 B.n394 10.6151
R1009 B.n394 B.n393 10.6151
R1010 B.n393 B.n390 10.6151
R1011 B.n390 B.n389 10.6151
R1012 B.n389 B.n386 10.6151
R1013 B.n386 B.n385 10.6151
R1014 B.n385 B.n382 10.6151
R1015 B.n382 B.n381 10.6151
R1016 B.n381 B.n378 10.6151
R1017 B.n378 B.n377 10.6151
R1018 B.n377 B.n374 10.6151
R1019 B.n374 B.n373 10.6151
R1020 B.n373 B.n370 10.6151
R1021 B.n370 B.n369 10.6151
R1022 B.n369 B.n366 10.6151
R1023 B.n366 B.n365 10.6151
R1024 B.n365 B.n362 10.6151
R1025 B.n362 B.n361 10.6151
R1026 B.n361 B.n358 10.6151
R1027 B.n358 B.n357 10.6151
R1028 B.n357 B.n354 10.6151
R1029 B.n354 B.n353 10.6151
R1030 B.n353 B.n350 10.6151
R1031 B.n350 B.n349 10.6151
R1032 B.n349 B.n346 10.6151
R1033 B.n346 B.n345 10.6151
R1034 B.n345 B.n342 10.6151
R1035 B.n340 B.n337 10.6151
R1036 B.n337 B.n336 10.6151
R1037 B.n336 B.n333 10.6151
R1038 B.n333 B.n332 10.6151
R1039 B.n332 B.n329 10.6151
R1040 B.n329 B.n328 10.6151
R1041 B.n328 B.n325 10.6151
R1042 B.n325 B.n324 10.6151
R1043 B.n321 B.n320 10.6151
R1044 B.n320 B.n317 10.6151
R1045 B.n317 B.n316 10.6151
R1046 B.n316 B.n313 10.6151
R1047 B.n313 B.n312 10.6151
R1048 B.n312 B.n309 10.6151
R1049 B.n309 B.n308 10.6151
R1050 B.n308 B.n305 10.6151
R1051 B.n305 B.n304 10.6151
R1052 B.n304 B.n301 10.6151
R1053 B.n301 B.n300 10.6151
R1054 B.n300 B.n297 10.6151
R1055 B.n297 B.n296 10.6151
R1056 B.n296 B.n293 10.6151
R1057 B.n293 B.n292 10.6151
R1058 B.n292 B.n289 10.6151
R1059 B.n289 B.n288 10.6151
R1060 B.n288 B.n285 10.6151
R1061 B.n285 B.n284 10.6151
R1062 B.n284 B.n281 10.6151
R1063 B.n281 B.n280 10.6151
R1064 B.n280 B.n277 10.6151
R1065 B.n277 B.n276 10.6151
R1066 B.n276 B.n273 10.6151
R1067 B.n273 B.n272 10.6151
R1068 B.n272 B.n269 10.6151
R1069 B.n269 B.n268 10.6151
R1070 B.n268 B.n265 10.6151
R1071 B.n265 B.n264 10.6151
R1072 B.n406 B.n218 10.6151
R1073 B.n407 B.n406 10.6151
R1074 B.n408 B.n407 10.6151
R1075 B.n408 B.n211 10.6151
R1076 B.n419 B.n211 10.6151
R1077 B.n420 B.n419 10.6151
R1078 B.n422 B.n420 10.6151
R1079 B.n422 B.n421 10.6151
R1080 B.n421 B.n203 10.6151
R1081 B.n433 B.n203 10.6151
R1082 B.n434 B.n433 10.6151
R1083 B.n435 B.n434 10.6151
R1084 B.n436 B.n435 10.6151
R1085 B.n437 B.n436 10.6151
R1086 B.n438 B.n437 10.6151
R1087 B.n439 B.n438 10.6151
R1088 B.n441 B.n439 10.6151
R1089 B.n442 B.n441 10.6151
R1090 B.n443 B.n442 10.6151
R1091 B.n444 B.n443 10.6151
R1092 B.n446 B.n444 10.6151
R1093 B.n447 B.n446 10.6151
R1094 B.n448 B.n447 10.6151
R1095 B.n9 B.n1 10.6151
R1096 B.n15 B.n9 10.6151
R1097 B.n465 B.n15 10.6151
R1098 B.n465 B.n464 10.6151
R1099 B.n464 B.n463 10.6151
R1100 B.n463 B.n16 10.6151
R1101 B.n457 B.n16 10.6151
R1102 B.n457 B.n456 10.6151
R1103 B.n456 B.n455 10.6151
R1104 B.n455 B.n23 10.6151
R1105 B.n69 B.n68 10.6151
R1106 B.n72 B.n69 10.6151
R1107 B.n73 B.n72 10.6151
R1108 B.n76 B.n73 10.6151
R1109 B.n77 B.n76 10.6151
R1110 B.n80 B.n77 10.6151
R1111 B.n81 B.n80 10.6151
R1112 B.n84 B.n81 10.6151
R1113 B.n85 B.n84 10.6151
R1114 B.n88 B.n85 10.6151
R1115 B.n89 B.n88 10.6151
R1116 B.n92 B.n89 10.6151
R1117 B.n93 B.n92 10.6151
R1118 B.n96 B.n93 10.6151
R1119 B.n97 B.n96 10.6151
R1120 B.n100 B.n97 10.6151
R1121 B.n101 B.n100 10.6151
R1122 B.n104 B.n101 10.6151
R1123 B.n105 B.n104 10.6151
R1124 B.n108 B.n105 10.6151
R1125 B.n109 B.n108 10.6151
R1126 B.n112 B.n109 10.6151
R1127 B.n113 B.n112 10.6151
R1128 B.n116 B.n113 10.6151
R1129 B.n117 B.n116 10.6151
R1130 B.n120 B.n117 10.6151
R1131 B.n121 B.n120 10.6151
R1132 B.n124 B.n121 10.6151
R1133 B.n125 B.n124 10.6151
R1134 B.n129 B.n128 10.6151
R1135 B.n132 B.n129 10.6151
R1136 B.n133 B.n132 10.6151
R1137 B.n136 B.n133 10.6151
R1138 B.n137 B.n136 10.6151
R1139 B.n140 B.n137 10.6151
R1140 B.n141 B.n140 10.6151
R1141 B.n144 B.n141 10.6151
R1142 B.n149 B.n146 10.6151
R1143 B.n150 B.n149 10.6151
R1144 B.n153 B.n150 10.6151
R1145 B.n154 B.n153 10.6151
R1146 B.n157 B.n154 10.6151
R1147 B.n158 B.n157 10.6151
R1148 B.n161 B.n158 10.6151
R1149 B.n162 B.n161 10.6151
R1150 B.n165 B.n162 10.6151
R1151 B.n166 B.n165 10.6151
R1152 B.n169 B.n166 10.6151
R1153 B.n170 B.n169 10.6151
R1154 B.n173 B.n170 10.6151
R1155 B.n174 B.n173 10.6151
R1156 B.n177 B.n174 10.6151
R1157 B.n178 B.n177 10.6151
R1158 B.n181 B.n178 10.6151
R1159 B.n182 B.n181 10.6151
R1160 B.n185 B.n182 10.6151
R1161 B.n186 B.n185 10.6151
R1162 B.n189 B.n186 10.6151
R1163 B.n190 B.n189 10.6151
R1164 B.n193 B.n190 10.6151
R1165 B.n194 B.n193 10.6151
R1166 B.n197 B.n194 10.6151
R1167 B.n198 B.n197 10.6151
R1168 B.n201 B.n198 10.6151
R1169 B.n202 B.n201 10.6151
R1170 B.n449 B.n202 10.6151
R1171 B.n477 B.n0 8.11757
R1172 B.n477 B.n1 8.11757
R1173 B.n341 B.n340 7.18099
R1174 B.n324 B.n262 7.18099
R1175 B.n128 B.n66 7.18099
R1176 B.n145 B.n144 7.18099
R1177 B.n430 B.t0 4.16244
R1178 B.n469 B.t1 4.16244
R1179 B.n342 B.n341 3.43465
R1180 B.n321 B.n262 3.43465
R1181 B.n125 B.n66 3.43465
R1182 B.n146 B.n145 3.43465
R1183 VP.n0 VP.t1 1186.79
R1184 VP.n0 VP.t0 1151.5
R1185 VP VP.n0 0.0516364
R1186 VDD1.n36 VDD1.n0 289.615
R1187 VDD1.n77 VDD1.n41 289.615
R1188 VDD1.n37 VDD1.n36 185
R1189 VDD1.n35 VDD1.n2 185
R1190 VDD1.n34 VDD1.n33 185
R1191 VDD1.n5 VDD1.n3 185
R1192 VDD1.n28 VDD1.n27 185
R1193 VDD1.n26 VDD1.n25 185
R1194 VDD1.n9 VDD1.n8 185
R1195 VDD1.n20 VDD1.n19 185
R1196 VDD1.n18 VDD1.n17 185
R1197 VDD1.n13 VDD1.n12 185
R1198 VDD1.n53 VDD1.n52 185
R1199 VDD1.n58 VDD1.n57 185
R1200 VDD1.n60 VDD1.n59 185
R1201 VDD1.n49 VDD1.n48 185
R1202 VDD1.n66 VDD1.n65 185
R1203 VDD1.n68 VDD1.n67 185
R1204 VDD1.n45 VDD1.n44 185
R1205 VDD1.n75 VDD1.n74 185
R1206 VDD1.n76 VDD1.n43 185
R1207 VDD1.n78 VDD1.n77 185
R1208 VDD1.n14 VDD1.t0 149.524
R1209 VDD1.n54 VDD1.t1 149.524
R1210 VDD1.n36 VDD1.n35 104.615
R1211 VDD1.n35 VDD1.n34 104.615
R1212 VDD1.n34 VDD1.n3 104.615
R1213 VDD1.n27 VDD1.n3 104.615
R1214 VDD1.n27 VDD1.n26 104.615
R1215 VDD1.n26 VDD1.n8 104.615
R1216 VDD1.n19 VDD1.n8 104.615
R1217 VDD1.n19 VDD1.n18 104.615
R1218 VDD1.n18 VDD1.n12 104.615
R1219 VDD1.n58 VDD1.n52 104.615
R1220 VDD1.n59 VDD1.n58 104.615
R1221 VDD1.n59 VDD1.n48 104.615
R1222 VDD1.n66 VDD1.n48 104.615
R1223 VDD1.n67 VDD1.n66 104.615
R1224 VDD1.n67 VDD1.n44 104.615
R1225 VDD1.n75 VDD1.n44 104.615
R1226 VDD1.n76 VDD1.n75 104.615
R1227 VDD1.n77 VDD1.n76 104.615
R1228 VDD1 VDD1.n81 83.3067
R1229 VDD1.t0 VDD1.n12 52.3082
R1230 VDD1.t1 VDD1.n52 52.3082
R1231 VDD1 VDD1.n40 51.3703
R1232 VDD1.n37 VDD1.n2 13.1884
R1233 VDD1.n78 VDD1.n43 13.1884
R1234 VDD1.n38 VDD1.n0 12.8005
R1235 VDD1.n33 VDD1.n4 12.8005
R1236 VDD1.n74 VDD1.n73 12.8005
R1237 VDD1.n79 VDD1.n41 12.8005
R1238 VDD1.n32 VDD1.n5 12.0247
R1239 VDD1.n72 VDD1.n45 12.0247
R1240 VDD1.n29 VDD1.n28 11.249
R1241 VDD1.n69 VDD1.n68 11.249
R1242 VDD1.n25 VDD1.n7 10.4732
R1243 VDD1.n65 VDD1.n47 10.4732
R1244 VDD1.n14 VDD1.n13 10.2747
R1245 VDD1.n54 VDD1.n53 10.2747
R1246 VDD1.n24 VDD1.n9 9.69747
R1247 VDD1.n64 VDD1.n49 9.69747
R1248 VDD1.n40 VDD1.n39 9.45567
R1249 VDD1.n81 VDD1.n80 9.45567
R1250 VDD1.n16 VDD1.n15 9.3005
R1251 VDD1.n11 VDD1.n10 9.3005
R1252 VDD1.n22 VDD1.n21 9.3005
R1253 VDD1.n24 VDD1.n23 9.3005
R1254 VDD1.n7 VDD1.n6 9.3005
R1255 VDD1.n30 VDD1.n29 9.3005
R1256 VDD1.n32 VDD1.n31 9.3005
R1257 VDD1.n4 VDD1.n1 9.3005
R1258 VDD1.n39 VDD1.n38 9.3005
R1259 VDD1.n80 VDD1.n79 9.3005
R1260 VDD1.n56 VDD1.n55 9.3005
R1261 VDD1.n51 VDD1.n50 9.3005
R1262 VDD1.n62 VDD1.n61 9.3005
R1263 VDD1.n64 VDD1.n63 9.3005
R1264 VDD1.n47 VDD1.n46 9.3005
R1265 VDD1.n70 VDD1.n69 9.3005
R1266 VDD1.n72 VDD1.n71 9.3005
R1267 VDD1.n73 VDD1.n42 9.3005
R1268 VDD1.n21 VDD1.n20 8.92171
R1269 VDD1.n61 VDD1.n60 8.92171
R1270 VDD1.n17 VDD1.n11 8.14595
R1271 VDD1.n57 VDD1.n51 8.14595
R1272 VDD1.n16 VDD1.n13 7.3702
R1273 VDD1.n56 VDD1.n53 7.3702
R1274 VDD1.n17 VDD1.n16 5.81868
R1275 VDD1.n57 VDD1.n56 5.81868
R1276 VDD1.n20 VDD1.n11 5.04292
R1277 VDD1.n60 VDD1.n51 5.04292
R1278 VDD1.n21 VDD1.n9 4.26717
R1279 VDD1.n61 VDD1.n49 4.26717
R1280 VDD1.n25 VDD1.n24 3.49141
R1281 VDD1.n65 VDD1.n64 3.49141
R1282 VDD1.n15 VDD1.n14 2.84304
R1283 VDD1.n55 VDD1.n54 2.84304
R1284 VDD1.n28 VDD1.n7 2.71565
R1285 VDD1.n68 VDD1.n47 2.71565
R1286 VDD1.n29 VDD1.n5 1.93989
R1287 VDD1.n69 VDD1.n45 1.93989
R1288 VDD1.n40 VDD1.n0 1.16414
R1289 VDD1.n33 VDD1.n32 1.16414
R1290 VDD1.n74 VDD1.n72 1.16414
R1291 VDD1.n81 VDD1.n41 1.16414
R1292 VDD1.n38 VDD1.n37 0.388379
R1293 VDD1.n4 VDD1.n2 0.388379
R1294 VDD1.n73 VDD1.n43 0.388379
R1295 VDD1.n79 VDD1.n78 0.388379
R1296 VDD1.n39 VDD1.n1 0.155672
R1297 VDD1.n31 VDD1.n1 0.155672
R1298 VDD1.n31 VDD1.n30 0.155672
R1299 VDD1.n30 VDD1.n6 0.155672
R1300 VDD1.n23 VDD1.n6 0.155672
R1301 VDD1.n23 VDD1.n22 0.155672
R1302 VDD1.n22 VDD1.n10 0.155672
R1303 VDD1.n15 VDD1.n10 0.155672
R1304 VDD1.n55 VDD1.n50 0.155672
R1305 VDD1.n62 VDD1.n50 0.155672
R1306 VDD1.n63 VDD1.n62 0.155672
R1307 VDD1.n63 VDD1.n46 0.155672
R1308 VDD1.n70 VDD1.n46 0.155672
R1309 VDD1.n71 VDD1.n70 0.155672
R1310 VDD1.n71 VDD1.n42 0.155672
R1311 VDD1.n80 VDD1.n42 0.155672
C0 VN VDD2 0.946296f
C1 VTAIL VP 0.56074f
C2 VDD1 VP 1.02928f
C3 VN VP 3.59743f
C4 VDD2 VP 0.235103f
C5 VDD1 VTAIL 5.29332f
C6 VN VTAIL 0.546181f
C7 VDD2 VTAIL 5.32483f
C8 VN VDD1 0.148693f
C9 VDD2 VDD1 0.419138f
C10 VDD2 B 2.838081f
C11 VDD1 B 4.75444f
C12 VTAIL B 4.238245f
C13 VN B 6.34518f
C14 VP B 3.218185f
C15 VDD1.n0 B 0.026755f
C16 VDD1.n1 B 0.020198f
C17 VDD1.n2 B 0.011173f
C18 VDD1.n3 B 0.025654f
C19 VDD1.n4 B 0.010854f
C20 VDD1.n5 B 0.011492f
C21 VDD1.n6 B 0.020198f
C22 VDD1.n7 B 0.010854f
C23 VDD1.n8 B 0.025654f
C24 VDD1.n9 B 0.011492f
C25 VDD1.n10 B 0.020198f
C26 VDD1.n11 B 0.010854f
C27 VDD1.n12 B 0.01924f
C28 VDD1.n13 B 0.018135f
C29 VDD1.t0 B 0.042897f
C30 VDD1.n14 B 0.114011f
C31 VDD1.n15 B 0.652375f
C32 VDD1.n16 B 0.010854f
C33 VDD1.n17 B 0.011492f
C34 VDD1.n18 B 0.025654f
C35 VDD1.n19 B 0.025654f
C36 VDD1.n20 B 0.011492f
C37 VDD1.n21 B 0.010854f
C38 VDD1.n22 B 0.020198f
C39 VDD1.n23 B 0.020198f
C40 VDD1.n24 B 0.010854f
C41 VDD1.n25 B 0.011492f
C42 VDD1.n26 B 0.025654f
C43 VDD1.n27 B 0.025654f
C44 VDD1.n28 B 0.011492f
C45 VDD1.n29 B 0.010854f
C46 VDD1.n30 B 0.020198f
C47 VDD1.n31 B 0.020198f
C48 VDD1.n32 B 0.010854f
C49 VDD1.n33 B 0.011492f
C50 VDD1.n34 B 0.025654f
C51 VDD1.n35 B 0.025654f
C52 VDD1.n36 B 0.052644f
C53 VDD1.n37 B 0.011173f
C54 VDD1.n38 B 0.010854f
C55 VDD1.n39 B 0.049998f
C56 VDD1.n40 B 0.043362f
C57 VDD1.n41 B 0.026755f
C58 VDD1.n42 B 0.020198f
C59 VDD1.n43 B 0.011173f
C60 VDD1.n44 B 0.025654f
C61 VDD1.n45 B 0.011492f
C62 VDD1.n46 B 0.020198f
C63 VDD1.n47 B 0.010854f
C64 VDD1.n48 B 0.025654f
C65 VDD1.n49 B 0.011492f
C66 VDD1.n50 B 0.020198f
C67 VDD1.n51 B 0.010854f
C68 VDD1.n52 B 0.01924f
C69 VDD1.n53 B 0.018135f
C70 VDD1.t1 B 0.042897f
C71 VDD1.n54 B 0.114011f
C72 VDD1.n55 B 0.652375f
C73 VDD1.n56 B 0.010854f
C74 VDD1.n57 B 0.011492f
C75 VDD1.n58 B 0.025654f
C76 VDD1.n59 B 0.025654f
C77 VDD1.n60 B 0.011492f
C78 VDD1.n61 B 0.010854f
C79 VDD1.n62 B 0.020198f
C80 VDD1.n63 B 0.020198f
C81 VDD1.n64 B 0.010854f
C82 VDD1.n65 B 0.011492f
C83 VDD1.n66 B 0.025654f
C84 VDD1.n67 B 0.025654f
C85 VDD1.n68 B 0.011492f
C86 VDD1.n69 B 0.010854f
C87 VDD1.n70 B 0.020198f
C88 VDD1.n71 B 0.020198f
C89 VDD1.n72 B 0.010854f
C90 VDD1.n73 B 0.010854f
C91 VDD1.n74 B 0.011492f
C92 VDD1.n75 B 0.025654f
C93 VDD1.n76 B 0.025654f
C94 VDD1.n77 B 0.052644f
C95 VDD1.n78 B 0.011173f
C96 VDD1.n79 B 0.010854f
C97 VDD1.n80 B 0.049998f
C98 VDD1.n81 B 0.381511f
C99 VP.t1 B 0.306131f
C100 VP.t0 B 0.261086f
C101 VP.n0 B 3.02713f
C102 VDD2.n0 B 0.027137f
C103 VDD2.n1 B 0.020486f
C104 VDD2.n2 B 0.011332f
C105 VDD2.n3 B 0.02602f
C106 VDD2.n4 B 0.011656f
C107 VDD2.n5 B 0.020486f
C108 VDD2.n6 B 0.011008f
C109 VDD2.n7 B 0.02602f
C110 VDD2.n8 B 0.011656f
C111 VDD2.n9 B 0.020486f
C112 VDD2.n10 B 0.011008f
C113 VDD2.n11 B 0.019515f
C114 VDD2.n12 B 0.018394f
C115 VDD2.t0 B 0.043509f
C116 VDD2.n13 B 0.115638f
C117 VDD2.n14 B 0.661689f
C118 VDD2.n15 B 0.011008f
C119 VDD2.n16 B 0.011656f
C120 VDD2.n17 B 0.02602f
C121 VDD2.n18 B 0.02602f
C122 VDD2.n19 B 0.011656f
C123 VDD2.n20 B 0.011008f
C124 VDD2.n21 B 0.020486f
C125 VDD2.n22 B 0.020486f
C126 VDD2.n23 B 0.011008f
C127 VDD2.n24 B 0.011656f
C128 VDD2.n25 B 0.02602f
C129 VDD2.n26 B 0.02602f
C130 VDD2.n27 B 0.011656f
C131 VDD2.n28 B 0.011008f
C132 VDD2.n29 B 0.020486f
C133 VDD2.n30 B 0.020486f
C134 VDD2.n31 B 0.011008f
C135 VDD2.n32 B 0.011008f
C136 VDD2.n33 B 0.011656f
C137 VDD2.n34 B 0.02602f
C138 VDD2.n35 B 0.02602f
C139 VDD2.n36 B 0.053396f
C140 VDD2.n37 B 0.011332f
C141 VDD2.n38 B 0.011008f
C142 VDD2.n39 B 0.050711f
C143 VDD2.n40 B 0.364848f
C144 VDD2.n41 B 0.027137f
C145 VDD2.n42 B 0.020486f
C146 VDD2.n43 B 0.011332f
C147 VDD2.n44 B 0.02602f
C148 VDD2.n45 B 0.011008f
C149 VDD2.n46 B 0.011656f
C150 VDD2.n47 B 0.020486f
C151 VDD2.n48 B 0.011008f
C152 VDD2.n49 B 0.02602f
C153 VDD2.n50 B 0.011656f
C154 VDD2.n51 B 0.020486f
C155 VDD2.n52 B 0.011008f
C156 VDD2.n53 B 0.019515f
C157 VDD2.n54 B 0.018394f
C158 VDD2.t1 B 0.043509f
C159 VDD2.n55 B 0.115638f
C160 VDD2.n56 B 0.661689f
C161 VDD2.n57 B 0.011008f
C162 VDD2.n58 B 0.011656f
C163 VDD2.n59 B 0.02602f
C164 VDD2.n60 B 0.02602f
C165 VDD2.n61 B 0.011656f
C166 VDD2.n62 B 0.011008f
C167 VDD2.n63 B 0.020486f
C168 VDD2.n64 B 0.020486f
C169 VDD2.n65 B 0.011008f
C170 VDD2.n66 B 0.011656f
C171 VDD2.n67 B 0.02602f
C172 VDD2.n68 B 0.02602f
C173 VDD2.n69 B 0.011656f
C174 VDD2.n70 B 0.011008f
C175 VDD2.n71 B 0.020486f
C176 VDD2.n72 B 0.020486f
C177 VDD2.n73 B 0.011008f
C178 VDD2.n74 B 0.011656f
C179 VDD2.n75 B 0.02602f
C180 VDD2.n76 B 0.02602f
C181 VDD2.n77 B 0.053396f
C182 VDD2.n78 B 0.011332f
C183 VDD2.n79 B 0.011008f
C184 VDD2.n80 B 0.050711f
C185 VDD2.n81 B 0.043796f
C186 VDD2.n82 B 1.77328f
C187 VTAIL.n0 B 0.02973f
C188 VTAIL.n1 B 0.022444f
C189 VTAIL.n2 B 0.012415f
C190 VTAIL.n3 B 0.028507f
C191 VTAIL.n4 B 0.01277f
C192 VTAIL.n5 B 0.022444f
C193 VTAIL.n6 B 0.012061f
C194 VTAIL.n7 B 0.028507f
C195 VTAIL.n8 B 0.01277f
C196 VTAIL.n9 B 0.022444f
C197 VTAIL.n10 B 0.012061f
C198 VTAIL.n11 B 0.02138f
C199 VTAIL.n12 B 0.020152f
C200 VTAIL.t0 B 0.047668f
C201 VTAIL.n13 B 0.12669f
C202 VTAIL.n14 B 0.72493f
C203 VTAIL.n15 B 0.012061f
C204 VTAIL.n16 B 0.01277f
C205 VTAIL.n17 B 0.028507f
C206 VTAIL.n18 B 0.028507f
C207 VTAIL.n19 B 0.01277f
C208 VTAIL.n20 B 0.012061f
C209 VTAIL.n21 B 0.022444f
C210 VTAIL.n22 B 0.022444f
C211 VTAIL.n23 B 0.012061f
C212 VTAIL.n24 B 0.01277f
C213 VTAIL.n25 B 0.028507f
C214 VTAIL.n26 B 0.028507f
C215 VTAIL.n27 B 0.01277f
C216 VTAIL.n28 B 0.012061f
C217 VTAIL.n29 B 0.022444f
C218 VTAIL.n30 B 0.022444f
C219 VTAIL.n31 B 0.012061f
C220 VTAIL.n32 B 0.012061f
C221 VTAIL.n33 B 0.01277f
C222 VTAIL.n34 B 0.028507f
C223 VTAIL.n35 B 0.028507f
C224 VTAIL.n36 B 0.058499f
C225 VTAIL.n37 B 0.012415f
C226 VTAIL.n38 B 0.012061f
C227 VTAIL.n39 B 0.055558f
C228 VTAIL.n40 B 0.032512f
C229 VTAIL.n41 B 0.937889f
C230 VTAIL.n42 B 0.02973f
C231 VTAIL.n43 B 0.022444f
C232 VTAIL.n44 B 0.012415f
C233 VTAIL.n45 B 0.028507f
C234 VTAIL.n46 B 0.012061f
C235 VTAIL.n47 B 0.01277f
C236 VTAIL.n48 B 0.022444f
C237 VTAIL.n49 B 0.012061f
C238 VTAIL.n50 B 0.028507f
C239 VTAIL.n51 B 0.01277f
C240 VTAIL.n52 B 0.022444f
C241 VTAIL.n53 B 0.012061f
C242 VTAIL.n54 B 0.02138f
C243 VTAIL.n55 B 0.020152f
C244 VTAIL.t1 B 0.047668f
C245 VTAIL.n56 B 0.12669f
C246 VTAIL.n57 B 0.72493f
C247 VTAIL.n58 B 0.012061f
C248 VTAIL.n59 B 0.01277f
C249 VTAIL.n60 B 0.028507f
C250 VTAIL.n61 B 0.028507f
C251 VTAIL.n62 B 0.01277f
C252 VTAIL.n63 B 0.012061f
C253 VTAIL.n64 B 0.022444f
C254 VTAIL.n65 B 0.022444f
C255 VTAIL.n66 B 0.012061f
C256 VTAIL.n67 B 0.01277f
C257 VTAIL.n68 B 0.028507f
C258 VTAIL.n69 B 0.028507f
C259 VTAIL.n70 B 0.01277f
C260 VTAIL.n71 B 0.012061f
C261 VTAIL.n72 B 0.022444f
C262 VTAIL.n73 B 0.022444f
C263 VTAIL.n74 B 0.012061f
C264 VTAIL.n75 B 0.01277f
C265 VTAIL.n76 B 0.028507f
C266 VTAIL.n77 B 0.028507f
C267 VTAIL.n78 B 0.058499f
C268 VTAIL.n79 B 0.012415f
C269 VTAIL.n80 B 0.012061f
C270 VTAIL.n81 B 0.055558f
C271 VTAIL.n82 B 0.032512f
C272 VTAIL.n83 B 0.942409f
C273 VTAIL.n84 B 0.02973f
C274 VTAIL.n85 B 0.022444f
C275 VTAIL.n86 B 0.012415f
C276 VTAIL.n87 B 0.028507f
C277 VTAIL.n88 B 0.012061f
C278 VTAIL.n89 B 0.01277f
C279 VTAIL.n90 B 0.022444f
C280 VTAIL.n91 B 0.012061f
C281 VTAIL.n92 B 0.028507f
C282 VTAIL.n93 B 0.01277f
C283 VTAIL.n94 B 0.022444f
C284 VTAIL.n95 B 0.012061f
C285 VTAIL.n96 B 0.02138f
C286 VTAIL.n97 B 0.020152f
C287 VTAIL.t3 B 0.047668f
C288 VTAIL.n98 B 0.12669f
C289 VTAIL.n99 B 0.72493f
C290 VTAIL.n100 B 0.012061f
C291 VTAIL.n101 B 0.01277f
C292 VTAIL.n102 B 0.028507f
C293 VTAIL.n103 B 0.028507f
C294 VTAIL.n104 B 0.01277f
C295 VTAIL.n105 B 0.012061f
C296 VTAIL.n106 B 0.022444f
C297 VTAIL.n107 B 0.022444f
C298 VTAIL.n108 B 0.012061f
C299 VTAIL.n109 B 0.01277f
C300 VTAIL.n110 B 0.028507f
C301 VTAIL.n111 B 0.028507f
C302 VTAIL.n112 B 0.01277f
C303 VTAIL.n113 B 0.012061f
C304 VTAIL.n114 B 0.022444f
C305 VTAIL.n115 B 0.022444f
C306 VTAIL.n116 B 0.012061f
C307 VTAIL.n117 B 0.01277f
C308 VTAIL.n118 B 0.028507f
C309 VTAIL.n119 B 0.028507f
C310 VTAIL.n120 B 0.058499f
C311 VTAIL.n121 B 0.012415f
C312 VTAIL.n122 B 0.012061f
C313 VTAIL.n123 B 0.055558f
C314 VTAIL.n124 B 0.032512f
C315 VTAIL.n125 B 0.907496f
C316 VTAIL.n126 B 0.02973f
C317 VTAIL.n127 B 0.022444f
C318 VTAIL.n128 B 0.012415f
C319 VTAIL.n129 B 0.028507f
C320 VTAIL.n130 B 0.01277f
C321 VTAIL.n131 B 0.022444f
C322 VTAIL.n132 B 0.012061f
C323 VTAIL.n133 B 0.028507f
C324 VTAIL.n134 B 0.01277f
C325 VTAIL.n135 B 0.022444f
C326 VTAIL.n136 B 0.012061f
C327 VTAIL.n137 B 0.02138f
C328 VTAIL.n138 B 0.020152f
C329 VTAIL.t2 B 0.047668f
C330 VTAIL.n139 B 0.12669f
C331 VTAIL.n140 B 0.72493f
C332 VTAIL.n141 B 0.012061f
C333 VTAIL.n142 B 0.01277f
C334 VTAIL.n143 B 0.028507f
C335 VTAIL.n144 B 0.028507f
C336 VTAIL.n145 B 0.01277f
C337 VTAIL.n146 B 0.012061f
C338 VTAIL.n147 B 0.022444f
C339 VTAIL.n148 B 0.022444f
C340 VTAIL.n149 B 0.012061f
C341 VTAIL.n150 B 0.01277f
C342 VTAIL.n151 B 0.028507f
C343 VTAIL.n152 B 0.028507f
C344 VTAIL.n153 B 0.01277f
C345 VTAIL.n154 B 0.012061f
C346 VTAIL.n155 B 0.022444f
C347 VTAIL.n156 B 0.022444f
C348 VTAIL.n157 B 0.012061f
C349 VTAIL.n158 B 0.012061f
C350 VTAIL.n159 B 0.01277f
C351 VTAIL.n160 B 0.028507f
C352 VTAIL.n161 B 0.028507f
C353 VTAIL.n162 B 0.058499f
C354 VTAIL.n163 B 0.012415f
C355 VTAIL.n164 B 0.012061f
C356 VTAIL.n165 B 0.055558f
C357 VTAIL.n166 B 0.032512f
C358 VTAIL.n167 B 0.860581f
C359 VN.t1 B 0.256383f
C360 VN.t0 B 0.301995f
.ends

