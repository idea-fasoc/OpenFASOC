* NGSPICE file created from diff_pair_sample_1732.ext - technology: sky130A

.subckt diff_pair_sample_1732 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t9 VN.t0 VDD2.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.0593 pd=6.75 as=1.0593 ps=6.75 w=6.42 l=1.33
X1 VDD2.t5 VN.t1 VTAIL.t8 B.t3 sky130_fd_pr__nfet_01v8 ad=1.0593 pd=6.75 as=2.5038 ps=13.62 w=6.42 l=1.33
X2 VDD2.t3 VN.t2 VTAIL.t7 B.t19 sky130_fd_pr__nfet_01v8 ad=2.5038 pd=13.62 as=1.0593 ps=6.75 w=6.42 l=1.33
X3 VTAIL.t6 VN.t3 VDD2.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.0593 pd=6.75 as=1.0593 ps=6.75 w=6.42 l=1.33
X4 VTAIL.t0 VP.t0 VDD1.t5 B.t0 sky130_fd_pr__nfet_01v8 ad=1.0593 pd=6.75 as=1.0593 ps=6.75 w=6.42 l=1.33
X5 B.t17 B.t15 B.t16 B.t5 sky130_fd_pr__nfet_01v8 ad=2.5038 pd=13.62 as=0 ps=0 w=6.42 l=1.33
X6 VDD1.t4 VP.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.0593 pd=6.75 as=2.5038 ps=13.62 w=6.42 l=1.33
X7 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=2.5038 pd=13.62 as=0 ps=0 w=6.42 l=1.33
X8 VDD1.t3 VP.t2 VTAIL.t11 B.t19 sky130_fd_pr__nfet_01v8 ad=2.5038 pd=13.62 as=1.0593 ps=6.75 w=6.42 l=1.33
X9 VDD2.t4 VN.t4 VTAIL.t5 B.t1 sky130_fd_pr__nfet_01v8 ad=1.0593 pd=6.75 as=2.5038 ps=13.62 w=6.42 l=1.33
X10 VDD2.t1 VN.t5 VTAIL.t4 B.t18 sky130_fd_pr__nfet_01v8 ad=2.5038 pd=13.62 as=1.0593 ps=6.75 w=6.42 l=1.33
X11 VDD1.t2 VP.t3 VTAIL.t10 B.t18 sky130_fd_pr__nfet_01v8 ad=2.5038 pd=13.62 as=1.0593 ps=6.75 w=6.42 l=1.33
X12 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=2.5038 pd=13.62 as=0 ps=0 w=6.42 l=1.33
X13 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=2.5038 pd=13.62 as=0 ps=0 w=6.42 l=1.33
X14 VTAIL.t2 VP.t4 VDD1.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=1.0593 pd=6.75 as=1.0593 ps=6.75 w=6.42 l=1.33
X15 VDD1.t0 VP.t5 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.0593 pd=6.75 as=2.5038 ps=13.62 w=6.42 l=1.33
R0 VN.n9 VN.n8 178.023
R1 VN.n19 VN.n18 178.023
R2 VN.n17 VN.n10 161.3
R3 VN.n16 VN.n15 161.3
R4 VN.n14 VN.n11 161.3
R5 VN.n7 VN.n0 161.3
R6 VN.n6 VN.n5 161.3
R7 VN.n4 VN.n1 161.3
R8 VN.n3 VN.t5 148.995
R9 VN.n13 VN.t4 148.995
R10 VN.n2 VN.t0 116.332
R11 VN.n8 VN.t1 116.332
R12 VN.n12 VN.t3 116.332
R13 VN.n18 VN.t2 116.332
R14 VN.n6 VN.n1 56.5617
R15 VN.n16 VN.n11 56.5617
R16 VN.n3 VN.n2 41.7772
R17 VN.n13 VN.n12 41.7772
R18 VN VN.n19 39.6994
R19 VN.n2 VN.n1 24.5923
R20 VN.n7 VN.n6 24.5923
R21 VN.n12 VN.n11 24.5923
R22 VN.n17 VN.n16 24.5923
R23 VN.n14 VN.n13 17.9746
R24 VN.n4 VN.n3 17.9746
R25 VN.n8 VN.n7 7.86989
R26 VN.n18 VN.n17 7.86989
R27 VN.n19 VN.n10 0.189894
R28 VN.n15 VN.n10 0.189894
R29 VN.n15 VN.n14 0.189894
R30 VN.n5 VN.n4 0.189894
R31 VN.n5 VN.n0 0.189894
R32 VN.n9 VN.n0 0.189894
R33 VN VN.n9 0.0516364
R34 VDD2.n1 VDD2.t1 71.8616
R35 VDD2.n2 VDD2.t3 70.8437
R36 VDD2.n1 VDD2.n0 68.0619
R37 VDD2 VDD2.n3 68.0591
R38 VDD2.n2 VDD2.n1 33.9006
R39 VDD2.n3 VDD2.t2 3.08461
R40 VDD2.n3 VDD2.t4 3.08461
R41 VDD2.n0 VDD2.t0 3.08461
R42 VDD2.n0 VDD2.t5 3.08461
R43 VDD2 VDD2.n2 1.13197
R44 VTAIL.n7 VTAIL.t5 54.165
R45 VTAIL.n10 VTAIL.t3 54.1649
R46 VTAIL.n11 VTAIL.t8 54.1648
R47 VTAIL.n2 VTAIL.t1 54.1648
R48 VTAIL.n9 VTAIL.n8 51.0809
R49 VTAIL.n6 VTAIL.n5 51.0809
R50 VTAIL.n1 VTAIL.n0 51.0807
R51 VTAIL.n4 VTAIL.n3 51.0807
R52 VTAIL.n6 VTAIL.n4 20.7634
R53 VTAIL.n11 VTAIL.n10 19.3324
R54 VTAIL.n0 VTAIL.t4 3.08461
R55 VTAIL.n0 VTAIL.t9 3.08461
R56 VTAIL.n3 VTAIL.t11 3.08461
R57 VTAIL.n3 VTAIL.t2 3.08461
R58 VTAIL.n8 VTAIL.t10 3.08461
R59 VTAIL.n8 VTAIL.t0 3.08461
R60 VTAIL.n5 VTAIL.t7 3.08461
R61 VTAIL.n5 VTAIL.t6 3.08461
R62 VTAIL.n7 VTAIL.n6 1.43153
R63 VTAIL.n10 VTAIL.n9 1.43153
R64 VTAIL.n4 VTAIL.n2 1.43153
R65 VTAIL.n9 VTAIL.n7 1.18584
R66 VTAIL.n2 VTAIL.n1 1.18584
R67 VTAIL VTAIL.n11 1.01559
R68 VTAIL VTAIL.n1 0.416448
R69 B.n529 B.n528 585
R70 B.n202 B.n82 585
R71 B.n201 B.n200 585
R72 B.n199 B.n198 585
R73 B.n197 B.n196 585
R74 B.n195 B.n194 585
R75 B.n193 B.n192 585
R76 B.n191 B.n190 585
R77 B.n189 B.n188 585
R78 B.n187 B.n186 585
R79 B.n185 B.n184 585
R80 B.n183 B.n182 585
R81 B.n181 B.n180 585
R82 B.n179 B.n178 585
R83 B.n177 B.n176 585
R84 B.n175 B.n174 585
R85 B.n173 B.n172 585
R86 B.n171 B.n170 585
R87 B.n169 B.n168 585
R88 B.n167 B.n166 585
R89 B.n165 B.n164 585
R90 B.n163 B.n162 585
R91 B.n161 B.n160 585
R92 B.n159 B.n158 585
R93 B.n157 B.n156 585
R94 B.n154 B.n153 585
R95 B.n152 B.n151 585
R96 B.n150 B.n149 585
R97 B.n148 B.n147 585
R98 B.n146 B.n145 585
R99 B.n144 B.n143 585
R100 B.n142 B.n141 585
R101 B.n140 B.n139 585
R102 B.n138 B.n137 585
R103 B.n136 B.n135 585
R104 B.n133 B.n132 585
R105 B.n131 B.n130 585
R106 B.n129 B.n128 585
R107 B.n127 B.n126 585
R108 B.n125 B.n124 585
R109 B.n123 B.n122 585
R110 B.n121 B.n120 585
R111 B.n119 B.n118 585
R112 B.n117 B.n116 585
R113 B.n115 B.n114 585
R114 B.n113 B.n112 585
R115 B.n111 B.n110 585
R116 B.n109 B.n108 585
R117 B.n107 B.n106 585
R118 B.n105 B.n104 585
R119 B.n103 B.n102 585
R120 B.n101 B.n100 585
R121 B.n99 B.n98 585
R122 B.n97 B.n96 585
R123 B.n95 B.n94 585
R124 B.n93 B.n92 585
R125 B.n91 B.n90 585
R126 B.n89 B.n88 585
R127 B.n53 B.n52 585
R128 B.n534 B.n533 585
R129 B.n527 B.n83 585
R130 B.n83 B.n50 585
R131 B.n526 B.n49 585
R132 B.n538 B.n49 585
R133 B.n525 B.n48 585
R134 B.n539 B.n48 585
R135 B.n524 B.n47 585
R136 B.n540 B.n47 585
R137 B.n523 B.n522 585
R138 B.n522 B.n43 585
R139 B.n521 B.n42 585
R140 B.n546 B.n42 585
R141 B.n520 B.n41 585
R142 B.n547 B.n41 585
R143 B.n519 B.n40 585
R144 B.n548 B.n40 585
R145 B.n518 B.n517 585
R146 B.n517 B.n36 585
R147 B.n516 B.n35 585
R148 B.n554 B.n35 585
R149 B.n515 B.n34 585
R150 B.n555 B.n34 585
R151 B.n514 B.n33 585
R152 B.n556 B.n33 585
R153 B.n513 B.n512 585
R154 B.n512 B.n29 585
R155 B.n511 B.n28 585
R156 B.n562 B.n28 585
R157 B.n510 B.n27 585
R158 B.n563 B.n27 585
R159 B.n509 B.n26 585
R160 B.n564 B.n26 585
R161 B.n508 B.n507 585
R162 B.n507 B.n22 585
R163 B.n506 B.n21 585
R164 B.n570 B.n21 585
R165 B.n505 B.n20 585
R166 B.n571 B.n20 585
R167 B.n504 B.n19 585
R168 B.n572 B.n19 585
R169 B.n503 B.n502 585
R170 B.n502 B.n15 585
R171 B.n501 B.n14 585
R172 B.n578 B.n14 585
R173 B.n500 B.n13 585
R174 B.n579 B.n13 585
R175 B.n499 B.n12 585
R176 B.n580 B.n12 585
R177 B.n498 B.n497 585
R178 B.n497 B.n496 585
R179 B.n495 B.n494 585
R180 B.n495 B.n8 585
R181 B.n493 B.n7 585
R182 B.n587 B.n7 585
R183 B.n492 B.n6 585
R184 B.n588 B.n6 585
R185 B.n491 B.n5 585
R186 B.n589 B.n5 585
R187 B.n490 B.n489 585
R188 B.n489 B.n4 585
R189 B.n488 B.n203 585
R190 B.n488 B.n487 585
R191 B.n478 B.n204 585
R192 B.n205 B.n204 585
R193 B.n480 B.n479 585
R194 B.n481 B.n480 585
R195 B.n477 B.n210 585
R196 B.n210 B.n209 585
R197 B.n476 B.n475 585
R198 B.n475 B.n474 585
R199 B.n212 B.n211 585
R200 B.n213 B.n212 585
R201 B.n467 B.n466 585
R202 B.n468 B.n467 585
R203 B.n465 B.n217 585
R204 B.n221 B.n217 585
R205 B.n464 B.n463 585
R206 B.n463 B.n462 585
R207 B.n219 B.n218 585
R208 B.n220 B.n219 585
R209 B.n455 B.n454 585
R210 B.n456 B.n455 585
R211 B.n453 B.n226 585
R212 B.n226 B.n225 585
R213 B.n452 B.n451 585
R214 B.n451 B.n450 585
R215 B.n228 B.n227 585
R216 B.n229 B.n228 585
R217 B.n443 B.n442 585
R218 B.n444 B.n443 585
R219 B.n441 B.n234 585
R220 B.n234 B.n233 585
R221 B.n440 B.n439 585
R222 B.n439 B.n438 585
R223 B.n236 B.n235 585
R224 B.n237 B.n236 585
R225 B.n431 B.n430 585
R226 B.n432 B.n431 585
R227 B.n429 B.n242 585
R228 B.n242 B.n241 585
R229 B.n428 B.n427 585
R230 B.n427 B.n426 585
R231 B.n244 B.n243 585
R232 B.n245 B.n244 585
R233 B.n419 B.n418 585
R234 B.n420 B.n419 585
R235 B.n417 B.n250 585
R236 B.n250 B.n249 585
R237 B.n416 B.n415 585
R238 B.n415 B.n414 585
R239 B.n252 B.n251 585
R240 B.n253 B.n252 585
R241 B.n410 B.n409 585
R242 B.n256 B.n255 585
R243 B.n406 B.n405 585
R244 B.n407 B.n406 585
R245 B.n404 B.n286 585
R246 B.n403 B.n402 585
R247 B.n401 B.n400 585
R248 B.n399 B.n398 585
R249 B.n397 B.n396 585
R250 B.n395 B.n394 585
R251 B.n393 B.n392 585
R252 B.n391 B.n390 585
R253 B.n389 B.n388 585
R254 B.n387 B.n386 585
R255 B.n385 B.n384 585
R256 B.n383 B.n382 585
R257 B.n381 B.n380 585
R258 B.n379 B.n378 585
R259 B.n377 B.n376 585
R260 B.n375 B.n374 585
R261 B.n373 B.n372 585
R262 B.n371 B.n370 585
R263 B.n369 B.n368 585
R264 B.n367 B.n366 585
R265 B.n365 B.n364 585
R266 B.n363 B.n362 585
R267 B.n361 B.n360 585
R268 B.n359 B.n358 585
R269 B.n357 B.n356 585
R270 B.n355 B.n354 585
R271 B.n353 B.n352 585
R272 B.n351 B.n350 585
R273 B.n349 B.n348 585
R274 B.n347 B.n346 585
R275 B.n345 B.n344 585
R276 B.n343 B.n342 585
R277 B.n341 B.n340 585
R278 B.n339 B.n338 585
R279 B.n337 B.n336 585
R280 B.n335 B.n334 585
R281 B.n333 B.n332 585
R282 B.n331 B.n330 585
R283 B.n329 B.n328 585
R284 B.n327 B.n326 585
R285 B.n325 B.n324 585
R286 B.n323 B.n322 585
R287 B.n321 B.n320 585
R288 B.n319 B.n318 585
R289 B.n317 B.n316 585
R290 B.n315 B.n314 585
R291 B.n313 B.n312 585
R292 B.n311 B.n310 585
R293 B.n309 B.n308 585
R294 B.n307 B.n306 585
R295 B.n305 B.n304 585
R296 B.n303 B.n302 585
R297 B.n301 B.n300 585
R298 B.n299 B.n298 585
R299 B.n297 B.n296 585
R300 B.n295 B.n294 585
R301 B.n293 B.n285 585
R302 B.n407 B.n285 585
R303 B.n411 B.n254 585
R304 B.n254 B.n253 585
R305 B.n413 B.n412 585
R306 B.n414 B.n413 585
R307 B.n248 B.n247 585
R308 B.n249 B.n248 585
R309 B.n422 B.n421 585
R310 B.n421 B.n420 585
R311 B.n423 B.n246 585
R312 B.n246 B.n245 585
R313 B.n425 B.n424 585
R314 B.n426 B.n425 585
R315 B.n240 B.n239 585
R316 B.n241 B.n240 585
R317 B.n434 B.n433 585
R318 B.n433 B.n432 585
R319 B.n435 B.n238 585
R320 B.n238 B.n237 585
R321 B.n437 B.n436 585
R322 B.n438 B.n437 585
R323 B.n232 B.n231 585
R324 B.n233 B.n232 585
R325 B.n446 B.n445 585
R326 B.n445 B.n444 585
R327 B.n447 B.n230 585
R328 B.n230 B.n229 585
R329 B.n449 B.n448 585
R330 B.n450 B.n449 585
R331 B.n224 B.n223 585
R332 B.n225 B.n224 585
R333 B.n458 B.n457 585
R334 B.n457 B.n456 585
R335 B.n459 B.n222 585
R336 B.n222 B.n220 585
R337 B.n461 B.n460 585
R338 B.n462 B.n461 585
R339 B.n216 B.n215 585
R340 B.n221 B.n216 585
R341 B.n470 B.n469 585
R342 B.n469 B.n468 585
R343 B.n471 B.n214 585
R344 B.n214 B.n213 585
R345 B.n473 B.n472 585
R346 B.n474 B.n473 585
R347 B.n208 B.n207 585
R348 B.n209 B.n208 585
R349 B.n483 B.n482 585
R350 B.n482 B.n481 585
R351 B.n484 B.n206 585
R352 B.n206 B.n205 585
R353 B.n486 B.n485 585
R354 B.n487 B.n486 585
R355 B.n3 B.n0 585
R356 B.n4 B.n3 585
R357 B.n586 B.n1 585
R358 B.n587 B.n586 585
R359 B.n585 B.n584 585
R360 B.n585 B.n8 585
R361 B.n583 B.n9 585
R362 B.n496 B.n9 585
R363 B.n582 B.n581 585
R364 B.n581 B.n580 585
R365 B.n11 B.n10 585
R366 B.n579 B.n11 585
R367 B.n577 B.n576 585
R368 B.n578 B.n577 585
R369 B.n575 B.n16 585
R370 B.n16 B.n15 585
R371 B.n574 B.n573 585
R372 B.n573 B.n572 585
R373 B.n18 B.n17 585
R374 B.n571 B.n18 585
R375 B.n569 B.n568 585
R376 B.n570 B.n569 585
R377 B.n567 B.n23 585
R378 B.n23 B.n22 585
R379 B.n566 B.n565 585
R380 B.n565 B.n564 585
R381 B.n25 B.n24 585
R382 B.n563 B.n25 585
R383 B.n561 B.n560 585
R384 B.n562 B.n561 585
R385 B.n559 B.n30 585
R386 B.n30 B.n29 585
R387 B.n558 B.n557 585
R388 B.n557 B.n556 585
R389 B.n32 B.n31 585
R390 B.n555 B.n32 585
R391 B.n553 B.n552 585
R392 B.n554 B.n553 585
R393 B.n551 B.n37 585
R394 B.n37 B.n36 585
R395 B.n550 B.n549 585
R396 B.n549 B.n548 585
R397 B.n39 B.n38 585
R398 B.n547 B.n39 585
R399 B.n545 B.n544 585
R400 B.n546 B.n545 585
R401 B.n543 B.n44 585
R402 B.n44 B.n43 585
R403 B.n542 B.n541 585
R404 B.n541 B.n540 585
R405 B.n46 B.n45 585
R406 B.n539 B.n46 585
R407 B.n537 B.n536 585
R408 B.n538 B.n537 585
R409 B.n535 B.n51 585
R410 B.n51 B.n50 585
R411 B.n590 B.n589 585
R412 B.n588 B.n2 585
R413 B.n533 B.n51 521.33
R414 B.n529 B.n83 521.33
R415 B.n285 B.n252 521.33
R416 B.n409 B.n254 521.33
R417 B.n86 B.t15 321.079
R418 B.n84 B.t4 321.079
R419 B.n290 B.t8 321.079
R420 B.n287 B.t12 321.079
R421 B.n531 B.n530 256.663
R422 B.n531 B.n81 256.663
R423 B.n531 B.n80 256.663
R424 B.n531 B.n79 256.663
R425 B.n531 B.n78 256.663
R426 B.n531 B.n77 256.663
R427 B.n531 B.n76 256.663
R428 B.n531 B.n75 256.663
R429 B.n531 B.n74 256.663
R430 B.n531 B.n73 256.663
R431 B.n531 B.n72 256.663
R432 B.n531 B.n71 256.663
R433 B.n531 B.n70 256.663
R434 B.n531 B.n69 256.663
R435 B.n531 B.n68 256.663
R436 B.n531 B.n67 256.663
R437 B.n531 B.n66 256.663
R438 B.n531 B.n65 256.663
R439 B.n531 B.n64 256.663
R440 B.n531 B.n63 256.663
R441 B.n531 B.n62 256.663
R442 B.n531 B.n61 256.663
R443 B.n531 B.n60 256.663
R444 B.n531 B.n59 256.663
R445 B.n531 B.n58 256.663
R446 B.n531 B.n57 256.663
R447 B.n531 B.n56 256.663
R448 B.n531 B.n55 256.663
R449 B.n531 B.n54 256.663
R450 B.n532 B.n531 256.663
R451 B.n408 B.n407 256.663
R452 B.n407 B.n257 256.663
R453 B.n407 B.n258 256.663
R454 B.n407 B.n259 256.663
R455 B.n407 B.n260 256.663
R456 B.n407 B.n261 256.663
R457 B.n407 B.n262 256.663
R458 B.n407 B.n263 256.663
R459 B.n407 B.n264 256.663
R460 B.n407 B.n265 256.663
R461 B.n407 B.n266 256.663
R462 B.n407 B.n267 256.663
R463 B.n407 B.n268 256.663
R464 B.n407 B.n269 256.663
R465 B.n407 B.n270 256.663
R466 B.n407 B.n271 256.663
R467 B.n407 B.n272 256.663
R468 B.n407 B.n273 256.663
R469 B.n407 B.n274 256.663
R470 B.n407 B.n275 256.663
R471 B.n407 B.n276 256.663
R472 B.n407 B.n277 256.663
R473 B.n407 B.n278 256.663
R474 B.n407 B.n279 256.663
R475 B.n407 B.n280 256.663
R476 B.n407 B.n281 256.663
R477 B.n407 B.n282 256.663
R478 B.n407 B.n283 256.663
R479 B.n407 B.n284 256.663
R480 B.n592 B.n591 256.663
R481 B.n88 B.n53 163.367
R482 B.n92 B.n91 163.367
R483 B.n96 B.n95 163.367
R484 B.n100 B.n99 163.367
R485 B.n104 B.n103 163.367
R486 B.n108 B.n107 163.367
R487 B.n112 B.n111 163.367
R488 B.n116 B.n115 163.367
R489 B.n120 B.n119 163.367
R490 B.n124 B.n123 163.367
R491 B.n128 B.n127 163.367
R492 B.n132 B.n131 163.367
R493 B.n137 B.n136 163.367
R494 B.n141 B.n140 163.367
R495 B.n145 B.n144 163.367
R496 B.n149 B.n148 163.367
R497 B.n153 B.n152 163.367
R498 B.n158 B.n157 163.367
R499 B.n162 B.n161 163.367
R500 B.n166 B.n165 163.367
R501 B.n170 B.n169 163.367
R502 B.n174 B.n173 163.367
R503 B.n178 B.n177 163.367
R504 B.n182 B.n181 163.367
R505 B.n186 B.n185 163.367
R506 B.n190 B.n189 163.367
R507 B.n194 B.n193 163.367
R508 B.n198 B.n197 163.367
R509 B.n200 B.n82 163.367
R510 B.n415 B.n252 163.367
R511 B.n415 B.n250 163.367
R512 B.n419 B.n250 163.367
R513 B.n419 B.n244 163.367
R514 B.n427 B.n244 163.367
R515 B.n427 B.n242 163.367
R516 B.n431 B.n242 163.367
R517 B.n431 B.n236 163.367
R518 B.n439 B.n236 163.367
R519 B.n439 B.n234 163.367
R520 B.n443 B.n234 163.367
R521 B.n443 B.n228 163.367
R522 B.n451 B.n228 163.367
R523 B.n451 B.n226 163.367
R524 B.n455 B.n226 163.367
R525 B.n455 B.n219 163.367
R526 B.n463 B.n219 163.367
R527 B.n463 B.n217 163.367
R528 B.n467 B.n217 163.367
R529 B.n467 B.n212 163.367
R530 B.n475 B.n212 163.367
R531 B.n475 B.n210 163.367
R532 B.n480 B.n210 163.367
R533 B.n480 B.n204 163.367
R534 B.n488 B.n204 163.367
R535 B.n489 B.n488 163.367
R536 B.n489 B.n5 163.367
R537 B.n6 B.n5 163.367
R538 B.n7 B.n6 163.367
R539 B.n495 B.n7 163.367
R540 B.n497 B.n495 163.367
R541 B.n497 B.n12 163.367
R542 B.n13 B.n12 163.367
R543 B.n14 B.n13 163.367
R544 B.n502 B.n14 163.367
R545 B.n502 B.n19 163.367
R546 B.n20 B.n19 163.367
R547 B.n21 B.n20 163.367
R548 B.n507 B.n21 163.367
R549 B.n507 B.n26 163.367
R550 B.n27 B.n26 163.367
R551 B.n28 B.n27 163.367
R552 B.n512 B.n28 163.367
R553 B.n512 B.n33 163.367
R554 B.n34 B.n33 163.367
R555 B.n35 B.n34 163.367
R556 B.n517 B.n35 163.367
R557 B.n517 B.n40 163.367
R558 B.n41 B.n40 163.367
R559 B.n42 B.n41 163.367
R560 B.n522 B.n42 163.367
R561 B.n522 B.n47 163.367
R562 B.n48 B.n47 163.367
R563 B.n49 B.n48 163.367
R564 B.n83 B.n49 163.367
R565 B.n406 B.n256 163.367
R566 B.n406 B.n286 163.367
R567 B.n402 B.n401 163.367
R568 B.n398 B.n397 163.367
R569 B.n394 B.n393 163.367
R570 B.n390 B.n389 163.367
R571 B.n386 B.n385 163.367
R572 B.n382 B.n381 163.367
R573 B.n378 B.n377 163.367
R574 B.n374 B.n373 163.367
R575 B.n370 B.n369 163.367
R576 B.n366 B.n365 163.367
R577 B.n362 B.n361 163.367
R578 B.n358 B.n357 163.367
R579 B.n354 B.n353 163.367
R580 B.n350 B.n349 163.367
R581 B.n346 B.n345 163.367
R582 B.n342 B.n341 163.367
R583 B.n338 B.n337 163.367
R584 B.n334 B.n333 163.367
R585 B.n330 B.n329 163.367
R586 B.n326 B.n325 163.367
R587 B.n322 B.n321 163.367
R588 B.n318 B.n317 163.367
R589 B.n314 B.n313 163.367
R590 B.n310 B.n309 163.367
R591 B.n306 B.n305 163.367
R592 B.n302 B.n301 163.367
R593 B.n298 B.n297 163.367
R594 B.n294 B.n285 163.367
R595 B.n413 B.n254 163.367
R596 B.n413 B.n248 163.367
R597 B.n421 B.n248 163.367
R598 B.n421 B.n246 163.367
R599 B.n425 B.n246 163.367
R600 B.n425 B.n240 163.367
R601 B.n433 B.n240 163.367
R602 B.n433 B.n238 163.367
R603 B.n437 B.n238 163.367
R604 B.n437 B.n232 163.367
R605 B.n445 B.n232 163.367
R606 B.n445 B.n230 163.367
R607 B.n449 B.n230 163.367
R608 B.n449 B.n224 163.367
R609 B.n457 B.n224 163.367
R610 B.n457 B.n222 163.367
R611 B.n461 B.n222 163.367
R612 B.n461 B.n216 163.367
R613 B.n469 B.n216 163.367
R614 B.n469 B.n214 163.367
R615 B.n473 B.n214 163.367
R616 B.n473 B.n208 163.367
R617 B.n482 B.n208 163.367
R618 B.n482 B.n206 163.367
R619 B.n486 B.n206 163.367
R620 B.n486 B.n3 163.367
R621 B.n590 B.n3 163.367
R622 B.n586 B.n2 163.367
R623 B.n586 B.n585 163.367
R624 B.n585 B.n9 163.367
R625 B.n581 B.n9 163.367
R626 B.n581 B.n11 163.367
R627 B.n577 B.n11 163.367
R628 B.n577 B.n16 163.367
R629 B.n573 B.n16 163.367
R630 B.n573 B.n18 163.367
R631 B.n569 B.n18 163.367
R632 B.n569 B.n23 163.367
R633 B.n565 B.n23 163.367
R634 B.n565 B.n25 163.367
R635 B.n561 B.n25 163.367
R636 B.n561 B.n30 163.367
R637 B.n557 B.n30 163.367
R638 B.n557 B.n32 163.367
R639 B.n553 B.n32 163.367
R640 B.n553 B.n37 163.367
R641 B.n549 B.n37 163.367
R642 B.n549 B.n39 163.367
R643 B.n545 B.n39 163.367
R644 B.n545 B.n44 163.367
R645 B.n541 B.n44 163.367
R646 B.n541 B.n46 163.367
R647 B.n537 B.n46 163.367
R648 B.n537 B.n51 163.367
R649 B.n407 B.n253 125.097
R650 B.n531 B.n50 125.097
R651 B.n84 B.t6 107.24
R652 B.n290 B.t11 107.24
R653 B.n86 B.t16 107.233
R654 B.n287 B.t14 107.233
R655 B.n85 B.t7 75.0454
R656 B.n291 B.t10 75.0454
R657 B.n87 B.t17 75.0386
R658 B.n288 B.t13 75.0386
R659 B.n533 B.n532 71.676
R660 B.n88 B.n54 71.676
R661 B.n92 B.n55 71.676
R662 B.n96 B.n56 71.676
R663 B.n100 B.n57 71.676
R664 B.n104 B.n58 71.676
R665 B.n108 B.n59 71.676
R666 B.n112 B.n60 71.676
R667 B.n116 B.n61 71.676
R668 B.n120 B.n62 71.676
R669 B.n124 B.n63 71.676
R670 B.n128 B.n64 71.676
R671 B.n132 B.n65 71.676
R672 B.n137 B.n66 71.676
R673 B.n141 B.n67 71.676
R674 B.n145 B.n68 71.676
R675 B.n149 B.n69 71.676
R676 B.n153 B.n70 71.676
R677 B.n158 B.n71 71.676
R678 B.n162 B.n72 71.676
R679 B.n166 B.n73 71.676
R680 B.n170 B.n74 71.676
R681 B.n174 B.n75 71.676
R682 B.n178 B.n76 71.676
R683 B.n182 B.n77 71.676
R684 B.n186 B.n78 71.676
R685 B.n190 B.n79 71.676
R686 B.n194 B.n80 71.676
R687 B.n198 B.n81 71.676
R688 B.n530 B.n82 71.676
R689 B.n530 B.n529 71.676
R690 B.n200 B.n81 71.676
R691 B.n197 B.n80 71.676
R692 B.n193 B.n79 71.676
R693 B.n189 B.n78 71.676
R694 B.n185 B.n77 71.676
R695 B.n181 B.n76 71.676
R696 B.n177 B.n75 71.676
R697 B.n173 B.n74 71.676
R698 B.n169 B.n73 71.676
R699 B.n165 B.n72 71.676
R700 B.n161 B.n71 71.676
R701 B.n157 B.n70 71.676
R702 B.n152 B.n69 71.676
R703 B.n148 B.n68 71.676
R704 B.n144 B.n67 71.676
R705 B.n140 B.n66 71.676
R706 B.n136 B.n65 71.676
R707 B.n131 B.n64 71.676
R708 B.n127 B.n63 71.676
R709 B.n123 B.n62 71.676
R710 B.n119 B.n61 71.676
R711 B.n115 B.n60 71.676
R712 B.n111 B.n59 71.676
R713 B.n107 B.n58 71.676
R714 B.n103 B.n57 71.676
R715 B.n99 B.n56 71.676
R716 B.n95 B.n55 71.676
R717 B.n91 B.n54 71.676
R718 B.n532 B.n53 71.676
R719 B.n409 B.n408 71.676
R720 B.n286 B.n257 71.676
R721 B.n401 B.n258 71.676
R722 B.n397 B.n259 71.676
R723 B.n393 B.n260 71.676
R724 B.n389 B.n261 71.676
R725 B.n385 B.n262 71.676
R726 B.n381 B.n263 71.676
R727 B.n377 B.n264 71.676
R728 B.n373 B.n265 71.676
R729 B.n369 B.n266 71.676
R730 B.n365 B.n267 71.676
R731 B.n361 B.n268 71.676
R732 B.n357 B.n269 71.676
R733 B.n353 B.n270 71.676
R734 B.n349 B.n271 71.676
R735 B.n345 B.n272 71.676
R736 B.n341 B.n273 71.676
R737 B.n337 B.n274 71.676
R738 B.n333 B.n275 71.676
R739 B.n329 B.n276 71.676
R740 B.n325 B.n277 71.676
R741 B.n321 B.n278 71.676
R742 B.n317 B.n279 71.676
R743 B.n313 B.n280 71.676
R744 B.n309 B.n281 71.676
R745 B.n305 B.n282 71.676
R746 B.n301 B.n283 71.676
R747 B.n297 B.n284 71.676
R748 B.n408 B.n256 71.676
R749 B.n402 B.n257 71.676
R750 B.n398 B.n258 71.676
R751 B.n394 B.n259 71.676
R752 B.n390 B.n260 71.676
R753 B.n386 B.n261 71.676
R754 B.n382 B.n262 71.676
R755 B.n378 B.n263 71.676
R756 B.n374 B.n264 71.676
R757 B.n370 B.n265 71.676
R758 B.n366 B.n266 71.676
R759 B.n362 B.n267 71.676
R760 B.n358 B.n268 71.676
R761 B.n354 B.n269 71.676
R762 B.n350 B.n270 71.676
R763 B.n346 B.n271 71.676
R764 B.n342 B.n272 71.676
R765 B.n338 B.n273 71.676
R766 B.n334 B.n274 71.676
R767 B.n330 B.n275 71.676
R768 B.n326 B.n276 71.676
R769 B.n322 B.n277 71.676
R770 B.n318 B.n278 71.676
R771 B.n314 B.n279 71.676
R772 B.n310 B.n280 71.676
R773 B.n306 B.n281 71.676
R774 B.n302 B.n282 71.676
R775 B.n298 B.n283 71.676
R776 B.n294 B.n284 71.676
R777 B.n591 B.n590 71.676
R778 B.n591 B.n2 71.676
R779 B.n414 B.n253 63.9595
R780 B.n414 B.n249 63.9595
R781 B.n420 B.n249 63.9595
R782 B.n420 B.n245 63.9595
R783 B.n426 B.n245 63.9595
R784 B.n432 B.n241 63.9595
R785 B.n432 B.n237 63.9595
R786 B.n438 B.n237 63.9595
R787 B.n438 B.n233 63.9595
R788 B.n444 B.n233 63.9595
R789 B.n444 B.n229 63.9595
R790 B.n450 B.n229 63.9595
R791 B.n456 B.n225 63.9595
R792 B.n456 B.n220 63.9595
R793 B.n462 B.n220 63.9595
R794 B.n462 B.n221 63.9595
R795 B.n468 B.n213 63.9595
R796 B.n474 B.n213 63.9595
R797 B.n474 B.n209 63.9595
R798 B.n481 B.n209 63.9595
R799 B.n487 B.n205 63.9595
R800 B.n487 B.n4 63.9595
R801 B.n589 B.n4 63.9595
R802 B.n589 B.n588 63.9595
R803 B.n588 B.n587 63.9595
R804 B.n587 B.n8 63.9595
R805 B.n496 B.n8 63.9595
R806 B.n580 B.n579 63.9595
R807 B.n579 B.n578 63.9595
R808 B.n578 B.n15 63.9595
R809 B.n572 B.n15 63.9595
R810 B.n571 B.n570 63.9595
R811 B.n570 B.n22 63.9595
R812 B.n564 B.n22 63.9595
R813 B.n564 B.n563 63.9595
R814 B.n562 B.n29 63.9595
R815 B.n556 B.n29 63.9595
R816 B.n556 B.n555 63.9595
R817 B.n555 B.n554 63.9595
R818 B.n554 B.n36 63.9595
R819 B.n548 B.n36 63.9595
R820 B.n548 B.n547 63.9595
R821 B.n546 B.n43 63.9595
R822 B.n540 B.n43 63.9595
R823 B.n540 B.n539 63.9595
R824 B.n539 B.n538 63.9595
R825 B.n538 B.n50 63.9595
R826 B.n134 B.n87 59.5399
R827 B.n155 B.n85 59.5399
R828 B.n292 B.n291 59.5399
R829 B.n289 B.n288 59.5399
R830 B.n450 B.t19 44.2074
R831 B.t3 B.n562 44.2074
R832 B.n426 B.t9 38.564
R833 B.t5 B.n546 38.564
R834 B.n221 B.t2 36.6828
R835 B.t0 B.n571 36.6828
R836 B.t1 B.n205 34.8017
R837 B.n496 B.t18 34.8017
R838 B.n411 B.n410 33.8737
R839 B.n293 B.n251 33.8737
R840 B.n528 B.n527 33.8737
R841 B.n535 B.n534 33.8737
R842 B.n87 B.n86 32.1944
R843 B.n85 B.n84 32.1944
R844 B.n291 B.n290 32.1944
R845 B.n288 B.n287 32.1944
R846 B.n481 B.t1 29.1583
R847 B.n580 B.t18 29.1583
R848 B.n468 B.t2 27.2771
R849 B.n572 B.t0 27.2771
R850 B.t9 B.n241 25.396
R851 B.n547 B.t5 25.396
R852 B.t19 B.n225 19.7525
R853 B.n563 B.t3 19.7525
R854 B B.n592 18.0485
R855 B.n412 B.n411 10.6151
R856 B.n412 B.n247 10.6151
R857 B.n422 B.n247 10.6151
R858 B.n423 B.n422 10.6151
R859 B.n424 B.n423 10.6151
R860 B.n424 B.n239 10.6151
R861 B.n434 B.n239 10.6151
R862 B.n435 B.n434 10.6151
R863 B.n436 B.n435 10.6151
R864 B.n436 B.n231 10.6151
R865 B.n446 B.n231 10.6151
R866 B.n447 B.n446 10.6151
R867 B.n448 B.n447 10.6151
R868 B.n448 B.n223 10.6151
R869 B.n458 B.n223 10.6151
R870 B.n459 B.n458 10.6151
R871 B.n460 B.n459 10.6151
R872 B.n460 B.n215 10.6151
R873 B.n470 B.n215 10.6151
R874 B.n471 B.n470 10.6151
R875 B.n472 B.n471 10.6151
R876 B.n472 B.n207 10.6151
R877 B.n483 B.n207 10.6151
R878 B.n484 B.n483 10.6151
R879 B.n485 B.n484 10.6151
R880 B.n485 B.n0 10.6151
R881 B.n410 B.n255 10.6151
R882 B.n405 B.n255 10.6151
R883 B.n405 B.n404 10.6151
R884 B.n404 B.n403 10.6151
R885 B.n403 B.n400 10.6151
R886 B.n400 B.n399 10.6151
R887 B.n399 B.n396 10.6151
R888 B.n396 B.n395 10.6151
R889 B.n395 B.n392 10.6151
R890 B.n392 B.n391 10.6151
R891 B.n391 B.n388 10.6151
R892 B.n388 B.n387 10.6151
R893 B.n387 B.n384 10.6151
R894 B.n384 B.n383 10.6151
R895 B.n383 B.n380 10.6151
R896 B.n380 B.n379 10.6151
R897 B.n379 B.n376 10.6151
R898 B.n376 B.n375 10.6151
R899 B.n375 B.n372 10.6151
R900 B.n372 B.n371 10.6151
R901 B.n371 B.n368 10.6151
R902 B.n368 B.n367 10.6151
R903 B.n367 B.n364 10.6151
R904 B.n364 B.n363 10.6151
R905 B.n360 B.n359 10.6151
R906 B.n359 B.n356 10.6151
R907 B.n356 B.n355 10.6151
R908 B.n355 B.n352 10.6151
R909 B.n352 B.n351 10.6151
R910 B.n351 B.n348 10.6151
R911 B.n348 B.n347 10.6151
R912 B.n347 B.n344 10.6151
R913 B.n344 B.n343 10.6151
R914 B.n340 B.n339 10.6151
R915 B.n339 B.n336 10.6151
R916 B.n336 B.n335 10.6151
R917 B.n335 B.n332 10.6151
R918 B.n332 B.n331 10.6151
R919 B.n331 B.n328 10.6151
R920 B.n328 B.n327 10.6151
R921 B.n327 B.n324 10.6151
R922 B.n324 B.n323 10.6151
R923 B.n323 B.n320 10.6151
R924 B.n320 B.n319 10.6151
R925 B.n319 B.n316 10.6151
R926 B.n316 B.n315 10.6151
R927 B.n315 B.n312 10.6151
R928 B.n312 B.n311 10.6151
R929 B.n311 B.n308 10.6151
R930 B.n308 B.n307 10.6151
R931 B.n307 B.n304 10.6151
R932 B.n304 B.n303 10.6151
R933 B.n303 B.n300 10.6151
R934 B.n300 B.n299 10.6151
R935 B.n299 B.n296 10.6151
R936 B.n296 B.n295 10.6151
R937 B.n295 B.n293 10.6151
R938 B.n416 B.n251 10.6151
R939 B.n417 B.n416 10.6151
R940 B.n418 B.n417 10.6151
R941 B.n418 B.n243 10.6151
R942 B.n428 B.n243 10.6151
R943 B.n429 B.n428 10.6151
R944 B.n430 B.n429 10.6151
R945 B.n430 B.n235 10.6151
R946 B.n440 B.n235 10.6151
R947 B.n441 B.n440 10.6151
R948 B.n442 B.n441 10.6151
R949 B.n442 B.n227 10.6151
R950 B.n452 B.n227 10.6151
R951 B.n453 B.n452 10.6151
R952 B.n454 B.n453 10.6151
R953 B.n454 B.n218 10.6151
R954 B.n464 B.n218 10.6151
R955 B.n465 B.n464 10.6151
R956 B.n466 B.n465 10.6151
R957 B.n466 B.n211 10.6151
R958 B.n476 B.n211 10.6151
R959 B.n477 B.n476 10.6151
R960 B.n479 B.n477 10.6151
R961 B.n479 B.n478 10.6151
R962 B.n478 B.n203 10.6151
R963 B.n490 B.n203 10.6151
R964 B.n491 B.n490 10.6151
R965 B.n492 B.n491 10.6151
R966 B.n493 B.n492 10.6151
R967 B.n494 B.n493 10.6151
R968 B.n498 B.n494 10.6151
R969 B.n499 B.n498 10.6151
R970 B.n500 B.n499 10.6151
R971 B.n501 B.n500 10.6151
R972 B.n503 B.n501 10.6151
R973 B.n504 B.n503 10.6151
R974 B.n505 B.n504 10.6151
R975 B.n506 B.n505 10.6151
R976 B.n508 B.n506 10.6151
R977 B.n509 B.n508 10.6151
R978 B.n510 B.n509 10.6151
R979 B.n511 B.n510 10.6151
R980 B.n513 B.n511 10.6151
R981 B.n514 B.n513 10.6151
R982 B.n515 B.n514 10.6151
R983 B.n516 B.n515 10.6151
R984 B.n518 B.n516 10.6151
R985 B.n519 B.n518 10.6151
R986 B.n520 B.n519 10.6151
R987 B.n521 B.n520 10.6151
R988 B.n523 B.n521 10.6151
R989 B.n524 B.n523 10.6151
R990 B.n525 B.n524 10.6151
R991 B.n526 B.n525 10.6151
R992 B.n527 B.n526 10.6151
R993 B.n584 B.n1 10.6151
R994 B.n584 B.n583 10.6151
R995 B.n583 B.n582 10.6151
R996 B.n582 B.n10 10.6151
R997 B.n576 B.n10 10.6151
R998 B.n576 B.n575 10.6151
R999 B.n575 B.n574 10.6151
R1000 B.n574 B.n17 10.6151
R1001 B.n568 B.n17 10.6151
R1002 B.n568 B.n567 10.6151
R1003 B.n567 B.n566 10.6151
R1004 B.n566 B.n24 10.6151
R1005 B.n560 B.n24 10.6151
R1006 B.n560 B.n559 10.6151
R1007 B.n559 B.n558 10.6151
R1008 B.n558 B.n31 10.6151
R1009 B.n552 B.n31 10.6151
R1010 B.n552 B.n551 10.6151
R1011 B.n551 B.n550 10.6151
R1012 B.n550 B.n38 10.6151
R1013 B.n544 B.n38 10.6151
R1014 B.n544 B.n543 10.6151
R1015 B.n543 B.n542 10.6151
R1016 B.n542 B.n45 10.6151
R1017 B.n536 B.n45 10.6151
R1018 B.n536 B.n535 10.6151
R1019 B.n534 B.n52 10.6151
R1020 B.n89 B.n52 10.6151
R1021 B.n90 B.n89 10.6151
R1022 B.n93 B.n90 10.6151
R1023 B.n94 B.n93 10.6151
R1024 B.n97 B.n94 10.6151
R1025 B.n98 B.n97 10.6151
R1026 B.n101 B.n98 10.6151
R1027 B.n102 B.n101 10.6151
R1028 B.n105 B.n102 10.6151
R1029 B.n106 B.n105 10.6151
R1030 B.n109 B.n106 10.6151
R1031 B.n110 B.n109 10.6151
R1032 B.n113 B.n110 10.6151
R1033 B.n114 B.n113 10.6151
R1034 B.n117 B.n114 10.6151
R1035 B.n118 B.n117 10.6151
R1036 B.n121 B.n118 10.6151
R1037 B.n122 B.n121 10.6151
R1038 B.n125 B.n122 10.6151
R1039 B.n126 B.n125 10.6151
R1040 B.n129 B.n126 10.6151
R1041 B.n130 B.n129 10.6151
R1042 B.n133 B.n130 10.6151
R1043 B.n138 B.n135 10.6151
R1044 B.n139 B.n138 10.6151
R1045 B.n142 B.n139 10.6151
R1046 B.n143 B.n142 10.6151
R1047 B.n146 B.n143 10.6151
R1048 B.n147 B.n146 10.6151
R1049 B.n150 B.n147 10.6151
R1050 B.n151 B.n150 10.6151
R1051 B.n154 B.n151 10.6151
R1052 B.n159 B.n156 10.6151
R1053 B.n160 B.n159 10.6151
R1054 B.n163 B.n160 10.6151
R1055 B.n164 B.n163 10.6151
R1056 B.n167 B.n164 10.6151
R1057 B.n168 B.n167 10.6151
R1058 B.n171 B.n168 10.6151
R1059 B.n172 B.n171 10.6151
R1060 B.n175 B.n172 10.6151
R1061 B.n176 B.n175 10.6151
R1062 B.n179 B.n176 10.6151
R1063 B.n180 B.n179 10.6151
R1064 B.n183 B.n180 10.6151
R1065 B.n184 B.n183 10.6151
R1066 B.n187 B.n184 10.6151
R1067 B.n188 B.n187 10.6151
R1068 B.n191 B.n188 10.6151
R1069 B.n192 B.n191 10.6151
R1070 B.n195 B.n192 10.6151
R1071 B.n196 B.n195 10.6151
R1072 B.n199 B.n196 10.6151
R1073 B.n201 B.n199 10.6151
R1074 B.n202 B.n201 10.6151
R1075 B.n528 B.n202 10.6151
R1076 B.n363 B.n289 9.36635
R1077 B.n340 B.n292 9.36635
R1078 B.n134 B.n133 9.36635
R1079 B.n156 B.n155 9.36635
R1080 B.n592 B.n0 8.11757
R1081 B.n592 B.n1 8.11757
R1082 B.n360 B.n289 1.24928
R1083 B.n343 B.n292 1.24928
R1084 B.n135 B.n134 1.24928
R1085 B.n155 B.n154 1.24928
R1086 VP.n15 VP.n14 178.023
R1087 VP.n27 VP.n26 178.023
R1088 VP.n13 VP.n12 178.023
R1089 VP.n8 VP.n5 161.3
R1090 VP.n10 VP.n9 161.3
R1091 VP.n11 VP.n4 161.3
R1092 VP.n25 VP.n0 161.3
R1093 VP.n24 VP.n23 161.3
R1094 VP.n22 VP.n1 161.3
R1095 VP.n21 VP.n20 161.3
R1096 VP.n19 VP.n2 161.3
R1097 VP.n18 VP.n17 161.3
R1098 VP.n16 VP.n3 161.3
R1099 VP.n7 VP.t3 148.995
R1100 VP.n20 VP.t4 116.332
R1101 VP.n14 VP.t2 116.332
R1102 VP.n26 VP.t1 116.332
R1103 VP.n6 VP.t0 116.332
R1104 VP.n12 VP.t5 116.332
R1105 VP.n19 VP.n18 56.5617
R1106 VP.n24 VP.n1 56.5617
R1107 VP.n10 VP.n5 56.5617
R1108 VP.n7 VP.n6 41.7772
R1109 VP.n15 VP.n13 39.3187
R1110 VP.n18 VP.n3 24.5923
R1111 VP.n20 VP.n19 24.5923
R1112 VP.n20 VP.n1 24.5923
R1113 VP.n25 VP.n24 24.5923
R1114 VP.n11 VP.n10 24.5923
R1115 VP.n6 VP.n5 24.5923
R1116 VP.n8 VP.n7 17.9746
R1117 VP.n14 VP.n3 7.86989
R1118 VP.n26 VP.n25 7.86989
R1119 VP.n12 VP.n11 7.86989
R1120 VP.n9 VP.n8 0.189894
R1121 VP.n9 VP.n4 0.189894
R1122 VP.n13 VP.n4 0.189894
R1123 VP.n16 VP.n15 0.189894
R1124 VP.n17 VP.n16 0.189894
R1125 VP.n17 VP.n2 0.189894
R1126 VP.n21 VP.n2 0.189894
R1127 VP.n22 VP.n21 0.189894
R1128 VP.n23 VP.n22 0.189894
R1129 VP.n23 VP.n0 0.189894
R1130 VP.n27 VP.n0 0.189894
R1131 VP VP.n27 0.0516364
R1132 VDD1 VDD1.t2 71.9752
R1133 VDD1.n1 VDD1.t3 71.8616
R1134 VDD1.n1 VDD1.n0 68.0619
R1135 VDD1.n3 VDD1.n2 67.7595
R1136 VDD1.n3 VDD1.n1 35.1992
R1137 VDD1.n2 VDD1.t5 3.08461
R1138 VDD1.n2 VDD1.t0 3.08461
R1139 VDD1.n0 VDD1.t1 3.08461
R1140 VDD1.n0 VDD1.t4 3.08461
R1141 VDD1 VDD1.n3 0.300069
C0 VDD1 VDD2 0.942571f
C1 VP VN 4.65957f
C2 VP VTAIL 3.37679f
C3 VTAIL VN 3.3625f
C4 VDD1 VP 3.39047f
C5 VDD1 VN 0.1494f
C6 VP VDD2 0.350539f
C7 VDD2 VN 3.19167f
C8 VDD1 VTAIL 5.47528f
C9 VTAIL VDD2 5.51776f
C10 VDD2 B 3.982267f
C11 VDD1 B 4.239837f
C12 VTAIL B 4.589112f
C13 VN B 8.68979f
C14 VP B 7.187768f
C15 VDD1.t2 B 1.22128f
C16 VDD1.t3 B 1.22066f
C17 VDD1.t1 B 0.113701f
C18 VDD1.t4 B 0.113701f
C19 VDD1.n0 B 0.957695f
C20 VDD1.n1 B 1.88167f
C21 VDD1.t5 B 0.113701f
C22 VDD1.t0 B 0.113701f
C23 VDD1.n2 B 0.956278f
C24 VDD1.n3 B 1.78581f
C25 VP.n0 B 0.037567f
C26 VP.t1 B 0.852281f
C27 VP.n1 B 0.062925f
C28 VP.n2 B 0.037567f
C29 VP.t4 B 0.852281f
C30 VP.n3 B 0.046279f
C31 VP.n4 B 0.037567f
C32 VP.t5 B 0.852281f
C33 VP.n5 B 0.062925f
C34 VP.t3 B 0.953903f
C35 VP.t0 B 0.852281f
C36 VP.n6 B 0.416379f
C37 VP.n7 B 0.407209f
C38 VP.n8 B 0.231506f
C39 VP.n9 B 0.037567f
C40 VP.n10 B 0.046295f
C41 VP.n11 B 0.046279f
C42 VP.n12 B 0.396542f
C43 VP.n13 B 1.39204f
C44 VP.t2 B 0.852281f
C45 VP.n14 B 0.396542f
C46 VP.n15 B 1.42649f
C47 VP.n16 B 0.037567f
C48 VP.n17 B 0.037567f
C49 VP.n18 B 0.046295f
C50 VP.n19 B 0.062925f
C51 VP.n20 B 0.369317f
C52 VP.n21 B 0.037567f
C53 VP.n22 B 0.037567f
C54 VP.n23 B 0.037567f
C55 VP.n24 B 0.046295f
C56 VP.n25 B 0.046279f
C57 VP.n26 B 0.396542f
C58 VP.n27 B 0.035593f
C59 VTAIL.t4 B 0.129543f
C60 VTAIL.t9 B 0.129543f
C61 VTAIL.n0 B 1.02317f
C62 VTAIL.n1 B 0.371471f
C63 VTAIL.t1 B 1.30546f
C64 VTAIL.n2 B 0.525991f
C65 VTAIL.t11 B 0.129543f
C66 VTAIL.t2 B 0.129543f
C67 VTAIL.n3 B 1.02317f
C68 VTAIL.n4 B 1.39516f
C69 VTAIL.t7 B 0.129543f
C70 VTAIL.t6 B 0.129543f
C71 VTAIL.n5 B 1.02317f
C72 VTAIL.n6 B 1.39516f
C73 VTAIL.t5 B 1.30547f
C74 VTAIL.n7 B 0.525983f
C75 VTAIL.t10 B 0.129543f
C76 VTAIL.t0 B 0.129543f
C77 VTAIL.n8 B 1.02317f
C78 VTAIL.n9 B 0.454985f
C79 VTAIL.t3 B 1.30546f
C80 VTAIL.n10 B 1.34842f
C81 VTAIL.t8 B 1.30546f
C82 VTAIL.n11 B 1.3142f
C83 VDD2.t1 B 1.20444f
C84 VDD2.t0 B 0.112189f
C85 VDD2.t5 B 0.112189f
C86 VDD2.n0 B 0.944962f
C87 VDD2.n1 B 1.77825f
C88 VDD2.t3 B 1.20003f
C89 VDD2.n2 B 1.76562f
C90 VDD2.t2 B 0.112189f
C91 VDD2.t4 B 0.112189f
C92 VDD2.n3 B 0.94494f
C93 VN.n0 B 0.036745f
C94 VN.t1 B 0.833631f
C95 VN.n1 B 0.061548f
C96 VN.t5 B 0.933028f
C97 VN.t0 B 0.833631f
C98 VN.n2 B 0.407267f
C99 VN.n3 B 0.398298f
C100 VN.n4 B 0.22644f
C101 VN.n5 B 0.036745f
C102 VN.n6 B 0.045282f
C103 VN.n7 B 0.045266f
C104 VN.n8 B 0.387864f
C105 VN.n9 B 0.034814f
C106 VN.n10 B 0.036745f
C107 VN.t2 B 0.833631f
C108 VN.n11 B 0.061548f
C109 VN.t4 B 0.933028f
C110 VN.t3 B 0.833631f
C111 VN.n12 B 0.407267f
C112 VN.n13 B 0.398298f
C113 VN.n14 B 0.22644f
C114 VN.n15 B 0.036745f
C115 VN.n16 B 0.045282f
C116 VN.n17 B 0.045266f
C117 VN.n18 B 0.387864f
C118 VN.n19 B 1.38581f
.ends

