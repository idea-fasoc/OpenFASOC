* NGSPICE file created from diff_pair_sample_1447.ext - technology: sky130A

.subckt diff_pair_sample_1447 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t7 VP.t0 VDD1.t1 w_n1654_n2582# sky130_fd_pr__pfet_01v8 ad=3.1473 pd=16.92 as=1.33155 ps=8.4 w=8.07 l=0.81
X1 B.t11 B.t9 B.t10 w_n1654_n2582# sky130_fd_pr__pfet_01v8 ad=3.1473 pd=16.92 as=0 ps=0 w=8.07 l=0.81
X2 B.t8 B.t6 B.t7 w_n1654_n2582# sky130_fd_pr__pfet_01v8 ad=3.1473 pd=16.92 as=0 ps=0 w=8.07 l=0.81
X3 VDD1.t3 VP.t1 VTAIL.t6 w_n1654_n2582# sky130_fd_pr__pfet_01v8 ad=1.33155 pd=8.4 as=3.1473 ps=16.92 w=8.07 l=0.81
X4 B.t5 B.t3 B.t4 w_n1654_n2582# sky130_fd_pr__pfet_01v8 ad=3.1473 pd=16.92 as=0 ps=0 w=8.07 l=0.81
X5 VDD1.t2 VP.t2 VTAIL.t5 w_n1654_n2582# sky130_fd_pr__pfet_01v8 ad=1.33155 pd=8.4 as=3.1473 ps=16.92 w=8.07 l=0.81
X6 VDD2.t3 VN.t0 VTAIL.t3 w_n1654_n2582# sky130_fd_pr__pfet_01v8 ad=1.33155 pd=8.4 as=3.1473 ps=16.92 w=8.07 l=0.81
X7 VDD2.t2 VN.t1 VTAIL.t0 w_n1654_n2582# sky130_fd_pr__pfet_01v8 ad=1.33155 pd=8.4 as=3.1473 ps=16.92 w=8.07 l=0.81
X8 VTAIL.t1 VN.t2 VDD2.t1 w_n1654_n2582# sky130_fd_pr__pfet_01v8 ad=3.1473 pd=16.92 as=1.33155 ps=8.4 w=8.07 l=0.81
X9 VTAIL.t2 VN.t3 VDD2.t0 w_n1654_n2582# sky130_fd_pr__pfet_01v8 ad=3.1473 pd=16.92 as=1.33155 ps=8.4 w=8.07 l=0.81
X10 B.t2 B.t0 B.t1 w_n1654_n2582# sky130_fd_pr__pfet_01v8 ad=3.1473 pd=16.92 as=0 ps=0 w=8.07 l=0.81
X11 VTAIL.t4 VP.t3 VDD1.t0 w_n1654_n2582# sky130_fd_pr__pfet_01v8 ad=3.1473 pd=16.92 as=1.33155 ps=8.4 w=8.07 l=0.81
R0 VP.n1 VP.t0 309.899
R1 VP.n1 VP.t2 309.849
R2 VP.n3 VP.t3 288.902
R3 VP.n5 VP.t1 288.902
R4 VP.n6 VP.n5 161.3
R5 VP.n4 VP.n0 161.3
R6 VP.n3 VP.n2 161.3
R7 VP.n2 VP.n1 82.5106
R8 VP.n4 VP.n3 24.1005
R9 VP.n5 VP.n4 24.1005
R10 VP.n2 VP.n0 0.189894
R11 VP.n6 VP.n0 0.189894
R12 VP VP.n6 0.0516364
R13 VDD1 VDD1.n1 115.186
R14 VDD1 VDD1.n0 81.0997
R15 VDD1.n0 VDD1.t1 4.02838
R16 VDD1.n0 VDD1.t2 4.02838
R17 VDD1.n1 VDD1.t0 4.02838
R18 VDD1.n1 VDD1.t3 4.02838
R19 VTAIL.n346 VTAIL.n308 756.745
R20 VTAIL.n38 VTAIL.n0 756.745
R21 VTAIL.n82 VTAIL.n44 756.745
R22 VTAIL.n126 VTAIL.n88 756.745
R23 VTAIL.n302 VTAIL.n264 756.745
R24 VTAIL.n258 VTAIL.n220 756.745
R25 VTAIL.n214 VTAIL.n176 756.745
R26 VTAIL.n170 VTAIL.n132 756.745
R27 VTAIL.n323 VTAIL.n322 585
R28 VTAIL.n320 VTAIL.n319 585
R29 VTAIL.n329 VTAIL.n328 585
R30 VTAIL.n331 VTAIL.n330 585
R31 VTAIL.n316 VTAIL.n315 585
R32 VTAIL.n337 VTAIL.n336 585
R33 VTAIL.n339 VTAIL.n338 585
R34 VTAIL.n312 VTAIL.n311 585
R35 VTAIL.n345 VTAIL.n344 585
R36 VTAIL.n347 VTAIL.n346 585
R37 VTAIL.n15 VTAIL.n14 585
R38 VTAIL.n12 VTAIL.n11 585
R39 VTAIL.n21 VTAIL.n20 585
R40 VTAIL.n23 VTAIL.n22 585
R41 VTAIL.n8 VTAIL.n7 585
R42 VTAIL.n29 VTAIL.n28 585
R43 VTAIL.n31 VTAIL.n30 585
R44 VTAIL.n4 VTAIL.n3 585
R45 VTAIL.n37 VTAIL.n36 585
R46 VTAIL.n39 VTAIL.n38 585
R47 VTAIL.n59 VTAIL.n58 585
R48 VTAIL.n56 VTAIL.n55 585
R49 VTAIL.n65 VTAIL.n64 585
R50 VTAIL.n67 VTAIL.n66 585
R51 VTAIL.n52 VTAIL.n51 585
R52 VTAIL.n73 VTAIL.n72 585
R53 VTAIL.n75 VTAIL.n74 585
R54 VTAIL.n48 VTAIL.n47 585
R55 VTAIL.n81 VTAIL.n80 585
R56 VTAIL.n83 VTAIL.n82 585
R57 VTAIL.n103 VTAIL.n102 585
R58 VTAIL.n100 VTAIL.n99 585
R59 VTAIL.n109 VTAIL.n108 585
R60 VTAIL.n111 VTAIL.n110 585
R61 VTAIL.n96 VTAIL.n95 585
R62 VTAIL.n117 VTAIL.n116 585
R63 VTAIL.n119 VTAIL.n118 585
R64 VTAIL.n92 VTAIL.n91 585
R65 VTAIL.n125 VTAIL.n124 585
R66 VTAIL.n127 VTAIL.n126 585
R67 VTAIL.n303 VTAIL.n302 585
R68 VTAIL.n301 VTAIL.n300 585
R69 VTAIL.n268 VTAIL.n267 585
R70 VTAIL.n295 VTAIL.n294 585
R71 VTAIL.n293 VTAIL.n292 585
R72 VTAIL.n272 VTAIL.n271 585
R73 VTAIL.n287 VTAIL.n286 585
R74 VTAIL.n285 VTAIL.n284 585
R75 VTAIL.n276 VTAIL.n275 585
R76 VTAIL.n279 VTAIL.n278 585
R77 VTAIL.n259 VTAIL.n258 585
R78 VTAIL.n257 VTAIL.n256 585
R79 VTAIL.n224 VTAIL.n223 585
R80 VTAIL.n251 VTAIL.n250 585
R81 VTAIL.n249 VTAIL.n248 585
R82 VTAIL.n228 VTAIL.n227 585
R83 VTAIL.n243 VTAIL.n242 585
R84 VTAIL.n241 VTAIL.n240 585
R85 VTAIL.n232 VTAIL.n231 585
R86 VTAIL.n235 VTAIL.n234 585
R87 VTAIL.n215 VTAIL.n214 585
R88 VTAIL.n213 VTAIL.n212 585
R89 VTAIL.n180 VTAIL.n179 585
R90 VTAIL.n207 VTAIL.n206 585
R91 VTAIL.n205 VTAIL.n204 585
R92 VTAIL.n184 VTAIL.n183 585
R93 VTAIL.n199 VTAIL.n198 585
R94 VTAIL.n197 VTAIL.n196 585
R95 VTAIL.n188 VTAIL.n187 585
R96 VTAIL.n191 VTAIL.n190 585
R97 VTAIL.n171 VTAIL.n170 585
R98 VTAIL.n169 VTAIL.n168 585
R99 VTAIL.n136 VTAIL.n135 585
R100 VTAIL.n163 VTAIL.n162 585
R101 VTAIL.n161 VTAIL.n160 585
R102 VTAIL.n140 VTAIL.n139 585
R103 VTAIL.n155 VTAIL.n154 585
R104 VTAIL.n153 VTAIL.n152 585
R105 VTAIL.n144 VTAIL.n143 585
R106 VTAIL.n147 VTAIL.n146 585
R107 VTAIL.t0 VTAIL.n321 327.473
R108 VTAIL.t2 VTAIL.n13 327.473
R109 VTAIL.t6 VTAIL.n57 327.473
R110 VTAIL.t4 VTAIL.n101 327.473
R111 VTAIL.t5 VTAIL.n277 327.473
R112 VTAIL.t7 VTAIL.n233 327.473
R113 VTAIL.t3 VTAIL.n189 327.473
R114 VTAIL.t1 VTAIL.n145 327.473
R115 VTAIL.n322 VTAIL.n319 171.744
R116 VTAIL.n329 VTAIL.n319 171.744
R117 VTAIL.n330 VTAIL.n329 171.744
R118 VTAIL.n330 VTAIL.n315 171.744
R119 VTAIL.n337 VTAIL.n315 171.744
R120 VTAIL.n338 VTAIL.n337 171.744
R121 VTAIL.n338 VTAIL.n311 171.744
R122 VTAIL.n345 VTAIL.n311 171.744
R123 VTAIL.n346 VTAIL.n345 171.744
R124 VTAIL.n14 VTAIL.n11 171.744
R125 VTAIL.n21 VTAIL.n11 171.744
R126 VTAIL.n22 VTAIL.n21 171.744
R127 VTAIL.n22 VTAIL.n7 171.744
R128 VTAIL.n29 VTAIL.n7 171.744
R129 VTAIL.n30 VTAIL.n29 171.744
R130 VTAIL.n30 VTAIL.n3 171.744
R131 VTAIL.n37 VTAIL.n3 171.744
R132 VTAIL.n38 VTAIL.n37 171.744
R133 VTAIL.n58 VTAIL.n55 171.744
R134 VTAIL.n65 VTAIL.n55 171.744
R135 VTAIL.n66 VTAIL.n65 171.744
R136 VTAIL.n66 VTAIL.n51 171.744
R137 VTAIL.n73 VTAIL.n51 171.744
R138 VTAIL.n74 VTAIL.n73 171.744
R139 VTAIL.n74 VTAIL.n47 171.744
R140 VTAIL.n81 VTAIL.n47 171.744
R141 VTAIL.n82 VTAIL.n81 171.744
R142 VTAIL.n102 VTAIL.n99 171.744
R143 VTAIL.n109 VTAIL.n99 171.744
R144 VTAIL.n110 VTAIL.n109 171.744
R145 VTAIL.n110 VTAIL.n95 171.744
R146 VTAIL.n117 VTAIL.n95 171.744
R147 VTAIL.n118 VTAIL.n117 171.744
R148 VTAIL.n118 VTAIL.n91 171.744
R149 VTAIL.n125 VTAIL.n91 171.744
R150 VTAIL.n126 VTAIL.n125 171.744
R151 VTAIL.n302 VTAIL.n301 171.744
R152 VTAIL.n301 VTAIL.n267 171.744
R153 VTAIL.n294 VTAIL.n267 171.744
R154 VTAIL.n294 VTAIL.n293 171.744
R155 VTAIL.n293 VTAIL.n271 171.744
R156 VTAIL.n286 VTAIL.n271 171.744
R157 VTAIL.n286 VTAIL.n285 171.744
R158 VTAIL.n285 VTAIL.n275 171.744
R159 VTAIL.n278 VTAIL.n275 171.744
R160 VTAIL.n258 VTAIL.n257 171.744
R161 VTAIL.n257 VTAIL.n223 171.744
R162 VTAIL.n250 VTAIL.n223 171.744
R163 VTAIL.n250 VTAIL.n249 171.744
R164 VTAIL.n249 VTAIL.n227 171.744
R165 VTAIL.n242 VTAIL.n227 171.744
R166 VTAIL.n242 VTAIL.n241 171.744
R167 VTAIL.n241 VTAIL.n231 171.744
R168 VTAIL.n234 VTAIL.n231 171.744
R169 VTAIL.n214 VTAIL.n213 171.744
R170 VTAIL.n213 VTAIL.n179 171.744
R171 VTAIL.n206 VTAIL.n179 171.744
R172 VTAIL.n206 VTAIL.n205 171.744
R173 VTAIL.n205 VTAIL.n183 171.744
R174 VTAIL.n198 VTAIL.n183 171.744
R175 VTAIL.n198 VTAIL.n197 171.744
R176 VTAIL.n197 VTAIL.n187 171.744
R177 VTAIL.n190 VTAIL.n187 171.744
R178 VTAIL.n170 VTAIL.n169 171.744
R179 VTAIL.n169 VTAIL.n135 171.744
R180 VTAIL.n162 VTAIL.n135 171.744
R181 VTAIL.n162 VTAIL.n161 171.744
R182 VTAIL.n161 VTAIL.n139 171.744
R183 VTAIL.n154 VTAIL.n139 171.744
R184 VTAIL.n154 VTAIL.n153 171.744
R185 VTAIL.n153 VTAIL.n143 171.744
R186 VTAIL.n146 VTAIL.n143 171.744
R187 VTAIL.n322 VTAIL.t0 85.8723
R188 VTAIL.n14 VTAIL.t2 85.8723
R189 VTAIL.n58 VTAIL.t6 85.8723
R190 VTAIL.n102 VTAIL.t4 85.8723
R191 VTAIL.n278 VTAIL.t5 85.8723
R192 VTAIL.n234 VTAIL.t7 85.8723
R193 VTAIL.n190 VTAIL.t3 85.8723
R194 VTAIL.n146 VTAIL.t1 85.8723
R195 VTAIL.n351 VTAIL.n350 30.4399
R196 VTAIL.n43 VTAIL.n42 30.4399
R197 VTAIL.n87 VTAIL.n86 30.4399
R198 VTAIL.n131 VTAIL.n130 30.4399
R199 VTAIL.n307 VTAIL.n306 30.4399
R200 VTAIL.n263 VTAIL.n262 30.4399
R201 VTAIL.n219 VTAIL.n218 30.4399
R202 VTAIL.n175 VTAIL.n174 30.4399
R203 VTAIL.n351 VTAIL.n307 20.3065
R204 VTAIL.n175 VTAIL.n131 20.3065
R205 VTAIL.n323 VTAIL.n321 16.3894
R206 VTAIL.n15 VTAIL.n13 16.3894
R207 VTAIL.n59 VTAIL.n57 16.3894
R208 VTAIL.n103 VTAIL.n101 16.3894
R209 VTAIL.n279 VTAIL.n277 16.3894
R210 VTAIL.n235 VTAIL.n233 16.3894
R211 VTAIL.n191 VTAIL.n189 16.3894
R212 VTAIL.n147 VTAIL.n145 16.3894
R213 VTAIL.n324 VTAIL.n320 12.8005
R214 VTAIL.n16 VTAIL.n12 12.8005
R215 VTAIL.n60 VTAIL.n56 12.8005
R216 VTAIL.n104 VTAIL.n100 12.8005
R217 VTAIL.n280 VTAIL.n276 12.8005
R218 VTAIL.n236 VTAIL.n232 12.8005
R219 VTAIL.n192 VTAIL.n188 12.8005
R220 VTAIL.n148 VTAIL.n144 12.8005
R221 VTAIL.n328 VTAIL.n327 12.0247
R222 VTAIL.n20 VTAIL.n19 12.0247
R223 VTAIL.n64 VTAIL.n63 12.0247
R224 VTAIL.n108 VTAIL.n107 12.0247
R225 VTAIL.n284 VTAIL.n283 12.0247
R226 VTAIL.n240 VTAIL.n239 12.0247
R227 VTAIL.n196 VTAIL.n195 12.0247
R228 VTAIL.n152 VTAIL.n151 12.0247
R229 VTAIL.n331 VTAIL.n318 11.249
R230 VTAIL.n23 VTAIL.n10 11.249
R231 VTAIL.n67 VTAIL.n54 11.249
R232 VTAIL.n111 VTAIL.n98 11.249
R233 VTAIL.n287 VTAIL.n274 11.249
R234 VTAIL.n243 VTAIL.n230 11.249
R235 VTAIL.n199 VTAIL.n186 11.249
R236 VTAIL.n155 VTAIL.n142 11.249
R237 VTAIL.n332 VTAIL.n316 10.4732
R238 VTAIL.n24 VTAIL.n8 10.4732
R239 VTAIL.n68 VTAIL.n52 10.4732
R240 VTAIL.n112 VTAIL.n96 10.4732
R241 VTAIL.n288 VTAIL.n272 10.4732
R242 VTAIL.n244 VTAIL.n228 10.4732
R243 VTAIL.n200 VTAIL.n184 10.4732
R244 VTAIL.n156 VTAIL.n140 10.4732
R245 VTAIL.n336 VTAIL.n335 9.69747
R246 VTAIL.n28 VTAIL.n27 9.69747
R247 VTAIL.n72 VTAIL.n71 9.69747
R248 VTAIL.n116 VTAIL.n115 9.69747
R249 VTAIL.n292 VTAIL.n291 9.69747
R250 VTAIL.n248 VTAIL.n247 9.69747
R251 VTAIL.n204 VTAIL.n203 9.69747
R252 VTAIL.n160 VTAIL.n159 9.69747
R253 VTAIL.n350 VTAIL.n349 9.45567
R254 VTAIL.n42 VTAIL.n41 9.45567
R255 VTAIL.n86 VTAIL.n85 9.45567
R256 VTAIL.n130 VTAIL.n129 9.45567
R257 VTAIL.n306 VTAIL.n305 9.45567
R258 VTAIL.n262 VTAIL.n261 9.45567
R259 VTAIL.n218 VTAIL.n217 9.45567
R260 VTAIL.n174 VTAIL.n173 9.45567
R261 VTAIL.n310 VTAIL.n309 9.3005
R262 VTAIL.n349 VTAIL.n348 9.3005
R263 VTAIL.n341 VTAIL.n340 9.3005
R264 VTAIL.n314 VTAIL.n313 9.3005
R265 VTAIL.n335 VTAIL.n334 9.3005
R266 VTAIL.n333 VTAIL.n332 9.3005
R267 VTAIL.n318 VTAIL.n317 9.3005
R268 VTAIL.n327 VTAIL.n326 9.3005
R269 VTAIL.n325 VTAIL.n324 9.3005
R270 VTAIL.n343 VTAIL.n342 9.3005
R271 VTAIL.n2 VTAIL.n1 9.3005
R272 VTAIL.n41 VTAIL.n40 9.3005
R273 VTAIL.n33 VTAIL.n32 9.3005
R274 VTAIL.n6 VTAIL.n5 9.3005
R275 VTAIL.n27 VTAIL.n26 9.3005
R276 VTAIL.n25 VTAIL.n24 9.3005
R277 VTAIL.n10 VTAIL.n9 9.3005
R278 VTAIL.n19 VTAIL.n18 9.3005
R279 VTAIL.n17 VTAIL.n16 9.3005
R280 VTAIL.n35 VTAIL.n34 9.3005
R281 VTAIL.n46 VTAIL.n45 9.3005
R282 VTAIL.n85 VTAIL.n84 9.3005
R283 VTAIL.n77 VTAIL.n76 9.3005
R284 VTAIL.n50 VTAIL.n49 9.3005
R285 VTAIL.n71 VTAIL.n70 9.3005
R286 VTAIL.n69 VTAIL.n68 9.3005
R287 VTAIL.n54 VTAIL.n53 9.3005
R288 VTAIL.n63 VTAIL.n62 9.3005
R289 VTAIL.n61 VTAIL.n60 9.3005
R290 VTAIL.n79 VTAIL.n78 9.3005
R291 VTAIL.n90 VTAIL.n89 9.3005
R292 VTAIL.n129 VTAIL.n128 9.3005
R293 VTAIL.n121 VTAIL.n120 9.3005
R294 VTAIL.n94 VTAIL.n93 9.3005
R295 VTAIL.n115 VTAIL.n114 9.3005
R296 VTAIL.n113 VTAIL.n112 9.3005
R297 VTAIL.n98 VTAIL.n97 9.3005
R298 VTAIL.n107 VTAIL.n106 9.3005
R299 VTAIL.n105 VTAIL.n104 9.3005
R300 VTAIL.n123 VTAIL.n122 9.3005
R301 VTAIL.n266 VTAIL.n265 9.3005
R302 VTAIL.n299 VTAIL.n298 9.3005
R303 VTAIL.n297 VTAIL.n296 9.3005
R304 VTAIL.n270 VTAIL.n269 9.3005
R305 VTAIL.n291 VTAIL.n290 9.3005
R306 VTAIL.n289 VTAIL.n288 9.3005
R307 VTAIL.n274 VTAIL.n273 9.3005
R308 VTAIL.n283 VTAIL.n282 9.3005
R309 VTAIL.n281 VTAIL.n280 9.3005
R310 VTAIL.n305 VTAIL.n304 9.3005
R311 VTAIL.n261 VTAIL.n260 9.3005
R312 VTAIL.n222 VTAIL.n221 9.3005
R313 VTAIL.n255 VTAIL.n254 9.3005
R314 VTAIL.n253 VTAIL.n252 9.3005
R315 VTAIL.n226 VTAIL.n225 9.3005
R316 VTAIL.n247 VTAIL.n246 9.3005
R317 VTAIL.n245 VTAIL.n244 9.3005
R318 VTAIL.n230 VTAIL.n229 9.3005
R319 VTAIL.n239 VTAIL.n238 9.3005
R320 VTAIL.n237 VTAIL.n236 9.3005
R321 VTAIL.n217 VTAIL.n216 9.3005
R322 VTAIL.n178 VTAIL.n177 9.3005
R323 VTAIL.n211 VTAIL.n210 9.3005
R324 VTAIL.n209 VTAIL.n208 9.3005
R325 VTAIL.n182 VTAIL.n181 9.3005
R326 VTAIL.n203 VTAIL.n202 9.3005
R327 VTAIL.n201 VTAIL.n200 9.3005
R328 VTAIL.n186 VTAIL.n185 9.3005
R329 VTAIL.n195 VTAIL.n194 9.3005
R330 VTAIL.n193 VTAIL.n192 9.3005
R331 VTAIL.n173 VTAIL.n172 9.3005
R332 VTAIL.n134 VTAIL.n133 9.3005
R333 VTAIL.n167 VTAIL.n166 9.3005
R334 VTAIL.n165 VTAIL.n164 9.3005
R335 VTAIL.n138 VTAIL.n137 9.3005
R336 VTAIL.n159 VTAIL.n158 9.3005
R337 VTAIL.n157 VTAIL.n156 9.3005
R338 VTAIL.n142 VTAIL.n141 9.3005
R339 VTAIL.n151 VTAIL.n150 9.3005
R340 VTAIL.n149 VTAIL.n148 9.3005
R341 VTAIL.n339 VTAIL.n314 8.92171
R342 VTAIL.n31 VTAIL.n6 8.92171
R343 VTAIL.n75 VTAIL.n50 8.92171
R344 VTAIL.n119 VTAIL.n94 8.92171
R345 VTAIL.n295 VTAIL.n270 8.92171
R346 VTAIL.n251 VTAIL.n226 8.92171
R347 VTAIL.n207 VTAIL.n182 8.92171
R348 VTAIL.n163 VTAIL.n138 8.92171
R349 VTAIL.n340 VTAIL.n312 8.14595
R350 VTAIL.n350 VTAIL.n308 8.14595
R351 VTAIL.n32 VTAIL.n4 8.14595
R352 VTAIL.n42 VTAIL.n0 8.14595
R353 VTAIL.n76 VTAIL.n48 8.14595
R354 VTAIL.n86 VTAIL.n44 8.14595
R355 VTAIL.n120 VTAIL.n92 8.14595
R356 VTAIL.n130 VTAIL.n88 8.14595
R357 VTAIL.n306 VTAIL.n264 8.14595
R358 VTAIL.n296 VTAIL.n268 8.14595
R359 VTAIL.n262 VTAIL.n220 8.14595
R360 VTAIL.n252 VTAIL.n224 8.14595
R361 VTAIL.n218 VTAIL.n176 8.14595
R362 VTAIL.n208 VTAIL.n180 8.14595
R363 VTAIL.n174 VTAIL.n132 8.14595
R364 VTAIL.n164 VTAIL.n136 8.14595
R365 VTAIL.n344 VTAIL.n343 7.3702
R366 VTAIL.n348 VTAIL.n347 7.3702
R367 VTAIL.n36 VTAIL.n35 7.3702
R368 VTAIL.n40 VTAIL.n39 7.3702
R369 VTAIL.n80 VTAIL.n79 7.3702
R370 VTAIL.n84 VTAIL.n83 7.3702
R371 VTAIL.n124 VTAIL.n123 7.3702
R372 VTAIL.n128 VTAIL.n127 7.3702
R373 VTAIL.n304 VTAIL.n303 7.3702
R374 VTAIL.n300 VTAIL.n299 7.3702
R375 VTAIL.n260 VTAIL.n259 7.3702
R376 VTAIL.n256 VTAIL.n255 7.3702
R377 VTAIL.n216 VTAIL.n215 7.3702
R378 VTAIL.n212 VTAIL.n211 7.3702
R379 VTAIL.n172 VTAIL.n171 7.3702
R380 VTAIL.n168 VTAIL.n167 7.3702
R381 VTAIL.n344 VTAIL.n310 6.59444
R382 VTAIL.n347 VTAIL.n310 6.59444
R383 VTAIL.n36 VTAIL.n2 6.59444
R384 VTAIL.n39 VTAIL.n2 6.59444
R385 VTAIL.n80 VTAIL.n46 6.59444
R386 VTAIL.n83 VTAIL.n46 6.59444
R387 VTAIL.n124 VTAIL.n90 6.59444
R388 VTAIL.n127 VTAIL.n90 6.59444
R389 VTAIL.n303 VTAIL.n266 6.59444
R390 VTAIL.n300 VTAIL.n266 6.59444
R391 VTAIL.n259 VTAIL.n222 6.59444
R392 VTAIL.n256 VTAIL.n222 6.59444
R393 VTAIL.n215 VTAIL.n178 6.59444
R394 VTAIL.n212 VTAIL.n178 6.59444
R395 VTAIL.n171 VTAIL.n134 6.59444
R396 VTAIL.n168 VTAIL.n134 6.59444
R397 VTAIL.n343 VTAIL.n312 5.81868
R398 VTAIL.n348 VTAIL.n308 5.81868
R399 VTAIL.n35 VTAIL.n4 5.81868
R400 VTAIL.n40 VTAIL.n0 5.81868
R401 VTAIL.n79 VTAIL.n48 5.81868
R402 VTAIL.n84 VTAIL.n44 5.81868
R403 VTAIL.n123 VTAIL.n92 5.81868
R404 VTAIL.n128 VTAIL.n88 5.81868
R405 VTAIL.n304 VTAIL.n264 5.81868
R406 VTAIL.n299 VTAIL.n268 5.81868
R407 VTAIL.n260 VTAIL.n220 5.81868
R408 VTAIL.n255 VTAIL.n224 5.81868
R409 VTAIL.n216 VTAIL.n176 5.81868
R410 VTAIL.n211 VTAIL.n180 5.81868
R411 VTAIL.n172 VTAIL.n132 5.81868
R412 VTAIL.n167 VTAIL.n136 5.81868
R413 VTAIL.n340 VTAIL.n339 5.04292
R414 VTAIL.n32 VTAIL.n31 5.04292
R415 VTAIL.n76 VTAIL.n75 5.04292
R416 VTAIL.n120 VTAIL.n119 5.04292
R417 VTAIL.n296 VTAIL.n295 5.04292
R418 VTAIL.n252 VTAIL.n251 5.04292
R419 VTAIL.n208 VTAIL.n207 5.04292
R420 VTAIL.n164 VTAIL.n163 5.04292
R421 VTAIL.n336 VTAIL.n314 4.26717
R422 VTAIL.n28 VTAIL.n6 4.26717
R423 VTAIL.n72 VTAIL.n50 4.26717
R424 VTAIL.n116 VTAIL.n94 4.26717
R425 VTAIL.n292 VTAIL.n270 4.26717
R426 VTAIL.n248 VTAIL.n226 4.26717
R427 VTAIL.n204 VTAIL.n182 4.26717
R428 VTAIL.n160 VTAIL.n138 4.26717
R429 VTAIL.n325 VTAIL.n321 3.70995
R430 VTAIL.n17 VTAIL.n13 3.70995
R431 VTAIL.n61 VTAIL.n57 3.70995
R432 VTAIL.n105 VTAIL.n101 3.70995
R433 VTAIL.n237 VTAIL.n233 3.70995
R434 VTAIL.n193 VTAIL.n189 3.70995
R435 VTAIL.n149 VTAIL.n145 3.70995
R436 VTAIL.n281 VTAIL.n277 3.70995
R437 VTAIL.n335 VTAIL.n316 3.49141
R438 VTAIL.n27 VTAIL.n8 3.49141
R439 VTAIL.n71 VTAIL.n52 3.49141
R440 VTAIL.n115 VTAIL.n96 3.49141
R441 VTAIL.n291 VTAIL.n272 3.49141
R442 VTAIL.n247 VTAIL.n228 3.49141
R443 VTAIL.n203 VTAIL.n184 3.49141
R444 VTAIL.n159 VTAIL.n140 3.49141
R445 VTAIL.n332 VTAIL.n331 2.71565
R446 VTAIL.n24 VTAIL.n23 2.71565
R447 VTAIL.n68 VTAIL.n67 2.71565
R448 VTAIL.n112 VTAIL.n111 2.71565
R449 VTAIL.n288 VTAIL.n287 2.71565
R450 VTAIL.n244 VTAIL.n243 2.71565
R451 VTAIL.n200 VTAIL.n199 2.71565
R452 VTAIL.n156 VTAIL.n155 2.71565
R453 VTAIL.n328 VTAIL.n318 1.93989
R454 VTAIL.n20 VTAIL.n10 1.93989
R455 VTAIL.n64 VTAIL.n54 1.93989
R456 VTAIL.n108 VTAIL.n98 1.93989
R457 VTAIL.n284 VTAIL.n274 1.93989
R458 VTAIL.n240 VTAIL.n230 1.93989
R459 VTAIL.n196 VTAIL.n186 1.93989
R460 VTAIL.n152 VTAIL.n142 1.93989
R461 VTAIL.n327 VTAIL.n320 1.16414
R462 VTAIL.n19 VTAIL.n12 1.16414
R463 VTAIL.n63 VTAIL.n56 1.16414
R464 VTAIL.n107 VTAIL.n100 1.16414
R465 VTAIL.n283 VTAIL.n276 1.16414
R466 VTAIL.n239 VTAIL.n232 1.16414
R467 VTAIL.n195 VTAIL.n188 1.16414
R468 VTAIL.n151 VTAIL.n144 1.16414
R469 VTAIL.n219 VTAIL.n175 0.983259
R470 VTAIL.n307 VTAIL.n263 0.983259
R471 VTAIL.n131 VTAIL.n87 0.983259
R472 VTAIL VTAIL.n43 0.550069
R473 VTAIL.n263 VTAIL.n219 0.470328
R474 VTAIL.n87 VTAIL.n43 0.470328
R475 VTAIL VTAIL.n351 0.43369
R476 VTAIL.n324 VTAIL.n323 0.388379
R477 VTAIL.n16 VTAIL.n15 0.388379
R478 VTAIL.n60 VTAIL.n59 0.388379
R479 VTAIL.n104 VTAIL.n103 0.388379
R480 VTAIL.n280 VTAIL.n279 0.388379
R481 VTAIL.n236 VTAIL.n235 0.388379
R482 VTAIL.n192 VTAIL.n191 0.388379
R483 VTAIL.n148 VTAIL.n147 0.388379
R484 VTAIL.n326 VTAIL.n325 0.155672
R485 VTAIL.n326 VTAIL.n317 0.155672
R486 VTAIL.n333 VTAIL.n317 0.155672
R487 VTAIL.n334 VTAIL.n333 0.155672
R488 VTAIL.n334 VTAIL.n313 0.155672
R489 VTAIL.n341 VTAIL.n313 0.155672
R490 VTAIL.n342 VTAIL.n341 0.155672
R491 VTAIL.n342 VTAIL.n309 0.155672
R492 VTAIL.n349 VTAIL.n309 0.155672
R493 VTAIL.n18 VTAIL.n17 0.155672
R494 VTAIL.n18 VTAIL.n9 0.155672
R495 VTAIL.n25 VTAIL.n9 0.155672
R496 VTAIL.n26 VTAIL.n25 0.155672
R497 VTAIL.n26 VTAIL.n5 0.155672
R498 VTAIL.n33 VTAIL.n5 0.155672
R499 VTAIL.n34 VTAIL.n33 0.155672
R500 VTAIL.n34 VTAIL.n1 0.155672
R501 VTAIL.n41 VTAIL.n1 0.155672
R502 VTAIL.n62 VTAIL.n61 0.155672
R503 VTAIL.n62 VTAIL.n53 0.155672
R504 VTAIL.n69 VTAIL.n53 0.155672
R505 VTAIL.n70 VTAIL.n69 0.155672
R506 VTAIL.n70 VTAIL.n49 0.155672
R507 VTAIL.n77 VTAIL.n49 0.155672
R508 VTAIL.n78 VTAIL.n77 0.155672
R509 VTAIL.n78 VTAIL.n45 0.155672
R510 VTAIL.n85 VTAIL.n45 0.155672
R511 VTAIL.n106 VTAIL.n105 0.155672
R512 VTAIL.n106 VTAIL.n97 0.155672
R513 VTAIL.n113 VTAIL.n97 0.155672
R514 VTAIL.n114 VTAIL.n113 0.155672
R515 VTAIL.n114 VTAIL.n93 0.155672
R516 VTAIL.n121 VTAIL.n93 0.155672
R517 VTAIL.n122 VTAIL.n121 0.155672
R518 VTAIL.n122 VTAIL.n89 0.155672
R519 VTAIL.n129 VTAIL.n89 0.155672
R520 VTAIL.n305 VTAIL.n265 0.155672
R521 VTAIL.n298 VTAIL.n265 0.155672
R522 VTAIL.n298 VTAIL.n297 0.155672
R523 VTAIL.n297 VTAIL.n269 0.155672
R524 VTAIL.n290 VTAIL.n269 0.155672
R525 VTAIL.n290 VTAIL.n289 0.155672
R526 VTAIL.n289 VTAIL.n273 0.155672
R527 VTAIL.n282 VTAIL.n273 0.155672
R528 VTAIL.n282 VTAIL.n281 0.155672
R529 VTAIL.n261 VTAIL.n221 0.155672
R530 VTAIL.n254 VTAIL.n221 0.155672
R531 VTAIL.n254 VTAIL.n253 0.155672
R532 VTAIL.n253 VTAIL.n225 0.155672
R533 VTAIL.n246 VTAIL.n225 0.155672
R534 VTAIL.n246 VTAIL.n245 0.155672
R535 VTAIL.n245 VTAIL.n229 0.155672
R536 VTAIL.n238 VTAIL.n229 0.155672
R537 VTAIL.n238 VTAIL.n237 0.155672
R538 VTAIL.n217 VTAIL.n177 0.155672
R539 VTAIL.n210 VTAIL.n177 0.155672
R540 VTAIL.n210 VTAIL.n209 0.155672
R541 VTAIL.n209 VTAIL.n181 0.155672
R542 VTAIL.n202 VTAIL.n181 0.155672
R543 VTAIL.n202 VTAIL.n201 0.155672
R544 VTAIL.n201 VTAIL.n185 0.155672
R545 VTAIL.n194 VTAIL.n185 0.155672
R546 VTAIL.n194 VTAIL.n193 0.155672
R547 VTAIL.n173 VTAIL.n133 0.155672
R548 VTAIL.n166 VTAIL.n133 0.155672
R549 VTAIL.n166 VTAIL.n165 0.155672
R550 VTAIL.n165 VTAIL.n137 0.155672
R551 VTAIL.n158 VTAIL.n137 0.155672
R552 VTAIL.n158 VTAIL.n157 0.155672
R553 VTAIL.n157 VTAIL.n141 0.155672
R554 VTAIL.n150 VTAIL.n141 0.155672
R555 VTAIL.n150 VTAIL.n149 0.155672
R556 B.n305 B.n50 585
R557 B.n307 B.n306 585
R558 B.n308 B.n49 585
R559 B.n310 B.n309 585
R560 B.n311 B.n48 585
R561 B.n313 B.n312 585
R562 B.n314 B.n47 585
R563 B.n316 B.n315 585
R564 B.n317 B.n46 585
R565 B.n319 B.n318 585
R566 B.n320 B.n45 585
R567 B.n322 B.n321 585
R568 B.n323 B.n44 585
R569 B.n325 B.n324 585
R570 B.n326 B.n43 585
R571 B.n328 B.n327 585
R572 B.n329 B.n42 585
R573 B.n331 B.n330 585
R574 B.n332 B.n41 585
R575 B.n334 B.n333 585
R576 B.n335 B.n40 585
R577 B.n337 B.n336 585
R578 B.n338 B.n39 585
R579 B.n340 B.n339 585
R580 B.n341 B.n38 585
R581 B.n343 B.n342 585
R582 B.n344 B.n37 585
R583 B.n346 B.n345 585
R584 B.n347 B.n36 585
R585 B.n349 B.n348 585
R586 B.n351 B.n33 585
R587 B.n353 B.n352 585
R588 B.n354 B.n32 585
R589 B.n356 B.n355 585
R590 B.n357 B.n31 585
R591 B.n359 B.n358 585
R592 B.n360 B.n30 585
R593 B.n362 B.n361 585
R594 B.n363 B.n29 585
R595 B.n365 B.n364 585
R596 B.n367 B.n366 585
R597 B.n368 B.n25 585
R598 B.n370 B.n369 585
R599 B.n371 B.n24 585
R600 B.n373 B.n372 585
R601 B.n374 B.n23 585
R602 B.n376 B.n375 585
R603 B.n377 B.n22 585
R604 B.n379 B.n378 585
R605 B.n380 B.n21 585
R606 B.n382 B.n381 585
R607 B.n383 B.n20 585
R608 B.n385 B.n384 585
R609 B.n386 B.n19 585
R610 B.n388 B.n387 585
R611 B.n389 B.n18 585
R612 B.n391 B.n390 585
R613 B.n392 B.n17 585
R614 B.n394 B.n393 585
R615 B.n395 B.n16 585
R616 B.n397 B.n396 585
R617 B.n398 B.n15 585
R618 B.n400 B.n399 585
R619 B.n401 B.n14 585
R620 B.n403 B.n402 585
R621 B.n404 B.n13 585
R622 B.n406 B.n405 585
R623 B.n407 B.n12 585
R624 B.n409 B.n408 585
R625 B.n410 B.n11 585
R626 B.n304 B.n303 585
R627 B.n302 B.n51 585
R628 B.n301 B.n300 585
R629 B.n299 B.n52 585
R630 B.n298 B.n297 585
R631 B.n296 B.n53 585
R632 B.n295 B.n294 585
R633 B.n293 B.n54 585
R634 B.n292 B.n291 585
R635 B.n290 B.n55 585
R636 B.n289 B.n288 585
R637 B.n287 B.n56 585
R638 B.n286 B.n285 585
R639 B.n284 B.n57 585
R640 B.n283 B.n282 585
R641 B.n281 B.n58 585
R642 B.n280 B.n279 585
R643 B.n278 B.n59 585
R644 B.n277 B.n276 585
R645 B.n275 B.n60 585
R646 B.n274 B.n273 585
R647 B.n272 B.n61 585
R648 B.n271 B.n270 585
R649 B.n269 B.n62 585
R650 B.n268 B.n267 585
R651 B.n266 B.n63 585
R652 B.n265 B.n264 585
R653 B.n263 B.n64 585
R654 B.n262 B.n261 585
R655 B.n260 B.n65 585
R656 B.n259 B.n258 585
R657 B.n257 B.n66 585
R658 B.n256 B.n255 585
R659 B.n254 B.n67 585
R660 B.n253 B.n252 585
R661 B.n251 B.n68 585
R662 B.n250 B.n249 585
R663 B.n143 B.n108 585
R664 B.n145 B.n144 585
R665 B.n146 B.n107 585
R666 B.n148 B.n147 585
R667 B.n149 B.n106 585
R668 B.n151 B.n150 585
R669 B.n152 B.n105 585
R670 B.n154 B.n153 585
R671 B.n155 B.n104 585
R672 B.n157 B.n156 585
R673 B.n158 B.n103 585
R674 B.n160 B.n159 585
R675 B.n161 B.n102 585
R676 B.n163 B.n162 585
R677 B.n164 B.n101 585
R678 B.n166 B.n165 585
R679 B.n167 B.n100 585
R680 B.n169 B.n168 585
R681 B.n170 B.n99 585
R682 B.n172 B.n171 585
R683 B.n173 B.n98 585
R684 B.n175 B.n174 585
R685 B.n176 B.n97 585
R686 B.n178 B.n177 585
R687 B.n179 B.n96 585
R688 B.n181 B.n180 585
R689 B.n182 B.n95 585
R690 B.n184 B.n183 585
R691 B.n185 B.n94 585
R692 B.n187 B.n186 585
R693 B.n189 B.n91 585
R694 B.n191 B.n190 585
R695 B.n192 B.n90 585
R696 B.n194 B.n193 585
R697 B.n195 B.n89 585
R698 B.n197 B.n196 585
R699 B.n198 B.n88 585
R700 B.n200 B.n199 585
R701 B.n201 B.n87 585
R702 B.n203 B.n202 585
R703 B.n205 B.n204 585
R704 B.n206 B.n83 585
R705 B.n208 B.n207 585
R706 B.n209 B.n82 585
R707 B.n211 B.n210 585
R708 B.n212 B.n81 585
R709 B.n214 B.n213 585
R710 B.n215 B.n80 585
R711 B.n217 B.n216 585
R712 B.n218 B.n79 585
R713 B.n220 B.n219 585
R714 B.n221 B.n78 585
R715 B.n223 B.n222 585
R716 B.n224 B.n77 585
R717 B.n226 B.n225 585
R718 B.n227 B.n76 585
R719 B.n229 B.n228 585
R720 B.n230 B.n75 585
R721 B.n232 B.n231 585
R722 B.n233 B.n74 585
R723 B.n235 B.n234 585
R724 B.n236 B.n73 585
R725 B.n238 B.n237 585
R726 B.n239 B.n72 585
R727 B.n241 B.n240 585
R728 B.n242 B.n71 585
R729 B.n244 B.n243 585
R730 B.n245 B.n70 585
R731 B.n247 B.n246 585
R732 B.n248 B.n69 585
R733 B.n142 B.n141 585
R734 B.n140 B.n109 585
R735 B.n139 B.n138 585
R736 B.n137 B.n110 585
R737 B.n136 B.n135 585
R738 B.n134 B.n111 585
R739 B.n133 B.n132 585
R740 B.n131 B.n112 585
R741 B.n130 B.n129 585
R742 B.n128 B.n113 585
R743 B.n127 B.n126 585
R744 B.n125 B.n114 585
R745 B.n124 B.n123 585
R746 B.n122 B.n115 585
R747 B.n121 B.n120 585
R748 B.n119 B.n116 585
R749 B.n118 B.n117 585
R750 B.n2 B.n0 585
R751 B.n437 B.n1 585
R752 B.n436 B.n435 585
R753 B.n434 B.n3 585
R754 B.n433 B.n432 585
R755 B.n431 B.n4 585
R756 B.n430 B.n429 585
R757 B.n428 B.n5 585
R758 B.n427 B.n426 585
R759 B.n425 B.n6 585
R760 B.n424 B.n423 585
R761 B.n422 B.n7 585
R762 B.n421 B.n420 585
R763 B.n419 B.n8 585
R764 B.n418 B.n417 585
R765 B.n416 B.n9 585
R766 B.n415 B.n414 585
R767 B.n413 B.n10 585
R768 B.n412 B.n411 585
R769 B.n439 B.n438 585
R770 B.n143 B.n142 502.111
R771 B.n412 B.n11 502.111
R772 B.n250 B.n69 502.111
R773 B.n305 B.n304 502.111
R774 B.n84 B.t9 441.904
R775 B.n92 B.t0 441.904
R776 B.n26 B.t6 441.904
R777 B.n34 B.t3 441.904
R778 B.n84 B.t11 327.156
R779 B.n34 B.t4 327.156
R780 B.n92 B.t2 327.156
R781 B.n26 B.t7 327.156
R782 B.n85 B.t10 305.048
R783 B.n35 B.t5 305.048
R784 B.n93 B.t1 305.048
R785 B.n27 B.t8 305.048
R786 B.n142 B.n109 163.367
R787 B.n138 B.n109 163.367
R788 B.n138 B.n137 163.367
R789 B.n137 B.n136 163.367
R790 B.n136 B.n111 163.367
R791 B.n132 B.n111 163.367
R792 B.n132 B.n131 163.367
R793 B.n131 B.n130 163.367
R794 B.n130 B.n113 163.367
R795 B.n126 B.n113 163.367
R796 B.n126 B.n125 163.367
R797 B.n125 B.n124 163.367
R798 B.n124 B.n115 163.367
R799 B.n120 B.n115 163.367
R800 B.n120 B.n119 163.367
R801 B.n119 B.n118 163.367
R802 B.n118 B.n2 163.367
R803 B.n438 B.n2 163.367
R804 B.n438 B.n437 163.367
R805 B.n437 B.n436 163.367
R806 B.n436 B.n3 163.367
R807 B.n432 B.n3 163.367
R808 B.n432 B.n431 163.367
R809 B.n431 B.n430 163.367
R810 B.n430 B.n5 163.367
R811 B.n426 B.n5 163.367
R812 B.n426 B.n425 163.367
R813 B.n425 B.n424 163.367
R814 B.n424 B.n7 163.367
R815 B.n420 B.n7 163.367
R816 B.n420 B.n419 163.367
R817 B.n419 B.n418 163.367
R818 B.n418 B.n9 163.367
R819 B.n414 B.n9 163.367
R820 B.n414 B.n413 163.367
R821 B.n413 B.n412 163.367
R822 B.n144 B.n143 163.367
R823 B.n144 B.n107 163.367
R824 B.n148 B.n107 163.367
R825 B.n149 B.n148 163.367
R826 B.n150 B.n149 163.367
R827 B.n150 B.n105 163.367
R828 B.n154 B.n105 163.367
R829 B.n155 B.n154 163.367
R830 B.n156 B.n155 163.367
R831 B.n156 B.n103 163.367
R832 B.n160 B.n103 163.367
R833 B.n161 B.n160 163.367
R834 B.n162 B.n161 163.367
R835 B.n162 B.n101 163.367
R836 B.n166 B.n101 163.367
R837 B.n167 B.n166 163.367
R838 B.n168 B.n167 163.367
R839 B.n168 B.n99 163.367
R840 B.n172 B.n99 163.367
R841 B.n173 B.n172 163.367
R842 B.n174 B.n173 163.367
R843 B.n174 B.n97 163.367
R844 B.n178 B.n97 163.367
R845 B.n179 B.n178 163.367
R846 B.n180 B.n179 163.367
R847 B.n180 B.n95 163.367
R848 B.n184 B.n95 163.367
R849 B.n185 B.n184 163.367
R850 B.n186 B.n185 163.367
R851 B.n186 B.n91 163.367
R852 B.n191 B.n91 163.367
R853 B.n192 B.n191 163.367
R854 B.n193 B.n192 163.367
R855 B.n193 B.n89 163.367
R856 B.n197 B.n89 163.367
R857 B.n198 B.n197 163.367
R858 B.n199 B.n198 163.367
R859 B.n199 B.n87 163.367
R860 B.n203 B.n87 163.367
R861 B.n204 B.n203 163.367
R862 B.n204 B.n83 163.367
R863 B.n208 B.n83 163.367
R864 B.n209 B.n208 163.367
R865 B.n210 B.n209 163.367
R866 B.n210 B.n81 163.367
R867 B.n214 B.n81 163.367
R868 B.n215 B.n214 163.367
R869 B.n216 B.n215 163.367
R870 B.n216 B.n79 163.367
R871 B.n220 B.n79 163.367
R872 B.n221 B.n220 163.367
R873 B.n222 B.n221 163.367
R874 B.n222 B.n77 163.367
R875 B.n226 B.n77 163.367
R876 B.n227 B.n226 163.367
R877 B.n228 B.n227 163.367
R878 B.n228 B.n75 163.367
R879 B.n232 B.n75 163.367
R880 B.n233 B.n232 163.367
R881 B.n234 B.n233 163.367
R882 B.n234 B.n73 163.367
R883 B.n238 B.n73 163.367
R884 B.n239 B.n238 163.367
R885 B.n240 B.n239 163.367
R886 B.n240 B.n71 163.367
R887 B.n244 B.n71 163.367
R888 B.n245 B.n244 163.367
R889 B.n246 B.n245 163.367
R890 B.n246 B.n69 163.367
R891 B.n251 B.n250 163.367
R892 B.n252 B.n251 163.367
R893 B.n252 B.n67 163.367
R894 B.n256 B.n67 163.367
R895 B.n257 B.n256 163.367
R896 B.n258 B.n257 163.367
R897 B.n258 B.n65 163.367
R898 B.n262 B.n65 163.367
R899 B.n263 B.n262 163.367
R900 B.n264 B.n263 163.367
R901 B.n264 B.n63 163.367
R902 B.n268 B.n63 163.367
R903 B.n269 B.n268 163.367
R904 B.n270 B.n269 163.367
R905 B.n270 B.n61 163.367
R906 B.n274 B.n61 163.367
R907 B.n275 B.n274 163.367
R908 B.n276 B.n275 163.367
R909 B.n276 B.n59 163.367
R910 B.n280 B.n59 163.367
R911 B.n281 B.n280 163.367
R912 B.n282 B.n281 163.367
R913 B.n282 B.n57 163.367
R914 B.n286 B.n57 163.367
R915 B.n287 B.n286 163.367
R916 B.n288 B.n287 163.367
R917 B.n288 B.n55 163.367
R918 B.n292 B.n55 163.367
R919 B.n293 B.n292 163.367
R920 B.n294 B.n293 163.367
R921 B.n294 B.n53 163.367
R922 B.n298 B.n53 163.367
R923 B.n299 B.n298 163.367
R924 B.n300 B.n299 163.367
R925 B.n300 B.n51 163.367
R926 B.n304 B.n51 163.367
R927 B.n408 B.n11 163.367
R928 B.n408 B.n407 163.367
R929 B.n407 B.n406 163.367
R930 B.n406 B.n13 163.367
R931 B.n402 B.n13 163.367
R932 B.n402 B.n401 163.367
R933 B.n401 B.n400 163.367
R934 B.n400 B.n15 163.367
R935 B.n396 B.n15 163.367
R936 B.n396 B.n395 163.367
R937 B.n395 B.n394 163.367
R938 B.n394 B.n17 163.367
R939 B.n390 B.n17 163.367
R940 B.n390 B.n389 163.367
R941 B.n389 B.n388 163.367
R942 B.n388 B.n19 163.367
R943 B.n384 B.n19 163.367
R944 B.n384 B.n383 163.367
R945 B.n383 B.n382 163.367
R946 B.n382 B.n21 163.367
R947 B.n378 B.n21 163.367
R948 B.n378 B.n377 163.367
R949 B.n377 B.n376 163.367
R950 B.n376 B.n23 163.367
R951 B.n372 B.n23 163.367
R952 B.n372 B.n371 163.367
R953 B.n371 B.n370 163.367
R954 B.n370 B.n25 163.367
R955 B.n366 B.n25 163.367
R956 B.n366 B.n365 163.367
R957 B.n365 B.n29 163.367
R958 B.n361 B.n29 163.367
R959 B.n361 B.n360 163.367
R960 B.n360 B.n359 163.367
R961 B.n359 B.n31 163.367
R962 B.n355 B.n31 163.367
R963 B.n355 B.n354 163.367
R964 B.n354 B.n353 163.367
R965 B.n353 B.n33 163.367
R966 B.n348 B.n33 163.367
R967 B.n348 B.n347 163.367
R968 B.n347 B.n346 163.367
R969 B.n346 B.n37 163.367
R970 B.n342 B.n37 163.367
R971 B.n342 B.n341 163.367
R972 B.n341 B.n340 163.367
R973 B.n340 B.n39 163.367
R974 B.n336 B.n39 163.367
R975 B.n336 B.n335 163.367
R976 B.n335 B.n334 163.367
R977 B.n334 B.n41 163.367
R978 B.n330 B.n41 163.367
R979 B.n330 B.n329 163.367
R980 B.n329 B.n328 163.367
R981 B.n328 B.n43 163.367
R982 B.n324 B.n43 163.367
R983 B.n324 B.n323 163.367
R984 B.n323 B.n322 163.367
R985 B.n322 B.n45 163.367
R986 B.n318 B.n45 163.367
R987 B.n318 B.n317 163.367
R988 B.n317 B.n316 163.367
R989 B.n316 B.n47 163.367
R990 B.n312 B.n47 163.367
R991 B.n312 B.n311 163.367
R992 B.n311 B.n310 163.367
R993 B.n310 B.n49 163.367
R994 B.n306 B.n49 163.367
R995 B.n306 B.n305 163.367
R996 B.n86 B.n85 59.5399
R997 B.n188 B.n93 59.5399
R998 B.n28 B.n27 59.5399
R999 B.n350 B.n35 59.5399
R1000 B.n411 B.n410 32.6249
R1001 B.n303 B.n50 32.6249
R1002 B.n249 B.n248 32.6249
R1003 B.n141 B.n108 32.6249
R1004 B.n85 B.n84 22.1096
R1005 B.n93 B.n92 22.1096
R1006 B.n27 B.n26 22.1096
R1007 B.n35 B.n34 22.1096
R1008 B B.n439 18.0485
R1009 B.n410 B.n409 10.6151
R1010 B.n409 B.n12 10.6151
R1011 B.n405 B.n12 10.6151
R1012 B.n405 B.n404 10.6151
R1013 B.n404 B.n403 10.6151
R1014 B.n403 B.n14 10.6151
R1015 B.n399 B.n14 10.6151
R1016 B.n399 B.n398 10.6151
R1017 B.n398 B.n397 10.6151
R1018 B.n397 B.n16 10.6151
R1019 B.n393 B.n16 10.6151
R1020 B.n393 B.n392 10.6151
R1021 B.n392 B.n391 10.6151
R1022 B.n391 B.n18 10.6151
R1023 B.n387 B.n18 10.6151
R1024 B.n387 B.n386 10.6151
R1025 B.n386 B.n385 10.6151
R1026 B.n385 B.n20 10.6151
R1027 B.n381 B.n20 10.6151
R1028 B.n381 B.n380 10.6151
R1029 B.n380 B.n379 10.6151
R1030 B.n379 B.n22 10.6151
R1031 B.n375 B.n22 10.6151
R1032 B.n375 B.n374 10.6151
R1033 B.n374 B.n373 10.6151
R1034 B.n373 B.n24 10.6151
R1035 B.n369 B.n24 10.6151
R1036 B.n369 B.n368 10.6151
R1037 B.n368 B.n367 10.6151
R1038 B.n364 B.n363 10.6151
R1039 B.n363 B.n362 10.6151
R1040 B.n362 B.n30 10.6151
R1041 B.n358 B.n30 10.6151
R1042 B.n358 B.n357 10.6151
R1043 B.n357 B.n356 10.6151
R1044 B.n356 B.n32 10.6151
R1045 B.n352 B.n32 10.6151
R1046 B.n352 B.n351 10.6151
R1047 B.n349 B.n36 10.6151
R1048 B.n345 B.n36 10.6151
R1049 B.n345 B.n344 10.6151
R1050 B.n344 B.n343 10.6151
R1051 B.n343 B.n38 10.6151
R1052 B.n339 B.n38 10.6151
R1053 B.n339 B.n338 10.6151
R1054 B.n338 B.n337 10.6151
R1055 B.n337 B.n40 10.6151
R1056 B.n333 B.n40 10.6151
R1057 B.n333 B.n332 10.6151
R1058 B.n332 B.n331 10.6151
R1059 B.n331 B.n42 10.6151
R1060 B.n327 B.n42 10.6151
R1061 B.n327 B.n326 10.6151
R1062 B.n326 B.n325 10.6151
R1063 B.n325 B.n44 10.6151
R1064 B.n321 B.n44 10.6151
R1065 B.n321 B.n320 10.6151
R1066 B.n320 B.n319 10.6151
R1067 B.n319 B.n46 10.6151
R1068 B.n315 B.n46 10.6151
R1069 B.n315 B.n314 10.6151
R1070 B.n314 B.n313 10.6151
R1071 B.n313 B.n48 10.6151
R1072 B.n309 B.n48 10.6151
R1073 B.n309 B.n308 10.6151
R1074 B.n308 B.n307 10.6151
R1075 B.n307 B.n50 10.6151
R1076 B.n249 B.n68 10.6151
R1077 B.n253 B.n68 10.6151
R1078 B.n254 B.n253 10.6151
R1079 B.n255 B.n254 10.6151
R1080 B.n255 B.n66 10.6151
R1081 B.n259 B.n66 10.6151
R1082 B.n260 B.n259 10.6151
R1083 B.n261 B.n260 10.6151
R1084 B.n261 B.n64 10.6151
R1085 B.n265 B.n64 10.6151
R1086 B.n266 B.n265 10.6151
R1087 B.n267 B.n266 10.6151
R1088 B.n267 B.n62 10.6151
R1089 B.n271 B.n62 10.6151
R1090 B.n272 B.n271 10.6151
R1091 B.n273 B.n272 10.6151
R1092 B.n273 B.n60 10.6151
R1093 B.n277 B.n60 10.6151
R1094 B.n278 B.n277 10.6151
R1095 B.n279 B.n278 10.6151
R1096 B.n279 B.n58 10.6151
R1097 B.n283 B.n58 10.6151
R1098 B.n284 B.n283 10.6151
R1099 B.n285 B.n284 10.6151
R1100 B.n285 B.n56 10.6151
R1101 B.n289 B.n56 10.6151
R1102 B.n290 B.n289 10.6151
R1103 B.n291 B.n290 10.6151
R1104 B.n291 B.n54 10.6151
R1105 B.n295 B.n54 10.6151
R1106 B.n296 B.n295 10.6151
R1107 B.n297 B.n296 10.6151
R1108 B.n297 B.n52 10.6151
R1109 B.n301 B.n52 10.6151
R1110 B.n302 B.n301 10.6151
R1111 B.n303 B.n302 10.6151
R1112 B.n145 B.n108 10.6151
R1113 B.n146 B.n145 10.6151
R1114 B.n147 B.n146 10.6151
R1115 B.n147 B.n106 10.6151
R1116 B.n151 B.n106 10.6151
R1117 B.n152 B.n151 10.6151
R1118 B.n153 B.n152 10.6151
R1119 B.n153 B.n104 10.6151
R1120 B.n157 B.n104 10.6151
R1121 B.n158 B.n157 10.6151
R1122 B.n159 B.n158 10.6151
R1123 B.n159 B.n102 10.6151
R1124 B.n163 B.n102 10.6151
R1125 B.n164 B.n163 10.6151
R1126 B.n165 B.n164 10.6151
R1127 B.n165 B.n100 10.6151
R1128 B.n169 B.n100 10.6151
R1129 B.n170 B.n169 10.6151
R1130 B.n171 B.n170 10.6151
R1131 B.n171 B.n98 10.6151
R1132 B.n175 B.n98 10.6151
R1133 B.n176 B.n175 10.6151
R1134 B.n177 B.n176 10.6151
R1135 B.n177 B.n96 10.6151
R1136 B.n181 B.n96 10.6151
R1137 B.n182 B.n181 10.6151
R1138 B.n183 B.n182 10.6151
R1139 B.n183 B.n94 10.6151
R1140 B.n187 B.n94 10.6151
R1141 B.n190 B.n189 10.6151
R1142 B.n190 B.n90 10.6151
R1143 B.n194 B.n90 10.6151
R1144 B.n195 B.n194 10.6151
R1145 B.n196 B.n195 10.6151
R1146 B.n196 B.n88 10.6151
R1147 B.n200 B.n88 10.6151
R1148 B.n201 B.n200 10.6151
R1149 B.n202 B.n201 10.6151
R1150 B.n206 B.n205 10.6151
R1151 B.n207 B.n206 10.6151
R1152 B.n207 B.n82 10.6151
R1153 B.n211 B.n82 10.6151
R1154 B.n212 B.n211 10.6151
R1155 B.n213 B.n212 10.6151
R1156 B.n213 B.n80 10.6151
R1157 B.n217 B.n80 10.6151
R1158 B.n218 B.n217 10.6151
R1159 B.n219 B.n218 10.6151
R1160 B.n219 B.n78 10.6151
R1161 B.n223 B.n78 10.6151
R1162 B.n224 B.n223 10.6151
R1163 B.n225 B.n224 10.6151
R1164 B.n225 B.n76 10.6151
R1165 B.n229 B.n76 10.6151
R1166 B.n230 B.n229 10.6151
R1167 B.n231 B.n230 10.6151
R1168 B.n231 B.n74 10.6151
R1169 B.n235 B.n74 10.6151
R1170 B.n236 B.n235 10.6151
R1171 B.n237 B.n236 10.6151
R1172 B.n237 B.n72 10.6151
R1173 B.n241 B.n72 10.6151
R1174 B.n242 B.n241 10.6151
R1175 B.n243 B.n242 10.6151
R1176 B.n243 B.n70 10.6151
R1177 B.n247 B.n70 10.6151
R1178 B.n248 B.n247 10.6151
R1179 B.n141 B.n140 10.6151
R1180 B.n140 B.n139 10.6151
R1181 B.n139 B.n110 10.6151
R1182 B.n135 B.n110 10.6151
R1183 B.n135 B.n134 10.6151
R1184 B.n134 B.n133 10.6151
R1185 B.n133 B.n112 10.6151
R1186 B.n129 B.n112 10.6151
R1187 B.n129 B.n128 10.6151
R1188 B.n128 B.n127 10.6151
R1189 B.n127 B.n114 10.6151
R1190 B.n123 B.n114 10.6151
R1191 B.n123 B.n122 10.6151
R1192 B.n122 B.n121 10.6151
R1193 B.n121 B.n116 10.6151
R1194 B.n117 B.n116 10.6151
R1195 B.n117 B.n0 10.6151
R1196 B.n435 B.n1 10.6151
R1197 B.n435 B.n434 10.6151
R1198 B.n434 B.n433 10.6151
R1199 B.n433 B.n4 10.6151
R1200 B.n429 B.n4 10.6151
R1201 B.n429 B.n428 10.6151
R1202 B.n428 B.n427 10.6151
R1203 B.n427 B.n6 10.6151
R1204 B.n423 B.n6 10.6151
R1205 B.n423 B.n422 10.6151
R1206 B.n422 B.n421 10.6151
R1207 B.n421 B.n8 10.6151
R1208 B.n417 B.n8 10.6151
R1209 B.n417 B.n416 10.6151
R1210 B.n416 B.n415 10.6151
R1211 B.n415 B.n10 10.6151
R1212 B.n411 B.n10 10.6151
R1213 B.n367 B.n28 9.36635
R1214 B.n350 B.n349 9.36635
R1215 B.n188 B.n187 9.36635
R1216 B.n205 B.n86 9.36635
R1217 B.n439 B.n0 2.81026
R1218 B.n439 B.n1 2.81026
R1219 B.n364 B.n28 1.24928
R1220 B.n351 B.n350 1.24928
R1221 B.n189 B.n188 1.24928
R1222 B.n202 B.n86 1.24928
R1223 VN.n0 VN.t3 309.899
R1224 VN.n1 VN.t0 309.899
R1225 VN.n0 VN.t1 309.849
R1226 VN.n1 VN.t2 309.849
R1227 VN VN.n1 82.8912
R1228 VN VN.n0 44.7132
R1229 VDD2.n2 VDD2.n0 114.662
R1230 VDD2.n2 VDD2.n1 81.0415
R1231 VDD2.n1 VDD2.t1 4.02838
R1232 VDD2.n1 VDD2.t3 4.02838
R1233 VDD2.n0 VDD2.t0 4.02838
R1234 VDD2.n0 VDD2.t2 4.02838
R1235 VDD2 VDD2.n2 0.0586897
C0 VDD1 VN 0.14719f
C1 VP w_n1654_n2582# 2.60368f
C2 w_n1654_n2582# VDD2 0.997166f
C3 VTAIL B 2.82245f
C4 VN w_n1654_n2582# 2.39558f
C5 VP B 1.05859f
C6 B VDD2 0.862874f
C7 VTAIL VP 2.15818f
C8 VTAIL VDD2 4.8849f
C9 VN B 0.721583f
C10 VDD1 w_n1654_n2582# 0.98043f
C11 VP VDD2 0.280212f
C12 VTAIL VN 2.14407f
C13 VDD1 B 0.839777f
C14 VN VP 4.17191f
C15 VN VDD2 2.36004f
C16 VTAIL VDD1 4.84269f
C17 VDD1 VP 2.49277f
C18 B w_n1654_n2582# 5.94115f
C19 VDD1 VDD2 0.591799f
C20 VTAIL w_n1654_n2582# 3.11593f
C21 VDD2 VSUBS 0.594486f
C22 VDD1 VSUBS 4.321982f
C23 VTAIL VSUBS 0.730327f
C24 VN VSUBS 5.3713f
C25 VP VSUBS 1.206629f
C26 B VSUBS 2.382494f
C27 w_n1654_n2582# VSUBS 52.9743f
C28 VDD2.t0 VSUBS 0.177494f
C29 VDD2.t2 VSUBS 0.177494f
C30 VDD2.n0 VSUBS 1.73758f
C31 VDD2.t1 VSUBS 0.177494f
C32 VDD2.t3 VSUBS 0.177494f
C33 VDD2.n1 VSUBS 1.26374f
C34 VDD2.n2 VSUBS 3.49458f
C35 VN.t3 VSUBS 1.17096f
C36 VN.t1 VSUBS 1.17087f
C37 VN.n0 VSUBS 0.913377f
C38 VN.t0 VSUBS 1.17096f
C39 VN.t2 VSUBS 1.17087f
C40 VN.n1 VSUBS 1.95719f
C41 B.n0 VSUBS 0.005463f
C42 B.n1 VSUBS 0.005463f
C43 B.n2 VSUBS 0.00864f
C44 B.n3 VSUBS 0.00864f
C45 B.n4 VSUBS 0.00864f
C46 B.n5 VSUBS 0.00864f
C47 B.n6 VSUBS 0.00864f
C48 B.n7 VSUBS 0.00864f
C49 B.n8 VSUBS 0.00864f
C50 B.n9 VSUBS 0.00864f
C51 B.n10 VSUBS 0.00864f
C52 B.n11 VSUBS 0.020962f
C53 B.n12 VSUBS 0.00864f
C54 B.n13 VSUBS 0.00864f
C55 B.n14 VSUBS 0.00864f
C56 B.n15 VSUBS 0.00864f
C57 B.n16 VSUBS 0.00864f
C58 B.n17 VSUBS 0.00864f
C59 B.n18 VSUBS 0.00864f
C60 B.n19 VSUBS 0.00864f
C61 B.n20 VSUBS 0.00864f
C62 B.n21 VSUBS 0.00864f
C63 B.n22 VSUBS 0.00864f
C64 B.n23 VSUBS 0.00864f
C65 B.n24 VSUBS 0.00864f
C66 B.n25 VSUBS 0.00864f
C67 B.t8 VSUBS 0.158165f
C68 B.t7 VSUBS 0.17278f
C69 B.t6 VSUBS 0.345483f
C70 B.n26 VSUBS 0.27971f
C71 B.n27 VSUBS 0.228592f
C72 B.n28 VSUBS 0.020017f
C73 B.n29 VSUBS 0.00864f
C74 B.n30 VSUBS 0.00864f
C75 B.n31 VSUBS 0.00864f
C76 B.n32 VSUBS 0.00864f
C77 B.n33 VSUBS 0.00864f
C78 B.t5 VSUBS 0.158168f
C79 B.t4 VSUBS 0.172783f
C80 B.t3 VSUBS 0.345483f
C81 B.n34 VSUBS 0.279707f
C82 B.n35 VSUBS 0.228589f
C83 B.n36 VSUBS 0.00864f
C84 B.n37 VSUBS 0.00864f
C85 B.n38 VSUBS 0.00864f
C86 B.n39 VSUBS 0.00864f
C87 B.n40 VSUBS 0.00864f
C88 B.n41 VSUBS 0.00864f
C89 B.n42 VSUBS 0.00864f
C90 B.n43 VSUBS 0.00864f
C91 B.n44 VSUBS 0.00864f
C92 B.n45 VSUBS 0.00864f
C93 B.n46 VSUBS 0.00864f
C94 B.n47 VSUBS 0.00864f
C95 B.n48 VSUBS 0.00864f
C96 B.n49 VSUBS 0.00864f
C97 B.n50 VSUBS 0.01994f
C98 B.n51 VSUBS 0.00864f
C99 B.n52 VSUBS 0.00864f
C100 B.n53 VSUBS 0.00864f
C101 B.n54 VSUBS 0.00864f
C102 B.n55 VSUBS 0.00864f
C103 B.n56 VSUBS 0.00864f
C104 B.n57 VSUBS 0.00864f
C105 B.n58 VSUBS 0.00864f
C106 B.n59 VSUBS 0.00864f
C107 B.n60 VSUBS 0.00864f
C108 B.n61 VSUBS 0.00864f
C109 B.n62 VSUBS 0.00864f
C110 B.n63 VSUBS 0.00864f
C111 B.n64 VSUBS 0.00864f
C112 B.n65 VSUBS 0.00864f
C113 B.n66 VSUBS 0.00864f
C114 B.n67 VSUBS 0.00864f
C115 B.n68 VSUBS 0.00864f
C116 B.n69 VSUBS 0.020962f
C117 B.n70 VSUBS 0.00864f
C118 B.n71 VSUBS 0.00864f
C119 B.n72 VSUBS 0.00864f
C120 B.n73 VSUBS 0.00864f
C121 B.n74 VSUBS 0.00864f
C122 B.n75 VSUBS 0.00864f
C123 B.n76 VSUBS 0.00864f
C124 B.n77 VSUBS 0.00864f
C125 B.n78 VSUBS 0.00864f
C126 B.n79 VSUBS 0.00864f
C127 B.n80 VSUBS 0.00864f
C128 B.n81 VSUBS 0.00864f
C129 B.n82 VSUBS 0.00864f
C130 B.n83 VSUBS 0.00864f
C131 B.t10 VSUBS 0.158168f
C132 B.t11 VSUBS 0.172783f
C133 B.t9 VSUBS 0.345483f
C134 B.n84 VSUBS 0.279707f
C135 B.n85 VSUBS 0.228589f
C136 B.n86 VSUBS 0.020017f
C137 B.n87 VSUBS 0.00864f
C138 B.n88 VSUBS 0.00864f
C139 B.n89 VSUBS 0.00864f
C140 B.n90 VSUBS 0.00864f
C141 B.n91 VSUBS 0.00864f
C142 B.t1 VSUBS 0.158165f
C143 B.t2 VSUBS 0.17278f
C144 B.t0 VSUBS 0.345483f
C145 B.n92 VSUBS 0.27971f
C146 B.n93 VSUBS 0.228592f
C147 B.n94 VSUBS 0.00864f
C148 B.n95 VSUBS 0.00864f
C149 B.n96 VSUBS 0.00864f
C150 B.n97 VSUBS 0.00864f
C151 B.n98 VSUBS 0.00864f
C152 B.n99 VSUBS 0.00864f
C153 B.n100 VSUBS 0.00864f
C154 B.n101 VSUBS 0.00864f
C155 B.n102 VSUBS 0.00864f
C156 B.n103 VSUBS 0.00864f
C157 B.n104 VSUBS 0.00864f
C158 B.n105 VSUBS 0.00864f
C159 B.n106 VSUBS 0.00864f
C160 B.n107 VSUBS 0.00864f
C161 B.n108 VSUBS 0.020962f
C162 B.n109 VSUBS 0.00864f
C163 B.n110 VSUBS 0.00864f
C164 B.n111 VSUBS 0.00864f
C165 B.n112 VSUBS 0.00864f
C166 B.n113 VSUBS 0.00864f
C167 B.n114 VSUBS 0.00864f
C168 B.n115 VSUBS 0.00864f
C169 B.n116 VSUBS 0.00864f
C170 B.n117 VSUBS 0.00864f
C171 B.n118 VSUBS 0.00864f
C172 B.n119 VSUBS 0.00864f
C173 B.n120 VSUBS 0.00864f
C174 B.n121 VSUBS 0.00864f
C175 B.n122 VSUBS 0.00864f
C176 B.n123 VSUBS 0.00864f
C177 B.n124 VSUBS 0.00864f
C178 B.n125 VSUBS 0.00864f
C179 B.n126 VSUBS 0.00864f
C180 B.n127 VSUBS 0.00864f
C181 B.n128 VSUBS 0.00864f
C182 B.n129 VSUBS 0.00864f
C183 B.n130 VSUBS 0.00864f
C184 B.n131 VSUBS 0.00864f
C185 B.n132 VSUBS 0.00864f
C186 B.n133 VSUBS 0.00864f
C187 B.n134 VSUBS 0.00864f
C188 B.n135 VSUBS 0.00864f
C189 B.n136 VSUBS 0.00864f
C190 B.n137 VSUBS 0.00864f
C191 B.n138 VSUBS 0.00864f
C192 B.n139 VSUBS 0.00864f
C193 B.n140 VSUBS 0.00864f
C194 B.n141 VSUBS 0.019441f
C195 B.n142 VSUBS 0.019441f
C196 B.n143 VSUBS 0.020962f
C197 B.n144 VSUBS 0.00864f
C198 B.n145 VSUBS 0.00864f
C199 B.n146 VSUBS 0.00864f
C200 B.n147 VSUBS 0.00864f
C201 B.n148 VSUBS 0.00864f
C202 B.n149 VSUBS 0.00864f
C203 B.n150 VSUBS 0.00864f
C204 B.n151 VSUBS 0.00864f
C205 B.n152 VSUBS 0.00864f
C206 B.n153 VSUBS 0.00864f
C207 B.n154 VSUBS 0.00864f
C208 B.n155 VSUBS 0.00864f
C209 B.n156 VSUBS 0.00864f
C210 B.n157 VSUBS 0.00864f
C211 B.n158 VSUBS 0.00864f
C212 B.n159 VSUBS 0.00864f
C213 B.n160 VSUBS 0.00864f
C214 B.n161 VSUBS 0.00864f
C215 B.n162 VSUBS 0.00864f
C216 B.n163 VSUBS 0.00864f
C217 B.n164 VSUBS 0.00864f
C218 B.n165 VSUBS 0.00864f
C219 B.n166 VSUBS 0.00864f
C220 B.n167 VSUBS 0.00864f
C221 B.n168 VSUBS 0.00864f
C222 B.n169 VSUBS 0.00864f
C223 B.n170 VSUBS 0.00864f
C224 B.n171 VSUBS 0.00864f
C225 B.n172 VSUBS 0.00864f
C226 B.n173 VSUBS 0.00864f
C227 B.n174 VSUBS 0.00864f
C228 B.n175 VSUBS 0.00864f
C229 B.n176 VSUBS 0.00864f
C230 B.n177 VSUBS 0.00864f
C231 B.n178 VSUBS 0.00864f
C232 B.n179 VSUBS 0.00864f
C233 B.n180 VSUBS 0.00864f
C234 B.n181 VSUBS 0.00864f
C235 B.n182 VSUBS 0.00864f
C236 B.n183 VSUBS 0.00864f
C237 B.n184 VSUBS 0.00864f
C238 B.n185 VSUBS 0.00864f
C239 B.n186 VSUBS 0.00864f
C240 B.n187 VSUBS 0.008132f
C241 B.n188 VSUBS 0.020017f
C242 B.n189 VSUBS 0.004828f
C243 B.n190 VSUBS 0.00864f
C244 B.n191 VSUBS 0.00864f
C245 B.n192 VSUBS 0.00864f
C246 B.n193 VSUBS 0.00864f
C247 B.n194 VSUBS 0.00864f
C248 B.n195 VSUBS 0.00864f
C249 B.n196 VSUBS 0.00864f
C250 B.n197 VSUBS 0.00864f
C251 B.n198 VSUBS 0.00864f
C252 B.n199 VSUBS 0.00864f
C253 B.n200 VSUBS 0.00864f
C254 B.n201 VSUBS 0.00864f
C255 B.n202 VSUBS 0.004828f
C256 B.n203 VSUBS 0.00864f
C257 B.n204 VSUBS 0.00864f
C258 B.n205 VSUBS 0.008132f
C259 B.n206 VSUBS 0.00864f
C260 B.n207 VSUBS 0.00864f
C261 B.n208 VSUBS 0.00864f
C262 B.n209 VSUBS 0.00864f
C263 B.n210 VSUBS 0.00864f
C264 B.n211 VSUBS 0.00864f
C265 B.n212 VSUBS 0.00864f
C266 B.n213 VSUBS 0.00864f
C267 B.n214 VSUBS 0.00864f
C268 B.n215 VSUBS 0.00864f
C269 B.n216 VSUBS 0.00864f
C270 B.n217 VSUBS 0.00864f
C271 B.n218 VSUBS 0.00864f
C272 B.n219 VSUBS 0.00864f
C273 B.n220 VSUBS 0.00864f
C274 B.n221 VSUBS 0.00864f
C275 B.n222 VSUBS 0.00864f
C276 B.n223 VSUBS 0.00864f
C277 B.n224 VSUBS 0.00864f
C278 B.n225 VSUBS 0.00864f
C279 B.n226 VSUBS 0.00864f
C280 B.n227 VSUBS 0.00864f
C281 B.n228 VSUBS 0.00864f
C282 B.n229 VSUBS 0.00864f
C283 B.n230 VSUBS 0.00864f
C284 B.n231 VSUBS 0.00864f
C285 B.n232 VSUBS 0.00864f
C286 B.n233 VSUBS 0.00864f
C287 B.n234 VSUBS 0.00864f
C288 B.n235 VSUBS 0.00864f
C289 B.n236 VSUBS 0.00864f
C290 B.n237 VSUBS 0.00864f
C291 B.n238 VSUBS 0.00864f
C292 B.n239 VSUBS 0.00864f
C293 B.n240 VSUBS 0.00864f
C294 B.n241 VSUBS 0.00864f
C295 B.n242 VSUBS 0.00864f
C296 B.n243 VSUBS 0.00864f
C297 B.n244 VSUBS 0.00864f
C298 B.n245 VSUBS 0.00864f
C299 B.n246 VSUBS 0.00864f
C300 B.n247 VSUBS 0.00864f
C301 B.n248 VSUBS 0.020962f
C302 B.n249 VSUBS 0.019441f
C303 B.n250 VSUBS 0.019441f
C304 B.n251 VSUBS 0.00864f
C305 B.n252 VSUBS 0.00864f
C306 B.n253 VSUBS 0.00864f
C307 B.n254 VSUBS 0.00864f
C308 B.n255 VSUBS 0.00864f
C309 B.n256 VSUBS 0.00864f
C310 B.n257 VSUBS 0.00864f
C311 B.n258 VSUBS 0.00864f
C312 B.n259 VSUBS 0.00864f
C313 B.n260 VSUBS 0.00864f
C314 B.n261 VSUBS 0.00864f
C315 B.n262 VSUBS 0.00864f
C316 B.n263 VSUBS 0.00864f
C317 B.n264 VSUBS 0.00864f
C318 B.n265 VSUBS 0.00864f
C319 B.n266 VSUBS 0.00864f
C320 B.n267 VSUBS 0.00864f
C321 B.n268 VSUBS 0.00864f
C322 B.n269 VSUBS 0.00864f
C323 B.n270 VSUBS 0.00864f
C324 B.n271 VSUBS 0.00864f
C325 B.n272 VSUBS 0.00864f
C326 B.n273 VSUBS 0.00864f
C327 B.n274 VSUBS 0.00864f
C328 B.n275 VSUBS 0.00864f
C329 B.n276 VSUBS 0.00864f
C330 B.n277 VSUBS 0.00864f
C331 B.n278 VSUBS 0.00864f
C332 B.n279 VSUBS 0.00864f
C333 B.n280 VSUBS 0.00864f
C334 B.n281 VSUBS 0.00864f
C335 B.n282 VSUBS 0.00864f
C336 B.n283 VSUBS 0.00864f
C337 B.n284 VSUBS 0.00864f
C338 B.n285 VSUBS 0.00864f
C339 B.n286 VSUBS 0.00864f
C340 B.n287 VSUBS 0.00864f
C341 B.n288 VSUBS 0.00864f
C342 B.n289 VSUBS 0.00864f
C343 B.n290 VSUBS 0.00864f
C344 B.n291 VSUBS 0.00864f
C345 B.n292 VSUBS 0.00864f
C346 B.n293 VSUBS 0.00864f
C347 B.n294 VSUBS 0.00864f
C348 B.n295 VSUBS 0.00864f
C349 B.n296 VSUBS 0.00864f
C350 B.n297 VSUBS 0.00864f
C351 B.n298 VSUBS 0.00864f
C352 B.n299 VSUBS 0.00864f
C353 B.n300 VSUBS 0.00864f
C354 B.n301 VSUBS 0.00864f
C355 B.n302 VSUBS 0.00864f
C356 B.n303 VSUBS 0.020463f
C357 B.n304 VSUBS 0.019441f
C358 B.n305 VSUBS 0.020962f
C359 B.n306 VSUBS 0.00864f
C360 B.n307 VSUBS 0.00864f
C361 B.n308 VSUBS 0.00864f
C362 B.n309 VSUBS 0.00864f
C363 B.n310 VSUBS 0.00864f
C364 B.n311 VSUBS 0.00864f
C365 B.n312 VSUBS 0.00864f
C366 B.n313 VSUBS 0.00864f
C367 B.n314 VSUBS 0.00864f
C368 B.n315 VSUBS 0.00864f
C369 B.n316 VSUBS 0.00864f
C370 B.n317 VSUBS 0.00864f
C371 B.n318 VSUBS 0.00864f
C372 B.n319 VSUBS 0.00864f
C373 B.n320 VSUBS 0.00864f
C374 B.n321 VSUBS 0.00864f
C375 B.n322 VSUBS 0.00864f
C376 B.n323 VSUBS 0.00864f
C377 B.n324 VSUBS 0.00864f
C378 B.n325 VSUBS 0.00864f
C379 B.n326 VSUBS 0.00864f
C380 B.n327 VSUBS 0.00864f
C381 B.n328 VSUBS 0.00864f
C382 B.n329 VSUBS 0.00864f
C383 B.n330 VSUBS 0.00864f
C384 B.n331 VSUBS 0.00864f
C385 B.n332 VSUBS 0.00864f
C386 B.n333 VSUBS 0.00864f
C387 B.n334 VSUBS 0.00864f
C388 B.n335 VSUBS 0.00864f
C389 B.n336 VSUBS 0.00864f
C390 B.n337 VSUBS 0.00864f
C391 B.n338 VSUBS 0.00864f
C392 B.n339 VSUBS 0.00864f
C393 B.n340 VSUBS 0.00864f
C394 B.n341 VSUBS 0.00864f
C395 B.n342 VSUBS 0.00864f
C396 B.n343 VSUBS 0.00864f
C397 B.n344 VSUBS 0.00864f
C398 B.n345 VSUBS 0.00864f
C399 B.n346 VSUBS 0.00864f
C400 B.n347 VSUBS 0.00864f
C401 B.n348 VSUBS 0.00864f
C402 B.n349 VSUBS 0.008132f
C403 B.n350 VSUBS 0.020017f
C404 B.n351 VSUBS 0.004828f
C405 B.n352 VSUBS 0.00864f
C406 B.n353 VSUBS 0.00864f
C407 B.n354 VSUBS 0.00864f
C408 B.n355 VSUBS 0.00864f
C409 B.n356 VSUBS 0.00864f
C410 B.n357 VSUBS 0.00864f
C411 B.n358 VSUBS 0.00864f
C412 B.n359 VSUBS 0.00864f
C413 B.n360 VSUBS 0.00864f
C414 B.n361 VSUBS 0.00864f
C415 B.n362 VSUBS 0.00864f
C416 B.n363 VSUBS 0.00864f
C417 B.n364 VSUBS 0.004828f
C418 B.n365 VSUBS 0.00864f
C419 B.n366 VSUBS 0.00864f
C420 B.n367 VSUBS 0.008132f
C421 B.n368 VSUBS 0.00864f
C422 B.n369 VSUBS 0.00864f
C423 B.n370 VSUBS 0.00864f
C424 B.n371 VSUBS 0.00864f
C425 B.n372 VSUBS 0.00864f
C426 B.n373 VSUBS 0.00864f
C427 B.n374 VSUBS 0.00864f
C428 B.n375 VSUBS 0.00864f
C429 B.n376 VSUBS 0.00864f
C430 B.n377 VSUBS 0.00864f
C431 B.n378 VSUBS 0.00864f
C432 B.n379 VSUBS 0.00864f
C433 B.n380 VSUBS 0.00864f
C434 B.n381 VSUBS 0.00864f
C435 B.n382 VSUBS 0.00864f
C436 B.n383 VSUBS 0.00864f
C437 B.n384 VSUBS 0.00864f
C438 B.n385 VSUBS 0.00864f
C439 B.n386 VSUBS 0.00864f
C440 B.n387 VSUBS 0.00864f
C441 B.n388 VSUBS 0.00864f
C442 B.n389 VSUBS 0.00864f
C443 B.n390 VSUBS 0.00864f
C444 B.n391 VSUBS 0.00864f
C445 B.n392 VSUBS 0.00864f
C446 B.n393 VSUBS 0.00864f
C447 B.n394 VSUBS 0.00864f
C448 B.n395 VSUBS 0.00864f
C449 B.n396 VSUBS 0.00864f
C450 B.n397 VSUBS 0.00864f
C451 B.n398 VSUBS 0.00864f
C452 B.n399 VSUBS 0.00864f
C453 B.n400 VSUBS 0.00864f
C454 B.n401 VSUBS 0.00864f
C455 B.n402 VSUBS 0.00864f
C456 B.n403 VSUBS 0.00864f
C457 B.n404 VSUBS 0.00864f
C458 B.n405 VSUBS 0.00864f
C459 B.n406 VSUBS 0.00864f
C460 B.n407 VSUBS 0.00864f
C461 B.n408 VSUBS 0.00864f
C462 B.n409 VSUBS 0.00864f
C463 B.n410 VSUBS 0.020962f
C464 B.n411 VSUBS 0.019441f
C465 B.n412 VSUBS 0.019441f
C466 B.n413 VSUBS 0.00864f
C467 B.n414 VSUBS 0.00864f
C468 B.n415 VSUBS 0.00864f
C469 B.n416 VSUBS 0.00864f
C470 B.n417 VSUBS 0.00864f
C471 B.n418 VSUBS 0.00864f
C472 B.n419 VSUBS 0.00864f
C473 B.n420 VSUBS 0.00864f
C474 B.n421 VSUBS 0.00864f
C475 B.n422 VSUBS 0.00864f
C476 B.n423 VSUBS 0.00864f
C477 B.n424 VSUBS 0.00864f
C478 B.n425 VSUBS 0.00864f
C479 B.n426 VSUBS 0.00864f
C480 B.n427 VSUBS 0.00864f
C481 B.n428 VSUBS 0.00864f
C482 B.n429 VSUBS 0.00864f
C483 B.n430 VSUBS 0.00864f
C484 B.n431 VSUBS 0.00864f
C485 B.n432 VSUBS 0.00864f
C486 B.n433 VSUBS 0.00864f
C487 B.n434 VSUBS 0.00864f
C488 B.n435 VSUBS 0.00864f
C489 B.n436 VSUBS 0.00864f
C490 B.n437 VSUBS 0.00864f
C491 B.n438 VSUBS 0.00864f
C492 B.n439 VSUBS 0.019563f
C493 VTAIL.n0 VSUBS 0.026804f
C494 VTAIL.n1 VSUBS 0.024206f
C495 VTAIL.n2 VSUBS 0.013007f
C496 VTAIL.n3 VSUBS 0.030744f
C497 VTAIL.n4 VSUBS 0.013772f
C498 VTAIL.n5 VSUBS 0.024206f
C499 VTAIL.n6 VSUBS 0.013007f
C500 VTAIL.n7 VSUBS 0.030744f
C501 VTAIL.n8 VSUBS 0.013772f
C502 VTAIL.n9 VSUBS 0.024206f
C503 VTAIL.n10 VSUBS 0.013007f
C504 VTAIL.n11 VSUBS 0.030744f
C505 VTAIL.n12 VSUBS 0.013772f
C506 VTAIL.n13 VSUBS 0.121303f
C507 VTAIL.t2 VSUBS 0.065553f
C508 VTAIL.n14 VSUBS 0.023058f
C509 VTAIL.n15 VSUBS 0.019558f
C510 VTAIL.n16 VSUBS 0.013007f
C511 VTAIL.n17 VSUBS 0.783766f
C512 VTAIL.n18 VSUBS 0.024206f
C513 VTAIL.n19 VSUBS 0.013007f
C514 VTAIL.n20 VSUBS 0.013772f
C515 VTAIL.n21 VSUBS 0.030744f
C516 VTAIL.n22 VSUBS 0.030744f
C517 VTAIL.n23 VSUBS 0.013772f
C518 VTAIL.n24 VSUBS 0.013007f
C519 VTAIL.n25 VSUBS 0.024206f
C520 VTAIL.n26 VSUBS 0.024206f
C521 VTAIL.n27 VSUBS 0.013007f
C522 VTAIL.n28 VSUBS 0.013772f
C523 VTAIL.n29 VSUBS 0.030744f
C524 VTAIL.n30 VSUBS 0.030744f
C525 VTAIL.n31 VSUBS 0.013772f
C526 VTAIL.n32 VSUBS 0.013007f
C527 VTAIL.n33 VSUBS 0.024206f
C528 VTAIL.n34 VSUBS 0.024206f
C529 VTAIL.n35 VSUBS 0.013007f
C530 VTAIL.n36 VSUBS 0.013772f
C531 VTAIL.n37 VSUBS 0.030744f
C532 VTAIL.n38 VSUBS 0.075132f
C533 VTAIL.n39 VSUBS 0.013772f
C534 VTAIL.n40 VSUBS 0.013007f
C535 VTAIL.n41 VSUBS 0.052975f
C536 VTAIL.n42 VSUBS 0.037721f
C537 VTAIL.n43 VSUBS 0.098506f
C538 VTAIL.n44 VSUBS 0.026804f
C539 VTAIL.n45 VSUBS 0.024206f
C540 VTAIL.n46 VSUBS 0.013007f
C541 VTAIL.n47 VSUBS 0.030744f
C542 VTAIL.n48 VSUBS 0.013772f
C543 VTAIL.n49 VSUBS 0.024206f
C544 VTAIL.n50 VSUBS 0.013007f
C545 VTAIL.n51 VSUBS 0.030744f
C546 VTAIL.n52 VSUBS 0.013772f
C547 VTAIL.n53 VSUBS 0.024206f
C548 VTAIL.n54 VSUBS 0.013007f
C549 VTAIL.n55 VSUBS 0.030744f
C550 VTAIL.n56 VSUBS 0.013772f
C551 VTAIL.n57 VSUBS 0.121303f
C552 VTAIL.t6 VSUBS 0.065553f
C553 VTAIL.n58 VSUBS 0.023058f
C554 VTAIL.n59 VSUBS 0.019558f
C555 VTAIL.n60 VSUBS 0.013007f
C556 VTAIL.n61 VSUBS 0.783766f
C557 VTAIL.n62 VSUBS 0.024206f
C558 VTAIL.n63 VSUBS 0.013007f
C559 VTAIL.n64 VSUBS 0.013772f
C560 VTAIL.n65 VSUBS 0.030744f
C561 VTAIL.n66 VSUBS 0.030744f
C562 VTAIL.n67 VSUBS 0.013772f
C563 VTAIL.n68 VSUBS 0.013007f
C564 VTAIL.n69 VSUBS 0.024206f
C565 VTAIL.n70 VSUBS 0.024206f
C566 VTAIL.n71 VSUBS 0.013007f
C567 VTAIL.n72 VSUBS 0.013772f
C568 VTAIL.n73 VSUBS 0.030744f
C569 VTAIL.n74 VSUBS 0.030744f
C570 VTAIL.n75 VSUBS 0.013772f
C571 VTAIL.n76 VSUBS 0.013007f
C572 VTAIL.n77 VSUBS 0.024206f
C573 VTAIL.n78 VSUBS 0.024206f
C574 VTAIL.n79 VSUBS 0.013007f
C575 VTAIL.n80 VSUBS 0.013772f
C576 VTAIL.n81 VSUBS 0.030744f
C577 VTAIL.n82 VSUBS 0.075132f
C578 VTAIL.n83 VSUBS 0.013772f
C579 VTAIL.n84 VSUBS 0.013007f
C580 VTAIL.n85 VSUBS 0.052975f
C581 VTAIL.n86 VSUBS 0.037721f
C582 VTAIL.n87 VSUBS 0.132293f
C583 VTAIL.n88 VSUBS 0.026804f
C584 VTAIL.n89 VSUBS 0.024206f
C585 VTAIL.n90 VSUBS 0.013007f
C586 VTAIL.n91 VSUBS 0.030744f
C587 VTAIL.n92 VSUBS 0.013772f
C588 VTAIL.n93 VSUBS 0.024206f
C589 VTAIL.n94 VSUBS 0.013007f
C590 VTAIL.n95 VSUBS 0.030744f
C591 VTAIL.n96 VSUBS 0.013772f
C592 VTAIL.n97 VSUBS 0.024206f
C593 VTAIL.n98 VSUBS 0.013007f
C594 VTAIL.n99 VSUBS 0.030744f
C595 VTAIL.n100 VSUBS 0.013772f
C596 VTAIL.n101 VSUBS 0.121303f
C597 VTAIL.t4 VSUBS 0.065553f
C598 VTAIL.n102 VSUBS 0.023058f
C599 VTAIL.n103 VSUBS 0.019558f
C600 VTAIL.n104 VSUBS 0.013007f
C601 VTAIL.n105 VSUBS 0.783766f
C602 VTAIL.n106 VSUBS 0.024206f
C603 VTAIL.n107 VSUBS 0.013007f
C604 VTAIL.n108 VSUBS 0.013772f
C605 VTAIL.n109 VSUBS 0.030744f
C606 VTAIL.n110 VSUBS 0.030744f
C607 VTAIL.n111 VSUBS 0.013772f
C608 VTAIL.n112 VSUBS 0.013007f
C609 VTAIL.n113 VSUBS 0.024206f
C610 VTAIL.n114 VSUBS 0.024206f
C611 VTAIL.n115 VSUBS 0.013007f
C612 VTAIL.n116 VSUBS 0.013772f
C613 VTAIL.n117 VSUBS 0.030744f
C614 VTAIL.n118 VSUBS 0.030744f
C615 VTAIL.n119 VSUBS 0.013772f
C616 VTAIL.n120 VSUBS 0.013007f
C617 VTAIL.n121 VSUBS 0.024206f
C618 VTAIL.n122 VSUBS 0.024206f
C619 VTAIL.n123 VSUBS 0.013007f
C620 VTAIL.n124 VSUBS 0.013772f
C621 VTAIL.n125 VSUBS 0.030744f
C622 VTAIL.n126 VSUBS 0.075132f
C623 VTAIL.n127 VSUBS 0.013772f
C624 VTAIL.n128 VSUBS 0.013007f
C625 VTAIL.n129 VSUBS 0.052975f
C626 VTAIL.n130 VSUBS 0.037721f
C627 VTAIL.n131 VSUBS 1.04372f
C628 VTAIL.n132 VSUBS 0.026804f
C629 VTAIL.n133 VSUBS 0.024206f
C630 VTAIL.n134 VSUBS 0.013007f
C631 VTAIL.n135 VSUBS 0.030744f
C632 VTAIL.n136 VSUBS 0.013772f
C633 VTAIL.n137 VSUBS 0.024206f
C634 VTAIL.n138 VSUBS 0.013007f
C635 VTAIL.n139 VSUBS 0.030744f
C636 VTAIL.n140 VSUBS 0.013772f
C637 VTAIL.n141 VSUBS 0.024206f
C638 VTAIL.n142 VSUBS 0.013007f
C639 VTAIL.n143 VSUBS 0.030744f
C640 VTAIL.n144 VSUBS 0.013772f
C641 VTAIL.n145 VSUBS 0.121303f
C642 VTAIL.t1 VSUBS 0.065553f
C643 VTAIL.n146 VSUBS 0.023058f
C644 VTAIL.n147 VSUBS 0.019558f
C645 VTAIL.n148 VSUBS 0.013007f
C646 VTAIL.n149 VSUBS 0.783766f
C647 VTAIL.n150 VSUBS 0.024206f
C648 VTAIL.n151 VSUBS 0.013007f
C649 VTAIL.n152 VSUBS 0.013772f
C650 VTAIL.n153 VSUBS 0.030744f
C651 VTAIL.n154 VSUBS 0.030744f
C652 VTAIL.n155 VSUBS 0.013772f
C653 VTAIL.n156 VSUBS 0.013007f
C654 VTAIL.n157 VSUBS 0.024206f
C655 VTAIL.n158 VSUBS 0.024206f
C656 VTAIL.n159 VSUBS 0.013007f
C657 VTAIL.n160 VSUBS 0.013772f
C658 VTAIL.n161 VSUBS 0.030744f
C659 VTAIL.n162 VSUBS 0.030744f
C660 VTAIL.n163 VSUBS 0.013772f
C661 VTAIL.n164 VSUBS 0.013007f
C662 VTAIL.n165 VSUBS 0.024206f
C663 VTAIL.n166 VSUBS 0.024206f
C664 VTAIL.n167 VSUBS 0.013007f
C665 VTAIL.n168 VSUBS 0.013772f
C666 VTAIL.n169 VSUBS 0.030744f
C667 VTAIL.n170 VSUBS 0.075132f
C668 VTAIL.n171 VSUBS 0.013772f
C669 VTAIL.n172 VSUBS 0.013007f
C670 VTAIL.n173 VSUBS 0.052975f
C671 VTAIL.n174 VSUBS 0.037721f
C672 VTAIL.n175 VSUBS 1.04372f
C673 VTAIL.n176 VSUBS 0.026804f
C674 VTAIL.n177 VSUBS 0.024206f
C675 VTAIL.n178 VSUBS 0.013007f
C676 VTAIL.n179 VSUBS 0.030744f
C677 VTAIL.n180 VSUBS 0.013772f
C678 VTAIL.n181 VSUBS 0.024206f
C679 VTAIL.n182 VSUBS 0.013007f
C680 VTAIL.n183 VSUBS 0.030744f
C681 VTAIL.n184 VSUBS 0.013772f
C682 VTAIL.n185 VSUBS 0.024206f
C683 VTAIL.n186 VSUBS 0.013007f
C684 VTAIL.n187 VSUBS 0.030744f
C685 VTAIL.n188 VSUBS 0.013772f
C686 VTAIL.n189 VSUBS 0.121303f
C687 VTAIL.t3 VSUBS 0.065553f
C688 VTAIL.n190 VSUBS 0.023058f
C689 VTAIL.n191 VSUBS 0.019558f
C690 VTAIL.n192 VSUBS 0.013007f
C691 VTAIL.n193 VSUBS 0.783766f
C692 VTAIL.n194 VSUBS 0.024206f
C693 VTAIL.n195 VSUBS 0.013007f
C694 VTAIL.n196 VSUBS 0.013772f
C695 VTAIL.n197 VSUBS 0.030744f
C696 VTAIL.n198 VSUBS 0.030744f
C697 VTAIL.n199 VSUBS 0.013772f
C698 VTAIL.n200 VSUBS 0.013007f
C699 VTAIL.n201 VSUBS 0.024206f
C700 VTAIL.n202 VSUBS 0.024206f
C701 VTAIL.n203 VSUBS 0.013007f
C702 VTAIL.n204 VSUBS 0.013772f
C703 VTAIL.n205 VSUBS 0.030744f
C704 VTAIL.n206 VSUBS 0.030744f
C705 VTAIL.n207 VSUBS 0.013772f
C706 VTAIL.n208 VSUBS 0.013007f
C707 VTAIL.n209 VSUBS 0.024206f
C708 VTAIL.n210 VSUBS 0.024206f
C709 VTAIL.n211 VSUBS 0.013007f
C710 VTAIL.n212 VSUBS 0.013772f
C711 VTAIL.n213 VSUBS 0.030744f
C712 VTAIL.n214 VSUBS 0.075132f
C713 VTAIL.n215 VSUBS 0.013772f
C714 VTAIL.n216 VSUBS 0.013007f
C715 VTAIL.n217 VSUBS 0.052975f
C716 VTAIL.n218 VSUBS 0.037721f
C717 VTAIL.n219 VSUBS 0.132293f
C718 VTAIL.n220 VSUBS 0.026804f
C719 VTAIL.n221 VSUBS 0.024206f
C720 VTAIL.n222 VSUBS 0.013007f
C721 VTAIL.n223 VSUBS 0.030744f
C722 VTAIL.n224 VSUBS 0.013772f
C723 VTAIL.n225 VSUBS 0.024206f
C724 VTAIL.n226 VSUBS 0.013007f
C725 VTAIL.n227 VSUBS 0.030744f
C726 VTAIL.n228 VSUBS 0.013772f
C727 VTAIL.n229 VSUBS 0.024206f
C728 VTAIL.n230 VSUBS 0.013007f
C729 VTAIL.n231 VSUBS 0.030744f
C730 VTAIL.n232 VSUBS 0.013772f
C731 VTAIL.n233 VSUBS 0.121303f
C732 VTAIL.t7 VSUBS 0.065553f
C733 VTAIL.n234 VSUBS 0.023058f
C734 VTAIL.n235 VSUBS 0.019558f
C735 VTAIL.n236 VSUBS 0.013007f
C736 VTAIL.n237 VSUBS 0.783766f
C737 VTAIL.n238 VSUBS 0.024206f
C738 VTAIL.n239 VSUBS 0.013007f
C739 VTAIL.n240 VSUBS 0.013772f
C740 VTAIL.n241 VSUBS 0.030744f
C741 VTAIL.n242 VSUBS 0.030744f
C742 VTAIL.n243 VSUBS 0.013772f
C743 VTAIL.n244 VSUBS 0.013007f
C744 VTAIL.n245 VSUBS 0.024206f
C745 VTAIL.n246 VSUBS 0.024206f
C746 VTAIL.n247 VSUBS 0.013007f
C747 VTAIL.n248 VSUBS 0.013772f
C748 VTAIL.n249 VSUBS 0.030744f
C749 VTAIL.n250 VSUBS 0.030744f
C750 VTAIL.n251 VSUBS 0.013772f
C751 VTAIL.n252 VSUBS 0.013007f
C752 VTAIL.n253 VSUBS 0.024206f
C753 VTAIL.n254 VSUBS 0.024206f
C754 VTAIL.n255 VSUBS 0.013007f
C755 VTAIL.n256 VSUBS 0.013772f
C756 VTAIL.n257 VSUBS 0.030744f
C757 VTAIL.n258 VSUBS 0.075132f
C758 VTAIL.n259 VSUBS 0.013772f
C759 VTAIL.n260 VSUBS 0.013007f
C760 VTAIL.n261 VSUBS 0.052975f
C761 VTAIL.n262 VSUBS 0.037721f
C762 VTAIL.n263 VSUBS 0.132293f
C763 VTAIL.n264 VSUBS 0.026804f
C764 VTAIL.n265 VSUBS 0.024206f
C765 VTAIL.n266 VSUBS 0.013007f
C766 VTAIL.n267 VSUBS 0.030744f
C767 VTAIL.n268 VSUBS 0.013772f
C768 VTAIL.n269 VSUBS 0.024206f
C769 VTAIL.n270 VSUBS 0.013007f
C770 VTAIL.n271 VSUBS 0.030744f
C771 VTAIL.n272 VSUBS 0.013772f
C772 VTAIL.n273 VSUBS 0.024206f
C773 VTAIL.n274 VSUBS 0.013007f
C774 VTAIL.n275 VSUBS 0.030744f
C775 VTAIL.n276 VSUBS 0.013772f
C776 VTAIL.n277 VSUBS 0.121303f
C777 VTAIL.t5 VSUBS 0.065553f
C778 VTAIL.n278 VSUBS 0.023058f
C779 VTAIL.n279 VSUBS 0.019558f
C780 VTAIL.n280 VSUBS 0.013007f
C781 VTAIL.n281 VSUBS 0.783766f
C782 VTAIL.n282 VSUBS 0.024206f
C783 VTAIL.n283 VSUBS 0.013007f
C784 VTAIL.n284 VSUBS 0.013772f
C785 VTAIL.n285 VSUBS 0.030744f
C786 VTAIL.n286 VSUBS 0.030744f
C787 VTAIL.n287 VSUBS 0.013772f
C788 VTAIL.n288 VSUBS 0.013007f
C789 VTAIL.n289 VSUBS 0.024206f
C790 VTAIL.n290 VSUBS 0.024206f
C791 VTAIL.n291 VSUBS 0.013007f
C792 VTAIL.n292 VSUBS 0.013772f
C793 VTAIL.n293 VSUBS 0.030744f
C794 VTAIL.n294 VSUBS 0.030744f
C795 VTAIL.n295 VSUBS 0.013772f
C796 VTAIL.n296 VSUBS 0.013007f
C797 VTAIL.n297 VSUBS 0.024206f
C798 VTAIL.n298 VSUBS 0.024206f
C799 VTAIL.n299 VSUBS 0.013007f
C800 VTAIL.n300 VSUBS 0.013772f
C801 VTAIL.n301 VSUBS 0.030744f
C802 VTAIL.n302 VSUBS 0.075132f
C803 VTAIL.n303 VSUBS 0.013772f
C804 VTAIL.n304 VSUBS 0.013007f
C805 VTAIL.n305 VSUBS 0.052975f
C806 VTAIL.n306 VSUBS 0.037721f
C807 VTAIL.n307 VSUBS 1.04372f
C808 VTAIL.n308 VSUBS 0.026804f
C809 VTAIL.n309 VSUBS 0.024206f
C810 VTAIL.n310 VSUBS 0.013007f
C811 VTAIL.n311 VSUBS 0.030744f
C812 VTAIL.n312 VSUBS 0.013772f
C813 VTAIL.n313 VSUBS 0.024206f
C814 VTAIL.n314 VSUBS 0.013007f
C815 VTAIL.n315 VSUBS 0.030744f
C816 VTAIL.n316 VSUBS 0.013772f
C817 VTAIL.n317 VSUBS 0.024206f
C818 VTAIL.n318 VSUBS 0.013007f
C819 VTAIL.n319 VSUBS 0.030744f
C820 VTAIL.n320 VSUBS 0.013772f
C821 VTAIL.n321 VSUBS 0.121303f
C822 VTAIL.t0 VSUBS 0.065553f
C823 VTAIL.n322 VSUBS 0.023058f
C824 VTAIL.n323 VSUBS 0.019558f
C825 VTAIL.n324 VSUBS 0.013007f
C826 VTAIL.n325 VSUBS 0.783766f
C827 VTAIL.n326 VSUBS 0.024206f
C828 VTAIL.n327 VSUBS 0.013007f
C829 VTAIL.n328 VSUBS 0.013772f
C830 VTAIL.n329 VSUBS 0.030744f
C831 VTAIL.n330 VSUBS 0.030744f
C832 VTAIL.n331 VSUBS 0.013772f
C833 VTAIL.n332 VSUBS 0.013007f
C834 VTAIL.n333 VSUBS 0.024206f
C835 VTAIL.n334 VSUBS 0.024206f
C836 VTAIL.n335 VSUBS 0.013007f
C837 VTAIL.n336 VSUBS 0.013772f
C838 VTAIL.n337 VSUBS 0.030744f
C839 VTAIL.n338 VSUBS 0.030744f
C840 VTAIL.n339 VSUBS 0.013772f
C841 VTAIL.n340 VSUBS 0.013007f
C842 VTAIL.n341 VSUBS 0.024206f
C843 VTAIL.n342 VSUBS 0.024206f
C844 VTAIL.n343 VSUBS 0.013007f
C845 VTAIL.n344 VSUBS 0.013772f
C846 VTAIL.n345 VSUBS 0.030744f
C847 VTAIL.n346 VSUBS 0.075132f
C848 VTAIL.n347 VSUBS 0.013772f
C849 VTAIL.n348 VSUBS 0.013007f
C850 VTAIL.n349 VSUBS 0.052975f
C851 VTAIL.n350 VSUBS 0.037721f
C852 VTAIL.n351 VSUBS 1.00086f
C853 VDD1.t1 VSUBS 0.175029f
C854 VDD1.t2 VSUBS 0.175029f
C855 VDD1.n0 VSUBS 1.24661f
C856 VDD1.t0 VSUBS 0.175029f
C857 VDD1.t3 VSUBS 0.175029f
C858 VDD1.n1 VSUBS 1.73521f
C859 VP.n0 VSUBS 0.063185f
C860 VP.t2 VSUBS 1.22244f
C861 VP.t0 VSUBS 1.22253f
C862 VP.n1 VSUBS 2.01835f
C863 VP.n2 VSUBS 3.49489f
C864 VP.t3 VSUBS 1.18808f
C865 VP.n3 VSUBS 0.503699f
C866 VP.n4 VSUBS 0.014338f
C867 VP.t1 VSUBS 1.18808f
C868 VP.n5 VSUBS 0.503699f
C869 VP.n6 VSUBS 0.048966f
.ends

