* NGSPICE file created from diff_pair_sample_0212.ext - technology: sky130A

.subckt diff_pair_sample_0212 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n4520_n3396# sky130_fd_pr__pfet_01v8 ad=4.7346 pd=25.06 as=0 ps=0 w=12.14 l=3.22
X1 VTAIL.t14 VN.t0 VDD2.t4 w_n4520_n3396# sky130_fd_pr__pfet_01v8 ad=2.0031 pd=12.47 as=2.0031 ps=12.47 w=12.14 l=3.22
X2 VDD1.t7 VP.t0 VTAIL.t6 w_n4520_n3396# sky130_fd_pr__pfet_01v8 ad=2.0031 pd=12.47 as=4.7346 ps=25.06 w=12.14 l=3.22
X3 B.t8 B.t6 B.t7 w_n4520_n3396# sky130_fd_pr__pfet_01v8 ad=4.7346 pd=25.06 as=0 ps=0 w=12.14 l=3.22
X4 VTAIL.t4 VP.t1 VDD1.t6 w_n4520_n3396# sky130_fd_pr__pfet_01v8 ad=4.7346 pd=25.06 as=2.0031 ps=12.47 w=12.14 l=3.22
X5 VTAIL.t13 VN.t1 VDD2.t3 w_n4520_n3396# sky130_fd_pr__pfet_01v8 ad=4.7346 pd=25.06 as=2.0031 ps=12.47 w=12.14 l=3.22
X6 VDD2.t7 VN.t2 VTAIL.t12 w_n4520_n3396# sky130_fd_pr__pfet_01v8 ad=2.0031 pd=12.47 as=4.7346 ps=25.06 w=12.14 l=3.22
X7 B.t5 B.t3 B.t4 w_n4520_n3396# sky130_fd_pr__pfet_01v8 ad=4.7346 pd=25.06 as=0 ps=0 w=12.14 l=3.22
X8 VTAIL.t11 VN.t3 VDD2.t6 w_n4520_n3396# sky130_fd_pr__pfet_01v8 ad=4.7346 pd=25.06 as=2.0031 ps=12.47 w=12.14 l=3.22
X9 VTAIL.t5 VP.t2 VDD1.t5 w_n4520_n3396# sky130_fd_pr__pfet_01v8 ad=2.0031 pd=12.47 as=2.0031 ps=12.47 w=12.14 l=3.22
X10 VDD2.t2 VN.t4 VTAIL.t10 w_n4520_n3396# sky130_fd_pr__pfet_01v8 ad=2.0031 pd=12.47 as=2.0031 ps=12.47 w=12.14 l=3.22
X11 VDD1.t4 VP.t3 VTAIL.t3 w_n4520_n3396# sky130_fd_pr__pfet_01v8 ad=2.0031 pd=12.47 as=2.0031 ps=12.47 w=12.14 l=3.22
X12 VDD2.t0 VN.t5 VTAIL.t9 w_n4520_n3396# sky130_fd_pr__pfet_01v8 ad=2.0031 pd=12.47 as=2.0031 ps=12.47 w=12.14 l=3.22
X13 VDD1.t3 VP.t4 VTAIL.t15 w_n4520_n3396# sky130_fd_pr__pfet_01v8 ad=2.0031 pd=12.47 as=4.7346 ps=25.06 w=12.14 l=3.22
X14 VTAIL.t8 VN.t6 VDD2.t5 w_n4520_n3396# sky130_fd_pr__pfet_01v8 ad=2.0031 pd=12.47 as=2.0031 ps=12.47 w=12.14 l=3.22
X15 VDD1.t2 VP.t5 VTAIL.t2 w_n4520_n3396# sky130_fd_pr__pfet_01v8 ad=2.0031 pd=12.47 as=2.0031 ps=12.47 w=12.14 l=3.22
X16 VTAIL.t0 VP.t6 VDD1.t1 w_n4520_n3396# sky130_fd_pr__pfet_01v8 ad=4.7346 pd=25.06 as=2.0031 ps=12.47 w=12.14 l=3.22
X17 B.t2 B.t0 B.t1 w_n4520_n3396# sky130_fd_pr__pfet_01v8 ad=4.7346 pd=25.06 as=0 ps=0 w=12.14 l=3.22
X18 VTAIL.t1 VP.t7 VDD1.t0 w_n4520_n3396# sky130_fd_pr__pfet_01v8 ad=2.0031 pd=12.47 as=2.0031 ps=12.47 w=12.14 l=3.22
X19 VDD2.t1 VN.t7 VTAIL.t7 w_n4520_n3396# sky130_fd_pr__pfet_01v8 ad=2.0031 pd=12.47 as=4.7346 ps=25.06 w=12.14 l=3.22
R0 B.n456 B.n455 585
R1 B.n454 B.n145 585
R2 B.n453 B.n452 585
R3 B.n451 B.n146 585
R4 B.n450 B.n449 585
R5 B.n448 B.n147 585
R6 B.n447 B.n446 585
R7 B.n445 B.n148 585
R8 B.n444 B.n443 585
R9 B.n442 B.n149 585
R10 B.n441 B.n440 585
R11 B.n439 B.n150 585
R12 B.n438 B.n437 585
R13 B.n436 B.n151 585
R14 B.n435 B.n434 585
R15 B.n433 B.n152 585
R16 B.n432 B.n431 585
R17 B.n430 B.n153 585
R18 B.n429 B.n428 585
R19 B.n427 B.n154 585
R20 B.n426 B.n425 585
R21 B.n424 B.n155 585
R22 B.n423 B.n422 585
R23 B.n421 B.n156 585
R24 B.n420 B.n419 585
R25 B.n418 B.n157 585
R26 B.n417 B.n416 585
R27 B.n415 B.n158 585
R28 B.n414 B.n413 585
R29 B.n412 B.n159 585
R30 B.n411 B.n410 585
R31 B.n409 B.n160 585
R32 B.n408 B.n407 585
R33 B.n406 B.n161 585
R34 B.n405 B.n404 585
R35 B.n403 B.n162 585
R36 B.n402 B.n401 585
R37 B.n400 B.n163 585
R38 B.n399 B.n398 585
R39 B.n397 B.n164 585
R40 B.n396 B.n395 585
R41 B.n394 B.n165 585
R42 B.n392 B.n391 585
R43 B.n390 B.n168 585
R44 B.n389 B.n388 585
R45 B.n387 B.n169 585
R46 B.n386 B.n385 585
R47 B.n384 B.n170 585
R48 B.n383 B.n382 585
R49 B.n381 B.n171 585
R50 B.n380 B.n379 585
R51 B.n378 B.n172 585
R52 B.n377 B.n376 585
R53 B.n372 B.n173 585
R54 B.n371 B.n370 585
R55 B.n369 B.n174 585
R56 B.n368 B.n367 585
R57 B.n366 B.n175 585
R58 B.n365 B.n364 585
R59 B.n363 B.n176 585
R60 B.n362 B.n361 585
R61 B.n360 B.n177 585
R62 B.n359 B.n358 585
R63 B.n357 B.n178 585
R64 B.n356 B.n355 585
R65 B.n354 B.n179 585
R66 B.n353 B.n352 585
R67 B.n351 B.n180 585
R68 B.n350 B.n349 585
R69 B.n348 B.n181 585
R70 B.n347 B.n346 585
R71 B.n345 B.n182 585
R72 B.n344 B.n343 585
R73 B.n342 B.n183 585
R74 B.n341 B.n340 585
R75 B.n339 B.n184 585
R76 B.n338 B.n337 585
R77 B.n336 B.n185 585
R78 B.n335 B.n334 585
R79 B.n333 B.n186 585
R80 B.n332 B.n331 585
R81 B.n330 B.n187 585
R82 B.n329 B.n328 585
R83 B.n327 B.n188 585
R84 B.n326 B.n325 585
R85 B.n324 B.n189 585
R86 B.n323 B.n322 585
R87 B.n321 B.n190 585
R88 B.n320 B.n319 585
R89 B.n318 B.n191 585
R90 B.n317 B.n316 585
R91 B.n315 B.n192 585
R92 B.n314 B.n313 585
R93 B.n312 B.n193 585
R94 B.n457 B.n144 585
R95 B.n459 B.n458 585
R96 B.n460 B.n143 585
R97 B.n462 B.n461 585
R98 B.n463 B.n142 585
R99 B.n465 B.n464 585
R100 B.n466 B.n141 585
R101 B.n468 B.n467 585
R102 B.n469 B.n140 585
R103 B.n471 B.n470 585
R104 B.n472 B.n139 585
R105 B.n474 B.n473 585
R106 B.n475 B.n138 585
R107 B.n477 B.n476 585
R108 B.n478 B.n137 585
R109 B.n480 B.n479 585
R110 B.n481 B.n136 585
R111 B.n483 B.n482 585
R112 B.n484 B.n135 585
R113 B.n486 B.n485 585
R114 B.n487 B.n134 585
R115 B.n489 B.n488 585
R116 B.n490 B.n133 585
R117 B.n492 B.n491 585
R118 B.n493 B.n132 585
R119 B.n495 B.n494 585
R120 B.n496 B.n131 585
R121 B.n498 B.n497 585
R122 B.n499 B.n130 585
R123 B.n501 B.n500 585
R124 B.n502 B.n129 585
R125 B.n504 B.n503 585
R126 B.n505 B.n128 585
R127 B.n507 B.n506 585
R128 B.n508 B.n127 585
R129 B.n510 B.n509 585
R130 B.n511 B.n126 585
R131 B.n513 B.n512 585
R132 B.n514 B.n125 585
R133 B.n516 B.n515 585
R134 B.n517 B.n124 585
R135 B.n519 B.n518 585
R136 B.n520 B.n123 585
R137 B.n522 B.n521 585
R138 B.n523 B.n122 585
R139 B.n525 B.n524 585
R140 B.n526 B.n121 585
R141 B.n528 B.n527 585
R142 B.n529 B.n120 585
R143 B.n531 B.n530 585
R144 B.n532 B.n119 585
R145 B.n534 B.n533 585
R146 B.n535 B.n118 585
R147 B.n537 B.n536 585
R148 B.n538 B.n117 585
R149 B.n540 B.n539 585
R150 B.n541 B.n116 585
R151 B.n543 B.n542 585
R152 B.n544 B.n115 585
R153 B.n546 B.n545 585
R154 B.n547 B.n114 585
R155 B.n549 B.n548 585
R156 B.n550 B.n113 585
R157 B.n552 B.n551 585
R158 B.n553 B.n112 585
R159 B.n555 B.n554 585
R160 B.n556 B.n111 585
R161 B.n558 B.n557 585
R162 B.n559 B.n110 585
R163 B.n561 B.n560 585
R164 B.n562 B.n109 585
R165 B.n564 B.n563 585
R166 B.n565 B.n108 585
R167 B.n567 B.n566 585
R168 B.n568 B.n107 585
R169 B.n570 B.n569 585
R170 B.n571 B.n106 585
R171 B.n573 B.n572 585
R172 B.n574 B.n105 585
R173 B.n576 B.n575 585
R174 B.n577 B.n104 585
R175 B.n579 B.n578 585
R176 B.n580 B.n103 585
R177 B.n582 B.n581 585
R178 B.n583 B.n102 585
R179 B.n585 B.n584 585
R180 B.n586 B.n101 585
R181 B.n588 B.n587 585
R182 B.n589 B.n100 585
R183 B.n591 B.n590 585
R184 B.n592 B.n99 585
R185 B.n594 B.n593 585
R186 B.n595 B.n98 585
R187 B.n597 B.n596 585
R188 B.n598 B.n97 585
R189 B.n600 B.n599 585
R190 B.n601 B.n96 585
R191 B.n603 B.n602 585
R192 B.n604 B.n95 585
R193 B.n606 B.n605 585
R194 B.n607 B.n94 585
R195 B.n609 B.n608 585
R196 B.n610 B.n93 585
R197 B.n612 B.n611 585
R198 B.n613 B.n92 585
R199 B.n615 B.n614 585
R200 B.n616 B.n91 585
R201 B.n618 B.n617 585
R202 B.n619 B.n90 585
R203 B.n621 B.n620 585
R204 B.n622 B.n89 585
R205 B.n624 B.n623 585
R206 B.n625 B.n88 585
R207 B.n627 B.n626 585
R208 B.n628 B.n87 585
R209 B.n630 B.n629 585
R210 B.n631 B.n86 585
R211 B.n633 B.n632 585
R212 B.n634 B.n85 585
R213 B.n636 B.n635 585
R214 B.n637 B.n84 585
R215 B.n639 B.n638 585
R216 B.n781 B.n32 585
R217 B.n780 B.n779 585
R218 B.n778 B.n33 585
R219 B.n777 B.n776 585
R220 B.n775 B.n34 585
R221 B.n774 B.n773 585
R222 B.n772 B.n35 585
R223 B.n771 B.n770 585
R224 B.n769 B.n36 585
R225 B.n768 B.n767 585
R226 B.n766 B.n37 585
R227 B.n765 B.n764 585
R228 B.n763 B.n38 585
R229 B.n762 B.n761 585
R230 B.n760 B.n39 585
R231 B.n759 B.n758 585
R232 B.n757 B.n40 585
R233 B.n756 B.n755 585
R234 B.n754 B.n41 585
R235 B.n753 B.n752 585
R236 B.n751 B.n42 585
R237 B.n750 B.n749 585
R238 B.n748 B.n43 585
R239 B.n747 B.n746 585
R240 B.n745 B.n44 585
R241 B.n744 B.n743 585
R242 B.n742 B.n45 585
R243 B.n741 B.n740 585
R244 B.n739 B.n46 585
R245 B.n738 B.n737 585
R246 B.n736 B.n47 585
R247 B.n735 B.n734 585
R248 B.n733 B.n48 585
R249 B.n732 B.n731 585
R250 B.n730 B.n49 585
R251 B.n729 B.n728 585
R252 B.n727 B.n50 585
R253 B.n726 B.n725 585
R254 B.n724 B.n51 585
R255 B.n723 B.n722 585
R256 B.n721 B.n52 585
R257 B.n720 B.n719 585
R258 B.n717 B.n53 585
R259 B.n716 B.n715 585
R260 B.n714 B.n56 585
R261 B.n713 B.n712 585
R262 B.n711 B.n57 585
R263 B.n710 B.n709 585
R264 B.n708 B.n58 585
R265 B.n707 B.n706 585
R266 B.n705 B.n59 585
R267 B.n704 B.n703 585
R268 B.n702 B.n701 585
R269 B.n700 B.n63 585
R270 B.n699 B.n698 585
R271 B.n697 B.n64 585
R272 B.n696 B.n695 585
R273 B.n694 B.n65 585
R274 B.n693 B.n692 585
R275 B.n691 B.n66 585
R276 B.n690 B.n689 585
R277 B.n688 B.n67 585
R278 B.n687 B.n686 585
R279 B.n685 B.n68 585
R280 B.n684 B.n683 585
R281 B.n682 B.n69 585
R282 B.n681 B.n680 585
R283 B.n679 B.n70 585
R284 B.n678 B.n677 585
R285 B.n676 B.n71 585
R286 B.n675 B.n674 585
R287 B.n673 B.n72 585
R288 B.n672 B.n671 585
R289 B.n670 B.n73 585
R290 B.n669 B.n668 585
R291 B.n667 B.n74 585
R292 B.n666 B.n665 585
R293 B.n664 B.n75 585
R294 B.n663 B.n662 585
R295 B.n661 B.n76 585
R296 B.n660 B.n659 585
R297 B.n658 B.n77 585
R298 B.n657 B.n656 585
R299 B.n655 B.n78 585
R300 B.n654 B.n653 585
R301 B.n652 B.n79 585
R302 B.n651 B.n650 585
R303 B.n649 B.n80 585
R304 B.n648 B.n647 585
R305 B.n646 B.n81 585
R306 B.n645 B.n644 585
R307 B.n643 B.n82 585
R308 B.n642 B.n641 585
R309 B.n640 B.n83 585
R310 B.n783 B.n782 585
R311 B.n784 B.n31 585
R312 B.n786 B.n785 585
R313 B.n787 B.n30 585
R314 B.n789 B.n788 585
R315 B.n790 B.n29 585
R316 B.n792 B.n791 585
R317 B.n793 B.n28 585
R318 B.n795 B.n794 585
R319 B.n796 B.n27 585
R320 B.n798 B.n797 585
R321 B.n799 B.n26 585
R322 B.n801 B.n800 585
R323 B.n802 B.n25 585
R324 B.n804 B.n803 585
R325 B.n805 B.n24 585
R326 B.n807 B.n806 585
R327 B.n808 B.n23 585
R328 B.n810 B.n809 585
R329 B.n811 B.n22 585
R330 B.n813 B.n812 585
R331 B.n814 B.n21 585
R332 B.n816 B.n815 585
R333 B.n817 B.n20 585
R334 B.n819 B.n818 585
R335 B.n820 B.n19 585
R336 B.n822 B.n821 585
R337 B.n823 B.n18 585
R338 B.n825 B.n824 585
R339 B.n826 B.n17 585
R340 B.n828 B.n827 585
R341 B.n829 B.n16 585
R342 B.n831 B.n830 585
R343 B.n832 B.n15 585
R344 B.n834 B.n833 585
R345 B.n835 B.n14 585
R346 B.n837 B.n836 585
R347 B.n838 B.n13 585
R348 B.n840 B.n839 585
R349 B.n841 B.n12 585
R350 B.n843 B.n842 585
R351 B.n844 B.n11 585
R352 B.n846 B.n845 585
R353 B.n847 B.n10 585
R354 B.n849 B.n848 585
R355 B.n850 B.n9 585
R356 B.n852 B.n851 585
R357 B.n853 B.n8 585
R358 B.n855 B.n854 585
R359 B.n856 B.n7 585
R360 B.n858 B.n857 585
R361 B.n859 B.n6 585
R362 B.n861 B.n860 585
R363 B.n862 B.n5 585
R364 B.n864 B.n863 585
R365 B.n865 B.n4 585
R366 B.n867 B.n866 585
R367 B.n868 B.n3 585
R368 B.n870 B.n869 585
R369 B.n871 B.n0 585
R370 B.n2 B.n1 585
R371 B.n224 B.n223 585
R372 B.n225 B.n222 585
R373 B.n227 B.n226 585
R374 B.n228 B.n221 585
R375 B.n230 B.n229 585
R376 B.n231 B.n220 585
R377 B.n233 B.n232 585
R378 B.n234 B.n219 585
R379 B.n236 B.n235 585
R380 B.n237 B.n218 585
R381 B.n239 B.n238 585
R382 B.n240 B.n217 585
R383 B.n242 B.n241 585
R384 B.n243 B.n216 585
R385 B.n245 B.n244 585
R386 B.n246 B.n215 585
R387 B.n248 B.n247 585
R388 B.n249 B.n214 585
R389 B.n251 B.n250 585
R390 B.n252 B.n213 585
R391 B.n254 B.n253 585
R392 B.n255 B.n212 585
R393 B.n257 B.n256 585
R394 B.n258 B.n211 585
R395 B.n260 B.n259 585
R396 B.n261 B.n210 585
R397 B.n263 B.n262 585
R398 B.n264 B.n209 585
R399 B.n266 B.n265 585
R400 B.n267 B.n208 585
R401 B.n269 B.n268 585
R402 B.n270 B.n207 585
R403 B.n272 B.n271 585
R404 B.n273 B.n206 585
R405 B.n275 B.n274 585
R406 B.n276 B.n205 585
R407 B.n278 B.n277 585
R408 B.n279 B.n204 585
R409 B.n281 B.n280 585
R410 B.n282 B.n203 585
R411 B.n284 B.n283 585
R412 B.n285 B.n202 585
R413 B.n287 B.n286 585
R414 B.n288 B.n201 585
R415 B.n290 B.n289 585
R416 B.n291 B.n200 585
R417 B.n293 B.n292 585
R418 B.n294 B.n199 585
R419 B.n296 B.n295 585
R420 B.n297 B.n198 585
R421 B.n299 B.n298 585
R422 B.n300 B.n197 585
R423 B.n302 B.n301 585
R424 B.n303 B.n196 585
R425 B.n305 B.n304 585
R426 B.n306 B.n195 585
R427 B.n308 B.n307 585
R428 B.n309 B.n194 585
R429 B.n311 B.n310 585
R430 B.n166 B.t1 447.094
R431 B.n60 B.t8 447.094
R432 B.n373 B.t10 447.094
R433 B.n54 B.t5 447.094
R434 B.n310 B.n193 439.647
R435 B.n457 B.n456 439.647
R436 B.n638 B.n83 439.647
R437 B.n782 B.n781 439.647
R438 B.n167 B.t2 378.245
R439 B.n61 B.t7 378.245
R440 B.n374 B.t11 378.245
R441 B.n55 B.t4 378.245
R442 B.n373 B.t9 299.685
R443 B.n166 B.t0 299.685
R444 B.n60 B.t6 299.685
R445 B.n54 B.t3 299.685
R446 B.n873 B.n872 256.663
R447 B.n872 B.n871 235.042
R448 B.n872 B.n2 235.042
R449 B.n314 B.n193 163.367
R450 B.n315 B.n314 163.367
R451 B.n316 B.n315 163.367
R452 B.n316 B.n191 163.367
R453 B.n320 B.n191 163.367
R454 B.n321 B.n320 163.367
R455 B.n322 B.n321 163.367
R456 B.n322 B.n189 163.367
R457 B.n326 B.n189 163.367
R458 B.n327 B.n326 163.367
R459 B.n328 B.n327 163.367
R460 B.n328 B.n187 163.367
R461 B.n332 B.n187 163.367
R462 B.n333 B.n332 163.367
R463 B.n334 B.n333 163.367
R464 B.n334 B.n185 163.367
R465 B.n338 B.n185 163.367
R466 B.n339 B.n338 163.367
R467 B.n340 B.n339 163.367
R468 B.n340 B.n183 163.367
R469 B.n344 B.n183 163.367
R470 B.n345 B.n344 163.367
R471 B.n346 B.n345 163.367
R472 B.n346 B.n181 163.367
R473 B.n350 B.n181 163.367
R474 B.n351 B.n350 163.367
R475 B.n352 B.n351 163.367
R476 B.n352 B.n179 163.367
R477 B.n356 B.n179 163.367
R478 B.n357 B.n356 163.367
R479 B.n358 B.n357 163.367
R480 B.n358 B.n177 163.367
R481 B.n362 B.n177 163.367
R482 B.n363 B.n362 163.367
R483 B.n364 B.n363 163.367
R484 B.n364 B.n175 163.367
R485 B.n368 B.n175 163.367
R486 B.n369 B.n368 163.367
R487 B.n370 B.n369 163.367
R488 B.n370 B.n173 163.367
R489 B.n377 B.n173 163.367
R490 B.n378 B.n377 163.367
R491 B.n379 B.n378 163.367
R492 B.n379 B.n171 163.367
R493 B.n383 B.n171 163.367
R494 B.n384 B.n383 163.367
R495 B.n385 B.n384 163.367
R496 B.n385 B.n169 163.367
R497 B.n389 B.n169 163.367
R498 B.n390 B.n389 163.367
R499 B.n391 B.n390 163.367
R500 B.n391 B.n165 163.367
R501 B.n396 B.n165 163.367
R502 B.n397 B.n396 163.367
R503 B.n398 B.n397 163.367
R504 B.n398 B.n163 163.367
R505 B.n402 B.n163 163.367
R506 B.n403 B.n402 163.367
R507 B.n404 B.n403 163.367
R508 B.n404 B.n161 163.367
R509 B.n408 B.n161 163.367
R510 B.n409 B.n408 163.367
R511 B.n410 B.n409 163.367
R512 B.n410 B.n159 163.367
R513 B.n414 B.n159 163.367
R514 B.n415 B.n414 163.367
R515 B.n416 B.n415 163.367
R516 B.n416 B.n157 163.367
R517 B.n420 B.n157 163.367
R518 B.n421 B.n420 163.367
R519 B.n422 B.n421 163.367
R520 B.n422 B.n155 163.367
R521 B.n426 B.n155 163.367
R522 B.n427 B.n426 163.367
R523 B.n428 B.n427 163.367
R524 B.n428 B.n153 163.367
R525 B.n432 B.n153 163.367
R526 B.n433 B.n432 163.367
R527 B.n434 B.n433 163.367
R528 B.n434 B.n151 163.367
R529 B.n438 B.n151 163.367
R530 B.n439 B.n438 163.367
R531 B.n440 B.n439 163.367
R532 B.n440 B.n149 163.367
R533 B.n444 B.n149 163.367
R534 B.n445 B.n444 163.367
R535 B.n446 B.n445 163.367
R536 B.n446 B.n147 163.367
R537 B.n450 B.n147 163.367
R538 B.n451 B.n450 163.367
R539 B.n452 B.n451 163.367
R540 B.n452 B.n145 163.367
R541 B.n456 B.n145 163.367
R542 B.n638 B.n637 163.367
R543 B.n637 B.n636 163.367
R544 B.n636 B.n85 163.367
R545 B.n632 B.n85 163.367
R546 B.n632 B.n631 163.367
R547 B.n631 B.n630 163.367
R548 B.n630 B.n87 163.367
R549 B.n626 B.n87 163.367
R550 B.n626 B.n625 163.367
R551 B.n625 B.n624 163.367
R552 B.n624 B.n89 163.367
R553 B.n620 B.n89 163.367
R554 B.n620 B.n619 163.367
R555 B.n619 B.n618 163.367
R556 B.n618 B.n91 163.367
R557 B.n614 B.n91 163.367
R558 B.n614 B.n613 163.367
R559 B.n613 B.n612 163.367
R560 B.n612 B.n93 163.367
R561 B.n608 B.n93 163.367
R562 B.n608 B.n607 163.367
R563 B.n607 B.n606 163.367
R564 B.n606 B.n95 163.367
R565 B.n602 B.n95 163.367
R566 B.n602 B.n601 163.367
R567 B.n601 B.n600 163.367
R568 B.n600 B.n97 163.367
R569 B.n596 B.n97 163.367
R570 B.n596 B.n595 163.367
R571 B.n595 B.n594 163.367
R572 B.n594 B.n99 163.367
R573 B.n590 B.n99 163.367
R574 B.n590 B.n589 163.367
R575 B.n589 B.n588 163.367
R576 B.n588 B.n101 163.367
R577 B.n584 B.n101 163.367
R578 B.n584 B.n583 163.367
R579 B.n583 B.n582 163.367
R580 B.n582 B.n103 163.367
R581 B.n578 B.n103 163.367
R582 B.n578 B.n577 163.367
R583 B.n577 B.n576 163.367
R584 B.n576 B.n105 163.367
R585 B.n572 B.n105 163.367
R586 B.n572 B.n571 163.367
R587 B.n571 B.n570 163.367
R588 B.n570 B.n107 163.367
R589 B.n566 B.n107 163.367
R590 B.n566 B.n565 163.367
R591 B.n565 B.n564 163.367
R592 B.n564 B.n109 163.367
R593 B.n560 B.n109 163.367
R594 B.n560 B.n559 163.367
R595 B.n559 B.n558 163.367
R596 B.n558 B.n111 163.367
R597 B.n554 B.n111 163.367
R598 B.n554 B.n553 163.367
R599 B.n553 B.n552 163.367
R600 B.n552 B.n113 163.367
R601 B.n548 B.n113 163.367
R602 B.n548 B.n547 163.367
R603 B.n547 B.n546 163.367
R604 B.n546 B.n115 163.367
R605 B.n542 B.n115 163.367
R606 B.n542 B.n541 163.367
R607 B.n541 B.n540 163.367
R608 B.n540 B.n117 163.367
R609 B.n536 B.n117 163.367
R610 B.n536 B.n535 163.367
R611 B.n535 B.n534 163.367
R612 B.n534 B.n119 163.367
R613 B.n530 B.n119 163.367
R614 B.n530 B.n529 163.367
R615 B.n529 B.n528 163.367
R616 B.n528 B.n121 163.367
R617 B.n524 B.n121 163.367
R618 B.n524 B.n523 163.367
R619 B.n523 B.n522 163.367
R620 B.n522 B.n123 163.367
R621 B.n518 B.n123 163.367
R622 B.n518 B.n517 163.367
R623 B.n517 B.n516 163.367
R624 B.n516 B.n125 163.367
R625 B.n512 B.n125 163.367
R626 B.n512 B.n511 163.367
R627 B.n511 B.n510 163.367
R628 B.n510 B.n127 163.367
R629 B.n506 B.n127 163.367
R630 B.n506 B.n505 163.367
R631 B.n505 B.n504 163.367
R632 B.n504 B.n129 163.367
R633 B.n500 B.n129 163.367
R634 B.n500 B.n499 163.367
R635 B.n499 B.n498 163.367
R636 B.n498 B.n131 163.367
R637 B.n494 B.n131 163.367
R638 B.n494 B.n493 163.367
R639 B.n493 B.n492 163.367
R640 B.n492 B.n133 163.367
R641 B.n488 B.n133 163.367
R642 B.n488 B.n487 163.367
R643 B.n487 B.n486 163.367
R644 B.n486 B.n135 163.367
R645 B.n482 B.n135 163.367
R646 B.n482 B.n481 163.367
R647 B.n481 B.n480 163.367
R648 B.n480 B.n137 163.367
R649 B.n476 B.n137 163.367
R650 B.n476 B.n475 163.367
R651 B.n475 B.n474 163.367
R652 B.n474 B.n139 163.367
R653 B.n470 B.n139 163.367
R654 B.n470 B.n469 163.367
R655 B.n469 B.n468 163.367
R656 B.n468 B.n141 163.367
R657 B.n464 B.n141 163.367
R658 B.n464 B.n463 163.367
R659 B.n463 B.n462 163.367
R660 B.n462 B.n143 163.367
R661 B.n458 B.n143 163.367
R662 B.n458 B.n457 163.367
R663 B.n781 B.n780 163.367
R664 B.n780 B.n33 163.367
R665 B.n776 B.n33 163.367
R666 B.n776 B.n775 163.367
R667 B.n775 B.n774 163.367
R668 B.n774 B.n35 163.367
R669 B.n770 B.n35 163.367
R670 B.n770 B.n769 163.367
R671 B.n769 B.n768 163.367
R672 B.n768 B.n37 163.367
R673 B.n764 B.n37 163.367
R674 B.n764 B.n763 163.367
R675 B.n763 B.n762 163.367
R676 B.n762 B.n39 163.367
R677 B.n758 B.n39 163.367
R678 B.n758 B.n757 163.367
R679 B.n757 B.n756 163.367
R680 B.n756 B.n41 163.367
R681 B.n752 B.n41 163.367
R682 B.n752 B.n751 163.367
R683 B.n751 B.n750 163.367
R684 B.n750 B.n43 163.367
R685 B.n746 B.n43 163.367
R686 B.n746 B.n745 163.367
R687 B.n745 B.n744 163.367
R688 B.n744 B.n45 163.367
R689 B.n740 B.n45 163.367
R690 B.n740 B.n739 163.367
R691 B.n739 B.n738 163.367
R692 B.n738 B.n47 163.367
R693 B.n734 B.n47 163.367
R694 B.n734 B.n733 163.367
R695 B.n733 B.n732 163.367
R696 B.n732 B.n49 163.367
R697 B.n728 B.n49 163.367
R698 B.n728 B.n727 163.367
R699 B.n727 B.n726 163.367
R700 B.n726 B.n51 163.367
R701 B.n722 B.n51 163.367
R702 B.n722 B.n721 163.367
R703 B.n721 B.n720 163.367
R704 B.n720 B.n53 163.367
R705 B.n715 B.n53 163.367
R706 B.n715 B.n714 163.367
R707 B.n714 B.n713 163.367
R708 B.n713 B.n57 163.367
R709 B.n709 B.n57 163.367
R710 B.n709 B.n708 163.367
R711 B.n708 B.n707 163.367
R712 B.n707 B.n59 163.367
R713 B.n703 B.n59 163.367
R714 B.n703 B.n702 163.367
R715 B.n702 B.n63 163.367
R716 B.n698 B.n63 163.367
R717 B.n698 B.n697 163.367
R718 B.n697 B.n696 163.367
R719 B.n696 B.n65 163.367
R720 B.n692 B.n65 163.367
R721 B.n692 B.n691 163.367
R722 B.n691 B.n690 163.367
R723 B.n690 B.n67 163.367
R724 B.n686 B.n67 163.367
R725 B.n686 B.n685 163.367
R726 B.n685 B.n684 163.367
R727 B.n684 B.n69 163.367
R728 B.n680 B.n69 163.367
R729 B.n680 B.n679 163.367
R730 B.n679 B.n678 163.367
R731 B.n678 B.n71 163.367
R732 B.n674 B.n71 163.367
R733 B.n674 B.n673 163.367
R734 B.n673 B.n672 163.367
R735 B.n672 B.n73 163.367
R736 B.n668 B.n73 163.367
R737 B.n668 B.n667 163.367
R738 B.n667 B.n666 163.367
R739 B.n666 B.n75 163.367
R740 B.n662 B.n75 163.367
R741 B.n662 B.n661 163.367
R742 B.n661 B.n660 163.367
R743 B.n660 B.n77 163.367
R744 B.n656 B.n77 163.367
R745 B.n656 B.n655 163.367
R746 B.n655 B.n654 163.367
R747 B.n654 B.n79 163.367
R748 B.n650 B.n79 163.367
R749 B.n650 B.n649 163.367
R750 B.n649 B.n648 163.367
R751 B.n648 B.n81 163.367
R752 B.n644 B.n81 163.367
R753 B.n644 B.n643 163.367
R754 B.n643 B.n642 163.367
R755 B.n642 B.n83 163.367
R756 B.n782 B.n31 163.367
R757 B.n786 B.n31 163.367
R758 B.n787 B.n786 163.367
R759 B.n788 B.n787 163.367
R760 B.n788 B.n29 163.367
R761 B.n792 B.n29 163.367
R762 B.n793 B.n792 163.367
R763 B.n794 B.n793 163.367
R764 B.n794 B.n27 163.367
R765 B.n798 B.n27 163.367
R766 B.n799 B.n798 163.367
R767 B.n800 B.n799 163.367
R768 B.n800 B.n25 163.367
R769 B.n804 B.n25 163.367
R770 B.n805 B.n804 163.367
R771 B.n806 B.n805 163.367
R772 B.n806 B.n23 163.367
R773 B.n810 B.n23 163.367
R774 B.n811 B.n810 163.367
R775 B.n812 B.n811 163.367
R776 B.n812 B.n21 163.367
R777 B.n816 B.n21 163.367
R778 B.n817 B.n816 163.367
R779 B.n818 B.n817 163.367
R780 B.n818 B.n19 163.367
R781 B.n822 B.n19 163.367
R782 B.n823 B.n822 163.367
R783 B.n824 B.n823 163.367
R784 B.n824 B.n17 163.367
R785 B.n828 B.n17 163.367
R786 B.n829 B.n828 163.367
R787 B.n830 B.n829 163.367
R788 B.n830 B.n15 163.367
R789 B.n834 B.n15 163.367
R790 B.n835 B.n834 163.367
R791 B.n836 B.n835 163.367
R792 B.n836 B.n13 163.367
R793 B.n840 B.n13 163.367
R794 B.n841 B.n840 163.367
R795 B.n842 B.n841 163.367
R796 B.n842 B.n11 163.367
R797 B.n846 B.n11 163.367
R798 B.n847 B.n846 163.367
R799 B.n848 B.n847 163.367
R800 B.n848 B.n9 163.367
R801 B.n852 B.n9 163.367
R802 B.n853 B.n852 163.367
R803 B.n854 B.n853 163.367
R804 B.n854 B.n7 163.367
R805 B.n858 B.n7 163.367
R806 B.n859 B.n858 163.367
R807 B.n860 B.n859 163.367
R808 B.n860 B.n5 163.367
R809 B.n864 B.n5 163.367
R810 B.n865 B.n864 163.367
R811 B.n866 B.n865 163.367
R812 B.n866 B.n3 163.367
R813 B.n870 B.n3 163.367
R814 B.n871 B.n870 163.367
R815 B.n224 B.n2 163.367
R816 B.n225 B.n224 163.367
R817 B.n226 B.n225 163.367
R818 B.n226 B.n221 163.367
R819 B.n230 B.n221 163.367
R820 B.n231 B.n230 163.367
R821 B.n232 B.n231 163.367
R822 B.n232 B.n219 163.367
R823 B.n236 B.n219 163.367
R824 B.n237 B.n236 163.367
R825 B.n238 B.n237 163.367
R826 B.n238 B.n217 163.367
R827 B.n242 B.n217 163.367
R828 B.n243 B.n242 163.367
R829 B.n244 B.n243 163.367
R830 B.n244 B.n215 163.367
R831 B.n248 B.n215 163.367
R832 B.n249 B.n248 163.367
R833 B.n250 B.n249 163.367
R834 B.n250 B.n213 163.367
R835 B.n254 B.n213 163.367
R836 B.n255 B.n254 163.367
R837 B.n256 B.n255 163.367
R838 B.n256 B.n211 163.367
R839 B.n260 B.n211 163.367
R840 B.n261 B.n260 163.367
R841 B.n262 B.n261 163.367
R842 B.n262 B.n209 163.367
R843 B.n266 B.n209 163.367
R844 B.n267 B.n266 163.367
R845 B.n268 B.n267 163.367
R846 B.n268 B.n207 163.367
R847 B.n272 B.n207 163.367
R848 B.n273 B.n272 163.367
R849 B.n274 B.n273 163.367
R850 B.n274 B.n205 163.367
R851 B.n278 B.n205 163.367
R852 B.n279 B.n278 163.367
R853 B.n280 B.n279 163.367
R854 B.n280 B.n203 163.367
R855 B.n284 B.n203 163.367
R856 B.n285 B.n284 163.367
R857 B.n286 B.n285 163.367
R858 B.n286 B.n201 163.367
R859 B.n290 B.n201 163.367
R860 B.n291 B.n290 163.367
R861 B.n292 B.n291 163.367
R862 B.n292 B.n199 163.367
R863 B.n296 B.n199 163.367
R864 B.n297 B.n296 163.367
R865 B.n298 B.n297 163.367
R866 B.n298 B.n197 163.367
R867 B.n302 B.n197 163.367
R868 B.n303 B.n302 163.367
R869 B.n304 B.n303 163.367
R870 B.n304 B.n195 163.367
R871 B.n308 B.n195 163.367
R872 B.n309 B.n308 163.367
R873 B.n310 B.n309 163.367
R874 B.n374 B.n373 68.849
R875 B.n167 B.n166 68.849
R876 B.n61 B.n60 68.849
R877 B.n55 B.n54 68.849
R878 B.n375 B.n374 59.5399
R879 B.n393 B.n167 59.5399
R880 B.n62 B.n61 59.5399
R881 B.n718 B.n55 59.5399
R882 B.n783 B.n32 28.5664
R883 B.n640 B.n639 28.5664
R884 B.n312 B.n311 28.5664
R885 B.n455 B.n144 28.5664
R886 B B.n873 18.0485
R887 B.n784 B.n783 10.6151
R888 B.n785 B.n784 10.6151
R889 B.n785 B.n30 10.6151
R890 B.n789 B.n30 10.6151
R891 B.n790 B.n789 10.6151
R892 B.n791 B.n790 10.6151
R893 B.n791 B.n28 10.6151
R894 B.n795 B.n28 10.6151
R895 B.n796 B.n795 10.6151
R896 B.n797 B.n796 10.6151
R897 B.n797 B.n26 10.6151
R898 B.n801 B.n26 10.6151
R899 B.n802 B.n801 10.6151
R900 B.n803 B.n802 10.6151
R901 B.n803 B.n24 10.6151
R902 B.n807 B.n24 10.6151
R903 B.n808 B.n807 10.6151
R904 B.n809 B.n808 10.6151
R905 B.n809 B.n22 10.6151
R906 B.n813 B.n22 10.6151
R907 B.n814 B.n813 10.6151
R908 B.n815 B.n814 10.6151
R909 B.n815 B.n20 10.6151
R910 B.n819 B.n20 10.6151
R911 B.n820 B.n819 10.6151
R912 B.n821 B.n820 10.6151
R913 B.n821 B.n18 10.6151
R914 B.n825 B.n18 10.6151
R915 B.n826 B.n825 10.6151
R916 B.n827 B.n826 10.6151
R917 B.n827 B.n16 10.6151
R918 B.n831 B.n16 10.6151
R919 B.n832 B.n831 10.6151
R920 B.n833 B.n832 10.6151
R921 B.n833 B.n14 10.6151
R922 B.n837 B.n14 10.6151
R923 B.n838 B.n837 10.6151
R924 B.n839 B.n838 10.6151
R925 B.n839 B.n12 10.6151
R926 B.n843 B.n12 10.6151
R927 B.n844 B.n843 10.6151
R928 B.n845 B.n844 10.6151
R929 B.n845 B.n10 10.6151
R930 B.n849 B.n10 10.6151
R931 B.n850 B.n849 10.6151
R932 B.n851 B.n850 10.6151
R933 B.n851 B.n8 10.6151
R934 B.n855 B.n8 10.6151
R935 B.n856 B.n855 10.6151
R936 B.n857 B.n856 10.6151
R937 B.n857 B.n6 10.6151
R938 B.n861 B.n6 10.6151
R939 B.n862 B.n861 10.6151
R940 B.n863 B.n862 10.6151
R941 B.n863 B.n4 10.6151
R942 B.n867 B.n4 10.6151
R943 B.n868 B.n867 10.6151
R944 B.n869 B.n868 10.6151
R945 B.n869 B.n0 10.6151
R946 B.n779 B.n32 10.6151
R947 B.n779 B.n778 10.6151
R948 B.n778 B.n777 10.6151
R949 B.n777 B.n34 10.6151
R950 B.n773 B.n34 10.6151
R951 B.n773 B.n772 10.6151
R952 B.n772 B.n771 10.6151
R953 B.n771 B.n36 10.6151
R954 B.n767 B.n36 10.6151
R955 B.n767 B.n766 10.6151
R956 B.n766 B.n765 10.6151
R957 B.n765 B.n38 10.6151
R958 B.n761 B.n38 10.6151
R959 B.n761 B.n760 10.6151
R960 B.n760 B.n759 10.6151
R961 B.n759 B.n40 10.6151
R962 B.n755 B.n40 10.6151
R963 B.n755 B.n754 10.6151
R964 B.n754 B.n753 10.6151
R965 B.n753 B.n42 10.6151
R966 B.n749 B.n42 10.6151
R967 B.n749 B.n748 10.6151
R968 B.n748 B.n747 10.6151
R969 B.n747 B.n44 10.6151
R970 B.n743 B.n44 10.6151
R971 B.n743 B.n742 10.6151
R972 B.n742 B.n741 10.6151
R973 B.n741 B.n46 10.6151
R974 B.n737 B.n46 10.6151
R975 B.n737 B.n736 10.6151
R976 B.n736 B.n735 10.6151
R977 B.n735 B.n48 10.6151
R978 B.n731 B.n48 10.6151
R979 B.n731 B.n730 10.6151
R980 B.n730 B.n729 10.6151
R981 B.n729 B.n50 10.6151
R982 B.n725 B.n50 10.6151
R983 B.n725 B.n724 10.6151
R984 B.n724 B.n723 10.6151
R985 B.n723 B.n52 10.6151
R986 B.n719 B.n52 10.6151
R987 B.n717 B.n716 10.6151
R988 B.n716 B.n56 10.6151
R989 B.n712 B.n56 10.6151
R990 B.n712 B.n711 10.6151
R991 B.n711 B.n710 10.6151
R992 B.n710 B.n58 10.6151
R993 B.n706 B.n58 10.6151
R994 B.n706 B.n705 10.6151
R995 B.n705 B.n704 10.6151
R996 B.n701 B.n700 10.6151
R997 B.n700 B.n699 10.6151
R998 B.n699 B.n64 10.6151
R999 B.n695 B.n64 10.6151
R1000 B.n695 B.n694 10.6151
R1001 B.n694 B.n693 10.6151
R1002 B.n693 B.n66 10.6151
R1003 B.n689 B.n66 10.6151
R1004 B.n689 B.n688 10.6151
R1005 B.n688 B.n687 10.6151
R1006 B.n687 B.n68 10.6151
R1007 B.n683 B.n68 10.6151
R1008 B.n683 B.n682 10.6151
R1009 B.n682 B.n681 10.6151
R1010 B.n681 B.n70 10.6151
R1011 B.n677 B.n70 10.6151
R1012 B.n677 B.n676 10.6151
R1013 B.n676 B.n675 10.6151
R1014 B.n675 B.n72 10.6151
R1015 B.n671 B.n72 10.6151
R1016 B.n671 B.n670 10.6151
R1017 B.n670 B.n669 10.6151
R1018 B.n669 B.n74 10.6151
R1019 B.n665 B.n74 10.6151
R1020 B.n665 B.n664 10.6151
R1021 B.n664 B.n663 10.6151
R1022 B.n663 B.n76 10.6151
R1023 B.n659 B.n76 10.6151
R1024 B.n659 B.n658 10.6151
R1025 B.n658 B.n657 10.6151
R1026 B.n657 B.n78 10.6151
R1027 B.n653 B.n78 10.6151
R1028 B.n653 B.n652 10.6151
R1029 B.n652 B.n651 10.6151
R1030 B.n651 B.n80 10.6151
R1031 B.n647 B.n80 10.6151
R1032 B.n647 B.n646 10.6151
R1033 B.n646 B.n645 10.6151
R1034 B.n645 B.n82 10.6151
R1035 B.n641 B.n82 10.6151
R1036 B.n641 B.n640 10.6151
R1037 B.n639 B.n84 10.6151
R1038 B.n635 B.n84 10.6151
R1039 B.n635 B.n634 10.6151
R1040 B.n634 B.n633 10.6151
R1041 B.n633 B.n86 10.6151
R1042 B.n629 B.n86 10.6151
R1043 B.n629 B.n628 10.6151
R1044 B.n628 B.n627 10.6151
R1045 B.n627 B.n88 10.6151
R1046 B.n623 B.n88 10.6151
R1047 B.n623 B.n622 10.6151
R1048 B.n622 B.n621 10.6151
R1049 B.n621 B.n90 10.6151
R1050 B.n617 B.n90 10.6151
R1051 B.n617 B.n616 10.6151
R1052 B.n616 B.n615 10.6151
R1053 B.n615 B.n92 10.6151
R1054 B.n611 B.n92 10.6151
R1055 B.n611 B.n610 10.6151
R1056 B.n610 B.n609 10.6151
R1057 B.n609 B.n94 10.6151
R1058 B.n605 B.n94 10.6151
R1059 B.n605 B.n604 10.6151
R1060 B.n604 B.n603 10.6151
R1061 B.n603 B.n96 10.6151
R1062 B.n599 B.n96 10.6151
R1063 B.n599 B.n598 10.6151
R1064 B.n598 B.n597 10.6151
R1065 B.n597 B.n98 10.6151
R1066 B.n593 B.n98 10.6151
R1067 B.n593 B.n592 10.6151
R1068 B.n592 B.n591 10.6151
R1069 B.n591 B.n100 10.6151
R1070 B.n587 B.n100 10.6151
R1071 B.n587 B.n586 10.6151
R1072 B.n586 B.n585 10.6151
R1073 B.n585 B.n102 10.6151
R1074 B.n581 B.n102 10.6151
R1075 B.n581 B.n580 10.6151
R1076 B.n580 B.n579 10.6151
R1077 B.n579 B.n104 10.6151
R1078 B.n575 B.n104 10.6151
R1079 B.n575 B.n574 10.6151
R1080 B.n574 B.n573 10.6151
R1081 B.n573 B.n106 10.6151
R1082 B.n569 B.n106 10.6151
R1083 B.n569 B.n568 10.6151
R1084 B.n568 B.n567 10.6151
R1085 B.n567 B.n108 10.6151
R1086 B.n563 B.n108 10.6151
R1087 B.n563 B.n562 10.6151
R1088 B.n562 B.n561 10.6151
R1089 B.n561 B.n110 10.6151
R1090 B.n557 B.n110 10.6151
R1091 B.n557 B.n556 10.6151
R1092 B.n556 B.n555 10.6151
R1093 B.n555 B.n112 10.6151
R1094 B.n551 B.n112 10.6151
R1095 B.n551 B.n550 10.6151
R1096 B.n550 B.n549 10.6151
R1097 B.n549 B.n114 10.6151
R1098 B.n545 B.n114 10.6151
R1099 B.n545 B.n544 10.6151
R1100 B.n544 B.n543 10.6151
R1101 B.n543 B.n116 10.6151
R1102 B.n539 B.n116 10.6151
R1103 B.n539 B.n538 10.6151
R1104 B.n538 B.n537 10.6151
R1105 B.n537 B.n118 10.6151
R1106 B.n533 B.n118 10.6151
R1107 B.n533 B.n532 10.6151
R1108 B.n532 B.n531 10.6151
R1109 B.n531 B.n120 10.6151
R1110 B.n527 B.n120 10.6151
R1111 B.n527 B.n526 10.6151
R1112 B.n526 B.n525 10.6151
R1113 B.n525 B.n122 10.6151
R1114 B.n521 B.n122 10.6151
R1115 B.n521 B.n520 10.6151
R1116 B.n520 B.n519 10.6151
R1117 B.n519 B.n124 10.6151
R1118 B.n515 B.n124 10.6151
R1119 B.n515 B.n514 10.6151
R1120 B.n514 B.n513 10.6151
R1121 B.n513 B.n126 10.6151
R1122 B.n509 B.n126 10.6151
R1123 B.n509 B.n508 10.6151
R1124 B.n508 B.n507 10.6151
R1125 B.n507 B.n128 10.6151
R1126 B.n503 B.n128 10.6151
R1127 B.n503 B.n502 10.6151
R1128 B.n502 B.n501 10.6151
R1129 B.n501 B.n130 10.6151
R1130 B.n497 B.n130 10.6151
R1131 B.n497 B.n496 10.6151
R1132 B.n496 B.n495 10.6151
R1133 B.n495 B.n132 10.6151
R1134 B.n491 B.n132 10.6151
R1135 B.n491 B.n490 10.6151
R1136 B.n490 B.n489 10.6151
R1137 B.n489 B.n134 10.6151
R1138 B.n485 B.n134 10.6151
R1139 B.n485 B.n484 10.6151
R1140 B.n484 B.n483 10.6151
R1141 B.n483 B.n136 10.6151
R1142 B.n479 B.n136 10.6151
R1143 B.n479 B.n478 10.6151
R1144 B.n478 B.n477 10.6151
R1145 B.n477 B.n138 10.6151
R1146 B.n473 B.n138 10.6151
R1147 B.n473 B.n472 10.6151
R1148 B.n472 B.n471 10.6151
R1149 B.n471 B.n140 10.6151
R1150 B.n467 B.n140 10.6151
R1151 B.n467 B.n466 10.6151
R1152 B.n466 B.n465 10.6151
R1153 B.n465 B.n142 10.6151
R1154 B.n461 B.n142 10.6151
R1155 B.n461 B.n460 10.6151
R1156 B.n460 B.n459 10.6151
R1157 B.n459 B.n144 10.6151
R1158 B.n223 B.n1 10.6151
R1159 B.n223 B.n222 10.6151
R1160 B.n227 B.n222 10.6151
R1161 B.n228 B.n227 10.6151
R1162 B.n229 B.n228 10.6151
R1163 B.n229 B.n220 10.6151
R1164 B.n233 B.n220 10.6151
R1165 B.n234 B.n233 10.6151
R1166 B.n235 B.n234 10.6151
R1167 B.n235 B.n218 10.6151
R1168 B.n239 B.n218 10.6151
R1169 B.n240 B.n239 10.6151
R1170 B.n241 B.n240 10.6151
R1171 B.n241 B.n216 10.6151
R1172 B.n245 B.n216 10.6151
R1173 B.n246 B.n245 10.6151
R1174 B.n247 B.n246 10.6151
R1175 B.n247 B.n214 10.6151
R1176 B.n251 B.n214 10.6151
R1177 B.n252 B.n251 10.6151
R1178 B.n253 B.n252 10.6151
R1179 B.n253 B.n212 10.6151
R1180 B.n257 B.n212 10.6151
R1181 B.n258 B.n257 10.6151
R1182 B.n259 B.n258 10.6151
R1183 B.n259 B.n210 10.6151
R1184 B.n263 B.n210 10.6151
R1185 B.n264 B.n263 10.6151
R1186 B.n265 B.n264 10.6151
R1187 B.n265 B.n208 10.6151
R1188 B.n269 B.n208 10.6151
R1189 B.n270 B.n269 10.6151
R1190 B.n271 B.n270 10.6151
R1191 B.n271 B.n206 10.6151
R1192 B.n275 B.n206 10.6151
R1193 B.n276 B.n275 10.6151
R1194 B.n277 B.n276 10.6151
R1195 B.n277 B.n204 10.6151
R1196 B.n281 B.n204 10.6151
R1197 B.n282 B.n281 10.6151
R1198 B.n283 B.n282 10.6151
R1199 B.n283 B.n202 10.6151
R1200 B.n287 B.n202 10.6151
R1201 B.n288 B.n287 10.6151
R1202 B.n289 B.n288 10.6151
R1203 B.n289 B.n200 10.6151
R1204 B.n293 B.n200 10.6151
R1205 B.n294 B.n293 10.6151
R1206 B.n295 B.n294 10.6151
R1207 B.n295 B.n198 10.6151
R1208 B.n299 B.n198 10.6151
R1209 B.n300 B.n299 10.6151
R1210 B.n301 B.n300 10.6151
R1211 B.n301 B.n196 10.6151
R1212 B.n305 B.n196 10.6151
R1213 B.n306 B.n305 10.6151
R1214 B.n307 B.n306 10.6151
R1215 B.n307 B.n194 10.6151
R1216 B.n311 B.n194 10.6151
R1217 B.n313 B.n312 10.6151
R1218 B.n313 B.n192 10.6151
R1219 B.n317 B.n192 10.6151
R1220 B.n318 B.n317 10.6151
R1221 B.n319 B.n318 10.6151
R1222 B.n319 B.n190 10.6151
R1223 B.n323 B.n190 10.6151
R1224 B.n324 B.n323 10.6151
R1225 B.n325 B.n324 10.6151
R1226 B.n325 B.n188 10.6151
R1227 B.n329 B.n188 10.6151
R1228 B.n330 B.n329 10.6151
R1229 B.n331 B.n330 10.6151
R1230 B.n331 B.n186 10.6151
R1231 B.n335 B.n186 10.6151
R1232 B.n336 B.n335 10.6151
R1233 B.n337 B.n336 10.6151
R1234 B.n337 B.n184 10.6151
R1235 B.n341 B.n184 10.6151
R1236 B.n342 B.n341 10.6151
R1237 B.n343 B.n342 10.6151
R1238 B.n343 B.n182 10.6151
R1239 B.n347 B.n182 10.6151
R1240 B.n348 B.n347 10.6151
R1241 B.n349 B.n348 10.6151
R1242 B.n349 B.n180 10.6151
R1243 B.n353 B.n180 10.6151
R1244 B.n354 B.n353 10.6151
R1245 B.n355 B.n354 10.6151
R1246 B.n355 B.n178 10.6151
R1247 B.n359 B.n178 10.6151
R1248 B.n360 B.n359 10.6151
R1249 B.n361 B.n360 10.6151
R1250 B.n361 B.n176 10.6151
R1251 B.n365 B.n176 10.6151
R1252 B.n366 B.n365 10.6151
R1253 B.n367 B.n366 10.6151
R1254 B.n367 B.n174 10.6151
R1255 B.n371 B.n174 10.6151
R1256 B.n372 B.n371 10.6151
R1257 B.n376 B.n372 10.6151
R1258 B.n380 B.n172 10.6151
R1259 B.n381 B.n380 10.6151
R1260 B.n382 B.n381 10.6151
R1261 B.n382 B.n170 10.6151
R1262 B.n386 B.n170 10.6151
R1263 B.n387 B.n386 10.6151
R1264 B.n388 B.n387 10.6151
R1265 B.n388 B.n168 10.6151
R1266 B.n392 B.n168 10.6151
R1267 B.n395 B.n394 10.6151
R1268 B.n395 B.n164 10.6151
R1269 B.n399 B.n164 10.6151
R1270 B.n400 B.n399 10.6151
R1271 B.n401 B.n400 10.6151
R1272 B.n401 B.n162 10.6151
R1273 B.n405 B.n162 10.6151
R1274 B.n406 B.n405 10.6151
R1275 B.n407 B.n406 10.6151
R1276 B.n407 B.n160 10.6151
R1277 B.n411 B.n160 10.6151
R1278 B.n412 B.n411 10.6151
R1279 B.n413 B.n412 10.6151
R1280 B.n413 B.n158 10.6151
R1281 B.n417 B.n158 10.6151
R1282 B.n418 B.n417 10.6151
R1283 B.n419 B.n418 10.6151
R1284 B.n419 B.n156 10.6151
R1285 B.n423 B.n156 10.6151
R1286 B.n424 B.n423 10.6151
R1287 B.n425 B.n424 10.6151
R1288 B.n425 B.n154 10.6151
R1289 B.n429 B.n154 10.6151
R1290 B.n430 B.n429 10.6151
R1291 B.n431 B.n430 10.6151
R1292 B.n431 B.n152 10.6151
R1293 B.n435 B.n152 10.6151
R1294 B.n436 B.n435 10.6151
R1295 B.n437 B.n436 10.6151
R1296 B.n437 B.n150 10.6151
R1297 B.n441 B.n150 10.6151
R1298 B.n442 B.n441 10.6151
R1299 B.n443 B.n442 10.6151
R1300 B.n443 B.n148 10.6151
R1301 B.n447 B.n148 10.6151
R1302 B.n448 B.n447 10.6151
R1303 B.n449 B.n448 10.6151
R1304 B.n449 B.n146 10.6151
R1305 B.n453 B.n146 10.6151
R1306 B.n454 B.n453 10.6151
R1307 B.n455 B.n454 10.6151
R1308 B.n719 B.n718 9.36635
R1309 B.n701 B.n62 9.36635
R1310 B.n376 B.n375 9.36635
R1311 B.n394 B.n393 9.36635
R1312 B.n873 B.n0 8.11757
R1313 B.n873 B.n1 8.11757
R1314 B.n718 B.n717 1.24928
R1315 B.n704 B.n62 1.24928
R1316 B.n375 B.n172 1.24928
R1317 B.n393 B.n392 1.24928
R1318 VN.n64 VN.n63 161.3
R1319 VN.n62 VN.n34 161.3
R1320 VN.n61 VN.n60 161.3
R1321 VN.n59 VN.n35 161.3
R1322 VN.n58 VN.n57 161.3
R1323 VN.n56 VN.n36 161.3
R1324 VN.n55 VN.n54 161.3
R1325 VN.n53 VN.n52 161.3
R1326 VN.n51 VN.n38 161.3
R1327 VN.n50 VN.n49 161.3
R1328 VN.n48 VN.n39 161.3
R1329 VN.n47 VN.n46 161.3
R1330 VN.n45 VN.n40 161.3
R1331 VN.n44 VN.n43 161.3
R1332 VN.n31 VN.n30 161.3
R1333 VN.n29 VN.n1 161.3
R1334 VN.n28 VN.n27 161.3
R1335 VN.n26 VN.n2 161.3
R1336 VN.n25 VN.n24 161.3
R1337 VN.n23 VN.n3 161.3
R1338 VN.n22 VN.n21 161.3
R1339 VN.n20 VN.n19 161.3
R1340 VN.n18 VN.n5 161.3
R1341 VN.n17 VN.n16 161.3
R1342 VN.n15 VN.n6 161.3
R1343 VN.n14 VN.n13 161.3
R1344 VN.n12 VN.n7 161.3
R1345 VN.n11 VN.n10 161.3
R1346 VN.n42 VN.t2 123.871
R1347 VN.n9 VN.t3 123.871
R1348 VN.n8 VN.t4 90.862
R1349 VN.n4 VN.t6 90.862
R1350 VN.n0 VN.t7 90.862
R1351 VN.n41 VN.t0 90.862
R1352 VN.n37 VN.t5 90.862
R1353 VN.n33 VN.t1 90.862
R1354 VN.n32 VN.n0 74.0678
R1355 VN.n65 VN.n33 74.0678
R1356 VN.n9 VN.n8 60.6108
R1357 VN.n42 VN.n41 60.6108
R1358 VN VN.n65 54.1797
R1359 VN.n28 VN.n2 45.2793
R1360 VN.n61 VN.n35 45.2793
R1361 VN.n13 VN.n6 40.4106
R1362 VN.n17 VN.n6 40.4106
R1363 VN.n46 VN.n39 40.4106
R1364 VN.n50 VN.n39 40.4106
R1365 VN.n24 VN.n2 35.5419
R1366 VN.n57 VN.n35 35.5419
R1367 VN.n12 VN.n11 24.3439
R1368 VN.n13 VN.n12 24.3439
R1369 VN.n18 VN.n17 24.3439
R1370 VN.n19 VN.n18 24.3439
R1371 VN.n23 VN.n22 24.3439
R1372 VN.n24 VN.n23 24.3439
R1373 VN.n29 VN.n28 24.3439
R1374 VN.n30 VN.n29 24.3439
R1375 VN.n46 VN.n45 24.3439
R1376 VN.n45 VN.n44 24.3439
R1377 VN.n57 VN.n56 24.3439
R1378 VN.n56 VN.n55 24.3439
R1379 VN.n52 VN.n51 24.3439
R1380 VN.n51 VN.n50 24.3439
R1381 VN.n63 VN.n62 24.3439
R1382 VN.n62 VN.n61 24.3439
R1383 VN.n30 VN.n0 15.8237
R1384 VN.n63 VN.n33 15.8237
R1385 VN.n11 VN.n8 13.3894
R1386 VN.n19 VN.n4 13.3894
R1387 VN.n44 VN.n41 13.3894
R1388 VN.n52 VN.n37 13.3894
R1389 VN.n22 VN.n4 10.955
R1390 VN.n55 VN.n37 10.955
R1391 VN.n43 VN.n42 4.11425
R1392 VN.n10 VN.n9 4.11425
R1393 VN.n65 VN.n64 0.355081
R1394 VN.n32 VN.n31 0.355081
R1395 VN VN.n32 0.26685
R1396 VN.n64 VN.n34 0.189894
R1397 VN.n60 VN.n34 0.189894
R1398 VN.n60 VN.n59 0.189894
R1399 VN.n59 VN.n58 0.189894
R1400 VN.n58 VN.n36 0.189894
R1401 VN.n54 VN.n36 0.189894
R1402 VN.n54 VN.n53 0.189894
R1403 VN.n53 VN.n38 0.189894
R1404 VN.n49 VN.n38 0.189894
R1405 VN.n49 VN.n48 0.189894
R1406 VN.n48 VN.n47 0.189894
R1407 VN.n47 VN.n40 0.189894
R1408 VN.n43 VN.n40 0.189894
R1409 VN.n10 VN.n7 0.189894
R1410 VN.n14 VN.n7 0.189894
R1411 VN.n15 VN.n14 0.189894
R1412 VN.n16 VN.n15 0.189894
R1413 VN.n16 VN.n5 0.189894
R1414 VN.n20 VN.n5 0.189894
R1415 VN.n21 VN.n20 0.189894
R1416 VN.n21 VN.n3 0.189894
R1417 VN.n25 VN.n3 0.189894
R1418 VN.n26 VN.n25 0.189894
R1419 VN.n27 VN.n26 0.189894
R1420 VN.n27 VN.n1 0.189894
R1421 VN.n31 VN.n1 0.189894
R1422 VDD2.n2 VDD2.n1 75.7017
R1423 VDD2.n2 VDD2.n0 75.7017
R1424 VDD2 VDD2.n5 75.6989
R1425 VDD2.n4 VDD2.n3 74.2271
R1426 VDD2.n4 VDD2.n2 47.9524
R1427 VDD2.n5 VDD2.t4 2.67801
R1428 VDD2.n5 VDD2.t7 2.67801
R1429 VDD2.n3 VDD2.t3 2.67801
R1430 VDD2.n3 VDD2.t0 2.67801
R1431 VDD2.n1 VDD2.t5 2.67801
R1432 VDD2.n1 VDD2.t1 2.67801
R1433 VDD2.n0 VDD2.t6 2.67801
R1434 VDD2.n0 VDD2.t2 2.67801
R1435 VDD2 VDD2.n4 1.58886
R1436 VTAIL.n530 VTAIL.n470 756.745
R1437 VTAIL.n62 VTAIL.n2 756.745
R1438 VTAIL.n128 VTAIL.n68 756.745
R1439 VTAIL.n196 VTAIL.n136 756.745
R1440 VTAIL.n464 VTAIL.n404 756.745
R1441 VTAIL.n396 VTAIL.n336 756.745
R1442 VTAIL.n330 VTAIL.n270 756.745
R1443 VTAIL.n262 VTAIL.n202 756.745
R1444 VTAIL.n490 VTAIL.n489 585
R1445 VTAIL.n495 VTAIL.n494 585
R1446 VTAIL.n497 VTAIL.n496 585
R1447 VTAIL.n486 VTAIL.n485 585
R1448 VTAIL.n503 VTAIL.n502 585
R1449 VTAIL.n505 VTAIL.n504 585
R1450 VTAIL.n482 VTAIL.n481 585
R1451 VTAIL.n512 VTAIL.n511 585
R1452 VTAIL.n513 VTAIL.n480 585
R1453 VTAIL.n515 VTAIL.n514 585
R1454 VTAIL.n478 VTAIL.n477 585
R1455 VTAIL.n521 VTAIL.n520 585
R1456 VTAIL.n523 VTAIL.n522 585
R1457 VTAIL.n474 VTAIL.n473 585
R1458 VTAIL.n529 VTAIL.n528 585
R1459 VTAIL.n531 VTAIL.n530 585
R1460 VTAIL.n22 VTAIL.n21 585
R1461 VTAIL.n27 VTAIL.n26 585
R1462 VTAIL.n29 VTAIL.n28 585
R1463 VTAIL.n18 VTAIL.n17 585
R1464 VTAIL.n35 VTAIL.n34 585
R1465 VTAIL.n37 VTAIL.n36 585
R1466 VTAIL.n14 VTAIL.n13 585
R1467 VTAIL.n44 VTAIL.n43 585
R1468 VTAIL.n45 VTAIL.n12 585
R1469 VTAIL.n47 VTAIL.n46 585
R1470 VTAIL.n10 VTAIL.n9 585
R1471 VTAIL.n53 VTAIL.n52 585
R1472 VTAIL.n55 VTAIL.n54 585
R1473 VTAIL.n6 VTAIL.n5 585
R1474 VTAIL.n61 VTAIL.n60 585
R1475 VTAIL.n63 VTAIL.n62 585
R1476 VTAIL.n88 VTAIL.n87 585
R1477 VTAIL.n93 VTAIL.n92 585
R1478 VTAIL.n95 VTAIL.n94 585
R1479 VTAIL.n84 VTAIL.n83 585
R1480 VTAIL.n101 VTAIL.n100 585
R1481 VTAIL.n103 VTAIL.n102 585
R1482 VTAIL.n80 VTAIL.n79 585
R1483 VTAIL.n110 VTAIL.n109 585
R1484 VTAIL.n111 VTAIL.n78 585
R1485 VTAIL.n113 VTAIL.n112 585
R1486 VTAIL.n76 VTAIL.n75 585
R1487 VTAIL.n119 VTAIL.n118 585
R1488 VTAIL.n121 VTAIL.n120 585
R1489 VTAIL.n72 VTAIL.n71 585
R1490 VTAIL.n127 VTAIL.n126 585
R1491 VTAIL.n129 VTAIL.n128 585
R1492 VTAIL.n156 VTAIL.n155 585
R1493 VTAIL.n161 VTAIL.n160 585
R1494 VTAIL.n163 VTAIL.n162 585
R1495 VTAIL.n152 VTAIL.n151 585
R1496 VTAIL.n169 VTAIL.n168 585
R1497 VTAIL.n171 VTAIL.n170 585
R1498 VTAIL.n148 VTAIL.n147 585
R1499 VTAIL.n178 VTAIL.n177 585
R1500 VTAIL.n179 VTAIL.n146 585
R1501 VTAIL.n181 VTAIL.n180 585
R1502 VTAIL.n144 VTAIL.n143 585
R1503 VTAIL.n187 VTAIL.n186 585
R1504 VTAIL.n189 VTAIL.n188 585
R1505 VTAIL.n140 VTAIL.n139 585
R1506 VTAIL.n195 VTAIL.n194 585
R1507 VTAIL.n197 VTAIL.n196 585
R1508 VTAIL.n465 VTAIL.n464 585
R1509 VTAIL.n463 VTAIL.n462 585
R1510 VTAIL.n408 VTAIL.n407 585
R1511 VTAIL.n457 VTAIL.n456 585
R1512 VTAIL.n455 VTAIL.n454 585
R1513 VTAIL.n412 VTAIL.n411 585
R1514 VTAIL.n449 VTAIL.n448 585
R1515 VTAIL.n447 VTAIL.n414 585
R1516 VTAIL.n446 VTAIL.n445 585
R1517 VTAIL.n417 VTAIL.n415 585
R1518 VTAIL.n440 VTAIL.n439 585
R1519 VTAIL.n438 VTAIL.n437 585
R1520 VTAIL.n421 VTAIL.n420 585
R1521 VTAIL.n432 VTAIL.n431 585
R1522 VTAIL.n430 VTAIL.n429 585
R1523 VTAIL.n425 VTAIL.n424 585
R1524 VTAIL.n397 VTAIL.n396 585
R1525 VTAIL.n395 VTAIL.n394 585
R1526 VTAIL.n340 VTAIL.n339 585
R1527 VTAIL.n389 VTAIL.n388 585
R1528 VTAIL.n387 VTAIL.n386 585
R1529 VTAIL.n344 VTAIL.n343 585
R1530 VTAIL.n381 VTAIL.n380 585
R1531 VTAIL.n379 VTAIL.n346 585
R1532 VTAIL.n378 VTAIL.n377 585
R1533 VTAIL.n349 VTAIL.n347 585
R1534 VTAIL.n372 VTAIL.n371 585
R1535 VTAIL.n370 VTAIL.n369 585
R1536 VTAIL.n353 VTAIL.n352 585
R1537 VTAIL.n364 VTAIL.n363 585
R1538 VTAIL.n362 VTAIL.n361 585
R1539 VTAIL.n357 VTAIL.n356 585
R1540 VTAIL.n331 VTAIL.n330 585
R1541 VTAIL.n329 VTAIL.n328 585
R1542 VTAIL.n274 VTAIL.n273 585
R1543 VTAIL.n323 VTAIL.n322 585
R1544 VTAIL.n321 VTAIL.n320 585
R1545 VTAIL.n278 VTAIL.n277 585
R1546 VTAIL.n315 VTAIL.n314 585
R1547 VTAIL.n313 VTAIL.n280 585
R1548 VTAIL.n312 VTAIL.n311 585
R1549 VTAIL.n283 VTAIL.n281 585
R1550 VTAIL.n306 VTAIL.n305 585
R1551 VTAIL.n304 VTAIL.n303 585
R1552 VTAIL.n287 VTAIL.n286 585
R1553 VTAIL.n298 VTAIL.n297 585
R1554 VTAIL.n296 VTAIL.n295 585
R1555 VTAIL.n291 VTAIL.n290 585
R1556 VTAIL.n263 VTAIL.n262 585
R1557 VTAIL.n261 VTAIL.n260 585
R1558 VTAIL.n206 VTAIL.n205 585
R1559 VTAIL.n255 VTAIL.n254 585
R1560 VTAIL.n253 VTAIL.n252 585
R1561 VTAIL.n210 VTAIL.n209 585
R1562 VTAIL.n247 VTAIL.n246 585
R1563 VTAIL.n245 VTAIL.n212 585
R1564 VTAIL.n244 VTAIL.n243 585
R1565 VTAIL.n215 VTAIL.n213 585
R1566 VTAIL.n238 VTAIL.n237 585
R1567 VTAIL.n236 VTAIL.n235 585
R1568 VTAIL.n219 VTAIL.n218 585
R1569 VTAIL.n230 VTAIL.n229 585
R1570 VTAIL.n228 VTAIL.n227 585
R1571 VTAIL.n223 VTAIL.n222 585
R1572 VTAIL.n491 VTAIL.t7 329.036
R1573 VTAIL.n23 VTAIL.t11 329.036
R1574 VTAIL.n89 VTAIL.t15 329.036
R1575 VTAIL.n157 VTAIL.t0 329.036
R1576 VTAIL.n426 VTAIL.t6 329.036
R1577 VTAIL.n358 VTAIL.t4 329.036
R1578 VTAIL.n292 VTAIL.t12 329.036
R1579 VTAIL.n224 VTAIL.t13 329.036
R1580 VTAIL.n495 VTAIL.n489 171.744
R1581 VTAIL.n496 VTAIL.n495 171.744
R1582 VTAIL.n496 VTAIL.n485 171.744
R1583 VTAIL.n503 VTAIL.n485 171.744
R1584 VTAIL.n504 VTAIL.n503 171.744
R1585 VTAIL.n504 VTAIL.n481 171.744
R1586 VTAIL.n512 VTAIL.n481 171.744
R1587 VTAIL.n513 VTAIL.n512 171.744
R1588 VTAIL.n514 VTAIL.n513 171.744
R1589 VTAIL.n514 VTAIL.n477 171.744
R1590 VTAIL.n521 VTAIL.n477 171.744
R1591 VTAIL.n522 VTAIL.n521 171.744
R1592 VTAIL.n522 VTAIL.n473 171.744
R1593 VTAIL.n529 VTAIL.n473 171.744
R1594 VTAIL.n530 VTAIL.n529 171.744
R1595 VTAIL.n27 VTAIL.n21 171.744
R1596 VTAIL.n28 VTAIL.n27 171.744
R1597 VTAIL.n28 VTAIL.n17 171.744
R1598 VTAIL.n35 VTAIL.n17 171.744
R1599 VTAIL.n36 VTAIL.n35 171.744
R1600 VTAIL.n36 VTAIL.n13 171.744
R1601 VTAIL.n44 VTAIL.n13 171.744
R1602 VTAIL.n45 VTAIL.n44 171.744
R1603 VTAIL.n46 VTAIL.n45 171.744
R1604 VTAIL.n46 VTAIL.n9 171.744
R1605 VTAIL.n53 VTAIL.n9 171.744
R1606 VTAIL.n54 VTAIL.n53 171.744
R1607 VTAIL.n54 VTAIL.n5 171.744
R1608 VTAIL.n61 VTAIL.n5 171.744
R1609 VTAIL.n62 VTAIL.n61 171.744
R1610 VTAIL.n93 VTAIL.n87 171.744
R1611 VTAIL.n94 VTAIL.n93 171.744
R1612 VTAIL.n94 VTAIL.n83 171.744
R1613 VTAIL.n101 VTAIL.n83 171.744
R1614 VTAIL.n102 VTAIL.n101 171.744
R1615 VTAIL.n102 VTAIL.n79 171.744
R1616 VTAIL.n110 VTAIL.n79 171.744
R1617 VTAIL.n111 VTAIL.n110 171.744
R1618 VTAIL.n112 VTAIL.n111 171.744
R1619 VTAIL.n112 VTAIL.n75 171.744
R1620 VTAIL.n119 VTAIL.n75 171.744
R1621 VTAIL.n120 VTAIL.n119 171.744
R1622 VTAIL.n120 VTAIL.n71 171.744
R1623 VTAIL.n127 VTAIL.n71 171.744
R1624 VTAIL.n128 VTAIL.n127 171.744
R1625 VTAIL.n161 VTAIL.n155 171.744
R1626 VTAIL.n162 VTAIL.n161 171.744
R1627 VTAIL.n162 VTAIL.n151 171.744
R1628 VTAIL.n169 VTAIL.n151 171.744
R1629 VTAIL.n170 VTAIL.n169 171.744
R1630 VTAIL.n170 VTAIL.n147 171.744
R1631 VTAIL.n178 VTAIL.n147 171.744
R1632 VTAIL.n179 VTAIL.n178 171.744
R1633 VTAIL.n180 VTAIL.n179 171.744
R1634 VTAIL.n180 VTAIL.n143 171.744
R1635 VTAIL.n187 VTAIL.n143 171.744
R1636 VTAIL.n188 VTAIL.n187 171.744
R1637 VTAIL.n188 VTAIL.n139 171.744
R1638 VTAIL.n195 VTAIL.n139 171.744
R1639 VTAIL.n196 VTAIL.n195 171.744
R1640 VTAIL.n464 VTAIL.n463 171.744
R1641 VTAIL.n463 VTAIL.n407 171.744
R1642 VTAIL.n456 VTAIL.n407 171.744
R1643 VTAIL.n456 VTAIL.n455 171.744
R1644 VTAIL.n455 VTAIL.n411 171.744
R1645 VTAIL.n448 VTAIL.n411 171.744
R1646 VTAIL.n448 VTAIL.n447 171.744
R1647 VTAIL.n447 VTAIL.n446 171.744
R1648 VTAIL.n446 VTAIL.n415 171.744
R1649 VTAIL.n439 VTAIL.n415 171.744
R1650 VTAIL.n439 VTAIL.n438 171.744
R1651 VTAIL.n438 VTAIL.n420 171.744
R1652 VTAIL.n431 VTAIL.n420 171.744
R1653 VTAIL.n431 VTAIL.n430 171.744
R1654 VTAIL.n430 VTAIL.n424 171.744
R1655 VTAIL.n396 VTAIL.n395 171.744
R1656 VTAIL.n395 VTAIL.n339 171.744
R1657 VTAIL.n388 VTAIL.n339 171.744
R1658 VTAIL.n388 VTAIL.n387 171.744
R1659 VTAIL.n387 VTAIL.n343 171.744
R1660 VTAIL.n380 VTAIL.n343 171.744
R1661 VTAIL.n380 VTAIL.n379 171.744
R1662 VTAIL.n379 VTAIL.n378 171.744
R1663 VTAIL.n378 VTAIL.n347 171.744
R1664 VTAIL.n371 VTAIL.n347 171.744
R1665 VTAIL.n371 VTAIL.n370 171.744
R1666 VTAIL.n370 VTAIL.n352 171.744
R1667 VTAIL.n363 VTAIL.n352 171.744
R1668 VTAIL.n363 VTAIL.n362 171.744
R1669 VTAIL.n362 VTAIL.n356 171.744
R1670 VTAIL.n330 VTAIL.n329 171.744
R1671 VTAIL.n329 VTAIL.n273 171.744
R1672 VTAIL.n322 VTAIL.n273 171.744
R1673 VTAIL.n322 VTAIL.n321 171.744
R1674 VTAIL.n321 VTAIL.n277 171.744
R1675 VTAIL.n314 VTAIL.n277 171.744
R1676 VTAIL.n314 VTAIL.n313 171.744
R1677 VTAIL.n313 VTAIL.n312 171.744
R1678 VTAIL.n312 VTAIL.n281 171.744
R1679 VTAIL.n305 VTAIL.n281 171.744
R1680 VTAIL.n305 VTAIL.n304 171.744
R1681 VTAIL.n304 VTAIL.n286 171.744
R1682 VTAIL.n297 VTAIL.n286 171.744
R1683 VTAIL.n297 VTAIL.n296 171.744
R1684 VTAIL.n296 VTAIL.n290 171.744
R1685 VTAIL.n262 VTAIL.n261 171.744
R1686 VTAIL.n261 VTAIL.n205 171.744
R1687 VTAIL.n254 VTAIL.n205 171.744
R1688 VTAIL.n254 VTAIL.n253 171.744
R1689 VTAIL.n253 VTAIL.n209 171.744
R1690 VTAIL.n246 VTAIL.n209 171.744
R1691 VTAIL.n246 VTAIL.n245 171.744
R1692 VTAIL.n245 VTAIL.n244 171.744
R1693 VTAIL.n244 VTAIL.n213 171.744
R1694 VTAIL.n237 VTAIL.n213 171.744
R1695 VTAIL.n237 VTAIL.n236 171.744
R1696 VTAIL.n236 VTAIL.n218 171.744
R1697 VTAIL.n229 VTAIL.n218 171.744
R1698 VTAIL.n229 VTAIL.n228 171.744
R1699 VTAIL.n228 VTAIL.n222 171.744
R1700 VTAIL.t7 VTAIL.n489 85.8723
R1701 VTAIL.t11 VTAIL.n21 85.8723
R1702 VTAIL.t15 VTAIL.n87 85.8723
R1703 VTAIL.t0 VTAIL.n155 85.8723
R1704 VTAIL.t6 VTAIL.n424 85.8723
R1705 VTAIL.t4 VTAIL.n356 85.8723
R1706 VTAIL.t12 VTAIL.n290 85.8723
R1707 VTAIL.t13 VTAIL.n222 85.8723
R1708 VTAIL.n403 VTAIL.n402 57.5483
R1709 VTAIL.n269 VTAIL.n268 57.5483
R1710 VTAIL.n1 VTAIL.n0 57.5481
R1711 VTAIL.n135 VTAIL.n134 57.5481
R1712 VTAIL.n535 VTAIL.n534 32.5732
R1713 VTAIL.n67 VTAIL.n66 32.5732
R1714 VTAIL.n133 VTAIL.n132 32.5732
R1715 VTAIL.n201 VTAIL.n200 32.5732
R1716 VTAIL.n469 VTAIL.n468 32.5732
R1717 VTAIL.n401 VTAIL.n400 32.5732
R1718 VTAIL.n335 VTAIL.n334 32.5732
R1719 VTAIL.n267 VTAIL.n266 32.5732
R1720 VTAIL.n535 VTAIL.n469 25.8927
R1721 VTAIL.n267 VTAIL.n201 25.8927
R1722 VTAIL.n515 VTAIL.n480 13.1884
R1723 VTAIL.n47 VTAIL.n12 13.1884
R1724 VTAIL.n113 VTAIL.n78 13.1884
R1725 VTAIL.n181 VTAIL.n146 13.1884
R1726 VTAIL.n449 VTAIL.n414 13.1884
R1727 VTAIL.n381 VTAIL.n346 13.1884
R1728 VTAIL.n315 VTAIL.n280 13.1884
R1729 VTAIL.n247 VTAIL.n212 13.1884
R1730 VTAIL.n511 VTAIL.n510 12.8005
R1731 VTAIL.n516 VTAIL.n478 12.8005
R1732 VTAIL.n43 VTAIL.n42 12.8005
R1733 VTAIL.n48 VTAIL.n10 12.8005
R1734 VTAIL.n109 VTAIL.n108 12.8005
R1735 VTAIL.n114 VTAIL.n76 12.8005
R1736 VTAIL.n177 VTAIL.n176 12.8005
R1737 VTAIL.n182 VTAIL.n144 12.8005
R1738 VTAIL.n450 VTAIL.n412 12.8005
R1739 VTAIL.n445 VTAIL.n416 12.8005
R1740 VTAIL.n382 VTAIL.n344 12.8005
R1741 VTAIL.n377 VTAIL.n348 12.8005
R1742 VTAIL.n316 VTAIL.n278 12.8005
R1743 VTAIL.n311 VTAIL.n282 12.8005
R1744 VTAIL.n248 VTAIL.n210 12.8005
R1745 VTAIL.n243 VTAIL.n214 12.8005
R1746 VTAIL.n509 VTAIL.n482 12.0247
R1747 VTAIL.n520 VTAIL.n519 12.0247
R1748 VTAIL.n41 VTAIL.n14 12.0247
R1749 VTAIL.n52 VTAIL.n51 12.0247
R1750 VTAIL.n107 VTAIL.n80 12.0247
R1751 VTAIL.n118 VTAIL.n117 12.0247
R1752 VTAIL.n175 VTAIL.n148 12.0247
R1753 VTAIL.n186 VTAIL.n185 12.0247
R1754 VTAIL.n454 VTAIL.n453 12.0247
R1755 VTAIL.n444 VTAIL.n417 12.0247
R1756 VTAIL.n386 VTAIL.n385 12.0247
R1757 VTAIL.n376 VTAIL.n349 12.0247
R1758 VTAIL.n320 VTAIL.n319 12.0247
R1759 VTAIL.n310 VTAIL.n283 12.0247
R1760 VTAIL.n252 VTAIL.n251 12.0247
R1761 VTAIL.n242 VTAIL.n215 12.0247
R1762 VTAIL.n506 VTAIL.n505 11.249
R1763 VTAIL.n523 VTAIL.n476 11.249
R1764 VTAIL.n38 VTAIL.n37 11.249
R1765 VTAIL.n55 VTAIL.n8 11.249
R1766 VTAIL.n104 VTAIL.n103 11.249
R1767 VTAIL.n121 VTAIL.n74 11.249
R1768 VTAIL.n172 VTAIL.n171 11.249
R1769 VTAIL.n189 VTAIL.n142 11.249
R1770 VTAIL.n457 VTAIL.n410 11.249
R1771 VTAIL.n441 VTAIL.n440 11.249
R1772 VTAIL.n389 VTAIL.n342 11.249
R1773 VTAIL.n373 VTAIL.n372 11.249
R1774 VTAIL.n323 VTAIL.n276 11.249
R1775 VTAIL.n307 VTAIL.n306 11.249
R1776 VTAIL.n255 VTAIL.n208 11.249
R1777 VTAIL.n239 VTAIL.n238 11.249
R1778 VTAIL.n491 VTAIL.n490 10.7239
R1779 VTAIL.n23 VTAIL.n22 10.7239
R1780 VTAIL.n89 VTAIL.n88 10.7239
R1781 VTAIL.n157 VTAIL.n156 10.7239
R1782 VTAIL.n426 VTAIL.n425 10.7239
R1783 VTAIL.n358 VTAIL.n357 10.7239
R1784 VTAIL.n292 VTAIL.n291 10.7239
R1785 VTAIL.n224 VTAIL.n223 10.7239
R1786 VTAIL.n502 VTAIL.n484 10.4732
R1787 VTAIL.n524 VTAIL.n474 10.4732
R1788 VTAIL.n34 VTAIL.n16 10.4732
R1789 VTAIL.n56 VTAIL.n6 10.4732
R1790 VTAIL.n100 VTAIL.n82 10.4732
R1791 VTAIL.n122 VTAIL.n72 10.4732
R1792 VTAIL.n168 VTAIL.n150 10.4732
R1793 VTAIL.n190 VTAIL.n140 10.4732
R1794 VTAIL.n458 VTAIL.n408 10.4732
R1795 VTAIL.n437 VTAIL.n419 10.4732
R1796 VTAIL.n390 VTAIL.n340 10.4732
R1797 VTAIL.n369 VTAIL.n351 10.4732
R1798 VTAIL.n324 VTAIL.n274 10.4732
R1799 VTAIL.n303 VTAIL.n285 10.4732
R1800 VTAIL.n256 VTAIL.n206 10.4732
R1801 VTAIL.n235 VTAIL.n217 10.4732
R1802 VTAIL.n501 VTAIL.n486 9.69747
R1803 VTAIL.n528 VTAIL.n527 9.69747
R1804 VTAIL.n33 VTAIL.n18 9.69747
R1805 VTAIL.n60 VTAIL.n59 9.69747
R1806 VTAIL.n99 VTAIL.n84 9.69747
R1807 VTAIL.n126 VTAIL.n125 9.69747
R1808 VTAIL.n167 VTAIL.n152 9.69747
R1809 VTAIL.n194 VTAIL.n193 9.69747
R1810 VTAIL.n462 VTAIL.n461 9.69747
R1811 VTAIL.n436 VTAIL.n421 9.69747
R1812 VTAIL.n394 VTAIL.n393 9.69747
R1813 VTAIL.n368 VTAIL.n353 9.69747
R1814 VTAIL.n328 VTAIL.n327 9.69747
R1815 VTAIL.n302 VTAIL.n287 9.69747
R1816 VTAIL.n260 VTAIL.n259 9.69747
R1817 VTAIL.n234 VTAIL.n219 9.69747
R1818 VTAIL.n534 VTAIL.n533 9.45567
R1819 VTAIL.n66 VTAIL.n65 9.45567
R1820 VTAIL.n132 VTAIL.n131 9.45567
R1821 VTAIL.n200 VTAIL.n199 9.45567
R1822 VTAIL.n468 VTAIL.n467 9.45567
R1823 VTAIL.n400 VTAIL.n399 9.45567
R1824 VTAIL.n334 VTAIL.n333 9.45567
R1825 VTAIL.n266 VTAIL.n265 9.45567
R1826 VTAIL.n533 VTAIL.n532 9.3005
R1827 VTAIL.n472 VTAIL.n471 9.3005
R1828 VTAIL.n527 VTAIL.n526 9.3005
R1829 VTAIL.n525 VTAIL.n524 9.3005
R1830 VTAIL.n476 VTAIL.n475 9.3005
R1831 VTAIL.n519 VTAIL.n518 9.3005
R1832 VTAIL.n517 VTAIL.n516 9.3005
R1833 VTAIL.n493 VTAIL.n492 9.3005
R1834 VTAIL.n488 VTAIL.n487 9.3005
R1835 VTAIL.n499 VTAIL.n498 9.3005
R1836 VTAIL.n501 VTAIL.n500 9.3005
R1837 VTAIL.n484 VTAIL.n483 9.3005
R1838 VTAIL.n507 VTAIL.n506 9.3005
R1839 VTAIL.n509 VTAIL.n508 9.3005
R1840 VTAIL.n510 VTAIL.n479 9.3005
R1841 VTAIL.n65 VTAIL.n64 9.3005
R1842 VTAIL.n4 VTAIL.n3 9.3005
R1843 VTAIL.n59 VTAIL.n58 9.3005
R1844 VTAIL.n57 VTAIL.n56 9.3005
R1845 VTAIL.n8 VTAIL.n7 9.3005
R1846 VTAIL.n51 VTAIL.n50 9.3005
R1847 VTAIL.n49 VTAIL.n48 9.3005
R1848 VTAIL.n25 VTAIL.n24 9.3005
R1849 VTAIL.n20 VTAIL.n19 9.3005
R1850 VTAIL.n31 VTAIL.n30 9.3005
R1851 VTAIL.n33 VTAIL.n32 9.3005
R1852 VTAIL.n16 VTAIL.n15 9.3005
R1853 VTAIL.n39 VTAIL.n38 9.3005
R1854 VTAIL.n41 VTAIL.n40 9.3005
R1855 VTAIL.n42 VTAIL.n11 9.3005
R1856 VTAIL.n131 VTAIL.n130 9.3005
R1857 VTAIL.n70 VTAIL.n69 9.3005
R1858 VTAIL.n125 VTAIL.n124 9.3005
R1859 VTAIL.n123 VTAIL.n122 9.3005
R1860 VTAIL.n74 VTAIL.n73 9.3005
R1861 VTAIL.n117 VTAIL.n116 9.3005
R1862 VTAIL.n115 VTAIL.n114 9.3005
R1863 VTAIL.n91 VTAIL.n90 9.3005
R1864 VTAIL.n86 VTAIL.n85 9.3005
R1865 VTAIL.n97 VTAIL.n96 9.3005
R1866 VTAIL.n99 VTAIL.n98 9.3005
R1867 VTAIL.n82 VTAIL.n81 9.3005
R1868 VTAIL.n105 VTAIL.n104 9.3005
R1869 VTAIL.n107 VTAIL.n106 9.3005
R1870 VTAIL.n108 VTAIL.n77 9.3005
R1871 VTAIL.n199 VTAIL.n198 9.3005
R1872 VTAIL.n138 VTAIL.n137 9.3005
R1873 VTAIL.n193 VTAIL.n192 9.3005
R1874 VTAIL.n191 VTAIL.n190 9.3005
R1875 VTAIL.n142 VTAIL.n141 9.3005
R1876 VTAIL.n185 VTAIL.n184 9.3005
R1877 VTAIL.n183 VTAIL.n182 9.3005
R1878 VTAIL.n159 VTAIL.n158 9.3005
R1879 VTAIL.n154 VTAIL.n153 9.3005
R1880 VTAIL.n165 VTAIL.n164 9.3005
R1881 VTAIL.n167 VTAIL.n166 9.3005
R1882 VTAIL.n150 VTAIL.n149 9.3005
R1883 VTAIL.n173 VTAIL.n172 9.3005
R1884 VTAIL.n175 VTAIL.n174 9.3005
R1885 VTAIL.n176 VTAIL.n145 9.3005
R1886 VTAIL.n428 VTAIL.n427 9.3005
R1887 VTAIL.n423 VTAIL.n422 9.3005
R1888 VTAIL.n434 VTAIL.n433 9.3005
R1889 VTAIL.n436 VTAIL.n435 9.3005
R1890 VTAIL.n419 VTAIL.n418 9.3005
R1891 VTAIL.n442 VTAIL.n441 9.3005
R1892 VTAIL.n444 VTAIL.n443 9.3005
R1893 VTAIL.n416 VTAIL.n413 9.3005
R1894 VTAIL.n467 VTAIL.n466 9.3005
R1895 VTAIL.n406 VTAIL.n405 9.3005
R1896 VTAIL.n461 VTAIL.n460 9.3005
R1897 VTAIL.n459 VTAIL.n458 9.3005
R1898 VTAIL.n410 VTAIL.n409 9.3005
R1899 VTAIL.n453 VTAIL.n452 9.3005
R1900 VTAIL.n451 VTAIL.n450 9.3005
R1901 VTAIL.n360 VTAIL.n359 9.3005
R1902 VTAIL.n355 VTAIL.n354 9.3005
R1903 VTAIL.n366 VTAIL.n365 9.3005
R1904 VTAIL.n368 VTAIL.n367 9.3005
R1905 VTAIL.n351 VTAIL.n350 9.3005
R1906 VTAIL.n374 VTAIL.n373 9.3005
R1907 VTAIL.n376 VTAIL.n375 9.3005
R1908 VTAIL.n348 VTAIL.n345 9.3005
R1909 VTAIL.n399 VTAIL.n398 9.3005
R1910 VTAIL.n338 VTAIL.n337 9.3005
R1911 VTAIL.n393 VTAIL.n392 9.3005
R1912 VTAIL.n391 VTAIL.n390 9.3005
R1913 VTAIL.n342 VTAIL.n341 9.3005
R1914 VTAIL.n385 VTAIL.n384 9.3005
R1915 VTAIL.n383 VTAIL.n382 9.3005
R1916 VTAIL.n294 VTAIL.n293 9.3005
R1917 VTAIL.n289 VTAIL.n288 9.3005
R1918 VTAIL.n300 VTAIL.n299 9.3005
R1919 VTAIL.n302 VTAIL.n301 9.3005
R1920 VTAIL.n285 VTAIL.n284 9.3005
R1921 VTAIL.n308 VTAIL.n307 9.3005
R1922 VTAIL.n310 VTAIL.n309 9.3005
R1923 VTAIL.n282 VTAIL.n279 9.3005
R1924 VTAIL.n333 VTAIL.n332 9.3005
R1925 VTAIL.n272 VTAIL.n271 9.3005
R1926 VTAIL.n327 VTAIL.n326 9.3005
R1927 VTAIL.n325 VTAIL.n324 9.3005
R1928 VTAIL.n276 VTAIL.n275 9.3005
R1929 VTAIL.n319 VTAIL.n318 9.3005
R1930 VTAIL.n317 VTAIL.n316 9.3005
R1931 VTAIL.n226 VTAIL.n225 9.3005
R1932 VTAIL.n221 VTAIL.n220 9.3005
R1933 VTAIL.n232 VTAIL.n231 9.3005
R1934 VTAIL.n234 VTAIL.n233 9.3005
R1935 VTAIL.n217 VTAIL.n216 9.3005
R1936 VTAIL.n240 VTAIL.n239 9.3005
R1937 VTAIL.n242 VTAIL.n241 9.3005
R1938 VTAIL.n214 VTAIL.n211 9.3005
R1939 VTAIL.n265 VTAIL.n264 9.3005
R1940 VTAIL.n204 VTAIL.n203 9.3005
R1941 VTAIL.n259 VTAIL.n258 9.3005
R1942 VTAIL.n257 VTAIL.n256 9.3005
R1943 VTAIL.n208 VTAIL.n207 9.3005
R1944 VTAIL.n251 VTAIL.n250 9.3005
R1945 VTAIL.n249 VTAIL.n248 9.3005
R1946 VTAIL.n498 VTAIL.n497 8.92171
R1947 VTAIL.n531 VTAIL.n472 8.92171
R1948 VTAIL.n30 VTAIL.n29 8.92171
R1949 VTAIL.n63 VTAIL.n4 8.92171
R1950 VTAIL.n96 VTAIL.n95 8.92171
R1951 VTAIL.n129 VTAIL.n70 8.92171
R1952 VTAIL.n164 VTAIL.n163 8.92171
R1953 VTAIL.n197 VTAIL.n138 8.92171
R1954 VTAIL.n465 VTAIL.n406 8.92171
R1955 VTAIL.n433 VTAIL.n432 8.92171
R1956 VTAIL.n397 VTAIL.n338 8.92171
R1957 VTAIL.n365 VTAIL.n364 8.92171
R1958 VTAIL.n331 VTAIL.n272 8.92171
R1959 VTAIL.n299 VTAIL.n298 8.92171
R1960 VTAIL.n263 VTAIL.n204 8.92171
R1961 VTAIL.n231 VTAIL.n230 8.92171
R1962 VTAIL.n494 VTAIL.n488 8.14595
R1963 VTAIL.n532 VTAIL.n470 8.14595
R1964 VTAIL.n26 VTAIL.n20 8.14595
R1965 VTAIL.n64 VTAIL.n2 8.14595
R1966 VTAIL.n92 VTAIL.n86 8.14595
R1967 VTAIL.n130 VTAIL.n68 8.14595
R1968 VTAIL.n160 VTAIL.n154 8.14595
R1969 VTAIL.n198 VTAIL.n136 8.14595
R1970 VTAIL.n466 VTAIL.n404 8.14595
R1971 VTAIL.n429 VTAIL.n423 8.14595
R1972 VTAIL.n398 VTAIL.n336 8.14595
R1973 VTAIL.n361 VTAIL.n355 8.14595
R1974 VTAIL.n332 VTAIL.n270 8.14595
R1975 VTAIL.n295 VTAIL.n289 8.14595
R1976 VTAIL.n264 VTAIL.n202 8.14595
R1977 VTAIL.n227 VTAIL.n221 8.14595
R1978 VTAIL.n493 VTAIL.n490 7.3702
R1979 VTAIL.n25 VTAIL.n22 7.3702
R1980 VTAIL.n91 VTAIL.n88 7.3702
R1981 VTAIL.n159 VTAIL.n156 7.3702
R1982 VTAIL.n428 VTAIL.n425 7.3702
R1983 VTAIL.n360 VTAIL.n357 7.3702
R1984 VTAIL.n294 VTAIL.n291 7.3702
R1985 VTAIL.n226 VTAIL.n223 7.3702
R1986 VTAIL.n494 VTAIL.n493 5.81868
R1987 VTAIL.n534 VTAIL.n470 5.81868
R1988 VTAIL.n26 VTAIL.n25 5.81868
R1989 VTAIL.n66 VTAIL.n2 5.81868
R1990 VTAIL.n92 VTAIL.n91 5.81868
R1991 VTAIL.n132 VTAIL.n68 5.81868
R1992 VTAIL.n160 VTAIL.n159 5.81868
R1993 VTAIL.n200 VTAIL.n136 5.81868
R1994 VTAIL.n468 VTAIL.n404 5.81868
R1995 VTAIL.n429 VTAIL.n428 5.81868
R1996 VTAIL.n400 VTAIL.n336 5.81868
R1997 VTAIL.n361 VTAIL.n360 5.81868
R1998 VTAIL.n334 VTAIL.n270 5.81868
R1999 VTAIL.n295 VTAIL.n294 5.81868
R2000 VTAIL.n266 VTAIL.n202 5.81868
R2001 VTAIL.n227 VTAIL.n226 5.81868
R2002 VTAIL.n497 VTAIL.n488 5.04292
R2003 VTAIL.n532 VTAIL.n531 5.04292
R2004 VTAIL.n29 VTAIL.n20 5.04292
R2005 VTAIL.n64 VTAIL.n63 5.04292
R2006 VTAIL.n95 VTAIL.n86 5.04292
R2007 VTAIL.n130 VTAIL.n129 5.04292
R2008 VTAIL.n163 VTAIL.n154 5.04292
R2009 VTAIL.n198 VTAIL.n197 5.04292
R2010 VTAIL.n466 VTAIL.n465 5.04292
R2011 VTAIL.n432 VTAIL.n423 5.04292
R2012 VTAIL.n398 VTAIL.n397 5.04292
R2013 VTAIL.n364 VTAIL.n355 5.04292
R2014 VTAIL.n332 VTAIL.n331 5.04292
R2015 VTAIL.n298 VTAIL.n289 5.04292
R2016 VTAIL.n264 VTAIL.n263 5.04292
R2017 VTAIL.n230 VTAIL.n221 5.04292
R2018 VTAIL.n498 VTAIL.n486 4.26717
R2019 VTAIL.n528 VTAIL.n472 4.26717
R2020 VTAIL.n30 VTAIL.n18 4.26717
R2021 VTAIL.n60 VTAIL.n4 4.26717
R2022 VTAIL.n96 VTAIL.n84 4.26717
R2023 VTAIL.n126 VTAIL.n70 4.26717
R2024 VTAIL.n164 VTAIL.n152 4.26717
R2025 VTAIL.n194 VTAIL.n138 4.26717
R2026 VTAIL.n462 VTAIL.n406 4.26717
R2027 VTAIL.n433 VTAIL.n421 4.26717
R2028 VTAIL.n394 VTAIL.n338 4.26717
R2029 VTAIL.n365 VTAIL.n353 4.26717
R2030 VTAIL.n328 VTAIL.n272 4.26717
R2031 VTAIL.n299 VTAIL.n287 4.26717
R2032 VTAIL.n260 VTAIL.n204 4.26717
R2033 VTAIL.n231 VTAIL.n219 4.26717
R2034 VTAIL.n502 VTAIL.n501 3.49141
R2035 VTAIL.n527 VTAIL.n474 3.49141
R2036 VTAIL.n34 VTAIL.n33 3.49141
R2037 VTAIL.n59 VTAIL.n6 3.49141
R2038 VTAIL.n100 VTAIL.n99 3.49141
R2039 VTAIL.n125 VTAIL.n72 3.49141
R2040 VTAIL.n168 VTAIL.n167 3.49141
R2041 VTAIL.n193 VTAIL.n140 3.49141
R2042 VTAIL.n461 VTAIL.n408 3.49141
R2043 VTAIL.n437 VTAIL.n436 3.49141
R2044 VTAIL.n393 VTAIL.n340 3.49141
R2045 VTAIL.n369 VTAIL.n368 3.49141
R2046 VTAIL.n327 VTAIL.n274 3.49141
R2047 VTAIL.n303 VTAIL.n302 3.49141
R2048 VTAIL.n259 VTAIL.n206 3.49141
R2049 VTAIL.n235 VTAIL.n234 3.49141
R2050 VTAIL.n269 VTAIL.n267 3.06084
R2051 VTAIL.n335 VTAIL.n269 3.06084
R2052 VTAIL.n403 VTAIL.n401 3.06084
R2053 VTAIL.n469 VTAIL.n403 3.06084
R2054 VTAIL.n201 VTAIL.n135 3.06084
R2055 VTAIL.n135 VTAIL.n133 3.06084
R2056 VTAIL.n67 VTAIL.n1 3.06084
R2057 VTAIL VTAIL.n535 3.00266
R2058 VTAIL.n505 VTAIL.n484 2.71565
R2059 VTAIL.n524 VTAIL.n523 2.71565
R2060 VTAIL.n37 VTAIL.n16 2.71565
R2061 VTAIL.n56 VTAIL.n55 2.71565
R2062 VTAIL.n103 VTAIL.n82 2.71565
R2063 VTAIL.n122 VTAIL.n121 2.71565
R2064 VTAIL.n171 VTAIL.n150 2.71565
R2065 VTAIL.n190 VTAIL.n189 2.71565
R2066 VTAIL.n458 VTAIL.n457 2.71565
R2067 VTAIL.n440 VTAIL.n419 2.71565
R2068 VTAIL.n390 VTAIL.n389 2.71565
R2069 VTAIL.n372 VTAIL.n351 2.71565
R2070 VTAIL.n324 VTAIL.n323 2.71565
R2071 VTAIL.n306 VTAIL.n285 2.71565
R2072 VTAIL.n256 VTAIL.n255 2.71565
R2073 VTAIL.n238 VTAIL.n217 2.71565
R2074 VTAIL.n0 VTAIL.t10 2.67801
R2075 VTAIL.n0 VTAIL.t8 2.67801
R2076 VTAIL.n134 VTAIL.t2 2.67801
R2077 VTAIL.n134 VTAIL.t1 2.67801
R2078 VTAIL.n402 VTAIL.t3 2.67801
R2079 VTAIL.n402 VTAIL.t5 2.67801
R2080 VTAIL.n268 VTAIL.t9 2.67801
R2081 VTAIL.n268 VTAIL.t14 2.67801
R2082 VTAIL.n427 VTAIL.n426 2.41282
R2083 VTAIL.n359 VTAIL.n358 2.41282
R2084 VTAIL.n293 VTAIL.n292 2.41282
R2085 VTAIL.n225 VTAIL.n224 2.41282
R2086 VTAIL.n492 VTAIL.n491 2.41282
R2087 VTAIL.n24 VTAIL.n23 2.41282
R2088 VTAIL.n90 VTAIL.n89 2.41282
R2089 VTAIL.n158 VTAIL.n157 2.41282
R2090 VTAIL.n506 VTAIL.n482 1.93989
R2091 VTAIL.n520 VTAIL.n476 1.93989
R2092 VTAIL.n38 VTAIL.n14 1.93989
R2093 VTAIL.n52 VTAIL.n8 1.93989
R2094 VTAIL.n104 VTAIL.n80 1.93989
R2095 VTAIL.n118 VTAIL.n74 1.93989
R2096 VTAIL.n172 VTAIL.n148 1.93989
R2097 VTAIL.n186 VTAIL.n142 1.93989
R2098 VTAIL.n454 VTAIL.n410 1.93989
R2099 VTAIL.n441 VTAIL.n417 1.93989
R2100 VTAIL.n386 VTAIL.n342 1.93989
R2101 VTAIL.n373 VTAIL.n349 1.93989
R2102 VTAIL.n320 VTAIL.n276 1.93989
R2103 VTAIL.n307 VTAIL.n283 1.93989
R2104 VTAIL.n252 VTAIL.n208 1.93989
R2105 VTAIL.n239 VTAIL.n215 1.93989
R2106 VTAIL.n511 VTAIL.n509 1.16414
R2107 VTAIL.n519 VTAIL.n478 1.16414
R2108 VTAIL.n43 VTAIL.n41 1.16414
R2109 VTAIL.n51 VTAIL.n10 1.16414
R2110 VTAIL.n109 VTAIL.n107 1.16414
R2111 VTAIL.n117 VTAIL.n76 1.16414
R2112 VTAIL.n177 VTAIL.n175 1.16414
R2113 VTAIL.n185 VTAIL.n144 1.16414
R2114 VTAIL.n453 VTAIL.n412 1.16414
R2115 VTAIL.n445 VTAIL.n444 1.16414
R2116 VTAIL.n385 VTAIL.n344 1.16414
R2117 VTAIL.n377 VTAIL.n376 1.16414
R2118 VTAIL.n319 VTAIL.n278 1.16414
R2119 VTAIL.n311 VTAIL.n310 1.16414
R2120 VTAIL.n251 VTAIL.n210 1.16414
R2121 VTAIL.n243 VTAIL.n242 1.16414
R2122 VTAIL.n401 VTAIL.n335 0.470328
R2123 VTAIL.n133 VTAIL.n67 0.470328
R2124 VTAIL.n510 VTAIL.n480 0.388379
R2125 VTAIL.n516 VTAIL.n515 0.388379
R2126 VTAIL.n42 VTAIL.n12 0.388379
R2127 VTAIL.n48 VTAIL.n47 0.388379
R2128 VTAIL.n108 VTAIL.n78 0.388379
R2129 VTAIL.n114 VTAIL.n113 0.388379
R2130 VTAIL.n176 VTAIL.n146 0.388379
R2131 VTAIL.n182 VTAIL.n181 0.388379
R2132 VTAIL.n450 VTAIL.n449 0.388379
R2133 VTAIL.n416 VTAIL.n414 0.388379
R2134 VTAIL.n382 VTAIL.n381 0.388379
R2135 VTAIL.n348 VTAIL.n346 0.388379
R2136 VTAIL.n316 VTAIL.n315 0.388379
R2137 VTAIL.n282 VTAIL.n280 0.388379
R2138 VTAIL.n248 VTAIL.n247 0.388379
R2139 VTAIL.n214 VTAIL.n212 0.388379
R2140 VTAIL.n492 VTAIL.n487 0.155672
R2141 VTAIL.n499 VTAIL.n487 0.155672
R2142 VTAIL.n500 VTAIL.n499 0.155672
R2143 VTAIL.n500 VTAIL.n483 0.155672
R2144 VTAIL.n507 VTAIL.n483 0.155672
R2145 VTAIL.n508 VTAIL.n507 0.155672
R2146 VTAIL.n508 VTAIL.n479 0.155672
R2147 VTAIL.n517 VTAIL.n479 0.155672
R2148 VTAIL.n518 VTAIL.n517 0.155672
R2149 VTAIL.n518 VTAIL.n475 0.155672
R2150 VTAIL.n525 VTAIL.n475 0.155672
R2151 VTAIL.n526 VTAIL.n525 0.155672
R2152 VTAIL.n526 VTAIL.n471 0.155672
R2153 VTAIL.n533 VTAIL.n471 0.155672
R2154 VTAIL.n24 VTAIL.n19 0.155672
R2155 VTAIL.n31 VTAIL.n19 0.155672
R2156 VTAIL.n32 VTAIL.n31 0.155672
R2157 VTAIL.n32 VTAIL.n15 0.155672
R2158 VTAIL.n39 VTAIL.n15 0.155672
R2159 VTAIL.n40 VTAIL.n39 0.155672
R2160 VTAIL.n40 VTAIL.n11 0.155672
R2161 VTAIL.n49 VTAIL.n11 0.155672
R2162 VTAIL.n50 VTAIL.n49 0.155672
R2163 VTAIL.n50 VTAIL.n7 0.155672
R2164 VTAIL.n57 VTAIL.n7 0.155672
R2165 VTAIL.n58 VTAIL.n57 0.155672
R2166 VTAIL.n58 VTAIL.n3 0.155672
R2167 VTAIL.n65 VTAIL.n3 0.155672
R2168 VTAIL.n90 VTAIL.n85 0.155672
R2169 VTAIL.n97 VTAIL.n85 0.155672
R2170 VTAIL.n98 VTAIL.n97 0.155672
R2171 VTAIL.n98 VTAIL.n81 0.155672
R2172 VTAIL.n105 VTAIL.n81 0.155672
R2173 VTAIL.n106 VTAIL.n105 0.155672
R2174 VTAIL.n106 VTAIL.n77 0.155672
R2175 VTAIL.n115 VTAIL.n77 0.155672
R2176 VTAIL.n116 VTAIL.n115 0.155672
R2177 VTAIL.n116 VTAIL.n73 0.155672
R2178 VTAIL.n123 VTAIL.n73 0.155672
R2179 VTAIL.n124 VTAIL.n123 0.155672
R2180 VTAIL.n124 VTAIL.n69 0.155672
R2181 VTAIL.n131 VTAIL.n69 0.155672
R2182 VTAIL.n158 VTAIL.n153 0.155672
R2183 VTAIL.n165 VTAIL.n153 0.155672
R2184 VTAIL.n166 VTAIL.n165 0.155672
R2185 VTAIL.n166 VTAIL.n149 0.155672
R2186 VTAIL.n173 VTAIL.n149 0.155672
R2187 VTAIL.n174 VTAIL.n173 0.155672
R2188 VTAIL.n174 VTAIL.n145 0.155672
R2189 VTAIL.n183 VTAIL.n145 0.155672
R2190 VTAIL.n184 VTAIL.n183 0.155672
R2191 VTAIL.n184 VTAIL.n141 0.155672
R2192 VTAIL.n191 VTAIL.n141 0.155672
R2193 VTAIL.n192 VTAIL.n191 0.155672
R2194 VTAIL.n192 VTAIL.n137 0.155672
R2195 VTAIL.n199 VTAIL.n137 0.155672
R2196 VTAIL.n467 VTAIL.n405 0.155672
R2197 VTAIL.n460 VTAIL.n405 0.155672
R2198 VTAIL.n460 VTAIL.n459 0.155672
R2199 VTAIL.n459 VTAIL.n409 0.155672
R2200 VTAIL.n452 VTAIL.n409 0.155672
R2201 VTAIL.n452 VTAIL.n451 0.155672
R2202 VTAIL.n451 VTAIL.n413 0.155672
R2203 VTAIL.n443 VTAIL.n413 0.155672
R2204 VTAIL.n443 VTAIL.n442 0.155672
R2205 VTAIL.n442 VTAIL.n418 0.155672
R2206 VTAIL.n435 VTAIL.n418 0.155672
R2207 VTAIL.n435 VTAIL.n434 0.155672
R2208 VTAIL.n434 VTAIL.n422 0.155672
R2209 VTAIL.n427 VTAIL.n422 0.155672
R2210 VTAIL.n399 VTAIL.n337 0.155672
R2211 VTAIL.n392 VTAIL.n337 0.155672
R2212 VTAIL.n392 VTAIL.n391 0.155672
R2213 VTAIL.n391 VTAIL.n341 0.155672
R2214 VTAIL.n384 VTAIL.n341 0.155672
R2215 VTAIL.n384 VTAIL.n383 0.155672
R2216 VTAIL.n383 VTAIL.n345 0.155672
R2217 VTAIL.n375 VTAIL.n345 0.155672
R2218 VTAIL.n375 VTAIL.n374 0.155672
R2219 VTAIL.n374 VTAIL.n350 0.155672
R2220 VTAIL.n367 VTAIL.n350 0.155672
R2221 VTAIL.n367 VTAIL.n366 0.155672
R2222 VTAIL.n366 VTAIL.n354 0.155672
R2223 VTAIL.n359 VTAIL.n354 0.155672
R2224 VTAIL.n333 VTAIL.n271 0.155672
R2225 VTAIL.n326 VTAIL.n271 0.155672
R2226 VTAIL.n326 VTAIL.n325 0.155672
R2227 VTAIL.n325 VTAIL.n275 0.155672
R2228 VTAIL.n318 VTAIL.n275 0.155672
R2229 VTAIL.n318 VTAIL.n317 0.155672
R2230 VTAIL.n317 VTAIL.n279 0.155672
R2231 VTAIL.n309 VTAIL.n279 0.155672
R2232 VTAIL.n309 VTAIL.n308 0.155672
R2233 VTAIL.n308 VTAIL.n284 0.155672
R2234 VTAIL.n301 VTAIL.n284 0.155672
R2235 VTAIL.n301 VTAIL.n300 0.155672
R2236 VTAIL.n300 VTAIL.n288 0.155672
R2237 VTAIL.n293 VTAIL.n288 0.155672
R2238 VTAIL.n265 VTAIL.n203 0.155672
R2239 VTAIL.n258 VTAIL.n203 0.155672
R2240 VTAIL.n258 VTAIL.n257 0.155672
R2241 VTAIL.n257 VTAIL.n207 0.155672
R2242 VTAIL.n250 VTAIL.n207 0.155672
R2243 VTAIL.n250 VTAIL.n249 0.155672
R2244 VTAIL.n249 VTAIL.n211 0.155672
R2245 VTAIL.n241 VTAIL.n211 0.155672
R2246 VTAIL.n241 VTAIL.n240 0.155672
R2247 VTAIL.n240 VTAIL.n216 0.155672
R2248 VTAIL.n233 VTAIL.n216 0.155672
R2249 VTAIL.n233 VTAIL.n232 0.155672
R2250 VTAIL.n232 VTAIL.n220 0.155672
R2251 VTAIL.n225 VTAIL.n220 0.155672
R2252 VTAIL VTAIL.n1 0.0586897
R2253 VP.n24 VP.n23 161.3
R2254 VP.n25 VP.n20 161.3
R2255 VP.n27 VP.n26 161.3
R2256 VP.n28 VP.n19 161.3
R2257 VP.n30 VP.n29 161.3
R2258 VP.n31 VP.n18 161.3
R2259 VP.n33 VP.n32 161.3
R2260 VP.n35 VP.n34 161.3
R2261 VP.n36 VP.n16 161.3
R2262 VP.n38 VP.n37 161.3
R2263 VP.n39 VP.n15 161.3
R2264 VP.n41 VP.n40 161.3
R2265 VP.n42 VP.n14 161.3
R2266 VP.n44 VP.n43 161.3
R2267 VP.n79 VP.n78 161.3
R2268 VP.n77 VP.n1 161.3
R2269 VP.n76 VP.n75 161.3
R2270 VP.n74 VP.n2 161.3
R2271 VP.n73 VP.n72 161.3
R2272 VP.n71 VP.n3 161.3
R2273 VP.n70 VP.n69 161.3
R2274 VP.n68 VP.n67 161.3
R2275 VP.n66 VP.n5 161.3
R2276 VP.n65 VP.n64 161.3
R2277 VP.n63 VP.n6 161.3
R2278 VP.n62 VP.n61 161.3
R2279 VP.n60 VP.n7 161.3
R2280 VP.n59 VP.n58 161.3
R2281 VP.n57 VP.n56 161.3
R2282 VP.n55 VP.n9 161.3
R2283 VP.n54 VP.n53 161.3
R2284 VP.n52 VP.n10 161.3
R2285 VP.n51 VP.n50 161.3
R2286 VP.n49 VP.n11 161.3
R2287 VP.n48 VP.n47 161.3
R2288 VP.n22 VP.t1 123.871
R2289 VP.n12 VP.t6 90.862
R2290 VP.n8 VP.t5 90.862
R2291 VP.n4 VP.t7 90.862
R2292 VP.n0 VP.t4 90.862
R2293 VP.n13 VP.t0 90.862
R2294 VP.n17 VP.t2 90.862
R2295 VP.n21 VP.t3 90.862
R2296 VP.n46 VP.n12 74.0678
R2297 VP.n80 VP.n0 74.0678
R2298 VP.n45 VP.n13 74.0678
R2299 VP.n22 VP.n21 60.6108
R2300 VP.n46 VP.n45 54.0143
R2301 VP.n50 VP.n10 45.2793
R2302 VP.n76 VP.n2 45.2793
R2303 VP.n41 VP.n15 45.2793
R2304 VP.n61 VP.n6 40.4106
R2305 VP.n65 VP.n6 40.4106
R2306 VP.n30 VP.n19 40.4106
R2307 VP.n26 VP.n19 40.4106
R2308 VP.n54 VP.n10 35.5419
R2309 VP.n72 VP.n2 35.5419
R2310 VP.n37 VP.n15 35.5419
R2311 VP.n49 VP.n48 24.3439
R2312 VP.n50 VP.n49 24.3439
R2313 VP.n55 VP.n54 24.3439
R2314 VP.n56 VP.n55 24.3439
R2315 VP.n60 VP.n59 24.3439
R2316 VP.n61 VP.n60 24.3439
R2317 VP.n66 VP.n65 24.3439
R2318 VP.n67 VP.n66 24.3439
R2319 VP.n71 VP.n70 24.3439
R2320 VP.n72 VP.n71 24.3439
R2321 VP.n77 VP.n76 24.3439
R2322 VP.n78 VP.n77 24.3439
R2323 VP.n42 VP.n41 24.3439
R2324 VP.n43 VP.n42 24.3439
R2325 VP.n31 VP.n30 24.3439
R2326 VP.n32 VP.n31 24.3439
R2327 VP.n36 VP.n35 24.3439
R2328 VP.n37 VP.n36 24.3439
R2329 VP.n25 VP.n24 24.3439
R2330 VP.n26 VP.n25 24.3439
R2331 VP.n48 VP.n12 15.8237
R2332 VP.n78 VP.n0 15.8237
R2333 VP.n43 VP.n13 15.8237
R2334 VP.n59 VP.n8 13.3894
R2335 VP.n67 VP.n4 13.3894
R2336 VP.n32 VP.n17 13.3894
R2337 VP.n24 VP.n21 13.3894
R2338 VP.n56 VP.n8 10.955
R2339 VP.n70 VP.n4 10.955
R2340 VP.n35 VP.n17 10.955
R2341 VP.n23 VP.n22 4.11423
R2342 VP.n45 VP.n44 0.355081
R2343 VP.n47 VP.n46 0.355081
R2344 VP.n80 VP.n79 0.355081
R2345 VP VP.n80 0.26685
R2346 VP.n23 VP.n20 0.189894
R2347 VP.n27 VP.n20 0.189894
R2348 VP.n28 VP.n27 0.189894
R2349 VP.n29 VP.n28 0.189894
R2350 VP.n29 VP.n18 0.189894
R2351 VP.n33 VP.n18 0.189894
R2352 VP.n34 VP.n33 0.189894
R2353 VP.n34 VP.n16 0.189894
R2354 VP.n38 VP.n16 0.189894
R2355 VP.n39 VP.n38 0.189894
R2356 VP.n40 VP.n39 0.189894
R2357 VP.n40 VP.n14 0.189894
R2358 VP.n44 VP.n14 0.189894
R2359 VP.n47 VP.n11 0.189894
R2360 VP.n51 VP.n11 0.189894
R2361 VP.n52 VP.n51 0.189894
R2362 VP.n53 VP.n52 0.189894
R2363 VP.n53 VP.n9 0.189894
R2364 VP.n57 VP.n9 0.189894
R2365 VP.n58 VP.n57 0.189894
R2366 VP.n58 VP.n7 0.189894
R2367 VP.n62 VP.n7 0.189894
R2368 VP.n63 VP.n62 0.189894
R2369 VP.n64 VP.n63 0.189894
R2370 VP.n64 VP.n5 0.189894
R2371 VP.n68 VP.n5 0.189894
R2372 VP.n69 VP.n68 0.189894
R2373 VP.n69 VP.n3 0.189894
R2374 VP.n73 VP.n3 0.189894
R2375 VP.n74 VP.n73 0.189894
R2376 VP.n75 VP.n74 0.189894
R2377 VP.n75 VP.n1 0.189894
R2378 VP.n79 VP.n1 0.189894
R2379 VDD1 VDD1.n0 75.8155
R2380 VDD1.n3 VDD1.n2 75.7017
R2381 VDD1.n3 VDD1.n1 75.7017
R2382 VDD1.n5 VDD1.n4 74.2269
R2383 VDD1.n5 VDD1.n3 48.5354
R2384 VDD1.n4 VDD1.t5 2.67801
R2385 VDD1.n4 VDD1.t7 2.67801
R2386 VDD1.n0 VDD1.t6 2.67801
R2387 VDD1.n0 VDD1.t4 2.67801
R2388 VDD1.n2 VDD1.t0 2.67801
R2389 VDD1.n2 VDD1.t3 2.67801
R2390 VDD1.n1 VDD1.t1 2.67801
R2391 VDD1.n1 VDD1.t2 2.67801
R2392 VDD1 VDD1.n5 1.47248
C0 VDD1 VN 0.152218f
C1 VTAIL w_n4520_n3396# 4.28866f
C2 VTAIL B 5.29679f
C3 VDD2 VN 9.136451f
C4 VN w_n4520_n3396# 9.39414f
C5 VTAIL VP 9.74692f
C6 VN B 1.36686f
C7 VN VP 8.4552f
C8 VN VTAIL 9.732821f
C9 VDD1 VDD2 2.09833f
C10 VDD1 w_n4520_n3396# 2.15407f
C11 VDD1 B 1.84202f
C12 VDD2 w_n4520_n3396# 2.29479f
C13 VDD2 B 1.95755f
C14 VDD1 VP 9.56754f
C15 w_n4520_n3396# B 11.1038f
C16 VDD2 VP 0.585014f
C17 VDD1 VTAIL 8.3289f
C18 w_n4520_n3396# VP 9.98276f
C19 B VP 2.35689f
C20 VDD2 VTAIL 8.387469f
C21 VDD2 VSUBS 2.19994f
C22 VDD1 VSUBS 2.96092f
C23 VTAIL VSUBS 1.453178f
C24 VN VSUBS 7.57256f
C25 VP VSUBS 4.23263f
C26 B VSUBS 5.707046f
C27 w_n4520_n3396# VSUBS 0.188918p
C28 VDD1.t6 VSUBS 0.291804f
C29 VDD1.t4 VSUBS 0.291804f
C30 VDD1.n0 VSUBS 2.3044f
C31 VDD1.t1 VSUBS 0.291804f
C32 VDD1.t2 VSUBS 0.291804f
C33 VDD1.n1 VSUBS 2.30266f
C34 VDD1.t0 VSUBS 0.291804f
C35 VDD1.t3 VSUBS 0.291804f
C36 VDD1.n2 VSUBS 2.30266f
C37 VDD1.n3 VSUBS 5.13275f
C38 VDD1.t5 VSUBS 0.291804f
C39 VDD1.t7 VSUBS 0.291804f
C40 VDD1.n4 VSUBS 2.28262f
C41 VDD1.n5 VSUBS 4.2231f
C42 VP.t4 VSUBS 3.02248f
C43 VP.n0 VSUBS 1.17429f
C44 VP.n1 VSUBS 0.028369f
C45 VP.n2 VSUBS 0.023888f
C46 VP.n3 VSUBS 0.028369f
C47 VP.t7 VSUBS 3.02248f
C48 VP.n4 VSUBS 1.06217f
C49 VP.n5 VSUBS 0.028369f
C50 VP.n6 VSUBS 0.022956f
C51 VP.n7 VSUBS 0.028369f
C52 VP.t5 VSUBS 3.02248f
C53 VP.n8 VSUBS 1.06217f
C54 VP.n9 VSUBS 0.028369f
C55 VP.n10 VSUBS 0.023888f
C56 VP.n11 VSUBS 0.028369f
C57 VP.t6 VSUBS 3.02248f
C58 VP.n12 VSUBS 1.17429f
C59 VP.t0 VSUBS 3.02248f
C60 VP.n13 VSUBS 1.17429f
C61 VP.n14 VSUBS 0.028369f
C62 VP.n15 VSUBS 0.023888f
C63 VP.n16 VSUBS 0.028369f
C64 VP.t2 VSUBS 3.02248f
C65 VP.n17 VSUBS 1.06217f
C66 VP.n18 VSUBS 0.028369f
C67 VP.n19 VSUBS 0.022956f
C68 VP.n20 VSUBS 0.028369f
C69 VP.t3 VSUBS 3.02248f
C70 VP.n21 VSUBS 1.15762f
C71 VP.t1 VSUBS 3.35954f
C72 VP.n22 VSUBS 1.10508f
C73 VP.n23 VSUBS 0.33015f
C74 VP.n24 VSUBS 0.041331f
C75 VP.n25 VSUBS 0.053137f
C76 VP.n26 VSUBS 0.056684f
C77 VP.n27 VSUBS 0.028369f
C78 VP.n28 VSUBS 0.028369f
C79 VP.n29 VSUBS 0.028369f
C80 VP.n30 VSUBS 0.056684f
C81 VP.n31 VSUBS 0.053137f
C82 VP.n32 VSUBS 0.041331f
C83 VP.n33 VSUBS 0.028369f
C84 VP.n34 VSUBS 0.028369f
C85 VP.n35 VSUBS 0.038707f
C86 VP.n36 VSUBS 0.053137f
C87 VP.n37 VSUBS 0.057601f
C88 VP.n38 VSUBS 0.028369f
C89 VP.n39 VSUBS 0.028369f
C90 VP.n40 VSUBS 0.028369f
C91 VP.n41 VSUBS 0.054835f
C92 VP.n42 VSUBS 0.053137f
C93 VP.n43 VSUBS 0.043955f
C94 VP.n44 VSUBS 0.045794f
C95 VP.n45 VSUBS 1.79755f
C96 VP.n46 VSUBS 1.81638f
C97 VP.n47 VSUBS 0.045794f
C98 VP.n48 VSUBS 0.043955f
C99 VP.n49 VSUBS 0.053137f
C100 VP.n50 VSUBS 0.054835f
C101 VP.n51 VSUBS 0.028369f
C102 VP.n52 VSUBS 0.028369f
C103 VP.n53 VSUBS 0.028369f
C104 VP.n54 VSUBS 0.057601f
C105 VP.n55 VSUBS 0.053137f
C106 VP.n56 VSUBS 0.038707f
C107 VP.n57 VSUBS 0.028369f
C108 VP.n58 VSUBS 0.028369f
C109 VP.n59 VSUBS 0.041331f
C110 VP.n60 VSUBS 0.053137f
C111 VP.n61 VSUBS 0.056684f
C112 VP.n62 VSUBS 0.028369f
C113 VP.n63 VSUBS 0.028369f
C114 VP.n64 VSUBS 0.028369f
C115 VP.n65 VSUBS 0.056684f
C116 VP.n66 VSUBS 0.053137f
C117 VP.n67 VSUBS 0.041331f
C118 VP.n68 VSUBS 0.028369f
C119 VP.n69 VSUBS 0.028369f
C120 VP.n70 VSUBS 0.038707f
C121 VP.n71 VSUBS 0.053137f
C122 VP.n72 VSUBS 0.057601f
C123 VP.n73 VSUBS 0.028369f
C124 VP.n74 VSUBS 0.028369f
C125 VP.n75 VSUBS 0.028369f
C126 VP.n76 VSUBS 0.054835f
C127 VP.n77 VSUBS 0.053137f
C128 VP.n78 VSUBS 0.043955f
C129 VP.n79 VSUBS 0.045794f
C130 VP.n80 VSUBS 0.06638f
C131 VTAIL.t10 VSUBS 0.245176f
C132 VTAIL.t8 VSUBS 0.245176f
C133 VTAIL.n0 VSUBS 1.78016f
C134 VTAIL.n1 VSUBS 0.839833f
C135 VTAIL.n2 VSUBS 0.028191f
C136 VTAIL.n3 VSUBS 0.025557f
C137 VTAIL.n4 VSUBS 0.013733f
C138 VTAIL.n5 VSUBS 0.03246f
C139 VTAIL.n6 VSUBS 0.014541f
C140 VTAIL.n7 VSUBS 0.025557f
C141 VTAIL.n8 VSUBS 0.013733f
C142 VTAIL.n9 VSUBS 0.03246f
C143 VTAIL.n10 VSUBS 0.014541f
C144 VTAIL.n11 VSUBS 0.025557f
C145 VTAIL.n12 VSUBS 0.014137f
C146 VTAIL.n13 VSUBS 0.03246f
C147 VTAIL.n14 VSUBS 0.014541f
C148 VTAIL.n15 VSUBS 0.025557f
C149 VTAIL.n16 VSUBS 0.013733f
C150 VTAIL.n17 VSUBS 0.03246f
C151 VTAIL.n18 VSUBS 0.014541f
C152 VTAIL.n19 VSUBS 0.025557f
C153 VTAIL.n20 VSUBS 0.013733f
C154 VTAIL.n21 VSUBS 0.024345f
C155 VTAIL.n22 VSUBS 0.024418f
C156 VTAIL.t11 VSUBS 0.06996f
C157 VTAIL.n23 VSUBS 0.202893f
C158 VTAIL.n24 VSUBS 1.27136f
C159 VTAIL.n25 VSUBS 0.013733f
C160 VTAIL.n26 VSUBS 0.014541f
C161 VTAIL.n27 VSUBS 0.03246f
C162 VTAIL.n28 VSUBS 0.03246f
C163 VTAIL.n29 VSUBS 0.014541f
C164 VTAIL.n30 VSUBS 0.013733f
C165 VTAIL.n31 VSUBS 0.025557f
C166 VTAIL.n32 VSUBS 0.025557f
C167 VTAIL.n33 VSUBS 0.013733f
C168 VTAIL.n34 VSUBS 0.014541f
C169 VTAIL.n35 VSUBS 0.03246f
C170 VTAIL.n36 VSUBS 0.03246f
C171 VTAIL.n37 VSUBS 0.014541f
C172 VTAIL.n38 VSUBS 0.013733f
C173 VTAIL.n39 VSUBS 0.025557f
C174 VTAIL.n40 VSUBS 0.025557f
C175 VTAIL.n41 VSUBS 0.013733f
C176 VTAIL.n42 VSUBS 0.013733f
C177 VTAIL.n43 VSUBS 0.014541f
C178 VTAIL.n44 VSUBS 0.03246f
C179 VTAIL.n45 VSUBS 0.03246f
C180 VTAIL.n46 VSUBS 0.03246f
C181 VTAIL.n47 VSUBS 0.014137f
C182 VTAIL.n48 VSUBS 0.013733f
C183 VTAIL.n49 VSUBS 0.025557f
C184 VTAIL.n50 VSUBS 0.025557f
C185 VTAIL.n51 VSUBS 0.013733f
C186 VTAIL.n52 VSUBS 0.014541f
C187 VTAIL.n53 VSUBS 0.03246f
C188 VTAIL.n54 VSUBS 0.03246f
C189 VTAIL.n55 VSUBS 0.014541f
C190 VTAIL.n56 VSUBS 0.013733f
C191 VTAIL.n57 VSUBS 0.025557f
C192 VTAIL.n58 VSUBS 0.025557f
C193 VTAIL.n59 VSUBS 0.013733f
C194 VTAIL.n60 VSUBS 0.014541f
C195 VTAIL.n61 VSUBS 0.03246f
C196 VTAIL.n62 VSUBS 0.078956f
C197 VTAIL.n63 VSUBS 0.014541f
C198 VTAIL.n64 VSUBS 0.013733f
C199 VTAIL.n65 VSUBS 0.059772f
C200 VTAIL.n66 VSUBS 0.039744f
C201 VTAIL.n67 VSUBS 0.31293f
C202 VTAIL.n68 VSUBS 0.028191f
C203 VTAIL.n69 VSUBS 0.025557f
C204 VTAIL.n70 VSUBS 0.013733f
C205 VTAIL.n71 VSUBS 0.03246f
C206 VTAIL.n72 VSUBS 0.014541f
C207 VTAIL.n73 VSUBS 0.025557f
C208 VTAIL.n74 VSUBS 0.013733f
C209 VTAIL.n75 VSUBS 0.03246f
C210 VTAIL.n76 VSUBS 0.014541f
C211 VTAIL.n77 VSUBS 0.025557f
C212 VTAIL.n78 VSUBS 0.014137f
C213 VTAIL.n79 VSUBS 0.03246f
C214 VTAIL.n80 VSUBS 0.014541f
C215 VTAIL.n81 VSUBS 0.025557f
C216 VTAIL.n82 VSUBS 0.013733f
C217 VTAIL.n83 VSUBS 0.03246f
C218 VTAIL.n84 VSUBS 0.014541f
C219 VTAIL.n85 VSUBS 0.025557f
C220 VTAIL.n86 VSUBS 0.013733f
C221 VTAIL.n87 VSUBS 0.024345f
C222 VTAIL.n88 VSUBS 0.024418f
C223 VTAIL.t15 VSUBS 0.06996f
C224 VTAIL.n89 VSUBS 0.202893f
C225 VTAIL.n90 VSUBS 1.27136f
C226 VTAIL.n91 VSUBS 0.013733f
C227 VTAIL.n92 VSUBS 0.014541f
C228 VTAIL.n93 VSUBS 0.03246f
C229 VTAIL.n94 VSUBS 0.03246f
C230 VTAIL.n95 VSUBS 0.014541f
C231 VTAIL.n96 VSUBS 0.013733f
C232 VTAIL.n97 VSUBS 0.025557f
C233 VTAIL.n98 VSUBS 0.025557f
C234 VTAIL.n99 VSUBS 0.013733f
C235 VTAIL.n100 VSUBS 0.014541f
C236 VTAIL.n101 VSUBS 0.03246f
C237 VTAIL.n102 VSUBS 0.03246f
C238 VTAIL.n103 VSUBS 0.014541f
C239 VTAIL.n104 VSUBS 0.013733f
C240 VTAIL.n105 VSUBS 0.025557f
C241 VTAIL.n106 VSUBS 0.025557f
C242 VTAIL.n107 VSUBS 0.013733f
C243 VTAIL.n108 VSUBS 0.013733f
C244 VTAIL.n109 VSUBS 0.014541f
C245 VTAIL.n110 VSUBS 0.03246f
C246 VTAIL.n111 VSUBS 0.03246f
C247 VTAIL.n112 VSUBS 0.03246f
C248 VTAIL.n113 VSUBS 0.014137f
C249 VTAIL.n114 VSUBS 0.013733f
C250 VTAIL.n115 VSUBS 0.025557f
C251 VTAIL.n116 VSUBS 0.025557f
C252 VTAIL.n117 VSUBS 0.013733f
C253 VTAIL.n118 VSUBS 0.014541f
C254 VTAIL.n119 VSUBS 0.03246f
C255 VTAIL.n120 VSUBS 0.03246f
C256 VTAIL.n121 VSUBS 0.014541f
C257 VTAIL.n122 VSUBS 0.013733f
C258 VTAIL.n123 VSUBS 0.025557f
C259 VTAIL.n124 VSUBS 0.025557f
C260 VTAIL.n125 VSUBS 0.013733f
C261 VTAIL.n126 VSUBS 0.014541f
C262 VTAIL.n127 VSUBS 0.03246f
C263 VTAIL.n128 VSUBS 0.078956f
C264 VTAIL.n129 VSUBS 0.014541f
C265 VTAIL.n130 VSUBS 0.013733f
C266 VTAIL.n131 VSUBS 0.059772f
C267 VTAIL.n132 VSUBS 0.039744f
C268 VTAIL.n133 VSUBS 0.31293f
C269 VTAIL.t2 VSUBS 0.245176f
C270 VTAIL.t1 VSUBS 0.245176f
C271 VTAIL.n134 VSUBS 1.78016f
C272 VTAIL.n135 VSUBS 1.08706f
C273 VTAIL.n136 VSUBS 0.028191f
C274 VTAIL.n137 VSUBS 0.025557f
C275 VTAIL.n138 VSUBS 0.013733f
C276 VTAIL.n139 VSUBS 0.03246f
C277 VTAIL.n140 VSUBS 0.014541f
C278 VTAIL.n141 VSUBS 0.025557f
C279 VTAIL.n142 VSUBS 0.013733f
C280 VTAIL.n143 VSUBS 0.03246f
C281 VTAIL.n144 VSUBS 0.014541f
C282 VTAIL.n145 VSUBS 0.025557f
C283 VTAIL.n146 VSUBS 0.014137f
C284 VTAIL.n147 VSUBS 0.03246f
C285 VTAIL.n148 VSUBS 0.014541f
C286 VTAIL.n149 VSUBS 0.025557f
C287 VTAIL.n150 VSUBS 0.013733f
C288 VTAIL.n151 VSUBS 0.03246f
C289 VTAIL.n152 VSUBS 0.014541f
C290 VTAIL.n153 VSUBS 0.025557f
C291 VTAIL.n154 VSUBS 0.013733f
C292 VTAIL.n155 VSUBS 0.024345f
C293 VTAIL.n156 VSUBS 0.024418f
C294 VTAIL.t0 VSUBS 0.06996f
C295 VTAIL.n157 VSUBS 0.202893f
C296 VTAIL.n158 VSUBS 1.27136f
C297 VTAIL.n159 VSUBS 0.013733f
C298 VTAIL.n160 VSUBS 0.014541f
C299 VTAIL.n161 VSUBS 0.03246f
C300 VTAIL.n162 VSUBS 0.03246f
C301 VTAIL.n163 VSUBS 0.014541f
C302 VTAIL.n164 VSUBS 0.013733f
C303 VTAIL.n165 VSUBS 0.025557f
C304 VTAIL.n166 VSUBS 0.025557f
C305 VTAIL.n167 VSUBS 0.013733f
C306 VTAIL.n168 VSUBS 0.014541f
C307 VTAIL.n169 VSUBS 0.03246f
C308 VTAIL.n170 VSUBS 0.03246f
C309 VTAIL.n171 VSUBS 0.014541f
C310 VTAIL.n172 VSUBS 0.013733f
C311 VTAIL.n173 VSUBS 0.025557f
C312 VTAIL.n174 VSUBS 0.025557f
C313 VTAIL.n175 VSUBS 0.013733f
C314 VTAIL.n176 VSUBS 0.013733f
C315 VTAIL.n177 VSUBS 0.014541f
C316 VTAIL.n178 VSUBS 0.03246f
C317 VTAIL.n179 VSUBS 0.03246f
C318 VTAIL.n180 VSUBS 0.03246f
C319 VTAIL.n181 VSUBS 0.014137f
C320 VTAIL.n182 VSUBS 0.013733f
C321 VTAIL.n183 VSUBS 0.025557f
C322 VTAIL.n184 VSUBS 0.025557f
C323 VTAIL.n185 VSUBS 0.013733f
C324 VTAIL.n186 VSUBS 0.014541f
C325 VTAIL.n187 VSUBS 0.03246f
C326 VTAIL.n188 VSUBS 0.03246f
C327 VTAIL.n189 VSUBS 0.014541f
C328 VTAIL.n190 VSUBS 0.013733f
C329 VTAIL.n191 VSUBS 0.025557f
C330 VTAIL.n192 VSUBS 0.025557f
C331 VTAIL.n193 VSUBS 0.013733f
C332 VTAIL.n194 VSUBS 0.014541f
C333 VTAIL.n195 VSUBS 0.03246f
C334 VTAIL.n196 VSUBS 0.078956f
C335 VTAIL.n197 VSUBS 0.014541f
C336 VTAIL.n198 VSUBS 0.013733f
C337 VTAIL.n199 VSUBS 0.059772f
C338 VTAIL.n200 VSUBS 0.039744f
C339 VTAIL.n201 VSUBS 1.73525f
C340 VTAIL.n202 VSUBS 0.028191f
C341 VTAIL.n203 VSUBS 0.025557f
C342 VTAIL.n204 VSUBS 0.013733f
C343 VTAIL.n205 VSUBS 0.03246f
C344 VTAIL.n206 VSUBS 0.014541f
C345 VTAIL.n207 VSUBS 0.025557f
C346 VTAIL.n208 VSUBS 0.013733f
C347 VTAIL.n209 VSUBS 0.03246f
C348 VTAIL.n210 VSUBS 0.014541f
C349 VTAIL.n211 VSUBS 0.025557f
C350 VTAIL.n212 VSUBS 0.014137f
C351 VTAIL.n213 VSUBS 0.03246f
C352 VTAIL.n214 VSUBS 0.013733f
C353 VTAIL.n215 VSUBS 0.014541f
C354 VTAIL.n216 VSUBS 0.025557f
C355 VTAIL.n217 VSUBS 0.013733f
C356 VTAIL.n218 VSUBS 0.03246f
C357 VTAIL.n219 VSUBS 0.014541f
C358 VTAIL.n220 VSUBS 0.025557f
C359 VTAIL.n221 VSUBS 0.013733f
C360 VTAIL.n222 VSUBS 0.024345f
C361 VTAIL.n223 VSUBS 0.024418f
C362 VTAIL.t13 VSUBS 0.06996f
C363 VTAIL.n224 VSUBS 0.202893f
C364 VTAIL.n225 VSUBS 1.27136f
C365 VTAIL.n226 VSUBS 0.013733f
C366 VTAIL.n227 VSUBS 0.014541f
C367 VTAIL.n228 VSUBS 0.03246f
C368 VTAIL.n229 VSUBS 0.03246f
C369 VTAIL.n230 VSUBS 0.014541f
C370 VTAIL.n231 VSUBS 0.013733f
C371 VTAIL.n232 VSUBS 0.025557f
C372 VTAIL.n233 VSUBS 0.025557f
C373 VTAIL.n234 VSUBS 0.013733f
C374 VTAIL.n235 VSUBS 0.014541f
C375 VTAIL.n236 VSUBS 0.03246f
C376 VTAIL.n237 VSUBS 0.03246f
C377 VTAIL.n238 VSUBS 0.014541f
C378 VTAIL.n239 VSUBS 0.013733f
C379 VTAIL.n240 VSUBS 0.025557f
C380 VTAIL.n241 VSUBS 0.025557f
C381 VTAIL.n242 VSUBS 0.013733f
C382 VTAIL.n243 VSUBS 0.014541f
C383 VTAIL.n244 VSUBS 0.03246f
C384 VTAIL.n245 VSUBS 0.03246f
C385 VTAIL.n246 VSUBS 0.03246f
C386 VTAIL.n247 VSUBS 0.014137f
C387 VTAIL.n248 VSUBS 0.013733f
C388 VTAIL.n249 VSUBS 0.025557f
C389 VTAIL.n250 VSUBS 0.025557f
C390 VTAIL.n251 VSUBS 0.013733f
C391 VTAIL.n252 VSUBS 0.014541f
C392 VTAIL.n253 VSUBS 0.03246f
C393 VTAIL.n254 VSUBS 0.03246f
C394 VTAIL.n255 VSUBS 0.014541f
C395 VTAIL.n256 VSUBS 0.013733f
C396 VTAIL.n257 VSUBS 0.025557f
C397 VTAIL.n258 VSUBS 0.025557f
C398 VTAIL.n259 VSUBS 0.013733f
C399 VTAIL.n260 VSUBS 0.014541f
C400 VTAIL.n261 VSUBS 0.03246f
C401 VTAIL.n262 VSUBS 0.078956f
C402 VTAIL.n263 VSUBS 0.014541f
C403 VTAIL.n264 VSUBS 0.013733f
C404 VTAIL.n265 VSUBS 0.059772f
C405 VTAIL.n266 VSUBS 0.039744f
C406 VTAIL.n267 VSUBS 1.73525f
C407 VTAIL.t9 VSUBS 0.245176f
C408 VTAIL.t14 VSUBS 0.245176f
C409 VTAIL.n268 VSUBS 1.78017f
C410 VTAIL.n269 VSUBS 1.08705f
C411 VTAIL.n270 VSUBS 0.028191f
C412 VTAIL.n271 VSUBS 0.025557f
C413 VTAIL.n272 VSUBS 0.013733f
C414 VTAIL.n273 VSUBS 0.03246f
C415 VTAIL.n274 VSUBS 0.014541f
C416 VTAIL.n275 VSUBS 0.025557f
C417 VTAIL.n276 VSUBS 0.013733f
C418 VTAIL.n277 VSUBS 0.03246f
C419 VTAIL.n278 VSUBS 0.014541f
C420 VTAIL.n279 VSUBS 0.025557f
C421 VTAIL.n280 VSUBS 0.014137f
C422 VTAIL.n281 VSUBS 0.03246f
C423 VTAIL.n282 VSUBS 0.013733f
C424 VTAIL.n283 VSUBS 0.014541f
C425 VTAIL.n284 VSUBS 0.025557f
C426 VTAIL.n285 VSUBS 0.013733f
C427 VTAIL.n286 VSUBS 0.03246f
C428 VTAIL.n287 VSUBS 0.014541f
C429 VTAIL.n288 VSUBS 0.025557f
C430 VTAIL.n289 VSUBS 0.013733f
C431 VTAIL.n290 VSUBS 0.024345f
C432 VTAIL.n291 VSUBS 0.024418f
C433 VTAIL.t12 VSUBS 0.06996f
C434 VTAIL.n292 VSUBS 0.202893f
C435 VTAIL.n293 VSUBS 1.27136f
C436 VTAIL.n294 VSUBS 0.013733f
C437 VTAIL.n295 VSUBS 0.014541f
C438 VTAIL.n296 VSUBS 0.03246f
C439 VTAIL.n297 VSUBS 0.03246f
C440 VTAIL.n298 VSUBS 0.014541f
C441 VTAIL.n299 VSUBS 0.013733f
C442 VTAIL.n300 VSUBS 0.025557f
C443 VTAIL.n301 VSUBS 0.025557f
C444 VTAIL.n302 VSUBS 0.013733f
C445 VTAIL.n303 VSUBS 0.014541f
C446 VTAIL.n304 VSUBS 0.03246f
C447 VTAIL.n305 VSUBS 0.03246f
C448 VTAIL.n306 VSUBS 0.014541f
C449 VTAIL.n307 VSUBS 0.013733f
C450 VTAIL.n308 VSUBS 0.025557f
C451 VTAIL.n309 VSUBS 0.025557f
C452 VTAIL.n310 VSUBS 0.013733f
C453 VTAIL.n311 VSUBS 0.014541f
C454 VTAIL.n312 VSUBS 0.03246f
C455 VTAIL.n313 VSUBS 0.03246f
C456 VTAIL.n314 VSUBS 0.03246f
C457 VTAIL.n315 VSUBS 0.014137f
C458 VTAIL.n316 VSUBS 0.013733f
C459 VTAIL.n317 VSUBS 0.025557f
C460 VTAIL.n318 VSUBS 0.025557f
C461 VTAIL.n319 VSUBS 0.013733f
C462 VTAIL.n320 VSUBS 0.014541f
C463 VTAIL.n321 VSUBS 0.03246f
C464 VTAIL.n322 VSUBS 0.03246f
C465 VTAIL.n323 VSUBS 0.014541f
C466 VTAIL.n324 VSUBS 0.013733f
C467 VTAIL.n325 VSUBS 0.025557f
C468 VTAIL.n326 VSUBS 0.025557f
C469 VTAIL.n327 VSUBS 0.013733f
C470 VTAIL.n328 VSUBS 0.014541f
C471 VTAIL.n329 VSUBS 0.03246f
C472 VTAIL.n330 VSUBS 0.078956f
C473 VTAIL.n331 VSUBS 0.014541f
C474 VTAIL.n332 VSUBS 0.013733f
C475 VTAIL.n333 VSUBS 0.059772f
C476 VTAIL.n334 VSUBS 0.039744f
C477 VTAIL.n335 VSUBS 0.31293f
C478 VTAIL.n336 VSUBS 0.028191f
C479 VTAIL.n337 VSUBS 0.025557f
C480 VTAIL.n338 VSUBS 0.013733f
C481 VTAIL.n339 VSUBS 0.03246f
C482 VTAIL.n340 VSUBS 0.014541f
C483 VTAIL.n341 VSUBS 0.025557f
C484 VTAIL.n342 VSUBS 0.013733f
C485 VTAIL.n343 VSUBS 0.03246f
C486 VTAIL.n344 VSUBS 0.014541f
C487 VTAIL.n345 VSUBS 0.025557f
C488 VTAIL.n346 VSUBS 0.014137f
C489 VTAIL.n347 VSUBS 0.03246f
C490 VTAIL.n348 VSUBS 0.013733f
C491 VTAIL.n349 VSUBS 0.014541f
C492 VTAIL.n350 VSUBS 0.025557f
C493 VTAIL.n351 VSUBS 0.013733f
C494 VTAIL.n352 VSUBS 0.03246f
C495 VTAIL.n353 VSUBS 0.014541f
C496 VTAIL.n354 VSUBS 0.025557f
C497 VTAIL.n355 VSUBS 0.013733f
C498 VTAIL.n356 VSUBS 0.024345f
C499 VTAIL.n357 VSUBS 0.024418f
C500 VTAIL.t4 VSUBS 0.06996f
C501 VTAIL.n358 VSUBS 0.202893f
C502 VTAIL.n359 VSUBS 1.27136f
C503 VTAIL.n360 VSUBS 0.013733f
C504 VTAIL.n361 VSUBS 0.014541f
C505 VTAIL.n362 VSUBS 0.03246f
C506 VTAIL.n363 VSUBS 0.03246f
C507 VTAIL.n364 VSUBS 0.014541f
C508 VTAIL.n365 VSUBS 0.013733f
C509 VTAIL.n366 VSUBS 0.025557f
C510 VTAIL.n367 VSUBS 0.025557f
C511 VTAIL.n368 VSUBS 0.013733f
C512 VTAIL.n369 VSUBS 0.014541f
C513 VTAIL.n370 VSUBS 0.03246f
C514 VTAIL.n371 VSUBS 0.03246f
C515 VTAIL.n372 VSUBS 0.014541f
C516 VTAIL.n373 VSUBS 0.013733f
C517 VTAIL.n374 VSUBS 0.025557f
C518 VTAIL.n375 VSUBS 0.025557f
C519 VTAIL.n376 VSUBS 0.013733f
C520 VTAIL.n377 VSUBS 0.014541f
C521 VTAIL.n378 VSUBS 0.03246f
C522 VTAIL.n379 VSUBS 0.03246f
C523 VTAIL.n380 VSUBS 0.03246f
C524 VTAIL.n381 VSUBS 0.014137f
C525 VTAIL.n382 VSUBS 0.013733f
C526 VTAIL.n383 VSUBS 0.025557f
C527 VTAIL.n384 VSUBS 0.025557f
C528 VTAIL.n385 VSUBS 0.013733f
C529 VTAIL.n386 VSUBS 0.014541f
C530 VTAIL.n387 VSUBS 0.03246f
C531 VTAIL.n388 VSUBS 0.03246f
C532 VTAIL.n389 VSUBS 0.014541f
C533 VTAIL.n390 VSUBS 0.013733f
C534 VTAIL.n391 VSUBS 0.025557f
C535 VTAIL.n392 VSUBS 0.025557f
C536 VTAIL.n393 VSUBS 0.013733f
C537 VTAIL.n394 VSUBS 0.014541f
C538 VTAIL.n395 VSUBS 0.03246f
C539 VTAIL.n396 VSUBS 0.078956f
C540 VTAIL.n397 VSUBS 0.014541f
C541 VTAIL.n398 VSUBS 0.013733f
C542 VTAIL.n399 VSUBS 0.059772f
C543 VTAIL.n400 VSUBS 0.039744f
C544 VTAIL.n401 VSUBS 0.31293f
C545 VTAIL.t3 VSUBS 0.245176f
C546 VTAIL.t5 VSUBS 0.245176f
C547 VTAIL.n402 VSUBS 1.78017f
C548 VTAIL.n403 VSUBS 1.08705f
C549 VTAIL.n404 VSUBS 0.028191f
C550 VTAIL.n405 VSUBS 0.025557f
C551 VTAIL.n406 VSUBS 0.013733f
C552 VTAIL.n407 VSUBS 0.03246f
C553 VTAIL.n408 VSUBS 0.014541f
C554 VTAIL.n409 VSUBS 0.025557f
C555 VTAIL.n410 VSUBS 0.013733f
C556 VTAIL.n411 VSUBS 0.03246f
C557 VTAIL.n412 VSUBS 0.014541f
C558 VTAIL.n413 VSUBS 0.025557f
C559 VTAIL.n414 VSUBS 0.014137f
C560 VTAIL.n415 VSUBS 0.03246f
C561 VTAIL.n416 VSUBS 0.013733f
C562 VTAIL.n417 VSUBS 0.014541f
C563 VTAIL.n418 VSUBS 0.025557f
C564 VTAIL.n419 VSUBS 0.013733f
C565 VTAIL.n420 VSUBS 0.03246f
C566 VTAIL.n421 VSUBS 0.014541f
C567 VTAIL.n422 VSUBS 0.025557f
C568 VTAIL.n423 VSUBS 0.013733f
C569 VTAIL.n424 VSUBS 0.024345f
C570 VTAIL.n425 VSUBS 0.024418f
C571 VTAIL.t6 VSUBS 0.06996f
C572 VTAIL.n426 VSUBS 0.202893f
C573 VTAIL.n427 VSUBS 1.27136f
C574 VTAIL.n428 VSUBS 0.013733f
C575 VTAIL.n429 VSUBS 0.014541f
C576 VTAIL.n430 VSUBS 0.03246f
C577 VTAIL.n431 VSUBS 0.03246f
C578 VTAIL.n432 VSUBS 0.014541f
C579 VTAIL.n433 VSUBS 0.013733f
C580 VTAIL.n434 VSUBS 0.025557f
C581 VTAIL.n435 VSUBS 0.025557f
C582 VTAIL.n436 VSUBS 0.013733f
C583 VTAIL.n437 VSUBS 0.014541f
C584 VTAIL.n438 VSUBS 0.03246f
C585 VTAIL.n439 VSUBS 0.03246f
C586 VTAIL.n440 VSUBS 0.014541f
C587 VTAIL.n441 VSUBS 0.013733f
C588 VTAIL.n442 VSUBS 0.025557f
C589 VTAIL.n443 VSUBS 0.025557f
C590 VTAIL.n444 VSUBS 0.013733f
C591 VTAIL.n445 VSUBS 0.014541f
C592 VTAIL.n446 VSUBS 0.03246f
C593 VTAIL.n447 VSUBS 0.03246f
C594 VTAIL.n448 VSUBS 0.03246f
C595 VTAIL.n449 VSUBS 0.014137f
C596 VTAIL.n450 VSUBS 0.013733f
C597 VTAIL.n451 VSUBS 0.025557f
C598 VTAIL.n452 VSUBS 0.025557f
C599 VTAIL.n453 VSUBS 0.013733f
C600 VTAIL.n454 VSUBS 0.014541f
C601 VTAIL.n455 VSUBS 0.03246f
C602 VTAIL.n456 VSUBS 0.03246f
C603 VTAIL.n457 VSUBS 0.014541f
C604 VTAIL.n458 VSUBS 0.013733f
C605 VTAIL.n459 VSUBS 0.025557f
C606 VTAIL.n460 VSUBS 0.025557f
C607 VTAIL.n461 VSUBS 0.013733f
C608 VTAIL.n462 VSUBS 0.014541f
C609 VTAIL.n463 VSUBS 0.03246f
C610 VTAIL.n464 VSUBS 0.078956f
C611 VTAIL.n465 VSUBS 0.014541f
C612 VTAIL.n466 VSUBS 0.013733f
C613 VTAIL.n467 VSUBS 0.059772f
C614 VTAIL.n468 VSUBS 0.039744f
C615 VTAIL.n469 VSUBS 1.73525f
C616 VTAIL.n470 VSUBS 0.028191f
C617 VTAIL.n471 VSUBS 0.025557f
C618 VTAIL.n472 VSUBS 0.013733f
C619 VTAIL.n473 VSUBS 0.03246f
C620 VTAIL.n474 VSUBS 0.014541f
C621 VTAIL.n475 VSUBS 0.025557f
C622 VTAIL.n476 VSUBS 0.013733f
C623 VTAIL.n477 VSUBS 0.03246f
C624 VTAIL.n478 VSUBS 0.014541f
C625 VTAIL.n479 VSUBS 0.025557f
C626 VTAIL.n480 VSUBS 0.014137f
C627 VTAIL.n481 VSUBS 0.03246f
C628 VTAIL.n482 VSUBS 0.014541f
C629 VTAIL.n483 VSUBS 0.025557f
C630 VTAIL.n484 VSUBS 0.013733f
C631 VTAIL.n485 VSUBS 0.03246f
C632 VTAIL.n486 VSUBS 0.014541f
C633 VTAIL.n487 VSUBS 0.025557f
C634 VTAIL.n488 VSUBS 0.013733f
C635 VTAIL.n489 VSUBS 0.024345f
C636 VTAIL.n490 VSUBS 0.024418f
C637 VTAIL.t7 VSUBS 0.06996f
C638 VTAIL.n491 VSUBS 0.202893f
C639 VTAIL.n492 VSUBS 1.27136f
C640 VTAIL.n493 VSUBS 0.013733f
C641 VTAIL.n494 VSUBS 0.014541f
C642 VTAIL.n495 VSUBS 0.03246f
C643 VTAIL.n496 VSUBS 0.03246f
C644 VTAIL.n497 VSUBS 0.014541f
C645 VTAIL.n498 VSUBS 0.013733f
C646 VTAIL.n499 VSUBS 0.025557f
C647 VTAIL.n500 VSUBS 0.025557f
C648 VTAIL.n501 VSUBS 0.013733f
C649 VTAIL.n502 VSUBS 0.014541f
C650 VTAIL.n503 VSUBS 0.03246f
C651 VTAIL.n504 VSUBS 0.03246f
C652 VTAIL.n505 VSUBS 0.014541f
C653 VTAIL.n506 VSUBS 0.013733f
C654 VTAIL.n507 VSUBS 0.025557f
C655 VTAIL.n508 VSUBS 0.025557f
C656 VTAIL.n509 VSUBS 0.013733f
C657 VTAIL.n510 VSUBS 0.013733f
C658 VTAIL.n511 VSUBS 0.014541f
C659 VTAIL.n512 VSUBS 0.03246f
C660 VTAIL.n513 VSUBS 0.03246f
C661 VTAIL.n514 VSUBS 0.03246f
C662 VTAIL.n515 VSUBS 0.014137f
C663 VTAIL.n516 VSUBS 0.013733f
C664 VTAIL.n517 VSUBS 0.025557f
C665 VTAIL.n518 VSUBS 0.025557f
C666 VTAIL.n519 VSUBS 0.013733f
C667 VTAIL.n520 VSUBS 0.014541f
C668 VTAIL.n521 VSUBS 0.03246f
C669 VTAIL.n522 VSUBS 0.03246f
C670 VTAIL.n523 VSUBS 0.014541f
C671 VTAIL.n524 VSUBS 0.013733f
C672 VTAIL.n525 VSUBS 0.025557f
C673 VTAIL.n526 VSUBS 0.025557f
C674 VTAIL.n527 VSUBS 0.013733f
C675 VTAIL.n528 VSUBS 0.014541f
C676 VTAIL.n529 VSUBS 0.03246f
C677 VTAIL.n530 VSUBS 0.078956f
C678 VTAIL.n531 VSUBS 0.014541f
C679 VTAIL.n532 VSUBS 0.013733f
C680 VTAIL.n533 VSUBS 0.059772f
C681 VTAIL.n534 VSUBS 0.039744f
C682 VTAIL.n535 VSUBS 1.73046f
C683 VDD2.t6 VSUBS 0.289325f
C684 VDD2.t2 VSUBS 0.289325f
C685 VDD2.n0 VSUBS 2.2831f
C686 VDD2.t5 VSUBS 0.289325f
C687 VDD2.t1 VSUBS 0.289325f
C688 VDD2.n1 VSUBS 2.2831f
C689 VDD2.n2 VSUBS 5.02673f
C690 VDD2.t3 VSUBS 0.289325f
C691 VDD2.t0 VSUBS 0.289325f
C692 VDD2.n3 VSUBS 2.26324f
C693 VDD2.n4 VSUBS 4.14954f
C694 VDD2.t4 VSUBS 0.289325f
C695 VDD2.t7 VSUBS 0.289325f
C696 VDD2.n5 VSUBS 2.28304f
C697 VN.t7 VSUBS 2.75659f
C698 VN.n0 VSUBS 1.07099f
C699 VN.n1 VSUBS 0.025873f
C700 VN.n2 VSUBS 0.021786f
C701 VN.n3 VSUBS 0.025873f
C702 VN.t6 VSUBS 2.75659f
C703 VN.n4 VSUBS 0.968735f
C704 VN.n5 VSUBS 0.025873f
C705 VN.n6 VSUBS 0.020937f
C706 VN.n7 VSUBS 0.025873f
C707 VN.t4 VSUBS 2.75659f
C708 VN.n8 VSUBS 1.05578f
C709 VN.t3 VSUBS 3.064f
C710 VN.n9 VSUBS 1.00787f
C711 VN.n10 VSUBS 0.301106f
C712 VN.n11 VSUBS 0.037695f
C713 VN.n12 VSUBS 0.048463f
C714 VN.n13 VSUBS 0.051697f
C715 VN.n14 VSUBS 0.025873f
C716 VN.n15 VSUBS 0.025873f
C717 VN.n16 VSUBS 0.025873f
C718 VN.n17 VSUBS 0.051697f
C719 VN.n18 VSUBS 0.048463f
C720 VN.n19 VSUBS 0.037695f
C721 VN.n20 VSUBS 0.025873f
C722 VN.n21 VSUBS 0.025873f
C723 VN.n22 VSUBS 0.035302f
C724 VN.n23 VSUBS 0.048463f
C725 VN.n24 VSUBS 0.052534f
C726 VN.n25 VSUBS 0.025873f
C727 VN.n26 VSUBS 0.025873f
C728 VN.n27 VSUBS 0.025873f
C729 VN.n28 VSUBS 0.050012f
C730 VN.n29 VSUBS 0.048463f
C731 VN.n30 VSUBS 0.040088f
C732 VN.n31 VSUBS 0.041765f
C733 VN.n32 VSUBS 0.060541f
C734 VN.t1 VSUBS 2.75659f
C735 VN.n33 VSUBS 1.07099f
C736 VN.n34 VSUBS 0.025873f
C737 VN.n35 VSUBS 0.021786f
C738 VN.n36 VSUBS 0.025873f
C739 VN.t5 VSUBS 2.75659f
C740 VN.n37 VSUBS 0.968735f
C741 VN.n38 VSUBS 0.025873f
C742 VN.n39 VSUBS 0.020937f
C743 VN.n40 VSUBS 0.025873f
C744 VN.t0 VSUBS 2.75659f
C745 VN.n41 VSUBS 1.05578f
C746 VN.t2 VSUBS 3.064f
C747 VN.n42 VSUBS 1.00787f
C748 VN.n43 VSUBS 0.301106f
C749 VN.n44 VSUBS 0.037695f
C750 VN.n45 VSUBS 0.048463f
C751 VN.n46 VSUBS 0.051697f
C752 VN.n47 VSUBS 0.025873f
C753 VN.n48 VSUBS 0.025873f
C754 VN.n49 VSUBS 0.025873f
C755 VN.n50 VSUBS 0.051697f
C756 VN.n51 VSUBS 0.048463f
C757 VN.n52 VSUBS 0.037695f
C758 VN.n53 VSUBS 0.025873f
C759 VN.n54 VSUBS 0.025873f
C760 VN.n55 VSUBS 0.035302f
C761 VN.n56 VSUBS 0.048463f
C762 VN.n57 VSUBS 0.052534f
C763 VN.n58 VSUBS 0.025873f
C764 VN.n59 VSUBS 0.025873f
C765 VN.n60 VSUBS 0.025873f
C766 VN.n61 VSUBS 0.050012f
C767 VN.n62 VSUBS 0.048463f
C768 VN.n63 VSUBS 0.040088f
C769 VN.n64 VSUBS 0.041765f
C770 VN.n65 VSUBS 1.64974f
C771 B.n0 VSUBS 0.006467f
C772 B.n1 VSUBS 0.006467f
C773 B.n2 VSUBS 0.009564f
C774 B.n3 VSUBS 0.007329f
C775 B.n4 VSUBS 0.007329f
C776 B.n5 VSUBS 0.007329f
C777 B.n6 VSUBS 0.007329f
C778 B.n7 VSUBS 0.007329f
C779 B.n8 VSUBS 0.007329f
C780 B.n9 VSUBS 0.007329f
C781 B.n10 VSUBS 0.007329f
C782 B.n11 VSUBS 0.007329f
C783 B.n12 VSUBS 0.007329f
C784 B.n13 VSUBS 0.007329f
C785 B.n14 VSUBS 0.007329f
C786 B.n15 VSUBS 0.007329f
C787 B.n16 VSUBS 0.007329f
C788 B.n17 VSUBS 0.007329f
C789 B.n18 VSUBS 0.007329f
C790 B.n19 VSUBS 0.007329f
C791 B.n20 VSUBS 0.007329f
C792 B.n21 VSUBS 0.007329f
C793 B.n22 VSUBS 0.007329f
C794 B.n23 VSUBS 0.007329f
C795 B.n24 VSUBS 0.007329f
C796 B.n25 VSUBS 0.007329f
C797 B.n26 VSUBS 0.007329f
C798 B.n27 VSUBS 0.007329f
C799 B.n28 VSUBS 0.007329f
C800 B.n29 VSUBS 0.007329f
C801 B.n30 VSUBS 0.007329f
C802 B.n31 VSUBS 0.007329f
C803 B.n32 VSUBS 0.016207f
C804 B.n33 VSUBS 0.007329f
C805 B.n34 VSUBS 0.007329f
C806 B.n35 VSUBS 0.007329f
C807 B.n36 VSUBS 0.007329f
C808 B.n37 VSUBS 0.007329f
C809 B.n38 VSUBS 0.007329f
C810 B.n39 VSUBS 0.007329f
C811 B.n40 VSUBS 0.007329f
C812 B.n41 VSUBS 0.007329f
C813 B.n42 VSUBS 0.007329f
C814 B.n43 VSUBS 0.007329f
C815 B.n44 VSUBS 0.007329f
C816 B.n45 VSUBS 0.007329f
C817 B.n46 VSUBS 0.007329f
C818 B.n47 VSUBS 0.007329f
C819 B.n48 VSUBS 0.007329f
C820 B.n49 VSUBS 0.007329f
C821 B.n50 VSUBS 0.007329f
C822 B.n51 VSUBS 0.007329f
C823 B.n52 VSUBS 0.007329f
C824 B.n53 VSUBS 0.007329f
C825 B.t4 VSUBS 0.224329f
C826 B.t5 VSUBS 0.264035f
C827 B.t3 VSUBS 1.88903f
C828 B.n54 VSUBS 0.420943f
C829 B.n55 VSUBS 0.268296f
C830 B.n56 VSUBS 0.007329f
C831 B.n57 VSUBS 0.007329f
C832 B.n58 VSUBS 0.007329f
C833 B.n59 VSUBS 0.007329f
C834 B.t7 VSUBS 0.224332f
C835 B.t8 VSUBS 0.264037f
C836 B.t6 VSUBS 1.88903f
C837 B.n60 VSUBS 0.42094f
C838 B.n61 VSUBS 0.268293f
C839 B.n62 VSUBS 0.016981f
C840 B.n63 VSUBS 0.007329f
C841 B.n64 VSUBS 0.007329f
C842 B.n65 VSUBS 0.007329f
C843 B.n66 VSUBS 0.007329f
C844 B.n67 VSUBS 0.007329f
C845 B.n68 VSUBS 0.007329f
C846 B.n69 VSUBS 0.007329f
C847 B.n70 VSUBS 0.007329f
C848 B.n71 VSUBS 0.007329f
C849 B.n72 VSUBS 0.007329f
C850 B.n73 VSUBS 0.007329f
C851 B.n74 VSUBS 0.007329f
C852 B.n75 VSUBS 0.007329f
C853 B.n76 VSUBS 0.007329f
C854 B.n77 VSUBS 0.007329f
C855 B.n78 VSUBS 0.007329f
C856 B.n79 VSUBS 0.007329f
C857 B.n80 VSUBS 0.007329f
C858 B.n81 VSUBS 0.007329f
C859 B.n82 VSUBS 0.007329f
C860 B.n83 VSUBS 0.016207f
C861 B.n84 VSUBS 0.007329f
C862 B.n85 VSUBS 0.007329f
C863 B.n86 VSUBS 0.007329f
C864 B.n87 VSUBS 0.007329f
C865 B.n88 VSUBS 0.007329f
C866 B.n89 VSUBS 0.007329f
C867 B.n90 VSUBS 0.007329f
C868 B.n91 VSUBS 0.007329f
C869 B.n92 VSUBS 0.007329f
C870 B.n93 VSUBS 0.007329f
C871 B.n94 VSUBS 0.007329f
C872 B.n95 VSUBS 0.007329f
C873 B.n96 VSUBS 0.007329f
C874 B.n97 VSUBS 0.007329f
C875 B.n98 VSUBS 0.007329f
C876 B.n99 VSUBS 0.007329f
C877 B.n100 VSUBS 0.007329f
C878 B.n101 VSUBS 0.007329f
C879 B.n102 VSUBS 0.007329f
C880 B.n103 VSUBS 0.007329f
C881 B.n104 VSUBS 0.007329f
C882 B.n105 VSUBS 0.007329f
C883 B.n106 VSUBS 0.007329f
C884 B.n107 VSUBS 0.007329f
C885 B.n108 VSUBS 0.007329f
C886 B.n109 VSUBS 0.007329f
C887 B.n110 VSUBS 0.007329f
C888 B.n111 VSUBS 0.007329f
C889 B.n112 VSUBS 0.007329f
C890 B.n113 VSUBS 0.007329f
C891 B.n114 VSUBS 0.007329f
C892 B.n115 VSUBS 0.007329f
C893 B.n116 VSUBS 0.007329f
C894 B.n117 VSUBS 0.007329f
C895 B.n118 VSUBS 0.007329f
C896 B.n119 VSUBS 0.007329f
C897 B.n120 VSUBS 0.007329f
C898 B.n121 VSUBS 0.007329f
C899 B.n122 VSUBS 0.007329f
C900 B.n123 VSUBS 0.007329f
C901 B.n124 VSUBS 0.007329f
C902 B.n125 VSUBS 0.007329f
C903 B.n126 VSUBS 0.007329f
C904 B.n127 VSUBS 0.007329f
C905 B.n128 VSUBS 0.007329f
C906 B.n129 VSUBS 0.007329f
C907 B.n130 VSUBS 0.007329f
C908 B.n131 VSUBS 0.007329f
C909 B.n132 VSUBS 0.007329f
C910 B.n133 VSUBS 0.007329f
C911 B.n134 VSUBS 0.007329f
C912 B.n135 VSUBS 0.007329f
C913 B.n136 VSUBS 0.007329f
C914 B.n137 VSUBS 0.007329f
C915 B.n138 VSUBS 0.007329f
C916 B.n139 VSUBS 0.007329f
C917 B.n140 VSUBS 0.007329f
C918 B.n141 VSUBS 0.007329f
C919 B.n142 VSUBS 0.007329f
C920 B.n143 VSUBS 0.007329f
C921 B.n144 VSUBS 0.016256f
C922 B.n145 VSUBS 0.007329f
C923 B.n146 VSUBS 0.007329f
C924 B.n147 VSUBS 0.007329f
C925 B.n148 VSUBS 0.007329f
C926 B.n149 VSUBS 0.007329f
C927 B.n150 VSUBS 0.007329f
C928 B.n151 VSUBS 0.007329f
C929 B.n152 VSUBS 0.007329f
C930 B.n153 VSUBS 0.007329f
C931 B.n154 VSUBS 0.007329f
C932 B.n155 VSUBS 0.007329f
C933 B.n156 VSUBS 0.007329f
C934 B.n157 VSUBS 0.007329f
C935 B.n158 VSUBS 0.007329f
C936 B.n159 VSUBS 0.007329f
C937 B.n160 VSUBS 0.007329f
C938 B.n161 VSUBS 0.007329f
C939 B.n162 VSUBS 0.007329f
C940 B.n163 VSUBS 0.007329f
C941 B.n164 VSUBS 0.007329f
C942 B.n165 VSUBS 0.007329f
C943 B.t2 VSUBS 0.224332f
C944 B.t1 VSUBS 0.264037f
C945 B.t0 VSUBS 1.88903f
C946 B.n166 VSUBS 0.42094f
C947 B.n167 VSUBS 0.268293f
C948 B.n168 VSUBS 0.007329f
C949 B.n169 VSUBS 0.007329f
C950 B.n170 VSUBS 0.007329f
C951 B.n171 VSUBS 0.007329f
C952 B.n172 VSUBS 0.004096f
C953 B.n173 VSUBS 0.007329f
C954 B.n174 VSUBS 0.007329f
C955 B.n175 VSUBS 0.007329f
C956 B.n176 VSUBS 0.007329f
C957 B.n177 VSUBS 0.007329f
C958 B.n178 VSUBS 0.007329f
C959 B.n179 VSUBS 0.007329f
C960 B.n180 VSUBS 0.007329f
C961 B.n181 VSUBS 0.007329f
C962 B.n182 VSUBS 0.007329f
C963 B.n183 VSUBS 0.007329f
C964 B.n184 VSUBS 0.007329f
C965 B.n185 VSUBS 0.007329f
C966 B.n186 VSUBS 0.007329f
C967 B.n187 VSUBS 0.007329f
C968 B.n188 VSUBS 0.007329f
C969 B.n189 VSUBS 0.007329f
C970 B.n190 VSUBS 0.007329f
C971 B.n191 VSUBS 0.007329f
C972 B.n192 VSUBS 0.007329f
C973 B.n193 VSUBS 0.016207f
C974 B.n194 VSUBS 0.007329f
C975 B.n195 VSUBS 0.007329f
C976 B.n196 VSUBS 0.007329f
C977 B.n197 VSUBS 0.007329f
C978 B.n198 VSUBS 0.007329f
C979 B.n199 VSUBS 0.007329f
C980 B.n200 VSUBS 0.007329f
C981 B.n201 VSUBS 0.007329f
C982 B.n202 VSUBS 0.007329f
C983 B.n203 VSUBS 0.007329f
C984 B.n204 VSUBS 0.007329f
C985 B.n205 VSUBS 0.007329f
C986 B.n206 VSUBS 0.007329f
C987 B.n207 VSUBS 0.007329f
C988 B.n208 VSUBS 0.007329f
C989 B.n209 VSUBS 0.007329f
C990 B.n210 VSUBS 0.007329f
C991 B.n211 VSUBS 0.007329f
C992 B.n212 VSUBS 0.007329f
C993 B.n213 VSUBS 0.007329f
C994 B.n214 VSUBS 0.007329f
C995 B.n215 VSUBS 0.007329f
C996 B.n216 VSUBS 0.007329f
C997 B.n217 VSUBS 0.007329f
C998 B.n218 VSUBS 0.007329f
C999 B.n219 VSUBS 0.007329f
C1000 B.n220 VSUBS 0.007329f
C1001 B.n221 VSUBS 0.007329f
C1002 B.n222 VSUBS 0.007329f
C1003 B.n223 VSUBS 0.007329f
C1004 B.n224 VSUBS 0.007329f
C1005 B.n225 VSUBS 0.007329f
C1006 B.n226 VSUBS 0.007329f
C1007 B.n227 VSUBS 0.007329f
C1008 B.n228 VSUBS 0.007329f
C1009 B.n229 VSUBS 0.007329f
C1010 B.n230 VSUBS 0.007329f
C1011 B.n231 VSUBS 0.007329f
C1012 B.n232 VSUBS 0.007329f
C1013 B.n233 VSUBS 0.007329f
C1014 B.n234 VSUBS 0.007329f
C1015 B.n235 VSUBS 0.007329f
C1016 B.n236 VSUBS 0.007329f
C1017 B.n237 VSUBS 0.007329f
C1018 B.n238 VSUBS 0.007329f
C1019 B.n239 VSUBS 0.007329f
C1020 B.n240 VSUBS 0.007329f
C1021 B.n241 VSUBS 0.007329f
C1022 B.n242 VSUBS 0.007329f
C1023 B.n243 VSUBS 0.007329f
C1024 B.n244 VSUBS 0.007329f
C1025 B.n245 VSUBS 0.007329f
C1026 B.n246 VSUBS 0.007329f
C1027 B.n247 VSUBS 0.007329f
C1028 B.n248 VSUBS 0.007329f
C1029 B.n249 VSUBS 0.007329f
C1030 B.n250 VSUBS 0.007329f
C1031 B.n251 VSUBS 0.007329f
C1032 B.n252 VSUBS 0.007329f
C1033 B.n253 VSUBS 0.007329f
C1034 B.n254 VSUBS 0.007329f
C1035 B.n255 VSUBS 0.007329f
C1036 B.n256 VSUBS 0.007329f
C1037 B.n257 VSUBS 0.007329f
C1038 B.n258 VSUBS 0.007329f
C1039 B.n259 VSUBS 0.007329f
C1040 B.n260 VSUBS 0.007329f
C1041 B.n261 VSUBS 0.007329f
C1042 B.n262 VSUBS 0.007329f
C1043 B.n263 VSUBS 0.007329f
C1044 B.n264 VSUBS 0.007329f
C1045 B.n265 VSUBS 0.007329f
C1046 B.n266 VSUBS 0.007329f
C1047 B.n267 VSUBS 0.007329f
C1048 B.n268 VSUBS 0.007329f
C1049 B.n269 VSUBS 0.007329f
C1050 B.n270 VSUBS 0.007329f
C1051 B.n271 VSUBS 0.007329f
C1052 B.n272 VSUBS 0.007329f
C1053 B.n273 VSUBS 0.007329f
C1054 B.n274 VSUBS 0.007329f
C1055 B.n275 VSUBS 0.007329f
C1056 B.n276 VSUBS 0.007329f
C1057 B.n277 VSUBS 0.007329f
C1058 B.n278 VSUBS 0.007329f
C1059 B.n279 VSUBS 0.007329f
C1060 B.n280 VSUBS 0.007329f
C1061 B.n281 VSUBS 0.007329f
C1062 B.n282 VSUBS 0.007329f
C1063 B.n283 VSUBS 0.007329f
C1064 B.n284 VSUBS 0.007329f
C1065 B.n285 VSUBS 0.007329f
C1066 B.n286 VSUBS 0.007329f
C1067 B.n287 VSUBS 0.007329f
C1068 B.n288 VSUBS 0.007329f
C1069 B.n289 VSUBS 0.007329f
C1070 B.n290 VSUBS 0.007329f
C1071 B.n291 VSUBS 0.007329f
C1072 B.n292 VSUBS 0.007329f
C1073 B.n293 VSUBS 0.007329f
C1074 B.n294 VSUBS 0.007329f
C1075 B.n295 VSUBS 0.007329f
C1076 B.n296 VSUBS 0.007329f
C1077 B.n297 VSUBS 0.007329f
C1078 B.n298 VSUBS 0.007329f
C1079 B.n299 VSUBS 0.007329f
C1080 B.n300 VSUBS 0.007329f
C1081 B.n301 VSUBS 0.007329f
C1082 B.n302 VSUBS 0.007329f
C1083 B.n303 VSUBS 0.007329f
C1084 B.n304 VSUBS 0.007329f
C1085 B.n305 VSUBS 0.007329f
C1086 B.n306 VSUBS 0.007329f
C1087 B.n307 VSUBS 0.007329f
C1088 B.n308 VSUBS 0.007329f
C1089 B.n309 VSUBS 0.007329f
C1090 B.n310 VSUBS 0.015266f
C1091 B.n311 VSUBS 0.015266f
C1092 B.n312 VSUBS 0.016207f
C1093 B.n313 VSUBS 0.007329f
C1094 B.n314 VSUBS 0.007329f
C1095 B.n315 VSUBS 0.007329f
C1096 B.n316 VSUBS 0.007329f
C1097 B.n317 VSUBS 0.007329f
C1098 B.n318 VSUBS 0.007329f
C1099 B.n319 VSUBS 0.007329f
C1100 B.n320 VSUBS 0.007329f
C1101 B.n321 VSUBS 0.007329f
C1102 B.n322 VSUBS 0.007329f
C1103 B.n323 VSUBS 0.007329f
C1104 B.n324 VSUBS 0.007329f
C1105 B.n325 VSUBS 0.007329f
C1106 B.n326 VSUBS 0.007329f
C1107 B.n327 VSUBS 0.007329f
C1108 B.n328 VSUBS 0.007329f
C1109 B.n329 VSUBS 0.007329f
C1110 B.n330 VSUBS 0.007329f
C1111 B.n331 VSUBS 0.007329f
C1112 B.n332 VSUBS 0.007329f
C1113 B.n333 VSUBS 0.007329f
C1114 B.n334 VSUBS 0.007329f
C1115 B.n335 VSUBS 0.007329f
C1116 B.n336 VSUBS 0.007329f
C1117 B.n337 VSUBS 0.007329f
C1118 B.n338 VSUBS 0.007329f
C1119 B.n339 VSUBS 0.007329f
C1120 B.n340 VSUBS 0.007329f
C1121 B.n341 VSUBS 0.007329f
C1122 B.n342 VSUBS 0.007329f
C1123 B.n343 VSUBS 0.007329f
C1124 B.n344 VSUBS 0.007329f
C1125 B.n345 VSUBS 0.007329f
C1126 B.n346 VSUBS 0.007329f
C1127 B.n347 VSUBS 0.007329f
C1128 B.n348 VSUBS 0.007329f
C1129 B.n349 VSUBS 0.007329f
C1130 B.n350 VSUBS 0.007329f
C1131 B.n351 VSUBS 0.007329f
C1132 B.n352 VSUBS 0.007329f
C1133 B.n353 VSUBS 0.007329f
C1134 B.n354 VSUBS 0.007329f
C1135 B.n355 VSUBS 0.007329f
C1136 B.n356 VSUBS 0.007329f
C1137 B.n357 VSUBS 0.007329f
C1138 B.n358 VSUBS 0.007329f
C1139 B.n359 VSUBS 0.007329f
C1140 B.n360 VSUBS 0.007329f
C1141 B.n361 VSUBS 0.007329f
C1142 B.n362 VSUBS 0.007329f
C1143 B.n363 VSUBS 0.007329f
C1144 B.n364 VSUBS 0.007329f
C1145 B.n365 VSUBS 0.007329f
C1146 B.n366 VSUBS 0.007329f
C1147 B.n367 VSUBS 0.007329f
C1148 B.n368 VSUBS 0.007329f
C1149 B.n369 VSUBS 0.007329f
C1150 B.n370 VSUBS 0.007329f
C1151 B.n371 VSUBS 0.007329f
C1152 B.n372 VSUBS 0.007329f
C1153 B.t11 VSUBS 0.224329f
C1154 B.t10 VSUBS 0.264035f
C1155 B.t9 VSUBS 1.88903f
C1156 B.n373 VSUBS 0.420943f
C1157 B.n374 VSUBS 0.268296f
C1158 B.n375 VSUBS 0.016981f
C1159 B.n376 VSUBS 0.006898f
C1160 B.n377 VSUBS 0.007329f
C1161 B.n378 VSUBS 0.007329f
C1162 B.n379 VSUBS 0.007329f
C1163 B.n380 VSUBS 0.007329f
C1164 B.n381 VSUBS 0.007329f
C1165 B.n382 VSUBS 0.007329f
C1166 B.n383 VSUBS 0.007329f
C1167 B.n384 VSUBS 0.007329f
C1168 B.n385 VSUBS 0.007329f
C1169 B.n386 VSUBS 0.007329f
C1170 B.n387 VSUBS 0.007329f
C1171 B.n388 VSUBS 0.007329f
C1172 B.n389 VSUBS 0.007329f
C1173 B.n390 VSUBS 0.007329f
C1174 B.n391 VSUBS 0.007329f
C1175 B.n392 VSUBS 0.004096f
C1176 B.n393 VSUBS 0.016981f
C1177 B.n394 VSUBS 0.006898f
C1178 B.n395 VSUBS 0.007329f
C1179 B.n396 VSUBS 0.007329f
C1180 B.n397 VSUBS 0.007329f
C1181 B.n398 VSUBS 0.007329f
C1182 B.n399 VSUBS 0.007329f
C1183 B.n400 VSUBS 0.007329f
C1184 B.n401 VSUBS 0.007329f
C1185 B.n402 VSUBS 0.007329f
C1186 B.n403 VSUBS 0.007329f
C1187 B.n404 VSUBS 0.007329f
C1188 B.n405 VSUBS 0.007329f
C1189 B.n406 VSUBS 0.007329f
C1190 B.n407 VSUBS 0.007329f
C1191 B.n408 VSUBS 0.007329f
C1192 B.n409 VSUBS 0.007329f
C1193 B.n410 VSUBS 0.007329f
C1194 B.n411 VSUBS 0.007329f
C1195 B.n412 VSUBS 0.007329f
C1196 B.n413 VSUBS 0.007329f
C1197 B.n414 VSUBS 0.007329f
C1198 B.n415 VSUBS 0.007329f
C1199 B.n416 VSUBS 0.007329f
C1200 B.n417 VSUBS 0.007329f
C1201 B.n418 VSUBS 0.007329f
C1202 B.n419 VSUBS 0.007329f
C1203 B.n420 VSUBS 0.007329f
C1204 B.n421 VSUBS 0.007329f
C1205 B.n422 VSUBS 0.007329f
C1206 B.n423 VSUBS 0.007329f
C1207 B.n424 VSUBS 0.007329f
C1208 B.n425 VSUBS 0.007329f
C1209 B.n426 VSUBS 0.007329f
C1210 B.n427 VSUBS 0.007329f
C1211 B.n428 VSUBS 0.007329f
C1212 B.n429 VSUBS 0.007329f
C1213 B.n430 VSUBS 0.007329f
C1214 B.n431 VSUBS 0.007329f
C1215 B.n432 VSUBS 0.007329f
C1216 B.n433 VSUBS 0.007329f
C1217 B.n434 VSUBS 0.007329f
C1218 B.n435 VSUBS 0.007329f
C1219 B.n436 VSUBS 0.007329f
C1220 B.n437 VSUBS 0.007329f
C1221 B.n438 VSUBS 0.007329f
C1222 B.n439 VSUBS 0.007329f
C1223 B.n440 VSUBS 0.007329f
C1224 B.n441 VSUBS 0.007329f
C1225 B.n442 VSUBS 0.007329f
C1226 B.n443 VSUBS 0.007329f
C1227 B.n444 VSUBS 0.007329f
C1228 B.n445 VSUBS 0.007329f
C1229 B.n446 VSUBS 0.007329f
C1230 B.n447 VSUBS 0.007329f
C1231 B.n448 VSUBS 0.007329f
C1232 B.n449 VSUBS 0.007329f
C1233 B.n450 VSUBS 0.007329f
C1234 B.n451 VSUBS 0.007329f
C1235 B.n452 VSUBS 0.007329f
C1236 B.n453 VSUBS 0.007329f
C1237 B.n454 VSUBS 0.007329f
C1238 B.n455 VSUBS 0.015217f
C1239 B.n456 VSUBS 0.016207f
C1240 B.n457 VSUBS 0.015266f
C1241 B.n458 VSUBS 0.007329f
C1242 B.n459 VSUBS 0.007329f
C1243 B.n460 VSUBS 0.007329f
C1244 B.n461 VSUBS 0.007329f
C1245 B.n462 VSUBS 0.007329f
C1246 B.n463 VSUBS 0.007329f
C1247 B.n464 VSUBS 0.007329f
C1248 B.n465 VSUBS 0.007329f
C1249 B.n466 VSUBS 0.007329f
C1250 B.n467 VSUBS 0.007329f
C1251 B.n468 VSUBS 0.007329f
C1252 B.n469 VSUBS 0.007329f
C1253 B.n470 VSUBS 0.007329f
C1254 B.n471 VSUBS 0.007329f
C1255 B.n472 VSUBS 0.007329f
C1256 B.n473 VSUBS 0.007329f
C1257 B.n474 VSUBS 0.007329f
C1258 B.n475 VSUBS 0.007329f
C1259 B.n476 VSUBS 0.007329f
C1260 B.n477 VSUBS 0.007329f
C1261 B.n478 VSUBS 0.007329f
C1262 B.n479 VSUBS 0.007329f
C1263 B.n480 VSUBS 0.007329f
C1264 B.n481 VSUBS 0.007329f
C1265 B.n482 VSUBS 0.007329f
C1266 B.n483 VSUBS 0.007329f
C1267 B.n484 VSUBS 0.007329f
C1268 B.n485 VSUBS 0.007329f
C1269 B.n486 VSUBS 0.007329f
C1270 B.n487 VSUBS 0.007329f
C1271 B.n488 VSUBS 0.007329f
C1272 B.n489 VSUBS 0.007329f
C1273 B.n490 VSUBS 0.007329f
C1274 B.n491 VSUBS 0.007329f
C1275 B.n492 VSUBS 0.007329f
C1276 B.n493 VSUBS 0.007329f
C1277 B.n494 VSUBS 0.007329f
C1278 B.n495 VSUBS 0.007329f
C1279 B.n496 VSUBS 0.007329f
C1280 B.n497 VSUBS 0.007329f
C1281 B.n498 VSUBS 0.007329f
C1282 B.n499 VSUBS 0.007329f
C1283 B.n500 VSUBS 0.007329f
C1284 B.n501 VSUBS 0.007329f
C1285 B.n502 VSUBS 0.007329f
C1286 B.n503 VSUBS 0.007329f
C1287 B.n504 VSUBS 0.007329f
C1288 B.n505 VSUBS 0.007329f
C1289 B.n506 VSUBS 0.007329f
C1290 B.n507 VSUBS 0.007329f
C1291 B.n508 VSUBS 0.007329f
C1292 B.n509 VSUBS 0.007329f
C1293 B.n510 VSUBS 0.007329f
C1294 B.n511 VSUBS 0.007329f
C1295 B.n512 VSUBS 0.007329f
C1296 B.n513 VSUBS 0.007329f
C1297 B.n514 VSUBS 0.007329f
C1298 B.n515 VSUBS 0.007329f
C1299 B.n516 VSUBS 0.007329f
C1300 B.n517 VSUBS 0.007329f
C1301 B.n518 VSUBS 0.007329f
C1302 B.n519 VSUBS 0.007329f
C1303 B.n520 VSUBS 0.007329f
C1304 B.n521 VSUBS 0.007329f
C1305 B.n522 VSUBS 0.007329f
C1306 B.n523 VSUBS 0.007329f
C1307 B.n524 VSUBS 0.007329f
C1308 B.n525 VSUBS 0.007329f
C1309 B.n526 VSUBS 0.007329f
C1310 B.n527 VSUBS 0.007329f
C1311 B.n528 VSUBS 0.007329f
C1312 B.n529 VSUBS 0.007329f
C1313 B.n530 VSUBS 0.007329f
C1314 B.n531 VSUBS 0.007329f
C1315 B.n532 VSUBS 0.007329f
C1316 B.n533 VSUBS 0.007329f
C1317 B.n534 VSUBS 0.007329f
C1318 B.n535 VSUBS 0.007329f
C1319 B.n536 VSUBS 0.007329f
C1320 B.n537 VSUBS 0.007329f
C1321 B.n538 VSUBS 0.007329f
C1322 B.n539 VSUBS 0.007329f
C1323 B.n540 VSUBS 0.007329f
C1324 B.n541 VSUBS 0.007329f
C1325 B.n542 VSUBS 0.007329f
C1326 B.n543 VSUBS 0.007329f
C1327 B.n544 VSUBS 0.007329f
C1328 B.n545 VSUBS 0.007329f
C1329 B.n546 VSUBS 0.007329f
C1330 B.n547 VSUBS 0.007329f
C1331 B.n548 VSUBS 0.007329f
C1332 B.n549 VSUBS 0.007329f
C1333 B.n550 VSUBS 0.007329f
C1334 B.n551 VSUBS 0.007329f
C1335 B.n552 VSUBS 0.007329f
C1336 B.n553 VSUBS 0.007329f
C1337 B.n554 VSUBS 0.007329f
C1338 B.n555 VSUBS 0.007329f
C1339 B.n556 VSUBS 0.007329f
C1340 B.n557 VSUBS 0.007329f
C1341 B.n558 VSUBS 0.007329f
C1342 B.n559 VSUBS 0.007329f
C1343 B.n560 VSUBS 0.007329f
C1344 B.n561 VSUBS 0.007329f
C1345 B.n562 VSUBS 0.007329f
C1346 B.n563 VSUBS 0.007329f
C1347 B.n564 VSUBS 0.007329f
C1348 B.n565 VSUBS 0.007329f
C1349 B.n566 VSUBS 0.007329f
C1350 B.n567 VSUBS 0.007329f
C1351 B.n568 VSUBS 0.007329f
C1352 B.n569 VSUBS 0.007329f
C1353 B.n570 VSUBS 0.007329f
C1354 B.n571 VSUBS 0.007329f
C1355 B.n572 VSUBS 0.007329f
C1356 B.n573 VSUBS 0.007329f
C1357 B.n574 VSUBS 0.007329f
C1358 B.n575 VSUBS 0.007329f
C1359 B.n576 VSUBS 0.007329f
C1360 B.n577 VSUBS 0.007329f
C1361 B.n578 VSUBS 0.007329f
C1362 B.n579 VSUBS 0.007329f
C1363 B.n580 VSUBS 0.007329f
C1364 B.n581 VSUBS 0.007329f
C1365 B.n582 VSUBS 0.007329f
C1366 B.n583 VSUBS 0.007329f
C1367 B.n584 VSUBS 0.007329f
C1368 B.n585 VSUBS 0.007329f
C1369 B.n586 VSUBS 0.007329f
C1370 B.n587 VSUBS 0.007329f
C1371 B.n588 VSUBS 0.007329f
C1372 B.n589 VSUBS 0.007329f
C1373 B.n590 VSUBS 0.007329f
C1374 B.n591 VSUBS 0.007329f
C1375 B.n592 VSUBS 0.007329f
C1376 B.n593 VSUBS 0.007329f
C1377 B.n594 VSUBS 0.007329f
C1378 B.n595 VSUBS 0.007329f
C1379 B.n596 VSUBS 0.007329f
C1380 B.n597 VSUBS 0.007329f
C1381 B.n598 VSUBS 0.007329f
C1382 B.n599 VSUBS 0.007329f
C1383 B.n600 VSUBS 0.007329f
C1384 B.n601 VSUBS 0.007329f
C1385 B.n602 VSUBS 0.007329f
C1386 B.n603 VSUBS 0.007329f
C1387 B.n604 VSUBS 0.007329f
C1388 B.n605 VSUBS 0.007329f
C1389 B.n606 VSUBS 0.007329f
C1390 B.n607 VSUBS 0.007329f
C1391 B.n608 VSUBS 0.007329f
C1392 B.n609 VSUBS 0.007329f
C1393 B.n610 VSUBS 0.007329f
C1394 B.n611 VSUBS 0.007329f
C1395 B.n612 VSUBS 0.007329f
C1396 B.n613 VSUBS 0.007329f
C1397 B.n614 VSUBS 0.007329f
C1398 B.n615 VSUBS 0.007329f
C1399 B.n616 VSUBS 0.007329f
C1400 B.n617 VSUBS 0.007329f
C1401 B.n618 VSUBS 0.007329f
C1402 B.n619 VSUBS 0.007329f
C1403 B.n620 VSUBS 0.007329f
C1404 B.n621 VSUBS 0.007329f
C1405 B.n622 VSUBS 0.007329f
C1406 B.n623 VSUBS 0.007329f
C1407 B.n624 VSUBS 0.007329f
C1408 B.n625 VSUBS 0.007329f
C1409 B.n626 VSUBS 0.007329f
C1410 B.n627 VSUBS 0.007329f
C1411 B.n628 VSUBS 0.007329f
C1412 B.n629 VSUBS 0.007329f
C1413 B.n630 VSUBS 0.007329f
C1414 B.n631 VSUBS 0.007329f
C1415 B.n632 VSUBS 0.007329f
C1416 B.n633 VSUBS 0.007329f
C1417 B.n634 VSUBS 0.007329f
C1418 B.n635 VSUBS 0.007329f
C1419 B.n636 VSUBS 0.007329f
C1420 B.n637 VSUBS 0.007329f
C1421 B.n638 VSUBS 0.015266f
C1422 B.n639 VSUBS 0.015266f
C1423 B.n640 VSUBS 0.016207f
C1424 B.n641 VSUBS 0.007329f
C1425 B.n642 VSUBS 0.007329f
C1426 B.n643 VSUBS 0.007329f
C1427 B.n644 VSUBS 0.007329f
C1428 B.n645 VSUBS 0.007329f
C1429 B.n646 VSUBS 0.007329f
C1430 B.n647 VSUBS 0.007329f
C1431 B.n648 VSUBS 0.007329f
C1432 B.n649 VSUBS 0.007329f
C1433 B.n650 VSUBS 0.007329f
C1434 B.n651 VSUBS 0.007329f
C1435 B.n652 VSUBS 0.007329f
C1436 B.n653 VSUBS 0.007329f
C1437 B.n654 VSUBS 0.007329f
C1438 B.n655 VSUBS 0.007329f
C1439 B.n656 VSUBS 0.007329f
C1440 B.n657 VSUBS 0.007329f
C1441 B.n658 VSUBS 0.007329f
C1442 B.n659 VSUBS 0.007329f
C1443 B.n660 VSUBS 0.007329f
C1444 B.n661 VSUBS 0.007329f
C1445 B.n662 VSUBS 0.007329f
C1446 B.n663 VSUBS 0.007329f
C1447 B.n664 VSUBS 0.007329f
C1448 B.n665 VSUBS 0.007329f
C1449 B.n666 VSUBS 0.007329f
C1450 B.n667 VSUBS 0.007329f
C1451 B.n668 VSUBS 0.007329f
C1452 B.n669 VSUBS 0.007329f
C1453 B.n670 VSUBS 0.007329f
C1454 B.n671 VSUBS 0.007329f
C1455 B.n672 VSUBS 0.007329f
C1456 B.n673 VSUBS 0.007329f
C1457 B.n674 VSUBS 0.007329f
C1458 B.n675 VSUBS 0.007329f
C1459 B.n676 VSUBS 0.007329f
C1460 B.n677 VSUBS 0.007329f
C1461 B.n678 VSUBS 0.007329f
C1462 B.n679 VSUBS 0.007329f
C1463 B.n680 VSUBS 0.007329f
C1464 B.n681 VSUBS 0.007329f
C1465 B.n682 VSUBS 0.007329f
C1466 B.n683 VSUBS 0.007329f
C1467 B.n684 VSUBS 0.007329f
C1468 B.n685 VSUBS 0.007329f
C1469 B.n686 VSUBS 0.007329f
C1470 B.n687 VSUBS 0.007329f
C1471 B.n688 VSUBS 0.007329f
C1472 B.n689 VSUBS 0.007329f
C1473 B.n690 VSUBS 0.007329f
C1474 B.n691 VSUBS 0.007329f
C1475 B.n692 VSUBS 0.007329f
C1476 B.n693 VSUBS 0.007329f
C1477 B.n694 VSUBS 0.007329f
C1478 B.n695 VSUBS 0.007329f
C1479 B.n696 VSUBS 0.007329f
C1480 B.n697 VSUBS 0.007329f
C1481 B.n698 VSUBS 0.007329f
C1482 B.n699 VSUBS 0.007329f
C1483 B.n700 VSUBS 0.007329f
C1484 B.n701 VSUBS 0.006898f
C1485 B.n702 VSUBS 0.007329f
C1486 B.n703 VSUBS 0.007329f
C1487 B.n704 VSUBS 0.004096f
C1488 B.n705 VSUBS 0.007329f
C1489 B.n706 VSUBS 0.007329f
C1490 B.n707 VSUBS 0.007329f
C1491 B.n708 VSUBS 0.007329f
C1492 B.n709 VSUBS 0.007329f
C1493 B.n710 VSUBS 0.007329f
C1494 B.n711 VSUBS 0.007329f
C1495 B.n712 VSUBS 0.007329f
C1496 B.n713 VSUBS 0.007329f
C1497 B.n714 VSUBS 0.007329f
C1498 B.n715 VSUBS 0.007329f
C1499 B.n716 VSUBS 0.007329f
C1500 B.n717 VSUBS 0.004096f
C1501 B.n718 VSUBS 0.016981f
C1502 B.n719 VSUBS 0.006898f
C1503 B.n720 VSUBS 0.007329f
C1504 B.n721 VSUBS 0.007329f
C1505 B.n722 VSUBS 0.007329f
C1506 B.n723 VSUBS 0.007329f
C1507 B.n724 VSUBS 0.007329f
C1508 B.n725 VSUBS 0.007329f
C1509 B.n726 VSUBS 0.007329f
C1510 B.n727 VSUBS 0.007329f
C1511 B.n728 VSUBS 0.007329f
C1512 B.n729 VSUBS 0.007329f
C1513 B.n730 VSUBS 0.007329f
C1514 B.n731 VSUBS 0.007329f
C1515 B.n732 VSUBS 0.007329f
C1516 B.n733 VSUBS 0.007329f
C1517 B.n734 VSUBS 0.007329f
C1518 B.n735 VSUBS 0.007329f
C1519 B.n736 VSUBS 0.007329f
C1520 B.n737 VSUBS 0.007329f
C1521 B.n738 VSUBS 0.007329f
C1522 B.n739 VSUBS 0.007329f
C1523 B.n740 VSUBS 0.007329f
C1524 B.n741 VSUBS 0.007329f
C1525 B.n742 VSUBS 0.007329f
C1526 B.n743 VSUBS 0.007329f
C1527 B.n744 VSUBS 0.007329f
C1528 B.n745 VSUBS 0.007329f
C1529 B.n746 VSUBS 0.007329f
C1530 B.n747 VSUBS 0.007329f
C1531 B.n748 VSUBS 0.007329f
C1532 B.n749 VSUBS 0.007329f
C1533 B.n750 VSUBS 0.007329f
C1534 B.n751 VSUBS 0.007329f
C1535 B.n752 VSUBS 0.007329f
C1536 B.n753 VSUBS 0.007329f
C1537 B.n754 VSUBS 0.007329f
C1538 B.n755 VSUBS 0.007329f
C1539 B.n756 VSUBS 0.007329f
C1540 B.n757 VSUBS 0.007329f
C1541 B.n758 VSUBS 0.007329f
C1542 B.n759 VSUBS 0.007329f
C1543 B.n760 VSUBS 0.007329f
C1544 B.n761 VSUBS 0.007329f
C1545 B.n762 VSUBS 0.007329f
C1546 B.n763 VSUBS 0.007329f
C1547 B.n764 VSUBS 0.007329f
C1548 B.n765 VSUBS 0.007329f
C1549 B.n766 VSUBS 0.007329f
C1550 B.n767 VSUBS 0.007329f
C1551 B.n768 VSUBS 0.007329f
C1552 B.n769 VSUBS 0.007329f
C1553 B.n770 VSUBS 0.007329f
C1554 B.n771 VSUBS 0.007329f
C1555 B.n772 VSUBS 0.007329f
C1556 B.n773 VSUBS 0.007329f
C1557 B.n774 VSUBS 0.007329f
C1558 B.n775 VSUBS 0.007329f
C1559 B.n776 VSUBS 0.007329f
C1560 B.n777 VSUBS 0.007329f
C1561 B.n778 VSUBS 0.007329f
C1562 B.n779 VSUBS 0.007329f
C1563 B.n780 VSUBS 0.007329f
C1564 B.n781 VSUBS 0.016207f
C1565 B.n782 VSUBS 0.015266f
C1566 B.n783 VSUBS 0.015266f
C1567 B.n784 VSUBS 0.007329f
C1568 B.n785 VSUBS 0.007329f
C1569 B.n786 VSUBS 0.007329f
C1570 B.n787 VSUBS 0.007329f
C1571 B.n788 VSUBS 0.007329f
C1572 B.n789 VSUBS 0.007329f
C1573 B.n790 VSUBS 0.007329f
C1574 B.n791 VSUBS 0.007329f
C1575 B.n792 VSUBS 0.007329f
C1576 B.n793 VSUBS 0.007329f
C1577 B.n794 VSUBS 0.007329f
C1578 B.n795 VSUBS 0.007329f
C1579 B.n796 VSUBS 0.007329f
C1580 B.n797 VSUBS 0.007329f
C1581 B.n798 VSUBS 0.007329f
C1582 B.n799 VSUBS 0.007329f
C1583 B.n800 VSUBS 0.007329f
C1584 B.n801 VSUBS 0.007329f
C1585 B.n802 VSUBS 0.007329f
C1586 B.n803 VSUBS 0.007329f
C1587 B.n804 VSUBS 0.007329f
C1588 B.n805 VSUBS 0.007329f
C1589 B.n806 VSUBS 0.007329f
C1590 B.n807 VSUBS 0.007329f
C1591 B.n808 VSUBS 0.007329f
C1592 B.n809 VSUBS 0.007329f
C1593 B.n810 VSUBS 0.007329f
C1594 B.n811 VSUBS 0.007329f
C1595 B.n812 VSUBS 0.007329f
C1596 B.n813 VSUBS 0.007329f
C1597 B.n814 VSUBS 0.007329f
C1598 B.n815 VSUBS 0.007329f
C1599 B.n816 VSUBS 0.007329f
C1600 B.n817 VSUBS 0.007329f
C1601 B.n818 VSUBS 0.007329f
C1602 B.n819 VSUBS 0.007329f
C1603 B.n820 VSUBS 0.007329f
C1604 B.n821 VSUBS 0.007329f
C1605 B.n822 VSUBS 0.007329f
C1606 B.n823 VSUBS 0.007329f
C1607 B.n824 VSUBS 0.007329f
C1608 B.n825 VSUBS 0.007329f
C1609 B.n826 VSUBS 0.007329f
C1610 B.n827 VSUBS 0.007329f
C1611 B.n828 VSUBS 0.007329f
C1612 B.n829 VSUBS 0.007329f
C1613 B.n830 VSUBS 0.007329f
C1614 B.n831 VSUBS 0.007329f
C1615 B.n832 VSUBS 0.007329f
C1616 B.n833 VSUBS 0.007329f
C1617 B.n834 VSUBS 0.007329f
C1618 B.n835 VSUBS 0.007329f
C1619 B.n836 VSUBS 0.007329f
C1620 B.n837 VSUBS 0.007329f
C1621 B.n838 VSUBS 0.007329f
C1622 B.n839 VSUBS 0.007329f
C1623 B.n840 VSUBS 0.007329f
C1624 B.n841 VSUBS 0.007329f
C1625 B.n842 VSUBS 0.007329f
C1626 B.n843 VSUBS 0.007329f
C1627 B.n844 VSUBS 0.007329f
C1628 B.n845 VSUBS 0.007329f
C1629 B.n846 VSUBS 0.007329f
C1630 B.n847 VSUBS 0.007329f
C1631 B.n848 VSUBS 0.007329f
C1632 B.n849 VSUBS 0.007329f
C1633 B.n850 VSUBS 0.007329f
C1634 B.n851 VSUBS 0.007329f
C1635 B.n852 VSUBS 0.007329f
C1636 B.n853 VSUBS 0.007329f
C1637 B.n854 VSUBS 0.007329f
C1638 B.n855 VSUBS 0.007329f
C1639 B.n856 VSUBS 0.007329f
C1640 B.n857 VSUBS 0.007329f
C1641 B.n858 VSUBS 0.007329f
C1642 B.n859 VSUBS 0.007329f
C1643 B.n860 VSUBS 0.007329f
C1644 B.n861 VSUBS 0.007329f
C1645 B.n862 VSUBS 0.007329f
C1646 B.n863 VSUBS 0.007329f
C1647 B.n864 VSUBS 0.007329f
C1648 B.n865 VSUBS 0.007329f
C1649 B.n866 VSUBS 0.007329f
C1650 B.n867 VSUBS 0.007329f
C1651 B.n868 VSUBS 0.007329f
C1652 B.n869 VSUBS 0.007329f
C1653 B.n870 VSUBS 0.007329f
C1654 B.n871 VSUBS 0.009564f
C1655 B.n872 VSUBS 0.010189f
C1656 B.n873 VSUBS 0.020261f
.ends

