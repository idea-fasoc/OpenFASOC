* NGSPICE file created from diff_pair_sample_0745.ext - technology: sky130A

.subckt diff_pair_sample_0745 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n1294_n2542# sky130_fd_pr__pfet_01v8 ad=3.0615 pd=16.48 as=0 ps=0 w=7.85 l=0.21
X1 VTAIL.t7 VP.t0 VDD1.t2 w_n1294_n2542# sky130_fd_pr__pfet_01v8 ad=3.0615 pd=16.48 as=1.29525 ps=8.18 w=7.85 l=0.21
X2 VDD1.t0 VP.t1 VTAIL.t6 w_n1294_n2542# sky130_fd_pr__pfet_01v8 ad=1.29525 pd=8.18 as=3.0615 ps=16.48 w=7.85 l=0.21
X3 VTAIL.t0 VN.t0 VDD2.t3 w_n1294_n2542# sky130_fd_pr__pfet_01v8 ad=3.0615 pd=16.48 as=1.29525 ps=8.18 w=7.85 l=0.21
X4 B.t8 B.t6 B.t7 w_n1294_n2542# sky130_fd_pr__pfet_01v8 ad=3.0615 pd=16.48 as=0 ps=0 w=7.85 l=0.21
X5 B.t5 B.t3 B.t4 w_n1294_n2542# sky130_fd_pr__pfet_01v8 ad=3.0615 pd=16.48 as=0 ps=0 w=7.85 l=0.21
X6 B.t2 B.t0 B.t1 w_n1294_n2542# sky130_fd_pr__pfet_01v8 ad=3.0615 pd=16.48 as=0 ps=0 w=7.85 l=0.21
X7 VDD2.t2 VN.t1 VTAIL.t3 w_n1294_n2542# sky130_fd_pr__pfet_01v8 ad=1.29525 pd=8.18 as=3.0615 ps=16.48 w=7.85 l=0.21
X8 VDD1.t3 VP.t2 VTAIL.t5 w_n1294_n2542# sky130_fd_pr__pfet_01v8 ad=1.29525 pd=8.18 as=3.0615 ps=16.48 w=7.85 l=0.21
X9 VDD2.t1 VN.t2 VTAIL.t1 w_n1294_n2542# sky130_fd_pr__pfet_01v8 ad=1.29525 pd=8.18 as=3.0615 ps=16.48 w=7.85 l=0.21
X10 VTAIL.t4 VP.t3 VDD1.t1 w_n1294_n2542# sky130_fd_pr__pfet_01v8 ad=3.0615 pd=16.48 as=1.29525 ps=8.18 w=7.85 l=0.21
X11 VTAIL.t2 VN.t3 VDD2.t0 w_n1294_n2542# sky130_fd_pr__pfet_01v8 ad=3.0615 pd=16.48 as=1.29525 ps=8.18 w=7.85 l=0.21
R0 B.n76 B.t6 1134.36
R1 B.n84 B.t0 1134.36
R2 B.n24 B.t9 1134.36
R3 B.n30 B.t3 1134.36
R4 B.n270 B.n47 585
R5 B.n272 B.n271 585
R6 B.n273 B.n46 585
R7 B.n275 B.n274 585
R8 B.n276 B.n45 585
R9 B.n278 B.n277 585
R10 B.n279 B.n44 585
R11 B.n281 B.n280 585
R12 B.n282 B.n43 585
R13 B.n284 B.n283 585
R14 B.n285 B.n42 585
R15 B.n287 B.n286 585
R16 B.n288 B.n41 585
R17 B.n290 B.n289 585
R18 B.n291 B.n40 585
R19 B.n293 B.n292 585
R20 B.n294 B.n39 585
R21 B.n296 B.n295 585
R22 B.n297 B.n38 585
R23 B.n299 B.n298 585
R24 B.n300 B.n37 585
R25 B.n302 B.n301 585
R26 B.n303 B.n36 585
R27 B.n305 B.n304 585
R28 B.n306 B.n35 585
R29 B.n308 B.n307 585
R30 B.n309 B.n34 585
R31 B.n311 B.n310 585
R32 B.n312 B.n33 585
R33 B.n314 B.n313 585
R34 B.n316 B.n315 585
R35 B.n317 B.n29 585
R36 B.n319 B.n318 585
R37 B.n320 B.n28 585
R38 B.n322 B.n321 585
R39 B.n323 B.n27 585
R40 B.n325 B.n324 585
R41 B.n326 B.n26 585
R42 B.n328 B.n327 585
R43 B.n330 B.n23 585
R44 B.n332 B.n331 585
R45 B.n333 B.n22 585
R46 B.n335 B.n334 585
R47 B.n336 B.n21 585
R48 B.n338 B.n337 585
R49 B.n339 B.n20 585
R50 B.n341 B.n340 585
R51 B.n342 B.n19 585
R52 B.n344 B.n343 585
R53 B.n345 B.n18 585
R54 B.n347 B.n346 585
R55 B.n348 B.n17 585
R56 B.n350 B.n349 585
R57 B.n351 B.n16 585
R58 B.n353 B.n352 585
R59 B.n354 B.n15 585
R60 B.n356 B.n355 585
R61 B.n357 B.n14 585
R62 B.n359 B.n358 585
R63 B.n360 B.n13 585
R64 B.n362 B.n361 585
R65 B.n363 B.n12 585
R66 B.n365 B.n364 585
R67 B.n366 B.n11 585
R68 B.n368 B.n367 585
R69 B.n369 B.n10 585
R70 B.n371 B.n370 585
R71 B.n372 B.n9 585
R72 B.n374 B.n373 585
R73 B.n269 B.n268 585
R74 B.n267 B.n48 585
R75 B.n266 B.n265 585
R76 B.n264 B.n49 585
R77 B.n263 B.n262 585
R78 B.n261 B.n50 585
R79 B.n260 B.n259 585
R80 B.n258 B.n51 585
R81 B.n257 B.n256 585
R82 B.n255 B.n52 585
R83 B.n254 B.n253 585
R84 B.n252 B.n53 585
R85 B.n251 B.n250 585
R86 B.n249 B.n54 585
R87 B.n248 B.n247 585
R88 B.n246 B.n55 585
R89 B.n245 B.n244 585
R90 B.n243 B.n56 585
R91 B.n242 B.n241 585
R92 B.n240 B.n57 585
R93 B.n239 B.n238 585
R94 B.n237 B.n58 585
R95 B.n236 B.n235 585
R96 B.n234 B.n59 585
R97 B.n233 B.n232 585
R98 B.n231 B.n60 585
R99 B.n230 B.n229 585
R100 B.n125 B.n124 585
R101 B.n126 B.n99 585
R102 B.n128 B.n127 585
R103 B.n129 B.n98 585
R104 B.n131 B.n130 585
R105 B.n132 B.n97 585
R106 B.n134 B.n133 585
R107 B.n135 B.n96 585
R108 B.n137 B.n136 585
R109 B.n138 B.n95 585
R110 B.n140 B.n139 585
R111 B.n141 B.n94 585
R112 B.n143 B.n142 585
R113 B.n144 B.n93 585
R114 B.n146 B.n145 585
R115 B.n147 B.n92 585
R116 B.n149 B.n148 585
R117 B.n150 B.n91 585
R118 B.n152 B.n151 585
R119 B.n153 B.n90 585
R120 B.n155 B.n154 585
R121 B.n156 B.n89 585
R122 B.n158 B.n157 585
R123 B.n159 B.n88 585
R124 B.n161 B.n160 585
R125 B.n162 B.n87 585
R126 B.n164 B.n163 585
R127 B.n165 B.n86 585
R128 B.n167 B.n166 585
R129 B.n168 B.n83 585
R130 B.n171 B.n170 585
R131 B.n172 B.n82 585
R132 B.n174 B.n173 585
R133 B.n175 B.n81 585
R134 B.n177 B.n176 585
R135 B.n178 B.n80 585
R136 B.n180 B.n179 585
R137 B.n181 B.n79 585
R138 B.n183 B.n182 585
R139 B.n185 B.n184 585
R140 B.n186 B.n75 585
R141 B.n188 B.n187 585
R142 B.n189 B.n74 585
R143 B.n191 B.n190 585
R144 B.n192 B.n73 585
R145 B.n194 B.n193 585
R146 B.n195 B.n72 585
R147 B.n197 B.n196 585
R148 B.n198 B.n71 585
R149 B.n200 B.n199 585
R150 B.n201 B.n70 585
R151 B.n203 B.n202 585
R152 B.n204 B.n69 585
R153 B.n206 B.n205 585
R154 B.n207 B.n68 585
R155 B.n209 B.n208 585
R156 B.n210 B.n67 585
R157 B.n212 B.n211 585
R158 B.n213 B.n66 585
R159 B.n215 B.n214 585
R160 B.n216 B.n65 585
R161 B.n218 B.n217 585
R162 B.n219 B.n64 585
R163 B.n221 B.n220 585
R164 B.n222 B.n63 585
R165 B.n224 B.n223 585
R166 B.n225 B.n62 585
R167 B.n227 B.n226 585
R168 B.n228 B.n61 585
R169 B.n123 B.n100 585
R170 B.n122 B.n121 585
R171 B.n120 B.n101 585
R172 B.n119 B.n118 585
R173 B.n117 B.n102 585
R174 B.n116 B.n115 585
R175 B.n114 B.n103 585
R176 B.n113 B.n112 585
R177 B.n111 B.n104 585
R178 B.n110 B.n109 585
R179 B.n108 B.n105 585
R180 B.n107 B.n106 585
R181 B.n2 B.n0 585
R182 B.n393 B.n1 585
R183 B.n392 B.n391 585
R184 B.n390 B.n3 585
R185 B.n389 B.n388 585
R186 B.n387 B.n4 585
R187 B.n386 B.n385 585
R188 B.n384 B.n5 585
R189 B.n383 B.n382 585
R190 B.n381 B.n6 585
R191 B.n380 B.n379 585
R192 B.n378 B.n7 585
R193 B.n377 B.n376 585
R194 B.n375 B.n8 585
R195 B.n395 B.n394 585
R196 B.n124 B.n123 439.647
R197 B.n375 B.n374 439.647
R198 B.n230 B.n61 439.647
R199 B.n268 B.n47 439.647
R200 B.n76 B.t8 311.253
R201 B.n30 B.t4 311.253
R202 B.n84 B.t2 311.253
R203 B.n24 B.t10 311.253
R204 B.n77 B.t7 300.781
R205 B.n31 B.t5 300.781
R206 B.n85 B.t1 300.781
R207 B.n25 B.t11 300.781
R208 B.n123 B.n122 163.367
R209 B.n122 B.n101 163.367
R210 B.n118 B.n101 163.367
R211 B.n118 B.n117 163.367
R212 B.n117 B.n116 163.367
R213 B.n116 B.n103 163.367
R214 B.n112 B.n103 163.367
R215 B.n112 B.n111 163.367
R216 B.n111 B.n110 163.367
R217 B.n110 B.n105 163.367
R218 B.n106 B.n105 163.367
R219 B.n106 B.n2 163.367
R220 B.n394 B.n2 163.367
R221 B.n394 B.n393 163.367
R222 B.n393 B.n392 163.367
R223 B.n392 B.n3 163.367
R224 B.n388 B.n3 163.367
R225 B.n388 B.n387 163.367
R226 B.n387 B.n386 163.367
R227 B.n386 B.n5 163.367
R228 B.n382 B.n5 163.367
R229 B.n382 B.n381 163.367
R230 B.n381 B.n380 163.367
R231 B.n380 B.n7 163.367
R232 B.n376 B.n7 163.367
R233 B.n376 B.n375 163.367
R234 B.n124 B.n99 163.367
R235 B.n128 B.n99 163.367
R236 B.n129 B.n128 163.367
R237 B.n130 B.n129 163.367
R238 B.n130 B.n97 163.367
R239 B.n134 B.n97 163.367
R240 B.n135 B.n134 163.367
R241 B.n136 B.n135 163.367
R242 B.n136 B.n95 163.367
R243 B.n140 B.n95 163.367
R244 B.n141 B.n140 163.367
R245 B.n142 B.n141 163.367
R246 B.n142 B.n93 163.367
R247 B.n146 B.n93 163.367
R248 B.n147 B.n146 163.367
R249 B.n148 B.n147 163.367
R250 B.n148 B.n91 163.367
R251 B.n152 B.n91 163.367
R252 B.n153 B.n152 163.367
R253 B.n154 B.n153 163.367
R254 B.n154 B.n89 163.367
R255 B.n158 B.n89 163.367
R256 B.n159 B.n158 163.367
R257 B.n160 B.n159 163.367
R258 B.n160 B.n87 163.367
R259 B.n164 B.n87 163.367
R260 B.n165 B.n164 163.367
R261 B.n166 B.n165 163.367
R262 B.n166 B.n83 163.367
R263 B.n171 B.n83 163.367
R264 B.n172 B.n171 163.367
R265 B.n173 B.n172 163.367
R266 B.n173 B.n81 163.367
R267 B.n177 B.n81 163.367
R268 B.n178 B.n177 163.367
R269 B.n179 B.n178 163.367
R270 B.n179 B.n79 163.367
R271 B.n183 B.n79 163.367
R272 B.n184 B.n183 163.367
R273 B.n184 B.n75 163.367
R274 B.n188 B.n75 163.367
R275 B.n189 B.n188 163.367
R276 B.n190 B.n189 163.367
R277 B.n190 B.n73 163.367
R278 B.n194 B.n73 163.367
R279 B.n195 B.n194 163.367
R280 B.n196 B.n195 163.367
R281 B.n196 B.n71 163.367
R282 B.n200 B.n71 163.367
R283 B.n201 B.n200 163.367
R284 B.n202 B.n201 163.367
R285 B.n202 B.n69 163.367
R286 B.n206 B.n69 163.367
R287 B.n207 B.n206 163.367
R288 B.n208 B.n207 163.367
R289 B.n208 B.n67 163.367
R290 B.n212 B.n67 163.367
R291 B.n213 B.n212 163.367
R292 B.n214 B.n213 163.367
R293 B.n214 B.n65 163.367
R294 B.n218 B.n65 163.367
R295 B.n219 B.n218 163.367
R296 B.n220 B.n219 163.367
R297 B.n220 B.n63 163.367
R298 B.n224 B.n63 163.367
R299 B.n225 B.n224 163.367
R300 B.n226 B.n225 163.367
R301 B.n226 B.n61 163.367
R302 B.n231 B.n230 163.367
R303 B.n232 B.n231 163.367
R304 B.n232 B.n59 163.367
R305 B.n236 B.n59 163.367
R306 B.n237 B.n236 163.367
R307 B.n238 B.n237 163.367
R308 B.n238 B.n57 163.367
R309 B.n242 B.n57 163.367
R310 B.n243 B.n242 163.367
R311 B.n244 B.n243 163.367
R312 B.n244 B.n55 163.367
R313 B.n248 B.n55 163.367
R314 B.n249 B.n248 163.367
R315 B.n250 B.n249 163.367
R316 B.n250 B.n53 163.367
R317 B.n254 B.n53 163.367
R318 B.n255 B.n254 163.367
R319 B.n256 B.n255 163.367
R320 B.n256 B.n51 163.367
R321 B.n260 B.n51 163.367
R322 B.n261 B.n260 163.367
R323 B.n262 B.n261 163.367
R324 B.n262 B.n49 163.367
R325 B.n266 B.n49 163.367
R326 B.n267 B.n266 163.367
R327 B.n268 B.n267 163.367
R328 B.n374 B.n9 163.367
R329 B.n370 B.n9 163.367
R330 B.n370 B.n369 163.367
R331 B.n369 B.n368 163.367
R332 B.n368 B.n11 163.367
R333 B.n364 B.n11 163.367
R334 B.n364 B.n363 163.367
R335 B.n363 B.n362 163.367
R336 B.n362 B.n13 163.367
R337 B.n358 B.n13 163.367
R338 B.n358 B.n357 163.367
R339 B.n357 B.n356 163.367
R340 B.n356 B.n15 163.367
R341 B.n352 B.n15 163.367
R342 B.n352 B.n351 163.367
R343 B.n351 B.n350 163.367
R344 B.n350 B.n17 163.367
R345 B.n346 B.n17 163.367
R346 B.n346 B.n345 163.367
R347 B.n345 B.n344 163.367
R348 B.n344 B.n19 163.367
R349 B.n340 B.n19 163.367
R350 B.n340 B.n339 163.367
R351 B.n339 B.n338 163.367
R352 B.n338 B.n21 163.367
R353 B.n334 B.n21 163.367
R354 B.n334 B.n333 163.367
R355 B.n333 B.n332 163.367
R356 B.n332 B.n23 163.367
R357 B.n327 B.n23 163.367
R358 B.n327 B.n326 163.367
R359 B.n326 B.n325 163.367
R360 B.n325 B.n27 163.367
R361 B.n321 B.n27 163.367
R362 B.n321 B.n320 163.367
R363 B.n320 B.n319 163.367
R364 B.n319 B.n29 163.367
R365 B.n315 B.n29 163.367
R366 B.n315 B.n314 163.367
R367 B.n314 B.n33 163.367
R368 B.n310 B.n33 163.367
R369 B.n310 B.n309 163.367
R370 B.n309 B.n308 163.367
R371 B.n308 B.n35 163.367
R372 B.n304 B.n35 163.367
R373 B.n304 B.n303 163.367
R374 B.n303 B.n302 163.367
R375 B.n302 B.n37 163.367
R376 B.n298 B.n37 163.367
R377 B.n298 B.n297 163.367
R378 B.n297 B.n296 163.367
R379 B.n296 B.n39 163.367
R380 B.n292 B.n39 163.367
R381 B.n292 B.n291 163.367
R382 B.n291 B.n290 163.367
R383 B.n290 B.n41 163.367
R384 B.n286 B.n41 163.367
R385 B.n286 B.n285 163.367
R386 B.n285 B.n284 163.367
R387 B.n284 B.n43 163.367
R388 B.n280 B.n43 163.367
R389 B.n280 B.n279 163.367
R390 B.n279 B.n278 163.367
R391 B.n278 B.n45 163.367
R392 B.n274 B.n45 163.367
R393 B.n274 B.n273 163.367
R394 B.n273 B.n272 163.367
R395 B.n272 B.n47 163.367
R396 B.n78 B.n77 59.5399
R397 B.n169 B.n85 59.5399
R398 B.n329 B.n25 59.5399
R399 B.n32 B.n31 59.5399
R400 B.n270 B.n269 28.5664
R401 B.n373 B.n8 28.5664
R402 B.n229 B.n228 28.5664
R403 B.n125 B.n100 28.5664
R404 B B.n395 18.0485
R405 B.n373 B.n372 10.6151
R406 B.n372 B.n371 10.6151
R407 B.n371 B.n10 10.6151
R408 B.n367 B.n10 10.6151
R409 B.n367 B.n366 10.6151
R410 B.n366 B.n365 10.6151
R411 B.n365 B.n12 10.6151
R412 B.n361 B.n12 10.6151
R413 B.n361 B.n360 10.6151
R414 B.n360 B.n359 10.6151
R415 B.n359 B.n14 10.6151
R416 B.n355 B.n14 10.6151
R417 B.n355 B.n354 10.6151
R418 B.n354 B.n353 10.6151
R419 B.n353 B.n16 10.6151
R420 B.n349 B.n16 10.6151
R421 B.n349 B.n348 10.6151
R422 B.n348 B.n347 10.6151
R423 B.n347 B.n18 10.6151
R424 B.n343 B.n18 10.6151
R425 B.n343 B.n342 10.6151
R426 B.n342 B.n341 10.6151
R427 B.n341 B.n20 10.6151
R428 B.n337 B.n20 10.6151
R429 B.n337 B.n336 10.6151
R430 B.n336 B.n335 10.6151
R431 B.n335 B.n22 10.6151
R432 B.n331 B.n22 10.6151
R433 B.n331 B.n330 10.6151
R434 B.n328 B.n26 10.6151
R435 B.n324 B.n26 10.6151
R436 B.n324 B.n323 10.6151
R437 B.n323 B.n322 10.6151
R438 B.n322 B.n28 10.6151
R439 B.n318 B.n28 10.6151
R440 B.n318 B.n317 10.6151
R441 B.n317 B.n316 10.6151
R442 B.n313 B.n312 10.6151
R443 B.n312 B.n311 10.6151
R444 B.n311 B.n34 10.6151
R445 B.n307 B.n34 10.6151
R446 B.n307 B.n306 10.6151
R447 B.n306 B.n305 10.6151
R448 B.n305 B.n36 10.6151
R449 B.n301 B.n36 10.6151
R450 B.n301 B.n300 10.6151
R451 B.n300 B.n299 10.6151
R452 B.n299 B.n38 10.6151
R453 B.n295 B.n38 10.6151
R454 B.n295 B.n294 10.6151
R455 B.n294 B.n293 10.6151
R456 B.n293 B.n40 10.6151
R457 B.n289 B.n40 10.6151
R458 B.n289 B.n288 10.6151
R459 B.n288 B.n287 10.6151
R460 B.n287 B.n42 10.6151
R461 B.n283 B.n42 10.6151
R462 B.n283 B.n282 10.6151
R463 B.n282 B.n281 10.6151
R464 B.n281 B.n44 10.6151
R465 B.n277 B.n44 10.6151
R466 B.n277 B.n276 10.6151
R467 B.n276 B.n275 10.6151
R468 B.n275 B.n46 10.6151
R469 B.n271 B.n46 10.6151
R470 B.n271 B.n270 10.6151
R471 B.n229 B.n60 10.6151
R472 B.n233 B.n60 10.6151
R473 B.n234 B.n233 10.6151
R474 B.n235 B.n234 10.6151
R475 B.n235 B.n58 10.6151
R476 B.n239 B.n58 10.6151
R477 B.n240 B.n239 10.6151
R478 B.n241 B.n240 10.6151
R479 B.n241 B.n56 10.6151
R480 B.n245 B.n56 10.6151
R481 B.n246 B.n245 10.6151
R482 B.n247 B.n246 10.6151
R483 B.n247 B.n54 10.6151
R484 B.n251 B.n54 10.6151
R485 B.n252 B.n251 10.6151
R486 B.n253 B.n252 10.6151
R487 B.n253 B.n52 10.6151
R488 B.n257 B.n52 10.6151
R489 B.n258 B.n257 10.6151
R490 B.n259 B.n258 10.6151
R491 B.n259 B.n50 10.6151
R492 B.n263 B.n50 10.6151
R493 B.n264 B.n263 10.6151
R494 B.n265 B.n264 10.6151
R495 B.n265 B.n48 10.6151
R496 B.n269 B.n48 10.6151
R497 B.n126 B.n125 10.6151
R498 B.n127 B.n126 10.6151
R499 B.n127 B.n98 10.6151
R500 B.n131 B.n98 10.6151
R501 B.n132 B.n131 10.6151
R502 B.n133 B.n132 10.6151
R503 B.n133 B.n96 10.6151
R504 B.n137 B.n96 10.6151
R505 B.n138 B.n137 10.6151
R506 B.n139 B.n138 10.6151
R507 B.n139 B.n94 10.6151
R508 B.n143 B.n94 10.6151
R509 B.n144 B.n143 10.6151
R510 B.n145 B.n144 10.6151
R511 B.n145 B.n92 10.6151
R512 B.n149 B.n92 10.6151
R513 B.n150 B.n149 10.6151
R514 B.n151 B.n150 10.6151
R515 B.n151 B.n90 10.6151
R516 B.n155 B.n90 10.6151
R517 B.n156 B.n155 10.6151
R518 B.n157 B.n156 10.6151
R519 B.n157 B.n88 10.6151
R520 B.n161 B.n88 10.6151
R521 B.n162 B.n161 10.6151
R522 B.n163 B.n162 10.6151
R523 B.n163 B.n86 10.6151
R524 B.n167 B.n86 10.6151
R525 B.n168 B.n167 10.6151
R526 B.n170 B.n82 10.6151
R527 B.n174 B.n82 10.6151
R528 B.n175 B.n174 10.6151
R529 B.n176 B.n175 10.6151
R530 B.n176 B.n80 10.6151
R531 B.n180 B.n80 10.6151
R532 B.n181 B.n180 10.6151
R533 B.n182 B.n181 10.6151
R534 B.n186 B.n185 10.6151
R535 B.n187 B.n186 10.6151
R536 B.n187 B.n74 10.6151
R537 B.n191 B.n74 10.6151
R538 B.n192 B.n191 10.6151
R539 B.n193 B.n192 10.6151
R540 B.n193 B.n72 10.6151
R541 B.n197 B.n72 10.6151
R542 B.n198 B.n197 10.6151
R543 B.n199 B.n198 10.6151
R544 B.n199 B.n70 10.6151
R545 B.n203 B.n70 10.6151
R546 B.n204 B.n203 10.6151
R547 B.n205 B.n204 10.6151
R548 B.n205 B.n68 10.6151
R549 B.n209 B.n68 10.6151
R550 B.n210 B.n209 10.6151
R551 B.n211 B.n210 10.6151
R552 B.n211 B.n66 10.6151
R553 B.n215 B.n66 10.6151
R554 B.n216 B.n215 10.6151
R555 B.n217 B.n216 10.6151
R556 B.n217 B.n64 10.6151
R557 B.n221 B.n64 10.6151
R558 B.n222 B.n221 10.6151
R559 B.n223 B.n222 10.6151
R560 B.n223 B.n62 10.6151
R561 B.n227 B.n62 10.6151
R562 B.n228 B.n227 10.6151
R563 B.n121 B.n100 10.6151
R564 B.n121 B.n120 10.6151
R565 B.n120 B.n119 10.6151
R566 B.n119 B.n102 10.6151
R567 B.n115 B.n102 10.6151
R568 B.n115 B.n114 10.6151
R569 B.n114 B.n113 10.6151
R570 B.n113 B.n104 10.6151
R571 B.n109 B.n104 10.6151
R572 B.n109 B.n108 10.6151
R573 B.n108 B.n107 10.6151
R574 B.n107 B.n0 10.6151
R575 B.n391 B.n1 10.6151
R576 B.n391 B.n390 10.6151
R577 B.n390 B.n389 10.6151
R578 B.n389 B.n4 10.6151
R579 B.n385 B.n4 10.6151
R580 B.n385 B.n384 10.6151
R581 B.n384 B.n383 10.6151
R582 B.n383 B.n6 10.6151
R583 B.n379 B.n6 10.6151
R584 B.n379 B.n378 10.6151
R585 B.n378 B.n377 10.6151
R586 B.n377 B.n8 10.6151
R587 B.n77 B.n76 10.4732
R588 B.n85 B.n84 10.4732
R589 B.n25 B.n24 10.4732
R590 B.n31 B.n30 10.4732
R591 B.n329 B.n328 7.18099
R592 B.n316 B.n32 7.18099
R593 B.n170 B.n169 7.18099
R594 B.n182 B.n78 7.18099
R595 B.n330 B.n329 3.43465
R596 B.n313 B.n32 3.43465
R597 B.n169 B.n168 3.43465
R598 B.n185 B.n78 3.43465
R599 B.n395 B.n0 2.81026
R600 B.n395 B.n1 2.81026
R601 VP.n1 VP.t2 1090.66
R602 VP.n1 VP.t3 1090.66
R603 VP.n0 VP.t0 1090.66
R604 VP.n0 VP.t1 1090.66
R605 VP.n2 VP.n0 197.103
R606 VP.n2 VP.n1 161.3
R607 VP VP.n2 0.0516364
R608 VDD1 VDD1.n1 115.749
R609 VDD1 VDD1.n0 83.387
R610 VDD1.n0 VDD1.t2 4.14126
R611 VDD1.n0 VDD1.t0 4.14126
R612 VDD1.n1 VDD1.t1 4.14126
R613 VDD1.n1 VDD1.t3 4.14126
R614 VTAIL.n330 VTAIL.n294 756.745
R615 VTAIL.n36 VTAIL.n0 756.745
R616 VTAIL.n78 VTAIL.n42 756.745
R617 VTAIL.n120 VTAIL.n84 756.745
R618 VTAIL.n288 VTAIL.n252 756.745
R619 VTAIL.n246 VTAIL.n210 756.745
R620 VTAIL.n204 VTAIL.n168 756.745
R621 VTAIL.n162 VTAIL.n126 756.745
R622 VTAIL.n306 VTAIL.n305 585
R623 VTAIL.n311 VTAIL.n310 585
R624 VTAIL.n313 VTAIL.n312 585
R625 VTAIL.n302 VTAIL.n301 585
R626 VTAIL.n319 VTAIL.n318 585
R627 VTAIL.n321 VTAIL.n320 585
R628 VTAIL.n298 VTAIL.n297 585
R629 VTAIL.n328 VTAIL.n327 585
R630 VTAIL.n329 VTAIL.n296 585
R631 VTAIL.n331 VTAIL.n330 585
R632 VTAIL.n12 VTAIL.n11 585
R633 VTAIL.n17 VTAIL.n16 585
R634 VTAIL.n19 VTAIL.n18 585
R635 VTAIL.n8 VTAIL.n7 585
R636 VTAIL.n25 VTAIL.n24 585
R637 VTAIL.n27 VTAIL.n26 585
R638 VTAIL.n4 VTAIL.n3 585
R639 VTAIL.n34 VTAIL.n33 585
R640 VTAIL.n35 VTAIL.n2 585
R641 VTAIL.n37 VTAIL.n36 585
R642 VTAIL.n54 VTAIL.n53 585
R643 VTAIL.n59 VTAIL.n58 585
R644 VTAIL.n61 VTAIL.n60 585
R645 VTAIL.n50 VTAIL.n49 585
R646 VTAIL.n67 VTAIL.n66 585
R647 VTAIL.n69 VTAIL.n68 585
R648 VTAIL.n46 VTAIL.n45 585
R649 VTAIL.n76 VTAIL.n75 585
R650 VTAIL.n77 VTAIL.n44 585
R651 VTAIL.n79 VTAIL.n78 585
R652 VTAIL.n96 VTAIL.n95 585
R653 VTAIL.n101 VTAIL.n100 585
R654 VTAIL.n103 VTAIL.n102 585
R655 VTAIL.n92 VTAIL.n91 585
R656 VTAIL.n109 VTAIL.n108 585
R657 VTAIL.n111 VTAIL.n110 585
R658 VTAIL.n88 VTAIL.n87 585
R659 VTAIL.n118 VTAIL.n117 585
R660 VTAIL.n119 VTAIL.n86 585
R661 VTAIL.n121 VTAIL.n120 585
R662 VTAIL.n289 VTAIL.n288 585
R663 VTAIL.n287 VTAIL.n254 585
R664 VTAIL.n286 VTAIL.n285 585
R665 VTAIL.n257 VTAIL.n255 585
R666 VTAIL.n280 VTAIL.n279 585
R667 VTAIL.n278 VTAIL.n277 585
R668 VTAIL.n261 VTAIL.n260 585
R669 VTAIL.n272 VTAIL.n271 585
R670 VTAIL.n270 VTAIL.n269 585
R671 VTAIL.n265 VTAIL.n264 585
R672 VTAIL.n247 VTAIL.n246 585
R673 VTAIL.n245 VTAIL.n212 585
R674 VTAIL.n244 VTAIL.n243 585
R675 VTAIL.n215 VTAIL.n213 585
R676 VTAIL.n238 VTAIL.n237 585
R677 VTAIL.n236 VTAIL.n235 585
R678 VTAIL.n219 VTAIL.n218 585
R679 VTAIL.n230 VTAIL.n229 585
R680 VTAIL.n228 VTAIL.n227 585
R681 VTAIL.n223 VTAIL.n222 585
R682 VTAIL.n205 VTAIL.n204 585
R683 VTAIL.n203 VTAIL.n170 585
R684 VTAIL.n202 VTAIL.n201 585
R685 VTAIL.n173 VTAIL.n171 585
R686 VTAIL.n196 VTAIL.n195 585
R687 VTAIL.n194 VTAIL.n193 585
R688 VTAIL.n177 VTAIL.n176 585
R689 VTAIL.n188 VTAIL.n187 585
R690 VTAIL.n186 VTAIL.n185 585
R691 VTAIL.n181 VTAIL.n180 585
R692 VTAIL.n163 VTAIL.n162 585
R693 VTAIL.n161 VTAIL.n128 585
R694 VTAIL.n160 VTAIL.n159 585
R695 VTAIL.n131 VTAIL.n129 585
R696 VTAIL.n154 VTAIL.n153 585
R697 VTAIL.n152 VTAIL.n151 585
R698 VTAIL.n135 VTAIL.n134 585
R699 VTAIL.n146 VTAIL.n145 585
R700 VTAIL.n144 VTAIL.n143 585
R701 VTAIL.n139 VTAIL.n138 585
R702 VTAIL.n307 VTAIL.t3 329.043
R703 VTAIL.n13 VTAIL.t0 329.043
R704 VTAIL.n55 VTAIL.t5 329.043
R705 VTAIL.n97 VTAIL.t4 329.043
R706 VTAIL.n266 VTAIL.t6 329.043
R707 VTAIL.n224 VTAIL.t7 329.043
R708 VTAIL.n182 VTAIL.t1 329.043
R709 VTAIL.n140 VTAIL.t2 329.043
R710 VTAIL.n311 VTAIL.n305 171.744
R711 VTAIL.n312 VTAIL.n311 171.744
R712 VTAIL.n312 VTAIL.n301 171.744
R713 VTAIL.n319 VTAIL.n301 171.744
R714 VTAIL.n320 VTAIL.n319 171.744
R715 VTAIL.n320 VTAIL.n297 171.744
R716 VTAIL.n328 VTAIL.n297 171.744
R717 VTAIL.n329 VTAIL.n328 171.744
R718 VTAIL.n330 VTAIL.n329 171.744
R719 VTAIL.n17 VTAIL.n11 171.744
R720 VTAIL.n18 VTAIL.n17 171.744
R721 VTAIL.n18 VTAIL.n7 171.744
R722 VTAIL.n25 VTAIL.n7 171.744
R723 VTAIL.n26 VTAIL.n25 171.744
R724 VTAIL.n26 VTAIL.n3 171.744
R725 VTAIL.n34 VTAIL.n3 171.744
R726 VTAIL.n35 VTAIL.n34 171.744
R727 VTAIL.n36 VTAIL.n35 171.744
R728 VTAIL.n59 VTAIL.n53 171.744
R729 VTAIL.n60 VTAIL.n59 171.744
R730 VTAIL.n60 VTAIL.n49 171.744
R731 VTAIL.n67 VTAIL.n49 171.744
R732 VTAIL.n68 VTAIL.n67 171.744
R733 VTAIL.n68 VTAIL.n45 171.744
R734 VTAIL.n76 VTAIL.n45 171.744
R735 VTAIL.n77 VTAIL.n76 171.744
R736 VTAIL.n78 VTAIL.n77 171.744
R737 VTAIL.n101 VTAIL.n95 171.744
R738 VTAIL.n102 VTAIL.n101 171.744
R739 VTAIL.n102 VTAIL.n91 171.744
R740 VTAIL.n109 VTAIL.n91 171.744
R741 VTAIL.n110 VTAIL.n109 171.744
R742 VTAIL.n110 VTAIL.n87 171.744
R743 VTAIL.n118 VTAIL.n87 171.744
R744 VTAIL.n119 VTAIL.n118 171.744
R745 VTAIL.n120 VTAIL.n119 171.744
R746 VTAIL.n288 VTAIL.n287 171.744
R747 VTAIL.n287 VTAIL.n286 171.744
R748 VTAIL.n286 VTAIL.n255 171.744
R749 VTAIL.n279 VTAIL.n255 171.744
R750 VTAIL.n279 VTAIL.n278 171.744
R751 VTAIL.n278 VTAIL.n260 171.744
R752 VTAIL.n271 VTAIL.n260 171.744
R753 VTAIL.n271 VTAIL.n270 171.744
R754 VTAIL.n270 VTAIL.n264 171.744
R755 VTAIL.n246 VTAIL.n245 171.744
R756 VTAIL.n245 VTAIL.n244 171.744
R757 VTAIL.n244 VTAIL.n213 171.744
R758 VTAIL.n237 VTAIL.n213 171.744
R759 VTAIL.n237 VTAIL.n236 171.744
R760 VTAIL.n236 VTAIL.n218 171.744
R761 VTAIL.n229 VTAIL.n218 171.744
R762 VTAIL.n229 VTAIL.n228 171.744
R763 VTAIL.n228 VTAIL.n222 171.744
R764 VTAIL.n204 VTAIL.n203 171.744
R765 VTAIL.n203 VTAIL.n202 171.744
R766 VTAIL.n202 VTAIL.n171 171.744
R767 VTAIL.n195 VTAIL.n171 171.744
R768 VTAIL.n195 VTAIL.n194 171.744
R769 VTAIL.n194 VTAIL.n176 171.744
R770 VTAIL.n187 VTAIL.n176 171.744
R771 VTAIL.n187 VTAIL.n186 171.744
R772 VTAIL.n186 VTAIL.n180 171.744
R773 VTAIL.n162 VTAIL.n161 171.744
R774 VTAIL.n161 VTAIL.n160 171.744
R775 VTAIL.n160 VTAIL.n129 171.744
R776 VTAIL.n153 VTAIL.n129 171.744
R777 VTAIL.n153 VTAIL.n152 171.744
R778 VTAIL.n152 VTAIL.n134 171.744
R779 VTAIL.n145 VTAIL.n134 171.744
R780 VTAIL.n145 VTAIL.n144 171.744
R781 VTAIL.n144 VTAIL.n138 171.744
R782 VTAIL.t3 VTAIL.n305 85.8723
R783 VTAIL.t0 VTAIL.n11 85.8723
R784 VTAIL.t5 VTAIL.n53 85.8723
R785 VTAIL.t4 VTAIL.n95 85.8723
R786 VTAIL.t6 VTAIL.n264 85.8723
R787 VTAIL.t7 VTAIL.n222 85.8723
R788 VTAIL.t1 VTAIL.n180 85.8723
R789 VTAIL.t2 VTAIL.n138 85.8723
R790 VTAIL.n335 VTAIL.n334 33.155
R791 VTAIL.n41 VTAIL.n40 33.155
R792 VTAIL.n83 VTAIL.n82 33.155
R793 VTAIL.n125 VTAIL.n124 33.155
R794 VTAIL.n293 VTAIL.n292 33.155
R795 VTAIL.n251 VTAIL.n250 33.155
R796 VTAIL.n209 VTAIL.n208 33.155
R797 VTAIL.n167 VTAIL.n166 33.155
R798 VTAIL.n335 VTAIL.n293 19.6169
R799 VTAIL.n167 VTAIL.n125 19.6169
R800 VTAIL.n331 VTAIL.n296 13.1884
R801 VTAIL.n37 VTAIL.n2 13.1884
R802 VTAIL.n79 VTAIL.n44 13.1884
R803 VTAIL.n121 VTAIL.n86 13.1884
R804 VTAIL.n289 VTAIL.n254 13.1884
R805 VTAIL.n247 VTAIL.n212 13.1884
R806 VTAIL.n205 VTAIL.n170 13.1884
R807 VTAIL.n163 VTAIL.n128 13.1884
R808 VTAIL.n327 VTAIL.n326 12.8005
R809 VTAIL.n332 VTAIL.n294 12.8005
R810 VTAIL.n33 VTAIL.n32 12.8005
R811 VTAIL.n38 VTAIL.n0 12.8005
R812 VTAIL.n75 VTAIL.n74 12.8005
R813 VTAIL.n80 VTAIL.n42 12.8005
R814 VTAIL.n117 VTAIL.n116 12.8005
R815 VTAIL.n122 VTAIL.n84 12.8005
R816 VTAIL.n290 VTAIL.n252 12.8005
R817 VTAIL.n285 VTAIL.n256 12.8005
R818 VTAIL.n248 VTAIL.n210 12.8005
R819 VTAIL.n243 VTAIL.n214 12.8005
R820 VTAIL.n206 VTAIL.n168 12.8005
R821 VTAIL.n201 VTAIL.n172 12.8005
R822 VTAIL.n164 VTAIL.n126 12.8005
R823 VTAIL.n159 VTAIL.n130 12.8005
R824 VTAIL.n325 VTAIL.n298 12.0247
R825 VTAIL.n31 VTAIL.n4 12.0247
R826 VTAIL.n73 VTAIL.n46 12.0247
R827 VTAIL.n115 VTAIL.n88 12.0247
R828 VTAIL.n284 VTAIL.n257 12.0247
R829 VTAIL.n242 VTAIL.n215 12.0247
R830 VTAIL.n200 VTAIL.n173 12.0247
R831 VTAIL.n158 VTAIL.n131 12.0247
R832 VTAIL.n322 VTAIL.n321 11.249
R833 VTAIL.n28 VTAIL.n27 11.249
R834 VTAIL.n70 VTAIL.n69 11.249
R835 VTAIL.n112 VTAIL.n111 11.249
R836 VTAIL.n281 VTAIL.n280 11.249
R837 VTAIL.n239 VTAIL.n238 11.249
R838 VTAIL.n197 VTAIL.n196 11.249
R839 VTAIL.n155 VTAIL.n154 11.249
R840 VTAIL.n307 VTAIL.n306 10.7238
R841 VTAIL.n13 VTAIL.n12 10.7238
R842 VTAIL.n55 VTAIL.n54 10.7238
R843 VTAIL.n97 VTAIL.n96 10.7238
R844 VTAIL.n266 VTAIL.n265 10.7238
R845 VTAIL.n224 VTAIL.n223 10.7238
R846 VTAIL.n182 VTAIL.n181 10.7238
R847 VTAIL.n140 VTAIL.n139 10.7238
R848 VTAIL.n318 VTAIL.n300 10.4732
R849 VTAIL.n24 VTAIL.n6 10.4732
R850 VTAIL.n66 VTAIL.n48 10.4732
R851 VTAIL.n108 VTAIL.n90 10.4732
R852 VTAIL.n277 VTAIL.n259 10.4732
R853 VTAIL.n235 VTAIL.n217 10.4732
R854 VTAIL.n193 VTAIL.n175 10.4732
R855 VTAIL.n151 VTAIL.n133 10.4732
R856 VTAIL.n317 VTAIL.n302 9.69747
R857 VTAIL.n23 VTAIL.n8 9.69747
R858 VTAIL.n65 VTAIL.n50 9.69747
R859 VTAIL.n107 VTAIL.n92 9.69747
R860 VTAIL.n276 VTAIL.n261 9.69747
R861 VTAIL.n234 VTAIL.n219 9.69747
R862 VTAIL.n192 VTAIL.n177 9.69747
R863 VTAIL.n150 VTAIL.n135 9.69747
R864 VTAIL.n334 VTAIL.n333 9.45567
R865 VTAIL.n40 VTAIL.n39 9.45567
R866 VTAIL.n82 VTAIL.n81 9.45567
R867 VTAIL.n124 VTAIL.n123 9.45567
R868 VTAIL.n292 VTAIL.n291 9.45567
R869 VTAIL.n250 VTAIL.n249 9.45567
R870 VTAIL.n208 VTAIL.n207 9.45567
R871 VTAIL.n166 VTAIL.n165 9.45567
R872 VTAIL.n333 VTAIL.n332 9.3005
R873 VTAIL.n309 VTAIL.n308 9.3005
R874 VTAIL.n304 VTAIL.n303 9.3005
R875 VTAIL.n315 VTAIL.n314 9.3005
R876 VTAIL.n317 VTAIL.n316 9.3005
R877 VTAIL.n300 VTAIL.n299 9.3005
R878 VTAIL.n323 VTAIL.n322 9.3005
R879 VTAIL.n325 VTAIL.n324 9.3005
R880 VTAIL.n326 VTAIL.n295 9.3005
R881 VTAIL.n39 VTAIL.n38 9.3005
R882 VTAIL.n15 VTAIL.n14 9.3005
R883 VTAIL.n10 VTAIL.n9 9.3005
R884 VTAIL.n21 VTAIL.n20 9.3005
R885 VTAIL.n23 VTAIL.n22 9.3005
R886 VTAIL.n6 VTAIL.n5 9.3005
R887 VTAIL.n29 VTAIL.n28 9.3005
R888 VTAIL.n31 VTAIL.n30 9.3005
R889 VTAIL.n32 VTAIL.n1 9.3005
R890 VTAIL.n81 VTAIL.n80 9.3005
R891 VTAIL.n57 VTAIL.n56 9.3005
R892 VTAIL.n52 VTAIL.n51 9.3005
R893 VTAIL.n63 VTAIL.n62 9.3005
R894 VTAIL.n65 VTAIL.n64 9.3005
R895 VTAIL.n48 VTAIL.n47 9.3005
R896 VTAIL.n71 VTAIL.n70 9.3005
R897 VTAIL.n73 VTAIL.n72 9.3005
R898 VTAIL.n74 VTAIL.n43 9.3005
R899 VTAIL.n123 VTAIL.n122 9.3005
R900 VTAIL.n99 VTAIL.n98 9.3005
R901 VTAIL.n94 VTAIL.n93 9.3005
R902 VTAIL.n105 VTAIL.n104 9.3005
R903 VTAIL.n107 VTAIL.n106 9.3005
R904 VTAIL.n90 VTAIL.n89 9.3005
R905 VTAIL.n113 VTAIL.n112 9.3005
R906 VTAIL.n115 VTAIL.n114 9.3005
R907 VTAIL.n116 VTAIL.n85 9.3005
R908 VTAIL.n268 VTAIL.n267 9.3005
R909 VTAIL.n263 VTAIL.n262 9.3005
R910 VTAIL.n274 VTAIL.n273 9.3005
R911 VTAIL.n276 VTAIL.n275 9.3005
R912 VTAIL.n259 VTAIL.n258 9.3005
R913 VTAIL.n282 VTAIL.n281 9.3005
R914 VTAIL.n284 VTAIL.n283 9.3005
R915 VTAIL.n256 VTAIL.n253 9.3005
R916 VTAIL.n291 VTAIL.n290 9.3005
R917 VTAIL.n226 VTAIL.n225 9.3005
R918 VTAIL.n221 VTAIL.n220 9.3005
R919 VTAIL.n232 VTAIL.n231 9.3005
R920 VTAIL.n234 VTAIL.n233 9.3005
R921 VTAIL.n217 VTAIL.n216 9.3005
R922 VTAIL.n240 VTAIL.n239 9.3005
R923 VTAIL.n242 VTAIL.n241 9.3005
R924 VTAIL.n214 VTAIL.n211 9.3005
R925 VTAIL.n249 VTAIL.n248 9.3005
R926 VTAIL.n184 VTAIL.n183 9.3005
R927 VTAIL.n179 VTAIL.n178 9.3005
R928 VTAIL.n190 VTAIL.n189 9.3005
R929 VTAIL.n192 VTAIL.n191 9.3005
R930 VTAIL.n175 VTAIL.n174 9.3005
R931 VTAIL.n198 VTAIL.n197 9.3005
R932 VTAIL.n200 VTAIL.n199 9.3005
R933 VTAIL.n172 VTAIL.n169 9.3005
R934 VTAIL.n207 VTAIL.n206 9.3005
R935 VTAIL.n142 VTAIL.n141 9.3005
R936 VTAIL.n137 VTAIL.n136 9.3005
R937 VTAIL.n148 VTAIL.n147 9.3005
R938 VTAIL.n150 VTAIL.n149 9.3005
R939 VTAIL.n133 VTAIL.n132 9.3005
R940 VTAIL.n156 VTAIL.n155 9.3005
R941 VTAIL.n158 VTAIL.n157 9.3005
R942 VTAIL.n130 VTAIL.n127 9.3005
R943 VTAIL.n165 VTAIL.n164 9.3005
R944 VTAIL.n314 VTAIL.n313 8.92171
R945 VTAIL.n20 VTAIL.n19 8.92171
R946 VTAIL.n62 VTAIL.n61 8.92171
R947 VTAIL.n104 VTAIL.n103 8.92171
R948 VTAIL.n273 VTAIL.n272 8.92171
R949 VTAIL.n231 VTAIL.n230 8.92171
R950 VTAIL.n189 VTAIL.n188 8.92171
R951 VTAIL.n147 VTAIL.n146 8.92171
R952 VTAIL.n310 VTAIL.n304 8.14595
R953 VTAIL.n16 VTAIL.n10 8.14595
R954 VTAIL.n58 VTAIL.n52 8.14595
R955 VTAIL.n100 VTAIL.n94 8.14595
R956 VTAIL.n269 VTAIL.n263 8.14595
R957 VTAIL.n227 VTAIL.n221 8.14595
R958 VTAIL.n185 VTAIL.n179 8.14595
R959 VTAIL.n143 VTAIL.n137 8.14595
R960 VTAIL.n309 VTAIL.n306 7.3702
R961 VTAIL.n15 VTAIL.n12 7.3702
R962 VTAIL.n57 VTAIL.n54 7.3702
R963 VTAIL.n99 VTAIL.n96 7.3702
R964 VTAIL.n268 VTAIL.n265 7.3702
R965 VTAIL.n226 VTAIL.n223 7.3702
R966 VTAIL.n184 VTAIL.n181 7.3702
R967 VTAIL.n142 VTAIL.n139 7.3702
R968 VTAIL.n310 VTAIL.n309 5.81868
R969 VTAIL.n16 VTAIL.n15 5.81868
R970 VTAIL.n58 VTAIL.n57 5.81868
R971 VTAIL.n100 VTAIL.n99 5.81868
R972 VTAIL.n269 VTAIL.n268 5.81868
R973 VTAIL.n227 VTAIL.n226 5.81868
R974 VTAIL.n185 VTAIL.n184 5.81868
R975 VTAIL.n143 VTAIL.n142 5.81868
R976 VTAIL.n313 VTAIL.n304 5.04292
R977 VTAIL.n19 VTAIL.n10 5.04292
R978 VTAIL.n61 VTAIL.n52 5.04292
R979 VTAIL.n103 VTAIL.n94 5.04292
R980 VTAIL.n272 VTAIL.n263 5.04292
R981 VTAIL.n230 VTAIL.n221 5.04292
R982 VTAIL.n188 VTAIL.n179 5.04292
R983 VTAIL.n146 VTAIL.n137 5.04292
R984 VTAIL.n314 VTAIL.n302 4.26717
R985 VTAIL.n20 VTAIL.n8 4.26717
R986 VTAIL.n62 VTAIL.n50 4.26717
R987 VTAIL.n104 VTAIL.n92 4.26717
R988 VTAIL.n273 VTAIL.n261 4.26717
R989 VTAIL.n231 VTAIL.n219 4.26717
R990 VTAIL.n189 VTAIL.n177 4.26717
R991 VTAIL.n147 VTAIL.n135 4.26717
R992 VTAIL.n318 VTAIL.n317 3.49141
R993 VTAIL.n24 VTAIL.n23 3.49141
R994 VTAIL.n66 VTAIL.n65 3.49141
R995 VTAIL.n108 VTAIL.n107 3.49141
R996 VTAIL.n277 VTAIL.n276 3.49141
R997 VTAIL.n235 VTAIL.n234 3.49141
R998 VTAIL.n193 VTAIL.n192 3.49141
R999 VTAIL.n151 VTAIL.n150 3.49141
R1000 VTAIL.n321 VTAIL.n300 2.71565
R1001 VTAIL.n27 VTAIL.n6 2.71565
R1002 VTAIL.n69 VTAIL.n48 2.71565
R1003 VTAIL.n111 VTAIL.n90 2.71565
R1004 VTAIL.n280 VTAIL.n259 2.71565
R1005 VTAIL.n238 VTAIL.n217 2.71565
R1006 VTAIL.n196 VTAIL.n175 2.71565
R1007 VTAIL.n154 VTAIL.n133 2.71565
R1008 VTAIL.n308 VTAIL.n307 2.4129
R1009 VTAIL.n14 VTAIL.n13 2.4129
R1010 VTAIL.n56 VTAIL.n55 2.4129
R1011 VTAIL.n98 VTAIL.n97 2.4129
R1012 VTAIL.n267 VTAIL.n266 2.4129
R1013 VTAIL.n225 VTAIL.n224 2.4129
R1014 VTAIL.n183 VTAIL.n182 2.4129
R1015 VTAIL.n141 VTAIL.n140 2.4129
R1016 VTAIL.n322 VTAIL.n298 1.93989
R1017 VTAIL.n28 VTAIL.n4 1.93989
R1018 VTAIL.n70 VTAIL.n46 1.93989
R1019 VTAIL.n112 VTAIL.n88 1.93989
R1020 VTAIL.n281 VTAIL.n257 1.93989
R1021 VTAIL.n239 VTAIL.n215 1.93989
R1022 VTAIL.n197 VTAIL.n173 1.93989
R1023 VTAIL.n155 VTAIL.n131 1.93989
R1024 VTAIL.n327 VTAIL.n325 1.16414
R1025 VTAIL.n334 VTAIL.n294 1.16414
R1026 VTAIL.n33 VTAIL.n31 1.16414
R1027 VTAIL.n40 VTAIL.n0 1.16414
R1028 VTAIL.n75 VTAIL.n73 1.16414
R1029 VTAIL.n82 VTAIL.n42 1.16414
R1030 VTAIL.n117 VTAIL.n115 1.16414
R1031 VTAIL.n124 VTAIL.n84 1.16414
R1032 VTAIL.n292 VTAIL.n252 1.16414
R1033 VTAIL.n285 VTAIL.n284 1.16414
R1034 VTAIL.n250 VTAIL.n210 1.16414
R1035 VTAIL.n243 VTAIL.n242 1.16414
R1036 VTAIL.n208 VTAIL.n168 1.16414
R1037 VTAIL.n201 VTAIL.n200 1.16414
R1038 VTAIL.n166 VTAIL.n126 1.16414
R1039 VTAIL.n159 VTAIL.n158 1.16414
R1040 VTAIL.n251 VTAIL.n209 0.470328
R1041 VTAIL.n83 VTAIL.n41 0.470328
R1042 VTAIL.n209 VTAIL.n167 0.466017
R1043 VTAIL.n293 VTAIL.n251 0.466017
R1044 VTAIL.n125 VTAIL.n83 0.466017
R1045 VTAIL.n326 VTAIL.n296 0.388379
R1046 VTAIL.n332 VTAIL.n331 0.388379
R1047 VTAIL.n32 VTAIL.n2 0.388379
R1048 VTAIL.n38 VTAIL.n37 0.388379
R1049 VTAIL.n74 VTAIL.n44 0.388379
R1050 VTAIL.n80 VTAIL.n79 0.388379
R1051 VTAIL.n116 VTAIL.n86 0.388379
R1052 VTAIL.n122 VTAIL.n121 0.388379
R1053 VTAIL.n290 VTAIL.n289 0.388379
R1054 VTAIL.n256 VTAIL.n254 0.388379
R1055 VTAIL.n248 VTAIL.n247 0.388379
R1056 VTAIL.n214 VTAIL.n212 0.388379
R1057 VTAIL.n206 VTAIL.n205 0.388379
R1058 VTAIL.n172 VTAIL.n170 0.388379
R1059 VTAIL.n164 VTAIL.n163 0.388379
R1060 VTAIL.n130 VTAIL.n128 0.388379
R1061 VTAIL VTAIL.n41 0.291448
R1062 VTAIL VTAIL.n335 0.175069
R1063 VTAIL.n308 VTAIL.n303 0.155672
R1064 VTAIL.n315 VTAIL.n303 0.155672
R1065 VTAIL.n316 VTAIL.n315 0.155672
R1066 VTAIL.n316 VTAIL.n299 0.155672
R1067 VTAIL.n323 VTAIL.n299 0.155672
R1068 VTAIL.n324 VTAIL.n323 0.155672
R1069 VTAIL.n324 VTAIL.n295 0.155672
R1070 VTAIL.n333 VTAIL.n295 0.155672
R1071 VTAIL.n14 VTAIL.n9 0.155672
R1072 VTAIL.n21 VTAIL.n9 0.155672
R1073 VTAIL.n22 VTAIL.n21 0.155672
R1074 VTAIL.n22 VTAIL.n5 0.155672
R1075 VTAIL.n29 VTAIL.n5 0.155672
R1076 VTAIL.n30 VTAIL.n29 0.155672
R1077 VTAIL.n30 VTAIL.n1 0.155672
R1078 VTAIL.n39 VTAIL.n1 0.155672
R1079 VTAIL.n56 VTAIL.n51 0.155672
R1080 VTAIL.n63 VTAIL.n51 0.155672
R1081 VTAIL.n64 VTAIL.n63 0.155672
R1082 VTAIL.n64 VTAIL.n47 0.155672
R1083 VTAIL.n71 VTAIL.n47 0.155672
R1084 VTAIL.n72 VTAIL.n71 0.155672
R1085 VTAIL.n72 VTAIL.n43 0.155672
R1086 VTAIL.n81 VTAIL.n43 0.155672
R1087 VTAIL.n98 VTAIL.n93 0.155672
R1088 VTAIL.n105 VTAIL.n93 0.155672
R1089 VTAIL.n106 VTAIL.n105 0.155672
R1090 VTAIL.n106 VTAIL.n89 0.155672
R1091 VTAIL.n113 VTAIL.n89 0.155672
R1092 VTAIL.n114 VTAIL.n113 0.155672
R1093 VTAIL.n114 VTAIL.n85 0.155672
R1094 VTAIL.n123 VTAIL.n85 0.155672
R1095 VTAIL.n291 VTAIL.n253 0.155672
R1096 VTAIL.n283 VTAIL.n253 0.155672
R1097 VTAIL.n283 VTAIL.n282 0.155672
R1098 VTAIL.n282 VTAIL.n258 0.155672
R1099 VTAIL.n275 VTAIL.n258 0.155672
R1100 VTAIL.n275 VTAIL.n274 0.155672
R1101 VTAIL.n274 VTAIL.n262 0.155672
R1102 VTAIL.n267 VTAIL.n262 0.155672
R1103 VTAIL.n249 VTAIL.n211 0.155672
R1104 VTAIL.n241 VTAIL.n211 0.155672
R1105 VTAIL.n241 VTAIL.n240 0.155672
R1106 VTAIL.n240 VTAIL.n216 0.155672
R1107 VTAIL.n233 VTAIL.n216 0.155672
R1108 VTAIL.n233 VTAIL.n232 0.155672
R1109 VTAIL.n232 VTAIL.n220 0.155672
R1110 VTAIL.n225 VTAIL.n220 0.155672
R1111 VTAIL.n207 VTAIL.n169 0.155672
R1112 VTAIL.n199 VTAIL.n169 0.155672
R1113 VTAIL.n199 VTAIL.n198 0.155672
R1114 VTAIL.n198 VTAIL.n174 0.155672
R1115 VTAIL.n191 VTAIL.n174 0.155672
R1116 VTAIL.n191 VTAIL.n190 0.155672
R1117 VTAIL.n190 VTAIL.n178 0.155672
R1118 VTAIL.n183 VTAIL.n178 0.155672
R1119 VTAIL.n165 VTAIL.n127 0.155672
R1120 VTAIL.n157 VTAIL.n127 0.155672
R1121 VTAIL.n157 VTAIL.n156 0.155672
R1122 VTAIL.n156 VTAIL.n132 0.155672
R1123 VTAIL.n149 VTAIL.n132 0.155672
R1124 VTAIL.n149 VTAIL.n148 0.155672
R1125 VTAIL.n148 VTAIL.n136 0.155672
R1126 VTAIL.n141 VTAIL.n136 0.155672
R1127 VN.n0 VN.t1 1090.66
R1128 VN.n0 VN.t0 1090.66
R1129 VN.n1 VN.t3 1090.66
R1130 VN.n1 VN.t2 1090.66
R1131 VN VN.n1 197.484
R1132 VN VN.n0 161.351
R1133 VDD2.n2 VDD2.n0 115.225
R1134 VDD2.n2 VDD2.n1 83.3288
R1135 VDD2.n1 VDD2.t0 4.14126
R1136 VDD2.n1 VDD2.t1 4.14126
R1137 VDD2.n0 VDD2.t3 4.14126
R1138 VDD2.n0 VDD2.t2 4.14126
R1139 VDD2 VDD2.n2 0.0586897
C0 VP VTAIL 0.874833f
C1 VDD1 w_n1294_n2542# 0.834914f
C2 VDD1 VDD2 0.460209f
C3 B VN 0.601459f
C4 VDD1 VTAIL 7.483541f
C5 VDD1 VP 1.32889f
C6 w_n1294_n2542# VN 1.681f
C7 VDD2 VN 1.23364f
C8 VTAIL VN 0.860726f
C9 w_n1294_n2542# B 5.19872f
C10 B VDD2 0.742035f
C11 VP VN 3.69784f
C12 B VTAIL 2.40435f
C13 VDD1 VN 0.147979f
C14 VP B 0.856354f
C15 w_n1294_n2542# VDD2 0.839991f
C16 w_n1294_n2542# VTAIL 3.18136f
C17 VDD2 VTAIL 7.52172f
C18 VDD1 B 0.727191f
C19 VP w_n1294_n2542# 1.8413f
C20 VP VDD2 0.243364f
C21 VDD2 VSUBS 0.510786f
C22 VDD1 VSUBS 4.241596f
C23 VTAIL VSUBS 0.223241f
C24 VN VSUBS 3.72891f
C25 VP VSUBS 0.877413f
C26 B VSUBS 1.852419f
C27 w_n1294_n2542# VSUBS 40.8231f
C28 VDD2.t3 VSUBS 0.186972f
C29 VDD2.t2 VSUBS 0.186972f
C30 VDD2.n0 VSUBS 1.80741f
C31 VDD2.t0 VSUBS 0.186972f
C32 VDD2.t1 VSUBS 0.186972f
C33 VDD2.n1 VSUBS 1.34545f
C34 VDD2.n2 VSUBS 3.54755f
C35 VN.t0 VSUBS 0.189723f
C36 VN.t1 VSUBS 0.189723f
C37 VN.n0 VSUBS 0.175154f
C38 VN.t3 VSUBS 0.189723f
C39 VN.t2 VSUBS 0.189723f
C40 VN.n1 VSUBS 0.408494f
C41 VTAIL.n0 VSUBS 0.026684f
C42 VTAIL.n1 VSUBS 0.026314f
C43 VTAIL.n2 VSUBS 0.014556f
C44 VTAIL.n3 VSUBS 0.033421f
C45 VTAIL.n4 VSUBS 0.014972f
C46 VTAIL.n5 VSUBS 0.026314f
C47 VTAIL.n6 VSUBS 0.01414f
C48 VTAIL.n7 VSUBS 0.033421f
C49 VTAIL.n8 VSUBS 0.014972f
C50 VTAIL.n9 VSUBS 0.026314f
C51 VTAIL.n10 VSUBS 0.01414f
C52 VTAIL.n11 VSUBS 0.025066f
C53 VTAIL.n12 VSUBS 0.025141f
C54 VTAIL.t0 VSUBS 0.071745f
C55 VTAIL.n13 VSUBS 0.157938f
C56 VTAIL.n14 VSUBS 0.814216f
C57 VTAIL.n15 VSUBS 0.01414f
C58 VTAIL.n16 VSUBS 0.014972f
C59 VTAIL.n17 VSUBS 0.033421f
C60 VTAIL.n18 VSUBS 0.033421f
C61 VTAIL.n19 VSUBS 0.014972f
C62 VTAIL.n20 VSUBS 0.01414f
C63 VTAIL.n21 VSUBS 0.026314f
C64 VTAIL.n22 VSUBS 0.026314f
C65 VTAIL.n23 VSUBS 0.01414f
C66 VTAIL.n24 VSUBS 0.014972f
C67 VTAIL.n25 VSUBS 0.033421f
C68 VTAIL.n26 VSUBS 0.033421f
C69 VTAIL.n27 VSUBS 0.014972f
C70 VTAIL.n28 VSUBS 0.01414f
C71 VTAIL.n29 VSUBS 0.026314f
C72 VTAIL.n30 VSUBS 0.026314f
C73 VTAIL.n31 VSUBS 0.01414f
C74 VTAIL.n32 VSUBS 0.01414f
C75 VTAIL.n33 VSUBS 0.014972f
C76 VTAIL.n34 VSUBS 0.033421f
C77 VTAIL.n35 VSUBS 0.033421f
C78 VTAIL.n36 VSUBS 0.073316f
C79 VTAIL.n37 VSUBS 0.014556f
C80 VTAIL.n38 VSUBS 0.01414f
C81 VTAIL.n39 VSUBS 0.06262f
C82 VTAIL.n40 VSUBS 0.036587f
C83 VTAIL.n41 VSUBS 0.087994f
C84 VTAIL.n42 VSUBS 0.026684f
C85 VTAIL.n43 VSUBS 0.026314f
C86 VTAIL.n44 VSUBS 0.014556f
C87 VTAIL.n45 VSUBS 0.033421f
C88 VTAIL.n46 VSUBS 0.014972f
C89 VTAIL.n47 VSUBS 0.026314f
C90 VTAIL.n48 VSUBS 0.01414f
C91 VTAIL.n49 VSUBS 0.033421f
C92 VTAIL.n50 VSUBS 0.014972f
C93 VTAIL.n51 VSUBS 0.026314f
C94 VTAIL.n52 VSUBS 0.01414f
C95 VTAIL.n53 VSUBS 0.025066f
C96 VTAIL.n54 VSUBS 0.025141f
C97 VTAIL.t5 VSUBS 0.071745f
C98 VTAIL.n55 VSUBS 0.157938f
C99 VTAIL.n56 VSUBS 0.814216f
C100 VTAIL.n57 VSUBS 0.01414f
C101 VTAIL.n58 VSUBS 0.014972f
C102 VTAIL.n59 VSUBS 0.033421f
C103 VTAIL.n60 VSUBS 0.033421f
C104 VTAIL.n61 VSUBS 0.014972f
C105 VTAIL.n62 VSUBS 0.01414f
C106 VTAIL.n63 VSUBS 0.026314f
C107 VTAIL.n64 VSUBS 0.026314f
C108 VTAIL.n65 VSUBS 0.01414f
C109 VTAIL.n66 VSUBS 0.014972f
C110 VTAIL.n67 VSUBS 0.033421f
C111 VTAIL.n68 VSUBS 0.033421f
C112 VTAIL.n69 VSUBS 0.014972f
C113 VTAIL.n70 VSUBS 0.01414f
C114 VTAIL.n71 VSUBS 0.026314f
C115 VTAIL.n72 VSUBS 0.026314f
C116 VTAIL.n73 VSUBS 0.01414f
C117 VTAIL.n74 VSUBS 0.01414f
C118 VTAIL.n75 VSUBS 0.014972f
C119 VTAIL.n76 VSUBS 0.033421f
C120 VTAIL.n77 VSUBS 0.033421f
C121 VTAIL.n78 VSUBS 0.073316f
C122 VTAIL.n79 VSUBS 0.014556f
C123 VTAIL.n80 VSUBS 0.01414f
C124 VTAIL.n81 VSUBS 0.06262f
C125 VTAIL.n82 VSUBS 0.036587f
C126 VTAIL.n83 VSUBS 0.102795f
C127 VTAIL.n84 VSUBS 0.026684f
C128 VTAIL.n85 VSUBS 0.026314f
C129 VTAIL.n86 VSUBS 0.014556f
C130 VTAIL.n87 VSUBS 0.033421f
C131 VTAIL.n88 VSUBS 0.014972f
C132 VTAIL.n89 VSUBS 0.026314f
C133 VTAIL.n90 VSUBS 0.01414f
C134 VTAIL.n91 VSUBS 0.033421f
C135 VTAIL.n92 VSUBS 0.014972f
C136 VTAIL.n93 VSUBS 0.026314f
C137 VTAIL.n94 VSUBS 0.01414f
C138 VTAIL.n95 VSUBS 0.025066f
C139 VTAIL.n96 VSUBS 0.025141f
C140 VTAIL.t4 VSUBS 0.071745f
C141 VTAIL.n97 VSUBS 0.157938f
C142 VTAIL.n98 VSUBS 0.814216f
C143 VTAIL.n99 VSUBS 0.01414f
C144 VTAIL.n100 VSUBS 0.014972f
C145 VTAIL.n101 VSUBS 0.033421f
C146 VTAIL.n102 VSUBS 0.033421f
C147 VTAIL.n103 VSUBS 0.014972f
C148 VTAIL.n104 VSUBS 0.01414f
C149 VTAIL.n105 VSUBS 0.026314f
C150 VTAIL.n106 VSUBS 0.026314f
C151 VTAIL.n107 VSUBS 0.01414f
C152 VTAIL.n108 VSUBS 0.014972f
C153 VTAIL.n109 VSUBS 0.033421f
C154 VTAIL.n110 VSUBS 0.033421f
C155 VTAIL.n111 VSUBS 0.014972f
C156 VTAIL.n112 VSUBS 0.01414f
C157 VTAIL.n113 VSUBS 0.026314f
C158 VTAIL.n114 VSUBS 0.026314f
C159 VTAIL.n115 VSUBS 0.01414f
C160 VTAIL.n116 VSUBS 0.01414f
C161 VTAIL.n117 VSUBS 0.014972f
C162 VTAIL.n118 VSUBS 0.033421f
C163 VTAIL.n119 VSUBS 0.033421f
C164 VTAIL.n120 VSUBS 0.073316f
C165 VTAIL.n121 VSUBS 0.014556f
C166 VTAIL.n122 VSUBS 0.01414f
C167 VTAIL.n123 VSUBS 0.06262f
C168 VTAIL.n124 VSUBS 0.036587f
C169 VTAIL.n125 VSUBS 1.03511f
C170 VTAIL.n126 VSUBS 0.026684f
C171 VTAIL.n127 VSUBS 0.026314f
C172 VTAIL.n128 VSUBS 0.014556f
C173 VTAIL.n129 VSUBS 0.033421f
C174 VTAIL.n130 VSUBS 0.01414f
C175 VTAIL.n131 VSUBS 0.014972f
C176 VTAIL.n132 VSUBS 0.026314f
C177 VTAIL.n133 VSUBS 0.01414f
C178 VTAIL.n134 VSUBS 0.033421f
C179 VTAIL.n135 VSUBS 0.014972f
C180 VTAIL.n136 VSUBS 0.026314f
C181 VTAIL.n137 VSUBS 0.01414f
C182 VTAIL.n138 VSUBS 0.025066f
C183 VTAIL.n139 VSUBS 0.025141f
C184 VTAIL.t2 VSUBS 0.071745f
C185 VTAIL.n140 VSUBS 0.157938f
C186 VTAIL.n141 VSUBS 0.814216f
C187 VTAIL.n142 VSUBS 0.01414f
C188 VTAIL.n143 VSUBS 0.014972f
C189 VTAIL.n144 VSUBS 0.033421f
C190 VTAIL.n145 VSUBS 0.033421f
C191 VTAIL.n146 VSUBS 0.014972f
C192 VTAIL.n147 VSUBS 0.01414f
C193 VTAIL.n148 VSUBS 0.026314f
C194 VTAIL.n149 VSUBS 0.026314f
C195 VTAIL.n150 VSUBS 0.01414f
C196 VTAIL.n151 VSUBS 0.014972f
C197 VTAIL.n152 VSUBS 0.033421f
C198 VTAIL.n153 VSUBS 0.033421f
C199 VTAIL.n154 VSUBS 0.014972f
C200 VTAIL.n155 VSUBS 0.01414f
C201 VTAIL.n156 VSUBS 0.026314f
C202 VTAIL.n157 VSUBS 0.026314f
C203 VTAIL.n158 VSUBS 0.01414f
C204 VTAIL.n159 VSUBS 0.014972f
C205 VTAIL.n160 VSUBS 0.033421f
C206 VTAIL.n161 VSUBS 0.033421f
C207 VTAIL.n162 VSUBS 0.073316f
C208 VTAIL.n163 VSUBS 0.014556f
C209 VTAIL.n164 VSUBS 0.01414f
C210 VTAIL.n165 VSUBS 0.06262f
C211 VTAIL.n166 VSUBS 0.036587f
C212 VTAIL.n167 VSUBS 1.03511f
C213 VTAIL.n168 VSUBS 0.026684f
C214 VTAIL.n169 VSUBS 0.026314f
C215 VTAIL.n170 VSUBS 0.014556f
C216 VTAIL.n171 VSUBS 0.033421f
C217 VTAIL.n172 VSUBS 0.01414f
C218 VTAIL.n173 VSUBS 0.014972f
C219 VTAIL.n174 VSUBS 0.026314f
C220 VTAIL.n175 VSUBS 0.01414f
C221 VTAIL.n176 VSUBS 0.033421f
C222 VTAIL.n177 VSUBS 0.014972f
C223 VTAIL.n178 VSUBS 0.026314f
C224 VTAIL.n179 VSUBS 0.01414f
C225 VTAIL.n180 VSUBS 0.025066f
C226 VTAIL.n181 VSUBS 0.025141f
C227 VTAIL.t1 VSUBS 0.071745f
C228 VTAIL.n182 VSUBS 0.157938f
C229 VTAIL.n183 VSUBS 0.814216f
C230 VTAIL.n184 VSUBS 0.01414f
C231 VTAIL.n185 VSUBS 0.014972f
C232 VTAIL.n186 VSUBS 0.033421f
C233 VTAIL.n187 VSUBS 0.033421f
C234 VTAIL.n188 VSUBS 0.014972f
C235 VTAIL.n189 VSUBS 0.01414f
C236 VTAIL.n190 VSUBS 0.026314f
C237 VTAIL.n191 VSUBS 0.026314f
C238 VTAIL.n192 VSUBS 0.01414f
C239 VTAIL.n193 VSUBS 0.014972f
C240 VTAIL.n194 VSUBS 0.033421f
C241 VTAIL.n195 VSUBS 0.033421f
C242 VTAIL.n196 VSUBS 0.014972f
C243 VTAIL.n197 VSUBS 0.01414f
C244 VTAIL.n198 VSUBS 0.026314f
C245 VTAIL.n199 VSUBS 0.026314f
C246 VTAIL.n200 VSUBS 0.01414f
C247 VTAIL.n201 VSUBS 0.014972f
C248 VTAIL.n202 VSUBS 0.033421f
C249 VTAIL.n203 VSUBS 0.033421f
C250 VTAIL.n204 VSUBS 0.073316f
C251 VTAIL.n205 VSUBS 0.014556f
C252 VTAIL.n206 VSUBS 0.01414f
C253 VTAIL.n207 VSUBS 0.06262f
C254 VTAIL.n208 VSUBS 0.036587f
C255 VTAIL.n209 VSUBS 0.102795f
C256 VTAIL.n210 VSUBS 0.026684f
C257 VTAIL.n211 VSUBS 0.026314f
C258 VTAIL.n212 VSUBS 0.014556f
C259 VTAIL.n213 VSUBS 0.033421f
C260 VTAIL.n214 VSUBS 0.01414f
C261 VTAIL.n215 VSUBS 0.014972f
C262 VTAIL.n216 VSUBS 0.026314f
C263 VTAIL.n217 VSUBS 0.01414f
C264 VTAIL.n218 VSUBS 0.033421f
C265 VTAIL.n219 VSUBS 0.014972f
C266 VTAIL.n220 VSUBS 0.026314f
C267 VTAIL.n221 VSUBS 0.01414f
C268 VTAIL.n222 VSUBS 0.025066f
C269 VTAIL.n223 VSUBS 0.025141f
C270 VTAIL.t7 VSUBS 0.071745f
C271 VTAIL.n224 VSUBS 0.157938f
C272 VTAIL.n225 VSUBS 0.814216f
C273 VTAIL.n226 VSUBS 0.01414f
C274 VTAIL.n227 VSUBS 0.014972f
C275 VTAIL.n228 VSUBS 0.033421f
C276 VTAIL.n229 VSUBS 0.033421f
C277 VTAIL.n230 VSUBS 0.014972f
C278 VTAIL.n231 VSUBS 0.01414f
C279 VTAIL.n232 VSUBS 0.026314f
C280 VTAIL.n233 VSUBS 0.026314f
C281 VTAIL.n234 VSUBS 0.01414f
C282 VTAIL.n235 VSUBS 0.014972f
C283 VTAIL.n236 VSUBS 0.033421f
C284 VTAIL.n237 VSUBS 0.033421f
C285 VTAIL.n238 VSUBS 0.014972f
C286 VTAIL.n239 VSUBS 0.01414f
C287 VTAIL.n240 VSUBS 0.026314f
C288 VTAIL.n241 VSUBS 0.026314f
C289 VTAIL.n242 VSUBS 0.01414f
C290 VTAIL.n243 VSUBS 0.014972f
C291 VTAIL.n244 VSUBS 0.033421f
C292 VTAIL.n245 VSUBS 0.033421f
C293 VTAIL.n246 VSUBS 0.073316f
C294 VTAIL.n247 VSUBS 0.014556f
C295 VTAIL.n248 VSUBS 0.01414f
C296 VTAIL.n249 VSUBS 0.06262f
C297 VTAIL.n250 VSUBS 0.036587f
C298 VTAIL.n251 VSUBS 0.102795f
C299 VTAIL.n252 VSUBS 0.026684f
C300 VTAIL.n253 VSUBS 0.026314f
C301 VTAIL.n254 VSUBS 0.014556f
C302 VTAIL.n255 VSUBS 0.033421f
C303 VTAIL.n256 VSUBS 0.01414f
C304 VTAIL.n257 VSUBS 0.014972f
C305 VTAIL.n258 VSUBS 0.026314f
C306 VTAIL.n259 VSUBS 0.01414f
C307 VTAIL.n260 VSUBS 0.033421f
C308 VTAIL.n261 VSUBS 0.014972f
C309 VTAIL.n262 VSUBS 0.026314f
C310 VTAIL.n263 VSUBS 0.01414f
C311 VTAIL.n264 VSUBS 0.025066f
C312 VTAIL.n265 VSUBS 0.025141f
C313 VTAIL.t6 VSUBS 0.071745f
C314 VTAIL.n266 VSUBS 0.157938f
C315 VTAIL.n267 VSUBS 0.814216f
C316 VTAIL.n268 VSUBS 0.01414f
C317 VTAIL.n269 VSUBS 0.014972f
C318 VTAIL.n270 VSUBS 0.033421f
C319 VTAIL.n271 VSUBS 0.033421f
C320 VTAIL.n272 VSUBS 0.014972f
C321 VTAIL.n273 VSUBS 0.01414f
C322 VTAIL.n274 VSUBS 0.026314f
C323 VTAIL.n275 VSUBS 0.026314f
C324 VTAIL.n276 VSUBS 0.01414f
C325 VTAIL.n277 VSUBS 0.014972f
C326 VTAIL.n278 VSUBS 0.033421f
C327 VTAIL.n279 VSUBS 0.033421f
C328 VTAIL.n280 VSUBS 0.014972f
C329 VTAIL.n281 VSUBS 0.01414f
C330 VTAIL.n282 VSUBS 0.026314f
C331 VTAIL.n283 VSUBS 0.026314f
C332 VTAIL.n284 VSUBS 0.01414f
C333 VTAIL.n285 VSUBS 0.014972f
C334 VTAIL.n286 VSUBS 0.033421f
C335 VTAIL.n287 VSUBS 0.033421f
C336 VTAIL.n288 VSUBS 0.073316f
C337 VTAIL.n289 VSUBS 0.014556f
C338 VTAIL.n290 VSUBS 0.01414f
C339 VTAIL.n291 VSUBS 0.06262f
C340 VTAIL.n292 VSUBS 0.036587f
C341 VTAIL.n293 VSUBS 1.03511f
C342 VTAIL.n294 VSUBS 0.026684f
C343 VTAIL.n295 VSUBS 0.026314f
C344 VTAIL.n296 VSUBS 0.014556f
C345 VTAIL.n297 VSUBS 0.033421f
C346 VTAIL.n298 VSUBS 0.014972f
C347 VTAIL.n299 VSUBS 0.026314f
C348 VTAIL.n300 VSUBS 0.01414f
C349 VTAIL.n301 VSUBS 0.033421f
C350 VTAIL.n302 VSUBS 0.014972f
C351 VTAIL.n303 VSUBS 0.026314f
C352 VTAIL.n304 VSUBS 0.01414f
C353 VTAIL.n305 VSUBS 0.025066f
C354 VTAIL.n306 VSUBS 0.025141f
C355 VTAIL.t3 VSUBS 0.071745f
C356 VTAIL.n307 VSUBS 0.157938f
C357 VTAIL.n308 VSUBS 0.814216f
C358 VTAIL.n309 VSUBS 0.01414f
C359 VTAIL.n310 VSUBS 0.014972f
C360 VTAIL.n311 VSUBS 0.033421f
C361 VTAIL.n312 VSUBS 0.033421f
C362 VTAIL.n313 VSUBS 0.014972f
C363 VTAIL.n314 VSUBS 0.01414f
C364 VTAIL.n315 VSUBS 0.026314f
C365 VTAIL.n316 VSUBS 0.026314f
C366 VTAIL.n317 VSUBS 0.01414f
C367 VTAIL.n318 VSUBS 0.014972f
C368 VTAIL.n319 VSUBS 0.033421f
C369 VTAIL.n320 VSUBS 0.033421f
C370 VTAIL.n321 VSUBS 0.014972f
C371 VTAIL.n322 VSUBS 0.01414f
C372 VTAIL.n323 VSUBS 0.026314f
C373 VTAIL.n324 VSUBS 0.026314f
C374 VTAIL.n325 VSUBS 0.01414f
C375 VTAIL.n326 VSUBS 0.01414f
C376 VTAIL.n327 VSUBS 0.014972f
C377 VTAIL.n328 VSUBS 0.033421f
C378 VTAIL.n329 VSUBS 0.033421f
C379 VTAIL.n330 VSUBS 0.073316f
C380 VTAIL.n331 VSUBS 0.014556f
C381 VTAIL.n332 VSUBS 0.01414f
C382 VTAIL.n333 VSUBS 0.06262f
C383 VTAIL.n334 VSUBS 0.036587f
C384 VTAIL.n335 VSUBS 1.01044f
C385 VDD1.t2 VSUBS 0.184238f
C386 VDD1.t0 VSUBS 0.184238f
C387 VDD1.n0 VSUBS 1.32617f
C388 VDD1.t1 VSUBS 0.184238f
C389 VDD1.t3 VSUBS 0.184238f
C390 VDD1.n1 VSUBS 1.80349f
C391 VP.t0 VSUBS 0.192642f
C392 VP.t1 VSUBS 0.192642f
C393 VP.n0 VSUBS 0.407858f
C394 VP.t3 VSUBS 0.192642f
C395 VP.t2 VSUBS 0.192642f
C396 VP.n1 VSUBS 0.177837f
C397 VP.n2 VSUBS 2.32838f
C398 B.n0 VSUBS 0.005971f
C399 B.n1 VSUBS 0.005971f
C400 B.n2 VSUBS 0.009442f
C401 B.n3 VSUBS 0.009442f
C402 B.n4 VSUBS 0.009442f
C403 B.n5 VSUBS 0.009442f
C404 B.n6 VSUBS 0.009442f
C405 B.n7 VSUBS 0.009442f
C406 B.n8 VSUBS 0.019542f
C407 B.n9 VSUBS 0.009442f
C408 B.n10 VSUBS 0.009442f
C409 B.n11 VSUBS 0.009442f
C410 B.n12 VSUBS 0.009442f
C411 B.n13 VSUBS 0.009442f
C412 B.n14 VSUBS 0.009442f
C413 B.n15 VSUBS 0.009442f
C414 B.n16 VSUBS 0.009442f
C415 B.n17 VSUBS 0.009442f
C416 B.n18 VSUBS 0.009442f
C417 B.n19 VSUBS 0.009442f
C418 B.n20 VSUBS 0.009442f
C419 B.n21 VSUBS 0.009442f
C420 B.n22 VSUBS 0.009442f
C421 B.n23 VSUBS 0.009442f
C422 B.t11 VSUBS 0.166519f
C423 B.t10 VSUBS 0.174212f
C424 B.t9 VSUBS 0.087606f
C425 B.n24 VSUBS 0.258394f
C426 B.n25 VSUBS 0.242086f
C427 B.n26 VSUBS 0.009442f
C428 B.n27 VSUBS 0.009442f
C429 B.n28 VSUBS 0.009442f
C430 B.n29 VSUBS 0.009442f
C431 B.t5 VSUBS 0.166523f
C432 B.t4 VSUBS 0.174215f
C433 B.t3 VSUBS 0.087606f
C434 B.n30 VSUBS 0.258391f
C435 B.n31 VSUBS 0.242083f
C436 B.n32 VSUBS 0.021877f
C437 B.n33 VSUBS 0.009442f
C438 B.n34 VSUBS 0.009442f
C439 B.n35 VSUBS 0.009442f
C440 B.n36 VSUBS 0.009442f
C441 B.n37 VSUBS 0.009442f
C442 B.n38 VSUBS 0.009442f
C443 B.n39 VSUBS 0.009442f
C444 B.n40 VSUBS 0.009442f
C445 B.n41 VSUBS 0.009442f
C446 B.n42 VSUBS 0.009442f
C447 B.n43 VSUBS 0.009442f
C448 B.n44 VSUBS 0.009442f
C449 B.n45 VSUBS 0.009442f
C450 B.n46 VSUBS 0.009442f
C451 B.n47 VSUBS 0.021004f
C452 B.n48 VSUBS 0.009442f
C453 B.n49 VSUBS 0.009442f
C454 B.n50 VSUBS 0.009442f
C455 B.n51 VSUBS 0.009442f
C456 B.n52 VSUBS 0.009442f
C457 B.n53 VSUBS 0.009442f
C458 B.n54 VSUBS 0.009442f
C459 B.n55 VSUBS 0.009442f
C460 B.n56 VSUBS 0.009442f
C461 B.n57 VSUBS 0.009442f
C462 B.n58 VSUBS 0.009442f
C463 B.n59 VSUBS 0.009442f
C464 B.n60 VSUBS 0.009442f
C465 B.n61 VSUBS 0.021004f
C466 B.n62 VSUBS 0.009442f
C467 B.n63 VSUBS 0.009442f
C468 B.n64 VSUBS 0.009442f
C469 B.n65 VSUBS 0.009442f
C470 B.n66 VSUBS 0.009442f
C471 B.n67 VSUBS 0.009442f
C472 B.n68 VSUBS 0.009442f
C473 B.n69 VSUBS 0.009442f
C474 B.n70 VSUBS 0.009442f
C475 B.n71 VSUBS 0.009442f
C476 B.n72 VSUBS 0.009442f
C477 B.n73 VSUBS 0.009442f
C478 B.n74 VSUBS 0.009442f
C479 B.n75 VSUBS 0.009442f
C480 B.t7 VSUBS 0.166523f
C481 B.t8 VSUBS 0.174215f
C482 B.t6 VSUBS 0.087606f
C483 B.n76 VSUBS 0.258391f
C484 B.n77 VSUBS 0.242083f
C485 B.n78 VSUBS 0.021877f
C486 B.n79 VSUBS 0.009442f
C487 B.n80 VSUBS 0.009442f
C488 B.n81 VSUBS 0.009442f
C489 B.n82 VSUBS 0.009442f
C490 B.n83 VSUBS 0.009442f
C491 B.t1 VSUBS 0.166519f
C492 B.t2 VSUBS 0.174212f
C493 B.t0 VSUBS 0.087606f
C494 B.n84 VSUBS 0.258394f
C495 B.n85 VSUBS 0.242086f
C496 B.n86 VSUBS 0.009442f
C497 B.n87 VSUBS 0.009442f
C498 B.n88 VSUBS 0.009442f
C499 B.n89 VSUBS 0.009442f
C500 B.n90 VSUBS 0.009442f
C501 B.n91 VSUBS 0.009442f
C502 B.n92 VSUBS 0.009442f
C503 B.n93 VSUBS 0.009442f
C504 B.n94 VSUBS 0.009442f
C505 B.n95 VSUBS 0.009442f
C506 B.n96 VSUBS 0.009442f
C507 B.n97 VSUBS 0.009442f
C508 B.n98 VSUBS 0.009442f
C509 B.n99 VSUBS 0.009442f
C510 B.n100 VSUBS 0.019542f
C511 B.n101 VSUBS 0.009442f
C512 B.n102 VSUBS 0.009442f
C513 B.n103 VSUBS 0.009442f
C514 B.n104 VSUBS 0.009442f
C515 B.n105 VSUBS 0.009442f
C516 B.n106 VSUBS 0.009442f
C517 B.n107 VSUBS 0.009442f
C518 B.n108 VSUBS 0.009442f
C519 B.n109 VSUBS 0.009442f
C520 B.n110 VSUBS 0.009442f
C521 B.n111 VSUBS 0.009442f
C522 B.n112 VSUBS 0.009442f
C523 B.n113 VSUBS 0.009442f
C524 B.n114 VSUBS 0.009442f
C525 B.n115 VSUBS 0.009442f
C526 B.n116 VSUBS 0.009442f
C527 B.n117 VSUBS 0.009442f
C528 B.n118 VSUBS 0.009442f
C529 B.n119 VSUBS 0.009442f
C530 B.n120 VSUBS 0.009442f
C531 B.n121 VSUBS 0.009442f
C532 B.n122 VSUBS 0.009442f
C533 B.n123 VSUBS 0.019542f
C534 B.n124 VSUBS 0.021004f
C535 B.n125 VSUBS 0.021004f
C536 B.n126 VSUBS 0.009442f
C537 B.n127 VSUBS 0.009442f
C538 B.n128 VSUBS 0.009442f
C539 B.n129 VSUBS 0.009442f
C540 B.n130 VSUBS 0.009442f
C541 B.n131 VSUBS 0.009442f
C542 B.n132 VSUBS 0.009442f
C543 B.n133 VSUBS 0.009442f
C544 B.n134 VSUBS 0.009442f
C545 B.n135 VSUBS 0.009442f
C546 B.n136 VSUBS 0.009442f
C547 B.n137 VSUBS 0.009442f
C548 B.n138 VSUBS 0.009442f
C549 B.n139 VSUBS 0.009442f
C550 B.n140 VSUBS 0.009442f
C551 B.n141 VSUBS 0.009442f
C552 B.n142 VSUBS 0.009442f
C553 B.n143 VSUBS 0.009442f
C554 B.n144 VSUBS 0.009442f
C555 B.n145 VSUBS 0.009442f
C556 B.n146 VSUBS 0.009442f
C557 B.n147 VSUBS 0.009442f
C558 B.n148 VSUBS 0.009442f
C559 B.n149 VSUBS 0.009442f
C560 B.n150 VSUBS 0.009442f
C561 B.n151 VSUBS 0.009442f
C562 B.n152 VSUBS 0.009442f
C563 B.n153 VSUBS 0.009442f
C564 B.n154 VSUBS 0.009442f
C565 B.n155 VSUBS 0.009442f
C566 B.n156 VSUBS 0.009442f
C567 B.n157 VSUBS 0.009442f
C568 B.n158 VSUBS 0.009442f
C569 B.n159 VSUBS 0.009442f
C570 B.n160 VSUBS 0.009442f
C571 B.n161 VSUBS 0.009442f
C572 B.n162 VSUBS 0.009442f
C573 B.n163 VSUBS 0.009442f
C574 B.n164 VSUBS 0.009442f
C575 B.n165 VSUBS 0.009442f
C576 B.n166 VSUBS 0.009442f
C577 B.n167 VSUBS 0.009442f
C578 B.n168 VSUBS 0.006249f
C579 B.n169 VSUBS 0.021877f
C580 B.n170 VSUBS 0.007915f
C581 B.n171 VSUBS 0.009442f
C582 B.n172 VSUBS 0.009442f
C583 B.n173 VSUBS 0.009442f
C584 B.n174 VSUBS 0.009442f
C585 B.n175 VSUBS 0.009442f
C586 B.n176 VSUBS 0.009442f
C587 B.n177 VSUBS 0.009442f
C588 B.n178 VSUBS 0.009442f
C589 B.n179 VSUBS 0.009442f
C590 B.n180 VSUBS 0.009442f
C591 B.n181 VSUBS 0.009442f
C592 B.n182 VSUBS 0.007915f
C593 B.n183 VSUBS 0.009442f
C594 B.n184 VSUBS 0.009442f
C595 B.n185 VSUBS 0.006249f
C596 B.n186 VSUBS 0.009442f
C597 B.n187 VSUBS 0.009442f
C598 B.n188 VSUBS 0.009442f
C599 B.n189 VSUBS 0.009442f
C600 B.n190 VSUBS 0.009442f
C601 B.n191 VSUBS 0.009442f
C602 B.n192 VSUBS 0.009442f
C603 B.n193 VSUBS 0.009442f
C604 B.n194 VSUBS 0.009442f
C605 B.n195 VSUBS 0.009442f
C606 B.n196 VSUBS 0.009442f
C607 B.n197 VSUBS 0.009442f
C608 B.n198 VSUBS 0.009442f
C609 B.n199 VSUBS 0.009442f
C610 B.n200 VSUBS 0.009442f
C611 B.n201 VSUBS 0.009442f
C612 B.n202 VSUBS 0.009442f
C613 B.n203 VSUBS 0.009442f
C614 B.n204 VSUBS 0.009442f
C615 B.n205 VSUBS 0.009442f
C616 B.n206 VSUBS 0.009442f
C617 B.n207 VSUBS 0.009442f
C618 B.n208 VSUBS 0.009442f
C619 B.n209 VSUBS 0.009442f
C620 B.n210 VSUBS 0.009442f
C621 B.n211 VSUBS 0.009442f
C622 B.n212 VSUBS 0.009442f
C623 B.n213 VSUBS 0.009442f
C624 B.n214 VSUBS 0.009442f
C625 B.n215 VSUBS 0.009442f
C626 B.n216 VSUBS 0.009442f
C627 B.n217 VSUBS 0.009442f
C628 B.n218 VSUBS 0.009442f
C629 B.n219 VSUBS 0.009442f
C630 B.n220 VSUBS 0.009442f
C631 B.n221 VSUBS 0.009442f
C632 B.n222 VSUBS 0.009442f
C633 B.n223 VSUBS 0.009442f
C634 B.n224 VSUBS 0.009442f
C635 B.n225 VSUBS 0.009442f
C636 B.n226 VSUBS 0.009442f
C637 B.n227 VSUBS 0.009442f
C638 B.n228 VSUBS 0.021004f
C639 B.n229 VSUBS 0.019542f
C640 B.n230 VSUBS 0.019542f
C641 B.n231 VSUBS 0.009442f
C642 B.n232 VSUBS 0.009442f
C643 B.n233 VSUBS 0.009442f
C644 B.n234 VSUBS 0.009442f
C645 B.n235 VSUBS 0.009442f
C646 B.n236 VSUBS 0.009442f
C647 B.n237 VSUBS 0.009442f
C648 B.n238 VSUBS 0.009442f
C649 B.n239 VSUBS 0.009442f
C650 B.n240 VSUBS 0.009442f
C651 B.n241 VSUBS 0.009442f
C652 B.n242 VSUBS 0.009442f
C653 B.n243 VSUBS 0.009442f
C654 B.n244 VSUBS 0.009442f
C655 B.n245 VSUBS 0.009442f
C656 B.n246 VSUBS 0.009442f
C657 B.n247 VSUBS 0.009442f
C658 B.n248 VSUBS 0.009442f
C659 B.n249 VSUBS 0.009442f
C660 B.n250 VSUBS 0.009442f
C661 B.n251 VSUBS 0.009442f
C662 B.n252 VSUBS 0.009442f
C663 B.n253 VSUBS 0.009442f
C664 B.n254 VSUBS 0.009442f
C665 B.n255 VSUBS 0.009442f
C666 B.n256 VSUBS 0.009442f
C667 B.n257 VSUBS 0.009442f
C668 B.n258 VSUBS 0.009442f
C669 B.n259 VSUBS 0.009442f
C670 B.n260 VSUBS 0.009442f
C671 B.n261 VSUBS 0.009442f
C672 B.n262 VSUBS 0.009442f
C673 B.n263 VSUBS 0.009442f
C674 B.n264 VSUBS 0.009442f
C675 B.n265 VSUBS 0.009442f
C676 B.n266 VSUBS 0.009442f
C677 B.n267 VSUBS 0.009442f
C678 B.n268 VSUBS 0.019542f
C679 B.n269 VSUBS 0.020818f
C680 B.n270 VSUBS 0.019729f
C681 B.n271 VSUBS 0.009442f
C682 B.n272 VSUBS 0.009442f
C683 B.n273 VSUBS 0.009442f
C684 B.n274 VSUBS 0.009442f
C685 B.n275 VSUBS 0.009442f
C686 B.n276 VSUBS 0.009442f
C687 B.n277 VSUBS 0.009442f
C688 B.n278 VSUBS 0.009442f
C689 B.n279 VSUBS 0.009442f
C690 B.n280 VSUBS 0.009442f
C691 B.n281 VSUBS 0.009442f
C692 B.n282 VSUBS 0.009442f
C693 B.n283 VSUBS 0.009442f
C694 B.n284 VSUBS 0.009442f
C695 B.n285 VSUBS 0.009442f
C696 B.n286 VSUBS 0.009442f
C697 B.n287 VSUBS 0.009442f
C698 B.n288 VSUBS 0.009442f
C699 B.n289 VSUBS 0.009442f
C700 B.n290 VSUBS 0.009442f
C701 B.n291 VSUBS 0.009442f
C702 B.n292 VSUBS 0.009442f
C703 B.n293 VSUBS 0.009442f
C704 B.n294 VSUBS 0.009442f
C705 B.n295 VSUBS 0.009442f
C706 B.n296 VSUBS 0.009442f
C707 B.n297 VSUBS 0.009442f
C708 B.n298 VSUBS 0.009442f
C709 B.n299 VSUBS 0.009442f
C710 B.n300 VSUBS 0.009442f
C711 B.n301 VSUBS 0.009442f
C712 B.n302 VSUBS 0.009442f
C713 B.n303 VSUBS 0.009442f
C714 B.n304 VSUBS 0.009442f
C715 B.n305 VSUBS 0.009442f
C716 B.n306 VSUBS 0.009442f
C717 B.n307 VSUBS 0.009442f
C718 B.n308 VSUBS 0.009442f
C719 B.n309 VSUBS 0.009442f
C720 B.n310 VSUBS 0.009442f
C721 B.n311 VSUBS 0.009442f
C722 B.n312 VSUBS 0.009442f
C723 B.n313 VSUBS 0.006249f
C724 B.n314 VSUBS 0.009442f
C725 B.n315 VSUBS 0.009442f
C726 B.n316 VSUBS 0.007915f
C727 B.n317 VSUBS 0.009442f
C728 B.n318 VSUBS 0.009442f
C729 B.n319 VSUBS 0.009442f
C730 B.n320 VSUBS 0.009442f
C731 B.n321 VSUBS 0.009442f
C732 B.n322 VSUBS 0.009442f
C733 B.n323 VSUBS 0.009442f
C734 B.n324 VSUBS 0.009442f
C735 B.n325 VSUBS 0.009442f
C736 B.n326 VSUBS 0.009442f
C737 B.n327 VSUBS 0.009442f
C738 B.n328 VSUBS 0.007915f
C739 B.n329 VSUBS 0.021877f
C740 B.n330 VSUBS 0.006249f
C741 B.n331 VSUBS 0.009442f
C742 B.n332 VSUBS 0.009442f
C743 B.n333 VSUBS 0.009442f
C744 B.n334 VSUBS 0.009442f
C745 B.n335 VSUBS 0.009442f
C746 B.n336 VSUBS 0.009442f
C747 B.n337 VSUBS 0.009442f
C748 B.n338 VSUBS 0.009442f
C749 B.n339 VSUBS 0.009442f
C750 B.n340 VSUBS 0.009442f
C751 B.n341 VSUBS 0.009442f
C752 B.n342 VSUBS 0.009442f
C753 B.n343 VSUBS 0.009442f
C754 B.n344 VSUBS 0.009442f
C755 B.n345 VSUBS 0.009442f
C756 B.n346 VSUBS 0.009442f
C757 B.n347 VSUBS 0.009442f
C758 B.n348 VSUBS 0.009442f
C759 B.n349 VSUBS 0.009442f
C760 B.n350 VSUBS 0.009442f
C761 B.n351 VSUBS 0.009442f
C762 B.n352 VSUBS 0.009442f
C763 B.n353 VSUBS 0.009442f
C764 B.n354 VSUBS 0.009442f
C765 B.n355 VSUBS 0.009442f
C766 B.n356 VSUBS 0.009442f
C767 B.n357 VSUBS 0.009442f
C768 B.n358 VSUBS 0.009442f
C769 B.n359 VSUBS 0.009442f
C770 B.n360 VSUBS 0.009442f
C771 B.n361 VSUBS 0.009442f
C772 B.n362 VSUBS 0.009442f
C773 B.n363 VSUBS 0.009442f
C774 B.n364 VSUBS 0.009442f
C775 B.n365 VSUBS 0.009442f
C776 B.n366 VSUBS 0.009442f
C777 B.n367 VSUBS 0.009442f
C778 B.n368 VSUBS 0.009442f
C779 B.n369 VSUBS 0.009442f
C780 B.n370 VSUBS 0.009442f
C781 B.n371 VSUBS 0.009442f
C782 B.n372 VSUBS 0.009442f
C783 B.n373 VSUBS 0.021004f
C784 B.n374 VSUBS 0.021004f
C785 B.n375 VSUBS 0.019542f
C786 B.n376 VSUBS 0.009442f
C787 B.n377 VSUBS 0.009442f
C788 B.n378 VSUBS 0.009442f
C789 B.n379 VSUBS 0.009442f
C790 B.n380 VSUBS 0.009442f
C791 B.n381 VSUBS 0.009442f
C792 B.n382 VSUBS 0.009442f
C793 B.n383 VSUBS 0.009442f
C794 B.n384 VSUBS 0.009442f
C795 B.n385 VSUBS 0.009442f
C796 B.n386 VSUBS 0.009442f
C797 B.n387 VSUBS 0.009442f
C798 B.n388 VSUBS 0.009442f
C799 B.n389 VSUBS 0.009442f
C800 B.n390 VSUBS 0.009442f
C801 B.n391 VSUBS 0.009442f
C802 B.n392 VSUBS 0.009442f
C803 B.n393 VSUBS 0.009442f
C804 B.n394 VSUBS 0.009442f
C805 B.n395 VSUBS 0.021381f
.ends

