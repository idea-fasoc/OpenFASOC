* NGSPICE file created from diff_pair_sample_0003.ext - technology: sky130A

.subckt diff_pair_sample_0003 VTAIL VN VP B VDD2 VDD1
X0 B.t18 B.t16 B.t17 B.t6 sky130_fd_pr__nfet_01v8 ad=3.705 pd=19.78 as=0 ps=0 w=9.5 l=1.61
X1 VDD2.t5 VN.t0 VTAIL.t9 B.t4 sky130_fd_pr__nfet_01v8 ad=3.705 pd=19.78 as=1.5675 ps=9.83 w=9.5 l=1.61
X2 VTAIL.t2 VP.t0 VDD1.t5 B.t0 sky130_fd_pr__nfet_01v8 ad=1.5675 pd=9.83 as=1.5675 ps=9.83 w=9.5 l=1.61
X3 VTAIL.t8 VN.t1 VDD2.t4 B.t19 sky130_fd_pr__nfet_01v8 ad=1.5675 pd=9.83 as=1.5675 ps=9.83 w=9.5 l=1.61
X4 VDD2.t3 VN.t2 VTAIL.t10 B.t1 sky130_fd_pr__nfet_01v8 ad=3.705 pd=19.78 as=1.5675 ps=9.83 w=9.5 l=1.61
X5 B.t15 B.t13 B.t14 B.t10 sky130_fd_pr__nfet_01v8 ad=3.705 pd=19.78 as=0 ps=0 w=9.5 l=1.61
X6 VDD1.t4 VP.t1 VTAIL.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=1.5675 pd=9.83 as=3.705 ps=19.78 w=9.5 l=1.61
X7 VDD1.t3 VP.t2 VTAIL.t5 B.t1 sky130_fd_pr__nfet_01v8 ad=3.705 pd=19.78 as=1.5675 ps=9.83 w=9.5 l=1.61
X8 VDD2.t2 VN.t3 VTAIL.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=1.5675 pd=9.83 as=3.705 ps=19.78 w=9.5 l=1.61
X9 VDD1.t2 VP.t3 VTAIL.t3 B.t4 sky130_fd_pr__nfet_01v8 ad=3.705 pd=19.78 as=1.5675 ps=9.83 w=9.5 l=1.61
X10 VDD2.t1 VN.t4 VTAIL.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=1.5675 pd=9.83 as=3.705 ps=19.78 w=9.5 l=1.61
X11 VDD1.t1 VP.t4 VTAIL.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=1.5675 pd=9.83 as=3.705 ps=19.78 w=9.5 l=1.61
X12 VTAIL.t7 VN.t5 VDD2.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.5675 pd=9.83 as=1.5675 ps=9.83 w=9.5 l=1.61
X13 B.t12 B.t9 B.t11 B.t10 sky130_fd_pr__nfet_01v8 ad=3.705 pd=19.78 as=0 ps=0 w=9.5 l=1.61
X14 VTAIL.t4 VP.t5 VDD1.t0 B.t19 sky130_fd_pr__nfet_01v8 ad=1.5675 pd=9.83 as=1.5675 ps=9.83 w=9.5 l=1.61
X15 B.t8 B.t5 B.t7 B.t6 sky130_fd_pr__nfet_01v8 ad=3.705 pd=19.78 as=0 ps=0 w=9.5 l=1.61
R0 B.n648 B.n647 585
R1 B.n254 B.n98 585
R2 B.n253 B.n252 585
R3 B.n251 B.n250 585
R4 B.n249 B.n248 585
R5 B.n247 B.n246 585
R6 B.n245 B.n244 585
R7 B.n243 B.n242 585
R8 B.n241 B.n240 585
R9 B.n239 B.n238 585
R10 B.n237 B.n236 585
R11 B.n235 B.n234 585
R12 B.n233 B.n232 585
R13 B.n231 B.n230 585
R14 B.n229 B.n228 585
R15 B.n227 B.n226 585
R16 B.n225 B.n224 585
R17 B.n223 B.n222 585
R18 B.n221 B.n220 585
R19 B.n219 B.n218 585
R20 B.n217 B.n216 585
R21 B.n215 B.n214 585
R22 B.n213 B.n212 585
R23 B.n211 B.n210 585
R24 B.n209 B.n208 585
R25 B.n207 B.n206 585
R26 B.n205 B.n204 585
R27 B.n203 B.n202 585
R28 B.n201 B.n200 585
R29 B.n199 B.n198 585
R30 B.n197 B.n196 585
R31 B.n195 B.n194 585
R32 B.n193 B.n192 585
R33 B.n191 B.n190 585
R34 B.n189 B.n188 585
R35 B.n187 B.n186 585
R36 B.n185 B.n184 585
R37 B.n183 B.n182 585
R38 B.n181 B.n180 585
R39 B.n179 B.n178 585
R40 B.n177 B.n176 585
R41 B.n175 B.n174 585
R42 B.n173 B.n172 585
R43 B.n171 B.n170 585
R44 B.n169 B.n168 585
R45 B.n167 B.n166 585
R46 B.n165 B.n164 585
R47 B.n163 B.n162 585
R48 B.n161 B.n160 585
R49 B.n159 B.n158 585
R50 B.n157 B.n156 585
R51 B.n155 B.n154 585
R52 B.n153 B.n152 585
R53 B.n151 B.n150 585
R54 B.n149 B.n148 585
R55 B.n147 B.n146 585
R56 B.n145 B.n144 585
R57 B.n143 B.n142 585
R58 B.n141 B.n140 585
R59 B.n139 B.n138 585
R60 B.n137 B.n136 585
R61 B.n135 B.n134 585
R62 B.n133 B.n132 585
R63 B.n131 B.n130 585
R64 B.n129 B.n128 585
R65 B.n127 B.n126 585
R66 B.n125 B.n124 585
R67 B.n123 B.n122 585
R68 B.n121 B.n120 585
R69 B.n119 B.n118 585
R70 B.n117 B.n116 585
R71 B.n115 B.n114 585
R72 B.n113 B.n112 585
R73 B.n111 B.n110 585
R74 B.n109 B.n108 585
R75 B.n107 B.n106 585
R76 B.n60 B.n59 585
R77 B.n653 B.n652 585
R78 B.n646 B.n99 585
R79 B.n99 B.n57 585
R80 B.n645 B.n56 585
R81 B.n657 B.n56 585
R82 B.n644 B.n55 585
R83 B.n658 B.n55 585
R84 B.n643 B.n54 585
R85 B.n659 B.n54 585
R86 B.n642 B.n641 585
R87 B.n641 B.n50 585
R88 B.n640 B.n49 585
R89 B.n665 B.n49 585
R90 B.n639 B.n48 585
R91 B.n666 B.n48 585
R92 B.n638 B.n47 585
R93 B.n667 B.n47 585
R94 B.n637 B.n636 585
R95 B.n636 B.n43 585
R96 B.n635 B.n42 585
R97 B.n673 B.n42 585
R98 B.n634 B.n41 585
R99 B.n674 B.n41 585
R100 B.n633 B.n40 585
R101 B.n675 B.n40 585
R102 B.n632 B.n631 585
R103 B.n631 B.n36 585
R104 B.n630 B.n35 585
R105 B.n681 B.n35 585
R106 B.n629 B.n34 585
R107 B.n682 B.n34 585
R108 B.n628 B.n33 585
R109 B.n683 B.n33 585
R110 B.n627 B.n626 585
R111 B.n626 B.n29 585
R112 B.n625 B.n28 585
R113 B.n689 B.n28 585
R114 B.n624 B.n27 585
R115 B.n690 B.n27 585
R116 B.n623 B.n26 585
R117 B.n691 B.n26 585
R118 B.n622 B.n621 585
R119 B.n621 B.n25 585
R120 B.n620 B.n21 585
R121 B.n697 B.n21 585
R122 B.n619 B.n20 585
R123 B.n698 B.n20 585
R124 B.n618 B.n19 585
R125 B.n699 B.n19 585
R126 B.n617 B.n616 585
R127 B.n616 B.n15 585
R128 B.n615 B.n14 585
R129 B.n705 B.n14 585
R130 B.n614 B.n13 585
R131 B.n706 B.n13 585
R132 B.n613 B.n12 585
R133 B.n707 B.n12 585
R134 B.n612 B.n611 585
R135 B.n611 B.n8 585
R136 B.n610 B.n7 585
R137 B.n713 B.n7 585
R138 B.n609 B.n6 585
R139 B.n714 B.n6 585
R140 B.n608 B.n5 585
R141 B.n715 B.n5 585
R142 B.n607 B.n606 585
R143 B.n606 B.n4 585
R144 B.n605 B.n255 585
R145 B.n605 B.n604 585
R146 B.n595 B.n256 585
R147 B.n257 B.n256 585
R148 B.n597 B.n596 585
R149 B.n598 B.n597 585
R150 B.n594 B.n261 585
R151 B.n265 B.n261 585
R152 B.n593 B.n592 585
R153 B.n592 B.n591 585
R154 B.n263 B.n262 585
R155 B.n264 B.n263 585
R156 B.n584 B.n583 585
R157 B.n585 B.n584 585
R158 B.n582 B.n270 585
R159 B.n270 B.n269 585
R160 B.n581 B.n580 585
R161 B.n580 B.n579 585
R162 B.n272 B.n271 585
R163 B.n572 B.n272 585
R164 B.n571 B.n570 585
R165 B.n573 B.n571 585
R166 B.n569 B.n277 585
R167 B.n277 B.n276 585
R168 B.n568 B.n567 585
R169 B.n567 B.n566 585
R170 B.n279 B.n278 585
R171 B.n280 B.n279 585
R172 B.n559 B.n558 585
R173 B.n560 B.n559 585
R174 B.n557 B.n285 585
R175 B.n285 B.n284 585
R176 B.n556 B.n555 585
R177 B.n555 B.n554 585
R178 B.n287 B.n286 585
R179 B.n288 B.n287 585
R180 B.n547 B.n546 585
R181 B.n548 B.n547 585
R182 B.n545 B.n293 585
R183 B.n293 B.n292 585
R184 B.n544 B.n543 585
R185 B.n543 B.n542 585
R186 B.n295 B.n294 585
R187 B.n296 B.n295 585
R188 B.n535 B.n534 585
R189 B.n536 B.n535 585
R190 B.n533 B.n300 585
R191 B.n304 B.n300 585
R192 B.n532 B.n531 585
R193 B.n531 B.n530 585
R194 B.n302 B.n301 585
R195 B.n303 B.n302 585
R196 B.n523 B.n522 585
R197 B.n524 B.n523 585
R198 B.n521 B.n309 585
R199 B.n309 B.n308 585
R200 B.n520 B.n519 585
R201 B.n519 B.n518 585
R202 B.n311 B.n310 585
R203 B.n312 B.n311 585
R204 B.n514 B.n513 585
R205 B.n315 B.n314 585
R206 B.n510 B.n509 585
R207 B.n511 B.n510 585
R208 B.n508 B.n354 585
R209 B.n507 B.n506 585
R210 B.n505 B.n504 585
R211 B.n503 B.n502 585
R212 B.n501 B.n500 585
R213 B.n499 B.n498 585
R214 B.n497 B.n496 585
R215 B.n495 B.n494 585
R216 B.n493 B.n492 585
R217 B.n491 B.n490 585
R218 B.n489 B.n488 585
R219 B.n487 B.n486 585
R220 B.n485 B.n484 585
R221 B.n483 B.n482 585
R222 B.n481 B.n480 585
R223 B.n479 B.n478 585
R224 B.n477 B.n476 585
R225 B.n475 B.n474 585
R226 B.n473 B.n472 585
R227 B.n471 B.n470 585
R228 B.n469 B.n468 585
R229 B.n467 B.n466 585
R230 B.n465 B.n464 585
R231 B.n463 B.n462 585
R232 B.n461 B.n460 585
R233 B.n459 B.n458 585
R234 B.n457 B.n456 585
R235 B.n455 B.n454 585
R236 B.n453 B.n452 585
R237 B.n451 B.n450 585
R238 B.n449 B.n448 585
R239 B.n446 B.n445 585
R240 B.n444 B.n443 585
R241 B.n442 B.n441 585
R242 B.n440 B.n439 585
R243 B.n438 B.n437 585
R244 B.n436 B.n435 585
R245 B.n434 B.n433 585
R246 B.n432 B.n431 585
R247 B.n430 B.n429 585
R248 B.n428 B.n427 585
R249 B.n425 B.n424 585
R250 B.n423 B.n422 585
R251 B.n421 B.n420 585
R252 B.n419 B.n418 585
R253 B.n417 B.n416 585
R254 B.n415 B.n414 585
R255 B.n413 B.n412 585
R256 B.n411 B.n410 585
R257 B.n409 B.n408 585
R258 B.n407 B.n406 585
R259 B.n405 B.n404 585
R260 B.n403 B.n402 585
R261 B.n401 B.n400 585
R262 B.n399 B.n398 585
R263 B.n397 B.n396 585
R264 B.n395 B.n394 585
R265 B.n393 B.n392 585
R266 B.n391 B.n390 585
R267 B.n389 B.n388 585
R268 B.n387 B.n386 585
R269 B.n385 B.n384 585
R270 B.n383 B.n382 585
R271 B.n381 B.n380 585
R272 B.n379 B.n378 585
R273 B.n377 B.n376 585
R274 B.n375 B.n374 585
R275 B.n373 B.n372 585
R276 B.n371 B.n370 585
R277 B.n369 B.n368 585
R278 B.n367 B.n366 585
R279 B.n365 B.n364 585
R280 B.n363 B.n362 585
R281 B.n361 B.n360 585
R282 B.n359 B.n353 585
R283 B.n511 B.n353 585
R284 B.n515 B.n313 585
R285 B.n313 B.n312 585
R286 B.n517 B.n516 585
R287 B.n518 B.n517 585
R288 B.n307 B.n306 585
R289 B.n308 B.n307 585
R290 B.n526 B.n525 585
R291 B.n525 B.n524 585
R292 B.n527 B.n305 585
R293 B.n305 B.n303 585
R294 B.n529 B.n528 585
R295 B.n530 B.n529 585
R296 B.n299 B.n298 585
R297 B.n304 B.n299 585
R298 B.n538 B.n537 585
R299 B.n537 B.n536 585
R300 B.n539 B.n297 585
R301 B.n297 B.n296 585
R302 B.n541 B.n540 585
R303 B.n542 B.n541 585
R304 B.n291 B.n290 585
R305 B.n292 B.n291 585
R306 B.n550 B.n549 585
R307 B.n549 B.n548 585
R308 B.n551 B.n289 585
R309 B.n289 B.n288 585
R310 B.n553 B.n552 585
R311 B.n554 B.n553 585
R312 B.n283 B.n282 585
R313 B.n284 B.n283 585
R314 B.n562 B.n561 585
R315 B.n561 B.n560 585
R316 B.n563 B.n281 585
R317 B.n281 B.n280 585
R318 B.n565 B.n564 585
R319 B.n566 B.n565 585
R320 B.n275 B.n274 585
R321 B.n276 B.n275 585
R322 B.n575 B.n574 585
R323 B.n574 B.n573 585
R324 B.n576 B.n273 585
R325 B.n572 B.n273 585
R326 B.n578 B.n577 585
R327 B.n579 B.n578 585
R328 B.n268 B.n267 585
R329 B.n269 B.n268 585
R330 B.n587 B.n586 585
R331 B.n586 B.n585 585
R332 B.n588 B.n266 585
R333 B.n266 B.n264 585
R334 B.n590 B.n589 585
R335 B.n591 B.n590 585
R336 B.n260 B.n259 585
R337 B.n265 B.n260 585
R338 B.n600 B.n599 585
R339 B.n599 B.n598 585
R340 B.n601 B.n258 585
R341 B.n258 B.n257 585
R342 B.n603 B.n602 585
R343 B.n604 B.n603 585
R344 B.n2 B.n0 585
R345 B.n4 B.n2 585
R346 B.n3 B.n1 585
R347 B.n714 B.n3 585
R348 B.n712 B.n711 585
R349 B.n713 B.n712 585
R350 B.n710 B.n9 585
R351 B.n9 B.n8 585
R352 B.n709 B.n708 585
R353 B.n708 B.n707 585
R354 B.n11 B.n10 585
R355 B.n706 B.n11 585
R356 B.n704 B.n703 585
R357 B.n705 B.n704 585
R358 B.n702 B.n16 585
R359 B.n16 B.n15 585
R360 B.n701 B.n700 585
R361 B.n700 B.n699 585
R362 B.n18 B.n17 585
R363 B.n698 B.n18 585
R364 B.n696 B.n695 585
R365 B.n697 B.n696 585
R366 B.n694 B.n22 585
R367 B.n25 B.n22 585
R368 B.n693 B.n692 585
R369 B.n692 B.n691 585
R370 B.n24 B.n23 585
R371 B.n690 B.n24 585
R372 B.n688 B.n687 585
R373 B.n689 B.n688 585
R374 B.n686 B.n30 585
R375 B.n30 B.n29 585
R376 B.n685 B.n684 585
R377 B.n684 B.n683 585
R378 B.n32 B.n31 585
R379 B.n682 B.n32 585
R380 B.n680 B.n679 585
R381 B.n681 B.n680 585
R382 B.n678 B.n37 585
R383 B.n37 B.n36 585
R384 B.n677 B.n676 585
R385 B.n676 B.n675 585
R386 B.n39 B.n38 585
R387 B.n674 B.n39 585
R388 B.n672 B.n671 585
R389 B.n673 B.n672 585
R390 B.n670 B.n44 585
R391 B.n44 B.n43 585
R392 B.n669 B.n668 585
R393 B.n668 B.n667 585
R394 B.n46 B.n45 585
R395 B.n666 B.n46 585
R396 B.n664 B.n663 585
R397 B.n665 B.n664 585
R398 B.n662 B.n51 585
R399 B.n51 B.n50 585
R400 B.n661 B.n660 585
R401 B.n660 B.n659 585
R402 B.n53 B.n52 585
R403 B.n658 B.n53 585
R404 B.n656 B.n655 585
R405 B.n657 B.n656 585
R406 B.n654 B.n58 585
R407 B.n58 B.n57 585
R408 B.n717 B.n716 585
R409 B.n716 B.n715 585
R410 B.n513 B.n313 497.305
R411 B.n652 B.n58 497.305
R412 B.n353 B.n311 497.305
R413 B.n648 B.n99 497.305
R414 B.n357 B.t9 348.033
R415 B.n355 B.t13 348.033
R416 B.n103 B.t16 348.033
R417 B.n100 B.t5 348.033
R418 B.n357 B.t12 277.05
R419 B.n100 B.t7 277.05
R420 B.n355 B.t15 277.05
R421 B.n103 B.t17 277.05
R422 B.n650 B.n649 256.663
R423 B.n650 B.n97 256.663
R424 B.n650 B.n96 256.663
R425 B.n650 B.n95 256.663
R426 B.n650 B.n94 256.663
R427 B.n650 B.n93 256.663
R428 B.n650 B.n92 256.663
R429 B.n650 B.n91 256.663
R430 B.n650 B.n90 256.663
R431 B.n650 B.n89 256.663
R432 B.n650 B.n88 256.663
R433 B.n650 B.n87 256.663
R434 B.n650 B.n86 256.663
R435 B.n650 B.n85 256.663
R436 B.n650 B.n84 256.663
R437 B.n650 B.n83 256.663
R438 B.n650 B.n82 256.663
R439 B.n650 B.n81 256.663
R440 B.n650 B.n80 256.663
R441 B.n650 B.n79 256.663
R442 B.n650 B.n78 256.663
R443 B.n650 B.n77 256.663
R444 B.n650 B.n76 256.663
R445 B.n650 B.n75 256.663
R446 B.n650 B.n74 256.663
R447 B.n650 B.n73 256.663
R448 B.n650 B.n72 256.663
R449 B.n650 B.n71 256.663
R450 B.n650 B.n70 256.663
R451 B.n650 B.n69 256.663
R452 B.n650 B.n68 256.663
R453 B.n650 B.n67 256.663
R454 B.n650 B.n66 256.663
R455 B.n650 B.n65 256.663
R456 B.n650 B.n64 256.663
R457 B.n650 B.n63 256.663
R458 B.n650 B.n62 256.663
R459 B.n650 B.n61 256.663
R460 B.n651 B.n650 256.663
R461 B.n512 B.n511 256.663
R462 B.n511 B.n316 256.663
R463 B.n511 B.n317 256.663
R464 B.n511 B.n318 256.663
R465 B.n511 B.n319 256.663
R466 B.n511 B.n320 256.663
R467 B.n511 B.n321 256.663
R468 B.n511 B.n322 256.663
R469 B.n511 B.n323 256.663
R470 B.n511 B.n324 256.663
R471 B.n511 B.n325 256.663
R472 B.n511 B.n326 256.663
R473 B.n511 B.n327 256.663
R474 B.n511 B.n328 256.663
R475 B.n511 B.n329 256.663
R476 B.n511 B.n330 256.663
R477 B.n511 B.n331 256.663
R478 B.n511 B.n332 256.663
R479 B.n511 B.n333 256.663
R480 B.n511 B.n334 256.663
R481 B.n511 B.n335 256.663
R482 B.n511 B.n336 256.663
R483 B.n511 B.n337 256.663
R484 B.n511 B.n338 256.663
R485 B.n511 B.n339 256.663
R486 B.n511 B.n340 256.663
R487 B.n511 B.n341 256.663
R488 B.n511 B.n342 256.663
R489 B.n511 B.n343 256.663
R490 B.n511 B.n344 256.663
R491 B.n511 B.n345 256.663
R492 B.n511 B.n346 256.663
R493 B.n511 B.n347 256.663
R494 B.n511 B.n348 256.663
R495 B.n511 B.n349 256.663
R496 B.n511 B.n350 256.663
R497 B.n511 B.n351 256.663
R498 B.n511 B.n352 256.663
R499 B.n358 B.t11 239.427
R500 B.n101 B.t8 239.427
R501 B.n356 B.t14 239.427
R502 B.n104 B.t18 239.427
R503 B.n517 B.n313 163.367
R504 B.n517 B.n307 163.367
R505 B.n525 B.n307 163.367
R506 B.n525 B.n305 163.367
R507 B.n529 B.n305 163.367
R508 B.n529 B.n299 163.367
R509 B.n537 B.n299 163.367
R510 B.n537 B.n297 163.367
R511 B.n541 B.n297 163.367
R512 B.n541 B.n291 163.367
R513 B.n549 B.n291 163.367
R514 B.n549 B.n289 163.367
R515 B.n553 B.n289 163.367
R516 B.n553 B.n283 163.367
R517 B.n561 B.n283 163.367
R518 B.n561 B.n281 163.367
R519 B.n565 B.n281 163.367
R520 B.n565 B.n275 163.367
R521 B.n574 B.n275 163.367
R522 B.n574 B.n273 163.367
R523 B.n578 B.n273 163.367
R524 B.n578 B.n268 163.367
R525 B.n586 B.n268 163.367
R526 B.n586 B.n266 163.367
R527 B.n590 B.n266 163.367
R528 B.n590 B.n260 163.367
R529 B.n599 B.n260 163.367
R530 B.n599 B.n258 163.367
R531 B.n603 B.n258 163.367
R532 B.n603 B.n2 163.367
R533 B.n716 B.n2 163.367
R534 B.n716 B.n3 163.367
R535 B.n712 B.n3 163.367
R536 B.n712 B.n9 163.367
R537 B.n708 B.n9 163.367
R538 B.n708 B.n11 163.367
R539 B.n704 B.n11 163.367
R540 B.n704 B.n16 163.367
R541 B.n700 B.n16 163.367
R542 B.n700 B.n18 163.367
R543 B.n696 B.n18 163.367
R544 B.n696 B.n22 163.367
R545 B.n692 B.n22 163.367
R546 B.n692 B.n24 163.367
R547 B.n688 B.n24 163.367
R548 B.n688 B.n30 163.367
R549 B.n684 B.n30 163.367
R550 B.n684 B.n32 163.367
R551 B.n680 B.n32 163.367
R552 B.n680 B.n37 163.367
R553 B.n676 B.n37 163.367
R554 B.n676 B.n39 163.367
R555 B.n672 B.n39 163.367
R556 B.n672 B.n44 163.367
R557 B.n668 B.n44 163.367
R558 B.n668 B.n46 163.367
R559 B.n664 B.n46 163.367
R560 B.n664 B.n51 163.367
R561 B.n660 B.n51 163.367
R562 B.n660 B.n53 163.367
R563 B.n656 B.n53 163.367
R564 B.n656 B.n58 163.367
R565 B.n510 B.n315 163.367
R566 B.n510 B.n354 163.367
R567 B.n506 B.n505 163.367
R568 B.n502 B.n501 163.367
R569 B.n498 B.n497 163.367
R570 B.n494 B.n493 163.367
R571 B.n490 B.n489 163.367
R572 B.n486 B.n485 163.367
R573 B.n482 B.n481 163.367
R574 B.n478 B.n477 163.367
R575 B.n474 B.n473 163.367
R576 B.n470 B.n469 163.367
R577 B.n466 B.n465 163.367
R578 B.n462 B.n461 163.367
R579 B.n458 B.n457 163.367
R580 B.n454 B.n453 163.367
R581 B.n450 B.n449 163.367
R582 B.n445 B.n444 163.367
R583 B.n441 B.n440 163.367
R584 B.n437 B.n436 163.367
R585 B.n433 B.n432 163.367
R586 B.n429 B.n428 163.367
R587 B.n424 B.n423 163.367
R588 B.n420 B.n419 163.367
R589 B.n416 B.n415 163.367
R590 B.n412 B.n411 163.367
R591 B.n408 B.n407 163.367
R592 B.n404 B.n403 163.367
R593 B.n400 B.n399 163.367
R594 B.n396 B.n395 163.367
R595 B.n392 B.n391 163.367
R596 B.n388 B.n387 163.367
R597 B.n384 B.n383 163.367
R598 B.n380 B.n379 163.367
R599 B.n376 B.n375 163.367
R600 B.n372 B.n371 163.367
R601 B.n368 B.n367 163.367
R602 B.n364 B.n363 163.367
R603 B.n360 B.n353 163.367
R604 B.n519 B.n311 163.367
R605 B.n519 B.n309 163.367
R606 B.n523 B.n309 163.367
R607 B.n523 B.n302 163.367
R608 B.n531 B.n302 163.367
R609 B.n531 B.n300 163.367
R610 B.n535 B.n300 163.367
R611 B.n535 B.n295 163.367
R612 B.n543 B.n295 163.367
R613 B.n543 B.n293 163.367
R614 B.n547 B.n293 163.367
R615 B.n547 B.n287 163.367
R616 B.n555 B.n287 163.367
R617 B.n555 B.n285 163.367
R618 B.n559 B.n285 163.367
R619 B.n559 B.n279 163.367
R620 B.n567 B.n279 163.367
R621 B.n567 B.n277 163.367
R622 B.n571 B.n277 163.367
R623 B.n571 B.n272 163.367
R624 B.n580 B.n272 163.367
R625 B.n580 B.n270 163.367
R626 B.n584 B.n270 163.367
R627 B.n584 B.n263 163.367
R628 B.n592 B.n263 163.367
R629 B.n592 B.n261 163.367
R630 B.n597 B.n261 163.367
R631 B.n597 B.n256 163.367
R632 B.n605 B.n256 163.367
R633 B.n606 B.n605 163.367
R634 B.n606 B.n5 163.367
R635 B.n6 B.n5 163.367
R636 B.n7 B.n6 163.367
R637 B.n611 B.n7 163.367
R638 B.n611 B.n12 163.367
R639 B.n13 B.n12 163.367
R640 B.n14 B.n13 163.367
R641 B.n616 B.n14 163.367
R642 B.n616 B.n19 163.367
R643 B.n20 B.n19 163.367
R644 B.n21 B.n20 163.367
R645 B.n621 B.n21 163.367
R646 B.n621 B.n26 163.367
R647 B.n27 B.n26 163.367
R648 B.n28 B.n27 163.367
R649 B.n626 B.n28 163.367
R650 B.n626 B.n33 163.367
R651 B.n34 B.n33 163.367
R652 B.n35 B.n34 163.367
R653 B.n631 B.n35 163.367
R654 B.n631 B.n40 163.367
R655 B.n41 B.n40 163.367
R656 B.n42 B.n41 163.367
R657 B.n636 B.n42 163.367
R658 B.n636 B.n47 163.367
R659 B.n48 B.n47 163.367
R660 B.n49 B.n48 163.367
R661 B.n641 B.n49 163.367
R662 B.n641 B.n54 163.367
R663 B.n55 B.n54 163.367
R664 B.n56 B.n55 163.367
R665 B.n99 B.n56 163.367
R666 B.n106 B.n60 163.367
R667 B.n110 B.n109 163.367
R668 B.n114 B.n113 163.367
R669 B.n118 B.n117 163.367
R670 B.n122 B.n121 163.367
R671 B.n126 B.n125 163.367
R672 B.n130 B.n129 163.367
R673 B.n134 B.n133 163.367
R674 B.n138 B.n137 163.367
R675 B.n142 B.n141 163.367
R676 B.n146 B.n145 163.367
R677 B.n150 B.n149 163.367
R678 B.n154 B.n153 163.367
R679 B.n158 B.n157 163.367
R680 B.n162 B.n161 163.367
R681 B.n166 B.n165 163.367
R682 B.n170 B.n169 163.367
R683 B.n174 B.n173 163.367
R684 B.n178 B.n177 163.367
R685 B.n182 B.n181 163.367
R686 B.n186 B.n185 163.367
R687 B.n190 B.n189 163.367
R688 B.n194 B.n193 163.367
R689 B.n198 B.n197 163.367
R690 B.n202 B.n201 163.367
R691 B.n206 B.n205 163.367
R692 B.n210 B.n209 163.367
R693 B.n214 B.n213 163.367
R694 B.n218 B.n217 163.367
R695 B.n222 B.n221 163.367
R696 B.n226 B.n225 163.367
R697 B.n230 B.n229 163.367
R698 B.n234 B.n233 163.367
R699 B.n238 B.n237 163.367
R700 B.n242 B.n241 163.367
R701 B.n246 B.n245 163.367
R702 B.n250 B.n249 163.367
R703 B.n252 B.n98 163.367
R704 B.n511 B.n312 88.5961
R705 B.n650 B.n57 88.5961
R706 B.n513 B.n512 71.676
R707 B.n354 B.n316 71.676
R708 B.n505 B.n317 71.676
R709 B.n501 B.n318 71.676
R710 B.n497 B.n319 71.676
R711 B.n493 B.n320 71.676
R712 B.n489 B.n321 71.676
R713 B.n485 B.n322 71.676
R714 B.n481 B.n323 71.676
R715 B.n477 B.n324 71.676
R716 B.n473 B.n325 71.676
R717 B.n469 B.n326 71.676
R718 B.n465 B.n327 71.676
R719 B.n461 B.n328 71.676
R720 B.n457 B.n329 71.676
R721 B.n453 B.n330 71.676
R722 B.n449 B.n331 71.676
R723 B.n444 B.n332 71.676
R724 B.n440 B.n333 71.676
R725 B.n436 B.n334 71.676
R726 B.n432 B.n335 71.676
R727 B.n428 B.n336 71.676
R728 B.n423 B.n337 71.676
R729 B.n419 B.n338 71.676
R730 B.n415 B.n339 71.676
R731 B.n411 B.n340 71.676
R732 B.n407 B.n341 71.676
R733 B.n403 B.n342 71.676
R734 B.n399 B.n343 71.676
R735 B.n395 B.n344 71.676
R736 B.n391 B.n345 71.676
R737 B.n387 B.n346 71.676
R738 B.n383 B.n347 71.676
R739 B.n379 B.n348 71.676
R740 B.n375 B.n349 71.676
R741 B.n371 B.n350 71.676
R742 B.n367 B.n351 71.676
R743 B.n363 B.n352 71.676
R744 B.n652 B.n651 71.676
R745 B.n106 B.n61 71.676
R746 B.n110 B.n62 71.676
R747 B.n114 B.n63 71.676
R748 B.n118 B.n64 71.676
R749 B.n122 B.n65 71.676
R750 B.n126 B.n66 71.676
R751 B.n130 B.n67 71.676
R752 B.n134 B.n68 71.676
R753 B.n138 B.n69 71.676
R754 B.n142 B.n70 71.676
R755 B.n146 B.n71 71.676
R756 B.n150 B.n72 71.676
R757 B.n154 B.n73 71.676
R758 B.n158 B.n74 71.676
R759 B.n162 B.n75 71.676
R760 B.n166 B.n76 71.676
R761 B.n170 B.n77 71.676
R762 B.n174 B.n78 71.676
R763 B.n178 B.n79 71.676
R764 B.n182 B.n80 71.676
R765 B.n186 B.n81 71.676
R766 B.n190 B.n82 71.676
R767 B.n194 B.n83 71.676
R768 B.n198 B.n84 71.676
R769 B.n202 B.n85 71.676
R770 B.n206 B.n86 71.676
R771 B.n210 B.n87 71.676
R772 B.n214 B.n88 71.676
R773 B.n218 B.n89 71.676
R774 B.n222 B.n90 71.676
R775 B.n226 B.n91 71.676
R776 B.n230 B.n92 71.676
R777 B.n234 B.n93 71.676
R778 B.n238 B.n94 71.676
R779 B.n242 B.n95 71.676
R780 B.n246 B.n96 71.676
R781 B.n250 B.n97 71.676
R782 B.n649 B.n98 71.676
R783 B.n649 B.n648 71.676
R784 B.n252 B.n97 71.676
R785 B.n249 B.n96 71.676
R786 B.n245 B.n95 71.676
R787 B.n241 B.n94 71.676
R788 B.n237 B.n93 71.676
R789 B.n233 B.n92 71.676
R790 B.n229 B.n91 71.676
R791 B.n225 B.n90 71.676
R792 B.n221 B.n89 71.676
R793 B.n217 B.n88 71.676
R794 B.n213 B.n87 71.676
R795 B.n209 B.n86 71.676
R796 B.n205 B.n85 71.676
R797 B.n201 B.n84 71.676
R798 B.n197 B.n83 71.676
R799 B.n193 B.n82 71.676
R800 B.n189 B.n81 71.676
R801 B.n185 B.n80 71.676
R802 B.n181 B.n79 71.676
R803 B.n177 B.n78 71.676
R804 B.n173 B.n77 71.676
R805 B.n169 B.n76 71.676
R806 B.n165 B.n75 71.676
R807 B.n161 B.n74 71.676
R808 B.n157 B.n73 71.676
R809 B.n153 B.n72 71.676
R810 B.n149 B.n71 71.676
R811 B.n145 B.n70 71.676
R812 B.n141 B.n69 71.676
R813 B.n137 B.n68 71.676
R814 B.n133 B.n67 71.676
R815 B.n129 B.n66 71.676
R816 B.n125 B.n65 71.676
R817 B.n121 B.n64 71.676
R818 B.n117 B.n63 71.676
R819 B.n113 B.n62 71.676
R820 B.n109 B.n61 71.676
R821 B.n651 B.n60 71.676
R822 B.n512 B.n315 71.676
R823 B.n506 B.n316 71.676
R824 B.n502 B.n317 71.676
R825 B.n498 B.n318 71.676
R826 B.n494 B.n319 71.676
R827 B.n490 B.n320 71.676
R828 B.n486 B.n321 71.676
R829 B.n482 B.n322 71.676
R830 B.n478 B.n323 71.676
R831 B.n474 B.n324 71.676
R832 B.n470 B.n325 71.676
R833 B.n466 B.n326 71.676
R834 B.n462 B.n327 71.676
R835 B.n458 B.n328 71.676
R836 B.n454 B.n329 71.676
R837 B.n450 B.n330 71.676
R838 B.n445 B.n331 71.676
R839 B.n441 B.n332 71.676
R840 B.n437 B.n333 71.676
R841 B.n433 B.n334 71.676
R842 B.n429 B.n335 71.676
R843 B.n424 B.n336 71.676
R844 B.n420 B.n337 71.676
R845 B.n416 B.n338 71.676
R846 B.n412 B.n339 71.676
R847 B.n408 B.n340 71.676
R848 B.n404 B.n341 71.676
R849 B.n400 B.n342 71.676
R850 B.n396 B.n343 71.676
R851 B.n392 B.n344 71.676
R852 B.n388 B.n345 71.676
R853 B.n384 B.n346 71.676
R854 B.n380 B.n347 71.676
R855 B.n376 B.n348 71.676
R856 B.n372 B.n349 71.676
R857 B.n368 B.n350 71.676
R858 B.n364 B.n351 71.676
R859 B.n360 B.n352 71.676
R860 B.n426 B.n358 59.5399
R861 B.n447 B.n356 59.5399
R862 B.n105 B.n104 59.5399
R863 B.n102 B.n101 59.5399
R864 B.n518 B.n312 50.6266
R865 B.n518 B.n308 50.6266
R866 B.n524 B.n308 50.6266
R867 B.n524 B.n303 50.6266
R868 B.n530 B.n303 50.6266
R869 B.n530 B.n304 50.6266
R870 B.n536 B.n296 50.6266
R871 B.n542 B.n296 50.6266
R872 B.n542 B.n292 50.6266
R873 B.n548 B.n292 50.6266
R874 B.n548 B.n288 50.6266
R875 B.n554 B.n288 50.6266
R876 B.n554 B.n284 50.6266
R877 B.n560 B.n284 50.6266
R878 B.n566 B.n280 50.6266
R879 B.n566 B.n276 50.6266
R880 B.n573 B.n276 50.6266
R881 B.n573 B.n572 50.6266
R882 B.n579 B.n269 50.6266
R883 B.n585 B.n269 50.6266
R884 B.n585 B.n264 50.6266
R885 B.n591 B.n264 50.6266
R886 B.n591 B.n265 50.6266
R887 B.n598 B.n257 50.6266
R888 B.n604 B.n257 50.6266
R889 B.n604 B.n4 50.6266
R890 B.n715 B.n4 50.6266
R891 B.n715 B.n714 50.6266
R892 B.n714 B.n713 50.6266
R893 B.n713 B.n8 50.6266
R894 B.n707 B.n8 50.6266
R895 B.n706 B.n705 50.6266
R896 B.n705 B.n15 50.6266
R897 B.n699 B.n15 50.6266
R898 B.n699 B.n698 50.6266
R899 B.n698 B.n697 50.6266
R900 B.n691 B.n25 50.6266
R901 B.n691 B.n690 50.6266
R902 B.n690 B.n689 50.6266
R903 B.n689 B.n29 50.6266
R904 B.n683 B.n682 50.6266
R905 B.n682 B.n681 50.6266
R906 B.n681 B.n36 50.6266
R907 B.n675 B.n36 50.6266
R908 B.n675 B.n674 50.6266
R909 B.n674 B.n673 50.6266
R910 B.n673 B.n43 50.6266
R911 B.n667 B.n43 50.6266
R912 B.n666 B.n665 50.6266
R913 B.n665 B.n50 50.6266
R914 B.n659 B.n50 50.6266
R915 B.n659 B.n658 50.6266
R916 B.n658 B.n657 50.6266
R917 B.n657 B.n57 50.6266
R918 B.t4 B.n280 43.9261
R919 B.t3 B.n29 43.9261
R920 B.n572 B.t19 42.437
R921 B.n25 B.t0 42.437
R922 B.n536 B.t10 39.459
R923 B.n667 B.t6 39.459
R924 B.n358 B.n357 37.6247
R925 B.n356 B.n355 37.6247
R926 B.n104 B.n103 37.6247
R927 B.n101 B.n100 37.6247
R928 B.n654 B.n653 32.3127
R929 B.n647 B.n646 32.3127
R930 B.n359 B.n310 32.3127
R931 B.n515 B.n514 32.3127
R932 B.n265 B.t2 27.547
R933 B.t1 B.n706 27.547
R934 B.n598 B.t2 23.08
R935 B.n707 B.t1 23.08
R936 B B.n717 18.0485
R937 B.n304 B.t10 11.168
R938 B.t6 B.n666 11.168
R939 B.n653 B.n59 10.6151
R940 B.n107 B.n59 10.6151
R941 B.n108 B.n107 10.6151
R942 B.n111 B.n108 10.6151
R943 B.n112 B.n111 10.6151
R944 B.n115 B.n112 10.6151
R945 B.n116 B.n115 10.6151
R946 B.n119 B.n116 10.6151
R947 B.n120 B.n119 10.6151
R948 B.n123 B.n120 10.6151
R949 B.n124 B.n123 10.6151
R950 B.n127 B.n124 10.6151
R951 B.n128 B.n127 10.6151
R952 B.n131 B.n128 10.6151
R953 B.n132 B.n131 10.6151
R954 B.n135 B.n132 10.6151
R955 B.n136 B.n135 10.6151
R956 B.n139 B.n136 10.6151
R957 B.n140 B.n139 10.6151
R958 B.n143 B.n140 10.6151
R959 B.n144 B.n143 10.6151
R960 B.n147 B.n144 10.6151
R961 B.n148 B.n147 10.6151
R962 B.n151 B.n148 10.6151
R963 B.n152 B.n151 10.6151
R964 B.n155 B.n152 10.6151
R965 B.n156 B.n155 10.6151
R966 B.n159 B.n156 10.6151
R967 B.n160 B.n159 10.6151
R968 B.n163 B.n160 10.6151
R969 B.n164 B.n163 10.6151
R970 B.n167 B.n164 10.6151
R971 B.n168 B.n167 10.6151
R972 B.n172 B.n171 10.6151
R973 B.n175 B.n172 10.6151
R974 B.n176 B.n175 10.6151
R975 B.n179 B.n176 10.6151
R976 B.n180 B.n179 10.6151
R977 B.n183 B.n180 10.6151
R978 B.n184 B.n183 10.6151
R979 B.n187 B.n184 10.6151
R980 B.n188 B.n187 10.6151
R981 B.n192 B.n191 10.6151
R982 B.n195 B.n192 10.6151
R983 B.n196 B.n195 10.6151
R984 B.n199 B.n196 10.6151
R985 B.n200 B.n199 10.6151
R986 B.n203 B.n200 10.6151
R987 B.n204 B.n203 10.6151
R988 B.n207 B.n204 10.6151
R989 B.n208 B.n207 10.6151
R990 B.n211 B.n208 10.6151
R991 B.n212 B.n211 10.6151
R992 B.n215 B.n212 10.6151
R993 B.n216 B.n215 10.6151
R994 B.n219 B.n216 10.6151
R995 B.n220 B.n219 10.6151
R996 B.n223 B.n220 10.6151
R997 B.n224 B.n223 10.6151
R998 B.n227 B.n224 10.6151
R999 B.n228 B.n227 10.6151
R1000 B.n231 B.n228 10.6151
R1001 B.n232 B.n231 10.6151
R1002 B.n235 B.n232 10.6151
R1003 B.n236 B.n235 10.6151
R1004 B.n239 B.n236 10.6151
R1005 B.n240 B.n239 10.6151
R1006 B.n243 B.n240 10.6151
R1007 B.n244 B.n243 10.6151
R1008 B.n247 B.n244 10.6151
R1009 B.n248 B.n247 10.6151
R1010 B.n251 B.n248 10.6151
R1011 B.n253 B.n251 10.6151
R1012 B.n254 B.n253 10.6151
R1013 B.n647 B.n254 10.6151
R1014 B.n520 B.n310 10.6151
R1015 B.n521 B.n520 10.6151
R1016 B.n522 B.n521 10.6151
R1017 B.n522 B.n301 10.6151
R1018 B.n532 B.n301 10.6151
R1019 B.n533 B.n532 10.6151
R1020 B.n534 B.n533 10.6151
R1021 B.n534 B.n294 10.6151
R1022 B.n544 B.n294 10.6151
R1023 B.n545 B.n544 10.6151
R1024 B.n546 B.n545 10.6151
R1025 B.n546 B.n286 10.6151
R1026 B.n556 B.n286 10.6151
R1027 B.n557 B.n556 10.6151
R1028 B.n558 B.n557 10.6151
R1029 B.n558 B.n278 10.6151
R1030 B.n568 B.n278 10.6151
R1031 B.n569 B.n568 10.6151
R1032 B.n570 B.n569 10.6151
R1033 B.n570 B.n271 10.6151
R1034 B.n581 B.n271 10.6151
R1035 B.n582 B.n581 10.6151
R1036 B.n583 B.n582 10.6151
R1037 B.n583 B.n262 10.6151
R1038 B.n593 B.n262 10.6151
R1039 B.n594 B.n593 10.6151
R1040 B.n596 B.n594 10.6151
R1041 B.n596 B.n595 10.6151
R1042 B.n595 B.n255 10.6151
R1043 B.n607 B.n255 10.6151
R1044 B.n608 B.n607 10.6151
R1045 B.n609 B.n608 10.6151
R1046 B.n610 B.n609 10.6151
R1047 B.n612 B.n610 10.6151
R1048 B.n613 B.n612 10.6151
R1049 B.n614 B.n613 10.6151
R1050 B.n615 B.n614 10.6151
R1051 B.n617 B.n615 10.6151
R1052 B.n618 B.n617 10.6151
R1053 B.n619 B.n618 10.6151
R1054 B.n620 B.n619 10.6151
R1055 B.n622 B.n620 10.6151
R1056 B.n623 B.n622 10.6151
R1057 B.n624 B.n623 10.6151
R1058 B.n625 B.n624 10.6151
R1059 B.n627 B.n625 10.6151
R1060 B.n628 B.n627 10.6151
R1061 B.n629 B.n628 10.6151
R1062 B.n630 B.n629 10.6151
R1063 B.n632 B.n630 10.6151
R1064 B.n633 B.n632 10.6151
R1065 B.n634 B.n633 10.6151
R1066 B.n635 B.n634 10.6151
R1067 B.n637 B.n635 10.6151
R1068 B.n638 B.n637 10.6151
R1069 B.n639 B.n638 10.6151
R1070 B.n640 B.n639 10.6151
R1071 B.n642 B.n640 10.6151
R1072 B.n643 B.n642 10.6151
R1073 B.n644 B.n643 10.6151
R1074 B.n645 B.n644 10.6151
R1075 B.n646 B.n645 10.6151
R1076 B.n514 B.n314 10.6151
R1077 B.n509 B.n314 10.6151
R1078 B.n509 B.n508 10.6151
R1079 B.n508 B.n507 10.6151
R1080 B.n507 B.n504 10.6151
R1081 B.n504 B.n503 10.6151
R1082 B.n503 B.n500 10.6151
R1083 B.n500 B.n499 10.6151
R1084 B.n499 B.n496 10.6151
R1085 B.n496 B.n495 10.6151
R1086 B.n495 B.n492 10.6151
R1087 B.n492 B.n491 10.6151
R1088 B.n491 B.n488 10.6151
R1089 B.n488 B.n487 10.6151
R1090 B.n487 B.n484 10.6151
R1091 B.n484 B.n483 10.6151
R1092 B.n483 B.n480 10.6151
R1093 B.n480 B.n479 10.6151
R1094 B.n479 B.n476 10.6151
R1095 B.n476 B.n475 10.6151
R1096 B.n475 B.n472 10.6151
R1097 B.n472 B.n471 10.6151
R1098 B.n471 B.n468 10.6151
R1099 B.n468 B.n467 10.6151
R1100 B.n467 B.n464 10.6151
R1101 B.n464 B.n463 10.6151
R1102 B.n463 B.n460 10.6151
R1103 B.n460 B.n459 10.6151
R1104 B.n459 B.n456 10.6151
R1105 B.n456 B.n455 10.6151
R1106 B.n455 B.n452 10.6151
R1107 B.n452 B.n451 10.6151
R1108 B.n451 B.n448 10.6151
R1109 B.n446 B.n443 10.6151
R1110 B.n443 B.n442 10.6151
R1111 B.n442 B.n439 10.6151
R1112 B.n439 B.n438 10.6151
R1113 B.n438 B.n435 10.6151
R1114 B.n435 B.n434 10.6151
R1115 B.n434 B.n431 10.6151
R1116 B.n431 B.n430 10.6151
R1117 B.n430 B.n427 10.6151
R1118 B.n425 B.n422 10.6151
R1119 B.n422 B.n421 10.6151
R1120 B.n421 B.n418 10.6151
R1121 B.n418 B.n417 10.6151
R1122 B.n417 B.n414 10.6151
R1123 B.n414 B.n413 10.6151
R1124 B.n413 B.n410 10.6151
R1125 B.n410 B.n409 10.6151
R1126 B.n409 B.n406 10.6151
R1127 B.n406 B.n405 10.6151
R1128 B.n405 B.n402 10.6151
R1129 B.n402 B.n401 10.6151
R1130 B.n401 B.n398 10.6151
R1131 B.n398 B.n397 10.6151
R1132 B.n397 B.n394 10.6151
R1133 B.n394 B.n393 10.6151
R1134 B.n393 B.n390 10.6151
R1135 B.n390 B.n389 10.6151
R1136 B.n389 B.n386 10.6151
R1137 B.n386 B.n385 10.6151
R1138 B.n385 B.n382 10.6151
R1139 B.n382 B.n381 10.6151
R1140 B.n381 B.n378 10.6151
R1141 B.n378 B.n377 10.6151
R1142 B.n377 B.n374 10.6151
R1143 B.n374 B.n373 10.6151
R1144 B.n373 B.n370 10.6151
R1145 B.n370 B.n369 10.6151
R1146 B.n369 B.n366 10.6151
R1147 B.n366 B.n365 10.6151
R1148 B.n365 B.n362 10.6151
R1149 B.n362 B.n361 10.6151
R1150 B.n361 B.n359 10.6151
R1151 B.n516 B.n515 10.6151
R1152 B.n516 B.n306 10.6151
R1153 B.n526 B.n306 10.6151
R1154 B.n527 B.n526 10.6151
R1155 B.n528 B.n527 10.6151
R1156 B.n528 B.n298 10.6151
R1157 B.n538 B.n298 10.6151
R1158 B.n539 B.n538 10.6151
R1159 B.n540 B.n539 10.6151
R1160 B.n540 B.n290 10.6151
R1161 B.n550 B.n290 10.6151
R1162 B.n551 B.n550 10.6151
R1163 B.n552 B.n551 10.6151
R1164 B.n552 B.n282 10.6151
R1165 B.n562 B.n282 10.6151
R1166 B.n563 B.n562 10.6151
R1167 B.n564 B.n563 10.6151
R1168 B.n564 B.n274 10.6151
R1169 B.n575 B.n274 10.6151
R1170 B.n576 B.n575 10.6151
R1171 B.n577 B.n576 10.6151
R1172 B.n577 B.n267 10.6151
R1173 B.n587 B.n267 10.6151
R1174 B.n588 B.n587 10.6151
R1175 B.n589 B.n588 10.6151
R1176 B.n589 B.n259 10.6151
R1177 B.n600 B.n259 10.6151
R1178 B.n601 B.n600 10.6151
R1179 B.n602 B.n601 10.6151
R1180 B.n602 B.n0 10.6151
R1181 B.n711 B.n1 10.6151
R1182 B.n711 B.n710 10.6151
R1183 B.n710 B.n709 10.6151
R1184 B.n709 B.n10 10.6151
R1185 B.n703 B.n10 10.6151
R1186 B.n703 B.n702 10.6151
R1187 B.n702 B.n701 10.6151
R1188 B.n701 B.n17 10.6151
R1189 B.n695 B.n17 10.6151
R1190 B.n695 B.n694 10.6151
R1191 B.n694 B.n693 10.6151
R1192 B.n693 B.n23 10.6151
R1193 B.n687 B.n23 10.6151
R1194 B.n687 B.n686 10.6151
R1195 B.n686 B.n685 10.6151
R1196 B.n685 B.n31 10.6151
R1197 B.n679 B.n31 10.6151
R1198 B.n679 B.n678 10.6151
R1199 B.n678 B.n677 10.6151
R1200 B.n677 B.n38 10.6151
R1201 B.n671 B.n38 10.6151
R1202 B.n671 B.n670 10.6151
R1203 B.n670 B.n669 10.6151
R1204 B.n669 B.n45 10.6151
R1205 B.n663 B.n45 10.6151
R1206 B.n663 B.n662 10.6151
R1207 B.n662 B.n661 10.6151
R1208 B.n661 B.n52 10.6151
R1209 B.n655 B.n52 10.6151
R1210 B.n655 B.n654 10.6151
R1211 B.n168 B.n105 9.36635
R1212 B.n191 B.n102 9.36635
R1213 B.n448 B.n447 9.36635
R1214 B.n426 B.n425 9.36635
R1215 B.n579 B.t19 8.19001
R1216 B.n697 B.t0 8.19001
R1217 B.n560 B.t4 6.70101
R1218 B.n683 B.t3 6.70101
R1219 B.n717 B.n0 2.81026
R1220 B.n717 B.n1 2.81026
R1221 B.n171 B.n105 1.24928
R1222 B.n188 B.n102 1.24928
R1223 B.n447 B.n446 1.24928
R1224 B.n427 B.n426 1.24928
R1225 VN.n11 VN.n10 176.548
R1226 VN.n23 VN.n22 176.548
R1227 VN.n2 VN.t2 175.653
R1228 VN.n14 VN.t4 175.653
R1229 VN.n21 VN.n12 161.3
R1230 VN.n20 VN.n19 161.3
R1231 VN.n18 VN.n13 161.3
R1232 VN.n17 VN.n16 161.3
R1233 VN.n9 VN.n0 161.3
R1234 VN.n8 VN.n7 161.3
R1235 VN.n6 VN.n1 161.3
R1236 VN.n5 VN.n4 161.3
R1237 VN.n3 VN.t5 142.206
R1238 VN.n10 VN.t3 142.206
R1239 VN.n15 VN.t1 142.206
R1240 VN.n22 VN.t0 142.206
R1241 VN.n8 VN.n1 56.5617
R1242 VN.n20 VN.n13 56.5617
R1243 VN.n3 VN.n2 54.2185
R1244 VN.n15 VN.n14 54.2185
R1245 VN VN.n23 43.2221
R1246 VN.n4 VN.n1 24.5923
R1247 VN.n9 VN.n8 24.5923
R1248 VN.n16 VN.n13 24.5923
R1249 VN.n21 VN.n20 24.5923
R1250 VN.n17 VN.n14 17.8292
R1251 VN.n5 VN.n2 17.8292
R1252 VN.n4 VN.n3 12.2964
R1253 VN.n16 VN.n15 12.2964
R1254 VN.n10 VN.n9 9.3454
R1255 VN.n22 VN.n21 9.3454
R1256 VN.n23 VN.n12 0.189894
R1257 VN.n19 VN.n12 0.189894
R1258 VN.n19 VN.n18 0.189894
R1259 VN.n18 VN.n17 0.189894
R1260 VN.n6 VN.n5 0.189894
R1261 VN.n7 VN.n6 0.189894
R1262 VN.n7 VN.n0 0.189894
R1263 VN.n11 VN.n0 0.189894
R1264 VN VN.n11 0.0516364
R1265 VTAIL.n210 VTAIL.n164 289.615
R1266 VTAIL.n48 VTAIL.n2 289.615
R1267 VTAIL.n158 VTAIL.n112 289.615
R1268 VTAIL.n104 VTAIL.n58 289.615
R1269 VTAIL.n180 VTAIL.n179 185
R1270 VTAIL.n185 VTAIL.n184 185
R1271 VTAIL.n187 VTAIL.n186 185
R1272 VTAIL.n176 VTAIL.n175 185
R1273 VTAIL.n193 VTAIL.n192 185
R1274 VTAIL.n195 VTAIL.n194 185
R1275 VTAIL.n172 VTAIL.n171 185
R1276 VTAIL.n201 VTAIL.n200 185
R1277 VTAIL.n203 VTAIL.n202 185
R1278 VTAIL.n168 VTAIL.n167 185
R1279 VTAIL.n209 VTAIL.n208 185
R1280 VTAIL.n211 VTAIL.n210 185
R1281 VTAIL.n18 VTAIL.n17 185
R1282 VTAIL.n23 VTAIL.n22 185
R1283 VTAIL.n25 VTAIL.n24 185
R1284 VTAIL.n14 VTAIL.n13 185
R1285 VTAIL.n31 VTAIL.n30 185
R1286 VTAIL.n33 VTAIL.n32 185
R1287 VTAIL.n10 VTAIL.n9 185
R1288 VTAIL.n39 VTAIL.n38 185
R1289 VTAIL.n41 VTAIL.n40 185
R1290 VTAIL.n6 VTAIL.n5 185
R1291 VTAIL.n47 VTAIL.n46 185
R1292 VTAIL.n49 VTAIL.n48 185
R1293 VTAIL.n159 VTAIL.n158 185
R1294 VTAIL.n157 VTAIL.n156 185
R1295 VTAIL.n116 VTAIL.n115 185
R1296 VTAIL.n151 VTAIL.n150 185
R1297 VTAIL.n149 VTAIL.n148 185
R1298 VTAIL.n120 VTAIL.n119 185
R1299 VTAIL.n143 VTAIL.n142 185
R1300 VTAIL.n141 VTAIL.n140 185
R1301 VTAIL.n124 VTAIL.n123 185
R1302 VTAIL.n135 VTAIL.n134 185
R1303 VTAIL.n133 VTAIL.n132 185
R1304 VTAIL.n128 VTAIL.n127 185
R1305 VTAIL.n105 VTAIL.n104 185
R1306 VTAIL.n103 VTAIL.n102 185
R1307 VTAIL.n62 VTAIL.n61 185
R1308 VTAIL.n97 VTAIL.n96 185
R1309 VTAIL.n95 VTAIL.n94 185
R1310 VTAIL.n66 VTAIL.n65 185
R1311 VTAIL.n89 VTAIL.n88 185
R1312 VTAIL.n87 VTAIL.n86 185
R1313 VTAIL.n70 VTAIL.n69 185
R1314 VTAIL.n81 VTAIL.n80 185
R1315 VTAIL.n79 VTAIL.n78 185
R1316 VTAIL.n74 VTAIL.n73 185
R1317 VTAIL.n129 VTAIL.t1 147.659
R1318 VTAIL.n181 VTAIL.t11 147.659
R1319 VTAIL.n19 VTAIL.t0 147.659
R1320 VTAIL.n75 VTAIL.t6 147.659
R1321 VTAIL.n185 VTAIL.n179 104.615
R1322 VTAIL.n186 VTAIL.n185 104.615
R1323 VTAIL.n186 VTAIL.n175 104.615
R1324 VTAIL.n193 VTAIL.n175 104.615
R1325 VTAIL.n194 VTAIL.n193 104.615
R1326 VTAIL.n194 VTAIL.n171 104.615
R1327 VTAIL.n201 VTAIL.n171 104.615
R1328 VTAIL.n202 VTAIL.n201 104.615
R1329 VTAIL.n202 VTAIL.n167 104.615
R1330 VTAIL.n209 VTAIL.n167 104.615
R1331 VTAIL.n210 VTAIL.n209 104.615
R1332 VTAIL.n23 VTAIL.n17 104.615
R1333 VTAIL.n24 VTAIL.n23 104.615
R1334 VTAIL.n24 VTAIL.n13 104.615
R1335 VTAIL.n31 VTAIL.n13 104.615
R1336 VTAIL.n32 VTAIL.n31 104.615
R1337 VTAIL.n32 VTAIL.n9 104.615
R1338 VTAIL.n39 VTAIL.n9 104.615
R1339 VTAIL.n40 VTAIL.n39 104.615
R1340 VTAIL.n40 VTAIL.n5 104.615
R1341 VTAIL.n47 VTAIL.n5 104.615
R1342 VTAIL.n48 VTAIL.n47 104.615
R1343 VTAIL.n158 VTAIL.n157 104.615
R1344 VTAIL.n157 VTAIL.n115 104.615
R1345 VTAIL.n150 VTAIL.n115 104.615
R1346 VTAIL.n150 VTAIL.n149 104.615
R1347 VTAIL.n149 VTAIL.n119 104.615
R1348 VTAIL.n142 VTAIL.n119 104.615
R1349 VTAIL.n142 VTAIL.n141 104.615
R1350 VTAIL.n141 VTAIL.n123 104.615
R1351 VTAIL.n134 VTAIL.n123 104.615
R1352 VTAIL.n134 VTAIL.n133 104.615
R1353 VTAIL.n133 VTAIL.n127 104.615
R1354 VTAIL.n104 VTAIL.n103 104.615
R1355 VTAIL.n103 VTAIL.n61 104.615
R1356 VTAIL.n96 VTAIL.n61 104.615
R1357 VTAIL.n96 VTAIL.n95 104.615
R1358 VTAIL.n95 VTAIL.n65 104.615
R1359 VTAIL.n88 VTAIL.n65 104.615
R1360 VTAIL.n88 VTAIL.n87 104.615
R1361 VTAIL.n87 VTAIL.n69 104.615
R1362 VTAIL.n80 VTAIL.n69 104.615
R1363 VTAIL.n80 VTAIL.n79 104.615
R1364 VTAIL.n79 VTAIL.n73 104.615
R1365 VTAIL.t11 VTAIL.n179 52.3082
R1366 VTAIL.t0 VTAIL.n17 52.3082
R1367 VTAIL.t1 VTAIL.n127 52.3082
R1368 VTAIL.t6 VTAIL.n73 52.3082
R1369 VTAIL.n1 VTAIL.n0 44.856
R1370 VTAIL.n55 VTAIL.n54 44.856
R1371 VTAIL.n111 VTAIL.n110 44.856
R1372 VTAIL.n57 VTAIL.n56 44.856
R1373 VTAIL.n215 VTAIL.n214 30.246
R1374 VTAIL.n53 VTAIL.n52 30.246
R1375 VTAIL.n163 VTAIL.n162 30.246
R1376 VTAIL.n109 VTAIL.n108 30.246
R1377 VTAIL.n57 VTAIL.n55 23.9014
R1378 VTAIL.n215 VTAIL.n163 22.2289
R1379 VTAIL.n181 VTAIL.n180 15.6677
R1380 VTAIL.n19 VTAIL.n18 15.6677
R1381 VTAIL.n129 VTAIL.n128 15.6677
R1382 VTAIL.n75 VTAIL.n74 15.6677
R1383 VTAIL.n184 VTAIL.n183 12.8005
R1384 VTAIL.n22 VTAIL.n21 12.8005
R1385 VTAIL.n132 VTAIL.n131 12.8005
R1386 VTAIL.n78 VTAIL.n77 12.8005
R1387 VTAIL.n187 VTAIL.n178 12.0247
R1388 VTAIL.n25 VTAIL.n16 12.0247
R1389 VTAIL.n135 VTAIL.n126 12.0247
R1390 VTAIL.n81 VTAIL.n72 12.0247
R1391 VTAIL.n188 VTAIL.n176 11.249
R1392 VTAIL.n26 VTAIL.n14 11.249
R1393 VTAIL.n136 VTAIL.n124 11.249
R1394 VTAIL.n82 VTAIL.n70 11.249
R1395 VTAIL.n192 VTAIL.n191 10.4732
R1396 VTAIL.n30 VTAIL.n29 10.4732
R1397 VTAIL.n140 VTAIL.n139 10.4732
R1398 VTAIL.n86 VTAIL.n85 10.4732
R1399 VTAIL.n195 VTAIL.n174 9.69747
R1400 VTAIL.n214 VTAIL.n164 9.69747
R1401 VTAIL.n33 VTAIL.n12 9.69747
R1402 VTAIL.n52 VTAIL.n2 9.69747
R1403 VTAIL.n162 VTAIL.n112 9.69747
R1404 VTAIL.n143 VTAIL.n122 9.69747
R1405 VTAIL.n108 VTAIL.n58 9.69747
R1406 VTAIL.n89 VTAIL.n68 9.69747
R1407 VTAIL.n214 VTAIL.n213 9.45567
R1408 VTAIL.n52 VTAIL.n51 9.45567
R1409 VTAIL.n162 VTAIL.n161 9.45567
R1410 VTAIL.n108 VTAIL.n107 9.45567
R1411 VTAIL.n205 VTAIL.n204 9.3005
R1412 VTAIL.n207 VTAIL.n206 9.3005
R1413 VTAIL.n166 VTAIL.n165 9.3005
R1414 VTAIL.n213 VTAIL.n212 9.3005
R1415 VTAIL.n199 VTAIL.n198 9.3005
R1416 VTAIL.n197 VTAIL.n196 9.3005
R1417 VTAIL.n174 VTAIL.n173 9.3005
R1418 VTAIL.n191 VTAIL.n190 9.3005
R1419 VTAIL.n189 VTAIL.n188 9.3005
R1420 VTAIL.n178 VTAIL.n177 9.3005
R1421 VTAIL.n183 VTAIL.n182 9.3005
R1422 VTAIL.n170 VTAIL.n169 9.3005
R1423 VTAIL.n43 VTAIL.n42 9.3005
R1424 VTAIL.n45 VTAIL.n44 9.3005
R1425 VTAIL.n4 VTAIL.n3 9.3005
R1426 VTAIL.n51 VTAIL.n50 9.3005
R1427 VTAIL.n37 VTAIL.n36 9.3005
R1428 VTAIL.n35 VTAIL.n34 9.3005
R1429 VTAIL.n12 VTAIL.n11 9.3005
R1430 VTAIL.n29 VTAIL.n28 9.3005
R1431 VTAIL.n27 VTAIL.n26 9.3005
R1432 VTAIL.n16 VTAIL.n15 9.3005
R1433 VTAIL.n21 VTAIL.n20 9.3005
R1434 VTAIL.n8 VTAIL.n7 9.3005
R1435 VTAIL.n114 VTAIL.n113 9.3005
R1436 VTAIL.n155 VTAIL.n154 9.3005
R1437 VTAIL.n153 VTAIL.n152 9.3005
R1438 VTAIL.n118 VTAIL.n117 9.3005
R1439 VTAIL.n147 VTAIL.n146 9.3005
R1440 VTAIL.n145 VTAIL.n144 9.3005
R1441 VTAIL.n122 VTAIL.n121 9.3005
R1442 VTAIL.n139 VTAIL.n138 9.3005
R1443 VTAIL.n137 VTAIL.n136 9.3005
R1444 VTAIL.n126 VTAIL.n125 9.3005
R1445 VTAIL.n131 VTAIL.n130 9.3005
R1446 VTAIL.n161 VTAIL.n160 9.3005
R1447 VTAIL.n101 VTAIL.n100 9.3005
R1448 VTAIL.n60 VTAIL.n59 9.3005
R1449 VTAIL.n107 VTAIL.n106 9.3005
R1450 VTAIL.n99 VTAIL.n98 9.3005
R1451 VTAIL.n64 VTAIL.n63 9.3005
R1452 VTAIL.n93 VTAIL.n92 9.3005
R1453 VTAIL.n91 VTAIL.n90 9.3005
R1454 VTAIL.n68 VTAIL.n67 9.3005
R1455 VTAIL.n85 VTAIL.n84 9.3005
R1456 VTAIL.n83 VTAIL.n82 9.3005
R1457 VTAIL.n72 VTAIL.n71 9.3005
R1458 VTAIL.n77 VTAIL.n76 9.3005
R1459 VTAIL.n196 VTAIL.n172 8.92171
R1460 VTAIL.n212 VTAIL.n211 8.92171
R1461 VTAIL.n34 VTAIL.n10 8.92171
R1462 VTAIL.n50 VTAIL.n49 8.92171
R1463 VTAIL.n160 VTAIL.n159 8.92171
R1464 VTAIL.n144 VTAIL.n120 8.92171
R1465 VTAIL.n106 VTAIL.n105 8.92171
R1466 VTAIL.n90 VTAIL.n66 8.92171
R1467 VTAIL.n200 VTAIL.n199 8.14595
R1468 VTAIL.n208 VTAIL.n166 8.14595
R1469 VTAIL.n38 VTAIL.n37 8.14595
R1470 VTAIL.n46 VTAIL.n4 8.14595
R1471 VTAIL.n156 VTAIL.n114 8.14595
R1472 VTAIL.n148 VTAIL.n147 8.14595
R1473 VTAIL.n102 VTAIL.n60 8.14595
R1474 VTAIL.n94 VTAIL.n93 8.14595
R1475 VTAIL.n203 VTAIL.n170 7.3702
R1476 VTAIL.n207 VTAIL.n168 7.3702
R1477 VTAIL.n41 VTAIL.n8 7.3702
R1478 VTAIL.n45 VTAIL.n6 7.3702
R1479 VTAIL.n155 VTAIL.n116 7.3702
R1480 VTAIL.n151 VTAIL.n118 7.3702
R1481 VTAIL.n101 VTAIL.n62 7.3702
R1482 VTAIL.n97 VTAIL.n64 7.3702
R1483 VTAIL.n204 VTAIL.n203 6.59444
R1484 VTAIL.n204 VTAIL.n168 6.59444
R1485 VTAIL.n42 VTAIL.n41 6.59444
R1486 VTAIL.n42 VTAIL.n6 6.59444
R1487 VTAIL.n152 VTAIL.n116 6.59444
R1488 VTAIL.n152 VTAIL.n151 6.59444
R1489 VTAIL.n98 VTAIL.n62 6.59444
R1490 VTAIL.n98 VTAIL.n97 6.59444
R1491 VTAIL.n200 VTAIL.n170 5.81868
R1492 VTAIL.n208 VTAIL.n207 5.81868
R1493 VTAIL.n38 VTAIL.n8 5.81868
R1494 VTAIL.n46 VTAIL.n45 5.81868
R1495 VTAIL.n156 VTAIL.n155 5.81868
R1496 VTAIL.n148 VTAIL.n118 5.81868
R1497 VTAIL.n102 VTAIL.n101 5.81868
R1498 VTAIL.n94 VTAIL.n64 5.81868
R1499 VTAIL.n199 VTAIL.n172 5.04292
R1500 VTAIL.n211 VTAIL.n166 5.04292
R1501 VTAIL.n37 VTAIL.n10 5.04292
R1502 VTAIL.n49 VTAIL.n4 5.04292
R1503 VTAIL.n159 VTAIL.n114 5.04292
R1504 VTAIL.n147 VTAIL.n120 5.04292
R1505 VTAIL.n105 VTAIL.n60 5.04292
R1506 VTAIL.n93 VTAIL.n66 5.04292
R1507 VTAIL.n182 VTAIL.n181 4.38563
R1508 VTAIL.n20 VTAIL.n19 4.38563
R1509 VTAIL.n130 VTAIL.n129 4.38563
R1510 VTAIL.n76 VTAIL.n75 4.38563
R1511 VTAIL.n196 VTAIL.n195 4.26717
R1512 VTAIL.n212 VTAIL.n164 4.26717
R1513 VTAIL.n34 VTAIL.n33 4.26717
R1514 VTAIL.n50 VTAIL.n2 4.26717
R1515 VTAIL.n160 VTAIL.n112 4.26717
R1516 VTAIL.n144 VTAIL.n143 4.26717
R1517 VTAIL.n106 VTAIL.n58 4.26717
R1518 VTAIL.n90 VTAIL.n89 4.26717
R1519 VTAIL.n192 VTAIL.n174 3.49141
R1520 VTAIL.n30 VTAIL.n12 3.49141
R1521 VTAIL.n140 VTAIL.n122 3.49141
R1522 VTAIL.n86 VTAIL.n68 3.49141
R1523 VTAIL.n191 VTAIL.n176 2.71565
R1524 VTAIL.n29 VTAIL.n14 2.71565
R1525 VTAIL.n139 VTAIL.n124 2.71565
R1526 VTAIL.n85 VTAIL.n70 2.71565
R1527 VTAIL.n0 VTAIL.t10 2.08471
R1528 VTAIL.n0 VTAIL.t7 2.08471
R1529 VTAIL.n54 VTAIL.t3 2.08471
R1530 VTAIL.n54 VTAIL.t4 2.08471
R1531 VTAIL.n110 VTAIL.t5 2.08471
R1532 VTAIL.n110 VTAIL.t2 2.08471
R1533 VTAIL.n56 VTAIL.t9 2.08471
R1534 VTAIL.n56 VTAIL.t8 2.08471
R1535 VTAIL.n188 VTAIL.n187 1.93989
R1536 VTAIL.n26 VTAIL.n25 1.93989
R1537 VTAIL.n136 VTAIL.n135 1.93989
R1538 VTAIL.n82 VTAIL.n81 1.93989
R1539 VTAIL.n109 VTAIL.n57 1.67291
R1540 VTAIL.n163 VTAIL.n111 1.67291
R1541 VTAIL.n55 VTAIL.n53 1.67291
R1542 VTAIL.n111 VTAIL.n109 1.30653
R1543 VTAIL.n53 VTAIL.n1 1.30653
R1544 VTAIL VTAIL.n215 1.19662
R1545 VTAIL.n184 VTAIL.n178 1.16414
R1546 VTAIL.n22 VTAIL.n16 1.16414
R1547 VTAIL.n132 VTAIL.n126 1.16414
R1548 VTAIL.n78 VTAIL.n72 1.16414
R1549 VTAIL VTAIL.n1 0.476793
R1550 VTAIL.n183 VTAIL.n180 0.388379
R1551 VTAIL.n21 VTAIL.n18 0.388379
R1552 VTAIL.n131 VTAIL.n128 0.388379
R1553 VTAIL.n77 VTAIL.n74 0.388379
R1554 VTAIL.n182 VTAIL.n177 0.155672
R1555 VTAIL.n189 VTAIL.n177 0.155672
R1556 VTAIL.n190 VTAIL.n189 0.155672
R1557 VTAIL.n190 VTAIL.n173 0.155672
R1558 VTAIL.n197 VTAIL.n173 0.155672
R1559 VTAIL.n198 VTAIL.n197 0.155672
R1560 VTAIL.n198 VTAIL.n169 0.155672
R1561 VTAIL.n205 VTAIL.n169 0.155672
R1562 VTAIL.n206 VTAIL.n205 0.155672
R1563 VTAIL.n206 VTAIL.n165 0.155672
R1564 VTAIL.n213 VTAIL.n165 0.155672
R1565 VTAIL.n20 VTAIL.n15 0.155672
R1566 VTAIL.n27 VTAIL.n15 0.155672
R1567 VTAIL.n28 VTAIL.n27 0.155672
R1568 VTAIL.n28 VTAIL.n11 0.155672
R1569 VTAIL.n35 VTAIL.n11 0.155672
R1570 VTAIL.n36 VTAIL.n35 0.155672
R1571 VTAIL.n36 VTAIL.n7 0.155672
R1572 VTAIL.n43 VTAIL.n7 0.155672
R1573 VTAIL.n44 VTAIL.n43 0.155672
R1574 VTAIL.n44 VTAIL.n3 0.155672
R1575 VTAIL.n51 VTAIL.n3 0.155672
R1576 VTAIL.n161 VTAIL.n113 0.155672
R1577 VTAIL.n154 VTAIL.n113 0.155672
R1578 VTAIL.n154 VTAIL.n153 0.155672
R1579 VTAIL.n153 VTAIL.n117 0.155672
R1580 VTAIL.n146 VTAIL.n117 0.155672
R1581 VTAIL.n146 VTAIL.n145 0.155672
R1582 VTAIL.n145 VTAIL.n121 0.155672
R1583 VTAIL.n138 VTAIL.n121 0.155672
R1584 VTAIL.n138 VTAIL.n137 0.155672
R1585 VTAIL.n137 VTAIL.n125 0.155672
R1586 VTAIL.n130 VTAIL.n125 0.155672
R1587 VTAIL.n107 VTAIL.n59 0.155672
R1588 VTAIL.n100 VTAIL.n59 0.155672
R1589 VTAIL.n100 VTAIL.n99 0.155672
R1590 VTAIL.n99 VTAIL.n63 0.155672
R1591 VTAIL.n92 VTAIL.n63 0.155672
R1592 VTAIL.n92 VTAIL.n91 0.155672
R1593 VTAIL.n91 VTAIL.n67 0.155672
R1594 VTAIL.n84 VTAIL.n67 0.155672
R1595 VTAIL.n84 VTAIL.n83 0.155672
R1596 VTAIL.n83 VTAIL.n71 0.155672
R1597 VTAIL.n76 VTAIL.n71 0.155672
R1598 VDD2.n99 VDD2.n53 289.615
R1599 VDD2.n46 VDD2.n0 289.615
R1600 VDD2.n100 VDD2.n99 185
R1601 VDD2.n98 VDD2.n97 185
R1602 VDD2.n57 VDD2.n56 185
R1603 VDD2.n92 VDD2.n91 185
R1604 VDD2.n90 VDD2.n89 185
R1605 VDD2.n61 VDD2.n60 185
R1606 VDD2.n84 VDD2.n83 185
R1607 VDD2.n82 VDD2.n81 185
R1608 VDD2.n65 VDD2.n64 185
R1609 VDD2.n76 VDD2.n75 185
R1610 VDD2.n74 VDD2.n73 185
R1611 VDD2.n69 VDD2.n68 185
R1612 VDD2.n16 VDD2.n15 185
R1613 VDD2.n21 VDD2.n20 185
R1614 VDD2.n23 VDD2.n22 185
R1615 VDD2.n12 VDD2.n11 185
R1616 VDD2.n29 VDD2.n28 185
R1617 VDD2.n31 VDD2.n30 185
R1618 VDD2.n8 VDD2.n7 185
R1619 VDD2.n37 VDD2.n36 185
R1620 VDD2.n39 VDD2.n38 185
R1621 VDD2.n4 VDD2.n3 185
R1622 VDD2.n45 VDD2.n44 185
R1623 VDD2.n47 VDD2.n46 185
R1624 VDD2.n70 VDD2.t5 147.659
R1625 VDD2.n17 VDD2.t3 147.659
R1626 VDD2.n99 VDD2.n98 104.615
R1627 VDD2.n98 VDD2.n56 104.615
R1628 VDD2.n91 VDD2.n56 104.615
R1629 VDD2.n91 VDD2.n90 104.615
R1630 VDD2.n90 VDD2.n60 104.615
R1631 VDD2.n83 VDD2.n60 104.615
R1632 VDD2.n83 VDD2.n82 104.615
R1633 VDD2.n82 VDD2.n64 104.615
R1634 VDD2.n75 VDD2.n64 104.615
R1635 VDD2.n75 VDD2.n74 104.615
R1636 VDD2.n74 VDD2.n68 104.615
R1637 VDD2.n21 VDD2.n15 104.615
R1638 VDD2.n22 VDD2.n21 104.615
R1639 VDD2.n22 VDD2.n11 104.615
R1640 VDD2.n29 VDD2.n11 104.615
R1641 VDD2.n30 VDD2.n29 104.615
R1642 VDD2.n30 VDD2.n7 104.615
R1643 VDD2.n37 VDD2.n7 104.615
R1644 VDD2.n38 VDD2.n37 104.615
R1645 VDD2.n38 VDD2.n3 104.615
R1646 VDD2.n45 VDD2.n3 104.615
R1647 VDD2.n46 VDD2.n45 104.615
R1648 VDD2.n52 VDD2.n51 61.8975
R1649 VDD2 VDD2.n105 61.8947
R1650 VDD2.t5 VDD2.n68 52.3082
R1651 VDD2.t3 VDD2.n15 52.3082
R1652 VDD2.n52 VDD2.n50 48.1237
R1653 VDD2.n104 VDD2.n103 46.9247
R1654 VDD2.n104 VDD2.n52 37.3403
R1655 VDD2.n70 VDD2.n69 15.6677
R1656 VDD2.n17 VDD2.n16 15.6677
R1657 VDD2.n73 VDD2.n72 12.8005
R1658 VDD2.n20 VDD2.n19 12.8005
R1659 VDD2.n76 VDD2.n67 12.0247
R1660 VDD2.n23 VDD2.n14 12.0247
R1661 VDD2.n77 VDD2.n65 11.249
R1662 VDD2.n24 VDD2.n12 11.249
R1663 VDD2.n81 VDD2.n80 10.4732
R1664 VDD2.n28 VDD2.n27 10.4732
R1665 VDD2.n103 VDD2.n53 9.69747
R1666 VDD2.n84 VDD2.n63 9.69747
R1667 VDD2.n31 VDD2.n10 9.69747
R1668 VDD2.n50 VDD2.n0 9.69747
R1669 VDD2.n103 VDD2.n102 9.45567
R1670 VDD2.n50 VDD2.n49 9.45567
R1671 VDD2.n96 VDD2.n95 9.3005
R1672 VDD2.n55 VDD2.n54 9.3005
R1673 VDD2.n102 VDD2.n101 9.3005
R1674 VDD2.n94 VDD2.n93 9.3005
R1675 VDD2.n59 VDD2.n58 9.3005
R1676 VDD2.n88 VDD2.n87 9.3005
R1677 VDD2.n86 VDD2.n85 9.3005
R1678 VDD2.n63 VDD2.n62 9.3005
R1679 VDD2.n80 VDD2.n79 9.3005
R1680 VDD2.n78 VDD2.n77 9.3005
R1681 VDD2.n67 VDD2.n66 9.3005
R1682 VDD2.n72 VDD2.n71 9.3005
R1683 VDD2.n41 VDD2.n40 9.3005
R1684 VDD2.n43 VDD2.n42 9.3005
R1685 VDD2.n2 VDD2.n1 9.3005
R1686 VDD2.n49 VDD2.n48 9.3005
R1687 VDD2.n35 VDD2.n34 9.3005
R1688 VDD2.n33 VDD2.n32 9.3005
R1689 VDD2.n10 VDD2.n9 9.3005
R1690 VDD2.n27 VDD2.n26 9.3005
R1691 VDD2.n25 VDD2.n24 9.3005
R1692 VDD2.n14 VDD2.n13 9.3005
R1693 VDD2.n19 VDD2.n18 9.3005
R1694 VDD2.n6 VDD2.n5 9.3005
R1695 VDD2.n101 VDD2.n100 8.92171
R1696 VDD2.n85 VDD2.n61 8.92171
R1697 VDD2.n32 VDD2.n8 8.92171
R1698 VDD2.n48 VDD2.n47 8.92171
R1699 VDD2.n97 VDD2.n55 8.14595
R1700 VDD2.n89 VDD2.n88 8.14595
R1701 VDD2.n36 VDD2.n35 8.14595
R1702 VDD2.n44 VDD2.n2 8.14595
R1703 VDD2.n96 VDD2.n57 7.3702
R1704 VDD2.n92 VDD2.n59 7.3702
R1705 VDD2.n39 VDD2.n6 7.3702
R1706 VDD2.n43 VDD2.n4 7.3702
R1707 VDD2.n93 VDD2.n57 6.59444
R1708 VDD2.n93 VDD2.n92 6.59444
R1709 VDD2.n40 VDD2.n39 6.59444
R1710 VDD2.n40 VDD2.n4 6.59444
R1711 VDD2.n97 VDD2.n96 5.81868
R1712 VDD2.n89 VDD2.n59 5.81868
R1713 VDD2.n36 VDD2.n6 5.81868
R1714 VDD2.n44 VDD2.n43 5.81868
R1715 VDD2.n100 VDD2.n55 5.04292
R1716 VDD2.n88 VDD2.n61 5.04292
R1717 VDD2.n35 VDD2.n8 5.04292
R1718 VDD2.n47 VDD2.n2 5.04292
R1719 VDD2.n71 VDD2.n70 4.38563
R1720 VDD2.n18 VDD2.n17 4.38563
R1721 VDD2.n101 VDD2.n53 4.26717
R1722 VDD2.n85 VDD2.n84 4.26717
R1723 VDD2.n32 VDD2.n31 4.26717
R1724 VDD2.n48 VDD2.n0 4.26717
R1725 VDD2.n81 VDD2.n63 3.49141
R1726 VDD2.n28 VDD2.n10 3.49141
R1727 VDD2.n80 VDD2.n65 2.71565
R1728 VDD2.n27 VDD2.n12 2.71565
R1729 VDD2.n105 VDD2.t4 2.08471
R1730 VDD2.n105 VDD2.t1 2.08471
R1731 VDD2.n51 VDD2.t0 2.08471
R1732 VDD2.n51 VDD2.t2 2.08471
R1733 VDD2.n77 VDD2.n76 1.93989
R1734 VDD2.n24 VDD2.n23 1.93989
R1735 VDD2 VDD2.n104 1.313
R1736 VDD2.n73 VDD2.n67 1.16414
R1737 VDD2.n20 VDD2.n14 1.16414
R1738 VDD2.n72 VDD2.n69 0.388379
R1739 VDD2.n19 VDD2.n16 0.388379
R1740 VDD2.n102 VDD2.n54 0.155672
R1741 VDD2.n95 VDD2.n54 0.155672
R1742 VDD2.n95 VDD2.n94 0.155672
R1743 VDD2.n94 VDD2.n58 0.155672
R1744 VDD2.n87 VDD2.n58 0.155672
R1745 VDD2.n87 VDD2.n86 0.155672
R1746 VDD2.n86 VDD2.n62 0.155672
R1747 VDD2.n79 VDD2.n62 0.155672
R1748 VDD2.n79 VDD2.n78 0.155672
R1749 VDD2.n78 VDD2.n66 0.155672
R1750 VDD2.n71 VDD2.n66 0.155672
R1751 VDD2.n18 VDD2.n13 0.155672
R1752 VDD2.n25 VDD2.n13 0.155672
R1753 VDD2.n26 VDD2.n25 0.155672
R1754 VDD2.n26 VDD2.n9 0.155672
R1755 VDD2.n33 VDD2.n9 0.155672
R1756 VDD2.n34 VDD2.n33 0.155672
R1757 VDD2.n34 VDD2.n5 0.155672
R1758 VDD2.n41 VDD2.n5 0.155672
R1759 VDD2.n42 VDD2.n41 0.155672
R1760 VDD2.n42 VDD2.n1 0.155672
R1761 VDD2.n49 VDD2.n1 0.155672
R1762 VP.n17 VP.n16 176.548
R1763 VP.n32 VP.n31 176.548
R1764 VP.n15 VP.n14 176.548
R1765 VP.n6 VP.t2 175.653
R1766 VP.n9 VP.n8 161.3
R1767 VP.n10 VP.n5 161.3
R1768 VP.n12 VP.n11 161.3
R1769 VP.n13 VP.n4 161.3
R1770 VP.n30 VP.n0 161.3
R1771 VP.n29 VP.n28 161.3
R1772 VP.n27 VP.n1 161.3
R1773 VP.n26 VP.n25 161.3
R1774 VP.n23 VP.n2 161.3
R1775 VP.n22 VP.n21 161.3
R1776 VP.n20 VP.n3 161.3
R1777 VP.n19 VP.n18 161.3
R1778 VP.n17 VP.t3 142.206
R1779 VP.n24 VP.t5 142.206
R1780 VP.n31 VP.t1 142.206
R1781 VP.n14 VP.t4 142.206
R1782 VP.n7 VP.t0 142.206
R1783 VP.n22 VP.n3 56.5617
R1784 VP.n29 VP.n1 56.5617
R1785 VP.n12 VP.n5 56.5617
R1786 VP.n7 VP.n6 54.2185
R1787 VP.n16 VP.n15 42.8414
R1788 VP.n18 VP.n3 24.5923
R1789 VP.n23 VP.n22 24.5923
R1790 VP.n25 VP.n1 24.5923
R1791 VP.n30 VP.n29 24.5923
R1792 VP.n13 VP.n12 24.5923
R1793 VP.n8 VP.n5 24.5923
R1794 VP.n9 VP.n6 17.8292
R1795 VP.n24 VP.n23 12.2964
R1796 VP.n25 VP.n24 12.2964
R1797 VP.n8 VP.n7 12.2964
R1798 VP.n18 VP.n17 9.3454
R1799 VP.n31 VP.n30 9.3454
R1800 VP.n14 VP.n13 9.3454
R1801 VP.n10 VP.n9 0.189894
R1802 VP.n11 VP.n10 0.189894
R1803 VP.n11 VP.n4 0.189894
R1804 VP.n15 VP.n4 0.189894
R1805 VP.n19 VP.n16 0.189894
R1806 VP.n20 VP.n19 0.189894
R1807 VP.n21 VP.n20 0.189894
R1808 VP.n21 VP.n2 0.189894
R1809 VP.n26 VP.n2 0.189894
R1810 VP.n27 VP.n26 0.189894
R1811 VP.n28 VP.n27 0.189894
R1812 VP.n28 VP.n0 0.189894
R1813 VP.n32 VP.n0 0.189894
R1814 VP VP.n32 0.0516364
R1815 VDD1.n46 VDD1.n0 289.615
R1816 VDD1.n97 VDD1.n51 289.615
R1817 VDD1.n47 VDD1.n46 185
R1818 VDD1.n45 VDD1.n44 185
R1819 VDD1.n4 VDD1.n3 185
R1820 VDD1.n39 VDD1.n38 185
R1821 VDD1.n37 VDD1.n36 185
R1822 VDD1.n8 VDD1.n7 185
R1823 VDD1.n31 VDD1.n30 185
R1824 VDD1.n29 VDD1.n28 185
R1825 VDD1.n12 VDD1.n11 185
R1826 VDD1.n23 VDD1.n22 185
R1827 VDD1.n21 VDD1.n20 185
R1828 VDD1.n16 VDD1.n15 185
R1829 VDD1.n67 VDD1.n66 185
R1830 VDD1.n72 VDD1.n71 185
R1831 VDD1.n74 VDD1.n73 185
R1832 VDD1.n63 VDD1.n62 185
R1833 VDD1.n80 VDD1.n79 185
R1834 VDD1.n82 VDD1.n81 185
R1835 VDD1.n59 VDD1.n58 185
R1836 VDD1.n88 VDD1.n87 185
R1837 VDD1.n90 VDD1.n89 185
R1838 VDD1.n55 VDD1.n54 185
R1839 VDD1.n96 VDD1.n95 185
R1840 VDD1.n98 VDD1.n97 185
R1841 VDD1.n17 VDD1.t3 147.659
R1842 VDD1.n68 VDD1.t2 147.659
R1843 VDD1.n46 VDD1.n45 104.615
R1844 VDD1.n45 VDD1.n3 104.615
R1845 VDD1.n38 VDD1.n3 104.615
R1846 VDD1.n38 VDD1.n37 104.615
R1847 VDD1.n37 VDD1.n7 104.615
R1848 VDD1.n30 VDD1.n7 104.615
R1849 VDD1.n30 VDD1.n29 104.615
R1850 VDD1.n29 VDD1.n11 104.615
R1851 VDD1.n22 VDD1.n11 104.615
R1852 VDD1.n22 VDD1.n21 104.615
R1853 VDD1.n21 VDD1.n15 104.615
R1854 VDD1.n72 VDD1.n66 104.615
R1855 VDD1.n73 VDD1.n72 104.615
R1856 VDD1.n73 VDD1.n62 104.615
R1857 VDD1.n80 VDD1.n62 104.615
R1858 VDD1.n81 VDD1.n80 104.615
R1859 VDD1.n81 VDD1.n58 104.615
R1860 VDD1.n88 VDD1.n58 104.615
R1861 VDD1.n89 VDD1.n88 104.615
R1862 VDD1.n89 VDD1.n54 104.615
R1863 VDD1.n96 VDD1.n54 104.615
R1864 VDD1.n97 VDD1.n96 104.615
R1865 VDD1.n103 VDD1.n102 61.8975
R1866 VDD1.n105 VDD1.n104 61.5347
R1867 VDD1.t3 VDD1.n15 52.3082
R1868 VDD1.t2 VDD1.n66 52.3082
R1869 VDD1 VDD1.n50 48.2372
R1870 VDD1.n103 VDD1.n101 48.1237
R1871 VDD1.n105 VDD1.n103 38.7595
R1872 VDD1.n17 VDD1.n16 15.6677
R1873 VDD1.n68 VDD1.n67 15.6677
R1874 VDD1.n20 VDD1.n19 12.8005
R1875 VDD1.n71 VDD1.n70 12.8005
R1876 VDD1.n23 VDD1.n14 12.0247
R1877 VDD1.n74 VDD1.n65 12.0247
R1878 VDD1.n24 VDD1.n12 11.249
R1879 VDD1.n75 VDD1.n63 11.249
R1880 VDD1.n28 VDD1.n27 10.4732
R1881 VDD1.n79 VDD1.n78 10.4732
R1882 VDD1.n50 VDD1.n0 9.69747
R1883 VDD1.n31 VDD1.n10 9.69747
R1884 VDD1.n82 VDD1.n61 9.69747
R1885 VDD1.n101 VDD1.n51 9.69747
R1886 VDD1.n50 VDD1.n49 9.45567
R1887 VDD1.n101 VDD1.n100 9.45567
R1888 VDD1.n43 VDD1.n42 9.3005
R1889 VDD1.n2 VDD1.n1 9.3005
R1890 VDD1.n49 VDD1.n48 9.3005
R1891 VDD1.n41 VDD1.n40 9.3005
R1892 VDD1.n6 VDD1.n5 9.3005
R1893 VDD1.n35 VDD1.n34 9.3005
R1894 VDD1.n33 VDD1.n32 9.3005
R1895 VDD1.n10 VDD1.n9 9.3005
R1896 VDD1.n27 VDD1.n26 9.3005
R1897 VDD1.n25 VDD1.n24 9.3005
R1898 VDD1.n14 VDD1.n13 9.3005
R1899 VDD1.n19 VDD1.n18 9.3005
R1900 VDD1.n92 VDD1.n91 9.3005
R1901 VDD1.n94 VDD1.n93 9.3005
R1902 VDD1.n53 VDD1.n52 9.3005
R1903 VDD1.n100 VDD1.n99 9.3005
R1904 VDD1.n86 VDD1.n85 9.3005
R1905 VDD1.n84 VDD1.n83 9.3005
R1906 VDD1.n61 VDD1.n60 9.3005
R1907 VDD1.n78 VDD1.n77 9.3005
R1908 VDD1.n76 VDD1.n75 9.3005
R1909 VDD1.n65 VDD1.n64 9.3005
R1910 VDD1.n70 VDD1.n69 9.3005
R1911 VDD1.n57 VDD1.n56 9.3005
R1912 VDD1.n48 VDD1.n47 8.92171
R1913 VDD1.n32 VDD1.n8 8.92171
R1914 VDD1.n83 VDD1.n59 8.92171
R1915 VDD1.n99 VDD1.n98 8.92171
R1916 VDD1.n44 VDD1.n2 8.14595
R1917 VDD1.n36 VDD1.n35 8.14595
R1918 VDD1.n87 VDD1.n86 8.14595
R1919 VDD1.n95 VDD1.n53 8.14595
R1920 VDD1.n43 VDD1.n4 7.3702
R1921 VDD1.n39 VDD1.n6 7.3702
R1922 VDD1.n90 VDD1.n57 7.3702
R1923 VDD1.n94 VDD1.n55 7.3702
R1924 VDD1.n40 VDD1.n4 6.59444
R1925 VDD1.n40 VDD1.n39 6.59444
R1926 VDD1.n91 VDD1.n90 6.59444
R1927 VDD1.n91 VDD1.n55 6.59444
R1928 VDD1.n44 VDD1.n43 5.81868
R1929 VDD1.n36 VDD1.n6 5.81868
R1930 VDD1.n87 VDD1.n57 5.81868
R1931 VDD1.n95 VDD1.n94 5.81868
R1932 VDD1.n47 VDD1.n2 5.04292
R1933 VDD1.n35 VDD1.n8 5.04292
R1934 VDD1.n86 VDD1.n59 5.04292
R1935 VDD1.n98 VDD1.n53 5.04292
R1936 VDD1.n18 VDD1.n17 4.38563
R1937 VDD1.n69 VDD1.n68 4.38563
R1938 VDD1.n48 VDD1.n0 4.26717
R1939 VDD1.n32 VDD1.n31 4.26717
R1940 VDD1.n83 VDD1.n82 4.26717
R1941 VDD1.n99 VDD1.n51 4.26717
R1942 VDD1.n28 VDD1.n10 3.49141
R1943 VDD1.n79 VDD1.n61 3.49141
R1944 VDD1.n27 VDD1.n12 2.71565
R1945 VDD1.n78 VDD1.n63 2.71565
R1946 VDD1.n104 VDD1.t5 2.08471
R1947 VDD1.n104 VDD1.t1 2.08471
R1948 VDD1.n102 VDD1.t0 2.08471
R1949 VDD1.n102 VDD1.t4 2.08471
R1950 VDD1.n24 VDD1.n23 1.93989
R1951 VDD1.n75 VDD1.n74 1.93989
R1952 VDD1.n20 VDD1.n14 1.16414
R1953 VDD1.n71 VDD1.n65 1.16414
R1954 VDD1.n19 VDD1.n16 0.388379
R1955 VDD1.n70 VDD1.n67 0.388379
R1956 VDD1 VDD1.n105 0.360414
R1957 VDD1.n49 VDD1.n1 0.155672
R1958 VDD1.n42 VDD1.n1 0.155672
R1959 VDD1.n42 VDD1.n41 0.155672
R1960 VDD1.n41 VDD1.n5 0.155672
R1961 VDD1.n34 VDD1.n5 0.155672
R1962 VDD1.n34 VDD1.n33 0.155672
R1963 VDD1.n33 VDD1.n9 0.155672
R1964 VDD1.n26 VDD1.n9 0.155672
R1965 VDD1.n26 VDD1.n25 0.155672
R1966 VDD1.n25 VDD1.n13 0.155672
R1967 VDD1.n18 VDD1.n13 0.155672
R1968 VDD1.n69 VDD1.n64 0.155672
R1969 VDD1.n76 VDD1.n64 0.155672
R1970 VDD1.n77 VDD1.n76 0.155672
R1971 VDD1.n77 VDD1.n60 0.155672
R1972 VDD1.n84 VDD1.n60 0.155672
R1973 VDD1.n85 VDD1.n84 0.155672
R1974 VDD1.n85 VDD1.n56 0.155672
R1975 VDD1.n92 VDD1.n56 0.155672
R1976 VDD1.n93 VDD1.n92 0.155672
R1977 VDD1.n93 VDD1.n52 0.155672
R1978 VDD1.n100 VDD1.n52 0.155672
C0 VDD1 VTAIL 6.79649f
C1 VP VDD1 5.04615f
C2 VDD2 VTAIL 6.8401f
C3 VP VDD2 0.374616f
C4 VDD1 VDD2 1.0487f
C5 VN VTAIL 4.85457f
C6 VP VN 5.49633f
C7 VDD1 VN 0.149787f
C8 VDD2 VN 4.82434f
C9 VP VTAIL 4.86891f
C10 VDD2 B 4.758522f
C11 VDD1 B 4.826814f
C12 VTAIL B 6.154915f
C13 VN B 9.83053f
C14 VP B 8.330711f
C15 VDD1.n0 B 0.032213f
C16 VDD1.n1 B 0.021868f
C17 VDD1.n2 B 0.011751f
C18 VDD1.n3 B 0.027775f
C19 VDD1.n4 B 0.012442f
C20 VDD1.n5 B 0.021868f
C21 VDD1.n6 B 0.011751f
C22 VDD1.n7 B 0.027775f
C23 VDD1.n8 B 0.012442f
C24 VDD1.n9 B 0.021868f
C25 VDD1.n10 B 0.011751f
C26 VDD1.n11 B 0.027775f
C27 VDD1.n12 B 0.012442f
C28 VDD1.n13 B 0.021868f
C29 VDD1.n14 B 0.011751f
C30 VDD1.n15 B 0.020831f
C31 VDD1.n16 B 0.016408f
C32 VDD1.t3 B 0.045391f
C33 VDD1.n17 B 0.112484f
C34 VDD1.n18 B 0.87154f
C35 VDD1.n19 B 0.011751f
C36 VDD1.n20 B 0.012442f
C37 VDD1.n21 B 0.027775f
C38 VDD1.n22 B 0.027775f
C39 VDD1.n23 B 0.012442f
C40 VDD1.n24 B 0.011751f
C41 VDD1.n25 B 0.021868f
C42 VDD1.n26 B 0.021868f
C43 VDD1.n27 B 0.011751f
C44 VDD1.n28 B 0.012442f
C45 VDD1.n29 B 0.027775f
C46 VDD1.n30 B 0.027775f
C47 VDD1.n31 B 0.012442f
C48 VDD1.n32 B 0.011751f
C49 VDD1.n33 B 0.021868f
C50 VDD1.n34 B 0.021868f
C51 VDD1.n35 B 0.011751f
C52 VDD1.n36 B 0.012442f
C53 VDD1.n37 B 0.027775f
C54 VDD1.n38 B 0.027775f
C55 VDD1.n39 B 0.012442f
C56 VDD1.n40 B 0.011751f
C57 VDD1.n41 B 0.021868f
C58 VDD1.n42 B 0.021868f
C59 VDD1.n43 B 0.011751f
C60 VDD1.n44 B 0.012442f
C61 VDD1.n45 B 0.027775f
C62 VDD1.n46 B 0.062738f
C63 VDD1.n47 B 0.012442f
C64 VDD1.n48 B 0.011751f
C65 VDD1.n49 B 0.04756f
C66 VDD1.n50 B 0.054019f
C67 VDD1.n51 B 0.032213f
C68 VDD1.n52 B 0.021868f
C69 VDD1.n53 B 0.011751f
C70 VDD1.n54 B 0.027775f
C71 VDD1.n55 B 0.012442f
C72 VDD1.n56 B 0.021868f
C73 VDD1.n57 B 0.011751f
C74 VDD1.n58 B 0.027775f
C75 VDD1.n59 B 0.012442f
C76 VDD1.n60 B 0.021868f
C77 VDD1.n61 B 0.011751f
C78 VDD1.n62 B 0.027775f
C79 VDD1.n63 B 0.012442f
C80 VDD1.n64 B 0.021868f
C81 VDD1.n65 B 0.011751f
C82 VDD1.n66 B 0.020831f
C83 VDD1.n67 B 0.016408f
C84 VDD1.t2 B 0.045391f
C85 VDD1.n68 B 0.112484f
C86 VDD1.n69 B 0.87154f
C87 VDD1.n70 B 0.011751f
C88 VDD1.n71 B 0.012442f
C89 VDD1.n72 B 0.027775f
C90 VDD1.n73 B 0.027775f
C91 VDD1.n74 B 0.012442f
C92 VDD1.n75 B 0.011751f
C93 VDD1.n76 B 0.021868f
C94 VDD1.n77 B 0.021868f
C95 VDD1.n78 B 0.011751f
C96 VDD1.n79 B 0.012442f
C97 VDD1.n80 B 0.027775f
C98 VDD1.n81 B 0.027775f
C99 VDD1.n82 B 0.012442f
C100 VDD1.n83 B 0.011751f
C101 VDD1.n84 B 0.021868f
C102 VDD1.n85 B 0.021868f
C103 VDD1.n86 B 0.011751f
C104 VDD1.n87 B 0.012442f
C105 VDD1.n88 B 0.027775f
C106 VDD1.n89 B 0.027775f
C107 VDD1.n90 B 0.012442f
C108 VDD1.n91 B 0.011751f
C109 VDD1.n92 B 0.021868f
C110 VDD1.n93 B 0.021868f
C111 VDD1.n94 B 0.011751f
C112 VDD1.n95 B 0.012442f
C113 VDD1.n96 B 0.027775f
C114 VDD1.n97 B 0.062738f
C115 VDD1.n98 B 0.012442f
C116 VDD1.n99 B 0.011751f
C117 VDD1.n100 B 0.04756f
C118 VDD1.n101 B 0.053525f
C119 VDD1.t0 B 0.164169f
C120 VDD1.t4 B 0.164169f
C121 VDD1.n102 B 1.43373f
C122 VDD1.n103 B 1.92374f
C123 VDD1.t5 B 0.164169f
C124 VDD1.t1 B 0.164169f
C125 VDD1.n104 B 1.43174f
C126 VDD1.n105 B 2.03249f
C127 VP.n0 B 0.032345f
C128 VP.t1 B 1.3378f
C129 VP.n1 B 0.044334f
C130 VP.n2 B 0.032345f
C131 VP.t5 B 1.3378f
C132 VP.n3 B 0.049704f
C133 VP.n4 B 0.032345f
C134 VP.t4 B 1.3378f
C135 VP.n5 B 0.044334f
C136 VP.t2 B 1.45663f
C137 VP.n6 B 0.565476f
C138 VP.t0 B 1.3378f
C139 VP.n7 B 0.554622f
C140 VP.n8 B 0.045176f
C141 VP.n9 B 0.207022f
C142 VP.n10 B 0.032345f
C143 VP.n11 B 0.032345f
C144 VP.n12 B 0.049704f
C145 VP.n13 B 0.041623f
C146 VP.n14 B 0.562795f
C147 VP.n15 B 1.38637f
C148 VP.n16 B 1.41359f
C149 VP.t3 B 1.3378f
C150 VP.n17 B 0.562795f
C151 VP.n18 B 0.041623f
C152 VP.n19 B 0.032345f
C153 VP.n20 B 0.032345f
C154 VP.n21 B 0.032345f
C155 VP.n22 B 0.044334f
C156 VP.n23 B 0.045176f
C157 VP.n24 B 0.491761f
C158 VP.n25 B 0.045176f
C159 VP.n26 B 0.032345f
C160 VP.n27 B 0.032345f
C161 VP.n28 B 0.032345f
C162 VP.n29 B 0.049704f
C163 VP.n30 B 0.041623f
C164 VP.n31 B 0.562795f
C165 VP.n32 B 0.031781f
C166 VDD2.n0 B 0.031886f
C167 VDD2.n1 B 0.021646f
C168 VDD2.n2 B 0.011631f
C169 VDD2.n3 B 0.027493f
C170 VDD2.n4 B 0.012316f
C171 VDD2.n5 B 0.021646f
C172 VDD2.n6 B 0.011631f
C173 VDD2.n7 B 0.027493f
C174 VDD2.n8 B 0.012316f
C175 VDD2.n9 B 0.021646f
C176 VDD2.n10 B 0.011631f
C177 VDD2.n11 B 0.027493f
C178 VDD2.n12 B 0.012316f
C179 VDD2.n13 B 0.021646f
C180 VDD2.n14 B 0.011631f
C181 VDD2.n15 B 0.020619f
C182 VDD2.n16 B 0.016241f
C183 VDD2.t3 B 0.044929f
C184 VDD2.n17 B 0.11134f
C185 VDD2.n18 B 0.862673f
C186 VDD2.n19 B 0.011631f
C187 VDD2.n20 B 0.012316f
C188 VDD2.n21 B 0.027493f
C189 VDD2.n22 B 0.027493f
C190 VDD2.n23 B 0.012316f
C191 VDD2.n24 B 0.011631f
C192 VDD2.n25 B 0.021646f
C193 VDD2.n26 B 0.021646f
C194 VDD2.n27 B 0.011631f
C195 VDD2.n28 B 0.012316f
C196 VDD2.n29 B 0.027493f
C197 VDD2.n30 B 0.027493f
C198 VDD2.n31 B 0.012316f
C199 VDD2.n32 B 0.011631f
C200 VDD2.n33 B 0.021646f
C201 VDD2.n34 B 0.021646f
C202 VDD2.n35 B 0.011631f
C203 VDD2.n36 B 0.012316f
C204 VDD2.n37 B 0.027493f
C205 VDD2.n38 B 0.027493f
C206 VDD2.n39 B 0.012316f
C207 VDD2.n40 B 0.011631f
C208 VDD2.n41 B 0.021646f
C209 VDD2.n42 B 0.021646f
C210 VDD2.n43 B 0.011631f
C211 VDD2.n44 B 0.012316f
C212 VDD2.n45 B 0.027493f
C213 VDD2.n46 B 0.062099f
C214 VDD2.n47 B 0.012316f
C215 VDD2.n48 B 0.011631f
C216 VDD2.n49 B 0.047076f
C217 VDD2.n50 B 0.05298f
C218 VDD2.t0 B 0.162499f
C219 VDD2.t2 B 0.162499f
C220 VDD2.n51 B 1.41914f
C221 VDD2.n52 B 1.81984f
C222 VDD2.n53 B 0.031886f
C223 VDD2.n54 B 0.021646f
C224 VDD2.n55 B 0.011631f
C225 VDD2.n56 B 0.027493f
C226 VDD2.n57 B 0.012316f
C227 VDD2.n58 B 0.021646f
C228 VDD2.n59 B 0.011631f
C229 VDD2.n60 B 0.027493f
C230 VDD2.n61 B 0.012316f
C231 VDD2.n62 B 0.021646f
C232 VDD2.n63 B 0.011631f
C233 VDD2.n64 B 0.027493f
C234 VDD2.n65 B 0.012316f
C235 VDD2.n66 B 0.021646f
C236 VDD2.n67 B 0.011631f
C237 VDD2.n68 B 0.020619f
C238 VDD2.n69 B 0.016241f
C239 VDD2.t5 B 0.044929f
C240 VDD2.n70 B 0.11134f
C241 VDD2.n71 B 0.862673f
C242 VDD2.n72 B 0.011631f
C243 VDD2.n73 B 0.012316f
C244 VDD2.n74 B 0.027493f
C245 VDD2.n75 B 0.027493f
C246 VDD2.n76 B 0.012316f
C247 VDD2.n77 B 0.011631f
C248 VDD2.n78 B 0.021646f
C249 VDD2.n79 B 0.021646f
C250 VDD2.n80 B 0.011631f
C251 VDD2.n81 B 0.012316f
C252 VDD2.n82 B 0.027493f
C253 VDD2.n83 B 0.027493f
C254 VDD2.n84 B 0.012316f
C255 VDD2.n85 B 0.011631f
C256 VDD2.n86 B 0.021646f
C257 VDD2.n87 B 0.021646f
C258 VDD2.n88 B 0.011631f
C259 VDD2.n89 B 0.012316f
C260 VDD2.n90 B 0.027493f
C261 VDD2.n91 B 0.027493f
C262 VDD2.n92 B 0.012316f
C263 VDD2.n93 B 0.011631f
C264 VDD2.n94 B 0.021646f
C265 VDD2.n95 B 0.021646f
C266 VDD2.n96 B 0.011631f
C267 VDD2.n97 B 0.012316f
C268 VDD2.n98 B 0.027493f
C269 VDD2.n99 B 0.062099f
C270 VDD2.n100 B 0.012316f
C271 VDD2.n101 B 0.011631f
C272 VDD2.n102 B 0.047076f
C273 VDD2.n103 B 0.04989f
C274 VDD2.n104 B 1.81316f
C275 VDD2.t4 B 0.162499f
C276 VDD2.t1 B 0.162499f
C277 VDD2.n105 B 1.41912f
C278 VTAIL.t10 B 0.180161f
C279 VTAIL.t7 B 0.180161f
C280 VTAIL.n0 B 1.49701f
C281 VTAIL.n1 B 0.383521f
C282 VTAIL.n2 B 0.035351f
C283 VTAIL.n3 B 0.023999f
C284 VTAIL.n4 B 0.012896f
C285 VTAIL.n5 B 0.030481f
C286 VTAIL.n6 B 0.013654f
C287 VTAIL.n7 B 0.023999f
C288 VTAIL.n8 B 0.012896f
C289 VTAIL.n9 B 0.030481f
C290 VTAIL.n10 B 0.013654f
C291 VTAIL.n11 B 0.023999f
C292 VTAIL.n12 B 0.012896f
C293 VTAIL.n13 B 0.030481f
C294 VTAIL.n14 B 0.013654f
C295 VTAIL.n15 B 0.023999f
C296 VTAIL.n16 B 0.012896f
C297 VTAIL.n17 B 0.022861f
C298 VTAIL.n18 B 0.018006f
C299 VTAIL.t0 B 0.049812f
C300 VTAIL.n19 B 0.123442f
C301 VTAIL.n20 B 0.956438f
C302 VTAIL.n21 B 0.012896f
C303 VTAIL.n22 B 0.013654f
C304 VTAIL.n23 B 0.030481f
C305 VTAIL.n24 B 0.030481f
C306 VTAIL.n25 B 0.013654f
C307 VTAIL.n26 B 0.012896f
C308 VTAIL.n27 B 0.023999f
C309 VTAIL.n28 B 0.023999f
C310 VTAIL.n29 B 0.012896f
C311 VTAIL.n30 B 0.013654f
C312 VTAIL.n31 B 0.030481f
C313 VTAIL.n32 B 0.030481f
C314 VTAIL.n33 B 0.013654f
C315 VTAIL.n34 B 0.012896f
C316 VTAIL.n35 B 0.023999f
C317 VTAIL.n36 B 0.023999f
C318 VTAIL.n37 B 0.012896f
C319 VTAIL.n38 B 0.013654f
C320 VTAIL.n39 B 0.030481f
C321 VTAIL.n40 B 0.030481f
C322 VTAIL.n41 B 0.013654f
C323 VTAIL.n42 B 0.012896f
C324 VTAIL.n43 B 0.023999f
C325 VTAIL.n44 B 0.023999f
C326 VTAIL.n45 B 0.012896f
C327 VTAIL.n46 B 0.013654f
C328 VTAIL.n47 B 0.030481f
C329 VTAIL.n48 B 0.068849f
C330 VTAIL.n49 B 0.013654f
C331 VTAIL.n50 B 0.012896f
C332 VTAIL.n51 B 0.052193f
C333 VTAIL.n52 B 0.038714f
C334 VTAIL.n53 B 0.248968f
C335 VTAIL.t3 B 0.180161f
C336 VTAIL.t4 B 0.180161f
C337 VTAIL.n54 B 1.49701f
C338 VTAIL.n55 B 1.59296f
C339 VTAIL.t9 B 0.180161f
C340 VTAIL.t8 B 0.180161f
C341 VTAIL.n56 B 1.49701f
C342 VTAIL.n57 B 1.59295f
C343 VTAIL.n58 B 0.035351f
C344 VTAIL.n59 B 0.023999f
C345 VTAIL.n60 B 0.012896f
C346 VTAIL.n61 B 0.030481f
C347 VTAIL.n62 B 0.013654f
C348 VTAIL.n63 B 0.023999f
C349 VTAIL.n64 B 0.012896f
C350 VTAIL.n65 B 0.030481f
C351 VTAIL.n66 B 0.013654f
C352 VTAIL.n67 B 0.023999f
C353 VTAIL.n68 B 0.012896f
C354 VTAIL.n69 B 0.030481f
C355 VTAIL.n70 B 0.013654f
C356 VTAIL.n71 B 0.023999f
C357 VTAIL.n72 B 0.012896f
C358 VTAIL.n73 B 0.022861f
C359 VTAIL.n74 B 0.018006f
C360 VTAIL.t6 B 0.049812f
C361 VTAIL.n75 B 0.123442f
C362 VTAIL.n76 B 0.956438f
C363 VTAIL.n77 B 0.012896f
C364 VTAIL.n78 B 0.013654f
C365 VTAIL.n79 B 0.030481f
C366 VTAIL.n80 B 0.030481f
C367 VTAIL.n81 B 0.013654f
C368 VTAIL.n82 B 0.012896f
C369 VTAIL.n83 B 0.023999f
C370 VTAIL.n84 B 0.023999f
C371 VTAIL.n85 B 0.012896f
C372 VTAIL.n86 B 0.013654f
C373 VTAIL.n87 B 0.030481f
C374 VTAIL.n88 B 0.030481f
C375 VTAIL.n89 B 0.013654f
C376 VTAIL.n90 B 0.012896f
C377 VTAIL.n91 B 0.023999f
C378 VTAIL.n92 B 0.023999f
C379 VTAIL.n93 B 0.012896f
C380 VTAIL.n94 B 0.013654f
C381 VTAIL.n95 B 0.030481f
C382 VTAIL.n96 B 0.030481f
C383 VTAIL.n97 B 0.013654f
C384 VTAIL.n98 B 0.012896f
C385 VTAIL.n99 B 0.023999f
C386 VTAIL.n100 B 0.023999f
C387 VTAIL.n101 B 0.012896f
C388 VTAIL.n102 B 0.013654f
C389 VTAIL.n103 B 0.030481f
C390 VTAIL.n104 B 0.068849f
C391 VTAIL.n105 B 0.013654f
C392 VTAIL.n106 B 0.012896f
C393 VTAIL.n107 B 0.052193f
C394 VTAIL.n108 B 0.038714f
C395 VTAIL.n109 B 0.248968f
C396 VTAIL.t5 B 0.180161f
C397 VTAIL.t2 B 0.180161f
C398 VTAIL.n110 B 1.49701f
C399 VTAIL.n111 B 0.47601f
C400 VTAIL.n112 B 0.035351f
C401 VTAIL.n113 B 0.023999f
C402 VTAIL.n114 B 0.012896f
C403 VTAIL.n115 B 0.030481f
C404 VTAIL.n116 B 0.013654f
C405 VTAIL.n117 B 0.023999f
C406 VTAIL.n118 B 0.012896f
C407 VTAIL.n119 B 0.030481f
C408 VTAIL.n120 B 0.013654f
C409 VTAIL.n121 B 0.023999f
C410 VTAIL.n122 B 0.012896f
C411 VTAIL.n123 B 0.030481f
C412 VTAIL.n124 B 0.013654f
C413 VTAIL.n125 B 0.023999f
C414 VTAIL.n126 B 0.012896f
C415 VTAIL.n127 B 0.022861f
C416 VTAIL.n128 B 0.018006f
C417 VTAIL.t1 B 0.049812f
C418 VTAIL.n129 B 0.123442f
C419 VTAIL.n130 B 0.956438f
C420 VTAIL.n131 B 0.012896f
C421 VTAIL.n132 B 0.013654f
C422 VTAIL.n133 B 0.030481f
C423 VTAIL.n134 B 0.030481f
C424 VTAIL.n135 B 0.013654f
C425 VTAIL.n136 B 0.012896f
C426 VTAIL.n137 B 0.023999f
C427 VTAIL.n138 B 0.023999f
C428 VTAIL.n139 B 0.012896f
C429 VTAIL.n140 B 0.013654f
C430 VTAIL.n141 B 0.030481f
C431 VTAIL.n142 B 0.030481f
C432 VTAIL.n143 B 0.013654f
C433 VTAIL.n144 B 0.012896f
C434 VTAIL.n145 B 0.023999f
C435 VTAIL.n146 B 0.023999f
C436 VTAIL.n147 B 0.012896f
C437 VTAIL.n148 B 0.013654f
C438 VTAIL.n149 B 0.030481f
C439 VTAIL.n150 B 0.030481f
C440 VTAIL.n151 B 0.013654f
C441 VTAIL.n152 B 0.012896f
C442 VTAIL.n153 B 0.023999f
C443 VTAIL.n154 B 0.023999f
C444 VTAIL.n155 B 0.012896f
C445 VTAIL.n156 B 0.013654f
C446 VTAIL.n157 B 0.030481f
C447 VTAIL.n158 B 0.068849f
C448 VTAIL.n159 B 0.013654f
C449 VTAIL.n160 B 0.012896f
C450 VTAIL.n161 B 0.052193f
C451 VTAIL.n162 B 0.038714f
C452 VTAIL.n163 B 1.23658f
C453 VTAIL.n164 B 0.035351f
C454 VTAIL.n165 B 0.023999f
C455 VTAIL.n166 B 0.012896f
C456 VTAIL.n167 B 0.030481f
C457 VTAIL.n168 B 0.013654f
C458 VTAIL.n169 B 0.023999f
C459 VTAIL.n170 B 0.012896f
C460 VTAIL.n171 B 0.030481f
C461 VTAIL.n172 B 0.013654f
C462 VTAIL.n173 B 0.023999f
C463 VTAIL.n174 B 0.012896f
C464 VTAIL.n175 B 0.030481f
C465 VTAIL.n176 B 0.013654f
C466 VTAIL.n177 B 0.023999f
C467 VTAIL.n178 B 0.012896f
C468 VTAIL.n179 B 0.022861f
C469 VTAIL.n180 B 0.018006f
C470 VTAIL.t11 B 0.049812f
C471 VTAIL.n181 B 0.123442f
C472 VTAIL.n182 B 0.956438f
C473 VTAIL.n183 B 0.012896f
C474 VTAIL.n184 B 0.013654f
C475 VTAIL.n185 B 0.030481f
C476 VTAIL.n186 B 0.030481f
C477 VTAIL.n187 B 0.013654f
C478 VTAIL.n188 B 0.012896f
C479 VTAIL.n189 B 0.023999f
C480 VTAIL.n190 B 0.023999f
C481 VTAIL.n191 B 0.012896f
C482 VTAIL.n192 B 0.013654f
C483 VTAIL.n193 B 0.030481f
C484 VTAIL.n194 B 0.030481f
C485 VTAIL.n195 B 0.013654f
C486 VTAIL.n196 B 0.012896f
C487 VTAIL.n197 B 0.023999f
C488 VTAIL.n198 B 0.023999f
C489 VTAIL.n199 B 0.012896f
C490 VTAIL.n200 B 0.013654f
C491 VTAIL.n201 B 0.030481f
C492 VTAIL.n202 B 0.030481f
C493 VTAIL.n203 B 0.013654f
C494 VTAIL.n204 B 0.012896f
C495 VTAIL.n205 B 0.023999f
C496 VTAIL.n206 B 0.023999f
C497 VTAIL.n207 B 0.012896f
C498 VTAIL.n208 B 0.013654f
C499 VTAIL.n209 B 0.030481f
C500 VTAIL.n210 B 0.068849f
C501 VTAIL.n211 B 0.013654f
C502 VTAIL.n212 B 0.012896f
C503 VTAIL.n213 B 0.052193f
C504 VTAIL.n214 B 0.038714f
C505 VTAIL.n215 B 1.19975f
C506 VN.n0 B 0.031831f
C507 VN.t3 B 1.31654f
C508 VN.n1 B 0.04363f
C509 VN.t2 B 1.43348f
C510 VN.n2 B 0.556489f
C511 VN.t5 B 1.31654f
C512 VN.n3 B 0.545808f
C513 VN.n4 B 0.044458f
C514 VN.n5 B 0.203732f
C515 VN.n6 B 0.031831f
C516 VN.n7 B 0.031831f
C517 VN.n8 B 0.048914f
C518 VN.n9 B 0.040961f
C519 VN.n10 B 0.553851f
C520 VN.n11 B 0.031276f
C521 VN.n12 B 0.031831f
C522 VN.t0 B 1.31654f
C523 VN.n13 B 0.04363f
C524 VN.t4 B 1.43348f
C525 VN.n14 B 0.556489f
C526 VN.t1 B 1.31654f
C527 VN.n15 B 0.545808f
C528 VN.n16 B 0.044458f
C529 VN.n17 B 0.203732f
C530 VN.n18 B 0.031831f
C531 VN.n19 B 0.031831f
C532 VN.n20 B 0.048914f
C533 VN.n21 B 0.040961f
C534 VN.n22 B 0.553851f
C535 VN.n23 B 1.38521f
.ends

