* NGSPICE file created from diff_pair_sample_0062.ext - technology: sky130A

.subckt diff_pair_sample_0062 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t7 VP.t0 VTAIL.t8 w_n4890_n2174# sky130_fd_pr__pfet_01v8 ad=0.99495 pd=6.36 as=0.99495 ps=6.36 w=6.03 l=3.59
X1 VDD1.t6 VP.t1 VTAIL.t10 w_n4890_n2174# sky130_fd_pr__pfet_01v8 ad=0.99495 pd=6.36 as=0.99495 ps=6.36 w=6.03 l=3.59
X2 VDD2.t7 VN.t0 VTAIL.t7 w_n4890_n2174# sky130_fd_pr__pfet_01v8 ad=0.99495 pd=6.36 as=0.99495 ps=6.36 w=6.03 l=3.59
X3 VTAIL.t6 VN.t1 VDD2.t6 w_n4890_n2174# sky130_fd_pr__pfet_01v8 ad=0.99495 pd=6.36 as=0.99495 ps=6.36 w=6.03 l=3.59
X4 VTAIL.t14 VP.t2 VDD1.t5 w_n4890_n2174# sky130_fd_pr__pfet_01v8 ad=2.3517 pd=12.84 as=0.99495 ps=6.36 w=6.03 l=3.59
X5 VDD1.t4 VP.t3 VTAIL.t12 w_n4890_n2174# sky130_fd_pr__pfet_01v8 ad=0.99495 pd=6.36 as=2.3517 ps=12.84 w=6.03 l=3.59
X6 VTAIL.t2 VN.t2 VDD2.t5 w_n4890_n2174# sky130_fd_pr__pfet_01v8 ad=0.99495 pd=6.36 as=0.99495 ps=6.36 w=6.03 l=3.59
X7 B.t11 B.t9 B.t10 w_n4890_n2174# sky130_fd_pr__pfet_01v8 ad=2.3517 pd=12.84 as=0 ps=0 w=6.03 l=3.59
X8 VDD2.t4 VN.t3 VTAIL.t0 w_n4890_n2174# sky130_fd_pr__pfet_01v8 ad=0.99495 pd=6.36 as=2.3517 ps=12.84 w=6.03 l=3.59
X9 VTAIL.t11 VP.t4 VDD1.t3 w_n4890_n2174# sky130_fd_pr__pfet_01v8 ad=2.3517 pd=12.84 as=0.99495 ps=6.36 w=6.03 l=3.59
X10 VDD2.t3 VN.t4 VTAIL.t1 w_n4890_n2174# sky130_fd_pr__pfet_01v8 ad=0.99495 pd=6.36 as=2.3517 ps=12.84 w=6.03 l=3.59
X11 VTAIL.t5 VN.t5 VDD2.t2 w_n4890_n2174# sky130_fd_pr__pfet_01v8 ad=2.3517 pd=12.84 as=0.99495 ps=6.36 w=6.03 l=3.59
X12 VDD1.t2 VP.t5 VTAIL.t15 w_n4890_n2174# sky130_fd_pr__pfet_01v8 ad=0.99495 pd=6.36 as=2.3517 ps=12.84 w=6.03 l=3.59
X13 VTAIL.t3 VN.t6 VDD2.t1 w_n4890_n2174# sky130_fd_pr__pfet_01v8 ad=2.3517 pd=12.84 as=0.99495 ps=6.36 w=6.03 l=3.59
X14 B.t8 B.t6 B.t7 w_n4890_n2174# sky130_fd_pr__pfet_01v8 ad=2.3517 pd=12.84 as=0 ps=0 w=6.03 l=3.59
X15 B.t5 B.t3 B.t4 w_n4890_n2174# sky130_fd_pr__pfet_01v8 ad=2.3517 pd=12.84 as=0 ps=0 w=6.03 l=3.59
X16 VTAIL.t13 VP.t6 VDD1.t1 w_n4890_n2174# sky130_fd_pr__pfet_01v8 ad=0.99495 pd=6.36 as=0.99495 ps=6.36 w=6.03 l=3.59
X17 VDD2.t0 VN.t7 VTAIL.t4 w_n4890_n2174# sky130_fd_pr__pfet_01v8 ad=0.99495 pd=6.36 as=0.99495 ps=6.36 w=6.03 l=3.59
X18 B.t2 B.t0 B.t1 w_n4890_n2174# sky130_fd_pr__pfet_01v8 ad=2.3517 pd=12.84 as=0 ps=0 w=6.03 l=3.59
X19 VTAIL.t9 VP.t7 VDD1.t0 w_n4890_n2174# sky130_fd_pr__pfet_01v8 ad=0.99495 pd=6.36 as=0.99495 ps=6.36 w=6.03 l=3.59
R0 VP.n24 VP.n21 161.3
R1 VP.n26 VP.n25 161.3
R2 VP.n27 VP.n20 161.3
R3 VP.n29 VP.n28 161.3
R4 VP.n30 VP.n19 161.3
R5 VP.n32 VP.n31 161.3
R6 VP.n33 VP.n18 161.3
R7 VP.n36 VP.n35 161.3
R8 VP.n37 VP.n17 161.3
R9 VP.n39 VP.n38 161.3
R10 VP.n40 VP.n16 161.3
R11 VP.n42 VP.n41 161.3
R12 VP.n43 VP.n15 161.3
R13 VP.n45 VP.n44 161.3
R14 VP.n46 VP.n14 161.3
R15 VP.n48 VP.n47 161.3
R16 VP.n89 VP.n88 161.3
R17 VP.n87 VP.n1 161.3
R18 VP.n86 VP.n85 161.3
R19 VP.n84 VP.n2 161.3
R20 VP.n83 VP.n82 161.3
R21 VP.n81 VP.n3 161.3
R22 VP.n80 VP.n79 161.3
R23 VP.n78 VP.n4 161.3
R24 VP.n77 VP.n76 161.3
R25 VP.n74 VP.n5 161.3
R26 VP.n73 VP.n72 161.3
R27 VP.n71 VP.n6 161.3
R28 VP.n70 VP.n69 161.3
R29 VP.n68 VP.n7 161.3
R30 VP.n67 VP.n66 161.3
R31 VP.n65 VP.n8 161.3
R32 VP.n64 VP.n63 161.3
R33 VP.n61 VP.n9 161.3
R34 VP.n60 VP.n59 161.3
R35 VP.n58 VP.n10 161.3
R36 VP.n57 VP.n56 161.3
R37 VP.n55 VP.n11 161.3
R38 VP.n54 VP.n53 161.3
R39 VP.n52 VP.n12 161.3
R40 VP.n51 VP.n50 83.706
R41 VP.n90 VP.n0 83.706
R42 VP.n49 VP.n13 83.706
R43 VP.n23 VP.t4 73.213
R44 VP.n23 VP.n22 64.2098
R45 VP.n56 VP.n10 56.5193
R46 VP.n82 VP.n2 56.5193
R47 VP.n41 VP.n15 56.5193
R48 VP.n69 VP.n6 56.5193
R49 VP.n28 VP.n19 56.5193
R50 VP.n51 VP.n49 51.0599
R51 VP.n50 VP.t2 40.4804
R52 VP.n62 VP.t1 40.4804
R53 VP.n75 VP.t7 40.4804
R54 VP.n0 VP.t5 40.4804
R55 VP.n13 VP.t3 40.4804
R56 VP.n34 VP.t6 40.4804
R57 VP.n22 VP.t0 40.4804
R58 VP.n54 VP.n12 24.4675
R59 VP.n55 VP.n54 24.4675
R60 VP.n56 VP.n55 24.4675
R61 VP.n60 VP.n10 24.4675
R62 VP.n61 VP.n60 24.4675
R63 VP.n63 VP.n61 24.4675
R64 VP.n67 VP.n8 24.4675
R65 VP.n68 VP.n67 24.4675
R66 VP.n69 VP.n68 24.4675
R67 VP.n73 VP.n6 24.4675
R68 VP.n74 VP.n73 24.4675
R69 VP.n76 VP.n74 24.4675
R70 VP.n80 VP.n4 24.4675
R71 VP.n81 VP.n80 24.4675
R72 VP.n82 VP.n81 24.4675
R73 VP.n86 VP.n2 24.4675
R74 VP.n87 VP.n86 24.4675
R75 VP.n88 VP.n87 24.4675
R76 VP.n45 VP.n15 24.4675
R77 VP.n46 VP.n45 24.4675
R78 VP.n47 VP.n46 24.4675
R79 VP.n32 VP.n19 24.4675
R80 VP.n33 VP.n32 24.4675
R81 VP.n35 VP.n33 24.4675
R82 VP.n39 VP.n17 24.4675
R83 VP.n40 VP.n39 24.4675
R84 VP.n41 VP.n40 24.4675
R85 VP.n26 VP.n21 24.4675
R86 VP.n27 VP.n26 24.4675
R87 VP.n28 VP.n27 24.4675
R88 VP.n63 VP.n62 14.1914
R89 VP.n75 VP.n4 14.1914
R90 VP.n34 VP.n17 14.1914
R91 VP.n62 VP.n8 10.2766
R92 VP.n76 VP.n75 10.2766
R93 VP.n35 VP.n34 10.2766
R94 VP.n22 VP.n21 10.2766
R95 VP.n50 VP.n12 6.36192
R96 VP.n88 VP.n0 6.36192
R97 VP.n47 VP.n13 6.36192
R98 VP.n24 VP.n23 3.27565
R99 VP.n49 VP.n48 0.354971
R100 VP.n52 VP.n51 0.354971
R101 VP.n90 VP.n89 0.354971
R102 VP VP.n90 0.26696
R103 VP.n25 VP.n24 0.189894
R104 VP.n25 VP.n20 0.189894
R105 VP.n29 VP.n20 0.189894
R106 VP.n30 VP.n29 0.189894
R107 VP.n31 VP.n30 0.189894
R108 VP.n31 VP.n18 0.189894
R109 VP.n36 VP.n18 0.189894
R110 VP.n37 VP.n36 0.189894
R111 VP.n38 VP.n37 0.189894
R112 VP.n38 VP.n16 0.189894
R113 VP.n42 VP.n16 0.189894
R114 VP.n43 VP.n42 0.189894
R115 VP.n44 VP.n43 0.189894
R116 VP.n44 VP.n14 0.189894
R117 VP.n48 VP.n14 0.189894
R118 VP.n53 VP.n52 0.189894
R119 VP.n53 VP.n11 0.189894
R120 VP.n57 VP.n11 0.189894
R121 VP.n58 VP.n57 0.189894
R122 VP.n59 VP.n58 0.189894
R123 VP.n59 VP.n9 0.189894
R124 VP.n64 VP.n9 0.189894
R125 VP.n65 VP.n64 0.189894
R126 VP.n66 VP.n65 0.189894
R127 VP.n66 VP.n7 0.189894
R128 VP.n70 VP.n7 0.189894
R129 VP.n71 VP.n70 0.189894
R130 VP.n72 VP.n71 0.189894
R131 VP.n72 VP.n5 0.189894
R132 VP.n77 VP.n5 0.189894
R133 VP.n78 VP.n77 0.189894
R134 VP.n79 VP.n78 0.189894
R135 VP.n79 VP.n3 0.189894
R136 VP.n83 VP.n3 0.189894
R137 VP.n84 VP.n83 0.189894
R138 VP.n85 VP.n84 0.189894
R139 VP.n85 VP.n1 0.189894
R140 VP.n89 VP.n1 0.189894
R141 VTAIL.n258 VTAIL.n232 756.745
R142 VTAIL.n28 VTAIL.n2 756.745
R143 VTAIL.n60 VTAIL.n34 756.745
R144 VTAIL.n94 VTAIL.n68 756.745
R145 VTAIL.n226 VTAIL.n200 756.745
R146 VTAIL.n192 VTAIL.n166 756.745
R147 VTAIL.n160 VTAIL.n134 756.745
R148 VTAIL.n126 VTAIL.n100 756.745
R149 VTAIL.n243 VTAIL.n242 585
R150 VTAIL.n240 VTAIL.n239 585
R151 VTAIL.n249 VTAIL.n248 585
R152 VTAIL.n251 VTAIL.n250 585
R153 VTAIL.n236 VTAIL.n235 585
R154 VTAIL.n257 VTAIL.n256 585
R155 VTAIL.n259 VTAIL.n258 585
R156 VTAIL.n13 VTAIL.n12 585
R157 VTAIL.n10 VTAIL.n9 585
R158 VTAIL.n19 VTAIL.n18 585
R159 VTAIL.n21 VTAIL.n20 585
R160 VTAIL.n6 VTAIL.n5 585
R161 VTAIL.n27 VTAIL.n26 585
R162 VTAIL.n29 VTAIL.n28 585
R163 VTAIL.n45 VTAIL.n44 585
R164 VTAIL.n42 VTAIL.n41 585
R165 VTAIL.n51 VTAIL.n50 585
R166 VTAIL.n53 VTAIL.n52 585
R167 VTAIL.n38 VTAIL.n37 585
R168 VTAIL.n59 VTAIL.n58 585
R169 VTAIL.n61 VTAIL.n60 585
R170 VTAIL.n79 VTAIL.n78 585
R171 VTAIL.n76 VTAIL.n75 585
R172 VTAIL.n85 VTAIL.n84 585
R173 VTAIL.n87 VTAIL.n86 585
R174 VTAIL.n72 VTAIL.n71 585
R175 VTAIL.n93 VTAIL.n92 585
R176 VTAIL.n95 VTAIL.n94 585
R177 VTAIL.n227 VTAIL.n226 585
R178 VTAIL.n225 VTAIL.n224 585
R179 VTAIL.n204 VTAIL.n203 585
R180 VTAIL.n219 VTAIL.n218 585
R181 VTAIL.n217 VTAIL.n216 585
R182 VTAIL.n208 VTAIL.n207 585
R183 VTAIL.n211 VTAIL.n210 585
R184 VTAIL.n193 VTAIL.n192 585
R185 VTAIL.n191 VTAIL.n190 585
R186 VTAIL.n170 VTAIL.n169 585
R187 VTAIL.n185 VTAIL.n184 585
R188 VTAIL.n183 VTAIL.n182 585
R189 VTAIL.n174 VTAIL.n173 585
R190 VTAIL.n177 VTAIL.n176 585
R191 VTAIL.n161 VTAIL.n160 585
R192 VTAIL.n159 VTAIL.n158 585
R193 VTAIL.n138 VTAIL.n137 585
R194 VTAIL.n153 VTAIL.n152 585
R195 VTAIL.n151 VTAIL.n150 585
R196 VTAIL.n142 VTAIL.n141 585
R197 VTAIL.n145 VTAIL.n144 585
R198 VTAIL.n127 VTAIL.n126 585
R199 VTAIL.n125 VTAIL.n124 585
R200 VTAIL.n104 VTAIL.n103 585
R201 VTAIL.n119 VTAIL.n118 585
R202 VTAIL.n117 VTAIL.n116 585
R203 VTAIL.n108 VTAIL.n107 585
R204 VTAIL.n111 VTAIL.n110 585
R205 VTAIL.t0 VTAIL.n241 327.601
R206 VTAIL.t5 VTAIL.n11 327.601
R207 VTAIL.t15 VTAIL.n43 327.601
R208 VTAIL.t14 VTAIL.n77 327.601
R209 VTAIL.t12 VTAIL.n209 327.601
R210 VTAIL.t11 VTAIL.n175 327.601
R211 VTAIL.t1 VTAIL.n143 327.601
R212 VTAIL.t3 VTAIL.n109 327.601
R213 VTAIL.n242 VTAIL.n239 171.744
R214 VTAIL.n249 VTAIL.n239 171.744
R215 VTAIL.n250 VTAIL.n249 171.744
R216 VTAIL.n250 VTAIL.n235 171.744
R217 VTAIL.n257 VTAIL.n235 171.744
R218 VTAIL.n258 VTAIL.n257 171.744
R219 VTAIL.n12 VTAIL.n9 171.744
R220 VTAIL.n19 VTAIL.n9 171.744
R221 VTAIL.n20 VTAIL.n19 171.744
R222 VTAIL.n20 VTAIL.n5 171.744
R223 VTAIL.n27 VTAIL.n5 171.744
R224 VTAIL.n28 VTAIL.n27 171.744
R225 VTAIL.n44 VTAIL.n41 171.744
R226 VTAIL.n51 VTAIL.n41 171.744
R227 VTAIL.n52 VTAIL.n51 171.744
R228 VTAIL.n52 VTAIL.n37 171.744
R229 VTAIL.n59 VTAIL.n37 171.744
R230 VTAIL.n60 VTAIL.n59 171.744
R231 VTAIL.n78 VTAIL.n75 171.744
R232 VTAIL.n85 VTAIL.n75 171.744
R233 VTAIL.n86 VTAIL.n85 171.744
R234 VTAIL.n86 VTAIL.n71 171.744
R235 VTAIL.n93 VTAIL.n71 171.744
R236 VTAIL.n94 VTAIL.n93 171.744
R237 VTAIL.n226 VTAIL.n225 171.744
R238 VTAIL.n225 VTAIL.n203 171.744
R239 VTAIL.n218 VTAIL.n203 171.744
R240 VTAIL.n218 VTAIL.n217 171.744
R241 VTAIL.n217 VTAIL.n207 171.744
R242 VTAIL.n210 VTAIL.n207 171.744
R243 VTAIL.n192 VTAIL.n191 171.744
R244 VTAIL.n191 VTAIL.n169 171.744
R245 VTAIL.n184 VTAIL.n169 171.744
R246 VTAIL.n184 VTAIL.n183 171.744
R247 VTAIL.n183 VTAIL.n173 171.744
R248 VTAIL.n176 VTAIL.n173 171.744
R249 VTAIL.n160 VTAIL.n159 171.744
R250 VTAIL.n159 VTAIL.n137 171.744
R251 VTAIL.n152 VTAIL.n137 171.744
R252 VTAIL.n152 VTAIL.n151 171.744
R253 VTAIL.n151 VTAIL.n141 171.744
R254 VTAIL.n144 VTAIL.n141 171.744
R255 VTAIL.n126 VTAIL.n125 171.744
R256 VTAIL.n125 VTAIL.n103 171.744
R257 VTAIL.n118 VTAIL.n103 171.744
R258 VTAIL.n118 VTAIL.n117 171.744
R259 VTAIL.n117 VTAIL.n107 171.744
R260 VTAIL.n110 VTAIL.n107 171.744
R261 VTAIL.n242 VTAIL.t0 85.8723
R262 VTAIL.n12 VTAIL.t5 85.8723
R263 VTAIL.n44 VTAIL.t15 85.8723
R264 VTAIL.n78 VTAIL.t14 85.8723
R265 VTAIL.n210 VTAIL.t12 85.8723
R266 VTAIL.n176 VTAIL.t11 85.8723
R267 VTAIL.n144 VTAIL.t1 85.8723
R268 VTAIL.n110 VTAIL.t3 85.8723
R269 VTAIL.n199 VTAIL.n198 76.1973
R270 VTAIL.n133 VTAIL.n132 76.1973
R271 VTAIL.n1 VTAIL.n0 76.1971
R272 VTAIL.n67 VTAIL.n66 76.1971
R273 VTAIL.n263 VTAIL.n262 32.7672
R274 VTAIL.n33 VTAIL.n32 32.7672
R275 VTAIL.n65 VTAIL.n64 32.7672
R276 VTAIL.n99 VTAIL.n98 32.7672
R277 VTAIL.n231 VTAIL.n230 32.7672
R278 VTAIL.n197 VTAIL.n196 32.7672
R279 VTAIL.n165 VTAIL.n164 32.7672
R280 VTAIL.n131 VTAIL.n130 32.7672
R281 VTAIL.n263 VTAIL.n231 20.9445
R282 VTAIL.n131 VTAIL.n99 20.9445
R283 VTAIL.n243 VTAIL.n241 16.3865
R284 VTAIL.n13 VTAIL.n11 16.3865
R285 VTAIL.n45 VTAIL.n43 16.3865
R286 VTAIL.n79 VTAIL.n77 16.3865
R287 VTAIL.n211 VTAIL.n209 16.3865
R288 VTAIL.n177 VTAIL.n175 16.3865
R289 VTAIL.n145 VTAIL.n143 16.3865
R290 VTAIL.n111 VTAIL.n109 16.3865
R291 VTAIL.n244 VTAIL.n240 12.8005
R292 VTAIL.n14 VTAIL.n10 12.8005
R293 VTAIL.n46 VTAIL.n42 12.8005
R294 VTAIL.n80 VTAIL.n76 12.8005
R295 VTAIL.n212 VTAIL.n208 12.8005
R296 VTAIL.n178 VTAIL.n174 12.8005
R297 VTAIL.n146 VTAIL.n142 12.8005
R298 VTAIL.n112 VTAIL.n108 12.8005
R299 VTAIL.n248 VTAIL.n247 12.0247
R300 VTAIL.n18 VTAIL.n17 12.0247
R301 VTAIL.n50 VTAIL.n49 12.0247
R302 VTAIL.n84 VTAIL.n83 12.0247
R303 VTAIL.n216 VTAIL.n215 12.0247
R304 VTAIL.n182 VTAIL.n181 12.0247
R305 VTAIL.n150 VTAIL.n149 12.0247
R306 VTAIL.n116 VTAIL.n115 12.0247
R307 VTAIL.n251 VTAIL.n238 11.249
R308 VTAIL.n21 VTAIL.n8 11.249
R309 VTAIL.n53 VTAIL.n40 11.249
R310 VTAIL.n87 VTAIL.n74 11.249
R311 VTAIL.n219 VTAIL.n206 11.249
R312 VTAIL.n185 VTAIL.n172 11.249
R313 VTAIL.n153 VTAIL.n140 11.249
R314 VTAIL.n119 VTAIL.n106 11.249
R315 VTAIL.n252 VTAIL.n236 10.4732
R316 VTAIL.n22 VTAIL.n6 10.4732
R317 VTAIL.n54 VTAIL.n38 10.4732
R318 VTAIL.n88 VTAIL.n72 10.4732
R319 VTAIL.n220 VTAIL.n204 10.4732
R320 VTAIL.n186 VTAIL.n170 10.4732
R321 VTAIL.n154 VTAIL.n138 10.4732
R322 VTAIL.n120 VTAIL.n104 10.4732
R323 VTAIL.n256 VTAIL.n255 9.69747
R324 VTAIL.n26 VTAIL.n25 9.69747
R325 VTAIL.n58 VTAIL.n57 9.69747
R326 VTAIL.n92 VTAIL.n91 9.69747
R327 VTAIL.n224 VTAIL.n223 9.69747
R328 VTAIL.n190 VTAIL.n189 9.69747
R329 VTAIL.n158 VTAIL.n157 9.69747
R330 VTAIL.n124 VTAIL.n123 9.69747
R331 VTAIL.n262 VTAIL.n261 9.45567
R332 VTAIL.n32 VTAIL.n31 9.45567
R333 VTAIL.n64 VTAIL.n63 9.45567
R334 VTAIL.n98 VTAIL.n97 9.45567
R335 VTAIL.n230 VTAIL.n229 9.45567
R336 VTAIL.n196 VTAIL.n195 9.45567
R337 VTAIL.n164 VTAIL.n163 9.45567
R338 VTAIL.n130 VTAIL.n129 9.45567
R339 VTAIL.n261 VTAIL.n260 9.3005
R340 VTAIL.n234 VTAIL.n233 9.3005
R341 VTAIL.n255 VTAIL.n254 9.3005
R342 VTAIL.n253 VTAIL.n252 9.3005
R343 VTAIL.n238 VTAIL.n237 9.3005
R344 VTAIL.n247 VTAIL.n246 9.3005
R345 VTAIL.n245 VTAIL.n244 9.3005
R346 VTAIL.n31 VTAIL.n30 9.3005
R347 VTAIL.n4 VTAIL.n3 9.3005
R348 VTAIL.n25 VTAIL.n24 9.3005
R349 VTAIL.n23 VTAIL.n22 9.3005
R350 VTAIL.n8 VTAIL.n7 9.3005
R351 VTAIL.n17 VTAIL.n16 9.3005
R352 VTAIL.n15 VTAIL.n14 9.3005
R353 VTAIL.n63 VTAIL.n62 9.3005
R354 VTAIL.n36 VTAIL.n35 9.3005
R355 VTAIL.n57 VTAIL.n56 9.3005
R356 VTAIL.n55 VTAIL.n54 9.3005
R357 VTAIL.n40 VTAIL.n39 9.3005
R358 VTAIL.n49 VTAIL.n48 9.3005
R359 VTAIL.n47 VTAIL.n46 9.3005
R360 VTAIL.n97 VTAIL.n96 9.3005
R361 VTAIL.n70 VTAIL.n69 9.3005
R362 VTAIL.n91 VTAIL.n90 9.3005
R363 VTAIL.n89 VTAIL.n88 9.3005
R364 VTAIL.n74 VTAIL.n73 9.3005
R365 VTAIL.n83 VTAIL.n82 9.3005
R366 VTAIL.n81 VTAIL.n80 9.3005
R367 VTAIL.n229 VTAIL.n228 9.3005
R368 VTAIL.n202 VTAIL.n201 9.3005
R369 VTAIL.n223 VTAIL.n222 9.3005
R370 VTAIL.n221 VTAIL.n220 9.3005
R371 VTAIL.n206 VTAIL.n205 9.3005
R372 VTAIL.n215 VTAIL.n214 9.3005
R373 VTAIL.n213 VTAIL.n212 9.3005
R374 VTAIL.n195 VTAIL.n194 9.3005
R375 VTAIL.n168 VTAIL.n167 9.3005
R376 VTAIL.n189 VTAIL.n188 9.3005
R377 VTAIL.n187 VTAIL.n186 9.3005
R378 VTAIL.n172 VTAIL.n171 9.3005
R379 VTAIL.n181 VTAIL.n180 9.3005
R380 VTAIL.n179 VTAIL.n178 9.3005
R381 VTAIL.n163 VTAIL.n162 9.3005
R382 VTAIL.n136 VTAIL.n135 9.3005
R383 VTAIL.n157 VTAIL.n156 9.3005
R384 VTAIL.n155 VTAIL.n154 9.3005
R385 VTAIL.n140 VTAIL.n139 9.3005
R386 VTAIL.n149 VTAIL.n148 9.3005
R387 VTAIL.n147 VTAIL.n146 9.3005
R388 VTAIL.n129 VTAIL.n128 9.3005
R389 VTAIL.n102 VTAIL.n101 9.3005
R390 VTAIL.n123 VTAIL.n122 9.3005
R391 VTAIL.n121 VTAIL.n120 9.3005
R392 VTAIL.n106 VTAIL.n105 9.3005
R393 VTAIL.n115 VTAIL.n114 9.3005
R394 VTAIL.n113 VTAIL.n112 9.3005
R395 VTAIL.n259 VTAIL.n234 8.92171
R396 VTAIL.n29 VTAIL.n4 8.92171
R397 VTAIL.n61 VTAIL.n36 8.92171
R398 VTAIL.n95 VTAIL.n70 8.92171
R399 VTAIL.n227 VTAIL.n202 8.92171
R400 VTAIL.n193 VTAIL.n168 8.92171
R401 VTAIL.n161 VTAIL.n136 8.92171
R402 VTAIL.n127 VTAIL.n102 8.92171
R403 VTAIL.n260 VTAIL.n232 8.14595
R404 VTAIL.n30 VTAIL.n2 8.14595
R405 VTAIL.n62 VTAIL.n34 8.14595
R406 VTAIL.n96 VTAIL.n68 8.14595
R407 VTAIL.n228 VTAIL.n200 8.14595
R408 VTAIL.n194 VTAIL.n166 8.14595
R409 VTAIL.n162 VTAIL.n134 8.14595
R410 VTAIL.n128 VTAIL.n100 8.14595
R411 VTAIL.n262 VTAIL.n232 5.81868
R412 VTAIL.n32 VTAIL.n2 5.81868
R413 VTAIL.n64 VTAIL.n34 5.81868
R414 VTAIL.n98 VTAIL.n68 5.81868
R415 VTAIL.n230 VTAIL.n200 5.81868
R416 VTAIL.n196 VTAIL.n166 5.81868
R417 VTAIL.n164 VTAIL.n134 5.81868
R418 VTAIL.n130 VTAIL.n100 5.81868
R419 VTAIL.n0 VTAIL.t4 5.39105
R420 VTAIL.n0 VTAIL.t6 5.39105
R421 VTAIL.n66 VTAIL.t10 5.39105
R422 VTAIL.n66 VTAIL.t9 5.39105
R423 VTAIL.n198 VTAIL.t8 5.39105
R424 VTAIL.n198 VTAIL.t13 5.39105
R425 VTAIL.n132 VTAIL.t7 5.39105
R426 VTAIL.n132 VTAIL.t2 5.39105
R427 VTAIL.n260 VTAIL.n259 5.04292
R428 VTAIL.n30 VTAIL.n29 5.04292
R429 VTAIL.n62 VTAIL.n61 5.04292
R430 VTAIL.n96 VTAIL.n95 5.04292
R431 VTAIL.n228 VTAIL.n227 5.04292
R432 VTAIL.n194 VTAIL.n193 5.04292
R433 VTAIL.n162 VTAIL.n161 5.04292
R434 VTAIL.n128 VTAIL.n127 5.04292
R435 VTAIL.n256 VTAIL.n234 4.26717
R436 VTAIL.n26 VTAIL.n4 4.26717
R437 VTAIL.n58 VTAIL.n36 4.26717
R438 VTAIL.n92 VTAIL.n70 4.26717
R439 VTAIL.n224 VTAIL.n202 4.26717
R440 VTAIL.n190 VTAIL.n168 4.26717
R441 VTAIL.n158 VTAIL.n136 4.26717
R442 VTAIL.n124 VTAIL.n102 4.26717
R443 VTAIL.n213 VTAIL.n209 3.71286
R444 VTAIL.n179 VTAIL.n175 3.71286
R445 VTAIL.n147 VTAIL.n143 3.71286
R446 VTAIL.n113 VTAIL.n109 3.71286
R447 VTAIL.n245 VTAIL.n241 3.71286
R448 VTAIL.n15 VTAIL.n11 3.71286
R449 VTAIL.n47 VTAIL.n43 3.71286
R450 VTAIL.n81 VTAIL.n77 3.71286
R451 VTAIL.n255 VTAIL.n236 3.49141
R452 VTAIL.n25 VTAIL.n6 3.49141
R453 VTAIL.n57 VTAIL.n38 3.49141
R454 VTAIL.n91 VTAIL.n72 3.49141
R455 VTAIL.n223 VTAIL.n204 3.49141
R456 VTAIL.n189 VTAIL.n170 3.49141
R457 VTAIL.n157 VTAIL.n138 3.49141
R458 VTAIL.n123 VTAIL.n104 3.49141
R459 VTAIL.n133 VTAIL.n131 3.37981
R460 VTAIL.n165 VTAIL.n133 3.37981
R461 VTAIL.n199 VTAIL.n197 3.37981
R462 VTAIL.n231 VTAIL.n199 3.37981
R463 VTAIL.n99 VTAIL.n67 3.37981
R464 VTAIL.n67 VTAIL.n65 3.37981
R465 VTAIL.n33 VTAIL.n1 3.37981
R466 VTAIL VTAIL.n263 3.32162
R467 VTAIL.n252 VTAIL.n251 2.71565
R468 VTAIL.n22 VTAIL.n21 2.71565
R469 VTAIL.n54 VTAIL.n53 2.71565
R470 VTAIL.n88 VTAIL.n87 2.71565
R471 VTAIL.n220 VTAIL.n219 2.71565
R472 VTAIL.n186 VTAIL.n185 2.71565
R473 VTAIL.n154 VTAIL.n153 2.71565
R474 VTAIL.n120 VTAIL.n119 2.71565
R475 VTAIL.n248 VTAIL.n238 1.93989
R476 VTAIL.n18 VTAIL.n8 1.93989
R477 VTAIL.n50 VTAIL.n40 1.93989
R478 VTAIL.n84 VTAIL.n74 1.93989
R479 VTAIL.n216 VTAIL.n206 1.93989
R480 VTAIL.n182 VTAIL.n172 1.93989
R481 VTAIL.n150 VTAIL.n140 1.93989
R482 VTAIL.n116 VTAIL.n106 1.93989
R483 VTAIL.n247 VTAIL.n240 1.16414
R484 VTAIL.n17 VTAIL.n10 1.16414
R485 VTAIL.n49 VTAIL.n42 1.16414
R486 VTAIL.n83 VTAIL.n76 1.16414
R487 VTAIL.n215 VTAIL.n208 1.16414
R488 VTAIL.n181 VTAIL.n174 1.16414
R489 VTAIL.n149 VTAIL.n142 1.16414
R490 VTAIL.n115 VTAIL.n108 1.16414
R491 VTAIL.n197 VTAIL.n165 0.470328
R492 VTAIL.n65 VTAIL.n33 0.470328
R493 VTAIL.n244 VTAIL.n243 0.388379
R494 VTAIL.n14 VTAIL.n13 0.388379
R495 VTAIL.n46 VTAIL.n45 0.388379
R496 VTAIL.n80 VTAIL.n79 0.388379
R497 VTAIL.n212 VTAIL.n211 0.388379
R498 VTAIL.n178 VTAIL.n177 0.388379
R499 VTAIL.n146 VTAIL.n145 0.388379
R500 VTAIL.n112 VTAIL.n111 0.388379
R501 VTAIL.n246 VTAIL.n245 0.155672
R502 VTAIL.n246 VTAIL.n237 0.155672
R503 VTAIL.n253 VTAIL.n237 0.155672
R504 VTAIL.n254 VTAIL.n253 0.155672
R505 VTAIL.n254 VTAIL.n233 0.155672
R506 VTAIL.n261 VTAIL.n233 0.155672
R507 VTAIL.n16 VTAIL.n15 0.155672
R508 VTAIL.n16 VTAIL.n7 0.155672
R509 VTAIL.n23 VTAIL.n7 0.155672
R510 VTAIL.n24 VTAIL.n23 0.155672
R511 VTAIL.n24 VTAIL.n3 0.155672
R512 VTAIL.n31 VTAIL.n3 0.155672
R513 VTAIL.n48 VTAIL.n47 0.155672
R514 VTAIL.n48 VTAIL.n39 0.155672
R515 VTAIL.n55 VTAIL.n39 0.155672
R516 VTAIL.n56 VTAIL.n55 0.155672
R517 VTAIL.n56 VTAIL.n35 0.155672
R518 VTAIL.n63 VTAIL.n35 0.155672
R519 VTAIL.n82 VTAIL.n81 0.155672
R520 VTAIL.n82 VTAIL.n73 0.155672
R521 VTAIL.n89 VTAIL.n73 0.155672
R522 VTAIL.n90 VTAIL.n89 0.155672
R523 VTAIL.n90 VTAIL.n69 0.155672
R524 VTAIL.n97 VTAIL.n69 0.155672
R525 VTAIL.n229 VTAIL.n201 0.155672
R526 VTAIL.n222 VTAIL.n201 0.155672
R527 VTAIL.n222 VTAIL.n221 0.155672
R528 VTAIL.n221 VTAIL.n205 0.155672
R529 VTAIL.n214 VTAIL.n205 0.155672
R530 VTAIL.n214 VTAIL.n213 0.155672
R531 VTAIL.n195 VTAIL.n167 0.155672
R532 VTAIL.n188 VTAIL.n167 0.155672
R533 VTAIL.n188 VTAIL.n187 0.155672
R534 VTAIL.n187 VTAIL.n171 0.155672
R535 VTAIL.n180 VTAIL.n171 0.155672
R536 VTAIL.n180 VTAIL.n179 0.155672
R537 VTAIL.n163 VTAIL.n135 0.155672
R538 VTAIL.n156 VTAIL.n135 0.155672
R539 VTAIL.n156 VTAIL.n155 0.155672
R540 VTAIL.n155 VTAIL.n139 0.155672
R541 VTAIL.n148 VTAIL.n139 0.155672
R542 VTAIL.n148 VTAIL.n147 0.155672
R543 VTAIL.n129 VTAIL.n101 0.155672
R544 VTAIL.n122 VTAIL.n101 0.155672
R545 VTAIL.n122 VTAIL.n121 0.155672
R546 VTAIL.n121 VTAIL.n105 0.155672
R547 VTAIL.n114 VTAIL.n105 0.155672
R548 VTAIL.n114 VTAIL.n113 0.155672
R549 VTAIL VTAIL.n1 0.0586897
R550 VDD1 VDD1.n0 94.6239
R551 VDD1.n3 VDD1.n2 94.5102
R552 VDD1.n3 VDD1.n1 94.5102
R553 VDD1.n5 VDD1.n4 92.8759
R554 VDD1.n5 VDD1.n3 44.7035
R555 VDD1.n4 VDD1.t1 5.39105
R556 VDD1.n4 VDD1.t4 5.39105
R557 VDD1.n0 VDD1.t3 5.39105
R558 VDD1.n0 VDD1.t7 5.39105
R559 VDD1.n2 VDD1.t0 5.39105
R560 VDD1.n2 VDD1.t2 5.39105
R561 VDD1.n1 VDD1.t5 5.39105
R562 VDD1.n1 VDD1.t6 5.39105
R563 VDD1 VDD1.n5 1.63197
R564 VN.n72 VN.n71 161.3
R565 VN.n70 VN.n38 161.3
R566 VN.n69 VN.n68 161.3
R567 VN.n67 VN.n39 161.3
R568 VN.n66 VN.n65 161.3
R569 VN.n64 VN.n40 161.3
R570 VN.n63 VN.n62 161.3
R571 VN.n61 VN.n41 161.3
R572 VN.n60 VN.n59 161.3
R573 VN.n58 VN.n42 161.3
R574 VN.n57 VN.n56 161.3
R575 VN.n55 VN.n44 161.3
R576 VN.n54 VN.n53 161.3
R577 VN.n52 VN.n45 161.3
R578 VN.n51 VN.n50 161.3
R579 VN.n49 VN.n46 161.3
R580 VN.n35 VN.n34 161.3
R581 VN.n33 VN.n1 161.3
R582 VN.n32 VN.n31 161.3
R583 VN.n30 VN.n2 161.3
R584 VN.n29 VN.n28 161.3
R585 VN.n27 VN.n3 161.3
R586 VN.n26 VN.n25 161.3
R587 VN.n24 VN.n4 161.3
R588 VN.n23 VN.n22 161.3
R589 VN.n20 VN.n5 161.3
R590 VN.n19 VN.n18 161.3
R591 VN.n17 VN.n6 161.3
R592 VN.n16 VN.n15 161.3
R593 VN.n14 VN.n7 161.3
R594 VN.n13 VN.n12 161.3
R595 VN.n11 VN.n8 161.3
R596 VN.n36 VN.n0 83.706
R597 VN.n73 VN.n37 83.706
R598 VN.n48 VN.t4 73.2132
R599 VN.n10 VN.t5 73.2132
R600 VN.n10 VN.n9 64.2098
R601 VN.n48 VN.n47 64.2098
R602 VN.n28 VN.n2 56.5193
R603 VN.n65 VN.n39 56.5193
R604 VN.n15 VN.n6 56.5193
R605 VN.n53 VN.n44 56.5193
R606 VN VN.n73 51.2253
R607 VN.n9 VN.t7 40.4804
R608 VN.n21 VN.t1 40.4804
R609 VN.n0 VN.t3 40.4804
R610 VN.n47 VN.t2 40.4804
R611 VN.n43 VN.t0 40.4804
R612 VN.n37 VN.t6 40.4804
R613 VN.n13 VN.n8 24.4675
R614 VN.n14 VN.n13 24.4675
R615 VN.n15 VN.n14 24.4675
R616 VN.n19 VN.n6 24.4675
R617 VN.n20 VN.n19 24.4675
R618 VN.n22 VN.n20 24.4675
R619 VN.n26 VN.n4 24.4675
R620 VN.n27 VN.n26 24.4675
R621 VN.n28 VN.n27 24.4675
R622 VN.n32 VN.n2 24.4675
R623 VN.n33 VN.n32 24.4675
R624 VN.n34 VN.n33 24.4675
R625 VN.n53 VN.n52 24.4675
R626 VN.n52 VN.n51 24.4675
R627 VN.n51 VN.n46 24.4675
R628 VN.n65 VN.n64 24.4675
R629 VN.n64 VN.n63 24.4675
R630 VN.n63 VN.n41 24.4675
R631 VN.n59 VN.n58 24.4675
R632 VN.n58 VN.n57 24.4675
R633 VN.n57 VN.n44 24.4675
R634 VN.n71 VN.n70 24.4675
R635 VN.n70 VN.n69 24.4675
R636 VN.n69 VN.n39 24.4675
R637 VN.n21 VN.n4 14.1914
R638 VN.n43 VN.n41 14.1914
R639 VN.n9 VN.n8 10.2766
R640 VN.n22 VN.n21 10.2766
R641 VN.n47 VN.n46 10.2766
R642 VN.n59 VN.n43 10.2766
R643 VN.n34 VN.n0 6.36192
R644 VN.n71 VN.n37 6.36192
R645 VN.n11 VN.n10 3.27566
R646 VN.n49 VN.n48 3.27566
R647 VN.n73 VN.n72 0.354971
R648 VN.n36 VN.n35 0.354971
R649 VN VN.n36 0.26696
R650 VN.n72 VN.n38 0.189894
R651 VN.n68 VN.n38 0.189894
R652 VN.n68 VN.n67 0.189894
R653 VN.n67 VN.n66 0.189894
R654 VN.n66 VN.n40 0.189894
R655 VN.n62 VN.n40 0.189894
R656 VN.n62 VN.n61 0.189894
R657 VN.n61 VN.n60 0.189894
R658 VN.n60 VN.n42 0.189894
R659 VN.n56 VN.n42 0.189894
R660 VN.n56 VN.n55 0.189894
R661 VN.n55 VN.n54 0.189894
R662 VN.n54 VN.n45 0.189894
R663 VN.n50 VN.n45 0.189894
R664 VN.n50 VN.n49 0.189894
R665 VN.n12 VN.n11 0.189894
R666 VN.n12 VN.n7 0.189894
R667 VN.n16 VN.n7 0.189894
R668 VN.n17 VN.n16 0.189894
R669 VN.n18 VN.n17 0.189894
R670 VN.n18 VN.n5 0.189894
R671 VN.n23 VN.n5 0.189894
R672 VN.n24 VN.n23 0.189894
R673 VN.n25 VN.n24 0.189894
R674 VN.n25 VN.n3 0.189894
R675 VN.n29 VN.n3 0.189894
R676 VN.n30 VN.n29 0.189894
R677 VN.n31 VN.n30 0.189894
R678 VN.n31 VN.n1 0.189894
R679 VN.n35 VN.n1 0.189894
R680 VDD2.n2 VDD2.n1 94.5102
R681 VDD2.n2 VDD2.n0 94.5102
R682 VDD2 VDD2.n5 94.5074
R683 VDD2.n4 VDD2.n3 92.8761
R684 VDD2.n4 VDD2.n2 44.1205
R685 VDD2.n5 VDD2.t5 5.39105
R686 VDD2.n5 VDD2.t3 5.39105
R687 VDD2.n3 VDD2.t1 5.39105
R688 VDD2.n3 VDD2.t7 5.39105
R689 VDD2.n1 VDD2.t6 5.39105
R690 VDD2.n1 VDD2.t4 5.39105
R691 VDD2.n0 VDD2.t2 5.39105
R692 VDD2.n0 VDD2.t0 5.39105
R693 VDD2 VDD2.n4 1.74834
R694 B.n384 B.n383 585
R695 B.n382 B.n135 585
R696 B.n381 B.n380 585
R697 B.n379 B.n136 585
R698 B.n378 B.n377 585
R699 B.n376 B.n137 585
R700 B.n375 B.n374 585
R701 B.n373 B.n138 585
R702 B.n372 B.n371 585
R703 B.n370 B.n139 585
R704 B.n369 B.n368 585
R705 B.n367 B.n140 585
R706 B.n366 B.n365 585
R707 B.n364 B.n141 585
R708 B.n363 B.n362 585
R709 B.n361 B.n142 585
R710 B.n360 B.n359 585
R711 B.n358 B.n143 585
R712 B.n357 B.n356 585
R713 B.n355 B.n144 585
R714 B.n354 B.n353 585
R715 B.n352 B.n145 585
R716 B.n351 B.n350 585
R717 B.n349 B.n146 585
R718 B.n347 B.n346 585
R719 B.n345 B.n149 585
R720 B.n344 B.n343 585
R721 B.n342 B.n150 585
R722 B.n341 B.n340 585
R723 B.n339 B.n151 585
R724 B.n338 B.n337 585
R725 B.n336 B.n152 585
R726 B.n335 B.n334 585
R727 B.n333 B.n153 585
R728 B.n332 B.n331 585
R729 B.n327 B.n154 585
R730 B.n326 B.n325 585
R731 B.n324 B.n155 585
R732 B.n323 B.n322 585
R733 B.n321 B.n156 585
R734 B.n320 B.n319 585
R735 B.n318 B.n157 585
R736 B.n317 B.n316 585
R737 B.n315 B.n158 585
R738 B.n314 B.n313 585
R739 B.n312 B.n159 585
R740 B.n311 B.n310 585
R741 B.n309 B.n160 585
R742 B.n308 B.n307 585
R743 B.n306 B.n161 585
R744 B.n305 B.n304 585
R745 B.n303 B.n162 585
R746 B.n302 B.n301 585
R747 B.n300 B.n163 585
R748 B.n299 B.n298 585
R749 B.n297 B.n164 585
R750 B.n296 B.n295 585
R751 B.n294 B.n165 585
R752 B.n385 B.n134 585
R753 B.n387 B.n386 585
R754 B.n388 B.n133 585
R755 B.n390 B.n389 585
R756 B.n391 B.n132 585
R757 B.n393 B.n392 585
R758 B.n394 B.n131 585
R759 B.n396 B.n395 585
R760 B.n397 B.n130 585
R761 B.n399 B.n398 585
R762 B.n400 B.n129 585
R763 B.n402 B.n401 585
R764 B.n403 B.n128 585
R765 B.n405 B.n404 585
R766 B.n406 B.n127 585
R767 B.n408 B.n407 585
R768 B.n409 B.n126 585
R769 B.n411 B.n410 585
R770 B.n412 B.n125 585
R771 B.n414 B.n413 585
R772 B.n415 B.n124 585
R773 B.n417 B.n416 585
R774 B.n418 B.n123 585
R775 B.n420 B.n419 585
R776 B.n421 B.n122 585
R777 B.n423 B.n422 585
R778 B.n424 B.n121 585
R779 B.n426 B.n425 585
R780 B.n427 B.n120 585
R781 B.n429 B.n428 585
R782 B.n430 B.n119 585
R783 B.n432 B.n431 585
R784 B.n433 B.n118 585
R785 B.n435 B.n434 585
R786 B.n436 B.n117 585
R787 B.n438 B.n437 585
R788 B.n439 B.n116 585
R789 B.n441 B.n440 585
R790 B.n442 B.n115 585
R791 B.n444 B.n443 585
R792 B.n445 B.n114 585
R793 B.n447 B.n446 585
R794 B.n448 B.n113 585
R795 B.n450 B.n449 585
R796 B.n451 B.n112 585
R797 B.n453 B.n452 585
R798 B.n454 B.n111 585
R799 B.n456 B.n455 585
R800 B.n457 B.n110 585
R801 B.n459 B.n458 585
R802 B.n460 B.n109 585
R803 B.n462 B.n461 585
R804 B.n463 B.n108 585
R805 B.n465 B.n464 585
R806 B.n466 B.n107 585
R807 B.n468 B.n467 585
R808 B.n469 B.n106 585
R809 B.n471 B.n470 585
R810 B.n472 B.n105 585
R811 B.n474 B.n473 585
R812 B.n475 B.n104 585
R813 B.n477 B.n476 585
R814 B.n478 B.n103 585
R815 B.n480 B.n479 585
R816 B.n481 B.n102 585
R817 B.n483 B.n482 585
R818 B.n484 B.n101 585
R819 B.n486 B.n485 585
R820 B.n487 B.n100 585
R821 B.n489 B.n488 585
R822 B.n490 B.n99 585
R823 B.n492 B.n491 585
R824 B.n493 B.n98 585
R825 B.n495 B.n494 585
R826 B.n496 B.n97 585
R827 B.n498 B.n497 585
R828 B.n499 B.n96 585
R829 B.n501 B.n500 585
R830 B.n502 B.n95 585
R831 B.n504 B.n503 585
R832 B.n505 B.n94 585
R833 B.n507 B.n506 585
R834 B.n508 B.n93 585
R835 B.n510 B.n509 585
R836 B.n511 B.n92 585
R837 B.n513 B.n512 585
R838 B.n514 B.n91 585
R839 B.n516 B.n515 585
R840 B.n517 B.n90 585
R841 B.n519 B.n518 585
R842 B.n520 B.n89 585
R843 B.n522 B.n521 585
R844 B.n523 B.n88 585
R845 B.n525 B.n524 585
R846 B.n526 B.n87 585
R847 B.n528 B.n527 585
R848 B.n529 B.n86 585
R849 B.n531 B.n530 585
R850 B.n532 B.n85 585
R851 B.n534 B.n533 585
R852 B.n535 B.n84 585
R853 B.n537 B.n536 585
R854 B.n538 B.n83 585
R855 B.n540 B.n539 585
R856 B.n541 B.n82 585
R857 B.n543 B.n542 585
R858 B.n544 B.n81 585
R859 B.n546 B.n545 585
R860 B.n547 B.n80 585
R861 B.n549 B.n548 585
R862 B.n550 B.n79 585
R863 B.n552 B.n551 585
R864 B.n553 B.n78 585
R865 B.n555 B.n554 585
R866 B.n556 B.n77 585
R867 B.n558 B.n557 585
R868 B.n559 B.n76 585
R869 B.n561 B.n560 585
R870 B.n562 B.n75 585
R871 B.n564 B.n563 585
R872 B.n565 B.n74 585
R873 B.n567 B.n566 585
R874 B.n568 B.n73 585
R875 B.n570 B.n569 585
R876 B.n571 B.n72 585
R877 B.n573 B.n572 585
R878 B.n574 B.n71 585
R879 B.n576 B.n575 585
R880 B.n577 B.n70 585
R881 B.n579 B.n578 585
R882 B.n580 B.n69 585
R883 B.n582 B.n581 585
R884 B.n670 B.n669 585
R885 B.n668 B.n35 585
R886 B.n667 B.n666 585
R887 B.n665 B.n36 585
R888 B.n664 B.n663 585
R889 B.n662 B.n37 585
R890 B.n661 B.n660 585
R891 B.n659 B.n38 585
R892 B.n658 B.n657 585
R893 B.n656 B.n39 585
R894 B.n655 B.n654 585
R895 B.n653 B.n40 585
R896 B.n652 B.n651 585
R897 B.n650 B.n41 585
R898 B.n649 B.n648 585
R899 B.n647 B.n42 585
R900 B.n646 B.n645 585
R901 B.n644 B.n43 585
R902 B.n643 B.n642 585
R903 B.n641 B.n44 585
R904 B.n640 B.n639 585
R905 B.n638 B.n45 585
R906 B.n637 B.n636 585
R907 B.n635 B.n46 585
R908 B.n634 B.n633 585
R909 B.n632 B.n47 585
R910 B.n631 B.n630 585
R911 B.n629 B.n51 585
R912 B.n628 B.n627 585
R913 B.n626 B.n52 585
R914 B.n625 B.n624 585
R915 B.n623 B.n53 585
R916 B.n622 B.n621 585
R917 B.n620 B.n54 585
R918 B.n618 B.n617 585
R919 B.n616 B.n57 585
R920 B.n615 B.n614 585
R921 B.n613 B.n58 585
R922 B.n612 B.n611 585
R923 B.n610 B.n59 585
R924 B.n609 B.n608 585
R925 B.n607 B.n60 585
R926 B.n606 B.n605 585
R927 B.n604 B.n61 585
R928 B.n603 B.n602 585
R929 B.n601 B.n62 585
R930 B.n600 B.n599 585
R931 B.n598 B.n63 585
R932 B.n597 B.n596 585
R933 B.n595 B.n64 585
R934 B.n594 B.n593 585
R935 B.n592 B.n65 585
R936 B.n591 B.n590 585
R937 B.n589 B.n66 585
R938 B.n588 B.n587 585
R939 B.n586 B.n67 585
R940 B.n585 B.n584 585
R941 B.n583 B.n68 585
R942 B.n671 B.n34 585
R943 B.n673 B.n672 585
R944 B.n674 B.n33 585
R945 B.n676 B.n675 585
R946 B.n677 B.n32 585
R947 B.n679 B.n678 585
R948 B.n680 B.n31 585
R949 B.n682 B.n681 585
R950 B.n683 B.n30 585
R951 B.n685 B.n684 585
R952 B.n686 B.n29 585
R953 B.n688 B.n687 585
R954 B.n689 B.n28 585
R955 B.n691 B.n690 585
R956 B.n692 B.n27 585
R957 B.n694 B.n693 585
R958 B.n695 B.n26 585
R959 B.n697 B.n696 585
R960 B.n698 B.n25 585
R961 B.n700 B.n699 585
R962 B.n701 B.n24 585
R963 B.n703 B.n702 585
R964 B.n704 B.n23 585
R965 B.n706 B.n705 585
R966 B.n707 B.n22 585
R967 B.n709 B.n708 585
R968 B.n710 B.n21 585
R969 B.n712 B.n711 585
R970 B.n713 B.n20 585
R971 B.n715 B.n714 585
R972 B.n716 B.n19 585
R973 B.n718 B.n717 585
R974 B.n719 B.n18 585
R975 B.n721 B.n720 585
R976 B.n722 B.n17 585
R977 B.n724 B.n723 585
R978 B.n725 B.n16 585
R979 B.n727 B.n726 585
R980 B.n728 B.n15 585
R981 B.n730 B.n729 585
R982 B.n731 B.n14 585
R983 B.n733 B.n732 585
R984 B.n734 B.n13 585
R985 B.n736 B.n735 585
R986 B.n737 B.n12 585
R987 B.n739 B.n738 585
R988 B.n740 B.n11 585
R989 B.n742 B.n741 585
R990 B.n743 B.n10 585
R991 B.n745 B.n744 585
R992 B.n746 B.n9 585
R993 B.n748 B.n747 585
R994 B.n749 B.n8 585
R995 B.n751 B.n750 585
R996 B.n752 B.n7 585
R997 B.n754 B.n753 585
R998 B.n755 B.n6 585
R999 B.n757 B.n756 585
R1000 B.n758 B.n5 585
R1001 B.n760 B.n759 585
R1002 B.n761 B.n4 585
R1003 B.n763 B.n762 585
R1004 B.n764 B.n3 585
R1005 B.n766 B.n765 585
R1006 B.n767 B.n0 585
R1007 B.n2 B.n1 585
R1008 B.n198 B.n197 585
R1009 B.n200 B.n199 585
R1010 B.n201 B.n196 585
R1011 B.n203 B.n202 585
R1012 B.n204 B.n195 585
R1013 B.n206 B.n205 585
R1014 B.n207 B.n194 585
R1015 B.n209 B.n208 585
R1016 B.n210 B.n193 585
R1017 B.n212 B.n211 585
R1018 B.n213 B.n192 585
R1019 B.n215 B.n214 585
R1020 B.n216 B.n191 585
R1021 B.n218 B.n217 585
R1022 B.n219 B.n190 585
R1023 B.n221 B.n220 585
R1024 B.n222 B.n189 585
R1025 B.n224 B.n223 585
R1026 B.n225 B.n188 585
R1027 B.n227 B.n226 585
R1028 B.n228 B.n187 585
R1029 B.n230 B.n229 585
R1030 B.n231 B.n186 585
R1031 B.n233 B.n232 585
R1032 B.n234 B.n185 585
R1033 B.n236 B.n235 585
R1034 B.n237 B.n184 585
R1035 B.n239 B.n238 585
R1036 B.n240 B.n183 585
R1037 B.n242 B.n241 585
R1038 B.n243 B.n182 585
R1039 B.n245 B.n244 585
R1040 B.n246 B.n181 585
R1041 B.n248 B.n247 585
R1042 B.n249 B.n180 585
R1043 B.n251 B.n250 585
R1044 B.n252 B.n179 585
R1045 B.n254 B.n253 585
R1046 B.n255 B.n178 585
R1047 B.n257 B.n256 585
R1048 B.n258 B.n177 585
R1049 B.n260 B.n259 585
R1050 B.n261 B.n176 585
R1051 B.n263 B.n262 585
R1052 B.n264 B.n175 585
R1053 B.n266 B.n265 585
R1054 B.n267 B.n174 585
R1055 B.n269 B.n268 585
R1056 B.n270 B.n173 585
R1057 B.n272 B.n271 585
R1058 B.n273 B.n172 585
R1059 B.n275 B.n274 585
R1060 B.n276 B.n171 585
R1061 B.n278 B.n277 585
R1062 B.n279 B.n170 585
R1063 B.n281 B.n280 585
R1064 B.n282 B.n169 585
R1065 B.n284 B.n283 585
R1066 B.n285 B.n168 585
R1067 B.n287 B.n286 585
R1068 B.n288 B.n167 585
R1069 B.n290 B.n289 585
R1070 B.n291 B.n166 585
R1071 B.n293 B.n292 585
R1072 B.n294 B.n293 516.524
R1073 B.n383 B.n134 516.524
R1074 B.n581 B.n68 516.524
R1075 B.n671 B.n670 516.524
R1076 B.n147 B.t1 344.8
R1077 B.n55 B.t5 344.8
R1078 B.n328 B.t10 344.798
R1079 B.n48 B.t8 344.798
R1080 B.n148 B.t2 268.774
R1081 B.n56 B.t4 268.774
R1082 B.n329 B.t11 268.774
R1083 B.n49 B.t7 268.774
R1084 B.n769 B.n768 256.663
R1085 B.n328 B.t9 249.653
R1086 B.n147 B.t0 249.653
R1087 B.n55 B.t3 249.653
R1088 B.n48 B.t6 249.653
R1089 B.n768 B.n767 235.042
R1090 B.n768 B.n2 235.042
R1091 B.n295 B.n294 163.367
R1092 B.n295 B.n164 163.367
R1093 B.n299 B.n164 163.367
R1094 B.n300 B.n299 163.367
R1095 B.n301 B.n300 163.367
R1096 B.n301 B.n162 163.367
R1097 B.n305 B.n162 163.367
R1098 B.n306 B.n305 163.367
R1099 B.n307 B.n306 163.367
R1100 B.n307 B.n160 163.367
R1101 B.n311 B.n160 163.367
R1102 B.n312 B.n311 163.367
R1103 B.n313 B.n312 163.367
R1104 B.n313 B.n158 163.367
R1105 B.n317 B.n158 163.367
R1106 B.n318 B.n317 163.367
R1107 B.n319 B.n318 163.367
R1108 B.n319 B.n156 163.367
R1109 B.n323 B.n156 163.367
R1110 B.n324 B.n323 163.367
R1111 B.n325 B.n324 163.367
R1112 B.n325 B.n154 163.367
R1113 B.n332 B.n154 163.367
R1114 B.n333 B.n332 163.367
R1115 B.n334 B.n333 163.367
R1116 B.n334 B.n152 163.367
R1117 B.n338 B.n152 163.367
R1118 B.n339 B.n338 163.367
R1119 B.n340 B.n339 163.367
R1120 B.n340 B.n150 163.367
R1121 B.n344 B.n150 163.367
R1122 B.n345 B.n344 163.367
R1123 B.n346 B.n345 163.367
R1124 B.n346 B.n146 163.367
R1125 B.n351 B.n146 163.367
R1126 B.n352 B.n351 163.367
R1127 B.n353 B.n352 163.367
R1128 B.n353 B.n144 163.367
R1129 B.n357 B.n144 163.367
R1130 B.n358 B.n357 163.367
R1131 B.n359 B.n358 163.367
R1132 B.n359 B.n142 163.367
R1133 B.n363 B.n142 163.367
R1134 B.n364 B.n363 163.367
R1135 B.n365 B.n364 163.367
R1136 B.n365 B.n140 163.367
R1137 B.n369 B.n140 163.367
R1138 B.n370 B.n369 163.367
R1139 B.n371 B.n370 163.367
R1140 B.n371 B.n138 163.367
R1141 B.n375 B.n138 163.367
R1142 B.n376 B.n375 163.367
R1143 B.n377 B.n376 163.367
R1144 B.n377 B.n136 163.367
R1145 B.n381 B.n136 163.367
R1146 B.n382 B.n381 163.367
R1147 B.n383 B.n382 163.367
R1148 B.n581 B.n580 163.367
R1149 B.n580 B.n579 163.367
R1150 B.n579 B.n70 163.367
R1151 B.n575 B.n70 163.367
R1152 B.n575 B.n574 163.367
R1153 B.n574 B.n573 163.367
R1154 B.n573 B.n72 163.367
R1155 B.n569 B.n72 163.367
R1156 B.n569 B.n568 163.367
R1157 B.n568 B.n567 163.367
R1158 B.n567 B.n74 163.367
R1159 B.n563 B.n74 163.367
R1160 B.n563 B.n562 163.367
R1161 B.n562 B.n561 163.367
R1162 B.n561 B.n76 163.367
R1163 B.n557 B.n76 163.367
R1164 B.n557 B.n556 163.367
R1165 B.n556 B.n555 163.367
R1166 B.n555 B.n78 163.367
R1167 B.n551 B.n78 163.367
R1168 B.n551 B.n550 163.367
R1169 B.n550 B.n549 163.367
R1170 B.n549 B.n80 163.367
R1171 B.n545 B.n80 163.367
R1172 B.n545 B.n544 163.367
R1173 B.n544 B.n543 163.367
R1174 B.n543 B.n82 163.367
R1175 B.n539 B.n82 163.367
R1176 B.n539 B.n538 163.367
R1177 B.n538 B.n537 163.367
R1178 B.n537 B.n84 163.367
R1179 B.n533 B.n84 163.367
R1180 B.n533 B.n532 163.367
R1181 B.n532 B.n531 163.367
R1182 B.n531 B.n86 163.367
R1183 B.n527 B.n86 163.367
R1184 B.n527 B.n526 163.367
R1185 B.n526 B.n525 163.367
R1186 B.n525 B.n88 163.367
R1187 B.n521 B.n88 163.367
R1188 B.n521 B.n520 163.367
R1189 B.n520 B.n519 163.367
R1190 B.n519 B.n90 163.367
R1191 B.n515 B.n90 163.367
R1192 B.n515 B.n514 163.367
R1193 B.n514 B.n513 163.367
R1194 B.n513 B.n92 163.367
R1195 B.n509 B.n92 163.367
R1196 B.n509 B.n508 163.367
R1197 B.n508 B.n507 163.367
R1198 B.n507 B.n94 163.367
R1199 B.n503 B.n94 163.367
R1200 B.n503 B.n502 163.367
R1201 B.n502 B.n501 163.367
R1202 B.n501 B.n96 163.367
R1203 B.n497 B.n96 163.367
R1204 B.n497 B.n496 163.367
R1205 B.n496 B.n495 163.367
R1206 B.n495 B.n98 163.367
R1207 B.n491 B.n98 163.367
R1208 B.n491 B.n490 163.367
R1209 B.n490 B.n489 163.367
R1210 B.n489 B.n100 163.367
R1211 B.n485 B.n100 163.367
R1212 B.n485 B.n484 163.367
R1213 B.n484 B.n483 163.367
R1214 B.n483 B.n102 163.367
R1215 B.n479 B.n102 163.367
R1216 B.n479 B.n478 163.367
R1217 B.n478 B.n477 163.367
R1218 B.n477 B.n104 163.367
R1219 B.n473 B.n104 163.367
R1220 B.n473 B.n472 163.367
R1221 B.n472 B.n471 163.367
R1222 B.n471 B.n106 163.367
R1223 B.n467 B.n106 163.367
R1224 B.n467 B.n466 163.367
R1225 B.n466 B.n465 163.367
R1226 B.n465 B.n108 163.367
R1227 B.n461 B.n108 163.367
R1228 B.n461 B.n460 163.367
R1229 B.n460 B.n459 163.367
R1230 B.n459 B.n110 163.367
R1231 B.n455 B.n110 163.367
R1232 B.n455 B.n454 163.367
R1233 B.n454 B.n453 163.367
R1234 B.n453 B.n112 163.367
R1235 B.n449 B.n112 163.367
R1236 B.n449 B.n448 163.367
R1237 B.n448 B.n447 163.367
R1238 B.n447 B.n114 163.367
R1239 B.n443 B.n114 163.367
R1240 B.n443 B.n442 163.367
R1241 B.n442 B.n441 163.367
R1242 B.n441 B.n116 163.367
R1243 B.n437 B.n116 163.367
R1244 B.n437 B.n436 163.367
R1245 B.n436 B.n435 163.367
R1246 B.n435 B.n118 163.367
R1247 B.n431 B.n118 163.367
R1248 B.n431 B.n430 163.367
R1249 B.n430 B.n429 163.367
R1250 B.n429 B.n120 163.367
R1251 B.n425 B.n120 163.367
R1252 B.n425 B.n424 163.367
R1253 B.n424 B.n423 163.367
R1254 B.n423 B.n122 163.367
R1255 B.n419 B.n122 163.367
R1256 B.n419 B.n418 163.367
R1257 B.n418 B.n417 163.367
R1258 B.n417 B.n124 163.367
R1259 B.n413 B.n124 163.367
R1260 B.n413 B.n412 163.367
R1261 B.n412 B.n411 163.367
R1262 B.n411 B.n126 163.367
R1263 B.n407 B.n126 163.367
R1264 B.n407 B.n406 163.367
R1265 B.n406 B.n405 163.367
R1266 B.n405 B.n128 163.367
R1267 B.n401 B.n128 163.367
R1268 B.n401 B.n400 163.367
R1269 B.n400 B.n399 163.367
R1270 B.n399 B.n130 163.367
R1271 B.n395 B.n130 163.367
R1272 B.n395 B.n394 163.367
R1273 B.n394 B.n393 163.367
R1274 B.n393 B.n132 163.367
R1275 B.n389 B.n132 163.367
R1276 B.n389 B.n388 163.367
R1277 B.n388 B.n387 163.367
R1278 B.n387 B.n134 163.367
R1279 B.n670 B.n35 163.367
R1280 B.n666 B.n35 163.367
R1281 B.n666 B.n665 163.367
R1282 B.n665 B.n664 163.367
R1283 B.n664 B.n37 163.367
R1284 B.n660 B.n37 163.367
R1285 B.n660 B.n659 163.367
R1286 B.n659 B.n658 163.367
R1287 B.n658 B.n39 163.367
R1288 B.n654 B.n39 163.367
R1289 B.n654 B.n653 163.367
R1290 B.n653 B.n652 163.367
R1291 B.n652 B.n41 163.367
R1292 B.n648 B.n41 163.367
R1293 B.n648 B.n647 163.367
R1294 B.n647 B.n646 163.367
R1295 B.n646 B.n43 163.367
R1296 B.n642 B.n43 163.367
R1297 B.n642 B.n641 163.367
R1298 B.n641 B.n640 163.367
R1299 B.n640 B.n45 163.367
R1300 B.n636 B.n45 163.367
R1301 B.n636 B.n635 163.367
R1302 B.n635 B.n634 163.367
R1303 B.n634 B.n47 163.367
R1304 B.n630 B.n47 163.367
R1305 B.n630 B.n629 163.367
R1306 B.n629 B.n628 163.367
R1307 B.n628 B.n52 163.367
R1308 B.n624 B.n52 163.367
R1309 B.n624 B.n623 163.367
R1310 B.n623 B.n622 163.367
R1311 B.n622 B.n54 163.367
R1312 B.n617 B.n54 163.367
R1313 B.n617 B.n616 163.367
R1314 B.n616 B.n615 163.367
R1315 B.n615 B.n58 163.367
R1316 B.n611 B.n58 163.367
R1317 B.n611 B.n610 163.367
R1318 B.n610 B.n609 163.367
R1319 B.n609 B.n60 163.367
R1320 B.n605 B.n60 163.367
R1321 B.n605 B.n604 163.367
R1322 B.n604 B.n603 163.367
R1323 B.n603 B.n62 163.367
R1324 B.n599 B.n62 163.367
R1325 B.n599 B.n598 163.367
R1326 B.n598 B.n597 163.367
R1327 B.n597 B.n64 163.367
R1328 B.n593 B.n64 163.367
R1329 B.n593 B.n592 163.367
R1330 B.n592 B.n591 163.367
R1331 B.n591 B.n66 163.367
R1332 B.n587 B.n66 163.367
R1333 B.n587 B.n586 163.367
R1334 B.n586 B.n585 163.367
R1335 B.n585 B.n68 163.367
R1336 B.n672 B.n671 163.367
R1337 B.n672 B.n33 163.367
R1338 B.n676 B.n33 163.367
R1339 B.n677 B.n676 163.367
R1340 B.n678 B.n677 163.367
R1341 B.n678 B.n31 163.367
R1342 B.n682 B.n31 163.367
R1343 B.n683 B.n682 163.367
R1344 B.n684 B.n683 163.367
R1345 B.n684 B.n29 163.367
R1346 B.n688 B.n29 163.367
R1347 B.n689 B.n688 163.367
R1348 B.n690 B.n689 163.367
R1349 B.n690 B.n27 163.367
R1350 B.n694 B.n27 163.367
R1351 B.n695 B.n694 163.367
R1352 B.n696 B.n695 163.367
R1353 B.n696 B.n25 163.367
R1354 B.n700 B.n25 163.367
R1355 B.n701 B.n700 163.367
R1356 B.n702 B.n701 163.367
R1357 B.n702 B.n23 163.367
R1358 B.n706 B.n23 163.367
R1359 B.n707 B.n706 163.367
R1360 B.n708 B.n707 163.367
R1361 B.n708 B.n21 163.367
R1362 B.n712 B.n21 163.367
R1363 B.n713 B.n712 163.367
R1364 B.n714 B.n713 163.367
R1365 B.n714 B.n19 163.367
R1366 B.n718 B.n19 163.367
R1367 B.n719 B.n718 163.367
R1368 B.n720 B.n719 163.367
R1369 B.n720 B.n17 163.367
R1370 B.n724 B.n17 163.367
R1371 B.n725 B.n724 163.367
R1372 B.n726 B.n725 163.367
R1373 B.n726 B.n15 163.367
R1374 B.n730 B.n15 163.367
R1375 B.n731 B.n730 163.367
R1376 B.n732 B.n731 163.367
R1377 B.n732 B.n13 163.367
R1378 B.n736 B.n13 163.367
R1379 B.n737 B.n736 163.367
R1380 B.n738 B.n737 163.367
R1381 B.n738 B.n11 163.367
R1382 B.n742 B.n11 163.367
R1383 B.n743 B.n742 163.367
R1384 B.n744 B.n743 163.367
R1385 B.n744 B.n9 163.367
R1386 B.n748 B.n9 163.367
R1387 B.n749 B.n748 163.367
R1388 B.n750 B.n749 163.367
R1389 B.n750 B.n7 163.367
R1390 B.n754 B.n7 163.367
R1391 B.n755 B.n754 163.367
R1392 B.n756 B.n755 163.367
R1393 B.n756 B.n5 163.367
R1394 B.n760 B.n5 163.367
R1395 B.n761 B.n760 163.367
R1396 B.n762 B.n761 163.367
R1397 B.n762 B.n3 163.367
R1398 B.n766 B.n3 163.367
R1399 B.n767 B.n766 163.367
R1400 B.n198 B.n2 163.367
R1401 B.n199 B.n198 163.367
R1402 B.n199 B.n196 163.367
R1403 B.n203 B.n196 163.367
R1404 B.n204 B.n203 163.367
R1405 B.n205 B.n204 163.367
R1406 B.n205 B.n194 163.367
R1407 B.n209 B.n194 163.367
R1408 B.n210 B.n209 163.367
R1409 B.n211 B.n210 163.367
R1410 B.n211 B.n192 163.367
R1411 B.n215 B.n192 163.367
R1412 B.n216 B.n215 163.367
R1413 B.n217 B.n216 163.367
R1414 B.n217 B.n190 163.367
R1415 B.n221 B.n190 163.367
R1416 B.n222 B.n221 163.367
R1417 B.n223 B.n222 163.367
R1418 B.n223 B.n188 163.367
R1419 B.n227 B.n188 163.367
R1420 B.n228 B.n227 163.367
R1421 B.n229 B.n228 163.367
R1422 B.n229 B.n186 163.367
R1423 B.n233 B.n186 163.367
R1424 B.n234 B.n233 163.367
R1425 B.n235 B.n234 163.367
R1426 B.n235 B.n184 163.367
R1427 B.n239 B.n184 163.367
R1428 B.n240 B.n239 163.367
R1429 B.n241 B.n240 163.367
R1430 B.n241 B.n182 163.367
R1431 B.n245 B.n182 163.367
R1432 B.n246 B.n245 163.367
R1433 B.n247 B.n246 163.367
R1434 B.n247 B.n180 163.367
R1435 B.n251 B.n180 163.367
R1436 B.n252 B.n251 163.367
R1437 B.n253 B.n252 163.367
R1438 B.n253 B.n178 163.367
R1439 B.n257 B.n178 163.367
R1440 B.n258 B.n257 163.367
R1441 B.n259 B.n258 163.367
R1442 B.n259 B.n176 163.367
R1443 B.n263 B.n176 163.367
R1444 B.n264 B.n263 163.367
R1445 B.n265 B.n264 163.367
R1446 B.n265 B.n174 163.367
R1447 B.n269 B.n174 163.367
R1448 B.n270 B.n269 163.367
R1449 B.n271 B.n270 163.367
R1450 B.n271 B.n172 163.367
R1451 B.n275 B.n172 163.367
R1452 B.n276 B.n275 163.367
R1453 B.n277 B.n276 163.367
R1454 B.n277 B.n170 163.367
R1455 B.n281 B.n170 163.367
R1456 B.n282 B.n281 163.367
R1457 B.n283 B.n282 163.367
R1458 B.n283 B.n168 163.367
R1459 B.n287 B.n168 163.367
R1460 B.n288 B.n287 163.367
R1461 B.n289 B.n288 163.367
R1462 B.n289 B.n166 163.367
R1463 B.n293 B.n166 163.367
R1464 B.n329 B.n328 76.0247
R1465 B.n148 B.n147 76.0247
R1466 B.n56 B.n55 76.0247
R1467 B.n49 B.n48 76.0247
R1468 B.n330 B.n329 59.5399
R1469 B.n348 B.n148 59.5399
R1470 B.n619 B.n56 59.5399
R1471 B.n50 B.n49 59.5399
R1472 B.n669 B.n34 33.5615
R1473 B.n583 B.n582 33.5615
R1474 B.n385 B.n384 33.5615
R1475 B.n292 B.n165 33.5615
R1476 B B.n769 18.0485
R1477 B.n673 B.n34 10.6151
R1478 B.n674 B.n673 10.6151
R1479 B.n675 B.n674 10.6151
R1480 B.n675 B.n32 10.6151
R1481 B.n679 B.n32 10.6151
R1482 B.n680 B.n679 10.6151
R1483 B.n681 B.n680 10.6151
R1484 B.n681 B.n30 10.6151
R1485 B.n685 B.n30 10.6151
R1486 B.n686 B.n685 10.6151
R1487 B.n687 B.n686 10.6151
R1488 B.n687 B.n28 10.6151
R1489 B.n691 B.n28 10.6151
R1490 B.n692 B.n691 10.6151
R1491 B.n693 B.n692 10.6151
R1492 B.n693 B.n26 10.6151
R1493 B.n697 B.n26 10.6151
R1494 B.n698 B.n697 10.6151
R1495 B.n699 B.n698 10.6151
R1496 B.n699 B.n24 10.6151
R1497 B.n703 B.n24 10.6151
R1498 B.n704 B.n703 10.6151
R1499 B.n705 B.n704 10.6151
R1500 B.n705 B.n22 10.6151
R1501 B.n709 B.n22 10.6151
R1502 B.n710 B.n709 10.6151
R1503 B.n711 B.n710 10.6151
R1504 B.n711 B.n20 10.6151
R1505 B.n715 B.n20 10.6151
R1506 B.n716 B.n715 10.6151
R1507 B.n717 B.n716 10.6151
R1508 B.n717 B.n18 10.6151
R1509 B.n721 B.n18 10.6151
R1510 B.n722 B.n721 10.6151
R1511 B.n723 B.n722 10.6151
R1512 B.n723 B.n16 10.6151
R1513 B.n727 B.n16 10.6151
R1514 B.n728 B.n727 10.6151
R1515 B.n729 B.n728 10.6151
R1516 B.n729 B.n14 10.6151
R1517 B.n733 B.n14 10.6151
R1518 B.n734 B.n733 10.6151
R1519 B.n735 B.n734 10.6151
R1520 B.n735 B.n12 10.6151
R1521 B.n739 B.n12 10.6151
R1522 B.n740 B.n739 10.6151
R1523 B.n741 B.n740 10.6151
R1524 B.n741 B.n10 10.6151
R1525 B.n745 B.n10 10.6151
R1526 B.n746 B.n745 10.6151
R1527 B.n747 B.n746 10.6151
R1528 B.n747 B.n8 10.6151
R1529 B.n751 B.n8 10.6151
R1530 B.n752 B.n751 10.6151
R1531 B.n753 B.n752 10.6151
R1532 B.n753 B.n6 10.6151
R1533 B.n757 B.n6 10.6151
R1534 B.n758 B.n757 10.6151
R1535 B.n759 B.n758 10.6151
R1536 B.n759 B.n4 10.6151
R1537 B.n763 B.n4 10.6151
R1538 B.n764 B.n763 10.6151
R1539 B.n765 B.n764 10.6151
R1540 B.n765 B.n0 10.6151
R1541 B.n669 B.n668 10.6151
R1542 B.n668 B.n667 10.6151
R1543 B.n667 B.n36 10.6151
R1544 B.n663 B.n36 10.6151
R1545 B.n663 B.n662 10.6151
R1546 B.n662 B.n661 10.6151
R1547 B.n661 B.n38 10.6151
R1548 B.n657 B.n38 10.6151
R1549 B.n657 B.n656 10.6151
R1550 B.n656 B.n655 10.6151
R1551 B.n655 B.n40 10.6151
R1552 B.n651 B.n40 10.6151
R1553 B.n651 B.n650 10.6151
R1554 B.n650 B.n649 10.6151
R1555 B.n649 B.n42 10.6151
R1556 B.n645 B.n42 10.6151
R1557 B.n645 B.n644 10.6151
R1558 B.n644 B.n643 10.6151
R1559 B.n643 B.n44 10.6151
R1560 B.n639 B.n44 10.6151
R1561 B.n639 B.n638 10.6151
R1562 B.n638 B.n637 10.6151
R1563 B.n637 B.n46 10.6151
R1564 B.n633 B.n632 10.6151
R1565 B.n632 B.n631 10.6151
R1566 B.n631 B.n51 10.6151
R1567 B.n627 B.n51 10.6151
R1568 B.n627 B.n626 10.6151
R1569 B.n626 B.n625 10.6151
R1570 B.n625 B.n53 10.6151
R1571 B.n621 B.n53 10.6151
R1572 B.n621 B.n620 10.6151
R1573 B.n618 B.n57 10.6151
R1574 B.n614 B.n57 10.6151
R1575 B.n614 B.n613 10.6151
R1576 B.n613 B.n612 10.6151
R1577 B.n612 B.n59 10.6151
R1578 B.n608 B.n59 10.6151
R1579 B.n608 B.n607 10.6151
R1580 B.n607 B.n606 10.6151
R1581 B.n606 B.n61 10.6151
R1582 B.n602 B.n61 10.6151
R1583 B.n602 B.n601 10.6151
R1584 B.n601 B.n600 10.6151
R1585 B.n600 B.n63 10.6151
R1586 B.n596 B.n63 10.6151
R1587 B.n596 B.n595 10.6151
R1588 B.n595 B.n594 10.6151
R1589 B.n594 B.n65 10.6151
R1590 B.n590 B.n65 10.6151
R1591 B.n590 B.n589 10.6151
R1592 B.n589 B.n588 10.6151
R1593 B.n588 B.n67 10.6151
R1594 B.n584 B.n67 10.6151
R1595 B.n584 B.n583 10.6151
R1596 B.n582 B.n69 10.6151
R1597 B.n578 B.n69 10.6151
R1598 B.n578 B.n577 10.6151
R1599 B.n577 B.n576 10.6151
R1600 B.n576 B.n71 10.6151
R1601 B.n572 B.n71 10.6151
R1602 B.n572 B.n571 10.6151
R1603 B.n571 B.n570 10.6151
R1604 B.n570 B.n73 10.6151
R1605 B.n566 B.n73 10.6151
R1606 B.n566 B.n565 10.6151
R1607 B.n565 B.n564 10.6151
R1608 B.n564 B.n75 10.6151
R1609 B.n560 B.n75 10.6151
R1610 B.n560 B.n559 10.6151
R1611 B.n559 B.n558 10.6151
R1612 B.n558 B.n77 10.6151
R1613 B.n554 B.n77 10.6151
R1614 B.n554 B.n553 10.6151
R1615 B.n553 B.n552 10.6151
R1616 B.n552 B.n79 10.6151
R1617 B.n548 B.n79 10.6151
R1618 B.n548 B.n547 10.6151
R1619 B.n547 B.n546 10.6151
R1620 B.n546 B.n81 10.6151
R1621 B.n542 B.n81 10.6151
R1622 B.n542 B.n541 10.6151
R1623 B.n541 B.n540 10.6151
R1624 B.n540 B.n83 10.6151
R1625 B.n536 B.n83 10.6151
R1626 B.n536 B.n535 10.6151
R1627 B.n535 B.n534 10.6151
R1628 B.n534 B.n85 10.6151
R1629 B.n530 B.n85 10.6151
R1630 B.n530 B.n529 10.6151
R1631 B.n529 B.n528 10.6151
R1632 B.n528 B.n87 10.6151
R1633 B.n524 B.n87 10.6151
R1634 B.n524 B.n523 10.6151
R1635 B.n523 B.n522 10.6151
R1636 B.n522 B.n89 10.6151
R1637 B.n518 B.n89 10.6151
R1638 B.n518 B.n517 10.6151
R1639 B.n517 B.n516 10.6151
R1640 B.n516 B.n91 10.6151
R1641 B.n512 B.n91 10.6151
R1642 B.n512 B.n511 10.6151
R1643 B.n511 B.n510 10.6151
R1644 B.n510 B.n93 10.6151
R1645 B.n506 B.n93 10.6151
R1646 B.n506 B.n505 10.6151
R1647 B.n505 B.n504 10.6151
R1648 B.n504 B.n95 10.6151
R1649 B.n500 B.n95 10.6151
R1650 B.n500 B.n499 10.6151
R1651 B.n499 B.n498 10.6151
R1652 B.n498 B.n97 10.6151
R1653 B.n494 B.n97 10.6151
R1654 B.n494 B.n493 10.6151
R1655 B.n493 B.n492 10.6151
R1656 B.n492 B.n99 10.6151
R1657 B.n488 B.n99 10.6151
R1658 B.n488 B.n487 10.6151
R1659 B.n487 B.n486 10.6151
R1660 B.n486 B.n101 10.6151
R1661 B.n482 B.n101 10.6151
R1662 B.n482 B.n481 10.6151
R1663 B.n481 B.n480 10.6151
R1664 B.n480 B.n103 10.6151
R1665 B.n476 B.n103 10.6151
R1666 B.n476 B.n475 10.6151
R1667 B.n475 B.n474 10.6151
R1668 B.n474 B.n105 10.6151
R1669 B.n470 B.n105 10.6151
R1670 B.n470 B.n469 10.6151
R1671 B.n469 B.n468 10.6151
R1672 B.n468 B.n107 10.6151
R1673 B.n464 B.n107 10.6151
R1674 B.n464 B.n463 10.6151
R1675 B.n463 B.n462 10.6151
R1676 B.n462 B.n109 10.6151
R1677 B.n458 B.n109 10.6151
R1678 B.n458 B.n457 10.6151
R1679 B.n457 B.n456 10.6151
R1680 B.n456 B.n111 10.6151
R1681 B.n452 B.n111 10.6151
R1682 B.n452 B.n451 10.6151
R1683 B.n451 B.n450 10.6151
R1684 B.n450 B.n113 10.6151
R1685 B.n446 B.n113 10.6151
R1686 B.n446 B.n445 10.6151
R1687 B.n445 B.n444 10.6151
R1688 B.n444 B.n115 10.6151
R1689 B.n440 B.n115 10.6151
R1690 B.n440 B.n439 10.6151
R1691 B.n439 B.n438 10.6151
R1692 B.n438 B.n117 10.6151
R1693 B.n434 B.n117 10.6151
R1694 B.n434 B.n433 10.6151
R1695 B.n433 B.n432 10.6151
R1696 B.n432 B.n119 10.6151
R1697 B.n428 B.n119 10.6151
R1698 B.n428 B.n427 10.6151
R1699 B.n427 B.n426 10.6151
R1700 B.n426 B.n121 10.6151
R1701 B.n422 B.n121 10.6151
R1702 B.n422 B.n421 10.6151
R1703 B.n421 B.n420 10.6151
R1704 B.n420 B.n123 10.6151
R1705 B.n416 B.n123 10.6151
R1706 B.n416 B.n415 10.6151
R1707 B.n415 B.n414 10.6151
R1708 B.n414 B.n125 10.6151
R1709 B.n410 B.n125 10.6151
R1710 B.n410 B.n409 10.6151
R1711 B.n409 B.n408 10.6151
R1712 B.n408 B.n127 10.6151
R1713 B.n404 B.n127 10.6151
R1714 B.n404 B.n403 10.6151
R1715 B.n403 B.n402 10.6151
R1716 B.n402 B.n129 10.6151
R1717 B.n398 B.n129 10.6151
R1718 B.n398 B.n397 10.6151
R1719 B.n397 B.n396 10.6151
R1720 B.n396 B.n131 10.6151
R1721 B.n392 B.n131 10.6151
R1722 B.n392 B.n391 10.6151
R1723 B.n391 B.n390 10.6151
R1724 B.n390 B.n133 10.6151
R1725 B.n386 B.n133 10.6151
R1726 B.n386 B.n385 10.6151
R1727 B.n197 B.n1 10.6151
R1728 B.n200 B.n197 10.6151
R1729 B.n201 B.n200 10.6151
R1730 B.n202 B.n201 10.6151
R1731 B.n202 B.n195 10.6151
R1732 B.n206 B.n195 10.6151
R1733 B.n207 B.n206 10.6151
R1734 B.n208 B.n207 10.6151
R1735 B.n208 B.n193 10.6151
R1736 B.n212 B.n193 10.6151
R1737 B.n213 B.n212 10.6151
R1738 B.n214 B.n213 10.6151
R1739 B.n214 B.n191 10.6151
R1740 B.n218 B.n191 10.6151
R1741 B.n219 B.n218 10.6151
R1742 B.n220 B.n219 10.6151
R1743 B.n220 B.n189 10.6151
R1744 B.n224 B.n189 10.6151
R1745 B.n225 B.n224 10.6151
R1746 B.n226 B.n225 10.6151
R1747 B.n226 B.n187 10.6151
R1748 B.n230 B.n187 10.6151
R1749 B.n231 B.n230 10.6151
R1750 B.n232 B.n231 10.6151
R1751 B.n232 B.n185 10.6151
R1752 B.n236 B.n185 10.6151
R1753 B.n237 B.n236 10.6151
R1754 B.n238 B.n237 10.6151
R1755 B.n238 B.n183 10.6151
R1756 B.n242 B.n183 10.6151
R1757 B.n243 B.n242 10.6151
R1758 B.n244 B.n243 10.6151
R1759 B.n244 B.n181 10.6151
R1760 B.n248 B.n181 10.6151
R1761 B.n249 B.n248 10.6151
R1762 B.n250 B.n249 10.6151
R1763 B.n250 B.n179 10.6151
R1764 B.n254 B.n179 10.6151
R1765 B.n255 B.n254 10.6151
R1766 B.n256 B.n255 10.6151
R1767 B.n256 B.n177 10.6151
R1768 B.n260 B.n177 10.6151
R1769 B.n261 B.n260 10.6151
R1770 B.n262 B.n261 10.6151
R1771 B.n262 B.n175 10.6151
R1772 B.n266 B.n175 10.6151
R1773 B.n267 B.n266 10.6151
R1774 B.n268 B.n267 10.6151
R1775 B.n268 B.n173 10.6151
R1776 B.n272 B.n173 10.6151
R1777 B.n273 B.n272 10.6151
R1778 B.n274 B.n273 10.6151
R1779 B.n274 B.n171 10.6151
R1780 B.n278 B.n171 10.6151
R1781 B.n279 B.n278 10.6151
R1782 B.n280 B.n279 10.6151
R1783 B.n280 B.n169 10.6151
R1784 B.n284 B.n169 10.6151
R1785 B.n285 B.n284 10.6151
R1786 B.n286 B.n285 10.6151
R1787 B.n286 B.n167 10.6151
R1788 B.n290 B.n167 10.6151
R1789 B.n291 B.n290 10.6151
R1790 B.n292 B.n291 10.6151
R1791 B.n296 B.n165 10.6151
R1792 B.n297 B.n296 10.6151
R1793 B.n298 B.n297 10.6151
R1794 B.n298 B.n163 10.6151
R1795 B.n302 B.n163 10.6151
R1796 B.n303 B.n302 10.6151
R1797 B.n304 B.n303 10.6151
R1798 B.n304 B.n161 10.6151
R1799 B.n308 B.n161 10.6151
R1800 B.n309 B.n308 10.6151
R1801 B.n310 B.n309 10.6151
R1802 B.n310 B.n159 10.6151
R1803 B.n314 B.n159 10.6151
R1804 B.n315 B.n314 10.6151
R1805 B.n316 B.n315 10.6151
R1806 B.n316 B.n157 10.6151
R1807 B.n320 B.n157 10.6151
R1808 B.n321 B.n320 10.6151
R1809 B.n322 B.n321 10.6151
R1810 B.n322 B.n155 10.6151
R1811 B.n326 B.n155 10.6151
R1812 B.n327 B.n326 10.6151
R1813 B.n331 B.n327 10.6151
R1814 B.n335 B.n153 10.6151
R1815 B.n336 B.n335 10.6151
R1816 B.n337 B.n336 10.6151
R1817 B.n337 B.n151 10.6151
R1818 B.n341 B.n151 10.6151
R1819 B.n342 B.n341 10.6151
R1820 B.n343 B.n342 10.6151
R1821 B.n343 B.n149 10.6151
R1822 B.n347 B.n149 10.6151
R1823 B.n350 B.n349 10.6151
R1824 B.n350 B.n145 10.6151
R1825 B.n354 B.n145 10.6151
R1826 B.n355 B.n354 10.6151
R1827 B.n356 B.n355 10.6151
R1828 B.n356 B.n143 10.6151
R1829 B.n360 B.n143 10.6151
R1830 B.n361 B.n360 10.6151
R1831 B.n362 B.n361 10.6151
R1832 B.n362 B.n141 10.6151
R1833 B.n366 B.n141 10.6151
R1834 B.n367 B.n366 10.6151
R1835 B.n368 B.n367 10.6151
R1836 B.n368 B.n139 10.6151
R1837 B.n372 B.n139 10.6151
R1838 B.n373 B.n372 10.6151
R1839 B.n374 B.n373 10.6151
R1840 B.n374 B.n137 10.6151
R1841 B.n378 B.n137 10.6151
R1842 B.n379 B.n378 10.6151
R1843 B.n380 B.n379 10.6151
R1844 B.n380 B.n135 10.6151
R1845 B.n384 B.n135 10.6151
R1846 B.n50 B.n46 9.36635
R1847 B.n619 B.n618 9.36635
R1848 B.n331 B.n330 9.36635
R1849 B.n349 B.n348 9.36635
R1850 B.n769 B.n0 8.11757
R1851 B.n769 B.n1 8.11757
R1852 B.n633 B.n50 1.24928
R1853 B.n620 B.n619 1.24928
R1854 B.n330 B.n153 1.24928
R1855 B.n348 B.n347 1.24928
C0 VN B 1.37977f
C1 VN VDD1 0.153658f
C2 B w_n4890_n2174# 9.97091f
C3 VDD1 w_n4890_n2174# 2.11523f
C4 VP B 2.45412f
C5 VP VDD1 5.31723f
C6 VTAIL B 3.3275f
C7 B VDD2 1.91822f
C8 VTAIL VDD1 6.77882f
C9 VDD1 VDD2 2.29169f
C10 VN w_n4890_n2174# 10.124901f
C11 VP VN 7.76987f
C12 VTAIL VN 6.08774f
C13 VN VDD2 4.84763f
C14 VP w_n4890_n2174# 10.7626f
C15 VTAIL w_n4890_n2174# 2.99481f
C16 VDD2 w_n4890_n2174# 2.27146f
C17 VP VTAIL 6.10185f
C18 VP VDD2 0.625158f
C19 VTAIL VDD2 6.83988f
C20 B VDD1 1.79104f
C21 VDD2 VSUBS 2.231621f
C22 VDD1 VSUBS 3.0638f
C23 VTAIL VSUBS 0.796423f
C24 VN VSUBS 7.842f
C25 VP VSUBS 4.143867f
C26 B VSUBS 5.603746f
C27 w_n4890_n2174# VSUBS 0.132675p
C28 B.n0 VSUBS 0.008127f
C29 B.n1 VSUBS 0.008127f
C30 B.n2 VSUBS 0.01202f
C31 B.n3 VSUBS 0.009211f
C32 B.n4 VSUBS 0.009211f
C33 B.n5 VSUBS 0.009211f
C34 B.n6 VSUBS 0.009211f
C35 B.n7 VSUBS 0.009211f
C36 B.n8 VSUBS 0.009211f
C37 B.n9 VSUBS 0.009211f
C38 B.n10 VSUBS 0.009211f
C39 B.n11 VSUBS 0.009211f
C40 B.n12 VSUBS 0.009211f
C41 B.n13 VSUBS 0.009211f
C42 B.n14 VSUBS 0.009211f
C43 B.n15 VSUBS 0.009211f
C44 B.n16 VSUBS 0.009211f
C45 B.n17 VSUBS 0.009211f
C46 B.n18 VSUBS 0.009211f
C47 B.n19 VSUBS 0.009211f
C48 B.n20 VSUBS 0.009211f
C49 B.n21 VSUBS 0.009211f
C50 B.n22 VSUBS 0.009211f
C51 B.n23 VSUBS 0.009211f
C52 B.n24 VSUBS 0.009211f
C53 B.n25 VSUBS 0.009211f
C54 B.n26 VSUBS 0.009211f
C55 B.n27 VSUBS 0.009211f
C56 B.n28 VSUBS 0.009211f
C57 B.n29 VSUBS 0.009211f
C58 B.n30 VSUBS 0.009211f
C59 B.n31 VSUBS 0.009211f
C60 B.n32 VSUBS 0.009211f
C61 B.n33 VSUBS 0.009211f
C62 B.n34 VSUBS 0.021079f
C63 B.n35 VSUBS 0.009211f
C64 B.n36 VSUBS 0.009211f
C65 B.n37 VSUBS 0.009211f
C66 B.n38 VSUBS 0.009211f
C67 B.n39 VSUBS 0.009211f
C68 B.n40 VSUBS 0.009211f
C69 B.n41 VSUBS 0.009211f
C70 B.n42 VSUBS 0.009211f
C71 B.n43 VSUBS 0.009211f
C72 B.n44 VSUBS 0.009211f
C73 B.n45 VSUBS 0.009211f
C74 B.n46 VSUBS 0.008669f
C75 B.n47 VSUBS 0.009211f
C76 B.t7 VSUBS 0.118541f
C77 B.t8 VSUBS 0.162364f
C78 B.t6 VSUBS 1.36623f
C79 B.n48 VSUBS 0.269055f
C80 B.n49 VSUBS 0.211896f
C81 B.n50 VSUBS 0.021341f
C82 B.n51 VSUBS 0.009211f
C83 B.n52 VSUBS 0.009211f
C84 B.n53 VSUBS 0.009211f
C85 B.n54 VSUBS 0.009211f
C86 B.t4 VSUBS 0.118543f
C87 B.t5 VSUBS 0.162366f
C88 B.t3 VSUBS 1.36623f
C89 B.n55 VSUBS 0.269053f
C90 B.n56 VSUBS 0.211894f
C91 B.n57 VSUBS 0.009211f
C92 B.n58 VSUBS 0.009211f
C93 B.n59 VSUBS 0.009211f
C94 B.n60 VSUBS 0.009211f
C95 B.n61 VSUBS 0.009211f
C96 B.n62 VSUBS 0.009211f
C97 B.n63 VSUBS 0.009211f
C98 B.n64 VSUBS 0.009211f
C99 B.n65 VSUBS 0.009211f
C100 B.n66 VSUBS 0.009211f
C101 B.n67 VSUBS 0.009211f
C102 B.n68 VSUBS 0.022809f
C103 B.n69 VSUBS 0.009211f
C104 B.n70 VSUBS 0.009211f
C105 B.n71 VSUBS 0.009211f
C106 B.n72 VSUBS 0.009211f
C107 B.n73 VSUBS 0.009211f
C108 B.n74 VSUBS 0.009211f
C109 B.n75 VSUBS 0.009211f
C110 B.n76 VSUBS 0.009211f
C111 B.n77 VSUBS 0.009211f
C112 B.n78 VSUBS 0.009211f
C113 B.n79 VSUBS 0.009211f
C114 B.n80 VSUBS 0.009211f
C115 B.n81 VSUBS 0.009211f
C116 B.n82 VSUBS 0.009211f
C117 B.n83 VSUBS 0.009211f
C118 B.n84 VSUBS 0.009211f
C119 B.n85 VSUBS 0.009211f
C120 B.n86 VSUBS 0.009211f
C121 B.n87 VSUBS 0.009211f
C122 B.n88 VSUBS 0.009211f
C123 B.n89 VSUBS 0.009211f
C124 B.n90 VSUBS 0.009211f
C125 B.n91 VSUBS 0.009211f
C126 B.n92 VSUBS 0.009211f
C127 B.n93 VSUBS 0.009211f
C128 B.n94 VSUBS 0.009211f
C129 B.n95 VSUBS 0.009211f
C130 B.n96 VSUBS 0.009211f
C131 B.n97 VSUBS 0.009211f
C132 B.n98 VSUBS 0.009211f
C133 B.n99 VSUBS 0.009211f
C134 B.n100 VSUBS 0.009211f
C135 B.n101 VSUBS 0.009211f
C136 B.n102 VSUBS 0.009211f
C137 B.n103 VSUBS 0.009211f
C138 B.n104 VSUBS 0.009211f
C139 B.n105 VSUBS 0.009211f
C140 B.n106 VSUBS 0.009211f
C141 B.n107 VSUBS 0.009211f
C142 B.n108 VSUBS 0.009211f
C143 B.n109 VSUBS 0.009211f
C144 B.n110 VSUBS 0.009211f
C145 B.n111 VSUBS 0.009211f
C146 B.n112 VSUBS 0.009211f
C147 B.n113 VSUBS 0.009211f
C148 B.n114 VSUBS 0.009211f
C149 B.n115 VSUBS 0.009211f
C150 B.n116 VSUBS 0.009211f
C151 B.n117 VSUBS 0.009211f
C152 B.n118 VSUBS 0.009211f
C153 B.n119 VSUBS 0.009211f
C154 B.n120 VSUBS 0.009211f
C155 B.n121 VSUBS 0.009211f
C156 B.n122 VSUBS 0.009211f
C157 B.n123 VSUBS 0.009211f
C158 B.n124 VSUBS 0.009211f
C159 B.n125 VSUBS 0.009211f
C160 B.n126 VSUBS 0.009211f
C161 B.n127 VSUBS 0.009211f
C162 B.n128 VSUBS 0.009211f
C163 B.n129 VSUBS 0.009211f
C164 B.n130 VSUBS 0.009211f
C165 B.n131 VSUBS 0.009211f
C166 B.n132 VSUBS 0.009211f
C167 B.n133 VSUBS 0.009211f
C168 B.n134 VSUBS 0.021079f
C169 B.n135 VSUBS 0.009211f
C170 B.n136 VSUBS 0.009211f
C171 B.n137 VSUBS 0.009211f
C172 B.n138 VSUBS 0.009211f
C173 B.n139 VSUBS 0.009211f
C174 B.n140 VSUBS 0.009211f
C175 B.n141 VSUBS 0.009211f
C176 B.n142 VSUBS 0.009211f
C177 B.n143 VSUBS 0.009211f
C178 B.n144 VSUBS 0.009211f
C179 B.n145 VSUBS 0.009211f
C180 B.n146 VSUBS 0.009211f
C181 B.t2 VSUBS 0.118543f
C182 B.t1 VSUBS 0.162366f
C183 B.t0 VSUBS 1.36623f
C184 B.n147 VSUBS 0.269053f
C185 B.n148 VSUBS 0.211894f
C186 B.n149 VSUBS 0.009211f
C187 B.n150 VSUBS 0.009211f
C188 B.n151 VSUBS 0.009211f
C189 B.n152 VSUBS 0.009211f
C190 B.n153 VSUBS 0.005147f
C191 B.n154 VSUBS 0.009211f
C192 B.n155 VSUBS 0.009211f
C193 B.n156 VSUBS 0.009211f
C194 B.n157 VSUBS 0.009211f
C195 B.n158 VSUBS 0.009211f
C196 B.n159 VSUBS 0.009211f
C197 B.n160 VSUBS 0.009211f
C198 B.n161 VSUBS 0.009211f
C199 B.n162 VSUBS 0.009211f
C200 B.n163 VSUBS 0.009211f
C201 B.n164 VSUBS 0.009211f
C202 B.n165 VSUBS 0.022809f
C203 B.n166 VSUBS 0.009211f
C204 B.n167 VSUBS 0.009211f
C205 B.n168 VSUBS 0.009211f
C206 B.n169 VSUBS 0.009211f
C207 B.n170 VSUBS 0.009211f
C208 B.n171 VSUBS 0.009211f
C209 B.n172 VSUBS 0.009211f
C210 B.n173 VSUBS 0.009211f
C211 B.n174 VSUBS 0.009211f
C212 B.n175 VSUBS 0.009211f
C213 B.n176 VSUBS 0.009211f
C214 B.n177 VSUBS 0.009211f
C215 B.n178 VSUBS 0.009211f
C216 B.n179 VSUBS 0.009211f
C217 B.n180 VSUBS 0.009211f
C218 B.n181 VSUBS 0.009211f
C219 B.n182 VSUBS 0.009211f
C220 B.n183 VSUBS 0.009211f
C221 B.n184 VSUBS 0.009211f
C222 B.n185 VSUBS 0.009211f
C223 B.n186 VSUBS 0.009211f
C224 B.n187 VSUBS 0.009211f
C225 B.n188 VSUBS 0.009211f
C226 B.n189 VSUBS 0.009211f
C227 B.n190 VSUBS 0.009211f
C228 B.n191 VSUBS 0.009211f
C229 B.n192 VSUBS 0.009211f
C230 B.n193 VSUBS 0.009211f
C231 B.n194 VSUBS 0.009211f
C232 B.n195 VSUBS 0.009211f
C233 B.n196 VSUBS 0.009211f
C234 B.n197 VSUBS 0.009211f
C235 B.n198 VSUBS 0.009211f
C236 B.n199 VSUBS 0.009211f
C237 B.n200 VSUBS 0.009211f
C238 B.n201 VSUBS 0.009211f
C239 B.n202 VSUBS 0.009211f
C240 B.n203 VSUBS 0.009211f
C241 B.n204 VSUBS 0.009211f
C242 B.n205 VSUBS 0.009211f
C243 B.n206 VSUBS 0.009211f
C244 B.n207 VSUBS 0.009211f
C245 B.n208 VSUBS 0.009211f
C246 B.n209 VSUBS 0.009211f
C247 B.n210 VSUBS 0.009211f
C248 B.n211 VSUBS 0.009211f
C249 B.n212 VSUBS 0.009211f
C250 B.n213 VSUBS 0.009211f
C251 B.n214 VSUBS 0.009211f
C252 B.n215 VSUBS 0.009211f
C253 B.n216 VSUBS 0.009211f
C254 B.n217 VSUBS 0.009211f
C255 B.n218 VSUBS 0.009211f
C256 B.n219 VSUBS 0.009211f
C257 B.n220 VSUBS 0.009211f
C258 B.n221 VSUBS 0.009211f
C259 B.n222 VSUBS 0.009211f
C260 B.n223 VSUBS 0.009211f
C261 B.n224 VSUBS 0.009211f
C262 B.n225 VSUBS 0.009211f
C263 B.n226 VSUBS 0.009211f
C264 B.n227 VSUBS 0.009211f
C265 B.n228 VSUBS 0.009211f
C266 B.n229 VSUBS 0.009211f
C267 B.n230 VSUBS 0.009211f
C268 B.n231 VSUBS 0.009211f
C269 B.n232 VSUBS 0.009211f
C270 B.n233 VSUBS 0.009211f
C271 B.n234 VSUBS 0.009211f
C272 B.n235 VSUBS 0.009211f
C273 B.n236 VSUBS 0.009211f
C274 B.n237 VSUBS 0.009211f
C275 B.n238 VSUBS 0.009211f
C276 B.n239 VSUBS 0.009211f
C277 B.n240 VSUBS 0.009211f
C278 B.n241 VSUBS 0.009211f
C279 B.n242 VSUBS 0.009211f
C280 B.n243 VSUBS 0.009211f
C281 B.n244 VSUBS 0.009211f
C282 B.n245 VSUBS 0.009211f
C283 B.n246 VSUBS 0.009211f
C284 B.n247 VSUBS 0.009211f
C285 B.n248 VSUBS 0.009211f
C286 B.n249 VSUBS 0.009211f
C287 B.n250 VSUBS 0.009211f
C288 B.n251 VSUBS 0.009211f
C289 B.n252 VSUBS 0.009211f
C290 B.n253 VSUBS 0.009211f
C291 B.n254 VSUBS 0.009211f
C292 B.n255 VSUBS 0.009211f
C293 B.n256 VSUBS 0.009211f
C294 B.n257 VSUBS 0.009211f
C295 B.n258 VSUBS 0.009211f
C296 B.n259 VSUBS 0.009211f
C297 B.n260 VSUBS 0.009211f
C298 B.n261 VSUBS 0.009211f
C299 B.n262 VSUBS 0.009211f
C300 B.n263 VSUBS 0.009211f
C301 B.n264 VSUBS 0.009211f
C302 B.n265 VSUBS 0.009211f
C303 B.n266 VSUBS 0.009211f
C304 B.n267 VSUBS 0.009211f
C305 B.n268 VSUBS 0.009211f
C306 B.n269 VSUBS 0.009211f
C307 B.n270 VSUBS 0.009211f
C308 B.n271 VSUBS 0.009211f
C309 B.n272 VSUBS 0.009211f
C310 B.n273 VSUBS 0.009211f
C311 B.n274 VSUBS 0.009211f
C312 B.n275 VSUBS 0.009211f
C313 B.n276 VSUBS 0.009211f
C314 B.n277 VSUBS 0.009211f
C315 B.n278 VSUBS 0.009211f
C316 B.n279 VSUBS 0.009211f
C317 B.n280 VSUBS 0.009211f
C318 B.n281 VSUBS 0.009211f
C319 B.n282 VSUBS 0.009211f
C320 B.n283 VSUBS 0.009211f
C321 B.n284 VSUBS 0.009211f
C322 B.n285 VSUBS 0.009211f
C323 B.n286 VSUBS 0.009211f
C324 B.n287 VSUBS 0.009211f
C325 B.n288 VSUBS 0.009211f
C326 B.n289 VSUBS 0.009211f
C327 B.n290 VSUBS 0.009211f
C328 B.n291 VSUBS 0.009211f
C329 B.n292 VSUBS 0.021079f
C330 B.n293 VSUBS 0.021079f
C331 B.n294 VSUBS 0.022809f
C332 B.n295 VSUBS 0.009211f
C333 B.n296 VSUBS 0.009211f
C334 B.n297 VSUBS 0.009211f
C335 B.n298 VSUBS 0.009211f
C336 B.n299 VSUBS 0.009211f
C337 B.n300 VSUBS 0.009211f
C338 B.n301 VSUBS 0.009211f
C339 B.n302 VSUBS 0.009211f
C340 B.n303 VSUBS 0.009211f
C341 B.n304 VSUBS 0.009211f
C342 B.n305 VSUBS 0.009211f
C343 B.n306 VSUBS 0.009211f
C344 B.n307 VSUBS 0.009211f
C345 B.n308 VSUBS 0.009211f
C346 B.n309 VSUBS 0.009211f
C347 B.n310 VSUBS 0.009211f
C348 B.n311 VSUBS 0.009211f
C349 B.n312 VSUBS 0.009211f
C350 B.n313 VSUBS 0.009211f
C351 B.n314 VSUBS 0.009211f
C352 B.n315 VSUBS 0.009211f
C353 B.n316 VSUBS 0.009211f
C354 B.n317 VSUBS 0.009211f
C355 B.n318 VSUBS 0.009211f
C356 B.n319 VSUBS 0.009211f
C357 B.n320 VSUBS 0.009211f
C358 B.n321 VSUBS 0.009211f
C359 B.n322 VSUBS 0.009211f
C360 B.n323 VSUBS 0.009211f
C361 B.n324 VSUBS 0.009211f
C362 B.n325 VSUBS 0.009211f
C363 B.n326 VSUBS 0.009211f
C364 B.n327 VSUBS 0.009211f
C365 B.t11 VSUBS 0.118541f
C366 B.t10 VSUBS 0.162364f
C367 B.t9 VSUBS 1.36623f
C368 B.n328 VSUBS 0.269055f
C369 B.n329 VSUBS 0.211896f
C370 B.n330 VSUBS 0.021341f
C371 B.n331 VSUBS 0.008669f
C372 B.n332 VSUBS 0.009211f
C373 B.n333 VSUBS 0.009211f
C374 B.n334 VSUBS 0.009211f
C375 B.n335 VSUBS 0.009211f
C376 B.n336 VSUBS 0.009211f
C377 B.n337 VSUBS 0.009211f
C378 B.n338 VSUBS 0.009211f
C379 B.n339 VSUBS 0.009211f
C380 B.n340 VSUBS 0.009211f
C381 B.n341 VSUBS 0.009211f
C382 B.n342 VSUBS 0.009211f
C383 B.n343 VSUBS 0.009211f
C384 B.n344 VSUBS 0.009211f
C385 B.n345 VSUBS 0.009211f
C386 B.n346 VSUBS 0.009211f
C387 B.n347 VSUBS 0.005147f
C388 B.n348 VSUBS 0.021341f
C389 B.n349 VSUBS 0.008669f
C390 B.n350 VSUBS 0.009211f
C391 B.n351 VSUBS 0.009211f
C392 B.n352 VSUBS 0.009211f
C393 B.n353 VSUBS 0.009211f
C394 B.n354 VSUBS 0.009211f
C395 B.n355 VSUBS 0.009211f
C396 B.n356 VSUBS 0.009211f
C397 B.n357 VSUBS 0.009211f
C398 B.n358 VSUBS 0.009211f
C399 B.n359 VSUBS 0.009211f
C400 B.n360 VSUBS 0.009211f
C401 B.n361 VSUBS 0.009211f
C402 B.n362 VSUBS 0.009211f
C403 B.n363 VSUBS 0.009211f
C404 B.n364 VSUBS 0.009211f
C405 B.n365 VSUBS 0.009211f
C406 B.n366 VSUBS 0.009211f
C407 B.n367 VSUBS 0.009211f
C408 B.n368 VSUBS 0.009211f
C409 B.n369 VSUBS 0.009211f
C410 B.n370 VSUBS 0.009211f
C411 B.n371 VSUBS 0.009211f
C412 B.n372 VSUBS 0.009211f
C413 B.n373 VSUBS 0.009211f
C414 B.n374 VSUBS 0.009211f
C415 B.n375 VSUBS 0.009211f
C416 B.n376 VSUBS 0.009211f
C417 B.n377 VSUBS 0.009211f
C418 B.n378 VSUBS 0.009211f
C419 B.n379 VSUBS 0.009211f
C420 B.n380 VSUBS 0.009211f
C421 B.n381 VSUBS 0.009211f
C422 B.n382 VSUBS 0.009211f
C423 B.n383 VSUBS 0.022809f
C424 B.n384 VSUBS 0.02175f
C425 B.n385 VSUBS 0.022138f
C426 B.n386 VSUBS 0.009211f
C427 B.n387 VSUBS 0.009211f
C428 B.n388 VSUBS 0.009211f
C429 B.n389 VSUBS 0.009211f
C430 B.n390 VSUBS 0.009211f
C431 B.n391 VSUBS 0.009211f
C432 B.n392 VSUBS 0.009211f
C433 B.n393 VSUBS 0.009211f
C434 B.n394 VSUBS 0.009211f
C435 B.n395 VSUBS 0.009211f
C436 B.n396 VSUBS 0.009211f
C437 B.n397 VSUBS 0.009211f
C438 B.n398 VSUBS 0.009211f
C439 B.n399 VSUBS 0.009211f
C440 B.n400 VSUBS 0.009211f
C441 B.n401 VSUBS 0.009211f
C442 B.n402 VSUBS 0.009211f
C443 B.n403 VSUBS 0.009211f
C444 B.n404 VSUBS 0.009211f
C445 B.n405 VSUBS 0.009211f
C446 B.n406 VSUBS 0.009211f
C447 B.n407 VSUBS 0.009211f
C448 B.n408 VSUBS 0.009211f
C449 B.n409 VSUBS 0.009211f
C450 B.n410 VSUBS 0.009211f
C451 B.n411 VSUBS 0.009211f
C452 B.n412 VSUBS 0.009211f
C453 B.n413 VSUBS 0.009211f
C454 B.n414 VSUBS 0.009211f
C455 B.n415 VSUBS 0.009211f
C456 B.n416 VSUBS 0.009211f
C457 B.n417 VSUBS 0.009211f
C458 B.n418 VSUBS 0.009211f
C459 B.n419 VSUBS 0.009211f
C460 B.n420 VSUBS 0.009211f
C461 B.n421 VSUBS 0.009211f
C462 B.n422 VSUBS 0.009211f
C463 B.n423 VSUBS 0.009211f
C464 B.n424 VSUBS 0.009211f
C465 B.n425 VSUBS 0.009211f
C466 B.n426 VSUBS 0.009211f
C467 B.n427 VSUBS 0.009211f
C468 B.n428 VSUBS 0.009211f
C469 B.n429 VSUBS 0.009211f
C470 B.n430 VSUBS 0.009211f
C471 B.n431 VSUBS 0.009211f
C472 B.n432 VSUBS 0.009211f
C473 B.n433 VSUBS 0.009211f
C474 B.n434 VSUBS 0.009211f
C475 B.n435 VSUBS 0.009211f
C476 B.n436 VSUBS 0.009211f
C477 B.n437 VSUBS 0.009211f
C478 B.n438 VSUBS 0.009211f
C479 B.n439 VSUBS 0.009211f
C480 B.n440 VSUBS 0.009211f
C481 B.n441 VSUBS 0.009211f
C482 B.n442 VSUBS 0.009211f
C483 B.n443 VSUBS 0.009211f
C484 B.n444 VSUBS 0.009211f
C485 B.n445 VSUBS 0.009211f
C486 B.n446 VSUBS 0.009211f
C487 B.n447 VSUBS 0.009211f
C488 B.n448 VSUBS 0.009211f
C489 B.n449 VSUBS 0.009211f
C490 B.n450 VSUBS 0.009211f
C491 B.n451 VSUBS 0.009211f
C492 B.n452 VSUBS 0.009211f
C493 B.n453 VSUBS 0.009211f
C494 B.n454 VSUBS 0.009211f
C495 B.n455 VSUBS 0.009211f
C496 B.n456 VSUBS 0.009211f
C497 B.n457 VSUBS 0.009211f
C498 B.n458 VSUBS 0.009211f
C499 B.n459 VSUBS 0.009211f
C500 B.n460 VSUBS 0.009211f
C501 B.n461 VSUBS 0.009211f
C502 B.n462 VSUBS 0.009211f
C503 B.n463 VSUBS 0.009211f
C504 B.n464 VSUBS 0.009211f
C505 B.n465 VSUBS 0.009211f
C506 B.n466 VSUBS 0.009211f
C507 B.n467 VSUBS 0.009211f
C508 B.n468 VSUBS 0.009211f
C509 B.n469 VSUBS 0.009211f
C510 B.n470 VSUBS 0.009211f
C511 B.n471 VSUBS 0.009211f
C512 B.n472 VSUBS 0.009211f
C513 B.n473 VSUBS 0.009211f
C514 B.n474 VSUBS 0.009211f
C515 B.n475 VSUBS 0.009211f
C516 B.n476 VSUBS 0.009211f
C517 B.n477 VSUBS 0.009211f
C518 B.n478 VSUBS 0.009211f
C519 B.n479 VSUBS 0.009211f
C520 B.n480 VSUBS 0.009211f
C521 B.n481 VSUBS 0.009211f
C522 B.n482 VSUBS 0.009211f
C523 B.n483 VSUBS 0.009211f
C524 B.n484 VSUBS 0.009211f
C525 B.n485 VSUBS 0.009211f
C526 B.n486 VSUBS 0.009211f
C527 B.n487 VSUBS 0.009211f
C528 B.n488 VSUBS 0.009211f
C529 B.n489 VSUBS 0.009211f
C530 B.n490 VSUBS 0.009211f
C531 B.n491 VSUBS 0.009211f
C532 B.n492 VSUBS 0.009211f
C533 B.n493 VSUBS 0.009211f
C534 B.n494 VSUBS 0.009211f
C535 B.n495 VSUBS 0.009211f
C536 B.n496 VSUBS 0.009211f
C537 B.n497 VSUBS 0.009211f
C538 B.n498 VSUBS 0.009211f
C539 B.n499 VSUBS 0.009211f
C540 B.n500 VSUBS 0.009211f
C541 B.n501 VSUBS 0.009211f
C542 B.n502 VSUBS 0.009211f
C543 B.n503 VSUBS 0.009211f
C544 B.n504 VSUBS 0.009211f
C545 B.n505 VSUBS 0.009211f
C546 B.n506 VSUBS 0.009211f
C547 B.n507 VSUBS 0.009211f
C548 B.n508 VSUBS 0.009211f
C549 B.n509 VSUBS 0.009211f
C550 B.n510 VSUBS 0.009211f
C551 B.n511 VSUBS 0.009211f
C552 B.n512 VSUBS 0.009211f
C553 B.n513 VSUBS 0.009211f
C554 B.n514 VSUBS 0.009211f
C555 B.n515 VSUBS 0.009211f
C556 B.n516 VSUBS 0.009211f
C557 B.n517 VSUBS 0.009211f
C558 B.n518 VSUBS 0.009211f
C559 B.n519 VSUBS 0.009211f
C560 B.n520 VSUBS 0.009211f
C561 B.n521 VSUBS 0.009211f
C562 B.n522 VSUBS 0.009211f
C563 B.n523 VSUBS 0.009211f
C564 B.n524 VSUBS 0.009211f
C565 B.n525 VSUBS 0.009211f
C566 B.n526 VSUBS 0.009211f
C567 B.n527 VSUBS 0.009211f
C568 B.n528 VSUBS 0.009211f
C569 B.n529 VSUBS 0.009211f
C570 B.n530 VSUBS 0.009211f
C571 B.n531 VSUBS 0.009211f
C572 B.n532 VSUBS 0.009211f
C573 B.n533 VSUBS 0.009211f
C574 B.n534 VSUBS 0.009211f
C575 B.n535 VSUBS 0.009211f
C576 B.n536 VSUBS 0.009211f
C577 B.n537 VSUBS 0.009211f
C578 B.n538 VSUBS 0.009211f
C579 B.n539 VSUBS 0.009211f
C580 B.n540 VSUBS 0.009211f
C581 B.n541 VSUBS 0.009211f
C582 B.n542 VSUBS 0.009211f
C583 B.n543 VSUBS 0.009211f
C584 B.n544 VSUBS 0.009211f
C585 B.n545 VSUBS 0.009211f
C586 B.n546 VSUBS 0.009211f
C587 B.n547 VSUBS 0.009211f
C588 B.n548 VSUBS 0.009211f
C589 B.n549 VSUBS 0.009211f
C590 B.n550 VSUBS 0.009211f
C591 B.n551 VSUBS 0.009211f
C592 B.n552 VSUBS 0.009211f
C593 B.n553 VSUBS 0.009211f
C594 B.n554 VSUBS 0.009211f
C595 B.n555 VSUBS 0.009211f
C596 B.n556 VSUBS 0.009211f
C597 B.n557 VSUBS 0.009211f
C598 B.n558 VSUBS 0.009211f
C599 B.n559 VSUBS 0.009211f
C600 B.n560 VSUBS 0.009211f
C601 B.n561 VSUBS 0.009211f
C602 B.n562 VSUBS 0.009211f
C603 B.n563 VSUBS 0.009211f
C604 B.n564 VSUBS 0.009211f
C605 B.n565 VSUBS 0.009211f
C606 B.n566 VSUBS 0.009211f
C607 B.n567 VSUBS 0.009211f
C608 B.n568 VSUBS 0.009211f
C609 B.n569 VSUBS 0.009211f
C610 B.n570 VSUBS 0.009211f
C611 B.n571 VSUBS 0.009211f
C612 B.n572 VSUBS 0.009211f
C613 B.n573 VSUBS 0.009211f
C614 B.n574 VSUBS 0.009211f
C615 B.n575 VSUBS 0.009211f
C616 B.n576 VSUBS 0.009211f
C617 B.n577 VSUBS 0.009211f
C618 B.n578 VSUBS 0.009211f
C619 B.n579 VSUBS 0.009211f
C620 B.n580 VSUBS 0.009211f
C621 B.n581 VSUBS 0.021079f
C622 B.n582 VSUBS 0.021079f
C623 B.n583 VSUBS 0.022809f
C624 B.n584 VSUBS 0.009211f
C625 B.n585 VSUBS 0.009211f
C626 B.n586 VSUBS 0.009211f
C627 B.n587 VSUBS 0.009211f
C628 B.n588 VSUBS 0.009211f
C629 B.n589 VSUBS 0.009211f
C630 B.n590 VSUBS 0.009211f
C631 B.n591 VSUBS 0.009211f
C632 B.n592 VSUBS 0.009211f
C633 B.n593 VSUBS 0.009211f
C634 B.n594 VSUBS 0.009211f
C635 B.n595 VSUBS 0.009211f
C636 B.n596 VSUBS 0.009211f
C637 B.n597 VSUBS 0.009211f
C638 B.n598 VSUBS 0.009211f
C639 B.n599 VSUBS 0.009211f
C640 B.n600 VSUBS 0.009211f
C641 B.n601 VSUBS 0.009211f
C642 B.n602 VSUBS 0.009211f
C643 B.n603 VSUBS 0.009211f
C644 B.n604 VSUBS 0.009211f
C645 B.n605 VSUBS 0.009211f
C646 B.n606 VSUBS 0.009211f
C647 B.n607 VSUBS 0.009211f
C648 B.n608 VSUBS 0.009211f
C649 B.n609 VSUBS 0.009211f
C650 B.n610 VSUBS 0.009211f
C651 B.n611 VSUBS 0.009211f
C652 B.n612 VSUBS 0.009211f
C653 B.n613 VSUBS 0.009211f
C654 B.n614 VSUBS 0.009211f
C655 B.n615 VSUBS 0.009211f
C656 B.n616 VSUBS 0.009211f
C657 B.n617 VSUBS 0.009211f
C658 B.n618 VSUBS 0.008669f
C659 B.n619 VSUBS 0.021341f
C660 B.n620 VSUBS 0.005147f
C661 B.n621 VSUBS 0.009211f
C662 B.n622 VSUBS 0.009211f
C663 B.n623 VSUBS 0.009211f
C664 B.n624 VSUBS 0.009211f
C665 B.n625 VSUBS 0.009211f
C666 B.n626 VSUBS 0.009211f
C667 B.n627 VSUBS 0.009211f
C668 B.n628 VSUBS 0.009211f
C669 B.n629 VSUBS 0.009211f
C670 B.n630 VSUBS 0.009211f
C671 B.n631 VSUBS 0.009211f
C672 B.n632 VSUBS 0.009211f
C673 B.n633 VSUBS 0.005147f
C674 B.n634 VSUBS 0.009211f
C675 B.n635 VSUBS 0.009211f
C676 B.n636 VSUBS 0.009211f
C677 B.n637 VSUBS 0.009211f
C678 B.n638 VSUBS 0.009211f
C679 B.n639 VSUBS 0.009211f
C680 B.n640 VSUBS 0.009211f
C681 B.n641 VSUBS 0.009211f
C682 B.n642 VSUBS 0.009211f
C683 B.n643 VSUBS 0.009211f
C684 B.n644 VSUBS 0.009211f
C685 B.n645 VSUBS 0.009211f
C686 B.n646 VSUBS 0.009211f
C687 B.n647 VSUBS 0.009211f
C688 B.n648 VSUBS 0.009211f
C689 B.n649 VSUBS 0.009211f
C690 B.n650 VSUBS 0.009211f
C691 B.n651 VSUBS 0.009211f
C692 B.n652 VSUBS 0.009211f
C693 B.n653 VSUBS 0.009211f
C694 B.n654 VSUBS 0.009211f
C695 B.n655 VSUBS 0.009211f
C696 B.n656 VSUBS 0.009211f
C697 B.n657 VSUBS 0.009211f
C698 B.n658 VSUBS 0.009211f
C699 B.n659 VSUBS 0.009211f
C700 B.n660 VSUBS 0.009211f
C701 B.n661 VSUBS 0.009211f
C702 B.n662 VSUBS 0.009211f
C703 B.n663 VSUBS 0.009211f
C704 B.n664 VSUBS 0.009211f
C705 B.n665 VSUBS 0.009211f
C706 B.n666 VSUBS 0.009211f
C707 B.n667 VSUBS 0.009211f
C708 B.n668 VSUBS 0.009211f
C709 B.n669 VSUBS 0.022809f
C710 B.n670 VSUBS 0.022809f
C711 B.n671 VSUBS 0.021079f
C712 B.n672 VSUBS 0.009211f
C713 B.n673 VSUBS 0.009211f
C714 B.n674 VSUBS 0.009211f
C715 B.n675 VSUBS 0.009211f
C716 B.n676 VSUBS 0.009211f
C717 B.n677 VSUBS 0.009211f
C718 B.n678 VSUBS 0.009211f
C719 B.n679 VSUBS 0.009211f
C720 B.n680 VSUBS 0.009211f
C721 B.n681 VSUBS 0.009211f
C722 B.n682 VSUBS 0.009211f
C723 B.n683 VSUBS 0.009211f
C724 B.n684 VSUBS 0.009211f
C725 B.n685 VSUBS 0.009211f
C726 B.n686 VSUBS 0.009211f
C727 B.n687 VSUBS 0.009211f
C728 B.n688 VSUBS 0.009211f
C729 B.n689 VSUBS 0.009211f
C730 B.n690 VSUBS 0.009211f
C731 B.n691 VSUBS 0.009211f
C732 B.n692 VSUBS 0.009211f
C733 B.n693 VSUBS 0.009211f
C734 B.n694 VSUBS 0.009211f
C735 B.n695 VSUBS 0.009211f
C736 B.n696 VSUBS 0.009211f
C737 B.n697 VSUBS 0.009211f
C738 B.n698 VSUBS 0.009211f
C739 B.n699 VSUBS 0.009211f
C740 B.n700 VSUBS 0.009211f
C741 B.n701 VSUBS 0.009211f
C742 B.n702 VSUBS 0.009211f
C743 B.n703 VSUBS 0.009211f
C744 B.n704 VSUBS 0.009211f
C745 B.n705 VSUBS 0.009211f
C746 B.n706 VSUBS 0.009211f
C747 B.n707 VSUBS 0.009211f
C748 B.n708 VSUBS 0.009211f
C749 B.n709 VSUBS 0.009211f
C750 B.n710 VSUBS 0.009211f
C751 B.n711 VSUBS 0.009211f
C752 B.n712 VSUBS 0.009211f
C753 B.n713 VSUBS 0.009211f
C754 B.n714 VSUBS 0.009211f
C755 B.n715 VSUBS 0.009211f
C756 B.n716 VSUBS 0.009211f
C757 B.n717 VSUBS 0.009211f
C758 B.n718 VSUBS 0.009211f
C759 B.n719 VSUBS 0.009211f
C760 B.n720 VSUBS 0.009211f
C761 B.n721 VSUBS 0.009211f
C762 B.n722 VSUBS 0.009211f
C763 B.n723 VSUBS 0.009211f
C764 B.n724 VSUBS 0.009211f
C765 B.n725 VSUBS 0.009211f
C766 B.n726 VSUBS 0.009211f
C767 B.n727 VSUBS 0.009211f
C768 B.n728 VSUBS 0.009211f
C769 B.n729 VSUBS 0.009211f
C770 B.n730 VSUBS 0.009211f
C771 B.n731 VSUBS 0.009211f
C772 B.n732 VSUBS 0.009211f
C773 B.n733 VSUBS 0.009211f
C774 B.n734 VSUBS 0.009211f
C775 B.n735 VSUBS 0.009211f
C776 B.n736 VSUBS 0.009211f
C777 B.n737 VSUBS 0.009211f
C778 B.n738 VSUBS 0.009211f
C779 B.n739 VSUBS 0.009211f
C780 B.n740 VSUBS 0.009211f
C781 B.n741 VSUBS 0.009211f
C782 B.n742 VSUBS 0.009211f
C783 B.n743 VSUBS 0.009211f
C784 B.n744 VSUBS 0.009211f
C785 B.n745 VSUBS 0.009211f
C786 B.n746 VSUBS 0.009211f
C787 B.n747 VSUBS 0.009211f
C788 B.n748 VSUBS 0.009211f
C789 B.n749 VSUBS 0.009211f
C790 B.n750 VSUBS 0.009211f
C791 B.n751 VSUBS 0.009211f
C792 B.n752 VSUBS 0.009211f
C793 B.n753 VSUBS 0.009211f
C794 B.n754 VSUBS 0.009211f
C795 B.n755 VSUBS 0.009211f
C796 B.n756 VSUBS 0.009211f
C797 B.n757 VSUBS 0.009211f
C798 B.n758 VSUBS 0.009211f
C799 B.n759 VSUBS 0.009211f
C800 B.n760 VSUBS 0.009211f
C801 B.n761 VSUBS 0.009211f
C802 B.n762 VSUBS 0.009211f
C803 B.n763 VSUBS 0.009211f
C804 B.n764 VSUBS 0.009211f
C805 B.n765 VSUBS 0.009211f
C806 B.n766 VSUBS 0.009211f
C807 B.n767 VSUBS 0.01202f
C808 B.n768 VSUBS 0.012804f
C809 B.n769 VSUBS 0.025463f
C810 VDD2.t2 VSUBS 0.158751f
C811 VDD2.t0 VSUBS 0.158751f
C812 VDD2.n0 VSUBS 1.07292f
C813 VDD2.t6 VSUBS 0.158751f
C814 VDD2.t4 VSUBS 0.158751f
C815 VDD2.n1 VSUBS 1.07292f
C816 VDD2.n2 VSUBS 5.17353f
C817 VDD2.t1 VSUBS 0.158751f
C818 VDD2.t7 VSUBS 0.158751f
C819 VDD2.n3 VSUBS 1.05402f
C820 VDD2.n4 VSUBS 4.04721f
C821 VDD2.t5 VSUBS 0.158751f
C822 VDD2.t3 VSUBS 0.158751f
C823 VDD2.n5 VSUBS 1.07288f
C824 VN.t3 VSUBS 1.83163f
C825 VN.n0 VSUBS 0.795219f
C826 VN.n1 VSUBS 0.031958f
C827 VN.n2 VSUBS 0.053778f
C828 VN.n3 VSUBS 0.031958f
C829 VN.n4 VSUBS 0.047211f
C830 VN.n5 VSUBS 0.031958f
C831 VN.n6 VSUBS 0.046653f
C832 VN.n7 VSUBS 0.031958f
C833 VN.n8 VSUBS 0.042506f
C834 VN.t7 VSUBS 1.83163f
C835 VN.n9 VSUBS 0.784131f
C836 VN.t5 VSUBS 2.2414f
C837 VN.n10 VSUBS 0.75586f
C838 VN.n11 VSUBS 0.40018f
C839 VN.n12 VSUBS 0.031958f
C840 VN.n13 VSUBS 0.059562f
C841 VN.n14 VSUBS 0.059562f
C842 VN.n15 VSUBS 0.046653f
C843 VN.n16 VSUBS 0.031958f
C844 VN.n17 VSUBS 0.031958f
C845 VN.n18 VSUBS 0.031958f
C846 VN.n19 VSUBS 0.059562f
C847 VN.n20 VSUBS 0.059562f
C848 VN.t1 VSUBS 1.83163f
C849 VN.n21 VSUBS 0.675675f
C850 VN.n22 VSUBS 0.042506f
C851 VN.n23 VSUBS 0.031958f
C852 VN.n24 VSUBS 0.031958f
C853 VN.n25 VSUBS 0.031958f
C854 VN.n26 VSUBS 0.059562f
C855 VN.n27 VSUBS 0.059562f
C856 VN.n28 VSUBS 0.039529f
C857 VN.n29 VSUBS 0.031958f
C858 VN.n30 VSUBS 0.031958f
C859 VN.n31 VSUBS 0.031958f
C860 VN.n32 VSUBS 0.059562f
C861 VN.n33 VSUBS 0.059562f
C862 VN.n34 VSUBS 0.037802f
C863 VN.n35 VSUBS 0.05158f
C864 VN.n36 VSUBS 0.091166f
C865 VN.t6 VSUBS 1.83163f
C866 VN.n37 VSUBS 0.795219f
C867 VN.n38 VSUBS 0.031958f
C868 VN.n39 VSUBS 0.053778f
C869 VN.n40 VSUBS 0.031958f
C870 VN.n41 VSUBS 0.047211f
C871 VN.n42 VSUBS 0.031958f
C872 VN.t0 VSUBS 1.83163f
C873 VN.n43 VSUBS 0.675675f
C874 VN.n44 VSUBS 0.046653f
C875 VN.n45 VSUBS 0.031958f
C876 VN.n46 VSUBS 0.042506f
C877 VN.t4 VSUBS 2.2414f
C878 VN.t2 VSUBS 1.83163f
C879 VN.n47 VSUBS 0.784131f
C880 VN.n48 VSUBS 0.75586f
C881 VN.n49 VSUBS 0.400181f
C882 VN.n50 VSUBS 0.031958f
C883 VN.n51 VSUBS 0.059562f
C884 VN.n52 VSUBS 0.059562f
C885 VN.n53 VSUBS 0.046653f
C886 VN.n54 VSUBS 0.031958f
C887 VN.n55 VSUBS 0.031958f
C888 VN.n56 VSUBS 0.031958f
C889 VN.n57 VSUBS 0.059562f
C890 VN.n58 VSUBS 0.059562f
C891 VN.n59 VSUBS 0.042506f
C892 VN.n60 VSUBS 0.031958f
C893 VN.n61 VSUBS 0.031958f
C894 VN.n62 VSUBS 0.031958f
C895 VN.n63 VSUBS 0.059562f
C896 VN.n64 VSUBS 0.059562f
C897 VN.n65 VSUBS 0.039529f
C898 VN.n66 VSUBS 0.031958f
C899 VN.n67 VSUBS 0.031958f
C900 VN.n68 VSUBS 0.031958f
C901 VN.n69 VSUBS 0.059562f
C902 VN.n70 VSUBS 0.059562f
C903 VN.n71 VSUBS 0.037802f
C904 VN.n72 VSUBS 0.05158f
C905 VN.n73 VSUBS 1.89979f
C906 VDD1.t3 VSUBS 0.160471f
C907 VDD1.t7 VSUBS 0.160471f
C908 VDD1.n0 VSUBS 1.08608f
C909 VDD1.t5 VSUBS 0.160471f
C910 VDD1.t6 VSUBS 0.160471f
C911 VDD1.n1 VSUBS 1.08455f
C912 VDD1.t0 VSUBS 0.160471f
C913 VDD1.t2 VSUBS 0.160471f
C914 VDD1.n2 VSUBS 1.08455f
C915 VDD1.n3 VSUBS 5.29927f
C916 VDD1.t1 VSUBS 0.160471f
C917 VDD1.t4 VSUBS 0.160471f
C918 VDD1.n4 VSUBS 1.06544f
C919 VDD1.n5 VSUBS 4.13318f
C920 VTAIL.t4 VSUBS 0.146293f
C921 VTAIL.t6 VSUBS 0.146293f
C922 VTAIL.n0 VSUBS 0.863398f
C923 VTAIL.n1 VSUBS 0.905054f
C924 VTAIL.n2 VSUBS 0.033996f
C925 VTAIL.n3 VSUBS 0.030701f
C926 VTAIL.n4 VSUBS 0.016497f
C927 VTAIL.n5 VSUBS 0.038994f
C928 VTAIL.n6 VSUBS 0.017468f
C929 VTAIL.n7 VSUBS 0.030701f
C930 VTAIL.n8 VSUBS 0.016497f
C931 VTAIL.n9 VSUBS 0.038994f
C932 VTAIL.n10 VSUBS 0.017468f
C933 VTAIL.n11 VSUBS 0.136066f
C934 VTAIL.t5 VSUBS 0.083723f
C935 VTAIL.n12 VSUBS 0.029245f
C936 VTAIL.n13 VSUBS 0.024793f
C937 VTAIL.n14 VSUBS 0.016497f
C938 VTAIL.n15 VSUBS 0.708344f
C939 VTAIL.n16 VSUBS 0.030701f
C940 VTAIL.n17 VSUBS 0.016497f
C941 VTAIL.n18 VSUBS 0.017468f
C942 VTAIL.n19 VSUBS 0.038994f
C943 VTAIL.n20 VSUBS 0.038994f
C944 VTAIL.n21 VSUBS 0.017468f
C945 VTAIL.n22 VSUBS 0.016497f
C946 VTAIL.n23 VSUBS 0.030701f
C947 VTAIL.n24 VSUBS 0.030701f
C948 VTAIL.n25 VSUBS 0.016497f
C949 VTAIL.n26 VSUBS 0.017468f
C950 VTAIL.n27 VSUBS 0.038994f
C951 VTAIL.n28 VSUBS 0.095293f
C952 VTAIL.n29 VSUBS 0.017468f
C953 VTAIL.n30 VSUBS 0.016497f
C954 VTAIL.n31 VSUBS 0.072222f
C955 VTAIL.n32 VSUBS 0.048f
C956 VTAIL.n33 VSUBS 0.40771f
C957 VTAIL.n34 VSUBS 0.033996f
C958 VTAIL.n35 VSUBS 0.030701f
C959 VTAIL.n36 VSUBS 0.016497f
C960 VTAIL.n37 VSUBS 0.038994f
C961 VTAIL.n38 VSUBS 0.017468f
C962 VTAIL.n39 VSUBS 0.030701f
C963 VTAIL.n40 VSUBS 0.016497f
C964 VTAIL.n41 VSUBS 0.038994f
C965 VTAIL.n42 VSUBS 0.017468f
C966 VTAIL.n43 VSUBS 0.136066f
C967 VTAIL.t15 VSUBS 0.083723f
C968 VTAIL.n44 VSUBS 0.029245f
C969 VTAIL.n45 VSUBS 0.024793f
C970 VTAIL.n46 VSUBS 0.016497f
C971 VTAIL.n47 VSUBS 0.708344f
C972 VTAIL.n48 VSUBS 0.030701f
C973 VTAIL.n49 VSUBS 0.016497f
C974 VTAIL.n50 VSUBS 0.017468f
C975 VTAIL.n51 VSUBS 0.038994f
C976 VTAIL.n52 VSUBS 0.038994f
C977 VTAIL.n53 VSUBS 0.017468f
C978 VTAIL.n54 VSUBS 0.016497f
C979 VTAIL.n55 VSUBS 0.030701f
C980 VTAIL.n56 VSUBS 0.030701f
C981 VTAIL.n57 VSUBS 0.016497f
C982 VTAIL.n58 VSUBS 0.017468f
C983 VTAIL.n59 VSUBS 0.038994f
C984 VTAIL.n60 VSUBS 0.095293f
C985 VTAIL.n61 VSUBS 0.017468f
C986 VTAIL.n62 VSUBS 0.016497f
C987 VTAIL.n63 VSUBS 0.072222f
C988 VTAIL.n64 VSUBS 0.048f
C989 VTAIL.n65 VSUBS 0.40771f
C990 VTAIL.t10 VSUBS 0.146293f
C991 VTAIL.t9 VSUBS 0.146293f
C992 VTAIL.n66 VSUBS 0.863398f
C993 VTAIL.n67 VSUBS 1.2336f
C994 VTAIL.n68 VSUBS 0.033996f
C995 VTAIL.n69 VSUBS 0.030701f
C996 VTAIL.n70 VSUBS 0.016497f
C997 VTAIL.n71 VSUBS 0.038994f
C998 VTAIL.n72 VSUBS 0.017468f
C999 VTAIL.n73 VSUBS 0.030701f
C1000 VTAIL.n74 VSUBS 0.016497f
C1001 VTAIL.n75 VSUBS 0.038994f
C1002 VTAIL.n76 VSUBS 0.017468f
C1003 VTAIL.n77 VSUBS 0.136066f
C1004 VTAIL.t14 VSUBS 0.083723f
C1005 VTAIL.n78 VSUBS 0.029245f
C1006 VTAIL.n79 VSUBS 0.024793f
C1007 VTAIL.n80 VSUBS 0.016497f
C1008 VTAIL.n81 VSUBS 0.708344f
C1009 VTAIL.n82 VSUBS 0.030701f
C1010 VTAIL.n83 VSUBS 0.016497f
C1011 VTAIL.n84 VSUBS 0.017468f
C1012 VTAIL.n85 VSUBS 0.038994f
C1013 VTAIL.n86 VSUBS 0.038994f
C1014 VTAIL.n87 VSUBS 0.017468f
C1015 VTAIL.n88 VSUBS 0.016497f
C1016 VTAIL.n89 VSUBS 0.030701f
C1017 VTAIL.n90 VSUBS 0.030701f
C1018 VTAIL.n91 VSUBS 0.016497f
C1019 VTAIL.n92 VSUBS 0.017468f
C1020 VTAIL.n93 VSUBS 0.038994f
C1021 VTAIL.n94 VSUBS 0.095293f
C1022 VTAIL.n95 VSUBS 0.017468f
C1023 VTAIL.n96 VSUBS 0.016497f
C1024 VTAIL.n97 VSUBS 0.072222f
C1025 VTAIL.n98 VSUBS 0.048f
C1026 VTAIL.n99 VSUBS 1.62681f
C1027 VTAIL.n100 VSUBS 0.033996f
C1028 VTAIL.n101 VSUBS 0.030701f
C1029 VTAIL.n102 VSUBS 0.016497f
C1030 VTAIL.n103 VSUBS 0.038994f
C1031 VTAIL.n104 VSUBS 0.017468f
C1032 VTAIL.n105 VSUBS 0.030701f
C1033 VTAIL.n106 VSUBS 0.016497f
C1034 VTAIL.n107 VSUBS 0.038994f
C1035 VTAIL.n108 VSUBS 0.017468f
C1036 VTAIL.n109 VSUBS 0.136066f
C1037 VTAIL.t3 VSUBS 0.083723f
C1038 VTAIL.n110 VSUBS 0.029245f
C1039 VTAIL.n111 VSUBS 0.024793f
C1040 VTAIL.n112 VSUBS 0.016497f
C1041 VTAIL.n113 VSUBS 0.708344f
C1042 VTAIL.n114 VSUBS 0.030701f
C1043 VTAIL.n115 VSUBS 0.016497f
C1044 VTAIL.n116 VSUBS 0.017468f
C1045 VTAIL.n117 VSUBS 0.038994f
C1046 VTAIL.n118 VSUBS 0.038994f
C1047 VTAIL.n119 VSUBS 0.017468f
C1048 VTAIL.n120 VSUBS 0.016497f
C1049 VTAIL.n121 VSUBS 0.030701f
C1050 VTAIL.n122 VSUBS 0.030701f
C1051 VTAIL.n123 VSUBS 0.016497f
C1052 VTAIL.n124 VSUBS 0.017468f
C1053 VTAIL.n125 VSUBS 0.038994f
C1054 VTAIL.n126 VSUBS 0.095293f
C1055 VTAIL.n127 VSUBS 0.017468f
C1056 VTAIL.n128 VSUBS 0.016497f
C1057 VTAIL.n129 VSUBS 0.072222f
C1058 VTAIL.n130 VSUBS 0.048f
C1059 VTAIL.n131 VSUBS 1.62681f
C1060 VTAIL.t7 VSUBS 0.146293f
C1061 VTAIL.t2 VSUBS 0.146293f
C1062 VTAIL.n132 VSUBS 0.863404f
C1063 VTAIL.n133 VSUBS 1.23359f
C1064 VTAIL.n134 VSUBS 0.033996f
C1065 VTAIL.n135 VSUBS 0.030701f
C1066 VTAIL.n136 VSUBS 0.016497f
C1067 VTAIL.n137 VSUBS 0.038994f
C1068 VTAIL.n138 VSUBS 0.017468f
C1069 VTAIL.n139 VSUBS 0.030701f
C1070 VTAIL.n140 VSUBS 0.016497f
C1071 VTAIL.n141 VSUBS 0.038994f
C1072 VTAIL.n142 VSUBS 0.017468f
C1073 VTAIL.n143 VSUBS 0.136066f
C1074 VTAIL.t1 VSUBS 0.083723f
C1075 VTAIL.n144 VSUBS 0.029245f
C1076 VTAIL.n145 VSUBS 0.024793f
C1077 VTAIL.n146 VSUBS 0.016497f
C1078 VTAIL.n147 VSUBS 0.708344f
C1079 VTAIL.n148 VSUBS 0.030701f
C1080 VTAIL.n149 VSUBS 0.016497f
C1081 VTAIL.n150 VSUBS 0.017468f
C1082 VTAIL.n151 VSUBS 0.038994f
C1083 VTAIL.n152 VSUBS 0.038994f
C1084 VTAIL.n153 VSUBS 0.017468f
C1085 VTAIL.n154 VSUBS 0.016497f
C1086 VTAIL.n155 VSUBS 0.030701f
C1087 VTAIL.n156 VSUBS 0.030701f
C1088 VTAIL.n157 VSUBS 0.016497f
C1089 VTAIL.n158 VSUBS 0.017468f
C1090 VTAIL.n159 VSUBS 0.038994f
C1091 VTAIL.n160 VSUBS 0.095293f
C1092 VTAIL.n161 VSUBS 0.017468f
C1093 VTAIL.n162 VSUBS 0.016497f
C1094 VTAIL.n163 VSUBS 0.072222f
C1095 VTAIL.n164 VSUBS 0.048f
C1096 VTAIL.n165 VSUBS 0.40771f
C1097 VTAIL.n166 VSUBS 0.033996f
C1098 VTAIL.n167 VSUBS 0.030701f
C1099 VTAIL.n168 VSUBS 0.016497f
C1100 VTAIL.n169 VSUBS 0.038994f
C1101 VTAIL.n170 VSUBS 0.017468f
C1102 VTAIL.n171 VSUBS 0.030701f
C1103 VTAIL.n172 VSUBS 0.016497f
C1104 VTAIL.n173 VSUBS 0.038994f
C1105 VTAIL.n174 VSUBS 0.017468f
C1106 VTAIL.n175 VSUBS 0.136066f
C1107 VTAIL.t11 VSUBS 0.083723f
C1108 VTAIL.n176 VSUBS 0.029245f
C1109 VTAIL.n177 VSUBS 0.024793f
C1110 VTAIL.n178 VSUBS 0.016497f
C1111 VTAIL.n179 VSUBS 0.708344f
C1112 VTAIL.n180 VSUBS 0.030701f
C1113 VTAIL.n181 VSUBS 0.016497f
C1114 VTAIL.n182 VSUBS 0.017468f
C1115 VTAIL.n183 VSUBS 0.038994f
C1116 VTAIL.n184 VSUBS 0.038994f
C1117 VTAIL.n185 VSUBS 0.017468f
C1118 VTAIL.n186 VSUBS 0.016497f
C1119 VTAIL.n187 VSUBS 0.030701f
C1120 VTAIL.n188 VSUBS 0.030701f
C1121 VTAIL.n189 VSUBS 0.016497f
C1122 VTAIL.n190 VSUBS 0.017468f
C1123 VTAIL.n191 VSUBS 0.038994f
C1124 VTAIL.n192 VSUBS 0.095293f
C1125 VTAIL.n193 VSUBS 0.017468f
C1126 VTAIL.n194 VSUBS 0.016497f
C1127 VTAIL.n195 VSUBS 0.072222f
C1128 VTAIL.n196 VSUBS 0.048f
C1129 VTAIL.n197 VSUBS 0.40771f
C1130 VTAIL.t8 VSUBS 0.146293f
C1131 VTAIL.t13 VSUBS 0.146293f
C1132 VTAIL.n198 VSUBS 0.863404f
C1133 VTAIL.n199 VSUBS 1.23359f
C1134 VTAIL.n200 VSUBS 0.033996f
C1135 VTAIL.n201 VSUBS 0.030701f
C1136 VTAIL.n202 VSUBS 0.016497f
C1137 VTAIL.n203 VSUBS 0.038994f
C1138 VTAIL.n204 VSUBS 0.017468f
C1139 VTAIL.n205 VSUBS 0.030701f
C1140 VTAIL.n206 VSUBS 0.016497f
C1141 VTAIL.n207 VSUBS 0.038994f
C1142 VTAIL.n208 VSUBS 0.017468f
C1143 VTAIL.n209 VSUBS 0.136066f
C1144 VTAIL.t12 VSUBS 0.083723f
C1145 VTAIL.n210 VSUBS 0.029245f
C1146 VTAIL.n211 VSUBS 0.024793f
C1147 VTAIL.n212 VSUBS 0.016497f
C1148 VTAIL.n213 VSUBS 0.708344f
C1149 VTAIL.n214 VSUBS 0.030701f
C1150 VTAIL.n215 VSUBS 0.016497f
C1151 VTAIL.n216 VSUBS 0.017468f
C1152 VTAIL.n217 VSUBS 0.038994f
C1153 VTAIL.n218 VSUBS 0.038994f
C1154 VTAIL.n219 VSUBS 0.017468f
C1155 VTAIL.n220 VSUBS 0.016497f
C1156 VTAIL.n221 VSUBS 0.030701f
C1157 VTAIL.n222 VSUBS 0.030701f
C1158 VTAIL.n223 VSUBS 0.016497f
C1159 VTAIL.n224 VSUBS 0.017468f
C1160 VTAIL.n225 VSUBS 0.038994f
C1161 VTAIL.n226 VSUBS 0.095293f
C1162 VTAIL.n227 VSUBS 0.017468f
C1163 VTAIL.n228 VSUBS 0.016497f
C1164 VTAIL.n229 VSUBS 0.072222f
C1165 VTAIL.n230 VSUBS 0.048f
C1166 VTAIL.n231 VSUBS 1.62681f
C1167 VTAIL.n232 VSUBS 0.033996f
C1168 VTAIL.n233 VSUBS 0.030701f
C1169 VTAIL.n234 VSUBS 0.016497f
C1170 VTAIL.n235 VSUBS 0.038994f
C1171 VTAIL.n236 VSUBS 0.017468f
C1172 VTAIL.n237 VSUBS 0.030701f
C1173 VTAIL.n238 VSUBS 0.016497f
C1174 VTAIL.n239 VSUBS 0.038994f
C1175 VTAIL.n240 VSUBS 0.017468f
C1176 VTAIL.n241 VSUBS 0.136066f
C1177 VTAIL.t0 VSUBS 0.083723f
C1178 VTAIL.n242 VSUBS 0.029245f
C1179 VTAIL.n243 VSUBS 0.024793f
C1180 VTAIL.n244 VSUBS 0.016497f
C1181 VTAIL.n245 VSUBS 0.708344f
C1182 VTAIL.n246 VSUBS 0.030701f
C1183 VTAIL.n247 VSUBS 0.016497f
C1184 VTAIL.n248 VSUBS 0.017468f
C1185 VTAIL.n249 VSUBS 0.038994f
C1186 VTAIL.n250 VSUBS 0.038994f
C1187 VTAIL.n251 VSUBS 0.017468f
C1188 VTAIL.n252 VSUBS 0.016497f
C1189 VTAIL.n253 VSUBS 0.030701f
C1190 VTAIL.n254 VSUBS 0.030701f
C1191 VTAIL.n255 VSUBS 0.016497f
C1192 VTAIL.n256 VSUBS 0.017468f
C1193 VTAIL.n257 VSUBS 0.038994f
C1194 VTAIL.n258 VSUBS 0.095293f
C1195 VTAIL.n259 VSUBS 0.017468f
C1196 VTAIL.n260 VSUBS 0.016497f
C1197 VTAIL.n261 VSUBS 0.072222f
C1198 VTAIL.n262 VSUBS 0.048f
C1199 VTAIL.n263 VSUBS 1.62106f
C1200 VP.t5 VSUBS 2.07017f
C1201 VP.n0 VSUBS 0.898784f
C1202 VP.n1 VSUBS 0.03612f
C1203 VP.n2 VSUBS 0.060781f
C1204 VP.n3 VSUBS 0.03612f
C1205 VP.n4 VSUBS 0.05336f
C1206 VP.n5 VSUBS 0.03612f
C1207 VP.n6 VSUBS 0.052729f
C1208 VP.n7 VSUBS 0.03612f
C1209 VP.n8 VSUBS 0.048042f
C1210 VP.n9 VSUBS 0.03612f
C1211 VP.n10 VSUBS 0.044677f
C1212 VP.n11 VSUBS 0.03612f
C1213 VP.n12 VSUBS 0.042725f
C1214 VP.t3 VSUBS 2.07017f
C1215 VP.n13 VSUBS 0.898784f
C1216 VP.n14 VSUBS 0.03612f
C1217 VP.n15 VSUBS 0.060781f
C1218 VP.n16 VSUBS 0.03612f
C1219 VP.n17 VSUBS 0.05336f
C1220 VP.n18 VSUBS 0.03612f
C1221 VP.n19 VSUBS 0.052729f
C1222 VP.n20 VSUBS 0.03612f
C1223 VP.n21 VSUBS 0.048042f
C1224 VP.t4 VSUBS 2.5333f
C1225 VP.t0 VSUBS 2.07017f
C1226 VP.n22 VSUBS 0.886253f
C1227 VP.n23 VSUBS 0.8543f
C1228 VP.n24 VSUBS 0.452299f
C1229 VP.n25 VSUBS 0.03612f
C1230 VP.n26 VSUBS 0.067319f
C1231 VP.n27 VSUBS 0.067319f
C1232 VP.n28 VSUBS 0.052729f
C1233 VP.n29 VSUBS 0.03612f
C1234 VP.n30 VSUBS 0.03612f
C1235 VP.n31 VSUBS 0.03612f
C1236 VP.n32 VSUBS 0.067319f
C1237 VP.n33 VSUBS 0.067319f
C1238 VP.t6 VSUBS 2.07017f
C1239 VP.n34 VSUBS 0.763671f
C1240 VP.n35 VSUBS 0.048042f
C1241 VP.n36 VSUBS 0.03612f
C1242 VP.n37 VSUBS 0.03612f
C1243 VP.n38 VSUBS 0.03612f
C1244 VP.n39 VSUBS 0.067319f
C1245 VP.n40 VSUBS 0.067319f
C1246 VP.n41 VSUBS 0.044677f
C1247 VP.n42 VSUBS 0.03612f
C1248 VP.n43 VSUBS 0.03612f
C1249 VP.n44 VSUBS 0.03612f
C1250 VP.n45 VSUBS 0.067319f
C1251 VP.n46 VSUBS 0.067319f
C1252 VP.n47 VSUBS 0.042725f
C1253 VP.n48 VSUBS 0.058297f
C1254 VP.n49 VSUBS 2.13254f
C1255 VP.t2 VSUBS 2.07017f
C1256 VP.n50 VSUBS 0.898784f
C1257 VP.n51 VSUBS 2.15797f
C1258 VP.n52 VSUBS 0.058297f
C1259 VP.n53 VSUBS 0.03612f
C1260 VP.n54 VSUBS 0.067319f
C1261 VP.n55 VSUBS 0.067319f
C1262 VP.n56 VSUBS 0.060781f
C1263 VP.n57 VSUBS 0.03612f
C1264 VP.n58 VSUBS 0.03612f
C1265 VP.n59 VSUBS 0.03612f
C1266 VP.n60 VSUBS 0.067319f
C1267 VP.n61 VSUBS 0.067319f
C1268 VP.t1 VSUBS 2.07017f
C1269 VP.n62 VSUBS 0.763671f
C1270 VP.n63 VSUBS 0.05336f
C1271 VP.n64 VSUBS 0.03612f
C1272 VP.n65 VSUBS 0.03612f
C1273 VP.n66 VSUBS 0.03612f
C1274 VP.n67 VSUBS 0.067319f
C1275 VP.n68 VSUBS 0.067319f
C1276 VP.n69 VSUBS 0.052729f
C1277 VP.n70 VSUBS 0.03612f
C1278 VP.n71 VSUBS 0.03612f
C1279 VP.n72 VSUBS 0.03612f
C1280 VP.n73 VSUBS 0.067319f
C1281 VP.n74 VSUBS 0.067319f
C1282 VP.t7 VSUBS 2.07017f
C1283 VP.n75 VSUBS 0.763671f
C1284 VP.n76 VSUBS 0.048042f
C1285 VP.n77 VSUBS 0.03612f
C1286 VP.n78 VSUBS 0.03612f
C1287 VP.n79 VSUBS 0.03612f
C1288 VP.n80 VSUBS 0.067319f
C1289 VP.n81 VSUBS 0.067319f
C1290 VP.n82 VSUBS 0.044677f
C1291 VP.n83 VSUBS 0.03612f
C1292 VP.n84 VSUBS 0.03612f
C1293 VP.n85 VSUBS 0.03612f
C1294 VP.n86 VSUBS 0.067319f
C1295 VP.n87 VSUBS 0.067319f
C1296 VP.n88 VSUBS 0.042725f
C1297 VP.n89 VSUBS 0.058297f
C1298 VP.n90 VSUBS 0.103039f
.ends

