* NGSPICE file created from diff_pair_sample_1679.ext - technology: sky130A

.subckt diff_pair_sample_1679 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t7 VP.t0 VDD1.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=7.6167 pd=39.84 as=3.22245 ps=19.86 w=19.53 l=1.91
X1 VTAIL.t2 VN.t0 VDD2.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=7.6167 pd=39.84 as=3.22245 ps=19.86 w=19.53 l=1.91
X2 VDD2.t2 VN.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=3.22245 pd=19.86 as=7.6167 ps=39.84 w=19.53 l=1.91
X3 B.t17 B.t15 B.t16 B.t12 sky130_fd_pr__nfet_01v8 ad=7.6167 pd=39.84 as=0 ps=0 w=19.53 l=1.91
X4 VDD1.t0 VP.t1 VTAIL.t6 B.t0 sky130_fd_pr__nfet_01v8 ad=3.22245 pd=19.86 as=7.6167 ps=39.84 w=19.53 l=1.91
X5 VDD1.t1 VP.t2 VTAIL.t5 B.t1 sky130_fd_pr__nfet_01v8 ad=3.22245 pd=19.86 as=7.6167 ps=39.84 w=19.53 l=1.91
X6 VTAIL.t4 VP.t3 VDD1.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=7.6167 pd=39.84 as=3.22245 ps=19.86 w=19.53 l=1.91
X7 VDD2.t1 VN.t2 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=3.22245 pd=19.86 as=7.6167 ps=39.84 w=19.53 l=1.91
X8 VTAIL.t3 VN.t3 VDD2.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=7.6167 pd=39.84 as=3.22245 ps=19.86 w=19.53 l=1.91
X9 B.t14 B.t11 B.t13 B.t12 sky130_fd_pr__nfet_01v8 ad=7.6167 pd=39.84 as=0 ps=0 w=19.53 l=1.91
X10 B.t10 B.t8 B.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=7.6167 pd=39.84 as=0 ps=0 w=19.53 l=1.91
X11 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=7.6167 pd=39.84 as=0 ps=0 w=19.53 l=1.91
R0 VP.n2 VP.t0 281.479
R1 VP.n2 VP.t1 280.962
R2 VP.n4 VP.t3 246.427
R3 VP.n11 VP.t2 246.427
R4 VP.n10 VP.n0 161.3
R5 VP.n9 VP.n8 161.3
R6 VP.n7 VP.n1 161.3
R7 VP.n6 VP.n5 161.3
R8 VP.n4 VP.n3 92.6509
R9 VP.n12 VP.n11 92.6509
R10 VP.n3 VP.n2 57.4222
R11 VP.n9 VP.n1 56.5193
R12 VP.n5 VP.n1 24.4675
R13 VP.n10 VP.n9 24.4675
R14 VP.n5 VP.n4 18.1061
R15 VP.n11 VP.n10 18.1061
R16 VP.n6 VP.n3 0.278367
R17 VP.n12 VP.n0 0.278367
R18 VP.n7 VP.n6 0.189894
R19 VP.n8 VP.n7 0.189894
R20 VP.n8 VP.n0 0.189894
R21 VP VP.n12 0.153454
R22 VDD1 VDD1.n1 111.144
R23 VDD1 VDD1.n0 64.3326
R24 VDD1.n0 VDD1.t2 1.01432
R25 VDD1.n0 VDD1.t0 1.01432
R26 VDD1.n1 VDD1.t3 1.01432
R27 VDD1.n1 VDD1.t1 1.01432
R28 VTAIL.n842 VTAIL.n742 214.453
R29 VTAIL.n100 VTAIL.n0 214.453
R30 VTAIL.n206 VTAIL.n106 214.453
R31 VTAIL.n312 VTAIL.n212 214.453
R32 VTAIL.n736 VTAIL.n636 214.453
R33 VTAIL.n630 VTAIL.n530 214.453
R34 VTAIL.n524 VTAIL.n424 214.453
R35 VTAIL.n418 VTAIL.n318 214.453
R36 VTAIL.n777 VTAIL.n776 185
R37 VTAIL.n774 VTAIL.n773 185
R38 VTAIL.n783 VTAIL.n782 185
R39 VTAIL.n785 VTAIL.n784 185
R40 VTAIL.n770 VTAIL.n769 185
R41 VTAIL.n791 VTAIL.n790 185
R42 VTAIL.n794 VTAIL.n793 185
R43 VTAIL.n792 VTAIL.n766 185
R44 VTAIL.n799 VTAIL.n765 185
R45 VTAIL.n801 VTAIL.n800 185
R46 VTAIL.n803 VTAIL.n802 185
R47 VTAIL.n762 VTAIL.n761 185
R48 VTAIL.n809 VTAIL.n808 185
R49 VTAIL.n811 VTAIL.n810 185
R50 VTAIL.n758 VTAIL.n757 185
R51 VTAIL.n817 VTAIL.n816 185
R52 VTAIL.n819 VTAIL.n818 185
R53 VTAIL.n754 VTAIL.n753 185
R54 VTAIL.n825 VTAIL.n824 185
R55 VTAIL.n827 VTAIL.n826 185
R56 VTAIL.n750 VTAIL.n749 185
R57 VTAIL.n833 VTAIL.n832 185
R58 VTAIL.n835 VTAIL.n834 185
R59 VTAIL.n746 VTAIL.n745 185
R60 VTAIL.n841 VTAIL.n840 185
R61 VTAIL.n843 VTAIL.n842 185
R62 VTAIL.n35 VTAIL.n34 185
R63 VTAIL.n32 VTAIL.n31 185
R64 VTAIL.n41 VTAIL.n40 185
R65 VTAIL.n43 VTAIL.n42 185
R66 VTAIL.n28 VTAIL.n27 185
R67 VTAIL.n49 VTAIL.n48 185
R68 VTAIL.n52 VTAIL.n51 185
R69 VTAIL.n50 VTAIL.n24 185
R70 VTAIL.n57 VTAIL.n23 185
R71 VTAIL.n59 VTAIL.n58 185
R72 VTAIL.n61 VTAIL.n60 185
R73 VTAIL.n20 VTAIL.n19 185
R74 VTAIL.n67 VTAIL.n66 185
R75 VTAIL.n69 VTAIL.n68 185
R76 VTAIL.n16 VTAIL.n15 185
R77 VTAIL.n75 VTAIL.n74 185
R78 VTAIL.n77 VTAIL.n76 185
R79 VTAIL.n12 VTAIL.n11 185
R80 VTAIL.n83 VTAIL.n82 185
R81 VTAIL.n85 VTAIL.n84 185
R82 VTAIL.n8 VTAIL.n7 185
R83 VTAIL.n91 VTAIL.n90 185
R84 VTAIL.n93 VTAIL.n92 185
R85 VTAIL.n4 VTAIL.n3 185
R86 VTAIL.n99 VTAIL.n98 185
R87 VTAIL.n101 VTAIL.n100 185
R88 VTAIL.n141 VTAIL.n140 185
R89 VTAIL.n138 VTAIL.n137 185
R90 VTAIL.n147 VTAIL.n146 185
R91 VTAIL.n149 VTAIL.n148 185
R92 VTAIL.n134 VTAIL.n133 185
R93 VTAIL.n155 VTAIL.n154 185
R94 VTAIL.n158 VTAIL.n157 185
R95 VTAIL.n156 VTAIL.n130 185
R96 VTAIL.n163 VTAIL.n129 185
R97 VTAIL.n165 VTAIL.n164 185
R98 VTAIL.n167 VTAIL.n166 185
R99 VTAIL.n126 VTAIL.n125 185
R100 VTAIL.n173 VTAIL.n172 185
R101 VTAIL.n175 VTAIL.n174 185
R102 VTAIL.n122 VTAIL.n121 185
R103 VTAIL.n181 VTAIL.n180 185
R104 VTAIL.n183 VTAIL.n182 185
R105 VTAIL.n118 VTAIL.n117 185
R106 VTAIL.n189 VTAIL.n188 185
R107 VTAIL.n191 VTAIL.n190 185
R108 VTAIL.n114 VTAIL.n113 185
R109 VTAIL.n197 VTAIL.n196 185
R110 VTAIL.n199 VTAIL.n198 185
R111 VTAIL.n110 VTAIL.n109 185
R112 VTAIL.n205 VTAIL.n204 185
R113 VTAIL.n207 VTAIL.n206 185
R114 VTAIL.n247 VTAIL.n246 185
R115 VTAIL.n244 VTAIL.n243 185
R116 VTAIL.n253 VTAIL.n252 185
R117 VTAIL.n255 VTAIL.n254 185
R118 VTAIL.n240 VTAIL.n239 185
R119 VTAIL.n261 VTAIL.n260 185
R120 VTAIL.n264 VTAIL.n263 185
R121 VTAIL.n262 VTAIL.n236 185
R122 VTAIL.n269 VTAIL.n235 185
R123 VTAIL.n271 VTAIL.n270 185
R124 VTAIL.n273 VTAIL.n272 185
R125 VTAIL.n232 VTAIL.n231 185
R126 VTAIL.n279 VTAIL.n278 185
R127 VTAIL.n281 VTAIL.n280 185
R128 VTAIL.n228 VTAIL.n227 185
R129 VTAIL.n287 VTAIL.n286 185
R130 VTAIL.n289 VTAIL.n288 185
R131 VTAIL.n224 VTAIL.n223 185
R132 VTAIL.n295 VTAIL.n294 185
R133 VTAIL.n297 VTAIL.n296 185
R134 VTAIL.n220 VTAIL.n219 185
R135 VTAIL.n303 VTAIL.n302 185
R136 VTAIL.n305 VTAIL.n304 185
R137 VTAIL.n216 VTAIL.n215 185
R138 VTAIL.n311 VTAIL.n310 185
R139 VTAIL.n313 VTAIL.n312 185
R140 VTAIL.n737 VTAIL.n736 185
R141 VTAIL.n735 VTAIL.n734 185
R142 VTAIL.n640 VTAIL.n639 185
R143 VTAIL.n729 VTAIL.n728 185
R144 VTAIL.n727 VTAIL.n726 185
R145 VTAIL.n644 VTAIL.n643 185
R146 VTAIL.n721 VTAIL.n720 185
R147 VTAIL.n719 VTAIL.n718 185
R148 VTAIL.n648 VTAIL.n647 185
R149 VTAIL.n713 VTAIL.n712 185
R150 VTAIL.n711 VTAIL.n710 185
R151 VTAIL.n652 VTAIL.n651 185
R152 VTAIL.n705 VTAIL.n704 185
R153 VTAIL.n703 VTAIL.n702 185
R154 VTAIL.n656 VTAIL.n655 185
R155 VTAIL.n697 VTAIL.n696 185
R156 VTAIL.n695 VTAIL.n694 185
R157 VTAIL.n693 VTAIL.n659 185
R158 VTAIL.n663 VTAIL.n660 185
R159 VTAIL.n688 VTAIL.n687 185
R160 VTAIL.n686 VTAIL.n685 185
R161 VTAIL.n665 VTAIL.n664 185
R162 VTAIL.n680 VTAIL.n679 185
R163 VTAIL.n678 VTAIL.n677 185
R164 VTAIL.n669 VTAIL.n668 185
R165 VTAIL.n672 VTAIL.n671 185
R166 VTAIL.n631 VTAIL.n630 185
R167 VTAIL.n629 VTAIL.n628 185
R168 VTAIL.n534 VTAIL.n533 185
R169 VTAIL.n623 VTAIL.n622 185
R170 VTAIL.n621 VTAIL.n620 185
R171 VTAIL.n538 VTAIL.n537 185
R172 VTAIL.n615 VTAIL.n614 185
R173 VTAIL.n613 VTAIL.n612 185
R174 VTAIL.n542 VTAIL.n541 185
R175 VTAIL.n607 VTAIL.n606 185
R176 VTAIL.n605 VTAIL.n604 185
R177 VTAIL.n546 VTAIL.n545 185
R178 VTAIL.n599 VTAIL.n598 185
R179 VTAIL.n597 VTAIL.n596 185
R180 VTAIL.n550 VTAIL.n549 185
R181 VTAIL.n591 VTAIL.n590 185
R182 VTAIL.n589 VTAIL.n588 185
R183 VTAIL.n587 VTAIL.n553 185
R184 VTAIL.n557 VTAIL.n554 185
R185 VTAIL.n582 VTAIL.n581 185
R186 VTAIL.n580 VTAIL.n579 185
R187 VTAIL.n559 VTAIL.n558 185
R188 VTAIL.n574 VTAIL.n573 185
R189 VTAIL.n572 VTAIL.n571 185
R190 VTAIL.n563 VTAIL.n562 185
R191 VTAIL.n566 VTAIL.n565 185
R192 VTAIL.n525 VTAIL.n524 185
R193 VTAIL.n523 VTAIL.n522 185
R194 VTAIL.n428 VTAIL.n427 185
R195 VTAIL.n517 VTAIL.n516 185
R196 VTAIL.n515 VTAIL.n514 185
R197 VTAIL.n432 VTAIL.n431 185
R198 VTAIL.n509 VTAIL.n508 185
R199 VTAIL.n507 VTAIL.n506 185
R200 VTAIL.n436 VTAIL.n435 185
R201 VTAIL.n501 VTAIL.n500 185
R202 VTAIL.n499 VTAIL.n498 185
R203 VTAIL.n440 VTAIL.n439 185
R204 VTAIL.n493 VTAIL.n492 185
R205 VTAIL.n491 VTAIL.n490 185
R206 VTAIL.n444 VTAIL.n443 185
R207 VTAIL.n485 VTAIL.n484 185
R208 VTAIL.n483 VTAIL.n482 185
R209 VTAIL.n481 VTAIL.n447 185
R210 VTAIL.n451 VTAIL.n448 185
R211 VTAIL.n476 VTAIL.n475 185
R212 VTAIL.n474 VTAIL.n473 185
R213 VTAIL.n453 VTAIL.n452 185
R214 VTAIL.n468 VTAIL.n467 185
R215 VTAIL.n466 VTAIL.n465 185
R216 VTAIL.n457 VTAIL.n456 185
R217 VTAIL.n460 VTAIL.n459 185
R218 VTAIL.n419 VTAIL.n418 185
R219 VTAIL.n417 VTAIL.n416 185
R220 VTAIL.n322 VTAIL.n321 185
R221 VTAIL.n411 VTAIL.n410 185
R222 VTAIL.n409 VTAIL.n408 185
R223 VTAIL.n326 VTAIL.n325 185
R224 VTAIL.n403 VTAIL.n402 185
R225 VTAIL.n401 VTAIL.n400 185
R226 VTAIL.n330 VTAIL.n329 185
R227 VTAIL.n395 VTAIL.n394 185
R228 VTAIL.n393 VTAIL.n392 185
R229 VTAIL.n334 VTAIL.n333 185
R230 VTAIL.n387 VTAIL.n386 185
R231 VTAIL.n385 VTAIL.n384 185
R232 VTAIL.n338 VTAIL.n337 185
R233 VTAIL.n379 VTAIL.n378 185
R234 VTAIL.n377 VTAIL.n376 185
R235 VTAIL.n375 VTAIL.n341 185
R236 VTAIL.n345 VTAIL.n342 185
R237 VTAIL.n370 VTAIL.n369 185
R238 VTAIL.n368 VTAIL.n367 185
R239 VTAIL.n347 VTAIL.n346 185
R240 VTAIL.n362 VTAIL.n361 185
R241 VTAIL.n360 VTAIL.n359 185
R242 VTAIL.n351 VTAIL.n350 185
R243 VTAIL.n354 VTAIL.n353 185
R244 VTAIL.t0 VTAIL.n775 149.524
R245 VTAIL.t2 VTAIL.n33 149.524
R246 VTAIL.t5 VTAIL.n139 149.524
R247 VTAIL.t4 VTAIL.n245 149.524
R248 VTAIL.t6 VTAIL.n670 149.524
R249 VTAIL.t7 VTAIL.n564 149.524
R250 VTAIL.t1 VTAIL.n458 149.524
R251 VTAIL.t3 VTAIL.n352 149.524
R252 VTAIL.n776 VTAIL.n773 104.615
R253 VTAIL.n783 VTAIL.n773 104.615
R254 VTAIL.n784 VTAIL.n783 104.615
R255 VTAIL.n784 VTAIL.n769 104.615
R256 VTAIL.n791 VTAIL.n769 104.615
R257 VTAIL.n793 VTAIL.n791 104.615
R258 VTAIL.n793 VTAIL.n792 104.615
R259 VTAIL.n792 VTAIL.n765 104.615
R260 VTAIL.n801 VTAIL.n765 104.615
R261 VTAIL.n802 VTAIL.n801 104.615
R262 VTAIL.n802 VTAIL.n761 104.615
R263 VTAIL.n809 VTAIL.n761 104.615
R264 VTAIL.n810 VTAIL.n809 104.615
R265 VTAIL.n810 VTAIL.n757 104.615
R266 VTAIL.n817 VTAIL.n757 104.615
R267 VTAIL.n818 VTAIL.n817 104.615
R268 VTAIL.n818 VTAIL.n753 104.615
R269 VTAIL.n825 VTAIL.n753 104.615
R270 VTAIL.n826 VTAIL.n825 104.615
R271 VTAIL.n826 VTAIL.n749 104.615
R272 VTAIL.n833 VTAIL.n749 104.615
R273 VTAIL.n834 VTAIL.n833 104.615
R274 VTAIL.n834 VTAIL.n745 104.615
R275 VTAIL.n841 VTAIL.n745 104.615
R276 VTAIL.n842 VTAIL.n841 104.615
R277 VTAIL.n34 VTAIL.n31 104.615
R278 VTAIL.n41 VTAIL.n31 104.615
R279 VTAIL.n42 VTAIL.n41 104.615
R280 VTAIL.n42 VTAIL.n27 104.615
R281 VTAIL.n49 VTAIL.n27 104.615
R282 VTAIL.n51 VTAIL.n49 104.615
R283 VTAIL.n51 VTAIL.n50 104.615
R284 VTAIL.n50 VTAIL.n23 104.615
R285 VTAIL.n59 VTAIL.n23 104.615
R286 VTAIL.n60 VTAIL.n59 104.615
R287 VTAIL.n60 VTAIL.n19 104.615
R288 VTAIL.n67 VTAIL.n19 104.615
R289 VTAIL.n68 VTAIL.n67 104.615
R290 VTAIL.n68 VTAIL.n15 104.615
R291 VTAIL.n75 VTAIL.n15 104.615
R292 VTAIL.n76 VTAIL.n75 104.615
R293 VTAIL.n76 VTAIL.n11 104.615
R294 VTAIL.n83 VTAIL.n11 104.615
R295 VTAIL.n84 VTAIL.n83 104.615
R296 VTAIL.n84 VTAIL.n7 104.615
R297 VTAIL.n91 VTAIL.n7 104.615
R298 VTAIL.n92 VTAIL.n91 104.615
R299 VTAIL.n92 VTAIL.n3 104.615
R300 VTAIL.n99 VTAIL.n3 104.615
R301 VTAIL.n100 VTAIL.n99 104.615
R302 VTAIL.n140 VTAIL.n137 104.615
R303 VTAIL.n147 VTAIL.n137 104.615
R304 VTAIL.n148 VTAIL.n147 104.615
R305 VTAIL.n148 VTAIL.n133 104.615
R306 VTAIL.n155 VTAIL.n133 104.615
R307 VTAIL.n157 VTAIL.n155 104.615
R308 VTAIL.n157 VTAIL.n156 104.615
R309 VTAIL.n156 VTAIL.n129 104.615
R310 VTAIL.n165 VTAIL.n129 104.615
R311 VTAIL.n166 VTAIL.n165 104.615
R312 VTAIL.n166 VTAIL.n125 104.615
R313 VTAIL.n173 VTAIL.n125 104.615
R314 VTAIL.n174 VTAIL.n173 104.615
R315 VTAIL.n174 VTAIL.n121 104.615
R316 VTAIL.n181 VTAIL.n121 104.615
R317 VTAIL.n182 VTAIL.n181 104.615
R318 VTAIL.n182 VTAIL.n117 104.615
R319 VTAIL.n189 VTAIL.n117 104.615
R320 VTAIL.n190 VTAIL.n189 104.615
R321 VTAIL.n190 VTAIL.n113 104.615
R322 VTAIL.n197 VTAIL.n113 104.615
R323 VTAIL.n198 VTAIL.n197 104.615
R324 VTAIL.n198 VTAIL.n109 104.615
R325 VTAIL.n205 VTAIL.n109 104.615
R326 VTAIL.n206 VTAIL.n205 104.615
R327 VTAIL.n246 VTAIL.n243 104.615
R328 VTAIL.n253 VTAIL.n243 104.615
R329 VTAIL.n254 VTAIL.n253 104.615
R330 VTAIL.n254 VTAIL.n239 104.615
R331 VTAIL.n261 VTAIL.n239 104.615
R332 VTAIL.n263 VTAIL.n261 104.615
R333 VTAIL.n263 VTAIL.n262 104.615
R334 VTAIL.n262 VTAIL.n235 104.615
R335 VTAIL.n271 VTAIL.n235 104.615
R336 VTAIL.n272 VTAIL.n271 104.615
R337 VTAIL.n272 VTAIL.n231 104.615
R338 VTAIL.n279 VTAIL.n231 104.615
R339 VTAIL.n280 VTAIL.n279 104.615
R340 VTAIL.n280 VTAIL.n227 104.615
R341 VTAIL.n287 VTAIL.n227 104.615
R342 VTAIL.n288 VTAIL.n287 104.615
R343 VTAIL.n288 VTAIL.n223 104.615
R344 VTAIL.n295 VTAIL.n223 104.615
R345 VTAIL.n296 VTAIL.n295 104.615
R346 VTAIL.n296 VTAIL.n219 104.615
R347 VTAIL.n303 VTAIL.n219 104.615
R348 VTAIL.n304 VTAIL.n303 104.615
R349 VTAIL.n304 VTAIL.n215 104.615
R350 VTAIL.n311 VTAIL.n215 104.615
R351 VTAIL.n312 VTAIL.n311 104.615
R352 VTAIL.n736 VTAIL.n735 104.615
R353 VTAIL.n735 VTAIL.n639 104.615
R354 VTAIL.n728 VTAIL.n639 104.615
R355 VTAIL.n728 VTAIL.n727 104.615
R356 VTAIL.n727 VTAIL.n643 104.615
R357 VTAIL.n720 VTAIL.n643 104.615
R358 VTAIL.n720 VTAIL.n719 104.615
R359 VTAIL.n719 VTAIL.n647 104.615
R360 VTAIL.n712 VTAIL.n647 104.615
R361 VTAIL.n712 VTAIL.n711 104.615
R362 VTAIL.n711 VTAIL.n651 104.615
R363 VTAIL.n704 VTAIL.n651 104.615
R364 VTAIL.n704 VTAIL.n703 104.615
R365 VTAIL.n703 VTAIL.n655 104.615
R366 VTAIL.n696 VTAIL.n655 104.615
R367 VTAIL.n696 VTAIL.n695 104.615
R368 VTAIL.n695 VTAIL.n659 104.615
R369 VTAIL.n663 VTAIL.n659 104.615
R370 VTAIL.n687 VTAIL.n663 104.615
R371 VTAIL.n687 VTAIL.n686 104.615
R372 VTAIL.n686 VTAIL.n664 104.615
R373 VTAIL.n679 VTAIL.n664 104.615
R374 VTAIL.n679 VTAIL.n678 104.615
R375 VTAIL.n678 VTAIL.n668 104.615
R376 VTAIL.n671 VTAIL.n668 104.615
R377 VTAIL.n630 VTAIL.n629 104.615
R378 VTAIL.n629 VTAIL.n533 104.615
R379 VTAIL.n622 VTAIL.n533 104.615
R380 VTAIL.n622 VTAIL.n621 104.615
R381 VTAIL.n621 VTAIL.n537 104.615
R382 VTAIL.n614 VTAIL.n537 104.615
R383 VTAIL.n614 VTAIL.n613 104.615
R384 VTAIL.n613 VTAIL.n541 104.615
R385 VTAIL.n606 VTAIL.n541 104.615
R386 VTAIL.n606 VTAIL.n605 104.615
R387 VTAIL.n605 VTAIL.n545 104.615
R388 VTAIL.n598 VTAIL.n545 104.615
R389 VTAIL.n598 VTAIL.n597 104.615
R390 VTAIL.n597 VTAIL.n549 104.615
R391 VTAIL.n590 VTAIL.n549 104.615
R392 VTAIL.n590 VTAIL.n589 104.615
R393 VTAIL.n589 VTAIL.n553 104.615
R394 VTAIL.n557 VTAIL.n553 104.615
R395 VTAIL.n581 VTAIL.n557 104.615
R396 VTAIL.n581 VTAIL.n580 104.615
R397 VTAIL.n580 VTAIL.n558 104.615
R398 VTAIL.n573 VTAIL.n558 104.615
R399 VTAIL.n573 VTAIL.n572 104.615
R400 VTAIL.n572 VTAIL.n562 104.615
R401 VTAIL.n565 VTAIL.n562 104.615
R402 VTAIL.n524 VTAIL.n523 104.615
R403 VTAIL.n523 VTAIL.n427 104.615
R404 VTAIL.n516 VTAIL.n427 104.615
R405 VTAIL.n516 VTAIL.n515 104.615
R406 VTAIL.n515 VTAIL.n431 104.615
R407 VTAIL.n508 VTAIL.n431 104.615
R408 VTAIL.n508 VTAIL.n507 104.615
R409 VTAIL.n507 VTAIL.n435 104.615
R410 VTAIL.n500 VTAIL.n435 104.615
R411 VTAIL.n500 VTAIL.n499 104.615
R412 VTAIL.n499 VTAIL.n439 104.615
R413 VTAIL.n492 VTAIL.n439 104.615
R414 VTAIL.n492 VTAIL.n491 104.615
R415 VTAIL.n491 VTAIL.n443 104.615
R416 VTAIL.n484 VTAIL.n443 104.615
R417 VTAIL.n484 VTAIL.n483 104.615
R418 VTAIL.n483 VTAIL.n447 104.615
R419 VTAIL.n451 VTAIL.n447 104.615
R420 VTAIL.n475 VTAIL.n451 104.615
R421 VTAIL.n475 VTAIL.n474 104.615
R422 VTAIL.n474 VTAIL.n452 104.615
R423 VTAIL.n467 VTAIL.n452 104.615
R424 VTAIL.n467 VTAIL.n466 104.615
R425 VTAIL.n466 VTAIL.n456 104.615
R426 VTAIL.n459 VTAIL.n456 104.615
R427 VTAIL.n418 VTAIL.n417 104.615
R428 VTAIL.n417 VTAIL.n321 104.615
R429 VTAIL.n410 VTAIL.n321 104.615
R430 VTAIL.n410 VTAIL.n409 104.615
R431 VTAIL.n409 VTAIL.n325 104.615
R432 VTAIL.n402 VTAIL.n325 104.615
R433 VTAIL.n402 VTAIL.n401 104.615
R434 VTAIL.n401 VTAIL.n329 104.615
R435 VTAIL.n394 VTAIL.n329 104.615
R436 VTAIL.n394 VTAIL.n393 104.615
R437 VTAIL.n393 VTAIL.n333 104.615
R438 VTAIL.n386 VTAIL.n333 104.615
R439 VTAIL.n386 VTAIL.n385 104.615
R440 VTAIL.n385 VTAIL.n337 104.615
R441 VTAIL.n378 VTAIL.n337 104.615
R442 VTAIL.n378 VTAIL.n377 104.615
R443 VTAIL.n377 VTAIL.n341 104.615
R444 VTAIL.n345 VTAIL.n341 104.615
R445 VTAIL.n369 VTAIL.n345 104.615
R446 VTAIL.n369 VTAIL.n368 104.615
R447 VTAIL.n368 VTAIL.n346 104.615
R448 VTAIL.n361 VTAIL.n346 104.615
R449 VTAIL.n361 VTAIL.n360 104.615
R450 VTAIL.n360 VTAIL.n350 104.615
R451 VTAIL.n353 VTAIL.n350 104.615
R452 VTAIL.n776 VTAIL.t0 52.3082
R453 VTAIL.n34 VTAIL.t2 52.3082
R454 VTAIL.n140 VTAIL.t5 52.3082
R455 VTAIL.n246 VTAIL.t4 52.3082
R456 VTAIL.n671 VTAIL.t6 52.3082
R457 VTAIL.n565 VTAIL.t7 52.3082
R458 VTAIL.n459 VTAIL.t1 52.3082
R459 VTAIL.n353 VTAIL.t3 52.3082
R460 VTAIL.n847 VTAIL.n846 36.2581
R461 VTAIL.n105 VTAIL.n104 36.2581
R462 VTAIL.n211 VTAIL.n210 36.2581
R463 VTAIL.n317 VTAIL.n316 36.2581
R464 VTAIL.n741 VTAIL.n740 36.2581
R465 VTAIL.n635 VTAIL.n634 36.2581
R466 VTAIL.n529 VTAIL.n528 36.2581
R467 VTAIL.n423 VTAIL.n422 36.2581
R468 VTAIL.n847 VTAIL.n741 31.1341
R469 VTAIL.n423 VTAIL.n317 31.1341
R470 VTAIL.n800 VTAIL.n799 13.1884
R471 VTAIL.n58 VTAIL.n57 13.1884
R472 VTAIL.n164 VTAIL.n163 13.1884
R473 VTAIL.n270 VTAIL.n269 13.1884
R474 VTAIL.n694 VTAIL.n693 13.1884
R475 VTAIL.n588 VTAIL.n587 13.1884
R476 VTAIL.n482 VTAIL.n481 13.1884
R477 VTAIL.n376 VTAIL.n375 13.1884
R478 VTAIL.n798 VTAIL.n766 12.8005
R479 VTAIL.n803 VTAIL.n764 12.8005
R480 VTAIL.n844 VTAIL.n843 12.8005
R481 VTAIL.n56 VTAIL.n24 12.8005
R482 VTAIL.n61 VTAIL.n22 12.8005
R483 VTAIL.n102 VTAIL.n101 12.8005
R484 VTAIL.n162 VTAIL.n130 12.8005
R485 VTAIL.n167 VTAIL.n128 12.8005
R486 VTAIL.n208 VTAIL.n207 12.8005
R487 VTAIL.n268 VTAIL.n236 12.8005
R488 VTAIL.n273 VTAIL.n234 12.8005
R489 VTAIL.n314 VTAIL.n313 12.8005
R490 VTAIL.n738 VTAIL.n737 12.8005
R491 VTAIL.n697 VTAIL.n658 12.8005
R492 VTAIL.n692 VTAIL.n660 12.8005
R493 VTAIL.n632 VTAIL.n631 12.8005
R494 VTAIL.n591 VTAIL.n552 12.8005
R495 VTAIL.n586 VTAIL.n554 12.8005
R496 VTAIL.n526 VTAIL.n525 12.8005
R497 VTAIL.n485 VTAIL.n446 12.8005
R498 VTAIL.n480 VTAIL.n448 12.8005
R499 VTAIL.n420 VTAIL.n419 12.8005
R500 VTAIL.n379 VTAIL.n340 12.8005
R501 VTAIL.n374 VTAIL.n342 12.8005
R502 VTAIL.n795 VTAIL.n794 12.0247
R503 VTAIL.n804 VTAIL.n762 12.0247
R504 VTAIL.n840 VTAIL.n744 12.0247
R505 VTAIL.n53 VTAIL.n52 12.0247
R506 VTAIL.n62 VTAIL.n20 12.0247
R507 VTAIL.n98 VTAIL.n2 12.0247
R508 VTAIL.n159 VTAIL.n158 12.0247
R509 VTAIL.n168 VTAIL.n126 12.0247
R510 VTAIL.n204 VTAIL.n108 12.0247
R511 VTAIL.n265 VTAIL.n264 12.0247
R512 VTAIL.n274 VTAIL.n232 12.0247
R513 VTAIL.n310 VTAIL.n214 12.0247
R514 VTAIL.n734 VTAIL.n638 12.0247
R515 VTAIL.n698 VTAIL.n656 12.0247
R516 VTAIL.n689 VTAIL.n688 12.0247
R517 VTAIL.n628 VTAIL.n532 12.0247
R518 VTAIL.n592 VTAIL.n550 12.0247
R519 VTAIL.n583 VTAIL.n582 12.0247
R520 VTAIL.n522 VTAIL.n426 12.0247
R521 VTAIL.n486 VTAIL.n444 12.0247
R522 VTAIL.n477 VTAIL.n476 12.0247
R523 VTAIL.n416 VTAIL.n320 12.0247
R524 VTAIL.n380 VTAIL.n338 12.0247
R525 VTAIL.n371 VTAIL.n370 12.0247
R526 VTAIL.n790 VTAIL.n768 11.249
R527 VTAIL.n808 VTAIL.n807 11.249
R528 VTAIL.n839 VTAIL.n746 11.249
R529 VTAIL.n48 VTAIL.n26 11.249
R530 VTAIL.n66 VTAIL.n65 11.249
R531 VTAIL.n97 VTAIL.n4 11.249
R532 VTAIL.n154 VTAIL.n132 11.249
R533 VTAIL.n172 VTAIL.n171 11.249
R534 VTAIL.n203 VTAIL.n110 11.249
R535 VTAIL.n260 VTAIL.n238 11.249
R536 VTAIL.n278 VTAIL.n277 11.249
R537 VTAIL.n309 VTAIL.n216 11.249
R538 VTAIL.n733 VTAIL.n640 11.249
R539 VTAIL.n702 VTAIL.n701 11.249
R540 VTAIL.n685 VTAIL.n662 11.249
R541 VTAIL.n627 VTAIL.n534 11.249
R542 VTAIL.n596 VTAIL.n595 11.249
R543 VTAIL.n579 VTAIL.n556 11.249
R544 VTAIL.n521 VTAIL.n428 11.249
R545 VTAIL.n490 VTAIL.n489 11.249
R546 VTAIL.n473 VTAIL.n450 11.249
R547 VTAIL.n415 VTAIL.n322 11.249
R548 VTAIL.n384 VTAIL.n383 11.249
R549 VTAIL.n367 VTAIL.n344 11.249
R550 VTAIL.n789 VTAIL.n770 10.4732
R551 VTAIL.n811 VTAIL.n760 10.4732
R552 VTAIL.n836 VTAIL.n835 10.4732
R553 VTAIL.n47 VTAIL.n28 10.4732
R554 VTAIL.n69 VTAIL.n18 10.4732
R555 VTAIL.n94 VTAIL.n93 10.4732
R556 VTAIL.n153 VTAIL.n134 10.4732
R557 VTAIL.n175 VTAIL.n124 10.4732
R558 VTAIL.n200 VTAIL.n199 10.4732
R559 VTAIL.n259 VTAIL.n240 10.4732
R560 VTAIL.n281 VTAIL.n230 10.4732
R561 VTAIL.n306 VTAIL.n305 10.4732
R562 VTAIL.n730 VTAIL.n729 10.4732
R563 VTAIL.n705 VTAIL.n654 10.4732
R564 VTAIL.n684 VTAIL.n665 10.4732
R565 VTAIL.n624 VTAIL.n623 10.4732
R566 VTAIL.n599 VTAIL.n548 10.4732
R567 VTAIL.n578 VTAIL.n559 10.4732
R568 VTAIL.n518 VTAIL.n517 10.4732
R569 VTAIL.n493 VTAIL.n442 10.4732
R570 VTAIL.n472 VTAIL.n453 10.4732
R571 VTAIL.n412 VTAIL.n411 10.4732
R572 VTAIL.n387 VTAIL.n336 10.4732
R573 VTAIL.n366 VTAIL.n347 10.4732
R574 VTAIL.n777 VTAIL.n775 10.2747
R575 VTAIL.n35 VTAIL.n33 10.2747
R576 VTAIL.n141 VTAIL.n139 10.2747
R577 VTAIL.n247 VTAIL.n245 10.2747
R578 VTAIL.n672 VTAIL.n670 10.2747
R579 VTAIL.n566 VTAIL.n564 10.2747
R580 VTAIL.n460 VTAIL.n458 10.2747
R581 VTAIL.n354 VTAIL.n352 10.2747
R582 VTAIL.n786 VTAIL.n785 9.69747
R583 VTAIL.n812 VTAIL.n758 9.69747
R584 VTAIL.n832 VTAIL.n748 9.69747
R585 VTAIL.n44 VTAIL.n43 9.69747
R586 VTAIL.n70 VTAIL.n16 9.69747
R587 VTAIL.n90 VTAIL.n6 9.69747
R588 VTAIL.n150 VTAIL.n149 9.69747
R589 VTAIL.n176 VTAIL.n122 9.69747
R590 VTAIL.n196 VTAIL.n112 9.69747
R591 VTAIL.n256 VTAIL.n255 9.69747
R592 VTAIL.n282 VTAIL.n228 9.69747
R593 VTAIL.n302 VTAIL.n218 9.69747
R594 VTAIL.n726 VTAIL.n642 9.69747
R595 VTAIL.n706 VTAIL.n652 9.69747
R596 VTAIL.n681 VTAIL.n680 9.69747
R597 VTAIL.n620 VTAIL.n536 9.69747
R598 VTAIL.n600 VTAIL.n546 9.69747
R599 VTAIL.n575 VTAIL.n574 9.69747
R600 VTAIL.n514 VTAIL.n430 9.69747
R601 VTAIL.n494 VTAIL.n440 9.69747
R602 VTAIL.n469 VTAIL.n468 9.69747
R603 VTAIL.n408 VTAIL.n324 9.69747
R604 VTAIL.n388 VTAIL.n334 9.69747
R605 VTAIL.n363 VTAIL.n362 9.69747
R606 VTAIL.n846 VTAIL.n845 9.45567
R607 VTAIL.n104 VTAIL.n103 9.45567
R608 VTAIL.n210 VTAIL.n209 9.45567
R609 VTAIL.n316 VTAIL.n315 9.45567
R610 VTAIL.n740 VTAIL.n739 9.45567
R611 VTAIL.n634 VTAIL.n633 9.45567
R612 VTAIL.n528 VTAIL.n527 9.45567
R613 VTAIL.n422 VTAIL.n421 9.45567
R614 VTAIL.n821 VTAIL.n820 9.3005
R615 VTAIL.n756 VTAIL.n755 9.3005
R616 VTAIL.n815 VTAIL.n814 9.3005
R617 VTAIL.n813 VTAIL.n812 9.3005
R618 VTAIL.n760 VTAIL.n759 9.3005
R619 VTAIL.n807 VTAIL.n806 9.3005
R620 VTAIL.n805 VTAIL.n804 9.3005
R621 VTAIL.n764 VTAIL.n763 9.3005
R622 VTAIL.n779 VTAIL.n778 9.3005
R623 VTAIL.n781 VTAIL.n780 9.3005
R624 VTAIL.n772 VTAIL.n771 9.3005
R625 VTAIL.n787 VTAIL.n786 9.3005
R626 VTAIL.n789 VTAIL.n788 9.3005
R627 VTAIL.n768 VTAIL.n767 9.3005
R628 VTAIL.n796 VTAIL.n795 9.3005
R629 VTAIL.n798 VTAIL.n797 9.3005
R630 VTAIL.n823 VTAIL.n822 9.3005
R631 VTAIL.n752 VTAIL.n751 9.3005
R632 VTAIL.n829 VTAIL.n828 9.3005
R633 VTAIL.n831 VTAIL.n830 9.3005
R634 VTAIL.n748 VTAIL.n747 9.3005
R635 VTAIL.n837 VTAIL.n836 9.3005
R636 VTAIL.n839 VTAIL.n838 9.3005
R637 VTAIL.n744 VTAIL.n743 9.3005
R638 VTAIL.n845 VTAIL.n844 9.3005
R639 VTAIL.n79 VTAIL.n78 9.3005
R640 VTAIL.n14 VTAIL.n13 9.3005
R641 VTAIL.n73 VTAIL.n72 9.3005
R642 VTAIL.n71 VTAIL.n70 9.3005
R643 VTAIL.n18 VTAIL.n17 9.3005
R644 VTAIL.n65 VTAIL.n64 9.3005
R645 VTAIL.n63 VTAIL.n62 9.3005
R646 VTAIL.n22 VTAIL.n21 9.3005
R647 VTAIL.n37 VTAIL.n36 9.3005
R648 VTAIL.n39 VTAIL.n38 9.3005
R649 VTAIL.n30 VTAIL.n29 9.3005
R650 VTAIL.n45 VTAIL.n44 9.3005
R651 VTAIL.n47 VTAIL.n46 9.3005
R652 VTAIL.n26 VTAIL.n25 9.3005
R653 VTAIL.n54 VTAIL.n53 9.3005
R654 VTAIL.n56 VTAIL.n55 9.3005
R655 VTAIL.n81 VTAIL.n80 9.3005
R656 VTAIL.n10 VTAIL.n9 9.3005
R657 VTAIL.n87 VTAIL.n86 9.3005
R658 VTAIL.n89 VTAIL.n88 9.3005
R659 VTAIL.n6 VTAIL.n5 9.3005
R660 VTAIL.n95 VTAIL.n94 9.3005
R661 VTAIL.n97 VTAIL.n96 9.3005
R662 VTAIL.n2 VTAIL.n1 9.3005
R663 VTAIL.n103 VTAIL.n102 9.3005
R664 VTAIL.n185 VTAIL.n184 9.3005
R665 VTAIL.n120 VTAIL.n119 9.3005
R666 VTAIL.n179 VTAIL.n178 9.3005
R667 VTAIL.n177 VTAIL.n176 9.3005
R668 VTAIL.n124 VTAIL.n123 9.3005
R669 VTAIL.n171 VTAIL.n170 9.3005
R670 VTAIL.n169 VTAIL.n168 9.3005
R671 VTAIL.n128 VTAIL.n127 9.3005
R672 VTAIL.n143 VTAIL.n142 9.3005
R673 VTAIL.n145 VTAIL.n144 9.3005
R674 VTAIL.n136 VTAIL.n135 9.3005
R675 VTAIL.n151 VTAIL.n150 9.3005
R676 VTAIL.n153 VTAIL.n152 9.3005
R677 VTAIL.n132 VTAIL.n131 9.3005
R678 VTAIL.n160 VTAIL.n159 9.3005
R679 VTAIL.n162 VTAIL.n161 9.3005
R680 VTAIL.n187 VTAIL.n186 9.3005
R681 VTAIL.n116 VTAIL.n115 9.3005
R682 VTAIL.n193 VTAIL.n192 9.3005
R683 VTAIL.n195 VTAIL.n194 9.3005
R684 VTAIL.n112 VTAIL.n111 9.3005
R685 VTAIL.n201 VTAIL.n200 9.3005
R686 VTAIL.n203 VTAIL.n202 9.3005
R687 VTAIL.n108 VTAIL.n107 9.3005
R688 VTAIL.n209 VTAIL.n208 9.3005
R689 VTAIL.n291 VTAIL.n290 9.3005
R690 VTAIL.n226 VTAIL.n225 9.3005
R691 VTAIL.n285 VTAIL.n284 9.3005
R692 VTAIL.n283 VTAIL.n282 9.3005
R693 VTAIL.n230 VTAIL.n229 9.3005
R694 VTAIL.n277 VTAIL.n276 9.3005
R695 VTAIL.n275 VTAIL.n274 9.3005
R696 VTAIL.n234 VTAIL.n233 9.3005
R697 VTAIL.n249 VTAIL.n248 9.3005
R698 VTAIL.n251 VTAIL.n250 9.3005
R699 VTAIL.n242 VTAIL.n241 9.3005
R700 VTAIL.n257 VTAIL.n256 9.3005
R701 VTAIL.n259 VTAIL.n258 9.3005
R702 VTAIL.n238 VTAIL.n237 9.3005
R703 VTAIL.n266 VTAIL.n265 9.3005
R704 VTAIL.n268 VTAIL.n267 9.3005
R705 VTAIL.n293 VTAIL.n292 9.3005
R706 VTAIL.n222 VTAIL.n221 9.3005
R707 VTAIL.n299 VTAIL.n298 9.3005
R708 VTAIL.n301 VTAIL.n300 9.3005
R709 VTAIL.n218 VTAIL.n217 9.3005
R710 VTAIL.n307 VTAIL.n306 9.3005
R711 VTAIL.n309 VTAIL.n308 9.3005
R712 VTAIL.n214 VTAIL.n213 9.3005
R713 VTAIL.n315 VTAIL.n314 9.3005
R714 VTAIL.n674 VTAIL.n673 9.3005
R715 VTAIL.n676 VTAIL.n675 9.3005
R716 VTAIL.n667 VTAIL.n666 9.3005
R717 VTAIL.n682 VTAIL.n681 9.3005
R718 VTAIL.n684 VTAIL.n683 9.3005
R719 VTAIL.n662 VTAIL.n661 9.3005
R720 VTAIL.n690 VTAIL.n689 9.3005
R721 VTAIL.n692 VTAIL.n691 9.3005
R722 VTAIL.n646 VTAIL.n645 9.3005
R723 VTAIL.n723 VTAIL.n722 9.3005
R724 VTAIL.n725 VTAIL.n724 9.3005
R725 VTAIL.n642 VTAIL.n641 9.3005
R726 VTAIL.n731 VTAIL.n730 9.3005
R727 VTAIL.n733 VTAIL.n732 9.3005
R728 VTAIL.n638 VTAIL.n637 9.3005
R729 VTAIL.n739 VTAIL.n738 9.3005
R730 VTAIL.n717 VTAIL.n716 9.3005
R731 VTAIL.n715 VTAIL.n714 9.3005
R732 VTAIL.n650 VTAIL.n649 9.3005
R733 VTAIL.n709 VTAIL.n708 9.3005
R734 VTAIL.n707 VTAIL.n706 9.3005
R735 VTAIL.n654 VTAIL.n653 9.3005
R736 VTAIL.n701 VTAIL.n700 9.3005
R737 VTAIL.n699 VTAIL.n698 9.3005
R738 VTAIL.n658 VTAIL.n657 9.3005
R739 VTAIL.n568 VTAIL.n567 9.3005
R740 VTAIL.n570 VTAIL.n569 9.3005
R741 VTAIL.n561 VTAIL.n560 9.3005
R742 VTAIL.n576 VTAIL.n575 9.3005
R743 VTAIL.n578 VTAIL.n577 9.3005
R744 VTAIL.n556 VTAIL.n555 9.3005
R745 VTAIL.n584 VTAIL.n583 9.3005
R746 VTAIL.n586 VTAIL.n585 9.3005
R747 VTAIL.n540 VTAIL.n539 9.3005
R748 VTAIL.n617 VTAIL.n616 9.3005
R749 VTAIL.n619 VTAIL.n618 9.3005
R750 VTAIL.n536 VTAIL.n535 9.3005
R751 VTAIL.n625 VTAIL.n624 9.3005
R752 VTAIL.n627 VTAIL.n626 9.3005
R753 VTAIL.n532 VTAIL.n531 9.3005
R754 VTAIL.n633 VTAIL.n632 9.3005
R755 VTAIL.n611 VTAIL.n610 9.3005
R756 VTAIL.n609 VTAIL.n608 9.3005
R757 VTAIL.n544 VTAIL.n543 9.3005
R758 VTAIL.n603 VTAIL.n602 9.3005
R759 VTAIL.n601 VTAIL.n600 9.3005
R760 VTAIL.n548 VTAIL.n547 9.3005
R761 VTAIL.n595 VTAIL.n594 9.3005
R762 VTAIL.n593 VTAIL.n592 9.3005
R763 VTAIL.n552 VTAIL.n551 9.3005
R764 VTAIL.n462 VTAIL.n461 9.3005
R765 VTAIL.n464 VTAIL.n463 9.3005
R766 VTAIL.n455 VTAIL.n454 9.3005
R767 VTAIL.n470 VTAIL.n469 9.3005
R768 VTAIL.n472 VTAIL.n471 9.3005
R769 VTAIL.n450 VTAIL.n449 9.3005
R770 VTAIL.n478 VTAIL.n477 9.3005
R771 VTAIL.n480 VTAIL.n479 9.3005
R772 VTAIL.n434 VTAIL.n433 9.3005
R773 VTAIL.n511 VTAIL.n510 9.3005
R774 VTAIL.n513 VTAIL.n512 9.3005
R775 VTAIL.n430 VTAIL.n429 9.3005
R776 VTAIL.n519 VTAIL.n518 9.3005
R777 VTAIL.n521 VTAIL.n520 9.3005
R778 VTAIL.n426 VTAIL.n425 9.3005
R779 VTAIL.n527 VTAIL.n526 9.3005
R780 VTAIL.n505 VTAIL.n504 9.3005
R781 VTAIL.n503 VTAIL.n502 9.3005
R782 VTAIL.n438 VTAIL.n437 9.3005
R783 VTAIL.n497 VTAIL.n496 9.3005
R784 VTAIL.n495 VTAIL.n494 9.3005
R785 VTAIL.n442 VTAIL.n441 9.3005
R786 VTAIL.n489 VTAIL.n488 9.3005
R787 VTAIL.n487 VTAIL.n486 9.3005
R788 VTAIL.n446 VTAIL.n445 9.3005
R789 VTAIL.n356 VTAIL.n355 9.3005
R790 VTAIL.n358 VTAIL.n357 9.3005
R791 VTAIL.n349 VTAIL.n348 9.3005
R792 VTAIL.n364 VTAIL.n363 9.3005
R793 VTAIL.n366 VTAIL.n365 9.3005
R794 VTAIL.n344 VTAIL.n343 9.3005
R795 VTAIL.n372 VTAIL.n371 9.3005
R796 VTAIL.n374 VTAIL.n373 9.3005
R797 VTAIL.n328 VTAIL.n327 9.3005
R798 VTAIL.n405 VTAIL.n404 9.3005
R799 VTAIL.n407 VTAIL.n406 9.3005
R800 VTAIL.n324 VTAIL.n323 9.3005
R801 VTAIL.n413 VTAIL.n412 9.3005
R802 VTAIL.n415 VTAIL.n414 9.3005
R803 VTAIL.n320 VTAIL.n319 9.3005
R804 VTAIL.n421 VTAIL.n420 9.3005
R805 VTAIL.n399 VTAIL.n398 9.3005
R806 VTAIL.n397 VTAIL.n396 9.3005
R807 VTAIL.n332 VTAIL.n331 9.3005
R808 VTAIL.n391 VTAIL.n390 9.3005
R809 VTAIL.n389 VTAIL.n388 9.3005
R810 VTAIL.n336 VTAIL.n335 9.3005
R811 VTAIL.n383 VTAIL.n382 9.3005
R812 VTAIL.n381 VTAIL.n380 9.3005
R813 VTAIL.n340 VTAIL.n339 9.3005
R814 VTAIL.n782 VTAIL.n772 8.92171
R815 VTAIL.n816 VTAIL.n815 8.92171
R816 VTAIL.n831 VTAIL.n750 8.92171
R817 VTAIL.n40 VTAIL.n30 8.92171
R818 VTAIL.n74 VTAIL.n73 8.92171
R819 VTAIL.n89 VTAIL.n8 8.92171
R820 VTAIL.n146 VTAIL.n136 8.92171
R821 VTAIL.n180 VTAIL.n179 8.92171
R822 VTAIL.n195 VTAIL.n114 8.92171
R823 VTAIL.n252 VTAIL.n242 8.92171
R824 VTAIL.n286 VTAIL.n285 8.92171
R825 VTAIL.n301 VTAIL.n220 8.92171
R826 VTAIL.n725 VTAIL.n644 8.92171
R827 VTAIL.n710 VTAIL.n709 8.92171
R828 VTAIL.n677 VTAIL.n667 8.92171
R829 VTAIL.n619 VTAIL.n538 8.92171
R830 VTAIL.n604 VTAIL.n603 8.92171
R831 VTAIL.n571 VTAIL.n561 8.92171
R832 VTAIL.n513 VTAIL.n432 8.92171
R833 VTAIL.n498 VTAIL.n497 8.92171
R834 VTAIL.n465 VTAIL.n455 8.92171
R835 VTAIL.n407 VTAIL.n326 8.92171
R836 VTAIL.n392 VTAIL.n391 8.92171
R837 VTAIL.n359 VTAIL.n349 8.92171
R838 VTAIL.n846 VTAIL.n742 8.2187
R839 VTAIL.n104 VTAIL.n0 8.2187
R840 VTAIL.n210 VTAIL.n106 8.2187
R841 VTAIL.n316 VTAIL.n212 8.2187
R842 VTAIL.n740 VTAIL.n636 8.2187
R843 VTAIL.n634 VTAIL.n530 8.2187
R844 VTAIL.n528 VTAIL.n424 8.2187
R845 VTAIL.n422 VTAIL.n318 8.2187
R846 VTAIL.n781 VTAIL.n774 8.14595
R847 VTAIL.n819 VTAIL.n756 8.14595
R848 VTAIL.n828 VTAIL.n827 8.14595
R849 VTAIL.n39 VTAIL.n32 8.14595
R850 VTAIL.n77 VTAIL.n14 8.14595
R851 VTAIL.n86 VTAIL.n85 8.14595
R852 VTAIL.n145 VTAIL.n138 8.14595
R853 VTAIL.n183 VTAIL.n120 8.14595
R854 VTAIL.n192 VTAIL.n191 8.14595
R855 VTAIL.n251 VTAIL.n244 8.14595
R856 VTAIL.n289 VTAIL.n226 8.14595
R857 VTAIL.n298 VTAIL.n297 8.14595
R858 VTAIL.n722 VTAIL.n721 8.14595
R859 VTAIL.n713 VTAIL.n650 8.14595
R860 VTAIL.n676 VTAIL.n669 8.14595
R861 VTAIL.n616 VTAIL.n615 8.14595
R862 VTAIL.n607 VTAIL.n544 8.14595
R863 VTAIL.n570 VTAIL.n563 8.14595
R864 VTAIL.n510 VTAIL.n509 8.14595
R865 VTAIL.n501 VTAIL.n438 8.14595
R866 VTAIL.n464 VTAIL.n457 8.14595
R867 VTAIL.n404 VTAIL.n403 8.14595
R868 VTAIL.n395 VTAIL.n332 8.14595
R869 VTAIL.n358 VTAIL.n351 8.14595
R870 VTAIL.n778 VTAIL.n777 7.3702
R871 VTAIL.n820 VTAIL.n754 7.3702
R872 VTAIL.n824 VTAIL.n752 7.3702
R873 VTAIL.n36 VTAIL.n35 7.3702
R874 VTAIL.n78 VTAIL.n12 7.3702
R875 VTAIL.n82 VTAIL.n10 7.3702
R876 VTAIL.n142 VTAIL.n141 7.3702
R877 VTAIL.n184 VTAIL.n118 7.3702
R878 VTAIL.n188 VTAIL.n116 7.3702
R879 VTAIL.n248 VTAIL.n247 7.3702
R880 VTAIL.n290 VTAIL.n224 7.3702
R881 VTAIL.n294 VTAIL.n222 7.3702
R882 VTAIL.n718 VTAIL.n646 7.3702
R883 VTAIL.n714 VTAIL.n648 7.3702
R884 VTAIL.n673 VTAIL.n672 7.3702
R885 VTAIL.n612 VTAIL.n540 7.3702
R886 VTAIL.n608 VTAIL.n542 7.3702
R887 VTAIL.n567 VTAIL.n566 7.3702
R888 VTAIL.n506 VTAIL.n434 7.3702
R889 VTAIL.n502 VTAIL.n436 7.3702
R890 VTAIL.n461 VTAIL.n460 7.3702
R891 VTAIL.n400 VTAIL.n328 7.3702
R892 VTAIL.n396 VTAIL.n330 7.3702
R893 VTAIL.n355 VTAIL.n354 7.3702
R894 VTAIL.n823 VTAIL.n754 6.59444
R895 VTAIL.n824 VTAIL.n823 6.59444
R896 VTAIL.n81 VTAIL.n12 6.59444
R897 VTAIL.n82 VTAIL.n81 6.59444
R898 VTAIL.n187 VTAIL.n118 6.59444
R899 VTAIL.n188 VTAIL.n187 6.59444
R900 VTAIL.n293 VTAIL.n224 6.59444
R901 VTAIL.n294 VTAIL.n293 6.59444
R902 VTAIL.n718 VTAIL.n717 6.59444
R903 VTAIL.n717 VTAIL.n648 6.59444
R904 VTAIL.n612 VTAIL.n611 6.59444
R905 VTAIL.n611 VTAIL.n542 6.59444
R906 VTAIL.n506 VTAIL.n505 6.59444
R907 VTAIL.n505 VTAIL.n436 6.59444
R908 VTAIL.n400 VTAIL.n399 6.59444
R909 VTAIL.n399 VTAIL.n330 6.59444
R910 VTAIL.n778 VTAIL.n774 5.81868
R911 VTAIL.n820 VTAIL.n819 5.81868
R912 VTAIL.n827 VTAIL.n752 5.81868
R913 VTAIL.n36 VTAIL.n32 5.81868
R914 VTAIL.n78 VTAIL.n77 5.81868
R915 VTAIL.n85 VTAIL.n10 5.81868
R916 VTAIL.n142 VTAIL.n138 5.81868
R917 VTAIL.n184 VTAIL.n183 5.81868
R918 VTAIL.n191 VTAIL.n116 5.81868
R919 VTAIL.n248 VTAIL.n244 5.81868
R920 VTAIL.n290 VTAIL.n289 5.81868
R921 VTAIL.n297 VTAIL.n222 5.81868
R922 VTAIL.n721 VTAIL.n646 5.81868
R923 VTAIL.n714 VTAIL.n713 5.81868
R924 VTAIL.n673 VTAIL.n669 5.81868
R925 VTAIL.n615 VTAIL.n540 5.81868
R926 VTAIL.n608 VTAIL.n607 5.81868
R927 VTAIL.n567 VTAIL.n563 5.81868
R928 VTAIL.n509 VTAIL.n434 5.81868
R929 VTAIL.n502 VTAIL.n501 5.81868
R930 VTAIL.n461 VTAIL.n457 5.81868
R931 VTAIL.n403 VTAIL.n328 5.81868
R932 VTAIL.n396 VTAIL.n395 5.81868
R933 VTAIL.n355 VTAIL.n351 5.81868
R934 VTAIL.n844 VTAIL.n742 5.3904
R935 VTAIL.n102 VTAIL.n0 5.3904
R936 VTAIL.n208 VTAIL.n106 5.3904
R937 VTAIL.n314 VTAIL.n212 5.3904
R938 VTAIL.n738 VTAIL.n636 5.3904
R939 VTAIL.n632 VTAIL.n530 5.3904
R940 VTAIL.n526 VTAIL.n424 5.3904
R941 VTAIL.n420 VTAIL.n318 5.3904
R942 VTAIL.n782 VTAIL.n781 5.04292
R943 VTAIL.n816 VTAIL.n756 5.04292
R944 VTAIL.n828 VTAIL.n750 5.04292
R945 VTAIL.n40 VTAIL.n39 5.04292
R946 VTAIL.n74 VTAIL.n14 5.04292
R947 VTAIL.n86 VTAIL.n8 5.04292
R948 VTAIL.n146 VTAIL.n145 5.04292
R949 VTAIL.n180 VTAIL.n120 5.04292
R950 VTAIL.n192 VTAIL.n114 5.04292
R951 VTAIL.n252 VTAIL.n251 5.04292
R952 VTAIL.n286 VTAIL.n226 5.04292
R953 VTAIL.n298 VTAIL.n220 5.04292
R954 VTAIL.n722 VTAIL.n644 5.04292
R955 VTAIL.n710 VTAIL.n650 5.04292
R956 VTAIL.n677 VTAIL.n676 5.04292
R957 VTAIL.n616 VTAIL.n538 5.04292
R958 VTAIL.n604 VTAIL.n544 5.04292
R959 VTAIL.n571 VTAIL.n570 5.04292
R960 VTAIL.n510 VTAIL.n432 5.04292
R961 VTAIL.n498 VTAIL.n438 5.04292
R962 VTAIL.n465 VTAIL.n464 5.04292
R963 VTAIL.n404 VTAIL.n326 5.04292
R964 VTAIL.n392 VTAIL.n332 5.04292
R965 VTAIL.n359 VTAIL.n358 5.04292
R966 VTAIL.n785 VTAIL.n772 4.26717
R967 VTAIL.n815 VTAIL.n758 4.26717
R968 VTAIL.n832 VTAIL.n831 4.26717
R969 VTAIL.n43 VTAIL.n30 4.26717
R970 VTAIL.n73 VTAIL.n16 4.26717
R971 VTAIL.n90 VTAIL.n89 4.26717
R972 VTAIL.n149 VTAIL.n136 4.26717
R973 VTAIL.n179 VTAIL.n122 4.26717
R974 VTAIL.n196 VTAIL.n195 4.26717
R975 VTAIL.n255 VTAIL.n242 4.26717
R976 VTAIL.n285 VTAIL.n228 4.26717
R977 VTAIL.n302 VTAIL.n301 4.26717
R978 VTAIL.n726 VTAIL.n725 4.26717
R979 VTAIL.n709 VTAIL.n652 4.26717
R980 VTAIL.n680 VTAIL.n667 4.26717
R981 VTAIL.n620 VTAIL.n619 4.26717
R982 VTAIL.n603 VTAIL.n546 4.26717
R983 VTAIL.n574 VTAIL.n561 4.26717
R984 VTAIL.n514 VTAIL.n513 4.26717
R985 VTAIL.n497 VTAIL.n440 4.26717
R986 VTAIL.n468 VTAIL.n455 4.26717
R987 VTAIL.n408 VTAIL.n407 4.26717
R988 VTAIL.n391 VTAIL.n334 4.26717
R989 VTAIL.n362 VTAIL.n349 4.26717
R990 VTAIL.n786 VTAIL.n770 3.49141
R991 VTAIL.n812 VTAIL.n811 3.49141
R992 VTAIL.n835 VTAIL.n748 3.49141
R993 VTAIL.n44 VTAIL.n28 3.49141
R994 VTAIL.n70 VTAIL.n69 3.49141
R995 VTAIL.n93 VTAIL.n6 3.49141
R996 VTAIL.n150 VTAIL.n134 3.49141
R997 VTAIL.n176 VTAIL.n175 3.49141
R998 VTAIL.n199 VTAIL.n112 3.49141
R999 VTAIL.n256 VTAIL.n240 3.49141
R1000 VTAIL.n282 VTAIL.n281 3.49141
R1001 VTAIL.n305 VTAIL.n218 3.49141
R1002 VTAIL.n729 VTAIL.n642 3.49141
R1003 VTAIL.n706 VTAIL.n705 3.49141
R1004 VTAIL.n681 VTAIL.n665 3.49141
R1005 VTAIL.n623 VTAIL.n536 3.49141
R1006 VTAIL.n600 VTAIL.n599 3.49141
R1007 VTAIL.n575 VTAIL.n559 3.49141
R1008 VTAIL.n517 VTAIL.n430 3.49141
R1009 VTAIL.n494 VTAIL.n493 3.49141
R1010 VTAIL.n469 VTAIL.n453 3.49141
R1011 VTAIL.n411 VTAIL.n324 3.49141
R1012 VTAIL.n388 VTAIL.n387 3.49141
R1013 VTAIL.n363 VTAIL.n347 3.49141
R1014 VTAIL.n779 VTAIL.n775 2.84303
R1015 VTAIL.n37 VTAIL.n33 2.84303
R1016 VTAIL.n143 VTAIL.n139 2.84303
R1017 VTAIL.n249 VTAIL.n245 2.84303
R1018 VTAIL.n674 VTAIL.n670 2.84303
R1019 VTAIL.n568 VTAIL.n564 2.84303
R1020 VTAIL.n462 VTAIL.n458 2.84303
R1021 VTAIL.n356 VTAIL.n352 2.84303
R1022 VTAIL.n790 VTAIL.n789 2.71565
R1023 VTAIL.n808 VTAIL.n760 2.71565
R1024 VTAIL.n836 VTAIL.n746 2.71565
R1025 VTAIL.n48 VTAIL.n47 2.71565
R1026 VTAIL.n66 VTAIL.n18 2.71565
R1027 VTAIL.n94 VTAIL.n4 2.71565
R1028 VTAIL.n154 VTAIL.n153 2.71565
R1029 VTAIL.n172 VTAIL.n124 2.71565
R1030 VTAIL.n200 VTAIL.n110 2.71565
R1031 VTAIL.n260 VTAIL.n259 2.71565
R1032 VTAIL.n278 VTAIL.n230 2.71565
R1033 VTAIL.n306 VTAIL.n216 2.71565
R1034 VTAIL.n730 VTAIL.n640 2.71565
R1035 VTAIL.n702 VTAIL.n654 2.71565
R1036 VTAIL.n685 VTAIL.n684 2.71565
R1037 VTAIL.n624 VTAIL.n534 2.71565
R1038 VTAIL.n596 VTAIL.n548 2.71565
R1039 VTAIL.n579 VTAIL.n578 2.71565
R1040 VTAIL.n518 VTAIL.n428 2.71565
R1041 VTAIL.n490 VTAIL.n442 2.71565
R1042 VTAIL.n473 VTAIL.n472 2.71565
R1043 VTAIL.n412 VTAIL.n322 2.71565
R1044 VTAIL.n384 VTAIL.n336 2.71565
R1045 VTAIL.n367 VTAIL.n366 2.71565
R1046 VTAIL.n794 VTAIL.n768 1.93989
R1047 VTAIL.n807 VTAIL.n762 1.93989
R1048 VTAIL.n840 VTAIL.n839 1.93989
R1049 VTAIL.n52 VTAIL.n26 1.93989
R1050 VTAIL.n65 VTAIL.n20 1.93989
R1051 VTAIL.n98 VTAIL.n97 1.93989
R1052 VTAIL.n158 VTAIL.n132 1.93989
R1053 VTAIL.n171 VTAIL.n126 1.93989
R1054 VTAIL.n204 VTAIL.n203 1.93989
R1055 VTAIL.n264 VTAIL.n238 1.93989
R1056 VTAIL.n277 VTAIL.n232 1.93989
R1057 VTAIL.n310 VTAIL.n309 1.93989
R1058 VTAIL.n734 VTAIL.n733 1.93989
R1059 VTAIL.n701 VTAIL.n656 1.93989
R1060 VTAIL.n688 VTAIL.n662 1.93989
R1061 VTAIL.n628 VTAIL.n627 1.93989
R1062 VTAIL.n595 VTAIL.n550 1.93989
R1063 VTAIL.n582 VTAIL.n556 1.93989
R1064 VTAIL.n522 VTAIL.n521 1.93989
R1065 VTAIL.n489 VTAIL.n444 1.93989
R1066 VTAIL.n476 VTAIL.n450 1.93989
R1067 VTAIL.n416 VTAIL.n415 1.93989
R1068 VTAIL.n383 VTAIL.n338 1.93989
R1069 VTAIL.n370 VTAIL.n344 1.93989
R1070 VTAIL.n529 VTAIL.n423 1.93153
R1071 VTAIL.n741 VTAIL.n635 1.93153
R1072 VTAIL.n317 VTAIL.n211 1.93153
R1073 VTAIL.n795 VTAIL.n766 1.16414
R1074 VTAIL.n804 VTAIL.n803 1.16414
R1075 VTAIL.n843 VTAIL.n744 1.16414
R1076 VTAIL.n53 VTAIL.n24 1.16414
R1077 VTAIL.n62 VTAIL.n61 1.16414
R1078 VTAIL.n101 VTAIL.n2 1.16414
R1079 VTAIL.n159 VTAIL.n130 1.16414
R1080 VTAIL.n168 VTAIL.n167 1.16414
R1081 VTAIL.n207 VTAIL.n108 1.16414
R1082 VTAIL.n265 VTAIL.n236 1.16414
R1083 VTAIL.n274 VTAIL.n273 1.16414
R1084 VTAIL.n313 VTAIL.n214 1.16414
R1085 VTAIL.n737 VTAIL.n638 1.16414
R1086 VTAIL.n698 VTAIL.n697 1.16414
R1087 VTAIL.n689 VTAIL.n660 1.16414
R1088 VTAIL.n631 VTAIL.n532 1.16414
R1089 VTAIL.n592 VTAIL.n591 1.16414
R1090 VTAIL.n583 VTAIL.n554 1.16414
R1091 VTAIL.n525 VTAIL.n426 1.16414
R1092 VTAIL.n486 VTAIL.n485 1.16414
R1093 VTAIL.n477 VTAIL.n448 1.16414
R1094 VTAIL.n419 VTAIL.n320 1.16414
R1095 VTAIL.n380 VTAIL.n379 1.16414
R1096 VTAIL.n371 VTAIL.n342 1.16414
R1097 VTAIL VTAIL.n105 1.02421
R1098 VTAIL VTAIL.n847 0.907828
R1099 VTAIL.n635 VTAIL.n529 0.470328
R1100 VTAIL.n211 VTAIL.n105 0.470328
R1101 VTAIL.n799 VTAIL.n798 0.388379
R1102 VTAIL.n800 VTAIL.n764 0.388379
R1103 VTAIL.n57 VTAIL.n56 0.388379
R1104 VTAIL.n58 VTAIL.n22 0.388379
R1105 VTAIL.n163 VTAIL.n162 0.388379
R1106 VTAIL.n164 VTAIL.n128 0.388379
R1107 VTAIL.n269 VTAIL.n268 0.388379
R1108 VTAIL.n270 VTAIL.n234 0.388379
R1109 VTAIL.n694 VTAIL.n658 0.388379
R1110 VTAIL.n693 VTAIL.n692 0.388379
R1111 VTAIL.n588 VTAIL.n552 0.388379
R1112 VTAIL.n587 VTAIL.n586 0.388379
R1113 VTAIL.n482 VTAIL.n446 0.388379
R1114 VTAIL.n481 VTAIL.n480 0.388379
R1115 VTAIL.n376 VTAIL.n340 0.388379
R1116 VTAIL.n375 VTAIL.n374 0.388379
R1117 VTAIL.n780 VTAIL.n779 0.155672
R1118 VTAIL.n780 VTAIL.n771 0.155672
R1119 VTAIL.n787 VTAIL.n771 0.155672
R1120 VTAIL.n788 VTAIL.n787 0.155672
R1121 VTAIL.n788 VTAIL.n767 0.155672
R1122 VTAIL.n796 VTAIL.n767 0.155672
R1123 VTAIL.n797 VTAIL.n796 0.155672
R1124 VTAIL.n797 VTAIL.n763 0.155672
R1125 VTAIL.n805 VTAIL.n763 0.155672
R1126 VTAIL.n806 VTAIL.n805 0.155672
R1127 VTAIL.n806 VTAIL.n759 0.155672
R1128 VTAIL.n813 VTAIL.n759 0.155672
R1129 VTAIL.n814 VTAIL.n813 0.155672
R1130 VTAIL.n814 VTAIL.n755 0.155672
R1131 VTAIL.n821 VTAIL.n755 0.155672
R1132 VTAIL.n822 VTAIL.n821 0.155672
R1133 VTAIL.n822 VTAIL.n751 0.155672
R1134 VTAIL.n829 VTAIL.n751 0.155672
R1135 VTAIL.n830 VTAIL.n829 0.155672
R1136 VTAIL.n830 VTAIL.n747 0.155672
R1137 VTAIL.n837 VTAIL.n747 0.155672
R1138 VTAIL.n838 VTAIL.n837 0.155672
R1139 VTAIL.n838 VTAIL.n743 0.155672
R1140 VTAIL.n845 VTAIL.n743 0.155672
R1141 VTAIL.n38 VTAIL.n37 0.155672
R1142 VTAIL.n38 VTAIL.n29 0.155672
R1143 VTAIL.n45 VTAIL.n29 0.155672
R1144 VTAIL.n46 VTAIL.n45 0.155672
R1145 VTAIL.n46 VTAIL.n25 0.155672
R1146 VTAIL.n54 VTAIL.n25 0.155672
R1147 VTAIL.n55 VTAIL.n54 0.155672
R1148 VTAIL.n55 VTAIL.n21 0.155672
R1149 VTAIL.n63 VTAIL.n21 0.155672
R1150 VTAIL.n64 VTAIL.n63 0.155672
R1151 VTAIL.n64 VTAIL.n17 0.155672
R1152 VTAIL.n71 VTAIL.n17 0.155672
R1153 VTAIL.n72 VTAIL.n71 0.155672
R1154 VTAIL.n72 VTAIL.n13 0.155672
R1155 VTAIL.n79 VTAIL.n13 0.155672
R1156 VTAIL.n80 VTAIL.n79 0.155672
R1157 VTAIL.n80 VTAIL.n9 0.155672
R1158 VTAIL.n87 VTAIL.n9 0.155672
R1159 VTAIL.n88 VTAIL.n87 0.155672
R1160 VTAIL.n88 VTAIL.n5 0.155672
R1161 VTAIL.n95 VTAIL.n5 0.155672
R1162 VTAIL.n96 VTAIL.n95 0.155672
R1163 VTAIL.n96 VTAIL.n1 0.155672
R1164 VTAIL.n103 VTAIL.n1 0.155672
R1165 VTAIL.n144 VTAIL.n143 0.155672
R1166 VTAIL.n144 VTAIL.n135 0.155672
R1167 VTAIL.n151 VTAIL.n135 0.155672
R1168 VTAIL.n152 VTAIL.n151 0.155672
R1169 VTAIL.n152 VTAIL.n131 0.155672
R1170 VTAIL.n160 VTAIL.n131 0.155672
R1171 VTAIL.n161 VTAIL.n160 0.155672
R1172 VTAIL.n161 VTAIL.n127 0.155672
R1173 VTAIL.n169 VTAIL.n127 0.155672
R1174 VTAIL.n170 VTAIL.n169 0.155672
R1175 VTAIL.n170 VTAIL.n123 0.155672
R1176 VTAIL.n177 VTAIL.n123 0.155672
R1177 VTAIL.n178 VTAIL.n177 0.155672
R1178 VTAIL.n178 VTAIL.n119 0.155672
R1179 VTAIL.n185 VTAIL.n119 0.155672
R1180 VTAIL.n186 VTAIL.n185 0.155672
R1181 VTAIL.n186 VTAIL.n115 0.155672
R1182 VTAIL.n193 VTAIL.n115 0.155672
R1183 VTAIL.n194 VTAIL.n193 0.155672
R1184 VTAIL.n194 VTAIL.n111 0.155672
R1185 VTAIL.n201 VTAIL.n111 0.155672
R1186 VTAIL.n202 VTAIL.n201 0.155672
R1187 VTAIL.n202 VTAIL.n107 0.155672
R1188 VTAIL.n209 VTAIL.n107 0.155672
R1189 VTAIL.n250 VTAIL.n249 0.155672
R1190 VTAIL.n250 VTAIL.n241 0.155672
R1191 VTAIL.n257 VTAIL.n241 0.155672
R1192 VTAIL.n258 VTAIL.n257 0.155672
R1193 VTAIL.n258 VTAIL.n237 0.155672
R1194 VTAIL.n266 VTAIL.n237 0.155672
R1195 VTAIL.n267 VTAIL.n266 0.155672
R1196 VTAIL.n267 VTAIL.n233 0.155672
R1197 VTAIL.n275 VTAIL.n233 0.155672
R1198 VTAIL.n276 VTAIL.n275 0.155672
R1199 VTAIL.n276 VTAIL.n229 0.155672
R1200 VTAIL.n283 VTAIL.n229 0.155672
R1201 VTAIL.n284 VTAIL.n283 0.155672
R1202 VTAIL.n284 VTAIL.n225 0.155672
R1203 VTAIL.n291 VTAIL.n225 0.155672
R1204 VTAIL.n292 VTAIL.n291 0.155672
R1205 VTAIL.n292 VTAIL.n221 0.155672
R1206 VTAIL.n299 VTAIL.n221 0.155672
R1207 VTAIL.n300 VTAIL.n299 0.155672
R1208 VTAIL.n300 VTAIL.n217 0.155672
R1209 VTAIL.n307 VTAIL.n217 0.155672
R1210 VTAIL.n308 VTAIL.n307 0.155672
R1211 VTAIL.n308 VTAIL.n213 0.155672
R1212 VTAIL.n315 VTAIL.n213 0.155672
R1213 VTAIL.n739 VTAIL.n637 0.155672
R1214 VTAIL.n732 VTAIL.n637 0.155672
R1215 VTAIL.n732 VTAIL.n731 0.155672
R1216 VTAIL.n731 VTAIL.n641 0.155672
R1217 VTAIL.n724 VTAIL.n641 0.155672
R1218 VTAIL.n724 VTAIL.n723 0.155672
R1219 VTAIL.n723 VTAIL.n645 0.155672
R1220 VTAIL.n716 VTAIL.n645 0.155672
R1221 VTAIL.n716 VTAIL.n715 0.155672
R1222 VTAIL.n715 VTAIL.n649 0.155672
R1223 VTAIL.n708 VTAIL.n649 0.155672
R1224 VTAIL.n708 VTAIL.n707 0.155672
R1225 VTAIL.n707 VTAIL.n653 0.155672
R1226 VTAIL.n700 VTAIL.n653 0.155672
R1227 VTAIL.n700 VTAIL.n699 0.155672
R1228 VTAIL.n699 VTAIL.n657 0.155672
R1229 VTAIL.n691 VTAIL.n657 0.155672
R1230 VTAIL.n691 VTAIL.n690 0.155672
R1231 VTAIL.n690 VTAIL.n661 0.155672
R1232 VTAIL.n683 VTAIL.n661 0.155672
R1233 VTAIL.n683 VTAIL.n682 0.155672
R1234 VTAIL.n682 VTAIL.n666 0.155672
R1235 VTAIL.n675 VTAIL.n666 0.155672
R1236 VTAIL.n675 VTAIL.n674 0.155672
R1237 VTAIL.n633 VTAIL.n531 0.155672
R1238 VTAIL.n626 VTAIL.n531 0.155672
R1239 VTAIL.n626 VTAIL.n625 0.155672
R1240 VTAIL.n625 VTAIL.n535 0.155672
R1241 VTAIL.n618 VTAIL.n535 0.155672
R1242 VTAIL.n618 VTAIL.n617 0.155672
R1243 VTAIL.n617 VTAIL.n539 0.155672
R1244 VTAIL.n610 VTAIL.n539 0.155672
R1245 VTAIL.n610 VTAIL.n609 0.155672
R1246 VTAIL.n609 VTAIL.n543 0.155672
R1247 VTAIL.n602 VTAIL.n543 0.155672
R1248 VTAIL.n602 VTAIL.n601 0.155672
R1249 VTAIL.n601 VTAIL.n547 0.155672
R1250 VTAIL.n594 VTAIL.n547 0.155672
R1251 VTAIL.n594 VTAIL.n593 0.155672
R1252 VTAIL.n593 VTAIL.n551 0.155672
R1253 VTAIL.n585 VTAIL.n551 0.155672
R1254 VTAIL.n585 VTAIL.n584 0.155672
R1255 VTAIL.n584 VTAIL.n555 0.155672
R1256 VTAIL.n577 VTAIL.n555 0.155672
R1257 VTAIL.n577 VTAIL.n576 0.155672
R1258 VTAIL.n576 VTAIL.n560 0.155672
R1259 VTAIL.n569 VTAIL.n560 0.155672
R1260 VTAIL.n569 VTAIL.n568 0.155672
R1261 VTAIL.n527 VTAIL.n425 0.155672
R1262 VTAIL.n520 VTAIL.n425 0.155672
R1263 VTAIL.n520 VTAIL.n519 0.155672
R1264 VTAIL.n519 VTAIL.n429 0.155672
R1265 VTAIL.n512 VTAIL.n429 0.155672
R1266 VTAIL.n512 VTAIL.n511 0.155672
R1267 VTAIL.n511 VTAIL.n433 0.155672
R1268 VTAIL.n504 VTAIL.n433 0.155672
R1269 VTAIL.n504 VTAIL.n503 0.155672
R1270 VTAIL.n503 VTAIL.n437 0.155672
R1271 VTAIL.n496 VTAIL.n437 0.155672
R1272 VTAIL.n496 VTAIL.n495 0.155672
R1273 VTAIL.n495 VTAIL.n441 0.155672
R1274 VTAIL.n488 VTAIL.n441 0.155672
R1275 VTAIL.n488 VTAIL.n487 0.155672
R1276 VTAIL.n487 VTAIL.n445 0.155672
R1277 VTAIL.n479 VTAIL.n445 0.155672
R1278 VTAIL.n479 VTAIL.n478 0.155672
R1279 VTAIL.n478 VTAIL.n449 0.155672
R1280 VTAIL.n471 VTAIL.n449 0.155672
R1281 VTAIL.n471 VTAIL.n470 0.155672
R1282 VTAIL.n470 VTAIL.n454 0.155672
R1283 VTAIL.n463 VTAIL.n454 0.155672
R1284 VTAIL.n463 VTAIL.n462 0.155672
R1285 VTAIL.n421 VTAIL.n319 0.155672
R1286 VTAIL.n414 VTAIL.n319 0.155672
R1287 VTAIL.n414 VTAIL.n413 0.155672
R1288 VTAIL.n413 VTAIL.n323 0.155672
R1289 VTAIL.n406 VTAIL.n323 0.155672
R1290 VTAIL.n406 VTAIL.n405 0.155672
R1291 VTAIL.n405 VTAIL.n327 0.155672
R1292 VTAIL.n398 VTAIL.n327 0.155672
R1293 VTAIL.n398 VTAIL.n397 0.155672
R1294 VTAIL.n397 VTAIL.n331 0.155672
R1295 VTAIL.n390 VTAIL.n331 0.155672
R1296 VTAIL.n390 VTAIL.n389 0.155672
R1297 VTAIL.n389 VTAIL.n335 0.155672
R1298 VTAIL.n382 VTAIL.n335 0.155672
R1299 VTAIL.n382 VTAIL.n381 0.155672
R1300 VTAIL.n381 VTAIL.n339 0.155672
R1301 VTAIL.n373 VTAIL.n339 0.155672
R1302 VTAIL.n373 VTAIL.n372 0.155672
R1303 VTAIL.n372 VTAIL.n343 0.155672
R1304 VTAIL.n365 VTAIL.n343 0.155672
R1305 VTAIL.n365 VTAIL.n364 0.155672
R1306 VTAIL.n364 VTAIL.n348 0.155672
R1307 VTAIL.n357 VTAIL.n348 0.155672
R1308 VTAIL.n357 VTAIL.n356 0.155672
R1309 B.n922 B.n921 585
R1310 B.n923 B.n922 585
R1311 B.n398 B.n123 585
R1312 B.n397 B.n396 585
R1313 B.n395 B.n394 585
R1314 B.n393 B.n392 585
R1315 B.n391 B.n390 585
R1316 B.n389 B.n388 585
R1317 B.n387 B.n386 585
R1318 B.n385 B.n384 585
R1319 B.n383 B.n382 585
R1320 B.n381 B.n380 585
R1321 B.n379 B.n378 585
R1322 B.n377 B.n376 585
R1323 B.n375 B.n374 585
R1324 B.n373 B.n372 585
R1325 B.n371 B.n370 585
R1326 B.n369 B.n368 585
R1327 B.n367 B.n366 585
R1328 B.n365 B.n364 585
R1329 B.n363 B.n362 585
R1330 B.n361 B.n360 585
R1331 B.n359 B.n358 585
R1332 B.n357 B.n356 585
R1333 B.n355 B.n354 585
R1334 B.n353 B.n352 585
R1335 B.n351 B.n350 585
R1336 B.n349 B.n348 585
R1337 B.n347 B.n346 585
R1338 B.n345 B.n344 585
R1339 B.n343 B.n342 585
R1340 B.n341 B.n340 585
R1341 B.n339 B.n338 585
R1342 B.n337 B.n336 585
R1343 B.n335 B.n334 585
R1344 B.n333 B.n332 585
R1345 B.n331 B.n330 585
R1346 B.n329 B.n328 585
R1347 B.n327 B.n326 585
R1348 B.n325 B.n324 585
R1349 B.n323 B.n322 585
R1350 B.n321 B.n320 585
R1351 B.n319 B.n318 585
R1352 B.n317 B.n316 585
R1353 B.n315 B.n314 585
R1354 B.n313 B.n312 585
R1355 B.n311 B.n310 585
R1356 B.n309 B.n308 585
R1357 B.n307 B.n306 585
R1358 B.n305 B.n304 585
R1359 B.n303 B.n302 585
R1360 B.n301 B.n300 585
R1361 B.n299 B.n298 585
R1362 B.n297 B.n296 585
R1363 B.n295 B.n294 585
R1364 B.n293 B.n292 585
R1365 B.n291 B.n290 585
R1366 B.n289 B.n288 585
R1367 B.n287 B.n286 585
R1368 B.n285 B.n284 585
R1369 B.n283 B.n282 585
R1370 B.n281 B.n280 585
R1371 B.n279 B.n278 585
R1372 B.n277 B.n276 585
R1373 B.n275 B.n274 585
R1374 B.n272 B.n271 585
R1375 B.n270 B.n269 585
R1376 B.n268 B.n267 585
R1377 B.n266 B.n265 585
R1378 B.n264 B.n263 585
R1379 B.n262 B.n261 585
R1380 B.n260 B.n259 585
R1381 B.n258 B.n257 585
R1382 B.n256 B.n255 585
R1383 B.n254 B.n253 585
R1384 B.n252 B.n251 585
R1385 B.n250 B.n249 585
R1386 B.n248 B.n247 585
R1387 B.n246 B.n245 585
R1388 B.n244 B.n243 585
R1389 B.n242 B.n241 585
R1390 B.n240 B.n239 585
R1391 B.n238 B.n237 585
R1392 B.n236 B.n235 585
R1393 B.n234 B.n233 585
R1394 B.n232 B.n231 585
R1395 B.n230 B.n229 585
R1396 B.n228 B.n227 585
R1397 B.n226 B.n225 585
R1398 B.n224 B.n223 585
R1399 B.n222 B.n221 585
R1400 B.n220 B.n219 585
R1401 B.n218 B.n217 585
R1402 B.n216 B.n215 585
R1403 B.n214 B.n213 585
R1404 B.n212 B.n211 585
R1405 B.n210 B.n209 585
R1406 B.n208 B.n207 585
R1407 B.n206 B.n205 585
R1408 B.n204 B.n203 585
R1409 B.n202 B.n201 585
R1410 B.n200 B.n199 585
R1411 B.n198 B.n197 585
R1412 B.n196 B.n195 585
R1413 B.n194 B.n193 585
R1414 B.n192 B.n191 585
R1415 B.n190 B.n189 585
R1416 B.n188 B.n187 585
R1417 B.n186 B.n185 585
R1418 B.n184 B.n183 585
R1419 B.n182 B.n181 585
R1420 B.n180 B.n179 585
R1421 B.n178 B.n177 585
R1422 B.n176 B.n175 585
R1423 B.n174 B.n173 585
R1424 B.n172 B.n171 585
R1425 B.n170 B.n169 585
R1426 B.n168 B.n167 585
R1427 B.n166 B.n165 585
R1428 B.n164 B.n163 585
R1429 B.n162 B.n161 585
R1430 B.n160 B.n159 585
R1431 B.n158 B.n157 585
R1432 B.n156 B.n155 585
R1433 B.n154 B.n153 585
R1434 B.n152 B.n151 585
R1435 B.n150 B.n149 585
R1436 B.n148 B.n147 585
R1437 B.n146 B.n145 585
R1438 B.n144 B.n143 585
R1439 B.n142 B.n141 585
R1440 B.n140 B.n139 585
R1441 B.n138 B.n137 585
R1442 B.n136 B.n135 585
R1443 B.n134 B.n133 585
R1444 B.n132 B.n131 585
R1445 B.n130 B.n129 585
R1446 B.n53 B.n52 585
R1447 B.n920 B.n54 585
R1448 B.n924 B.n54 585
R1449 B.n919 B.n918 585
R1450 B.n918 B.n50 585
R1451 B.n917 B.n49 585
R1452 B.n930 B.n49 585
R1453 B.n916 B.n48 585
R1454 B.n931 B.n48 585
R1455 B.n915 B.n47 585
R1456 B.n932 B.n47 585
R1457 B.n914 B.n913 585
R1458 B.n913 B.n43 585
R1459 B.n912 B.n42 585
R1460 B.n938 B.n42 585
R1461 B.n911 B.n41 585
R1462 B.n939 B.n41 585
R1463 B.n910 B.n40 585
R1464 B.n940 B.n40 585
R1465 B.n909 B.n908 585
R1466 B.n908 B.n36 585
R1467 B.n907 B.n35 585
R1468 B.n946 B.n35 585
R1469 B.n906 B.n34 585
R1470 B.n947 B.n34 585
R1471 B.n905 B.n33 585
R1472 B.n948 B.n33 585
R1473 B.n904 B.n903 585
R1474 B.n903 B.n29 585
R1475 B.n902 B.n28 585
R1476 B.n954 B.n28 585
R1477 B.n901 B.n27 585
R1478 B.n955 B.n27 585
R1479 B.n900 B.n26 585
R1480 B.n956 B.n26 585
R1481 B.n899 B.n898 585
R1482 B.n898 B.n22 585
R1483 B.n897 B.n21 585
R1484 B.n962 B.n21 585
R1485 B.n896 B.n20 585
R1486 B.n963 B.n20 585
R1487 B.n895 B.n19 585
R1488 B.n964 B.n19 585
R1489 B.n894 B.n893 585
R1490 B.n893 B.n15 585
R1491 B.n892 B.n14 585
R1492 B.n970 B.n14 585
R1493 B.n891 B.n13 585
R1494 B.n971 B.n13 585
R1495 B.n890 B.n12 585
R1496 B.n972 B.n12 585
R1497 B.n889 B.n888 585
R1498 B.n888 B.n8 585
R1499 B.n887 B.n7 585
R1500 B.n978 B.n7 585
R1501 B.n886 B.n6 585
R1502 B.n979 B.n6 585
R1503 B.n885 B.n5 585
R1504 B.n980 B.n5 585
R1505 B.n884 B.n883 585
R1506 B.n883 B.n4 585
R1507 B.n882 B.n399 585
R1508 B.n882 B.n881 585
R1509 B.n872 B.n400 585
R1510 B.n401 B.n400 585
R1511 B.n874 B.n873 585
R1512 B.n875 B.n874 585
R1513 B.n871 B.n405 585
R1514 B.n409 B.n405 585
R1515 B.n870 B.n869 585
R1516 B.n869 B.n868 585
R1517 B.n407 B.n406 585
R1518 B.n408 B.n407 585
R1519 B.n861 B.n860 585
R1520 B.n862 B.n861 585
R1521 B.n859 B.n414 585
R1522 B.n414 B.n413 585
R1523 B.n858 B.n857 585
R1524 B.n857 B.n856 585
R1525 B.n416 B.n415 585
R1526 B.n417 B.n416 585
R1527 B.n849 B.n848 585
R1528 B.n850 B.n849 585
R1529 B.n847 B.n422 585
R1530 B.n422 B.n421 585
R1531 B.n846 B.n845 585
R1532 B.n845 B.n844 585
R1533 B.n424 B.n423 585
R1534 B.n425 B.n424 585
R1535 B.n837 B.n836 585
R1536 B.n838 B.n837 585
R1537 B.n835 B.n430 585
R1538 B.n430 B.n429 585
R1539 B.n834 B.n833 585
R1540 B.n833 B.n832 585
R1541 B.n432 B.n431 585
R1542 B.n433 B.n432 585
R1543 B.n825 B.n824 585
R1544 B.n826 B.n825 585
R1545 B.n823 B.n438 585
R1546 B.n438 B.n437 585
R1547 B.n822 B.n821 585
R1548 B.n821 B.n820 585
R1549 B.n440 B.n439 585
R1550 B.n441 B.n440 585
R1551 B.n813 B.n812 585
R1552 B.n814 B.n813 585
R1553 B.n811 B.n446 585
R1554 B.n446 B.n445 585
R1555 B.n810 B.n809 585
R1556 B.n809 B.n808 585
R1557 B.n448 B.n447 585
R1558 B.n449 B.n448 585
R1559 B.n801 B.n800 585
R1560 B.n802 B.n801 585
R1561 B.n452 B.n451 585
R1562 B.n528 B.n526 585
R1563 B.n529 B.n525 585
R1564 B.n529 B.n453 585
R1565 B.n532 B.n531 585
R1566 B.n533 B.n524 585
R1567 B.n535 B.n534 585
R1568 B.n537 B.n523 585
R1569 B.n540 B.n539 585
R1570 B.n541 B.n522 585
R1571 B.n543 B.n542 585
R1572 B.n545 B.n521 585
R1573 B.n548 B.n547 585
R1574 B.n549 B.n520 585
R1575 B.n551 B.n550 585
R1576 B.n553 B.n519 585
R1577 B.n556 B.n555 585
R1578 B.n557 B.n518 585
R1579 B.n559 B.n558 585
R1580 B.n561 B.n517 585
R1581 B.n564 B.n563 585
R1582 B.n565 B.n516 585
R1583 B.n567 B.n566 585
R1584 B.n569 B.n515 585
R1585 B.n572 B.n571 585
R1586 B.n573 B.n514 585
R1587 B.n575 B.n574 585
R1588 B.n577 B.n513 585
R1589 B.n580 B.n579 585
R1590 B.n581 B.n512 585
R1591 B.n583 B.n582 585
R1592 B.n585 B.n511 585
R1593 B.n588 B.n587 585
R1594 B.n589 B.n510 585
R1595 B.n591 B.n590 585
R1596 B.n593 B.n509 585
R1597 B.n596 B.n595 585
R1598 B.n597 B.n508 585
R1599 B.n599 B.n598 585
R1600 B.n601 B.n507 585
R1601 B.n604 B.n603 585
R1602 B.n605 B.n506 585
R1603 B.n607 B.n606 585
R1604 B.n609 B.n505 585
R1605 B.n612 B.n611 585
R1606 B.n613 B.n504 585
R1607 B.n615 B.n614 585
R1608 B.n617 B.n503 585
R1609 B.n620 B.n619 585
R1610 B.n621 B.n502 585
R1611 B.n623 B.n622 585
R1612 B.n625 B.n501 585
R1613 B.n628 B.n627 585
R1614 B.n629 B.n500 585
R1615 B.n631 B.n630 585
R1616 B.n633 B.n499 585
R1617 B.n636 B.n635 585
R1618 B.n637 B.n498 585
R1619 B.n639 B.n638 585
R1620 B.n641 B.n497 585
R1621 B.n644 B.n643 585
R1622 B.n645 B.n496 585
R1623 B.n647 B.n646 585
R1624 B.n649 B.n495 585
R1625 B.n652 B.n651 585
R1626 B.n654 B.n492 585
R1627 B.n656 B.n655 585
R1628 B.n658 B.n491 585
R1629 B.n661 B.n660 585
R1630 B.n662 B.n490 585
R1631 B.n664 B.n663 585
R1632 B.n666 B.n489 585
R1633 B.n669 B.n668 585
R1634 B.n670 B.n486 585
R1635 B.n673 B.n672 585
R1636 B.n675 B.n485 585
R1637 B.n678 B.n677 585
R1638 B.n679 B.n484 585
R1639 B.n681 B.n680 585
R1640 B.n683 B.n483 585
R1641 B.n686 B.n685 585
R1642 B.n687 B.n482 585
R1643 B.n689 B.n688 585
R1644 B.n691 B.n481 585
R1645 B.n694 B.n693 585
R1646 B.n695 B.n480 585
R1647 B.n697 B.n696 585
R1648 B.n699 B.n479 585
R1649 B.n702 B.n701 585
R1650 B.n703 B.n478 585
R1651 B.n705 B.n704 585
R1652 B.n707 B.n477 585
R1653 B.n710 B.n709 585
R1654 B.n711 B.n476 585
R1655 B.n713 B.n712 585
R1656 B.n715 B.n475 585
R1657 B.n718 B.n717 585
R1658 B.n719 B.n474 585
R1659 B.n721 B.n720 585
R1660 B.n723 B.n473 585
R1661 B.n726 B.n725 585
R1662 B.n727 B.n472 585
R1663 B.n729 B.n728 585
R1664 B.n731 B.n471 585
R1665 B.n734 B.n733 585
R1666 B.n735 B.n470 585
R1667 B.n737 B.n736 585
R1668 B.n739 B.n469 585
R1669 B.n742 B.n741 585
R1670 B.n743 B.n468 585
R1671 B.n745 B.n744 585
R1672 B.n747 B.n467 585
R1673 B.n750 B.n749 585
R1674 B.n751 B.n466 585
R1675 B.n753 B.n752 585
R1676 B.n755 B.n465 585
R1677 B.n758 B.n757 585
R1678 B.n759 B.n464 585
R1679 B.n761 B.n760 585
R1680 B.n763 B.n463 585
R1681 B.n766 B.n765 585
R1682 B.n767 B.n462 585
R1683 B.n769 B.n768 585
R1684 B.n771 B.n461 585
R1685 B.n774 B.n773 585
R1686 B.n775 B.n460 585
R1687 B.n777 B.n776 585
R1688 B.n779 B.n459 585
R1689 B.n782 B.n781 585
R1690 B.n783 B.n458 585
R1691 B.n785 B.n784 585
R1692 B.n787 B.n457 585
R1693 B.n790 B.n789 585
R1694 B.n791 B.n456 585
R1695 B.n793 B.n792 585
R1696 B.n795 B.n455 585
R1697 B.n798 B.n797 585
R1698 B.n799 B.n454 585
R1699 B.n804 B.n803 585
R1700 B.n803 B.n802 585
R1701 B.n805 B.n450 585
R1702 B.n450 B.n449 585
R1703 B.n807 B.n806 585
R1704 B.n808 B.n807 585
R1705 B.n444 B.n443 585
R1706 B.n445 B.n444 585
R1707 B.n816 B.n815 585
R1708 B.n815 B.n814 585
R1709 B.n817 B.n442 585
R1710 B.n442 B.n441 585
R1711 B.n819 B.n818 585
R1712 B.n820 B.n819 585
R1713 B.n436 B.n435 585
R1714 B.n437 B.n436 585
R1715 B.n828 B.n827 585
R1716 B.n827 B.n826 585
R1717 B.n829 B.n434 585
R1718 B.n434 B.n433 585
R1719 B.n831 B.n830 585
R1720 B.n832 B.n831 585
R1721 B.n428 B.n427 585
R1722 B.n429 B.n428 585
R1723 B.n840 B.n839 585
R1724 B.n839 B.n838 585
R1725 B.n841 B.n426 585
R1726 B.n426 B.n425 585
R1727 B.n843 B.n842 585
R1728 B.n844 B.n843 585
R1729 B.n420 B.n419 585
R1730 B.n421 B.n420 585
R1731 B.n852 B.n851 585
R1732 B.n851 B.n850 585
R1733 B.n853 B.n418 585
R1734 B.n418 B.n417 585
R1735 B.n855 B.n854 585
R1736 B.n856 B.n855 585
R1737 B.n412 B.n411 585
R1738 B.n413 B.n412 585
R1739 B.n864 B.n863 585
R1740 B.n863 B.n862 585
R1741 B.n865 B.n410 585
R1742 B.n410 B.n408 585
R1743 B.n867 B.n866 585
R1744 B.n868 B.n867 585
R1745 B.n404 B.n403 585
R1746 B.n409 B.n404 585
R1747 B.n877 B.n876 585
R1748 B.n876 B.n875 585
R1749 B.n878 B.n402 585
R1750 B.n402 B.n401 585
R1751 B.n880 B.n879 585
R1752 B.n881 B.n880 585
R1753 B.n2 B.n0 585
R1754 B.n4 B.n2 585
R1755 B.n3 B.n1 585
R1756 B.n979 B.n3 585
R1757 B.n977 B.n976 585
R1758 B.n978 B.n977 585
R1759 B.n975 B.n9 585
R1760 B.n9 B.n8 585
R1761 B.n974 B.n973 585
R1762 B.n973 B.n972 585
R1763 B.n11 B.n10 585
R1764 B.n971 B.n11 585
R1765 B.n969 B.n968 585
R1766 B.n970 B.n969 585
R1767 B.n967 B.n16 585
R1768 B.n16 B.n15 585
R1769 B.n966 B.n965 585
R1770 B.n965 B.n964 585
R1771 B.n18 B.n17 585
R1772 B.n963 B.n18 585
R1773 B.n961 B.n960 585
R1774 B.n962 B.n961 585
R1775 B.n959 B.n23 585
R1776 B.n23 B.n22 585
R1777 B.n958 B.n957 585
R1778 B.n957 B.n956 585
R1779 B.n25 B.n24 585
R1780 B.n955 B.n25 585
R1781 B.n953 B.n952 585
R1782 B.n954 B.n953 585
R1783 B.n951 B.n30 585
R1784 B.n30 B.n29 585
R1785 B.n950 B.n949 585
R1786 B.n949 B.n948 585
R1787 B.n32 B.n31 585
R1788 B.n947 B.n32 585
R1789 B.n945 B.n944 585
R1790 B.n946 B.n945 585
R1791 B.n943 B.n37 585
R1792 B.n37 B.n36 585
R1793 B.n942 B.n941 585
R1794 B.n941 B.n940 585
R1795 B.n39 B.n38 585
R1796 B.n939 B.n39 585
R1797 B.n937 B.n936 585
R1798 B.n938 B.n937 585
R1799 B.n935 B.n44 585
R1800 B.n44 B.n43 585
R1801 B.n934 B.n933 585
R1802 B.n933 B.n932 585
R1803 B.n46 B.n45 585
R1804 B.n931 B.n46 585
R1805 B.n929 B.n928 585
R1806 B.n930 B.n929 585
R1807 B.n927 B.n51 585
R1808 B.n51 B.n50 585
R1809 B.n926 B.n925 585
R1810 B.n925 B.n924 585
R1811 B.n982 B.n981 585
R1812 B.n981 B.n980 585
R1813 B.n803 B.n452 487.695
R1814 B.n925 B.n53 487.695
R1815 B.n801 B.n454 487.695
R1816 B.n922 B.n54 487.695
R1817 B.n487 B.t10 455.257
R1818 B.n493 B.t7 455.257
R1819 B.n126 B.t16 455.257
R1820 B.n124 B.t13 455.257
R1821 B.n487 B.t8 453.125
R1822 B.n493 B.t4 453.125
R1823 B.n126 B.t15 453.125
R1824 B.n124 B.t11 453.125
R1825 B.n488 B.t9 411.815
R1826 B.n125 B.t14 411.815
R1827 B.n494 B.t6 411.815
R1828 B.n127 B.t17 411.815
R1829 B.n923 B.n122 256.663
R1830 B.n923 B.n121 256.663
R1831 B.n923 B.n120 256.663
R1832 B.n923 B.n119 256.663
R1833 B.n923 B.n118 256.663
R1834 B.n923 B.n117 256.663
R1835 B.n923 B.n116 256.663
R1836 B.n923 B.n115 256.663
R1837 B.n923 B.n114 256.663
R1838 B.n923 B.n113 256.663
R1839 B.n923 B.n112 256.663
R1840 B.n923 B.n111 256.663
R1841 B.n923 B.n110 256.663
R1842 B.n923 B.n109 256.663
R1843 B.n923 B.n108 256.663
R1844 B.n923 B.n107 256.663
R1845 B.n923 B.n106 256.663
R1846 B.n923 B.n105 256.663
R1847 B.n923 B.n104 256.663
R1848 B.n923 B.n103 256.663
R1849 B.n923 B.n102 256.663
R1850 B.n923 B.n101 256.663
R1851 B.n923 B.n100 256.663
R1852 B.n923 B.n99 256.663
R1853 B.n923 B.n98 256.663
R1854 B.n923 B.n97 256.663
R1855 B.n923 B.n96 256.663
R1856 B.n923 B.n95 256.663
R1857 B.n923 B.n94 256.663
R1858 B.n923 B.n93 256.663
R1859 B.n923 B.n92 256.663
R1860 B.n923 B.n91 256.663
R1861 B.n923 B.n90 256.663
R1862 B.n923 B.n89 256.663
R1863 B.n923 B.n88 256.663
R1864 B.n923 B.n87 256.663
R1865 B.n923 B.n86 256.663
R1866 B.n923 B.n85 256.663
R1867 B.n923 B.n84 256.663
R1868 B.n923 B.n83 256.663
R1869 B.n923 B.n82 256.663
R1870 B.n923 B.n81 256.663
R1871 B.n923 B.n80 256.663
R1872 B.n923 B.n79 256.663
R1873 B.n923 B.n78 256.663
R1874 B.n923 B.n77 256.663
R1875 B.n923 B.n76 256.663
R1876 B.n923 B.n75 256.663
R1877 B.n923 B.n74 256.663
R1878 B.n923 B.n73 256.663
R1879 B.n923 B.n72 256.663
R1880 B.n923 B.n71 256.663
R1881 B.n923 B.n70 256.663
R1882 B.n923 B.n69 256.663
R1883 B.n923 B.n68 256.663
R1884 B.n923 B.n67 256.663
R1885 B.n923 B.n66 256.663
R1886 B.n923 B.n65 256.663
R1887 B.n923 B.n64 256.663
R1888 B.n923 B.n63 256.663
R1889 B.n923 B.n62 256.663
R1890 B.n923 B.n61 256.663
R1891 B.n923 B.n60 256.663
R1892 B.n923 B.n59 256.663
R1893 B.n923 B.n58 256.663
R1894 B.n923 B.n57 256.663
R1895 B.n923 B.n56 256.663
R1896 B.n923 B.n55 256.663
R1897 B.n527 B.n453 256.663
R1898 B.n530 B.n453 256.663
R1899 B.n536 B.n453 256.663
R1900 B.n538 B.n453 256.663
R1901 B.n544 B.n453 256.663
R1902 B.n546 B.n453 256.663
R1903 B.n552 B.n453 256.663
R1904 B.n554 B.n453 256.663
R1905 B.n560 B.n453 256.663
R1906 B.n562 B.n453 256.663
R1907 B.n568 B.n453 256.663
R1908 B.n570 B.n453 256.663
R1909 B.n576 B.n453 256.663
R1910 B.n578 B.n453 256.663
R1911 B.n584 B.n453 256.663
R1912 B.n586 B.n453 256.663
R1913 B.n592 B.n453 256.663
R1914 B.n594 B.n453 256.663
R1915 B.n600 B.n453 256.663
R1916 B.n602 B.n453 256.663
R1917 B.n608 B.n453 256.663
R1918 B.n610 B.n453 256.663
R1919 B.n616 B.n453 256.663
R1920 B.n618 B.n453 256.663
R1921 B.n624 B.n453 256.663
R1922 B.n626 B.n453 256.663
R1923 B.n632 B.n453 256.663
R1924 B.n634 B.n453 256.663
R1925 B.n640 B.n453 256.663
R1926 B.n642 B.n453 256.663
R1927 B.n648 B.n453 256.663
R1928 B.n650 B.n453 256.663
R1929 B.n657 B.n453 256.663
R1930 B.n659 B.n453 256.663
R1931 B.n665 B.n453 256.663
R1932 B.n667 B.n453 256.663
R1933 B.n674 B.n453 256.663
R1934 B.n676 B.n453 256.663
R1935 B.n682 B.n453 256.663
R1936 B.n684 B.n453 256.663
R1937 B.n690 B.n453 256.663
R1938 B.n692 B.n453 256.663
R1939 B.n698 B.n453 256.663
R1940 B.n700 B.n453 256.663
R1941 B.n706 B.n453 256.663
R1942 B.n708 B.n453 256.663
R1943 B.n714 B.n453 256.663
R1944 B.n716 B.n453 256.663
R1945 B.n722 B.n453 256.663
R1946 B.n724 B.n453 256.663
R1947 B.n730 B.n453 256.663
R1948 B.n732 B.n453 256.663
R1949 B.n738 B.n453 256.663
R1950 B.n740 B.n453 256.663
R1951 B.n746 B.n453 256.663
R1952 B.n748 B.n453 256.663
R1953 B.n754 B.n453 256.663
R1954 B.n756 B.n453 256.663
R1955 B.n762 B.n453 256.663
R1956 B.n764 B.n453 256.663
R1957 B.n770 B.n453 256.663
R1958 B.n772 B.n453 256.663
R1959 B.n778 B.n453 256.663
R1960 B.n780 B.n453 256.663
R1961 B.n786 B.n453 256.663
R1962 B.n788 B.n453 256.663
R1963 B.n794 B.n453 256.663
R1964 B.n796 B.n453 256.663
R1965 B.n803 B.n450 163.367
R1966 B.n807 B.n450 163.367
R1967 B.n807 B.n444 163.367
R1968 B.n815 B.n444 163.367
R1969 B.n815 B.n442 163.367
R1970 B.n819 B.n442 163.367
R1971 B.n819 B.n436 163.367
R1972 B.n827 B.n436 163.367
R1973 B.n827 B.n434 163.367
R1974 B.n831 B.n434 163.367
R1975 B.n831 B.n428 163.367
R1976 B.n839 B.n428 163.367
R1977 B.n839 B.n426 163.367
R1978 B.n843 B.n426 163.367
R1979 B.n843 B.n420 163.367
R1980 B.n851 B.n420 163.367
R1981 B.n851 B.n418 163.367
R1982 B.n855 B.n418 163.367
R1983 B.n855 B.n412 163.367
R1984 B.n863 B.n412 163.367
R1985 B.n863 B.n410 163.367
R1986 B.n867 B.n410 163.367
R1987 B.n867 B.n404 163.367
R1988 B.n876 B.n404 163.367
R1989 B.n876 B.n402 163.367
R1990 B.n880 B.n402 163.367
R1991 B.n880 B.n2 163.367
R1992 B.n981 B.n2 163.367
R1993 B.n981 B.n3 163.367
R1994 B.n977 B.n3 163.367
R1995 B.n977 B.n9 163.367
R1996 B.n973 B.n9 163.367
R1997 B.n973 B.n11 163.367
R1998 B.n969 B.n11 163.367
R1999 B.n969 B.n16 163.367
R2000 B.n965 B.n16 163.367
R2001 B.n965 B.n18 163.367
R2002 B.n961 B.n18 163.367
R2003 B.n961 B.n23 163.367
R2004 B.n957 B.n23 163.367
R2005 B.n957 B.n25 163.367
R2006 B.n953 B.n25 163.367
R2007 B.n953 B.n30 163.367
R2008 B.n949 B.n30 163.367
R2009 B.n949 B.n32 163.367
R2010 B.n945 B.n32 163.367
R2011 B.n945 B.n37 163.367
R2012 B.n941 B.n37 163.367
R2013 B.n941 B.n39 163.367
R2014 B.n937 B.n39 163.367
R2015 B.n937 B.n44 163.367
R2016 B.n933 B.n44 163.367
R2017 B.n933 B.n46 163.367
R2018 B.n929 B.n46 163.367
R2019 B.n929 B.n51 163.367
R2020 B.n925 B.n51 163.367
R2021 B.n529 B.n528 163.367
R2022 B.n531 B.n529 163.367
R2023 B.n535 B.n524 163.367
R2024 B.n539 B.n537 163.367
R2025 B.n543 B.n522 163.367
R2026 B.n547 B.n545 163.367
R2027 B.n551 B.n520 163.367
R2028 B.n555 B.n553 163.367
R2029 B.n559 B.n518 163.367
R2030 B.n563 B.n561 163.367
R2031 B.n567 B.n516 163.367
R2032 B.n571 B.n569 163.367
R2033 B.n575 B.n514 163.367
R2034 B.n579 B.n577 163.367
R2035 B.n583 B.n512 163.367
R2036 B.n587 B.n585 163.367
R2037 B.n591 B.n510 163.367
R2038 B.n595 B.n593 163.367
R2039 B.n599 B.n508 163.367
R2040 B.n603 B.n601 163.367
R2041 B.n607 B.n506 163.367
R2042 B.n611 B.n609 163.367
R2043 B.n615 B.n504 163.367
R2044 B.n619 B.n617 163.367
R2045 B.n623 B.n502 163.367
R2046 B.n627 B.n625 163.367
R2047 B.n631 B.n500 163.367
R2048 B.n635 B.n633 163.367
R2049 B.n639 B.n498 163.367
R2050 B.n643 B.n641 163.367
R2051 B.n647 B.n496 163.367
R2052 B.n651 B.n649 163.367
R2053 B.n656 B.n492 163.367
R2054 B.n660 B.n658 163.367
R2055 B.n664 B.n490 163.367
R2056 B.n668 B.n666 163.367
R2057 B.n673 B.n486 163.367
R2058 B.n677 B.n675 163.367
R2059 B.n681 B.n484 163.367
R2060 B.n685 B.n683 163.367
R2061 B.n689 B.n482 163.367
R2062 B.n693 B.n691 163.367
R2063 B.n697 B.n480 163.367
R2064 B.n701 B.n699 163.367
R2065 B.n705 B.n478 163.367
R2066 B.n709 B.n707 163.367
R2067 B.n713 B.n476 163.367
R2068 B.n717 B.n715 163.367
R2069 B.n721 B.n474 163.367
R2070 B.n725 B.n723 163.367
R2071 B.n729 B.n472 163.367
R2072 B.n733 B.n731 163.367
R2073 B.n737 B.n470 163.367
R2074 B.n741 B.n739 163.367
R2075 B.n745 B.n468 163.367
R2076 B.n749 B.n747 163.367
R2077 B.n753 B.n466 163.367
R2078 B.n757 B.n755 163.367
R2079 B.n761 B.n464 163.367
R2080 B.n765 B.n763 163.367
R2081 B.n769 B.n462 163.367
R2082 B.n773 B.n771 163.367
R2083 B.n777 B.n460 163.367
R2084 B.n781 B.n779 163.367
R2085 B.n785 B.n458 163.367
R2086 B.n789 B.n787 163.367
R2087 B.n793 B.n456 163.367
R2088 B.n797 B.n795 163.367
R2089 B.n801 B.n448 163.367
R2090 B.n809 B.n448 163.367
R2091 B.n809 B.n446 163.367
R2092 B.n813 B.n446 163.367
R2093 B.n813 B.n440 163.367
R2094 B.n821 B.n440 163.367
R2095 B.n821 B.n438 163.367
R2096 B.n825 B.n438 163.367
R2097 B.n825 B.n432 163.367
R2098 B.n833 B.n432 163.367
R2099 B.n833 B.n430 163.367
R2100 B.n837 B.n430 163.367
R2101 B.n837 B.n424 163.367
R2102 B.n845 B.n424 163.367
R2103 B.n845 B.n422 163.367
R2104 B.n849 B.n422 163.367
R2105 B.n849 B.n416 163.367
R2106 B.n857 B.n416 163.367
R2107 B.n857 B.n414 163.367
R2108 B.n861 B.n414 163.367
R2109 B.n861 B.n407 163.367
R2110 B.n869 B.n407 163.367
R2111 B.n869 B.n405 163.367
R2112 B.n874 B.n405 163.367
R2113 B.n874 B.n400 163.367
R2114 B.n882 B.n400 163.367
R2115 B.n883 B.n882 163.367
R2116 B.n883 B.n5 163.367
R2117 B.n6 B.n5 163.367
R2118 B.n7 B.n6 163.367
R2119 B.n888 B.n7 163.367
R2120 B.n888 B.n12 163.367
R2121 B.n13 B.n12 163.367
R2122 B.n14 B.n13 163.367
R2123 B.n893 B.n14 163.367
R2124 B.n893 B.n19 163.367
R2125 B.n20 B.n19 163.367
R2126 B.n21 B.n20 163.367
R2127 B.n898 B.n21 163.367
R2128 B.n898 B.n26 163.367
R2129 B.n27 B.n26 163.367
R2130 B.n28 B.n27 163.367
R2131 B.n903 B.n28 163.367
R2132 B.n903 B.n33 163.367
R2133 B.n34 B.n33 163.367
R2134 B.n35 B.n34 163.367
R2135 B.n908 B.n35 163.367
R2136 B.n908 B.n40 163.367
R2137 B.n41 B.n40 163.367
R2138 B.n42 B.n41 163.367
R2139 B.n913 B.n42 163.367
R2140 B.n913 B.n47 163.367
R2141 B.n48 B.n47 163.367
R2142 B.n49 B.n48 163.367
R2143 B.n918 B.n49 163.367
R2144 B.n918 B.n54 163.367
R2145 B.n131 B.n130 163.367
R2146 B.n135 B.n134 163.367
R2147 B.n139 B.n138 163.367
R2148 B.n143 B.n142 163.367
R2149 B.n147 B.n146 163.367
R2150 B.n151 B.n150 163.367
R2151 B.n155 B.n154 163.367
R2152 B.n159 B.n158 163.367
R2153 B.n163 B.n162 163.367
R2154 B.n167 B.n166 163.367
R2155 B.n171 B.n170 163.367
R2156 B.n175 B.n174 163.367
R2157 B.n179 B.n178 163.367
R2158 B.n183 B.n182 163.367
R2159 B.n187 B.n186 163.367
R2160 B.n191 B.n190 163.367
R2161 B.n195 B.n194 163.367
R2162 B.n199 B.n198 163.367
R2163 B.n203 B.n202 163.367
R2164 B.n207 B.n206 163.367
R2165 B.n211 B.n210 163.367
R2166 B.n215 B.n214 163.367
R2167 B.n219 B.n218 163.367
R2168 B.n223 B.n222 163.367
R2169 B.n227 B.n226 163.367
R2170 B.n231 B.n230 163.367
R2171 B.n235 B.n234 163.367
R2172 B.n239 B.n238 163.367
R2173 B.n243 B.n242 163.367
R2174 B.n247 B.n246 163.367
R2175 B.n251 B.n250 163.367
R2176 B.n255 B.n254 163.367
R2177 B.n259 B.n258 163.367
R2178 B.n263 B.n262 163.367
R2179 B.n267 B.n266 163.367
R2180 B.n271 B.n270 163.367
R2181 B.n276 B.n275 163.367
R2182 B.n280 B.n279 163.367
R2183 B.n284 B.n283 163.367
R2184 B.n288 B.n287 163.367
R2185 B.n292 B.n291 163.367
R2186 B.n296 B.n295 163.367
R2187 B.n300 B.n299 163.367
R2188 B.n304 B.n303 163.367
R2189 B.n308 B.n307 163.367
R2190 B.n312 B.n311 163.367
R2191 B.n316 B.n315 163.367
R2192 B.n320 B.n319 163.367
R2193 B.n324 B.n323 163.367
R2194 B.n328 B.n327 163.367
R2195 B.n332 B.n331 163.367
R2196 B.n336 B.n335 163.367
R2197 B.n340 B.n339 163.367
R2198 B.n344 B.n343 163.367
R2199 B.n348 B.n347 163.367
R2200 B.n352 B.n351 163.367
R2201 B.n356 B.n355 163.367
R2202 B.n360 B.n359 163.367
R2203 B.n364 B.n363 163.367
R2204 B.n368 B.n367 163.367
R2205 B.n372 B.n371 163.367
R2206 B.n376 B.n375 163.367
R2207 B.n380 B.n379 163.367
R2208 B.n384 B.n383 163.367
R2209 B.n388 B.n387 163.367
R2210 B.n392 B.n391 163.367
R2211 B.n396 B.n395 163.367
R2212 B.n922 B.n123 163.367
R2213 B.n527 B.n452 71.676
R2214 B.n531 B.n530 71.676
R2215 B.n536 B.n535 71.676
R2216 B.n539 B.n538 71.676
R2217 B.n544 B.n543 71.676
R2218 B.n547 B.n546 71.676
R2219 B.n552 B.n551 71.676
R2220 B.n555 B.n554 71.676
R2221 B.n560 B.n559 71.676
R2222 B.n563 B.n562 71.676
R2223 B.n568 B.n567 71.676
R2224 B.n571 B.n570 71.676
R2225 B.n576 B.n575 71.676
R2226 B.n579 B.n578 71.676
R2227 B.n584 B.n583 71.676
R2228 B.n587 B.n586 71.676
R2229 B.n592 B.n591 71.676
R2230 B.n595 B.n594 71.676
R2231 B.n600 B.n599 71.676
R2232 B.n603 B.n602 71.676
R2233 B.n608 B.n607 71.676
R2234 B.n611 B.n610 71.676
R2235 B.n616 B.n615 71.676
R2236 B.n619 B.n618 71.676
R2237 B.n624 B.n623 71.676
R2238 B.n627 B.n626 71.676
R2239 B.n632 B.n631 71.676
R2240 B.n635 B.n634 71.676
R2241 B.n640 B.n639 71.676
R2242 B.n643 B.n642 71.676
R2243 B.n648 B.n647 71.676
R2244 B.n651 B.n650 71.676
R2245 B.n657 B.n656 71.676
R2246 B.n660 B.n659 71.676
R2247 B.n665 B.n664 71.676
R2248 B.n668 B.n667 71.676
R2249 B.n674 B.n673 71.676
R2250 B.n677 B.n676 71.676
R2251 B.n682 B.n681 71.676
R2252 B.n685 B.n684 71.676
R2253 B.n690 B.n689 71.676
R2254 B.n693 B.n692 71.676
R2255 B.n698 B.n697 71.676
R2256 B.n701 B.n700 71.676
R2257 B.n706 B.n705 71.676
R2258 B.n709 B.n708 71.676
R2259 B.n714 B.n713 71.676
R2260 B.n717 B.n716 71.676
R2261 B.n722 B.n721 71.676
R2262 B.n725 B.n724 71.676
R2263 B.n730 B.n729 71.676
R2264 B.n733 B.n732 71.676
R2265 B.n738 B.n737 71.676
R2266 B.n741 B.n740 71.676
R2267 B.n746 B.n745 71.676
R2268 B.n749 B.n748 71.676
R2269 B.n754 B.n753 71.676
R2270 B.n757 B.n756 71.676
R2271 B.n762 B.n761 71.676
R2272 B.n765 B.n764 71.676
R2273 B.n770 B.n769 71.676
R2274 B.n773 B.n772 71.676
R2275 B.n778 B.n777 71.676
R2276 B.n781 B.n780 71.676
R2277 B.n786 B.n785 71.676
R2278 B.n789 B.n788 71.676
R2279 B.n794 B.n793 71.676
R2280 B.n797 B.n796 71.676
R2281 B.n55 B.n53 71.676
R2282 B.n131 B.n56 71.676
R2283 B.n135 B.n57 71.676
R2284 B.n139 B.n58 71.676
R2285 B.n143 B.n59 71.676
R2286 B.n147 B.n60 71.676
R2287 B.n151 B.n61 71.676
R2288 B.n155 B.n62 71.676
R2289 B.n159 B.n63 71.676
R2290 B.n163 B.n64 71.676
R2291 B.n167 B.n65 71.676
R2292 B.n171 B.n66 71.676
R2293 B.n175 B.n67 71.676
R2294 B.n179 B.n68 71.676
R2295 B.n183 B.n69 71.676
R2296 B.n187 B.n70 71.676
R2297 B.n191 B.n71 71.676
R2298 B.n195 B.n72 71.676
R2299 B.n199 B.n73 71.676
R2300 B.n203 B.n74 71.676
R2301 B.n207 B.n75 71.676
R2302 B.n211 B.n76 71.676
R2303 B.n215 B.n77 71.676
R2304 B.n219 B.n78 71.676
R2305 B.n223 B.n79 71.676
R2306 B.n227 B.n80 71.676
R2307 B.n231 B.n81 71.676
R2308 B.n235 B.n82 71.676
R2309 B.n239 B.n83 71.676
R2310 B.n243 B.n84 71.676
R2311 B.n247 B.n85 71.676
R2312 B.n251 B.n86 71.676
R2313 B.n255 B.n87 71.676
R2314 B.n259 B.n88 71.676
R2315 B.n263 B.n89 71.676
R2316 B.n267 B.n90 71.676
R2317 B.n271 B.n91 71.676
R2318 B.n276 B.n92 71.676
R2319 B.n280 B.n93 71.676
R2320 B.n284 B.n94 71.676
R2321 B.n288 B.n95 71.676
R2322 B.n292 B.n96 71.676
R2323 B.n296 B.n97 71.676
R2324 B.n300 B.n98 71.676
R2325 B.n304 B.n99 71.676
R2326 B.n308 B.n100 71.676
R2327 B.n312 B.n101 71.676
R2328 B.n316 B.n102 71.676
R2329 B.n320 B.n103 71.676
R2330 B.n324 B.n104 71.676
R2331 B.n328 B.n105 71.676
R2332 B.n332 B.n106 71.676
R2333 B.n336 B.n107 71.676
R2334 B.n340 B.n108 71.676
R2335 B.n344 B.n109 71.676
R2336 B.n348 B.n110 71.676
R2337 B.n352 B.n111 71.676
R2338 B.n356 B.n112 71.676
R2339 B.n360 B.n113 71.676
R2340 B.n364 B.n114 71.676
R2341 B.n368 B.n115 71.676
R2342 B.n372 B.n116 71.676
R2343 B.n376 B.n117 71.676
R2344 B.n380 B.n118 71.676
R2345 B.n384 B.n119 71.676
R2346 B.n388 B.n120 71.676
R2347 B.n392 B.n121 71.676
R2348 B.n396 B.n122 71.676
R2349 B.n123 B.n122 71.676
R2350 B.n395 B.n121 71.676
R2351 B.n391 B.n120 71.676
R2352 B.n387 B.n119 71.676
R2353 B.n383 B.n118 71.676
R2354 B.n379 B.n117 71.676
R2355 B.n375 B.n116 71.676
R2356 B.n371 B.n115 71.676
R2357 B.n367 B.n114 71.676
R2358 B.n363 B.n113 71.676
R2359 B.n359 B.n112 71.676
R2360 B.n355 B.n111 71.676
R2361 B.n351 B.n110 71.676
R2362 B.n347 B.n109 71.676
R2363 B.n343 B.n108 71.676
R2364 B.n339 B.n107 71.676
R2365 B.n335 B.n106 71.676
R2366 B.n331 B.n105 71.676
R2367 B.n327 B.n104 71.676
R2368 B.n323 B.n103 71.676
R2369 B.n319 B.n102 71.676
R2370 B.n315 B.n101 71.676
R2371 B.n311 B.n100 71.676
R2372 B.n307 B.n99 71.676
R2373 B.n303 B.n98 71.676
R2374 B.n299 B.n97 71.676
R2375 B.n295 B.n96 71.676
R2376 B.n291 B.n95 71.676
R2377 B.n287 B.n94 71.676
R2378 B.n283 B.n93 71.676
R2379 B.n279 B.n92 71.676
R2380 B.n275 B.n91 71.676
R2381 B.n270 B.n90 71.676
R2382 B.n266 B.n89 71.676
R2383 B.n262 B.n88 71.676
R2384 B.n258 B.n87 71.676
R2385 B.n254 B.n86 71.676
R2386 B.n250 B.n85 71.676
R2387 B.n246 B.n84 71.676
R2388 B.n242 B.n83 71.676
R2389 B.n238 B.n82 71.676
R2390 B.n234 B.n81 71.676
R2391 B.n230 B.n80 71.676
R2392 B.n226 B.n79 71.676
R2393 B.n222 B.n78 71.676
R2394 B.n218 B.n77 71.676
R2395 B.n214 B.n76 71.676
R2396 B.n210 B.n75 71.676
R2397 B.n206 B.n74 71.676
R2398 B.n202 B.n73 71.676
R2399 B.n198 B.n72 71.676
R2400 B.n194 B.n71 71.676
R2401 B.n190 B.n70 71.676
R2402 B.n186 B.n69 71.676
R2403 B.n182 B.n68 71.676
R2404 B.n178 B.n67 71.676
R2405 B.n174 B.n66 71.676
R2406 B.n170 B.n65 71.676
R2407 B.n166 B.n64 71.676
R2408 B.n162 B.n63 71.676
R2409 B.n158 B.n62 71.676
R2410 B.n154 B.n61 71.676
R2411 B.n150 B.n60 71.676
R2412 B.n146 B.n59 71.676
R2413 B.n142 B.n58 71.676
R2414 B.n138 B.n57 71.676
R2415 B.n134 B.n56 71.676
R2416 B.n130 B.n55 71.676
R2417 B.n528 B.n527 71.676
R2418 B.n530 B.n524 71.676
R2419 B.n537 B.n536 71.676
R2420 B.n538 B.n522 71.676
R2421 B.n545 B.n544 71.676
R2422 B.n546 B.n520 71.676
R2423 B.n553 B.n552 71.676
R2424 B.n554 B.n518 71.676
R2425 B.n561 B.n560 71.676
R2426 B.n562 B.n516 71.676
R2427 B.n569 B.n568 71.676
R2428 B.n570 B.n514 71.676
R2429 B.n577 B.n576 71.676
R2430 B.n578 B.n512 71.676
R2431 B.n585 B.n584 71.676
R2432 B.n586 B.n510 71.676
R2433 B.n593 B.n592 71.676
R2434 B.n594 B.n508 71.676
R2435 B.n601 B.n600 71.676
R2436 B.n602 B.n506 71.676
R2437 B.n609 B.n608 71.676
R2438 B.n610 B.n504 71.676
R2439 B.n617 B.n616 71.676
R2440 B.n618 B.n502 71.676
R2441 B.n625 B.n624 71.676
R2442 B.n626 B.n500 71.676
R2443 B.n633 B.n632 71.676
R2444 B.n634 B.n498 71.676
R2445 B.n641 B.n640 71.676
R2446 B.n642 B.n496 71.676
R2447 B.n649 B.n648 71.676
R2448 B.n650 B.n492 71.676
R2449 B.n658 B.n657 71.676
R2450 B.n659 B.n490 71.676
R2451 B.n666 B.n665 71.676
R2452 B.n667 B.n486 71.676
R2453 B.n675 B.n674 71.676
R2454 B.n676 B.n484 71.676
R2455 B.n683 B.n682 71.676
R2456 B.n684 B.n482 71.676
R2457 B.n691 B.n690 71.676
R2458 B.n692 B.n480 71.676
R2459 B.n699 B.n698 71.676
R2460 B.n700 B.n478 71.676
R2461 B.n707 B.n706 71.676
R2462 B.n708 B.n476 71.676
R2463 B.n715 B.n714 71.676
R2464 B.n716 B.n474 71.676
R2465 B.n723 B.n722 71.676
R2466 B.n724 B.n472 71.676
R2467 B.n731 B.n730 71.676
R2468 B.n732 B.n470 71.676
R2469 B.n739 B.n738 71.676
R2470 B.n740 B.n468 71.676
R2471 B.n747 B.n746 71.676
R2472 B.n748 B.n466 71.676
R2473 B.n755 B.n754 71.676
R2474 B.n756 B.n464 71.676
R2475 B.n763 B.n762 71.676
R2476 B.n764 B.n462 71.676
R2477 B.n771 B.n770 71.676
R2478 B.n772 B.n460 71.676
R2479 B.n779 B.n778 71.676
R2480 B.n780 B.n458 71.676
R2481 B.n787 B.n786 71.676
R2482 B.n788 B.n456 71.676
R2483 B.n795 B.n794 71.676
R2484 B.n796 B.n454 71.676
R2485 B.n671 B.n488 59.5399
R2486 B.n653 B.n494 59.5399
R2487 B.n128 B.n127 59.5399
R2488 B.n273 B.n125 59.5399
R2489 B.n802 B.n453 50.9983
R2490 B.n924 B.n923 50.9983
R2491 B.n488 B.n487 43.4429
R2492 B.n494 B.n493 43.4429
R2493 B.n127 B.n126 43.4429
R2494 B.n125 B.n124 43.4429
R2495 B.n926 B.n52 31.6883
R2496 B.n921 B.n920 31.6883
R2497 B.n800 B.n799 31.6883
R2498 B.n804 B.n451 31.6883
R2499 B.n802 B.n449 30.1557
R2500 B.n808 B.n449 30.1557
R2501 B.n808 B.n445 30.1557
R2502 B.n814 B.n445 30.1557
R2503 B.n814 B.n441 30.1557
R2504 B.n820 B.n441 30.1557
R2505 B.n826 B.n437 30.1557
R2506 B.n826 B.n433 30.1557
R2507 B.n832 B.n433 30.1557
R2508 B.n832 B.n429 30.1557
R2509 B.n838 B.n429 30.1557
R2510 B.n838 B.n425 30.1557
R2511 B.n844 B.n425 30.1557
R2512 B.n844 B.n421 30.1557
R2513 B.n850 B.n421 30.1557
R2514 B.n856 B.n417 30.1557
R2515 B.n856 B.n413 30.1557
R2516 B.n862 B.n413 30.1557
R2517 B.n862 B.n408 30.1557
R2518 B.n868 B.n408 30.1557
R2519 B.n868 B.n409 30.1557
R2520 B.n875 B.n401 30.1557
R2521 B.n881 B.n401 30.1557
R2522 B.n881 B.n4 30.1557
R2523 B.n980 B.n4 30.1557
R2524 B.n980 B.n979 30.1557
R2525 B.n979 B.n978 30.1557
R2526 B.n978 B.n8 30.1557
R2527 B.n972 B.n8 30.1557
R2528 B.n971 B.n970 30.1557
R2529 B.n970 B.n15 30.1557
R2530 B.n964 B.n15 30.1557
R2531 B.n964 B.n963 30.1557
R2532 B.n963 B.n962 30.1557
R2533 B.n962 B.n22 30.1557
R2534 B.n956 B.n955 30.1557
R2535 B.n955 B.n954 30.1557
R2536 B.n954 B.n29 30.1557
R2537 B.n948 B.n29 30.1557
R2538 B.n948 B.n947 30.1557
R2539 B.n947 B.n946 30.1557
R2540 B.n946 B.n36 30.1557
R2541 B.n940 B.n36 30.1557
R2542 B.n940 B.n939 30.1557
R2543 B.n938 B.n43 30.1557
R2544 B.n932 B.n43 30.1557
R2545 B.n932 B.n931 30.1557
R2546 B.n931 B.n930 30.1557
R2547 B.n930 B.n50 30.1557
R2548 B.n924 B.n50 30.1557
R2549 B.n875 B.t1 27.0515
R2550 B.n972 B.t2 27.0515
R2551 B.n820 B.t5 21.73
R2552 B.t12 B.n938 21.73
R2553 B B.n982 18.0485
R2554 B.n850 B.t3 15.5216
R2555 B.n956 B.t0 15.5216
R2556 B.t3 B.n417 14.6346
R2557 B.t0 B.n22 14.6346
R2558 B.n129 B.n52 10.6151
R2559 B.n132 B.n129 10.6151
R2560 B.n133 B.n132 10.6151
R2561 B.n136 B.n133 10.6151
R2562 B.n137 B.n136 10.6151
R2563 B.n140 B.n137 10.6151
R2564 B.n141 B.n140 10.6151
R2565 B.n144 B.n141 10.6151
R2566 B.n145 B.n144 10.6151
R2567 B.n148 B.n145 10.6151
R2568 B.n149 B.n148 10.6151
R2569 B.n152 B.n149 10.6151
R2570 B.n153 B.n152 10.6151
R2571 B.n156 B.n153 10.6151
R2572 B.n157 B.n156 10.6151
R2573 B.n160 B.n157 10.6151
R2574 B.n161 B.n160 10.6151
R2575 B.n164 B.n161 10.6151
R2576 B.n165 B.n164 10.6151
R2577 B.n168 B.n165 10.6151
R2578 B.n169 B.n168 10.6151
R2579 B.n172 B.n169 10.6151
R2580 B.n173 B.n172 10.6151
R2581 B.n176 B.n173 10.6151
R2582 B.n177 B.n176 10.6151
R2583 B.n180 B.n177 10.6151
R2584 B.n181 B.n180 10.6151
R2585 B.n184 B.n181 10.6151
R2586 B.n185 B.n184 10.6151
R2587 B.n188 B.n185 10.6151
R2588 B.n189 B.n188 10.6151
R2589 B.n192 B.n189 10.6151
R2590 B.n193 B.n192 10.6151
R2591 B.n196 B.n193 10.6151
R2592 B.n197 B.n196 10.6151
R2593 B.n200 B.n197 10.6151
R2594 B.n201 B.n200 10.6151
R2595 B.n204 B.n201 10.6151
R2596 B.n205 B.n204 10.6151
R2597 B.n208 B.n205 10.6151
R2598 B.n209 B.n208 10.6151
R2599 B.n212 B.n209 10.6151
R2600 B.n213 B.n212 10.6151
R2601 B.n216 B.n213 10.6151
R2602 B.n217 B.n216 10.6151
R2603 B.n220 B.n217 10.6151
R2604 B.n221 B.n220 10.6151
R2605 B.n224 B.n221 10.6151
R2606 B.n225 B.n224 10.6151
R2607 B.n228 B.n225 10.6151
R2608 B.n229 B.n228 10.6151
R2609 B.n232 B.n229 10.6151
R2610 B.n233 B.n232 10.6151
R2611 B.n236 B.n233 10.6151
R2612 B.n237 B.n236 10.6151
R2613 B.n240 B.n237 10.6151
R2614 B.n241 B.n240 10.6151
R2615 B.n244 B.n241 10.6151
R2616 B.n245 B.n244 10.6151
R2617 B.n248 B.n245 10.6151
R2618 B.n249 B.n248 10.6151
R2619 B.n252 B.n249 10.6151
R2620 B.n253 B.n252 10.6151
R2621 B.n257 B.n256 10.6151
R2622 B.n260 B.n257 10.6151
R2623 B.n261 B.n260 10.6151
R2624 B.n264 B.n261 10.6151
R2625 B.n265 B.n264 10.6151
R2626 B.n268 B.n265 10.6151
R2627 B.n269 B.n268 10.6151
R2628 B.n272 B.n269 10.6151
R2629 B.n277 B.n274 10.6151
R2630 B.n278 B.n277 10.6151
R2631 B.n281 B.n278 10.6151
R2632 B.n282 B.n281 10.6151
R2633 B.n285 B.n282 10.6151
R2634 B.n286 B.n285 10.6151
R2635 B.n289 B.n286 10.6151
R2636 B.n290 B.n289 10.6151
R2637 B.n293 B.n290 10.6151
R2638 B.n294 B.n293 10.6151
R2639 B.n297 B.n294 10.6151
R2640 B.n298 B.n297 10.6151
R2641 B.n301 B.n298 10.6151
R2642 B.n302 B.n301 10.6151
R2643 B.n305 B.n302 10.6151
R2644 B.n306 B.n305 10.6151
R2645 B.n309 B.n306 10.6151
R2646 B.n310 B.n309 10.6151
R2647 B.n313 B.n310 10.6151
R2648 B.n314 B.n313 10.6151
R2649 B.n317 B.n314 10.6151
R2650 B.n318 B.n317 10.6151
R2651 B.n321 B.n318 10.6151
R2652 B.n322 B.n321 10.6151
R2653 B.n325 B.n322 10.6151
R2654 B.n326 B.n325 10.6151
R2655 B.n329 B.n326 10.6151
R2656 B.n330 B.n329 10.6151
R2657 B.n333 B.n330 10.6151
R2658 B.n334 B.n333 10.6151
R2659 B.n337 B.n334 10.6151
R2660 B.n338 B.n337 10.6151
R2661 B.n341 B.n338 10.6151
R2662 B.n342 B.n341 10.6151
R2663 B.n345 B.n342 10.6151
R2664 B.n346 B.n345 10.6151
R2665 B.n349 B.n346 10.6151
R2666 B.n350 B.n349 10.6151
R2667 B.n353 B.n350 10.6151
R2668 B.n354 B.n353 10.6151
R2669 B.n357 B.n354 10.6151
R2670 B.n358 B.n357 10.6151
R2671 B.n361 B.n358 10.6151
R2672 B.n362 B.n361 10.6151
R2673 B.n365 B.n362 10.6151
R2674 B.n366 B.n365 10.6151
R2675 B.n369 B.n366 10.6151
R2676 B.n370 B.n369 10.6151
R2677 B.n373 B.n370 10.6151
R2678 B.n374 B.n373 10.6151
R2679 B.n377 B.n374 10.6151
R2680 B.n378 B.n377 10.6151
R2681 B.n381 B.n378 10.6151
R2682 B.n382 B.n381 10.6151
R2683 B.n385 B.n382 10.6151
R2684 B.n386 B.n385 10.6151
R2685 B.n389 B.n386 10.6151
R2686 B.n390 B.n389 10.6151
R2687 B.n393 B.n390 10.6151
R2688 B.n394 B.n393 10.6151
R2689 B.n397 B.n394 10.6151
R2690 B.n398 B.n397 10.6151
R2691 B.n921 B.n398 10.6151
R2692 B.n800 B.n447 10.6151
R2693 B.n810 B.n447 10.6151
R2694 B.n811 B.n810 10.6151
R2695 B.n812 B.n811 10.6151
R2696 B.n812 B.n439 10.6151
R2697 B.n822 B.n439 10.6151
R2698 B.n823 B.n822 10.6151
R2699 B.n824 B.n823 10.6151
R2700 B.n824 B.n431 10.6151
R2701 B.n834 B.n431 10.6151
R2702 B.n835 B.n834 10.6151
R2703 B.n836 B.n835 10.6151
R2704 B.n836 B.n423 10.6151
R2705 B.n846 B.n423 10.6151
R2706 B.n847 B.n846 10.6151
R2707 B.n848 B.n847 10.6151
R2708 B.n848 B.n415 10.6151
R2709 B.n858 B.n415 10.6151
R2710 B.n859 B.n858 10.6151
R2711 B.n860 B.n859 10.6151
R2712 B.n860 B.n406 10.6151
R2713 B.n870 B.n406 10.6151
R2714 B.n871 B.n870 10.6151
R2715 B.n873 B.n871 10.6151
R2716 B.n873 B.n872 10.6151
R2717 B.n872 B.n399 10.6151
R2718 B.n884 B.n399 10.6151
R2719 B.n885 B.n884 10.6151
R2720 B.n886 B.n885 10.6151
R2721 B.n887 B.n886 10.6151
R2722 B.n889 B.n887 10.6151
R2723 B.n890 B.n889 10.6151
R2724 B.n891 B.n890 10.6151
R2725 B.n892 B.n891 10.6151
R2726 B.n894 B.n892 10.6151
R2727 B.n895 B.n894 10.6151
R2728 B.n896 B.n895 10.6151
R2729 B.n897 B.n896 10.6151
R2730 B.n899 B.n897 10.6151
R2731 B.n900 B.n899 10.6151
R2732 B.n901 B.n900 10.6151
R2733 B.n902 B.n901 10.6151
R2734 B.n904 B.n902 10.6151
R2735 B.n905 B.n904 10.6151
R2736 B.n906 B.n905 10.6151
R2737 B.n907 B.n906 10.6151
R2738 B.n909 B.n907 10.6151
R2739 B.n910 B.n909 10.6151
R2740 B.n911 B.n910 10.6151
R2741 B.n912 B.n911 10.6151
R2742 B.n914 B.n912 10.6151
R2743 B.n915 B.n914 10.6151
R2744 B.n916 B.n915 10.6151
R2745 B.n917 B.n916 10.6151
R2746 B.n919 B.n917 10.6151
R2747 B.n920 B.n919 10.6151
R2748 B.n526 B.n451 10.6151
R2749 B.n526 B.n525 10.6151
R2750 B.n532 B.n525 10.6151
R2751 B.n533 B.n532 10.6151
R2752 B.n534 B.n533 10.6151
R2753 B.n534 B.n523 10.6151
R2754 B.n540 B.n523 10.6151
R2755 B.n541 B.n540 10.6151
R2756 B.n542 B.n541 10.6151
R2757 B.n542 B.n521 10.6151
R2758 B.n548 B.n521 10.6151
R2759 B.n549 B.n548 10.6151
R2760 B.n550 B.n549 10.6151
R2761 B.n550 B.n519 10.6151
R2762 B.n556 B.n519 10.6151
R2763 B.n557 B.n556 10.6151
R2764 B.n558 B.n557 10.6151
R2765 B.n558 B.n517 10.6151
R2766 B.n564 B.n517 10.6151
R2767 B.n565 B.n564 10.6151
R2768 B.n566 B.n565 10.6151
R2769 B.n566 B.n515 10.6151
R2770 B.n572 B.n515 10.6151
R2771 B.n573 B.n572 10.6151
R2772 B.n574 B.n573 10.6151
R2773 B.n574 B.n513 10.6151
R2774 B.n580 B.n513 10.6151
R2775 B.n581 B.n580 10.6151
R2776 B.n582 B.n581 10.6151
R2777 B.n582 B.n511 10.6151
R2778 B.n588 B.n511 10.6151
R2779 B.n589 B.n588 10.6151
R2780 B.n590 B.n589 10.6151
R2781 B.n590 B.n509 10.6151
R2782 B.n596 B.n509 10.6151
R2783 B.n597 B.n596 10.6151
R2784 B.n598 B.n597 10.6151
R2785 B.n598 B.n507 10.6151
R2786 B.n604 B.n507 10.6151
R2787 B.n605 B.n604 10.6151
R2788 B.n606 B.n605 10.6151
R2789 B.n606 B.n505 10.6151
R2790 B.n612 B.n505 10.6151
R2791 B.n613 B.n612 10.6151
R2792 B.n614 B.n613 10.6151
R2793 B.n614 B.n503 10.6151
R2794 B.n620 B.n503 10.6151
R2795 B.n621 B.n620 10.6151
R2796 B.n622 B.n621 10.6151
R2797 B.n622 B.n501 10.6151
R2798 B.n628 B.n501 10.6151
R2799 B.n629 B.n628 10.6151
R2800 B.n630 B.n629 10.6151
R2801 B.n630 B.n499 10.6151
R2802 B.n636 B.n499 10.6151
R2803 B.n637 B.n636 10.6151
R2804 B.n638 B.n637 10.6151
R2805 B.n638 B.n497 10.6151
R2806 B.n644 B.n497 10.6151
R2807 B.n645 B.n644 10.6151
R2808 B.n646 B.n645 10.6151
R2809 B.n646 B.n495 10.6151
R2810 B.n652 B.n495 10.6151
R2811 B.n655 B.n654 10.6151
R2812 B.n655 B.n491 10.6151
R2813 B.n661 B.n491 10.6151
R2814 B.n662 B.n661 10.6151
R2815 B.n663 B.n662 10.6151
R2816 B.n663 B.n489 10.6151
R2817 B.n669 B.n489 10.6151
R2818 B.n670 B.n669 10.6151
R2819 B.n672 B.n485 10.6151
R2820 B.n678 B.n485 10.6151
R2821 B.n679 B.n678 10.6151
R2822 B.n680 B.n679 10.6151
R2823 B.n680 B.n483 10.6151
R2824 B.n686 B.n483 10.6151
R2825 B.n687 B.n686 10.6151
R2826 B.n688 B.n687 10.6151
R2827 B.n688 B.n481 10.6151
R2828 B.n694 B.n481 10.6151
R2829 B.n695 B.n694 10.6151
R2830 B.n696 B.n695 10.6151
R2831 B.n696 B.n479 10.6151
R2832 B.n702 B.n479 10.6151
R2833 B.n703 B.n702 10.6151
R2834 B.n704 B.n703 10.6151
R2835 B.n704 B.n477 10.6151
R2836 B.n710 B.n477 10.6151
R2837 B.n711 B.n710 10.6151
R2838 B.n712 B.n711 10.6151
R2839 B.n712 B.n475 10.6151
R2840 B.n718 B.n475 10.6151
R2841 B.n719 B.n718 10.6151
R2842 B.n720 B.n719 10.6151
R2843 B.n720 B.n473 10.6151
R2844 B.n726 B.n473 10.6151
R2845 B.n727 B.n726 10.6151
R2846 B.n728 B.n727 10.6151
R2847 B.n728 B.n471 10.6151
R2848 B.n734 B.n471 10.6151
R2849 B.n735 B.n734 10.6151
R2850 B.n736 B.n735 10.6151
R2851 B.n736 B.n469 10.6151
R2852 B.n742 B.n469 10.6151
R2853 B.n743 B.n742 10.6151
R2854 B.n744 B.n743 10.6151
R2855 B.n744 B.n467 10.6151
R2856 B.n750 B.n467 10.6151
R2857 B.n751 B.n750 10.6151
R2858 B.n752 B.n751 10.6151
R2859 B.n752 B.n465 10.6151
R2860 B.n758 B.n465 10.6151
R2861 B.n759 B.n758 10.6151
R2862 B.n760 B.n759 10.6151
R2863 B.n760 B.n463 10.6151
R2864 B.n766 B.n463 10.6151
R2865 B.n767 B.n766 10.6151
R2866 B.n768 B.n767 10.6151
R2867 B.n768 B.n461 10.6151
R2868 B.n774 B.n461 10.6151
R2869 B.n775 B.n774 10.6151
R2870 B.n776 B.n775 10.6151
R2871 B.n776 B.n459 10.6151
R2872 B.n782 B.n459 10.6151
R2873 B.n783 B.n782 10.6151
R2874 B.n784 B.n783 10.6151
R2875 B.n784 B.n457 10.6151
R2876 B.n790 B.n457 10.6151
R2877 B.n791 B.n790 10.6151
R2878 B.n792 B.n791 10.6151
R2879 B.n792 B.n455 10.6151
R2880 B.n798 B.n455 10.6151
R2881 B.n799 B.n798 10.6151
R2882 B.n805 B.n804 10.6151
R2883 B.n806 B.n805 10.6151
R2884 B.n806 B.n443 10.6151
R2885 B.n816 B.n443 10.6151
R2886 B.n817 B.n816 10.6151
R2887 B.n818 B.n817 10.6151
R2888 B.n818 B.n435 10.6151
R2889 B.n828 B.n435 10.6151
R2890 B.n829 B.n828 10.6151
R2891 B.n830 B.n829 10.6151
R2892 B.n830 B.n427 10.6151
R2893 B.n840 B.n427 10.6151
R2894 B.n841 B.n840 10.6151
R2895 B.n842 B.n841 10.6151
R2896 B.n842 B.n419 10.6151
R2897 B.n852 B.n419 10.6151
R2898 B.n853 B.n852 10.6151
R2899 B.n854 B.n853 10.6151
R2900 B.n854 B.n411 10.6151
R2901 B.n864 B.n411 10.6151
R2902 B.n865 B.n864 10.6151
R2903 B.n866 B.n865 10.6151
R2904 B.n866 B.n403 10.6151
R2905 B.n877 B.n403 10.6151
R2906 B.n878 B.n877 10.6151
R2907 B.n879 B.n878 10.6151
R2908 B.n879 B.n0 10.6151
R2909 B.n976 B.n1 10.6151
R2910 B.n976 B.n975 10.6151
R2911 B.n975 B.n974 10.6151
R2912 B.n974 B.n10 10.6151
R2913 B.n968 B.n10 10.6151
R2914 B.n968 B.n967 10.6151
R2915 B.n967 B.n966 10.6151
R2916 B.n966 B.n17 10.6151
R2917 B.n960 B.n17 10.6151
R2918 B.n960 B.n959 10.6151
R2919 B.n959 B.n958 10.6151
R2920 B.n958 B.n24 10.6151
R2921 B.n952 B.n24 10.6151
R2922 B.n952 B.n951 10.6151
R2923 B.n951 B.n950 10.6151
R2924 B.n950 B.n31 10.6151
R2925 B.n944 B.n31 10.6151
R2926 B.n944 B.n943 10.6151
R2927 B.n943 B.n942 10.6151
R2928 B.n942 B.n38 10.6151
R2929 B.n936 B.n38 10.6151
R2930 B.n936 B.n935 10.6151
R2931 B.n935 B.n934 10.6151
R2932 B.n934 B.n45 10.6151
R2933 B.n928 B.n45 10.6151
R2934 B.n928 B.n927 10.6151
R2935 B.n927 B.n926 10.6151
R2936 B.t5 B.n437 8.42622
R2937 B.n939 B.t12 8.42622
R2938 B.n256 B.n128 6.5566
R2939 B.n273 B.n272 6.5566
R2940 B.n654 B.n653 6.5566
R2941 B.n671 B.n670 6.5566
R2942 B.n253 B.n128 4.05904
R2943 B.n274 B.n273 4.05904
R2944 B.n653 B.n652 4.05904
R2945 B.n672 B.n671 4.05904
R2946 B.n409 B.t1 3.10471
R2947 B.t2 B.n971 3.10471
R2948 B.n982 B.n0 2.81026
R2949 B.n982 B.n1 2.81026
R2950 VN.n0 VN.t0 281.479
R2951 VN.n1 VN.t2 281.479
R2952 VN.n0 VN.t1 280.962
R2953 VN.n1 VN.t3 280.962
R2954 VN VN.n1 57.701
R2955 VN VN.n0 7.62148
R2956 VDD2.n2 VDD2.n0 110.618
R2957 VDD2.n2 VDD2.n1 64.2744
R2958 VDD2.n1 VDD2.t0 1.01432
R2959 VDD2.n1 VDD2.t1 1.01432
R2960 VDD2.n0 VDD2.t3 1.01432
R2961 VDD2.n0 VDD2.t2 1.01432
R2962 VDD2 VDD2.n2 0.0586897
C0 VTAIL VDD1 7.42601f
C1 VN VTAIL 6.56727f
C2 VDD1 VDD2 0.8613f
C3 VN VDD2 7.05954f
C4 VTAIL VDD2 7.47559f
C5 VP VDD1 7.261f
C6 VN VP 7.09235f
C7 VTAIL VP 6.58138f
C8 VP VDD2 0.350524f
C9 VN VDD1 0.148501f
C10 VDD2 B 3.965792f
C11 VDD1 B 8.670111f
C12 VTAIL B 14.138347f
C13 VN B 10.19354f
C14 VP B 7.99093f
C15 VDD2.t3 B 0.409839f
C16 VDD2.t2 B 0.409839f
C17 VDD2.n0 B 4.63849f
C18 VDD2.t0 B 0.409839f
C19 VDD2.t1 B 0.409839f
C20 VDD2.n1 B 3.75537f
C21 VDD2.n2 B 4.39583f
C22 VN.t0 B 3.18623f
C23 VN.t1 B 3.18399f
C24 VN.n0 B 2.17694f
C25 VN.t2 B 3.18623f
C26 VN.t3 B 3.18399f
C27 VN.n1 B 3.77585f
C28 VTAIL.n0 B 0.021059f
C29 VTAIL.n1 B 0.015002f
C30 VTAIL.n2 B 0.008062f
C31 VTAIL.n3 B 0.019055f
C32 VTAIL.n4 B 0.008536f
C33 VTAIL.n5 B 0.015002f
C34 VTAIL.n6 B 0.008062f
C35 VTAIL.n7 B 0.019055f
C36 VTAIL.n8 B 0.008536f
C37 VTAIL.n9 B 0.015002f
C38 VTAIL.n10 B 0.008062f
C39 VTAIL.n11 B 0.019055f
C40 VTAIL.n12 B 0.008536f
C41 VTAIL.n13 B 0.015002f
C42 VTAIL.n14 B 0.008062f
C43 VTAIL.n15 B 0.019055f
C44 VTAIL.n16 B 0.008536f
C45 VTAIL.n17 B 0.015002f
C46 VTAIL.n18 B 0.008062f
C47 VTAIL.n19 B 0.019055f
C48 VTAIL.n20 B 0.008536f
C49 VTAIL.n21 B 0.015002f
C50 VTAIL.n22 B 0.008062f
C51 VTAIL.n23 B 0.019055f
C52 VTAIL.n24 B 0.008536f
C53 VTAIL.n25 B 0.015002f
C54 VTAIL.n26 B 0.008062f
C55 VTAIL.n27 B 0.019055f
C56 VTAIL.n28 B 0.008536f
C57 VTAIL.n29 B 0.015002f
C58 VTAIL.n30 B 0.008062f
C59 VTAIL.n31 B 0.019055f
C60 VTAIL.n32 B 0.008536f
C61 VTAIL.n33 B 0.151534f
C62 VTAIL.t2 B 0.03279f
C63 VTAIL.n34 B 0.014291f
C64 VTAIL.n35 B 0.01347f
C65 VTAIL.n36 B 0.008062f
C66 VTAIL.n37 B 1.2593f
C67 VTAIL.n38 B 0.015002f
C68 VTAIL.n39 B 0.008062f
C69 VTAIL.n40 B 0.008536f
C70 VTAIL.n41 B 0.019055f
C71 VTAIL.n42 B 0.019055f
C72 VTAIL.n43 B 0.008536f
C73 VTAIL.n44 B 0.008062f
C74 VTAIL.n45 B 0.015002f
C75 VTAIL.n46 B 0.015002f
C76 VTAIL.n47 B 0.008062f
C77 VTAIL.n48 B 0.008536f
C78 VTAIL.n49 B 0.019055f
C79 VTAIL.n50 B 0.019055f
C80 VTAIL.n51 B 0.019055f
C81 VTAIL.n52 B 0.008536f
C82 VTAIL.n53 B 0.008062f
C83 VTAIL.n54 B 0.015002f
C84 VTAIL.n55 B 0.015002f
C85 VTAIL.n56 B 0.008062f
C86 VTAIL.n57 B 0.008299f
C87 VTAIL.n58 B 0.008299f
C88 VTAIL.n59 B 0.019055f
C89 VTAIL.n60 B 0.019055f
C90 VTAIL.n61 B 0.008536f
C91 VTAIL.n62 B 0.008062f
C92 VTAIL.n63 B 0.015002f
C93 VTAIL.n64 B 0.015002f
C94 VTAIL.n65 B 0.008062f
C95 VTAIL.n66 B 0.008536f
C96 VTAIL.n67 B 0.019055f
C97 VTAIL.n68 B 0.019055f
C98 VTAIL.n69 B 0.008536f
C99 VTAIL.n70 B 0.008062f
C100 VTAIL.n71 B 0.015002f
C101 VTAIL.n72 B 0.015002f
C102 VTAIL.n73 B 0.008062f
C103 VTAIL.n74 B 0.008536f
C104 VTAIL.n75 B 0.019055f
C105 VTAIL.n76 B 0.019055f
C106 VTAIL.n77 B 0.008536f
C107 VTAIL.n78 B 0.008062f
C108 VTAIL.n79 B 0.015002f
C109 VTAIL.n80 B 0.015002f
C110 VTAIL.n81 B 0.008062f
C111 VTAIL.n82 B 0.008536f
C112 VTAIL.n83 B 0.019055f
C113 VTAIL.n84 B 0.019055f
C114 VTAIL.n85 B 0.008536f
C115 VTAIL.n86 B 0.008062f
C116 VTAIL.n87 B 0.015002f
C117 VTAIL.n88 B 0.015002f
C118 VTAIL.n89 B 0.008062f
C119 VTAIL.n90 B 0.008536f
C120 VTAIL.n91 B 0.019055f
C121 VTAIL.n92 B 0.019055f
C122 VTAIL.n93 B 0.008536f
C123 VTAIL.n94 B 0.008062f
C124 VTAIL.n95 B 0.015002f
C125 VTAIL.n96 B 0.015002f
C126 VTAIL.n97 B 0.008062f
C127 VTAIL.n98 B 0.008536f
C128 VTAIL.n99 B 0.019055f
C129 VTAIL.n100 B 0.03954f
C130 VTAIL.n101 B 0.008536f
C131 VTAIL.n102 B 0.015763f
C132 VTAIL.n103 B 0.038981f
C133 VTAIL.n104 B 0.041567f
C134 VTAIL.n105 B 0.087447f
C135 VTAIL.n106 B 0.021059f
C136 VTAIL.n107 B 0.015002f
C137 VTAIL.n108 B 0.008062f
C138 VTAIL.n109 B 0.019055f
C139 VTAIL.n110 B 0.008536f
C140 VTAIL.n111 B 0.015002f
C141 VTAIL.n112 B 0.008062f
C142 VTAIL.n113 B 0.019055f
C143 VTAIL.n114 B 0.008536f
C144 VTAIL.n115 B 0.015002f
C145 VTAIL.n116 B 0.008062f
C146 VTAIL.n117 B 0.019055f
C147 VTAIL.n118 B 0.008536f
C148 VTAIL.n119 B 0.015002f
C149 VTAIL.n120 B 0.008062f
C150 VTAIL.n121 B 0.019055f
C151 VTAIL.n122 B 0.008536f
C152 VTAIL.n123 B 0.015002f
C153 VTAIL.n124 B 0.008062f
C154 VTAIL.n125 B 0.019055f
C155 VTAIL.n126 B 0.008536f
C156 VTAIL.n127 B 0.015002f
C157 VTAIL.n128 B 0.008062f
C158 VTAIL.n129 B 0.019055f
C159 VTAIL.n130 B 0.008536f
C160 VTAIL.n131 B 0.015002f
C161 VTAIL.n132 B 0.008062f
C162 VTAIL.n133 B 0.019055f
C163 VTAIL.n134 B 0.008536f
C164 VTAIL.n135 B 0.015002f
C165 VTAIL.n136 B 0.008062f
C166 VTAIL.n137 B 0.019055f
C167 VTAIL.n138 B 0.008536f
C168 VTAIL.n139 B 0.151534f
C169 VTAIL.t5 B 0.03279f
C170 VTAIL.n140 B 0.014291f
C171 VTAIL.n141 B 0.01347f
C172 VTAIL.n142 B 0.008062f
C173 VTAIL.n143 B 1.2593f
C174 VTAIL.n144 B 0.015002f
C175 VTAIL.n145 B 0.008062f
C176 VTAIL.n146 B 0.008536f
C177 VTAIL.n147 B 0.019055f
C178 VTAIL.n148 B 0.019055f
C179 VTAIL.n149 B 0.008536f
C180 VTAIL.n150 B 0.008062f
C181 VTAIL.n151 B 0.015002f
C182 VTAIL.n152 B 0.015002f
C183 VTAIL.n153 B 0.008062f
C184 VTAIL.n154 B 0.008536f
C185 VTAIL.n155 B 0.019055f
C186 VTAIL.n156 B 0.019055f
C187 VTAIL.n157 B 0.019055f
C188 VTAIL.n158 B 0.008536f
C189 VTAIL.n159 B 0.008062f
C190 VTAIL.n160 B 0.015002f
C191 VTAIL.n161 B 0.015002f
C192 VTAIL.n162 B 0.008062f
C193 VTAIL.n163 B 0.008299f
C194 VTAIL.n164 B 0.008299f
C195 VTAIL.n165 B 0.019055f
C196 VTAIL.n166 B 0.019055f
C197 VTAIL.n167 B 0.008536f
C198 VTAIL.n168 B 0.008062f
C199 VTAIL.n169 B 0.015002f
C200 VTAIL.n170 B 0.015002f
C201 VTAIL.n171 B 0.008062f
C202 VTAIL.n172 B 0.008536f
C203 VTAIL.n173 B 0.019055f
C204 VTAIL.n174 B 0.019055f
C205 VTAIL.n175 B 0.008536f
C206 VTAIL.n176 B 0.008062f
C207 VTAIL.n177 B 0.015002f
C208 VTAIL.n178 B 0.015002f
C209 VTAIL.n179 B 0.008062f
C210 VTAIL.n180 B 0.008536f
C211 VTAIL.n181 B 0.019055f
C212 VTAIL.n182 B 0.019055f
C213 VTAIL.n183 B 0.008536f
C214 VTAIL.n184 B 0.008062f
C215 VTAIL.n185 B 0.015002f
C216 VTAIL.n186 B 0.015002f
C217 VTAIL.n187 B 0.008062f
C218 VTAIL.n188 B 0.008536f
C219 VTAIL.n189 B 0.019055f
C220 VTAIL.n190 B 0.019055f
C221 VTAIL.n191 B 0.008536f
C222 VTAIL.n192 B 0.008062f
C223 VTAIL.n193 B 0.015002f
C224 VTAIL.n194 B 0.015002f
C225 VTAIL.n195 B 0.008062f
C226 VTAIL.n196 B 0.008536f
C227 VTAIL.n197 B 0.019055f
C228 VTAIL.n198 B 0.019055f
C229 VTAIL.n199 B 0.008536f
C230 VTAIL.n200 B 0.008062f
C231 VTAIL.n201 B 0.015002f
C232 VTAIL.n202 B 0.015002f
C233 VTAIL.n203 B 0.008062f
C234 VTAIL.n204 B 0.008536f
C235 VTAIL.n205 B 0.019055f
C236 VTAIL.n206 B 0.03954f
C237 VTAIL.n207 B 0.008536f
C238 VTAIL.n208 B 0.015763f
C239 VTAIL.n209 B 0.038981f
C240 VTAIL.n210 B 0.041567f
C241 VTAIL.n211 B 0.131308f
C242 VTAIL.n212 B 0.021059f
C243 VTAIL.n213 B 0.015002f
C244 VTAIL.n214 B 0.008062f
C245 VTAIL.n215 B 0.019055f
C246 VTAIL.n216 B 0.008536f
C247 VTAIL.n217 B 0.015002f
C248 VTAIL.n218 B 0.008062f
C249 VTAIL.n219 B 0.019055f
C250 VTAIL.n220 B 0.008536f
C251 VTAIL.n221 B 0.015002f
C252 VTAIL.n222 B 0.008062f
C253 VTAIL.n223 B 0.019055f
C254 VTAIL.n224 B 0.008536f
C255 VTAIL.n225 B 0.015002f
C256 VTAIL.n226 B 0.008062f
C257 VTAIL.n227 B 0.019055f
C258 VTAIL.n228 B 0.008536f
C259 VTAIL.n229 B 0.015002f
C260 VTAIL.n230 B 0.008062f
C261 VTAIL.n231 B 0.019055f
C262 VTAIL.n232 B 0.008536f
C263 VTAIL.n233 B 0.015002f
C264 VTAIL.n234 B 0.008062f
C265 VTAIL.n235 B 0.019055f
C266 VTAIL.n236 B 0.008536f
C267 VTAIL.n237 B 0.015002f
C268 VTAIL.n238 B 0.008062f
C269 VTAIL.n239 B 0.019055f
C270 VTAIL.n240 B 0.008536f
C271 VTAIL.n241 B 0.015002f
C272 VTAIL.n242 B 0.008062f
C273 VTAIL.n243 B 0.019055f
C274 VTAIL.n244 B 0.008536f
C275 VTAIL.n245 B 0.151534f
C276 VTAIL.t4 B 0.03279f
C277 VTAIL.n246 B 0.014291f
C278 VTAIL.n247 B 0.01347f
C279 VTAIL.n248 B 0.008062f
C280 VTAIL.n249 B 1.2593f
C281 VTAIL.n250 B 0.015002f
C282 VTAIL.n251 B 0.008062f
C283 VTAIL.n252 B 0.008536f
C284 VTAIL.n253 B 0.019055f
C285 VTAIL.n254 B 0.019055f
C286 VTAIL.n255 B 0.008536f
C287 VTAIL.n256 B 0.008062f
C288 VTAIL.n257 B 0.015002f
C289 VTAIL.n258 B 0.015002f
C290 VTAIL.n259 B 0.008062f
C291 VTAIL.n260 B 0.008536f
C292 VTAIL.n261 B 0.019055f
C293 VTAIL.n262 B 0.019055f
C294 VTAIL.n263 B 0.019055f
C295 VTAIL.n264 B 0.008536f
C296 VTAIL.n265 B 0.008062f
C297 VTAIL.n266 B 0.015002f
C298 VTAIL.n267 B 0.015002f
C299 VTAIL.n268 B 0.008062f
C300 VTAIL.n269 B 0.008299f
C301 VTAIL.n270 B 0.008299f
C302 VTAIL.n271 B 0.019055f
C303 VTAIL.n272 B 0.019055f
C304 VTAIL.n273 B 0.008536f
C305 VTAIL.n274 B 0.008062f
C306 VTAIL.n275 B 0.015002f
C307 VTAIL.n276 B 0.015002f
C308 VTAIL.n277 B 0.008062f
C309 VTAIL.n278 B 0.008536f
C310 VTAIL.n279 B 0.019055f
C311 VTAIL.n280 B 0.019055f
C312 VTAIL.n281 B 0.008536f
C313 VTAIL.n282 B 0.008062f
C314 VTAIL.n283 B 0.015002f
C315 VTAIL.n284 B 0.015002f
C316 VTAIL.n285 B 0.008062f
C317 VTAIL.n286 B 0.008536f
C318 VTAIL.n287 B 0.019055f
C319 VTAIL.n288 B 0.019055f
C320 VTAIL.n289 B 0.008536f
C321 VTAIL.n290 B 0.008062f
C322 VTAIL.n291 B 0.015002f
C323 VTAIL.n292 B 0.015002f
C324 VTAIL.n293 B 0.008062f
C325 VTAIL.n294 B 0.008536f
C326 VTAIL.n295 B 0.019055f
C327 VTAIL.n296 B 0.019055f
C328 VTAIL.n297 B 0.008536f
C329 VTAIL.n298 B 0.008062f
C330 VTAIL.n299 B 0.015002f
C331 VTAIL.n300 B 0.015002f
C332 VTAIL.n301 B 0.008062f
C333 VTAIL.n302 B 0.008536f
C334 VTAIL.n303 B 0.019055f
C335 VTAIL.n304 B 0.019055f
C336 VTAIL.n305 B 0.008536f
C337 VTAIL.n306 B 0.008062f
C338 VTAIL.n307 B 0.015002f
C339 VTAIL.n308 B 0.015002f
C340 VTAIL.n309 B 0.008062f
C341 VTAIL.n310 B 0.008536f
C342 VTAIL.n311 B 0.019055f
C343 VTAIL.n312 B 0.03954f
C344 VTAIL.n313 B 0.008536f
C345 VTAIL.n314 B 0.015763f
C346 VTAIL.n315 B 0.038981f
C347 VTAIL.n316 B 0.041567f
C348 VTAIL.n317 B 1.2196f
C349 VTAIL.n318 B 0.021059f
C350 VTAIL.n319 B 0.015002f
C351 VTAIL.n320 B 0.008062f
C352 VTAIL.n321 B 0.019055f
C353 VTAIL.n322 B 0.008536f
C354 VTAIL.n323 B 0.015002f
C355 VTAIL.n324 B 0.008062f
C356 VTAIL.n325 B 0.019055f
C357 VTAIL.n326 B 0.008536f
C358 VTAIL.n327 B 0.015002f
C359 VTAIL.n328 B 0.008062f
C360 VTAIL.n329 B 0.019055f
C361 VTAIL.n330 B 0.008536f
C362 VTAIL.n331 B 0.015002f
C363 VTAIL.n332 B 0.008062f
C364 VTAIL.n333 B 0.019055f
C365 VTAIL.n334 B 0.008536f
C366 VTAIL.n335 B 0.015002f
C367 VTAIL.n336 B 0.008062f
C368 VTAIL.n337 B 0.019055f
C369 VTAIL.n338 B 0.008536f
C370 VTAIL.n339 B 0.015002f
C371 VTAIL.n340 B 0.008062f
C372 VTAIL.n341 B 0.019055f
C373 VTAIL.n342 B 0.008536f
C374 VTAIL.n343 B 0.015002f
C375 VTAIL.n344 B 0.008062f
C376 VTAIL.n345 B 0.019055f
C377 VTAIL.n346 B 0.019055f
C378 VTAIL.n347 B 0.008536f
C379 VTAIL.n348 B 0.015002f
C380 VTAIL.n349 B 0.008062f
C381 VTAIL.n350 B 0.019055f
C382 VTAIL.n351 B 0.008536f
C383 VTAIL.n352 B 0.151534f
C384 VTAIL.t3 B 0.03279f
C385 VTAIL.n353 B 0.014291f
C386 VTAIL.n354 B 0.01347f
C387 VTAIL.n355 B 0.008062f
C388 VTAIL.n356 B 1.2593f
C389 VTAIL.n357 B 0.015002f
C390 VTAIL.n358 B 0.008062f
C391 VTAIL.n359 B 0.008536f
C392 VTAIL.n360 B 0.019055f
C393 VTAIL.n361 B 0.019055f
C394 VTAIL.n362 B 0.008536f
C395 VTAIL.n363 B 0.008062f
C396 VTAIL.n364 B 0.015002f
C397 VTAIL.n365 B 0.015002f
C398 VTAIL.n366 B 0.008062f
C399 VTAIL.n367 B 0.008536f
C400 VTAIL.n368 B 0.019055f
C401 VTAIL.n369 B 0.019055f
C402 VTAIL.n370 B 0.008536f
C403 VTAIL.n371 B 0.008062f
C404 VTAIL.n372 B 0.015002f
C405 VTAIL.n373 B 0.015002f
C406 VTAIL.n374 B 0.008062f
C407 VTAIL.n375 B 0.008299f
C408 VTAIL.n376 B 0.008299f
C409 VTAIL.n377 B 0.019055f
C410 VTAIL.n378 B 0.019055f
C411 VTAIL.n379 B 0.008536f
C412 VTAIL.n380 B 0.008062f
C413 VTAIL.n381 B 0.015002f
C414 VTAIL.n382 B 0.015002f
C415 VTAIL.n383 B 0.008062f
C416 VTAIL.n384 B 0.008536f
C417 VTAIL.n385 B 0.019055f
C418 VTAIL.n386 B 0.019055f
C419 VTAIL.n387 B 0.008536f
C420 VTAIL.n388 B 0.008062f
C421 VTAIL.n389 B 0.015002f
C422 VTAIL.n390 B 0.015002f
C423 VTAIL.n391 B 0.008062f
C424 VTAIL.n392 B 0.008536f
C425 VTAIL.n393 B 0.019055f
C426 VTAIL.n394 B 0.019055f
C427 VTAIL.n395 B 0.008536f
C428 VTAIL.n396 B 0.008062f
C429 VTAIL.n397 B 0.015002f
C430 VTAIL.n398 B 0.015002f
C431 VTAIL.n399 B 0.008062f
C432 VTAIL.n400 B 0.008536f
C433 VTAIL.n401 B 0.019055f
C434 VTAIL.n402 B 0.019055f
C435 VTAIL.n403 B 0.008536f
C436 VTAIL.n404 B 0.008062f
C437 VTAIL.n405 B 0.015002f
C438 VTAIL.n406 B 0.015002f
C439 VTAIL.n407 B 0.008062f
C440 VTAIL.n408 B 0.008536f
C441 VTAIL.n409 B 0.019055f
C442 VTAIL.n410 B 0.019055f
C443 VTAIL.n411 B 0.008536f
C444 VTAIL.n412 B 0.008062f
C445 VTAIL.n413 B 0.015002f
C446 VTAIL.n414 B 0.015002f
C447 VTAIL.n415 B 0.008062f
C448 VTAIL.n416 B 0.008536f
C449 VTAIL.n417 B 0.019055f
C450 VTAIL.n418 B 0.03954f
C451 VTAIL.n419 B 0.008536f
C452 VTAIL.n420 B 0.015763f
C453 VTAIL.n421 B 0.038981f
C454 VTAIL.n422 B 0.041567f
C455 VTAIL.n423 B 1.2196f
C456 VTAIL.n424 B 0.021059f
C457 VTAIL.n425 B 0.015002f
C458 VTAIL.n426 B 0.008062f
C459 VTAIL.n427 B 0.019055f
C460 VTAIL.n428 B 0.008536f
C461 VTAIL.n429 B 0.015002f
C462 VTAIL.n430 B 0.008062f
C463 VTAIL.n431 B 0.019055f
C464 VTAIL.n432 B 0.008536f
C465 VTAIL.n433 B 0.015002f
C466 VTAIL.n434 B 0.008062f
C467 VTAIL.n435 B 0.019055f
C468 VTAIL.n436 B 0.008536f
C469 VTAIL.n437 B 0.015002f
C470 VTAIL.n438 B 0.008062f
C471 VTAIL.n439 B 0.019055f
C472 VTAIL.n440 B 0.008536f
C473 VTAIL.n441 B 0.015002f
C474 VTAIL.n442 B 0.008062f
C475 VTAIL.n443 B 0.019055f
C476 VTAIL.n444 B 0.008536f
C477 VTAIL.n445 B 0.015002f
C478 VTAIL.n446 B 0.008062f
C479 VTAIL.n447 B 0.019055f
C480 VTAIL.n448 B 0.008536f
C481 VTAIL.n449 B 0.015002f
C482 VTAIL.n450 B 0.008062f
C483 VTAIL.n451 B 0.019055f
C484 VTAIL.n452 B 0.019055f
C485 VTAIL.n453 B 0.008536f
C486 VTAIL.n454 B 0.015002f
C487 VTAIL.n455 B 0.008062f
C488 VTAIL.n456 B 0.019055f
C489 VTAIL.n457 B 0.008536f
C490 VTAIL.n458 B 0.151534f
C491 VTAIL.t1 B 0.03279f
C492 VTAIL.n459 B 0.014291f
C493 VTAIL.n460 B 0.01347f
C494 VTAIL.n461 B 0.008062f
C495 VTAIL.n462 B 1.2593f
C496 VTAIL.n463 B 0.015002f
C497 VTAIL.n464 B 0.008062f
C498 VTAIL.n465 B 0.008536f
C499 VTAIL.n466 B 0.019055f
C500 VTAIL.n467 B 0.019055f
C501 VTAIL.n468 B 0.008536f
C502 VTAIL.n469 B 0.008062f
C503 VTAIL.n470 B 0.015002f
C504 VTAIL.n471 B 0.015002f
C505 VTAIL.n472 B 0.008062f
C506 VTAIL.n473 B 0.008536f
C507 VTAIL.n474 B 0.019055f
C508 VTAIL.n475 B 0.019055f
C509 VTAIL.n476 B 0.008536f
C510 VTAIL.n477 B 0.008062f
C511 VTAIL.n478 B 0.015002f
C512 VTAIL.n479 B 0.015002f
C513 VTAIL.n480 B 0.008062f
C514 VTAIL.n481 B 0.008299f
C515 VTAIL.n482 B 0.008299f
C516 VTAIL.n483 B 0.019055f
C517 VTAIL.n484 B 0.019055f
C518 VTAIL.n485 B 0.008536f
C519 VTAIL.n486 B 0.008062f
C520 VTAIL.n487 B 0.015002f
C521 VTAIL.n488 B 0.015002f
C522 VTAIL.n489 B 0.008062f
C523 VTAIL.n490 B 0.008536f
C524 VTAIL.n491 B 0.019055f
C525 VTAIL.n492 B 0.019055f
C526 VTAIL.n493 B 0.008536f
C527 VTAIL.n494 B 0.008062f
C528 VTAIL.n495 B 0.015002f
C529 VTAIL.n496 B 0.015002f
C530 VTAIL.n497 B 0.008062f
C531 VTAIL.n498 B 0.008536f
C532 VTAIL.n499 B 0.019055f
C533 VTAIL.n500 B 0.019055f
C534 VTAIL.n501 B 0.008536f
C535 VTAIL.n502 B 0.008062f
C536 VTAIL.n503 B 0.015002f
C537 VTAIL.n504 B 0.015002f
C538 VTAIL.n505 B 0.008062f
C539 VTAIL.n506 B 0.008536f
C540 VTAIL.n507 B 0.019055f
C541 VTAIL.n508 B 0.019055f
C542 VTAIL.n509 B 0.008536f
C543 VTAIL.n510 B 0.008062f
C544 VTAIL.n511 B 0.015002f
C545 VTAIL.n512 B 0.015002f
C546 VTAIL.n513 B 0.008062f
C547 VTAIL.n514 B 0.008536f
C548 VTAIL.n515 B 0.019055f
C549 VTAIL.n516 B 0.019055f
C550 VTAIL.n517 B 0.008536f
C551 VTAIL.n518 B 0.008062f
C552 VTAIL.n519 B 0.015002f
C553 VTAIL.n520 B 0.015002f
C554 VTAIL.n521 B 0.008062f
C555 VTAIL.n522 B 0.008536f
C556 VTAIL.n523 B 0.019055f
C557 VTAIL.n524 B 0.03954f
C558 VTAIL.n525 B 0.008536f
C559 VTAIL.n526 B 0.015763f
C560 VTAIL.n527 B 0.038981f
C561 VTAIL.n528 B 0.041567f
C562 VTAIL.n529 B 0.131308f
C563 VTAIL.n530 B 0.021059f
C564 VTAIL.n531 B 0.015002f
C565 VTAIL.n532 B 0.008062f
C566 VTAIL.n533 B 0.019055f
C567 VTAIL.n534 B 0.008536f
C568 VTAIL.n535 B 0.015002f
C569 VTAIL.n536 B 0.008062f
C570 VTAIL.n537 B 0.019055f
C571 VTAIL.n538 B 0.008536f
C572 VTAIL.n539 B 0.015002f
C573 VTAIL.n540 B 0.008062f
C574 VTAIL.n541 B 0.019055f
C575 VTAIL.n542 B 0.008536f
C576 VTAIL.n543 B 0.015002f
C577 VTAIL.n544 B 0.008062f
C578 VTAIL.n545 B 0.019055f
C579 VTAIL.n546 B 0.008536f
C580 VTAIL.n547 B 0.015002f
C581 VTAIL.n548 B 0.008062f
C582 VTAIL.n549 B 0.019055f
C583 VTAIL.n550 B 0.008536f
C584 VTAIL.n551 B 0.015002f
C585 VTAIL.n552 B 0.008062f
C586 VTAIL.n553 B 0.019055f
C587 VTAIL.n554 B 0.008536f
C588 VTAIL.n555 B 0.015002f
C589 VTAIL.n556 B 0.008062f
C590 VTAIL.n557 B 0.019055f
C591 VTAIL.n558 B 0.019055f
C592 VTAIL.n559 B 0.008536f
C593 VTAIL.n560 B 0.015002f
C594 VTAIL.n561 B 0.008062f
C595 VTAIL.n562 B 0.019055f
C596 VTAIL.n563 B 0.008536f
C597 VTAIL.n564 B 0.151534f
C598 VTAIL.t7 B 0.03279f
C599 VTAIL.n565 B 0.014291f
C600 VTAIL.n566 B 0.01347f
C601 VTAIL.n567 B 0.008062f
C602 VTAIL.n568 B 1.2593f
C603 VTAIL.n569 B 0.015002f
C604 VTAIL.n570 B 0.008062f
C605 VTAIL.n571 B 0.008536f
C606 VTAIL.n572 B 0.019055f
C607 VTAIL.n573 B 0.019055f
C608 VTAIL.n574 B 0.008536f
C609 VTAIL.n575 B 0.008062f
C610 VTAIL.n576 B 0.015002f
C611 VTAIL.n577 B 0.015002f
C612 VTAIL.n578 B 0.008062f
C613 VTAIL.n579 B 0.008536f
C614 VTAIL.n580 B 0.019055f
C615 VTAIL.n581 B 0.019055f
C616 VTAIL.n582 B 0.008536f
C617 VTAIL.n583 B 0.008062f
C618 VTAIL.n584 B 0.015002f
C619 VTAIL.n585 B 0.015002f
C620 VTAIL.n586 B 0.008062f
C621 VTAIL.n587 B 0.008299f
C622 VTAIL.n588 B 0.008299f
C623 VTAIL.n589 B 0.019055f
C624 VTAIL.n590 B 0.019055f
C625 VTAIL.n591 B 0.008536f
C626 VTAIL.n592 B 0.008062f
C627 VTAIL.n593 B 0.015002f
C628 VTAIL.n594 B 0.015002f
C629 VTAIL.n595 B 0.008062f
C630 VTAIL.n596 B 0.008536f
C631 VTAIL.n597 B 0.019055f
C632 VTAIL.n598 B 0.019055f
C633 VTAIL.n599 B 0.008536f
C634 VTAIL.n600 B 0.008062f
C635 VTAIL.n601 B 0.015002f
C636 VTAIL.n602 B 0.015002f
C637 VTAIL.n603 B 0.008062f
C638 VTAIL.n604 B 0.008536f
C639 VTAIL.n605 B 0.019055f
C640 VTAIL.n606 B 0.019055f
C641 VTAIL.n607 B 0.008536f
C642 VTAIL.n608 B 0.008062f
C643 VTAIL.n609 B 0.015002f
C644 VTAIL.n610 B 0.015002f
C645 VTAIL.n611 B 0.008062f
C646 VTAIL.n612 B 0.008536f
C647 VTAIL.n613 B 0.019055f
C648 VTAIL.n614 B 0.019055f
C649 VTAIL.n615 B 0.008536f
C650 VTAIL.n616 B 0.008062f
C651 VTAIL.n617 B 0.015002f
C652 VTAIL.n618 B 0.015002f
C653 VTAIL.n619 B 0.008062f
C654 VTAIL.n620 B 0.008536f
C655 VTAIL.n621 B 0.019055f
C656 VTAIL.n622 B 0.019055f
C657 VTAIL.n623 B 0.008536f
C658 VTAIL.n624 B 0.008062f
C659 VTAIL.n625 B 0.015002f
C660 VTAIL.n626 B 0.015002f
C661 VTAIL.n627 B 0.008062f
C662 VTAIL.n628 B 0.008536f
C663 VTAIL.n629 B 0.019055f
C664 VTAIL.n630 B 0.03954f
C665 VTAIL.n631 B 0.008536f
C666 VTAIL.n632 B 0.015763f
C667 VTAIL.n633 B 0.038981f
C668 VTAIL.n634 B 0.041567f
C669 VTAIL.n635 B 0.131308f
C670 VTAIL.n636 B 0.021059f
C671 VTAIL.n637 B 0.015002f
C672 VTAIL.n638 B 0.008062f
C673 VTAIL.n639 B 0.019055f
C674 VTAIL.n640 B 0.008536f
C675 VTAIL.n641 B 0.015002f
C676 VTAIL.n642 B 0.008062f
C677 VTAIL.n643 B 0.019055f
C678 VTAIL.n644 B 0.008536f
C679 VTAIL.n645 B 0.015002f
C680 VTAIL.n646 B 0.008062f
C681 VTAIL.n647 B 0.019055f
C682 VTAIL.n648 B 0.008536f
C683 VTAIL.n649 B 0.015002f
C684 VTAIL.n650 B 0.008062f
C685 VTAIL.n651 B 0.019055f
C686 VTAIL.n652 B 0.008536f
C687 VTAIL.n653 B 0.015002f
C688 VTAIL.n654 B 0.008062f
C689 VTAIL.n655 B 0.019055f
C690 VTAIL.n656 B 0.008536f
C691 VTAIL.n657 B 0.015002f
C692 VTAIL.n658 B 0.008062f
C693 VTAIL.n659 B 0.019055f
C694 VTAIL.n660 B 0.008536f
C695 VTAIL.n661 B 0.015002f
C696 VTAIL.n662 B 0.008062f
C697 VTAIL.n663 B 0.019055f
C698 VTAIL.n664 B 0.019055f
C699 VTAIL.n665 B 0.008536f
C700 VTAIL.n666 B 0.015002f
C701 VTAIL.n667 B 0.008062f
C702 VTAIL.n668 B 0.019055f
C703 VTAIL.n669 B 0.008536f
C704 VTAIL.n670 B 0.151534f
C705 VTAIL.t6 B 0.03279f
C706 VTAIL.n671 B 0.014291f
C707 VTAIL.n672 B 0.01347f
C708 VTAIL.n673 B 0.008062f
C709 VTAIL.n674 B 1.2593f
C710 VTAIL.n675 B 0.015002f
C711 VTAIL.n676 B 0.008062f
C712 VTAIL.n677 B 0.008536f
C713 VTAIL.n678 B 0.019055f
C714 VTAIL.n679 B 0.019055f
C715 VTAIL.n680 B 0.008536f
C716 VTAIL.n681 B 0.008062f
C717 VTAIL.n682 B 0.015002f
C718 VTAIL.n683 B 0.015002f
C719 VTAIL.n684 B 0.008062f
C720 VTAIL.n685 B 0.008536f
C721 VTAIL.n686 B 0.019055f
C722 VTAIL.n687 B 0.019055f
C723 VTAIL.n688 B 0.008536f
C724 VTAIL.n689 B 0.008062f
C725 VTAIL.n690 B 0.015002f
C726 VTAIL.n691 B 0.015002f
C727 VTAIL.n692 B 0.008062f
C728 VTAIL.n693 B 0.008299f
C729 VTAIL.n694 B 0.008299f
C730 VTAIL.n695 B 0.019055f
C731 VTAIL.n696 B 0.019055f
C732 VTAIL.n697 B 0.008536f
C733 VTAIL.n698 B 0.008062f
C734 VTAIL.n699 B 0.015002f
C735 VTAIL.n700 B 0.015002f
C736 VTAIL.n701 B 0.008062f
C737 VTAIL.n702 B 0.008536f
C738 VTAIL.n703 B 0.019055f
C739 VTAIL.n704 B 0.019055f
C740 VTAIL.n705 B 0.008536f
C741 VTAIL.n706 B 0.008062f
C742 VTAIL.n707 B 0.015002f
C743 VTAIL.n708 B 0.015002f
C744 VTAIL.n709 B 0.008062f
C745 VTAIL.n710 B 0.008536f
C746 VTAIL.n711 B 0.019055f
C747 VTAIL.n712 B 0.019055f
C748 VTAIL.n713 B 0.008536f
C749 VTAIL.n714 B 0.008062f
C750 VTAIL.n715 B 0.015002f
C751 VTAIL.n716 B 0.015002f
C752 VTAIL.n717 B 0.008062f
C753 VTAIL.n718 B 0.008536f
C754 VTAIL.n719 B 0.019055f
C755 VTAIL.n720 B 0.019055f
C756 VTAIL.n721 B 0.008536f
C757 VTAIL.n722 B 0.008062f
C758 VTAIL.n723 B 0.015002f
C759 VTAIL.n724 B 0.015002f
C760 VTAIL.n725 B 0.008062f
C761 VTAIL.n726 B 0.008536f
C762 VTAIL.n727 B 0.019055f
C763 VTAIL.n728 B 0.019055f
C764 VTAIL.n729 B 0.008536f
C765 VTAIL.n730 B 0.008062f
C766 VTAIL.n731 B 0.015002f
C767 VTAIL.n732 B 0.015002f
C768 VTAIL.n733 B 0.008062f
C769 VTAIL.n734 B 0.008536f
C770 VTAIL.n735 B 0.019055f
C771 VTAIL.n736 B 0.03954f
C772 VTAIL.n737 B 0.008536f
C773 VTAIL.n738 B 0.015763f
C774 VTAIL.n739 B 0.038981f
C775 VTAIL.n740 B 0.041567f
C776 VTAIL.n741 B 1.2196f
C777 VTAIL.n742 B 0.021059f
C778 VTAIL.n743 B 0.015002f
C779 VTAIL.n744 B 0.008062f
C780 VTAIL.n745 B 0.019055f
C781 VTAIL.n746 B 0.008536f
C782 VTAIL.n747 B 0.015002f
C783 VTAIL.n748 B 0.008062f
C784 VTAIL.n749 B 0.019055f
C785 VTAIL.n750 B 0.008536f
C786 VTAIL.n751 B 0.015002f
C787 VTAIL.n752 B 0.008062f
C788 VTAIL.n753 B 0.019055f
C789 VTAIL.n754 B 0.008536f
C790 VTAIL.n755 B 0.015002f
C791 VTAIL.n756 B 0.008062f
C792 VTAIL.n757 B 0.019055f
C793 VTAIL.n758 B 0.008536f
C794 VTAIL.n759 B 0.015002f
C795 VTAIL.n760 B 0.008062f
C796 VTAIL.n761 B 0.019055f
C797 VTAIL.n762 B 0.008536f
C798 VTAIL.n763 B 0.015002f
C799 VTAIL.n764 B 0.008062f
C800 VTAIL.n765 B 0.019055f
C801 VTAIL.n766 B 0.008536f
C802 VTAIL.n767 B 0.015002f
C803 VTAIL.n768 B 0.008062f
C804 VTAIL.n769 B 0.019055f
C805 VTAIL.n770 B 0.008536f
C806 VTAIL.n771 B 0.015002f
C807 VTAIL.n772 B 0.008062f
C808 VTAIL.n773 B 0.019055f
C809 VTAIL.n774 B 0.008536f
C810 VTAIL.n775 B 0.151534f
C811 VTAIL.t0 B 0.03279f
C812 VTAIL.n776 B 0.014291f
C813 VTAIL.n777 B 0.01347f
C814 VTAIL.n778 B 0.008062f
C815 VTAIL.n779 B 1.2593f
C816 VTAIL.n780 B 0.015002f
C817 VTAIL.n781 B 0.008062f
C818 VTAIL.n782 B 0.008536f
C819 VTAIL.n783 B 0.019055f
C820 VTAIL.n784 B 0.019055f
C821 VTAIL.n785 B 0.008536f
C822 VTAIL.n786 B 0.008062f
C823 VTAIL.n787 B 0.015002f
C824 VTAIL.n788 B 0.015002f
C825 VTAIL.n789 B 0.008062f
C826 VTAIL.n790 B 0.008536f
C827 VTAIL.n791 B 0.019055f
C828 VTAIL.n792 B 0.019055f
C829 VTAIL.n793 B 0.019055f
C830 VTAIL.n794 B 0.008536f
C831 VTAIL.n795 B 0.008062f
C832 VTAIL.n796 B 0.015002f
C833 VTAIL.n797 B 0.015002f
C834 VTAIL.n798 B 0.008062f
C835 VTAIL.n799 B 0.008299f
C836 VTAIL.n800 B 0.008299f
C837 VTAIL.n801 B 0.019055f
C838 VTAIL.n802 B 0.019055f
C839 VTAIL.n803 B 0.008536f
C840 VTAIL.n804 B 0.008062f
C841 VTAIL.n805 B 0.015002f
C842 VTAIL.n806 B 0.015002f
C843 VTAIL.n807 B 0.008062f
C844 VTAIL.n808 B 0.008536f
C845 VTAIL.n809 B 0.019055f
C846 VTAIL.n810 B 0.019055f
C847 VTAIL.n811 B 0.008536f
C848 VTAIL.n812 B 0.008062f
C849 VTAIL.n813 B 0.015002f
C850 VTAIL.n814 B 0.015002f
C851 VTAIL.n815 B 0.008062f
C852 VTAIL.n816 B 0.008536f
C853 VTAIL.n817 B 0.019055f
C854 VTAIL.n818 B 0.019055f
C855 VTAIL.n819 B 0.008536f
C856 VTAIL.n820 B 0.008062f
C857 VTAIL.n821 B 0.015002f
C858 VTAIL.n822 B 0.015002f
C859 VTAIL.n823 B 0.008062f
C860 VTAIL.n824 B 0.008536f
C861 VTAIL.n825 B 0.019055f
C862 VTAIL.n826 B 0.019055f
C863 VTAIL.n827 B 0.008536f
C864 VTAIL.n828 B 0.008062f
C865 VTAIL.n829 B 0.015002f
C866 VTAIL.n830 B 0.015002f
C867 VTAIL.n831 B 0.008062f
C868 VTAIL.n832 B 0.008536f
C869 VTAIL.n833 B 0.019055f
C870 VTAIL.n834 B 0.019055f
C871 VTAIL.n835 B 0.008536f
C872 VTAIL.n836 B 0.008062f
C873 VTAIL.n837 B 0.015002f
C874 VTAIL.n838 B 0.015002f
C875 VTAIL.n839 B 0.008062f
C876 VTAIL.n840 B 0.008536f
C877 VTAIL.n841 B 0.019055f
C878 VTAIL.n842 B 0.03954f
C879 VTAIL.n843 B 0.008536f
C880 VTAIL.n844 B 0.015763f
C881 VTAIL.n845 B 0.038981f
C882 VTAIL.n846 B 0.041567f
C883 VTAIL.n847 B 1.17011f
C884 VDD1.t2 B 0.409892f
C885 VDD1.t0 B 0.409892f
C886 VDD1.n0 B 3.75621f
C887 VDD1.t3 B 0.409892f
C888 VDD1.t1 B 0.409892f
C889 VDD1.n1 B 4.66697f
C890 VP.n0 B 0.039409f
C891 VP.t2 B 3.0715f
C892 VP.n1 B 0.043637f
C893 VP.t1 B 3.22104f
C894 VP.t0 B 3.22331f
C895 VP.n2 B 3.80464f
C896 VP.n3 B 1.90978f
C897 VP.t3 B 3.0715f
C898 VP.n4 B 1.15377f
C899 VP.n5 B 0.04856f
C900 VP.n6 B 0.039409f
C901 VP.n7 B 0.029892f
C902 VP.n8 B 0.029892f
C903 VP.n9 B 0.043637f
C904 VP.n10 B 0.04856f
C905 VP.n11 B 1.15377f
C906 VP.n12 B 0.037176f
.ends

