* NGSPICE file created from diff_pair_sample_0098.ext - technology: sky130A

.subckt diff_pair_sample_0098 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t16 B.t1 sky130_fd_pr__nfet_01v8 ad=2.94525 pd=18.18 as=2.94525 ps=18.18 w=17.85 l=2.46
X1 VTAIL.t5 VN.t0 VDD2.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=2.94525 pd=18.18 as=2.94525 ps=18.18 w=17.85 l=2.46
X2 VDD2.t8 VN.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.94525 pd=18.18 as=6.9615 ps=36.48 w=17.85 l=2.46
X3 VDD1.t8 VP.t1 VTAIL.t19 B.t9 sky130_fd_pr__nfet_01v8 ad=2.94525 pd=18.18 as=6.9615 ps=36.48 w=17.85 l=2.46
X4 VTAIL.t18 VP.t2 VDD1.t7 B.t4 sky130_fd_pr__nfet_01v8 ad=2.94525 pd=18.18 as=2.94525 ps=18.18 w=17.85 l=2.46
X5 VTAIL.t15 VP.t3 VDD1.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=2.94525 pd=18.18 as=2.94525 ps=18.18 w=17.85 l=2.46
X6 VDD2.t7 VN.t2 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=2.94525 pd=18.18 as=2.94525 ps=18.18 w=17.85 l=2.46
X7 VTAIL.t4 VN.t3 VDD2.t6 B.t4 sky130_fd_pr__nfet_01v8 ad=2.94525 pd=18.18 as=2.94525 ps=18.18 w=17.85 l=2.46
X8 VDD1.t5 VP.t4 VTAIL.t11 B.t0 sky130_fd_pr__nfet_01v8 ad=2.94525 pd=18.18 as=6.9615 ps=36.48 w=17.85 l=2.46
X9 B.t23 B.t21 B.t22 B.t15 sky130_fd_pr__nfet_01v8 ad=6.9615 pd=36.48 as=0 ps=0 w=17.85 l=2.46
X10 VTAIL.t3 VN.t4 VDD2.t5 B.t3 sky130_fd_pr__nfet_01v8 ad=2.94525 pd=18.18 as=2.94525 ps=18.18 w=17.85 l=2.46
X11 B.t20 B.t18 B.t19 B.t11 sky130_fd_pr__nfet_01v8 ad=6.9615 pd=36.48 as=0 ps=0 w=17.85 l=2.46
X12 VDD2.t4 VN.t5 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=6.9615 pd=36.48 as=2.94525 ps=18.18 w=17.85 l=2.46
X13 VTAIL.t2 VN.t6 VDD2.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=2.94525 pd=18.18 as=2.94525 ps=18.18 w=17.85 l=2.46
X14 VDD1.t4 VP.t5 VTAIL.t17 B.t6 sky130_fd_pr__nfet_01v8 ad=6.9615 pd=36.48 as=2.94525 ps=18.18 w=17.85 l=2.46
X15 VDD2.t2 VN.t7 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.94525 pd=18.18 as=2.94525 ps=18.18 w=17.85 l=2.46
X16 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=6.9615 pd=36.48 as=0 ps=0 w=17.85 l=2.46
X17 VDD2.t1 VN.t8 VTAIL.t8 B.t8 sky130_fd_pr__nfet_01v8 ad=6.9615 pd=36.48 as=2.94525 ps=18.18 w=17.85 l=2.46
X18 VDD1.t3 VP.t6 VTAIL.t14 B.t8 sky130_fd_pr__nfet_01v8 ad=6.9615 pd=36.48 as=2.94525 ps=18.18 w=17.85 l=2.46
X19 VDD2.t0 VN.t9 VTAIL.t9 B.t9 sky130_fd_pr__nfet_01v8 ad=2.94525 pd=18.18 as=6.9615 ps=36.48 w=17.85 l=2.46
X20 VTAIL.t10 VP.t7 VDD1.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=2.94525 pd=18.18 as=2.94525 ps=18.18 w=17.85 l=2.46
X21 VDD1.t1 VP.t8 VTAIL.t13 B.t7 sky130_fd_pr__nfet_01v8 ad=2.94525 pd=18.18 as=2.94525 ps=18.18 w=17.85 l=2.46
X22 VTAIL.t12 VP.t9 VDD1.t0 B.t5 sky130_fd_pr__nfet_01v8 ad=2.94525 pd=18.18 as=2.94525 ps=18.18 w=17.85 l=2.46
X23 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=6.9615 pd=36.48 as=0 ps=0 w=17.85 l=2.46
R0 VP.n23 VP.t6 206.546
R1 VP.n71 VP.t8 174.873
R2 VP.n53 VP.t5 174.873
R3 VP.n9 VP.t9 174.873
R4 VP.n3 VP.t3 174.873
R5 VP.n89 VP.t1 174.873
R6 VP.n32 VP.t0 174.873
R7 VP.n50 VP.t4 174.873
R8 VP.n16 VP.t7 174.873
R9 VP.n22 VP.t2 174.873
R10 VP.n25 VP.n24 161.3
R11 VP.n26 VP.n21 161.3
R12 VP.n28 VP.n27 161.3
R13 VP.n29 VP.n20 161.3
R14 VP.n31 VP.n30 161.3
R15 VP.n32 VP.n19 161.3
R16 VP.n34 VP.n33 161.3
R17 VP.n35 VP.n18 161.3
R18 VP.n37 VP.n36 161.3
R19 VP.n38 VP.n17 161.3
R20 VP.n40 VP.n39 161.3
R21 VP.n42 VP.n41 161.3
R22 VP.n43 VP.n15 161.3
R23 VP.n45 VP.n44 161.3
R24 VP.n46 VP.n14 161.3
R25 VP.n48 VP.n47 161.3
R26 VP.n49 VP.n13 161.3
R27 VP.n88 VP.n0 161.3
R28 VP.n87 VP.n86 161.3
R29 VP.n85 VP.n1 161.3
R30 VP.n84 VP.n83 161.3
R31 VP.n82 VP.n2 161.3
R32 VP.n81 VP.n80 161.3
R33 VP.n79 VP.n78 161.3
R34 VP.n77 VP.n4 161.3
R35 VP.n76 VP.n75 161.3
R36 VP.n74 VP.n5 161.3
R37 VP.n73 VP.n72 161.3
R38 VP.n71 VP.n6 161.3
R39 VP.n70 VP.n69 161.3
R40 VP.n68 VP.n7 161.3
R41 VP.n67 VP.n66 161.3
R42 VP.n65 VP.n8 161.3
R43 VP.n64 VP.n63 161.3
R44 VP.n62 VP.n61 161.3
R45 VP.n60 VP.n10 161.3
R46 VP.n59 VP.n58 161.3
R47 VP.n57 VP.n11 161.3
R48 VP.n56 VP.n55 161.3
R49 VP.n54 VP.n12 161.3
R50 VP.n53 VP.n52 106.841
R51 VP.n90 VP.n89 106.841
R52 VP.n51 VP.n50 106.841
R53 VP.n23 VP.n22 57.8794
R54 VP.n52 VP.n51 56.6776
R55 VP.n59 VP.n11 56.5193
R56 VP.n83 VP.n1 56.5193
R57 VP.n44 VP.n14 56.5193
R58 VP.n66 VP.n7 50.6917
R59 VP.n76 VP.n5 50.6917
R60 VP.n37 VP.n18 50.6917
R61 VP.n27 VP.n20 50.6917
R62 VP.n66 VP.n65 30.2951
R63 VP.n77 VP.n76 30.2951
R64 VP.n38 VP.n37 30.2951
R65 VP.n27 VP.n26 30.2951
R66 VP.n55 VP.n54 24.4675
R67 VP.n55 VP.n11 24.4675
R68 VP.n60 VP.n59 24.4675
R69 VP.n61 VP.n60 24.4675
R70 VP.n65 VP.n64 24.4675
R71 VP.n70 VP.n7 24.4675
R72 VP.n71 VP.n70 24.4675
R73 VP.n72 VP.n71 24.4675
R74 VP.n72 VP.n5 24.4675
R75 VP.n78 VP.n77 24.4675
R76 VP.n82 VP.n81 24.4675
R77 VP.n83 VP.n82 24.4675
R78 VP.n87 VP.n1 24.4675
R79 VP.n88 VP.n87 24.4675
R80 VP.n48 VP.n14 24.4675
R81 VP.n49 VP.n48 24.4675
R82 VP.n39 VP.n38 24.4675
R83 VP.n43 VP.n42 24.4675
R84 VP.n44 VP.n43 24.4675
R85 VP.n31 VP.n20 24.4675
R86 VP.n32 VP.n31 24.4675
R87 VP.n33 VP.n32 24.4675
R88 VP.n33 VP.n18 24.4675
R89 VP.n26 VP.n25 24.4675
R90 VP.n64 VP.n9 14.1914
R91 VP.n78 VP.n3 14.1914
R92 VP.n39 VP.n16 14.1914
R93 VP.n25 VP.n22 14.1914
R94 VP.n61 VP.n9 10.2766
R95 VP.n81 VP.n3 10.2766
R96 VP.n42 VP.n16 10.2766
R97 VP.n24 VP.n23 7.2327
R98 VP.n54 VP.n53 3.91522
R99 VP.n89 VP.n88 3.91522
R100 VP.n50 VP.n49 3.91522
R101 VP.n51 VP.n13 0.278367
R102 VP.n52 VP.n12 0.278367
R103 VP.n90 VP.n0 0.278367
R104 VP.n24 VP.n21 0.189894
R105 VP.n28 VP.n21 0.189894
R106 VP.n29 VP.n28 0.189894
R107 VP.n30 VP.n29 0.189894
R108 VP.n30 VP.n19 0.189894
R109 VP.n34 VP.n19 0.189894
R110 VP.n35 VP.n34 0.189894
R111 VP.n36 VP.n35 0.189894
R112 VP.n36 VP.n17 0.189894
R113 VP.n40 VP.n17 0.189894
R114 VP.n41 VP.n40 0.189894
R115 VP.n41 VP.n15 0.189894
R116 VP.n45 VP.n15 0.189894
R117 VP.n46 VP.n45 0.189894
R118 VP.n47 VP.n46 0.189894
R119 VP.n47 VP.n13 0.189894
R120 VP.n56 VP.n12 0.189894
R121 VP.n57 VP.n56 0.189894
R122 VP.n58 VP.n57 0.189894
R123 VP.n58 VP.n10 0.189894
R124 VP.n62 VP.n10 0.189894
R125 VP.n63 VP.n62 0.189894
R126 VP.n63 VP.n8 0.189894
R127 VP.n67 VP.n8 0.189894
R128 VP.n68 VP.n67 0.189894
R129 VP.n69 VP.n68 0.189894
R130 VP.n69 VP.n6 0.189894
R131 VP.n73 VP.n6 0.189894
R132 VP.n74 VP.n73 0.189894
R133 VP.n75 VP.n74 0.189894
R134 VP.n75 VP.n4 0.189894
R135 VP.n79 VP.n4 0.189894
R136 VP.n80 VP.n79 0.189894
R137 VP.n80 VP.n2 0.189894
R138 VP.n84 VP.n2 0.189894
R139 VP.n85 VP.n84 0.189894
R140 VP.n86 VP.n85 0.189894
R141 VP.n86 VP.n0 0.189894
R142 VP VP.n90 0.153454
R143 VTAIL.n11 VTAIL.t9 44.5126
R144 VTAIL.n17 VTAIL.t0 44.5124
R145 VTAIL.n2 VTAIL.t19 44.5124
R146 VTAIL.n16 VTAIL.t11 44.5124
R147 VTAIL.n15 VTAIL.n14 43.4034
R148 VTAIL.n13 VTAIL.n12 43.4034
R149 VTAIL.n10 VTAIL.n9 43.4034
R150 VTAIL.n8 VTAIL.n7 43.4034
R151 VTAIL.n19 VTAIL.n18 43.4032
R152 VTAIL.n1 VTAIL.n0 43.4032
R153 VTAIL.n4 VTAIL.n3 43.4032
R154 VTAIL.n6 VTAIL.n5 43.4032
R155 VTAIL.n8 VTAIL.n6 32.5652
R156 VTAIL.n17 VTAIL.n16 30.16
R157 VTAIL.n10 VTAIL.n8 2.40567
R158 VTAIL.n11 VTAIL.n10 2.40567
R159 VTAIL.n15 VTAIL.n13 2.40567
R160 VTAIL.n16 VTAIL.n15 2.40567
R161 VTAIL.n6 VTAIL.n4 2.40567
R162 VTAIL.n4 VTAIL.n2 2.40567
R163 VTAIL.n19 VTAIL.n17 2.40567
R164 VTAIL VTAIL.n1 1.86257
R165 VTAIL.n13 VTAIL.n11 1.67291
R166 VTAIL.n2 VTAIL.n1 1.67291
R167 VTAIL.n18 VTAIL.t1 1.10974
R168 VTAIL.n18 VTAIL.t3 1.10974
R169 VTAIL.n0 VTAIL.t8 1.10974
R170 VTAIL.n0 VTAIL.t4 1.10974
R171 VTAIL.n3 VTAIL.t13 1.10974
R172 VTAIL.n3 VTAIL.t15 1.10974
R173 VTAIL.n5 VTAIL.t17 1.10974
R174 VTAIL.n5 VTAIL.t12 1.10974
R175 VTAIL.n14 VTAIL.t16 1.10974
R176 VTAIL.n14 VTAIL.t10 1.10974
R177 VTAIL.n12 VTAIL.t14 1.10974
R178 VTAIL.n12 VTAIL.t18 1.10974
R179 VTAIL.n9 VTAIL.t7 1.10974
R180 VTAIL.n9 VTAIL.t2 1.10974
R181 VTAIL.n7 VTAIL.t6 1.10974
R182 VTAIL.n7 VTAIL.t5 1.10974
R183 VTAIL VTAIL.n19 0.543603
R184 VDD1.n1 VDD1.t3 63.5966
R185 VDD1.n3 VDD1.t4 63.5964
R186 VDD1.n5 VDD1.n4 61.8305
R187 VDD1.n1 VDD1.n0 60.0822
R188 VDD1.n7 VDD1.n6 60.082
R189 VDD1.n3 VDD1.n2 60.0819
R190 VDD1.n7 VDD1.n5 52.3134
R191 VDD1 VDD1.n7 1.74619
R192 VDD1.n6 VDD1.t2 1.10974
R193 VDD1.n6 VDD1.t5 1.10974
R194 VDD1.n0 VDD1.t7 1.10974
R195 VDD1.n0 VDD1.t9 1.10974
R196 VDD1.n4 VDD1.t6 1.10974
R197 VDD1.n4 VDD1.t8 1.10974
R198 VDD1.n2 VDD1.t0 1.10974
R199 VDD1.n2 VDD1.t1 1.10974
R200 VDD1 VDD1.n1 0.659983
R201 VDD1.n5 VDD1.n3 0.546447
R202 B.n1108 B.n1107 585
R203 B.n1109 B.n1108 585
R204 B.n426 B.n169 585
R205 B.n425 B.n424 585
R206 B.n423 B.n422 585
R207 B.n421 B.n420 585
R208 B.n419 B.n418 585
R209 B.n417 B.n416 585
R210 B.n415 B.n414 585
R211 B.n413 B.n412 585
R212 B.n411 B.n410 585
R213 B.n409 B.n408 585
R214 B.n407 B.n406 585
R215 B.n405 B.n404 585
R216 B.n403 B.n402 585
R217 B.n401 B.n400 585
R218 B.n399 B.n398 585
R219 B.n397 B.n396 585
R220 B.n395 B.n394 585
R221 B.n393 B.n392 585
R222 B.n391 B.n390 585
R223 B.n389 B.n388 585
R224 B.n387 B.n386 585
R225 B.n385 B.n384 585
R226 B.n383 B.n382 585
R227 B.n381 B.n380 585
R228 B.n379 B.n378 585
R229 B.n377 B.n376 585
R230 B.n375 B.n374 585
R231 B.n373 B.n372 585
R232 B.n371 B.n370 585
R233 B.n369 B.n368 585
R234 B.n367 B.n366 585
R235 B.n365 B.n364 585
R236 B.n363 B.n362 585
R237 B.n361 B.n360 585
R238 B.n359 B.n358 585
R239 B.n357 B.n356 585
R240 B.n355 B.n354 585
R241 B.n353 B.n352 585
R242 B.n351 B.n350 585
R243 B.n349 B.n348 585
R244 B.n347 B.n346 585
R245 B.n345 B.n344 585
R246 B.n343 B.n342 585
R247 B.n341 B.n340 585
R248 B.n339 B.n338 585
R249 B.n337 B.n336 585
R250 B.n335 B.n334 585
R251 B.n333 B.n332 585
R252 B.n331 B.n330 585
R253 B.n329 B.n328 585
R254 B.n327 B.n326 585
R255 B.n325 B.n324 585
R256 B.n323 B.n322 585
R257 B.n321 B.n320 585
R258 B.n319 B.n318 585
R259 B.n317 B.n316 585
R260 B.n315 B.n314 585
R261 B.n313 B.n312 585
R262 B.n311 B.n310 585
R263 B.n309 B.n308 585
R264 B.n307 B.n306 585
R265 B.n305 B.n304 585
R266 B.n303 B.n302 585
R267 B.n301 B.n300 585
R268 B.n299 B.n298 585
R269 B.n297 B.n296 585
R270 B.n295 B.n294 585
R271 B.n292 B.n291 585
R272 B.n290 B.n289 585
R273 B.n288 B.n287 585
R274 B.n286 B.n285 585
R275 B.n284 B.n283 585
R276 B.n282 B.n281 585
R277 B.n280 B.n279 585
R278 B.n278 B.n277 585
R279 B.n276 B.n275 585
R280 B.n274 B.n273 585
R281 B.n272 B.n271 585
R282 B.n270 B.n269 585
R283 B.n268 B.n267 585
R284 B.n266 B.n265 585
R285 B.n264 B.n263 585
R286 B.n262 B.n261 585
R287 B.n260 B.n259 585
R288 B.n258 B.n257 585
R289 B.n256 B.n255 585
R290 B.n254 B.n253 585
R291 B.n252 B.n251 585
R292 B.n250 B.n249 585
R293 B.n248 B.n247 585
R294 B.n246 B.n245 585
R295 B.n244 B.n243 585
R296 B.n242 B.n241 585
R297 B.n240 B.n239 585
R298 B.n238 B.n237 585
R299 B.n236 B.n235 585
R300 B.n234 B.n233 585
R301 B.n232 B.n231 585
R302 B.n230 B.n229 585
R303 B.n228 B.n227 585
R304 B.n226 B.n225 585
R305 B.n224 B.n223 585
R306 B.n222 B.n221 585
R307 B.n220 B.n219 585
R308 B.n218 B.n217 585
R309 B.n216 B.n215 585
R310 B.n214 B.n213 585
R311 B.n212 B.n211 585
R312 B.n210 B.n209 585
R313 B.n208 B.n207 585
R314 B.n206 B.n205 585
R315 B.n204 B.n203 585
R316 B.n202 B.n201 585
R317 B.n200 B.n199 585
R318 B.n198 B.n197 585
R319 B.n196 B.n195 585
R320 B.n194 B.n193 585
R321 B.n192 B.n191 585
R322 B.n190 B.n189 585
R323 B.n188 B.n187 585
R324 B.n186 B.n185 585
R325 B.n184 B.n183 585
R326 B.n182 B.n181 585
R327 B.n180 B.n179 585
R328 B.n178 B.n177 585
R329 B.n176 B.n175 585
R330 B.n1106 B.n105 585
R331 B.n1110 B.n105 585
R332 B.n1105 B.n104 585
R333 B.n1111 B.n104 585
R334 B.n1104 B.n1103 585
R335 B.n1103 B.n100 585
R336 B.n1102 B.n99 585
R337 B.n1117 B.n99 585
R338 B.n1101 B.n98 585
R339 B.n1118 B.n98 585
R340 B.n1100 B.n97 585
R341 B.n1119 B.n97 585
R342 B.n1099 B.n1098 585
R343 B.n1098 B.n93 585
R344 B.n1097 B.n92 585
R345 B.n1125 B.n92 585
R346 B.n1096 B.n91 585
R347 B.n1126 B.n91 585
R348 B.n1095 B.n90 585
R349 B.n1127 B.n90 585
R350 B.n1094 B.n1093 585
R351 B.n1093 B.n86 585
R352 B.n1092 B.n85 585
R353 B.n1133 B.n85 585
R354 B.n1091 B.n84 585
R355 B.n1134 B.n84 585
R356 B.n1090 B.n83 585
R357 B.n1135 B.n83 585
R358 B.n1089 B.n1088 585
R359 B.n1088 B.n79 585
R360 B.n1087 B.n78 585
R361 B.n1141 B.n78 585
R362 B.n1086 B.n77 585
R363 B.n1142 B.n77 585
R364 B.n1085 B.n76 585
R365 B.n1143 B.n76 585
R366 B.n1084 B.n1083 585
R367 B.n1083 B.n75 585
R368 B.n1082 B.n71 585
R369 B.n1149 B.n71 585
R370 B.n1081 B.n70 585
R371 B.n1150 B.n70 585
R372 B.n1080 B.n69 585
R373 B.n1151 B.n69 585
R374 B.n1079 B.n1078 585
R375 B.n1078 B.n65 585
R376 B.n1077 B.n64 585
R377 B.n1157 B.n64 585
R378 B.n1076 B.n63 585
R379 B.n1158 B.n63 585
R380 B.n1075 B.n62 585
R381 B.n1159 B.n62 585
R382 B.n1074 B.n1073 585
R383 B.n1073 B.n58 585
R384 B.n1072 B.n57 585
R385 B.n1165 B.n57 585
R386 B.n1071 B.n56 585
R387 B.n1166 B.n56 585
R388 B.n1070 B.n55 585
R389 B.n1167 B.n55 585
R390 B.n1069 B.n1068 585
R391 B.n1068 B.n51 585
R392 B.n1067 B.n50 585
R393 B.n1173 B.n50 585
R394 B.n1066 B.n49 585
R395 B.n1174 B.n49 585
R396 B.n1065 B.n48 585
R397 B.n1175 B.n48 585
R398 B.n1064 B.n1063 585
R399 B.n1063 B.n44 585
R400 B.n1062 B.n43 585
R401 B.n1181 B.n43 585
R402 B.n1061 B.n42 585
R403 B.n1182 B.n42 585
R404 B.n1060 B.n41 585
R405 B.n1183 B.n41 585
R406 B.n1059 B.n1058 585
R407 B.n1058 B.n37 585
R408 B.n1057 B.n36 585
R409 B.n1189 B.n36 585
R410 B.n1056 B.n35 585
R411 B.n1190 B.n35 585
R412 B.n1055 B.n34 585
R413 B.n1191 B.n34 585
R414 B.n1054 B.n1053 585
R415 B.n1053 B.n30 585
R416 B.n1052 B.n29 585
R417 B.n1197 B.n29 585
R418 B.n1051 B.n28 585
R419 B.n1198 B.n28 585
R420 B.n1050 B.n27 585
R421 B.n1199 B.n27 585
R422 B.n1049 B.n1048 585
R423 B.n1048 B.n23 585
R424 B.n1047 B.n22 585
R425 B.n1205 B.n22 585
R426 B.n1046 B.n21 585
R427 B.n1206 B.n21 585
R428 B.n1045 B.n20 585
R429 B.n1207 B.n20 585
R430 B.n1044 B.n1043 585
R431 B.n1043 B.n16 585
R432 B.n1042 B.n15 585
R433 B.n1213 B.n15 585
R434 B.n1041 B.n14 585
R435 B.n1214 B.n14 585
R436 B.n1040 B.n13 585
R437 B.n1215 B.n13 585
R438 B.n1039 B.n1038 585
R439 B.n1038 B.n12 585
R440 B.n1037 B.n1036 585
R441 B.n1037 B.n8 585
R442 B.n1035 B.n7 585
R443 B.n1222 B.n7 585
R444 B.n1034 B.n6 585
R445 B.n1223 B.n6 585
R446 B.n1033 B.n5 585
R447 B.n1224 B.n5 585
R448 B.n1032 B.n1031 585
R449 B.n1031 B.n4 585
R450 B.n1030 B.n427 585
R451 B.n1030 B.n1029 585
R452 B.n1020 B.n428 585
R453 B.n429 B.n428 585
R454 B.n1022 B.n1021 585
R455 B.n1023 B.n1022 585
R456 B.n1019 B.n434 585
R457 B.n434 B.n433 585
R458 B.n1018 B.n1017 585
R459 B.n1017 B.n1016 585
R460 B.n436 B.n435 585
R461 B.n437 B.n436 585
R462 B.n1009 B.n1008 585
R463 B.n1010 B.n1009 585
R464 B.n1007 B.n442 585
R465 B.n442 B.n441 585
R466 B.n1006 B.n1005 585
R467 B.n1005 B.n1004 585
R468 B.n444 B.n443 585
R469 B.n445 B.n444 585
R470 B.n997 B.n996 585
R471 B.n998 B.n997 585
R472 B.n995 B.n450 585
R473 B.n450 B.n449 585
R474 B.n994 B.n993 585
R475 B.n993 B.n992 585
R476 B.n452 B.n451 585
R477 B.n453 B.n452 585
R478 B.n985 B.n984 585
R479 B.n986 B.n985 585
R480 B.n983 B.n458 585
R481 B.n458 B.n457 585
R482 B.n982 B.n981 585
R483 B.n981 B.n980 585
R484 B.n460 B.n459 585
R485 B.n461 B.n460 585
R486 B.n973 B.n972 585
R487 B.n974 B.n973 585
R488 B.n971 B.n466 585
R489 B.n466 B.n465 585
R490 B.n970 B.n969 585
R491 B.n969 B.n968 585
R492 B.n468 B.n467 585
R493 B.n469 B.n468 585
R494 B.n961 B.n960 585
R495 B.n962 B.n961 585
R496 B.n959 B.n474 585
R497 B.n474 B.n473 585
R498 B.n958 B.n957 585
R499 B.n957 B.n956 585
R500 B.n476 B.n475 585
R501 B.n477 B.n476 585
R502 B.n949 B.n948 585
R503 B.n950 B.n949 585
R504 B.n947 B.n482 585
R505 B.n482 B.n481 585
R506 B.n946 B.n945 585
R507 B.n945 B.n944 585
R508 B.n484 B.n483 585
R509 B.n485 B.n484 585
R510 B.n937 B.n936 585
R511 B.n938 B.n937 585
R512 B.n935 B.n490 585
R513 B.n490 B.n489 585
R514 B.n934 B.n933 585
R515 B.n933 B.n932 585
R516 B.n492 B.n491 585
R517 B.n493 B.n492 585
R518 B.n925 B.n924 585
R519 B.n926 B.n925 585
R520 B.n923 B.n498 585
R521 B.n498 B.n497 585
R522 B.n922 B.n921 585
R523 B.n921 B.n920 585
R524 B.n500 B.n499 585
R525 B.n913 B.n500 585
R526 B.n912 B.n911 585
R527 B.n914 B.n912 585
R528 B.n910 B.n505 585
R529 B.n505 B.n504 585
R530 B.n909 B.n908 585
R531 B.n908 B.n907 585
R532 B.n507 B.n506 585
R533 B.n508 B.n507 585
R534 B.n900 B.n899 585
R535 B.n901 B.n900 585
R536 B.n898 B.n513 585
R537 B.n513 B.n512 585
R538 B.n897 B.n896 585
R539 B.n896 B.n895 585
R540 B.n515 B.n514 585
R541 B.n516 B.n515 585
R542 B.n888 B.n887 585
R543 B.n889 B.n888 585
R544 B.n886 B.n521 585
R545 B.n521 B.n520 585
R546 B.n885 B.n884 585
R547 B.n884 B.n883 585
R548 B.n523 B.n522 585
R549 B.n524 B.n523 585
R550 B.n876 B.n875 585
R551 B.n877 B.n876 585
R552 B.n874 B.n529 585
R553 B.n529 B.n528 585
R554 B.n873 B.n872 585
R555 B.n872 B.n871 585
R556 B.n531 B.n530 585
R557 B.n532 B.n531 585
R558 B.n864 B.n863 585
R559 B.n865 B.n864 585
R560 B.n862 B.n537 585
R561 B.n537 B.n536 585
R562 B.n856 B.n855 585
R563 B.n854 B.n602 585
R564 B.n853 B.n601 585
R565 B.n858 B.n601 585
R566 B.n852 B.n851 585
R567 B.n850 B.n849 585
R568 B.n848 B.n847 585
R569 B.n846 B.n845 585
R570 B.n844 B.n843 585
R571 B.n842 B.n841 585
R572 B.n840 B.n839 585
R573 B.n838 B.n837 585
R574 B.n836 B.n835 585
R575 B.n834 B.n833 585
R576 B.n832 B.n831 585
R577 B.n830 B.n829 585
R578 B.n828 B.n827 585
R579 B.n826 B.n825 585
R580 B.n824 B.n823 585
R581 B.n822 B.n821 585
R582 B.n820 B.n819 585
R583 B.n818 B.n817 585
R584 B.n816 B.n815 585
R585 B.n814 B.n813 585
R586 B.n812 B.n811 585
R587 B.n810 B.n809 585
R588 B.n808 B.n807 585
R589 B.n806 B.n805 585
R590 B.n804 B.n803 585
R591 B.n802 B.n801 585
R592 B.n800 B.n799 585
R593 B.n798 B.n797 585
R594 B.n796 B.n795 585
R595 B.n794 B.n793 585
R596 B.n792 B.n791 585
R597 B.n790 B.n789 585
R598 B.n788 B.n787 585
R599 B.n786 B.n785 585
R600 B.n784 B.n783 585
R601 B.n782 B.n781 585
R602 B.n780 B.n779 585
R603 B.n778 B.n777 585
R604 B.n776 B.n775 585
R605 B.n774 B.n773 585
R606 B.n772 B.n771 585
R607 B.n770 B.n769 585
R608 B.n768 B.n767 585
R609 B.n766 B.n765 585
R610 B.n764 B.n763 585
R611 B.n762 B.n761 585
R612 B.n760 B.n759 585
R613 B.n758 B.n757 585
R614 B.n756 B.n755 585
R615 B.n754 B.n753 585
R616 B.n752 B.n751 585
R617 B.n750 B.n749 585
R618 B.n748 B.n747 585
R619 B.n746 B.n745 585
R620 B.n744 B.n743 585
R621 B.n742 B.n741 585
R622 B.n740 B.n739 585
R623 B.n738 B.n737 585
R624 B.n736 B.n735 585
R625 B.n734 B.n733 585
R626 B.n732 B.n731 585
R627 B.n730 B.n729 585
R628 B.n728 B.n727 585
R629 B.n726 B.n725 585
R630 B.n724 B.n723 585
R631 B.n721 B.n720 585
R632 B.n719 B.n718 585
R633 B.n717 B.n716 585
R634 B.n715 B.n714 585
R635 B.n713 B.n712 585
R636 B.n711 B.n710 585
R637 B.n709 B.n708 585
R638 B.n707 B.n706 585
R639 B.n705 B.n704 585
R640 B.n703 B.n702 585
R641 B.n701 B.n700 585
R642 B.n699 B.n698 585
R643 B.n697 B.n696 585
R644 B.n695 B.n694 585
R645 B.n693 B.n692 585
R646 B.n691 B.n690 585
R647 B.n689 B.n688 585
R648 B.n687 B.n686 585
R649 B.n685 B.n684 585
R650 B.n683 B.n682 585
R651 B.n681 B.n680 585
R652 B.n679 B.n678 585
R653 B.n677 B.n676 585
R654 B.n675 B.n674 585
R655 B.n673 B.n672 585
R656 B.n671 B.n670 585
R657 B.n669 B.n668 585
R658 B.n667 B.n666 585
R659 B.n665 B.n664 585
R660 B.n663 B.n662 585
R661 B.n661 B.n660 585
R662 B.n659 B.n658 585
R663 B.n657 B.n656 585
R664 B.n655 B.n654 585
R665 B.n653 B.n652 585
R666 B.n651 B.n650 585
R667 B.n649 B.n648 585
R668 B.n647 B.n646 585
R669 B.n645 B.n644 585
R670 B.n643 B.n642 585
R671 B.n641 B.n640 585
R672 B.n639 B.n638 585
R673 B.n637 B.n636 585
R674 B.n635 B.n634 585
R675 B.n633 B.n632 585
R676 B.n631 B.n630 585
R677 B.n629 B.n628 585
R678 B.n627 B.n626 585
R679 B.n625 B.n624 585
R680 B.n623 B.n622 585
R681 B.n621 B.n620 585
R682 B.n619 B.n618 585
R683 B.n617 B.n616 585
R684 B.n615 B.n614 585
R685 B.n613 B.n612 585
R686 B.n611 B.n610 585
R687 B.n609 B.n608 585
R688 B.n539 B.n538 585
R689 B.n861 B.n860 585
R690 B.n535 B.n534 585
R691 B.n536 B.n535 585
R692 B.n867 B.n866 585
R693 B.n866 B.n865 585
R694 B.n868 B.n533 585
R695 B.n533 B.n532 585
R696 B.n870 B.n869 585
R697 B.n871 B.n870 585
R698 B.n527 B.n526 585
R699 B.n528 B.n527 585
R700 B.n879 B.n878 585
R701 B.n878 B.n877 585
R702 B.n880 B.n525 585
R703 B.n525 B.n524 585
R704 B.n882 B.n881 585
R705 B.n883 B.n882 585
R706 B.n519 B.n518 585
R707 B.n520 B.n519 585
R708 B.n891 B.n890 585
R709 B.n890 B.n889 585
R710 B.n892 B.n517 585
R711 B.n517 B.n516 585
R712 B.n894 B.n893 585
R713 B.n895 B.n894 585
R714 B.n511 B.n510 585
R715 B.n512 B.n511 585
R716 B.n903 B.n902 585
R717 B.n902 B.n901 585
R718 B.n904 B.n509 585
R719 B.n509 B.n508 585
R720 B.n906 B.n905 585
R721 B.n907 B.n906 585
R722 B.n503 B.n502 585
R723 B.n504 B.n503 585
R724 B.n916 B.n915 585
R725 B.n915 B.n914 585
R726 B.n917 B.n501 585
R727 B.n913 B.n501 585
R728 B.n919 B.n918 585
R729 B.n920 B.n919 585
R730 B.n496 B.n495 585
R731 B.n497 B.n496 585
R732 B.n928 B.n927 585
R733 B.n927 B.n926 585
R734 B.n929 B.n494 585
R735 B.n494 B.n493 585
R736 B.n931 B.n930 585
R737 B.n932 B.n931 585
R738 B.n488 B.n487 585
R739 B.n489 B.n488 585
R740 B.n940 B.n939 585
R741 B.n939 B.n938 585
R742 B.n941 B.n486 585
R743 B.n486 B.n485 585
R744 B.n943 B.n942 585
R745 B.n944 B.n943 585
R746 B.n480 B.n479 585
R747 B.n481 B.n480 585
R748 B.n952 B.n951 585
R749 B.n951 B.n950 585
R750 B.n953 B.n478 585
R751 B.n478 B.n477 585
R752 B.n955 B.n954 585
R753 B.n956 B.n955 585
R754 B.n472 B.n471 585
R755 B.n473 B.n472 585
R756 B.n964 B.n963 585
R757 B.n963 B.n962 585
R758 B.n965 B.n470 585
R759 B.n470 B.n469 585
R760 B.n967 B.n966 585
R761 B.n968 B.n967 585
R762 B.n464 B.n463 585
R763 B.n465 B.n464 585
R764 B.n976 B.n975 585
R765 B.n975 B.n974 585
R766 B.n977 B.n462 585
R767 B.n462 B.n461 585
R768 B.n979 B.n978 585
R769 B.n980 B.n979 585
R770 B.n456 B.n455 585
R771 B.n457 B.n456 585
R772 B.n988 B.n987 585
R773 B.n987 B.n986 585
R774 B.n989 B.n454 585
R775 B.n454 B.n453 585
R776 B.n991 B.n990 585
R777 B.n992 B.n991 585
R778 B.n448 B.n447 585
R779 B.n449 B.n448 585
R780 B.n1000 B.n999 585
R781 B.n999 B.n998 585
R782 B.n1001 B.n446 585
R783 B.n446 B.n445 585
R784 B.n1003 B.n1002 585
R785 B.n1004 B.n1003 585
R786 B.n440 B.n439 585
R787 B.n441 B.n440 585
R788 B.n1012 B.n1011 585
R789 B.n1011 B.n1010 585
R790 B.n1013 B.n438 585
R791 B.n438 B.n437 585
R792 B.n1015 B.n1014 585
R793 B.n1016 B.n1015 585
R794 B.n432 B.n431 585
R795 B.n433 B.n432 585
R796 B.n1025 B.n1024 585
R797 B.n1024 B.n1023 585
R798 B.n1026 B.n430 585
R799 B.n430 B.n429 585
R800 B.n1028 B.n1027 585
R801 B.n1029 B.n1028 585
R802 B.n3 B.n0 585
R803 B.n4 B.n3 585
R804 B.n1221 B.n1 585
R805 B.n1222 B.n1221 585
R806 B.n1220 B.n1219 585
R807 B.n1220 B.n8 585
R808 B.n1218 B.n9 585
R809 B.n12 B.n9 585
R810 B.n1217 B.n1216 585
R811 B.n1216 B.n1215 585
R812 B.n11 B.n10 585
R813 B.n1214 B.n11 585
R814 B.n1212 B.n1211 585
R815 B.n1213 B.n1212 585
R816 B.n1210 B.n17 585
R817 B.n17 B.n16 585
R818 B.n1209 B.n1208 585
R819 B.n1208 B.n1207 585
R820 B.n19 B.n18 585
R821 B.n1206 B.n19 585
R822 B.n1204 B.n1203 585
R823 B.n1205 B.n1204 585
R824 B.n1202 B.n24 585
R825 B.n24 B.n23 585
R826 B.n1201 B.n1200 585
R827 B.n1200 B.n1199 585
R828 B.n26 B.n25 585
R829 B.n1198 B.n26 585
R830 B.n1196 B.n1195 585
R831 B.n1197 B.n1196 585
R832 B.n1194 B.n31 585
R833 B.n31 B.n30 585
R834 B.n1193 B.n1192 585
R835 B.n1192 B.n1191 585
R836 B.n33 B.n32 585
R837 B.n1190 B.n33 585
R838 B.n1188 B.n1187 585
R839 B.n1189 B.n1188 585
R840 B.n1186 B.n38 585
R841 B.n38 B.n37 585
R842 B.n1185 B.n1184 585
R843 B.n1184 B.n1183 585
R844 B.n40 B.n39 585
R845 B.n1182 B.n40 585
R846 B.n1180 B.n1179 585
R847 B.n1181 B.n1180 585
R848 B.n1178 B.n45 585
R849 B.n45 B.n44 585
R850 B.n1177 B.n1176 585
R851 B.n1176 B.n1175 585
R852 B.n47 B.n46 585
R853 B.n1174 B.n47 585
R854 B.n1172 B.n1171 585
R855 B.n1173 B.n1172 585
R856 B.n1170 B.n52 585
R857 B.n52 B.n51 585
R858 B.n1169 B.n1168 585
R859 B.n1168 B.n1167 585
R860 B.n54 B.n53 585
R861 B.n1166 B.n54 585
R862 B.n1164 B.n1163 585
R863 B.n1165 B.n1164 585
R864 B.n1162 B.n59 585
R865 B.n59 B.n58 585
R866 B.n1161 B.n1160 585
R867 B.n1160 B.n1159 585
R868 B.n61 B.n60 585
R869 B.n1158 B.n61 585
R870 B.n1156 B.n1155 585
R871 B.n1157 B.n1156 585
R872 B.n1154 B.n66 585
R873 B.n66 B.n65 585
R874 B.n1153 B.n1152 585
R875 B.n1152 B.n1151 585
R876 B.n68 B.n67 585
R877 B.n1150 B.n68 585
R878 B.n1148 B.n1147 585
R879 B.n1149 B.n1148 585
R880 B.n1146 B.n72 585
R881 B.n75 B.n72 585
R882 B.n1145 B.n1144 585
R883 B.n1144 B.n1143 585
R884 B.n74 B.n73 585
R885 B.n1142 B.n74 585
R886 B.n1140 B.n1139 585
R887 B.n1141 B.n1140 585
R888 B.n1138 B.n80 585
R889 B.n80 B.n79 585
R890 B.n1137 B.n1136 585
R891 B.n1136 B.n1135 585
R892 B.n82 B.n81 585
R893 B.n1134 B.n82 585
R894 B.n1132 B.n1131 585
R895 B.n1133 B.n1132 585
R896 B.n1130 B.n87 585
R897 B.n87 B.n86 585
R898 B.n1129 B.n1128 585
R899 B.n1128 B.n1127 585
R900 B.n89 B.n88 585
R901 B.n1126 B.n89 585
R902 B.n1124 B.n1123 585
R903 B.n1125 B.n1124 585
R904 B.n1122 B.n94 585
R905 B.n94 B.n93 585
R906 B.n1121 B.n1120 585
R907 B.n1120 B.n1119 585
R908 B.n96 B.n95 585
R909 B.n1118 B.n96 585
R910 B.n1116 B.n1115 585
R911 B.n1117 B.n1116 585
R912 B.n1114 B.n101 585
R913 B.n101 B.n100 585
R914 B.n1113 B.n1112 585
R915 B.n1112 B.n1111 585
R916 B.n103 B.n102 585
R917 B.n1110 B.n103 585
R918 B.n1225 B.n1224 585
R919 B.n1223 B.n2 585
R920 B.n175 B.n103 492.5
R921 B.n1108 B.n105 492.5
R922 B.n860 B.n537 492.5
R923 B.n856 B.n535 492.5
R924 B.n173 B.t18 382.697
R925 B.n170 B.t10 382.697
R926 B.n606 B.t21 382.697
R927 B.n603 B.t14 382.697
R928 B.n1109 B.n168 256.663
R929 B.n1109 B.n167 256.663
R930 B.n1109 B.n166 256.663
R931 B.n1109 B.n165 256.663
R932 B.n1109 B.n164 256.663
R933 B.n1109 B.n163 256.663
R934 B.n1109 B.n162 256.663
R935 B.n1109 B.n161 256.663
R936 B.n1109 B.n160 256.663
R937 B.n1109 B.n159 256.663
R938 B.n1109 B.n158 256.663
R939 B.n1109 B.n157 256.663
R940 B.n1109 B.n156 256.663
R941 B.n1109 B.n155 256.663
R942 B.n1109 B.n154 256.663
R943 B.n1109 B.n153 256.663
R944 B.n1109 B.n152 256.663
R945 B.n1109 B.n151 256.663
R946 B.n1109 B.n150 256.663
R947 B.n1109 B.n149 256.663
R948 B.n1109 B.n148 256.663
R949 B.n1109 B.n147 256.663
R950 B.n1109 B.n146 256.663
R951 B.n1109 B.n145 256.663
R952 B.n1109 B.n144 256.663
R953 B.n1109 B.n143 256.663
R954 B.n1109 B.n142 256.663
R955 B.n1109 B.n141 256.663
R956 B.n1109 B.n140 256.663
R957 B.n1109 B.n139 256.663
R958 B.n1109 B.n138 256.663
R959 B.n1109 B.n137 256.663
R960 B.n1109 B.n136 256.663
R961 B.n1109 B.n135 256.663
R962 B.n1109 B.n134 256.663
R963 B.n1109 B.n133 256.663
R964 B.n1109 B.n132 256.663
R965 B.n1109 B.n131 256.663
R966 B.n1109 B.n130 256.663
R967 B.n1109 B.n129 256.663
R968 B.n1109 B.n128 256.663
R969 B.n1109 B.n127 256.663
R970 B.n1109 B.n126 256.663
R971 B.n1109 B.n125 256.663
R972 B.n1109 B.n124 256.663
R973 B.n1109 B.n123 256.663
R974 B.n1109 B.n122 256.663
R975 B.n1109 B.n121 256.663
R976 B.n1109 B.n120 256.663
R977 B.n1109 B.n119 256.663
R978 B.n1109 B.n118 256.663
R979 B.n1109 B.n117 256.663
R980 B.n1109 B.n116 256.663
R981 B.n1109 B.n115 256.663
R982 B.n1109 B.n114 256.663
R983 B.n1109 B.n113 256.663
R984 B.n1109 B.n112 256.663
R985 B.n1109 B.n111 256.663
R986 B.n1109 B.n110 256.663
R987 B.n1109 B.n109 256.663
R988 B.n1109 B.n108 256.663
R989 B.n1109 B.n107 256.663
R990 B.n1109 B.n106 256.663
R991 B.n858 B.n857 256.663
R992 B.n858 B.n540 256.663
R993 B.n858 B.n541 256.663
R994 B.n858 B.n542 256.663
R995 B.n858 B.n543 256.663
R996 B.n858 B.n544 256.663
R997 B.n858 B.n545 256.663
R998 B.n858 B.n546 256.663
R999 B.n858 B.n547 256.663
R1000 B.n858 B.n548 256.663
R1001 B.n858 B.n549 256.663
R1002 B.n858 B.n550 256.663
R1003 B.n858 B.n551 256.663
R1004 B.n858 B.n552 256.663
R1005 B.n858 B.n553 256.663
R1006 B.n858 B.n554 256.663
R1007 B.n858 B.n555 256.663
R1008 B.n858 B.n556 256.663
R1009 B.n858 B.n557 256.663
R1010 B.n858 B.n558 256.663
R1011 B.n858 B.n559 256.663
R1012 B.n858 B.n560 256.663
R1013 B.n858 B.n561 256.663
R1014 B.n858 B.n562 256.663
R1015 B.n858 B.n563 256.663
R1016 B.n858 B.n564 256.663
R1017 B.n858 B.n565 256.663
R1018 B.n858 B.n566 256.663
R1019 B.n858 B.n567 256.663
R1020 B.n858 B.n568 256.663
R1021 B.n858 B.n569 256.663
R1022 B.n858 B.n570 256.663
R1023 B.n858 B.n571 256.663
R1024 B.n858 B.n572 256.663
R1025 B.n858 B.n573 256.663
R1026 B.n858 B.n574 256.663
R1027 B.n858 B.n575 256.663
R1028 B.n858 B.n576 256.663
R1029 B.n858 B.n577 256.663
R1030 B.n858 B.n578 256.663
R1031 B.n858 B.n579 256.663
R1032 B.n858 B.n580 256.663
R1033 B.n858 B.n581 256.663
R1034 B.n858 B.n582 256.663
R1035 B.n858 B.n583 256.663
R1036 B.n858 B.n584 256.663
R1037 B.n858 B.n585 256.663
R1038 B.n858 B.n586 256.663
R1039 B.n858 B.n587 256.663
R1040 B.n858 B.n588 256.663
R1041 B.n858 B.n589 256.663
R1042 B.n858 B.n590 256.663
R1043 B.n858 B.n591 256.663
R1044 B.n858 B.n592 256.663
R1045 B.n858 B.n593 256.663
R1046 B.n858 B.n594 256.663
R1047 B.n858 B.n595 256.663
R1048 B.n858 B.n596 256.663
R1049 B.n858 B.n597 256.663
R1050 B.n858 B.n598 256.663
R1051 B.n858 B.n599 256.663
R1052 B.n858 B.n600 256.663
R1053 B.n859 B.n858 256.663
R1054 B.n1227 B.n1226 256.663
R1055 B.n179 B.n178 163.367
R1056 B.n183 B.n182 163.367
R1057 B.n187 B.n186 163.367
R1058 B.n191 B.n190 163.367
R1059 B.n195 B.n194 163.367
R1060 B.n199 B.n198 163.367
R1061 B.n203 B.n202 163.367
R1062 B.n207 B.n206 163.367
R1063 B.n211 B.n210 163.367
R1064 B.n215 B.n214 163.367
R1065 B.n219 B.n218 163.367
R1066 B.n223 B.n222 163.367
R1067 B.n227 B.n226 163.367
R1068 B.n231 B.n230 163.367
R1069 B.n235 B.n234 163.367
R1070 B.n239 B.n238 163.367
R1071 B.n243 B.n242 163.367
R1072 B.n247 B.n246 163.367
R1073 B.n251 B.n250 163.367
R1074 B.n255 B.n254 163.367
R1075 B.n259 B.n258 163.367
R1076 B.n263 B.n262 163.367
R1077 B.n267 B.n266 163.367
R1078 B.n271 B.n270 163.367
R1079 B.n275 B.n274 163.367
R1080 B.n279 B.n278 163.367
R1081 B.n283 B.n282 163.367
R1082 B.n287 B.n286 163.367
R1083 B.n291 B.n290 163.367
R1084 B.n296 B.n295 163.367
R1085 B.n300 B.n299 163.367
R1086 B.n304 B.n303 163.367
R1087 B.n308 B.n307 163.367
R1088 B.n312 B.n311 163.367
R1089 B.n316 B.n315 163.367
R1090 B.n320 B.n319 163.367
R1091 B.n324 B.n323 163.367
R1092 B.n328 B.n327 163.367
R1093 B.n332 B.n331 163.367
R1094 B.n336 B.n335 163.367
R1095 B.n340 B.n339 163.367
R1096 B.n344 B.n343 163.367
R1097 B.n348 B.n347 163.367
R1098 B.n352 B.n351 163.367
R1099 B.n356 B.n355 163.367
R1100 B.n360 B.n359 163.367
R1101 B.n364 B.n363 163.367
R1102 B.n368 B.n367 163.367
R1103 B.n372 B.n371 163.367
R1104 B.n376 B.n375 163.367
R1105 B.n380 B.n379 163.367
R1106 B.n384 B.n383 163.367
R1107 B.n388 B.n387 163.367
R1108 B.n392 B.n391 163.367
R1109 B.n396 B.n395 163.367
R1110 B.n400 B.n399 163.367
R1111 B.n404 B.n403 163.367
R1112 B.n408 B.n407 163.367
R1113 B.n412 B.n411 163.367
R1114 B.n416 B.n415 163.367
R1115 B.n420 B.n419 163.367
R1116 B.n424 B.n423 163.367
R1117 B.n1108 B.n169 163.367
R1118 B.n864 B.n537 163.367
R1119 B.n864 B.n531 163.367
R1120 B.n872 B.n531 163.367
R1121 B.n872 B.n529 163.367
R1122 B.n876 B.n529 163.367
R1123 B.n876 B.n523 163.367
R1124 B.n884 B.n523 163.367
R1125 B.n884 B.n521 163.367
R1126 B.n888 B.n521 163.367
R1127 B.n888 B.n515 163.367
R1128 B.n896 B.n515 163.367
R1129 B.n896 B.n513 163.367
R1130 B.n900 B.n513 163.367
R1131 B.n900 B.n507 163.367
R1132 B.n908 B.n507 163.367
R1133 B.n908 B.n505 163.367
R1134 B.n912 B.n505 163.367
R1135 B.n912 B.n500 163.367
R1136 B.n921 B.n500 163.367
R1137 B.n921 B.n498 163.367
R1138 B.n925 B.n498 163.367
R1139 B.n925 B.n492 163.367
R1140 B.n933 B.n492 163.367
R1141 B.n933 B.n490 163.367
R1142 B.n937 B.n490 163.367
R1143 B.n937 B.n484 163.367
R1144 B.n945 B.n484 163.367
R1145 B.n945 B.n482 163.367
R1146 B.n949 B.n482 163.367
R1147 B.n949 B.n476 163.367
R1148 B.n957 B.n476 163.367
R1149 B.n957 B.n474 163.367
R1150 B.n961 B.n474 163.367
R1151 B.n961 B.n468 163.367
R1152 B.n969 B.n468 163.367
R1153 B.n969 B.n466 163.367
R1154 B.n973 B.n466 163.367
R1155 B.n973 B.n460 163.367
R1156 B.n981 B.n460 163.367
R1157 B.n981 B.n458 163.367
R1158 B.n985 B.n458 163.367
R1159 B.n985 B.n452 163.367
R1160 B.n993 B.n452 163.367
R1161 B.n993 B.n450 163.367
R1162 B.n997 B.n450 163.367
R1163 B.n997 B.n444 163.367
R1164 B.n1005 B.n444 163.367
R1165 B.n1005 B.n442 163.367
R1166 B.n1009 B.n442 163.367
R1167 B.n1009 B.n436 163.367
R1168 B.n1017 B.n436 163.367
R1169 B.n1017 B.n434 163.367
R1170 B.n1022 B.n434 163.367
R1171 B.n1022 B.n428 163.367
R1172 B.n1030 B.n428 163.367
R1173 B.n1031 B.n1030 163.367
R1174 B.n1031 B.n5 163.367
R1175 B.n6 B.n5 163.367
R1176 B.n7 B.n6 163.367
R1177 B.n1037 B.n7 163.367
R1178 B.n1038 B.n1037 163.367
R1179 B.n1038 B.n13 163.367
R1180 B.n14 B.n13 163.367
R1181 B.n15 B.n14 163.367
R1182 B.n1043 B.n15 163.367
R1183 B.n1043 B.n20 163.367
R1184 B.n21 B.n20 163.367
R1185 B.n22 B.n21 163.367
R1186 B.n1048 B.n22 163.367
R1187 B.n1048 B.n27 163.367
R1188 B.n28 B.n27 163.367
R1189 B.n29 B.n28 163.367
R1190 B.n1053 B.n29 163.367
R1191 B.n1053 B.n34 163.367
R1192 B.n35 B.n34 163.367
R1193 B.n36 B.n35 163.367
R1194 B.n1058 B.n36 163.367
R1195 B.n1058 B.n41 163.367
R1196 B.n42 B.n41 163.367
R1197 B.n43 B.n42 163.367
R1198 B.n1063 B.n43 163.367
R1199 B.n1063 B.n48 163.367
R1200 B.n49 B.n48 163.367
R1201 B.n50 B.n49 163.367
R1202 B.n1068 B.n50 163.367
R1203 B.n1068 B.n55 163.367
R1204 B.n56 B.n55 163.367
R1205 B.n57 B.n56 163.367
R1206 B.n1073 B.n57 163.367
R1207 B.n1073 B.n62 163.367
R1208 B.n63 B.n62 163.367
R1209 B.n64 B.n63 163.367
R1210 B.n1078 B.n64 163.367
R1211 B.n1078 B.n69 163.367
R1212 B.n70 B.n69 163.367
R1213 B.n71 B.n70 163.367
R1214 B.n1083 B.n71 163.367
R1215 B.n1083 B.n76 163.367
R1216 B.n77 B.n76 163.367
R1217 B.n78 B.n77 163.367
R1218 B.n1088 B.n78 163.367
R1219 B.n1088 B.n83 163.367
R1220 B.n84 B.n83 163.367
R1221 B.n85 B.n84 163.367
R1222 B.n1093 B.n85 163.367
R1223 B.n1093 B.n90 163.367
R1224 B.n91 B.n90 163.367
R1225 B.n92 B.n91 163.367
R1226 B.n1098 B.n92 163.367
R1227 B.n1098 B.n97 163.367
R1228 B.n98 B.n97 163.367
R1229 B.n99 B.n98 163.367
R1230 B.n1103 B.n99 163.367
R1231 B.n1103 B.n104 163.367
R1232 B.n105 B.n104 163.367
R1233 B.n602 B.n601 163.367
R1234 B.n851 B.n601 163.367
R1235 B.n849 B.n848 163.367
R1236 B.n845 B.n844 163.367
R1237 B.n841 B.n840 163.367
R1238 B.n837 B.n836 163.367
R1239 B.n833 B.n832 163.367
R1240 B.n829 B.n828 163.367
R1241 B.n825 B.n824 163.367
R1242 B.n821 B.n820 163.367
R1243 B.n817 B.n816 163.367
R1244 B.n813 B.n812 163.367
R1245 B.n809 B.n808 163.367
R1246 B.n805 B.n804 163.367
R1247 B.n801 B.n800 163.367
R1248 B.n797 B.n796 163.367
R1249 B.n793 B.n792 163.367
R1250 B.n789 B.n788 163.367
R1251 B.n785 B.n784 163.367
R1252 B.n781 B.n780 163.367
R1253 B.n777 B.n776 163.367
R1254 B.n773 B.n772 163.367
R1255 B.n769 B.n768 163.367
R1256 B.n765 B.n764 163.367
R1257 B.n761 B.n760 163.367
R1258 B.n757 B.n756 163.367
R1259 B.n753 B.n752 163.367
R1260 B.n749 B.n748 163.367
R1261 B.n745 B.n744 163.367
R1262 B.n741 B.n740 163.367
R1263 B.n737 B.n736 163.367
R1264 B.n733 B.n732 163.367
R1265 B.n729 B.n728 163.367
R1266 B.n725 B.n724 163.367
R1267 B.n720 B.n719 163.367
R1268 B.n716 B.n715 163.367
R1269 B.n712 B.n711 163.367
R1270 B.n708 B.n707 163.367
R1271 B.n704 B.n703 163.367
R1272 B.n700 B.n699 163.367
R1273 B.n696 B.n695 163.367
R1274 B.n692 B.n691 163.367
R1275 B.n688 B.n687 163.367
R1276 B.n684 B.n683 163.367
R1277 B.n680 B.n679 163.367
R1278 B.n676 B.n675 163.367
R1279 B.n672 B.n671 163.367
R1280 B.n668 B.n667 163.367
R1281 B.n664 B.n663 163.367
R1282 B.n660 B.n659 163.367
R1283 B.n656 B.n655 163.367
R1284 B.n652 B.n651 163.367
R1285 B.n648 B.n647 163.367
R1286 B.n644 B.n643 163.367
R1287 B.n640 B.n639 163.367
R1288 B.n636 B.n635 163.367
R1289 B.n632 B.n631 163.367
R1290 B.n628 B.n627 163.367
R1291 B.n624 B.n623 163.367
R1292 B.n620 B.n619 163.367
R1293 B.n616 B.n615 163.367
R1294 B.n612 B.n611 163.367
R1295 B.n608 B.n539 163.367
R1296 B.n866 B.n535 163.367
R1297 B.n866 B.n533 163.367
R1298 B.n870 B.n533 163.367
R1299 B.n870 B.n527 163.367
R1300 B.n878 B.n527 163.367
R1301 B.n878 B.n525 163.367
R1302 B.n882 B.n525 163.367
R1303 B.n882 B.n519 163.367
R1304 B.n890 B.n519 163.367
R1305 B.n890 B.n517 163.367
R1306 B.n894 B.n517 163.367
R1307 B.n894 B.n511 163.367
R1308 B.n902 B.n511 163.367
R1309 B.n902 B.n509 163.367
R1310 B.n906 B.n509 163.367
R1311 B.n906 B.n503 163.367
R1312 B.n915 B.n503 163.367
R1313 B.n915 B.n501 163.367
R1314 B.n919 B.n501 163.367
R1315 B.n919 B.n496 163.367
R1316 B.n927 B.n496 163.367
R1317 B.n927 B.n494 163.367
R1318 B.n931 B.n494 163.367
R1319 B.n931 B.n488 163.367
R1320 B.n939 B.n488 163.367
R1321 B.n939 B.n486 163.367
R1322 B.n943 B.n486 163.367
R1323 B.n943 B.n480 163.367
R1324 B.n951 B.n480 163.367
R1325 B.n951 B.n478 163.367
R1326 B.n955 B.n478 163.367
R1327 B.n955 B.n472 163.367
R1328 B.n963 B.n472 163.367
R1329 B.n963 B.n470 163.367
R1330 B.n967 B.n470 163.367
R1331 B.n967 B.n464 163.367
R1332 B.n975 B.n464 163.367
R1333 B.n975 B.n462 163.367
R1334 B.n979 B.n462 163.367
R1335 B.n979 B.n456 163.367
R1336 B.n987 B.n456 163.367
R1337 B.n987 B.n454 163.367
R1338 B.n991 B.n454 163.367
R1339 B.n991 B.n448 163.367
R1340 B.n999 B.n448 163.367
R1341 B.n999 B.n446 163.367
R1342 B.n1003 B.n446 163.367
R1343 B.n1003 B.n440 163.367
R1344 B.n1011 B.n440 163.367
R1345 B.n1011 B.n438 163.367
R1346 B.n1015 B.n438 163.367
R1347 B.n1015 B.n432 163.367
R1348 B.n1024 B.n432 163.367
R1349 B.n1024 B.n430 163.367
R1350 B.n1028 B.n430 163.367
R1351 B.n1028 B.n3 163.367
R1352 B.n1225 B.n3 163.367
R1353 B.n1221 B.n2 163.367
R1354 B.n1221 B.n1220 163.367
R1355 B.n1220 B.n9 163.367
R1356 B.n1216 B.n9 163.367
R1357 B.n1216 B.n11 163.367
R1358 B.n1212 B.n11 163.367
R1359 B.n1212 B.n17 163.367
R1360 B.n1208 B.n17 163.367
R1361 B.n1208 B.n19 163.367
R1362 B.n1204 B.n19 163.367
R1363 B.n1204 B.n24 163.367
R1364 B.n1200 B.n24 163.367
R1365 B.n1200 B.n26 163.367
R1366 B.n1196 B.n26 163.367
R1367 B.n1196 B.n31 163.367
R1368 B.n1192 B.n31 163.367
R1369 B.n1192 B.n33 163.367
R1370 B.n1188 B.n33 163.367
R1371 B.n1188 B.n38 163.367
R1372 B.n1184 B.n38 163.367
R1373 B.n1184 B.n40 163.367
R1374 B.n1180 B.n40 163.367
R1375 B.n1180 B.n45 163.367
R1376 B.n1176 B.n45 163.367
R1377 B.n1176 B.n47 163.367
R1378 B.n1172 B.n47 163.367
R1379 B.n1172 B.n52 163.367
R1380 B.n1168 B.n52 163.367
R1381 B.n1168 B.n54 163.367
R1382 B.n1164 B.n54 163.367
R1383 B.n1164 B.n59 163.367
R1384 B.n1160 B.n59 163.367
R1385 B.n1160 B.n61 163.367
R1386 B.n1156 B.n61 163.367
R1387 B.n1156 B.n66 163.367
R1388 B.n1152 B.n66 163.367
R1389 B.n1152 B.n68 163.367
R1390 B.n1148 B.n68 163.367
R1391 B.n1148 B.n72 163.367
R1392 B.n1144 B.n72 163.367
R1393 B.n1144 B.n74 163.367
R1394 B.n1140 B.n74 163.367
R1395 B.n1140 B.n80 163.367
R1396 B.n1136 B.n80 163.367
R1397 B.n1136 B.n82 163.367
R1398 B.n1132 B.n82 163.367
R1399 B.n1132 B.n87 163.367
R1400 B.n1128 B.n87 163.367
R1401 B.n1128 B.n89 163.367
R1402 B.n1124 B.n89 163.367
R1403 B.n1124 B.n94 163.367
R1404 B.n1120 B.n94 163.367
R1405 B.n1120 B.n96 163.367
R1406 B.n1116 B.n96 163.367
R1407 B.n1116 B.n101 163.367
R1408 B.n1112 B.n101 163.367
R1409 B.n1112 B.n103 163.367
R1410 B.n170 B.t12 124.663
R1411 B.n606 B.t23 124.663
R1412 B.n173 B.t19 124.639
R1413 B.n603 B.t17 124.639
R1414 B.n175 B.n106 71.676
R1415 B.n179 B.n107 71.676
R1416 B.n183 B.n108 71.676
R1417 B.n187 B.n109 71.676
R1418 B.n191 B.n110 71.676
R1419 B.n195 B.n111 71.676
R1420 B.n199 B.n112 71.676
R1421 B.n203 B.n113 71.676
R1422 B.n207 B.n114 71.676
R1423 B.n211 B.n115 71.676
R1424 B.n215 B.n116 71.676
R1425 B.n219 B.n117 71.676
R1426 B.n223 B.n118 71.676
R1427 B.n227 B.n119 71.676
R1428 B.n231 B.n120 71.676
R1429 B.n235 B.n121 71.676
R1430 B.n239 B.n122 71.676
R1431 B.n243 B.n123 71.676
R1432 B.n247 B.n124 71.676
R1433 B.n251 B.n125 71.676
R1434 B.n255 B.n126 71.676
R1435 B.n259 B.n127 71.676
R1436 B.n263 B.n128 71.676
R1437 B.n267 B.n129 71.676
R1438 B.n271 B.n130 71.676
R1439 B.n275 B.n131 71.676
R1440 B.n279 B.n132 71.676
R1441 B.n283 B.n133 71.676
R1442 B.n287 B.n134 71.676
R1443 B.n291 B.n135 71.676
R1444 B.n296 B.n136 71.676
R1445 B.n300 B.n137 71.676
R1446 B.n304 B.n138 71.676
R1447 B.n308 B.n139 71.676
R1448 B.n312 B.n140 71.676
R1449 B.n316 B.n141 71.676
R1450 B.n320 B.n142 71.676
R1451 B.n324 B.n143 71.676
R1452 B.n328 B.n144 71.676
R1453 B.n332 B.n145 71.676
R1454 B.n336 B.n146 71.676
R1455 B.n340 B.n147 71.676
R1456 B.n344 B.n148 71.676
R1457 B.n348 B.n149 71.676
R1458 B.n352 B.n150 71.676
R1459 B.n356 B.n151 71.676
R1460 B.n360 B.n152 71.676
R1461 B.n364 B.n153 71.676
R1462 B.n368 B.n154 71.676
R1463 B.n372 B.n155 71.676
R1464 B.n376 B.n156 71.676
R1465 B.n380 B.n157 71.676
R1466 B.n384 B.n158 71.676
R1467 B.n388 B.n159 71.676
R1468 B.n392 B.n160 71.676
R1469 B.n396 B.n161 71.676
R1470 B.n400 B.n162 71.676
R1471 B.n404 B.n163 71.676
R1472 B.n408 B.n164 71.676
R1473 B.n412 B.n165 71.676
R1474 B.n416 B.n166 71.676
R1475 B.n420 B.n167 71.676
R1476 B.n424 B.n168 71.676
R1477 B.n169 B.n168 71.676
R1478 B.n423 B.n167 71.676
R1479 B.n419 B.n166 71.676
R1480 B.n415 B.n165 71.676
R1481 B.n411 B.n164 71.676
R1482 B.n407 B.n163 71.676
R1483 B.n403 B.n162 71.676
R1484 B.n399 B.n161 71.676
R1485 B.n395 B.n160 71.676
R1486 B.n391 B.n159 71.676
R1487 B.n387 B.n158 71.676
R1488 B.n383 B.n157 71.676
R1489 B.n379 B.n156 71.676
R1490 B.n375 B.n155 71.676
R1491 B.n371 B.n154 71.676
R1492 B.n367 B.n153 71.676
R1493 B.n363 B.n152 71.676
R1494 B.n359 B.n151 71.676
R1495 B.n355 B.n150 71.676
R1496 B.n351 B.n149 71.676
R1497 B.n347 B.n148 71.676
R1498 B.n343 B.n147 71.676
R1499 B.n339 B.n146 71.676
R1500 B.n335 B.n145 71.676
R1501 B.n331 B.n144 71.676
R1502 B.n327 B.n143 71.676
R1503 B.n323 B.n142 71.676
R1504 B.n319 B.n141 71.676
R1505 B.n315 B.n140 71.676
R1506 B.n311 B.n139 71.676
R1507 B.n307 B.n138 71.676
R1508 B.n303 B.n137 71.676
R1509 B.n299 B.n136 71.676
R1510 B.n295 B.n135 71.676
R1511 B.n290 B.n134 71.676
R1512 B.n286 B.n133 71.676
R1513 B.n282 B.n132 71.676
R1514 B.n278 B.n131 71.676
R1515 B.n274 B.n130 71.676
R1516 B.n270 B.n129 71.676
R1517 B.n266 B.n128 71.676
R1518 B.n262 B.n127 71.676
R1519 B.n258 B.n126 71.676
R1520 B.n254 B.n125 71.676
R1521 B.n250 B.n124 71.676
R1522 B.n246 B.n123 71.676
R1523 B.n242 B.n122 71.676
R1524 B.n238 B.n121 71.676
R1525 B.n234 B.n120 71.676
R1526 B.n230 B.n119 71.676
R1527 B.n226 B.n118 71.676
R1528 B.n222 B.n117 71.676
R1529 B.n218 B.n116 71.676
R1530 B.n214 B.n115 71.676
R1531 B.n210 B.n114 71.676
R1532 B.n206 B.n113 71.676
R1533 B.n202 B.n112 71.676
R1534 B.n198 B.n111 71.676
R1535 B.n194 B.n110 71.676
R1536 B.n190 B.n109 71.676
R1537 B.n186 B.n108 71.676
R1538 B.n182 B.n107 71.676
R1539 B.n178 B.n106 71.676
R1540 B.n857 B.n856 71.676
R1541 B.n851 B.n540 71.676
R1542 B.n848 B.n541 71.676
R1543 B.n844 B.n542 71.676
R1544 B.n840 B.n543 71.676
R1545 B.n836 B.n544 71.676
R1546 B.n832 B.n545 71.676
R1547 B.n828 B.n546 71.676
R1548 B.n824 B.n547 71.676
R1549 B.n820 B.n548 71.676
R1550 B.n816 B.n549 71.676
R1551 B.n812 B.n550 71.676
R1552 B.n808 B.n551 71.676
R1553 B.n804 B.n552 71.676
R1554 B.n800 B.n553 71.676
R1555 B.n796 B.n554 71.676
R1556 B.n792 B.n555 71.676
R1557 B.n788 B.n556 71.676
R1558 B.n784 B.n557 71.676
R1559 B.n780 B.n558 71.676
R1560 B.n776 B.n559 71.676
R1561 B.n772 B.n560 71.676
R1562 B.n768 B.n561 71.676
R1563 B.n764 B.n562 71.676
R1564 B.n760 B.n563 71.676
R1565 B.n756 B.n564 71.676
R1566 B.n752 B.n565 71.676
R1567 B.n748 B.n566 71.676
R1568 B.n744 B.n567 71.676
R1569 B.n740 B.n568 71.676
R1570 B.n736 B.n569 71.676
R1571 B.n732 B.n570 71.676
R1572 B.n728 B.n571 71.676
R1573 B.n724 B.n572 71.676
R1574 B.n719 B.n573 71.676
R1575 B.n715 B.n574 71.676
R1576 B.n711 B.n575 71.676
R1577 B.n707 B.n576 71.676
R1578 B.n703 B.n577 71.676
R1579 B.n699 B.n578 71.676
R1580 B.n695 B.n579 71.676
R1581 B.n691 B.n580 71.676
R1582 B.n687 B.n581 71.676
R1583 B.n683 B.n582 71.676
R1584 B.n679 B.n583 71.676
R1585 B.n675 B.n584 71.676
R1586 B.n671 B.n585 71.676
R1587 B.n667 B.n586 71.676
R1588 B.n663 B.n587 71.676
R1589 B.n659 B.n588 71.676
R1590 B.n655 B.n589 71.676
R1591 B.n651 B.n590 71.676
R1592 B.n647 B.n591 71.676
R1593 B.n643 B.n592 71.676
R1594 B.n639 B.n593 71.676
R1595 B.n635 B.n594 71.676
R1596 B.n631 B.n595 71.676
R1597 B.n627 B.n596 71.676
R1598 B.n623 B.n597 71.676
R1599 B.n619 B.n598 71.676
R1600 B.n615 B.n599 71.676
R1601 B.n611 B.n600 71.676
R1602 B.n859 B.n539 71.676
R1603 B.n857 B.n602 71.676
R1604 B.n849 B.n540 71.676
R1605 B.n845 B.n541 71.676
R1606 B.n841 B.n542 71.676
R1607 B.n837 B.n543 71.676
R1608 B.n833 B.n544 71.676
R1609 B.n829 B.n545 71.676
R1610 B.n825 B.n546 71.676
R1611 B.n821 B.n547 71.676
R1612 B.n817 B.n548 71.676
R1613 B.n813 B.n549 71.676
R1614 B.n809 B.n550 71.676
R1615 B.n805 B.n551 71.676
R1616 B.n801 B.n552 71.676
R1617 B.n797 B.n553 71.676
R1618 B.n793 B.n554 71.676
R1619 B.n789 B.n555 71.676
R1620 B.n785 B.n556 71.676
R1621 B.n781 B.n557 71.676
R1622 B.n777 B.n558 71.676
R1623 B.n773 B.n559 71.676
R1624 B.n769 B.n560 71.676
R1625 B.n765 B.n561 71.676
R1626 B.n761 B.n562 71.676
R1627 B.n757 B.n563 71.676
R1628 B.n753 B.n564 71.676
R1629 B.n749 B.n565 71.676
R1630 B.n745 B.n566 71.676
R1631 B.n741 B.n567 71.676
R1632 B.n737 B.n568 71.676
R1633 B.n733 B.n569 71.676
R1634 B.n729 B.n570 71.676
R1635 B.n725 B.n571 71.676
R1636 B.n720 B.n572 71.676
R1637 B.n716 B.n573 71.676
R1638 B.n712 B.n574 71.676
R1639 B.n708 B.n575 71.676
R1640 B.n704 B.n576 71.676
R1641 B.n700 B.n577 71.676
R1642 B.n696 B.n578 71.676
R1643 B.n692 B.n579 71.676
R1644 B.n688 B.n580 71.676
R1645 B.n684 B.n581 71.676
R1646 B.n680 B.n582 71.676
R1647 B.n676 B.n583 71.676
R1648 B.n672 B.n584 71.676
R1649 B.n668 B.n585 71.676
R1650 B.n664 B.n586 71.676
R1651 B.n660 B.n587 71.676
R1652 B.n656 B.n588 71.676
R1653 B.n652 B.n589 71.676
R1654 B.n648 B.n590 71.676
R1655 B.n644 B.n591 71.676
R1656 B.n640 B.n592 71.676
R1657 B.n636 B.n593 71.676
R1658 B.n632 B.n594 71.676
R1659 B.n628 B.n595 71.676
R1660 B.n624 B.n596 71.676
R1661 B.n620 B.n597 71.676
R1662 B.n616 B.n598 71.676
R1663 B.n612 B.n599 71.676
R1664 B.n608 B.n600 71.676
R1665 B.n860 B.n859 71.676
R1666 B.n1226 B.n1225 71.676
R1667 B.n1226 B.n2 71.676
R1668 B.n171 B.t13 70.5546
R1669 B.n607 B.t22 70.5546
R1670 B.n174 B.t20 70.5309
R1671 B.n604 B.t16 70.5309
R1672 B.n293 B.n174 59.5399
R1673 B.n172 B.n171 59.5399
R1674 B.n722 B.n607 59.5399
R1675 B.n605 B.n604 59.5399
R1676 B.n174 B.n173 54.1096
R1677 B.n171 B.n170 54.1096
R1678 B.n607 B.n606 54.1096
R1679 B.n604 B.n603 54.1096
R1680 B.n858 B.n536 53.7519
R1681 B.n1110 B.n1109 53.7519
R1682 B.n865 B.n536 32.3464
R1683 B.n865 B.n532 32.3464
R1684 B.n871 B.n532 32.3464
R1685 B.n871 B.n528 32.3464
R1686 B.n877 B.n528 32.3464
R1687 B.n877 B.n524 32.3464
R1688 B.n883 B.n524 32.3464
R1689 B.n889 B.n520 32.3464
R1690 B.n889 B.n516 32.3464
R1691 B.n895 B.n516 32.3464
R1692 B.n895 B.n512 32.3464
R1693 B.n901 B.n512 32.3464
R1694 B.n901 B.n508 32.3464
R1695 B.n907 B.n508 32.3464
R1696 B.n907 B.n504 32.3464
R1697 B.n914 B.n504 32.3464
R1698 B.n914 B.n913 32.3464
R1699 B.n920 B.n497 32.3464
R1700 B.n926 B.n497 32.3464
R1701 B.n926 B.n493 32.3464
R1702 B.n932 B.n493 32.3464
R1703 B.n932 B.n489 32.3464
R1704 B.n938 B.n489 32.3464
R1705 B.n938 B.n485 32.3464
R1706 B.n944 B.n485 32.3464
R1707 B.n950 B.n481 32.3464
R1708 B.n950 B.n477 32.3464
R1709 B.n956 B.n477 32.3464
R1710 B.n956 B.n473 32.3464
R1711 B.n962 B.n473 32.3464
R1712 B.n962 B.n469 32.3464
R1713 B.n968 B.n469 32.3464
R1714 B.n974 B.n465 32.3464
R1715 B.n974 B.n461 32.3464
R1716 B.n980 B.n461 32.3464
R1717 B.n980 B.n457 32.3464
R1718 B.n986 B.n457 32.3464
R1719 B.n986 B.n453 32.3464
R1720 B.n992 B.n453 32.3464
R1721 B.n998 B.n449 32.3464
R1722 B.n998 B.n445 32.3464
R1723 B.n1004 B.n445 32.3464
R1724 B.n1004 B.n441 32.3464
R1725 B.n1010 B.n441 32.3464
R1726 B.n1010 B.n437 32.3464
R1727 B.n1016 B.n437 32.3464
R1728 B.n1023 B.n433 32.3464
R1729 B.n1023 B.n429 32.3464
R1730 B.n1029 B.n429 32.3464
R1731 B.n1029 B.n4 32.3464
R1732 B.n1224 B.n4 32.3464
R1733 B.n1224 B.n1223 32.3464
R1734 B.n1223 B.n1222 32.3464
R1735 B.n1222 B.n8 32.3464
R1736 B.n12 B.n8 32.3464
R1737 B.n1215 B.n12 32.3464
R1738 B.n1215 B.n1214 32.3464
R1739 B.n1213 B.n16 32.3464
R1740 B.n1207 B.n16 32.3464
R1741 B.n1207 B.n1206 32.3464
R1742 B.n1206 B.n1205 32.3464
R1743 B.n1205 B.n23 32.3464
R1744 B.n1199 B.n23 32.3464
R1745 B.n1199 B.n1198 32.3464
R1746 B.n1197 B.n30 32.3464
R1747 B.n1191 B.n30 32.3464
R1748 B.n1191 B.n1190 32.3464
R1749 B.n1190 B.n1189 32.3464
R1750 B.n1189 B.n37 32.3464
R1751 B.n1183 B.n37 32.3464
R1752 B.n1183 B.n1182 32.3464
R1753 B.n1181 B.n44 32.3464
R1754 B.n1175 B.n44 32.3464
R1755 B.n1175 B.n1174 32.3464
R1756 B.n1174 B.n1173 32.3464
R1757 B.n1173 B.n51 32.3464
R1758 B.n1167 B.n51 32.3464
R1759 B.n1167 B.n1166 32.3464
R1760 B.n1165 B.n58 32.3464
R1761 B.n1159 B.n58 32.3464
R1762 B.n1159 B.n1158 32.3464
R1763 B.n1158 B.n1157 32.3464
R1764 B.n1157 B.n65 32.3464
R1765 B.n1151 B.n65 32.3464
R1766 B.n1151 B.n1150 32.3464
R1767 B.n1150 B.n1149 32.3464
R1768 B.n1143 B.n75 32.3464
R1769 B.n1143 B.n1142 32.3464
R1770 B.n1142 B.n1141 32.3464
R1771 B.n1141 B.n79 32.3464
R1772 B.n1135 B.n79 32.3464
R1773 B.n1135 B.n1134 32.3464
R1774 B.n1134 B.n1133 32.3464
R1775 B.n1133 B.n86 32.3464
R1776 B.n1127 B.n86 32.3464
R1777 B.n1127 B.n1126 32.3464
R1778 B.n1125 B.n93 32.3464
R1779 B.n1119 B.n93 32.3464
R1780 B.n1119 B.n1118 32.3464
R1781 B.n1118 B.n1117 32.3464
R1782 B.n1117 B.n100 32.3464
R1783 B.n1111 B.n100 32.3464
R1784 B.n1111 B.n1110 32.3464
R1785 B.n855 B.n534 32.0005
R1786 B.n862 B.n861 32.0005
R1787 B.n1107 B.n1106 32.0005
R1788 B.n176 B.n102 32.0005
R1789 B.n913 B.t6 31.3951
R1790 B.n75 B.t0 31.3951
R1791 B.t5 B.n481 26.6383
R1792 B.n1166 B.t3 26.6383
R1793 B.n1016 B.t9 25.687
R1794 B.t8 B.n1213 25.687
R1795 B.t7 B.n465 19.9789
R1796 B.n1182 B.t1 19.9789
R1797 B.n992 B.t2 19.0275
R1798 B.t4 B.n1197 19.0275
R1799 B.n883 B.t15 18.0762
R1800 B.t11 B.n1125 18.0762
R1801 B B.n1227 18.0485
R1802 B.t15 B.n520 14.2708
R1803 B.n1126 B.t11 14.2708
R1804 B.t2 B.n449 13.3194
R1805 B.n1198 B.t4 13.3194
R1806 B.n968 B.t7 12.3681
R1807 B.t1 B.n1181 12.3681
R1808 B.n867 B.n534 10.6151
R1809 B.n868 B.n867 10.6151
R1810 B.n869 B.n868 10.6151
R1811 B.n869 B.n526 10.6151
R1812 B.n879 B.n526 10.6151
R1813 B.n880 B.n879 10.6151
R1814 B.n881 B.n880 10.6151
R1815 B.n881 B.n518 10.6151
R1816 B.n891 B.n518 10.6151
R1817 B.n892 B.n891 10.6151
R1818 B.n893 B.n892 10.6151
R1819 B.n893 B.n510 10.6151
R1820 B.n903 B.n510 10.6151
R1821 B.n904 B.n903 10.6151
R1822 B.n905 B.n904 10.6151
R1823 B.n905 B.n502 10.6151
R1824 B.n916 B.n502 10.6151
R1825 B.n917 B.n916 10.6151
R1826 B.n918 B.n917 10.6151
R1827 B.n918 B.n495 10.6151
R1828 B.n928 B.n495 10.6151
R1829 B.n929 B.n928 10.6151
R1830 B.n930 B.n929 10.6151
R1831 B.n930 B.n487 10.6151
R1832 B.n940 B.n487 10.6151
R1833 B.n941 B.n940 10.6151
R1834 B.n942 B.n941 10.6151
R1835 B.n942 B.n479 10.6151
R1836 B.n952 B.n479 10.6151
R1837 B.n953 B.n952 10.6151
R1838 B.n954 B.n953 10.6151
R1839 B.n954 B.n471 10.6151
R1840 B.n964 B.n471 10.6151
R1841 B.n965 B.n964 10.6151
R1842 B.n966 B.n965 10.6151
R1843 B.n966 B.n463 10.6151
R1844 B.n976 B.n463 10.6151
R1845 B.n977 B.n976 10.6151
R1846 B.n978 B.n977 10.6151
R1847 B.n978 B.n455 10.6151
R1848 B.n988 B.n455 10.6151
R1849 B.n989 B.n988 10.6151
R1850 B.n990 B.n989 10.6151
R1851 B.n990 B.n447 10.6151
R1852 B.n1000 B.n447 10.6151
R1853 B.n1001 B.n1000 10.6151
R1854 B.n1002 B.n1001 10.6151
R1855 B.n1002 B.n439 10.6151
R1856 B.n1012 B.n439 10.6151
R1857 B.n1013 B.n1012 10.6151
R1858 B.n1014 B.n1013 10.6151
R1859 B.n1014 B.n431 10.6151
R1860 B.n1025 B.n431 10.6151
R1861 B.n1026 B.n1025 10.6151
R1862 B.n1027 B.n1026 10.6151
R1863 B.n1027 B.n0 10.6151
R1864 B.n855 B.n854 10.6151
R1865 B.n854 B.n853 10.6151
R1866 B.n853 B.n852 10.6151
R1867 B.n852 B.n850 10.6151
R1868 B.n850 B.n847 10.6151
R1869 B.n847 B.n846 10.6151
R1870 B.n846 B.n843 10.6151
R1871 B.n843 B.n842 10.6151
R1872 B.n842 B.n839 10.6151
R1873 B.n839 B.n838 10.6151
R1874 B.n838 B.n835 10.6151
R1875 B.n835 B.n834 10.6151
R1876 B.n834 B.n831 10.6151
R1877 B.n831 B.n830 10.6151
R1878 B.n830 B.n827 10.6151
R1879 B.n827 B.n826 10.6151
R1880 B.n826 B.n823 10.6151
R1881 B.n823 B.n822 10.6151
R1882 B.n822 B.n819 10.6151
R1883 B.n819 B.n818 10.6151
R1884 B.n818 B.n815 10.6151
R1885 B.n815 B.n814 10.6151
R1886 B.n814 B.n811 10.6151
R1887 B.n811 B.n810 10.6151
R1888 B.n810 B.n807 10.6151
R1889 B.n807 B.n806 10.6151
R1890 B.n806 B.n803 10.6151
R1891 B.n803 B.n802 10.6151
R1892 B.n802 B.n799 10.6151
R1893 B.n799 B.n798 10.6151
R1894 B.n798 B.n795 10.6151
R1895 B.n795 B.n794 10.6151
R1896 B.n794 B.n791 10.6151
R1897 B.n791 B.n790 10.6151
R1898 B.n790 B.n787 10.6151
R1899 B.n787 B.n786 10.6151
R1900 B.n786 B.n783 10.6151
R1901 B.n783 B.n782 10.6151
R1902 B.n782 B.n779 10.6151
R1903 B.n779 B.n778 10.6151
R1904 B.n778 B.n775 10.6151
R1905 B.n775 B.n774 10.6151
R1906 B.n774 B.n771 10.6151
R1907 B.n771 B.n770 10.6151
R1908 B.n770 B.n767 10.6151
R1909 B.n767 B.n766 10.6151
R1910 B.n766 B.n763 10.6151
R1911 B.n763 B.n762 10.6151
R1912 B.n762 B.n759 10.6151
R1913 B.n759 B.n758 10.6151
R1914 B.n758 B.n755 10.6151
R1915 B.n755 B.n754 10.6151
R1916 B.n754 B.n751 10.6151
R1917 B.n751 B.n750 10.6151
R1918 B.n750 B.n747 10.6151
R1919 B.n747 B.n746 10.6151
R1920 B.n746 B.n743 10.6151
R1921 B.n743 B.n742 10.6151
R1922 B.n739 B.n738 10.6151
R1923 B.n738 B.n735 10.6151
R1924 B.n735 B.n734 10.6151
R1925 B.n734 B.n731 10.6151
R1926 B.n731 B.n730 10.6151
R1927 B.n730 B.n727 10.6151
R1928 B.n727 B.n726 10.6151
R1929 B.n726 B.n723 10.6151
R1930 B.n721 B.n718 10.6151
R1931 B.n718 B.n717 10.6151
R1932 B.n717 B.n714 10.6151
R1933 B.n714 B.n713 10.6151
R1934 B.n713 B.n710 10.6151
R1935 B.n710 B.n709 10.6151
R1936 B.n709 B.n706 10.6151
R1937 B.n706 B.n705 10.6151
R1938 B.n705 B.n702 10.6151
R1939 B.n702 B.n701 10.6151
R1940 B.n701 B.n698 10.6151
R1941 B.n698 B.n697 10.6151
R1942 B.n697 B.n694 10.6151
R1943 B.n694 B.n693 10.6151
R1944 B.n693 B.n690 10.6151
R1945 B.n690 B.n689 10.6151
R1946 B.n689 B.n686 10.6151
R1947 B.n686 B.n685 10.6151
R1948 B.n685 B.n682 10.6151
R1949 B.n682 B.n681 10.6151
R1950 B.n681 B.n678 10.6151
R1951 B.n678 B.n677 10.6151
R1952 B.n677 B.n674 10.6151
R1953 B.n674 B.n673 10.6151
R1954 B.n673 B.n670 10.6151
R1955 B.n670 B.n669 10.6151
R1956 B.n669 B.n666 10.6151
R1957 B.n666 B.n665 10.6151
R1958 B.n665 B.n662 10.6151
R1959 B.n662 B.n661 10.6151
R1960 B.n661 B.n658 10.6151
R1961 B.n658 B.n657 10.6151
R1962 B.n657 B.n654 10.6151
R1963 B.n654 B.n653 10.6151
R1964 B.n653 B.n650 10.6151
R1965 B.n650 B.n649 10.6151
R1966 B.n649 B.n646 10.6151
R1967 B.n646 B.n645 10.6151
R1968 B.n645 B.n642 10.6151
R1969 B.n642 B.n641 10.6151
R1970 B.n641 B.n638 10.6151
R1971 B.n638 B.n637 10.6151
R1972 B.n637 B.n634 10.6151
R1973 B.n634 B.n633 10.6151
R1974 B.n633 B.n630 10.6151
R1975 B.n630 B.n629 10.6151
R1976 B.n629 B.n626 10.6151
R1977 B.n626 B.n625 10.6151
R1978 B.n625 B.n622 10.6151
R1979 B.n622 B.n621 10.6151
R1980 B.n621 B.n618 10.6151
R1981 B.n618 B.n617 10.6151
R1982 B.n617 B.n614 10.6151
R1983 B.n614 B.n613 10.6151
R1984 B.n613 B.n610 10.6151
R1985 B.n610 B.n609 10.6151
R1986 B.n609 B.n538 10.6151
R1987 B.n861 B.n538 10.6151
R1988 B.n863 B.n862 10.6151
R1989 B.n863 B.n530 10.6151
R1990 B.n873 B.n530 10.6151
R1991 B.n874 B.n873 10.6151
R1992 B.n875 B.n874 10.6151
R1993 B.n875 B.n522 10.6151
R1994 B.n885 B.n522 10.6151
R1995 B.n886 B.n885 10.6151
R1996 B.n887 B.n886 10.6151
R1997 B.n887 B.n514 10.6151
R1998 B.n897 B.n514 10.6151
R1999 B.n898 B.n897 10.6151
R2000 B.n899 B.n898 10.6151
R2001 B.n899 B.n506 10.6151
R2002 B.n909 B.n506 10.6151
R2003 B.n910 B.n909 10.6151
R2004 B.n911 B.n910 10.6151
R2005 B.n911 B.n499 10.6151
R2006 B.n922 B.n499 10.6151
R2007 B.n923 B.n922 10.6151
R2008 B.n924 B.n923 10.6151
R2009 B.n924 B.n491 10.6151
R2010 B.n934 B.n491 10.6151
R2011 B.n935 B.n934 10.6151
R2012 B.n936 B.n935 10.6151
R2013 B.n936 B.n483 10.6151
R2014 B.n946 B.n483 10.6151
R2015 B.n947 B.n946 10.6151
R2016 B.n948 B.n947 10.6151
R2017 B.n948 B.n475 10.6151
R2018 B.n958 B.n475 10.6151
R2019 B.n959 B.n958 10.6151
R2020 B.n960 B.n959 10.6151
R2021 B.n960 B.n467 10.6151
R2022 B.n970 B.n467 10.6151
R2023 B.n971 B.n970 10.6151
R2024 B.n972 B.n971 10.6151
R2025 B.n972 B.n459 10.6151
R2026 B.n982 B.n459 10.6151
R2027 B.n983 B.n982 10.6151
R2028 B.n984 B.n983 10.6151
R2029 B.n984 B.n451 10.6151
R2030 B.n994 B.n451 10.6151
R2031 B.n995 B.n994 10.6151
R2032 B.n996 B.n995 10.6151
R2033 B.n996 B.n443 10.6151
R2034 B.n1006 B.n443 10.6151
R2035 B.n1007 B.n1006 10.6151
R2036 B.n1008 B.n1007 10.6151
R2037 B.n1008 B.n435 10.6151
R2038 B.n1018 B.n435 10.6151
R2039 B.n1019 B.n1018 10.6151
R2040 B.n1021 B.n1019 10.6151
R2041 B.n1021 B.n1020 10.6151
R2042 B.n1020 B.n427 10.6151
R2043 B.n1032 B.n427 10.6151
R2044 B.n1033 B.n1032 10.6151
R2045 B.n1034 B.n1033 10.6151
R2046 B.n1035 B.n1034 10.6151
R2047 B.n1036 B.n1035 10.6151
R2048 B.n1039 B.n1036 10.6151
R2049 B.n1040 B.n1039 10.6151
R2050 B.n1041 B.n1040 10.6151
R2051 B.n1042 B.n1041 10.6151
R2052 B.n1044 B.n1042 10.6151
R2053 B.n1045 B.n1044 10.6151
R2054 B.n1046 B.n1045 10.6151
R2055 B.n1047 B.n1046 10.6151
R2056 B.n1049 B.n1047 10.6151
R2057 B.n1050 B.n1049 10.6151
R2058 B.n1051 B.n1050 10.6151
R2059 B.n1052 B.n1051 10.6151
R2060 B.n1054 B.n1052 10.6151
R2061 B.n1055 B.n1054 10.6151
R2062 B.n1056 B.n1055 10.6151
R2063 B.n1057 B.n1056 10.6151
R2064 B.n1059 B.n1057 10.6151
R2065 B.n1060 B.n1059 10.6151
R2066 B.n1061 B.n1060 10.6151
R2067 B.n1062 B.n1061 10.6151
R2068 B.n1064 B.n1062 10.6151
R2069 B.n1065 B.n1064 10.6151
R2070 B.n1066 B.n1065 10.6151
R2071 B.n1067 B.n1066 10.6151
R2072 B.n1069 B.n1067 10.6151
R2073 B.n1070 B.n1069 10.6151
R2074 B.n1071 B.n1070 10.6151
R2075 B.n1072 B.n1071 10.6151
R2076 B.n1074 B.n1072 10.6151
R2077 B.n1075 B.n1074 10.6151
R2078 B.n1076 B.n1075 10.6151
R2079 B.n1077 B.n1076 10.6151
R2080 B.n1079 B.n1077 10.6151
R2081 B.n1080 B.n1079 10.6151
R2082 B.n1081 B.n1080 10.6151
R2083 B.n1082 B.n1081 10.6151
R2084 B.n1084 B.n1082 10.6151
R2085 B.n1085 B.n1084 10.6151
R2086 B.n1086 B.n1085 10.6151
R2087 B.n1087 B.n1086 10.6151
R2088 B.n1089 B.n1087 10.6151
R2089 B.n1090 B.n1089 10.6151
R2090 B.n1091 B.n1090 10.6151
R2091 B.n1092 B.n1091 10.6151
R2092 B.n1094 B.n1092 10.6151
R2093 B.n1095 B.n1094 10.6151
R2094 B.n1096 B.n1095 10.6151
R2095 B.n1097 B.n1096 10.6151
R2096 B.n1099 B.n1097 10.6151
R2097 B.n1100 B.n1099 10.6151
R2098 B.n1101 B.n1100 10.6151
R2099 B.n1102 B.n1101 10.6151
R2100 B.n1104 B.n1102 10.6151
R2101 B.n1105 B.n1104 10.6151
R2102 B.n1106 B.n1105 10.6151
R2103 B.n1219 B.n1 10.6151
R2104 B.n1219 B.n1218 10.6151
R2105 B.n1218 B.n1217 10.6151
R2106 B.n1217 B.n10 10.6151
R2107 B.n1211 B.n10 10.6151
R2108 B.n1211 B.n1210 10.6151
R2109 B.n1210 B.n1209 10.6151
R2110 B.n1209 B.n18 10.6151
R2111 B.n1203 B.n18 10.6151
R2112 B.n1203 B.n1202 10.6151
R2113 B.n1202 B.n1201 10.6151
R2114 B.n1201 B.n25 10.6151
R2115 B.n1195 B.n25 10.6151
R2116 B.n1195 B.n1194 10.6151
R2117 B.n1194 B.n1193 10.6151
R2118 B.n1193 B.n32 10.6151
R2119 B.n1187 B.n32 10.6151
R2120 B.n1187 B.n1186 10.6151
R2121 B.n1186 B.n1185 10.6151
R2122 B.n1185 B.n39 10.6151
R2123 B.n1179 B.n39 10.6151
R2124 B.n1179 B.n1178 10.6151
R2125 B.n1178 B.n1177 10.6151
R2126 B.n1177 B.n46 10.6151
R2127 B.n1171 B.n46 10.6151
R2128 B.n1171 B.n1170 10.6151
R2129 B.n1170 B.n1169 10.6151
R2130 B.n1169 B.n53 10.6151
R2131 B.n1163 B.n53 10.6151
R2132 B.n1163 B.n1162 10.6151
R2133 B.n1162 B.n1161 10.6151
R2134 B.n1161 B.n60 10.6151
R2135 B.n1155 B.n60 10.6151
R2136 B.n1155 B.n1154 10.6151
R2137 B.n1154 B.n1153 10.6151
R2138 B.n1153 B.n67 10.6151
R2139 B.n1147 B.n67 10.6151
R2140 B.n1147 B.n1146 10.6151
R2141 B.n1146 B.n1145 10.6151
R2142 B.n1145 B.n73 10.6151
R2143 B.n1139 B.n73 10.6151
R2144 B.n1139 B.n1138 10.6151
R2145 B.n1138 B.n1137 10.6151
R2146 B.n1137 B.n81 10.6151
R2147 B.n1131 B.n81 10.6151
R2148 B.n1131 B.n1130 10.6151
R2149 B.n1130 B.n1129 10.6151
R2150 B.n1129 B.n88 10.6151
R2151 B.n1123 B.n88 10.6151
R2152 B.n1123 B.n1122 10.6151
R2153 B.n1122 B.n1121 10.6151
R2154 B.n1121 B.n95 10.6151
R2155 B.n1115 B.n95 10.6151
R2156 B.n1115 B.n1114 10.6151
R2157 B.n1114 B.n1113 10.6151
R2158 B.n1113 B.n102 10.6151
R2159 B.n177 B.n176 10.6151
R2160 B.n180 B.n177 10.6151
R2161 B.n181 B.n180 10.6151
R2162 B.n184 B.n181 10.6151
R2163 B.n185 B.n184 10.6151
R2164 B.n188 B.n185 10.6151
R2165 B.n189 B.n188 10.6151
R2166 B.n192 B.n189 10.6151
R2167 B.n193 B.n192 10.6151
R2168 B.n196 B.n193 10.6151
R2169 B.n197 B.n196 10.6151
R2170 B.n200 B.n197 10.6151
R2171 B.n201 B.n200 10.6151
R2172 B.n204 B.n201 10.6151
R2173 B.n205 B.n204 10.6151
R2174 B.n208 B.n205 10.6151
R2175 B.n209 B.n208 10.6151
R2176 B.n212 B.n209 10.6151
R2177 B.n213 B.n212 10.6151
R2178 B.n216 B.n213 10.6151
R2179 B.n217 B.n216 10.6151
R2180 B.n220 B.n217 10.6151
R2181 B.n221 B.n220 10.6151
R2182 B.n224 B.n221 10.6151
R2183 B.n225 B.n224 10.6151
R2184 B.n228 B.n225 10.6151
R2185 B.n229 B.n228 10.6151
R2186 B.n232 B.n229 10.6151
R2187 B.n233 B.n232 10.6151
R2188 B.n236 B.n233 10.6151
R2189 B.n237 B.n236 10.6151
R2190 B.n240 B.n237 10.6151
R2191 B.n241 B.n240 10.6151
R2192 B.n244 B.n241 10.6151
R2193 B.n245 B.n244 10.6151
R2194 B.n248 B.n245 10.6151
R2195 B.n249 B.n248 10.6151
R2196 B.n252 B.n249 10.6151
R2197 B.n253 B.n252 10.6151
R2198 B.n256 B.n253 10.6151
R2199 B.n257 B.n256 10.6151
R2200 B.n260 B.n257 10.6151
R2201 B.n261 B.n260 10.6151
R2202 B.n264 B.n261 10.6151
R2203 B.n265 B.n264 10.6151
R2204 B.n268 B.n265 10.6151
R2205 B.n269 B.n268 10.6151
R2206 B.n272 B.n269 10.6151
R2207 B.n273 B.n272 10.6151
R2208 B.n276 B.n273 10.6151
R2209 B.n277 B.n276 10.6151
R2210 B.n280 B.n277 10.6151
R2211 B.n281 B.n280 10.6151
R2212 B.n284 B.n281 10.6151
R2213 B.n285 B.n284 10.6151
R2214 B.n288 B.n285 10.6151
R2215 B.n289 B.n288 10.6151
R2216 B.n292 B.n289 10.6151
R2217 B.n297 B.n294 10.6151
R2218 B.n298 B.n297 10.6151
R2219 B.n301 B.n298 10.6151
R2220 B.n302 B.n301 10.6151
R2221 B.n305 B.n302 10.6151
R2222 B.n306 B.n305 10.6151
R2223 B.n309 B.n306 10.6151
R2224 B.n310 B.n309 10.6151
R2225 B.n314 B.n313 10.6151
R2226 B.n317 B.n314 10.6151
R2227 B.n318 B.n317 10.6151
R2228 B.n321 B.n318 10.6151
R2229 B.n322 B.n321 10.6151
R2230 B.n325 B.n322 10.6151
R2231 B.n326 B.n325 10.6151
R2232 B.n329 B.n326 10.6151
R2233 B.n330 B.n329 10.6151
R2234 B.n333 B.n330 10.6151
R2235 B.n334 B.n333 10.6151
R2236 B.n337 B.n334 10.6151
R2237 B.n338 B.n337 10.6151
R2238 B.n341 B.n338 10.6151
R2239 B.n342 B.n341 10.6151
R2240 B.n345 B.n342 10.6151
R2241 B.n346 B.n345 10.6151
R2242 B.n349 B.n346 10.6151
R2243 B.n350 B.n349 10.6151
R2244 B.n353 B.n350 10.6151
R2245 B.n354 B.n353 10.6151
R2246 B.n357 B.n354 10.6151
R2247 B.n358 B.n357 10.6151
R2248 B.n361 B.n358 10.6151
R2249 B.n362 B.n361 10.6151
R2250 B.n365 B.n362 10.6151
R2251 B.n366 B.n365 10.6151
R2252 B.n369 B.n366 10.6151
R2253 B.n370 B.n369 10.6151
R2254 B.n373 B.n370 10.6151
R2255 B.n374 B.n373 10.6151
R2256 B.n377 B.n374 10.6151
R2257 B.n378 B.n377 10.6151
R2258 B.n381 B.n378 10.6151
R2259 B.n382 B.n381 10.6151
R2260 B.n385 B.n382 10.6151
R2261 B.n386 B.n385 10.6151
R2262 B.n389 B.n386 10.6151
R2263 B.n390 B.n389 10.6151
R2264 B.n393 B.n390 10.6151
R2265 B.n394 B.n393 10.6151
R2266 B.n397 B.n394 10.6151
R2267 B.n398 B.n397 10.6151
R2268 B.n401 B.n398 10.6151
R2269 B.n402 B.n401 10.6151
R2270 B.n405 B.n402 10.6151
R2271 B.n406 B.n405 10.6151
R2272 B.n409 B.n406 10.6151
R2273 B.n410 B.n409 10.6151
R2274 B.n413 B.n410 10.6151
R2275 B.n414 B.n413 10.6151
R2276 B.n417 B.n414 10.6151
R2277 B.n418 B.n417 10.6151
R2278 B.n421 B.n418 10.6151
R2279 B.n422 B.n421 10.6151
R2280 B.n425 B.n422 10.6151
R2281 B.n426 B.n425 10.6151
R2282 B.n1107 B.n426 10.6151
R2283 B.n1227 B.n0 8.11757
R2284 B.n1227 B.n1 8.11757
R2285 B.t9 B.n433 6.65996
R2286 B.n1214 B.t8 6.65996
R2287 B.n739 B.n605 6.5566
R2288 B.n723 B.n722 6.5566
R2289 B.n294 B.n293 6.5566
R2290 B.n310 B.n172 6.5566
R2291 B.n944 B.t5 5.70861
R2292 B.t3 B.n1165 5.70861
R2293 B.n742 B.n605 4.05904
R2294 B.n722 B.n721 4.05904
R2295 B.n293 B.n292 4.05904
R2296 B.n313 B.n172 4.05904
R2297 B.n920 B.t6 0.951851
R2298 B.n1149 B.t0 0.951851
R2299 VN.n10 VN.t8 206.546
R2300 VN.n49 VN.t9 206.546
R2301 VN.n19 VN.t7 174.873
R2302 VN.n9 VN.t3 174.873
R2303 VN.n3 VN.t4 174.873
R2304 VN.n37 VN.t1 174.873
R2305 VN.n58 VN.t2 174.873
R2306 VN.n48 VN.t6 174.873
R2307 VN.n42 VN.t0 174.873
R2308 VN.n76 VN.t5 174.873
R2309 VN.n75 VN.n39 161.3
R2310 VN.n74 VN.n73 161.3
R2311 VN.n72 VN.n40 161.3
R2312 VN.n71 VN.n70 161.3
R2313 VN.n69 VN.n41 161.3
R2314 VN.n68 VN.n67 161.3
R2315 VN.n66 VN.n65 161.3
R2316 VN.n64 VN.n43 161.3
R2317 VN.n63 VN.n62 161.3
R2318 VN.n61 VN.n44 161.3
R2319 VN.n60 VN.n59 161.3
R2320 VN.n58 VN.n45 161.3
R2321 VN.n57 VN.n56 161.3
R2322 VN.n55 VN.n46 161.3
R2323 VN.n54 VN.n53 161.3
R2324 VN.n52 VN.n47 161.3
R2325 VN.n51 VN.n50 161.3
R2326 VN.n36 VN.n0 161.3
R2327 VN.n35 VN.n34 161.3
R2328 VN.n33 VN.n1 161.3
R2329 VN.n32 VN.n31 161.3
R2330 VN.n30 VN.n2 161.3
R2331 VN.n29 VN.n28 161.3
R2332 VN.n27 VN.n26 161.3
R2333 VN.n25 VN.n4 161.3
R2334 VN.n24 VN.n23 161.3
R2335 VN.n22 VN.n5 161.3
R2336 VN.n21 VN.n20 161.3
R2337 VN.n19 VN.n6 161.3
R2338 VN.n18 VN.n17 161.3
R2339 VN.n16 VN.n7 161.3
R2340 VN.n15 VN.n14 161.3
R2341 VN.n13 VN.n8 161.3
R2342 VN.n12 VN.n11 161.3
R2343 VN.n38 VN.n37 106.841
R2344 VN.n77 VN.n76 106.841
R2345 VN.n10 VN.n9 57.8794
R2346 VN.n49 VN.n48 57.8794
R2347 VN VN.n77 56.9565
R2348 VN.n31 VN.n1 56.5193
R2349 VN.n70 VN.n40 56.5193
R2350 VN.n14 VN.n7 50.6917
R2351 VN.n24 VN.n5 50.6917
R2352 VN.n53 VN.n46 50.6917
R2353 VN.n63 VN.n44 50.6917
R2354 VN.n14 VN.n13 30.2951
R2355 VN.n25 VN.n24 30.2951
R2356 VN.n53 VN.n52 30.2951
R2357 VN.n64 VN.n63 30.2951
R2358 VN.n13 VN.n12 24.4675
R2359 VN.n18 VN.n7 24.4675
R2360 VN.n19 VN.n18 24.4675
R2361 VN.n20 VN.n19 24.4675
R2362 VN.n20 VN.n5 24.4675
R2363 VN.n26 VN.n25 24.4675
R2364 VN.n30 VN.n29 24.4675
R2365 VN.n31 VN.n30 24.4675
R2366 VN.n35 VN.n1 24.4675
R2367 VN.n36 VN.n35 24.4675
R2368 VN.n52 VN.n51 24.4675
R2369 VN.n59 VN.n44 24.4675
R2370 VN.n59 VN.n58 24.4675
R2371 VN.n58 VN.n57 24.4675
R2372 VN.n57 VN.n46 24.4675
R2373 VN.n70 VN.n69 24.4675
R2374 VN.n69 VN.n68 24.4675
R2375 VN.n65 VN.n64 24.4675
R2376 VN.n75 VN.n74 24.4675
R2377 VN.n74 VN.n40 24.4675
R2378 VN.n12 VN.n9 14.1914
R2379 VN.n26 VN.n3 14.1914
R2380 VN.n51 VN.n48 14.1914
R2381 VN.n65 VN.n42 14.1914
R2382 VN.n29 VN.n3 10.2766
R2383 VN.n68 VN.n42 10.2766
R2384 VN.n50 VN.n49 7.2327
R2385 VN.n11 VN.n10 7.2327
R2386 VN.n37 VN.n36 3.91522
R2387 VN.n76 VN.n75 3.91522
R2388 VN.n77 VN.n39 0.278367
R2389 VN.n38 VN.n0 0.278367
R2390 VN.n73 VN.n39 0.189894
R2391 VN.n73 VN.n72 0.189894
R2392 VN.n72 VN.n71 0.189894
R2393 VN.n71 VN.n41 0.189894
R2394 VN.n67 VN.n41 0.189894
R2395 VN.n67 VN.n66 0.189894
R2396 VN.n66 VN.n43 0.189894
R2397 VN.n62 VN.n43 0.189894
R2398 VN.n62 VN.n61 0.189894
R2399 VN.n61 VN.n60 0.189894
R2400 VN.n60 VN.n45 0.189894
R2401 VN.n56 VN.n45 0.189894
R2402 VN.n56 VN.n55 0.189894
R2403 VN.n55 VN.n54 0.189894
R2404 VN.n54 VN.n47 0.189894
R2405 VN.n50 VN.n47 0.189894
R2406 VN.n11 VN.n8 0.189894
R2407 VN.n15 VN.n8 0.189894
R2408 VN.n16 VN.n15 0.189894
R2409 VN.n17 VN.n16 0.189894
R2410 VN.n17 VN.n6 0.189894
R2411 VN.n21 VN.n6 0.189894
R2412 VN.n22 VN.n21 0.189894
R2413 VN.n23 VN.n22 0.189894
R2414 VN.n23 VN.n4 0.189894
R2415 VN.n27 VN.n4 0.189894
R2416 VN.n28 VN.n27 0.189894
R2417 VN.n28 VN.n2 0.189894
R2418 VN.n32 VN.n2 0.189894
R2419 VN.n33 VN.n32 0.189894
R2420 VN.n34 VN.n33 0.189894
R2421 VN.n34 VN.n0 0.189894
R2422 VN VN.n38 0.153454
R2423 VDD2.n1 VDD2.t1 63.5964
R2424 VDD2.n3 VDD2.n2 61.8305
R2425 VDD2 VDD2.n7 61.8277
R2426 VDD2.n4 VDD2.t4 61.1914
R2427 VDD2.n6 VDD2.n5 60.0822
R2428 VDD2.n1 VDD2.n0 60.0819
R2429 VDD2.n4 VDD2.n3 50.5278
R2430 VDD2.n6 VDD2.n4 2.40567
R2431 VDD2.n7 VDD2.t3 1.10974
R2432 VDD2.n7 VDD2.t0 1.10974
R2433 VDD2.n5 VDD2.t9 1.10974
R2434 VDD2.n5 VDD2.t7 1.10974
R2435 VDD2.n2 VDD2.t5 1.10974
R2436 VDD2.n2 VDD2.t8 1.10974
R2437 VDD2.n0 VDD2.t6 1.10974
R2438 VDD2.n0 VDD2.t2 1.10974
R2439 VDD2 VDD2.n6 0.659983
R2440 VDD2.n3 VDD2.n1 0.546447
C0 VP VN 9.28051f
C1 VTAIL VP 15.778199f
C2 VDD2 VP 0.566252f
C3 VTAIL VN 15.7638f
C4 VDD2 VN 15.4394f
C5 VDD1 VP 15.8477f
C6 VDD2 VTAIL 13.1946f
C7 VDD1 VN 0.153082f
C8 VTAIL VDD1 13.1462f
C9 VDD2 VDD1 2.08431f
C10 VDD2 B 8.082314f
C11 VDD1 B 8.055098f
C12 VTAIL B 10.420218f
C13 VN B 17.98317f
C14 VP B 16.397028f
C15 VDD2.t1 B 3.86458f
C16 VDD2.t6 B 0.330686f
C17 VDD2.t2 B 0.330686f
C18 VDD2.n0 B 3.01055f
C19 VDD2.n1 B 0.854164f
C20 VDD2.t5 B 0.330686f
C21 VDD2.t8 B 0.330686f
C22 VDD2.n2 B 3.02524f
C23 VDD2.n3 B 3.00111f
C24 VDD2.t4 B 3.8475f
C25 VDD2.n4 B 3.30279f
C26 VDD2.t9 B 0.330686f
C27 VDD2.t7 B 0.330686f
C28 VDD2.n5 B 3.01056f
C29 VDD2.n6 B 0.427134f
C30 VDD2.t3 B 0.330686f
C31 VDD2.t0 B 0.330686f
C32 VDD2.n7 B 3.02519f
C33 VN.n0 B 0.028148f
C34 VN.t1 B 2.57825f
C35 VN.n1 B 0.035036f
C36 VN.n2 B 0.02135f
C37 VN.t4 B 2.57825f
C38 VN.n3 B 0.895417f
C39 VN.n4 B 0.02135f
C40 VN.n5 B 0.038978f
C41 VN.n6 B 0.02135f
C42 VN.t7 B 2.57825f
C43 VN.n7 B 0.038978f
C44 VN.n8 B 0.02135f
C45 VN.t3 B 2.57825f
C46 VN.n9 B 0.956542f
C47 VN.t8 B 2.73478f
C48 VN.n10 B 0.94355f
C49 VN.n11 B 0.202707f
C50 VN.n12 B 0.03154f
C51 VN.n13 B 0.042663f
C52 VN.n14 B 0.020488f
C53 VN.n15 B 0.02135f
C54 VN.n16 B 0.02135f
C55 VN.n17 B 0.02135f
C56 VN.n18 B 0.039791f
C57 VN.n19 B 0.915563f
C58 VN.n20 B 0.039791f
C59 VN.n21 B 0.02135f
C60 VN.n22 B 0.02135f
C61 VN.n23 B 0.02135f
C62 VN.n24 B 0.020488f
C63 VN.n25 B 0.042663f
C64 VN.n26 B 0.03154f
C65 VN.n27 B 0.02135f
C66 VN.n28 B 0.02135f
C67 VN.n29 B 0.028397f
C68 VN.n30 B 0.039791f
C69 VN.n31 B 0.027302f
C70 VN.n32 B 0.02135f
C71 VN.n33 B 0.02135f
C72 VN.n34 B 0.02135f
C73 VN.n35 B 0.039791f
C74 VN.n36 B 0.023289f
C75 VN.n37 B 0.956225f
C76 VN.n38 B 0.036527f
C77 VN.n39 B 0.028148f
C78 VN.t5 B 2.57825f
C79 VN.n40 B 0.035036f
C80 VN.n41 B 0.02135f
C81 VN.t0 B 2.57825f
C82 VN.n42 B 0.895417f
C83 VN.n43 B 0.02135f
C84 VN.n44 B 0.038978f
C85 VN.n45 B 0.02135f
C86 VN.t2 B 2.57825f
C87 VN.n46 B 0.038978f
C88 VN.n47 B 0.02135f
C89 VN.t6 B 2.57825f
C90 VN.n48 B 0.956542f
C91 VN.t9 B 2.73478f
C92 VN.n49 B 0.94355f
C93 VN.n50 B 0.202707f
C94 VN.n51 B 0.03154f
C95 VN.n52 B 0.042663f
C96 VN.n53 B 0.020488f
C97 VN.n54 B 0.02135f
C98 VN.n55 B 0.02135f
C99 VN.n56 B 0.02135f
C100 VN.n57 B 0.039791f
C101 VN.n58 B 0.915563f
C102 VN.n59 B 0.039791f
C103 VN.n60 B 0.02135f
C104 VN.n61 B 0.02135f
C105 VN.n62 B 0.02135f
C106 VN.n63 B 0.020488f
C107 VN.n64 B 0.042663f
C108 VN.n65 B 0.03154f
C109 VN.n66 B 0.02135f
C110 VN.n67 B 0.02135f
C111 VN.n68 B 0.028397f
C112 VN.n69 B 0.039791f
C113 VN.n70 B 0.027302f
C114 VN.n71 B 0.02135f
C115 VN.n72 B 0.02135f
C116 VN.n73 B 0.02135f
C117 VN.n74 B 0.039791f
C118 VN.n75 B 0.023289f
C119 VN.n76 B 0.956225f
C120 VN.n77 B 1.43277f
C121 VDD1.t3 B 3.89137f
C122 VDD1.t7 B 0.332979f
C123 VDD1.t9 B 0.332979f
C124 VDD1.n0 B 3.03143f
C125 VDD1.n1 B 0.867713f
C126 VDD1.t4 B 3.89137f
C127 VDD1.t0 B 0.332979f
C128 VDD1.t1 B 0.332979f
C129 VDD1.n2 B 3.03142f
C130 VDD1.n3 B 0.860085f
C131 VDD1.t6 B 0.332979f
C132 VDD1.t8 B 0.332979f
C133 VDD1.n4 B 3.04621f
C134 VDD1.n5 B 3.13968f
C135 VDD1.t2 B 0.332979f
C136 VDD1.t5 B 0.332979f
C137 VDD1.n6 B 3.03142f
C138 VDD1.n7 B 3.36253f
C139 VTAIL.t8 B 0.333472f
C140 VTAIL.t4 B 0.333472f
C141 VTAIL.n0 B 2.96184f
C142 VTAIL.n1 B 0.508474f
C143 VTAIL.t19 B 3.78314f
C144 VTAIL.n2 B 0.638009f
C145 VTAIL.t13 B 0.333472f
C146 VTAIL.t15 B 0.333472f
C147 VTAIL.n3 B 2.96184f
C148 VTAIL.n4 B 0.605665f
C149 VTAIL.t17 B 0.333472f
C150 VTAIL.t12 B 0.333472f
C151 VTAIL.n5 B 2.96184f
C152 VTAIL.n6 B 2.28223f
C153 VTAIL.t6 B 0.333472f
C154 VTAIL.t5 B 0.333472f
C155 VTAIL.n7 B 2.96184f
C156 VTAIL.n8 B 2.28222f
C157 VTAIL.t7 B 0.333472f
C158 VTAIL.t2 B 0.333472f
C159 VTAIL.n9 B 2.96184f
C160 VTAIL.n10 B 0.605661f
C161 VTAIL.t9 B 3.78315f
C162 VTAIL.n11 B 0.638005f
C163 VTAIL.t14 B 0.333472f
C164 VTAIL.t18 B 0.333472f
C165 VTAIL.n12 B 2.96184f
C166 VTAIL.n13 B 0.549842f
C167 VTAIL.t16 B 0.333472f
C168 VTAIL.t10 B 0.333472f
C169 VTAIL.n14 B 2.96184f
C170 VTAIL.n15 B 0.605661f
C171 VTAIL.t11 B 3.78314f
C172 VTAIL.n16 B 2.18717f
C173 VTAIL.t0 B 3.78314f
C174 VTAIL.n17 B 2.18717f
C175 VTAIL.t1 B 0.333472f
C176 VTAIL.t3 B 0.333472f
C177 VTAIL.n18 B 2.96184f
C178 VTAIL.n19 B 0.463818f
C179 VP.n0 B 0.028447f
C180 VP.t1 B 2.60565f
C181 VP.n1 B 0.035409f
C182 VP.n2 B 0.021577f
C183 VP.t3 B 2.60565f
C184 VP.n3 B 0.904931f
C185 VP.n4 B 0.021577f
C186 VP.n5 B 0.039392f
C187 VP.n6 B 0.021577f
C188 VP.t8 B 2.60565f
C189 VP.n7 B 0.039392f
C190 VP.n8 B 0.021577f
C191 VP.t9 B 2.60565f
C192 VP.n9 B 0.904931f
C193 VP.n10 B 0.021577f
C194 VP.n11 B 0.035409f
C195 VP.n12 B 0.028447f
C196 VP.t5 B 2.60565f
C197 VP.n13 B 0.028447f
C198 VP.t4 B 2.60565f
C199 VP.n14 B 0.035409f
C200 VP.n15 B 0.021577f
C201 VP.t7 B 2.60565f
C202 VP.n16 B 0.904931f
C203 VP.n17 B 0.021577f
C204 VP.n18 B 0.039392f
C205 VP.n19 B 0.021577f
C206 VP.t0 B 2.60565f
C207 VP.n20 B 0.039392f
C208 VP.n21 B 0.021577f
C209 VP.t2 B 2.60565f
C210 VP.n22 B 0.966706f
C211 VP.t6 B 2.76383f
C212 VP.n23 B 0.953576f
C213 VP.n24 B 0.204861f
C214 VP.n25 B 0.031875f
C215 VP.n26 B 0.043116f
C216 VP.n27 B 0.020706f
C217 VP.n28 B 0.021577f
C218 VP.n29 B 0.021577f
C219 VP.n30 B 0.021577f
C220 VP.n31 B 0.040214f
C221 VP.n32 B 0.925291f
C222 VP.n33 B 0.040214f
C223 VP.n34 B 0.021577f
C224 VP.n35 B 0.021577f
C225 VP.n36 B 0.021577f
C226 VP.n37 B 0.020706f
C227 VP.n38 B 0.043116f
C228 VP.n39 B 0.031875f
C229 VP.n40 B 0.021577f
C230 VP.n41 B 0.021577f
C231 VP.n42 B 0.028699f
C232 VP.n43 B 0.040214f
C233 VP.n44 B 0.027592f
C234 VP.n45 B 0.021577f
C235 VP.n46 B 0.021577f
C236 VP.n47 B 0.021577f
C237 VP.n48 B 0.040214f
C238 VP.n49 B 0.023537f
C239 VP.n50 B 0.966386f
C240 VP.n51 B 1.43661f
C241 VP.n52 B 1.4503f
C242 VP.n53 B 0.966386f
C243 VP.n54 B 0.023537f
C244 VP.n55 B 0.040214f
C245 VP.n56 B 0.021577f
C246 VP.n57 B 0.021577f
C247 VP.n58 B 0.021577f
C248 VP.n59 B 0.027592f
C249 VP.n60 B 0.040214f
C250 VP.n61 B 0.028699f
C251 VP.n62 B 0.021577f
C252 VP.n63 B 0.021577f
C253 VP.n64 B 0.031875f
C254 VP.n65 B 0.043116f
C255 VP.n66 B 0.020706f
C256 VP.n67 B 0.021577f
C257 VP.n68 B 0.021577f
C258 VP.n69 B 0.021577f
C259 VP.n70 B 0.040214f
C260 VP.n71 B 0.925291f
C261 VP.n72 B 0.040214f
C262 VP.n73 B 0.021577f
C263 VP.n74 B 0.021577f
C264 VP.n75 B 0.021577f
C265 VP.n76 B 0.020706f
C266 VP.n77 B 0.043116f
C267 VP.n78 B 0.031875f
C268 VP.n79 B 0.021577f
C269 VP.n80 B 0.021577f
C270 VP.n81 B 0.028699f
C271 VP.n82 B 0.040214f
C272 VP.n83 B 0.027592f
C273 VP.n84 B 0.021577f
C274 VP.n85 B 0.021577f
C275 VP.n86 B 0.021577f
C276 VP.n87 B 0.040214f
C277 VP.n88 B 0.023537f
C278 VP.n89 B 0.966386f
C279 VP.n90 B 0.036915f
.ends

