* NGSPICE file created from diff_pair_sample_1714.ext - technology: sky130A

.subckt diff_pair_sample_1714 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n1794_n3680# sky130_fd_pr__pfet_01v8 ad=5.2884 pd=27.9 as=0 ps=0 w=13.56 l=1.73
X1 VDD2.t1 VN.t0 VTAIL.t3 w_n1794_n3680# sky130_fd_pr__pfet_01v8 ad=5.2884 pd=27.9 as=5.2884 ps=27.9 w=13.56 l=1.73
X2 B.t8 B.t6 B.t7 w_n1794_n3680# sky130_fd_pr__pfet_01v8 ad=5.2884 pd=27.9 as=0 ps=0 w=13.56 l=1.73
X3 VDD2.t0 VN.t1 VTAIL.t2 w_n1794_n3680# sky130_fd_pr__pfet_01v8 ad=5.2884 pd=27.9 as=5.2884 ps=27.9 w=13.56 l=1.73
X4 VDD1.t1 VP.t0 VTAIL.t0 w_n1794_n3680# sky130_fd_pr__pfet_01v8 ad=5.2884 pd=27.9 as=5.2884 ps=27.9 w=13.56 l=1.73
X5 B.t5 B.t3 B.t4 w_n1794_n3680# sky130_fd_pr__pfet_01v8 ad=5.2884 pd=27.9 as=0 ps=0 w=13.56 l=1.73
X6 B.t2 B.t0 B.t1 w_n1794_n3680# sky130_fd_pr__pfet_01v8 ad=5.2884 pd=27.9 as=0 ps=0 w=13.56 l=1.73
X7 VDD1.t0 VP.t1 VTAIL.t1 w_n1794_n3680# sky130_fd_pr__pfet_01v8 ad=5.2884 pd=27.9 as=5.2884 ps=27.9 w=13.56 l=1.73
R0 B.n398 B.n67 585
R1 B.n400 B.n399 585
R2 B.n401 B.n66 585
R3 B.n403 B.n402 585
R4 B.n404 B.n65 585
R5 B.n406 B.n405 585
R6 B.n407 B.n64 585
R7 B.n409 B.n408 585
R8 B.n410 B.n63 585
R9 B.n412 B.n411 585
R10 B.n413 B.n62 585
R11 B.n415 B.n414 585
R12 B.n416 B.n61 585
R13 B.n418 B.n417 585
R14 B.n419 B.n60 585
R15 B.n421 B.n420 585
R16 B.n422 B.n59 585
R17 B.n424 B.n423 585
R18 B.n425 B.n58 585
R19 B.n427 B.n426 585
R20 B.n428 B.n57 585
R21 B.n430 B.n429 585
R22 B.n431 B.n56 585
R23 B.n433 B.n432 585
R24 B.n434 B.n55 585
R25 B.n436 B.n435 585
R26 B.n437 B.n54 585
R27 B.n439 B.n438 585
R28 B.n440 B.n53 585
R29 B.n442 B.n441 585
R30 B.n443 B.n52 585
R31 B.n445 B.n444 585
R32 B.n446 B.n51 585
R33 B.n448 B.n447 585
R34 B.n449 B.n50 585
R35 B.n451 B.n450 585
R36 B.n452 B.n49 585
R37 B.n454 B.n453 585
R38 B.n455 B.n48 585
R39 B.n457 B.n456 585
R40 B.n458 B.n47 585
R41 B.n460 B.n459 585
R42 B.n461 B.n46 585
R43 B.n463 B.n462 585
R44 B.n464 B.n45 585
R45 B.n466 B.n465 585
R46 B.n468 B.n467 585
R47 B.n469 B.n41 585
R48 B.n471 B.n470 585
R49 B.n472 B.n40 585
R50 B.n474 B.n473 585
R51 B.n475 B.n39 585
R52 B.n477 B.n476 585
R53 B.n478 B.n38 585
R54 B.n480 B.n479 585
R55 B.n481 B.n35 585
R56 B.n484 B.n483 585
R57 B.n485 B.n34 585
R58 B.n487 B.n486 585
R59 B.n488 B.n33 585
R60 B.n490 B.n489 585
R61 B.n491 B.n32 585
R62 B.n493 B.n492 585
R63 B.n494 B.n31 585
R64 B.n496 B.n495 585
R65 B.n497 B.n30 585
R66 B.n499 B.n498 585
R67 B.n500 B.n29 585
R68 B.n502 B.n501 585
R69 B.n503 B.n28 585
R70 B.n505 B.n504 585
R71 B.n506 B.n27 585
R72 B.n508 B.n507 585
R73 B.n509 B.n26 585
R74 B.n511 B.n510 585
R75 B.n512 B.n25 585
R76 B.n514 B.n513 585
R77 B.n515 B.n24 585
R78 B.n517 B.n516 585
R79 B.n518 B.n23 585
R80 B.n520 B.n519 585
R81 B.n521 B.n22 585
R82 B.n523 B.n522 585
R83 B.n524 B.n21 585
R84 B.n526 B.n525 585
R85 B.n527 B.n20 585
R86 B.n529 B.n528 585
R87 B.n530 B.n19 585
R88 B.n532 B.n531 585
R89 B.n533 B.n18 585
R90 B.n535 B.n534 585
R91 B.n536 B.n17 585
R92 B.n538 B.n537 585
R93 B.n539 B.n16 585
R94 B.n541 B.n540 585
R95 B.n542 B.n15 585
R96 B.n544 B.n543 585
R97 B.n545 B.n14 585
R98 B.n547 B.n546 585
R99 B.n548 B.n13 585
R100 B.n550 B.n549 585
R101 B.n551 B.n12 585
R102 B.n397 B.n396 585
R103 B.n395 B.n68 585
R104 B.n394 B.n393 585
R105 B.n392 B.n69 585
R106 B.n391 B.n390 585
R107 B.n389 B.n70 585
R108 B.n388 B.n387 585
R109 B.n386 B.n71 585
R110 B.n385 B.n384 585
R111 B.n383 B.n72 585
R112 B.n382 B.n381 585
R113 B.n380 B.n73 585
R114 B.n379 B.n378 585
R115 B.n377 B.n74 585
R116 B.n376 B.n375 585
R117 B.n374 B.n75 585
R118 B.n373 B.n372 585
R119 B.n371 B.n76 585
R120 B.n370 B.n369 585
R121 B.n368 B.n77 585
R122 B.n367 B.n366 585
R123 B.n365 B.n78 585
R124 B.n364 B.n363 585
R125 B.n362 B.n79 585
R126 B.n361 B.n360 585
R127 B.n359 B.n80 585
R128 B.n358 B.n357 585
R129 B.n356 B.n81 585
R130 B.n355 B.n354 585
R131 B.n353 B.n82 585
R132 B.n352 B.n351 585
R133 B.n350 B.n83 585
R134 B.n349 B.n348 585
R135 B.n347 B.n84 585
R136 B.n346 B.n345 585
R137 B.n344 B.n85 585
R138 B.n343 B.n342 585
R139 B.n341 B.n86 585
R140 B.n340 B.n339 585
R141 B.n338 B.n87 585
R142 B.n337 B.n336 585
R143 B.n182 B.n143 585
R144 B.n184 B.n183 585
R145 B.n185 B.n142 585
R146 B.n187 B.n186 585
R147 B.n188 B.n141 585
R148 B.n190 B.n189 585
R149 B.n191 B.n140 585
R150 B.n193 B.n192 585
R151 B.n194 B.n139 585
R152 B.n196 B.n195 585
R153 B.n197 B.n138 585
R154 B.n199 B.n198 585
R155 B.n200 B.n137 585
R156 B.n202 B.n201 585
R157 B.n203 B.n136 585
R158 B.n205 B.n204 585
R159 B.n206 B.n135 585
R160 B.n208 B.n207 585
R161 B.n209 B.n134 585
R162 B.n211 B.n210 585
R163 B.n212 B.n133 585
R164 B.n214 B.n213 585
R165 B.n215 B.n132 585
R166 B.n217 B.n216 585
R167 B.n218 B.n131 585
R168 B.n220 B.n219 585
R169 B.n221 B.n130 585
R170 B.n223 B.n222 585
R171 B.n224 B.n129 585
R172 B.n226 B.n225 585
R173 B.n227 B.n128 585
R174 B.n229 B.n228 585
R175 B.n230 B.n127 585
R176 B.n232 B.n231 585
R177 B.n233 B.n126 585
R178 B.n235 B.n234 585
R179 B.n236 B.n125 585
R180 B.n238 B.n237 585
R181 B.n239 B.n124 585
R182 B.n241 B.n240 585
R183 B.n242 B.n123 585
R184 B.n244 B.n243 585
R185 B.n245 B.n122 585
R186 B.n247 B.n246 585
R187 B.n248 B.n121 585
R188 B.n250 B.n249 585
R189 B.n252 B.n251 585
R190 B.n253 B.n117 585
R191 B.n255 B.n254 585
R192 B.n256 B.n116 585
R193 B.n258 B.n257 585
R194 B.n259 B.n115 585
R195 B.n261 B.n260 585
R196 B.n262 B.n114 585
R197 B.n264 B.n263 585
R198 B.n265 B.n111 585
R199 B.n268 B.n267 585
R200 B.n269 B.n110 585
R201 B.n271 B.n270 585
R202 B.n272 B.n109 585
R203 B.n274 B.n273 585
R204 B.n275 B.n108 585
R205 B.n277 B.n276 585
R206 B.n278 B.n107 585
R207 B.n280 B.n279 585
R208 B.n281 B.n106 585
R209 B.n283 B.n282 585
R210 B.n284 B.n105 585
R211 B.n286 B.n285 585
R212 B.n287 B.n104 585
R213 B.n289 B.n288 585
R214 B.n290 B.n103 585
R215 B.n292 B.n291 585
R216 B.n293 B.n102 585
R217 B.n295 B.n294 585
R218 B.n296 B.n101 585
R219 B.n298 B.n297 585
R220 B.n299 B.n100 585
R221 B.n301 B.n300 585
R222 B.n302 B.n99 585
R223 B.n304 B.n303 585
R224 B.n305 B.n98 585
R225 B.n307 B.n306 585
R226 B.n308 B.n97 585
R227 B.n310 B.n309 585
R228 B.n311 B.n96 585
R229 B.n313 B.n312 585
R230 B.n314 B.n95 585
R231 B.n316 B.n315 585
R232 B.n317 B.n94 585
R233 B.n319 B.n318 585
R234 B.n320 B.n93 585
R235 B.n322 B.n321 585
R236 B.n323 B.n92 585
R237 B.n325 B.n324 585
R238 B.n326 B.n91 585
R239 B.n328 B.n327 585
R240 B.n329 B.n90 585
R241 B.n331 B.n330 585
R242 B.n332 B.n89 585
R243 B.n334 B.n333 585
R244 B.n335 B.n88 585
R245 B.n181 B.n180 585
R246 B.n179 B.n144 585
R247 B.n178 B.n177 585
R248 B.n176 B.n145 585
R249 B.n175 B.n174 585
R250 B.n173 B.n146 585
R251 B.n172 B.n171 585
R252 B.n170 B.n147 585
R253 B.n169 B.n168 585
R254 B.n167 B.n148 585
R255 B.n166 B.n165 585
R256 B.n164 B.n149 585
R257 B.n163 B.n162 585
R258 B.n161 B.n150 585
R259 B.n160 B.n159 585
R260 B.n158 B.n151 585
R261 B.n157 B.n156 585
R262 B.n155 B.n152 585
R263 B.n154 B.n153 585
R264 B.n2 B.n0 585
R265 B.n581 B.n1 585
R266 B.n580 B.n579 585
R267 B.n578 B.n3 585
R268 B.n577 B.n576 585
R269 B.n575 B.n4 585
R270 B.n574 B.n573 585
R271 B.n572 B.n5 585
R272 B.n571 B.n570 585
R273 B.n569 B.n6 585
R274 B.n568 B.n567 585
R275 B.n566 B.n7 585
R276 B.n565 B.n564 585
R277 B.n563 B.n8 585
R278 B.n562 B.n561 585
R279 B.n560 B.n9 585
R280 B.n559 B.n558 585
R281 B.n557 B.n10 585
R282 B.n556 B.n555 585
R283 B.n554 B.n11 585
R284 B.n553 B.n552 585
R285 B.n583 B.n582 585
R286 B.n180 B.n143 535.745
R287 B.n552 B.n551 535.745
R288 B.n336 B.n335 535.745
R289 B.n396 B.n67 535.745
R290 B.n112 B.t5 443.854
R291 B.n42 B.t7 443.854
R292 B.n118 B.t2 443.854
R293 B.n36 B.t10 443.854
R294 B.n113 B.t4 403.904
R295 B.n43 B.t8 403.904
R296 B.n119 B.t1 403.902
R297 B.n37 B.t11 403.902
R298 B.n112 B.t3 395.104
R299 B.n118 B.t0 395.104
R300 B.n36 B.t9 395.104
R301 B.n42 B.t6 395.104
R302 B.n180 B.n179 163.367
R303 B.n179 B.n178 163.367
R304 B.n178 B.n145 163.367
R305 B.n174 B.n145 163.367
R306 B.n174 B.n173 163.367
R307 B.n173 B.n172 163.367
R308 B.n172 B.n147 163.367
R309 B.n168 B.n147 163.367
R310 B.n168 B.n167 163.367
R311 B.n167 B.n166 163.367
R312 B.n166 B.n149 163.367
R313 B.n162 B.n149 163.367
R314 B.n162 B.n161 163.367
R315 B.n161 B.n160 163.367
R316 B.n160 B.n151 163.367
R317 B.n156 B.n151 163.367
R318 B.n156 B.n155 163.367
R319 B.n155 B.n154 163.367
R320 B.n154 B.n2 163.367
R321 B.n582 B.n2 163.367
R322 B.n582 B.n581 163.367
R323 B.n581 B.n580 163.367
R324 B.n580 B.n3 163.367
R325 B.n576 B.n3 163.367
R326 B.n576 B.n575 163.367
R327 B.n575 B.n574 163.367
R328 B.n574 B.n5 163.367
R329 B.n570 B.n5 163.367
R330 B.n570 B.n569 163.367
R331 B.n569 B.n568 163.367
R332 B.n568 B.n7 163.367
R333 B.n564 B.n7 163.367
R334 B.n564 B.n563 163.367
R335 B.n563 B.n562 163.367
R336 B.n562 B.n9 163.367
R337 B.n558 B.n9 163.367
R338 B.n558 B.n557 163.367
R339 B.n557 B.n556 163.367
R340 B.n556 B.n11 163.367
R341 B.n552 B.n11 163.367
R342 B.n184 B.n143 163.367
R343 B.n185 B.n184 163.367
R344 B.n186 B.n185 163.367
R345 B.n186 B.n141 163.367
R346 B.n190 B.n141 163.367
R347 B.n191 B.n190 163.367
R348 B.n192 B.n191 163.367
R349 B.n192 B.n139 163.367
R350 B.n196 B.n139 163.367
R351 B.n197 B.n196 163.367
R352 B.n198 B.n197 163.367
R353 B.n198 B.n137 163.367
R354 B.n202 B.n137 163.367
R355 B.n203 B.n202 163.367
R356 B.n204 B.n203 163.367
R357 B.n204 B.n135 163.367
R358 B.n208 B.n135 163.367
R359 B.n209 B.n208 163.367
R360 B.n210 B.n209 163.367
R361 B.n210 B.n133 163.367
R362 B.n214 B.n133 163.367
R363 B.n215 B.n214 163.367
R364 B.n216 B.n215 163.367
R365 B.n216 B.n131 163.367
R366 B.n220 B.n131 163.367
R367 B.n221 B.n220 163.367
R368 B.n222 B.n221 163.367
R369 B.n222 B.n129 163.367
R370 B.n226 B.n129 163.367
R371 B.n227 B.n226 163.367
R372 B.n228 B.n227 163.367
R373 B.n228 B.n127 163.367
R374 B.n232 B.n127 163.367
R375 B.n233 B.n232 163.367
R376 B.n234 B.n233 163.367
R377 B.n234 B.n125 163.367
R378 B.n238 B.n125 163.367
R379 B.n239 B.n238 163.367
R380 B.n240 B.n239 163.367
R381 B.n240 B.n123 163.367
R382 B.n244 B.n123 163.367
R383 B.n245 B.n244 163.367
R384 B.n246 B.n245 163.367
R385 B.n246 B.n121 163.367
R386 B.n250 B.n121 163.367
R387 B.n251 B.n250 163.367
R388 B.n251 B.n117 163.367
R389 B.n255 B.n117 163.367
R390 B.n256 B.n255 163.367
R391 B.n257 B.n256 163.367
R392 B.n257 B.n115 163.367
R393 B.n261 B.n115 163.367
R394 B.n262 B.n261 163.367
R395 B.n263 B.n262 163.367
R396 B.n263 B.n111 163.367
R397 B.n268 B.n111 163.367
R398 B.n269 B.n268 163.367
R399 B.n270 B.n269 163.367
R400 B.n270 B.n109 163.367
R401 B.n274 B.n109 163.367
R402 B.n275 B.n274 163.367
R403 B.n276 B.n275 163.367
R404 B.n276 B.n107 163.367
R405 B.n280 B.n107 163.367
R406 B.n281 B.n280 163.367
R407 B.n282 B.n281 163.367
R408 B.n282 B.n105 163.367
R409 B.n286 B.n105 163.367
R410 B.n287 B.n286 163.367
R411 B.n288 B.n287 163.367
R412 B.n288 B.n103 163.367
R413 B.n292 B.n103 163.367
R414 B.n293 B.n292 163.367
R415 B.n294 B.n293 163.367
R416 B.n294 B.n101 163.367
R417 B.n298 B.n101 163.367
R418 B.n299 B.n298 163.367
R419 B.n300 B.n299 163.367
R420 B.n300 B.n99 163.367
R421 B.n304 B.n99 163.367
R422 B.n305 B.n304 163.367
R423 B.n306 B.n305 163.367
R424 B.n306 B.n97 163.367
R425 B.n310 B.n97 163.367
R426 B.n311 B.n310 163.367
R427 B.n312 B.n311 163.367
R428 B.n312 B.n95 163.367
R429 B.n316 B.n95 163.367
R430 B.n317 B.n316 163.367
R431 B.n318 B.n317 163.367
R432 B.n318 B.n93 163.367
R433 B.n322 B.n93 163.367
R434 B.n323 B.n322 163.367
R435 B.n324 B.n323 163.367
R436 B.n324 B.n91 163.367
R437 B.n328 B.n91 163.367
R438 B.n329 B.n328 163.367
R439 B.n330 B.n329 163.367
R440 B.n330 B.n89 163.367
R441 B.n334 B.n89 163.367
R442 B.n335 B.n334 163.367
R443 B.n336 B.n87 163.367
R444 B.n340 B.n87 163.367
R445 B.n341 B.n340 163.367
R446 B.n342 B.n341 163.367
R447 B.n342 B.n85 163.367
R448 B.n346 B.n85 163.367
R449 B.n347 B.n346 163.367
R450 B.n348 B.n347 163.367
R451 B.n348 B.n83 163.367
R452 B.n352 B.n83 163.367
R453 B.n353 B.n352 163.367
R454 B.n354 B.n353 163.367
R455 B.n354 B.n81 163.367
R456 B.n358 B.n81 163.367
R457 B.n359 B.n358 163.367
R458 B.n360 B.n359 163.367
R459 B.n360 B.n79 163.367
R460 B.n364 B.n79 163.367
R461 B.n365 B.n364 163.367
R462 B.n366 B.n365 163.367
R463 B.n366 B.n77 163.367
R464 B.n370 B.n77 163.367
R465 B.n371 B.n370 163.367
R466 B.n372 B.n371 163.367
R467 B.n372 B.n75 163.367
R468 B.n376 B.n75 163.367
R469 B.n377 B.n376 163.367
R470 B.n378 B.n377 163.367
R471 B.n378 B.n73 163.367
R472 B.n382 B.n73 163.367
R473 B.n383 B.n382 163.367
R474 B.n384 B.n383 163.367
R475 B.n384 B.n71 163.367
R476 B.n388 B.n71 163.367
R477 B.n389 B.n388 163.367
R478 B.n390 B.n389 163.367
R479 B.n390 B.n69 163.367
R480 B.n394 B.n69 163.367
R481 B.n395 B.n394 163.367
R482 B.n396 B.n395 163.367
R483 B.n551 B.n550 163.367
R484 B.n550 B.n13 163.367
R485 B.n546 B.n13 163.367
R486 B.n546 B.n545 163.367
R487 B.n545 B.n544 163.367
R488 B.n544 B.n15 163.367
R489 B.n540 B.n15 163.367
R490 B.n540 B.n539 163.367
R491 B.n539 B.n538 163.367
R492 B.n538 B.n17 163.367
R493 B.n534 B.n17 163.367
R494 B.n534 B.n533 163.367
R495 B.n533 B.n532 163.367
R496 B.n532 B.n19 163.367
R497 B.n528 B.n19 163.367
R498 B.n528 B.n527 163.367
R499 B.n527 B.n526 163.367
R500 B.n526 B.n21 163.367
R501 B.n522 B.n21 163.367
R502 B.n522 B.n521 163.367
R503 B.n521 B.n520 163.367
R504 B.n520 B.n23 163.367
R505 B.n516 B.n23 163.367
R506 B.n516 B.n515 163.367
R507 B.n515 B.n514 163.367
R508 B.n514 B.n25 163.367
R509 B.n510 B.n25 163.367
R510 B.n510 B.n509 163.367
R511 B.n509 B.n508 163.367
R512 B.n508 B.n27 163.367
R513 B.n504 B.n27 163.367
R514 B.n504 B.n503 163.367
R515 B.n503 B.n502 163.367
R516 B.n502 B.n29 163.367
R517 B.n498 B.n29 163.367
R518 B.n498 B.n497 163.367
R519 B.n497 B.n496 163.367
R520 B.n496 B.n31 163.367
R521 B.n492 B.n31 163.367
R522 B.n492 B.n491 163.367
R523 B.n491 B.n490 163.367
R524 B.n490 B.n33 163.367
R525 B.n486 B.n33 163.367
R526 B.n486 B.n485 163.367
R527 B.n485 B.n484 163.367
R528 B.n484 B.n35 163.367
R529 B.n479 B.n35 163.367
R530 B.n479 B.n478 163.367
R531 B.n478 B.n477 163.367
R532 B.n477 B.n39 163.367
R533 B.n473 B.n39 163.367
R534 B.n473 B.n472 163.367
R535 B.n472 B.n471 163.367
R536 B.n471 B.n41 163.367
R537 B.n467 B.n41 163.367
R538 B.n467 B.n466 163.367
R539 B.n466 B.n45 163.367
R540 B.n462 B.n45 163.367
R541 B.n462 B.n461 163.367
R542 B.n461 B.n460 163.367
R543 B.n460 B.n47 163.367
R544 B.n456 B.n47 163.367
R545 B.n456 B.n455 163.367
R546 B.n455 B.n454 163.367
R547 B.n454 B.n49 163.367
R548 B.n450 B.n49 163.367
R549 B.n450 B.n449 163.367
R550 B.n449 B.n448 163.367
R551 B.n448 B.n51 163.367
R552 B.n444 B.n51 163.367
R553 B.n444 B.n443 163.367
R554 B.n443 B.n442 163.367
R555 B.n442 B.n53 163.367
R556 B.n438 B.n53 163.367
R557 B.n438 B.n437 163.367
R558 B.n437 B.n436 163.367
R559 B.n436 B.n55 163.367
R560 B.n432 B.n55 163.367
R561 B.n432 B.n431 163.367
R562 B.n431 B.n430 163.367
R563 B.n430 B.n57 163.367
R564 B.n426 B.n57 163.367
R565 B.n426 B.n425 163.367
R566 B.n425 B.n424 163.367
R567 B.n424 B.n59 163.367
R568 B.n420 B.n59 163.367
R569 B.n420 B.n419 163.367
R570 B.n419 B.n418 163.367
R571 B.n418 B.n61 163.367
R572 B.n414 B.n61 163.367
R573 B.n414 B.n413 163.367
R574 B.n413 B.n412 163.367
R575 B.n412 B.n63 163.367
R576 B.n408 B.n63 163.367
R577 B.n408 B.n407 163.367
R578 B.n407 B.n406 163.367
R579 B.n406 B.n65 163.367
R580 B.n402 B.n65 163.367
R581 B.n402 B.n401 163.367
R582 B.n401 B.n400 163.367
R583 B.n400 B.n67 163.367
R584 B.n266 B.n113 59.5399
R585 B.n120 B.n119 59.5399
R586 B.n482 B.n37 59.5399
R587 B.n44 B.n43 59.5399
R588 B.n113 B.n112 39.952
R589 B.n119 B.n118 39.952
R590 B.n37 B.n36 39.952
R591 B.n43 B.n42 39.952
R592 B.n553 B.n12 34.8103
R593 B.n398 B.n397 34.8103
R594 B.n337 B.n88 34.8103
R595 B.n182 B.n181 34.8103
R596 B B.n583 18.0485
R597 B.n549 B.n12 10.6151
R598 B.n549 B.n548 10.6151
R599 B.n548 B.n547 10.6151
R600 B.n547 B.n14 10.6151
R601 B.n543 B.n14 10.6151
R602 B.n543 B.n542 10.6151
R603 B.n542 B.n541 10.6151
R604 B.n541 B.n16 10.6151
R605 B.n537 B.n16 10.6151
R606 B.n537 B.n536 10.6151
R607 B.n536 B.n535 10.6151
R608 B.n535 B.n18 10.6151
R609 B.n531 B.n18 10.6151
R610 B.n531 B.n530 10.6151
R611 B.n530 B.n529 10.6151
R612 B.n529 B.n20 10.6151
R613 B.n525 B.n20 10.6151
R614 B.n525 B.n524 10.6151
R615 B.n524 B.n523 10.6151
R616 B.n523 B.n22 10.6151
R617 B.n519 B.n22 10.6151
R618 B.n519 B.n518 10.6151
R619 B.n518 B.n517 10.6151
R620 B.n517 B.n24 10.6151
R621 B.n513 B.n24 10.6151
R622 B.n513 B.n512 10.6151
R623 B.n512 B.n511 10.6151
R624 B.n511 B.n26 10.6151
R625 B.n507 B.n26 10.6151
R626 B.n507 B.n506 10.6151
R627 B.n506 B.n505 10.6151
R628 B.n505 B.n28 10.6151
R629 B.n501 B.n28 10.6151
R630 B.n501 B.n500 10.6151
R631 B.n500 B.n499 10.6151
R632 B.n499 B.n30 10.6151
R633 B.n495 B.n30 10.6151
R634 B.n495 B.n494 10.6151
R635 B.n494 B.n493 10.6151
R636 B.n493 B.n32 10.6151
R637 B.n489 B.n32 10.6151
R638 B.n489 B.n488 10.6151
R639 B.n488 B.n487 10.6151
R640 B.n487 B.n34 10.6151
R641 B.n483 B.n34 10.6151
R642 B.n481 B.n480 10.6151
R643 B.n480 B.n38 10.6151
R644 B.n476 B.n38 10.6151
R645 B.n476 B.n475 10.6151
R646 B.n475 B.n474 10.6151
R647 B.n474 B.n40 10.6151
R648 B.n470 B.n40 10.6151
R649 B.n470 B.n469 10.6151
R650 B.n469 B.n468 10.6151
R651 B.n465 B.n464 10.6151
R652 B.n464 B.n463 10.6151
R653 B.n463 B.n46 10.6151
R654 B.n459 B.n46 10.6151
R655 B.n459 B.n458 10.6151
R656 B.n458 B.n457 10.6151
R657 B.n457 B.n48 10.6151
R658 B.n453 B.n48 10.6151
R659 B.n453 B.n452 10.6151
R660 B.n452 B.n451 10.6151
R661 B.n451 B.n50 10.6151
R662 B.n447 B.n50 10.6151
R663 B.n447 B.n446 10.6151
R664 B.n446 B.n445 10.6151
R665 B.n445 B.n52 10.6151
R666 B.n441 B.n52 10.6151
R667 B.n441 B.n440 10.6151
R668 B.n440 B.n439 10.6151
R669 B.n439 B.n54 10.6151
R670 B.n435 B.n54 10.6151
R671 B.n435 B.n434 10.6151
R672 B.n434 B.n433 10.6151
R673 B.n433 B.n56 10.6151
R674 B.n429 B.n56 10.6151
R675 B.n429 B.n428 10.6151
R676 B.n428 B.n427 10.6151
R677 B.n427 B.n58 10.6151
R678 B.n423 B.n58 10.6151
R679 B.n423 B.n422 10.6151
R680 B.n422 B.n421 10.6151
R681 B.n421 B.n60 10.6151
R682 B.n417 B.n60 10.6151
R683 B.n417 B.n416 10.6151
R684 B.n416 B.n415 10.6151
R685 B.n415 B.n62 10.6151
R686 B.n411 B.n62 10.6151
R687 B.n411 B.n410 10.6151
R688 B.n410 B.n409 10.6151
R689 B.n409 B.n64 10.6151
R690 B.n405 B.n64 10.6151
R691 B.n405 B.n404 10.6151
R692 B.n404 B.n403 10.6151
R693 B.n403 B.n66 10.6151
R694 B.n399 B.n66 10.6151
R695 B.n399 B.n398 10.6151
R696 B.n338 B.n337 10.6151
R697 B.n339 B.n338 10.6151
R698 B.n339 B.n86 10.6151
R699 B.n343 B.n86 10.6151
R700 B.n344 B.n343 10.6151
R701 B.n345 B.n344 10.6151
R702 B.n345 B.n84 10.6151
R703 B.n349 B.n84 10.6151
R704 B.n350 B.n349 10.6151
R705 B.n351 B.n350 10.6151
R706 B.n351 B.n82 10.6151
R707 B.n355 B.n82 10.6151
R708 B.n356 B.n355 10.6151
R709 B.n357 B.n356 10.6151
R710 B.n357 B.n80 10.6151
R711 B.n361 B.n80 10.6151
R712 B.n362 B.n361 10.6151
R713 B.n363 B.n362 10.6151
R714 B.n363 B.n78 10.6151
R715 B.n367 B.n78 10.6151
R716 B.n368 B.n367 10.6151
R717 B.n369 B.n368 10.6151
R718 B.n369 B.n76 10.6151
R719 B.n373 B.n76 10.6151
R720 B.n374 B.n373 10.6151
R721 B.n375 B.n374 10.6151
R722 B.n375 B.n74 10.6151
R723 B.n379 B.n74 10.6151
R724 B.n380 B.n379 10.6151
R725 B.n381 B.n380 10.6151
R726 B.n381 B.n72 10.6151
R727 B.n385 B.n72 10.6151
R728 B.n386 B.n385 10.6151
R729 B.n387 B.n386 10.6151
R730 B.n387 B.n70 10.6151
R731 B.n391 B.n70 10.6151
R732 B.n392 B.n391 10.6151
R733 B.n393 B.n392 10.6151
R734 B.n393 B.n68 10.6151
R735 B.n397 B.n68 10.6151
R736 B.n183 B.n182 10.6151
R737 B.n183 B.n142 10.6151
R738 B.n187 B.n142 10.6151
R739 B.n188 B.n187 10.6151
R740 B.n189 B.n188 10.6151
R741 B.n189 B.n140 10.6151
R742 B.n193 B.n140 10.6151
R743 B.n194 B.n193 10.6151
R744 B.n195 B.n194 10.6151
R745 B.n195 B.n138 10.6151
R746 B.n199 B.n138 10.6151
R747 B.n200 B.n199 10.6151
R748 B.n201 B.n200 10.6151
R749 B.n201 B.n136 10.6151
R750 B.n205 B.n136 10.6151
R751 B.n206 B.n205 10.6151
R752 B.n207 B.n206 10.6151
R753 B.n207 B.n134 10.6151
R754 B.n211 B.n134 10.6151
R755 B.n212 B.n211 10.6151
R756 B.n213 B.n212 10.6151
R757 B.n213 B.n132 10.6151
R758 B.n217 B.n132 10.6151
R759 B.n218 B.n217 10.6151
R760 B.n219 B.n218 10.6151
R761 B.n219 B.n130 10.6151
R762 B.n223 B.n130 10.6151
R763 B.n224 B.n223 10.6151
R764 B.n225 B.n224 10.6151
R765 B.n225 B.n128 10.6151
R766 B.n229 B.n128 10.6151
R767 B.n230 B.n229 10.6151
R768 B.n231 B.n230 10.6151
R769 B.n231 B.n126 10.6151
R770 B.n235 B.n126 10.6151
R771 B.n236 B.n235 10.6151
R772 B.n237 B.n236 10.6151
R773 B.n237 B.n124 10.6151
R774 B.n241 B.n124 10.6151
R775 B.n242 B.n241 10.6151
R776 B.n243 B.n242 10.6151
R777 B.n243 B.n122 10.6151
R778 B.n247 B.n122 10.6151
R779 B.n248 B.n247 10.6151
R780 B.n249 B.n248 10.6151
R781 B.n253 B.n252 10.6151
R782 B.n254 B.n253 10.6151
R783 B.n254 B.n116 10.6151
R784 B.n258 B.n116 10.6151
R785 B.n259 B.n258 10.6151
R786 B.n260 B.n259 10.6151
R787 B.n260 B.n114 10.6151
R788 B.n264 B.n114 10.6151
R789 B.n265 B.n264 10.6151
R790 B.n267 B.n110 10.6151
R791 B.n271 B.n110 10.6151
R792 B.n272 B.n271 10.6151
R793 B.n273 B.n272 10.6151
R794 B.n273 B.n108 10.6151
R795 B.n277 B.n108 10.6151
R796 B.n278 B.n277 10.6151
R797 B.n279 B.n278 10.6151
R798 B.n279 B.n106 10.6151
R799 B.n283 B.n106 10.6151
R800 B.n284 B.n283 10.6151
R801 B.n285 B.n284 10.6151
R802 B.n285 B.n104 10.6151
R803 B.n289 B.n104 10.6151
R804 B.n290 B.n289 10.6151
R805 B.n291 B.n290 10.6151
R806 B.n291 B.n102 10.6151
R807 B.n295 B.n102 10.6151
R808 B.n296 B.n295 10.6151
R809 B.n297 B.n296 10.6151
R810 B.n297 B.n100 10.6151
R811 B.n301 B.n100 10.6151
R812 B.n302 B.n301 10.6151
R813 B.n303 B.n302 10.6151
R814 B.n303 B.n98 10.6151
R815 B.n307 B.n98 10.6151
R816 B.n308 B.n307 10.6151
R817 B.n309 B.n308 10.6151
R818 B.n309 B.n96 10.6151
R819 B.n313 B.n96 10.6151
R820 B.n314 B.n313 10.6151
R821 B.n315 B.n314 10.6151
R822 B.n315 B.n94 10.6151
R823 B.n319 B.n94 10.6151
R824 B.n320 B.n319 10.6151
R825 B.n321 B.n320 10.6151
R826 B.n321 B.n92 10.6151
R827 B.n325 B.n92 10.6151
R828 B.n326 B.n325 10.6151
R829 B.n327 B.n326 10.6151
R830 B.n327 B.n90 10.6151
R831 B.n331 B.n90 10.6151
R832 B.n332 B.n331 10.6151
R833 B.n333 B.n332 10.6151
R834 B.n333 B.n88 10.6151
R835 B.n181 B.n144 10.6151
R836 B.n177 B.n144 10.6151
R837 B.n177 B.n176 10.6151
R838 B.n176 B.n175 10.6151
R839 B.n175 B.n146 10.6151
R840 B.n171 B.n146 10.6151
R841 B.n171 B.n170 10.6151
R842 B.n170 B.n169 10.6151
R843 B.n169 B.n148 10.6151
R844 B.n165 B.n148 10.6151
R845 B.n165 B.n164 10.6151
R846 B.n164 B.n163 10.6151
R847 B.n163 B.n150 10.6151
R848 B.n159 B.n150 10.6151
R849 B.n159 B.n158 10.6151
R850 B.n158 B.n157 10.6151
R851 B.n157 B.n152 10.6151
R852 B.n153 B.n152 10.6151
R853 B.n153 B.n0 10.6151
R854 B.n579 B.n1 10.6151
R855 B.n579 B.n578 10.6151
R856 B.n578 B.n577 10.6151
R857 B.n577 B.n4 10.6151
R858 B.n573 B.n4 10.6151
R859 B.n573 B.n572 10.6151
R860 B.n572 B.n571 10.6151
R861 B.n571 B.n6 10.6151
R862 B.n567 B.n6 10.6151
R863 B.n567 B.n566 10.6151
R864 B.n566 B.n565 10.6151
R865 B.n565 B.n8 10.6151
R866 B.n561 B.n8 10.6151
R867 B.n561 B.n560 10.6151
R868 B.n560 B.n559 10.6151
R869 B.n559 B.n10 10.6151
R870 B.n555 B.n10 10.6151
R871 B.n555 B.n554 10.6151
R872 B.n554 B.n553 10.6151
R873 B.n483 B.n482 9.36635
R874 B.n465 B.n44 9.36635
R875 B.n249 B.n120 9.36635
R876 B.n267 B.n266 9.36635
R877 B.n583 B.n0 2.81026
R878 B.n583 B.n1 2.81026
R879 B.n482 B.n481 1.24928
R880 B.n468 B.n44 1.24928
R881 B.n252 B.n120 1.24928
R882 B.n266 B.n265 1.24928
R883 VN VN.t1 291.459
R884 VN VN.t0 247.976
R885 VTAIL.n290 VTAIL.n222 756.745
R886 VTAIL.n68 VTAIL.n0 756.745
R887 VTAIL.n216 VTAIL.n148 756.745
R888 VTAIL.n142 VTAIL.n74 756.745
R889 VTAIL.n247 VTAIL.n246 585
R890 VTAIL.n249 VTAIL.n248 585
R891 VTAIL.n242 VTAIL.n241 585
R892 VTAIL.n255 VTAIL.n254 585
R893 VTAIL.n257 VTAIL.n256 585
R894 VTAIL.n238 VTAIL.n237 585
R895 VTAIL.n264 VTAIL.n263 585
R896 VTAIL.n265 VTAIL.n236 585
R897 VTAIL.n267 VTAIL.n266 585
R898 VTAIL.n234 VTAIL.n233 585
R899 VTAIL.n273 VTAIL.n272 585
R900 VTAIL.n275 VTAIL.n274 585
R901 VTAIL.n230 VTAIL.n229 585
R902 VTAIL.n281 VTAIL.n280 585
R903 VTAIL.n283 VTAIL.n282 585
R904 VTAIL.n226 VTAIL.n225 585
R905 VTAIL.n289 VTAIL.n288 585
R906 VTAIL.n291 VTAIL.n290 585
R907 VTAIL.n25 VTAIL.n24 585
R908 VTAIL.n27 VTAIL.n26 585
R909 VTAIL.n20 VTAIL.n19 585
R910 VTAIL.n33 VTAIL.n32 585
R911 VTAIL.n35 VTAIL.n34 585
R912 VTAIL.n16 VTAIL.n15 585
R913 VTAIL.n42 VTAIL.n41 585
R914 VTAIL.n43 VTAIL.n14 585
R915 VTAIL.n45 VTAIL.n44 585
R916 VTAIL.n12 VTAIL.n11 585
R917 VTAIL.n51 VTAIL.n50 585
R918 VTAIL.n53 VTAIL.n52 585
R919 VTAIL.n8 VTAIL.n7 585
R920 VTAIL.n59 VTAIL.n58 585
R921 VTAIL.n61 VTAIL.n60 585
R922 VTAIL.n4 VTAIL.n3 585
R923 VTAIL.n67 VTAIL.n66 585
R924 VTAIL.n69 VTAIL.n68 585
R925 VTAIL.n217 VTAIL.n216 585
R926 VTAIL.n215 VTAIL.n214 585
R927 VTAIL.n152 VTAIL.n151 585
R928 VTAIL.n209 VTAIL.n208 585
R929 VTAIL.n207 VTAIL.n206 585
R930 VTAIL.n156 VTAIL.n155 585
R931 VTAIL.n201 VTAIL.n200 585
R932 VTAIL.n199 VTAIL.n198 585
R933 VTAIL.n160 VTAIL.n159 585
R934 VTAIL.n164 VTAIL.n162 585
R935 VTAIL.n193 VTAIL.n192 585
R936 VTAIL.n191 VTAIL.n190 585
R937 VTAIL.n166 VTAIL.n165 585
R938 VTAIL.n185 VTAIL.n184 585
R939 VTAIL.n183 VTAIL.n182 585
R940 VTAIL.n170 VTAIL.n169 585
R941 VTAIL.n177 VTAIL.n176 585
R942 VTAIL.n175 VTAIL.n174 585
R943 VTAIL.n143 VTAIL.n142 585
R944 VTAIL.n141 VTAIL.n140 585
R945 VTAIL.n78 VTAIL.n77 585
R946 VTAIL.n135 VTAIL.n134 585
R947 VTAIL.n133 VTAIL.n132 585
R948 VTAIL.n82 VTAIL.n81 585
R949 VTAIL.n127 VTAIL.n126 585
R950 VTAIL.n125 VTAIL.n124 585
R951 VTAIL.n86 VTAIL.n85 585
R952 VTAIL.n90 VTAIL.n88 585
R953 VTAIL.n119 VTAIL.n118 585
R954 VTAIL.n117 VTAIL.n116 585
R955 VTAIL.n92 VTAIL.n91 585
R956 VTAIL.n111 VTAIL.n110 585
R957 VTAIL.n109 VTAIL.n108 585
R958 VTAIL.n96 VTAIL.n95 585
R959 VTAIL.n103 VTAIL.n102 585
R960 VTAIL.n101 VTAIL.n100 585
R961 VTAIL.n245 VTAIL.t3 329.036
R962 VTAIL.n23 VTAIL.t1 329.036
R963 VTAIL.n173 VTAIL.t0 329.036
R964 VTAIL.n99 VTAIL.t2 329.036
R965 VTAIL.n248 VTAIL.n247 171.744
R966 VTAIL.n248 VTAIL.n241 171.744
R967 VTAIL.n255 VTAIL.n241 171.744
R968 VTAIL.n256 VTAIL.n255 171.744
R969 VTAIL.n256 VTAIL.n237 171.744
R970 VTAIL.n264 VTAIL.n237 171.744
R971 VTAIL.n265 VTAIL.n264 171.744
R972 VTAIL.n266 VTAIL.n265 171.744
R973 VTAIL.n266 VTAIL.n233 171.744
R974 VTAIL.n273 VTAIL.n233 171.744
R975 VTAIL.n274 VTAIL.n273 171.744
R976 VTAIL.n274 VTAIL.n229 171.744
R977 VTAIL.n281 VTAIL.n229 171.744
R978 VTAIL.n282 VTAIL.n281 171.744
R979 VTAIL.n282 VTAIL.n225 171.744
R980 VTAIL.n289 VTAIL.n225 171.744
R981 VTAIL.n290 VTAIL.n289 171.744
R982 VTAIL.n26 VTAIL.n25 171.744
R983 VTAIL.n26 VTAIL.n19 171.744
R984 VTAIL.n33 VTAIL.n19 171.744
R985 VTAIL.n34 VTAIL.n33 171.744
R986 VTAIL.n34 VTAIL.n15 171.744
R987 VTAIL.n42 VTAIL.n15 171.744
R988 VTAIL.n43 VTAIL.n42 171.744
R989 VTAIL.n44 VTAIL.n43 171.744
R990 VTAIL.n44 VTAIL.n11 171.744
R991 VTAIL.n51 VTAIL.n11 171.744
R992 VTAIL.n52 VTAIL.n51 171.744
R993 VTAIL.n52 VTAIL.n7 171.744
R994 VTAIL.n59 VTAIL.n7 171.744
R995 VTAIL.n60 VTAIL.n59 171.744
R996 VTAIL.n60 VTAIL.n3 171.744
R997 VTAIL.n67 VTAIL.n3 171.744
R998 VTAIL.n68 VTAIL.n67 171.744
R999 VTAIL.n216 VTAIL.n215 171.744
R1000 VTAIL.n215 VTAIL.n151 171.744
R1001 VTAIL.n208 VTAIL.n151 171.744
R1002 VTAIL.n208 VTAIL.n207 171.744
R1003 VTAIL.n207 VTAIL.n155 171.744
R1004 VTAIL.n200 VTAIL.n155 171.744
R1005 VTAIL.n200 VTAIL.n199 171.744
R1006 VTAIL.n199 VTAIL.n159 171.744
R1007 VTAIL.n164 VTAIL.n159 171.744
R1008 VTAIL.n192 VTAIL.n164 171.744
R1009 VTAIL.n192 VTAIL.n191 171.744
R1010 VTAIL.n191 VTAIL.n165 171.744
R1011 VTAIL.n184 VTAIL.n165 171.744
R1012 VTAIL.n184 VTAIL.n183 171.744
R1013 VTAIL.n183 VTAIL.n169 171.744
R1014 VTAIL.n176 VTAIL.n169 171.744
R1015 VTAIL.n176 VTAIL.n175 171.744
R1016 VTAIL.n142 VTAIL.n141 171.744
R1017 VTAIL.n141 VTAIL.n77 171.744
R1018 VTAIL.n134 VTAIL.n77 171.744
R1019 VTAIL.n134 VTAIL.n133 171.744
R1020 VTAIL.n133 VTAIL.n81 171.744
R1021 VTAIL.n126 VTAIL.n81 171.744
R1022 VTAIL.n126 VTAIL.n125 171.744
R1023 VTAIL.n125 VTAIL.n85 171.744
R1024 VTAIL.n90 VTAIL.n85 171.744
R1025 VTAIL.n118 VTAIL.n90 171.744
R1026 VTAIL.n118 VTAIL.n117 171.744
R1027 VTAIL.n117 VTAIL.n91 171.744
R1028 VTAIL.n110 VTAIL.n91 171.744
R1029 VTAIL.n110 VTAIL.n109 171.744
R1030 VTAIL.n109 VTAIL.n95 171.744
R1031 VTAIL.n102 VTAIL.n95 171.744
R1032 VTAIL.n102 VTAIL.n101 171.744
R1033 VTAIL.n247 VTAIL.t3 85.8723
R1034 VTAIL.n25 VTAIL.t1 85.8723
R1035 VTAIL.n175 VTAIL.t0 85.8723
R1036 VTAIL.n101 VTAIL.t2 85.8723
R1037 VTAIL.n295 VTAIL.n294 32.1853
R1038 VTAIL.n73 VTAIL.n72 32.1853
R1039 VTAIL.n221 VTAIL.n220 32.1853
R1040 VTAIL.n147 VTAIL.n146 32.1853
R1041 VTAIL.n147 VTAIL.n73 27.6083
R1042 VTAIL.n295 VTAIL.n221 25.8324
R1043 VTAIL.n267 VTAIL.n234 13.1884
R1044 VTAIL.n45 VTAIL.n12 13.1884
R1045 VTAIL.n162 VTAIL.n160 13.1884
R1046 VTAIL.n88 VTAIL.n86 13.1884
R1047 VTAIL.n268 VTAIL.n236 12.8005
R1048 VTAIL.n272 VTAIL.n271 12.8005
R1049 VTAIL.n46 VTAIL.n14 12.8005
R1050 VTAIL.n50 VTAIL.n49 12.8005
R1051 VTAIL.n198 VTAIL.n197 12.8005
R1052 VTAIL.n194 VTAIL.n193 12.8005
R1053 VTAIL.n124 VTAIL.n123 12.8005
R1054 VTAIL.n120 VTAIL.n119 12.8005
R1055 VTAIL.n263 VTAIL.n262 12.0247
R1056 VTAIL.n275 VTAIL.n232 12.0247
R1057 VTAIL.n41 VTAIL.n40 12.0247
R1058 VTAIL.n53 VTAIL.n10 12.0247
R1059 VTAIL.n201 VTAIL.n158 12.0247
R1060 VTAIL.n190 VTAIL.n163 12.0247
R1061 VTAIL.n127 VTAIL.n84 12.0247
R1062 VTAIL.n116 VTAIL.n89 12.0247
R1063 VTAIL.n261 VTAIL.n238 11.249
R1064 VTAIL.n276 VTAIL.n230 11.249
R1065 VTAIL.n39 VTAIL.n16 11.249
R1066 VTAIL.n54 VTAIL.n8 11.249
R1067 VTAIL.n202 VTAIL.n156 11.249
R1068 VTAIL.n189 VTAIL.n166 11.249
R1069 VTAIL.n128 VTAIL.n82 11.249
R1070 VTAIL.n115 VTAIL.n92 11.249
R1071 VTAIL.n246 VTAIL.n245 10.7239
R1072 VTAIL.n24 VTAIL.n23 10.7239
R1073 VTAIL.n174 VTAIL.n173 10.7239
R1074 VTAIL.n100 VTAIL.n99 10.7239
R1075 VTAIL.n258 VTAIL.n257 10.4732
R1076 VTAIL.n280 VTAIL.n279 10.4732
R1077 VTAIL.n36 VTAIL.n35 10.4732
R1078 VTAIL.n58 VTAIL.n57 10.4732
R1079 VTAIL.n206 VTAIL.n205 10.4732
R1080 VTAIL.n186 VTAIL.n185 10.4732
R1081 VTAIL.n132 VTAIL.n131 10.4732
R1082 VTAIL.n112 VTAIL.n111 10.4732
R1083 VTAIL.n254 VTAIL.n240 9.69747
R1084 VTAIL.n283 VTAIL.n228 9.69747
R1085 VTAIL.n32 VTAIL.n18 9.69747
R1086 VTAIL.n61 VTAIL.n6 9.69747
R1087 VTAIL.n209 VTAIL.n154 9.69747
R1088 VTAIL.n182 VTAIL.n168 9.69747
R1089 VTAIL.n135 VTAIL.n80 9.69747
R1090 VTAIL.n108 VTAIL.n94 9.69747
R1091 VTAIL.n294 VTAIL.n293 9.45567
R1092 VTAIL.n72 VTAIL.n71 9.45567
R1093 VTAIL.n220 VTAIL.n219 9.45567
R1094 VTAIL.n146 VTAIL.n145 9.45567
R1095 VTAIL.n293 VTAIL.n292 9.3005
R1096 VTAIL.n287 VTAIL.n286 9.3005
R1097 VTAIL.n285 VTAIL.n284 9.3005
R1098 VTAIL.n228 VTAIL.n227 9.3005
R1099 VTAIL.n279 VTAIL.n278 9.3005
R1100 VTAIL.n277 VTAIL.n276 9.3005
R1101 VTAIL.n232 VTAIL.n231 9.3005
R1102 VTAIL.n271 VTAIL.n270 9.3005
R1103 VTAIL.n244 VTAIL.n243 9.3005
R1104 VTAIL.n251 VTAIL.n250 9.3005
R1105 VTAIL.n253 VTAIL.n252 9.3005
R1106 VTAIL.n240 VTAIL.n239 9.3005
R1107 VTAIL.n259 VTAIL.n258 9.3005
R1108 VTAIL.n261 VTAIL.n260 9.3005
R1109 VTAIL.n262 VTAIL.n235 9.3005
R1110 VTAIL.n269 VTAIL.n268 9.3005
R1111 VTAIL.n224 VTAIL.n223 9.3005
R1112 VTAIL.n71 VTAIL.n70 9.3005
R1113 VTAIL.n65 VTAIL.n64 9.3005
R1114 VTAIL.n63 VTAIL.n62 9.3005
R1115 VTAIL.n6 VTAIL.n5 9.3005
R1116 VTAIL.n57 VTAIL.n56 9.3005
R1117 VTAIL.n55 VTAIL.n54 9.3005
R1118 VTAIL.n10 VTAIL.n9 9.3005
R1119 VTAIL.n49 VTAIL.n48 9.3005
R1120 VTAIL.n22 VTAIL.n21 9.3005
R1121 VTAIL.n29 VTAIL.n28 9.3005
R1122 VTAIL.n31 VTAIL.n30 9.3005
R1123 VTAIL.n18 VTAIL.n17 9.3005
R1124 VTAIL.n37 VTAIL.n36 9.3005
R1125 VTAIL.n39 VTAIL.n38 9.3005
R1126 VTAIL.n40 VTAIL.n13 9.3005
R1127 VTAIL.n47 VTAIL.n46 9.3005
R1128 VTAIL.n2 VTAIL.n1 9.3005
R1129 VTAIL.n172 VTAIL.n171 9.3005
R1130 VTAIL.n179 VTAIL.n178 9.3005
R1131 VTAIL.n181 VTAIL.n180 9.3005
R1132 VTAIL.n168 VTAIL.n167 9.3005
R1133 VTAIL.n187 VTAIL.n186 9.3005
R1134 VTAIL.n189 VTAIL.n188 9.3005
R1135 VTAIL.n163 VTAIL.n161 9.3005
R1136 VTAIL.n195 VTAIL.n194 9.3005
R1137 VTAIL.n219 VTAIL.n218 9.3005
R1138 VTAIL.n150 VTAIL.n149 9.3005
R1139 VTAIL.n213 VTAIL.n212 9.3005
R1140 VTAIL.n211 VTAIL.n210 9.3005
R1141 VTAIL.n154 VTAIL.n153 9.3005
R1142 VTAIL.n205 VTAIL.n204 9.3005
R1143 VTAIL.n203 VTAIL.n202 9.3005
R1144 VTAIL.n158 VTAIL.n157 9.3005
R1145 VTAIL.n197 VTAIL.n196 9.3005
R1146 VTAIL.n98 VTAIL.n97 9.3005
R1147 VTAIL.n105 VTAIL.n104 9.3005
R1148 VTAIL.n107 VTAIL.n106 9.3005
R1149 VTAIL.n94 VTAIL.n93 9.3005
R1150 VTAIL.n113 VTAIL.n112 9.3005
R1151 VTAIL.n115 VTAIL.n114 9.3005
R1152 VTAIL.n89 VTAIL.n87 9.3005
R1153 VTAIL.n121 VTAIL.n120 9.3005
R1154 VTAIL.n145 VTAIL.n144 9.3005
R1155 VTAIL.n76 VTAIL.n75 9.3005
R1156 VTAIL.n139 VTAIL.n138 9.3005
R1157 VTAIL.n137 VTAIL.n136 9.3005
R1158 VTAIL.n80 VTAIL.n79 9.3005
R1159 VTAIL.n131 VTAIL.n130 9.3005
R1160 VTAIL.n129 VTAIL.n128 9.3005
R1161 VTAIL.n84 VTAIL.n83 9.3005
R1162 VTAIL.n123 VTAIL.n122 9.3005
R1163 VTAIL.n253 VTAIL.n242 8.92171
R1164 VTAIL.n284 VTAIL.n226 8.92171
R1165 VTAIL.n31 VTAIL.n20 8.92171
R1166 VTAIL.n62 VTAIL.n4 8.92171
R1167 VTAIL.n210 VTAIL.n152 8.92171
R1168 VTAIL.n181 VTAIL.n170 8.92171
R1169 VTAIL.n136 VTAIL.n78 8.92171
R1170 VTAIL.n107 VTAIL.n96 8.92171
R1171 VTAIL.n250 VTAIL.n249 8.14595
R1172 VTAIL.n288 VTAIL.n287 8.14595
R1173 VTAIL.n28 VTAIL.n27 8.14595
R1174 VTAIL.n66 VTAIL.n65 8.14595
R1175 VTAIL.n214 VTAIL.n213 8.14595
R1176 VTAIL.n178 VTAIL.n177 8.14595
R1177 VTAIL.n140 VTAIL.n139 8.14595
R1178 VTAIL.n104 VTAIL.n103 8.14595
R1179 VTAIL.n246 VTAIL.n244 7.3702
R1180 VTAIL.n291 VTAIL.n224 7.3702
R1181 VTAIL.n294 VTAIL.n222 7.3702
R1182 VTAIL.n24 VTAIL.n22 7.3702
R1183 VTAIL.n69 VTAIL.n2 7.3702
R1184 VTAIL.n72 VTAIL.n0 7.3702
R1185 VTAIL.n220 VTAIL.n148 7.3702
R1186 VTAIL.n217 VTAIL.n150 7.3702
R1187 VTAIL.n174 VTAIL.n172 7.3702
R1188 VTAIL.n146 VTAIL.n74 7.3702
R1189 VTAIL.n143 VTAIL.n76 7.3702
R1190 VTAIL.n100 VTAIL.n98 7.3702
R1191 VTAIL.n292 VTAIL.n291 6.59444
R1192 VTAIL.n292 VTAIL.n222 6.59444
R1193 VTAIL.n70 VTAIL.n69 6.59444
R1194 VTAIL.n70 VTAIL.n0 6.59444
R1195 VTAIL.n218 VTAIL.n148 6.59444
R1196 VTAIL.n218 VTAIL.n217 6.59444
R1197 VTAIL.n144 VTAIL.n74 6.59444
R1198 VTAIL.n144 VTAIL.n143 6.59444
R1199 VTAIL.n249 VTAIL.n244 5.81868
R1200 VTAIL.n288 VTAIL.n224 5.81868
R1201 VTAIL.n27 VTAIL.n22 5.81868
R1202 VTAIL.n66 VTAIL.n2 5.81868
R1203 VTAIL.n214 VTAIL.n150 5.81868
R1204 VTAIL.n177 VTAIL.n172 5.81868
R1205 VTAIL.n140 VTAIL.n76 5.81868
R1206 VTAIL.n103 VTAIL.n98 5.81868
R1207 VTAIL.n250 VTAIL.n242 5.04292
R1208 VTAIL.n287 VTAIL.n226 5.04292
R1209 VTAIL.n28 VTAIL.n20 5.04292
R1210 VTAIL.n65 VTAIL.n4 5.04292
R1211 VTAIL.n213 VTAIL.n152 5.04292
R1212 VTAIL.n178 VTAIL.n170 5.04292
R1213 VTAIL.n139 VTAIL.n78 5.04292
R1214 VTAIL.n104 VTAIL.n96 5.04292
R1215 VTAIL.n254 VTAIL.n253 4.26717
R1216 VTAIL.n284 VTAIL.n283 4.26717
R1217 VTAIL.n32 VTAIL.n31 4.26717
R1218 VTAIL.n62 VTAIL.n61 4.26717
R1219 VTAIL.n210 VTAIL.n209 4.26717
R1220 VTAIL.n182 VTAIL.n181 4.26717
R1221 VTAIL.n136 VTAIL.n135 4.26717
R1222 VTAIL.n108 VTAIL.n107 4.26717
R1223 VTAIL.n257 VTAIL.n240 3.49141
R1224 VTAIL.n280 VTAIL.n228 3.49141
R1225 VTAIL.n35 VTAIL.n18 3.49141
R1226 VTAIL.n58 VTAIL.n6 3.49141
R1227 VTAIL.n206 VTAIL.n154 3.49141
R1228 VTAIL.n185 VTAIL.n168 3.49141
R1229 VTAIL.n132 VTAIL.n80 3.49141
R1230 VTAIL.n111 VTAIL.n94 3.49141
R1231 VTAIL.n258 VTAIL.n238 2.71565
R1232 VTAIL.n279 VTAIL.n230 2.71565
R1233 VTAIL.n36 VTAIL.n16 2.71565
R1234 VTAIL.n57 VTAIL.n8 2.71565
R1235 VTAIL.n205 VTAIL.n156 2.71565
R1236 VTAIL.n186 VTAIL.n166 2.71565
R1237 VTAIL.n131 VTAIL.n82 2.71565
R1238 VTAIL.n112 VTAIL.n92 2.71565
R1239 VTAIL.n245 VTAIL.n243 2.41282
R1240 VTAIL.n23 VTAIL.n21 2.41282
R1241 VTAIL.n173 VTAIL.n171 2.41282
R1242 VTAIL.n99 VTAIL.n97 2.41282
R1243 VTAIL.n263 VTAIL.n261 1.93989
R1244 VTAIL.n276 VTAIL.n275 1.93989
R1245 VTAIL.n41 VTAIL.n39 1.93989
R1246 VTAIL.n54 VTAIL.n53 1.93989
R1247 VTAIL.n202 VTAIL.n201 1.93989
R1248 VTAIL.n190 VTAIL.n189 1.93989
R1249 VTAIL.n128 VTAIL.n127 1.93989
R1250 VTAIL.n116 VTAIL.n115 1.93989
R1251 VTAIL.n221 VTAIL.n147 1.35826
R1252 VTAIL.n262 VTAIL.n236 1.16414
R1253 VTAIL.n272 VTAIL.n232 1.16414
R1254 VTAIL.n40 VTAIL.n14 1.16414
R1255 VTAIL.n50 VTAIL.n10 1.16414
R1256 VTAIL.n198 VTAIL.n158 1.16414
R1257 VTAIL.n193 VTAIL.n163 1.16414
R1258 VTAIL.n124 VTAIL.n84 1.16414
R1259 VTAIL.n119 VTAIL.n89 1.16414
R1260 VTAIL VTAIL.n73 0.972483
R1261 VTAIL.n268 VTAIL.n267 0.388379
R1262 VTAIL.n271 VTAIL.n234 0.388379
R1263 VTAIL.n46 VTAIL.n45 0.388379
R1264 VTAIL.n49 VTAIL.n12 0.388379
R1265 VTAIL.n197 VTAIL.n160 0.388379
R1266 VTAIL.n194 VTAIL.n162 0.388379
R1267 VTAIL.n123 VTAIL.n86 0.388379
R1268 VTAIL.n120 VTAIL.n88 0.388379
R1269 VTAIL VTAIL.n295 0.386276
R1270 VTAIL.n251 VTAIL.n243 0.155672
R1271 VTAIL.n252 VTAIL.n251 0.155672
R1272 VTAIL.n252 VTAIL.n239 0.155672
R1273 VTAIL.n259 VTAIL.n239 0.155672
R1274 VTAIL.n260 VTAIL.n259 0.155672
R1275 VTAIL.n260 VTAIL.n235 0.155672
R1276 VTAIL.n269 VTAIL.n235 0.155672
R1277 VTAIL.n270 VTAIL.n269 0.155672
R1278 VTAIL.n270 VTAIL.n231 0.155672
R1279 VTAIL.n277 VTAIL.n231 0.155672
R1280 VTAIL.n278 VTAIL.n277 0.155672
R1281 VTAIL.n278 VTAIL.n227 0.155672
R1282 VTAIL.n285 VTAIL.n227 0.155672
R1283 VTAIL.n286 VTAIL.n285 0.155672
R1284 VTAIL.n286 VTAIL.n223 0.155672
R1285 VTAIL.n293 VTAIL.n223 0.155672
R1286 VTAIL.n29 VTAIL.n21 0.155672
R1287 VTAIL.n30 VTAIL.n29 0.155672
R1288 VTAIL.n30 VTAIL.n17 0.155672
R1289 VTAIL.n37 VTAIL.n17 0.155672
R1290 VTAIL.n38 VTAIL.n37 0.155672
R1291 VTAIL.n38 VTAIL.n13 0.155672
R1292 VTAIL.n47 VTAIL.n13 0.155672
R1293 VTAIL.n48 VTAIL.n47 0.155672
R1294 VTAIL.n48 VTAIL.n9 0.155672
R1295 VTAIL.n55 VTAIL.n9 0.155672
R1296 VTAIL.n56 VTAIL.n55 0.155672
R1297 VTAIL.n56 VTAIL.n5 0.155672
R1298 VTAIL.n63 VTAIL.n5 0.155672
R1299 VTAIL.n64 VTAIL.n63 0.155672
R1300 VTAIL.n64 VTAIL.n1 0.155672
R1301 VTAIL.n71 VTAIL.n1 0.155672
R1302 VTAIL.n219 VTAIL.n149 0.155672
R1303 VTAIL.n212 VTAIL.n149 0.155672
R1304 VTAIL.n212 VTAIL.n211 0.155672
R1305 VTAIL.n211 VTAIL.n153 0.155672
R1306 VTAIL.n204 VTAIL.n153 0.155672
R1307 VTAIL.n204 VTAIL.n203 0.155672
R1308 VTAIL.n203 VTAIL.n157 0.155672
R1309 VTAIL.n196 VTAIL.n157 0.155672
R1310 VTAIL.n196 VTAIL.n195 0.155672
R1311 VTAIL.n195 VTAIL.n161 0.155672
R1312 VTAIL.n188 VTAIL.n161 0.155672
R1313 VTAIL.n188 VTAIL.n187 0.155672
R1314 VTAIL.n187 VTAIL.n167 0.155672
R1315 VTAIL.n180 VTAIL.n167 0.155672
R1316 VTAIL.n180 VTAIL.n179 0.155672
R1317 VTAIL.n179 VTAIL.n171 0.155672
R1318 VTAIL.n145 VTAIL.n75 0.155672
R1319 VTAIL.n138 VTAIL.n75 0.155672
R1320 VTAIL.n138 VTAIL.n137 0.155672
R1321 VTAIL.n137 VTAIL.n79 0.155672
R1322 VTAIL.n130 VTAIL.n79 0.155672
R1323 VTAIL.n130 VTAIL.n129 0.155672
R1324 VTAIL.n129 VTAIL.n83 0.155672
R1325 VTAIL.n122 VTAIL.n83 0.155672
R1326 VTAIL.n122 VTAIL.n121 0.155672
R1327 VTAIL.n121 VTAIL.n87 0.155672
R1328 VTAIL.n114 VTAIL.n87 0.155672
R1329 VTAIL.n114 VTAIL.n113 0.155672
R1330 VTAIL.n113 VTAIL.n93 0.155672
R1331 VTAIL.n106 VTAIL.n93 0.155672
R1332 VTAIL.n106 VTAIL.n105 0.155672
R1333 VTAIL.n105 VTAIL.n97 0.155672
R1334 VDD2.n141 VDD2.n73 756.745
R1335 VDD2.n68 VDD2.n0 756.745
R1336 VDD2.n142 VDD2.n141 585
R1337 VDD2.n140 VDD2.n139 585
R1338 VDD2.n77 VDD2.n76 585
R1339 VDD2.n134 VDD2.n133 585
R1340 VDD2.n132 VDD2.n131 585
R1341 VDD2.n81 VDD2.n80 585
R1342 VDD2.n126 VDD2.n125 585
R1343 VDD2.n124 VDD2.n123 585
R1344 VDD2.n85 VDD2.n84 585
R1345 VDD2.n89 VDD2.n87 585
R1346 VDD2.n118 VDD2.n117 585
R1347 VDD2.n116 VDD2.n115 585
R1348 VDD2.n91 VDD2.n90 585
R1349 VDD2.n110 VDD2.n109 585
R1350 VDD2.n108 VDD2.n107 585
R1351 VDD2.n95 VDD2.n94 585
R1352 VDD2.n102 VDD2.n101 585
R1353 VDD2.n100 VDD2.n99 585
R1354 VDD2.n25 VDD2.n24 585
R1355 VDD2.n27 VDD2.n26 585
R1356 VDD2.n20 VDD2.n19 585
R1357 VDD2.n33 VDD2.n32 585
R1358 VDD2.n35 VDD2.n34 585
R1359 VDD2.n16 VDD2.n15 585
R1360 VDD2.n42 VDD2.n41 585
R1361 VDD2.n43 VDD2.n14 585
R1362 VDD2.n45 VDD2.n44 585
R1363 VDD2.n12 VDD2.n11 585
R1364 VDD2.n51 VDD2.n50 585
R1365 VDD2.n53 VDD2.n52 585
R1366 VDD2.n8 VDD2.n7 585
R1367 VDD2.n59 VDD2.n58 585
R1368 VDD2.n61 VDD2.n60 585
R1369 VDD2.n4 VDD2.n3 585
R1370 VDD2.n67 VDD2.n66 585
R1371 VDD2.n69 VDD2.n68 585
R1372 VDD2.n98 VDD2.t0 329.036
R1373 VDD2.n23 VDD2.t1 329.036
R1374 VDD2.n141 VDD2.n140 171.744
R1375 VDD2.n140 VDD2.n76 171.744
R1376 VDD2.n133 VDD2.n76 171.744
R1377 VDD2.n133 VDD2.n132 171.744
R1378 VDD2.n132 VDD2.n80 171.744
R1379 VDD2.n125 VDD2.n80 171.744
R1380 VDD2.n125 VDD2.n124 171.744
R1381 VDD2.n124 VDD2.n84 171.744
R1382 VDD2.n89 VDD2.n84 171.744
R1383 VDD2.n117 VDD2.n89 171.744
R1384 VDD2.n117 VDD2.n116 171.744
R1385 VDD2.n116 VDD2.n90 171.744
R1386 VDD2.n109 VDD2.n90 171.744
R1387 VDD2.n109 VDD2.n108 171.744
R1388 VDD2.n108 VDD2.n94 171.744
R1389 VDD2.n101 VDD2.n94 171.744
R1390 VDD2.n101 VDD2.n100 171.744
R1391 VDD2.n26 VDD2.n25 171.744
R1392 VDD2.n26 VDD2.n19 171.744
R1393 VDD2.n33 VDD2.n19 171.744
R1394 VDD2.n34 VDD2.n33 171.744
R1395 VDD2.n34 VDD2.n15 171.744
R1396 VDD2.n42 VDD2.n15 171.744
R1397 VDD2.n43 VDD2.n42 171.744
R1398 VDD2.n44 VDD2.n43 171.744
R1399 VDD2.n44 VDD2.n11 171.744
R1400 VDD2.n51 VDD2.n11 171.744
R1401 VDD2.n52 VDD2.n51 171.744
R1402 VDD2.n52 VDD2.n7 171.744
R1403 VDD2.n59 VDD2.n7 171.744
R1404 VDD2.n60 VDD2.n59 171.744
R1405 VDD2.n60 VDD2.n3 171.744
R1406 VDD2.n67 VDD2.n3 171.744
R1407 VDD2.n68 VDD2.n67 171.744
R1408 VDD2.n146 VDD2.n72 87.765
R1409 VDD2.n100 VDD2.t0 85.8723
R1410 VDD2.n25 VDD2.t1 85.8723
R1411 VDD2.n146 VDD2.n145 48.8641
R1412 VDD2.n87 VDD2.n85 13.1884
R1413 VDD2.n45 VDD2.n12 13.1884
R1414 VDD2.n123 VDD2.n122 12.8005
R1415 VDD2.n119 VDD2.n118 12.8005
R1416 VDD2.n46 VDD2.n14 12.8005
R1417 VDD2.n50 VDD2.n49 12.8005
R1418 VDD2.n126 VDD2.n83 12.0247
R1419 VDD2.n115 VDD2.n88 12.0247
R1420 VDD2.n41 VDD2.n40 12.0247
R1421 VDD2.n53 VDD2.n10 12.0247
R1422 VDD2.n127 VDD2.n81 11.249
R1423 VDD2.n114 VDD2.n91 11.249
R1424 VDD2.n39 VDD2.n16 11.249
R1425 VDD2.n54 VDD2.n8 11.249
R1426 VDD2.n99 VDD2.n98 10.7239
R1427 VDD2.n24 VDD2.n23 10.7239
R1428 VDD2.n131 VDD2.n130 10.4732
R1429 VDD2.n111 VDD2.n110 10.4732
R1430 VDD2.n36 VDD2.n35 10.4732
R1431 VDD2.n58 VDD2.n57 10.4732
R1432 VDD2.n134 VDD2.n79 9.69747
R1433 VDD2.n107 VDD2.n93 9.69747
R1434 VDD2.n32 VDD2.n18 9.69747
R1435 VDD2.n61 VDD2.n6 9.69747
R1436 VDD2.n145 VDD2.n144 9.45567
R1437 VDD2.n72 VDD2.n71 9.45567
R1438 VDD2.n97 VDD2.n96 9.3005
R1439 VDD2.n104 VDD2.n103 9.3005
R1440 VDD2.n106 VDD2.n105 9.3005
R1441 VDD2.n93 VDD2.n92 9.3005
R1442 VDD2.n112 VDD2.n111 9.3005
R1443 VDD2.n114 VDD2.n113 9.3005
R1444 VDD2.n88 VDD2.n86 9.3005
R1445 VDD2.n120 VDD2.n119 9.3005
R1446 VDD2.n144 VDD2.n143 9.3005
R1447 VDD2.n75 VDD2.n74 9.3005
R1448 VDD2.n138 VDD2.n137 9.3005
R1449 VDD2.n136 VDD2.n135 9.3005
R1450 VDD2.n79 VDD2.n78 9.3005
R1451 VDD2.n130 VDD2.n129 9.3005
R1452 VDD2.n128 VDD2.n127 9.3005
R1453 VDD2.n83 VDD2.n82 9.3005
R1454 VDD2.n122 VDD2.n121 9.3005
R1455 VDD2.n71 VDD2.n70 9.3005
R1456 VDD2.n65 VDD2.n64 9.3005
R1457 VDD2.n63 VDD2.n62 9.3005
R1458 VDD2.n6 VDD2.n5 9.3005
R1459 VDD2.n57 VDD2.n56 9.3005
R1460 VDD2.n55 VDD2.n54 9.3005
R1461 VDD2.n10 VDD2.n9 9.3005
R1462 VDD2.n49 VDD2.n48 9.3005
R1463 VDD2.n22 VDD2.n21 9.3005
R1464 VDD2.n29 VDD2.n28 9.3005
R1465 VDD2.n31 VDD2.n30 9.3005
R1466 VDD2.n18 VDD2.n17 9.3005
R1467 VDD2.n37 VDD2.n36 9.3005
R1468 VDD2.n39 VDD2.n38 9.3005
R1469 VDD2.n40 VDD2.n13 9.3005
R1470 VDD2.n47 VDD2.n46 9.3005
R1471 VDD2.n2 VDD2.n1 9.3005
R1472 VDD2.n135 VDD2.n77 8.92171
R1473 VDD2.n106 VDD2.n95 8.92171
R1474 VDD2.n31 VDD2.n20 8.92171
R1475 VDD2.n62 VDD2.n4 8.92171
R1476 VDD2.n139 VDD2.n138 8.14595
R1477 VDD2.n103 VDD2.n102 8.14595
R1478 VDD2.n28 VDD2.n27 8.14595
R1479 VDD2.n66 VDD2.n65 8.14595
R1480 VDD2.n145 VDD2.n73 7.3702
R1481 VDD2.n142 VDD2.n75 7.3702
R1482 VDD2.n99 VDD2.n97 7.3702
R1483 VDD2.n24 VDD2.n22 7.3702
R1484 VDD2.n69 VDD2.n2 7.3702
R1485 VDD2.n72 VDD2.n0 7.3702
R1486 VDD2.n143 VDD2.n73 6.59444
R1487 VDD2.n143 VDD2.n142 6.59444
R1488 VDD2.n70 VDD2.n69 6.59444
R1489 VDD2.n70 VDD2.n0 6.59444
R1490 VDD2.n139 VDD2.n75 5.81868
R1491 VDD2.n102 VDD2.n97 5.81868
R1492 VDD2.n27 VDD2.n22 5.81868
R1493 VDD2.n66 VDD2.n2 5.81868
R1494 VDD2.n138 VDD2.n77 5.04292
R1495 VDD2.n103 VDD2.n95 5.04292
R1496 VDD2.n28 VDD2.n20 5.04292
R1497 VDD2.n65 VDD2.n4 5.04292
R1498 VDD2.n135 VDD2.n134 4.26717
R1499 VDD2.n107 VDD2.n106 4.26717
R1500 VDD2.n32 VDD2.n31 4.26717
R1501 VDD2.n62 VDD2.n61 4.26717
R1502 VDD2.n131 VDD2.n79 3.49141
R1503 VDD2.n110 VDD2.n93 3.49141
R1504 VDD2.n35 VDD2.n18 3.49141
R1505 VDD2.n58 VDD2.n6 3.49141
R1506 VDD2.n130 VDD2.n81 2.71565
R1507 VDD2.n111 VDD2.n91 2.71565
R1508 VDD2.n36 VDD2.n16 2.71565
R1509 VDD2.n57 VDD2.n8 2.71565
R1510 VDD2.n98 VDD2.n96 2.41282
R1511 VDD2.n23 VDD2.n21 2.41282
R1512 VDD2.n127 VDD2.n126 1.93989
R1513 VDD2.n115 VDD2.n114 1.93989
R1514 VDD2.n41 VDD2.n39 1.93989
R1515 VDD2.n54 VDD2.n53 1.93989
R1516 VDD2.n123 VDD2.n83 1.16414
R1517 VDD2.n118 VDD2.n88 1.16414
R1518 VDD2.n40 VDD2.n14 1.16414
R1519 VDD2.n50 VDD2.n10 1.16414
R1520 VDD2 VDD2.n146 0.502655
R1521 VDD2.n122 VDD2.n85 0.388379
R1522 VDD2.n119 VDD2.n87 0.388379
R1523 VDD2.n46 VDD2.n45 0.388379
R1524 VDD2.n49 VDD2.n12 0.388379
R1525 VDD2.n144 VDD2.n74 0.155672
R1526 VDD2.n137 VDD2.n74 0.155672
R1527 VDD2.n137 VDD2.n136 0.155672
R1528 VDD2.n136 VDD2.n78 0.155672
R1529 VDD2.n129 VDD2.n78 0.155672
R1530 VDD2.n129 VDD2.n128 0.155672
R1531 VDD2.n128 VDD2.n82 0.155672
R1532 VDD2.n121 VDD2.n82 0.155672
R1533 VDD2.n121 VDD2.n120 0.155672
R1534 VDD2.n120 VDD2.n86 0.155672
R1535 VDD2.n113 VDD2.n86 0.155672
R1536 VDD2.n113 VDD2.n112 0.155672
R1537 VDD2.n112 VDD2.n92 0.155672
R1538 VDD2.n105 VDD2.n92 0.155672
R1539 VDD2.n105 VDD2.n104 0.155672
R1540 VDD2.n104 VDD2.n96 0.155672
R1541 VDD2.n29 VDD2.n21 0.155672
R1542 VDD2.n30 VDD2.n29 0.155672
R1543 VDD2.n30 VDD2.n17 0.155672
R1544 VDD2.n37 VDD2.n17 0.155672
R1545 VDD2.n38 VDD2.n37 0.155672
R1546 VDD2.n38 VDD2.n13 0.155672
R1547 VDD2.n47 VDD2.n13 0.155672
R1548 VDD2.n48 VDD2.n47 0.155672
R1549 VDD2.n48 VDD2.n9 0.155672
R1550 VDD2.n55 VDD2.n9 0.155672
R1551 VDD2.n56 VDD2.n55 0.155672
R1552 VDD2.n56 VDD2.n5 0.155672
R1553 VDD2.n63 VDD2.n5 0.155672
R1554 VDD2.n64 VDD2.n63 0.155672
R1555 VDD2.n64 VDD2.n1 0.155672
R1556 VDD2.n71 VDD2.n1 0.155672
R1557 VP.n0 VP.t0 291.267
R1558 VP.n0 VP.t1 247.736
R1559 VP VP.n0 0.241678
R1560 VDD1.n68 VDD1.n0 756.745
R1561 VDD1.n141 VDD1.n73 756.745
R1562 VDD1.n69 VDD1.n68 585
R1563 VDD1.n67 VDD1.n66 585
R1564 VDD1.n4 VDD1.n3 585
R1565 VDD1.n61 VDD1.n60 585
R1566 VDD1.n59 VDD1.n58 585
R1567 VDD1.n8 VDD1.n7 585
R1568 VDD1.n53 VDD1.n52 585
R1569 VDD1.n51 VDD1.n50 585
R1570 VDD1.n12 VDD1.n11 585
R1571 VDD1.n16 VDD1.n14 585
R1572 VDD1.n45 VDD1.n44 585
R1573 VDD1.n43 VDD1.n42 585
R1574 VDD1.n18 VDD1.n17 585
R1575 VDD1.n37 VDD1.n36 585
R1576 VDD1.n35 VDD1.n34 585
R1577 VDD1.n22 VDD1.n21 585
R1578 VDD1.n29 VDD1.n28 585
R1579 VDD1.n27 VDD1.n26 585
R1580 VDD1.n98 VDD1.n97 585
R1581 VDD1.n100 VDD1.n99 585
R1582 VDD1.n93 VDD1.n92 585
R1583 VDD1.n106 VDD1.n105 585
R1584 VDD1.n108 VDD1.n107 585
R1585 VDD1.n89 VDD1.n88 585
R1586 VDD1.n115 VDD1.n114 585
R1587 VDD1.n116 VDD1.n87 585
R1588 VDD1.n118 VDD1.n117 585
R1589 VDD1.n85 VDD1.n84 585
R1590 VDD1.n124 VDD1.n123 585
R1591 VDD1.n126 VDD1.n125 585
R1592 VDD1.n81 VDD1.n80 585
R1593 VDD1.n132 VDD1.n131 585
R1594 VDD1.n134 VDD1.n133 585
R1595 VDD1.n77 VDD1.n76 585
R1596 VDD1.n140 VDD1.n139 585
R1597 VDD1.n142 VDD1.n141 585
R1598 VDD1.n25 VDD1.t1 329.036
R1599 VDD1.n96 VDD1.t0 329.036
R1600 VDD1.n68 VDD1.n67 171.744
R1601 VDD1.n67 VDD1.n3 171.744
R1602 VDD1.n60 VDD1.n3 171.744
R1603 VDD1.n60 VDD1.n59 171.744
R1604 VDD1.n59 VDD1.n7 171.744
R1605 VDD1.n52 VDD1.n7 171.744
R1606 VDD1.n52 VDD1.n51 171.744
R1607 VDD1.n51 VDD1.n11 171.744
R1608 VDD1.n16 VDD1.n11 171.744
R1609 VDD1.n44 VDD1.n16 171.744
R1610 VDD1.n44 VDD1.n43 171.744
R1611 VDD1.n43 VDD1.n17 171.744
R1612 VDD1.n36 VDD1.n17 171.744
R1613 VDD1.n36 VDD1.n35 171.744
R1614 VDD1.n35 VDD1.n21 171.744
R1615 VDD1.n28 VDD1.n21 171.744
R1616 VDD1.n28 VDD1.n27 171.744
R1617 VDD1.n99 VDD1.n98 171.744
R1618 VDD1.n99 VDD1.n92 171.744
R1619 VDD1.n106 VDD1.n92 171.744
R1620 VDD1.n107 VDD1.n106 171.744
R1621 VDD1.n107 VDD1.n88 171.744
R1622 VDD1.n115 VDD1.n88 171.744
R1623 VDD1.n116 VDD1.n115 171.744
R1624 VDD1.n117 VDD1.n116 171.744
R1625 VDD1.n117 VDD1.n84 171.744
R1626 VDD1.n124 VDD1.n84 171.744
R1627 VDD1.n125 VDD1.n124 171.744
R1628 VDD1.n125 VDD1.n80 171.744
R1629 VDD1.n132 VDD1.n80 171.744
R1630 VDD1.n133 VDD1.n132 171.744
R1631 VDD1.n133 VDD1.n76 171.744
R1632 VDD1.n140 VDD1.n76 171.744
R1633 VDD1.n141 VDD1.n140 171.744
R1634 VDD1 VDD1.n145 88.7338
R1635 VDD1.n27 VDD1.t1 85.8723
R1636 VDD1.n98 VDD1.t0 85.8723
R1637 VDD1 VDD1.n72 49.3663
R1638 VDD1.n14 VDD1.n12 13.1884
R1639 VDD1.n118 VDD1.n85 13.1884
R1640 VDD1.n50 VDD1.n49 12.8005
R1641 VDD1.n46 VDD1.n45 12.8005
R1642 VDD1.n119 VDD1.n87 12.8005
R1643 VDD1.n123 VDD1.n122 12.8005
R1644 VDD1.n53 VDD1.n10 12.0247
R1645 VDD1.n42 VDD1.n15 12.0247
R1646 VDD1.n114 VDD1.n113 12.0247
R1647 VDD1.n126 VDD1.n83 12.0247
R1648 VDD1.n54 VDD1.n8 11.249
R1649 VDD1.n41 VDD1.n18 11.249
R1650 VDD1.n112 VDD1.n89 11.249
R1651 VDD1.n127 VDD1.n81 11.249
R1652 VDD1.n26 VDD1.n25 10.7239
R1653 VDD1.n97 VDD1.n96 10.7239
R1654 VDD1.n58 VDD1.n57 10.4732
R1655 VDD1.n38 VDD1.n37 10.4732
R1656 VDD1.n109 VDD1.n108 10.4732
R1657 VDD1.n131 VDD1.n130 10.4732
R1658 VDD1.n61 VDD1.n6 9.69747
R1659 VDD1.n34 VDD1.n20 9.69747
R1660 VDD1.n105 VDD1.n91 9.69747
R1661 VDD1.n134 VDD1.n79 9.69747
R1662 VDD1.n72 VDD1.n71 9.45567
R1663 VDD1.n145 VDD1.n144 9.45567
R1664 VDD1.n24 VDD1.n23 9.3005
R1665 VDD1.n31 VDD1.n30 9.3005
R1666 VDD1.n33 VDD1.n32 9.3005
R1667 VDD1.n20 VDD1.n19 9.3005
R1668 VDD1.n39 VDD1.n38 9.3005
R1669 VDD1.n41 VDD1.n40 9.3005
R1670 VDD1.n15 VDD1.n13 9.3005
R1671 VDD1.n47 VDD1.n46 9.3005
R1672 VDD1.n71 VDD1.n70 9.3005
R1673 VDD1.n2 VDD1.n1 9.3005
R1674 VDD1.n65 VDD1.n64 9.3005
R1675 VDD1.n63 VDD1.n62 9.3005
R1676 VDD1.n6 VDD1.n5 9.3005
R1677 VDD1.n57 VDD1.n56 9.3005
R1678 VDD1.n55 VDD1.n54 9.3005
R1679 VDD1.n10 VDD1.n9 9.3005
R1680 VDD1.n49 VDD1.n48 9.3005
R1681 VDD1.n144 VDD1.n143 9.3005
R1682 VDD1.n138 VDD1.n137 9.3005
R1683 VDD1.n136 VDD1.n135 9.3005
R1684 VDD1.n79 VDD1.n78 9.3005
R1685 VDD1.n130 VDD1.n129 9.3005
R1686 VDD1.n128 VDD1.n127 9.3005
R1687 VDD1.n83 VDD1.n82 9.3005
R1688 VDD1.n122 VDD1.n121 9.3005
R1689 VDD1.n95 VDD1.n94 9.3005
R1690 VDD1.n102 VDD1.n101 9.3005
R1691 VDD1.n104 VDD1.n103 9.3005
R1692 VDD1.n91 VDD1.n90 9.3005
R1693 VDD1.n110 VDD1.n109 9.3005
R1694 VDD1.n112 VDD1.n111 9.3005
R1695 VDD1.n113 VDD1.n86 9.3005
R1696 VDD1.n120 VDD1.n119 9.3005
R1697 VDD1.n75 VDD1.n74 9.3005
R1698 VDD1.n62 VDD1.n4 8.92171
R1699 VDD1.n33 VDD1.n22 8.92171
R1700 VDD1.n104 VDD1.n93 8.92171
R1701 VDD1.n135 VDD1.n77 8.92171
R1702 VDD1.n66 VDD1.n65 8.14595
R1703 VDD1.n30 VDD1.n29 8.14595
R1704 VDD1.n101 VDD1.n100 8.14595
R1705 VDD1.n139 VDD1.n138 8.14595
R1706 VDD1.n72 VDD1.n0 7.3702
R1707 VDD1.n69 VDD1.n2 7.3702
R1708 VDD1.n26 VDD1.n24 7.3702
R1709 VDD1.n97 VDD1.n95 7.3702
R1710 VDD1.n142 VDD1.n75 7.3702
R1711 VDD1.n145 VDD1.n73 7.3702
R1712 VDD1.n70 VDD1.n0 6.59444
R1713 VDD1.n70 VDD1.n69 6.59444
R1714 VDD1.n143 VDD1.n142 6.59444
R1715 VDD1.n143 VDD1.n73 6.59444
R1716 VDD1.n66 VDD1.n2 5.81868
R1717 VDD1.n29 VDD1.n24 5.81868
R1718 VDD1.n100 VDD1.n95 5.81868
R1719 VDD1.n139 VDD1.n75 5.81868
R1720 VDD1.n65 VDD1.n4 5.04292
R1721 VDD1.n30 VDD1.n22 5.04292
R1722 VDD1.n101 VDD1.n93 5.04292
R1723 VDD1.n138 VDD1.n77 5.04292
R1724 VDD1.n62 VDD1.n61 4.26717
R1725 VDD1.n34 VDD1.n33 4.26717
R1726 VDD1.n105 VDD1.n104 4.26717
R1727 VDD1.n135 VDD1.n134 4.26717
R1728 VDD1.n58 VDD1.n6 3.49141
R1729 VDD1.n37 VDD1.n20 3.49141
R1730 VDD1.n108 VDD1.n91 3.49141
R1731 VDD1.n131 VDD1.n79 3.49141
R1732 VDD1.n57 VDD1.n8 2.71565
R1733 VDD1.n38 VDD1.n18 2.71565
R1734 VDD1.n109 VDD1.n89 2.71565
R1735 VDD1.n130 VDD1.n81 2.71565
R1736 VDD1.n25 VDD1.n23 2.41282
R1737 VDD1.n96 VDD1.n94 2.41282
R1738 VDD1.n54 VDD1.n53 1.93989
R1739 VDD1.n42 VDD1.n41 1.93989
R1740 VDD1.n114 VDD1.n112 1.93989
R1741 VDD1.n127 VDD1.n126 1.93989
R1742 VDD1.n50 VDD1.n10 1.16414
R1743 VDD1.n45 VDD1.n15 1.16414
R1744 VDD1.n113 VDD1.n87 1.16414
R1745 VDD1.n123 VDD1.n83 1.16414
R1746 VDD1.n49 VDD1.n12 0.388379
R1747 VDD1.n46 VDD1.n14 0.388379
R1748 VDD1.n119 VDD1.n118 0.388379
R1749 VDD1.n122 VDD1.n85 0.388379
R1750 VDD1.n71 VDD1.n1 0.155672
R1751 VDD1.n64 VDD1.n1 0.155672
R1752 VDD1.n64 VDD1.n63 0.155672
R1753 VDD1.n63 VDD1.n5 0.155672
R1754 VDD1.n56 VDD1.n5 0.155672
R1755 VDD1.n56 VDD1.n55 0.155672
R1756 VDD1.n55 VDD1.n9 0.155672
R1757 VDD1.n48 VDD1.n9 0.155672
R1758 VDD1.n48 VDD1.n47 0.155672
R1759 VDD1.n47 VDD1.n13 0.155672
R1760 VDD1.n40 VDD1.n13 0.155672
R1761 VDD1.n40 VDD1.n39 0.155672
R1762 VDD1.n39 VDD1.n19 0.155672
R1763 VDD1.n32 VDD1.n19 0.155672
R1764 VDD1.n32 VDD1.n31 0.155672
R1765 VDD1.n31 VDD1.n23 0.155672
R1766 VDD1.n102 VDD1.n94 0.155672
R1767 VDD1.n103 VDD1.n102 0.155672
R1768 VDD1.n103 VDD1.n90 0.155672
R1769 VDD1.n110 VDD1.n90 0.155672
R1770 VDD1.n111 VDD1.n110 0.155672
R1771 VDD1.n111 VDD1.n86 0.155672
R1772 VDD1.n120 VDD1.n86 0.155672
R1773 VDD1.n121 VDD1.n120 0.155672
R1774 VDD1.n121 VDD1.n82 0.155672
R1775 VDD1.n128 VDD1.n82 0.155672
R1776 VDD1.n129 VDD1.n128 0.155672
R1777 VDD1.n129 VDD1.n78 0.155672
R1778 VDD1.n136 VDD1.n78 0.155672
R1779 VDD1.n137 VDD1.n136 0.155672
R1780 VDD1.n137 VDD1.n74 0.155672
R1781 VDD1.n144 VDD1.n74 0.155672
C0 w_n1794_n3680# VN 2.43932f
C1 w_n1794_n3680# VDD1 1.79464f
C2 VDD1 VN 0.147389f
C3 w_n1794_n3680# VDD2 1.81007f
C4 VDD2 VN 2.88443f
C5 VDD1 VDD2 0.572445f
C6 VTAIL B 3.5964f
C7 VTAIL VP 2.43644f
C8 B VP 1.28725f
C9 w_n1794_n3680# VTAIL 3.0141f
C10 VTAIL VN 2.42203f
C11 VTAIL VDD1 5.47729f
C12 VTAIL VDD2 5.52033f
C13 w_n1794_n3680# B 8.30617f
C14 B VN 0.918123f
C15 w_n1794_n3680# VP 2.66597f
C16 B VDD1 1.70332f
C17 VN VP 5.34103f
C18 B VDD2 1.72571f
C19 VDD1 VP 3.03f
C20 VDD2 VP 0.296435f
C21 VDD2 VSUBS 0.870059f
C22 VDD1 VSUBS 3.58192f
C23 VTAIL VSUBS 0.964255f
C24 VN VSUBS 8.03138f
C25 VP VSUBS 1.489623f
C26 B VSUBS 3.38066f
C27 w_n1794_n3680# VSUBS 81.096f
C28 VDD1.n0 VSUBS 0.022758f
C29 VDD1.n1 VSUBS 0.020166f
C30 VDD1.n2 VSUBS 0.010836f
C31 VDD1.n3 VSUBS 0.025613f
C32 VDD1.n4 VSUBS 0.011474f
C33 VDD1.n5 VSUBS 0.020166f
C34 VDD1.n6 VSUBS 0.010836f
C35 VDD1.n7 VSUBS 0.025613f
C36 VDD1.n8 VSUBS 0.011474f
C37 VDD1.n9 VSUBS 0.020166f
C38 VDD1.n10 VSUBS 0.010836f
C39 VDD1.n11 VSUBS 0.025613f
C40 VDD1.n12 VSUBS 0.011155f
C41 VDD1.n13 VSUBS 0.020166f
C42 VDD1.n14 VSUBS 0.011155f
C43 VDD1.n15 VSUBS 0.010836f
C44 VDD1.n16 VSUBS 0.025613f
C45 VDD1.n17 VSUBS 0.025613f
C46 VDD1.n18 VSUBS 0.011474f
C47 VDD1.n19 VSUBS 0.020166f
C48 VDD1.n20 VSUBS 0.010836f
C49 VDD1.n21 VSUBS 0.025613f
C50 VDD1.n22 VSUBS 0.011474f
C51 VDD1.n23 VSUBS 1.12866f
C52 VDD1.n24 VSUBS 0.010836f
C53 VDD1.t1 VSUBS 0.055298f
C54 VDD1.n25 VSUBS 0.173042f
C55 VDD1.n26 VSUBS 0.019267f
C56 VDD1.n27 VSUBS 0.01921f
C57 VDD1.n28 VSUBS 0.025613f
C58 VDD1.n29 VSUBS 0.011474f
C59 VDD1.n30 VSUBS 0.010836f
C60 VDD1.n31 VSUBS 0.020166f
C61 VDD1.n32 VSUBS 0.020166f
C62 VDD1.n33 VSUBS 0.010836f
C63 VDD1.n34 VSUBS 0.011474f
C64 VDD1.n35 VSUBS 0.025613f
C65 VDD1.n36 VSUBS 0.025613f
C66 VDD1.n37 VSUBS 0.011474f
C67 VDD1.n38 VSUBS 0.010836f
C68 VDD1.n39 VSUBS 0.020166f
C69 VDD1.n40 VSUBS 0.020166f
C70 VDD1.n41 VSUBS 0.010836f
C71 VDD1.n42 VSUBS 0.011474f
C72 VDD1.n43 VSUBS 0.025613f
C73 VDD1.n44 VSUBS 0.025613f
C74 VDD1.n45 VSUBS 0.011474f
C75 VDD1.n46 VSUBS 0.010836f
C76 VDD1.n47 VSUBS 0.020166f
C77 VDD1.n48 VSUBS 0.020166f
C78 VDD1.n49 VSUBS 0.010836f
C79 VDD1.n50 VSUBS 0.011474f
C80 VDD1.n51 VSUBS 0.025613f
C81 VDD1.n52 VSUBS 0.025613f
C82 VDD1.n53 VSUBS 0.011474f
C83 VDD1.n54 VSUBS 0.010836f
C84 VDD1.n55 VSUBS 0.020166f
C85 VDD1.n56 VSUBS 0.020166f
C86 VDD1.n57 VSUBS 0.010836f
C87 VDD1.n58 VSUBS 0.011474f
C88 VDD1.n59 VSUBS 0.025613f
C89 VDD1.n60 VSUBS 0.025613f
C90 VDD1.n61 VSUBS 0.011474f
C91 VDD1.n62 VSUBS 0.010836f
C92 VDD1.n63 VSUBS 0.020166f
C93 VDD1.n64 VSUBS 0.020166f
C94 VDD1.n65 VSUBS 0.010836f
C95 VDD1.n66 VSUBS 0.011474f
C96 VDD1.n67 VSUBS 0.025613f
C97 VDD1.n68 VSUBS 0.064049f
C98 VDD1.n69 VSUBS 0.011474f
C99 VDD1.n70 VSUBS 0.010836f
C100 VDD1.n71 VSUBS 0.046613f
C101 VDD1.n72 VSUBS 0.046951f
C102 VDD1.n73 VSUBS 0.022758f
C103 VDD1.n74 VSUBS 0.020166f
C104 VDD1.n75 VSUBS 0.010836f
C105 VDD1.n76 VSUBS 0.025613f
C106 VDD1.n77 VSUBS 0.011474f
C107 VDD1.n78 VSUBS 0.020166f
C108 VDD1.n79 VSUBS 0.010836f
C109 VDD1.n80 VSUBS 0.025613f
C110 VDD1.n81 VSUBS 0.011474f
C111 VDD1.n82 VSUBS 0.020166f
C112 VDD1.n83 VSUBS 0.010836f
C113 VDD1.n84 VSUBS 0.025613f
C114 VDD1.n85 VSUBS 0.011155f
C115 VDD1.n86 VSUBS 0.020166f
C116 VDD1.n87 VSUBS 0.011474f
C117 VDD1.n88 VSUBS 0.025613f
C118 VDD1.n89 VSUBS 0.011474f
C119 VDD1.n90 VSUBS 0.020166f
C120 VDD1.n91 VSUBS 0.010836f
C121 VDD1.n92 VSUBS 0.025613f
C122 VDD1.n93 VSUBS 0.011474f
C123 VDD1.n94 VSUBS 1.12866f
C124 VDD1.n95 VSUBS 0.010836f
C125 VDD1.t0 VSUBS 0.055298f
C126 VDD1.n96 VSUBS 0.173042f
C127 VDD1.n97 VSUBS 0.019267f
C128 VDD1.n98 VSUBS 0.01921f
C129 VDD1.n99 VSUBS 0.025613f
C130 VDD1.n100 VSUBS 0.011474f
C131 VDD1.n101 VSUBS 0.010836f
C132 VDD1.n102 VSUBS 0.020166f
C133 VDD1.n103 VSUBS 0.020166f
C134 VDD1.n104 VSUBS 0.010836f
C135 VDD1.n105 VSUBS 0.011474f
C136 VDD1.n106 VSUBS 0.025613f
C137 VDD1.n107 VSUBS 0.025613f
C138 VDD1.n108 VSUBS 0.011474f
C139 VDD1.n109 VSUBS 0.010836f
C140 VDD1.n110 VSUBS 0.020166f
C141 VDD1.n111 VSUBS 0.020166f
C142 VDD1.n112 VSUBS 0.010836f
C143 VDD1.n113 VSUBS 0.010836f
C144 VDD1.n114 VSUBS 0.011474f
C145 VDD1.n115 VSUBS 0.025613f
C146 VDD1.n116 VSUBS 0.025613f
C147 VDD1.n117 VSUBS 0.025613f
C148 VDD1.n118 VSUBS 0.011155f
C149 VDD1.n119 VSUBS 0.010836f
C150 VDD1.n120 VSUBS 0.020166f
C151 VDD1.n121 VSUBS 0.020166f
C152 VDD1.n122 VSUBS 0.010836f
C153 VDD1.n123 VSUBS 0.011474f
C154 VDD1.n124 VSUBS 0.025613f
C155 VDD1.n125 VSUBS 0.025613f
C156 VDD1.n126 VSUBS 0.011474f
C157 VDD1.n127 VSUBS 0.010836f
C158 VDD1.n128 VSUBS 0.020166f
C159 VDD1.n129 VSUBS 0.020166f
C160 VDD1.n130 VSUBS 0.010836f
C161 VDD1.n131 VSUBS 0.011474f
C162 VDD1.n132 VSUBS 0.025613f
C163 VDD1.n133 VSUBS 0.025613f
C164 VDD1.n134 VSUBS 0.011474f
C165 VDD1.n135 VSUBS 0.010836f
C166 VDD1.n136 VSUBS 0.020166f
C167 VDD1.n137 VSUBS 0.020166f
C168 VDD1.n138 VSUBS 0.010836f
C169 VDD1.n139 VSUBS 0.011474f
C170 VDD1.n140 VSUBS 0.025613f
C171 VDD1.n141 VSUBS 0.064049f
C172 VDD1.n142 VSUBS 0.011474f
C173 VDD1.n143 VSUBS 0.010836f
C174 VDD1.n144 VSUBS 0.046613f
C175 VDD1.n145 VSUBS 0.62728f
C176 VP.t0 VSUBS 3.914f
C177 VP.t1 VSUBS 3.42795f
C178 VP.n0 VSUBS 5.98701f
C179 VDD2.n0 VSUBS 0.022689f
C180 VDD2.n1 VSUBS 0.020105f
C181 VDD2.n2 VSUBS 0.010804f
C182 VDD2.n3 VSUBS 0.025535f
C183 VDD2.n4 VSUBS 0.011439f
C184 VDD2.n5 VSUBS 0.020105f
C185 VDD2.n6 VSUBS 0.010804f
C186 VDD2.n7 VSUBS 0.025535f
C187 VDD2.n8 VSUBS 0.011439f
C188 VDD2.n9 VSUBS 0.020105f
C189 VDD2.n10 VSUBS 0.010804f
C190 VDD2.n11 VSUBS 0.025535f
C191 VDD2.n12 VSUBS 0.011121f
C192 VDD2.n13 VSUBS 0.020105f
C193 VDD2.n14 VSUBS 0.011439f
C194 VDD2.n15 VSUBS 0.025535f
C195 VDD2.n16 VSUBS 0.011439f
C196 VDD2.n17 VSUBS 0.020105f
C197 VDD2.n18 VSUBS 0.010804f
C198 VDD2.n19 VSUBS 0.025535f
C199 VDD2.n20 VSUBS 0.011439f
C200 VDD2.n21 VSUBS 1.12524f
C201 VDD2.n22 VSUBS 0.010804f
C202 VDD2.t1 VSUBS 0.05513f
C203 VDD2.n23 VSUBS 0.172518f
C204 VDD2.n24 VSUBS 0.019209f
C205 VDD2.n25 VSUBS 0.019152f
C206 VDD2.n26 VSUBS 0.025535f
C207 VDD2.n27 VSUBS 0.011439f
C208 VDD2.n28 VSUBS 0.010804f
C209 VDD2.n29 VSUBS 0.020105f
C210 VDD2.n30 VSUBS 0.020105f
C211 VDD2.n31 VSUBS 0.010804f
C212 VDD2.n32 VSUBS 0.011439f
C213 VDD2.n33 VSUBS 0.025535f
C214 VDD2.n34 VSUBS 0.025535f
C215 VDD2.n35 VSUBS 0.011439f
C216 VDD2.n36 VSUBS 0.010804f
C217 VDD2.n37 VSUBS 0.020105f
C218 VDD2.n38 VSUBS 0.020105f
C219 VDD2.n39 VSUBS 0.010804f
C220 VDD2.n40 VSUBS 0.010804f
C221 VDD2.n41 VSUBS 0.011439f
C222 VDD2.n42 VSUBS 0.025535f
C223 VDD2.n43 VSUBS 0.025535f
C224 VDD2.n44 VSUBS 0.025535f
C225 VDD2.n45 VSUBS 0.011121f
C226 VDD2.n46 VSUBS 0.010804f
C227 VDD2.n47 VSUBS 0.020105f
C228 VDD2.n48 VSUBS 0.020105f
C229 VDD2.n49 VSUBS 0.010804f
C230 VDD2.n50 VSUBS 0.011439f
C231 VDD2.n51 VSUBS 0.025535f
C232 VDD2.n52 VSUBS 0.025535f
C233 VDD2.n53 VSUBS 0.011439f
C234 VDD2.n54 VSUBS 0.010804f
C235 VDD2.n55 VSUBS 0.020105f
C236 VDD2.n56 VSUBS 0.020105f
C237 VDD2.n57 VSUBS 0.010804f
C238 VDD2.n58 VSUBS 0.011439f
C239 VDD2.n59 VSUBS 0.025535f
C240 VDD2.n60 VSUBS 0.025535f
C241 VDD2.n61 VSUBS 0.011439f
C242 VDD2.n62 VSUBS 0.010804f
C243 VDD2.n63 VSUBS 0.020105f
C244 VDD2.n64 VSUBS 0.020105f
C245 VDD2.n65 VSUBS 0.010804f
C246 VDD2.n66 VSUBS 0.011439f
C247 VDD2.n67 VSUBS 0.025535f
C248 VDD2.n68 VSUBS 0.063855f
C249 VDD2.n69 VSUBS 0.011439f
C250 VDD2.n70 VSUBS 0.010804f
C251 VDD2.n71 VSUBS 0.046471f
C252 VDD2.n72 VSUBS 0.591031f
C253 VDD2.n73 VSUBS 0.022689f
C254 VDD2.n74 VSUBS 0.020105f
C255 VDD2.n75 VSUBS 0.010804f
C256 VDD2.n76 VSUBS 0.025535f
C257 VDD2.n77 VSUBS 0.011439f
C258 VDD2.n78 VSUBS 0.020105f
C259 VDD2.n79 VSUBS 0.010804f
C260 VDD2.n80 VSUBS 0.025535f
C261 VDD2.n81 VSUBS 0.011439f
C262 VDD2.n82 VSUBS 0.020105f
C263 VDD2.n83 VSUBS 0.010804f
C264 VDD2.n84 VSUBS 0.025535f
C265 VDD2.n85 VSUBS 0.011121f
C266 VDD2.n86 VSUBS 0.020105f
C267 VDD2.n87 VSUBS 0.011121f
C268 VDD2.n88 VSUBS 0.010804f
C269 VDD2.n89 VSUBS 0.025535f
C270 VDD2.n90 VSUBS 0.025535f
C271 VDD2.n91 VSUBS 0.011439f
C272 VDD2.n92 VSUBS 0.020105f
C273 VDD2.n93 VSUBS 0.010804f
C274 VDD2.n94 VSUBS 0.025535f
C275 VDD2.n95 VSUBS 0.011439f
C276 VDD2.n96 VSUBS 1.12524f
C277 VDD2.n97 VSUBS 0.010804f
C278 VDD2.t0 VSUBS 0.05513f
C279 VDD2.n98 VSUBS 0.172518f
C280 VDD2.n99 VSUBS 0.019209f
C281 VDD2.n100 VSUBS 0.019152f
C282 VDD2.n101 VSUBS 0.025535f
C283 VDD2.n102 VSUBS 0.011439f
C284 VDD2.n103 VSUBS 0.010804f
C285 VDD2.n104 VSUBS 0.020105f
C286 VDD2.n105 VSUBS 0.020105f
C287 VDD2.n106 VSUBS 0.010804f
C288 VDD2.n107 VSUBS 0.011439f
C289 VDD2.n108 VSUBS 0.025535f
C290 VDD2.n109 VSUBS 0.025535f
C291 VDD2.n110 VSUBS 0.011439f
C292 VDD2.n111 VSUBS 0.010804f
C293 VDD2.n112 VSUBS 0.020105f
C294 VDD2.n113 VSUBS 0.020105f
C295 VDD2.n114 VSUBS 0.010804f
C296 VDD2.n115 VSUBS 0.011439f
C297 VDD2.n116 VSUBS 0.025535f
C298 VDD2.n117 VSUBS 0.025535f
C299 VDD2.n118 VSUBS 0.011439f
C300 VDD2.n119 VSUBS 0.010804f
C301 VDD2.n120 VSUBS 0.020105f
C302 VDD2.n121 VSUBS 0.020105f
C303 VDD2.n122 VSUBS 0.010804f
C304 VDD2.n123 VSUBS 0.011439f
C305 VDD2.n124 VSUBS 0.025535f
C306 VDD2.n125 VSUBS 0.025535f
C307 VDD2.n126 VSUBS 0.011439f
C308 VDD2.n127 VSUBS 0.010804f
C309 VDD2.n128 VSUBS 0.020105f
C310 VDD2.n129 VSUBS 0.020105f
C311 VDD2.n130 VSUBS 0.010804f
C312 VDD2.n131 VSUBS 0.011439f
C313 VDD2.n132 VSUBS 0.025535f
C314 VDD2.n133 VSUBS 0.025535f
C315 VDD2.n134 VSUBS 0.011439f
C316 VDD2.n135 VSUBS 0.010804f
C317 VDD2.n136 VSUBS 0.020105f
C318 VDD2.n137 VSUBS 0.020105f
C319 VDD2.n138 VSUBS 0.010804f
C320 VDD2.n139 VSUBS 0.011439f
C321 VDD2.n140 VSUBS 0.025535f
C322 VDD2.n141 VSUBS 0.063855f
C323 VDD2.n142 VSUBS 0.011439f
C324 VDD2.n143 VSUBS 0.010804f
C325 VDD2.n144 VSUBS 0.046471f
C326 VDD2.n145 VSUBS 0.046084f
C327 VDD2.n146 VSUBS 2.44848f
C328 VTAIL.n0 VSUBS 0.032148f
C329 VTAIL.n1 VSUBS 0.028487f
C330 VTAIL.n2 VSUBS 0.015308f
C331 VTAIL.n3 VSUBS 0.036182f
C332 VTAIL.n4 VSUBS 0.016208f
C333 VTAIL.n5 VSUBS 0.028487f
C334 VTAIL.n6 VSUBS 0.015308f
C335 VTAIL.n7 VSUBS 0.036182f
C336 VTAIL.n8 VSUBS 0.016208f
C337 VTAIL.n9 VSUBS 0.028487f
C338 VTAIL.n10 VSUBS 0.015308f
C339 VTAIL.n11 VSUBS 0.036182f
C340 VTAIL.n12 VSUBS 0.015758f
C341 VTAIL.n13 VSUBS 0.028487f
C342 VTAIL.n14 VSUBS 0.016208f
C343 VTAIL.n15 VSUBS 0.036182f
C344 VTAIL.n16 VSUBS 0.016208f
C345 VTAIL.n17 VSUBS 0.028487f
C346 VTAIL.n18 VSUBS 0.015308f
C347 VTAIL.n19 VSUBS 0.036182f
C348 VTAIL.n20 VSUBS 0.016208f
C349 VTAIL.n21 VSUBS 1.5944f
C350 VTAIL.n22 VSUBS 0.015308f
C351 VTAIL.t1 VSUBS 0.078116f
C352 VTAIL.n23 VSUBS 0.244447f
C353 VTAIL.n24 VSUBS 0.027218f
C354 VTAIL.n25 VSUBS 0.027137f
C355 VTAIL.n26 VSUBS 0.036182f
C356 VTAIL.n27 VSUBS 0.016208f
C357 VTAIL.n28 VSUBS 0.015308f
C358 VTAIL.n29 VSUBS 0.028487f
C359 VTAIL.n30 VSUBS 0.028487f
C360 VTAIL.n31 VSUBS 0.015308f
C361 VTAIL.n32 VSUBS 0.016208f
C362 VTAIL.n33 VSUBS 0.036182f
C363 VTAIL.n34 VSUBS 0.036182f
C364 VTAIL.n35 VSUBS 0.016208f
C365 VTAIL.n36 VSUBS 0.015308f
C366 VTAIL.n37 VSUBS 0.028487f
C367 VTAIL.n38 VSUBS 0.028487f
C368 VTAIL.n39 VSUBS 0.015308f
C369 VTAIL.n40 VSUBS 0.015308f
C370 VTAIL.n41 VSUBS 0.016208f
C371 VTAIL.n42 VSUBS 0.036182f
C372 VTAIL.n43 VSUBS 0.036182f
C373 VTAIL.n44 VSUBS 0.036182f
C374 VTAIL.n45 VSUBS 0.015758f
C375 VTAIL.n46 VSUBS 0.015308f
C376 VTAIL.n47 VSUBS 0.028487f
C377 VTAIL.n48 VSUBS 0.028487f
C378 VTAIL.n49 VSUBS 0.015308f
C379 VTAIL.n50 VSUBS 0.016208f
C380 VTAIL.n51 VSUBS 0.036182f
C381 VTAIL.n52 VSUBS 0.036182f
C382 VTAIL.n53 VSUBS 0.016208f
C383 VTAIL.n54 VSUBS 0.015308f
C384 VTAIL.n55 VSUBS 0.028487f
C385 VTAIL.n56 VSUBS 0.028487f
C386 VTAIL.n57 VSUBS 0.015308f
C387 VTAIL.n58 VSUBS 0.016208f
C388 VTAIL.n59 VSUBS 0.036182f
C389 VTAIL.n60 VSUBS 0.036182f
C390 VTAIL.n61 VSUBS 0.016208f
C391 VTAIL.n62 VSUBS 0.015308f
C392 VTAIL.n63 VSUBS 0.028487f
C393 VTAIL.n64 VSUBS 0.028487f
C394 VTAIL.n65 VSUBS 0.015308f
C395 VTAIL.n66 VSUBS 0.016208f
C396 VTAIL.n67 VSUBS 0.036182f
C397 VTAIL.n68 VSUBS 0.090478f
C398 VTAIL.n69 VSUBS 0.016208f
C399 VTAIL.n70 VSUBS 0.015308f
C400 VTAIL.n71 VSUBS 0.065847f
C401 VTAIL.n72 VSUBS 0.045629f
C402 VTAIL.n73 VSUBS 1.89957f
C403 VTAIL.n74 VSUBS 0.032148f
C404 VTAIL.n75 VSUBS 0.028487f
C405 VTAIL.n76 VSUBS 0.015308f
C406 VTAIL.n77 VSUBS 0.036182f
C407 VTAIL.n78 VSUBS 0.016208f
C408 VTAIL.n79 VSUBS 0.028487f
C409 VTAIL.n80 VSUBS 0.015308f
C410 VTAIL.n81 VSUBS 0.036182f
C411 VTAIL.n82 VSUBS 0.016208f
C412 VTAIL.n83 VSUBS 0.028487f
C413 VTAIL.n84 VSUBS 0.015308f
C414 VTAIL.n85 VSUBS 0.036182f
C415 VTAIL.n86 VSUBS 0.015758f
C416 VTAIL.n87 VSUBS 0.028487f
C417 VTAIL.n88 VSUBS 0.015758f
C418 VTAIL.n89 VSUBS 0.015308f
C419 VTAIL.n90 VSUBS 0.036182f
C420 VTAIL.n91 VSUBS 0.036182f
C421 VTAIL.n92 VSUBS 0.016208f
C422 VTAIL.n93 VSUBS 0.028487f
C423 VTAIL.n94 VSUBS 0.015308f
C424 VTAIL.n95 VSUBS 0.036182f
C425 VTAIL.n96 VSUBS 0.016208f
C426 VTAIL.n97 VSUBS 1.5944f
C427 VTAIL.n98 VSUBS 0.015308f
C428 VTAIL.t2 VSUBS 0.078116f
C429 VTAIL.n99 VSUBS 0.244447f
C430 VTAIL.n100 VSUBS 0.027218f
C431 VTAIL.n101 VSUBS 0.027137f
C432 VTAIL.n102 VSUBS 0.036182f
C433 VTAIL.n103 VSUBS 0.016208f
C434 VTAIL.n104 VSUBS 0.015308f
C435 VTAIL.n105 VSUBS 0.028487f
C436 VTAIL.n106 VSUBS 0.028487f
C437 VTAIL.n107 VSUBS 0.015308f
C438 VTAIL.n108 VSUBS 0.016208f
C439 VTAIL.n109 VSUBS 0.036182f
C440 VTAIL.n110 VSUBS 0.036182f
C441 VTAIL.n111 VSUBS 0.016208f
C442 VTAIL.n112 VSUBS 0.015308f
C443 VTAIL.n113 VSUBS 0.028487f
C444 VTAIL.n114 VSUBS 0.028487f
C445 VTAIL.n115 VSUBS 0.015308f
C446 VTAIL.n116 VSUBS 0.016208f
C447 VTAIL.n117 VSUBS 0.036182f
C448 VTAIL.n118 VSUBS 0.036182f
C449 VTAIL.n119 VSUBS 0.016208f
C450 VTAIL.n120 VSUBS 0.015308f
C451 VTAIL.n121 VSUBS 0.028487f
C452 VTAIL.n122 VSUBS 0.028487f
C453 VTAIL.n123 VSUBS 0.015308f
C454 VTAIL.n124 VSUBS 0.016208f
C455 VTAIL.n125 VSUBS 0.036182f
C456 VTAIL.n126 VSUBS 0.036182f
C457 VTAIL.n127 VSUBS 0.016208f
C458 VTAIL.n128 VSUBS 0.015308f
C459 VTAIL.n129 VSUBS 0.028487f
C460 VTAIL.n130 VSUBS 0.028487f
C461 VTAIL.n131 VSUBS 0.015308f
C462 VTAIL.n132 VSUBS 0.016208f
C463 VTAIL.n133 VSUBS 0.036182f
C464 VTAIL.n134 VSUBS 0.036182f
C465 VTAIL.n135 VSUBS 0.016208f
C466 VTAIL.n136 VSUBS 0.015308f
C467 VTAIL.n137 VSUBS 0.028487f
C468 VTAIL.n138 VSUBS 0.028487f
C469 VTAIL.n139 VSUBS 0.015308f
C470 VTAIL.n140 VSUBS 0.016208f
C471 VTAIL.n141 VSUBS 0.036182f
C472 VTAIL.n142 VSUBS 0.090478f
C473 VTAIL.n143 VSUBS 0.016208f
C474 VTAIL.n144 VSUBS 0.015308f
C475 VTAIL.n145 VSUBS 0.065847f
C476 VTAIL.n146 VSUBS 0.045629f
C477 VTAIL.n147 VSUBS 1.93498f
C478 VTAIL.n148 VSUBS 0.032148f
C479 VTAIL.n149 VSUBS 0.028487f
C480 VTAIL.n150 VSUBS 0.015308f
C481 VTAIL.n151 VSUBS 0.036182f
C482 VTAIL.n152 VSUBS 0.016208f
C483 VTAIL.n153 VSUBS 0.028487f
C484 VTAIL.n154 VSUBS 0.015308f
C485 VTAIL.n155 VSUBS 0.036182f
C486 VTAIL.n156 VSUBS 0.016208f
C487 VTAIL.n157 VSUBS 0.028487f
C488 VTAIL.n158 VSUBS 0.015308f
C489 VTAIL.n159 VSUBS 0.036182f
C490 VTAIL.n160 VSUBS 0.015758f
C491 VTAIL.n161 VSUBS 0.028487f
C492 VTAIL.n162 VSUBS 0.015758f
C493 VTAIL.n163 VSUBS 0.015308f
C494 VTAIL.n164 VSUBS 0.036182f
C495 VTAIL.n165 VSUBS 0.036182f
C496 VTAIL.n166 VSUBS 0.016208f
C497 VTAIL.n167 VSUBS 0.028487f
C498 VTAIL.n168 VSUBS 0.015308f
C499 VTAIL.n169 VSUBS 0.036182f
C500 VTAIL.n170 VSUBS 0.016208f
C501 VTAIL.n171 VSUBS 1.5944f
C502 VTAIL.n172 VSUBS 0.015308f
C503 VTAIL.t0 VSUBS 0.078116f
C504 VTAIL.n173 VSUBS 0.244447f
C505 VTAIL.n174 VSUBS 0.027218f
C506 VTAIL.n175 VSUBS 0.027137f
C507 VTAIL.n176 VSUBS 0.036182f
C508 VTAIL.n177 VSUBS 0.016208f
C509 VTAIL.n178 VSUBS 0.015308f
C510 VTAIL.n179 VSUBS 0.028487f
C511 VTAIL.n180 VSUBS 0.028487f
C512 VTAIL.n181 VSUBS 0.015308f
C513 VTAIL.n182 VSUBS 0.016208f
C514 VTAIL.n183 VSUBS 0.036182f
C515 VTAIL.n184 VSUBS 0.036182f
C516 VTAIL.n185 VSUBS 0.016208f
C517 VTAIL.n186 VSUBS 0.015308f
C518 VTAIL.n187 VSUBS 0.028487f
C519 VTAIL.n188 VSUBS 0.028487f
C520 VTAIL.n189 VSUBS 0.015308f
C521 VTAIL.n190 VSUBS 0.016208f
C522 VTAIL.n191 VSUBS 0.036182f
C523 VTAIL.n192 VSUBS 0.036182f
C524 VTAIL.n193 VSUBS 0.016208f
C525 VTAIL.n194 VSUBS 0.015308f
C526 VTAIL.n195 VSUBS 0.028487f
C527 VTAIL.n196 VSUBS 0.028487f
C528 VTAIL.n197 VSUBS 0.015308f
C529 VTAIL.n198 VSUBS 0.016208f
C530 VTAIL.n199 VSUBS 0.036182f
C531 VTAIL.n200 VSUBS 0.036182f
C532 VTAIL.n201 VSUBS 0.016208f
C533 VTAIL.n202 VSUBS 0.015308f
C534 VTAIL.n203 VSUBS 0.028487f
C535 VTAIL.n204 VSUBS 0.028487f
C536 VTAIL.n205 VSUBS 0.015308f
C537 VTAIL.n206 VSUBS 0.016208f
C538 VTAIL.n207 VSUBS 0.036182f
C539 VTAIL.n208 VSUBS 0.036182f
C540 VTAIL.n209 VSUBS 0.016208f
C541 VTAIL.n210 VSUBS 0.015308f
C542 VTAIL.n211 VSUBS 0.028487f
C543 VTAIL.n212 VSUBS 0.028487f
C544 VTAIL.n213 VSUBS 0.015308f
C545 VTAIL.n214 VSUBS 0.016208f
C546 VTAIL.n215 VSUBS 0.036182f
C547 VTAIL.n216 VSUBS 0.090478f
C548 VTAIL.n217 VSUBS 0.016208f
C549 VTAIL.n218 VSUBS 0.015308f
C550 VTAIL.n219 VSUBS 0.065847f
C551 VTAIL.n220 VSUBS 0.045629f
C552 VTAIL.n221 VSUBS 1.77197f
C553 VTAIL.n222 VSUBS 0.032148f
C554 VTAIL.n223 VSUBS 0.028487f
C555 VTAIL.n224 VSUBS 0.015308f
C556 VTAIL.n225 VSUBS 0.036182f
C557 VTAIL.n226 VSUBS 0.016208f
C558 VTAIL.n227 VSUBS 0.028487f
C559 VTAIL.n228 VSUBS 0.015308f
C560 VTAIL.n229 VSUBS 0.036182f
C561 VTAIL.n230 VSUBS 0.016208f
C562 VTAIL.n231 VSUBS 0.028487f
C563 VTAIL.n232 VSUBS 0.015308f
C564 VTAIL.n233 VSUBS 0.036182f
C565 VTAIL.n234 VSUBS 0.015758f
C566 VTAIL.n235 VSUBS 0.028487f
C567 VTAIL.n236 VSUBS 0.016208f
C568 VTAIL.n237 VSUBS 0.036182f
C569 VTAIL.n238 VSUBS 0.016208f
C570 VTAIL.n239 VSUBS 0.028487f
C571 VTAIL.n240 VSUBS 0.015308f
C572 VTAIL.n241 VSUBS 0.036182f
C573 VTAIL.n242 VSUBS 0.016208f
C574 VTAIL.n243 VSUBS 1.5944f
C575 VTAIL.n244 VSUBS 0.015308f
C576 VTAIL.t3 VSUBS 0.078116f
C577 VTAIL.n245 VSUBS 0.244447f
C578 VTAIL.n246 VSUBS 0.027218f
C579 VTAIL.n247 VSUBS 0.027137f
C580 VTAIL.n248 VSUBS 0.036182f
C581 VTAIL.n249 VSUBS 0.016208f
C582 VTAIL.n250 VSUBS 0.015308f
C583 VTAIL.n251 VSUBS 0.028487f
C584 VTAIL.n252 VSUBS 0.028487f
C585 VTAIL.n253 VSUBS 0.015308f
C586 VTAIL.n254 VSUBS 0.016208f
C587 VTAIL.n255 VSUBS 0.036182f
C588 VTAIL.n256 VSUBS 0.036182f
C589 VTAIL.n257 VSUBS 0.016208f
C590 VTAIL.n258 VSUBS 0.015308f
C591 VTAIL.n259 VSUBS 0.028487f
C592 VTAIL.n260 VSUBS 0.028487f
C593 VTAIL.n261 VSUBS 0.015308f
C594 VTAIL.n262 VSUBS 0.015308f
C595 VTAIL.n263 VSUBS 0.016208f
C596 VTAIL.n264 VSUBS 0.036182f
C597 VTAIL.n265 VSUBS 0.036182f
C598 VTAIL.n266 VSUBS 0.036182f
C599 VTAIL.n267 VSUBS 0.015758f
C600 VTAIL.n268 VSUBS 0.015308f
C601 VTAIL.n269 VSUBS 0.028487f
C602 VTAIL.n270 VSUBS 0.028487f
C603 VTAIL.n271 VSUBS 0.015308f
C604 VTAIL.n272 VSUBS 0.016208f
C605 VTAIL.n273 VSUBS 0.036182f
C606 VTAIL.n274 VSUBS 0.036182f
C607 VTAIL.n275 VSUBS 0.016208f
C608 VTAIL.n276 VSUBS 0.015308f
C609 VTAIL.n277 VSUBS 0.028487f
C610 VTAIL.n278 VSUBS 0.028487f
C611 VTAIL.n279 VSUBS 0.015308f
C612 VTAIL.n280 VSUBS 0.016208f
C613 VTAIL.n281 VSUBS 0.036182f
C614 VTAIL.n282 VSUBS 0.036182f
C615 VTAIL.n283 VSUBS 0.016208f
C616 VTAIL.n284 VSUBS 0.015308f
C617 VTAIL.n285 VSUBS 0.028487f
C618 VTAIL.n286 VSUBS 0.028487f
C619 VTAIL.n287 VSUBS 0.015308f
C620 VTAIL.n288 VSUBS 0.016208f
C621 VTAIL.n289 VSUBS 0.036182f
C622 VTAIL.n290 VSUBS 0.090478f
C623 VTAIL.n291 VSUBS 0.016208f
C624 VTAIL.n292 VSUBS 0.015308f
C625 VTAIL.n293 VSUBS 0.065847f
C626 VTAIL.n294 VSUBS 0.045629f
C627 VTAIL.n295 VSUBS 1.68275f
C628 VN.t0 VSUBS 3.30987f
C629 VN.t1 VSUBS 3.78291f
C630 B.n0 VSUBS 0.004016f
C631 B.n1 VSUBS 0.004016f
C632 B.n2 VSUBS 0.006351f
C633 B.n3 VSUBS 0.006351f
C634 B.n4 VSUBS 0.006351f
C635 B.n5 VSUBS 0.006351f
C636 B.n6 VSUBS 0.006351f
C637 B.n7 VSUBS 0.006351f
C638 B.n8 VSUBS 0.006351f
C639 B.n9 VSUBS 0.006351f
C640 B.n10 VSUBS 0.006351f
C641 B.n11 VSUBS 0.006351f
C642 B.n12 VSUBS 0.015976f
C643 B.n13 VSUBS 0.006351f
C644 B.n14 VSUBS 0.006351f
C645 B.n15 VSUBS 0.006351f
C646 B.n16 VSUBS 0.006351f
C647 B.n17 VSUBS 0.006351f
C648 B.n18 VSUBS 0.006351f
C649 B.n19 VSUBS 0.006351f
C650 B.n20 VSUBS 0.006351f
C651 B.n21 VSUBS 0.006351f
C652 B.n22 VSUBS 0.006351f
C653 B.n23 VSUBS 0.006351f
C654 B.n24 VSUBS 0.006351f
C655 B.n25 VSUBS 0.006351f
C656 B.n26 VSUBS 0.006351f
C657 B.n27 VSUBS 0.006351f
C658 B.n28 VSUBS 0.006351f
C659 B.n29 VSUBS 0.006351f
C660 B.n30 VSUBS 0.006351f
C661 B.n31 VSUBS 0.006351f
C662 B.n32 VSUBS 0.006351f
C663 B.n33 VSUBS 0.006351f
C664 B.n34 VSUBS 0.006351f
C665 B.n35 VSUBS 0.006351f
C666 B.t11 VSUBS 0.223614f
C667 B.t10 VSUBS 0.244782f
C668 B.t9 VSUBS 0.933328f
C669 B.n36 VSUBS 0.369874f
C670 B.n37 VSUBS 0.244226f
C671 B.n38 VSUBS 0.006351f
C672 B.n39 VSUBS 0.006351f
C673 B.n40 VSUBS 0.006351f
C674 B.n41 VSUBS 0.006351f
C675 B.t8 VSUBS 0.223617f
C676 B.t7 VSUBS 0.244784f
C677 B.t6 VSUBS 0.933328f
C678 B.n42 VSUBS 0.369871f
C679 B.n43 VSUBS 0.244223f
C680 B.n44 VSUBS 0.014714f
C681 B.n45 VSUBS 0.006351f
C682 B.n46 VSUBS 0.006351f
C683 B.n47 VSUBS 0.006351f
C684 B.n48 VSUBS 0.006351f
C685 B.n49 VSUBS 0.006351f
C686 B.n50 VSUBS 0.006351f
C687 B.n51 VSUBS 0.006351f
C688 B.n52 VSUBS 0.006351f
C689 B.n53 VSUBS 0.006351f
C690 B.n54 VSUBS 0.006351f
C691 B.n55 VSUBS 0.006351f
C692 B.n56 VSUBS 0.006351f
C693 B.n57 VSUBS 0.006351f
C694 B.n58 VSUBS 0.006351f
C695 B.n59 VSUBS 0.006351f
C696 B.n60 VSUBS 0.006351f
C697 B.n61 VSUBS 0.006351f
C698 B.n62 VSUBS 0.006351f
C699 B.n63 VSUBS 0.006351f
C700 B.n64 VSUBS 0.006351f
C701 B.n65 VSUBS 0.006351f
C702 B.n66 VSUBS 0.006351f
C703 B.n67 VSUBS 0.015976f
C704 B.n68 VSUBS 0.006351f
C705 B.n69 VSUBS 0.006351f
C706 B.n70 VSUBS 0.006351f
C707 B.n71 VSUBS 0.006351f
C708 B.n72 VSUBS 0.006351f
C709 B.n73 VSUBS 0.006351f
C710 B.n74 VSUBS 0.006351f
C711 B.n75 VSUBS 0.006351f
C712 B.n76 VSUBS 0.006351f
C713 B.n77 VSUBS 0.006351f
C714 B.n78 VSUBS 0.006351f
C715 B.n79 VSUBS 0.006351f
C716 B.n80 VSUBS 0.006351f
C717 B.n81 VSUBS 0.006351f
C718 B.n82 VSUBS 0.006351f
C719 B.n83 VSUBS 0.006351f
C720 B.n84 VSUBS 0.006351f
C721 B.n85 VSUBS 0.006351f
C722 B.n86 VSUBS 0.006351f
C723 B.n87 VSUBS 0.006351f
C724 B.n88 VSUBS 0.015976f
C725 B.n89 VSUBS 0.006351f
C726 B.n90 VSUBS 0.006351f
C727 B.n91 VSUBS 0.006351f
C728 B.n92 VSUBS 0.006351f
C729 B.n93 VSUBS 0.006351f
C730 B.n94 VSUBS 0.006351f
C731 B.n95 VSUBS 0.006351f
C732 B.n96 VSUBS 0.006351f
C733 B.n97 VSUBS 0.006351f
C734 B.n98 VSUBS 0.006351f
C735 B.n99 VSUBS 0.006351f
C736 B.n100 VSUBS 0.006351f
C737 B.n101 VSUBS 0.006351f
C738 B.n102 VSUBS 0.006351f
C739 B.n103 VSUBS 0.006351f
C740 B.n104 VSUBS 0.006351f
C741 B.n105 VSUBS 0.006351f
C742 B.n106 VSUBS 0.006351f
C743 B.n107 VSUBS 0.006351f
C744 B.n108 VSUBS 0.006351f
C745 B.n109 VSUBS 0.006351f
C746 B.n110 VSUBS 0.006351f
C747 B.n111 VSUBS 0.006351f
C748 B.t4 VSUBS 0.223617f
C749 B.t5 VSUBS 0.244784f
C750 B.t3 VSUBS 0.933328f
C751 B.n112 VSUBS 0.369871f
C752 B.n113 VSUBS 0.244223f
C753 B.n114 VSUBS 0.006351f
C754 B.n115 VSUBS 0.006351f
C755 B.n116 VSUBS 0.006351f
C756 B.n117 VSUBS 0.006351f
C757 B.t1 VSUBS 0.223614f
C758 B.t2 VSUBS 0.244782f
C759 B.t0 VSUBS 0.933328f
C760 B.n118 VSUBS 0.369874f
C761 B.n119 VSUBS 0.244226f
C762 B.n120 VSUBS 0.014714f
C763 B.n121 VSUBS 0.006351f
C764 B.n122 VSUBS 0.006351f
C765 B.n123 VSUBS 0.006351f
C766 B.n124 VSUBS 0.006351f
C767 B.n125 VSUBS 0.006351f
C768 B.n126 VSUBS 0.006351f
C769 B.n127 VSUBS 0.006351f
C770 B.n128 VSUBS 0.006351f
C771 B.n129 VSUBS 0.006351f
C772 B.n130 VSUBS 0.006351f
C773 B.n131 VSUBS 0.006351f
C774 B.n132 VSUBS 0.006351f
C775 B.n133 VSUBS 0.006351f
C776 B.n134 VSUBS 0.006351f
C777 B.n135 VSUBS 0.006351f
C778 B.n136 VSUBS 0.006351f
C779 B.n137 VSUBS 0.006351f
C780 B.n138 VSUBS 0.006351f
C781 B.n139 VSUBS 0.006351f
C782 B.n140 VSUBS 0.006351f
C783 B.n141 VSUBS 0.006351f
C784 B.n142 VSUBS 0.006351f
C785 B.n143 VSUBS 0.015976f
C786 B.n144 VSUBS 0.006351f
C787 B.n145 VSUBS 0.006351f
C788 B.n146 VSUBS 0.006351f
C789 B.n147 VSUBS 0.006351f
C790 B.n148 VSUBS 0.006351f
C791 B.n149 VSUBS 0.006351f
C792 B.n150 VSUBS 0.006351f
C793 B.n151 VSUBS 0.006351f
C794 B.n152 VSUBS 0.006351f
C795 B.n153 VSUBS 0.006351f
C796 B.n154 VSUBS 0.006351f
C797 B.n155 VSUBS 0.006351f
C798 B.n156 VSUBS 0.006351f
C799 B.n157 VSUBS 0.006351f
C800 B.n158 VSUBS 0.006351f
C801 B.n159 VSUBS 0.006351f
C802 B.n160 VSUBS 0.006351f
C803 B.n161 VSUBS 0.006351f
C804 B.n162 VSUBS 0.006351f
C805 B.n163 VSUBS 0.006351f
C806 B.n164 VSUBS 0.006351f
C807 B.n165 VSUBS 0.006351f
C808 B.n166 VSUBS 0.006351f
C809 B.n167 VSUBS 0.006351f
C810 B.n168 VSUBS 0.006351f
C811 B.n169 VSUBS 0.006351f
C812 B.n170 VSUBS 0.006351f
C813 B.n171 VSUBS 0.006351f
C814 B.n172 VSUBS 0.006351f
C815 B.n173 VSUBS 0.006351f
C816 B.n174 VSUBS 0.006351f
C817 B.n175 VSUBS 0.006351f
C818 B.n176 VSUBS 0.006351f
C819 B.n177 VSUBS 0.006351f
C820 B.n178 VSUBS 0.006351f
C821 B.n179 VSUBS 0.006351f
C822 B.n180 VSUBS 0.015031f
C823 B.n181 VSUBS 0.015031f
C824 B.n182 VSUBS 0.015976f
C825 B.n183 VSUBS 0.006351f
C826 B.n184 VSUBS 0.006351f
C827 B.n185 VSUBS 0.006351f
C828 B.n186 VSUBS 0.006351f
C829 B.n187 VSUBS 0.006351f
C830 B.n188 VSUBS 0.006351f
C831 B.n189 VSUBS 0.006351f
C832 B.n190 VSUBS 0.006351f
C833 B.n191 VSUBS 0.006351f
C834 B.n192 VSUBS 0.006351f
C835 B.n193 VSUBS 0.006351f
C836 B.n194 VSUBS 0.006351f
C837 B.n195 VSUBS 0.006351f
C838 B.n196 VSUBS 0.006351f
C839 B.n197 VSUBS 0.006351f
C840 B.n198 VSUBS 0.006351f
C841 B.n199 VSUBS 0.006351f
C842 B.n200 VSUBS 0.006351f
C843 B.n201 VSUBS 0.006351f
C844 B.n202 VSUBS 0.006351f
C845 B.n203 VSUBS 0.006351f
C846 B.n204 VSUBS 0.006351f
C847 B.n205 VSUBS 0.006351f
C848 B.n206 VSUBS 0.006351f
C849 B.n207 VSUBS 0.006351f
C850 B.n208 VSUBS 0.006351f
C851 B.n209 VSUBS 0.006351f
C852 B.n210 VSUBS 0.006351f
C853 B.n211 VSUBS 0.006351f
C854 B.n212 VSUBS 0.006351f
C855 B.n213 VSUBS 0.006351f
C856 B.n214 VSUBS 0.006351f
C857 B.n215 VSUBS 0.006351f
C858 B.n216 VSUBS 0.006351f
C859 B.n217 VSUBS 0.006351f
C860 B.n218 VSUBS 0.006351f
C861 B.n219 VSUBS 0.006351f
C862 B.n220 VSUBS 0.006351f
C863 B.n221 VSUBS 0.006351f
C864 B.n222 VSUBS 0.006351f
C865 B.n223 VSUBS 0.006351f
C866 B.n224 VSUBS 0.006351f
C867 B.n225 VSUBS 0.006351f
C868 B.n226 VSUBS 0.006351f
C869 B.n227 VSUBS 0.006351f
C870 B.n228 VSUBS 0.006351f
C871 B.n229 VSUBS 0.006351f
C872 B.n230 VSUBS 0.006351f
C873 B.n231 VSUBS 0.006351f
C874 B.n232 VSUBS 0.006351f
C875 B.n233 VSUBS 0.006351f
C876 B.n234 VSUBS 0.006351f
C877 B.n235 VSUBS 0.006351f
C878 B.n236 VSUBS 0.006351f
C879 B.n237 VSUBS 0.006351f
C880 B.n238 VSUBS 0.006351f
C881 B.n239 VSUBS 0.006351f
C882 B.n240 VSUBS 0.006351f
C883 B.n241 VSUBS 0.006351f
C884 B.n242 VSUBS 0.006351f
C885 B.n243 VSUBS 0.006351f
C886 B.n244 VSUBS 0.006351f
C887 B.n245 VSUBS 0.006351f
C888 B.n246 VSUBS 0.006351f
C889 B.n247 VSUBS 0.006351f
C890 B.n248 VSUBS 0.006351f
C891 B.n249 VSUBS 0.005977f
C892 B.n250 VSUBS 0.006351f
C893 B.n251 VSUBS 0.006351f
C894 B.n252 VSUBS 0.003549f
C895 B.n253 VSUBS 0.006351f
C896 B.n254 VSUBS 0.006351f
C897 B.n255 VSUBS 0.006351f
C898 B.n256 VSUBS 0.006351f
C899 B.n257 VSUBS 0.006351f
C900 B.n258 VSUBS 0.006351f
C901 B.n259 VSUBS 0.006351f
C902 B.n260 VSUBS 0.006351f
C903 B.n261 VSUBS 0.006351f
C904 B.n262 VSUBS 0.006351f
C905 B.n263 VSUBS 0.006351f
C906 B.n264 VSUBS 0.006351f
C907 B.n265 VSUBS 0.003549f
C908 B.n266 VSUBS 0.014714f
C909 B.n267 VSUBS 0.005977f
C910 B.n268 VSUBS 0.006351f
C911 B.n269 VSUBS 0.006351f
C912 B.n270 VSUBS 0.006351f
C913 B.n271 VSUBS 0.006351f
C914 B.n272 VSUBS 0.006351f
C915 B.n273 VSUBS 0.006351f
C916 B.n274 VSUBS 0.006351f
C917 B.n275 VSUBS 0.006351f
C918 B.n276 VSUBS 0.006351f
C919 B.n277 VSUBS 0.006351f
C920 B.n278 VSUBS 0.006351f
C921 B.n279 VSUBS 0.006351f
C922 B.n280 VSUBS 0.006351f
C923 B.n281 VSUBS 0.006351f
C924 B.n282 VSUBS 0.006351f
C925 B.n283 VSUBS 0.006351f
C926 B.n284 VSUBS 0.006351f
C927 B.n285 VSUBS 0.006351f
C928 B.n286 VSUBS 0.006351f
C929 B.n287 VSUBS 0.006351f
C930 B.n288 VSUBS 0.006351f
C931 B.n289 VSUBS 0.006351f
C932 B.n290 VSUBS 0.006351f
C933 B.n291 VSUBS 0.006351f
C934 B.n292 VSUBS 0.006351f
C935 B.n293 VSUBS 0.006351f
C936 B.n294 VSUBS 0.006351f
C937 B.n295 VSUBS 0.006351f
C938 B.n296 VSUBS 0.006351f
C939 B.n297 VSUBS 0.006351f
C940 B.n298 VSUBS 0.006351f
C941 B.n299 VSUBS 0.006351f
C942 B.n300 VSUBS 0.006351f
C943 B.n301 VSUBS 0.006351f
C944 B.n302 VSUBS 0.006351f
C945 B.n303 VSUBS 0.006351f
C946 B.n304 VSUBS 0.006351f
C947 B.n305 VSUBS 0.006351f
C948 B.n306 VSUBS 0.006351f
C949 B.n307 VSUBS 0.006351f
C950 B.n308 VSUBS 0.006351f
C951 B.n309 VSUBS 0.006351f
C952 B.n310 VSUBS 0.006351f
C953 B.n311 VSUBS 0.006351f
C954 B.n312 VSUBS 0.006351f
C955 B.n313 VSUBS 0.006351f
C956 B.n314 VSUBS 0.006351f
C957 B.n315 VSUBS 0.006351f
C958 B.n316 VSUBS 0.006351f
C959 B.n317 VSUBS 0.006351f
C960 B.n318 VSUBS 0.006351f
C961 B.n319 VSUBS 0.006351f
C962 B.n320 VSUBS 0.006351f
C963 B.n321 VSUBS 0.006351f
C964 B.n322 VSUBS 0.006351f
C965 B.n323 VSUBS 0.006351f
C966 B.n324 VSUBS 0.006351f
C967 B.n325 VSUBS 0.006351f
C968 B.n326 VSUBS 0.006351f
C969 B.n327 VSUBS 0.006351f
C970 B.n328 VSUBS 0.006351f
C971 B.n329 VSUBS 0.006351f
C972 B.n330 VSUBS 0.006351f
C973 B.n331 VSUBS 0.006351f
C974 B.n332 VSUBS 0.006351f
C975 B.n333 VSUBS 0.006351f
C976 B.n334 VSUBS 0.006351f
C977 B.n335 VSUBS 0.015976f
C978 B.n336 VSUBS 0.015031f
C979 B.n337 VSUBS 0.015031f
C980 B.n338 VSUBS 0.006351f
C981 B.n339 VSUBS 0.006351f
C982 B.n340 VSUBS 0.006351f
C983 B.n341 VSUBS 0.006351f
C984 B.n342 VSUBS 0.006351f
C985 B.n343 VSUBS 0.006351f
C986 B.n344 VSUBS 0.006351f
C987 B.n345 VSUBS 0.006351f
C988 B.n346 VSUBS 0.006351f
C989 B.n347 VSUBS 0.006351f
C990 B.n348 VSUBS 0.006351f
C991 B.n349 VSUBS 0.006351f
C992 B.n350 VSUBS 0.006351f
C993 B.n351 VSUBS 0.006351f
C994 B.n352 VSUBS 0.006351f
C995 B.n353 VSUBS 0.006351f
C996 B.n354 VSUBS 0.006351f
C997 B.n355 VSUBS 0.006351f
C998 B.n356 VSUBS 0.006351f
C999 B.n357 VSUBS 0.006351f
C1000 B.n358 VSUBS 0.006351f
C1001 B.n359 VSUBS 0.006351f
C1002 B.n360 VSUBS 0.006351f
C1003 B.n361 VSUBS 0.006351f
C1004 B.n362 VSUBS 0.006351f
C1005 B.n363 VSUBS 0.006351f
C1006 B.n364 VSUBS 0.006351f
C1007 B.n365 VSUBS 0.006351f
C1008 B.n366 VSUBS 0.006351f
C1009 B.n367 VSUBS 0.006351f
C1010 B.n368 VSUBS 0.006351f
C1011 B.n369 VSUBS 0.006351f
C1012 B.n370 VSUBS 0.006351f
C1013 B.n371 VSUBS 0.006351f
C1014 B.n372 VSUBS 0.006351f
C1015 B.n373 VSUBS 0.006351f
C1016 B.n374 VSUBS 0.006351f
C1017 B.n375 VSUBS 0.006351f
C1018 B.n376 VSUBS 0.006351f
C1019 B.n377 VSUBS 0.006351f
C1020 B.n378 VSUBS 0.006351f
C1021 B.n379 VSUBS 0.006351f
C1022 B.n380 VSUBS 0.006351f
C1023 B.n381 VSUBS 0.006351f
C1024 B.n382 VSUBS 0.006351f
C1025 B.n383 VSUBS 0.006351f
C1026 B.n384 VSUBS 0.006351f
C1027 B.n385 VSUBS 0.006351f
C1028 B.n386 VSUBS 0.006351f
C1029 B.n387 VSUBS 0.006351f
C1030 B.n388 VSUBS 0.006351f
C1031 B.n389 VSUBS 0.006351f
C1032 B.n390 VSUBS 0.006351f
C1033 B.n391 VSUBS 0.006351f
C1034 B.n392 VSUBS 0.006351f
C1035 B.n393 VSUBS 0.006351f
C1036 B.n394 VSUBS 0.006351f
C1037 B.n395 VSUBS 0.006351f
C1038 B.n396 VSUBS 0.015031f
C1039 B.n397 VSUBS 0.015735f
C1040 B.n398 VSUBS 0.015272f
C1041 B.n399 VSUBS 0.006351f
C1042 B.n400 VSUBS 0.006351f
C1043 B.n401 VSUBS 0.006351f
C1044 B.n402 VSUBS 0.006351f
C1045 B.n403 VSUBS 0.006351f
C1046 B.n404 VSUBS 0.006351f
C1047 B.n405 VSUBS 0.006351f
C1048 B.n406 VSUBS 0.006351f
C1049 B.n407 VSUBS 0.006351f
C1050 B.n408 VSUBS 0.006351f
C1051 B.n409 VSUBS 0.006351f
C1052 B.n410 VSUBS 0.006351f
C1053 B.n411 VSUBS 0.006351f
C1054 B.n412 VSUBS 0.006351f
C1055 B.n413 VSUBS 0.006351f
C1056 B.n414 VSUBS 0.006351f
C1057 B.n415 VSUBS 0.006351f
C1058 B.n416 VSUBS 0.006351f
C1059 B.n417 VSUBS 0.006351f
C1060 B.n418 VSUBS 0.006351f
C1061 B.n419 VSUBS 0.006351f
C1062 B.n420 VSUBS 0.006351f
C1063 B.n421 VSUBS 0.006351f
C1064 B.n422 VSUBS 0.006351f
C1065 B.n423 VSUBS 0.006351f
C1066 B.n424 VSUBS 0.006351f
C1067 B.n425 VSUBS 0.006351f
C1068 B.n426 VSUBS 0.006351f
C1069 B.n427 VSUBS 0.006351f
C1070 B.n428 VSUBS 0.006351f
C1071 B.n429 VSUBS 0.006351f
C1072 B.n430 VSUBS 0.006351f
C1073 B.n431 VSUBS 0.006351f
C1074 B.n432 VSUBS 0.006351f
C1075 B.n433 VSUBS 0.006351f
C1076 B.n434 VSUBS 0.006351f
C1077 B.n435 VSUBS 0.006351f
C1078 B.n436 VSUBS 0.006351f
C1079 B.n437 VSUBS 0.006351f
C1080 B.n438 VSUBS 0.006351f
C1081 B.n439 VSUBS 0.006351f
C1082 B.n440 VSUBS 0.006351f
C1083 B.n441 VSUBS 0.006351f
C1084 B.n442 VSUBS 0.006351f
C1085 B.n443 VSUBS 0.006351f
C1086 B.n444 VSUBS 0.006351f
C1087 B.n445 VSUBS 0.006351f
C1088 B.n446 VSUBS 0.006351f
C1089 B.n447 VSUBS 0.006351f
C1090 B.n448 VSUBS 0.006351f
C1091 B.n449 VSUBS 0.006351f
C1092 B.n450 VSUBS 0.006351f
C1093 B.n451 VSUBS 0.006351f
C1094 B.n452 VSUBS 0.006351f
C1095 B.n453 VSUBS 0.006351f
C1096 B.n454 VSUBS 0.006351f
C1097 B.n455 VSUBS 0.006351f
C1098 B.n456 VSUBS 0.006351f
C1099 B.n457 VSUBS 0.006351f
C1100 B.n458 VSUBS 0.006351f
C1101 B.n459 VSUBS 0.006351f
C1102 B.n460 VSUBS 0.006351f
C1103 B.n461 VSUBS 0.006351f
C1104 B.n462 VSUBS 0.006351f
C1105 B.n463 VSUBS 0.006351f
C1106 B.n464 VSUBS 0.006351f
C1107 B.n465 VSUBS 0.005977f
C1108 B.n466 VSUBS 0.006351f
C1109 B.n467 VSUBS 0.006351f
C1110 B.n468 VSUBS 0.003549f
C1111 B.n469 VSUBS 0.006351f
C1112 B.n470 VSUBS 0.006351f
C1113 B.n471 VSUBS 0.006351f
C1114 B.n472 VSUBS 0.006351f
C1115 B.n473 VSUBS 0.006351f
C1116 B.n474 VSUBS 0.006351f
C1117 B.n475 VSUBS 0.006351f
C1118 B.n476 VSUBS 0.006351f
C1119 B.n477 VSUBS 0.006351f
C1120 B.n478 VSUBS 0.006351f
C1121 B.n479 VSUBS 0.006351f
C1122 B.n480 VSUBS 0.006351f
C1123 B.n481 VSUBS 0.003549f
C1124 B.n482 VSUBS 0.014714f
C1125 B.n483 VSUBS 0.005977f
C1126 B.n484 VSUBS 0.006351f
C1127 B.n485 VSUBS 0.006351f
C1128 B.n486 VSUBS 0.006351f
C1129 B.n487 VSUBS 0.006351f
C1130 B.n488 VSUBS 0.006351f
C1131 B.n489 VSUBS 0.006351f
C1132 B.n490 VSUBS 0.006351f
C1133 B.n491 VSUBS 0.006351f
C1134 B.n492 VSUBS 0.006351f
C1135 B.n493 VSUBS 0.006351f
C1136 B.n494 VSUBS 0.006351f
C1137 B.n495 VSUBS 0.006351f
C1138 B.n496 VSUBS 0.006351f
C1139 B.n497 VSUBS 0.006351f
C1140 B.n498 VSUBS 0.006351f
C1141 B.n499 VSUBS 0.006351f
C1142 B.n500 VSUBS 0.006351f
C1143 B.n501 VSUBS 0.006351f
C1144 B.n502 VSUBS 0.006351f
C1145 B.n503 VSUBS 0.006351f
C1146 B.n504 VSUBS 0.006351f
C1147 B.n505 VSUBS 0.006351f
C1148 B.n506 VSUBS 0.006351f
C1149 B.n507 VSUBS 0.006351f
C1150 B.n508 VSUBS 0.006351f
C1151 B.n509 VSUBS 0.006351f
C1152 B.n510 VSUBS 0.006351f
C1153 B.n511 VSUBS 0.006351f
C1154 B.n512 VSUBS 0.006351f
C1155 B.n513 VSUBS 0.006351f
C1156 B.n514 VSUBS 0.006351f
C1157 B.n515 VSUBS 0.006351f
C1158 B.n516 VSUBS 0.006351f
C1159 B.n517 VSUBS 0.006351f
C1160 B.n518 VSUBS 0.006351f
C1161 B.n519 VSUBS 0.006351f
C1162 B.n520 VSUBS 0.006351f
C1163 B.n521 VSUBS 0.006351f
C1164 B.n522 VSUBS 0.006351f
C1165 B.n523 VSUBS 0.006351f
C1166 B.n524 VSUBS 0.006351f
C1167 B.n525 VSUBS 0.006351f
C1168 B.n526 VSUBS 0.006351f
C1169 B.n527 VSUBS 0.006351f
C1170 B.n528 VSUBS 0.006351f
C1171 B.n529 VSUBS 0.006351f
C1172 B.n530 VSUBS 0.006351f
C1173 B.n531 VSUBS 0.006351f
C1174 B.n532 VSUBS 0.006351f
C1175 B.n533 VSUBS 0.006351f
C1176 B.n534 VSUBS 0.006351f
C1177 B.n535 VSUBS 0.006351f
C1178 B.n536 VSUBS 0.006351f
C1179 B.n537 VSUBS 0.006351f
C1180 B.n538 VSUBS 0.006351f
C1181 B.n539 VSUBS 0.006351f
C1182 B.n540 VSUBS 0.006351f
C1183 B.n541 VSUBS 0.006351f
C1184 B.n542 VSUBS 0.006351f
C1185 B.n543 VSUBS 0.006351f
C1186 B.n544 VSUBS 0.006351f
C1187 B.n545 VSUBS 0.006351f
C1188 B.n546 VSUBS 0.006351f
C1189 B.n547 VSUBS 0.006351f
C1190 B.n548 VSUBS 0.006351f
C1191 B.n549 VSUBS 0.006351f
C1192 B.n550 VSUBS 0.006351f
C1193 B.n551 VSUBS 0.015976f
C1194 B.n552 VSUBS 0.015031f
C1195 B.n553 VSUBS 0.015031f
C1196 B.n554 VSUBS 0.006351f
C1197 B.n555 VSUBS 0.006351f
C1198 B.n556 VSUBS 0.006351f
C1199 B.n557 VSUBS 0.006351f
C1200 B.n558 VSUBS 0.006351f
C1201 B.n559 VSUBS 0.006351f
C1202 B.n560 VSUBS 0.006351f
C1203 B.n561 VSUBS 0.006351f
C1204 B.n562 VSUBS 0.006351f
C1205 B.n563 VSUBS 0.006351f
C1206 B.n564 VSUBS 0.006351f
C1207 B.n565 VSUBS 0.006351f
C1208 B.n566 VSUBS 0.006351f
C1209 B.n567 VSUBS 0.006351f
C1210 B.n568 VSUBS 0.006351f
C1211 B.n569 VSUBS 0.006351f
C1212 B.n570 VSUBS 0.006351f
C1213 B.n571 VSUBS 0.006351f
C1214 B.n572 VSUBS 0.006351f
C1215 B.n573 VSUBS 0.006351f
C1216 B.n574 VSUBS 0.006351f
C1217 B.n575 VSUBS 0.006351f
C1218 B.n576 VSUBS 0.006351f
C1219 B.n577 VSUBS 0.006351f
C1220 B.n578 VSUBS 0.006351f
C1221 B.n579 VSUBS 0.006351f
C1222 B.n580 VSUBS 0.006351f
C1223 B.n581 VSUBS 0.006351f
C1224 B.n582 VSUBS 0.006351f
C1225 B.n583 VSUBS 0.014381f
.ends

