* NGSPICE file created from diff_pair_sample_0662.ext - technology: sky130A

.subckt diff_pair_sample_0662 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t1 VN.t0 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=2.5233 pd=13.72 as=2.5233 ps=13.72 w=6.47 l=0.76
X1 B.t15 B.t13 B.t14 B.t7 sky130_fd_pr__nfet_01v8 ad=2.5233 pd=13.72 as=0 ps=0 w=6.47 l=0.76
X2 B.t12 B.t10 B.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=2.5233 pd=13.72 as=0 ps=0 w=6.47 l=0.76
X3 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=2.5233 pd=13.72 as=0 ps=0 w=6.47 l=0.76
X4 VDD1.t1 VP.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.5233 pd=13.72 as=2.5233 ps=13.72 w=6.47 l=0.76
X5 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=2.5233 pd=13.72 as=0 ps=0 w=6.47 l=0.76
X6 VDD1.t0 VP.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.5233 pd=13.72 as=2.5233 ps=13.72 w=6.47 l=0.76
X7 VDD2.t0 VN.t1 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=2.5233 pd=13.72 as=2.5233 ps=13.72 w=6.47 l=0.76
R0 VN VN.t0 454.455
R1 VN VN.t1 418.524
R2 VTAIL.n134 VTAIL.n133 289.615
R3 VTAIL.n32 VTAIL.n31 289.615
R4 VTAIL.n100 VTAIL.n99 289.615
R5 VTAIL.n66 VTAIL.n65 289.615
R6 VTAIL.n112 VTAIL.n111 185
R7 VTAIL.n117 VTAIL.n116 185
R8 VTAIL.n119 VTAIL.n118 185
R9 VTAIL.n108 VTAIL.n107 185
R10 VTAIL.n125 VTAIL.n124 185
R11 VTAIL.n127 VTAIL.n126 185
R12 VTAIL.n104 VTAIL.n103 185
R13 VTAIL.n133 VTAIL.n132 185
R14 VTAIL.n10 VTAIL.n9 185
R15 VTAIL.n15 VTAIL.n14 185
R16 VTAIL.n17 VTAIL.n16 185
R17 VTAIL.n6 VTAIL.n5 185
R18 VTAIL.n23 VTAIL.n22 185
R19 VTAIL.n25 VTAIL.n24 185
R20 VTAIL.n2 VTAIL.n1 185
R21 VTAIL.n31 VTAIL.n30 185
R22 VTAIL.n99 VTAIL.n98 185
R23 VTAIL.n70 VTAIL.n69 185
R24 VTAIL.n93 VTAIL.n92 185
R25 VTAIL.n91 VTAIL.n90 185
R26 VTAIL.n74 VTAIL.n73 185
R27 VTAIL.n85 VTAIL.n84 185
R28 VTAIL.n83 VTAIL.n82 185
R29 VTAIL.n78 VTAIL.n77 185
R30 VTAIL.n65 VTAIL.n64 185
R31 VTAIL.n36 VTAIL.n35 185
R32 VTAIL.n59 VTAIL.n58 185
R33 VTAIL.n57 VTAIL.n56 185
R34 VTAIL.n40 VTAIL.n39 185
R35 VTAIL.n51 VTAIL.n50 185
R36 VTAIL.n49 VTAIL.n48 185
R37 VTAIL.n44 VTAIL.n43 185
R38 VTAIL.n45 VTAIL.t2 149.525
R39 VTAIL.n113 VTAIL.t3 149.525
R40 VTAIL.n11 VTAIL.t0 149.525
R41 VTAIL.n79 VTAIL.t1 149.525
R42 VTAIL.n117 VTAIL.n111 104.615
R43 VTAIL.n118 VTAIL.n117 104.615
R44 VTAIL.n118 VTAIL.n107 104.615
R45 VTAIL.n125 VTAIL.n107 104.615
R46 VTAIL.n126 VTAIL.n125 104.615
R47 VTAIL.n126 VTAIL.n103 104.615
R48 VTAIL.n133 VTAIL.n103 104.615
R49 VTAIL.n15 VTAIL.n9 104.615
R50 VTAIL.n16 VTAIL.n15 104.615
R51 VTAIL.n16 VTAIL.n5 104.615
R52 VTAIL.n23 VTAIL.n5 104.615
R53 VTAIL.n24 VTAIL.n23 104.615
R54 VTAIL.n24 VTAIL.n1 104.615
R55 VTAIL.n31 VTAIL.n1 104.615
R56 VTAIL.n99 VTAIL.n69 104.615
R57 VTAIL.n92 VTAIL.n69 104.615
R58 VTAIL.n92 VTAIL.n91 104.615
R59 VTAIL.n91 VTAIL.n73 104.615
R60 VTAIL.n84 VTAIL.n73 104.615
R61 VTAIL.n84 VTAIL.n83 104.615
R62 VTAIL.n83 VTAIL.n77 104.615
R63 VTAIL.n65 VTAIL.n35 104.615
R64 VTAIL.n58 VTAIL.n35 104.615
R65 VTAIL.n58 VTAIL.n57 104.615
R66 VTAIL.n57 VTAIL.n39 104.615
R67 VTAIL.n50 VTAIL.n39 104.615
R68 VTAIL.n50 VTAIL.n49 104.615
R69 VTAIL.n49 VTAIL.n43 104.615
R70 VTAIL.t3 VTAIL.n111 52.3082
R71 VTAIL.t0 VTAIL.n9 52.3082
R72 VTAIL.t1 VTAIL.n77 52.3082
R73 VTAIL.t2 VTAIL.n43 52.3082
R74 VTAIL.n135 VTAIL.n134 33.9308
R75 VTAIL.n33 VTAIL.n32 33.9308
R76 VTAIL.n101 VTAIL.n100 33.9308
R77 VTAIL.n67 VTAIL.n66 33.9308
R78 VTAIL.n67 VTAIL.n33 19.841
R79 VTAIL.n135 VTAIL.n101 18.9014
R80 VTAIL.n132 VTAIL.n102 12.8005
R81 VTAIL.n30 VTAIL.n0 12.8005
R82 VTAIL.n98 VTAIL.n68 12.8005
R83 VTAIL.n64 VTAIL.n34 12.8005
R84 VTAIL.n131 VTAIL.n104 12.0247
R85 VTAIL.n29 VTAIL.n2 12.0247
R86 VTAIL.n97 VTAIL.n70 12.0247
R87 VTAIL.n63 VTAIL.n36 12.0247
R88 VTAIL.n128 VTAIL.n127 11.249
R89 VTAIL.n26 VTAIL.n25 11.249
R90 VTAIL.n94 VTAIL.n93 11.249
R91 VTAIL.n60 VTAIL.n59 11.249
R92 VTAIL.n124 VTAIL.n106 10.4732
R93 VTAIL.n22 VTAIL.n4 10.4732
R94 VTAIL.n90 VTAIL.n72 10.4732
R95 VTAIL.n56 VTAIL.n38 10.4732
R96 VTAIL.n113 VTAIL.n112 10.2746
R97 VTAIL.n11 VTAIL.n10 10.2746
R98 VTAIL.n79 VTAIL.n78 10.2746
R99 VTAIL.n45 VTAIL.n44 10.2746
R100 VTAIL.n123 VTAIL.n108 9.69747
R101 VTAIL.n21 VTAIL.n6 9.69747
R102 VTAIL.n89 VTAIL.n74 9.69747
R103 VTAIL.n55 VTAIL.n40 9.69747
R104 VTAIL.n130 VTAIL.n102 9.45567
R105 VTAIL.n28 VTAIL.n0 9.45567
R106 VTAIL.n96 VTAIL.n68 9.45567
R107 VTAIL.n62 VTAIL.n34 9.45567
R108 VTAIL.n115 VTAIL.n114 9.3005
R109 VTAIL.n110 VTAIL.n109 9.3005
R110 VTAIL.n121 VTAIL.n120 9.3005
R111 VTAIL.n123 VTAIL.n122 9.3005
R112 VTAIL.n106 VTAIL.n105 9.3005
R113 VTAIL.n129 VTAIL.n128 9.3005
R114 VTAIL.n131 VTAIL.n130 9.3005
R115 VTAIL.n13 VTAIL.n12 9.3005
R116 VTAIL.n8 VTAIL.n7 9.3005
R117 VTAIL.n19 VTAIL.n18 9.3005
R118 VTAIL.n21 VTAIL.n20 9.3005
R119 VTAIL.n4 VTAIL.n3 9.3005
R120 VTAIL.n27 VTAIL.n26 9.3005
R121 VTAIL.n29 VTAIL.n28 9.3005
R122 VTAIL.n97 VTAIL.n96 9.3005
R123 VTAIL.n95 VTAIL.n94 9.3005
R124 VTAIL.n72 VTAIL.n71 9.3005
R125 VTAIL.n89 VTAIL.n88 9.3005
R126 VTAIL.n87 VTAIL.n86 9.3005
R127 VTAIL.n76 VTAIL.n75 9.3005
R128 VTAIL.n81 VTAIL.n80 9.3005
R129 VTAIL.n42 VTAIL.n41 9.3005
R130 VTAIL.n53 VTAIL.n52 9.3005
R131 VTAIL.n55 VTAIL.n54 9.3005
R132 VTAIL.n38 VTAIL.n37 9.3005
R133 VTAIL.n61 VTAIL.n60 9.3005
R134 VTAIL.n63 VTAIL.n62 9.3005
R135 VTAIL.n47 VTAIL.n46 9.3005
R136 VTAIL.n120 VTAIL.n119 8.92171
R137 VTAIL.n18 VTAIL.n17 8.92171
R138 VTAIL.n86 VTAIL.n85 8.92171
R139 VTAIL.n52 VTAIL.n51 8.92171
R140 VTAIL.n116 VTAIL.n110 8.14595
R141 VTAIL.n14 VTAIL.n8 8.14595
R142 VTAIL.n82 VTAIL.n76 8.14595
R143 VTAIL.n48 VTAIL.n42 8.14595
R144 VTAIL.n115 VTAIL.n112 7.3702
R145 VTAIL.n13 VTAIL.n10 7.3702
R146 VTAIL.n81 VTAIL.n78 7.3702
R147 VTAIL.n47 VTAIL.n44 7.3702
R148 VTAIL.n116 VTAIL.n115 5.81868
R149 VTAIL.n14 VTAIL.n13 5.81868
R150 VTAIL.n82 VTAIL.n81 5.81868
R151 VTAIL.n48 VTAIL.n47 5.81868
R152 VTAIL.n119 VTAIL.n110 5.04292
R153 VTAIL.n17 VTAIL.n8 5.04292
R154 VTAIL.n85 VTAIL.n76 5.04292
R155 VTAIL.n51 VTAIL.n42 5.04292
R156 VTAIL.n120 VTAIL.n108 4.26717
R157 VTAIL.n18 VTAIL.n6 4.26717
R158 VTAIL.n86 VTAIL.n74 4.26717
R159 VTAIL.n52 VTAIL.n40 4.26717
R160 VTAIL.n124 VTAIL.n123 3.49141
R161 VTAIL.n22 VTAIL.n21 3.49141
R162 VTAIL.n90 VTAIL.n89 3.49141
R163 VTAIL.n56 VTAIL.n55 3.49141
R164 VTAIL.n46 VTAIL.n45 2.84308
R165 VTAIL.n114 VTAIL.n113 2.84308
R166 VTAIL.n12 VTAIL.n11 2.84308
R167 VTAIL.n80 VTAIL.n79 2.84308
R168 VTAIL.n127 VTAIL.n106 2.71565
R169 VTAIL.n25 VTAIL.n4 2.71565
R170 VTAIL.n93 VTAIL.n72 2.71565
R171 VTAIL.n59 VTAIL.n38 2.71565
R172 VTAIL.n128 VTAIL.n104 1.93989
R173 VTAIL.n26 VTAIL.n2 1.93989
R174 VTAIL.n94 VTAIL.n70 1.93989
R175 VTAIL.n60 VTAIL.n36 1.93989
R176 VTAIL.n132 VTAIL.n131 1.16414
R177 VTAIL.n30 VTAIL.n29 1.16414
R178 VTAIL.n98 VTAIL.n97 1.16414
R179 VTAIL.n64 VTAIL.n63 1.16414
R180 VTAIL.n101 VTAIL.n67 0.940155
R181 VTAIL VTAIL.n33 0.763431
R182 VTAIL.n134 VTAIL.n102 0.388379
R183 VTAIL.n32 VTAIL.n0 0.388379
R184 VTAIL.n100 VTAIL.n68 0.388379
R185 VTAIL.n66 VTAIL.n34 0.388379
R186 VTAIL VTAIL.n135 0.177224
R187 VTAIL.n114 VTAIL.n109 0.155672
R188 VTAIL.n121 VTAIL.n109 0.155672
R189 VTAIL.n122 VTAIL.n121 0.155672
R190 VTAIL.n122 VTAIL.n105 0.155672
R191 VTAIL.n129 VTAIL.n105 0.155672
R192 VTAIL.n130 VTAIL.n129 0.155672
R193 VTAIL.n12 VTAIL.n7 0.155672
R194 VTAIL.n19 VTAIL.n7 0.155672
R195 VTAIL.n20 VTAIL.n19 0.155672
R196 VTAIL.n20 VTAIL.n3 0.155672
R197 VTAIL.n27 VTAIL.n3 0.155672
R198 VTAIL.n28 VTAIL.n27 0.155672
R199 VTAIL.n96 VTAIL.n95 0.155672
R200 VTAIL.n95 VTAIL.n71 0.155672
R201 VTAIL.n88 VTAIL.n71 0.155672
R202 VTAIL.n88 VTAIL.n87 0.155672
R203 VTAIL.n87 VTAIL.n75 0.155672
R204 VTAIL.n80 VTAIL.n75 0.155672
R205 VTAIL.n62 VTAIL.n61 0.155672
R206 VTAIL.n61 VTAIL.n37 0.155672
R207 VTAIL.n54 VTAIL.n37 0.155672
R208 VTAIL.n54 VTAIL.n53 0.155672
R209 VTAIL.n53 VTAIL.n41 0.155672
R210 VTAIL.n46 VTAIL.n41 0.155672
R211 VDD2.n65 VDD2.n64 289.615
R212 VDD2.n32 VDD2.n31 289.615
R213 VDD2.n64 VDD2.n63 185
R214 VDD2.n35 VDD2.n34 185
R215 VDD2.n58 VDD2.n57 185
R216 VDD2.n56 VDD2.n55 185
R217 VDD2.n39 VDD2.n38 185
R218 VDD2.n50 VDD2.n49 185
R219 VDD2.n48 VDD2.n47 185
R220 VDD2.n43 VDD2.n42 185
R221 VDD2.n10 VDD2.n9 185
R222 VDD2.n15 VDD2.n14 185
R223 VDD2.n17 VDD2.n16 185
R224 VDD2.n6 VDD2.n5 185
R225 VDD2.n23 VDD2.n22 185
R226 VDD2.n25 VDD2.n24 185
R227 VDD2.n2 VDD2.n1 185
R228 VDD2.n31 VDD2.n30 185
R229 VDD2.n44 VDD2.t1 149.525
R230 VDD2.n11 VDD2.t0 149.525
R231 VDD2.n64 VDD2.n34 104.615
R232 VDD2.n57 VDD2.n34 104.615
R233 VDD2.n57 VDD2.n56 104.615
R234 VDD2.n56 VDD2.n38 104.615
R235 VDD2.n49 VDD2.n38 104.615
R236 VDD2.n49 VDD2.n48 104.615
R237 VDD2.n48 VDD2.n42 104.615
R238 VDD2.n15 VDD2.n9 104.615
R239 VDD2.n16 VDD2.n15 104.615
R240 VDD2.n16 VDD2.n5 104.615
R241 VDD2.n23 VDD2.n5 104.615
R242 VDD2.n24 VDD2.n23 104.615
R243 VDD2.n24 VDD2.n1 104.615
R244 VDD2.n31 VDD2.n1 104.615
R245 VDD2.n66 VDD2.n32 81.7432
R246 VDD2.t1 VDD2.n42 52.3082
R247 VDD2.t0 VDD2.n9 52.3082
R248 VDD2.n66 VDD2.n65 50.6096
R249 VDD2.n63 VDD2.n33 12.8005
R250 VDD2.n30 VDD2.n0 12.8005
R251 VDD2.n62 VDD2.n35 12.0247
R252 VDD2.n29 VDD2.n2 12.0247
R253 VDD2.n59 VDD2.n58 11.249
R254 VDD2.n26 VDD2.n25 11.249
R255 VDD2.n55 VDD2.n37 10.4732
R256 VDD2.n22 VDD2.n4 10.4732
R257 VDD2.n44 VDD2.n43 10.2746
R258 VDD2.n11 VDD2.n10 10.2746
R259 VDD2.n54 VDD2.n39 9.69747
R260 VDD2.n21 VDD2.n6 9.69747
R261 VDD2.n61 VDD2.n33 9.45567
R262 VDD2.n28 VDD2.n0 9.45567
R263 VDD2.n62 VDD2.n61 9.3005
R264 VDD2.n60 VDD2.n59 9.3005
R265 VDD2.n37 VDD2.n36 9.3005
R266 VDD2.n54 VDD2.n53 9.3005
R267 VDD2.n52 VDD2.n51 9.3005
R268 VDD2.n41 VDD2.n40 9.3005
R269 VDD2.n46 VDD2.n45 9.3005
R270 VDD2.n13 VDD2.n12 9.3005
R271 VDD2.n8 VDD2.n7 9.3005
R272 VDD2.n19 VDD2.n18 9.3005
R273 VDD2.n21 VDD2.n20 9.3005
R274 VDD2.n4 VDD2.n3 9.3005
R275 VDD2.n27 VDD2.n26 9.3005
R276 VDD2.n29 VDD2.n28 9.3005
R277 VDD2.n51 VDD2.n50 8.92171
R278 VDD2.n18 VDD2.n17 8.92171
R279 VDD2.n47 VDD2.n41 8.14595
R280 VDD2.n14 VDD2.n8 8.14595
R281 VDD2.n46 VDD2.n43 7.3702
R282 VDD2.n13 VDD2.n10 7.3702
R283 VDD2.n47 VDD2.n46 5.81868
R284 VDD2.n14 VDD2.n13 5.81868
R285 VDD2.n50 VDD2.n41 5.04292
R286 VDD2.n17 VDD2.n8 5.04292
R287 VDD2.n51 VDD2.n39 4.26717
R288 VDD2.n18 VDD2.n6 4.26717
R289 VDD2.n55 VDD2.n54 3.49141
R290 VDD2.n22 VDD2.n21 3.49141
R291 VDD2.n45 VDD2.n44 2.84308
R292 VDD2.n12 VDD2.n11 2.84308
R293 VDD2.n58 VDD2.n37 2.71565
R294 VDD2.n25 VDD2.n4 2.71565
R295 VDD2.n59 VDD2.n35 1.93989
R296 VDD2.n26 VDD2.n2 1.93989
R297 VDD2.n63 VDD2.n62 1.16414
R298 VDD2.n30 VDD2.n29 1.16414
R299 VDD2.n65 VDD2.n33 0.388379
R300 VDD2.n32 VDD2.n0 0.388379
R301 VDD2 VDD2.n66 0.293603
R302 VDD2.n61 VDD2.n60 0.155672
R303 VDD2.n60 VDD2.n36 0.155672
R304 VDD2.n53 VDD2.n36 0.155672
R305 VDD2.n53 VDD2.n52 0.155672
R306 VDD2.n52 VDD2.n40 0.155672
R307 VDD2.n45 VDD2.n40 0.155672
R308 VDD2.n12 VDD2.n7 0.155672
R309 VDD2.n19 VDD2.n7 0.155672
R310 VDD2.n20 VDD2.n19 0.155672
R311 VDD2.n20 VDD2.n3 0.155672
R312 VDD2.n27 VDD2.n3 0.155672
R313 VDD2.n28 VDD2.n27 0.155672
R314 B.n310 B.n309 585
R315 B.n312 B.n65 585
R316 B.n315 B.n314 585
R317 B.n316 B.n64 585
R318 B.n318 B.n317 585
R319 B.n320 B.n63 585
R320 B.n323 B.n322 585
R321 B.n324 B.n62 585
R322 B.n326 B.n325 585
R323 B.n328 B.n61 585
R324 B.n331 B.n330 585
R325 B.n332 B.n60 585
R326 B.n334 B.n333 585
R327 B.n336 B.n59 585
R328 B.n339 B.n338 585
R329 B.n340 B.n58 585
R330 B.n342 B.n341 585
R331 B.n344 B.n57 585
R332 B.n347 B.n346 585
R333 B.n348 B.n56 585
R334 B.n350 B.n349 585
R335 B.n352 B.n55 585
R336 B.n355 B.n354 585
R337 B.n356 B.n51 585
R338 B.n358 B.n357 585
R339 B.n360 B.n50 585
R340 B.n363 B.n362 585
R341 B.n364 B.n49 585
R342 B.n366 B.n365 585
R343 B.n368 B.n48 585
R344 B.n371 B.n370 585
R345 B.n372 B.n47 585
R346 B.n374 B.n373 585
R347 B.n376 B.n46 585
R348 B.n379 B.n378 585
R349 B.n381 B.n43 585
R350 B.n383 B.n382 585
R351 B.n385 B.n42 585
R352 B.n388 B.n387 585
R353 B.n389 B.n41 585
R354 B.n391 B.n390 585
R355 B.n393 B.n40 585
R356 B.n396 B.n395 585
R357 B.n397 B.n39 585
R358 B.n399 B.n398 585
R359 B.n401 B.n38 585
R360 B.n404 B.n403 585
R361 B.n405 B.n37 585
R362 B.n407 B.n406 585
R363 B.n409 B.n36 585
R364 B.n412 B.n411 585
R365 B.n413 B.n35 585
R366 B.n415 B.n414 585
R367 B.n417 B.n34 585
R368 B.n420 B.n419 585
R369 B.n421 B.n33 585
R370 B.n423 B.n422 585
R371 B.n425 B.n32 585
R372 B.n428 B.n427 585
R373 B.n429 B.n31 585
R374 B.n308 B.n29 585
R375 B.n432 B.n29 585
R376 B.n307 B.n28 585
R377 B.n433 B.n28 585
R378 B.n306 B.n27 585
R379 B.n434 B.n27 585
R380 B.n305 B.n304 585
R381 B.n304 B.n23 585
R382 B.n303 B.n22 585
R383 B.n440 B.n22 585
R384 B.n302 B.n21 585
R385 B.n441 B.n21 585
R386 B.n301 B.n20 585
R387 B.n442 B.n20 585
R388 B.n300 B.n299 585
R389 B.n299 B.n16 585
R390 B.n298 B.n15 585
R391 B.n448 B.n15 585
R392 B.n297 B.n14 585
R393 B.n449 B.n14 585
R394 B.n296 B.n13 585
R395 B.n450 B.n13 585
R396 B.n295 B.n294 585
R397 B.n294 B.n12 585
R398 B.n293 B.n292 585
R399 B.n293 B.n8 585
R400 B.n291 B.n7 585
R401 B.n457 B.n7 585
R402 B.n290 B.n6 585
R403 B.n458 B.n6 585
R404 B.n289 B.n5 585
R405 B.n459 B.n5 585
R406 B.n288 B.n287 585
R407 B.n287 B.n4 585
R408 B.n286 B.n66 585
R409 B.n286 B.n285 585
R410 B.n275 B.n67 585
R411 B.n278 B.n67 585
R412 B.n277 B.n276 585
R413 B.n279 B.n277 585
R414 B.n274 B.n72 585
R415 B.n72 B.n71 585
R416 B.n273 B.n272 585
R417 B.n272 B.n271 585
R418 B.n74 B.n73 585
R419 B.n75 B.n74 585
R420 B.n264 B.n263 585
R421 B.n265 B.n264 585
R422 B.n262 B.n80 585
R423 B.n80 B.n79 585
R424 B.n261 B.n260 585
R425 B.n260 B.n259 585
R426 B.n82 B.n81 585
R427 B.n83 B.n82 585
R428 B.n252 B.n251 585
R429 B.n253 B.n252 585
R430 B.n250 B.n88 585
R431 B.n88 B.n87 585
R432 B.n249 B.n248 585
R433 B.n248 B.n247 585
R434 B.n244 B.n92 585
R435 B.n243 B.n242 585
R436 B.n240 B.n93 585
R437 B.n240 B.n91 585
R438 B.n239 B.n238 585
R439 B.n237 B.n236 585
R440 B.n235 B.n95 585
R441 B.n233 B.n232 585
R442 B.n231 B.n96 585
R443 B.n230 B.n229 585
R444 B.n227 B.n97 585
R445 B.n225 B.n224 585
R446 B.n223 B.n98 585
R447 B.n222 B.n221 585
R448 B.n219 B.n99 585
R449 B.n217 B.n216 585
R450 B.n215 B.n100 585
R451 B.n214 B.n213 585
R452 B.n211 B.n101 585
R453 B.n209 B.n208 585
R454 B.n207 B.n102 585
R455 B.n206 B.n205 585
R456 B.n203 B.n103 585
R457 B.n201 B.n200 585
R458 B.n199 B.n104 585
R459 B.n198 B.n197 585
R460 B.n195 B.n194 585
R461 B.n193 B.n192 585
R462 B.n191 B.n109 585
R463 B.n189 B.n188 585
R464 B.n187 B.n110 585
R465 B.n186 B.n185 585
R466 B.n183 B.n111 585
R467 B.n181 B.n180 585
R468 B.n179 B.n112 585
R469 B.n178 B.n177 585
R470 B.n175 B.n174 585
R471 B.n173 B.n172 585
R472 B.n171 B.n117 585
R473 B.n169 B.n168 585
R474 B.n167 B.n118 585
R475 B.n166 B.n165 585
R476 B.n163 B.n119 585
R477 B.n161 B.n160 585
R478 B.n159 B.n120 585
R479 B.n158 B.n157 585
R480 B.n155 B.n121 585
R481 B.n153 B.n152 585
R482 B.n151 B.n122 585
R483 B.n150 B.n149 585
R484 B.n147 B.n123 585
R485 B.n145 B.n144 585
R486 B.n143 B.n124 585
R487 B.n142 B.n141 585
R488 B.n139 B.n125 585
R489 B.n137 B.n136 585
R490 B.n135 B.n126 585
R491 B.n134 B.n133 585
R492 B.n131 B.n127 585
R493 B.n129 B.n128 585
R494 B.n90 B.n89 585
R495 B.n91 B.n90 585
R496 B.n246 B.n245 585
R497 B.n247 B.n246 585
R498 B.n86 B.n85 585
R499 B.n87 B.n86 585
R500 B.n255 B.n254 585
R501 B.n254 B.n253 585
R502 B.n256 B.n84 585
R503 B.n84 B.n83 585
R504 B.n258 B.n257 585
R505 B.n259 B.n258 585
R506 B.n78 B.n77 585
R507 B.n79 B.n78 585
R508 B.n267 B.n266 585
R509 B.n266 B.n265 585
R510 B.n268 B.n76 585
R511 B.n76 B.n75 585
R512 B.n270 B.n269 585
R513 B.n271 B.n270 585
R514 B.n70 B.n69 585
R515 B.n71 B.n70 585
R516 B.n281 B.n280 585
R517 B.n280 B.n279 585
R518 B.n282 B.n68 585
R519 B.n278 B.n68 585
R520 B.n284 B.n283 585
R521 B.n285 B.n284 585
R522 B.n3 B.n0 585
R523 B.n4 B.n3 585
R524 B.n456 B.n1 585
R525 B.n457 B.n456 585
R526 B.n455 B.n454 585
R527 B.n455 B.n8 585
R528 B.n453 B.n9 585
R529 B.n12 B.n9 585
R530 B.n452 B.n451 585
R531 B.n451 B.n450 585
R532 B.n11 B.n10 585
R533 B.n449 B.n11 585
R534 B.n447 B.n446 585
R535 B.n448 B.n447 585
R536 B.n445 B.n17 585
R537 B.n17 B.n16 585
R538 B.n444 B.n443 585
R539 B.n443 B.n442 585
R540 B.n19 B.n18 585
R541 B.n441 B.n19 585
R542 B.n439 B.n438 585
R543 B.n440 B.n439 585
R544 B.n437 B.n24 585
R545 B.n24 B.n23 585
R546 B.n436 B.n435 585
R547 B.n435 B.n434 585
R548 B.n26 B.n25 585
R549 B.n433 B.n26 585
R550 B.n431 B.n430 585
R551 B.n432 B.n431 585
R552 B.n460 B.n459 585
R553 B.n458 B.n2 585
R554 B.n431 B.n31 535.745
R555 B.n310 B.n29 535.745
R556 B.n248 B.n90 535.745
R557 B.n246 B.n92 535.745
R558 B.n44 B.t13 407.452
R559 B.n52 B.t6 407.452
R560 B.n113 B.t2 407.452
R561 B.n105 B.t10 407.452
R562 B.n311 B.n30 256.663
R563 B.n313 B.n30 256.663
R564 B.n319 B.n30 256.663
R565 B.n321 B.n30 256.663
R566 B.n327 B.n30 256.663
R567 B.n329 B.n30 256.663
R568 B.n335 B.n30 256.663
R569 B.n337 B.n30 256.663
R570 B.n343 B.n30 256.663
R571 B.n345 B.n30 256.663
R572 B.n351 B.n30 256.663
R573 B.n353 B.n30 256.663
R574 B.n359 B.n30 256.663
R575 B.n361 B.n30 256.663
R576 B.n367 B.n30 256.663
R577 B.n369 B.n30 256.663
R578 B.n375 B.n30 256.663
R579 B.n377 B.n30 256.663
R580 B.n384 B.n30 256.663
R581 B.n386 B.n30 256.663
R582 B.n392 B.n30 256.663
R583 B.n394 B.n30 256.663
R584 B.n400 B.n30 256.663
R585 B.n402 B.n30 256.663
R586 B.n408 B.n30 256.663
R587 B.n410 B.n30 256.663
R588 B.n416 B.n30 256.663
R589 B.n418 B.n30 256.663
R590 B.n424 B.n30 256.663
R591 B.n426 B.n30 256.663
R592 B.n241 B.n91 256.663
R593 B.n94 B.n91 256.663
R594 B.n234 B.n91 256.663
R595 B.n228 B.n91 256.663
R596 B.n226 B.n91 256.663
R597 B.n220 B.n91 256.663
R598 B.n218 B.n91 256.663
R599 B.n212 B.n91 256.663
R600 B.n210 B.n91 256.663
R601 B.n204 B.n91 256.663
R602 B.n202 B.n91 256.663
R603 B.n196 B.n91 256.663
R604 B.n108 B.n91 256.663
R605 B.n190 B.n91 256.663
R606 B.n184 B.n91 256.663
R607 B.n182 B.n91 256.663
R608 B.n176 B.n91 256.663
R609 B.n116 B.n91 256.663
R610 B.n170 B.n91 256.663
R611 B.n164 B.n91 256.663
R612 B.n162 B.n91 256.663
R613 B.n156 B.n91 256.663
R614 B.n154 B.n91 256.663
R615 B.n148 B.n91 256.663
R616 B.n146 B.n91 256.663
R617 B.n140 B.n91 256.663
R618 B.n138 B.n91 256.663
R619 B.n132 B.n91 256.663
R620 B.n130 B.n91 256.663
R621 B.n462 B.n461 256.663
R622 B.n52 B.t8 207.732
R623 B.n113 B.t5 207.732
R624 B.n44 B.t14 207.732
R625 B.n105 B.t12 207.732
R626 B.n53 B.t9 186.593
R627 B.n114 B.t4 186.593
R628 B.n45 B.t15 186.593
R629 B.n106 B.t11 186.593
R630 B.n427 B.n425 163.367
R631 B.n423 B.n33 163.367
R632 B.n419 B.n417 163.367
R633 B.n415 B.n35 163.367
R634 B.n411 B.n409 163.367
R635 B.n407 B.n37 163.367
R636 B.n403 B.n401 163.367
R637 B.n399 B.n39 163.367
R638 B.n395 B.n393 163.367
R639 B.n391 B.n41 163.367
R640 B.n387 B.n385 163.367
R641 B.n383 B.n43 163.367
R642 B.n378 B.n376 163.367
R643 B.n374 B.n47 163.367
R644 B.n370 B.n368 163.367
R645 B.n366 B.n49 163.367
R646 B.n362 B.n360 163.367
R647 B.n358 B.n51 163.367
R648 B.n354 B.n352 163.367
R649 B.n350 B.n56 163.367
R650 B.n346 B.n344 163.367
R651 B.n342 B.n58 163.367
R652 B.n338 B.n336 163.367
R653 B.n334 B.n60 163.367
R654 B.n330 B.n328 163.367
R655 B.n326 B.n62 163.367
R656 B.n322 B.n320 163.367
R657 B.n318 B.n64 163.367
R658 B.n314 B.n312 163.367
R659 B.n248 B.n88 163.367
R660 B.n252 B.n88 163.367
R661 B.n252 B.n82 163.367
R662 B.n260 B.n82 163.367
R663 B.n260 B.n80 163.367
R664 B.n264 B.n80 163.367
R665 B.n264 B.n74 163.367
R666 B.n272 B.n74 163.367
R667 B.n272 B.n72 163.367
R668 B.n277 B.n72 163.367
R669 B.n277 B.n67 163.367
R670 B.n286 B.n67 163.367
R671 B.n287 B.n286 163.367
R672 B.n287 B.n5 163.367
R673 B.n6 B.n5 163.367
R674 B.n7 B.n6 163.367
R675 B.n293 B.n7 163.367
R676 B.n294 B.n293 163.367
R677 B.n294 B.n13 163.367
R678 B.n14 B.n13 163.367
R679 B.n15 B.n14 163.367
R680 B.n299 B.n15 163.367
R681 B.n299 B.n20 163.367
R682 B.n21 B.n20 163.367
R683 B.n22 B.n21 163.367
R684 B.n304 B.n22 163.367
R685 B.n304 B.n27 163.367
R686 B.n28 B.n27 163.367
R687 B.n29 B.n28 163.367
R688 B.n242 B.n240 163.367
R689 B.n240 B.n239 163.367
R690 B.n236 B.n235 163.367
R691 B.n233 B.n96 163.367
R692 B.n229 B.n227 163.367
R693 B.n225 B.n98 163.367
R694 B.n221 B.n219 163.367
R695 B.n217 B.n100 163.367
R696 B.n213 B.n211 163.367
R697 B.n209 B.n102 163.367
R698 B.n205 B.n203 163.367
R699 B.n201 B.n104 163.367
R700 B.n197 B.n195 163.367
R701 B.n192 B.n191 163.367
R702 B.n189 B.n110 163.367
R703 B.n185 B.n183 163.367
R704 B.n181 B.n112 163.367
R705 B.n177 B.n175 163.367
R706 B.n172 B.n171 163.367
R707 B.n169 B.n118 163.367
R708 B.n165 B.n163 163.367
R709 B.n161 B.n120 163.367
R710 B.n157 B.n155 163.367
R711 B.n153 B.n122 163.367
R712 B.n149 B.n147 163.367
R713 B.n145 B.n124 163.367
R714 B.n141 B.n139 163.367
R715 B.n137 B.n126 163.367
R716 B.n133 B.n131 163.367
R717 B.n129 B.n90 163.367
R718 B.n246 B.n86 163.367
R719 B.n254 B.n86 163.367
R720 B.n254 B.n84 163.367
R721 B.n258 B.n84 163.367
R722 B.n258 B.n78 163.367
R723 B.n266 B.n78 163.367
R724 B.n266 B.n76 163.367
R725 B.n270 B.n76 163.367
R726 B.n270 B.n70 163.367
R727 B.n280 B.n70 163.367
R728 B.n280 B.n68 163.367
R729 B.n284 B.n68 163.367
R730 B.n284 B.n3 163.367
R731 B.n460 B.n3 163.367
R732 B.n456 B.n2 163.367
R733 B.n456 B.n455 163.367
R734 B.n455 B.n9 163.367
R735 B.n451 B.n9 163.367
R736 B.n451 B.n11 163.367
R737 B.n447 B.n11 163.367
R738 B.n447 B.n17 163.367
R739 B.n443 B.n17 163.367
R740 B.n443 B.n19 163.367
R741 B.n439 B.n19 163.367
R742 B.n439 B.n24 163.367
R743 B.n435 B.n24 163.367
R744 B.n435 B.n26 163.367
R745 B.n431 B.n26 163.367
R746 B.n247 B.n91 116.873
R747 B.n432 B.n30 116.873
R748 B.n426 B.n31 71.676
R749 B.n425 B.n424 71.676
R750 B.n418 B.n33 71.676
R751 B.n417 B.n416 71.676
R752 B.n410 B.n35 71.676
R753 B.n409 B.n408 71.676
R754 B.n402 B.n37 71.676
R755 B.n401 B.n400 71.676
R756 B.n394 B.n39 71.676
R757 B.n393 B.n392 71.676
R758 B.n386 B.n41 71.676
R759 B.n385 B.n384 71.676
R760 B.n377 B.n43 71.676
R761 B.n376 B.n375 71.676
R762 B.n369 B.n47 71.676
R763 B.n368 B.n367 71.676
R764 B.n361 B.n49 71.676
R765 B.n360 B.n359 71.676
R766 B.n353 B.n51 71.676
R767 B.n352 B.n351 71.676
R768 B.n345 B.n56 71.676
R769 B.n344 B.n343 71.676
R770 B.n337 B.n58 71.676
R771 B.n336 B.n335 71.676
R772 B.n329 B.n60 71.676
R773 B.n328 B.n327 71.676
R774 B.n321 B.n62 71.676
R775 B.n320 B.n319 71.676
R776 B.n313 B.n64 71.676
R777 B.n312 B.n311 71.676
R778 B.n311 B.n310 71.676
R779 B.n314 B.n313 71.676
R780 B.n319 B.n318 71.676
R781 B.n322 B.n321 71.676
R782 B.n327 B.n326 71.676
R783 B.n330 B.n329 71.676
R784 B.n335 B.n334 71.676
R785 B.n338 B.n337 71.676
R786 B.n343 B.n342 71.676
R787 B.n346 B.n345 71.676
R788 B.n351 B.n350 71.676
R789 B.n354 B.n353 71.676
R790 B.n359 B.n358 71.676
R791 B.n362 B.n361 71.676
R792 B.n367 B.n366 71.676
R793 B.n370 B.n369 71.676
R794 B.n375 B.n374 71.676
R795 B.n378 B.n377 71.676
R796 B.n384 B.n383 71.676
R797 B.n387 B.n386 71.676
R798 B.n392 B.n391 71.676
R799 B.n395 B.n394 71.676
R800 B.n400 B.n399 71.676
R801 B.n403 B.n402 71.676
R802 B.n408 B.n407 71.676
R803 B.n411 B.n410 71.676
R804 B.n416 B.n415 71.676
R805 B.n419 B.n418 71.676
R806 B.n424 B.n423 71.676
R807 B.n427 B.n426 71.676
R808 B.n241 B.n92 71.676
R809 B.n239 B.n94 71.676
R810 B.n235 B.n234 71.676
R811 B.n228 B.n96 71.676
R812 B.n227 B.n226 71.676
R813 B.n220 B.n98 71.676
R814 B.n219 B.n218 71.676
R815 B.n212 B.n100 71.676
R816 B.n211 B.n210 71.676
R817 B.n204 B.n102 71.676
R818 B.n203 B.n202 71.676
R819 B.n196 B.n104 71.676
R820 B.n195 B.n108 71.676
R821 B.n191 B.n190 71.676
R822 B.n184 B.n110 71.676
R823 B.n183 B.n182 71.676
R824 B.n176 B.n112 71.676
R825 B.n175 B.n116 71.676
R826 B.n171 B.n170 71.676
R827 B.n164 B.n118 71.676
R828 B.n163 B.n162 71.676
R829 B.n156 B.n120 71.676
R830 B.n155 B.n154 71.676
R831 B.n148 B.n122 71.676
R832 B.n147 B.n146 71.676
R833 B.n140 B.n124 71.676
R834 B.n139 B.n138 71.676
R835 B.n132 B.n126 71.676
R836 B.n131 B.n130 71.676
R837 B.n242 B.n241 71.676
R838 B.n236 B.n94 71.676
R839 B.n234 B.n233 71.676
R840 B.n229 B.n228 71.676
R841 B.n226 B.n225 71.676
R842 B.n221 B.n220 71.676
R843 B.n218 B.n217 71.676
R844 B.n213 B.n212 71.676
R845 B.n210 B.n209 71.676
R846 B.n205 B.n204 71.676
R847 B.n202 B.n201 71.676
R848 B.n197 B.n196 71.676
R849 B.n192 B.n108 71.676
R850 B.n190 B.n189 71.676
R851 B.n185 B.n184 71.676
R852 B.n182 B.n181 71.676
R853 B.n177 B.n176 71.676
R854 B.n172 B.n116 71.676
R855 B.n170 B.n169 71.676
R856 B.n165 B.n164 71.676
R857 B.n162 B.n161 71.676
R858 B.n157 B.n156 71.676
R859 B.n154 B.n153 71.676
R860 B.n149 B.n148 71.676
R861 B.n146 B.n145 71.676
R862 B.n141 B.n140 71.676
R863 B.n138 B.n137 71.676
R864 B.n133 B.n132 71.676
R865 B.n130 B.n129 71.676
R866 B.n461 B.n460 71.676
R867 B.n461 B.n2 71.676
R868 B.n247 B.n87 63.5789
R869 B.n253 B.n87 63.5789
R870 B.n253 B.n83 63.5789
R871 B.n259 B.n83 63.5789
R872 B.n265 B.n79 63.5789
R873 B.n265 B.n75 63.5789
R874 B.n271 B.n75 63.5789
R875 B.n271 B.n71 63.5789
R876 B.n279 B.n71 63.5789
R877 B.n279 B.n278 63.5789
R878 B.n285 B.n4 63.5789
R879 B.n459 B.n4 63.5789
R880 B.n459 B.n458 63.5789
R881 B.n458 B.n457 63.5789
R882 B.n457 B.n8 63.5789
R883 B.n450 B.n12 63.5789
R884 B.n450 B.n449 63.5789
R885 B.n449 B.n448 63.5789
R886 B.n448 B.n16 63.5789
R887 B.n442 B.n16 63.5789
R888 B.n442 B.n441 63.5789
R889 B.n440 B.n23 63.5789
R890 B.n434 B.n23 63.5789
R891 B.n434 B.n433 63.5789
R892 B.n433 B.n432 63.5789
R893 B.n380 B.n45 59.5399
R894 B.n54 B.n53 59.5399
R895 B.n115 B.n114 59.5399
R896 B.n107 B.n106 59.5399
R897 B.n259 B.t3 56.0991
R898 B.t7 B.n440 56.0991
R899 B.n285 B.t0 44.8794
R900 B.t1 B.n8 44.8794
R901 B.n245 B.n244 34.8103
R902 B.n249 B.n89 34.8103
R903 B.n309 B.n308 34.8103
R904 B.n430 B.n429 34.8103
R905 B.n45 B.n44 21.1399
R906 B.n53 B.n52 21.1399
R907 B.n114 B.n113 21.1399
R908 B.n106 B.n105 21.1399
R909 B.n278 B.t0 18.7
R910 B.n12 B.t1 18.7
R911 B B.n462 18.0485
R912 B.n245 B.n85 10.6151
R913 B.n255 B.n85 10.6151
R914 B.n256 B.n255 10.6151
R915 B.n257 B.n256 10.6151
R916 B.n257 B.n77 10.6151
R917 B.n267 B.n77 10.6151
R918 B.n268 B.n267 10.6151
R919 B.n269 B.n268 10.6151
R920 B.n269 B.n69 10.6151
R921 B.n281 B.n69 10.6151
R922 B.n282 B.n281 10.6151
R923 B.n283 B.n282 10.6151
R924 B.n283 B.n0 10.6151
R925 B.n244 B.n243 10.6151
R926 B.n243 B.n93 10.6151
R927 B.n238 B.n93 10.6151
R928 B.n238 B.n237 10.6151
R929 B.n237 B.n95 10.6151
R930 B.n232 B.n95 10.6151
R931 B.n232 B.n231 10.6151
R932 B.n231 B.n230 10.6151
R933 B.n230 B.n97 10.6151
R934 B.n224 B.n97 10.6151
R935 B.n224 B.n223 10.6151
R936 B.n223 B.n222 10.6151
R937 B.n222 B.n99 10.6151
R938 B.n216 B.n99 10.6151
R939 B.n216 B.n215 10.6151
R940 B.n215 B.n214 10.6151
R941 B.n214 B.n101 10.6151
R942 B.n208 B.n101 10.6151
R943 B.n208 B.n207 10.6151
R944 B.n207 B.n206 10.6151
R945 B.n206 B.n103 10.6151
R946 B.n200 B.n103 10.6151
R947 B.n200 B.n199 10.6151
R948 B.n199 B.n198 10.6151
R949 B.n194 B.n193 10.6151
R950 B.n193 B.n109 10.6151
R951 B.n188 B.n109 10.6151
R952 B.n188 B.n187 10.6151
R953 B.n187 B.n186 10.6151
R954 B.n186 B.n111 10.6151
R955 B.n180 B.n111 10.6151
R956 B.n180 B.n179 10.6151
R957 B.n179 B.n178 10.6151
R958 B.n174 B.n173 10.6151
R959 B.n173 B.n117 10.6151
R960 B.n168 B.n117 10.6151
R961 B.n168 B.n167 10.6151
R962 B.n167 B.n166 10.6151
R963 B.n166 B.n119 10.6151
R964 B.n160 B.n119 10.6151
R965 B.n160 B.n159 10.6151
R966 B.n159 B.n158 10.6151
R967 B.n158 B.n121 10.6151
R968 B.n152 B.n121 10.6151
R969 B.n152 B.n151 10.6151
R970 B.n151 B.n150 10.6151
R971 B.n150 B.n123 10.6151
R972 B.n144 B.n123 10.6151
R973 B.n144 B.n143 10.6151
R974 B.n143 B.n142 10.6151
R975 B.n142 B.n125 10.6151
R976 B.n136 B.n125 10.6151
R977 B.n136 B.n135 10.6151
R978 B.n135 B.n134 10.6151
R979 B.n134 B.n127 10.6151
R980 B.n128 B.n127 10.6151
R981 B.n128 B.n89 10.6151
R982 B.n250 B.n249 10.6151
R983 B.n251 B.n250 10.6151
R984 B.n251 B.n81 10.6151
R985 B.n261 B.n81 10.6151
R986 B.n262 B.n261 10.6151
R987 B.n263 B.n262 10.6151
R988 B.n263 B.n73 10.6151
R989 B.n273 B.n73 10.6151
R990 B.n274 B.n273 10.6151
R991 B.n276 B.n274 10.6151
R992 B.n276 B.n275 10.6151
R993 B.n275 B.n66 10.6151
R994 B.n288 B.n66 10.6151
R995 B.n289 B.n288 10.6151
R996 B.n290 B.n289 10.6151
R997 B.n291 B.n290 10.6151
R998 B.n292 B.n291 10.6151
R999 B.n295 B.n292 10.6151
R1000 B.n296 B.n295 10.6151
R1001 B.n297 B.n296 10.6151
R1002 B.n298 B.n297 10.6151
R1003 B.n300 B.n298 10.6151
R1004 B.n301 B.n300 10.6151
R1005 B.n302 B.n301 10.6151
R1006 B.n303 B.n302 10.6151
R1007 B.n305 B.n303 10.6151
R1008 B.n306 B.n305 10.6151
R1009 B.n307 B.n306 10.6151
R1010 B.n308 B.n307 10.6151
R1011 B.n454 B.n1 10.6151
R1012 B.n454 B.n453 10.6151
R1013 B.n453 B.n452 10.6151
R1014 B.n452 B.n10 10.6151
R1015 B.n446 B.n10 10.6151
R1016 B.n446 B.n445 10.6151
R1017 B.n445 B.n444 10.6151
R1018 B.n444 B.n18 10.6151
R1019 B.n438 B.n18 10.6151
R1020 B.n438 B.n437 10.6151
R1021 B.n437 B.n436 10.6151
R1022 B.n436 B.n25 10.6151
R1023 B.n430 B.n25 10.6151
R1024 B.n429 B.n428 10.6151
R1025 B.n428 B.n32 10.6151
R1026 B.n422 B.n32 10.6151
R1027 B.n422 B.n421 10.6151
R1028 B.n421 B.n420 10.6151
R1029 B.n420 B.n34 10.6151
R1030 B.n414 B.n34 10.6151
R1031 B.n414 B.n413 10.6151
R1032 B.n413 B.n412 10.6151
R1033 B.n412 B.n36 10.6151
R1034 B.n406 B.n36 10.6151
R1035 B.n406 B.n405 10.6151
R1036 B.n405 B.n404 10.6151
R1037 B.n404 B.n38 10.6151
R1038 B.n398 B.n38 10.6151
R1039 B.n398 B.n397 10.6151
R1040 B.n397 B.n396 10.6151
R1041 B.n396 B.n40 10.6151
R1042 B.n390 B.n40 10.6151
R1043 B.n390 B.n389 10.6151
R1044 B.n389 B.n388 10.6151
R1045 B.n388 B.n42 10.6151
R1046 B.n382 B.n42 10.6151
R1047 B.n382 B.n381 10.6151
R1048 B.n379 B.n46 10.6151
R1049 B.n373 B.n46 10.6151
R1050 B.n373 B.n372 10.6151
R1051 B.n372 B.n371 10.6151
R1052 B.n371 B.n48 10.6151
R1053 B.n365 B.n48 10.6151
R1054 B.n365 B.n364 10.6151
R1055 B.n364 B.n363 10.6151
R1056 B.n363 B.n50 10.6151
R1057 B.n357 B.n356 10.6151
R1058 B.n356 B.n355 10.6151
R1059 B.n355 B.n55 10.6151
R1060 B.n349 B.n55 10.6151
R1061 B.n349 B.n348 10.6151
R1062 B.n348 B.n347 10.6151
R1063 B.n347 B.n57 10.6151
R1064 B.n341 B.n57 10.6151
R1065 B.n341 B.n340 10.6151
R1066 B.n340 B.n339 10.6151
R1067 B.n339 B.n59 10.6151
R1068 B.n333 B.n59 10.6151
R1069 B.n333 B.n332 10.6151
R1070 B.n332 B.n331 10.6151
R1071 B.n331 B.n61 10.6151
R1072 B.n325 B.n61 10.6151
R1073 B.n325 B.n324 10.6151
R1074 B.n324 B.n323 10.6151
R1075 B.n323 B.n63 10.6151
R1076 B.n317 B.n63 10.6151
R1077 B.n317 B.n316 10.6151
R1078 B.n316 B.n315 10.6151
R1079 B.n315 B.n65 10.6151
R1080 B.n309 B.n65 10.6151
R1081 B.n198 B.n107 8.74196
R1082 B.n174 B.n115 8.74196
R1083 B.n381 B.n380 8.74196
R1084 B.n357 B.n54 8.74196
R1085 B.n462 B.n0 8.11757
R1086 B.n462 B.n1 8.11757
R1087 B.t3 B.n79 7.48031
R1088 B.n441 B.t7 7.48031
R1089 B.n194 B.n107 1.87367
R1090 B.n178 B.n115 1.87367
R1091 B.n380 B.n379 1.87367
R1092 B.n54 B.n50 1.87367
R1093 VP.n0 VP.t1 454.075
R1094 VP.n0 VP.t0 418.473
R1095 VP VP.n0 0.0516364
R1096 VDD1.n32 VDD1.n31 289.615
R1097 VDD1.n65 VDD1.n64 289.615
R1098 VDD1.n31 VDD1.n30 185
R1099 VDD1.n2 VDD1.n1 185
R1100 VDD1.n25 VDD1.n24 185
R1101 VDD1.n23 VDD1.n22 185
R1102 VDD1.n6 VDD1.n5 185
R1103 VDD1.n17 VDD1.n16 185
R1104 VDD1.n15 VDD1.n14 185
R1105 VDD1.n10 VDD1.n9 185
R1106 VDD1.n43 VDD1.n42 185
R1107 VDD1.n48 VDD1.n47 185
R1108 VDD1.n50 VDD1.n49 185
R1109 VDD1.n39 VDD1.n38 185
R1110 VDD1.n56 VDD1.n55 185
R1111 VDD1.n58 VDD1.n57 185
R1112 VDD1.n35 VDD1.n34 185
R1113 VDD1.n64 VDD1.n63 185
R1114 VDD1.n11 VDD1.t0 149.525
R1115 VDD1.n44 VDD1.t1 149.525
R1116 VDD1.n31 VDD1.n1 104.615
R1117 VDD1.n24 VDD1.n1 104.615
R1118 VDD1.n24 VDD1.n23 104.615
R1119 VDD1.n23 VDD1.n5 104.615
R1120 VDD1.n16 VDD1.n5 104.615
R1121 VDD1.n16 VDD1.n15 104.615
R1122 VDD1.n15 VDD1.n9 104.615
R1123 VDD1.n48 VDD1.n42 104.615
R1124 VDD1.n49 VDD1.n48 104.615
R1125 VDD1.n49 VDD1.n38 104.615
R1126 VDD1.n56 VDD1.n38 104.615
R1127 VDD1.n57 VDD1.n56 104.615
R1128 VDD1.n57 VDD1.n34 104.615
R1129 VDD1.n64 VDD1.n34 104.615
R1130 VDD1 VDD1.n65 82.5029
R1131 VDD1.t0 VDD1.n9 52.3082
R1132 VDD1.t1 VDD1.n42 52.3082
R1133 VDD1 VDD1.n32 50.9027
R1134 VDD1.n30 VDD1.n0 12.8005
R1135 VDD1.n63 VDD1.n33 12.8005
R1136 VDD1.n29 VDD1.n2 12.0247
R1137 VDD1.n62 VDD1.n35 12.0247
R1138 VDD1.n26 VDD1.n25 11.249
R1139 VDD1.n59 VDD1.n58 11.249
R1140 VDD1.n22 VDD1.n4 10.4732
R1141 VDD1.n55 VDD1.n37 10.4732
R1142 VDD1.n11 VDD1.n10 10.2746
R1143 VDD1.n44 VDD1.n43 10.2746
R1144 VDD1.n21 VDD1.n6 9.69747
R1145 VDD1.n54 VDD1.n39 9.69747
R1146 VDD1.n28 VDD1.n0 9.45567
R1147 VDD1.n61 VDD1.n33 9.45567
R1148 VDD1.n29 VDD1.n28 9.3005
R1149 VDD1.n27 VDD1.n26 9.3005
R1150 VDD1.n4 VDD1.n3 9.3005
R1151 VDD1.n21 VDD1.n20 9.3005
R1152 VDD1.n19 VDD1.n18 9.3005
R1153 VDD1.n8 VDD1.n7 9.3005
R1154 VDD1.n13 VDD1.n12 9.3005
R1155 VDD1.n46 VDD1.n45 9.3005
R1156 VDD1.n41 VDD1.n40 9.3005
R1157 VDD1.n52 VDD1.n51 9.3005
R1158 VDD1.n54 VDD1.n53 9.3005
R1159 VDD1.n37 VDD1.n36 9.3005
R1160 VDD1.n60 VDD1.n59 9.3005
R1161 VDD1.n62 VDD1.n61 9.3005
R1162 VDD1.n18 VDD1.n17 8.92171
R1163 VDD1.n51 VDD1.n50 8.92171
R1164 VDD1.n14 VDD1.n8 8.14595
R1165 VDD1.n47 VDD1.n41 8.14595
R1166 VDD1.n13 VDD1.n10 7.3702
R1167 VDD1.n46 VDD1.n43 7.3702
R1168 VDD1.n14 VDD1.n13 5.81868
R1169 VDD1.n47 VDD1.n46 5.81868
R1170 VDD1.n17 VDD1.n8 5.04292
R1171 VDD1.n50 VDD1.n41 5.04292
R1172 VDD1.n18 VDD1.n6 4.26717
R1173 VDD1.n51 VDD1.n39 4.26717
R1174 VDD1.n22 VDD1.n21 3.49141
R1175 VDD1.n55 VDD1.n54 3.49141
R1176 VDD1.n12 VDD1.n11 2.84308
R1177 VDD1.n45 VDD1.n44 2.84308
R1178 VDD1.n25 VDD1.n4 2.71565
R1179 VDD1.n58 VDD1.n37 2.71565
R1180 VDD1.n26 VDD1.n2 1.93989
R1181 VDD1.n59 VDD1.n35 1.93989
R1182 VDD1.n30 VDD1.n29 1.16414
R1183 VDD1.n63 VDD1.n62 1.16414
R1184 VDD1.n32 VDD1.n0 0.388379
R1185 VDD1.n65 VDD1.n33 0.388379
R1186 VDD1.n28 VDD1.n27 0.155672
R1187 VDD1.n27 VDD1.n3 0.155672
R1188 VDD1.n20 VDD1.n3 0.155672
R1189 VDD1.n20 VDD1.n19 0.155672
R1190 VDD1.n19 VDD1.n7 0.155672
R1191 VDD1.n12 VDD1.n7 0.155672
R1192 VDD1.n45 VDD1.n40 0.155672
R1193 VDD1.n52 VDD1.n40 0.155672
R1194 VDD1.n53 VDD1.n52 0.155672
R1195 VDD1.n53 VDD1.n36 0.155672
R1196 VDD1.n60 VDD1.n36 0.155672
R1197 VDD1.n61 VDD1.n60 0.155672
C0 VDD1 VTAIL 3.5753f
C1 VDD1 VN 0.148616f
C2 VP VTAIL 1.0152f
C3 VN VP 3.56481f
C4 VN VTAIL 1.00084f
C5 VDD1 VDD2 0.466442f
C6 VP VDD2 0.256669f
C7 VTAIL VDD2 3.61276f
C8 VN VDD2 1.21258f
C9 VDD1 VP 1.31825f
C10 VDD2 B 2.764505f
C11 VDD1 B 4.23975f
C12 VTAIL B 4.196293f
C13 VN B 6.12019f
C14 VP B 3.670115f
C15 VDD1.n0 B 0.008682f
C16 VDD1.n1 B 0.019631f
C17 VDD1.n2 B 0.008794f
C18 VDD1.n3 B 0.015456f
C19 VDD1.n4 B 0.008305f
C20 VDD1.n5 B 0.019631f
C21 VDD1.n6 B 0.008794f
C22 VDD1.n7 B 0.015456f
C23 VDD1.n8 B 0.008305f
C24 VDD1.n9 B 0.014723f
C25 VDD1.n10 B 0.013877f
C26 VDD1.t0 B 0.032731f
C27 VDD1.n11 B 0.078685f
C28 VDD1.n12 B 0.399468f
C29 VDD1.n13 B 0.008305f
C30 VDD1.n14 B 0.008794f
C31 VDD1.n15 B 0.019631f
C32 VDD1.n16 B 0.019631f
C33 VDD1.n17 B 0.008794f
C34 VDD1.n18 B 0.008305f
C35 VDD1.n19 B 0.015456f
C36 VDD1.n20 B 0.015456f
C37 VDD1.n21 B 0.008305f
C38 VDD1.n22 B 0.008794f
C39 VDD1.n23 B 0.019631f
C40 VDD1.n24 B 0.019631f
C41 VDD1.n25 B 0.008794f
C42 VDD1.n26 B 0.008305f
C43 VDD1.n27 B 0.015456f
C44 VDD1.n28 B 0.038049f
C45 VDD1.n29 B 0.008305f
C46 VDD1.n30 B 0.008794f
C47 VDD1.n31 B 0.038625f
C48 VDD1.n32 B 0.042806f
C49 VDD1.n33 B 0.008682f
C50 VDD1.n34 B 0.019631f
C51 VDD1.n35 B 0.008794f
C52 VDD1.n36 B 0.015456f
C53 VDD1.n37 B 0.008305f
C54 VDD1.n38 B 0.019631f
C55 VDD1.n39 B 0.008794f
C56 VDD1.n40 B 0.015456f
C57 VDD1.n41 B 0.008305f
C58 VDD1.n42 B 0.014723f
C59 VDD1.n43 B 0.013877f
C60 VDD1.t1 B 0.032731f
C61 VDD1.n44 B 0.078685f
C62 VDD1.n45 B 0.399468f
C63 VDD1.n46 B 0.008305f
C64 VDD1.n47 B 0.008794f
C65 VDD1.n48 B 0.019631f
C66 VDD1.n49 B 0.019631f
C67 VDD1.n50 B 0.008794f
C68 VDD1.n51 B 0.008305f
C69 VDD1.n52 B 0.015456f
C70 VDD1.n53 B 0.015456f
C71 VDD1.n54 B 0.008305f
C72 VDD1.n55 B 0.008794f
C73 VDD1.n56 B 0.019631f
C74 VDD1.n57 B 0.019631f
C75 VDD1.n58 B 0.008794f
C76 VDD1.n59 B 0.008305f
C77 VDD1.n60 B 0.015456f
C78 VDD1.n61 B 0.038049f
C79 VDD1.n62 B 0.008305f
C80 VDD1.n63 B 0.008794f
C81 VDD1.n64 B 0.038625f
C82 VDD1.n65 B 0.296869f
C83 VP.t1 B 0.671342f
C84 VP.t0 B 0.576825f
C85 VP.n0 B 2.33848f
C86 VDD2.n0 B 0.008822f
C87 VDD2.n1 B 0.019947f
C88 VDD2.n2 B 0.008936f
C89 VDD2.n3 B 0.015705f
C90 VDD2.n4 B 0.008439f
C91 VDD2.n5 B 0.019947f
C92 VDD2.n6 B 0.008936f
C93 VDD2.n7 B 0.015705f
C94 VDD2.n8 B 0.008439f
C95 VDD2.n9 B 0.01496f
C96 VDD2.n10 B 0.014101f
C97 VDD2.t0 B 0.033258f
C98 VDD2.n11 B 0.079953f
C99 VDD2.n12 B 0.405904f
C100 VDD2.n13 B 0.008439f
C101 VDD2.n14 B 0.008936f
C102 VDD2.n15 B 0.019947f
C103 VDD2.n16 B 0.019947f
C104 VDD2.n17 B 0.008936f
C105 VDD2.n18 B 0.008439f
C106 VDD2.n19 B 0.015705f
C107 VDD2.n20 B 0.015705f
C108 VDD2.n21 B 0.008439f
C109 VDD2.n22 B 0.008936f
C110 VDD2.n23 B 0.019947f
C111 VDD2.n24 B 0.019947f
C112 VDD2.n25 B 0.008936f
C113 VDD2.n26 B 0.008439f
C114 VDD2.n27 B 0.015705f
C115 VDD2.n28 B 0.038662f
C116 VDD2.n29 B 0.008439f
C117 VDD2.n30 B 0.008936f
C118 VDD2.n31 B 0.039248f
C119 VDD2.n32 B 0.282964f
C120 VDD2.n33 B 0.008822f
C121 VDD2.n34 B 0.019947f
C122 VDD2.n35 B 0.008936f
C123 VDD2.n36 B 0.015705f
C124 VDD2.n37 B 0.008439f
C125 VDD2.n38 B 0.019947f
C126 VDD2.n39 B 0.008936f
C127 VDD2.n40 B 0.015705f
C128 VDD2.n41 B 0.008439f
C129 VDD2.n42 B 0.01496f
C130 VDD2.n43 B 0.014101f
C131 VDD2.t1 B 0.033258f
C132 VDD2.n44 B 0.079953f
C133 VDD2.n45 B 0.405904f
C134 VDD2.n46 B 0.008439f
C135 VDD2.n47 B 0.008936f
C136 VDD2.n48 B 0.019947f
C137 VDD2.n49 B 0.019947f
C138 VDD2.n50 B 0.008936f
C139 VDD2.n51 B 0.008439f
C140 VDD2.n52 B 0.015705f
C141 VDD2.n53 B 0.015705f
C142 VDD2.n54 B 0.008439f
C143 VDD2.n55 B 0.008936f
C144 VDD2.n56 B 0.019947f
C145 VDD2.n57 B 0.019947f
C146 VDD2.n58 B 0.008936f
C147 VDD2.n59 B 0.008439f
C148 VDD2.n60 B 0.015705f
C149 VDD2.n61 B 0.038662f
C150 VDD2.n62 B 0.008439f
C151 VDD2.n63 B 0.008936f
C152 VDD2.n64 B 0.039248f
C153 VDD2.n65 B 0.04323f
C154 VDD2.n66 B 1.32527f
C155 VTAIL.n0 B 0.009821f
C156 VTAIL.n1 B 0.022205f
C157 VTAIL.n2 B 0.009947f
C158 VTAIL.n3 B 0.017483f
C159 VTAIL.n4 B 0.009394f
C160 VTAIL.n5 B 0.022205f
C161 VTAIL.n6 B 0.009947f
C162 VTAIL.n7 B 0.017483f
C163 VTAIL.n8 B 0.009394f
C164 VTAIL.n9 B 0.016654f
C165 VTAIL.n10 B 0.015697f
C166 VTAIL.t0 B 0.037022f
C167 VTAIL.n11 B 0.089002f
C168 VTAIL.n12 B 0.451843f
C169 VTAIL.n13 B 0.009394f
C170 VTAIL.n14 B 0.009947f
C171 VTAIL.n15 B 0.022205f
C172 VTAIL.n16 B 0.022205f
C173 VTAIL.n17 B 0.009947f
C174 VTAIL.n18 B 0.009394f
C175 VTAIL.n19 B 0.017483f
C176 VTAIL.n20 B 0.017483f
C177 VTAIL.n21 B 0.009394f
C178 VTAIL.n22 B 0.009947f
C179 VTAIL.n23 B 0.022205f
C180 VTAIL.n24 B 0.022205f
C181 VTAIL.n25 B 0.009947f
C182 VTAIL.n26 B 0.009394f
C183 VTAIL.n27 B 0.017483f
C184 VTAIL.n28 B 0.043037f
C185 VTAIL.n29 B 0.009394f
C186 VTAIL.n30 B 0.009947f
C187 VTAIL.n31 B 0.04369f
C188 VTAIL.n32 B 0.036068f
C189 VTAIL.n33 B 0.717645f
C190 VTAIL.n34 B 0.009821f
C191 VTAIL.n35 B 0.022205f
C192 VTAIL.n36 B 0.009947f
C193 VTAIL.n37 B 0.017483f
C194 VTAIL.n38 B 0.009394f
C195 VTAIL.n39 B 0.022205f
C196 VTAIL.n40 B 0.009947f
C197 VTAIL.n41 B 0.017483f
C198 VTAIL.n42 B 0.009394f
C199 VTAIL.n43 B 0.016654f
C200 VTAIL.n44 B 0.015697f
C201 VTAIL.t2 B 0.037022f
C202 VTAIL.n45 B 0.089002f
C203 VTAIL.n46 B 0.451843f
C204 VTAIL.n47 B 0.009394f
C205 VTAIL.n48 B 0.009947f
C206 VTAIL.n49 B 0.022205f
C207 VTAIL.n50 B 0.022205f
C208 VTAIL.n51 B 0.009947f
C209 VTAIL.n52 B 0.009394f
C210 VTAIL.n53 B 0.017483f
C211 VTAIL.n54 B 0.017483f
C212 VTAIL.n55 B 0.009394f
C213 VTAIL.n56 B 0.009947f
C214 VTAIL.n57 B 0.022205f
C215 VTAIL.n58 B 0.022205f
C216 VTAIL.n59 B 0.009947f
C217 VTAIL.n60 B 0.009394f
C218 VTAIL.n61 B 0.017483f
C219 VTAIL.n62 B 0.043037f
C220 VTAIL.n63 B 0.009394f
C221 VTAIL.n64 B 0.009947f
C222 VTAIL.n65 B 0.04369f
C223 VTAIL.n66 B 0.036068f
C224 VTAIL.n67 B 0.727601f
C225 VTAIL.n68 B 0.009821f
C226 VTAIL.n69 B 0.022205f
C227 VTAIL.n70 B 0.009947f
C228 VTAIL.n71 B 0.017483f
C229 VTAIL.n72 B 0.009394f
C230 VTAIL.n73 B 0.022205f
C231 VTAIL.n74 B 0.009947f
C232 VTAIL.n75 B 0.017483f
C233 VTAIL.n76 B 0.009394f
C234 VTAIL.n77 B 0.016654f
C235 VTAIL.n78 B 0.015697f
C236 VTAIL.t1 B 0.037022f
C237 VTAIL.n79 B 0.089002f
C238 VTAIL.n80 B 0.451843f
C239 VTAIL.n81 B 0.009394f
C240 VTAIL.n82 B 0.009947f
C241 VTAIL.n83 B 0.022205f
C242 VTAIL.n84 B 0.022205f
C243 VTAIL.n85 B 0.009947f
C244 VTAIL.n86 B 0.009394f
C245 VTAIL.n87 B 0.017483f
C246 VTAIL.n88 B 0.017483f
C247 VTAIL.n89 B 0.009394f
C248 VTAIL.n90 B 0.009947f
C249 VTAIL.n91 B 0.022205f
C250 VTAIL.n92 B 0.022205f
C251 VTAIL.n93 B 0.009947f
C252 VTAIL.n94 B 0.009394f
C253 VTAIL.n95 B 0.017483f
C254 VTAIL.n96 B 0.043037f
C255 VTAIL.n97 B 0.009394f
C256 VTAIL.n98 B 0.009947f
C257 VTAIL.n99 B 0.04369f
C258 VTAIL.n100 B 0.036068f
C259 VTAIL.n101 B 0.674667f
C260 VTAIL.n102 B 0.009821f
C261 VTAIL.n103 B 0.022205f
C262 VTAIL.n104 B 0.009947f
C263 VTAIL.n105 B 0.017483f
C264 VTAIL.n106 B 0.009394f
C265 VTAIL.n107 B 0.022205f
C266 VTAIL.n108 B 0.009947f
C267 VTAIL.n109 B 0.017483f
C268 VTAIL.n110 B 0.009394f
C269 VTAIL.n111 B 0.016654f
C270 VTAIL.n112 B 0.015697f
C271 VTAIL.t3 B 0.037022f
C272 VTAIL.n113 B 0.089002f
C273 VTAIL.n114 B 0.451843f
C274 VTAIL.n115 B 0.009394f
C275 VTAIL.n116 B 0.009947f
C276 VTAIL.n117 B 0.022205f
C277 VTAIL.n118 B 0.022205f
C278 VTAIL.n119 B 0.009947f
C279 VTAIL.n120 B 0.009394f
C280 VTAIL.n121 B 0.017483f
C281 VTAIL.n122 B 0.017483f
C282 VTAIL.n123 B 0.009394f
C283 VTAIL.n124 B 0.009947f
C284 VTAIL.n125 B 0.022205f
C285 VTAIL.n126 B 0.022205f
C286 VTAIL.n127 B 0.009947f
C287 VTAIL.n128 B 0.009394f
C288 VTAIL.n129 B 0.017483f
C289 VTAIL.n130 B 0.043037f
C290 VTAIL.n131 B 0.009394f
C291 VTAIL.n132 B 0.009947f
C292 VTAIL.n133 B 0.04369f
C293 VTAIL.n134 B 0.036068f
C294 VTAIL.n135 B 0.631689f
C295 VN.t1 B 0.569143f
C296 VN.t0 B 0.665094f
.ends

