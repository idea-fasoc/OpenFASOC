* NGSPICE file created from diff_pair_sample_0253.ext - technology: sky130A

.subckt diff_pair_sample_0253 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n2746_n2548# sky130_fd_pr__pfet_01v8 ad=3.081 pd=16.58 as=0 ps=0 w=7.9 l=1.15
X1 VDD2.t9 VN.t0 VTAIL.t13 w_n2746_n2548# sky130_fd_pr__pfet_01v8 ad=3.081 pd=16.58 as=1.3035 ps=8.23 w=7.9 l=1.15
X2 VTAIL.t3 VP.t0 VDD1.t9 w_n2746_n2548# sky130_fd_pr__pfet_01v8 ad=1.3035 pd=8.23 as=1.3035 ps=8.23 w=7.9 l=1.15
X3 VDD2.t8 VN.t1 VTAIL.t14 w_n2746_n2548# sky130_fd_pr__pfet_01v8 ad=3.081 pd=16.58 as=1.3035 ps=8.23 w=7.9 l=1.15
X4 VDD2.t7 VN.t2 VTAIL.t15 w_n2746_n2548# sky130_fd_pr__pfet_01v8 ad=1.3035 pd=8.23 as=1.3035 ps=8.23 w=7.9 l=1.15
X5 B.t8 B.t6 B.t7 w_n2746_n2548# sky130_fd_pr__pfet_01v8 ad=3.081 pd=16.58 as=0 ps=0 w=7.9 l=1.15
X6 VDD2.t6 VN.t3 VTAIL.t10 w_n2746_n2548# sky130_fd_pr__pfet_01v8 ad=1.3035 pd=8.23 as=1.3035 ps=8.23 w=7.9 l=1.15
X7 B.t5 B.t3 B.t4 w_n2746_n2548# sky130_fd_pr__pfet_01v8 ad=3.081 pd=16.58 as=0 ps=0 w=7.9 l=1.15
X8 VDD2.t5 VN.t4 VTAIL.t16 w_n2746_n2548# sky130_fd_pr__pfet_01v8 ad=1.3035 pd=8.23 as=3.081 ps=16.58 w=7.9 l=1.15
X9 VTAIL.t17 VN.t5 VDD2.t4 w_n2746_n2548# sky130_fd_pr__pfet_01v8 ad=1.3035 pd=8.23 as=1.3035 ps=8.23 w=7.9 l=1.15
X10 VTAIL.t18 VN.t6 VDD2.t3 w_n2746_n2548# sky130_fd_pr__pfet_01v8 ad=1.3035 pd=8.23 as=1.3035 ps=8.23 w=7.9 l=1.15
X11 VTAIL.t2 VP.t1 VDD1.t8 w_n2746_n2548# sky130_fd_pr__pfet_01v8 ad=1.3035 pd=8.23 as=1.3035 ps=8.23 w=7.9 l=1.15
X12 VDD2.t2 VN.t7 VTAIL.t11 w_n2746_n2548# sky130_fd_pr__pfet_01v8 ad=1.3035 pd=8.23 as=3.081 ps=16.58 w=7.9 l=1.15
X13 VDD1.t7 VP.t2 VTAIL.t1 w_n2746_n2548# sky130_fd_pr__pfet_01v8 ad=1.3035 pd=8.23 as=3.081 ps=16.58 w=7.9 l=1.15
X14 VTAIL.t7 VP.t3 VDD1.t6 w_n2746_n2548# sky130_fd_pr__pfet_01v8 ad=1.3035 pd=8.23 as=1.3035 ps=8.23 w=7.9 l=1.15
X15 B.t2 B.t0 B.t1 w_n2746_n2548# sky130_fd_pr__pfet_01v8 ad=3.081 pd=16.58 as=0 ps=0 w=7.9 l=1.15
X16 VDD1.t5 VP.t4 VTAIL.t6 w_n2746_n2548# sky130_fd_pr__pfet_01v8 ad=1.3035 pd=8.23 as=3.081 ps=16.58 w=7.9 l=1.15
X17 VDD1.t4 VP.t5 VTAIL.t9 w_n2746_n2548# sky130_fd_pr__pfet_01v8 ad=3.081 pd=16.58 as=1.3035 ps=8.23 w=7.9 l=1.15
X18 VTAIL.t12 VN.t8 VDD2.t1 w_n2746_n2548# sky130_fd_pr__pfet_01v8 ad=1.3035 pd=8.23 as=1.3035 ps=8.23 w=7.9 l=1.15
X19 VDD1.t3 VP.t6 VTAIL.t4 w_n2746_n2548# sky130_fd_pr__pfet_01v8 ad=1.3035 pd=8.23 as=1.3035 ps=8.23 w=7.9 l=1.15
X20 VDD1.t2 VP.t7 VTAIL.t5 w_n2746_n2548# sky130_fd_pr__pfet_01v8 ad=1.3035 pd=8.23 as=1.3035 ps=8.23 w=7.9 l=1.15
X21 VTAIL.t19 VN.t9 VDD2.t0 w_n2746_n2548# sky130_fd_pr__pfet_01v8 ad=1.3035 pd=8.23 as=1.3035 ps=8.23 w=7.9 l=1.15
X22 VTAIL.t8 VP.t8 VDD1.t1 w_n2746_n2548# sky130_fd_pr__pfet_01v8 ad=1.3035 pd=8.23 as=1.3035 ps=8.23 w=7.9 l=1.15
X23 VDD1.t0 VP.t9 VTAIL.t0 w_n2746_n2548# sky130_fd_pr__pfet_01v8 ad=3.081 pd=16.58 as=1.3035 ps=8.23 w=7.9 l=1.15
R0 B.n407 B.n406 585
R1 B.n408 B.n57 585
R2 B.n410 B.n409 585
R3 B.n411 B.n56 585
R4 B.n413 B.n412 585
R5 B.n414 B.n55 585
R6 B.n416 B.n415 585
R7 B.n417 B.n54 585
R8 B.n419 B.n418 585
R9 B.n420 B.n53 585
R10 B.n422 B.n421 585
R11 B.n423 B.n52 585
R12 B.n425 B.n424 585
R13 B.n426 B.n51 585
R14 B.n428 B.n427 585
R15 B.n429 B.n50 585
R16 B.n431 B.n430 585
R17 B.n432 B.n49 585
R18 B.n434 B.n433 585
R19 B.n435 B.n48 585
R20 B.n437 B.n436 585
R21 B.n438 B.n47 585
R22 B.n440 B.n439 585
R23 B.n441 B.n46 585
R24 B.n443 B.n442 585
R25 B.n444 B.n45 585
R26 B.n446 B.n445 585
R27 B.n447 B.n44 585
R28 B.n449 B.n448 585
R29 B.n450 B.n41 585
R30 B.n453 B.n452 585
R31 B.n454 B.n40 585
R32 B.n456 B.n455 585
R33 B.n457 B.n39 585
R34 B.n459 B.n458 585
R35 B.n460 B.n38 585
R36 B.n462 B.n461 585
R37 B.n463 B.n37 585
R38 B.n465 B.n464 585
R39 B.n467 B.n466 585
R40 B.n468 B.n33 585
R41 B.n470 B.n469 585
R42 B.n471 B.n32 585
R43 B.n473 B.n472 585
R44 B.n474 B.n31 585
R45 B.n476 B.n475 585
R46 B.n477 B.n30 585
R47 B.n479 B.n478 585
R48 B.n480 B.n29 585
R49 B.n482 B.n481 585
R50 B.n483 B.n28 585
R51 B.n485 B.n484 585
R52 B.n486 B.n27 585
R53 B.n488 B.n487 585
R54 B.n489 B.n26 585
R55 B.n491 B.n490 585
R56 B.n492 B.n25 585
R57 B.n494 B.n493 585
R58 B.n495 B.n24 585
R59 B.n497 B.n496 585
R60 B.n498 B.n23 585
R61 B.n500 B.n499 585
R62 B.n501 B.n22 585
R63 B.n503 B.n502 585
R64 B.n504 B.n21 585
R65 B.n506 B.n505 585
R66 B.n507 B.n20 585
R67 B.n509 B.n508 585
R68 B.n510 B.n19 585
R69 B.n405 B.n58 585
R70 B.n404 B.n403 585
R71 B.n402 B.n59 585
R72 B.n401 B.n400 585
R73 B.n399 B.n60 585
R74 B.n398 B.n397 585
R75 B.n396 B.n61 585
R76 B.n395 B.n394 585
R77 B.n393 B.n62 585
R78 B.n392 B.n391 585
R79 B.n390 B.n63 585
R80 B.n389 B.n388 585
R81 B.n387 B.n64 585
R82 B.n386 B.n385 585
R83 B.n384 B.n65 585
R84 B.n383 B.n382 585
R85 B.n381 B.n66 585
R86 B.n380 B.n379 585
R87 B.n378 B.n67 585
R88 B.n377 B.n376 585
R89 B.n375 B.n68 585
R90 B.n374 B.n373 585
R91 B.n372 B.n69 585
R92 B.n371 B.n370 585
R93 B.n369 B.n70 585
R94 B.n368 B.n367 585
R95 B.n366 B.n71 585
R96 B.n365 B.n364 585
R97 B.n363 B.n72 585
R98 B.n362 B.n361 585
R99 B.n360 B.n73 585
R100 B.n359 B.n358 585
R101 B.n357 B.n74 585
R102 B.n356 B.n355 585
R103 B.n354 B.n75 585
R104 B.n353 B.n352 585
R105 B.n351 B.n76 585
R106 B.n350 B.n349 585
R107 B.n348 B.n77 585
R108 B.n347 B.n346 585
R109 B.n345 B.n78 585
R110 B.n344 B.n343 585
R111 B.n342 B.n79 585
R112 B.n341 B.n340 585
R113 B.n339 B.n80 585
R114 B.n338 B.n337 585
R115 B.n336 B.n81 585
R116 B.n335 B.n334 585
R117 B.n333 B.n82 585
R118 B.n332 B.n331 585
R119 B.n330 B.n83 585
R120 B.n329 B.n328 585
R121 B.n327 B.n84 585
R122 B.n326 B.n325 585
R123 B.n324 B.n85 585
R124 B.n323 B.n322 585
R125 B.n321 B.n86 585
R126 B.n320 B.n319 585
R127 B.n318 B.n87 585
R128 B.n317 B.n316 585
R129 B.n315 B.n88 585
R130 B.n314 B.n313 585
R131 B.n312 B.n89 585
R132 B.n311 B.n310 585
R133 B.n309 B.n90 585
R134 B.n308 B.n307 585
R135 B.n306 B.n91 585
R136 B.n305 B.n304 585
R137 B.n303 B.n92 585
R138 B.n198 B.n131 585
R139 B.n200 B.n199 585
R140 B.n201 B.n130 585
R141 B.n203 B.n202 585
R142 B.n204 B.n129 585
R143 B.n206 B.n205 585
R144 B.n207 B.n128 585
R145 B.n209 B.n208 585
R146 B.n210 B.n127 585
R147 B.n212 B.n211 585
R148 B.n213 B.n126 585
R149 B.n215 B.n214 585
R150 B.n216 B.n125 585
R151 B.n218 B.n217 585
R152 B.n219 B.n124 585
R153 B.n221 B.n220 585
R154 B.n222 B.n123 585
R155 B.n224 B.n223 585
R156 B.n225 B.n122 585
R157 B.n227 B.n226 585
R158 B.n228 B.n121 585
R159 B.n230 B.n229 585
R160 B.n231 B.n120 585
R161 B.n233 B.n232 585
R162 B.n234 B.n119 585
R163 B.n236 B.n235 585
R164 B.n237 B.n118 585
R165 B.n239 B.n238 585
R166 B.n240 B.n117 585
R167 B.n242 B.n241 585
R168 B.n244 B.n243 585
R169 B.n245 B.n113 585
R170 B.n247 B.n246 585
R171 B.n248 B.n112 585
R172 B.n250 B.n249 585
R173 B.n251 B.n111 585
R174 B.n253 B.n252 585
R175 B.n254 B.n110 585
R176 B.n256 B.n255 585
R177 B.n258 B.n107 585
R178 B.n260 B.n259 585
R179 B.n261 B.n106 585
R180 B.n263 B.n262 585
R181 B.n264 B.n105 585
R182 B.n266 B.n265 585
R183 B.n267 B.n104 585
R184 B.n269 B.n268 585
R185 B.n270 B.n103 585
R186 B.n272 B.n271 585
R187 B.n273 B.n102 585
R188 B.n275 B.n274 585
R189 B.n276 B.n101 585
R190 B.n278 B.n277 585
R191 B.n279 B.n100 585
R192 B.n281 B.n280 585
R193 B.n282 B.n99 585
R194 B.n284 B.n283 585
R195 B.n285 B.n98 585
R196 B.n287 B.n286 585
R197 B.n288 B.n97 585
R198 B.n290 B.n289 585
R199 B.n291 B.n96 585
R200 B.n293 B.n292 585
R201 B.n294 B.n95 585
R202 B.n296 B.n295 585
R203 B.n297 B.n94 585
R204 B.n299 B.n298 585
R205 B.n300 B.n93 585
R206 B.n302 B.n301 585
R207 B.n197 B.n196 585
R208 B.n195 B.n132 585
R209 B.n194 B.n193 585
R210 B.n192 B.n133 585
R211 B.n191 B.n190 585
R212 B.n189 B.n134 585
R213 B.n188 B.n187 585
R214 B.n186 B.n135 585
R215 B.n185 B.n184 585
R216 B.n183 B.n136 585
R217 B.n182 B.n181 585
R218 B.n180 B.n137 585
R219 B.n179 B.n178 585
R220 B.n177 B.n138 585
R221 B.n176 B.n175 585
R222 B.n174 B.n139 585
R223 B.n173 B.n172 585
R224 B.n171 B.n140 585
R225 B.n170 B.n169 585
R226 B.n168 B.n141 585
R227 B.n167 B.n166 585
R228 B.n165 B.n142 585
R229 B.n164 B.n163 585
R230 B.n162 B.n143 585
R231 B.n161 B.n160 585
R232 B.n159 B.n144 585
R233 B.n158 B.n157 585
R234 B.n156 B.n145 585
R235 B.n155 B.n154 585
R236 B.n153 B.n146 585
R237 B.n152 B.n151 585
R238 B.n150 B.n147 585
R239 B.n149 B.n148 585
R240 B.n2 B.n0 585
R241 B.n561 B.n1 585
R242 B.n560 B.n559 585
R243 B.n558 B.n3 585
R244 B.n557 B.n556 585
R245 B.n555 B.n4 585
R246 B.n554 B.n553 585
R247 B.n552 B.n5 585
R248 B.n551 B.n550 585
R249 B.n549 B.n6 585
R250 B.n548 B.n547 585
R251 B.n546 B.n7 585
R252 B.n545 B.n544 585
R253 B.n543 B.n8 585
R254 B.n542 B.n541 585
R255 B.n540 B.n9 585
R256 B.n539 B.n538 585
R257 B.n537 B.n10 585
R258 B.n536 B.n535 585
R259 B.n534 B.n11 585
R260 B.n533 B.n532 585
R261 B.n531 B.n12 585
R262 B.n530 B.n529 585
R263 B.n528 B.n13 585
R264 B.n527 B.n526 585
R265 B.n525 B.n14 585
R266 B.n524 B.n523 585
R267 B.n522 B.n15 585
R268 B.n521 B.n520 585
R269 B.n519 B.n16 585
R270 B.n518 B.n517 585
R271 B.n516 B.n17 585
R272 B.n515 B.n514 585
R273 B.n513 B.n18 585
R274 B.n512 B.n511 585
R275 B.n563 B.n562 585
R276 B.n196 B.n131 511.721
R277 B.n512 B.n19 511.721
R278 B.n303 B.n302 511.721
R279 B.n406 B.n405 511.721
R280 B.n108 B.t0 369.404
R281 B.n114 B.t9 369.404
R282 B.n34 B.t6 369.404
R283 B.n42 B.t3 369.404
R284 B.n108 B.t2 330.454
R285 B.n42 B.t4 330.454
R286 B.n114 B.t11 330.454
R287 B.n34 B.t7 330.454
R288 B.n109 B.t1 301.75
R289 B.n43 B.t5 301.75
R290 B.n115 B.t10 301.75
R291 B.n35 B.t8 301.75
R292 B.n196 B.n195 163.367
R293 B.n195 B.n194 163.367
R294 B.n194 B.n133 163.367
R295 B.n190 B.n133 163.367
R296 B.n190 B.n189 163.367
R297 B.n189 B.n188 163.367
R298 B.n188 B.n135 163.367
R299 B.n184 B.n135 163.367
R300 B.n184 B.n183 163.367
R301 B.n183 B.n182 163.367
R302 B.n182 B.n137 163.367
R303 B.n178 B.n137 163.367
R304 B.n178 B.n177 163.367
R305 B.n177 B.n176 163.367
R306 B.n176 B.n139 163.367
R307 B.n172 B.n139 163.367
R308 B.n172 B.n171 163.367
R309 B.n171 B.n170 163.367
R310 B.n170 B.n141 163.367
R311 B.n166 B.n141 163.367
R312 B.n166 B.n165 163.367
R313 B.n165 B.n164 163.367
R314 B.n164 B.n143 163.367
R315 B.n160 B.n143 163.367
R316 B.n160 B.n159 163.367
R317 B.n159 B.n158 163.367
R318 B.n158 B.n145 163.367
R319 B.n154 B.n145 163.367
R320 B.n154 B.n153 163.367
R321 B.n153 B.n152 163.367
R322 B.n152 B.n147 163.367
R323 B.n148 B.n147 163.367
R324 B.n148 B.n2 163.367
R325 B.n562 B.n2 163.367
R326 B.n562 B.n561 163.367
R327 B.n561 B.n560 163.367
R328 B.n560 B.n3 163.367
R329 B.n556 B.n3 163.367
R330 B.n556 B.n555 163.367
R331 B.n555 B.n554 163.367
R332 B.n554 B.n5 163.367
R333 B.n550 B.n5 163.367
R334 B.n550 B.n549 163.367
R335 B.n549 B.n548 163.367
R336 B.n548 B.n7 163.367
R337 B.n544 B.n7 163.367
R338 B.n544 B.n543 163.367
R339 B.n543 B.n542 163.367
R340 B.n542 B.n9 163.367
R341 B.n538 B.n9 163.367
R342 B.n538 B.n537 163.367
R343 B.n537 B.n536 163.367
R344 B.n536 B.n11 163.367
R345 B.n532 B.n11 163.367
R346 B.n532 B.n531 163.367
R347 B.n531 B.n530 163.367
R348 B.n530 B.n13 163.367
R349 B.n526 B.n13 163.367
R350 B.n526 B.n525 163.367
R351 B.n525 B.n524 163.367
R352 B.n524 B.n15 163.367
R353 B.n520 B.n15 163.367
R354 B.n520 B.n519 163.367
R355 B.n519 B.n518 163.367
R356 B.n518 B.n17 163.367
R357 B.n514 B.n17 163.367
R358 B.n514 B.n513 163.367
R359 B.n513 B.n512 163.367
R360 B.n200 B.n131 163.367
R361 B.n201 B.n200 163.367
R362 B.n202 B.n201 163.367
R363 B.n202 B.n129 163.367
R364 B.n206 B.n129 163.367
R365 B.n207 B.n206 163.367
R366 B.n208 B.n207 163.367
R367 B.n208 B.n127 163.367
R368 B.n212 B.n127 163.367
R369 B.n213 B.n212 163.367
R370 B.n214 B.n213 163.367
R371 B.n214 B.n125 163.367
R372 B.n218 B.n125 163.367
R373 B.n219 B.n218 163.367
R374 B.n220 B.n219 163.367
R375 B.n220 B.n123 163.367
R376 B.n224 B.n123 163.367
R377 B.n225 B.n224 163.367
R378 B.n226 B.n225 163.367
R379 B.n226 B.n121 163.367
R380 B.n230 B.n121 163.367
R381 B.n231 B.n230 163.367
R382 B.n232 B.n231 163.367
R383 B.n232 B.n119 163.367
R384 B.n236 B.n119 163.367
R385 B.n237 B.n236 163.367
R386 B.n238 B.n237 163.367
R387 B.n238 B.n117 163.367
R388 B.n242 B.n117 163.367
R389 B.n243 B.n242 163.367
R390 B.n243 B.n113 163.367
R391 B.n247 B.n113 163.367
R392 B.n248 B.n247 163.367
R393 B.n249 B.n248 163.367
R394 B.n249 B.n111 163.367
R395 B.n253 B.n111 163.367
R396 B.n254 B.n253 163.367
R397 B.n255 B.n254 163.367
R398 B.n255 B.n107 163.367
R399 B.n260 B.n107 163.367
R400 B.n261 B.n260 163.367
R401 B.n262 B.n261 163.367
R402 B.n262 B.n105 163.367
R403 B.n266 B.n105 163.367
R404 B.n267 B.n266 163.367
R405 B.n268 B.n267 163.367
R406 B.n268 B.n103 163.367
R407 B.n272 B.n103 163.367
R408 B.n273 B.n272 163.367
R409 B.n274 B.n273 163.367
R410 B.n274 B.n101 163.367
R411 B.n278 B.n101 163.367
R412 B.n279 B.n278 163.367
R413 B.n280 B.n279 163.367
R414 B.n280 B.n99 163.367
R415 B.n284 B.n99 163.367
R416 B.n285 B.n284 163.367
R417 B.n286 B.n285 163.367
R418 B.n286 B.n97 163.367
R419 B.n290 B.n97 163.367
R420 B.n291 B.n290 163.367
R421 B.n292 B.n291 163.367
R422 B.n292 B.n95 163.367
R423 B.n296 B.n95 163.367
R424 B.n297 B.n296 163.367
R425 B.n298 B.n297 163.367
R426 B.n298 B.n93 163.367
R427 B.n302 B.n93 163.367
R428 B.n304 B.n303 163.367
R429 B.n304 B.n91 163.367
R430 B.n308 B.n91 163.367
R431 B.n309 B.n308 163.367
R432 B.n310 B.n309 163.367
R433 B.n310 B.n89 163.367
R434 B.n314 B.n89 163.367
R435 B.n315 B.n314 163.367
R436 B.n316 B.n315 163.367
R437 B.n316 B.n87 163.367
R438 B.n320 B.n87 163.367
R439 B.n321 B.n320 163.367
R440 B.n322 B.n321 163.367
R441 B.n322 B.n85 163.367
R442 B.n326 B.n85 163.367
R443 B.n327 B.n326 163.367
R444 B.n328 B.n327 163.367
R445 B.n328 B.n83 163.367
R446 B.n332 B.n83 163.367
R447 B.n333 B.n332 163.367
R448 B.n334 B.n333 163.367
R449 B.n334 B.n81 163.367
R450 B.n338 B.n81 163.367
R451 B.n339 B.n338 163.367
R452 B.n340 B.n339 163.367
R453 B.n340 B.n79 163.367
R454 B.n344 B.n79 163.367
R455 B.n345 B.n344 163.367
R456 B.n346 B.n345 163.367
R457 B.n346 B.n77 163.367
R458 B.n350 B.n77 163.367
R459 B.n351 B.n350 163.367
R460 B.n352 B.n351 163.367
R461 B.n352 B.n75 163.367
R462 B.n356 B.n75 163.367
R463 B.n357 B.n356 163.367
R464 B.n358 B.n357 163.367
R465 B.n358 B.n73 163.367
R466 B.n362 B.n73 163.367
R467 B.n363 B.n362 163.367
R468 B.n364 B.n363 163.367
R469 B.n364 B.n71 163.367
R470 B.n368 B.n71 163.367
R471 B.n369 B.n368 163.367
R472 B.n370 B.n369 163.367
R473 B.n370 B.n69 163.367
R474 B.n374 B.n69 163.367
R475 B.n375 B.n374 163.367
R476 B.n376 B.n375 163.367
R477 B.n376 B.n67 163.367
R478 B.n380 B.n67 163.367
R479 B.n381 B.n380 163.367
R480 B.n382 B.n381 163.367
R481 B.n382 B.n65 163.367
R482 B.n386 B.n65 163.367
R483 B.n387 B.n386 163.367
R484 B.n388 B.n387 163.367
R485 B.n388 B.n63 163.367
R486 B.n392 B.n63 163.367
R487 B.n393 B.n392 163.367
R488 B.n394 B.n393 163.367
R489 B.n394 B.n61 163.367
R490 B.n398 B.n61 163.367
R491 B.n399 B.n398 163.367
R492 B.n400 B.n399 163.367
R493 B.n400 B.n59 163.367
R494 B.n404 B.n59 163.367
R495 B.n405 B.n404 163.367
R496 B.n508 B.n19 163.367
R497 B.n508 B.n507 163.367
R498 B.n507 B.n506 163.367
R499 B.n506 B.n21 163.367
R500 B.n502 B.n21 163.367
R501 B.n502 B.n501 163.367
R502 B.n501 B.n500 163.367
R503 B.n500 B.n23 163.367
R504 B.n496 B.n23 163.367
R505 B.n496 B.n495 163.367
R506 B.n495 B.n494 163.367
R507 B.n494 B.n25 163.367
R508 B.n490 B.n25 163.367
R509 B.n490 B.n489 163.367
R510 B.n489 B.n488 163.367
R511 B.n488 B.n27 163.367
R512 B.n484 B.n27 163.367
R513 B.n484 B.n483 163.367
R514 B.n483 B.n482 163.367
R515 B.n482 B.n29 163.367
R516 B.n478 B.n29 163.367
R517 B.n478 B.n477 163.367
R518 B.n477 B.n476 163.367
R519 B.n476 B.n31 163.367
R520 B.n472 B.n31 163.367
R521 B.n472 B.n471 163.367
R522 B.n471 B.n470 163.367
R523 B.n470 B.n33 163.367
R524 B.n466 B.n33 163.367
R525 B.n466 B.n465 163.367
R526 B.n465 B.n37 163.367
R527 B.n461 B.n37 163.367
R528 B.n461 B.n460 163.367
R529 B.n460 B.n459 163.367
R530 B.n459 B.n39 163.367
R531 B.n455 B.n39 163.367
R532 B.n455 B.n454 163.367
R533 B.n454 B.n453 163.367
R534 B.n453 B.n41 163.367
R535 B.n448 B.n41 163.367
R536 B.n448 B.n447 163.367
R537 B.n447 B.n446 163.367
R538 B.n446 B.n45 163.367
R539 B.n442 B.n45 163.367
R540 B.n442 B.n441 163.367
R541 B.n441 B.n440 163.367
R542 B.n440 B.n47 163.367
R543 B.n436 B.n47 163.367
R544 B.n436 B.n435 163.367
R545 B.n435 B.n434 163.367
R546 B.n434 B.n49 163.367
R547 B.n430 B.n49 163.367
R548 B.n430 B.n429 163.367
R549 B.n429 B.n428 163.367
R550 B.n428 B.n51 163.367
R551 B.n424 B.n51 163.367
R552 B.n424 B.n423 163.367
R553 B.n423 B.n422 163.367
R554 B.n422 B.n53 163.367
R555 B.n418 B.n53 163.367
R556 B.n418 B.n417 163.367
R557 B.n417 B.n416 163.367
R558 B.n416 B.n55 163.367
R559 B.n412 B.n55 163.367
R560 B.n412 B.n411 163.367
R561 B.n411 B.n410 163.367
R562 B.n410 B.n57 163.367
R563 B.n406 B.n57 163.367
R564 B.n257 B.n109 59.5399
R565 B.n116 B.n115 59.5399
R566 B.n36 B.n35 59.5399
R567 B.n451 B.n43 59.5399
R568 B.n511 B.n510 33.2493
R569 B.n407 B.n58 33.2493
R570 B.n301 B.n92 33.2493
R571 B.n198 B.n197 33.2493
R572 B.n109 B.n108 28.7035
R573 B.n115 B.n114 28.7035
R574 B.n35 B.n34 28.7035
R575 B.n43 B.n42 28.7035
R576 B B.n563 18.0485
R577 B.n510 B.n509 10.6151
R578 B.n509 B.n20 10.6151
R579 B.n505 B.n20 10.6151
R580 B.n505 B.n504 10.6151
R581 B.n504 B.n503 10.6151
R582 B.n503 B.n22 10.6151
R583 B.n499 B.n22 10.6151
R584 B.n499 B.n498 10.6151
R585 B.n498 B.n497 10.6151
R586 B.n497 B.n24 10.6151
R587 B.n493 B.n24 10.6151
R588 B.n493 B.n492 10.6151
R589 B.n492 B.n491 10.6151
R590 B.n491 B.n26 10.6151
R591 B.n487 B.n26 10.6151
R592 B.n487 B.n486 10.6151
R593 B.n486 B.n485 10.6151
R594 B.n485 B.n28 10.6151
R595 B.n481 B.n28 10.6151
R596 B.n481 B.n480 10.6151
R597 B.n480 B.n479 10.6151
R598 B.n479 B.n30 10.6151
R599 B.n475 B.n30 10.6151
R600 B.n475 B.n474 10.6151
R601 B.n474 B.n473 10.6151
R602 B.n473 B.n32 10.6151
R603 B.n469 B.n32 10.6151
R604 B.n469 B.n468 10.6151
R605 B.n468 B.n467 10.6151
R606 B.n464 B.n463 10.6151
R607 B.n463 B.n462 10.6151
R608 B.n462 B.n38 10.6151
R609 B.n458 B.n38 10.6151
R610 B.n458 B.n457 10.6151
R611 B.n457 B.n456 10.6151
R612 B.n456 B.n40 10.6151
R613 B.n452 B.n40 10.6151
R614 B.n450 B.n449 10.6151
R615 B.n449 B.n44 10.6151
R616 B.n445 B.n44 10.6151
R617 B.n445 B.n444 10.6151
R618 B.n444 B.n443 10.6151
R619 B.n443 B.n46 10.6151
R620 B.n439 B.n46 10.6151
R621 B.n439 B.n438 10.6151
R622 B.n438 B.n437 10.6151
R623 B.n437 B.n48 10.6151
R624 B.n433 B.n48 10.6151
R625 B.n433 B.n432 10.6151
R626 B.n432 B.n431 10.6151
R627 B.n431 B.n50 10.6151
R628 B.n427 B.n50 10.6151
R629 B.n427 B.n426 10.6151
R630 B.n426 B.n425 10.6151
R631 B.n425 B.n52 10.6151
R632 B.n421 B.n52 10.6151
R633 B.n421 B.n420 10.6151
R634 B.n420 B.n419 10.6151
R635 B.n419 B.n54 10.6151
R636 B.n415 B.n54 10.6151
R637 B.n415 B.n414 10.6151
R638 B.n414 B.n413 10.6151
R639 B.n413 B.n56 10.6151
R640 B.n409 B.n56 10.6151
R641 B.n409 B.n408 10.6151
R642 B.n408 B.n407 10.6151
R643 B.n305 B.n92 10.6151
R644 B.n306 B.n305 10.6151
R645 B.n307 B.n306 10.6151
R646 B.n307 B.n90 10.6151
R647 B.n311 B.n90 10.6151
R648 B.n312 B.n311 10.6151
R649 B.n313 B.n312 10.6151
R650 B.n313 B.n88 10.6151
R651 B.n317 B.n88 10.6151
R652 B.n318 B.n317 10.6151
R653 B.n319 B.n318 10.6151
R654 B.n319 B.n86 10.6151
R655 B.n323 B.n86 10.6151
R656 B.n324 B.n323 10.6151
R657 B.n325 B.n324 10.6151
R658 B.n325 B.n84 10.6151
R659 B.n329 B.n84 10.6151
R660 B.n330 B.n329 10.6151
R661 B.n331 B.n330 10.6151
R662 B.n331 B.n82 10.6151
R663 B.n335 B.n82 10.6151
R664 B.n336 B.n335 10.6151
R665 B.n337 B.n336 10.6151
R666 B.n337 B.n80 10.6151
R667 B.n341 B.n80 10.6151
R668 B.n342 B.n341 10.6151
R669 B.n343 B.n342 10.6151
R670 B.n343 B.n78 10.6151
R671 B.n347 B.n78 10.6151
R672 B.n348 B.n347 10.6151
R673 B.n349 B.n348 10.6151
R674 B.n349 B.n76 10.6151
R675 B.n353 B.n76 10.6151
R676 B.n354 B.n353 10.6151
R677 B.n355 B.n354 10.6151
R678 B.n355 B.n74 10.6151
R679 B.n359 B.n74 10.6151
R680 B.n360 B.n359 10.6151
R681 B.n361 B.n360 10.6151
R682 B.n361 B.n72 10.6151
R683 B.n365 B.n72 10.6151
R684 B.n366 B.n365 10.6151
R685 B.n367 B.n366 10.6151
R686 B.n367 B.n70 10.6151
R687 B.n371 B.n70 10.6151
R688 B.n372 B.n371 10.6151
R689 B.n373 B.n372 10.6151
R690 B.n373 B.n68 10.6151
R691 B.n377 B.n68 10.6151
R692 B.n378 B.n377 10.6151
R693 B.n379 B.n378 10.6151
R694 B.n379 B.n66 10.6151
R695 B.n383 B.n66 10.6151
R696 B.n384 B.n383 10.6151
R697 B.n385 B.n384 10.6151
R698 B.n385 B.n64 10.6151
R699 B.n389 B.n64 10.6151
R700 B.n390 B.n389 10.6151
R701 B.n391 B.n390 10.6151
R702 B.n391 B.n62 10.6151
R703 B.n395 B.n62 10.6151
R704 B.n396 B.n395 10.6151
R705 B.n397 B.n396 10.6151
R706 B.n397 B.n60 10.6151
R707 B.n401 B.n60 10.6151
R708 B.n402 B.n401 10.6151
R709 B.n403 B.n402 10.6151
R710 B.n403 B.n58 10.6151
R711 B.n199 B.n198 10.6151
R712 B.n199 B.n130 10.6151
R713 B.n203 B.n130 10.6151
R714 B.n204 B.n203 10.6151
R715 B.n205 B.n204 10.6151
R716 B.n205 B.n128 10.6151
R717 B.n209 B.n128 10.6151
R718 B.n210 B.n209 10.6151
R719 B.n211 B.n210 10.6151
R720 B.n211 B.n126 10.6151
R721 B.n215 B.n126 10.6151
R722 B.n216 B.n215 10.6151
R723 B.n217 B.n216 10.6151
R724 B.n217 B.n124 10.6151
R725 B.n221 B.n124 10.6151
R726 B.n222 B.n221 10.6151
R727 B.n223 B.n222 10.6151
R728 B.n223 B.n122 10.6151
R729 B.n227 B.n122 10.6151
R730 B.n228 B.n227 10.6151
R731 B.n229 B.n228 10.6151
R732 B.n229 B.n120 10.6151
R733 B.n233 B.n120 10.6151
R734 B.n234 B.n233 10.6151
R735 B.n235 B.n234 10.6151
R736 B.n235 B.n118 10.6151
R737 B.n239 B.n118 10.6151
R738 B.n240 B.n239 10.6151
R739 B.n241 B.n240 10.6151
R740 B.n245 B.n244 10.6151
R741 B.n246 B.n245 10.6151
R742 B.n246 B.n112 10.6151
R743 B.n250 B.n112 10.6151
R744 B.n251 B.n250 10.6151
R745 B.n252 B.n251 10.6151
R746 B.n252 B.n110 10.6151
R747 B.n256 B.n110 10.6151
R748 B.n259 B.n258 10.6151
R749 B.n259 B.n106 10.6151
R750 B.n263 B.n106 10.6151
R751 B.n264 B.n263 10.6151
R752 B.n265 B.n264 10.6151
R753 B.n265 B.n104 10.6151
R754 B.n269 B.n104 10.6151
R755 B.n270 B.n269 10.6151
R756 B.n271 B.n270 10.6151
R757 B.n271 B.n102 10.6151
R758 B.n275 B.n102 10.6151
R759 B.n276 B.n275 10.6151
R760 B.n277 B.n276 10.6151
R761 B.n277 B.n100 10.6151
R762 B.n281 B.n100 10.6151
R763 B.n282 B.n281 10.6151
R764 B.n283 B.n282 10.6151
R765 B.n283 B.n98 10.6151
R766 B.n287 B.n98 10.6151
R767 B.n288 B.n287 10.6151
R768 B.n289 B.n288 10.6151
R769 B.n289 B.n96 10.6151
R770 B.n293 B.n96 10.6151
R771 B.n294 B.n293 10.6151
R772 B.n295 B.n294 10.6151
R773 B.n295 B.n94 10.6151
R774 B.n299 B.n94 10.6151
R775 B.n300 B.n299 10.6151
R776 B.n301 B.n300 10.6151
R777 B.n197 B.n132 10.6151
R778 B.n193 B.n132 10.6151
R779 B.n193 B.n192 10.6151
R780 B.n192 B.n191 10.6151
R781 B.n191 B.n134 10.6151
R782 B.n187 B.n134 10.6151
R783 B.n187 B.n186 10.6151
R784 B.n186 B.n185 10.6151
R785 B.n185 B.n136 10.6151
R786 B.n181 B.n136 10.6151
R787 B.n181 B.n180 10.6151
R788 B.n180 B.n179 10.6151
R789 B.n179 B.n138 10.6151
R790 B.n175 B.n138 10.6151
R791 B.n175 B.n174 10.6151
R792 B.n174 B.n173 10.6151
R793 B.n173 B.n140 10.6151
R794 B.n169 B.n140 10.6151
R795 B.n169 B.n168 10.6151
R796 B.n168 B.n167 10.6151
R797 B.n167 B.n142 10.6151
R798 B.n163 B.n142 10.6151
R799 B.n163 B.n162 10.6151
R800 B.n162 B.n161 10.6151
R801 B.n161 B.n144 10.6151
R802 B.n157 B.n144 10.6151
R803 B.n157 B.n156 10.6151
R804 B.n156 B.n155 10.6151
R805 B.n155 B.n146 10.6151
R806 B.n151 B.n146 10.6151
R807 B.n151 B.n150 10.6151
R808 B.n150 B.n149 10.6151
R809 B.n149 B.n0 10.6151
R810 B.n559 B.n1 10.6151
R811 B.n559 B.n558 10.6151
R812 B.n558 B.n557 10.6151
R813 B.n557 B.n4 10.6151
R814 B.n553 B.n4 10.6151
R815 B.n553 B.n552 10.6151
R816 B.n552 B.n551 10.6151
R817 B.n551 B.n6 10.6151
R818 B.n547 B.n6 10.6151
R819 B.n547 B.n546 10.6151
R820 B.n546 B.n545 10.6151
R821 B.n545 B.n8 10.6151
R822 B.n541 B.n8 10.6151
R823 B.n541 B.n540 10.6151
R824 B.n540 B.n539 10.6151
R825 B.n539 B.n10 10.6151
R826 B.n535 B.n10 10.6151
R827 B.n535 B.n534 10.6151
R828 B.n534 B.n533 10.6151
R829 B.n533 B.n12 10.6151
R830 B.n529 B.n12 10.6151
R831 B.n529 B.n528 10.6151
R832 B.n528 B.n527 10.6151
R833 B.n527 B.n14 10.6151
R834 B.n523 B.n14 10.6151
R835 B.n523 B.n522 10.6151
R836 B.n522 B.n521 10.6151
R837 B.n521 B.n16 10.6151
R838 B.n517 B.n16 10.6151
R839 B.n517 B.n516 10.6151
R840 B.n516 B.n515 10.6151
R841 B.n515 B.n18 10.6151
R842 B.n511 B.n18 10.6151
R843 B.n464 B.n36 6.5566
R844 B.n452 B.n451 6.5566
R845 B.n244 B.n116 6.5566
R846 B.n257 B.n256 6.5566
R847 B.n467 B.n36 4.05904
R848 B.n451 B.n450 4.05904
R849 B.n241 B.n116 4.05904
R850 B.n258 B.n257 4.05904
R851 B.n563 B.n0 2.81026
R852 B.n563 B.n1 2.81026
R853 VN.n4 VN.t0 223.238
R854 VN.n23 VN.t7 223.238
R855 VN.n17 VN.t4 200.136
R856 VN.n36 VN.t1 200.136
R857 VN.n10 VN.t2 165.558
R858 VN.n5 VN.t5 165.558
R859 VN.n1 VN.t6 165.558
R860 VN.n29 VN.t3 165.558
R861 VN.n24 VN.t9 165.558
R862 VN.n20 VN.t8 165.558
R863 VN.n35 VN.n19 161.3
R864 VN.n34 VN.n33 161.3
R865 VN.n32 VN.n31 161.3
R866 VN.n30 VN.n21 161.3
R867 VN.n29 VN.n28 161.3
R868 VN.n27 VN.n22 161.3
R869 VN.n26 VN.n25 161.3
R870 VN.n16 VN.n0 161.3
R871 VN.n15 VN.n14 161.3
R872 VN.n13 VN.n12 161.3
R873 VN.n11 VN.n2 161.3
R874 VN.n10 VN.n9 161.3
R875 VN.n8 VN.n3 161.3
R876 VN.n7 VN.n6 161.3
R877 VN.n37 VN.n36 80.6037
R878 VN.n18 VN.n17 80.6037
R879 VN.n6 VN.n3 56.4773
R880 VN.n12 VN.n11 56.4773
R881 VN.n25 VN.n22 56.4773
R882 VN.n31 VN.n30 56.4773
R883 VN.n17 VN.n16 50.8783
R884 VN.n36 VN.n35 50.8783
R885 VN VN.n37 42.6354
R886 VN.n5 VN.n4 33.6563
R887 VN.n24 VN.n23 33.6563
R888 VN.n26 VN.n23 28.104
R889 VN.n7 VN.n4 28.104
R890 VN.n10 VN.n3 24.3439
R891 VN.n11 VN.n10 24.3439
R892 VN.n16 VN.n15 24.3439
R893 VN.n30 VN.n29 24.3439
R894 VN.n29 VN.n22 24.3439
R895 VN.n35 VN.n34 24.3439
R896 VN.n6 VN.n5 23.3702
R897 VN.n12 VN.n1 23.3702
R898 VN.n25 VN.n24 23.3702
R899 VN.n31 VN.n20 23.3702
R900 VN.n15 VN.n1 0.974237
R901 VN.n34 VN.n20 0.974237
R902 VN.n37 VN.n19 0.285035
R903 VN.n18 VN.n0 0.285035
R904 VN.n33 VN.n19 0.189894
R905 VN.n33 VN.n32 0.189894
R906 VN.n32 VN.n21 0.189894
R907 VN.n28 VN.n21 0.189894
R908 VN.n28 VN.n27 0.189894
R909 VN.n27 VN.n26 0.189894
R910 VN.n8 VN.n7 0.189894
R911 VN.n9 VN.n8 0.189894
R912 VN.n9 VN.n2 0.189894
R913 VN.n13 VN.n2 0.189894
R914 VN.n14 VN.n13 0.189894
R915 VN.n14 VN.n0 0.189894
R916 VN VN.n18 0.146778
R917 VTAIL.n176 VTAIL.n140 756.745
R918 VTAIL.n38 VTAIL.n2 756.745
R919 VTAIL.n134 VTAIL.n98 756.745
R920 VTAIL.n88 VTAIL.n52 756.745
R921 VTAIL.n152 VTAIL.n151 585
R922 VTAIL.n157 VTAIL.n156 585
R923 VTAIL.n159 VTAIL.n158 585
R924 VTAIL.n148 VTAIL.n147 585
R925 VTAIL.n165 VTAIL.n164 585
R926 VTAIL.n167 VTAIL.n166 585
R927 VTAIL.n144 VTAIL.n143 585
R928 VTAIL.n174 VTAIL.n173 585
R929 VTAIL.n175 VTAIL.n142 585
R930 VTAIL.n177 VTAIL.n176 585
R931 VTAIL.n14 VTAIL.n13 585
R932 VTAIL.n19 VTAIL.n18 585
R933 VTAIL.n21 VTAIL.n20 585
R934 VTAIL.n10 VTAIL.n9 585
R935 VTAIL.n27 VTAIL.n26 585
R936 VTAIL.n29 VTAIL.n28 585
R937 VTAIL.n6 VTAIL.n5 585
R938 VTAIL.n36 VTAIL.n35 585
R939 VTAIL.n37 VTAIL.n4 585
R940 VTAIL.n39 VTAIL.n38 585
R941 VTAIL.n135 VTAIL.n134 585
R942 VTAIL.n133 VTAIL.n100 585
R943 VTAIL.n132 VTAIL.n131 585
R944 VTAIL.n103 VTAIL.n101 585
R945 VTAIL.n126 VTAIL.n125 585
R946 VTAIL.n124 VTAIL.n123 585
R947 VTAIL.n107 VTAIL.n106 585
R948 VTAIL.n118 VTAIL.n117 585
R949 VTAIL.n116 VTAIL.n115 585
R950 VTAIL.n111 VTAIL.n110 585
R951 VTAIL.n89 VTAIL.n88 585
R952 VTAIL.n87 VTAIL.n54 585
R953 VTAIL.n86 VTAIL.n85 585
R954 VTAIL.n57 VTAIL.n55 585
R955 VTAIL.n80 VTAIL.n79 585
R956 VTAIL.n78 VTAIL.n77 585
R957 VTAIL.n61 VTAIL.n60 585
R958 VTAIL.n72 VTAIL.n71 585
R959 VTAIL.n70 VTAIL.n69 585
R960 VTAIL.n65 VTAIL.n64 585
R961 VTAIL.n153 VTAIL.t16 329.043
R962 VTAIL.n15 VTAIL.t6 329.043
R963 VTAIL.n112 VTAIL.t1 329.043
R964 VTAIL.n66 VTAIL.t11 329.043
R965 VTAIL.n157 VTAIL.n151 171.744
R966 VTAIL.n158 VTAIL.n157 171.744
R967 VTAIL.n158 VTAIL.n147 171.744
R968 VTAIL.n165 VTAIL.n147 171.744
R969 VTAIL.n166 VTAIL.n165 171.744
R970 VTAIL.n166 VTAIL.n143 171.744
R971 VTAIL.n174 VTAIL.n143 171.744
R972 VTAIL.n175 VTAIL.n174 171.744
R973 VTAIL.n176 VTAIL.n175 171.744
R974 VTAIL.n19 VTAIL.n13 171.744
R975 VTAIL.n20 VTAIL.n19 171.744
R976 VTAIL.n20 VTAIL.n9 171.744
R977 VTAIL.n27 VTAIL.n9 171.744
R978 VTAIL.n28 VTAIL.n27 171.744
R979 VTAIL.n28 VTAIL.n5 171.744
R980 VTAIL.n36 VTAIL.n5 171.744
R981 VTAIL.n37 VTAIL.n36 171.744
R982 VTAIL.n38 VTAIL.n37 171.744
R983 VTAIL.n134 VTAIL.n133 171.744
R984 VTAIL.n133 VTAIL.n132 171.744
R985 VTAIL.n132 VTAIL.n101 171.744
R986 VTAIL.n125 VTAIL.n101 171.744
R987 VTAIL.n125 VTAIL.n124 171.744
R988 VTAIL.n124 VTAIL.n106 171.744
R989 VTAIL.n117 VTAIL.n106 171.744
R990 VTAIL.n117 VTAIL.n116 171.744
R991 VTAIL.n116 VTAIL.n110 171.744
R992 VTAIL.n88 VTAIL.n87 171.744
R993 VTAIL.n87 VTAIL.n86 171.744
R994 VTAIL.n86 VTAIL.n55 171.744
R995 VTAIL.n79 VTAIL.n55 171.744
R996 VTAIL.n79 VTAIL.n78 171.744
R997 VTAIL.n78 VTAIL.n60 171.744
R998 VTAIL.n71 VTAIL.n60 171.744
R999 VTAIL.n71 VTAIL.n70 171.744
R1000 VTAIL.n70 VTAIL.n64 171.744
R1001 VTAIL.t16 VTAIL.n151 85.8723
R1002 VTAIL.t6 VTAIL.n13 85.8723
R1003 VTAIL.t1 VTAIL.n110 85.8723
R1004 VTAIL.t11 VTAIL.n64 85.8723
R1005 VTAIL.n97 VTAIL.n96 67.6198
R1006 VTAIL.n95 VTAIL.n94 67.6198
R1007 VTAIL.n51 VTAIL.n50 67.6198
R1008 VTAIL.n49 VTAIL.n48 67.6198
R1009 VTAIL.n183 VTAIL.n182 67.6197
R1010 VTAIL.n1 VTAIL.n0 67.6197
R1011 VTAIL.n45 VTAIL.n44 67.6197
R1012 VTAIL.n47 VTAIL.n46 67.6197
R1013 VTAIL.n181 VTAIL.n180 34.1247
R1014 VTAIL.n43 VTAIL.n42 34.1247
R1015 VTAIL.n139 VTAIL.n138 34.1247
R1016 VTAIL.n93 VTAIL.n92 34.1247
R1017 VTAIL.n49 VTAIL.n47 21.7289
R1018 VTAIL.n181 VTAIL.n139 20.4531
R1019 VTAIL.n177 VTAIL.n142 13.1884
R1020 VTAIL.n39 VTAIL.n4 13.1884
R1021 VTAIL.n135 VTAIL.n100 13.1884
R1022 VTAIL.n89 VTAIL.n54 13.1884
R1023 VTAIL.n173 VTAIL.n172 12.8005
R1024 VTAIL.n178 VTAIL.n140 12.8005
R1025 VTAIL.n35 VTAIL.n34 12.8005
R1026 VTAIL.n40 VTAIL.n2 12.8005
R1027 VTAIL.n136 VTAIL.n98 12.8005
R1028 VTAIL.n131 VTAIL.n102 12.8005
R1029 VTAIL.n90 VTAIL.n52 12.8005
R1030 VTAIL.n85 VTAIL.n56 12.8005
R1031 VTAIL.n171 VTAIL.n144 12.0247
R1032 VTAIL.n33 VTAIL.n6 12.0247
R1033 VTAIL.n130 VTAIL.n103 12.0247
R1034 VTAIL.n84 VTAIL.n57 12.0247
R1035 VTAIL.n168 VTAIL.n167 11.249
R1036 VTAIL.n30 VTAIL.n29 11.249
R1037 VTAIL.n127 VTAIL.n126 11.249
R1038 VTAIL.n81 VTAIL.n80 11.249
R1039 VTAIL.n153 VTAIL.n152 10.7238
R1040 VTAIL.n15 VTAIL.n14 10.7238
R1041 VTAIL.n112 VTAIL.n111 10.7238
R1042 VTAIL.n66 VTAIL.n65 10.7238
R1043 VTAIL.n164 VTAIL.n146 10.4732
R1044 VTAIL.n26 VTAIL.n8 10.4732
R1045 VTAIL.n123 VTAIL.n105 10.4732
R1046 VTAIL.n77 VTAIL.n59 10.4732
R1047 VTAIL.n163 VTAIL.n148 9.69747
R1048 VTAIL.n25 VTAIL.n10 9.69747
R1049 VTAIL.n122 VTAIL.n107 9.69747
R1050 VTAIL.n76 VTAIL.n61 9.69747
R1051 VTAIL.n180 VTAIL.n179 9.45567
R1052 VTAIL.n42 VTAIL.n41 9.45567
R1053 VTAIL.n138 VTAIL.n137 9.45567
R1054 VTAIL.n92 VTAIL.n91 9.45567
R1055 VTAIL.n179 VTAIL.n178 9.3005
R1056 VTAIL.n155 VTAIL.n154 9.3005
R1057 VTAIL.n150 VTAIL.n149 9.3005
R1058 VTAIL.n161 VTAIL.n160 9.3005
R1059 VTAIL.n163 VTAIL.n162 9.3005
R1060 VTAIL.n146 VTAIL.n145 9.3005
R1061 VTAIL.n169 VTAIL.n168 9.3005
R1062 VTAIL.n171 VTAIL.n170 9.3005
R1063 VTAIL.n172 VTAIL.n141 9.3005
R1064 VTAIL.n41 VTAIL.n40 9.3005
R1065 VTAIL.n17 VTAIL.n16 9.3005
R1066 VTAIL.n12 VTAIL.n11 9.3005
R1067 VTAIL.n23 VTAIL.n22 9.3005
R1068 VTAIL.n25 VTAIL.n24 9.3005
R1069 VTAIL.n8 VTAIL.n7 9.3005
R1070 VTAIL.n31 VTAIL.n30 9.3005
R1071 VTAIL.n33 VTAIL.n32 9.3005
R1072 VTAIL.n34 VTAIL.n3 9.3005
R1073 VTAIL.n114 VTAIL.n113 9.3005
R1074 VTAIL.n109 VTAIL.n108 9.3005
R1075 VTAIL.n120 VTAIL.n119 9.3005
R1076 VTAIL.n122 VTAIL.n121 9.3005
R1077 VTAIL.n105 VTAIL.n104 9.3005
R1078 VTAIL.n128 VTAIL.n127 9.3005
R1079 VTAIL.n130 VTAIL.n129 9.3005
R1080 VTAIL.n102 VTAIL.n99 9.3005
R1081 VTAIL.n137 VTAIL.n136 9.3005
R1082 VTAIL.n68 VTAIL.n67 9.3005
R1083 VTAIL.n63 VTAIL.n62 9.3005
R1084 VTAIL.n74 VTAIL.n73 9.3005
R1085 VTAIL.n76 VTAIL.n75 9.3005
R1086 VTAIL.n59 VTAIL.n58 9.3005
R1087 VTAIL.n82 VTAIL.n81 9.3005
R1088 VTAIL.n84 VTAIL.n83 9.3005
R1089 VTAIL.n56 VTAIL.n53 9.3005
R1090 VTAIL.n91 VTAIL.n90 9.3005
R1091 VTAIL.n160 VTAIL.n159 8.92171
R1092 VTAIL.n22 VTAIL.n21 8.92171
R1093 VTAIL.n119 VTAIL.n118 8.92171
R1094 VTAIL.n73 VTAIL.n72 8.92171
R1095 VTAIL.n156 VTAIL.n150 8.14595
R1096 VTAIL.n18 VTAIL.n12 8.14595
R1097 VTAIL.n115 VTAIL.n109 8.14595
R1098 VTAIL.n69 VTAIL.n63 8.14595
R1099 VTAIL.n155 VTAIL.n152 7.3702
R1100 VTAIL.n17 VTAIL.n14 7.3702
R1101 VTAIL.n114 VTAIL.n111 7.3702
R1102 VTAIL.n68 VTAIL.n65 7.3702
R1103 VTAIL.n156 VTAIL.n155 5.81868
R1104 VTAIL.n18 VTAIL.n17 5.81868
R1105 VTAIL.n115 VTAIL.n114 5.81868
R1106 VTAIL.n69 VTAIL.n68 5.81868
R1107 VTAIL.n159 VTAIL.n150 5.04292
R1108 VTAIL.n21 VTAIL.n12 5.04292
R1109 VTAIL.n118 VTAIL.n109 5.04292
R1110 VTAIL.n72 VTAIL.n63 5.04292
R1111 VTAIL.n160 VTAIL.n148 4.26717
R1112 VTAIL.n22 VTAIL.n10 4.26717
R1113 VTAIL.n119 VTAIL.n107 4.26717
R1114 VTAIL.n73 VTAIL.n61 4.26717
R1115 VTAIL.n182 VTAIL.t15 4.11506
R1116 VTAIL.n182 VTAIL.t18 4.11506
R1117 VTAIL.n0 VTAIL.t13 4.11506
R1118 VTAIL.n0 VTAIL.t17 4.11506
R1119 VTAIL.n44 VTAIL.t5 4.11506
R1120 VTAIL.n44 VTAIL.t8 4.11506
R1121 VTAIL.n46 VTAIL.t9 4.11506
R1122 VTAIL.n46 VTAIL.t7 4.11506
R1123 VTAIL.n96 VTAIL.t4 4.11506
R1124 VTAIL.n96 VTAIL.t3 4.11506
R1125 VTAIL.n94 VTAIL.t0 4.11506
R1126 VTAIL.n94 VTAIL.t2 4.11506
R1127 VTAIL.n50 VTAIL.t10 4.11506
R1128 VTAIL.n50 VTAIL.t19 4.11506
R1129 VTAIL.n48 VTAIL.t14 4.11506
R1130 VTAIL.n48 VTAIL.t12 4.11506
R1131 VTAIL.n164 VTAIL.n163 3.49141
R1132 VTAIL.n26 VTAIL.n25 3.49141
R1133 VTAIL.n123 VTAIL.n122 3.49141
R1134 VTAIL.n77 VTAIL.n76 3.49141
R1135 VTAIL.n167 VTAIL.n146 2.71565
R1136 VTAIL.n29 VTAIL.n8 2.71565
R1137 VTAIL.n126 VTAIL.n105 2.71565
R1138 VTAIL.n80 VTAIL.n59 2.71565
R1139 VTAIL.n154 VTAIL.n153 2.4129
R1140 VTAIL.n16 VTAIL.n15 2.4129
R1141 VTAIL.n113 VTAIL.n112 2.4129
R1142 VTAIL.n67 VTAIL.n66 2.4129
R1143 VTAIL.n168 VTAIL.n144 1.93989
R1144 VTAIL.n30 VTAIL.n6 1.93989
R1145 VTAIL.n127 VTAIL.n103 1.93989
R1146 VTAIL.n81 VTAIL.n57 1.93989
R1147 VTAIL.n51 VTAIL.n49 1.27636
R1148 VTAIL.n93 VTAIL.n51 1.27636
R1149 VTAIL.n97 VTAIL.n95 1.27636
R1150 VTAIL.n139 VTAIL.n97 1.27636
R1151 VTAIL.n47 VTAIL.n45 1.27636
R1152 VTAIL.n45 VTAIL.n43 1.27636
R1153 VTAIL.n183 VTAIL.n181 1.27636
R1154 VTAIL.n173 VTAIL.n171 1.16414
R1155 VTAIL.n180 VTAIL.n140 1.16414
R1156 VTAIL.n35 VTAIL.n33 1.16414
R1157 VTAIL.n42 VTAIL.n2 1.16414
R1158 VTAIL.n138 VTAIL.n98 1.16414
R1159 VTAIL.n131 VTAIL.n130 1.16414
R1160 VTAIL.n92 VTAIL.n52 1.16414
R1161 VTAIL.n85 VTAIL.n84 1.16414
R1162 VTAIL.n95 VTAIL.n93 1.10826
R1163 VTAIL.n43 VTAIL.n1 1.10826
R1164 VTAIL VTAIL.n1 1.01559
R1165 VTAIL.n172 VTAIL.n142 0.388379
R1166 VTAIL.n178 VTAIL.n177 0.388379
R1167 VTAIL.n34 VTAIL.n4 0.388379
R1168 VTAIL.n40 VTAIL.n39 0.388379
R1169 VTAIL.n136 VTAIL.n135 0.388379
R1170 VTAIL.n102 VTAIL.n100 0.388379
R1171 VTAIL.n90 VTAIL.n89 0.388379
R1172 VTAIL.n56 VTAIL.n54 0.388379
R1173 VTAIL VTAIL.n183 0.261276
R1174 VTAIL.n154 VTAIL.n149 0.155672
R1175 VTAIL.n161 VTAIL.n149 0.155672
R1176 VTAIL.n162 VTAIL.n161 0.155672
R1177 VTAIL.n162 VTAIL.n145 0.155672
R1178 VTAIL.n169 VTAIL.n145 0.155672
R1179 VTAIL.n170 VTAIL.n169 0.155672
R1180 VTAIL.n170 VTAIL.n141 0.155672
R1181 VTAIL.n179 VTAIL.n141 0.155672
R1182 VTAIL.n16 VTAIL.n11 0.155672
R1183 VTAIL.n23 VTAIL.n11 0.155672
R1184 VTAIL.n24 VTAIL.n23 0.155672
R1185 VTAIL.n24 VTAIL.n7 0.155672
R1186 VTAIL.n31 VTAIL.n7 0.155672
R1187 VTAIL.n32 VTAIL.n31 0.155672
R1188 VTAIL.n32 VTAIL.n3 0.155672
R1189 VTAIL.n41 VTAIL.n3 0.155672
R1190 VTAIL.n137 VTAIL.n99 0.155672
R1191 VTAIL.n129 VTAIL.n99 0.155672
R1192 VTAIL.n129 VTAIL.n128 0.155672
R1193 VTAIL.n128 VTAIL.n104 0.155672
R1194 VTAIL.n121 VTAIL.n104 0.155672
R1195 VTAIL.n121 VTAIL.n120 0.155672
R1196 VTAIL.n120 VTAIL.n108 0.155672
R1197 VTAIL.n113 VTAIL.n108 0.155672
R1198 VTAIL.n91 VTAIL.n53 0.155672
R1199 VTAIL.n83 VTAIL.n53 0.155672
R1200 VTAIL.n83 VTAIL.n82 0.155672
R1201 VTAIL.n82 VTAIL.n58 0.155672
R1202 VTAIL.n75 VTAIL.n58 0.155672
R1203 VTAIL.n75 VTAIL.n74 0.155672
R1204 VTAIL.n74 VTAIL.n62 0.155672
R1205 VTAIL.n67 VTAIL.n62 0.155672
R1206 VDD2.n81 VDD2.n45 756.745
R1207 VDD2.n36 VDD2.n0 756.745
R1208 VDD2.n82 VDD2.n81 585
R1209 VDD2.n80 VDD2.n47 585
R1210 VDD2.n79 VDD2.n78 585
R1211 VDD2.n50 VDD2.n48 585
R1212 VDD2.n73 VDD2.n72 585
R1213 VDD2.n71 VDD2.n70 585
R1214 VDD2.n54 VDD2.n53 585
R1215 VDD2.n65 VDD2.n64 585
R1216 VDD2.n63 VDD2.n62 585
R1217 VDD2.n58 VDD2.n57 585
R1218 VDD2.n12 VDD2.n11 585
R1219 VDD2.n17 VDD2.n16 585
R1220 VDD2.n19 VDD2.n18 585
R1221 VDD2.n8 VDD2.n7 585
R1222 VDD2.n25 VDD2.n24 585
R1223 VDD2.n27 VDD2.n26 585
R1224 VDD2.n4 VDD2.n3 585
R1225 VDD2.n34 VDD2.n33 585
R1226 VDD2.n35 VDD2.n2 585
R1227 VDD2.n37 VDD2.n36 585
R1228 VDD2.n59 VDD2.t8 329.043
R1229 VDD2.n13 VDD2.t9 329.043
R1230 VDD2.n81 VDD2.n80 171.744
R1231 VDD2.n80 VDD2.n79 171.744
R1232 VDD2.n79 VDD2.n48 171.744
R1233 VDD2.n72 VDD2.n48 171.744
R1234 VDD2.n72 VDD2.n71 171.744
R1235 VDD2.n71 VDD2.n53 171.744
R1236 VDD2.n64 VDD2.n53 171.744
R1237 VDD2.n64 VDD2.n63 171.744
R1238 VDD2.n63 VDD2.n57 171.744
R1239 VDD2.n17 VDD2.n11 171.744
R1240 VDD2.n18 VDD2.n17 171.744
R1241 VDD2.n18 VDD2.n7 171.744
R1242 VDD2.n25 VDD2.n7 171.744
R1243 VDD2.n26 VDD2.n25 171.744
R1244 VDD2.n26 VDD2.n3 171.744
R1245 VDD2.n34 VDD2.n3 171.744
R1246 VDD2.n35 VDD2.n34 171.744
R1247 VDD2.n36 VDD2.n35 171.744
R1248 VDD2.t8 VDD2.n57 85.8723
R1249 VDD2.t9 VDD2.n11 85.8723
R1250 VDD2.n44 VDD2.n43 85.2
R1251 VDD2 VDD2.n89 85.1972
R1252 VDD2.n88 VDD2.n87 84.2986
R1253 VDD2.n42 VDD2.n41 84.2985
R1254 VDD2.n42 VDD2.n40 52.0794
R1255 VDD2.n86 VDD2.n85 50.8035
R1256 VDD2.n86 VDD2.n44 36.586
R1257 VDD2.n82 VDD2.n47 13.1884
R1258 VDD2.n37 VDD2.n2 13.1884
R1259 VDD2.n83 VDD2.n45 12.8005
R1260 VDD2.n78 VDD2.n49 12.8005
R1261 VDD2.n33 VDD2.n32 12.8005
R1262 VDD2.n38 VDD2.n0 12.8005
R1263 VDD2.n77 VDD2.n50 12.0247
R1264 VDD2.n31 VDD2.n4 12.0247
R1265 VDD2.n74 VDD2.n73 11.249
R1266 VDD2.n28 VDD2.n27 11.249
R1267 VDD2.n59 VDD2.n58 10.7238
R1268 VDD2.n13 VDD2.n12 10.7238
R1269 VDD2.n70 VDD2.n52 10.4732
R1270 VDD2.n24 VDD2.n6 10.4732
R1271 VDD2.n69 VDD2.n54 9.69747
R1272 VDD2.n23 VDD2.n8 9.69747
R1273 VDD2.n85 VDD2.n84 9.45567
R1274 VDD2.n40 VDD2.n39 9.45567
R1275 VDD2.n61 VDD2.n60 9.3005
R1276 VDD2.n56 VDD2.n55 9.3005
R1277 VDD2.n67 VDD2.n66 9.3005
R1278 VDD2.n69 VDD2.n68 9.3005
R1279 VDD2.n52 VDD2.n51 9.3005
R1280 VDD2.n75 VDD2.n74 9.3005
R1281 VDD2.n77 VDD2.n76 9.3005
R1282 VDD2.n49 VDD2.n46 9.3005
R1283 VDD2.n84 VDD2.n83 9.3005
R1284 VDD2.n39 VDD2.n38 9.3005
R1285 VDD2.n15 VDD2.n14 9.3005
R1286 VDD2.n10 VDD2.n9 9.3005
R1287 VDD2.n21 VDD2.n20 9.3005
R1288 VDD2.n23 VDD2.n22 9.3005
R1289 VDD2.n6 VDD2.n5 9.3005
R1290 VDD2.n29 VDD2.n28 9.3005
R1291 VDD2.n31 VDD2.n30 9.3005
R1292 VDD2.n32 VDD2.n1 9.3005
R1293 VDD2.n66 VDD2.n65 8.92171
R1294 VDD2.n20 VDD2.n19 8.92171
R1295 VDD2.n62 VDD2.n56 8.14595
R1296 VDD2.n16 VDD2.n10 8.14595
R1297 VDD2.n61 VDD2.n58 7.3702
R1298 VDD2.n15 VDD2.n12 7.3702
R1299 VDD2.n62 VDD2.n61 5.81868
R1300 VDD2.n16 VDD2.n15 5.81868
R1301 VDD2.n65 VDD2.n56 5.04292
R1302 VDD2.n19 VDD2.n10 5.04292
R1303 VDD2.n66 VDD2.n54 4.26717
R1304 VDD2.n20 VDD2.n8 4.26717
R1305 VDD2.n89 VDD2.t0 4.11506
R1306 VDD2.n89 VDD2.t2 4.11506
R1307 VDD2.n87 VDD2.t1 4.11506
R1308 VDD2.n87 VDD2.t6 4.11506
R1309 VDD2.n43 VDD2.t3 4.11506
R1310 VDD2.n43 VDD2.t5 4.11506
R1311 VDD2.n41 VDD2.t4 4.11506
R1312 VDD2.n41 VDD2.t7 4.11506
R1313 VDD2.n70 VDD2.n69 3.49141
R1314 VDD2.n24 VDD2.n23 3.49141
R1315 VDD2.n73 VDD2.n52 2.71565
R1316 VDD2.n27 VDD2.n6 2.71565
R1317 VDD2.n60 VDD2.n59 2.4129
R1318 VDD2.n14 VDD2.n13 2.4129
R1319 VDD2.n74 VDD2.n50 1.93989
R1320 VDD2.n28 VDD2.n4 1.93989
R1321 VDD2.n88 VDD2.n86 1.27636
R1322 VDD2.n85 VDD2.n45 1.16414
R1323 VDD2.n78 VDD2.n77 1.16414
R1324 VDD2.n33 VDD2.n31 1.16414
R1325 VDD2.n40 VDD2.n0 1.16414
R1326 VDD2.n83 VDD2.n82 0.388379
R1327 VDD2.n49 VDD2.n47 0.388379
R1328 VDD2.n32 VDD2.n2 0.388379
R1329 VDD2.n38 VDD2.n37 0.388379
R1330 VDD2 VDD2.n88 0.377655
R1331 VDD2.n44 VDD2.n42 0.26412
R1332 VDD2.n84 VDD2.n46 0.155672
R1333 VDD2.n76 VDD2.n46 0.155672
R1334 VDD2.n76 VDD2.n75 0.155672
R1335 VDD2.n75 VDD2.n51 0.155672
R1336 VDD2.n68 VDD2.n51 0.155672
R1337 VDD2.n68 VDD2.n67 0.155672
R1338 VDD2.n67 VDD2.n55 0.155672
R1339 VDD2.n60 VDD2.n55 0.155672
R1340 VDD2.n14 VDD2.n9 0.155672
R1341 VDD2.n21 VDD2.n9 0.155672
R1342 VDD2.n22 VDD2.n21 0.155672
R1343 VDD2.n22 VDD2.n5 0.155672
R1344 VDD2.n29 VDD2.n5 0.155672
R1345 VDD2.n30 VDD2.n29 0.155672
R1346 VDD2.n30 VDD2.n1 0.155672
R1347 VDD2.n39 VDD2.n1 0.155672
R1348 VP.n10 VP.t9 223.238
R1349 VP.n5 VP.t5 200.136
R1350 VP.n41 VP.t4 200.136
R1351 VP.n23 VP.t2 200.136
R1352 VP.n34 VP.t7 165.558
R1353 VP.n29 VP.t3 165.558
R1354 VP.n1 VP.t8 165.558
R1355 VP.n16 VP.t6 165.558
R1356 VP.n7 VP.t0 165.558
R1357 VP.n11 VP.t1 165.558
R1358 VP.n13 VP.n12 161.3
R1359 VP.n14 VP.n9 161.3
R1360 VP.n16 VP.n15 161.3
R1361 VP.n17 VP.n8 161.3
R1362 VP.n19 VP.n18 161.3
R1363 VP.n21 VP.n20 161.3
R1364 VP.n22 VP.n6 161.3
R1365 VP.n40 VP.n0 161.3
R1366 VP.n39 VP.n38 161.3
R1367 VP.n37 VP.n36 161.3
R1368 VP.n35 VP.n2 161.3
R1369 VP.n34 VP.n33 161.3
R1370 VP.n32 VP.n3 161.3
R1371 VP.n31 VP.n30 161.3
R1372 VP.n28 VP.n4 161.3
R1373 VP.n27 VP.n26 161.3
R1374 VP.n24 VP.n23 80.6037
R1375 VP.n42 VP.n41 80.6037
R1376 VP.n25 VP.n5 80.6037
R1377 VP.n30 VP.n3 56.4773
R1378 VP.n36 VP.n35 56.4773
R1379 VP.n18 VP.n17 56.4773
R1380 VP.n12 VP.n9 56.4773
R1381 VP.n27 VP.n5 50.8783
R1382 VP.n41 VP.n40 50.8783
R1383 VP.n23 VP.n22 50.8783
R1384 VP.n25 VP.n24 42.3499
R1385 VP.n11 VP.n10 33.6563
R1386 VP.n13 VP.n10 28.104
R1387 VP.n28 VP.n27 24.3439
R1388 VP.n34 VP.n3 24.3439
R1389 VP.n35 VP.n34 24.3439
R1390 VP.n40 VP.n39 24.3439
R1391 VP.n22 VP.n21 24.3439
R1392 VP.n16 VP.n9 24.3439
R1393 VP.n17 VP.n16 24.3439
R1394 VP.n30 VP.n29 23.3702
R1395 VP.n36 VP.n1 23.3702
R1396 VP.n18 VP.n7 23.3702
R1397 VP.n12 VP.n11 23.3702
R1398 VP.n29 VP.n28 0.974237
R1399 VP.n39 VP.n1 0.974237
R1400 VP.n21 VP.n7 0.974237
R1401 VP.n24 VP.n6 0.285035
R1402 VP.n26 VP.n25 0.285035
R1403 VP.n42 VP.n0 0.285035
R1404 VP.n14 VP.n13 0.189894
R1405 VP.n15 VP.n14 0.189894
R1406 VP.n15 VP.n8 0.189894
R1407 VP.n19 VP.n8 0.189894
R1408 VP.n20 VP.n19 0.189894
R1409 VP.n20 VP.n6 0.189894
R1410 VP.n26 VP.n4 0.189894
R1411 VP.n31 VP.n4 0.189894
R1412 VP.n32 VP.n31 0.189894
R1413 VP.n33 VP.n32 0.189894
R1414 VP.n33 VP.n2 0.189894
R1415 VP.n37 VP.n2 0.189894
R1416 VP.n38 VP.n37 0.189894
R1417 VP.n38 VP.n0 0.189894
R1418 VP VP.n42 0.146778
R1419 VDD1.n36 VDD1.n0 756.745
R1420 VDD1.n79 VDD1.n43 756.745
R1421 VDD1.n37 VDD1.n36 585
R1422 VDD1.n35 VDD1.n2 585
R1423 VDD1.n34 VDD1.n33 585
R1424 VDD1.n5 VDD1.n3 585
R1425 VDD1.n28 VDD1.n27 585
R1426 VDD1.n26 VDD1.n25 585
R1427 VDD1.n9 VDD1.n8 585
R1428 VDD1.n20 VDD1.n19 585
R1429 VDD1.n18 VDD1.n17 585
R1430 VDD1.n13 VDD1.n12 585
R1431 VDD1.n55 VDD1.n54 585
R1432 VDD1.n60 VDD1.n59 585
R1433 VDD1.n62 VDD1.n61 585
R1434 VDD1.n51 VDD1.n50 585
R1435 VDD1.n68 VDD1.n67 585
R1436 VDD1.n70 VDD1.n69 585
R1437 VDD1.n47 VDD1.n46 585
R1438 VDD1.n77 VDD1.n76 585
R1439 VDD1.n78 VDD1.n45 585
R1440 VDD1.n80 VDD1.n79 585
R1441 VDD1.n14 VDD1.t0 329.043
R1442 VDD1.n56 VDD1.t4 329.043
R1443 VDD1.n36 VDD1.n35 171.744
R1444 VDD1.n35 VDD1.n34 171.744
R1445 VDD1.n34 VDD1.n3 171.744
R1446 VDD1.n27 VDD1.n3 171.744
R1447 VDD1.n27 VDD1.n26 171.744
R1448 VDD1.n26 VDD1.n8 171.744
R1449 VDD1.n19 VDD1.n8 171.744
R1450 VDD1.n19 VDD1.n18 171.744
R1451 VDD1.n18 VDD1.n12 171.744
R1452 VDD1.n60 VDD1.n54 171.744
R1453 VDD1.n61 VDD1.n60 171.744
R1454 VDD1.n61 VDD1.n50 171.744
R1455 VDD1.n68 VDD1.n50 171.744
R1456 VDD1.n69 VDD1.n68 171.744
R1457 VDD1.n69 VDD1.n46 171.744
R1458 VDD1.n77 VDD1.n46 171.744
R1459 VDD1.n78 VDD1.n77 171.744
R1460 VDD1.n79 VDD1.n78 171.744
R1461 VDD1.t0 VDD1.n12 85.8723
R1462 VDD1.t4 VDD1.n54 85.8723
R1463 VDD1.n87 VDD1.n86 85.2
R1464 VDD1.n42 VDD1.n41 84.2986
R1465 VDD1.n89 VDD1.n88 84.2985
R1466 VDD1.n85 VDD1.n84 84.2985
R1467 VDD1.n42 VDD1.n40 52.0794
R1468 VDD1.n85 VDD1.n83 52.0794
R1469 VDD1.n89 VDD1.n87 37.8069
R1470 VDD1.n37 VDD1.n2 13.1884
R1471 VDD1.n80 VDD1.n45 13.1884
R1472 VDD1.n38 VDD1.n0 12.8005
R1473 VDD1.n33 VDD1.n4 12.8005
R1474 VDD1.n76 VDD1.n75 12.8005
R1475 VDD1.n81 VDD1.n43 12.8005
R1476 VDD1.n32 VDD1.n5 12.0247
R1477 VDD1.n74 VDD1.n47 12.0247
R1478 VDD1.n29 VDD1.n28 11.249
R1479 VDD1.n71 VDD1.n70 11.249
R1480 VDD1.n14 VDD1.n13 10.7238
R1481 VDD1.n56 VDD1.n55 10.7238
R1482 VDD1.n25 VDD1.n7 10.4732
R1483 VDD1.n67 VDD1.n49 10.4732
R1484 VDD1.n24 VDD1.n9 9.69747
R1485 VDD1.n66 VDD1.n51 9.69747
R1486 VDD1.n40 VDD1.n39 9.45567
R1487 VDD1.n83 VDD1.n82 9.45567
R1488 VDD1.n16 VDD1.n15 9.3005
R1489 VDD1.n11 VDD1.n10 9.3005
R1490 VDD1.n22 VDD1.n21 9.3005
R1491 VDD1.n24 VDD1.n23 9.3005
R1492 VDD1.n7 VDD1.n6 9.3005
R1493 VDD1.n30 VDD1.n29 9.3005
R1494 VDD1.n32 VDD1.n31 9.3005
R1495 VDD1.n4 VDD1.n1 9.3005
R1496 VDD1.n39 VDD1.n38 9.3005
R1497 VDD1.n82 VDD1.n81 9.3005
R1498 VDD1.n58 VDD1.n57 9.3005
R1499 VDD1.n53 VDD1.n52 9.3005
R1500 VDD1.n64 VDD1.n63 9.3005
R1501 VDD1.n66 VDD1.n65 9.3005
R1502 VDD1.n49 VDD1.n48 9.3005
R1503 VDD1.n72 VDD1.n71 9.3005
R1504 VDD1.n74 VDD1.n73 9.3005
R1505 VDD1.n75 VDD1.n44 9.3005
R1506 VDD1.n21 VDD1.n20 8.92171
R1507 VDD1.n63 VDD1.n62 8.92171
R1508 VDD1.n17 VDD1.n11 8.14595
R1509 VDD1.n59 VDD1.n53 8.14595
R1510 VDD1.n16 VDD1.n13 7.3702
R1511 VDD1.n58 VDD1.n55 7.3702
R1512 VDD1.n17 VDD1.n16 5.81868
R1513 VDD1.n59 VDD1.n58 5.81868
R1514 VDD1.n20 VDD1.n11 5.04292
R1515 VDD1.n62 VDD1.n53 5.04292
R1516 VDD1.n21 VDD1.n9 4.26717
R1517 VDD1.n63 VDD1.n51 4.26717
R1518 VDD1.n88 VDD1.t9 4.11506
R1519 VDD1.n88 VDD1.t7 4.11506
R1520 VDD1.n41 VDD1.t8 4.11506
R1521 VDD1.n41 VDD1.t3 4.11506
R1522 VDD1.n86 VDD1.t1 4.11506
R1523 VDD1.n86 VDD1.t5 4.11506
R1524 VDD1.n84 VDD1.t6 4.11506
R1525 VDD1.n84 VDD1.t2 4.11506
R1526 VDD1.n25 VDD1.n24 3.49141
R1527 VDD1.n67 VDD1.n66 3.49141
R1528 VDD1.n28 VDD1.n7 2.71565
R1529 VDD1.n70 VDD1.n49 2.71565
R1530 VDD1.n15 VDD1.n14 2.4129
R1531 VDD1.n57 VDD1.n56 2.4129
R1532 VDD1.n29 VDD1.n5 1.93989
R1533 VDD1.n71 VDD1.n47 1.93989
R1534 VDD1.n40 VDD1.n0 1.16414
R1535 VDD1.n33 VDD1.n32 1.16414
R1536 VDD1.n76 VDD1.n74 1.16414
R1537 VDD1.n83 VDD1.n43 1.16414
R1538 VDD1 VDD1.n89 0.899207
R1539 VDD1.n38 VDD1.n37 0.388379
R1540 VDD1.n4 VDD1.n2 0.388379
R1541 VDD1.n75 VDD1.n45 0.388379
R1542 VDD1.n81 VDD1.n80 0.388379
R1543 VDD1 VDD1.n42 0.377655
R1544 VDD1.n87 VDD1.n85 0.26412
R1545 VDD1.n39 VDD1.n1 0.155672
R1546 VDD1.n31 VDD1.n1 0.155672
R1547 VDD1.n31 VDD1.n30 0.155672
R1548 VDD1.n30 VDD1.n6 0.155672
R1549 VDD1.n23 VDD1.n6 0.155672
R1550 VDD1.n23 VDD1.n22 0.155672
R1551 VDD1.n22 VDD1.n10 0.155672
R1552 VDD1.n15 VDD1.n10 0.155672
R1553 VDD1.n57 VDD1.n52 0.155672
R1554 VDD1.n64 VDD1.n52 0.155672
R1555 VDD1.n65 VDD1.n64 0.155672
R1556 VDD1.n65 VDD1.n48 0.155672
R1557 VDD1.n72 VDD1.n48 0.155672
R1558 VDD1.n73 VDD1.n72 0.155672
R1559 VDD1.n73 VDD1.n44 0.155672
R1560 VDD1.n82 VDD1.n44 0.155672
C0 VTAIL VDD1 8.775579f
C1 VTAIL w_n2746_n2548# 2.43681f
C2 VP VN 5.50263f
C3 w_n2746_n2548# VDD1 1.93649f
C4 VN B 0.863469f
C5 VDD2 VTAIL 8.816059f
C6 VDD2 VDD1 1.24808f
C7 VDD2 w_n2746_n2548# 2.00462f
C8 VP B 1.44913f
C9 VTAIL VN 5.88829f
C10 VDD1 VN 0.149849f
C11 w_n2746_n2548# VN 5.34904f
C12 VDD2 VN 5.69185f
C13 VTAIL VP 5.90265f
C14 VTAIL B 2.22646f
C15 VP VDD1 5.93698f
C16 w_n2746_n2548# VP 5.70208f
C17 VDD1 B 1.58891f
C18 w_n2746_n2548# B 6.95859f
C19 VDD2 VP 0.398088f
C20 VDD2 B 1.65046f
C21 VDD2 VSUBS 1.411783f
C22 VDD1 VSUBS 1.206487f
C23 VTAIL VSUBS 0.795743f
C24 VN VSUBS 5.27602f
C25 VP VSUBS 2.264711f
C26 B VSUBS 3.220737f
C27 w_n2746_n2548# VSUBS 86.8285f
C28 VDD1.n0 VSUBS 0.024068f
C29 VDD1.n1 VSUBS 0.023248f
C30 VDD1.n2 VSUBS 0.01286f
C31 VDD1.n3 VSUBS 0.029528f
C32 VDD1.n4 VSUBS 0.012493f
C33 VDD1.n5 VSUBS 0.013228f
C34 VDD1.n6 VSUBS 0.023248f
C35 VDD1.n7 VSUBS 0.012493f
C36 VDD1.n8 VSUBS 0.029528f
C37 VDD1.n9 VSUBS 0.013228f
C38 VDD1.n10 VSUBS 0.023248f
C39 VDD1.n11 VSUBS 0.012493f
C40 VDD1.n12 VSUBS 0.022146f
C41 VDD1.n13 VSUBS 0.022212f
C42 VDD1.t0 VSUBS 0.063405f
C43 VDD1.n14 VSUBS 0.140078f
C44 VDD1.n15 VSUBS 0.724444f
C45 VDD1.n16 VSUBS 0.012493f
C46 VDD1.n17 VSUBS 0.013228f
C47 VDD1.n18 VSUBS 0.029528f
C48 VDD1.n19 VSUBS 0.029528f
C49 VDD1.n20 VSUBS 0.013228f
C50 VDD1.n21 VSUBS 0.012493f
C51 VDD1.n22 VSUBS 0.023248f
C52 VDD1.n23 VSUBS 0.023248f
C53 VDD1.n24 VSUBS 0.012493f
C54 VDD1.n25 VSUBS 0.013228f
C55 VDD1.n26 VSUBS 0.029528f
C56 VDD1.n27 VSUBS 0.029528f
C57 VDD1.n28 VSUBS 0.013228f
C58 VDD1.n29 VSUBS 0.012493f
C59 VDD1.n30 VSUBS 0.023248f
C60 VDD1.n31 VSUBS 0.023248f
C61 VDD1.n32 VSUBS 0.012493f
C62 VDD1.n33 VSUBS 0.013228f
C63 VDD1.n34 VSUBS 0.029528f
C64 VDD1.n35 VSUBS 0.029528f
C65 VDD1.n36 VSUBS 0.066454f
C66 VDD1.n37 VSUBS 0.01286f
C67 VDD1.n38 VSUBS 0.012493f
C68 VDD1.n39 VSUBS 0.056914f
C69 VDD1.n40 VSUBS 0.052803f
C70 VDD1.t8 VSUBS 0.145136f
C71 VDD1.t3 VSUBS 0.145136f
C72 VDD1.n41 VSUBS 1.04777f
C73 VDD1.n42 VSUBS 0.654887f
C74 VDD1.n43 VSUBS 0.024068f
C75 VDD1.n44 VSUBS 0.023248f
C76 VDD1.n45 VSUBS 0.01286f
C77 VDD1.n46 VSUBS 0.029528f
C78 VDD1.n47 VSUBS 0.013228f
C79 VDD1.n48 VSUBS 0.023248f
C80 VDD1.n49 VSUBS 0.012493f
C81 VDD1.n50 VSUBS 0.029528f
C82 VDD1.n51 VSUBS 0.013228f
C83 VDD1.n52 VSUBS 0.023248f
C84 VDD1.n53 VSUBS 0.012493f
C85 VDD1.n54 VSUBS 0.022146f
C86 VDD1.n55 VSUBS 0.022212f
C87 VDD1.t4 VSUBS 0.063405f
C88 VDD1.n56 VSUBS 0.140078f
C89 VDD1.n57 VSUBS 0.724444f
C90 VDD1.n58 VSUBS 0.012493f
C91 VDD1.n59 VSUBS 0.013228f
C92 VDD1.n60 VSUBS 0.029528f
C93 VDD1.n61 VSUBS 0.029528f
C94 VDD1.n62 VSUBS 0.013228f
C95 VDD1.n63 VSUBS 0.012493f
C96 VDD1.n64 VSUBS 0.023248f
C97 VDD1.n65 VSUBS 0.023248f
C98 VDD1.n66 VSUBS 0.012493f
C99 VDD1.n67 VSUBS 0.013228f
C100 VDD1.n68 VSUBS 0.029528f
C101 VDD1.n69 VSUBS 0.029528f
C102 VDD1.n70 VSUBS 0.013228f
C103 VDD1.n71 VSUBS 0.012493f
C104 VDD1.n72 VSUBS 0.023248f
C105 VDD1.n73 VSUBS 0.023248f
C106 VDD1.n74 VSUBS 0.012493f
C107 VDD1.n75 VSUBS 0.012493f
C108 VDD1.n76 VSUBS 0.013228f
C109 VDD1.n77 VSUBS 0.029528f
C110 VDD1.n78 VSUBS 0.029528f
C111 VDD1.n79 VSUBS 0.066454f
C112 VDD1.n80 VSUBS 0.01286f
C113 VDD1.n81 VSUBS 0.012493f
C114 VDD1.n82 VSUBS 0.056914f
C115 VDD1.n83 VSUBS 0.052803f
C116 VDD1.t6 VSUBS 0.145136f
C117 VDD1.t2 VSUBS 0.145136f
C118 VDD1.n84 VSUBS 1.04777f
C119 VDD1.n85 VSUBS 0.648431f
C120 VDD1.t1 VSUBS 0.145136f
C121 VDD1.t5 VSUBS 0.145136f
C122 VDD1.n86 VSUBS 1.05375f
C123 VDD1.n87 VSUBS 2.04273f
C124 VDD1.t9 VSUBS 0.145136f
C125 VDD1.t7 VSUBS 0.145136f
C126 VDD1.n88 VSUBS 1.04777f
C127 VDD1.n89 VSUBS 2.29574f
C128 VP.n0 VSUBS 0.063441f
C129 VP.t8 VSUBS 1.1594f
C130 VP.n1 VSUBS 0.447461f
C131 VP.n2 VSUBS 0.047543f
C132 VP.t7 VSUBS 1.1594f
C133 VP.n3 VSUBS 0.068373f
C134 VP.n4 VSUBS 0.047543f
C135 VP.t3 VSUBS 1.1594f
C136 VP.t5 VSUBS 1.24367f
C137 VP.n5 VSUBS 0.534143f
C138 VP.n6 VSUBS 0.063441f
C139 VP.t2 VSUBS 1.24367f
C140 VP.t0 VSUBS 1.1594f
C141 VP.n7 VSUBS 0.447461f
C142 VP.n8 VSUBS 0.047543f
C143 VP.t6 VSUBS 1.1594f
C144 VP.n9 VSUBS 0.068373f
C145 VP.t9 VSUBS 1.30022f
C146 VP.n10 VSUBS 0.511948f
C147 VP.t1 VSUBS 1.1594f
C148 VP.n11 VSUBS 0.526022f
C149 VP.n12 VSUBS 0.069282f
C150 VP.n13 VSUBS 0.252027f
C151 VP.n14 VSUBS 0.047543f
C152 VP.n15 VSUBS 0.047543f
C153 VP.n16 VSUBS 0.492545f
C154 VP.n17 VSUBS 0.068373f
C155 VP.n18 VSUBS 0.069282f
C156 VP.n19 VSUBS 0.047543f
C157 VP.n20 VSUBS 0.047543f
C158 VP.n21 VSUBS 0.046843f
C159 VP.n22 VSUBS 0.063667f
C160 VP.n23 VSUBS 0.534143f
C161 VP.n24 VSUBS 2.00667f
C162 VP.n25 VSUBS 2.04691f
C163 VP.n26 VSUBS 0.063441f
C164 VP.n27 VSUBS 0.063667f
C165 VP.n28 VSUBS 0.046843f
C166 VP.n29 VSUBS 0.447461f
C167 VP.n30 VSUBS 0.069282f
C168 VP.n31 VSUBS 0.047543f
C169 VP.n32 VSUBS 0.047543f
C170 VP.n33 VSUBS 0.047543f
C171 VP.n34 VSUBS 0.492545f
C172 VP.n35 VSUBS 0.068373f
C173 VP.n36 VSUBS 0.069282f
C174 VP.n37 VSUBS 0.047543f
C175 VP.n38 VSUBS 0.047543f
C176 VP.n39 VSUBS 0.046843f
C177 VP.n40 VSUBS 0.063667f
C178 VP.t4 VSUBS 1.24367f
C179 VP.n41 VSUBS 0.534143f
C180 VP.n42 VSUBS 0.044526f
C181 VDD2.n0 VSUBS 0.027174f
C182 VDD2.n1 VSUBS 0.026249f
C183 VDD2.n2 VSUBS 0.01452f
C184 VDD2.n3 VSUBS 0.033339f
C185 VDD2.n4 VSUBS 0.014935f
C186 VDD2.n5 VSUBS 0.026249f
C187 VDD2.n6 VSUBS 0.014105f
C188 VDD2.n7 VSUBS 0.033339f
C189 VDD2.n8 VSUBS 0.014935f
C190 VDD2.n9 VSUBS 0.026249f
C191 VDD2.n10 VSUBS 0.014105f
C192 VDD2.n11 VSUBS 0.025004f
C193 VDD2.n12 VSUBS 0.025079f
C194 VDD2.t9 VSUBS 0.071587f
C195 VDD2.n13 VSUBS 0.158154f
C196 VDD2.n14 VSUBS 0.81793f
C197 VDD2.n15 VSUBS 0.014105f
C198 VDD2.n16 VSUBS 0.014935f
C199 VDD2.n17 VSUBS 0.033339f
C200 VDD2.n18 VSUBS 0.033339f
C201 VDD2.n19 VSUBS 0.014935f
C202 VDD2.n20 VSUBS 0.014105f
C203 VDD2.n21 VSUBS 0.026249f
C204 VDD2.n22 VSUBS 0.026249f
C205 VDD2.n23 VSUBS 0.014105f
C206 VDD2.n24 VSUBS 0.014935f
C207 VDD2.n25 VSUBS 0.033339f
C208 VDD2.n26 VSUBS 0.033339f
C209 VDD2.n27 VSUBS 0.014935f
C210 VDD2.n28 VSUBS 0.014105f
C211 VDD2.n29 VSUBS 0.026249f
C212 VDD2.n30 VSUBS 0.026249f
C213 VDD2.n31 VSUBS 0.014105f
C214 VDD2.n32 VSUBS 0.014105f
C215 VDD2.n33 VSUBS 0.014935f
C216 VDD2.n34 VSUBS 0.033339f
C217 VDD2.n35 VSUBS 0.033339f
C218 VDD2.n36 VSUBS 0.07503f
C219 VDD2.n37 VSUBS 0.01452f
C220 VDD2.n38 VSUBS 0.014105f
C221 VDD2.n39 VSUBS 0.064258f
C222 VDD2.n40 VSUBS 0.059617f
C223 VDD2.t4 VSUBS 0.163865f
C224 VDD2.t7 VSUBS 0.163865f
C225 VDD2.n41 VSUBS 1.18298f
C226 VDD2.n42 VSUBS 0.732108f
C227 VDD2.t3 VSUBS 0.163865f
C228 VDD2.t5 VSUBS 0.163865f
C229 VDD2.n43 VSUBS 1.18973f
C230 VDD2.n44 VSUBS 2.21634f
C231 VDD2.n45 VSUBS 0.027174f
C232 VDD2.n46 VSUBS 0.026249f
C233 VDD2.n47 VSUBS 0.01452f
C234 VDD2.n48 VSUBS 0.033339f
C235 VDD2.n49 VSUBS 0.014105f
C236 VDD2.n50 VSUBS 0.014935f
C237 VDD2.n51 VSUBS 0.026249f
C238 VDD2.n52 VSUBS 0.014105f
C239 VDD2.n53 VSUBS 0.033339f
C240 VDD2.n54 VSUBS 0.014935f
C241 VDD2.n55 VSUBS 0.026249f
C242 VDD2.n56 VSUBS 0.014105f
C243 VDD2.n57 VSUBS 0.025004f
C244 VDD2.n58 VSUBS 0.025079f
C245 VDD2.t8 VSUBS 0.071587f
C246 VDD2.n59 VSUBS 0.158154f
C247 VDD2.n60 VSUBS 0.81793f
C248 VDD2.n61 VSUBS 0.014105f
C249 VDD2.n62 VSUBS 0.014935f
C250 VDD2.n63 VSUBS 0.033339f
C251 VDD2.n64 VSUBS 0.033339f
C252 VDD2.n65 VSUBS 0.014935f
C253 VDD2.n66 VSUBS 0.014105f
C254 VDD2.n67 VSUBS 0.026249f
C255 VDD2.n68 VSUBS 0.026249f
C256 VDD2.n69 VSUBS 0.014105f
C257 VDD2.n70 VSUBS 0.014935f
C258 VDD2.n71 VSUBS 0.033339f
C259 VDD2.n72 VSUBS 0.033339f
C260 VDD2.n73 VSUBS 0.014935f
C261 VDD2.n74 VSUBS 0.014105f
C262 VDD2.n75 VSUBS 0.026249f
C263 VDD2.n76 VSUBS 0.026249f
C264 VDD2.n77 VSUBS 0.014105f
C265 VDD2.n78 VSUBS 0.014935f
C266 VDD2.n79 VSUBS 0.033339f
C267 VDD2.n80 VSUBS 0.033339f
C268 VDD2.n81 VSUBS 0.07503f
C269 VDD2.n82 VSUBS 0.01452f
C270 VDD2.n83 VSUBS 0.014105f
C271 VDD2.n84 VSUBS 0.064258f
C272 VDD2.n85 VSUBS 0.055684f
C273 VDD2.n86 VSUBS 2.10804f
C274 VDD2.t1 VSUBS 0.163865f
C275 VDD2.t6 VSUBS 0.163865f
C276 VDD2.n87 VSUBS 1.18298f
C277 VDD2.n88 VSUBS 0.582821f
C278 VDD2.t0 VSUBS 0.163865f
C279 VDD2.t2 VSUBS 0.163865f
C280 VDD2.n89 VSUBS 1.1897f
C281 VTAIL.t13 VSUBS 0.185885f
C282 VTAIL.t17 VSUBS 0.185885f
C283 VTAIL.n0 VSUBS 1.21939f
C284 VTAIL.n1 VSUBS 0.788311f
C285 VTAIL.n2 VSUBS 0.030826f
C286 VTAIL.n3 VSUBS 0.029776f
C287 VTAIL.n4 VSUBS 0.016471f
C288 VTAIL.n5 VSUBS 0.037819f
C289 VTAIL.n6 VSUBS 0.016941f
C290 VTAIL.n7 VSUBS 0.029776f
C291 VTAIL.n8 VSUBS 0.016f
C292 VTAIL.n9 VSUBS 0.037819f
C293 VTAIL.n10 VSUBS 0.016941f
C294 VTAIL.n11 VSUBS 0.029776f
C295 VTAIL.n12 VSUBS 0.016f
C296 VTAIL.n13 VSUBS 0.028364f
C297 VTAIL.n14 VSUBS 0.028449f
C298 VTAIL.t6 VSUBS 0.081207f
C299 VTAIL.n15 VSUBS 0.179406f
C300 VTAIL.n16 VSUBS 0.927842f
C301 VTAIL.n17 VSUBS 0.016f
C302 VTAIL.n18 VSUBS 0.016941f
C303 VTAIL.n19 VSUBS 0.037819f
C304 VTAIL.n20 VSUBS 0.037819f
C305 VTAIL.n21 VSUBS 0.016941f
C306 VTAIL.n22 VSUBS 0.016f
C307 VTAIL.n23 VSUBS 0.029776f
C308 VTAIL.n24 VSUBS 0.029776f
C309 VTAIL.n25 VSUBS 0.016f
C310 VTAIL.n26 VSUBS 0.016941f
C311 VTAIL.n27 VSUBS 0.037819f
C312 VTAIL.n28 VSUBS 0.037819f
C313 VTAIL.n29 VSUBS 0.016941f
C314 VTAIL.n30 VSUBS 0.016f
C315 VTAIL.n31 VSUBS 0.029776f
C316 VTAIL.n32 VSUBS 0.029776f
C317 VTAIL.n33 VSUBS 0.016f
C318 VTAIL.n34 VSUBS 0.016f
C319 VTAIL.n35 VSUBS 0.016941f
C320 VTAIL.n36 VSUBS 0.037819f
C321 VTAIL.n37 VSUBS 0.037819f
C322 VTAIL.n38 VSUBS 0.085112f
C323 VTAIL.n39 VSUBS 0.016471f
C324 VTAIL.n40 VSUBS 0.016f
C325 VTAIL.n41 VSUBS 0.072893f
C326 VTAIL.n42 VSUBS 0.042638f
C327 VTAIL.n43 VSUBS 0.256425f
C328 VTAIL.t5 VSUBS 0.185885f
C329 VTAIL.t8 VSUBS 0.185885f
C330 VTAIL.n44 VSUBS 1.21939f
C331 VTAIL.n45 VSUBS 0.82946f
C332 VTAIL.t9 VSUBS 0.185885f
C333 VTAIL.t7 VSUBS 0.185885f
C334 VTAIL.n46 VSUBS 1.21939f
C335 VTAIL.n47 VSUBS 2.00976f
C336 VTAIL.t14 VSUBS 0.185885f
C337 VTAIL.t12 VSUBS 0.185885f
C338 VTAIL.n48 VSUBS 1.21939f
C339 VTAIL.n49 VSUBS 2.00975f
C340 VTAIL.t10 VSUBS 0.185885f
C341 VTAIL.t19 VSUBS 0.185885f
C342 VTAIL.n50 VSUBS 1.21939f
C343 VTAIL.n51 VSUBS 0.829451f
C344 VTAIL.n52 VSUBS 0.030826f
C345 VTAIL.n53 VSUBS 0.029776f
C346 VTAIL.n54 VSUBS 0.016471f
C347 VTAIL.n55 VSUBS 0.037819f
C348 VTAIL.n56 VSUBS 0.016f
C349 VTAIL.n57 VSUBS 0.016941f
C350 VTAIL.n58 VSUBS 0.029776f
C351 VTAIL.n59 VSUBS 0.016f
C352 VTAIL.n60 VSUBS 0.037819f
C353 VTAIL.n61 VSUBS 0.016941f
C354 VTAIL.n62 VSUBS 0.029776f
C355 VTAIL.n63 VSUBS 0.016f
C356 VTAIL.n64 VSUBS 0.028364f
C357 VTAIL.n65 VSUBS 0.028449f
C358 VTAIL.t11 VSUBS 0.081207f
C359 VTAIL.n66 VSUBS 0.179406f
C360 VTAIL.n67 VSUBS 0.927842f
C361 VTAIL.n68 VSUBS 0.016f
C362 VTAIL.n69 VSUBS 0.016941f
C363 VTAIL.n70 VSUBS 0.037819f
C364 VTAIL.n71 VSUBS 0.037819f
C365 VTAIL.n72 VSUBS 0.016941f
C366 VTAIL.n73 VSUBS 0.016f
C367 VTAIL.n74 VSUBS 0.029776f
C368 VTAIL.n75 VSUBS 0.029776f
C369 VTAIL.n76 VSUBS 0.016f
C370 VTAIL.n77 VSUBS 0.016941f
C371 VTAIL.n78 VSUBS 0.037819f
C372 VTAIL.n79 VSUBS 0.037819f
C373 VTAIL.n80 VSUBS 0.016941f
C374 VTAIL.n81 VSUBS 0.016f
C375 VTAIL.n82 VSUBS 0.029776f
C376 VTAIL.n83 VSUBS 0.029776f
C377 VTAIL.n84 VSUBS 0.016f
C378 VTAIL.n85 VSUBS 0.016941f
C379 VTAIL.n86 VSUBS 0.037819f
C380 VTAIL.n87 VSUBS 0.037819f
C381 VTAIL.n88 VSUBS 0.085112f
C382 VTAIL.n89 VSUBS 0.016471f
C383 VTAIL.n90 VSUBS 0.016f
C384 VTAIL.n91 VSUBS 0.072893f
C385 VTAIL.n92 VSUBS 0.042638f
C386 VTAIL.n93 VSUBS 0.256425f
C387 VTAIL.t0 VSUBS 0.185885f
C388 VTAIL.t2 VSUBS 0.185885f
C389 VTAIL.n94 VSUBS 1.21939f
C390 VTAIL.n95 VSUBS 0.813322f
C391 VTAIL.t4 VSUBS 0.185885f
C392 VTAIL.t3 VSUBS 0.185885f
C393 VTAIL.n96 VSUBS 1.21939f
C394 VTAIL.n97 VSUBS 0.829451f
C395 VTAIL.n98 VSUBS 0.030826f
C396 VTAIL.n99 VSUBS 0.029776f
C397 VTAIL.n100 VSUBS 0.016471f
C398 VTAIL.n101 VSUBS 0.037819f
C399 VTAIL.n102 VSUBS 0.016f
C400 VTAIL.n103 VSUBS 0.016941f
C401 VTAIL.n104 VSUBS 0.029776f
C402 VTAIL.n105 VSUBS 0.016f
C403 VTAIL.n106 VSUBS 0.037819f
C404 VTAIL.n107 VSUBS 0.016941f
C405 VTAIL.n108 VSUBS 0.029776f
C406 VTAIL.n109 VSUBS 0.016f
C407 VTAIL.n110 VSUBS 0.028364f
C408 VTAIL.n111 VSUBS 0.028449f
C409 VTAIL.t1 VSUBS 0.081207f
C410 VTAIL.n112 VSUBS 0.179406f
C411 VTAIL.n113 VSUBS 0.927842f
C412 VTAIL.n114 VSUBS 0.016f
C413 VTAIL.n115 VSUBS 0.016941f
C414 VTAIL.n116 VSUBS 0.037819f
C415 VTAIL.n117 VSUBS 0.037819f
C416 VTAIL.n118 VSUBS 0.016941f
C417 VTAIL.n119 VSUBS 0.016f
C418 VTAIL.n120 VSUBS 0.029776f
C419 VTAIL.n121 VSUBS 0.029776f
C420 VTAIL.n122 VSUBS 0.016f
C421 VTAIL.n123 VSUBS 0.016941f
C422 VTAIL.n124 VSUBS 0.037819f
C423 VTAIL.n125 VSUBS 0.037819f
C424 VTAIL.n126 VSUBS 0.016941f
C425 VTAIL.n127 VSUBS 0.016f
C426 VTAIL.n128 VSUBS 0.029776f
C427 VTAIL.n129 VSUBS 0.029776f
C428 VTAIL.n130 VSUBS 0.016f
C429 VTAIL.n131 VSUBS 0.016941f
C430 VTAIL.n132 VSUBS 0.037819f
C431 VTAIL.n133 VSUBS 0.037819f
C432 VTAIL.n134 VSUBS 0.085112f
C433 VTAIL.n135 VSUBS 0.016471f
C434 VTAIL.n136 VSUBS 0.016f
C435 VTAIL.n137 VSUBS 0.072893f
C436 VTAIL.n138 VSUBS 0.042638f
C437 VTAIL.n139 VSUBS 1.33044f
C438 VTAIL.n140 VSUBS 0.030826f
C439 VTAIL.n141 VSUBS 0.029776f
C440 VTAIL.n142 VSUBS 0.016471f
C441 VTAIL.n143 VSUBS 0.037819f
C442 VTAIL.n144 VSUBS 0.016941f
C443 VTAIL.n145 VSUBS 0.029776f
C444 VTAIL.n146 VSUBS 0.016f
C445 VTAIL.n147 VSUBS 0.037819f
C446 VTAIL.n148 VSUBS 0.016941f
C447 VTAIL.n149 VSUBS 0.029776f
C448 VTAIL.n150 VSUBS 0.016f
C449 VTAIL.n151 VSUBS 0.028364f
C450 VTAIL.n152 VSUBS 0.028449f
C451 VTAIL.t16 VSUBS 0.081207f
C452 VTAIL.n153 VSUBS 0.179406f
C453 VTAIL.n154 VSUBS 0.927842f
C454 VTAIL.n155 VSUBS 0.016f
C455 VTAIL.n156 VSUBS 0.016941f
C456 VTAIL.n157 VSUBS 0.037819f
C457 VTAIL.n158 VSUBS 0.037819f
C458 VTAIL.n159 VSUBS 0.016941f
C459 VTAIL.n160 VSUBS 0.016f
C460 VTAIL.n161 VSUBS 0.029776f
C461 VTAIL.n162 VSUBS 0.029776f
C462 VTAIL.n163 VSUBS 0.016f
C463 VTAIL.n164 VSUBS 0.016941f
C464 VTAIL.n165 VSUBS 0.037819f
C465 VTAIL.n166 VSUBS 0.037819f
C466 VTAIL.n167 VSUBS 0.016941f
C467 VTAIL.n168 VSUBS 0.016f
C468 VTAIL.n169 VSUBS 0.029776f
C469 VTAIL.n170 VSUBS 0.029776f
C470 VTAIL.n171 VSUBS 0.016f
C471 VTAIL.n172 VSUBS 0.016f
C472 VTAIL.n173 VSUBS 0.016941f
C473 VTAIL.n174 VSUBS 0.037819f
C474 VTAIL.n175 VSUBS 0.037819f
C475 VTAIL.n176 VSUBS 0.085112f
C476 VTAIL.n177 VSUBS 0.016471f
C477 VTAIL.n178 VSUBS 0.016f
C478 VTAIL.n179 VSUBS 0.072893f
C479 VTAIL.n180 VSUBS 0.042638f
C480 VTAIL.n181 VSUBS 1.33044f
C481 VTAIL.t15 VSUBS 0.185885f
C482 VTAIL.t18 VSUBS 0.185885f
C483 VTAIL.n182 VSUBS 1.21939f
C484 VTAIL.n183 VSUBS 0.732068f
C485 VN.n0 VSUBS 0.061607f
C486 VN.t6 VSUBS 1.12588f
C487 VN.n1 VSUBS 0.434525f
C488 VN.n2 VSUBS 0.046169f
C489 VN.t2 VSUBS 1.12588f
C490 VN.n3 VSUBS 0.066396f
C491 VN.t0 VSUBS 1.26263f
C492 VN.n4 VSUBS 0.497149f
C493 VN.t5 VSUBS 1.12588f
C494 VN.n5 VSUBS 0.510815f
C495 VN.n6 VSUBS 0.067279f
C496 VN.n7 VSUBS 0.244741f
C497 VN.n8 VSUBS 0.046169f
C498 VN.n9 VSUBS 0.046169f
C499 VN.n10 VSUBS 0.478306f
C500 VN.n11 VSUBS 0.066396f
C501 VN.n12 VSUBS 0.067279f
C502 VN.n13 VSUBS 0.046169f
C503 VN.n14 VSUBS 0.046169f
C504 VN.n15 VSUBS 0.045489f
C505 VN.n16 VSUBS 0.061826f
C506 VN.t4 VSUBS 1.20772f
C507 VN.n17 VSUBS 0.518701f
C508 VN.n18 VSUBS 0.043239f
C509 VN.n19 VSUBS 0.061607f
C510 VN.t8 VSUBS 1.12588f
C511 VN.n20 VSUBS 0.434525f
C512 VN.n21 VSUBS 0.046169f
C513 VN.t3 VSUBS 1.12588f
C514 VN.n22 VSUBS 0.066396f
C515 VN.t7 VSUBS 1.26263f
C516 VN.n23 VSUBS 0.497149f
C517 VN.t9 VSUBS 1.12588f
C518 VN.n24 VSUBS 0.510815f
C519 VN.n25 VSUBS 0.067279f
C520 VN.n26 VSUBS 0.244741f
C521 VN.n27 VSUBS 0.046169f
C522 VN.n28 VSUBS 0.046169f
C523 VN.n29 VSUBS 0.478306f
C524 VN.n30 VSUBS 0.066396f
C525 VN.n31 VSUBS 0.067279f
C526 VN.n32 VSUBS 0.046169f
C527 VN.n33 VSUBS 0.046169f
C528 VN.n34 VSUBS 0.045489f
C529 VN.n35 VSUBS 0.061826f
C530 VN.t1 VSUBS 1.20772f
C531 VN.n36 VSUBS 0.518701f
C532 VN.n37 VSUBS 1.97452f
C533 B.n0 VSUBS 0.004845f
C534 B.n1 VSUBS 0.004845f
C535 B.n2 VSUBS 0.007662f
C536 B.n3 VSUBS 0.007662f
C537 B.n4 VSUBS 0.007662f
C538 B.n5 VSUBS 0.007662f
C539 B.n6 VSUBS 0.007662f
C540 B.n7 VSUBS 0.007662f
C541 B.n8 VSUBS 0.007662f
C542 B.n9 VSUBS 0.007662f
C543 B.n10 VSUBS 0.007662f
C544 B.n11 VSUBS 0.007662f
C545 B.n12 VSUBS 0.007662f
C546 B.n13 VSUBS 0.007662f
C547 B.n14 VSUBS 0.007662f
C548 B.n15 VSUBS 0.007662f
C549 B.n16 VSUBS 0.007662f
C550 B.n17 VSUBS 0.007662f
C551 B.n18 VSUBS 0.007662f
C552 B.n19 VSUBS 0.018845f
C553 B.n20 VSUBS 0.007662f
C554 B.n21 VSUBS 0.007662f
C555 B.n22 VSUBS 0.007662f
C556 B.n23 VSUBS 0.007662f
C557 B.n24 VSUBS 0.007662f
C558 B.n25 VSUBS 0.007662f
C559 B.n26 VSUBS 0.007662f
C560 B.n27 VSUBS 0.007662f
C561 B.n28 VSUBS 0.007662f
C562 B.n29 VSUBS 0.007662f
C563 B.n30 VSUBS 0.007662f
C564 B.n31 VSUBS 0.007662f
C565 B.n32 VSUBS 0.007662f
C566 B.n33 VSUBS 0.007662f
C567 B.t8 VSUBS 0.136281f
C568 B.t7 VSUBS 0.152835f
C569 B.t6 VSUBS 0.438651f
C570 B.n34 VSUBS 0.254122f
C571 B.n35 VSUBS 0.201513f
C572 B.n36 VSUBS 0.017752f
C573 B.n37 VSUBS 0.007662f
C574 B.n38 VSUBS 0.007662f
C575 B.n39 VSUBS 0.007662f
C576 B.n40 VSUBS 0.007662f
C577 B.n41 VSUBS 0.007662f
C578 B.t5 VSUBS 0.136283f
C579 B.t4 VSUBS 0.152837f
C580 B.t3 VSUBS 0.438651f
C581 B.n42 VSUBS 0.25412f
C582 B.n43 VSUBS 0.20151f
C583 B.n44 VSUBS 0.007662f
C584 B.n45 VSUBS 0.007662f
C585 B.n46 VSUBS 0.007662f
C586 B.n47 VSUBS 0.007662f
C587 B.n48 VSUBS 0.007662f
C588 B.n49 VSUBS 0.007662f
C589 B.n50 VSUBS 0.007662f
C590 B.n51 VSUBS 0.007662f
C591 B.n52 VSUBS 0.007662f
C592 B.n53 VSUBS 0.007662f
C593 B.n54 VSUBS 0.007662f
C594 B.n55 VSUBS 0.007662f
C595 B.n56 VSUBS 0.007662f
C596 B.n57 VSUBS 0.007662f
C597 B.n58 VSUBS 0.018325f
C598 B.n59 VSUBS 0.007662f
C599 B.n60 VSUBS 0.007662f
C600 B.n61 VSUBS 0.007662f
C601 B.n62 VSUBS 0.007662f
C602 B.n63 VSUBS 0.007662f
C603 B.n64 VSUBS 0.007662f
C604 B.n65 VSUBS 0.007662f
C605 B.n66 VSUBS 0.007662f
C606 B.n67 VSUBS 0.007662f
C607 B.n68 VSUBS 0.007662f
C608 B.n69 VSUBS 0.007662f
C609 B.n70 VSUBS 0.007662f
C610 B.n71 VSUBS 0.007662f
C611 B.n72 VSUBS 0.007662f
C612 B.n73 VSUBS 0.007662f
C613 B.n74 VSUBS 0.007662f
C614 B.n75 VSUBS 0.007662f
C615 B.n76 VSUBS 0.007662f
C616 B.n77 VSUBS 0.007662f
C617 B.n78 VSUBS 0.007662f
C618 B.n79 VSUBS 0.007662f
C619 B.n80 VSUBS 0.007662f
C620 B.n81 VSUBS 0.007662f
C621 B.n82 VSUBS 0.007662f
C622 B.n83 VSUBS 0.007662f
C623 B.n84 VSUBS 0.007662f
C624 B.n85 VSUBS 0.007662f
C625 B.n86 VSUBS 0.007662f
C626 B.n87 VSUBS 0.007662f
C627 B.n88 VSUBS 0.007662f
C628 B.n89 VSUBS 0.007662f
C629 B.n90 VSUBS 0.007662f
C630 B.n91 VSUBS 0.007662f
C631 B.n92 VSUBS 0.017436f
C632 B.n93 VSUBS 0.007662f
C633 B.n94 VSUBS 0.007662f
C634 B.n95 VSUBS 0.007662f
C635 B.n96 VSUBS 0.007662f
C636 B.n97 VSUBS 0.007662f
C637 B.n98 VSUBS 0.007662f
C638 B.n99 VSUBS 0.007662f
C639 B.n100 VSUBS 0.007662f
C640 B.n101 VSUBS 0.007662f
C641 B.n102 VSUBS 0.007662f
C642 B.n103 VSUBS 0.007662f
C643 B.n104 VSUBS 0.007662f
C644 B.n105 VSUBS 0.007662f
C645 B.n106 VSUBS 0.007662f
C646 B.n107 VSUBS 0.007662f
C647 B.t1 VSUBS 0.136283f
C648 B.t2 VSUBS 0.152837f
C649 B.t0 VSUBS 0.438651f
C650 B.n108 VSUBS 0.25412f
C651 B.n109 VSUBS 0.20151f
C652 B.n110 VSUBS 0.007662f
C653 B.n111 VSUBS 0.007662f
C654 B.n112 VSUBS 0.007662f
C655 B.n113 VSUBS 0.007662f
C656 B.t10 VSUBS 0.136281f
C657 B.t11 VSUBS 0.152835f
C658 B.t9 VSUBS 0.438651f
C659 B.n114 VSUBS 0.254122f
C660 B.n115 VSUBS 0.201513f
C661 B.n116 VSUBS 0.017752f
C662 B.n117 VSUBS 0.007662f
C663 B.n118 VSUBS 0.007662f
C664 B.n119 VSUBS 0.007662f
C665 B.n120 VSUBS 0.007662f
C666 B.n121 VSUBS 0.007662f
C667 B.n122 VSUBS 0.007662f
C668 B.n123 VSUBS 0.007662f
C669 B.n124 VSUBS 0.007662f
C670 B.n125 VSUBS 0.007662f
C671 B.n126 VSUBS 0.007662f
C672 B.n127 VSUBS 0.007662f
C673 B.n128 VSUBS 0.007662f
C674 B.n129 VSUBS 0.007662f
C675 B.n130 VSUBS 0.007662f
C676 B.n131 VSUBS 0.018845f
C677 B.n132 VSUBS 0.007662f
C678 B.n133 VSUBS 0.007662f
C679 B.n134 VSUBS 0.007662f
C680 B.n135 VSUBS 0.007662f
C681 B.n136 VSUBS 0.007662f
C682 B.n137 VSUBS 0.007662f
C683 B.n138 VSUBS 0.007662f
C684 B.n139 VSUBS 0.007662f
C685 B.n140 VSUBS 0.007662f
C686 B.n141 VSUBS 0.007662f
C687 B.n142 VSUBS 0.007662f
C688 B.n143 VSUBS 0.007662f
C689 B.n144 VSUBS 0.007662f
C690 B.n145 VSUBS 0.007662f
C691 B.n146 VSUBS 0.007662f
C692 B.n147 VSUBS 0.007662f
C693 B.n148 VSUBS 0.007662f
C694 B.n149 VSUBS 0.007662f
C695 B.n150 VSUBS 0.007662f
C696 B.n151 VSUBS 0.007662f
C697 B.n152 VSUBS 0.007662f
C698 B.n153 VSUBS 0.007662f
C699 B.n154 VSUBS 0.007662f
C700 B.n155 VSUBS 0.007662f
C701 B.n156 VSUBS 0.007662f
C702 B.n157 VSUBS 0.007662f
C703 B.n158 VSUBS 0.007662f
C704 B.n159 VSUBS 0.007662f
C705 B.n160 VSUBS 0.007662f
C706 B.n161 VSUBS 0.007662f
C707 B.n162 VSUBS 0.007662f
C708 B.n163 VSUBS 0.007662f
C709 B.n164 VSUBS 0.007662f
C710 B.n165 VSUBS 0.007662f
C711 B.n166 VSUBS 0.007662f
C712 B.n167 VSUBS 0.007662f
C713 B.n168 VSUBS 0.007662f
C714 B.n169 VSUBS 0.007662f
C715 B.n170 VSUBS 0.007662f
C716 B.n171 VSUBS 0.007662f
C717 B.n172 VSUBS 0.007662f
C718 B.n173 VSUBS 0.007662f
C719 B.n174 VSUBS 0.007662f
C720 B.n175 VSUBS 0.007662f
C721 B.n176 VSUBS 0.007662f
C722 B.n177 VSUBS 0.007662f
C723 B.n178 VSUBS 0.007662f
C724 B.n179 VSUBS 0.007662f
C725 B.n180 VSUBS 0.007662f
C726 B.n181 VSUBS 0.007662f
C727 B.n182 VSUBS 0.007662f
C728 B.n183 VSUBS 0.007662f
C729 B.n184 VSUBS 0.007662f
C730 B.n185 VSUBS 0.007662f
C731 B.n186 VSUBS 0.007662f
C732 B.n187 VSUBS 0.007662f
C733 B.n188 VSUBS 0.007662f
C734 B.n189 VSUBS 0.007662f
C735 B.n190 VSUBS 0.007662f
C736 B.n191 VSUBS 0.007662f
C737 B.n192 VSUBS 0.007662f
C738 B.n193 VSUBS 0.007662f
C739 B.n194 VSUBS 0.007662f
C740 B.n195 VSUBS 0.007662f
C741 B.n196 VSUBS 0.017436f
C742 B.n197 VSUBS 0.017436f
C743 B.n198 VSUBS 0.018845f
C744 B.n199 VSUBS 0.007662f
C745 B.n200 VSUBS 0.007662f
C746 B.n201 VSUBS 0.007662f
C747 B.n202 VSUBS 0.007662f
C748 B.n203 VSUBS 0.007662f
C749 B.n204 VSUBS 0.007662f
C750 B.n205 VSUBS 0.007662f
C751 B.n206 VSUBS 0.007662f
C752 B.n207 VSUBS 0.007662f
C753 B.n208 VSUBS 0.007662f
C754 B.n209 VSUBS 0.007662f
C755 B.n210 VSUBS 0.007662f
C756 B.n211 VSUBS 0.007662f
C757 B.n212 VSUBS 0.007662f
C758 B.n213 VSUBS 0.007662f
C759 B.n214 VSUBS 0.007662f
C760 B.n215 VSUBS 0.007662f
C761 B.n216 VSUBS 0.007662f
C762 B.n217 VSUBS 0.007662f
C763 B.n218 VSUBS 0.007662f
C764 B.n219 VSUBS 0.007662f
C765 B.n220 VSUBS 0.007662f
C766 B.n221 VSUBS 0.007662f
C767 B.n222 VSUBS 0.007662f
C768 B.n223 VSUBS 0.007662f
C769 B.n224 VSUBS 0.007662f
C770 B.n225 VSUBS 0.007662f
C771 B.n226 VSUBS 0.007662f
C772 B.n227 VSUBS 0.007662f
C773 B.n228 VSUBS 0.007662f
C774 B.n229 VSUBS 0.007662f
C775 B.n230 VSUBS 0.007662f
C776 B.n231 VSUBS 0.007662f
C777 B.n232 VSUBS 0.007662f
C778 B.n233 VSUBS 0.007662f
C779 B.n234 VSUBS 0.007662f
C780 B.n235 VSUBS 0.007662f
C781 B.n236 VSUBS 0.007662f
C782 B.n237 VSUBS 0.007662f
C783 B.n238 VSUBS 0.007662f
C784 B.n239 VSUBS 0.007662f
C785 B.n240 VSUBS 0.007662f
C786 B.n241 VSUBS 0.005296f
C787 B.n242 VSUBS 0.007662f
C788 B.n243 VSUBS 0.007662f
C789 B.n244 VSUBS 0.006197f
C790 B.n245 VSUBS 0.007662f
C791 B.n246 VSUBS 0.007662f
C792 B.n247 VSUBS 0.007662f
C793 B.n248 VSUBS 0.007662f
C794 B.n249 VSUBS 0.007662f
C795 B.n250 VSUBS 0.007662f
C796 B.n251 VSUBS 0.007662f
C797 B.n252 VSUBS 0.007662f
C798 B.n253 VSUBS 0.007662f
C799 B.n254 VSUBS 0.007662f
C800 B.n255 VSUBS 0.007662f
C801 B.n256 VSUBS 0.006197f
C802 B.n257 VSUBS 0.017752f
C803 B.n258 VSUBS 0.005296f
C804 B.n259 VSUBS 0.007662f
C805 B.n260 VSUBS 0.007662f
C806 B.n261 VSUBS 0.007662f
C807 B.n262 VSUBS 0.007662f
C808 B.n263 VSUBS 0.007662f
C809 B.n264 VSUBS 0.007662f
C810 B.n265 VSUBS 0.007662f
C811 B.n266 VSUBS 0.007662f
C812 B.n267 VSUBS 0.007662f
C813 B.n268 VSUBS 0.007662f
C814 B.n269 VSUBS 0.007662f
C815 B.n270 VSUBS 0.007662f
C816 B.n271 VSUBS 0.007662f
C817 B.n272 VSUBS 0.007662f
C818 B.n273 VSUBS 0.007662f
C819 B.n274 VSUBS 0.007662f
C820 B.n275 VSUBS 0.007662f
C821 B.n276 VSUBS 0.007662f
C822 B.n277 VSUBS 0.007662f
C823 B.n278 VSUBS 0.007662f
C824 B.n279 VSUBS 0.007662f
C825 B.n280 VSUBS 0.007662f
C826 B.n281 VSUBS 0.007662f
C827 B.n282 VSUBS 0.007662f
C828 B.n283 VSUBS 0.007662f
C829 B.n284 VSUBS 0.007662f
C830 B.n285 VSUBS 0.007662f
C831 B.n286 VSUBS 0.007662f
C832 B.n287 VSUBS 0.007662f
C833 B.n288 VSUBS 0.007662f
C834 B.n289 VSUBS 0.007662f
C835 B.n290 VSUBS 0.007662f
C836 B.n291 VSUBS 0.007662f
C837 B.n292 VSUBS 0.007662f
C838 B.n293 VSUBS 0.007662f
C839 B.n294 VSUBS 0.007662f
C840 B.n295 VSUBS 0.007662f
C841 B.n296 VSUBS 0.007662f
C842 B.n297 VSUBS 0.007662f
C843 B.n298 VSUBS 0.007662f
C844 B.n299 VSUBS 0.007662f
C845 B.n300 VSUBS 0.007662f
C846 B.n301 VSUBS 0.018845f
C847 B.n302 VSUBS 0.018845f
C848 B.n303 VSUBS 0.017436f
C849 B.n304 VSUBS 0.007662f
C850 B.n305 VSUBS 0.007662f
C851 B.n306 VSUBS 0.007662f
C852 B.n307 VSUBS 0.007662f
C853 B.n308 VSUBS 0.007662f
C854 B.n309 VSUBS 0.007662f
C855 B.n310 VSUBS 0.007662f
C856 B.n311 VSUBS 0.007662f
C857 B.n312 VSUBS 0.007662f
C858 B.n313 VSUBS 0.007662f
C859 B.n314 VSUBS 0.007662f
C860 B.n315 VSUBS 0.007662f
C861 B.n316 VSUBS 0.007662f
C862 B.n317 VSUBS 0.007662f
C863 B.n318 VSUBS 0.007662f
C864 B.n319 VSUBS 0.007662f
C865 B.n320 VSUBS 0.007662f
C866 B.n321 VSUBS 0.007662f
C867 B.n322 VSUBS 0.007662f
C868 B.n323 VSUBS 0.007662f
C869 B.n324 VSUBS 0.007662f
C870 B.n325 VSUBS 0.007662f
C871 B.n326 VSUBS 0.007662f
C872 B.n327 VSUBS 0.007662f
C873 B.n328 VSUBS 0.007662f
C874 B.n329 VSUBS 0.007662f
C875 B.n330 VSUBS 0.007662f
C876 B.n331 VSUBS 0.007662f
C877 B.n332 VSUBS 0.007662f
C878 B.n333 VSUBS 0.007662f
C879 B.n334 VSUBS 0.007662f
C880 B.n335 VSUBS 0.007662f
C881 B.n336 VSUBS 0.007662f
C882 B.n337 VSUBS 0.007662f
C883 B.n338 VSUBS 0.007662f
C884 B.n339 VSUBS 0.007662f
C885 B.n340 VSUBS 0.007662f
C886 B.n341 VSUBS 0.007662f
C887 B.n342 VSUBS 0.007662f
C888 B.n343 VSUBS 0.007662f
C889 B.n344 VSUBS 0.007662f
C890 B.n345 VSUBS 0.007662f
C891 B.n346 VSUBS 0.007662f
C892 B.n347 VSUBS 0.007662f
C893 B.n348 VSUBS 0.007662f
C894 B.n349 VSUBS 0.007662f
C895 B.n350 VSUBS 0.007662f
C896 B.n351 VSUBS 0.007662f
C897 B.n352 VSUBS 0.007662f
C898 B.n353 VSUBS 0.007662f
C899 B.n354 VSUBS 0.007662f
C900 B.n355 VSUBS 0.007662f
C901 B.n356 VSUBS 0.007662f
C902 B.n357 VSUBS 0.007662f
C903 B.n358 VSUBS 0.007662f
C904 B.n359 VSUBS 0.007662f
C905 B.n360 VSUBS 0.007662f
C906 B.n361 VSUBS 0.007662f
C907 B.n362 VSUBS 0.007662f
C908 B.n363 VSUBS 0.007662f
C909 B.n364 VSUBS 0.007662f
C910 B.n365 VSUBS 0.007662f
C911 B.n366 VSUBS 0.007662f
C912 B.n367 VSUBS 0.007662f
C913 B.n368 VSUBS 0.007662f
C914 B.n369 VSUBS 0.007662f
C915 B.n370 VSUBS 0.007662f
C916 B.n371 VSUBS 0.007662f
C917 B.n372 VSUBS 0.007662f
C918 B.n373 VSUBS 0.007662f
C919 B.n374 VSUBS 0.007662f
C920 B.n375 VSUBS 0.007662f
C921 B.n376 VSUBS 0.007662f
C922 B.n377 VSUBS 0.007662f
C923 B.n378 VSUBS 0.007662f
C924 B.n379 VSUBS 0.007662f
C925 B.n380 VSUBS 0.007662f
C926 B.n381 VSUBS 0.007662f
C927 B.n382 VSUBS 0.007662f
C928 B.n383 VSUBS 0.007662f
C929 B.n384 VSUBS 0.007662f
C930 B.n385 VSUBS 0.007662f
C931 B.n386 VSUBS 0.007662f
C932 B.n387 VSUBS 0.007662f
C933 B.n388 VSUBS 0.007662f
C934 B.n389 VSUBS 0.007662f
C935 B.n390 VSUBS 0.007662f
C936 B.n391 VSUBS 0.007662f
C937 B.n392 VSUBS 0.007662f
C938 B.n393 VSUBS 0.007662f
C939 B.n394 VSUBS 0.007662f
C940 B.n395 VSUBS 0.007662f
C941 B.n396 VSUBS 0.007662f
C942 B.n397 VSUBS 0.007662f
C943 B.n398 VSUBS 0.007662f
C944 B.n399 VSUBS 0.007662f
C945 B.n400 VSUBS 0.007662f
C946 B.n401 VSUBS 0.007662f
C947 B.n402 VSUBS 0.007662f
C948 B.n403 VSUBS 0.007662f
C949 B.n404 VSUBS 0.007662f
C950 B.n405 VSUBS 0.017436f
C951 B.n406 VSUBS 0.018845f
C952 B.n407 VSUBS 0.017956f
C953 B.n408 VSUBS 0.007662f
C954 B.n409 VSUBS 0.007662f
C955 B.n410 VSUBS 0.007662f
C956 B.n411 VSUBS 0.007662f
C957 B.n412 VSUBS 0.007662f
C958 B.n413 VSUBS 0.007662f
C959 B.n414 VSUBS 0.007662f
C960 B.n415 VSUBS 0.007662f
C961 B.n416 VSUBS 0.007662f
C962 B.n417 VSUBS 0.007662f
C963 B.n418 VSUBS 0.007662f
C964 B.n419 VSUBS 0.007662f
C965 B.n420 VSUBS 0.007662f
C966 B.n421 VSUBS 0.007662f
C967 B.n422 VSUBS 0.007662f
C968 B.n423 VSUBS 0.007662f
C969 B.n424 VSUBS 0.007662f
C970 B.n425 VSUBS 0.007662f
C971 B.n426 VSUBS 0.007662f
C972 B.n427 VSUBS 0.007662f
C973 B.n428 VSUBS 0.007662f
C974 B.n429 VSUBS 0.007662f
C975 B.n430 VSUBS 0.007662f
C976 B.n431 VSUBS 0.007662f
C977 B.n432 VSUBS 0.007662f
C978 B.n433 VSUBS 0.007662f
C979 B.n434 VSUBS 0.007662f
C980 B.n435 VSUBS 0.007662f
C981 B.n436 VSUBS 0.007662f
C982 B.n437 VSUBS 0.007662f
C983 B.n438 VSUBS 0.007662f
C984 B.n439 VSUBS 0.007662f
C985 B.n440 VSUBS 0.007662f
C986 B.n441 VSUBS 0.007662f
C987 B.n442 VSUBS 0.007662f
C988 B.n443 VSUBS 0.007662f
C989 B.n444 VSUBS 0.007662f
C990 B.n445 VSUBS 0.007662f
C991 B.n446 VSUBS 0.007662f
C992 B.n447 VSUBS 0.007662f
C993 B.n448 VSUBS 0.007662f
C994 B.n449 VSUBS 0.007662f
C995 B.n450 VSUBS 0.005296f
C996 B.n451 VSUBS 0.017752f
C997 B.n452 VSUBS 0.006197f
C998 B.n453 VSUBS 0.007662f
C999 B.n454 VSUBS 0.007662f
C1000 B.n455 VSUBS 0.007662f
C1001 B.n456 VSUBS 0.007662f
C1002 B.n457 VSUBS 0.007662f
C1003 B.n458 VSUBS 0.007662f
C1004 B.n459 VSUBS 0.007662f
C1005 B.n460 VSUBS 0.007662f
C1006 B.n461 VSUBS 0.007662f
C1007 B.n462 VSUBS 0.007662f
C1008 B.n463 VSUBS 0.007662f
C1009 B.n464 VSUBS 0.006197f
C1010 B.n465 VSUBS 0.007662f
C1011 B.n466 VSUBS 0.007662f
C1012 B.n467 VSUBS 0.005296f
C1013 B.n468 VSUBS 0.007662f
C1014 B.n469 VSUBS 0.007662f
C1015 B.n470 VSUBS 0.007662f
C1016 B.n471 VSUBS 0.007662f
C1017 B.n472 VSUBS 0.007662f
C1018 B.n473 VSUBS 0.007662f
C1019 B.n474 VSUBS 0.007662f
C1020 B.n475 VSUBS 0.007662f
C1021 B.n476 VSUBS 0.007662f
C1022 B.n477 VSUBS 0.007662f
C1023 B.n478 VSUBS 0.007662f
C1024 B.n479 VSUBS 0.007662f
C1025 B.n480 VSUBS 0.007662f
C1026 B.n481 VSUBS 0.007662f
C1027 B.n482 VSUBS 0.007662f
C1028 B.n483 VSUBS 0.007662f
C1029 B.n484 VSUBS 0.007662f
C1030 B.n485 VSUBS 0.007662f
C1031 B.n486 VSUBS 0.007662f
C1032 B.n487 VSUBS 0.007662f
C1033 B.n488 VSUBS 0.007662f
C1034 B.n489 VSUBS 0.007662f
C1035 B.n490 VSUBS 0.007662f
C1036 B.n491 VSUBS 0.007662f
C1037 B.n492 VSUBS 0.007662f
C1038 B.n493 VSUBS 0.007662f
C1039 B.n494 VSUBS 0.007662f
C1040 B.n495 VSUBS 0.007662f
C1041 B.n496 VSUBS 0.007662f
C1042 B.n497 VSUBS 0.007662f
C1043 B.n498 VSUBS 0.007662f
C1044 B.n499 VSUBS 0.007662f
C1045 B.n500 VSUBS 0.007662f
C1046 B.n501 VSUBS 0.007662f
C1047 B.n502 VSUBS 0.007662f
C1048 B.n503 VSUBS 0.007662f
C1049 B.n504 VSUBS 0.007662f
C1050 B.n505 VSUBS 0.007662f
C1051 B.n506 VSUBS 0.007662f
C1052 B.n507 VSUBS 0.007662f
C1053 B.n508 VSUBS 0.007662f
C1054 B.n509 VSUBS 0.007662f
C1055 B.n510 VSUBS 0.018845f
C1056 B.n511 VSUBS 0.017436f
C1057 B.n512 VSUBS 0.017436f
C1058 B.n513 VSUBS 0.007662f
C1059 B.n514 VSUBS 0.007662f
C1060 B.n515 VSUBS 0.007662f
C1061 B.n516 VSUBS 0.007662f
C1062 B.n517 VSUBS 0.007662f
C1063 B.n518 VSUBS 0.007662f
C1064 B.n519 VSUBS 0.007662f
C1065 B.n520 VSUBS 0.007662f
C1066 B.n521 VSUBS 0.007662f
C1067 B.n522 VSUBS 0.007662f
C1068 B.n523 VSUBS 0.007662f
C1069 B.n524 VSUBS 0.007662f
C1070 B.n525 VSUBS 0.007662f
C1071 B.n526 VSUBS 0.007662f
C1072 B.n527 VSUBS 0.007662f
C1073 B.n528 VSUBS 0.007662f
C1074 B.n529 VSUBS 0.007662f
C1075 B.n530 VSUBS 0.007662f
C1076 B.n531 VSUBS 0.007662f
C1077 B.n532 VSUBS 0.007662f
C1078 B.n533 VSUBS 0.007662f
C1079 B.n534 VSUBS 0.007662f
C1080 B.n535 VSUBS 0.007662f
C1081 B.n536 VSUBS 0.007662f
C1082 B.n537 VSUBS 0.007662f
C1083 B.n538 VSUBS 0.007662f
C1084 B.n539 VSUBS 0.007662f
C1085 B.n540 VSUBS 0.007662f
C1086 B.n541 VSUBS 0.007662f
C1087 B.n542 VSUBS 0.007662f
C1088 B.n543 VSUBS 0.007662f
C1089 B.n544 VSUBS 0.007662f
C1090 B.n545 VSUBS 0.007662f
C1091 B.n546 VSUBS 0.007662f
C1092 B.n547 VSUBS 0.007662f
C1093 B.n548 VSUBS 0.007662f
C1094 B.n549 VSUBS 0.007662f
C1095 B.n550 VSUBS 0.007662f
C1096 B.n551 VSUBS 0.007662f
C1097 B.n552 VSUBS 0.007662f
C1098 B.n553 VSUBS 0.007662f
C1099 B.n554 VSUBS 0.007662f
C1100 B.n555 VSUBS 0.007662f
C1101 B.n556 VSUBS 0.007662f
C1102 B.n557 VSUBS 0.007662f
C1103 B.n558 VSUBS 0.007662f
C1104 B.n559 VSUBS 0.007662f
C1105 B.n560 VSUBS 0.007662f
C1106 B.n561 VSUBS 0.007662f
C1107 B.n562 VSUBS 0.007662f
C1108 B.n563 VSUBS 0.017349f
.ends

