* NGSPICE file created from diff_pair_sample_1662.ext - technology: sky130A

.subckt diff_pair_sample_1662 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t7 VP.t0 VTAIL.t14 w_n2150_n2704# sky130_fd_pr__pfet_01v8 ad=1.4322 pd=9.01 as=3.3852 ps=18.14 w=8.68 l=0.85
X1 VDD2.t7 VN.t0 VTAIL.t7 w_n2150_n2704# sky130_fd_pr__pfet_01v8 ad=1.4322 pd=9.01 as=1.4322 ps=9.01 w=8.68 l=0.85
X2 B.t11 B.t9 B.t10 w_n2150_n2704# sky130_fd_pr__pfet_01v8 ad=3.3852 pd=18.14 as=0 ps=0 w=8.68 l=0.85
X3 VTAIL.t6 VN.t1 VDD2.t6 w_n2150_n2704# sky130_fd_pr__pfet_01v8 ad=1.4322 pd=9.01 as=1.4322 ps=9.01 w=8.68 l=0.85
X4 VDD2.t5 VN.t2 VTAIL.t5 w_n2150_n2704# sky130_fd_pr__pfet_01v8 ad=1.4322 pd=9.01 as=1.4322 ps=9.01 w=8.68 l=0.85
X5 VTAIL.t4 VN.t3 VDD2.t4 w_n2150_n2704# sky130_fd_pr__pfet_01v8 ad=1.4322 pd=9.01 as=1.4322 ps=9.01 w=8.68 l=0.85
X6 VDD1.t6 VP.t1 VTAIL.t9 w_n2150_n2704# sky130_fd_pr__pfet_01v8 ad=1.4322 pd=9.01 as=1.4322 ps=9.01 w=8.68 l=0.85
X7 B.t8 B.t6 B.t7 w_n2150_n2704# sky130_fd_pr__pfet_01v8 ad=3.3852 pd=18.14 as=0 ps=0 w=8.68 l=0.85
X8 VTAIL.t10 VP.t2 VDD1.t5 w_n2150_n2704# sky130_fd_pr__pfet_01v8 ad=1.4322 pd=9.01 as=1.4322 ps=9.01 w=8.68 l=0.85
X9 VDD2.t3 VN.t4 VTAIL.t0 w_n2150_n2704# sky130_fd_pr__pfet_01v8 ad=1.4322 pd=9.01 as=3.3852 ps=18.14 w=8.68 l=0.85
X10 VTAIL.t12 VP.t3 VDD1.t4 w_n2150_n2704# sky130_fd_pr__pfet_01v8 ad=3.3852 pd=18.14 as=1.4322 ps=9.01 w=8.68 l=0.85
X11 VDD1.t3 VP.t4 VTAIL.t11 w_n2150_n2704# sky130_fd_pr__pfet_01v8 ad=1.4322 pd=9.01 as=1.4322 ps=9.01 w=8.68 l=0.85
X12 VTAIL.t1 VN.t5 VDD2.t2 w_n2150_n2704# sky130_fd_pr__pfet_01v8 ad=3.3852 pd=18.14 as=1.4322 ps=9.01 w=8.68 l=0.85
X13 VTAIL.t15 VP.t5 VDD1.t2 w_n2150_n2704# sky130_fd_pr__pfet_01v8 ad=3.3852 pd=18.14 as=1.4322 ps=9.01 w=8.68 l=0.85
X14 VDD1.t1 VP.t6 VTAIL.t13 w_n2150_n2704# sky130_fd_pr__pfet_01v8 ad=1.4322 pd=9.01 as=3.3852 ps=18.14 w=8.68 l=0.85
X15 B.t5 B.t3 B.t4 w_n2150_n2704# sky130_fd_pr__pfet_01v8 ad=3.3852 pd=18.14 as=0 ps=0 w=8.68 l=0.85
X16 VDD2.t1 VN.t6 VTAIL.t2 w_n2150_n2704# sky130_fd_pr__pfet_01v8 ad=1.4322 pd=9.01 as=3.3852 ps=18.14 w=8.68 l=0.85
X17 VTAIL.t3 VN.t7 VDD2.t0 w_n2150_n2704# sky130_fd_pr__pfet_01v8 ad=3.3852 pd=18.14 as=1.4322 ps=9.01 w=8.68 l=0.85
X18 VTAIL.t8 VP.t7 VDD1.t0 w_n2150_n2704# sky130_fd_pr__pfet_01v8 ad=1.4322 pd=9.01 as=1.4322 ps=9.01 w=8.68 l=0.85
X19 B.t2 B.t0 B.t1 w_n2150_n2704# sky130_fd_pr__pfet_01v8 ad=3.3852 pd=18.14 as=0 ps=0 w=8.68 l=0.85
R0 VP.n7 VP.t3 313.279
R1 VP.n17 VP.t5 292.32
R2 VP.n29 VP.t0 292.32
R3 VP.n15 VP.t6 292.32
R4 VP.n22 VP.t4 246.105
R5 VP.n1 VP.t2 246.105
R6 VP.n5 VP.t7 246.105
R7 VP.n8 VP.t1 246.105
R8 VP.n30 VP.n29 161.3
R9 VP.n9 VP.n6 161.3
R10 VP.n11 VP.n10 161.3
R11 VP.n13 VP.n12 161.3
R12 VP.n14 VP.n4 161.3
R13 VP.n16 VP.n15 161.3
R14 VP.n28 VP.n0 161.3
R15 VP.n27 VP.n26 161.3
R16 VP.n25 VP.n24 161.3
R17 VP.n23 VP.n2 161.3
R18 VP.n21 VP.n20 161.3
R19 VP.n19 VP.n3 161.3
R20 VP.n18 VP.n17 161.3
R21 VP.n24 VP.n23 56.5617
R22 VP.n10 VP.n9 56.5617
R23 VP.n21 VP.n3 47.3584
R24 VP.n28 VP.n27 47.3584
R25 VP.n14 VP.n13 47.3584
R26 VP.n7 VP.n6 42.9081
R27 VP.n18 VP.n16 40.1975
R28 VP.n8 VP.n7 37.615
R29 VP.n23 VP.n22 16.7229
R30 VP.n24 VP.n1 16.7229
R31 VP.n10 VP.n5 16.7229
R32 VP.n9 VP.n8 16.7229
R33 VP.n17 VP.n3 13.8763
R34 VP.n29 VP.n28 13.8763
R35 VP.n15 VP.n14 13.8763
R36 VP.n22 VP.n21 7.86989
R37 VP.n27 VP.n1 7.86989
R38 VP.n13 VP.n5 7.86989
R39 VP.n11 VP.n6 0.189894
R40 VP.n12 VP.n11 0.189894
R41 VP.n12 VP.n4 0.189894
R42 VP.n16 VP.n4 0.189894
R43 VP.n19 VP.n18 0.189894
R44 VP.n20 VP.n19 0.189894
R45 VP.n20 VP.n2 0.189894
R46 VP.n25 VP.n2 0.189894
R47 VP.n26 VP.n25 0.189894
R48 VP.n26 VP.n0 0.189894
R49 VP.n30 VP.n0 0.189894
R50 VP VP.n30 0.0516364
R51 VTAIL.n370 VTAIL.n330 756.745
R52 VTAIL.n42 VTAIL.n2 756.745
R53 VTAIL.n88 VTAIL.n48 756.745
R54 VTAIL.n136 VTAIL.n96 756.745
R55 VTAIL.n324 VTAIL.n284 756.745
R56 VTAIL.n276 VTAIL.n236 756.745
R57 VTAIL.n230 VTAIL.n190 756.745
R58 VTAIL.n182 VTAIL.n142 756.745
R59 VTAIL.n345 VTAIL.n344 585
R60 VTAIL.n342 VTAIL.n341 585
R61 VTAIL.n351 VTAIL.n350 585
R62 VTAIL.n353 VTAIL.n352 585
R63 VTAIL.n338 VTAIL.n337 585
R64 VTAIL.n359 VTAIL.n358 585
R65 VTAIL.n362 VTAIL.n361 585
R66 VTAIL.n360 VTAIL.n334 585
R67 VTAIL.n367 VTAIL.n333 585
R68 VTAIL.n369 VTAIL.n368 585
R69 VTAIL.n371 VTAIL.n370 585
R70 VTAIL.n17 VTAIL.n16 585
R71 VTAIL.n14 VTAIL.n13 585
R72 VTAIL.n23 VTAIL.n22 585
R73 VTAIL.n25 VTAIL.n24 585
R74 VTAIL.n10 VTAIL.n9 585
R75 VTAIL.n31 VTAIL.n30 585
R76 VTAIL.n34 VTAIL.n33 585
R77 VTAIL.n32 VTAIL.n6 585
R78 VTAIL.n39 VTAIL.n5 585
R79 VTAIL.n41 VTAIL.n40 585
R80 VTAIL.n43 VTAIL.n42 585
R81 VTAIL.n63 VTAIL.n62 585
R82 VTAIL.n60 VTAIL.n59 585
R83 VTAIL.n69 VTAIL.n68 585
R84 VTAIL.n71 VTAIL.n70 585
R85 VTAIL.n56 VTAIL.n55 585
R86 VTAIL.n77 VTAIL.n76 585
R87 VTAIL.n80 VTAIL.n79 585
R88 VTAIL.n78 VTAIL.n52 585
R89 VTAIL.n85 VTAIL.n51 585
R90 VTAIL.n87 VTAIL.n86 585
R91 VTAIL.n89 VTAIL.n88 585
R92 VTAIL.n111 VTAIL.n110 585
R93 VTAIL.n108 VTAIL.n107 585
R94 VTAIL.n117 VTAIL.n116 585
R95 VTAIL.n119 VTAIL.n118 585
R96 VTAIL.n104 VTAIL.n103 585
R97 VTAIL.n125 VTAIL.n124 585
R98 VTAIL.n128 VTAIL.n127 585
R99 VTAIL.n126 VTAIL.n100 585
R100 VTAIL.n133 VTAIL.n99 585
R101 VTAIL.n135 VTAIL.n134 585
R102 VTAIL.n137 VTAIL.n136 585
R103 VTAIL.n325 VTAIL.n324 585
R104 VTAIL.n323 VTAIL.n322 585
R105 VTAIL.n321 VTAIL.n287 585
R106 VTAIL.n291 VTAIL.n288 585
R107 VTAIL.n316 VTAIL.n315 585
R108 VTAIL.n314 VTAIL.n313 585
R109 VTAIL.n293 VTAIL.n292 585
R110 VTAIL.n308 VTAIL.n307 585
R111 VTAIL.n306 VTAIL.n305 585
R112 VTAIL.n297 VTAIL.n296 585
R113 VTAIL.n300 VTAIL.n299 585
R114 VTAIL.n277 VTAIL.n276 585
R115 VTAIL.n275 VTAIL.n274 585
R116 VTAIL.n273 VTAIL.n239 585
R117 VTAIL.n243 VTAIL.n240 585
R118 VTAIL.n268 VTAIL.n267 585
R119 VTAIL.n266 VTAIL.n265 585
R120 VTAIL.n245 VTAIL.n244 585
R121 VTAIL.n260 VTAIL.n259 585
R122 VTAIL.n258 VTAIL.n257 585
R123 VTAIL.n249 VTAIL.n248 585
R124 VTAIL.n252 VTAIL.n251 585
R125 VTAIL.n231 VTAIL.n230 585
R126 VTAIL.n229 VTAIL.n228 585
R127 VTAIL.n227 VTAIL.n193 585
R128 VTAIL.n197 VTAIL.n194 585
R129 VTAIL.n222 VTAIL.n221 585
R130 VTAIL.n220 VTAIL.n219 585
R131 VTAIL.n199 VTAIL.n198 585
R132 VTAIL.n214 VTAIL.n213 585
R133 VTAIL.n212 VTAIL.n211 585
R134 VTAIL.n203 VTAIL.n202 585
R135 VTAIL.n206 VTAIL.n205 585
R136 VTAIL.n183 VTAIL.n182 585
R137 VTAIL.n181 VTAIL.n180 585
R138 VTAIL.n179 VTAIL.n145 585
R139 VTAIL.n149 VTAIL.n146 585
R140 VTAIL.n174 VTAIL.n173 585
R141 VTAIL.n172 VTAIL.n171 585
R142 VTAIL.n151 VTAIL.n150 585
R143 VTAIL.n166 VTAIL.n165 585
R144 VTAIL.n164 VTAIL.n163 585
R145 VTAIL.n155 VTAIL.n154 585
R146 VTAIL.n158 VTAIL.n157 585
R147 VTAIL.t13 VTAIL.n298 329.039
R148 VTAIL.t12 VTAIL.n250 329.039
R149 VTAIL.t0 VTAIL.n204 329.039
R150 VTAIL.t1 VTAIL.n156 329.039
R151 VTAIL.t2 VTAIL.n343 329.038
R152 VTAIL.t3 VTAIL.n15 329.038
R153 VTAIL.t14 VTAIL.n61 329.038
R154 VTAIL.t15 VTAIL.n109 329.038
R155 VTAIL.n344 VTAIL.n341 171.744
R156 VTAIL.n351 VTAIL.n341 171.744
R157 VTAIL.n352 VTAIL.n351 171.744
R158 VTAIL.n352 VTAIL.n337 171.744
R159 VTAIL.n359 VTAIL.n337 171.744
R160 VTAIL.n361 VTAIL.n359 171.744
R161 VTAIL.n361 VTAIL.n360 171.744
R162 VTAIL.n360 VTAIL.n333 171.744
R163 VTAIL.n369 VTAIL.n333 171.744
R164 VTAIL.n370 VTAIL.n369 171.744
R165 VTAIL.n16 VTAIL.n13 171.744
R166 VTAIL.n23 VTAIL.n13 171.744
R167 VTAIL.n24 VTAIL.n23 171.744
R168 VTAIL.n24 VTAIL.n9 171.744
R169 VTAIL.n31 VTAIL.n9 171.744
R170 VTAIL.n33 VTAIL.n31 171.744
R171 VTAIL.n33 VTAIL.n32 171.744
R172 VTAIL.n32 VTAIL.n5 171.744
R173 VTAIL.n41 VTAIL.n5 171.744
R174 VTAIL.n42 VTAIL.n41 171.744
R175 VTAIL.n62 VTAIL.n59 171.744
R176 VTAIL.n69 VTAIL.n59 171.744
R177 VTAIL.n70 VTAIL.n69 171.744
R178 VTAIL.n70 VTAIL.n55 171.744
R179 VTAIL.n77 VTAIL.n55 171.744
R180 VTAIL.n79 VTAIL.n77 171.744
R181 VTAIL.n79 VTAIL.n78 171.744
R182 VTAIL.n78 VTAIL.n51 171.744
R183 VTAIL.n87 VTAIL.n51 171.744
R184 VTAIL.n88 VTAIL.n87 171.744
R185 VTAIL.n110 VTAIL.n107 171.744
R186 VTAIL.n117 VTAIL.n107 171.744
R187 VTAIL.n118 VTAIL.n117 171.744
R188 VTAIL.n118 VTAIL.n103 171.744
R189 VTAIL.n125 VTAIL.n103 171.744
R190 VTAIL.n127 VTAIL.n125 171.744
R191 VTAIL.n127 VTAIL.n126 171.744
R192 VTAIL.n126 VTAIL.n99 171.744
R193 VTAIL.n135 VTAIL.n99 171.744
R194 VTAIL.n136 VTAIL.n135 171.744
R195 VTAIL.n324 VTAIL.n323 171.744
R196 VTAIL.n323 VTAIL.n287 171.744
R197 VTAIL.n291 VTAIL.n287 171.744
R198 VTAIL.n315 VTAIL.n291 171.744
R199 VTAIL.n315 VTAIL.n314 171.744
R200 VTAIL.n314 VTAIL.n292 171.744
R201 VTAIL.n307 VTAIL.n292 171.744
R202 VTAIL.n307 VTAIL.n306 171.744
R203 VTAIL.n306 VTAIL.n296 171.744
R204 VTAIL.n299 VTAIL.n296 171.744
R205 VTAIL.n276 VTAIL.n275 171.744
R206 VTAIL.n275 VTAIL.n239 171.744
R207 VTAIL.n243 VTAIL.n239 171.744
R208 VTAIL.n267 VTAIL.n243 171.744
R209 VTAIL.n267 VTAIL.n266 171.744
R210 VTAIL.n266 VTAIL.n244 171.744
R211 VTAIL.n259 VTAIL.n244 171.744
R212 VTAIL.n259 VTAIL.n258 171.744
R213 VTAIL.n258 VTAIL.n248 171.744
R214 VTAIL.n251 VTAIL.n248 171.744
R215 VTAIL.n230 VTAIL.n229 171.744
R216 VTAIL.n229 VTAIL.n193 171.744
R217 VTAIL.n197 VTAIL.n193 171.744
R218 VTAIL.n221 VTAIL.n197 171.744
R219 VTAIL.n221 VTAIL.n220 171.744
R220 VTAIL.n220 VTAIL.n198 171.744
R221 VTAIL.n213 VTAIL.n198 171.744
R222 VTAIL.n213 VTAIL.n212 171.744
R223 VTAIL.n212 VTAIL.n202 171.744
R224 VTAIL.n205 VTAIL.n202 171.744
R225 VTAIL.n182 VTAIL.n181 171.744
R226 VTAIL.n181 VTAIL.n145 171.744
R227 VTAIL.n149 VTAIL.n145 171.744
R228 VTAIL.n173 VTAIL.n149 171.744
R229 VTAIL.n173 VTAIL.n172 171.744
R230 VTAIL.n172 VTAIL.n150 171.744
R231 VTAIL.n165 VTAIL.n150 171.744
R232 VTAIL.n165 VTAIL.n164 171.744
R233 VTAIL.n164 VTAIL.n154 171.744
R234 VTAIL.n157 VTAIL.n154 171.744
R235 VTAIL.n344 VTAIL.t2 85.8723
R236 VTAIL.n16 VTAIL.t3 85.8723
R237 VTAIL.n62 VTAIL.t14 85.8723
R238 VTAIL.n110 VTAIL.t15 85.8723
R239 VTAIL.n299 VTAIL.t13 85.8723
R240 VTAIL.n251 VTAIL.t12 85.8723
R241 VTAIL.n205 VTAIL.t0 85.8723
R242 VTAIL.n157 VTAIL.t1 85.8723
R243 VTAIL.n283 VTAIL.n282 66.7285
R244 VTAIL.n189 VTAIL.n188 66.7285
R245 VTAIL.n1 VTAIL.n0 66.7283
R246 VTAIL.n95 VTAIL.n94 66.7283
R247 VTAIL.n375 VTAIL.n374 35.2884
R248 VTAIL.n47 VTAIL.n46 35.2884
R249 VTAIL.n93 VTAIL.n92 35.2884
R250 VTAIL.n141 VTAIL.n140 35.2884
R251 VTAIL.n329 VTAIL.n328 35.2884
R252 VTAIL.n281 VTAIL.n280 35.2884
R253 VTAIL.n235 VTAIL.n234 35.2884
R254 VTAIL.n187 VTAIL.n186 35.2884
R255 VTAIL.n375 VTAIL.n329 20.8669
R256 VTAIL.n187 VTAIL.n141 20.8669
R257 VTAIL.n368 VTAIL.n367 13.1884
R258 VTAIL.n40 VTAIL.n39 13.1884
R259 VTAIL.n86 VTAIL.n85 13.1884
R260 VTAIL.n134 VTAIL.n133 13.1884
R261 VTAIL.n322 VTAIL.n321 13.1884
R262 VTAIL.n274 VTAIL.n273 13.1884
R263 VTAIL.n228 VTAIL.n227 13.1884
R264 VTAIL.n180 VTAIL.n179 13.1884
R265 VTAIL.n366 VTAIL.n334 12.8005
R266 VTAIL.n371 VTAIL.n332 12.8005
R267 VTAIL.n38 VTAIL.n6 12.8005
R268 VTAIL.n43 VTAIL.n4 12.8005
R269 VTAIL.n84 VTAIL.n52 12.8005
R270 VTAIL.n89 VTAIL.n50 12.8005
R271 VTAIL.n132 VTAIL.n100 12.8005
R272 VTAIL.n137 VTAIL.n98 12.8005
R273 VTAIL.n325 VTAIL.n286 12.8005
R274 VTAIL.n320 VTAIL.n288 12.8005
R275 VTAIL.n277 VTAIL.n238 12.8005
R276 VTAIL.n272 VTAIL.n240 12.8005
R277 VTAIL.n231 VTAIL.n192 12.8005
R278 VTAIL.n226 VTAIL.n194 12.8005
R279 VTAIL.n183 VTAIL.n144 12.8005
R280 VTAIL.n178 VTAIL.n146 12.8005
R281 VTAIL.n363 VTAIL.n362 12.0247
R282 VTAIL.n372 VTAIL.n330 12.0247
R283 VTAIL.n35 VTAIL.n34 12.0247
R284 VTAIL.n44 VTAIL.n2 12.0247
R285 VTAIL.n81 VTAIL.n80 12.0247
R286 VTAIL.n90 VTAIL.n48 12.0247
R287 VTAIL.n129 VTAIL.n128 12.0247
R288 VTAIL.n138 VTAIL.n96 12.0247
R289 VTAIL.n326 VTAIL.n284 12.0247
R290 VTAIL.n317 VTAIL.n316 12.0247
R291 VTAIL.n278 VTAIL.n236 12.0247
R292 VTAIL.n269 VTAIL.n268 12.0247
R293 VTAIL.n232 VTAIL.n190 12.0247
R294 VTAIL.n223 VTAIL.n222 12.0247
R295 VTAIL.n184 VTAIL.n142 12.0247
R296 VTAIL.n175 VTAIL.n174 12.0247
R297 VTAIL.n358 VTAIL.n336 11.249
R298 VTAIL.n30 VTAIL.n8 11.249
R299 VTAIL.n76 VTAIL.n54 11.249
R300 VTAIL.n124 VTAIL.n102 11.249
R301 VTAIL.n313 VTAIL.n290 11.249
R302 VTAIL.n265 VTAIL.n242 11.249
R303 VTAIL.n219 VTAIL.n196 11.249
R304 VTAIL.n171 VTAIL.n148 11.249
R305 VTAIL.n345 VTAIL.n343 10.7239
R306 VTAIL.n17 VTAIL.n15 10.7239
R307 VTAIL.n63 VTAIL.n61 10.7239
R308 VTAIL.n111 VTAIL.n109 10.7239
R309 VTAIL.n300 VTAIL.n298 10.7239
R310 VTAIL.n252 VTAIL.n250 10.7239
R311 VTAIL.n206 VTAIL.n204 10.7239
R312 VTAIL.n158 VTAIL.n156 10.7239
R313 VTAIL.n357 VTAIL.n338 10.4732
R314 VTAIL.n29 VTAIL.n10 10.4732
R315 VTAIL.n75 VTAIL.n56 10.4732
R316 VTAIL.n123 VTAIL.n104 10.4732
R317 VTAIL.n312 VTAIL.n293 10.4732
R318 VTAIL.n264 VTAIL.n245 10.4732
R319 VTAIL.n218 VTAIL.n199 10.4732
R320 VTAIL.n170 VTAIL.n151 10.4732
R321 VTAIL.n354 VTAIL.n353 9.69747
R322 VTAIL.n26 VTAIL.n25 9.69747
R323 VTAIL.n72 VTAIL.n71 9.69747
R324 VTAIL.n120 VTAIL.n119 9.69747
R325 VTAIL.n309 VTAIL.n308 9.69747
R326 VTAIL.n261 VTAIL.n260 9.69747
R327 VTAIL.n215 VTAIL.n214 9.69747
R328 VTAIL.n167 VTAIL.n166 9.69747
R329 VTAIL.n374 VTAIL.n373 9.45567
R330 VTAIL.n46 VTAIL.n45 9.45567
R331 VTAIL.n92 VTAIL.n91 9.45567
R332 VTAIL.n140 VTAIL.n139 9.45567
R333 VTAIL.n328 VTAIL.n327 9.45567
R334 VTAIL.n280 VTAIL.n279 9.45567
R335 VTAIL.n234 VTAIL.n233 9.45567
R336 VTAIL.n186 VTAIL.n185 9.45567
R337 VTAIL.n373 VTAIL.n372 9.3005
R338 VTAIL.n332 VTAIL.n331 9.3005
R339 VTAIL.n347 VTAIL.n346 9.3005
R340 VTAIL.n349 VTAIL.n348 9.3005
R341 VTAIL.n340 VTAIL.n339 9.3005
R342 VTAIL.n355 VTAIL.n354 9.3005
R343 VTAIL.n357 VTAIL.n356 9.3005
R344 VTAIL.n336 VTAIL.n335 9.3005
R345 VTAIL.n364 VTAIL.n363 9.3005
R346 VTAIL.n366 VTAIL.n365 9.3005
R347 VTAIL.n45 VTAIL.n44 9.3005
R348 VTAIL.n4 VTAIL.n3 9.3005
R349 VTAIL.n19 VTAIL.n18 9.3005
R350 VTAIL.n21 VTAIL.n20 9.3005
R351 VTAIL.n12 VTAIL.n11 9.3005
R352 VTAIL.n27 VTAIL.n26 9.3005
R353 VTAIL.n29 VTAIL.n28 9.3005
R354 VTAIL.n8 VTAIL.n7 9.3005
R355 VTAIL.n36 VTAIL.n35 9.3005
R356 VTAIL.n38 VTAIL.n37 9.3005
R357 VTAIL.n91 VTAIL.n90 9.3005
R358 VTAIL.n50 VTAIL.n49 9.3005
R359 VTAIL.n65 VTAIL.n64 9.3005
R360 VTAIL.n67 VTAIL.n66 9.3005
R361 VTAIL.n58 VTAIL.n57 9.3005
R362 VTAIL.n73 VTAIL.n72 9.3005
R363 VTAIL.n75 VTAIL.n74 9.3005
R364 VTAIL.n54 VTAIL.n53 9.3005
R365 VTAIL.n82 VTAIL.n81 9.3005
R366 VTAIL.n84 VTAIL.n83 9.3005
R367 VTAIL.n139 VTAIL.n138 9.3005
R368 VTAIL.n98 VTAIL.n97 9.3005
R369 VTAIL.n113 VTAIL.n112 9.3005
R370 VTAIL.n115 VTAIL.n114 9.3005
R371 VTAIL.n106 VTAIL.n105 9.3005
R372 VTAIL.n121 VTAIL.n120 9.3005
R373 VTAIL.n123 VTAIL.n122 9.3005
R374 VTAIL.n102 VTAIL.n101 9.3005
R375 VTAIL.n130 VTAIL.n129 9.3005
R376 VTAIL.n132 VTAIL.n131 9.3005
R377 VTAIL.n302 VTAIL.n301 9.3005
R378 VTAIL.n304 VTAIL.n303 9.3005
R379 VTAIL.n295 VTAIL.n294 9.3005
R380 VTAIL.n310 VTAIL.n309 9.3005
R381 VTAIL.n312 VTAIL.n311 9.3005
R382 VTAIL.n290 VTAIL.n289 9.3005
R383 VTAIL.n318 VTAIL.n317 9.3005
R384 VTAIL.n320 VTAIL.n319 9.3005
R385 VTAIL.n327 VTAIL.n326 9.3005
R386 VTAIL.n286 VTAIL.n285 9.3005
R387 VTAIL.n254 VTAIL.n253 9.3005
R388 VTAIL.n256 VTAIL.n255 9.3005
R389 VTAIL.n247 VTAIL.n246 9.3005
R390 VTAIL.n262 VTAIL.n261 9.3005
R391 VTAIL.n264 VTAIL.n263 9.3005
R392 VTAIL.n242 VTAIL.n241 9.3005
R393 VTAIL.n270 VTAIL.n269 9.3005
R394 VTAIL.n272 VTAIL.n271 9.3005
R395 VTAIL.n279 VTAIL.n278 9.3005
R396 VTAIL.n238 VTAIL.n237 9.3005
R397 VTAIL.n208 VTAIL.n207 9.3005
R398 VTAIL.n210 VTAIL.n209 9.3005
R399 VTAIL.n201 VTAIL.n200 9.3005
R400 VTAIL.n216 VTAIL.n215 9.3005
R401 VTAIL.n218 VTAIL.n217 9.3005
R402 VTAIL.n196 VTAIL.n195 9.3005
R403 VTAIL.n224 VTAIL.n223 9.3005
R404 VTAIL.n226 VTAIL.n225 9.3005
R405 VTAIL.n233 VTAIL.n232 9.3005
R406 VTAIL.n192 VTAIL.n191 9.3005
R407 VTAIL.n160 VTAIL.n159 9.3005
R408 VTAIL.n162 VTAIL.n161 9.3005
R409 VTAIL.n153 VTAIL.n152 9.3005
R410 VTAIL.n168 VTAIL.n167 9.3005
R411 VTAIL.n170 VTAIL.n169 9.3005
R412 VTAIL.n148 VTAIL.n147 9.3005
R413 VTAIL.n176 VTAIL.n175 9.3005
R414 VTAIL.n178 VTAIL.n177 9.3005
R415 VTAIL.n185 VTAIL.n184 9.3005
R416 VTAIL.n144 VTAIL.n143 9.3005
R417 VTAIL.n350 VTAIL.n340 8.92171
R418 VTAIL.n22 VTAIL.n12 8.92171
R419 VTAIL.n68 VTAIL.n58 8.92171
R420 VTAIL.n116 VTAIL.n106 8.92171
R421 VTAIL.n305 VTAIL.n295 8.92171
R422 VTAIL.n257 VTAIL.n247 8.92171
R423 VTAIL.n211 VTAIL.n201 8.92171
R424 VTAIL.n163 VTAIL.n153 8.92171
R425 VTAIL.n349 VTAIL.n342 8.14595
R426 VTAIL.n21 VTAIL.n14 8.14595
R427 VTAIL.n67 VTAIL.n60 8.14595
R428 VTAIL.n115 VTAIL.n108 8.14595
R429 VTAIL.n304 VTAIL.n297 8.14595
R430 VTAIL.n256 VTAIL.n249 8.14595
R431 VTAIL.n210 VTAIL.n203 8.14595
R432 VTAIL.n162 VTAIL.n155 8.14595
R433 VTAIL.n346 VTAIL.n345 7.3702
R434 VTAIL.n18 VTAIL.n17 7.3702
R435 VTAIL.n64 VTAIL.n63 7.3702
R436 VTAIL.n112 VTAIL.n111 7.3702
R437 VTAIL.n301 VTAIL.n300 7.3702
R438 VTAIL.n253 VTAIL.n252 7.3702
R439 VTAIL.n207 VTAIL.n206 7.3702
R440 VTAIL.n159 VTAIL.n158 7.3702
R441 VTAIL.n346 VTAIL.n342 5.81868
R442 VTAIL.n18 VTAIL.n14 5.81868
R443 VTAIL.n64 VTAIL.n60 5.81868
R444 VTAIL.n112 VTAIL.n108 5.81868
R445 VTAIL.n301 VTAIL.n297 5.81868
R446 VTAIL.n253 VTAIL.n249 5.81868
R447 VTAIL.n207 VTAIL.n203 5.81868
R448 VTAIL.n159 VTAIL.n155 5.81868
R449 VTAIL.n350 VTAIL.n349 5.04292
R450 VTAIL.n22 VTAIL.n21 5.04292
R451 VTAIL.n68 VTAIL.n67 5.04292
R452 VTAIL.n116 VTAIL.n115 5.04292
R453 VTAIL.n305 VTAIL.n304 5.04292
R454 VTAIL.n257 VTAIL.n256 5.04292
R455 VTAIL.n211 VTAIL.n210 5.04292
R456 VTAIL.n163 VTAIL.n162 5.04292
R457 VTAIL.n353 VTAIL.n340 4.26717
R458 VTAIL.n25 VTAIL.n12 4.26717
R459 VTAIL.n71 VTAIL.n58 4.26717
R460 VTAIL.n119 VTAIL.n106 4.26717
R461 VTAIL.n308 VTAIL.n295 4.26717
R462 VTAIL.n260 VTAIL.n247 4.26717
R463 VTAIL.n214 VTAIL.n201 4.26717
R464 VTAIL.n166 VTAIL.n153 4.26717
R465 VTAIL.n0 VTAIL.t5 3.74532
R466 VTAIL.n0 VTAIL.t4 3.74532
R467 VTAIL.n94 VTAIL.t11 3.74532
R468 VTAIL.n94 VTAIL.t10 3.74532
R469 VTAIL.n282 VTAIL.t9 3.74532
R470 VTAIL.n282 VTAIL.t8 3.74532
R471 VTAIL.n188 VTAIL.t7 3.74532
R472 VTAIL.n188 VTAIL.t6 3.74532
R473 VTAIL.n354 VTAIL.n338 3.49141
R474 VTAIL.n26 VTAIL.n10 3.49141
R475 VTAIL.n72 VTAIL.n56 3.49141
R476 VTAIL.n120 VTAIL.n104 3.49141
R477 VTAIL.n309 VTAIL.n293 3.49141
R478 VTAIL.n261 VTAIL.n245 3.49141
R479 VTAIL.n215 VTAIL.n199 3.49141
R480 VTAIL.n167 VTAIL.n151 3.49141
R481 VTAIL.n358 VTAIL.n357 2.71565
R482 VTAIL.n30 VTAIL.n29 2.71565
R483 VTAIL.n76 VTAIL.n75 2.71565
R484 VTAIL.n124 VTAIL.n123 2.71565
R485 VTAIL.n313 VTAIL.n312 2.71565
R486 VTAIL.n265 VTAIL.n264 2.71565
R487 VTAIL.n219 VTAIL.n218 2.71565
R488 VTAIL.n171 VTAIL.n170 2.71565
R489 VTAIL.n347 VTAIL.n343 2.41285
R490 VTAIL.n19 VTAIL.n15 2.41285
R491 VTAIL.n65 VTAIL.n61 2.41285
R492 VTAIL.n113 VTAIL.n109 2.41285
R493 VTAIL.n302 VTAIL.n298 2.41285
R494 VTAIL.n254 VTAIL.n250 2.41285
R495 VTAIL.n208 VTAIL.n204 2.41285
R496 VTAIL.n160 VTAIL.n156 2.41285
R497 VTAIL.n362 VTAIL.n336 1.93989
R498 VTAIL.n374 VTAIL.n330 1.93989
R499 VTAIL.n34 VTAIL.n8 1.93989
R500 VTAIL.n46 VTAIL.n2 1.93989
R501 VTAIL.n80 VTAIL.n54 1.93989
R502 VTAIL.n92 VTAIL.n48 1.93989
R503 VTAIL.n128 VTAIL.n102 1.93989
R504 VTAIL.n140 VTAIL.n96 1.93989
R505 VTAIL.n328 VTAIL.n284 1.93989
R506 VTAIL.n316 VTAIL.n290 1.93989
R507 VTAIL.n280 VTAIL.n236 1.93989
R508 VTAIL.n268 VTAIL.n242 1.93989
R509 VTAIL.n234 VTAIL.n190 1.93989
R510 VTAIL.n222 VTAIL.n196 1.93989
R511 VTAIL.n186 VTAIL.n142 1.93989
R512 VTAIL.n174 VTAIL.n148 1.93989
R513 VTAIL.n363 VTAIL.n334 1.16414
R514 VTAIL.n372 VTAIL.n371 1.16414
R515 VTAIL.n35 VTAIL.n6 1.16414
R516 VTAIL.n44 VTAIL.n43 1.16414
R517 VTAIL.n81 VTAIL.n52 1.16414
R518 VTAIL.n90 VTAIL.n89 1.16414
R519 VTAIL.n129 VTAIL.n100 1.16414
R520 VTAIL.n138 VTAIL.n137 1.16414
R521 VTAIL.n326 VTAIL.n325 1.16414
R522 VTAIL.n317 VTAIL.n288 1.16414
R523 VTAIL.n278 VTAIL.n277 1.16414
R524 VTAIL.n269 VTAIL.n240 1.16414
R525 VTAIL.n232 VTAIL.n231 1.16414
R526 VTAIL.n223 VTAIL.n194 1.16414
R527 VTAIL.n184 VTAIL.n183 1.16414
R528 VTAIL.n175 VTAIL.n146 1.16414
R529 VTAIL.n189 VTAIL.n187 1.01774
R530 VTAIL.n235 VTAIL.n189 1.01774
R531 VTAIL.n283 VTAIL.n281 1.01774
R532 VTAIL.n329 VTAIL.n283 1.01774
R533 VTAIL.n141 VTAIL.n95 1.01774
R534 VTAIL.n95 VTAIL.n93 1.01774
R535 VTAIL.n47 VTAIL.n1 1.01774
R536 VTAIL VTAIL.n375 0.959552
R537 VTAIL.n281 VTAIL.n235 0.470328
R538 VTAIL.n93 VTAIL.n47 0.470328
R539 VTAIL.n367 VTAIL.n366 0.388379
R540 VTAIL.n368 VTAIL.n332 0.388379
R541 VTAIL.n39 VTAIL.n38 0.388379
R542 VTAIL.n40 VTAIL.n4 0.388379
R543 VTAIL.n85 VTAIL.n84 0.388379
R544 VTAIL.n86 VTAIL.n50 0.388379
R545 VTAIL.n133 VTAIL.n132 0.388379
R546 VTAIL.n134 VTAIL.n98 0.388379
R547 VTAIL.n322 VTAIL.n286 0.388379
R548 VTAIL.n321 VTAIL.n320 0.388379
R549 VTAIL.n274 VTAIL.n238 0.388379
R550 VTAIL.n273 VTAIL.n272 0.388379
R551 VTAIL.n228 VTAIL.n192 0.388379
R552 VTAIL.n227 VTAIL.n226 0.388379
R553 VTAIL.n180 VTAIL.n144 0.388379
R554 VTAIL.n179 VTAIL.n178 0.388379
R555 VTAIL.n348 VTAIL.n347 0.155672
R556 VTAIL.n348 VTAIL.n339 0.155672
R557 VTAIL.n355 VTAIL.n339 0.155672
R558 VTAIL.n356 VTAIL.n355 0.155672
R559 VTAIL.n356 VTAIL.n335 0.155672
R560 VTAIL.n364 VTAIL.n335 0.155672
R561 VTAIL.n365 VTAIL.n364 0.155672
R562 VTAIL.n365 VTAIL.n331 0.155672
R563 VTAIL.n373 VTAIL.n331 0.155672
R564 VTAIL.n20 VTAIL.n19 0.155672
R565 VTAIL.n20 VTAIL.n11 0.155672
R566 VTAIL.n27 VTAIL.n11 0.155672
R567 VTAIL.n28 VTAIL.n27 0.155672
R568 VTAIL.n28 VTAIL.n7 0.155672
R569 VTAIL.n36 VTAIL.n7 0.155672
R570 VTAIL.n37 VTAIL.n36 0.155672
R571 VTAIL.n37 VTAIL.n3 0.155672
R572 VTAIL.n45 VTAIL.n3 0.155672
R573 VTAIL.n66 VTAIL.n65 0.155672
R574 VTAIL.n66 VTAIL.n57 0.155672
R575 VTAIL.n73 VTAIL.n57 0.155672
R576 VTAIL.n74 VTAIL.n73 0.155672
R577 VTAIL.n74 VTAIL.n53 0.155672
R578 VTAIL.n82 VTAIL.n53 0.155672
R579 VTAIL.n83 VTAIL.n82 0.155672
R580 VTAIL.n83 VTAIL.n49 0.155672
R581 VTAIL.n91 VTAIL.n49 0.155672
R582 VTAIL.n114 VTAIL.n113 0.155672
R583 VTAIL.n114 VTAIL.n105 0.155672
R584 VTAIL.n121 VTAIL.n105 0.155672
R585 VTAIL.n122 VTAIL.n121 0.155672
R586 VTAIL.n122 VTAIL.n101 0.155672
R587 VTAIL.n130 VTAIL.n101 0.155672
R588 VTAIL.n131 VTAIL.n130 0.155672
R589 VTAIL.n131 VTAIL.n97 0.155672
R590 VTAIL.n139 VTAIL.n97 0.155672
R591 VTAIL.n327 VTAIL.n285 0.155672
R592 VTAIL.n319 VTAIL.n285 0.155672
R593 VTAIL.n319 VTAIL.n318 0.155672
R594 VTAIL.n318 VTAIL.n289 0.155672
R595 VTAIL.n311 VTAIL.n289 0.155672
R596 VTAIL.n311 VTAIL.n310 0.155672
R597 VTAIL.n310 VTAIL.n294 0.155672
R598 VTAIL.n303 VTAIL.n294 0.155672
R599 VTAIL.n303 VTAIL.n302 0.155672
R600 VTAIL.n279 VTAIL.n237 0.155672
R601 VTAIL.n271 VTAIL.n237 0.155672
R602 VTAIL.n271 VTAIL.n270 0.155672
R603 VTAIL.n270 VTAIL.n241 0.155672
R604 VTAIL.n263 VTAIL.n241 0.155672
R605 VTAIL.n263 VTAIL.n262 0.155672
R606 VTAIL.n262 VTAIL.n246 0.155672
R607 VTAIL.n255 VTAIL.n246 0.155672
R608 VTAIL.n255 VTAIL.n254 0.155672
R609 VTAIL.n233 VTAIL.n191 0.155672
R610 VTAIL.n225 VTAIL.n191 0.155672
R611 VTAIL.n225 VTAIL.n224 0.155672
R612 VTAIL.n224 VTAIL.n195 0.155672
R613 VTAIL.n217 VTAIL.n195 0.155672
R614 VTAIL.n217 VTAIL.n216 0.155672
R615 VTAIL.n216 VTAIL.n200 0.155672
R616 VTAIL.n209 VTAIL.n200 0.155672
R617 VTAIL.n209 VTAIL.n208 0.155672
R618 VTAIL.n185 VTAIL.n143 0.155672
R619 VTAIL.n177 VTAIL.n143 0.155672
R620 VTAIL.n177 VTAIL.n176 0.155672
R621 VTAIL.n176 VTAIL.n147 0.155672
R622 VTAIL.n169 VTAIL.n147 0.155672
R623 VTAIL.n169 VTAIL.n168 0.155672
R624 VTAIL.n168 VTAIL.n152 0.155672
R625 VTAIL.n161 VTAIL.n152 0.155672
R626 VTAIL.n161 VTAIL.n160 0.155672
R627 VTAIL VTAIL.n1 0.0586897
R628 VDD1 VDD1.n0 83.9741
R629 VDD1.n3 VDD1.n2 83.8604
R630 VDD1.n3 VDD1.n1 83.8604
R631 VDD1.n5 VDD1.n4 83.4071
R632 VDD1.n5 VDD1.n3 36.3587
R633 VDD1.n4 VDD1.t0 3.74532
R634 VDD1.n4 VDD1.t1 3.74532
R635 VDD1.n0 VDD1.t4 3.74532
R636 VDD1.n0 VDD1.t6 3.74532
R637 VDD1.n2 VDD1.t5 3.74532
R638 VDD1.n2 VDD1.t7 3.74532
R639 VDD1.n1 VDD1.t2 3.74532
R640 VDD1.n1 VDD1.t3 3.74532
R641 VDD1 VDD1.n5 0.450931
R642 VN.n3 VN.t7 313.279
R643 VN.n16 VN.t4 313.279
R644 VN.n11 VN.t6 292.32
R645 VN.n24 VN.t5 292.32
R646 VN.n4 VN.t2 246.105
R647 VN.n1 VN.t3 246.105
R648 VN.n17 VN.t1 246.105
R649 VN.n14 VN.t0 246.105
R650 VN.n12 VN.n11 161.3
R651 VN.n25 VN.n24 161.3
R652 VN.n23 VN.n13 161.3
R653 VN.n22 VN.n21 161.3
R654 VN.n20 VN.n19 161.3
R655 VN.n18 VN.n15 161.3
R656 VN.n10 VN.n0 161.3
R657 VN.n9 VN.n8 161.3
R658 VN.n7 VN.n6 161.3
R659 VN.n5 VN.n2 161.3
R660 VN.n6 VN.n5 56.5617
R661 VN.n19 VN.n18 56.5617
R662 VN.n10 VN.n9 47.3584
R663 VN.n23 VN.n22 47.3584
R664 VN.n16 VN.n15 42.9081
R665 VN.n3 VN.n2 42.9081
R666 VN VN.n25 40.5781
R667 VN.n4 VN.n3 37.615
R668 VN.n17 VN.n16 37.615
R669 VN.n5 VN.n4 16.7229
R670 VN.n6 VN.n1 16.7229
R671 VN.n18 VN.n17 16.7229
R672 VN.n19 VN.n14 16.7229
R673 VN.n11 VN.n10 13.8763
R674 VN.n24 VN.n23 13.8763
R675 VN.n9 VN.n1 7.86989
R676 VN.n22 VN.n14 7.86989
R677 VN.n25 VN.n13 0.189894
R678 VN.n21 VN.n13 0.189894
R679 VN.n21 VN.n20 0.189894
R680 VN.n20 VN.n15 0.189894
R681 VN.n7 VN.n2 0.189894
R682 VN.n8 VN.n7 0.189894
R683 VN.n8 VN.n0 0.189894
R684 VN.n12 VN.n0 0.189894
R685 VN VN.n12 0.0516364
R686 VDD2.n2 VDD2.n1 83.8604
R687 VDD2.n2 VDD2.n0 83.8604
R688 VDD2 VDD2.n5 83.8576
R689 VDD2.n4 VDD2.n3 83.4073
R690 VDD2.n4 VDD2.n2 35.7756
R691 VDD2.n5 VDD2.t6 3.74532
R692 VDD2.n5 VDD2.t3 3.74532
R693 VDD2.n3 VDD2.t2 3.74532
R694 VDD2.n3 VDD2.t7 3.74532
R695 VDD2.n1 VDD2.t4 3.74532
R696 VDD2.n1 VDD2.t1 3.74532
R697 VDD2.n0 VDD2.t0 3.74532
R698 VDD2.n0 VDD2.t5 3.74532
R699 VDD2 VDD2.n4 0.56731
R700 B.n281 B.n82 585
R701 B.n280 B.n279 585
R702 B.n278 B.n83 585
R703 B.n277 B.n276 585
R704 B.n275 B.n84 585
R705 B.n274 B.n273 585
R706 B.n272 B.n85 585
R707 B.n271 B.n270 585
R708 B.n269 B.n86 585
R709 B.n268 B.n267 585
R710 B.n266 B.n87 585
R711 B.n265 B.n264 585
R712 B.n263 B.n88 585
R713 B.n262 B.n261 585
R714 B.n260 B.n89 585
R715 B.n259 B.n258 585
R716 B.n257 B.n90 585
R717 B.n256 B.n255 585
R718 B.n254 B.n91 585
R719 B.n253 B.n252 585
R720 B.n251 B.n92 585
R721 B.n250 B.n249 585
R722 B.n248 B.n93 585
R723 B.n247 B.n246 585
R724 B.n245 B.n94 585
R725 B.n244 B.n243 585
R726 B.n242 B.n95 585
R727 B.n241 B.n240 585
R728 B.n239 B.n96 585
R729 B.n238 B.n237 585
R730 B.n236 B.n97 585
R731 B.n235 B.n234 585
R732 B.n232 B.n98 585
R733 B.n231 B.n230 585
R734 B.n229 B.n101 585
R735 B.n228 B.n227 585
R736 B.n226 B.n102 585
R737 B.n225 B.n224 585
R738 B.n223 B.n103 585
R739 B.n222 B.n221 585
R740 B.n220 B.n104 585
R741 B.n218 B.n217 585
R742 B.n216 B.n107 585
R743 B.n215 B.n214 585
R744 B.n213 B.n108 585
R745 B.n212 B.n211 585
R746 B.n210 B.n109 585
R747 B.n209 B.n208 585
R748 B.n207 B.n110 585
R749 B.n206 B.n205 585
R750 B.n204 B.n111 585
R751 B.n203 B.n202 585
R752 B.n201 B.n112 585
R753 B.n200 B.n199 585
R754 B.n198 B.n113 585
R755 B.n197 B.n196 585
R756 B.n195 B.n114 585
R757 B.n194 B.n193 585
R758 B.n192 B.n115 585
R759 B.n191 B.n190 585
R760 B.n189 B.n116 585
R761 B.n188 B.n187 585
R762 B.n186 B.n117 585
R763 B.n185 B.n184 585
R764 B.n183 B.n118 585
R765 B.n182 B.n181 585
R766 B.n180 B.n119 585
R767 B.n179 B.n178 585
R768 B.n177 B.n120 585
R769 B.n176 B.n175 585
R770 B.n174 B.n121 585
R771 B.n173 B.n172 585
R772 B.n171 B.n122 585
R773 B.n283 B.n282 585
R774 B.n284 B.n81 585
R775 B.n286 B.n285 585
R776 B.n287 B.n80 585
R777 B.n289 B.n288 585
R778 B.n290 B.n79 585
R779 B.n292 B.n291 585
R780 B.n293 B.n78 585
R781 B.n295 B.n294 585
R782 B.n296 B.n77 585
R783 B.n298 B.n297 585
R784 B.n299 B.n76 585
R785 B.n301 B.n300 585
R786 B.n302 B.n75 585
R787 B.n304 B.n303 585
R788 B.n305 B.n74 585
R789 B.n307 B.n306 585
R790 B.n308 B.n73 585
R791 B.n310 B.n309 585
R792 B.n311 B.n72 585
R793 B.n313 B.n312 585
R794 B.n314 B.n71 585
R795 B.n316 B.n315 585
R796 B.n317 B.n70 585
R797 B.n319 B.n318 585
R798 B.n320 B.n69 585
R799 B.n322 B.n321 585
R800 B.n323 B.n68 585
R801 B.n325 B.n324 585
R802 B.n326 B.n67 585
R803 B.n328 B.n327 585
R804 B.n329 B.n66 585
R805 B.n331 B.n330 585
R806 B.n332 B.n65 585
R807 B.n334 B.n333 585
R808 B.n335 B.n64 585
R809 B.n337 B.n336 585
R810 B.n338 B.n63 585
R811 B.n340 B.n339 585
R812 B.n341 B.n62 585
R813 B.n343 B.n342 585
R814 B.n344 B.n61 585
R815 B.n346 B.n345 585
R816 B.n347 B.n60 585
R817 B.n349 B.n348 585
R818 B.n350 B.n59 585
R819 B.n352 B.n351 585
R820 B.n353 B.n58 585
R821 B.n355 B.n354 585
R822 B.n356 B.n57 585
R823 B.n358 B.n357 585
R824 B.n359 B.n56 585
R825 B.n470 B.n469 585
R826 B.n468 B.n15 585
R827 B.n467 B.n466 585
R828 B.n465 B.n16 585
R829 B.n464 B.n463 585
R830 B.n462 B.n17 585
R831 B.n461 B.n460 585
R832 B.n459 B.n18 585
R833 B.n458 B.n457 585
R834 B.n456 B.n19 585
R835 B.n455 B.n454 585
R836 B.n453 B.n20 585
R837 B.n452 B.n451 585
R838 B.n450 B.n21 585
R839 B.n449 B.n448 585
R840 B.n447 B.n22 585
R841 B.n446 B.n445 585
R842 B.n444 B.n23 585
R843 B.n443 B.n442 585
R844 B.n441 B.n24 585
R845 B.n440 B.n439 585
R846 B.n438 B.n25 585
R847 B.n437 B.n436 585
R848 B.n435 B.n26 585
R849 B.n434 B.n433 585
R850 B.n432 B.n27 585
R851 B.n431 B.n430 585
R852 B.n429 B.n28 585
R853 B.n428 B.n427 585
R854 B.n426 B.n29 585
R855 B.n425 B.n424 585
R856 B.n423 B.n30 585
R857 B.n422 B.n421 585
R858 B.n420 B.n31 585
R859 B.n419 B.n418 585
R860 B.n417 B.n35 585
R861 B.n416 B.n415 585
R862 B.n414 B.n36 585
R863 B.n413 B.n412 585
R864 B.n411 B.n37 585
R865 B.n410 B.n409 585
R866 B.n407 B.n38 585
R867 B.n406 B.n405 585
R868 B.n404 B.n41 585
R869 B.n403 B.n402 585
R870 B.n401 B.n42 585
R871 B.n400 B.n399 585
R872 B.n398 B.n43 585
R873 B.n397 B.n396 585
R874 B.n395 B.n44 585
R875 B.n394 B.n393 585
R876 B.n392 B.n45 585
R877 B.n391 B.n390 585
R878 B.n389 B.n46 585
R879 B.n388 B.n387 585
R880 B.n386 B.n47 585
R881 B.n385 B.n384 585
R882 B.n383 B.n48 585
R883 B.n382 B.n381 585
R884 B.n380 B.n49 585
R885 B.n379 B.n378 585
R886 B.n377 B.n50 585
R887 B.n376 B.n375 585
R888 B.n374 B.n51 585
R889 B.n373 B.n372 585
R890 B.n371 B.n52 585
R891 B.n370 B.n369 585
R892 B.n368 B.n53 585
R893 B.n367 B.n366 585
R894 B.n365 B.n54 585
R895 B.n364 B.n363 585
R896 B.n362 B.n55 585
R897 B.n361 B.n360 585
R898 B.n471 B.n14 585
R899 B.n473 B.n472 585
R900 B.n474 B.n13 585
R901 B.n476 B.n475 585
R902 B.n477 B.n12 585
R903 B.n479 B.n478 585
R904 B.n480 B.n11 585
R905 B.n482 B.n481 585
R906 B.n483 B.n10 585
R907 B.n485 B.n484 585
R908 B.n486 B.n9 585
R909 B.n488 B.n487 585
R910 B.n489 B.n8 585
R911 B.n491 B.n490 585
R912 B.n492 B.n7 585
R913 B.n494 B.n493 585
R914 B.n495 B.n6 585
R915 B.n497 B.n496 585
R916 B.n498 B.n5 585
R917 B.n500 B.n499 585
R918 B.n501 B.n4 585
R919 B.n503 B.n502 585
R920 B.n504 B.n3 585
R921 B.n506 B.n505 585
R922 B.n507 B.n0 585
R923 B.n2 B.n1 585
R924 B.n135 B.n134 585
R925 B.n137 B.n136 585
R926 B.n138 B.n133 585
R927 B.n140 B.n139 585
R928 B.n141 B.n132 585
R929 B.n143 B.n142 585
R930 B.n144 B.n131 585
R931 B.n146 B.n145 585
R932 B.n147 B.n130 585
R933 B.n149 B.n148 585
R934 B.n150 B.n129 585
R935 B.n152 B.n151 585
R936 B.n153 B.n128 585
R937 B.n155 B.n154 585
R938 B.n156 B.n127 585
R939 B.n158 B.n157 585
R940 B.n159 B.n126 585
R941 B.n161 B.n160 585
R942 B.n162 B.n125 585
R943 B.n164 B.n163 585
R944 B.n165 B.n124 585
R945 B.n167 B.n166 585
R946 B.n168 B.n123 585
R947 B.n170 B.n169 585
R948 B.n169 B.n122 516.524
R949 B.n283 B.n82 516.524
R950 B.n361 B.n56 516.524
R951 B.n471 B.n470 516.524
R952 B.n105 B.t0 447.892
R953 B.n99 B.t3 447.892
R954 B.n39 B.t9 447.892
R955 B.n32 B.t6 447.892
R956 B.n99 B.t4 338.779
R957 B.n39 B.t11 338.779
R958 B.n105 B.t1 338.779
R959 B.n32 B.t8 338.779
R960 B.n100 B.t5 315.894
R961 B.n40 B.t10 315.894
R962 B.n106 B.t2 315.894
R963 B.n33 B.t7 315.894
R964 B.n509 B.n508 256.663
R965 B.n508 B.n507 235.042
R966 B.n508 B.n2 235.042
R967 B.n173 B.n122 163.367
R968 B.n174 B.n173 163.367
R969 B.n175 B.n174 163.367
R970 B.n175 B.n120 163.367
R971 B.n179 B.n120 163.367
R972 B.n180 B.n179 163.367
R973 B.n181 B.n180 163.367
R974 B.n181 B.n118 163.367
R975 B.n185 B.n118 163.367
R976 B.n186 B.n185 163.367
R977 B.n187 B.n186 163.367
R978 B.n187 B.n116 163.367
R979 B.n191 B.n116 163.367
R980 B.n192 B.n191 163.367
R981 B.n193 B.n192 163.367
R982 B.n193 B.n114 163.367
R983 B.n197 B.n114 163.367
R984 B.n198 B.n197 163.367
R985 B.n199 B.n198 163.367
R986 B.n199 B.n112 163.367
R987 B.n203 B.n112 163.367
R988 B.n204 B.n203 163.367
R989 B.n205 B.n204 163.367
R990 B.n205 B.n110 163.367
R991 B.n209 B.n110 163.367
R992 B.n210 B.n209 163.367
R993 B.n211 B.n210 163.367
R994 B.n211 B.n108 163.367
R995 B.n215 B.n108 163.367
R996 B.n216 B.n215 163.367
R997 B.n217 B.n216 163.367
R998 B.n217 B.n104 163.367
R999 B.n222 B.n104 163.367
R1000 B.n223 B.n222 163.367
R1001 B.n224 B.n223 163.367
R1002 B.n224 B.n102 163.367
R1003 B.n228 B.n102 163.367
R1004 B.n229 B.n228 163.367
R1005 B.n230 B.n229 163.367
R1006 B.n230 B.n98 163.367
R1007 B.n235 B.n98 163.367
R1008 B.n236 B.n235 163.367
R1009 B.n237 B.n236 163.367
R1010 B.n237 B.n96 163.367
R1011 B.n241 B.n96 163.367
R1012 B.n242 B.n241 163.367
R1013 B.n243 B.n242 163.367
R1014 B.n243 B.n94 163.367
R1015 B.n247 B.n94 163.367
R1016 B.n248 B.n247 163.367
R1017 B.n249 B.n248 163.367
R1018 B.n249 B.n92 163.367
R1019 B.n253 B.n92 163.367
R1020 B.n254 B.n253 163.367
R1021 B.n255 B.n254 163.367
R1022 B.n255 B.n90 163.367
R1023 B.n259 B.n90 163.367
R1024 B.n260 B.n259 163.367
R1025 B.n261 B.n260 163.367
R1026 B.n261 B.n88 163.367
R1027 B.n265 B.n88 163.367
R1028 B.n266 B.n265 163.367
R1029 B.n267 B.n266 163.367
R1030 B.n267 B.n86 163.367
R1031 B.n271 B.n86 163.367
R1032 B.n272 B.n271 163.367
R1033 B.n273 B.n272 163.367
R1034 B.n273 B.n84 163.367
R1035 B.n277 B.n84 163.367
R1036 B.n278 B.n277 163.367
R1037 B.n279 B.n278 163.367
R1038 B.n279 B.n82 163.367
R1039 B.n357 B.n56 163.367
R1040 B.n357 B.n356 163.367
R1041 B.n356 B.n355 163.367
R1042 B.n355 B.n58 163.367
R1043 B.n351 B.n58 163.367
R1044 B.n351 B.n350 163.367
R1045 B.n350 B.n349 163.367
R1046 B.n349 B.n60 163.367
R1047 B.n345 B.n60 163.367
R1048 B.n345 B.n344 163.367
R1049 B.n344 B.n343 163.367
R1050 B.n343 B.n62 163.367
R1051 B.n339 B.n62 163.367
R1052 B.n339 B.n338 163.367
R1053 B.n338 B.n337 163.367
R1054 B.n337 B.n64 163.367
R1055 B.n333 B.n64 163.367
R1056 B.n333 B.n332 163.367
R1057 B.n332 B.n331 163.367
R1058 B.n331 B.n66 163.367
R1059 B.n327 B.n66 163.367
R1060 B.n327 B.n326 163.367
R1061 B.n326 B.n325 163.367
R1062 B.n325 B.n68 163.367
R1063 B.n321 B.n68 163.367
R1064 B.n321 B.n320 163.367
R1065 B.n320 B.n319 163.367
R1066 B.n319 B.n70 163.367
R1067 B.n315 B.n70 163.367
R1068 B.n315 B.n314 163.367
R1069 B.n314 B.n313 163.367
R1070 B.n313 B.n72 163.367
R1071 B.n309 B.n72 163.367
R1072 B.n309 B.n308 163.367
R1073 B.n308 B.n307 163.367
R1074 B.n307 B.n74 163.367
R1075 B.n303 B.n74 163.367
R1076 B.n303 B.n302 163.367
R1077 B.n302 B.n301 163.367
R1078 B.n301 B.n76 163.367
R1079 B.n297 B.n76 163.367
R1080 B.n297 B.n296 163.367
R1081 B.n296 B.n295 163.367
R1082 B.n295 B.n78 163.367
R1083 B.n291 B.n78 163.367
R1084 B.n291 B.n290 163.367
R1085 B.n290 B.n289 163.367
R1086 B.n289 B.n80 163.367
R1087 B.n285 B.n80 163.367
R1088 B.n285 B.n284 163.367
R1089 B.n284 B.n283 163.367
R1090 B.n470 B.n15 163.367
R1091 B.n466 B.n15 163.367
R1092 B.n466 B.n465 163.367
R1093 B.n465 B.n464 163.367
R1094 B.n464 B.n17 163.367
R1095 B.n460 B.n17 163.367
R1096 B.n460 B.n459 163.367
R1097 B.n459 B.n458 163.367
R1098 B.n458 B.n19 163.367
R1099 B.n454 B.n19 163.367
R1100 B.n454 B.n453 163.367
R1101 B.n453 B.n452 163.367
R1102 B.n452 B.n21 163.367
R1103 B.n448 B.n21 163.367
R1104 B.n448 B.n447 163.367
R1105 B.n447 B.n446 163.367
R1106 B.n446 B.n23 163.367
R1107 B.n442 B.n23 163.367
R1108 B.n442 B.n441 163.367
R1109 B.n441 B.n440 163.367
R1110 B.n440 B.n25 163.367
R1111 B.n436 B.n25 163.367
R1112 B.n436 B.n435 163.367
R1113 B.n435 B.n434 163.367
R1114 B.n434 B.n27 163.367
R1115 B.n430 B.n27 163.367
R1116 B.n430 B.n429 163.367
R1117 B.n429 B.n428 163.367
R1118 B.n428 B.n29 163.367
R1119 B.n424 B.n29 163.367
R1120 B.n424 B.n423 163.367
R1121 B.n423 B.n422 163.367
R1122 B.n422 B.n31 163.367
R1123 B.n418 B.n31 163.367
R1124 B.n418 B.n417 163.367
R1125 B.n417 B.n416 163.367
R1126 B.n416 B.n36 163.367
R1127 B.n412 B.n36 163.367
R1128 B.n412 B.n411 163.367
R1129 B.n411 B.n410 163.367
R1130 B.n410 B.n38 163.367
R1131 B.n405 B.n38 163.367
R1132 B.n405 B.n404 163.367
R1133 B.n404 B.n403 163.367
R1134 B.n403 B.n42 163.367
R1135 B.n399 B.n42 163.367
R1136 B.n399 B.n398 163.367
R1137 B.n398 B.n397 163.367
R1138 B.n397 B.n44 163.367
R1139 B.n393 B.n44 163.367
R1140 B.n393 B.n392 163.367
R1141 B.n392 B.n391 163.367
R1142 B.n391 B.n46 163.367
R1143 B.n387 B.n46 163.367
R1144 B.n387 B.n386 163.367
R1145 B.n386 B.n385 163.367
R1146 B.n385 B.n48 163.367
R1147 B.n381 B.n48 163.367
R1148 B.n381 B.n380 163.367
R1149 B.n380 B.n379 163.367
R1150 B.n379 B.n50 163.367
R1151 B.n375 B.n50 163.367
R1152 B.n375 B.n374 163.367
R1153 B.n374 B.n373 163.367
R1154 B.n373 B.n52 163.367
R1155 B.n369 B.n52 163.367
R1156 B.n369 B.n368 163.367
R1157 B.n368 B.n367 163.367
R1158 B.n367 B.n54 163.367
R1159 B.n363 B.n54 163.367
R1160 B.n363 B.n362 163.367
R1161 B.n362 B.n361 163.367
R1162 B.n472 B.n471 163.367
R1163 B.n472 B.n13 163.367
R1164 B.n476 B.n13 163.367
R1165 B.n477 B.n476 163.367
R1166 B.n478 B.n477 163.367
R1167 B.n478 B.n11 163.367
R1168 B.n482 B.n11 163.367
R1169 B.n483 B.n482 163.367
R1170 B.n484 B.n483 163.367
R1171 B.n484 B.n9 163.367
R1172 B.n488 B.n9 163.367
R1173 B.n489 B.n488 163.367
R1174 B.n490 B.n489 163.367
R1175 B.n490 B.n7 163.367
R1176 B.n494 B.n7 163.367
R1177 B.n495 B.n494 163.367
R1178 B.n496 B.n495 163.367
R1179 B.n496 B.n5 163.367
R1180 B.n500 B.n5 163.367
R1181 B.n501 B.n500 163.367
R1182 B.n502 B.n501 163.367
R1183 B.n502 B.n3 163.367
R1184 B.n506 B.n3 163.367
R1185 B.n507 B.n506 163.367
R1186 B.n134 B.n2 163.367
R1187 B.n137 B.n134 163.367
R1188 B.n138 B.n137 163.367
R1189 B.n139 B.n138 163.367
R1190 B.n139 B.n132 163.367
R1191 B.n143 B.n132 163.367
R1192 B.n144 B.n143 163.367
R1193 B.n145 B.n144 163.367
R1194 B.n145 B.n130 163.367
R1195 B.n149 B.n130 163.367
R1196 B.n150 B.n149 163.367
R1197 B.n151 B.n150 163.367
R1198 B.n151 B.n128 163.367
R1199 B.n155 B.n128 163.367
R1200 B.n156 B.n155 163.367
R1201 B.n157 B.n156 163.367
R1202 B.n157 B.n126 163.367
R1203 B.n161 B.n126 163.367
R1204 B.n162 B.n161 163.367
R1205 B.n163 B.n162 163.367
R1206 B.n163 B.n124 163.367
R1207 B.n167 B.n124 163.367
R1208 B.n168 B.n167 163.367
R1209 B.n169 B.n168 163.367
R1210 B.n219 B.n106 59.5399
R1211 B.n233 B.n100 59.5399
R1212 B.n408 B.n40 59.5399
R1213 B.n34 B.n33 59.5399
R1214 B.n469 B.n14 33.5615
R1215 B.n360 B.n359 33.5615
R1216 B.n282 B.n281 33.5615
R1217 B.n171 B.n170 33.5615
R1218 B.n106 B.n105 22.8853
R1219 B.n100 B.n99 22.8853
R1220 B.n40 B.n39 22.8853
R1221 B.n33 B.n32 22.8853
R1222 B B.n509 18.0485
R1223 B.n473 B.n14 10.6151
R1224 B.n474 B.n473 10.6151
R1225 B.n475 B.n474 10.6151
R1226 B.n475 B.n12 10.6151
R1227 B.n479 B.n12 10.6151
R1228 B.n480 B.n479 10.6151
R1229 B.n481 B.n480 10.6151
R1230 B.n481 B.n10 10.6151
R1231 B.n485 B.n10 10.6151
R1232 B.n486 B.n485 10.6151
R1233 B.n487 B.n486 10.6151
R1234 B.n487 B.n8 10.6151
R1235 B.n491 B.n8 10.6151
R1236 B.n492 B.n491 10.6151
R1237 B.n493 B.n492 10.6151
R1238 B.n493 B.n6 10.6151
R1239 B.n497 B.n6 10.6151
R1240 B.n498 B.n497 10.6151
R1241 B.n499 B.n498 10.6151
R1242 B.n499 B.n4 10.6151
R1243 B.n503 B.n4 10.6151
R1244 B.n504 B.n503 10.6151
R1245 B.n505 B.n504 10.6151
R1246 B.n505 B.n0 10.6151
R1247 B.n469 B.n468 10.6151
R1248 B.n468 B.n467 10.6151
R1249 B.n467 B.n16 10.6151
R1250 B.n463 B.n16 10.6151
R1251 B.n463 B.n462 10.6151
R1252 B.n462 B.n461 10.6151
R1253 B.n461 B.n18 10.6151
R1254 B.n457 B.n18 10.6151
R1255 B.n457 B.n456 10.6151
R1256 B.n456 B.n455 10.6151
R1257 B.n455 B.n20 10.6151
R1258 B.n451 B.n20 10.6151
R1259 B.n451 B.n450 10.6151
R1260 B.n450 B.n449 10.6151
R1261 B.n449 B.n22 10.6151
R1262 B.n445 B.n22 10.6151
R1263 B.n445 B.n444 10.6151
R1264 B.n444 B.n443 10.6151
R1265 B.n443 B.n24 10.6151
R1266 B.n439 B.n24 10.6151
R1267 B.n439 B.n438 10.6151
R1268 B.n438 B.n437 10.6151
R1269 B.n437 B.n26 10.6151
R1270 B.n433 B.n26 10.6151
R1271 B.n433 B.n432 10.6151
R1272 B.n432 B.n431 10.6151
R1273 B.n431 B.n28 10.6151
R1274 B.n427 B.n28 10.6151
R1275 B.n427 B.n426 10.6151
R1276 B.n426 B.n425 10.6151
R1277 B.n425 B.n30 10.6151
R1278 B.n421 B.n420 10.6151
R1279 B.n420 B.n419 10.6151
R1280 B.n419 B.n35 10.6151
R1281 B.n415 B.n35 10.6151
R1282 B.n415 B.n414 10.6151
R1283 B.n414 B.n413 10.6151
R1284 B.n413 B.n37 10.6151
R1285 B.n409 B.n37 10.6151
R1286 B.n407 B.n406 10.6151
R1287 B.n406 B.n41 10.6151
R1288 B.n402 B.n41 10.6151
R1289 B.n402 B.n401 10.6151
R1290 B.n401 B.n400 10.6151
R1291 B.n400 B.n43 10.6151
R1292 B.n396 B.n43 10.6151
R1293 B.n396 B.n395 10.6151
R1294 B.n395 B.n394 10.6151
R1295 B.n394 B.n45 10.6151
R1296 B.n390 B.n45 10.6151
R1297 B.n390 B.n389 10.6151
R1298 B.n389 B.n388 10.6151
R1299 B.n388 B.n47 10.6151
R1300 B.n384 B.n47 10.6151
R1301 B.n384 B.n383 10.6151
R1302 B.n383 B.n382 10.6151
R1303 B.n382 B.n49 10.6151
R1304 B.n378 B.n49 10.6151
R1305 B.n378 B.n377 10.6151
R1306 B.n377 B.n376 10.6151
R1307 B.n376 B.n51 10.6151
R1308 B.n372 B.n51 10.6151
R1309 B.n372 B.n371 10.6151
R1310 B.n371 B.n370 10.6151
R1311 B.n370 B.n53 10.6151
R1312 B.n366 B.n53 10.6151
R1313 B.n366 B.n365 10.6151
R1314 B.n365 B.n364 10.6151
R1315 B.n364 B.n55 10.6151
R1316 B.n360 B.n55 10.6151
R1317 B.n359 B.n358 10.6151
R1318 B.n358 B.n57 10.6151
R1319 B.n354 B.n57 10.6151
R1320 B.n354 B.n353 10.6151
R1321 B.n353 B.n352 10.6151
R1322 B.n352 B.n59 10.6151
R1323 B.n348 B.n59 10.6151
R1324 B.n348 B.n347 10.6151
R1325 B.n347 B.n346 10.6151
R1326 B.n346 B.n61 10.6151
R1327 B.n342 B.n61 10.6151
R1328 B.n342 B.n341 10.6151
R1329 B.n341 B.n340 10.6151
R1330 B.n340 B.n63 10.6151
R1331 B.n336 B.n63 10.6151
R1332 B.n336 B.n335 10.6151
R1333 B.n335 B.n334 10.6151
R1334 B.n334 B.n65 10.6151
R1335 B.n330 B.n65 10.6151
R1336 B.n330 B.n329 10.6151
R1337 B.n329 B.n328 10.6151
R1338 B.n328 B.n67 10.6151
R1339 B.n324 B.n67 10.6151
R1340 B.n324 B.n323 10.6151
R1341 B.n323 B.n322 10.6151
R1342 B.n322 B.n69 10.6151
R1343 B.n318 B.n69 10.6151
R1344 B.n318 B.n317 10.6151
R1345 B.n317 B.n316 10.6151
R1346 B.n316 B.n71 10.6151
R1347 B.n312 B.n71 10.6151
R1348 B.n312 B.n311 10.6151
R1349 B.n311 B.n310 10.6151
R1350 B.n310 B.n73 10.6151
R1351 B.n306 B.n73 10.6151
R1352 B.n306 B.n305 10.6151
R1353 B.n305 B.n304 10.6151
R1354 B.n304 B.n75 10.6151
R1355 B.n300 B.n75 10.6151
R1356 B.n300 B.n299 10.6151
R1357 B.n299 B.n298 10.6151
R1358 B.n298 B.n77 10.6151
R1359 B.n294 B.n77 10.6151
R1360 B.n294 B.n293 10.6151
R1361 B.n293 B.n292 10.6151
R1362 B.n292 B.n79 10.6151
R1363 B.n288 B.n79 10.6151
R1364 B.n288 B.n287 10.6151
R1365 B.n287 B.n286 10.6151
R1366 B.n286 B.n81 10.6151
R1367 B.n282 B.n81 10.6151
R1368 B.n135 B.n1 10.6151
R1369 B.n136 B.n135 10.6151
R1370 B.n136 B.n133 10.6151
R1371 B.n140 B.n133 10.6151
R1372 B.n141 B.n140 10.6151
R1373 B.n142 B.n141 10.6151
R1374 B.n142 B.n131 10.6151
R1375 B.n146 B.n131 10.6151
R1376 B.n147 B.n146 10.6151
R1377 B.n148 B.n147 10.6151
R1378 B.n148 B.n129 10.6151
R1379 B.n152 B.n129 10.6151
R1380 B.n153 B.n152 10.6151
R1381 B.n154 B.n153 10.6151
R1382 B.n154 B.n127 10.6151
R1383 B.n158 B.n127 10.6151
R1384 B.n159 B.n158 10.6151
R1385 B.n160 B.n159 10.6151
R1386 B.n160 B.n125 10.6151
R1387 B.n164 B.n125 10.6151
R1388 B.n165 B.n164 10.6151
R1389 B.n166 B.n165 10.6151
R1390 B.n166 B.n123 10.6151
R1391 B.n170 B.n123 10.6151
R1392 B.n172 B.n171 10.6151
R1393 B.n172 B.n121 10.6151
R1394 B.n176 B.n121 10.6151
R1395 B.n177 B.n176 10.6151
R1396 B.n178 B.n177 10.6151
R1397 B.n178 B.n119 10.6151
R1398 B.n182 B.n119 10.6151
R1399 B.n183 B.n182 10.6151
R1400 B.n184 B.n183 10.6151
R1401 B.n184 B.n117 10.6151
R1402 B.n188 B.n117 10.6151
R1403 B.n189 B.n188 10.6151
R1404 B.n190 B.n189 10.6151
R1405 B.n190 B.n115 10.6151
R1406 B.n194 B.n115 10.6151
R1407 B.n195 B.n194 10.6151
R1408 B.n196 B.n195 10.6151
R1409 B.n196 B.n113 10.6151
R1410 B.n200 B.n113 10.6151
R1411 B.n201 B.n200 10.6151
R1412 B.n202 B.n201 10.6151
R1413 B.n202 B.n111 10.6151
R1414 B.n206 B.n111 10.6151
R1415 B.n207 B.n206 10.6151
R1416 B.n208 B.n207 10.6151
R1417 B.n208 B.n109 10.6151
R1418 B.n212 B.n109 10.6151
R1419 B.n213 B.n212 10.6151
R1420 B.n214 B.n213 10.6151
R1421 B.n214 B.n107 10.6151
R1422 B.n218 B.n107 10.6151
R1423 B.n221 B.n220 10.6151
R1424 B.n221 B.n103 10.6151
R1425 B.n225 B.n103 10.6151
R1426 B.n226 B.n225 10.6151
R1427 B.n227 B.n226 10.6151
R1428 B.n227 B.n101 10.6151
R1429 B.n231 B.n101 10.6151
R1430 B.n232 B.n231 10.6151
R1431 B.n234 B.n97 10.6151
R1432 B.n238 B.n97 10.6151
R1433 B.n239 B.n238 10.6151
R1434 B.n240 B.n239 10.6151
R1435 B.n240 B.n95 10.6151
R1436 B.n244 B.n95 10.6151
R1437 B.n245 B.n244 10.6151
R1438 B.n246 B.n245 10.6151
R1439 B.n246 B.n93 10.6151
R1440 B.n250 B.n93 10.6151
R1441 B.n251 B.n250 10.6151
R1442 B.n252 B.n251 10.6151
R1443 B.n252 B.n91 10.6151
R1444 B.n256 B.n91 10.6151
R1445 B.n257 B.n256 10.6151
R1446 B.n258 B.n257 10.6151
R1447 B.n258 B.n89 10.6151
R1448 B.n262 B.n89 10.6151
R1449 B.n263 B.n262 10.6151
R1450 B.n264 B.n263 10.6151
R1451 B.n264 B.n87 10.6151
R1452 B.n268 B.n87 10.6151
R1453 B.n269 B.n268 10.6151
R1454 B.n270 B.n269 10.6151
R1455 B.n270 B.n85 10.6151
R1456 B.n274 B.n85 10.6151
R1457 B.n275 B.n274 10.6151
R1458 B.n276 B.n275 10.6151
R1459 B.n276 B.n83 10.6151
R1460 B.n280 B.n83 10.6151
R1461 B.n281 B.n280 10.6151
R1462 B.n509 B.n0 8.11757
R1463 B.n509 B.n1 8.11757
R1464 B.n421 B.n34 6.5566
R1465 B.n409 B.n408 6.5566
R1466 B.n220 B.n219 6.5566
R1467 B.n233 B.n232 6.5566
R1468 B.n34 B.n30 4.05904
R1469 B.n408 B.n407 4.05904
R1470 B.n219 B.n218 4.05904
R1471 B.n234 B.n233 4.05904
C0 w_n2150_n2704# VN 3.81983f
C1 VP VTAIL 4.44968f
C2 VP VN 4.90379f
C3 VDD2 VTAIL 8.04513f
C4 VDD1 VTAIL 8.00244f
C5 VDD2 VN 4.49432f
C6 VDD1 VN 0.148591f
C7 B VTAIL 3.03957f
C8 B VN 0.780034f
C9 w_n2150_n2704# VP 4.09379f
C10 VDD2 w_n2150_n2704# 1.30501f
C11 w_n2150_n2704# VDD1 1.26395f
C12 VN VTAIL 4.43558f
C13 VDD2 VP 0.333479f
C14 VDD1 VP 4.6787f
C15 B w_n2150_n2704# 6.50654f
C16 B VP 1.22995f
C17 VDD2 VDD1 0.898604f
C18 VDD2 B 1.06769f
C19 B VDD1 1.02639f
C20 w_n2150_n2704# VTAIL 3.36112f
C21 VDD2 VSUBS 1.233564f
C22 VDD1 VSUBS 1.570296f
C23 VTAIL VSUBS 0.810194f
C24 VN VSUBS 4.55054f
C25 VP VSUBS 1.67356f
C26 B VSUBS 2.773225f
C27 w_n2150_n2704# VSUBS 72.0078f
C28 B.n0 VSUBS 0.007422f
C29 B.n1 VSUBS 0.007422f
C30 B.n2 VSUBS 0.010977f
C31 B.n3 VSUBS 0.008412f
C32 B.n4 VSUBS 0.008412f
C33 B.n5 VSUBS 0.008412f
C34 B.n6 VSUBS 0.008412f
C35 B.n7 VSUBS 0.008412f
C36 B.n8 VSUBS 0.008412f
C37 B.n9 VSUBS 0.008412f
C38 B.n10 VSUBS 0.008412f
C39 B.n11 VSUBS 0.008412f
C40 B.n12 VSUBS 0.008412f
C41 B.n13 VSUBS 0.008412f
C42 B.n14 VSUBS 0.019721f
C43 B.n15 VSUBS 0.008412f
C44 B.n16 VSUBS 0.008412f
C45 B.n17 VSUBS 0.008412f
C46 B.n18 VSUBS 0.008412f
C47 B.n19 VSUBS 0.008412f
C48 B.n20 VSUBS 0.008412f
C49 B.n21 VSUBS 0.008412f
C50 B.n22 VSUBS 0.008412f
C51 B.n23 VSUBS 0.008412f
C52 B.n24 VSUBS 0.008412f
C53 B.n25 VSUBS 0.008412f
C54 B.n26 VSUBS 0.008412f
C55 B.n27 VSUBS 0.008412f
C56 B.n28 VSUBS 0.008412f
C57 B.n29 VSUBS 0.008412f
C58 B.n30 VSUBS 0.005814f
C59 B.n31 VSUBS 0.008412f
C60 B.t7 VSUBS 0.168481f
C61 B.t8 VSUBS 0.183528f
C62 B.t6 VSUBS 0.379167f
C63 B.n32 VSUBS 0.292062f
C64 B.n33 VSUBS 0.23476f
C65 B.n34 VSUBS 0.019489f
C66 B.n35 VSUBS 0.008412f
C67 B.n36 VSUBS 0.008412f
C68 B.n37 VSUBS 0.008412f
C69 B.n38 VSUBS 0.008412f
C70 B.t10 VSUBS 0.168484f
C71 B.t11 VSUBS 0.183531f
C72 B.t9 VSUBS 0.379167f
C73 B.n39 VSUBS 0.292059f
C74 B.n40 VSUBS 0.234757f
C75 B.n41 VSUBS 0.008412f
C76 B.n42 VSUBS 0.008412f
C77 B.n43 VSUBS 0.008412f
C78 B.n44 VSUBS 0.008412f
C79 B.n45 VSUBS 0.008412f
C80 B.n46 VSUBS 0.008412f
C81 B.n47 VSUBS 0.008412f
C82 B.n48 VSUBS 0.008412f
C83 B.n49 VSUBS 0.008412f
C84 B.n50 VSUBS 0.008412f
C85 B.n51 VSUBS 0.008412f
C86 B.n52 VSUBS 0.008412f
C87 B.n53 VSUBS 0.008412f
C88 B.n54 VSUBS 0.008412f
C89 B.n55 VSUBS 0.008412f
C90 B.n56 VSUBS 0.019721f
C91 B.n57 VSUBS 0.008412f
C92 B.n58 VSUBS 0.008412f
C93 B.n59 VSUBS 0.008412f
C94 B.n60 VSUBS 0.008412f
C95 B.n61 VSUBS 0.008412f
C96 B.n62 VSUBS 0.008412f
C97 B.n63 VSUBS 0.008412f
C98 B.n64 VSUBS 0.008412f
C99 B.n65 VSUBS 0.008412f
C100 B.n66 VSUBS 0.008412f
C101 B.n67 VSUBS 0.008412f
C102 B.n68 VSUBS 0.008412f
C103 B.n69 VSUBS 0.008412f
C104 B.n70 VSUBS 0.008412f
C105 B.n71 VSUBS 0.008412f
C106 B.n72 VSUBS 0.008412f
C107 B.n73 VSUBS 0.008412f
C108 B.n74 VSUBS 0.008412f
C109 B.n75 VSUBS 0.008412f
C110 B.n76 VSUBS 0.008412f
C111 B.n77 VSUBS 0.008412f
C112 B.n78 VSUBS 0.008412f
C113 B.n79 VSUBS 0.008412f
C114 B.n80 VSUBS 0.008412f
C115 B.n81 VSUBS 0.008412f
C116 B.n82 VSUBS 0.020358f
C117 B.n83 VSUBS 0.008412f
C118 B.n84 VSUBS 0.008412f
C119 B.n85 VSUBS 0.008412f
C120 B.n86 VSUBS 0.008412f
C121 B.n87 VSUBS 0.008412f
C122 B.n88 VSUBS 0.008412f
C123 B.n89 VSUBS 0.008412f
C124 B.n90 VSUBS 0.008412f
C125 B.n91 VSUBS 0.008412f
C126 B.n92 VSUBS 0.008412f
C127 B.n93 VSUBS 0.008412f
C128 B.n94 VSUBS 0.008412f
C129 B.n95 VSUBS 0.008412f
C130 B.n96 VSUBS 0.008412f
C131 B.n97 VSUBS 0.008412f
C132 B.n98 VSUBS 0.008412f
C133 B.t5 VSUBS 0.168484f
C134 B.t4 VSUBS 0.183531f
C135 B.t3 VSUBS 0.379167f
C136 B.n99 VSUBS 0.292059f
C137 B.n100 VSUBS 0.234757f
C138 B.n101 VSUBS 0.008412f
C139 B.n102 VSUBS 0.008412f
C140 B.n103 VSUBS 0.008412f
C141 B.n104 VSUBS 0.008412f
C142 B.t2 VSUBS 0.168481f
C143 B.t1 VSUBS 0.183528f
C144 B.t0 VSUBS 0.379167f
C145 B.n105 VSUBS 0.292062f
C146 B.n106 VSUBS 0.23476f
C147 B.n107 VSUBS 0.008412f
C148 B.n108 VSUBS 0.008412f
C149 B.n109 VSUBS 0.008412f
C150 B.n110 VSUBS 0.008412f
C151 B.n111 VSUBS 0.008412f
C152 B.n112 VSUBS 0.008412f
C153 B.n113 VSUBS 0.008412f
C154 B.n114 VSUBS 0.008412f
C155 B.n115 VSUBS 0.008412f
C156 B.n116 VSUBS 0.008412f
C157 B.n117 VSUBS 0.008412f
C158 B.n118 VSUBS 0.008412f
C159 B.n119 VSUBS 0.008412f
C160 B.n120 VSUBS 0.008412f
C161 B.n121 VSUBS 0.008412f
C162 B.n122 VSUBS 0.020358f
C163 B.n123 VSUBS 0.008412f
C164 B.n124 VSUBS 0.008412f
C165 B.n125 VSUBS 0.008412f
C166 B.n126 VSUBS 0.008412f
C167 B.n127 VSUBS 0.008412f
C168 B.n128 VSUBS 0.008412f
C169 B.n129 VSUBS 0.008412f
C170 B.n130 VSUBS 0.008412f
C171 B.n131 VSUBS 0.008412f
C172 B.n132 VSUBS 0.008412f
C173 B.n133 VSUBS 0.008412f
C174 B.n134 VSUBS 0.008412f
C175 B.n135 VSUBS 0.008412f
C176 B.n136 VSUBS 0.008412f
C177 B.n137 VSUBS 0.008412f
C178 B.n138 VSUBS 0.008412f
C179 B.n139 VSUBS 0.008412f
C180 B.n140 VSUBS 0.008412f
C181 B.n141 VSUBS 0.008412f
C182 B.n142 VSUBS 0.008412f
C183 B.n143 VSUBS 0.008412f
C184 B.n144 VSUBS 0.008412f
C185 B.n145 VSUBS 0.008412f
C186 B.n146 VSUBS 0.008412f
C187 B.n147 VSUBS 0.008412f
C188 B.n148 VSUBS 0.008412f
C189 B.n149 VSUBS 0.008412f
C190 B.n150 VSUBS 0.008412f
C191 B.n151 VSUBS 0.008412f
C192 B.n152 VSUBS 0.008412f
C193 B.n153 VSUBS 0.008412f
C194 B.n154 VSUBS 0.008412f
C195 B.n155 VSUBS 0.008412f
C196 B.n156 VSUBS 0.008412f
C197 B.n157 VSUBS 0.008412f
C198 B.n158 VSUBS 0.008412f
C199 B.n159 VSUBS 0.008412f
C200 B.n160 VSUBS 0.008412f
C201 B.n161 VSUBS 0.008412f
C202 B.n162 VSUBS 0.008412f
C203 B.n163 VSUBS 0.008412f
C204 B.n164 VSUBS 0.008412f
C205 B.n165 VSUBS 0.008412f
C206 B.n166 VSUBS 0.008412f
C207 B.n167 VSUBS 0.008412f
C208 B.n168 VSUBS 0.008412f
C209 B.n169 VSUBS 0.019721f
C210 B.n170 VSUBS 0.019721f
C211 B.n171 VSUBS 0.020358f
C212 B.n172 VSUBS 0.008412f
C213 B.n173 VSUBS 0.008412f
C214 B.n174 VSUBS 0.008412f
C215 B.n175 VSUBS 0.008412f
C216 B.n176 VSUBS 0.008412f
C217 B.n177 VSUBS 0.008412f
C218 B.n178 VSUBS 0.008412f
C219 B.n179 VSUBS 0.008412f
C220 B.n180 VSUBS 0.008412f
C221 B.n181 VSUBS 0.008412f
C222 B.n182 VSUBS 0.008412f
C223 B.n183 VSUBS 0.008412f
C224 B.n184 VSUBS 0.008412f
C225 B.n185 VSUBS 0.008412f
C226 B.n186 VSUBS 0.008412f
C227 B.n187 VSUBS 0.008412f
C228 B.n188 VSUBS 0.008412f
C229 B.n189 VSUBS 0.008412f
C230 B.n190 VSUBS 0.008412f
C231 B.n191 VSUBS 0.008412f
C232 B.n192 VSUBS 0.008412f
C233 B.n193 VSUBS 0.008412f
C234 B.n194 VSUBS 0.008412f
C235 B.n195 VSUBS 0.008412f
C236 B.n196 VSUBS 0.008412f
C237 B.n197 VSUBS 0.008412f
C238 B.n198 VSUBS 0.008412f
C239 B.n199 VSUBS 0.008412f
C240 B.n200 VSUBS 0.008412f
C241 B.n201 VSUBS 0.008412f
C242 B.n202 VSUBS 0.008412f
C243 B.n203 VSUBS 0.008412f
C244 B.n204 VSUBS 0.008412f
C245 B.n205 VSUBS 0.008412f
C246 B.n206 VSUBS 0.008412f
C247 B.n207 VSUBS 0.008412f
C248 B.n208 VSUBS 0.008412f
C249 B.n209 VSUBS 0.008412f
C250 B.n210 VSUBS 0.008412f
C251 B.n211 VSUBS 0.008412f
C252 B.n212 VSUBS 0.008412f
C253 B.n213 VSUBS 0.008412f
C254 B.n214 VSUBS 0.008412f
C255 B.n215 VSUBS 0.008412f
C256 B.n216 VSUBS 0.008412f
C257 B.n217 VSUBS 0.008412f
C258 B.n218 VSUBS 0.005814f
C259 B.n219 VSUBS 0.019489f
C260 B.n220 VSUBS 0.006803f
C261 B.n221 VSUBS 0.008412f
C262 B.n222 VSUBS 0.008412f
C263 B.n223 VSUBS 0.008412f
C264 B.n224 VSUBS 0.008412f
C265 B.n225 VSUBS 0.008412f
C266 B.n226 VSUBS 0.008412f
C267 B.n227 VSUBS 0.008412f
C268 B.n228 VSUBS 0.008412f
C269 B.n229 VSUBS 0.008412f
C270 B.n230 VSUBS 0.008412f
C271 B.n231 VSUBS 0.008412f
C272 B.n232 VSUBS 0.006803f
C273 B.n233 VSUBS 0.019489f
C274 B.n234 VSUBS 0.005814f
C275 B.n235 VSUBS 0.008412f
C276 B.n236 VSUBS 0.008412f
C277 B.n237 VSUBS 0.008412f
C278 B.n238 VSUBS 0.008412f
C279 B.n239 VSUBS 0.008412f
C280 B.n240 VSUBS 0.008412f
C281 B.n241 VSUBS 0.008412f
C282 B.n242 VSUBS 0.008412f
C283 B.n243 VSUBS 0.008412f
C284 B.n244 VSUBS 0.008412f
C285 B.n245 VSUBS 0.008412f
C286 B.n246 VSUBS 0.008412f
C287 B.n247 VSUBS 0.008412f
C288 B.n248 VSUBS 0.008412f
C289 B.n249 VSUBS 0.008412f
C290 B.n250 VSUBS 0.008412f
C291 B.n251 VSUBS 0.008412f
C292 B.n252 VSUBS 0.008412f
C293 B.n253 VSUBS 0.008412f
C294 B.n254 VSUBS 0.008412f
C295 B.n255 VSUBS 0.008412f
C296 B.n256 VSUBS 0.008412f
C297 B.n257 VSUBS 0.008412f
C298 B.n258 VSUBS 0.008412f
C299 B.n259 VSUBS 0.008412f
C300 B.n260 VSUBS 0.008412f
C301 B.n261 VSUBS 0.008412f
C302 B.n262 VSUBS 0.008412f
C303 B.n263 VSUBS 0.008412f
C304 B.n264 VSUBS 0.008412f
C305 B.n265 VSUBS 0.008412f
C306 B.n266 VSUBS 0.008412f
C307 B.n267 VSUBS 0.008412f
C308 B.n268 VSUBS 0.008412f
C309 B.n269 VSUBS 0.008412f
C310 B.n270 VSUBS 0.008412f
C311 B.n271 VSUBS 0.008412f
C312 B.n272 VSUBS 0.008412f
C313 B.n273 VSUBS 0.008412f
C314 B.n274 VSUBS 0.008412f
C315 B.n275 VSUBS 0.008412f
C316 B.n276 VSUBS 0.008412f
C317 B.n277 VSUBS 0.008412f
C318 B.n278 VSUBS 0.008412f
C319 B.n279 VSUBS 0.008412f
C320 B.n280 VSUBS 0.008412f
C321 B.n281 VSUBS 0.01939f
C322 B.n282 VSUBS 0.020688f
C323 B.n283 VSUBS 0.019721f
C324 B.n284 VSUBS 0.008412f
C325 B.n285 VSUBS 0.008412f
C326 B.n286 VSUBS 0.008412f
C327 B.n287 VSUBS 0.008412f
C328 B.n288 VSUBS 0.008412f
C329 B.n289 VSUBS 0.008412f
C330 B.n290 VSUBS 0.008412f
C331 B.n291 VSUBS 0.008412f
C332 B.n292 VSUBS 0.008412f
C333 B.n293 VSUBS 0.008412f
C334 B.n294 VSUBS 0.008412f
C335 B.n295 VSUBS 0.008412f
C336 B.n296 VSUBS 0.008412f
C337 B.n297 VSUBS 0.008412f
C338 B.n298 VSUBS 0.008412f
C339 B.n299 VSUBS 0.008412f
C340 B.n300 VSUBS 0.008412f
C341 B.n301 VSUBS 0.008412f
C342 B.n302 VSUBS 0.008412f
C343 B.n303 VSUBS 0.008412f
C344 B.n304 VSUBS 0.008412f
C345 B.n305 VSUBS 0.008412f
C346 B.n306 VSUBS 0.008412f
C347 B.n307 VSUBS 0.008412f
C348 B.n308 VSUBS 0.008412f
C349 B.n309 VSUBS 0.008412f
C350 B.n310 VSUBS 0.008412f
C351 B.n311 VSUBS 0.008412f
C352 B.n312 VSUBS 0.008412f
C353 B.n313 VSUBS 0.008412f
C354 B.n314 VSUBS 0.008412f
C355 B.n315 VSUBS 0.008412f
C356 B.n316 VSUBS 0.008412f
C357 B.n317 VSUBS 0.008412f
C358 B.n318 VSUBS 0.008412f
C359 B.n319 VSUBS 0.008412f
C360 B.n320 VSUBS 0.008412f
C361 B.n321 VSUBS 0.008412f
C362 B.n322 VSUBS 0.008412f
C363 B.n323 VSUBS 0.008412f
C364 B.n324 VSUBS 0.008412f
C365 B.n325 VSUBS 0.008412f
C366 B.n326 VSUBS 0.008412f
C367 B.n327 VSUBS 0.008412f
C368 B.n328 VSUBS 0.008412f
C369 B.n329 VSUBS 0.008412f
C370 B.n330 VSUBS 0.008412f
C371 B.n331 VSUBS 0.008412f
C372 B.n332 VSUBS 0.008412f
C373 B.n333 VSUBS 0.008412f
C374 B.n334 VSUBS 0.008412f
C375 B.n335 VSUBS 0.008412f
C376 B.n336 VSUBS 0.008412f
C377 B.n337 VSUBS 0.008412f
C378 B.n338 VSUBS 0.008412f
C379 B.n339 VSUBS 0.008412f
C380 B.n340 VSUBS 0.008412f
C381 B.n341 VSUBS 0.008412f
C382 B.n342 VSUBS 0.008412f
C383 B.n343 VSUBS 0.008412f
C384 B.n344 VSUBS 0.008412f
C385 B.n345 VSUBS 0.008412f
C386 B.n346 VSUBS 0.008412f
C387 B.n347 VSUBS 0.008412f
C388 B.n348 VSUBS 0.008412f
C389 B.n349 VSUBS 0.008412f
C390 B.n350 VSUBS 0.008412f
C391 B.n351 VSUBS 0.008412f
C392 B.n352 VSUBS 0.008412f
C393 B.n353 VSUBS 0.008412f
C394 B.n354 VSUBS 0.008412f
C395 B.n355 VSUBS 0.008412f
C396 B.n356 VSUBS 0.008412f
C397 B.n357 VSUBS 0.008412f
C398 B.n358 VSUBS 0.008412f
C399 B.n359 VSUBS 0.019721f
C400 B.n360 VSUBS 0.020358f
C401 B.n361 VSUBS 0.020358f
C402 B.n362 VSUBS 0.008412f
C403 B.n363 VSUBS 0.008412f
C404 B.n364 VSUBS 0.008412f
C405 B.n365 VSUBS 0.008412f
C406 B.n366 VSUBS 0.008412f
C407 B.n367 VSUBS 0.008412f
C408 B.n368 VSUBS 0.008412f
C409 B.n369 VSUBS 0.008412f
C410 B.n370 VSUBS 0.008412f
C411 B.n371 VSUBS 0.008412f
C412 B.n372 VSUBS 0.008412f
C413 B.n373 VSUBS 0.008412f
C414 B.n374 VSUBS 0.008412f
C415 B.n375 VSUBS 0.008412f
C416 B.n376 VSUBS 0.008412f
C417 B.n377 VSUBS 0.008412f
C418 B.n378 VSUBS 0.008412f
C419 B.n379 VSUBS 0.008412f
C420 B.n380 VSUBS 0.008412f
C421 B.n381 VSUBS 0.008412f
C422 B.n382 VSUBS 0.008412f
C423 B.n383 VSUBS 0.008412f
C424 B.n384 VSUBS 0.008412f
C425 B.n385 VSUBS 0.008412f
C426 B.n386 VSUBS 0.008412f
C427 B.n387 VSUBS 0.008412f
C428 B.n388 VSUBS 0.008412f
C429 B.n389 VSUBS 0.008412f
C430 B.n390 VSUBS 0.008412f
C431 B.n391 VSUBS 0.008412f
C432 B.n392 VSUBS 0.008412f
C433 B.n393 VSUBS 0.008412f
C434 B.n394 VSUBS 0.008412f
C435 B.n395 VSUBS 0.008412f
C436 B.n396 VSUBS 0.008412f
C437 B.n397 VSUBS 0.008412f
C438 B.n398 VSUBS 0.008412f
C439 B.n399 VSUBS 0.008412f
C440 B.n400 VSUBS 0.008412f
C441 B.n401 VSUBS 0.008412f
C442 B.n402 VSUBS 0.008412f
C443 B.n403 VSUBS 0.008412f
C444 B.n404 VSUBS 0.008412f
C445 B.n405 VSUBS 0.008412f
C446 B.n406 VSUBS 0.008412f
C447 B.n407 VSUBS 0.005814f
C448 B.n408 VSUBS 0.019489f
C449 B.n409 VSUBS 0.006803f
C450 B.n410 VSUBS 0.008412f
C451 B.n411 VSUBS 0.008412f
C452 B.n412 VSUBS 0.008412f
C453 B.n413 VSUBS 0.008412f
C454 B.n414 VSUBS 0.008412f
C455 B.n415 VSUBS 0.008412f
C456 B.n416 VSUBS 0.008412f
C457 B.n417 VSUBS 0.008412f
C458 B.n418 VSUBS 0.008412f
C459 B.n419 VSUBS 0.008412f
C460 B.n420 VSUBS 0.008412f
C461 B.n421 VSUBS 0.006803f
C462 B.n422 VSUBS 0.008412f
C463 B.n423 VSUBS 0.008412f
C464 B.n424 VSUBS 0.008412f
C465 B.n425 VSUBS 0.008412f
C466 B.n426 VSUBS 0.008412f
C467 B.n427 VSUBS 0.008412f
C468 B.n428 VSUBS 0.008412f
C469 B.n429 VSUBS 0.008412f
C470 B.n430 VSUBS 0.008412f
C471 B.n431 VSUBS 0.008412f
C472 B.n432 VSUBS 0.008412f
C473 B.n433 VSUBS 0.008412f
C474 B.n434 VSUBS 0.008412f
C475 B.n435 VSUBS 0.008412f
C476 B.n436 VSUBS 0.008412f
C477 B.n437 VSUBS 0.008412f
C478 B.n438 VSUBS 0.008412f
C479 B.n439 VSUBS 0.008412f
C480 B.n440 VSUBS 0.008412f
C481 B.n441 VSUBS 0.008412f
C482 B.n442 VSUBS 0.008412f
C483 B.n443 VSUBS 0.008412f
C484 B.n444 VSUBS 0.008412f
C485 B.n445 VSUBS 0.008412f
C486 B.n446 VSUBS 0.008412f
C487 B.n447 VSUBS 0.008412f
C488 B.n448 VSUBS 0.008412f
C489 B.n449 VSUBS 0.008412f
C490 B.n450 VSUBS 0.008412f
C491 B.n451 VSUBS 0.008412f
C492 B.n452 VSUBS 0.008412f
C493 B.n453 VSUBS 0.008412f
C494 B.n454 VSUBS 0.008412f
C495 B.n455 VSUBS 0.008412f
C496 B.n456 VSUBS 0.008412f
C497 B.n457 VSUBS 0.008412f
C498 B.n458 VSUBS 0.008412f
C499 B.n459 VSUBS 0.008412f
C500 B.n460 VSUBS 0.008412f
C501 B.n461 VSUBS 0.008412f
C502 B.n462 VSUBS 0.008412f
C503 B.n463 VSUBS 0.008412f
C504 B.n464 VSUBS 0.008412f
C505 B.n465 VSUBS 0.008412f
C506 B.n466 VSUBS 0.008412f
C507 B.n467 VSUBS 0.008412f
C508 B.n468 VSUBS 0.008412f
C509 B.n469 VSUBS 0.020358f
C510 B.n470 VSUBS 0.020358f
C511 B.n471 VSUBS 0.019721f
C512 B.n472 VSUBS 0.008412f
C513 B.n473 VSUBS 0.008412f
C514 B.n474 VSUBS 0.008412f
C515 B.n475 VSUBS 0.008412f
C516 B.n476 VSUBS 0.008412f
C517 B.n477 VSUBS 0.008412f
C518 B.n478 VSUBS 0.008412f
C519 B.n479 VSUBS 0.008412f
C520 B.n480 VSUBS 0.008412f
C521 B.n481 VSUBS 0.008412f
C522 B.n482 VSUBS 0.008412f
C523 B.n483 VSUBS 0.008412f
C524 B.n484 VSUBS 0.008412f
C525 B.n485 VSUBS 0.008412f
C526 B.n486 VSUBS 0.008412f
C527 B.n487 VSUBS 0.008412f
C528 B.n488 VSUBS 0.008412f
C529 B.n489 VSUBS 0.008412f
C530 B.n490 VSUBS 0.008412f
C531 B.n491 VSUBS 0.008412f
C532 B.n492 VSUBS 0.008412f
C533 B.n493 VSUBS 0.008412f
C534 B.n494 VSUBS 0.008412f
C535 B.n495 VSUBS 0.008412f
C536 B.n496 VSUBS 0.008412f
C537 B.n497 VSUBS 0.008412f
C538 B.n498 VSUBS 0.008412f
C539 B.n499 VSUBS 0.008412f
C540 B.n500 VSUBS 0.008412f
C541 B.n501 VSUBS 0.008412f
C542 B.n502 VSUBS 0.008412f
C543 B.n503 VSUBS 0.008412f
C544 B.n504 VSUBS 0.008412f
C545 B.n505 VSUBS 0.008412f
C546 B.n506 VSUBS 0.008412f
C547 B.n507 VSUBS 0.010977f
C548 B.n508 VSUBS 0.011693f
C549 B.n509 VSUBS 0.023252f
C550 VDD2.t0 VSUBS 0.180254f
C551 VDD2.t5 VSUBS 0.180254f
C552 VDD2.n0 VSUBS 1.33385f
C553 VDD2.t4 VSUBS 0.180254f
C554 VDD2.t1 VSUBS 0.180254f
C555 VDD2.n1 VSUBS 1.33385f
C556 VDD2.n2 VSUBS 2.63239f
C557 VDD2.t2 VSUBS 0.180254f
C558 VDD2.t7 VSUBS 0.180254f
C559 VDD2.n3 VSUBS 1.33068f
C560 VDD2.n4 VSUBS 2.42419f
C561 VDD2.t6 VSUBS 0.180254f
C562 VDD2.t3 VSUBS 0.180254f
C563 VDD2.n5 VSUBS 1.33382f
C564 VN.n0 VSUBS 0.052483f
C565 VN.t3 VSUBS 1.0435f
C566 VN.n1 VSUBS 0.409773f
C567 VN.n2 VSUBS 0.221441f
C568 VN.t2 VSUBS 1.0435f
C569 VN.t7 VSUBS 1.14317f
C570 VN.n3 VSUBS 0.463624f
C571 VN.n4 VSUBS 0.464042f
C572 VN.n5 VSUBS 0.060918f
C573 VN.n6 VSUBS 0.060918f
C574 VN.n7 VSUBS 0.052483f
C575 VN.n8 VSUBS 0.052483f
C576 VN.n9 VSUBS 0.066039f
C577 VN.n10 VSUBS 0.021011f
C578 VN.t6 VSUBS 1.11143f
C579 VN.n11 VSUBS 0.461464f
C580 VN.n12 VSUBS 0.040673f
C581 VN.n13 VSUBS 0.052483f
C582 VN.t0 VSUBS 1.0435f
C583 VN.n14 VSUBS 0.409773f
C584 VN.n15 VSUBS 0.221441f
C585 VN.t1 VSUBS 1.0435f
C586 VN.t4 VSUBS 1.14317f
C587 VN.n16 VSUBS 0.463624f
C588 VN.n17 VSUBS 0.464042f
C589 VN.n18 VSUBS 0.060918f
C590 VN.n19 VSUBS 0.060918f
C591 VN.n20 VSUBS 0.052483f
C592 VN.n21 VSUBS 0.052483f
C593 VN.n22 VSUBS 0.066039f
C594 VN.n23 VSUBS 0.021011f
C595 VN.t5 VSUBS 1.11143f
C596 VN.n24 VSUBS 0.461464f
C597 VN.n25 VSUBS 2.04584f
C598 VDD1.t4 VSUBS 0.181727f
C599 VDD1.t6 VSUBS 0.181727f
C600 VDD1.n0 VSUBS 1.34561f
C601 VDD1.t2 VSUBS 0.181727f
C602 VDD1.t3 VSUBS 0.181727f
C603 VDD1.n1 VSUBS 1.34475f
C604 VDD1.t5 VSUBS 0.181727f
C605 VDD1.t7 VSUBS 0.181727f
C606 VDD1.n2 VSUBS 1.34475f
C607 VDD1.n3 VSUBS 2.71047f
C608 VDD1.t0 VSUBS 0.181727f
C609 VDD1.t1 VSUBS 0.181727f
C610 VDD1.n4 VSUBS 1.34155f
C611 VDD1.n5 VSUBS 2.47535f
C612 VTAIL.t5 VSUBS 0.174794f
C613 VTAIL.t4 VSUBS 0.174794f
C614 VTAIL.n0 VSUBS 1.18219f
C615 VTAIL.n1 VSUBS 0.599516f
C616 VTAIL.n2 VSUBS 0.027462f
C617 VTAIL.n3 VSUBS 0.025483f
C618 VTAIL.n4 VSUBS 0.013693f
C619 VTAIL.n5 VSUBS 0.032367f
C620 VTAIL.n6 VSUBS 0.014499f
C621 VTAIL.n7 VSUBS 0.025483f
C622 VTAIL.n8 VSUBS 0.013693f
C623 VTAIL.n9 VSUBS 0.032367f
C624 VTAIL.n10 VSUBS 0.014499f
C625 VTAIL.n11 VSUBS 0.025483f
C626 VTAIL.n12 VSUBS 0.013693f
C627 VTAIL.n13 VSUBS 0.032367f
C628 VTAIL.n14 VSUBS 0.014499f
C629 VTAIL.n15 VSUBS 0.162504f
C630 VTAIL.t3 VSUBS 0.069536f
C631 VTAIL.n16 VSUBS 0.024275f
C632 VTAIL.n17 VSUBS 0.024348f
C633 VTAIL.n18 VSUBS 0.013693f
C634 VTAIL.n19 VSUBS 0.881224f
C635 VTAIL.n20 VSUBS 0.025483f
C636 VTAIL.n21 VSUBS 0.013693f
C637 VTAIL.n22 VSUBS 0.014499f
C638 VTAIL.n23 VSUBS 0.032367f
C639 VTAIL.n24 VSUBS 0.032367f
C640 VTAIL.n25 VSUBS 0.014499f
C641 VTAIL.n26 VSUBS 0.013693f
C642 VTAIL.n27 VSUBS 0.025483f
C643 VTAIL.n28 VSUBS 0.025483f
C644 VTAIL.n29 VSUBS 0.013693f
C645 VTAIL.n30 VSUBS 0.014499f
C646 VTAIL.n31 VSUBS 0.032367f
C647 VTAIL.n32 VSUBS 0.032367f
C648 VTAIL.n33 VSUBS 0.032367f
C649 VTAIL.n34 VSUBS 0.014499f
C650 VTAIL.n35 VSUBS 0.013693f
C651 VTAIL.n36 VSUBS 0.025483f
C652 VTAIL.n37 VSUBS 0.025483f
C653 VTAIL.n38 VSUBS 0.013693f
C654 VTAIL.n39 VSUBS 0.014096f
C655 VTAIL.n40 VSUBS 0.014096f
C656 VTAIL.n41 VSUBS 0.032367f
C657 VTAIL.n42 VSUBS 0.076521f
C658 VTAIL.n43 VSUBS 0.014499f
C659 VTAIL.n44 VSUBS 0.013693f
C660 VTAIL.n45 VSUBS 0.064473f
C661 VTAIL.n46 VSUBS 0.038565f
C662 VTAIL.n47 VSUBS 0.147022f
C663 VTAIL.n48 VSUBS 0.027462f
C664 VTAIL.n49 VSUBS 0.025483f
C665 VTAIL.n50 VSUBS 0.013693f
C666 VTAIL.n51 VSUBS 0.032367f
C667 VTAIL.n52 VSUBS 0.014499f
C668 VTAIL.n53 VSUBS 0.025483f
C669 VTAIL.n54 VSUBS 0.013693f
C670 VTAIL.n55 VSUBS 0.032367f
C671 VTAIL.n56 VSUBS 0.014499f
C672 VTAIL.n57 VSUBS 0.025483f
C673 VTAIL.n58 VSUBS 0.013693f
C674 VTAIL.n59 VSUBS 0.032367f
C675 VTAIL.n60 VSUBS 0.014499f
C676 VTAIL.n61 VSUBS 0.162504f
C677 VTAIL.t14 VSUBS 0.069536f
C678 VTAIL.n62 VSUBS 0.024275f
C679 VTAIL.n63 VSUBS 0.024348f
C680 VTAIL.n64 VSUBS 0.013693f
C681 VTAIL.n65 VSUBS 0.881224f
C682 VTAIL.n66 VSUBS 0.025483f
C683 VTAIL.n67 VSUBS 0.013693f
C684 VTAIL.n68 VSUBS 0.014499f
C685 VTAIL.n69 VSUBS 0.032367f
C686 VTAIL.n70 VSUBS 0.032367f
C687 VTAIL.n71 VSUBS 0.014499f
C688 VTAIL.n72 VSUBS 0.013693f
C689 VTAIL.n73 VSUBS 0.025483f
C690 VTAIL.n74 VSUBS 0.025483f
C691 VTAIL.n75 VSUBS 0.013693f
C692 VTAIL.n76 VSUBS 0.014499f
C693 VTAIL.n77 VSUBS 0.032367f
C694 VTAIL.n78 VSUBS 0.032367f
C695 VTAIL.n79 VSUBS 0.032367f
C696 VTAIL.n80 VSUBS 0.014499f
C697 VTAIL.n81 VSUBS 0.013693f
C698 VTAIL.n82 VSUBS 0.025483f
C699 VTAIL.n83 VSUBS 0.025483f
C700 VTAIL.n84 VSUBS 0.013693f
C701 VTAIL.n85 VSUBS 0.014096f
C702 VTAIL.n86 VSUBS 0.014096f
C703 VTAIL.n87 VSUBS 0.032367f
C704 VTAIL.n88 VSUBS 0.076521f
C705 VTAIL.n89 VSUBS 0.014499f
C706 VTAIL.n90 VSUBS 0.013693f
C707 VTAIL.n91 VSUBS 0.064473f
C708 VTAIL.n92 VSUBS 0.038565f
C709 VTAIL.n93 VSUBS 0.147022f
C710 VTAIL.t11 VSUBS 0.174794f
C711 VTAIL.t10 VSUBS 0.174794f
C712 VTAIL.n94 VSUBS 1.18219f
C713 VTAIL.n95 VSUBS 0.678266f
C714 VTAIL.n96 VSUBS 0.027462f
C715 VTAIL.n97 VSUBS 0.025483f
C716 VTAIL.n98 VSUBS 0.013693f
C717 VTAIL.n99 VSUBS 0.032367f
C718 VTAIL.n100 VSUBS 0.014499f
C719 VTAIL.n101 VSUBS 0.025483f
C720 VTAIL.n102 VSUBS 0.013693f
C721 VTAIL.n103 VSUBS 0.032367f
C722 VTAIL.n104 VSUBS 0.014499f
C723 VTAIL.n105 VSUBS 0.025483f
C724 VTAIL.n106 VSUBS 0.013693f
C725 VTAIL.n107 VSUBS 0.032367f
C726 VTAIL.n108 VSUBS 0.014499f
C727 VTAIL.n109 VSUBS 0.162504f
C728 VTAIL.t15 VSUBS 0.069536f
C729 VTAIL.n110 VSUBS 0.024275f
C730 VTAIL.n111 VSUBS 0.024348f
C731 VTAIL.n112 VSUBS 0.013693f
C732 VTAIL.n113 VSUBS 0.881224f
C733 VTAIL.n114 VSUBS 0.025483f
C734 VTAIL.n115 VSUBS 0.013693f
C735 VTAIL.n116 VSUBS 0.014499f
C736 VTAIL.n117 VSUBS 0.032367f
C737 VTAIL.n118 VSUBS 0.032367f
C738 VTAIL.n119 VSUBS 0.014499f
C739 VTAIL.n120 VSUBS 0.013693f
C740 VTAIL.n121 VSUBS 0.025483f
C741 VTAIL.n122 VSUBS 0.025483f
C742 VTAIL.n123 VSUBS 0.013693f
C743 VTAIL.n124 VSUBS 0.014499f
C744 VTAIL.n125 VSUBS 0.032367f
C745 VTAIL.n126 VSUBS 0.032367f
C746 VTAIL.n127 VSUBS 0.032367f
C747 VTAIL.n128 VSUBS 0.014499f
C748 VTAIL.n129 VSUBS 0.013693f
C749 VTAIL.n130 VSUBS 0.025483f
C750 VTAIL.n131 VSUBS 0.025483f
C751 VTAIL.n132 VSUBS 0.013693f
C752 VTAIL.n133 VSUBS 0.014096f
C753 VTAIL.n134 VSUBS 0.014096f
C754 VTAIL.n135 VSUBS 0.032367f
C755 VTAIL.n136 VSUBS 0.076521f
C756 VTAIL.n137 VSUBS 0.014499f
C757 VTAIL.n138 VSUBS 0.013693f
C758 VTAIL.n139 VSUBS 0.064473f
C759 VTAIL.n140 VSUBS 0.038565f
C760 VTAIL.n141 VSUBS 1.15256f
C761 VTAIL.n142 VSUBS 0.027462f
C762 VTAIL.n143 VSUBS 0.025483f
C763 VTAIL.n144 VSUBS 0.013693f
C764 VTAIL.n145 VSUBS 0.032367f
C765 VTAIL.n146 VSUBS 0.014499f
C766 VTAIL.n147 VSUBS 0.025483f
C767 VTAIL.n148 VSUBS 0.013693f
C768 VTAIL.n149 VSUBS 0.032367f
C769 VTAIL.n150 VSUBS 0.032367f
C770 VTAIL.n151 VSUBS 0.014499f
C771 VTAIL.n152 VSUBS 0.025483f
C772 VTAIL.n153 VSUBS 0.013693f
C773 VTAIL.n154 VSUBS 0.032367f
C774 VTAIL.n155 VSUBS 0.014499f
C775 VTAIL.n156 VSUBS 0.162504f
C776 VTAIL.t1 VSUBS 0.069536f
C777 VTAIL.n157 VSUBS 0.024275f
C778 VTAIL.n158 VSUBS 0.024348f
C779 VTAIL.n159 VSUBS 0.013693f
C780 VTAIL.n160 VSUBS 0.881224f
C781 VTAIL.n161 VSUBS 0.025483f
C782 VTAIL.n162 VSUBS 0.013693f
C783 VTAIL.n163 VSUBS 0.014499f
C784 VTAIL.n164 VSUBS 0.032367f
C785 VTAIL.n165 VSUBS 0.032367f
C786 VTAIL.n166 VSUBS 0.014499f
C787 VTAIL.n167 VSUBS 0.013693f
C788 VTAIL.n168 VSUBS 0.025483f
C789 VTAIL.n169 VSUBS 0.025483f
C790 VTAIL.n170 VSUBS 0.013693f
C791 VTAIL.n171 VSUBS 0.014499f
C792 VTAIL.n172 VSUBS 0.032367f
C793 VTAIL.n173 VSUBS 0.032367f
C794 VTAIL.n174 VSUBS 0.014499f
C795 VTAIL.n175 VSUBS 0.013693f
C796 VTAIL.n176 VSUBS 0.025483f
C797 VTAIL.n177 VSUBS 0.025483f
C798 VTAIL.n178 VSUBS 0.013693f
C799 VTAIL.n179 VSUBS 0.014096f
C800 VTAIL.n180 VSUBS 0.014096f
C801 VTAIL.n181 VSUBS 0.032367f
C802 VTAIL.n182 VSUBS 0.076521f
C803 VTAIL.n183 VSUBS 0.014499f
C804 VTAIL.n184 VSUBS 0.013693f
C805 VTAIL.n185 VSUBS 0.064473f
C806 VTAIL.n186 VSUBS 0.038565f
C807 VTAIL.n187 VSUBS 1.15256f
C808 VTAIL.t7 VSUBS 0.174794f
C809 VTAIL.t6 VSUBS 0.174794f
C810 VTAIL.n188 VSUBS 1.18219f
C811 VTAIL.n189 VSUBS 0.678258f
C812 VTAIL.n190 VSUBS 0.027462f
C813 VTAIL.n191 VSUBS 0.025483f
C814 VTAIL.n192 VSUBS 0.013693f
C815 VTAIL.n193 VSUBS 0.032367f
C816 VTAIL.n194 VSUBS 0.014499f
C817 VTAIL.n195 VSUBS 0.025483f
C818 VTAIL.n196 VSUBS 0.013693f
C819 VTAIL.n197 VSUBS 0.032367f
C820 VTAIL.n198 VSUBS 0.032367f
C821 VTAIL.n199 VSUBS 0.014499f
C822 VTAIL.n200 VSUBS 0.025483f
C823 VTAIL.n201 VSUBS 0.013693f
C824 VTAIL.n202 VSUBS 0.032367f
C825 VTAIL.n203 VSUBS 0.014499f
C826 VTAIL.n204 VSUBS 0.162504f
C827 VTAIL.t0 VSUBS 0.069536f
C828 VTAIL.n205 VSUBS 0.024275f
C829 VTAIL.n206 VSUBS 0.024348f
C830 VTAIL.n207 VSUBS 0.013693f
C831 VTAIL.n208 VSUBS 0.881224f
C832 VTAIL.n209 VSUBS 0.025483f
C833 VTAIL.n210 VSUBS 0.013693f
C834 VTAIL.n211 VSUBS 0.014499f
C835 VTAIL.n212 VSUBS 0.032367f
C836 VTAIL.n213 VSUBS 0.032367f
C837 VTAIL.n214 VSUBS 0.014499f
C838 VTAIL.n215 VSUBS 0.013693f
C839 VTAIL.n216 VSUBS 0.025483f
C840 VTAIL.n217 VSUBS 0.025483f
C841 VTAIL.n218 VSUBS 0.013693f
C842 VTAIL.n219 VSUBS 0.014499f
C843 VTAIL.n220 VSUBS 0.032367f
C844 VTAIL.n221 VSUBS 0.032367f
C845 VTAIL.n222 VSUBS 0.014499f
C846 VTAIL.n223 VSUBS 0.013693f
C847 VTAIL.n224 VSUBS 0.025483f
C848 VTAIL.n225 VSUBS 0.025483f
C849 VTAIL.n226 VSUBS 0.013693f
C850 VTAIL.n227 VSUBS 0.014096f
C851 VTAIL.n228 VSUBS 0.014096f
C852 VTAIL.n229 VSUBS 0.032367f
C853 VTAIL.n230 VSUBS 0.076521f
C854 VTAIL.n231 VSUBS 0.014499f
C855 VTAIL.n232 VSUBS 0.013693f
C856 VTAIL.n233 VSUBS 0.064473f
C857 VTAIL.n234 VSUBS 0.038565f
C858 VTAIL.n235 VSUBS 0.147022f
C859 VTAIL.n236 VSUBS 0.027462f
C860 VTAIL.n237 VSUBS 0.025483f
C861 VTAIL.n238 VSUBS 0.013693f
C862 VTAIL.n239 VSUBS 0.032367f
C863 VTAIL.n240 VSUBS 0.014499f
C864 VTAIL.n241 VSUBS 0.025483f
C865 VTAIL.n242 VSUBS 0.013693f
C866 VTAIL.n243 VSUBS 0.032367f
C867 VTAIL.n244 VSUBS 0.032367f
C868 VTAIL.n245 VSUBS 0.014499f
C869 VTAIL.n246 VSUBS 0.025483f
C870 VTAIL.n247 VSUBS 0.013693f
C871 VTAIL.n248 VSUBS 0.032367f
C872 VTAIL.n249 VSUBS 0.014499f
C873 VTAIL.n250 VSUBS 0.162504f
C874 VTAIL.t12 VSUBS 0.069536f
C875 VTAIL.n251 VSUBS 0.024275f
C876 VTAIL.n252 VSUBS 0.024348f
C877 VTAIL.n253 VSUBS 0.013693f
C878 VTAIL.n254 VSUBS 0.881224f
C879 VTAIL.n255 VSUBS 0.025483f
C880 VTAIL.n256 VSUBS 0.013693f
C881 VTAIL.n257 VSUBS 0.014499f
C882 VTAIL.n258 VSUBS 0.032367f
C883 VTAIL.n259 VSUBS 0.032367f
C884 VTAIL.n260 VSUBS 0.014499f
C885 VTAIL.n261 VSUBS 0.013693f
C886 VTAIL.n262 VSUBS 0.025483f
C887 VTAIL.n263 VSUBS 0.025483f
C888 VTAIL.n264 VSUBS 0.013693f
C889 VTAIL.n265 VSUBS 0.014499f
C890 VTAIL.n266 VSUBS 0.032367f
C891 VTAIL.n267 VSUBS 0.032367f
C892 VTAIL.n268 VSUBS 0.014499f
C893 VTAIL.n269 VSUBS 0.013693f
C894 VTAIL.n270 VSUBS 0.025483f
C895 VTAIL.n271 VSUBS 0.025483f
C896 VTAIL.n272 VSUBS 0.013693f
C897 VTAIL.n273 VSUBS 0.014096f
C898 VTAIL.n274 VSUBS 0.014096f
C899 VTAIL.n275 VSUBS 0.032367f
C900 VTAIL.n276 VSUBS 0.076521f
C901 VTAIL.n277 VSUBS 0.014499f
C902 VTAIL.n278 VSUBS 0.013693f
C903 VTAIL.n279 VSUBS 0.064473f
C904 VTAIL.n280 VSUBS 0.038565f
C905 VTAIL.n281 VSUBS 0.147022f
C906 VTAIL.t9 VSUBS 0.174794f
C907 VTAIL.t8 VSUBS 0.174794f
C908 VTAIL.n282 VSUBS 1.18219f
C909 VTAIL.n283 VSUBS 0.678258f
C910 VTAIL.n284 VSUBS 0.027462f
C911 VTAIL.n285 VSUBS 0.025483f
C912 VTAIL.n286 VSUBS 0.013693f
C913 VTAIL.n287 VSUBS 0.032367f
C914 VTAIL.n288 VSUBS 0.014499f
C915 VTAIL.n289 VSUBS 0.025483f
C916 VTAIL.n290 VSUBS 0.013693f
C917 VTAIL.n291 VSUBS 0.032367f
C918 VTAIL.n292 VSUBS 0.032367f
C919 VTAIL.n293 VSUBS 0.014499f
C920 VTAIL.n294 VSUBS 0.025483f
C921 VTAIL.n295 VSUBS 0.013693f
C922 VTAIL.n296 VSUBS 0.032367f
C923 VTAIL.n297 VSUBS 0.014499f
C924 VTAIL.n298 VSUBS 0.162504f
C925 VTAIL.t13 VSUBS 0.069536f
C926 VTAIL.n299 VSUBS 0.024275f
C927 VTAIL.n300 VSUBS 0.024348f
C928 VTAIL.n301 VSUBS 0.013693f
C929 VTAIL.n302 VSUBS 0.881224f
C930 VTAIL.n303 VSUBS 0.025483f
C931 VTAIL.n304 VSUBS 0.013693f
C932 VTAIL.n305 VSUBS 0.014499f
C933 VTAIL.n306 VSUBS 0.032367f
C934 VTAIL.n307 VSUBS 0.032367f
C935 VTAIL.n308 VSUBS 0.014499f
C936 VTAIL.n309 VSUBS 0.013693f
C937 VTAIL.n310 VSUBS 0.025483f
C938 VTAIL.n311 VSUBS 0.025483f
C939 VTAIL.n312 VSUBS 0.013693f
C940 VTAIL.n313 VSUBS 0.014499f
C941 VTAIL.n314 VSUBS 0.032367f
C942 VTAIL.n315 VSUBS 0.032367f
C943 VTAIL.n316 VSUBS 0.014499f
C944 VTAIL.n317 VSUBS 0.013693f
C945 VTAIL.n318 VSUBS 0.025483f
C946 VTAIL.n319 VSUBS 0.025483f
C947 VTAIL.n320 VSUBS 0.013693f
C948 VTAIL.n321 VSUBS 0.014096f
C949 VTAIL.n322 VSUBS 0.014096f
C950 VTAIL.n323 VSUBS 0.032367f
C951 VTAIL.n324 VSUBS 0.076521f
C952 VTAIL.n325 VSUBS 0.014499f
C953 VTAIL.n326 VSUBS 0.013693f
C954 VTAIL.n327 VSUBS 0.064473f
C955 VTAIL.n328 VSUBS 0.038565f
C956 VTAIL.n329 VSUBS 1.15256f
C957 VTAIL.n330 VSUBS 0.027462f
C958 VTAIL.n331 VSUBS 0.025483f
C959 VTAIL.n332 VSUBS 0.013693f
C960 VTAIL.n333 VSUBS 0.032367f
C961 VTAIL.n334 VSUBS 0.014499f
C962 VTAIL.n335 VSUBS 0.025483f
C963 VTAIL.n336 VSUBS 0.013693f
C964 VTAIL.n337 VSUBS 0.032367f
C965 VTAIL.n338 VSUBS 0.014499f
C966 VTAIL.n339 VSUBS 0.025483f
C967 VTAIL.n340 VSUBS 0.013693f
C968 VTAIL.n341 VSUBS 0.032367f
C969 VTAIL.n342 VSUBS 0.014499f
C970 VTAIL.n343 VSUBS 0.162504f
C971 VTAIL.t2 VSUBS 0.069536f
C972 VTAIL.n344 VSUBS 0.024275f
C973 VTAIL.n345 VSUBS 0.024348f
C974 VTAIL.n346 VSUBS 0.013693f
C975 VTAIL.n347 VSUBS 0.881224f
C976 VTAIL.n348 VSUBS 0.025483f
C977 VTAIL.n349 VSUBS 0.013693f
C978 VTAIL.n350 VSUBS 0.014499f
C979 VTAIL.n351 VSUBS 0.032367f
C980 VTAIL.n352 VSUBS 0.032367f
C981 VTAIL.n353 VSUBS 0.014499f
C982 VTAIL.n354 VSUBS 0.013693f
C983 VTAIL.n355 VSUBS 0.025483f
C984 VTAIL.n356 VSUBS 0.025483f
C985 VTAIL.n357 VSUBS 0.013693f
C986 VTAIL.n358 VSUBS 0.014499f
C987 VTAIL.n359 VSUBS 0.032367f
C988 VTAIL.n360 VSUBS 0.032367f
C989 VTAIL.n361 VSUBS 0.032367f
C990 VTAIL.n362 VSUBS 0.014499f
C991 VTAIL.n363 VSUBS 0.013693f
C992 VTAIL.n364 VSUBS 0.025483f
C993 VTAIL.n365 VSUBS 0.025483f
C994 VTAIL.n366 VSUBS 0.013693f
C995 VTAIL.n367 VSUBS 0.014096f
C996 VTAIL.n368 VSUBS 0.014096f
C997 VTAIL.n369 VSUBS 0.032367f
C998 VTAIL.n370 VSUBS 0.076521f
C999 VTAIL.n371 VSUBS 0.014499f
C1000 VTAIL.n372 VSUBS 0.013693f
C1001 VTAIL.n373 VSUBS 0.064473f
C1002 VTAIL.n374 VSUBS 0.038565f
C1003 VTAIL.n375 VSUBS 1.14778f
C1004 VP.n0 VSUBS 0.054201f
C1005 VP.t2 VSUBS 1.07767f
C1006 VP.n1 VSUBS 0.423188f
C1007 VP.n2 VSUBS 0.054201f
C1008 VP.t4 VSUBS 1.07767f
C1009 VP.n3 VSUBS 0.021699f
C1010 VP.n4 VSUBS 0.054201f
C1011 VP.t6 VSUBS 1.14782f
C1012 VP.t7 VSUBS 1.07767f
C1013 VP.n5 VSUBS 0.423188f
C1014 VP.n6 VSUBS 0.22869f
C1015 VP.t1 VSUBS 1.07767f
C1016 VP.t3 VSUBS 1.18059f
C1017 VP.n7 VSUBS 0.478803f
C1018 VP.n8 VSUBS 0.479233f
C1019 VP.n9 VSUBS 0.062912f
C1020 VP.n10 VSUBS 0.062912f
C1021 VP.n11 VSUBS 0.054201f
C1022 VP.n12 VSUBS 0.054201f
C1023 VP.n13 VSUBS 0.068201f
C1024 VP.n14 VSUBS 0.021699f
C1025 VP.n15 VSUBS 0.476571f
C1026 VP.n16 VSUBS 2.07714f
C1027 VP.t5 VSUBS 1.14782f
C1028 VP.n17 VSUBS 0.476571f
C1029 VP.n18 VSUBS 2.12575f
C1030 VP.n19 VSUBS 0.054201f
C1031 VP.n20 VSUBS 0.054201f
C1032 VP.n21 VSUBS 0.068201f
C1033 VP.n22 VSUBS 0.423188f
C1034 VP.n23 VSUBS 0.062912f
C1035 VP.n24 VSUBS 0.062912f
C1036 VP.n25 VSUBS 0.054201f
C1037 VP.n26 VSUBS 0.054201f
C1038 VP.n27 VSUBS 0.068201f
C1039 VP.n28 VSUBS 0.021699f
C1040 VP.t0 VSUBS 1.14782f
C1041 VP.n29 VSUBS 0.476571f
C1042 VP.n30 VSUBS 0.042004f
.ends

