* NGSPICE file created from diff_pair_sample_1526.ext - technology: sky130A

.subckt diff_pair_sample_1526 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t7 VN.t0 VTAIL.t7 B.t1 sky130_fd_pr__nfet_01v8 ad=0.60555 pd=4 as=0.60555 ps=4 w=3.67 l=2.56
X1 VTAIL.t3 VP.t0 VDD1.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=1.4313 pd=8.12 as=0.60555 ps=4 w=3.67 l=2.56
X2 VTAIL.t4 VP.t1 VDD1.t6 B.t4 sky130_fd_pr__nfet_01v8 ad=0.60555 pd=4 as=0.60555 ps=4 w=3.67 l=2.56
X3 VDD2.t6 VN.t1 VTAIL.t11 B.t2 sky130_fd_pr__nfet_01v8 ad=0.60555 pd=4 as=0.60555 ps=4 w=3.67 l=2.56
X4 B.t19 B.t17 B.t18 B.t14 sky130_fd_pr__nfet_01v8 ad=1.4313 pd=8.12 as=0 ps=0 w=3.67 l=2.56
X5 B.t16 B.t13 B.t15 B.t14 sky130_fd_pr__nfet_01v8 ad=1.4313 pd=8.12 as=0 ps=0 w=3.67 l=2.56
X6 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=1.4313 pd=8.12 as=0 ps=0 w=3.67 l=2.56
X7 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=1.4313 pd=8.12 as=0 ps=0 w=3.67 l=2.56
X8 VDD1.t5 VP.t2 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.60555 pd=4 as=0.60555 ps=4 w=3.67 l=2.56
X9 VDD1.t4 VP.t3 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.60555 pd=4 as=0.60555 ps=4 w=3.67 l=2.56
X10 VTAIL.t12 VN.t2 VDD2.t5 B.t3 sky130_fd_pr__nfet_01v8 ad=1.4313 pd=8.12 as=0.60555 ps=4 w=3.67 l=2.56
X11 VDD1.t3 VP.t4 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.60555 pd=4 as=1.4313 ps=8.12 w=3.67 l=2.56
X12 VTAIL.t13 VN.t3 VDD2.t4 B.t20 sky130_fd_pr__nfet_01v8 ad=1.4313 pd=8.12 as=0.60555 ps=4 w=3.67 l=2.56
X13 VDD2.t3 VN.t4 VTAIL.t14 B.t0 sky130_fd_pr__nfet_01v8 ad=0.60555 pd=4 as=1.4313 ps=8.12 w=3.67 l=2.56
X14 VDD1.t2 VP.t5 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=0.60555 pd=4 as=1.4313 ps=8.12 w=3.67 l=2.56
X15 VTAIL.t15 VP.t6 VDD1.t1 B.t21 sky130_fd_pr__nfet_01v8 ad=0.60555 pd=4 as=0.60555 ps=4 w=3.67 l=2.56
X16 VTAIL.t8 VN.t5 VDD2.t2 B.t21 sky130_fd_pr__nfet_01v8 ad=0.60555 pd=4 as=0.60555 ps=4 w=3.67 l=2.56
X17 VTAIL.t6 VP.t7 VDD1.t0 B.t20 sky130_fd_pr__nfet_01v8 ad=1.4313 pd=8.12 as=0.60555 ps=4 w=3.67 l=2.56
X18 VDD2.t1 VN.t6 VTAIL.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=0.60555 pd=4 as=1.4313 ps=8.12 w=3.67 l=2.56
X19 VTAIL.t10 VN.t7 VDD2.t0 B.t4 sky130_fd_pr__nfet_01v8 ad=0.60555 pd=4 as=0.60555 ps=4 w=3.67 l=2.56
R0 VN.n55 VN.n29 161.3
R1 VN.n54 VN.n53 161.3
R2 VN.n52 VN.n30 161.3
R3 VN.n51 VN.n50 161.3
R4 VN.n49 VN.n31 161.3
R5 VN.n48 VN.n47 161.3
R6 VN.n46 VN.n45 161.3
R7 VN.n44 VN.n33 161.3
R8 VN.n43 VN.n42 161.3
R9 VN.n41 VN.n34 161.3
R10 VN.n40 VN.n39 161.3
R11 VN.n38 VN.n35 161.3
R12 VN.n26 VN.n0 161.3
R13 VN.n25 VN.n24 161.3
R14 VN.n23 VN.n1 161.3
R15 VN.n22 VN.n21 161.3
R16 VN.n20 VN.n2 161.3
R17 VN.n19 VN.n18 161.3
R18 VN.n17 VN.n16 161.3
R19 VN.n15 VN.n4 161.3
R20 VN.n14 VN.n13 161.3
R21 VN.n12 VN.n5 161.3
R22 VN.n11 VN.n10 161.3
R23 VN.n9 VN.n6 161.3
R24 VN.n28 VN.n27 106.597
R25 VN.n57 VN.n56 106.597
R26 VN.n7 VN.t2 66.272
R27 VN.n36 VN.t4 66.272
R28 VN.n8 VN.n7 62.8231
R29 VN.n37 VN.n36 62.8231
R30 VN.n14 VN.n5 56.5193
R31 VN.n43 VN.n34 56.5193
R32 VN.n21 VN.n1 54.0911
R33 VN.n50 VN.n30 54.0911
R34 VN VN.n57 44.5966
R35 VN.n8 VN.t0 34.5501
R36 VN.n3 VN.t5 34.5501
R37 VN.n27 VN.t6 34.5501
R38 VN.n37 VN.t7 34.5501
R39 VN.n32 VN.t1 34.5501
R40 VN.n56 VN.t3 34.5501
R41 VN.n21 VN.n20 26.8957
R42 VN.n50 VN.n49 26.8957
R43 VN.n10 VN.n9 24.4675
R44 VN.n10 VN.n5 24.4675
R45 VN.n15 VN.n14 24.4675
R46 VN.n16 VN.n15 24.4675
R47 VN.n20 VN.n19 24.4675
R48 VN.n25 VN.n1 24.4675
R49 VN.n26 VN.n25 24.4675
R50 VN.n39 VN.n34 24.4675
R51 VN.n39 VN.n38 24.4675
R52 VN.n49 VN.n48 24.4675
R53 VN.n45 VN.n44 24.4675
R54 VN.n44 VN.n43 24.4675
R55 VN.n55 VN.n54 24.4675
R56 VN.n54 VN.n30 24.4675
R57 VN.n19 VN.n3 14.9254
R58 VN.n48 VN.n32 14.9254
R59 VN.n9 VN.n8 9.54263
R60 VN.n16 VN.n3 9.54263
R61 VN.n38 VN.n37 9.54263
R62 VN.n45 VN.n32 9.54263
R63 VN.n36 VN.n35 7.21701
R64 VN.n7 VN.n6 7.21701
R65 VN.n27 VN.n26 4.15989
R66 VN.n56 VN.n55 4.15989
R67 VN.n57 VN.n29 0.278367
R68 VN.n28 VN.n0 0.278367
R69 VN.n53 VN.n29 0.189894
R70 VN.n53 VN.n52 0.189894
R71 VN.n52 VN.n51 0.189894
R72 VN.n51 VN.n31 0.189894
R73 VN.n47 VN.n31 0.189894
R74 VN.n47 VN.n46 0.189894
R75 VN.n46 VN.n33 0.189894
R76 VN.n42 VN.n33 0.189894
R77 VN.n42 VN.n41 0.189894
R78 VN.n41 VN.n40 0.189894
R79 VN.n40 VN.n35 0.189894
R80 VN.n11 VN.n6 0.189894
R81 VN.n12 VN.n11 0.189894
R82 VN.n13 VN.n12 0.189894
R83 VN.n13 VN.n4 0.189894
R84 VN.n17 VN.n4 0.189894
R85 VN.n18 VN.n17 0.189894
R86 VN.n18 VN.n2 0.189894
R87 VN.n22 VN.n2 0.189894
R88 VN.n23 VN.n22 0.189894
R89 VN.n24 VN.n23 0.189894
R90 VN.n24 VN.n0 0.189894
R91 VN VN.n28 0.153454
R92 VTAIL.n11 VTAIL.t3 67.7617
R93 VTAIL.n10 VTAIL.t14 67.7617
R94 VTAIL.n7 VTAIL.t13 67.7617
R95 VTAIL.n15 VTAIL.t9 67.7617
R96 VTAIL.n2 VTAIL.t12 67.7617
R97 VTAIL.n3 VTAIL.t0 67.7617
R98 VTAIL.n6 VTAIL.t6 67.7617
R99 VTAIL.n14 VTAIL.t5 67.7617
R100 VTAIL.n13 VTAIL.n12 62.3667
R101 VTAIL.n9 VTAIL.n8 62.3667
R102 VTAIL.n1 VTAIL.n0 62.3665
R103 VTAIL.n5 VTAIL.n4 62.3665
R104 VTAIL.n15 VTAIL.n14 18.0221
R105 VTAIL.n7 VTAIL.n6 18.0221
R106 VTAIL.n0 VTAIL.t7 5.3956
R107 VTAIL.n0 VTAIL.t8 5.3956
R108 VTAIL.n4 VTAIL.t2 5.3956
R109 VTAIL.n4 VTAIL.t4 5.3956
R110 VTAIL.n12 VTAIL.t1 5.3956
R111 VTAIL.n12 VTAIL.t15 5.3956
R112 VTAIL.n8 VTAIL.t11 5.3956
R113 VTAIL.n8 VTAIL.t10 5.3956
R114 VTAIL.n9 VTAIL.n7 2.49188
R115 VTAIL.n10 VTAIL.n9 2.49188
R116 VTAIL.n13 VTAIL.n11 2.49188
R117 VTAIL.n14 VTAIL.n13 2.49188
R118 VTAIL.n6 VTAIL.n5 2.49188
R119 VTAIL.n5 VTAIL.n3 2.49188
R120 VTAIL.n2 VTAIL.n1 2.49188
R121 VTAIL VTAIL.n15 2.43369
R122 VTAIL.n11 VTAIL.n10 0.470328
R123 VTAIL.n3 VTAIL.n2 0.470328
R124 VTAIL VTAIL.n1 0.0586897
R125 VDD2.n2 VDD2.n1 80.2356
R126 VDD2.n2 VDD2.n0 80.2356
R127 VDD2 VDD2.n5 80.2329
R128 VDD2.n4 VDD2.n3 79.0455
R129 VDD2.n4 VDD2.n2 38.0903
R130 VDD2.n5 VDD2.t0 5.3956
R131 VDD2.n5 VDD2.t3 5.3956
R132 VDD2.n3 VDD2.t4 5.3956
R133 VDD2.n3 VDD2.t6 5.3956
R134 VDD2.n1 VDD2.t2 5.3956
R135 VDD2.n1 VDD2.t1 5.3956
R136 VDD2.n0 VDD2.t5 5.3956
R137 VDD2.n0 VDD2.t7 5.3956
R138 VDD2 VDD2.n4 1.30438
R139 B.n550 B.n549 585
R140 B.n552 B.n120 585
R141 B.n555 B.n554 585
R142 B.n556 B.n119 585
R143 B.n558 B.n557 585
R144 B.n560 B.n118 585
R145 B.n563 B.n562 585
R146 B.n564 B.n117 585
R147 B.n566 B.n565 585
R148 B.n568 B.n116 585
R149 B.n571 B.n570 585
R150 B.n572 B.n115 585
R151 B.n574 B.n573 585
R152 B.n576 B.n114 585
R153 B.n579 B.n578 585
R154 B.n580 B.n110 585
R155 B.n582 B.n581 585
R156 B.n584 B.n109 585
R157 B.n587 B.n586 585
R158 B.n588 B.n108 585
R159 B.n590 B.n589 585
R160 B.n592 B.n107 585
R161 B.n595 B.n594 585
R162 B.n596 B.n106 585
R163 B.n598 B.n597 585
R164 B.n600 B.n105 585
R165 B.n603 B.n602 585
R166 B.n605 B.n102 585
R167 B.n607 B.n606 585
R168 B.n609 B.n101 585
R169 B.n612 B.n611 585
R170 B.n613 B.n100 585
R171 B.n615 B.n614 585
R172 B.n617 B.n99 585
R173 B.n620 B.n619 585
R174 B.n621 B.n98 585
R175 B.n623 B.n622 585
R176 B.n625 B.n97 585
R177 B.n628 B.n627 585
R178 B.n629 B.n96 585
R179 B.n631 B.n630 585
R180 B.n633 B.n95 585
R181 B.n636 B.n635 585
R182 B.n637 B.n94 585
R183 B.n548 B.n92 585
R184 B.n640 B.n92 585
R185 B.n547 B.n91 585
R186 B.n641 B.n91 585
R187 B.n546 B.n90 585
R188 B.n642 B.n90 585
R189 B.n545 B.n544 585
R190 B.n544 B.n86 585
R191 B.n543 B.n85 585
R192 B.n648 B.n85 585
R193 B.n542 B.n84 585
R194 B.n649 B.n84 585
R195 B.n541 B.n83 585
R196 B.n650 B.n83 585
R197 B.n540 B.n539 585
R198 B.n539 B.n82 585
R199 B.n538 B.n78 585
R200 B.n656 B.n78 585
R201 B.n537 B.n77 585
R202 B.n657 B.n77 585
R203 B.n536 B.n76 585
R204 B.n658 B.n76 585
R205 B.n535 B.n534 585
R206 B.n534 B.n72 585
R207 B.n533 B.n71 585
R208 B.n664 B.n71 585
R209 B.n532 B.n70 585
R210 B.n665 B.n70 585
R211 B.n531 B.n69 585
R212 B.n666 B.n69 585
R213 B.n530 B.n529 585
R214 B.n529 B.n65 585
R215 B.n528 B.n64 585
R216 B.n672 B.n64 585
R217 B.n527 B.n63 585
R218 B.n673 B.n63 585
R219 B.n526 B.n62 585
R220 B.n674 B.n62 585
R221 B.n525 B.n524 585
R222 B.n524 B.n61 585
R223 B.n523 B.n57 585
R224 B.n680 B.n57 585
R225 B.n522 B.n56 585
R226 B.n681 B.n56 585
R227 B.n521 B.n55 585
R228 B.n682 B.n55 585
R229 B.n520 B.n519 585
R230 B.n519 B.n51 585
R231 B.n518 B.n50 585
R232 B.n688 B.n50 585
R233 B.n517 B.n49 585
R234 B.n689 B.n49 585
R235 B.n516 B.n48 585
R236 B.n690 B.n48 585
R237 B.n515 B.n514 585
R238 B.n514 B.n47 585
R239 B.n513 B.n43 585
R240 B.n696 B.n43 585
R241 B.n512 B.n42 585
R242 B.n697 B.n42 585
R243 B.n511 B.n41 585
R244 B.n698 B.n41 585
R245 B.n510 B.n509 585
R246 B.n509 B.n37 585
R247 B.n508 B.n36 585
R248 B.n704 B.n36 585
R249 B.n507 B.n35 585
R250 B.n705 B.n35 585
R251 B.n506 B.n34 585
R252 B.n706 B.n34 585
R253 B.n505 B.n504 585
R254 B.n504 B.n30 585
R255 B.n503 B.n29 585
R256 B.n712 B.n29 585
R257 B.n502 B.n28 585
R258 B.n713 B.n28 585
R259 B.n501 B.n27 585
R260 B.n714 B.n27 585
R261 B.n500 B.n499 585
R262 B.n499 B.n23 585
R263 B.n498 B.n22 585
R264 B.n720 B.n22 585
R265 B.n497 B.n21 585
R266 B.n721 B.n21 585
R267 B.n496 B.n20 585
R268 B.n722 B.n20 585
R269 B.n495 B.n494 585
R270 B.n494 B.n16 585
R271 B.n493 B.n15 585
R272 B.n728 B.n15 585
R273 B.n492 B.n14 585
R274 B.n729 B.n14 585
R275 B.n491 B.n13 585
R276 B.n730 B.n13 585
R277 B.n490 B.n489 585
R278 B.n489 B.n12 585
R279 B.n488 B.n487 585
R280 B.n488 B.n8 585
R281 B.n486 B.n7 585
R282 B.n737 B.n7 585
R283 B.n485 B.n6 585
R284 B.n738 B.n6 585
R285 B.n484 B.n5 585
R286 B.n739 B.n5 585
R287 B.n483 B.n482 585
R288 B.n482 B.n4 585
R289 B.n481 B.n121 585
R290 B.n481 B.n480 585
R291 B.n471 B.n122 585
R292 B.n123 B.n122 585
R293 B.n473 B.n472 585
R294 B.n474 B.n473 585
R295 B.n470 B.n128 585
R296 B.n128 B.n127 585
R297 B.n469 B.n468 585
R298 B.n468 B.n467 585
R299 B.n130 B.n129 585
R300 B.n131 B.n130 585
R301 B.n460 B.n459 585
R302 B.n461 B.n460 585
R303 B.n458 B.n136 585
R304 B.n136 B.n135 585
R305 B.n457 B.n456 585
R306 B.n456 B.n455 585
R307 B.n138 B.n137 585
R308 B.n139 B.n138 585
R309 B.n448 B.n447 585
R310 B.n449 B.n448 585
R311 B.n446 B.n144 585
R312 B.n144 B.n143 585
R313 B.n445 B.n444 585
R314 B.n444 B.n443 585
R315 B.n146 B.n145 585
R316 B.n147 B.n146 585
R317 B.n436 B.n435 585
R318 B.n437 B.n436 585
R319 B.n434 B.n152 585
R320 B.n152 B.n151 585
R321 B.n433 B.n432 585
R322 B.n432 B.n431 585
R323 B.n154 B.n153 585
R324 B.n155 B.n154 585
R325 B.n424 B.n423 585
R326 B.n425 B.n424 585
R327 B.n422 B.n160 585
R328 B.n160 B.n159 585
R329 B.n421 B.n420 585
R330 B.n420 B.n419 585
R331 B.n162 B.n161 585
R332 B.n412 B.n162 585
R333 B.n411 B.n410 585
R334 B.n413 B.n411 585
R335 B.n409 B.n167 585
R336 B.n167 B.n166 585
R337 B.n408 B.n407 585
R338 B.n407 B.n406 585
R339 B.n169 B.n168 585
R340 B.n170 B.n169 585
R341 B.n399 B.n398 585
R342 B.n400 B.n399 585
R343 B.n397 B.n175 585
R344 B.n175 B.n174 585
R345 B.n396 B.n395 585
R346 B.n395 B.n394 585
R347 B.n177 B.n176 585
R348 B.n387 B.n177 585
R349 B.n386 B.n385 585
R350 B.n388 B.n386 585
R351 B.n384 B.n182 585
R352 B.n182 B.n181 585
R353 B.n383 B.n382 585
R354 B.n382 B.n381 585
R355 B.n184 B.n183 585
R356 B.n185 B.n184 585
R357 B.n374 B.n373 585
R358 B.n375 B.n374 585
R359 B.n372 B.n190 585
R360 B.n190 B.n189 585
R361 B.n371 B.n370 585
R362 B.n370 B.n369 585
R363 B.n192 B.n191 585
R364 B.n193 B.n192 585
R365 B.n362 B.n361 585
R366 B.n363 B.n362 585
R367 B.n360 B.n198 585
R368 B.n198 B.n197 585
R369 B.n359 B.n358 585
R370 B.n358 B.n357 585
R371 B.n200 B.n199 585
R372 B.n350 B.n200 585
R373 B.n349 B.n348 585
R374 B.n351 B.n349 585
R375 B.n347 B.n205 585
R376 B.n205 B.n204 585
R377 B.n346 B.n345 585
R378 B.n345 B.n344 585
R379 B.n207 B.n206 585
R380 B.n208 B.n207 585
R381 B.n337 B.n336 585
R382 B.n338 B.n337 585
R383 B.n335 B.n213 585
R384 B.n213 B.n212 585
R385 B.n334 B.n333 585
R386 B.n333 B.n332 585
R387 B.n329 B.n217 585
R388 B.n328 B.n327 585
R389 B.n325 B.n218 585
R390 B.n325 B.n216 585
R391 B.n324 B.n323 585
R392 B.n322 B.n321 585
R393 B.n320 B.n220 585
R394 B.n318 B.n317 585
R395 B.n316 B.n221 585
R396 B.n315 B.n314 585
R397 B.n312 B.n222 585
R398 B.n310 B.n309 585
R399 B.n308 B.n223 585
R400 B.n307 B.n306 585
R401 B.n304 B.n224 585
R402 B.n302 B.n301 585
R403 B.n300 B.n225 585
R404 B.n299 B.n298 585
R405 B.n296 B.n295 585
R406 B.n294 B.n293 585
R407 B.n292 B.n230 585
R408 B.n290 B.n289 585
R409 B.n288 B.n231 585
R410 B.n287 B.n286 585
R411 B.n284 B.n232 585
R412 B.n282 B.n281 585
R413 B.n280 B.n233 585
R414 B.n279 B.n278 585
R415 B.n276 B.n275 585
R416 B.n274 B.n273 585
R417 B.n272 B.n238 585
R418 B.n270 B.n269 585
R419 B.n268 B.n239 585
R420 B.n267 B.n266 585
R421 B.n264 B.n240 585
R422 B.n262 B.n261 585
R423 B.n260 B.n241 585
R424 B.n259 B.n258 585
R425 B.n256 B.n242 585
R426 B.n254 B.n253 585
R427 B.n252 B.n243 585
R428 B.n251 B.n250 585
R429 B.n248 B.n244 585
R430 B.n246 B.n245 585
R431 B.n215 B.n214 585
R432 B.n216 B.n215 585
R433 B.n331 B.n330 585
R434 B.n332 B.n331 585
R435 B.n211 B.n210 585
R436 B.n212 B.n211 585
R437 B.n340 B.n339 585
R438 B.n339 B.n338 585
R439 B.n341 B.n209 585
R440 B.n209 B.n208 585
R441 B.n343 B.n342 585
R442 B.n344 B.n343 585
R443 B.n203 B.n202 585
R444 B.n204 B.n203 585
R445 B.n353 B.n352 585
R446 B.n352 B.n351 585
R447 B.n354 B.n201 585
R448 B.n350 B.n201 585
R449 B.n356 B.n355 585
R450 B.n357 B.n356 585
R451 B.n196 B.n195 585
R452 B.n197 B.n196 585
R453 B.n365 B.n364 585
R454 B.n364 B.n363 585
R455 B.n366 B.n194 585
R456 B.n194 B.n193 585
R457 B.n368 B.n367 585
R458 B.n369 B.n368 585
R459 B.n188 B.n187 585
R460 B.n189 B.n188 585
R461 B.n377 B.n376 585
R462 B.n376 B.n375 585
R463 B.n378 B.n186 585
R464 B.n186 B.n185 585
R465 B.n380 B.n379 585
R466 B.n381 B.n380 585
R467 B.n180 B.n179 585
R468 B.n181 B.n180 585
R469 B.n390 B.n389 585
R470 B.n389 B.n388 585
R471 B.n391 B.n178 585
R472 B.n387 B.n178 585
R473 B.n393 B.n392 585
R474 B.n394 B.n393 585
R475 B.n173 B.n172 585
R476 B.n174 B.n173 585
R477 B.n402 B.n401 585
R478 B.n401 B.n400 585
R479 B.n403 B.n171 585
R480 B.n171 B.n170 585
R481 B.n405 B.n404 585
R482 B.n406 B.n405 585
R483 B.n165 B.n164 585
R484 B.n166 B.n165 585
R485 B.n415 B.n414 585
R486 B.n414 B.n413 585
R487 B.n416 B.n163 585
R488 B.n412 B.n163 585
R489 B.n418 B.n417 585
R490 B.n419 B.n418 585
R491 B.n158 B.n157 585
R492 B.n159 B.n158 585
R493 B.n427 B.n426 585
R494 B.n426 B.n425 585
R495 B.n428 B.n156 585
R496 B.n156 B.n155 585
R497 B.n430 B.n429 585
R498 B.n431 B.n430 585
R499 B.n150 B.n149 585
R500 B.n151 B.n150 585
R501 B.n439 B.n438 585
R502 B.n438 B.n437 585
R503 B.n440 B.n148 585
R504 B.n148 B.n147 585
R505 B.n442 B.n441 585
R506 B.n443 B.n442 585
R507 B.n142 B.n141 585
R508 B.n143 B.n142 585
R509 B.n451 B.n450 585
R510 B.n450 B.n449 585
R511 B.n452 B.n140 585
R512 B.n140 B.n139 585
R513 B.n454 B.n453 585
R514 B.n455 B.n454 585
R515 B.n134 B.n133 585
R516 B.n135 B.n134 585
R517 B.n463 B.n462 585
R518 B.n462 B.n461 585
R519 B.n464 B.n132 585
R520 B.n132 B.n131 585
R521 B.n466 B.n465 585
R522 B.n467 B.n466 585
R523 B.n126 B.n125 585
R524 B.n127 B.n126 585
R525 B.n476 B.n475 585
R526 B.n475 B.n474 585
R527 B.n477 B.n124 585
R528 B.n124 B.n123 585
R529 B.n479 B.n478 585
R530 B.n480 B.n479 585
R531 B.n3 B.n0 585
R532 B.n4 B.n3 585
R533 B.n736 B.n1 585
R534 B.n737 B.n736 585
R535 B.n735 B.n734 585
R536 B.n735 B.n8 585
R537 B.n733 B.n9 585
R538 B.n12 B.n9 585
R539 B.n732 B.n731 585
R540 B.n731 B.n730 585
R541 B.n11 B.n10 585
R542 B.n729 B.n11 585
R543 B.n727 B.n726 585
R544 B.n728 B.n727 585
R545 B.n725 B.n17 585
R546 B.n17 B.n16 585
R547 B.n724 B.n723 585
R548 B.n723 B.n722 585
R549 B.n19 B.n18 585
R550 B.n721 B.n19 585
R551 B.n719 B.n718 585
R552 B.n720 B.n719 585
R553 B.n717 B.n24 585
R554 B.n24 B.n23 585
R555 B.n716 B.n715 585
R556 B.n715 B.n714 585
R557 B.n26 B.n25 585
R558 B.n713 B.n26 585
R559 B.n711 B.n710 585
R560 B.n712 B.n711 585
R561 B.n709 B.n31 585
R562 B.n31 B.n30 585
R563 B.n708 B.n707 585
R564 B.n707 B.n706 585
R565 B.n33 B.n32 585
R566 B.n705 B.n33 585
R567 B.n703 B.n702 585
R568 B.n704 B.n703 585
R569 B.n701 B.n38 585
R570 B.n38 B.n37 585
R571 B.n700 B.n699 585
R572 B.n699 B.n698 585
R573 B.n40 B.n39 585
R574 B.n697 B.n40 585
R575 B.n695 B.n694 585
R576 B.n696 B.n695 585
R577 B.n693 B.n44 585
R578 B.n47 B.n44 585
R579 B.n692 B.n691 585
R580 B.n691 B.n690 585
R581 B.n46 B.n45 585
R582 B.n689 B.n46 585
R583 B.n687 B.n686 585
R584 B.n688 B.n687 585
R585 B.n685 B.n52 585
R586 B.n52 B.n51 585
R587 B.n684 B.n683 585
R588 B.n683 B.n682 585
R589 B.n54 B.n53 585
R590 B.n681 B.n54 585
R591 B.n679 B.n678 585
R592 B.n680 B.n679 585
R593 B.n677 B.n58 585
R594 B.n61 B.n58 585
R595 B.n676 B.n675 585
R596 B.n675 B.n674 585
R597 B.n60 B.n59 585
R598 B.n673 B.n60 585
R599 B.n671 B.n670 585
R600 B.n672 B.n671 585
R601 B.n669 B.n66 585
R602 B.n66 B.n65 585
R603 B.n668 B.n667 585
R604 B.n667 B.n666 585
R605 B.n68 B.n67 585
R606 B.n665 B.n68 585
R607 B.n663 B.n662 585
R608 B.n664 B.n663 585
R609 B.n661 B.n73 585
R610 B.n73 B.n72 585
R611 B.n660 B.n659 585
R612 B.n659 B.n658 585
R613 B.n75 B.n74 585
R614 B.n657 B.n75 585
R615 B.n655 B.n654 585
R616 B.n656 B.n655 585
R617 B.n653 B.n79 585
R618 B.n82 B.n79 585
R619 B.n652 B.n651 585
R620 B.n651 B.n650 585
R621 B.n81 B.n80 585
R622 B.n649 B.n81 585
R623 B.n647 B.n646 585
R624 B.n648 B.n647 585
R625 B.n645 B.n87 585
R626 B.n87 B.n86 585
R627 B.n644 B.n643 585
R628 B.n643 B.n642 585
R629 B.n89 B.n88 585
R630 B.n641 B.n89 585
R631 B.n639 B.n638 585
R632 B.n640 B.n639 585
R633 B.n740 B.n739 585
R634 B.n738 B.n2 585
R635 B.n639 B.n94 502.111
R636 B.n550 B.n92 502.111
R637 B.n333 B.n215 502.111
R638 B.n331 B.n217 502.111
R639 B.n551 B.n93 256.663
R640 B.n553 B.n93 256.663
R641 B.n559 B.n93 256.663
R642 B.n561 B.n93 256.663
R643 B.n567 B.n93 256.663
R644 B.n569 B.n93 256.663
R645 B.n575 B.n93 256.663
R646 B.n577 B.n93 256.663
R647 B.n583 B.n93 256.663
R648 B.n585 B.n93 256.663
R649 B.n591 B.n93 256.663
R650 B.n593 B.n93 256.663
R651 B.n599 B.n93 256.663
R652 B.n601 B.n93 256.663
R653 B.n608 B.n93 256.663
R654 B.n610 B.n93 256.663
R655 B.n616 B.n93 256.663
R656 B.n618 B.n93 256.663
R657 B.n624 B.n93 256.663
R658 B.n626 B.n93 256.663
R659 B.n632 B.n93 256.663
R660 B.n634 B.n93 256.663
R661 B.n326 B.n216 256.663
R662 B.n219 B.n216 256.663
R663 B.n319 B.n216 256.663
R664 B.n313 B.n216 256.663
R665 B.n311 B.n216 256.663
R666 B.n305 B.n216 256.663
R667 B.n303 B.n216 256.663
R668 B.n297 B.n216 256.663
R669 B.n229 B.n216 256.663
R670 B.n291 B.n216 256.663
R671 B.n285 B.n216 256.663
R672 B.n283 B.n216 256.663
R673 B.n277 B.n216 256.663
R674 B.n237 B.n216 256.663
R675 B.n271 B.n216 256.663
R676 B.n265 B.n216 256.663
R677 B.n263 B.n216 256.663
R678 B.n257 B.n216 256.663
R679 B.n255 B.n216 256.663
R680 B.n249 B.n216 256.663
R681 B.n247 B.n216 256.663
R682 B.n742 B.n741 256.663
R683 B.n103 B.t10 242.536
R684 B.n111 B.t6 242.536
R685 B.n234 B.t13 242.536
R686 B.n226 B.t17 242.536
R687 B.n635 B.n633 163.367
R688 B.n631 B.n96 163.367
R689 B.n627 B.n625 163.367
R690 B.n623 B.n98 163.367
R691 B.n619 B.n617 163.367
R692 B.n615 B.n100 163.367
R693 B.n611 B.n609 163.367
R694 B.n607 B.n102 163.367
R695 B.n602 B.n600 163.367
R696 B.n598 B.n106 163.367
R697 B.n594 B.n592 163.367
R698 B.n590 B.n108 163.367
R699 B.n586 B.n584 163.367
R700 B.n582 B.n110 163.367
R701 B.n578 B.n576 163.367
R702 B.n574 B.n115 163.367
R703 B.n570 B.n568 163.367
R704 B.n566 B.n117 163.367
R705 B.n562 B.n560 163.367
R706 B.n558 B.n119 163.367
R707 B.n554 B.n552 163.367
R708 B.n333 B.n213 163.367
R709 B.n337 B.n213 163.367
R710 B.n337 B.n207 163.367
R711 B.n345 B.n207 163.367
R712 B.n345 B.n205 163.367
R713 B.n349 B.n205 163.367
R714 B.n349 B.n200 163.367
R715 B.n358 B.n200 163.367
R716 B.n358 B.n198 163.367
R717 B.n362 B.n198 163.367
R718 B.n362 B.n192 163.367
R719 B.n370 B.n192 163.367
R720 B.n370 B.n190 163.367
R721 B.n374 B.n190 163.367
R722 B.n374 B.n184 163.367
R723 B.n382 B.n184 163.367
R724 B.n382 B.n182 163.367
R725 B.n386 B.n182 163.367
R726 B.n386 B.n177 163.367
R727 B.n395 B.n177 163.367
R728 B.n395 B.n175 163.367
R729 B.n399 B.n175 163.367
R730 B.n399 B.n169 163.367
R731 B.n407 B.n169 163.367
R732 B.n407 B.n167 163.367
R733 B.n411 B.n167 163.367
R734 B.n411 B.n162 163.367
R735 B.n420 B.n162 163.367
R736 B.n420 B.n160 163.367
R737 B.n424 B.n160 163.367
R738 B.n424 B.n154 163.367
R739 B.n432 B.n154 163.367
R740 B.n432 B.n152 163.367
R741 B.n436 B.n152 163.367
R742 B.n436 B.n146 163.367
R743 B.n444 B.n146 163.367
R744 B.n444 B.n144 163.367
R745 B.n448 B.n144 163.367
R746 B.n448 B.n138 163.367
R747 B.n456 B.n138 163.367
R748 B.n456 B.n136 163.367
R749 B.n460 B.n136 163.367
R750 B.n460 B.n130 163.367
R751 B.n468 B.n130 163.367
R752 B.n468 B.n128 163.367
R753 B.n473 B.n128 163.367
R754 B.n473 B.n122 163.367
R755 B.n481 B.n122 163.367
R756 B.n482 B.n481 163.367
R757 B.n482 B.n5 163.367
R758 B.n6 B.n5 163.367
R759 B.n7 B.n6 163.367
R760 B.n488 B.n7 163.367
R761 B.n489 B.n488 163.367
R762 B.n489 B.n13 163.367
R763 B.n14 B.n13 163.367
R764 B.n15 B.n14 163.367
R765 B.n494 B.n15 163.367
R766 B.n494 B.n20 163.367
R767 B.n21 B.n20 163.367
R768 B.n22 B.n21 163.367
R769 B.n499 B.n22 163.367
R770 B.n499 B.n27 163.367
R771 B.n28 B.n27 163.367
R772 B.n29 B.n28 163.367
R773 B.n504 B.n29 163.367
R774 B.n504 B.n34 163.367
R775 B.n35 B.n34 163.367
R776 B.n36 B.n35 163.367
R777 B.n509 B.n36 163.367
R778 B.n509 B.n41 163.367
R779 B.n42 B.n41 163.367
R780 B.n43 B.n42 163.367
R781 B.n514 B.n43 163.367
R782 B.n514 B.n48 163.367
R783 B.n49 B.n48 163.367
R784 B.n50 B.n49 163.367
R785 B.n519 B.n50 163.367
R786 B.n519 B.n55 163.367
R787 B.n56 B.n55 163.367
R788 B.n57 B.n56 163.367
R789 B.n524 B.n57 163.367
R790 B.n524 B.n62 163.367
R791 B.n63 B.n62 163.367
R792 B.n64 B.n63 163.367
R793 B.n529 B.n64 163.367
R794 B.n529 B.n69 163.367
R795 B.n70 B.n69 163.367
R796 B.n71 B.n70 163.367
R797 B.n534 B.n71 163.367
R798 B.n534 B.n76 163.367
R799 B.n77 B.n76 163.367
R800 B.n78 B.n77 163.367
R801 B.n539 B.n78 163.367
R802 B.n539 B.n83 163.367
R803 B.n84 B.n83 163.367
R804 B.n85 B.n84 163.367
R805 B.n544 B.n85 163.367
R806 B.n544 B.n90 163.367
R807 B.n91 B.n90 163.367
R808 B.n92 B.n91 163.367
R809 B.n327 B.n325 163.367
R810 B.n325 B.n324 163.367
R811 B.n321 B.n320 163.367
R812 B.n318 B.n221 163.367
R813 B.n314 B.n312 163.367
R814 B.n310 B.n223 163.367
R815 B.n306 B.n304 163.367
R816 B.n302 B.n225 163.367
R817 B.n298 B.n296 163.367
R818 B.n293 B.n292 163.367
R819 B.n290 B.n231 163.367
R820 B.n286 B.n284 163.367
R821 B.n282 B.n233 163.367
R822 B.n278 B.n276 163.367
R823 B.n273 B.n272 163.367
R824 B.n270 B.n239 163.367
R825 B.n266 B.n264 163.367
R826 B.n262 B.n241 163.367
R827 B.n258 B.n256 163.367
R828 B.n254 B.n243 163.367
R829 B.n250 B.n248 163.367
R830 B.n246 B.n215 163.367
R831 B.n331 B.n211 163.367
R832 B.n339 B.n211 163.367
R833 B.n339 B.n209 163.367
R834 B.n343 B.n209 163.367
R835 B.n343 B.n203 163.367
R836 B.n352 B.n203 163.367
R837 B.n352 B.n201 163.367
R838 B.n356 B.n201 163.367
R839 B.n356 B.n196 163.367
R840 B.n364 B.n196 163.367
R841 B.n364 B.n194 163.367
R842 B.n368 B.n194 163.367
R843 B.n368 B.n188 163.367
R844 B.n376 B.n188 163.367
R845 B.n376 B.n186 163.367
R846 B.n380 B.n186 163.367
R847 B.n380 B.n180 163.367
R848 B.n389 B.n180 163.367
R849 B.n389 B.n178 163.367
R850 B.n393 B.n178 163.367
R851 B.n393 B.n173 163.367
R852 B.n401 B.n173 163.367
R853 B.n401 B.n171 163.367
R854 B.n405 B.n171 163.367
R855 B.n405 B.n165 163.367
R856 B.n414 B.n165 163.367
R857 B.n414 B.n163 163.367
R858 B.n418 B.n163 163.367
R859 B.n418 B.n158 163.367
R860 B.n426 B.n158 163.367
R861 B.n426 B.n156 163.367
R862 B.n430 B.n156 163.367
R863 B.n430 B.n150 163.367
R864 B.n438 B.n150 163.367
R865 B.n438 B.n148 163.367
R866 B.n442 B.n148 163.367
R867 B.n442 B.n142 163.367
R868 B.n450 B.n142 163.367
R869 B.n450 B.n140 163.367
R870 B.n454 B.n140 163.367
R871 B.n454 B.n134 163.367
R872 B.n462 B.n134 163.367
R873 B.n462 B.n132 163.367
R874 B.n466 B.n132 163.367
R875 B.n466 B.n126 163.367
R876 B.n475 B.n126 163.367
R877 B.n475 B.n124 163.367
R878 B.n479 B.n124 163.367
R879 B.n479 B.n3 163.367
R880 B.n740 B.n3 163.367
R881 B.n736 B.n2 163.367
R882 B.n736 B.n735 163.367
R883 B.n735 B.n9 163.367
R884 B.n731 B.n9 163.367
R885 B.n731 B.n11 163.367
R886 B.n727 B.n11 163.367
R887 B.n727 B.n17 163.367
R888 B.n723 B.n17 163.367
R889 B.n723 B.n19 163.367
R890 B.n719 B.n19 163.367
R891 B.n719 B.n24 163.367
R892 B.n715 B.n24 163.367
R893 B.n715 B.n26 163.367
R894 B.n711 B.n26 163.367
R895 B.n711 B.n31 163.367
R896 B.n707 B.n31 163.367
R897 B.n707 B.n33 163.367
R898 B.n703 B.n33 163.367
R899 B.n703 B.n38 163.367
R900 B.n699 B.n38 163.367
R901 B.n699 B.n40 163.367
R902 B.n695 B.n40 163.367
R903 B.n695 B.n44 163.367
R904 B.n691 B.n44 163.367
R905 B.n691 B.n46 163.367
R906 B.n687 B.n46 163.367
R907 B.n687 B.n52 163.367
R908 B.n683 B.n52 163.367
R909 B.n683 B.n54 163.367
R910 B.n679 B.n54 163.367
R911 B.n679 B.n58 163.367
R912 B.n675 B.n58 163.367
R913 B.n675 B.n60 163.367
R914 B.n671 B.n60 163.367
R915 B.n671 B.n66 163.367
R916 B.n667 B.n66 163.367
R917 B.n667 B.n68 163.367
R918 B.n663 B.n68 163.367
R919 B.n663 B.n73 163.367
R920 B.n659 B.n73 163.367
R921 B.n659 B.n75 163.367
R922 B.n655 B.n75 163.367
R923 B.n655 B.n79 163.367
R924 B.n651 B.n79 163.367
R925 B.n651 B.n81 163.367
R926 B.n647 B.n81 163.367
R927 B.n647 B.n87 163.367
R928 B.n643 B.n87 163.367
R929 B.n643 B.n89 163.367
R930 B.n639 B.n89 163.367
R931 B.n332 B.n216 161.096
R932 B.n640 B.n93 161.096
R933 B.n111 B.t8 133.642
R934 B.n234 B.t16 133.642
R935 B.n103 B.t11 133.638
R936 B.n226 B.t19 133.638
R937 B.n332 B.n212 83.6226
R938 B.n338 B.n212 83.6226
R939 B.n338 B.n208 83.6226
R940 B.n344 B.n208 83.6226
R941 B.n344 B.n204 83.6226
R942 B.n351 B.n204 83.6226
R943 B.n351 B.n350 83.6226
R944 B.n357 B.n197 83.6226
R945 B.n363 B.n197 83.6226
R946 B.n363 B.n193 83.6226
R947 B.n369 B.n193 83.6226
R948 B.n369 B.n189 83.6226
R949 B.n375 B.n189 83.6226
R950 B.n375 B.n185 83.6226
R951 B.n381 B.n185 83.6226
R952 B.n381 B.n181 83.6226
R953 B.n388 B.n181 83.6226
R954 B.n388 B.n387 83.6226
R955 B.n394 B.n174 83.6226
R956 B.n400 B.n174 83.6226
R957 B.n400 B.n170 83.6226
R958 B.n406 B.n170 83.6226
R959 B.n406 B.n166 83.6226
R960 B.n413 B.n166 83.6226
R961 B.n413 B.n412 83.6226
R962 B.n419 B.n159 83.6226
R963 B.n425 B.n159 83.6226
R964 B.n425 B.n155 83.6226
R965 B.n431 B.n155 83.6226
R966 B.n431 B.n151 83.6226
R967 B.n437 B.n151 83.6226
R968 B.n437 B.n147 83.6226
R969 B.n443 B.n147 83.6226
R970 B.n449 B.n143 83.6226
R971 B.n449 B.n139 83.6226
R972 B.n455 B.n139 83.6226
R973 B.n455 B.n135 83.6226
R974 B.n461 B.n135 83.6226
R975 B.n461 B.n131 83.6226
R976 B.n467 B.n131 83.6226
R977 B.n474 B.n127 83.6226
R978 B.n474 B.n123 83.6226
R979 B.n480 B.n123 83.6226
R980 B.n480 B.n4 83.6226
R981 B.n739 B.n4 83.6226
R982 B.n739 B.n738 83.6226
R983 B.n738 B.n737 83.6226
R984 B.n737 B.n8 83.6226
R985 B.n12 B.n8 83.6226
R986 B.n730 B.n12 83.6226
R987 B.n730 B.n729 83.6226
R988 B.n728 B.n16 83.6226
R989 B.n722 B.n16 83.6226
R990 B.n722 B.n721 83.6226
R991 B.n721 B.n720 83.6226
R992 B.n720 B.n23 83.6226
R993 B.n714 B.n23 83.6226
R994 B.n714 B.n713 83.6226
R995 B.n712 B.n30 83.6226
R996 B.n706 B.n30 83.6226
R997 B.n706 B.n705 83.6226
R998 B.n705 B.n704 83.6226
R999 B.n704 B.n37 83.6226
R1000 B.n698 B.n37 83.6226
R1001 B.n698 B.n697 83.6226
R1002 B.n697 B.n696 83.6226
R1003 B.n690 B.n47 83.6226
R1004 B.n690 B.n689 83.6226
R1005 B.n689 B.n688 83.6226
R1006 B.n688 B.n51 83.6226
R1007 B.n682 B.n51 83.6226
R1008 B.n682 B.n681 83.6226
R1009 B.n681 B.n680 83.6226
R1010 B.n674 B.n61 83.6226
R1011 B.n674 B.n673 83.6226
R1012 B.n673 B.n672 83.6226
R1013 B.n672 B.n65 83.6226
R1014 B.n666 B.n65 83.6226
R1015 B.n666 B.n665 83.6226
R1016 B.n665 B.n664 83.6226
R1017 B.n664 B.n72 83.6226
R1018 B.n658 B.n72 83.6226
R1019 B.n658 B.n657 83.6226
R1020 B.n657 B.n656 83.6226
R1021 B.n650 B.n82 83.6226
R1022 B.n650 B.n649 83.6226
R1023 B.n649 B.n648 83.6226
R1024 B.n648 B.n86 83.6226
R1025 B.n642 B.n86 83.6226
R1026 B.n642 B.n641 83.6226
R1027 B.n641 B.n640 83.6226
R1028 B.n112 B.t9 77.593
R1029 B.n235 B.t15 77.593
R1030 B.n104 B.t12 77.5901
R1031 B.n227 B.t18 77.5901
R1032 B.n634 B.n94 71.676
R1033 B.n633 B.n632 71.676
R1034 B.n626 B.n96 71.676
R1035 B.n625 B.n624 71.676
R1036 B.n618 B.n98 71.676
R1037 B.n617 B.n616 71.676
R1038 B.n610 B.n100 71.676
R1039 B.n609 B.n608 71.676
R1040 B.n601 B.n102 71.676
R1041 B.n600 B.n599 71.676
R1042 B.n593 B.n106 71.676
R1043 B.n592 B.n591 71.676
R1044 B.n585 B.n108 71.676
R1045 B.n584 B.n583 71.676
R1046 B.n577 B.n110 71.676
R1047 B.n576 B.n575 71.676
R1048 B.n569 B.n115 71.676
R1049 B.n568 B.n567 71.676
R1050 B.n561 B.n117 71.676
R1051 B.n560 B.n559 71.676
R1052 B.n553 B.n119 71.676
R1053 B.n552 B.n551 71.676
R1054 B.n551 B.n550 71.676
R1055 B.n554 B.n553 71.676
R1056 B.n559 B.n558 71.676
R1057 B.n562 B.n561 71.676
R1058 B.n567 B.n566 71.676
R1059 B.n570 B.n569 71.676
R1060 B.n575 B.n574 71.676
R1061 B.n578 B.n577 71.676
R1062 B.n583 B.n582 71.676
R1063 B.n586 B.n585 71.676
R1064 B.n591 B.n590 71.676
R1065 B.n594 B.n593 71.676
R1066 B.n599 B.n598 71.676
R1067 B.n602 B.n601 71.676
R1068 B.n608 B.n607 71.676
R1069 B.n611 B.n610 71.676
R1070 B.n616 B.n615 71.676
R1071 B.n619 B.n618 71.676
R1072 B.n624 B.n623 71.676
R1073 B.n627 B.n626 71.676
R1074 B.n632 B.n631 71.676
R1075 B.n635 B.n634 71.676
R1076 B.n326 B.n217 71.676
R1077 B.n324 B.n219 71.676
R1078 B.n320 B.n319 71.676
R1079 B.n313 B.n221 71.676
R1080 B.n312 B.n311 71.676
R1081 B.n305 B.n223 71.676
R1082 B.n304 B.n303 71.676
R1083 B.n297 B.n225 71.676
R1084 B.n296 B.n229 71.676
R1085 B.n292 B.n291 71.676
R1086 B.n285 B.n231 71.676
R1087 B.n284 B.n283 71.676
R1088 B.n277 B.n233 71.676
R1089 B.n276 B.n237 71.676
R1090 B.n272 B.n271 71.676
R1091 B.n265 B.n239 71.676
R1092 B.n264 B.n263 71.676
R1093 B.n257 B.n241 71.676
R1094 B.n256 B.n255 71.676
R1095 B.n249 B.n243 71.676
R1096 B.n248 B.n247 71.676
R1097 B.n327 B.n326 71.676
R1098 B.n321 B.n219 71.676
R1099 B.n319 B.n318 71.676
R1100 B.n314 B.n313 71.676
R1101 B.n311 B.n310 71.676
R1102 B.n306 B.n305 71.676
R1103 B.n303 B.n302 71.676
R1104 B.n298 B.n297 71.676
R1105 B.n293 B.n229 71.676
R1106 B.n291 B.n290 71.676
R1107 B.n286 B.n285 71.676
R1108 B.n283 B.n282 71.676
R1109 B.n278 B.n277 71.676
R1110 B.n273 B.n237 71.676
R1111 B.n271 B.n270 71.676
R1112 B.n266 B.n265 71.676
R1113 B.n263 B.n262 71.676
R1114 B.n258 B.n257 71.676
R1115 B.n255 B.n254 71.676
R1116 B.n250 B.n249 71.676
R1117 B.n247 B.n246 71.676
R1118 B.n741 B.n740 71.676
R1119 B.n741 B.n2 71.676
R1120 B.n394 B.t20 71.3253
R1121 B.t4 B.n143 71.3253
R1122 B.n713 B.t1 71.3253
R1123 B.n680 B.t5 71.3253
R1124 B.n604 B.n104 59.5399
R1125 B.n113 B.n112 59.5399
R1126 B.n236 B.n235 59.5399
R1127 B.n228 B.n227 59.5399
R1128 B.n104 B.n103 56.049
R1129 B.n112 B.n111 56.049
R1130 B.n235 B.n234 56.049
R1131 B.n227 B.n226 56.049
R1132 B.n412 B.t2 54.1089
R1133 B.n467 B.t0 54.1089
R1134 B.t3 B.n728 54.1089
R1135 B.n47 B.t21 54.1089
R1136 B.n357 B.t14 46.7305
R1137 B.n656 B.t7 46.7305
R1138 B.n350 B.t14 36.8926
R1139 B.n82 B.t7 36.8926
R1140 B.n330 B.n329 32.6249
R1141 B.n334 B.n214 32.6249
R1142 B.n549 B.n548 32.6249
R1143 B.n638 B.n637 32.6249
R1144 B.n419 B.t2 29.5142
R1145 B.t0 B.n127 29.5142
R1146 B.n729 B.t3 29.5142
R1147 B.n696 B.t21 29.5142
R1148 B B.n742 18.0485
R1149 B.n387 B.t20 12.2979
R1150 B.n443 B.t4 12.2979
R1151 B.t1 B.n712 12.2979
R1152 B.n61 B.t5 12.2979
R1153 B.n330 B.n210 10.6151
R1154 B.n340 B.n210 10.6151
R1155 B.n341 B.n340 10.6151
R1156 B.n342 B.n341 10.6151
R1157 B.n342 B.n202 10.6151
R1158 B.n353 B.n202 10.6151
R1159 B.n354 B.n353 10.6151
R1160 B.n355 B.n354 10.6151
R1161 B.n355 B.n195 10.6151
R1162 B.n365 B.n195 10.6151
R1163 B.n366 B.n365 10.6151
R1164 B.n367 B.n366 10.6151
R1165 B.n367 B.n187 10.6151
R1166 B.n377 B.n187 10.6151
R1167 B.n378 B.n377 10.6151
R1168 B.n379 B.n378 10.6151
R1169 B.n379 B.n179 10.6151
R1170 B.n390 B.n179 10.6151
R1171 B.n391 B.n390 10.6151
R1172 B.n392 B.n391 10.6151
R1173 B.n392 B.n172 10.6151
R1174 B.n402 B.n172 10.6151
R1175 B.n403 B.n402 10.6151
R1176 B.n404 B.n403 10.6151
R1177 B.n404 B.n164 10.6151
R1178 B.n415 B.n164 10.6151
R1179 B.n416 B.n415 10.6151
R1180 B.n417 B.n416 10.6151
R1181 B.n417 B.n157 10.6151
R1182 B.n427 B.n157 10.6151
R1183 B.n428 B.n427 10.6151
R1184 B.n429 B.n428 10.6151
R1185 B.n429 B.n149 10.6151
R1186 B.n439 B.n149 10.6151
R1187 B.n440 B.n439 10.6151
R1188 B.n441 B.n440 10.6151
R1189 B.n441 B.n141 10.6151
R1190 B.n451 B.n141 10.6151
R1191 B.n452 B.n451 10.6151
R1192 B.n453 B.n452 10.6151
R1193 B.n453 B.n133 10.6151
R1194 B.n463 B.n133 10.6151
R1195 B.n464 B.n463 10.6151
R1196 B.n465 B.n464 10.6151
R1197 B.n465 B.n125 10.6151
R1198 B.n476 B.n125 10.6151
R1199 B.n477 B.n476 10.6151
R1200 B.n478 B.n477 10.6151
R1201 B.n478 B.n0 10.6151
R1202 B.n329 B.n328 10.6151
R1203 B.n328 B.n218 10.6151
R1204 B.n323 B.n218 10.6151
R1205 B.n323 B.n322 10.6151
R1206 B.n322 B.n220 10.6151
R1207 B.n317 B.n220 10.6151
R1208 B.n317 B.n316 10.6151
R1209 B.n316 B.n315 10.6151
R1210 B.n315 B.n222 10.6151
R1211 B.n309 B.n222 10.6151
R1212 B.n309 B.n308 10.6151
R1213 B.n308 B.n307 10.6151
R1214 B.n307 B.n224 10.6151
R1215 B.n301 B.n224 10.6151
R1216 B.n301 B.n300 10.6151
R1217 B.n300 B.n299 10.6151
R1218 B.n295 B.n294 10.6151
R1219 B.n294 B.n230 10.6151
R1220 B.n289 B.n230 10.6151
R1221 B.n289 B.n288 10.6151
R1222 B.n288 B.n287 10.6151
R1223 B.n287 B.n232 10.6151
R1224 B.n281 B.n232 10.6151
R1225 B.n281 B.n280 10.6151
R1226 B.n280 B.n279 10.6151
R1227 B.n275 B.n274 10.6151
R1228 B.n274 B.n238 10.6151
R1229 B.n269 B.n238 10.6151
R1230 B.n269 B.n268 10.6151
R1231 B.n268 B.n267 10.6151
R1232 B.n267 B.n240 10.6151
R1233 B.n261 B.n240 10.6151
R1234 B.n261 B.n260 10.6151
R1235 B.n260 B.n259 10.6151
R1236 B.n259 B.n242 10.6151
R1237 B.n253 B.n242 10.6151
R1238 B.n253 B.n252 10.6151
R1239 B.n252 B.n251 10.6151
R1240 B.n251 B.n244 10.6151
R1241 B.n245 B.n244 10.6151
R1242 B.n245 B.n214 10.6151
R1243 B.n335 B.n334 10.6151
R1244 B.n336 B.n335 10.6151
R1245 B.n336 B.n206 10.6151
R1246 B.n346 B.n206 10.6151
R1247 B.n347 B.n346 10.6151
R1248 B.n348 B.n347 10.6151
R1249 B.n348 B.n199 10.6151
R1250 B.n359 B.n199 10.6151
R1251 B.n360 B.n359 10.6151
R1252 B.n361 B.n360 10.6151
R1253 B.n361 B.n191 10.6151
R1254 B.n371 B.n191 10.6151
R1255 B.n372 B.n371 10.6151
R1256 B.n373 B.n372 10.6151
R1257 B.n373 B.n183 10.6151
R1258 B.n383 B.n183 10.6151
R1259 B.n384 B.n383 10.6151
R1260 B.n385 B.n384 10.6151
R1261 B.n385 B.n176 10.6151
R1262 B.n396 B.n176 10.6151
R1263 B.n397 B.n396 10.6151
R1264 B.n398 B.n397 10.6151
R1265 B.n398 B.n168 10.6151
R1266 B.n408 B.n168 10.6151
R1267 B.n409 B.n408 10.6151
R1268 B.n410 B.n409 10.6151
R1269 B.n410 B.n161 10.6151
R1270 B.n421 B.n161 10.6151
R1271 B.n422 B.n421 10.6151
R1272 B.n423 B.n422 10.6151
R1273 B.n423 B.n153 10.6151
R1274 B.n433 B.n153 10.6151
R1275 B.n434 B.n433 10.6151
R1276 B.n435 B.n434 10.6151
R1277 B.n435 B.n145 10.6151
R1278 B.n445 B.n145 10.6151
R1279 B.n446 B.n445 10.6151
R1280 B.n447 B.n446 10.6151
R1281 B.n447 B.n137 10.6151
R1282 B.n457 B.n137 10.6151
R1283 B.n458 B.n457 10.6151
R1284 B.n459 B.n458 10.6151
R1285 B.n459 B.n129 10.6151
R1286 B.n469 B.n129 10.6151
R1287 B.n470 B.n469 10.6151
R1288 B.n472 B.n470 10.6151
R1289 B.n472 B.n471 10.6151
R1290 B.n471 B.n121 10.6151
R1291 B.n483 B.n121 10.6151
R1292 B.n484 B.n483 10.6151
R1293 B.n485 B.n484 10.6151
R1294 B.n486 B.n485 10.6151
R1295 B.n487 B.n486 10.6151
R1296 B.n490 B.n487 10.6151
R1297 B.n491 B.n490 10.6151
R1298 B.n492 B.n491 10.6151
R1299 B.n493 B.n492 10.6151
R1300 B.n495 B.n493 10.6151
R1301 B.n496 B.n495 10.6151
R1302 B.n497 B.n496 10.6151
R1303 B.n498 B.n497 10.6151
R1304 B.n500 B.n498 10.6151
R1305 B.n501 B.n500 10.6151
R1306 B.n502 B.n501 10.6151
R1307 B.n503 B.n502 10.6151
R1308 B.n505 B.n503 10.6151
R1309 B.n506 B.n505 10.6151
R1310 B.n507 B.n506 10.6151
R1311 B.n508 B.n507 10.6151
R1312 B.n510 B.n508 10.6151
R1313 B.n511 B.n510 10.6151
R1314 B.n512 B.n511 10.6151
R1315 B.n513 B.n512 10.6151
R1316 B.n515 B.n513 10.6151
R1317 B.n516 B.n515 10.6151
R1318 B.n517 B.n516 10.6151
R1319 B.n518 B.n517 10.6151
R1320 B.n520 B.n518 10.6151
R1321 B.n521 B.n520 10.6151
R1322 B.n522 B.n521 10.6151
R1323 B.n523 B.n522 10.6151
R1324 B.n525 B.n523 10.6151
R1325 B.n526 B.n525 10.6151
R1326 B.n527 B.n526 10.6151
R1327 B.n528 B.n527 10.6151
R1328 B.n530 B.n528 10.6151
R1329 B.n531 B.n530 10.6151
R1330 B.n532 B.n531 10.6151
R1331 B.n533 B.n532 10.6151
R1332 B.n535 B.n533 10.6151
R1333 B.n536 B.n535 10.6151
R1334 B.n537 B.n536 10.6151
R1335 B.n538 B.n537 10.6151
R1336 B.n540 B.n538 10.6151
R1337 B.n541 B.n540 10.6151
R1338 B.n542 B.n541 10.6151
R1339 B.n543 B.n542 10.6151
R1340 B.n545 B.n543 10.6151
R1341 B.n546 B.n545 10.6151
R1342 B.n547 B.n546 10.6151
R1343 B.n548 B.n547 10.6151
R1344 B.n734 B.n1 10.6151
R1345 B.n734 B.n733 10.6151
R1346 B.n733 B.n732 10.6151
R1347 B.n732 B.n10 10.6151
R1348 B.n726 B.n10 10.6151
R1349 B.n726 B.n725 10.6151
R1350 B.n725 B.n724 10.6151
R1351 B.n724 B.n18 10.6151
R1352 B.n718 B.n18 10.6151
R1353 B.n718 B.n717 10.6151
R1354 B.n717 B.n716 10.6151
R1355 B.n716 B.n25 10.6151
R1356 B.n710 B.n25 10.6151
R1357 B.n710 B.n709 10.6151
R1358 B.n709 B.n708 10.6151
R1359 B.n708 B.n32 10.6151
R1360 B.n702 B.n32 10.6151
R1361 B.n702 B.n701 10.6151
R1362 B.n701 B.n700 10.6151
R1363 B.n700 B.n39 10.6151
R1364 B.n694 B.n39 10.6151
R1365 B.n694 B.n693 10.6151
R1366 B.n693 B.n692 10.6151
R1367 B.n692 B.n45 10.6151
R1368 B.n686 B.n45 10.6151
R1369 B.n686 B.n685 10.6151
R1370 B.n685 B.n684 10.6151
R1371 B.n684 B.n53 10.6151
R1372 B.n678 B.n53 10.6151
R1373 B.n678 B.n677 10.6151
R1374 B.n677 B.n676 10.6151
R1375 B.n676 B.n59 10.6151
R1376 B.n670 B.n59 10.6151
R1377 B.n670 B.n669 10.6151
R1378 B.n669 B.n668 10.6151
R1379 B.n668 B.n67 10.6151
R1380 B.n662 B.n67 10.6151
R1381 B.n662 B.n661 10.6151
R1382 B.n661 B.n660 10.6151
R1383 B.n660 B.n74 10.6151
R1384 B.n654 B.n74 10.6151
R1385 B.n654 B.n653 10.6151
R1386 B.n653 B.n652 10.6151
R1387 B.n652 B.n80 10.6151
R1388 B.n646 B.n80 10.6151
R1389 B.n646 B.n645 10.6151
R1390 B.n645 B.n644 10.6151
R1391 B.n644 B.n88 10.6151
R1392 B.n638 B.n88 10.6151
R1393 B.n637 B.n636 10.6151
R1394 B.n636 B.n95 10.6151
R1395 B.n630 B.n95 10.6151
R1396 B.n630 B.n629 10.6151
R1397 B.n629 B.n628 10.6151
R1398 B.n628 B.n97 10.6151
R1399 B.n622 B.n97 10.6151
R1400 B.n622 B.n621 10.6151
R1401 B.n621 B.n620 10.6151
R1402 B.n620 B.n99 10.6151
R1403 B.n614 B.n99 10.6151
R1404 B.n614 B.n613 10.6151
R1405 B.n613 B.n612 10.6151
R1406 B.n612 B.n101 10.6151
R1407 B.n606 B.n101 10.6151
R1408 B.n606 B.n605 10.6151
R1409 B.n603 B.n105 10.6151
R1410 B.n597 B.n105 10.6151
R1411 B.n597 B.n596 10.6151
R1412 B.n596 B.n595 10.6151
R1413 B.n595 B.n107 10.6151
R1414 B.n589 B.n107 10.6151
R1415 B.n589 B.n588 10.6151
R1416 B.n588 B.n587 10.6151
R1417 B.n587 B.n109 10.6151
R1418 B.n581 B.n580 10.6151
R1419 B.n580 B.n579 10.6151
R1420 B.n579 B.n114 10.6151
R1421 B.n573 B.n114 10.6151
R1422 B.n573 B.n572 10.6151
R1423 B.n572 B.n571 10.6151
R1424 B.n571 B.n116 10.6151
R1425 B.n565 B.n116 10.6151
R1426 B.n565 B.n564 10.6151
R1427 B.n564 B.n563 10.6151
R1428 B.n563 B.n118 10.6151
R1429 B.n557 B.n118 10.6151
R1430 B.n557 B.n556 10.6151
R1431 B.n556 B.n555 10.6151
R1432 B.n555 B.n120 10.6151
R1433 B.n549 B.n120 10.6151
R1434 B.n299 B.n228 9.36635
R1435 B.n275 B.n236 9.36635
R1436 B.n605 B.n604 9.36635
R1437 B.n581 B.n113 9.36635
R1438 B.n742 B.n0 8.11757
R1439 B.n742 B.n1 8.11757
R1440 B.n295 B.n228 1.24928
R1441 B.n279 B.n236 1.24928
R1442 B.n604 B.n603 1.24928
R1443 B.n113 B.n109 1.24928
R1444 VP.n19 VP.n16 161.3
R1445 VP.n21 VP.n20 161.3
R1446 VP.n22 VP.n15 161.3
R1447 VP.n24 VP.n23 161.3
R1448 VP.n25 VP.n14 161.3
R1449 VP.n27 VP.n26 161.3
R1450 VP.n29 VP.n28 161.3
R1451 VP.n30 VP.n12 161.3
R1452 VP.n32 VP.n31 161.3
R1453 VP.n33 VP.n11 161.3
R1454 VP.n35 VP.n34 161.3
R1455 VP.n36 VP.n10 161.3
R1456 VP.n68 VP.n0 161.3
R1457 VP.n67 VP.n66 161.3
R1458 VP.n65 VP.n1 161.3
R1459 VP.n64 VP.n63 161.3
R1460 VP.n62 VP.n2 161.3
R1461 VP.n61 VP.n60 161.3
R1462 VP.n59 VP.n58 161.3
R1463 VP.n57 VP.n4 161.3
R1464 VP.n56 VP.n55 161.3
R1465 VP.n54 VP.n5 161.3
R1466 VP.n53 VP.n52 161.3
R1467 VP.n51 VP.n6 161.3
R1468 VP.n49 VP.n48 161.3
R1469 VP.n47 VP.n7 161.3
R1470 VP.n46 VP.n45 161.3
R1471 VP.n44 VP.n8 161.3
R1472 VP.n43 VP.n42 161.3
R1473 VP.n41 VP.n9 161.3
R1474 VP.n40 VP.n39 106.597
R1475 VP.n70 VP.n69 106.597
R1476 VP.n38 VP.n37 106.597
R1477 VP.n17 VP.t0 66.272
R1478 VP.n18 VP.n17 62.8231
R1479 VP.n56 VP.n5 56.5193
R1480 VP.n24 VP.n15 56.5193
R1481 VP.n45 VP.n44 54.0911
R1482 VP.n63 VP.n1 54.0911
R1483 VP.n31 VP.n11 54.0911
R1484 VP.n40 VP.n38 44.3178
R1485 VP.n39 VP.t7 34.5501
R1486 VP.n50 VP.t2 34.5501
R1487 VP.n3 VP.t1 34.5501
R1488 VP.n69 VP.t4 34.5501
R1489 VP.n37 VP.t5 34.5501
R1490 VP.n13 VP.t6 34.5501
R1491 VP.n18 VP.t3 34.5501
R1492 VP.n45 VP.n7 26.8957
R1493 VP.n63 VP.n62 26.8957
R1494 VP.n31 VP.n30 26.8957
R1495 VP.n43 VP.n9 24.4675
R1496 VP.n44 VP.n43 24.4675
R1497 VP.n49 VP.n7 24.4675
R1498 VP.n52 VP.n51 24.4675
R1499 VP.n52 VP.n5 24.4675
R1500 VP.n57 VP.n56 24.4675
R1501 VP.n58 VP.n57 24.4675
R1502 VP.n62 VP.n61 24.4675
R1503 VP.n67 VP.n1 24.4675
R1504 VP.n68 VP.n67 24.4675
R1505 VP.n35 VP.n11 24.4675
R1506 VP.n36 VP.n35 24.4675
R1507 VP.n25 VP.n24 24.4675
R1508 VP.n26 VP.n25 24.4675
R1509 VP.n30 VP.n29 24.4675
R1510 VP.n20 VP.n19 24.4675
R1511 VP.n20 VP.n15 24.4675
R1512 VP.n50 VP.n49 14.9254
R1513 VP.n61 VP.n3 14.9254
R1514 VP.n29 VP.n13 14.9254
R1515 VP.n51 VP.n50 9.54263
R1516 VP.n58 VP.n3 9.54263
R1517 VP.n26 VP.n13 9.54263
R1518 VP.n19 VP.n18 9.54263
R1519 VP.n17 VP.n16 7.21701
R1520 VP.n39 VP.n9 4.15989
R1521 VP.n69 VP.n68 4.15989
R1522 VP.n37 VP.n36 4.15989
R1523 VP.n38 VP.n10 0.278367
R1524 VP.n41 VP.n40 0.278367
R1525 VP.n70 VP.n0 0.278367
R1526 VP.n21 VP.n16 0.189894
R1527 VP.n22 VP.n21 0.189894
R1528 VP.n23 VP.n22 0.189894
R1529 VP.n23 VP.n14 0.189894
R1530 VP.n27 VP.n14 0.189894
R1531 VP.n28 VP.n27 0.189894
R1532 VP.n28 VP.n12 0.189894
R1533 VP.n32 VP.n12 0.189894
R1534 VP.n33 VP.n32 0.189894
R1535 VP.n34 VP.n33 0.189894
R1536 VP.n34 VP.n10 0.189894
R1537 VP.n42 VP.n41 0.189894
R1538 VP.n42 VP.n8 0.189894
R1539 VP.n46 VP.n8 0.189894
R1540 VP.n47 VP.n46 0.189894
R1541 VP.n48 VP.n47 0.189894
R1542 VP.n48 VP.n6 0.189894
R1543 VP.n53 VP.n6 0.189894
R1544 VP.n54 VP.n53 0.189894
R1545 VP.n55 VP.n54 0.189894
R1546 VP.n55 VP.n4 0.189894
R1547 VP.n59 VP.n4 0.189894
R1548 VP.n60 VP.n59 0.189894
R1549 VP.n60 VP.n2 0.189894
R1550 VP.n64 VP.n2 0.189894
R1551 VP.n65 VP.n64 0.189894
R1552 VP.n66 VP.n65 0.189894
R1553 VP.n66 VP.n0 0.189894
R1554 VP VP.n70 0.153454
R1555 VDD1 VDD1.n0 80.3494
R1556 VDD1.n3 VDD1.n2 80.2356
R1557 VDD1.n3 VDD1.n1 80.2356
R1558 VDD1.n5 VDD1.n4 79.0454
R1559 VDD1.n5 VDD1.n3 38.6733
R1560 VDD1.n4 VDD1.t1 5.3956
R1561 VDD1.n4 VDD1.t2 5.3956
R1562 VDD1.n0 VDD1.t7 5.3956
R1563 VDD1.n0 VDD1.t4 5.3956
R1564 VDD1.n2 VDD1.t6 5.3956
R1565 VDD1.n2 VDD1.t3 5.3956
R1566 VDD1.n1 VDD1.t0 5.3956
R1567 VDD1.n1 VDD1.t5 5.3956
R1568 VDD1 VDD1.n5 1.188
C0 VTAIL VN 3.92528f
C1 VDD2 VP 0.520577f
C2 VDD1 VP 3.3255f
C3 VDD1 VDD2 1.75652f
C4 VN VP 6.08039f
C5 VTAIL VP 3.93938f
C6 VN VDD2 2.96327f
C7 VTAIL VDD2 5.29906f
C8 VDD1 VN 0.15616f
C9 VDD1 VTAIL 5.24491f
C10 VDD2 B 4.645095f
C11 VDD1 B 5.078581f
C12 VTAIL B 5.082615f
C13 VN B 14.56684f
C14 VP B 13.138449f
C15 VDD1.t7 B 0.071418f
C16 VDD1.t4 B 0.071418f
C17 VDD1.n0 B 0.559548f
C18 VDD1.t0 B 0.071418f
C19 VDD1.t5 B 0.071418f
C20 VDD1.n1 B 0.558721f
C21 VDD1.t6 B 0.071418f
C22 VDD1.t3 B 0.071418f
C23 VDD1.n2 B 0.558721f
C24 VDD1.n3 B 2.73591f
C25 VDD1.t1 B 0.071418f
C26 VDD1.t2 B 0.071418f
C27 VDD1.n4 B 0.551401f
C28 VDD1.n5 B 2.27292f
C29 VP.n0 B 0.03706f
C30 VP.t4 B 0.672902f
C31 VP.n1 B 0.049271f
C32 VP.n2 B 0.02811f
C33 VP.t1 B 0.672902f
C34 VP.n3 B 0.272571f
C35 VP.n4 B 0.02811f
C36 VP.n5 B 0.041035f
C37 VP.n6 B 0.02811f
C38 VP.t2 B 0.672902f
C39 VP.n7 B 0.05449f
C40 VP.n8 B 0.02811f
C41 VP.n9 B 0.03092f
C42 VP.n10 B 0.03706f
C43 VP.t5 B 0.672902f
C44 VP.n11 B 0.049271f
C45 VP.n12 B 0.02811f
C46 VP.t6 B 0.672902f
C47 VP.n13 B 0.272571f
C48 VP.n14 B 0.02811f
C49 VP.n15 B 0.041035f
C50 VP.n16 B 0.27001f
C51 VP.t3 B 0.672902f
C52 VP.t0 B 0.884565f
C53 VP.n17 B 0.34248f
C54 VP.n18 B 0.350312f
C55 VP.n19 B 0.036611f
C56 VP.n20 B 0.05239f
C57 VP.n21 B 0.02811f
C58 VP.n22 B 0.02811f
C59 VP.n23 B 0.02811f
C60 VP.n24 B 0.041035f
C61 VP.n25 B 0.05239f
C62 VP.n26 B 0.036611f
C63 VP.n27 B 0.02811f
C64 VP.n28 B 0.02811f
C65 VP.n29 B 0.042301f
C66 VP.n30 B 0.05449f
C67 VP.n31 B 0.030699f
C68 VP.n32 B 0.02811f
C69 VP.n33 B 0.02811f
C70 VP.n34 B 0.02811f
C71 VP.n35 B 0.05239f
C72 VP.n36 B 0.03092f
C73 VP.n37 B 0.356605f
C74 VP.n38 B 1.30505f
C75 VP.t7 B 0.672902f
C76 VP.n39 B 0.356605f
C77 VP.n40 B 1.32785f
C78 VP.n41 B 0.03706f
C79 VP.n42 B 0.02811f
C80 VP.n43 B 0.05239f
C81 VP.n44 B 0.049271f
C82 VP.n45 B 0.030699f
C83 VP.n46 B 0.02811f
C84 VP.n47 B 0.02811f
C85 VP.n48 B 0.02811f
C86 VP.n49 B 0.042301f
C87 VP.n50 B 0.272571f
C88 VP.n51 B 0.036611f
C89 VP.n52 B 0.05239f
C90 VP.n53 B 0.02811f
C91 VP.n54 B 0.02811f
C92 VP.n55 B 0.02811f
C93 VP.n56 B 0.041035f
C94 VP.n57 B 0.05239f
C95 VP.n58 B 0.036611f
C96 VP.n59 B 0.02811f
C97 VP.n60 B 0.02811f
C98 VP.n61 B 0.042301f
C99 VP.n62 B 0.05449f
C100 VP.n63 B 0.030699f
C101 VP.n64 B 0.02811f
C102 VP.n65 B 0.02811f
C103 VP.n66 B 0.02811f
C104 VP.n67 B 0.05239f
C105 VP.n68 B 0.03092f
C106 VP.n69 B 0.356605f
C107 VP.n70 B 0.04905f
C108 VDD2.t5 B 0.070492f
C109 VDD2.t7 B 0.070492f
C110 VDD2.n0 B 0.551476f
C111 VDD2.t2 B 0.070492f
C112 VDD2.t1 B 0.070492f
C113 VDD2.n1 B 0.551476f
C114 VDD2.n2 B 2.64958f
C115 VDD2.t4 B 0.070492f
C116 VDD2.t6 B 0.070492f
C117 VDD2.n3 B 0.544253f
C118 VDD2.n4 B 2.21364f
C119 VDD2.t0 B 0.070492f
C120 VDD2.t3 B 0.070492f
C121 VDD2.n5 B 0.551448f
C122 VTAIL.t7 B 0.076521f
C123 VTAIL.t8 B 0.076521f
C124 VTAIL.n0 B 0.537465f
C125 VTAIL.n1 B 0.438682f
C126 VTAIL.t12 B 0.692842f
C127 VTAIL.n2 B 0.526996f
C128 VTAIL.t0 B 0.692842f
C129 VTAIL.n3 B 0.526996f
C130 VTAIL.t2 B 0.076521f
C131 VTAIL.t4 B 0.076521f
C132 VTAIL.n4 B 0.537465f
C133 VTAIL.n5 B 0.64555f
C134 VTAIL.t6 B 0.692842f
C135 VTAIL.n6 B 1.32626f
C136 VTAIL.t13 B 0.692846f
C137 VTAIL.n7 B 1.32626f
C138 VTAIL.t11 B 0.076521f
C139 VTAIL.t10 B 0.076521f
C140 VTAIL.n8 B 0.537468f
C141 VTAIL.n9 B 0.645547f
C142 VTAIL.t14 B 0.692846f
C143 VTAIL.n10 B 0.526992f
C144 VTAIL.t3 B 0.692846f
C145 VTAIL.n11 B 0.526992f
C146 VTAIL.t1 B 0.076521f
C147 VTAIL.t15 B 0.076521f
C148 VTAIL.n12 B 0.537468f
C149 VTAIL.n13 B 0.645547f
C150 VTAIL.t5 B 0.692842f
C151 VTAIL.n14 B 1.32626f
C152 VTAIL.t9 B 0.692842f
C153 VTAIL.n15 B 1.32132f
C154 VN.n0 B 0.036117f
C155 VN.t6 B 0.655775f
C156 VN.n1 B 0.048017f
C157 VN.n2 B 0.027394f
C158 VN.t5 B 0.655775f
C159 VN.n3 B 0.265633f
C160 VN.n4 B 0.027394f
C161 VN.n5 B 0.039991f
C162 VN.n6 B 0.263138f
C163 VN.t0 B 0.655775f
C164 VN.t2 B 0.862052f
C165 VN.n7 B 0.333763f
C166 VN.n8 B 0.341396f
C167 VN.n9 B 0.035679f
C168 VN.n10 B 0.051056f
C169 VN.n11 B 0.027394f
C170 VN.n12 B 0.027394f
C171 VN.n13 B 0.027394f
C172 VN.n14 B 0.039991f
C173 VN.n15 B 0.051056f
C174 VN.n16 B 0.035679f
C175 VN.n17 B 0.027394f
C176 VN.n18 B 0.027394f
C177 VN.n19 B 0.041224f
C178 VN.n20 B 0.053103f
C179 VN.n21 B 0.029918f
C180 VN.n22 B 0.027394f
C181 VN.n23 B 0.027394f
C182 VN.n24 B 0.027394f
C183 VN.n25 B 0.051056f
C184 VN.n26 B 0.030133f
C185 VN.n27 B 0.347529f
C186 VN.n28 B 0.047802f
C187 VN.n29 B 0.036117f
C188 VN.t3 B 0.655775f
C189 VN.n30 B 0.048017f
C190 VN.n31 B 0.027394f
C191 VN.t1 B 0.655775f
C192 VN.n32 B 0.265633f
C193 VN.n33 B 0.027394f
C194 VN.n34 B 0.039991f
C195 VN.n35 B 0.263138f
C196 VN.t7 B 0.655775f
C197 VN.t4 B 0.862052f
C198 VN.n36 B 0.333763f
C199 VN.n37 B 0.341396f
C200 VN.n38 B 0.035679f
C201 VN.n39 B 0.051056f
C202 VN.n40 B 0.027394f
C203 VN.n41 B 0.027394f
C204 VN.n42 B 0.027394f
C205 VN.n43 B 0.039991f
C206 VN.n44 B 0.051056f
C207 VN.n45 B 0.035679f
C208 VN.n46 B 0.027394f
C209 VN.n47 B 0.027394f
C210 VN.n48 B 0.041224f
C211 VN.n49 B 0.053103f
C212 VN.n50 B 0.029918f
C213 VN.n51 B 0.027394f
C214 VN.n52 B 0.027394f
C215 VN.n53 B 0.027394f
C216 VN.n54 B 0.051056f
C217 VN.n55 B 0.030133f
C218 VN.n56 B 0.347529f
C219 VN.n57 B 1.28686f
.ends

