* NGSPICE file created from diff_pair_sample_0085.ext - technology: sky130A

.subckt diff_pair_sample_0085 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t3 VN.t0 VTAIL.t7 w_n3058_n4482# sky130_fd_pr__pfet_01v8 ad=2.89905 pd=17.9 as=6.8523 ps=35.92 w=17.57 l=3.15
X1 VTAIL.t1 VP.t0 VDD1.t3 w_n3058_n4482# sky130_fd_pr__pfet_01v8 ad=6.8523 pd=35.92 as=2.89905 ps=17.9 w=17.57 l=3.15
X2 B.t11 B.t9 B.t10 w_n3058_n4482# sky130_fd_pr__pfet_01v8 ad=6.8523 pd=35.92 as=0 ps=0 w=17.57 l=3.15
X3 VDD2.t2 VN.t1 VTAIL.t5 w_n3058_n4482# sky130_fd_pr__pfet_01v8 ad=2.89905 pd=17.9 as=6.8523 ps=35.92 w=17.57 l=3.15
X4 VDD1.t2 VP.t1 VTAIL.t3 w_n3058_n4482# sky130_fd_pr__pfet_01v8 ad=2.89905 pd=17.9 as=6.8523 ps=35.92 w=17.57 l=3.15
X5 VTAIL.t4 VN.t2 VDD2.t1 w_n3058_n4482# sky130_fd_pr__pfet_01v8 ad=6.8523 pd=35.92 as=2.89905 ps=17.9 w=17.57 l=3.15
X6 B.t8 B.t6 B.t7 w_n3058_n4482# sky130_fd_pr__pfet_01v8 ad=6.8523 pd=35.92 as=0 ps=0 w=17.57 l=3.15
X7 B.t5 B.t3 B.t4 w_n3058_n4482# sky130_fd_pr__pfet_01v8 ad=6.8523 pd=35.92 as=0 ps=0 w=17.57 l=3.15
X8 B.t2 B.t0 B.t1 w_n3058_n4482# sky130_fd_pr__pfet_01v8 ad=6.8523 pd=35.92 as=0 ps=0 w=17.57 l=3.15
X9 VTAIL.t6 VN.t3 VDD2.t0 w_n3058_n4482# sky130_fd_pr__pfet_01v8 ad=6.8523 pd=35.92 as=2.89905 ps=17.9 w=17.57 l=3.15
X10 VTAIL.t0 VP.t2 VDD1.t1 w_n3058_n4482# sky130_fd_pr__pfet_01v8 ad=6.8523 pd=35.92 as=2.89905 ps=17.9 w=17.57 l=3.15
X11 VDD1.t0 VP.t3 VTAIL.t2 w_n3058_n4482# sky130_fd_pr__pfet_01v8 ad=2.89905 pd=17.9 as=6.8523 ps=35.92 w=17.57 l=3.15
R0 VN.n1 VN.t1 168.899
R1 VN.n0 VN.t2 168.899
R2 VN.n0 VN.t0 167.815
R3 VN.n1 VN.t3 167.815
R4 VN VN.n1 55.0359
R5 VN VN.n0 2.69121
R6 VTAIL.n778 VTAIL.n686 756.745
R7 VTAIL.n92 VTAIL.n0 756.745
R8 VTAIL.n190 VTAIL.n98 756.745
R9 VTAIL.n288 VTAIL.n196 756.745
R10 VTAIL.n680 VTAIL.n588 756.745
R11 VTAIL.n582 VTAIL.n490 756.745
R12 VTAIL.n484 VTAIL.n392 756.745
R13 VTAIL.n386 VTAIL.n294 756.745
R14 VTAIL.n719 VTAIL.n718 585
R15 VTAIL.n721 VTAIL.n720 585
R16 VTAIL.n714 VTAIL.n713 585
R17 VTAIL.n727 VTAIL.n726 585
R18 VTAIL.n729 VTAIL.n728 585
R19 VTAIL.n710 VTAIL.n709 585
R20 VTAIL.n735 VTAIL.n734 585
R21 VTAIL.n737 VTAIL.n736 585
R22 VTAIL.n706 VTAIL.n705 585
R23 VTAIL.n743 VTAIL.n742 585
R24 VTAIL.n745 VTAIL.n744 585
R25 VTAIL.n702 VTAIL.n701 585
R26 VTAIL.n751 VTAIL.n750 585
R27 VTAIL.n753 VTAIL.n752 585
R28 VTAIL.n698 VTAIL.n697 585
R29 VTAIL.n760 VTAIL.n759 585
R30 VTAIL.n761 VTAIL.n696 585
R31 VTAIL.n763 VTAIL.n762 585
R32 VTAIL.n694 VTAIL.n693 585
R33 VTAIL.n769 VTAIL.n768 585
R34 VTAIL.n771 VTAIL.n770 585
R35 VTAIL.n690 VTAIL.n689 585
R36 VTAIL.n777 VTAIL.n776 585
R37 VTAIL.n779 VTAIL.n778 585
R38 VTAIL.n33 VTAIL.n32 585
R39 VTAIL.n35 VTAIL.n34 585
R40 VTAIL.n28 VTAIL.n27 585
R41 VTAIL.n41 VTAIL.n40 585
R42 VTAIL.n43 VTAIL.n42 585
R43 VTAIL.n24 VTAIL.n23 585
R44 VTAIL.n49 VTAIL.n48 585
R45 VTAIL.n51 VTAIL.n50 585
R46 VTAIL.n20 VTAIL.n19 585
R47 VTAIL.n57 VTAIL.n56 585
R48 VTAIL.n59 VTAIL.n58 585
R49 VTAIL.n16 VTAIL.n15 585
R50 VTAIL.n65 VTAIL.n64 585
R51 VTAIL.n67 VTAIL.n66 585
R52 VTAIL.n12 VTAIL.n11 585
R53 VTAIL.n74 VTAIL.n73 585
R54 VTAIL.n75 VTAIL.n10 585
R55 VTAIL.n77 VTAIL.n76 585
R56 VTAIL.n8 VTAIL.n7 585
R57 VTAIL.n83 VTAIL.n82 585
R58 VTAIL.n85 VTAIL.n84 585
R59 VTAIL.n4 VTAIL.n3 585
R60 VTAIL.n91 VTAIL.n90 585
R61 VTAIL.n93 VTAIL.n92 585
R62 VTAIL.n131 VTAIL.n130 585
R63 VTAIL.n133 VTAIL.n132 585
R64 VTAIL.n126 VTAIL.n125 585
R65 VTAIL.n139 VTAIL.n138 585
R66 VTAIL.n141 VTAIL.n140 585
R67 VTAIL.n122 VTAIL.n121 585
R68 VTAIL.n147 VTAIL.n146 585
R69 VTAIL.n149 VTAIL.n148 585
R70 VTAIL.n118 VTAIL.n117 585
R71 VTAIL.n155 VTAIL.n154 585
R72 VTAIL.n157 VTAIL.n156 585
R73 VTAIL.n114 VTAIL.n113 585
R74 VTAIL.n163 VTAIL.n162 585
R75 VTAIL.n165 VTAIL.n164 585
R76 VTAIL.n110 VTAIL.n109 585
R77 VTAIL.n172 VTAIL.n171 585
R78 VTAIL.n173 VTAIL.n108 585
R79 VTAIL.n175 VTAIL.n174 585
R80 VTAIL.n106 VTAIL.n105 585
R81 VTAIL.n181 VTAIL.n180 585
R82 VTAIL.n183 VTAIL.n182 585
R83 VTAIL.n102 VTAIL.n101 585
R84 VTAIL.n189 VTAIL.n188 585
R85 VTAIL.n191 VTAIL.n190 585
R86 VTAIL.n229 VTAIL.n228 585
R87 VTAIL.n231 VTAIL.n230 585
R88 VTAIL.n224 VTAIL.n223 585
R89 VTAIL.n237 VTAIL.n236 585
R90 VTAIL.n239 VTAIL.n238 585
R91 VTAIL.n220 VTAIL.n219 585
R92 VTAIL.n245 VTAIL.n244 585
R93 VTAIL.n247 VTAIL.n246 585
R94 VTAIL.n216 VTAIL.n215 585
R95 VTAIL.n253 VTAIL.n252 585
R96 VTAIL.n255 VTAIL.n254 585
R97 VTAIL.n212 VTAIL.n211 585
R98 VTAIL.n261 VTAIL.n260 585
R99 VTAIL.n263 VTAIL.n262 585
R100 VTAIL.n208 VTAIL.n207 585
R101 VTAIL.n270 VTAIL.n269 585
R102 VTAIL.n271 VTAIL.n206 585
R103 VTAIL.n273 VTAIL.n272 585
R104 VTAIL.n204 VTAIL.n203 585
R105 VTAIL.n279 VTAIL.n278 585
R106 VTAIL.n281 VTAIL.n280 585
R107 VTAIL.n200 VTAIL.n199 585
R108 VTAIL.n287 VTAIL.n286 585
R109 VTAIL.n289 VTAIL.n288 585
R110 VTAIL.n681 VTAIL.n680 585
R111 VTAIL.n679 VTAIL.n678 585
R112 VTAIL.n592 VTAIL.n591 585
R113 VTAIL.n673 VTAIL.n672 585
R114 VTAIL.n671 VTAIL.n670 585
R115 VTAIL.n596 VTAIL.n595 585
R116 VTAIL.n600 VTAIL.n598 585
R117 VTAIL.n665 VTAIL.n664 585
R118 VTAIL.n663 VTAIL.n662 585
R119 VTAIL.n602 VTAIL.n601 585
R120 VTAIL.n657 VTAIL.n656 585
R121 VTAIL.n655 VTAIL.n654 585
R122 VTAIL.n606 VTAIL.n605 585
R123 VTAIL.n649 VTAIL.n648 585
R124 VTAIL.n647 VTAIL.n646 585
R125 VTAIL.n610 VTAIL.n609 585
R126 VTAIL.n641 VTAIL.n640 585
R127 VTAIL.n639 VTAIL.n638 585
R128 VTAIL.n614 VTAIL.n613 585
R129 VTAIL.n633 VTAIL.n632 585
R130 VTAIL.n631 VTAIL.n630 585
R131 VTAIL.n618 VTAIL.n617 585
R132 VTAIL.n625 VTAIL.n624 585
R133 VTAIL.n623 VTAIL.n622 585
R134 VTAIL.n583 VTAIL.n582 585
R135 VTAIL.n581 VTAIL.n580 585
R136 VTAIL.n494 VTAIL.n493 585
R137 VTAIL.n575 VTAIL.n574 585
R138 VTAIL.n573 VTAIL.n572 585
R139 VTAIL.n498 VTAIL.n497 585
R140 VTAIL.n502 VTAIL.n500 585
R141 VTAIL.n567 VTAIL.n566 585
R142 VTAIL.n565 VTAIL.n564 585
R143 VTAIL.n504 VTAIL.n503 585
R144 VTAIL.n559 VTAIL.n558 585
R145 VTAIL.n557 VTAIL.n556 585
R146 VTAIL.n508 VTAIL.n507 585
R147 VTAIL.n551 VTAIL.n550 585
R148 VTAIL.n549 VTAIL.n548 585
R149 VTAIL.n512 VTAIL.n511 585
R150 VTAIL.n543 VTAIL.n542 585
R151 VTAIL.n541 VTAIL.n540 585
R152 VTAIL.n516 VTAIL.n515 585
R153 VTAIL.n535 VTAIL.n534 585
R154 VTAIL.n533 VTAIL.n532 585
R155 VTAIL.n520 VTAIL.n519 585
R156 VTAIL.n527 VTAIL.n526 585
R157 VTAIL.n525 VTAIL.n524 585
R158 VTAIL.n485 VTAIL.n484 585
R159 VTAIL.n483 VTAIL.n482 585
R160 VTAIL.n396 VTAIL.n395 585
R161 VTAIL.n477 VTAIL.n476 585
R162 VTAIL.n475 VTAIL.n474 585
R163 VTAIL.n400 VTAIL.n399 585
R164 VTAIL.n404 VTAIL.n402 585
R165 VTAIL.n469 VTAIL.n468 585
R166 VTAIL.n467 VTAIL.n466 585
R167 VTAIL.n406 VTAIL.n405 585
R168 VTAIL.n461 VTAIL.n460 585
R169 VTAIL.n459 VTAIL.n458 585
R170 VTAIL.n410 VTAIL.n409 585
R171 VTAIL.n453 VTAIL.n452 585
R172 VTAIL.n451 VTAIL.n450 585
R173 VTAIL.n414 VTAIL.n413 585
R174 VTAIL.n445 VTAIL.n444 585
R175 VTAIL.n443 VTAIL.n442 585
R176 VTAIL.n418 VTAIL.n417 585
R177 VTAIL.n437 VTAIL.n436 585
R178 VTAIL.n435 VTAIL.n434 585
R179 VTAIL.n422 VTAIL.n421 585
R180 VTAIL.n429 VTAIL.n428 585
R181 VTAIL.n427 VTAIL.n426 585
R182 VTAIL.n387 VTAIL.n386 585
R183 VTAIL.n385 VTAIL.n384 585
R184 VTAIL.n298 VTAIL.n297 585
R185 VTAIL.n379 VTAIL.n378 585
R186 VTAIL.n377 VTAIL.n376 585
R187 VTAIL.n302 VTAIL.n301 585
R188 VTAIL.n306 VTAIL.n304 585
R189 VTAIL.n371 VTAIL.n370 585
R190 VTAIL.n369 VTAIL.n368 585
R191 VTAIL.n308 VTAIL.n307 585
R192 VTAIL.n363 VTAIL.n362 585
R193 VTAIL.n361 VTAIL.n360 585
R194 VTAIL.n312 VTAIL.n311 585
R195 VTAIL.n355 VTAIL.n354 585
R196 VTAIL.n353 VTAIL.n352 585
R197 VTAIL.n316 VTAIL.n315 585
R198 VTAIL.n347 VTAIL.n346 585
R199 VTAIL.n345 VTAIL.n344 585
R200 VTAIL.n320 VTAIL.n319 585
R201 VTAIL.n339 VTAIL.n338 585
R202 VTAIL.n337 VTAIL.n336 585
R203 VTAIL.n324 VTAIL.n323 585
R204 VTAIL.n331 VTAIL.n330 585
R205 VTAIL.n329 VTAIL.n328 585
R206 VTAIL.n717 VTAIL.t7 327.466
R207 VTAIL.n31 VTAIL.t4 327.466
R208 VTAIL.n129 VTAIL.t3 327.466
R209 VTAIL.n227 VTAIL.t1 327.466
R210 VTAIL.n621 VTAIL.t2 327.466
R211 VTAIL.n523 VTAIL.t0 327.466
R212 VTAIL.n425 VTAIL.t5 327.466
R213 VTAIL.n327 VTAIL.t6 327.466
R214 VTAIL.n720 VTAIL.n719 171.744
R215 VTAIL.n720 VTAIL.n713 171.744
R216 VTAIL.n727 VTAIL.n713 171.744
R217 VTAIL.n728 VTAIL.n727 171.744
R218 VTAIL.n728 VTAIL.n709 171.744
R219 VTAIL.n735 VTAIL.n709 171.744
R220 VTAIL.n736 VTAIL.n735 171.744
R221 VTAIL.n736 VTAIL.n705 171.744
R222 VTAIL.n743 VTAIL.n705 171.744
R223 VTAIL.n744 VTAIL.n743 171.744
R224 VTAIL.n744 VTAIL.n701 171.744
R225 VTAIL.n751 VTAIL.n701 171.744
R226 VTAIL.n752 VTAIL.n751 171.744
R227 VTAIL.n752 VTAIL.n697 171.744
R228 VTAIL.n760 VTAIL.n697 171.744
R229 VTAIL.n761 VTAIL.n760 171.744
R230 VTAIL.n762 VTAIL.n761 171.744
R231 VTAIL.n762 VTAIL.n693 171.744
R232 VTAIL.n769 VTAIL.n693 171.744
R233 VTAIL.n770 VTAIL.n769 171.744
R234 VTAIL.n770 VTAIL.n689 171.744
R235 VTAIL.n777 VTAIL.n689 171.744
R236 VTAIL.n778 VTAIL.n777 171.744
R237 VTAIL.n34 VTAIL.n33 171.744
R238 VTAIL.n34 VTAIL.n27 171.744
R239 VTAIL.n41 VTAIL.n27 171.744
R240 VTAIL.n42 VTAIL.n41 171.744
R241 VTAIL.n42 VTAIL.n23 171.744
R242 VTAIL.n49 VTAIL.n23 171.744
R243 VTAIL.n50 VTAIL.n49 171.744
R244 VTAIL.n50 VTAIL.n19 171.744
R245 VTAIL.n57 VTAIL.n19 171.744
R246 VTAIL.n58 VTAIL.n57 171.744
R247 VTAIL.n58 VTAIL.n15 171.744
R248 VTAIL.n65 VTAIL.n15 171.744
R249 VTAIL.n66 VTAIL.n65 171.744
R250 VTAIL.n66 VTAIL.n11 171.744
R251 VTAIL.n74 VTAIL.n11 171.744
R252 VTAIL.n75 VTAIL.n74 171.744
R253 VTAIL.n76 VTAIL.n75 171.744
R254 VTAIL.n76 VTAIL.n7 171.744
R255 VTAIL.n83 VTAIL.n7 171.744
R256 VTAIL.n84 VTAIL.n83 171.744
R257 VTAIL.n84 VTAIL.n3 171.744
R258 VTAIL.n91 VTAIL.n3 171.744
R259 VTAIL.n92 VTAIL.n91 171.744
R260 VTAIL.n132 VTAIL.n131 171.744
R261 VTAIL.n132 VTAIL.n125 171.744
R262 VTAIL.n139 VTAIL.n125 171.744
R263 VTAIL.n140 VTAIL.n139 171.744
R264 VTAIL.n140 VTAIL.n121 171.744
R265 VTAIL.n147 VTAIL.n121 171.744
R266 VTAIL.n148 VTAIL.n147 171.744
R267 VTAIL.n148 VTAIL.n117 171.744
R268 VTAIL.n155 VTAIL.n117 171.744
R269 VTAIL.n156 VTAIL.n155 171.744
R270 VTAIL.n156 VTAIL.n113 171.744
R271 VTAIL.n163 VTAIL.n113 171.744
R272 VTAIL.n164 VTAIL.n163 171.744
R273 VTAIL.n164 VTAIL.n109 171.744
R274 VTAIL.n172 VTAIL.n109 171.744
R275 VTAIL.n173 VTAIL.n172 171.744
R276 VTAIL.n174 VTAIL.n173 171.744
R277 VTAIL.n174 VTAIL.n105 171.744
R278 VTAIL.n181 VTAIL.n105 171.744
R279 VTAIL.n182 VTAIL.n181 171.744
R280 VTAIL.n182 VTAIL.n101 171.744
R281 VTAIL.n189 VTAIL.n101 171.744
R282 VTAIL.n190 VTAIL.n189 171.744
R283 VTAIL.n230 VTAIL.n229 171.744
R284 VTAIL.n230 VTAIL.n223 171.744
R285 VTAIL.n237 VTAIL.n223 171.744
R286 VTAIL.n238 VTAIL.n237 171.744
R287 VTAIL.n238 VTAIL.n219 171.744
R288 VTAIL.n245 VTAIL.n219 171.744
R289 VTAIL.n246 VTAIL.n245 171.744
R290 VTAIL.n246 VTAIL.n215 171.744
R291 VTAIL.n253 VTAIL.n215 171.744
R292 VTAIL.n254 VTAIL.n253 171.744
R293 VTAIL.n254 VTAIL.n211 171.744
R294 VTAIL.n261 VTAIL.n211 171.744
R295 VTAIL.n262 VTAIL.n261 171.744
R296 VTAIL.n262 VTAIL.n207 171.744
R297 VTAIL.n270 VTAIL.n207 171.744
R298 VTAIL.n271 VTAIL.n270 171.744
R299 VTAIL.n272 VTAIL.n271 171.744
R300 VTAIL.n272 VTAIL.n203 171.744
R301 VTAIL.n279 VTAIL.n203 171.744
R302 VTAIL.n280 VTAIL.n279 171.744
R303 VTAIL.n280 VTAIL.n199 171.744
R304 VTAIL.n287 VTAIL.n199 171.744
R305 VTAIL.n288 VTAIL.n287 171.744
R306 VTAIL.n680 VTAIL.n679 171.744
R307 VTAIL.n679 VTAIL.n591 171.744
R308 VTAIL.n672 VTAIL.n591 171.744
R309 VTAIL.n672 VTAIL.n671 171.744
R310 VTAIL.n671 VTAIL.n595 171.744
R311 VTAIL.n600 VTAIL.n595 171.744
R312 VTAIL.n664 VTAIL.n600 171.744
R313 VTAIL.n664 VTAIL.n663 171.744
R314 VTAIL.n663 VTAIL.n601 171.744
R315 VTAIL.n656 VTAIL.n601 171.744
R316 VTAIL.n656 VTAIL.n655 171.744
R317 VTAIL.n655 VTAIL.n605 171.744
R318 VTAIL.n648 VTAIL.n605 171.744
R319 VTAIL.n648 VTAIL.n647 171.744
R320 VTAIL.n647 VTAIL.n609 171.744
R321 VTAIL.n640 VTAIL.n609 171.744
R322 VTAIL.n640 VTAIL.n639 171.744
R323 VTAIL.n639 VTAIL.n613 171.744
R324 VTAIL.n632 VTAIL.n613 171.744
R325 VTAIL.n632 VTAIL.n631 171.744
R326 VTAIL.n631 VTAIL.n617 171.744
R327 VTAIL.n624 VTAIL.n617 171.744
R328 VTAIL.n624 VTAIL.n623 171.744
R329 VTAIL.n582 VTAIL.n581 171.744
R330 VTAIL.n581 VTAIL.n493 171.744
R331 VTAIL.n574 VTAIL.n493 171.744
R332 VTAIL.n574 VTAIL.n573 171.744
R333 VTAIL.n573 VTAIL.n497 171.744
R334 VTAIL.n502 VTAIL.n497 171.744
R335 VTAIL.n566 VTAIL.n502 171.744
R336 VTAIL.n566 VTAIL.n565 171.744
R337 VTAIL.n565 VTAIL.n503 171.744
R338 VTAIL.n558 VTAIL.n503 171.744
R339 VTAIL.n558 VTAIL.n557 171.744
R340 VTAIL.n557 VTAIL.n507 171.744
R341 VTAIL.n550 VTAIL.n507 171.744
R342 VTAIL.n550 VTAIL.n549 171.744
R343 VTAIL.n549 VTAIL.n511 171.744
R344 VTAIL.n542 VTAIL.n511 171.744
R345 VTAIL.n542 VTAIL.n541 171.744
R346 VTAIL.n541 VTAIL.n515 171.744
R347 VTAIL.n534 VTAIL.n515 171.744
R348 VTAIL.n534 VTAIL.n533 171.744
R349 VTAIL.n533 VTAIL.n519 171.744
R350 VTAIL.n526 VTAIL.n519 171.744
R351 VTAIL.n526 VTAIL.n525 171.744
R352 VTAIL.n484 VTAIL.n483 171.744
R353 VTAIL.n483 VTAIL.n395 171.744
R354 VTAIL.n476 VTAIL.n395 171.744
R355 VTAIL.n476 VTAIL.n475 171.744
R356 VTAIL.n475 VTAIL.n399 171.744
R357 VTAIL.n404 VTAIL.n399 171.744
R358 VTAIL.n468 VTAIL.n404 171.744
R359 VTAIL.n468 VTAIL.n467 171.744
R360 VTAIL.n467 VTAIL.n405 171.744
R361 VTAIL.n460 VTAIL.n405 171.744
R362 VTAIL.n460 VTAIL.n459 171.744
R363 VTAIL.n459 VTAIL.n409 171.744
R364 VTAIL.n452 VTAIL.n409 171.744
R365 VTAIL.n452 VTAIL.n451 171.744
R366 VTAIL.n451 VTAIL.n413 171.744
R367 VTAIL.n444 VTAIL.n413 171.744
R368 VTAIL.n444 VTAIL.n443 171.744
R369 VTAIL.n443 VTAIL.n417 171.744
R370 VTAIL.n436 VTAIL.n417 171.744
R371 VTAIL.n436 VTAIL.n435 171.744
R372 VTAIL.n435 VTAIL.n421 171.744
R373 VTAIL.n428 VTAIL.n421 171.744
R374 VTAIL.n428 VTAIL.n427 171.744
R375 VTAIL.n386 VTAIL.n385 171.744
R376 VTAIL.n385 VTAIL.n297 171.744
R377 VTAIL.n378 VTAIL.n297 171.744
R378 VTAIL.n378 VTAIL.n377 171.744
R379 VTAIL.n377 VTAIL.n301 171.744
R380 VTAIL.n306 VTAIL.n301 171.744
R381 VTAIL.n370 VTAIL.n306 171.744
R382 VTAIL.n370 VTAIL.n369 171.744
R383 VTAIL.n369 VTAIL.n307 171.744
R384 VTAIL.n362 VTAIL.n307 171.744
R385 VTAIL.n362 VTAIL.n361 171.744
R386 VTAIL.n361 VTAIL.n311 171.744
R387 VTAIL.n354 VTAIL.n311 171.744
R388 VTAIL.n354 VTAIL.n353 171.744
R389 VTAIL.n353 VTAIL.n315 171.744
R390 VTAIL.n346 VTAIL.n315 171.744
R391 VTAIL.n346 VTAIL.n345 171.744
R392 VTAIL.n345 VTAIL.n319 171.744
R393 VTAIL.n338 VTAIL.n319 171.744
R394 VTAIL.n338 VTAIL.n337 171.744
R395 VTAIL.n337 VTAIL.n323 171.744
R396 VTAIL.n330 VTAIL.n323 171.744
R397 VTAIL.n330 VTAIL.n329 171.744
R398 VTAIL.n719 VTAIL.t7 85.8723
R399 VTAIL.n33 VTAIL.t4 85.8723
R400 VTAIL.n131 VTAIL.t3 85.8723
R401 VTAIL.n229 VTAIL.t1 85.8723
R402 VTAIL.n623 VTAIL.t2 85.8723
R403 VTAIL.n525 VTAIL.t0 85.8723
R404 VTAIL.n427 VTAIL.t5 85.8723
R405 VTAIL.n329 VTAIL.t6 85.8723
R406 VTAIL.n783 VTAIL.n782 33.155
R407 VTAIL.n97 VTAIL.n96 33.155
R408 VTAIL.n195 VTAIL.n194 33.155
R409 VTAIL.n293 VTAIL.n292 33.155
R410 VTAIL.n685 VTAIL.n684 33.155
R411 VTAIL.n587 VTAIL.n586 33.155
R412 VTAIL.n489 VTAIL.n488 33.155
R413 VTAIL.n391 VTAIL.n390 33.155
R414 VTAIL.n783 VTAIL.n685 30.5134
R415 VTAIL.n391 VTAIL.n293 30.5134
R416 VTAIL.n718 VTAIL.n717 16.3895
R417 VTAIL.n32 VTAIL.n31 16.3895
R418 VTAIL.n130 VTAIL.n129 16.3895
R419 VTAIL.n228 VTAIL.n227 16.3895
R420 VTAIL.n622 VTAIL.n621 16.3895
R421 VTAIL.n524 VTAIL.n523 16.3895
R422 VTAIL.n426 VTAIL.n425 16.3895
R423 VTAIL.n328 VTAIL.n327 16.3895
R424 VTAIL.n763 VTAIL.n694 13.1884
R425 VTAIL.n77 VTAIL.n8 13.1884
R426 VTAIL.n175 VTAIL.n106 13.1884
R427 VTAIL.n273 VTAIL.n204 13.1884
R428 VTAIL.n598 VTAIL.n596 13.1884
R429 VTAIL.n500 VTAIL.n498 13.1884
R430 VTAIL.n402 VTAIL.n400 13.1884
R431 VTAIL.n304 VTAIL.n302 13.1884
R432 VTAIL.n721 VTAIL.n716 12.8005
R433 VTAIL.n764 VTAIL.n696 12.8005
R434 VTAIL.n768 VTAIL.n767 12.8005
R435 VTAIL.n35 VTAIL.n30 12.8005
R436 VTAIL.n78 VTAIL.n10 12.8005
R437 VTAIL.n82 VTAIL.n81 12.8005
R438 VTAIL.n133 VTAIL.n128 12.8005
R439 VTAIL.n176 VTAIL.n108 12.8005
R440 VTAIL.n180 VTAIL.n179 12.8005
R441 VTAIL.n231 VTAIL.n226 12.8005
R442 VTAIL.n274 VTAIL.n206 12.8005
R443 VTAIL.n278 VTAIL.n277 12.8005
R444 VTAIL.n670 VTAIL.n669 12.8005
R445 VTAIL.n666 VTAIL.n665 12.8005
R446 VTAIL.n625 VTAIL.n620 12.8005
R447 VTAIL.n572 VTAIL.n571 12.8005
R448 VTAIL.n568 VTAIL.n567 12.8005
R449 VTAIL.n527 VTAIL.n522 12.8005
R450 VTAIL.n474 VTAIL.n473 12.8005
R451 VTAIL.n470 VTAIL.n469 12.8005
R452 VTAIL.n429 VTAIL.n424 12.8005
R453 VTAIL.n376 VTAIL.n375 12.8005
R454 VTAIL.n372 VTAIL.n371 12.8005
R455 VTAIL.n331 VTAIL.n326 12.8005
R456 VTAIL.n722 VTAIL.n714 12.0247
R457 VTAIL.n759 VTAIL.n758 12.0247
R458 VTAIL.n771 VTAIL.n692 12.0247
R459 VTAIL.n36 VTAIL.n28 12.0247
R460 VTAIL.n73 VTAIL.n72 12.0247
R461 VTAIL.n85 VTAIL.n6 12.0247
R462 VTAIL.n134 VTAIL.n126 12.0247
R463 VTAIL.n171 VTAIL.n170 12.0247
R464 VTAIL.n183 VTAIL.n104 12.0247
R465 VTAIL.n232 VTAIL.n224 12.0247
R466 VTAIL.n269 VTAIL.n268 12.0247
R467 VTAIL.n281 VTAIL.n202 12.0247
R468 VTAIL.n673 VTAIL.n594 12.0247
R469 VTAIL.n662 VTAIL.n599 12.0247
R470 VTAIL.n626 VTAIL.n618 12.0247
R471 VTAIL.n575 VTAIL.n496 12.0247
R472 VTAIL.n564 VTAIL.n501 12.0247
R473 VTAIL.n528 VTAIL.n520 12.0247
R474 VTAIL.n477 VTAIL.n398 12.0247
R475 VTAIL.n466 VTAIL.n403 12.0247
R476 VTAIL.n430 VTAIL.n422 12.0247
R477 VTAIL.n379 VTAIL.n300 12.0247
R478 VTAIL.n368 VTAIL.n305 12.0247
R479 VTAIL.n332 VTAIL.n324 12.0247
R480 VTAIL.n726 VTAIL.n725 11.249
R481 VTAIL.n757 VTAIL.n698 11.249
R482 VTAIL.n772 VTAIL.n690 11.249
R483 VTAIL.n40 VTAIL.n39 11.249
R484 VTAIL.n71 VTAIL.n12 11.249
R485 VTAIL.n86 VTAIL.n4 11.249
R486 VTAIL.n138 VTAIL.n137 11.249
R487 VTAIL.n169 VTAIL.n110 11.249
R488 VTAIL.n184 VTAIL.n102 11.249
R489 VTAIL.n236 VTAIL.n235 11.249
R490 VTAIL.n267 VTAIL.n208 11.249
R491 VTAIL.n282 VTAIL.n200 11.249
R492 VTAIL.n674 VTAIL.n592 11.249
R493 VTAIL.n661 VTAIL.n602 11.249
R494 VTAIL.n630 VTAIL.n629 11.249
R495 VTAIL.n576 VTAIL.n494 11.249
R496 VTAIL.n563 VTAIL.n504 11.249
R497 VTAIL.n532 VTAIL.n531 11.249
R498 VTAIL.n478 VTAIL.n396 11.249
R499 VTAIL.n465 VTAIL.n406 11.249
R500 VTAIL.n434 VTAIL.n433 11.249
R501 VTAIL.n380 VTAIL.n298 11.249
R502 VTAIL.n367 VTAIL.n308 11.249
R503 VTAIL.n336 VTAIL.n335 11.249
R504 VTAIL.n729 VTAIL.n712 10.4732
R505 VTAIL.n754 VTAIL.n753 10.4732
R506 VTAIL.n776 VTAIL.n775 10.4732
R507 VTAIL.n43 VTAIL.n26 10.4732
R508 VTAIL.n68 VTAIL.n67 10.4732
R509 VTAIL.n90 VTAIL.n89 10.4732
R510 VTAIL.n141 VTAIL.n124 10.4732
R511 VTAIL.n166 VTAIL.n165 10.4732
R512 VTAIL.n188 VTAIL.n187 10.4732
R513 VTAIL.n239 VTAIL.n222 10.4732
R514 VTAIL.n264 VTAIL.n263 10.4732
R515 VTAIL.n286 VTAIL.n285 10.4732
R516 VTAIL.n678 VTAIL.n677 10.4732
R517 VTAIL.n658 VTAIL.n657 10.4732
R518 VTAIL.n633 VTAIL.n616 10.4732
R519 VTAIL.n580 VTAIL.n579 10.4732
R520 VTAIL.n560 VTAIL.n559 10.4732
R521 VTAIL.n535 VTAIL.n518 10.4732
R522 VTAIL.n482 VTAIL.n481 10.4732
R523 VTAIL.n462 VTAIL.n461 10.4732
R524 VTAIL.n437 VTAIL.n420 10.4732
R525 VTAIL.n384 VTAIL.n383 10.4732
R526 VTAIL.n364 VTAIL.n363 10.4732
R527 VTAIL.n339 VTAIL.n322 10.4732
R528 VTAIL.n730 VTAIL.n710 9.69747
R529 VTAIL.n750 VTAIL.n700 9.69747
R530 VTAIL.n779 VTAIL.n688 9.69747
R531 VTAIL.n44 VTAIL.n24 9.69747
R532 VTAIL.n64 VTAIL.n14 9.69747
R533 VTAIL.n93 VTAIL.n2 9.69747
R534 VTAIL.n142 VTAIL.n122 9.69747
R535 VTAIL.n162 VTAIL.n112 9.69747
R536 VTAIL.n191 VTAIL.n100 9.69747
R537 VTAIL.n240 VTAIL.n220 9.69747
R538 VTAIL.n260 VTAIL.n210 9.69747
R539 VTAIL.n289 VTAIL.n198 9.69747
R540 VTAIL.n681 VTAIL.n590 9.69747
R541 VTAIL.n654 VTAIL.n604 9.69747
R542 VTAIL.n634 VTAIL.n614 9.69747
R543 VTAIL.n583 VTAIL.n492 9.69747
R544 VTAIL.n556 VTAIL.n506 9.69747
R545 VTAIL.n536 VTAIL.n516 9.69747
R546 VTAIL.n485 VTAIL.n394 9.69747
R547 VTAIL.n458 VTAIL.n408 9.69747
R548 VTAIL.n438 VTAIL.n418 9.69747
R549 VTAIL.n387 VTAIL.n296 9.69747
R550 VTAIL.n360 VTAIL.n310 9.69747
R551 VTAIL.n340 VTAIL.n320 9.69747
R552 VTAIL.n782 VTAIL.n781 9.45567
R553 VTAIL.n96 VTAIL.n95 9.45567
R554 VTAIL.n194 VTAIL.n193 9.45567
R555 VTAIL.n292 VTAIL.n291 9.45567
R556 VTAIL.n684 VTAIL.n683 9.45567
R557 VTAIL.n586 VTAIL.n585 9.45567
R558 VTAIL.n488 VTAIL.n487 9.45567
R559 VTAIL.n390 VTAIL.n389 9.45567
R560 VTAIL.n781 VTAIL.n780 9.3005
R561 VTAIL.n688 VTAIL.n687 9.3005
R562 VTAIL.n775 VTAIL.n774 9.3005
R563 VTAIL.n773 VTAIL.n772 9.3005
R564 VTAIL.n692 VTAIL.n691 9.3005
R565 VTAIL.n767 VTAIL.n766 9.3005
R566 VTAIL.n739 VTAIL.n738 9.3005
R567 VTAIL.n708 VTAIL.n707 9.3005
R568 VTAIL.n733 VTAIL.n732 9.3005
R569 VTAIL.n731 VTAIL.n730 9.3005
R570 VTAIL.n712 VTAIL.n711 9.3005
R571 VTAIL.n725 VTAIL.n724 9.3005
R572 VTAIL.n723 VTAIL.n722 9.3005
R573 VTAIL.n716 VTAIL.n715 9.3005
R574 VTAIL.n741 VTAIL.n740 9.3005
R575 VTAIL.n704 VTAIL.n703 9.3005
R576 VTAIL.n747 VTAIL.n746 9.3005
R577 VTAIL.n749 VTAIL.n748 9.3005
R578 VTAIL.n700 VTAIL.n699 9.3005
R579 VTAIL.n755 VTAIL.n754 9.3005
R580 VTAIL.n757 VTAIL.n756 9.3005
R581 VTAIL.n758 VTAIL.n695 9.3005
R582 VTAIL.n765 VTAIL.n764 9.3005
R583 VTAIL.n95 VTAIL.n94 9.3005
R584 VTAIL.n2 VTAIL.n1 9.3005
R585 VTAIL.n89 VTAIL.n88 9.3005
R586 VTAIL.n87 VTAIL.n86 9.3005
R587 VTAIL.n6 VTAIL.n5 9.3005
R588 VTAIL.n81 VTAIL.n80 9.3005
R589 VTAIL.n53 VTAIL.n52 9.3005
R590 VTAIL.n22 VTAIL.n21 9.3005
R591 VTAIL.n47 VTAIL.n46 9.3005
R592 VTAIL.n45 VTAIL.n44 9.3005
R593 VTAIL.n26 VTAIL.n25 9.3005
R594 VTAIL.n39 VTAIL.n38 9.3005
R595 VTAIL.n37 VTAIL.n36 9.3005
R596 VTAIL.n30 VTAIL.n29 9.3005
R597 VTAIL.n55 VTAIL.n54 9.3005
R598 VTAIL.n18 VTAIL.n17 9.3005
R599 VTAIL.n61 VTAIL.n60 9.3005
R600 VTAIL.n63 VTAIL.n62 9.3005
R601 VTAIL.n14 VTAIL.n13 9.3005
R602 VTAIL.n69 VTAIL.n68 9.3005
R603 VTAIL.n71 VTAIL.n70 9.3005
R604 VTAIL.n72 VTAIL.n9 9.3005
R605 VTAIL.n79 VTAIL.n78 9.3005
R606 VTAIL.n193 VTAIL.n192 9.3005
R607 VTAIL.n100 VTAIL.n99 9.3005
R608 VTAIL.n187 VTAIL.n186 9.3005
R609 VTAIL.n185 VTAIL.n184 9.3005
R610 VTAIL.n104 VTAIL.n103 9.3005
R611 VTAIL.n179 VTAIL.n178 9.3005
R612 VTAIL.n151 VTAIL.n150 9.3005
R613 VTAIL.n120 VTAIL.n119 9.3005
R614 VTAIL.n145 VTAIL.n144 9.3005
R615 VTAIL.n143 VTAIL.n142 9.3005
R616 VTAIL.n124 VTAIL.n123 9.3005
R617 VTAIL.n137 VTAIL.n136 9.3005
R618 VTAIL.n135 VTAIL.n134 9.3005
R619 VTAIL.n128 VTAIL.n127 9.3005
R620 VTAIL.n153 VTAIL.n152 9.3005
R621 VTAIL.n116 VTAIL.n115 9.3005
R622 VTAIL.n159 VTAIL.n158 9.3005
R623 VTAIL.n161 VTAIL.n160 9.3005
R624 VTAIL.n112 VTAIL.n111 9.3005
R625 VTAIL.n167 VTAIL.n166 9.3005
R626 VTAIL.n169 VTAIL.n168 9.3005
R627 VTAIL.n170 VTAIL.n107 9.3005
R628 VTAIL.n177 VTAIL.n176 9.3005
R629 VTAIL.n291 VTAIL.n290 9.3005
R630 VTAIL.n198 VTAIL.n197 9.3005
R631 VTAIL.n285 VTAIL.n284 9.3005
R632 VTAIL.n283 VTAIL.n282 9.3005
R633 VTAIL.n202 VTAIL.n201 9.3005
R634 VTAIL.n277 VTAIL.n276 9.3005
R635 VTAIL.n249 VTAIL.n248 9.3005
R636 VTAIL.n218 VTAIL.n217 9.3005
R637 VTAIL.n243 VTAIL.n242 9.3005
R638 VTAIL.n241 VTAIL.n240 9.3005
R639 VTAIL.n222 VTAIL.n221 9.3005
R640 VTAIL.n235 VTAIL.n234 9.3005
R641 VTAIL.n233 VTAIL.n232 9.3005
R642 VTAIL.n226 VTAIL.n225 9.3005
R643 VTAIL.n251 VTAIL.n250 9.3005
R644 VTAIL.n214 VTAIL.n213 9.3005
R645 VTAIL.n257 VTAIL.n256 9.3005
R646 VTAIL.n259 VTAIL.n258 9.3005
R647 VTAIL.n210 VTAIL.n209 9.3005
R648 VTAIL.n265 VTAIL.n264 9.3005
R649 VTAIL.n267 VTAIL.n266 9.3005
R650 VTAIL.n268 VTAIL.n205 9.3005
R651 VTAIL.n275 VTAIL.n274 9.3005
R652 VTAIL.n608 VTAIL.n607 9.3005
R653 VTAIL.n651 VTAIL.n650 9.3005
R654 VTAIL.n653 VTAIL.n652 9.3005
R655 VTAIL.n604 VTAIL.n603 9.3005
R656 VTAIL.n659 VTAIL.n658 9.3005
R657 VTAIL.n661 VTAIL.n660 9.3005
R658 VTAIL.n599 VTAIL.n597 9.3005
R659 VTAIL.n667 VTAIL.n666 9.3005
R660 VTAIL.n683 VTAIL.n682 9.3005
R661 VTAIL.n590 VTAIL.n589 9.3005
R662 VTAIL.n677 VTAIL.n676 9.3005
R663 VTAIL.n675 VTAIL.n674 9.3005
R664 VTAIL.n594 VTAIL.n593 9.3005
R665 VTAIL.n669 VTAIL.n668 9.3005
R666 VTAIL.n645 VTAIL.n644 9.3005
R667 VTAIL.n643 VTAIL.n642 9.3005
R668 VTAIL.n612 VTAIL.n611 9.3005
R669 VTAIL.n637 VTAIL.n636 9.3005
R670 VTAIL.n635 VTAIL.n634 9.3005
R671 VTAIL.n616 VTAIL.n615 9.3005
R672 VTAIL.n629 VTAIL.n628 9.3005
R673 VTAIL.n627 VTAIL.n626 9.3005
R674 VTAIL.n620 VTAIL.n619 9.3005
R675 VTAIL.n510 VTAIL.n509 9.3005
R676 VTAIL.n553 VTAIL.n552 9.3005
R677 VTAIL.n555 VTAIL.n554 9.3005
R678 VTAIL.n506 VTAIL.n505 9.3005
R679 VTAIL.n561 VTAIL.n560 9.3005
R680 VTAIL.n563 VTAIL.n562 9.3005
R681 VTAIL.n501 VTAIL.n499 9.3005
R682 VTAIL.n569 VTAIL.n568 9.3005
R683 VTAIL.n585 VTAIL.n584 9.3005
R684 VTAIL.n492 VTAIL.n491 9.3005
R685 VTAIL.n579 VTAIL.n578 9.3005
R686 VTAIL.n577 VTAIL.n576 9.3005
R687 VTAIL.n496 VTAIL.n495 9.3005
R688 VTAIL.n571 VTAIL.n570 9.3005
R689 VTAIL.n547 VTAIL.n546 9.3005
R690 VTAIL.n545 VTAIL.n544 9.3005
R691 VTAIL.n514 VTAIL.n513 9.3005
R692 VTAIL.n539 VTAIL.n538 9.3005
R693 VTAIL.n537 VTAIL.n536 9.3005
R694 VTAIL.n518 VTAIL.n517 9.3005
R695 VTAIL.n531 VTAIL.n530 9.3005
R696 VTAIL.n529 VTAIL.n528 9.3005
R697 VTAIL.n522 VTAIL.n521 9.3005
R698 VTAIL.n412 VTAIL.n411 9.3005
R699 VTAIL.n455 VTAIL.n454 9.3005
R700 VTAIL.n457 VTAIL.n456 9.3005
R701 VTAIL.n408 VTAIL.n407 9.3005
R702 VTAIL.n463 VTAIL.n462 9.3005
R703 VTAIL.n465 VTAIL.n464 9.3005
R704 VTAIL.n403 VTAIL.n401 9.3005
R705 VTAIL.n471 VTAIL.n470 9.3005
R706 VTAIL.n487 VTAIL.n486 9.3005
R707 VTAIL.n394 VTAIL.n393 9.3005
R708 VTAIL.n481 VTAIL.n480 9.3005
R709 VTAIL.n479 VTAIL.n478 9.3005
R710 VTAIL.n398 VTAIL.n397 9.3005
R711 VTAIL.n473 VTAIL.n472 9.3005
R712 VTAIL.n449 VTAIL.n448 9.3005
R713 VTAIL.n447 VTAIL.n446 9.3005
R714 VTAIL.n416 VTAIL.n415 9.3005
R715 VTAIL.n441 VTAIL.n440 9.3005
R716 VTAIL.n439 VTAIL.n438 9.3005
R717 VTAIL.n420 VTAIL.n419 9.3005
R718 VTAIL.n433 VTAIL.n432 9.3005
R719 VTAIL.n431 VTAIL.n430 9.3005
R720 VTAIL.n424 VTAIL.n423 9.3005
R721 VTAIL.n314 VTAIL.n313 9.3005
R722 VTAIL.n357 VTAIL.n356 9.3005
R723 VTAIL.n359 VTAIL.n358 9.3005
R724 VTAIL.n310 VTAIL.n309 9.3005
R725 VTAIL.n365 VTAIL.n364 9.3005
R726 VTAIL.n367 VTAIL.n366 9.3005
R727 VTAIL.n305 VTAIL.n303 9.3005
R728 VTAIL.n373 VTAIL.n372 9.3005
R729 VTAIL.n389 VTAIL.n388 9.3005
R730 VTAIL.n296 VTAIL.n295 9.3005
R731 VTAIL.n383 VTAIL.n382 9.3005
R732 VTAIL.n381 VTAIL.n380 9.3005
R733 VTAIL.n300 VTAIL.n299 9.3005
R734 VTAIL.n375 VTAIL.n374 9.3005
R735 VTAIL.n351 VTAIL.n350 9.3005
R736 VTAIL.n349 VTAIL.n348 9.3005
R737 VTAIL.n318 VTAIL.n317 9.3005
R738 VTAIL.n343 VTAIL.n342 9.3005
R739 VTAIL.n341 VTAIL.n340 9.3005
R740 VTAIL.n322 VTAIL.n321 9.3005
R741 VTAIL.n335 VTAIL.n334 9.3005
R742 VTAIL.n333 VTAIL.n332 9.3005
R743 VTAIL.n326 VTAIL.n325 9.3005
R744 VTAIL.n734 VTAIL.n733 8.92171
R745 VTAIL.n749 VTAIL.n702 8.92171
R746 VTAIL.n780 VTAIL.n686 8.92171
R747 VTAIL.n48 VTAIL.n47 8.92171
R748 VTAIL.n63 VTAIL.n16 8.92171
R749 VTAIL.n94 VTAIL.n0 8.92171
R750 VTAIL.n146 VTAIL.n145 8.92171
R751 VTAIL.n161 VTAIL.n114 8.92171
R752 VTAIL.n192 VTAIL.n98 8.92171
R753 VTAIL.n244 VTAIL.n243 8.92171
R754 VTAIL.n259 VTAIL.n212 8.92171
R755 VTAIL.n290 VTAIL.n196 8.92171
R756 VTAIL.n682 VTAIL.n588 8.92171
R757 VTAIL.n653 VTAIL.n606 8.92171
R758 VTAIL.n638 VTAIL.n637 8.92171
R759 VTAIL.n584 VTAIL.n490 8.92171
R760 VTAIL.n555 VTAIL.n508 8.92171
R761 VTAIL.n540 VTAIL.n539 8.92171
R762 VTAIL.n486 VTAIL.n392 8.92171
R763 VTAIL.n457 VTAIL.n410 8.92171
R764 VTAIL.n442 VTAIL.n441 8.92171
R765 VTAIL.n388 VTAIL.n294 8.92171
R766 VTAIL.n359 VTAIL.n312 8.92171
R767 VTAIL.n344 VTAIL.n343 8.92171
R768 VTAIL.n737 VTAIL.n708 8.14595
R769 VTAIL.n746 VTAIL.n745 8.14595
R770 VTAIL.n51 VTAIL.n22 8.14595
R771 VTAIL.n60 VTAIL.n59 8.14595
R772 VTAIL.n149 VTAIL.n120 8.14595
R773 VTAIL.n158 VTAIL.n157 8.14595
R774 VTAIL.n247 VTAIL.n218 8.14595
R775 VTAIL.n256 VTAIL.n255 8.14595
R776 VTAIL.n650 VTAIL.n649 8.14595
R777 VTAIL.n641 VTAIL.n612 8.14595
R778 VTAIL.n552 VTAIL.n551 8.14595
R779 VTAIL.n543 VTAIL.n514 8.14595
R780 VTAIL.n454 VTAIL.n453 8.14595
R781 VTAIL.n445 VTAIL.n416 8.14595
R782 VTAIL.n356 VTAIL.n355 8.14595
R783 VTAIL.n347 VTAIL.n318 8.14595
R784 VTAIL.n738 VTAIL.n706 7.3702
R785 VTAIL.n742 VTAIL.n704 7.3702
R786 VTAIL.n52 VTAIL.n20 7.3702
R787 VTAIL.n56 VTAIL.n18 7.3702
R788 VTAIL.n150 VTAIL.n118 7.3702
R789 VTAIL.n154 VTAIL.n116 7.3702
R790 VTAIL.n248 VTAIL.n216 7.3702
R791 VTAIL.n252 VTAIL.n214 7.3702
R792 VTAIL.n646 VTAIL.n608 7.3702
R793 VTAIL.n642 VTAIL.n610 7.3702
R794 VTAIL.n548 VTAIL.n510 7.3702
R795 VTAIL.n544 VTAIL.n512 7.3702
R796 VTAIL.n450 VTAIL.n412 7.3702
R797 VTAIL.n446 VTAIL.n414 7.3702
R798 VTAIL.n352 VTAIL.n314 7.3702
R799 VTAIL.n348 VTAIL.n316 7.3702
R800 VTAIL.n741 VTAIL.n706 6.59444
R801 VTAIL.n742 VTAIL.n741 6.59444
R802 VTAIL.n55 VTAIL.n20 6.59444
R803 VTAIL.n56 VTAIL.n55 6.59444
R804 VTAIL.n153 VTAIL.n118 6.59444
R805 VTAIL.n154 VTAIL.n153 6.59444
R806 VTAIL.n251 VTAIL.n216 6.59444
R807 VTAIL.n252 VTAIL.n251 6.59444
R808 VTAIL.n646 VTAIL.n645 6.59444
R809 VTAIL.n645 VTAIL.n610 6.59444
R810 VTAIL.n548 VTAIL.n547 6.59444
R811 VTAIL.n547 VTAIL.n512 6.59444
R812 VTAIL.n450 VTAIL.n449 6.59444
R813 VTAIL.n449 VTAIL.n414 6.59444
R814 VTAIL.n352 VTAIL.n351 6.59444
R815 VTAIL.n351 VTAIL.n316 6.59444
R816 VTAIL.n738 VTAIL.n737 5.81868
R817 VTAIL.n745 VTAIL.n704 5.81868
R818 VTAIL.n52 VTAIL.n51 5.81868
R819 VTAIL.n59 VTAIL.n18 5.81868
R820 VTAIL.n150 VTAIL.n149 5.81868
R821 VTAIL.n157 VTAIL.n116 5.81868
R822 VTAIL.n248 VTAIL.n247 5.81868
R823 VTAIL.n255 VTAIL.n214 5.81868
R824 VTAIL.n649 VTAIL.n608 5.81868
R825 VTAIL.n642 VTAIL.n641 5.81868
R826 VTAIL.n551 VTAIL.n510 5.81868
R827 VTAIL.n544 VTAIL.n543 5.81868
R828 VTAIL.n453 VTAIL.n412 5.81868
R829 VTAIL.n446 VTAIL.n445 5.81868
R830 VTAIL.n355 VTAIL.n314 5.81868
R831 VTAIL.n348 VTAIL.n347 5.81868
R832 VTAIL.n734 VTAIL.n708 5.04292
R833 VTAIL.n746 VTAIL.n702 5.04292
R834 VTAIL.n782 VTAIL.n686 5.04292
R835 VTAIL.n48 VTAIL.n22 5.04292
R836 VTAIL.n60 VTAIL.n16 5.04292
R837 VTAIL.n96 VTAIL.n0 5.04292
R838 VTAIL.n146 VTAIL.n120 5.04292
R839 VTAIL.n158 VTAIL.n114 5.04292
R840 VTAIL.n194 VTAIL.n98 5.04292
R841 VTAIL.n244 VTAIL.n218 5.04292
R842 VTAIL.n256 VTAIL.n212 5.04292
R843 VTAIL.n292 VTAIL.n196 5.04292
R844 VTAIL.n684 VTAIL.n588 5.04292
R845 VTAIL.n650 VTAIL.n606 5.04292
R846 VTAIL.n638 VTAIL.n612 5.04292
R847 VTAIL.n586 VTAIL.n490 5.04292
R848 VTAIL.n552 VTAIL.n508 5.04292
R849 VTAIL.n540 VTAIL.n514 5.04292
R850 VTAIL.n488 VTAIL.n392 5.04292
R851 VTAIL.n454 VTAIL.n410 5.04292
R852 VTAIL.n442 VTAIL.n416 5.04292
R853 VTAIL.n390 VTAIL.n294 5.04292
R854 VTAIL.n356 VTAIL.n312 5.04292
R855 VTAIL.n344 VTAIL.n318 5.04292
R856 VTAIL.n733 VTAIL.n710 4.26717
R857 VTAIL.n750 VTAIL.n749 4.26717
R858 VTAIL.n780 VTAIL.n779 4.26717
R859 VTAIL.n47 VTAIL.n24 4.26717
R860 VTAIL.n64 VTAIL.n63 4.26717
R861 VTAIL.n94 VTAIL.n93 4.26717
R862 VTAIL.n145 VTAIL.n122 4.26717
R863 VTAIL.n162 VTAIL.n161 4.26717
R864 VTAIL.n192 VTAIL.n191 4.26717
R865 VTAIL.n243 VTAIL.n220 4.26717
R866 VTAIL.n260 VTAIL.n259 4.26717
R867 VTAIL.n290 VTAIL.n289 4.26717
R868 VTAIL.n682 VTAIL.n681 4.26717
R869 VTAIL.n654 VTAIL.n653 4.26717
R870 VTAIL.n637 VTAIL.n614 4.26717
R871 VTAIL.n584 VTAIL.n583 4.26717
R872 VTAIL.n556 VTAIL.n555 4.26717
R873 VTAIL.n539 VTAIL.n516 4.26717
R874 VTAIL.n486 VTAIL.n485 4.26717
R875 VTAIL.n458 VTAIL.n457 4.26717
R876 VTAIL.n441 VTAIL.n418 4.26717
R877 VTAIL.n388 VTAIL.n387 4.26717
R878 VTAIL.n360 VTAIL.n359 4.26717
R879 VTAIL.n343 VTAIL.n320 4.26717
R880 VTAIL.n717 VTAIL.n715 3.70982
R881 VTAIL.n31 VTAIL.n29 3.70982
R882 VTAIL.n129 VTAIL.n127 3.70982
R883 VTAIL.n227 VTAIL.n225 3.70982
R884 VTAIL.n621 VTAIL.n619 3.70982
R885 VTAIL.n523 VTAIL.n521 3.70982
R886 VTAIL.n425 VTAIL.n423 3.70982
R887 VTAIL.n327 VTAIL.n325 3.70982
R888 VTAIL.n730 VTAIL.n729 3.49141
R889 VTAIL.n753 VTAIL.n700 3.49141
R890 VTAIL.n776 VTAIL.n688 3.49141
R891 VTAIL.n44 VTAIL.n43 3.49141
R892 VTAIL.n67 VTAIL.n14 3.49141
R893 VTAIL.n90 VTAIL.n2 3.49141
R894 VTAIL.n142 VTAIL.n141 3.49141
R895 VTAIL.n165 VTAIL.n112 3.49141
R896 VTAIL.n188 VTAIL.n100 3.49141
R897 VTAIL.n240 VTAIL.n239 3.49141
R898 VTAIL.n263 VTAIL.n210 3.49141
R899 VTAIL.n286 VTAIL.n198 3.49141
R900 VTAIL.n678 VTAIL.n590 3.49141
R901 VTAIL.n657 VTAIL.n604 3.49141
R902 VTAIL.n634 VTAIL.n633 3.49141
R903 VTAIL.n580 VTAIL.n492 3.49141
R904 VTAIL.n559 VTAIL.n506 3.49141
R905 VTAIL.n536 VTAIL.n535 3.49141
R906 VTAIL.n482 VTAIL.n394 3.49141
R907 VTAIL.n461 VTAIL.n408 3.49141
R908 VTAIL.n438 VTAIL.n437 3.49141
R909 VTAIL.n384 VTAIL.n296 3.49141
R910 VTAIL.n363 VTAIL.n310 3.49141
R911 VTAIL.n340 VTAIL.n339 3.49141
R912 VTAIL.n489 VTAIL.n391 3.0005
R913 VTAIL.n685 VTAIL.n587 3.0005
R914 VTAIL.n293 VTAIL.n195 3.0005
R915 VTAIL.n726 VTAIL.n712 2.71565
R916 VTAIL.n754 VTAIL.n698 2.71565
R917 VTAIL.n775 VTAIL.n690 2.71565
R918 VTAIL.n40 VTAIL.n26 2.71565
R919 VTAIL.n68 VTAIL.n12 2.71565
R920 VTAIL.n89 VTAIL.n4 2.71565
R921 VTAIL.n138 VTAIL.n124 2.71565
R922 VTAIL.n166 VTAIL.n110 2.71565
R923 VTAIL.n187 VTAIL.n102 2.71565
R924 VTAIL.n236 VTAIL.n222 2.71565
R925 VTAIL.n264 VTAIL.n208 2.71565
R926 VTAIL.n285 VTAIL.n200 2.71565
R927 VTAIL.n677 VTAIL.n592 2.71565
R928 VTAIL.n658 VTAIL.n602 2.71565
R929 VTAIL.n630 VTAIL.n616 2.71565
R930 VTAIL.n579 VTAIL.n494 2.71565
R931 VTAIL.n560 VTAIL.n504 2.71565
R932 VTAIL.n532 VTAIL.n518 2.71565
R933 VTAIL.n481 VTAIL.n396 2.71565
R934 VTAIL.n462 VTAIL.n406 2.71565
R935 VTAIL.n434 VTAIL.n420 2.71565
R936 VTAIL.n383 VTAIL.n298 2.71565
R937 VTAIL.n364 VTAIL.n308 2.71565
R938 VTAIL.n336 VTAIL.n322 2.71565
R939 VTAIL.n725 VTAIL.n714 1.93989
R940 VTAIL.n759 VTAIL.n757 1.93989
R941 VTAIL.n772 VTAIL.n771 1.93989
R942 VTAIL.n39 VTAIL.n28 1.93989
R943 VTAIL.n73 VTAIL.n71 1.93989
R944 VTAIL.n86 VTAIL.n85 1.93989
R945 VTAIL.n137 VTAIL.n126 1.93989
R946 VTAIL.n171 VTAIL.n169 1.93989
R947 VTAIL.n184 VTAIL.n183 1.93989
R948 VTAIL.n235 VTAIL.n224 1.93989
R949 VTAIL.n269 VTAIL.n267 1.93989
R950 VTAIL.n282 VTAIL.n281 1.93989
R951 VTAIL.n674 VTAIL.n673 1.93989
R952 VTAIL.n662 VTAIL.n661 1.93989
R953 VTAIL.n629 VTAIL.n618 1.93989
R954 VTAIL.n576 VTAIL.n575 1.93989
R955 VTAIL.n564 VTAIL.n563 1.93989
R956 VTAIL.n531 VTAIL.n520 1.93989
R957 VTAIL.n478 VTAIL.n477 1.93989
R958 VTAIL.n466 VTAIL.n465 1.93989
R959 VTAIL.n433 VTAIL.n422 1.93989
R960 VTAIL.n380 VTAIL.n379 1.93989
R961 VTAIL.n368 VTAIL.n367 1.93989
R962 VTAIL.n335 VTAIL.n324 1.93989
R963 VTAIL VTAIL.n97 1.55869
R964 VTAIL VTAIL.n783 1.44231
R965 VTAIL.n722 VTAIL.n721 1.16414
R966 VTAIL.n758 VTAIL.n696 1.16414
R967 VTAIL.n768 VTAIL.n692 1.16414
R968 VTAIL.n36 VTAIL.n35 1.16414
R969 VTAIL.n72 VTAIL.n10 1.16414
R970 VTAIL.n82 VTAIL.n6 1.16414
R971 VTAIL.n134 VTAIL.n133 1.16414
R972 VTAIL.n170 VTAIL.n108 1.16414
R973 VTAIL.n180 VTAIL.n104 1.16414
R974 VTAIL.n232 VTAIL.n231 1.16414
R975 VTAIL.n268 VTAIL.n206 1.16414
R976 VTAIL.n278 VTAIL.n202 1.16414
R977 VTAIL.n670 VTAIL.n594 1.16414
R978 VTAIL.n665 VTAIL.n599 1.16414
R979 VTAIL.n626 VTAIL.n625 1.16414
R980 VTAIL.n572 VTAIL.n496 1.16414
R981 VTAIL.n567 VTAIL.n501 1.16414
R982 VTAIL.n528 VTAIL.n527 1.16414
R983 VTAIL.n474 VTAIL.n398 1.16414
R984 VTAIL.n469 VTAIL.n403 1.16414
R985 VTAIL.n430 VTAIL.n429 1.16414
R986 VTAIL.n376 VTAIL.n300 1.16414
R987 VTAIL.n371 VTAIL.n305 1.16414
R988 VTAIL.n332 VTAIL.n331 1.16414
R989 VTAIL.n587 VTAIL.n489 0.470328
R990 VTAIL.n195 VTAIL.n97 0.470328
R991 VTAIL.n718 VTAIL.n716 0.388379
R992 VTAIL.n764 VTAIL.n763 0.388379
R993 VTAIL.n767 VTAIL.n694 0.388379
R994 VTAIL.n32 VTAIL.n30 0.388379
R995 VTAIL.n78 VTAIL.n77 0.388379
R996 VTAIL.n81 VTAIL.n8 0.388379
R997 VTAIL.n130 VTAIL.n128 0.388379
R998 VTAIL.n176 VTAIL.n175 0.388379
R999 VTAIL.n179 VTAIL.n106 0.388379
R1000 VTAIL.n228 VTAIL.n226 0.388379
R1001 VTAIL.n274 VTAIL.n273 0.388379
R1002 VTAIL.n277 VTAIL.n204 0.388379
R1003 VTAIL.n669 VTAIL.n596 0.388379
R1004 VTAIL.n666 VTAIL.n598 0.388379
R1005 VTAIL.n622 VTAIL.n620 0.388379
R1006 VTAIL.n571 VTAIL.n498 0.388379
R1007 VTAIL.n568 VTAIL.n500 0.388379
R1008 VTAIL.n524 VTAIL.n522 0.388379
R1009 VTAIL.n473 VTAIL.n400 0.388379
R1010 VTAIL.n470 VTAIL.n402 0.388379
R1011 VTAIL.n426 VTAIL.n424 0.388379
R1012 VTAIL.n375 VTAIL.n302 0.388379
R1013 VTAIL.n372 VTAIL.n304 0.388379
R1014 VTAIL.n328 VTAIL.n326 0.388379
R1015 VTAIL.n723 VTAIL.n715 0.155672
R1016 VTAIL.n724 VTAIL.n723 0.155672
R1017 VTAIL.n724 VTAIL.n711 0.155672
R1018 VTAIL.n731 VTAIL.n711 0.155672
R1019 VTAIL.n732 VTAIL.n731 0.155672
R1020 VTAIL.n732 VTAIL.n707 0.155672
R1021 VTAIL.n739 VTAIL.n707 0.155672
R1022 VTAIL.n740 VTAIL.n739 0.155672
R1023 VTAIL.n740 VTAIL.n703 0.155672
R1024 VTAIL.n747 VTAIL.n703 0.155672
R1025 VTAIL.n748 VTAIL.n747 0.155672
R1026 VTAIL.n748 VTAIL.n699 0.155672
R1027 VTAIL.n755 VTAIL.n699 0.155672
R1028 VTAIL.n756 VTAIL.n755 0.155672
R1029 VTAIL.n756 VTAIL.n695 0.155672
R1030 VTAIL.n765 VTAIL.n695 0.155672
R1031 VTAIL.n766 VTAIL.n765 0.155672
R1032 VTAIL.n766 VTAIL.n691 0.155672
R1033 VTAIL.n773 VTAIL.n691 0.155672
R1034 VTAIL.n774 VTAIL.n773 0.155672
R1035 VTAIL.n774 VTAIL.n687 0.155672
R1036 VTAIL.n781 VTAIL.n687 0.155672
R1037 VTAIL.n37 VTAIL.n29 0.155672
R1038 VTAIL.n38 VTAIL.n37 0.155672
R1039 VTAIL.n38 VTAIL.n25 0.155672
R1040 VTAIL.n45 VTAIL.n25 0.155672
R1041 VTAIL.n46 VTAIL.n45 0.155672
R1042 VTAIL.n46 VTAIL.n21 0.155672
R1043 VTAIL.n53 VTAIL.n21 0.155672
R1044 VTAIL.n54 VTAIL.n53 0.155672
R1045 VTAIL.n54 VTAIL.n17 0.155672
R1046 VTAIL.n61 VTAIL.n17 0.155672
R1047 VTAIL.n62 VTAIL.n61 0.155672
R1048 VTAIL.n62 VTAIL.n13 0.155672
R1049 VTAIL.n69 VTAIL.n13 0.155672
R1050 VTAIL.n70 VTAIL.n69 0.155672
R1051 VTAIL.n70 VTAIL.n9 0.155672
R1052 VTAIL.n79 VTAIL.n9 0.155672
R1053 VTAIL.n80 VTAIL.n79 0.155672
R1054 VTAIL.n80 VTAIL.n5 0.155672
R1055 VTAIL.n87 VTAIL.n5 0.155672
R1056 VTAIL.n88 VTAIL.n87 0.155672
R1057 VTAIL.n88 VTAIL.n1 0.155672
R1058 VTAIL.n95 VTAIL.n1 0.155672
R1059 VTAIL.n135 VTAIL.n127 0.155672
R1060 VTAIL.n136 VTAIL.n135 0.155672
R1061 VTAIL.n136 VTAIL.n123 0.155672
R1062 VTAIL.n143 VTAIL.n123 0.155672
R1063 VTAIL.n144 VTAIL.n143 0.155672
R1064 VTAIL.n144 VTAIL.n119 0.155672
R1065 VTAIL.n151 VTAIL.n119 0.155672
R1066 VTAIL.n152 VTAIL.n151 0.155672
R1067 VTAIL.n152 VTAIL.n115 0.155672
R1068 VTAIL.n159 VTAIL.n115 0.155672
R1069 VTAIL.n160 VTAIL.n159 0.155672
R1070 VTAIL.n160 VTAIL.n111 0.155672
R1071 VTAIL.n167 VTAIL.n111 0.155672
R1072 VTAIL.n168 VTAIL.n167 0.155672
R1073 VTAIL.n168 VTAIL.n107 0.155672
R1074 VTAIL.n177 VTAIL.n107 0.155672
R1075 VTAIL.n178 VTAIL.n177 0.155672
R1076 VTAIL.n178 VTAIL.n103 0.155672
R1077 VTAIL.n185 VTAIL.n103 0.155672
R1078 VTAIL.n186 VTAIL.n185 0.155672
R1079 VTAIL.n186 VTAIL.n99 0.155672
R1080 VTAIL.n193 VTAIL.n99 0.155672
R1081 VTAIL.n233 VTAIL.n225 0.155672
R1082 VTAIL.n234 VTAIL.n233 0.155672
R1083 VTAIL.n234 VTAIL.n221 0.155672
R1084 VTAIL.n241 VTAIL.n221 0.155672
R1085 VTAIL.n242 VTAIL.n241 0.155672
R1086 VTAIL.n242 VTAIL.n217 0.155672
R1087 VTAIL.n249 VTAIL.n217 0.155672
R1088 VTAIL.n250 VTAIL.n249 0.155672
R1089 VTAIL.n250 VTAIL.n213 0.155672
R1090 VTAIL.n257 VTAIL.n213 0.155672
R1091 VTAIL.n258 VTAIL.n257 0.155672
R1092 VTAIL.n258 VTAIL.n209 0.155672
R1093 VTAIL.n265 VTAIL.n209 0.155672
R1094 VTAIL.n266 VTAIL.n265 0.155672
R1095 VTAIL.n266 VTAIL.n205 0.155672
R1096 VTAIL.n275 VTAIL.n205 0.155672
R1097 VTAIL.n276 VTAIL.n275 0.155672
R1098 VTAIL.n276 VTAIL.n201 0.155672
R1099 VTAIL.n283 VTAIL.n201 0.155672
R1100 VTAIL.n284 VTAIL.n283 0.155672
R1101 VTAIL.n284 VTAIL.n197 0.155672
R1102 VTAIL.n291 VTAIL.n197 0.155672
R1103 VTAIL.n683 VTAIL.n589 0.155672
R1104 VTAIL.n676 VTAIL.n589 0.155672
R1105 VTAIL.n676 VTAIL.n675 0.155672
R1106 VTAIL.n675 VTAIL.n593 0.155672
R1107 VTAIL.n668 VTAIL.n593 0.155672
R1108 VTAIL.n668 VTAIL.n667 0.155672
R1109 VTAIL.n667 VTAIL.n597 0.155672
R1110 VTAIL.n660 VTAIL.n597 0.155672
R1111 VTAIL.n660 VTAIL.n659 0.155672
R1112 VTAIL.n659 VTAIL.n603 0.155672
R1113 VTAIL.n652 VTAIL.n603 0.155672
R1114 VTAIL.n652 VTAIL.n651 0.155672
R1115 VTAIL.n651 VTAIL.n607 0.155672
R1116 VTAIL.n644 VTAIL.n607 0.155672
R1117 VTAIL.n644 VTAIL.n643 0.155672
R1118 VTAIL.n643 VTAIL.n611 0.155672
R1119 VTAIL.n636 VTAIL.n611 0.155672
R1120 VTAIL.n636 VTAIL.n635 0.155672
R1121 VTAIL.n635 VTAIL.n615 0.155672
R1122 VTAIL.n628 VTAIL.n615 0.155672
R1123 VTAIL.n628 VTAIL.n627 0.155672
R1124 VTAIL.n627 VTAIL.n619 0.155672
R1125 VTAIL.n585 VTAIL.n491 0.155672
R1126 VTAIL.n578 VTAIL.n491 0.155672
R1127 VTAIL.n578 VTAIL.n577 0.155672
R1128 VTAIL.n577 VTAIL.n495 0.155672
R1129 VTAIL.n570 VTAIL.n495 0.155672
R1130 VTAIL.n570 VTAIL.n569 0.155672
R1131 VTAIL.n569 VTAIL.n499 0.155672
R1132 VTAIL.n562 VTAIL.n499 0.155672
R1133 VTAIL.n562 VTAIL.n561 0.155672
R1134 VTAIL.n561 VTAIL.n505 0.155672
R1135 VTAIL.n554 VTAIL.n505 0.155672
R1136 VTAIL.n554 VTAIL.n553 0.155672
R1137 VTAIL.n553 VTAIL.n509 0.155672
R1138 VTAIL.n546 VTAIL.n509 0.155672
R1139 VTAIL.n546 VTAIL.n545 0.155672
R1140 VTAIL.n545 VTAIL.n513 0.155672
R1141 VTAIL.n538 VTAIL.n513 0.155672
R1142 VTAIL.n538 VTAIL.n537 0.155672
R1143 VTAIL.n537 VTAIL.n517 0.155672
R1144 VTAIL.n530 VTAIL.n517 0.155672
R1145 VTAIL.n530 VTAIL.n529 0.155672
R1146 VTAIL.n529 VTAIL.n521 0.155672
R1147 VTAIL.n487 VTAIL.n393 0.155672
R1148 VTAIL.n480 VTAIL.n393 0.155672
R1149 VTAIL.n480 VTAIL.n479 0.155672
R1150 VTAIL.n479 VTAIL.n397 0.155672
R1151 VTAIL.n472 VTAIL.n397 0.155672
R1152 VTAIL.n472 VTAIL.n471 0.155672
R1153 VTAIL.n471 VTAIL.n401 0.155672
R1154 VTAIL.n464 VTAIL.n401 0.155672
R1155 VTAIL.n464 VTAIL.n463 0.155672
R1156 VTAIL.n463 VTAIL.n407 0.155672
R1157 VTAIL.n456 VTAIL.n407 0.155672
R1158 VTAIL.n456 VTAIL.n455 0.155672
R1159 VTAIL.n455 VTAIL.n411 0.155672
R1160 VTAIL.n448 VTAIL.n411 0.155672
R1161 VTAIL.n448 VTAIL.n447 0.155672
R1162 VTAIL.n447 VTAIL.n415 0.155672
R1163 VTAIL.n440 VTAIL.n415 0.155672
R1164 VTAIL.n440 VTAIL.n439 0.155672
R1165 VTAIL.n439 VTAIL.n419 0.155672
R1166 VTAIL.n432 VTAIL.n419 0.155672
R1167 VTAIL.n432 VTAIL.n431 0.155672
R1168 VTAIL.n431 VTAIL.n423 0.155672
R1169 VTAIL.n389 VTAIL.n295 0.155672
R1170 VTAIL.n382 VTAIL.n295 0.155672
R1171 VTAIL.n382 VTAIL.n381 0.155672
R1172 VTAIL.n381 VTAIL.n299 0.155672
R1173 VTAIL.n374 VTAIL.n299 0.155672
R1174 VTAIL.n374 VTAIL.n373 0.155672
R1175 VTAIL.n373 VTAIL.n303 0.155672
R1176 VTAIL.n366 VTAIL.n303 0.155672
R1177 VTAIL.n366 VTAIL.n365 0.155672
R1178 VTAIL.n365 VTAIL.n309 0.155672
R1179 VTAIL.n358 VTAIL.n309 0.155672
R1180 VTAIL.n358 VTAIL.n357 0.155672
R1181 VTAIL.n357 VTAIL.n313 0.155672
R1182 VTAIL.n350 VTAIL.n313 0.155672
R1183 VTAIL.n350 VTAIL.n349 0.155672
R1184 VTAIL.n349 VTAIL.n317 0.155672
R1185 VTAIL.n342 VTAIL.n317 0.155672
R1186 VTAIL.n342 VTAIL.n341 0.155672
R1187 VTAIL.n341 VTAIL.n321 0.155672
R1188 VTAIL.n334 VTAIL.n321 0.155672
R1189 VTAIL.n334 VTAIL.n333 0.155672
R1190 VTAIL.n333 VTAIL.n325 0.155672
R1191 VDD2.n2 VDD2.n0 117.853
R1192 VDD2.n2 VDD2.n1 69.9917
R1193 VDD2.n1 VDD2.t0 1.85053
R1194 VDD2.n1 VDD2.t2 1.85053
R1195 VDD2.n0 VDD2.t1 1.85053
R1196 VDD2.n0 VDD2.t3 1.85053
R1197 VDD2 VDD2.n2 0.0586897
R1198 VP.n5 VP.t2 168.899
R1199 VP.n5 VP.t3 167.815
R1200 VP.n17 VP.n16 161.3
R1201 VP.n15 VP.n1 161.3
R1202 VP.n14 VP.n13 161.3
R1203 VP.n12 VP.n2 161.3
R1204 VP.n11 VP.n10 161.3
R1205 VP.n9 VP.n3 161.3
R1206 VP.n8 VP.n7 161.3
R1207 VP.n4 VP.t0 134.424
R1208 VP.n0 VP.t1 134.424
R1209 VP.n6 VP.n4 78.3232
R1210 VP.n18 VP.n0 78.3232
R1211 VP.n6 VP.n5 54.8705
R1212 VP.n10 VP.n2 40.4934
R1213 VP.n14 VP.n2 40.4934
R1214 VP.n9 VP.n8 24.4675
R1215 VP.n10 VP.n9 24.4675
R1216 VP.n15 VP.n14 24.4675
R1217 VP.n16 VP.n15 24.4675
R1218 VP.n8 VP.n4 11.7447
R1219 VP.n16 VP.n0 11.7447
R1220 VP.n7 VP.n6 0.354971
R1221 VP.n18 VP.n17 0.354971
R1222 VP VP.n18 0.26696
R1223 VP.n7 VP.n3 0.189894
R1224 VP.n11 VP.n3 0.189894
R1225 VP.n12 VP.n11 0.189894
R1226 VP.n13 VP.n12 0.189894
R1227 VP.n13 VP.n1 0.189894
R1228 VP.n17 VP.n1 0.189894
R1229 VDD1 VDD1.n1 118.377
R1230 VDD1 VDD1.n0 70.0499
R1231 VDD1.n0 VDD1.t1 1.85053
R1232 VDD1.n0 VDD1.t0 1.85053
R1233 VDD1.n1 VDD1.t3 1.85053
R1234 VDD1.n1 VDD1.t2 1.85053
R1235 B.n582 B.n89 585
R1236 B.n584 B.n583 585
R1237 B.n585 B.n88 585
R1238 B.n587 B.n586 585
R1239 B.n588 B.n87 585
R1240 B.n590 B.n589 585
R1241 B.n591 B.n86 585
R1242 B.n593 B.n592 585
R1243 B.n594 B.n85 585
R1244 B.n596 B.n595 585
R1245 B.n597 B.n84 585
R1246 B.n599 B.n598 585
R1247 B.n600 B.n83 585
R1248 B.n602 B.n601 585
R1249 B.n603 B.n82 585
R1250 B.n605 B.n604 585
R1251 B.n606 B.n81 585
R1252 B.n608 B.n607 585
R1253 B.n609 B.n80 585
R1254 B.n611 B.n610 585
R1255 B.n612 B.n79 585
R1256 B.n614 B.n613 585
R1257 B.n615 B.n78 585
R1258 B.n617 B.n616 585
R1259 B.n618 B.n77 585
R1260 B.n620 B.n619 585
R1261 B.n621 B.n76 585
R1262 B.n623 B.n622 585
R1263 B.n624 B.n75 585
R1264 B.n626 B.n625 585
R1265 B.n627 B.n74 585
R1266 B.n629 B.n628 585
R1267 B.n630 B.n73 585
R1268 B.n632 B.n631 585
R1269 B.n633 B.n72 585
R1270 B.n635 B.n634 585
R1271 B.n636 B.n71 585
R1272 B.n638 B.n637 585
R1273 B.n639 B.n70 585
R1274 B.n641 B.n640 585
R1275 B.n642 B.n69 585
R1276 B.n644 B.n643 585
R1277 B.n645 B.n68 585
R1278 B.n647 B.n646 585
R1279 B.n648 B.n67 585
R1280 B.n650 B.n649 585
R1281 B.n651 B.n66 585
R1282 B.n653 B.n652 585
R1283 B.n654 B.n65 585
R1284 B.n656 B.n655 585
R1285 B.n657 B.n64 585
R1286 B.n659 B.n658 585
R1287 B.n660 B.n63 585
R1288 B.n662 B.n661 585
R1289 B.n663 B.n62 585
R1290 B.n665 B.n664 585
R1291 B.n666 B.n61 585
R1292 B.n668 B.n667 585
R1293 B.n670 B.n58 585
R1294 B.n672 B.n671 585
R1295 B.n673 B.n57 585
R1296 B.n675 B.n674 585
R1297 B.n676 B.n56 585
R1298 B.n678 B.n677 585
R1299 B.n679 B.n55 585
R1300 B.n681 B.n680 585
R1301 B.n682 B.n51 585
R1302 B.n684 B.n683 585
R1303 B.n685 B.n50 585
R1304 B.n687 B.n686 585
R1305 B.n688 B.n49 585
R1306 B.n690 B.n689 585
R1307 B.n691 B.n48 585
R1308 B.n693 B.n692 585
R1309 B.n694 B.n47 585
R1310 B.n696 B.n695 585
R1311 B.n697 B.n46 585
R1312 B.n699 B.n698 585
R1313 B.n700 B.n45 585
R1314 B.n702 B.n701 585
R1315 B.n703 B.n44 585
R1316 B.n705 B.n704 585
R1317 B.n706 B.n43 585
R1318 B.n708 B.n707 585
R1319 B.n709 B.n42 585
R1320 B.n711 B.n710 585
R1321 B.n712 B.n41 585
R1322 B.n714 B.n713 585
R1323 B.n715 B.n40 585
R1324 B.n717 B.n716 585
R1325 B.n718 B.n39 585
R1326 B.n720 B.n719 585
R1327 B.n721 B.n38 585
R1328 B.n723 B.n722 585
R1329 B.n724 B.n37 585
R1330 B.n726 B.n725 585
R1331 B.n727 B.n36 585
R1332 B.n729 B.n728 585
R1333 B.n730 B.n35 585
R1334 B.n732 B.n731 585
R1335 B.n733 B.n34 585
R1336 B.n735 B.n734 585
R1337 B.n736 B.n33 585
R1338 B.n738 B.n737 585
R1339 B.n739 B.n32 585
R1340 B.n741 B.n740 585
R1341 B.n742 B.n31 585
R1342 B.n744 B.n743 585
R1343 B.n745 B.n30 585
R1344 B.n747 B.n746 585
R1345 B.n748 B.n29 585
R1346 B.n750 B.n749 585
R1347 B.n751 B.n28 585
R1348 B.n753 B.n752 585
R1349 B.n754 B.n27 585
R1350 B.n756 B.n755 585
R1351 B.n757 B.n26 585
R1352 B.n759 B.n758 585
R1353 B.n760 B.n25 585
R1354 B.n762 B.n761 585
R1355 B.n763 B.n24 585
R1356 B.n765 B.n764 585
R1357 B.n766 B.n23 585
R1358 B.n768 B.n767 585
R1359 B.n769 B.n22 585
R1360 B.n771 B.n770 585
R1361 B.n581 B.n580 585
R1362 B.n579 B.n90 585
R1363 B.n578 B.n577 585
R1364 B.n576 B.n91 585
R1365 B.n575 B.n574 585
R1366 B.n573 B.n92 585
R1367 B.n572 B.n571 585
R1368 B.n570 B.n93 585
R1369 B.n569 B.n568 585
R1370 B.n567 B.n94 585
R1371 B.n566 B.n565 585
R1372 B.n564 B.n95 585
R1373 B.n563 B.n562 585
R1374 B.n561 B.n96 585
R1375 B.n560 B.n559 585
R1376 B.n558 B.n97 585
R1377 B.n557 B.n556 585
R1378 B.n555 B.n98 585
R1379 B.n554 B.n553 585
R1380 B.n552 B.n99 585
R1381 B.n551 B.n550 585
R1382 B.n549 B.n100 585
R1383 B.n548 B.n547 585
R1384 B.n546 B.n101 585
R1385 B.n545 B.n544 585
R1386 B.n543 B.n102 585
R1387 B.n542 B.n541 585
R1388 B.n540 B.n103 585
R1389 B.n539 B.n538 585
R1390 B.n537 B.n104 585
R1391 B.n536 B.n535 585
R1392 B.n534 B.n105 585
R1393 B.n533 B.n532 585
R1394 B.n531 B.n106 585
R1395 B.n530 B.n529 585
R1396 B.n528 B.n107 585
R1397 B.n527 B.n526 585
R1398 B.n525 B.n108 585
R1399 B.n524 B.n523 585
R1400 B.n522 B.n109 585
R1401 B.n521 B.n520 585
R1402 B.n519 B.n110 585
R1403 B.n518 B.n517 585
R1404 B.n516 B.n111 585
R1405 B.n515 B.n514 585
R1406 B.n513 B.n112 585
R1407 B.n512 B.n511 585
R1408 B.n510 B.n113 585
R1409 B.n509 B.n508 585
R1410 B.n507 B.n114 585
R1411 B.n506 B.n505 585
R1412 B.n504 B.n115 585
R1413 B.n503 B.n502 585
R1414 B.n501 B.n116 585
R1415 B.n500 B.n499 585
R1416 B.n498 B.n117 585
R1417 B.n497 B.n496 585
R1418 B.n495 B.n118 585
R1419 B.n494 B.n493 585
R1420 B.n492 B.n119 585
R1421 B.n491 B.n490 585
R1422 B.n489 B.n120 585
R1423 B.n488 B.n487 585
R1424 B.n486 B.n121 585
R1425 B.n485 B.n484 585
R1426 B.n483 B.n122 585
R1427 B.n482 B.n481 585
R1428 B.n480 B.n123 585
R1429 B.n479 B.n478 585
R1430 B.n477 B.n124 585
R1431 B.n476 B.n475 585
R1432 B.n474 B.n125 585
R1433 B.n473 B.n472 585
R1434 B.n471 B.n126 585
R1435 B.n470 B.n469 585
R1436 B.n468 B.n127 585
R1437 B.n467 B.n466 585
R1438 B.n465 B.n128 585
R1439 B.n464 B.n463 585
R1440 B.n273 B.n196 585
R1441 B.n275 B.n274 585
R1442 B.n276 B.n195 585
R1443 B.n278 B.n277 585
R1444 B.n279 B.n194 585
R1445 B.n281 B.n280 585
R1446 B.n282 B.n193 585
R1447 B.n284 B.n283 585
R1448 B.n285 B.n192 585
R1449 B.n287 B.n286 585
R1450 B.n288 B.n191 585
R1451 B.n290 B.n289 585
R1452 B.n291 B.n190 585
R1453 B.n293 B.n292 585
R1454 B.n294 B.n189 585
R1455 B.n296 B.n295 585
R1456 B.n297 B.n188 585
R1457 B.n299 B.n298 585
R1458 B.n300 B.n187 585
R1459 B.n302 B.n301 585
R1460 B.n303 B.n186 585
R1461 B.n305 B.n304 585
R1462 B.n306 B.n185 585
R1463 B.n308 B.n307 585
R1464 B.n309 B.n184 585
R1465 B.n311 B.n310 585
R1466 B.n312 B.n183 585
R1467 B.n314 B.n313 585
R1468 B.n315 B.n182 585
R1469 B.n317 B.n316 585
R1470 B.n318 B.n181 585
R1471 B.n320 B.n319 585
R1472 B.n321 B.n180 585
R1473 B.n323 B.n322 585
R1474 B.n324 B.n179 585
R1475 B.n326 B.n325 585
R1476 B.n327 B.n178 585
R1477 B.n329 B.n328 585
R1478 B.n330 B.n177 585
R1479 B.n332 B.n331 585
R1480 B.n333 B.n176 585
R1481 B.n335 B.n334 585
R1482 B.n336 B.n175 585
R1483 B.n338 B.n337 585
R1484 B.n339 B.n174 585
R1485 B.n341 B.n340 585
R1486 B.n342 B.n173 585
R1487 B.n344 B.n343 585
R1488 B.n345 B.n172 585
R1489 B.n347 B.n346 585
R1490 B.n348 B.n171 585
R1491 B.n350 B.n349 585
R1492 B.n351 B.n170 585
R1493 B.n353 B.n352 585
R1494 B.n354 B.n169 585
R1495 B.n356 B.n355 585
R1496 B.n357 B.n168 585
R1497 B.n359 B.n358 585
R1498 B.n361 B.n360 585
R1499 B.n362 B.n164 585
R1500 B.n364 B.n363 585
R1501 B.n365 B.n163 585
R1502 B.n367 B.n366 585
R1503 B.n368 B.n162 585
R1504 B.n370 B.n369 585
R1505 B.n371 B.n161 585
R1506 B.n373 B.n372 585
R1507 B.n374 B.n158 585
R1508 B.n377 B.n376 585
R1509 B.n378 B.n157 585
R1510 B.n380 B.n379 585
R1511 B.n381 B.n156 585
R1512 B.n383 B.n382 585
R1513 B.n384 B.n155 585
R1514 B.n386 B.n385 585
R1515 B.n387 B.n154 585
R1516 B.n389 B.n388 585
R1517 B.n390 B.n153 585
R1518 B.n392 B.n391 585
R1519 B.n393 B.n152 585
R1520 B.n395 B.n394 585
R1521 B.n396 B.n151 585
R1522 B.n398 B.n397 585
R1523 B.n399 B.n150 585
R1524 B.n401 B.n400 585
R1525 B.n402 B.n149 585
R1526 B.n404 B.n403 585
R1527 B.n405 B.n148 585
R1528 B.n407 B.n406 585
R1529 B.n408 B.n147 585
R1530 B.n410 B.n409 585
R1531 B.n411 B.n146 585
R1532 B.n413 B.n412 585
R1533 B.n414 B.n145 585
R1534 B.n416 B.n415 585
R1535 B.n417 B.n144 585
R1536 B.n419 B.n418 585
R1537 B.n420 B.n143 585
R1538 B.n422 B.n421 585
R1539 B.n423 B.n142 585
R1540 B.n425 B.n424 585
R1541 B.n426 B.n141 585
R1542 B.n428 B.n427 585
R1543 B.n429 B.n140 585
R1544 B.n431 B.n430 585
R1545 B.n432 B.n139 585
R1546 B.n434 B.n433 585
R1547 B.n435 B.n138 585
R1548 B.n437 B.n436 585
R1549 B.n438 B.n137 585
R1550 B.n440 B.n439 585
R1551 B.n441 B.n136 585
R1552 B.n443 B.n442 585
R1553 B.n444 B.n135 585
R1554 B.n446 B.n445 585
R1555 B.n447 B.n134 585
R1556 B.n449 B.n448 585
R1557 B.n450 B.n133 585
R1558 B.n452 B.n451 585
R1559 B.n453 B.n132 585
R1560 B.n455 B.n454 585
R1561 B.n456 B.n131 585
R1562 B.n458 B.n457 585
R1563 B.n459 B.n130 585
R1564 B.n461 B.n460 585
R1565 B.n462 B.n129 585
R1566 B.n272 B.n271 585
R1567 B.n270 B.n197 585
R1568 B.n269 B.n268 585
R1569 B.n267 B.n198 585
R1570 B.n266 B.n265 585
R1571 B.n264 B.n199 585
R1572 B.n263 B.n262 585
R1573 B.n261 B.n200 585
R1574 B.n260 B.n259 585
R1575 B.n258 B.n201 585
R1576 B.n257 B.n256 585
R1577 B.n255 B.n202 585
R1578 B.n254 B.n253 585
R1579 B.n252 B.n203 585
R1580 B.n251 B.n250 585
R1581 B.n249 B.n204 585
R1582 B.n248 B.n247 585
R1583 B.n246 B.n205 585
R1584 B.n245 B.n244 585
R1585 B.n243 B.n206 585
R1586 B.n242 B.n241 585
R1587 B.n240 B.n207 585
R1588 B.n239 B.n238 585
R1589 B.n237 B.n208 585
R1590 B.n236 B.n235 585
R1591 B.n234 B.n209 585
R1592 B.n233 B.n232 585
R1593 B.n231 B.n210 585
R1594 B.n230 B.n229 585
R1595 B.n228 B.n211 585
R1596 B.n227 B.n226 585
R1597 B.n225 B.n212 585
R1598 B.n224 B.n223 585
R1599 B.n222 B.n213 585
R1600 B.n221 B.n220 585
R1601 B.n219 B.n214 585
R1602 B.n218 B.n217 585
R1603 B.n216 B.n215 585
R1604 B.n2 B.n0 585
R1605 B.n829 B.n1 585
R1606 B.n828 B.n827 585
R1607 B.n826 B.n3 585
R1608 B.n825 B.n824 585
R1609 B.n823 B.n4 585
R1610 B.n822 B.n821 585
R1611 B.n820 B.n5 585
R1612 B.n819 B.n818 585
R1613 B.n817 B.n6 585
R1614 B.n816 B.n815 585
R1615 B.n814 B.n7 585
R1616 B.n813 B.n812 585
R1617 B.n811 B.n8 585
R1618 B.n810 B.n809 585
R1619 B.n808 B.n9 585
R1620 B.n807 B.n806 585
R1621 B.n805 B.n10 585
R1622 B.n804 B.n803 585
R1623 B.n802 B.n11 585
R1624 B.n801 B.n800 585
R1625 B.n799 B.n12 585
R1626 B.n798 B.n797 585
R1627 B.n796 B.n13 585
R1628 B.n795 B.n794 585
R1629 B.n793 B.n14 585
R1630 B.n792 B.n791 585
R1631 B.n790 B.n15 585
R1632 B.n789 B.n788 585
R1633 B.n787 B.n16 585
R1634 B.n786 B.n785 585
R1635 B.n784 B.n17 585
R1636 B.n783 B.n782 585
R1637 B.n781 B.n18 585
R1638 B.n780 B.n779 585
R1639 B.n778 B.n19 585
R1640 B.n777 B.n776 585
R1641 B.n775 B.n20 585
R1642 B.n774 B.n773 585
R1643 B.n772 B.n21 585
R1644 B.n831 B.n830 585
R1645 B.n159 B.t5 543.525
R1646 B.n59 B.t1 543.525
R1647 B.n165 B.t8 543.525
R1648 B.n52 B.t10 543.525
R1649 B.n160 B.t4 476.034
R1650 B.n60 B.t2 476.034
R1651 B.n166 B.t7 476.034
R1652 B.n53 B.t11 476.034
R1653 B.n271 B.n196 434.841
R1654 B.n770 B.n21 434.841
R1655 B.n463 B.n462 434.841
R1656 B.n582 B.n581 434.841
R1657 B.n159 B.t3 343.173
R1658 B.n165 B.t6 343.173
R1659 B.n52 B.t9 343.173
R1660 B.n59 B.t0 343.173
R1661 B.n271 B.n270 163.367
R1662 B.n270 B.n269 163.367
R1663 B.n269 B.n198 163.367
R1664 B.n265 B.n198 163.367
R1665 B.n265 B.n264 163.367
R1666 B.n264 B.n263 163.367
R1667 B.n263 B.n200 163.367
R1668 B.n259 B.n200 163.367
R1669 B.n259 B.n258 163.367
R1670 B.n258 B.n257 163.367
R1671 B.n257 B.n202 163.367
R1672 B.n253 B.n202 163.367
R1673 B.n253 B.n252 163.367
R1674 B.n252 B.n251 163.367
R1675 B.n251 B.n204 163.367
R1676 B.n247 B.n204 163.367
R1677 B.n247 B.n246 163.367
R1678 B.n246 B.n245 163.367
R1679 B.n245 B.n206 163.367
R1680 B.n241 B.n206 163.367
R1681 B.n241 B.n240 163.367
R1682 B.n240 B.n239 163.367
R1683 B.n239 B.n208 163.367
R1684 B.n235 B.n208 163.367
R1685 B.n235 B.n234 163.367
R1686 B.n234 B.n233 163.367
R1687 B.n233 B.n210 163.367
R1688 B.n229 B.n210 163.367
R1689 B.n229 B.n228 163.367
R1690 B.n228 B.n227 163.367
R1691 B.n227 B.n212 163.367
R1692 B.n223 B.n212 163.367
R1693 B.n223 B.n222 163.367
R1694 B.n222 B.n221 163.367
R1695 B.n221 B.n214 163.367
R1696 B.n217 B.n214 163.367
R1697 B.n217 B.n216 163.367
R1698 B.n216 B.n2 163.367
R1699 B.n830 B.n2 163.367
R1700 B.n830 B.n829 163.367
R1701 B.n829 B.n828 163.367
R1702 B.n828 B.n3 163.367
R1703 B.n824 B.n3 163.367
R1704 B.n824 B.n823 163.367
R1705 B.n823 B.n822 163.367
R1706 B.n822 B.n5 163.367
R1707 B.n818 B.n5 163.367
R1708 B.n818 B.n817 163.367
R1709 B.n817 B.n816 163.367
R1710 B.n816 B.n7 163.367
R1711 B.n812 B.n7 163.367
R1712 B.n812 B.n811 163.367
R1713 B.n811 B.n810 163.367
R1714 B.n810 B.n9 163.367
R1715 B.n806 B.n9 163.367
R1716 B.n806 B.n805 163.367
R1717 B.n805 B.n804 163.367
R1718 B.n804 B.n11 163.367
R1719 B.n800 B.n11 163.367
R1720 B.n800 B.n799 163.367
R1721 B.n799 B.n798 163.367
R1722 B.n798 B.n13 163.367
R1723 B.n794 B.n13 163.367
R1724 B.n794 B.n793 163.367
R1725 B.n793 B.n792 163.367
R1726 B.n792 B.n15 163.367
R1727 B.n788 B.n15 163.367
R1728 B.n788 B.n787 163.367
R1729 B.n787 B.n786 163.367
R1730 B.n786 B.n17 163.367
R1731 B.n782 B.n17 163.367
R1732 B.n782 B.n781 163.367
R1733 B.n781 B.n780 163.367
R1734 B.n780 B.n19 163.367
R1735 B.n776 B.n19 163.367
R1736 B.n776 B.n775 163.367
R1737 B.n775 B.n774 163.367
R1738 B.n774 B.n21 163.367
R1739 B.n275 B.n196 163.367
R1740 B.n276 B.n275 163.367
R1741 B.n277 B.n276 163.367
R1742 B.n277 B.n194 163.367
R1743 B.n281 B.n194 163.367
R1744 B.n282 B.n281 163.367
R1745 B.n283 B.n282 163.367
R1746 B.n283 B.n192 163.367
R1747 B.n287 B.n192 163.367
R1748 B.n288 B.n287 163.367
R1749 B.n289 B.n288 163.367
R1750 B.n289 B.n190 163.367
R1751 B.n293 B.n190 163.367
R1752 B.n294 B.n293 163.367
R1753 B.n295 B.n294 163.367
R1754 B.n295 B.n188 163.367
R1755 B.n299 B.n188 163.367
R1756 B.n300 B.n299 163.367
R1757 B.n301 B.n300 163.367
R1758 B.n301 B.n186 163.367
R1759 B.n305 B.n186 163.367
R1760 B.n306 B.n305 163.367
R1761 B.n307 B.n306 163.367
R1762 B.n307 B.n184 163.367
R1763 B.n311 B.n184 163.367
R1764 B.n312 B.n311 163.367
R1765 B.n313 B.n312 163.367
R1766 B.n313 B.n182 163.367
R1767 B.n317 B.n182 163.367
R1768 B.n318 B.n317 163.367
R1769 B.n319 B.n318 163.367
R1770 B.n319 B.n180 163.367
R1771 B.n323 B.n180 163.367
R1772 B.n324 B.n323 163.367
R1773 B.n325 B.n324 163.367
R1774 B.n325 B.n178 163.367
R1775 B.n329 B.n178 163.367
R1776 B.n330 B.n329 163.367
R1777 B.n331 B.n330 163.367
R1778 B.n331 B.n176 163.367
R1779 B.n335 B.n176 163.367
R1780 B.n336 B.n335 163.367
R1781 B.n337 B.n336 163.367
R1782 B.n337 B.n174 163.367
R1783 B.n341 B.n174 163.367
R1784 B.n342 B.n341 163.367
R1785 B.n343 B.n342 163.367
R1786 B.n343 B.n172 163.367
R1787 B.n347 B.n172 163.367
R1788 B.n348 B.n347 163.367
R1789 B.n349 B.n348 163.367
R1790 B.n349 B.n170 163.367
R1791 B.n353 B.n170 163.367
R1792 B.n354 B.n353 163.367
R1793 B.n355 B.n354 163.367
R1794 B.n355 B.n168 163.367
R1795 B.n359 B.n168 163.367
R1796 B.n360 B.n359 163.367
R1797 B.n360 B.n164 163.367
R1798 B.n364 B.n164 163.367
R1799 B.n365 B.n364 163.367
R1800 B.n366 B.n365 163.367
R1801 B.n366 B.n162 163.367
R1802 B.n370 B.n162 163.367
R1803 B.n371 B.n370 163.367
R1804 B.n372 B.n371 163.367
R1805 B.n372 B.n158 163.367
R1806 B.n377 B.n158 163.367
R1807 B.n378 B.n377 163.367
R1808 B.n379 B.n378 163.367
R1809 B.n379 B.n156 163.367
R1810 B.n383 B.n156 163.367
R1811 B.n384 B.n383 163.367
R1812 B.n385 B.n384 163.367
R1813 B.n385 B.n154 163.367
R1814 B.n389 B.n154 163.367
R1815 B.n390 B.n389 163.367
R1816 B.n391 B.n390 163.367
R1817 B.n391 B.n152 163.367
R1818 B.n395 B.n152 163.367
R1819 B.n396 B.n395 163.367
R1820 B.n397 B.n396 163.367
R1821 B.n397 B.n150 163.367
R1822 B.n401 B.n150 163.367
R1823 B.n402 B.n401 163.367
R1824 B.n403 B.n402 163.367
R1825 B.n403 B.n148 163.367
R1826 B.n407 B.n148 163.367
R1827 B.n408 B.n407 163.367
R1828 B.n409 B.n408 163.367
R1829 B.n409 B.n146 163.367
R1830 B.n413 B.n146 163.367
R1831 B.n414 B.n413 163.367
R1832 B.n415 B.n414 163.367
R1833 B.n415 B.n144 163.367
R1834 B.n419 B.n144 163.367
R1835 B.n420 B.n419 163.367
R1836 B.n421 B.n420 163.367
R1837 B.n421 B.n142 163.367
R1838 B.n425 B.n142 163.367
R1839 B.n426 B.n425 163.367
R1840 B.n427 B.n426 163.367
R1841 B.n427 B.n140 163.367
R1842 B.n431 B.n140 163.367
R1843 B.n432 B.n431 163.367
R1844 B.n433 B.n432 163.367
R1845 B.n433 B.n138 163.367
R1846 B.n437 B.n138 163.367
R1847 B.n438 B.n437 163.367
R1848 B.n439 B.n438 163.367
R1849 B.n439 B.n136 163.367
R1850 B.n443 B.n136 163.367
R1851 B.n444 B.n443 163.367
R1852 B.n445 B.n444 163.367
R1853 B.n445 B.n134 163.367
R1854 B.n449 B.n134 163.367
R1855 B.n450 B.n449 163.367
R1856 B.n451 B.n450 163.367
R1857 B.n451 B.n132 163.367
R1858 B.n455 B.n132 163.367
R1859 B.n456 B.n455 163.367
R1860 B.n457 B.n456 163.367
R1861 B.n457 B.n130 163.367
R1862 B.n461 B.n130 163.367
R1863 B.n462 B.n461 163.367
R1864 B.n463 B.n128 163.367
R1865 B.n467 B.n128 163.367
R1866 B.n468 B.n467 163.367
R1867 B.n469 B.n468 163.367
R1868 B.n469 B.n126 163.367
R1869 B.n473 B.n126 163.367
R1870 B.n474 B.n473 163.367
R1871 B.n475 B.n474 163.367
R1872 B.n475 B.n124 163.367
R1873 B.n479 B.n124 163.367
R1874 B.n480 B.n479 163.367
R1875 B.n481 B.n480 163.367
R1876 B.n481 B.n122 163.367
R1877 B.n485 B.n122 163.367
R1878 B.n486 B.n485 163.367
R1879 B.n487 B.n486 163.367
R1880 B.n487 B.n120 163.367
R1881 B.n491 B.n120 163.367
R1882 B.n492 B.n491 163.367
R1883 B.n493 B.n492 163.367
R1884 B.n493 B.n118 163.367
R1885 B.n497 B.n118 163.367
R1886 B.n498 B.n497 163.367
R1887 B.n499 B.n498 163.367
R1888 B.n499 B.n116 163.367
R1889 B.n503 B.n116 163.367
R1890 B.n504 B.n503 163.367
R1891 B.n505 B.n504 163.367
R1892 B.n505 B.n114 163.367
R1893 B.n509 B.n114 163.367
R1894 B.n510 B.n509 163.367
R1895 B.n511 B.n510 163.367
R1896 B.n511 B.n112 163.367
R1897 B.n515 B.n112 163.367
R1898 B.n516 B.n515 163.367
R1899 B.n517 B.n516 163.367
R1900 B.n517 B.n110 163.367
R1901 B.n521 B.n110 163.367
R1902 B.n522 B.n521 163.367
R1903 B.n523 B.n522 163.367
R1904 B.n523 B.n108 163.367
R1905 B.n527 B.n108 163.367
R1906 B.n528 B.n527 163.367
R1907 B.n529 B.n528 163.367
R1908 B.n529 B.n106 163.367
R1909 B.n533 B.n106 163.367
R1910 B.n534 B.n533 163.367
R1911 B.n535 B.n534 163.367
R1912 B.n535 B.n104 163.367
R1913 B.n539 B.n104 163.367
R1914 B.n540 B.n539 163.367
R1915 B.n541 B.n540 163.367
R1916 B.n541 B.n102 163.367
R1917 B.n545 B.n102 163.367
R1918 B.n546 B.n545 163.367
R1919 B.n547 B.n546 163.367
R1920 B.n547 B.n100 163.367
R1921 B.n551 B.n100 163.367
R1922 B.n552 B.n551 163.367
R1923 B.n553 B.n552 163.367
R1924 B.n553 B.n98 163.367
R1925 B.n557 B.n98 163.367
R1926 B.n558 B.n557 163.367
R1927 B.n559 B.n558 163.367
R1928 B.n559 B.n96 163.367
R1929 B.n563 B.n96 163.367
R1930 B.n564 B.n563 163.367
R1931 B.n565 B.n564 163.367
R1932 B.n565 B.n94 163.367
R1933 B.n569 B.n94 163.367
R1934 B.n570 B.n569 163.367
R1935 B.n571 B.n570 163.367
R1936 B.n571 B.n92 163.367
R1937 B.n575 B.n92 163.367
R1938 B.n576 B.n575 163.367
R1939 B.n577 B.n576 163.367
R1940 B.n577 B.n90 163.367
R1941 B.n581 B.n90 163.367
R1942 B.n770 B.n769 163.367
R1943 B.n769 B.n768 163.367
R1944 B.n768 B.n23 163.367
R1945 B.n764 B.n23 163.367
R1946 B.n764 B.n763 163.367
R1947 B.n763 B.n762 163.367
R1948 B.n762 B.n25 163.367
R1949 B.n758 B.n25 163.367
R1950 B.n758 B.n757 163.367
R1951 B.n757 B.n756 163.367
R1952 B.n756 B.n27 163.367
R1953 B.n752 B.n27 163.367
R1954 B.n752 B.n751 163.367
R1955 B.n751 B.n750 163.367
R1956 B.n750 B.n29 163.367
R1957 B.n746 B.n29 163.367
R1958 B.n746 B.n745 163.367
R1959 B.n745 B.n744 163.367
R1960 B.n744 B.n31 163.367
R1961 B.n740 B.n31 163.367
R1962 B.n740 B.n739 163.367
R1963 B.n739 B.n738 163.367
R1964 B.n738 B.n33 163.367
R1965 B.n734 B.n33 163.367
R1966 B.n734 B.n733 163.367
R1967 B.n733 B.n732 163.367
R1968 B.n732 B.n35 163.367
R1969 B.n728 B.n35 163.367
R1970 B.n728 B.n727 163.367
R1971 B.n727 B.n726 163.367
R1972 B.n726 B.n37 163.367
R1973 B.n722 B.n37 163.367
R1974 B.n722 B.n721 163.367
R1975 B.n721 B.n720 163.367
R1976 B.n720 B.n39 163.367
R1977 B.n716 B.n39 163.367
R1978 B.n716 B.n715 163.367
R1979 B.n715 B.n714 163.367
R1980 B.n714 B.n41 163.367
R1981 B.n710 B.n41 163.367
R1982 B.n710 B.n709 163.367
R1983 B.n709 B.n708 163.367
R1984 B.n708 B.n43 163.367
R1985 B.n704 B.n43 163.367
R1986 B.n704 B.n703 163.367
R1987 B.n703 B.n702 163.367
R1988 B.n702 B.n45 163.367
R1989 B.n698 B.n45 163.367
R1990 B.n698 B.n697 163.367
R1991 B.n697 B.n696 163.367
R1992 B.n696 B.n47 163.367
R1993 B.n692 B.n47 163.367
R1994 B.n692 B.n691 163.367
R1995 B.n691 B.n690 163.367
R1996 B.n690 B.n49 163.367
R1997 B.n686 B.n49 163.367
R1998 B.n686 B.n685 163.367
R1999 B.n685 B.n684 163.367
R2000 B.n684 B.n51 163.367
R2001 B.n680 B.n51 163.367
R2002 B.n680 B.n679 163.367
R2003 B.n679 B.n678 163.367
R2004 B.n678 B.n56 163.367
R2005 B.n674 B.n56 163.367
R2006 B.n674 B.n673 163.367
R2007 B.n673 B.n672 163.367
R2008 B.n672 B.n58 163.367
R2009 B.n667 B.n58 163.367
R2010 B.n667 B.n666 163.367
R2011 B.n666 B.n665 163.367
R2012 B.n665 B.n62 163.367
R2013 B.n661 B.n62 163.367
R2014 B.n661 B.n660 163.367
R2015 B.n660 B.n659 163.367
R2016 B.n659 B.n64 163.367
R2017 B.n655 B.n64 163.367
R2018 B.n655 B.n654 163.367
R2019 B.n654 B.n653 163.367
R2020 B.n653 B.n66 163.367
R2021 B.n649 B.n66 163.367
R2022 B.n649 B.n648 163.367
R2023 B.n648 B.n647 163.367
R2024 B.n647 B.n68 163.367
R2025 B.n643 B.n68 163.367
R2026 B.n643 B.n642 163.367
R2027 B.n642 B.n641 163.367
R2028 B.n641 B.n70 163.367
R2029 B.n637 B.n70 163.367
R2030 B.n637 B.n636 163.367
R2031 B.n636 B.n635 163.367
R2032 B.n635 B.n72 163.367
R2033 B.n631 B.n72 163.367
R2034 B.n631 B.n630 163.367
R2035 B.n630 B.n629 163.367
R2036 B.n629 B.n74 163.367
R2037 B.n625 B.n74 163.367
R2038 B.n625 B.n624 163.367
R2039 B.n624 B.n623 163.367
R2040 B.n623 B.n76 163.367
R2041 B.n619 B.n76 163.367
R2042 B.n619 B.n618 163.367
R2043 B.n618 B.n617 163.367
R2044 B.n617 B.n78 163.367
R2045 B.n613 B.n78 163.367
R2046 B.n613 B.n612 163.367
R2047 B.n612 B.n611 163.367
R2048 B.n611 B.n80 163.367
R2049 B.n607 B.n80 163.367
R2050 B.n607 B.n606 163.367
R2051 B.n606 B.n605 163.367
R2052 B.n605 B.n82 163.367
R2053 B.n601 B.n82 163.367
R2054 B.n601 B.n600 163.367
R2055 B.n600 B.n599 163.367
R2056 B.n599 B.n84 163.367
R2057 B.n595 B.n84 163.367
R2058 B.n595 B.n594 163.367
R2059 B.n594 B.n593 163.367
R2060 B.n593 B.n86 163.367
R2061 B.n589 B.n86 163.367
R2062 B.n589 B.n588 163.367
R2063 B.n588 B.n587 163.367
R2064 B.n587 B.n88 163.367
R2065 B.n583 B.n88 163.367
R2066 B.n583 B.n582 163.367
R2067 B.n160 B.n159 67.4914
R2068 B.n166 B.n165 67.4914
R2069 B.n53 B.n52 67.4914
R2070 B.n60 B.n59 67.4914
R2071 B.n375 B.n160 59.5399
R2072 B.n167 B.n166 59.5399
R2073 B.n54 B.n53 59.5399
R2074 B.n669 B.n60 59.5399
R2075 B.n772 B.n771 28.2542
R2076 B.n580 B.n89 28.2542
R2077 B.n464 B.n129 28.2542
R2078 B.n273 B.n272 28.2542
R2079 B B.n831 18.0485
R2080 B.n771 B.n22 10.6151
R2081 B.n767 B.n22 10.6151
R2082 B.n767 B.n766 10.6151
R2083 B.n766 B.n765 10.6151
R2084 B.n765 B.n24 10.6151
R2085 B.n761 B.n24 10.6151
R2086 B.n761 B.n760 10.6151
R2087 B.n760 B.n759 10.6151
R2088 B.n759 B.n26 10.6151
R2089 B.n755 B.n26 10.6151
R2090 B.n755 B.n754 10.6151
R2091 B.n754 B.n753 10.6151
R2092 B.n753 B.n28 10.6151
R2093 B.n749 B.n28 10.6151
R2094 B.n749 B.n748 10.6151
R2095 B.n748 B.n747 10.6151
R2096 B.n747 B.n30 10.6151
R2097 B.n743 B.n30 10.6151
R2098 B.n743 B.n742 10.6151
R2099 B.n742 B.n741 10.6151
R2100 B.n741 B.n32 10.6151
R2101 B.n737 B.n32 10.6151
R2102 B.n737 B.n736 10.6151
R2103 B.n736 B.n735 10.6151
R2104 B.n735 B.n34 10.6151
R2105 B.n731 B.n34 10.6151
R2106 B.n731 B.n730 10.6151
R2107 B.n730 B.n729 10.6151
R2108 B.n729 B.n36 10.6151
R2109 B.n725 B.n36 10.6151
R2110 B.n725 B.n724 10.6151
R2111 B.n724 B.n723 10.6151
R2112 B.n723 B.n38 10.6151
R2113 B.n719 B.n38 10.6151
R2114 B.n719 B.n718 10.6151
R2115 B.n718 B.n717 10.6151
R2116 B.n717 B.n40 10.6151
R2117 B.n713 B.n40 10.6151
R2118 B.n713 B.n712 10.6151
R2119 B.n712 B.n711 10.6151
R2120 B.n711 B.n42 10.6151
R2121 B.n707 B.n42 10.6151
R2122 B.n707 B.n706 10.6151
R2123 B.n706 B.n705 10.6151
R2124 B.n705 B.n44 10.6151
R2125 B.n701 B.n44 10.6151
R2126 B.n701 B.n700 10.6151
R2127 B.n700 B.n699 10.6151
R2128 B.n699 B.n46 10.6151
R2129 B.n695 B.n46 10.6151
R2130 B.n695 B.n694 10.6151
R2131 B.n694 B.n693 10.6151
R2132 B.n693 B.n48 10.6151
R2133 B.n689 B.n48 10.6151
R2134 B.n689 B.n688 10.6151
R2135 B.n688 B.n687 10.6151
R2136 B.n687 B.n50 10.6151
R2137 B.n683 B.n682 10.6151
R2138 B.n682 B.n681 10.6151
R2139 B.n681 B.n55 10.6151
R2140 B.n677 B.n55 10.6151
R2141 B.n677 B.n676 10.6151
R2142 B.n676 B.n675 10.6151
R2143 B.n675 B.n57 10.6151
R2144 B.n671 B.n57 10.6151
R2145 B.n671 B.n670 10.6151
R2146 B.n668 B.n61 10.6151
R2147 B.n664 B.n61 10.6151
R2148 B.n664 B.n663 10.6151
R2149 B.n663 B.n662 10.6151
R2150 B.n662 B.n63 10.6151
R2151 B.n658 B.n63 10.6151
R2152 B.n658 B.n657 10.6151
R2153 B.n657 B.n656 10.6151
R2154 B.n656 B.n65 10.6151
R2155 B.n652 B.n65 10.6151
R2156 B.n652 B.n651 10.6151
R2157 B.n651 B.n650 10.6151
R2158 B.n650 B.n67 10.6151
R2159 B.n646 B.n67 10.6151
R2160 B.n646 B.n645 10.6151
R2161 B.n645 B.n644 10.6151
R2162 B.n644 B.n69 10.6151
R2163 B.n640 B.n69 10.6151
R2164 B.n640 B.n639 10.6151
R2165 B.n639 B.n638 10.6151
R2166 B.n638 B.n71 10.6151
R2167 B.n634 B.n71 10.6151
R2168 B.n634 B.n633 10.6151
R2169 B.n633 B.n632 10.6151
R2170 B.n632 B.n73 10.6151
R2171 B.n628 B.n73 10.6151
R2172 B.n628 B.n627 10.6151
R2173 B.n627 B.n626 10.6151
R2174 B.n626 B.n75 10.6151
R2175 B.n622 B.n75 10.6151
R2176 B.n622 B.n621 10.6151
R2177 B.n621 B.n620 10.6151
R2178 B.n620 B.n77 10.6151
R2179 B.n616 B.n77 10.6151
R2180 B.n616 B.n615 10.6151
R2181 B.n615 B.n614 10.6151
R2182 B.n614 B.n79 10.6151
R2183 B.n610 B.n79 10.6151
R2184 B.n610 B.n609 10.6151
R2185 B.n609 B.n608 10.6151
R2186 B.n608 B.n81 10.6151
R2187 B.n604 B.n81 10.6151
R2188 B.n604 B.n603 10.6151
R2189 B.n603 B.n602 10.6151
R2190 B.n602 B.n83 10.6151
R2191 B.n598 B.n83 10.6151
R2192 B.n598 B.n597 10.6151
R2193 B.n597 B.n596 10.6151
R2194 B.n596 B.n85 10.6151
R2195 B.n592 B.n85 10.6151
R2196 B.n592 B.n591 10.6151
R2197 B.n591 B.n590 10.6151
R2198 B.n590 B.n87 10.6151
R2199 B.n586 B.n87 10.6151
R2200 B.n586 B.n585 10.6151
R2201 B.n585 B.n584 10.6151
R2202 B.n584 B.n89 10.6151
R2203 B.n465 B.n464 10.6151
R2204 B.n466 B.n465 10.6151
R2205 B.n466 B.n127 10.6151
R2206 B.n470 B.n127 10.6151
R2207 B.n471 B.n470 10.6151
R2208 B.n472 B.n471 10.6151
R2209 B.n472 B.n125 10.6151
R2210 B.n476 B.n125 10.6151
R2211 B.n477 B.n476 10.6151
R2212 B.n478 B.n477 10.6151
R2213 B.n478 B.n123 10.6151
R2214 B.n482 B.n123 10.6151
R2215 B.n483 B.n482 10.6151
R2216 B.n484 B.n483 10.6151
R2217 B.n484 B.n121 10.6151
R2218 B.n488 B.n121 10.6151
R2219 B.n489 B.n488 10.6151
R2220 B.n490 B.n489 10.6151
R2221 B.n490 B.n119 10.6151
R2222 B.n494 B.n119 10.6151
R2223 B.n495 B.n494 10.6151
R2224 B.n496 B.n495 10.6151
R2225 B.n496 B.n117 10.6151
R2226 B.n500 B.n117 10.6151
R2227 B.n501 B.n500 10.6151
R2228 B.n502 B.n501 10.6151
R2229 B.n502 B.n115 10.6151
R2230 B.n506 B.n115 10.6151
R2231 B.n507 B.n506 10.6151
R2232 B.n508 B.n507 10.6151
R2233 B.n508 B.n113 10.6151
R2234 B.n512 B.n113 10.6151
R2235 B.n513 B.n512 10.6151
R2236 B.n514 B.n513 10.6151
R2237 B.n514 B.n111 10.6151
R2238 B.n518 B.n111 10.6151
R2239 B.n519 B.n518 10.6151
R2240 B.n520 B.n519 10.6151
R2241 B.n520 B.n109 10.6151
R2242 B.n524 B.n109 10.6151
R2243 B.n525 B.n524 10.6151
R2244 B.n526 B.n525 10.6151
R2245 B.n526 B.n107 10.6151
R2246 B.n530 B.n107 10.6151
R2247 B.n531 B.n530 10.6151
R2248 B.n532 B.n531 10.6151
R2249 B.n532 B.n105 10.6151
R2250 B.n536 B.n105 10.6151
R2251 B.n537 B.n536 10.6151
R2252 B.n538 B.n537 10.6151
R2253 B.n538 B.n103 10.6151
R2254 B.n542 B.n103 10.6151
R2255 B.n543 B.n542 10.6151
R2256 B.n544 B.n543 10.6151
R2257 B.n544 B.n101 10.6151
R2258 B.n548 B.n101 10.6151
R2259 B.n549 B.n548 10.6151
R2260 B.n550 B.n549 10.6151
R2261 B.n550 B.n99 10.6151
R2262 B.n554 B.n99 10.6151
R2263 B.n555 B.n554 10.6151
R2264 B.n556 B.n555 10.6151
R2265 B.n556 B.n97 10.6151
R2266 B.n560 B.n97 10.6151
R2267 B.n561 B.n560 10.6151
R2268 B.n562 B.n561 10.6151
R2269 B.n562 B.n95 10.6151
R2270 B.n566 B.n95 10.6151
R2271 B.n567 B.n566 10.6151
R2272 B.n568 B.n567 10.6151
R2273 B.n568 B.n93 10.6151
R2274 B.n572 B.n93 10.6151
R2275 B.n573 B.n572 10.6151
R2276 B.n574 B.n573 10.6151
R2277 B.n574 B.n91 10.6151
R2278 B.n578 B.n91 10.6151
R2279 B.n579 B.n578 10.6151
R2280 B.n580 B.n579 10.6151
R2281 B.n274 B.n273 10.6151
R2282 B.n274 B.n195 10.6151
R2283 B.n278 B.n195 10.6151
R2284 B.n279 B.n278 10.6151
R2285 B.n280 B.n279 10.6151
R2286 B.n280 B.n193 10.6151
R2287 B.n284 B.n193 10.6151
R2288 B.n285 B.n284 10.6151
R2289 B.n286 B.n285 10.6151
R2290 B.n286 B.n191 10.6151
R2291 B.n290 B.n191 10.6151
R2292 B.n291 B.n290 10.6151
R2293 B.n292 B.n291 10.6151
R2294 B.n292 B.n189 10.6151
R2295 B.n296 B.n189 10.6151
R2296 B.n297 B.n296 10.6151
R2297 B.n298 B.n297 10.6151
R2298 B.n298 B.n187 10.6151
R2299 B.n302 B.n187 10.6151
R2300 B.n303 B.n302 10.6151
R2301 B.n304 B.n303 10.6151
R2302 B.n304 B.n185 10.6151
R2303 B.n308 B.n185 10.6151
R2304 B.n309 B.n308 10.6151
R2305 B.n310 B.n309 10.6151
R2306 B.n310 B.n183 10.6151
R2307 B.n314 B.n183 10.6151
R2308 B.n315 B.n314 10.6151
R2309 B.n316 B.n315 10.6151
R2310 B.n316 B.n181 10.6151
R2311 B.n320 B.n181 10.6151
R2312 B.n321 B.n320 10.6151
R2313 B.n322 B.n321 10.6151
R2314 B.n322 B.n179 10.6151
R2315 B.n326 B.n179 10.6151
R2316 B.n327 B.n326 10.6151
R2317 B.n328 B.n327 10.6151
R2318 B.n328 B.n177 10.6151
R2319 B.n332 B.n177 10.6151
R2320 B.n333 B.n332 10.6151
R2321 B.n334 B.n333 10.6151
R2322 B.n334 B.n175 10.6151
R2323 B.n338 B.n175 10.6151
R2324 B.n339 B.n338 10.6151
R2325 B.n340 B.n339 10.6151
R2326 B.n340 B.n173 10.6151
R2327 B.n344 B.n173 10.6151
R2328 B.n345 B.n344 10.6151
R2329 B.n346 B.n345 10.6151
R2330 B.n346 B.n171 10.6151
R2331 B.n350 B.n171 10.6151
R2332 B.n351 B.n350 10.6151
R2333 B.n352 B.n351 10.6151
R2334 B.n352 B.n169 10.6151
R2335 B.n356 B.n169 10.6151
R2336 B.n357 B.n356 10.6151
R2337 B.n358 B.n357 10.6151
R2338 B.n362 B.n361 10.6151
R2339 B.n363 B.n362 10.6151
R2340 B.n363 B.n163 10.6151
R2341 B.n367 B.n163 10.6151
R2342 B.n368 B.n367 10.6151
R2343 B.n369 B.n368 10.6151
R2344 B.n369 B.n161 10.6151
R2345 B.n373 B.n161 10.6151
R2346 B.n374 B.n373 10.6151
R2347 B.n376 B.n157 10.6151
R2348 B.n380 B.n157 10.6151
R2349 B.n381 B.n380 10.6151
R2350 B.n382 B.n381 10.6151
R2351 B.n382 B.n155 10.6151
R2352 B.n386 B.n155 10.6151
R2353 B.n387 B.n386 10.6151
R2354 B.n388 B.n387 10.6151
R2355 B.n388 B.n153 10.6151
R2356 B.n392 B.n153 10.6151
R2357 B.n393 B.n392 10.6151
R2358 B.n394 B.n393 10.6151
R2359 B.n394 B.n151 10.6151
R2360 B.n398 B.n151 10.6151
R2361 B.n399 B.n398 10.6151
R2362 B.n400 B.n399 10.6151
R2363 B.n400 B.n149 10.6151
R2364 B.n404 B.n149 10.6151
R2365 B.n405 B.n404 10.6151
R2366 B.n406 B.n405 10.6151
R2367 B.n406 B.n147 10.6151
R2368 B.n410 B.n147 10.6151
R2369 B.n411 B.n410 10.6151
R2370 B.n412 B.n411 10.6151
R2371 B.n412 B.n145 10.6151
R2372 B.n416 B.n145 10.6151
R2373 B.n417 B.n416 10.6151
R2374 B.n418 B.n417 10.6151
R2375 B.n418 B.n143 10.6151
R2376 B.n422 B.n143 10.6151
R2377 B.n423 B.n422 10.6151
R2378 B.n424 B.n423 10.6151
R2379 B.n424 B.n141 10.6151
R2380 B.n428 B.n141 10.6151
R2381 B.n429 B.n428 10.6151
R2382 B.n430 B.n429 10.6151
R2383 B.n430 B.n139 10.6151
R2384 B.n434 B.n139 10.6151
R2385 B.n435 B.n434 10.6151
R2386 B.n436 B.n435 10.6151
R2387 B.n436 B.n137 10.6151
R2388 B.n440 B.n137 10.6151
R2389 B.n441 B.n440 10.6151
R2390 B.n442 B.n441 10.6151
R2391 B.n442 B.n135 10.6151
R2392 B.n446 B.n135 10.6151
R2393 B.n447 B.n446 10.6151
R2394 B.n448 B.n447 10.6151
R2395 B.n448 B.n133 10.6151
R2396 B.n452 B.n133 10.6151
R2397 B.n453 B.n452 10.6151
R2398 B.n454 B.n453 10.6151
R2399 B.n454 B.n131 10.6151
R2400 B.n458 B.n131 10.6151
R2401 B.n459 B.n458 10.6151
R2402 B.n460 B.n459 10.6151
R2403 B.n460 B.n129 10.6151
R2404 B.n272 B.n197 10.6151
R2405 B.n268 B.n197 10.6151
R2406 B.n268 B.n267 10.6151
R2407 B.n267 B.n266 10.6151
R2408 B.n266 B.n199 10.6151
R2409 B.n262 B.n199 10.6151
R2410 B.n262 B.n261 10.6151
R2411 B.n261 B.n260 10.6151
R2412 B.n260 B.n201 10.6151
R2413 B.n256 B.n201 10.6151
R2414 B.n256 B.n255 10.6151
R2415 B.n255 B.n254 10.6151
R2416 B.n254 B.n203 10.6151
R2417 B.n250 B.n203 10.6151
R2418 B.n250 B.n249 10.6151
R2419 B.n249 B.n248 10.6151
R2420 B.n248 B.n205 10.6151
R2421 B.n244 B.n205 10.6151
R2422 B.n244 B.n243 10.6151
R2423 B.n243 B.n242 10.6151
R2424 B.n242 B.n207 10.6151
R2425 B.n238 B.n207 10.6151
R2426 B.n238 B.n237 10.6151
R2427 B.n237 B.n236 10.6151
R2428 B.n236 B.n209 10.6151
R2429 B.n232 B.n209 10.6151
R2430 B.n232 B.n231 10.6151
R2431 B.n231 B.n230 10.6151
R2432 B.n230 B.n211 10.6151
R2433 B.n226 B.n211 10.6151
R2434 B.n226 B.n225 10.6151
R2435 B.n225 B.n224 10.6151
R2436 B.n224 B.n213 10.6151
R2437 B.n220 B.n213 10.6151
R2438 B.n220 B.n219 10.6151
R2439 B.n219 B.n218 10.6151
R2440 B.n218 B.n215 10.6151
R2441 B.n215 B.n0 10.6151
R2442 B.n827 B.n1 10.6151
R2443 B.n827 B.n826 10.6151
R2444 B.n826 B.n825 10.6151
R2445 B.n825 B.n4 10.6151
R2446 B.n821 B.n4 10.6151
R2447 B.n821 B.n820 10.6151
R2448 B.n820 B.n819 10.6151
R2449 B.n819 B.n6 10.6151
R2450 B.n815 B.n6 10.6151
R2451 B.n815 B.n814 10.6151
R2452 B.n814 B.n813 10.6151
R2453 B.n813 B.n8 10.6151
R2454 B.n809 B.n8 10.6151
R2455 B.n809 B.n808 10.6151
R2456 B.n808 B.n807 10.6151
R2457 B.n807 B.n10 10.6151
R2458 B.n803 B.n10 10.6151
R2459 B.n803 B.n802 10.6151
R2460 B.n802 B.n801 10.6151
R2461 B.n801 B.n12 10.6151
R2462 B.n797 B.n12 10.6151
R2463 B.n797 B.n796 10.6151
R2464 B.n796 B.n795 10.6151
R2465 B.n795 B.n14 10.6151
R2466 B.n791 B.n14 10.6151
R2467 B.n791 B.n790 10.6151
R2468 B.n790 B.n789 10.6151
R2469 B.n789 B.n16 10.6151
R2470 B.n785 B.n16 10.6151
R2471 B.n785 B.n784 10.6151
R2472 B.n784 B.n783 10.6151
R2473 B.n783 B.n18 10.6151
R2474 B.n779 B.n18 10.6151
R2475 B.n779 B.n778 10.6151
R2476 B.n778 B.n777 10.6151
R2477 B.n777 B.n20 10.6151
R2478 B.n773 B.n20 10.6151
R2479 B.n773 B.n772 10.6151
R2480 B.n54 B.n50 9.36635
R2481 B.n669 B.n668 9.36635
R2482 B.n358 B.n167 9.36635
R2483 B.n376 B.n375 9.36635
R2484 B.n831 B.n0 2.81026
R2485 B.n831 B.n1 2.81026
R2486 B.n683 B.n54 1.24928
R2487 B.n670 B.n669 1.24928
R2488 B.n361 B.n167 1.24928
R2489 B.n375 B.n374 1.24928
C0 VDD1 VTAIL 6.76435f
C1 w_n3058_n4482# VP 5.79423f
C2 B VP 1.93579f
C3 VDD2 VTAIL 6.82224f
C4 VDD1 VN 0.149341f
C5 VDD2 VN 7.03441f
C6 VTAIL w_n3058_n4482# 5.22152f
C7 VTAIL B 7.06134f
C8 VTAIL VP 6.78155f
C9 VN w_n3058_n4482# 5.39972f
C10 VN B 1.27856f
C11 VDD1 VDD2 1.15992f
C12 VN VP 7.62397f
C13 VDD1 w_n3058_n4482# 1.70392f
C14 VDD1 B 1.50875f
C15 VN VTAIL 6.76745f
C16 VDD2 w_n3058_n4482# 1.77222f
C17 VDD1 VP 7.31334f
C18 VDD2 B 1.57003f
C19 VDD2 VP 0.429146f
C20 w_n3058_n4482# B 11.4835f
C21 VDD2 VSUBS 1.1628f
C22 VDD1 VSUBS 6.74302f
C23 VTAIL VSUBS 1.539109f
C24 VN VSUBS 5.93655f
C25 VP VSUBS 2.779254f
C26 B VSUBS 5.220204f
C27 w_n3058_n4482# VSUBS 0.167664p
C28 B.n0 VSUBS 0.003663f
C29 B.n1 VSUBS 0.003663f
C30 B.n2 VSUBS 0.005793f
C31 B.n3 VSUBS 0.005793f
C32 B.n4 VSUBS 0.005793f
C33 B.n5 VSUBS 0.005793f
C34 B.n6 VSUBS 0.005793f
C35 B.n7 VSUBS 0.005793f
C36 B.n8 VSUBS 0.005793f
C37 B.n9 VSUBS 0.005793f
C38 B.n10 VSUBS 0.005793f
C39 B.n11 VSUBS 0.005793f
C40 B.n12 VSUBS 0.005793f
C41 B.n13 VSUBS 0.005793f
C42 B.n14 VSUBS 0.005793f
C43 B.n15 VSUBS 0.005793f
C44 B.n16 VSUBS 0.005793f
C45 B.n17 VSUBS 0.005793f
C46 B.n18 VSUBS 0.005793f
C47 B.n19 VSUBS 0.005793f
C48 B.n20 VSUBS 0.005793f
C49 B.n21 VSUBS 0.011957f
C50 B.n22 VSUBS 0.005793f
C51 B.n23 VSUBS 0.005793f
C52 B.n24 VSUBS 0.005793f
C53 B.n25 VSUBS 0.005793f
C54 B.n26 VSUBS 0.005793f
C55 B.n27 VSUBS 0.005793f
C56 B.n28 VSUBS 0.005793f
C57 B.n29 VSUBS 0.005793f
C58 B.n30 VSUBS 0.005793f
C59 B.n31 VSUBS 0.005793f
C60 B.n32 VSUBS 0.005793f
C61 B.n33 VSUBS 0.005793f
C62 B.n34 VSUBS 0.005793f
C63 B.n35 VSUBS 0.005793f
C64 B.n36 VSUBS 0.005793f
C65 B.n37 VSUBS 0.005793f
C66 B.n38 VSUBS 0.005793f
C67 B.n39 VSUBS 0.005793f
C68 B.n40 VSUBS 0.005793f
C69 B.n41 VSUBS 0.005793f
C70 B.n42 VSUBS 0.005793f
C71 B.n43 VSUBS 0.005793f
C72 B.n44 VSUBS 0.005793f
C73 B.n45 VSUBS 0.005793f
C74 B.n46 VSUBS 0.005793f
C75 B.n47 VSUBS 0.005793f
C76 B.n48 VSUBS 0.005793f
C77 B.n49 VSUBS 0.005793f
C78 B.n50 VSUBS 0.005452f
C79 B.n51 VSUBS 0.005793f
C80 B.t11 VSUBS 0.282006f
C81 B.t10 VSUBS 0.314452f
C82 B.t9 VSUBS 2.06345f
C83 B.n52 VSUBS 0.493655f
C84 B.n53 VSUBS 0.269562f
C85 B.n54 VSUBS 0.013421f
C86 B.n55 VSUBS 0.005793f
C87 B.n56 VSUBS 0.005793f
C88 B.n57 VSUBS 0.005793f
C89 B.n58 VSUBS 0.005793f
C90 B.t2 VSUBS 0.282009f
C91 B.t1 VSUBS 0.314455f
C92 B.t0 VSUBS 2.06345f
C93 B.n59 VSUBS 0.493652f
C94 B.n60 VSUBS 0.269559f
C95 B.n61 VSUBS 0.005793f
C96 B.n62 VSUBS 0.005793f
C97 B.n63 VSUBS 0.005793f
C98 B.n64 VSUBS 0.005793f
C99 B.n65 VSUBS 0.005793f
C100 B.n66 VSUBS 0.005793f
C101 B.n67 VSUBS 0.005793f
C102 B.n68 VSUBS 0.005793f
C103 B.n69 VSUBS 0.005793f
C104 B.n70 VSUBS 0.005793f
C105 B.n71 VSUBS 0.005793f
C106 B.n72 VSUBS 0.005793f
C107 B.n73 VSUBS 0.005793f
C108 B.n74 VSUBS 0.005793f
C109 B.n75 VSUBS 0.005793f
C110 B.n76 VSUBS 0.005793f
C111 B.n77 VSUBS 0.005793f
C112 B.n78 VSUBS 0.005793f
C113 B.n79 VSUBS 0.005793f
C114 B.n80 VSUBS 0.005793f
C115 B.n81 VSUBS 0.005793f
C116 B.n82 VSUBS 0.005793f
C117 B.n83 VSUBS 0.005793f
C118 B.n84 VSUBS 0.005793f
C119 B.n85 VSUBS 0.005793f
C120 B.n86 VSUBS 0.005793f
C121 B.n87 VSUBS 0.005793f
C122 B.n88 VSUBS 0.005793f
C123 B.n89 VSUBS 0.011957f
C124 B.n90 VSUBS 0.005793f
C125 B.n91 VSUBS 0.005793f
C126 B.n92 VSUBS 0.005793f
C127 B.n93 VSUBS 0.005793f
C128 B.n94 VSUBS 0.005793f
C129 B.n95 VSUBS 0.005793f
C130 B.n96 VSUBS 0.005793f
C131 B.n97 VSUBS 0.005793f
C132 B.n98 VSUBS 0.005793f
C133 B.n99 VSUBS 0.005793f
C134 B.n100 VSUBS 0.005793f
C135 B.n101 VSUBS 0.005793f
C136 B.n102 VSUBS 0.005793f
C137 B.n103 VSUBS 0.005793f
C138 B.n104 VSUBS 0.005793f
C139 B.n105 VSUBS 0.005793f
C140 B.n106 VSUBS 0.005793f
C141 B.n107 VSUBS 0.005793f
C142 B.n108 VSUBS 0.005793f
C143 B.n109 VSUBS 0.005793f
C144 B.n110 VSUBS 0.005793f
C145 B.n111 VSUBS 0.005793f
C146 B.n112 VSUBS 0.005793f
C147 B.n113 VSUBS 0.005793f
C148 B.n114 VSUBS 0.005793f
C149 B.n115 VSUBS 0.005793f
C150 B.n116 VSUBS 0.005793f
C151 B.n117 VSUBS 0.005793f
C152 B.n118 VSUBS 0.005793f
C153 B.n119 VSUBS 0.005793f
C154 B.n120 VSUBS 0.005793f
C155 B.n121 VSUBS 0.005793f
C156 B.n122 VSUBS 0.005793f
C157 B.n123 VSUBS 0.005793f
C158 B.n124 VSUBS 0.005793f
C159 B.n125 VSUBS 0.005793f
C160 B.n126 VSUBS 0.005793f
C161 B.n127 VSUBS 0.005793f
C162 B.n128 VSUBS 0.005793f
C163 B.n129 VSUBS 0.012748f
C164 B.n130 VSUBS 0.005793f
C165 B.n131 VSUBS 0.005793f
C166 B.n132 VSUBS 0.005793f
C167 B.n133 VSUBS 0.005793f
C168 B.n134 VSUBS 0.005793f
C169 B.n135 VSUBS 0.005793f
C170 B.n136 VSUBS 0.005793f
C171 B.n137 VSUBS 0.005793f
C172 B.n138 VSUBS 0.005793f
C173 B.n139 VSUBS 0.005793f
C174 B.n140 VSUBS 0.005793f
C175 B.n141 VSUBS 0.005793f
C176 B.n142 VSUBS 0.005793f
C177 B.n143 VSUBS 0.005793f
C178 B.n144 VSUBS 0.005793f
C179 B.n145 VSUBS 0.005793f
C180 B.n146 VSUBS 0.005793f
C181 B.n147 VSUBS 0.005793f
C182 B.n148 VSUBS 0.005793f
C183 B.n149 VSUBS 0.005793f
C184 B.n150 VSUBS 0.005793f
C185 B.n151 VSUBS 0.005793f
C186 B.n152 VSUBS 0.005793f
C187 B.n153 VSUBS 0.005793f
C188 B.n154 VSUBS 0.005793f
C189 B.n155 VSUBS 0.005793f
C190 B.n156 VSUBS 0.005793f
C191 B.n157 VSUBS 0.005793f
C192 B.n158 VSUBS 0.005793f
C193 B.t4 VSUBS 0.282009f
C194 B.t5 VSUBS 0.314455f
C195 B.t3 VSUBS 2.06345f
C196 B.n159 VSUBS 0.493652f
C197 B.n160 VSUBS 0.269559f
C198 B.n161 VSUBS 0.005793f
C199 B.n162 VSUBS 0.005793f
C200 B.n163 VSUBS 0.005793f
C201 B.n164 VSUBS 0.005793f
C202 B.t7 VSUBS 0.282006f
C203 B.t8 VSUBS 0.314452f
C204 B.t6 VSUBS 2.06345f
C205 B.n165 VSUBS 0.493655f
C206 B.n166 VSUBS 0.269562f
C207 B.n167 VSUBS 0.013421f
C208 B.n168 VSUBS 0.005793f
C209 B.n169 VSUBS 0.005793f
C210 B.n170 VSUBS 0.005793f
C211 B.n171 VSUBS 0.005793f
C212 B.n172 VSUBS 0.005793f
C213 B.n173 VSUBS 0.005793f
C214 B.n174 VSUBS 0.005793f
C215 B.n175 VSUBS 0.005793f
C216 B.n176 VSUBS 0.005793f
C217 B.n177 VSUBS 0.005793f
C218 B.n178 VSUBS 0.005793f
C219 B.n179 VSUBS 0.005793f
C220 B.n180 VSUBS 0.005793f
C221 B.n181 VSUBS 0.005793f
C222 B.n182 VSUBS 0.005793f
C223 B.n183 VSUBS 0.005793f
C224 B.n184 VSUBS 0.005793f
C225 B.n185 VSUBS 0.005793f
C226 B.n186 VSUBS 0.005793f
C227 B.n187 VSUBS 0.005793f
C228 B.n188 VSUBS 0.005793f
C229 B.n189 VSUBS 0.005793f
C230 B.n190 VSUBS 0.005793f
C231 B.n191 VSUBS 0.005793f
C232 B.n192 VSUBS 0.005793f
C233 B.n193 VSUBS 0.005793f
C234 B.n194 VSUBS 0.005793f
C235 B.n195 VSUBS 0.005793f
C236 B.n196 VSUBS 0.012748f
C237 B.n197 VSUBS 0.005793f
C238 B.n198 VSUBS 0.005793f
C239 B.n199 VSUBS 0.005793f
C240 B.n200 VSUBS 0.005793f
C241 B.n201 VSUBS 0.005793f
C242 B.n202 VSUBS 0.005793f
C243 B.n203 VSUBS 0.005793f
C244 B.n204 VSUBS 0.005793f
C245 B.n205 VSUBS 0.005793f
C246 B.n206 VSUBS 0.005793f
C247 B.n207 VSUBS 0.005793f
C248 B.n208 VSUBS 0.005793f
C249 B.n209 VSUBS 0.005793f
C250 B.n210 VSUBS 0.005793f
C251 B.n211 VSUBS 0.005793f
C252 B.n212 VSUBS 0.005793f
C253 B.n213 VSUBS 0.005793f
C254 B.n214 VSUBS 0.005793f
C255 B.n215 VSUBS 0.005793f
C256 B.n216 VSUBS 0.005793f
C257 B.n217 VSUBS 0.005793f
C258 B.n218 VSUBS 0.005793f
C259 B.n219 VSUBS 0.005793f
C260 B.n220 VSUBS 0.005793f
C261 B.n221 VSUBS 0.005793f
C262 B.n222 VSUBS 0.005793f
C263 B.n223 VSUBS 0.005793f
C264 B.n224 VSUBS 0.005793f
C265 B.n225 VSUBS 0.005793f
C266 B.n226 VSUBS 0.005793f
C267 B.n227 VSUBS 0.005793f
C268 B.n228 VSUBS 0.005793f
C269 B.n229 VSUBS 0.005793f
C270 B.n230 VSUBS 0.005793f
C271 B.n231 VSUBS 0.005793f
C272 B.n232 VSUBS 0.005793f
C273 B.n233 VSUBS 0.005793f
C274 B.n234 VSUBS 0.005793f
C275 B.n235 VSUBS 0.005793f
C276 B.n236 VSUBS 0.005793f
C277 B.n237 VSUBS 0.005793f
C278 B.n238 VSUBS 0.005793f
C279 B.n239 VSUBS 0.005793f
C280 B.n240 VSUBS 0.005793f
C281 B.n241 VSUBS 0.005793f
C282 B.n242 VSUBS 0.005793f
C283 B.n243 VSUBS 0.005793f
C284 B.n244 VSUBS 0.005793f
C285 B.n245 VSUBS 0.005793f
C286 B.n246 VSUBS 0.005793f
C287 B.n247 VSUBS 0.005793f
C288 B.n248 VSUBS 0.005793f
C289 B.n249 VSUBS 0.005793f
C290 B.n250 VSUBS 0.005793f
C291 B.n251 VSUBS 0.005793f
C292 B.n252 VSUBS 0.005793f
C293 B.n253 VSUBS 0.005793f
C294 B.n254 VSUBS 0.005793f
C295 B.n255 VSUBS 0.005793f
C296 B.n256 VSUBS 0.005793f
C297 B.n257 VSUBS 0.005793f
C298 B.n258 VSUBS 0.005793f
C299 B.n259 VSUBS 0.005793f
C300 B.n260 VSUBS 0.005793f
C301 B.n261 VSUBS 0.005793f
C302 B.n262 VSUBS 0.005793f
C303 B.n263 VSUBS 0.005793f
C304 B.n264 VSUBS 0.005793f
C305 B.n265 VSUBS 0.005793f
C306 B.n266 VSUBS 0.005793f
C307 B.n267 VSUBS 0.005793f
C308 B.n268 VSUBS 0.005793f
C309 B.n269 VSUBS 0.005793f
C310 B.n270 VSUBS 0.005793f
C311 B.n271 VSUBS 0.011957f
C312 B.n272 VSUBS 0.011957f
C313 B.n273 VSUBS 0.012748f
C314 B.n274 VSUBS 0.005793f
C315 B.n275 VSUBS 0.005793f
C316 B.n276 VSUBS 0.005793f
C317 B.n277 VSUBS 0.005793f
C318 B.n278 VSUBS 0.005793f
C319 B.n279 VSUBS 0.005793f
C320 B.n280 VSUBS 0.005793f
C321 B.n281 VSUBS 0.005793f
C322 B.n282 VSUBS 0.005793f
C323 B.n283 VSUBS 0.005793f
C324 B.n284 VSUBS 0.005793f
C325 B.n285 VSUBS 0.005793f
C326 B.n286 VSUBS 0.005793f
C327 B.n287 VSUBS 0.005793f
C328 B.n288 VSUBS 0.005793f
C329 B.n289 VSUBS 0.005793f
C330 B.n290 VSUBS 0.005793f
C331 B.n291 VSUBS 0.005793f
C332 B.n292 VSUBS 0.005793f
C333 B.n293 VSUBS 0.005793f
C334 B.n294 VSUBS 0.005793f
C335 B.n295 VSUBS 0.005793f
C336 B.n296 VSUBS 0.005793f
C337 B.n297 VSUBS 0.005793f
C338 B.n298 VSUBS 0.005793f
C339 B.n299 VSUBS 0.005793f
C340 B.n300 VSUBS 0.005793f
C341 B.n301 VSUBS 0.005793f
C342 B.n302 VSUBS 0.005793f
C343 B.n303 VSUBS 0.005793f
C344 B.n304 VSUBS 0.005793f
C345 B.n305 VSUBS 0.005793f
C346 B.n306 VSUBS 0.005793f
C347 B.n307 VSUBS 0.005793f
C348 B.n308 VSUBS 0.005793f
C349 B.n309 VSUBS 0.005793f
C350 B.n310 VSUBS 0.005793f
C351 B.n311 VSUBS 0.005793f
C352 B.n312 VSUBS 0.005793f
C353 B.n313 VSUBS 0.005793f
C354 B.n314 VSUBS 0.005793f
C355 B.n315 VSUBS 0.005793f
C356 B.n316 VSUBS 0.005793f
C357 B.n317 VSUBS 0.005793f
C358 B.n318 VSUBS 0.005793f
C359 B.n319 VSUBS 0.005793f
C360 B.n320 VSUBS 0.005793f
C361 B.n321 VSUBS 0.005793f
C362 B.n322 VSUBS 0.005793f
C363 B.n323 VSUBS 0.005793f
C364 B.n324 VSUBS 0.005793f
C365 B.n325 VSUBS 0.005793f
C366 B.n326 VSUBS 0.005793f
C367 B.n327 VSUBS 0.005793f
C368 B.n328 VSUBS 0.005793f
C369 B.n329 VSUBS 0.005793f
C370 B.n330 VSUBS 0.005793f
C371 B.n331 VSUBS 0.005793f
C372 B.n332 VSUBS 0.005793f
C373 B.n333 VSUBS 0.005793f
C374 B.n334 VSUBS 0.005793f
C375 B.n335 VSUBS 0.005793f
C376 B.n336 VSUBS 0.005793f
C377 B.n337 VSUBS 0.005793f
C378 B.n338 VSUBS 0.005793f
C379 B.n339 VSUBS 0.005793f
C380 B.n340 VSUBS 0.005793f
C381 B.n341 VSUBS 0.005793f
C382 B.n342 VSUBS 0.005793f
C383 B.n343 VSUBS 0.005793f
C384 B.n344 VSUBS 0.005793f
C385 B.n345 VSUBS 0.005793f
C386 B.n346 VSUBS 0.005793f
C387 B.n347 VSUBS 0.005793f
C388 B.n348 VSUBS 0.005793f
C389 B.n349 VSUBS 0.005793f
C390 B.n350 VSUBS 0.005793f
C391 B.n351 VSUBS 0.005793f
C392 B.n352 VSUBS 0.005793f
C393 B.n353 VSUBS 0.005793f
C394 B.n354 VSUBS 0.005793f
C395 B.n355 VSUBS 0.005793f
C396 B.n356 VSUBS 0.005793f
C397 B.n357 VSUBS 0.005793f
C398 B.n358 VSUBS 0.005452f
C399 B.n359 VSUBS 0.005793f
C400 B.n360 VSUBS 0.005793f
C401 B.n361 VSUBS 0.003237f
C402 B.n362 VSUBS 0.005793f
C403 B.n363 VSUBS 0.005793f
C404 B.n364 VSUBS 0.005793f
C405 B.n365 VSUBS 0.005793f
C406 B.n366 VSUBS 0.005793f
C407 B.n367 VSUBS 0.005793f
C408 B.n368 VSUBS 0.005793f
C409 B.n369 VSUBS 0.005793f
C410 B.n370 VSUBS 0.005793f
C411 B.n371 VSUBS 0.005793f
C412 B.n372 VSUBS 0.005793f
C413 B.n373 VSUBS 0.005793f
C414 B.n374 VSUBS 0.003237f
C415 B.n375 VSUBS 0.013421f
C416 B.n376 VSUBS 0.005452f
C417 B.n377 VSUBS 0.005793f
C418 B.n378 VSUBS 0.005793f
C419 B.n379 VSUBS 0.005793f
C420 B.n380 VSUBS 0.005793f
C421 B.n381 VSUBS 0.005793f
C422 B.n382 VSUBS 0.005793f
C423 B.n383 VSUBS 0.005793f
C424 B.n384 VSUBS 0.005793f
C425 B.n385 VSUBS 0.005793f
C426 B.n386 VSUBS 0.005793f
C427 B.n387 VSUBS 0.005793f
C428 B.n388 VSUBS 0.005793f
C429 B.n389 VSUBS 0.005793f
C430 B.n390 VSUBS 0.005793f
C431 B.n391 VSUBS 0.005793f
C432 B.n392 VSUBS 0.005793f
C433 B.n393 VSUBS 0.005793f
C434 B.n394 VSUBS 0.005793f
C435 B.n395 VSUBS 0.005793f
C436 B.n396 VSUBS 0.005793f
C437 B.n397 VSUBS 0.005793f
C438 B.n398 VSUBS 0.005793f
C439 B.n399 VSUBS 0.005793f
C440 B.n400 VSUBS 0.005793f
C441 B.n401 VSUBS 0.005793f
C442 B.n402 VSUBS 0.005793f
C443 B.n403 VSUBS 0.005793f
C444 B.n404 VSUBS 0.005793f
C445 B.n405 VSUBS 0.005793f
C446 B.n406 VSUBS 0.005793f
C447 B.n407 VSUBS 0.005793f
C448 B.n408 VSUBS 0.005793f
C449 B.n409 VSUBS 0.005793f
C450 B.n410 VSUBS 0.005793f
C451 B.n411 VSUBS 0.005793f
C452 B.n412 VSUBS 0.005793f
C453 B.n413 VSUBS 0.005793f
C454 B.n414 VSUBS 0.005793f
C455 B.n415 VSUBS 0.005793f
C456 B.n416 VSUBS 0.005793f
C457 B.n417 VSUBS 0.005793f
C458 B.n418 VSUBS 0.005793f
C459 B.n419 VSUBS 0.005793f
C460 B.n420 VSUBS 0.005793f
C461 B.n421 VSUBS 0.005793f
C462 B.n422 VSUBS 0.005793f
C463 B.n423 VSUBS 0.005793f
C464 B.n424 VSUBS 0.005793f
C465 B.n425 VSUBS 0.005793f
C466 B.n426 VSUBS 0.005793f
C467 B.n427 VSUBS 0.005793f
C468 B.n428 VSUBS 0.005793f
C469 B.n429 VSUBS 0.005793f
C470 B.n430 VSUBS 0.005793f
C471 B.n431 VSUBS 0.005793f
C472 B.n432 VSUBS 0.005793f
C473 B.n433 VSUBS 0.005793f
C474 B.n434 VSUBS 0.005793f
C475 B.n435 VSUBS 0.005793f
C476 B.n436 VSUBS 0.005793f
C477 B.n437 VSUBS 0.005793f
C478 B.n438 VSUBS 0.005793f
C479 B.n439 VSUBS 0.005793f
C480 B.n440 VSUBS 0.005793f
C481 B.n441 VSUBS 0.005793f
C482 B.n442 VSUBS 0.005793f
C483 B.n443 VSUBS 0.005793f
C484 B.n444 VSUBS 0.005793f
C485 B.n445 VSUBS 0.005793f
C486 B.n446 VSUBS 0.005793f
C487 B.n447 VSUBS 0.005793f
C488 B.n448 VSUBS 0.005793f
C489 B.n449 VSUBS 0.005793f
C490 B.n450 VSUBS 0.005793f
C491 B.n451 VSUBS 0.005793f
C492 B.n452 VSUBS 0.005793f
C493 B.n453 VSUBS 0.005793f
C494 B.n454 VSUBS 0.005793f
C495 B.n455 VSUBS 0.005793f
C496 B.n456 VSUBS 0.005793f
C497 B.n457 VSUBS 0.005793f
C498 B.n458 VSUBS 0.005793f
C499 B.n459 VSUBS 0.005793f
C500 B.n460 VSUBS 0.005793f
C501 B.n461 VSUBS 0.005793f
C502 B.n462 VSUBS 0.012748f
C503 B.n463 VSUBS 0.011957f
C504 B.n464 VSUBS 0.011957f
C505 B.n465 VSUBS 0.005793f
C506 B.n466 VSUBS 0.005793f
C507 B.n467 VSUBS 0.005793f
C508 B.n468 VSUBS 0.005793f
C509 B.n469 VSUBS 0.005793f
C510 B.n470 VSUBS 0.005793f
C511 B.n471 VSUBS 0.005793f
C512 B.n472 VSUBS 0.005793f
C513 B.n473 VSUBS 0.005793f
C514 B.n474 VSUBS 0.005793f
C515 B.n475 VSUBS 0.005793f
C516 B.n476 VSUBS 0.005793f
C517 B.n477 VSUBS 0.005793f
C518 B.n478 VSUBS 0.005793f
C519 B.n479 VSUBS 0.005793f
C520 B.n480 VSUBS 0.005793f
C521 B.n481 VSUBS 0.005793f
C522 B.n482 VSUBS 0.005793f
C523 B.n483 VSUBS 0.005793f
C524 B.n484 VSUBS 0.005793f
C525 B.n485 VSUBS 0.005793f
C526 B.n486 VSUBS 0.005793f
C527 B.n487 VSUBS 0.005793f
C528 B.n488 VSUBS 0.005793f
C529 B.n489 VSUBS 0.005793f
C530 B.n490 VSUBS 0.005793f
C531 B.n491 VSUBS 0.005793f
C532 B.n492 VSUBS 0.005793f
C533 B.n493 VSUBS 0.005793f
C534 B.n494 VSUBS 0.005793f
C535 B.n495 VSUBS 0.005793f
C536 B.n496 VSUBS 0.005793f
C537 B.n497 VSUBS 0.005793f
C538 B.n498 VSUBS 0.005793f
C539 B.n499 VSUBS 0.005793f
C540 B.n500 VSUBS 0.005793f
C541 B.n501 VSUBS 0.005793f
C542 B.n502 VSUBS 0.005793f
C543 B.n503 VSUBS 0.005793f
C544 B.n504 VSUBS 0.005793f
C545 B.n505 VSUBS 0.005793f
C546 B.n506 VSUBS 0.005793f
C547 B.n507 VSUBS 0.005793f
C548 B.n508 VSUBS 0.005793f
C549 B.n509 VSUBS 0.005793f
C550 B.n510 VSUBS 0.005793f
C551 B.n511 VSUBS 0.005793f
C552 B.n512 VSUBS 0.005793f
C553 B.n513 VSUBS 0.005793f
C554 B.n514 VSUBS 0.005793f
C555 B.n515 VSUBS 0.005793f
C556 B.n516 VSUBS 0.005793f
C557 B.n517 VSUBS 0.005793f
C558 B.n518 VSUBS 0.005793f
C559 B.n519 VSUBS 0.005793f
C560 B.n520 VSUBS 0.005793f
C561 B.n521 VSUBS 0.005793f
C562 B.n522 VSUBS 0.005793f
C563 B.n523 VSUBS 0.005793f
C564 B.n524 VSUBS 0.005793f
C565 B.n525 VSUBS 0.005793f
C566 B.n526 VSUBS 0.005793f
C567 B.n527 VSUBS 0.005793f
C568 B.n528 VSUBS 0.005793f
C569 B.n529 VSUBS 0.005793f
C570 B.n530 VSUBS 0.005793f
C571 B.n531 VSUBS 0.005793f
C572 B.n532 VSUBS 0.005793f
C573 B.n533 VSUBS 0.005793f
C574 B.n534 VSUBS 0.005793f
C575 B.n535 VSUBS 0.005793f
C576 B.n536 VSUBS 0.005793f
C577 B.n537 VSUBS 0.005793f
C578 B.n538 VSUBS 0.005793f
C579 B.n539 VSUBS 0.005793f
C580 B.n540 VSUBS 0.005793f
C581 B.n541 VSUBS 0.005793f
C582 B.n542 VSUBS 0.005793f
C583 B.n543 VSUBS 0.005793f
C584 B.n544 VSUBS 0.005793f
C585 B.n545 VSUBS 0.005793f
C586 B.n546 VSUBS 0.005793f
C587 B.n547 VSUBS 0.005793f
C588 B.n548 VSUBS 0.005793f
C589 B.n549 VSUBS 0.005793f
C590 B.n550 VSUBS 0.005793f
C591 B.n551 VSUBS 0.005793f
C592 B.n552 VSUBS 0.005793f
C593 B.n553 VSUBS 0.005793f
C594 B.n554 VSUBS 0.005793f
C595 B.n555 VSUBS 0.005793f
C596 B.n556 VSUBS 0.005793f
C597 B.n557 VSUBS 0.005793f
C598 B.n558 VSUBS 0.005793f
C599 B.n559 VSUBS 0.005793f
C600 B.n560 VSUBS 0.005793f
C601 B.n561 VSUBS 0.005793f
C602 B.n562 VSUBS 0.005793f
C603 B.n563 VSUBS 0.005793f
C604 B.n564 VSUBS 0.005793f
C605 B.n565 VSUBS 0.005793f
C606 B.n566 VSUBS 0.005793f
C607 B.n567 VSUBS 0.005793f
C608 B.n568 VSUBS 0.005793f
C609 B.n569 VSUBS 0.005793f
C610 B.n570 VSUBS 0.005793f
C611 B.n571 VSUBS 0.005793f
C612 B.n572 VSUBS 0.005793f
C613 B.n573 VSUBS 0.005793f
C614 B.n574 VSUBS 0.005793f
C615 B.n575 VSUBS 0.005793f
C616 B.n576 VSUBS 0.005793f
C617 B.n577 VSUBS 0.005793f
C618 B.n578 VSUBS 0.005793f
C619 B.n579 VSUBS 0.005793f
C620 B.n580 VSUBS 0.012748f
C621 B.n581 VSUBS 0.011957f
C622 B.n582 VSUBS 0.012748f
C623 B.n583 VSUBS 0.005793f
C624 B.n584 VSUBS 0.005793f
C625 B.n585 VSUBS 0.005793f
C626 B.n586 VSUBS 0.005793f
C627 B.n587 VSUBS 0.005793f
C628 B.n588 VSUBS 0.005793f
C629 B.n589 VSUBS 0.005793f
C630 B.n590 VSUBS 0.005793f
C631 B.n591 VSUBS 0.005793f
C632 B.n592 VSUBS 0.005793f
C633 B.n593 VSUBS 0.005793f
C634 B.n594 VSUBS 0.005793f
C635 B.n595 VSUBS 0.005793f
C636 B.n596 VSUBS 0.005793f
C637 B.n597 VSUBS 0.005793f
C638 B.n598 VSUBS 0.005793f
C639 B.n599 VSUBS 0.005793f
C640 B.n600 VSUBS 0.005793f
C641 B.n601 VSUBS 0.005793f
C642 B.n602 VSUBS 0.005793f
C643 B.n603 VSUBS 0.005793f
C644 B.n604 VSUBS 0.005793f
C645 B.n605 VSUBS 0.005793f
C646 B.n606 VSUBS 0.005793f
C647 B.n607 VSUBS 0.005793f
C648 B.n608 VSUBS 0.005793f
C649 B.n609 VSUBS 0.005793f
C650 B.n610 VSUBS 0.005793f
C651 B.n611 VSUBS 0.005793f
C652 B.n612 VSUBS 0.005793f
C653 B.n613 VSUBS 0.005793f
C654 B.n614 VSUBS 0.005793f
C655 B.n615 VSUBS 0.005793f
C656 B.n616 VSUBS 0.005793f
C657 B.n617 VSUBS 0.005793f
C658 B.n618 VSUBS 0.005793f
C659 B.n619 VSUBS 0.005793f
C660 B.n620 VSUBS 0.005793f
C661 B.n621 VSUBS 0.005793f
C662 B.n622 VSUBS 0.005793f
C663 B.n623 VSUBS 0.005793f
C664 B.n624 VSUBS 0.005793f
C665 B.n625 VSUBS 0.005793f
C666 B.n626 VSUBS 0.005793f
C667 B.n627 VSUBS 0.005793f
C668 B.n628 VSUBS 0.005793f
C669 B.n629 VSUBS 0.005793f
C670 B.n630 VSUBS 0.005793f
C671 B.n631 VSUBS 0.005793f
C672 B.n632 VSUBS 0.005793f
C673 B.n633 VSUBS 0.005793f
C674 B.n634 VSUBS 0.005793f
C675 B.n635 VSUBS 0.005793f
C676 B.n636 VSUBS 0.005793f
C677 B.n637 VSUBS 0.005793f
C678 B.n638 VSUBS 0.005793f
C679 B.n639 VSUBS 0.005793f
C680 B.n640 VSUBS 0.005793f
C681 B.n641 VSUBS 0.005793f
C682 B.n642 VSUBS 0.005793f
C683 B.n643 VSUBS 0.005793f
C684 B.n644 VSUBS 0.005793f
C685 B.n645 VSUBS 0.005793f
C686 B.n646 VSUBS 0.005793f
C687 B.n647 VSUBS 0.005793f
C688 B.n648 VSUBS 0.005793f
C689 B.n649 VSUBS 0.005793f
C690 B.n650 VSUBS 0.005793f
C691 B.n651 VSUBS 0.005793f
C692 B.n652 VSUBS 0.005793f
C693 B.n653 VSUBS 0.005793f
C694 B.n654 VSUBS 0.005793f
C695 B.n655 VSUBS 0.005793f
C696 B.n656 VSUBS 0.005793f
C697 B.n657 VSUBS 0.005793f
C698 B.n658 VSUBS 0.005793f
C699 B.n659 VSUBS 0.005793f
C700 B.n660 VSUBS 0.005793f
C701 B.n661 VSUBS 0.005793f
C702 B.n662 VSUBS 0.005793f
C703 B.n663 VSUBS 0.005793f
C704 B.n664 VSUBS 0.005793f
C705 B.n665 VSUBS 0.005793f
C706 B.n666 VSUBS 0.005793f
C707 B.n667 VSUBS 0.005793f
C708 B.n668 VSUBS 0.005452f
C709 B.n669 VSUBS 0.013421f
C710 B.n670 VSUBS 0.003237f
C711 B.n671 VSUBS 0.005793f
C712 B.n672 VSUBS 0.005793f
C713 B.n673 VSUBS 0.005793f
C714 B.n674 VSUBS 0.005793f
C715 B.n675 VSUBS 0.005793f
C716 B.n676 VSUBS 0.005793f
C717 B.n677 VSUBS 0.005793f
C718 B.n678 VSUBS 0.005793f
C719 B.n679 VSUBS 0.005793f
C720 B.n680 VSUBS 0.005793f
C721 B.n681 VSUBS 0.005793f
C722 B.n682 VSUBS 0.005793f
C723 B.n683 VSUBS 0.003237f
C724 B.n684 VSUBS 0.005793f
C725 B.n685 VSUBS 0.005793f
C726 B.n686 VSUBS 0.005793f
C727 B.n687 VSUBS 0.005793f
C728 B.n688 VSUBS 0.005793f
C729 B.n689 VSUBS 0.005793f
C730 B.n690 VSUBS 0.005793f
C731 B.n691 VSUBS 0.005793f
C732 B.n692 VSUBS 0.005793f
C733 B.n693 VSUBS 0.005793f
C734 B.n694 VSUBS 0.005793f
C735 B.n695 VSUBS 0.005793f
C736 B.n696 VSUBS 0.005793f
C737 B.n697 VSUBS 0.005793f
C738 B.n698 VSUBS 0.005793f
C739 B.n699 VSUBS 0.005793f
C740 B.n700 VSUBS 0.005793f
C741 B.n701 VSUBS 0.005793f
C742 B.n702 VSUBS 0.005793f
C743 B.n703 VSUBS 0.005793f
C744 B.n704 VSUBS 0.005793f
C745 B.n705 VSUBS 0.005793f
C746 B.n706 VSUBS 0.005793f
C747 B.n707 VSUBS 0.005793f
C748 B.n708 VSUBS 0.005793f
C749 B.n709 VSUBS 0.005793f
C750 B.n710 VSUBS 0.005793f
C751 B.n711 VSUBS 0.005793f
C752 B.n712 VSUBS 0.005793f
C753 B.n713 VSUBS 0.005793f
C754 B.n714 VSUBS 0.005793f
C755 B.n715 VSUBS 0.005793f
C756 B.n716 VSUBS 0.005793f
C757 B.n717 VSUBS 0.005793f
C758 B.n718 VSUBS 0.005793f
C759 B.n719 VSUBS 0.005793f
C760 B.n720 VSUBS 0.005793f
C761 B.n721 VSUBS 0.005793f
C762 B.n722 VSUBS 0.005793f
C763 B.n723 VSUBS 0.005793f
C764 B.n724 VSUBS 0.005793f
C765 B.n725 VSUBS 0.005793f
C766 B.n726 VSUBS 0.005793f
C767 B.n727 VSUBS 0.005793f
C768 B.n728 VSUBS 0.005793f
C769 B.n729 VSUBS 0.005793f
C770 B.n730 VSUBS 0.005793f
C771 B.n731 VSUBS 0.005793f
C772 B.n732 VSUBS 0.005793f
C773 B.n733 VSUBS 0.005793f
C774 B.n734 VSUBS 0.005793f
C775 B.n735 VSUBS 0.005793f
C776 B.n736 VSUBS 0.005793f
C777 B.n737 VSUBS 0.005793f
C778 B.n738 VSUBS 0.005793f
C779 B.n739 VSUBS 0.005793f
C780 B.n740 VSUBS 0.005793f
C781 B.n741 VSUBS 0.005793f
C782 B.n742 VSUBS 0.005793f
C783 B.n743 VSUBS 0.005793f
C784 B.n744 VSUBS 0.005793f
C785 B.n745 VSUBS 0.005793f
C786 B.n746 VSUBS 0.005793f
C787 B.n747 VSUBS 0.005793f
C788 B.n748 VSUBS 0.005793f
C789 B.n749 VSUBS 0.005793f
C790 B.n750 VSUBS 0.005793f
C791 B.n751 VSUBS 0.005793f
C792 B.n752 VSUBS 0.005793f
C793 B.n753 VSUBS 0.005793f
C794 B.n754 VSUBS 0.005793f
C795 B.n755 VSUBS 0.005793f
C796 B.n756 VSUBS 0.005793f
C797 B.n757 VSUBS 0.005793f
C798 B.n758 VSUBS 0.005793f
C799 B.n759 VSUBS 0.005793f
C800 B.n760 VSUBS 0.005793f
C801 B.n761 VSUBS 0.005793f
C802 B.n762 VSUBS 0.005793f
C803 B.n763 VSUBS 0.005793f
C804 B.n764 VSUBS 0.005793f
C805 B.n765 VSUBS 0.005793f
C806 B.n766 VSUBS 0.005793f
C807 B.n767 VSUBS 0.005793f
C808 B.n768 VSUBS 0.005793f
C809 B.n769 VSUBS 0.005793f
C810 B.n770 VSUBS 0.012748f
C811 B.n771 VSUBS 0.012748f
C812 B.n772 VSUBS 0.011957f
C813 B.n773 VSUBS 0.005793f
C814 B.n774 VSUBS 0.005793f
C815 B.n775 VSUBS 0.005793f
C816 B.n776 VSUBS 0.005793f
C817 B.n777 VSUBS 0.005793f
C818 B.n778 VSUBS 0.005793f
C819 B.n779 VSUBS 0.005793f
C820 B.n780 VSUBS 0.005793f
C821 B.n781 VSUBS 0.005793f
C822 B.n782 VSUBS 0.005793f
C823 B.n783 VSUBS 0.005793f
C824 B.n784 VSUBS 0.005793f
C825 B.n785 VSUBS 0.005793f
C826 B.n786 VSUBS 0.005793f
C827 B.n787 VSUBS 0.005793f
C828 B.n788 VSUBS 0.005793f
C829 B.n789 VSUBS 0.005793f
C830 B.n790 VSUBS 0.005793f
C831 B.n791 VSUBS 0.005793f
C832 B.n792 VSUBS 0.005793f
C833 B.n793 VSUBS 0.005793f
C834 B.n794 VSUBS 0.005793f
C835 B.n795 VSUBS 0.005793f
C836 B.n796 VSUBS 0.005793f
C837 B.n797 VSUBS 0.005793f
C838 B.n798 VSUBS 0.005793f
C839 B.n799 VSUBS 0.005793f
C840 B.n800 VSUBS 0.005793f
C841 B.n801 VSUBS 0.005793f
C842 B.n802 VSUBS 0.005793f
C843 B.n803 VSUBS 0.005793f
C844 B.n804 VSUBS 0.005793f
C845 B.n805 VSUBS 0.005793f
C846 B.n806 VSUBS 0.005793f
C847 B.n807 VSUBS 0.005793f
C848 B.n808 VSUBS 0.005793f
C849 B.n809 VSUBS 0.005793f
C850 B.n810 VSUBS 0.005793f
C851 B.n811 VSUBS 0.005793f
C852 B.n812 VSUBS 0.005793f
C853 B.n813 VSUBS 0.005793f
C854 B.n814 VSUBS 0.005793f
C855 B.n815 VSUBS 0.005793f
C856 B.n816 VSUBS 0.005793f
C857 B.n817 VSUBS 0.005793f
C858 B.n818 VSUBS 0.005793f
C859 B.n819 VSUBS 0.005793f
C860 B.n820 VSUBS 0.005793f
C861 B.n821 VSUBS 0.005793f
C862 B.n822 VSUBS 0.005793f
C863 B.n823 VSUBS 0.005793f
C864 B.n824 VSUBS 0.005793f
C865 B.n825 VSUBS 0.005793f
C866 B.n826 VSUBS 0.005793f
C867 B.n827 VSUBS 0.005793f
C868 B.n828 VSUBS 0.005793f
C869 B.n829 VSUBS 0.005793f
C870 B.n830 VSUBS 0.005793f
C871 B.n831 VSUBS 0.013117f
C872 VDD1.t1 VSUBS 0.373502f
C873 VDD1.t0 VSUBS 0.373502f
C874 VDD1.n0 VSUBS 3.09818f
C875 VDD1.t3 VSUBS 0.373502f
C876 VDD1.t2 VSUBS 0.373502f
C877 VDD1.n1 VSUBS 4.099f
C878 VP.t1 VSUBS 4.17016f
C879 VP.n0 VSUBS 1.54078f
C880 VP.n1 VSUBS 0.027406f
C881 VP.n2 VSUBS 0.022155f
C882 VP.n3 VSUBS 0.027406f
C883 VP.t0 VSUBS 4.17016f
C884 VP.n4 VSUBS 1.54078f
C885 VP.t2 VSUBS 4.5049f
C886 VP.t3 VSUBS 4.49464f
C887 VP.n5 VSUBS 4.65435f
C888 VP.n6 VSUBS 1.77291f
C889 VP.n7 VSUBS 0.044233f
C890 VP.n8 VSUBS 0.037965f
C891 VP.n9 VSUBS 0.051078f
C892 VP.n10 VSUBS 0.05447f
C893 VP.n11 VSUBS 0.027406f
C894 VP.n12 VSUBS 0.027406f
C895 VP.n13 VSUBS 0.027406f
C896 VP.n14 VSUBS 0.05447f
C897 VP.n15 VSUBS 0.051078f
C898 VP.n16 VSUBS 0.037965f
C899 VP.n17 VSUBS 0.044233f
C900 VP.n18 VSUBS 0.067512f
C901 VDD2.t1 VSUBS 0.36815f
C902 VDD2.t3 VSUBS 0.36815f
C903 VDD2.n0 VSUBS 4.0128f
C904 VDD2.t0 VSUBS 0.36815f
C905 VDD2.t2 VSUBS 0.36815f
C906 VDD2.n1 VSUBS 3.05312f
C907 VDD2.n2 VSUBS 4.99945f
C908 VTAIL.n0 VSUBS 0.024932f
C909 VTAIL.n1 VSUBS 0.022689f
C910 VTAIL.n2 VSUBS 0.012192f
C911 VTAIL.n3 VSUBS 0.028818f
C912 VTAIL.n4 VSUBS 0.012909f
C913 VTAIL.n5 VSUBS 0.022689f
C914 VTAIL.n6 VSUBS 0.012192f
C915 VTAIL.n7 VSUBS 0.028818f
C916 VTAIL.n8 VSUBS 0.012551f
C917 VTAIL.n9 VSUBS 0.022689f
C918 VTAIL.n10 VSUBS 0.012909f
C919 VTAIL.n11 VSUBS 0.028818f
C920 VTAIL.n12 VSUBS 0.012909f
C921 VTAIL.n13 VSUBS 0.022689f
C922 VTAIL.n14 VSUBS 0.012192f
C923 VTAIL.n15 VSUBS 0.028818f
C924 VTAIL.n16 VSUBS 0.012909f
C925 VTAIL.n17 VSUBS 0.022689f
C926 VTAIL.n18 VSUBS 0.012192f
C927 VTAIL.n19 VSUBS 0.028818f
C928 VTAIL.n20 VSUBS 0.012909f
C929 VTAIL.n21 VSUBS 0.022689f
C930 VTAIL.n22 VSUBS 0.012192f
C931 VTAIL.n23 VSUBS 0.028818f
C932 VTAIL.n24 VSUBS 0.012909f
C933 VTAIL.n25 VSUBS 0.022689f
C934 VTAIL.n26 VSUBS 0.012192f
C935 VTAIL.n27 VSUBS 0.028818f
C936 VTAIL.n28 VSUBS 0.012909f
C937 VTAIL.n29 VSUBS 1.71346f
C938 VTAIL.n30 VSUBS 0.012192f
C939 VTAIL.t4 VSUBS 0.061838f
C940 VTAIL.n31 VSUBS 0.177138f
C941 VTAIL.n32 VSUBS 0.018333f
C942 VTAIL.n33 VSUBS 0.021613f
C943 VTAIL.n34 VSUBS 0.028818f
C944 VTAIL.n35 VSUBS 0.012909f
C945 VTAIL.n36 VSUBS 0.012192f
C946 VTAIL.n37 VSUBS 0.022689f
C947 VTAIL.n38 VSUBS 0.022689f
C948 VTAIL.n39 VSUBS 0.012192f
C949 VTAIL.n40 VSUBS 0.012909f
C950 VTAIL.n41 VSUBS 0.028818f
C951 VTAIL.n42 VSUBS 0.028818f
C952 VTAIL.n43 VSUBS 0.012909f
C953 VTAIL.n44 VSUBS 0.012192f
C954 VTAIL.n45 VSUBS 0.022689f
C955 VTAIL.n46 VSUBS 0.022689f
C956 VTAIL.n47 VSUBS 0.012192f
C957 VTAIL.n48 VSUBS 0.012909f
C958 VTAIL.n49 VSUBS 0.028818f
C959 VTAIL.n50 VSUBS 0.028818f
C960 VTAIL.n51 VSUBS 0.012909f
C961 VTAIL.n52 VSUBS 0.012192f
C962 VTAIL.n53 VSUBS 0.022689f
C963 VTAIL.n54 VSUBS 0.022689f
C964 VTAIL.n55 VSUBS 0.012192f
C965 VTAIL.n56 VSUBS 0.012909f
C966 VTAIL.n57 VSUBS 0.028818f
C967 VTAIL.n58 VSUBS 0.028818f
C968 VTAIL.n59 VSUBS 0.012909f
C969 VTAIL.n60 VSUBS 0.012192f
C970 VTAIL.n61 VSUBS 0.022689f
C971 VTAIL.n62 VSUBS 0.022689f
C972 VTAIL.n63 VSUBS 0.012192f
C973 VTAIL.n64 VSUBS 0.012909f
C974 VTAIL.n65 VSUBS 0.028818f
C975 VTAIL.n66 VSUBS 0.028818f
C976 VTAIL.n67 VSUBS 0.012909f
C977 VTAIL.n68 VSUBS 0.012192f
C978 VTAIL.n69 VSUBS 0.022689f
C979 VTAIL.n70 VSUBS 0.022689f
C980 VTAIL.n71 VSUBS 0.012192f
C981 VTAIL.n72 VSUBS 0.012192f
C982 VTAIL.n73 VSUBS 0.012909f
C983 VTAIL.n74 VSUBS 0.028818f
C984 VTAIL.n75 VSUBS 0.028818f
C985 VTAIL.n76 VSUBS 0.028818f
C986 VTAIL.n77 VSUBS 0.012551f
C987 VTAIL.n78 VSUBS 0.012192f
C988 VTAIL.n79 VSUBS 0.022689f
C989 VTAIL.n80 VSUBS 0.022689f
C990 VTAIL.n81 VSUBS 0.012192f
C991 VTAIL.n82 VSUBS 0.012909f
C992 VTAIL.n83 VSUBS 0.028818f
C993 VTAIL.n84 VSUBS 0.028818f
C994 VTAIL.n85 VSUBS 0.012909f
C995 VTAIL.n86 VSUBS 0.012192f
C996 VTAIL.n87 VSUBS 0.022689f
C997 VTAIL.n88 VSUBS 0.022689f
C998 VTAIL.n89 VSUBS 0.012192f
C999 VTAIL.n90 VSUBS 0.012909f
C1000 VTAIL.n91 VSUBS 0.028818f
C1001 VTAIL.n92 VSUBS 0.069769f
C1002 VTAIL.n93 VSUBS 0.012909f
C1003 VTAIL.n94 VSUBS 0.012192f
C1004 VTAIL.n95 VSUBS 0.053995f
C1005 VTAIL.n96 VSUBS 0.035134f
C1006 VTAIL.n97 VSUBS 0.168521f
C1007 VTAIL.n98 VSUBS 0.024932f
C1008 VTAIL.n99 VSUBS 0.022689f
C1009 VTAIL.n100 VSUBS 0.012192f
C1010 VTAIL.n101 VSUBS 0.028818f
C1011 VTAIL.n102 VSUBS 0.012909f
C1012 VTAIL.n103 VSUBS 0.022689f
C1013 VTAIL.n104 VSUBS 0.012192f
C1014 VTAIL.n105 VSUBS 0.028818f
C1015 VTAIL.n106 VSUBS 0.012551f
C1016 VTAIL.n107 VSUBS 0.022689f
C1017 VTAIL.n108 VSUBS 0.012909f
C1018 VTAIL.n109 VSUBS 0.028818f
C1019 VTAIL.n110 VSUBS 0.012909f
C1020 VTAIL.n111 VSUBS 0.022689f
C1021 VTAIL.n112 VSUBS 0.012192f
C1022 VTAIL.n113 VSUBS 0.028818f
C1023 VTAIL.n114 VSUBS 0.012909f
C1024 VTAIL.n115 VSUBS 0.022689f
C1025 VTAIL.n116 VSUBS 0.012192f
C1026 VTAIL.n117 VSUBS 0.028818f
C1027 VTAIL.n118 VSUBS 0.012909f
C1028 VTAIL.n119 VSUBS 0.022689f
C1029 VTAIL.n120 VSUBS 0.012192f
C1030 VTAIL.n121 VSUBS 0.028818f
C1031 VTAIL.n122 VSUBS 0.012909f
C1032 VTAIL.n123 VSUBS 0.022689f
C1033 VTAIL.n124 VSUBS 0.012192f
C1034 VTAIL.n125 VSUBS 0.028818f
C1035 VTAIL.n126 VSUBS 0.012909f
C1036 VTAIL.n127 VSUBS 1.71346f
C1037 VTAIL.n128 VSUBS 0.012192f
C1038 VTAIL.t3 VSUBS 0.061838f
C1039 VTAIL.n129 VSUBS 0.177138f
C1040 VTAIL.n130 VSUBS 0.018333f
C1041 VTAIL.n131 VSUBS 0.021613f
C1042 VTAIL.n132 VSUBS 0.028818f
C1043 VTAIL.n133 VSUBS 0.012909f
C1044 VTAIL.n134 VSUBS 0.012192f
C1045 VTAIL.n135 VSUBS 0.022689f
C1046 VTAIL.n136 VSUBS 0.022689f
C1047 VTAIL.n137 VSUBS 0.012192f
C1048 VTAIL.n138 VSUBS 0.012909f
C1049 VTAIL.n139 VSUBS 0.028818f
C1050 VTAIL.n140 VSUBS 0.028818f
C1051 VTAIL.n141 VSUBS 0.012909f
C1052 VTAIL.n142 VSUBS 0.012192f
C1053 VTAIL.n143 VSUBS 0.022689f
C1054 VTAIL.n144 VSUBS 0.022689f
C1055 VTAIL.n145 VSUBS 0.012192f
C1056 VTAIL.n146 VSUBS 0.012909f
C1057 VTAIL.n147 VSUBS 0.028818f
C1058 VTAIL.n148 VSUBS 0.028818f
C1059 VTAIL.n149 VSUBS 0.012909f
C1060 VTAIL.n150 VSUBS 0.012192f
C1061 VTAIL.n151 VSUBS 0.022689f
C1062 VTAIL.n152 VSUBS 0.022689f
C1063 VTAIL.n153 VSUBS 0.012192f
C1064 VTAIL.n154 VSUBS 0.012909f
C1065 VTAIL.n155 VSUBS 0.028818f
C1066 VTAIL.n156 VSUBS 0.028818f
C1067 VTAIL.n157 VSUBS 0.012909f
C1068 VTAIL.n158 VSUBS 0.012192f
C1069 VTAIL.n159 VSUBS 0.022689f
C1070 VTAIL.n160 VSUBS 0.022689f
C1071 VTAIL.n161 VSUBS 0.012192f
C1072 VTAIL.n162 VSUBS 0.012909f
C1073 VTAIL.n163 VSUBS 0.028818f
C1074 VTAIL.n164 VSUBS 0.028818f
C1075 VTAIL.n165 VSUBS 0.012909f
C1076 VTAIL.n166 VSUBS 0.012192f
C1077 VTAIL.n167 VSUBS 0.022689f
C1078 VTAIL.n168 VSUBS 0.022689f
C1079 VTAIL.n169 VSUBS 0.012192f
C1080 VTAIL.n170 VSUBS 0.012192f
C1081 VTAIL.n171 VSUBS 0.012909f
C1082 VTAIL.n172 VSUBS 0.028818f
C1083 VTAIL.n173 VSUBS 0.028818f
C1084 VTAIL.n174 VSUBS 0.028818f
C1085 VTAIL.n175 VSUBS 0.012551f
C1086 VTAIL.n176 VSUBS 0.012192f
C1087 VTAIL.n177 VSUBS 0.022689f
C1088 VTAIL.n178 VSUBS 0.022689f
C1089 VTAIL.n179 VSUBS 0.012192f
C1090 VTAIL.n180 VSUBS 0.012909f
C1091 VTAIL.n181 VSUBS 0.028818f
C1092 VTAIL.n182 VSUBS 0.028818f
C1093 VTAIL.n183 VSUBS 0.012909f
C1094 VTAIL.n184 VSUBS 0.012192f
C1095 VTAIL.n185 VSUBS 0.022689f
C1096 VTAIL.n186 VSUBS 0.022689f
C1097 VTAIL.n187 VSUBS 0.012192f
C1098 VTAIL.n188 VSUBS 0.012909f
C1099 VTAIL.n189 VSUBS 0.028818f
C1100 VTAIL.n190 VSUBS 0.069769f
C1101 VTAIL.n191 VSUBS 0.012909f
C1102 VTAIL.n192 VSUBS 0.012192f
C1103 VTAIL.n193 VSUBS 0.053995f
C1104 VTAIL.n194 VSUBS 0.035134f
C1105 VTAIL.n195 VSUBS 0.273931f
C1106 VTAIL.n196 VSUBS 0.024932f
C1107 VTAIL.n197 VSUBS 0.022689f
C1108 VTAIL.n198 VSUBS 0.012192f
C1109 VTAIL.n199 VSUBS 0.028818f
C1110 VTAIL.n200 VSUBS 0.012909f
C1111 VTAIL.n201 VSUBS 0.022689f
C1112 VTAIL.n202 VSUBS 0.012192f
C1113 VTAIL.n203 VSUBS 0.028818f
C1114 VTAIL.n204 VSUBS 0.012551f
C1115 VTAIL.n205 VSUBS 0.022689f
C1116 VTAIL.n206 VSUBS 0.012909f
C1117 VTAIL.n207 VSUBS 0.028818f
C1118 VTAIL.n208 VSUBS 0.012909f
C1119 VTAIL.n209 VSUBS 0.022689f
C1120 VTAIL.n210 VSUBS 0.012192f
C1121 VTAIL.n211 VSUBS 0.028818f
C1122 VTAIL.n212 VSUBS 0.012909f
C1123 VTAIL.n213 VSUBS 0.022689f
C1124 VTAIL.n214 VSUBS 0.012192f
C1125 VTAIL.n215 VSUBS 0.028818f
C1126 VTAIL.n216 VSUBS 0.012909f
C1127 VTAIL.n217 VSUBS 0.022689f
C1128 VTAIL.n218 VSUBS 0.012192f
C1129 VTAIL.n219 VSUBS 0.028818f
C1130 VTAIL.n220 VSUBS 0.012909f
C1131 VTAIL.n221 VSUBS 0.022689f
C1132 VTAIL.n222 VSUBS 0.012192f
C1133 VTAIL.n223 VSUBS 0.028818f
C1134 VTAIL.n224 VSUBS 0.012909f
C1135 VTAIL.n225 VSUBS 1.71346f
C1136 VTAIL.n226 VSUBS 0.012192f
C1137 VTAIL.t1 VSUBS 0.061838f
C1138 VTAIL.n227 VSUBS 0.177138f
C1139 VTAIL.n228 VSUBS 0.018333f
C1140 VTAIL.n229 VSUBS 0.021613f
C1141 VTAIL.n230 VSUBS 0.028818f
C1142 VTAIL.n231 VSUBS 0.012909f
C1143 VTAIL.n232 VSUBS 0.012192f
C1144 VTAIL.n233 VSUBS 0.022689f
C1145 VTAIL.n234 VSUBS 0.022689f
C1146 VTAIL.n235 VSUBS 0.012192f
C1147 VTAIL.n236 VSUBS 0.012909f
C1148 VTAIL.n237 VSUBS 0.028818f
C1149 VTAIL.n238 VSUBS 0.028818f
C1150 VTAIL.n239 VSUBS 0.012909f
C1151 VTAIL.n240 VSUBS 0.012192f
C1152 VTAIL.n241 VSUBS 0.022689f
C1153 VTAIL.n242 VSUBS 0.022689f
C1154 VTAIL.n243 VSUBS 0.012192f
C1155 VTAIL.n244 VSUBS 0.012909f
C1156 VTAIL.n245 VSUBS 0.028818f
C1157 VTAIL.n246 VSUBS 0.028818f
C1158 VTAIL.n247 VSUBS 0.012909f
C1159 VTAIL.n248 VSUBS 0.012192f
C1160 VTAIL.n249 VSUBS 0.022689f
C1161 VTAIL.n250 VSUBS 0.022689f
C1162 VTAIL.n251 VSUBS 0.012192f
C1163 VTAIL.n252 VSUBS 0.012909f
C1164 VTAIL.n253 VSUBS 0.028818f
C1165 VTAIL.n254 VSUBS 0.028818f
C1166 VTAIL.n255 VSUBS 0.012909f
C1167 VTAIL.n256 VSUBS 0.012192f
C1168 VTAIL.n257 VSUBS 0.022689f
C1169 VTAIL.n258 VSUBS 0.022689f
C1170 VTAIL.n259 VSUBS 0.012192f
C1171 VTAIL.n260 VSUBS 0.012909f
C1172 VTAIL.n261 VSUBS 0.028818f
C1173 VTAIL.n262 VSUBS 0.028818f
C1174 VTAIL.n263 VSUBS 0.012909f
C1175 VTAIL.n264 VSUBS 0.012192f
C1176 VTAIL.n265 VSUBS 0.022689f
C1177 VTAIL.n266 VSUBS 0.022689f
C1178 VTAIL.n267 VSUBS 0.012192f
C1179 VTAIL.n268 VSUBS 0.012192f
C1180 VTAIL.n269 VSUBS 0.012909f
C1181 VTAIL.n270 VSUBS 0.028818f
C1182 VTAIL.n271 VSUBS 0.028818f
C1183 VTAIL.n272 VSUBS 0.028818f
C1184 VTAIL.n273 VSUBS 0.012551f
C1185 VTAIL.n274 VSUBS 0.012192f
C1186 VTAIL.n275 VSUBS 0.022689f
C1187 VTAIL.n276 VSUBS 0.022689f
C1188 VTAIL.n277 VSUBS 0.012192f
C1189 VTAIL.n278 VSUBS 0.012909f
C1190 VTAIL.n279 VSUBS 0.028818f
C1191 VTAIL.n280 VSUBS 0.028818f
C1192 VTAIL.n281 VSUBS 0.012909f
C1193 VTAIL.n282 VSUBS 0.012192f
C1194 VTAIL.n283 VSUBS 0.022689f
C1195 VTAIL.n284 VSUBS 0.022689f
C1196 VTAIL.n285 VSUBS 0.012192f
C1197 VTAIL.n286 VSUBS 0.012909f
C1198 VTAIL.n287 VSUBS 0.028818f
C1199 VTAIL.n288 VSUBS 0.069769f
C1200 VTAIL.n289 VSUBS 0.012909f
C1201 VTAIL.n290 VSUBS 0.012192f
C1202 VTAIL.n291 VSUBS 0.053995f
C1203 VTAIL.n292 VSUBS 0.035134f
C1204 VTAIL.n293 VSUBS 1.87447f
C1205 VTAIL.n294 VSUBS 0.024932f
C1206 VTAIL.n295 VSUBS 0.022689f
C1207 VTAIL.n296 VSUBS 0.012192f
C1208 VTAIL.n297 VSUBS 0.028818f
C1209 VTAIL.n298 VSUBS 0.012909f
C1210 VTAIL.n299 VSUBS 0.022689f
C1211 VTAIL.n300 VSUBS 0.012192f
C1212 VTAIL.n301 VSUBS 0.028818f
C1213 VTAIL.n302 VSUBS 0.012551f
C1214 VTAIL.n303 VSUBS 0.022689f
C1215 VTAIL.n304 VSUBS 0.012551f
C1216 VTAIL.n305 VSUBS 0.012192f
C1217 VTAIL.n306 VSUBS 0.028818f
C1218 VTAIL.n307 VSUBS 0.028818f
C1219 VTAIL.n308 VSUBS 0.012909f
C1220 VTAIL.n309 VSUBS 0.022689f
C1221 VTAIL.n310 VSUBS 0.012192f
C1222 VTAIL.n311 VSUBS 0.028818f
C1223 VTAIL.n312 VSUBS 0.012909f
C1224 VTAIL.n313 VSUBS 0.022689f
C1225 VTAIL.n314 VSUBS 0.012192f
C1226 VTAIL.n315 VSUBS 0.028818f
C1227 VTAIL.n316 VSUBS 0.012909f
C1228 VTAIL.n317 VSUBS 0.022689f
C1229 VTAIL.n318 VSUBS 0.012192f
C1230 VTAIL.n319 VSUBS 0.028818f
C1231 VTAIL.n320 VSUBS 0.012909f
C1232 VTAIL.n321 VSUBS 0.022689f
C1233 VTAIL.n322 VSUBS 0.012192f
C1234 VTAIL.n323 VSUBS 0.028818f
C1235 VTAIL.n324 VSUBS 0.012909f
C1236 VTAIL.n325 VSUBS 1.71346f
C1237 VTAIL.n326 VSUBS 0.012192f
C1238 VTAIL.t6 VSUBS 0.061838f
C1239 VTAIL.n327 VSUBS 0.177138f
C1240 VTAIL.n328 VSUBS 0.018333f
C1241 VTAIL.n329 VSUBS 0.021613f
C1242 VTAIL.n330 VSUBS 0.028818f
C1243 VTAIL.n331 VSUBS 0.012909f
C1244 VTAIL.n332 VSUBS 0.012192f
C1245 VTAIL.n333 VSUBS 0.022689f
C1246 VTAIL.n334 VSUBS 0.022689f
C1247 VTAIL.n335 VSUBS 0.012192f
C1248 VTAIL.n336 VSUBS 0.012909f
C1249 VTAIL.n337 VSUBS 0.028818f
C1250 VTAIL.n338 VSUBS 0.028818f
C1251 VTAIL.n339 VSUBS 0.012909f
C1252 VTAIL.n340 VSUBS 0.012192f
C1253 VTAIL.n341 VSUBS 0.022689f
C1254 VTAIL.n342 VSUBS 0.022689f
C1255 VTAIL.n343 VSUBS 0.012192f
C1256 VTAIL.n344 VSUBS 0.012909f
C1257 VTAIL.n345 VSUBS 0.028818f
C1258 VTAIL.n346 VSUBS 0.028818f
C1259 VTAIL.n347 VSUBS 0.012909f
C1260 VTAIL.n348 VSUBS 0.012192f
C1261 VTAIL.n349 VSUBS 0.022689f
C1262 VTAIL.n350 VSUBS 0.022689f
C1263 VTAIL.n351 VSUBS 0.012192f
C1264 VTAIL.n352 VSUBS 0.012909f
C1265 VTAIL.n353 VSUBS 0.028818f
C1266 VTAIL.n354 VSUBS 0.028818f
C1267 VTAIL.n355 VSUBS 0.012909f
C1268 VTAIL.n356 VSUBS 0.012192f
C1269 VTAIL.n357 VSUBS 0.022689f
C1270 VTAIL.n358 VSUBS 0.022689f
C1271 VTAIL.n359 VSUBS 0.012192f
C1272 VTAIL.n360 VSUBS 0.012909f
C1273 VTAIL.n361 VSUBS 0.028818f
C1274 VTAIL.n362 VSUBS 0.028818f
C1275 VTAIL.n363 VSUBS 0.012909f
C1276 VTAIL.n364 VSUBS 0.012192f
C1277 VTAIL.n365 VSUBS 0.022689f
C1278 VTAIL.n366 VSUBS 0.022689f
C1279 VTAIL.n367 VSUBS 0.012192f
C1280 VTAIL.n368 VSUBS 0.012909f
C1281 VTAIL.n369 VSUBS 0.028818f
C1282 VTAIL.n370 VSUBS 0.028818f
C1283 VTAIL.n371 VSUBS 0.012909f
C1284 VTAIL.n372 VSUBS 0.012192f
C1285 VTAIL.n373 VSUBS 0.022689f
C1286 VTAIL.n374 VSUBS 0.022689f
C1287 VTAIL.n375 VSUBS 0.012192f
C1288 VTAIL.n376 VSUBS 0.012909f
C1289 VTAIL.n377 VSUBS 0.028818f
C1290 VTAIL.n378 VSUBS 0.028818f
C1291 VTAIL.n379 VSUBS 0.012909f
C1292 VTAIL.n380 VSUBS 0.012192f
C1293 VTAIL.n381 VSUBS 0.022689f
C1294 VTAIL.n382 VSUBS 0.022689f
C1295 VTAIL.n383 VSUBS 0.012192f
C1296 VTAIL.n384 VSUBS 0.012909f
C1297 VTAIL.n385 VSUBS 0.028818f
C1298 VTAIL.n386 VSUBS 0.069769f
C1299 VTAIL.n387 VSUBS 0.012909f
C1300 VTAIL.n388 VSUBS 0.012192f
C1301 VTAIL.n389 VSUBS 0.053995f
C1302 VTAIL.n390 VSUBS 0.035134f
C1303 VTAIL.n391 VSUBS 1.87447f
C1304 VTAIL.n392 VSUBS 0.024932f
C1305 VTAIL.n393 VSUBS 0.022689f
C1306 VTAIL.n394 VSUBS 0.012192f
C1307 VTAIL.n395 VSUBS 0.028818f
C1308 VTAIL.n396 VSUBS 0.012909f
C1309 VTAIL.n397 VSUBS 0.022689f
C1310 VTAIL.n398 VSUBS 0.012192f
C1311 VTAIL.n399 VSUBS 0.028818f
C1312 VTAIL.n400 VSUBS 0.012551f
C1313 VTAIL.n401 VSUBS 0.022689f
C1314 VTAIL.n402 VSUBS 0.012551f
C1315 VTAIL.n403 VSUBS 0.012192f
C1316 VTAIL.n404 VSUBS 0.028818f
C1317 VTAIL.n405 VSUBS 0.028818f
C1318 VTAIL.n406 VSUBS 0.012909f
C1319 VTAIL.n407 VSUBS 0.022689f
C1320 VTAIL.n408 VSUBS 0.012192f
C1321 VTAIL.n409 VSUBS 0.028818f
C1322 VTAIL.n410 VSUBS 0.012909f
C1323 VTAIL.n411 VSUBS 0.022689f
C1324 VTAIL.n412 VSUBS 0.012192f
C1325 VTAIL.n413 VSUBS 0.028818f
C1326 VTAIL.n414 VSUBS 0.012909f
C1327 VTAIL.n415 VSUBS 0.022689f
C1328 VTAIL.n416 VSUBS 0.012192f
C1329 VTAIL.n417 VSUBS 0.028818f
C1330 VTAIL.n418 VSUBS 0.012909f
C1331 VTAIL.n419 VSUBS 0.022689f
C1332 VTAIL.n420 VSUBS 0.012192f
C1333 VTAIL.n421 VSUBS 0.028818f
C1334 VTAIL.n422 VSUBS 0.012909f
C1335 VTAIL.n423 VSUBS 1.71346f
C1336 VTAIL.n424 VSUBS 0.012192f
C1337 VTAIL.t5 VSUBS 0.061838f
C1338 VTAIL.n425 VSUBS 0.177138f
C1339 VTAIL.n426 VSUBS 0.018333f
C1340 VTAIL.n427 VSUBS 0.021613f
C1341 VTAIL.n428 VSUBS 0.028818f
C1342 VTAIL.n429 VSUBS 0.012909f
C1343 VTAIL.n430 VSUBS 0.012192f
C1344 VTAIL.n431 VSUBS 0.022689f
C1345 VTAIL.n432 VSUBS 0.022689f
C1346 VTAIL.n433 VSUBS 0.012192f
C1347 VTAIL.n434 VSUBS 0.012909f
C1348 VTAIL.n435 VSUBS 0.028818f
C1349 VTAIL.n436 VSUBS 0.028818f
C1350 VTAIL.n437 VSUBS 0.012909f
C1351 VTAIL.n438 VSUBS 0.012192f
C1352 VTAIL.n439 VSUBS 0.022689f
C1353 VTAIL.n440 VSUBS 0.022689f
C1354 VTAIL.n441 VSUBS 0.012192f
C1355 VTAIL.n442 VSUBS 0.012909f
C1356 VTAIL.n443 VSUBS 0.028818f
C1357 VTAIL.n444 VSUBS 0.028818f
C1358 VTAIL.n445 VSUBS 0.012909f
C1359 VTAIL.n446 VSUBS 0.012192f
C1360 VTAIL.n447 VSUBS 0.022689f
C1361 VTAIL.n448 VSUBS 0.022689f
C1362 VTAIL.n449 VSUBS 0.012192f
C1363 VTAIL.n450 VSUBS 0.012909f
C1364 VTAIL.n451 VSUBS 0.028818f
C1365 VTAIL.n452 VSUBS 0.028818f
C1366 VTAIL.n453 VSUBS 0.012909f
C1367 VTAIL.n454 VSUBS 0.012192f
C1368 VTAIL.n455 VSUBS 0.022689f
C1369 VTAIL.n456 VSUBS 0.022689f
C1370 VTAIL.n457 VSUBS 0.012192f
C1371 VTAIL.n458 VSUBS 0.012909f
C1372 VTAIL.n459 VSUBS 0.028818f
C1373 VTAIL.n460 VSUBS 0.028818f
C1374 VTAIL.n461 VSUBS 0.012909f
C1375 VTAIL.n462 VSUBS 0.012192f
C1376 VTAIL.n463 VSUBS 0.022689f
C1377 VTAIL.n464 VSUBS 0.022689f
C1378 VTAIL.n465 VSUBS 0.012192f
C1379 VTAIL.n466 VSUBS 0.012909f
C1380 VTAIL.n467 VSUBS 0.028818f
C1381 VTAIL.n468 VSUBS 0.028818f
C1382 VTAIL.n469 VSUBS 0.012909f
C1383 VTAIL.n470 VSUBS 0.012192f
C1384 VTAIL.n471 VSUBS 0.022689f
C1385 VTAIL.n472 VSUBS 0.022689f
C1386 VTAIL.n473 VSUBS 0.012192f
C1387 VTAIL.n474 VSUBS 0.012909f
C1388 VTAIL.n475 VSUBS 0.028818f
C1389 VTAIL.n476 VSUBS 0.028818f
C1390 VTAIL.n477 VSUBS 0.012909f
C1391 VTAIL.n478 VSUBS 0.012192f
C1392 VTAIL.n479 VSUBS 0.022689f
C1393 VTAIL.n480 VSUBS 0.022689f
C1394 VTAIL.n481 VSUBS 0.012192f
C1395 VTAIL.n482 VSUBS 0.012909f
C1396 VTAIL.n483 VSUBS 0.028818f
C1397 VTAIL.n484 VSUBS 0.069769f
C1398 VTAIL.n485 VSUBS 0.012909f
C1399 VTAIL.n486 VSUBS 0.012192f
C1400 VTAIL.n487 VSUBS 0.053995f
C1401 VTAIL.n488 VSUBS 0.035134f
C1402 VTAIL.n489 VSUBS 0.273931f
C1403 VTAIL.n490 VSUBS 0.024932f
C1404 VTAIL.n491 VSUBS 0.022689f
C1405 VTAIL.n492 VSUBS 0.012192f
C1406 VTAIL.n493 VSUBS 0.028818f
C1407 VTAIL.n494 VSUBS 0.012909f
C1408 VTAIL.n495 VSUBS 0.022689f
C1409 VTAIL.n496 VSUBS 0.012192f
C1410 VTAIL.n497 VSUBS 0.028818f
C1411 VTAIL.n498 VSUBS 0.012551f
C1412 VTAIL.n499 VSUBS 0.022689f
C1413 VTAIL.n500 VSUBS 0.012551f
C1414 VTAIL.n501 VSUBS 0.012192f
C1415 VTAIL.n502 VSUBS 0.028818f
C1416 VTAIL.n503 VSUBS 0.028818f
C1417 VTAIL.n504 VSUBS 0.012909f
C1418 VTAIL.n505 VSUBS 0.022689f
C1419 VTAIL.n506 VSUBS 0.012192f
C1420 VTAIL.n507 VSUBS 0.028818f
C1421 VTAIL.n508 VSUBS 0.012909f
C1422 VTAIL.n509 VSUBS 0.022689f
C1423 VTAIL.n510 VSUBS 0.012192f
C1424 VTAIL.n511 VSUBS 0.028818f
C1425 VTAIL.n512 VSUBS 0.012909f
C1426 VTAIL.n513 VSUBS 0.022689f
C1427 VTAIL.n514 VSUBS 0.012192f
C1428 VTAIL.n515 VSUBS 0.028818f
C1429 VTAIL.n516 VSUBS 0.012909f
C1430 VTAIL.n517 VSUBS 0.022689f
C1431 VTAIL.n518 VSUBS 0.012192f
C1432 VTAIL.n519 VSUBS 0.028818f
C1433 VTAIL.n520 VSUBS 0.012909f
C1434 VTAIL.n521 VSUBS 1.71346f
C1435 VTAIL.n522 VSUBS 0.012192f
C1436 VTAIL.t0 VSUBS 0.061838f
C1437 VTAIL.n523 VSUBS 0.177138f
C1438 VTAIL.n524 VSUBS 0.018333f
C1439 VTAIL.n525 VSUBS 0.021613f
C1440 VTAIL.n526 VSUBS 0.028818f
C1441 VTAIL.n527 VSUBS 0.012909f
C1442 VTAIL.n528 VSUBS 0.012192f
C1443 VTAIL.n529 VSUBS 0.022689f
C1444 VTAIL.n530 VSUBS 0.022689f
C1445 VTAIL.n531 VSUBS 0.012192f
C1446 VTAIL.n532 VSUBS 0.012909f
C1447 VTAIL.n533 VSUBS 0.028818f
C1448 VTAIL.n534 VSUBS 0.028818f
C1449 VTAIL.n535 VSUBS 0.012909f
C1450 VTAIL.n536 VSUBS 0.012192f
C1451 VTAIL.n537 VSUBS 0.022689f
C1452 VTAIL.n538 VSUBS 0.022689f
C1453 VTAIL.n539 VSUBS 0.012192f
C1454 VTAIL.n540 VSUBS 0.012909f
C1455 VTAIL.n541 VSUBS 0.028818f
C1456 VTAIL.n542 VSUBS 0.028818f
C1457 VTAIL.n543 VSUBS 0.012909f
C1458 VTAIL.n544 VSUBS 0.012192f
C1459 VTAIL.n545 VSUBS 0.022689f
C1460 VTAIL.n546 VSUBS 0.022689f
C1461 VTAIL.n547 VSUBS 0.012192f
C1462 VTAIL.n548 VSUBS 0.012909f
C1463 VTAIL.n549 VSUBS 0.028818f
C1464 VTAIL.n550 VSUBS 0.028818f
C1465 VTAIL.n551 VSUBS 0.012909f
C1466 VTAIL.n552 VSUBS 0.012192f
C1467 VTAIL.n553 VSUBS 0.022689f
C1468 VTAIL.n554 VSUBS 0.022689f
C1469 VTAIL.n555 VSUBS 0.012192f
C1470 VTAIL.n556 VSUBS 0.012909f
C1471 VTAIL.n557 VSUBS 0.028818f
C1472 VTAIL.n558 VSUBS 0.028818f
C1473 VTAIL.n559 VSUBS 0.012909f
C1474 VTAIL.n560 VSUBS 0.012192f
C1475 VTAIL.n561 VSUBS 0.022689f
C1476 VTAIL.n562 VSUBS 0.022689f
C1477 VTAIL.n563 VSUBS 0.012192f
C1478 VTAIL.n564 VSUBS 0.012909f
C1479 VTAIL.n565 VSUBS 0.028818f
C1480 VTAIL.n566 VSUBS 0.028818f
C1481 VTAIL.n567 VSUBS 0.012909f
C1482 VTAIL.n568 VSUBS 0.012192f
C1483 VTAIL.n569 VSUBS 0.022689f
C1484 VTAIL.n570 VSUBS 0.022689f
C1485 VTAIL.n571 VSUBS 0.012192f
C1486 VTAIL.n572 VSUBS 0.012909f
C1487 VTAIL.n573 VSUBS 0.028818f
C1488 VTAIL.n574 VSUBS 0.028818f
C1489 VTAIL.n575 VSUBS 0.012909f
C1490 VTAIL.n576 VSUBS 0.012192f
C1491 VTAIL.n577 VSUBS 0.022689f
C1492 VTAIL.n578 VSUBS 0.022689f
C1493 VTAIL.n579 VSUBS 0.012192f
C1494 VTAIL.n580 VSUBS 0.012909f
C1495 VTAIL.n581 VSUBS 0.028818f
C1496 VTAIL.n582 VSUBS 0.069769f
C1497 VTAIL.n583 VSUBS 0.012909f
C1498 VTAIL.n584 VSUBS 0.012192f
C1499 VTAIL.n585 VSUBS 0.053995f
C1500 VTAIL.n586 VSUBS 0.035134f
C1501 VTAIL.n587 VSUBS 0.273931f
C1502 VTAIL.n588 VSUBS 0.024932f
C1503 VTAIL.n589 VSUBS 0.022689f
C1504 VTAIL.n590 VSUBS 0.012192f
C1505 VTAIL.n591 VSUBS 0.028818f
C1506 VTAIL.n592 VSUBS 0.012909f
C1507 VTAIL.n593 VSUBS 0.022689f
C1508 VTAIL.n594 VSUBS 0.012192f
C1509 VTAIL.n595 VSUBS 0.028818f
C1510 VTAIL.n596 VSUBS 0.012551f
C1511 VTAIL.n597 VSUBS 0.022689f
C1512 VTAIL.n598 VSUBS 0.012551f
C1513 VTAIL.n599 VSUBS 0.012192f
C1514 VTAIL.n600 VSUBS 0.028818f
C1515 VTAIL.n601 VSUBS 0.028818f
C1516 VTAIL.n602 VSUBS 0.012909f
C1517 VTAIL.n603 VSUBS 0.022689f
C1518 VTAIL.n604 VSUBS 0.012192f
C1519 VTAIL.n605 VSUBS 0.028818f
C1520 VTAIL.n606 VSUBS 0.012909f
C1521 VTAIL.n607 VSUBS 0.022689f
C1522 VTAIL.n608 VSUBS 0.012192f
C1523 VTAIL.n609 VSUBS 0.028818f
C1524 VTAIL.n610 VSUBS 0.012909f
C1525 VTAIL.n611 VSUBS 0.022689f
C1526 VTAIL.n612 VSUBS 0.012192f
C1527 VTAIL.n613 VSUBS 0.028818f
C1528 VTAIL.n614 VSUBS 0.012909f
C1529 VTAIL.n615 VSUBS 0.022689f
C1530 VTAIL.n616 VSUBS 0.012192f
C1531 VTAIL.n617 VSUBS 0.028818f
C1532 VTAIL.n618 VSUBS 0.012909f
C1533 VTAIL.n619 VSUBS 1.71346f
C1534 VTAIL.n620 VSUBS 0.012192f
C1535 VTAIL.t2 VSUBS 0.061838f
C1536 VTAIL.n621 VSUBS 0.177138f
C1537 VTAIL.n622 VSUBS 0.018333f
C1538 VTAIL.n623 VSUBS 0.021613f
C1539 VTAIL.n624 VSUBS 0.028818f
C1540 VTAIL.n625 VSUBS 0.012909f
C1541 VTAIL.n626 VSUBS 0.012192f
C1542 VTAIL.n627 VSUBS 0.022689f
C1543 VTAIL.n628 VSUBS 0.022689f
C1544 VTAIL.n629 VSUBS 0.012192f
C1545 VTAIL.n630 VSUBS 0.012909f
C1546 VTAIL.n631 VSUBS 0.028818f
C1547 VTAIL.n632 VSUBS 0.028818f
C1548 VTAIL.n633 VSUBS 0.012909f
C1549 VTAIL.n634 VSUBS 0.012192f
C1550 VTAIL.n635 VSUBS 0.022689f
C1551 VTAIL.n636 VSUBS 0.022689f
C1552 VTAIL.n637 VSUBS 0.012192f
C1553 VTAIL.n638 VSUBS 0.012909f
C1554 VTAIL.n639 VSUBS 0.028818f
C1555 VTAIL.n640 VSUBS 0.028818f
C1556 VTAIL.n641 VSUBS 0.012909f
C1557 VTAIL.n642 VSUBS 0.012192f
C1558 VTAIL.n643 VSUBS 0.022689f
C1559 VTAIL.n644 VSUBS 0.022689f
C1560 VTAIL.n645 VSUBS 0.012192f
C1561 VTAIL.n646 VSUBS 0.012909f
C1562 VTAIL.n647 VSUBS 0.028818f
C1563 VTAIL.n648 VSUBS 0.028818f
C1564 VTAIL.n649 VSUBS 0.012909f
C1565 VTAIL.n650 VSUBS 0.012192f
C1566 VTAIL.n651 VSUBS 0.022689f
C1567 VTAIL.n652 VSUBS 0.022689f
C1568 VTAIL.n653 VSUBS 0.012192f
C1569 VTAIL.n654 VSUBS 0.012909f
C1570 VTAIL.n655 VSUBS 0.028818f
C1571 VTAIL.n656 VSUBS 0.028818f
C1572 VTAIL.n657 VSUBS 0.012909f
C1573 VTAIL.n658 VSUBS 0.012192f
C1574 VTAIL.n659 VSUBS 0.022689f
C1575 VTAIL.n660 VSUBS 0.022689f
C1576 VTAIL.n661 VSUBS 0.012192f
C1577 VTAIL.n662 VSUBS 0.012909f
C1578 VTAIL.n663 VSUBS 0.028818f
C1579 VTAIL.n664 VSUBS 0.028818f
C1580 VTAIL.n665 VSUBS 0.012909f
C1581 VTAIL.n666 VSUBS 0.012192f
C1582 VTAIL.n667 VSUBS 0.022689f
C1583 VTAIL.n668 VSUBS 0.022689f
C1584 VTAIL.n669 VSUBS 0.012192f
C1585 VTAIL.n670 VSUBS 0.012909f
C1586 VTAIL.n671 VSUBS 0.028818f
C1587 VTAIL.n672 VSUBS 0.028818f
C1588 VTAIL.n673 VSUBS 0.012909f
C1589 VTAIL.n674 VSUBS 0.012192f
C1590 VTAIL.n675 VSUBS 0.022689f
C1591 VTAIL.n676 VSUBS 0.022689f
C1592 VTAIL.n677 VSUBS 0.012192f
C1593 VTAIL.n678 VSUBS 0.012909f
C1594 VTAIL.n679 VSUBS 0.028818f
C1595 VTAIL.n680 VSUBS 0.069769f
C1596 VTAIL.n681 VSUBS 0.012909f
C1597 VTAIL.n682 VSUBS 0.012192f
C1598 VTAIL.n683 VSUBS 0.053995f
C1599 VTAIL.n684 VSUBS 0.035134f
C1600 VTAIL.n685 VSUBS 1.87447f
C1601 VTAIL.n686 VSUBS 0.024932f
C1602 VTAIL.n687 VSUBS 0.022689f
C1603 VTAIL.n688 VSUBS 0.012192f
C1604 VTAIL.n689 VSUBS 0.028818f
C1605 VTAIL.n690 VSUBS 0.012909f
C1606 VTAIL.n691 VSUBS 0.022689f
C1607 VTAIL.n692 VSUBS 0.012192f
C1608 VTAIL.n693 VSUBS 0.028818f
C1609 VTAIL.n694 VSUBS 0.012551f
C1610 VTAIL.n695 VSUBS 0.022689f
C1611 VTAIL.n696 VSUBS 0.012909f
C1612 VTAIL.n697 VSUBS 0.028818f
C1613 VTAIL.n698 VSUBS 0.012909f
C1614 VTAIL.n699 VSUBS 0.022689f
C1615 VTAIL.n700 VSUBS 0.012192f
C1616 VTAIL.n701 VSUBS 0.028818f
C1617 VTAIL.n702 VSUBS 0.012909f
C1618 VTAIL.n703 VSUBS 0.022689f
C1619 VTAIL.n704 VSUBS 0.012192f
C1620 VTAIL.n705 VSUBS 0.028818f
C1621 VTAIL.n706 VSUBS 0.012909f
C1622 VTAIL.n707 VSUBS 0.022689f
C1623 VTAIL.n708 VSUBS 0.012192f
C1624 VTAIL.n709 VSUBS 0.028818f
C1625 VTAIL.n710 VSUBS 0.012909f
C1626 VTAIL.n711 VSUBS 0.022689f
C1627 VTAIL.n712 VSUBS 0.012192f
C1628 VTAIL.n713 VSUBS 0.028818f
C1629 VTAIL.n714 VSUBS 0.012909f
C1630 VTAIL.n715 VSUBS 1.71346f
C1631 VTAIL.n716 VSUBS 0.012192f
C1632 VTAIL.t7 VSUBS 0.061838f
C1633 VTAIL.n717 VSUBS 0.177138f
C1634 VTAIL.n718 VSUBS 0.018333f
C1635 VTAIL.n719 VSUBS 0.021613f
C1636 VTAIL.n720 VSUBS 0.028818f
C1637 VTAIL.n721 VSUBS 0.012909f
C1638 VTAIL.n722 VSUBS 0.012192f
C1639 VTAIL.n723 VSUBS 0.022689f
C1640 VTAIL.n724 VSUBS 0.022689f
C1641 VTAIL.n725 VSUBS 0.012192f
C1642 VTAIL.n726 VSUBS 0.012909f
C1643 VTAIL.n727 VSUBS 0.028818f
C1644 VTAIL.n728 VSUBS 0.028818f
C1645 VTAIL.n729 VSUBS 0.012909f
C1646 VTAIL.n730 VSUBS 0.012192f
C1647 VTAIL.n731 VSUBS 0.022689f
C1648 VTAIL.n732 VSUBS 0.022689f
C1649 VTAIL.n733 VSUBS 0.012192f
C1650 VTAIL.n734 VSUBS 0.012909f
C1651 VTAIL.n735 VSUBS 0.028818f
C1652 VTAIL.n736 VSUBS 0.028818f
C1653 VTAIL.n737 VSUBS 0.012909f
C1654 VTAIL.n738 VSUBS 0.012192f
C1655 VTAIL.n739 VSUBS 0.022689f
C1656 VTAIL.n740 VSUBS 0.022689f
C1657 VTAIL.n741 VSUBS 0.012192f
C1658 VTAIL.n742 VSUBS 0.012909f
C1659 VTAIL.n743 VSUBS 0.028818f
C1660 VTAIL.n744 VSUBS 0.028818f
C1661 VTAIL.n745 VSUBS 0.012909f
C1662 VTAIL.n746 VSUBS 0.012192f
C1663 VTAIL.n747 VSUBS 0.022689f
C1664 VTAIL.n748 VSUBS 0.022689f
C1665 VTAIL.n749 VSUBS 0.012192f
C1666 VTAIL.n750 VSUBS 0.012909f
C1667 VTAIL.n751 VSUBS 0.028818f
C1668 VTAIL.n752 VSUBS 0.028818f
C1669 VTAIL.n753 VSUBS 0.012909f
C1670 VTAIL.n754 VSUBS 0.012192f
C1671 VTAIL.n755 VSUBS 0.022689f
C1672 VTAIL.n756 VSUBS 0.022689f
C1673 VTAIL.n757 VSUBS 0.012192f
C1674 VTAIL.n758 VSUBS 0.012192f
C1675 VTAIL.n759 VSUBS 0.012909f
C1676 VTAIL.n760 VSUBS 0.028818f
C1677 VTAIL.n761 VSUBS 0.028818f
C1678 VTAIL.n762 VSUBS 0.028818f
C1679 VTAIL.n763 VSUBS 0.012551f
C1680 VTAIL.n764 VSUBS 0.012192f
C1681 VTAIL.n765 VSUBS 0.022689f
C1682 VTAIL.n766 VSUBS 0.022689f
C1683 VTAIL.n767 VSUBS 0.012192f
C1684 VTAIL.n768 VSUBS 0.012909f
C1685 VTAIL.n769 VSUBS 0.028818f
C1686 VTAIL.n770 VSUBS 0.028818f
C1687 VTAIL.n771 VSUBS 0.012909f
C1688 VTAIL.n772 VSUBS 0.012192f
C1689 VTAIL.n773 VSUBS 0.022689f
C1690 VTAIL.n774 VSUBS 0.022689f
C1691 VTAIL.n775 VSUBS 0.012192f
C1692 VTAIL.n776 VSUBS 0.012909f
C1693 VTAIL.n777 VSUBS 0.028818f
C1694 VTAIL.n778 VSUBS 0.069769f
C1695 VTAIL.n779 VSUBS 0.012909f
C1696 VTAIL.n780 VSUBS 0.012192f
C1697 VTAIL.n781 VSUBS 0.053995f
C1698 VTAIL.n782 VSUBS 0.035134f
C1699 VTAIL.n783 VSUBS 1.76055f
C1700 VN.t0 VSUBS 4.3741f
C1701 VN.t2 VSUBS 4.38408f
C1702 VN.n0 VSUBS 2.73872f
C1703 VN.t3 VSUBS 4.3741f
C1704 VN.t1 VSUBS 4.38408f
C1705 VN.n1 VSUBS 4.54006f
.ends

