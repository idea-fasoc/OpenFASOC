* NGSPICE file created from diff_pair_sample_0082.ext - technology: sky130A

.subckt diff_pair_sample_0082 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t9 VN.t0 VTAIL.t12 B.t3 sky130_fd_pr__nfet_01v8 ad=2.2581 pd=12.36 as=0.95535 ps=6.12 w=5.79 l=0.57
X1 VDD1.t9 VP.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.95535 pd=6.12 as=2.2581 ps=12.36 w=5.79 l=0.57
X2 VDD1.t8 VP.t1 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=0.95535 pd=6.12 as=2.2581 ps=12.36 w=5.79 l=0.57
X3 VTAIL.t11 VN.t1 VDD2.t8 B.t6 sky130_fd_pr__nfet_01v8 ad=0.95535 pd=6.12 as=0.95535 ps=6.12 w=5.79 l=0.57
X4 VTAIL.t2 VP.t2 VDD1.t7 B.t2 sky130_fd_pr__nfet_01v8 ad=0.95535 pd=6.12 as=0.95535 ps=6.12 w=5.79 l=0.57
X5 VTAIL.t10 VN.t2 VDD2.t7 B.t9 sky130_fd_pr__nfet_01v8 ad=0.95535 pd=6.12 as=0.95535 ps=6.12 w=5.79 l=0.57
X6 VTAIL.t7 VP.t3 VDD1.t6 B.t7 sky130_fd_pr__nfet_01v8 ad=0.95535 pd=6.12 as=0.95535 ps=6.12 w=5.79 l=0.57
X7 VTAIL.t9 VN.t3 VDD2.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=0.95535 pd=6.12 as=0.95535 ps=6.12 w=5.79 l=0.57
X8 VDD2.t5 VN.t4 VTAIL.t13 B.t4 sky130_fd_pr__nfet_01v8 ad=0.95535 pd=6.12 as=0.95535 ps=6.12 w=5.79 l=0.57
X9 B.t23 B.t21 B.t22 B.t15 sky130_fd_pr__nfet_01v8 ad=2.2581 pd=12.36 as=0 ps=0 w=5.79 l=0.57
X10 VDD2.t4 VN.t5 VTAIL.t16 B.t8 sky130_fd_pr__nfet_01v8 ad=0.95535 pd=6.12 as=0.95535 ps=6.12 w=5.79 l=0.57
X11 VDD1.t5 VP.t4 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=0.95535 pd=6.12 as=0.95535 ps=6.12 w=5.79 l=0.57
X12 VTAIL.t17 VN.t6 VDD2.t3 B.t7 sky130_fd_pr__nfet_01v8 ad=0.95535 pd=6.12 as=0.95535 ps=6.12 w=5.79 l=0.57
X13 B.t20 B.t18 B.t19 B.t11 sky130_fd_pr__nfet_01v8 ad=2.2581 pd=12.36 as=0 ps=0 w=5.79 l=0.57
X14 VTAIL.t18 VP.t5 VDD1.t4 B.t9 sky130_fd_pr__nfet_01v8 ad=0.95535 pd=6.12 as=0.95535 ps=6.12 w=5.79 l=0.57
X15 VDD2.t2 VN.t7 VTAIL.t14 B.t5 sky130_fd_pr__nfet_01v8 ad=0.95535 pd=6.12 as=2.2581 ps=12.36 w=5.79 l=0.57
X16 VTAIL.t6 VP.t6 VDD1.t3 B.t6 sky130_fd_pr__nfet_01v8 ad=0.95535 pd=6.12 as=0.95535 ps=6.12 w=5.79 l=0.57
X17 VDD1.t2 VP.t7 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.2581 pd=12.36 as=0.95535 ps=6.12 w=5.79 l=0.57
X18 VDD1.t1 VP.t8 VTAIL.t19 B.t8 sky130_fd_pr__nfet_01v8 ad=0.95535 pd=6.12 as=0.95535 ps=6.12 w=5.79 l=0.57
X19 VDD2.t1 VN.t8 VTAIL.t8 B.t1 sky130_fd_pr__nfet_01v8 ad=0.95535 pd=6.12 as=2.2581 ps=12.36 w=5.79 l=0.57
X20 VDD2.t0 VN.t9 VTAIL.t15 B.t0 sky130_fd_pr__nfet_01v8 ad=2.2581 pd=12.36 as=0.95535 ps=6.12 w=5.79 l=0.57
X21 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=2.2581 pd=12.36 as=0 ps=0 w=5.79 l=0.57
X22 VDD1.t0 VP.t9 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.2581 pd=12.36 as=0.95535 ps=6.12 w=5.79 l=0.57
X23 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=2.2581 pd=12.36 as=0 ps=0 w=5.79 l=0.57
R0 VN.n3 VN.t9 338.866
R1 VN.n13 VN.t7 338.866
R2 VN.n2 VN.t2 314.147
R3 VN.n1 VN.t4 314.147
R4 VN.n6 VN.t3 314.147
R5 VN.n8 VN.t8 314.147
R6 VN.n12 VN.t6 314.147
R7 VN.n11 VN.t5 314.147
R8 VN.n16 VN.t1 314.147
R9 VN.n18 VN.t0 314.147
R10 VN.n9 VN.n8 161.3
R11 VN.n19 VN.n18 161.3
R12 VN.n17 VN.n10 161.3
R13 VN.n16 VN.n15 161.3
R14 VN.n7 VN.n0 161.3
R15 VN.n6 VN.n5 161.3
R16 VN.n14 VN.n11 80.6037
R17 VN.n4 VN.n1 80.6037
R18 VN.n2 VN.n1 48.2005
R19 VN.n6 VN.n1 48.2005
R20 VN.n12 VN.n11 48.2005
R21 VN.n16 VN.n11 48.2005
R22 VN.n14 VN.n13 45.0526
R23 VN.n4 VN.n3 45.0526
R24 VN.n8 VN.n7 38.7066
R25 VN.n18 VN.n17 38.7066
R26 VN VN.n19 37.7145
R27 VN.n3 VN.n2 16.5858
R28 VN.n13 VN.n12 16.5858
R29 VN.n7 VN.n6 9.49444
R30 VN.n17 VN.n16 9.49444
R31 VN.n15 VN.n14 0.285035
R32 VN.n5 VN.n4 0.285035
R33 VN.n19 VN.n10 0.189894
R34 VN.n15 VN.n10 0.189894
R35 VN.n5 VN.n0 0.189894
R36 VN.n9 VN.n0 0.189894
R37 VN VN.n9 0.0516364
R38 VTAIL.n132 VTAIL.n131 289.615
R39 VTAIL.n30 VTAIL.n29 289.615
R40 VTAIL.n102 VTAIL.n101 289.615
R41 VTAIL.n68 VTAIL.n67 289.615
R42 VTAIL.n115 VTAIL.n114 185
R43 VTAIL.n117 VTAIL.n116 185
R44 VTAIL.n110 VTAIL.n109 185
R45 VTAIL.n123 VTAIL.n122 185
R46 VTAIL.n125 VTAIL.n124 185
R47 VTAIL.n106 VTAIL.n105 185
R48 VTAIL.n131 VTAIL.n130 185
R49 VTAIL.n13 VTAIL.n12 185
R50 VTAIL.n15 VTAIL.n14 185
R51 VTAIL.n8 VTAIL.n7 185
R52 VTAIL.n21 VTAIL.n20 185
R53 VTAIL.n23 VTAIL.n22 185
R54 VTAIL.n4 VTAIL.n3 185
R55 VTAIL.n29 VTAIL.n28 185
R56 VTAIL.n101 VTAIL.n100 185
R57 VTAIL.n76 VTAIL.n75 185
R58 VTAIL.n95 VTAIL.n94 185
R59 VTAIL.n93 VTAIL.n92 185
R60 VTAIL.n80 VTAIL.n79 185
R61 VTAIL.n87 VTAIL.n86 185
R62 VTAIL.n85 VTAIL.n84 185
R63 VTAIL.n67 VTAIL.n66 185
R64 VTAIL.n42 VTAIL.n41 185
R65 VTAIL.n61 VTAIL.n60 185
R66 VTAIL.n59 VTAIL.n58 185
R67 VTAIL.n46 VTAIL.n45 185
R68 VTAIL.n53 VTAIL.n52 185
R69 VTAIL.n51 VTAIL.n50 185
R70 VTAIL.n113 VTAIL.t8 149.528
R71 VTAIL.n11 VTAIL.t5 149.528
R72 VTAIL.n83 VTAIL.t1 149.528
R73 VTAIL.n49 VTAIL.t14 149.528
R74 VTAIL.n116 VTAIL.n115 104.615
R75 VTAIL.n116 VTAIL.n109 104.615
R76 VTAIL.n123 VTAIL.n109 104.615
R77 VTAIL.n124 VTAIL.n123 104.615
R78 VTAIL.n124 VTAIL.n105 104.615
R79 VTAIL.n131 VTAIL.n105 104.615
R80 VTAIL.n14 VTAIL.n13 104.615
R81 VTAIL.n14 VTAIL.n7 104.615
R82 VTAIL.n21 VTAIL.n7 104.615
R83 VTAIL.n22 VTAIL.n21 104.615
R84 VTAIL.n22 VTAIL.n3 104.615
R85 VTAIL.n29 VTAIL.n3 104.615
R86 VTAIL.n101 VTAIL.n75 104.615
R87 VTAIL.n94 VTAIL.n75 104.615
R88 VTAIL.n94 VTAIL.n93 104.615
R89 VTAIL.n93 VTAIL.n79 104.615
R90 VTAIL.n86 VTAIL.n79 104.615
R91 VTAIL.n86 VTAIL.n85 104.615
R92 VTAIL.n67 VTAIL.n41 104.615
R93 VTAIL.n60 VTAIL.n41 104.615
R94 VTAIL.n60 VTAIL.n59 104.615
R95 VTAIL.n59 VTAIL.n45 104.615
R96 VTAIL.n52 VTAIL.n45 104.615
R97 VTAIL.n52 VTAIL.n51 104.615
R98 VTAIL.n73 VTAIL.n72 52.6055
R99 VTAIL.n71 VTAIL.n70 52.6055
R100 VTAIL.n39 VTAIL.n38 52.6055
R101 VTAIL.n37 VTAIL.n36 52.6055
R102 VTAIL.n135 VTAIL.n134 52.6045
R103 VTAIL.n1 VTAIL.n0 52.6045
R104 VTAIL.n33 VTAIL.n32 52.6045
R105 VTAIL.n35 VTAIL.n34 52.6045
R106 VTAIL.n115 VTAIL.t8 52.3082
R107 VTAIL.n13 VTAIL.t5 52.3082
R108 VTAIL.n85 VTAIL.t1 52.3082
R109 VTAIL.n51 VTAIL.t14 52.3082
R110 VTAIL.n133 VTAIL.n132 33.9308
R111 VTAIL.n31 VTAIL.n30 33.9308
R112 VTAIL.n103 VTAIL.n102 33.9308
R113 VTAIL.n69 VTAIL.n68 33.9308
R114 VTAIL.n37 VTAIL.n35 18.91
R115 VTAIL.n133 VTAIL.n103 18.1341
R116 VTAIL.n130 VTAIL.n104 12.0247
R117 VTAIL.n28 VTAIL.n2 12.0247
R118 VTAIL.n100 VTAIL.n74 12.0247
R119 VTAIL.n66 VTAIL.n40 12.0247
R120 VTAIL.n129 VTAIL.n106 11.249
R121 VTAIL.n27 VTAIL.n4 11.249
R122 VTAIL.n99 VTAIL.n76 11.249
R123 VTAIL.n65 VTAIL.n42 11.249
R124 VTAIL.n126 VTAIL.n125 10.4732
R125 VTAIL.n24 VTAIL.n23 10.4732
R126 VTAIL.n96 VTAIL.n95 10.4732
R127 VTAIL.n62 VTAIL.n61 10.4732
R128 VTAIL.n114 VTAIL.n113 10.2745
R129 VTAIL.n12 VTAIL.n11 10.2745
R130 VTAIL.n84 VTAIL.n83 10.2745
R131 VTAIL.n50 VTAIL.n49 10.2745
R132 VTAIL.n122 VTAIL.n108 9.69747
R133 VTAIL.n20 VTAIL.n6 9.69747
R134 VTAIL.n92 VTAIL.n78 9.69747
R135 VTAIL.n58 VTAIL.n44 9.69747
R136 VTAIL.n128 VTAIL.n104 9.45567
R137 VTAIL.n26 VTAIL.n2 9.45567
R138 VTAIL.n98 VTAIL.n74 9.45567
R139 VTAIL.n64 VTAIL.n40 9.45567
R140 VTAIL.n112 VTAIL.n111 9.3005
R141 VTAIL.n119 VTAIL.n118 9.3005
R142 VTAIL.n121 VTAIL.n120 9.3005
R143 VTAIL.n108 VTAIL.n107 9.3005
R144 VTAIL.n127 VTAIL.n126 9.3005
R145 VTAIL.n129 VTAIL.n128 9.3005
R146 VTAIL.n10 VTAIL.n9 9.3005
R147 VTAIL.n17 VTAIL.n16 9.3005
R148 VTAIL.n19 VTAIL.n18 9.3005
R149 VTAIL.n6 VTAIL.n5 9.3005
R150 VTAIL.n25 VTAIL.n24 9.3005
R151 VTAIL.n27 VTAIL.n26 9.3005
R152 VTAIL.n99 VTAIL.n98 9.3005
R153 VTAIL.n97 VTAIL.n96 9.3005
R154 VTAIL.n78 VTAIL.n77 9.3005
R155 VTAIL.n91 VTAIL.n90 9.3005
R156 VTAIL.n89 VTAIL.n88 9.3005
R157 VTAIL.n82 VTAIL.n81 9.3005
R158 VTAIL.n55 VTAIL.n54 9.3005
R159 VTAIL.n57 VTAIL.n56 9.3005
R160 VTAIL.n44 VTAIL.n43 9.3005
R161 VTAIL.n63 VTAIL.n62 9.3005
R162 VTAIL.n65 VTAIL.n64 9.3005
R163 VTAIL.n48 VTAIL.n47 9.3005
R164 VTAIL.n121 VTAIL.n110 8.92171
R165 VTAIL.n19 VTAIL.n8 8.92171
R166 VTAIL.n91 VTAIL.n80 8.92171
R167 VTAIL.n57 VTAIL.n46 8.92171
R168 VTAIL.n118 VTAIL.n117 8.14595
R169 VTAIL.n16 VTAIL.n15 8.14595
R170 VTAIL.n88 VTAIL.n87 8.14595
R171 VTAIL.n54 VTAIL.n53 8.14595
R172 VTAIL.n114 VTAIL.n112 7.3702
R173 VTAIL.n12 VTAIL.n10 7.3702
R174 VTAIL.n84 VTAIL.n82 7.3702
R175 VTAIL.n50 VTAIL.n48 7.3702
R176 VTAIL.n117 VTAIL.n112 5.81868
R177 VTAIL.n15 VTAIL.n10 5.81868
R178 VTAIL.n87 VTAIL.n82 5.81868
R179 VTAIL.n53 VTAIL.n48 5.81868
R180 VTAIL.n118 VTAIL.n110 5.04292
R181 VTAIL.n16 VTAIL.n8 5.04292
R182 VTAIL.n88 VTAIL.n80 5.04292
R183 VTAIL.n54 VTAIL.n46 5.04292
R184 VTAIL.n122 VTAIL.n121 4.26717
R185 VTAIL.n20 VTAIL.n19 4.26717
R186 VTAIL.n92 VTAIL.n91 4.26717
R187 VTAIL.n58 VTAIL.n57 4.26717
R188 VTAIL.n125 VTAIL.n108 3.49141
R189 VTAIL.n23 VTAIL.n6 3.49141
R190 VTAIL.n95 VTAIL.n78 3.49141
R191 VTAIL.n61 VTAIL.n44 3.49141
R192 VTAIL.n134 VTAIL.t13 3.42019
R193 VTAIL.n134 VTAIL.t9 3.42019
R194 VTAIL.n0 VTAIL.t15 3.42019
R195 VTAIL.n0 VTAIL.t10 3.42019
R196 VTAIL.n32 VTAIL.t19 3.42019
R197 VTAIL.n32 VTAIL.t7 3.42019
R198 VTAIL.n34 VTAIL.t3 3.42019
R199 VTAIL.n34 VTAIL.t6 3.42019
R200 VTAIL.n72 VTAIL.t4 3.42019
R201 VTAIL.n72 VTAIL.t2 3.42019
R202 VTAIL.n70 VTAIL.t0 3.42019
R203 VTAIL.n70 VTAIL.t18 3.42019
R204 VTAIL.n38 VTAIL.t16 3.42019
R205 VTAIL.n38 VTAIL.t17 3.42019
R206 VTAIL.n36 VTAIL.t12 3.42019
R207 VTAIL.n36 VTAIL.t11 3.42019
R208 VTAIL.n83 VTAIL.n81 2.84323
R209 VTAIL.n49 VTAIL.n47 2.84323
R210 VTAIL.n113 VTAIL.n111 2.84323
R211 VTAIL.n11 VTAIL.n9 2.84323
R212 VTAIL.n126 VTAIL.n106 2.71565
R213 VTAIL.n24 VTAIL.n4 2.71565
R214 VTAIL.n96 VTAIL.n76 2.71565
R215 VTAIL.n62 VTAIL.n42 2.71565
R216 VTAIL.n130 VTAIL.n129 1.93989
R217 VTAIL.n28 VTAIL.n27 1.93989
R218 VTAIL.n100 VTAIL.n99 1.93989
R219 VTAIL.n66 VTAIL.n65 1.93989
R220 VTAIL.n132 VTAIL.n104 1.16414
R221 VTAIL.n30 VTAIL.n2 1.16414
R222 VTAIL.n102 VTAIL.n74 1.16414
R223 VTAIL.n68 VTAIL.n40 1.16414
R224 VTAIL.n71 VTAIL.n69 0.858259
R225 VTAIL.n31 VTAIL.n1 0.858259
R226 VTAIL.n39 VTAIL.n37 0.776362
R227 VTAIL.n69 VTAIL.n39 0.776362
R228 VTAIL.n73 VTAIL.n71 0.776362
R229 VTAIL.n103 VTAIL.n73 0.776362
R230 VTAIL.n35 VTAIL.n33 0.776362
R231 VTAIL.n33 VTAIL.n31 0.776362
R232 VTAIL.n135 VTAIL.n133 0.776362
R233 VTAIL VTAIL.n1 0.640586
R234 VTAIL.n119 VTAIL.n111 0.155672
R235 VTAIL.n120 VTAIL.n119 0.155672
R236 VTAIL.n120 VTAIL.n107 0.155672
R237 VTAIL.n127 VTAIL.n107 0.155672
R238 VTAIL.n128 VTAIL.n127 0.155672
R239 VTAIL.n17 VTAIL.n9 0.155672
R240 VTAIL.n18 VTAIL.n17 0.155672
R241 VTAIL.n18 VTAIL.n5 0.155672
R242 VTAIL.n25 VTAIL.n5 0.155672
R243 VTAIL.n26 VTAIL.n25 0.155672
R244 VTAIL.n98 VTAIL.n97 0.155672
R245 VTAIL.n97 VTAIL.n77 0.155672
R246 VTAIL.n90 VTAIL.n77 0.155672
R247 VTAIL.n90 VTAIL.n89 0.155672
R248 VTAIL.n89 VTAIL.n81 0.155672
R249 VTAIL.n64 VTAIL.n63 0.155672
R250 VTAIL.n63 VTAIL.n43 0.155672
R251 VTAIL.n56 VTAIL.n43 0.155672
R252 VTAIL.n56 VTAIL.n55 0.155672
R253 VTAIL.n55 VTAIL.n47 0.155672
R254 VTAIL VTAIL.n135 0.136276
R255 VDD2.n61 VDD2.n60 289.615
R256 VDD2.n28 VDD2.n27 289.615
R257 VDD2.n60 VDD2.n59 185
R258 VDD2.n35 VDD2.n34 185
R259 VDD2.n54 VDD2.n53 185
R260 VDD2.n52 VDD2.n51 185
R261 VDD2.n39 VDD2.n38 185
R262 VDD2.n46 VDD2.n45 185
R263 VDD2.n44 VDD2.n43 185
R264 VDD2.n11 VDD2.n10 185
R265 VDD2.n13 VDD2.n12 185
R266 VDD2.n6 VDD2.n5 185
R267 VDD2.n19 VDD2.n18 185
R268 VDD2.n21 VDD2.n20 185
R269 VDD2.n2 VDD2.n1 185
R270 VDD2.n27 VDD2.n26 185
R271 VDD2.n42 VDD2.t9 149.528
R272 VDD2.n9 VDD2.t0 149.528
R273 VDD2.n60 VDD2.n34 104.615
R274 VDD2.n53 VDD2.n34 104.615
R275 VDD2.n53 VDD2.n52 104.615
R276 VDD2.n52 VDD2.n38 104.615
R277 VDD2.n45 VDD2.n38 104.615
R278 VDD2.n45 VDD2.n44 104.615
R279 VDD2.n12 VDD2.n11 104.615
R280 VDD2.n12 VDD2.n5 104.615
R281 VDD2.n19 VDD2.n5 104.615
R282 VDD2.n20 VDD2.n19 104.615
R283 VDD2.n20 VDD2.n1 104.615
R284 VDD2.n27 VDD2.n1 104.615
R285 VDD2.n32 VDD2.n31 69.8098
R286 VDD2 VDD2.n65 69.8068
R287 VDD2.n64 VDD2.n63 69.2843
R288 VDD2.n30 VDD2.n29 69.2833
R289 VDD2.n44 VDD2.t9 52.3082
R290 VDD2.n11 VDD2.t0 52.3082
R291 VDD2.n30 VDD2.n28 51.3855
R292 VDD2.n62 VDD2.n61 50.6096
R293 VDD2.n62 VDD2.n32 32.392
R294 VDD2.n59 VDD2.n33 12.0247
R295 VDD2.n26 VDD2.n0 12.0247
R296 VDD2.n58 VDD2.n35 11.249
R297 VDD2.n25 VDD2.n2 11.249
R298 VDD2.n55 VDD2.n54 10.4732
R299 VDD2.n22 VDD2.n21 10.4732
R300 VDD2.n43 VDD2.n42 10.2745
R301 VDD2.n10 VDD2.n9 10.2745
R302 VDD2.n51 VDD2.n37 9.69747
R303 VDD2.n18 VDD2.n4 9.69747
R304 VDD2.n57 VDD2.n33 9.45567
R305 VDD2.n24 VDD2.n0 9.45567
R306 VDD2.n48 VDD2.n47 9.3005
R307 VDD2.n50 VDD2.n49 9.3005
R308 VDD2.n37 VDD2.n36 9.3005
R309 VDD2.n56 VDD2.n55 9.3005
R310 VDD2.n58 VDD2.n57 9.3005
R311 VDD2.n41 VDD2.n40 9.3005
R312 VDD2.n8 VDD2.n7 9.3005
R313 VDD2.n15 VDD2.n14 9.3005
R314 VDD2.n17 VDD2.n16 9.3005
R315 VDD2.n4 VDD2.n3 9.3005
R316 VDD2.n23 VDD2.n22 9.3005
R317 VDD2.n25 VDD2.n24 9.3005
R318 VDD2.n50 VDD2.n39 8.92171
R319 VDD2.n17 VDD2.n6 8.92171
R320 VDD2.n47 VDD2.n46 8.14595
R321 VDD2.n14 VDD2.n13 8.14595
R322 VDD2.n43 VDD2.n41 7.3702
R323 VDD2.n10 VDD2.n8 7.3702
R324 VDD2.n46 VDD2.n41 5.81868
R325 VDD2.n13 VDD2.n8 5.81868
R326 VDD2.n47 VDD2.n39 5.04292
R327 VDD2.n14 VDD2.n6 5.04292
R328 VDD2.n51 VDD2.n50 4.26717
R329 VDD2.n18 VDD2.n17 4.26717
R330 VDD2.n54 VDD2.n37 3.49141
R331 VDD2.n21 VDD2.n4 3.49141
R332 VDD2.n65 VDD2.t3 3.42019
R333 VDD2.n65 VDD2.t2 3.42019
R334 VDD2.n63 VDD2.t8 3.42019
R335 VDD2.n63 VDD2.t4 3.42019
R336 VDD2.n31 VDD2.t6 3.42019
R337 VDD2.n31 VDD2.t1 3.42019
R338 VDD2.n29 VDD2.t7 3.42019
R339 VDD2.n29 VDD2.t5 3.42019
R340 VDD2.n42 VDD2.n40 2.84323
R341 VDD2.n9 VDD2.n7 2.84323
R342 VDD2.n55 VDD2.n35 2.71565
R343 VDD2.n22 VDD2.n2 2.71565
R344 VDD2.n59 VDD2.n58 1.93989
R345 VDD2.n26 VDD2.n25 1.93989
R346 VDD2.n61 VDD2.n33 1.16414
R347 VDD2.n28 VDD2.n0 1.16414
R348 VDD2.n64 VDD2.n62 0.776362
R349 VDD2 VDD2.n64 0.252655
R350 VDD2.n57 VDD2.n56 0.155672
R351 VDD2.n56 VDD2.n36 0.155672
R352 VDD2.n49 VDD2.n36 0.155672
R353 VDD2.n49 VDD2.n48 0.155672
R354 VDD2.n48 VDD2.n40 0.155672
R355 VDD2.n15 VDD2.n7 0.155672
R356 VDD2.n16 VDD2.n15 0.155672
R357 VDD2.n16 VDD2.n3 0.155672
R358 VDD2.n23 VDD2.n3 0.155672
R359 VDD2.n24 VDD2.n23 0.155672
R360 VDD2.n32 VDD2.n30 0.139119
R361 B.n484 B.n483 585
R362 B.n188 B.n75 585
R363 B.n187 B.n186 585
R364 B.n185 B.n184 585
R365 B.n183 B.n182 585
R366 B.n181 B.n180 585
R367 B.n179 B.n178 585
R368 B.n177 B.n176 585
R369 B.n175 B.n174 585
R370 B.n173 B.n172 585
R371 B.n171 B.n170 585
R372 B.n169 B.n168 585
R373 B.n167 B.n166 585
R374 B.n165 B.n164 585
R375 B.n163 B.n162 585
R376 B.n161 B.n160 585
R377 B.n159 B.n158 585
R378 B.n157 B.n156 585
R379 B.n155 B.n154 585
R380 B.n153 B.n152 585
R381 B.n151 B.n150 585
R382 B.n149 B.n148 585
R383 B.n147 B.n146 585
R384 B.n144 B.n143 585
R385 B.n142 B.n141 585
R386 B.n140 B.n139 585
R387 B.n138 B.n137 585
R388 B.n136 B.n135 585
R389 B.n134 B.n133 585
R390 B.n132 B.n131 585
R391 B.n130 B.n129 585
R392 B.n128 B.n127 585
R393 B.n126 B.n125 585
R394 B.n123 B.n122 585
R395 B.n121 B.n120 585
R396 B.n119 B.n118 585
R397 B.n117 B.n116 585
R398 B.n115 B.n114 585
R399 B.n113 B.n112 585
R400 B.n111 B.n110 585
R401 B.n109 B.n108 585
R402 B.n107 B.n106 585
R403 B.n105 B.n104 585
R404 B.n103 B.n102 585
R405 B.n101 B.n100 585
R406 B.n99 B.n98 585
R407 B.n97 B.n96 585
R408 B.n95 B.n94 585
R409 B.n93 B.n92 585
R410 B.n91 B.n90 585
R411 B.n89 B.n88 585
R412 B.n87 B.n86 585
R413 B.n85 B.n84 585
R414 B.n83 B.n82 585
R415 B.n81 B.n80 585
R416 B.n46 B.n45 585
R417 B.n482 B.n47 585
R418 B.n487 B.n47 585
R419 B.n481 B.n480 585
R420 B.n480 B.n43 585
R421 B.n479 B.n42 585
R422 B.n493 B.n42 585
R423 B.n478 B.n41 585
R424 B.n494 B.n41 585
R425 B.n477 B.n40 585
R426 B.n495 B.n40 585
R427 B.n476 B.n475 585
R428 B.n475 B.n36 585
R429 B.n474 B.n35 585
R430 B.n501 B.n35 585
R431 B.n473 B.n34 585
R432 B.n502 B.n34 585
R433 B.n472 B.n33 585
R434 B.n503 B.n33 585
R435 B.n471 B.n470 585
R436 B.n470 B.n29 585
R437 B.n469 B.n28 585
R438 B.n509 B.n28 585
R439 B.n468 B.n27 585
R440 B.n510 B.n27 585
R441 B.n467 B.n26 585
R442 B.n511 B.n26 585
R443 B.n466 B.n465 585
R444 B.n465 B.n25 585
R445 B.n464 B.n21 585
R446 B.n517 B.n21 585
R447 B.n463 B.n20 585
R448 B.n518 B.n20 585
R449 B.n462 B.n19 585
R450 B.n519 B.n19 585
R451 B.n461 B.n460 585
R452 B.n460 B.n15 585
R453 B.n459 B.n14 585
R454 B.n525 B.n14 585
R455 B.n458 B.n13 585
R456 B.n526 B.n13 585
R457 B.n457 B.n12 585
R458 B.n527 B.n12 585
R459 B.n456 B.n455 585
R460 B.n455 B.n11 585
R461 B.n454 B.n7 585
R462 B.n533 B.n7 585
R463 B.n453 B.n6 585
R464 B.n534 B.n6 585
R465 B.n452 B.n5 585
R466 B.n535 B.n5 585
R467 B.n451 B.n450 585
R468 B.n450 B.n4 585
R469 B.n449 B.n189 585
R470 B.n449 B.n448 585
R471 B.n438 B.n190 585
R472 B.n441 B.n190 585
R473 B.n440 B.n439 585
R474 B.n442 B.n440 585
R475 B.n437 B.n195 585
R476 B.n195 B.n194 585
R477 B.n436 B.n435 585
R478 B.n435 B.n434 585
R479 B.n197 B.n196 585
R480 B.n198 B.n197 585
R481 B.n427 B.n426 585
R482 B.n428 B.n427 585
R483 B.n425 B.n202 585
R484 B.n205 B.n202 585
R485 B.n424 B.n423 585
R486 B.n423 B.n422 585
R487 B.n204 B.n203 585
R488 B.n415 B.n204 585
R489 B.n414 B.n413 585
R490 B.n416 B.n414 585
R491 B.n412 B.n210 585
R492 B.n210 B.n209 585
R493 B.n411 B.n410 585
R494 B.n410 B.n409 585
R495 B.n212 B.n211 585
R496 B.n213 B.n212 585
R497 B.n402 B.n401 585
R498 B.n403 B.n402 585
R499 B.n400 B.n218 585
R500 B.n218 B.n217 585
R501 B.n399 B.n398 585
R502 B.n398 B.n397 585
R503 B.n220 B.n219 585
R504 B.n221 B.n220 585
R505 B.n390 B.n389 585
R506 B.n391 B.n390 585
R507 B.n388 B.n226 585
R508 B.n226 B.n225 585
R509 B.n387 B.n386 585
R510 B.n386 B.n385 585
R511 B.n228 B.n227 585
R512 B.n229 B.n228 585
R513 B.n378 B.n377 585
R514 B.n379 B.n378 585
R515 B.n232 B.n231 585
R516 B.n269 B.n268 585
R517 B.n270 B.n266 585
R518 B.n266 B.n233 585
R519 B.n272 B.n271 585
R520 B.n274 B.n265 585
R521 B.n277 B.n276 585
R522 B.n278 B.n264 585
R523 B.n280 B.n279 585
R524 B.n282 B.n263 585
R525 B.n285 B.n284 585
R526 B.n286 B.n262 585
R527 B.n288 B.n287 585
R528 B.n290 B.n261 585
R529 B.n293 B.n292 585
R530 B.n294 B.n260 585
R531 B.n296 B.n295 585
R532 B.n298 B.n259 585
R533 B.n301 B.n300 585
R534 B.n302 B.n258 585
R535 B.n304 B.n303 585
R536 B.n306 B.n257 585
R537 B.n309 B.n308 585
R538 B.n310 B.n254 585
R539 B.n313 B.n312 585
R540 B.n315 B.n253 585
R541 B.n318 B.n317 585
R542 B.n319 B.n252 585
R543 B.n321 B.n320 585
R544 B.n323 B.n251 585
R545 B.n326 B.n325 585
R546 B.n327 B.n250 585
R547 B.n329 B.n328 585
R548 B.n331 B.n249 585
R549 B.n334 B.n333 585
R550 B.n335 B.n245 585
R551 B.n337 B.n336 585
R552 B.n339 B.n244 585
R553 B.n342 B.n341 585
R554 B.n343 B.n243 585
R555 B.n345 B.n344 585
R556 B.n347 B.n242 585
R557 B.n350 B.n349 585
R558 B.n351 B.n241 585
R559 B.n353 B.n352 585
R560 B.n355 B.n240 585
R561 B.n358 B.n357 585
R562 B.n359 B.n239 585
R563 B.n361 B.n360 585
R564 B.n363 B.n238 585
R565 B.n366 B.n365 585
R566 B.n367 B.n237 585
R567 B.n369 B.n368 585
R568 B.n371 B.n236 585
R569 B.n372 B.n235 585
R570 B.n375 B.n374 585
R571 B.n376 B.n234 585
R572 B.n234 B.n233 585
R573 B.n381 B.n380 585
R574 B.n380 B.n379 585
R575 B.n382 B.n230 585
R576 B.n230 B.n229 585
R577 B.n384 B.n383 585
R578 B.n385 B.n384 585
R579 B.n224 B.n223 585
R580 B.n225 B.n224 585
R581 B.n393 B.n392 585
R582 B.n392 B.n391 585
R583 B.n394 B.n222 585
R584 B.n222 B.n221 585
R585 B.n396 B.n395 585
R586 B.n397 B.n396 585
R587 B.n216 B.n215 585
R588 B.n217 B.n216 585
R589 B.n405 B.n404 585
R590 B.n404 B.n403 585
R591 B.n406 B.n214 585
R592 B.n214 B.n213 585
R593 B.n408 B.n407 585
R594 B.n409 B.n408 585
R595 B.n208 B.n207 585
R596 B.n209 B.n208 585
R597 B.n418 B.n417 585
R598 B.n417 B.n416 585
R599 B.n419 B.n206 585
R600 B.n415 B.n206 585
R601 B.n421 B.n420 585
R602 B.n422 B.n421 585
R603 B.n201 B.n200 585
R604 B.n205 B.n201 585
R605 B.n430 B.n429 585
R606 B.n429 B.n428 585
R607 B.n431 B.n199 585
R608 B.n199 B.n198 585
R609 B.n433 B.n432 585
R610 B.n434 B.n433 585
R611 B.n193 B.n192 585
R612 B.n194 B.n193 585
R613 B.n444 B.n443 585
R614 B.n443 B.n442 585
R615 B.n445 B.n191 585
R616 B.n441 B.n191 585
R617 B.n447 B.n446 585
R618 B.n448 B.n447 585
R619 B.n2 B.n0 585
R620 B.n4 B.n2 585
R621 B.n3 B.n1 585
R622 B.n534 B.n3 585
R623 B.n532 B.n531 585
R624 B.n533 B.n532 585
R625 B.n530 B.n8 585
R626 B.n11 B.n8 585
R627 B.n529 B.n528 585
R628 B.n528 B.n527 585
R629 B.n10 B.n9 585
R630 B.n526 B.n10 585
R631 B.n524 B.n523 585
R632 B.n525 B.n524 585
R633 B.n522 B.n16 585
R634 B.n16 B.n15 585
R635 B.n521 B.n520 585
R636 B.n520 B.n519 585
R637 B.n18 B.n17 585
R638 B.n518 B.n18 585
R639 B.n516 B.n515 585
R640 B.n517 B.n516 585
R641 B.n514 B.n22 585
R642 B.n25 B.n22 585
R643 B.n513 B.n512 585
R644 B.n512 B.n511 585
R645 B.n24 B.n23 585
R646 B.n510 B.n24 585
R647 B.n508 B.n507 585
R648 B.n509 B.n508 585
R649 B.n506 B.n30 585
R650 B.n30 B.n29 585
R651 B.n505 B.n504 585
R652 B.n504 B.n503 585
R653 B.n32 B.n31 585
R654 B.n502 B.n32 585
R655 B.n500 B.n499 585
R656 B.n501 B.n500 585
R657 B.n498 B.n37 585
R658 B.n37 B.n36 585
R659 B.n497 B.n496 585
R660 B.n496 B.n495 585
R661 B.n39 B.n38 585
R662 B.n494 B.n39 585
R663 B.n492 B.n491 585
R664 B.n493 B.n492 585
R665 B.n490 B.n44 585
R666 B.n44 B.n43 585
R667 B.n489 B.n488 585
R668 B.n488 B.n487 585
R669 B.n537 B.n536 585
R670 B.n536 B.n535 585
R671 B.n380 B.n232 521.33
R672 B.n488 B.n46 521.33
R673 B.n378 B.n234 521.33
R674 B.n484 B.n47 521.33
R675 B.n246 B.t10 449.733
R676 B.n255 B.t18 449.733
R677 B.n78 B.t21 449.733
R678 B.n76 B.t14 449.733
R679 B.n486 B.n485 256.663
R680 B.n486 B.n74 256.663
R681 B.n486 B.n73 256.663
R682 B.n486 B.n72 256.663
R683 B.n486 B.n71 256.663
R684 B.n486 B.n70 256.663
R685 B.n486 B.n69 256.663
R686 B.n486 B.n68 256.663
R687 B.n486 B.n67 256.663
R688 B.n486 B.n66 256.663
R689 B.n486 B.n65 256.663
R690 B.n486 B.n64 256.663
R691 B.n486 B.n63 256.663
R692 B.n486 B.n62 256.663
R693 B.n486 B.n61 256.663
R694 B.n486 B.n60 256.663
R695 B.n486 B.n59 256.663
R696 B.n486 B.n58 256.663
R697 B.n486 B.n57 256.663
R698 B.n486 B.n56 256.663
R699 B.n486 B.n55 256.663
R700 B.n486 B.n54 256.663
R701 B.n486 B.n53 256.663
R702 B.n486 B.n52 256.663
R703 B.n486 B.n51 256.663
R704 B.n486 B.n50 256.663
R705 B.n486 B.n49 256.663
R706 B.n486 B.n48 256.663
R707 B.n267 B.n233 256.663
R708 B.n273 B.n233 256.663
R709 B.n275 B.n233 256.663
R710 B.n281 B.n233 256.663
R711 B.n283 B.n233 256.663
R712 B.n289 B.n233 256.663
R713 B.n291 B.n233 256.663
R714 B.n297 B.n233 256.663
R715 B.n299 B.n233 256.663
R716 B.n305 B.n233 256.663
R717 B.n307 B.n233 256.663
R718 B.n314 B.n233 256.663
R719 B.n316 B.n233 256.663
R720 B.n322 B.n233 256.663
R721 B.n324 B.n233 256.663
R722 B.n330 B.n233 256.663
R723 B.n332 B.n233 256.663
R724 B.n338 B.n233 256.663
R725 B.n340 B.n233 256.663
R726 B.n346 B.n233 256.663
R727 B.n348 B.n233 256.663
R728 B.n354 B.n233 256.663
R729 B.n356 B.n233 256.663
R730 B.n362 B.n233 256.663
R731 B.n364 B.n233 256.663
R732 B.n370 B.n233 256.663
R733 B.n373 B.n233 256.663
R734 B.n246 B.t13 192.369
R735 B.n76 B.t16 192.369
R736 B.n255 B.t20 192.369
R737 B.n78 B.t22 192.369
R738 B.n247 B.t12 174.913
R739 B.n77 B.t17 174.913
R740 B.n256 B.t19 174.913
R741 B.n79 B.t23 174.913
R742 B.n380 B.n230 163.367
R743 B.n384 B.n230 163.367
R744 B.n384 B.n224 163.367
R745 B.n392 B.n224 163.367
R746 B.n392 B.n222 163.367
R747 B.n396 B.n222 163.367
R748 B.n396 B.n216 163.367
R749 B.n404 B.n216 163.367
R750 B.n404 B.n214 163.367
R751 B.n408 B.n214 163.367
R752 B.n408 B.n208 163.367
R753 B.n417 B.n208 163.367
R754 B.n417 B.n206 163.367
R755 B.n421 B.n206 163.367
R756 B.n421 B.n201 163.367
R757 B.n429 B.n201 163.367
R758 B.n429 B.n199 163.367
R759 B.n433 B.n199 163.367
R760 B.n433 B.n193 163.367
R761 B.n443 B.n193 163.367
R762 B.n443 B.n191 163.367
R763 B.n447 B.n191 163.367
R764 B.n447 B.n2 163.367
R765 B.n536 B.n2 163.367
R766 B.n536 B.n3 163.367
R767 B.n532 B.n3 163.367
R768 B.n532 B.n8 163.367
R769 B.n528 B.n8 163.367
R770 B.n528 B.n10 163.367
R771 B.n524 B.n10 163.367
R772 B.n524 B.n16 163.367
R773 B.n520 B.n16 163.367
R774 B.n520 B.n18 163.367
R775 B.n516 B.n18 163.367
R776 B.n516 B.n22 163.367
R777 B.n512 B.n22 163.367
R778 B.n512 B.n24 163.367
R779 B.n508 B.n24 163.367
R780 B.n508 B.n30 163.367
R781 B.n504 B.n30 163.367
R782 B.n504 B.n32 163.367
R783 B.n500 B.n32 163.367
R784 B.n500 B.n37 163.367
R785 B.n496 B.n37 163.367
R786 B.n496 B.n39 163.367
R787 B.n492 B.n39 163.367
R788 B.n492 B.n44 163.367
R789 B.n488 B.n44 163.367
R790 B.n268 B.n266 163.367
R791 B.n272 B.n266 163.367
R792 B.n276 B.n274 163.367
R793 B.n280 B.n264 163.367
R794 B.n284 B.n282 163.367
R795 B.n288 B.n262 163.367
R796 B.n292 B.n290 163.367
R797 B.n296 B.n260 163.367
R798 B.n300 B.n298 163.367
R799 B.n304 B.n258 163.367
R800 B.n308 B.n306 163.367
R801 B.n313 B.n254 163.367
R802 B.n317 B.n315 163.367
R803 B.n321 B.n252 163.367
R804 B.n325 B.n323 163.367
R805 B.n329 B.n250 163.367
R806 B.n333 B.n331 163.367
R807 B.n337 B.n245 163.367
R808 B.n341 B.n339 163.367
R809 B.n345 B.n243 163.367
R810 B.n349 B.n347 163.367
R811 B.n353 B.n241 163.367
R812 B.n357 B.n355 163.367
R813 B.n361 B.n239 163.367
R814 B.n365 B.n363 163.367
R815 B.n369 B.n237 163.367
R816 B.n372 B.n371 163.367
R817 B.n374 B.n234 163.367
R818 B.n378 B.n228 163.367
R819 B.n386 B.n228 163.367
R820 B.n386 B.n226 163.367
R821 B.n390 B.n226 163.367
R822 B.n390 B.n220 163.367
R823 B.n398 B.n220 163.367
R824 B.n398 B.n218 163.367
R825 B.n402 B.n218 163.367
R826 B.n402 B.n212 163.367
R827 B.n410 B.n212 163.367
R828 B.n410 B.n210 163.367
R829 B.n414 B.n210 163.367
R830 B.n414 B.n204 163.367
R831 B.n423 B.n204 163.367
R832 B.n423 B.n202 163.367
R833 B.n427 B.n202 163.367
R834 B.n427 B.n197 163.367
R835 B.n435 B.n197 163.367
R836 B.n435 B.n195 163.367
R837 B.n440 B.n195 163.367
R838 B.n440 B.n190 163.367
R839 B.n449 B.n190 163.367
R840 B.n450 B.n449 163.367
R841 B.n450 B.n5 163.367
R842 B.n6 B.n5 163.367
R843 B.n7 B.n6 163.367
R844 B.n455 B.n7 163.367
R845 B.n455 B.n12 163.367
R846 B.n13 B.n12 163.367
R847 B.n14 B.n13 163.367
R848 B.n460 B.n14 163.367
R849 B.n460 B.n19 163.367
R850 B.n20 B.n19 163.367
R851 B.n21 B.n20 163.367
R852 B.n465 B.n21 163.367
R853 B.n465 B.n26 163.367
R854 B.n27 B.n26 163.367
R855 B.n28 B.n27 163.367
R856 B.n470 B.n28 163.367
R857 B.n470 B.n33 163.367
R858 B.n34 B.n33 163.367
R859 B.n35 B.n34 163.367
R860 B.n475 B.n35 163.367
R861 B.n475 B.n40 163.367
R862 B.n41 B.n40 163.367
R863 B.n42 B.n41 163.367
R864 B.n480 B.n42 163.367
R865 B.n480 B.n47 163.367
R866 B.n82 B.n81 163.367
R867 B.n86 B.n85 163.367
R868 B.n90 B.n89 163.367
R869 B.n94 B.n93 163.367
R870 B.n98 B.n97 163.367
R871 B.n102 B.n101 163.367
R872 B.n106 B.n105 163.367
R873 B.n110 B.n109 163.367
R874 B.n114 B.n113 163.367
R875 B.n118 B.n117 163.367
R876 B.n122 B.n121 163.367
R877 B.n127 B.n126 163.367
R878 B.n131 B.n130 163.367
R879 B.n135 B.n134 163.367
R880 B.n139 B.n138 163.367
R881 B.n143 B.n142 163.367
R882 B.n148 B.n147 163.367
R883 B.n152 B.n151 163.367
R884 B.n156 B.n155 163.367
R885 B.n160 B.n159 163.367
R886 B.n164 B.n163 163.367
R887 B.n168 B.n167 163.367
R888 B.n172 B.n171 163.367
R889 B.n176 B.n175 163.367
R890 B.n180 B.n179 163.367
R891 B.n184 B.n183 163.367
R892 B.n186 B.n75 163.367
R893 B.n379 B.n233 122.278
R894 B.n487 B.n486 122.278
R895 B.n267 B.n232 71.676
R896 B.n273 B.n272 71.676
R897 B.n276 B.n275 71.676
R898 B.n281 B.n280 71.676
R899 B.n284 B.n283 71.676
R900 B.n289 B.n288 71.676
R901 B.n292 B.n291 71.676
R902 B.n297 B.n296 71.676
R903 B.n300 B.n299 71.676
R904 B.n305 B.n304 71.676
R905 B.n308 B.n307 71.676
R906 B.n314 B.n313 71.676
R907 B.n317 B.n316 71.676
R908 B.n322 B.n321 71.676
R909 B.n325 B.n324 71.676
R910 B.n330 B.n329 71.676
R911 B.n333 B.n332 71.676
R912 B.n338 B.n337 71.676
R913 B.n341 B.n340 71.676
R914 B.n346 B.n345 71.676
R915 B.n349 B.n348 71.676
R916 B.n354 B.n353 71.676
R917 B.n357 B.n356 71.676
R918 B.n362 B.n361 71.676
R919 B.n365 B.n364 71.676
R920 B.n370 B.n369 71.676
R921 B.n373 B.n372 71.676
R922 B.n48 B.n46 71.676
R923 B.n82 B.n49 71.676
R924 B.n86 B.n50 71.676
R925 B.n90 B.n51 71.676
R926 B.n94 B.n52 71.676
R927 B.n98 B.n53 71.676
R928 B.n102 B.n54 71.676
R929 B.n106 B.n55 71.676
R930 B.n110 B.n56 71.676
R931 B.n114 B.n57 71.676
R932 B.n118 B.n58 71.676
R933 B.n122 B.n59 71.676
R934 B.n127 B.n60 71.676
R935 B.n131 B.n61 71.676
R936 B.n135 B.n62 71.676
R937 B.n139 B.n63 71.676
R938 B.n143 B.n64 71.676
R939 B.n148 B.n65 71.676
R940 B.n152 B.n66 71.676
R941 B.n156 B.n67 71.676
R942 B.n160 B.n68 71.676
R943 B.n164 B.n69 71.676
R944 B.n168 B.n70 71.676
R945 B.n172 B.n71 71.676
R946 B.n176 B.n72 71.676
R947 B.n180 B.n73 71.676
R948 B.n184 B.n74 71.676
R949 B.n485 B.n75 71.676
R950 B.n485 B.n484 71.676
R951 B.n186 B.n74 71.676
R952 B.n183 B.n73 71.676
R953 B.n179 B.n72 71.676
R954 B.n175 B.n71 71.676
R955 B.n171 B.n70 71.676
R956 B.n167 B.n69 71.676
R957 B.n163 B.n68 71.676
R958 B.n159 B.n67 71.676
R959 B.n155 B.n66 71.676
R960 B.n151 B.n65 71.676
R961 B.n147 B.n64 71.676
R962 B.n142 B.n63 71.676
R963 B.n138 B.n62 71.676
R964 B.n134 B.n61 71.676
R965 B.n130 B.n60 71.676
R966 B.n126 B.n59 71.676
R967 B.n121 B.n58 71.676
R968 B.n117 B.n57 71.676
R969 B.n113 B.n56 71.676
R970 B.n109 B.n55 71.676
R971 B.n105 B.n54 71.676
R972 B.n101 B.n53 71.676
R973 B.n97 B.n52 71.676
R974 B.n93 B.n51 71.676
R975 B.n89 B.n50 71.676
R976 B.n85 B.n49 71.676
R977 B.n81 B.n48 71.676
R978 B.n268 B.n267 71.676
R979 B.n274 B.n273 71.676
R980 B.n275 B.n264 71.676
R981 B.n282 B.n281 71.676
R982 B.n283 B.n262 71.676
R983 B.n290 B.n289 71.676
R984 B.n291 B.n260 71.676
R985 B.n298 B.n297 71.676
R986 B.n299 B.n258 71.676
R987 B.n306 B.n305 71.676
R988 B.n307 B.n254 71.676
R989 B.n315 B.n314 71.676
R990 B.n316 B.n252 71.676
R991 B.n323 B.n322 71.676
R992 B.n324 B.n250 71.676
R993 B.n331 B.n330 71.676
R994 B.n332 B.n245 71.676
R995 B.n339 B.n338 71.676
R996 B.n340 B.n243 71.676
R997 B.n347 B.n346 71.676
R998 B.n348 B.n241 71.676
R999 B.n355 B.n354 71.676
R1000 B.n356 B.n239 71.676
R1001 B.n363 B.n362 71.676
R1002 B.n364 B.n237 71.676
R1003 B.n371 B.n370 71.676
R1004 B.n374 B.n373 71.676
R1005 B.n379 B.n229 67.601
R1006 B.n385 B.n229 67.601
R1007 B.n385 B.n225 67.601
R1008 B.n391 B.n225 67.601
R1009 B.n397 B.n221 67.601
R1010 B.n397 B.n217 67.601
R1011 B.n403 B.n217 67.601
R1012 B.n403 B.n213 67.601
R1013 B.n409 B.n213 67.601
R1014 B.n416 B.n209 67.601
R1015 B.n416 B.n415 67.601
R1016 B.n422 B.n205 67.601
R1017 B.n428 B.n198 67.601
R1018 B.n434 B.n198 67.601
R1019 B.n442 B.n194 67.601
R1020 B.n442 B.n441 67.601
R1021 B.n448 B.n4 67.601
R1022 B.n535 B.n4 67.601
R1023 B.n535 B.n534 67.601
R1024 B.n534 B.n533 67.601
R1025 B.n527 B.n11 67.601
R1026 B.n527 B.n526 67.601
R1027 B.n525 B.n15 67.601
R1028 B.n519 B.n15 67.601
R1029 B.n518 B.n517 67.601
R1030 B.n511 B.n25 67.601
R1031 B.n511 B.n510 67.601
R1032 B.n509 B.n29 67.601
R1033 B.n503 B.n29 67.601
R1034 B.n503 B.n502 67.601
R1035 B.n502 B.n501 67.601
R1036 B.n501 B.n36 67.601
R1037 B.n495 B.n494 67.601
R1038 B.n494 B.n493 67.601
R1039 B.n493 B.n43 67.601
R1040 B.n487 B.n43 67.601
R1041 B.n448 B.t5 62.6304
R1042 B.n533 B.t0 62.6304
R1043 B.n248 B.n247 59.5399
R1044 B.n311 B.n256 59.5399
R1045 B.n124 B.n79 59.5399
R1046 B.n145 B.n77 59.5399
R1047 B.n422 B.t6 58.6539
R1048 B.n517 B.t2 58.6539
R1049 B.n205 B.t8 52.6892
R1050 B.t4 B.n518 52.6892
R1051 B.n391 B.t11 42.7479
R1052 B.n495 B.t15 42.7479
R1053 B.t7 B.n194 38.7714
R1054 B.n526 B.t9 38.7714
R1055 B.t3 B.n209 34.7949
R1056 B.n510 B.t1 34.7949
R1057 B.n489 B.n45 33.8737
R1058 B.n483 B.n482 33.8737
R1059 B.n377 B.n376 33.8737
R1060 B.n381 B.n231 33.8737
R1061 B.n409 B.t3 32.8066
R1062 B.t1 B.n509 32.8066
R1063 B.n434 B.t7 28.8301
R1064 B.t9 B.n525 28.8301
R1065 B.t11 B.n221 24.8536
R1066 B.t15 B.n36 24.8536
R1067 B B.n537 18.0485
R1068 B.n247 B.n246 17.455
R1069 B.n256 B.n255 17.455
R1070 B.n79 B.n78 17.455
R1071 B.n77 B.n76 17.455
R1072 B.n428 B.t8 14.9124
R1073 B.n519 B.t4 14.9124
R1074 B.n80 B.n45 10.6151
R1075 B.n83 B.n80 10.6151
R1076 B.n84 B.n83 10.6151
R1077 B.n87 B.n84 10.6151
R1078 B.n88 B.n87 10.6151
R1079 B.n91 B.n88 10.6151
R1080 B.n92 B.n91 10.6151
R1081 B.n95 B.n92 10.6151
R1082 B.n96 B.n95 10.6151
R1083 B.n99 B.n96 10.6151
R1084 B.n100 B.n99 10.6151
R1085 B.n103 B.n100 10.6151
R1086 B.n104 B.n103 10.6151
R1087 B.n107 B.n104 10.6151
R1088 B.n108 B.n107 10.6151
R1089 B.n111 B.n108 10.6151
R1090 B.n112 B.n111 10.6151
R1091 B.n115 B.n112 10.6151
R1092 B.n116 B.n115 10.6151
R1093 B.n119 B.n116 10.6151
R1094 B.n120 B.n119 10.6151
R1095 B.n123 B.n120 10.6151
R1096 B.n128 B.n125 10.6151
R1097 B.n129 B.n128 10.6151
R1098 B.n132 B.n129 10.6151
R1099 B.n133 B.n132 10.6151
R1100 B.n136 B.n133 10.6151
R1101 B.n137 B.n136 10.6151
R1102 B.n140 B.n137 10.6151
R1103 B.n141 B.n140 10.6151
R1104 B.n144 B.n141 10.6151
R1105 B.n149 B.n146 10.6151
R1106 B.n150 B.n149 10.6151
R1107 B.n153 B.n150 10.6151
R1108 B.n154 B.n153 10.6151
R1109 B.n157 B.n154 10.6151
R1110 B.n158 B.n157 10.6151
R1111 B.n161 B.n158 10.6151
R1112 B.n162 B.n161 10.6151
R1113 B.n165 B.n162 10.6151
R1114 B.n166 B.n165 10.6151
R1115 B.n169 B.n166 10.6151
R1116 B.n170 B.n169 10.6151
R1117 B.n173 B.n170 10.6151
R1118 B.n174 B.n173 10.6151
R1119 B.n177 B.n174 10.6151
R1120 B.n178 B.n177 10.6151
R1121 B.n181 B.n178 10.6151
R1122 B.n182 B.n181 10.6151
R1123 B.n185 B.n182 10.6151
R1124 B.n187 B.n185 10.6151
R1125 B.n188 B.n187 10.6151
R1126 B.n483 B.n188 10.6151
R1127 B.n377 B.n227 10.6151
R1128 B.n387 B.n227 10.6151
R1129 B.n388 B.n387 10.6151
R1130 B.n389 B.n388 10.6151
R1131 B.n389 B.n219 10.6151
R1132 B.n399 B.n219 10.6151
R1133 B.n400 B.n399 10.6151
R1134 B.n401 B.n400 10.6151
R1135 B.n401 B.n211 10.6151
R1136 B.n411 B.n211 10.6151
R1137 B.n412 B.n411 10.6151
R1138 B.n413 B.n412 10.6151
R1139 B.n413 B.n203 10.6151
R1140 B.n424 B.n203 10.6151
R1141 B.n425 B.n424 10.6151
R1142 B.n426 B.n425 10.6151
R1143 B.n426 B.n196 10.6151
R1144 B.n436 B.n196 10.6151
R1145 B.n437 B.n436 10.6151
R1146 B.n439 B.n437 10.6151
R1147 B.n439 B.n438 10.6151
R1148 B.n438 B.n189 10.6151
R1149 B.n451 B.n189 10.6151
R1150 B.n452 B.n451 10.6151
R1151 B.n453 B.n452 10.6151
R1152 B.n454 B.n453 10.6151
R1153 B.n456 B.n454 10.6151
R1154 B.n457 B.n456 10.6151
R1155 B.n458 B.n457 10.6151
R1156 B.n459 B.n458 10.6151
R1157 B.n461 B.n459 10.6151
R1158 B.n462 B.n461 10.6151
R1159 B.n463 B.n462 10.6151
R1160 B.n464 B.n463 10.6151
R1161 B.n466 B.n464 10.6151
R1162 B.n467 B.n466 10.6151
R1163 B.n468 B.n467 10.6151
R1164 B.n469 B.n468 10.6151
R1165 B.n471 B.n469 10.6151
R1166 B.n472 B.n471 10.6151
R1167 B.n473 B.n472 10.6151
R1168 B.n474 B.n473 10.6151
R1169 B.n476 B.n474 10.6151
R1170 B.n477 B.n476 10.6151
R1171 B.n478 B.n477 10.6151
R1172 B.n479 B.n478 10.6151
R1173 B.n481 B.n479 10.6151
R1174 B.n482 B.n481 10.6151
R1175 B.n269 B.n231 10.6151
R1176 B.n270 B.n269 10.6151
R1177 B.n271 B.n270 10.6151
R1178 B.n271 B.n265 10.6151
R1179 B.n277 B.n265 10.6151
R1180 B.n278 B.n277 10.6151
R1181 B.n279 B.n278 10.6151
R1182 B.n279 B.n263 10.6151
R1183 B.n285 B.n263 10.6151
R1184 B.n286 B.n285 10.6151
R1185 B.n287 B.n286 10.6151
R1186 B.n287 B.n261 10.6151
R1187 B.n293 B.n261 10.6151
R1188 B.n294 B.n293 10.6151
R1189 B.n295 B.n294 10.6151
R1190 B.n295 B.n259 10.6151
R1191 B.n301 B.n259 10.6151
R1192 B.n302 B.n301 10.6151
R1193 B.n303 B.n302 10.6151
R1194 B.n303 B.n257 10.6151
R1195 B.n309 B.n257 10.6151
R1196 B.n310 B.n309 10.6151
R1197 B.n312 B.n253 10.6151
R1198 B.n318 B.n253 10.6151
R1199 B.n319 B.n318 10.6151
R1200 B.n320 B.n319 10.6151
R1201 B.n320 B.n251 10.6151
R1202 B.n326 B.n251 10.6151
R1203 B.n327 B.n326 10.6151
R1204 B.n328 B.n327 10.6151
R1205 B.n328 B.n249 10.6151
R1206 B.n335 B.n334 10.6151
R1207 B.n336 B.n335 10.6151
R1208 B.n336 B.n244 10.6151
R1209 B.n342 B.n244 10.6151
R1210 B.n343 B.n342 10.6151
R1211 B.n344 B.n343 10.6151
R1212 B.n344 B.n242 10.6151
R1213 B.n350 B.n242 10.6151
R1214 B.n351 B.n350 10.6151
R1215 B.n352 B.n351 10.6151
R1216 B.n352 B.n240 10.6151
R1217 B.n358 B.n240 10.6151
R1218 B.n359 B.n358 10.6151
R1219 B.n360 B.n359 10.6151
R1220 B.n360 B.n238 10.6151
R1221 B.n366 B.n238 10.6151
R1222 B.n367 B.n366 10.6151
R1223 B.n368 B.n367 10.6151
R1224 B.n368 B.n236 10.6151
R1225 B.n236 B.n235 10.6151
R1226 B.n375 B.n235 10.6151
R1227 B.n376 B.n375 10.6151
R1228 B.n382 B.n381 10.6151
R1229 B.n383 B.n382 10.6151
R1230 B.n383 B.n223 10.6151
R1231 B.n393 B.n223 10.6151
R1232 B.n394 B.n393 10.6151
R1233 B.n395 B.n394 10.6151
R1234 B.n395 B.n215 10.6151
R1235 B.n405 B.n215 10.6151
R1236 B.n406 B.n405 10.6151
R1237 B.n407 B.n406 10.6151
R1238 B.n407 B.n207 10.6151
R1239 B.n418 B.n207 10.6151
R1240 B.n419 B.n418 10.6151
R1241 B.n420 B.n419 10.6151
R1242 B.n420 B.n200 10.6151
R1243 B.n430 B.n200 10.6151
R1244 B.n431 B.n430 10.6151
R1245 B.n432 B.n431 10.6151
R1246 B.n432 B.n192 10.6151
R1247 B.n444 B.n192 10.6151
R1248 B.n445 B.n444 10.6151
R1249 B.n446 B.n445 10.6151
R1250 B.n446 B.n0 10.6151
R1251 B.n531 B.n1 10.6151
R1252 B.n531 B.n530 10.6151
R1253 B.n530 B.n529 10.6151
R1254 B.n529 B.n9 10.6151
R1255 B.n523 B.n9 10.6151
R1256 B.n523 B.n522 10.6151
R1257 B.n522 B.n521 10.6151
R1258 B.n521 B.n17 10.6151
R1259 B.n515 B.n17 10.6151
R1260 B.n515 B.n514 10.6151
R1261 B.n514 B.n513 10.6151
R1262 B.n513 B.n23 10.6151
R1263 B.n507 B.n23 10.6151
R1264 B.n507 B.n506 10.6151
R1265 B.n506 B.n505 10.6151
R1266 B.n505 B.n31 10.6151
R1267 B.n499 B.n31 10.6151
R1268 B.n499 B.n498 10.6151
R1269 B.n498 B.n497 10.6151
R1270 B.n497 B.n38 10.6151
R1271 B.n491 B.n38 10.6151
R1272 B.n491 B.n490 10.6151
R1273 B.n490 B.n489 10.6151
R1274 B.n124 B.n123 9.36635
R1275 B.n146 B.n145 9.36635
R1276 B.n311 B.n310 9.36635
R1277 B.n334 B.n248 9.36635
R1278 B.n415 B.t6 8.94763
R1279 B.n25 B.t2 8.94763
R1280 B.n441 B.t5 4.97113
R1281 B.n11 B.t0 4.97113
R1282 B.n537 B.n0 2.81026
R1283 B.n537 B.n1 2.81026
R1284 B.n125 B.n124 1.24928
R1285 B.n145 B.n144 1.24928
R1286 B.n312 B.n311 1.24928
R1287 B.n249 B.n248 1.24928
R1288 VP.n6 VP.t7 338.866
R1289 VP.n14 VP.t9 314.147
R1290 VP.n16 VP.t6 314.147
R1291 VP.n1 VP.t8 314.147
R1292 VP.n20 VP.t3 314.147
R1293 VP.n22 VP.t1 314.147
R1294 VP.n11 VP.t0 314.147
R1295 VP.n9 VP.t2 314.147
R1296 VP.n8 VP.t4 314.147
R1297 VP.n7 VP.t5 314.147
R1298 VP.n23 VP.n22 161.3
R1299 VP.n9 VP.n4 161.3
R1300 VP.n10 VP.n3 161.3
R1301 VP.n12 VP.n11 161.3
R1302 VP.n21 VP.n0 161.3
R1303 VP.n20 VP.n19 161.3
R1304 VP.n17 VP.n16 161.3
R1305 VP.n15 VP.n2 161.3
R1306 VP.n14 VP.n13 161.3
R1307 VP.n8 VP.n5 80.6037
R1308 VP.n18 VP.n1 80.6037
R1309 VP.n16 VP.n1 48.2005
R1310 VP.n20 VP.n1 48.2005
R1311 VP.n9 VP.n8 48.2005
R1312 VP.n8 VP.n7 48.2005
R1313 VP.n6 VP.n5 45.0526
R1314 VP.n15 VP.n14 38.7066
R1315 VP.n22 VP.n21 38.7066
R1316 VP.n11 VP.n10 38.7066
R1317 VP.n13 VP.n12 37.3338
R1318 VP.n7 VP.n6 16.5858
R1319 VP.n16 VP.n15 9.49444
R1320 VP.n21 VP.n20 9.49444
R1321 VP.n10 VP.n9 9.49444
R1322 VP.n5 VP.n4 0.285035
R1323 VP.n18 VP.n17 0.285035
R1324 VP.n19 VP.n18 0.285035
R1325 VP.n4 VP.n3 0.189894
R1326 VP.n12 VP.n3 0.189894
R1327 VP.n13 VP.n2 0.189894
R1328 VP.n17 VP.n2 0.189894
R1329 VP.n19 VP.n0 0.189894
R1330 VP.n23 VP.n0 0.189894
R1331 VP VP.n23 0.0516364
R1332 VDD1.n28 VDD1.n27 289.615
R1333 VDD1.n59 VDD1.n58 289.615
R1334 VDD1.n27 VDD1.n26 185
R1335 VDD1.n2 VDD1.n1 185
R1336 VDD1.n21 VDD1.n20 185
R1337 VDD1.n19 VDD1.n18 185
R1338 VDD1.n6 VDD1.n5 185
R1339 VDD1.n13 VDD1.n12 185
R1340 VDD1.n11 VDD1.n10 185
R1341 VDD1.n42 VDD1.n41 185
R1342 VDD1.n44 VDD1.n43 185
R1343 VDD1.n37 VDD1.n36 185
R1344 VDD1.n50 VDD1.n49 185
R1345 VDD1.n52 VDD1.n51 185
R1346 VDD1.n33 VDD1.n32 185
R1347 VDD1.n58 VDD1.n57 185
R1348 VDD1.n9 VDD1.t2 149.528
R1349 VDD1.n40 VDD1.t0 149.528
R1350 VDD1.n27 VDD1.n1 104.615
R1351 VDD1.n20 VDD1.n1 104.615
R1352 VDD1.n20 VDD1.n19 104.615
R1353 VDD1.n19 VDD1.n5 104.615
R1354 VDD1.n12 VDD1.n5 104.615
R1355 VDD1.n12 VDD1.n11 104.615
R1356 VDD1.n43 VDD1.n42 104.615
R1357 VDD1.n43 VDD1.n36 104.615
R1358 VDD1.n50 VDD1.n36 104.615
R1359 VDD1.n51 VDD1.n50 104.615
R1360 VDD1.n51 VDD1.n32 104.615
R1361 VDD1.n58 VDD1.n32 104.615
R1362 VDD1.n63 VDD1.n62 69.8098
R1363 VDD1.n30 VDD1.n29 69.2843
R1364 VDD1.n61 VDD1.n60 69.2833
R1365 VDD1.n65 VDD1.n64 69.2831
R1366 VDD1.n11 VDD1.t2 52.3082
R1367 VDD1.n42 VDD1.t0 52.3082
R1368 VDD1.n30 VDD1.n28 51.3855
R1369 VDD1.n61 VDD1.n59 51.3855
R1370 VDD1.n65 VDD1.n63 33.363
R1371 VDD1.n26 VDD1.n0 12.0247
R1372 VDD1.n57 VDD1.n31 12.0247
R1373 VDD1.n25 VDD1.n2 11.249
R1374 VDD1.n56 VDD1.n33 11.249
R1375 VDD1.n22 VDD1.n21 10.4732
R1376 VDD1.n53 VDD1.n52 10.4732
R1377 VDD1.n10 VDD1.n9 10.2745
R1378 VDD1.n41 VDD1.n40 10.2745
R1379 VDD1.n18 VDD1.n4 9.69747
R1380 VDD1.n49 VDD1.n35 9.69747
R1381 VDD1.n24 VDD1.n0 9.45567
R1382 VDD1.n55 VDD1.n31 9.45567
R1383 VDD1.n15 VDD1.n14 9.3005
R1384 VDD1.n17 VDD1.n16 9.3005
R1385 VDD1.n4 VDD1.n3 9.3005
R1386 VDD1.n23 VDD1.n22 9.3005
R1387 VDD1.n25 VDD1.n24 9.3005
R1388 VDD1.n8 VDD1.n7 9.3005
R1389 VDD1.n39 VDD1.n38 9.3005
R1390 VDD1.n46 VDD1.n45 9.3005
R1391 VDD1.n48 VDD1.n47 9.3005
R1392 VDD1.n35 VDD1.n34 9.3005
R1393 VDD1.n54 VDD1.n53 9.3005
R1394 VDD1.n56 VDD1.n55 9.3005
R1395 VDD1.n17 VDD1.n6 8.92171
R1396 VDD1.n48 VDD1.n37 8.92171
R1397 VDD1.n14 VDD1.n13 8.14595
R1398 VDD1.n45 VDD1.n44 8.14595
R1399 VDD1.n10 VDD1.n8 7.3702
R1400 VDD1.n41 VDD1.n39 7.3702
R1401 VDD1.n13 VDD1.n8 5.81868
R1402 VDD1.n44 VDD1.n39 5.81868
R1403 VDD1.n14 VDD1.n6 5.04292
R1404 VDD1.n45 VDD1.n37 5.04292
R1405 VDD1.n18 VDD1.n17 4.26717
R1406 VDD1.n49 VDD1.n48 4.26717
R1407 VDD1.n21 VDD1.n4 3.49141
R1408 VDD1.n52 VDD1.n35 3.49141
R1409 VDD1.n64 VDD1.t7 3.42019
R1410 VDD1.n64 VDD1.t9 3.42019
R1411 VDD1.n29 VDD1.t4 3.42019
R1412 VDD1.n29 VDD1.t5 3.42019
R1413 VDD1.n62 VDD1.t6 3.42019
R1414 VDD1.n62 VDD1.t8 3.42019
R1415 VDD1.n60 VDD1.t3 3.42019
R1416 VDD1.n60 VDD1.t1 3.42019
R1417 VDD1.n9 VDD1.n7 2.84323
R1418 VDD1.n40 VDD1.n38 2.84323
R1419 VDD1.n22 VDD1.n2 2.71565
R1420 VDD1.n53 VDD1.n33 2.71565
R1421 VDD1.n26 VDD1.n25 1.93989
R1422 VDD1.n57 VDD1.n56 1.93989
R1423 VDD1.n28 VDD1.n0 1.16414
R1424 VDD1.n59 VDD1.n31 1.16414
R1425 VDD1 VDD1.n65 0.524207
R1426 VDD1 VDD1.n30 0.252655
R1427 VDD1.n24 VDD1.n23 0.155672
R1428 VDD1.n23 VDD1.n3 0.155672
R1429 VDD1.n16 VDD1.n3 0.155672
R1430 VDD1.n16 VDD1.n15 0.155672
R1431 VDD1.n15 VDD1.n7 0.155672
R1432 VDD1.n46 VDD1.n38 0.155672
R1433 VDD1.n47 VDD1.n46 0.155672
R1434 VDD1.n47 VDD1.n34 0.155672
R1435 VDD1.n54 VDD1.n34 0.155672
R1436 VDD1.n55 VDD1.n54 0.155672
R1437 VDD1.n63 VDD1.n61 0.139119
C0 VP VN 4.25878f
C1 VTAIL VDD2 8.7807f
C2 VTAIL VDD1 8.7442f
C3 VDD2 VP 0.324066f
C4 VP VDD1 3.27018f
C5 VTAIL VP 3.18588f
C6 VDD2 VN 3.09742f
C7 VDD1 VN 0.148722f
C8 VDD2 VDD1 0.889709f
C9 VTAIL VN 3.17151f
C10 VDD2 B 3.705568f
C11 VDD1 B 3.630112f
C12 VTAIL B 4.017012f
C13 VN B 8.09712f
C14 VP B 6.376791f
C15 VDD1.n0 B 0.014319f
C16 VDD1.n1 B 0.032323f
C17 VDD1.n2 B 0.01448f
C18 VDD1.n3 B 0.025449f
C19 VDD1.n4 B 0.013675f
C20 VDD1.n5 B 0.032323f
C21 VDD1.n6 B 0.01448f
C22 VDD1.n7 B 0.580584f
C23 VDD1.n8 B 0.013675f
C24 VDD1.t2 B 0.053863f
C25 VDD1.n9 B 0.123029f
C26 VDD1.n10 B 0.022849f
C27 VDD1.n11 B 0.024242f
C28 VDD1.n12 B 0.032323f
C29 VDD1.n13 B 0.01448f
C30 VDD1.n14 B 0.013675f
C31 VDD1.n15 B 0.025449f
C32 VDD1.n16 B 0.025449f
C33 VDD1.n17 B 0.013675f
C34 VDD1.n18 B 0.01448f
C35 VDD1.n19 B 0.032323f
C36 VDD1.n20 B 0.032323f
C37 VDD1.n21 B 0.01448f
C38 VDD1.n22 B 0.013675f
C39 VDD1.n23 B 0.025449f
C40 VDD1.n24 B 0.064039f
C41 VDD1.n25 B 0.013675f
C42 VDD1.n26 B 0.01448f
C43 VDD1.n27 B 0.063598f
C44 VDD1.n28 B 0.072583f
C45 VDD1.t4 B 0.11644f
C46 VDD1.t5 B 0.11644f
C47 VDD1.n29 B 0.977655f
C48 VDD1.n30 B 0.392033f
C49 VDD1.n31 B 0.014319f
C50 VDD1.n32 B 0.032323f
C51 VDD1.n33 B 0.01448f
C52 VDD1.n34 B 0.025449f
C53 VDD1.n35 B 0.013675f
C54 VDD1.n36 B 0.032323f
C55 VDD1.n37 B 0.01448f
C56 VDD1.n38 B 0.580584f
C57 VDD1.n39 B 0.013675f
C58 VDD1.t0 B 0.053863f
C59 VDD1.n40 B 0.123029f
C60 VDD1.n41 B 0.022849f
C61 VDD1.n42 B 0.024242f
C62 VDD1.n43 B 0.032323f
C63 VDD1.n44 B 0.01448f
C64 VDD1.n45 B 0.013675f
C65 VDD1.n46 B 0.025449f
C66 VDD1.n47 B 0.025449f
C67 VDD1.n48 B 0.013675f
C68 VDD1.n49 B 0.01448f
C69 VDD1.n50 B 0.032323f
C70 VDD1.n51 B 0.032323f
C71 VDD1.n52 B 0.01448f
C72 VDD1.n53 B 0.013675f
C73 VDD1.n54 B 0.025449f
C74 VDD1.n55 B 0.064039f
C75 VDD1.n56 B 0.013675f
C76 VDD1.n57 B 0.01448f
C77 VDD1.n58 B 0.063598f
C78 VDD1.n59 B 0.072583f
C79 VDD1.t3 B 0.11644f
C80 VDD1.t1 B 0.11644f
C81 VDD1.n60 B 0.977657f
C82 VDD1.n61 B 0.386977f
C83 VDD1.t6 B 0.11644f
C84 VDD1.t8 B 0.11644f
C85 VDD1.n62 B 0.980019f
C86 VDD1.n63 B 1.55025f
C87 VDD1.t7 B 0.11644f
C88 VDD1.t9 B 0.11644f
C89 VDD1.n64 B 0.977653f
C90 VDD1.n65 B 1.85972f
C91 VP.n0 B 0.047993f
C92 VP.t8 B 0.460238f
C93 VP.n1 B 0.228518f
C94 VP.n2 B 0.047993f
C95 VP.n3 B 0.047993f
C96 VP.t0 B 0.460238f
C97 VP.t2 B 0.460238f
C98 VP.n4 B 0.06404f
C99 VP.t4 B 0.460238f
C100 VP.n5 B 0.227579f
C101 VP.t5 B 0.460238f
C102 VP.t7 B 0.476069f
C103 VP.n6 B 0.205103f
C104 VP.n7 B 0.226578f
C105 VP.n8 B 0.228518f
C106 VP.n9 B 0.219551f
C107 VP.n10 B 0.010891f
C108 VP.n11 B 0.215704f
C109 VP.n12 B 1.61392f
C110 VP.n13 B 1.66013f
C111 VP.t9 B 0.460238f
C112 VP.n14 B 0.215704f
C113 VP.n15 B 0.010891f
C114 VP.t6 B 0.460238f
C115 VP.n16 B 0.219551f
C116 VP.n17 B 0.06404f
C117 VP.n18 B 0.06389f
C118 VP.n19 B 0.06404f
C119 VP.t3 B 0.460238f
C120 VP.n20 B 0.219551f
C121 VP.n21 B 0.010891f
C122 VP.t1 B 0.460238f
C123 VP.n22 B 0.215704f
C124 VP.n23 B 0.037193f
C125 VDD2.n0 B 0.014312f
C126 VDD2.n1 B 0.032307f
C127 VDD2.n2 B 0.014472f
C128 VDD2.n3 B 0.025436f
C129 VDD2.n4 B 0.013668f
C130 VDD2.n5 B 0.032307f
C131 VDD2.n6 B 0.014472f
C132 VDD2.n7 B 0.580291f
C133 VDD2.n8 B 0.013668f
C134 VDD2.t0 B 0.053836f
C135 VDD2.n9 B 0.122967f
C136 VDD2.n10 B 0.022837f
C137 VDD2.n11 B 0.02423f
C138 VDD2.n12 B 0.032307f
C139 VDD2.n13 B 0.014472f
C140 VDD2.n14 B 0.013668f
C141 VDD2.n15 B 0.025436f
C142 VDD2.n16 B 0.025436f
C143 VDD2.n17 B 0.013668f
C144 VDD2.n18 B 0.014472f
C145 VDD2.n19 B 0.032307f
C146 VDD2.n20 B 0.032307f
C147 VDD2.n21 B 0.014472f
C148 VDD2.n22 B 0.013668f
C149 VDD2.n23 B 0.025436f
C150 VDD2.n24 B 0.064006f
C151 VDD2.n25 B 0.013668f
C152 VDD2.n26 B 0.014472f
C153 VDD2.n27 B 0.063566f
C154 VDD2.n28 B 0.072546f
C155 VDD2.t7 B 0.116381f
C156 VDD2.t5 B 0.116381f
C157 VDD2.n29 B 0.977164f
C158 VDD2.n30 B 0.386782f
C159 VDD2.t6 B 0.116381f
C160 VDD2.t1 B 0.116381f
C161 VDD2.n31 B 0.979525f
C162 VDD2.n32 B 1.4765f
C163 VDD2.n33 B 0.014312f
C164 VDD2.n34 B 0.032307f
C165 VDD2.n35 B 0.014472f
C166 VDD2.n36 B 0.025436f
C167 VDD2.n37 B 0.013668f
C168 VDD2.n38 B 0.032307f
C169 VDD2.n39 B 0.014472f
C170 VDD2.n40 B 0.580291f
C171 VDD2.n41 B 0.013668f
C172 VDD2.t9 B 0.053836f
C173 VDD2.n42 B 0.122967f
C174 VDD2.n43 B 0.022837f
C175 VDD2.n44 B 0.02423f
C176 VDD2.n45 B 0.032307f
C177 VDD2.n46 B 0.014472f
C178 VDD2.n47 B 0.013668f
C179 VDD2.n48 B 0.025436f
C180 VDD2.n49 B 0.025436f
C181 VDD2.n50 B 0.013668f
C182 VDD2.n51 B 0.014472f
C183 VDD2.n52 B 0.032307f
C184 VDD2.n53 B 0.032307f
C185 VDD2.n54 B 0.014472f
C186 VDD2.n55 B 0.013668f
C187 VDD2.n56 B 0.025436f
C188 VDD2.n57 B 0.064006f
C189 VDD2.n58 B 0.013668f
C190 VDD2.n59 B 0.014472f
C191 VDD2.n60 B 0.063566f
C192 VDD2.n61 B 0.07082f
C193 VDD2.n62 B 1.64046f
C194 VDD2.t8 B 0.116381f
C195 VDD2.t4 B 0.116381f
C196 VDD2.n63 B 0.977162f
C197 VDD2.n64 B 0.279202f
C198 VDD2.t3 B 0.116381f
C199 VDD2.t2 B 0.116381f
C200 VDD2.n65 B 0.979498f
C201 VTAIL.t15 B 0.129488f
C202 VTAIL.t10 B 0.129488f
C203 VTAIL.n0 B 1.02015f
C204 VTAIL.n1 B 0.382085f
C205 VTAIL.n2 B 0.015924f
C206 VTAIL.n3 B 0.035945f
C207 VTAIL.n4 B 0.016102f
C208 VTAIL.n5 B 0.028301f
C209 VTAIL.n6 B 0.015208f
C210 VTAIL.n7 B 0.035945f
C211 VTAIL.n8 B 0.016102f
C212 VTAIL.n9 B 0.645644f
C213 VTAIL.n10 B 0.015208f
C214 VTAIL.t5 B 0.059899f
C215 VTAIL.n11 B 0.136816f
C216 VTAIL.n12 B 0.025409f
C217 VTAIL.n13 B 0.026959f
C218 VTAIL.n14 B 0.035945f
C219 VTAIL.n15 B 0.016102f
C220 VTAIL.n16 B 0.015208f
C221 VTAIL.n17 B 0.028301f
C222 VTAIL.n18 B 0.028301f
C223 VTAIL.n19 B 0.015208f
C224 VTAIL.n20 B 0.016102f
C225 VTAIL.n21 B 0.035945f
C226 VTAIL.n22 B 0.035945f
C227 VTAIL.n23 B 0.016102f
C228 VTAIL.n24 B 0.015208f
C229 VTAIL.n25 B 0.028301f
C230 VTAIL.n26 B 0.071215f
C231 VTAIL.n27 B 0.015208f
C232 VTAIL.n28 B 0.016102f
C233 VTAIL.n29 B 0.070724f
C234 VTAIL.n30 B 0.05928f
C235 VTAIL.n31 B 0.175109f
C236 VTAIL.t19 B 0.129488f
C237 VTAIL.t7 B 0.129488f
C238 VTAIL.n32 B 1.02015f
C239 VTAIL.n33 B 0.386998f
C240 VTAIL.t3 B 0.129488f
C241 VTAIL.t6 B 0.129488f
C242 VTAIL.n34 B 1.02015f
C243 VTAIL.n35 B 1.29735f
C244 VTAIL.t12 B 0.129488f
C245 VTAIL.t11 B 0.129488f
C246 VTAIL.n36 B 1.02015f
C247 VTAIL.n37 B 1.29735f
C248 VTAIL.t16 B 0.129488f
C249 VTAIL.t17 B 0.129488f
C250 VTAIL.n38 B 1.02015f
C251 VTAIL.n39 B 0.386999f
C252 VTAIL.n40 B 0.015924f
C253 VTAIL.n41 B 0.035945f
C254 VTAIL.n42 B 0.016102f
C255 VTAIL.n43 B 0.028301f
C256 VTAIL.n44 B 0.015208f
C257 VTAIL.n45 B 0.035945f
C258 VTAIL.n46 B 0.016102f
C259 VTAIL.n47 B 0.645644f
C260 VTAIL.n48 B 0.015208f
C261 VTAIL.t14 B 0.059899f
C262 VTAIL.n49 B 0.136816f
C263 VTAIL.n50 B 0.025409f
C264 VTAIL.n51 B 0.026959f
C265 VTAIL.n52 B 0.035945f
C266 VTAIL.n53 B 0.016102f
C267 VTAIL.n54 B 0.015208f
C268 VTAIL.n55 B 0.028301f
C269 VTAIL.n56 B 0.028301f
C270 VTAIL.n57 B 0.015208f
C271 VTAIL.n58 B 0.016102f
C272 VTAIL.n59 B 0.035945f
C273 VTAIL.n60 B 0.035945f
C274 VTAIL.n61 B 0.016102f
C275 VTAIL.n62 B 0.015208f
C276 VTAIL.n63 B 0.028301f
C277 VTAIL.n64 B 0.071215f
C278 VTAIL.n65 B 0.015208f
C279 VTAIL.n66 B 0.016102f
C280 VTAIL.n67 B 0.070724f
C281 VTAIL.n68 B 0.05928f
C282 VTAIL.n69 B 0.175109f
C283 VTAIL.t0 B 0.129488f
C284 VTAIL.t18 B 0.129488f
C285 VTAIL.n70 B 1.02015f
C286 VTAIL.n71 B 0.394467f
C287 VTAIL.t4 B 0.129488f
C288 VTAIL.t2 B 0.129488f
C289 VTAIL.n72 B 1.02015f
C290 VTAIL.n73 B 0.386999f
C291 VTAIL.n74 B 0.015924f
C292 VTAIL.n75 B 0.035945f
C293 VTAIL.n76 B 0.016102f
C294 VTAIL.n77 B 0.028301f
C295 VTAIL.n78 B 0.015208f
C296 VTAIL.n79 B 0.035945f
C297 VTAIL.n80 B 0.016102f
C298 VTAIL.n81 B 0.645644f
C299 VTAIL.n82 B 0.015208f
C300 VTAIL.t1 B 0.059899f
C301 VTAIL.n83 B 0.136816f
C302 VTAIL.n84 B 0.025409f
C303 VTAIL.n85 B 0.026959f
C304 VTAIL.n86 B 0.035945f
C305 VTAIL.n87 B 0.016102f
C306 VTAIL.n88 B 0.015208f
C307 VTAIL.n89 B 0.028301f
C308 VTAIL.n90 B 0.028301f
C309 VTAIL.n91 B 0.015208f
C310 VTAIL.n92 B 0.016102f
C311 VTAIL.n93 B 0.035945f
C312 VTAIL.n94 B 0.035945f
C313 VTAIL.n95 B 0.016102f
C314 VTAIL.n96 B 0.015208f
C315 VTAIL.n97 B 0.028301f
C316 VTAIL.n98 B 0.071215f
C317 VTAIL.n99 B 0.015208f
C318 VTAIL.n100 B 0.016102f
C319 VTAIL.n101 B 0.070724f
C320 VTAIL.n102 B 0.05928f
C321 VTAIL.n103 B 1.00724f
C322 VTAIL.n104 B 0.015924f
C323 VTAIL.n105 B 0.035945f
C324 VTAIL.n106 B 0.016102f
C325 VTAIL.n107 B 0.028301f
C326 VTAIL.n108 B 0.015208f
C327 VTAIL.n109 B 0.035945f
C328 VTAIL.n110 B 0.016102f
C329 VTAIL.n111 B 0.645644f
C330 VTAIL.n112 B 0.015208f
C331 VTAIL.t8 B 0.059899f
C332 VTAIL.n113 B 0.136816f
C333 VTAIL.n114 B 0.025409f
C334 VTAIL.n115 B 0.026959f
C335 VTAIL.n116 B 0.035945f
C336 VTAIL.n117 B 0.016102f
C337 VTAIL.n118 B 0.015208f
C338 VTAIL.n119 B 0.028301f
C339 VTAIL.n120 B 0.028301f
C340 VTAIL.n121 B 0.015208f
C341 VTAIL.n122 B 0.016102f
C342 VTAIL.n123 B 0.035945f
C343 VTAIL.n124 B 0.035945f
C344 VTAIL.n125 B 0.016102f
C345 VTAIL.n126 B 0.015208f
C346 VTAIL.n127 B 0.028301f
C347 VTAIL.n128 B 0.071215f
C348 VTAIL.n129 B 0.015208f
C349 VTAIL.n130 B 0.016102f
C350 VTAIL.n131 B 0.070724f
C351 VTAIL.n132 B 0.05928f
C352 VTAIL.n133 B 1.00724f
C353 VTAIL.t13 B 0.129488f
C354 VTAIL.t9 B 0.129488f
C355 VTAIL.n134 B 1.02015f
C356 VTAIL.n135 B 0.328628f
C357 VN.n0 B 0.046812f
C358 VN.t4 B 0.448911f
C359 VN.n1 B 0.222894f
C360 VN.t9 B 0.464352f
C361 VN.t2 B 0.448911f
C362 VN.n2 B 0.221002f
C363 VN.n3 B 0.200056f
C364 VN.n4 B 0.221978f
C365 VN.n5 B 0.062464f
C366 VN.t3 B 0.448911f
C367 VN.n6 B 0.214147f
C368 VN.n7 B 0.010623f
C369 VN.t8 B 0.448911f
C370 VN.n8 B 0.210395f
C371 VN.n9 B 0.036277f
C372 VN.n10 B 0.046812f
C373 VN.t5 B 0.448911f
C374 VN.n11 B 0.222894f
C375 VN.t1 B 0.448911f
C376 VN.t7 B 0.464352f
C377 VN.t6 B 0.448911f
C378 VN.n12 B 0.221002f
C379 VN.n13 B 0.200056f
C380 VN.n14 B 0.221978f
C381 VN.n15 B 0.062464f
C382 VN.n16 B 0.214147f
C383 VN.n17 B 0.010623f
C384 VN.t0 B 0.448911f
C385 VN.n18 B 0.210395f
C386 VN.n19 B 1.60517f
.ends

