* NGSPICE file created from diff_pair_sample_1328.ext - technology: sky130A

.subckt diff_pair_sample_1328 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t5 VP.t0 VTAIL.t8 w_n1410_n4554# sky130_fd_pr__pfet_01v8 ad=6.9927 pd=36.64 as=2.95845 ps=18.26 w=17.93 l=0.22
X1 VDD2.t5 VN.t0 VTAIL.t5 w_n1410_n4554# sky130_fd_pr__pfet_01v8 ad=6.9927 pd=36.64 as=2.95845 ps=18.26 w=17.93 l=0.22
X2 B.t11 B.t9 B.t10 w_n1410_n4554# sky130_fd_pr__pfet_01v8 ad=6.9927 pd=36.64 as=0 ps=0 w=17.93 l=0.22
X3 VDD1.t4 VP.t1 VTAIL.t10 w_n1410_n4554# sky130_fd_pr__pfet_01v8 ad=2.95845 pd=18.26 as=6.9927 ps=36.64 w=17.93 l=0.22
X4 B.t8 B.t6 B.t7 w_n1410_n4554# sky130_fd_pr__pfet_01v8 ad=6.9927 pd=36.64 as=0 ps=0 w=17.93 l=0.22
X5 VDD1.t3 VP.t2 VTAIL.t11 w_n1410_n4554# sky130_fd_pr__pfet_01v8 ad=6.9927 pd=36.64 as=2.95845 ps=18.26 w=17.93 l=0.22
X6 VDD2.t4 VN.t1 VTAIL.t4 w_n1410_n4554# sky130_fd_pr__pfet_01v8 ad=6.9927 pd=36.64 as=2.95845 ps=18.26 w=17.93 l=0.22
X7 B.t5 B.t3 B.t4 w_n1410_n4554# sky130_fd_pr__pfet_01v8 ad=6.9927 pd=36.64 as=0 ps=0 w=17.93 l=0.22
X8 VDD2.t3 VN.t2 VTAIL.t0 w_n1410_n4554# sky130_fd_pr__pfet_01v8 ad=2.95845 pd=18.26 as=6.9927 ps=36.64 w=17.93 l=0.22
X9 VTAIL.t9 VP.t3 VDD1.t2 w_n1410_n4554# sky130_fd_pr__pfet_01v8 ad=2.95845 pd=18.26 as=2.95845 ps=18.26 w=17.93 l=0.22
X10 VTAIL.t6 VP.t4 VDD1.t1 w_n1410_n4554# sky130_fd_pr__pfet_01v8 ad=2.95845 pd=18.26 as=2.95845 ps=18.26 w=17.93 l=0.22
X11 VDD2.t2 VN.t3 VTAIL.t1 w_n1410_n4554# sky130_fd_pr__pfet_01v8 ad=2.95845 pd=18.26 as=6.9927 ps=36.64 w=17.93 l=0.22
X12 VTAIL.t2 VN.t4 VDD2.t1 w_n1410_n4554# sky130_fd_pr__pfet_01v8 ad=2.95845 pd=18.26 as=2.95845 ps=18.26 w=17.93 l=0.22
X13 VTAIL.t3 VN.t5 VDD2.t0 w_n1410_n4554# sky130_fd_pr__pfet_01v8 ad=2.95845 pd=18.26 as=2.95845 ps=18.26 w=17.93 l=0.22
X14 B.t2 B.t0 B.t1 w_n1410_n4554# sky130_fd_pr__pfet_01v8 ad=6.9927 pd=36.64 as=0 ps=0 w=17.93 l=0.22
X15 VDD1.t0 VP.t5 VTAIL.t7 w_n1410_n4554# sky130_fd_pr__pfet_01v8 ad=2.95845 pd=18.26 as=6.9927 ps=36.64 w=17.93 l=0.22
R0 VP.n7 VP.t5 2151.47
R1 VP.n5 VP.t2 2151.47
R2 VP.n0 VP.t0 2151.47
R3 VP.n2 VP.t1 2151.47
R4 VP.n6 VP.t4 2107.65
R5 VP.n1 VP.t3 2107.65
R6 VP.n3 VP.n0 161.489
R7 VP.n8 VP.n7 161.3
R8 VP.n3 VP.n2 161.3
R9 VP.n5 VP.n4 161.3
R10 VP.n4 VP.n3 43.8982
R11 VP.n6 VP.n5 36.5157
R12 VP.n7 VP.n6 36.5157
R13 VP.n1 VP.n0 36.5157
R14 VP.n2 VP.n1 36.5157
R15 VP.n8 VP.n4 0.189894
R16 VP VP.n8 0.0516364
R17 VTAIL.n7 VTAIL.t0 54.9545
R18 VTAIL.n11 VTAIL.t1 54.9542
R19 VTAIL.n2 VTAIL.t7 54.9542
R20 VTAIL.n10 VTAIL.t10 54.9542
R21 VTAIL.n9 VTAIL.n8 53.1416
R22 VTAIL.n6 VTAIL.n5 53.1416
R23 VTAIL.n1 VTAIL.n0 53.1414
R24 VTAIL.n4 VTAIL.n3 53.1414
R25 VTAIL.n6 VTAIL.n4 28.7721
R26 VTAIL.n11 VTAIL.n10 28.2979
R27 VTAIL.n0 VTAIL.t5 1.81338
R28 VTAIL.n0 VTAIL.t2 1.81338
R29 VTAIL.n3 VTAIL.t11 1.81338
R30 VTAIL.n3 VTAIL.t6 1.81338
R31 VTAIL.n8 VTAIL.t8 1.81338
R32 VTAIL.n8 VTAIL.t9 1.81338
R33 VTAIL.n5 VTAIL.t4 1.81338
R34 VTAIL.n5 VTAIL.t3 1.81338
R35 VTAIL.n9 VTAIL.n7 0.707397
R36 VTAIL.n2 VTAIL.n1 0.707397
R37 VTAIL.n7 VTAIL.n6 0.474638
R38 VTAIL.n10 VTAIL.n9 0.474638
R39 VTAIL.n4 VTAIL.n2 0.474638
R40 VTAIL VTAIL.n11 0.297914
R41 VTAIL VTAIL.n1 0.177224
R42 VDD1 VDD1.t5 72.0471
R43 VDD1.n1 VDD1.t3 71.9333
R44 VDD1.n1 VDD1.n0 69.8833
R45 VDD1.n3 VDD1.n2 69.8202
R46 VDD1.n3 VDD1.n1 41.5332
R47 VDD1.n2 VDD1.t2 1.81338
R48 VDD1.n2 VDD1.t4 1.81338
R49 VDD1.n0 VDD1.t1 1.81338
R50 VDD1.n0 VDD1.t0 1.81338
R51 VDD1 VDD1.n3 0.0608448
R52 VN.n2 VN.t3 2151.47
R53 VN.n0 VN.t0 2151.47
R54 VN.n6 VN.t1 2151.47
R55 VN.n4 VN.t2 2151.47
R56 VN.n1 VN.t4 2107.65
R57 VN.n5 VN.t5 2107.65
R58 VN.n7 VN.n4 161.489
R59 VN.n3 VN.n0 161.489
R60 VN.n3 VN.n2 161.3
R61 VN.n7 VN.n6 161.3
R62 VN VN.n7 44.2789
R63 VN.n1 VN.n0 36.5157
R64 VN.n2 VN.n1 36.5157
R65 VN.n6 VN.n5 36.5157
R66 VN.n5 VN.n4 36.5157
R67 VN VN.n3 0.0516364
R68 VDD2.n1 VDD2.t5 71.9333
R69 VDD2.n2 VDD2.t4 71.6333
R70 VDD2.n1 VDD2.n0 69.8833
R71 VDD2 VDD2.n3 69.8805
R72 VDD2.n2 VDD2.n1 40.7131
R73 VDD2.n3 VDD2.t0 1.81338
R74 VDD2.n3 VDD2.t3 1.81338
R75 VDD2.n0 VDD2.t1 1.81338
R76 VDD2.n0 VDD2.t2 1.81338
R77 VDD2 VDD2.n2 0.414293
R78 B.n272 B.t9 2195.02
R79 B.n123 B.t3 2195.02
R80 B.n47 B.t0 2195.02
R81 B.n40 B.t6 2195.02
R82 B.n380 B.n93 585
R83 B.n379 B.n378 585
R84 B.n377 B.n94 585
R85 B.n376 B.n375 585
R86 B.n374 B.n95 585
R87 B.n373 B.n372 585
R88 B.n371 B.n96 585
R89 B.n370 B.n369 585
R90 B.n368 B.n97 585
R91 B.n367 B.n366 585
R92 B.n365 B.n98 585
R93 B.n364 B.n363 585
R94 B.n362 B.n99 585
R95 B.n361 B.n360 585
R96 B.n359 B.n100 585
R97 B.n358 B.n357 585
R98 B.n356 B.n101 585
R99 B.n355 B.n354 585
R100 B.n353 B.n102 585
R101 B.n352 B.n351 585
R102 B.n350 B.n103 585
R103 B.n349 B.n348 585
R104 B.n347 B.n104 585
R105 B.n346 B.n345 585
R106 B.n344 B.n105 585
R107 B.n343 B.n342 585
R108 B.n341 B.n106 585
R109 B.n340 B.n339 585
R110 B.n338 B.n107 585
R111 B.n337 B.n336 585
R112 B.n335 B.n108 585
R113 B.n334 B.n333 585
R114 B.n332 B.n109 585
R115 B.n331 B.n330 585
R116 B.n329 B.n110 585
R117 B.n328 B.n327 585
R118 B.n326 B.n111 585
R119 B.n325 B.n324 585
R120 B.n323 B.n112 585
R121 B.n322 B.n321 585
R122 B.n320 B.n113 585
R123 B.n319 B.n318 585
R124 B.n317 B.n114 585
R125 B.n316 B.n315 585
R126 B.n314 B.n115 585
R127 B.n313 B.n312 585
R128 B.n311 B.n116 585
R129 B.n310 B.n309 585
R130 B.n308 B.n117 585
R131 B.n307 B.n306 585
R132 B.n305 B.n118 585
R133 B.n304 B.n303 585
R134 B.n302 B.n119 585
R135 B.n301 B.n300 585
R136 B.n299 B.n120 585
R137 B.n298 B.n297 585
R138 B.n296 B.n121 585
R139 B.n295 B.n294 585
R140 B.n293 B.n122 585
R141 B.n291 B.n290 585
R142 B.n289 B.n125 585
R143 B.n288 B.n287 585
R144 B.n286 B.n126 585
R145 B.n285 B.n284 585
R146 B.n283 B.n127 585
R147 B.n282 B.n281 585
R148 B.n280 B.n128 585
R149 B.n279 B.n278 585
R150 B.n277 B.n129 585
R151 B.n276 B.n275 585
R152 B.n271 B.n130 585
R153 B.n270 B.n269 585
R154 B.n268 B.n131 585
R155 B.n267 B.n266 585
R156 B.n265 B.n132 585
R157 B.n264 B.n263 585
R158 B.n262 B.n133 585
R159 B.n261 B.n260 585
R160 B.n259 B.n134 585
R161 B.n258 B.n257 585
R162 B.n256 B.n135 585
R163 B.n255 B.n254 585
R164 B.n253 B.n136 585
R165 B.n252 B.n251 585
R166 B.n250 B.n137 585
R167 B.n249 B.n248 585
R168 B.n247 B.n138 585
R169 B.n246 B.n245 585
R170 B.n244 B.n139 585
R171 B.n243 B.n242 585
R172 B.n241 B.n140 585
R173 B.n240 B.n239 585
R174 B.n238 B.n141 585
R175 B.n237 B.n236 585
R176 B.n235 B.n142 585
R177 B.n234 B.n233 585
R178 B.n232 B.n143 585
R179 B.n231 B.n230 585
R180 B.n229 B.n144 585
R181 B.n228 B.n227 585
R182 B.n226 B.n145 585
R183 B.n225 B.n224 585
R184 B.n223 B.n146 585
R185 B.n222 B.n221 585
R186 B.n220 B.n147 585
R187 B.n219 B.n218 585
R188 B.n217 B.n148 585
R189 B.n216 B.n215 585
R190 B.n214 B.n149 585
R191 B.n213 B.n212 585
R192 B.n211 B.n150 585
R193 B.n210 B.n209 585
R194 B.n208 B.n151 585
R195 B.n207 B.n206 585
R196 B.n205 B.n152 585
R197 B.n204 B.n203 585
R198 B.n202 B.n153 585
R199 B.n201 B.n200 585
R200 B.n199 B.n154 585
R201 B.n198 B.n197 585
R202 B.n196 B.n155 585
R203 B.n195 B.n194 585
R204 B.n193 B.n156 585
R205 B.n192 B.n191 585
R206 B.n190 B.n157 585
R207 B.n189 B.n188 585
R208 B.n187 B.n158 585
R209 B.n186 B.n185 585
R210 B.n382 B.n381 585
R211 B.n383 B.n92 585
R212 B.n385 B.n384 585
R213 B.n386 B.n91 585
R214 B.n388 B.n387 585
R215 B.n389 B.n90 585
R216 B.n391 B.n390 585
R217 B.n392 B.n89 585
R218 B.n394 B.n393 585
R219 B.n395 B.n88 585
R220 B.n397 B.n396 585
R221 B.n398 B.n87 585
R222 B.n400 B.n399 585
R223 B.n401 B.n86 585
R224 B.n403 B.n402 585
R225 B.n404 B.n85 585
R226 B.n406 B.n405 585
R227 B.n407 B.n84 585
R228 B.n409 B.n408 585
R229 B.n410 B.n83 585
R230 B.n412 B.n411 585
R231 B.n413 B.n82 585
R232 B.n415 B.n414 585
R233 B.n416 B.n81 585
R234 B.n418 B.n417 585
R235 B.n419 B.n80 585
R236 B.n421 B.n420 585
R237 B.n422 B.n79 585
R238 B.n424 B.n423 585
R239 B.n425 B.n78 585
R240 B.n618 B.n9 585
R241 B.n617 B.n616 585
R242 B.n615 B.n10 585
R243 B.n614 B.n613 585
R244 B.n612 B.n11 585
R245 B.n611 B.n610 585
R246 B.n609 B.n12 585
R247 B.n608 B.n607 585
R248 B.n606 B.n13 585
R249 B.n605 B.n604 585
R250 B.n603 B.n14 585
R251 B.n602 B.n601 585
R252 B.n600 B.n15 585
R253 B.n599 B.n598 585
R254 B.n597 B.n16 585
R255 B.n596 B.n595 585
R256 B.n594 B.n17 585
R257 B.n593 B.n592 585
R258 B.n591 B.n18 585
R259 B.n590 B.n589 585
R260 B.n588 B.n19 585
R261 B.n587 B.n586 585
R262 B.n585 B.n20 585
R263 B.n584 B.n583 585
R264 B.n582 B.n21 585
R265 B.n581 B.n580 585
R266 B.n579 B.n22 585
R267 B.n578 B.n577 585
R268 B.n576 B.n23 585
R269 B.n575 B.n574 585
R270 B.n573 B.n24 585
R271 B.n572 B.n571 585
R272 B.n570 B.n25 585
R273 B.n569 B.n568 585
R274 B.n567 B.n26 585
R275 B.n566 B.n565 585
R276 B.n564 B.n27 585
R277 B.n563 B.n562 585
R278 B.n561 B.n28 585
R279 B.n560 B.n559 585
R280 B.n558 B.n29 585
R281 B.n557 B.n556 585
R282 B.n555 B.n30 585
R283 B.n554 B.n553 585
R284 B.n552 B.n31 585
R285 B.n551 B.n550 585
R286 B.n549 B.n32 585
R287 B.n548 B.n547 585
R288 B.n546 B.n33 585
R289 B.n545 B.n544 585
R290 B.n543 B.n34 585
R291 B.n542 B.n541 585
R292 B.n540 B.n35 585
R293 B.n539 B.n538 585
R294 B.n537 B.n36 585
R295 B.n536 B.n535 585
R296 B.n534 B.n37 585
R297 B.n533 B.n532 585
R298 B.n531 B.n38 585
R299 B.n530 B.n529 585
R300 B.n528 B.n39 585
R301 B.n527 B.n526 585
R302 B.n525 B.n43 585
R303 B.n524 B.n523 585
R304 B.n522 B.n44 585
R305 B.n521 B.n520 585
R306 B.n519 B.n45 585
R307 B.n518 B.n517 585
R308 B.n516 B.n46 585
R309 B.n514 B.n513 585
R310 B.n512 B.n49 585
R311 B.n511 B.n510 585
R312 B.n509 B.n50 585
R313 B.n508 B.n507 585
R314 B.n506 B.n51 585
R315 B.n505 B.n504 585
R316 B.n503 B.n52 585
R317 B.n502 B.n501 585
R318 B.n500 B.n53 585
R319 B.n499 B.n498 585
R320 B.n497 B.n54 585
R321 B.n496 B.n495 585
R322 B.n494 B.n55 585
R323 B.n493 B.n492 585
R324 B.n491 B.n56 585
R325 B.n490 B.n489 585
R326 B.n488 B.n57 585
R327 B.n487 B.n486 585
R328 B.n485 B.n58 585
R329 B.n484 B.n483 585
R330 B.n482 B.n59 585
R331 B.n481 B.n480 585
R332 B.n479 B.n60 585
R333 B.n478 B.n477 585
R334 B.n476 B.n61 585
R335 B.n475 B.n474 585
R336 B.n473 B.n62 585
R337 B.n472 B.n471 585
R338 B.n470 B.n63 585
R339 B.n469 B.n468 585
R340 B.n467 B.n64 585
R341 B.n466 B.n465 585
R342 B.n464 B.n65 585
R343 B.n463 B.n462 585
R344 B.n461 B.n66 585
R345 B.n460 B.n459 585
R346 B.n458 B.n67 585
R347 B.n457 B.n456 585
R348 B.n455 B.n68 585
R349 B.n454 B.n453 585
R350 B.n452 B.n69 585
R351 B.n451 B.n450 585
R352 B.n449 B.n70 585
R353 B.n448 B.n447 585
R354 B.n446 B.n71 585
R355 B.n445 B.n444 585
R356 B.n443 B.n72 585
R357 B.n442 B.n441 585
R358 B.n440 B.n73 585
R359 B.n439 B.n438 585
R360 B.n437 B.n74 585
R361 B.n436 B.n435 585
R362 B.n434 B.n75 585
R363 B.n433 B.n432 585
R364 B.n431 B.n76 585
R365 B.n430 B.n429 585
R366 B.n428 B.n77 585
R367 B.n427 B.n426 585
R368 B.n620 B.n619 585
R369 B.n621 B.n8 585
R370 B.n623 B.n622 585
R371 B.n624 B.n7 585
R372 B.n626 B.n625 585
R373 B.n627 B.n6 585
R374 B.n629 B.n628 585
R375 B.n630 B.n5 585
R376 B.n632 B.n631 585
R377 B.n633 B.n4 585
R378 B.n635 B.n634 585
R379 B.n636 B.n3 585
R380 B.n638 B.n637 585
R381 B.n639 B.n0 585
R382 B.n2 B.n1 585
R383 B.n166 B.n165 585
R384 B.n168 B.n167 585
R385 B.n169 B.n164 585
R386 B.n171 B.n170 585
R387 B.n172 B.n163 585
R388 B.n174 B.n173 585
R389 B.n175 B.n162 585
R390 B.n177 B.n176 585
R391 B.n178 B.n161 585
R392 B.n180 B.n179 585
R393 B.n181 B.n160 585
R394 B.n183 B.n182 585
R395 B.n184 B.n159 585
R396 B.n185 B.n184 487.695
R397 B.n381 B.n380 487.695
R398 B.n427 B.n78 487.695
R399 B.n620 B.n9 487.695
R400 B.n641 B.n640 256.663
R401 B.n640 B.n639 235.042
R402 B.n640 B.n2 235.042
R403 B.n185 B.n158 163.367
R404 B.n189 B.n158 163.367
R405 B.n190 B.n189 163.367
R406 B.n191 B.n190 163.367
R407 B.n191 B.n156 163.367
R408 B.n195 B.n156 163.367
R409 B.n196 B.n195 163.367
R410 B.n197 B.n196 163.367
R411 B.n197 B.n154 163.367
R412 B.n201 B.n154 163.367
R413 B.n202 B.n201 163.367
R414 B.n203 B.n202 163.367
R415 B.n203 B.n152 163.367
R416 B.n207 B.n152 163.367
R417 B.n208 B.n207 163.367
R418 B.n209 B.n208 163.367
R419 B.n209 B.n150 163.367
R420 B.n213 B.n150 163.367
R421 B.n214 B.n213 163.367
R422 B.n215 B.n214 163.367
R423 B.n215 B.n148 163.367
R424 B.n219 B.n148 163.367
R425 B.n220 B.n219 163.367
R426 B.n221 B.n220 163.367
R427 B.n221 B.n146 163.367
R428 B.n225 B.n146 163.367
R429 B.n226 B.n225 163.367
R430 B.n227 B.n226 163.367
R431 B.n227 B.n144 163.367
R432 B.n231 B.n144 163.367
R433 B.n232 B.n231 163.367
R434 B.n233 B.n232 163.367
R435 B.n233 B.n142 163.367
R436 B.n237 B.n142 163.367
R437 B.n238 B.n237 163.367
R438 B.n239 B.n238 163.367
R439 B.n239 B.n140 163.367
R440 B.n243 B.n140 163.367
R441 B.n244 B.n243 163.367
R442 B.n245 B.n244 163.367
R443 B.n245 B.n138 163.367
R444 B.n249 B.n138 163.367
R445 B.n250 B.n249 163.367
R446 B.n251 B.n250 163.367
R447 B.n251 B.n136 163.367
R448 B.n255 B.n136 163.367
R449 B.n256 B.n255 163.367
R450 B.n257 B.n256 163.367
R451 B.n257 B.n134 163.367
R452 B.n261 B.n134 163.367
R453 B.n262 B.n261 163.367
R454 B.n263 B.n262 163.367
R455 B.n263 B.n132 163.367
R456 B.n267 B.n132 163.367
R457 B.n268 B.n267 163.367
R458 B.n269 B.n268 163.367
R459 B.n269 B.n130 163.367
R460 B.n276 B.n130 163.367
R461 B.n277 B.n276 163.367
R462 B.n278 B.n277 163.367
R463 B.n278 B.n128 163.367
R464 B.n282 B.n128 163.367
R465 B.n283 B.n282 163.367
R466 B.n284 B.n283 163.367
R467 B.n284 B.n126 163.367
R468 B.n288 B.n126 163.367
R469 B.n289 B.n288 163.367
R470 B.n290 B.n289 163.367
R471 B.n290 B.n122 163.367
R472 B.n295 B.n122 163.367
R473 B.n296 B.n295 163.367
R474 B.n297 B.n296 163.367
R475 B.n297 B.n120 163.367
R476 B.n301 B.n120 163.367
R477 B.n302 B.n301 163.367
R478 B.n303 B.n302 163.367
R479 B.n303 B.n118 163.367
R480 B.n307 B.n118 163.367
R481 B.n308 B.n307 163.367
R482 B.n309 B.n308 163.367
R483 B.n309 B.n116 163.367
R484 B.n313 B.n116 163.367
R485 B.n314 B.n313 163.367
R486 B.n315 B.n314 163.367
R487 B.n315 B.n114 163.367
R488 B.n319 B.n114 163.367
R489 B.n320 B.n319 163.367
R490 B.n321 B.n320 163.367
R491 B.n321 B.n112 163.367
R492 B.n325 B.n112 163.367
R493 B.n326 B.n325 163.367
R494 B.n327 B.n326 163.367
R495 B.n327 B.n110 163.367
R496 B.n331 B.n110 163.367
R497 B.n332 B.n331 163.367
R498 B.n333 B.n332 163.367
R499 B.n333 B.n108 163.367
R500 B.n337 B.n108 163.367
R501 B.n338 B.n337 163.367
R502 B.n339 B.n338 163.367
R503 B.n339 B.n106 163.367
R504 B.n343 B.n106 163.367
R505 B.n344 B.n343 163.367
R506 B.n345 B.n344 163.367
R507 B.n345 B.n104 163.367
R508 B.n349 B.n104 163.367
R509 B.n350 B.n349 163.367
R510 B.n351 B.n350 163.367
R511 B.n351 B.n102 163.367
R512 B.n355 B.n102 163.367
R513 B.n356 B.n355 163.367
R514 B.n357 B.n356 163.367
R515 B.n357 B.n100 163.367
R516 B.n361 B.n100 163.367
R517 B.n362 B.n361 163.367
R518 B.n363 B.n362 163.367
R519 B.n363 B.n98 163.367
R520 B.n367 B.n98 163.367
R521 B.n368 B.n367 163.367
R522 B.n369 B.n368 163.367
R523 B.n369 B.n96 163.367
R524 B.n373 B.n96 163.367
R525 B.n374 B.n373 163.367
R526 B.n375 B.n374 163.367
R527 B.n375 B.n94 163.367
R528 B.n379 B.n94 163.367
R529 B.n380 B.n379 163.367
R530 B.n423 B.n78 163.367
R531 B.n423 B.n422 163.367
R532 B.n422 B.n421 163.367
R533 B.n421 B.n80 163.367
R534 B.n417 B.n80 163.367
R535 B.n417 B.n416 163.367
R536 B.n416 B.n415 163.367
R537 B.n415 B.n82 163.367
R538 B.n411 B.n82 163.367
R539 B.n411 B.n410 163.367
R540 B.n410 B.n409 163.367
R541 B.n409 B.n84 163.367
R542 B.n405 B.n84 163.367
R543 B.n405 B.n404 163.367
R544 B.n404 B.n403 163.367
R545 B.n403 B.n86 163.367
R546 B.n399 B.n86 163.367
R547 B.n399 B.n398 163.367
R548 B.n398 B.n397 163.367
R549 B.n397 B.n88 163.367
R550 B.n393 B.n88 163.367
R551 B.n393 B.n392 163.367
R552 B.n392 B.n391 163.367
R553 B.n391 B.n90 163.367
R554 B.n387 B.n90 163.367
R555 B.n387 B.n386 163.367
R556 B.n386 B.n385 163.367
R557 B.n385 B.n92 163.367
R558 B.n381 B.n92 163.367
R559 B.n616 B.n9 163.367
R560 B.n616 B.n615 163.367
R561 B.n615 B.n614 163.367
R562 B.n614 B.n11 163.367
R563 B.n610 B.n11 163.367
R564 B.n610 B.n609 163.367
R565 B.n609 B.n608 163.367
R566 B.n608 B.n13 163.367
R567 B.n604 B.n13 163.367
R568 B.n604 B.n603 163.367
R569 B.n603 B.n602 163.367
R570 B.n602 B.n15 163.367
R571 B.n598 B.n15 163.367
R572 B.n598 B.n597 163.367
R573 B.n597 B.n596 163.367
R574 B.n596 B.n17 163.367
R575 B.n592 B.n17 163.367
R576 B.n592 B.n591 163.367
R577 B.n591 B.n590 163.367
R578 B.n590 B.n19 163.367
R579 B.n586 B.n19 163.367
R580 B.n586 B.n585 163.367
R581 B.n585 B.n584 163.367
R582 B.n584 B.n21 163.367
R583 B.n580 B.n21 163.367
R584 B.n580 B.n579 163.367
R585 B.n579 B.n578 163.367
R586 B.n578 B.n23 163.367
R587 B.n574 B.n23 163.367
R588 B.n574 B.n573 163.367
R589 B.n573 B.n572 163.367
R590 B.n572 B.n25 163.367
R591 B.n568 B.n25 163.367
R592 B.n568 B.n567 163.367
R593 B.n567 B.n566 163.367
R594 B.n566 B.n27 163.367
R595 B.n562 B.n27 163.367
R596 B.n562 B.n561 163.367
R597 B.n561 B.n560 163.367
R598 B.n560 B.n29 163.367
R599 B.n556 B.n29 163.367
R600 B.n556 B.n555 163.367
R601 B.n555 B.n554 163.367
R602 B.n554 B.n31 163.367
R603 B.n550 B.n31 163.367
R604 B.n550 B.n549 163.367
R605 B.n549 B.n548 163.367
R606 B.n548 B.n33 163.367
R607 B.n544 B.n33 163.367
R608 B.n544 B.n543 163.367
R609 B.n543 B.n542 163.367
R610 B.n542 B.n35 163.367
R611 B.n538 B.n35 163.367
R612 B.n538 B.n537 163.367
R613 B.n537 B.n536 163.367
R614 B.n536 B.n37 163.367
R615 B.n532 B.n37 163.367
R616 B.n532 B.n531 163.367
R617 B.n531 B.n530 163.367
R618 B.n530 B.n39 163.367
R619 B.n526 B.n39 163.367
R620 B.n526 B.n525 163.367
R621 B.n525 B.n524 163.367
R622 B.n524 B.n44 163.367
R623 B.n520 B.n44 163.367
R624 B.n520 B.n519 163.367
R625 B.n519 B.n518 163.367
R626 B.n518 B.n46 163.367
R627 B.n513 B.n46 163.367
R628 B.n513 B.n512 163.367
R629 B.n512 B.n511 163.367
R630 B.n511 B.n50 163.367
R631 B.n507 B.n50 163.367
R632 B.n507 B.n506 163.367
R633 B.n506 B.n505 163.367
R634 B.n505 B.n52 163.367
R635 B.n501 B.n52 163.367
R636 B.n501 B.n500 163.367
R637 B.n500 B.n499 163.367
R638 B.n499 B.n54 163.367
R639 B.n495 B.n54 163.367
R640 B.n495 B.n494 163.367
R641 B.n494 B.n493 163.367
R642 B.n493 B.n56 163.367
R643 B.n489 B.n56 163.367
R644 B.n489 B.n488 163.367
R645 B.n488 B.n487 163.367
R646 B.n487 B.n58 163.367
R647 B.n483 B.n58 163.367
R648 B.n483 B.n482 163.367
R649 B.n482 B.n481 163.367
R650 B.n481 B.n60 163.367
R651 B.n477 B.n60 163.367
R652 B.n477 B.n476 163.367
R653 B.n476 B.n475 163.367
R654 B.n475 B.n62 163.367
R655 B.n471 B.n62 163.367
R656 B.n471 B.n470 163.367
R657 B.n470 B.n469 163.367
R658 B.n469 B.n64 163.367
R659 B.n465 B.n64 163.367
R660 B.n465 B.n464 163.367
R661 B.n464 B.n463 163.367
R662 B.n463 B.n66 163.367
R663 B.n459 B.n66 163.367
R664 B.n459 B.n458 163.367
R665 B.n458 B.n457 163.367
R666 B.n457 B.n68 163.367
R667 B.n453 B.n68 163.367
R668 B.n453 B.n452 163.367
R669 B.n452 B.n451 163.367
R670 B.n451 B.n70 163.367
R671 B.n447 B.n70 163.367
R672 B.n447 B.n446 163.367
R673 B.n446 B.n445 163.367
R674 B.n445 B.n72 163.367
R675 B.n441 B.n72 163.367
R676 B.n441 B.n440 163.367
R677 B.n440 B.n439 163.367
R678 B.n439 B.n74 163.367
R679 B.n435 B.n74 163.367
R680 B.n435 B.n434 163.367
R681 B.n434 B.n433 163.367
R682 B.n433 B.n76 163.367
R683 B.n429 B.n76 163.367
R684 B.n429 B.n428 163.367
R685 B.n428 B.n427 163.367
R686 B.n621 B.n620 163.367
R687 B.n622 B.n621 163.367
R688 B.n622 B.n7 163.367
R689 B.n626 B.n7 163.367
R690 B.n627 B.n626 163.367
R691 B.n628 B.n627 163.367
R692 B.n628 B.n5 163.367
R693 B.n632 B.n5 163.367
R694 B.n633 B.n632 163.367
R695 B.n634 B.n633 163.367
R696 B.n634 B.n3 163.367
R697 B.n638 B.n3 163.367
R698 B.n639 B.n638 163.367
R699 B.n166 B.n2 163.367
R700 B.n167 B.n166 163.367
R701 B.n167 B.n164 163.367
R702 B.n171 B.n164 163.367
R703 B.n172 B.n171 163.367
R704 B.n173 B.n172 163.367
R705 B.n173 B.n162 163.367
R706 B.n177 B.n162 163.367
R707 B.n178 B.n177 163.367
R708 B.n179 B.n178 163.367
R709 B.n179 B.n160 163.367
R710 B.n183 B.n160 163.367
R711 B.n184 B.n183 163.367
R712 B.n123 B.t4 121.725
R713 B.n47 B.t2 121.725
R714 B.n272 B.t10 121.703
R715 B.n40 B.t8 121.703
R716 B.n124 B.t5 111.059
R717 B.n48 B.t1 111.059
R718 B.n273 B.t11 111.037
R719 B.n41 B.t7 111.037
R720 B.n274 B.n273 59.5399
R721 B.n292 B.n124 59.5399
R722 B.n515 B.n48 59.5399
R723 B.n42 B.n41 59.5399
R724 B.n619 B.n618 31.6883
R725 B.n426 B.n425 31.6883
R726 B.n382 B.n93 31.6883
R727 B.n186 B.n159 31.6883
R728 B B.n641 18.0485
R729 B.n273 B.n272 10.6672
R730 B.n124 B.n123 10.6672
R731 B.n48 B.n47 10.6672
R732 B.n41 B.n40 10.6672
R733 B.n619 B.n8 10.6151
R734 B.n623 B.n8 10.6151
R735 B.n624 B.n623 10.6151
R736 B.n625 B.n624 10.6151
R737 B.n625 B.n6 10.6151
R738 B.n629 B.n6 10.6151
R739 B.n630 B.n629 10.6151
R740 B.n631 B.n630 10.6151
R741 B.n631 B.n4 10.6151
R742 B.n635 B.n4 10.6151
R743 B.n636 B.n635 10.6151
R744 B.n637 B.n636 10.6151
R745 B.n637 B.n0 10.6151
R746 B.n618 B.n617 10.6151
R747 B.n617 B.n10 10.6151
R748 B.n613 B.n10 10.6151
R749 B.n613 B.n612 10.6151
R750 B.n612 B.n611 10.6151
R751 B.n611 B.n12 10.6151
R752 B.n607 B.n12 10.6151
R753 B.n607 B.n606 10.6151
R754 B.n606 B.n605 10.6151
R755 B.n605 B.n14 10.6151
R756 B.n601 B.n14 10.6151
R757 B.n601 B.n600 10.6151
R758 B.n600 B.n599 10.6151
R759 B.n599 B.n16 10.6151
R760 B.n595 B.n16 10.6151
R761 B.n595 B.n594 10.6151
R762 B.n594 B.n593 10.6151
R763 B.n593 B.n18 10.6151
R764 B.n589 B.n18 10.6151
R765 B.n589 B.n588 10.6151
R766 B.n588 B.n587 10.6151
R767 B.n587 B.n20 10.6151
R768 B.n583 B.n20 10.6151
R769 B.n583 B.n582 10.6151
R770 B.n582 B.n581 10.6151
R771 B.n581 B.n22 10.6151
R772 B.n577 B.n22 10.6151
R773 B.n577 B.n576 10.6151
R774 B.n576 B.n575 10.6151
R775 B.n575 B.n24 10.6151
R776 B.n571 B.n24 10.6151
R777 B.n571 B.n570 10.6151
R778 B.n570 B.n569 10.6151
R779 B.n569 B.n26 10.6151
R780 B.n565 B.n26 10.6151
R781 B.n565 B.n564 10.6151
R782 B.n564 B.n563 10.6151
R783 B.n563 B.n28 10.6151
R784 B.n559 B.n28 10.6151
R785 B.n559 B.n558 10.6151
R786 B.n558 B.n557 10.6151
R787 B.n557 B.n30 10.6151
R788 B.n553 B.n30 10.6151
R789 B.n553 B.n552 10.6151
R790 B.n552 B.n551 10.6151
R791 B.n551 B.n32 10.6151
R792 B.n547 B.n32 10.6151
R793 B.n547 B.n546 10.6151
R794 B.n546 B.n545 10.6151
R795 B.n545 B.n34 10.6151
R796 B.n541 B.n34 10.6151
R797 B.n541 B.n540 10.6151
R798 B.n540 B.n539 10.6151
R799 B.n539 B.n36 10.6151
R800 B.n535 B.n36 10.6151
R801 B.n535 B.n534 10.6151
R802 B.n534 B.n533 10.6151
R803 B.n533 B.n38 10.6151
R804 B.n529 B.n528 10.6151
R805 B.n528 B.n527 10.6151
R806 B.n527 B.n43 10.6151
R807 B.n523 B.n43 10.6151
R808 B.n523 B.n522 10.6151
R809 B.n522 B.n521 10.6151
R810 B.n521 B.n45 10.6151
R811 B.n517 B.n45 10.6151
R812 B.n517 B.n516 10.6151
R813 B.n514 B.n49 10.6151
R814 B.n510 B.n49 10.6151
R815 B.n510 B.n509 10.6151
R816 B.n509 B.n508 10.6151
R817 B.n508 B.n51 10.6151
R818 B.n504 B.n51 10.6151
R819 B.n504 B.n503 10.6151
R820 B.n503 B.n502 10.6151
R821 B.n502 B.n53 10.6151
R822 B.n498 B.n53 10.6151
R823 B.n498 B.n497 10.6151
R824 B.n497 B.n496 10.6151
R825 B.n496 B.n55 10.6151
R826 B.n492 B.n55 10.6151
R827 B.n492 B.n491 10.6151
R828 B.n491 B.n490 10.6151
R829 B.n490 B.n57 10.6151
R830 B.n486 B.n57 10.6151
R831 B.n486 B.n485 10.6151
R832 B.n485 B.n484 10.6151
R833 B.n484 B.n59 10.6151
R834 B.n480 B.n59 10.6151
R835 B.n480 B.n479 10.6151
R836 B.n479 B.n478 10.6151
R837 B.n478 B.n61 10.6151
R838 B.n474 B.n61 10.6151
R839 B.n474 B.n473 10.6151
R840 B.n473 B.n472 10.6151
R841 B.n472 B.n63 10.6151
R842 B.n468 B.n63 10.6151
R843 B.n468 B.n467 10.6151
R844 B.n467 B.n466 10.6151
R845 B.n466 B.n65 10.6151
R846 B.n462 B.n65 10.6151
R847 B.n462 B.n461 10.6151
R848 B.n461 B.n460 10.6151
R849 B.n460 B.n67 10.6151
R850 B.n456 B.n67 10.6151
R851 B.n456 B.n455 10.6151
R852 B.n455 B.n454 10.6151
R853 B.n454 B.n69 10.6151
R854 B.n450 B.n69 10.6151
R855 B.n450 B.n449 10.6151
R856 B.n449 B.n448 10.6151
R857 B.n448 B.n71 10.6151
R858 B.n444 B.n71 10.6151
R859 B.n444 B.n443 10.6151
R860 B.n443 B.n442 10.6151
R861 B.n442 B.n73 10.6151
R862 B.n438 B.n73 10.6151
R863 B.n438 B.n437 10.6151
R864 B.n437 B.n436 10.6151
R865 B.n436 B.n75 10.6151
R866 B.n432 B.n75 10.6151
R867 B.n432 B.n431 10.6151
R868 B.n431 B.n430 10.6151
R869 B.n430 B.n77 10.6151
R870 B.n426 B.n77 10.6151
R871 B.n425 B.n424 10.6151
R872 B.n424 B.n79 10.6151
R873 B.n420 B.n79 10.6151
R874 B.n420 B.n419 10.6151
R875 B.n419 B.n418 10.6151
R876 B.n418 B.n81 10.6151
R877 B.n414 B.n81 10.6151
R878 B.n414 B.n413 10.6151
R879 B.n413 B.n412 10.6151
R880 B.n412 B.n83 10.6151
R881 B.n408 B.n83 10.6151
R882 B.n408 B.n407 10.6151
R883 B.n407 B.n406 10.6151
R884 B.n406 B.n85 10.6151
R885 B.n402 B.n85 10.6151
R886 B.n402 B.n401 10.6151
R887 B.n401 B.n400 10.6151
R888 B.n400 B.n87 10.6151
R889 B.n396 B.n87 10.6151
R890 B.n396 B.n395 10.6151
R891 B.n395 B.n394 10.6151
R892 B.n394 B.n89 10.6151
R893 B.n390 B.n89 10.6151
R894 B.n390 B.n389 10.6151
R895 B.n389 B.n388 10.6151
R896 B.n388 B.n91 10.6151
R897 B.n384 B.n91 10.6151
R898 B.n384 B.n383 10.6151
R899 B.n383 B.n382 10.6151
R900 B.n165 B.n1 10.6151
R901 B.n168 B.n165 10.6151
R902 B.n169 B.n168 10.6151
R903 B.n170 B.n169 10.6151
R904 B.n170 B.n163 10.6151
R905 B.n174 B.n163 10.6151
R906 B.n175 B.n174 10.6151
R907 B.n176 B.n175 10.6151
R908 B.n176 B.n161 10.6151
R909 B.n180 B.n161 10.6151
R910 B.n181 B.n180 10.6151
R911 B.n182 B.n181 10.6151
R912 B.n182 B.n159 10.6151
R913 B.n187 B.n186 10.6151
R914 B.n188 B.n187 10.6151
R915 B.n188 B.n157 10.6151
R916 B.n192 B.n157 10.6151
R917 B.n193 B.n192 10.6151
R918 B.n194 B.n193 10.6151
R919 B.n194 B.n155 10.6151
R920 B.n198 B.n155 10.6151
R921 B.n199 B.n198 10.6151
R922 B.n200 B.n199 10.6151
R923 B.n200 B.n153 10.6151
R924 B.n204 B.n153 10.6151
R925 B.n205 B.n204 10.6151
R926 B.n206 B.n205 10.6151
R927 B.n206 B.n151 10.6151
R928 B.n210 B.n151 10.6151
R929 B.n211 B.n210 10.6151
R930 B.n212 B.n211 10.6151
R931 B.n212 B.n149 10.6151
R932 B.n216 B.n149 10.6151
R933 B.n217 B.n216 10.6151
R934 B.n218 B.n217 10.6151
R935 B.n218 B.n147 10.6151
R936 B.n222 B.n147 10.6151
R937 B.n223 B.n222 10.6151
R938 B.n224 B.n223 10.6151
R939 B.n224 B.n145 10.6151
R940 B.n228 B.n145 10.6151
R941 B.n229 B.n228 10.6151
R942 B.n230 B.n229 10.6151
R943 B.n230 B.n143 10.6151
R944 B.n234 B.n143 10.6151
R945 B.n235 B.n234 10.6151
R946 B.n236 B.n235 10.6151
R947 B.n236 B.n141 10.6151
R948 B.n240 B.n141 10.6151
R949 B.n241 B.n240 10.6151
R950 B.n242 B.n241 10.6151
R951 B.n242 B.n139 10.6151
R952 B.n246 B.n139 10.6151
R953 B.n247 B.n246 10.6151
R954 B.n248 B.n247 10.6151
R955 B.n248 B.n137 10.6151
R956 B.n252 B.n137 10.6151
R957 B.n253 B.n252 10.6151
R958 B.n254 B.n253 10.6151
R959 B.n254 B.n135 10.6151
R960 B.n258 B.n135 10.6151
R961 B.n259 B.n258 10.6151
R962 B.n260 B.n259 10.6151
R963 B.n260 B.n133 10.6151
R964 B.n264 B.n133 10.6151
R965 B.n265 B.n264 10.6151
R966 B.n266 B.n265 10.6151
R967 B.n266 B.n131 10.6151
R968 B.n270 B.n131 10.6151
R969 B.n271 B.n270 10.6151
R970 B.n275 B.n271 10.6151
R971 B.n279 B.n129 10.6151
R972 B.n280 B.n279 10.6151
R973 B.n281 B.n280 10.6151
R974 B.n281 B.n127 10.6151
R975 B.n285 B.n127 10.6151
R976 B.n286 B.n285 10.6151
R977 B.n287 B.n286 10.6151
R978 B.n287 B.n125 10.6151
R979 B.n291 B.n125 10.6151
R980 B.n294 B.n293 10.6151
R981 B.n294 B.n121 10.6151
R982 B.n298 B.n121 10.6151
R983 B.n299 B.n298 10.6151
R984 B.n300 B.n299 10.6151
R985 B.n300 B.n119 10.6151
R986 B.n304 B.n119 10.6151
R987 B.n305 B.n304 10.6151
R988 B.n306 B.n305 10.6151
R989 B.n306 B.n117 10.6151
R990 B.n310 B.n117 10.6151
R991 B.n311 B.n310 10.6151
R992 B.n312 B.n311 10.6151
R993 B.n312 B.n115 10.6151
R994 B.n316 B.n115 10.6151
R995 B.n317 B.n316 10.6151
R996 B.n318 B.n317 10.6151
R997 B.n318 B.n113 10.6151
R998 B.n322 B.n113 10.6151
R999 B.n323 B.n322 10.6151
R1000 B.n324 B.n323 10.6151
R1001 B.n324 B.n111 10.6151
R1002 B.n328 B.n111 10.6151
R1003 B.n329 B.n328 10.6151
R1004 B.n330 B.n329 10.6151
R1005 B.n330 B.n109 10.6151
R1006 B.n334 B.n109 10.6151
R1007 B.n335 B.n334 10.6151
R1008 B.n336 B.n335 10.6151
R1009 B.n336 B.n107 10.6151
R1010 B.n340 B.n107 10.6151
R1011 B.n341 B.n340 10.6151
R1012 B.n342 B.n341 10.6151
R1013 B.n342 B.n105 10.6151
R1014 B.n346 B.n105 10.6151
R1015 B.n347 B.n346 10.6151
R1016 B.n348 B.n347 10.6151
R1017 B.n348 B.n103 10.6151
R1018 B.n352 B.n103 10.6151
R1019 B.n353 B.n352 10.6151
R1020 B.n354 B.n353 10.6151
R1021 B.n354 B.n101 10.6151
R1022 B.n358 B.n101 10.6151
R1023 B.n359 B.n358 10.6151
R1024 B.n360 B.n359 10.6151
R1025 B.n360 B.n99 10.6151
R1026 B.n364 B.n99 10.6151
R1027 B.n365 B.n364 10.6151
R1028 B.n366 B.n365 10.6151
R1029 B.n366 B.n97 10.6151
R1030 B.n370 B.n97 10.6151
R1031 B.n371 B.n370 10.6151
R1032 B.n372 B.n371 10.6151
R1033 B.n372 B.n95 10.6151
R1034 B.n376 B.n95 10.6151
R1035 B.n377 B.n376 10.6151
R1036 B.n378 B.n377 10.6151
R1037 B.n378 B.n93 10.6151
R1038 B.n42 B.n38 9.36635
R1039 B.n515 B.n514 9.36635
R1040 B.n275 B.n274 9.36635
R1041 B.n293 B.n292 9.36635
R1042 B.n641 B.n0 8.11757
R1043 B.n641 B.n1 8.11757
R1044 B.n529 B.n42 1.24928
R1045 B.n516 B.n515 1.24928
R1046 B.n274 B.n129 1.24928
R1047 B.n292 B.n291 1.24928
C0 VP VN 5.71247f
C1 VDD2 w_n1410_n4554# 2.12723f
C2 VN VDD1 0.147281f
C3 VP VDD2 0.258119f
C4 B w_n1410_n4554# 8.10323f
C5 B VP 1.01014f
C6 VTAIL VN 2.47479f
C7 VDD2 VDD1 0.544608f
C8 B VDD1 1.8184f
C9 VTAIL VDD2 22.705801f
C10 VP w_n1410_n4554# 2.38569f
C11 B VTAIL 3.33236f
C12 VDD1 w_n1410_n4554# 2.1173f
C13 VP VDD1 3.35333f
C14 VTAIL w_n1410_n4554# 4.03061f
C15 VTAIL VP 2.48993f
C16 VDD2 VN 3.2503f
C17 B VN 0.728835f
C18 VTAIL VDD1 22.6818f
C19 B VDD2 1.83695f
C20 VN w_n1410_n4554# 2.21002f
C21 VDD2 VSUBS 1.658854f
C22 VDD1 VSUBS 1.933471f
C23 VTAIL VSUBS 0.679067f
C24 VN VSUBS 5.15984f
C25 VP VSUBS 1.329838f
C26 B VSUBS 2.773073f
C27 w_n1410_n4554# VSUBS 78.5257f
C28 B.n0 VSUBS 0.006541f
C29 B.n1 VSUBS 0.006541f
C30 B.n2 VSUBS 0.009674f
C31 B.n3 VSUBS 0.007414f
C32 B.n4 VSUBS 0.007414f
C33 B.n5 VSUBS 0.007414f
C34 B.n6 VSUBS 0.007414f
C35 B.n7 VSUBS 0.007414f
C36 B.n8 VSUBS 0.007414f
C37 B.n9 VSUBS 0.017613f
C38 B.n10 VSUBS 0.007414f
C39 B.n11 VSUBS 0.007414f
C40 B.n12 VSUBS 0.007414f
C41 B.n13 VSUBS 0.007414f
C42 B.n14 VSUBS 0.007414f
C43 B.n15 VSUBS 0.007414f
C44 B.n16 VSUBS 0.007414f
C45 B.n17 VSUBS 0.007414f
C46 B.n18 VSUBS 0.007414f
C47 B.n19 VSUBS 0.007414f
C48 B.n20 VSUBS 0.007414f
C49 B.n21 VSUBS 0.007414f
C50 B.n22 VSUBS 0.007414f
C51 B.n23 VSUBS 0.007414f
C52 B.n24 VSUBS 0.007414f
C53 B.n25 VSUBS 0.007414f
C54 B.n26 VSUBS 0.007414f
C55 B.n27 VSUBS 0.007414f
C56 B.n28 VSUBS 0.007414f
C57 B.n29 VSUBS 0.007414f
C58 B.n30 VSUBS 0.007414f
C59 B.n31 VSUBS 0.007414f
C60 B.n32 VSUBS 0.007414f
C61 B.n33 VSUBS 0.007414f
C62 B.n34 VSUBS 0.007414f
C63 B.n35 VSUBS 0.007414f
C64 B.n36 VSUBS 0.007414f
C65 B.n37 VSUBS 0.007414f
C66 B.n38 VSUBS 0.006977f
C67 B.n39 VSUBS 0.007414f
C68 B.t7 VSUBS 0.640922f
C69 B.t8 VSUBS 0.645771f
C70 B.t6 VSUBS 0.160616f
C71 B.n40 VSUBS 0.110268f
C72 B.n41 VSUBS 0.065908f
C73 B.n42 VSUBS 0.017176f
C74 B.n43 VSUBS 0.007414f
C75 B.n44 VSUBS 0.007414f
C76 B.n45 VSUBS 0.007414f
C77 B.n46 VSUBS 0.007414f
C78 B.t1 VSUBS 0.640899f
C79 B.t2 VSUBS 0.645749f
C80 B.t0 VSUBS 0.160616f
C81 B.n47 VSUBS 0.11029f
C82 B.n48 VSUBS 0.065931f
C83 B.n49 VSUBS 0.007414f
C84 B.n50 VSUBS 0.007414f
C85 B.n51 VSUBS 0.007414f
C86 B.n52 VSUBS 0.007414f
C87 B.n53 VSUBS 0.007414f
C88 B.n54 VSUBS 0.007414f
C89 B.n55 VSUBS 0.007414f
C90 B.n56 VSUBS 0.007414f
C91 B.n57 VSUBS 0.007414f
C92 B.n58 VSUBS 0.007414f
C93 B.n59 VSUBS 0.007414f
C94 B.n60 VSUBS 0.007414f
C95 B.n61 VSUBS 0.007414f
C96 B.n62 VSUBS 0.007414f
C97 B.n63 VSUBS 0.007414f
C98 B.n64 VSUBS 0.007414f
C99 B.n65 VSUBS 0.007414f
C100 B.n66 VSUBS 0.007414f
C101 B.n67 VSUBS 0.007414f
C102 B.n68 VSUBS 0.007414f
C103 B.n69 VSUBS 0.007414f
C104 B.n70 VSUBS 0.007414f
C105 B.n71 VSUBS 0.007414f
C106 B.n72 VSUBS 0.007414f
C107 B.n73 VSUBS 0.007414f
C108 B.n74 VSUBS 0.007414f
C109 B.n75 VSUBS 0.007414f
C110 B.n76 VSUBS 0.007414f
C111 B.n77 VSUBS 0.007414f
C112 B.n78 VSUBS 0.016402f
C113 B.n79 VSUBS 0.007414f
C114 B.n80 VSUBS 0.007414f
C115 B.n81 VSUBS 0.007414f
C116 B.n82 VSUBS 0.007414f
C117 B.n83 VSUBS 0.007414f
C118 B.n84 VSUBS 0.007414f
C119 B.n85 VSUBS 0.007414f
C120 B.n86 VSUBS 0.007414f
C121 B.n87 VSUBS 0.007414f
C122 B.n88 VSUBS 0.007414f
C123 B.n89 VSUBS 0.007414f
C124 B.n90 VSUBS 0.007414f
C125 B.n91 VSUBS 0.007414f
C126 B.n92 VSUBS 0.007414f
C127 B.n93 VSUBS 0.01671f
C128 B.n94 VSUBS 0.007414f
C129 B.n95 VSUBS 0.007414f
C130 B.n96 VSUBS 0.007414f
C131 B.n97 VSUBS 0.007414f
C132 B.n98 VSUBS 0.007414f
C133 B.n99 VSUBS 0.007414f
C134 B.n100 VSUBS 0.007414f
C135 B.n101 VSUBS 0.007414f
C136 B.n102 VSUBS 0.007414f
C137 B.n103 VSUBS 0.007414f
C138 B.n104 VSUBS 0.007414f
C139 B.n105 VSUBS 0.007414f
C140 B.n106 VSUBS 0.007414f
C141 B.n107 VSUBS 0.007414f
C142 B.n108 VSUBS 0.007414f
C143 B.n109 VSUBS 0.007414f
C144 B.n110 VSUBS 0.007414f
C145 B.n111 VSUBS 0.007414f
C146 B.n112 VSUBS 0.007414f
C147 B.n113 VSUBS 0.007414f
C148 B.n114 VSUBS 0.007414f
C149 B.n115 VSUBS 0.007414f
C150 B.n116 VSUBS 0.007414f
C151 B.n117 VSUBS 0.007414f
C152 B.n118 VSUBS 0.007414f
C153 B.n119 VSUBS 0.007414f
C154 B.n120 VSUBS 0.007414f
C155 B.n121 VSUBS 0.007414f
C156 B.n122 VSUBS 0.007414f
C157 B.t5 VSUBS 0.640899f
C158 B.t4 VSUBS 0.645749f
C159 B.t3 VSUBS 0.160616f
C160 B.n123 VSUBS 0.11029f
C161 B.n124 VSUBS 0.065931f
C162 B.n125 VSUBS 0.007414f
C163 B.n126 VSUBS 0.007414f
C164 B.n127 VSUBS 0.007414f
C165 B.n128 VSUBS 0.007414f
C166 B.n129 VSUBS 0.004143f
C167 B.n130 VSUBS 0.007414f
C168 B.n131 VSUBS 0.007414f
C169 B.n132 VSUBS 0.007414f
C170 B.n133 VSUBS 0.007414f
C171 B.n134 VSUBS 0.007414f
C172 B.n135 VSUBS 0.007414f
C173 B.n136 VSUBS 0.007414f
C174 B.n137 VSUBS 0.007414f
C175 B.n138 VSUBS 0.007414f
C176 B.n139 VSUBS 0.007414f
C177 B.n140 VSUBS 0.007414f
C178 B.n141 VSUBS 0.007414f
C179 B.n142 VSUBS 0.007414f
C180 B.n143 VSUBS 0.007414f
C181 B.n144 VSUBS 0.007414f
C182 B.n145 VSUBS 0.007414f
C183 B.n146 VSUBS 0.007414f
C184 B.n147 VSUBS 0.007414f
C185 B.n148 VSUBS 0.007414f
C186 B.n149 VSUBS 0.007414f
C187 B.n150 VSUBS 0.007414f
C188 B.n151 VSUBS 0.007414f
C189 B.n152 VSUBS 0.007414f
C190 B.n153 VSUBS 0.007414f
C191 B.n154 VSUBS 0.007414f
C192 B.n155 VSUBS 0.007414f
C193 B.n156 VSUBS 0.007414f
C194 B.n157 VSUBS 0.007414f
C195 B.n158 VSUBS 0.007414f
C196 B.n159 VSUBS 0.016402f
C197 B.n160 VSUBS 0.007414f
C198 B.n161 VSUBS 0.007414f
C199 B.n162 VSUBS 0.007414f
C200 B.n163 VSUBS 0.007414f
C201 B.n164 VSUBS 0.007414f
C202 B.n165 VSUBS 0.007414f
C203 B.n166 VSUBS 0.007414f
C204 B.n167 VSUBS 0.007414f
C205 B.n168 VSUBS 0.007414f
C206 B.n169 VSUBS 0.007414f
C207 B.n170 VSUBS 0.007414f
C208 B.n171 VSUBS 0.007414f
C209 B.n172 VSUBS 0.007414f
C210 B.n173 VSUBS 0.007414f
C211 B.n174 VSUBS 0.007414f
C212 B.n175 VSUBS 0.007414f
C213 B.n176 VSUBS 0.007414f
C214 B.n177 VSUBS 0.007414f
C215 B.n178 VSUBS 0.007414f
C216 B.n179 VSUBS 0.007414f
C217 B.n180 VSUBS 0.007414f
C218 B.n181 VSUBS 0.007414f
C219 B.n182 VSUBS 0.007414f
C220 B.n183 VSUBS 0.007414f
C221 B.n184 VSUBS 0.016402f
C222 B.n185 VSUBS 0.017613f
C223 B.n186 VSUBS 0.017613f
C224 B.n187 VSUBS 0.007414f
C225 B.n188 VSUBS 0.007414f
C226 B.n189 VSUBS 0.007414f
C227 B.n190 VSUBS 0.007414f
C228 B.n191 VSUBS 0.007414f
C229 B.n192 VSUBS 0.007414f
C230 B.n193 VSUBS 0.007414f
C231 B.n194 VSUBS 0.007414f
C232 B.n195 VSUBS 0.007414f
C233 B.n196 VSUBS 0.007414f
C234 B.n197 VSUBS 0.007414f
C235 B.n198 VSUBS 0.007414f
C236 B.n199 VSUBS 0.007414f
C237 B.n200 VSUBS 0.007414f
C238 B.n201 VSUBS 0.007414f
C239 B.n202 VSUBS 0.007414f
C240 B.n203 VSUBS 0.007414f
C241 B.n204 VSUBS 0.007414f
C242 B.n205 VSUBS 0.007414f
C243 B.n206 VSUBS 0.007414f
C244 B.n207 VSUBS 0.007414f
C245 B.n208 VSUBS 0.007414f
C246 B.n209 VSUBS 0.007414f
C247 B.n210 VSUBS 0.007414f
C248 B.n211 VSUBS 0.007414f
C249 B.n212 VSUBS 0.007414f
C250 B.n213 VSUBS 0.007414f
C251 B.n214 VSUBS 0.007414f
C252 B.n215 VSUBS 0.007414f
C253 B.n216 VSUBS 0.007414f
C254 B.n217 VSUBS 0.007414f
C255 B.n218 VSUBS 0.007414f
C256 B.n219 VSUBS 0.007414f
C257 B.n220 VSUBS 0.007414f
C258 B.n221 VSUBS 0.007414f
C259 B.n222 VSUBS 0.007414f
C260 B.n223 VSUBS 0.007414f
C261 B.n224 VSUBS 0.007414f
C262 B.n225 VSUBS 0.007414f
C263 B.n226 VSUBS 0.007414f
C264 B.n227 VSUBS 0.007414f
C265 B.n228 VSUBS 0.007414f
C266 B.n229 VSUBS 0.007414f
C267 B.n230 VSUBS 0.007414f
C268 B.n231 VSUBS 0.007414f
C269 B.n232 VSUBS 0.007414f
C270 B.n233 VSUBS 0.007414f
C271 B.n234 VSUBS 0.007414f
C272 B.n235 VSUBS 0.007414f
C273 B.n236 VSUBS 0.007414f
C274 B.n237 VSUBS 0.007414f
C275 B.n238 VSUBS 0.007414f
C276 B.n239 VSUBS 0.007414f
C277 B.n240 VSUBS 0.007414f
C278 B.n241 VSUBS 0.007414f
C279 B.n242 VSUBS 0.007414f
C280 B.n243 VSUBS 0.007414f
C281 B.n244 VSUBS 0.007414f
C282 B.n245 VSUBS 0.007414f
C283 B.n246 VSUBS 0.007414f
C284 B.n247 VSUBS 0.007414f
C285 B.n248 VSUBS 0.007414f
C286 B.n249 VSUBS 0.007414f
C287 B.n250 VSUBS 0.007414f
C288 B.n251 VSUBS 0.007414f
C289 B.n252 VSUBS 0.007414f
C290 B.n253 VSUBS 0.007414f
C291 B.n254 VSUBS 0.007414f
C292 B.n255 VSUBS 0.007414f
C293 B.n256 VSUBS 0.007414f
C294 B.n257 VSUBS 0.007414f
C295 B.n258 VSUBS 0.007414f
C296 B.n259 VSUBS 0.007414f
C297 B.n260 VSUBS 0.007414f
C298 B.n261 VSUBS 0.007414f
C299 B.n262 VSUBS 0.007414f
C300 B.n263 VSUBS 0.007414f
C301 B.n264 VSUBS 0.007414f
C302 B.n265 VSUBS 0.007414f
C303 B.n266 VSUBS 0.007414f
C304 B.n267 VSUBS 0.007414f
C305 B.n268 VSUBS 0.007414f
C306 B.n269 VSUBS 0.007414f
C307 B.n270 VSUBS 0.007414f
C308 B.n271 VSUBS 0.007414f
C309 B.t11 VSUBS 0.640922f
C310 B.t10 VSUBS 0.645771f
C311 B.t9 VSUBS 0.160616f
C312 B.n272 VSUBS 0.110268f
C313 B.n273 VSUBS 0.065908f
C314 B.n274 VSUBS 0.017176f
C315 B.n275 VSUBS 0.006977f
C316 B.n276 VSUBS 0.007414f
C317 B.n277 VSUBS 0.007414f
C318 B.n278 VSUBS 0.007414f
C319 B.n279 VSUBS 0.007414f
C320 B.n280 VSUBS 0.007414f
C321 B.n281 VSUBS 0.007414f
C322 B.n282 VSUBS 0.007414f
C323 B.n283 VSUBS 0.007414f
C324 B.n284 VSUBS 0.007414f
C325 B.n285 VSUBS 0.007414f
C326 B.n286 VSUBS 0.007414f
C327 B.n287 VSUBS 0.007414f
C328 B.n288 VSUBS 0.007414f
C329 B.n289 VSUBS 0.007414f
C330 B.n290 VSUBS 0.007414f
C331 B.n291 VSUBS 0.004143f
C332 B.n292 VSUBS 0.017176f
C333 B.n293 VSUBS 0.006977f
C334 B.n294 VSUBS 0.007414f
C335 B.n295 VSUBS 0.007414f
C336 B.n296 VSUBS 0.007414f
C337 B.n297 VSUBS 0.007414f
C338 B.n298 VSUBS 0.007414f
C339 B.n299 VSUBS 0.007414f
C340 B.n300 VSUBS 0.007414f
C341 B.n301 VSUBS 0.007414f
C342 B.n302 VSUBS 0.007414f
C343 B.n303 VSUBS 0.007414f
C344 B.n304 VSUBS 0.007414f
C345 B.n305 VSUBS 0.007414f
C346 B.n306 VSUBS 0.007414f
C347 B.n307 VSUBS 0.007414f
C348 B.n308 VSUBS 0.007414f
C349 B.n309 VSUBS 0.007414f
C350 B.n310 VSUBS 0.007414f
C351 B.n311 VSUBS 0.007414f
C352 B.n312 VSUBS 0.007414f
C353 B.n313 VSUBS 0.007414f
C354 B.n314 VSUBS 0.007414f
C355 B.n315 VSUBS 0.007414f
C356 B.n316 VSUBS 0.007414f
C357 B.n317 VSUBS 0.007414f
C358 B.n318 VSUBS 0.007414f
C359 B.n319 VSUBS 0.007414f
C360 B.n320 VSUBS 0.007414f
C361 B.n321 VSUBS 0.007414f
C362 B.n322 VSUBS 0.007414f
C363 B.n323 VSUBS 0.007414f
C364 B.n324 VSUBS 0.007414f
C365 B.n325 VSUBS 0.007414f
C366 B.n326 VSUBS 0.007414f
C367 B.n327 VSUBS 0.007414f
C368 B.n328 VSUBS 0.007414f
C369 B.n329 VSUBS 0.007414f
C370 B.n330 VSUBS 0.007414f
C371 B.n331 VSUBS 0.007414f
C372 B.n332 VSUBS 0.007414f
C373 B.n333 VSUBS 0.007414f
C374 B.n334 VSUBS 0.007414f
C375 B.n335 VSUBS 0.007414f
C376 B.n336 VSUBS 0.007414f
C377 B.n337 VSUBS 0.007414f
C378 B.n338 VSUBS 0.007414f
C379 B.n339 VSUBS 0.007414f
C380 B.n340 VSUBS 0.007414f
C381 B.n341 VSUBS 0.007414f
C382 B.n342 VSUBS 0.007414f
C383 B.n343 VSUBS 0.007414f
C384 B.n344 VSUBS 0.007414f
C385 B.n345 VSUBS 0.007414f
C386 B.n346 VSUBS 0.007414f
C387 B.n347 VSUBS 0.007414f
C388 B.n348 VSUBS 0.007414f
C389 B.n349 VSUBS 0.007414f
C390 B.n350 VSUBS 0.007414f
C391 B.n351 VSUBS 0.007414f
C392 B.n352 VSUBS 0.007414f
C393 B.n353 VSUBS 0.007414f
C394 B.n354 VSUBS 0.007414f
C395 B.n355 VSUBS 0.007414f
C396 B.n356 VSUBS 0.007414f
C397 B.n357 VSUBS 0.007414f
C398 B.n358 VSUBS 0.007414f
C399 B.n359 VSUBS 0.007414f
C400 B.n360 VSUBS 0.007414f
C401 B.n361 VSUBS 0.007414f
C402 B.n362 VSUBS 0.007414f
C403 B.n363 VSUBS 0.007414f
C404 B.n364 VSUBS 0.007414f
C405 B.n365 VSUBS 0.007414f
C406 B.n366 VSUBS 0.007414f
C407 B.n367 VSUBS 0.007414f
C408 B.n368 VSUBS 0.007414f
C409 B.n369 VSUBS 0.007414f
C410 B.n370 VSUBS 0.007414f
C411 B.n371 VSUBS 0.007414f
C412 B.n372 VSUBS 0.007414f
C413 B.n373 VSUBS 0.007414f
C414 B.n374 VSUBS 0.007414f
C415 B.n375 VSUBS 0.007414f
C416 B.n376 VSUBS 0.007414f
C417 B.n377 VSUBS 0.007414f
C418 B.n378 VSUBS 0.007414f
C419 B.n379 VSUBS 0.007414f
C420 B.n380 VSUBS 0.017613f
C421 B.n381 VSUBS 0.016402f
C422 B.n382 VSUBS 0.017305f
C423 B.n383 VSUBS 0.007414f
C424 B.n384 VSUBS 0.007414f
C425 B.n385 VSUBS 0.007414f
C426 B.n386 VSUBS 0.007414f
C427 B.n387 VSUBS 0.007414f
C428 B.n388 VSUBS 0.007414f
C429 B.n389 VSUBS 0.007414f
C430 B.n390 VSUBS 0.007414f
C431 B.n391 VSUBS 0.007414f
C432 B.n392 VSUBS 0.007414f
C433 B.n393 VSUBS 0.007414f
C434 B.n394 VSUBS 0.007414f
C435 B.n395 VSUBS 0.007414f
C436 B.n396 VSUBS 0.007414f
C437 B.n397 VSUBS 0.007414f
C438 B.n398 VSUBS 0.007414f
C439 B.n399 VSUBS 0.007414f
C440 B.n400 VSUBS 0.007414f
C441 B.n401 VSUBS 0.007414f
C442 B.n402 VSUBS 0.007414f
C443 B.n403 VSUBS 0.007414f
C444 B.n404 VSUBS 0.007414f
C445 B.n405 VSUBS 0.007414f
C446 B.n406 VSUBS 0.007414f
C447 B.n407 VSUBS 0.007414f
C448 B.n408 VSUBS 0.007414f
C449 B.n409 VSUBS 0.007414f
C450 B.n410 VSUBS 0.007414f
C451 B.n411 VSUBS 0.007414f
C452 B.n412 VSUBS 0.007414f
C453 B.n413 VSUBS 0.007414f
C454 B.n414 VSUBS 0.007414f
C455 B.n415 VSUBS 0.007414f
C456 B.n416 VSUBS 0.007414f
C457 B.n417 VSUBS 0.007414f
C458 B.n418 VSUBS 0.007414f
C459 B.n419 VSUBS 0.007414f
C460 B.n420 VSUBS 0.007414f
C461 B.n421 VSUBS 0.007414f
C462 B.n422 VSUBS 0.007414f
C463 B.n423 VSUBS 0.007414f
C464 B.n424 VSUBS 0.007414f
C465 B.n425 VSUBS 0.016402f
C466 B.n426 VSUBS 0.017613f
C467 B.n427 VSUBS 0.017613f
C468 B.n428 VSUBS 0.007414f
C469 B.n429 VSUBS 0.007414f
C470 B.n430 VSUBS 0.007414f
C471 B.n431 VSUBS 0.007414f
C472 B.n432 VSUBS 0.007414f
C473 B.n433 VSUBS 0.007414f
C474 B.n434 VSUBS 0.007414f
C475 B.n435 VSUBS 0.007414f
C476 B.n436 VSUBS 0.007414f
C477 B.n437 VSUBS 0.007414f
C478 B.n438 VSUBS 0.007414f
C479 B.n439 VSUBS 0.007414f
C480 B.n440 VSUBS 0.007414f
C481 B.n441 VSUBS 0.007414f
C482 B.n442 VSUBS 0.007414f
C483 B.n443 VSUBS 0.007414f
C484 B.n444 VSUBS 0.007414f
C485 B.n445 VSUBS 0.007414f
C486 B.n446 VSUBS 0.007414f
C487 B.n447 VSUBS 0.007414f
C488 B.n448 VSUBS 0.007414f
C489 B.n449 VSUBS 0.007414f
C490 B.n450 VSUBS 0.007414f
C491 B.n451 VSUBS 0.007414f
C492 B.n452 VSUBS 0.007414f
C493 B.n453 VSUBS 0.007414f
C494 B.n454 VSUBS 0.007414f
C495 B.n455 VSUBS 0.007414f
C496 B.n456 VSUBS 0.007414f
C497 B.n457 VSUBS 0.007414f
C498 B.n458 VSUBS 0.007414f
C499 B.n459 VSUBS 0.007414f
C500 B.n460 VSUBS 0.007414f
C501 B.n461 VSUBS 0.007414f
C502 B.n462 VSUBS 0.007414f
C503 B.n463 VSUBS 0.007414f
C504 B.n464 VSUBS 0.007414f
C505 B.n465 VSUBS 0.007414f
C506 B.n466 VSUBS 0.007414f
C507 B.n467 VSUBS 0.007414f
C508 B.n468 VSUBS 0.007414f
C509 B.n469 VSUBS 0.007414f
C510 B.n470 VSUBS 0.007414f
C511 B.n471 VSUBS 0.007414f
C512 B.n472 VSUBS 0.007414f
C513 B.n473 VSUBS 0.007414f
C514 B.n474 VSUBS 0.007414f
C515 B.n475 VSUBS 0.007414f
C516 B.n476 VSUBS 0.007414f
C517 B.n477 VSUBS 0.007414f
C518 B.n478 VSUBS 0.007414f
C519 B.n479 VSUBS 0.007414f
C520 B.n480 VSUBS 0.007414f
C521 B.n481 VSUBS 0.007414f
C522 B.n482 VSUBS 0.007414f
C523 B.n483 VSUBS 0.007414f
C524 B.n484 VSUBS 0.007414f
C525 B.n485 VSUBS 0.007414f
C526 B.n486 VSUBS 0.007414f
C527 B.n487 VSUBS 0.007414f
C528 B.n488 VSUBS 0.007414f
C529 B.n489 VSUBS 0.007414f
C530 B.n490 VSUBS 0.007414f
C531 B.n491 VSUBS 0.007414f
C532 B.n492 VSUBS 0.007414f
C533 B.n493 VSUBS 0.007414f
C534 B.n494 VSUBS 0.007414f
C535 B.n495 VSUBS 0.007414f
C536 B.n496 VSUBS 0.007414f
C537 B.n497 VSUBS 0.007414f
C538 B.n498 VSUBS 0.007414f
C539 B.n499 VSUBS 0.007414f
C540 B.n500 VSUBS 0.007414f
C541 B.n501 VSUBS 0.007414f
C542 B.n502 VSUBS 0.007414f
C543 B.n503 VSUBS 0.007414f
C544 B.n504 VSUBS 0.007414f
C545 B.n505 VSUBS 0.007414f
C546 B.n506 VSUBS 0.007414f
C547 B.n507 VSUBS 0.007414f
C548 B.n508 VSUBS 0.007414f
C549 B.n509 VSUBS 0.007414f
C550 B.n510 VSUBS 0.007414f
C551 B.n511 VSUBS 0.007414f
C552 B.n512 VSUBS 0.007414f
C553 B.n513 VSUBS 0.007414f
C554 B.n514 VSUBS 0.006977f
C555 B.n515 VSUBS 0.017176f
C556 B.n516 VSUBS 0.004143f
C557 B.n517 VSUBS 0.007414f
C558 B.n518 VSUBS 0.007414f
C559 B.n519 VSUBS 0.007414f
C560 B.n520 VSUBS 0.007414f
C561 B.n521 VSUBS 0.007414f
C562 B.n522 VSUBS 0.007414f
C563 B.n523 VSUBS 0.007414f
C564 B.n524 VSUBS 0.007414f
C565 B.n525 VSUBS 0.007414f
C566 B.n526 VSUBS 0.007414f
C567 B.n527 VSUBS 0.007414f
C568 B.n528 VSUBS 0.007414f
C569 B.n529 VSUBS 0.004143f
C570 B.n530 VSUBS 0.007414f
C571 B.n531 VSUBS 0.007414f
C572 B.n532 VSUBS 0.007414f
C573 B.n533 VSUBS 0.007414f
C574 B.n534 VSUBS 0.007414f
C575 B.n535 VSUBS 0.007414f
C576 B.n536 VSUBS 0.007414f
C577 B.n537 VSUBS 0.007414f
C578 B.n538 VSUBS 0.007414f
C579 B.n539 VSUBS 0.007414f
C580 B.n540 VSUBS 0.007414f
C581 B.n541 VSUBS 0.007414f
C582 B.n542 VSUBS 0.007414f
C583 B.n543 VSUBS 0.007414f
C584 B.n544 VSUBS 0.007414f
C585 B.n545 VSUBS 0.007414f
C586 B.n546 VSUBS 0.007414f
C587 B.n547 VSUBS 0.007414f
C588 B.n548 VSUBS 0.007414f
C589 B.n549 VSUBS 0.007414f
C590 B.n550 VSUBS 0.007414f
C591 B.n551 VSUBS 0.007414f
C592 B.n552 VSUBS 0.007414f
C593 B.n553 VSUBS 0.007414f
C594 B.n554 VSUBS 0.007414f
C595 B.n555 VSUBS 0.007414f
C596 B.n556 VSUBS 0.007414f
C597 B.n557 VSUBS 0.007414f
C598 B.n558 VSUBS 0.007414f
C599 B.n559 VSUBS 0.007414f
C600 B.n560 VSUBS 0.007414f
C601 B.n561 VSUBS 0.007414f
C602 B.n562 VSUBS 0.007414f
C603 B.n563 VSUBS 0.007414f
C604 B.n564 VSUBS 0.007414f
C605 B.n565 VSUBS 0.007414f
C606 B.n566 VSUBS 0.007414f
C607 B.n567 VSUBS 0.007414f
C608 B.n568 VSUBS 0.007414f
C609 B.n569 VSUBS 0.007414f
C610 B.n570 VSUBS 0.007414f
C611 B.n571 VSUBS 0.007414f
C612 B.n572 VSUBS 0.007414f
C613 B.n573 VSUBS 0.007414f
C614 B.n574 VSUBS 0.007414f
C615 B.n575 VSUBS 0.007414f
C616 B.n576 VSUBS 0.007414f
C617 B.n577 VSUBS 0.007414f
C618 B.n578 VSUBS 0.007414f
C619 B.n579 VSUBS 0.007414f
C620 B.n580 VSUBS 0.007414f
C621 B.n581 VSUBS 0.007414f
C622 B.n582 VSUBS 0.007414f
C623 B.n583 VSUBS 0.007414f
C624 B.n584 VSUBS 0.007414f
C625 B.n585 VSUBS 0.007414f
C626 B.n586 VSUBS 0.007414f
C627 B.n587 VSUBS 0.007414f
C628 B.n588 VSUBS 0.007414f
C629 B.n589 VSUBS 0.007414f
C630 B.n590 VSUBS 0.007414f
C631 B.n591 VSUBS 0.007414f
C632 B.n592 VSUBS 0.007414f
C633 B.n593 VSUBS 0.007414f
C634 B.n594 VSUBS 0.007414f
C635 B.n595 VSUBS 0.007414f
C636 B.n596 VSUBS 0.007414f
C637 B.n597 VSUBS 0.007414f
C638 B.n598 VSUBS 0.007414f
C639 B.n599 VSUBS 0.007414f
C640 B.n600 VSUBS 0.007414f
C641 B.n601 VSUBS 0.007414f
C642 B.n602 VSUBS 0.007414f
C643 B.n603 VSUBS 0.007414f
C644 B.n604 VSUBS 0.007414f
C645 B.n605 VSUBS 0.007414f
C646 B.n606 VSUBS 0.007414f
C647 B.n607 VSUBS 0.007414f
C648 B.n608 VSUBS 0.007414f
C649 B.n609 VSUBS 0.007414f
C650 B.n610 VSUBS 0.007414f
C651 B.n611 VSUBS 0.007414f
C652 B.n612 VSUBS 0.007414f
C653 B.n613 VSUBS 0.007414f
C654 B.n614 VSUBS 0.007414f
C655 B.n615 VSUBS 0.007414f
C656 B.n616 VSUBS 0.007414f
C657 B.n617 VSUBS 0.007414f
C658 B.n618 VSUBS 0.017613f
C659 B.n619 VSUBS 0.016402f
C660 B.n620 VSUBS 0.016402f
C661 B.n621 VSUBS 0.007414f
C662 B.n622 VSUBS 0.007414f
C663 B.n623 VSUBS 0.007414f
C664 B.n624 VSUBS 0.007414f
C665 B.n625 VSUBS 0.007414f
C666 B.n626 VSUBS 0.007414f
C667 B.n627 VSUBS 0.007414f
C668 B.n628 VSUBS 0.007414f
C669 B.n629 VSUBS 0.007414f
C670 B.n630 VSUBS 0.007414f
C671 B.n631 VSUBS 0.007414f
C672 B.n632 VSUBS 0.007414f
C673 B.n633 VSUBS 0.007414f
C674 B.n634 VSUBS 0.007414f
C675 B.n635 VSUBS 0.007414f
C676 B.n636 VSUBS 0.007414f
C677 B.n637 VSUBS 0.007414f
C678 B.n638 VSUBS 0.007414f
C679 B.n639 VSUBS 0.009674f
C680 B.n640 VSUBS 0.010306f
C681 B.n641 VSUBS 0.020494f
C682 VDD2.t5 VSUBS 5.05001f
C683 VDD2.t1 VSUBS 0.467854f
C684 VDD2.t2 VSUBS 0.467854f
C685 VDD2.n0 VSUBS 3.8902f
C686 VDD2.n1 VSUBS 3.73777f
C687 VDD2.t4 VSUBS 5.04663f
C688 VDD2.n2 VSUBS 3.84762f
C689 VDD2.t0 VSUBS 0.467854f
C690 VDD2.t3 VSUBS 0.467854f
C691 VDD2.n3 VSUBS 3.89015f
C692 VN.t0 VSUBS 0.82017f
C693 VN.n0 VSUBS 0.333151f
C694 VN.t4 VSUBS 0.813798f
C695 VN.n1 VSUBS 0.311981f
C696 VN.t3 VSUBS 0.82017f
C697 VN.n2 VSUBS 0.333048f
C698 VN.n3 VSUBS 0.144255f
C699 VN.t2 VSUBS 0.82017f
C700 VN.n4 VSUBS 0.333151f
C701 VN.t1 VSUBS 0.82017f
C702 VN.t5 VSUBS 0.813798f
C703 VN.n5 VSUBS 0.311981f
C704 VN.n6 VSUBS 0.333048f
C705 VN.n7 VSUBS 3.38419f
C706 VDD1.t5 VSUBS 5.04742f
C707 VDD1.t3 VSUBS 5.04608f
C708 VDD1.t1 VSUBS 0.46749f
C709 VDD1.t0 VSUBS 0.46749f
C710 VDD1.n0 VSUBS 3.88718f
C711 VDD1.n1 VSUBS 3.82316f
C712 VDD1.t2 VSUBS 0.46749f
C713 VDD1.t4 VSUBS 0.46749f
C714 VDD1.n2 VSUBS 3.88651f
C715 VDD1.n3 VSUBS 3.77226f
C716 VTAIL.t5 VSUBS 0.498498f
C717 VTAIL.t2 VSUBS 0.498498f
C718 VTAIL.n0 VSUBS 3.93031f
C719 VTAIL.n1 VSUBS 0.954853f
C720 VTAIL.t7 VSUBS 5.13179f
C721 VTAIL.n2 VSUBS 1.14663f
C722 VTAIL.t11 VSUBS 0.498498f
C723 VTAIL.t6 VSUBS 0.498498f
C724 VTAIL.n3 VSUBS 3.93031f
C725 VTAIL.n4 VSUBS 3.24615f
C726 VTAIL.t4 VSUBS 0.498498f
C727 VTAIL.t3 VSUBS 0.498498f
C728 VTAIL.n5 VSUBS 3.93032f
C729 VTAIL.n6 VSUBS 3.24614f
C730 VTAIL.t0 VSUBS 5.1318f
C731 VTAIL.n7 VSUBS 1.14662f
C732 VTAIL.t8 VSUBS 0.498498f
C733 VTAIL.t9 VSUBS 0.498498f
C734 VTAIL.n8 VSUBS 3.93032f
C735 VTAIL.n9 VSUBS 0.988561f
C736 VTAIL.t10 VSUBS 5.13179f
C737 VTAIL.n10 VSUBS 3.35046f
C738 VTAIL.t1 VSUBS 5.13179f
C739 VTAIL.n11 VSUBS 3.33042f
C740 VP.t0 VSUBS 0.844472f
C741 VP.n0 VSUBS 0.343023f
C742 VP.t3 VSUBS 0.837911f
C743 VP.n1 VSUBS 0.321225f
C744 VP.t1 VSUBS 0.844472f
C745 VP.n2 VSUBS 0.342917f
C746 VP.n3 VSUBS 3.43512f
C747 VP.n4 VSUBS 3.40671f
C748 VP.t4 VSUBS 0.837911f
C749 VP.t2 VSUBS 0.844472f
C750 VP.n5 VSUBS 0.342917f
C751 VP.n6 VSUBS 0.321225f
C752 VP.t5 VSUBS 0.844472f
C753 VP.n7 VSUBS 0.342917f
C754 VP.n8 VSUBS 0.058403f
.ends

