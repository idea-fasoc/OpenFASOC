* NGSPICE file created from diff_pair_sample_0939.ext - technology: sky130A

.subckt diff_pair_sample_0939 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t3 VP.t0 VTAIL.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=0.1815 pd=1.43 as=0.429 ps=2.98 w=1.1 l=3.6
X1 B.t17 B.t15 B.t16 B.t5 sky130_fd_pr__nfet_01v8 ad=0.429 pd=2.98 as=0 ps=0 w=1.1 l=3.6
X2 VTAIL.t1 VN.t0 VDD2.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=0.429 pd=2.98 as=0.1815 ps=1.43 w=1.1 l=3.6
X3 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=0.429 pd=2.98 as=0 ps=0 w=1.1 l=3.6
X4 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=0.429 pd=2.98 as=0 ps=0 w=1.1 l=3.6
X5 VDD2.t2 VN.t1 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.1815 pd=1.43 as=0.429 ps=2.98 w=1.1 l=3.6
X6 VDD1.t2 VP.t1 VTAIL.t7 B.t2 sky130_fd_pr__nfet_01v8 ad=0.1815 pd=1.43 as=0.429 ps=2.98 w=1.1 l=3.6
X7 VDD2.t1 VN.t2 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.1815 pd=1.43 as=0.429 ps=2.98 w=1.1 l=3.6
X8 VTAIL.t6 VP.t2 VDD1.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=0.429 pd=2.98 as=0.1815 ps=1.43 w=1.1 l=3.6
X9 VTAIL.t0 VN.t3 VDD2.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.429 pd=2.98 as=0.1815 ps=1.43 w=1.1 l=3.6
X10 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=0.429 pd=2.98 as=0 ps=0 w=1.1 l=3.6
X11 VTAIL.t5 VP.t3 VDD1.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=0.429 pd=2.98 as=0.1815 ps=1.43 w=1.1 l=3.6
R0 VP.n19 VP.n18 161.3
R1 VP.n17 VP.n1 161.3
R2 VP.n16 VP.n15 161.3
R3 VP.n14 VP.n2 161.3
R4 VP.n13 VP.n12 161.3
R5 VP.n11 VP.n3 161.3
R6 VP.n10 VP.n9 161.3
R7 VP.n8 VP.n4 161.3
R8 VP.n7 VP.n6 79.4233
R9 VP.n20 VP.n0 79.4233
R10 VP.n12 VP.n2 56.4773
R11 VP.n7 VP.n5 43.3237
R12 VP.n5 VP.t3 42.158
R13 VP.n5 VP.t0 40.9152
R14 VP.n10 VP.n4 24.3439
R15 VP.n11 VP.n10 24.3439
R16 VP.n12 VP.n11 24.3439
R17 VP.n16 VP.n2 24.3439
R18 VP.n17 VP.n16 24.3439
R19 VP.n18 VP.n17 24.3439
R20 VP.n6 VP.n4 10.4682
R21 VP.n18 VP.n0 10.4682
R22 VP.n6 VP.t2 7.36439
R23 VP.n0 VP.t1 7.36439
R24 VP.n8 VP.n7 0.355081
R25 VP.n20 VP.n19 0.355081
R26 VP VP.n20 0.26685
R27 VP.n9 VP.n8 0.189894
R28 VP.n9 VP.n3 0.189894
R29 VP.n13 VP.n3 0.189894
R30 VP.n14 VP.n13 0.189894
R31 VP.n15 VP.n14 0.189894
R32 VP.n15 VP.n1 0.189894
R33 VP.n19 VP.n1 0.189894
R34 VTAIL.n7 VTAIL.t3 155.721
R35 VTAIL.n0 VTAIL.t1 155.721
R36 VTAIL.n1 VTAIL.t7 155.721
R37 VTAIL.n2 VTAIL.t6 155.721
R38 VTAIL.n6 VTAIL.t4 155.721
R39 VTAIL.n5 VTAIL.t5 155.721
R40 VTAIL.n4 VTAIL.t2 155.721
R41 VTAIL.n3 VTAIL.t0 155.721
R42 VTAIL.n7 VTAIL.n6 16.7031
R43 VTAIL.n3 VTAIL.n2 16.7031
R44 VTAIL.n4 VTAIL.n3 3.38843
R45 VTAIL.n6 VTAIL.n5 3.38843
R46 VTAIL.n2 VTAIL.n1 3.38843
R47 VTAIL VTAIL.n0 1.75266
R48 VTAIL VTAIL.n7 1.63628
R49 VTAIL.n5 VTAIL.n4 0.470328
R50 VTAIL.n1 VTAIL.n0 0.470328
R51 VDD1 VDD1.n1 181.589
R52 VDD1 VDD1.n0 146.297
R53 VDD1.n0 VDD1.t0 18.0005
R54 VDD1.n0 VDD1.t3 18.0005
R55 VDD1.n1 VDD1.t1 18.0005
R56 VDD1.n1 VDD1.t2 18.0005
R57 B.n500 B.n499 585
R58 B.n501 B.n500 585
R59 B.n153 B.n95 585
R60 B.n152 B.n151 585
R61 B.n150 B.n149 585
R62 B.n148 B.n147 585
R63 B.n146 B.n145 585
R64 B.n144 B.n143 585
R65 B.n142 B.n141 585
R66 B.n140 B.n139 585
R67 B.n138 B.n137 585
R68 B.n135 B.n134 585
R69 B.n133 B.n132 585
R70 B.n131 B.n130 585
R71 B.n129 B.n128 585
R72 B.n127 B.n126 585
R73 B.n125 B.n124 585
R74 B.n123 B.n122 585
R75 B.n121 B.n120 585
R76 B.n119 B.n118 585
R77 B.n117 B.n116 585
R78 B.n115 B.n114 585
R79 B.n113 B.n112 585
R80 B.n111 B.n110 585
R81 B.n109 B.n108 585
R82 B.n107 B.n106 585
R83 B.n105 B.n104 585
R84 B.n103 B.n102 585
R85 B.n81 B.n80 585
R86 B.n504 B.n503 585
R87 B.n498 B.n96 585
R88 B.n96 B.n78 585
R89 B.n497 B.n77 585
R90 B.n508 B.n77 585
R91 B.n496 B.n76 585
R92 B.n509 B.n76 585
R93 B.n495 B.n75 585
R94 B.n510 B.n75 585
R95 B.n494 B.n493 585
R96 B.n493 B.n71 585
R97 B.n492 B.n70 585
R98 B.n516 B.n70 585
R99 B.n491 B.n69 585
R100 B.n517 B.n69 585
R101 B.n490 B.n68 585
R102 B.n518 B.n68 585
R103 B.n489 B.n488 585
R104 B.n488 B.n64 585
R105 B.n487 B.n63 585
R106 B.n524 B.n63 585
R107 B.n486 B.n62 585
R108 B.n525 B.n62 585
R109 B.n485 B.n61 585
R110 B.n526 B.n61 585
R111 B.n484 B.n483 585
R112 B.n483 B.n57 585
R113 B.n482 B.n56 585
R114 B.n532 B.n56 585
R115 B.n481 B.n55 585
R116 B.n533 B.n55 585
R117 B.n480 B.n54 585
R118 B.n534 B.n54 585
R119 B.n479 B.n478 585
R120 B.n478 B.n50 585
R121 B.n477 B.n49 585
R122 B.n540 B.n49 585
R123 B.n476 B.n48 585
R124 B.n541 B.n48 585
R125 B.n475 B.n47 585
R126 B.n542 B.n47 585
R127 B.n474 B.n473 585
R128 B.n473 B.n43 585
R129 B.n472 B.n42 585
R130 B.n548 B.n42 585
R131 B.n471 B.n41 585
R132 B.n549 B.n41 585
R133 B.n470 B.n40 585
R134 B.n550 B.n40 585
R135 B.n469 B.n468 585
R136 B.n468 B.n39 585
R137 B.n467 B.n35 585
R138 B.n556 B.n35 585
R139 B.n466 B.n34 585
R140 B.n557 B.n34 585
R141 B.n465 B.n33 585
R142 B.n558 B.n33 585
R143 B.n464 B.n463 585
R144 B.n463 B.n29 585
R145 B.n462 B.n28 585
R146 B.n564 B.n28 585
R147 B.n461 B.n27 585
R148 B.n565 B.n27 585
R149 B.n460 B.n26 585
R150 B.n566 B.n26 585
R151 B.n459 B.n458 585
R152 B.n458 B.n22 585
R153 B.n457 B.n21 585
R154 B.n572 B.n21 585
R155 B.n456 B.n20 585
R156 B.n573 B.n20 585
R157 B.n455 B.n19 585
R158 B.n574 B.n19 585
R159 B.n454 B.n453 585
R160 B.n453 B.n15 585
R161 B.n452 B.n14 585
R162 B.n580 B.n14 585
R163 B.n451 B.n13 585
R164 B.n581 B.n13 585
R165 B.n450 B.n12 585
R166 B.n582 B.n12 585
R167 B.n449 B.n448 585
R168 B.n448 B.n8 585
R169 B.n447 B.n7 585
R170 B.n588 B.n7 585
R171 B.n446 B.n6 585
R172 B.n589 B.n6 585
R173 B.n445 B.n5 585
R174 B.n590 B.n5 585
R175 B.n444 B.n443 585
R176 B.n443 B.n4 585
R177 B.n442 B.n154 585
R178 B.n442 B.n441 585
R179 B.n432 B.n155 585
R180 B.n156 B.n155 585
R181 B.n434 B.n433 585
R182 B.n435 B.n434 585
R183 B.n431 B.n161 585
R184 B.n161 B.n160 585
R185 B.n430 B.n429 585
R186 B.n429 B.n428 585
R187 B.n163 B.n162 585
R188 B.n164 B.n163 585
R189 B.n421 B.n420 585
R190 B.n422 B.n421 585
R191 B.n419 B.n169 585
R192 B.n169 B.n168 585
R193 B.n418 B.n417 585
R194 B.n417 B.n416 585
R195 B.n171 B.n170 585
R196 B.n172 B.n171 585
R197 B.n409 B.n408 585
R198 B.n410 B.n409 585
R199 B.n407 B.n177 585
R200 B.n177 B.n176 585
R201 B.n406 B.n405 585
R202 B.n405 B.n404 585
R203 B.n179 B.n178 585
R204 B.n180 B.n179 585
R205 B.n397 B.n396 585
R206 B.n398 B.n397 585
R207 B.n395 B.n185 585
R208 B.n185 B.n184 585
R209 B.n394 B.n393 585
R210 B.n393 B.n392 585
R211 B.n187 B.n186 585
R212 B.n385 B.n187 585
R213 B.n384 B.n383 585
R214 B.n386 B.n384 585
R215 B.n382 B.n192 585
R216 B.n192 B.n191 585
R217 B.n381 B.n380 585
R218 B.n380 B.n379 585
R219 B.n194 B.n193 585
R220 B.n195 B.n194 585
R221 B.n372 B.n371 585
R222 B.n373 B.n372 585
R223 B.n370 B.n200 585
R224 B.n200 B.n199 585
R225 B.n369 B.n368 585
R226 B.n368 B.n367 585
R227 B.n202 B.n201 585
R228 B.n203 B.n202 585
R229 B.n360 B.n359 585
R230 B.n361 B.n360 585
R231 B.n358 B.n208 585
R232 B.n208 B.n207 585
R233 B.n357 B.n356 585
R234 B.n356 B.n355 585
R235 B.n210 B.n209 585
R236 B.n211 B.n210 585
R237 B.n348 B.n347 585
R238 B.n349 B.n348 585
R239 B.n346 B.n216 585
R240 B.n216 B.n215 585
R241 B.n345 B.n344 585
R242 B.n344 B.n343 585
R243 B.n218 B.n217 585
R244 B.n219 B.n218 585
R245 B.n336 B.n335 585
R246 B.n337 B.n336 585
R247 B.n334 B.n224 585
R248 B.n224 B.n223 585
R249 B.n333 B.n332 585
R250 B.n332 B.n331 585
R251 B.n226 B.n225 585
R252 B.n227 B.n226 585
R253 B.n324 B.n323 585
R254 B.n325 B.n324 585
R255 B.n322 B.n232 585
R256 B.n232 B.n231 585
R257 B.n321 B.n320 585
R258 B.n320 B.n319 585
R259 B.n234 B.n233 585
R260 B.n235 B.n234 585
R261 B.n315 B.n314 585
R262 B.n238 B.n237 585
R263 B.n311 B.n310 585
R264 B.n312 B.n311 585
R265 B.n309 B.n252 585
R266 B.n308 B.n307 585
R267 B.n306 B.n305 585
R268 B.n304 B.n303 585
R269 B.n302 B.n301 585
R270 B.n300 B.n299 585
R271 B.n298 B.n297 585
R272 B.n295 B.n294 585
R273 B.n293 B.n292 585
R274 B.n291 B.n290 585
R275 B.n289 B.n288 585
R276 B.n287 B.n286 585
R277 B.n285 B.n284 585
R278 B.n283 B.n282 585
R279 B.n281 B.n280 585
R280 B.n279 B.n278 585
R281 B.n277 B.n276 585
R282 B.n275 B.n274 585
R283 B.n273 B.n272 585
R284 B.n271 B.n270 585
R285 B.n269 B.n268 585
R286 B.n267 B.n266 585
R287 B.n265 B.n264 585
R288 B.n263 B.n262 585
R289 B.n261 B.n260 585
R290 B.n259 B.n258 585
R291 B.n316 B.n236 585
R292 B.n236 B.n235 585
R293 B.n318 B.n317 585
R294 B.n319 B.n318 585
R295 B.n230 B.n229 585
R296 B.n231 B.n230 585
R297 B.n327 B.n326 585
R298 B.n326 B.n325 585
R299 B.n328 B.n228 585
R300 B.n228 B.n227 585
R301 B.n330 B.n329 585
R302 B.n331 B.n330 585
R303 B.n222 B.n221 585
R304 B.n223 B.n222 585
R305 B.n339 B.n338 585
R306 B.n338 B.n337 585
R307 B.n340 B.n220 585
R308 B.n220 B.n219 585
R309 B.n342 B.n341 585
R310 B.n343 B.n342 585
R311 B.n214 B.n213 585
R312 B.n215 B.n214 585
R313 B.n351 B.n350 585
R314 B.n350 B.n349 585
R315 B.n352 B.n212 585
R316 B.n212 B.n211 585
R317 B.n354 B.n353 585
R318 B.n355 B.n354 585
R319 B.n206 B.n205 585
R320 B.n207 B.n206 585
R321 B.n363 B.n362 585
R322 B.n362 B.n361 585
R323 B.n364 B.n204 585
R324 B.n204 B.n203 585
R325 B.n366 B.n365 585
R326 B.n367 B.n366 585
R327 B.n198 B.n197 585
R328 B.n199 B.n198 585
R329 B.n375 B.n374 585
R330 B.n374 B.n373 585
R331 B.n376 B.n196 585
R332 B.n196 B.n195 585
R333 B.n378 B.n377 585
R334 B.n379 B.n378 585
R335 B.n190 B.n189 585
R336 B.n191 B.n190 585
R337 B.n388 B.n387 585
R338 B.n387 B.n386 585
R339 B.n389 B.n188 585
R340 B.n385 B.n188 585
R341 B.n391 B.n390 585
R342 B.n392 B.n391 585
R343 B.n183 B.n182 585
R344 B.n184 B.n183 585
R345 B.n400 B.n399 585
R346 B.n399 B.n398 585
R347 B.n401 B.n181 585
R348 B.n181 B.n180 585
R349 B.n403 B.n402 585
R350 B.n404 B.n403 585
R351 B.n175 B.n174 585
R352 B.n176 B.n175 585
R353 B.n412 B.n411 585
R354 B.n411 B.n410 585
R355 B.n413 B.n173 585
R356 B.n173 B.n172 585
R357 B.n415 B.n414 585
R358 B.n416 B.n415 585
R359 B.n167 B.n166 585
R360 B.n168 B.n167 585
R361 B.n424 B.n423 585
R362 B.n423 B.n422 585
R363 B.n425 B.n165 585
R364 B.n165 B.n164 585
R365 B.n427 B.n426 585
R366 B.n428 B.n427 585
R367 B.n159 B.n158 585
R368 B.n160 B.n159 585
R369 B.n437 B.n436 585
R370 B.n436 B.n435 585
R371 B.n438 B.n157 585
R372 B.n157 B.n156 585
R373 B.n440 B.n439 585
R374 B.n441 B.n440 585
R375 B.n2 B.n0 585
R376 B.n4 B.n2 585
R377 B.n3 B.n1 585
R378 B.n589 B.n3 585
R379 B.n587 B.n586 585
R380 B.n588 B.n587 585
R381 B.n585 B.n9 585
R382 B.n9 B.n8 585
R383 B.n584 B.n583 585
R384 B.n583 B.n582 585
R385 B.n11 B.n10 585
R386 B.n581 B.n11 585
R387 B.n579 B.n578 585
R388 B.n580 B.n579 585
R389 B.n577 B.n16 585
R390 B.n16 B.n15 585
R391 B.n576 B.n575 585
R392 B.n575 B.n574 585
R393 B.n18 B.n17 585
R394 B.n573 B.n18 585
R395 B.n571 B.n570 585
R396 B.n572 B.n571 585
R397 B.n569 B.n23 585
R398 B.n23 B.n22 585
R399 B.n568 B.n567 585
R400 B.n567 B.n566 585
R401 B.n25 B.n24 585
R402 B.n565 B.n25 585
R403 B.n563 B.n562 585
R404 B.n564 B.n563 585
R405 B.n561 B.n30 585
R406 B.n30 B.n29 585
R407 B.n560 B.n559 585
R408 B.n559 B.n558 585
R409 B.n32 B.n31 585
R410 B.n557 B.n32 585
R411 B.n555 B.n554 585
R412 B.n556 B.n555 585
R413 B.n553 B.n36 585
R414 B.n39 B.n36 585
R415 B.n552 B.n551 585
R416 B.n551 B.n550 585
R417 B.n38 B.n37 585
R418 B.n549 B.n38 585
R419 B.n547 B.n546 585
R420 B.n548 B.n547 585
R421 B.n545 B.n44 585
R422 B.n44 B.n43 585
R423 B.n544 B.n543 585
R424 B.n543 B.n542 585
R425 B.n46 B.n45 585
R426 B.n541 B.n46 585
R427 B.n539 B.n538 585
R428 B.n540 B.n539 585
R429 B.n537 B.n51 585
R430 B.n51 B.n50 585
R431 B.n536 B.n535 585
R432 B.n535 B.n534 585
R433 B.n53 B.n52 585
R434 B.n533 B.n53 585
R435 B.n531 B.n530 585
R436 B.n532 B.n531 585
R437 B.n529 B.n58 585
R438 B.n58 B.n57 585
R439 B.n528 B.n527 585
R440 B.n527 B.n526 585
R441 B.n60 B.n59 585
R442 B.n525 B.n60 585
R443 B.n523 B.n522 585
R444 B.n524 B.n523 585
R445 B.n521 B.n65 585
R446 B.n65 B.n64 585
R447 B.n520 B.n519 585
R448 B.n519 B.n518 585
R449 B.n67 B.n66 585
R450 B.n517 B.n67 585
R451 B.n515 B.n514 585
R452 B.n516 B.n515 585
R453 B.n513 B.n72 585
R454 B.n72 B.n71 585
R455 B.n512 B.n511 585
R456 B.n511 B.n510 585
R457 B.n74 B.n73 585
R458 B.n509 B.n74 585
R459 B.n507 B.n506 585
R460 B.n508 B.n507 585
R461 B.n505 B.n79 585
R462 B.n79 B.n78 585
R463 B.n592 B.n591 585
R464 B.n591 B.n590 585
R465 B.n314 B.n236 439.647
R466 B.n503 B.n79 439.647
R467 B.n258 B.n234 439.647
R468 B.n500 B.n96 439.647
R469 B.n501 B.n94 256.663
R470 B.n501 B.n93 256.663
R471 B.n501 B.n92 256.663
R472 B.n501 B.n91 256.663
R473 B.n501 B.n90 256.663
R474 B.n501 B.n89 256.663
R475 B.n501 B.n88 256.663
R476 B.n501 B.n87 256.663
R477 B.n501 B.n86 256.663
R478 B.n501 B.n85 256.663
R479 B.n501 B.n84 256.663
R480 B.n501 B.n83 256.663
R481 B.n501 B.n82 256.663
R482 B.n502 B.n501 256.663
R483 B.n313 B.n312 256.663
R484 B.n312 B.n239 256.663
R485 B.n312 B.n240 256.663
R486 B.n312 B.n241 256.663
R487 B.n312 B.n242 256.663
R488 B.n312 B.n243 256.663
R489 B.n312 B.n244 256.663
R490 B.n312 B.n245 256.663
R491 B.n312 B.n246 256.663
R492 B.n312 B.n247 256.663
R493 B.n312 B.n248 256.663
R494 B.n312 B.n249 256.663
R495 B.n312 B.n250 256.663
R496 B.n312 B.n251 256.663
R497 B.n253 B.t14 222.518
R498 B.n99 B.t16 222.518
R499 B.n255 B.t11 222.518
R500 B.n97 B.t6 222.518
R501 B.n255 B.t8 209.804
R502 B.n253 B.t12 209.804
R503 B.n99 B.t15 209.804
R504 B.n97 B.t4 209.804
R505 B.n312 B.n235 188.078
R506 B.n501 B.n78 188.078
R507 B.n318 B.n236 163.367
R508 B.n318 B.n230 163.367
R509 B.n326 B.n230 163.367
R510 B.n326 B.n228 163.367
R511 B.n330 B.n228 163.367
R512 B.n330 B.n222 163.367
R513 B.n338 B.n222 163.367
R514 B.n338 B.n220 163.367
R515 B.n342 B.n220 163.367
R516 B.n342 B.n214 163.367
R517 B.n350 B.n214 163.367
R518 B.n350 B.n212 163.367
R519 B.n354 B.n212 163.367
R520 B.n354 B.n206 163.367
R521 B.n362 B.n206 163.367
R522 B.n362 B.n204 163.367
R523 B.n366 B.n204 163.367
R524 B.n366 B.n198 163.367
R525 B.n374 B.n198 163.367
R526 B.n374 B.n196 163.367
R527 B.n378 B.n196 163.367
R528 B.n378 B.n190 163.367
R529 B.n387 B.n190 163.367
R530 B.n387 B.n188 163.367
R531 B.n391 B.n188 163.367
R532 B.n391 B.n183 163.367
R533 B.n399 B.n183 163.367
R534 B.n399 B.n181 163.367
R535 B.n403 B.n181 163.367
R536 B.n403 B.n175 163.367
R537 B.n411 B.n175 163.367
R538 B.n411 B.n173 163.367
R539 B.n415 B.n173 163.367
R540 B.n415 B.n167 163.367
R541 B.n423 B.n167 163.367
R542 B.n423 B.n165 163.367
R543 B.n427 B.n165 163.367
R544 B.n427 B.n159 163.367
R545 B.n436 B.n159 163.367
R546 B.n436 B.n157 163.367
R547 B.n440 B.n157 163.367
R548 B.n440 B.n2 163.367
R549 B.n591 B.n2 163.367
R550 B.n591 B.n3 163.367
R551 B.n587 B.n3 163.367
R552 B.n587 B.n9 163.367
R553 B.n583 B.n9 163.367
R554 B.n583 B.n11 163.367
R555 B.n579 B.n11 163.367
R556 B.n579 B.n16 163.367
R557 B.n575 B.n16 163.367
R558 B.n575 B.n18 163.367
R559 B.n571 B.n18 163.367
R560 B.n571 B.n23 163.367
R561 B.n567 B.n23 163.367
R562 B.n567 B.n25 163.367
R563 B.n563 B.n25 163.367
R564 B.n563 B.n30 163.367
R565 B.n559 B.n30 163.367
R566 B.n559 B.n32 163.367
R567 B.n555 B.n32 163.367
R568 B.n555 B.n36 163.367
R569 B.n551 B.n36 163.367
R570 B.n551 B.n38 163.367
R571 B.n547 B.n38 163.367
R572 B.n547 B.n44 163.367
R573 B.n543 B.n44 163.367
R574 B.n543 B.n46 163.367
R575 B.n539 B.n46 163.367
R576 B.n539 B.n51 163.367
R577 B.n535 B.n51 163.367
R578 B.n535 B.n53 163.367
R579 B.n531 B.n53 163.367
R580 B.n531 B.n58 163.367
R581 B.n527 B.n58 163.367
R582 B.n527 B.n60 163.367
R583 B.n523 B.n60 163.367
R584 B.n523 B.n65 163.367
R585 B.n519 B.n65 163.367
R586 B.n519 B.n67 163.367
R587 B.n515 B.n67 163.367
R588 B.n515 B.n72 163.367
R589 B.n511 B.n72 163.367
R590 B.n511 B.n74 163.367
R591 B.n507 B.n74 163.367
R592 B.n507 B.n79 163.367
R593 B.n311 B.n238 163.367
R594 B.n311 B.n252 163.367
R595 B.n307 B.n306 163.367
R596 B.n303 B.n302 163.367
R597 B.n299 B.n298 163.367
R598 B.n294 B.n293 163.367
R599 B.n290 B.n289 163.367
R600 B.n286 B.n285 163.367
R601 B.n282 B.n281 163.367
R602 B.n278 B.n277 163.367
R603 B.n274 B.n273 163.367
R604 B.n270 B.n269 163.367
R605 B.n266 B.n265 163.367
R606 B.n262 B.n261 163.367
R607 B.n320 B.n234 163.367
R608 B.n320 B.n232 163.367
R609 B.n324 B.n232 163.367
R610 B.n324 B.n226 163.367
R611 B.n332 B.n226 163.367
R612 B.n332 B.n224 163.367
R613 B.n336 B.n224 163.367
R614 B.n336 B.n218 163.367
R615 B.n344 B.n218 163.367
R616 B.n344 B.n216 163.367
R617 B.n348 B.n216 163.367
R618 B.n348 B.n210 163.367
R619 B.n356 B.n210 163.367
R620 B.n356 B.n208 163.367
R621 B.n360 B.n208 163.367
R622 B.n360 B.n202 163.367
R623 B.n368 B.n202 163.367
R624 B.n368 B.n200 163.367
R625 B.n372 B.n200 163.367
R626 B.n372 B.n194 163.367
R627 B.n380 B.n194 163.367
R628 B.n380 B.n192 163.367
R629 B.n384 B.n192 163.367
R630 B.n384 B.n187 163.367
R631 B.n393 B.n187 163.367
R632 B.n393 B.n185 163.367
R633 B.n397 B.n185 163.367
R634 B.n397 B.n179 163.367
R635 B.n405 B.n179 163.367
R636 B.n405 B.n177 163.367
R637 B.n409 B.n177 163.367
R638 B.n409 B.n171 163.367
R639 B.n417 B.n171 163.367
R640 B.n417 B.n169 163.367
R641 B.n421 B.n169 163.367
R642 B.n421 B.n163 163.367
R643 B.n429 B.n163 163.367
R644 B.n429 B.n161 163.367
R645 B.n434 B.n161 163.367
R646 B.n434 B.n155 163.367
R647 B.n442 B.n155 163.367
R648 B.n443 B.n442 163.367
R649 B.n443 B.n5 163.367
R650 B.n6 B.n5 163.367
R651 B.n7 B.n6 163.367
R652 B.n448 B.n7 163.367
R653 B.n448 B.n12 163.367
R654 B.n13 B.n12 163.367
R655 B.n14 B.n13 163.367
R656 B.n453 B.n14 163.367
R657 B.n453 B.n19 163.367
R658 B.n20 B.n19 163.367
R659 B.n21 B.n20 163.367
R660 B.n458 B.n21 163.367
R661 B.n458 B.n26 163.367
R662 B.n27 B.n26 163.367
R663 B.n28 B.n27 163.367
R664 B.n463 B.n28 163.367
R665 B.n463 B.n33 163.367
R666 B.n34 B.n33 163.367
R667 B.n35 B.n34 163.367
R668 B.n468 B.n35 163.367
R669 B.n468 B.n40 163.367
R670 B.n41 B.n40 163.367
R671 B.n42 B.n41 163.367
R672 B.n473 B.n42 163.367
R673 B.n473 B.n47 163.367
R674 B.n48 B.n47 163.367
R675 B.n49 B.n48 163.367
R676 B.n478 B.n49 163.367
R677 B.n478 B.n54 163.367
R678 B.n55 B.n54 163.367
R679 B.n56 B.n55 163.367
R680 B.n483 B.n56 163.367
R681 B.n483 B.n61 163.367
R682 B.n62 B.n61 163.367
R683 B.n63 B.n62 163.367
R684 B.n488 B.n63 163.367
R685 B.n488 B.n68 163.367
R686 B.n69 B.n68 163.367
R687 B.n70 B.n69 163.367
R688 B.n493 B.n70 163.367
R689 B.n493 B.n75 163.367
R690 B.n76 B.n75 163.367
R691 B.n77 B.n76 163.367
R692 B.n96 B.n77 163.367
R693 B.n102 B.n81 163.367
R694 B.n106 B.n105 163.367
R695 B.n110 B.n109 163.367
R696 B.n114 B.n113 163.367
R697 B.n118 B.n117 163.367
R698 B.n122 B.n121 163.367
R699 B.n126 B.n125 163.367
R700 B.n130 B.n129 163.367
R701 B.n134 B.n133 163.367
R702 B.n139 B.n138 163.367
R703 B.n143 B.n142 163.367
R704 B.n147 B.n146 163.367
R705 B.n151 B.n150 163.367
R706 B.n500 B.n95 163.367
R707 B.n256 B.t10 146.299
R708 B.n254 B.t13 146.299
R709 B.n100 B.t17 146.299
R710 B.n98 B.t7 146.299
R711 B.n319 B.n235 117.334
R712 B.n319 B.n231 117.334
R713 B.n325 B.n231 117.334
R714 B.n325 B.n227 117.334
R715 B.n331 B.n227 117.334
R716 B.n331 B.n223 117.334
R717 B.n337 B.n223 117.334
R718 B.n337 B.n219 117.334
R719 B.n343 B.n219 117.334
R720 B.n349 B.n215 117.334
R721 B.n349 B.n211 117.334
R722 B.n355 B.n211 117.334
R723 B.n355 B.n207 117.334
R724 B.n361 B.n207 117.334
R725 B.n361 B.n203 117.334
R726 B.n367 B.n203 117.334
R727 B.n367 B.n199 117.334
R728 B.n373 B.n199 117.334
R729 B.n373 B.n195 117.334
R730 B.n379 B.n195 117.334
R731 B.n379 B.n191 117.334
R732 B.n386 B.n191 117.334
R733 B.n386 B.n385 117.334
R734 B.n392 B.n184 117.334
R735 B.n398 B.n184 117.334
R736 B.n398 B.n180 117.334
R737 B.n404 B.n180 117.334
R738 B.n404 B.n176 117.334
R739 B.n410 B.n176 117.334
R740 B.n410 B.n172 117.334
R741 B.n416 B.n172 117.334
R742 B.n416 B.n168 117.334
R743 B.n422 B.n168 117.334
R744 B.n428 B.n164 117.334
R745 B.n428 B.n160 117.334
R746 B.n435 B.n160 117.334
R747 B.n435 B.n156 117.334
R748 B.n441 B.n156 117.334
R749 B.n441 B.n4 117.334
R750 B.n590 B.n4 117.334
R751 B.n590 B.n589 117.334
R752 B.n589 B.n588 117.334
R753 B.n588 B.n8 117.334
R754 B.n582 B.n8 117.334
R755 B.n582 B.n581 117.334
R756 B.n581 B.n580 117.334
R757 B.n580 B.n15 117.334
R758 B.n574 B.n573 117.334
R759 B.n573 B.n572 117.334
R760 B.n572 B.n22 117.334
R761 B.n566 B.n22 117.334
R762 B.n566 B.n565 117.334
R763 B.n565 B.n564 117.334
R764 B.n564 B.n29 117.334
R765 B.n558 B.n29 117.334
R766 B.n558 B.n557 117.334
R767 B.n557 B.n556 117.334
R768 B.n550 B.n39 117.334
R769 B.n550 B.n549 117.334
R770 B.n549 B.n548 117.334
R771 B.n548 B.n43 117.334
R772 B.n542 B.n43 117.334
R773 B.n542 B.n541 117.334
R774 B.n541 B.n540 117.334
R775 B.n540 B.n50 117.334
R776 B.n534 B.n50 117.334
R777 B.n534 B.n533 117.334
R778 B.n533 B.n532 117.334
R779 B.n532 B.n57 117.334
R780 B.n526 B.n57 117.334
R781 B.n526 B.n525 117.334
R782 B.n524 B.n64 117.334
R783 B.n518 B.n64 117.334
R784 B.n518 B.n517 117.334
R785 B.n517 B.n516 117.334
R786 B.n516 B.n71 117.334
R787 B.n510 B.n71 117.334
R788 B.n510 B.n509 117.334
R789 B.n509 B.n508 117.334
R790 B.n508 B.n78 117.334
R791 B.n392 B.t0 110.431
R792 B.n556 B.t3 110.431
R793 B.t9 B.n215 82.824
R794 B.n525 B.t5 82.824
R795 B.n256 B.n255 76.2187
R796 B.n254 B.n253 76.2187
R797 B.n100 B.n99 76.2187
R798 B.n98 B.n97 76.2187
R799 B.n422 B.t2 72.4711
R800 B.n574 B.t1 72.4711
R801 B.n314 B.n313 71.676
R802 B.n252 B.n239 71.676
R803 B.n306 B.n240 71.676
R804 B.n302 B.n241 71.676
R805 B.n298 B.n242 71.676
R806 B.n293 B.n243 71.676
R807 B.n289 B.n244 71.676
R808 B.n285 B.n245 71.676
R809 B.n281 B.n246 71.676
R810 B.n277 B.n247 71.676
R811 B.n273 B.n248 71.676
R812 B.n269 B.n249 71.676
R813 B.n265 B.n250 71.676
R814 B.n261 B.n251 71.676
R815 B.n503 B.n502 71.676
R816 B.n102 B.n82 71.676
R817 B.n106 B.n83 71.676
R818 B.n110 B.n84 71.676
R819 B.n114 B.n85 71.676
R820 B.n118 B.n86 71.676
R821 B.n122 B.n87 71.676
R822 B.n126 B.n88 71.676
R823 B.n130 B.n89 71.676
R824 B.n134 B.n90 71.676
R825 B.n139 B.n91 71.676
R826 B.n143 B.n92 71.676
R827 B.n147 B.n93 71.676
R828 B.n151 B.n94 71.676
R829 B.n95 B.n94 71.676
R830 B.n150 B.n93 71.676
R831 B.n146 B.n92 71.676
R832 B.n142 B.n91 71.676
R833 B.n138 B.n90 71.676
R834 B.n133 B.n89 71.676
R835 B.n129 B.n88 71.676
R836 B.n125 B.n87 71.676
R837 B.n121 B.n86 71.676
R838 B.n117 B.n85 71.676
R839 B.n113 B.n84 71.676
R840 B.n109 B.n83 71.676
R841 B.n105 B.n82 71.676
R842 B.n502 B.n81 71.676
R843 B.n313 B.n238 71.676
R844 B.n307 B.n239 71.676
R845 B.n303 B.n240 71.676
R846 B.n299 B.n241 71.676
R847 B.n294 B.n242 71.676
R848 B.n290 B.n243 71.676
R849 B.n286 B.n244 71.676
R850 B.n282 B.n245 71.676
R851 B.n278 B.n246 71.676
R852 B.n274 B.n247 71.676
R853 B.n270 B.n248 71.676
R854 B.n266 B.n249 71.676
R855 B.n262 B.n250 71.676
R856 B.n258 B.n251 71.676
R857 B.n257 B.n256 59.5399
R858 B.n296 B.n254 59.5399
R859 B.n101 B.n100 59.5399
R860 B.n136 B.n98 59.5399
R861 B.t2 B.n164 44.8632
R862 B.t1 B.n15 44.8632
R863 B.n343 B.t9 34.5103
R864 B.t5 B.n524 34.5103
R865 B.n505 B.n504 28.5664
R866 B.n259 B.n233 28.5664
R867 B.n316 B.n315 28.5664
R868 B.n499 B.n498 28.5664
R869 B B.n592 18.0485
R870 B.n504 B.n80 10.6151
R871 B.n103 B.n80 10.6151
R872 B.n104 B.n103 10.6151
R873 B.n107 B.n104 10.6151
R874 B.n108 B.n107 10.6151
R875 B.n111 B.n108 10.6151
R876 B.n112 B.n111 10.6151
R877 B.n115 B.n112 10.6151
R878 B.n116 B.n115 10.6151
R879 B.n120 B.n119 10.6151
R880 B.n123 B.n120 10.6151
R881 B.n124 B.n123 10.6151
R882 B.n127 B.n124 10.6151
R883 B.n128 B.n127 10.6151
R884 B.n131 B.n128 10.6151
R885 B.n132 B.n131 10.6151
R886 B.n135 B.n132 10.6151
R887 B.n140 B.n137 10.6151
R888 B.n141 B.n140 10.6151
R889 B.n144 B.n141 10.6151
R890 B.n145 B.n144 10.6151
R891 B.n148 B.n145 10.6151
R892 B.n149 B.n148 10.6151
R893 B.n152 B.n149 10.6151
R894 B.n153 B.n152 10.6151
R895 B.n499 B.n153 10.6151
R896 B.n321 B.n233 10.6151
R897 B.n322 B.n321 10.6151
R898 B.n323 B.n322 10.6151
R899 B.n323 B.n225 10.6151
R900 B.n333 B.n225 10.6151
R901 B.n334 B.n333 10.6151
R902 B.n335 B.n334 10.6151
R903 B.n335 B.n217 10.6151
R904 B.n345 B.n217 10.6151
R905 B.n346 B.n345 10.6151
R906 B.n347 B.n346 10.6151
R907 B.n347 B.n209 10.6151
R908 B.n357 B.n209 10.6151
R909 B.n358 B.n357 10.6151
R910 B.n359 B.n358 10.6151
R911 B.n359 B.n201 10.6151
R912 B.n369 B.n201 10.6151
R913 B.n370 B.n369 10.6151
R914 B.n371 B.n370 10.6151
R915 B.n371 B.n193 10.6151
R916 B.n381 B.n193 10.6151
R917 B.n382 B.n381 10.6151
R918 B.n383 B.n382 10.6151
R919 B.n383 B.n186 10.6151
R920 B.n394 B.n186 10.6151
R921 B.n395 B.n394 10.6151
R922 B.n396 B.n395 10.6151
R923 B.n396 B.n178 10.6151
R924 B.n406 B.n178 10.6151
R925 B.n407 B.n406 10.6151
R926 B.n408 B.n407 10.6151
R927 B.n408 B.n170 10.6151
R928 B.n418 B.n170 10.6151
R929 B.n419 B.n418 10.6151
R930 B.n420 B.n419 10.6151
R931 B.n420 B.n162 10.6151
R932 B.n430 B.n162 10.6151
R933 B.n431 B.n430 10.6151
R934 B.n433 B.n431 10.6151
R935 B.n433 B.n432 10.6151
R936 B.n432 B.n154 10.6151
R937 B.n444 B.n154 10.6151
R938 B.n445 B.n444 10.6151
R939 B.n446 B.n445 10.6151
R940 B.n447 B.n446 10.6151
R941 B.n449 B.n447 10.6151
R942 B.n450 B.n449 10.6151
R943 B.n451 B.n450 10.6151
R944 B.n452 B.n451 10.6151
R945 B.n454 B.n452 10.6151
R946 B.n455 B.n454 10.6151
R947 B.n456 B.n455 10.6151
R948 B.n457 B.n456 10.6151
R949 B.n459 B.n457 10.6151
R950 B.n460 B.n459 10.6151
R951 B.n461 B.n460 10.6151
R952 B.n462 B.n461 10.6151
R953 B.n464 B.n462 10.6151
R954 B.n465 B.n464 10.6151
R955 B.n466 B.n465 10.6151
R956 B.n467 B.n466 10.6151
R957 B.n469 B.n467 10.6151
R958 B.n470 B.n469 10.6151
R959 B.n471 B.n470 10.6151
R960 B.n472 B.n471 10.6151
R961 B.n474 B.n472 10.6151
R962 B.n475 B.n474 10.6151
R963 B.n476 B.n475 10.6151
R964 B.n477 B.n476 10.6151
R965 B.n479 B.n477 10.6151
R966 B.n480 B.n479 10.6151
R967 B.n481 B.n480 10.6151
R968 B.n482 B.n481 10.6151
R969 B.n484 B.n482 10.6151
R970 B.n485 B.n484 10.6151
R971 B.n486 B.n485 10.6151
R972 B.n487 B.n486 10.6151
R973 B.n489 B.n487 10.6151
R974 B.n490 B.n489 10.6151
R975 B.n491 B.n490 10.6151
R976 B.n492 B.n491 10.6151
R977 B.n494 B.n492 10.6151
R978 B.n495 B.n494 10.6151
R979 B.n496 B.n495 10.6151
R980 B.n497 B.n496 10.6151
R981 B.n498 B.n497 10.6151
R982 B.n315 B.n237 10.6151
R983 B.n310 B.n237 10.6151
R984 B.n310 B.n309 10.6151
R985 B.n309 B.n308 10.6151
R986 B.n308 B.n305 10.6151
R987 B.n305 B.n304 10.6151
R988 B.n304 B.n301 10.6151
R989 B.n301 B.n300 10.6151
R990 B.n300 B.n297 10.6151
R991 B.n295 B.n292 10.6151
R992 B.n292 B.n291 10.6151
R993 B.n291 B.n288 10.6151
R994 B.n288 B.n287 10.6151
R995 B.n287 B.n284 10.6151
R996 B.n284 B.n283 10.6151
R997 B.n283 B.n280 10.6151
R998 B.n280 B.n279 10.6151
R999 B.n276 B.n275 10.6151
R1000 B.n275 B.n272 10.6151
R1001 B.n272 B.n271 10.6151
R1002 B.n271 B.n268 10.6151
R1003 B.n268 B.n267 10.6151
R1004 B.n267 B.n264 10.6151
R1005 B.n264 B.n263 10.6151
R1006 B.n263 B.n260 10.6151
R1007 B.n260 B.n259 10.6151
R1008 B.n317 B.n316 10.6151
R1009 B.n317 B.n229 10.6151
R1010 B.n327 B.n229 10.6151
R1011 B.n328 B.n327 10.6151
R1012 B.n329 B.n328 10.6151
R1013 B.n329 B.n221 10.6151
R1014 B.n339 B.n221 10.6151
R1015 B.n340 B.n339 10.6151
R1016 B.n341 B.n340 10.6151
R1017 B.n341 B.n213 10.6151
R1018 B.n351 B.n213 10.6151
R1019 B.n352 B.n351 10.6151
R1020 B.n353 B.n352 10.6151
R1021 B.n353 B.n205 10.6151
R1022 B.n363 B.n205 10.6151
R1023 B.n364 B.n363 10.6151
R1024 B.n365 B.n364 10.6151
R1025 B.n365 B.n197 10.6151
R1026 B.n375 B.n197 10.6151
R1027 B.n376 B.n375 10.6151
R1028 B.n377 B.n376 10.6151
R1029 B.n377 B.n189 10.6151
R1030 B.n388 B.n189 10.6151
R1031 B.n389 B.n388 10.6151
R1032 B.n390 B.n389 10.6151
R1033 B.n390 B.n182 10.6151
R1034 B.n400 B.n182 10.6151
R1035 B.n401 B.n400 10.6151
R1036 B.n402 B.n401 10.6151
R1037 B.n402 B.n174 10.6151
R1038 B.n412 B.n174 10.6151
R1039 B.n413 B.n412 10.6151
R1040 B.n414 B.n413 10.6151
R1041 B.n414 B.n166 10.6151
R1042 B.n424 B.n166 10.6151
R1043 B.n425 B.n424 10.6151
R1044 B.n426 B.n425 10.6151
R1045 B.n426 B.n158 10.6151
R1046 B.n437 B.n158 10.6151
R1047 B.n438 B.n437 10.6151
R1048 B.n439 B.n438 10.6151
R1049 B.n439 B.n0 10.6151
R1050 B.n586 B.n1 10.6151
R1051 B.n586 B.n585 10.6151
R1052 B.n585 B.n584 10.6151
R1053 B.n584 B.n10 10.6151
R1054 B.n578 B.n10 10.6151
R1055 B.n578 B.n577 10.6151
R1056 B.n577 B.n576 10.6151
R1057 B.n576 B.n17 10.6151
R1058 B.n570 B.n17 10.6151
R1059 B.n570 B.n569 10.6151
R1060 B.n569 B.n568 10.6151
R1061 B.n568 B.n24 10.6151
R1062 B.n562 B.n24 10.6151
R1063 B.n562 B.n561 10.6151
R1064 B.n561 B.n560 10.6151
R1065 B.n560 B.n31 10.6151
R1066 B.n554 B.n31 10.6151
R1067 B.n554 B.n553 10.6151
R1068 B.n553 B.n552 10.6151
R1069 B.n552 B.n37 10.6151
R1070 B.n546 B.n37 10.6151
R1071 B.n546 B.n545 10.6151
R1072 B.n545 B.n544 10.6151
R1073 B.n544 B.n45 10.6151
R1074 B.n538 B.n45 10.6151
R1075 B.n538 B.n537 10.6151
R1076 B.n537 B.n536 10.6151
R1077 B.n536 B.n52 10.6151
R1078 B.n530 B.n52 10.6151
R1079 B.n530 B.n529 10.6151
R1080 B.n529 B.n528 10.6151
R1081 B.n528 B.n59 10.6151
R1082 B.n522 B.n59 10.6151
R1083 B.n522 B.n521 10.6151
R1084 B.n521 B.n520 10.6151
R1085 B.n520 B.n66 10.6151
R1086 B.n514 B.n66 10.6151
R1087 B.n514 B.n513 10.6151
R1088 B.n513 B.n512 10.6151
R1089 B.n512 B.n73 10.6151
R1090 B.n506 B.n73 10.6151
R1091 B.n506 B.n505 10.6151
R1092 B.n385 B.t0 6.90246
R1093 B.n39 B.t3 6.90246
R1094 B.n119 B.n101 6.5566
R1095 B.n136 B.n135 6.5566
R1096 B.n296 B.n295 6.5566
R1097 B.n279 B.n257 6.5566
R1098 B.n116 B.n101 4.05904
R1099 B.n137 B.n136 4.05904
R1100 B.n297 B.n296 4.05904
R1101 B.n276 B.n257 4.05904
R1102 B.n592 B.n0 2.81026
R1103 B.n592 B.n1 2.81026
R1104 VN VN.n1 43.4892
R1105 VN.n1 VN.t1 42.1582
R1106 VN.n0 VN.t0 42.1582
R1107 VN.n0 VN.t2 40.9152
R1108 VN.n1 VN.t3 40.9152
R1109 VN VN.n0 2.10662
R1110 VDD2.n2 VDD2.n0 181.065
R1111 VDD2.n2 VDD2.n1 146.238
R1112 VDD2.n1 VDD2.t0 18.0005
R1113 VDD2.n1 VDD2.t2 18.0005
R1114 VDD2.n0 VDD2.t3 18.0005
R1115 VDD2.n0 VDD2.t1 18.0005
R1116 VDD2 VDD2.n2 0.0586897
C0 VN VTAIL 1.69702f
C1 VDD1 VTAIL 3.36628f
C2 VDD1 VN 0.156575f
C3 VDD2 VP 0.466122f
C4 VP VTAIL 1.71112f
C5 VP VN 4.9055f
C6 VP VDD1 1.07116f
C7 VDD2 VTAIL 3.42719f
C8 VDD2 VN 0.76442f
C9 VDD2 VDD1 1.26814f
C10 VDD2 B 3.456769f
C11 VDD1 B 6.42067f
C12 VTAIL B 3.424703f
C13 VN B 11.49025f
C14 VP B 10.022605f
C15 VDD2.t3 B 0.021818f
C16 VDD2.t1 B 0.021818f
C17 VDD2.n0 B 0.286882f
C18 VDD2.t0 B 0.021818f
C19 VDD2.t2 B 0.021818f
C20 VDD2.n1 B 0.111782f
C21 VDD2.n2 B 2.63466f
C22 VN.t2 B 0.416341f
C23 VN.t0 B 0.426471f
C24 VN.n0 B 0.338072f
C25 VN.t1 B 0.426471f
C26 VN.t3 B 0.416341f
C27 VN.n1 B 1.53606f
C28 VDD1.t0 B 0.021239f
C29 VDD1.t3 B 0.021239f
C30 VDD1.n0 B 0.108988f
C31 VDD1.t1 B 0.021239f
C32 VDD1.t2 B 0.021239f
C33 VDD1.n1 B 0.290898f
C34 VTAIL.t1 B 0.11683f
C35 VTAIL.n0 B 0.316092f
C36 VTAIL.t7 B 0.11683f
C37 VTAIL.n1 B 0.436273f
C38 VTAIL.t6 B 0.11683f
C39 VTAIL.n2 B 1.03007f
C40 VTAIL.t0 B 0.11683f
C41 VTAIL.n3 B 1.03007f
C42 VTAIL.t2 B 0.11683f
C43 VTAIL.n4 B 0.436273f
C44 VTAIL.t5 B 0.11683f
C45 VTAIL.n5 B 0.436273f
C46 VTAIL.t4 B 0.11683f
C47 VTAIL.n6 B 1.03007f
C48 VTAIL.t3 B 0.11683f
C49 VTAIL.n7 B 0.901334f
C50 VP.t1 B 0.18269f
C51 VP.n0 B 0.204143f
C52 VP.n1 B 0.023619f
C53 VP.n2 B 0.03463f
C54 VP.n3 B 0.023619f
C55 VP.n4 B 0.03179f
C56 VP.t3 B 0.42936f
C57 VP.t0 B 0.419162f
C58 VP.n5 B 1.53636f
C59 VP.t2 B 0.18269f
C60 VP.n6 B 0.204143f
C61 VP.n7 B 1.09806f
C62 VP.n8 B 0.038127f
C63 VP.n9 B 0.023619f
C64 VP.n10 B 0.044241f
C65 VP.n11 B 0.044241f
C66 VP.n12 B 0.03463f
C67 VP.n13 B 0.023619f
C68 VP.n14 B 0.023619f
C69 VP.n15 B 0.023619f
C70 VP.n16 B 0.044241f
C71 VP.n17 B 0.044241f
C72 VP.n18 B 0.03179f
C73 VP.n19 B 0.038127f
C74 VP.n20 B 0.064172f
.ends

