* NGSPICE file created from diff_pair_sample_1147.ext - technology: sky130A

.subckt diff_pair_sample_1147 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VP.t0 VDD1.t1 w_n2030_n4702# sky130_fd_pr__pfet_01v8 ad=7.2813 pd=38.12 as=3.08055 ps=19 w=18.67 l=0.73
X1 VTAIL.t14 VP.t1 VDD1.t0 w_n2030_n4702# sky130_fd_pr__pfet_01v8 ad=7.2813 pd=38.12 as=3.08055 ps=19 w=18.67 l=0.73
X2 VDD1.t3 VP.t2 VTAIL.t13 w_n2030_n4702# sky130_fd_pr__pfet_01v8 ad=3.08055 pd=19 as=3.08055 ps=19 w=18.67 l=0.73
X3 VTAIL.t12 VP.t3 VDD1.t2 w_n2030_n4702# sky130_fd_pr__pfet_01v8 ad=3.08055 pd=19 as=3.08055 ps=19 w=18.67 l=0.73
X4 B.t11 B.t9 B.t10 w_n2030_n4702# sky130_fd_pr__pfet_01v8 ad=7.2813 pd=38.12 as=0 ps=0 w=18.67 l=0.73
X5 VDD1.t7 VP.t4 VTAIL.t11 w_n2030_n4702# sky130_fd_pr__pfet_01v8 ad=3.08055 pd=19 as=7.2813 ps=38.12 w=18.67 l=0.73
X6 VTAIL.t10 VP.t5 VDD1.t6 w_n2030_n4702# sky130_fd_pr__pfet_01v8 ad=3.08055 pd=19 as=3.08055 ps=19 w=18.67 l=0.73
X7 B.t8 B.t6 B.t7 w_n2030_n4702# sky130_fd_pr__pfet_01v8 ad=7.2813 pd=38.12 as=0 ps=0 w=18.67 l=0.73
X8 VDD2.t7 VN.t0 VTAIL.t2 w_n2030_n4702# sky130_fd_pr__pfet_01v8 ad=3.08055 pd=19 as=7.2813 ps=38.12 w=18.67 l=0.73
X9 VDD2.t6 VN.t1 VTAIL.t7 w_n2030_n4702# sky130_fd_pr__pfet_01v8 ad=3.08055 pd=19 as=3.08055 ps=19 w=18.67 l=0.73
X10 VDD1.t5 VP.t6 VTAIL.t9 w_n2030_n4702# sky130_fd_pr__pfet_01v8 ad=3.08055 pd=19 as=3.08055 ps=19 w=18.67 l=0.73
X11 B.t5 B.t3 B.t4 w_n2030_n4702# sky130_fd_pr__pfet_01v8 ad=7.2813 pd=38.12 as=0 ps=0 w=18.67 l=0.73
X12 VDD2.t5 VN.t2 VTAIL.t6 w_n2030_n4702# sky130_fd_pr__pfet_01v8 ad=3.08055 pd=19 as=3.08055 ps=19 w=18.67 l=0.73
X13 VDD2.t4 VN.t3 VTAIL.t5 w_n2030_n4702# sky130_fd_pr__pfet_01v8 ad=3.08055 pd=19 as=7.2813 ps=38.12 w=18.67 l=0.73
X14 VTAIL.t3 VN.t4 VDD2.t3 w_n2030_n4702# sky130_fd_pr__pfet_01v8 ad=7.2813 pd=38.12 as=3.08055 ps=19 w=18.67 l=0.73
X15 VTAIL.t4 VN.t5 VDD2.t2 w_n2030_n4702# sky130_fd_pr__pfet_01v8 ad=3.08055 pd=19 as=3.08055 ps=19 w=18.67 l=0.73
X16 B.t2 B.t0 B.t1 w_n2030_n4702# sky130_fd_pr__pfet_01v8 ad=7.2813 pd=38.12 as=0 ps=0 w=18.67 l=0.73
X17 VDD1.t4 VP.t7 VTAIL.t8 w_n2030_n4702# sky130_fd_pr__pfet_01v8 ad=3.08055 pd=19 as=7.2813 ps=38.12 w=18.67 l=0.73
X18 VTAIL.t1 VN.t6 VDD2.t1 w_n2030_n4702# sky130_fd_pr__pfet_01v8 ad=3.08055 pd=19 as=3.08055 ps=19 w=18.67 l=0.73
X19 VTAIL.t0 VN.t7 VDD2.t0 w_n2030_n4702# sky130_fd_pr__pfet_01v8 ad=7.2813 pd=38.12 as=3.08055 ps=19 w=18.67 l=0.73
R0 VP.n6 VP.t0 693.812
R1 VP.n14 VP.t1 670.509
R2 VP.n16 VP.t2 670.509
R3 VP.n20 VP.t3 670.509
R4 VP.n22 VP.t4 670.509
R5 VP.n11 VP.t7 670.509
R6 VP.n9 VP.t5 670.509
R7 VP.n5 VP.t6 670.509
R8 VP.n23 VP.n22 161.3
R9 VP.n8 VP.n7 161.3
R10 VP.n9 VP.n4 161.3
R11 VP.n10 VP.n3 161.3
R12 VP.n12 VP.n11 161.3
R13 VP.n21 VP.n0 161.3
R14 VP.n20 VP.n19 161.3
R15 VP.n18 VP.n1 161.3
R16 VP.n17 VP.n16 161.3
R17 VP.n15 VP.n2 161.3
R18 VP.n14 VP.n13 161.3
R19 VP.n13 VP.n12 47.2278
R20 VP.n7 VP.n6 44.8907
R21 VP.n15 VP.n14 32.8641
R22 VP.n22 VP.n21 32.8641
R23 VP.n11 VP.n10 32.8641
R24 VP.n16 VP.n1 24.1005
R25 VP.n20 VP.n1 24.1005
R26 VP.n8 VP.n5 24.1005
R27 VP.n9 VP.n8 24.1005
R28 VP.n6 VP.n5 18.4104
R29 VP.n16 VP.n15 15.3369
R30 VP.n21 VP.n20 15.3369
R31 VP.n10 VP.n9 15.3369
R32 VP.n7 VP.n4 0.189894
R33 VP.n4 VP.n3 0.189894
R34 VP.n12 VP.n3 0.189894
R35 VP.n13 VP.n2 0.189894
R36 VP.n17 VP.n2 0.189894
R37 VP.n18 VP.n17 0.189894
R38 VP.n19 VP.n18 0.189894
R39 VP.n19 VP.n0 0.189894
R40 VP.n23 VP.n0 0.189894
R41 VP VP.n23 0.0516364
R42 VDD1 VDD1.n0 70.4052
R43 VDD1.n3 VDD1.n2 70.2914
R44 VDD1.n3 VDD1.n1 70.2914
R45 VDD1.n5 VDD1.n4 69.8899
R46 VDD1.n5 VDD1.n3 44.5052
R47 VDD1.n4 VDD1.t6 1.74153
R48 VDD1.n4 VDD1.t4 1.74153
R49 VDD1.n0 VDD1.t1 1.74153
R50 VDD1.n0 VDD1.t5 1.74153
R51 VDD1.n2 VDD1.t2 1.74153
R52 VDD1.n2 VDD1.t7 1.74153
R53 VDD1.n1 VDD1.t0 1.74153
R54 VDD1.n1 VDD1.t3 1.74153
R55 VDD1 VDD1.n5 0.399207
R56 VTAIL.n11 VTAIL.t15 54.9523
R57 VTAIL.n10 VTAIL.t2 54.9523
R58 VTAIL.n7 VTAIL.t0 54.9523
R59 VTAIL.n14 VTAIL.t8 54.9522
R60 VTAIL.n15 VTAIL.t5 54.9521
R61 VTAIL.n2 VTAIL.t3 54.9521
R62 VTAIL.n3 VTAIL.t11 54.9521
R63 VTAIL.n6 VTAIL.t14 54.9521
R64 VTAIL.n13 VTAIL.n12 53.2113
R65 VTAIL.n9 VTAIL.n8 53.2113
R66 VTAIL.n1 VTAIL.n0 53.2111
R67 VTAIL.n5 VTAIL.n4 53.2111
R68 VTAIL.n15 VTAIL.n14 29.3755
R69 VTAIL.n7 VTAIL.n6 29.3755
R70 VTAIL.n0 VTAIL.t6 1.74153
R71 VTAIL.n0 VTAIL.t4 1.74153
R72 VTAIL.n4 VTAIL.t13 1.74153
R73 VTAIL.n4 VTAIL.t12 1.74153
R74 VTAIL.n12 VTAIL.t9 1.74153
R75 VTAIL.n12 VTAIL.t10 1.74153
R76 VTAIL.n8 VTAIL.t7 1.74153
R77 VTAIL.n8 VTAIL.t1 1.74153
R78 VTAIL.n9 VTAIL.n7 0.914293
R79 VTAIL.n10 VTAIL.n9 0.914293
R80 VTAIL.n13 VTAIL.n11 0.914293
R81 VTAIL.n14 VTAIL.n13 0.914293
R82 VTAIL.n6 VTAIL.n5 0.914293
R83 VTAIL.n5 VTAIL.n3 0.914293
R84 VTAIL.n2 VTAIL.n1 0.914293
R85 VTAIL VTAIL.n15 0.856103
R86 VTAIL.n11 VTAIL.n10 0.470328
R87 VTAIL.n3 VTAIL.n2 0.470328
R88 VTAIL VTAIL.n1 0.0586897
R89 B.n144 B.t0 818.977
R90 B.n326 B.t3 818.977
R91 B.n52 B.t9 818.977
R92 B.n44 B.t6 818.977
R93 B.n421 B.n108 585
R94 B.n420 B.n419 585
R95 B.n418 B.n109 585
R96 B.n417 B.n416 585
R97 B.n415 B.n110 585
R98 B.n414 B.n413 585
R99 B.n412 B.n111 585
R100 B.n411 B.n410 585
R101 B.n409 B.n112 585
R102 B.n408 B.n407 585
R103 B.n406 B.n113 585
R104 B.n405 B.n404 585
R105 B.n403 B.n114 585
R106 B.n402 B.n401 585
R107 B.n400 B.n115 585
R108 B.n399 B.n398 585
R109 B.n397 B.n116 585
R110 B.n396 B.n395 585
R111 B.n394 B.n117 585
R112 B.n393 B.n392 585
R113 B.n391 B.n118 585
R114 B.n390 B.n389 585
R115 B.n388 B.n119 585
R116 B.n387 B.n386 585
R117 B.n385 B.n120 585
R118 B.n384 B.n383 585
R119 B.n382 B.n121 585
R120 B.n381 B.n380 585
R121 B.n379 B.n122 585
R122 B.n378 B.n377 585
R123 B.n376 B.n123 585
R124 B.n375 B.n374 585
R125 B.n373 B.n124 585
R126 B.n372 B.n371 585
R127 B.n370 B.n125 585
R128 B.n369 B.n368 585
R129 B.n367 B.n126 585
R130 B.n366 B.n365 585
R131 B.n364 B.n127 585
R132 B.n363 B.n362 585
R133 B.n361 B.n128 585
R134 B.n360 B.n359 585
R135 B.n358 B.n129 585
R136 B.n357 B.n356 585
R137 B.n355 B.n130 585
R138 B.n354 B.n353 585
R139 B.n352 B.n131 585
R140 B.n351 B.n350 585
R141 B.n349 B.n132 585
R142 B.n348 B.n347 585
R143 B.n346 B.n133 585
R144 B.n345 B.n344 585
R145 B.n343 B.n134 585
R146 B.n342 B.n341 585
R147 B.n340 B.n135 585
R148 B.n339 B.n338 585
R149 B.n337 B.n136 585
R150 B.n336 B.n335 585
R151 B.n334 B.n137 585
R152 B.n333 B.n332 585
R153 B.n331 B.n138 585
R154 B.n330 B.n329 585
R155 B.n325 B.n139 585
R156 B.n324 B.n323 585
R157 B.n322 B.n140 585
R158 B.n321 B.n320 585
R159 B.n319 B.n141 585
R160 B.n318 B.n317 585
R161 B.n316 B.n142 585
R162 B.n315 B.n314 585
R163 B.n313 B.n143 585
R164 B.n311 B.n310 585
R165 B.n309 B.n146 585
R166 B.n308 B.n307 585
R167 B.n306 B.n147 585
R168 B.n305 B.n304 585
R169 B.n303 B.n148 585
R170 B.n302 B.n301 585
R171 B.n300 B.n149 585
R172 B.n299 B.n298 585
R173 B.n297 B.n150 585
R174 B.n296 B.n295 585
R175 B.n294 B.n151 585
R176 B.n293 B.n292 585
R177 B.n291 B.n152 585
R178 B.n290 B.n289 585
R179 B.n288 B.n153 585
R180 B.n287 B.n286 585
R181 B.n285 B.n154 585
R182 B.n284 B.n283 585
R183 B.n282 B.n155 585
R184 B.n281 B.n280 585
R185 B.n279 B.n156 585
R186 B.n278 B.n277 585
R187 B.n276 B.n157 585
R188 B.n275 B.n274 585
R189 B.n273 B.n158 585
R190 B.n272 B.n271 585
R191 B.n270 B.n159 585
R192 B.n269 B.n268 585
R193 B.n267 B.n160 585
R194 B.n266 B.n265 585
R195 B.n264 B.n161 585
R196 B.n263 B.n262 585
R197 B.n261 B.n162 585
R198 B.n260 B.n259 585
R199 B.n258 B.n163 585
R200 B.n257 B.n256 585
R201 B.n255 B.n164 585
R202 B.n254 B.n253 585
R203 B.n252 B.n165 585
R204 B.n251 B.n250 585
R205 B.n249 B.n166 585
R206 B.n248 B.n247 585
R207 B.n246 B.n167 585
R208 B.n245 B.n244 585
R209 B.n243 B.n168 585
R210 B.n242 B.n241 585
R211 B.n240 B.n169 585
R212 B.n239 B.n238 585
R213 B.n237 B.n170 585
R214 B.n236 B.n235 585
R215 B.n234 B.n171 585
R216 B.n233 B.n232 585
R217 B.n231 B.n172 585
R218 B.n230 B.n229 585
R219 B.n228 B.n173 585
R220 B.n227 B.n226 585
R221 B.n225 B.n174 585
R222 B.n224 B.n223 585
R223 B.n222 B.n175 585
R224 B.n221 B.n220 585
R225 B.n423 B.n422 585
R226 B.n424 B.n107 585
R227 B.n426 B.n425 585
R228 B.n427 B.n106 585
R229 B.n429 B.n428 585
R230 B.n430 B.n105 585
R231 B.n432 B.n431 585
R232 B.n433 B.n104 585
R233 B.n435 B.n434 585
R234 B.n436 B.n103 585
R235 B.n438 B.n437 585
R236 B.n439 B.n102 585
R237 B.n441 B.n440 585
R238 B.n442 B.n101 585
R239 B.n444 B.n443 585
R240 B.n445 B.n100 585
R241 B.n447 B.n446 585
R242 B.n448 B.n99 585
R243 B.n450 B.n449 585
R244 B.n451 B.n98 585
R245 B.n453 B.n452 585
R246 B.n454 B.n97 585
R247 B.n456 B.n455 585
R248 B.n457 B.n96 585
R249 B.n459 B.n458 585
R250 B.n460 B.n95 585
R251 B.n462 B.n461 585
R252 B.n463 B.n94 585
R253 B.n465 B.n464 585
R254 B.n466 B.n93 585
R255 B.n468 B.n467 585
R256 B.n469 B.n92 585
R257 B.n471 B.n470 585
R258 B.n472 B.n91 585
R259 B.n474 B.n473 585
R260 B.n475 B.n90 585
R261 B.n477 B.n476 585
R262 B.n478 B.n89 585
R263 B.n480 B.n479 585
R264 B.n481 B.n88 585
R265 B.n483 B.n482 585
R266 B.n484 B.n87 585
R267 B.n486 B.n485 585
R268 B.n487 B.n86 585
R269 B.n489 B.n488 585
R270 B.n490 B.n85 585
R271 B.n492 B.n491 585
R272 B.n493 B.n84 585
R273 B.n693 B.n692 585
R274 B.n691 B.n14 585
R275 B.n690 B.n689 585
R276 B.n688 B.n15 585
R277 B.n687 B.n686 585
R278 B.n685 B.n16 585
R279 B.n684 B.n683 585
R280 B.n682 B.n17 585
R281 B.n681 B.n680 585
R282 B.n679 B.n18 585
R283 B.n678 B.n677 585
R284 B.n676 B.n19 585
R285 B.n675 B.n674 585
R286 B.n673 B.n20 585
R287 B.n672 B.n671 585
R288 B.n670 B.n21 585
R289 B.n669 B.n668 585
R290 B.n667 B.n22 585
R291 B.n666 B.n665 585
R292 B.n664 B.n23 585
R293 B.n663 B.n662 585
R294 B.n661 B.n24 585
R295 B.n660 B.n659 585
R296 B.n658 B.n25 585
R297 B.n657 B.n656 585
R298 B.n655 B.n26 585
R299 B.n654 B.n653 585
R300 B.n652 B.n27 585
R301 B.n651 B.n650 585
R302 B.n649 B.n28 585
R303 B.n648 B.n647 585
R304 B.n646 B.n29 585
R305 B.n645 B.n644 585
R306 B.n643 B.n30 585
R307 B.n642 B.n641 585
R308 B.n640 B.n31 585
R309 B.n639 B.n638 585
R310 B.n637 B.n32 585
R311 B.n636 B.n635 585
R312 B.n634 B.n33 585
R313 B.n633 B.n632 585
R314 B.n631 B.n34 585
R315 B.n630 B.n629 585
R316 B.n628 B.n35 585
R317 B.n627 B.n626 585
R318 B.n625 B.n36 585
R319 B.n624 B.n623 585
R320 B.n622 B.n37 585
R321 B.n621 B.n620 585
R322 B.n619 B.n38 585
R323 B.n618 B.n617 585
R324 B.n616 B.n39 585
R325 B.n615 B.n614 585
R326 B.n613 B.n40 585
R327 B.n612 B.n611 585
R328 B.n610 B.n41 585
R329 B.n609 B.n608 585
R330 B.n607 B.n42 585
R331 B.n606 B.n605 585
R332 B.n604 B.n43 585
R333 B.n603 B.n602 585
R334 B.n601 B.n600 585
R335 B.n599 B.n47 585
R336 B.n598 B.n597 585
R337 B.n596 B.n48 585
R338 B.n595 B.n594 585
R339 B.n593 B.n49 585
R340 B.n592 B.n591 585
R341 B.n590 B.n50 585
R342 B.n589 B.n588 585
R343 B.n587 B.n51 585
R344 B.n585 B.n584 585
R345 B.n583 B.n54 585
R346 B.n582 B.n581 585
R347 B.n580 B.n55 585
R348 B.n579 B.n578 585
R349 B.n577 B.n56 585
R350 B.n576 B.n575 585
R351 B.n574 B.n57 585
R352 B.n573 B.n572 585
R353 B.n571 B.n58 585
R354 B.n570 B.n569 585
R355 B.n568 B.n59 585
R356 B.n567 B.n566 585
R357 B.n565 B.n60 585
R358 B.n564 B.n563 585
R359 B.n562 B.n61 585
R360 B.n561 B.n560 585
R361 B.n559 B.n62 585
R362 B.n558 B.n557 585
R363 B.n556 B.n63 585
R364 B.n555 B.n554 585
R365 B.n553 B.n64 585
R366 B.n552 B.n551 585
R367 B.n550 B.n65 585
R368 B.n549 B.n548 585
R369 B.n547 B.n66 585
R370 B.n546 B.n545 585
R371 B.n544 B.n67 585
R372 B.n543 B.n542 585
R373 B.n541 B.n68 585
R374 B.n540 B.n539 585
R375 B.n538 B.n69 585
R376 B.n537 B.n536 585
R377 B.n535 B.n70 585
R378 B.n534 B.n533 585
R379 B.n532 B.n71 585
R380 B.n531 B.n530 585
R381 B.n529 B.n72 585
R382 B.n528 B.n527 585
R383 B.n526 B.n73 585
R384 B.n525 B.n524 585
R385 B.n523 B.n74 585
R386 B.n522 B.n521 585
R387 B.n520 B.n75 585
R388 B.n519 B.n518 585
R389 B.n517 B.n76 585
R390 B.n516 B.n515 585
R391 B.n514 B.n77 585
R392 B.n513 B.n512 585
R393 B.n511 B.n78 585
R394 B.n510 B.n509 585
R395 B.n508 B.n79 585
R396 B.n507 B.n506 585
R397 B.n505 B.n80 585
R398 B.n504 B.n503 585
R399 B.n502 B.n81 585
R400 B.n501 B.n500 585
R401 B.n499 B.n82 585
R402 B.n498 B.n497 585
R403 B.n496 B.n83 585
R404 B.n495 B.n494 585
R405 B.n694 B.n13 585
R406 B.n696 B.n695 585
R407 B.n697 B.n12 585
R408 B.n699 B.n698 585
R409 B.n700 B.n11 585
R410 B.n702 B.n701 585
R411 B.n703 B.n10 585
R412 B.n705 B.n704 585
R413 B.n706 B.n9 585
R414 B.n708 B.n707 585
R415 B.n709 B.n8 585
R416 B.n711 B.n710 585
R417 B.n712 B.n7 585
R418 B.n714 B.n713 585
R419 B.n715 B.n6 585
R420 B.n717 B.n716 585
R421 B.n718 B.n5 585
R422 B.n720 B.n719 585
R423 B.n721 B.n4 585
R424 B.n723 B.n722 585
R425 B.n724 B.n3 585
R426 B.n726 B.n725 585
R427 B.n727 B.n0 585
R428 B.n2 B.n1 585
R429 B.n188 B.n187 585
R430 B.n189 B.n186 585
R431 B.n191 B.n190 585
R432 B.n192 B.n185 585
R433 B.n194 B.n193 585
R434 B.n195 B.n184 585
R435 B.n197 B.n196 585
R436 B.n198 B.n183 585
R437 B.n200 B.n199 585
R438 B.n201 B.n182 585
R439 B.n203 B.n202 585
R440 B.n204 B.n181 585
R441 B.n206 B.n205 585
R442 B.n207 B.n180 585
R443 B.n209 B.n208 585
R444 B.n210 B.n179 585
R445 B.n212 B.n211 585
R446 B.n213 B.n178 585
R447 B.n215 B.n214 585
R448 B.n216 B.n177 585
R449 B.n218 B.n217 585
R450 B.n219 B.n176 585
R451 B.n220 B.n219 535.745
R452 B.n422 B.n421 535.745
R453 B.n494 B.n493 535.745
R454 B.n692 B.n13 535.745
R455 B.n729 B.n728 256.663
R456 B.n728 B.n727 235.042
R457 B.n728 B.n2 235.042
R458 B.n220 B.n175 163.367
R459 B.n224 B.n175 163.367
R460 B.n225 B.n224 163.367
R461 B.n226 B.n225 163.367
R462 B.n226 B.n173 163.367
R463 B.n230 B.n173 163.367
R464 B.n231 B.n230 163.367
R465 B.n232 B.n231 163.367
R466 B.n232 B.n171 163.367
R467 B.n236 B.n171 163.367
R468 B.n237 B.n236 163.367
R469 B.n238 B.n237 163.367
R470 B.n238 B.n169 163.367
R471 B.n242 B.n169 163.367
R472 B.n243 B.n242 163.367
R473 B.n244 B.n243 163.367
R474 B.n244 B.n167 163.367
R475 B.n248 B.n167 163.367
R476 B.n249 B.n248 163.367
R477 B.n250 B.n249 163.367
R478 B.n250 B.n165 163.367
R479 B.n254 B.n165 163.367
R480 B.n255 B.n254 163.367
R481 B.n256 B.n255 163.367
R482 B.n256 B.n163 163.367
R483 B.n260 B.n163 163.367
R484 B.n261 B.n260 163.367
R485 B.n262 B.n261 163.367
R486 B.n262 B.n161 163.367
R487 B.n266 B.n161 163.367
R488 B.n267 B.n266 163.367
R489 B.n268 B.n267 163.367
R490 B.n268 B.n159 163.367
R491 B.n272 B.n159 163.367
R492 B.n273 B.n272 163.367
R493 B.n274 B.n273 163.367
R494 B.n274 B.n157 163.367
R495 B.n278 B.n157 163.367
R496 B.n279 B.n278 163.367
R497 B.n280 B.n279 163.367
R498 B.n280 B.n155 163.367
R499 B.n284 B.n155 163.367
R500 B.n285 B.n284 163.367
R501 B.n286 B.n285 163.367
R502 B.n286 B.n153 163.367
R503 B.n290 B.n153 163.367
R504 B.n291 B.n290 163.367
R505 B.n292 B.n291 163.367
R506 B.n292 B.n151 163.367
R507 B.n296 B.n151 163.367
R508 B.n297 B.n296 163.367
R509 B.n298 B.n297 163.367
R510 B.n298 B.n149 163.367
R511 B.n302 B.n149 163.367
R512 B.n303 B.n302 163.367
R513 B.n304 B.n303 163.367
R514 B.n304 B.n147 163.367
R515 B.n308 B.n147 163.367
R516 B.n309 B.n308 163.367
R517 B.n310 B.n309 163.367
R518 B.n310 B.n143 163.367
R519 B.n315 B.n143 163.367
R520 B.n316 B.n315 163.367
R521 B.n317 B.n316 163.367
R522 B.n317 B.n141 163.367
R523 B.n321 B.n141 163.367
R524 B.n322 B.n321 163.367
R525 B.n323 B.n322 163.367
R526 B.n323 B.n139 163.367
R527 B.n330 B.n139 163.367
R528 B.n331 B.n330 163.367
R529 B.n332 B.n331 163.367
R530 B.n332 B.n137 163.367
R531 B.n336 B.n137 163.367
R532 B.n337 B.n336 163.367
R533 B.n338 B.n337 163.367
R534 B.n338 B.n135 163.367
R535 B.n342 B.n135 163.367
R536 B.n343 B.n342 163.367
R537 B.n344 B.n343 163.367
R538 B.n344 B.n133 163.367
R539 B.n348 B.n133 163.367
R540 B.n349 B.n348 163.367
R541 B.n350 B.n349 163.367
R542 B.n350 B.n131 163.367
R543 B.n354 B.n131 163.367
R544 B.n355 B.n354 163.367
R545 B.n356 B.n355 163.367
R546 B.n356 B.n129 163.367
R547 B.n360 B.n129 163.367
R548 B.n361 B.n360 163.367
R549 B.n362 B.n361 163.367
R550 B.n362 B.n127 163.367
R551 B.n366 B.n127 163.367
R552 B.n367 B.n366 163.367
R553 B.n368 B.n367 163.367
R554 B.n368 B.n125 163.367
R555 B.n372 B.n125 163.367
R556 B.n373 B.n372 163.367
R557 B.n374 B.n373 163.367
R558 B.n374 B.n123 163.367
R559 B.n378 B.n123 163.367
R560 B.n379 B.n378 163.367
R561 B.n380 B.n379 163.367
R562 B.n380 B.n121 163.367
R563 B.n384 B.n121 163.367
R564 B.n385 B.n384 163.367
R565 B.n386 B.n385 163.367
R566 B.n386 B.n119 163.367
R567 B.n390 B.n119 163.367
R568 B.n391 B.n390 163.367
R569 B.n392 B.n391 163.367
R570 B.n392 B.n117 163.367
R571 B.n396 B.n117 163.367
R572 B.n397 B.n396 163.367
R573 B.n398 B.n397 163.367
R574 B.n398 B.n115 163.367
R575 B.n402 B.n115 163.367
R576 B.n403 B.n402 163.367
R577 B.n404 B.n403 163.367
R578 B.n404 B.n113 163.367
R579 B.n408 B.n113 163.367
R580 B.n409 B.n408 163.367
R581 B.n410 B.n409 163.367
R582 B.n410 B.n111 163.367
R583 B.n414 B.n111 163.367
R584 B.n415 B.n414 163.367
R585 B.n416 B.n415 163.367
R586 B.n416 B.n109 163.367
R587 B.n420 B.n109 163.367
R588 B.n421 B.n420 163.367
R589 B.n493 B.n492 163.367
R590 B.n492 B.n85 163.367
R591 B.n488 B.n85 163.367
R592 B.n488 B.n487 163.367
R593 B.n487 B.n486 163.367
R594 B.n486 B.n87 163.367
R595 B.n482 B.n87 163.367
R596 B.n482 B.n481 163.367
R597 B.n481 B.n480 163.367
R598 B.n480 B.n89 163.367
R599 B.n476 B.n89 163.367
R600 B.n476 B.n475 163.367
R601 B.n475 B.n474 163.367
R602 B.n474 B.n91 163.367
R603 B.n470 B.n91 163.367
R604 B.n470 B.n469 163.367
R605 B.n469 B.n468 163.367
R606 B.n468 B.n93 163.367
R607 B.n464 B.n93 163.367
R608 B.n464 B.n463 163.367
R609 B.n463 B.n462 163.367
R610 B.n462 B.n95 163.367
R611 B.n458 B.n95 163.367
R612 B.n458 B.n457 163.367
R613 B.n457 B.n456 163.367
R614 B.n456 B.n97 163.367
R615 B.n452 B.n97 163.367
R616 B.n452 B.n451 163.367
R617 B.n451 B.n450 163.367
R618 B.n450 B.n99 163.367
R619 B.n446 B.n99 163.367
R620 B.n446 B.n445 163.367
R621 B.n445 B.n444 163.367
R622 B.n444 B.n101 163.367
R623 B.n440 B.n101 163.367
R624 B.n440 B.n439 163.367
R625 B.n439 B.n438 163.367
R626 B.n438 B.n103 163.367
R627 B.n434 B.n103 163.367
R628 B.n434 B.n433 163.367
R629 B.n433 B.n432 163.367
R630 B.n432 B.n105 163.367
R631 B.n428 B.n105 163.367
R632 B.n428 B.n427 163.367
R633 B.n427 B.n426 163.367
R634 B.n426 B.n107 163.367
R635 B.n422 B.n107 163.367
R636 B.n692 B.n691 163.367
R637 B.n691 B.n690 163.367
R638 B.n690 B.n15 163.367
R639 B.n686 B.n15 163.367
R640 B.n686 B.n685 163.367
R641 B.n685 B.n684 163.367
R642 B.n684 B.n17 163.367
R643 B.n680 B.n17 163.367
R644 B.n680 B.n679 163.367
R645 B.n679 B.n678 163.367
R646 B.n678 B.n19 163.367
R647 B.n674 B.n19 163.367
R648 B.n674 B.n673 163.367
R649 B.n673 B.n672 163.367
R650 B.n672 B.n21 163.367
R651 B.n668 B.n21 163.367
R652 B.n668 B.n667 163.367
R653 B.n667 B.n666 163.367
R654 B.n666 B.n23 163.367
R655 B.n662 B.n23 163.367
R656 B.n662 B.n661 163.367
R657 B.n661 B.n660 163.367
R658 B.n660 B.n25 163.367
R659 B.n656 B.n25 163.367
R660 B.n656 B.n655 163.367
R661 B.n655 B.n654 163.367
R662 B.n654 B.n27 163.367
R663 B.n650 B.n27 163.367
R664 B.n650 B.n649 163.367
R665 B.n649 B.n648 163.367
R666 B.n648 B.n29 163.367
R667 B.n644 B.n29 163.367
R668 B.n644 B.n643 163.367
R669 B.n643 B.n642 163.367
R670 B.n642 B.n31 163.367
R671 B.n638 B.n31 163.367
R672 B.n638 B.n637 163.367
R673 B.n637 B.n636 163.367
R674 B.n636 B.n33 163.367
R675 B.n632 B.n33 163.367
R676 B.n632 B.n631 163.367
R677 B.n631 B.n630 163.367
R678 B.n630 B.n35 163.367
R679 B.n626 B.n35 163.367
R680 B.n626 B.n625 163.367
R681 B.n625 B.n624 163.367
R682 B.n624 B.n37 163.367
R683 B.n620 B.n37 163.367
R684 B.n620 B.n619 163.367
R685 B.n619 B.n618 163.367
R686 B.n618 B.n39 163.367
R687 B.n614 B.n39 163.367
R688 B.n614 B.n613 163.367
R689 B.n613 B.n612 163.367
R690 B.n612 B.n41 163.367
R691 B.n608 B.n41 163.367
R692 B.n608 B.n607 163.367
R693 B.n607 B.n606 163.367
R694 B.n606 B.n43 163.367
R695 B.n602 B.n43 163.367
R696 B.n602 B.n601 163.367
R697 B.n601 B.n47 163.367
R698 B.n597 B.n47 163.367
R699 B.n597 B.n596 163.367
R700 B.n596 B.n595 163.367
R701 B.n595 B.n49 163.367
R702 B.n591 B.n49 163.367
R703 B.n591 B.n590 163.367
R704 B.n590 B.n589 163.367
R705 B.n589 B.n51 163.367
R706 B.n584 B.n51 163.367
R707 B.n584 B.n583 163.367
R708 B.n583 B.n582 163.367
R709 B.n582 B.n55 163.367
R710 B.n578 B.n55 163.367
R711 B.n578 B.n577 163.367
R712 B.n577 B.n576 163.367
R713 B.n576 B.n57 163.367
R714 B.n572 B.n57 163.367
R715 B.n572 B.n571 163.367
R716 B.n571 B.n570 163.367
R717 B.n570 B.n59 163.367
R718 B.n566 B.n59 163.367
R719 B.n566 B.n565 163.367
R720 B.n565 B.n564 163.367
R721 B.n564 B.n61 163.367
R722 B.n560 B.n61 163.367
R723 B.n560 B.n559 163.367
R724 B.n559 B.n558 163.367
R725 B.n558 B.n63 163.367
R726 B.n554 B.n63 163.367
R727 B.n554 B.n553 163.367
R728 B.n553 B.n552 163.367
R729 B.n552 B.n65 163.367
R730 B.n548 B.n65 163.367
R731 B.n548 B.n547 163.367
R732 B.n547 B.n546 163.367
R733 B.n546 B.n67 163.367
R734 B.n542 B.n67 163.367
R735 B.n542 B.n541 163.367
R736 B.n541 B.n540 163.367
R737 B.n540 B.n69 163.367
R738 B.n536 B.n69 163.367
R739 B.n536 B.n535 163.367
R740 B.n535 B.n534 163.367
R741 B.n534 B.n71 163.367
R742 B.n530 B.n71 163.367
R743 B.n530 B.n529 163.367
R744 B.n529 B.n528 163.367
R745 B.n528 B.n73 163.367
R746 B.n524 B.n73 163.367
R747 B.n524 B.n523 163.367
R748 B.n523 B.n522 163.367
R749 B.n522 B.n75 163.367
R750 B.n518 B.n75 163.367
R751 B.n518 B.n517 163.367
R752 B.n517 B.n516 163.367
R753 B.n516 B.n77 163.367
R754 B.n512 B.n77 163.367
R755 B.n512 B.n511 163.367
R756 B.n511 B.n510 163.367
R757 B.n510 B.n79 163.367
R758 B.n506 B.n79 163.367
R759 B.n506 B.n505 163.367
R760 B.n505 B.n504 163.367
R761 B.n504 B.n81 163.367
R762 B.n500 B.n81 163.367
R763 B.n500 B.n499 163.367
R764 B.n499 B.n498 163.367
R765 B.n498 B.n83 163.367
R766 B.n494 B.n83 163.367
R767 B.n696 B.n13 163.367
R768 B.n697 B.n696 163.367
R769 B.n698 B.n697 163.367
R770 B.n698 B.n11 163.367
R771 B.n702 B.n11 163.367
R772 B.n703 B.n702 163.367
R773 B.n704 B.n703 163.367
R774 B.n704 B.n9 163.367
R775 B.n708 B.n9 163.367
R776 B.n709 B.n708 163.367
R777 B.n710 B.n709 163.367
R778 B.n710 B.n7 163.367
R779 B.n714 B.n7 163.367
R780 B.n715 B.n714 163.367
R781 B.n716 B.n715 163.367
R782 B.n716 B.n5 163.367
R783 B.n720 B.n5 163.367
R784 B.n721 B.n720 163.367
R785 B.n722 B.n721 163.367
R786 B.n722 B.n3 163.367
R787 B.n726 B.n3 163.367
R788 B.n727 B.n726 163.367
R789 B.n188 B.n2 163.367
R790 B.n189 B.n188 163.367
R791 B.n190 B.n189 163.367
R792 B.n190 B.n185 163.367
R793 B.n194 B.n185 163.367
R794 B.n195 B.n194 163.367
R795 B.n196 B.n195 163.367
R796 B.n196 B.n183 163.367
R797 B.n200 B.n183 163.367
R798 B.n201 B.n200 163.367
R799 B.n202 B.n201 163.367
R800 B.n202 B.n181 163.367
R801 B.n206 B.n181 163.367
R802 B.n207 B.n206 163.367
R803 B.n208 B.n207 163.367
R804 B.n208 B.n179 163.367
R805 B.n212 B.n179 163.367
R806 B.n213 B.n212 163.367
R807 B.n214 B.n213 163.367
R808 B.n214 B.n177 163.367
R809 B.n218 B.n177 163.367
R810 B.n219 B.n218 163.367
R811 B.n326 B.t4 132.709
R812 B.n52 B.t11 132.709
R813 B.n144 B.t1 132.685
R814 B.n44 B.t8 132.685
R815 B.n327 B.t5 112.153
R816 B.n53 B.t10 112.153
R817 B.n145 B.t2 112.129
R818 B.n45 B.t7 112.129
R819 B.n312 B.n145 59.5399
R820 B.n328 B.n327 59.5399
R821 B.n586 B.n53 59.5399
R822 B.n46 B.n45 59.5399
R823 B.n694 B.n693 34.8103
R824 B.n495 B.n84 34.8103
R825 B.n423 B.n108 34.8103
R826 B.n221 B.n176 34.8103
R827 B.n145 B.n144 20.5581
R828 B.n327 B.n326 20.5581
R829 B.n53 B.n52 20.5581
R830 B.n45 B.n44 20.5581
R831 B B.n729 18.0485
R832 B.n695 B.n694 10.6151
R833 B.n695 B.n12 10.6151
R834 B.n699 B.n12 10.6151
R835 B.n700 B.n699 10.6151
R836 B.n701 B.n700 10.6151
R837 B.n701 B.n10 10.6151
R838 B.n705 B.n10 10.6151
R839 B.n706 B.n705 10.6151
R840 B.n707 B.n706 10.6151
R841 B.n707 B.n8 10.6151
R842 B.n711 B.n8 10.6151
R843 B.n712 B.n711 10.6151
R844 B.n713 B.n712 10.6151
R845 B.n713 B.n6 10.6151
R846 B.n717 B.n6 10.6151
R847 B.n718 B.n717 10.6151
R848 B.n719 B.n718 10.6151
R849 B.n719 B.n4 10.6151
R850 B.n723 B.n4 10.6151
R851 B.n724 B.n723 10.6151
R852 B.n725 B.n724 10.6151
R853 B.n725 B.n0 10.6151
R854 B.n693 B.n14 10.6151
R855 B.n689 B.n14 10.6151
R856 B.n689 B.n688 10.6151
R857 B.n688 B.n687 10.6151
R858 B.n687 B.n16 10.6151
R859 B.n683 B.n16 10.6151
R860 B.n683 B.n682 10.6151
R861 B.n682 B.n681 10.6151
R862 B.n681 B.n18 10.6151
R863 B.n677 B.n18 10.6151
R864 B.n677 B.n676 10.6151
R865 B.n676 B.n675 10.6151
R866 B.n675 B.n20 10.6151
R867 B.n671 B.n20 10.6151
R868 B.n671 B.n670 10.6151
R869 B.n670 B.n669 10.6151
R870 B.n669 B.n22 10.6151
R871 B.n665 B.n22 10.6151
R872 B.n665 B.n664 10.6151
R873 B.n664 B.n663 10.6151
R874 B.n663 B.n24 10.6151
R875 B.n659 B.n24 10.6151
R876 B.n659 B.n658 10.6151
R877 B.n658 B.n657 10.6151
R878 B.n657 B.n26 10.6151
R879 B.n653 B.n26 10.6151
R880 B.n653 B.n652 10.6151
R881 B.n652 B.n651 10.6151
R882 B.n651 B.n28 10.6151
R883 B.n647 B.n28 10.6151
R884 B.n647 B.n646 10.6151
R885 B.n646 B.n645 10.6151
R886 B.n645 B.n30 10.6151
R887 B.n641 B.n30 10.6151
R888 B.n641 B.n640 10.6151
R889 B.n640 B.n639 10.6151
R890 B.n639 B.n32 10.6151
R891 B.n635 B.n32 10.6151
R892 B.n635 B.n634 10.6151
R893 B.n634 B.n633 10.6151
R894 B.n633 B.n34 10.6151
R895 B.n629 B.n34 10.6151
R896 B.n629 B.n628 10.6151
R897 B.n628 B.n627 10.6151
R898 B.n627 B.n36 10.6151
R899 B.n623 B.n36 10.6151
R900 B.n623 B.n622 10.6151
R901 B.n622 B.n621 10.6151
R902 B.n621 B.n38 10.6151
R903 B.n617 B.n38 10.6151
R904 B.n617 B.n616 10.6151
R905 B.n616 B.n615 10.6151
R906 B.n615 B.n40 10.6151
R907 B.n611 B.n40 10.6151
R908 B.n611 B.n610 10.6151
R909 B.n610 B.n609 10.6151
R910 B.n609 B.n42 10.6151
R911 B.n605 B.n42 10.6151
R912 B.n605 B.n604 10.6151
R913 B.n604 B.n603 10.6151
R914 B.n600 B.n599 10.6151
R915 B.n599 B.n598 10.6151
R916 B.n598 B.n48 10.6151
R917 B.n594 B.n48 10.6151
R918 B.n594 B.n593 10.6151
R919 B.n593 B.n592 10.6151
R920 B.n592 B.n50 10.6151
R921 B.n588 B.n50 10.6151
R922 B.n588 B.n587 10.6151
R923 B.n585 B.n54 10.6151
R924 B.n581 B.n54 10.6151
R925 B.n581 B.n580 10.6151
R926 B.n580 B.n579 10.6151
R927 B.n579 B.n56 10.6151
R928 B.n575 B.n56 10.6151
R929 B.n575 B.n574 10.6151
R930 B.n574 B.n573 10.6151
R931 B.n573 B.n58 10.6151
R932 B.n569 B.n58 10.6151
R933 B.n569 B.n568 10.6151
R934 B.n568 B.n567 10.6151
R935 B.n567 B.n60 10.6151
R936 B.n563 B.n60 10.6151
R937 B.n563 B.n562 10.6151
R938 B.n562 B.n561 10.6151
R939 B.n561 B.n62 10.6151
R940 B.n557 B.n62 10.6151
R941 B.n557 B.n556 10.6151
R942 B.n556 B.n555 10.6151
R943 B.n555 B.n64 10.6151
R944 B.n551 B.n64 10.6151
R945 B.n551 B.n550 10.6151
R946 B.n550 B.n549 10.6151
R947 B.n549 B.n66 10.6151
R948 B.n545 B.n66 10.6151
R949 B.n545 B.n544 10.6151
R950 B.n544 B.n543 10.6151
R951 B.n543 B.n68 10.6151
R952 B.n539 B.n68 10.6151
R953 B.n539 B.n538 10.6151
R954 B.n538 B.n537 10.6151
R955 B.n537 B.n70 10.6151
R956 B.n533 B.n70 10.6151
R957 B.n533 B.n532 10.6151
R958 B.n532 B.n531 10.6151
R959 B.n531 B.n72 10.6151
R960 B.n527 B.n72 10.6151
R961 B.n527 B.n526 10.6151
R962 B.n526 B.n525 10.6151
R963 B.n525 B.n74 10.6151
R964 B.n521 B.n74 10.6151
R965 B.n521 B.n520 10.6151
R966 B.n520 B.n519 10.6151
R967 B.n519 B.n76 10.6151
R968 B.n515 B.n76 10.6151
R969 B.n515 B.n514 10.6151
R970 B.n514 B.n513 10.6151
R971 B.n513 B.n78 10.6151
R972 B.n509 B.n78 10.6151
R973 B.n509 B.n508 10.6151
R974 B.n508 B.n507 10.6151
R975 B.n507 B.n80 10.6151
R976 B.n503 B.n80 10.6151
R977 B.n503 B.n502 10.6151
R978 B.n502 B.n501 10.6151
R979 B.n501 B.n82 10.6151
R980 B.n497 B.n82 10.6151
R981 B.n497 B.n496 10.6151
R982 B.n496 B.n495 10.6151
R983 B.n491 B.n84 10.6151
R984 B.n491 B.n490 10.6151
R985 B.n490 B.n489 10.6151
R986 B.n489 B.n86 10.6151
R987 B.n485 B.n86 10.6151
R988 B.n485 B.n484 10.6151
R989 B.n484 B.n483 10.6151
R990 B.n483 B.n88 10.6151
R991 B.n479 B.n88 10.6151
R992 B.n479 B.n478 10.6151
R993 B.n478 B.n477 10.6151
R994 B.n477 B.n90 10.6151
R995 B.n473 B.n90 10.6151
R996 B.n473 B.n472 10.6151
R997 B.n472 B.n471 10.6151
R998 B.n471 B.n92 10.6151
R999 B.n467 B.n92 10.6151
R1000 B.n467 B.n466 10.6151
R1001 B.n466 B.n465 10.6151
R1002 B.n465 B.n94 10.6151
R1003 B.n461 B.n94 10.6151
R1004 B.n461 B.n460 10.6151
R1005 B.n460 B.n459 10.6151
R1006 B.n459 B.n96 10.6151
R1007 B.n455 B.n96 10.6151
R1008 B.n455 B.n454 10.6151
R1009 B.n454 B.n453 10.6151
R1010 B.n453 B.n98 10.6151
R1011 B.n449 B.n98 10.6151
R1012 B.n449 B.n448 10.6151
R1013 B.n448 B.n447 10.6151
R1014 B.n447 B.n100 10.6151
R1015 B.n443 B.n100 10.6151
R1016 B.n443 B.n442 10.6151
R1017 B.n442 B.n441 10.6151
R1018 B.n441 B.n102 10.6151
R1019 B.n437 B.n102 10.6151
R1020 B.n437 B.n436 10.6151
R1021 B.n436 B.n435 10.6151
R1022 B.n435 B.n104 10.6151
R1023 B.n431 B.n104 10.6151
R1024 B.n431 B.n430 10.6151
R1025 B.n430 B.n429 10.6151
R1026 B.n429 B.n106 10.6151
R1027 B.n425 B.n106 10.6151
R1028 B.n425 B.n424 10.6151
R1029 B.n424 B.n423 10.6151
R1030 B.n187 B.n1 10.6151
R1031 B.n187 B.n186 10.6151
R1032 B.n191 B.n186 10.6151
R1033 B.n192 B.n191 10.6151
R1034 B.n193 B.n192 10.6151
R1035 B.n193 B.n184 10.6151
R1036 B.n197 B.n184 10.6151
R1037 B.n198 B.n197 10.6151
R1038 B.n199 B.n198 10.6151
R1039 B.n199 B.n182 10.6151
R1040 B.n203 B.n182 10.6151
R1041 B.n204 B.n203 10.6151
R1042 B.n205 B.n204 10.6151
R1043 B.n205 B.n180 10.6151
R1044 B.n209 B.n180 10.6151
R1045 B.n210 B.n209 10.6151
R1046 B.n211 B.n210 10.6151
R1047 B.n211 B.n178 10.6151
R1048 B.n215 B.n178 10.6151
R1049 B.n216 B.n215 10.6151
R1050 B.n217 B.n216 10.6151
R1051 B.n217 B.n176 10.6151
R1052 B.n222 B.n221 10.6151
R1053 B.n223 B.n222 10.6151
R1054 B.n223 B.n174 10.6151
R1055 B.n227 B.n174 10.6151
R1056 B.n228 B.n227 10.6151
R1057 B.n229 B.n228 10.6151
R1058 B.n229 B.n172 10.6151
R1059 B.n233 B.n172 10.6151
R1060 B.n234 B.n233 10.6151
R1061 B.n235 B.n234 10.6151
R1062 B.n235 B.n170 10.6151
R1063 B.n239 B.n170 10.6151
R1064 B.n240 B.n239 10.6151
R1065 B.n241 B.n240 10.6151
R1066 B.n241 B.n168 10.6151
R1067 B.n245 B.n168 10.6151
R1068 B.n246 B.n245 10.6151
R1069 B.n247 B.n246 10.6151
R1070 B.n247 B.n166 10.6151
R1071 B.n251 B.n166 10.6151
R1072 B.n252 B.n251 10.6151
R1073 B.n253 B.n252 10.6151
R1074 B.n253 B.n164 10.6151
R1075 B.n257 B.n164 10.6151
R1076 B.n258 B.n257 10.6151
R1077 B.n259 B.n258 10.6151
R1078 B.n259 B.n162 10.6151
R1079 B.n263 B.n162 10.6151
R1080 B.n264 B.n263 10.6151
R1081 B.n265 B.n264 10.6151
R1082 B.n265 B.n160 10.6151
R1083 B.n269 B.n160 10.6151
R1084 B.n270 B.n269 10.6151
R1085 B.n271 B.n270 10.6151
R1086 B.n271 B.n158 10.6151
R1087 B.n275 B.n158 10.6151
R1088 B.n276 B.n275 10.6151
R1089 B.n277 B.n276 10.6151
R1090 B.n277 B.n156 10.6151
R1091 B.n281 B.n156 10.6151
R1092 B.n282 B.n281 10.6151
R1093 B.n283 B.n282 10.6151
R1094 B.n283 B.n154 10.6151
R1095 B.n287 B.n154 10.6151
R1096 B.n288 B.n287 10.6151
R1097 B.n289 B.n288 10.6151
R1098 B.n289 B.n152 10.6151
R1099 B.n293 B.n152 10.6151
R1100 B.n294 B.n293 10.6151
R1101 B.n295 B.n294 10.6151
R1102 B.n295 B.n150 10.6151
R1103 B.n299 B.n150 10.6151
R1104 B.n300 B.n299 10.6151
R1105 B.n301 B.n300 10.6151
R1106 B.n301 B.n148 10.6151
R1107 B.n305 B.n148 10.6151
R1108 B.n306 B.n305 10.6151
R1109 B.n307 B.n306 10.6151
R1110 B.n307 B.n146 10.6151
R1111 B.n311 B.n146 10.6151
R1112 B.n314 B.n313 10.6151
R1113 B.n314 B.n142 10.6151
R1114 B.n318 B.n142 10.6151
R1115 B.n319 B.n318 10.6151
R1116 B.n320 B.n319 10.6151
R1117 B.n320 B.n140 10.6151
R1118 B.n324 B.n140 10.6151
R1119 B.n325 B.n324 10.6151
R1120 B.n329 B.n325 10.6151
R1121 B.n333 B.n138 10.6151
R1122 B.n334 B.n333 10.6151
R1123 B.n335 B.n334 10.6151
R1124 B.n335 B.n136 10.6151
R1125 B.n339 B.n136 10.6151
R1126 B.n340 B.n339 10.6151
R1127 B.n341 B.n340 10.6151
R1128 B.n341 B.n134 10.6151
R1129 B.n345 B.n134 10.6151
R1130 B.n346 B.n345 10.6151
R1131 B.n347 B.n346 10.6151
R1132 B.n347 B.n132 10.6151
R1133 B.n351 B.n132 10.6151
R1134 B.n352 B.n351 10.6151
R1135 B.n353 B.n352 10.6151
R1136 B.n353 B.n130 10.6151
R1137 B.n357 B.n130 10.6151
R1138 B.n358 B.n357 10.6151
R1139 B.n359 B.n358 10.6151
R1140 B.n359 B.n128 10.6151
R1141 B.n363 B.n128 10.6151
R1142 B.n364 B.n363 10.6151
R1143 B.n365 B.n364 10.6151
R1144 B.n365 B.n126 10.6151
R1145 B.n369 B.n126 10.6151
R1146 B.n370 B.n369 10.6151
R1147 B.n371 B.n370 10.6151
R1148 B.n371 B.n124 10.6151
R1149 B.n375 B.n124 10.6151
R1150 B.n376 B.n375 10.6151
R1151 B.n377 B.n376 10.6151
R1152 B.n377 B.n122 10.6151
R1153 B.n381 B.n122 10.6151
R1154 B.n382 B.n381 10.6151
R1155 B.n383 B.n382 10.6151
R1156 B.n383 B.n120 10.6151
R1157 B.n387 B.n120 10.6151
R1158 B.n388 B.n387 10.6151
R1159 B.n389 B.n388 10.6151
R1160 B.n389 B.n118 10.6151
R1161 B.n393 B.n118 10.6151
R1162 B.n394 B.n393 10.6151
R1163 B.n395 B.n394 10.6151
R1164 B.n395 B.n116 10.6151
R1165 B.n399 B.n116 10.6151
R1166 B.n400 B.n399 10.6151
R1167 B.n401 B.n400 10.6151
R1168 B.n401 B.n114 10.6151
R1169 B.n405 B.n114 10.6151
R1170 B.n406 B.n405 10.6151
R1171 B.n407 B.n406 10.6151
R1172 B.n407 B.n112 10.6151
R1173 B.n411 B.n112 10.6151
R1174 B.n412 B.n411 10.6151
R1175 B.n413 B.n412 10.6151
R1176 B.n413 B.n110 10.6151
R1177 B.n417 B.n110 10.6151
R1178 B.n418 B.n417 10.6151
R1179 B.n419 B.n418 10.6151
R1180 B.n419 B.n108 10.6151
R1181 B.n603 B.n46 9.36635
R1182 B.n586 B.n585 9.36635
R1183 B.n312 B.n311 9.36635
R1184 B.n328 B.n138 9.36635
R1185 B.n729 B.n0 8.11757
R1186 B.n729 B.n1 8.11757
R1187 B.n600 B.n46 1.24928
R1188 B.n587 B.n586 1.24928
R1189 B.n313 B.n312 1.24928
R1190 B.n329 B.n328 1.24928
R1191 VN.n3 VN.t4 693.812
R1192 VN.n13 VN.t0 693.812
R1193 VN.n2 VN.t2 670.509
R1194 VN.n6 VN.t5 670.509
R1195 VN.n8 VN.t3 670.509
R1196 VN.n12 VN.t6 670.509
R1197 VN.n16 VN.t1 670.509
R1198 VN.n18 VN.t7 670.509
R1199 VN.n9 VN.n8 161.3
R1200 VN.n19 VN.n18 161.3
R1201 VN.n17 VN.n10 161.3
R1202 VN.n16 VN.n15 161.3
R1203 VN.n14 VN.n11 161.3
R1204 VN.n7 VN.n0 161.3
R1205 VN.n6 VN.n5 161.3
R1206 VN.n4 VN.n1 161.3
R1207 VN VN.n19 47.6085
R1208 VN.n14 VN.n13 44.8907
R1209 VN.n4 VN.n3 44.8907
R1210 VN.n8 VN.n7 32.8641
R1211 VN.n18 VN.n17 32.8641
R1212 VN.n2 VN.n1 24.1005
R1213 VN.n6 VN.n1 24.1005
R1214 VN.n16 VN.n11 24.1005
R1215 VN.n12 VN.n11 24.1005
R1216 VN.n3 VN.n2 18.4104
R1217 VN.n13 VN.n12 18.4104
R1218 VN.n7 VN.n6 15.3369
R1219 VN.n17 VN.n16 15.3369
R1220 VN.n19 VN.n10 0.189894
R1221 VN.n15 VN.n10 0.189894
R1222 VN.n15 VN.n14 0.189894
R1223 VN.n5 VN.n4 0.189894
R1224 VN.n5 VN.n0 0.189894
R1225 VN.n9 VN.n0 0.189894
R1226 VN VN.n9 0.0516364
R1227 VDD2.n2 VDD2.n1 70.2914
R1228 VDD2.n2 VDD2.n0 70.2914
R1229 VDD2 VDD2.n5 70.2886
R1230 VDD2.n4 VDD2.n3 69.8901
R1231 VDD2.n4 VDD2.n2 43.9222
R1232 VDD2.n5 VDD2.t1 1.74153
R1233 VDD2.n5 VDD2.t7 1.74153
R1234 VDD2.n3 VDD2.t0 1.74153
R1235 VDD2.n3 VDD2.t6 1.74153
R1236 VDD2.n1 VDD2.t2 1.74153
R1237 VDD2.n1 VDD2.t4 1.74153
R1238 VDD2.n0 VDD2.t3 1.74153
R1239 VDD2.n0 VDD2.t5 1.74153
R1240 VDD2 VDD2.n4 0.515586
C0 VDD1 w_n2030_n4702# 1.48541f
C1 VTAIL B 5.67336f
C2 B w_n2030_n4702# 9.12407f
C3 VTAIL w_n2030_n4702# 5.87317f
C4 VDD2 VP 0.320338f
C5 VN VP 6.60996f
C6 VDD1 VP 8.72172f
C7 VDD2 VN 8.54983f
C8 VP B 1.28935f
C9 VDD2 VDD1 0.838674f
C10 VDD2 B 1.29646f
C11 VDD1 VN 0.148002f
C12 VN B 0.86678f
C13 VTAIL VP 8.07104f
C14 VP w_n2030_n4702# 3.99462f
C15 VDD1 B 1.25888f
C16 VDD2 VTAIL 15.7674f
C17 VDD2 w_n2030_n4702# 1.5215f
C18 VTAIL VN 8.05693f
C19 VN w_n2030_n4702# 3.7366f
C20 VDD1 VTAIL 15.7255f
C21 VDD2 VSUBS 1.525318f
C22 VDD1 VSUBS 1.83556f
C23 VTAIL VSUBS 1.19951f
C24 VN VSUBS 5.21281f
C25 VP VSUBS 1.922233f
C26 B VSUBS 3.484318f
C27 w_n2030_n4702# VSUBS 0.11666p
C28 VDD2.t3 VSUBS 0.403072f
C29 VDD2.t5 VSUBS 0.403072f
C30 VDD2.n0 VSUBS 3.37273f
C31 VDD2.t2 VSUBS 0.403072f
C32 VDD2.t4 VSUBS 0.403072f
C33 VDD2.n1 VSUBS 3.37273f
C34 VDD2.n2 VSUBS 3.46562f
C35 VDD2.t0 VSUBS 0.403072f
C36 VDD2.t6 VSUBS 0.403072f
C37 VDD2.n3 VSUBS 3.36894f
C38 VDD2.n4 VSUBS 3.3836f
C39 VDD2.t1 VSUBS 0.403072f
C40 VDD2.t7 VSUBS 0.403072f
C41 VDD2.n5 VSUBS 3.37269f
C42 VN.n0 VSUBS 0.049763f
C43 VN.n1 VSUBS 0.011292f
C44 VN.t4 VSUBS 1.94667f
C45 VN.t2 VSUBS 1.92242f
C46 VN.n2 VSUBS 0.726635f
C47 VN.n3 VSUBS 0.702211f
C48 VN.n4 VSUBS 0.210587f
C49 VN.n5 VSUBS 0.049763f
C50 VN.t5 VSUBS 1.92242f
C51 VN.n6 VSUBS 0.721069f
C52 VN.n7 VSUBS 0.011292f
C53 VN.t3 VSUBS 1.92242f
C54 VN.n8 VSUBS 0.719689f
C55 VN.n9 VSUBS 0.038564f
C56 VN.n10 VSUBS 0.049763f
C57 VN.n11 VSUBS 0.011292f
C58 VN.t1 VSUBS 1.92242f
C59 VN.t0 VSUBS 1.94667f
C60 VN.t6 VSUBS 1.92242f
C61 VN.n12 VSUBS 0.726635f
C62 VN.n13 VSUBS 0.702211f
C63 VN.n14 VSUBS 0.210587f
C64 VN.n15 VSUBS 0.049763f
C65 VN.n16 VSUBS 0.721069f
C66 VN.n17 VSUBS 0.011292f
C67 VN.t7 VSUBS 1.92242f
C68 VN.n18 VSUBS 0.719689f
C69 VN.n19 VSUBS 2.5123f
C70 B.n0 VSUBS 0.006727f
C71 B.n1 VSUBS 0.006727f
C72 B.n2 VSUBS 0.009948f
C73 B.n3 VSUBS 0.007623f
C74 B.n4 VSUBS 0.007623f
C75 B.n5 VSUBS 0.007623f
C76 B.n6 VSUBS 0.007623f
C77 B.n7 VSUBS 0.007623f
C78 B.n8 VSUBS 0.007623f
C79 B.n9 VSUBS 0.007623f
C80 B.n10 VSUBS 0.007623f
C81 B.n11 VSUBS 0.007623f
C82 B.n12 VSUBS 0.007623f
C83 B.n13 VSUBS 0.018085f
C84 B.n14 VSUBS 0.007623f
C85 B.n15 VSUBS 0.007623f
C86 B.n16 VSUBS 0.007623f
C87 B.n17 VSUBS 0.007623f
C88 B.n18 VSUBS 0.007623f
C89 B.n19 VSUBS 0.007623f
C90 B.n20 VSUBS 0.007623f
C91 B.n21 VSUBS 0.007623f
C92 B.n22 VSUBS 0.007623f
C93 B.n23 VSUBS 0.007623f
C94 B.n24 VSUBS 0.007623f
C95 B.n25 VSUBS 0.007623f
C96 B.n26 VSUBS 0.007623f
C97 B.n27 VSUBS 0.007623f
C98 B.n28 VSUBS 0.007623f
C99 B.n29 VSUBS 0.007623f
C100 B.n30 VSUBS 0.007623f
C101 B.n31 VSUBS 0.007623f
C102 B.n32 VSUBS 0.007623f
C103 B.n33 VSUBS 0.007623f
C104 B.n34 VSUBS 0.007623f
C105 B.n35 VSUBS 0.007623f
C106 B.n36 VSUBS 0.007623f
C107 B.n37 VSUBS 0.007623f
C108 B.n38 VSUBS 0.007623f
C109 B.n39 VSUBS 0.007623f
C110 B.n40 VSUBS 0.007623f
C111 B.n41 VSUBS 0.007623f
C112 B.n42 VSUBS 0.007623f
C113 B.n43 VSUBS 0.007623f
C114 B.t7 VSUBS 0.688181f
C115 B.t8 VSUBS 0.697357f
C116 B.t6 VSUBS 0.598646f
C117 B.n44 VSUBS 0.212272f
C118 B.n45 VSUBS 0.070101f
C119 B.n46 VSUBS 0.017663f
C120 B.n47 VSUBS 0.007623f
C121 B.n48 VSUBS 0.007623f
C122 B.n49 VSUBS 0.007623f
C123 B.n50 VSUBS 0.007623f
C124 B.n51 VSUBS 0.007623f
C125 B.t10 VSUBS 0.688155f
C126 B.t11 VSUBS 0.697333f
C127 B.t9 VSUBS 0.598646f
C128 B.n52 VSUBS 0.212296f
C129 B.n53 VSUBS 0.070127f
C130 B.n54 VSUBS 0.007623f
C131 B.n55 VSUBS 0.007623f
C132 B.n56 VSUBS 0.007623f
C133 B.n57 VSUBS 0.007623f
C134 B.n58 VSUBS 0.007623f
C135 B.n59 VSUBS 0.007623f
C136 B.n60 VSUBS 0.007623f
C137 B.n61 VSUBS 0.007623f
C138 B.n62 VSUBS 0.007623f
C139 B.n63 VSUBS 0.007623f
C140 B.n64 VSUBS 0.007623f
C141 B.n65 VSUBS 0.007623f
C142 B.n66 VSUBS 0.007623f
C143 B.n67 VSUBS 0.007623f
C144 B.n68 VSUBS 0.007623f
C145 B.n69 VSUBS 0.007623f
C146 B.n70 VSUBS 0.007623f
C147 B.n71 VSUBS 0.007623f
C148 B.n72 VSUBS 0.007623f
C149 B.n73 VSUBS 0.007623f
C150 B.n74 VSUBS 0.007623f
C151 B.n75 VSUBS 0.007623f
C152 B.n76 VSUBS 0.007623f
C153 B.n77 VSUBS 0.007623f
C154 B.n78 VSUBS 0.007623f
C155 B.n79 VSUBS 0.007623f
C156 B.n80 VSUBS 0.007623f
C157 B.n81 VSUBS 0.007623f
C158 B.n82 VSUBS 0.007623f
C159 B.n83 VSUBS 0.007623f
C160 B.n84 VSUBS 0.018085f
C161 B.n85 VSUBS 0.007623f
C162 B.n86 VSUBS 0.007623f
C163 B.n87 VSUBS 0.007623f
C164 B.n88 VSUBS 0.007623f
C165 B.n89 VSUBS 0.007623f
C166 B.n90 VSUBS 0.007623f
C167 B.n91 VSUBS 0.007623f
C168 B.n92 VSUBS 0.007623f
C169 B.n93 VSUBS 0.007623f
C170 B.n94 VSUBS 0.007623f
C171 B.n95 VSUBS 0.007623f
C172 B.n96 VSUBS 0.007623f
C173 B.n97 VSUBS 0.007623f
C174 B.n98 VSUBS 0.007623f
C175 B.n99 VSUBS 0.007623f
C176 B.n100 VSUBS 0.007623f
C177 B.n101 VSUBS 0.007623f
C178 B.n102 VSUBS 0.007623f
C179 B.n103 VSUBS 0.007623f
C180 B.n104 VSUBS 0.007623f
C181 B.n105 VSUBS 0.007623f
C182 B.n106 VSUBS 0.007623f
C183 B.n107 VSUBS 0.007623f
C184 B.n108 VSUBS 0.018291f
C185 B.n109 VSUBS 0.007623f
C186 B.n110 VSUBS 0.007623f
C187 B.n111 VSUBS 0.007623f
C188 B.n112 VSUBS 0.007623f
C189 B.n113 VSUBS 0.007623f
C190 B.n114 VSUBS 0.007623f
C191 B.n115 VSUBS 0.007623f
C192 B.n116 VSUBS 0.007623f
C193 B.n117 VSUBS 0.007623f
C194 B.n118 VSUBS 0.007623f
C195 B.n119 VSUBS 0.007623f
C196 B.n120 VSUBS 0.007623f
C197 B.n121 VSUBS 0.007623f
C198 B.n122 VSUBS 0.007623f
C199 B.n123 VSUBS 0.007623f
C200 B.n124 VSUBS 0.007623f
C201 B.n125 VSUBS 0.007623f
C202 B.n126 VSUBS 0.007623f
C203 B.n127 VSUBS 0.007623f
C204 B.n128 VSUBS 0.007623f
C205 B.n129 VSUBS 0.007623f
C206 B.n130 VSUBS 0.007623f
C207 B.n131 VSUBS 0.007623f
C208 B.n132 VSUBS 0.007623f
C209 B.n133 VSUBS 0.007623f
C210 B.n134 VSUBS 0.007623f
C211 B.n135 VSUBS 0.007623f
C212 B.n136 VSUBS 0.007623f
C213 B.n137 VSUBS 0.007623f
C214 B.n138 VSUBS 0.007175f
C215 B.n139 VSUBS 0.007623f
C216 B.n140 VSUBS 0.007623f
C217 B.n141 VSUBS 0.007623f
C218 B.n142 VSUBS 0.007623f
C219 B.n143 VSUBS 0.007623f
C220 B.t2 VSUBS 0.688181f
C221 B.t1 VSUBS 0.697357f
C222 B.t0 VSUBS 0.598646f
C223 B.n144 VSUBS 0.212272f
C224 B.n145 VSUBS 0.070101f
C225 B.n146 VSUBS 0.007623f
C226 B.n147 VSUBS 0.007623f
C227 B.n148 VSUBS 0.007623f
C228 B.n149 VSUBS 0.007623f
C229 B.n150 VSUBS 0.007623f
C230 B.n151 VSUBS 0.007623f
C231 B.n152 VSUBS 0.007623f
C232 B.n153 VSUBS 0.007623f
C233 B.n154 VSUBS 0.007623f
C234 B.n155 VSUBS 0.007623f
C235 B.n156 VSUBS 0.007623f
C236 B.n157 VSUBS 0.007623f
C237 B.n158 VSUBS 0.007623f
C238 B.n159 VSUBS 0.007623f
C239 B.n160 VSUBS 0.007623f
C240 B.n161 VSUBS 0.007623f
C241 B.n162 VSUBS 0.007623f
C242 B.n163 VSUBS 0.007623f
C243 B.n164 VSUBS 0.007623f
C244 B.n165 VSUBS 0.007623f
C245 B.n166 VSUBS 0.007623f
C246 B.n167 VSUBS 0.007623f
C247 B.n168 VSUBS 0.007623f
C248 B.n169 VSUBS 0.007623f
C249 B.n170 VSUBS 0.007623f
C250 B.n171 VSUBS 0.007623f
C251 B.n172 VSUBS 0.007623f
C252 B.n173 VSUBS 0.007623f
C253 B.n174 VSUBS 0.007623f
C254 B.n175 VSUBS 0.007623f
C255 B.n176 VSUBS 0.018085f
C256 B.n177 VSUBS 0.007623f
C257 B.n178 VSUBS 0.007623f
C258 B.n179 VSUBS 0.007623f
C259 B.n180 VSUBS 0.007623f
C260 B.n181 VSUBS 0.007623f
C261 B.n182 VSUBS 0.007623f
C262 B.n183 VSUBS 0.007623f
C263 B.n184 VSUBS 0.007623f
C264 B.n185 VSUBS 0.007623f
C265 B.n186 VSUBS 0.007623f
C266 B.n187 VSUBS 0.007623f
C267 B.n188 VSUBS 0.007623f
C268 B.n189 VSUBS 0.007623f
C269 B.n190 VSUBS 0.007623f
C270 B.n191 VSUBS 0.007623f
C271 B.n192 VSUBS 0.007623f
C272 B.n193 VSUBS 0.007623f
C273 B.n194 VSUBS 0.007623f
C274 B.n195 VSUBS 0.007623f
C275 B.n196 VSUBS 0.007623f
C276 B.n197 VSUBS 0.007623f
C277 B.n198 VSUBS 0.007623f
C278 B.n199 VSUBS 0.007623f
C279 B.n200 VSUBS 0.007623f
C280 B.n201 VSUBS 0.007623f
C281 B.n202 VSUBS 0.007623f
C282 B.n203 VSUBS 0.007623f
C283 B.n204 VSUBS 0.007623f
C284 B.n205 VSUBS 0.007623f
C285 B.n206 VSUBS 0.007623f
C286 B.n207 VSUBS 0.007623f
C287 B.n208 VSUBS 0.007623f
C288 B.n209 VSUBS 0.007623f
C289 B.n210 VSUBS 0.007623f
C290 B.n211 VSUBS 0.007623f
C291 B.n212 VSUBS 0.007623f
C292 B.n213 VSUBS 0.007623f
C293 B.n214 VSUBS 0.007623f
C294 B.n215 VSUBS 0.007623f
C295 B.n216 VSUBS 0.007623f
C296 B.n217 VSUBS 0.007623f
C297 B.n218 VSUBS 0.007623f
C298 B.n219 VSUBS 0.018085f
C299 B.n220 VSUBS 0.019136f
C300 B.n221 VSUBS 0.019136f
C301 B.n222 VSUBS 0.007623f
C302 B.n223 VSUBS 0.007623f
C303 B.n224 VSUBS 0.007623f
C304 B.n225 VSUBS 0.007623f
C305 B.n226 VSUBS 0.007623f
C306 B.n227 VSUBS 0.007623f
C307 B.n228 VSUBS 0.007623f
C308 B.n229 VSUBS 0.007623f
C309 B.n230 VSUBS 0.007623f
C310 B.n231 VSUBS 0.007623f
C311 B.n232 VSUBS 0.007623f
C312 B.n233 VSUBS 0.007623f
C313 B.n234 VSUBS 0.007623f
C314 B.n235 VSUBS 0.007623f
C315 B.n236 VSUBS 0.007623f
C316 B.n237 VSUBS 0.007623f
C317 B.n238 VSUBS 0.007623f
C318 B.n239 VSUBS 0.007623f
C319 B.n240 VSUBS 0.007623f
C320 B.n241 VSUBS 0.007623f
C321 B.n242 VSUBS 0.007623f
C322 B.n243 VSUBS 0.007623f
C323 B.n244 VSUBS 0.007623f
C324 B.n245 VSUBS 0.007623f
C325 B.n246 VSUBS 0.007623f
C326 B.n247 VSUBS 0.007623f
C327 B.n248 VSUBS 0.007623f
C328 B.n249 VSUBS 0.007623f
C329 B.n250 VSUBS 0.007623f
C330 B.n251 VSUBS 0.007623f
C331 B.n252 VSUBS 0.007623f
C332 B.n253 VSUBS 0.007623f
C333 B.n254 VSUBS 0.007623f
C334 B.n255 VSUBS 0.007623f
C335 B.n256 VSUBS 0.007623f
C336 B.n257 VSUBS 0.007623f
C337 B.n258 VSUBS 0.007623f
C338 B.n259 VSUBS 0.007623f
C339 B.n260 VSUBS 0.007623f
C340 B.n261 VSUBS 0.007623f
C341 B.n262 VSUBS 0.007623f
C342 B.n263 VSUBS 0.007623f
C343 B.n264 VSUBS 0.007623f
C344 B.n265 VSUBS 0.007623f
C345 B.n266 VSUBS 0.007623f
C346 B.n267 VSUBS 0.007623f
C347 B.n268 VSUBS 0.007623f
C348 B.n269 VSUBS 0.007623f
C349 B.n270 VSUBS 0.007623f
C350 B.n271 VSUBS 0.007623f
C351 B.n272 VSUBS 0.007623f
C352 B.n273 VSUBS 0.007623f
C353 B.n274 VSUBS 0.007623f
C354 B.n275 VSUBS 0.007623f
C355 B.n276 VSUBS 0.007623f
C356 B.n277 VSUBS 0.007623f
C357 B.n278 VSUBS 0.007623f
C358 B.n279 VSUBS 0.007623f
C359 B.n280 VSUBS 0.007623f
C360 B.n281 VSUBS 0.007623f
C361 B.n282 VSUBS 0.007623f
C362 B.n283 VSUBS 0.007623f
C363 B.n284 VSUBS 0.007623f
C364 B.n285 VSUBS 0.007623f
C365 B.n286 VSUBS 0.007623f
C366 B.n287 VSUBS 0.007623f
C367 B.n288 VSUBS 0.007623f
C368 B.n289 VSUBS 0.007623f
C369 B.n290 VSUBS 0.007623f
C370 B.n291 VSUBS 0.007623f
C371 B.n292 VSUBS 0.007623f
C372 B.n293 VSUBS 0.007623f
C373 B.n294 VSUBS 0.007623f
C374 B.n295 VSUBS 0.007623f
C375 B.n296 VSUBS 0.007623f
C376 B.n297 VSUBS 0.007623f
C377 B.n298 VSUBS 0.007623f
C378 B.n299 VSUBS 0.007623f
C379 B.n300 VSUBS 0.007623f
C380 B.n301 VSUBS 0.007623f
C381 B.n302 VSUBS 0.007623f
C382 B.n303 VSUBS 0.007623f
C383 B.n304 VSUBS 0.007623f
C384 B.n305 VSUBS 0.007623f
C385 B.n306 VSUBS 0.007623f
C386 B.n307 VSUBS 0.007623f
C387 B.n308 VSUBS 0.007623f
C388 B.n309 VSUBS 0.007623f
C389 B.n310 VSUBS 0.007623f
C390 B.n311 VSUBS 0.007175f
C391 B.n312 VSUBS 0.017663f
C392 B.n313 VSUBS 0.00426f
C393 B.n314 VSUBS 0.007623f
C394 B.n315 VSUBS 0.007623f
C395 B.n316 VSUBS 0.007623f
C396 B.n317 VSUBS 0.007623f
C397 B.n318 VSUBS 0.007623f
C398 B.n319 VSUBS 0.007623f
C399 B.n320 VSUBS 0.007623f
C400 B.n321 VSUBS 0.007623f
C401 B.n322 VSUBS 0.007623f
C402 B.n323 VSUBS 0.007623f
C403 B.n324 VSUBS 0.007623f
C404 B.n325 VSUBS 0.007623f
C405 B.t5 VSUBS 0.688155f
C406 B.t4 VSUBS 0.697333f
C407 B.t3 VSUBS 0.598646f
C408 B.n326 VSUBS 0.212296f
C409 B.n327 VSUBS 0.070127f
C410 B.n328 VSUBS 0.017663f
C411 B.n329 VSUBS 0.00426f
C412 B.n330 VSUBS 0.007623f
C413 B.n331 VSUBS 0.007623f
C414 B.n332 VSUBS 0.007623f
C415 B.n333 VSUBS 0.007623f
C416 B.n334 VSUBS 0.007623f
C417 B.n335 VSUBS 0.007623f
C418 B.n336 VSUBS 0.007623f
C419 B.n337 VSUBS 0.007623f
C420 B.n338 VSUBS 0.007623f
C421 B.n339 VSUBS 0.007623f
C422 B.n340 VSUBS 0.007623f
C423 B.n341 VSUBS 0.007623f
C424 B.n342 VSUBS 0.007623f
C425 B.n343 VSUBS 0.007623f
C426 B.n344 VSUBS 0.007623f
C427 B.n345 VSUBS 0.007623f
C428 B.n346 VSUBS 0.007623f
C429 B.n347 VSUBS 0.007623f
C430 B.n348 VSUBS 0.007623f
C431 B.n349 VSUBS 0.007623f
C432 B.n350 VSUBS 0.007623f
C433 B.n351 VSUBS 0.007623f
C434 B.n352 VSUBS 0.007623f
C435 B.n353 VSUBS 0.007623f
C436 B.n354 VSUBS 0.007623f
C437 B.n355 VSUBS 0.007623f
C438 B.n356 VSUBS 0.007623f
C439 B.n357 VSUBS 0.007623f
C440 B.n358 VSUBS 0.007623f
C441 B.n359 VSUBS 0.007623f
C442 B.n360 VSUBS 0.007623f
C443 B.n361 VSUBS 0.007623f
C444 B.n362 VSUBS 0.007623f
C445 B.n363 VSUBS 0.007623f
C446 B.n364 VSUBS 0.007623f
C447 B.n365 VSUBS 0.007623f
C448 B.n366 VSUBS 0.007623f
C449 B.n367 VSUBS 0.007623f
C450 B.n368 VSUBS 0.007623f
C451 B.n369 VSUBS 0.007623f
C452 B.n370 VSUBS 0.007623f
C453 B.n371 VSUBS 0.007623f
C454 B.n372 VSUBS 0.007623f
C455 B.n373 VSUBS 0.007623f
C456 B.n374 VSUBS 0.007623f
C457 B.n375 VSUBS 0.007623f
C458 B.n376 VSUBS 0.007623f
C459 B.n377 VSUBS 0.007623f
C460 B.n378 VSUBS 0.007623f
C461 B.n379 VSUBS 0.007623f
C462 B.n380 VSUBS 0.007623f
C463 B.n381 VSUBS 0.007623f
C464 B.n382 VSUBS 0.007623f
C465 B.n383 VSUBS 0.007623f
C466 B.n384 VSUBS 0.007623f
C467 B.n385 VSUBS 0.007623f
C468 B.n386 VSUBS 0.007623f
C469 B.n387 VSUBS 0.007623f
C470 B.n388 VSUBS 0.007623f
C471 B.n389 VSUBS 0.007623f
C472 B.n390 VSUBS 0.007623f
C473 B.n391 VSUBS 0.007623f
C474 B.n392 VSUBS 0.007623f
C475 B.n393 VSUBS 0.007623f
C476 B.n394 VSUBS 0.007623f
C477 B.n395 VSUBS 0.007623f
C478 B.n396 VSUBS 0.007623f
C479 B.n397 VSUBS 0.007623f
C480 B.n398 VSUBS 0.007623f
C481 B.n399 VSUBS 0.007623f
C482 B.n400 VSUBS 0.007623f
C483 B.n401 VSUBS 0.007623f
C484 B.n402 VSUBS 0.007623f
C485 B.n403 VSUBS 0.007623f
C486 B.n404 VSUBS 0.007623f
C487 B.n405 VSUBS 0.007623f
C488 B.n406 VSUBS 0.007623f
C489 B.n407 VSUBS 0.007623f
C490 B.n408 VSUBS 0.007623f
C491 B.n409 VSUBS 0.007623f
C492 B.n410 VSUBS 0.007623f
C493 B.n411 VSUBS 0.007623f
C494 B.n412 VSUBS 0.007623f
C495 B.n413 VSUBS 0.007623f
C496 B.n414 VSUBS 0.007623f
C497 B.n415 VSUBS 0.007623f
C498 B.n416 VSUBS 0.007623f
C499 B.n417 VSUBS 0.007623f
C500 B.n418 VSUBS 0.007623f
C501 B.n419 VSUBS 0.007623f
C502 B.n420 VSUBS 0.007623f
C503 B.n421 VSUBS 0.019136f
C504 B.n422 VSUBS 0.018085f
C505 B.n423 VSUBS 0.01893f
C506 B.n424 VSUBS 0.007623f
C507 B.n425 VSUBS 0.007623f
C508 B.n426 VSUBS 0.007623f
C509 B.n427 VSUBS 0.007623f
C510 B.n428 VSUBS 0.007623f
C511 B.n429 VSUBS 0.007623f
C512 B.n430 VSUBS 0.007623f
C513 B.n431 VSUBS 0.007623f
C514 B.n432 VSUBS 0.007623f
C515 B.n433 VSUBS 0.007623f
C516 B.n434 VSUBS 0.007623f
C517 B.n435 VSUBS 0.007623f
C518 B.n436 VSUBS 0.007623f
C519 B.n437 VSUBS 0.007623f
C520 B.n438 VSUBS 0.007623f
C521 B.n439 VSUBS 0.007623f
C522 B.n440 VSUBS 0.007623f
C523 B.n441 VSUBS 0.007623f
C524 B.n442 VSUBS 0.007623f
C525 B.n443 VSUBS 0.007623f
C526 B.n444 VSUBS 0.007623f
C527 B.n445 VSUBS 0.007623f
C528 B.n446 VSUBS 0.007623f
C529 B.n447 VSUBS 0.007623f
C530 B.n448 VSUBS 0.007623f
C531 B.n449 VSUBS 0.007623f
C532 B.n450 VSUBS 0.007623f
C533 B.n451 VSUBS 0.007623f
C534 B.n452 VSUBS 0.007623f
C535 B.n453 VSUBS 0.007623f
C536 B.n454 VSUBS 0.007623f
C537 B.n455 VSUBS 0.007623f
C538 B.n456 VSUBS 0.007623f
C539 B.n457 VSUBS 0.007623f
C540 B.n458 VSUBS 0.007623f
C541 B.n459 VSUBS 0.007623f
C542 B.n460 VSUBS 0.007623f
C543 B.n461 VSUBS 0.007623f
C544 B.n462 VSUBS 0.007623f
C545 B.n463 VSUBS 0.007623f
C546 B.n464 VSUBS 0.007623f
C547 B.n465 VSUBS 0.007623f
C548 B.n466 VSUBS 0.007623f
C549 B.n467 VSUBS 0.007623f
C550 B.n468 VSUBS 0.007623f
C551 B.n469 VSUBS 0.007623f
C552 B.n470 VSUBS 0.007623f
C553 B.n471 VSUBS 0.007623f
C554 B.n472 VSUBS 0.007623f
C555 B.n473 VSUBS 0.007623f
C556 B.n474 VSUBS 0.007623f
C557 B.n475 VSUBS 0.007623f
C558 B.n476 VSUBS 0.007623f
C559 B.n477 VSUBS 0.007623f
C560 B.n478 VSUBS 0.007623f
C561 B.n479 VSUBS 0.007623f
C562 B.n480 VSUBS 0.007623f
C563 B.n481 VSUBS 0.007623f
C564 B.n482 VSUBS 0.007623f
C565 B.n483 VSUBS 0.007623f
C566 B.n484 VSUBS 0.007623f
C567 B.n485 VSUBS 0.007623f
C568 B.n486 VSUBS 0.007623f
C569 B.n487 VSUBS 0.007623f
C570 B.n488 VSUBS 0.007623f
C571 B.n489 VSUBS 0.007623f
C572 B.n490 VSUBS 0.007623f
C573 B.n491 VSUBS 0.007623f
C574 B.n492 VSUBS 0.007623f
C575 B.n493 VSUBS 0.018085f
C576 B.n494 VSUBS 0.019136f
C577 B.n495 VSUBS 0.019136f
C578 B.n496 VSUBS 0.007623f
C579 B.n497 VSUBS 0.007623f
C580 B.n498 VSUBS 0.007623f
C581 B.n499 VSUBS 0.007623f
C582 B.n500 VSUBS 0.007623f
C583 B.n501 VSUBS 0.007623f
C584 B.n502 VSUBS 0.007623f
C585 B.n503 VSUBS 0.007623f
C586 B.n504 VSUBS 0.007623f
C587 B.n505 VSUBS 0.007623f
C588 B.n506 VSUBS 0.007623f
C589 B.n507 VSUBS 0.007623f
C590 B.n508 VSUBS 0.007623f
C591 B.n509 VSUBS 0.007623f
C592 B.n510 VSUBS 0.007623f
C593 B.n511 VSUBS 0.007623f
C594 B.n512 VSUBS 0.007623f
C595 B.n513 VSUBS 0.007623f
C596 B.n514 VSUBS 0.007623f
C597 B.n515 VSUBS 0.007623f
C598 B.n516 VSUBS 0.007623f
C599 B.n517 VSUBS 0.007623f
C600 B.n518 VSUBS 0.007623f
C601 B.n519 VSUBS 0.007623f
C602 B.n520 VSUBS 0.007623f
C603 B.n521 VSUBS 0.007623f
C604 B.n522 VSUBS 0.007623f
C605 B.n523 VSUBS 0.007623f
C606 B.n524 VSUBS 0.007623f
C607 B.n525 VSUBS 0.007623f
C608 B.n526 VSUBS 0.007623f
C609 B.n527 VSUBS 0.007623f
C610 B.n528 VSUBS 0.007623f
C611 B.n529 VSUBS 0.007623f
C612 B.n530 VSUBS 0.007623f
C613 B.n531 VSUBS 0.007623f
C614 B.n532 VSUBS 0.007623f
C615 B.n533 VSUBS 0.007623f
C616 B.n534 VSUBS 0.007623f
C617 B.n535 VSUBS 0.007623f
C618 B.n536 VSUBS 0.007623f
C619 B.n537 VSUBS 0.007623f
C620 B.n538 VSUBS 0.007623f
C621 B.n539 VSUBS 0.007623f
C622 B.n540 VSUBS 0.007623f
C623 B.n541 VSUBS 0.007623f
C624 B.n542 VSUBS 0.007623f
C625 B.n543 VSUBS 0.007623f
C626 B.n544 VSUBS 0.007623f
C627 B.n545 VSUBS 0.007623f
C628 B.n546 VSUBS 0.007623f
C629 B.n547 VSUBS 0.007623f
C630 B.n548 VSUBS 0.007623f
C631 B.n549 VSUBS 0.007623f
C632 B.n550 VSUBS 0.007623f
C633 B.n551 VSUBS 0.007623f
C634 B.n552 VSUBS 0.007623f
C635 B.n553 VSUBS 0.007623f
C636 B.n554 VSUBS 0.007623f
C637 B.n555 VSUBS 0.007623f
C638 B.n556 VSUBS 0.007623f
C639 B.n557 VSUBS 0.007623f
C640 B.n558 VSUBS 0.007623f
C641 B.n559 VSUBS 0.007623f
C642 B.n560 VSUBS 0.007623f
C643 B.n561 VSUBS 0.007623f
C644 B.n562 VSUBS 0.007623f
C645 B.n563 VSUBS 0.007623f
C646 B.n564 VSUBS 0.007623f
C647 B.n565 VSUBS 0.007623f
C648 B.n566 VSUBS 0.007623f
C649 B.n567 VSUBS 0.007623f
C650 B.n568 VSUBS 0.007623f
C651 B.n569 VSUBS 0.007623f
C652 B.n570 VSUBS 0.007623f
C653 B.n571 VSUBS 0.007623f
C654 B.n572 VSUBS 0.007623f
C655 B.n573 VSUBS 0.007623f
C656 B.n574 VSUBS 0.007623f
C657 B.n575 VSUBS 0.007623f
C658 B.n576 VSUBS 0.007623f
C659 B.n577 VSUBS 0.007623f
C660 B.n578 VSUBS 0.007623f
C661 B.n579 VSUBS 0.007623f
C662 B.n580 VSUBS 0.007623f
C663 B.n581 VSUBS 0.007623f
C664 B.n582 VSUBS 0.007623f
C665 B.n583 VSUBS 0.007623f
C666 B.n584 VSUBS 0.007623f
C667 B.n585 VSUBS 0.007175f
C668 B.n586 VSUBS 0.017663f
C669 B.n587 VSUBS 0.00426f
C670 B.n588 VSUBS 0.007623f
C671 B.n589 VSUBS 0.007623f
C672 B.n590 VSUBS 0.007623f
C673 B.n591 VSUBS 0.007623f
C674 B.n592 VSUBS 0.007623f
C675 B.n593 VSUBS 0.007623f
C676 B.n594 VSUBS 0.007623f
C677 B.n595 VSUBS 0.007623f
C678 B.n596 VSUBS 0.007623f
C679 B.n597 VSUBS 0.007623f
C680 B.n598 VSUBS 0.007623f
C681 B.n599 VSUBS 0.007623f
C682 B.n600 VSUBS 0.00426f
C683 B.n601 VSUBS 0.007623f
C684 B.n602 VSUBS 0.007623f
C685 B.n603 VSUBS 0.007175f
C686 B.n604 VSUBS 0.007623f
C687 B.n605 VSUBS 0.007623f
C688 B.n606 VSUBS 0.007623f
C689 B.n607 VSUBS 0.007623f
C690 B.n608 VSUBS 0.007623f
C691 B.n609 VSUBS 0.007623f
C692 B.n610 VSUBS 0.007623f
C693 B.n611 VSUBS 0.007623f
C694 B.n612 VSUBS 0.007623f
C695 B.n613 VSUBS 0.007623f
C696 B.n614 VSUBS 0.007623f
C697 B.n615 VSUBS 0.007623f
C698 B.n616 VSUBS 0.007623f
C699 B.n617 VSUBS 0.007623f
C700 B.n618 VSUBS 0.007623f
C701 B.n619 VSUBS 0.007623f
C702 B.n620 VSUBS 0.007623f
C703 B.n621 VSUBS 0.007623f
C704 B.n622 VSUBS 0.007623f
C705 B.n623 VSUBS 0.007623f
C706 B.n624 VSUBS 0.007623f
C707 B.n625 VSUBS 0.007623f
C708 B.n626 VSUBS 0.007623f
C709 B.n627 VSUBS 0.007623f
C710 B.n628 VSUBS 0.007623f
C711 B.n629 VSUBS 0.007623f
C712 B.n630 VSUBS 0.007623f
C713 B.n631 VSUBS 0.007623f
C714 B.n632 VSUBS 0.007623f
C715 B.n633 VSUBS 0.007623f
C716 B.n634 VSUBS 0.007623f
C717 B.n635 VSUBS 0.007623f
C718 B.n636 VSUBS 0.007623f
C719 B.n637 VSUBS 0.007623f
C720 B.n638 VSUBS 0.007623f
C721 B.n639 VSUBS 0.007623f
C722 B.n640 VSUBS 0.007623f
C723 B.n641 VSUBS 0.007623f
C724 B.n642 VSUBS 0.007623f
C725 B.n643 VSUBS 0.007623f
C726 B.n644 VSUBS 0.007623f
C727 B.n645 VSUBS 0.007623f
C728 B.n646 VSUBS 0.007623f
C729 B.n647 VSUBS 0.007623f
C730 B.n648 VSUBS 0.007623f
C731 B.n649 VSUBS 0.007623f
C732 B.n650 VSUBS 0.007623f
C733 B.n651 VSUBS 0.007623f
C734 B.n652 VSUBS 0.007623f
C735 B.n653 VSUBS 0.007623f
C736 B.n654 VSUBS 0.007623f
C737 B.n655 VSUBS 0.007623f
C738 B.n656 VSUBS 0.007623f
C739 B.n657 VSUBS 0.007623f
C740 B.n658 VSUBS 0.007623f
C741 B.n659 VSUBS 0.007623f
C742 B.n660 VSUBS 0.007623f
C743 B.n661 VSUBS 0.007623f
C744 B.n662 VSUBS 0.007623f
C745 B.n663 VSUBS 0.007623f
C746 B.n664 VSUBS 0.007623f
C747 B.n665 VSUBS 0.007623f
C748 B.n666 VSUBS 0.007623f
C749 B.n667 VSUBS 0.007623f
C750 B.n668 VSUBS 0.007623f
C751 B.n669 VSUBS 0.007623f
C752 B.n670 VSUBS 0.007623f
C753 B.n671 VSUBS 0.007623f
C754 B.n672 VSUBS 0.007623f
C755 B.n673 VSUBS 0.007623f
C756 B.n674 VSUBS 0.007623f
C757 B.n675 VSUBS 0.007623f
C758 B.n676 VSUBS 0.007623f
C759 B.n677 VSUBS 0.007623f
C760 B.n678 VSUBS 0.007623f
C761 B.n679 VSUBS 0.007623f
C762 B.n680 VSUBS 0.007623f
C763 B.n681 VSUBS 0.007623f
C764 B.n682 VSUBS 0.007623f
C765 B.n683 VSUBS 0.007623f
C766 B.n684 VSUBS 0.007623f
C767 B.n685 VSUBS 0.007623f
C768 B.n686 VSUBS 0.007623f
C769 B.n687 VSUBS 0.007623f
C770 B.n688 VSUBS 0.007623f
C771 B.n689 VSUBS 0.007623f
C772 B.n690 VSUBS 0.007623f
C773 B.n691 VSUBS 0.007623f
C774 B.n692 VSUBS 0.019136f
C775 B.n693 VSUBS 0.019136f
C776 B.n694 VSUBS 0.018085f
C777 B.n695 VSUBS 0.007623f
C778 B.n696 VSUBS 0.007623f
C779 B.n697 VSUBS 0.007623f
C780 B.n698 VSUBS 0.007623f
C781 B.n699 VSUBS 0.007623f
C782 B.n700 VSUBS 0.007623f
C783 B.n701 VSUBS 0.007623f
C784 B.n702 VSUBS 0.007623f
C785 B.n703 VSUBS 0.007623f
C786 B.n704 VSUBS 0.007623f
C787 B.n705 VSUBS 0.007623f
C788 B.n706 VSUBS 0.007623f
C789 B.n707 VSUBS 0.007623f
C790 B.n708 VSUBS 0.007623f
C791 B.n709 VSUBS 0.007623f
C792 B.n710 VSUBS 0.007623f
C793 B.n711 VSUBS 0.007623f
C794 B.n712 VSUBS 0.007623f
C795 B.n713 VSUBS 0.007623f
C796 B.n714 VSUBS 0.007623f
C797 B.n715 VSUBS 0.007623f
C798 B.n716 VSUBS 0.007623f
C799 B.n717 VSUBS 0.007623f
C800 B.n718 VSUBS 0.007623f
C801 B.n719 VSUBS 0.007623f
C802 B.n720 VSUBS 0.007623f
C803 B.n721 VSUBS 0.007623f
C804 B.n722 VSUBS 0.007623f
C805 B.n723 VSUBS 0.007623f
C806 B.n724 VSUBS 0.007623f
C807 B.n725 VSUBS 0.007623f
C808 B.n726 VSUBS 0.007623f
C809 B.n727 VSUBS 0.009948f
C810 B.n728 VSUBS 0.010597f
C811 B.n729 VSUBS 0.021074f
C812 VTAIL.t6 VSUBS 0.354857f
C813 VTAIL.t4 VSUBS 0.354857f
C814 VTAIL.n0 VSUBS 2.81951f
C815 VTAIL.n1 VSUBS 0.660849f
C816 VTAIL.t3 VSUBS 3.67854f
C817 VTAIL.n2 VSUBS 0.801512f
C818 VTAIL.t11 VSUBS 3.67854f
C819 VTAIL.n3 VSUBS 0.801512f
C820 VTAIL.t13 VSUBS 0.354857f
C821 VTAIL.t12 VSUBS 0.354857f
C822 VTAIL.n4 VSUBS 2.81951f
C823 VTAIL.n5 VSUBS 0.72716f
C824 VTAIL.t14 VSUBS 3.67854f
C825 VTAIL.n6 VSUBS 2.41002f
C826 VTAIL.t0 VSUBS 3.67857f
C827 VTAIL.n7 VSUBS 2.40999f
C828 VTAIL.t7 VSUBS 0.354857f
C829 VTAIL.t1 VSUBS 0.354857f
C830 VTAIL.n8 VSUBS 2.81952f
C831 VTAIL.n9 VSUBS 0.727154f
C832 VTAIL.t2 VSUBS 3.67857f
C833 VTAIL.n10 VSUBS 0.801486f
C834 VTAIL.t15 VSUBS 3.67857f
C835 VTAIL.n11 VSUBS 0.801486f
C836 VTAIL.t9 VSUBS 0.354857f
C837 VTAIL.t10 VSUBS 0.354857f
C838 VTAIL.n12 VSUBS 2.81952f
C839 VTAIL.n13 VSUBS 0.727154f
C840 VTAIL.t8 VSUBS 3.67854f
C841 VTAIL.n14 VSUBS 2.41002f
C842 VTAIL.t5 VSUBS 3.67854f
C843 VTAIL.n15 VSUBS 2.40551f
C844 VDD1.t1 VSUBS 0.403057f
C845 VDD1.t5 VSUBS 0.403057f
C846 VDD1.n0 VSUBS 3.37374f
C847 VDD1.t0 VSUBS 0.403057f
C848 VDD1.t3 VSUBS 0.403057f
C849 VDD1.n1 VSUBS 3.37261f
C850 VDD1.t2 VSUBS 0.403057f
C851 VDD1.t7 VSUBS 0.403057f
C852 VDD1.n2 VSUBS 3.37261f
C853 VDD1.n3 VSUBS 3.52333f
C854 VDD1.t6 VSUBS 0.403057f
C855 VDD1.t4 VSUBS 0.403057f
C856 VDD1.n4 VSUBS 3.3688f
C857 VDD1.n5 VSUBS 3.41632f
C858 VP.n0 VSUBS 0.05082f
C859 VP.n1 VSUBS 0.011532f
C860 VP.n2 VSUBS 0.05082f
C861 VP.n3 VSUBS 0.05082f
C862 VP.t7 VSUBS 1.96326f
C863 VP.t5 VSUBS 1.96326f
C864 VP.n4 VSUBS 0.05082f
C865 VP.t6 VSUBS 1.96326f
C866 VP.n5 VSUBS 0.742071f
C867 VP.t0 VSUBS 1.98802f
C868 VP.n6 VSUBS 0.717128f
C869 VP.n7 VSUBS 0.215061f
C870 VP.n8 VSUBS 0.011532f
C871 VP.n9 VSUBS 0.736387f
C872 VP.n10 VSUBS 0.011532f
C873 VP.n11 VSUBS 0.734977f
C874 VP.n12 VSUBS 2.53254f
C875 VP.n13 VSUBS 2.57122f
C876 VP.t1 VSUBS 1.96326f
C877 VP.n14 VSUBS 0.734977f
C878 VP.n15 VSUBS 0.011532f
C879 VP.t2 VSUBS 1.96326f
C880 VP.n16 VSUBS 0.736387f
C881 VP.n17 VSUBS 0.05082f
C882 VP.n18 VSUBS 0.05082f
C883 VP.n19 VSUBS 0.05082f
C884 VP.t3 VSUBS 1.96326f
C885 VP.n20 VSUBS 0.736387f
C886 VP.n21 VSUBS 0.011532f
C887 VP.t4 VSUBS 1.96326f
C888 VP.n22 VSUBS 0.734977f
C889 VP.n23 VSUBS 0.039384f
.ends

