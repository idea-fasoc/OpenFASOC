* NGSPICE file created from diff_pair_sample_0496.ext - technology: sky130A

.subckt diff_pair_sample_0496 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VP.t0 VDD1.t3 B.t7 sky130_fd_pr__nfet_01v8 ad=2.3133 pd=14.35 as=2.3133 ps=14.35 w=14.02 l=1.5
X1 B.t21 B.t19 B.t20 B.t13 sky130_fd_pr__nfet_01v8 ad=5.4678 pd=28.82 as=0 ps=0 w=14.02 l=1.5
X2 VTAIL.t3 VN.t0 VDD2.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=5.4678 pd=28.82 as=2.3133 ps=14.35 w=14.02 l=1.5
X3 VDD2.t6 VN.t1 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=2.3133 pd=14.35 as=2.3133 ps=14.35 w=14.02 l=1.5
X4 VTAIL.t1 VN.t2 VDD2.t5 B.t1 sky130_fd_pr__nfet_01v8 ad=5.4678 pd=28.82 as=2.3133 ps=14.35 w=14.02 l=1.5
X5 VDD1.t4 VP.t1 VTAIL.t14 B.t0 sky130_fd_pr__nfet_01v8 ad=2.3133 pd=14.35 as=5.4678 ps=28.82 w=14.02 l=1.5
X6 VTAIL.t7 VN.t3 VDD2.t4 B.t7 sky130_fd_pr__nfet_01v8 ad=2.3133 pd=14.35 as=2.3133 ps=14.35 w=14.02 l=1.5
X7 VDD1.t2 VP.t2 VTAIL.t13 B.t5 sky130_fd_pr__nfet_01v8 ad=2.3133 pd=14.35 as=2.3133 ps=14.35 w=14.02 l=1.5
X8 B.t18 B.t16 B.t17 B.t9 sky130_fd_pr__nfet_01v8 ad=5.4678 pd=28.82 as=0 ps=0 w=14.02 l=1.5
X9 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=5.4678 pd=28.82 as=0 ps=0 w=14.02 l=1.5
X10 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=5.4678 pd=28.82 as=0 ps=0 w=14.02 l=1.5
X11 VDD1.t6 VP.t3 VTAIL.t12 B.t4 sky130_fd_pr__nfet_01v8 ad=2.3133 pd=14.35 as=2.3133 ps=14.35 w=14.02 l=1.5
X12 VTAIL.t2 VN.t4 VDD2.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=2.3133 pd=14.35 as=2.3133 ps=14.35 w=14.02 l=1.5
X13 VTAIL.t11 VP.t4 VDD1.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=5.4678 pd=28.82 as=2.3133 ps=14.35 w=14.02 l=1.5
X14 VTAIL.t10 VP.t5 VDD1.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=5.4678 pd=28.82 as=2.3133 ps=14.35 w=14.02 l=1.5
X15 VDD2.t2 VN.t5 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.3133 pd=14.35 as=5.4678 ps=28.82 w=14.02 l=1.5
X16 VDD2.t1 VN.t6 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=2.3133 pd=14.35 as=2.3133 ps=14.35 w=14.02 l=1.5
X17 VTAIL.t9 VP.t6 VDD1.t5 B.t2 sky130_fd_pr__nfet_01v8 ad=2.3133 pd=14.35 as=2.3133 ps=14.35 w=14.02 l=1.5
X18 VDD1.t0 VP.t7 VTAIL.t8 B.t6 sky130_fd_pr__nfet_01v8 ad=2.3133 pd=14.35 as=5.4678 ps=28.82 w=14.02 l=1.5
X19 VDD2.t0 VN.t7 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=2.3133 pd=14.35 as=5.4678 ps=28.82 w=14.02 l=1.5
R0 VP.n11 VP.t5 260.092
R1 VP.n25 VP.t4 225.256
R2 VP.n31 VP.t2 225.256
R3 VP.n38 VP.t6 225.256
R4 VP.n45 VP.t1 225.256
R5 VP.n23 VP.t7 225.256
R6 VP.n16 VP.t0 225.256
R7 VP.n10 VP.t3 225.256
R8 VP.n26 VP.n25 173.843
R9 VP.n46 VP.n45 173.843
R10 VP.n24 VP.n23 173.843
R11 VP.n12 VP.n9 161.3
R12 VP.n14 VP.n13 161.3
R13 VP.n15 VP.n8 161.3
R14 VP.n18 VP.n17 161.3
R15 VP.n19 VP.n7 161.3
R16 VP.n21 VP.n20 161.3
R17 VP.n22 VP.n6 161.3
R18 VP.n44 VP.n0 161.3
R19 VP.n43 VP.n42 161.3
R20 VP.n41 VP.n1 161.3
R21 VP.n40 VP.n39 161.3
R22 VP.n37 VP.n2 161.3
R23 VP.n36 VP.n35 161.3
R24 VP.n34 VP.n3 161.3
R25 VP.n33 VP.n32 161.3
R26 VP.n30 VP.n4 161.3
R27 VP.n29 VP.n28 161.3
R28 VP.n27 VP.n5 161.3
R29 VP.n30 VP.n29 56.5617
R30 VP.n43 VP.n1 56.5617
R31 VP.n21 VP.n7 56.5617
R32 VP.n26 VP.n24 47.2354
R33 VP.n11 VP.n10 46.3697
R34 VP.n36 VP.n3 40.577
R35 VP.n37 VP.n36 40.577
R36 VP.n15 VP.n14 40.577
R37 VP.n14 VP.n9 40.577
R38 VP.n29 VP.n5 24.5923
R39 VP.n32 VP.n30 24.5923
R40 VP.n39 VP.n1 24.5923
R41 VP.n44 VP.n43 24.5923
R42 VP.n22 VP.n21 24.5923
R43 VP.n17 VP.n7 24.5923
R44 VP.n31 VP.n3 20.4117
R45 VP.n38 VP.n37 20.4117
R46 VP.n16 VP.n15 20.4117
R47 VP.n10 VP.n9 20.4117
R48 VP.n12 VP.n11 17.5628
R49 VP.n25 VP.n5 12.0505
R50 VP.n45 VP.n44 12.0505
R51 VP.n23 VP.n22 12.0505
R52 VP.n32 VP.n31 4.18111
R53 VP.n39 VP.n38 4.18111
R54 VP.n17 VP.n16 4.18111
R55 VP.n13 VP.n12 0.189894
R56 VP.n13 VP.n8 0.189894
R57 VP.n18 VP.n8 0.189894
R58 VP.n19 VP.n18 0.189894
R59 VP.n20 VP.n19 0.189894
R60 VP.n20 VP.n6 0.189894
R61 VP.n24 VP.n6 0.189894
R62 VP.n27 VP.n26 0.189894
R63 VP.n28 VP.n27 0.189894
R64 VP.n28 VP.n4 0.189894
R65 VP.n33 VP.n4 0.189894
R66 VP.n34 VP.n33 0.189894
R67 VP.n35 VP.n34 0.189894
R68 VP.n35 VP.n2 0.189894
R69 VP.n40 VP.n2 0.189894
R70 VP.n41 VP.n40 0.189894
R71 VP.n42 VP.n41 0.189894
R72 VP.n42 VP.n0 0.189894
R73 VP.n46 VP.n0 0.189894
R74 VP VP.n46 0.0516364
R75 VDD1 VDD1.n0 63.8008
R76 VDD1.n3 VDD1.n2 63.6871
R77 VDD1.n3 VDD1.n1 63.6871
R78 VDD1.n5 VDD1.n4 62.9536
R79 VDD1.n5 VDD1.n3 43.4836
R80 VDD1.n4 VDD1.t3 1.41277
R81 VDD1.n4 VDD1.t0 1.41277
R82 VDD1.n0 VDD1.t1 1.41277
R83 VDD1.n0 VDD1.t6 1.41277
R84 VDD1.n2 VDD1.t5 1.41277
R85 VDD1.n2 VDD1.t4 1.41277
R86 VDD1.n1 VDD1.t7 1.41277
R87 VDD1.n1 VDD1.t2 1.41277
R88 VDD1 VDD1.n5 0.731103
R89 VTAIL.n626 VTAIL.n554 289.615
R90 VTAIL.n74 VTAIL.n2 289.615
R91 VTAIL.n152 VTAIL.n80 289.615
R92 VTAIL.n232 VTAIL.n160 289.615
R93 VTAIL.n548 VTAIL.n476 289.615
R94 VTAIL.n468 VTAIL.n396 289.615
R95 VTAIL.n390 VTAIL.n318 289.615
R96 VTAIL.n310 VTAIL.n238 289.615
R97 VTAIL.n578 VTAIL.n577 185
R98 VTAIL.n583 VTAIL.n582 185
R99 VTAIL.n585 VTAIL.n584 185
R100 VTAIL.n574 VTAIL.n573 185
R101 VTAIL.n591 VTAIL.n590 185
R102 VTAIL.n593 VTAIL.n592 185
R103 VTAIL.n570 VTAIL.n569 185
R104 VTAIL.n599 VTAIL.n598 185
R105 VTAIL.n601 VTAIL.n600 185
R106 VTAIL.n566 VTAIL.n565 185
R107 VTAIL.n607 VTAIL.n606 185
R108 VTAIL.n609 VTAIL.n608 185
R109 VTAIL.n562 VTAIL.n561 185
R110 VTAIL.n615 VTAIL.n614 185
R111 VTAIL.n617 VTAIL.n616 185
R112 VTAIL.n558 VTAIL.n557 185
R113 VTAIL.n624 VTAIL.n623 185
R114 VTAIL.n625 VTAIL.n556 185
R115 VTAIL.n627 VTAIL.n626 185
R116 VTAIL.n26 VTAIL.n25 185
R117 VTAIL.n31 VTAIL.n30 185
R118 VTAIL.n33 VTAIL.n32 185
R119 VTAIL.n22 VTAIL.n21 185
R120 VTAIL.n39 VTAIL.n38 185
R121 VTAIL.n41 VTAIL.n40 185
R122 VTAIL.n18 VTAIL.n17 185
R123 VTAIL.n47 VTAIL.n46 185
R124 VTAIL.n49 VTAIL.n48 185
R125 VTAIL.n14 VTAIL.n13 185
R126 VTAIL.n55 VTAIL.n54 185
R127 VTAIL.n57 VTAIL.n56 185
R128 VTAIL.n10 VTAIL.n9 185
R129 VTAIL.n63 VTAIL.n62 185
R130 VTAIL.n65 VTAIL.n64 185
R131 VTAIL.n6 VTAIL.n5 185
R132 VTAIL.n72 VTAIL.n71 185
R133 VTAIL.n73 VTAIL.n4 185
R134 VTAIL.n75 VTAIL.n74 185
R135 VTAIL.n104 VTAIL.n103 185
R136 VTAIL.n109 VTAIL.n108 185
R137 VTAIL.n111 VTAIL.n110 185
R138 VTAIL.n100 VTAIL.n99 185
R139 VTAIL.n117 VTAIL.n116 185
R140 VTAIL.n119 VTAIL.n118 185
R141 VTAIL.n96 VTAIL.n95 185
R142 VTAIL.n125 VTAIL.n124 185
R143 VTAIL.n127 VTAIL.n126 185
R144 VTAIL.n92 VTAIL.n91 185
R145 VTAIL.n133 VTAIL.n132 185
R146 VTAIL.n135 VTAIL.n134 185
R147 VTAIL.n88 VTAIL.n87 185
R148 VTAIL.n141 VTAIL.n140 185
R149 VTAIL.n143 VTAIL.n142 185
R150 VTAIL.n84 VTAIL.n83 185
R151 VTAIL.n150 VTAIL.n149 185
R152 VTAIL.n151 VTAIL.n82 185
R153 VTAIL.n153 VTAIL.n152 185
R154 VTAIL.n184 VTAIL.n183 185
R155 VTAIL.n189 VTAIL.n188 185
R156 VTAIL.n191 VTAIL.n190 185
R157 VTAIL.n180 VTAIL.n179 185
R158 VTAIL.n197 VTAIL.n196 185
R159 VTAIL.n199 VTAIL.n198 185
R160 VTAIL.n176 VTAIL.n175 185
R161 VTAIL.n205 VTAIL.n204 185
R162 VTAIL.n207 VTAIL.n206 185
R163 VTAIL.n172 VTAIL.n171 185
R164 VTAIL.n213 VTAIL.n212 185
R165 VTAIL.n215 VTAIL.n214 185
R166 VTAIL.n168 VTAIL.n167 185
R167 VTAIL.n221 VTAIL.n220 185
R168 VTAIL.n223 VTAIL.n222 185
R169 VTAIL.n164 VTAIL.n163 185
R170 VTAIL.n230 VTAIL.n229 185
R171 VTAIL.n231 VTAIL.n162 185
R172 VTAIL.n233 VTAIL.n232 185
R173 VTAIL.n549 VTAIL.n548 185
R174 VTAIL.n547 VTAIL.n478 185
R175 VTAIL.n546 VTAIL.n545 185
R176 VTAIL.n481 VTAIL.n479 185
R177 VTAIL.n540 VTAIL.n539 185
R178 VTAIL.n538 VTAIL.n537 185
R179 VTAIL.n485 VTAIL.n484 185
R180 VTAIL.n532 VTAIL.n531 185
R181 VTAIL.n530 VTAIL.n529 185
R182 VTAIL.n489 VTAIL.n488 185
R183 VTAIL.n524 VTAIL.n523 185
R184 VTAIL.n522 VTAIL.n521 185
R185 VTAIL.n493 VTAIL.n492 185
R186 VTAIL.n516 VTAIL.n515 185
R187 VTAIL.n514 VTAIL.n513 185
R188 VTAIL.n497 VTAIL.n496 185
R189 VTAIL.n508 VTAIL.n507 185
R190 VTAIL.n506 VTAIL.n505 185
R191 VTAIL.n501 VTAIL.n500 185
R192 VTAIL.n469 VTAIL.n468 185
R193 VTAIL.n467 VTAIL.n398 185
R194 VTAIL.n466 VTAIL.n465 185
R195 VTAIL.n401 VTAIL.n399 185
R196 VTAIL.n460 VTAIL.n459 185
R197 VTAIL.n458 VTAIL.n457 185
R198 VTAIL.n405 VTAIL.n404 185
R199 VTAIL.n452 VTAIL.n451 185
R200 VTAIL.n450 VTAIL.n449 185
R201 VTAIL.n409 VTAIL.n408 185
R202 VTAIL.n444 VTAIL.n443 185
R203 VTAIL.n442 VTAIL.n441 185
R204 VTAIL.n413 VTAIL.n412 185
R205 VTAIL.n436 VTAIL.n435 185
R206 VTAIL.n434 VTAIL.n433 185
R207 VTAIL.n417 VTAIL.n416 185
R208 VTAIL.n428 VTAIL.n427 185
R209 VTAIL.n426 VTAIL.n425 185
R210 VTAIL.n421 VTAIL.n420 185
R211 VTAIL.n391 VTAIL.n390 185
R212 VTAIL.n389 VTAIL.n320 185
R213 VTAIL.n388 VTAIL.n387 185
R214 VTAIL.n323 VTAIL.n321 185
R215 VTAIL.n382 VTAIL.n381 185
R216 VTAIL.n380 VTAIL.n379 185
R217 VTAIL.n327 VTAIL.n326 185
R218 VTAIL.n374 VTAIL.n373 185
R219 VTAIL.n372 VTAIL.n371 185
R220 VTAIL.n331 VTAIL.n330 185
R221 VTAIL.n366 VTAIL.n365 185
R222 VTAIL.n364 VTAIL.n363 185
R223 VTAIL.n335 VTAIL.n334 185
R224 VTAIL.n358 VTAIL.n357 185
R225 VTAIL.n356 VTAIL.n355 185
R226 VTAIL.n339 VTAIL.n338 185
R227 VTAIL.n350 VTAIL.n349 185
R228 VTAIL.n348 VTAIL.n347 185
R229 VTAIL.n343 VTAIL.n342 185
R230 VTAIL.n311 VTAIL.n310 185
R231 VTAIL.n309 VTAIL.n240 185
R232 VTAIL.n308 VTAIL.n307 185
R233 VTAIL.n243 VTAIL.n241 185
R234 VTAIL.n302 VTAIL.n301 185
R235 VTAIL.n300 VTAIL.n299 185
R236 VTAIL.n247 VTAIL.n246 185
R237 VTAIL.n294 VTAIL.n293 185
R238 VTAIL.n292 VTAIL.n291 185
R239 VTAIL.n251 VTAIL.n250 185
R240 VTAIL.n286 VTAIL.n285 185
R241 VTAIL.n284 VTAIL.n283 185
R242 VTAIL.n255 VTAIL.n254 185
R243 VTAIL.n278 VTAIL.n277 185
R244 VTAIL.n276 VTAIL.n275 185
R245 VTAIL.n259 VTAIL.n258 185
R246 VTAIL.n270 VTAIL.n269 185
R247 VTAIL.n268 VTAIL.n267 185
R248 VTAIL.n263 VTAIL.n262 185
R249 VTAIL.n579 VTAIL.t6 147.659
R250 VTAIL.n27 VTAIL.t1 147.659
R251 VTAIL.n105 VTAIL.t14 147.659
R252 VTAIL.n185 VTAIL.t11 147.659
R253 VTAIL.n502 VTAIL.t8 147.659
R254 VTAIL.n422 VTAIL.t10 147.659
R255 VTAIL.n344 VTAIL.t0 147.659
R256 VTAIL.n264 VTAIL.t3 147.659
R257 VTAIL.n583 VTAIL.n577 104.615
R258 VTAIL.n584 VTAIL.n583 104.615
R259 VTAIL.n584 VTAIL.n573 104.615
R260 VTAIL.n591 VTAIL.n573 104.615
R261 VTAIL.n592 VTAIL.n591 104.615
R262 VTAIL.n592 VTAIL.n569 104.615
R263 VTAIL.n599 VTAIL.n569 104.615
R264 VTAIL.n600 VTAIL.n599 104.615
R265 VTAIL.n600 VTAIL.n565 104.615
R266 VTAIL.n607 VTAIL.n565 104.615
R267 VTAIL.n608 VTAIL.n607 104.615
R268 VTAIL.n608 VTAIL.n561 104.615
R269 VTAIL.n615 VTAIL.n561 104.615
R270 VTAIL.n616 VTAIL.n615 104.615
R271 VTAIL.n616 VTAIL.n557 104.615
R272 VTAIL.n624 VTAIL.n557 104.615
R273 VTAIL.n625 VTAIL.n624 104.615
R274 VTAIL.n626 VTAIL.n625 104.615
R275 VTAIL.n31 VTAIL.n25 104.615
R276 VTAIL.n32 VTAIL.n31 104.615
R277 VTAIL.n32 VTAIL.n21 104.615
R278 VTAIL.n39 VTAIL.n21 104.615
R279 VTAIL.n40 VTAIL.n39 104.615
R280 VTAIL.n40 VTAIL.n17 104.615
R281 VTAIL.n47 VTAIL.n17 104.615
R282 VTAIL.n48 VTAIL.n47 104.615
R283 VTAIL.n48 VTAIL.n13 104.615
R284 VTAIL.n55 VTAIL.n13 104.615
R285 VTAIL.n56 VTAIL.n55 104.615
R286 VTAIL.n56 VTAIL.n9 104.615
R287 VTAIL.n63 VTAIL.n9 104.615
R288 VTAIL.n64 VTAIL.n63 104.615
R289 VTAIL.n64 VTAIL.n5 104.615
R290 VTAIL.n72 VTAIL.n5 104.615
R291 VTAIL.n73 VTAIL.n72 104.615
R292 VTAIL.n74 VTAIL.n73 104.615
R293 VTAIL.n109 VTAIL.n103 104.615
R294 VTAIL.n110 VTAIL.n109 104.615
R295 VTAIL.n110 VTAIL.n99 104.615
R296 VTAIL.n117 VTAIL.n99 104.615
R297 VTAIL.n118 VTAIL.n117 104.615
R298 VTAIL.n118 VTAIL.n95 104.615
R299 VTAIL.n125 VTAIL.n95 104.615
R300 VTAIL.n126 VTAIL.n125 104.615
R301 VTAIL.n126 VTAIL.n91 104.615
R302 VTAIL.n133 VTAIL.n91 104.615
R303 VTAIL.n134 VTAIL.n133 104.615
R304 VTAIL.n134 VTAIL.n87 104.615
R305 VTAIL.n141 VTAIL.n87 104.615
R306 VTAIL.n142 VTAIL.n141 104.615
R307 VTAIL.n142 VTAIL.n83 104.615
R308 VTAIL.n150 VTAIL.n83 104.615
R309 VTAIL.n151 VTAIL.n150 104.615
R310 VTAIL.n152 VTAIL.n151 104.615
R311 VTAIL.n189 VTAIL.n183 104.615
R312 VTAIL.n190 VTAIL.n189 104.615
R313 VTAIL.n190 VTAIL.n179 104.615
R314 VTAIL.n197 VTAIL.n179 104.615
R315 VTAIL.n198 VTAIL.n197 104.615
R316 VTAIL.n198 VTAIL.n175 104.615
R317 VTAIL.n205 VTAIL.n175 104.615
R318 VTAIL.n206 VTAIL.n205 104.615
R319 VTAIL.n206 VTAIL.n171 104.615
R320 VTAIL.n213 VTAIL.n171 104.615
R321 VTAIL.n214 VTAIL.n213 104.615
R322 VTAIL.n214 VTAIL.n167 104.615
R323 VTAIL.n221 VTAIL.n167 104.615
R324 VTAIL.n222 VTAIL.n221 104.615
R325 VTAIL.n222 VTAIL.n163 104.615
R326 VTAIL.n230 VTAIL.n163 104.615
R327 VTAIL.n231 VTAIL.n230 104.615
R328 VTAIL.n232 VTAIL.n231 104.615
R329 VTAIL.n548 VTAIL.n547 104.615
R330 VTAIL.n547 VTAIL.n546 104.615
R331 VTAIL.n546 VTAIL.n479 104.615
R332 VTAIL.n539 VTAIL.n479 104.615
R333 VTAIL.n539 VTAIL.n538 104.615
R334 VTAIL.n538 VTAIL.n484 104.615
R335 VTAIL.n531 VTAIL.n484 104.615
R336 VTAIL.n531 VTAIL.n530 104.615
R337 VTAIL.n530 VTAIL.n488 104.615
R338 VTAIL.n523 VTAIL.n488 104.615
R339 VTAIL.n523 VTAIL.n522 104.615
R340 VTAIL.n522 VTAIL.n492 104.615
R341 VTAIL.n515 VTAIL.n492 104.615
R342 VTAIL.n515 VTAIL.n514 104.615
R343 VTAIL.n514 VTAIL.n496 104.615
R344 VTAIL.n507 VTAIL.n496 104.615
R345 VTAIL.n507 VTAIL.n506 104.615
R346 VTAIL.n506 VTAIL.n500 104.615
R347 VTAIL.n468 VTAIL.n467 104.615
R348 VTAIL.n467 VTAIL.n466 104.615
R349 VTAIL.n466 VTAIL.n399 104.615
R350 VTAIL.n459 VTAIL.n399 104.615
R351 VTAIL.n459 VTAIL.n458 104.615
R352 VTAIL.n458 VTAIL.n404 104.615
R353 VTAIL.n451 VTAIL.n404 104.615
R354 VTAIL.n451 VTAIL.n450 104.615
R355 VTAIL.n450 VTAIL.n408 104.615
R356 VTAIL.n443 VTAIL.n408 104.615
R357 VTAIL.n443 VTAIL.n442 104.615
R358 VTAIL.n442 VTAIL.n412 104.615
R359 VTAIL.n435 VTAIL.n412 104.615
R360 VTAIL.n435 VTAIL.n434 104.615
R361 VTAIL.n434 VTAIL.n416 104.615
R362 VTAIL.n427 VTAIL.n416 104.615
R363 VTAIL.n427 VTAIL.n426 104.615
R364 VTAIL.n426 VTAIL.n420 104.615
R365 VTAIL.n390 VTAIL.n389 104.615
R366 VTAIL.n389 VTAIL.n388 104.615
R367 VTAIL.n388 VTAIL.n321 104.615
R368 VTAIL.n381 VTAIL.n321 104.615
R369 VTAIL.n381 VTAIL.n380 104.615
R370 VTAIL.n380 VTAIL.n326 104.615
R371 VTAIL.n373 VTAIL.n326 104.615
R372 VTAIL.n373 VTAIL.n372 104.615
R373 VTAIL.n372 VTAIL.n330 104.615
R374 VTAIL.n365 VTAIL.n330 104.615
R375 VTAIL.n365 VTAIL.n364 104.615
R376 VTAIL.n364 VTAIL.n334 104.615
R377 VTAIL.n357 VTAIL.n334 104.615
R378 VTAIL.n357 VTAIL.n356 104.615
R379 VTAIL.n356 VTAIL.n338 104.615
R380 VTAIL.n349 VTAIL.n338 104.615
R381 VTAIL.n349 VTAIL.n348 104.615
R382 VTAIL.n348 VTAIL.n342 104.615
R383 VTAIL.n310 VTAIL.n309 104.615
R384 VTAIL.n309 VTAIL.n308 104.615
R385 VTAIL.n308 VTAIL.n241 104.615
R386 VTAIL.n301 VTAIL.n241 104.615
R387 VTAIL.n301 VTAIL.n300 104.615
R388 VTAIL.n300 VTAIL.n246 104.615
R389 VTAIL.n293 VTAIL.n246 104.615
R390 VTAIL.n293 VTAIL.n292 104.615
R391 VTAIL.n292 VTAIL.n250 104.615
R392 VTAIL.n285 VTAIL.n250 104.615
R393 VTAIL.n285 VTAIL.n284 104.615
R394 VTAIL.n284 VTAIL.n254 104.615
R395 VTAIL.n277 VTAIL.n254 104.615
R396 VTAIL.n277 VTAIL.n276 104.615
R397 VTAIL.n276 VTAIL.n258 104.615
R398 VTAIL.n269 VTAIL.n258 104.615
R399 VTAIL.n269 VTAIL.n268 104.615
R400 VTAIL.n268 VTAIL.n262 104.615
R401 VTAIL.t6 VTAIL.n577 52.3082
R402 VTAIL.t1 VTAIL.n25 52.3082
R403 VTAIL.t14 VTAIL.n103 52.3082
R404 VTAIL.t11 VTAIL.n183 52.3082
R405 VTAIL.t8 VTAIL.n500 52.3082
R406 VTAIL.t10 VTAIL.n420 52.3082
R407 VTAIL.t0 VTAIL.n342 52.3082
R408 VTAIL.t3 VTAIL.n262 52.3082
R409 VTAIL.n475 VTAIL.n474 46.275
R410 VTAIL.n317 VTAIL.n316 46.275
R411 VTAIL.n1 VTAIL.n0 46.2748
R412 VTAIL.n159 VTAIL.n158 46.2748
R413 VTAIL.n631 VTAIL.n630 34.1247
R414 VTAIL.n79 VTAIL.n78 34.1247
R415 VTAIL.n157 VTAIL.n156 34.1247
R416 VTAIL.n237 VTAIL.n236 34.1247
R417 VTAIL.n553 VTAIL.n552 34.1247
R418 VTAIL.n473 VTAIL.n472 34.1247
R419 VTAIL.n395 VTAIL.n394 34.1247
R420 VTAIL.n315 VTAIL.n314 34.1247
R421 VTAIL.n631 VTAIL.n553 26.0307
R422 VTAIL.n315 VTAIL.n237 26.0307
R423 VTAIL.n579 VTAIL.n578 15.6677
R424 VTAIL.n27 VTAIL.n26 15.6677
R425 VTAIL.n105 VTAIL.n104 15.6677
R426 VTAIL.n185 VTAIL.n184 15.6677
R427 VTAIL.n502 VTAIL.n501 15.6677
R428 VTAIL.n422 VTAIL.n421 15.6677
R429 VTAIL.n344 VTAIL.n343 15.6677
R430 VTAIL.n264 VTAIL.n263 15.6677
R431 VTAIL.n627 VTAIL.n556 13.1884
R432 VTAIL.n75 VTAIL.n4 13.1884
R433 VTAIL.n153 VTAIL.n82 13.1884
R434 VTAIL.n233 VTAIL.n162 13.1884
R435 VTAIL.n549 VTAIL.n478 13.1884
R436 VTAIL.n469 VTAIL.n398 13.1884
R437 VTAIL.n391 VTAIL.n320 13.1884
R438 VTAIL.n311 VTAIL.n240 13.1884
R439 VTAIL.n582 VTAIL.n581 12.8005
R440 VTAIL.n623 VTAIL.n622 12.8005
R441 VTAIL.n628 VTAIL.n554 12.8005
R442 VTAIL.n30 VTAIL.n29 12.8005
R443 VTAIL.n71 VTAIL.n70 12.8005
R444 VTAIL.n76 VTAIL.n2 12.8005
R445 VTAIL.n108 VTAIL.n107 12.8005
R446 VTAIL.n149 VTAIL.n148 12.8005
R447 VTAIL.n154 VTAIL.n80 12.8005
R448 VTAIL.n188 VTAIL.n187 12.8005
R449 VTAIL.n229 VTAIL.n228 12.8005
R450 VTAIL.n234 VTAIL.n160 12.8005
R451 VTAIL.n550 VTAIL.n476 12.8005
R452 VTAIL.n545 VTAIL.n480 12.8005
R453 VTAIL.n505 VTAIL.n504 12.8005
R454 VTAIL.n470 VTAIL.n396 12.8005
R455 VTAIL.n465 VTAIL.n400 12.8005
R456 VTAIL.n425 VTAIL.n424 12.8005
R457 VTAIL.n392 VTAIL.n318 12.8005
R458 VTAIL.n387 VTAIL.n322 12.8005
R459 VTAIL.n347 VTAIL.n346 12.8005
R460 VTAIL.n312 VTAIL.n238 12.8005
R461 VTAIL.n307 VTAIL.n242 12.8005
R462 VTAIL.n267 VTAIL.n266 12.8005
R463 VTAIL.n585 VTAIL.n576 12.0247
R464 VTAIL.n621 VTAIL.n558 12.0247
R465 VTAIL.n33 VTAIL.n24 12.0247
R466 VTAIL.n69 VTAIL.n6 12.0247
R467 VTAIL.n111 VTAIL.n102 12.0247
R468 VTAIL.n147 VTAIL.n84 12.0247
R469 VTAIL.n191 VTAIL.n182 12.0247
R470 VTAIL.n227 VTAIL.n164 12.0247
R471 VTAIL.n544 VTAIL.n481 12.0247
R472 VTAIL.n508 VTAIL.n499 12.0247
R473 VTAIL.n464 VTAIL.n401 12.0247
R474 VTAIL.n428 VTAIL.n419 12.0247
R475 VTAIL.n386 VTAIL.n323 12.0247
R476 VTAIL.n350 VTAIL.n341 12.0247
R477 VTAIL.n306 VTAIL.n243 12.0247
R478 VTAIL.n270 VTAIL.n261 12.0247
R479 VTAIL.n586 VTAIL.n574 11.249
R480 VTAIL.n618 VTAIL.n617 11.249
R481 VTAIL.n34 VTAIL.n22 11.249
R482 VTAIL.n66 VTAIL.n65 11.249
R483 VTAIL.n112 VTAIL.n100 11.249
R484 VTAIL.n144 VTAIL.n143 11.249
R485 VTAIL.n192 VTAIL.n180 11.249
R486 VTAIL.n224 VTAIL.n223 11.249
R487 VTAIL.n541 VTAIL.n540 11.249
R488 VTAIL.n509 VTAIL.n497 11.249
R489 VTAIL.n461 VTAIL.n460 11.249
R490 VTAIL.n429 VTAIL.n417 11.249
R491 VTAIL.n383 VTAIL.n382 11.249
R492 VTAIL.n351 VTAIL.n339 11.249
R493 VTAIL.n303 VTAIL.n302 11.249
R494 VTAIL.n271 VTAIL.n259 11.249
R495 VTAIL.n590 VTAIL.n589 10.4732
R496 VTAIL.n614 VTAIL.n560 10.4732
R497 VTAIL.n38 VTAIL.n37 10.4732
R498 VTAIL.n62 VTAIL.n8 10.4732
R499 VTAIL.n116 VTAIL.n115 10.4732
R500 VTAIL.n140 VTAIL.n86 10.4732
R501 VTAIL.n196 VTAIL.n195 10.4732
R502 VTAIL.n220 VTAIL.n166 10.4732
R503 VTAIL.n537 VTAIL.n483 10.4732
R504 VTAIL.n513 VTAIL.n512 10.4732
R505 VTAIL.n457 VTAIL.n403 10.4732
R506 VTAIL.n433 VTAIL.n432 10.4732
R507 VTAIL.n379 VTAIL.n325 10.4732
R508 VTAIL.n355 VTAIL.n354 10.4732
R509 VTAIL.n299 VTAIL.n245 10.4732
R510 VTAIL.n275 VTAIL.n274 10.4732
R511 VTAIL.n593 VTAIL.n572 9.69747
R512 VTAIL.n613 VTAIL.n562 9.69747
R513 VTAIL.n41 VTAIL.n20 9.69747
R514 VTAIL.n61 VTAIL.n10 9.69747
R515 VTAIL.n119 VTAIL.n98 9.69747
R516 VTAIL.n139 VTAIL.n88 9.69747
R517 VTAIL.n199 VTAIL.n178 9.69747
R518 VTAIL.n219 VTAIL.n168 9.69747
R519 VTAIL.n536 VTAIL.n485 9.69747
R520 VTAIL.n516 VTAIL.n495 9.69747
R521 VTAIL.n456 VTAIL.n405 9.69747
R522 VTAIL.n436 VTAIL.n415 9.69747
R523 VTAIL.n378 VTAIL.n327 9.69747
R524 VTAIL.n358 VTAIL.n337 9.69747
R525 VTAIL.n298 VTAIL.n247 9.69747
R526 VTAIL.n278 VTAIL.n257 9.69747
R527 VTAIL.n630 VTAIL.n629 9.45567
R528 VTAIL.n78 VTAIL.n77 9.45567
R529 VTAIL.n156 VTAIL.n155 9.45567
R530 VTAIL.n236 VTAIL.n235 9.45567
R531 VTAIL.n552 VTAIL.n551 9.45567
R532 VTAIL.n472 VTAIL.n471 9.45567
R533 VTAIL.n394 VTAIL.n393 9.45567
R534 VTAIL.n314 VTAIL.n313 9.45567
R535 VTAIL.n629 VTAIL.n628 9.3005
R536 VTAIL.n568 VTAIL.n567 9.3005
R537 VTAIL.n597 VTAIL.n596 9.3005
R538 VTAIL.n595 VTAIL.n594 9.3005
R539 VTAIL.n572 VTAIL.n571 9.3005
R540 VTAIL.n589 VTAIL.n588 9.3005
R541 VTAIL.n587 VTAIL.n586 9.3005
R542 VTAIL.n576 VTAIL.n575 9.3005
R543 VTAIL.n581 VTAIL.n580 9.3005
R544 VTAIL.n603 VTAIL.n602 9.3005
R545 VTAIL.n605 VTAIL.n604 9.3005
R546 VTAIL.n564 VTAIL.n563 9.3005
R547 VTAIL.n611 VTAIL.n610 9.3005
R548 VTAIL.n613 VTAIL.n612 9.3005
R549 VTAIL.n560 VTAIL.n559 9.3005
R550 VTAIL.n619 VTAIL.n618 9.3005
R551 VTAIL.n621 VTAIL.n620 9.3005
R552 VTAIL.n622 VTAIL.n555 9.3005
R553 VTAIL.n77 VTAIL.n76 9.3005
R554 VTAIL.n16 VTAIL.n15 9.3005
R555 VTAIL.n45 VTAIL.n44 9.3005
R556 VTAIL.n43 VTAIL.n42 9.3005
R557 VTAIL.n20 VTAIL.n19 9.3005
R558 VTAIL.n37 VTAIL.n36 9.3005
R559 VTAIL.n35 VTAIL.n34 9.3005
R560 VTAIL.n24 VTAIL.n23 9.3005
R561 VTAIL.n29 VTAIL.n28 9.3005
R562 VTAIL.n51 VTAIL.n50 9.3005
R563 VTAIL.n53 VTAIL.n52 9.3005
R564 VTAIL.n12 VTAIL.n11 9.3005
R565 VTAIL.n59 VTAIL.n58 9.3005
R566 VTAIL.n61 VTAIL.n60 9.3005
R567 VTAIL.n8 VTAIL.n7 9.3005
R568 VTAIL.n67 VTAIL.n66 9.3005
R569 VTAIL.n69 VTAIL.n68 9.3005
R570 VTAIL.n70 VTAIL.n3 9.3005
R571 VTAIL.n155 VTAIL.n154 9.3005
R572 VTAIL.n94 VTAIL.n93 9.3005
R573 VTAIL.n123 VTAIL.n122 9.3005
R574 VTAIL.n121 VTAIL.n120 9.3005
R575 VTAIL.n98 VTAIL.n97 9.3005
R576 VTAIL.n115 VTAIL.n114 9.3005
R577 VTAIL.n113 VTAIL.n112 9.3005
R578 VTAIL.n102 VTAIL.n101 9.3005
R579 VTAIL.n107 VTAIL.n106 9.3005
R580 VTAIL.n129 VTAIL.n128 9.3005
R581 VTAIL.n131 VTAIL.n130 9.3005
R582 VTAIL.n90 VTAIL.n89 9.3005
R583 VTAIL.n137 VTAIL.n136 9.3005
R584 VTAIL.n139 VTAIL.n138 9.3005
R585 VTAIL.n86 VTAIL.n85 9.3005
R586 VTAIL.n145 VTAIL.n144 9.3005
R587 VTAIL.n147 VTAIL.n146 9.3005
R588 VTAIL.n148 VTAIL.n81 9.3005
R589 VTAIL.n235 VTAIL.n234 9.3005
R590 VTAIL.n174 VTAIL.n173 9.3005
R591 VTAIL.n203 VTAIL.n202 9.3005
R592 VTAIL.n201 VTAIL.n200 9.3005
R593 VTAIL.n178 VTAIL.n177 9.3005
R594 VTAIL.n195 VTAIL.n194 9.3005
R595 VTAIL.n193 VTAIL.n192 9.3005
R596 VTAIL.n182 VTAIL.n181 9.3005
R597 VTAIL.n187 VTAIL.n186 9.3005
R598 VTAIL.n209 VTAIL.n208 9.3005
R599 VTAIL.n211 VTAIL.n210 9.3005
R600 VTAIL.n170 VTAIL.n169 9.3005
R601 VTAIL.n217 VTAIL.n216 9.3005
R602 VTAIL.n219 VTAIL.n218 9.3005
R603 VTAIL.n166 VTAIL.n165 9.3005
R604 VTAIL.n225 VTAIL.n224 9.3005
R605 VTAIL.n227 VTAIL.n226 9.3005
R606 VTAIL.n228 VTAIL.n161 9.3005
R607 VTAIL.n528 VTAIL.n527 9.3005
R608 VTAIL.n487 VTAIL.n486 9.3005
R609 VTAIL.n534 VTAIL.n533 9.3005
R610 VTAIL.n536 VTAIL.n535 9.3005
R611 VTAIL.n483 VTAIL.n482 9.3005
R612 VTAIL.n542 VTAIL.n541 9.3005
R613 VTAIL.n544 VTAIL.n543 9.3005
R614 VTAIL.n480 VTAIL.n477 9.3005
R615 VTAIL.n551 VTAIL.n550 9.3005
R616 VTAIL.n526 VTAIL.n525 9.3005
R617 VTAIL.n491 VTAIL.n490 9.3005
R618 VTAIL.n520 VTAIL.n519 9.3005
R619 VTAIL.n518 VTAIL.n517 9.3005
R620 VTAIL.n495 VTAIL.n494 9.3005
R621 VTAIL.n512 VTAIL.n511 9.3005
R622 VTAIL.n510 VTAIL.n509 9.3005
R623 VTAIL.n499 VTAIL.n498 9.3005
R624 VTAIL.n504 VTAIL.n503 9.3005
R625 VTAIL.n448 VTAIL.n447 9.3005
R626 VTAIL.n407 VTAIL.n406 9.3005
R627 VTAIL.n454 VTAIL.n453 9.3005
R628 VTAIL.n456 VTAIL.n455 9.3005
R629 VTAIL.n403 VTAIL.n402 9.3005
R630 VTAIL.n462 VTAIL.n461 9.3005
R631 VTAIL.n464 VTAIL.n463 9.3005
R632 VTAIL.n400 VTAIL.n397 9.3005
R633 VTAIL.n471 VTAIL.n470 9.3005
R634 VTAIL.n446 VTAIL.n445 9.3005
R635 VTAIL.n411 VTAIL.n410 9.3005
R636 VTAIL.n440 VTAIL.n439 9.3005
R637 VTAIL.n438 VTAIL.n437 9.3005
R638 VTAIL.n415 VTAIL.n414 9.3005
R639 VTAIL.n432 VTAIL.n431 9.3005
R640 VTAIL.n430 VTAIL.n429 9.3005
R641 VTAIL.n419 VTAIL.n418 9.3005
R642 VTAIL.n424 VTAIL.n423 9.3005
R643 VTAIL.n370 VTAIL.n369 9.3005
R644 VTAIL.n329 VTAIL.n328 9.3005
R645 VTAIL.n376 VTAIL.n375 9.3005
R646 VTAIL.n378 VTAIL.n377 9.3005
R647 VTAIL.n325 VTAIL.n324 9.3005
R648 VTAIL.n384 VTAIL.n383 9.3005
R649 VTAIL.n386 VTAIL.n385 9.3005
R650 VTAIL.n322 VTAIL.n319 9.3005
R651 VTAIL.n393 VTAIL.n392 9.3005
R652 VTAIL.n368 VTAIL.n367 9.3005
R653 VTAIL.n333 VTAIL.n332 9.3005
R654 VTAIL.n362 VTAIL.n361 9.3005
R655 VTAIL.n360 VTAIL.n359 9.3005
R656 VTAIL.n337 VTAIL.n336 9.3005
R657 VTAIL.n354 VTAIL.n353 9.3005
R658 VTAIL.n352 VTAIL.n351 9.3005
R659 VTAIL.n341 VTAIL.n340 9.3005
R660 VTAIL.n346 VTAIL.n345 9.3005
R661 VTAIL.n290 VTAIL.n289 9.3005
R662 VTAIL.n249 VTAIL.n248 9.3005
R663 VTAIL.n296 VTAIL.n295 9.3005
R664 VTAIL.n298 VTAIL.n297 9.3005
R665 VTAIL.n245 VTAIL.n244 9.3005
R666 VTAIL.n304 VTAIL.n303 9.3005
R667 VTAIL.n306 VTAIL.n305 9.3005
R668 VTAIL.n242 VTAIL.n239 9.3005
R669 VTAIL.n313 VTAIL.n312 9.3005
R670 VTAIL.n288 VTAIL.n287 9.3005
R671 VTAIL.n253 VTAIL.n252 9.3005
R672 VTAIL.n282 VTAIL.n281 9.3005
R673 VTAIL.n280 VTAIL.n279 9.3005
R674 VTAIL.n257 VTAIL.n256 9.3005
R675 VTAIL.n274 VTAIL.n273 9.3005
R676 VTAIL.n272 VTAIL.n271 9.3005
R677 VTAIL.n261 VTAIL.n260 9.3005
R678 VTAIL.n266 VTAIL.n265 9.3005
R679 VTAIL.n594 VTAIL.n570 8.92171
R680 VTAIL.n610 VTAIL.n609 8.92171
R681 VTAIL.n42 VTAIL.n18 8.92171
R682 VTAIL.n58 VTAIL.n57 8.92171
R683 VTAIL.n120 VTAIL.n96 8.92171
R684 VTAIL.n136 VTAIL.n135 8.92171
R685 VTAIL.n200 VTAIL.n176 8.92171
R686 VTAIL.n216 VTAIL.n215 8.92171
R687 VTAIL.n533 VTAIL.n532 8.92171
R688 VTAIL.n517 VTAIL.n493 8.92171
R689 VTAIL.n453 VTAIL.n452 8.92171
R690 VTAIL.n437 VTAIL.n413 8.92171
R691 VTAIL.n375 VTAIL.n374 8.92171
R692 VTAIL.n359 VTAIL.n335 8.92171
R693 VTAIL.n295 VTAIL.n294 8.92171
R694 VTAIL.n279 VTAIL.n255 8.92171
R695 VTAIL.n598 VTAIL.n597 8.14595
R696 VTAIL.n606 VTAIL.n564 8.14595
R697 VTAIL.n46 VTAIL.n45 8.14595
R698 VTAIL.n54 VTAIL.n12 8.14595
R699 VTAIL.n124 VTAIL.n123 8.14595
R700 VTAIL.n132 VTAIL.n90 8.14595
R701 VTAIL.n204 VTAIL.n203 8.14595
R702 VTAIL.n212 VTAIL.n170 8.14595
R703 VTAIL.n529 VTAIL.n487 8.14595
R704 VTAIL.n521 VTAIL.n520 8.14595
R705 VTAIL.n449 VTAIL.n407 8.14595
R706 VTAIL.n441 VTAIL.n440 8.14595
R707 VTAIL.n371 VTAIL.n329 8.14595
R708 VTAIL.n363 VTAIL.n362 8.14595
R709 VTAIL.n291 VTAIL.n249 8.14595
R710 VTAIL.n283 VTAIL.n282 8.14595
R711 VTAIL.n601 VTAIL.n568 7.3702
R712 VTAIL.n605 VTAIL.n566 7.3702
R713 VTAIL.n49 VTAIL.n16 7.3702
R714 VTAIL.n53 VTAIL.n14 7.3702
R715 VTAIL.n127 VTAIL.n94 7.3702
R716 VTAIL.n131 VTAIL.n92 7.3702
R717 VTAIL.n207 VTAIL.n174 7.3702
R718 VTAIL.n211 VTAIL.n172 7.3702
R719 VTAIL.n528 VTAIL.n489 7.3702
R720 VTAIL.n524 VTAIL.n491 7.3702
R721 VTAIL.n448 VTAIL.n409 7.3702
R722 VTAIL.n444 VTAIL.n411 7.3702
R723 VTAIL.n370 VTAIL.n331 7.3702
R724 VTAIL.n366 VTAIL.n333 7.3702
R725 VTAIL.n290 VTAIL.n251 7.3702
R726 VTAIL.n286 VTAIL.n253 7.3702
R727 VTAIL.n602 VTAIL.n601 6.59444
R728 VTAIL.n602 VTAIL.n566 6.59444
R729 VTAIL.n50 VTAIL.n49 6.59444
R730 VTAIL.n50 VTAIL.n14 6.59444
R731 VTAIL.n128 VTAIL.n127 6.59444
R732 VTAIL.n128 VTAIL.n92 6.59444
R733 VTAIL.n208 VTAIL.n207 6.59444
R734 VTAIL.n208 VTAIL.n172 6.59444
R735 VTAIL.n525 VTAIL.n489 6.59444
R736 VTAIL.n525 VTAIL.n524 6.59444
R737 VTAIL.n445 VTAIL.n409 6.59444
R738 VTAIL.n445 VTAIL.n444 6.59444
R739 VTAIL.n367 VTAIL.n331 6.59444
R740 VTAIL.n367 VTAIL.n366 6.59444
R741 VTAIL.n287 VTAIL.n251 6.59444
R742 VTAIL.n287 VTAIL.n286 6.59444
R743 VTAIL.n598 VTAIL.n568 5.81868
R744 VTAIL.n606 VTAIL.n605 5.81868
R745 VTAIL.n46 VTAIL.n16 5.81868
R746 VTAIL.n54 VTAIL.n53 5.81868
R747 VTAIL.n124 VTAIL.n94 5.81868
R748 VTAIL.n132 VTAIL.n131 5.81868
R749 VTAIL.n204 VTAIL.n174 5.81868
R750 VTAIL.n212 VTAIL.n211 5.81868
R751 VTAIL.n529 VTAIL.n528 5.81868
R752 VTAIL.n521 VTAIL.n491 5.81868
R753 VTAIL.n449 VTAIL.n448 5.81868
R754 VTAIL.n441 VTAIL.n411 5.81868
R755 VTAIL.n371 VTAIL.n370 5.81868
R756 VTAIL.n363 VTAIL.n333 5.81868
R757 VTAIL.n291 VTAIL.n290 5.81868
R758 VTAIL.n283 VTAIL.n253 5.81868
R759 VTAIL.n597 VTAIL.n570 5.04292
R760 VTAIL.n609 VTAIL.n564 5.04292
R761 VTAIL.n45 VTAIL.n18 5.04292
R762 VTAIL.n57 VTAIL.n12 5.04292
R763 VTAIL.n123 VTAIL.n96 5.04292
R764 VTAIL.n135 VTAIL.n90 5.04292
R765 VTAIL.n203 VTAIL.n176 5.04292
R766 VTAIL.n215 VTAIL.n170 5.04292
R767 VTAIL.n532 VTAIL.n487 5.04292
R768 VTAIL.n520 VTAIL.n493 5.04292
R769 VTAIL.n452 VTAIL.n407 5.04292
R770 VTAIL.n440 VTAIL.n413 5.04292
R771 VTAIL.n374 VTAIL.n329 5.04292
R772 VTAIL.n362 VTAIL.n335 5.04292
R773 VTAIL.n294 VTAIL.n249 5.04292
R774 VTAIL.n282 VTAIL.n255 5.04292
R775 VTAIL.n580 VTAIL.n579 4.38563
R776 VTAIL.n28 VTAIL.n27 4.38563
R777 VTAIL.n106 VTAIL.n105 4.38563
R778 VTAIL.n186 VTAIL.n185 4.38563
R779 VTAIL.n503 VTAIL.n502 4.38563
R780 VTAIL.n423 VTAIL.n422 4.38563
R781 VTAIL.n345 VTAIL.n344 4.38563
R782 VTAIL.n265 VTAIL.n264 4.38563
R783 VTAIL.n594 VTAIL.n593 4.26717
R784 VTAIL.n610 VTAIL.n562 4.26717
R785 VTAIL.n42 VTAIL.n41 4.26717
R786 VTAIL.n58 VTAIL.n10 4.26717
R787 VTAIL.n120 VTAIL.n119 4.26717
R788 VTAIL.n136 VTAIL.n88 4.26717
R789 VTAIL.n200 VTAIL.n199 4.26717
R790 VTAIL.n216 VTAIL.n168 4.26717
R791 VTAIL.n533 VTAIL.n485 4.26717
R792 VTAIL.n517 VTAIL.n516 4.26717
R793 VTAIL.n453 VTAIL.n405 4.26717
R794 VTAIL.n437 VTAIL.n436 4.26717
R795 VTAIL.n375 VTAIL.n327 4.26717
R796 VTAIL.n359 VTAIL.n358 4.26717
R797 VTAIL.n295 VTAIL.n247 4.26717
R798 VTAIL.n279 VTAIL.n278 4.26717
R799 VTAIL.n590 VTAIL.n572 3.49141
R800 VTAIL.n614 VTAIL.n613 3.49141
R801 VTAIL.n38 VTAIL.n20 3.49141
R802 VTAIL.n62 VTAIL.n61 3.49141
R803 VTAIL.n116 VTAIL.n98 3.49141
R804 VTAIL.n140 VTAIL.n139 3.49141
R805 VTAIL.n196 VTAIL.n178 3.49141
R806 VTAIL.n220 VTAIL.n219 3.49141
R807 VTAIL.n537 VTAIL.n536 3.49141
R808 VTAIL.n513 VTAIL.n495 3.49141
R809 VTAIL.n457 VTAIL.n456 3.49141
R810 VTAIL.n433 VTAIL.n415 3.49141
R811 VTAIL.n379 VTAIL.n378 3.49141
R812 VTAIL.n355 VTAIL.n337 3.49141
R813 VTAIL.n299 VTAIL.n298 3.49141
R814 VTAIL.n275 VTAIL.n257 3.49141
R815 VTAIL.n589 VTAIL.n574 2.71565
R816 VTAIL.n617 VTAIL.n560 2.71565
R817 VTAIL.n37 VTAIL.n22 2.71565
R818 VTAIL.n65 VTAIL.n8 2.71565
R819 VTAIL.n115 VTAIL.n100 2.71565
R820 VTAIL.n143 VTAIL.n86 2.71565
R821 VTAIL.n195 VTAIL.n180 2.71565
R822 VTAIL.n223 VTAIL.n166 2.71565
R823 VTAIL.n540 VTAIL.n483 2.71565
R824 VTAIL.n512 VTAIL.n497 2.71565
R825 VTAIL.n460 VTAIL.n403 2.71565
R826 VTAIL.n432 VTAIL.n417 2.71565
R827 VTAIL.n382 VTAIL.n325 2.71565
R828 VTAIL.n354 VTAIL.n339 2.71565
R829 VTAIL.n302 VTAIL.n245 2.71565
R830 VTAIL.n274 VTAIL.n259 2.71565
R831 VTAIL.n586 VTAIL.n585 1.93989
R832 VTAIL.n618 VTAIL.n558 1.93989
R833 VTAIL.n34 VTAIL.n33 1.93989
R834 VTAIL.n66 VTAIL.n6 1.93989
R835 VTAIL.n112 VTAIL.n111 1.93989
R836 VTAIL.n144 VTAIL.n84 1.93989
R837 VTAIL.n192 VTAIL.n191 1.93989
R838 VTAIL.n224 VTAIL.n164 1.93989
R839 VTAIL.n541 VTAIL.n481 1.93989
R840 VTAIL.n509 VTAIL.n508 1.93989
R841 VTAIL.n461 VTAIL.n401 1.93989
R842 VTAIL.n429 VTAIL.n428 1.93989
R843 VTAIL.n383 VTAIL.n323 1.93989
R844 VTAIL.n351 VTAIL.n350 1.93989
R845 VTAIL.n303 VTAIL.n243 1.93989
R846 VTAIL.n271 VTAIL.n270 1.93989
R847 VTAIL.n317 VTAIL.n315 1.57809
R848 VTAIL.n395 VTAIL.n317 1.57809
R849 VTAIL.n475 VTAIL.n473 1.57809
R850 VTAIL.n553 VTAIL.n475 1.57809
R851 VTAIL.n237 VTAIL.n159 1.57809
R852 VTAIL.n159 VTAIL.n157 1.57809
R853 VTAIL.n79 VTAIL.n1 1.57809
R854 VTAIL VTAIL.n631 1.5199
R855 VTAIL.n0 VTAIL.t4 1.41277
R856 VTAIL.n0 VTAIL.t7 1.41277
R857 VTAIL.n158 VTAIL.t13 1.41277
R858 VTAIL.n158 VTAIL.t9 1.41277
R859 VTAIL.n474 VTAIL.t12 1.41277
R860 VTAIL.n474 VTAIL.t15 1.41277
R861 VTAIL.n316 VTAIL.t5 1.41277
R862 VTAIL.n316 VTAIL.t2 1.41277
R863 VTAIL.n582 VTAIL.n576 1.16414
R864 VTAIL.n623 VTAIL.n621 1.16414
R865 VTAIL.n630 VTAIL.n554 1.16414
R866 VTAIL.n30 VTAIL.n24 1.16414
R867 VTAIL.n71 VTAIL.n69 1.16414
R868 VTAIL.n78 VTAIL.n2 1.16414
R869 VTAIL.n108 VTAIL.n102 1.16414
R870 VTAIL.n149 VTAIL.n147 1.16414
R871 VTAIL.n156 VTAIL.n80 1.16414
R872 VTAIL.n188 VTAIL.n182 1.16414
R873 VTAIL.n229 VTAIL.n227 1.16414
R874 VTAIL.n236 VTAIL.n160 1.16414
R875 VTAIL.n552 VTAIL.n476 1.16414
R876 VTAIL.n545 VTAIL.n544 1.16414
R877 VTAIL.n505 VTAIL.n499 1.16414
R878 VTAIL.n472 VTAIL.n396 1.16414
R879 VTAIL.n465 VTAIL.n464 1.16414
R880 VTAIL.n425 VTAIL.n419 1.16414
R881 VTAIL.n394 VTAIL.n318 1.16414
R882 VTAIL.n387 VTAIL.n386 1.16414
R883 VTAIL.n347 VTAIL.n341 1.16414
R884 VTAIL.n314 VTAIL.n238 1.16414
R885 VTAIL.n307 VTAIL.n306 1.16414
R886 VTAIL.n267 VTAIL.n261 1.16414
R887 VTAIL.n473 VTAIL.n395 0.470328
R888 VTAIL.n157 VTAIL.n79 0.470328
R889 VTAIL.n581 VTAIL.n578 0.388379
R890 VTAIL.n622 VTAIL.n556 0.388379
R891 VTAIL.n628 VTAIL.n627 0.388379
R892 VTAIL.n29 VTAIL.n26 0.388379
R893 VTAIL.n70 VTAIL.n4 0.388379
R894 VTAIL.n76 VTAIL.n75 0.388379
R895 VTAIL.n107 VTAIL.n104 0.388379
R896 VTAIL.n148 VTAIL.n82 0.388379
R897 VTAIL.n154 VTAIL.n153 0.388379
R898 VTAIL.n187 VTAIL.n184 0.388379
R899 VTAIL.n228 VTAIL.n162 0.388379
R900 VTAIL.n234 VTAIL.n233 0.388379
R901 VTAIL.n550 VTAIL.n549 0.388379
R902 VTAIL.n480 VTAIL.n478 0.388379
R903 VTAIL.n504 VTAIL.n501 0.388379
R904 VTAIL.n470 VTAIL.n469 0.388379
R905 VTAIL.n400 VTAIL.n398 0.388379
R906 VTAIL.n424 VTAIL.n421 0.388379
R907 VTAIL.n392 VTAIL.n391 0.388379
R908 VTAIL.n322 VTAIL.n320 0.388379
R909 VTAIL.n346 VTAIL.n343 0.388379
R910 VTAIL.n312 VTAIL.n311 0.388379
R911 VTAIL.n242 VTAIL.n240 0.388379
R912 VTAIL.n266 VTAIL.n263 0.388379
R913 VTAIL.n580 VTAIL.n575 0.155672
R914 VTAIL.n587 VTAIL.n575 0.155672
R915 VTAIL.n588 VTAIL.n587 0.155672
R916 VTAIL.n588 VTAIL.n571 0.155672
R917 VTAIL.n595 VTAIL.n571 0.155672
R918 VTAIL.n596 VTAIL.n595 0.155672
R919 VTAIL.n596 VTAIL.n567 0.155672
R920 VTAIL.n603 VTAIL.n567 0.155672
R921 VTAIL.n604 VTAIL.n603 0.155672
R922 VTAIL.n604 VTAIL.n563 0.155672
R923 VTAIL.n611 VTAIL.n563 0.155672
R924 VTAIL.n612 VTAIL.n611 0.155672
R925 VTAIL.n612 VTAIL.n559 0.155672
R926 VTAIL.n619 VTAIL.n559 0.155672
R927 VTAIL.n620 VTAIL.n619 0.155672
R928 VTAIL.n620 VTAIL.n555 0.155672
R929 VTAIL.n629 VTAIL.n555 0.155672
R930 VTAIL.n28 VTAIL.n23 0.155672
R931 VTAIL.n35 VTAIL.n23 0.155672
R932 VTAIL.n36 VTAIL.n35 0.155672
R933 VTAIL.n36 VTAIL.n19 0.155672
R934 VTAIL.n43 VTAIL.n19 0.155672
R935 VTAIL.n44 VTAIL.n43 0.155672
R936 VTAIL.n44 VTAIL.n15 0.155672
R937 VTAIL.n51 VTAIL.n15 0.155672
R938 VTAIL.n52 VTAIL.n51 0.155672
R939 VTAIL.n52 VTAIL.n11 0.155672
R940 VTAIL.n59 VTAIL.n11 0.155672
R941 VTAIL.n60 VTAIL.n59 0.155672
R942 VTAIL.n60 VTAIL.n7 0.155672
R943 VTAIL.n67 VTAIL.n7 0.155672
R944 VTAIL.n68 VTAIL.n67 0.155672
R945 VTAIL.n68 VTAIL.n3 0.155672
R946 VTAIL.n77 VTAIL.n3 0.155672
R947 VTAIL.n106 VTAIL.n101 0.155672
R948 VTAIL.n113 VTAIL.n101 0.155672
R949 VTAIL.n114 VTAIL.n113 0.155672
R950 VTAIL.n114 VTAIL.n97 0.155672
R951 VTAIL.n121 VTAIL.n97 0.155672
R952 VTAIL.n122 VTAIL.n121 0.155672
R953 VTAIL.n122 VTAIL.n93 0.155672
R954 VTAIL.n129 VTAIL.n93 0.155672
R955 VTAIL.n130 VTAIL.n129 0.155672
R956 VTAIL.n130 VTAIL.n89 0.155672
R957 VTAIL.n137 VTAIL.n89 0.155672
R958 VTAIL.n138 VTAIL.n137 0.155672
R959 VTAIL.n138 VTAIL.n85 0.155672
R960 VTAIL.n145 VTAIL.n85 0.155672
R961 VTAIL.n146 VTAIL.n145 0.155672
R962 VTAIL.n146 VTAIL.n81 0.155672
R963 VTAIL.n155 VTAIL.n81 0.155672
R964 VTAIL.n186 VTAIL.n181 0.155672
R965 VTAIL.n193 VTAIL.n181 0.155672
R966 VTAIL.n194 VTAIL.n193 0.155672
R967 VTAIL.n194 VTAIL.n177 0.155672
R968 VTAIL.n201 VTAIL.n177 0.155672
R969 VTAIL.n202 VTAIL.n201 0.155672
R970 VTAIL.n202 VTAIL.n173 0.155672
R971 VTAIL.n209 VTAIL.n173 0.155672
R972 VTAIL.n210 VTAIL.n209 0.155672
R973 VTAIL.n210 VTAIL.n169 0.155672
R974 VTAIL.n217 VTAIL.n169 0.155672
R975 VTAIL.n218 VTAIL.n217 0.155672
R976 VTAIL.n218 VTAIL.n165 0.155672
R977 VTAIL.n225 VTAIL.n165 0.155672
R978 VTAIL.n226 VTAIL.n225 0.155672
R979 VTAIL.n226 VTAIL.n161 0.155672
R980 VTAIL.n235 VTAIL.n161 0.155672
R981 VTAIL.n551 VTAIL.n477 0.155672
R982 VTAIL.n543 VTAIL.n477 0.155672
R983 VTAIL.n543 VTAIL.n542 0.155672
R984 VTAIL.n542 VTAIL.n482 0.155672
R985 VTAIL.n535 VTAIL.n482 0.155672
R986 VTAIL.n535 VTAIL.n534 0.155672
R987 VTAIL.n534 VTAIL.n486 0.155672
R988 VTAIL.n527 VTAIL.n486 0.155672
R989 VTAIL.n527 VTAIL.n526 0.155672
R990 VTAIL.n526 VTAIL.n490 0.155672
R991 VTAIL.n519 VTAIL.n490 0.155672
R992 VTAIL.n519 VTAIL.n518 0.155672
R993 VTAIL.n518 VTAIL.n494 0.155672
R994 VTAIL.n511 VTAIL.n494 0.155672
R995 VTAIL.n511 VTAIL.n510 0.155672
R996 VTAIL.n510 VTAIL.n498 0.155672
R997 VTAIL.n503 VTAIL.n498 0.155672
R998 VTAIL.n471 VTAIL.n397 0.155672
R999 VTAIL.n463 VTAIL.n397 0.155672
R1000 VTAIL.n463 VTAIL.n462 0.155672
R1001 VTAIL.n462 VTAIL.n402 0.155672
R1002 VTAIL.n455 VTAIL.n402 0.155672
R1003 VTAIL.n455 VTAIL.n454 0.155672
R1004 VTAIL.n454 VTAIL.n406 0.155672
R1005 VTAIL.n447 VTAIL.n406 0.155672
R1006 VTAIL.n447 VTAIL.n446 0.155672
R1007 VTAIL.n446 VTAIL.n410 0.155672
R1008 VTAIL.n439 VTAIL.n410 0.155672
R1009 VTAIL.n439 VTAIL.n438 0.155672
R1010 VTAIL.n438 VTAIL.n414 0.155672
R1011 VTAIL.n431 VTAIL.n414 0.155672
R1012 VTAIL.n431 VTAIL.n430 0.155672
R1013 VTAIL.n430 VTAIL.n418 0.155672
R1014 VTAIL.n423 VTAIL.n418 0.155672
R1015 VTAIL.n393 VTAIL.n319 0.155672
R1016 VTAIL.n385 VTAIL.n319 0.155672
R1017 VTAIL.n385 VTAIL.n384 0.155672
R1018 VTAIL.n384 VTAIL.n324 0.155672
R1019 VTAIL.n377 VTAIL.n324 0.155672
R1020 VTAIL.n377 VTAIL.n376 0.155672
R1021 VTAIL.n376 VTAIL.n328 0.155672
R1022 VTAIL.n369 VTAIL.n328 0.155672
R1023 VTAIL.n369 VTAIL.n368 0.155672
R1024 VTAIL.n368 VTAIL.n332 0.155672
R1025 VTAIL.n361 VTAIL.n332 0.155672
R1026 VTAIL.n361 VTAIL.n360 0.155672
R1027 VTAIL.n360 VTAIL.n336 0.155672
R1028 VTAIL.n353 VTAIL.n336 0.155672
R1029 VTAIL.n353 VTAIL.n352 0.155672
R1030 VTAIL.n352 VTAIL.n340 0.155672
R1031 VTAIL.n345 VTAIL.n340 0.155672
R1032 VTAIL.n313 VTAIL.n239 0.155672
R1033 VTAIL.n305 VTAIL.n239 0.155672
R1034 VTAIL.n305 VTAIL.n304 0.155672
R1035 VTAIL.n304 VTAIL.n244 0.155672
R1036 VTAIL.n297 VTAIL.n244 0.155672
R1037 VTAIL.n297 VTAIL.n296 0.155672
R1038 VTAIL.n296 VTAIL.n248 0.155672
R1039 VTAIL.n289 VTAIL.n248 0.155672
R1040 VTAIL.n289 VTAIL.n288 0.155672
R1041 VTAIL.n288 VTAIL.n252 0.155672
R1042 VTAIL.n281 VTAIL.n252 0.155672
R1043 VTAIL.n281 VTAIL.n280 0.155672
R1044 VTAIL.n280 VTAIL.n256 0.155672
R1045 VTAIL.n273 VTAIL.n256 0.155672
R1046 VTAIL.n273 VTAIL.n272 0.155672
R1047 VTAIL.n272 VTAIL.n260 0.155672
R1048 VTAIL.n265 VTAIL.n260 0.155672
R1049 VTAIL VTAIL.n1 0.0586897
R1050 B.n816 B.n815 585
R1051 B.n817 B.n816 585
R1052 B.n329 B.n119 585
R1053 B.n328 B.n327 585
R1054 B.n326 B.n325 585
R1055 B.n324 B.n323 585
R1056 B.n322 B.n321 585
R1057 B.n320 B.n319 585
R1058 B.n318 B.n317 585
R1059 B.n316 B.n315 585
R1060 B.n314 B.n313 585
R1061 B.n312 B.n311 585
R1062 B.n310 B.n309 585
R1063 B.n308 B.n307 585
R1064 B.n306 B.n305 585
R1065 B.n304 B.n303 585
R1066 B.n302 B.n301 585
R1067 B.n300 B.n299 585
R1068 B.n298 B.n297 585
R1069 B.n296 B.n295 585
R1070 B.n294 B.n293 585
R1071 B.n292 B.n291 585
R1072 B.n290 B.n289 585
R1073 B.n288 B.n287 585
R1074 B.n286 B.n285 585
R1075 B.n284 B.n283 585
R1076 B.n282 B.n281 585
R1077 B.n280 B.n279 585
R1078 B.n278 B.n277 585
R1079 B.n276 B.n275 585
R1080 B.n274 B.n273 585
R1081 B.n272 B.n271 585
R1082 B.n270 B.n269 585
R1083 B.n268 B.n267 585
R1084 B.n266 B.n265 585
R1085 B.n264 B.n263 585
R1086 B.n262 B.n261 585
R1087 B.n260 B.n259 585
R1088 B.n258 B.n257 585
R1089 B.n256 B.n255 585
R1090 B.n254 B.n253 585
R1091 B.n252 B.n251 585
R1092 B.n250 B.n249 585
R1093 B.n248 B.n247 585
R1094 B.n246 B.n245 585
R1095 B.n244 B.n243 585
R1096 B.n242 B.n241 585
R1097 B.n240 B.n239 585
R1098 B.n238 B.n237 585
R1099 B.n235 B.n234 585
R1100 B.n233 B.n232 585
R1101 B.n231 B.n230 585
R1102 B.n229 B.n228 585
R1103 B.n227 B.n226 585
R1104 B.n225 B.n224 585
R1105 B.n223 B.n222 585
R1106 B.n221 B.n220 585
R1107 B.n219 B.n218 585
R1108 B.n217 B.n216 585
R1109 B.n215 B.n214 585
R1110 B.n213 B.n212 585
R1111 B.n211 B.n210 585
R1112 B.n209 B.n208 585
R1113 B.n207 B.n206 585
R1114 B.n205 B.n204 585
R1115 B.n203 B.n202 585
R1116 B.n201 B.n200 585
R1117 B.n199 B.n198 585
R1118 B.n197 B.n196 585
R1119 B.n195 B.n194 585
R1120 B.n193 B.n192 585
R1121 B.n191 B.n190 585
R1122 B.n189 B.n188 585
R1123 B.n187 B.n186 585
R1124 B.n185 B.n184 585
R1125 B.n183 B.n182 585
R1126 B.n181 B.n180 585
R1127 B.n179 B.n178 585
R1128 B.n177 B.n176 585
R1129 B.n175 B.n174 585
R1130 B.n173 B.n172 585
R1131 B.n171 B.n170 585
R1132 B.n169 B.n168 585
R1133 B.n167 B.n166 585
R1134 B.n165 B.n164 585
R1135 B.n163 B.n162 585
R1136 B.n161 B.n160 585
R1137 B.n159 B.n158 585
R1138 B.n157 B.n156 585
R1139 B.n155 B.n154 585
R1140 B.n153 B.n152 585
R1141 B.n151 B.n150 585
R1142 B.n149 B.n148 585
R1143 B.n147 B.n146 585
R1144 B.n145 B.n144 585
R1145 B.n143 B.n142 585
R1146 B.n141 B.n140 585
R1147 B.n139 B.n138 585
R1148 B.n137 B.n136 585
R1149 B.n135 B.n134 585
R1150 B.n133 B.n132 585
R1151 B.n131 B.n130 585
R1152 B.n129 B.n128 585
R1153 B.n127 B.n126 585
R1154 B.n67 B.n66 585
R1155 B.n820 B.n819 585
R1156 B.n814 B.n120 585
R1157 B.n120 B.n64 585
R1158 B.n813 B.n63 585
R1159 B.n824 B.n63 585
R1160 B.n812 B.n62 585
R1161 B.n825 B.n62 585
R1162 B.n811 B.n61 585
R1163 B.n826 B.n61 585
R1164 B.n810 B.n809 585
R1165 B.n809 B.n57 585
R1166 B.n808 B.n56 585
R1167 B.n832 B.n56 585
R1168 B.n807 B.n55 585
R1169 B.n833 B.n55 585
R1170 B.n806 B.n54 585
R1171 B.n834 B.n54 585
R1172 B.n805 B.n804 585
R1173 B.n804 B.n50 585
R1174 B.n803 B.n49 585
R1175 B.n840 B.n49 585
R1176 B.n802 B.n48 585
R1177 B.n841 B.n48 585
R1178 B.n801 B.n47 585
R1179 B.n842 B.n47 585
R1180 B.n800 B.n799 585
R1181 B.n799 B.n43 585
R1182 B.n798 B.n42 585
R1183 B.n848 B.n42 585
R1184 B.n797 B.n41 585
R1185 B.n849 B.n41 585
R1186 B.n796 B.n40 585
R1187 B.n850 B.n40 585
R1188 B.n795 B.n794 585
R1189 B.n794 B.n36 585
R1190 B.n793 B.n35 585
R1191 B.n856 B.n35 585
R1192 B.n792 B.n34 585
R1193 B.n857 B.n34 585
R1194 B.n791 B.n33 585
R1195 B.n858 B.n33 585
R1196 B.n790 B.n789 585
R1197 B.n789 B.n29 585
R1198 B.n788 B.n28 585
R1199 B.n864 B.n28 585
R1200 B.n787 B.n27 585
R1201 B.n865 B.n27 585
R1202 B.n786 B.n26 585
R1203 B.n866 B.n26 585
R1204 B.n785 B.n784 585
R1205 B.n784 B.n22 585
R1206 B.n783 B.n21 585
R1207 B.n872 B.n21 585
R1208 B.n782 B.n20 585
R1209 B.n873 B.n20 585
R1210 B.n781 B.n19 585
R1211 B.n874 B.n19 585
R1212 B.n780 B.n779 585
R1213 B.n779 B.n15 585
R1214 B.n778 B.n14 585
R1215 B.n880 B.n14 585
R1216 B.n777 B.n13 585
R1217 B.n881 B.n13 585
R1218 B.n776 B.n12 585
R1219 B.n882 B.n12 585
R1220 B.n775 B.n774 585
R1221 B.n774 B.n8 585
R1222 B.n773 B.n7 585
R1223 B.n888 B.n7 585
R1224 B.n772 B.n6 585
R1225 B.n889 B.n6 585
R1226 B.n771 B.n5 585
R1227 B.n890 B.n5 585
R1228 B.n770 B.n769 585
R1229 B.n769 B.n4 585
R1230 B.n768 B.n330 585
R1231 B.n768 B.n767 585
R1232 B.n758 B.n331 585
R1233 B.n332 B.n331 585
R1234 B.n760 B.n759 585
R1235 B.n761 B.n760 585
R1236 B.n757 B.n336 585
R1237 B.n340 B.n336 585
R1238 B.n756 B.n755 585
R1239 B.n755 B.n754 585
R1240 B.n338 B.n337 585
R1241 B.n339 B.n338 585
R1242 B.n747 B.n746 585
R1243 B.n748 B.n747 585
R1244 B.n745 B.n345 585
R1245 B.n345 B.n344 585
R1246 B.n744 B.n743 585
R1247 B.n743 B.n742 585
R1248 B.n347 B.n346 585
R1249 B.n348 B.n347 585
R1250 B.n735 B.n734 585
R1251 B.n736 B.n735 585
R1252 B.n733 B.n353 585
R1253 B.n353 B.n352 585
R1254 B.n732 B.n731 585
R1255 B.n731 B.n730 585
R1256 B.n355 B.n354 585
R1257 B.n356 B.n355 585
R1258 B.n723 B.n722 585
R1259 B.n724 B.n723 585
R1260 B.n721 B.n361 585
R1261 B.n361 B.n360 585
R1262 B.n720 B.n719 585
R1263 B.n719 B.n718 585
R1264 B.n363 B.n362 585
R1265 B.n364 B.n363 585
R1266 B.n711 B.n710 585
R1267 B.n712 B.n711 585
R1268 B.n709 B.n368 585
R1269 B.n372 B.n368 585
R1270 B.n708 B.n707 585
R1271 B.n707 B.n706 585
R1272 B.n370 B.n369 585
R1273 B.n371 B.n370 585
R1274 B.n699 B.n698 585
R1275 B.n700 B.n699 585
R1276 B.n697 B.n377 585
R1277 B.n377 B.n376 585
R1278 B.n696 B.n695 585
R1279 B.n695 B.n694 585
R1280 B.n379 B.n378 585
R1281 B.n380 B.n379 585
R1282 B.n687 B.n686 585
R1283 B.n688 B.n687 585
R1284 B.n685 B.n385 585
R1285 B.n385 B.n384 585
R1286 B.n684 B.n683 585
R1287 B.n683 B.n682 585
R1288 B.n387 B.n386 585
R1289 B.n388 B.n387 585
R1290 B.n675 B.n674 585
R1291 B.n676 B.n675 585
R1292 B.n673 B.n393 585
R1293 B.n393 B.n392 585
R1294 B.n672 B.n671 585
R1295 B.n671 B.n670 585
R1296 B.n395 B.n394 585
R1297 B.n396 B.n395 585
R1298 B.n666 B.n665 585
R1299 B.n399 B.n398 585
R1300 B.n662 B.n661 585
R1301 B.n663 B.n662 585
R1302 B.n660 B.n451 585
R1303 B.n659 B.n658 585
R1304 B.n657 B.n656 585
R1305 B.n655 B.n654 585
R1306 B.n653 B.n652 585
R1307 B.n651 B.n650 585
R1308 B.n649 B.n648 585
R1309 B.n647 B.n646 585
R1310 B.n645 B.n644 585
R1311 B.n643 B.n642 585
R1312 B.n641 B.n640 585
R1313 B.n639 B.n638 585
R1314 B.n637 B.n636 585
R1315 B.n635 B.n634 585
R1316 B.n633 B.n632 585
R1317 B.n631 B.n630 585
R1318 B.n629 B.n628 585
R1319 B.n627 B.n626 585
R1320 B.n625 B.n624 585
R1321 B.n623 B.n622 585
R1322 B.n621 B.n620 585
R1323 B.n619 B.n618 585
R1324 B.n617 B.n616 585
R1325 B.n615 B.n614 585
R1326 B.n613 B.n612 585
R1327 B.n611 B.n610 585
R1328 B.n609 B.n608 585
R1329 B.n607 B.n606 585
R1330 B.n605 B.n604 585
R1331 B.n603 B.n602 585
R1332 B.n601 B.n600 585
R1333 B.n599 B.n598 585
R1334 B.n597 B.n596 585
R1335 B.n595 B.n594 585
R1336 B.n593 B.n592 585
R1337 B.n591 B.n590 585
R1338 B.n589 B.n588 585
R1339 B.n587 B.n586 585
R1340 B.n585 B.n584 585
R1341 B.n583 B.n582 585
R1342 B.n581 B.n580 585
R1343 B.n579 B.n578 585
R1344 B.n577 B.n576 585
R1345 B.n575 B.n574 585
R1346 B.n573 B.n572 585
R1347 B.n570 B.n569 585
R1348 B.n568 B.n567 585
R1349 B.n566 B.n565 585
R1350 B.n564 B.n563 585
R1351 B.n562 B.n561 585
R1352 B.n560 B.n559 585
R1353 B.n558 B.n557 585
R1354 B.n556 B.n555 585
R1355 B.n554 B.n553 585
R1356 B.n552 B.n551 585
R1357 B.n550 B.n549 585
R1358 B.n548 B.n547 585
R1359 B.n546 B.n545 585
R1360 B.n544 B.n543 585
R1361 B.n542 B.n541 585
R1362 B.n540 B.n539 585
R1363 B.n538 B.n537 585
R1364 B.n536 B.n535 585
R1365 B.n534 B.n533 585
R1366 B.n532 B.n531 585
R1367 B.n530 B.n529 585
R1368 B.n528 B.n527 585
R1369 B.n526 B.n525 585
R1370 B.n524 B.n523 585
R1371 B.n522 B.n521 585
R1372 B.n520 B.n519 585
R1373 B.n518 B.n517 585
R1374 B.n516 B.n515 585
R1375 B.n514 B.n513 585
R1376 B.n512 B.n511 585
R1377 B.n510 B.n509 585
R1378 B.n508 B.n507 585
R1379 B.n506 B.n505 585
R1380 B.n504 B.n503 585
R1381 B.n502 B.n501 585
R1382 B.n500 B.n499 585
R1383 B.n498 B.n497 585
R1384 B.n496 B.n495 585
R1385 B.n494 B.n493 585
R1386 B.n492 B.n491 585
R1387 B.n490 B.n489 585
R1388 B.n488 B.n487 585
R1389 B.n486 B.n485 585
R1390 B.n484 B.n483 585
R1391 B.n482 B.n481 585
R1392 B.n480 B.n479 585
R1393 B.n478 B.n477 585
R1394 B.n476 B.n475 585
R1395 B.n474 B.n473 585
R1396 B.n472 B.n471 585
R1397 B.n470 B.n469 585
R1398 B.n468 B.n467 585
R1399 B.n466 B.n465 585
R1400 B.n464 B.n463 585
R1401 B.n462 B.n461 585
R1402 B.n460 B.n459 585
R1403 B.n458 B.n457 585
R1404 B.n667 B.n397 585
R1405 B.n397 B.n396 585
R1406 B.n669 B.n668 585
R1407 B.n670 B.n669 585
R1408 B.n391 B.n390 585
R1409 B.n392 B.n391 585
R1410 B.n678 B.n677 585
R1411 B.n677 B.n676 585
R1412 B.n679 B.n389 585
R1413 B.n389 B.n388 585
R1414 B.n681 B.n680 585
R1415 B.n682 B.n681 585
R1416 B.n383 B.n382 585
R1417 B.n384 B.n383 585
R1418 B.n690 B.n689 585
R1419 B.n689 B.n688 585
R1420 B.n691 B.n381 585
R1421 B.n381 B.n380 585
R1422 B.n693 B.n692 585
R1423 B.n694 B.n693 585
R1424 B.n375 B.n374 585
R1425 B.n376 B.n375 585
R1426 B.n702 B.n701 585
R1427 B.n701 B.n700 585
R1428 B.n703 B.n373 585
R1429 B.n373 B.n371 585
R1430 B.n705 B.n704 585
R1431 B.n706 B.n705 585
R1432 B.n367 B.n366 585
R1433 B.n372 B.n367 585
R1434 B.n714 B.n713 585
R1435 B.n713 B.n712 585
R1436 B.n715 B.n365 585
R1437 B.n365 B.n364 585
R1438 B.n717 B.n716 585
R1439 B.n718 B.n717 585
R1440 B.n359 B.n358 585
R1441 B.n360 B.n359 585
R1442 B.n726 B.n725 585
R1443 B.n725 B.n724 585
R1444 B.n727 B.n357 585
R1445 B.n357 B.n356 585
R1446 B.n729 B.n728 585
R1447 B.n730 B.n729 585
R1448 B.n351 B.n350 585
R1449 B.n352 B.n351 585
R1450 B.n738 B.n737 585
R1451 B.n737 B.n736 585
R1452 B.n739 B.n349 585
R1453 B.n349 B.n348 585
R1454 B.n741 B.n740 585
R1455 B.n742 B.n741 585
R1456 B.n343 B.n342 585
R1457 B.n344 B.n343 585
R1458 B.n750 B.n749 585
R1459 B.n749 B.n748 585
R1460 B.n751 B.n341 585
R1461 B.n341 B.n339 585
R1462 B.n753 B.n752 585
R1463 B.n754 B.n753 585
R1464 B.n335 B.n334 585
R1465 B.n340 B.n335 585
R1466 B.n763 B.n762 585
R1467 B.n762 B.n761 585
R1468 B.n764 B.n333 585
R1469 B.n333 B.n332 585
R1470 B.n766 B.n765 585
R1471 B.n767 B.n766 585
R1472 B.n2 B.n0 585
R1473 B.n4 B.n2 585
R1474 B.n3 B.n1 585
R1475 B.n889 B.n3 585
R1476 B.n887 B.n886 585
R1477 B.n888 B.n887 585
R1478 B.n885 B.n9 585
R1479 B.n9 B.n8 585
R1480 B.n884 B.n883 585
R1481 B.n883 B.n882 585
R1482 B.n11 B.n10 585
R1483 B.n881 B.n11 585
R1484 B.n879 B.n878 585
R1485 B.n880 B.n879 585
R1486 B.n877 B.n16 585
R1487 B.n16 B.n15 585
R1488 B.n876 B.n875 585
R1489 B.n875 B.n874 585
R1490 B.n18 B.n17 585
R1491 B.n873 B.n18 585
R1492 B.n871 B.n870 585
R1493 B.n872 B.n871 585
R1494 B.n869 B.n23 585
R1495 B.n23 B.n22 585
R1496 B.n868 B.n867 585
R1497 B.n867 B.n866 585
R1498 B.n25 B.n24 585
R1499 B.n865 B.n25 585
R1500 B.n863 B.n862 585
R1501 B.n864 B.n863 585
R1502 B.n861 B.n30 585
R1503 B.n30 B.n29 585
R1504 B.n860 B.n859 585
R1505 B.n859 B.n858 585
R1506 B.n32 B.n31 585
R1507 B.n857 B.n32 585
R1508 B.n855 B.n854 585
R1509 B.n856 B.n855 585
R1510 B.n853 B.n37 585
R1511 B.n37 B.n36 585
R1512 B.n852 B.n851 585
R1513 B.n851 B.n850 585
R1514 B.n39 B.n38 585
R1515 B.n849 B.n39 585
R1516 B.n847 B.n846 585
R1517 B.n848 B.n847 585
R1518 B.n845 B.n44 585
R1519 B.n44 B.n43 585
R1520 B.n844 B.n843 585
R1521 B.n843 B.n842 585
R1522 B.n46 B.n45 585
R1523 B.n841 B.n46 585
R1524 B.n839 B.n838 585
R1525 B.n840 B.n839 585
R1526 B.n837 B.n51 585
R1527 B.n51 B.n50 585
R1528 B.n836 B.n835 585
R1529 B.n835 B.n834 585
R1530 B.n53 B.n52 585
R1531 B.n833 B.n53 585
R1532 B.n831 B.n830 585
R1533 B.n832 B.n831 585
R1534 B.n829 B.n58 585
R1535 B.n58 B.n57 585
R1536 B.n828 B.n827 585
R1537 B.n827 B.n826 585
R1538 B.n60 B.n59 585
R1539 B.n825 B.n60 585
R1540 B.n823 B.n822 585
R1541 B.n824 B.n823 585
R1542 B.n821 B.n65 585
R1543 B.n65 B.n64 585
R1544 B.n892 B.n891 585
R1545 B.n891 B.n890 585
R1546 B.n665 B.n397 478.086
R1547 B.n819 B.n65 478.086
R1548 B.n457 B.n395 478.086
R1549 B.n816 B.n120 478.086
R1550 B.n454 B.t16 430.695
R1551 B.n452 B.t8 430.695
R1552 B.n123 B.t19 430.695
R1553 B.n121 B.t12 430.695
R1554 B.n454 B.t18 352.248
R1555 B.n121 B.t14 352.248
R1556 B.n452 B.t11 352.248
R1557 B.n123 B.t20 352.248
R1558 B.n455 B.t17 316.757
R1559 B.n122 B.t15 316.757
R1560 B.n453 B.t10 316.757
R1561 B.n124 B.t21 316.757
R1562 B.n817 B.n118 256.663
R1563 B.n817 B.n117 256.663
R1564 B.n817 B.n116 256.663
R1565 B.n817 B.n115 256.663
R1566 B.n817 B.n114 256.663
R1567 B.n817 B.n113 256.663
R1568 B.n817 B.n112 256.663
R1569 B.n817 B.n111 256.663
R1570 B.n817 B.n110 256.663
R1571 B.n817 B.n109 256.663
R1572 B.n817 B.n108 256.663
R1573 B.n817 B.n107 256.663
R1574 B.n817 B.n106 256.663
R1575 B.n817 B.n105 256.663
R1576 B.n817 B.n104 256.663
R1577 B.n817 B.n103 256.663
R1578 B.n817 B.n102 256.663
R1579 B.n817 B.n101 256.663
R1580 B.n817 B.n100 256.663
R1581 B.n817 B.n99 256.663
R1582 B.n817 B.n98 256.663
R1583 B.n817 B.n97 256.663
R1584 B.n817 B.n96 256.663
R1585 B.n817 B.n95 256.663
R1586 B.n817 B.n94 256.663
R1587 B.n817 B.n93 256.663
R1588 B.n817 B.n92 256.663
R1589 B.n817 B.n91 256.663
R1590 B.n817 B.n90 256.663
R1591 B.n817 B.n89 256.663
R1592 B.n817 B.n88 256.663
R1593 B.n817 B.n87 256.663
R1594 B.n817 B.n86 256.663
R1595 B.n817 B.n85 256.663
R1596 B.n817 B.n84 256.663
R1597 B.n817 B.n83 256.663
R1598 B.n817 B.n82 256.663
R1599 B.n817 B.n81 256.663
R1600 B.n817 B.n80 256.663
R1601 B.n817 B.n79 256.663
R1602 B.n817 B.n78 256.663
R1603 B.n817 B.n77 256.663
R1604 B.n817 B.n76 256.663
R1605 B.n817 B.n75 256.663
R1606 B.n817 B.n74 256.663
R1607 B.n817 B.n73 256.663
R1608 B.n817 B.n72 256.663
R1609 B.n817 B.n71 256.663
R1610 B.n817 B.n70 256.663
R1611 B.n817 B.n69 256.663
R1612 B.n817 B.n68 256.663
R1613 B.n818 B.n817 256.663
R1614 B.n664 B.n663 256.663
R1615 B.n663 B.n400 256.663
R1616 B.n663 B.n401 256.663
R1617 B.n663 B.n402 256.663
R1618 B.n663 B.n403 256.663
R1619 B.n663 B.n404 256.663
R1620 B.n663 B.n405 256.663
R1621 B.n663 B.n406 256.663
R1622 B.n663 B.n407 256.663
R1623 B.n663 B.n408 256.663
R1624 B.n663 B.n409 256.663
R1625 B.n663 B.n410 256.663
R1626 B.n663 B.n411 256.663
R1627 B.n663 B.n412 256.663
R1628 B.n663 B.n413 256.663
R1629 B.n663 B.n414 256.663
R1630 B.n663 B.n415 256.663
R1631 B.n663 B.n416 256.663
R1632 B.n663 B.n417 256.663
R1633 B.n663 B.n418 256.663
R1634 B.n663 B.n419 256.663
R1635 B.n663 B.n420 256.663
R1636 B.n663 B.n421 256.663
R1637 B.n663 B.n422 256.663
R1638 B.n663 B.n423 256.663
R1639 B.n663 B.n424 256.663
R1640 B.n663 B.n425 256.663
R1641 B.n663 B.n426 256.663
R1642 B.n663 B.n427 256.663
R1643 B.n663 B.n428 256.663
R1644 B.n663 B.n429 256.663
R1645 B.n663 B.n430 256.663
R1646 B.n663 B.n431 256.663
R1647 B.n663 B.n432 256.663
R1648 B.n663 B.n433 256.663
R1649 B.n663 B.n434 256.663
R1650 B.n663 B.n435 256.663
R1651 B.n663 B.n436 256.663
R1652 B.n663 B.n437 256.663
R1653 B.n663 B.n438 256.663
R1654 B.n663 B.n439 256.663
R1655 B.n663 B.n440 256.663
R1656 B.n663 B.n441 256.663
R1657 B.n663 B.n442 256.663
R1658 B.n663 B.n443 256.663
R1659 B.n663 B.n444 256.663
R1660 B.n663 B.n445 256.663
R1661 B.n663 B.n446 256.663
R1662 B.n663 B.n447 256.663
R1663 B.n663 B.n448 256.663
R1664 B.n663 B.n449 256.663
R1665 B.n663 B.n450 256.663
R1666 B.n669 B.n397 163.367
R1667 B.n669 B.n391 163.367
R1668 B.n677 B.n391 163.367
R1669 B.n677 B.n389 163.367
R1670 B.n681 B.n389 163.367
R1671 B.n681 B.n383 163.367
R1672 B.n689 B.n383 163.367
R1673 B.n689 B.n381 163.367
R1674 B.n693 B.n381 163.367
R1675 B.n693 B.n375 163.367
R1676 B.n701 B.n375 163.367
R1677 B.n701 B.n373 163.367
R1678 B.n705 B.n373 163.367
R1679 B.n705 B.n367 163.367
R1680 B.n713 B.n367 163.367
R1681 B.n713 B.n365 163.367
R1682 B.n717 B.n365 163.367
R1683 B.n717 B.n359 163.367
R1684 B.n725 B.n359 163.367
R1685 B.n725 B.n357 163.367
R1686 B.n729 B.n357 163.367
R1687 B.n729 B.n351 163.367
R1688 B.n737 B.n351 163.367
R1689 B.n737 B.n349 163.367
R1690 B.n741 B.n349 163.367
R1691 B.n741 B.n343 163.367
R1692 B.n749 B.n343 163.367
R1693 B.n749 B.n341 163.367
R1694 B.n753 B.n341 163.367
R1695 B.n753 B.n335 163.367
R1696 B.n762 B.n335 163.367
R1697 B.n762 B.n333 163.367
R1698 B.n766 B.n333 163.367
R1699 B.n766 B.n2 163.367
R1700 B.n891 B.n2 163.367
R1701 B.n891 B.n3 163.367
R1702 B.n887 B.n3 163.367
R1703 B.n887 B.n9 163.367
R1704 B.n883 B.n9 163.367
R1705 B.n883 B.n11 163.367
R1706 B.n879 B.n11 163.367
R1707 B.n879 B.n16 163.367
R1708 B.n875 B.n16 163.367
R1709 B.n875 B.n18 163.367
R1710 B.n871 B.n18 163.367
R1711 B.n871 B.n23 163.367
R1712 B.n867 B.n23 163.367
R1713 B.n867 B.n25 163.367
R1714 B.n863 B.n25 163.367
R1715 B.n863 B.n30 163.367
R1716 B.n859 B.n30 163.367
R1717 B.n859 B.n32 163.367
R1718 B.n855 B.n32 163.367
R1719 B.n855 B.n37 163.367
R1720 B.n851 B.n37 163.367
R1721 B.n851 B.n39 163.367
R1722 B.n847 B.n39 163.367
R1723 B.n847 B.n44 163.367
R1724 B.n843 B.n44 163.367
R1725 B.n843 B.n46 163.367
R1726 B.n839 B.n46 163.367
R1727 B.n839 B.n51 163.367
R1728 B.n835 B.n51 163.367
R1729 B.n835 B.n53 163.367
R1730 B.n831 B.n53 163.367
R1731 B.n831 B.n58 163.367
R1732 B.n827 B.n58 163.367
R1733 B.n827 B.n60 163.367
R1734 B.n823 B.n60 163.367
R1735 B.n823 B.n65 163.367
R1736 B.n662 B.n399 163.367
R1737 B.n662 B.n451 163.367
R1738 B.n658 B.n657 163.367
R1739 B.n654 B.n653 163.367
R1740 B.n650 B.n649 163.367
R1741 B.n646 B.n645 163.367
R1742 B.n642 B.n641 163.367
R1743 B.n638 B.n637 163.367
R1744 B.n634 B.n633 163.367
R1745 B.n630 B.n629 163.367
R1746 B.n626 B.n625 163.367
R1747 B.n622 B.n621 163.367
R1748 B.n618 B.n617 163.367
R1749 B.n614 B.n613 163.367
R1750 B.n610 B.n609 163.367
R1751 B.n606 B.n605 163.367
R1752 B.n602 B.n601 163.367
R1753 B.n598 B.n597 163.367
R1754 B.n594 B.n593 163.367
R1755 B.n590 B.n589 163.367
R1756 B.n586 B.n585 163.367
R1757 B.n582 B.n581 163.367
R1758 B.n578 B.n577 163.367
R1759 B.n574 B.n573 163.367
R1760 B.n569 B.n568 163.367
R1761 B.n565 B.n564 163.367
R1762 B.n561 B.n560 163.367
R1763 B.n557 B.n556 163.367
R1764 B.n553 B.n552 163.367
R1765 B.n549 B.n548 163.367
R1766 B.n545 B.n544 163.367
R1767 B.n541 B.n540 163.367
R1768 B.n537 B.n536 163.367
R1769 B.n533 B.n532 163.367
R1770 B.n529 B.n528 163.367
R1771 B.n525 B.n524 163.367
R1772 B.n521 B.n520 163.367
R1773 B.n517 B.n516 163.367
R1774 B.n513 B.n512 163.367
R1775 B.n509 B.n508 163.367
R1776 B.n505 B.n504 163.367
R1777 B.n501 B.n500 163.367
R1778 B.n497 B.n496 163.367
R1779 B.n493 B.n492 163.367
R1780 B.n489 B.n488 163.367
R1781 B.n485 B.n484 163.367
R1782 B.n481 B.n480 163.367
R1783 B.n477 B.n476 163.367
R1784 B.n473 B.n472 163.367
R1785 B.n469 B.n468 163.367
R1786 B.n465 B.n464 163.367
R1787 B.n461 B.n460 163.367
R1788 B.n671 B.n395 163.367
R1789 B.n671 B.n393 163.367
R1790 B.n675 B.n393 163.367
R1791 B.n675 B.n387 163.367
R1792 B.n683 B.n387 163.367
R1793 B.n683 B.n385 163.367
R1794 B.n687 B.n385 163.367
R1795 B.n687 B.n379 163.367
R1796 B.n695 B.n379 163.367
R1797 B.n695 B.n377 163.367
R1798 B.n699 B.n377 163.367
R1799 B.n699 B.n370 163.367
R1800 B.n707 B.n370 163.367
R1801 B.n707 B.n368 163.367
R1802 B.n711 B.n368 163.367
R1803 B.n711 B.n363 163.367
R1804 B.n719 B.n363 163.367
R1805 B.n719 B.n361 163.367
R1806 B.n723 B.n361 163.367
R1807 B.n723 B.n355 163.367
R1808 B.n731 B.n355 163.367
R1809 B.n731 B.n353 163.367
R1810 B.n735 B.n353 163.367
R1811 B.n735 B.n347 163.367
R1812 B.n743 B.n347 163.367
R1813 B.n743 B.n345 163.367
R1814 B.n747 B.n345 163.367
R1815 B.n747 B.n338 163.367
R1816 B.n755 B.n338 163.367
R1817 B.n755 B.n336 163.367
R1818 B.n760 B.n336 163.367
R1819 B.n760 B.n331 163.367
R1820 B.n768 B.n331 163.367
R1821 B.n769 B.n768 163.367
R1822 B.n769 B.n5 163.367
R1823 B.n6 B.n5 163.367
R1824 B.n7 B.n6 163.367
R1825 B.n774 B.n7 163.367
R1826 B.n774 B.n12 163.367
R1827 B.n13 B.n12 163.367
R1828 B.n14 B.n13 163.367
R1829 B.n779 B.n14 163.367
R1830 B.n779 B.n19 163.367
R1831 B.n20 B.n19 163.367
R1832 B.n21 B.n20 163.367
R1833 B.n784 B.n21 163.367
R1834 B.n784 B.n26 163.367
R1835 B.n27 B.n26 163.367
R1836 B.n28 B.n27 163.367
R1837 B.n789 B.n28 163.367
R1838 B.n789 B.n33 163.367
R1839 B.n34 B.n33 163.367
R1840 B.n35 B.n34 163.367
R1841 B.n794 B.n35 163.367
R1842 B.n794 B.n40 163.367
R1843 B.n41 B.n40 163.367
R1844 B.n42 B.n41 163.367
R1845 B.n799 B.n42 163.367
R1846 B.n799 B.n47 163.367
R1847 B.n48 B.n47 163.367
R1848 B.n49 B.n48 163.367
R1849 B.n804 B.n49 163.367
R1850 B.n804 B.n54 163.367
R1851 B.n55 B.n54 163.367
R1852 B.n56 B.n55 163.367
R1853 B.n809 B.n56 163.367
R1854 B.n809 B.n61 163.367
R1855 B.n62 B.n61 163.367
R1856 B.n63 B.n62 163.367
R1857 B.n120 B.n63 163.367
R1858 B.n126 B.n67 163.367
R1859 B.n130 B.n129 163.367
R1860 B.n134 B.n133 163.367
R1861 B.n138 B.n137 163.367
R1862 B.n142 B.n141 163.367
R1863 B.n146 B.n145 163.367
R1864 B.n150 B.n149 163.367
R1865 B.n154 B.n153 163.367
R1866 B.n158 B.n157 163.367
R1867 B.n162 B.n161 163.367
R1868 B.n166 B.n165 163.367
R1869 B.n170 B.n169 163.367
R1870 B.n174 B.n173 163.367
R1871 B.n178 B.n177 163.367
R1872 B.n182 B.n181 163.367
R1873 B.n186 B.n185 163.367
R1874 B.n190 B.n189 163.367
R1875 B.n194 B.n193 163.367
R1876 B.n198 B.n197 163.367
R1877 B.n202 B.n201 163.367
R1878 B.n206 B.n205 163.367
R1879 B.n210 B.n209 163.367
R1880 B.n214 B.n213 163.367
R1881 B.n218 B.n217 163.367
R1882 B.n222 B.n221 163.367
R1883 B.n226 B.n225 163.367
R1884 B.n230 B.n229 163.367
R1885 B.n234 B.n233 163.367
R1886 B.n239 B.n238 163.367
R1887 B.n243 B.n242 163.367
R1888 B.n247 B.n246 163.367
R1889 B.n251 B.n250 163.367
R1890 B.n255 B.n254 163.367
R1891 B.n259 B.n258 163.367
R1892 B.n263 B.n262 163.367
R1893 B.n267 B.n266 163.367
R1894 B.n271 B.n270 163.367
R1895 B.n275 B.n274 163.367
R1896 B.n279 B.n278 163.367
R1897 B.n283 B.n282 163.367
R1898 B.n287 B.n286 163.367
R1899 B.n291 B.n290 163.367
R1900 B.n295 B.n294 163.367
R1901 B.n299 B.n298 163.367
R1902 B.n303 B.n302 163.367
R1903 B.n307 B.n306 163.367
R1904 B.n311 B.n310 163.367
R1905 B.n315 B.n314 163.367
R1906 B.n319 B.n318 163.367
R1907 B.n323 B.n322 163.367
R1908 B.n327 B.n326 163.367
R1909 B.n816 B.n119 163.367
R1910 B.n665 B.n664 71.676
R1911 B.n451 B.n400 71.676
R1912 B.n657 B.n401 71.676
R1913 B.n653 B.n402 71.676
R1914 B.n649 B.n403 71.676
R1915 B.n645 B.n404 71.676
R1916 B.n641 B.n405 71.676
R1917 B.n637 B.n406 71.676
R1918 B.n633 B.n407 71.676
R1919 B.n629 B.n408 71.676
R1920 B.n625 B.n409 71.676
R1921 B.n621 B.n410 71.676
R1922 B.n617 B.n411 71.676
R1923 B.n613 B.n412 71.676
R1924 B.n609 B.n413 71.676
R1925 B.n605 B.n414 71.676
R1926 B.n601 B.n415 71.676
R1927 B.n597 B.n416 71.676
R1928 B.n593 B.n417 71.676
R1929 B.n589 B.n418 71.676
R1930 B.n585 B.n419 71.676
R1931 B.n581 B.n420 71.676
R1932 B.n577 B.n421 71.676
R1933 B.n573 B.n422 71.676
R1934 B.n568 B.n423 71.676
R1935 B.n564 B.n424 71.676
R1936 B.n560 B.n425 71.676
R1937 B.n556 B.n426 71.676
R1938 B.n552 B.n427 71.676
R1939 B.n548 B.n428 71.676
R1940 B.n544 B.n429 71.676
R1941 B.n540 B.n430 71.676
R1942 B.n536 B.n431 71.676
R1943 B.n532 B.n432 71.676
R1944 B.n528 B.n433 71.676
R1945 B.n524 B.n434 71.676
R1946 B.n520 B.n435 71.676
R1947 B.n516 B.n436 71.676
R1948 B.n512 B.n437 71.676
R1949 B.n508 B.n438 71.676
R1950 B.n504 B.n439 71.676
R1951 B.n500 B.n440 71.676
R1952 B.n496 B.n441 71.676
R1953 B.n492 B.n442 71.676
R1954 B.n488 B.n443 71.676
R1955 B.n484 B.n444 71.676
R1956 B.n480 B.n445 71.676
R1957 B.n476 B.n446 71.676
R1958 B.n472 B.n447 71.676
R1959 B.n468 B.n448 71.676
R1960 B.n464 B.n449 71.676
R1961 B.n460 B.n450 71.676
R1962 B.n819 B.n818 71.676
R1963 B.n126 B.n68 71.676
R1964 B.n130 B.n69 71.676
R1965 B.n134 B.n70 71.676
R1966 B.n138 B.n71 71.676
R1967 B.n142 B.n72 71.676
R1968 B.n146 B.n73 71.676
R1969 B.n150 B.n74 71.676
R1970 B.n154 B.n75 71.676
R1971 B.n158 B.n76 71.676
R1972 B.n162 B.n77 71.676
R1973 B.n166 B.n78 71.676
R1974 B.n170 B.n79 71.676
R1975 B.n174 B.n80 71.676
R1976 B.n178 B.n81 71.676
R1977 B.n182 B.n82 71.676
R1978 B.n186 B.n83 71.676
R1979 B.n190 B.n84 71.676
R1980 B.n194 B.n85 71.676
R1981 B.n198 B.n86 71.676
R1982 B.n202 B.n87 71.676
R1983 B.n206 B.n88 71.676
R1984 B.n210 B.n89 71.676
R1985 B.n214 B.n90 71.676
R1986 B.n218 B.n91 71.676
R1987 B.n222 B.n92 71.676
R1988 B.n226 B.n93 71.676
R1989 B.n230 B.n94 71.676
R1990 B.n234 B.n95 71.676
R1991 B.n239 B.n96 71.676
R1992 B.n243 B.n97 71.676
R1993 B.n247 B.n98 71.676
R1994 B.n251 B.n99 71.676
R1995 B.n255 B.n100 71.676
R1996 B.n259 B.n101 71.676
R1997 B.n263 B.n102 71.676
R1998 B.n267 B.n103 71.676
R1999 B.n271 B.n104 71.676
R2000 B.n275 B.n105 71.676
R2001 B.n279 B.n106 71.676
R2002 B.n283 B.n107 71.676
R2003 B.n287 B.n108 71.676
R2004 B.n291 B.n109 71.676
R2005 B.n295 B.n110 71.676
R2006 B.n299 B.n111 71.676
R2007 B.n303 B.n112 71.676
R2008 B.n307 B.n113 71.676
R2009 B.n311 B.n114 71.676
R2010 B.n315 B.n115 71.676
R2011 B.n319 B.n116 71.676
R2012 B.n323 B.n117 71.676
R2013 B.n327 B.n118 71.676
R2014 B.n119 B.n118 71.676
R2015 B.n326 B.n117 71.676
R2016 B.n322 B.n116 71.676
R2017 B.n318 B.n115 71.676
R2018 B.n314 B.n114 71.676
R2019 B.n310 B.n113 71.676
R2020 B.n306 B.n112 71.676
R2021 B.n302 B.n111 71.676
R2022 B.n298 B.n110 71.676
R2023 B.n294 B.n109 71.676
R2024 B.n290 B.n108 71.676
R2025 B.n286 B.n107 71.676
R2026 B.n282 B.n106 71.676
R2027 B.n278 B.n105 71.676
R2028 B.n274 B.n104 71.676
R2029 B.n270 B.n103 71.676
R2030 B.n266 B.n102 71.676
R2031 B.n262 B.n101 71.676
R2032 B.n258 B.n100 71.676
R2033 B.n254 B.n99 71.676
R2034 B.n250 B.n98 71.676
R2035 B.n246 B.n97 71.676
R2036 B.n242 B.n96 71.676
R2037 B.n238 B.n95 71.676
R2038 B.n233 B.n94 71.676
R2039 B.n229 B.n93 71.676
R2040 B.n225 B.n92 71.676
R2041 B.n221 B.n91 71.676
R2042 B.n217 B.n90 71.676
R2043 B.n213 B.n89 71.676
R2044 B.n209 B.n88 71.676
R2045 B.n205 B.n87 71.676
R2046 B.n201 B.n86 71.676
R2047 B.n197 B.n85 71.676
R2048 B.n193 B.n84 71.676
R2049 B.n189 B.n83 71.676
R2050 B.n185 B.n82 71.676
R2051 B.n181 B.n81 71.676
R2052 B.n177 B.n80 71.676
R2053 B.n173 B.n79 71.676
R2054 B.n169 B.n78 71.676
R2055 B.n165 B.n77 71.676
R2056 B.n161 B.n76 71.676
R2057 B.n157 B.n75 71.676
R2058 B.n153 B.n74 71.676
R2059 B.n149 B.n73 71.676
R2060 B.n145 B.n72 71.676
R2061 B.n141 B.n71 71.676
R2062 B.n137 B.n70 71.676
R2063 B.n133 B.n69 71.676
R2064 B.n129 B.n68 71.676
R2065 B.n818 B.n67 71.676
R2066 B.n664 B.n399 71.676
R2067 B.n658 B.n400 71.676
R2068 B.n654 B.n401 71.676
R2069 B.n650 B.n402 71.676
R2070 B.n646 B.n403 71.676
R2071 B.n642 B.n404 71.676
R2072 B.n638 B.n405 71.676
R2073 B.n634 B.n406 71.676
R2074 B.n630 B.n407 71.676
R2075 B.n626 B.n408 71.676
R2076 B.n622 B.n409 71.676
R2077 B.n618 B.n410 71.676
R2078 B.n614 B.n411 71.676
R2079 B.n610 B.n412 71.676
R2080 B.n606 B.n413 71.676
R2081 B.n602 B.n414 71.676
R2082 B.n598 B.n415 71.676
R2083 B.n594 B.n416 71.676
R2084 B.n590 B.n417 71.676
R2085 B.n586 B.n418 71.676
R2086 B.n582 B.n419 71.676
R2087 B.n578 B.n420 71.676
R2088 B.n574 B.n421 71.676
R2089 B.n569 B.n422 71.676
R2090 B.n565 B.n423 71.676
R2091 B.n561 B.n424 71.676
R2092 B.n557 B.n425 71.676
R2093 B.n553 B.n426 71.676
R2094 B.n549 B.n427 71.676
R2095 B.n545 B.n428 71.676
R2096 B.n541 B.n429 71.676
R2097 B.n537 B.n430 71.676
R2098 B.n533 B.n431 71.676
R2099 B.n529 B.n432 71.676
R2100 B.n525 B.n433 71.676
R2101 B.n521 B.n434 71.676
R2102 B.n517 B.n435 71.676
R2103 B.n513 B.n436 71.676
R2104 B.n509 B.n437 71.676
R2105 B.n505 B.n438 71.676
R2106 B.n501 B.n439 71.676
R2107 B.n497 B.n440 71.676
R2108 B.n493 B.n441 71.676
R2109 B.n489 B.n442 71.676
R2110 B.n485 B.n443 71.676
R2111 B.n481 B.n444 71.676
R2112 B.n477 B.n445 71.676
R2113 B.n473 B.n446 71.676
R2114 B.n469 B.n447 71.676
R2115 B.n465 B.n448 71.676
R2116 B.n461 B.n449 71.676
R2117 B.n457 B.n450 71.676
R2118 B.n663 B.n396 71.2625
R2119 B.n817 B.n64 71.2625
R2120 B.n456 B.n455 59.5399
R2121 B.n571 B.n453 59.5399
R2122 B.n125 B.n124 59.5399
R2123 B.n236 B.n122 59.5399
R2124 B.n670 B.n396 38.767
R2125 B.n670 B.n392 38.767
R2126 B.n676 B.n392 38.767
R2127 B.n676 B.n388 38.767
R2128 B.n682 B.n388 38.767
R2129 B.n688 B.n384 38.767
R2130 B.n688 B.n380 38.767
R2131 B.n694 B.n380 38.767
R2132 B.n694 B.n376 38.767
R2133 B.n700 B.n376 38.767
R2134 B.n700 B.n371 38.767
R2135 B.n706 B.n371 38.767
R2136 B.n706 B.n372 38.767
R2137 B.n712 B.n364 38.767
R2138 B.n718 B.n364 38.767
R2139 B.n718 B.n360 38.767
R2140 B.n724 B.n360 38.767
R2141 B.n730 B.n356 38.767
R2142 B.n730 B.n352 38.767
R2143 B.n736 B.n352 38.767
R2144 B.n736 B.n348 38.767
R2145 B.n742 B.n348 38.767
R2146 B.n748 B.n344 38.767
R2147 B.n748 B.n339 38.767
R2148 B.n754 B.n339 38.767
R2149 B.n754 B.n340 38.767
R2150 B.n761 B.n332 38.767
R2151 B.n767 B.n332 38.767
R2152 B.n767 B.n4 38.767
R2153 B.n890 B.n4 38.767
R2154 B.n890 B.n889 38.767
R2155 B.n889 B.n888 38.767
R2156 B.n888 B.n8 38.767
R2157 B.n882 B.n8 38.767
R2158 B.n881 B.n880 38.767
R2159 B.n880 B.n15 38.767
R2160 B.n874 B.n15 38.767
R2161 B.n874 B.n873 38.767
R2162 B.n872 B.n22 38.767
R2163 B.n866 B.n22 38.767
R2164 B.n866 B.n865 38.767
R2165 B.n865 B.n864 38.767
R2166 B.n864 B.n29 38.767
R2167 B.n858 B.n857 38.767
R2168 B.n857 B.n856 38.767
R2169 B.n856 B.n36 38.767
R2170 B.n850 B.n36 38.767
R2171 B.n849 B.n848 38.767
R2172 B.n848 B.n43 38.767
R2173 B.n842 B.n43 38.767
R2174 B.n842 B.n841 38.767
R2175 B.n841 B.n840 38.767
R2176 B.n840 B.n50 38.767
R2177 B.n834 B.n50 38.767
R2178 B.n834 B.n833 38.767
R2179 B.n832 B.n57 38.767
R2180 B.n826 B.n57 38.767
R2181 B.n826 B.n825 38.767
R2182 B.n825 B.n824 38.767
R2183 B.n824 B.n64 38.767
R2184 B.n682 B.t9 37.6268
R2185 B.t13 B.n832 37.6268
R2186 B.n724 B.t5 36.4866
R2187 B.n858 B.t7 36.4866
R2188 B.n455 B.n454 35.4914
R2189 B.n453 B.n452 35.4914
R2190 B.n124 B.n123 35.4914
R2191 B.n122 B.n121 35.4914
R2192 B.n821 B.n820 31.0639
R2193 B.n815 B.n814 31.0639
R2194 B.n458 B.n394 31.0639
R2195 B.n667 B.n666 31.0639
R2196 B.n340 B.t0 27.3651
R2197 B.t1 B.n881 27.3651
R2198 B.t2 B.n344 26.2249
R2199 B.n873 B.t4 26.2249
R2200 B.n372 B.t3 21.6641
R2201 B.t6 B.n849 21.6641
R2202 B B.n892 18.0485
R2203 B.n712 B.t3 17.1034
R2204 B.n850 B.t6 17.1034
R2205 B.n742 B.t2 12.5426
R2206 B.t4 B.n872 12.5426
R2207 B.n761 B.t0 11.4024
R2208 B.n882 B.t1 11.4024
R2209 B.n820 B.n66 10.6151
R2210 B.n127 B.n66 10.6151
R2211 B.n128 B.n127 10.6151
R2212 B.n131 B.n128 10.6151
R2213 B.n132 B.n131 10.6151
R2214 B.n135 B.n132 10.6151
R2215 B.n136 B.n135 10.6151
R2216 B.n139 B.n136 10.6151
R2217 B.n140 B.n139 10.6151
R2218 B.n143 B.n140 10.6151
R2219 B.n144 B.n143 10.6151
R2220 B.n147 B.n144 10.6151
R2221 B.n148 B.n147 10.6151
R2222 B.n151 B.n148 10.6151
R2223 B.n152 B.n151 10.6151
R2224 B.n155 B.n152 10.6151
R2225 B.n156 B.n155 10.6151
R2226 B.n159 B.n156 10.6151
R2227 B.n160 B.n159 10.6151
R2228 B.n163 B.n160 10.6151
R2229 B.n164 B.n163 10.6151
R2230 B.n167 B.n164 10.6151
R2231 B.n168 B.n167 10.6151
R2232 B.n171 B.n168 10.6151
R2233 B.n172 B.n171 10.6151
R2234 B.n175 B.n172 10.6151
R2235 B.n176 B.n175 10.6151
R2236 B.n179 B.n176 10.6151
R2237 B.n180 B.n179 10.6151
R2238 B.n183 B.n180 10.6151
R2239 B.n184 B.n183 10.6151
R2240 B.n187 B.n184 10.6151
R2241 B.n188 B.n187 10.6151
R2242 B.n191 B.n188 10.6151
R2243 B.n192 B.n191 10.6151
R2244 B.n195 B.n192 10.6151
R2245 B.n196 B.n195 10.6151
R2246 B.n199 B.n196 10.6151
R2247 B.n200 B.n199 10.6151
R2248 B.n203 B.n200 10.6151
R2249 B.n204 B.n203 10.6151
R2250 B.n207 B.n204 10.6151
R2251 B.n208 B.n207 10.6151
R2252 B.n211 B.n208 10.6151
R2253 B.n212 B.n211 10.6151
R2254 B.n215 B.n212 10.6151
R2255 B.n216 B.n215 10.6151
R2256 B.n220 B.n219 10.6151
R2257 B.n223 B.n220 10.6151
R2258 B.n224 B.n223 10.6151
R2259 B.n227 B.n224 10.6151
R2260 B.n228 B.n227 10.6151
R2261 B.n231 B.n228 10.6151
R2262 B.n232 B.n231 10.6151
R2263 B.n235 B.n232 10.6151
R2264 B.n240 B.n237 10.6151
R2265 B.n241 B.n240 10.6151
R2266 B.n244 B.n241 10.6151
R2267 B.n245 B.n244 10.6151
R2268 B.n248 B.n245 10.6151
R2269 B.n249 B.n248 10.6151
R2270 B.n252 B.n249 10.6151
R2271 B.n253 B.n252 10.6151
R2272 B.n256 B.n253 10.6151
R2273 B.n257 B.n256 10.6151
R2274 B.n260 B.n257 10.6151
R2275 B.n261 B.n260 10.6151
R2276 B.n264 B.n261 10.6151
R2277 B.n265 B.n264 10.6151
R2278 B.n268 B.n265 10.6151
R2279 B.n269 B.n268 10.6151
R2280 B.n272 B.n269 10.6151
R2281 B.n273 B.n272 10.6151
R2282 B.n276 B.n273 10.6151
R2283 B.n277 B.n276 10.6151
R2284 B.n280 B.n277 10.6151
R2285 B.n281 B.n280 10.6151
R2286 B.n284 B.n281 10.6151
R2287 B.n285 B.n284 10.6151
R2288 B.n288 B.n285 10.6151
R2289 B.n289 B.n288 10.6151
R2290 B.n292 B.n289 10.6151
R2291 B.n293 B.n292 10.6151
R2292 B.n296 B.n293 10.6151
R2293 B.n297 B.n296 10.6151
R2294 B.n300 B.n297 10.6151
R2295 B.n301 B.n300 10.6151
R2296 B.n304 B.n301 10.6151
R2297 B.n305 B.n304 10.6151
R2298 B.n308 B.n305 10.6151
R2299 B.n309 B.n308 10.6151
R2300 B.n312 B.n309 10.6151
R2301 B.n313 B.n312 10.6151
R2302 B.n316 B.n313 10.6151
R2303 B.n317 B.n316 10.6151
R2304 B.n320 B.n317 10.6151
R2305 B.n321 B.n320 10.6151
R2306 B.n324 B.n321 10.6151
R2307 B.n325 B.n324 10.6151
R2308 B.n328 B.n325 10.6151
R2309 B.n329 B.n328 10.6151
R2310 B.n815 B.n329 10.6151
R2311 B.n672 B.n394 10.6151
R2312 B.n673 B.n672 10.6151
R2313 B.n674 B.n673 10.6151
R2314 B.n674 B.n386 10.6151
R2315 B.n684 B.n386 10.6151
R2316 B.n685 B.n684 10.6151
R2317 B.n686 B.n685 10.6151
R2318 B.n686 B.n378 10.6151
R2319 B.n696 B.n378 10.6151
R2320 B.n697 B.n696 10.6151
R2321 B.n698 B.n697 10.6151
R2322 B.n698 B.n369 10.6151
R2323 B.n708 B.n369 10.6151
R2324 B.n709 B.n708 10.6151
R2325 B.n710 B.n709 10.6151
R2326 B.n710 B.n362 10.6151
R2327 B.n720 B.n362 10.6151
R2328 B.n721 B.n720 10.6151
R2329 B.n722 B.n721 10.6151
R2330 B.n722 B.n354 10.6151
R2331 B.n732 B.n354 10.6151
R2332 B.n733 B.n732 10.6151
R2333 B.n734 B.n733 10.6151
R2334 B.n734 B.n346 10.6151
R2335 B.n744 B.n346 10.6151
R2336 B.n745 B.n744 10.6151
R2337 B.n746 B.n745 10.6151
R2338 B.n746 B.n337 10.6151
R2339 B.n756 B.n337 10.6151
R2340 B.n757 B.n756 10.6151
R2341 B.n759 B.n757 10.6151
R2342 B.n759 B.n758 10.6151
R2343 B.n758 B.n330 10.6151
R2344 B.n770 B.n330 10.6151
R2345 B.n771 B.n770 10.6151
R2346 B.n772 B.n771 10.6151
R2347 B.n773 B.n772 10.6151
R2348 B.n775 B.n773 10.6151
R2349 B.n776 B.n775 10.6151
R2350 B.n777 B.n776 10.6151
R2351 B.n778 B.n777 10.6151
R2352 B.n780 B.n778 10.6151
R2353 B.n781 B.n780 10.6151
R2354 B.n782 B.n781 10.6151
R2355 B.n783 B.n782 10.6151
R2356 B.n785 B.n783 10.6151
R2357 B.n786 B.n785 10.6151
R2358 B.n787 B.n786 10.6151
R2359 B.n788 B.n787 10.6151
R2360 B.n790 B.n788 10.6151
R2361 B.n791 B.n790 10.6151
R2362 B.n792 B.n791 10.6151
R2363 B.n793 B.n792 10.6151
R2364 B.n795 B.n793 10.6151
R2365 B.n796 B.n795 10.6151
R2366 B.n797 B.n796 10.6151
R2367 B.n798 B.n797 10.6151
R2368 B.n800 B.n798 10.6151
R2369 B.n801 B.n800 10.6151
R2370 B.n802 B.n801 10.6151
R2371 B.n803 B.n802 10.6151
R2372 B.n805 B.n803 10.6151
R2373 B.n806 B.n805 10.6151
R2374 B.n807 B.n806 10.6151
R2375 B.n808 B.n807 10.6151
R2376 B.n810 B.n808 10.6151
R2377 B.n811 B.n810 10.6151
R2378 B.n812 B.n811 10.6151
R2379 B.n813 B.n812 10.6151
R2380 B.n814 B.n813 10.6151
R2381 B.n666 B.n398 10.6151
R2382 B.n661 B.n398 10.6151
R2383 B.n661 B.n660 10.6151
R2384 B.n660 B.n659 10.6151
R2385 B.n659 B.n656 10.6151
R2386 B.n656 B.n655 10.6151
R2387 B.n655 B.n652 10.6151
R2388 B.n652 B.n651 10.6151
R2389 B.n651 B.n648 10.6151
R2390 B.n648 B.n647 10.6151
R2391 B.n647 B.n644 10.6151
R2392 B.n644 B.n643 10.6151
R2393 B.n643 B.n640 10.6151
R2394 B.n640 B.n639 10.6151
R2395 B.n639 B.n636 10.6151
R2396 B.n636 B.n635 10.6151
R2397 B.n635 B.n632 10.6151
R2398 B.n632 B.n631 10.6151
R2399 B.n631 B.n628 10.6151
R2400 B.n628 B.n627 10.6151
R2401 B.n627 B.n624 10.6151
R2402 B.n624 B.n623 10.6151
R2403 B.n623 B.n620 10.6151
R2404 B.n620 B.n619 10.6151
R2405 B.n619 B.n616 10.6151
R2406 B.n616 B.n615 10.6151
R2407 B.n615 B.n612 10.6151
R2408 B.n612 B.n611 10.6151
R2409 B.n611 B.n608 10.6151
R2410 B.n608 B.n607 10.6151
R2411 B.n607 B.n604 10.6151
R2412 B.n604 B.n603 10.6151
R2413 B.n603 B.n600 10.6151
R2414 B.n600 B.n599 10.6151
R2415 B.n599 B.n596 10.6151
R2416 B.n596 B.n595 10.6151
R2417 B.n595 B.n592 10.6151
R2418 B.n592 B.n591 10.6151
R2419 B.n591 B.n588 10.6151
R2420 B.n588 B.n587 10.6151
R2421 B.n587 B.n584 10.6151
R2422 B.n584 B.n583 10.6151
R2423 B.n583 B.n580 10.6151
R2424 B.n580 B.n579 10.6151
R2425 B.n579 B.n576 10.6151
R2426 B.n576 B.n575 10.6151
R2427 B.n575 B.n572 10.6151
R2428 B.n570 B.n567 10.6151
R2429 B.n567 B.n566 10.6151
R2430 B.n566 B.n563 10.6151
R2431 B.n563 B.n562 10.6151
R2432 B.n562 B.n559 10.6151
R2433 B.n559 B.n558 10.6151
R2434 B.n558 B.n555 10.6151
R2435 B.n555 B.n554 10.6151
R2436 B.n551 B.n550 10.6151
R2437 B.n550 B.n547 10.6151
R2438 B.n547 B.n546 10.6151
R2439 B.n546 B.n543 10.6151
R2440 B.n543 B.n542 10.6151
R2441 B.n542 B.n539 10.6151
R2442 B.n539 B.n538 10.6151
R2443 B.n538 B.n535 10.6151
R2444 B.n535 B.n534 10.6151
R2445 B.n534 B.n531 10.6151
R2446 B.n531 B.n530 10.6151
R2447 B.n530 B.n527 10.6151
R2448 B.n527 B.n526 10.6151
R2449 B.n526 B.n523 10.6151
R2450 B.n523 B.n522 10.6151
R2451 B.n522 B.n519 10.6151
R2452 B.n519 B.n518 10.6151
R2453 B.n518 B.n515 10.6151
R2454 B.n515 B.n514 10.6151
R2455 B.n514 B.n511 10.6151
R2456 B.n511 B.n510 10.6151
R2457 B.n510 B.n507 10.6151
R2458 B.n507 B.n506 10.6151
R2459 B.n506 B.n503 10.6151
R2460 B.n503 B.n502 10.6151
R2461 B.n502 B.n499 10.6151
R2462 B.n499 B.n498 10.6151
R2463 B.n498 B.n495 10.6151
R2464 B.n495 B.n494 10.6151
R2465 B.n494 B.n491 10.6151
R2466 B.n491 B.n490 10.6151
R2467 B.n490 B.n487 10.6151
R2468 B.n487 B.n486 10.6151
R2469 B.n486 B.n483 10.6151
R2470 B.n483 B.n482 10.6151
R2471 B.n482 B.n479 10.6151
R2472 B.n479 B.n478 10.6151
R2473 B.n478 B.n475 10.6151
R2474 B.n475 B.n474 10.6151
R2475 B.n474 B.n471 10.6151
R2476 B.n471 B.n470 10.6151
R2477 B.n470 B.n467 10.6151
R2478 B.n467 B.n466 10.6151
R2479 B.n466 B.n463 10.6151
R2480 B.n463 B.n462 10.6151
R2481 B.n462 B.n459 10.6151
R2482 B.n459 B.n458 10.6151
R2483 B.n668 B.n667 10.6151
R2484 B.n668 B.n390 10.6151
R2485 B.n678 B.n390 10.6151
R2486 B.n679 B.n678 10.6151
R2487 B.n680 B.n679 10.6151
R2488 B.n680 B.n382 10.6151
R2489 B.n690 B.n382 10.6151
R2490 B.n691 B.n690 10.6151
R2491 B.n692 B.n691 10.6151
R2492 B.n692 B.n374 10.6151
R2493 B.n702 B.n374 10.6151
R2494 B.n703 B.n702 10.6151
R2495 B.n704 B.n703 10.6151
R2496 B.n704 B.n366 10.6151
R2497 B.n714 B.n366 10.6151
R2498 B.n715 B.n714 10.6151
R2499 B.n716 B.n715 10.6151
R2500 B.n716 B.n358 10.6151
R2501 B.n726 B.n358 10.6151
R2502 B.n727 B.n726 10.6151
R2503 B.n728 B.n727 10.6151
R2504 B.n728 B.n350 10.6151
R2505 B.n738 B.n350 10.6151
R2506 B.n739 B.n738 10.6151
R2507 B.n740 B.n739 10.6151
R2508 B.n740 B.n342 10.6151
R2509 B.n750 B.n342 10.6151
R2510 B.n751 B.n750 10.6151
R2511 B.n752 B.n751 10.6151
R2512 B.n752 B.n334 10.6151
R2513 B.n763 B.n334 10.6151
R2514 B.n764 B.n763 10.6151
R2515 B.n765 B.n764 10.6151
R2516 B.n765 B.n0 10.6151
R2517 B.n886 B.n1 10.6151
R2518 B.n886 B.n885 10.6151
R2519 B.n885 B.n884 10.6151
R2520 B.n884 B.n10 10.6151
R2521 B.n878 B.n10 10.6151
R2522 B.n878 B.n877 10.6151
R2523 B.n877 B.n876 10.6151
R2524 B.n876 B.n17 10.6151
R2525 B.n870 B.n17 10.6151
R2526 B.n870 B.n869 10.6151
R2527 B.n869 B.n868 10.6151
R2528 B.n868 B.n24 10.6151
R2529 B.n862 B.n24 10.6151
R2530 B.n862 B.n861 10.6151
R2531 B.n861 B.n860 10.6151
R2532 B.n860 B.n31 10.6151
R2533 B.n854 B.n31 10.6151
R2534 B.n854 B.n853 10.6151
R2535 B.n853 B.n852 10.6151
R2536 B.n852 B.n38 10.6151
R2537 B.n846 B.n38 10.6151
R2538 B.n846 B.n845 10.6151
R2539 B.n845 B.n844 10.6151
R2540 B.n844 B.n45 10.6151
R2541 B.n838 B.n45 10.6151
R2542 B.n838 B.n837 10.6151
R2543 B.n837 B.n836 10.6151
R2544 B.n836 B.n52 10.6151
R2545 B.n830 B.n52 10.6151
R2546 B.n830 B.n829 10.6151
R2547 B.n829 B.n828 10.6151
R2548 B.n828 B.n59 10.6151
R2549 B.n822 B.n59 10.6151
R2550 B.n822 B.n821 10.6151
R2551 B.n219 B.n125 6.5566
R2552 B.n236 B.n235 6.5566
R2553 B.n571 B.n570 6.5566
R2554 B.n554 B.n456 6.5566
R2555 B.n216 B.n125 4.05904
R2556 B.n237 B.n236 4.05904
R2557 B.n572 B.n571 4.05904
R2558 B.n551 B.n456 4.05904
R2559 B.n892 B.n0 2.81026
R2560 B.n892 B.n1 2.81026
R2561 B.t5 B.n356 2.28088
R2562 B.t7 B.n29 2.28088
R2563 B.t9 B.n384 1.14069
R2564 B.n833 B.t13 1.14069
R2565 VN.n5 VN.t2 260.092
R2566 VN.n24 VN.t5 260.092
R2567 VN.n4 VN.t6 225.256
R2568 VN.n10 VN.t3 225.256
R2569 VN.n17 VN.t7 225.256
R2570 VN.n23 VN.t4 225.256
R2571 VN.n29 VN.t1 225.256
R2572 VN.n36 VN.t0 225.256
R2573 VN.n18 VN.n17 173.843
R2574 VN.n37 VN.n36 173.843
R2575 VN.n35 VN.n19 161.3
R2576 VN.n34 VN.n33 161.3
R2577 VN.n32 VN.n20 161.3
R2578 VN.n31 VN.n30 161.3
R2579 VN.n28 VN.n21 161.3
R2580 VN.n27 VN.n26 161.3
R2581 VN.n25 VN.n22 161.3
R2582 VN.n16 VN.n0 161.3
R2583 VN.n15 VN.n14 161.3
R2584 VN.n13 VN.n1 161.3
R2585 VN.n12 VN.n11 161.3
R2586 VN.n9 VN.n2 161.3
R2587 VN.n8 VN.n7 161.3
R2588 VN.n6 VN.n3 161.3
R2589 VN.n15 VN.n1 56.5617
R2590 VN.n34 VN.n20 56.5617
R2591 VN VN.n37 47.616
R2592 VN.n5 VN.n4 46.3697
R2593 VN.n24 VN.n23 46.3697
R2594 VN.n8 VN.n3 40.577
R2595 VN.n9 VN.n8 40.577
R2596 VN.n27 VN.n22 40.577
R2597 VN.n28 VN.n27 40.577
R2598 VN.n11 VN.n1 24.5923
R2599 VN.n16 VN.n15 24.5923
R2600 VN.n30 VN.n20 24.5923
R2601 VN.n35 VN.n34 24.5923
R2602 VN.n4 VN.n3 20.4117
R2603 VN.n10 VN.n9 20.4117
R2604 VN.n23 VN.n22 20.4117
R2605 VN.n29 VN.n28 20.4117
R2606 VN.n25 VN.n24 17.5628
R2607 VN.n6 VN.n5 17.5628
R2608 VN.n17 VN.n16 12.0505
R2609 VN.n36 VN.n35 12.0505
R2610 VN.n11 VN.n10 4.18111
R2611 VN.n30 VN.n29 4.18111
R2612 VN.n37 VN.n19 0.189894
R2613 VN.n33 VN.n19 0.189894
R2614 VN.n33 VN.n32 0.189894
R2615 VN.n32 VN.n31 0.189894
R2616 VN.n31 VN.n21 0.189894
R2617 VN.n26 VN.n21 0.189894
R2618 VN.n26 VN.n25 0.189894
R2619 VN.n7 VN.n6 0.189894
R2620 VN.n7 VN.n2 0.189894
R2621 VN.n12 VN.n2 0.189894
R2622 VN.n13 VN.n12 0.189894
R2623 VN.n14 VN.n13 0.189894
R2624 VN.n14 VN.n0 0.189894
R2625 VN.n18 VN.n0 0.189894
R2626 VN VN.n18 0.0516364
R2627 VDD2.n2 VDD2.n1 63.6871
R2628 VDD2.n2 VDD2.n0 63.6871
R2629 VDD2 VDD2.n5 63.6842
R2630 VDD2.n4 VDD2.n3 62.9538
R2631 VDD2.n4 VDD2.n2 42.9006
R2632 VDD2.n5 VDD2.t3 1.41277
R2633 VDD2.n5 VDD2.t2 1.41277
R2634 VDD2.n3 VDD2.t7 1.41277
R2635 VDD2.n3 VDD2.t6 1.41277
R2636 VDD2.n1 VDD2.t4 1.41277
R2637 VDD2.n1 VDD2.t0 1.41277
R2638 VDD2.n0 VDD2.t5 1.41277
R2639 VDD2.n0 VDD2.t1 1.41277
R2640 VDD2 VDD2.n4 0.847483
C0 VDD1 VP 9.015161f
C1 VDD2 VP 0.40302f
C2 VTAIL VP 8.74612f
C3 VN VP 6.68545f
C4 VDD1 VDD2 1.22323f
C5 VTAIL VDD1 9.405981f
C6 VTAIL VDD2 9.45302f
C7 VN VDD1 0.15014f
C8 VN VDD2 8.76312f
C9 VN VTAIL 8.73201f
C10 VDD2 B 4.427595f
C11 VDD1 B 4.743109f
C12 VTAIL B 10.817836f
C13 VN B 11.56756f
C14 VP B 9.893922f
C15 VDD2.t5 B 0.278273f
C16 VDD2.t1 B 0.278273f
C17 VDD2.n0 B 2.51391f
C18 VDD2.t4 B 0.278273f
C19 VDD2.t0 B 0.278273f
C20 VDD2.n1 B 2.51391f
C21 VDD2.n2 B 2.76876f
C22 VDD2.t7 B 0.278273f
C23 VDD2.t6 B 0.278273f
C24 VDD2.n3 B 2.50931f
C25 VDD2.n4 B 2.73159f
C26 VDD2.t3 B 0.278273f
C27 VDD2.t2 B 0.278273f
C28 VDD2.n5 B 2.51388f
C29 VN.n0 B 0.030598f
C30 VN.t7 B 1.76046f
C31 VN.n1 B 0.051252f
C32 VN.n2 B 0.030598f
C33 VN.t3 B 1.76046f
C34 VN.n3 B 0.055731f
C35 VN.t2 B 1.86067f
C36 VN.t6 B 1.76046f
C37 VN.n4 B 0.695376f
C38 VN.n5 B 0.696311f
C39 VN.n6 B 0.194552f
C40 VN.n7 B 0.030598f
C41 VN.n8 B 0.024713f
C42 VN.n9 B 0.055731f
C43 VN.n10 B 0.629122f
C44 VN.n11 B 0.033492f
C45 VN.n12 B 0.030598f
C46 VN.n13 B 0.030598f
C47 VN.n14 B 0.030598f
C48 VN.n15 B 0.037707f
C49 VN.n16 B 0.042456f
C50 VN.n17 B 0.694506f
C51 VN.n18 B 0.028796f
C52 VN.n19 B 0.030598f
C53 VN.t0 B 1.76046f
C54 VN.n20 B 0.051252f
C55 VN.n21 B 0.030598f
C56 VN.t1 B 1.76046f
C57 VN.n22 B 0.055731f
C58 VN.t5 B 1.86067f
C59 VN.t4 B 1.76046f
C60 VN.n23 B 0.695376f
C61 VN.n24 B 0.696311f
C62 VN.n25 B 0.194552f
C63 VN.n26 B 0.030598f
C64 VN.n27 B 0.024713f
C65 VN.n28 B 0.055731f
C66 VN.n29 B 0.629122f
C67 VN.n30 B 0.033492f
C68 VN.n31 B 0.030598f
C69 VN.n32 B 0.030598f
C70 VN.n33 B 0.030598f
C71 VN.n34 B 0.037707f
C72 VN.n35 B 0.042456f
C73 VN.n36 B 0.694506f
C74 VN.n37 B 1.55019f
C75 VTAIL.t4 B 0.208654f
C76 VTAIL.t7 B 0.208654f
C77 VTAIL.n0 B 1.82811f
C78 VTAIL.n1 B 0.278863f
C79 VTAIL.n2 B 0.024693f
C80 VTAIL.n3 B 0.018833f
C81 VTAIL.n4 B 0.010418f
C82 VTAIL.n5 B 0.02392f
C83 VTAIL.n6 B 0.010715f
C84 VTAIL.n7 B 0.018833f
C85 VTAIL.n8 B 0.01012f
C86 VTAIL.n9 B 0.02392f
C87 VTAIL.n10 B 0.010715f
C88 VTAIL.n11 B 0.018833f
C89 VTAIL.n12 B 0.01012f
C90 VTAIL.n13 B 0.02392f
C91 VTAIL.n14 B 0.010715f
C92 VTAIL.n15 B 0.018833f
C93 VTAIL.n16 B 0.01012f
C94 VTAIL.n17 B 0.02392f
C95 VTAIL.n18 B 0.010715f
C96 VTAIL.n19 B 0.018833f
C97 VTAIL.n20 B 0.01012f
C98 VTAIL.n21 B 0.02392f
C99 VTAIL.n22 B 0.010715f
C100 VTAIL.n23 B 0.018833f
C101 VTAIL.n24 B 0.01012f
C102 VTAIL.n25 B 0.01794f
C103 VTAIL.n26 B 0.014131f
C104 VTAIL.t1 B 0.039379f
C105 VTAIL.n27 B 0.118207f
C106 VTAIL.n28 B 1.14073f
C107 VTAIL.n29 B 0.01012f
C108 VTAIL.n30 B 0.010715f
C109 VTAIL.n31 B 0.02392f
C110 VTAIL.n32 B 0.02392f
C111 VTAIL.n33 B 0.010715f
C112 VTAIL.n34 B 0.01012f
C113 VTAIL.n35 B 0.018833f
C114 VTAIL.n36 B 0.018833f
C115 VTAIL.n37 B 0.01012f
C116 VTAIL.n38 B 0.010715f
C117 VTAIL.n39 B 0.02392f
C118 VTAIL.n40 B 0.02392f
C119 VTAIL.n41 B 0.010715f
C120 VTAIL.n42 B 0.01012f
C121 VTAIL.n43 B 0.018833f
C122 VTAIL.n44 B 0.018833f
C123 VTAIL.n45 B 0.01012f
C124 VTAIL.n46 B 0.010715f
C125 VTAIL.n47 B 0.02392f
C126 VTAIL.n48 B 0.02392f
C127 VTAIL.n49 B 0.010715f
C128 VTAIL.n50 B 0.01012f
C129 VTAIL.n51 B 0.018833f
C130 VTAIL.n52 B 0.018833f
C131 VTAIL.n53 B 0.01012f
C132 VTAIL.n54 B 0.010715f
C133 VTAIL.n55 B 0.02392f
C134 VTAIL.n56 B 0.02392f
C135 VTAIL.n57 B 0.010715f
C136 VTAIL.n58 B 0.01012f
C137 VTAIL.n59 B 0.018833f
C138 VTAIL.n60 B 0.018833f
C139 VTAIL.n61 B 0.01012f
C140 VTAIL.n62 B 0.010715f
C141 VTAIL.n63 B 0.02392f
C142 VTAIL.n64 B 0.02392f
C143 VTAIL.n65 B 0.010715f
C144 VTAIL.n66 B 0.01012f
C145 VTAIL.n67 B 0.018833f
C146 VTAIL.n68 B 0.018833f
C147 VTAIL.n69 B 0.01012f
C148 VTAIL.n70 B 0.01012f
C149 VTAIL.n71 B 0.010715f
C150 VTAIL.n72 B 0.02392f
C151 VTAIL.n73 B 0.02392f
C152 VTAIL.n74 B 0.048638f
C153 VTAIL.n75 B 0.010418f
C154 VTAIL.n76 B 0.01012f
C155 VTAIL.n77 B 0.046105f
C156 VTAIL.n78 B 0.026968f
C157 VTAIL.n79 B 0.141786f
C158 VTAIL.n80 B 0.024693f
C159 VTAIL.n81 B 0.018833f
C160 VTAIL.n82 B 0.010418f
C161 VTAIL.n83 B 0.02392f
C162 VTAIL.n84 B 0.010715f
C163 VTAIL.n85 B 0.018833f
C164 VTAIL.n86 B 0.01012f
C165 VTAIL.n87 B 0.02392f
C166 VTAIL.n88 B 0.010715f
C167 VTAIL.n89 B 0.018833f
C168 VTAIL.n90 B 0.01012f
C169 VTAIL.n91 B 0.02392f
C170 VTAIL.n92 B 0.010715f
C171 VTAIL.n93 B 0.018833f
C172 VTAIL.n94 B 0.01012f
C173 VTAIL.n95 B 0.02392f
C174 VTAIL.n96 B 0.010715f
C175 VTAIL.n97 B 0.018833f
C176 VTAIL.n98 B 0.01012f
C177 VTAIL.n99 B 0.02392f
C178 VTAIL.n100 B 0.010715f
C179 VTAIL.n101 B 0.018833f
C180 VTAIL.n102 B 0.01012f
C181 VTAIL.n103 B 0.01794f
C182 VTAIL.n104 B 0.014131f
C183 VTAIL.t14 B 0.039379f
C184 VTAIL.n105 B 0.118207f
C185 VTAIL.n106 B 1.14073f
C186 VTAIL.n107 B 0.01012f
C187 VTAIL.n108 B 0.010715f
C188 VTAIL.n109 B 0.02392f
C189 VTAIL.n110 B 0.02392f
C190 VTAIL.n111 B 0.010715f
C191 VTAIL.n112 B 0.01012f
C192 VTAIL.n113 B 0.018833f
C193 VTAIL.n114 B 0.018833f
C194 VTAIL.n115 B 0.01012f
C195 VTAIL.n116 B 0.010715f
C196 VTAIL.n117 B 0.02392f
C197 VTAIL.n118 B 0.02392f
C198 VTAIL.n119 B 0.010715f
C199 VTAIL.n120 B 0.01012f
C200 VTAIL.n121 B 0.018833f
C201 VTAIL.n122 B 0.018833f
C202 VTAIL.n123 B 0.01012f
C203 VTAIL.n124 B 0.010715f
C204 VTAIL.n125 B 0.02392f
C205 VTAIL.n126 B 0.02392f
C206 VTAIL.n127 B 0.010715f
C207 VTAIL.n128 B 0.01012f
C208 VTAIL.n129 B 0.018833f
C209 VTAIL.n130 B 0.018833f
C210 VTAIL.n131 B 0.01012f
C211 VTAIL.n132 B 0.010715f
C212 VTAIL.n133 B 0.02392f
C213 VTAIL.n134 B 0.02392f
C214 VTAIL.n135 B 0.010715f
C215 VTAIL.n136 B 0.01012f
C216 VTAIL.n137 B 0.018833f
C217 VTAIL.n138 B 0.018833f
C218 VTAIL.n139 B 0.01012f
C219 VTAIL.n140 B 0.010715f
C220 VTAIL.n141 B 0.02392f
C221 VTAIL.n142 B 0.02392f
C222 VTAIL.n143 B 0.010715f
C223 VTAIL.n144 B 0.01012f
C224 VTAIL.n145 B 0.018833f
C225 VTAIL.n146 B 0.018833f
C226 VTAIL.n147 B 0.01012f
C227 VTAIL.n148 B 0.01012f
C228 VTAIL.n149 B 0.010715f
C229 VTAIL.n150 B 0.02392f
C230 VTAIL.n151 B 0.02392f
C231 VTAIL.n152 B 0.048638f
C232 VTAIL.n153 B 0.010418f
C233 VTAIL.n154 B 0.01012f
C234 VTAIL.n155 B 0.046105f
C235 VTAIL.n156 B 0.026968f
C236 VTAIL.n157 B 0.141786f
C237 VTAIL.t13 B 0.208654f
C238 VTAIL.t9 B 0.208654f
C239 VTAIL.n158 B 1.82811f
C240 VTAIL.n159 B 0.371068f
C241 VTAIL.n160 B 0.024693f
C242 VTAIL.n161 B 0.018833f
C243 VTAIL.n162 B 0.010418f
C244 VTAIL.n163 B 0.02392f
C245 VTAIL.n164 B 0.010715f
C246 VTAIL.n165 B 0.018833f
C247 VTAIL.n166 B 0.01012f
C248 VTAIL.n167 B 0.02392f
C249 VTAIL.n168 B 0.010715f
C250 VTAIL.n169 B 0.018833f
C251 VTAIL.n170 B 0.01012f
C252 VTAIL.n171 B 0.02392f
C253 VTAIL.n172 B 0.010715f
C254 VTAIL.n173 B 0.018833f
C255 VTAIL.n174 B 0.01012f
C256 VTAIL.n175 B 0.02392f
C257 VTAIL.n176 B 0.010715f
C258 VTAIL.n177 B 0.018833f
C259 VTAIL.n178 B 0.01012f
C260 VTAIL.n179 B 0.02392f
C261 VTAIL.n180 B 0.010715f
C262 VTAIL.n181 B 0.018833f
C263 VTAIL.n182 B 0.01012f
C264 VTAIL.n183 B 0.01794f
C265 VTAIL.n184 B 0.014131f
C266 VTAIL.t11 B 0.039379f
C267 VTAIL.n185 B 0.118207f
C268 VTAIL.n186 B 1.14073f
C269 VTAIL.n187 B 0.01012f
C270 VTAIL.n188 B 0.010715f
C271 VTAIL.n189 B 0.02392f
C272 VTAIL.n190 B 0.02392f
C273 VTAIL.n191 B 0.010715f
C274 VTAIL.n192 B 0.01012f
C275 VTAIL.n193 B 0.018833f
C276 VTAIL.n194 B 0.018833f
C277 VTAIL.n195 B 0.01012f
C278 VTAIL.n196 B 0.010715f
C279 VTAIL.n197 B 0.02392f
C280 VTAIL.n198 B 0.02392f
C281 VTAIL.n199 B 0.010715f
C282 VTAIL.n200 B 0.01012f
C283 VTAIL.n201 B 0.018833f
C284 VTAIL.n202 B 0.018833f
C285 VTAIL.n203 B 0.01012f
C286 VTAIL.n204 B 0.010715f
C287 VTAIL.n205 B 0.02392f
C288 VTAIL.n206 B 0.02392f
C289 VTAIL.n207 B 0.010715f
C290 VTAIL.n208 B 0.01012f
C291 VTAIL.n209 B 0.018833f
C292 VTAIL.n210 B 0.018833f
C293 VTAIL.n211 B 0.01012f
C294 VTAIL.n212 B 0.010715f
C295 VTAIL.n213 B 0.02392f
C296 VTAIL.n214 B 0.02392f
C297 VTAIL.n215 B 0.010715f
C298 VTAIL.n216 B 0.01012f
C299 VTAIL.n217 B 0.018833f
C300 VTAIL.n218 B 0.018833f
C301 VTAIL.n219 B 0.01012f
C302 VTAIL.n220 B 0.010715f
C303 VTAIL.n221 B 0.02392f
C304 VTAIL.n222 B 0.02392f
C305 VTAIL.n223 B 0.010715f
C306 VTAIL.n224 B 0.01012f
C307 VTAIL.n225 B 0.018833f
C308 VTAIL.n226 B 0.018833f
C309 VTAIL.n227 B 0.01012f
C310 VTAIL.n228 B 0.01012f
C311 VTAIL.n229 B 0.010715f
C312 VTAIL.n230 B 0.02392f
C313 VTAIL.n231 B 0.02392f
C314 VTAIL.n232 B 0.048638f
C315 VTAIL.n233 B 0.010418f
C316 VTAIL.n234 B 0.01012f
C317 VTAIL.n235 B 0.046105f
C318 VTAIL.n236 B 0.026968f
C319 VTAIL.n237 B 1.19829f
C320 VTAIL.n238 B 0.024693f
C321 VTAIL.n239 B 0.018833f
C322 VTAIL.n240 B 0.010418f
C323 VTAIL.n241 B 0.02392f
C324 VTAIL.n242 B 0.01012f
C325 VTAIL.n243 B 0.010715f
C326 VTAIL.n244 B 0.018833f
C327 VTAIL.n245 B 0.01012f
C328 VTAIL.n246 B 0.02392f
C329 VTAIL.n247 B 0.010715f
C330 VTAIL.n248 B 0.018833f
C331 VTAIL.n249 B 0.01012f
C332 VTAIL.n250 B 0.02392f
C333 VTAIL.n251 B 0.010715f
C334 VTAIL.n252 B 0.018833f
C335 VTAIL.n253 B 0.01012f
C336 VTAIL.n254 B 0.02392f
C337 VTAIL.n255 B 0.010715f
C338 VTAIL.n256 B 0.018833f
C339 VTAIL.n257 B 0.01012f
C340 VTAIL.n258 B 0.02392f
C341 VTAIL.n259 B 0.010715f
C342 VTAIL.n260 B 0.018833f
C343 VTAIL.n261 B 0.01012f
C344 VTAIL.n262 B 0.01794f
C345 VTAIL.n263 B 0.014131f
C346 VTAIL.t3 B 0.039379f
C347 VTAIL.n264 B 0.118207f
C348 VTAIL.n265 B 1.14073f
C349 VTAIL.n266 B 0.01012f
C350 VTAIL.n267 B 0.010715f
C351 VTAIL.n268 B 0.02392f
C352 VTAIL.n269 B 0.02392f
C353 VTAIL.n270 B 0.010715f
C354 VTAIL.n271 B 0.01012f
C355 VTAIL.n272 B 0.018833f
C356 VTAIL.n273 B 0.018833f
C357 VTAIL.n274 B 0.01012f
C358 VTAIL.n275 B 0.010715f
C359 VTAIL.n276 B 0.02392f
C360 VTAIL.n277 B 0.02392f
C361 VTAIL.n278 B 0.010715f
C362 VTAIL.n279 B 0.01012f
C363 VTAIL.n280 B 0.018833f
C364 VTAIL.n281 B 0.018833f
C365 VTAIL.n282 B 0.01012f
C366 VTAIL.n283 B 0.010715f
C367 VTAIL.n284 B 0.02392f
C368 VTAIL.n285 B 0.02392f
C369 VTAIL.n286 B 0.010715f
C370 VTAIL.n287 B 0.01012f
C371 VTAIL.n288 B 0.018833f
C372 VTAIL.n289 B 0.018833f
C373 VTAIL.n290 B 0.01012f
C374 VTAIL.n291 B 0.010715f
C375 VTAIL.n292 B 0.02392f
C376 VTAIL.n293 B 0.02392f
C377 VTAIL.n294 B 0.010715f
C378 VTAIL.n295 B 0.01012f
C379 VTAIL.n296 B 0.018833f
C380 VTAIL.n297 B 0.018833f
C381 VTAIL.n298 B 0.01012f
C382 VTAIL.n299 B 0.010715f
C383 VTAIL.n300 B 0.02392f
C384 VTAIL.n301 B 0.02392f
C385 VTAIL.n302 B 0.010715f
C386 VTAIL.n303 B 0.01012f
C387 VTAIL.n304 B 0.018833f
C388 VTAIL.n305 B 0.018833f
C389 VTAIL.n306 B 0.01012f
C390 VTAIL.n307 B 0.010715f
C391 VTAIL.n308 B 0.02392f
C392 VTAIL.n309 B 0.02392f
C393 VTAIL.n310 B 0.048638f
C394 VTAIL.n311 B 0.010418f
C395 VTAIL.n312 B 0.01012f
C396 VTAIL.n313 B 0.046105f
C397 VTAIL.n314 B 0.026968f
C398 VTAIL.n315 B 1.19829f
C399 VTAIL.t5 B 0.208654f
C400 VTAIL.t2 B 0.208654f
C401 VTAIL.n316 B 1.82812f
C402 VTAIL.n317 B 0.371058f
C403 VTAIL.n318 B 0.024693f
C404 VTAIL.n319 B 0.018833f
C405 VTAIL.n320 B 0.010418f
C406 VTAIL.n321 B 0.02392f
C407 VTAIL.n322 B 0.01012f
C408 VTAIL.n323 B 0.010715f
C409 VTAIL.n324 B 0.018833f
C410 VTAIL.n325 B 0.01012f
C411 VTAIL.n326 B 0.02392f
C412 VTAIL.n327 B 0.010715f
C413 VTAIL.n328 B 0.018833f
C414 VTAIL.n329 B 0.01012f
C415 VTAIL.n330 B 0.02392f
C416 VTAIL.n331 B 0.010715f
C417 VTAIL.n332 B 0.018833f
C418 VTAIL.n333 B 0.01012f
C419 VTAIL.n334 B 0.02392f
C420 VTAIL.n335 B 0.010715f
C421 VTAIL.n336 B 0.018833f
C422 VTAIL.n337 B 0.01012f
C423 VTAIL.n338 B 0.02392f
C424 VTAIL.n339 B 0.010715f
C425 VTAIL.n340 B 0.018833f
C426 VTAIL.n341 B 0.01012f
C427 VTAIL.n342 B 0.01794f
C428 VTAIL.n343 B 0.014131f
C429 VTAIL.t0 B 0.039379f
C430 VTAIL.n344 B 0.118207f
C431 VTAIL.n345 B 1.14073f
C432 VTAIL.n346 B 0.01012f
C433 VTAIL.n347 B 0.010715f
C434 VTAIL.n348 B 0.02392f
C435 VTAIL.n349 B 0.02392f
C436 VTAIL.n350 B 0.010715f
C437 VTAIL.n351 B 0.01012f
C438 VTAIL.n352 B 0.018833f
C439 VTAIL.n353 B 0.018833f
C440 VTAIL.n354 B 0.01012f
C441 VTAIL.n355 B 0.010715f
C442 VTAIL.n356 B 0.02392f
C443 VTAIL.n357 B 0.02392f
C444 VTAIL.n358 B 0.010715f
C445 VTAIL.n359 B 0.01012f
C446 VTAIL.n360 B 0.018833f
C447 VTAIL.n361 B 0.018833f
C448 VTAIL.n362 B 0.01012f
C449 VTAIL.n363 B 0.010715f
C450 VTAIL.n364 B 0.02392f
C451 VTAIL.n365 B 0.02392f
C452 VTAIL.n366 B 0.010715f
C453 VTAIL.n367 B 0.01012f
C454 VTAIL.n368 B 0.018833f
C455 VTAIL.n369 B 0.018833f
C456 VTAIL.n370 B 0.01012f
C457 VTAIL.n371 B 0.010715f
C458 VTAIL.n372 B 0.02392f
C459 VTAIL.n373 B 0.02392f
C460 VTAIL.n374 B 0.010715f
C461 VTAIL.n375 B 0.01012f
C462 VTAIL.n376 B 0.018833f
C463 VTAIL.n377 B 0.018833f
C464 VTAIL.n378 B 0.01012f
C465 VTAIL.n379 B 0.010715f
C466 VTAIL.n380 B 0.02392f
C467 VTAIL.n381 B 0.02392f
C468 VTAIL.n382 B 0.010715f
C469 VTAIL.n383 B 0.01012f
C470 VTAIL.n384 B 0.018833f
C471 VTAIL.n385 B 0.018833f
C472 VTAIL.n386 B 0.01012f
C473 VTAIL.n387 B 0.010715f
C474 VTAIL.n388 B 0.02392f
C475 VTAIL.n389 B 0.02392f
C476 VTAIL.n390 B 0.048638f
C477 VTAIL.n391 B 0.010418f
C478 VTAIL.n392 B 0.01012f
C479 VTAIL.n393 B 0.046105f
C480 VTAIL.n394 B 0.026968f
C481 VTAIL.n395 B 0.141786f
C482 VTAIL.n396 B 0.024693f
C483 VTAIL.n397 B 0.018833f
C484 VTAIL.n398 B 0.010418f
C485 VTAIL.n399 B 0.02392f
C486 VTAIL.n400 B 0.01012f
C487 VTAIL.n401 B 0.010715f
C488 VTAIL.n402 B 0.018833f
C489 VTAIL.n403 B 0.01012f
C490 VTAIL.n404 B 0.02392f
C491 VTAIL.n405 B 0.010715f
C492 VTAIL.n406 B 0.018833f
C493 VTAIL.n407 B 0.01012f
C494 VTAIL.n408 B 0.02392f
C495 VTAIL.n409 B 0.010715f
C496 VTAIL.n410 B 0.018833f
C497 VTAIL.n411 B 0.01012f
C498 VTAIL.n412 B 0.02392f
C499 VTAIL.n413 B 0.010715f
C500 VTAIL.n414 B 0.018833f
C501 VTAIL.n415 B 0.01012f
C502 VTAIL.n416 B 0.02392f
C503 VTAIL.n417 B 0.010715f
C504 VTAIL.n418 B 0.018833f
C505 VTAIL.n419 B 0.01012f
C506 VTAIL.n420 B 0.01794f
C507 VTAIL.n421 B 0.014131f
C508 VTAIL.t10 B 0.039379f
C509 VTAIL.n422 B 0.118207f
C510 VTAIL.n423 B 1.14073f
C511 VTAIL.n424 B 0.01012f
C512 VTAIL.n425 B 0.010715f
C513 VTAIL.n426 B 0.02392f
C514 VTAIL.n427 B 0.02392f
C515 VTAIL.n428 B 0.010715f
C516 VTAIL.n429 B 0.01012f
C517 VTAIL.n430 B 0.018833f
C518 VTAIL.n431 B 0.018833f
C519 VTAIL.n432 B 0.01012f
C520 VTAIL.n433 B 0.010715f
C521 VTAIL.n434 B 0.02392f
C522 VTAIL.n435 B 0.02392f
C523 VTAIL.n436 B 0.010715f
C524 VTAIL.n437 B 0.01012f
C525 VTAIL.n438 B 0.018833f
C526 VTAIL.n439 B 0.018833f
C527 VTAIL.n440 B 0.01012f
C528 VTAIL.n441 B 0.010715f
C529 VTAIL.n442 B 0.02392f
C530 VTAIL.n443 B 0.02392f
C531 VTAIL.n444 B 0.010715f
C532 VTAIL.n445 B 0.01012f
C533 VTAIL.n446 B 0.018833f
C534 VTAIL.n447 B 0.018833f
C535 VTAIL.n448 B 0.01012f
C536 VTAIL.n449 B 0.010715f
C537 VTAIL.n450 B 0.02392f
C538 VTAIL.n451 B 0.02392f
C539 VTAIL.n452 B 0.010715f
C540 VTAIL.n453 B 0.01012f
C541 VTAIL.n454 B 0.018833f
C542 VTAIL.n455 B 0.018833f
C543 VTAIL.n456 B 0.01012f
C544 VTAIL.n457 B 0.010715f
C545 VTAIL.n458 B 0.02392f
C546 VTAIL.n459 B 0.02392f
C547 VTAIL.n460 B 0.010715f
C548 VTAIL.n461 B 0.01012f
C549 VTAIL.n462 B 0.018833f
C550 VTAIL.n463 B 0.018833f
C551 VTAIL.n464 B 0.01012f
C552 VTAIL.n465 B 0.010715f
C553 VTAIL.n466 B 0.02392f
C554 VTAIL.n467 B 0.02392f
C555 VTAIL.n468 B 0.048638f
C556 VTAIL.n469 B 0.010418f
C557 VTAIL.n470 B 0.01012f
C558 VTAIL.n471 B 0.046105f
C559 VTAIL.n472 B 0.026968f
C560 VTAIL.n473 B 0.141786f
C561 VTAIL.t12 B 0.208654f
C562 VTAIL.t15 B 0.208654f
C563 VTAIL.n474 B 1.82812f
C564 VTAIL.n475 B 0.371058f
C565 VTAIL.n476 B 0.024693f
C566 VTAIL.n477 B 0.018833f
C567 VTAIL.n478 B 0.010418f
C568 VTAIL.n479 B 0.02392f
C569 VTAIL.n480 B 0.01012f
C570 VTAIL.n481 B 0.010715f
C571 VTAIL.n482 B 0.018833f
C572 VTAIL.n483 B 0.01012f
C573 VTAIL.n484 B 0.02392f
C574 VTAIL.n485 B 0.010715f
C575 VTAIL.n486 B 0.018833f
C576 VTAIL.n487 B 0.01012f
C577 VTAIL.n488 B 0.02392f
C578 VTAIL.n489 B 0.010715f
C579 VTAIL.n490 B 0.018833f
C580 VTAIL.n491 B 0.01012f
C581 VTAIL.n492 B 0.02392f
C582 VTAIL.n493 B 0.010715f
C583 VTAIL.n494 B 0.018833f
C584 VTAIL.n495 B 0.01012f
C585 VTAIL.n496 B 0.02392f
C586 VTAIL.n497 B 0.010715f
C587 VTAIL.n498 B 0.018833f
C588 VTAIL.n499 B 0.01012f
C589 VTAIL.n500 B 0.01794f
C590 VTAIL.n501 B 0.014131f
C591 VTAIL.t8 B 0.039379f
C592 VTAIL.n502 B 0.118207f
C593 VTAIL.n503 B 1.14073f
C594 VTAIL.n504 B 0.01012f
C595 VTAIL.n505 B 0.010715f
C596 VTAIL.n506 B 0.02392f
C597 VTAIL.n507 B 0.02392f
C598 VTAIL.n508 B 0.010715f
C599 VTAIL.n509 B 0.01012f
C600 VTAIL.n510 B 0.018833f
C601 VTAIL.n511 B 0.018833f
C602 VTAIL.n512 B 0.01012f
C603 VTAIL.n513 B 0.010715f
C604 VTAIL.n514 B 0.02392f
C605 VTAIL.n515 B 0.02392f
C606 VTAIL.n516 B 0.010715f
C607 VTAIL.n517 B 0.01012f
C608 VTAIL.n518 B 0.018833f
C609 VTAIL.n519 B 0.018833f
C610 VTAIL.n520 B 0.01012f
C611 VTAIL.n521 B 0.010715f
C612 VTAIL.n522 B 0.02392f
C613 VTAIL.n523 B 0.02392f
C614 VTAIL.n524 B 0.010715f
C615 VTAIL.n525 B 0.01012f
C616 VTAIL.n526 B 0.018833f
C617 VTAIL.n527 B 0.018833f
C618 VTAIL.n528 B 0.01012f
C619 VTAIL.n529 B 0.010715f
C620 VTAIL.n530 B 0.02392f
C621 VTAIL.n531 B 0.02392f
C622 VTAIL.n532 B 0.010715f
C623 VTAIL.n533 B 0.01012f
C624 VTAIL.n534 B 0.018833f
C625 VTAIL.n535 B 0.018833f
C626 VTAIL.n536 B 0.01012f
C627 VTAIL.n537 B 0.010715f
C628 VTAIL.n538 B 0.02392f
C629 VTAIL.n539 B 0.02392f
C630 VTAIL.n540 B 0.010715f
C631 VTAIL.n541 B 0.01012f
C632 VTAIL.n542 B 0.018833f
C633 VTAIL.n543 B 0.018833f
C634 VTAIL.n544 B 0.01012f
C635 VTAIL.n545 B 0.010715f
C636 VTAIL.n546 B 0.02392f
C637 VTAIL.n547 B 0.02392f
C638 VTAIL.n548 B 0.048638f
C639 VTAIL.n549 B 0.010418f
C640 VTAIL.n550 B 0.01012f
C641 VTAIL.n551 B 0.046105f
C642 VTAIL.n552 B 0.026968f
C643 VTAIL.n553 B 1.19829f
C644 VTAIL.n554 B 0.024693f
C645 VTAIL.n555 B 0.018833f
C646 VTAIL.n556 B 0.010418f
C647 VTAIL.n557 B 0.02392f
C648 VTAIL.n558 B 0.010715f
C649 VTAIL.n559 B 0.018833f
C650 VTAIL.n560 B 0.01012f
C651 VTAIL.n561 B 0.02392f
C652 VTAIL.n562 B 0.010715f
C653 VTAIL.n563 B 0.018833f
C654 VTAIL.n564 B 0.01012f
C655 VTAIL.n565 B 0.02392f
C656 VTAIL.n566 B 0.010715f
C657 VTAIL.n567 B 0.018833f
C658 VTAIL.n568 B 0.01012f
C659 VTAIL.n569 B 0.02392f
C660 VTAIL.n570 B 0.010715f
C661 VTAIL.n571 B 0.018833f
C662 VTAIL.n572 B 0.01012f
C663 VTAIL.n573 B 0.02392f
C664 VTAIL.n574 B 0.010715f
C665 VTAIL.n575 B 0.018833f
C666 VTAIL.n576 B 0.01012f
C667 VTAIL.n577 B 0.01794f
C668 VTAIL.n578 B 0.014131f
C669 VTAIL.t6 B 0.039379f
C670 VTAIL.n579 B 0.118207f
C671 VTAIL.n580 B 1.14073f
C672 VTAIL.n581 B 0.01012f
C673 VTAIL.n582 B 0.010715f
C674 VTAIL.n583 B 0.02392f
C675 VTAIL.n584 B 0.02392f
C676 VTAIL.n585 B 0.010715f
C677 VTAIL.n586 B 0.01012f
C678 VTAIL.n587 B 0.018833f
C679 VTAIL.n588 B 0.018833f
C680 VTAIL.n589 B 0.01012f
C681 VTAIL.n590 B 0.010715f
C682 VTAIL.n591 B 0.02392f
C683 VTAIL.n592 B 0.02392f
C684 VTAIL.n593 B 0.010715f
C685 VTAIL.n594 B 0.01012f
C686 VTAIL.n595 B 0.018833f
C687 VTAIL.n596 B 0.018833f
C688 VTAIL.n597 B 0.01012f
C689 VTAIL.n598 B 0.010715f
C690 VTAIL.n599 B 0.02392f
C691 VTAIL.n600 B 0.02392f
C692 VTAIL.n601 B 0.010715f
C693 VTAIL.n602 B 0.01012f
C694 VTAIL.n603 B 0.018833f
C695 VTAIL.n604 B 0.018833f
C696 VTAIL.n605 B 0.01012f
C697 VTAIL.n606 B 0.010715f
C698 VTAIL.n607 B 0.02392f
C699 VTAIL.n608 B 0.02392f
C700 VTAIL.n609 B 0.010715f
C701 VTAIL.n610 B 0.01012f
C702 VTAIL.n611 B 0.018833f
C703 VTAIL.n612 B 0.018833f
C704 VTAIL.n613 B 0.01012f
C705 VTAIL.n614 B 0.010715f
C706 VTAIL.n615 B 0.02392f
C707 VTAIL.n616 B 0.02392f
C708 VTAIL.n617 B 0.010715f
C709 VTAIL.n618 B 0.01012f
C710 VTAIL.n619 B 0.018833f
C711 VTAIL.n620 B 0.018833f
C712 VTAIL.n621 B 0.01012f
C713 VTAIL.n622 B 0.01012f
C714 VTAIL.n623 B 0.010715f
C715 VTAIL.n624 B 0.02392f
C716 VTAIL.n625 B 0.02392f
C717 VTAIL.n626 B 0.048638f
C718 VTAIL.n627 B 0.010418f
C719 VTAIL.n628 B 0.01012f
C720 VTAIL.n629 B 0.046105f
C721 VTAIL.n630 B 0.026968f
C722 VTAIL.n631 B 1.19476f
C723 VDD1.t1 B 0.278383f
C724 VDD1.t6 B 0.278383f
C725 VDD1.n0 B 2.51573f
C726 VDD1.t7 B 0.278383f
C727 VDD1.t2 B 0.278383f
C728 VDD1.n1 B 2.5149f
C729 VDD1.t5 B 0.278383f
C730 VDD1.t4 B 0.278383f
C731 VDD1.n2 B 2.5149f
C732 VDD1.n3 B 2.82277f
C733 VDD1.t3 B 0.278383f
C734 VDD1.t0 B 0.278383f
C735 VDD1.n4 B 2.51029f
C736 VDD1.n5 B 2.76313f
C737 VP.n0 B 0.030906f
C738 VP.t1 B 1.77817f
C739 VP.n1 B 0.051767f
C740 VP.n2 B 0.030906f
C741 VP.t6 B 1.77817f
C742 VP.n3 B 0.056292f
C743 VP.n4 B 0.030906f
C744 VP.n5 B 0.042883f
C745 VP.n6 B 0.030906f
C746 VP.t7 B 1.77817f
C747 VP.n7 B 0.051767f
C748 VP.n8 B 0.030906f
C749 VP.t0 B 1.77817f
C750 VP.n9 B 0.056292f
C751 VP.t5 B 1.87939f
C752 VP.t3 B 1.77817f
C753 VP.n10 B 0.702371f
C754 VP.n11 B 0.703316f
C755 VP.n12 B 0.196509f
C756 VP.n13 B 0.030906f
C757 VP.n14 B 0.024962f
C758 VP.n15 B 0.056292f
C759 VP.n16 B 0.635451f
C760 VP.n17 B 0.033829f
C761 VP.n18 B 0.030906f
C762 VP.n19 B 0.030906f
C763 VP.n20 B 0.030906f
C764 VP.n21 B 0.038086f
C765 VP.n22 B 0.042883f
C766 VP.n23 B 0.701492f
C767 VP.n24 B 1.54563f
C768 VP.t4 B 1.77817f
C769 VP.n25 B 0.701492f
C770 VP.n26 B 1.56922f
C771 VP.n27 B 0.030906f
C772 VP.n28 B 0.030906f
C773 VP.n29 B 0.038086f
C774 VP.n30 B 0.051767f
C775 VP.t2 B 1.77817f
C776 VP.n31 B 0.635451f
C777 VP.n32 B 0.033829f
C778 VP.n33 B 0.030906f
C779 VP.n34 B 0.030906f
C780 VP.n35 B 0.030906f
C781 VP.n36 B 0.024962f
C782 VP.n37 B 0.056292f
C783 VP.n38 B 0.635451f
C784 VP.n39 B 0.033829f
C785 VP.n40 B 0.030906f
C786 VP.n41 B 0.030906f
C787 VP.n42 B 0.030906f
C788 VP.n43 B 0.038086f
C789 VP.n44 B 0.042883f
C790 VP.n45 B 0.701492f
C791 VP.n46 B 0.029086f
.ends

