* NGSPICE file created from diff_pair_sample_1620.ext - technology: sky130A

.subckt diff_pair_sample_1620 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n3010_n2136# sky130_fd_pr__pfet_01v8 ad=2.2776 pd=12.46 as=0 ps=0 w=5.84 l=2.22
X1 VDD2.t5 VN.t0 VTAIL.t4 w_n3010_n2136# sky130_fd_pr__pfet_01v8 ad=2.2776 pd=12.46 as=0.9636 ps=6.17 w=5.84 l=2.22
X2 B.t8 B.t6 B.t7 w_n3010_n2136# sky130_fd_pr__pfet_01v8 ad=2.2776 pd=12.46 as=0 ps=0 w=5.84 l=2.22
X3 VDD2.t4 VN.t1 VTAIL.t5 w_n3010_n2136# sky130_fd_pr__pfet_01v8 ad=0.9636 pd=6.17 as=2.2776 ps=12.46 w=5.84 l=2.22
X4 VDD2.t3 VN.t2 VTAIL.t7 w_n3010_n2136# sky130_fd_pr__pfet_01v8 ad=2.2776 pd=12.46 as=0.9636 ps=6.17 w=5.84 l=2.22
X5 B.t5 B.t3 B.t4 w_n3010_n2136# sky130_fd_pr__pfet_01v8 ad=2.2776 pd=12.46 as=0 ps=0 w=5.84 l=2.22
X6 VDD2.t2 VN.t3 VTAIL.t9 w_n3010_n2136# sky130_fd_pr__pfet_01v8 ad=0.9636 pd=6.17 as=2.2776 ps=12.46 w=5.84 l=2.22
X7 VDD1.t5 VP.t0 VTAIL.t2 w_n3010_n2136# sky130_fd_pr__pfet_01v8 ad=0.9636 pd=6.17 as=2.2776 ps=12.46 w=5.84 l=2.22
X8 VDD1.t4 VP.t1 VTAIL.t3 w_n3010_n2136# sky130_fd_pr__pfet_01v8 ad=0.9636 pd=6.17 as=2.2776 ps=12.46 w=5.84 l=2.22
X9 VTAIL.t6 VN.t4 VDD2.t1 w_n3010_n2136# sky130_fd_pr__pfet_01v8 ad=0.9636 pd=6.17 as=0.9636 ps=6.17 w=5.84 l=2.22
X10 VTAIL.t8 VN.t5 VDD2.t0 w_n3010_n2136# sky130_fd_pr__pfet_01v8 ad=0.9636 pd=6.17 as=0.9636 ps=6.17 w=5.84 l=2.22
X11 B.t2 B.t0 B.t1 w_n3010_n2136# sky130_fd_pr__pfet_01v8 ad=2.2776 pd=12.46 as=0 ps=0 w=5.84 l=2.22
X12 VDD1.t3 VP.t2 VTAIL.t1 w_n3010_n2136# sky130_fd_pr__pfet_01v8 ad=2.2776 pd=12.46 as=0.9636 ps=6.17 w=5.84 l=2.22
X13 VTAIL.t10 VP.t3 VDD1.t2 w_n3010_n2136# sky130_fd_pr__pfet_01v8 ad=0.9636 pd=6.17 as=0.9636 ps=6.17 w=5.84 l=2.22
X14 VTAIL.t0 VP.t4 VDD1.t1 w_n3010_n2136# sky130_fd_pr__pfet_01v8 ad=0.9636 pd=6.17 as=0.9636 ps=6.17 w=5.84 l=2.22
X15 VDD1.t0 VP.t5 VTAIL.t11 w_n3010_n2136# sky130_fd_pr__pfet_01v8 ad=2.2776 pd=12.46 as=0.9636 ps=6.17 w=5.84 l=2.22
R0 B.n402 B.n53 585
R1 B.n404 B.n403 585
R2 B.n405 B.n52 585
R3 B.n407 B.n406 585
R4 B.n408 B.n51 585
R5 B.n410 B.n409 585
R6 B.n411 B.n50 585
R7 B.n413 B.n412 585
R8 B.n414 B.n49 585
R9 B.n416 B.n415 585
R10 B.n417 B.n48 585
R11 B.n419 B.n418 585
R12 B.n420 B.n47 585
R13 B.n422 B.n421 585
R14 B.n423 B.n46 585
R15 B.n425 B.n424 585
R16 B.n426 B.n45 585
R17 B.n428 B.n427 585
R18 B.n429 B.n44 585
R19 B.n431 B.n430 585
R20 B.n432 B.n43 585
R21 B.n434 B.n433 585
R22 B.n435 B.n42 585
R23 B.n437 B.n436 585
R24 B.n439 B.n39 585
R25 B.n441 B.n440 585
R26 B.n442 B.n38 585
R27 B.n444 B.n443 585
R28 B.n445 B.n37 585
R29 B.n447 B.n446 585
R30 B.n448 B.n36 585
R31 B.n450 B.n449 585
R32 B.n451 B.n33 585
R33 B.n454 B.n453 585
R34 B.n455 B.n32 585
R35 B.n457 B.n456 585
R36 B.n458 B.n31 585
R37 B.n460 B.n459 585
R38 B.n461 B.n30 585
R39 B.n463 B.n462 585
R40 B.n464 B.n29 585
R41 B.n466 B.n465 585
R42 B.n467 B.n28 585
R43 B.n469 B.n468 585
R44 B.n470 B.n27 585
R45 B.n472 B.n471 585
R46 B.n473 B.n26 585
R47 B.n475 B.n474 585
R48 B.n476 B.n25 585
R49 B.n478 B.n477 585
R50 B.n479 B.n24 585
R51 B.n481 B.n480 585
R52 B.n482 B.n23 585
R53 B.n484 B.n483 585
R54 B.n485 B.n22 585
R55 B.n487 B.n486 585
R56 B.n488 B.n21 585
R57 B.n401 B.n400 585
R58 B.n399 B.n54 585
R59 B.n398 B.n397 585
R60 B.n396 B.n55 585
R61 B.n395 B.n394 585
R62 B.n393 B.n56 585
R63 B.n392 B.n391 585
R64 B.n390 B.n57 585
R65 B.n389 B.n388 585
R66 B.n387 B.n58 585
R67 B.n386 B.n385 585
R68 B.n384 B.n59 585
R69 B.n383 B.n382 585
R70 B.n381 B.n60 585
R71 B.n380 B.n379 585
R72 B.n378 B.n61 585
R73 B.n377 B.n376 585
R74 B.n375 B.n62 585
R75 B.n374 B.n373 585
R76 B.n372 B.n63 585
R77 B.n371 B.n370 585
R78 B.n369 B.n64 585
R79 B.n368 B.n367 585
R80 B.n366 B.n65 585
R81 B.n365 B.n364 585
R82 B.n363 B.n66 585
R83 B.n362 B.n361 585
R84 B.n360 B.n67 585
R85 B.n359 B.n358 585
R86 B.n357 B.n68 585
R87 B.n356 B.n355 585
R88 B.n354 B.n69 585
R89 B.n353 B.n352 585
R90 B.n351 B.n70 585
R91 B.n350 B.n349 585
R92 B.n348 B.n71 585
R93 B.n347 B.n346 585
R94 B.n345 B.n72 585
R95 B.n344 B.n343 585
R96 B.n342 B.n73 585
R97 B.n341 B.n340 585
R98 B.n339 B.n74 585
R99 B.n338 B.n337 585
R100 B.n336 B.n75 585
R101 B.n335 B.n334 585
R102 B.n333 B.n76 585
R103 B.n332 B.n331 585
R104 B.n330 B.n77 585
R105 B.n329 B.n328 585
R106 B.n327 B.n78 585
R107 B.n326 B.n325 585
R108 B.n324 B.n79 585
R109 B.n323 B.n322 585
R110 B.n321 B.n80 585
R111 B.n320 B.n319 585
R112 B.n318 B.n81 585
R113 B.n317 B.n316 585
R114 B.n315 B.n82 585
R115 B.n314 B.n313 585
R116 B.n312 B.n83 585
R117 B.n311 B.n310 585
R118 B.n309 B.n84 585
R119 B.n308 B.n307 585
R120 B.n306 B.n85 585
R121 B.n305 B.n304 585
R122 B.n303 B.n86 585
R123 B.n302 B.n301 585
R124 B.n300 B.n87 585
R125 B.n299 B.n298 585
R126 B.n297 B.n88 585
R127 B.n296 B.n295 585
R128 B.n294 B.n89 585
R129 B.n293 B.n292 585
R130 B.n291 B.n90 585
R131 B.n290 B.n289 585
R132 B.n288 B.n91 585
R133 B.n287 B.n286 585
R134 B.n200 B.n199 585
R135 B.n201 B.n124 585
R136 B.n203 B.n202 585
R137 B.n204 B.n123 585
R138 B.n206 B.n205 585
R139 B.n207 B.n122 585
R140 B.n209 B.n208 585
R141 B.n210 B.n121 585
R142 B.n212 B.n211 585
R143 B.n213 B.n120 585
R144 B.n215 B.n214 585
R145 B.n216 B.n119 585
R146 B.n218 B.n217 585
R147 B.n219 B.n118 585
R148 B.n221 B.n220 585
R149 B.n222 B.n117 585
R150 B.n224 B.n223 585
R151 B.n225 B.n116 585
R152 B.n227 B.n226 585
R153 B.n228 B.n115 585
R154 B.n230 B.n229 585
R155 B.n231 B.n114 585
R156 B.n233 B.n232 585
R157 B.n234 B.n111 585
R158 B.n237 B.n236 585
R159 B.n238 B.n110 585
R160 B.n240 B.n239 585
R161 B.n241 B.n109 585
R162 B.n243 B.n242 585
R163 B.n244 B.n108 585
R164 B.n246 B.n245 585
R165 B.n247 B.n107 585
R166 B.n249 B.n248 585
R167 B.n251 B.n250 585
R168 B.n252 B.n103 585
R169 B.n254 B.n253 585
R170 B.n255 B.n102 585
R171 B.n257 B.n256 585
R172 B.n258 B.n101 585
R173 B.n260 B.n259 585
R174 B.n261 B.n100 585
R175 B.n263 B.n262 585
R176 B.n264 B.n99 585
R177 B.n266 B.n265 585
R178 B.n267 B.n98 585
R179 B.n269 B.n268 585
R180 B.n270 B.n97 585
R181 B.n272 B.n271 585
R182 B.n273 B.n96 585
R183 B.n275 B.n274 585
R184 B.n276 B.n95 585
R185 B.n278 B.n277 585
R186 B.n279 B.n94 585
R187 B.n281 B.n280 585
R188 B.n282 B.n93 585
R189 B.n284 B.n283 585
R190 B.n285 B.n92 585
R191 B.n198 B.n125 585
R192 B.n197 B.n196 585
R193 B.n195 B.n126 585
R194 B.n194 B.n193 585
R195 B.n192 B.n127 585
R196 B.n191 B.n190 585
R197 B.n189 B.n128 585
R198 B.n188 B.n187 585
R199 B.n186 B.n129 585
R200 B.n185 B.n184 585
R201 B.n183 B.n130 585
R202 B.n182 B.n181 585
R203 B.n180 B.n131 585
R204 B.n179 B.n178 585
R205 B.n177 B.n132 585
R206 B.n176 B.n175 585
R207 B.n174 B.n133 585
R208 B.n173 B.n172 585
R209 B.n171 B.n134 585
R210 B.n170 B.n169 585
R211 B.n168 B.n135 585
R212 B.n167 B.n166 585
R213 B.n165 B.n136 585
R214 B.n164 B.n163 585
R215 B.n162 B.n137 585
R216 B.n161 B.n160 585
R217 B.n159 B.n138 585
R218 B.n158 B.n157 585
R219 B.n156 B.n139 585
R220 B.n155 B.n154 585
R221 B.n153 B.n140 585
R222 B.n152 B.n151 585
R223 B.n150 B.n141 585
R224 B.n149 B.n148 585
R225 B.n147 B.n142 585
R226 B.n146 B.n145 585
R227 B.n144 B.n143 585
R228 B.n2 B.n0 585
R229 B.n545 B.n1 585
R230 B.n544 B.n543 585
R231 B.n542 B.n3 585
R232 B.n541 B.n540 585
R233 B.n539 B.n4 585
R234 B.n538 B.n537 585
R235 B.n536 B.n5 585
R236 B.n535 B.n534 585
R237 B.n533 B.n6 585
R238 B.n532 B.n531 585
R239 B.n530 B.n7 585
R240 B.n529 B.n528 585
R241 B.n527 B.n8 585
R242 B.n526 B.n525 585
R243 B.n524 B.n9 585
R244 B.n523 B.n522 585
R245 B.n521 B.n10 585
R246 B.n520 B.n519 585
R247 B.n518 B.n11 585
R248 B.n517 B.n516 585
R249 B.n515 B.n12 585
R250 B.n514 B.n513 585
R251 B.n512 B.n13 585
R252 B.n511 B.n510 585
R253 B.n509 B.n14 585
R254 B.n508 B.n507 585
R255 B.n506 B.n15 585
R256 B.n505 B.n504 585
R257 B.n503 B.n16 585
R258 B.n502 B.n501 585
R259 B.n500 B.n17 585
R260 B.n499 B.n498 585
R261 B.n497 B.n18 585
R262 B.n496 B.n495 585
R263 B.n494 B.n19 585
R264 B.n493 B.n492 585
R265 B.n491 B.n20 585
R266 B.n490 B.n489 585
R267 B.n547 B.n546 585
R268 B.n200 B.n125 482.89
R269 B.n490 B.n21 482.89
R270 B.n286 B.n285 482.89
R271 B.n400 B.n53 482.89
R272 B.n104 B.t8 314.545
R273 B.n40 B.t4 314.545
R274 B.n112 B.t2 314.545
R275 B.n34 B.t10 314.545
R276 B.n104 B.t6 270.789
R277 B.n112 B.t0 270.789
R278 B.n34 B.t9 270.789
R279 B.n40 B.t3 270.789
R280 B.n105 B.t7 265.089
R281 B.n41 B.t5 265.089
R282 B.n113 B.t1 265.089
R283 B.n35 B.t11 265.089
R284 B.n196 B.n125 163.367
R285 B.n196 B.n195 163.367
R286 B.n195 B.n194 163.367
R287 B.n194 B.n127 163.367
R288 B.n190 B.n127 163.367
R289 B.n190 B.n189 163.367
R290 B.n189 B.n188 163.367
R291 B.n188 B.n129 163.367
R292 B.n184 B.n129 163.367
R293 B.n184 B.n183 163.367
R294 B.n183 B.n182 163.367
R295 B.n182 B.n131 163.367
R296 B.n178 B.n131 163.367
R297 B.n178 B.n177 163.367
R298 B.n177 B.n176 163.367
R299 B.n176 B.n133 163.367
R300 B.n172 B.n133 163.367
R301 B.n172 B.n171 163.367
R302 B.n171 B.n170 163.367
R303 B.n170 B.n135 163.367
R304 B.n166 B.n135 163.367
R305 B.n166 B.n165 163.367
R306 B.n165 B.n164 163.367
R307 B.n164 B.n137 163.367
R308 B.n160 B.n137 163.367
R309 B.n160 B.n159 163.367
R310 B.n159 B.n158 163.367
R311 B.n158 B.n139 163.367
R312 B.n154 B.n139 163.367
R313 B.n154 B.n153 163.367
R314 B.n153 B.n152 163.367
R315 B.n152 B.n141 163.367
R316 B.n148 B.n141 163.367
R317 B.n148 B.n147 163.367
R318 B.n147 B.n146 163.367
R319 B.n146 B.n143 163.367
R320 B.n143 B.n2 163.367
R321 B.n546 B.n2 163.367
R322 B.n546 B.n545 163.367
R323 B.n545 B.n544 163.367
R324 B.n544 B.n3 163.367
R325 B.n540 B.n3 163.367
R326 B.n540 B.n539 163.367
R327 B.n539 B.n538 163.367
R328 B.n538 B.n5 163.367
R329 B.n534 B.n5 163.367
R330 B.n534 B.n533 163.367
R331 B.n533 B.n532 163.367
R332 B.n532 B.n7 163.367
R333 B.n528 B.n7 163.367
R334 B.n528 B.n527 163.367
R335 B.n527 B.n526 163.367
R336 B.n526 B.n9 163.367
R337 B.n522 B.n9 163.367
R338 B.n522 B.n521 163.367
R339 B.n521 B.n520 163.367
R340 B.n520 B.n11 163.367
R341 B.n516 B.n11 163.367
R342 B.n516 B.n515 163.367
R343 B.n515 B.n514 163.367
R344 B.n514 B.n13 163.367
R345 B.n510 B.n13 163.367
R346 B.n510 B.n509 163.367
R347 B.n509 B.n508 163.367
R348 B.n508 B.n15 163.367
R349 B.n504 B.n15 163.367
R350 B.n504 B.n503 163.367
R351 B.n503 B.n502 163.367
R352 B.n502 B.n17 163.367
R353 B.n498 B.n17 163.367
R354 B.n498 B.n497 163.367
R355 B.n497 B.n496 163.367
R356 B.n496 B.n19 163.367
R357 B.n492 B.n19 163.367
R358 B.n492 B.n491 163.367
R359 B.n491 B.n490 163.367
R360 B.n201 B.n200 163.367
R361 B.n202 B.n201 163.367
R362 B.n202 B.n123 163.367
R363 B.n206 B.n123 163.367
R364 B.n207 B.n206 163.367
R365 B.n208 B.n207 163.367
R366 B.n208 B.n121 163.367
R367 B.n212 B.n121 163.367
R368 B.n213 B.n212 163.367
R369 B.n214 B.n213 163.367
R370 B.n214 B.n119 163.367
R371 B.n218 B.n119 163.367
R372 B.n219 B.n218 163.367
R373 B.n220 B.n219 163.367
R374 B.n220 B.n117 163.367
R375 B.n224 B.n117 163.367
R376 B.n225 B.n224 163.367
R377 B.n226 B.n225 163.367
R378 B.n226 B.n115 163.367
R379 B.n230 B.n115 163.367
R380 B.n231 B.n230 163.367
R381 B.n232 B.n231 163.367
R382 B.n232 B.n111 163.367
R383 B.n237 B.n111 163.367
R384 B.n238 B.n237 163.367
R385 B.n239 B.n238 163.367
R386 B.n239 B.n109 163.367
R387 B.n243 B.n109 163.367
R388 B.n244 B.n243 163.367
R389 B.n245 B.n244 163.367
R390 B.n245 B.n107 163.367
R391 B.n249 B.n107 163.367
R392 B.n250 B.n249 163.367
R393 B.n250 B.n103 163.367
R394 B.n254 B.n103 163.367
R395 B.n255 B.n254 163.367
R396 B.n256 B.n255 163.367
R397 B.n256 B.n101 163.367
R398 B.n260 B.n101 163.367
R399 B.n261 B.n260 163.367
R400 B.n262 B.n261 163.367
R401 B.n262 B.n99 163.367
R402 B.n266 B.n99 163.367
R403 B.n267 B.n266 163.367
R404 B.n268 B.n267 163.367
R405 B.n268 B.n97 163.367
R406 B.n272 B.n97 163.367
R407 B.n273 B.n272 163.367
R408 B.n274 B.n273 163.367
R409 B.n274 B.n95 163.367
R410 B.n278 B.n95 163.367
R411 B.n279 B.n278 163.367
R412 B.n280 B.n279 163.367
R413 B.n280 B.n93 163.367
R414 B.n284 B.n93 163.367
R415 B.n285 B.n284 163.367
R416 B.n286 B.n91 163.367
R417 B.n290 B.n91 163.367
R418 B.n291 B.n290 163.367
R419 B.n292 B.n291 163.367
R420 B.n292 B.n89 163.367
R421 B.n296 B.n89 163.367
R422 B.n297 B.n296 163.367
R423 B.n298 B.n297 163.367
R424 B.n298 B.n87 163.367
R425 B.n302 B.n87 163.367
R426 B.n303 B.n302 163.367
R427 B.n304 B.n303 163.367
R428 B.n304 B.n85 163.367
R429 B.n308 B.n85 163.367
R430 B.n309 B.n308 163.367
R431 B.n310 B.n309 163.367
R432 B.n310 B.n83 163.367
R433 B.n314 B.n83 163.367
R434 B.n315 B.n314 163.367
R435 B.n316 B.n315 163.367
R436 B.n316 B.n81 163.367
R437 B.n320 B.n81 163.367
R438 B.n321 B.n320 163.367
R439 B.n322 B.n321 163.367
R440 B.n322 B.n79 163.367
R441 B.n326 B.n79 163.367
R442 B.n327 B.n326 163.367
R443 B.n328 B.n327 163.367
R444 B.n328 B.n77 163.367
R445 B.n332 B.n77 163.367
R446 B.n333 B.n332 163.367
R447 B.n334 B.n333 163.367
R448 B.n334 B.n75 163.367
R449 B.n338 B.n75 163.367
R450 B.n339 B.n338 163.367
R451 B.n340 B.n339 163.367
R452 B.n340 B.n73 163.367
R453 B.n344 B.n73 163.367
R454 B.n345 B.n344 163.367
R455 B.n346 B.n345 163.367
R456 B.n346 B.n71 163.367
R457 B.n350 B.n71 163.367
R458 B.n351 B.n350 163.367
R459 B.n352 B.n351 163.367
R460 B.n352 B.n69 163.367
R461 B.n356 B.n69 163.367
R462 B.n357 B.n356 163.367
R463 B.n358 B.n357 163.367
R464 B.n358 B.n67 163.367
R465 B.n362 B.n67 163.367
R466 B.n363 B.n362 163.367
R467 B.n364 B.n363 163.367
R468 B.n364 B.n65 163.367
R469 B.n368 B.n65 163.367
R470 B.n369 B.n368 163.367
R471 B.n370 B.n369 163.367
R472 B.n370 B.n63 163.367
R473 B.n374 B.n63 163.367
R474 B.n375 B.n374 163.367
R475 B.n376 B.n375 163.367
R476 B.n376 B.n61 163.367
R477 B.n380 B.n61 163.367
R478 B.n381 B.n380 163.367
R479 B.n382 B.n381 163.367
R480 B.n382 B.n59 163.367
R481 B.n386 B.n59 163.367
R482 B.n387 B.n386 163.367
R483 B.n388 B.n387 163.367
R484 B.n388 B.n57 163.367
R485 B.n392 B.n57 163.367
R486 B.n393 B.n392 163.367
R487 B.n394 B.n393 163.367
R488 B.n394 B.n55 163.367
R489 B.n398 B.n55 163.367
R490 B.n399 B.n398 163.367
R491 B.n400 B.n399 163.367
R492 B.n486 B.n21 163.367
R493 B.n486 B.n485 163.367
R494 B.n485 B.n484 163.367
R495 B.n484 B.n23 163.367
R496 B.n480 B.n23 163.367
R497 B.n480 B.n479 163.367
R498 B.n479 B.n478 163.367
R499 B.n478 B.n25 163.367
R500 B.n474 B.n25 163.367
R501 B.n474 B.n473 163.367
R502 B.n473 B.n472 163.367
R503 B.n472 B.n27 163.367
R504 B.n468 B.n27 163.367
R505 B.n468 B.n467 163.367
R506 B.n467 B.n466 163.367
R507 B.n466 B.n29 163.367
R508 B.n462 B.n29 163.367
R509 B.n462 B.n461 163.367
R510 B.n461 B.n460 163.367
R511 B.n460 B.n31 163.367
R512 B.n456 B.n31 163.367
R513 B.n456 B.n455 163.367
R514 B.n455 B.n454 163.367
R515 B.n454 B.n33 163.367
R516 B.n449 B.n33 163.367
R517 B.n449 B.n448 163.367
R518 B.n448 B.n447 163.367
R519 B.n447 B.n37 163.367
R520 B.n443 B.n37 163.367
R521 B.n443 B.n442 163.367
R522 B.n442 B.n441 163.367
R523 B.n441 B.n39 163.367
R524 B.n436 B.n39 163.367
R525 B.n436 B.n435 163.367
R526 B.n435 B.n434 163.367
R527 B.n434 B.n43 163.367
R528 B.n430 B.n43 163.367
R529 B.n430 B.n429 163.367
R530 B.n429 B.n428 163.367
R531 B.n428 B.n45 163.367
R532 B.n424 B.n45 163.367
R533 B.n424 B.n423 163.367
R534 B.n423 B.n422 163.367
R535 B.n422 B.n47 163.367
R536 B.n418 B.n47 163.367
R537 B.n418 B.n417 163.367
R538 B.n417 B.n416 163.367
R539 B.n416 B.n49 163.367
R540 B.n412 B.n49 163.367
R541 B.n412 B.n411 163.367
R542 B.n411 B.n410 163.367
R543 B.n410 B.n51 163.367
R544 B.n406 B.n51 163.367
R545 B.n406 B.n405 163.367
R546 B.n405 B.n404 163.367
R547 B.n404 B.n53 163.367
R548 B.n106 B.n105 59.5399
R549 B.n235 B.n113 59.5399
R550 B.n452 B.n35 59.5399
R551 B.n438 B.n41 59.5399
R552 B.n105 B.n104 49.455
R553 B.n113 B.n112 49.455
R554 B.n35 B.n34 49.455
R555 B.n41 B.n40 49.455
R556 B.n489 B.n488 31.3761
R557 B.n402 B.n401 31.3761
R558 B.n287 B.n92 31.3761
R559 B.n199 B.n198 31.3761
R560 B B.n547 18.0485
R561 B.n488 B.n487 10.6151
R562 B.n487 B.n22 10.6151
R563 B.n483 B.n22 10.6151
R564 B.n483 B.n482 10.6151
R565 B.n482 B.n481 10.6151
R566 B.n481 B.n24 10.6151
R567 B.n477 B.n24 10.6151
R568 B.n477 B.n476 10.6151
R569 B.n476 B.n475 10.6151
R570 B.n475 B.n26 10.6151
R571 B.n471 B.n26 10.6151
R572 B.n471 B.n470 10.6151
R573 B.n470 B.n469 10.6151
R574 B.n469 B.n28 10.6151
R575 B.n465 B.n28 10.6151
R576 B.n465 B.n464 10.6151
R577 B.n464 B.n463 10.6151
R578 B.n463 B.n30 10.6151
R579 B.n459 B.n30 10.6151
R580 B.n459 B.n458 10.6151
R581 B.n458 B.n457 10.6151
R582 B.n457 B.n32 10.6151
R583 B.n453 B.n32 10.6151
R584 B.n451 B.n450 10.6151
R585 B.n450 B.n36 10.6151
R586 B.n446 B.n36 10.6151
R587 B.n446 B.n445 10.6151
R588 B.n445 B.n444 10.6151
R589 B.n444 B.n38 10.6151
R590 B.n440 B.n38 10.6151
R591 B.n440 B.n439 10.6151
R592 B.n437 B.n42 10.6151
R593 B.n433 B.n42 10.6151
R594 B.n433 B.n432 10.6151
R595 B.n432 B.n431 10.6151
R596 B.n431 B.n44 10.6151
R597 B.n427 B.n44 10.6151
R598 B.n427 B.n426 10.6151
R599 B.n426 B.n425 10.6151
R600 B.n425 B.n46 10.6151
R601 B.n421 B.n46 10.6151
R602 B.n421 B.n420 10.6151
R603 B.n420 B.n419 10.6151
R604 B.n419 B.n48 10.6151
R605 B.n415 B.n48 10.6151
R606 B.n415 B.n414 10.6151
R607 B.n414 B.n413 10.6151
R608 B.n413 B.n50 10.6151
R609 B.n409 B.n50 10.6151
R610 B.n409 B.n408 10.6151
R611 B.n408 B.n407 10.6151
R612 B.n407 B.n52 10.6151
R613 B.n403 B.n52 10.6151
R614 B.n403 B.n402 10.6151
R615 B.n288 B.n287 10.6151
R616 B.n289 B.n288 10.6151
R617 B.n289 B.n90 10.6151
R618 B.n293 B.n90 10.6151
R619 B.n294 B.n293 10.6151
R620 B.n295 B.n294 10.6151
R621 B.n295 B.n88 10.6151
R622 B.n299 B.n88 10.6151
R623 B.n300 B.n299 10.6151
R624 B.n301 B.n300 10.6151
R625 B.n301 B.n86 10.6151
R626 B.n305 B.n86 10.6151
R627 B.n306 B.n305 10.6151
R628 B.n307 B.n306 10.6151
R629 B.n307 B.n84 10.6151
R630 B.n311 B.n84 10.6151
R631 B.n312 B.n311 10.6151
R632 B.n313 B.n312 10.6151
R633 B.n313 B.n82 10.6151
R634 B.n317 B.n82 10.6151
R635 B.n318 B.n317 10.6151
R636 B.n319 B.n318 10.6151
R637 B.n319 B.n80 10.6151
R638 B.n323 B.n80 10.6151
R639 B.n324 B.n323 10.6151
R640 B.n325 B.n324 10.6151
R641 B.n325 B.n78 10.6151
R642 B.n329 B.n78 10.6151
R643 B.n330 B.n329 10.6151
R644 B.n331 B.n330 10.6151
R645 B.n331 B.n76 10.6151
R646 B.n335 B.n76 10.6151
R647 B.n336 B.n335 10.6151
R648 B.n337 B.n336 10.6151
R649 B.n337 B.n74 10.6151
R650 B.n341 B.n74 10.6151
R651 B.n342 B.n341 10.6151
R652 B.n343 B.n342 10.6151
R653 B.n343 B.n72 10.6151
R654 B.n347 B.n72 10.6151
R655 B.n348 B.n347 10.6151
R656 B.n349 B.n348 10.6151
R657 B.n349 B.n70 10.6151
R658 B.n353 B.n70 10.6151
R659 B.n354 B.n353 10.6151
R660 B.n355 B.n354 10.6151
R661 B.n355 B.n68 10.6151
R662 B.n359 B.n68 10.6151
R663 B.n360 B.n359 10.6151
R664 B.n361 B.n360 10.6151
R665 B.n361 B.n66 10.6151
R666 B.n365 B.n66 10.6151
R667 B.n366 B.n365 10.6151
R668 B.n367 B.n366 10.6151
R669 B.n367 B.n64 10.6151
R670 B.n371 B.n64 10.6151
R671 B.n372 B.n371 10.6151
R672 B.n373 B.n372 10.6151
R673 B.n373 B.n62 10.6151
R674 B.n377 B.n62 10.6151
R675 B.n378 B.n377 10.6151
R676 B.n379 B.n378 10.6151
R677 B.n379 B.n60 10.6151
R678 B.n383 B.n60 10.6151
R679 B.n384 B.n383 10.6151
R680 B.n385 B.n384 10.6151
R681 B.n385 B.n58 10.6151
R682 B.n389 B.n58 10.6151
R683 B.n390 B.n389 10.6151
R684 B.n391 B.n390 10.6151
R685 B.n391 B.n56 10.6151
R686 B.n395 B.n56 10.6151
R687 B.n396 B.n395 10.6151
R688 B.n397 B.n396 10.6151
R689 B.n397 B.n54 10.6151
R690 B.n401 B.n54 10.6151
R691 B.n199 B.n124 10.6151
R692 B.n203 B.n124 10.6151
R693 B.n204 B.n203 10.6151
R694 B.n205 B.n204 10.6151
R695 B.n205 B.n122 10.6151
R696 B.n209 B.n122 10.6151
R697 B.n210 B.n209 10.6151
R698 B.n211 B.n210 10.6151
R699 B.n211 B.n120 10.6151
R700 B.n215 B.n120 10.6151
R701 B.n216 B.n215 10.6151
R702 B.n217 B.n216 10.6151
R703 B.n217 B.n118 10.6151
R704 B.n221 B.n118 10.6151
R705 B.n222 B.n221 10.6151
R706 B.n223 B.n222 10.6151
R707 B.n223 B.n116 10.6151
R708 B.n227 B.n116 10.6151
R709 B.n228 B.n227 10.6151
R710 B.n229 B.n228 10.6151
R711 B.n229 B.n114 10.6151
R712 B.n233 B.n114 10.6151
R713 B.n234 B.n233 10.6151
R714 B.n236 B.n110 10.6151
R715 B.n240 B.n110 10.6151
R716 B.n241 B.n240 10.6151
R717 B.n242 B.n241 10.6151
R718 B.n242 B.n108 10.6151
R719 B.n246 B.n108 10.6151
R720 B.n247 B.n246 10.6151
R721 B.n248 B.n247 10.6151
R722 B.n252 B.n251 10.6151
R723 B.n253 B.n252 10.6151
R724 B.n253 B.n102 10.6151
R725 B.n257 B.n102 10.6151
R726 B.n258 B.n257 10.6151
R727 B.n259 B.n258 10.6151
R728 B.n259 B.n100 10.6151
R729 B.n263 B.n100 10.6151
R730 B.n264 B.n263 10.6151
R731 B.n265 B.n264 10.6151
R732 B.n265 B.n98 10.6151
R733 B.n269 B.n98 10.6151
R734 B.n270 B.n269 10.6151
R735 B.n271 B.n270 10.6151
R736 B.n271 B.n96 10.6151
R737 B.n275 B.n96 10.6151
R738 B.n276 B.n275 10.6151
R739 B.n277 B.n276 10.6151
R740 B.n277 B.n94 10.6151
R741 B.n281 B.n94 10.6151
R742 B.n282 B.n281 10.6151
R743 B.n283 B.n282 10.6151
R744 B.n283 B.n92 10.6151
R745 B.n198 B.n197 10.6151
R746 B.n197 B.n126 10.6151
R747 B.n193 B.n126 10.6151
R748 B.n193 B.n192 10.6151
R749 B.n192 B.n191 10.6151
R750 B.n191 B.n128 10.6151
R751 B.n187 B.n128 10.6151
R752 B.n187 B.n186 10.6151
R753 B.n186 B.n185 10.6151
R754 B.n185 B.n130 10.6151
R755 B.n181 B.n130 10.6151
R756 B.n181 B.n180 10.6151
R757 B.n180 B.n179 10.6151
R758 B.n179 B.n132 10.6151
R759 B.n175 B.n132 10.6151
R760 B.n175 B.n174 10.6151
R761 B.n174 B.n173 10.6151
R762 B.n173 B.n134 10.6151
R763 B.n169 B.n134 10.6151
R764 B.n169 B.n168 10.6151
R765 B.n168 B.n167 10.6151
R766 B.n167 B.n136 10.6151
R767 B.n163 B.n136 10.6151
R768 B.n163 B.n162 10.6151
R769 B.n162 B.n161 10.6151
R770 B.n161 B.n138 10.6151
R771 B.n157 B.n138 10.6151
R772 B.n157 B.n156 10.6151
R773 B.n156 B.n155 10.6151
R774 B.n155 B.n140 10.6151
R775 B.n151 B.n140 10.6151
R776 B.n151 B.n150 10.6151
R777 B.n150 B.n149 10.6151
R778 B.n149 B.n142 10.6151
R779 B.n145 B.n142 10.6151
R780 B.n145 B.n144 10.6151
R781 B.n144 B.n0 10.6151
R782 B.n543 B.n1 10.6151
R783 B.n543 B.n542 10.6151
R784 B.n542 B.n541 10.6151
R785 B.n541 B.n4 10.6151
R786 B.n537 B.n4 10.6151
R787 B.n537 B.n536 10.6151
R788 B.n536 B.n535 10.6151
R789 B.n535 B.n6 10.6151
R790 B.n531 B.n6 10.6151
R791 B.n531 B.n530 10.6151
R792 B.n530 B.n529 10.6151
R793 B.n529 B.n8 10.6151
R794 B.n525 B.n8 10.6151
R795 B.n525 B.n524 10.6151
R796 B.n524 B.n523 10.6151
R797 B.n523 B.n10 10.6151
R798 B.n519 B.n10 10.6151
R799 B.n519 B.n518 10.6151
R800 B.n518 B.n517 10.6151
R801 B.n517 B.n12 10.6151
R802 B.n513 B.n12 10.6151
R803 B.n513 B.n512 10.6151
R804 B.n512 B.n511 10.6151
R805 B.n511 B.n14 10.6151
R806 B.n507 B.n14 10.6151
R807 B.n507 B.n506 10.6151
R808 B.n506 B.n505 10.6151
R809 B.n505 B.n16 10.6151
R810 B.n501 B.n16 10.6151
R811 B.n501 B.n500 10.6151
R812 B.n500 B.n499 10.6151
R813 B.n499 B.n18 10.6151
R814 B.n495 B.n18 10.6151
R815 B.n495 B.n494 10.6151
R816 B.n494 B.n493 10.6151
R817 B.n493 B.n20 10.6151
R818 B.n489 B.n20 10.6151
R819 B.n452 B.n451 6.5566
R820 B.n439 B.n438 6.5566
R821 B.n236 B.n235 6.5566
R822 B.n248 B.n106 6.5566
R823 B.n453 B.n452 4.05904
R824 B.n438 B.n437 4.05904
R825 B.n235 B.n234 4.05904
R826 B.n251 B.n106 4.05904
R827 B.n547 B.n0 2.81026
R828 B.n547 B.n1 2.81026
R829 VN.n25 VN.n14 161.3
R830 VN.n24 VN.n23 161.3
R831 VN.n22 VN.n15 161.3
R832 VN.n21 VN.n20 161.3
R833 VN.n19 VN.n16 161.3
R834 VN.n11 VN.n0 161.3
R835 VN.n10 VN.n9 161.3
R836 VN.n8 VN.n1 161.3
R837 VN.n7 VN.n6 161.3
R838 VN.n5 VN.n2 161.3
R839 VN.n3 VN.t2 96.179
R840 VN.n17 VN.t3 96.179
R841 VN.n13 VN.n12 96.1531
R842 VN.n27 VN.n26 96.1531
R843 VN.n4 VN.t4 63.3987
R844 VN.n12 VN.t1 63.3987
R845 VN.n18 VN.t5 63.3987
R846 VN.n26 VN.t0 63.3987
R847 VN.n4 VN.n3 59.4177
R848 VN.n18 VN.n17 59.4177
R849 VN.n10 VN.n1 42.999
R850 VN.n24 VN.n15 42.999
R851 VN VN.n27 42.7974
R852 VN.n6 VN.n1 38.1551
R853 VN.n20 VN.n15 38.1551
R854 VN.n6 VN.n5 24.5923
R855 VN.n11 VN.n10 24.5923
R856 VN.n20 VN.n19 24.5923
R857 VN.n25 VN.n24 24.5923
R858 VN.n12 VN.n11 14.7556
R859 VN.n26 VN.n25 14.7556
R860 VN.n5 VN.n4 12.2964
R861 VN.n19 VN.n18 12.2964
R862 VN.n17 VN.n16 9.46545
R863 VN.n3 VN.n2 9.46545
R864 VN.n27 VN.n14 0.278335
R865 VN.n13 VN.n0 0.278335
R866 VN.n23 VN.n14 0.189894
R867 VN.n23 VN.n22 0.189894
R868 VN.n22 VN.n21 0.189894
R869 VN.n21 VN.n16 0.189894
R870 VN.n7 VN.n2 0.189894
R871 VN.n8 VN.n7 0.189894
R872 VN.n9 VN.n8 0.189894
R873 VN.n9 VN.n0 0.189894
R874 VN VN.n13 0.153485
R875 VTAIL.n126 VTAIL.n125 756.745
R876 VTAIL.n30 VTAIL.n29 756.745
R877 VTAIL.n96 VTAIL.n95 756.745
R878 VTAIL.n64 VTAIL.n63 756.745
R879 VTAIL.n109 VTAIL.n108 585
R880 VTAIL.n111 VTAIL.n110 585
R881 VTAIL.n104 VTAIL.n103 585
R882 VTAIL.n117 VTAIL.n116 585
R883 VTAIL.n119 VTAIL.n118 585
R884 VTAIL.n100 VTAIL.n99 585
R885 VTAIL.n125 VTAIL.n124 585
R886 VTAIL.n13 VTAIL.n12 585
R887 VTAIL.n15 VTAIL.n14 585
R888 VTAIL.n8 VTAIL.n7 585
R889 VTAIL.n21 VTAIL.n20 585
R890 VTAIL.n23 VTAIL.n22 585
R891 VTAIL.n4 VTAIL.n3 585
R892 VTAIL.n29 VTAIL.n28 585
R893 VTAIL.n95 VTAIL.n94 585
R894 VTAIL.n70 VTAIL.n69 585
R895 VTAIL.n89 VTAIL.n88 585
R896 VTAIL.n87 VTAIL.n86 585
R897 VTAIL.n74 VTAIL.n73 585
R898 VTAIL.n81 VTAIL.n80 585
R899 VTAIL.n79 VTAIL.n78 585
R900 VTAIL.n63 VTAIL.n62 585
R901 VTAIL.n38 VTAIL.n37 585
R902 VTAIL.n57 VTAIL.n56 585
R903 VTAIL.n55 VTAIL.n54 585
R904 VTAIL.n42 VTAIL.n41 585
R905 VTAIL.n49 VTAIL.n48 585
R906 VTAIL.n47 VTAIL.n46 585
R907 VTAIL.n107 VTAIL.t5 329.175
R908 VTAIL.n11 VTAIL.t3 329.175
R909 VTAIL.n77 VTAIL.t2 329.175
R910 VTAIL.n45 VTAIL.t9 329.175
R911 VTAIL.n110 VTAIL.n109 171.744
R912 VTAIL.n110 VTAIL.n103 171.744
R913 VTAIL.n117 VTAIL.n103 171.744
R914 VTAIL.n118 VTAIL.n117 171.744
R915 VTAIL.n118 VTAIL.n99 171.744
R916 VTAIL.n125 VTAIL.n99 171.744
R917 VTAIL.n14 VTAIL.n13 171.744
R918 VTAIL.n14 VTAIL.n7 171.744
R919 VTAIL.n21 VTAIL.n7 171.744
R920 VTAIL.n22 VTAIL.n21 171.744
R921 VTAIL.n22 VTAIL.n3 171.744
R922 VTAIL.n29 VTAIL.n3 171.744
R923 VTAIL.n95 VTAIL.n69 171.744
R924 VTAIL.n88 VTAIL.n69 171.744
R925 VTAIL.n88 VTAIL.n87 171.744
R926 VTAIL.n87 VTAIL.n73 171.744
R927 VTAIL.n80 VTAIL.n73 171.744
R928 VTAIL.n80 VTAIL.n79 171.744
R929 VTAIL.n63 VTAIL.n37 171.744
R930 VTAIL.n56 VTAIL.n37 171.744
R931 VTAIL.n56 VTAIL.n55 171.744
R932 VTAIL.n55 VTAIL.n41 171.744
R933 VTAIL.n48 VTAIL.n41 171.744
R934 VTAIL.n48 VTAIL.n47 171.744
R935 VTAIL.n109 VTAIL.t5 85.8723
R936 VTAIL.n13 VTAIL.t3 85.8723
R937 VTAIL.n79 VTAIL.t2 85.8723
R938 VTAIL.n47 VTAIL.t9 85.8723
R939 VTAIL.n67 VTAIL.n66 78.822
R940 VTAIL.n35 VTAIL.n34 78.822
R941 VTAIL.n1 VTAIL.n0 78.821
R942 VTAIL.n33 VTAIL.n32 78.821
R943 VTAIL.n127 VTAIL.n126 34.9005
R944 VTAIL.n31 VTAIL.n30 34.9005
R945 VTAIL.n97 VTAIL.n96 34.9005
R946 VTAIL.n65 VTAIL.n64 34.9005
R947 VTAIL.n35 VTAIL.n33 21.7979
R948 VTAIL.n127 VTAIL.n97 19.5996
R949 VTAIL.n124 VTAIL.n98 12.0247
R950 VTAIL.n28 VTAIL.n2 12.0247
R951 VTAIL.n94 VTAIL.n68 12.0247
R952 VTAIL.n62 VTAIL.n36 12.0247
R953 VTAIL.n123 VTAIL.n100 11.249
R954 VTAIL.n27 VTAIL.n4 11.249
R955 VTAIL.n93 VTAIL.n70 11.249
R956 VTAIL.n61 VTAIL.n38 11.249
R957 VTAIL.n108 VTAIL.n107 10.722
R958 VTAIL.n12 VTAIL.n11 10.722
R959 VTAIL.n78 VTAIL.n77 10.722
R960 VTAIL.n46 VTAIL.n45 10.722
R961 VTAIL.n120 VTAIL.n119 10.4732
R962 VTAIL.n24 VTAIL.n23 10.4732
R963 VTAIL.n90 VTAIL.n89 10.4732
R964 VTAIL.n58 VTAIL.n57 10.4732
R965 VTAIL.n116 VTAIL.n102 9.69747
R966 VTAIL.n20 VTAIL.n6 9.69747
R967 VTAIL.n86 VTAIL.n72 9.69747
R968 VTAIL.n54 VTAIL.n40 9.69747
R969 VTAIL.n122 VTAIL.n98 9.45567
R970 VTAIL.n26 VTAIL.n2 9.45567
R971 VTAIL.n92 VTAIL.n68 9.45567
R972 VTAIL.n60 VTAIL.n36 9.45567
R973 VTAIL.n106 VTAIL.n105 9.3005
R974 VTAIL.n113 VTAIL.n112 9.3005
R975 VTAIL.n115 VTAIL.n114 9.3005
R976 VTAIL.n102 VTAIL.n101 9.3005
R977 VTAIL.n121 VTAIL.n120 9.3005
R978 VTAIL.n123 VTAIL.n122 9.3005
R979 VTAIL.n10 VTAIL.n9 9.3005
R980 VTAIL.n17 VTAIL.n16 9.3005
R981 VTAIL.n19 VTAIL.n18 9.3005
R982 VTAIL.n6 VTAIL.n5 9.3005
R983 VTAIL.n25 VTAIL.n24 9.3005
R984 VTAIL.n27 VTAIL.n26 9.3005
R985 VTAIL.n93 VTAIL.n92 9.3005
R986 VTAIL.n91 VTAIL.n90 9.3005
R987 VTAIL.n72 VTAIL.n71 9.3005
R988 VTAIL.n85 VTAIL.n84 9.3005
R989 VTAIL.n83 VTAIL.n82 9.3005
R990 VTAIL.n76 VTAIL.n75 9.3005
R991 VTAIL.n51 VTAIL.n50 9.3005
R992 VTAIL.n53 VTAIL.n52 9.3005
R993 VTAIL.n40 VTAIL.n39 9.3005
R994 VTAIL.n59 VTAIL.n58 9.3005
R995 VTAIL.n61 VTAIL.n60 9.3005
R996 VTAIL.n44 VTAIL.n43 9.3005
R997 VTAIL.n115 VTAIL.n104 8.92171
R998 VTAIL.n19 VTAIL.n8 8.92171
R999 VTAIL.n85 VTAIL.n74 8.92171
R1000 VTAIL.n53 VTAIL.n42 8.92171
R1001 VTAIL.n112 VTAIL.n111 8.14595
R1002 VTAIL.n16 VTAIL.n15 8.14595
R1003 VTAIL.n82 VTAIL.n81 8.14595
R1004 VTAIL.n50 VTAIL.n49 8.14595
R1005 VTAIL.n108 VTAIL.n106 7.3702
R1006 VTAIL.n12 VTAIL.n10 7.3702
R1007 VTAIL.n78 VTAIL.n76 7.3702
R1008 VTAIL.n46 VTAIL.n44 7.3702
R1009 VTAIL.n111 VTAIL.n106 5.81868
R1010 VTAIL.n15 VTAIL.n10 5.81868
R1011 VTAIL.n81 VTAIL.n76 5.81868
R1012 VTAIL.n49 VTAIL.n44 5.81868
R1013 VTAIL.n0 VTAIL.t7 5.56642
R1014 VTAIL.n0 VTAIL.t6 5.56642
R1015 VTAIL.n32 VTAIL.t11 5.56642
R1016 VTAIL.n32 VTAIL.t10 5.56642
R1017 VTAIL.n66 VTAIL.t1 5.56642
R1018 VTAIL.n66 VTAIL.t0 5.56642
R1019 VTAIL.n34 VTAIL.t4 5.56642
R1020 VTAIL.n34 VTAIL.t8 5.56642
R1021 VTAIL.n112 VTAIL.n104 5.04292
R1022 VTAIL.n16 VTAIL.n8 5.04292
R1023 VTAIL.n82 VTAIL.n74 5.04292
R1024 VTAIL.n50 VTAIL.n42 5.04292
R1025 VTAIL.n116 VTAIL.n115 4.26717
R1026 VTAIL.n20 VTAIL.n19 4.26717
R1027 VTAIL.n86 VTAIL.n85 4.26717
R1028 VTAIL.n54 VTAIL.n53 4.26717
R1029 VTAIL.n119 VTAIL.n102 3.49141
R1030 VTAIL.n23 VTAIL.n6 3.49141
R1031 VTAIL.n89 VTAIL.n72 3.49141
R1032 VTAIL.n57 VTAIL.n40 3.49141
R1033 VTAIL.n120 VTAIL.n100 2.71565
R1034 VTAIL.n24 VTAIL.n4 2.71565
R1035 VTAIL.n90 VTAIL.n70 2.71565
R1036 VTAIL.n58 VTAIL.n38 2.71565
R1037 VTAIL.n107 VTAIL.n105 2.4147
R1038 VTAIL.n11 VTAIL.n9 2.4147
R1039 VTAIL.n77 VTAIL.n75 2.4147
R1040 VTAIL.n45 VTAIL.n43 2.4147
R1041 VTAIL.n65 VTAIL.n35 2.19878
R1042 VTAIL.n97 VTAIL.n67 2.19878
R1043 VTAIL.n33 VTAIL.n31 2.19878
R1044 VTAIL.n124 VTAIL.n123 1.93989
R1045 VTAIL.n28 VTAIL.n27 1.93989
R1046 VTAIL.n94 VTAIL.n93 1.93989
R1047 VTAIL.n62 VTAIL.n61 1.93989
R1048 VTAIL VTAIL.n127 1.59102
R1049 VTAIL.n67 VTAIL.n65 1.56947
R1050 VTAIL.n31 VTAIL.n1 1.56947
R1051 VTAIL.n126 VTAIL.n98 1.16414
R1052 VTAIL.n30 VTAIL.n2 1.16414
R1053 VTAIL.n96 VTAIL.n68 1.16414
R1054 VTAIL.n64 VTAIL.n36 1.16414
R1055 VTAIL VTAIL.n1 0.608259
R1056 VTAIL.n113 VTAIL.n105 0.155672
R1057 VTAIL.n114 VTAIL.n113 0.155672
R1058 VTAIL.n114 VTAIL.n101 0.155672
R1059 VTAIL.n121 VTAIL.n101 0.155672
R1060 VTAIL.n122 VTAIL.n121 0.155672
R1061 VTAIL.n17 VTAIL.n9 0.155672
R1062 VTAIL.n18 VTAIL.n17 0.155672
R1063 VTAIL.n18 VTAIL.n5 0.155672
R1064 VTAIL.n25 VTAIL.n5 0.155672
R1065 VTAIL.n26 VTAIL.n25 0.155672
R1066 VTAIL.n92 VTAIL.n91 0.155672
R1067 VTAIL.n91 VTAIL.n71 0.155672
R1068 VTAIL.n84 VTAIL.n71 0.155672
R1069 VTAIL.n84 VTAIL.n83 0.155672
R1070 VTAIL.n83 VTAIL.n75 0.155672
R1071 VTAIL.n60 VTAIL.n59 0.155672
R1072 VTAIL.n59 VTAIL.n39 0.155672
R1073 VTAIL.n52 VTAIL.n39 0.155672
R1074 VTAIL.n52 VTAIL.n51 0.155672
R1075 VTAIL.n51 VTAIL.n43 0.155672
R1076 VDD2.n59 VDD2.n58 756.745
R1077 VDD2.n28 VDD2.n27 756.745
R1078 VDD2.n58 VDD2.n57 585
R1079 VDD2.n33 VDD2.n32 585
R1080 VDD2.n52 VDD2.n51 585
R1081 VDD2.n50 VDD2.n49 585
R1082 VDD2.n37 VDD2.n36 585
R1083 VDD2.n44 VDD2.n43 585
R1084 VDD2.n42 VDD2.n41 585
R1085 VDD2.n11 VDD2.n10 585
R1086 VDD2.n13 VDD2.n12 585
R1087 VDD2.n6 VDD2.n5 585
R1088 VDD2.n19 VDD2.n18 585
R1089 VDD2.n21 VDD2.n20 585
R1090 VDD2.n2 VDD2.n1 585
R1091 VDD2.n27 VDD2.n26 585
R1092 VDD2.n9 VDD2.t3 329.175
R1093 VDD2.n40 VDD2.t5 329.175
R1094 VDD2.n58 VDD2.n32 171.744
R1095 VDD2.n51 VDD2.n32 171.744
R1096 VDD2.n51 VDD2.n50 171.744
R1097 VDD2.n50 VDD2.n36 171.744
R1098 VDD2.n43 VDD2.n36 171.744
R1099 VDD2.n43 VDD2.n42 171.744
R1100 VDD2.n12 VDD2.n11 171.744
R1101 VDD2.n12 VDD2.n5 171.744
R1102 VDD2.n19 VDD2.n5 171.744
R1103 VDD2.n20 VDD2.n19 171.744
R1104 VDD2.n20 VDD2.n1 171.744
R1105 VDD2.n27 VDD2.n1 171.744
R1106 VDD2.n30 VDD2.n29 95.994
R1107 VDD2 VDD2.n61 95.991
R1108 VDD2.n42 VDD2.t5 85.8723
R1109 VDD2.n11 VDD2.t3 85.8723
R1110 VDD2.n30 VDD2.n28 53.1726
R1111 VDD2.n60 VDD2.n59 51.5793
R1112 VDD2.n60 VDD2.n30 35.8942
R1113 VDD2.n57 VDD2.n31 12.0247
R1114 VDD2.n26 VDD2.n0 12.0247
R1115 VDD2.n56 VDD2.n33 11.249
R1116 VDD2.n25 VDD2.n2 11.249
R1117 VDD2.n10 VDD2.n9 10.722
R1118 VDD2.n41 VDD2.n40 10.722
R1119 VDD2.n53 VDD2.n52 10.4732
R1120 VDD2.n22 VDD2.n21 10.4732
R1121 VDD2.n49 VDD2.n35 9.69747
R1122 VDD2.n18 VDD2.n4 9.69747
R1123 VDD2.n55 VDD2.n31 9.45567
R1124 VDD2.n24 VDD2.n0 9.45567
R1125 VDD2.n46 VDD2.n45 9.3005
R1126 VDD2.n48 VDD2.n47 9.3005
R1127 VDD2.n35 VDD2.n34 9.3005
R1128 VDD2.n54 VDD2.n53 9.3005
R1129 VDD2.n56 VDD2.n55 9.3005
R1130 VDD2.n39 VDD2.n38 9.3005
R1131 VDD2.n8 VDD2.n7 9.3005
R1132 VDD2.n15 VDD2.n14 9.3005
R1133 VDD2.n17 VDD2.n16 9.3005
R1134 VDD2.n4 VDD2.n3 9.3005
R1135 VDD2.n23 VDD2.n22 9.3005
R1136 VDD2.n25 VDD2.n24 9.3005
R1137 VDD2.n48 VDD2.n37 8.92171
R1138 VDD2.n17 VDD2.n6 8.92171
R1139 VDD2.n45 VDD2.n44 8.14595
R1140 VDD2.n14 VDD2.n13 8.14595
R1141 VDD2.n41 VDD2.n39 7.3702
R1142 VDD2.n10 VDD2.n8 7.3702
R1143 VDD2.n44 VDD2.n39 5.81868
R1144 VDD2.n13 VDD2.n8 5.81868
R1145 VDD2.n61 VDD2.t0 5.56642
R1146 VDD2.n61 VDD2.t2 5.56642
R1147 VDD2.n29 VDD2.t1 5.56642
R1148 VDD2.n29 VDD2.t4 5.56642
R1149 VDD2.n45 VDD2.n37 5.04292
R1150 VDD2.n14 VDD2.n6 5.04292
R1151 VDD2.n49 VDD2.n48 4.26717
R1152 VDD2.n18 VDD2.n17 4.26717
R1153 VDD2.n52 VDD2.n35 3.49141
R1154 VDD2.n21 VDD2.n4 3.49141
R1155 VDD2.n53 VDD2.n33 2.71565
R1156 VDD2.n22 VDD2.n2 2.71565
R1157 VDD2.n9 VDD2.n7 2.4147
R1158 VDD2.n40 VDD2.n38 2.4147
R1159 VDD2.n57 VDD2.n56 1.93989
R1160 VDD2.n26 VDD2.n25 1.93989
R1161 VDD2 VDD2.n60 1.7074
R1162 VDD2.n59 VDD2.n31 1.16414
R1163 VDD2.n28 VDD2.n0 1.16414
R1164 VDD2.n55 VDD2.n54 0.155672
R1165 VDD2.n54 VDD2.n34 0.155672
R1166 VDD2.n47 VDD2.n34 0.155672
R1167 VDD2.n47 VDD2.n46 0.155672
R1168 VDD2.n46 VDD2.n38 0.155672
R1169 VDD2.n15 VDD2.n7 0.155672
R1170 VDD2.n16 VDD2.n15 0.155672
R1171 VDD2.n16 VDD2.n3 0.155672
R1172 VDD2.n23 VDD2.n3 0.155672
R1173 VDD2.n24 VDD2.n23 0.155672
R1174 VP.n11 VP.n8 161.3
R1175 VP.n13 VP.n12 161.3
R1176 VP.n14 VP.n7 161.3
R1177 VP.n16 VP.n15 161.3
R1178 VP.n17 VP.n6 161.3
R1179 VP.n36 VP.n0 161.3
R1180 VP.n35 VP.n34 161.3
R1181 VP.n33 VP.n1 161.3
R1182 VP.n32 VP.n31 161.3
R1183 VP.n30 VP.n2 161.3
R1184 VP.n28 VP.n27 161.3
R1185 VP.n26 VP.n3 161.3
R1186 VP.n25 VP.n24 161.3
R1187 VP.n23 VP.n4 161.3
R1188 VP.n22 VP.n21 161.3
R1189 VP.n9 VP.t2 96.179
R1190 VP.n20 VP.n5 96.1531
R1191 VP.n38 VP.n37 96.1531
R1192 VP.n19 VP.n18 96.1531
R1193 VP.n5 VP.t5 63.3987
R1194 VP.n29 VP.t3 63.3987
R1195 VP.n37 VP.t1 63.3987
R1196 VP.n18 VP.t0 63.3987
R1197 VP.n10 VP.t4 63.3987
R1198 VP.n10 VP.n9 59.4177
R1199 VP.n24 VP.n23 42.999
R1200 VP.n35 VP.n1 42.999
R1201 VP.n16 VP.n7 42.999
R1202 VP.n20 VP.n19 42.5186
R1203 VP.n24 VP.n3 38.1551
R1204 VP.n31 VP.n1 38.1551
R1205 VP.n12 VP.n7 38.1551
R1206 VP.n23 VP.n22 24.5923
R1207 VP.n28 VP.n3 24.5923
R1208 VP.n31 VP.n30 24.5923
R1209 VP.n36 VP.n35 24.5923
R1210 VP.n17 VP.n16 24.5923
R1211 VP.n12 VP.n11 24.5923
R1212 VP.n22 VP.n5 14.7556
R1213 VP.n37 VP.n36 14.7556
R1214 VP.n18 VP.n17 14.7556
R1215 VP.n29 VP.n28 12.2964
R1216 VP.n30 VP.n29 12.2964
R1217 VP.n11 VP.n10 12.2964
R1218 VP.n9 VP.n8 9.46545
R1219 VP.n19 VP.n6 0.278335
R1220 VP.n21 VP.n20 0.278335
R1221 VP.n38 VP.n0 0.278335
R1222 VP.n13 VP.n8 0.189894
R1223 VP.n14 VP.n13 0.189894
R1224 VP.n15 VP.n14 0.189894
R1225 VP.n15 VP.n6 0.189894
R1226 VP.n21 VP.n4 0.189894
R1227 VP.n25 VP.n4 0.189894
R1228 VP.n26 VP.n25 0.189894
R1229 VP.n27 VP.n26 0.189894
R1230 VP.n27 VP.n2 0.189894
R1231 VP.n32 VP.n2 0.189894
R1232 VP.n33 VP.n32 0.189894
R1233 VP.n34 VP.n33 0.189894
R1234 VP.n34 VP.n0 0.189894
R1235 VP VP.n38 0.153485
R1236 VDD1.n28 VDD1.n27 756.745
R1237 VDD1.n57 VDD1.n56 756.745
R1238 VDD1.n27 VDD1.n26 585
R1239 VDD1.n2 VDD1.n1 585
R1240 VDD1.n21 VDD1.n20 585
R1241 VDD1.n19 VDD1.n18 585
R1242 VDD1.n6 VDD1.n5 585
R1243 VDD1.n13 VDD1.n12 585
R1244 VDD1.n11 VDD1.n10 585
R1245 VDD1.n40 VDD1.n39 585
R1246 VDD1.n42 VDD1.n41 585
R1247 VDD1.n35 VDD1.n34 585
R1248 VDD1.n48 VDD1.n47 585
R1249 VDD1.n50 VDD1.n49 585
R1250 VDD1.n31 VDD1.n30 585
R1251 VDD1.n56 VDD1.n55 585
R1252 VDD1.n38 VDD1.t0 329.175
R1253 VDD1.n9 VDD1.t3 329.175
R1254 VDD1.n27 VDD1.n1 171.744
R1255 VDD1.n20 VDD1.n1 171.744
R1256 VDD1.n20 VDD1.n19 171.744
R1257 VDD1.n19 VDD1.n5 171.744
R1258 VDD1.n12 VDD1.n5 171.744
R1259 VDD1.n12 VDD1.n11 171.744
R1260 VDD1.n41 VDD1.n40 171.744
R1261 VDD1.n41 VDD1.n34 171.744
R1262 VDD1.n48 VDD1.n34 171.744
R1263 VDD1.n49 VDD1.n48 171.744
R1264 VDD1.n49 VDD1.n30 171.744
R1265 VDD1.n56 VDD1.n30 171.744
R1266 VDD1.n59 VDD1.n58 95.994
R1267 VDD1.n61 VDD1.n60 95.4997
R1268 VDD1.n11 VDD1.t3 85.8723
R1269 VDD1.n40 VDD1.t0 85.8723
R1270 VDD1 VDD1.n28 53.2862
R1271 VDD1.n59 VDD1.n57 53.1726
R1272 VDD1.n61 VDD1.n59 37.5763
R1273 VDD1.n26 VDD1.n0 12.0247
R1274 VDD1.n55 VDD1.n29 12.0247
R1275 VDD1.n25 VDD1.n2 11.249
R1276 VDD1.n54 VDD1.n31 11.249
R1277 VDD1.n39 VDD1.n38 10.722
R1278 VDD1.n10 VDD1.n9 10.722
R1279 VDD1.n22 VDD1.n21 10.4732
R1280 VDD1.n51 VDD1.n50 10.4732
R1281 VDD1.n18 VDD1.n4 9.69747
R1282 VDD1.n47 VDD1.n33 9.69747
R1283 VDD1.n24 VDD1.n0 9.45567
R1284 VDD1.n53 VDD1.n29 9.45567
R1285 VDD1.n15 VDD1.n14 9.3005
R1286 VDD1.n17 VDD1.n16 9.3005
R1287 VDD1.n4 VDD1.n3 9.3005
R1288 VDD1.n23 VDD1.n22 9.3005
R1289 VDD1.n25 VDD1.n24 9.3005
R1290 VDD1.n8 VDD1.n7 9.3005
R1291 VDD1.n37 VDD1.n36 9.3005
R1292 VDD1.n44 VDD1.n43 9.3005
R1293 VDD1.n46 VDD1.n45 9.3005
R1294 VDD1.n33 VDD1.n32 9.3005
R1295 VDD1.n52 VDD1.n51 9.3005
R1296 VDD1.n54 VDD1.n53 9.3005
R1297 VDD1.n17 VDD1.n6 8.92171
R1298 VDD1.n46 VDD1.n35 8.92171
R1299 VDD1.n14 VDD1.n13 8.14595
R1300 VDD1.n43 VDD1.n42 8.14595
R1301 VDD1.n10 VDD1.n8 7.3702
R1302 VDD1.n39 VDD1.n37 7.3702
R1303 VDD1.n13 VDD1.n8 5.81868
R1304 VDD1.n42 VDD1.n37 5.81868
R1305 VDD1.n60 VDD1.t1 5.56642
R1306 VDD1.n60 VDD1.t5 5.56642
R1307 VDD1.n58 VDD1.t2 5.56642
R1308 VDD1.n58 VDD1.t4 5.56642
R1309 VDD1.n14 VDD1.n6 5.04292
R1310 VDD1.n43 VDD1.n35 5.04292
R1311 VDD1.n18 VDD1.n17 4.26717
R1312 VDD1.n47 VDD1.n46 4.26717
R1313 VDD1.n21 VDD1.n4 3.49141
R1314 VDD1.n50 VDD1.n33 3.49141
R1315 VDD1.n22 VDD1.n2 2.71565
R1316 VDD1.n51 VDD1.n31 2.71565
R1317 VDD1.n38 VDD1.n36 2.4147
R1318 VDD1.n9 VDD1.n7 2.4147
R1319 VDD1.n26 VDD1.n25 1.93989
R1320 VDD1.n55 VDD1.n54 1.93989
R1321 VDD1.n28 VDD1.n0 1.16414
R1322 VDD1.n57 VDD1.n29 1.16414
R1323 VDD1 VDD1.n61 0.491879
R1324 VDD1.n24 VDD1.n23 0.155672
R1325 VDD1.n23 VDD1.n3 0.155672
R1326 VDD1.n16 VDD1.n3 0.155672
R1327 VDD1.n16 VDD1.n15 0.155672
R1328 VDD1.n15 VDD1.n7 0.155672
R1329 VDD1.n44 VDD1.n36 0.155672
R1330 VDD1.n45 VDD1.n44 0.155672
R1331 VDD1.n45 VDD1.n32 0.155672
R1332 VDD1.n52 VDD1.n32 0.155672
R1333 VDD1.n53 VDD1.n52 0.155672
C0 VP VN 5.41384f
C1 w_n3010_n2136# VDD1 1.76473f
C2 w_n3010_n2136# VDD2 1.83767f
C3 VTAIL B 2.18185f
C4 VDD1 VP 3.64146f
C5 VDD2 VP 0.425726f
C6 VDD1 VN 0.150373f
C7 VDD2 VN 3.36821f
C8 w_n3010_n2136# B 7.434081f
C9 VTAIL w_n3010_n2136# 2.06335f
C10 VDD1 VDD2 1.25693f
C11 B VP 1.65948f
C12 VTAIL VP 3.84572f
C13 B VN 1.01343f
C14 VTAIL VN 3.83151f
C15 VDD1 B 1.51098f
C16 VDD2 B 1.57599f
C17 VTAIL VDD1 5.32573f
C18 w_n3010_n2136# VP 5.88753f
C19 VTAIL VDD2 5.37522f
C20 w_n3010_n2136# VN 5.49944f
C21 VDD2 VSUBS 1.348453f
C22 VDD1 VSUBS 1.429535f
C23 VTAIL VSUBS 0.634939f
C24 VN VSUBS 5.19312f
C25 VP VSUBS 2.278127f
C26 B VSUBS 3.739241f
C27 w_n3010_n2136# VSUBS 80.2948f
C28 VDD1.n0 VSUBS 0.012451f
C29 VDD1.n1 VSUBS 0.028049f
C30 VDD1.n2 VSUBS 0.012565f
C31 VDD1.n3 VSUBS 0.022083f
C32 VDD1.n4 VSUBS 0.011867f
C33 VDD1.n5 VSUBS 0.028049f
C34 VDD1.n6 VSUBS 0.012565f
C35 VDD1.n7 VSUBS 0.488172f
C36 VDD1.n8 VSUBS 0.011867f
C37 VDD1.t3 VSUBS 0.060436f
C38 VDD1.n9 VSUBS 0.112774f
C39 VDD1.n10 VSUBS 0.021091f
C40 VDD1.n11 VSUBS 0.021036f
C41 VDD1.n12 VSUBS 0.028049f
C42 VDD1.n13 VSUBS 0.012565f
C43 VDD1.n14 VSUBS 0.011867f
C44 VDD1.n15 VSUBS 0.022083f
C45 VDD1.n16 VSUBS 0.022083f
C46 VDD1.n17 VSUBS 0.011867f
C47 VDD1.n18 VSUBS 0.012565f
C48 VDD1.n19 VSUBS 0.028049f
C49 VDD1.n20 VSUBS 0.028049f
C50 VDD1.n21 VSUBS 0.012565f
C51 VDD1.n22 VSUBS 0.011867f
C52 VDD1.n23 VSUBS 0.022083f
C53 VDD1.n24 VSUBS 0.057078f
C54 VDD1.n25 VSUBS 0.011867f
C55 VDD1.n26 VSUBS 0.012565f
C56 VDD1.n27 VSUBS 0.062486f
C57 VDD1.n28 VSUBS 0.06246f
C58 VDD1.n29 VSUBS 0.012451f
C59 VDD1.n30 VSUBS 0.028049f
C60 VDD1.n31 VSUBS 0.012565f
C61 VDD1.n32 VSUBS 0.022083f
C62 VDD1.n33 VSUBS 0.011867f
C63 VDD1.n34 VSUBS 0.028049f
C64 VDD1.n35 VSUBS 0.012565f
C65 VDD1.n36 VSUBS 0.488172f
C66 VDD1.n37 VSUBS 0.011867f
C67 VDD1.t0 VSUBS 0.060436f
C68 VDD1.n38 VSUBS 0.112774f
C69 VDD1.n39 VSUBS 0.021091f
C70 VDD1.n40 VSUBS 0.021036f
C71 VDD1.n41 VSUBS 0.028049f
C72 VDD1.n42 VSUBS 0.012565f
C73 VDD1.n43 VSUBS 0.011867f
C74 VDD1.n44 VSUBS 0.022083f
C75 VDD1.n45 VSUBS 0.022083f
C76 VDD1.n46 VSUBS 0.011867f
C77 VDD1.n47 VSUBS 0.012565f
C78 VDD1.n48 VSUBS 0.028049f
C79 VDD1.n49 VSUBS 0.028049f
C80 VDD1.n50 VSUBS 0.012565f
C81 VDD1.n51 VSUBS 0.011867f
C82 VDD1.n52 VSUBS 0.022083f
C83 VDD1.n53 VSUBS 0.057078f
C84 VDD1.n54 VSUBS 0.011867f
C85 VDD1.n55 VSUBS 0.012565f
C86 VDD1.n56 VSUBS 0.062486f
C87 VDD1.n57 VSUBS 0.061883f
C88 VDD1.t2 VSUBS 0.101914f
C89 VDD1.t4 VSUBS 0.101914f
C90 VDD1.n58 VSUBS 0.688781f
C91 VDD1.n59 VSUBS 2.14948f
C92 VDD1.t1 VSUBS 0.101914f
C93 VDD1.t5 VSUBS 0.101914f
C94 VDD1.n60 VSUBS 0.685991f
C95 VDD1.n61 VSUBS 2.10488f
C96 VP.n0 VSUBS 0.056014f
C97 VP.t1 VSUBS 1.45565f
C98 VP.n1 VSUBS 0.034657f
C99 VP.n2 VSUBS 0.042489f
C100 VP.t3 VSUBS 1.45565f
C101 VP.n3 VSUBS 0.084876f
C102 VP.n4 VSUBS 0.042489f
C103 VP.t5 VSUBS 1.45565f
C104 VP.n5 VSUBS 0.684032f
C105 VP.n6 VSUBS 0.056014f
C106 VP.t0 VSUBS 1.45565f
C107 VP.n7 VSUBS 0.034657f
C108 VP.n8 VSUBS 0.362563f
C109 VP.t4 VSUBS 1.45565f
C110 VP.t2 VSUBS 1.72237f
C111 VP.n9 VSUBS 0.646986f
C112 VP.n10 VSUBS 0.663039f
C113 VP.n11 VSUBS 0.059343f
C114 VP.n12 VSUBS 0.084876f
C115 VP.n13 VSUBS 0.042489f
C116 VP.n14 VSUBS 0.042489f
C117 VP.n15 VSUBS 0.042489f
C118 VP.n16 VSUBS 0.082788f
C119 VP.n17 VSUBS 0.063233f
C120 VP.n18 VSUBS 0.684032f
C121 VP.n19 VSUBS 1.83332f
C122 VP.n20 VSUBS 1.86934f
C123 VP.n21 VSUBS 0.056014f
C124 VP.n22 VSUBS 0.063233f
C125 VP.n23 VSUBS 0.082788f
C126 VP.n24 VSUBS 0.034657f
C127 VP.n25 VSUBS 0.042489f
C128 VP.n26 VSUBS 0.042489f
C129 VP.n27 VSUBS 0.042489f
C130 VP.n28 VSUBS 0.059343f
C131 VP.n29 VSUBS 0.553487f
C132 VP.n30 VSUBS 0.059343f
C133 VP.n31 VSUBS 0.084876f
C134 VP.n32 VSUBS 0.042489f
C135 VP.n33 VSUBS 0.042489f
C136 VP.n34 VSUBS 0.042489f
C137 VP.n35 VSUBS 0.082788f
C138 VP.n36 VSUBS 0.063233f
C139 VP.n37 VSUBS 0.684032f
C140 VP.n38 VSUBS 0.059432f
C141 VDD2.n0 VSUBS 0.012425f
C142 VDD2.n1 VSUBS 0.02799f
C143 VDD2.n2 VSUBS 0.012539f
C144 VDD2.n3 VSUBS 0.022037f
C145 VDD2.n4 VSUBS 0.011842f
C146 VDD2.n5 VSUBS 0.02799f
C147 VDD2.n6 VSUBS 0.012539f
C148 VDD2.n7 VSUBS 0.487151f
C149 VDD2.n8 VSUBS 0.011842f
C150 VDD2.t3 VSUBS 0.060309f
C151 VDD2.n9 VSUBS 0.112538f
C152 VDD2.n10 VSUBS 0.021046f
C153 VDD2.n11 VSUBS 0.020992f
C154 VDD2.n12 VSUBS 0.02799f
C155 VDD2.n13 VSUBS 0.012539f
C156 VDD2.n14 VSUBS 0.011842f
C157 VDD2.n15 VSUBS 0.022037f
C158 VDD2.n16 VSUBS 0.022037f
C159 VDD2.n17 VSUBS 0.011842f
C160 VDD2.n18 VSUBS 0.012539f
C161 VDD2.n19 VSUBS 0.02799f
C162 VDD2.n20 VSUBS 0.02799f
C163 VDD2.n21 VSUBS 0.012539f
C164 VDD2.n22 VSUBS 0.011842f
C165 VDD2.n23 VSUBS 0.022037f
C166 VDD2.n24 VSUBS 0.056959f
C167 VDD2.n25 VSUBS 0.011842f
C168 VDD2.n26 VSUBS 0.012539f
C169 VDD2.n27 VSUBS 0.062355f
C170 VDD2.n28 VSUBS 0.061754f
C171 VDD2.t1 VSUBS 0.101701f
C172 VDD2.t4 VSUBS 0.101701f
C173 VDD2.n29 VSUBS 0.687341f
C174 VDD2.n30 VSUBS 2.04888f
C175 VDD2.n31 VSUBS 0.012425f
C176 VDD2.n32 VSUBS 0.02799f
C177 VDD2.n33 VSUBS 0.012539f
C178 VDD2.n34 VSUBS 0.022037f
C179 VDD2.n35 VSUBS 0.011842f
C180 VDD2.n36 VSUBS 0.02799f
C181 VDD2.n37 VSUBS 0.012539f
C182 VDD2.n38 VSUBS 0.487151f
C183 VDD2.n39 VSUBS 0.011842f
C184 VDD2.t5 VSUBS 0.060309f
C185 VDD2.n40 VSUBS 0.112538f
C186 VDD2.n41 VSUBS 0.021046f
C187 VDD2.n42 VSUBS 0.020992f
C188 VDD2.n43 VSUBS 0.02799f
C189 VDD2.n44 VSUBS 0.012539f
C190 VDD2.n45 VSUBS 0.011842f
C191 VDD2.n46 VSUBS 0.022037f
C192 VDD2.n47 VSUBS 0.022037f
C193 VDD2.n48 VSUBS 0.011842f
C194 VDD2.n49 VSUBS 0.012539f
C195 VDD2.n50 VSUBS 0.02799f
C196 VDD2.n51 VSUBS 0.02799f
C197 VDD2.n52 VSUBS 0.012539f
C198 VDD2.n53 VSUBS 0.011842f
C199 VDD2.n54 VSUBS 0.022037f
C200 VDD2.n55 VSUBS 0.056959f
C201 VDD2.n56 VSUBS 0.011842f
C202 VDD2.n57 VSUBS 0.012539f
C203 VDD2.n58 VSUBS 0.062355f
C204 VDD2.n59 VSUBS 0.05701f
C205 VDD2.n60 VSUBS 1.74216f
C206 VDD2.t0 VSUBS 0.101701f
C207 VDD2.t2 VSUBS 0.101701f
C208 VDD2.n61 VSUBS 0.687317f
C209 VTAIL.t7 VSUBS 0.151892f
C210 VTAIL.t6 VSUBS 0.151892f
C211 VTAIL.n0 VSUBS 0.916527f
C212 VTAIL.n1 VSUBS 0.798615f
C213 VTAIL.n2 VSUBS 0.018556f
C214 VTAIL.n3 VSUBS 0.041804f
C215 VTAIL.n4 VSUBS 0.018726f
C216 VTAIL.n5 VSUBS 0.032913f
C217 VTAIL.n6 VSUBS 0.017686f
C218 VTAIL.n7 VSUBS 0.041804f
C219 VTAIL.n8 VSUBS 0.018726f
C220 VTAIL.n9 VSUBS 0.727571f
C221 VTAIL.n10 VSUBS 0.017686f
C222 VTAIL.t3 VSUBS 0.090073f
C223 VTAIL.n11 VSUBS 0.168078f
C224 VTAIL.n12 VSUBS 0.031434f
C225 VTAIL.n13 VSUBS 0.031353f
C226 VTAIL.n14 VSUBS 0.041804f
C227 VTAIL.n15 VSUBS 0.018726f
C228 VTAIL.n16 VSUBS 0.017686f
C229 VTAIL.n17 VSUBS 0.032913f
C230 VTAIL.n18 VSUBS 0.032913f
C231 VTAIL.n19 VSUBS 0.017686f
C232 VTAIL.n20 VSUBS 0.018726f
C233 VTAIL.n21 VSUBS 0.041804f
C234 VTAIL.n22 VSUBS 0.041804f
C235 VTAIL.n23 VSUBS 0.018726f
C236 VTAIL.n24 VSUBS 0.017686f
C237 VTAIL.n25 VSUBS 0.032913f
C238 VTAIL.n26 VSUBS 0.08507f
C239 VTAIL.n27 VSUBS 0.017686f
C240 VTAIL.n28 VSUBS 0.018726f
C241 VTAIL.n29 VSUBS 0.093129f
C242 VTAIL.n30 VSUBS 0.062466f
C243 VTAIL.n31 VSUBS 0.431199f
C244 VTAIL.t11 VSUBS 0.151892f
C245 VTAIL.t10 VSUBS 0.151892f
C246 VTAIL.n32 VSUBS 0.916527f
C247 VTAIL.n33 VSUBS 2.24818f
C248 VTAIL.t4 VSUBS 0.151892f
C249 VTAIL.t8 VSUBS 0.151892f
C250 VTAIL.n34 VSUBS 0.916531f
C251 VTAIL.n35 VSUBS 2.24818f
C252 VTAIL.n36 VSUBS 0.018556f
C253 VTAIL.n37 VSUBS 0.041804f
C254 VTAIL.n38 VSUBS 0.018726f
C255 VTAIL.n39 VSUBS 0.032913f
C256 VTAIL.n40 VSUBS 0.017686f
C257 VTAIL.n41 VSUBS 0.041804f
C258 VTAIL.n42 VSUBS 0.018726f
C259 VTAIL.n43 VSUBS 0.727571f
C260 VTAIL.n44 VSUBS 0.017686f
C261 VTAIL.t9 VSUBS 0.090073f
C262 VTAIL.n45 VSUBS 0.168078f
C263 VTAIL.n46 VSUBS 0.031434f
C264 VTAIL.n47 VSUBS 0.031353f
C265 VTAIL.n48 VSUBS 0.041804f
C266 VTAIL.n49 VSUBS 0.018726f
C267 VTAIL.n50 VSUBS 0.017686f
C268 VTAIL.n51 VSUBS 0.032913f
C269 VTAIL.n52 VSUBS 0.032913f
C270 VTAIL.n53 VSUBS 0.017686f
C271 VTAIL.n54 VSUBS 0.018726f
C272 VTAIL.n55 VSUBS 0.041804f
C273 VTAIL.n56 VSUBS 0.041804f
C274 VTAIL.n57 VSUBS 0.018726f
C275 VTAIL.n58 VSUBS 0.017686f
C276 VTAIL.n59 VSUBS 0.032913f
C277 VTAIL.n60 VSUBS 0.08507f
C278 VTAIL.n61 VSUBS 0.017686f
C279 VTAIL.n62 VSUBS 0.018726f
C280 VTAIL.n63 VSUBS 0.093129f
C281 VTAIL.n64 VSUBS 0.062466f
C282 VTAIL.n65 VSUBS 0.431199f
C283 VTAIL.t1 VSUBS 0.151892f
C284 VTAIL.t0 VSUBS 0.151892f
C285 VTAIL.n66 VSUBS 0.916531f
C286 VTAIL.n67 VSUBS 0.967292f
C287 VTAIL.n68 VSUBS 0.018556f
C288 VTAIL.n69 VSUBS 0.041804f
C289 VTAIL.n70 VSUBS 0.018726f
C290 VTAIL.n71 VSUBS 0.032913f
C291 VTAIL.n72 VSUBS 0.017686f
C292 VTAIL.n73 VSUBS 0.041804f
C293 VTAIL.n74 VSUBS 0.018726f
C294 VTAIL.n75 VSUBS 0.727571f
C295 VTAIL.n76 VSUBS 0.017686f
C296 VTAIL.t2 VSUBS 0.090073f
C297 VTAIL.n77 VSUBS 0.168078f
C298 VTAIL.n78 VSUBS 0.031434f
C299 VTAIL.n79 VSUBS 0.031353f
C300 VTAIL.n80 VSUBS 0.041804f
C301 VTAIL.n81 VSUBS 0.018726f
C302 VTAIL.n82 VSUBS 0.017686f
C303 VTAIL.n83 VSUBS 0.032913f
C304 VTAIL.n84 VSUBS 0.032913f
C305 VTAIL.n85 VSUBS 0.017686f
C306 VTAIL.n86 VSUBS 0.018726f
C307 VTAIL.n87 VSUBS 0.041804f
C308 VTAIL.n88 VSUBS 0.041804f
C309 VTAIL.n89 VSUBS 0.018726f
C310 VTAIL.n90 VSUBS 0.017686f
C311 VTAIL.n91 VSUBS 0.032913f
C312 VTAIL.n92 VSUBS 0.08507f
C313 VTAIL.n93 VSUBS 0.017686f
C314 VTAIL.n94 VSUBS 0.018726f
C315 VTAIL.n95 VSUBS 0.093129f
C316 VTAIL.n96 VSUBS 0.062466f
C317 VTAIL.n97 VSUBS 1.47895f
C318 VTAIL.n98 VSUBS 0.018556f
C319 VTAIL.n99 VSUBS 0.041804f
C320 VTAIL.n100 VSUBS 0.018726f
C321 VTAIL.n101 VSUBS 0.032913f
C322 VTAIL.n102 VSUBS 0.017686f
C323 VTAIL.n103 VSUBS 0.041804f
C324 VTAIL.n104 VSUBS 0.018726f
C325 VTAIL.n105 VSUBS 0.727571f
C326 VTAIL.n106 VSUBS 0.017686f
C327 VTAIL.t5 VSUBS 0.090073f
C328 VTAIL.n107 VSUBS 0.168078f
C329 VTAIL.n108 VSUBS 0.031434f
C330 VTAIL.n109 VSUBS 0.031353f
C331 VTAIL.n110 VSUBS 0.041804f
C332 VTAIL.n111 VSUBS 0.018726f
C333 VTAIL.n112 VSUBS 0.017686f
C334 VTAIL.n113 VSUBS 0.032913f
C335 VTAIL.n114 VSUBS 0.032913f
C336 VTAIL.n115 VSUBS 0.017686f
C337 VTAIL.n116 VSUBS 0.018726f
C338 VTAIL.n117 VSUBS 0.041804f
C339 VTAIL.n118 VSUBS 0.041804f
C340 VTAIL.n119 VSUBS 0.018726f
C341 VTAIL.n120 VSUBS 0.017686f
C342 VTAIL.n121 VSUBS 0.032913f
C343 VTAIL.n122 VSUBS 0.08507f
C344 VTAIL.n123 VSUBS 0.017686f
C345 VTAIL.n124 VSUBS 0.018726f
C346 VTAIL.n125 VSUBS 0.093129f
C347 VTAIL.n126 VSUBS 0.062466f
C348 VTAIL.n127 VSUBS 1.4145f
C349 VN.n0 VSUBS 0.054044f
C350 VN.t1 VSUBS 1.40446f
C351 VN.n1 VSUBS 0.033438f
C352 VN.n2 VSUBS 0.349812f
C353 VN.t4 VSUBS 1.40446f
C354 VN.t2 VSUBS 1.6618f
C355 VN.n3 VSUBS 0.624233f
C356 VN.n4 VSUBS 0.639722f
C357 VN.n5 VSUBS 0.057256f
C358 VN.n6 VSUBS 0.081891f
C359 VN.n7 VSUBS 0.040995f
C360 VN.n8 VSUBS 0.040995f
C361 VN.n9 VSUBS 0.040995f
C362 VN.n10 VSUBS 0.079877f
C363 VN.n11 VSUBS 0.061009f
C364 VN.n12 VSUBS 0.659977f
C365 VN.n13 VSUBS 0.057342f
C366 VN.n14 VSUBS 0.054044f
C367 VN.t0 VSUBS 1.40446f
C368 VN.n15 VSUBS 0.033438f
C369 VN.n16 VSUBS 0.349812f
C370 VN.t5 VSUBS 1.40446f
C371 VN.t3 VSUBS 1.6618f
C372 VN.n17 VSUBS 0.624233f
C373 VN.n18 VSUBS 0.639722f
C374 VN.n19 VSUBS 0.057256f
C375 VN.n20 VSUBS 0.081891f
C376 VN.n21 VSUBS 0.040995f
C377 VN.n22 VSUBS 0.040995f
C378 VN.n23 VSUBS 0.040995f
C379 VN.n24 VSUBS 0.079877f
C380 VN.n25 VSUBS 0.061009f
C381 VN.n26 VSUBS 0.659977f
C382 VN.n27 VSUBS 1.79149f
C383 B.n0 VSUBS 0.004977f
C384 B.n1 VSUBS 0.004977f
C385 B.n2 VSUBS 0.007871f
C386 B.n3 VSUBS 0.007871f
C387 B.n4 VSUBS 0.007871f
C388 B.n5 VSUBS 0.007871f
C389 B.n6 VSUBS 0.007871f
C390 B.n7 VSUBS 0.007871f
C391 B.n8 VSUBS 0.007871f
C392 B.n9 VSUBS 0.007871f
C393 B.n10 VSUBS 0.007871f
C394 B.n11 VSUBS 0.007871f
C395 B.n12 VSUBS 0.007871f
C396 B.n13 VSUBS 0.007871f
C397 B.n14 VSUBS 0.007871f
C398 B.n15 VSUBS 0.007871f
C399 B.n16 VSUBS 0.007871f
C400 B.n17 VSUBS 0.007871f
C401 B.n18 VSUBS 0.007871f
C402 B.n19 VSUBS 0.007871f
C403 B.n20 VSUBS 0.007871f
C404 B.n21 VSUBS 0.018661f
C405 B.n22 VSUBS 0.007871f
C406 B.n23 VSUBS 0.007871f
C407 B.n24 VSUBS 0.007871f
C408 B.n25 VSUBS 0.007871f
C409 B.n26 VSUBS 0.007871f
C410 B.n27 VSUBS 0.007871f
C411 B.n28 VSUBS 0.007871f
C412 B.n29 VSUBS 0.007871f
C413 B.n30 VSUBS 0.007871f
C414 B.n31 VSUBS 0.007871f
C415 B.n32 VSUBS 0.007871f
C416 B.n33 VSUBS 0.007871f
C417 B.t11 VSUBS 0.097144f
C418 B.t10 VSUBS 0.122281f
C419 B.t9 VSUBS 0.684859f
C420 B.n34 VSUBS 0.211809f
C421 B.n35 VSUBS 0.171106f
C422 B.n36 VSUBS 0.007871f
C423 B.n37 VSUBS 0.007871f
C424 B.n38 VSUBS 0.007871f
C425 B.n39 VSUBS 0.007871f
C426 B.t5 VSUBS 0.097146f
C427 B.t4 VSUBS 0.122283f
C428 B.t3 VSUBS 0.684859f
C429 B.n40 VSUBS 0.211808f
C430 B.n41 VSUBS 0.171104f
C431 B.n42 VSUBS 0.007871f
C432 B.n43 VSUBS 0.007871f
C433 B.n44 VSUBS 0.007871f
C434 B.n45 VSUBS 0.007871f
C435 B.n46 VSUBS 0.007871f
C436 B.n47 VSUBS 0.007871f
C437 B.n48 VSUBS 0.007871f
C438 B.n49 VSUBS 0.007871f
C439 B.n50 VSUBS 0.007871f
C440 B.n51 VSUBS 0.007871f
C441 B.n52 VSUBS 0.007871f
C442 B.n53 VSUBS 0.018661f
C443 B.n54 VSUBS 0.007871f
C444 B.n55 VSUBS 0.007871f
C445 B.n56 VSUBS 0.007871f
C446 B.n57 VSUBS 0.007871f
C447 B.n58 VSUBS 0.007871f
C448 B.n59 VSUBS 0.007871f
C449 B.n60 VSUBS 0.007871f
C450 B.n61 VSUBS 0.007871f
C451 B.n62 VSUBS 0.007871f
C452 B.n63 VSUBS 0.007871f
C453 B.n64 VSUBS 0.007871f
C454 B.n65 VSUBS 0.007871f
C455 B.n66 VSUBS 0.007871f
C456 B.n67 VSUBS 0.007871f
C457 B.n68 VSUBS 0.007871f
C458 B.n69 VSUBS 0.007871f
C459 B.n70 VSUBS 0.007871f
C460 B.n71 VSUBS 0.007871f
C461 B.n72 VSUBS 0.007871f
C462 B.n73 VSUBS 0.007871f
C463 B.n74 VSUBS 0.007871f
C464 B.n75 VSUBS 0.007871f
C465 B.n76 VSUBS 0.007871f
C466 B.n77 VSUBS 0.007871f
C467 B.n78 VSUBS 0.007871f
C468 B.n79 VSUBS 0.007871f
C469 B.n80 VSUBS 0.007871f
C470 B.n81 VSUBS 0.007871f
C471 B.n82 VSUBS 0.007871f
C472 B.n83 VSUBS 0.007871f
C473 B.n84 VSUBS 0.007871f
C474 B.n85 VSUBS 0.007871f
C475 B.n86 VSUBS 0.007871f
C476 B.n87 VSUBS 0.007871f
C477 B.n88 VSUBS 0.007871f
C478 B.n89 VSUBS 0.007871f
C479 B.n90 VSUBS 0.007871f
C480 B.n91 VSUBS 0.007871f
C481 B.n92 VSUBS 0.018661f
C482 B.n93 VSUBS 0.007871f
C483 B.n94 VSUBS 0.007871f
C484 B.n95 VSUBS 0.007871f
C485 B.n96 VSUBS 0.007871f
C486 B.n97 VSUBS 0.007871f
C487 B.n98 VSUBS 0.007871f
C488 B.n99 VSUBS 0.007871f
C489 B.n100 VSUBS 0.007871f
C490 B.n101 VSUBS 0.007871f
C491 B.n102 VSUBS 0.007871f
C492 B.n103 VSUBS 0.007871f
C493 B.t7 VSUBS 0.097146f
C494 B.t8 VSUBS 0.122283f
C495 B.t6 VSUBS 0.684859f
C496 B.n104 VSUBS 0.211808f
C497 B.n105 VSUBS 0.171104f
C498 B.n106 VSUBS 0.018236f
C499 B.n107 VSUBS 0.007871f
C500 B.n108 VSUBS 0.007871f
C501 B.n109 VSUBS 0.007871f
C502 B.n110 VSUBS 0.007871f
C503 B.n111 VSUBS 0.007871f
C504 B.t1 VSUBS 0.097144f
C505 B.t2 VSUBS 0.122281f
C506 B.t0 VSUBS 0.684859f
C507 B.n112 VSUBS 0.211809f
C508 B.n113 VSUBS 0.171106f
C509 B.n114 VSUBS 0.007871f
C510 B.n115 VSUBS 0.007871f
C511 B.n116 VSUBS 0.007871f
C512 B.n117 VSUBS 0.007871f
C513 B.n118 VSUBS 0.007871f
C514 B.n119 VSUBS 0.007871f
C515 B.n120 VSUBS 0.007871f
C516 B.n121 VSUBS 0.007871f
C517 B.n122 VSUBS 0.007871f
C518 B.n123 VSUBS 0.007871f
C519 B.n124 VSUBS 0.007871f
C520 B.n125 VSUBS 0.017221f
C521 B.n126 VSUBS 0.007871f
C522 B.n127 VSUBS 0.007871f
C523 B.n128 VSUBS 0.007871f
C524 B.n129 VSUBS 0.007871f
C525 B.n130 VSUBS 0.007871f
C526 B.n131 VSUBS 0.007871f
C527 B.n132 VSUBS 0.007871f
C528 B.n133 VSUBS 0.007871f
C529 B.n134 VSUBS 0.007871f
C530 B.n135 VSUBS 0.007871f
C531 B.n136 VSUBS 0.007871f
C532 B.n137 VSUBS 0.007871f
C533 B.n138 VSUBS 0.007871f
C534 B.n139 VSUBS 0.007871f
C535 B.n140 VSUBS 0.007871f
C536 B.n141 VSUBS 0.007871f
C537 B.n142 VSUBS 0.007871f
C538 B.n143 VSUBS 0.007871f
C539 B.n144 VSUBS 0.007871f
C540 B.n145 VSUBS 0.007871f
C541 B.n146 VSUBS 0.007871f
C542 B.n147 VSUBS 0.007871f
C543 B.n148 VSUBS 0.007871f
C544 B.n149 VSUBS 0.007871f
C545 B.n150 VSUBS 0.007871f
C546 B.n151 VSUBS 0.007871f
C547 B.n152 VSUBS 0.007871f
C548 B.n153 VSUBS 0.007871f
C549 B.n154 VSUBS 0.007871f
C550 B.n155 VSUBS 0.007871f
C551 B.n156 VSUBS 0.007871f
C552 B.n157 VSUBS 0.007871f
C553 B.n158 VSUBS 0.007871f
C554 B.n159 VSUBS 0.007871f
C555 B.n160 VSUBS 0.007871f
C556 B.n161 VSUBS 0.007871f
C557 B.n162 VSUBS 0.007871f
C558 B.n163 VSUBS 0.007871f
C559 B.n164 VSUBS 0.007871f
C560 B.n165 VSUBS 0.007871f
C561 B.n166 VSUBS 0.007871f
C562 B.n167 VSUBS 0.007871f
C563 B.n168 VSUBS 0.007871f
C564 B.n169 VSUBS 0.007871f
C565 B.n170 VSUBS 0.007871f
C566 B.n171 VSUBS 0.007871f
C567 B.n172 VSUBS 0.007871f
C568 B.n173 VSUBS 0.007871f
C569 B.n174 VSUBS 0.007871f
C570 B.n175 VSUBS 0.007871f
C571 B.n176 VSUBS 0.007871f
C572 B.n177 VSUBS 0.007871f
C573 B.n178 VSUBS 0.007871f
C574 B.n179 VSUBS 0.007871f
C575 B.n180 VSUBS 0.007871f
C576 B.n181 VSUBS 0.007871f
C577 B.n182 VSUBS 0.007871f
C578 B.n183 VSUBS 0.007871f
C579 B.n184 VSUBS 0.007871f
C580 B.n185 VSUBS 0.007871f
C581 B.n186 VSUBS 0.007871f
C582 B.n187 VSUBS 0.007871f
C583 B.n188 VSUBS 0.007871f
C584 B.n189 VSUBS 0.007871f
C585 B.n190 VSUBS 0.007871f
C586 B.n191 VSUBS 0.007871f
C587 B.n192 VSUBS 0.007871f
C588 B.n193 VSUBS 0.007871f
C589 B.n194 VSUBS 0.007871f
C590 B.n195 VSUBS 0.007871f
C591 B.n196 VSUBS 0.007871f
C592 B.n197 VSUBS 0.007871f
C593 B.n198 VSUBS 0.017221f
C594 B.n199 VSUBS 0.018661f
C595 B.n200 VSUBS 0.018661f
C596 B.n201 VSUBS 0.007871f
C597 B.n202 VSUBS 0.007871f
C598 B.n203 VSUBS 0.007871f
C599 B.n204 VSUBS 0.007871f
C600 B.n205 VSUBS 0.007871f
C601 B.n206 VSUBS 0.007871f
C602 B.n207 VSUBS 0.007871f
C603 B.n208 VSUBS 0.007871f
C604 B.n209 VSUBS 0.007871f
C605 B.n210 VSUBS 0.007871f
C606 B.n211 VSUBS 0.007871f
C607 B.n212 VSUBS 0.007871f
C608 B.n213 VSUBS 0.007871f
C609 B.n214 VSUBS 0.007871f
C610 B.n215 VSUBS 0.007871f
C611 B.n216 VSUBS 0.007871f
C612 B.n217 VSUBS 0.007871f
C613 B.n218 VSUBS 0.007871f
C614 B.n219 VSUBS 0.007871f
C615 B.n220 VSUBS 0.007871f
C616 B.n221 VSUBS 0.007871f
C617 B.n222 VSUBS 0.007871f
C618 B.n223 VSUBS 0.007871f
C619 B.n224 VSUBS 0.007871f
C620 B.n225 VSUBS 0.007871f
C621 B.n226 VSUBS 0.007871f
C622 B.n227 VSUBS 0.007871f
C623 B.n228 VSUBS 0.007871f
C624 B.n229 VSUBS 0.007871f
C625 B.n230 VSUBS 0.007871f
C626 B.n231 VSUBS 0.007871f
C627 B.n232 VSUBS 0.007871f
C628 B.n233 VSUBS 0.007871f
C629 B.n234 VSUBS 0.00544f
C630 B.n235 VSUBS 0.018236f
C631 B.n236 VSUBS 0.006366f
C632 B.n237 VSUBS 0.007871f
C633 B.n238 VSUBS 0.007871f
C634 B.n239 VSUBS 0.007871f
C635 B.n240 VSUBS 0.007871f
C636 B.n241 VSUBS 0.007871f
C637 B.n242 VSUBS 0.007871f
C638 B.n243 VSUBS 0.007871f
C639 B.n244 VSUBS 0.007871f
C640 B.n245 VSUBS 0.007871f
C641 B.n246 VSUBS 0.007871f
C642 B.n247 VSUBS 0.007871f
C643 B.n248 VSUBS 0.006366f
C644 B.n249 VSUBS 0.007871f
C645 B.n250 VSUBS 0.007871f
C646 B.n251 VSUBS 0.00544f
C647 B.n252 VSUBS 0.007871f
C648 B.n253 VSUBS 0.007871f
C649 B.n254 VSUBS 0.007871f
C650 B.n255 VSUBS 0.007871f
C651 B.n256 VSUBS 0.007871f
C652 B.n257 VSUBS 0.007871f
C653 B.n258 VSUBS 0.007871f
C654 B.n259 VSUBS 0.007871f
C655 B.n260 VSUBS 0.007871f
C656 B.n261 VSUBS 0.007871f
C657 B.n262 VSUBS 0.007871f
C658 B.n263 VSUBS 0.007871f
C659 B.n264 VSUBS 0.007871f
C660 B.n265 VSUBS 0.007871f
C661 B.n266 VSUBS 0.007871f
C662 B.n267 VSUBS 0.007871f
C663 B.n268 VSUBS 0.007871f
C664 B.n269 VSUBS 0.007871f
C665 B.n270 VSUBS 0.007871f
C666 B.n271 VSUBS 0.007871f
C667 B.n272 VSUBS 0.007871f
C668 B.n273 VSUBS 0.007871f
C669 B.n274 VSUBS 0.007871f
C670 B.n275 VSUBS 0.007871f
C671 B.n276 VSUBS 0.007871f
C672 B.n277 VSUBS 0.007871f
C673 B.n278 VSUBS 0.007871f
C674 B.n279 VSUBS 0.007871f
C675 B.n280 VSUBS 0.007871f
C676 B.n281 VSUBS 0.007871f
C677 B.n282 VSUBS 0.007871f
C678 B.n283 VSUBS 0.007871f
C679 B.n284 VSUBS 0.007871f
C680 B.n285 VSUBS 0.018661f
C681 B.n286 VSUBS 0.017221f
C682 B.n287 VSUBS 0.017221f
C683 B.n288 VSUBS 0.007871f
C684 B.n289 VSUBS 0.007871f
C685 B.n290 VSUBS 0.007871f
C686 B.n291 VSUBS 0.007871f
C687 B.n292 VSUBS 0.007871f
C688 B.n293 VSUBS 0.007871f
C689 B.n294 VSUBS 0.007871f
C690 B.n295 VSUBS 0.007871f
C691 B.n296 VSUBS 0.007871f
C692 B.n297 VSUBS 0.007871f
C693 B.n298 VSUBS 0.007871f
C694 B.n299 VSUBS 0.007871f
C695 B.n300 VSUBS 0.007871f
C696 B.n301 VSUBS 0.007871f
C697 B.n302 VSUBS 0.007871f
C698 B.n303 VSUBS 0.007871f
C699 B.n304 VSUBS 0.007871f
C700 B.n305 VSUBS 0.007871f
C701 B.n306 VSUBS 0.007871f
C702 B.n307 VSUBS 0.007871f
C703 B.n308 VSUBS 0.007871f
C704 B.n309 VSUBS 0.007871f
C705 B.n310 VSUBS 0.007871f
C706 B.n311 VSUBS 0.007871f
C707 B.n312 VSUBS 0.007871f
C708 B.n313 VSUBS 0.007871f
C709 B.n314 VSUBS 0.007871f
C710 B.n315 VSUBS 0.007871f
C711 B.n316 VSUBS 0.007871f
C712 B.n317 VSUBS 0.007871f
C713 B.n318 VSUBS 0.007871f
C714 B.n319 VSUBS 0.007871f
C715 B.n320 VSUBS 0.007871f
C716 B.n321 VSUBS 0.007871f
C717 B.n322 VSUBS 0.007871f
C718 B.n323 VSUBS 0.007871f
C719 B.n324 VSUBS 0.007871f
C720 B.n325 VSUBS 0.007871f
C721 B.n326 VSUBS 0.007871f
C722 B.n327 VSUBS 0.007871f
C723 B.n328 VSUBS 0.007871f
C724 B.n329 VSUBS 0.007871f
C725 B.n330 VSUBS 0.007871f
C726 B.n331 VSUBS 0.007871f
C727 B.n332 VSUBS 0.007871f
C728 B.n333 VSUBS 0.007871f
C729 B.n334 VSUBS 0.007871f
C730 B.n335 VSUBS 0.007871f
C731 B.n336 VSUBS 0.007871f
C732 B.n337 VSUBS 0.007871f
C733 B.n338 VSUBS 0.007871f
C734 B.n339 VSUBS 0.007871f
C735 B.n340 VSUBS 0.007871f
C736 B.n341 VSUBS 0.007871f
C737 B.n342 VSUBS 0.007871f
C738 B.n343 VSUBS 0.007871f
C739 B.n344 VSUBS 0.007871f
C740 B.n345 VSUBS 0.007871f
C741 B.n346 VSUBS 0.007871f
C742 B.n347 VSUBS 0.007871f
C743 B.n348 VSUBS 0.007871f
C744 B.n349 VSUBS 0.007871f
C745 B.n350 VSUBS 0.007871f
C746 B.n351 VSUBS 0.007871f
C747 B.n352 VSUBS 0.007871f
C748 B.n353 VSUBS 0.007871f
C749 B.n354 VSUBS 0.007871f
C750 B.n355 VSUBS 0.007871f
C751 B.n356 VSUBS 0.007871f
C752 B.n357 VSUBS 0.007871f
C753 B.n358 VSUBS 0.007871f
C754 B.n359 VSUBS 0.007871f
C755 B.n360 VSUBS 0.007871f
C756 B.n361 VSUBS 0.007871f
C757 B.n362 VSUBS 0.007871f
C758 B.n363 VSUBS 0.007871f
C759 B.n364 VSUBS 0.007871f
C760 B.n365 VSUBS 0.007871f
C761 B.n366 VSUBS 0.007871f
C762 B.n367 VSUBS 0.007871f
C763 B.n368 VSUBS 0.007871f
C764 B.n369 VSUBS 0.007871f
C765 B.n370 VSUBS 0.007871f
C766 B.n371 VSUBS 0.007871f
C767 B.n372 VSUBS 0.007871f
C768 B.n373 VSUBS 0.007871f
C769 B.n374 VSUBS 0.007871f
C770 B.n375 VSUBS 0.007871f
C771 B.n376 VSUBS 0.007871f
C772 B.n377 VSUBS 0.007871f
C773 B.n378 VSUBS 0.007871f
C774 B.n379 VSUBS 0.007871f
C775 B.n380 VSUBS 0.007871f
C776 B.n381 VSUBS 0.007871f
C777 B.n382 VSUBS 0.007871f
C778 B.n383 VSUBS 0.007871f
C779 B.n384 VSUBS 0.007871f
C780 B.n385 VSUBS 0.007871f
C781 B.n386 VSUBS 0.007871f
C782 B.n387 VSUBS 0.007871f
C783 B.n388 VSUBS 0.007871f
C784 B.n389 VSUBS 0.007871f
C785 B.n390 VSUBS 0.007871f
C786 B.n391 VSUBS 0.007871f
C787 B.n392 VSUBS 0.007871f
C788 B.n393 VSUBS 0.007871f
C789 B.n394 VSUBS 0.007871f
C790 B.n395 VSUBS 0.007871f
C791 B.n396 VSUBS 0.007871f
C792 B.n397 VSUBS 0.007871f
C793 B.n398 VSUBS 0.007871f
C794 B.n399 VSUBS 0.007871f
C795 B.n400 VSUBS 0.017221f
C796 B.n401 VSUBS 0.018189f
C797 B.n402 VSUBS 0.017693f
C798 B.n403 VSUBS 0.007871f
C799 B.n404 VSUBS 0.007871f
C800 B.n405 VSUBS 0.007871f
C801 B.n406 VSUBS 0.007871f
C802 B.n407 VSUBS 0.007871f
C803 B.n408 VSUBS 0.007871f
C804 B.n409 VSUBS 0.007871f
C805 B.n410 VSUBS 0.007871f
C806 B.n411 VSUBS 0.007871f
C807 B.n412 VSUBS 0.007871f
C808 B.n413 VSUBS 0.007871f
C809 B.n414 VSUBS 0.007871f
C810 B.n415 VSUBS 0.007871f
C811 B.n416 VSUBS 0.007871f
C812 B.n417 VSUBS 0.007871f
C813 B.n418 VSUBS 0.007871f
C814 B.n419 VSUBS 0.007871f
C815 B.n420 VSUBS 0.007871f
C816 B.n421 VSUBS 0.007871f
C817 B.n422 VSUBS 0.007871f
C818 B.n423 VSUBS 0.007871f
C819 B.n424 VSUBS 0.007871f
C820 B.n425 VSUBS 0.007871f
C821 B.n426 VSUBS 0.007871f
C822 B.n427 VSUBS 0.007871f
C823 B.n428 VSUBS 0.007871f
C824 B.n429 VSUBS 0.007871f
C825 B.n430 VSUBS 0.007871f
C826 B.n431 VSUBS 0.007871f
C827 B.n432 VSUBS 0.007871f
C828 B.n433 VSUBS 0.007871f
C829 B.n434 VSUBS 0.007871f
C830 B.n435 VSUBS 0.007871f
C831 B.n436 VSUBS 0.007871f
C832 B.n437 VSUBS 0.00544f
C833 B.n438 VSUBS 0.018236f
C834 B.n439 VSUBS 0.006366f
C835 B.n440 VSUBS 0.007871f
C836 B.n441 VSUBS 0.007871f
C837 B.n442 VSUBS 0.007871f
C838 B.n443 VSUBS 0.007871f
C839 B.n444 VSUBS 0.007871f
C840 B.n445 VSUBS 0.007871f
C841 B.n446 VSUBS 0.007871f
C842 B.n447 VSUBS 0.007871f
C843 B.n448 VSUBS 0.007871f
C844 B.n449 VSUBS 0.007871f
C845 B.n450 VSUBS 0.007871f
C846 B.n451 VSUBS 0.006366f
C847 B.n452 VSUBS 0.018236f
C848 B.n453 VSUBS 0.00544f
C849 B.n454 VSUBS 0.007871f
C850 B.n455 VSUBS 0.007871f
C851 B.n456 VSUBS 0.007871f
C852 B.n457 VSUBS 0.007871f
C853 B.n458 VSUBS 0.007871f
C854 B.n459 VSUBS 0.007871f
C855 B.n460 VSUBS 0.007871f
C856 B.n461 VSUBS 0.007871f
C857 B.n462 VSUBS 0.007871f
C858 B.n463 VSUBS 0.007871f
C859 B.n464 VSUBS 0.007871f
C860 B.n465 VSUBS 0.007871f
C861 B.n466 VSUBS 0.007871f
C862 B.n467 VSUBS 0.007871f
C863 B.n468 VSUBS 0.007871f
C864 B.n469 VSUBS 0.007871f
C865 B.n470 VSUBS 0.007871f
C866 B.n471 VSUBS 0.007871f
C867 B.n472 VSUBS 0.007871f
C868 B.n473 VSUBS 0.007871f
C869 B.n474 VSUBS 0.007871f
C870 B.n475 VSUBS 0.007871f
C871 B.n476 VSUBS 0.007871f
C872 B.n477 VSUBS 0.007871f
C873 B.n478 VSUBS 0.007871f
C874 B.n479 VSUBS 0.007871f
C875 B.n480 VSUBS 0.007871f
C876 B.n481 VSUBS 0.007871f
C877 B.n482 VSUBS 0.007871f
C878 B.n483 VSUBS 0.007871f
C879 B.n484 VSUBS 0.007871f
C880 B.n485 VSUBS 0.007871f
C881 B.n486 VSUBS 0.007871f
C882 B.n487 VSUBS 0.007871f
C883 B.n488 VSUBS 0.018661f
C884 B.n489 VSUBS 0.017221f
C885 B.n490 VSUBS 0.017221f
C886 B.n491 VSUBS 0.007871f
C887 B.n492 VSUBS 0.007871f
C888 B.n493 VSUBS 0.007871f
C889 B.n494 VSUBS 0.007871f
C890 B.n495 VSUBS 0.007871f
C891 B.n496 VSUBS 0.007871f
C892 B.n497 VSUBS 0.007871f
C893 B.n498 VSUBS 0.007871f
C894 B.n499 VSUBS 0.007871f
C895 B.n500 VSUBS 0.007871f
C896 B.n501 VSUBS 0.007871f
C897 B.n502 VSUBS 0.007871f
C898 B.n503 VSUBS 0.007871f
C899 B.n504 VSUBS 0.007871f
C900 B.n505 VSUBS 0.007871f
C901 B.n506 VSUBS 0.007871f
C902 B.n507 VSUBS 0.007871f
C903 B.n508 VSUBS 0.007871f
C904 B.n509 VSUBS 0.007871f
C905 B.n510 VSUBS 0.007871f
C906 B.n511 VSUBS 0.007871f
C907 B.n512 VSUBS 0.007871f
C908 B.n513 VSUBS 0.007871f
C909 B.n514 VSUBS 0.007871f
C910 B.n515 VSUBS 0.007871f
C911 B.n516 VSUBS 0.007871f
C912 B.n517 VSUBS 0.007871f
C913 B.n518 VSUBS 0.007871f
C914 B.n519 VSUBS 0.007871f
C915 B.n520 VSUBS 0.007871f
C916 B.n521 VSUBS 0.007871f
C917 B.n522 VSUBS 0.007871f
C918 B.n523 VSUBS 0.007871f
C919 B.n524 VSUBS 0.007871f
C920 B.n525 VSUBS 0.007871f
C921 B.n526 VSUBS 0.007871f
C922 B.n527 VSUBS 0.007871f
C923 B.n528 VSUBS 0.007871f
C924 B.n529 VSUBS 0.007871f
C925 B.n530 VSUBS 0.007871f
C926 B.n531 VSUBS 0.007871f
C927 B.n532 VSUBS 0.007871f
C928 B.n533 VSUBS 0.007871f
C929 B.n534 VSUBS 0.007871f
C930 B.n535 VSUBS 0.007871f
C931 B.n536 VSUBS 0.007871f
C932 B.n537 VSUBS 0.007871f
C933 B.n538 VSUBS 0.007871f
C934 B.n539 VSUBS 0.007871f
C935 B.n540 VSUBS 0.007871f
C936 B.n541 VSUBS 0.007871f
C937 B.n542 VSUBS 0.007871f
C938 B.n543 VSUBS 0.007871f
C939 B.n544 VSUBS 0.007871f
C940 B.n545 VSUBS 0.007871f
C941 B.n546 VSUBS 0.007871f
C942 B.n547 VSUBS 0.017822f
.ends

