* NGSPICE file created from diff_pair_sample_0490.ext - technology: sky130A

.subckt diff_pair_sample_0490 VTAIL VN VP B VDD2 VDD1
X0 B.t21 B.t19 B.t20 B.t13 sky130_fd_pr__nfet_01v8 ad=3.0147 pd=16.24 as=0 ps=0 w=7.73 l=0.57
X1 VTAIL.t15 VP.t0 VDD1.t0 B.t6 sky130_fd_pr__nfet_01v8 ad=3.0147 pd=16.24 as=1.27545 ps=8.06 w=7.73 l=0.57
X2 VDD1.t1 VP.t1 VTAIL.t14 B.t4 sky130_fd_pr__nfet_01v8 ad=1.27545 pd=8.06 as=1.27545 ps=8.06 w=7.73 l=0.57
X3 B.t18 B.t16 B.t17 B.t9 sky130_fd_pr__nfet_01v8 ad=3.0147 pd=16.24 as=0 ps=0 w=7.73 l=0.57
X4 VTAIL.t3 VN.t0 VDD2.t7 B.t6 sky130_fd_pr__nfet_01v8 ad=3.0147 pd=16.24 as=1.27545 ps=8.06 w=7.73 l=0.57
X5 VDD1.t2 VP.t2 VTAIL.t13 B.t7 sky130_fd_pr__nfet_01v8 ad=1.27545 pd=8.06 as=3.0147 ps=16.24 w=7.73 l=0.57
X6 VTAIL.t1 VN.t1 VDD2.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=3.0147 pd=16.24 as=1.27545 ps=8.06 w=7.73 l=0.57
X7 VDD2.t5 VN.t2 VTAIL.t2 B.t4 sky130_fd_pr__nfet_01v8 ad=1.27545 pd=8.06 as=1.27545 ps=8.06 w=7.73 l=0.57
X8 VDD1.t3 VP.t3 VTAIL.t12 B.t0 sky130_fd_pr__nfet_01v8 ad=1.27545 pd=8.06 as=3.0147 ps=16.24 w=7.73 l=0.57
X9 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=3.0147 pd=16.24 as=0 ps=0 w=7.73 l=0.57
X10 VTAIL.t11 VP.t4 VDD1.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=1.27545 pd=8.06 as=1.27545 ps=8.06 w=7.73 l=0.57
X11 VDD2.t4 VN.t3 VTAIL.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=1.27545 pd=8.06 as=1.27545 ps=8.06 w=7.73 l=0.57
X12 VTAIL.t6 VN.t4 VDD2.t3 B.t5 sky130_fd_pr__nfet_01v8 ad=1.27545 pd=8.06 as=1.27545 ps=8.06 w=7.73 l=0.57
X13 VDD1.t5 VP.t5 VTAIL.t10 B.t1 sky130_fd_pr__nfet_01v8 ad=1.27545 pd=8.06 as=1.27545 ps=8.06 w=7.73 l=0.57
X14 VDD2.t2 VN.t5 VTAIL.t5 B.t0 sky130_fd_pr__nfet_01v8 ad=1.27545 pd=8.06 as=3.0147 ps=16.24 w=7.73 l=0.57
X15 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=3.0147 pd=16.24 as=0 ps=0 w=7.73 l=0.57
X16 VTAIL.t9 VP.t6 VDD1.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=3.0147 pd=16.24 as=1.27545 ps=8.06 w=7.73 l=0.57
X17 VTAIL.t8 VP.t7 VDD1.t7 B.t5 sky130_fd_pr__nfet_01v8 ad=1.27545 pd=8.06 as=1.27545 ps=8.06 w=7.73 l=0.57
X18 VDD2.t1 VN.t6 VTAIL.t4 B.t7 sky130_fd_pr__nfet_01v8 ad=1.27545 pd=8.06 as=3.0147 ps=16.24 w=7.73 l=0.57
X19 VTAIL.t7 VN.t7 VDD2.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=1.27545 pd=8.06 as=1.27545 ps=8.06 w=7.73 l=0.57
R0 B.n524 B.n523 585
R1 B.n215 B.n76 585
R2 B.n214 B.n213 585
R3 B.n212 B.n211 585
R4 B.n210 B.n209 585
R5 B.n208 B.n207 585
R6 B.n206 B.n205 585
R7 B.n204 B.n203 585
R8 B.n202 B.n201 585
R9 B.n200 B.n199 585
R10 B.n198 B.n197 585
R11 B.n196 B.n195 585
R12 B.n194 B.n193 585
R13 B.n192 B.n191 585
R14 B.n190 B.n189 585
R15 B.n188 B.n187 585
R16 B.n186 B.n185 585
R17 B.n184 B.n183 585
R18 B.n182 B.n181 585
R19 B.n180 B.n179 585
R20 B.n178 B.n177 585
R21 B.n176 B.n175 585
R22 B.n174 B.n173 585
R23 B.n172 B.n171 585
R24 B.n170 B.n169 585
R25 B.n168 B.n167 585
R26 B.n166 B.n165 585
R27 B.n164 B.n163 585
R28 B.n162 B.n161 585
R29 B.n159 B.n158 585
R30 B.n157 B.n156 585
R31 B.n155 B.n154 585
R32 B.n153 B.n152 585
R33 B.n151 B.n150 585
R34 B.n149 B.n148 585
R35 B.n147 B.n146 585
R36 B.n145 B.n144 585
R37 B.n143 B.n142 585
R38 B.n141 B.n140 585
R39 B.n138 B.n137 585
R40 B.n136 B.n135 585
R41 B.n134 B.n133 585
R42 B.n132 B.n131 585
R43 B.n130 B.n129 585
R44 B.n128 B.n127 585
R45 B.n126 B.n125 585
R46 B.n124 B.n123 585
R47 B.n122 B.n121 585
R48 B.n120 B.n119 585
R49 B.n118 B.n117 585
R50 B.n116 B.n115 585
R51 B.n114 B.n113 585
R52 B.n112 B.n111 585
R53 B.n110 B.n109 585
R54 B.n108 B.n107 585
R55 B.n106 B.n105 585
R56 B.n104 B.n103 585
R57 B.n102 B.n101 585
R58 B.n100 B.n99 585
R59 B.n98 B.n97 585
R60 B.n96 B.n95 585
R61 B.n94 B.n93 585
R62 B.n92 B.n91 585
R63 B.n90 B.n89 585
R64 B.n88 B.n87 585
R65 B.n86 B.n85 585
R66 B.n84 B.n83 585
R67 B.n82 B.n81 585
R68 B.n522 B.n42 585
R69 B.n527 B.n42 585
R70 B.n521 B.n41 585
R71 B.n528 B.n41 585
R72 B.n520 B.n519 585
R73 B.n519 B.n37 585
R74 B.n518 B.n36 585
R75 B.n534 B.n36 585
R76 B.n517 B.n35 585
R77 B.n535 B.n35 585
R78 B.n516 B.n34 585
R79 B.n536 B.n34 585
R80 B.n515 B.n514 585
R81 B.n514 B.n30 585
R82 B.n513 B.n29 585
R83 B.n542 B.n29 585
R84 B.n512 B.n28 585
R85 B.n543 B.n28 585
R86 B.n511 B.n27 585
R87 B.n544 B.n27 585
R88 B.n510 B.n509 585
R89 B.n509 B.n26 585
R90 B.n508 B.n22 585
R91 B.n550 B.n22 585
R92 B.n507 B.n21 585
R93 B.n551 B.n21 585
R94 B.n506 B.n20 585
R95 B.n552 B.n20 585
R96 B.n505 B.n504 585
R97 B.n504 B.n16 585
R98 B.n503 B.n15 585
R99 B.n558 B.n15 585
R100 B.n502 B.n14 585
R101 B.n559 B.n14 585
R102 B.n501 B.n13 585
R103 B.n560 B.n13 585
R104 B.n500 B.n499 585
R105 B.n499 B.n12 585
R106 B.n498 B.n497 585
R107 B.n498 B.n8 585
R108 B.n496 B.n7 585
R109 B.n567 B.n7 585
R110 B.n495 B.n6 585
R111 B.n568 B.n6 585
R112 B.n494 B.n5 585
R113 B.n569 B.n5 585
R114 B.n493 B.n492 585
R115 B.n492 B.n4 585
R116 B.n491 B.n216 585
R117 B.n491 B.n490 585
R118 B.n480 B.n217 585
R119 B.n483 B.n217 585
R120 B.n482 B.n481 585
R121 B.n484 B.n482 585
R122 B.n479 B.n222 585
R123 B.n222 B.n221 585
R124 B.n478 B.n477 585
R125 B.n477 B.n476 585
R126 B.n224 B.n223 585
R127 B.n225 B.n224 585
R128 B.n469 B.n468 585
R129 B.n470 B.n469 585
R130 B.n467 B.n230 585
R131 B.n230 B.n229 585
R132 B.n466 B.n465 585
R133 B.n465 B.n464 585
R134 B.n232 B.n231 585
R135 B.n457 B.n232 585
R136 B.n456 B.n455 585
R137 B.n458 B.n456 585
R138 B.n454 B.n237 585
R139 B.n237 B.n236 585
R140 B.n453 B.n452 585
R141 B.n452 B.n451 585
R142 B.n239 B.n238 585
R143 B.n240 B.n239 585
R144 B.n444 B.n443 585
R145 B.n445 B.n444 585
R146 B.n442 B.n244 585
R147 B.n248 B.n244 585
R148 B.n441 B.n440 585
R149 B.n440 B.n439 585
R150 B.n246 B.n245 585
R151 B.n247 B.n246 585
R152 B.n432 B.n431 585
R153 B.n433 B.n432 585
R154 B.n430 B.n253 585
R155 B.n253 B.n252 585
R156 B.n425 B.n424 585
R157 B.n423 B.n289 585
R158 B.n422 B.n288 585
R159 B.n427 B.n288 585
R160 B.n421 B.n420 585
R161 B.n419 B.n418 585
R162 B.n417 B.n416 585
R163 B.n415 B.n414 585
R164 B.n413 B.n412 585
R165 B.n411 B.n410 585
R166 B.n409 B.n408 585
R167 B.n407 B.n406 585
R168 B.n405 B.n404 585
R169 B.n403 B.n402 585
R170 B.n401 B.n400 585
R171 B.n399 B.n398 585
R172 B.n397 B.n396 585
R173 B.n395 B.n394 585
R174 B.n393 B.n392 585
R175 B.n391 B.n390 585
R176 B.n389 B.n388 585
R177 B.n387 B.n386 585
R178 B.n385 B.n384 585
R179 B.n383 B.n382 585
R180 B.n381 B.n380 585
R181 B.n379 B.n378 585
R182 B.n377 B.n376 585
R183 B.n375 B.n374 585
R184 B.n373 B.n372 585
R185 B.n371 B.n370 585
R186 B.n369 B.n368 585
R187 B.n367 B.n366 585
R188 B.n365 B.n364 585
R189 B.n363 B.n362 585
R190 B.n361 B.n360 585
R191 B.n359 B.n358 585
R192 B.n357 B.n356 585
R193 B.n355 B.n354 585
R194 B.n353 B.n352 585
R195 B.n351 B.n350 585
R196 B.n349 B.n348 585
R197 B.n347 B.n346 585
R198 B.n345 B.n344 585
R199 B.n343 B.n342 585
R200 B.n341 B.n340 585
R201 B.n339 B.n338 585
R202 B.n337 B.n336 585
R203 B.n335 B.n334 585
R204 B.n333 B.n332 585
R205 B.n331 B.n330 585
R206 B.n329 B.n328 585
R207 B.n327 B.n326 585
R208 B.n325 B.n324 585
R209 B.n323 B.n322 585
R210 B.n321 B.n320 585
R211 B.n319 B.n318 585
R212 B.n317 B.n316 585
R213 B.n315 B.n314 585
R214 B.n313 B.n312 585
R215 B.n311 B.n310 585
R216 B.n309 B.n308 585
R217 B.n307 B.n306 585
R218 B.n305 B.n304 585
R219 B.n303 B.n302 585
R220 B.n301 B.n300 585
R221 B.n299 B.n298 585
R222 B.n297 B.n296 585
R223 B.n255 B.n254 585
R224 B.n429 B.n428 585
R225 B.n428 B.n427 585
R226 B.n251 B.n250 585
R227 B.n252 B.n251 585
R228 B.n435 B.n434 585
R229 B.n434 B.n433 585
R230 B.n436 B.n249 585
R231 B.n249 B.n247 585
R232 B.n438 B.n437 585
R233 B.n439 B.n438 585
R234 B.n243 B.n242 585
R235 B.n248 B.n243 585
R236 B.n447 B.n446 585
R237 B.n446 B.n445 585
R238 B.n448 B.n241 585
R239 B.n241 B.n240 585
R240 B.n450 B.n449 585
R241 B.n451 B.n450 585
R242 B.n235 B.n234 585
R243 B.n236 B.n235 585
R244 B.n460 B.n459 585
R245 B.n459 B.n458 585
R246 B.n461 B.n233 585
R247 B.n457 B.n233 585
R248 B.n463 B.n462 585
R249 B.n464 B.n463 585
R250 B.n228 B.n227 585
R251 B.n229 B.n228 585
R252 B.n472 B.n471 585
R253 B.n471 B.n470 585
R254 B.n473 B.n226 585
R255 B.n226 B.n225 585
R256 B.n475 B.n474 585
R257 B.n476 B.n475 585
R258 B.n220 B.n219 585
R259 B.n221 B.n220 585
R260 B.n486 B.n485 585
R261 B.n485 B.n484 585
R262 B.n487 B.n218 585
R263 B.n483 B.n218 585
R264 B.n489 B.n488 585
R265 B.n490 B.n489 585
R266 B.n3 B.n0 585
R267 B.n4 B.n3 585
R268 B.n566 B.n1 585
R269 B.n567 B.n566 585
R270 B.n565 B.n564 585
R271 B.n565 B.n8 585
R272 B.n563 B.n9 585
R273 B.n12 B.n9 585
R274 B.n562 B.n561 585
R275 B.n561 B.n560 585
R276 B.n11 B.n10 585
R277 B.n559 B.n11 585
R278 B.n557 B.n556 585
R279 B.n558 B.n557 585
R280 B.n555 B.n17 585
R281 B.n17 B.n16 585
R282 B.n554 B.n553 585
R283 B.n553 B.n552 585
R284 B.n19 B.n18 585
R285 B.n551 B.n19 585
R286 B.n549 B.n548 585
R287 B.n550 B.n549 585
R288 B.n547 B.n23 585
R289 B.n26 B.n23 585
R290 B.n546 B.n545 585
R291 B.n545 B.n544 585
R292 B.n25 B.n24 585
R293 B.n543 B.n25 585
R294 B.n541 B.n540 585
R295 B.n542 B.n541 585
R296 B.n539 B.n31 585
R297 B.n31 B.n30 585
R298 B.n538 B.n537 585
R299 B.n537 B.n536 585
R300 B.n33 B.n32 585
R301 B.n535 B.n33 585
R302 B.n533 B.n532 585
R303 B.n534 B.n533 585
R304 B.n531 B.n38 585
R305 B.n38 B.n37 585
R306 B.n530 B.n529 585
R307 B.n529 B.n528 585
R308 B.n40 B.n39 585
R309 B.n527 B.n40 585
R310 B.n570 B.n569 585
R311 B.n568 B.n2 585
R312 B.n79 B.t12 531.759
R313 B.n77 B.t19 531.759
R314 B.n293 B.t16 531.759
R315 B.n290 B.t8 531.759
R316 B.n81 B.n40 449.257
R317 B.n524 B.n42 449.257
R318 B.n428 B.n253 449.257
R319 B.n425 B.n251 449.257
R320 B.n526 B.n525 256.663
R321 B.n526 B.n75 256.663
R322 B.n526 B.n74 256.663
R323 B.n526 B.n73 256.663
R324 B.n526 B.n72 256.663
R325 B.n526 B.n71 256.663
R326 B.n526 B.n70 256.663
R327 B.n526 B.n69 256.663
R328 B.n526 B.n68 256.663
R329 B.n526 B.n67 256.663
R330 B.n526 B.n66 256.663
R331 B.n526 B.n65 256.663
R332 B.n526 B.n64 256.663
R333 B.n526 B.n63 256.663
R334 B.n526 B.n62 256.663
R335 B.n526 B.n61 256.663
R336 B.n526 B.n60 256.663
R337 B.n526 B.n59 256.663
R338 B.n526 B.n58 256.663
R339 B.n526 B.n57 256.663
R340 B.n526 B.n56 256.663
R341 B.n526 B.n55 256.663
R342 B.n526 B.n54 256.663
R343 B.n526 B.n53 256.663
R344 B.n526 B.n52 256.663
R345 B.n526 B.n51 256.663
R346 B.n526 B.n50 256.663
R347 B.n526 B.n49 256.663
R348 B.n526 B.n48 256.663
R349 B.n526 B.n47 256.663
R350 B.n526 B.n46 256.663
R351 B.n526 B.n45 256.663
R352 B.n526 B.n44 256.663
R353 B.n526 B.n43 256.663
R354 B.n427 B.n426 256.663
R355 B.n427 B.n256 256.663
R356 B.n427 B.n257 256.663
R357 B.n427 B.n258 256.663
R358 B.n427 B.n259 256.663
R359 B.n427 B.n260 256.663
R360 B.n427 B.n261 256.663
R361 B.n427 B.n262 256.663
R362 B.n427 B.n263 256.663
R363 B.n427 B.n264 256.663
R364 B.n427 B.n265 256.663
R365 B.n427 B.n266 256.663
R366 B.n427 B.n267 256.663
R367 B.n427 B.n268 256.663
R368 B.n427 B.n269 256.663
R369 B.n427 B.n270 256.663
R370 B.n427 B.n271 256.663
R371 B.n427 B.n272 256.663
R372 B.n427 B.n273 256.663
R373 B.n427 B.n274 256.663
R374 B.n427 B.n275 256.663
R375 B.n427 B.n276 256.663
R376 B.n427 B.n277 256.663
R377 B.n427 B.n278 256.663
R378 B.n427 B.n279 256.663
R379 B.n427 B.n280 256.663
R380 B.n427 B.n281 256.663
R381 B.n427 B.n282 256.663
R382 B.n427 B.n283 256.663
R383 B.n427 B.n284 256.663
R384 B.n427 B.n285 256.663
R385 B.n427 B.n286 256.663
R386 B.n427 B.n287 256.663
R387 B.n572 B.n571 256.663
R388 B.n85 B.n84 163.367
R389 B.n89 B.n88 163.367
R390 B.n93 B.n92 163.367
R391 B.n97 B.n96 163.367
R392 B.n101 B.n100 163.367
R393 B.n105 B.n104 163.367
R394 B.n109 B.n108 163.367
R395 B.n113 B.n112 163.367
R396 B.n117 B.n116 163.367
R397 B.n121 B.n120 163.367
R398 B.n125 B.n124 163.367
R399 B.n129 B.n128 163.367
R400 B.n133 B.n132 163.367
R401 B.n137 B.n136 163.367
R402 B.n142 B.n141 163.367
R403 B.n146 B.n145 163.367
R404 B.n150 B.n149 163.367
R405 B.n154 B.n153 163.367
R406 B.n158 B.n157 163.367
R407 B.n163 B.n162 163.367
R408 B.n167 B.n166 163.367
R409 B.n171 B.n170 163.367
R410 B.n175 B.n174 163.367
R411 B.n179 B.n178 163.367
R412 B.n183 B.n182 163.367
R413 B.n187 B.n186 163.367
R414 B.n191 B.n190 163.367
R415 B.n195 B.n194 163.367
R416 B.n199 B.n198 163.367
R417 B.n203 B.n202 163.367
R418 B.n207 B.n206 163.367
R419 B.n211 B.n210 163.367
R420 B.n213 B.n76 163.367
R421 B.n432 B.n253 163.367
R422 B.n432 B.n246 163.367
R423 B.n440 B.n246 163.367
R424 B.n440 B.n244 163.367
R425 B.n444 B.n244 163.367
R426 B.n444 B.n239 163.367
R427 B.n452 B.n239 163.367
R428 B.n452 B.n237 163.367
R429 B.n456 B.n237 163.367
R430 B.n456 B.n232 163.367
R431 B.n465 B.n232 163.367
R432 B.n465 B.n230 163.367
R433 B.n469 B.n230 163.367
R434 B.n469 B.n224 163.367
R435 B.n477 B.n224 163.367
R436 B.n477 B.n222 163.367
R437 B.n482 B.n222 163.367
R438 B.n482 B.n217 163.367
R439 B.n491 B.n217 163.367
R440 B.n492 B.n491 163.367
R441 B.n492 B.n5 163.367
R442 B.n6 B.n5 163.367
R443 B.n7 B.n6 163.367
R444 B.n498 B.n7 163.367
R445 B.n499 B.n498 163.367
R446 B.n499 B.n13 163.367
R447 B.n14 B.n13 163.367
R448 B.n15 B.n14 163.367
R449 B.n504 B.n15 163.367
R450 B.n504 B.n20 163.367
R451 B.n21 B.n20 163.367
R452 B.n22 B.n21 163.367
R453 B.n509 B.n22 163.367
R454 B.n509 B.n27 163.367
R455 B.n28 B.n27 163.367
R456 B.n29 B.n28 163.367
R457 B.n514 B.n29 163.367
R458 B.n514 B.n34 163.367
R459 B.n35 B.n34 163.367
R460 B.n36 B.n35 163.367
R461 B.n519 B.n36 163.367
R462 B.n519 B.n41 163.367
R463 B.n42 B.n41 163.367
R464 B.n289 B.n288 163.367
R465 B.n420 B.n288 163.367
R466 B.n418 B.n417 163.367
R467 B.n414 B.n413 163.367
R468 B.n410 B.n409 163.367
R469 B.n406 B.n405 163.367
R470 B.n402 B.n401 163.367
R471 B.n398 B.n397 163.367
R472 B.n394 B.n393 163.367
R473 B.n390 B.n389 163.367
R474 B.n386 B.n385 163.367
R475 B.n382 B.n381 163.367
R476 B.n378 B.n377 163.367
R477 B.n374 B.n373 163.367
R478 B.n370 B.n369 163.367
R479 B.n366 B.n365 163.367
R480 B.n362 B.n361 163.367
R481 B.n358 B.n357 163.367
R482 B.n354 B.n353 163.367
R483 B.n350 B.n349 163.367
R484 B.n346 B.n345 163.367
R485 B.n342 B.n341 163.367
R486 B.n338 B.n337 163.367
R487 B.n334 B.n333 163.367
R488 B.n330 B.n329 163.367
R489 B.n326 B.n325 163.367
R490 B.n322 B.n321 163.367
R491 B.n318 B.n317 163.367
R492 B.n314 B.n313 163.367
R493 B.n310 B.n309 163.367
R494 B.n306 B.n305 163.367
R495 B.n302 B.n301 163.367
R496 B.n298 B.n297 163.367
R497 B.n428 B.n255 163.367
R498 B.n434 B.n251 163.367
R499 B.n434 B.n249 163.367
R500 B.n438 B.n249 163.367
R501 B.n438 B.n243 163.367
R502 B.n446 B.n243 163.367
R503 B.n446 B.n241 163.367
R504 B.n450 B.n241 163.367
R505 B.n450 B.n235 163.367
R506 B.n459 B.n235 163.367
R507 B.n459 B.n233 163.367
R508 B.n463 B.n233 163.367
R509 B.n463 B.n228 163.367
R510 B.n471 B.n228 163.367
R511 B.n471 B.n226 163.367
R512 B.n475 B.n226 163.367
R513 B.n475 B.n220 163.367
R514 B.n485 B.n220 163.367
R515 B.n485 B.n218 163.367
R516 B.n489 B.n218 163.367
R517 B.n489 B.n3 163.367
R518 B.n570 B.n3 163.367
R519 B.n566 B.n2 163.367
R520 B.n566 B.n565 163.367
R521 B.n565 B.n9 163.367
R522 B.n561 B.n9 163.367
R523 B.n561 B.n11 163.367
R524 B.n557 B.n11 163.367
R525 B.n557 B.n17 163.367
R526 B.n553 B.n17 163.367
R527 B.n553 B.n19 163.367
R528 B.n549 B.n19 163.367
R529 B.n549 B.n23 163.367
R530 B.n545 B.n23 163.367
R531 B.n545 B.n25 163.367
R532 B.n541 B.n25 163.367
R533 B.n541 B.n31 163.367
R534 B.n537 B.n31 163.367
R535 B.n537 B.n33 163.367
R536 B.n533 B.n33 163.367
R537 B.n533 B.n38 163.367
R538 B.n529 B.n38 163.367
R539 B.n529 B.n40 163.367
R540 B.n427 B.n252 95.5791
R541 B.n527 B.n526 95.5791
R542 B.n77 B.t20 90.9993
R543 B.n293 B.t18 90.9993
R544 B.n79 B.t14 90.9905
R545 B.n290 B.t11 90.9905
R546 B.n78 B.t21 73.5447
R547 B.n294 B.t17 73.5447
R548 B.n80 B.t15 73.536
R549 B.n291 B.t10 73.536
R550 B.n81 B.n43 71.676
R551 B.n85 B.n44 71.676
R552 B.n89 B.n45 71.676
R553 B.n93 B.n46 71.676
R554 B.n97 B.n47 71.676
R555 B.n101 B.n48 71.676
R556 B.n105 B.n49 71.676
R557 B.n109 B.n50 71.676
R558 B.n113 B.n51 71.676
R559 B.n117 B.n52 71.676
R560 B.n121 B.n53 71.676
R561 B.n125 B.n54 71.676
R562 B.n129 B.n55 71.676
R563 B.n133 B.n56 71.676
R564 B.n137 B.n57 71.676
R565 B.n142 B.n58 71.676
R566 B.n146 B.n59 71.676
R567 B.n150 B.n60 71.676
R568 B.n154 B.n61 71.676
R569 B.n158 B.n62 71.676
R570 B.n163 B.n63 71.676
R571 B.n167 B.n64 71.676
R572 B.n171 B.n65 71.676
R573 B.n175 B.n66 71.676
R574 B.n179 B.n67 71.676
R575 B.n183 B.n68 71.676
R576 B.n187 B.n69 71.676
R577 B.n191 B.n70 71.676
R578 B.n195 B.n71 71.676
R579 B.n199 B.n72 71.676
R580 B.n203 B.n73 71.676
R581 B.n207 B.n74 71.676
R582 B.n211 B.n75 71.676
R583 B.n525 B.n76 71.676
R584 B.n525 B.n524 71.676
R585 B.n213 B.n75 71.676
R586 B.n210 B.n74 71.676
R587 B.n206 B.n73 71.676
R588 B.n202 B.n72 71.676
R589 B.n198 B.n71 71.676
R590 B.n194 B.n70 71.676
R591 B.n190 B.n69 71.676
R592 B.n186 B.n68 71.676
R593 B.n182 B.n67 71.676
R594 B.n178 B.n66 71.676
R595 B.n174 B.n65 71.676
R596 B.n170 B.n64 71.676
R597 B.n166 B.n63 71.676
R598 B.n162 B.n62 71.676
R599 B.n157 B.n61 71.676
R600 B.n153 B.n60 71.676
R601 B.n149 B.n59 71.676
R602 B.n145 B.n58 71.676
R603 B.n141 B.n57 71.676
R604 B.n136 B.n56 71.676
R605 B.n132 B.n55 71.676
R606 B.n128 B.n54 71.676
R607 B.n124 B.n53 71.676
R608 B.n120 B.n52 71.676
R609 B.n116 B.n51 71.676
R610 B.n112 B.n50 71.676
R611 B.n108 B.n49 71.676
R612 B.n104 B.n48 71.676
R613 B.n100 B.n47 71.676
R614 B.n96 B.n46 71.676
R615 B.n92 B.n45 71.676
R616 B.n88 B.n44 71.676
R617 B.n84 B.n43 71.676
R618 B.n426 B.n425 71.676
R619 B.n420 B.n256 71.676
R620 B.n417 B.n257 71.676
R621 B.n413 B.n258 71.676
R622 B.n409 B.n259 71.676
R623 B.n405 B.n260 71.676
R624 B.n401 B.n261 71.676
R625 B.n397 B.n262 71.676
R626 B.n393 B.n263 71.676
R627 B.n389 B.n264 71.676
R628 B.n385 B.n265 71.676
R629 B.n381 B.n266 71.676
R630 B.n377 B.n267 71.676
R631 B.n373 B.n268 71.676
R632 B.n369 B.n269 71.676
R633 B.n365 B.n270 71.676
R634 B.n361 B.n271 71.676
R635 B.n357 B.n272 71.676
R636 B.n353 B.n273 71.676
R637 B.n349 B.n274 71.676
R638 B.n345 B.n275 71.676
R639 B.n341 B.n276 71.676
R640 B.n337 B.n277 71.676
R641 B.n333 B.n278 71.676
R642 B.n329 B.n279 71.676
R643 B.n325 B.n280 71.676
R644 B.n321 B.n281 71.676
R645 B.n317 B.n282 71.676
R646 B.n313 B.n283 71.676
R647 B.n309 B.n284 71.676
R648 B.n305 B.n285 71.676
R649 B.n301 B.n286 71.676
R650 B.n297 B.n287 71.676
R651 B.n426 B.n289 71.676
R652 B.n418 B.n256 71.676
R653 B.n414 B.n257 71.676
R654 B.n410 B.n258 71.676
R655 B.n406 B.n259 71.676
R656 B.n402 B.n260 71.676
R657 B.n398 B.n261 71.676
R658 B.n394 B.n262 71.676
R659 B.n390 B.n263 71.676
R660 B.n386 B.n264 71.676
R661 B.n382 B.n265 71.676
R662 B.n378 B.n266 71.676
R663 B.n374 B.n267 71.676
R664 B.n370 B.n268 71.676
R665 B.n366 B.n269 71.676
R666 B.n362 B.n270 71.676
R667 B.n358 B.n271 71.676
R668 B.n354 B.n272 71.676
R669 B.n350 B.n273 71.676
R670 B.n346 B.n274 71.676
R671 B.n342 B.n275 71.676
R672 B.n338 B.n276 71.676
R673 B.n334 B.n277 71.676
R674 B.n330 B.n278 71.676
R675 B.n326 B.n279 71.676
R676 B.n322 B.n280 71.676
R677 B.n318 B.n281 71.676
R678 B.n314 B.n282 71.676
R679 B.n310 B.n283 71.676
R680 B.n306 B.n284 71.676
R681 B.n302 B.n285 71.676
R682 B.n298 B.n286 71.676
R683 B.n287 B.n255 71.676
R684 B.n571 B.n570 71.676
R685 B.n571 B.n2 71.676
R686 B.n139 B.n80 59.5399
R687 B.n160 B.n78 59.5399
R688 B.n295 B.n294 59.5399
R689 B.n292 B.n291 59.5399
R690 B.n433 B.n252 57.5168
R691 B.n433 B.n247 57.5168
R692 B.n439 B.n247 57.5168
R693 B.n439 B.n248 57.5168
R694 B.n445 B.n240 57.5168
R695 B.n451 B.n240 57.5168
R696 B.n451 B.n236 57.5168
R697 B.n458 B.n236 57.5168
R698 B.n458 B.n457 57.5168
R699 B.n464 B.n229 57.5168
R700 B.n470 B.n229 57.5168
R701 B.n476 B.n225 57.5168
R702 B.n484 B.n221 57.5168
R703 B.n484 B.n483 57.5168
R704 B.n490 B.n4 57.5168
R705 B.n569 B.n4 57.5168
R706 B.n569 B.n568 57.5168
R707 B.n568 B.n567 57.5168
R708 B.n567 B.n8 57.5168
R709 B.n560 B.n12 57.5168
R710 B.n560 B.n559 57.5168
R711 B.n558 B.n16 57.5168
R712 B.n552 B.n551 57.5168
R713 B.n551 B.n550 57.5168
R714 B.n544 B.n26 57.5168
R715 B.n544 B.n543 57.5168
R716 B.n543 B.n542 57.5168
R717 B.n542 B.n30 57.5168
R718 B.n536 B.n30 57.5168
R719 B.n535 B.n534 57.5168
R720 B.n534 B.n37 57.5168
R721 B.n528 B.n37 57.5168
R722 B.n528 B.n527 57.5168
R723 B.n476 B.t5 53.2877
R724 B.t1 B.n558 53.2877
R725 B.n248 B.t9 44.8294
R726 B.t13 B.n535 44.8294
R727 B.t4 B.n225 41.4461
R728 B.t3 B.n16 41.4461
R729 B.n457 B.t6 36.3711
R730 B.n26 B.t7 36.3711
R731 B.n483 B.t0 32.9878
R732 B.n12 B.t2 32.9878
R733 B.n424 B.n250 29.1907
R734 B.n430 B.n429 29.1907
R735 B.n523 B.n522 29.1907
R736 B.n82 B.n39 29.1907
R737 B.n490 B.t0 24.5295
R738 B.t2 B.n8 24.5295
R739 B.n464 B.t6 21.1462
R740 B.n550 B.t7 21.1462
R741 B B.n572 18.0485
R742 B.n80 B.n79 17.455
R743 B.n78 B.n77 17.455
R744 B.n294 B.n293 17.455
R745 B.n291 B.n290 17.455
R746 B.n470 B.t4 16.0712
R747 B.n552 B.t3 16.0712
R748 B.n445 B.t9 12.6879
R749 B.n536 B.t13 12.6879
R750 B.n435 B.n250 10.6151
R751 B.n436 B.n435 10.6151
R752 B.n437 B.n436 10.6151
R753 B.n437 B.n242 10.6151
R754 B.n447 B.n242 10.6151
R755 B.n448 B.n447 10.6151
R756 B.n449 B.n448 10.6151
R757 B.n449 B.n234 10.6151
R758 B.n460 B.n234 10.6151
R759 B.n461 B.n460 10.6151
R760 B.n462 B.n461 10.6151
R761 B.n462 B.n227 10.6151
R762 B.n472 B.n227 10.6151
R763 B.n473 B.n472 10.6151
R764 B.n474 B.n473 10.6151
R765 B.n474 B.n219 10.6151
R766 B.n486 B.n219 10.6151
R767 B.n487 B.n486 10.6151
R768 B.n488 B.n487 10.6151
R769 B.n488 B.n0 10.6151
R770 B.n424 B.n423 10.6151
R771 B.n423 B.n422 10.6151
R772 B.n422 B.n421 10.6151
R773 B.n421 B.n419 10.6151
R774 B.n419 B.n416 10.6151
R775 B.n416 B.n415 10.6151
R776 B.n415 B.n412 10.6151
R777 B.n412 B.n411 10.6151
R778 B.n411 B.n408 10.6151
R779 B.n408 B.n407 10.6151
R780 B.n407 B.n404 10.6151
R781 B.n404 B.n403 10.6151
R782 B.n403 B.n400 10.6151
R783 B.n400 B.n399 10.6151
R784 B.n399 B.n396 10.6151
R785 B.n396 B.n395 10.6151
R786 B.n395 B.n392 10.6151
R787 B.n392 B.n391 10.6151
R788 B.n391 B.n388 10.6151
R789 B.n388 B.n387 10.6151
R790 B.n387 B.n384 10.6151
R791 B.n384 B.n383 10.6151
R792 B.n383 B.n380 10.6151
R793 B.n380 B.n379 10.6151
R794 B.n379 B.n376 10.6151
R795 B.n376 B.n375 10.6151
R796 B.n375 B.n372 10.6151
R797 B.n372 B.n371 10.6151
R798 B.n368 B.n367 10.6151
R799 B.n367 B.n364 10.6151
R800 B.n364 B.n363 10.6151
R801 B.n363 B.n360 10.6151
R802 B.n360 B.n359 10.6151
R803 B.n359 B.n356 10.6151
R804 B.n356 B.n355 10.6151
R805 B.n355 B.n352 10.6151
R806 B.n352 B.n351 10.6151
R807 B.n348 B.n347 10.6151
R808 B.n347 B.n344 10.6151
R809 B.n344 B.n343 10.6151
R810 B.n343 B.n340 10.6151
R811 B.n340 B.n339 10.6151
R812 B.n339 B.n336 10.6151
R813 B.n336 B.n335 10.6151
R814 B.n335 B.n332 10.6151
R815 B.n332 B.n331 10.6151
R816 B.n331 B.n328 10.6151
R817 B.n328 B.n327 10.6151
R818 B.n327 B.n324 10.6151
R819 B.n324 B.n323 10.6151
R820 B.n323 B.n320 10.6151
R821 B.n320 B.n319 10.6151
R822 B.n319 B.n316 10.6151
R823 B.n316 B.n315 10.6151
R824 B.n315 B.n312 10.6151
R825 B.n312 B.n311 10.6151
R826 B.n311 B.n308 10.6151
R827 B.n308 B.n307 10.6151
R828 B.n307 B.n304 10.6151
R829 B.n304 B.n303 10.6151
R830 B.n303 B.n300 10.6151
R831 B.n300 B.n299 10.6151
R832 B.n299 B.n296 10.6151
R833 B.n296 B.n254 10.6151
R834 B.n429 B.n254 10.6151
R835 B.n431 B.n430 10.6151
R836 B.n431 B.n245 10.6151
R837 B.n441 B.n245 10.6151
R838 B.n442 B.n441 10.6151
R839 B.n443 B.n442 10.6151
R840 B.n443 B.n238 10.6151
R841 B.n453 B.n238 10.6151
R842 B.n454 B.n453 10.6151
R843 B.n455 B.n454 10.6151
R844 B.n455 B.n231 10.6151
R845 B.n466 B.n231 10.6151
R846 B.n467 B.n466 10.6151
R847 B.n468 B.n467 10.6151
R848 B.n468 B.n223 10.6151
R849 B.n478 B.n223 10.6151
R850 B.n479 B.n478 10.6151
R851 B.n481 B.n479 10.6151
R852 B.n481 B.n480 10.6151
R853 B.n480 B.n216 10.6151
R854 B.n493 B.n216 10.6151
R855 B.n494 B.n493 10.6151
R856 B.n495 B.n494 10.6151
R857 B.n496 B.n495 10.6151
R858 B.n497 B.n496 10.6151
R859 B.n500 B.n497 10.6151
R860 B.n501 B.n500 10.6151
R861 B.n502 B.n501 10.6151
R862 B.n503 B.n502 10.6151
R863 B.n505 B.n503 10.6151
R864 B.n506 B.n505 10.6151
R865 B.n507 B.n506 10.6151
R866 B.n508 B.n507 10.6151
R867 B.n510 B.n508 10.6151
R868 B.n511 B.n510 10.6151
R869 B.n512 B.n511 10.6151
R870 B.n513 B.n512 10.6151
R871 B.n515 B.n513 10.6151
R872 B.n516 B.n515 10.6151
R873 B.n517 B.n516 10.6151
R874 B.n518 B.n517 10.6151
R875 B.n520 B.n518 10.6151
R876 B.n521 B.n520 10.6151
R877 B.n522 B.n521 10.6151
R878 B.n564 B.n1 10.6151
R879 B.n564 B.n563 10.6151
R880 B.n563 B.n562 10.6151
R881 B.n562 B.n10 10.6151
R882 B.n556 B.n10 10.6151
R883 B.n556 B.n555 10.6151
R884 B.n555 B.n554 10.6151
R885 B.n554 B.n18 10.6151
R886 B.n548 B.n18 10.6151
R887 B.n548 B.n547 10.6151
R888 B.n547 B.n546 10.6151
R889 B.n546 B.n24 10.6151
R890 B.n540 B.n24 10.6151
R891 B.n540 B.n539 10.6151
R892 B.n539 B.n538 10.6151
R893 B.n538 B.n32 10.6151
R894 B.n532 B.n32 10.6151
R895 B.n532 B.n531 10.6151
R896 B.n531 B.n530 10.6151
R897 B.n530 B.n39 10.6151
R898 B.n83 B.n82 10.6151
R899 B.n86 B.n83 10.6151
R900 B.n87 B.n86 10.6151
R901 B.n90 B.n87 10.6151
R902 B.n91 B.n90 10.6151
R903 B.n94 B.n91 10.6151
R904 B.n95 B.n94 10.6151
R905 B.n98 B.n95 10.6151
R906 B.n99 B.n98 10.6151
R907 B.n102 B.n99 10.6151
R908 B.n103 B.n102 10.6151
R909 B.n106 B.n103 10.6151
R910 B.n107 B.n106 10.6151
R911 B.n110 B.n107 10.6151
R912 B.n111 B.n110 10.6151
R913 B.n114 B.n111 10.6151
R914 B.n115 B.n114 10.6151
R915 B.n118 B.n115 10.6151
R916 B.n119 B.n118 10.6151
R917 B.n122 B.n119 10.6151
R918 B.n123 B.n122 10.6151
R919 B.n126 B.n123 10.6151
R920 B.n127 B.n126 10.6151
R921 B.n130 B.n127 10.6151
R922 B.n131 B.n130 10.6151
R923 B.n134 B.n131 10.6151
R924 B.n135 B.n134 10.6151
R925 B.n138 B.n135 10.6151
R926 B.n143 B.n140 10.6151
R927 B.n144 B.n143 10.6151
R928 B.n147 B.n144 10.6151
R929 B.n148 B.n147 10.6151
R930 B.n151 B.n148 10.6151
R931 B.n152 B.n151 10.6151
R932 B.n155 B.n152 10.6151
R933 B.n156 B.n155 10.6151
R934 B.n159 B.n156 10.6151
R935 B.n164 B.n161 10.6151
R936 B.n165 B.n164 10.6151
R937 B.n168 B.n165 10.6151
R938 B.n169 B.n168 10.6151
R939 B.n172 B.n169 10.6151
R940 B.n173 B.n172 10.6151
R941 B.n176 B.n173 10.6151
R942 B.n177 B.n176 10.6151
R943 B.n180 B.n177 10.6151
R944 B.n181 B.n180 10.6151
R945 B.n184 B.n181 10.6151
R946 B.n185 B.n184 10.6151
R947 B.n188 B.n185 10.6151
R948 B.n189 B.n188 10.6151
R949 B.n192 B.n189 10.6151
R950 B.n193 B.n192 10.6151
R951 B.n196 B.n193 10.6151
R952 B.n197 B.n196 10.6151
R953 B.n200 B.n197 10.6151
R954 B.n201 B.n200 10.6151
R955 B.n204 B.n201 10.6151
R956 B.n205 B.n204 10.6151
R957 B.n208 B.n205 10.6151
R958 B.n209 B.n208 10.6151
R959 B.n212 B.n209 10.6151
R960 B.n214 B.n212 10.6151
R961 B.n215 B.n214 10.6151
R962 B.n523 B.n215 10.6151
R963 B.n371 B.n292 9.36635
R964 B.n348 B.n295 9.36635
R965 B.n139 B.n138 9.36635
R966 B.n161 B.n160 9.36635
R967 B.n572 B.n0 8.11757
R968 B.n572 B.n1 8.11757
R969 B.t5 B.n221 4.22964
R970 B.n559 B.t1 4.22964
R971 B.n368 B.n292 1.24928
R972 B.n351 B.n295 1.24928
R973 B.n140 B.n139 1.24928
R974 B.n160 B.n159 1.24928
R975 VP.n4 VP.t6 422.529
R976 VP.n11 VP.t0 396.171
R977 VP.n1 VP.t1 396.171
R978 VP.n16 VP.t7 396.171
R979 VP.n18 VP.t3 396.171
R980 VP.n8 VP.t2 396.171
R981 VP.n6 VP.t4 396.171
R982 VP.n5 VP.t5 396.171
R983 VP.n19 VP.n18 161.3
R984 VP.n6 VP.n3 161.3
R985 VP.n7 VP.n2 161.3
R986 VP.n9 VP.n8 161.3
R987 VP.n17 VP.n0 161.3
R988 VP.n16 VP.n15 161.3
R989 VP.n14 VP.n1 161.3
R990 VP.n13 VP.n12 161.3
R991 VP.n11 VP.n10 161.3
R992 VP.n16 VP.n1 48.2005
R993 VP.n6 VP.n5 48.2005
R994 VP.n12 VP.n11 46.0096
R995 VP.n18 VP.n17 46.0096
R996 VP.n8 VP.n7 46.0096
R997 VP.n4 VP.n3 45.0871
R998 VP.n10 VP.n9 38.1596
R999 VP.n5 VP.n4 14.1472
R1000 VP.n12 VP.n1 2.19141
R1001 VP.n17 VP.n16 2.19141
R1002 VP.n7 VP.n6 2.19141
R1003 VP.n3 VP.n2 0.189894
R1004 VP.n9 VP.n2 0.189894
R1005 VP.n13 VP.n10 0.189894
R1006 VP.n14 VP.n13 0.189894
R1007 VP.n15 VP.n14 0.189894
R1008 VP.n15 VP.n0 0.189894
R1009 VP.n19 VP.n0 0.189894
R1010 VP VP.n19 0.0516364
R1011 VDD1 VDD1.n0 63.9212
R1012 VDD1.n3 VDD1.n2 63.8076
R1013 VDD1.n3 VDD1.n1 63.8076
R1014 VDD1.n5 VDD1.n4 63.475
R1015 VDD1.n5 VDD1.n3 34.4535
R1016 VDD1.n4 VDD1.t4 2.56195
R1017 VDD1.n4 VDD1.t2 2.56195
R1018 VDD1.n0 VDD1.t6 2.56195
R1019 VDD1.n0 VDD1.t5 2.56195
R1020 VDD1.n2 VDD1.t7 2.56195
R1021 VDD1.n2 VDD1.t3 2.56195
R1022 VDD1.n1 VDD1.t0 2.56195
R1023 VDD1.n1 VDD1.t1 2.56195
R1024 VDD1 VDD1.n5 0.330241
R1025 VTAIL.n14 VTAIL.t13 49.3577
R1026 VTAIL.n11 VTAIL.t9 49.3577
R1027 VTAIL.n10 VTAIL.t5 49.3577
R1028 VTAIL.n7 VTAIL.t3 49.3577
R1029 VTAIL.n15 VTAIL.t4 49.3575
R1030 VTAIL.n2 VTAIL.t1 49.3575
R1031 VTAIL.n3 VTAIL.t12 49.3575
R1032 VTAIL.n6 VTAIL.t15 49.3575
R1033 VTAIL.n13 VTAIL.n12 46.7963
R1034 VTAIL.n9 VTAIL.n8 46.7963
R1035 VTAIL.n1 VTAIL.n0 46.7962
R1036 VTAIL.n5 VTAIL.n4 46.7962
R1037 VTAIL.n15 VTAIL.n14 19.8065
R1038 VTAIL.n7 VTAIL.n6 19.8065
R1039 VTAIL.n0 VTAIL.t0 2.56195
R1040 VTAIL.n0 VTAIL.t7 2.56195
R1041 VTAIL.n4 VTAIL.t14 2.56195
R1042 VTAIL.n4 VTAIL.t8 2.56195
R1043 VTAIL.n12 VTAIL.t10 2.56195
R1044 VTAIL.n12 VTAIL.t11 2.56195
R1045 VTAIL.n8 VTAIL.t2 2.56195
R1046 VTAIL.n8 VTAIL.t6 2.56195
R1047 VTAIL.n9 VTAIL.n7 0.776362
R1048 VTAIL.n10 VTAIL.n9 0.776362
R1049 VTAIL.n13 VTAIL.n11 0.776362
R1050 VTAIL.n14 VTAIL.n13 0.776362
R1051 VTAIL.n6 VTAIL.n5 0.776362
R1052 VTAIL.n5 VTAIL.n3 0.776362
R1053 VTAIL.n2 VTAIL.n1 0.776362
R1054 VTAIL VTAIL.n15 0.718172
R1055 VTAIL.n11 VTAIL.n10 0.470328
R1056 VTAIL.n3 VTAIL.n2 0.470328
R1057 VTAIL VTAIL.n1 0.0586897
R1058 VN.n2 VN.t1 422.529
R1059 VN.n10 VN.t5 422.529
R1060 VN.n1 VN.t3 396.171
R1061 VN.n4 VN.t7 396.171
R1062 VN.n6 VN.t6 396.171
R1063 VN.n9 VN.t4 396.171
R1064 VN.n12 VN.t2 396.171
R1065 VN.n14 VN.t0 396.171
R1066 VN.n7 VN.n6 161.3
R1067 VN.n15 VN.n14 161.3
R1068 VN.n13 VN.n8 161.3
R1069 VN.n12 VN.n11 161.3
R1070 VN.n5 VN.n0 161.3
R1071 VN.n4 VN.n3 161.3
R1072 VN.n4 VN.n1 48.2005
R1073 VN.n12 VN.n9 48.2005
R1074 VN.n6 VN.n5 46.0096
R1075 VN.n14 VN.n13 46.0096
R1076 VN.n11 VN.n10 45.0871
R1077 VN.n3 VN.n2 45.0871
R1078 VN VN.n15 38.5403
R1079 VN.n2 VN.n1 14.1472
R1080 VN.n10 VN.n9 14.1472
R1081 VN.n5 VN.n4 2.19141
R1082 VN.n13 VN.n12 2.19141
R1083 VN.n15 VN.n8 0.189894
R1084 VN.n11 VN.n8 0.189894
R1085 VN.n3 VN.n0 0.189894
R1086 VN.n7 VN.n0 0.189894
R1087 VN VN.n7 0.0516364
R1088 VDD2.n2 VDD2.n1 63.8076
R1089 VDD2.n2 VDD2.n0 63.8076
R1090 VDD2 VDD2.n5 63.8048
R1091 VDD2.n4 VDD2.n3 63.475
R1092 VDD2.n4 VDD2.n2 33.8705
R1093 VDD2.n5 VDD2.t3 2.56195
R1094 VDD2.n5 VDD2.t2 2.56195
R1095 VDD2.n3 VDD2.t7 2.56195
R1096 VDD2.n3 VDD2.t5 2.56195
R1097 VDD2.n1 VDD2.t0 2.56195
R1098 VDD2.n1 VDD2.t1 2.56195
R1099 VDD2.n0 VDD2.t6 2.56195
R1100 VDD2.n0 VDD2.t4 2.56195
R1101 VDD2 VDD2.n4 0.446621
C0 VN VDD2 3.30503f
C1 VP VDD2 0.303626f
C2 VTAIL VDD1 8.54857f
C3 VN VTAIL 3.1779f
C4 VP VTAIL 3.192f
C5 VTAIL VDD2 8.58937f
C6 VN VDD1 0.148026f
C7 VP VDD1 3.46026f
C8 VDD1 VDD2 0.762046f
C9 VN VP 4.39056f
C10 VDD2 B 3.043018f
C11 VDD1 B 3.263824f
C12 VTAIL B 6.420433f
C13 VN B 7.63042f
C14 VP B 5.832883f
C15 VDD2.t6 B 0.171699f
C16 VDD2.t4 B 0.171699f
C17 VDD2.n0 B 1.47269f
C18 VDD2.t0 B 0.171699f
C19 VDD2.t1 B 0.171699f
C20 VDD2.n1 B 1.47269f
C21 VDD2.n2 B 2.07384f
C22 VDD2.t7 B 0.171699f
C23 VDD2.t5 B 0.171699f
C24 VDD2.n3 B 1.47088f
C25 VDD2.n4 B 2.14931f
C26 VDD2.t3 B 0.171699f
C27 VDD2.t2 B 0.171699f
C28 VDD2.n5 B 1.47267f
C29 VN.n0 B 0.047473f
C30 VN.t3 B 0.602371f
C31 VN.n1 B 0.274463f
C32 VN.t1 B 0.618856f
C33 VN.n2 B 0.249413f
C34 VN.n3 B 0.196824f
C35 VN.t7 B 0.602371f
C36 VN.n4 B 0.264748f
C37 VN.n5 B 0.010773f
C38 VN.t6 B 0.602371f
C39 VN.n6 B 0.26387f
C40 VN.n7 B 0.03679f
C41 VN.n8 B 0.047473f
C42 VN.t4 B 0.602371f
C43 VN.n9 B 0.274463f
C44 VN.t2 B 0.602371f
C45 VN.t5 B 0.618856f
C46 VN.n10 B 0.249413f
C47 VN.n11 B 0.196824f
C48 VN.n12 B 0.264748f
C49 VN.n13 B 0.010773f
C50 VN.t0 B 0.602371f
C51 VN.n14 B 0.26387f
C52 VN.n15 B 1.6921f
C53 VTAIL.t0 B 0.131681f
C54 VTAIL.t7 B 0.131681f
C55 VTAIL.n0 B 1.06545f
C56 VTAIL.n1 B 0.271002f
C57 VTAIL.t1 B 1.35748f
C58 VTAIL.n2 B 0.366697f
C59 VTAIL.t12 B 1.35748f
C60 VTAIL.n3 B 0.366697f
C61 VTAIL.t14 B 0.131681f
C62 VTAIL.t8 B 0.131681f
C63 VTAIL.n4 B 1.06545f
C64 VTAIL.n5 B 0.320853f
C65 VTAIL.t15 B 1.35748f
C66 VTAIL.n6 B 1.14366f
C67 VTAIL.t3 B 1.35749f
C68 VTAIL.n7 B 1.14366f
C69 VTAIL.t2 B 0.131681f
C70 VTAIL.t6 B 0.131681f
C71 VTAIL.n8 B 1.06546f
C72 VTAIL.n9 B 0.320851f
C73 VTAIL.t5 B 1.35749f
C74 VTAIL.n10 B 0.366689f
C75 VTAIL.t9 B 1.35749f
C76 VTAIL.n11 B 0.366689f
C77 VTAIL.t10 B 0.131681f
C78 VTAIL.t11 B 0.131681f
C79 VTAIL.n12 B 1.06546f
C80 VTAIL.n13 B 0.320851f
C81 VTAIL.t13 B 1.35749f
C82 VTAIL.n14 B 1.14366f
C83 VTAIL.t4 B 1.35748f
C84 VTAIL.n15 B 1.13962f
C85 VDD1.t6 B 0.171645f
C86 VDD1.t5 B 0.171645f
C87 VDD1.n0 B 1.4729f
C88 VDD1.t0 B 0.171645f
C89 VDD1.t1 B 0.171645f
C90 VDD1.n1 B 1.47222f
C91 VDD1.t7 B 0.171645f
C92 VDD1.t3 B 0.171645f
C93 VDD1.n2 B 1.47222f
C94 VDD1.n3 B 2.13348f
C95 VDD1.t4 B 0.171645f
C96 VDD1.t2 B 0.171645f
C97 VDD1.n4 B 1.47041f
C98 VDD1.n5 B 2.18158f
C99 VP.n0 B 0.048642f
C100 VP.t1 B 0.617202f
C101 VP.n1 B 0.271267f
C102 VP.n2 B 0.048642f
C103 VP.t2 B 0.617202f
C104 VP.t4 B 0.617202f
C105 VP.n3 B 0.201671f
C106 VP.t5 B 0.617202f
C107 VP.t6 B 0.634093f
C108 VP.n4 B 0.255554f
C109 VP.n5 B 0.281221f
C110 VP.n6 B 0.271267f
C111 VP.n7 B 0.011038f
C112 VP.n8 B 0.270367f
C113 VP.n9 B 1.70163f
C114 VP.n10 B 1.74745f
C115 VP.t0 B 0.617202f
C116 VP.n11 B 0.270367f
C117 VP.n12 B 0.011038f
C118 VP.n13 B 0.048642f
C119 VP.n14 B 0.048642f
C120 VP.n15 B 0.048642f
C121 VP.t7 B 0.617202f
C122 VP.n16 B 0.271267f
C123 VP.n17 B 0.011038f
C124 VP.t3 B 0.617202f
C125 VP.n18 B 0.270367f
C126 VP.n19 B 0.037696f
.ends

