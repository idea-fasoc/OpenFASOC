* NGSPICE file created from diff_pair_sample_0994.ext - technology: sky130A

.subckt diff_pair_sample_0994 VTAIL VN VP B VDD2 VDD1
X0 B.t15 B.t13 B.t14 B.t3 sky130_fd_pr__nfet_01v8 ad=5.1831 pd=27.36 as=0 ps=0 w=13.29 l=3.82
X1 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=5.1831 pd=27.36 as=0 ps=0 w=13.29 l=3.82
X2 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=5.1831 pd=27.36 as=0 ps=0 w=13.29 l=3.82
X3 VDD1.t1 VP.t0 VTAIL.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=5.1831 pd=27.36 as=5.1831 ps=27.36 w=13.29 l=3.82
X4 VDD2.t1 VN.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=5.1831 pd=27.36 as=5.1831 ps=27.36 w=13.29 l=3.82
X5 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=5.1831 pd=27.36 as=0 ps=0 w=13.29 l=3.82
X6 VDD1.t0 VP.t1 VTAIL.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=5.1831 pd=27.36 as=5.1831 ps=27.36 w=13.29 l=3.82
X7 VDD2.t0 VN.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=5.1831 pd=27.36 as=5.1831 ps=27.36 w=13.29 l=3.82
R0 B.n771 B.n770 585
R1 B.n313 B.n112 585
R2 B.n312 B.n311 585
R3 B.n310 B.n309 585
R4 B.n308 B.n307 585
R5 B.n306 B.n305 585
R6 B.n304 B.n303 585
R7 B.n302 B.n301 585
R8 B.n300 B.n299 585
R9 B.n298 B.n297 585
R10 B.n296 B.n295 585
R11 B.n294 B.n293 585
R12 B.n292 B.n291 585
R13 B.n290 B.n289 585
R14 B.n288 B.n287 585
R15 B.n286 B.n285 585
R16 B.n284 B.n283 585
R17 B.n282 B.n281 585
R18 B.n280 B.n279 585
R19 B.n278 B.n277 585
R20 B.n276 B.n275 585
R21 B.n274 B.n273 585
R22 B.n272 B.n271 585
R23 B.n270 B.n269 585
R24 B.n268 B.n267 585
R25 B.n266 B.n265 585
R26 B.n264 B.n263 585
R27 B.n262 B.n261 585
R28 B.n260 B.n259 585
R29 B.n258 B.n257 585
R30 B.n256 B.n255 585
R31 B.n254 B.n253 585
R32 B.n252 B.n251 585
R33 B.n250 B.n249 585
R34 B.n248 B.n247 585
R35 B.n246 B.n245 585
R36 B.n244 B.n243 585
R37 B.n242 B.n241 585
R38 B.n240 B.n239 585
R39 B.n238 B.n237 585
R40 B.n236 B.n235 585
R41 B.n234 B.n233 585
R42 B.n232 B.n231 585
R43 B.n230 B.n229 585
R44 B.n228 B.n227 585
R45 B.n225 B.n224 585
R46 B.n223 B.n222 585
R47 B.n221 B.n220 585
R48 B.n219 B.n218 585
R49 B.n217 B.n216 585
R50 B.n215 B.n214 585
R51 B.n213 B.n212 585
R52 B.n211 B.n210 585
R53 B.n209 B.n208 585
R54 B.n207 B.n206 585
R55 B.n204 B.n203 585
R56 B.n202 B.n201 585
R57 B.n200 B.n199 585
R58 B.n198 B.n197 585
R59 B.n196 B.n195 585
R60 B.n194 B.n193 585
R61 B.n192 B.n191 585
R62 B.n190 B.n189 585
R63 B.n188 B.n187 585
R64 B.n186 B.n185 585
R65 B.n184 B.n183 585
R66 B.n182 B.n181 585
R67 B.n180 B.n179 585
R68 B.n178 B.n177 585
R69 B.n176 B.n175 585
R70 B.n174 B.n173 585
R71 B.n172 B.n171 585
R72 B.n170 B.n169 585
R73 B.n168 B.n167 585
R74 B.n166 B.n165 585
R75 B.n164 B.n163 585
R76 B.n162 B.n161 585
R77 B.n160 B.n159 585
R78 B.n158 B.n157 585
R79 B.n156 B.n155 585
R80 B.n154 B.n153 585
R81 B.n152 B.n151 585
R82 B.n150 B.n149 585
R83 B.n148 B.n147 585
R84 B.n146 B.n145 585
R85 B.n144 B.n143 585
R86 B.n142 B.n141 585
R87 B.n140 B.n139 585
R88 B.n138 B.n137 585
R89 B.n136 B.n135 585
R90 B.n134 B.n133 585
R91 B.n132 B.n131 585
R92 B.n130 B.n129 585
R93 B.n128 B.n127 585
R94 B.n126 B.n125 585
R95 B.n124 B.n123 585
R96 B.n122 B.n121 585
R97 B.n120 B.n119 585
R98 B.n118 B.n117 585
R99 B.n61 B.n60 585
R100 B.n769 B.n62 585
R101 B.n774 B.n62 585
R102 B.n768 B.n767 585
R103 B.n767 B.n58 585
R104 B.n766 B.n57 585
R105 B.n780 B.n57 585
R106 B.n765 B.n56 585
R107 B.n781 B.n56 585
R108 B.n764 B.n55 585
R109 B.n782 B.n55 585
R110 B.n763 B.n762 585
R111 B.n762 B.n51 585
R112 B.n761 B.n50 585
R113 B.n788 B.n50 585
R114 B.n760 B.n49 585
R115 B.n789 B.n49 585
R116 B.n759 B.n48 585
R117 B.n790 B.n48 585
R118 B.n758 B.n757 585
R119 B.n757 B.n47 585
R120 B.n756 B.n43 585
R121 B.n796 B.n43 585
R122 B.n755 B.n42 585
R123 B.n797 B.n42 585
R124 B.n754 B.n41 585
R125 B.n798 B.n41 585
R126 B.n753 B.n752 585
R127 B.n752 B.n37 585
R128 B.n751 B.n36 585
R129 B.n804 B.n36 585
R130 B.n750 B.n35 585
R131 B.n805 B.n35 585
R132 B.n749 B.n34 585
R133 B.n806 B.n34 585
R134 B.n748 B.n747 585
R135 B.n747 B.n30 585
R136 B.n746 B.n29 585
R137 B.n812 B.n29 585
R138 B.n745 B.n28 585
R139 B.n813 B.n28 585
R140 B.n744 B.n27 585
R141 B.n814 B.n27 585
R142 B.n743 B.n742 585
R143 B.n742 B.n23 585
R144 B.n741 B.n22 585
R145 B.n820 B.n22 585
R146 B.n740 B.n21 585
R147 B.n821 B.n21 585
R148 B.n739 B.n20 585
R149 B.n822 B.n20 585
R150 B.n738 B.n737 585
R151 B.n737 B.n16 585
R152 B.n736 B.n15 585
R153 B.n828 B.n15 585
R154 B.n735 B.n14 585
R155 B.n829 B.n14 585
R156 B.n734 B.n13 585
R157 B.n830 B.n13 585
R158 B.n733 B.n732 585
R159 B.n732 B.n12 585
R160 B.n731 B.n730 585
R161 B.n731 B.n8 585
R162 B.n729 B.n7 585
R163 B.n837 B.n7 585
R164 B.n728 B.n6 585
R165 B.n838 B.n6 585
R166 B.n727 B.n5 585
R167 B.n839 B.n5 585
R168 B.n726 B.n725 585
R169 B.n725 B.n4 585
R170 B.n724 B.n314 585
R171 B.n724 B.n723 585
R172 B.n714 B.n315 585
R173 B.n316 B.n315 585
R174 B.n716 B.n715 585
R175 B.n717 B.n716 585
R176 B.n713 B.n321 585
R177 B.n321 B.n320 585
R178 B.n712 B.n711 585
R179 B.n711 B.n710 585
R180 B.n323 B.n322 585
R181 B.n324 B.n323 585
R182 B.n703 B.n702 585
R183 B.n704 B.n703 585
R184 B.n701 B.n329 585
R185 B.n329 B.n328 585
R186 B.n700 B.n699 585
R187 B.n699 B.n698 585
R188 B.n331 B.n330 585
R189 B.n332 B.n331 585
R190 B.n691 B.n690 585
R191 B.n692 B.n691 585
R192 B.n689 B.n337 585
R193 B.n337 B.n336 585
R194 B.n688 B.n687 585
R195 B.n687 B.n686 585
R196 B.n339 B.n338 585
R197 B.n340 B.n339 585
R198 B.n679 B.n678 585
R199 B.n680 B.n679 585
R200 B.n677 B.n345 585
R201 B.n345 B.n344 585
R202 B.n676 B.n675 585
R203 B.n675 B.n674 585
R204 B.n347 B.n346 585
R205 B.n348 B.n347 585
R206 B.n667 B.n666 585
R207 B.n668 B.n667 585
R208 B.n665 B.n353 585
R209 B.n353 B.n352 585
R210 B.n664 B.n663 585
R211 B.n663 B.n662 585
R212 B.n355 B.n354 585
R213 B.n655 B.n355 585
R214 B.n654 B.n653 585
R215 B.n656 B.n654 585
R216 B.n652 B.n360 585
R217 B.n360 B.n359 585
R218 B.n651 B.n650 585
R219 B.n650 B.n649 585
R220 B.n362 B.n361 585
R221 B.n363 B.n362 585
R222 B.n642 B.n641 585
R223 B.n643 B.n642 585
R224 B.n640 B.n368 585
R225 B.n368 B.n367 585
R226 B.n639 B.n638 585
R227 B.n638 B.n637 585
R228 B.n370 B.n369 585
R229 B.n371 B.n370 585
R230 B.n630 B.n629 585
R231 B.n631 B.n630 585
R232 B.n374 B.n373 585
R233 B.n433 B.n432 585
R234 B.n434 B.n430 585
R235 B.n430 B.n375 585
R236 B.n436 B.n435 585
R237 B.n438 B.n429 585
R238 B.n441 B.n440 585
R239 B.n442 B.n428 585
R240 B.n444 B.n443 585
R241 B.n446 B.n427 585
R242 B.n449 B.n448 585
R243 B.n450 B.n426 585
R244 B.n452 B.n451 585
R245 B.n454 B.n425 585
R246 B.n457 B.n456 585
R247 B.n458 B.n424 585
R248 B.n460 B.n459 585
R249 B.n462 B.n423 585
R250 B.n465 B.n464 585
R251 B.n466 B.n422 585
R252 B.n468 B.n467 585
R253 B.n470 B.n421 585
R254 B.n473 B.n472 585
R255 B.n474 B.n420 585
R256 B.n476 B.n475 585
R257 B.n478 B.n419 585
R258 B.n481 B.n480 585
R259 B.n482 B.n418 585
R260 B.n484 B.n483 585
R261 B.n486 B.n417 585
R262 B.n489 B.n488 585
R263 B.n490 B.n416 585
R264 B.n492 B.n491 585
R265 B.n494 B.n415 585
R266 B.n497 B.n496 585
R267 B.n498 B.n414 585
R268 B.n500 B.n499 585
R269 B.n502 B.n413 585
R270 B.n505 B.n504 585
R271 B.n506 B.n412 585
R272 B.n508 B.n507 585
R273 B.n510 B.n411 585
R274 B.n513 B.n512 585
R275 B.n514 B.n410 585
R276 B.n516 B.n515 585
R277 B.n518 B.n409 585
R278 B.n521 B.n520 585
R279 B.n522 B.n405 585
R280 B.n524 B.n523 585
R281 B.n526 B.n404 585
R282 B.n529 B.n528 585
R283 B.n530 B.n403 585
R284 B.n532 B.n531 585
R285 B.n534 B.n402 585
R286 B.n537 B.n536 585
R287 B.n538 B.n399 585
R288 B.n541 B.n540 585
R289 B.n543 B.n398 585
R290 B.n546 B.n545 585
R291 B.n547 B.n397 585
R292 B.n549 B.n548 585
R293 B.n551 B.n396 585
R294 B.n554 B.n553 585
R295 B.n555 B.n395 585
R296 B.n557 B.n556 585
R297 B.n559 B.n394 585
R298 B.n562 B.n561 585
R299 B.n563 B.n393 585
R300 B.n565 B.n564 585
R301 B.n567 B.n392 585
R302 B.n570 B.n569 585
R303 B.n571 B.n391 585
R304 B.n573 B.n572 585
R305 B.n575 B.n390 585
R306 B.n578 B.n577 585
R307 B.n579 B.n389 585
R308 B.n581 B.n580 585
R309 B.n583 B.n388 585
R310 B.n586 B.n585 585
R311 B.n587 B.n387 585
R312 B.n589 B.n588 585
R313 B.n591 B.n386 585
R314 B.n594 B.n593 585
R315 B.n595 B.n385 585
R316 B.n597 B.n596 585
R317 B.n599 B.n384 585
R318 B.n602 B.n601 585
R319 B.n603 B.n383 585
R320 B.n605 B.n604 585
R321 B.n607 B.n382 585
R322 B.n610 B.n609 585
R323 B.n611 B.n381 585
R324 B.n613 B.n612 585
R325 B.n615 B.n380 585
R326 B.n618 B.n617 585
R327 B.n619 B.n379 585
R328 B.n621 B.n620 585
R329 B.n623 B.n378 585
R330 B.n624 B.n377 585
R331 B.n627 B.n626 585
R332 B.n628 B.n376 585
R333 B.n376 B.n375 585
R334 B.n633 B.n632 585
R335 B.n632 B.n631 585
R336 B.n634 B.n372 585
R337 B.n372 B.n371 585
R338 B.n636 B.n635 585
R339 B.n637 B.n636 585
R340 B.n366 B.n365 585
R341 B.n367 B.n366 585
R342 B.n645 B.n644 585
R343 B.n644 B.n643 585
R344 B.n646 B.n364 585
R345 B.n364 B.n363 585
R346 B.n648 B.n647 585
R347 B.n649 B.n648 585
R348 B.n358 B.n357 585
R349 B.n359 B.n358 585
R350 B.n658 B.n657 585
R351 B.n657 B.n656 585
R352 B.n659 B.n356 585
R353 B.n655 B.n356 585
R354 B.n661 B.n660 585
R355 B.n662 B.n661 585
R356 B.n351 B.n350 585
R357 B.n352 B.n351 585
R358 B.n670 B.n669 585
R359 B.n669 B.n668 585
R360 B.n671 B.n349 585
R361 B.n349 B.n348 585
R362 B.n673 B.n672 585
R363 B.n674 B.n673 585
R364 B.n343 B.n342 585
R365 B.n344 B.n343 585
R366 B.n682 B.n681 585
R367 B.n681 B.n680 585
R368 B.n683 B.n341 585
R369 B.n341 B.n340 585
R370 B.n685 B.n684 585
R371 B.n686 B.n685 585
R372 B.n335 B.n334 585
R373 B.n336 B.n335 585
R374 B.n694 B.n693 585
R375 B.n693 B.n692 585
R376 B.n695 B.n333 585
R377 B.n333 B.n332 585
R378 B.n697 B.n696 585
R379 B.n698 B.n697 585
R380 B.n327 B.n326 585
R381 B.n328 B.n327 585
R382 B.n706 B.n705 585
R383 B.n705 B.n704 585
R384 B.n707 B.n325 585
R385 B.n325 B.n324 585
R386 B.n709 B.n708 585
R387 B.n710 B.n709 585
R388 B.n319 B.n318 585
R389 B.n320 B.n319 585
R390 B.n719 B.n718 585
R391 B.n718 B.n717 585
R392 B.n720 B.n317 585
R393 B.n317 B.n316 585
R394 B.n722 B.n721 585
R395 B.n723 B.n722 585
R396 B.n3 B.n0 585
R397 B.n4 B.n3 585
R398 B.n836 B.n1 585
R399 B.n837 B.n836 585
R400 B.n835 B.n834 585
R401 B.n835 B.n8 585
R402 B.n833 B.n9 585
R403 B.n12 B.n9 585
R404 B.n832 B.n831 585
R405 B.n831 B.n830 585
R406 B.n11 B.n10 585
R407 B.n829 B.n11 585
R408 B.n827 B.n826 585
R409 B.n828 B.n827 585
R410 B.n825 B.n17 585
R411 B.n17 B.n16 585
R412 B.n824 B.n823 585
R413 B.n823 B.n822 585
R414 B.n19 B.n18 585
R415 B.n821 B.n19 585
R416 B.n819 B.n818 585
R417 B.n820 B.n819 585
R418 B.n817 B.n24 585
R419 B.n24 B.n23 585
R420 B.n816 B.n815 585
R421 B.n815 B.n814 585
R422 B.n26 B.n25 585
R423 B.n813 B.n26 585
R424 B.n811 B.n810 585
R425 B.n812 B.n811 585
R426 B.n809 B.n31 585
R427 B.n31 B.n30 585
R428 B.n808 B.n807 585
R429 B.n807 B.n806 585
R430 B.n33 B.n32 585
R431 B.n805 B.n33 585
R432 B.n803 B.n802 585
R433 B.n804 B.n803 585
R434 B.n801 B.n38 585
R435 B.n38 B.n37 585
R436 B.n800 B.n799 585
R437 B.n799 B.n798 585
R438 B.n40 B.n39 585
R439 B.n797 B.n40 585
R440 B.n795 B.n794 585
R441 B.n796 B.n795 585
R442 B.n793 B.n44 585
R443 B.n47 B.n44 585
R444 B.n792 B.n791 585
R445 B.n791 B.n790 585
R446 B.n46 B.n45 585
R447 B.n789 B.n46 585
R448 B.n787 B.n786 585
R449 B.n788 B.n787 585
R450 B.n785 B.n52 585
R451 B.n52 B.n51 585
R452 B.n784 B.n783 585
R453 B.n783 B.n782 585
R454 B.n54 B.n53 585
R455 B.n781 B.n54 585
R456 B.n779 B.n778 585
R457 B.n780 B.n779 585
R458 B.n777 B.n59 585
R459 B.n59 B.n58 585
R460 B.n776 B.n775 585
R461 B.n775 B.n774 585
R462 B.n840 B.n839 585
R463 B.n838 B.n2 585
R464 B.n775 B.n61 535.745
R465 B.n771 B.n62 535.745
R466 B.n630 B.n376 535.745
R467 B.n632 B.n374 535.745
R468 B.n113 B.t8 384.56
R469 B.n400 B.t5 384.56
R470 B.n115 B.t11 384.56
R471 B.n406 B.t15 384.56
R472 B.n114 B.t9 304.075
R473 B.n401 B.t4 304.075
R474 B.n116 B.t12 304.075
R475 B.n407 B.t14 304.075
R476 B.n115 B.t10 293.204
R477 B.n113 B.t6 293.204
R478 B.n400 B.t2 293.204
R479 B.n406 B.t13 293.204
R480 B.n773 B.n772 256.663
R481 B.n773 B.n111 256.663
R482 B.n773 B.n110 256.663
R483 B.n773 B.n109 256.663
R484 B.n773 B.n108 256.663
R485 B.n773 B.n107 256.663
R486 B.n773 B.n106 256.663
R487 B.n773 B.n105 256.663
R488 B.n773 B.n104 256.663
R489 B.n773 B.n103 256.663
R490 B.n773 B.n102 256.663
R491 B.n773 B.n101 256.663
R492 B.n773 B.n100 256.663
R493 B.n773 B.n99 256.663
R494 B.n773 B.n98 256.663
R495 B.n773 B.n97 256.663
R496 B.n773 B.n96 256.663
R497 B.n773 B.n95 256.663
R498 B.n773 B.n94 256.663
R499 B.n773 B.n93 256.663
R500 B.n773 B.n92 256.663
R501 B.n773 B.n91 256.663
R502 B.n773 B.n90 256.663
R503 B.n773 B.n89 256.663
R504 B.n773 B.n88 256.663
R505 B.n773 B.n87 256.663
R506 B.n773 B.n86 256.663
R507 B.n773 B.n85 256.663
R508 B.n773 B.n84 256.663
R509 B.n773 B.n83 256.663
R510 B.n773 B.n82 256.663
R511 B.n773 B.n81 256.663
R512 B.n773 B.n80 256.663
R513 B.n773 B.n79 256.663
R514 B.n773 B.n78 256.663
R515 B.n773 B.n77 256.663
R516 B.n773 B.n76 256.663
R517 B.n773 B.n75 256.663
R518 B.n773 B.n74 256.663
R519 B.n773 B.n73 256.663
R520 B.n773 B.n72 256.663
R521 B.n773 B.n71 256.663
R522 B.n773 B.n70 256.663
R523 B.n773 B.n69 256.663
R524 B.n773 B.n68 256.663
R525 B.n773 B.n67 256.663
R526 B.n773 B.n66 256.663
R527 B.n773 B.n65 256.663
R528 B.n773 B.n64 256.663
R529 B.n773 B.n63 256.663
R530 B.n431 B.n375 256.663
R531 B.n437 B.n375 256.663
R532 B.n439 B.n375 256.663
R533 B.n445 B.n375 256.663
R534 B.n447 B.n375 256.663
R535 B.n453 B.n375 256.663
R536 B.n455 B.n375 256.663
R537 B.n461 B.n375 256.663
R538 B.n463 B.n375 256.663
R539 B.n469 B.n375 256.663
R540 B.n471 B.n375 256.663
R541 B.n477 B.n375 256.663
R542 B.n479 B.n375 256.663
R543 B.n485 B.n375 256.663
R544 B.n487 B.n375 256.663
R545 B.n493 B.n375 256.663
R546 B.n495 B.n375 256.663
R547 B.n501 B.n375 256.663
R548 B.n503 B.n375 256.663
R549 B.n509 B.n375 256.663
R550 B.n511 B.n375 256.663
R551 B.n517 B.n375 256.663
R552 B.n519 B.n375 256.663
R553 B.n525 B.n375 256.663
R554 B.n527 B.n375 256.663
R555 B.n533 B.n375 256.663
R556 B.n535 B.n375 256.663
R557 B.n542 B.n375 256.663
R558 B.n544 B.n375 256.663
R559 B.n550 B.n375 256.663
R560 B.n552 B.n375 256.663
R561 B.n558 B.n375 256.663
R562 B.n560 B.n375 256.663
R563 B.n566 B.n375 256.663
R564 B.n568 B.n375 256.663
R565 B.n574 B.n375 256.663
R566 B.n576 B.n375 256.663
R567 B.n582 B.n375 256.663
R568 B.n584 B.n375 256.663
R569 B.n590 B.n375 256.663
R570 B.n592 B.n375 256.663
R571 B.n598 B.n375 256.663
R572 B.n600 B.n375 256.663
R573 B.n606 B.n375 256.663
R574 B.n608 B.n375 256.663
R575 B.n614 B.n375 256.663
R576 B.n616 B.n375 256.663
R577 B.n622 B.n375 256.663
R578 B.n625 B.n375 256.663
R579 B.n842 B.n841 256.663
R580 B.n119 B.n118 163.367
R581 B.n123 B.n122 163.367
R582 B.n127 B.n126 163.367
R583 B.n131 B.n130 163.367
R584 B.n135 B.n134 163.367
R585 B.n139 B.n138 163.367
R586 B.n143 B.n142 163.367
R587 B.n147 B.n146 163.367
R588 B.n151 B.n150 163.367
R589 B.n155 B.n154 163.367
R590 B.n159 B.n158 163.367
R591 B.n163 B.n162 163.367
R592 B.n167 B.n166 163.367
R593 B.n171 B.n170 163.367
R594 B.n175 B.n174 163.367
R595 B.n179 B.n178 163.367
R596 B.n183 B.n182 163.367
R597 B.n187 B.n186 163.367
R598 B.n191 B.n190 163.367
R599 B.n195 B.n194 163.367
R600 B.n199 B.n198 163.367
R601 B.n203 B.n202 163.367
R602 B.n208 B.n207 163.367
R603 B.n212 B.n211 163.367
R604 B.n216 B.n215 163.367
R605 B.n220 B.n219 163.367
R606 B.n224 B.n223 163.367
R607 B.n229 B.n228 163.367
R608 B.n233 B.n232 163.367
R609 B.n237 B.n236 163.367
R610 B.n241 B.n240 163.367
R611 B.n245 B.n244 163.367
R612 B.n249 B.n248 163.367
R613 B.n253 B.n252 163.367
R614 B.n257 B.n256 163.367
R615 B.n261 B.n260 163.367
R616 B.n265 B.n264 163.367
R617 B.n269 B.n268 163.367
R618 B.n273 B.n272 163.367
R619 B.n277 B.n276 163.367
R620 B.n281 B.n280 163.367
R621 B.n285 B.n284 163.367
R622 B.n289 B.n288 163.367
R623 B.n293 B.n292 163.367
R624 B.n297 B.n296 163.367
R625 B.n301 B.n300 163.367
R626 B.n305 B.n304 163.367
R627 B.n309 B.n308 163.367
R628 B.n311 B.n112 163.367
R629 B.n630 B.n370 163.367
R630 B.n638 B.n370 163.367
R631 B.n638 B.n368 163.367
R632 B.n642 B.n368 163.367
R633 B.n642 B.n362 163.367
R634 B.n650 B.n362 163.367
R635 B.n650 B.n360 163.367
R636 B.n654 B.n360 163.367
R637 B.n654 B.n355 163.367
R638 B.n663 B.n355 163.367
R639 B.n663 B.n353 163.367
R640 B.n667 B.n353 163.367
R641 B.n667 B.n347 163.367
R642 B.n675 B.n347 163.367
R643 B.n675 B.n345 163.367
R644 B.n679 B.n345 163.367
R645 B.n679 B.n339 163.367
R646 B.n687 B.n339 163.367
R647 B.n687 B.n337 163.367
R648 B.n691 B.n337 163.367
R649 B.n691 B.n331 163.367
R650 B.n699 B.n331 163.367
R651 B.n699 B.n329 163.367
R652 B.n703 B.n329 163.367
R653 B.n703 B.n323 163.367
R654 B.n711 B.n323 163.367
R655 B.n711 B.n321 163.367
R656 B.n716 B.n321 163.367
R657 B.n716 B.n315 163.367
R658 B.n724 B.n315 163.367
R659 B.n725 B.n724 163.367
R660 B.n725 B.n5 163.367
R661 B.n6 B.n5 163.367
R662 B.n7 B.n6 163.367
R663 B.n731 B.n7 163.367
R664 B.n732 B.n731 163.367
R665 B.n732 B.n13 163.367
R666 B.n14 B.n13 163.367
R667 B.n15 B.n14 163.367
R668 B.n737 B.n15 163.367
R669 B.n737 B.n20 163.367
R670 B.n21 B.n20 163.367
R671 B.n22 B.n21 163.367
R672 B.n742 B.n22 163.367
R673 B.n742 B.n27 163.367
R674 B.n28 B.n27 163.367
R675 B.n29 B.n28 163.367
R676 B.n747 B.n29 163.367
R677 B.n747 B.n34 163.367
R678 B.n35 B.n34 163.367
R679 B.n36 B.n35 163.367
R680 B.n752 B.n36 163.367
R681 B.n752 B.n41 163.367
R682 B.n42 B.n41 163.367
R683 B.n43 B.n42 163.367
R684 B.n757 B.n43 163.367
R685 B.n757 B.n48 163.367
R686 B.n49 B.n48 163.367
R687 B.n50 B.n49 163.367
R688 B.n762 B.n50 163.367
R689 B.n762 B.n55 163.367
R690 B.n56 B.n55 163.367
R691 B.n57 B.n56 163.367
R692 B.n767 B.n57 163.367
R693 B.n767 B.n62 163.367
R694 B.n432 B.n430 163.367
R695 B.n436 B.n430 163.367
R696 B.n440 B.n438 163.367
R697 B.n444 B.n428 163.367
R698 B.n448 B.n446 163.367
R699 B.n452 B.n426 163.367
R700 B.n456 B.n454 163.367
R701 B.n460 B.n424 163.367
R702 B.n464 B.n462 163.367
R703 B.n468 B.n422 163.367
R704 B.n472 B.n470 163.367
R705 B.n476 B.n420 163.367
R706 B.n480 B.n478 163.367
R707 B.n484 B.n418 163.367
R708 B.n488 B.n486 163.367
R709 B.n492 B.n416 163.367
R710 B.n496 B.n494 163.367
R711 B.n500 B.n414 163.367
R712 B.n504 B.n502 163.367
R713 B.n508 B.n412 163.367
R714 B.n512 B.n510 163.367
R715 B.n516 B.n410 163.367
R716 B.n520 B.n518 163.367
R717 B.n524 B.n405 163.367
R718 B.n528 B.n526 163.367
R719 B.n532 B.n403 163.367
R720 B.n536 B.n534 163.367
R721 B.n541 B.n399 163.367
R722 B.n545 B.n543 163.367
R723 B.n549 B.n397 163.367
R724 B.n553 B.n551 163.367
R725 B.n557 B.n395 163.367
R726 B.n561 B.n559 163.367
R727 B.n565 B.n393 163.367
R728 B.n569 B.n567 163.367
R729 B.n573 B.n391 163.367
R730 B.n577 B.n575 163.367
R731 B.n581 B.n389 163.367
R732 B.n585 B.n583 163.367
R733 B.n589 B.n387 163.367
R734 B.n593 B.n591 163.367
R735 B.n597 B.n385 163.367
R736 B.n601 B.n599 163.367
R737 B.n605 B.n383 163.367
R738 B.n609 B.n607 163.367
R739 B.n613 B.n381 163.367
R740 B.n617 B.n615 163.367
R741 B.n621 B.n379 163.367
R742 B.n624 B.n623 163.367
R743 B.n626 B.n376 163.367
R744 B.n632 B.n372 163.367
R745 B.n636 B.n372 163.367
R746 B.n636 B.n366 163.367
R747 B.n644 B.n366 163.367
R748 B.n644 B.n364 163.367
R749 B.n648 B.n364 163.367
R750 B.n648 B.n358 163.367
R751 B.n657 B.n358 163.367
R752 B.n657 B.n356 163.367
R753 B.n661 B.n356 163.367
R754 B.n661 B.n351 163.367
R755 B.n669 B.n351 163.367
R756 B.n669 B.n349 163.367
R757 B.n673 B.n349 163.367
R758 B.n673 B.n343 163.367
R759 B.n681 B.n343 163.367
R760 B.n681 B.n341 163.367
R761 B.n685 B.n341 163.367
R762 B.n685 B.n335 163.367
R763 B.n693 B.n335 163.367
R764 B.n693 B.n333 163.367
R765 B.n697 B.n333 163.367
R766 B.n697 B.n327 163.367
R767 B.n705 B.n327 163.367
R768 B.n705 B.n325 163.367
R769 B.n709 B.n325 163.367
R770 B.n709 B.n319 163.367
R771 B.n718 B.n319 163.367
R772 B.n718 B.n317 163.367
R773 B.n722 B.n317 163.367
R774 B.n722 B.n3 163.367
R775 B.n840 B.n3 163.367
R776 B.n836 B.n2 163.367
R777 B.n836 B.n835 163.367
R778 B.n835 B.n9 163.367
R779 B.n831 B.n9 163.367
R780 B.n831 B.n11 163.367
R781 B.n827 B.n11 163.367
R782 B.n827 B.n17 163.367
R783 B.n823 B.n17 163.367
R784 B.n823 B.n19 163.367
R785 B.n819 B.n19 163.367
R786 B.n819 B.n24 163.367
R787 B.n815 B.n24 163.367
R788 B.n815 B.n26 163.367
R789 B.n811 B.n26 163.367
R790 B.n811 B.n31 163.367
R791 B.n807 B.n31 163.367
R792 B.n807 B.n33 163.367
R793 B.n803 B.n33 163.367
R794 B.n803 B.n38 163.367
R795 B.n799 B.n38 163.367
R796 B.n799 B.n40 163.367
R797 B.n795 B.n40 163.367
R798 B.n795 B.n44 163.367
R799 B.n791 B.n44 163.367
R800 B.n791 B.n46 163.367
R801 B.n787 B.n46 163.367
R802 B.n787 B.n52 163.367
R803 B.n783 B.n52 163.367
R804 B.n783 B.n54 163.367
R805 B.n779 B.n54 163.367
R806 B.n779 B.n59 163.367
R807 B.n775 B.n59 163.367
R808 B.n116 B.n115 80.4853
R809 B.n114 B.n113 80.4853
R810 B.n401 B.n400 80.4853
R811 B.n407 B.n406 80.4853
R812 B.n631 B.n375 74.0646
R813 B.n774 B.n773 74.0646
R814 B.n63 B.n61 71.676
R815 B.n119 B.n64 71.676
R816 B.n123 B.n65 71.676
R817 B.n127 B.n66 71.676
R818 B.n131 B.n67 71.676
R819 B.n135 B.n68 71.676
R820 B.n139 B.n69 71.676
R821 B.n143 B.n70 71.676
R822 B.n147 B.n71 71.676
R823 B.n151 B.n72 71.676
R824 B.n155 B.n73 71.676
R825 B.n159 B.n74 71.676
R826 B.n163 B.n75 71.676
R827 B.n167 B.n76 71.676
R828 B.n171 B.n77 71.676
R829 B.n175 B.n78 71.676
R830 B.n179 B.n79 71.676
R831 B.n183 B.n80 71.676
R832 B.n187 B.n81 71.676
R833 B.n191 B.n82 71.676
R834 B.n195 B.n83 71.676
R835 B.n199 B.n84 71.676
R836 B.n203 B.n85 71.676
R837 B.n208 B.n86 71.676
R838 B.n212 B.n87 71.676
R839 B.n216 B.n88 71.676
R840 B.n220 B.n89 71.676
R841 B.n224 B.n90 71.676
R842 B.n229 B.n91 71.676
R843 B.n233 B.n92 71.676
R844 B.n237 B.n93 71.676
R845 B.n241 B.n94 71.676
R846 B.n245 B.n95 71.676
R847 B.n249 B.n96 71.676
R848 B.n253 B.n97 71.676
R849 B.n257 B.n98 71.676
R850 B.n261 B.n99 71.676
R851 B.n265 B.n100 71.676
R852 B.n269 B.n101 71.676
R853 B.n273 B.n102 71.676
R854 B.n277 B.n103 71.676
R855 B.n281 B.n104 71.676
R856 B.n285 B.n105 71.676
R857 B.n289 B.n106 71.676
R858 B.n293 B.n107 71.676
R859 B.n297 B.n108 71.676
R860 B.n301 B.n109 71.676
R861 B.n305 B.n110 71.676
R862 B.n309 B.n111 71.676
R863 B.n772 B.n112 71.676
R864 B.n772 B.n771 71.676
R865 B.n311 B.n111 71.676
R866 B.n308 B.n110 71.676
R867 B.n304 B.n109 71.676
R868 B.n300 B.n108 71.676
R869 B.n296 B.n107 71.676
R870 B.n292 B.n106 71.676
R871 B.n288 B.n105 71.676
R872 B.n284 B.n104 71.676
R873 B.n280 B.n103 71.676
R874 B.n276 B.n102 71.676
R875 B.n272 B.n101 71.676
R876 B.n268 B.n100 71.676
R877 B.n264 B.n99 71.676
R878 B.n260 B.n98 71.676
R879 B.n256 B.n97 71.676
R880 B.n252 B.n96 71.676
R881 B.n248 B.n95 71.676
R882 B.n244 B.n94 71.676
R883 B.n240 B.n93 71.676
R884 B.n236 B.n92 71.676
R885 B.n232 B.n91 71.676
R886 B.n228 B.n90 71.676
R887 B.n223 B.n89 71.676
R888 B.n219 B.n88 71.676
R889 B.n215 B.n87 71.676
R890 B.n211 B.n86 71.676
R891 B.n207 B.n85 71.676
R892 B.n202 B.n84 71.676
R893 B.n198 B.n83 71.676
R894 B.n194 B.n82 71.676
R895 B.n190 B.n81 71.676
R896 B.n186 B.n80 71.676
R897 B.n182 B.n79 71.676
R898 B.n178 B.n78 71.676
R899 B.n174 B.n77 71.676
R900 B.n170 B.n76 71.676
R901 B.n166 B.n75 71.676
R902 B.n162 B.n74 71.676
R903 B.n158 B.n73 71.676
R904 B.n154 B.n72 71.676
R905 B.n150 B.n71 71.676
R906 B.n146 B.n70 71.676
R907 B.n142 B.n69 71.676
R908 B.n138 B.n68 71.676
R909 B.n134 B.n67 71.676
R910 B.n130 B.n66 71.676
R911 B.n126 B.n65 71.676
R912 B.n122 B.n64 71.676
R913 B.n118 B.n63 71.676
R914 B.n431 B.n374 71.676
R915 B.n437 B.n436 71.676
R916 B.n440 B.n439 71.676
R917 B.n445 B.n444 71.676
R918 B.n448 B.n447 71.676
R919 B.n453 B.n452 71.676
R920 B.n456 B.n455 71.676
R921 B.n461 B.n460 71.676
R922 B.n464 B.n463 71.676
R923 B.n469 B.n468 71.676
R924 B.n472 B.n471 71.676
R925 B.n477 B.n476 71.676
R926 B.n480 B.n479 71.676
R927 B.n485 B.n484 71.676
R928 B.n488 B.n487 71.676
R929 B.n493 B.n492 71.676
R930 B.n496 B.n495 71.676
R931 B.n501 B.n500 71.676
R932 B.n504 B.n503 71.676
R933 B.n509 B.n508 71.676
R934 B.n512 B.n511 71.676
R935 B.n517 B.n516 71.676
R936 B.n520 B.n519 71.676
R937 B.n525 B.n524 71.676
R938 B.n528 B.n527 71.676
R939 B.n533 B.n532 71.676
R940 B.n536 B.n535 71.676
R941 B.n542 B.n541 71.676
R942 B.n545 B.n544 71.676
R943 B.n550 B.n549 71.676
R944 B.n553 B.n552 71.676
R945 B.n558 B.n557 71.676
R946 B.n561 B.n560 71.676
R947 B.n566 B.n565 71.676
R948 B.n569 B.n568 71.676
R949 B.n574 B.n573 71.676
R950 B.n577 B.n576 71.676
R951 B.n582 B.n581 71.676
R952 B.n585 B.n584 71.676
R953 B.n590 B.n589 71.676
R954 B.n593 B.n592 71.676
R955 B.n598 B.n597 71.676
R956 B.n601 B.n600 71.676
R957 B.n606 B.n605 71.676
R958 B.n609 B.n608 71.676
R959 B.n614 B.n613 71.676
R960 B.n617 B.n616 71.676
R961 B.n622 B.n621 71.676
R962 B.n625 B.n624 71.676
R963 B.n432 B.n431 71.676
R964 B.n438 B.n437 71.676
R965 B.n439 B.n428 71.676
R966 B.n446 B.n445 71.676
R967 B.n447 B.n426 71.676
R968 B.n454 B.n453 71.676
R969 B.n455 B.n424 71.676
R970 B.n462 B.n461 71.676
R971 B.n463 B.n422 71.676
R972 B.n470 B.n469 71.676
R973 B.n471 B.n420 71.676
R974 B.n478 B.n477 71.676
R975 B.n479 B.n418 71.676
R976 B.n486 B.n485 71.676
R977 B.n487 B.n416 71.676
R978 B.n494 B.n493 71.676
R979 B.n495 B.n414 71.676
R980 B.n502 B.n501 71.676
R981 B.n503 B.n412 71.676
R982 B.n510 B.n509 71.676
R983 B.n511 B.n410 71.676
R984 B.n518 B.n517 71.676
R985 B.n519 B.n405 71.676
R986 B.n526 B.n525 71.676
R987 B.n527 B.n403 71.676
R988 B.n534 B.n533 71.676
R989 B.n535 B.n399 71.676
R990 B.n543 B.n542 71.676
R991 B.n544 B.n397 71.676
R992 B.n551 B.n550 71.676
R993 B.n552 B.n395 71.676
R994 B.n559 B.n558 71.676
R995 B.n560 B.n393 71.676
R996 B.n567 B.n566 71.676
R997 B.n568 B.n391 71.676
R998 B.n575 B.n574 71.676
R999 B.n576 B.n389 71.676
R1000 B.n583 B.n582 71.676
R1001 B.n584 B.n387 71.676
R1002 B.n591 B.n590 71.676
R1003 B.n592 B.n385 71.676
R1004 B.n599 B.n598 71.676
R1005 B.n600 B.n383 71.676
R1006 B.n607 B.n606 71.676
R1007 B.n608 B.n381 71.676
R1008 B.n615 B.n614 71.676
R1009 B.n616 B.n379 71.676
R1010 B.n623 B.n622 71.676
R1011 B.n626 B.n625 71.676
R1012 B.n841 B.n840 71.676
R1013 B.n841 B.n2 71.676
R1014 B.n205 B.n116 59.5399
R1015 B.n226 B.n114 59.5399
R1016 B.n539 B.n401 59.5399
R1017 B.n408 B.n407 59.5399
R1018 B.n631 B.n371 40.2914
R1019 B.n637 B.n371 40.2914
R1020 B.n637 B.n367 40.2914
R1021 B.n643 B.n367 40.2914
R1022 B.n643 B.n363 40.2914
R1023 B.n649 B.n363 40.2914
R1024 B.n649 B.n359 40.2914
R1025 B.n656 B.n359 40.2914
R1026 B.n656 B.n655 40.2914
R1027 B.n662 B.n352 40.2914
R1028 B.n668 B.n352 40.2914
R1029 B.n668 B.n348 40.2914
R1030 B.n674 B.n348 40.2914
R1031 B.n674 B.n344 40.2914
R1032 B.n680 B.n344 40.2914
R1033 B.n680 B.n340 40.2914
R1034 B.n686 B.n340 40.2914
R1035 B.n686 B.n336 40.2914
R1036 B.n692 B.n336 40.2914
R1037 B.n692 B.n332 40.2914
R1038 B.n698 B.n332 40.2914
R1039 B.n698 B.n328 40.2914
R1040 B.n704 B.n328 40.2914
R1041 B.n710 B.n324 40.2914
R1042 B.n710 B.n320 40.2914
R1043 B.n717 B.n320 40.2914
R1044 B.n717 B.n316 40.2914
R1045 B.n723 B.n316 40.2914
R1046 B.n723 B.n4 40.2914
R1047 B.n839 B.n4 40.2914
R1048 B.n839 B.n838 40.2914
R1049 B.n838 B.n837 40.2914
R1050 B.n837 B.n8 40.2914
R1051 B.n12 B.n8 40.2914
R1052 B.n830 B.n12 40.2914
R1053 B.n830 B.n829 40.2914
R1054 B.n829 B.n828 40.2914
R1055 B.n828 B.n16 40.2914
R1056 B.n822 B.n821 40.2914
R1057 B.n821 B.n820 40.2914
R1058 B.n820 B.n23 40.2914
R1059 B.n814 B.n23 40.2914
R1060 B.n814 B.n813 40.2914
R1061 B.n813 B.n812 40.2914
R1062 B.n812 B.n30 40.2914
R1063 B.n806 B.n30 40.2914
R1064 B.n806 B.n805 40.2914
R1065 B.n805 B.n804 40.2914
R1066 B.n804 B.n37 40.2914
R1067 B.n798 B.n37 40.2914
R1068 B.n798 B.n797 40.2914
R1069 B.n797 B.n796 40.2914
R1070 B.n790 B.n47 40.2914
R1071 B.n790 B.n789 40.2914
R1072 B.n789 B.n788 40.2914
R1073 B.n788 B.n51 40.2914
R1074 B.n782 B.n51 40.2914
R1075 B.n782 B.n781 40.2914
R1076 B.n781 B.n780 40.2914
R1077 B.n780 B.n58 40.2914
R1078 B.n774 B.n58 40.2914
R1079 B.n633 B.n373 34.8103
R1080 B.n629 B.n628 34.8103
R1081 B.n770 B.n769 34.8103
R1082 B.n776 B.n60 34.8103
R1083 B.n704 B.t0 31.9962
R1084 B.n822 B.t1 31.9962
R1085 B.n662 B.t3 24.886
R1086 B.n796 B.t7 24.886
R1087 B B.n842 18.0485
R1088 B.n655 B.t3 15.4058
R1089 B.n47 B.t7 15.4058
R1090 B.n634 B.n633 10.6151
R1091 B.n635 B.n634 10.6151
R1092 B.n635 B.n365 10.6151
R1093 B.n645 B.n365 10.6151
R1094 B.n646 B.n645 10.6151
R1095 B.n647 B.n646 10.6151
R1096 B.n647 B.n357 10.6151
R1097 B.n658 B.n357 10.6151
R1098 B.n659 B.n658 10.6151
R1099 B.n660 B.n659 10.6151
R1100 B.n660 B.n350 10.6151
R1101 B.n670 B.n350 10.6151
R1102 B.n671 B.n670 10.6151
R1103 B.n672 B.n671 10.6151
R1104 B.n672 B.n342 10.6151
R1105 B.n682 B.n342 10.6151
R1106 B.n683 B.n682 10.6151
R1107 B.n684 B.n683 10.6151
R1108 B.n684 B.n334 10.6151
R1109 B.n694 B.n334 10.6151
R1110 B.n695 B.n694 10.6151
R1111 B.n696 B.n695 10.6151
R1112 B.n696 B.n326 10.6151
R1113 B.n706 B.n326 10.6151
R1114 B.n707 B.n706 10.6151
R1115 B.n708 B.n707 10.6151
R1116 B.n708 B.n318 10.6151
R1117 B.n719 B.n318 10.6151
R1118 B.n720 B.n719 10.6151
R1119 B.n721 B.n720 10.6151
R1120 B.n721 B.n0 10.6151
R1121 B.n433 B.n373 10.6151
R1122 B.n434 B.n433 10.6151
R1123 B.n435 B.n434 10.6151
R1124 B.n435 B.n429 10.6151
R1125 B.n441 B.n429 10.6151
R1126 B.n442 B.n441 10.6151
R1127 B.n443 B.n442 10.6151
R1128 B.n443 B.n427 10.6151
R1129 B.n449 B.n427 10.6151
R1130 B.n450 B.n449 10.6151
R1131 B.n451 B.n450 10.6151
R1132 B.n451 B.n425 10.6151
R1133 B.n457 B.n425 10.6151
R1134 B.n458 B.n457 10.6151
R1135 B.n459 B.n458 10.6151
R1136 B.n459 B.n423 10.6151
R1137 B.n465 B.n423 10.6151
R1138 B.n466 B.n465 10.6151
R1139 B.n467 B.n466 10.6151
R1140 B.n467 B.n421 10.6151
R1141 B.n473 B.n421 10.6151
R1142 B.n474 B.n473 10.6151
R1143 B.n475 B.n474 10.6151
R1144 B.n475 B.n419 10.6151
R1145 B.n481 B.n419 10.6151
R1146 B.n482 B.n481 10.6151
R1147 B.n483 B.n482 10.6151
R1148 B.n483 B.n417 10.6151
R1149 B.n489 B.n417 10.6151
R1150 B.n490 B.n489 10.6151
R1151 B.n491 B.n490 10.6151
R1152 B.n491 B.n415 10.6151
R1153 B.n497 B.n415 10.6151
R1154 B.n498 B.n497 10.6151
R1155 B.n499 B.n498 10.6151
R1156 B.n499 B.n413 10.6151
R1157 B.n505 B.n413 10.6151
R1158 B.n506 B.n505 10.6151
R1159 B.n507 B.n506 10.6151
R1160 B.n507 B.n411 10.6151
R1161 B.n513 B.n411 10.6151
R1162 B.n514 B.n513 10.6151
R1163 B.n515 B.n514 10.6151
R1164 B.n515 B.n409 10.6151
R1165 B.n522 B.n521 10.6151
R1166 B.n523 B.n522 10.6151
R1167 B.n523 B.n404 10.6151
R1168 B.n529 B.n404 10.6151
R1169 B.n530 B.n529 10.6151
R1170 B.n531 B.n530 10.6151
R1171 B.n531 B.n402 10.6151
R1172 B.n537 B.n402 10.6151
R1173 B.n538 B.n537 10.6151
R1174 B.n540 B.n398 10.6151
R1175 B.n546 B.n398 10.6151
R1176 B.n547 B.n546 10.6151
R1177 B.n548 B.n547 10.6151
R1178 B.n548 B.n396 10.6151
R1179 B.n554 B.n396 10.6151
R1180 B.n555 B.n554 10.6151
R1181 B.n556 B.n555 10.6151
R1182 B.n556 B.n394 10.6151
R1183 B.n562 B.n394 10.6151
R1184 B.n563 B.n562 10.6151
R1185 B.n564 B.n563 10.6151
R1186 B.n564 B.n392 10.6151
R1187 B.n570 B.n392 10.6151
R1188 B.n571 B.n570 10.6151
R1189 B.n572 B.n571 10.6151
R1190 B.n572 B.n390 10.6151
R1191 B.n578 B.n390 10.6151
R1192 B.n579 B.n578 10.6151
R1193 B.n580 B.n579 10.6151
R1194 B.n580 B.n388 10.6151
R1195 B.n586 B.n388 10.6151
R1196 B.n587 B.n586 10.6151
R1197 B.n588 B.n587 10.6151
R1198 B.n588 B.n386 10.6151
R1199 B.n594 B.n386 10.6151
R1200 B.n595 B.n594 10.6151
R1201 B.n596 B.n595 10.6151
R1202 B.n596 B.n384 10.6151
R1203 B.n602 B.n384 10.6151
R1204 B.n603 B.n602 10.6151
R1205 B.n604 B.n603 10.6151
R1206 B.n604 B.n382 10.6151
R1207 B.n610 B.n382 10.6151
R1208 B.n611 B.n610 10.6151
R1209 B.n612 B.n611 10.6151
R1210 B.n612 B.n380 10.6151
R1211 B.n618 B.n380 10.6151
R1212 B.n619 B.n618 10.6151
R1213 B.n620 B.n619 10.6151
R1214 B.n620 B.n378 10.6151
R1215 B.n378 B.n377 10.6151
R1216 B.n627 B.n377 10.6151
R1217 B.n628 B.n627 10.6151
R1218 B.n629 B.n369 10.6151
R1219 B.n639 B.n369 10.6151
R1220 B.n640 B.n639 10.6151
R1221 B.n641 B.n640 10.6151
R1222 B.n641 B.n361 10.6151
R1223 B.n651 B.n361 10.6151
R1224 B.n652 B.n651 10.6151
R1225 B.n653 B.n652 10.6151
R1226 B.n653 B.n354 10.6151
R1227 B.n664 B.n354 10.6151
R1228 B.n665 B.n664 10.6151
R1229 B.n666 B.n665 10.6151
R1230 B.n666 B.n346 10.6151
R1231 B.n676 B.n346 10.6151
R1232 B.n677 B.n676 10.6151
R1233 B.n678 B.n677 10.6151
R1234 B.n678 B.n338 10.6151
R1235 B.n688 B.n338 10.6151
R1236 B.n689 B.n688 10.6151
R1237 B.n690 B.n689 10.6151
R1238 B.n690 B.n330 10.6151
R1239 B.n700 B.n330 10.6151
R1240 B.n701 B.n700 10.6151
R1241 B.n702 B.n701 10.6151
R1242 B.n702 B.n322 10.6151
R1243 B.n712 B.n322 10.6151
R1244 B.n713 B.n712 10.6151
R1245 B.n715 B.n713 10.6151
R1246 B.n715 B.n714 10.6151
R1247 B.n714 B.n314 10.6151
R1248 B.n726 B.n314 10.6151
R1249 B.n727 B.n726 10.6151
R1250 B.n728 B.n727 10.6151
R1251 B.n729 B.n728 10.6151
R1252 B.n730 B.n729 10.6151
R1253 B.n733 B.n730 10.6151
R1254 B.n734 B.n733 10.6151
R1255 B.n735 B.n734 10.6151
R1256 B.n736 B.n735 10.6151
R1257 B.n738 B.n736 10.6151
R1258 B.n739 B.n738 10.6151
R1259 B.n740 B.n739 10.6151
R1260 B.n741 B.n740 10.6151
R1261 B.n743 B.n741 10.6151
R1262 B.n744 B.n743 10.6151
R1263 B.n745 B.n744 10.6151
R1264 B.n746 B.n745 10.6151
R1265 B.n748 B.n746 10.6151
R1266 B.n749 B.n748 10.6151
R1267 B.n750 B.n749 10.6151
R1268 B.n751 B.n750 10.6151
R1269 B.n753 B.n751 10.6151
R1270 B.n754 B.n753 10.6151
R1271 B.n755 B.n754 10.6151
R1272 B.n756 B.n755 10.6151
R1273 B.n758 B.n756 10.6151
R1274 B.n759 B.n758 10.6151
R1275 B.n760 B.n759 10.6151
R1276 B.n761 B.n760 10.6151
R1277 B.n763 B.n761 10.6151
R1278 B.n764 B.n763 10.6151
R1279 B.n765 B.n764 10.6151
R1280 B.n766 B.n765 10.6151
R1281 B.n768 B.n766 10.6151
R1282 B.n769 B.n768 10.6151
R1283 B.n834 B.n1 10.6151
R1284 B.n834 B.n833 10.6151
R1285 B.n833 B.n832 10.6151
R1286 B.n832 B.n10 10.6151
R1287 B.n826 B.n10 10.6151
R1288 B.n826 B.n825 10.6151
R1289 B.n825 B.n824 10.6151
R1290 B.n824 B.n18 10.6151
R1291 B.n818 B.n18 10.6151
R1292 B.n818 B.n817 10.6151
R1293 B.n817 B.n816 10.6151
R1294 B.n816 B.n25 10.6151
R1295 B.n810 B.n25 10.6151
R1296 B.n810 B.n809 10.6151
R1297 B.n809 B.n808 10.6151
R1298 B.n808 B.n32 10.6151
R1299 B.n802 B.n32 10.6151
R1300 B.n802 B.n801 10.6151
R1301 B.n801 B.n800 10.6151
R1302 B.n800 B.n39 10.6151
R1303 B.n794 B.n39 10.6151
R1304 B.n794 B.n793 10.6151
R1305 B.n793 B.n792 10.6151
R1306 B.n792 B.n45 10.6151
R1307 B.n786 B.n45 10.6151
R1308 B.n786 B.n785 10.6151
R1309 B.n785 B.n784 10.6151
R1310 B.n784 B.n53 10.6151
R1311 B.n778 B.n53 10.6151
R1312 B.n778 B.n777 10.6151
R1313 B.n777 B.n776 10.6151
R1314 B.n117 B.n60 10.6151
R1315 B.n120 B.n117 10.6151
R1316 B.n121 B.n120 10.6151
R1317 B.n124 B.n121 10.6151
R1318 B.n125 B.n124 10.6151
R1319 B.n128 B.n125 10.6151
R1320 B.n129 B.n128 10.6151
R1321 B.n132 B.n129 10.6151
R1322 B.n133 B.n132 10.6151
R1323 B.n136 B.n133 10.6151
R1324 B.n137 B.n136 10.6151
R1325 B.n140 B.n137 10.6151
R1326 B.n141 B.n140 10.6151
R1327 B.n144 B.n141 10.6151
R1328 B.n145 B.n144 10.6151
R1329 B.n148 B.n145 10.6151
R1330 B.n149 B.n148 10.6151
R1331 B.n152 B.n149 10.6151
R1332 B.n153 B.n152 10.6151
R1333 B.n156 B.n153 10.6151
R1334 B.n157 B.n156 10.6151
R1335 B.n160 B.n157 10.6151
R1336 B.n161 B.n160 10.6151
R1337 B.n164 B.n161 10.6151
R1338 B.n165 B.n164 10.6151
R1339 B.n168 B.n165 10.6151
R1340 B.n169 B.n168 10.6151
R1341 B.n172 B.n169 10.6151
R1342 B.n173 B.n172 10.6151
R1343 B.n176 B.n173 10.6151
R1344 B.n177 B.n176 10.6151
R1345 B.n180 B.n177 10.6151
R1346 B.n181 B.n180 10.6151
R1347 B.n184 B.n181 10.6151
R1348 B.n185 B.n184 10.6151
R1349 B.n188 B.n185 10.6151
R1350 B.n189 B.n188 10.6151
R1351 B.n192 B.n189 10.6151
R1352 B.n193 B.n192 10.6151
R1353 B.n196 B.n193 10.6151
R1354 B.n197 B.n196 10.6151
R1355 B.n200 B.n197 10.6151
R1356 B.n201 B.n200 10.6151
R1357 B.n204 B.n201 10.6151
R1358 B.n209 B.n206 10.6151
R1359 B.n210 B.n209 10.6151
R1360 B.n213 B.n210 10.6151
R1361 B.n214 B.n213 10.6151
R1362 B.n217 B.n214 10.6151
R1363 B.n218 B.n217 10.6151
R1364 B.n221 B.n218 10.6151
R1365 B.n222 B.n221 10.6151
R1366 B.n225 B.n222 10.6151
R1367 B.n230 B.n227 10.6151
R1368 B.n231 B.n230 10.6151
R1369 B.n234 B.n231 10.6151
R1370 B.n235 B.n234 10.6151
R1371 B.n238 B.n235 10.6151
R1372 B.n239 B.n238 10.6151
R1373 B.n242 B.n239 10.6151
R1374 B.n243 B.n242 10.6151
R1375 B.n246 B.n243 10.6151
R1376 B.n247 B.n246 10.6151
R1377 B.n250 B.n247 10.6151
R1378 B.n251 B.n250 10.6151
R1379 B.n254 B.n251 10.6151
R1380 B.n255 B.n254 10.6151
R1381 B.n258 B.n255 10.6151
R1382 B.n259 B.n258 10.6151
R1383 B.n262 B.n259 10.6151
R1384 B.n263 B.n262 10.6151
R1385 B.n266 B.n263 10.6151
R1386 B.n267 B.n266 10.6151
R1387 B.n270 B.n267 10.6151
R1388 B.n271 B.n270 10.6151
R1389 B.n274 B.n271 10.6151
R1390 B.n275 B.n274 10.6151
R1391 B.n278 B.n275 10.6151
R1392 B.n279 B.n278 10.6151
R1393 B.n282 B.n279 10.6151
R1394 B.n283 B.n282 10.6151
R1395 B.n286 B.n283 10.6151
R1396 B.n287 B.n286 10.6151
R1397 B.n290 B.n287 10.6151
R1398 B.n291 B.n290 10.6151
R1399 B.n294 B.n291 10.6151
R1400 B.n295 B.n294 10.6151
R1401 B.n298 B.n295 10.6151
R1402 B.n299 B.n298 10.6151
R1403 B.n302 B.n299 10.6151
R1404 B.n303 B.n302 10.6151
R1405 B.n306 B.n303 10.6151
R1406 B.n307 B.n306 10.6151
R1407 B.n310 B.n307 10.6151
R1408 B.n312 B.n310 10.6151
R1409 B.n313 B.n312 10.6151
R1410 B.n770 B.n313 10.6151
R1411 B.n409 B.n408 9.36635
R1412 B.n540 B.n539 9.36635
R1413 B.n205 B.n204 9.36635
R1414 B.n227 B.n226 9.36635
R1415 B.t0 B.n324 8.29568
R1416 B.t1 B.n16 8.29568
R1417 B.n842 B.n0 8.11757
R1418 B.n842 B.n1 8.11757
R1419 B.n521 B.n408 1.24928
R1420 B.n539 B.n538 1.24928
R1421 B.n206 B.n205 1.24928
R1422 B.n226 B.n225 1.24928
R1423 VP.n0 VP.t1 167.751
R1424 VP.n0 VP.t0 118.882
R1425 VP VP.n0 0.621237
R1426 VTAIL.n282 VTAIL.n216 214.453
R1427 VTAIL.n66 VTAIL.n0 214.453
R1428 VTAIL.n210 VTAIL.n144 214.453
R1429 VTAIL.n138 VTAIL.n72 214.453
R1430 VTAIL.n241 VTAIL.n240 185
R1431 VTAIL.n243 VTAIL.n242 185
R1432 VTAIL.n236 VTAIL.n235 185
R1433 VTAIL.n249 VTAIL.n248 185
R1434 VTAIL.n251 VTAIL.n250 185
R1435 VTAIL.n232 VTAIL.n231 185
R1436 VTAIL.n257 VTAIL.n256 185
R1437 VTAIL.n259 VTAIL.n258 185
R1438 VTAIL.n228 VTAIL.n227 185
R1439 VTAIL.n265 VTAIL.n264 185
R1440 VTAIL.n267 VTAIL.n266 185
R1441 VTAIL.n224 VTAIL.n223 185
R1442 VTAIL.n273 VTAIL.n272 185
R1443 VTAIL.n275 VTAIL.n274 185
R1444 VTAIL.n220 VTAIL.n219 185
R1445 VTAIL.n281 VTAIL.n280 185
R1446 VTAIL.n283 VTAIL.n282 185
R1447 VTAIL.n25 VTAIL.n24 185
R1448 VTAIL.n27 VTAIL.n26 185
R1449 VTAIL.n20 VTAIL.n19 185
R1450 VTAIL.n33 VTAIL.n32 185
R1451 VTAIL.n35 VTAIL.n34 185
R1452 VTAIL.n16 VTAIL.n15 185
R1453 VTAIL.n41 VTAIL.n40 185
R1454 VTAIL.n43 VTAIL.n42 185
R1455 VTAIL.n12 VTAIL.n11 185
R1456 VTAIL.n49 VTAIL.n48 185
R1457 VTAIL.n51 VTAIL.n50 185
R1458 VTAIL.n8 VTAIL.n7 185
R1459 VTAIL.n57 VTAIL.n56 185
R1460 VTAIL.n59 VTAIL.n58 185
R1461 VTAIL.n4 VTAIL.n3 185
R1462 VTAIL.n65 VTAIL.n64 185
R1463 VTAIL.n67 VTAIL.n66 185
R1464 VTAIL.n211 VTAIL.n210 185
R1465 VTAIL.n209 VTAIL.n208 185
R1466 VTAIL.n148 VTAIL.n147 185
R1467 VTAIL.n203 VTAIL.n202 185
R1468 VTAIL.n201 VTAIL.n200 185
R1469 VTAIL.n152 VTAIL.n151 185
R1470 VTAIL.n195 VTAIL.n194 185
R1471 VTAIL.n193 VTAIL.n192 185
R1472 VTAIL.n156 VTAIL.n155 185
R1473 VTAIL.n187 VTAIL.n186 185
R1474 VTAIL.n185 VTAIL.n184 185
R1475 VTAIL.n160 VTAIL.n159 185
R1476 VTAIL.n179 VTAIL.n178 185
R1477 VTAIL.n177 VTAIL.n176 185
R1478 VTAIL.n164 VTAIL.n163 185
R1479 VTAIL.n171 VTAIL.n170 185
R1480 VTAIL.n169 VTAIL.n168 185
R1481 VTAIL.n139 VTAIL.n138 185
R1482 VTAIL.n137 VTAIL.n136 185
R1483 VTAIL.n76 VTAIL.n75 185
R1484 VTAIL.n131 VTAIL.n130 185
R1485 VTAIL.n129 VTAIL.n128 185
R1486 VTAIL.n80 VTAIL.n79 185
R1487 VTAIL.n123 VTAIL.n122 185
R1488 VTAIL.n121 VTAIL.n120 185
R1489 VTAIL.n84 VTAIL.n83 185
R1490 VTAIL.n115 VTAIL.n114 185
R1491 VTAIL.n113 VTAIL.n112 185
R1492 VTAIL.n88 VTAIL.n87 185
R1493 VTAIL.n107 VTAIL.n106 185
R1494 VTAIL.n105 VTAIL.n104 185
R1495 VTAIL.n92 VTAIL.n91 185
R1496 VTAIL.n99 VTAIL.n98 185
R1497 VTAIL.n97 VTAIL.n96 185
R1498 VTAIL.n239 VTAIL.t1 147.659
R1499 VTAIL.n23 VTAIL.t3 147.659
R1500 VTAIL.n167 VTAIL.t2 147.659
R1501 VTAIL.n95 VTAIL.t0 147.659
R1502 VTAIL.n242 VTAIL.n241 104.615
R1503 VTAIL.n242 VTAIL.n235 104.615
R1504 VTAIL.n249 VTAIL.n235 104.615
R1505 VTAIL.n250 VTAIL.n249 104.615
R1506 VTAIL.n250 VTAIL.n231 104.615
R1507 VTAIL.n257 VTAIL.n231 104.615
R1508 VTAIL.n258 VTAIL.n257 104.615
R1509 VTAIL.n258 VTAIL.n227 104.615
R1510 VTAIL.n265 VTAIL.n227 104.615
R1511 VTAIL.n266 VTAIL.n265 104.615
R1512 VTAIL.n266 VTAIL.n223 104.615
R1513 VTAIL.n273 VTAIL.n223 104.615
R1514 VTAIL.n274 VTAIL.n273 104.615
R1515 VTAIL.n274 VTAIL.n219 104.615
R1516 VTAIL.n281 VTAIL.n219 104.615
R1517 VTAIL.n282 VTAIL.n281 104.615
R1518 VTAIL.n26 VTAIL.n25 104.615
R1519 VTAIL.n26 VTAIL.n19 104.615
R1520 VTAIL.n33 VTAIL.n19 104.615
R1521 VTAIL.n34 VTAIL.n33 104.615
R1522 VTAIL.n34 VTAIL.n15 104.615
R1523 VTAIL.n41 VTAIL.n15 104.615
R1524 VTAIL.n42 VTAIL.n41 104.615
R1525 VTAIL.n42 VTAIL.n11 104.615
R1526 VTAIL.n49 VTAIL.n11 104.615
R1527 VTAIL.n50 VTAIL.n49 104.615
R1528 VTAIL.n50 VTAIL.n7 104.615
R1529 VTAIL.n57 VTAIL.n7 104.615
R1530 VTAIL.n58 VTAIL.n57 104.615
R1531 VTAIL.n58 VTAIL.n3 104.615
R1532 VTAIL.n65 VTAIL.n3 104.615
R1533 VTAIL.n66 VTAIL.n65 104.615
R1534 VTAIL.n210 VTAIL.n209 104.615
R1535 VTAIL.n209 VTAIL.n147 104.615
R1536 VTAIL.n202 VTAIL.n147 104.615
R1537 VTAIL.n202 VTAIL.n201 104.615
R1538 VTAIL.n201 VTAIL.n151 104.615
R1539 VTAIL.n194 VTAIL.n151 104.615
R1540 VTAIL.n194 VTAIL.n193 104.615
R1541 VTAIL.n193 VTAIL.n155 104.615
R1542 VTAIL.n186 VTAIL.n155 104.615
R1543 VTAIL.n186 VTAIL.n185 104.615
R1544 VTAIL.n185 VTAIL.n159 104.615
R1545 VTAIL.n178 VTAIL.n159 104.615
R1546 VTAIL.n178 VTAIL.n177 104.615
R1547 VTAIL.n177 VTAIL.n163 104.615
R1548 VTAIL.n170 VTAIL.n163 104.615
R1549 VTAIL.n170 VTAIL.n169 104.615
R1550 VTAIL.n138 VTAIL.n137 104.615
R1551 VTAIL.n137 VTAIL.n75 104.615
R1552 VTAIL.n130 VTAIL.n75 104.615
R1553 VTAIL.n130 VTAIL.n129 104.615
R1554 VTAIL.n129 VTAIL.n79 104.615
R1555 VTAIL.n122 VTAIL.n79 104.615
R1556 VTAIL.n122 VTAIL.n121 104.615
R1557 VTAIL.n121 VTAIL.n83 104.615
R1558 VTAIL.n114 VTAIL.n83 104.615
R1559 VTAIL.n114 VTAIL.n113 104.615
R1560 VTAIL.n113 VTAIL.n87 104.615
R1561 VTAIL.n106 VTAIL.n87 104.615
R1562 VTAIL.n106 VTAIL.n105 104.615
R1563 VTAIL.n105 VTAIL.n91 104.615
R1564 VTAIL.n98 VTAIL.n91 104.615
R1565 VTAIL.n98 VTAIL.n97 104.615
R1566 VTAIL.n241 VTAIL.t1 52.3082
R1567 VTAIL.n25 VTAIL.t3 52.3082
R1568 VTAIL.n169 VTAIL.t2 52.3082
R1569 VTAIL.n97 VTAIL.t0 52.3082
R1570 VTAIL.n287 VTAIL.n286 33.9308
R1571 VTAIL.n71 VTAIL.n70 33.9308
R1572 VTAIL.n215 VTAIL.n214 33.9308
R1573 VTAIL.n143 VTAIL.n142 33.9308
R1574 VTAIL.n143 VTAIL.n71 30.9789
R1575 VTAIL.n287 VTAIL.n215 27.4014
R1576 VTAIL.n240 VTAIL.n239 15.6677
R1577 VTAIL.n24 VTAIL.n23 15.6677
R1578 VTAIL.n168 VTAIL.n167 15.6677
R1579 VTAIL.n96 VTAIL.n95 15.6677
R1580 VTAIL.n243 VTAIL.n238 12.8005
R1581 VTAIL.n284 VTAIL.n283 12.8005
R1582 VTAIL.n27 VTAIL.n22 12.8005
R1583 VTAIL.n68 VTAIL.n67 12.8005
R1584 VTAIL.n212 VTAIL.n211 12.8005
R1585 VTAIL.n171 VTAIL.n166 12.8005
R1586 VTAIL.n140 VTAIL.n139 12.8005
R1587 VTAIL.n99 VTAIL.n94 12.8005
R1588 VTAIL.n244 VTAIL.n236 12.0247
R1589 VTAIL.n280 VTAIL.n218 12.0247
R1590 VTAIL.n28 VTAIL.n20 12.0247
R1591 VTAIL.n64 VTAIL.n2 12.0247
R1592 VTAIL.n208 VTAIL.n146 12.0247
R1593 VTAIL.n172 VTAIL.n164 12.0247
R1594 VTAIL.n136 VTAIL.n74 12.0247
R1595 VTAIL.n100 VTAIL.n92 12.0247
R1596 VTAIL.n248 VTAIL.n247 11.249
R1597 VTAIL.n279 VTAIL.n220 11.249
R1598 VTAIL.n32 VTAIL.n31 11.249
R1599 VTAIL.n63 VTAIL.n4 11.249
R1600 VTAIL.n207 VTAIL.n148 11.249
R1601 VTAIL.n176 VTAIL.n175 11.249
R1602 VTAIL.n135 VTAIL.n76 11.249
R1603 VTAIL.n104 VTAIL.n103 11.249
R1604 VTAIL.n251 VTAIL.n234 10.4732
R1605 VTAIL.n276 VTAIL.n275 10.4732
R1606 VTAIL.n35 VTAIL.n18 10.4732
R1607 VTAIL.n60 VTAIL.n59 10.4732
R1608 VTAIL.n204 VTAIL.n203 10.4732
R1609 VTAIL.n179 VTAIL.n162 10.4732
R1610 VTAIL.n132 VTAIL.n131 10.4732
R1611 VTAIL.n107 VTAIL.n90 10.4732
R1612 VTAIL.n252 VTAIL.n232 9.69747
R1613 VTAIL.n272 VTAIL.n222 9.69747
R1614 VTAIL.n36 VTAIL.n16 9.69747
R1615 VTAIL.n56 VTAIL.n6 9.69747
R1616 VTAIL.n200 VTAIL.n150 9.69747
R1617 VTAIL.n180 VTAIL.n160 9.69747
R1618 VTAIL.n128 VTAIL.n78 9.69747
R1619 VTAIL.n108 VTAIL.n88 9.69747
R1620 VTAIL.n286 VTAIL.n285 9.45567
R1621 VTAIL.n70 VTAIL.n69 9.45567
R1622 VTAIL.n214 VTAIL.n213 9.45567
R1623 VTAIL.n142 VTAIL.n141 9.45567
R1624 VTAIL.n261 VTAIL.n260 9.3005
R1625 VTAIL.n230 VTAIL.n229 9.3005
R1626 VTAIL.n255 VTAIL.n254 9.3005
R1627 VTAIL.n253 VTAIL.n252 9.3005
R1628 VTAIL.n234 VTAIL.n233 9.3005
R1629 VTAIL.n247 VTAIL.n246 9.3005
R1630 VTAIL.n245 VTAIL.n244 9.3005
R1631 VTAIL.n238 VTAIL.n237 9.3005
R1632 VTAIL.n263 VTAIL.n262 9.3005
R1633 VTAIL.n226 VTAIL.n225 9.3005
R1634 VTAIL.n269 VTAIL.n268 9.3005
R1635 VTAIL.n271 VTAIL.n270 9.3005
R1636 VTAIL.n222 VTAIL.n221 9.3005
R1637 VTAIL.n277 VTAIL.n276 9.3005
R1638 VTAIL.n279 VTAIL.n278 9.3005
R1639 VTAIL.n218 VTAIL.n217 9.3005
R1640 VTAIL.n285 VTAIL.n284 9.3005
R1641 VTAIL.n45 VTAIL.n44 9.3005
R1642 VTAIL.n14 VTAIL.n13 9.3005
R1643 VTAIL.n39 VTAIL.n38 9.3005
R1644 VTAIL.n37 VTAIL.n36 9.3005
R1645 VTAIL.n18 VTAIL.n17 9.3005
R1646 VTAIL.n31 VTAIL.n30 9.3005
R1647 VTAIL.n29 VTAIL.n28 9.3005
R1648 VTAIL.n22 VTAIL.n21 9.3005
R1649 VTAIL.n47 VTAIL.n46 9.3005
R1650 VTAIL.n10 VTAIL.n9 9.3005
R1651 VTAIL.n53 VTAIL.n52 9.3005
R1652 VTAIL.n55 VTAIL.n54 9.3005
R1653 VTAIL.n6 VTAIL.n5 9.3005
R1654 VTAIL.n61 VTAIL.n60 9.3005
R1655 VTAIL.n63 VTAIL.n62 9.3005
R1656 VTAIL.n2 VTAIL.n1 9.3005
R1657 VTAIL.n69 VTAIL.n68 9.3005
R1658 VTAIL.n154 VTAIL.n153 9.3005
R1659 VTAIL.n197 VTAIL.n196 9.3005
R1660 VTAIL.n199 VTAIL.n198 9.3005
R1661 VTAIL.n150 VTAIL.n149 9.3005
R1662 VTAIL.n205 VTAIL.n204 9.3005
R1663 VTAIL.n207 VTAIL.n206 9.3005
R1664 VTAIL.n146 VTAIL.n145 9.3005
R1665 VTAIL.n213 VTAIL.n212 9.3005
R1666 VTAIL.n191 VTAIL.n190 9.3005
R1667 VTAIL.n189 VTAIL.n188 9.3005
R1668 VTAIL.n158 VTAIL.n157 9.3005
R1669 VTAIL.n183 VTAIL.n182 9.3005
R1670 VTAIL.n181 VTAIL.n180 9.3005
R1671 VTAIL.n162 VTAIL.n161 9.3005
R1672 VTAIL.n175 VTAIL.n174 9.3005
R1673 VTAIL.n173 VTAIL.n172 9.3005
R1674 VTAIL.n166 VTAIL.n165 9.3005
R1675 VTAIL.n82 VTAIL.n81 9.3005
R1676 VTAIL.n125 VTAIL.n124 9.3005
R1677 VTAIL.n127 VTAIL.n126 9.3005
R1678 VTAIL.n78 VTAIL.n77 9.3005
R1679 VTAIL.n133 VTAIL.n132 9.3005
R1680 VTAIL.n135 VTAIL.n134 9.3005
R1681 VTAIL.n74 VTAIL.n73 9.3005
R1682 VTAIL.n141 VTAIL.n140 9.3005
R1683 VTAIL.n119 VTAIL.n118 9.3005
R1684 VTAIL.n117 VTAIL.n116 9.3005
R1685 VTAIL.n86 VTAIL.n85 9.3005
R1686 VTAIL.n111 VTAIL.n110 9.3005
R1687 VTAIL.n109 VTAIL.n108 9.3005
R1688 VTAIL.n90 VTAIL.n89 9.3005
R1689 VTAIL.n103 VTAIL.n102 9.3005
R1690 VTAIL.n101 VTAIL.n100 9.3005
R1691 VTAIL.n94 VTAIL.n93 9.3005
R1692 VTAIL.n256 VTAIL.n255 8.92171
R1693 VTAIL.n271 VTAIL.n224 8.92171
R1694 VTAIL.n40 VTAIL.n39 8.92171
R1695 VTAIL.n55 VTAIL.n8 8.92171
R1696 VTAIL.n199 VTAIL.n152 8.92171
R1697 VTAIL.n184 VTAIL.n183 8.92171
R1698 VTAIL.n127 VTAIL.n80 8.92171
R1699 VTAIL.n112 VTAIL.n111 8.92171
R1700 VTAIL.n286 VTAIL.n216 8.2187
R1701 VTAIL.n70 VTAIL.n0 8.2187
R1702 VTAIL.n214 VTAIL.n144 8.2187
R1703 VTAIL.n142 VTAIL.n72 8.2187
R1704 VTAIL.n259 VTAIL.n230 8.14595
R1705 VTAIL.n268 VTAIL.n267 8.14595
R1706 VTAIL.n43 VTAIL.n14 8.14595
R1707 VTAIL.n52 VTAIL.n51 8.14595
R1708 VTAIL.n196 VTAIL.n195 8.14595
R1709 VTAIL.n187 VTAIL.n158 8.14595
R1710 VTAIL.n124 VTAIL.n123 8.14595
R1711 VTAIL.n115 VTAIL.n86 8.14595
R1712 VTAIL.n260 VTAIL.n228 7.3702
R1713 VTAIL.n264 VTAIL.n226 7.3702
R1714 VTAIL.n44 VTAIL.n12 7.3702
R1715 VTAIL.n48 VTAIL.n10 7.3702
R1716 VTAIL.n192 VTAIL.n154 7.3702
R1717 VTAIL.n188 VTAIL.n156 7.3702
R1718 VTAIL.n120 VTAIL.n82 7.3702
R1719 VTAIL.n116 VTAIL.n84 7.3702
R1720 VTAIL.n263 VTAIL.n228 6.59444
R1721 VTAIL.n264 VTAIL.n263 6.59444
R1722 VTAIL.n47 VTAIL.n12 6.59444
R1723 VTAIL.n48 VTAIL.n47 6.59444
R1724 VTAIL.n192 VTAIL.n191 6.59444
R1725 VTAIL.n191 VTAIL.n156 6.59444
R1726 VTAIL.n120 VTAIL.n119 6.59444
R1727 VTAIL.n119 VTAIL.n84 6.59444
R1728 VTAIL.n260 VTAIL.n259 5.81868
R1729 VTAIL.n267 VTAIL.n226 5.81868
R1730 VTAIL.n44 VTAIL.n43 5.81868
R1731 VTAIL.n51 VTAIL.n10 5.81868
R1732 VTAIL.n195 VTAIL.n154 5.81868
R1733 VTAIL.n188 VTAIL.n187 5.81868
R1734 VTAIL.n123 VTAIL.n82 5.81868
R1735 VTAIL.n116 VTAIL.n115 5.81868
R1736 VTAIL.n284 VTAIL.n216 5.3904
R1737 VTAIL.n68 VTAIL.n0 5.3904
R1738 VTAIL.n212 VTAIL.n144 5.3904
R1739 VTAIL.n140 VTAIL.n72 5.3904
R1740 VTAIL.n256 VTAIL.n230 5.04292
R1741 VTAIL.n268 VTAIL.n224 5.04292
R1742 VTAIL.n40 VTAIL.n14 5.04292
R1743 VTAIL.n52 VTAIL.n8 5.04292
R1744 VTAIL.n196 VTAIL.n152 5.04292
R1745 VTAIL.n184 VTAIL.n158 5.04292
R1746 VTAIL.n124 VTAIL.n80 5.04292
R1747 VTAIL.n112 VTAIL.n86 5.04292
R1748 VTAIL.n239 VTAIL.n237 4.38563
R1749 VTAIL.n23 VTAIL.n21 4.38563
R1750 VTAIL.n167 VTAIL.n165 4.38563
R1751 VTAIL.n95 VTAIL.n93 4.38563
R1752 VTAIL.n255 VTAIL.n232 4.26717
R1753 VTAIL.n272 VTAIL.n271 4.26717
R1754 VTAIL.n39 VTAIL.n16 4.26717
R1755 VTAIL.n56 VTAIL.n55 4.26717
R1756 VTAIL.n200 VTAIL.n199 4.26717
R1757 VTAIL.n183 VTAIL.n160 4.26717
R1758 VTAIL.n128 VTAIL.n127 4.26717
R1759 VTAIL.n111 VTAIL.n88 4.26717
R1760 VTAIL.n252 VTAIL.n251 3.49141
R1761 VTAIL.n275 VTAIL.n222 3.49141
R1762 VTAIL.n36 VTAIL.n35 3.49141
R1763 VTAIL.n59 VTAIL.n6 3.49141
R1764 VTAIL.n203 VTAIL.n150 3.49141
R1765 VTAIL.n180 VTAIL.n179 3.49141
R1766 VTAIL.n131 VTAIL.n78 3.49141
R1767 VTAIL.n108 VTAIL.n107 3.49141
R1768 VTAIL.n248 VTAIL.n234 2.71565
R1769 VTAIL.n276 VTAIL.n220 2.71565
R1770 VTAIL.n32 VTAIL.n18 2.71565
R1771 VTAIL.n60 VTAIL.n4 2.71565
R1772 VTAIL.n204 VTAIL.n148 2.71565
R1773 VTAIL.n176 VTAIL.n162 2.71565
R1774 VTAIL.n132 VTAIL.n76 2.71565
R1775 VTAIL.n104 VTAIL.n90 2.71565
R1776 VTAIL.n215 VTAIL.n143 2.25912
R1777 VTAIL.n247 VTAIL.n236 1.93989
R1778 VTAIL.n280 VTAIL.n279 1.93989
R1779 VTAIL.n31 VTAIL.n20 1.93989
R1780 VTAIL.n64 VTAIL.n63 1.93989
R1781 VTAIL.n208 VTAIL.n207 1.93989
R1782 VTAIL.n175 VTAIL.n164 1.93989
R1783 VTAIL.n136 VTAIL.n135 1.93989
R1784 VTAIL.n103 VTAIL.n92 1.93989
R1785 VTAIL VTAIL.n71 1.42291
R1786 VTAIL.n244 VTAIL.n243 1.16414
R1787 VTAIL.n283 VTAIL.n218 1.16414
R1788 VTAIL.n28 VTAIL.n27 1.16414
R1789 VTAIL.n67 VTAIL.n2 1.16414
R1790 VTAIL.n211 VTAIL.n146 1.16414
R1791 VTAIL.n172 VTAIL.n171 1.16414
R1792 VTAIL.n139 VTAIL.n74 1.16414
R1793 VTAIL.n100 VTAIL.n99 1.16414
R1794 VTAIL VTAIL.n287 0.836707
R1795 VTAIL.n240 VTAIL.n238 0.388379
R1796 VTAIL.n24 VTAIL.n22 0.388379
R1797 VTAIL.n168 VTAIL.n166 0.388379
R1798 VTAIL.n96 VTAIL.n94 0.388379
R1799 VTAIL.n245 VTAIL.n237 0.155672
R1800 VTAIL.n246 VTAIL.n245 0.155672
R1801 VTAIL.n246 VTAIL.n233 0.155672
R1802 VTAIL.n253 VTAIL.n233 0.155672
R1803 VTAIL.n254 VTAIL.n253 0.155672
R1804 VTAIL.n254 VTAIL.n229 0.155672
R1805 VTAIL.n261 VTAIL.n229 0.155672
R1806 VTAIL.n262 VTAIL.n261 0.155672
R1807 VTAIL.n262 VTAIL.n225 0.155672
R1808 VTAIL.n269 VTAIL.n225 0.155672
R1809 VTAIL.n270 VTAIL.n269 0.155672
R1810 VTAIL.n270 VTAIL.n221 0.155672
R1811 VTAIL.n277 VTAIL.n221 0.155672
R1812 VTAIL.n278 VTAIL.n277 0.155672
R1813 VTAIL.n278 VTAIL.n217 0.155672
R1814 VTAIL.n285 VTAIL.n217 0.155672
R1815 VTAIL.n29 VTAIL.n21 0.155672
R1816 VTAIL.n30 VTAIL.n29 0.155672
R1817 VTAIL.n30 VTAIL.n17 0.155672
R1818 VTAIL.n37 VTAIL.n17 0.155672
R1819 VTAIL.n38 VTAIL.n37 0.155672
R1820 VTAIL.n38 VTAIL.n13 0.155672
R1821 VTAIL.n45 VTAIL.n13 0.155672
R1822 VTAIL.n46 VTAIL.n45 0.155672
R1823 VTAIL.n46 VTAIL.n9 0.155672
R1824 VTAIL.n53 VTAIL.n9 0.155672
R1825 VTAIL.n54 VTAIL.n53 0.155672
R1826 VTAIL.n54 VTAIL.n5 0.155672
R1827 VTAIL.n61 VTAIL.n5 0.155672
R1828 VTAIL.n62 VTAIL.n61 0.155672
R1829 VTAIL.n62 VTAIL.n1 0.155672
R1830 VTAIL.n69 VTAIL.n1 0.155672
R1831 VTAIL.n213 VTAIL.n145 0.155672
R1832 VTAIL.n206 VTAIL.n145 0.155672
R1833 VTAIL.n206 VTAIL.n205 0.155672
R1834 VTAIL.n205 VTAIL.n149 0.155672
R1835 VTAIL.n198 VTAIL.n149 0.155672
R1836 VTAIL.n198 VTAIL.n197 0.155672
R1837 VTAIL.n197 VTAIL.n153 0.155672
R1838 VTAIL.n190 VTAIL.n153 0.155672
R1839 VTAIL.n190 VTAIL.n189 0.155672
R1840 VTAIL.n189 VTAIL.n157 0.155672
R1841 VTAIL.n182 VTAIL.n157 0.155672
R1842 VTAIL.n182 VTAIL.n181 0.155672
R1843 VTAIL.n181 VTAIL.n161 0.155672
R1844 VTAIL.n174 VTAIL.n161 0.155672
R1845 VTAIL.n174 VTAIL.n173 0.155672
R1846 VTAIL.n173 VTAIL.n165 0.155672
R1847 VTAIL.n141 VTAIL.n73 0.155672
R1848 VTAIL.n134 VTAIL.n73 0.155672
R1849 VTAIL.n134 VTAIL.n133 0.155672
R1850 VTAIL.n133 VTAIL.n77 0.155672
R1851 VTAIL.n126 VTAIL.n77 0.155672
R1852 VTAIL.n126 VTAIL.n125 0.155672
R1853 VTAIL.n125 VTAIL.n81 0.155672
R1854 VTAIL.n118 VTAIL.n81 0.155672
R1855 VTAIL.n118 VTAIL.n117 0.155672
R1856 VTAIL.n117 VTAIL.n85 0.155672
R1857 VTAIL.n110 VTAIL.n85 0.155672
R1858 VTAIL.n110 VTAIL.n109 0.155672
R1859 VTAIL.n109 VTAIL.n89 0.155672
R1860 VTAIL.n102 VTAIL.n89 0.155672
R1861 VTAIL.n102 VTAIL.n101 0.155672
R1862 VTAIL.n101 VTAIL.n93 0.155672
R1863 VDD1.n66 VDD1.n0 214.453
R1864 VDD1.n137 VDD1.n71 214.453
R1865 VDD1.n67 VDD1.n66 185
R1866 VDD1.n65 VDD1.n64 185
R1867 VDD1.n4 VDD1.n3 185
R1868 VDD1.n59 VDD1.n58 185
R1869 VDD1.n57 VDD1.n56 185
R1870 VDD1.n8 VDD1.n7 185
R1871 VDD1.n51 VDD1.n50 185
R1872 VDD1.n49 VDD1.n48 185
R1873 VDD1.n12 VDD1.n11 185
R1874 VDD1.n43 VDD1.n42 185
R1875 VDD1.n41 VDD1.n40 185
R1876 VDD1.n16 VDD1.n15 185
R1877 VDD1.n35 VDD1.n34 185
R1878 VDD1.n33 VDD1.n32 185
R1879 VDD1.n20 VDD1.n19 185
R1880 VDD1.n27 VDD1.n26 185
R1881 VDD1.n25 VDD1.n24 185
R1882 VDD1.n96 VDD1.n95 185
R1883 VDD1.n98 VDD1.n97 185
R1884 VDD1.n91 VDD1.n90 185
R1885 VDD1.n104 VDD1.n103 185
R1886 VDD1.n106 VDD1.n105 185
R1887 VDD1.n87 VDD1.n86 185
R1888 VDD1.n112 VDD1.n111 185
R1889 VDD1.n114 VDD1.n113 185
R1890 VDD1.n83 VDD1.n82 185
R1891 VDD1.n120 VDD1.n119 185
R1892 VDD1.n122 VDD1.n121 185
R1893 VDD1.n79 VDD1.n78 185
R1894 VDD1.n128 VDD1.n127 185
R1895 VDD1.n130 VDD1.n129 185
R1896 VDD1.n75 VDD1.n74 185
R1897 VDD1.n136 VDD1.n135 185
R1898 VDD1.n138 VDD1.n137 185
R1899 VDD1.n94 VDD1.t1 147.659
R1900 VDD1.n23 VDD1.t0 147.659
R1901 VDD1.n66 VDD1.n65 104.615
R1902 VDD1.n65 VDD1.n3 104.615
R1903 VDD1.n58 VDD1.n3 104.615
R1904 VDD1.n58 VDD1.n57 104.615
R1905 VDD1.n57 VDD1.n7 104.615
R1906 VDD1.n50 VDD1.n7 104.615
R1907 VDD1.n50 VDD1.n49 104.615
R1908 VDD1.n49 VDD1.n11 104.615
R1909 VDD1.n42 VDD1.n11 104.615
R1910 VDD1.n42 VDD1.n41 104.615
R1911 VDD1.n41 VDD1.n15 104.615
R1912 VDD1.n34 VDD1.n15 104.615
R1913 VDD1.n34 VDD1.n33 104.615
R1914 VDD1.n33 VDD1.n19 104.615
R1915 VDD1.n26 VDD1.n19 104.615
R1916 VDD1.n26 VDD1.n25 104.615
R1917 VDD1.n97 VDD1.n96 104.615
R1918 VDD1.n97 VDD1.n90 104.615
R1919 VDD1.n104 VDD1.n90 104.615
R1920 VDD1.n105 VDD1.n104 104.615
R1921 VDD1.n105 VDD1.n86 104.615
R1922 VDD1.n112 VDD1.n86 104.615
R1923 VDD1.n113 VDD1.n112 104.615
R1924 VDD1.n113 VDD1.n82 104.615
R1925 VDD1.n120 VDD1.n82 104.615
R1926 VDD1.n121 VDD1.n120 104.615
R1927 VDD1.n121 VDD1.n78 104.615
R1928 VDD1.n128 VDD1.n78 104.615
R1929 VDD1.n129 VDD1.n128 104.615
R1930 VDD1.n129 VDD1.n74 104.615
R1931 VDD1.n136 VDD1.n74 104.615
R1932 VDD1.n137 VDD1.n136 104.615
R1933 VDD1 VDD1.n141 94.3003
R1934 VDD1.n25 VDD1.t0 52.3082
R1935 VDD1.n96 VDD1.t1 52.3082
R1936 VDD1 VDD1.n70 51.5622
R1937 VDD1.n24 VDD1.n23 15.6677
R1938 VDD1.n95 VDD1.n94 15.6677
R1939 VDD1.n68 VDD1.n67 12.8005
R1940 VDD1.n27 VDD1.n22 12.8005
R1941 VDD1.n98 VDD1.n93 12.8005
R1942 VDD1.n139 VDD1.n138 12.8005
R1943 VDD1.n64 VDD1.n2 12.0247
R1944 VDD1.n28 VDD1.n20 12.0247
R1945 VDD1.n99 VDD1.n91 12.0247
R1946 VDD1.n135 VDD1.n73 12.0247
R1947 VDD1.n63 VDD1.n4 11.249
R1948 VDD1.n32 VDD1.n31 11.249
R1949 VDD1.n103 VDD1.n102 11.249
R1950 VDD1.n134 VDD1.n75 11.249
R1951 VDD1.n60 VDD1.n59 10.4732
R1952 VDD1.n35 VDD1.n18 10.4732
R1953 VDD1.n106 VDD1.n89 10.4732
R1954 VDD1.n131 VDD1.n130 10.4732
R1955 VDD1.n56 VDD1.n6 9.69747
R1956 VDD1.n36 VDD1.n16 9.69747
R1957 VDD1.n107 VDD1.n87 9.69747
R1958 VDD1.n127 VDD1.n77 9.69747
R1959 VDD1.n70 VDD1.n69 9.45567
R1960 VDD1.n141 VDD1.n140 9.45567
R1961 VDD1.n10 VDD1.n9 9.3005
R1962 VDD1.n53 VDD1.n52 9.3005
R1963 VDD1.n55 VDD1.n54 9.3005
R1964 VDD1.n6 VDD1.n5 9.3005
R1965 VDD1.n61 VDD1.n60 9.3005
R1966 VDD1.n63 VDD1.n62 9.3005
R1967 VDD1.n2 VDD1.n1 9.3005
R1968 VDD1.n69 VDD1.n68 9.3005
R1969 VDD1.n47 VDD1.n46 9.3005
R1970 VDD1.n45 VDD1.n44 9.3005
R1971 VDD1.n14 VDD1.n13 9.3005
R1972 VDD1.n39 VDD1.n38 9.3005
R1973 VDD1.n37 VDD1.n36 9.3005
R1974 VDD1.n18 VDD1.n17 9.3005
R1975 VDD1.n31 VDD1.n30 9.3005
R1976 VDD1.n29 VDD1.n28 9.3005
R1977 VDD1.n22 VDD1.n21 9.3005
R1978 VDD1.n116 VDD1.n115 9.3005
R1979 VDD1.n85 VDD1.n84 9.3005
R1980 VDD1.n110 VDD1.n109 9.3005
R1981 VDD1.n108 VDD1.n107 9.3005
R1982 VDD1.n89 VDD1.n88 9.3005
R1983 VDD1.n102 VDD1.n101 9.3005
R1984 VDD1.n100 VDD1.n99 9.3005
R1985 VDD1.n93 VDD1.n92 9.3005
R1986 VDD1.n118 VDD1.n117 9.3005
R1987 VDD1.n81 VDD1.n80 9.3005
R1988 VDD1.n124 VDD1.n123 9.3005
R1989 VDD1.n126 VDD1.n125 9.3005
R1990 VDD1.n77 VDD1.n76 9.3005
R1991 VDD1.n132 VDD1.n131 9.3005
R1992 VDD1.n134 VDD1.n133 9.3005
R1993 VDD1.n73 VDD1.n72 9.3005
R1994 VDD1.n140 VDD1.n139 9.3005
R1995 VDD1.n55 VDD1.n8 8.92171
R1996 VDD1.n40 VDD1.n39 8.92171
R1997 VDD1.n111 VDD1.n110 8.92171
R1998 VDD1.n126 VDD1.n79 8.92171
R1999 VDD1.n70 VDD1.n0 8.2187
R2000 VDD1.n141 VDD1.n71 8.2187
R2001 VDD1.n52 VDD1.n51 8.14595
R2002 VDD1.n43 VDD1.n14 8.14595
R2003 VDD1.n114 VDD1.n85 8.14595
R2004 VDD1.n123 VDD1.n122 8.14595
R2005 VDD1.n48 VDD1.n10 7.3702
R2006 VDD1.n44 VDD1.n12 7.3702
R2007 VDD1.n115 VDD1.n83 7.3702
R2008 VDD1.n119 VDD1.n81 7.3702
R2009 VDD1.n48 VDD1.n47 6.59444
R2010 VDD1.n47 VDD1.n12 6.59444
R2011 VDD1.n118 VDD1.n83 6.59444
R2012 VDD1.n119 VDD1.n118 6.59444
R2013 VDD1.n51 VDD1.n10 5.81868
R2014 VDD1.n44 VDD1.n43 5.81868
R2015 VDD1.n115 VDD1.n114 5.81868
R2016 VDD1.n122 VDD1.n81 5.81868
R2017 VDD1.n68 VDD1.n0 5.3904
R2018 VDD1.n139 VDD1.n71 5.3904
R2019 VDD1.n52 VDD1.n8 5.04292
R2020 VDD1.n40 VDD1.n14 5.04292
R2021 VDD1.n111 VDD1.n85 5.04292
R2022 VDD1.n123 VDD1.n79 5.04292
R2023 VDD1.n94 VDD1.n92 4.38563
R2024 VDD1.n23 VDD1.n21 4.38563
R2025 VDD1.n56 VDD1.n55 4.26717
R2026 VDD1.n39 VDD1.n16 4.26717
R2027 VDD1.n110 VDD1.n87 4.26717
R2028 VDD1.n127 VDD1.n126 4.26717
R2029 VDD1.n59 VDD1.n6 3.49141
R2030 VDD1.n36 VDD1.n35 3.49141
R2031 VDD1.n107 VDD1.n106 3.49141
R2032 VDD1.n130 VDD1.n77 3.49141
R2033 VDD1.n60 VDD1.n4 2.71565
R2034 VDD1.n32 VDD1.n18 2.71565
R2035 VDD1.n103 VDD1.n89 2.71565
R2036 VDD1.n131 VDD1.n75 2.71565
R2037 VDD1.n64 VDD1.n63 1.93989
R2038 VDD1.n31 VDD1.n20 1.93989
R2039 VDD1.n102 VDD1.n91 1.93989
R2040 VDD1.n135 VDD1.n134 1.93989
R2041 VDD1.n67 VDD1.n2 1.16414
R2042 VDD1.n28 VDD1.n27 1.16414
R2043 VDD1.n99 VDD1.n98 1.16414
R2044 VDD1.n138 VDD1.n73 1.16414
R2045 VDD1.n24 VDD1.n22 0.388379
R2046 VDD1.n95 VDD1.n93 0.388379
R2047 VDD1.n69 VDD1.n1 0.155672
R2048 VDD1.n62 VDD1.n1 0.155672
R2049 VDD1.n62 VDD1.n61 0.155672
R2050 VDD1.n61 VDD1.n5 0.155672
R2051 VDD1.n54 VDD1.n5 0.155672
R2052 VDD1.n54 VDD1.n53 0.155672
R2053 VDD1.n53 VDD1.n9 0.155672
R2054 VDD1.n46 VDD1.n9 0.155672
R2055 VDD1.n46 VDD1.n45 0.155672
R2056 VDD1.n45 VDD1.n13 0.155672
R2057 VDD1.n38 VDD1.n13 0.155672
R2058 VDD1.n38 VDD1.n37 0.155672
R2059 VDD1.n37 VDD1.n17 0.155672
R2060 VDD1.n30 VDD1.n17 0.155672
R2061 VDD1.n30 VDD1.n29 0.155672
R2062 VDD1.n29 VDD1.n21 0.155672
R2063 VDD1.n100 VDD1.n92 0.155672
R2064 VDD1.n101 VDD1.n100 0.155672
R2065 VDD1.n101 VDD1.n88 0.155672
R2066 VDD1.n108 VDD1.n88 0.155672
R2067 VDD1.n109 VDD1.n108 0.155672
R2068 VDD1.n109 VDD1.n84 0.155672
R2069 VDD1.n116 VDD1.n84 0.155672
R2070 VDD1.n117 VDD1.n116 0.155672
R2071 VDD1.n117 VDD1.n80 0.155672
R2072 VDD1.n124 VDD1.n80 0.155672
R2073 VDD1.n125 VDD1.n124 0.155672
R2074 VDD1.n125 VDD1.n76 0.155672
R2075 VDD1.n132 VDD1.n76 0.155672
R2076 VDD1.n133 VDD1.n132 0.155672
R2077 VDD1.n133 VDD1.n72 0.155672
R2078 VDD1.n140 VDD1.n72 0.155672
R2079 VN VN.t0 167.565
R2080 VN VN.t1 119.504
R2081 VDD2.n137 VDD2.n71 214.453
R2082 VDD2.n66 VDD2.n0 214.453
R2083 VDD2.n138 VDD2.n137 185
R2084 VDD2.n136 VDD2.n135 185
R2085 VDD2.n75 VDD2.n74 185
R2086 VDD2.n130 VDD2.n129 185
R2087 VDD2.n128 VDD2.n127 185
R2088 VDD2.n79 VDD2.n78 185
R2089 VDD2.n122 VDD2.n121 185
R2090 VDD2.n120 VDD2.n119 185
R2091 VDD2.n83 VDD2.n82 185
R2092 VDD2.n114 VDD2.n113 185
R2093 VDD2.n112 VDD2.n111 185
R2094 VDD2.n87 VDD2.n86 185
R2095 VDD2.n106 VDD2.n105 185
R2096 VDD2.n104 VDD2.n103 185
R2097 VDD2.n91 VDD2.n90 185
R2098 VDD2.n98 VDD2.n97 185
R2099 VDD2.n96 VDD2.n95 185
R2100 VDD2.n25 VDD2.n24 185
R2101 VDD2.n27 VDD2.n26 185
R2102 VDD2.n20 VDD2.n19 185
R2103 VDD2.n33 VDD2.n32 185
R2104 VDD2.n35 VDD2.n34 185
R2105 VDD2.n16 VDD2.n15 185
R2106 VDD2.n41 VDD2.n40 185
R2107 VDD2.n43 VDD2.n42 185
R2108 VDD2.n12 VDD2.n11 185
R2109 VDD2.n49 VDD2.n48 185
R2110 VDD2.n51 VDD2.n50 185
R2111 VDD2.n8 VDD2.n7 185
R2112 VDD2.n57 VDD2.n56 185
R2113 VDD2.n59 VDD2.n58 185
R2114 VDD2.n4 VDD2.n3 185
R2115 VDD2.n65 VDD2.n64 185
R2116 VDD2.n67 VDD2.n66 185
R2117 VDD2.n23 VDD2.t0 147.659
R2118 VDD2.n94 VDD2.t1 147.659
R2119 VDD2.n137 VDD2.n136 104.615
R2120 VDD2.n136 VDD2.n74 104.615
R2121 VDD2.n129 VDD2.n74 104.615
R2122 VDD2.n129 VDD2.n128 104.615
R2123 VDD2.n128 VDD2.n78 104.615
R2124 VDD2.n121 VDD2.n78 104.615
R2125 VDD2.n121 VDD2.n120 104.615
R2126 VDD2.n120 VDD2.n82 104.615
R2127 VDD2.n113 VDD2.n82 104.615
R2128 VDD2.n113 VDD2.n112 104.615
R2129 VDD2.n112 VDD2.n86 104.615
R2130 VDD2.n105 VDD2.n86 104.615
R2131 VDD2.n105 VDD2.n104 104.615
R2132 VDD2.n104 VDD2.n90 104.615
R2133 VDD2.n97 VDD2.n90 104.615
R2134 VDD2.n97 VDD2.n96 104.615
R2135 VDD2.n26 VDD2.n25 104.615
R2136 VDD2.n26 VDD2.n19 104.615
R2137 VDD2.n33 VDD2.n19 104.615
R2138 VDD2.n34 VDD2.n33 104.615
R2139 VDD2.n34 VDD2.n15 104.615
R2140 VDD2.n41 VDD2.n15 104.615
R2141 VDD2.n42 VDD2.n41 104.615
R2142 VDD2.n42 VDD2.n11 104.615
R2143 VDD2.n49 VDD2.n11 104.615
R2144 VDD2.n50 VDD2.n49 104.615
R2145 VDD2.n50 VDD2.n7 104.615
R2146 VDD2.n57 VDD2.n7 104.615
R2147 VDD2.n58 VDD2.n57 104.615
R2148 VDD2.n58 VDD2.n3 104.615
R2149 VDD2.n65 VDD2.n3 104.615
R2150 VDD2.n66 VDD2.n65 104.615
R2151 VDD2.n142 VDD2.n70 92.8811
R2152 VDD2.n96 VDD2.t1 52.3082
R2153 VDD2.n25 VDD2.t0 52.3082
R2154 VDD2.n142 VDD2.n141 50.6096
R2155 VDD2.n95 VDD2.n94 15.6677
R2156 VDD2.n24 VDD2.n23 15.6677
R2157 VDD2.n139 VDD2.n138 12.8005
R2158 VDD2.n98 VDD2.n93 12.8005
R2159 VDD2.n27 VDD2.n22 12.8005
R2160 VDD2.n68 VDD2.n67 12.8005
R2161 VDD2.n135 VDD2.n73 12.0247
R2162 VDD2.n99 VDD2.n91 12.0247
R2163 VDD2.n28 VDD2.n20 12.0247
R2164 VDD2.n64 VDD2.n2 12.0247
R2165 VDD2.n134 VDD2.n75 11.249
R2166 VDD2.n103 VDD2.n102 11.249
R2167 VDD2.n32 VDD2.n31 11.249
R2168 VDD2.n63 VDD2.n4 11.249
R2169 VDD2.n131 VDD2.n130 10.4732
R2170 VDD2.n106 VDD2.n89 10.4732
R2171 VDD2.n35 VDD2.n18 10.4732
R2172 VDD2.n60 VDD2.n59 10.4732
R2173 VDD2.n127 VDD2.n77 9.69747
R2174 VDD2.n107 VDD2.n87 9.69747
R2175 VDD2.n36 VDD2.n16 9.69747
R2176 VDD2.n56 VDD2.n6 9.69747
R2177 VDD2.n141 VDD2.n140 9.45567
R2178 VDD2.n70 VDD2.n69 9.45567
R2179 VDD2.n81 VDD2.n80 9.3005
R2180 VDD2.n124 VDD2.n123 9.3005
R2181 VDD2.n126 VDD2.n125 9.3005
R2182 VDD2.n77 VDD2.n76 9.3005
R2183 VDD2.n132 VDD2.n131 9.3005
R2184 VDD2.n134 VDD2.n133 9.3005
R2185 VDD2.n73 VDD2.n72 9.3005
R2186 VDD2.n140 VDD2.n139 9.3005
R2187 VDD2.n118 VDD2.n117 9.3005
R2188 VDD2.n116 VDD2.n115 9.3005
R2189 VDD2.n85 VDD2.n84 9.3005
R2190 VDD2.n110 VDD2.n109 9.3005
R2191 VDD2.n108 VDD2.n107 9.3005
R2192 VDD2.n89 VDD2.n88 9.3005
R2193 VDD2.n102 VDD2.n101 9.3005
R2194 VDD2.n100 VDD2.n99 9.3005
R2195 VDD2.n93 VDD2.n92 9.3005
R2196 VDD2.n45 VDD2.n44 9.3005
R2197 VDD2.n14 VDD2.n13 9.3005
R2198 VDD2.n39 VDD2.n38 9.3005
R2199 VDD2.n37 VDD2.n36 9.3005
R2200 VDD2.n18 VDD2.n17 9.3005
R2201 VDD2.n31 VDD2.n30 9.3005
R2202 VDD2.n29 VDD2.n28 9.3005
R2203 VDD2.n22 VDD2.n21 9.3005
R2204 VDD2.n47 VDD2.n46 9.3005
R2205 VDD2.n10 VDD2.n9 9.3005
R2206 VDD2.n53 VDD2.n52 9.3005
R2207 VDD2.n55 VDD2.n54 9.3005
R2208 VDD2.n6 VDD2.n5 9.3005
R2209 VDD2.n61 VDD2.n60 9.3005
R2210 VDD2.n63 VDD2.n62 9.3005
R2211 VDD2.n2 VDD2.n1 9.3005
R2212 VDD2.n69 VDD2.n68 9.3005
R2213 VDD2.n126 VDD2.n79 8.92171
R2214 VDD2.n111 VDD2.n110 8.92171
R2215 VDD2.n40 VDD2.n39 8.92171
R2216 VDD2.n55 VDD2.n8 8.92171
R2217 VDD2.n141 VDD2.n71 8.2187
R2218 VDD2.n70 VDD2.n0 8.2187
R2219 VDD2.n123 VDD2.n122 8.14595
R2220 VDD2.n114 VDD2.n85 8.14595
R2221 VDD2.n43 VDD2.n14 8.14595
R2222 VDD2.n52 VDD2.n51 8.14595
R2223 VDD2.n119 VDD2.n81 7.3702
R2224 VDD2.n115 VDD2.n83 7.3702
R2225 VDD2.n44 VDD2.n12 7.3702
R2226 VDD2.n48 VDD2.n10 7.3702
R2227 VDD2.n119 VDD2.n118 6.59444
R2228 VDD2.n118 VDD2.n83 6.59444
R2229 VDD2.n47 VDD2.n12 6.59444
R2230 VDD2.n48 VDD2.n47 6.59444
R2231 VDD2.n122 VDD2.n81 5.81868
R2232 VDD2.n115 VDD2.n114 5.81868
R2233 VDD2.n44 VDD2.n43 5.81868
R2234 VDD2.n51 VDD2.n10 5.81868
R2235 VDD2.n139 VDD2.n71 5.3904
R2236 VDD2.n68 VDD2.n0 5.3904
R2237 VDD2.n123 VDD2.n79 5.04292
R2238 VDD2.n111 VDD2.n85 5.04292
R2239 VDD2.n40 VDD2.n14 5.04292
R2240 VDD2.n52 VDD2.n8 5.04292
R2241 VDD2.n23 VDD2.n21 4.38563
R2242 VDD2.n94 VDD2.n92 4.38563
R2243 VDD2.n127 VDD2.n126 4.26717
R2244 VDD2.n110 VDD2.n87 4.26717
R2245 VDD2.n39 VDD2.n16 4.26717
R2246 VDD2.n56 VDD2.n55 4.26717
R2247 VDD2.n130 VDD2.n77 3.49141
R2248 VDD2.n107 VDD2.n106 3.49141
R2249 VDD2.n36 VDD2.n35 3.49141
R2250 VDD2.n59 VDD2.n6 3.49141
R2251 VDD2.n131 VDD2.n75 2.71565
R2252 VDD2.n103 VDD2.n89 2.71565
R2253 VDD2.n32 VDD2.n18 2.71565
R2254 VDD2.n60 VDD2.n4 2.71565
R2255 VDD2.n135 VDD2.n134 1.93989
R2256 VDD2.n102 VDD2.n91 1.93989
R2257 VDD2.n31 VDD2.n20 1.93989
R2258 VDD2.n64 VDD2.n63 1.93989
R2259 VDD2.n138 VDD2.n73 1.16414
R2260 VDD2.n99 VDD2.n98 1.16414
R2261 VDD2.n28 VDD2.n27 1.16414
R2262 VDD2.n67 VDD2.n2 1.16414
R2263 VDD2 VDD2.n142 0.953086
R2264 VDD2.n95 VDD2.n93 0.388379
R2265 VDD2.n24 VDD2.n22 0.388379
R2266 VDD2.n140 VDD2.n72 0.155672
R2267 VDD2.n133 VDD2.n72 0.155672
R2268 VDD2.n133 VDD2.n132 0.155672
R2269 VDD2.n132 VDD2.n76 0.155672
R2270 VDD2.n125 VDD2.n76 0.155672
R2271 VDD2.n125 VDD2.n124 0.155672
R2272 VDD2.n124 VDD2.n80 0.155672
R2273 VDD2.n117 VDD2.n80 0.155672
R2274 VDD2.n117 VDD2.n116 0.155672
R2275 VDD2.n116 VDD2.n84 0.155672
R2276 VDD2.n109 VDD2.n84 0.155672
R2277 VDD2.n109 VDD2.n108 0.155672
R2278 VDD2.n108 VDD2.n88 0.155672
R2279 VDD2.n101 VDD2.n88 0.155672
R2280 VDD2.n101 VDD2.n100 0.155672
R2281 VDD2.n100 VDD2.n92 0.155672
R2282 VDD2.n29 VDD2.n21 0.155672
R2283 VDD2.n30 VDD2.n29 0.155672
R2284 VDD2.n30 VDD2.n17 0.155672
R2285 VDD2.n37 VDD2.n17 0.155672
R2286 VDD2.n38 VDD2.n37 0.155672
R2287 VDD2.n38 VDD2.n13 0.155672
R2288 VDD2.n45 VDD2.n13 0.155672
R2289 VDD2.n46 VDD2.n45 0.155672
R2290 VDD2.n46 VDD2.n9 0.155672
R2291 VDD2.n53 VDD2.n9 0.155672
R2292 VDD2.n54 VDD2.n53 0.155672
R2293 VDD2.n54 VDD2.n5 0.155672
R2294 VDD2.n61 VDD2.n5 0.155672
R2295 VDD2.n62 VDD2.n61 0.155672
R2296 VDD2.n62 VDD2.n1 0.155672
R2297 VDD2.n69 VDD2.n1 0.155672
C0 VTAIL VP 2.90325f
C1 VDD1 VP 3.44261f
C2 VTAIL VDD1 5.639471f
C3 VDD2 VP 0.383821f
C4 VDD2 VTAIL 5.69904f
C5 VDD2 VDD1 0.810601f
C6 VN VP 6.26902f
C7 VTAIL VN 2.88842f
C8 VN VDD1 0.148683f
C9 VDD2 VN 3.20911f
C10 VDD2 B 5.10418f
C11 VDD1 B 8.17385f
C12 VTAIL B 8.468237f
C13 VN B 12.260631f
C14 VP B 8.004513f
C15 VDD2.n0 B 0.027076f
C16 VDD2.n1 B 0.020356f
C17 VDD2.n2 B 0.010939f
C18 VDD2.n3 B 0.025855f
C19 VDD2.n4 B 0.011582f
C20 VDD2.n5 B 0.020356f
C21 VDD2.n6 B 0.010939f
C22 VDD2.n7 B 0.025855f
C23 VDD2.n8 B 0.011582f
C24 VDD2.n9 B 0.020356f
C25 VDD2.n10 B 0.010939f
C26 VDD2.n11 B 0.025855f
C27 VDD2.n12 B 0.011582f
C28 VDD2.n13 B 0.020356f
C29 VDD2.n14 B 0.010939f
C30 VDD2.n15 B 0.025855f
C31 VDD2.n16 B 0.011582f
C32 VDD2.n17 B 0.020356f
C33 VDD2.n18 B 0.010939f
C34 VDD2.n19 B 0.025855f
C35 VDD2.n20 B 0.011582f
C36 VDD2.n21 B 1.16488f
C37 VDD2.n22 B 0.010939f
C38 VDD2.t0 B 0.042512f
C39 VDD2.n23 B 0.124041f
C40 VDD2.n24 B 0.015273f
C41 VDD2.n25 B 0.019391f
C42 VDD2.n26 B 0.025855f
C43 VDD2.n27 B 0.011582f
C44 VDD2.n28 B 0.010939f
C45 VDD2.n29 B 0.020356f
C46 VDD2.n30 B 0.020356f
C47 VDD2.n31 B 0.010939f
C48 VDD2.n32 B 0.011582f
C49 VDD2.n33 B 0.025855f
C50 VDD2.n34 B 0.025855f
C51 VDD2.n35 B 0.011582f
C52 VDD2.n36 B 0.010939f
C53 VDD2.n37 B 0.020356f
C54 VDD2.n38 B 0.020356f
C55 VDD2.n39 B 0.010939f
C56 VDD2.n40 B 0.011582f
C57 VDD2.n41 B 0.025855f
C58 VDD2.n42 B 0.025855f
C59 VDD2.n43 B 0.011582f
C60 VDD2.n44 B 0.010939f
C61 VDD2.n45 B 0.020356f
C62 VDD2.n46 B 0.020356f
C63 VDD2.n47 B 0.010939f
C64 VDD2.n48 B 0.011582f
C65 VDD2.n49 B 0.025855f
C66 VDD2.n50 B 0.025855f
C67 VDD2.n51 B 0.011582f
C68 VDD2.n52 B 0.010939f
C69 VDD2.n53 B 0.020356f
C70 VDD2.n54 B 0.020356f
C71 VDD2.n55 B 0.010939f
C72 VDD2.n56 B 0.011582f
C73 VDD2.n57 B 0.025855f
C74 VDD2.n58 B 0.025855f
C75 VDD2.n59 B 0.011582f
C76 VDD2.n60 B 0.010939f
C77 VDD2.n61 B 0.020356f
C78 VDD2.n62 B 0.020356f
C79 VDD2.n63 B 0.010939f
C80 VDD2.n64 B 0.011582f
C81 VDD2.n65 B 0.025855f
C82 VDD2.n66 B 0.052159f
C83 VDD2.n67 B 0.011582f
C84 VDD2.n68 B 0.021389f
C85 VDD2.n69 B 0.049556f
C86 VDD2.n70 B 0.713339f
C87 VDD2.n71 B 0.027076f
C88 VDD2.n72 B 0.020356f
C89 VDD2.n73 B 0.010939f
C90 VDD2.n74 B 0.025855f
C91 VDD2.n75 B 0.011582f
C92 VDD2.n76 B 0.020356f
C93 VDD2.n77 B 0.010939f
C94 VDD2.n78 B 0.025855f
C95 VDD2.n79 B 0.011582f
C96 VDD2.n80 B 0.020356f
C97 VDD2.n81 B 0.010939f
C98 VDD2.n82 B 0.025855f
C99 VDD2.n83 B 0.011582f
C100 VDD2.n84 B 0.020356f
C101 VDD2.n85 B 0.010939f
C102 VDD2.n86 B 0.025855f
C103 VDD2.n87 B 0.011582f
C104 VDD2.n88 B 0.020356f
C105 VDD2.n89 B 0.010939f
C106 VDD2.n90 B 0.025855f
C107 VDD2.n91 B 0.011582f
C108 VDD2.n92 B 1.16488f
C109 VDD2.n93 B 0.010939f
C110 VDD2.t1 B 0.042512f
C111 VDD2.n94 B 0.124041f
C112 VDD2.n95 B 0.015273f
C113 VDD2.n96 B 0.019391f
C114 VDD2.n97 B 0.025855f
C115 VDD2.n98 B 0.011582f
C116 VDD2.n99 B 0.010939f
C117 VDD2.n100 B 0.020356f
C118 VDD2.n101 B 0.020356f
C119 VDD2.n102 B 0.010939f
C120 VDD2.n103 B 0.011582f
C121 VDD2.n104 B 0.025855f
C122 VDD2.n105 B 0.025855f
C123 VDD2.n106 B 0.011582f
C124 VDD2.n107 B 0.010939f
C125 VDD2.n108 B 0.020356f
C126 VDD2.n109 B 0.020356f
C127 VDD2.n110 B 0.010939f
C128 VDD2.n111 B 0.011582f
C129 VDD2.n112 B 0.025855f
C130 VDD2.n113 B 0.025855f
C131 VDD2.n114 B 0.011582f
C132 VDD2.n115 B 0.010939f
C133 VDD2.n116 B 0.020356f
C134 VDD2.n117 B 0.020356f
C135 VDD2.n118 B 0.010939f
C136 VDD2.n119 B 0.011582f
C137 VDD2.n120 B 0.025855f
C138 VDD2.n121 B 0.025855f
C139 VDD2.n122 B 0.011582f
C140 VDD2.n123 B 0.010939f
C141 VDD2.n124 B 0.020356f
C142 VDD2.n125 B 0.020356f
C143 VDD2.n126 B 0.010939f
C144 VDD2.n127 B 0.011582f
C145 VDD2.n128 B 0.025855f
C146 VDD2.n129 B 0.025855f
C147 VDD2.n130 B 0.011582f
C148 VDD2.n131 B 0.010939f
C149 VDD2.n132 B 0.020356f
C150 VDD2.n133 B 0.020356f
C151 VDD2.n134 B 0.010939f
C152 VDD2.n135 B 0.011582f
C153 VDD2.n136 B 0.025855f
C154 VDD2.n137 B 0.052159f
C155 VDD2.n138 B 0.011582f
C156 VDD2.n139 B 0.021389f
C157 VDD2.n140 B 0.049556f
C158 VDD2.n141 B 0.066843f
C159 VDD2.n142 B 2.79988f
C160 VN.t1 B 3.73548f
C161 VN.t0 B 4.43978f
C162 VDD1.n0 B 0.02715f
C163 VDD1.n1 B 0.020413f
C164 VDD1.n2 B 0.010969f
C165 VDD1.n3 B 0.025926f
C166 VDD1.n4 B 0.011614f
C167 VDD1.n5 B 0.020413f
C168 VDD1.n6 B 0.010969f
C169 VDD1.n7 B 0.025926f
C170 VDD1.n8 B 0.011614f
C171 VDD1.n9 B 0.020413f
C172 VDD1.n10 B 0.010969f
C173 VDD1.n11 B 0.025926f
C174 VDD1.n12 B 0.011614f
C175 VDD1.n13 B 0.020413f
C176 VDD1.n14 B 0.010969f
C177 VDD1.n15 B 0.025926f
C178 VDD1.n16 B 0.011614f
C179 VDD1.n17 B 0.020413f
C180 VDD1.n18 B 0.010969f
C181 VDD1.n19 B 0.025926f
C182 VDD1.n20 B 0.011614f
C183 VDD1.n21 B 1.1681f
C184 VDD1.n22 B 0.010969f
C185 VDD1.t0 B 0.04263f
C186 VDD1.n23 B 0.124384f
C187 VDD1.n24 B 0.015316f
C188 VDD1.n25 B 0.019445f
C189 VDD1.n26 B 0.025926f
C190 VDD1.n27 B 0.011614f
C191 VDD1.n28 B 0.010969f
C192 VDD1.n29 B 0.020413f
C193 VDD1.n30 B 0.020413f
C194 VDD1.n31 B 0.010969f
C195 VDD1.n32 B 0.011614f
C196 VDD1.n33 B 0.025926f
C197 VDD1.n34 B 0.025926f
C198 VDD1.n35 B 0.011614f
C199 VDD1.n36 B 0.010969f
C200 VDD1.n37 B 0.020413f
C201 VDD1.n38 B 0.020413f
C202 VDD1.n39 B 0.010969f
C203 VDD1.n40 B 0.011614f
C204 VDD1.n41 B 0.025926f
C205 VDD1.n42 B 0.025926f
C206 VDD1.n43 B 0.011614f
C207 VDD1.n44 B 0.010969f
C208 VDD1.n45 B 0.020413f
C209 VDD1.n46 B 0.020413f
C210 VDD1.n47 B 0.010969f
C211 VDD1.n48 B 0.011614f
C212 VDD1.n49 B 0.025926f
C213 VDD1.n50 B 0.025926f
C214 VDD1.n51 B 0.011614f
C215 VDD1.n52 B 0.010969f
C216 VDD1.n53 B 0.020413f
C217 VDD1.n54 B 0.020413f
C218 VDD1.n55 B 0.010969f
C219 VDD1.n56 B 0.011614f
C220 VDD1.n57 B 0.025926f
C221 VDD1.n58 B 0.025926f
C222 VDD1.n59 B 0.011614f
C223 VDD1.n60 B 0.010969f
C224 VDD1.n61 B 0.020413f
C225 VDD1.n62 B 0.020413f
C226 VDD1.n63 B 0.010969f
C227 VDD1.n64 B 0.011614f
C228 VDD1.n65 B 0.025926f
C229 VDD1.n66 B 0.052303f
C230 VDD1.n67 B 0.011614f
C231 VDD1.n68 B 0.021448f
C232 VDD1.n69 B 0.049693f
C233 VDD1.n70 B 0.068938f
C234 VDD1.n71 B 0.02715f
C235 VDD1.n72 B 0.020413f
C236 VDD1.n73 B 0.010969f
C237 VDD1.n74 B 0.025926f
C238 VDD1.n75 B 0.011614f
C239 VDD1.n76 B 0.020413f
C240 VDD1.n77 B 0.010969f
C241 VDD1.n78 B 0.025926f
C242 VDD1.n79 B 0.011614f
C243 VDD1.n80 B 0.020413f
C244 VDD1.n81 B 0.010969f
C245 VDD1.n82 B 0.025926f
C246 VDD1.n83 B 0.011614f
C247 VDD1.n84 B 0.020413f
C248 VDD1.n85 B 0.010969f
C249 VDD1.n86 B 0.025926f
C250 VDD1.n87 B 0.011614f
C251 VDD1.n88 B 0.020413f
C252 VDD1.n89 B 0.010969f
C253 VDD1.n90 B 0.025926f
C254 VDD1.n91 B 0.011614f
C255 VDD1.n92 B 1.1681f
C256 VDD1.n93 B 0.010969f
C257 VDD1.t1 B 0.04263f
C258 VDD1.n94 B 0.124384f
C259 VDD1.n95 B 0.015316f
C260 VDD1.n96 B 0.019445f
C261 VDD1.n97 B 0.025926f
C262 VDD1.n98 B 0.011614f
C263 VDD1.n99 B 0.010969f
C264 VDD1.n100 B 0.020413f
C265 VDD1.n101 B 0.020413f
C266 VDD1.n102 B 0.010969f
C267 VDD1.n103 B 0.011614f
C268 VDD1.n104 B 0.025926f
C269 VDD1.n105 B 0.025926f
C270 VDD1.n106 B 0.011614f
C271 VDD1.n107 B 0.010969f
C272 VDD1.n108 B 0.020413f
C273 VDD1.n109 B 0.020413f
C274 VDD1.n110 B 0.010969f
C275 VDD1.n111 B 0.011614f
C276 VDD1.n112 B 0.025926f
C277 VDD1.n113 B 0.025926f
C278 VDD1.n114 B 0.011614f
C279 VDD1.n115 B 0.010969f
C280 VDD1.n116 B 0.020413f
C281 VDD1.n117 B 0.020413f
C282 VDD1.n118 B 0.010969f
C283 VDD1.n119 B 0.011614f
C284 VDD1.n120 B 0.025926f
C285 VDD1.n121 B 0.025926f
C286 VDD1.n122 B 0.011614f
C287 VDD1.n123 B 0.010969f
C288 VDD1.n124 B 0.020413f
C289 VDD1.n125 B 0.020413f
C290 VDD1.n126 B 0.010969f
C291 VDD1.n127 B 0.011614f
C292 VDD1.n128 B 0.025926f
C293 VDD1.n129 B 0.025926f
C294 VDD1.n130 B 0.011614f
C295 VDD1.n131 B 0.010969f
C296 VDD1.n132 B 0.020413f
C297 VDD1.n133 B 0.020413f
C298 VDD1.n134 B 0.010969f
C299 VDD1.n135 B 0.011614f
C300 VDD1.n136 B 0.025926f
C301 VDD1.n137 B 0.052303f
C302 VDD1.n138 B 0.011614f
C303 VDD1.n139 B 0.021448f
C304 VDD1.n140 B 0.049693f
C305 VDD1.n141 B 0.764773f
C306 VTAIL.n0 B 0.02776f
C307 VTAIL.n1 B 0.020871f
C308 VTAIL.n2 B 0.011215f
C309 VTAIL.n3 B 0.026509f
C310 VTAIL.n4 B 0.011875f
C311 VTAIL.n5 B 0.020871f
C312 VTAIL.n6 B 0.011215f
C313 VTAIL.n7 B 0.026509f
C314 VTAIL.n8 B 0.011875f
C315 VTAIL.n9 B 0.020871f
C316 VTAIL.n10 B 0.011215f
C317 VTAIL.n11 B 0.026509f
C318 VTAIL.n12 B 0.011875f
C319 VTAIL.n13 B 0.020871f
C320 VTAIL.n14 B 0.011215f
C321 VTAIL.n15 B 0.026509f
C322 VTAIL.n16 B 0.011875f
C323 VTAIL.n17 B 0.020871f
C324 VTAIL.n18 B 0.011215f
C325 VTAIL.n19 B 0.026509f
C326 VTAIL.n20 B 0.011875f
C327 VTAIL.n21 B 1.19435f
C328 VTAIL.n22 B 0.011215f
C329 VTAIL.t3 B 0.043588f
C330 VTAIL.n23 B 0.127178f
C331 VTAIL.n24 B 0.01566f
C332 VTAIL.n25 B 0.019882f
C333 VTAIL.n26 B 0.026509f
C334 VTAIL.n27 B 0.011875f
C335 VTAIL.n28 B 0.011215f
C336 VTAIL.n29 B 0.020871f
C337 VTAIL.n30 B 0.020871f
C338 VTAIL.n31 B 0.011215f
C339 VTAIL.n32 B 0.011875f
C340 VTAIL.n33 B 0.026509f
C341 VTAIL.n34 B 0.026509f
C342 VTAIL.n35 B 0.011875f
C343 VTAIL.n36 B 0.011215f
C344 VTAIL.n37 B 0.020871f
C345 VTAIL.n38 B 0.020871f
C346 VTAIL.n39 B 0.011215f
C347 VTAIL.n40 B 0.011875f
C348 VTAIL.n41 B 0.026509f
C349 VTAIL.n42 B 0.026509f
C350 VTAIL.n43 B 0.011875f
C351 VTAIL.n44 B 0.011215f
C352 VTAIL.n45 B 0.020871f
C353 VTAIL.n46 B 0.020871f
C354 VTAIL.n47 B 0.011215f
C355 VTAIL.n48 B 0.011875f
C356 VTAIL.n49 B 0.026509f
C357 VTAIL.n50 B 0.026509f
C358 VTAIL.n51 B 0.011875f
C359 VTAIL.n52 B 0.011215f
C360 VTAIL.n53 B 0.020871f
C361 VTAIL.n54 B 0.020871f
C362 VTAIL.n55 B 0.011215f
C363 VTAIL.n56 B 0.011875f
C364 VTAIL.n57 B 0.026509f
C365 VTAIL.n58 B 0.026509f
C366 VTAIL.n59 B 0.011875f
C367 VTAIL.n60 B 0.011215f
C368 VTAIL.n61 B 0.020871f
C369 VTAIL.n62 B 0.020871f
C370 VTAIL.n63 B 0.011215f
C371 VTAIL.n64 B 0.011875f
C372 VTAIL.n65 B 0.026509f
C373 VTAIL.n66 B 0.053478f
C374 VTAIL.n67 B 0.011875f
C375 VTAIL.n68 B 0.02193f
C376 VTAIL.n69 B 0.050809f
C377 VTAIL.n70 B 0.054142f
C378 VTAIL.n71 B 1.65014f
C379 VTAIL.n72 B 0.02776f
C380 VTAIL.n73 B 0.020871f
C381 VTAIL.n74 B 0.011215f
C382 VTAIL.n75 B 0.026509f
C383 VTAIL.n76 B 0.011875f
C384 VTAIL.n77 B 0.020871f
C385 VTAIL.n78 B 0.011215f
C386 VTAIL.n79 B 0.026509f
C387 VTAIL.n80 B 0.011875f
C388 VTAIL.n81 B 0.020871f
C389 VTAIL.n82 B 0.011215f
C390 VTAIL.n83 B 0.026509f
C391 VTAIL.n84 B 0.011875f
C392 VTAIL.n85 B 0.020871f
C393 VTAIL.n86 B 0.011215f
C394 VTAIL.n87 B 0.026509f
C395 VTAIL.n88 B 0.011875f
C396 VTAIL.n89 B 0.020871f
C397 VTAIL.n90 B 0.011215f
C398 VTAIL.n91 B 0.026509f
C399 VTAIL.n92 B 0.011875f
C400 VTAIL.n93 B 1.19435f
C401 VTAIL.n94 B 0.011215f
C402 VTAIL.t0 B 0.043588f
C403 VTAIL.n95 B 0.127178f
C404 VTAIL.n96 B 0.01566f
C405 VTAIL.n97 B 0.019882f
C406 VTAIL.n98 B 0.026509f
C407 VTAIL.n99 B 0.011875f
C408 VTAIL.n100 B 0.011215f
C409 VTAIL.n101 B 0.020871f
C410 VTAIL.n102 B 0.020871f
C411 VTAIL.n103 B 0.011215f
C412 VTAIL.n104 B 0.011875f
C413 VTAIL.n105 B 0.026509f
C414 VTAIL.n106 B 0.026509f
C415 VTAIL.n107 B 0.011875f
C416 VTAIL.n108 B 0.011215f
C417 VTAIL.n109 B 0.020871f
C418 VTAIL.n110 B 0.020871f
C419 VTAIL.n111 B 0.011215f
C420 VTAIL.n112 B 0.011875f
C421 VTAIL.n113 B 0.026509f
C422 VTAIL.n114 B 0.026509f
C423 VTAIL.n115 B 0.011875f
C424 VTAIL.n116 B 0.011215f
C425 VTAIL.n117 B 0.020871f
C426 VTAIL.n118 B 0.020871f
C427 VTAIL.n119 B 0.011215f
C428 VTAIL.n120 B 0.011875f
C429 VTAIL.n121 B 0.026509f
C430 VTAIL.n122 B 0.026509f
C431 VTAIL.n123 B 0.011875f
C432 VTAIL.n124 B 0.011215f
C433 VTAIL.n125 B 0.020871f
C434 VTAIL.n126 B 0.020871f
C435 VTAIL.n127 B 0.011215f
C436 VTAIL.n128 B 0.011875f
C437 VTAIL.n129 B 0.026509f
C438 VTAIL.n130 B 0.026509f
C439 VTAIL.n131 B 0.011875f
C440 VTAIL.n132 B 0.011215f
C441 VTAIL.n133 B 0.020871f
C442 VTAIL.n134 B 0.020871f
C443 VTAIL.n135 B 0.011215f
C444 VTAIL.n136 B 0.011875f
C445 VTAIL.n137 B 0.026509f
C446 VTAIL.n138 B 0.053478f
C447 VTAIL.n139 B 0.011875f
C448 VTAIL.n140 B 0.02193f
C449 VTAIL.n141 B 0.050809f
C450 VTAIL.n142 B 0.054142f
C451 VTAIL.n143 B 1.70638f
C452 VTAIL.n144 B 0.02776f
C453 VTAIL.n145 B 0.020871f
C454 VTAIL.n146 B 0.011215f
C455 VTAIL.n147 B 0.026509f
C456 VTAIL.n148 B 0.011875f
C457 VTAIL.n149 B 0.020871f
C458 VTAIL.n150 B 0.011215f
C459 VTAIL.n151 B 0.026509f
C460 VTAIL.n152 B 0.011875f
C461 VTAIL.n153 B 0.020871f
C462 VTAIL.n154 B 0.011215f
C463 VTAIL.n155 B 0.026509f
C464 VTAIL.n156 B 0.011875f
C465 VTAIL.n157 B 0.020871f
C466 VTAIL.n158 B 0.011215f
C467 VTAIL.n159 B 0.026509f
C468 VTAIL.n160 B 0.011875f
C469 VTAIL.n161 B 0.020871f
C470 VTAIL.n162 B 0.011215f
C471 VTAIL.n163 B 0.026509f
C472 VTAIL.n164 B 0.011875f
C473 VTAIL.n165 B 1.19435f
C474 VTAIL.n166 B 0.011215f
C475 VTAIL.t2 B 0.043588f
C476 VTAIL.n167 B 0.127178f
C477 VTAIL.n168 B 0.01566f
C478 VTAIL.n169 B 0.019882f
C479 VTAIL.n170 B 0.026509f
C480 VTAIL.n171 B 0.011875f
C481 VTAIL.n172 B 0.011215f
C482 VTAIL.n173 B 0.020871f
C483 VTAIL.n174 B 0.020871f
C484 VTAIL.n175 B 0.011215f
C485 VTAIL.n176 B 0.011875f
C486 VTAIL.n177 B 0.026509f
C487 VTAIL.n178 B 0.026509f
C488 VTAIL.n179 B 0.011875f
C489 VTAIL.n180 B 0.011215f
C490 VTAIL.n181 B 0.020871f
C491 VTAIL.n182 B 0.020871f
C492 VTAIL.n183 B 0.011215f
C493 VTAIL.n184 B 0.011875f
C494 VTAIL.n185 B 0.026509f
C495 VTAIL.n186 B 0.026509f
C496 VTAIL.n187 B 0.011875f
C497 VTAIL.n188 B 0.011215f
C498 VTAIL.n189 B 0.020871f
C499 VTAIL.n190 B 0.020871f
C500 VTAIL.n191 B 0.011215f
C501 VTAIL.n192 B 0.011875f
C502 VTAIL.n193 B 0.026509f
C503 VTAIL.n194 B 0.026509f
C504 VTAIL.n195 B 0.011875f
C505 VTAIL.n196 B 0.011215f
C506 VTAIL.n197 B 0.020871f
C507 VTAIL.n198 B 0.020871f
C508 VTAIL.n199 B 0.011215f
C509 VTAIL.n200 B 0.011875f
C510 VTAIL.n201 B 0.026509f
C511 VTAIL.n202 B 0.026509f
C512 VTAIL.n203 B 0.011875f
C513 VTAIL.n204 B 0.011215f
C514 VTAIL.n205 B 0.020871f
C515 VTAIL.n206 B 0.020871f
C516 VTAIL.n207 B 0.011215f
C517 VTAIL.n208 B 0.011875f
C518 VTAIL.n209 B 0.026509f
C519 VTAIL.n210 B 0.053478f
C520 VTAIL.n211 B 0.011875f
C521 VTAIL.n212 B 0.02193f
C522 VTAIL.n213 B 0.050809f
C523 VTAIL.n214 B 0.054142f
C524 VTAIL.n215 B 1.46578f
C525 VTAIL.n216 B 0.02776f
C526 VTAIL.n217 B 0.020871f
C527 VTAIL.n218 B 0.011215f
C528 VTAIL.n219 B 0.026509f
C529 VTAIL.n220 B 0.011875f
C530 VTAIL.n221 B 0.020871f
C531 VTAIL.n222 B 0.011215f
C532 VTAIL.n223 B 0.026509f
C533 VTAIL.n224 B 0.011875f
C534 VTAIL.n225 B 0.020871f
C535 VTAIL.n226 B 0.011215f
C536 VTAIL.n227 B 0.026509f
C537 VTAIL.n228 B 0.011875f
C538 VTAIL.n229 B 0.020871f
C539 VTAIL.n230 B 0.011215f
C540 VTAIL.n231 B 0.026509f
C541 VTAIL.n232 B 0.011875f
C542 VTAIL.n233 B 0.020871f
C543 VTAIL.n234 B 0.011215f
C544 VTAIL.n235 B 0.026509f
C545 VTAIL.n236 B 0.011875f
C546 VTAIL.n237 B 1.19435f
C547 VTAIL.n238 B 0.011215f
C548 VTAIL.t1 B 0.043588f
C549 VTAIL.n239 B 0.127178f
C550 VTAIL.n240 B 0.01566f
C551 VTAIL.n241 B 0.019882f
C552 VTAIL.n242 B 0.026509f
C553 VTAIL.n243 B 0.011875f
C554 VTAIL.n244 B 0.011215f
C555 VTAIL.n245 B 0.020871f
C556 VTAIL.n246 B 0.020871f
C557 VTAIL.n247 B 0.011215f
C558 VTAIL.n248 B 0.011875f
C559 VTAIL.n249 B 0.026509f
C560 VTAIL.n250 B 0.026509f
C561 VTAIL.n251 B 0.011875f
C562 VTAIL.n252 B 0.011215f
C563 VTAIL.n253 B 0.020871f
C564 VTAIL.n254 B 0.020871f
C565 VTAIL.n255 B 0.011215f
C566 VTAIL.n256 B 0.011875f
C567 VTAIL.n257 B 0.026509f
C568 VTAIL.n258 B 0.026509f
C569 VTAIL.n259 B 0.011875f
C570 VTAIL.n260 B 0.011215f
C571 VTAIL.n261 B 0.020871f
C572 VTAIL.n262 B 0.020871f
C573 VTAIL.n263 B 0.011215f
C574 VTAIL.n264 B 0.011875f
C575 VTAIL.n265 B 0.026509f
C576 VTAIL.n266 B 0.026509f
C577 VTAIL.n267 B 0.011875f
C578 VTAIL.n268 B 0.011215f
C579 VTAIL.n269 B 0.020871f
C580 VTAIL.n270 B 0.020871f
C581 VTAIL.n271 B 0.011215f
C582 VTAIL.n272 B 0.011875f
C583 VTAIL.n273 B 0.026509f
C584 VTAIL.n274 B 0.026509f
C585 VTAIL.n275 B 0.011875f
C586 VTAIL.n276 B 0.011215f
C587 VTAIL.n277 B 0.020871f
C588 VTAIL.n278 B 0.020871f
C589 VTAIL.n279 B 0.011215f
C590 VTAIL.n280 B 0.011875f
C591 VTAIL.n281 B 0.026509f
C592 VTAIL.n282 B 0.053478f
C593 VTAIL.n283 B 0.011875f
C594 VTAIL.n284 B 0.02193f
C595 VTAIL.n285 B 0.050809f
C596 VTAIL.n286 B 0.054142f
C597 VTAIL.n287 B 1.37012f
C598 VP.t1 B 4.52566f
C599 VP.t0 B 3.79998f
C600 VP.n0 B 4.16974f
.ends

