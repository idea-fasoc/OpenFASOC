* NGSPICE file created from diff_pair_sample_0890.ext - technology: sky130A

.subckt diff_pair_sample_0890 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t1 VN.t0 VTAIL.t2 w_n2178_n2686# sky130_fd_pr__pfet_01v8 ad=3.3501 pd=17.96 as=3.3501 ps=17.96 w=8.59 l=2.69
X1 B.t11 B.t9 B.t10 w_n2178_n2686# sky130_fd_pr__pfet_01v8 ad=3.3501 pd=17.96 as=0 ps=0 w=8.59 l=2.69
X2 B.t8 B.t6 B.t7 w_n2178_n2686# sky130_fd_pr__pfet_01v8 ad=3.3501 pd=17.96 as=0 ps=0 w=8.59 l=2.69
X3 VDD1.t1 VP.t0 VTAIL.t1 w_n2178_n2686# sky130_fd_pr__pfet_01v8 ad=3.3501 pd=17.96 as=3.3501 ps=17.96 w=8.59 l=2.69
X4 VDD2.t0 VN.t1 VTAIL.t3 w_n2178_n2686# sky130_fd_pr__pfet_01v8 ad=3.3501 pd=17.96 as=3.3501 ps=17.96 w=8.59 l=2.69
X5 VDD1.t0 VP.t1 VTAIL.t0 w_n2178_n2686# sky130_fd_pr__pfet_01v8 ad=3.3501 pd=17.96 as=3.3501 ps=17.96 w=8.59 l=2.69
X6 B.t5 B.t3 B.t4 w_n2178_n2686# sky130_fd_pr__pfet_01v8 ad=3.3501 pd=17.96 as=0 ps=0 w=8.59 l=2.69
X7 B.t2 B.t0 B.t1 w_n2178_n2686# sky130_fd_pr__pfet_01v8 ad=3.3501 pd=17.96 as=0 ps=0 w=8.59 l=2.69
R0 VN VN.t1 160.369
R1 VN VN.t0 118.487
R2 VTAIL.n178 VTAIL.n138 756.745
R3 VTAIL.n40 VTAIL.n0 756.745
R4 VTAIL.n132 VTAIL.n92 756.745
R5 VTAIL.n86 VTAIL.n46 756.745
R6 VTAIL.n153 VTAIL.n152 585
R7 VTAIL.n150 VTAIL.n149 585
R8 VTAIL.n159 VTAIL.n158 585
R9 VTAIL.n161 VTAIL.n160 585
R10 VTAIL.n146 VTAIL.n145 585
R11 VTAIL.n167 VTAIL.n166 585
R12 VTAIL.n170 VTAIL.n169 585
R13 VTAIL.n168 VTAIL.n142 585
R14 VTAIL.n175 VTAIL.n141 585
R15 VTAIL.n177 VTAIL.n176 585
R16 VTAIL.n179 VTAIL.n178 585
R17 VTAIL.n15 VTAIL.n14 585
R18 VTAIL.n12 VTAIL.n11 585
R19 VTAIL.n21 VTAIL.n20 585
R20 VTAIL.n23 VTAIL.n22 585
R21 VTAIL.n8 VTAIL.n7 585
R22 VTAIL.n29 VTAIL.n28 585
R23 VTAIL.n32 VTAIL.n31 585
R24 VTAIL.n30 VTAIL.n4 585
R25 VTAIL.n37 VTAIL.n3 585
R26 VTAIL.n39 VTAIL.n38 585
R27 VTAIL.n41 VTAIL.n40 585
R28 VTAIL.n133 VTAIL.n132 585
R29 VTAIL.n131 VTAIL.n130 585
R30 VTAIL.n129 VTAIL.n95 585
R31 VTAIL.n99 VTAIL.n96 585
R32 VTAIL.n124 VTAIL.n123 585
R33 VTAIL.n122 VTAIL.n121 585
R34 VTAIL.n101 VTAIL.n100 585
R35 VTAIL.n116 VTAIL.n115 585
R36 VTAIL.n114 VTAIL.n113 585
R37 VTAIL.n105 VTAIL.n104 585
R38 VTAIL.n108 VTAIL.n107 585
R39 VTAIL.n87 VTAIL.n86 585
R40 VTAIL.n85 VTAIL.n84 585
R41 VTAIL.n83 VTAIL.n49 585
R42 VTAIL.n53 VTAIL.n50 585
R43 VTAIL.n78 VTAIL.n77 585
R44 VTAIL.n76 VTAIL.n75 585
R45 VTAIL.n55 VTAIL.n54 585
R46 VTAIL.n70 VTAIL.n69 585
R47 VTAIL.n68 VTAIL.n67 585
R48 VTAIL.n59 VTAIL.n58 585
R49 VTAIL.n62 VTAIL.n61 585
R50 VTAIL.t0 VTAIL.n106 329.039
R51 VTAIL.t3 VTAIL.n60 329.039
R52 VTAIL.t2 VTAIL.n151 329.038
R53 VTAIL.t1 VTAIL.n13 329.038
R54 VTAIL.n152 VTAIL.n149 171.744
R55 VTAIL.n159 VTAIL.n149 171.744
R56 VTAIL.n160 VTAIL.n159 171.744
R57 VTAIL.n160 VTAIL.n145 171.744
R58 VTAIL.n167 VTAIL.n145 171.744
R59 VTAIL.n169 VTAIL.n167 171.744
R60 VTAIL.n169 VTAIL.n168 171.744
R61 VTAIL.n168 VTAIL.n141 171.744
R62 VTAIL.n177 VTAIL.n141 171.744
R63 VTAIL.n178 VTAIL.n177 171.744
R64 VTAIL.n14 VTAIL.n11 171.744
R65 VTAIL.n21 VTAIL.n11 171.744
R66 VTAIL.n22 VTAIL.n21 171.744
R67 VTAIL.n22 VTAIL.n7 171.744
R68 VTAIL.n29 VTAIL.n7 171.744
R69 VTAIL.n31 VTAIL.n29 171.744
R70 VTAIL.n31 VTAIL.n30 171.744
R71 VTAIL.n30 VTAIL.n3 171.744
R72 VTAIL.n39 VTAIL.n3 171.744
R73 VTAIL.n40 VTAIL.n39 171.744
R74 VTAIL.n132 VTAIL.n131 171.744
R75 VTAIL.n131 VTAIL.n95 171.744
R76 VTAIL.n99 VTAIL.n95 171.744
R77 VTAIL.n123 VTAIL.n99 171.744
R78 VTAIL.n123 VTAIL.n122 171.744
R79 VTAIL.n122 VTAIL.n100 171.744
R80 VTAIL.n115 VTAIL.n100 171.744
R81 VTAIL.n115 VTAIL.n114 171.744
R82 VTAIL.n114 VTAIL.n104 171.744
R83 VTAIL.n107 VTAIL.n104 171.744
R84 VTAIL.n86 VTAIL.n85 171.744
R85 VTAIL.n85 VTAIL.n49 171.744
R86 VTAIL.n53 VTAIL.n49 171.744
R87 VTAIL.n77 VTAIL.n53 171.744
R88 VTAIL.n77 VTAIL.n76 171.744
R89 VTAIL.n76 VTAIL.n54 171.744
R90 VTAIL.n69 VTAIL.n54 171.744
R91 VTAIL.n69 VTAIL.n68 171.744
R92 VTAIL.n68 VTAIL.n58 171.744
R93 VTAIL.n61 VTAIL.n58 171.744
R94 VTAIL.n152 VTAIL.t2 85.8723
R95 VTAIL.n14 VTAIL.t1 85.8723
R96 VTAIL.n107 VTAIL.t0 85.8723
R97 VTAIL.n61 VTAIL.t3 85.8723
R98 VTAIL.n183 VTAIL.n182 33.5429
R99 VTAIL.n45 VTAIL.n44 33.5429
R100 VTAIL.n137 VTAIL.n136 33.5429
R101 VTAIL.n91 VTAIL.n90 33.5429
R102 VTAIL.n91 VTAIL.n45 24.9789
R103 VTAIL.n183 VTAIL.n137 22.3755
R104 VTAIL.n176 VTAIL.n175 13.1884
R105 VTAIL.n38 VTAIL.n37 13.1884
R106 VTAIL.n130 VTAIL.n129 13.1884
R107 VTAIL.n84 VTAIL.n83 13.1884
R108 VTAIL.n174 VTAIL.n142 12.8005
R109 VTAIL.n179 VTAIL.n140 12.8005
R110 VTAIL.n36 VTAIL.n4 12.8005
R111 VTAIL.n41 VTAIL.n2 12.8005
R112 VTAIL.n133 VTAIL.n94 12.8005
R113 VTAIL.n128 VTAIL.n96 12.8005
R114 VTAIL.n87 VTAIL.n48 12.8005
R115 VTAIL.n82 VTAIL.n50 12.8005
R116 VTAIL.n171 VTAIL.n170 12.0247
R117 VTAIL.n180 VTAIL.n138 12.0247
R118 VTAIL.n33 VTAIL.n32 12.0247
R119 VTAIL.n42 VTAIL.n0 12.0247
R120 VTAIL.n134 VTAIL.n92 12.0247
R121 VTAIL.n125 VTAIL.n124 12.0247
R122 VTAIL.n88 VTAIL.n46 12.0247
R123 VTAIL.n79 VTAIL.n78 12.0247
R124 VTAIL.n166 VTAIL.n144 11.249
R125 VTAIL.n28 VTAIL.n6 11.249
R126 VTAIL.n121 VTAIL.n98 11.249
R127 VTAIL.n75 VTAIL.n52 11.249
R128 VTAIL.n153 VTAIL.n151 10.7239
R129 VTAIL.n15 VTAIL.n13 10.7239
R130 VTAIL.n108 VTAIL.n106 10.7239
R131 VTAIL.n62 VTAIL.n60 10.7239
R132 VTAIL.n165 VTAIL.n146 10.4732
R133 VTAIL.n27 VTAIL.n8 10.4732
R134 VTAIL.n120 VTAIL.n101 10.4732
R135 VTAIL.n74 VTAIL.n55 10.4732
R136 VTAIL.n162 VTAIL.n161 9.69747
R137 VTAIL.n24 VTAIL.n23 9.69747
R138 VTAIL.n117 VTAIL.n116 9.69747
R139 VTAIL.n71 VTAIL.n70 9.69747
R140 VTAIL.n182 VTAIL.n181 9.45567
R141 VTAIL.n44 VTAIL.n43 9.45567
R142 VTAIL.n136 VTAIL.n135 9.45567
R143 VTAIL.n90 VTAIL.n89 9.45567
R144 VTAIL.n181 VTAIL.n180 9.3005
R145 VTAIL.n140 VTAIL.n139 9.3005
R146 VTAIL.n155 VTAIL.n154 9.3005
R147 VTAIL.n157 VTAIL.n156 9.3005
R148 VTAIL.n148 VTAIL.n147 9.3005
R149 VTAIL.n163 VTAIL.n162 9.3005
R150 VTAIL.n165 VTAIL.n164 9.3005
R151 VTAIL.n144 VTAIL.n143 9.3005
R152 VTAIL.n172 VTAIL.n171 9.3005
R153 VTAIL.n174 VTAIL.n173 9.3005
R154 VTAIL.n43 VTAIL.n42 9.3005
R155 VTAIL.n2 VTAIL.n1 9.3005
R156 VTAIL.n17 VTAIL.n16 9.3005
R157 VTAIL.n19 VTAIL.n18 9.3005
R158 VTAIL.n10 VTAIL.n9 9.3005
R159 VTAIL.n25 VTAIL.n24 9.3005
R160 VTAIL.n27 VTAIL.n26 9.3005
R161 VTAIL.n6 VTAIL.n5 9.3005
R162 VTAIL.n34 VTAIL.n33 9.3005
R163 VTAIL.n36 VTAIL.n35 9.3005
R164 VTAIL.n110 VTAIL.n109 9.3005
R165 VTAIL.n112 VTAIL.n111 9.3005
R166 VTAIL.n103 VTAIL.n102 9.3005
R167 VTAIL.n118 VTAIL.n117 9.3005
R168 VTAIL.n120 VTAIL.n119 9.3005
R169 VTAIL.n98 VTAIL.n97 9.3005
R170 VTAIL.n126 VTAIL.n125 9.3005
R171 VTAIL.n128 VTAIL.n127 9.3005
R172 VTAIL.n135 VTAIL.n134 9.3005
R173 VTAIL.n94 VTAIL.n93 9.3005
R174 VTAIL.n64 VTAIL.n63 9.3005
R175 VTAIL.n66 VTAIL.n65 9.3005
R176 VTAIL.n57 VTAIL.n56 9.3005
R177 VTAIL.n72 VTAIL.n71 9.3005
R178 VTAIL.n74 VTAIL.n73 9.3005
R179 VTAIL.n52 VTAIL.n51 9.3005
R180 VTAIL.n80 VTAIL.n79 9.3005
R181 VTAIL.n82 VTAIL.n81 9.3005
R182 VTAIL.n89 VTAIL.n88 9.3005
R183 VTAIL.n48 VTAIL.n47 9.3005
R184 VTAIL.n158 VTAIL.n148 8.92171
R185 VTAIL.n20 VTAIL.n10 8.92171
R186 VTAIL.n113 VTAIL.n103 8.92171
R187 VTAIL.n67 VTAIL.n57 8.92171
R188 VTAIL.n157 VTAIL.n150 8.14595
R189 VTAIL.n19 VTAIL.n12 8.14595
R190 VTAIL.n112 VTAIL.n105 8.14595
R191 VTAIL.n66 VTAIL.n59 8.14595
R192 VTAIL.n154 VTAIL.n153 7.3702
R193 VTAIL.n16 VTAIL.n15 7.3702
R194 VTAIL.n109 VTAIL.n108 7.3702
R195 VTAIL.n63 VTAIL.n62 7.3702
R196 VTAIL.n154 VTAIL.n150 5.81868
R197 VTAIL.n16 VTAIL.n12 5.81868
R198 VTAIL.n109 VTAIL.n105 5.81868
R199 VTAIL.n63 VTAIL.n59 5.81868
R200 VTAIL.n158 VTAIL.n157 5.04292
R201 VTAIL.n20 VTAIL.n19 5.04292
R202 VTAIL.n113 VTAIL.n112 5.04292
R203 VTAIL.n67 VTAIL.n66 5.04292
R204 VTAIL.n161 VTAIL.n148 4.26717
R205 VTAIL.n23 VTAIL.n10 4.26717
R206 VTAIL.n116 VTAIL.n103 4.26717
R207 VTAIL.n70 VTAIL.n57 4.26717
R208 VTAIL.n162 VTAIL.n146 3.49141
R209 VTAIL.n24 VTAIL.n8 3.49141
R210 VTAIL.n117 VTAIL.n101 3.49141
R211 VTAIL.n71 VTAIL.n55 3.49141
R212 VTAIL.n166 VTAIL.n165 2.71565
R213 VTAIL.n28 VTAIL.n27 2.71565
R214 VTAIL.n121 VTAIL.n120 2.71565
R215 VTAIL.n75 VTAIL.n74 2.71565
R216 VTAIL.n155 VTAIL.n151 2.41285
R217 VTAIL.n17 VTAIL.n13 2.41285
R218 VTAIL.n110 VTAIL.n106 2.41285
R219 VTAIL.n64 VTAIL.n60 2.41285
R220 VTAIL.n170 VTAIL.n144 1.93989
R221 VTAIL.n182 VTAIL.n138 1.93989
R222 VTAIL.n32 VTAIL.n6 1.93989
R223 VTAIL.n44 VTAIL.n0 1.93989
R224 VTAIL.n136 VTAIL.n92 1.93989
R225 VTAIL.n124 VTAIL.n98 1.93989
R226 VTAIL.n90 VTAIL.n46 1.93989
R227 VTAIL.n78 VTAIL.n52 1.93989
R228 VTAIL.n137 VTAIL.n91 1.77205
R229 VTAIL VTAIL.n45 1.17938
R230 VTAIL.n171 VTAIL.n142 1.16414
R231 VTAIL.n180 VTAIL.n179 1.16414
R232 VTAIL.n33 VTAIL.n4 1.16414
R233 VTAIL.n42 VTAIL.n41 1.16414
R234 VTAIL.n134 VTAIL.n133 1.16414
R235 VTAIL.n125 VTAIL.n96 1.16414
R236 VTAIL.n88 VTAIL.n87 1.16414
R237 VTAIL.n79 VTAIL.n50 1.16414
R238 VTAIL VTAIL.n183 0.593172
R239 VTAIL.n175 VTAIL.n174 0.388379
R240 VTAIL.n176 VTAIL.n140 0.388379
R241 VTAIL.n37 VTAIL.n36 0.388379
R242 VTAIL.n38 VTAIL.n2 0.388379
R243 VTAIL.n130 VTAIL.n94 0.388379
R244 VTAIL.n129 VTAIL.n128 0.388379
R245 VTAIL.n84 VTAIL.n48 0.388379
R246 VTAIL.n83 VTAIL.n82 0.388379
R247 VTAIL.n156 VTAIL.n155 0.155672
R248 VTAIL.n156 VTAIL.n147 0.155672
R249 VTAIL.n163 VTAIL.n147 0.155672
R250 VTAIL.n164 VTAIL.n163 0.155672
R251 VTAIL.n164 VTAIL.n143 0.155672
R252 VTAIL.n172 VTAIL.n143 0.155672
R253 VTAIL.n173 VTAIL.n172 0.155672
R254 VTAIL.n173 VTAIL.n139 0.155672
R255 VTAIL.n181 VTAIL.n139 0.155672
R256 VTAIL.n18 VTAIL.n17 0.155672
R257 VTAIL.n18 VTAIL.n9 0.155672
R258 VTAIL.n25 VTAIL.n9 0.155672
R259 VTAIL.n26 VTAIL.n25 0.155672
R260 VTAIL.n26 VTAIL.n5 0.155672
R261 VTAIL.n34 VTAIL.n5 0.155672
R262 VTAIL.n35 VTAIL.n34 0.155672
R263 VTAIL.n35 VTAIL.n1 0.155672
R264 VTAIL.n43 VTAIL.n1 0.155672
R265 VTAIL.n135 VTAIL.n93 0.155672
R266 VTAIL.n127 VTAIL.n93 0.155672
R267 VTAIL.n127 VTAIL.n126 0.155672
R268 VTAIL.n126 VTAIL.n97 0.155672
R269 VTAIL.n119 VTAIL.n97 0.155672
R270 VTAIL.n119 VTAIL.n118 0.155672
R271 VTAIL.n118 VTAIL.n102 0.155672
R272 VTAIL.n111 VTAIL.n102 0.155672
R273 VTAIL.n111 VTAIL.n110 0.155672
R274 VTAIL.n89 VTAIL.n47 0.155672
R275 VTAIL.n81 VTAIL.n47 0.155672
R276 VTAIL.n81 VTAIL.n80 0.155672
R277 VTAIL.n80 VTAIL.n51 0.155672
R278 VTAIL.n73 VTAIL.n51 0.155672
R279 VTAIL.n73 VTAIL.n72 0.155672
R280 VTAIL.n72 VTAIL.n56 0.155672
R281 VTAIL.n65 VTAIL.n56 0.155672
R282 VTAIL.n65 VTAIL.n64 0.155672
R283 VDD2.n85 VDD2.n45 756.745
R284 VDD2.n40 VDD2.n0 756.745
R285 VDD2.n86 VDD2.n85 585
R286 VDD2.n84 VDD2.n83 585
R287 VDD2.n82 VDD2.n48 585
R288 VDD2.n52 VDD2.n49 585
R289 VDD2.n77 VDD2.n76 585
R290 VDD2.n75 VDD2.n74 585
R291 VDD2.n54 VDD2.n53 585
R292 VDD2.n69 VDD2.n68 585
R293 VDD2.n67 VDD2.n66 585
R294 VDD2.n58 VDD2.n57 585
R295 VDD2.n61 VDD2.n60 585
R296 VDD2.n15 VDD2.n14 585
R297 VDD2.n12 VDD2.n11 585
R298 VDD2.n21 VDD2.n20 585
R299 VDD2.n23 VDD2.n22 585
R300 VDD2.n8 VDD2.n7 585
R301 VDD2.n29 VDD2.n28 585
R302 VDD2.n32 VDD2.n31 585
R303 VDD2.n30 VDD2.n4 585
R304 VDD2.n37 VDD2.n3 585
R305 VDD2.n39 VDD2.n38 585
R306 VDD2.n41 VDD2.n40 585
R307 VDD2.t0 VDD2.n59 329.039
R308 VDD2.t1 VDD2.n13 329.038
R309 VDD2.n85 VDD2.n84 171.744
R310 VDD2.n84 VDD2.n48 171.744
R311 VDD2.n52 VDD2.n48 171.744
R312 VDD2.n76 VDD2.n52 171.744
R313 VDD2.n76 VDD2.n75 171.744
R314 VDD2.n75 VDD2.n53 171.744
R315 VDD2.n68 VDD2.n53 171.744
R316 VDD2.n68 VDD2.n67 171.744
R317 VDD2.n67 VDD2.n57 171.744
R318 VDD2.n60 VDD2.n57 171.744
R319 VDD2.n14 VDD2.n11 171.744
R320 VDD2.n21 VDD2.n11 171.744
R321 VDD2.n22 VDD2.n21 171.744
R322 VDD2.n22 VDD2.n7 171.744
R323 VDD2.n29 VDD2.n7 171.744
R324 VDD2.n31 VDD2.n29 171.744
R325 VDD2.n31 VDD2.n30 171.744
R326 VDD2.n30 VDD2.n3 171.744
R327 VDD2.n39 VDD2.n3 171.744
R328 VDD2.n40 VDD2.n39 171.744
R329 VDD2.n90 VDD2.n44 86.4932
R330 VDD2.n60 VDD2.t0 85.8723
R331 VDD2.n14 VDD2.t1 85.8723
R332 VDD2.n90 VDD2.n89 50.2217
R333 VDD2.n83 VDD2.n82 13.1884
R334 VDD2.n38 VDD2.n37 13.1884
R335 VDD2.n86 VDD2.n47 12.8005
R336 VDD2.n81 VDD2.n49 12.8005
R337 VDD2.n36 VDD2.n4 12.8005
R338 VDD2.n41 VDD2.n2 12.8005
R339 VDD2.n87 VDD2.n45 12.0247
R340 VDD2.n78 VDD2.n77 12.0247
R341 VDD2.n33 VDD2.n32 12.0247
R342 VDD2.n42 VDD2.n0 12.0247
R343 VDD2.n74 VDD2.n51 11.249
R344 VDD2.n28 VDD2.n6 11.249
R345 VDD2.n61 VDD2.n59 10.7239
R346 VDD2.n15 VDD2.n13 10.7239
R347 VDD2.n73 VDD2.n54 10.4732
R348 VDD2.n27 VDD2.n8 10.4732
R349 VDD2.n70 VDD2.n69 9.69747
R350 VDD2.n24 VDD2.n23 9.69747
R351 VDD2.n89 VDD2.n88 9.45567
R352 VDD2.n44 VDD2.n43 9.45567
R353 VDD2.n63 VDD2.n62 9.3005
R354 VDD2.n65 VDD2.n64 9.3005
R355 VDD2.n56 VDD2.n55 9.3005
R356 VDD2.n71 VDD2.n70 9.3005
R357 VDD2.n73 VDD2.n72 9.3005
R358 VDD2.n51 VDD2.n50 9.3005
R359 VDD2.n79 VDD2.n78 9.3005
R360 VDD2.n81 VDD2.n80 9.3005
R361 VDD2.n88 VDD2.n87 9.3005
R362 VDD2.n47 VDD2.n46 9.3005
R363 VDD2.n43 VDD2.n42 9.3005
R364 VDD2.n2 VDD2.n1 9.3005
R365 VDD2.n17 VDD2.n16 9.3005
R366 VDD2.n19 VDD2.n18 9.3005
R367 VDD2.n10 VDD2.n9 9.3005
R368 VDD2.n25 VDD2.n24 9.3005
R369 VDD2.n27 VDD2.n26 9.3005
R370 VDD2.n6 VDD2.n5 9.3005
R371 VDD2.n34 VDD2.n33 9.3005
R372 VDD2.n36 VDD2.n35 9.3005
R373 VDD2.n66 VDD2.n56 8.92171
R374 VDD2.n20 VDD2.n10 8.92171
R375 VDD2.n65 VDD2.n58 8.14595
R376 VDD2.n19 VDD2.n12 8.14595
R377 VDD2.n62 VDD2.n61 7.3702
R378 VDD2.n16 VDD2.n15 7.3702
R379 VDD2.n62 VDD2.n58 5.81868
R380 VDD2.n16 VDD2.n12 5.81868
R381 VDD2.n66 VDD2.n65 5.04292
R382 VDD2.n20 VDD2.n19 5.04292
R383 VDD2.n69 VDD2.n56 4.26717
R384 VDD2.n23 VDD2.n10 4.26717
R385 VDD2.n70 VDD2.n54 3.49141
R386 VDD2.n24 VDD2.n8 3.49141
R387 VDD2.n74 VDD2.n73 2.71565
R388 VDD2.n28 VDD2.n27 2.71565
R389 VDD2.n63 VDD2.n59 2.41285
R390 VDD2.n17 VDD2.n13 2.41285
R391 VDD2.n89 VDD2.n45 1.93989
R392 VDD2.n77 VDD2.n51 1.93989
R393 VDD2.n32 VDD2.n6 1.93989
R394 VDD2.n44 VDD2.n0 1.93989
R395 VDD2.n87 VDD2.n86 1.16414
R396 VDD2.n78 VDD2.n49 1.16414
R397 VDD2.n33 VDD2.n4 1.16414
R398 VDD2.n42 VDD2.n41 1.16414
R399 VDD2 VDD2.n90 0.709552
R400 VDD2.n83 VDD2.n47 0.388379
R401 VDD2.n82 VDD2.n81 0.388379
R402 VDD2.n37 VDD2.n36 0.388379
R403 VDD2.n38 VDD2.n2 0.388379
R404 VDD2.n88 VDD2.n46 0.155672
R405 VDD2.n80 VDD2.n46 0.155672
R406 VDD2.n80 VDD2.n79 0.155672
R407 VDD2.n79 VDD2.n50 0.155672
R408 VDD2.n72 VDD2.n50 0.155672
R409 VDD2.n72 VDD2.n71 0.155672
R410 VDD2.n71 VDD2.n55 0.155672
R411 VDD2.n64 VDD2.n55 0.155672
R412 VDD2.n64 VDD2.n63 0.155672
R413 VDD2.n18 VDD2.n17 0.155672
R414 VDD2.n18 VDD2.n9 0.155672
R415 VDD2.n25 VDD2.n9 0.155672
R416 VDD2.n26 VDD2.n25 0.155672
R417 VDD2.n26 VDD2.n5 0.155672
R418 VDD2.n34 VDD2.n5 0.155672
R419 VDD2.n35 VDD2.n34 0.155672
R420 VDD2.n35 VDD2.n1 0.155672
R421 VDD2.n43 VDD2.n1 0.155672
R422 B.n364 B.n55 585
R423 B.n366 B.n365 585
R424 B.n367 B.n54 585
R425 B.n369 B.n368 585
R426 B.n370 B.n53 585
R427 B.n372 B.n371 585
R428 B.n373 B.n52 585
R429 B.n375 B.n374 585
R430 B.n376 B.n51 585
R431 B.n378 B.n377 585
R432 B.n379 B.n50 585
R433 B.n381 B.n380 585
R434 B.n382 B.n49 585
R435 B.n384 B.n383 585
R436 B.n385 B.n48 585
R437 B.n387 B.n386 585
R438 B.n388 B.n47 585
R439 B.n390 B.n389 585
R440 B.n391 B.n46 585
R441 B.n393 B.n392 585
R442 B.n394 B.n45 585
R443 B.n396 B.n395 585
R444 B.n397 B.n44 585
R445 B.n399 B.n398 585
R446 B.n400 B.n43 585
R447 B.n402 B.n401 585
R448 B.n403 B.n42 585
R449 B.n405 B.n404 585
R450 B.n406 B.n41 585
R451 B.n408 B.n407 585
R452 B.n409 B.n40 585
R453 B.n411 B.n410 585
R454 B.n413 B.n37 585
R455 B.n415 B.n414 585
R456 B.n416 B.n36 585
R457 B.n418 B.n417 585
R458 B.n419 B.n35 585
R459 B.n421 B.n420 585
R460 B.n422 B.n34 585
R461 B.n424 B.n423 585
R462 B.n425 B.n31 585
R463 B.n428 B.n427 585
R464 B.n429 B.n30 585
R465 B.n431 B.n430 585
R466 B.n432 B.n29 585
R467 B.n434 B.n433 585
R468 B.n435 B.n28 585
R469 B.n437 B.n436 585
R470 B.n438 B.n27 585
R471 B.n440 B.n439 585
R472 B.n441 B.n26 585
R473 B.n443 B.n442 585
R474 B.n444 B.n25 585
R475 B.n446 B.n445 585
R476 B.n447 B.n24 585
R477 B.n449 B.n448 585
R478 B.n450 B.n23 585
R479 B.n452 B.n451 585
R480 B.n453 B.n22 585
R481 B.n455 B.n454 585
R482 B.n456 B.n21 585
R483 B.n458 B.n457 585
R484 B.n459 B.n20 585
R485 B.n461 B.n460 585
R486 B.n462 B.n19 585
R487 B.n464 B.n463 585
R488 B.n465 B.n18 585
R489 B.n467 B.n466 585
R490 B.n468 B.n17 585
R491 B.n470 B.n469 585
R492 B.n471 B.n16 585
R493 B.n473 B.n472 585
R494 B.n474 B.n15 585
R495 B.n363 B.n362 585
R496 B.n361 B.n56 585
R497 B.n360 B.n359 585
R498 B.n358 B.n57 585
R499 B.n357 B.n356 585
R500 B.n355 B.n58 585
R501 B.n354 B.n353 585
R502 B.n352 B.n59 585
R503 B.n351 B.n350 585
R504 B.n349 B.n60 585
R505 B.n348 B.n347 585
R506 B.n346 B.n61 585
R507 B.n345 B.n344 585
R508 B.n343 B.n62 585
R509 B.n342 B.n341 585
R510 B.n340 B.n63 585
R511 B.n339 B.n338 585
R512 B.n337 B.n64 585
R513 B.n336 B.n335 585
R514 B.n334 B.n65 585
R515 B.n333 B.n332 585
R516 B.n331 B.n66 585
R517 B.n330 B.n329 585
R518 B.n328 B.n67 585
R519 B.n327 B.n326 585
R520 B.n325 B.n68 585
R521 B.n324 B.n323 585
R522 B.n322 B.n69 585
R523 B.n321 B.n320 585
R524 B.n319 B.n70 585
R525 B.n318 B.n317 585
R526 B.n316 B.n71 585
R527 B.n315 B.n314 585
R528 B.n313 B.n72 585
R529 B.n312 B.n311 585
R530 B.n310 B.n73 585
R531 B.n309 B.n308 585
R532 B.n307 B.n74 585
R533 B.n306 B.n305 585
R534 B.n304 B.n75 585
R535 B.n303 B.n302 585
R536 B.n301 B.n76 585
R537 B.n300 B.n299 585
R538 B.n298 B.n77 585
R539 B.n297 B.n296 585
R540 B.n295 B.n78 585
R541 B.n294 B.n293 585
R542 B.n292 B.n79 585
R543 B.n291 B.n290 585
R544 B.n289 B.n80 585
R545 B.n288 B.n287 585
R546 B.n286 B.n81 585
R547 B.n285 B.n284 585
R548 B.n174 B.n173 585
R549 B.n175 B.n122 585
R550 B.n177 B.n176 585
R551 B.n178 B.n121 585
R552 B.n180 B.n179 585
R553 B.n181 B.n120 585
R554 B.n183 B.n182 585
R555 B.n184 B.n119 585
R556 B.n186 B.n185 585
R557 B.n187 B.n118 585
R558 B.n189 B.n188 585
R559 B.n190 B.n117 585
R560 B.n192 B.n191 585
R561 B.n193 B.n116 585
R562 B.n195 B.n194 585
R563 B.n196 B.n115 585
R564 B.n198 B.n197 585
R565 B.n199 B.n114 585
R566 B.n201 B.n200 585
R567 B.n202 B.n113 585
R568 B.n204 B.n203 585
R569 B.n205 B.n112 585
R570 B.n207 B.n206 585
R571 B.n208 B.n111 585
R572 B.n210 B.n209 585
R573 B.n211 B.n110 585
R574 B.n213 B.n212 585
R575 B.n214 B.n109 585
R576 B.n216 B.n215 585
R577 B.n217 B.n108 585
R578 B.n219 B.n218 585
R579 B.n220 B.n105 585
R580 B.n223 B.n222 585
R581 B.n224 B.n104 585
R582 B.n226 B.n225 585
R583 B.n227 B.n103 585
R584 B.n229 B.n228 585
R585 B.n230 B.n102 585
R586 B.n232 B.n231 585
R587 B.n233 B.n101 585
R588 B.n235 B.n234 585
R589 B.n237 B.n236 585
R590 B.n238 B.n97 585
R591 B.n240 B.n239 585
R592 B.n241 B.n96 585
R593 B.n243 B.n242 585
R594 B.n244 B.n95 585
R595 B.n246 B.n245 585
R596 B.n247 B.n94 585
R597 B.n249 B.n248 585
R598 B.n250 B.n93 585
R599 B.n252 B.n251 585
R600 B.n253 B.n92 585
R601 B.n255 B.n254 585
R602 B.n256 B.n91 585
R603 B.n258 B.n257 585
R604 B.n259 B.n90 585
R605 B.n261 B.n260 585
R606 B.n262 B.n89 585
R607 B.n264 B.n263 585
R608 B.n265 B.n88 585
R609 B.n267 B.n266 585
R610 B.n268 B.n87 585
R611 B.n270 B.n269 585
R612 B.n271 B.n86 585
R613 B.n273 B.n272 585
R614 B.n274 B.n85 585
R615 B.n276 B.n275 585
R616 B.n277 B.n84 585
R617 B.n279 B.n278 585
R618 B.n280 B.n83 585
R619 B.n282 B.n281 585
R620 B.n283 B.n82 585
R621 B.n172 B.n123 585
R622 B.n171 B.n170 585
R623 B.n169 B.n124 585
R624 B.n168 B.n167 585
R625 B.n166 B.n125 585
R626 B.n165 B.n164 585
R627 B.n163 B.n126 585
R628 B.n162 B.n161 585
R629 B.n160 B.n127 585
R630 B.n159 B.n158 585
R631 B.n157 B.n128 585
R632 B.n156 B.n155 585
R633 B.n154 B.n129 585
R634 B.n153 B.n152 585
R635 B.n151 B.n130 585
R636 B.n150 B.n149 585
R637 B.n148 B.n131 585
R638 B.n147 B.n146 585
R639 B.n145 B.n132 585
R640 B.n144 B.n143 585
R641 B.n142 B.n133 585
R642 B.n141 B.n140 585
R643 B.n139 B.n134 585
R644 B.n138 B.n137 585
R645 B.n136 B.n135 585
R646 B.n2 B.n0 585
R647 B.n513 B.n1 585
R648 B.n512 B.n511 585
R649 B.n510 B.n3 585
R650 B.n509 B.n508 585
R651 B.n507 B.n4 585
R652 B.n506 B.n505 585
R653 B.n504 B.n5 585
R654 B.n503 B.n502 585
R655 B.n501 B.n6 585
R656 B.n500 B.n499 585
R657 B.n498 B.n7 585
R658 B.n497 B.n496 585
R659 B.n495 B.n8 585
R660 B.n494 B.n493 585
R661 B.n492 B.n9 585
R662 B.n491 B.n490 585
R663 B.n489 B.n10 585
R664 B.n488 B.n487 585
R665 B.n486 B.n11 585
R666 B.n485 B.n484 585
R667 B.n483 B.n12 585
R668 B.n482 B.n481 585
R669 B.n480 B.n13 585
R670 B.n479 B.n478 585
R671 B.n477 B.n14 585
R672 B.n476 B.n475 585
R673 B.n515 B.n514 585
R674 B.n174 B.n123 458.866
R675 B.n476 B.n15 458.866
R676 B.n284 B.n283 458.866
R677 B.n362 B.n55 458.866
R678 B.n98 B.t5 372.719
R679 B.n38 B.t7 372.719
R680 B.n106 B.t2 372.719
R681 B.n32 B.t10 372.719
R682 B.n99 B.t4 314.149
R683 B.n39 B.t8 314.149
R684 B.n107 B.t1 314.149
R685 B.n33 B.t11 314.149
R686 B.n98 B.t3 285.137
R687 B.n106 B.t0 285.137
R688 B.n32 B.t9 285.137
R689 B.n38 B.t6 285.137
R690 B.n170 B.n123 163.367
R691 B.n170 B.n169 163.367
R692 B.n169 B.n168 163.367
R693 B.n168 B.n125 163.367
R694 B.n164 B.n125 163.367
R695 B.n164 B.n163 163.367
R696 B.n163 B.n162 163.367
R697 B.n162 B.n127 163.367
R698 B.n158 B.n127 163.367
R699 B.n158 B.n157 163.367
R700 B.n157 B.n156 163.367
R701 B.n156 B.n129 163.367
R702 B.n152 B.n129 163.367
R703 B.n152 B.n151 163.367
R704 B.n151 B.n150 163.367
R705 B.n150 B.n131 163.367
R706 B.n146 B.n131 163.367
R707 B.n146 B.n145 163.367
R708 B.n145 B.n144 163.367
R709 B.n144 B.n133 163.367
R710 B.n140 B.n133 163.367
R711 B.n140 B.n139 163.367
R712 B.n139 B.n138 163.367
R713 B.n138 B.n135 163.367
R714 B.n135 B.n2 163.367
R715 B.n514 B.n2 163.367
R716 B.n514 B.n513 163.367
R717 B.n513 B.n512 163.367
R718 B.n512 B.n3 163.367
R719 B.n508 B.n3 163.367
R720 B.n508 B.n507 163.367
R721 B.n507 B.n506 163.367
R722 B.n506 B.n5 163.367
R723 B.n502 B.n5 163.367
R724 B.n502 B.n501 163.367
R725 B.n501 B.n500 163.367
R726 B.n500 B.n7 163.367
R727 B.n496 B.n7 163.367
R728 B.n496 B.n495 163.367
R729 B.n495 B.n494 163.367
R730 B.n494 B.n9 163.367
R731 B.n490 B.n9 163.367
R732 B.n490 B.n489 163.367
R733 B.n489 B.n488 163.367
R734 B.n488 B.n11 163.367
R735 B.n484 B.n11 163.367
R736 B.n484 B.n483 163.367
R737 B.n483 B.n482 163.367
R738 B.n482 B.n13 163.367
R739 B.n478 B.n13 163.367
R740 B.n478 B.n477 163.367
R741 B.n477 B.n476 163.367
R742 B.n175 B.n174 163.367
R743 B.n176 B.n175 163.367
R744 B.n176 B.n121 163.367
R745 B.n180 B.n121 163.367
R746 B.n181 B.n180 163.367
R747 B.n182 B.n181 163.367
R748 B.n182 B.n119 163.367
R749 B.n186 B.n119 163.367
R750 B.n187 B.n186 163.367
R751 B.n188 B.n187 163.367
R752 B.n188 B.n117 163.367
R753 B.n192 B.n117 163.367
R754 B.n193 B.n192 163.367
R755 B.n194 B.n193 163.367
R756 B.n194 B.n115 163.367
R757 B.n198 B.n115 163.367
R758 B.n199 B.n198 163.367
R759 B.n200 B.n199 163.367
R760 B.n200 B.n113 163.367
R761 B.n204 B.n113 163.367
R762 B.n205 B.n204 163.367
R763 B.n206 B.n205 163.367
R764 B.n206 B.n111 163.367
R765 B.n210 B.n111 163.367
R766 B.n211 B.n210 163.367
R767 B.n212 B.n211 163.367
R768 B.n212 B.n109 163.367
R769 B.n216 B.n109 163.367
R770 B.n217 B.n216 163.367
R771 B.n218 B.n217 163.367
R772 B.n218 B.n105 163.367
R773 B.n223 B.n105 163.367
R774 B.n224 B.n223 163.367
R775 B.n225 B.n224 163.367
R776 B.n225 B.n103 163.367
R777 B.n229 B.n103 163.367
R778 B.n230 B.n229 163.367
R779 B.n231 B.n230 163.367
R780 B.n231 B.n101 163.367
R781 B.n235 B.n101 163.367
R782 B.n236 B.n235 163.367
R783 B.n236 B.n97 163.367
R784 B.n240 B.n97 163.367
R785 B.n241 B.n240 163.367
R786 B.n242 B.n241 163.367
R787 B.n242 B.n95 163.367
R788 B.n246 B.n95 163.367
R789 B.n247 B.n246 163.367
R790 B.n248 B.n247 163.367
R791 B.n248 B.n93 163.367
R792 B.n252 B.n93 163.367
R793 B.n253 B.n252 163.367
R794 B.n254 B.n253 163.367
R795 B.n254 B.n91 163.367
R796 B.n258 B.n91 163.367
R797 B.n259 B.n258 163.367
R798 B.n260 B.n259 163.367
R799 B.n260 B.n89 163.367
R800 B.n264 B.n89 163.367
R801 B.n265 B.n264 163.367
R802 B.n266 B.n265 163.367
R803 B.n266 B.n87 163.367
R804 B.n270 B.n87 163.367
R805 B.n271 B.n270 163.367
R806 B.n272 B.n271 163.367
R807 B.n272 B.n85 163.367
R808 B.n276 B.n85 163.367
R809 B.n277 B.n276 163.367
R810 B.n278 B.n277 163.367
R811 B.n278 B.n83 163.367
R812 B.n282 B.n83 163.367
R813 B.n283 B.n282 163.367
R814 B.n284 B.n81 163.367
R815 B.n288 B.n81 163.367
R816 B.n289 B.n288 163.367
R817 B.n290 B.n289 163.367
R818 B.n290 B.n79 163.367
R819 B.n294 B.n79 163.367
R820 B.n295 B.n294 163.367
R821 B.n296 B.n295 163.367
R822 B.n296 B.n77 163.367
R823 B.n300 B.n77 163.367
R824 B.n301 B.n300 163.367
R825 B.n302 B.n301 163.367
R826 B.n302 B.n75 163.367
R827 B.n306 B.n75 163.367
R828 B.n307 B.n306 163.367
R829 B.n308 B.n307 163.367
R830 B.n308 B.n73 163.367
R831 B.n312 B.n73 163.367
R832 B.n313 B.n312 163.367
R833 B.n314 B.n313 163.367
R834 B.n314 B.n71 163.367
R835 B.n318 B.n71 163.367
R836 B.n319 B.n318 163.367
R837 B.n320 B.n319 163.367
R838 B.n320 B.n69 163.367
R839 B.n324 B.n69 163.367
R840 B.n325 B.n324 163.367
R841 B.n326 B.n325 163.367
R842 B.n326 B.n67 163.367
R843 B.n330 B.n67 163.367
R844 B.n331 B.n330 163.367
R845 B.n332 B.n331 163.367
R846 B.n332 B.n65 163.367
R847 B.n336 B.n65 163.367
R848 B.n337 B.n336 163.367
R849 B.n338 B.n337 163.367
R850 B.n338 B.n63 163.367
R851 B.n342 B.n63 163.367
R852 B.n343 B.n342 163.367
R853 B.n344 B.n343 163.367
R854 B.n344 B.n61 163.367
R855 B.n348 B.n61 163.367
R856 B.n349 B.n348 163.367
R857 B.n350 B.n349 163.367
R858 B.n350 B.n59 163.367
R859 B.n354 B.n59 163.367
R860 B.n355 B.n354 163.367
R861 B.n356 B.n355 163.367
R862 B.n356 B.n57 163.367
R863 B.n360 B.n57 163.367
R864 B.n361 B.n360 163.367
R865 B.n362 B.n361 163.367
R866 B.n472 B.n15 163.367
R867 B.n472 B.n471 163.367
R868 B.n471 B.n470 163.367
R869 B.n470 B.n17 163.367
R870 B.n466 B.n17 163.367
R871 B.n466 B.n465 163.367
R872 B.n465 B.n464 163.367
R873 B.n464 B.n19 163.367
R874 B.n460 B.n19 163.367
R875 B.n460 B.n459 163.367
R876 B.n459 B.n458 163.367
R877 B.n458 B.n21 163.367
R878 B.n454 B.n21 163.367
R879 B.n454 B.n453 163.367
R880 B.n453 B.n452 163.367
R881 B.n452 B.n23 163.367
R882 B.n448 B.n23 163.367
R883 B.n448 B.n447 163.367
R884 B.n447 B.n446 163.367
R885 B.n446 B.n25 163.367
R886 B.n442 B.n25 163.367
R887 B.n442 B.n441 163.367
R888 B.n441 B.n440 163.367
R889 B.n440 B.n27 163.367
R890 B.n436 B.n27 163.367
R891 B.n436 B.n435 163.367
R892 B.n435 B.n434 163.367
R893 B.n434 B.n29 163.367
R894 B.n430 B.n29 163.367
R895 B.n430 B.n429 163.367
R896 B.n429 B.n428 163.367
R897 B.n428 B.n31 163.367
R898 B.n423 B.n31 163.367
R899 B.n423 B.n422 163.367
R900 B.n422 B.n421 163.367
R901 B.n421 B.n35 163.367
R902 B.n417 B.n35 163.367
R903 B.n417 B.n416 163.367
R904 B.n416 B.n415 163.367
R905 B.n415 B.n37 163.367
R906 B.n410 B.n37 163.367
R907 B.n410 B.n409 163.367
R908 B.n409 B.n408 163.367
R909 B.n408 B.n41 163.367
R910 B.n404 B.n41 163.367
R911 B.n404 B.n403 163.367
R912 B.n403 B.n402 163.367
R913 B.n402 B.n43 163.367
R914 B.n398 B.n43 163.367
R915 B.n398 B.n397 163.367
R916 B.n397 B.n396 163.367
R917 B.n396 B.n45 163.367
R918 B.n392 B.n45 163.367
R919 B.n392 B.n391 163.367
R920 B.n391 B.n390 163.367
R921 B.n390 B.n47 163.367
R922 B.n386 B.n47 163.367
R923 B.n386 B.n385 163.367
R924 B.n385 B.n384 163.367
R925 B.n384 B.n49 163.367
R926 B.n380 B.n49 163.367
R927 B.n380 B.n379 163.367
R928 B.n379 B.n378 163.367
R929 B.n378 B.n51 163.367
R930 B.n374 B.n51 163.367
R931 B.n374 B.n373 163.367
R932 B.n373 B.n372 163.367
R933 B.n372 B.n53 163.367
R934 B.n368 B.n53 163.367
R935 B.n368 B.n367 163.367
R936 B.n367 B.n366 163.367
R937 B.n366 B.n55 163.367
R938 B.n100 B.n99 59.5399
R939 B.n221 B.n107 59.5399
R940 B.n426 B.n33 59.5399
R941 B.n412 B.n39 59.5399
R942 B.n99 B.n98 58.5702
R943 B.n107 B.n106 58.5702
R944 B.n33 B.n32 58.5702
R945 B.n39 B.n38 58.5702
R946 B.n475 B.n474 29.8151
R947 B.n364 B.n363 29.8151
R948 B.n285 B.n82 29.8151
R949 B.n173 B.n172 29.8151
R950 B B.n515 18.0485
R951 B.n474 B.n473 10.6151
R952 B.n473 B.n16 10.6151
R953 B.n469 B.n16 10.6151
R954 B.n469 B.n468 10.6151
R955 B.n468 B.n467 10.6151
R956 B.n467 B.n18 10.6151
R957 B.n463 B.n18 10.6151
R958 B.n463 B.n462 10.6151
R959 B.n462 B.n461 10.6151
R960 B.n461 B.n20 10.6151
R961 B.n457 B.n20 10.6151
R962 B.n457 B.n456 10.6151
R963 B.n456 B.n455 10.6151
R964 B.n455 B.n22 10.6151
R965 B.n451 B.n22 10.6151
R966 B.n451 B.n450 10.6151
R967 B.n450 B.n449 10.6151
R968 B.n449 B.n24 10.6151
R969 B.n445 B.n24 10.6151
R970 B.n445 B.n444 10.6151
R971 B.n444 B.n443 10.6151
R972 B.n443 B.n26 10.6151
R973 B.n439 B.n26 10.6151
R974 B.n439 B.n438 10.6151
R975 B.n438 B.n437 10.6151
R976 B.n437 B.n28 10.6151
R977 B.n433 B.n28 10.6151
R978 B.n433 B.n432 10.6151
R979 B.n432 B.n431 10.6151
R980 B.n431 B.n30 10.6151
R981 B.n427 B.n30 10.6151
R982 B.n425 B.n424 10.6151
R983 B.n424 B.n34 10.6151
R984 B.n420 B.n34 10.6151
R985 B.n420 B.n419 10.6151
R986 B.n419 B.n418 10.6151
R987 B.n418 B.n36 10.6151
R988 B.n414 B.n36 10.6151
R989 B.n414 B.n413 10.6151
R990 B.n411 B.n40 10.6151
R991 B.n407 B.n40 10.6151
R992 B.n407 B.n406 10.6151
R993 B.n406 B.n405 10.6151
R994 B.n405 B.n42 10.6151
R995 B.n401 B.n42 10.6151
R996 B.n401 B.n400 10.6151
R997 B.n400 B.n399 10.6151
R998 B.n399 B.n44 10.6151
R999 B.n395 B.n44 10.6151
R1000 B.n395 B.n394 10.6151
R1001 B.n394 B.n393 10.6151
R1002 B.n393 B.n46 10.6151
R1003 B.n389 B.n46 10.6151
R1004 B.n389 B.n388 10.6151
R1005 B.n388 B.n387 10.6151
R1006 B.n387 B.n48 10.6151
R1007 B.n383 B.n48 10.6151
R1008 B.n383 B.n382 10.6151
R1009 B.n382 B.n381 10.6151
R1010 B.n381 B.n50 10.6151
R1011 B.n377 B.n50 10.6151
R1012 B.n377 B.n376 10.6151
R1013 B.n376 B.n375 10.6151
R1014 B.n375 B.n52 10.6151
R1015 B.n371 B.n52 10.6151
R1016 B.n371 B.n370 10.6151
R1017 B.n370 B.n369 10.6151
R1018 B.n369 B.n54 10.6151
R1019 B.n365 B.n54 10.6151
R1020 B.n365 B.n364 10.6151
R1021 B.n286 B.n285 10.6151
R1022 B.n287 B.n286 10.6151
R1023 B.n287 B.n80 10.6151
R1024 B.n291 B.n80 10.6151
R1025 B.n292 B.n291 10.6151
R1026 B.n293 B.n292 10.6151
R1027 B.n293 B.n78 10.6151
R1028 B.n297 B.n78 10.6151
R1029 B.n298 B.n297 10.6151
R1030 B.n299 B.n298 10.6151
R1031 B.n299 B.n76 10.6151
R1032 B.n303 B.n76 10.6151
R1033 B.n304 B.n303 10.6151
R1034 B.n305 B.n304 10.6151
R1035 B.n305 B.n74 10.6151
R1036 B.n309 B.n74 10.6151
R1037 B.n310 B.n309 10.6151
R1038 B.n311 B.n310 10.6151
R1039 B.n311 B.n72 10.6151
R1040 B.n315 B.n72 10.6151
R1041 B.n316 B.n315 10.6151
R1042 B.n317 B.n316 10.6151
R1043 B.n317 B.n70 10.6151
R1044 B.n321 B.n70 10.6151
R1045 B.n322 B.n321 10.6151
R1046 B.n323 B.n322 10.6151
R1047 B.n323 B.n68 10.6151
R1048 B.n327 B.n68 10.6151
R1049 B.n328 B.n327 10.6151
R1050 B.n329 B.n328 10.6151
R1051 B.n329 B.n66 10.6151
R1052 B.n333 B.n66 10.6151
R1053 B.n334 B.n333 10.6151
R1054 B.n335 B.n334 10.6151
R1055 B.n335 B.n64 10.6151
R1056 B.n339 B.n64 10.6151
R1057 B.n340 B.n339 10.6151
R1058 B.n341 B.n340 10.6151
R1059 B.n341 B.n62 10.6151
R1060 B.n345 B.n62 10.6151
R1061 B.n346 B.n345 10.6151
R1062 B.n347 B.n346 10.6151
R1063 B.n347 B.n60 10.6151
R1064 B.n351 B.n60 10.6151
R1065 B.n352 B.n351 10.6151
R1066 B.n353 B.n352 10.6151
R1067 B.n353 B.n58 10.6151
R1068 B.n357 B.n58 10.6151
R1069 B.n358 B.n357 10.6151
R1070 B.n359 B.n358 10.6151
R1071 B.n359 B.n56 10.6151
R1072 B.n363 B.n56 10.6151
R1073 B.n173 B.n122 10.6151
R1074 B.n177 B.n122 10.6151
R1075 B.n178 B.n177 10.6151
R1076 B.n179 B.n178 10.6151
R1077 B.n179 B.n120 10.6151
R1078 B.n183 B.n120 10.6151
R1079 B.n184 B.n183 10.6151
R1080 B.n185 B.n184 10.6151
R1081 B.n185 B.n118 10.6151
R1082 B.n189 B.n118 10.6151
R1083 B.n190 B.n189 10.6151
R1084 B.n191 B.n190 10.6151
R1085 B.n191 B.n116 10.6151
R1086 B.n195 B.n116 10.6151
R1087 B.n196 B.n195 10.6151
R1088 B.n197 B.n196 10.6151
R1089 B.n197 B.n114 10.6151
R1090 B.n201 B.n114 10.6151
R1091 B.n202 B.n201 10.6151
R1092 B.n203 B.n202 10.6151
R1093 B.n203 B.n112 10.6151
R1094 B.n207 B.n112 10.6151
R1095 B.n208 B.n207 10.6151
R1096 B.n209 B.n208 10.6151
R1097 B.n209 B.n110 10.6151
R1098 B.n213 B.n110 10.6151
R1099 B.n214 B.n213 10.6151
R1100 B.n215 B.n214 10.6151
R1101 B.n215 B.n108 10.6151
R1102 B.n219 B.n108 10.6151
R1103 B.n220 B.n219 10.6151
R1104 B.n222 B.n104 10.6151
R1105 B.n226 B.n104 10.6151
R1106 B.n227 B.n226 10.6151
R1107 B.n228 B.n227 10.6151
R1108 B.n228 B.n102 10.6151
R1109 B.n232 B.n102 10.6151
R1110 B.n233 B.n232 10.6151
R1111 B.n234 B.n233 10.6151
R1112 B.n238 B.n237 10.6151
R1113 B.n239 B.n238 10.6151
R1114 B.n239 B.n96 10.6151
R1115 B.n243 B.n96 10.6151
R1116 B.n244 B.n243 10.6151
R1117 B.n245 B.n244 10.6151
R1118 B.n245 B.n94 10.6151
R1119 B.n249 B.n94 10.6151
R1120 B.n250 B.n249 10.6151
R1121 B.n251 B.n250 10.6151
R1122 B.n251 B.n92 10.6151
R1123 B.n255 B.n92 10.6151
R1124 B.n256 B.n255 10.6151
R1125 B.n257 B.n256 10.6151
R1126 B.n257 B.n90 10.6151
R1127 B.n261 B.n90 10.6151
R1128 B.n262 B.n261 10.6151
R1129 B.n263 B.n262 10.6151
R1130 B.n263 B.n88 10.6151
R1131 B.n267 B.n88 10.6151
R1132 B.n268 B.n267 10.6151
R1133 B.n269 B.n268 10.6151
R1134 B.n269 B.n86 10.6151
R1135 B.n273 B.n86 10.6151
R1136 B.n274 B.n273 10.6151
R1137 B.n275 B.n274 10.6151
R1138 B.n275 B.n84 10.6151
R1139 B.n279 B.n84 10.6151
R1140 B.n280 B.n279 10.6151
R1141 B.n281 B.n280 10.6151
R1142 B.n281 B.n82 10.6151
R1143 B.n172 B.n171 10.6151
R1144 B.n171 B.n124 10.6151
R1145 B.n167 B.n124 10.6151
R1146 B.n167 B.n166 10.6151
R1147 B.n166 B.n165 10.6151
R1148 B.n165 B.n126 10.6151
R1149 B.n161 B.n126 10.6151
R1150 B.n161 B.n160 10.6151
R1151 B.n160 B.n159 10.6151
R1152 B.n159 B.n128 10.6151
R1153 B.n155 B.n128 10.6151
R1154 B.n155 B.n154 10.6151
R1155 B.n154 B.n153 10.6151
R1156 B.n153 B.n130 10.6151
R1157 B.n149 B.n130 10.6151
R1158 B.n149 B.n148 10.6151
R1159 B.n148 B.n147 10.6151
R1160 B.n147 B.n132 10.6151
R1161 B.n143 B.n132 10.6151
R1162 B.n143 B.n142 10.6151
R1163 B.n142 B.n141 10.6151
R1164 B.n141 B.n134 10.6151
R1165 B.n137 B.n134 10.6151
R1166 B.n137 B.n136 10.6151
R1167 B.n136 B.n0 10.6151
R1168 B.n511 B.n1 10.6151
R1169 B.n511 B.n510 10.6151
R1170 B.n510 B.n509 10.6151
R1171 B.n509 B.n4 10.6151
R1172 B.n505 B.n4 10.6151
R1173 B.n505 B.n504 10.6151
R1174 B.n504 B.n503 10.6151
R1175 B.n503 B.n6 10.6151
R1176 B.n499 B.n6 10.6151
R1177 B.n499 B.n498 10.6151
R1178 B.n498 B.n497 10.6151
R1179 B.n497 B.n8 10.6151
R1180 B.n493 B.n8 10.6151
R1181 B.n493 B.n492 10.6151
R1182 B.n492 B.n491 10.6151
R1183 B.n491 B.n10 10.6151
R1184 B.n487 B.n10 10.6151
R1185 B.n487 B.n486 10.6151
R1186 B.n486 B.n485 10.6151
R1187 B.n485 B.n12 10.6151
R1188 B.n481 B.n12 10.6151
R1189 B.n481 B.n480 10.6151
R1190 B.n480 B.n479 10.6151
R1191 B.n479 B.n14 10.6151
R1192 B.n475 B.n14 10.6151
R1193 B.n426 B.n425 6.5566
R1194 B.n413 B.n412 6.5566
R1195 B.n222 B.n221 6.5566
R1196 B.n234 B.n100 6.5566
R1197 B.n427 B.n426 4.05904
R1198 B.n412 B.n411 4.05904
R1199 B.n221 B.n220 4.05904
R1200 B.n237 B.n100 4.05904
R1201 B.n515 B.n0 2.81026
R1202 B.n515 B.n1 2.81026
R1203 VP.n0 VP.t1 160.368
R1204 VP.n0 VP.t0 118.055
R1205 VP VP.n0 0.431811
R1206 VDD1.n40 VDD1.n0 756.745
R1207 VDD1.n85 VDD1.n45 756.745
R1208 VDD1.n41 VDD1.n40 585
R1209 VDD1.n39 VDD1.n38 585
R1210 VDD1.n37 VDD1.n3 585
R1211 VDD1.n7 VDD1.n4 585
R1212 VDD1.n32 VDD1.n31 585
R1213 VDD1.n30 VDD1.n29 585
R1214 VDD1.n9 VDD1.n8 585
R1215 VDD1.n24 VDD1.n23 585
R1216 VDD1.n22 VDD1.n21 585
R1217 VDD1.n13 VDD1.n12 585
R1218 VDD1.n16 VDD1.n15 585
R1219 VDD1.n60 VDD1.n59 585
R1220 VDD1.n57 VDD1.n56 585
R1221 VDD1.n66 VDD1.n65 585
R1222 VDD1.n68 VDD1.n67 585
R1223 VDD1.n53 VDD1.n52 585
R1224 VDD1.n74 VDD1.n73 585
R1225 VDD1.n77 VDD1.n76 585
R1226 VDD1.n75 VDD1.n49 585
R1227 VDD1.n82 VDD1.n48 585
R1228 VDD1.n84 VDD1.n83 585
R1229 VDD1.n86 VDD1.n85 585
R1230 VDD1.t0 VDD1.n14 329.039
R1231 VDD1.t1 VDD1.n58 329.038
R1232 VDD1.n40 VDD1.n39 171.744
R1233 VDD1.n39 VDD1.n3 171.744
R1234 VDD1.n7 VDD1.n3 171.744
R1235 VDD1.n31 VDD1.n7 171.744
R1236 VDD1.n31 VDD1.n30 171.744
R1237 VDD1.n30 VDD1.n8 171.744
R1238 VDD1.n23 VDD1.n8 171.744
R1239 VDD1.n23 VDD1.n22 171.744
R1240 VDD1.n22 VDD1.n12 171.744
R1241 VDD1.n15 VDD1.n12 171.744
R1242 VDD1.n59 VDD1.n56 171.744
R1243 VDD1.n66 VDD1.n56 171.744
R1244 VDD1.n67 VDD1.n66 171.744
R1245 VDD1.n67 VDD1.n52 171.744
R1246 VDD1.n74 VDD1.n52 171.744
R1247 VDD1.n76 VDD1.n74 171.744
R1248 VDD1.n76 VDD1.n75 171.744
R1249 VDD1.n75 VDD1.n48 171.744
R1250 VDD1.n84 VDD1.n48 171.744
R1251 VDD1.n85 VDD1.n84 171.744
R1252 VDD1 VDD1.n89 87.6689
R1253 VDD1.n15 VDD1.t0 85.8723
R1254 VDD1.n59 VDD1.t1 85.8723
R1255 VDD1 VDD1.n44 50.9308
R1256 VDD1.n38 VDD1.n37 13.1884
R1257 VDD1.n83 VDD1.n82 13.1884
R1258 VDD1.n41 VDD1.n2 12.8005
R1259 VDD1.n36 VDD1.n4 12.8005
R1260 VDD1.n81 VDD1.n49 12.8005
R1261 VDD1.n86 VDD1.n47 12.8005
R1262 VDD1.n42 VDD1.n0 12.0247
R1263 VDD1.n33 VDD1.n32 12.0247
R1264 VDD1.n78 VDD1.n77 12.0247
R1265 VDD1.n87 VDD1.n45 12.0247
R1266 VDD1.n29 VDD1.n6 11.249
R1267 VDD1.n73 VDD1.n51 11.249
R1268 VDD1.n16 VDD1.n14 10.7239
R1269 VDD1.n60 VDD1.n58 10.7239
R1270 VDD1.n28 VDD1.n9 10.4732
R1271 VDD1.n72 VDD1.n53 10.4732
R1272 VDD1.n25 VDD1.n24 9.69747
R1273 VDD1.n69 VDD1.n68 9.69747
R1274 VDD1.n44 VDD1.n43 9.45567
R1275 VDD1.n89 VDD1.n88 9.45567
R1276 VDD1.n18 VDD1.n17 9.3005
R1277 VDD1.n20 VDD1.n19 9.3005
R1278 VDD1.n11 VDD1.n10 9.3005
R1279 VDD1.n26 VDD1.n25 9.3005
R1280 VDD1.n28 VDD1.n27 9.3005
R1281 VDD1.n6 VDD1.n5 9.3005
R1282 VDD1.n34 VDD1.n33 9.3005
R1283 VDD1.n36 VDD1.n35 9.3005
R1284 VDD1.n43 VDD1.n42 9.3005
R1285 VDD1.n2 VDD1.n1 9.3005
R1286 VDD1.n88 VDD1.n87 9.3005
R1287 VDD1.n47 VDD1.n46 9.3005
R1288 VDD1.n62 VDD1.n61 9.3005
R1289 VDD1.n64 VDD1.n63 9.3005
R1290 VDD1.n55 VDD1.n54 9.3005
R1291 VDD1.n70 VDD1.n69 9.3005
R1292 VDD1.n72 VDD1.n71 9.3005
R1293 VDD1.n51 VDD1.n50 9.3005
R1294 VDD1.n79 VDD1.n78 9.3005
R1295 VDD1.n81 VDD1.n80 9.3005
R1296 VDD1.n21 VDD1.n11 8.92171
R1297 VDD1.n65 VDD1.n55 8.92171
R1298 VDD1.n20 VDD1.n13 8.14595
R1299 VDD1.n64 VDD1.n57 8.14595
R1300 VDD1.n17 VDD1.n16 7.3702
R1301 VDD1.n61 VDD1.n60 7.3702
R1302 VDD1.n17 VDD1.n13 5.81868
R1303 VDD1.n61 VDD1.n57 5.81868
R1304 VDD1.n21 VDD1.n20 5.04292
R1305 VDD1.n65 VDD1.n64 5.04292
R1306 VDD1.n24 VDD1.n11 4.26717
R1307 VDD1.n68 VDD1.n55 4.26717
R1308 VDD1.n25 VDD1.n9 3.49141
R1309 VDD1.n69 VDD1.n53 3.49141
R1310 VDD1.n29 VDD1.n28 2.71565
R1311 VDD1.n73 VDD1.n72 2.71565
R1312 VDD1.n18 VDD1.n14 2.41285
R1313 VDD1.n62 VDD1.n58 2.41285
R1314 VDD1.n44 VDD1.n0 1.93989
R1315 VDD1.n32 VDD1.n6 1.93989
R1316 VDD1.n77 VDD1.n51 1.93989
R1317 VDD1.n89 VDD1.n45 1.93989
R1318 VDD1.n42 VDD1.n41 1.16414
R1319 VDD1.n33 VDD1.n4 1.16414
R1320 VDD1.n78 VDD1.n49 1.16414
R1321 VDD1.n87 VDD1.n86 1.16414
R1322 VDD1.n38 VDD1.n2 0.388379
R1323 VDD1.n37 VDD1.n36 0.388379
R1324 VDD1.n82 VDD1.n81 0.388379
R1325 VDD1.n83 VDD1.n47 0.388379
R1326 VDD1.n43 VDD1.n1 0.155672
R1327 VDD1.n35 VDD1.n1 0.155672
R1328 VDD1.n35 VDD1.n34 0.155672
R1329 VDD1.n34 VDD1.n5 0.155672
R1330 VDD1.n27 VDD1.n5 0.155672
R1331 VDD1.n27 VDD1.n26 0.155672
R1332 VDD1.n26 VDD1.n10 0.155672
R1333 VDD1.n19 VDD1.n10 0.155672
R1334 VDD1.n19 VDD1.n18 0.155672
R1335 VDD1.n63 VDD1.n62 0.155672
R1336 VDD1.n63 VDD1.n54 0.155672
R1337 VDD1.n70 VDD1.n54 0.155672
R1338 VDD1.n71 VDD1.n70 0.155672
R1339 VDD1.n71 VDD1.n50 0.155672
R1340 VDD1.n79 VDD1.n50 0.155672
R1341 VDD1.n80 VDD1.n79 0.155672
R1342 VDD1.n80 VDD1.n46 0.155672
R1343 VDD1.n88 VDD1.n46 0.155672
C0 w_n2178_n2686# VP 3.24321f
C1 VDD2 VN 2.07082f
C2 VTAIL B 2.92464f
C3 VN VDD1 0.148163f
C4 VN VP 4.86979f
C5 VDD2 B 1.4786f
C6 w_n2178_n2686# VN 2.96558f
C7 VDD2 VTAIL 4.23679f
C8 B VDD1 1.44772f
C9 B VP 1.48183f
C10 VTAIL VDD1 4.18471f
C11 VTAIL VP 1.91275f
C12 w_n2178_n2686# B 7.94999f
C13 w_n2178_n2686# VTAIL 2.26932f
C14 VDD2 VDD1 0.685083f
C15 VDD2 VP 0.336579f
C16 VDD2 w_n2178_n2686# 1.58179f
C17 B VN 1.02504f
C18 VDD1 VP 2.25733f
C19 VTAIL VN 1.89852f
C20 w_n2178_n2686# VDD1 1.55479f
C21 VDD2 VSUBS 0.791271f
C22 VDD1 VSUBS 3.382489f
C23 VTAIL VSUBS 0.84308f
C24 VN VSUBS 6.52279f
C25 VP VSUBS 1.584387f
C26 B VSUBS 3.687038f
C27 w_n2178_n2686# VSUBS 72.4751f
C28 VDD1.n0 VSUBS 0.021815f
C29 VDD1.n1 VSUBS 0.020986f
C30 VDD1.n2 VSUBS 0.011277f
C31 VDD1.n3 VSUBS 0.026655f
C32 VDD1.n4 VSUBS 0.01194f
C33 VDD1.n5 VSUBS 0.020986f
C34 VDD1.n6 VSUBS 0.011277f
C35 VDD1.n7 VSUBS 0.026655f
C36 VDD1.n8 VSUBS 0.026655f
C37 VDD1.n9 VSUBS 0.01194f
C38 VDD1.n10 VSUBS 0.020986f
C39 VDD1.n11 VSUBS 0.011277f
C40 VDD1.n12 VSUBS 0.026655f
C41 VDD1.n13 VSUBS 0.01194f
C42 VDD1.n14 VSUBS 0.132963f
C43 VDD1.t0 VSUBS 0.057246f
C44 VDD1.n15 VSUBS 0.019991f
C45 VDD1.n16 VSUBS 0.020051f
C46 VDD1.n17 VSUBS 0.011277f
C47 VDD1.n18 VSUBS 0.717463f
C48 VDD1.n19 VSUBS 0.020986f
C49 VDD1.n20 VSUBS 0.011277f
C50 VDD1.n21 VSUBS 0.01194f
C51 VDD1.n22 VSUBS 0.026655f
C52 VDD1.n23 VSUBS 0.026655f
C53 VDD1.n24 VSUBS 0.01194f
C54 VDD1.n25 VSUBS 0.011277f
C55 VDD1.n26 VSUBS 0.020986f
C56 VDD1.n27 VSUBS 0.020986f
C57 VDD1.n28 VSUBS 0.011277f
C58 VDD1.n29 VSUBS 0.01194f
C59 VDD1.n30 VSUBS 0.026655f
C60 VDD1.n31 VSUBS 0.026655f
C61 VDD1.n32 VSUBS 0.01194f
C62 VDD1.n33 VSUBS 0.011277f
C63 VDD1.n34 VSUBS 0.020986f
C64 VDD1.n35 VSUBS 0.020986f
C65 VDD1.n36 VSUBS 0.011277f
C66 VDD1.n37 VSUBS 0.011609f
C67 VDD1.n38 VSUBS 0.011609f
C68 VDD1.n39 VSUBS 0.026655f
C69 VDD1.n40 VSUBS 0.06029f
C70 VDD1.n41 VSUBS 0.01194f
C71 VDD1.n42 VSUBS 0.011277f
C72 VDD1.n43 VSUBS 0.050515f
C73 VDD1.n44 VSUBS 0.045913f
C74 VDD1.n45 VSUBS 0.021815f
C75 VDD1.n46 VSUBS 0.020986f
C76 VDD1.n47 VSUBS 0.011277f
C77 VDD1.n48 VSUBS 0.026655f
C78 VDD1.n49 VSUBS 0.01194f
C79 VDD1.n50 VSUBS 0.020986f
C80 VDD1.n51 VSUBS 0.011277f
C81 VDD1.n52 VSUBS 0.026655f
C82 VDD1.n53 VSUBS 0.01194f
C83 VDD1.n54 VSUBS 0.020986f
C84 VDD1.n55 VSUBS 0.011277f
C85 VDD1.n56 VSUBS 0.026655f
C86 VDD1.n57 VSUBS 0.01194f
C87 VDD1.n58 VSUBS 0.132963f
C88 VDD1.t1 VSUBS 0.057246f
C89 VDD1.n59 VSUBS 0.019991f
C90 VDD1.n60 VSUBS 0.020051f
C91 VDD1.n61 VSUBS 0.011277f
C92 VDD1.n62 VSUBS 0.717462f
C93 VDD1.n63 VSUBS 0.020986f
C94 VDD1.n64 VSUBS 0.011277f
C95 VDD1.n65 VSUBS 0.01194f
C96 VDD1.n66 VSUBS 0.026655f
C97 VDD1.n67 VSUBS 0.026655f
C98 VDD1.n68 VSUBS 0.01194f
C99 VDD1.n69 VSUBS 0.011277f
C100 VDD1.n70 VSUBS 0.020986f
C101 VDD1.n71 VSUBS 0.020986f
C102 VDD1.n72 VSUBS 0.011277f
C103 VDD1.n73 VSUBS 0.01194f
C104 VDD1.n74 VSUBS 0.026655f
C105 VDD1.n75 VSUBS 0.026655f
C106 VDD1.n76 VSUBS 0.026655f
C107 VDD1.n77 VSUBS 0.01194f
C108 VDD1.n78 VSUBS 0.011277f
C109 VDD1.n79 VSUBS 0.020986f
C110 VDD1.n80 VSUBS 0.020986f
C111 VDD1.n81 VSUBS 0.011277f
C112 VDD1.n82 VSUBS 0.011609f
C113 VDD1.n83 VSUBS 0.011609f
C114 VDD1.n84 VSUBS 0.026655f
C115 VDD1.n85 VSUBS 0.06029f
C116 VDD1.n86 VSUBS 0.01194f
C117 VDD1.n87 VSUBS 0.011277f
C118 VDD1.n88 VSUBS 0.050515f
C119 VDD1.n89 VSUBS 0.553221f
C120 VP.t0 VSUBS 2.71186f
C121 VP.t1 VSUBS 3.36416f
C122 VP.n0 VSUBS 4.22465f
C123 B.n0 VSUBS 0.00428f
C124 B.n1 VSUBS 0.00428f
C125 B.n2 VSUBS 0.006769f
C126 B.n3 VSUBS 0.006769f
C127 B.n4 VSUBS 0.006769f
C128 B.n5 VSUBS 0.006769f
C129 B.n6 VSUBS 0.006769f
C130 B.n7 VSUBS 0.006769f
C131 B.n8 VSUBS 0.006769f
C132 B.n9 VSUBS 0.006769f
C133 B.n10 VSUBS 0.006769f
C134 B.n11 VSUBS 0.006769f
C135 B.n12 VSUBS 0.006769f
C136 B.n13 VSUBS 0.006769f
C137 B.n14 VSUBS 0.006769f
C138 B.n15 VSUBS 0.015347f
C139 B.n16 VSUBS 0.006769f
C140 B.n17 VSUBS 0.006769f
C141 B.n18 VSUBS 0.006769f
C142 B.n19 VSUBS 0.006769f
C143 B.n20 VSUBS 0.006769f
C144 B.n21 VSUBS 0.006769f
C145 B.n22 VSUBS 0.006769f
C146 B.n23 VSUBS 0.006769f
C147 B.n24 VSUBS 0.006769f
C148 B.n25 VSUBS 0.006769f
C149 B.n26 VSUBS 0.006769f
C150 B.n27 VSUBS 0.006769f
C151 B.n28 VSUBS 0.006769f
C152 B.n29 VSUBS 0.006769f
C153 B.n30 VSUBS 0.006769f
C154 B.n31 VSUBS 0.006769f
C155 B.t11 VSUBS 0.133667f
C156 B.t10 VSUBS 0.162798f
C157 B.t9 VSUBS 1.03981f
C158 B.n32 VSUBS 0.267876f
C159 B.n33 VSUBS 0.195035f
C160 B.n34 VSUBS 0.006769f
C161 B.n35 VSUBS 0.006769f
C162 B.n36 VSUBS 0.006769f
C163 B.n37 VSUBS 0.006769f
C164 B.t8 VSUBS 0.133669f
C165 B.t7 VSUBS 0.1628f
C166 B.t6 VSUBS 1.03981f
C167 B.n38 VSUBS 0.267874f
C168 B.n39 VSUBS 0.195032f
C169 B.n40 VSUBS 0.006769f
C170 B.n41 VSUBS 0.006769f
C171 B.n42 VSUBS 0.006769f
C172 B.n43 VSUBS 0.006769f
C173 B.n44 VSUBS 0.006769f
C174 B.n45 VSUBS 0.006769f
C175 B.n46 VSUBS 0.006769f
C176 B.n47 VSUBS 0.006769f
C177 B.n48 VSUBS 0.006769f
C178 B.n49 VSUBS 0.006769f
C179 B.n50 VSUBS 0.006769f
C180 B.n51 VSUBS 0.006769f
C181 B.n52 VSUBS 0.006769f
C182 B.n53 VSUBS 0.006769f
C183 B.n54 VSUBS 0.006769f
C184 B.n55 VSUBS 0.015347f
C185 B.n56 VSUBS 0.006769f
C186 B.n57 VSUBS 0.006769f
C187 B.n58 VSUBS 0.006769f
C188 B.n59 VSUBS 0.006769f
C189 B.n60 VSUBS 0.006769f
C190 B.n61 VSUBS 0.006769f
C191 B.n62 VSUBS 0.006769f
C192 B.n63 VSUBS 0.006769f
C193 B.n64 VSUBS 0.006769f
C194 B.n65 VSUBS 0.006769f
C195 B.n66 VSUBS 0.006769f
C196 B.n67 VSUBS 0.006769f
C197 B.n68 VSUBS 0.006769f
C198 B.n69 VSUBS 0.006769f
C199 B.n70 VSUBS 0.006769f
C200 B.n71 VSUBS 0.006769f
C201 B.n72 VSUBS 0.006769f
C202 B.n73 VSUBS 0.006769f
C203 B.n74 VSUBS 0.006769f
C204 B.n75 VSUBS 0.006769f
C205 B.n76 VSUBS 0.006769f
C206 B.n77 VSUBS 0.006769f
C207 B.n78 VSUBS 0.006769f
C208 B.n79 VSUBS 0.006769f
C209 B.n80 VSUBS 0.006769f
C210 B.n81 VSUBS 0.006769f
C211 B.n82 VSUBS 0.015347f
C212 B.n83 VSUBS 0.006769f
C213 B.n84 VSUBS 0.006769f
C214 B.n85 VSUBS 0.006769f
C215 B.n86 VSUBS 0.006769f
C216 B.n87 VSUBS 0.006769f
C217 B.n88 VSUBS 0.006769f
C218 B.n89 VSUBS 0.006769f
C219 B.n90 VSUBS 0.006769f
C220 B.n91 VSUBS 0.006769f
C221 B.n92 VSUBS 0.006769f
C222 B.n93 VSUBS 0.006769f
C223 B.n94 VSUBS 0.006769f
C224 B.n95 VSUBS 0.006769f
C225 B.n96 VSUBS 0.006769f
C226 B.n97 VSUBS 0.006769f
C227 B.t4 VSUBS 0.133669f
C228 B.t5 VSUBS 0.1628f
C229 B.t3 VSUBS 1.03981f
C230 B.n98 VSUBS 0.267874f
C231 B.n99 VSUBS 0.195032f
C232 B.n100 VSUBS 0.015682f
C233 B.n101 VSUBS 0.006769f
C234 B.n102 VSUBS 0.006769f
C235 B.n103 VSUBS 0.006769f
C236 B.n104 VSUBS 0.006769f
C237 B.n105 VSUBS 0.006769f
C238 B.t1 VSUBS 0.133667f
C239 B.t2 VSUBS 0.162798f
C240 B.t0 VSUBS 1.03981f
C241 B.n106 VSUBS 0.267876f
C242 B.n107 VSUBS 0.195035f
C243 B.n108 VSUBS 0.006769f
C244 B.n109 VSUBS 0.006769f
C245 B.n110 VSUBS 0.006769f
C246 B.n111 VSUBS 0.006769f
C247 B.n112 VSUBS 0.006769f
C248 B.n113 VSUBS 0.006769f
C249 B.n114 VSUBS 0.006769f
C250 B.n115 VSUBS 0.006769f
C251 B.n116 VSUBS 0.006769f
C252 B.n117 VSUBS 0.006769f
C253 B.n118 VSUBS 0.006769f
C254 B.n119 VSUBS 0.006769f
C255 B.n120 VSUBS 0.006769f
C256 B.n121 VSUBS 0.006769f
C257 B.n122 VSUBS 0.006769f
C258 B.n123 VSUBS 0.014514f
C259 B.n124 VSUBS 0.006769f
C260 B.n125 VSUBS 0.006769f
C261 B.n126 VSUBS 0.006769f
C262 B.n127 VSUBS 0.006769f
C263 B.n128 VSUBS 0.006769f
C264 B.n129 VSUBS 0.006769f
C265 B.n130 VSUBS 0.006769f
C266 B.n131 VSUBS 0.006769f
C267 B.n132 VSUBS 0.006769f
C268 B.n133 VSUBS 0.006769f
C269 B.n134 VSUBS 0.006769f
C270 B.n135 VSUBS 0.006769f
C271 B.n136 VSUBS 0.006769f
C272 B.n137 VSUBS 0.006769f
C273 B.n138 VSUBS 0.006769f
C274 B.n139 VSUBS 0.006769f
C275 B.n140 VSUBS 0.006769f
C276 B.n141 VSUBS 0.006769f
C277 B.n142 VSUBS 0.006769f
C278 B.n143 VSUBS 0.006769f
C279 B.n144 VSUBS 0.006769f
C280 B.n145 VSUBS 0.006769f
C281 B.n146 VSUBS 0.006769f
C282 B.n147 VSUBS 0.006769f
C283 B.n148 VSUBS 0.006769f
C284 B.n149 VSUBS 0.006769f
C285 B.n150 VSUBS 0.006769f
C286 B.n151 VSUBS 0.006769f
C287 B.n152 VSUBS 0.006769f
C288 B.n153 VSUBS 0.006769f
C289 B.n154 VSUBS 0.006769f
C290 B.n155 VSUBS 0.006769f
C291 B.n156 VSUBS 0.006769f
C292 B.n157 VSUBS 0.006769f
C293 B.n158 VSUBS 0.006769f
C294 B.n159 VSUBS 0.006769f
C295 B.n160 VSUBS 0.006769f
C296 B.n161 VSUBS 0.006769f
C297 B.n162 VSUBS 0.006769f
C298 B.n163 VSUBS 0.006769f
C299 B.n164 VSUBS 0.006769f
C300 B.n165 VSUBS 0.006769f
C301 B.n166 VSUBS 0.006769f
C302 B.n167 VSUBS 0.006769f
C303 B.n168 VSUBS 0.006769f
C304 B.n169 VSUBS 0.006769f
C305 B.n170 VSUBS 0.006769f
C306 B.n171 VSUBS 0.006769f
C307 B.n172 VSUBS 0.014514f
C308 B.n173 VSUBS 0.015347f
C309 B.n174 VSUBS 0.015347f
C310 B.n175 VSUBS 0.006769f
C311 B.n176 VSUBS 0.006769f
C312 B.n177 VSUBS 0.006769f
C313 B.n178 VSUBS 0.006769f
C314 B.n179 VSUBS 0.006769f
C315 B.n180 VSUBS 0.006769f
C316 B.n181 VSUBS 0.006769f
C317 B.n182 VSUBS 0.006769f
C318 B.n183 VSUBS 0.006769f
C319 B.n184 VSUBS 0.006769f
C320 B.n185 VSUBS 0.006769f
C321 B.n186 VSUBS 0.006769f
C322 B.n187 VSUBS 0.006769f
C323 B.n188 VSUBS 0.006769f
C324 B.n189 VSUBS 0.006769f
C325 B.n190 VSUBS 0.006769f
C326 B.n191 VSUBS 0.006769f
C327 B.n192 VSUBS 0.006769f
C328 B.n193 VSUBS 0.006769f
C329 B.n194 VSUBS 0.006769f
C330 B.n195 VSUBS 0.006769f
C331 B.n196 VSUBS 0.006769f
C332 B.n197 VSUBS 0.006769f
C333 B.n198 VSUBS 0.006769f
C334 B.n199 VSUBS 0.006769f
C335 B.n200 VSUBS 0.006769f
C336 B.n201 VSUBS 0.006769f
C337 B.n202 VSUBS 0.006769f
C338 B.n203 VSUBS 0.006769f
C339 B.n204 VSUBS 0.006769f
C340 B.n205 VSUBS 0.006769f
C341 B.n206 VSUBS 0.006769f
C342 B.n207 VSUBS 0.006769f
C343 B.n208 VSUBS 0.006769f
C344 B.n209 VSUBS 0.006769f
C345 B.n210 VSUBS 0.006769f
C346 B.n211 VSUBS 0.006769f
C347 B.n212 VSUBS 0.006769f
C348 B.n213 VSUBS 0.006769f
C349 B.n214 VSUBS 0.006769f
C350 B.n215 VSUBS 0.006769f
C351 B.n216 VSUBS 0.006769f
C352 B.n217 VSUBS 0.006769f
C353 B.n218 VSUBS 0.006769f
C354 B.n219 VSUBS 0.006769f
C355 B.n220 VSUBS 0.004678f
C356 B.n221 VSUBS 0.015682f
C357 B.n222 VSUBS 0.005475f
C358 B.n223 VSUBS 0.006769f
C359 B.n224 VSUBS 0.006769f
C360 B.n225 VSUBS 0.006769f
C361 B.n226 VSUBS 0.006769f
C362 B.n227 VSUBS 0.006769f
C363 B.n228 VSUBS 0.006769f
C364 B.n229 VSUBS 0.006769f
C365 B.n230 VSUBS 0.006769f
C366 B.n231 VSUBS 0.006769f
C367 B.n232 VSUBS 0.006769f
C368 B.n233 VSUBS 0.006769f
C369 B.n234 VSUBS 0.005475f
C370 B.n235 VSUBS 0.006769f
C371 B.n236 VSUBS 0.006769f
C372 B.n237 VSUBS 0.004678f
C373 B.n238 VSUBS 0.006769f
C374 B.n239 VSUBS 0.006769f
C375 B.n240 VSUBS 0.006769f
C376 B.n241 VSUBS 0.006769f
C377 B.n242 VSUBS 0.006769f
C378 B.n243 VSUBS 0.006769f
C379 B.n244 VSUBS 0.006769f
C380 B.n245 VSUBS 0.006769f
C381 B.n246 VSUBS 0.006769f
C382 B.n247 VSUBS 0.006769f
C383 B.n248 VSUBS 0.006769f
C384 B.n249 VSUBS 0.006769f
C385 B.n250 VSUBS 0.006769f
C386 B.n251 VSUBS 0.006769f
C387 B.n252 VSUBS 0.006769f
C388 B.n253 VSUBS 0.006769f
C389 B.n254 VSUBS 0.006769f
C390 B.n255 VSUBS 0.006769f
C391 B.n256 VSUBS 0.006769f
C392 B.n257 VSUBS 0.006769f
C393 B.n258 VSUBS 0.006769f
C394 B.n259 VSUBS 0.006769f
C395 B.n260 VSUBS 0.006769f
C396 B.n261 VSUBS 0.006769f
C397 B.n262 VSUBS 0.006769f
C398 B.n263 VSUBS 0.006769f
C399 B.n264 VSUBS 0.006769f
C400 B.n265 VSUBS 0.006769f
C401 B.n266 VSUBS 0.006769f
C402 B.n267 VSUBS 0.006769f
C403 B.n268 VSUBS 0.006769f
C404 B.n269 VSUBS 0.006769f
C405 B.n270 VSUBS 0.006769f
C406 B.n271 VSUBS 0.006769f
C407 B.n272 VSUBS 0.006769f
C408 B.n273 VSUBS 0.006769f
C409 B.n274 VSUBS 0.006769f
C410 B.n275 VSUBS 0.006769f
C411 B.n276 VSUBS 0.006769f
C412 B.n277 VSUBS 0.006769f
C413 B.n278 VSUBS 0.006769f
C414 B.n279 VSUBS 0.006769f
C415 B.n280 VSUBS 0.006769f
C416 B.n281 VSUBS 0.006769f
C417 B.n282 VSUBS 0.006769f
C418 B.n283 VSUBS 0.015347f
C419 B.n284 VSUBS 0.014514f
C420 B.n285 VSUBS 0.014514f
C421 B.n286 VSUBS 0.006769f
C422 B.n287 VSUBS 0.006769f
C423 B.n288 VSUBS 0.006769f
C424 B.n289 VSUBS 0.006769f
C425 B.n290 VSUBS 0.006769f
C426 B.n291 VSUBS 0.006769f
C427 B.n292 VSUBS 0.006769f
C428 B.n293 VSUBS 0.006769f
C429 B.n294 VSUBS 0.006769f
C430 B.n295 VSUBS 0.006769f
C431 B.n296 VSUBS 0.006769f
C432 B.n297 VSUBS 0.006769f
C433 B.n298 VSUBS 0.006769f
C434 B.n299 VSUBS 0.006769f
C435 B.n300 VSUBS 0.006769f
C436 B.n301 VSUBS 0.006769f
C437 B.n302 VSUBS 0.006769f
C438 B.n303 VSUBS 0.006769f
C439 B.n304 VSUBS 0.006769f
C440 B.n305 VSUBS 0.006769f
C441 B.n306 VSUBS 0.006769f
C442 B.n307 VSUBS 0.006769f
C443 B.n308 VSUBS 0.006769f
C444 B.n309 VSUBS 0.006769f
C445 B.n310 VSUBS 0.006769f
C446 B.n311 VSUBS 0.006769f
C447 B.n312 VSUBS 0.006769f
C448 B.n313 VSUBS 0.006769f
C449 B.n314 VSUBS 0.006769f
C450 B.n315 VSUBS 0.006769f
C451 B.n316 VSUBS 0.006769f
C452 B.n317 VSUBS 0.006769f
C453 B.n318 VSUBS 0.006769f
C454 B.n319 VSUBS 0.006769f
C455 B.n320 VSUBS 0.006769f
C456 B.n321 VSUBS 0.006769f
C457 B.n322 VSUBS 0.006769f
C458 B.n323 VSUBS 0.006769f
C459 B.n324 VSUBS 0.006769f
C460 B.n325 VSUBS 0.006769f
C461 B.n326 VSUBS 0.006769f
C462 B.n327 VSUBS 0.006769f
C463 B.n328 VSUBS 0.006769f
C464 B.n329 VSUBS 0.006769f
C465 B.n330 VSUBS 0.006769f
C466 B.n331 VSUBS 0.006769f
C467 B.n332 VSUBS 0.006769f
C468 B.n333 VSUBS 0.006769f
C469 B.n334 VSUBS 0.006769f
C470 B.n335 VSUBS 0.006769f
C471 B.n336 VSUBS 0.006769f
C472 B.n337 VSUBS 0.006769f
C473 B.n338 VSUBS 0.006769f
C474 B.n339 VSUBS 0.006769f
C475 B.n340 VSUBS 0.006769f
C476 B.n341 VSUBS 0.006769f
C477 B.n342 VSUBS 0.006769f
C478 B.n343 VSUBS 0.006769f
C479 B.n344 VSUBS 0.006769f
C480 B.n345 VSUBS 0.006769f
C481 B.n346 VSUBS 0.006769f
C482 B.n347 VSUBS 0.006769f
C483 B.n348 VSUBS 0.006769f
C484 B.n349 VSUBS 0.006769f
C485 B.n350 VSUBS 0.006769f
C486 B.n351 VSUBS 0.006769f
C487 B.n352 VSUBS 0.006769f
C488 B.n353 VSUBS 0.006769f
C489 B.n354 VSUBS 0.006769f
C490 B.n355 VSUBS 0.006769f
C491 B.n356 VSUBS 0.006769f
C492 B.n357 VSUBS 0.006769f
C493 B.n358 VSUBS 0.006769f
C494 B.n359 VSUBS 0.006769f
C495 B.n360 VSUBS 0.006769f
C496 B.n361 VSUBS 0.006769f
C497 B.n362 VSUBS 0.014514f
C498 B.n363 VSUBS 0.01539f
C499 B.n364 VSUBS 0.014471f
C500 B.n365 VSUBS 0.006769f
C501 B.n366 VSUBS 0.006769f
C502 B.n367 VSUBS 0.006769f
C503 B.n368 VSUBS 0.006769f
C504 B.n369 VSUBS 0.006769f
C505 B.n370 VSUBS 0.006769f
C506 B.n371 VSUBS 0.006769f
C507 B.n372 VSUBS 0.006769f
C508 B.n373 VSUBS 0.006769f
C509 B.n374 VSUBS 0.006769f
C510 B.n375 VSUBS 0.006769f
C511 B.n376 VSUBS 0.006769f
C512 B.n377 VSUBS 0.006769f
C513 B.n378 VSUBS 0.006769f
C514 B.n379 VSUBS 0.006769f
C515 B.n380 VSUBS 0.006769f
C516 B.n381 VSUBS 0.006769f
C517 B.n382 VSUBS 0.006769f
C518 B.n383 VSUBS 0.006769f
C519 B.n384 VSUBS 0.006769f
C520 B.n385 VSUBS 0.006769f
C521 B.n386 VSUBS 0.006769f
C522 B.n387 VSUBS 0.006769f
C523 B.n388 VSUBS 0.006769f
C524 B.n389 VSUBS 0.006769f
C525 B.n390 VSUBS 0.006769f
C526 B.n391 VSUBS 0.006769f
C527 B.n392 VSUBS 0.006769f
C528 B.n393 VSUBS 0.006769f
C529 B.n394 VSUBS 0.006769f
C530 B.n395 VSUBS 0.006769f
C531 B.n396 VSUBS 0.006769f
C532 B.n397 VSUBS 0.006769f
C533 B.n398 VSUBS 0.006769f
C534 B.n399 VSUBS 0.006769f
C535 B.n400 VSUBS 0.006769f
C536 B.n401 VSUBS 0.006769f
C537 B.n402 VSUBS 0.006769f
C538 B.n403 VSUBS 0.006769f
C539 B.n404 VSUBS 0.006769f
C540 B.n405 VSUBS 0.006769f
C541 B.n406 VSUBS 0.006769f
C542 B.n407 VSUBS 0.006769f
C543 B.n408 VSUBS 0.006769f
C544 B.n409 VSUBS 0.006769f
C545 B.n410 VSUBS 0.006769f
C546 B.n411 VSUBS 0.004678f
C547 B.n412 VSUBS 0.015682f
C548 B.n413 VSUBS 0.005475f
C549 B.n414 VSUBS 0.006769f
C550 B.n415 VSUBS 0.006769f
C551 B.n416 VSUBS 0.006769f
C552 B.n417 VSUBS 0.006769f
C553 B.n418 VSUBS 0.006769f
C554 B.n419 VSUBS 0.006769f
C555 B.n420 VSUBS 0.006769f
C556 B.n421 VSUBS 0.006769f
C557 B.n422 VSUBS 0.006769f
C558 B.n423 VSUBS 0.006769f
C559 B.n424 VSUBS 0.006769f
C560 B.n425 VSUBS 0.005475f
C561 B.n426 VSUBS 0.015682f
C562 B.n427 VSUBS 0.004678f
C563 B.n428 VSUBS 0.006769f
C564 B.n429 VSUBS 0.006769f
C565 B.n430 VSUBS 0.006769f
C566 B.n431 VSUBS 0.006769f
C567 B.n432 VSUBS 0.006769f
C568 B.n433 VSUBS 0.006769f
C569 B.n434 VSUBS 0.006769f
C570 B.n435 VSUBS 0.006769f
C571 B.n436 VSUBS 0.006769f
C572 B.n437 VSUBS 0.006769f
C573 B.n438 VSUBS 0.006769f
C574 B.n439 VSUBS 0.006769f
C575 B.n440 VSUBS 0.006769f
C576 B.n441 VSUBS 0.006769f
C577 B.n442 VSUBS 0.006769f
C578 B.n443 VSUBS 0.006769f
C579 B.n444 VSUBS 0.006769f
C580 B.n445 VSUBS 0.006769f
C581 B.n446 VSUBS 0.006769f
C582 B.n447 VSUBS 0.006769f
C583 B.n448 VSUBS 0.006769f
C584 B.n449 VSUBS 0.006769f
C585 B.n450 VSUBS 0.006769f
C586 B.n451 VSUBS 0.006769f
C587 B.n452 VSUBS 0.006769f
C588 B.n453 VSUBS 0.006769f
C589 B.n454 VSUBS 0.006769f
C590 B.n455 VSUBS 0.006769f
C591 B.n456 VSUBS 0.006769f
C592 B.n457 VSUBS 0.006769f
C593 B.n458 VSUBS 0.006769f
C594 B.n459 VSUBS 0.006769f
C595 B.n460 VSUBS 0.006769f
C596 B.n461 VSUBS 0.006769f
C597 B.n462 VSUBS 0.006769f
C598 B.n463 VSUBS 0.006769f
C599 B.n464 VSUBS 0.006769f
C600 B.n465 VSUBS 0.006769f
C601 B.n466 VSUBS 0.006769f
C602 B.n467 VSUBS 0.006769f
C603 B.n468 VSUBS 0.006769f
C604 B.n469 VSUBS 0.006769f
C605 B.n470 VSUBS 0.006769f
C606 B.n471 VSUBS 0.006769f
C607 B.n472 VSUBS 0.006769f
C608 B.n473 VSUBS 0.006769f
C609 B.n474 VSUBS 0.015347f
C610 B.n475 VSUBS 0.014514f
C611 B.n476 VSUBS 0.014514f
C612 B.n477 VSUBS 0.006769f
C613 B.n478 VSUBS 0.006769f
C614 B.n479 VSUBS 0.006769f
C615 B.n480 VSUBS 0.006769f
C616 B.n481 VSUBS 0.006769f
C617 B.n482 VSUBS 0.006769f
C618 B.n483 VSUBS 0.006769f
C619 B.n484 VSUBS 0.006769f
C620 B.n485 VSUBS 0.006769f
C621 B.n486 VSUBS 0.006769f
C622 B.n487 VSUBS 0.006769f
C623 B.n488 VSUBS 0.006769f
C624 B.n489 VSUBS 0.006769f
C625 B.n490 VSUBS 0.006769f
C626 B.n491 VSUBS 0.006769f
C627 B.n492 VSUBS 0.006769f
C628 B.n493 VSUBS 0.006769f
C629 B.n494 VSUBS 0.006769f
C630 B.n495 VSUBS 0.006769f
C631 B.n496 VSUBS 0.006769f
C632 B.n497 VSUBS 0.006769f
C633 B.n498 VSUBS 0.006769f
C634 B.n499 VSUBS 0.006769f
C635 B.n500 VSUBS 0.006769f
C636 B.n501 VSUBS 0.006769f
C637 B.n502 VSUBS 0.006769f
C638 B.n503 VSUBS 0.006769f
C639 B.n504 VSUBS 0.006769f
C640 B.n505 VSUBS 0.006769f
C641 B.n506 VSUBS 0.006769f
C642 B.n507 VSUBS 0.006769f
C643 B.n508 VSUBS 0.006769f
C644 B.n509 VSUBS 0.006769f
C645 B.n510 VSUBS 0.006769f
C646 B.n511 VSUBS 0.006769f
C647 B.n512 VSUBS 0.006769f
C648 B.n513 VSUBS 0.006769f
C649 B.n514 VSUBS 0.006769f
C650 B.n515 VSUBS 0.015326f
C651 VDD2.n0 VSUBS 0.021399f
C652 VDD2.n1 VSUBS 0.020586f
C653 VDD2.n2 VSUBS 0.011062f
C654 VDD2.n3 VSUBS 0.026146f
C655 VDD2.n4 VSUBS 0.011713f
C656 VDD2.n5 VSUBS 0.020586f
C657 VDD2.n6 VSUBS 0.011062f
C658 VDD2.n7 VSUBS 0.026146f
C659 VDD2.n8 VSUBS 0.011713f
C660 VDD2.n9 VSUBS 0.020586f
C661 VDD2.n10 VSUBS 0.011062f
C662 VDD2.n11 VSUBS 0.026146f
C663 VDD2.n12 VSUBS 0.011713f
C664 VDD2.n13 VSUBS 0.130427f
C665 VDD2.t1 VSUBS 0.056155f
C666 VDD2.n14 VSUBS 0.01961f
C667 VDD2.n15 VSUBS 0.019669f
C668 VDD2.n16 VSUBS 0.011062f
C669 VDD2.n17 VSUBS 0.703779f
C670 VDD2.n18 VSUBS 0.020586f
C671 VDD2.n19 VSUBS 0.011062f
C672 VDD2.n20 VSUBS 0.011713f
C673 VDD2.n21 VSUBS 0.026146f
C674 VDD2.n22 VSUBS 0.026146f
C675 VDD2.n23 VSUBS 0.011713f
C676 VDD2.n24 VSUBS 0.011062f
C677 VDD2.n25 VSUBS 0.020586f
C678 VDD2.n26 VSUBS 0.020586f
C679 VDD2.n27 VSUBS 0.011062f
C680 VDD2.n28 VSUBS 0.011713f
C681 VDD2.n29 VSUBS 0.026146f
C682 VDD2.n30 VSUBS 0.026146f
C683 VDD2.n31 VSUBS 0.026146f
C684 VDD2.n32 VSUBS 0.011713f
C685 VDD2.n33 VSUBS 0.011062f
C686 VDD2.n34 VSUBS 0.020586f
C687 VDD2.n35 VSUBS 0.020586f
C688 VDD2.n36 VSUBS 0.011062f
C689 VDD2.n37 VSUBS 0.011387f
C690 VDD2.n38 VSUBS 0.011387f
C691 VDD2.n39 VSUBS 0.026146f
C692 VDD2.n40 VSUBS 0.05914f
C693 VDD2.n41 VSUBS 0.011713f
C694 VDD2.n42 VSUBS 0.011062f
C695 VDD2.n43 VSUBS 0.049552f
C696 VDD2.n44 VSUBS 0.504661f
C697 VDD2.n45 VSUBS 0.021399f
C698 VDD2.n46 VSUBS 0.020586f
C699 VDD2.n47 VSUBS 0.011062f
C700 VDD2.n48 VSUBS 0.026146f
C701 VDD2.n49 VSUBS 0.011713f
C702 VDD2.n50 VSUBS 0.020586f
C703 VDD2.n51 VSUBS 0.011062f
C704 VDD2.n52 VSUBS 0.026146f
C705 VDD2.n53 VSUBS 0.026146f
C706 VDD2.n54 VSUBS 0.011713f
C707 VDD2.n55 VSUBS 0.020586f
C708 VDD2.n56 VSUBS 0.011062f
C709 VDD2.n57 VSUBS 0.026146f
C710 VDD2.n58 VSUBS 0.011713f
C711 VDD2.n59 VSUBS 0.130427f
C712 VDD2.t0 VSUBS 0.056155f
C713 VDD2.n60 VSUBS 0.01961f
C714 VDD2.n61 VSUBS 0.019669f
C715 VDD2.n62 VSUBS 0.011062f
C716 VDD2.n63 VSUBS 0.703779f
C717 VDD2.n64 VSUBS 0.020586f
C718 VDD2.n65 VSUBS 0.011062f
C719 VDD2.n66 VSUBS 0.011713f
C720 VDD2.n67 VSUBS 0.026146f
C721 VDD2.n68 VSUBS 0.026146f
C722 VDD2.n69 VSUBS 0.011713f
C723 VDD2.n70 VSUBS 0.011062f
C724 VDD2.n71 VSUBS 0.020586f
C725 VDD2.n72 VSUBS 0.020586f
C726 VDD2.n73 VSUBS 0.011062f
C727 VDD2.n74 VSUBS 0.011713f
C728 VDD2.n75 VSUBS 0.026146f
C729 VDD2.n76 VSUBS 0.026146f
C730 VDD2.n77 VSUBS 0.011713f
C731 VDD2.n78 VSUBS 0.011062f
C732 VDD2.n79 VSUBS 0.020586f
C733 VDD2.n80 VSUBS 0.020586f
C734 VDD2.n81 VSUBS 0.011062f
C735 VDD2.n82 VSUBS 0.011387f
C736 VDD2.n83 VSUBS 0.011387f
C737 VDD2.n84 VSUBS 0.026146f
C738 VDD2.n85 VSUBS 0.05914f
C739 VDD2.n86 VSUBS 0.011713f
C740 VDD2.n87 VSUBS 0.011062f
C741 VDD2.n88 VSUBS 0.049552f
C742 VDD2.n89 VSUBS 0.043815f
C743 VDD2.n90 VSUBS 2.24391f
C744 VTAIL.n0 VSUBS 0.02524f
C745 VTAIL.n1 VSUBS 0.024281f
C746 VTAIL.n2 VSUBS 0.013048f
C747 VTAIL.n3 VSUBS 0.03084f
C748 VTAIL.n4 VSUBS 0.013815f
C749 VTAIL.n5 VSUBS 0.024281f
C750 VTAIL.n6 VSUBS 0.013048f
C751 VTAIL.n7 VSUBS 0.03084f
C752 VTAIL.n8 VSUBS 0.013815f
C753 VTAIL.n9 VSUBS 0.024281f
C754 VTAIL.n10 VSUBS 0.013048f
C755 VTAIL.n11 VSUBS 0.03084f
C756 VTAIL.n12 VSUBS 0.013815f
C757 VTAIL.n13 VSUBS 0.153841f
C758 VTAIL.t1 VSUBS 0.066235f
C759 VTAIL.n14 VSUBS 0.02313f
C760 VTAIL.n15 VSUBS 0.0232f
C761 VTAIL.n16 VSUBS 0.013048f
C762 VTAIL.n17 VSUBS 0.830121f
C763 VTAIL.n18 VSUBS 0.024281f
C764 VTAIL.n19 VSUBS 0.013048f
C765 VTAIL.n20 VSUBS 0.013815f
C766 VTAIL.n21 VSUBS 0.03084f
C767 VTAIL.n22 VSUBS 0.03084f
C768 VTAIL.n23 VSUBS 0.013815f
C769 VTAIL.n24 VSUBS 0.013048f
C770 VTAIL.n25 VSUBS 0.024281f
C771 VTAIL.n26 VSUBS 0.024281f
C772 VTAIL.n27 VSUBS 0.013048f
C773 VTAIL.n28 VSUBS 0.013815f
C774 VTAIL.n29 VSUBS 0.03084f
C775 VTAIL.n30 VSUBS 0.03084f
C776 VTAIL.n31 VSUBS 0.03084f
C777 VTAIL.n32 VSUBS 0.013815f
C778 VTAIL.n33 VSUBS 0.013048f
C779 VTAIL.n34 VSUBS 0.024281f
C780 VTAIL.n35 VSUBS 0.024281f
C781 VTAIL.n36 VSUBS 0.013048f
C782 VTAIL.n37 VSUBS 0.013432f
C783 VTAIL.n38 VSUBS 0.013432f
C784 VTAIL.n39 VSUBS 0.03084f
C785 VTAIL.n40 VSUBS 0.069757f
C786 VTAIL.n41 VSUBS 0.013815f
C787 VTAIL.n42 VSUBS 0.013048f
C788 VTAIL.n43 VSUBS 0.058447f
C789 VTAIL.n44 VSUBS 0.034933f
C790 VTAIL.n45 VSUBS 1.43089f
C791 VTAIL.n46 VSUBS 0.02524f
C792 VTAIL.n47 VSUBS 0.024281f
C793 VTAIL.n48 VSUBS 0.013048f
C794 VTAIL.n49 VSUBS 0.03084f
C795 VTAIL.n50 VSUBS 0.013815f
C796 VTAIL.n51 VSUBS 0.024281f
C797 VTAIL.n52 VSUBS 0.013048f
C798 VTAIL.n53 VSUBS 0.03084f
C799 VTAIL.n54 VSUBS 0.03084f
C800 VTAIL.n55 VSUBS 0.013815f
C801 VTAIL.n56 VSUBS 0.024281f
C802 VTAIL.n57 VSUBS 0.013048f
C803 VTAIL.n58 VSUBS 0.03084f
C804 VTAIL.n59 VSUBS 0.013815f
C805 VTAIL.n60 VSUBS 0.153841f
C806 VTAIL.t3 VSUBS 0.066235f
C807 VTAIL.n61 VSUBS 0.02313f
C808 VTAIL.n62 VSUBS 0.0232f
C809 VTAIL.n63 VSUBS 0.013048f
C810 VTAIL.n64 VSUBS 0.830121f
C811 VTAIL.n65 VSUBS 0.024281f
C812 VTAIL.n66 VSUBS 0.013048f
C813 VTAIL.n67 VSUBS 0.013815f
C814 VTAIL.n68 VSUBS 0.03084f
C815 VTAIL.n69 VSUBS 0.03084f
C816 VTAIL.n70 VSUBS 0.013815f
C817 VTAIL.n71 VSUBS 0.013048f
C818 VTAIL.n72 VSUBS 0.024281f
C819 VTAIL.n73 VSUBS 0.024281f
C820 VTAIL.n74 VSUBS 0.013048f
C821 VTAIL.n75 VSUBS 0.013815f
C822 VTAIL.n76 VSUBS 0.03084f
C823 VTAIL.n77 VSUBS 0.03084f
C824 VTAIL.n78 VSUBS 0.013815f
C825 VTAIL.n79 VSUBS 0.013048f
C826 VTAIL.n80 VSUBS 0.024281f
C827 VTAIL.n81 VSUBS 0.024281f
C828 VTAIL.n82 VSUBS 0.013048f
C829 VTAIL.n83 VSUBS 0.013432f
C830 VTAIL.n84 VSUBS 0.013432f
C831 VTAIL.n85 VSUBS 0.03084f
C832 VTAIL.n86 VSUBS 0.069757f
C833 VTAIL.n87 VSUBS 0.013815f
C834 VTAIL.n88 VSUBS 0.013048f
C835 VTAIL.n89 VSUBS 0.058447f
C836 VTAIL.n90 VSUBS 0.034933f
C837 VTAIL.n91 VSUBS 1.47726f
C838 VTAIL.n92 VSUBS 0.02524f
C839 VTAIL.n93 VSUBS 0.024281f
C840 VTAIL.n94 VSUBS 0.013048f
C841 VTAIL.n95 VSUBS 0.03084f
C842 VTAIL.n96 VSUBS 0.013815f
C843 VTAIL.n97 VSUBS 0.024281f
C844 VTAIL.n98 VSUBS 0.013048f
C845 VTAIL.n99 VSUBS 0.03084f
C846 VTAIL.n100 VSUBS 0.03084f
C847 VTAIL.n101 VSUBS 0.013815f
C848 VTAIL.n102 VSUBS 0.024281f
C849 VTAIL.n103 VSUBS 0.013048f
C850 VTAIL.n104 VSUBS 0.03084f
C851 VTAIL.n105 VSUBS 0.013815f
C852 VTAIL.n106 VSUBS 0.153841f
C853 VTAIL.t0 VSUBS 0.066235f
C854 VTAIL.n107 VSUBS 0.02313f
C855 VTAIL.n108 VSUBS 0.0232f
C856 VTAIL.n109 VSUBS 0.013048f
C857 VTAIL.n110 VSUBS 0.830121f
C858 VTAIL.n111 VSUBS 0.024281f
C859 VTAIL.n112 VSUBS 0.013048f
C860 VTAIL.n113 VSUBS 0.013815f
C861 VTAIL.n114 VSUBS 0.03084f
C862 VTAIL.n115 VSUBS 0.03084f
C863 VTAIL.n116 VSUBS 0.013815f
C864 VTAIL.n117 VSUBS 0.013048f
C865 VTAIL.n118 VSUBS 0.024281f
C866 VTAIL.n119 VSUBS 0.024281f
C867 VTAIL.n120 VSUBS 0.013048f
C868 VTAIL.n121 VSUBS 0.013815f
C869 VTAIL.n122 VSUBS 0.03084f
C870 VTAIL.n123 VSUBS 0.03084f
C871 VTAIL.n124 VSUBS 0.013815f
C872 VTAIL.n125 VSUBS 0.013048f
C873 VTAIL.n126 VSUBS 0.024281f
C874 VTAIL.n127 VSUBS 0.024281f
C875 VTAIL.n128 VSUBS 0.013048f
C876 VTAIL.n129 VSUBS 0.013432f
C877 VTAIL.n130 VSUBS 0.013432f
C878 VTAIL.n131 VSUBS 0.03084f
C879 VTAIL.n132 VSUBS 0.069757f
C880 VTAIL.n133 VSUBS 0.013815f
C881 VTAIL.n134 VSUBS 0.013048f
C882 VTAIL.n135 VSUBS 0.058447f
C883 VTAIL.n136 VSUBS 0.034933f
C884 VTAIL.n137 VSUBS 1.27357f
C885 VTAIL.n138 VSUBS 0.02524f
C886 VTAIL.n139 VSUBS 0.024281f
C887 VTAIL.n140 VSUBS 0.013048f
C888 VTAIL.n141 VSUBS 0.03084f
C889 VTAIL.n142 VSUBS 0.013815f
C890 VTAIL.n143 VSUBS 0.024281f
C891 VTAIL.n144 VSUBS 0.013048f
C892 VTAIL.n145 VSUBS 0.03084f
C893 VTAIL.n146 VSUBS 0.013815f
C894 VTAIL.n147 VSUBS 0.024281f
C895 VTAIL.n148 VSUBS 0.013048f
C896 VTAIL.n149 VSUBS 0.03084f
C897 VTAIL.n150 VSUBS 0.013815f
C898 VTAIL.n151 VSUBS 0.153841f
C899 VTAIL.t2 VSUBS 0.066235f
C900 VTAIL.n152 VSUBS 0.02313f
C901 VTAIL.n153 VSUBS 0.0232f
C902 VTAIL.n154 VSUBS 0.013048f
C903 VTAIL.n155 VSUBS 0.830121f
C904 VTAIL.n156 VSUBS 0.024281f
C905 VTAIL.n157 VSUBS 0.013048f
C906 VTAIL.n158 VSUBS 0.013815f
C907 VTAIL.n159 VSUBS 0.03084f
C908 VTAIL.n160 VSUBS 0.03084f
C909 VTAIL.n161 VSUBS 0.013815f
C910 VTAIL.n162 VSUBS 0.013048f
C911 VTAIL.n163 VSUBS 0.024281f
C912 VTAIL.n164 VSUBS 0.024281f
C913 VTAIL.n165 VSUBS 0.013048f
C914 VTAIL.n166 VSUBS 0.013815f
C915 VTAIL.n167 VSUBS 0.03084f
C916 VTAIL.n168 VSUBS 0.03084f
C917 VTAIL.n169 VSUBS 0.03084f
C918 VTAIL.n170 VSUBS 0.013815f
C919 VTAIL.n171 VSUBS 0.013048f
C920 VTAIL.n172 VSUBS 0.024281f
C921 VTAIL.n173 VSUBS 0.024281f
C922 VTAIL.n174 VSUBS 0.013048f
C923 VTAIL.n175 VSUBS 0.013432f
C924 VTAIL.n176 VSUBS 0.013432f
C925 VTAIL.n177 VSUBS 0.03084f
C926 VTAIL.n178 VSUBS 0.069757f
C927 VTAIL.n179 VSUBS 0.013815f
C928 VTAIL.n180 VSUBS 0.013048f
C929 VTAIL.n181 VSUBS 0.058447f
C930 VTAIL.n182 VSUBS 0.034933f
C931 VTAIL.n183 VSUBS 1.18133f
C932 VN.t0 VSUBS 2.59756f
C933 VN.t1 VSUBS 3.22098f
.ends

