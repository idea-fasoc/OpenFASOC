* NGSPICE file created from diff_pair_sample_0046.ext - technology: sky130A

.subckt diff_pair_sample_0046 VTAIL VN VP B VDD2 VDD1
X0 B.t16 B.t14 B.t15 B.t8 sky130_fd_pr__nfet_01v8 ad=5.4444 pd=28.7 as=0 ps=0 w=13.96 l=0.97
X1 VDD2.t3 VN.t0 VTAIL.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=2.3034 pd=14.29 as=5.4444 ps=28.7 w=13.96 l=0.97
X2 B.t13 B.t11 B.t12 B.t4 sky130_fd_pr__nfet_01v8 ad=5.4444 pd=28.7 as=0 ps=0 w=13.96 l=0.97
X3 VTAIL.t7 VP.t0 VDD1.t3 B.t17 sky130_fd_pr__nfet_01v8 ad=5.4444 pd=28.7 as=2.3034 ps=14.29 w=13.96 l=0.97
X4 VDD2.t2 VN.t1 VTAIL.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=2.3034 pd=14.29 as=5.4444 ps=28.7 w=13.96 l=0.97
X5 VDD1.t2 VP.t1 VTAIL.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=2.3034 pd=14.29 as=5.4444 ps=28.7 w=13.96 l=0.97
X6 B.t10 B.t7 B.t9 B.t8 sky130_fd_pr__nfet_01v8 ad=5.4444 pd=28.7 as=0 ps=0 w=13.96 l=0.97
X7 VDD1.t1 VP.t2 VTAIL.t5 B.t1 sky130_fd_pr__nfet_01v8 ad=2.3034 pd=14.29 as=5.4444 ps=28.7 w=13.96 l=0.97
X8 VTAIL.t0 VN.t2 VDD2.t1 B.t17 sky130_fd_pr__nfet_01v8 ad=5.4444 pd=28.7 as=2.3034 ps=14.29 w=13.96 l=0.97
X9 B.t6 B.t3 B.t5 B.t4 sky130_fd_pr__nfet_01v8 ad=5.4444 pd=28.7 as=0 ps=0 w=13.96 l=0.97
X10 VTAIL.t1 VN.t3 VDD2.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=5.4444 pd=28.7 as=2.3034 ps=14.29 w=13.96 l=0.97
X11 VTAIL.t4 VP.t3 VDD1.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=5.4444 pd=28.7 as=2.3034 ps=14.29 w=13.96 l=0.97
R0 B.n685 B.n684 585
R1 B.n298 B.n90 585
R2 B.n297 B.n296 585
R3 B.n295 B.n294 585
R4 B.n293 B.n292 585
R5 B.n291 B.n290 585
R6 B.n289 B.n288 585
R7 B.n287 B.n286 585
R8 B.n285 B.n284 585
R9 B.n283 B.n282 585
R10 B.n281 B.n280 585
R11 B.n279 B.n278 585
R12 B.n277 B.n276 585
R13 B.n275 B.n274 585
R14 B.n273 B.n272 585
R15 B.n271 B.n270 585
R16 B.n269 B.n268 585
R17 B.n267 B.n266 585
R18 B.n265 B.n264 585
R19 B.n263 B.n262 585
R20 B.n261 B.n260 585
R21 B.n259 B.n258 585
R22 B.n257 B.n256 585
R23 B.n255 B.n254 585
R24 B.n253 B.n252 585
R25 B.n251 B.n250 585
R26 B.n249 B.n248 585
R27 B.n247 B.n246 585
R28 B.n245 B.n244 585
R29 B.n243 B.n242 585
R30 B.n241 B.n240 585
R31 B.n239 B.n238 585
R32 B.n237 B.n236 585
R33 B.n235 B.n234 585
R34 B.n233 B.n232 585
R35 B.n231 B.n230 585
R36 B.n229 B.n228 585
R37 B.n227 B.n226 585
R38 B.n225 B.n224 585
R39 B.n223 B.n222 585
R40 B.n221 B.n220 585
R41 B.n219 B.n218 585
R42 B.n217 B.n216 585
R43 B.n215 B.n214 585
R44 B.n213 B.n212 585
R45 B.n211 B.n210 585
R46 B.n209 B.n208 585
R47 B.n206 B.n205 585
R48 B.n204 B.n203 585
R49 B.n202 B.n201 585
R50 B.n200 B.n199 585
R51 B.n198 B.n197 585
R52 B.n196 B.n195 585
R53 B.n194 B.n193 585
R54 B.n192 B.n191 585
R55 B.n190 B.n189 585
R56 B.n188 B.n187 585
R57 B.n185 B.n184 585
R58 B.n183 B.n182 585
R59 B.n181 B.n180 585
R60 B.n179 B.n178 585
R61 B.n177 B.n176 585
R62 B.n175 B.n174 585
R63 B.n173 B.n172 585
R64 B.n171 B.n170 585
R65 B.n169 B.n168 585
R66 B.n167 B.n166 585
R67 B.n165 B.n164 585
R68 B.n163 B.n162 585
R69 B.n161 B.n160 585
R70 B.n159 B.n158 585
R71 B.n157 B.n156 585
R72 B.n155 B.n154 585
R73 B.n153 B.n152 585
R74 B.n151 B.n150 585
R75 B.n149 B.n148 585
R76 B.n147 B.n146 585
R77 B.n145 B.n144 585
R78 B.n143 B.n142 585
R79 B.n141 B.n140 585
R80 B.n139 B.n138 585
R81 B.n137 B.n136 585
R82 B.n135 B.n134 585
R83 B.n133 B.n132 585
R84 B.n131 B.n130 585
R85 B.n129 B.n128 585
R86 B.n127 B.n126 585
R87 B.n125 B.n124 585
R88 B.n123 B.n122 585
R89 B.n121 B.n120 585
R90 B.n119 B.n118 585
R91 B.n117 B.n116 585
R92 B.n115 B.n114 585
R93 B.n113 B.n112 585
R94 B.n111 B.n110 585
R95 B.n109 B.n108 585
R96 B.n107 B.n106 585
R97 B.n105 B.n104 585
R98 B.n103 B.n102 585
R99 B.n101 B.n100 585
R100 B.n99 B.n98 585
R101 B.n97 B.n96 585
R102 B.n39 B.n38 585
R103 B.n690 B.n689 585
R104 B.n683 B.n91 585
R105 B.n91 B.n36 585
R106 B.n682 B.n35 585
R107 B.n694 B.n35 585
R108 B.n681 B.n34 585
R109 B.n695 B.n34 585
R110 B.n680 B.n33 585
R111 B.n696 B.n33 585
R112 B.n679 B.n678 585
R113 B.n678 B.n29 585
R114 B.n677 B.n28 585
R115 B.n702 B.n28 585
R116 B.n676 B.n27 585
R117 B.n703 B.n27 585
R118 B.n675 B.n26 585
R119 B.n704 B.n26 585
R120 B.n674 B.n673 585
R121 B.n673 B.n22 585
R122 B.n672 B.n21 585
R123 B.n710 B.n21 585
R124 B.n671 B.n20 585
R125 B.n711 B.n20 585
R126 B.n670 B.n19 585
R127 B.n712 B.n19 585
R128 B.n669 B.n668 585
R129 B.n668 B.n18 585
R130 B.n667 B.n14 585
R131 B.n718 B.n14 585
R132 B.n666 B.n13 585
R133 B.n719 B.n13 585
R134 B.n665 B.n12 585
R135 B.n720 B.n12 585
R136 B.n664 B.n663 585
R137 B.n663 B.n662 585
R138 B.n661 B.n660 585
R139 B.n661 B.n8 585
R140 B.n659 B.n7 585
R141 B.n727 B.n7 585
R142 B.n658 B.n6 585
R143 B.n728 B.n6 585
R144 B.n657 B.n5 585
R145 B.n729 B.n5 585
R146 B.n656 B.n655 585
R147 B.n655 B.n4 585
R148 B.n654 B.n299 585
R149 B.n654 B.n653 585
R150 B.n644 B.n300 585
R151 B.n301 B.n300 585
R152 B.n646 B.n645 585
R153 B.n647 B.n646 585
R154 B.n643 B.n306 585
R155 B.n306 B.n305 585
R156 B.n642 B.n641 585
R157 B.n641 B.n640 585
R158 B.n308 B.n307 585
R159 B.n633 B.n308 585
R160 B.n632 B.n631 585
R161 B.n634 B.n632 585
R162 B.n630 B.n313 585
R163 B.n313 B.n312 585
R164 B.n629 B.n628 585
R165 B.n628 B.n627 585
R166 B.n315 B.n314 585
R167 B.n316 B.n315 585
R168 B.n620 B.n619 585
R169 B.n621 B.n620 585
R170 B.n618 B.n321 585
R171 B.n321 B.n320 585
R172 B.n617 B.n616 585
R173 B.n616 B.n615 585
R174 B.n323 B.n322 585
R175 B.n324 B.n323 585
R176 B.n608 B.n607 585
R177 B.n609 B.n608 585
R178 B.n606 B.n329 585
R179 B.n329 B.n328 585
R180 B.n605 B.n604 585
R181 B.n604 B.n603 585
R182 B.n331 B.n330 585
R183 B.n332 B.n331 585
R184 B.n599 B.n598 585
R185 B.n335 B.n334 585
R186 B.n595 B.n594 585
R187 B.n596 B.n595 585
R188 B.n593 B.n387 585
R189 B.n592 B.n591 585
R190 B.n590 B.n589 585
R191 B.n588 B.n587 585
R192 B.n586 B.n585 585
R193 B.n584 B.n583 585
R194 B.n582 B.n581 585
R195 B.n580 B.n579 585
R196 B.n578 B.n577 585
R197 B.n576 B.n575 585
R198 B.n574 B.n573 585
R199 B.n572 B.n571 585
R200 B.n570 B.n569 585
R201 B.n568 B.n567 585
R202 B.n566 B.n565 585
R203 B.n564 B.n563 585
R204 B.n562 B.n561 585
R205 B.n560 B.n559 585
R206 B.n558 B.n557 585
R207 B.n556 B.n555 585
R208 B.n554 B.n553 585
R209 B.n552 B.n551 585
R210 B.n550 B.n549 585
R211 B.n548 B.n547 585
R212 B.n546 B.n545 585
R213 B.n544 B.n543 585
R214 B.n542 B.n541 585
R215 B.n540 B.n539 585
R216 B.n538 B.n537 585
R217 B.n536 B.n535 585
R218 B.n534 B.n533 585
R219 B.n532 B.n531 585
R220 B.n530 B.n529 585
R221 B.n528 B.n527 585
R222 B.n526 B.n525 585
R223 B.n524 B.n523 585
R224 B.n522 B.n521 585
R225 B.n520 B.n519 585
R226 B.n518 B.n517 585
R227 B.n516 B.n515 585
R228 B.n514 B.n513 585
R229 B.n512 B.n511 585
R230 B.n510 B.n509 585
R231 B.n508 B.n507 585
R232 B.n506 B.n505 585
R233 B.n504 B.n503 585
R234 B.n502 B.n501 585
R235 B.n500 B.n499 585
R236 B.n498 B.n497 585
R237 B.n496 B.n495 585
R238 B.n494 B.n493 585
R239 B.n492 B.n491 585
R240 B.n490 B.n489 585
R241 B.n488 B.n487 585
R242 B.n486 B.n485 585
R243 B.n484 B.n483 585
R244 B.n482 B.n481 585
R245 B.n480 B.n479 585
R246 B.n478 B.n477 585
R247 B.n476 B.n475 585
R248 B.n474 B.n473 585
R249 B.n472 B.n471 585
R250 B.n470 B.n469 585
R251 B.n468 B.n467 585
R252 B.n466 B.n465 585
R253 B.n464 B.n463 585
R254 B.n462 B.n461 585
R255 B.n460 B.n459 585
R256 B.n458 B.n457 585
R257 B.n456 B.n455 585
R258 B.n454 B.n453 585
R259 B.n452 B.n451 585
R260 B.n450 B.n449 585
R261 B.n448 B.n447 585
R262 B.n446 B.n445 585
R263 B.n444 B.n443 585
R264 B.n442 B.n441 585
R265 B.n440 B.n439 585
R266 B.n438 B.n437 585
R267 B.n436 B.n435 585
R268 B.n434 B.n433 585
R269 B.n432 B.n431 585
R270 B.n430 B.n429 585
R271 B.n428 B.n427 585
R272 B.n426 B.n425 585
R273 B.n424 B.n423 585
R274 B.n422 B.n421 585
R275 B.n420 B.n419 585
R276 B.n418 B.n417 585
R277 B.n416 B.n415 585
R278 B.n414 B.n413 585
R279 B.n412 B.n411 585
R280 B.n410 B.n409 585
R281 B.n408 B.n407 585
R282 B.n406 B.n405 585
R283 B.n404 B.n403 585
R284 B.n402 B.n401 585
R285 B.n400 B.n399 585
R286 B.n398 B.n397 585
R287 B.n396 B.n395 585
R288 B.n394 B.n386 585
R289 B.n596 B.n386 585
R290 B.n600 B.n333 585
R291 B.n333 B.n332 585
R292 B.n602 B.n601 585
R293 B.n603 B.n602 585
R294 B.n327 B.n326 585
R295 B.n328 B.n327 585
R296 B.n611 B.n610 585
R297 B.n610 B.n609 585
R298 B.n612 B.n325 585
R299 B.n325 B.n324 585
R300 B.n614 B.n613 585
R301 B.n615 B.n614 585
R302 B.n319 B.n318 585
R303 B.n320 B.n319 585
R304 B.n623 B.n622 585
R305 B.n622 B.n621 585
R306 B.n624 B.n317 585
R307 B.n317 B.n316 585
R308 B.n626 B.n625 585
R309 B.n627 B.n626 585
R310 B.n311 B.n310 585
R311 B.n312 B.n311 585
R312 B.n636 B.n635 585
R313 B.n635 B.n634 585
R314 B.n637 B.n309 585
R315 B.n633 B.n309 585
R316 B.n639 B.n638 585
R317 B.n640 B.n639 585
R318 B.n304 B.n303 585
R319 B.n305 B.n304 585
R320 B.n649 B.n648 585
R321 B.n648 B.n647 585
R322 B.n650 B.n302 585
R323 B.n302 B.n301 585
R324 B.n652 B.n651 585
R325 B.n653 B.n652 585
R326 B.n3 B.n0 585
R327 B.n4 B.n3 585
R328 B.n726 B.n1 585
R329 B.n727 B.n726 585
R330 B.n725 B.n724 585
R331 B.n725 B.n8 585
R332 B.n723 B.n9 585
R333 B.n662 B.n9 585
R334 B.n722 B.n721 585
R335 B.n721 B.n720 585
R336 B.n11 B.n10 585
R337 B.n719 B.n11 585
R338 B.n717 B.n716 585
R339 B.n718 B.n717 585
R340 B.n715 B.n15 585
R341 B.n18 B.n15 585
R342 B.n714 B.n713 585
R343 B.n713 B.n712 585
R344 B.n17 B.n16 585
R345 B.n711 B.n17 585
R346 B.n709 B.n708 585
R347 B.n710 B.n709 585
R348 B.n707 B.n23 585
R349 B.n23 B.n22 585
R350 B.n706 B.n705 585
R351 B.n705 B.n704 585
R352 B.n25 B.n24 585
R353 B.n703 B.n25 585
R354 B.n701 B.n700 585
R355 B.n702 B.n701 585
R356 B.n699 B.n30 585
R357 B.n30 B.n29 585
R358 B.n698 B.n697 585
R359 B.n697 B.n696 585
R360 B.n32 B.n31 585
R361 B.n695 B.n32 585
R362 B.n693 B.n692 585
R363 B.n694 B.n693 585
R364 B.n691 B.n37 585
R365 B.n37 B.n36 585
R366 B.n730 B.n729 585
R367 B.n728 B.n2 585
R368 B.n94 B.t11 549.561
R369 B.n92 B.t3 549.561
R370 B.n391 B.t7 549.561
R371 B.n388 B.t14 549.561
R372 B.n689 B.n37 540.549
R373 B.n685 B.n91 540.549
R374 B.n386 B.n331 540.549
R375 B.n598 B.n333 540.549
R376 B.n92 B.t5 340.805
R377 B.n391 B.t10 340.805
R378 B.n94 B.t12 340.805
R379 B.n388 B.t16 340.805
R380 B.n93 B.t6 315.594
R381 B.n392 B.t9 315.594
R382 B.n95 B.t13 315.594
R383 B.n389 B.t15 315.594
R384 B.n687 B.n686 256.663
R385 B.n687 B.n89 256.663
R386 B.n687 B.n88 256.663
R387 B.n687 B.n87 256.663
R388 B.n687 B.n86 256.663
R389 B.n687 B.n85 256.663
R390 B.n687 B.n84 256.663
R391 B.n687 B.n83 256.663
R392 B.n687 B.n82 256.663
R393 B.n687 B.n81 256.663
R394 B.n687 B.n80 256.663
R395 B.n687 B.n79 256.663
R396 B.n687 B.n78 256.663
R397 B.n687 B.n77 256.663
R398 B.n687 B.n76 256.663
R399 B.n687 B.n75 256.663
R400 B.n687 B.n74 256.663
R401 B.n687 B.n73 256.663
R402 B.n687 B.n72 256.663
R403 B.n687 B.n71 256.663
R404 B.n687 B.n70 256.663
R405 B.n687 B.n69 256.663
R406 B.n687 B.n68 256.663
R407 B.n687 B.n67 256.663
R408 B.n687 B.n66 256.663
R409 B.n687 B.n65 256.663
R410 B.n687 B.n64 256.663
R411 B.n687 B.n63 256.663
R412 B.n687 B.n62 256.663
R413 B.n687 B.n61 256.663
R414 B.n687 B.n60 256.663
R415 B.n687 B.n59 256.663
R416 B.n687 B.n58 256.663
R417 B.n687 B.n57 256.663
R418 B.n687 B.n56 256.663
R419 B.n687 B.n55 256.663
R420 B.n687 B.n54 256.663
R421 B.n687 B.n53 256.663
R422 B.n687 B.n52 256.663
R423 B.n687 B.n51 256.663
R424 B.n687 B.n50 256.663
R425 B.n687 B.n49 256.663
R426 B.n687 B.n48 256.663
R427 B.n687 B.n47 256.663
R428 B.n687 B.n46 256.663
R429 B.n687 B.n45 256.663
R430 B.n687 B.n44 256.663
R431 B.n687 B.n43 256.663
R432 B.n687 B.n42 256.663
R433 B.n687 B.n41 256.663
R434 B.n687 B.n40 256.663
R435 B.n688 B.n687 256.663
R436 B.n597 B.n596 256.663
R437 B.n596 B.n336 256.663
R438 B.n596 B.n337 256.663
R439 B.n596 B.n338 256.663
R440 B.n596 B.n339 256.663
R441 B.n596 B.n340 256.663
R442 B.n596 B.n341 256.663
R443 B.n596 B.n342 256.663
R444 B.n596 B.n343 256.663
R445 B.n596 B.n344 256.663
R446 B.n596 B.n345 256.663
R447 B.n596 B.n346 256.663
R448 B.n596 B.n347 256.663
R449 B.n596 B.n348 256.663
R450 B.n596 B.n349 256.663
R451 B.n596 B.n350 256.663
R452 B.n596 B.n351 256.663
R453 B.n596 B.n352 256.663
R454 B.n596 B.n353 256.663
R455 B.n596 B.n354 256.663
R456 B.n596 B.n355 256.663
R457 B.n596 B.n356 256.663
R458 B.n596 B.n357 256.663
R459 B.n596 B.n358 256.663
R460 B.n596 B.n359 256.663
R461 B.n596 B.n360 256.663
R462 B.n596 B.n361 256.663
R463 B.n596 B.n362 256.663
R464 B.n596 B.n363 256.663
R465 B.n596 B.n364 256.663
R466 B.n596 B.n365 256.663
R467 B.n596 B.n366 256.663
R468 B.n596 B.n367 256.663
R469 B.n596 B.n368 256.663
R470 B.n596 B.n369 256.663
R471 B.n596 B.n370 256.663
R472 B.n596 B.n371 256.663
R473 B.n596 B.n372 256.663
R474 B.n596 B.n373 256.663
R475 B.n596 B.n374 256.663
R476 B.n596 B.n375 256.663
R477 B.n596 B.n376 256.663
R478 B.n596 B.n377 256.663
R479 B.n596 B.n378 256.663
R480 B.n596 B.n379 256.663
R481 B.n596 B.n380 256.663
R482 B.n596 B.n381 256.663
R483 B.n596 B.n382 256.663
R484 B.n596 B.n383 256.663
R485 B.n596 B.n384 256.663
R486 B.n596 B.n385 256.663
R487 B.n732 B.n731 256.663
R488 B.n96 B.n39 163.367
R489 B.n100 B.n99 163.367
R490 B.n104 B.n103 163.367
R491 B.n108 B.n107 163.367
R492 B.n112 B.n111 163.367
R493 B.n116 B.n115 163.367
R494 B.n120 B.n119 163.367
R495 B.n124 B.n123 163.367
R496 B.n128 B.n127 163.367
R497 B.n132 B.n131 163.367
R498 B.n136 B.n135 163.367
R499 B.n140 B.n139 163.367
R500 B.n144 B.n143 163.367
R501 B.n148 B.n147 163.367
R502 B.n152 B.n151 163.367
R503 B.n156 B.n155 163.367
R504 B.n160 B.n159 163.367
R505 B.n164 B.n163 163.367
R506 B.n168 B.n167 163.367
R507 B.n172 B.n171 163.367
R508 B.n176 B.n175 163.367
R509 B.n180 B.n179 163.367
R510 B.n184 B.n183 163.367
R511 B.n189 B.n188 163.367
R512 B.n193 B.n192 163.367
R513 B.n197 B.n196 163.367
R514 B.n201 B.n200 163.367
R515 B.n205 B.n204 163.367
R516 B.n210 B.n209 163.367
R517 B.n214 B.n213 163.367
R518 B.n218 B.n217 163.367
R519 B.n222 B.n221 163.367
R520 B.n226 B.n225 163.367
R521 B.n230 B.n229 163.367
R522 B.n234 B.n233 163.367
R523 B.n238 B.n237 163.367
R524 B.n242 B.n241 163.367
R525 B.n246 B.n245 163.367
R526 B.n250 B.n249 163.367
R527 B.n254 B.n253 163.367
R528 B.n258 B.n257 163.367
R529 B.n262 B.n261 163.367
R530 B.n266 B.n265 163.367
R531 B.n270 B.n269 163.367
R532 B.n274 B.n273 163.367
R533 B.n278 B.n277 163.367
R534 B.n282 B.n281 163.367
R535 B.n286 B.n285 163.367
R536 B.n290 B.n289 163.367
R537 B.n294 B.n293 163.367
R538 B.n296 B.n90 163.367
R539 B.n604 B.n331 163.367
R540 B.n604 B.n329 163.367
R541 B.n608 B.n329 163.367
R542 B.n608 B.n323 163.367
R543 B.n616 B.n323 163.367
R544 B.n616 B.n321 163.367
R545 B.n620 B.n321 163.367
R546 B.n620 B.n315 163.367
R547 B.n628 B.n315 163.367
R548 B.n628 B.n313 163.367
R549 B.n632 B.n313 163.367
R550 B.n632 B.n308 163.367
R551 B.n641 B.n308 163.367
R552 B.n641 B.n306 163.367
R553 B.n646 B.n306 163.367
R554 B.n646 B.n300 163.367
R555 B.n654 B.n300 163.367
R556 B.n655 B.n654 163.367
R557 B.n655 B.n5 163.367
R558 B.n6 B.n5 163.367
R559 B.n7 B.n6 163.367
R560 B.n661 B.n7 163.367
R561 B.n663 B.n661 163.367
R562 B.n663 B.n12 163.367
R563 B.n13 B.n12 163.367
R564 B.n14 B.n13 163.367
R565 B.n668 B.n14 163.367
R566 B.n668 B.n19 163.367
R567 B.n20 B.n19 163.367
R568 B.n21 B.n20 163.367
R569 B.n673 B.n21 163.367
R570 B.n673 B.n26 163.367
R571 B.n27 B.n26 163.367
R572 B.n28 B.n27 163.367
R573 B.n678 B.n28 163.367
R574 B.n678 B.n33 163.367
R575 B.n34 B.n33 163.367
R576 B.n35 B.n34 163.367
R577 B.n91 B.n35 163.367
R578 B.n595 B.n335 163.367
R579 B.n595 B.n387 163.367
R580 B.n591 B.n590 163.367
R581 B.n587 B.n586 163.367
R582 B.n583 B.n582 163.367
R583 B.n579 B.n578 163.367
R584 B.n575 B.n574 163.367
R585 B.n571 B.n570 163.367
R586 B.n567 B.n566 163.367
R587 B.n563 B.n562 163.367
R588 B.n559 B.n558 163.367
R589 B.n555 B.n554 163.367
R590 B.n551 B.n550 163.367
R591 B.n547 B.n546 163.367
R592 B.n543 B.n542 163.367
R593 B.n539 B.n538 163.367
R594 B.n535 B.n534 163.367
R595 B.n531 B.n530 163.367
R596 B.n527 B.n526 163.367
R597 B.n523 B.n522 163.367
R598 B.n519 B.n518 163.367
R599 B.n515 B.n514 163.367
R600 B.n511 B.n510 163.367
R601 B.n507 B.n506 163.367
R602 B.n503 B.n502 163.367
R603 B.n499 B.n498 163.367
R604 B.n495 B.n494 163.367
R605 B.n491 B.n490 163.367
R606 B.n487 B.n486 163.367
R607 B.n483 B.n482 163.367
R608 B.n479 B.n478 163.367
R609 B.n475 B.n474 163.367
R610 B.n471 B.n470 163.367
R611 B.n467 B.n466 163.367
R612 B.n463 B.n462 163.367
R613 B.n459 B.n458 163.367
R614 B.n455 B.n454 163.367
R615 B.n451 B.n450 163.367
R616 B.n447 B.n446 163.367
R617 B.n443 B.n442 163.367
R618 B.n439 B.n438 163.367
R619 B.n435 B.n434 163.367
R620 B.n431 B.n430 163.367
R621 B.n427 B.n426 163.367
R622 B.n423 B.n422 163.367
R623 B.n419 B.n418 163.367
R624 B.n415 B.n414 163.367
R625 B.n411 B.n410 163.367
R626 B.n407 B.n406 163.367
R627 B.n403 B.n402 163.367
R628 B.n399 B.n398 163.367
R629 B.n395 B.n386 163.367
R630 B.n602 B.n333 163.367
R631 B.n602 B.n327 163.367
R632 B.n610 B.n327 163.367
R633 B.n610 B.n325 163.367
R634 B.n614 B.n325 163.367
R635 B.n614 B.n319 163.367
R636 B.n622 B.n319 163.367
R637 B.n622 B.n317 163.367
R638 B.n626 B.n317 163.367
R639 B.n626 B.n311 163.367
R640 B.n635 B.n311 163.367
R641 B.n635 B.n309 163.367
R642 B.n639 B.n309 163.367
R643 B.n639 B.n304 163.367
R644 B.n648 B.n304 163.367
R645 B.n648 B.n302 163.367
R646 B.n652 B.n302 163.367
R647 B.n652 B.n3 163.367
R648 B.n730 B.n3 163.367
R649 B.n726 B.n2 163.367
R650 B.n726 B.n725 163.367
R651 B.n725 B.n9 163.367
R652 B.n721 B.n9 163.367
R653 B.n721 B.n11 163.367
R654 B.n717 B.n11 163.367
R655 B.n717 B.n15 163.367
R656 B.n713 B.n15 163.367
R657 B.n713 B.n17 163.367
R658 B.n709 B.n17 163.367
R659 B.n709 B.n23 163.367
R660 B.n705 B.n23 163.367
R661 B.n705 B.n25 163.367
R662 B.n701 B.n25 163.367
R663 B.n701 B.n30 163.367
R664 B.n697 B.n30 163.367
R665 B.n697 B.n32 163.367
R666 B.n693 B.n32 163.367
R667 B.n693 B.n37 163.367
R668 B.n596 B.n332 73.7723
R669 B.n687 B.n36 73.7723
R670 B.n689 B.n688 71.676
R671 B.n96 B.n40 71.676
R672 B.n100 B.n41 71.676
R673 B.n104 B.n42 71.676
R674 B.n108 B.n43 71.676
R675 B.n112 B.n44 71.676
R676 B.n116 B.n45 71.676
R677 B.n120 B.n46 71.676
R678 B.n124 B.n47 71.676
R679 B.n128 B.n48 71.676
R680 B.n132 B.n49 71.676
R681 B.n136 B.n50 71.676
R682 B.n140 B.n51 71.676
R683 B.n144 B.n52 71.676
R684 B.n148 B.n53 71.676
R685 B.n152 B.n54 71.676
R686 B.n156 B.n55 71.676
R687 B.n160 B.n56 71.676
R688 B.n164 B.n57 71.676
R689 B.n168 B.n58 71.676
R690 B.n172 B.n59 71.676
R691 B.n176 B.n60 71.676
R692 B.n180 B.n61 71.676
R693 B.n184 B.n62 71.676
R694 B.n189 B.n63 71.676
R695 B.n193 B.n64 71.676
R696 B.n197 B.n65 71.676
R697 B.n201 B.n66 71.676
R698 B.n205 B.n67 71.676
R699 B.n210 B.n68 71.676
R700 B.n214 B.n69 71.676
R701 B.n218 B.n70 71.676
R702 B.n222 B.n71 71.676
R703 B.n226 B.n72 71.676
R704 B.n230 B.n73 71.676
R705 B.n234 B.n74 71.676
R706 B.n238 B.n75 71.676
R707 B.n242 B.n76 71.676
R708 B.n246 B.n77 71.676
R709 B.n250 B.n78 71.676
R710 B.n254 B.n79 71.676
R711 B.n258 B.n80 71.676
R712 B.n262 B.n81 71.676
R713 B.n266 B.n82 71.676
R714 B.n270 B.n83 71.676
R715 B.n274 B.n84 71.676
R716 B.n278 B.n85 71.676
R717 B.n282 B.n86 71.676
R718 B.n286 B.n87 71.676
R719 B.n290 B.n88 71.676
R720 B.n294 B.n89 71.676
R721 B.n686 B.n90 71.676
R722 B.n686 B.n685 71.676
R723 B.n296 B.n89 71.676
R724 B.n293 B.n88 71.676
R725 B.n289 B.n87 71.676
R726 B.n285 B.n86 71.676
R727 B.n281 B.n85 71.676
R728 B.n277 B.n84 71.676
R729 B.n273 B.n83 71.676
R730 B.n269 B.n82 71.676
R731 B.n265 B.n81 71.676
R732 B.n261 B.n80 71.676
R733 B.n257 B.n79 71.676
R734 B.n253 B.n78 71.676
R735 B.n249 B.n77 71.676
R736 B.n245 B.n76 71.676
R737 B.n241 B.n75 71.676
R738 B.n237 B.n74 71.676
R739 B.n233 B.n73 71.676
R740 B.n229 B.n72 71.676
R741 B.n225 B.n71 71.676
R742 B.n221 B.n70 71.676
R743 B.n217 B.n69 71.676
R744 B.n213 B.n68 71.676
R745 B.n209 B.n67 71.676
R746 B.n204 B.n66 71.676
R747 B.n200 B.n65 71.676
R748 B.n196 B.n64 71.676
R749 B.n192 B.n63 71.676
R750 B.n188 B.n62 71.676
R751 B.n183 B.n61 71.676
R752 B.n179 B.n60 71.676
R753 B.n175 B.n59 71.676
R754 B.n171 B.n58 71.676
R755 B.n167 B.n57 71.676
R756 B.n163 B.n56 71.676
R757 B.n159 B.n55 71.676
R758 B.n155 B.n54 71.676
R759 B.n151 B.n53 71.676
R760 B.n147 B.n52 71.676
R761 B.n143 B.n51 71.676
R762 B.n139 B.n50 71.676
R763 B.n135 B.n49 71.676
R764 B.n131 B.n48 71.676
R765 B.n127 B.n47 71.676
R766 B.n123 B.n46 71.676
R767 B.n119 B.n45 71.676
R768 B.n115 B.n44 71.676
R769 B.n111 B.n43 71.676
R770 B.n107 B.n42 71.676
R771 B.n103 B.n41 71.676
R772 B.n99 B.n40 71.676
R773 B.n688 B.n39 71.676
R774 B.n598 B.n597 71.676
R775 B.n387 B.n336 71.676
R776 B.n590 B.n337 71.676
R777 B.n586 B.n338 71.676
R778 B.n582 B.n339 71.676
R779 B.n578 B.n340 71.676
R780 B.n574 B.n341 71.676
R781 B.n570 B.n342 71.676
R782 B.n566 B.n343 71.676
R783 B.n562 B.n344 71.676
R784 B.n558 B.n345 71.676
R785 B.n554 B.n346 71.676
R786 B.n550 B.n347 71.676
R787 B.n546 B.n348 71.676
R788 B.n542 B.n349 71.676
R789 B.n538 B.n350 71.676
R790 B.n534 B.n351 71.676
R791 B.n530 B.n352 71.676
R792 B.n526 B.n353 71.676
R793 B.n522 B.n354 71.676
R794 B.n518 B.n355 71.676
R795 B.n514 B.n356 71.676
R796 B.n510 B.n357 71.676
R797 B.n506 B.n358 71.676
R798 B.n502 B.n359 71.676
R799 B.n498 B.n360 71.676
R800 B.n494 B.n361 71.676
R801 B.n490 B.n362 71.676
R802 B.n486 B.n363 71.676
R803 B.n482 B.n364 71.676
R804 B.n478 B.n365 71.676
R805 B.n474 B.n366 71.676
R806 B.n470 B.n367 71.676
R807 B.n466 B.n368 71.676
R808 B.n462 B.n369 71.676
R809 B.n458 B.n370 71.676
R810 B.n454 B.n371 71.676
R811 B.n450 B.n372 71.676
R812 B.n446 B.n373 71.676
R813 B.n442 B.n374 71.676
R814 B.n438 B.n375 71.676
R815 B.n434 B.n376 71.676
R816 B.n430 B.n377 71.676
R817 B.n426 B.n378 71.676
R818 B.n422 B.n379 71.676
R819 B.n418 B.n380 71.676
R820 B.n414 B.n381 71.676
R821 B.n410 B.n382 71.676
R822 B.n406 B.n383 71.676
R823 B.n402 B.n384 71.676
R824 B.n398 B.n385 71.676
R825 B.n597 B.n335 71.676
R826 B.n591 B.n336 71.676
R827 B.n587 B.n337 71.676
R828 B.n583 B.n338 71.676
R829 B.n579 B.n339 71.676
R830 B.n575 B.n340 71.676
R831 B.n571 B.n341 71.676
R832 B.n567 B.n342 71.676
R833 B.n563 B.n343 71.676
R834 B.n559 B.n344 71.676
R835 B.n555 B.n345 71.676
R836 B.n551 B.n346 71.676
R837 B.n547 B.n347 71.676
R838 B.n543 B.n348 71.676
R839 B.n539 B.n349 71.676
R840 B.n535 B.n350 71.676
R841 B.n531 B.n351 71.676
R842 B.n527 B.n352 71.676
R843 B.n523 B.n353 71.676
R844 B.n519 B.n354 71.676
R845 B.n515 B.n355 71.676
R846 B.n511 B.n356 71.676
R847 B.n507 B.n357 71.676
R848 B.n503 B.n358 71.676
R849 B.n499 B.n359 71.676
R850 B.n495 B.n360 71.676
R851 B.n491 B.n361 71.676
R852 B.n487 B.n362 71.676
R853 B.n483 B.n363 71.676
R854 B.n479 B.n364 71.676
R855 B.n475 B.n365 71.676
R856 B.n471 B.n366 71.676
R857 B.n467 B.n367 71.676
R858 B.n463 B.n368 71.676
R859 B.n459 B.n369 71.676
R860 B.n455 B.n370 71.676
R861 B.n451 B.n371 71.676
R862 B.n447 B.n372 71.676
R863 B.n443 B.n373 71.676
R864 B.n439 B.n374 71.676
R865 B.n435 B.n375 71.676
R866 B.n431 B.n376 71.676
R867 B.n427 B.n377 71.676
R868 B.n423 B.n378 71.676
R869 B.n419 B.n379 71.676
R870 B.n415 B.n380 71.676
R871 B.n411 B.n381 71.676
R872 B.n407 B.n382 71.676
R873 B.n403 B.n383 71.676
R874 B.n399 B.n384 71.676
R875 B.n395 B.n385 71.676
R876 B.n731 B.n730 71.676
R877 B.n731 B.n2 71.676
R878 B.n186 B.n95 59.5399
R879 B.n207 B.n93 59.5399
R880 B.n393 B.n392 59.5399
R881 B.n390 B.n389 59.5399
R882 B.n603 B.n332 38.8879
R883 B.n603 B.n328 38.8879
R884 B.n609 B.n328 38.8879
R885 B.n609 B.n324 38.8879
R886 B.n615 B.n324 38.8879
R887 B.n621 B.n320 38.8879
R888 B.n621 B.n316 38.8879
R889 B.n627 B.n316 38.8879
R890 B.n627 B.n312 38.8879
R891 B.n634 B.n312 38.8879
R892 B.n634 B.n633 38.8879
R893 B.n640 B.n305 38.8879
R894 B.n647 B.n305 38.8879
R895 B.n653 B.n301 38.8879
R896 B.n653 B.n4 38.8879
R897 B.n729 B.n4 38.8879
R898 B.n729 B.n728 38.8879
R899 B.n728 B.n727 38.8879
R900 B.n727 B.n8 38.8879
R901 B.n662 B.n8 38.8879
R902 B.n720 B.n719 38.8879
R903 B.n719 B.n718 38.8879
R904 B.n712 B.n18 38.8879
R905 B.n712 B.n711 38.8879
R906 B.n711 B.n710 38.8879
R907 B.n710 B.n22 38.8879
R908 B.n704 B.n22 38.8879
R909 B.n704 B.n703 38.8879
R910 B.n702 B.n29 38.8879
R911 B.n696 B.n29 38.8879
R912 B.n696 B.n695 38.8879
R913 B.n695 B.n694 38.8879
R914 B.n694 B.n36 38.8879
R915 B.n647 B.t2 38.3161
R916 B.n720 B.t0 38.3161
R917 B.n600 B.n599 35.1225
R918 B.n394 B.n330 35.1225
R919 B.n691 B.n690 35.1225
R920 B.n684 B.n683 35.1224
R921 B.t8 B.n320 33.7411
R922 B.n703 B.t4 33.7411
R923 B.n640 B.t17 32.5973
R924 B.n718 B.t1 32.5973
R925 B.n95 B.n94 25.2126
R926 B.n93 B.n92 25.2126
R927 B.n392 B.n391 25.2126
R928 B.n389 B.n388 25.2126
R929 B B.n732 18.0485
R930 B.n601 B.n600 10.6151
R931 B.n601 B.n326 10.6151
R932 B.n611 B.n326 10.6151
R933 B.n612 B.n611 10.6151
R934 B.n613 B.n612 10.6151
R935 B.n613 B.n318 10.6151
R936 B.n623 B.n318 10.6151
R937 B.n624 B.n623 10.6151
R938 B.n625 B.n624 10.6151
R939 B.n625 B.n310 10.6151
R940 B.n636 B.n310 10.6151
R941 B.n637 B.n636 10.6151
R942 B.n638 B.n637 10.6151
R943 B.n638 B.n303 10.6151
R944 B.n649 B.n303 10.6151
R945 B.n650 B.n649 10.6151
R946 B.n651 B.n650 10.6151
R947 B.n651 B.n0 10.6151
R948 B.n599 B.n334 10.6151
R949 B.n594 B.n334 10.6151
R950 B.n594 B.n593 10.6151
R951 B.n593 B.n592 10.6151
R952 B.n592 B.n589 10.6151
R953 B.n589 B.n588 10.6151
R954 B.n588 B.n585 10.6151
R955 B.n585 B.n584 10.6151
R956 B.n584 B.n581 10.6151
R957 B.n581 B.n580 10.6151
R958 B.n580 B.n577 10.6151
R959 B.n577 B.n576 10.6151
R960 B.n576 B.n573 10.6151
R961 B.n573 B.n572 10.6151
R962 B.n572 B.n569 10.6151
R963 B.n569 B.n568 10.6151
R964 B.n568 B.n565 10.6151
R965 B.n565 B.n564 10.6151
R966 B.n564 B.n561 10.6151
R967 B.n561 B.n560 10.6151
R968 B.n560 B.n557 10.6151
R969 B.n557 B.n556 10.6151
R970 B.n556 B.n553 10.6151
R971 B.n553 B.n552 10.6151
R972 B.n552 B.n549 10.6151
R973 B.n549 B.n548 10.6151
R974 B.n548 B.n545 10.6151
R975 B.n545 B.n544 10.6151
R976 B.n544 B.n541 10.6151
R977 B.n541 B.n540 10.6151
R978 B.n540 B.n537 10.6151
R979 B.n537 B.n536 10.6151
R980 B.n536 B.n533 10.6151
R981 B.n533 B.n532 10.6151
R982 B.n532 B.n529 10.6151
R983 B.n529 B.n528 10.6151
R984 B.n528 B.n525 10.6151
R985 B.n525 B.n524 10.6151
R986 B.n524 B.n521 10.6151
R987 B.n521 B.n520 10.6151
R988 B.n520 B.n517 10.6151
R989 B.n517 B.n516 10.6151
R990 B.n516 B.n513 10.6151
R991 B.n513 B.n512 10.6151
R992 B.n512 B.n509 10.6151
R993 B.n509 B.n508 10.6151
R994 B.n505 B.n504 10.6151
R995 B.n504 B.n501 10.6151
R996 B.n501 B.n500 10.6151
R997 B.n500 B.n497 10.6151
R998 B.n497 B.n496 10.6151
R999 B.n496 B.n493 10.6151
R1000 B.n493 B.n492 10.6151
R1001 B.n492 B.n489 10.6151
R1002 B.n489 B.n488 10.6151
R1003 B.n485 B.n484 10.6151
R1004 B.n484 B.n481 10.6151
R1005 B.n481 B.n480 10.6151
R1006 B.n480 B.n477 10.6151
R1007 B.n477 B.n476 10.6151
R1008 B.n476 B.n473 10.6151
R1009 B.n473 B.n472 10.6151
R1010 B.n472 B.n469 10.6151
R1011 B.n469 B.n468 10.6151
R1012 B.n468 B.n465 10.6151
R1013 B.n465 B.n464 10.6151
R1014 B.n464 B.n461 10.6151
R1015 B.n461 B.n460 10.6151
R1016 B.n460 B.n457 10.6151
R1017 B.n457 B.n456 10.6151
R1018 B.n456 B.n453 10.6151
R1019 B.n453 B.n452 10.6151
R1020 B.n452 B.n449 10.6151
R1021 B.n449 B.n448 10.6151
R1022 B.n448 B.n445 10.6151
R1023 B.n445 B.n444 10.6151
R1024 B.n444 B.n441 10.6151
R1025 B.n441 B.n440 10.6151
R1026 B.n440 B.n437 10.6151
R1027 B.n437 B.n436 10.6151
R1028 B.n436 B.n433 10.6151
R1029 B.n433 B.n432 10.6151
R1030 B.n432 B.n429 10.6151
R1031 B.n429 B.n428 10.6151
R1032 B.n428 B.n425 10.6151
R1033 B.n425 B.n424 10.6151
R1034 B.n424 B.n421 10.6151
R1035 B.n421 B.n420 10.6151
R1036 B.n420 B.n417 10.6151
R1037 B.n417 B.n416 10.6151
R1038 B.n416 B.n413 10.6151
R1039 B.n413 B.n412 10.6151
R1040 B.n412 B.n409 10.6151
R1041 B.n409 B.n408 10.6151
R1042 B.n408 B.n405 10.6151
R1043 B.n405 B.n404 10.6151
R1044 B.n404 B.n401 10.6151
R1045 B.n401 B.n400 10.6151
R1046 B.n400 B.n397 10.6151
R1047 B.n397 B.n396 10.6151
R1048 B.n396 B.n394 10.6151
R1049 B.n605 B.n330 10.6151
R1050 B.n606 B.n605 10.6151
R1051 B.n607 B.n606 10.6151
R1052 B.n607 B.n322 10.6151
R1053 B.n617 B.n322 10.6151
R1054 B.n618 B.n617 10.6151
R1055 B.n619 B.n618 10.6151
R1056 B.n619 B.n314 10.6151
R1057 B.n629 B.n314 10.6151
R1058 B.n630 B.n629 10.6151
R1059 B.n631 B.n630 10.6151
R1060 B.n631 B.n307 10.6151
R1061 B.n642 B.n307 10.6151
R1062 B.n643 B.n642 10.6151
R1063 B.n645 B.n643 10.6151
R1064 B.n645 B.n644 10.6151
R1065 B.n644 B.n299 10.6151
R1066 B.n656 B.n299 10.6151
R1067 B.n657 B.n656 10.6151
R1068 B.n658 B.n657 10.6151
R1069 B.n659 B.n658 10.6151
R1070 B.n660 B.n659 10.6151
R1071 B.n664 B.n660 10.6151
R1072 B.n665 B.n664 10.6151
R1073 B.n666 B.n665 10.6151
R1074 B.n667 B.n666 10.6151
R1075 B.n669 B.n667 10.6151
R1076 B.n670 B.n669 10.6151
R1077 B.n671 B.n670 10.6151
R1078 B.n672 B.n671 10.6151
R1079 B.n674 B.n672 10.6151
R1080 B.n675 B.n674 10.6151
R1081 B.n676 B.n675 10.6151
R1082 B.n677 B.n676 10.6151
R1083 B.n679 B.n677 10.6151
R1084 B.n680 B.n679 10.6151
R1085 B.n681 B.n680 10.6151
R1086 B.n682 B.n681 10.6151
R1087 B.n683 B.n682 10.6151
R1088 B.n724 B.n1 10.6151
R1089 B.n724 B.n723 10.6151
R1090 B.n723 B.n722 10.6151
R1091 B.n722 B.n10 10.6151
R1092 B.n716 B.n10 10.6151
R1093 B.n716 B.n715 10.6151
R1094 B.n715 B.n714 10.6151
R1095 B.n714 B.n16 10.6151
R1096 B.n708 B.n16 10.6151
R1097 B.n708 B.n707 10.6151
R1098 B.n707 B.n706 10.6151
R1099 B.n706 B.n24 10.6151
R1100 B.n700 B.n24 10.6151
R1101 B.n700 B.n699 10.6151
R1102 B.n699 B.n698 10.6151
R1103 B.n698 B.n31 10.6151
R1104 B.n692 B.n31 10.6151
R1105 B.n692 B.n691 10.6151
R1106 B.n690 B.n38 10.6151
R1107 B.n97 B.n38 10.6151
R1108 B.n98 B.n97 10.6151
R1109 B.n101 B.n98 10.6151
R1110 B.n102 B.n101 10.6151
R1111 B.n105 B.n102 10.6151
R1112 B.n106 B.n105 10.6151
R1113 B.n109 B.n106 10.6151
R1114 B.n110 B.n109 10.6151
R1115 B.n113 B.n110 10.6151
R1116 B.n114 B.n113 10.6151
R1117 B.n117 B.n114 10.6151
R1118 B.n118 B.n117 10.6151
R1119 B.n121 B.n118 10.6151
R1120 B.n122 B.n121 10.6151
R1121 B.n125 B.n122 10.6151
R1122 B.n126 B.n125 10.6151
R1123 B.n129 B.n126 10.6151
R1124 B.n130 B.n129 10.6151
R1125 B.n133 B.n130 10.6151
R1126 B.n134 B.n133 10.6151
R1127 B.n137 B.n134 10.6151
R1128 B.n138 B.n137 10.6151
R1129 B.n141 B.n138 10.6151
R1130 B.n142 B.n141 10.6151
R1131 B.n145 B.n142 10.6151
R1132 B.n146 B.n145 10.6151
R1133 B.n149 B.n146 10.6151
R1134 B.n150 B.n149 10.6151
R1135 B.n153 B.n150 10.6151
R1136 B.n154 B.n153 10.6151
R1137 B.n157 B.n154 10.6151
R1138 B.n158 B.n157 10.6151
R1139 B.n161 B.n158 10.6151
R1140 B.n162 B.n161 10.6151
R1141 B.n165 B.n162 10.6151
R1142 B.n166 B.n165 10.6151
R1143 B.n169 B.n166 10.6151
R1144 B.n170 B.n169 10.6151
R1145 B.n173 B.n170 10.6151
R1146 B.n174 B.n173 10.6151
R1147 B.n177 B.n174 10.6151
R1148 B.n178 B.n177 10.6151
R1149 B.n181 B.n178 10.6151
R1150 B.n182 B.n181 10.6151
R1151 B.n185 B.n182 10.6151
R1152 B.n190 B.n187 10.6151
R1153 B.n191 B.n190 10.6151
R1154 B.n194 B.n191 10.6151
R1155 B.n195 B.n194 10.6151
R1156 B.n198 B.n195 10.6151
R1157 B.n199 B.n198 10.6151
R1158 B.n202 B.n199 10.6151
R1159 B.n203 B.n202 10.6151
R1160 B.n206 B.n203 10.6151
R1161 B.n211 B.n208 10.6151
R1162 B.n212 B.n211 10.6151
R1163 B.n215 B.n212 10.6151
R1164 B.n216 B.n215 10.6151
R1165 B.n219 B.n216 10.6151
R1166 B.n220 B.n219 10.6151
R1167 B.n223 B.n220 10.6151
R1168 B.n224 B.n223 10.6151
R1169 B.n227 B.n224 10.6151
R1170 B.n228 B.n227 10.6151
R1171 B.n231 B.n228 10.6151
R1172 B.n232 B.n231 10.6151
R1173 B.n235 B.n232 10.6151
R1174 B.n236 B.n235 10.6151
R1175 B.n239 B.n236 10.6151
R1176 B.n240 B.n239 10.6151
R1177 B.n243 B.n240 10.6151
R1178 B.n244 B.n243 10.6151
R1179 B.n247 B.n244 10.6151
R1180 B.n248 B.n247 10.6151
R1181 B.n251 B.n248 10.6151
R1182 B.n252 B.n251 10.6151
R1183 B.n255 B.n252 10.6151
R1184 B.n256 B.n255 10.6151
R1185 B.n259 B.n256 10.6151
R1186 B.n260 B.n259 10.6151
R1187 B.n263 B.n260 10.6151
R1188 B.n264 B.n263 10.6151
R1189 B.n267 B.n264 10.6151
R1190 B.n268 B.n267 10.6151
R1191 B.n271 B.n268 10.6151
R1192 B.n272 B.n271 10.6151
R1193 B.n275 B.n272 10.6151
R1194 B.n276 B.n275 10.6151
R1195 B.n279 B.n276 10.6151
R1196 B.n280 B.n279 10.6151
R1197 B.n283 B.n280 10.6151
R1198 B.n284 B.n283 10.6151
R1199 B.n287 B.n284 10.6151
R1200 B.n288 B.n287 10.6151
R1201 B.n291 B.n288 10.6151
R1202 B.n292 B.n291 10.6151
R1203 B.n295 B.n292 10.6151
R1204 B.n297 B.n295 10.6151
R1205 B.n298 B.n297 10.6151
R1206 B.n684 B.n298 10.6151
R1207 B.n508 B.n390 9.36635
R1208 B.n485 B.n393 9.36635
R1209 B.n186 B.n185 9.36635
R1210 B.n208 B.n207 9.36635
R1211 B.n732 B.n0 8.11757
R1212 B.n732 B.n1 8.11757
R1213 B.n633 B.t17 6.29112
R1214 B.n18 B.t1 6.29112
R1215 B.n615 B.t8 5.14737
R1216 B.t4 B.n702 5.14737
R1217 B.n505 B.n390 1.24928
R1218 B.n488 B.n393 1.24928
R1219 B.n187 B.n186 1.24928
R1220 B.n207 B.n206 1.24928
R1221 B.t2 B.n301 0.572374
R1222 B.n662 B.t0 0.572374
R1223 VN.n0 VN.t3 406.443
R1224 VN.n1 VN.t1 406.443
R1225 VN.n1 VN.t2 406.356
R1226 VN.n0 VN.t0 406.356
R1227 VN VN.n1 74.319
R1228 VN VN.n0 31.2622
R1229 VTAIL.n618 VTAIL.n546 289.615
R1230 VTAIL.n72 VTAIL.n0 289.615
R1231 VTAIL.n150 VTAIL.n78 289.615
R1232 VTAIL.n228 VTAIL.n156 289.615
R1233 VTAIL.n540 VTAIL.n468 289.615
R1234 VTAIL.n462 VTAIL.n390 289.615
R1235 VTAIL.n384 VTAIL.n312 289.615
R1236 VTAIL.n306 VTAIL.n234 289.615
R1237 VTAIL.n570 VTAIL.n569 185
R1238 VTAIL.n575 VTAIL.n574 185
R1239 VTAIL.n577 VTAIL.n576 185
R1240 VTAIL.n566 VTAIL.n565 185
R1241 VTAIL.n583 VTAIL.n582 185
R1242 VTAIL.n585 VTAIL.n584 185
R1243 VTAIL.n562 VTAIL.n561 185
R1244 VTAIL.n591 VTAIL.n590 185
R1245 VTAIL.n593 VTAIL.n592 185
R1246 VTAIL.n558 VTAIL.n557 185
R1247 VTAIL.n599 VTAIL.n598 185
R1248 VTAIL.n601 VTAIL.n600 185
R1249 VTAIL.n554 VTAIL.n553 185
R1250 VTAIL.n607 VTAIL.n606 185
R1251 VTAIL.n609 VTAIL.n608 185
R1252 VTAIL.n550 VTAIL.n549 185
R1253 VTAIL.n616 VTAIL.n615 185
R1254 VTAIL.n617 VTAIL.n548 185
R1255 VTAIL.n619 VTAIL.n618 185
R1256 VTAIL.n24 VTAIL.n23 185
R1257 VTAIL.n29 VTAIL.n28 185
R1258 VTAIL.n31 VTAIL.n30 185
R1259 VTAIL.n20 VTAIL.n19 185
R1260 VTAIL.n37 VTAIL.n36 185
R1261 VTAIL.n39 VTAIL.n38 185
R1262 VTAIL.n16 VTAIL.n15 185
R1263 VTAIL.n45 VTAIL.n44 185
R1264 VTAIL.n47 VTAIL.n46 185
R1265 VTAIL.n12 VTAIL.n11 185
R1266 VTAIL.n53 VTAIL.n52 185
R1267 VTAIL.n55 VTAIL.n54 185
R1268 VTAIL.n8 VTAIL.n7 185
R1269 VTAIL.n61 VTAIL.n60 185
R1270 VTAIL.n63 VTAIL.n62 185
R1271 VTAIL.n4 VTAIL.n3 185
R1272 VTAIL.n70 VTAIL.n69 185
R1273 VTAIL.n71 VTAIL.n2 185
R1274 VTAIL.n73 VTAIL.n72 185
R1275 VTAIL.n102 VTAIL.n101 185
R1276 VTAIL.n107 VTAIL.n106 185
R1277 VTAIL.n109 VTAIL.n108 185
R1278 VTAIL.n98 VTAIL.n97 185
R1279 VTAIL.n115 VTAIL.n114 185
R1280 VTAIL.n117 VTAIL.n116 185
R1281 VTAIL.n94 VTAIL.n93 185
R1282 VTAIL.n123 VTAIL.n122 185
R1283 VTAIL.n125 VTAIL.n124 185
R1284 VTAIL.n90 VTAIL.n89 185
R1285 VTAIL.n131 VTAIL.n130 185
R1286 VTAIL.n133 VTAIL.n132 185
R1287 VTAIL.n86 VTAIL.n85 185
R1288 VTAIL.n139 VTAIL.n138 185
R1289 VTAIL.n141 VTAIL.n140 185
R1290 VTAIL.n82 VTAIL.n81 185
R1291 VTAIL.n148 VTAIL.n147 185
R1292 VTAIL.n149 VTAIL.n80 185
R1293 VTAIL.n151 VTAIL.n150 185
R1294 VTAIL.n180 VTAIL.n179 185
R1295 VTAIL.n185 VTAIL.n184 185
R1296 VTAIL.n187 VTAIL.n186 185
R1297 VTAIL.n176 VTAIL.n175 185
R1298 VTAIL.n193 VTAIL.n192 185
R1299 VTAIL.n195 VTAIL.n194 185
R1300 VTAIL.n172 VTAIL.n171 185
R1301 VTAIL.n201 VTAIL.n200 185
R1302 VTAIL.n203 VTAIL.n202 185
R1303 VTAIL.n168 VTAIL.n167 185
R1304 VTAIL.n209 VTAIL.n208 185
R1305 VTAIL.n211 VTAIL.n210 185
R1306 VTAIL.n164 VTAIL.n163 185
R1307 VTAIL.n217 VTAIL.n216 185
R1308 VTAIL.n219 VTAIL.n218 185
R1309 VTAIL.n160 VTAIL.n159 185
R1310 VTAIL.n226 VTAIL.n225 185
R1311 VTAIL.n227 VTAIL.n158 185
R1312 VTAIL.n229 VTAIL.n228 185
R1313 VTAIL.n541 VTAIL.n540 185
R1314 VTAIL.n539 VTAIL.n470 185
R1315 VTAIL.n538 VTAIL.n537 185
R1316 VTAIL.n473 VTAIL.n471 185
R1317 VTAIL.n532 VTAIL.n531 185
R1318 VTAIL.n530 VTAIL.n529 185
R1319 VTAIL.n477 VTAIL.n476 185
R1320 VTAIL.n524 VTAIL.n523 185
R1321 VTAIL.n522 VTAIL.n521 185
R1322 VTAIL.n481 VTAIL.n480 185
R1323 VTAIL.n516 VTAIL.n515 185
R1324 VTAIL.n514 VTAIL.n513 185
R1325 VTAIL.n485 VTAIL.n484 185
R1326 VTAIL.n508 VTAIL.n507 185
R1327 VTAIL.n506 VTAIL.n505 185
R1328 VTAIL.n489 VTAIL.n488 185
R1329 VTAIL.n500 VTAIL.n499 185
R1330 VTAIL.n498 VTAIL.n497 185
R1331 VTAIL.n493 VTAIL.n492 185
R1332 VTAIL.n463 VTAIL.n462 185
R1333 VTAIL.n461 VTAIL.n392 185
R1334 VTAIL.n460 VTAIL.n459 185
R1335 VTAIL.n395 VTAIL.n393 185
R1336 VTAIL.n454 VTAIL.n453 185
R1337 VTAIL.n452 VTAIL.n451 185
R1338 VTAIL.n399 VTAIL.n398 185
R1339 VTAIL.n446 VTAIL.n445 185
R1340 VTAIL.n444 VTAIL.n443 185
R1341 VTAIL.n403 VTAIL.n402 185
R1342 VTAIL.n438 VTAIL.n437 185
R1343 VTAIL.n436 VTAIL.n435 185
R1344 VTAIL.n407 VTAIL.n406 185
R1345 VTAIL.n430 VTAIL.n429 185
R1346 VTAIL.n428 VTAIL.n427 185
R1347 VTAIL.n411 VTAIL.n410 185
R1348 VTAIL.n422 VTAIL.n421 185
R1349 VTAIL.n420 VTAIL.n419 185
R1350 VTAIL.n415 VTAIL.n414 185
R1351 VTAIL.n385 VTAIL.n384 185
R1352 VTAIL.n383 VTAIL.n314 185
R1353 VTAIL.n382 VTAIL.n381 185
R1354 VTAIL.n317 VTAIL.n315 185
R1355 VTAIL.n376 VTAIL.n375 185
R1356 VTAIL.n374 VTAIL.n373 185
R1357 VTAIL.n321 VTAIL.n320 185
R1358 VTAIL.n368 VTAIL.n367 185
R1359 VTAIL.n366 VTAIL.n365 185
R1360 VTAIL.n325 VTAIL.n324 185
R1361 VTAIL.n360 VTAIL.n359 185
R1362 VTAIL.n358 VTAIL.n357 185
R1363 VTAIL.n329 VTAIL.n328 185
R1364 VTAIL.n352 VTAIL.n351 185
R1365 VTAIL.n350 VTAIL.n349 185
R1366 VTAIL.n333 VTAIL.n332 185
R1367 VTAIL.n344 VTAIL.n343 185
R1368 VTAIL.n342 VTAIL.n341 185
R1369 VTAIL.n337 VTAIL.n336 185
R1370 VTAIL.n307 VTAIL.n306 185
R1371 VTAIL.n305 VTAIL.n236 185
R1372 VTAIL.n304 VTAIL.n303 185
R1373 VTAIL.n239 VTAIL.n237 185
R1374 VTAIL.n298 VTAIL.n297 185
R1375 VTAIL.n296 VTAIL.n295 185
R1376 VTAIL.n243 VTAIL.n242 185
R1377 VTAIL.n290 VTAIL.n289 185
R1378 VTAIL.n288 VTAIL.n287 185
R1379 VTAIL.n247 VTAIL.n246 185
R1380 VTAIL.n282 VTAIL.n281 185
R1381 VTAIL.n280 VTAIL.n279 185
R1382 VTAIL.n251 VTAIL.n250 185
R1383 VTAIL.n274 VTAIL.n273 185
R1384 VTAIL.n272 VTAIL.n271 185
R1385 VTAIL.n255 VTAIL.n254 185
R1386 VTAIL.n266 VTAIL.n265 185
R1387 VTAIL.n264 VTAIL.n263 185
R1388 VTAIL.n259 VTAIL.n258 185
R1389 VTAIL.n571 VTAIL.t2 147.659
R1390 VTAIL.n25 VTAIL.t1 147.659
R1391 VTAIL.n103 VTAIL.t6 147.659
R1392 VTAIL.n181 VTAIL.t7 147.659
R1393 VTAIL.n494 VTAIL.t5 147.659
R1394 VTAIL.n416 VTAIL.t4 147.659
R1395 VTAIL.n338 VTAIL.t3 147.659
R1396 VTAIL.n260 VTAIL.t0 147.659
R1397 VTAIL.n575 VTAIL.n569 104.615
R1398 VTAIL.n576 VTAIL.n575 104.615
R1399 VTAIL.n576 VTAIL.n565 104.615
R1400 VTAIL.n583 VTAIL.n565 104.615
R1401 VTAIL.n584 VTAIL.n583 104.615
R1402 VTAIL.n584 VTAIL.n561 104.615
R1403 VTAIL.n591 VTAIL.n561 104.615
R1404 VTAIL.n592 VTAIL.n591 104.615
R1405 VTAIL.n592 VTAIL.n557 104.615
R1406 VTAIL.n599 VTAIL.n557 104.615
R1407 VTAIL.n600 VTAIL.n599 104.615
R1408 VTAIL.n600 VTAIL.n553 104.615
R1409 VTAIL.n607 VTAIL.n553 104.615
R1410 VTAIL.n608 VTAIL.n607 104.615
R1411 VTAIL.n608 VTAIL.n549 104.615
R1412 VTAIL.n616 VTAIL.n549 104.615
R1413 VTAIL.n617 VTAIL.n616 104.615
R1414 VTAIL.n618 VTAIL.n617 104.615
R1415 VTAIL.n29 VTAIL.n23 104.615
R1416 VTAIL.n30 VTAIL.n29 104.615
R1417 VTAIL.n30 VTAIL.n19 104.615
R1418 VTAIL.n37 VTAIL.n19 104.615
R1419 VTAIL.n38 VTAIL.n37 104.615
R1420 VTAIL.n38 VTAIL.n15 104.615
R1421 VTAIL.n45 VTAIL.n15 104.615
R1422 VTAIL.n46 VTAIL.n45 104.615
R1423 VTAIL.n46 VTAIL.n11 104.615
R1424 VTAIL.n53 VTAIL.n11 104.615
R1425 VTAIL.n54 VTAIL.n53 104.615
R1426 VTAIL.n54 VTAIL.n7 104.615
R1427 VTAIL.n61 VTAIL.n7 104.615
R1428 VTAIL.n62 VTAIL.n61 104.615
R1429 VTAIL.n62 VTAIL.n3 104.615
R1430 VTAIL.n70 VTAIL.n3 104.615
R1431 VTAIL.n71 VTAIL.n70 104.615
R1432 VTAIL.n72 VTAIL.n71 104.615
R1433 VTAIL.n107 VTAIL.n101 104.615
R1434 VTAIL.n108 VTAIL.n107 104.615
R1435 VTAIL.n108 VTAIL.n97 104.615
R1436 VTAIL.n115 VTAIL.n97 104.615
R1437 VTAIL.n116 VTAIL.n115 104.615
R1438 VTAIL.n116 VTAIL.n93 104.615
R1439 VTAIL.n123 VTAIL.n93 104.615
R1440 VTAIL.n124 VTAIL.n123 104.615
R1441 VTAIL.n124 VTAIL.n89 104.615
R1442 VTAIL.n131 VTAIL.n89 104.615
R1443 VTAIL.n132 VTAIL.n131 104.615
R1444 VTAIL.n132 VTAIL.n85 104.615
R1445 VTAIL.n139 VTAIL.n85 104.615
R1446 VTAIL.n140 VTAIL.n139 104.615
R1447 VTAIL.n140 VTAIL.n81 104.615
R1448 VTAIL.n148 VTAIL.n81 104.615
R1449 VTAIL.n149 VTAIL.n148 104.615
R1450 VTAIL.n150 VTAIL.n149 104.615
R1451 VTAIL.n185 VTAIL.n179 104.615
R1452 VTAIL.n186 VTAIL.n185 104.615
R1453 VTAIL.n186 VTAIL.n175 104.615
R1454 VTAIL.n193 VTAIL.n175 104.615
R1455 VTAIL.n194 VTAIL.n193 104.615
R1456 VTAIL.n194 VTAIL.n171 104.615
R1457 VTAIL.n201 VTAIL.n171 104.615
R1458 VTAIL.n202 VTAIL.n201 104.615
R1459 VTAIL.n202 VTAIL.n167 104.615
R1460 VTAIL.n209 VTAIL.n167 104.615
R1461 VTAIL.n210 VTAIL.n209 104.615
R1462 VTAIL.n210 VTAIL.n163 104.615
R1463 VTAIL.n217 VTAIL.n163 104.615
R1464 VTAIL.n218 VTAIL.n217 104.615
R1465 VTAIL.n218 VTAIL.n159 104.615
R1466 VTAIL.n226 VTAIL.n159 104.615
R1467 VTAIL.n227 VTAIL.n226 104.615
R1468 VTAIL.n228 VTAIL.n227 104.615
R1469 VTAIL.n540 VTAIL.n539 104.615
R1470 VTAIL.n539 VTAIL.n538 104.615
R1471 VTAIL.n538 VTAIL.n471 104.615
R1472 VTAIL.n531 VTAIL.n471 104.615
R1473 VTAIL.n531 VTAIL.n530 104.615
R1474 VTAIL.n530 VTAIL.n476 104.615
R1475 VTAIL.n523 VTAIL.n476 104.615
R1476 VTAIL.n523 VTAIL.n522 104.615
R1477 VTAIL.n522 VTAIL.n480 104.615
R1478 VTAIL.n515 VTAIL.n480 104.615
R1479 VTAIL.n515 VTAIL.n514 104.615
R1480 VTAIL.n514 VTAIL.n484 104.615
R1481 VTAIL.n507 VTAIL.n484 104.615
R1482 VTAIL.n507 VTAIL.n506 104.615
R1483 VTAIL.n506 VTAIL.n488 104.615
R1484 VTAIL.n499 VTAIL.n488 104.615
R1485 VTAIL.n499 VTAIL.n498 104.615
R1486 VTAIL.n498 VTAIL.n492 104.615
R1487 VTAIL.n462 VTAIL.n461 104.615
R1488 VTAIL.n461 VTAIL.n460 104.615
R1489 VTAIL.n460 VTAIL.n393 104.615
R1490 VTAIL.n453 VTAIL.n393 104.615
R1491 VTAIL.n453 VTAIL.n452 104.615
R1492 VTAIL.n452 VTAIL.n398 104.615
R1493 VTAIL.n445 VTAIL.n398 104.615
R1494 VTAIL.n445 VTAIL.n444 104.615
R1495 VTAIL.n444 VTAIL.n402 104.615
R1496 VTAIL.n437 VTAIL.n402 104.615
R1497 VTAIL.n437 VTAIL.n436 104.615
R1498 VTAIL.n436 VTAIL.n406 104.615
R1499 VTAIL.n429 VTAIL.n406 104.615
R1500 VTAIL.n429 VTAIL.n428 104.615
R1501 VTAIL.n428 VTAIL.n410 104.615
R1502 VTAIL.n421 VTAIL.n410 104.615
R1503 VTAIL.n421 VTAIL.n420 104.615
R1504 VTAIL.n420 VTAIL.n414 104.615
R1505 VTAIL.n384 VTAIL.n383 104.615
R1506 VTAIL.n383 VTAIL.n382 104.615
R1507 VTAIL.n382 VTAIL.n315 104.615
R1508 VTAIL.n375 VTAIL.n315 104.615
R1509 VTAIL.n375 VTAIL.n374 104.615
R1510 VTAIL.n374 VTAIL.n320 104.615
R1511 VTAIL.n367 VTAIL.n320 104.615
R1512 VTAIL.n367 VTAIL.n366 104.615
R1513 VTAIL.n366 VTAIL.n324 104.615
R1514 VTAIL.n359 VTAIL.n324 104.615
R1515 VTAIL.n359 VTAIL.n358 104.615
R1516 VTAIL.n358 VTAIL.n328 104.615
R1517 VTAIL.n351 VTAIL.n328 104.615
R1518 VTAIL.n351 VTAIL.n350 104.615
R1519 VTAIL.n350 VTAIL.n332 104.615
R1520 VTAIL.n343 VTAIL.n332 104.615
R1521 VTAIL.n343 VTAIL.n342 104.615
R1522 VTAIL.n342 VTAIL.n336 104.615
R1523 VTAIL.n306 VTAIL.n305 104.615
R1524 VTAIL.n305 VTAIL.n304 104.615
R1525 VTAIL.n304 VTAIL.n237 104.615
R1526 VTAIL.n297 VTAIL.n237 104.615
R1527 VTAIL.n297 VTAIL.n296 104.615
R1528 VTAIL.n296 VTAIL.n242 104.615
R1529 VTAIL.n289 VTAIL.n242 104.615
R1530 VTAIL.n289 VTAIL.n288 104.615
R1531 VTAIL.n288 VTAIL.n246 104.615
R1532 VTAIL.n281 VTAIL.n246 104.615
R1533 VTAIL.n281 VTAIL.n280 104.615
R1534 VTAIL.n280 VTAIL.n250 104.615
R1535 VTAIL.n273 VTAIL.n250 104.615
R1536 VTAIL.n273 VTAIL.n272 104.615
R1537 VTAIL.n272 VTAIL.n254 104.615
R1538 VTAIL.n265 VTAIL.n254 104.615
R1539 VTAIL.n265 VTAIL.n264 104.615
R1540 VTAIL.n264 VTAIL.n258 104.615
R1541 VTAIL.t2 VTAIL.n569 52.3082
R1542 VTAIL.t1 VTAIL.n23 52.3082
R1543 VTAIL.t6 VTAIL.n101 52.3082
R1544 VTAIL.t7 VTAIL.n179 52.3082
R1545 VTAIL.t5 VTAIL.n492 52.3082
R1546 VTAIL.t4 VTAIL.n414 52.3082
R1547 VTAIL.t3 VTAIL.n336 52.3082
R1548 VTAIL.t0 VTAIL.n258 52.3082
R1549 VTAIL.n623 VTAIL.n622 32.9611
R1550 VTAIL.n77 VTAIL.n76 32.9611
R1551 VTAIL.n155 VTAIL.n154 32.9611
R1552 VTAIL.n233 VTAIL.n232 32.9611
R1553 VTAIL.n545 VTAIL.n544 32.9611
R1554 VTAIL.n467 VTAIL.n466 32.9611
R1555 VTAIL.n389 VTAIL.n388 32.9611
R1556 VTAIL.n311 VTAIL.n310 32.9611
R1557 VTAIL.n623 VTAIL.n545 25.5221
R1558 VTAIL.n311 VTAIL.n233 25.5221
R1559 VTAIL.n571 VTAIL.n570 15.6677
R1560 VTAIL.n25 VTAIL.n24 15.6677
R1561 VTAIL.n103 VTAIL.n102 15.6677
R1562 VTAIL.n181 VTAIL.n180 15.6677
R1563 VTAIL.n494 VTAIL.n493 15.6677
R1564 VTAIL.n416 VTAIL.n415 15.6677
R1565 VTAIL.n338 VTAIL.n337 15.6677
R1566 VTAIL.n260 VTAIL.n259 15.6677
R1567 VTAIL.n619 VTAIL.n548 13.1884
R1568 VTAIL.n73 VTAIL.n2 13.1884
R1569 VTAIL.n151 VTAIL.n80 13.1884
R1570 VTAIL.n229 VTAIL.n158 13.1884
R1571 VTAIL.n541 VTAIL.n470 13.1884
R1572 VTAIL.n463 VTAIL.n392 13.1884
R1573 VTAIL.n385 VTAIL.n314 13.1884
R1574 VTAIL.n307 VTAIL.n236 13.1884
R1575 VTAIL.n574 VTAIL.n573 12.8005
R1576 VTAIL.n615 VTAIL.n614 12.8005
R1577 VTAIL.n620 VTAIL.n546 12.8005
R1578 VTAIL.n28 VTAIL.n27 12.8005
R1579 VTAIL.n69 VTAIL.n68 12.8005
R1580 VTAIL.n74 VTAIL.n0 12.8005
R1581 VTAIL.n106 VTAIL.n105 12.8005
R1582 VTAIL.n147 VTAIL.n146 12.8005
R1583 VTAIL.n152 VTAIL.n78 12.8005
R1584 VTAIL.n184 VTAIL.n183 12.8005
R1585 VTAIL.n225 VTAIL.n224 12.8005
R1586 VTAIL.n230 VTAIL.n156 12.8005
R1587 VTAIL.n542 VTAIL.n468 12.8005
R1588 VTAIL.n537 VTAIL.n472 12.8005
R1589 VTAIL.n497 VTAIL.n496 12.8005
R1590 VTAIL.n464 VTAIL.n390 12.8005
R1591 VTAIL.n459 VTAIL.n394 12.8005
R1592 VTAIL.n419 VTAIL.n418 12.8005
R1593 VTAIL.n386 VTAIL.n312 12.8005
R1594 VTAIL.n381 VTAIL.n316 12.8005
R1595 VTAIL.n341 VTAIL.n340 12.8005
R1596 VTAIL.n308 VTAIL.n234 12.8005
R1597 VTAIL.n303 VTAIL.n238 12.8005
R1598 VTAIL.n263 VTAIL.n262 12.8005
R1599 VTAIL.n577 VTAIL.n568 12.0247
R1600 VTAIL.n613 VTAIL.n550 12.0247
R1601 VTAIL.n31 VTAIL.n22 12.0247
R1602 VTAIL.n67 VTAIL.n4 12.0247
R1603 VTAIL.n109 VTAIL.n100 12.0247
R1604 VTAIL.n145 VTAIL.n82 12.0247
R1605 VTAIL.n187 VTAIL.n178 12.0247
R1606 VTAIL.n223 VTAIL.n160 12.0247
R1607 VTAIL.n536 VTAIL.n473 12.0247
R1608 VTAIL.n500 VTAIL.n491 12.0247
R1609 VTAIL.n458 VTAIL.n395 12.0247
R1610 VTAIL.n422 VTAIL.n413 12.0247
R1611 VTAIL.n380 VTAIL.n317 12.0247
R1612 VTAIL.n344 VTAIL.n335 12.0247
R1613 VTAIL.n302 VTAIL.n239 12.0247
R1614 VTAIL.n266 VTAIL.n257 12.0247
R1615 VTAIL.n578 VTAIL.n566 11.249
R1616 VTAIL.n610 VTAIL.n609 11.249
R1617 VTAIL.n32 VTAIL.n20 11.249
R1618 VTAIL.n64 VTAIL.n63 11.249
R1619 VTAIL.n110 VTAIL.n98 11.249
R1620 VTAIL.n142 VTAIL.n141 11.249
R1621 VTAIL.n188 VTAIL.n176 11.249
R1622 VTAIL.n220 VTAIL.n219 11.249
R1623 VTAIL.n533 VTAIL.n532 11.249
R1624 VTAIL.n501 VTAIL.n489 11.249
R1625 VTAIL.n455 VTAIL.n454 11.249
R1626 VTAIL.n423 VTAIL.n411 11.249
R1627 VTAIL.n377 VTAIL.n376 11.249
R1628 VTAIL.n345 VTAIL.n333 11.249
R1629 VTAIL.n299 VTAIL.n298 11.249
R1630 VTAIL.n267 VTAIL.n255 11.249
R1631 VTAIL.n582 VTAIL.n581 10.4732
R1632 VTAIL.n606 VTAIL.n552 10.4732
R1633 VTAIL.n36 VTAIL.n35 10.4732
R1634 VTAIL.n60 VTAIL.n6 10.4732
R1635 VTAIL.n114 VTAIL.n113 10.4732
R1636 VTAIL.n138 VTAIL.n84 10.4732
R1637 VTAIL.n192 VTAIL.n191 10.4732
R1638 VTAIL.n216 VTAIL.n162 10.4732
R1639 VTAIL.n529 VTAIL.n475 10.4732
R1640 VTAIL.n505 VTAIL.n504 10.4732
R1641 VTAIL.n451 VTAIL.n397 10.4732
R1642 VTAIL.n427 VTAIL.n426 10.4732
R1643 VTAIL.n373 VTAIL.n319 10.4732
R1644 VTAIL.n349 VTAIL.n348 10.4732
R1645 VTAIL.n295 VTAIL.n241 10.4732
R1646 VTAIL.n271 VTAIL.n270 10.4732
R1647 VTAIL.n585 VTAIL.n564 9.69747
R1648 VTAIL.n605 VTAIL.n554 9.69747
R1649 VTAIL.n39 VTAIL.n18 9.69747
R1650 VTAIL.n59 VTAIL.n8 9.69747
R1651 VTAIL.n117 VTAIL.n96 9.69747
R1652 VTAIL.n137 VTAIL.n86 9.69747
R1653 VTAIL.n195 VTAIL.n174 9.69747
R1654 VTAIL.n215 VTAIL.n164 9.69747
R1655 VTAIL.n528 VTAIL.n477 9.69747
R1656 VTAIL.n508 VTAIL.n487 9.69747
R1657 VTAIL.n450 VTAIL.n399 9.69747
R1658 VTAIL.n430 VTAIL.n409 9.69747
R1659 VTAIL.n372 VTAIL.n321 9.69747
R1660 VTAIL.n352 VTAIL.n331 9.69747
R1661 VTAIL.n294 VTAIL.n243 9.69747
R1662 VTAIL.n274 VTAIL.n253 9.69747
R1663 VTAIL.n622 VTAIL.n621 9.45567
R1664 VTAIL.n76 VTAIL.n75 9.45567
R1665 VTAIL.n154 VTAIL.n153 9.45567
R1666 VTAIL.n232 VTAIL.n231 9.45567
R1667 VTAIL.n544 VTAIL.n543 9.45567
R1668 VTAIL.n466 VTAIL.n465 9.45567
R1669 VTAIL.n388 VTAIL.n387 9.45567
R1670 VTAIL.n310 VTAIL.n309 9.45567
R1671 VTAIL.n621 VTAIL.n620 9.3005
R1672 VTAIL.n560 VTAIL.n559 9.3005
R1673 VTAIL.n589 VTAIL.n588 9.3005
R1674 VTAIL.n587 VTAIL.n586 9.3005
R1675 VTAIL.n564 VTAIL.n563 9.3005
R1676 VTAIL.n581 VTAIL.n580 9.3005
R1677 VTAIL.n579 VTAIL.n578 9.3005
R1678 VTAIL.n568 VTAIL.n567 9.3005
R1679 VTAIL.n573 VTAIL.n572 9.3005
R1680 VTAIL.n595 VTAIL.n594 9.3005
R1681 VTAIL.n597 VTAIL.n596 9.3005
R1682 VTAIL.n556 VTAIL.n555 9.3005
R1683 VTAIL.n603 VTAIL.n602 9.3005
R1684 VTAIL.n605 VTAIL.n604 9.3005
R1685 VTAIL.n552 VTAIL.n551 9.3005
R1686 VTAIL.n611 VTAIL.n610 9.3005
R1687 VTAIL.n613 VTAIL.n612 9.3005
R1688 VTAIL.n614 VTAIL.n547 9.3005
R1689 VTAIL.n75 VTAIL.n74 9.3005
R1690 VTAIL.n14 VTAIL.n13 9.3005
R1691 VTAIL.n43 VTAIL.n42 9.3005
R1692 VTAIL.n41 VTAIL.n40 9.3005
R1693 VTAIL.n18 VTAIL.n17 9.3005
R1694 VTAIL.n35 VTAIL.n34 9.3005
R1695 VTAIL.n33 VTAIL.n32 9.3005
R1696 VTAIL.n22 VTAIL.n21 9.3005
R1697 VTAIL.n27 VTAIL.n26 9.3005
R1698 VTAIL.n49 VTAIL.n48 9.3005
R1699 VTAIL.n51 VTAIL.n50 9.3005
R1700 VTAIL.n10 VTAIL.n9 9.3005
R1701 VTAIL.n57 VTAIL.n56 9.3005
R1702 VTAIL.n59 VTAIL.n58 9.3005
R1703 VTAIL.n6 VTAIL.n5 9.3005
R1704 VTAIL.n65 VTAIL.n64 9.3005
R1705 VTAIL.n67 VTAIL.n66 9.3005
R1706 VTAIL.n68 VTAIL.n1 9.3005
R1707 VTAIL.n153 VTAIL.n152 9.3005
R1708 VTAIL.n92 VTAIL.n91 9.3005
R1709 VTAIL.n121 VTAIL.n120 9.3005
R1710 VTAIL.n119 VTAIL.n118 9.3005
R1711 VTAIL.n96 VTAIL.n95 9.3005
R1712 VTAIL.n113 VTAIL.n112 9.3005
R1713 VTAIL.n111 VTAIL.n110 9.3005
R1714 VTAIL.n100 VTAIL.n99 9.3005
R1715 VTAIL.n105 VTAIL.n104 9.3005
R1716 VTAIL.n127 VTAIL.n126 9.3005
R1717 VTAIL.n129 VTAIL.n128 9.3005
R1718 VTAIL.n88 VTAIL.n87 9.3005
R1719 VTAIL.n135 VTAIL.n134 9.3005
R1720 VTAIL.n137 VTAIL.n136 9.3005
R1721 VTAIL.n84 VTAIL.n83 9.3005
R1722 VTAIL.n143 VTAIL.n142 9.3005
R1723 VTAIL.n145 VTAIL.n144 9.3005
R1724 VTAIL.n146 VTAIL.n79 9.3005
R1725 VTAIL.n231 VTAIL.n230 9.3005
R1726 VTAIL.n170 VTAIL.n169 9.3005
R1727 VTAIL.n199 VTAIL.n198 9.3005
R1728 VTAIL.n197 VTAIL.n196 9.3005
R1729 VTAIL.n174 VTAIL.n173 9.3005
R1730 VTAIL.n191 VTAIL.n190 9.3005
R1731 VTAIL.n189 VTAIL.n188 9.3005
R1732 VTAIL.n178 VTAIL.n177 9.3005
R1733 VTAIL.n183 VTAIL.n182 9.3005
R1734 VTAIL.n205 VTAIL.n204 9.3005
R1735 VTAIL.n207 VTAIL.n206 9.3005
R1736 VTAIL.n166 VTAIL.n165 9.3005
R1737 VTAIL.n213 VTAIL.n212 9.3005
R1738 VTAIL.n215 VTAIL.n214 9.3005
R1739 VTAIL.n162 VTAIL.n161 9.3005
R1740 VTAIL.n221 VTAIL.n220 9.3005
R1741 VTAIL.n223 VTAIL.n222 9.3005
R1742 VTAIL.n224 VTAIL.n157 9.3005
R1743 VTAIL.n520 VTAIL.n519 9.3005
R1744 VTAIL.n479 VTAIL.n478 9.3005
R1745 VTAIL.n526 VTAIL.n525 9.3005
R1746 VTAIL.n528 VTAIL.n527 9.3005
R1747 VTAIL.n475 VTAIL.n474 9.3005
R1748 VTAIL.n534 VTAIL.n533 9.3005
R1749 VTAIL.n536 VTAIL.n535 9.3005
R1750 VTAIL.n472 VTAIL.n469 9.3005
R1751 VTAIL.n543 VTAIL.n542 9.3005
R1752 VTAIL.n518 VTAIL.n517 9.3005
R1753 VTAIL.n483 VTAIL.n482 9.3005
R1754 VTAIL.n512 VTAIL.n511 9.3005
R1755 VTAIL.n510 VTAIL.n509 9.3005
R1756 VTAIL.n487 VTAIL.n486 9.3005
R1757 VTAIL.n504 VTAIL.n503 9.3005
R1758 VTAIL.n502 VTAIL.n501 9.3005
R1759 VTAIL.n491 VTAIL.n490 9.3005
R1760 VTAIL.n496 VTAIL.n495 9.3005
R1761 VTAIL.n442 VTAIL.n441 9.3005
R1762 VTAIL.n401 VTAIL.n400 9.3005
R1763 VTAIL.n448 VTAIL.n447 9.3005
R1764 VTAIL.n450 VTAIL.n449 9.3005
R1765 VTAIL.n397 VTAIL.n396 9.3005
R1766 VTAIL.n456 VTAIL.n455 9.3005
R1767 VTAIL.n458 VTAIL.n457 9.3005
R1768 VTAIL.n394 VTAIL.n391 9.3005
R1769 VTAIL.n465 VTAIL.n464 9.3005
R1770 VTAIL.n440 VTAIL.n439 9.3005
R1771 VTAIL.n405 VTAIL.n404 9.3005
R1772 VTAIL.n434 VTAIL.n433 9.3005
R1773 VTAIL.n432 VTAIL.n431 9.3005
R1774 VTAIL.n409 VTAIL.n408 9.3005
R1775 VTAIL.n426 VTAIL.n425 9.3005
R1776 VTAIL.n424 VTAIL.n423 9.3005
R1777 VTAIL.n413 VTAIL.n412 9.3005
R1778 VTAIL.n418 VTAIL.n417 9.3005
R1779 VTAIL.n364 VTAIL.n363 9.3005
R1780 VTAIL.n323 VTAIL.n322 9.3005
R1781 VTAIL.n370 VTAIL.n369 9.3005
R1782 VTAIL.n372 VTAIL.n371 9.3005
R1783 VTAIL.n319 VTAIL.n318 9.3005
R1784 VTAIL.n378 VTAIL.n377 9.3005
R1785 VTAIL.n380 VTAIL.n379 9.3005
R1786 VTAIL.n316 VTAIL.n313 9.3005
R1787 VTAIL.n387 VTAIL.n386 9.3005
R1788 VTAIL.n362 VTAIL.n361 9.3005
R1789 VTAIL.n327 VTAIL.n326 9.3005
R1790 VTAIL.n356 VTAIL.n355 9.3005
R1791 VTAIL.n354 VTAIL.n353 9.3005
R1792 VTAIL.n331 VTAIL.n330 9.3005
R1793 VTAIL.n348 VTAIL.n347 9.3005
R1794 VTAIL.n346 VTAIL.n345 9.3005
R1795 VTAIL.n335 VTAIL.n334 9.3005
R1796 VTAIL.n340 VTAIL.n339 9.3005
R1797 VTAIL.n286 VTAIL.n285 9.3005
R1798 VTAIL.n245 VTAIL.n244 9.3005
R1799 VTAIL.n292 VTAIL.n291 9.3005
R1800 VTAIL.n294 VTAIL.n293 9.3005
R1801 VTAIL.n241 VTAIL.n240 9.3005
R1802 VTAIL.n300 VTAIL.n299 9.3005
R1803 VTAIL.n302 VTAIL.n301 9.3005
R1804 VTAIL.n238 VTAIL.n235 9.3005
R1805 VTAIL.n309 VTAIL.n308 9.3005
R1806 VTAIL.n284 VTAIL.n283 9.3005
R1807 VTAIL.n249 VTAIL.n248 9.3005
R1808 VTAIL.n278 VTAIL.n277 9.3005
R1809 VTAIL.n276 VTAIL.n275 9.3005
R1810 VTAIL.n253 VTAIL.n252 9.3005
R1811 VTAIL.n270 VTAIL.n269 9.3005
R1812 VTAIL.n268 VTAIL.n267 9.3005
R1813 VTAIL.n257 VTAIL.n256 9.3005
R1814 VTAIL.n262 VTAIL.n261 9.3005
R1815 VTAIL.n586 VTAIL.n562 8.92171
R1816 VTAIL.n602 VTAIL.n601 8.92171
R1817 VTAIL.n40 VTAIL.n16 8.92171
R1818 VTAIL.n56 VTAIL.n55 8.92171
R1819 VTAIL.n118 VTAIL.n94 8.92171
R1820 VTAIL.n134 VTAIL.n133 8.92171
R1821 VTAIL.n196 VTAIL.n172 8.92171
R1822 VTAIL.n212 VTAIL.n211 8.92171
R1823 VTAIL.n525 VTAIL.n524 8.92171
R1824 VTAIL.n509 VTAIL.n485 8.92171
R1825 VTAIL.n447 VTAIL.n446 8.92171
R1826 VTAIL.n431 VTAIL.n407 8.92171
R1827 VTAIL.n369 VTAIL.n368 8.92171
R1828 VTAIL.n353 VTAIL.n329 8.92171
R1829 VTAIL.n291 VTAIL.n290 8.92171
R1830 VTAIL.n275 VTAIL.n251 8.92171
R1831 VTAIL.n590 VTAIL.n589 8.14595
R1832 VTAIL.n598 VTAIL.n556 8.14595
R1833 VTAIL.n44 VTAIL.n43 8.14595
R1834 VTAIL.n52 VTAIL.n10 8.14595
R1835 VTAIL.n122 VTAIL.n121 8.14595
R1836 VTAIL.n130 VTAIL.n88 8.14595
R1837 VTAIL.n200 VTAIL.n199 8.14595
R1838 VTAIL.n208 VTAIL.n166 8.14595
R1839 VTAIL.n521 VTAIL.n479 8.14595
R1840 VTAIL.n513 VTAIL.n512 8.14595
R1841 VTAIL.n443 VTAIL.n401 8.14595
R1842 VTAIL.n435 VTAIL.n434 8.14595
R1843 VTAIL.n365 VTAIL.n323 8.14595
R1844 VTAIL.n357 VTAIL.n356 8.14595
R1845 VTAIL.n287 VTAIL.n245 8.14595
R1846 VTAIL.n279 VTAIL.n278 8.14595
R1847 VTAIL.n593 VTAIL.n560 7.3702
R1848 VTAIL.n597 VTAIL.n558 7.3702
R1849 VTAIL.n47 VTAIL.n14 7.3702
R1850 VTAIL.n51 VTAIL.n12 7.3702
R1851 VTAIL.n125 VTAIL.n92 7.3702
R1852 VTAIL.n129 VTAIL.n90 7.3702
R1853 VTAIL.n203 VTAIL.n170 7.3702
R1854 VTAIL.n207 VTAIL.n168 7.3702
R1855 VTAIL.n520 VTAIL.n481 7.3702
R1856 VTAIL.n516 VTAIL.n483 7.3702
R1857 VTAIL.n442 VTAIL.n403 7.3702
R1858 VTAIL.n438 VTAIL.n405 7.3702
R1859 VTAIL.n364 VTAIL.n325 7.3702
R1860 VTAIL.n360 VTAIL.n327 7.3702
R1861 VTAIL.n286 VTAIL.n247 7.3702
R1862 VTAIL.n282 VTAIL.n249 7.3702
R1863 VTAIL.n594 VTAIL.n593 6.59444
R1864 VTAIL.n594 VTAIL.n558 6.59444
R1865 VTAIL.n48 VTAIL.n47 6.59444
R1866 VTAIL.n48 VTAIL.n12 6.59444
R1867 VTAIL.n126 VTAIL.n125 6.59444
R1868 VTAIL.n126 VTAIL.n90 6.59444
R1869 VTAIL.n204 VTAIL.n203 6.59444
R1870 VTAIL.n204 VTAIL.n168 6.59444
R1871 VTAIL.n517 VTAIL.n481 6.59444
R1872 VTAIL.n517 VTAIL.n516 6.59444
R1873 VTAIL.n439 VTAIL.n403 6.59444
R1874 VTAIL.n439 VTAIL.n438 6.59444
R1875 VTAIL.n361 VTAIL.n325 6.59444
R1876 VTAIL.n361 VTAIL.n360 6.59444
R1877 VTAIL.n283 VTAIL.n247 6.59444
R1878 VTAIL.n283 VTAIL.n282 6.59444
R1879 VTAIL.n590 VTAIL.n560 5.81868
R1880 VTAIL.n598 VTAIL.n597 5.81868
R1881 VTAIL.n44 VTAIL.n14 5.81868
R1882 VTAIL.n52 VTAIL.n51 5.81868
R1883 VTAIL.n122 VTAIL.n92 5.81868
R1884 VTAIL.n130 VTAIL.n129 5.81868
R1885 VTAIL.n200 VTAIL.n170 5.81868
R1886 VTAIL.n208 VTAIL.n207 5.81868
R1887 VTAIL.n521 VTAIL.n520 5.81868
R1888 VTAIL.n513 VTAIL.n483 5.81868
R1889 VTAIL.n443 VTAIL.n442 5.81868
R1890 VTAIL.n435 VTAIL.n405 5.81868
R1891 VTAIL.n365 VTAIL.n364 5.81868
R1892 VTAIL.n357 VTAIL.n327 5.81868
R1893 VTAIL.n287 VTAIL.n286 5.81868
R1894 VTAIL.n279 VTAIL.n249 5.81868
R1895 VTAIL.n589 VTAIL.n562 5.04292
R1896 VTAIL.n601 VTAIL.n556 5.04292
R1897 VTAIL.n43 VTAIL.n16 5.04292
R1898 VTAIL.n55 VTAIL.n10 5.04292
R1899 VTAIL.n121 VTAIL.n94 5.04292
R1900 VTAIL.n133 VTAIL.n88 5.04292
R1901 VTAIL.n199 VTAIL.n172 5.04292
R1902 VTAIL.n211 VTAIL.n166 5.04292
R1903 VTAIL.n524 VTAIL.n479 5.04292
R1904 VTAIL.n512 VTAIL.n485 5.04292
R1905 VTAIL.n446 VTAIL.n401 5.04292
R1906 VTAIL.n434 VTAIL.n407 5.04292
R1907 VTAIL.n368 VTAIL.n323 5.04292
R1908 VTAIL.n356 VTAIL.n329 5.04292
R1909 VTAIL.n290 VTAIL.n245 5.04292
R1910 VTAIL.n278 VTAIL.n251 5.04292
R1911 VTAIL.n572 VTAIL.n571 4.38563
R1912 VTAIL.n26 VTAIL.n25 4.38563
R1913 VTAIL.n104 VTAIL.n103 4.38563
R1914 VTAIL.n182 VTAIL.n181 4.38563
R1915 VTAIL.n495 VTAIL.n494 4.38563
R1916 VTAIL.n417 VTAIL.n416 4.38563
R1917 VTAIL.n339 VTAIL.n338 4.38563
R1918 VTAIL.n261 VTAIL.n260 4.38563
R1919 VTAIL.n586 VTAIL.n585 4.26717
R1920 VTAIL.n602 VTAIL.n554 4.26717
R1921 VTAIL.n40 VTAIL.n39 4.26717
R1922 VTAIL.n56 VTAIL.n8 4.26717
R1923 VTAIL.n118 VTAIL.n117 4.26717
R1924 VTAIL.n134 VTAIL.n86 4.26717
R1925 VTAIL.n196 VTAIL.n195 4.26717
R1926 VTAIL.n212 VTAIL.n164 4.26717
R1927 VTAIL.n525 VTAIL.n477 4.26717
R1928 VTAIL.n509 VTAIL.n508 4.26717
R1929 VTAIL.n447 VTAIL.n399 4.26717
R1930 VTAIL.n431 VTAIL.n430 4.26717
R1931 VTAIL.n369 VTAIL.n321 4.26717
R1932 VTAIL.n353 VTAIL.n352 4.26717
R1933 VTAIL.n291 VTAIL.n243 4.26717
R1934 VTAIL.n275 VTAIL.n274 4.26717
R1935 VTAIL.n582 VTAIL.n564 3.49141
R1936 VTAIL.n606 VTAIL.n605 3.49141
R1937 VTAIL.n36 VTAIL.n18 3.49141
R1938 VTAIL.n60 VTAIL.n59 3.49141
R1939 VTAIL.n114 VTAIL.n96 3.49141
R1940 VTAIL.n138 VTAIL.n137 3.49141
R1941 VTAIL.n192 VTAIL.n174 3.49141
R1942 VTAIL.n216 VTAIL.n215 3.49141
R1943 VTAIL.n529 VTAIL.n528 3.49141
R1944 VTAIL.n505 VTAIL.n487 3.49141
R1945 VTAIL.n451 VTAIL.n450 3.49141
R1946 VTAIL.n427 VTAIL.n409 3.49141
R1947 VTAIL.n373 VTAIL.n372 3.49141
R1948 VTAIL.n349 VTAIL.n331 3.49141
R1949 VTAIL.n295 VTAIL.n294 3.49141
R1950 VTAIL.n271 VTAIL.n253 3.49141
R1951 VTAIL.n581 VTAIL.n566 2.71565
R1952 VTAIL.n609 VTAIL.n552 2.71565
R1953 VTAIL.n35 VTAIL.n20 2.71565
R1954 VTAIL.n63 VTAIL.n6 2.71565
R1955 VTAIL.n113 VTAIL.n98 2.71565
R1956 VTAIL.n141 VTAIL.n84 2.71565
R1957 VTAIL.n191 VTAIL.n176 2.71565
R1958 VTAIL.n219 VTAIL.n162 2.71565
R1959 VTAIL.n532 VTAIL.n475 2.71565
R1960 VTAIL.n504 VTAIL.n489 2.71565
R1961 VTAIL.n454 VTAIL.n397 2.71565
R1962 VTAIL.n426 VTAIL.n411 2.71565
R1963 VTAIL.n376 VTAIL.n319 2.71565
R1964 VTAIL.n348 VTAIL.n333 2.71565
R1965 VTAIL.n298 VTAIL.n241 2.71565
R1966 VTAIL.n270 VTAIL.n255 2.71565
R1967 VTAIL.n578 VTAIL.n577 1.93989
R1968 VTAIL.n610 VTAIL.n550 1.93989
R1969 VTAIL.n32 VTAIL.n31 1.93989
R1970 VTAIL.n64 VTAIL.n4 1.93989
R1971 VTAIL.n110 VTAIL.n109 1.93989
R1972 VTAIL.n142 VTAIL.n82 1.93989
R1973 VTAIL.n188 VTAIL.n187 1.93989
R1974 VTAIL.n220 VTAIL.n160 1.93989
R1975 VTAIL.n533 VTAIL.n473 1.93989
R1976 VTAIL.n501 VTAIL.n500 1.93989
R1977 VTAIL.n455 VTAIL.n395 1.93989
R1978 VTAIL.n423 VTAIL.n422 1.93989
R1979 VTAIL.n377 VTAIL.n317 1.93989
R1980 VTAIL.n345 VTAIL.n344 1.93989
R1981 VTAIL.n299 VTAIL.n239 1.93989
R1982 VTAIL.n267 VTAIL.n266 1.93989
R1983 VTAIL.n574 VTAIL.n568 1.16414
R1984 VTAIL.n615 VTAIL.n613 1.16414
R1985 VTAIL.n622 VTAIL.n546 1.16414
R1986 VTAIL.n28 VTAIL.n22 1.16414
R1987 VTAIL.n69 VTAIL.n67 1.16414
R1988 VTAIL.n76 VTAIL.n0 1.16414
R1989 VTAIL.n106 VTAIL.n100 1.16414
R1990 VTAIL.n147 VTAIL.n145 1.16414
R1991 VTAIL.n154 VTAIL.n78 1.16414
R1992 VTAIL.n184 VTAIL.n178 1.16414
R1993 VTAIL.n225 VTAIL.n223 1.16414
R1994 VTAIL.n232 VTAIL.n156 1.16414
R1995 VTAIL.n544 VTAIL.n468 1.16414
R1996 VTAIL.n537 VTAIL.n536 1.16414
R1997 VTAIL.n497 VTAIL.n491 1.16414
R1998 VTAIL.n466 VTAIL.n390 1.16414
R1999 VTAIL.n459 VTAIL.n458 1.16414
R2000 VTAIL.n419 VTAIL.n413 1.16414
R2001 VTAIL.n388 VTAIL.n312 1.16414
R2002 VTAIL.n381 VTAIL.n380 1.16414
R2003 VTAIL.n341 VTAIL.n335 1.16414
R2004 VTAIL.n310 VTAIL.n234 1.16414
R2005 VTAIL.n303 VTAIL.n302 1.16414
R2006 VTAIL.n263 VTAIL.n257 1.16414
R2007 VTAIL.n389 VTAIL.n311 1.12119
R2008 VTAIL.n545 VTAIL.n467 1.12119
R2009 VTAIL.n233 VTAIL.n155 1.12119
R2010 VTAIL VTAIL.n77 0.619035
R2011 VTAIL VTAIL.n623 0.502655
R2012 VTAIL.n467 VTAIL.n389 0.470328
R2013 VTAIL.n155 VTAIL.n77 0.470328
R2014 VTAIL.n573 VTAIL.n570 0.388379
R2015 VTAIL.n614 VTAIL.n548 0.388379
R2016 VTAIL.n620 VTAIL.n619 0.388379
R2017 VTAIL.n27 VTAIL.n24 0.388379
R2018 VTAIL.n68 VTAIL.n2 0.388379
R2019 VTAIL.n74 VTAIL.n73 0.388379
R2020 VTAIL.n105 VTAIL.n102 0.388379
R2021 VTAIL.n146 VTAIL.n80 0.388379
R2022 VTAIL.n152 VTAIL.n151 0.388379
R2023 VTAIL.n183 VTAIL.n180 0.388379
R2024 VTAIL.n224 VTAIL.n158 0.388379
R2025 VTAIL.n230 VTAIL.n229 0.388379
R2026 VTAIL.n542 VTAIL.n541 0.388379
R2027 VTAIL.n472 VTAIL.n470 0.388379
R2028 VTAIL.n496 VTAIL.n493 0.388379
R2029 VTAIL.n464 VTAIL.n463 0.388379
R2030 VTAIL.n394 VTAIL.n392 0.388379
R2031 VTAIL.n418 VTAIL.n415 0.388379
R2032 VTAIL.n386 VTAIL.n385 0.388379
R2033 VTAIL.n316 VTAIL.n314 0.388379
R2034 VTAIL.n340 VTAIL.n337 0.388379
R2035 VTAIL.n308 VTAIL.n307 0.388379
R2036 VTAIL.n238 VTAIL.n236 0.388379
R2037 VTAIL.n262 VTAIL.n259 0.388379
R2038 VTAIL.n572 VTAIL.n567 0.155672
R2039 VTAIL.n579 VTAIL.n567 0.155672
R2040 VTAIL.n580 VTAIL.n579 0.155672
R2041 VTAIL.n580 VTAIL.n563 0.155672
R2042 VTAIL.n587 VTAIL.n563 0.155672
R2043 VTAIL.n588 VTAIL.n587 0.155672
R2044 VTAIL.n588 VTAIL.n559 0.155672
R2045 VTAIL.n595 VTAIL.n559 0.155672
R2046 VTAIL.n596 VTAIL.n595 0.155672
R2047 VTAIL.n596 VTAIL.n555 0.155672
R2048 VTAIL.n603 VTAIL.n555 0.155672
R2049 VTAIL.n604 VTAIL.n603 0.155672
R2050 VTAIL.n604 VTAIL.n551 0.155672
R2051 VTAIL.n611 VTAIL.n551 0.155672
R2052 VTAIL.n612 VTAIL.n611 0.155672
R2053 VTAIL.n612 VTAIL.n547 0.155672
R2054 VTAIL.n621 VTAIL.n547 0.155672
R2055 VTAIL.n26 VTAIL.n21 0.155672
R2056 VTAIL.n33 VTAIL.n21 0.155672
R2057 VTAIL.n34 VTAIL.n33 0.155672
R2058 VTAIL.n34 VTAIL.n17 0.155672
R2059 VTAIL.n41 VTAIL.n17 0.155672
R2060 VTAIL.n42 VTAIL.n41 0.155672
R2061 VTAIL.n42 VTAIL.n13 0.155672
R2062 VTAIL.n49 VTAIL.n13 0.155672
R2063 VTAIL.n50 VTAIL.n49 0.155672
R2064 VTAIL.n50 VTAIL.n9 0.155672
R2065 VTAIL.n57 VTAIL.n9 0.155672
R2066 VTAIL.n58 VTAIL.n57 0.155672
R2067 VTAIL.n58 VTAIL.n5 0.155672
R2068 VTAIL.n65 VTAIL.n5 0.155672
R2069 VTAIL.n66 VTAIL.n65 0.155672
R2070 VTAIL.n66 VTAIL.n1 0.155672
R2071 VTAIL.n75 VTAIL.n1 0.155672
R2072 VTAIL.n104 VTAIL.n99 0.155672
R2073 VTAIL.n111 VTAIL.n99 0.155672
R2074 VTAIL.n112 VTAIL.n111 0.155672
R2075 VTAIL.n112 VTAIL.n95 0.155672
R2076 VTAIL.n119 VTAIL.n95 0.155672
R2077 VTAIL.n120 VTAIL.n119 0.155672
R2078 VTAIL.n120 VTAIL.n91 0.155672
R2079 VTAIL.n127 VTAIL.n91 0.155672
R2080 VTAIL.n128 VTAIL.n127 0.155672
R2081 VTAIL.n128 VTAIL.n87 0.155672
R2082 VTAIL.n135 VTAIL.n87 0.155672
R2083 VTAIL.n136 VTAIL.n135 0.155672
R2084 VTAIL.n136 VTAIL.n83 0.155672
R2085 VTAIL.n143 VTAIL.n83 0.155672
R2086 VTAIL.n144 VTAIL.n143 0.155672
R2087 VTAIL.n144 VTAIL.n79 0.155672
R2088 VTAIL.n153 VTAIL.n79 0.155672
R2089 VTAIL.n182 VTAIL.n177 0.155672
R2090 VTAIL.n189 VTAIL.n177 0.155672
R2091 VTAIL.n190 VTAIL.n189 0.155672
R2092 VTAIL.n190 VTAIL.n173 0.155672
R2093 VTAIL.n197 VTAIL.n173 0.155672
R2094 VTAIL.n198 VTAIL.n197 0.155672
R2095 VTAIL.n198 VTAIL.n169 0.155672
R2096 VTAIL.n205 VTAIL.n169 0.155672
R2097 VTAIL.n206 VTAIL.n205 0.155672
R2098 VTAIL.n206 VTAIL.n165 0.155672
R2099 VTAIL.n213 VTAIL.n165 0.155672
R2100 VTAIL.n214 VTAIL.n213 0.155672
R2101 VTAIL.n214 VTAIL.n161 0.155672
R2102 VTAIL.n221 VTAIL.n161 0.155672
R2103 VTAIL.n222 VTAIL.n221 0.155672
R2104 VTAIL.n222 VTAIL.n157 0.155672
R2105 VTAIL.n231 VTAIL.n157 0.155672
R2106 VTAIL.n543 VTAIL.n469 0.155672
R2107 VTAIL.n535 VTAIL.n469 0.155672
R2108 VTAIL.n535 VTAIL.n534 0.155672
R2109 VTAIL.n534 VTAIL.n474 0.155672
R2110 VTAIL.n527 VTAIL.n474 0.155672
R2111 VTAIL.n527 VTAIL.n526 0.155672
R2112 VTAIL.n526 VTAIL.n478 0.155672
R2113 VTAIL.n519 VTAIL.n478 0.155672
R2114 VTAIL.n519 VTAIL.n518 0.155672
R2115 VTAIL.n518 VTAIL.n482 0.155672
R2116 VTAIL.n511 VTAIL.n482 0.155672
R2117 VTAIL.n511 VTAIL.n510 0.155672
R2118 VTAIL.n510 VTAIL.n486 0.155672
R2119 VTAIL.n503 VTAIL.n486 0.155672
R2120 VTAIL.n503 VTAIL.n502 0.155672
R2121 VTAIL.n502 VTAIL.n490 0.155672
R2122 VTAIL.n495 VTAIL.n490 0.155672
R2123 VTAIL.n465 VTAIL.n391 0.155672
R2124 VTAIL.n457 VTAIL.n391 0.155672
R2125 VTAIL.n457 VTAIL.n456 0.155672
R2126 VTAIL.n456 VTAIL.n396 0.155672
R2127 VTAIL.n449 VTAIL.n396 0.155672
R2128 VTAIL.n449 VTAIL.n448 0.155672
R2129 VTAIL.n448 VTAIL.n400 0.155672
R2130 VTAIL.n441 VTAIL.n400 0.155672
R2131 VTAIL.n441 VTAIL.n440 0.155672
R2132 VTAIL.n440 VTAIL.n404 0.155672
R2133 VTAIL.n433 VTAIL.n404 0.155672
R2134 VTAIL.n433 VTAIL.n432 0.155672
R2135 VTAIL.n432 VTAIL.n408 0.155672
R2136 VTAIL.n425 VTAIL.n408 0.155672
R2137 VTAIL.n425 VTAIL.n424 0.155672
R2138 VTAIL.n424 VTAIL.n412 0.155672
R2139 VTAIL.n417 VTAIL.n412 0.155672
R2140 VTAIL.n387 VTAIL.n313 0.155672
R2141 VTAIL.n379 VTAIL.n313 0.155672
R2142 VTAIL.n379 VTAIL.n378 0.155672
R2143 VTAIL.n378 VTAIL.n318 0.155672
R2144 VTAIL.n371 VTAIL.n318 0.155672
R2145 VTAIL.n371 VTAIL.n370 0.155672
R2146 VTAIL.n370 VTAIL.n322 0.155672
R2147 VTAIL.n363 VTAIL.n322 0.155672
R2148 VTAIL.n363 VTAIL.n362 0.155672
R2149 VTAIL.n362 VTAIL.n326 0.155672
R2150 VTAIL.n355 VTAIL.n326 0.155672
R2151 VTAIL.n355 VTAIL.n354 0.155672
R2152 VTAIL.n354 VTAIL.n330 0.155672
R2153 VTAIL.n347 VTAIL.n330 0.155672
R2154 VTAIL.n347 VTAIL.n346 0.155672
R2155 VTAIL.n346 VTAIL.n334 0.155672
R2156 VTAIL.n339 VTAIL.n334 0.155672
R2157 VTAIL.n309 VTAIL.n235 0.155672
R2158 VTAIL.n301 VTAIL.n235 0.155672
R2159 VTAIL.n301 VTAIL.n300 0.155672
R2160 VTAIL.n300 VTAIL.n240 0.155672
R2161 VTAIL.n293 VTAIL.n240 0.155672
R2162 VTAIL.n293 VTAIL.n292 0.155672
R2163 VTAIL.n292 VTAIL.n244 0.155672
R2164 VTAIL.n285 VTAIL.n244 0.155672
R2165 VTAIL.n285 VTAIL.n284 0.155672
R2166 VTAIL.n284 VTAIL.n248 0.155672
R2167 VTAIL.n277 VTAIL.n248 0.155672
R2168 VTAIL.n277 VTAIL.n276 0.155672
R2169 VTAIL.n276 VTAIL.n252 0.155672
R2170 VTAIL.n269 VTAIL.n252 0.155672
R2171 VTAIL.n269 VTAIL.n268 0.155672
R2172 VTAIL.n268 VTAIL.n256 0.155672
R2173 VTAIL.n261 VTAIL.n256 0.155672
R2174 VDD2.n2 VDD2.n0 100.901
R2175 VDD2.n2 VDD2.n1 61.79
R2176 VDD2.n1 VDD2.t1 1.41884
R2177 VDD2.n1 VDD2.t2 1.41884
R2178 VDD2.n0 VDD2.t0 1.41884
R2179 VDD2.n0 VDD2.t3 1.41884
R2180 VDD2 VDD2.n2 0.0586897
R2181 VP.n0 VP.t3 406.443
R2182 VP.n0 VP.t2 406.356
R2183 VP.n2 VP.t0 387.837
R2184 VP.n3 VP.t1 387.837
R2185 VP.n4 VP.n3 80.6037
R2186 VP.n2 VP.n1 80.6037
R2187 VP.n1 VP.n0 74.0335
R2188 VP.n3 VP.n2 48.2005
R2189 VP.n4 VP.n1 0.380177
R2190 VP VP.n4 0.146778
R2191 VDD1 VDD1.n1 101.427
R2192 VDD1 VDD1.n0 61.8482
R2193 VDD1.n0 VDD1.t0 1.41884
R2194 VDD1.n0 VDD1.t1 1.41884
R2195 VDD1.n1 VDD1.t3 1.41884
R2196 VDD1.n1 VDD1.t2 1.41884
C0 VP VDD2 0.290363f
C1 VN VDD1 0.147304f
C2 VN VTAIL 3.74113f
C3 VTAIL VDD1 6.8372f
C4 VN VDD2 4.15879f
C5 VDD1 VDD2 0.63147f
C6 VTAIL VDD2 6.88048f
C7 VN VP 5.38371f
C8 VDD1 VP 4.30152f
C9 VTAIL VP 3.75524f
C10 VDD2 B 3.009942f
C11 VDD1 B 6.89342f
C12 VTAIL B 10.13306f
C13 VN B 8.571671f
C14 VP B 5.621939f
C15 VDD1.t0 B 0.300042f
C16 VDD1.t1 B 0.300042f
C17 VDD1.n0 B 2.70403f
C18 VDD1.t3 B 0.300042f
C19 VDD1.t2 B 0.300042f
C20 VDD1.n1 B 3.3954f
C21 VP.t2 B 1.72901f
C22 VP.t3 B 1.72917f
C23 VP.n0 B 2.42801f
C24 VP.n1 B 2.79862f
C25 VP.t0 B 1.69889f
C26 VP.n2 B 0.660954f
C27 VP.t1 B 1.69889f
C28 VP.n3 B 0.660954f
C29 VP.n4 B 0.056027f
C30 VDD2.t0 B 0.302782f
C31 VDD2.t3 B 0.302782f
C32 VDD2.n0 B 3.39933f
C33 VDD2.t1 B 0.302782f
C34 VDD2.t2 B 0.302782f
C35 VDD2.n1 B 2.72841f
C36 VDD2.n2 B 3.65611f
C37 VTAIL.n0 B 0.019972f
C38 VTAIL.n1 B 0.015718f
C39 VTAIL.n2 B 0.008695f
C40 VTAIL.n3 B 0.019964f
C41 VTAIL.n4 B 0.008943f
C42 VTAIL.n5 B 0.015718f
C43 VTAIL.n6 B 0.008446f
C44 VTAIL.n7 B 0.019964f
C45 VTAIL.n8 B 0.008943f
C46 VTAIL.n9 B 0.015718f
C47 VTAIL.n10 B 0.008446f
C48 VTAIL.n11 B 0.019964f
C49 VTAIL.n12 B 0.008943f
C50 VTAIL.n13 B 0.015718f
C51 VTAIL.n14 B 0.008446f
C52 VTAIL.n15 B 0.019964f
C53 VTAIL.n16 B 0.008943f
C54 VTAIL.n17 B 0.015718f
C55 VTAIL.n18 B 0.008446f
C56 VTAIL.n19 B 0.019964f
C57 VTAIL.n20 B 0.008943f
C58 VTAIL.n21 B 0.015718f
C59 VTAIL.n22 B 0.008446f
C60 VTAIL.n23 B 0.014973f
C61 VTAIL.n24 B 0.011793f
C62 VTAIL.t1 B 0.032862f
C63 VTAIL.n25 B 0.098419f
C64 VTAIL.n26 B 0.947735f
C65 VTAIL.n27 B 0.008446f
C66 VTAIL.n28 B 0.008943f
C67 VTAIL.n29 B 0.019964f
C68 VTAIL.n30 B 0.019964f
C69 VTAIL.n31 B 0.008943f
C70 VTAIL.n32 B 0.008446f
C71 VTAIL.n33 B 0.015718f
C72 VTAIL.n34 B 0.015718f
C73 VTAIL.n35 B 0.008446f
C74 VTAIL.n36 B 0.008943f
C75 VTAIL.n37 B 0.019964f
C76 VTAIL.n38 B 0.019964f
C77 VTAIL.n39 B 0.008943f
C78 VTAIL.n40 B 0.008446f
C79 VTAIL.n41 B 0.015718f
C80 VTAIL.n42 B 0.015718f
C81 VTAIL.n43 B 0.008446f
C82 VTAIL.n44 B 0.008943f
C83 VTAIL.n45 B 0.019964f
C84 VTAIL.n46 B 0.019964f
C85 VTAIL.n47 B 0.008943f
C86 VTAIL.n48 B 0.008446f
C87 VTAIL.n49 B 0.015718f
C88 VTAIL.n50 B 0.015718f
C89 VTAIL.n51 B 0.008446f
C90 VTAIL.n52 B 0.008943f
C91 VTAIL.n53 B 0.019964f
C92 VTAIL.n54 B 0.019964f
C93 VTAIL.n55 B 0.008943f
C94 VTAIL.n56 B 0.008446f
C95 VTAIL.n57 B 0.015718f
C96 VTAIL.n58 B 0.015718f
C97 VTAIL.n59 B 0.008446f
C98 VTAIL.n60 B 0.008943f
C99 VTAIL.n61 B 0.019964f
C100 VTAIL.n62 B 0.019964f
C101 VTAIL.n63 B 0.008943f
C102 VTAIL.n64 B 0.008446f
C103 VTAIL.n65 B 0.015718f
C104 VTAIL.n66 B 0.015718f
C105 VTAIL.n67 B 0.008446f
C106 VTAIL.n68 B 0.008446f
C107 VTAIL.n69 B 0.008943f
C108 VTAIL.n70 B 0.019964f
C109 VTAIL.n71 B 0.019964f
C110 VTAIL.n72 B 0.039468f
C111 VTAIL.n73 B 0.008695f
C112 VTAIL.n74 B 0.008446f
C113 VTAIL.n75 B 0.037191f
C114 VTAIL.n76 B 0.021725f
C115 VTAIL.n77 B 0.069033f
C116 VTAIL.n78 B 0.019972f
C117 VTAIL.n79 B 0.015718f
C118 VTAIL.n80 B 0.008695f
C119 VTAIL.n81 B 0.019964f
C120 VTAIL.n82 B 0.008943f
C121 VTAIL.n83 B 0.015718f
C122 VTAIL.n84 B 0.008446f
C123 VTAIL.n85 B 0.019964f
C124 VTAIL.n86 B 0.008943f
C125 VTAIL.n87 B 0.015718f
C126 VTAIL.n88 B 0.008446f
C127 VTAIL.n89 B 0.019964f
C128 VTAIL.n90 B 0.008943f
C129 VTAIL.n91 B 0.015718f
C130 VTAIL.n92 B 0.008446f
C131 VTAIL.n93 B 0.019964f
C132 VTAIL.n94 B 0.008943f
C133 VTAIL.n95 B 0.015718f
C134 VTAIL.n96 B 0.008446f
C135 VTAIL.n97 B 0.019964f
C136 VTAIL.n98 B 0.008943f
C137 VTAIL.n99 B 0.015718f
C138 VTAIL.n100 B 0.008446f
C139 VTAIL.n101 B 0.014973f
C140 VTAIL.n102 B 0.011793f
C141 VTAIL.t6 B 0.032862f
C142 VTAIL.n103 B 0.098419f
C143 VTAIL.n104 B 0.947735f
C144 VTAIL.n105 B 0.008446f
C145 VTAIL.n106 B 0.008943f
C146 VTAIL.n107 B 0.019964f
C147 VTAIL.n108 B 0.019964f
C148 VTAIL.n109 B 0.008943f
C149 VTAIL.n110 B 0.008446f
C150 VTAIL.n111 B 0.015718f
C151 VTAIL.n112 B 0.015718f
C152 VTAIL.n113 B 0.008446f
C153 VTAIL.n114 B 0.008943f
C154 VTAIL.n115 B 0.019964f
C155 VTAIL.n116 B 0.019964f
C156 VTAIL.n117 B 0.008943f
C157 VTAIL.n118 B 0.008446f
C158 VTAIL.n119 B 0.015718f
C159 VTAIL.n120 B 0.015718f
C160 VTAIL.n121 B 0.008446f
C161 VTAIL.n122 B 0.008943f
C162 VTAIL.n123 B 0.019964f
C163 VTAIL.n124 B 0.019964f
C164 VTAIL.n125 B 0.008943f
C165 VTAIL.n126 B 0.008446f
C166 VTAIL.n127 B 0.015718f
C167 VTAIL.n128 B 0.015718f
C168 VTAIL.n129 B 0.008446f
C169 VTAIL.n130 B 0.008943f
C170 VTAIL.n131 B 0.019964f
C171 VTAIL.n132 B 0.019964f
C172 VTAIL.n133 B 0.008943f
C173 VTAIL.n134 B 0.008446f
C174 VTAIL.n135 B 0.015718f
C175 VTAIL.n136 B 0.015718f
C176 VTAIL.n137 B 0.008446f
C177 VTAIL.n138 B 0.008943f
C178 VTAIL.n139 B 0.019964f
C179 VTAIL.n140 B 0.019964f
C180 VTAIL.n141 B 0.008943f
C181 VTAIL.n142 B 0.008446f
C182 VTAIL.n143 B 0.015718f
C183 VTAIL.n144 B 0.015718f
C184 VTAIL.n145 B 0.008446f
C185 VTAIL.n146 B 0.008446f
C186 VTAIL.n147 B 0.008943f
C187 VTAIL.n148 B 0.019964f
C188 VTAIL.n149 B 0.019964f
C189 VTAIL.n150 B 0.039468f
C190 VTAIL.n151 B 0.008695f
C191 VTAIL.n152 B 0.008446f
C192 VTAIL.n153 B 0.037191f
C193 VTAIL.n154 B 0.021725f
C194 VTAIL.n155 B 0.094466f
C195 VTAIL.n156 B 0.019972f
C196 VTAIL.n157 B 0.015718f
C197 VTAIL.n158 B 0.008695f
C198 VTAIL.n159 B 0.019964f
C199 VTAIL.n160 B 0.008943f
C200 VTAIL.n161 B 0.015718f
C201 VTAIL.n162 B 0.008446f
C202 VTAIL.n163 B 0.019964f
C203 VTAIL.n164 B 0.008943f
C204 VTAIL.n165 B 0.015718f
C205 VTAIL.n166 B 0.008446f
C206 VTAIL.n167 B 0.019964f
C207 VTAIL.n168 B 0.008943f
C208 VTAIL.n169 B 0.015718f
C209 VTAIL.n170 B 0.008446f
C210 VTAIL.n171 B 0.019964f
C211 VTAIL.n172 B 0.008943f
C212 VTAIL.n173 B 0.015718f
C213 VTAIL.n174 B 0.008446f
C214 VTAIL.n175 B 0.019964f
C215 VTAIL.n176 B 0.008943f
C216 VTAIL.n177 B 0.015718f
C217 VTAIL.n178 B 0.008446f
C218 VTAIL.n179 B 0.014973f
C219 VTAIL.n180 B 0.011793f
C220 VTAIL.t7 B 0.032862f
C221 VTAIL.n181 B 0.098419f
C222 VTAIL.n182 B 0.947735f
C223 VTAIL.n183 B 0.008446f
C224 VTAIL.n184 B 0.008943f
C225 VTAIL.n185 B 0.019964f
C226 VTAIL.n186 B 0.019964f
C227 VTAIL.n187 B 0.008943f
C228 VTAIL.n188 B 0.008446f
C229 VTAIL.n189 B 0.015718f
C230 VTAIL.n190 B 0.015718f
C231 VTAIL.n191 B 0.008446f
C232 VTAIL.n192 B 0.008943f
C233 VTAIL.n193 B 0.019964f
C234 VTAIL.n194 B 0.019964f
C235 VTAIL.n195 B 0.008943f
C236 VTAIL.n196 B 0.008446f
C237 VTAIL.n197 B 0.015718f
C238 VTAIL.n198 B 0.015718f
C239 VTAIL.n199 B 0.008446f
C240 VTAIL.n200 B 0.008943f
C241 VTAIL.n201 B 0.019964f
C242 VTAIL.n202 B 0.019964f
C243 VTAIL.n203 B 0.008943f
C244 VTAIL.n204 B 0.008446f
C245 VTAIL.n205 B 0.015718f
C246 VTAIL.n206 B 0.015718f
C247 VTAIL.n207 B 0.008446f
C248 VTAIL.n208 B 0.008943f
C249 VTAIL.n209 B 0.019964f
C250 VTAIL.n210 B 0.019964f
C251 VTAIL.n211 B 0.008943f
C252 VTAIL.n212 B 0.008446f
C253 VTAIL.n213 B 0.015718f
C254 VTAIL.n214 B 0.015718f
C255 VTAIL.n215 B 0.008446f
C256 VTAIL.n216 B 0.008943f
C257 VTAIL.n217 B 0.019964f
C258 VTAIL.n218 B 0.019964f
C259 VTAIL.n219 B 0.008943f
C260 VTAIL.n220 B 0.008446f
C261 VTAIL.n221 B 0.015718f
C262 VTAIL.n222 B 0.015718f
C263 VTAIL.n223 B 0.008446f
C264 VTAIL.n224 B 0.008446f
C265 VTAIL.n225 B 0.008943f
C266 VTAIL.n226 B 0.019964f
C267 VTAIL.n227 B 0.019964f
C268 VTAIL.n228 B 0.039468f
C269 VTAIL.n229 B 0.008695f
C270 VTAIL.n230 B 0.008446f
C271 VTAIL.n231 B 0.037191f
C272 VTAIL.n232 B 0.021725f
C273 VTAIL.n233 B 0.950465f
C274 VTAIL.n234 B 0.019972f
C275 VTAIL.n235 B 0.015718f
C276 VTAIL.n236 B 0.008695f
C277 VTAIL.n237 B 0.019964f
C278 VTAIL.n238 B 0.008446f
C279 VTAIL.n239 B 0.008943f
C280 VTAIL.n240 B 0.015718f
C281 VTAIL.n241 B 0.008446f
C282 VTAIL.n242 B 0.019964f
C283 VTAIL.n243 B 0.008943f
C284 VTAIL.n244 B 0.015718f
C285 VTAIL.n245 B 0.008446f
C286 VTAIL.n246 B 0.019964f
C287 VTAIL.n247 B 0.008943f
C288 VTAIL.n248 B 0.015718f
C289 VTAIL.n249 B 0.008446f
C290 VTAIL.n250 B 0.019964f
C291 VTAIL.n251 B 0.008943f
C292 VTAIL.n252 B 0.015718f
C293 VTAIL.n253 B 0.008446f
C294 VTAIL.n254 B 0.019964f
C295 VTAIL.n255 B 0.008943f
C296 VTAIL.n256 B 0.015718f
C297 VTAIL.n257 B 0.008446f
C298 VTAIL.n258 B 0.014973f
C299 VTAIL.n259 B 0.011793f
C300 VTAIL.t0 B 0.032862f
C301 VTAIL.n260 B 0.098419f
C302 VTAIL.n261 B 0.947735f
C303 VTAIL.n262 B 0.008446f
C304 VTAIL.n263 B 0.008943f
C305 VTAIL.n264 B 0.019964f
C306 VTAIL.n265 B 0.019964f
C307 VTAIL.n266 B 0.008943f
C308 VTAIL.n267 B 0.008446f
C309 VTAIL.n268 B 0.015718f
C310 VTAIL.n269 B 0.015718f
C311 VTAIL.n270 B 0.008446f
C312 VTAIL.n271 B 0.008943f
C313 VTAIL.n272 B 0.019964f
C314 VTAIL.n273 B 0.019964f
C315 VTAIL.n274 B 0.008943f
C316 VTAIL.n275 B 0.008446f
C317 VTAIL.n276 B 0.015718f
C318 VTAIL.n277 B 0.015718f
C319 VTAIL.n278 B 0.008446f
C320 VTAIL.n279 B 0.008943f
C321 VTAIL.n280 B 0.019964f
C322 VTAIL.n281 B 0.019964f
C323 VTAIL.n282 B 0.008943f
C324 VTAIL.n283 B 0.008446f
C325 VTAIL.n284 B 0.015718f
C326 VTAIL.n285 B 0.015718f
C327 VTAIL.n286 B 0.008446f
C328 VTAIL.n287 B 0.008943f
C329 VTAIL.n288 B 0.019964f
C330 VTAIL.n289 B 0.019964f
C331 VTAIL.n290 B 0.008943f
C332 VTAIL.n291 B 0.008446f
C333 VTAIL.n292 B 0.015718f
C334 VTAIL.n293 B 0.015718f
C335 VTAIL.n294 B 0.008446f
C336 VTAIL.n295 B 0.008943f
C337 VTAIL.n296 B 0.019964f
C338 VTAIL.n297 B 0.019964f
C339 VTAIL.n298 B 0.008943f
C340 VTAIL.n299 B 0.008446f
C341 VTAIL.n300 B 0.015718f
C342 VTAIL.n301 B 0.015718f
C343 VTAIL.n302 B 0.008446f
C344 VTAIL.n303 B 0.008943f
C345 VTAIL.n304 B 0.019964f
C346 VTAIL.n305 B 0.019964f
C347 VTAIL.n306 B 0.039468f
C348 VTAIL.n307 B 0.008695f
C349 VTAIL.n308 B 0.008446f
C350 VTAIL.n309 B 0.037191f
C351 VTAIL.n310 B 0.021725f
C352 VTAIL.n311 B 0.950465f
C353 VTAIL.n312 B 0.019972f
C354 VTAIL.n313 B 0.015718f
C355 VTAIL.n314 B 0.008695f
C356 VTAIL.n315 B 0.019964f
C357 VTAIL.n316 B 0.008446f
C358 VTAIL.n317 B 0.008943f
C359 VTAIL.n318 B 0.015718f
C360 VTAIL.n319 B 0.008446f
C361 VTAIL.n320 B 0.019964f
C362 VTAIL.n321 B 0.008943f
C363 VTAIL.n322 B 0.015718f
C364 VTAIL.n323 B 0.008446f
C365 VTAIL.n324 B 0.019964f
C366 VTAIL.n325 B 0.008943f
C367 VTAIL.n326 B 0.015718f
C368 VTAIL.n327 B 0.008446f
C369 VTAIL.n328 B 0.019964f
C370 VTAIL.n329 B 0.008943f
C371 VTAIL.n330 B 0.015718f
C372 VTAIL.n331 B 0.008446f
C373 VTAIL.n332 B 0.019964f
C374 VTAIL.n333 B 0.008943f
C375 VTAIL.n334 B 0.015718f
C376 VTAIL.n335 B 0.008446f
C377 VTAIL.n336 B 0.014973f
C378 VTAIL.n337 B 0.011793f
C379 VTAIL.t3 B 0.032862f
C380 VTAIL.n338 B 0.098419f
C381 VTAIL.n339 B 0.947735f
C382 VTAIL.n340 B 0.008446f
C383 VTAIL.n341 B 0.008943f
C384 VTAIL.n342 B 0.019964f
C385 VTAIL.n343 B 0.019964f
C386 VTAIL.n344 B 0.008943f
C387 VTAIL.n345 B 0.008446f
C388 VTAIL.n346 B 0.015718f
C389 VTAIL.n347 B 0.015718f
C390 VTAIL.n348 B 0.008446f
C391 VTAIL.n349 B 0.008943f
C392 VTAIL.n350 B 0.019964f
C393 VTAIL.n351 B 0.019964f
C394 VTAIL.n352 B 0.008943f
C395 VTAIL.n353 B 0.008446f
C396 VTAIL.n354 B 0.015718f
C397 VTAIL.n355 B 0.015718f
C398 VTAIL.n356 B 0.008446f
C399 VTAIL.n357 B 0.008943f
C400 VTAIL.n358 B 0.019964f
C401 VTAIL.n359 B 0.019964f
C402 VTAIL.n360 B 0.008943f
C403 VTAIL.n361 B 0.008446f
C404 VTAIL.n362 B 0.015718f
C405 VTAIL.n363 B 0.015718f
C406 VTAIL.n364 B 0.008446f
C407 VTAIL.n365 B 0.008943f
C408 VTAIL.n366 B 0.019964f
C409 VTAIL.n367 B 0.019964f
C410 VTAIL.n368 B 0.008943f
C411 VTAIL.n369 B 0.008446f
C412 VTAIL.n370 B 0.015718f
C413 VTAIL.n371 B 0.015718f
C414 VTAIL.n372 B 0.008446f
C415 VTAIL.n373 B 0.008943f
C416 VTAIL.n374 B 0.019964f
C417 VTAIL.n375 B 0.019964f
C418 VTAIL.n376 B 0.008943f
C419 VTAIL.n377 B 0.008446f
C420 VTAIL.n378 B 0.015718f
C421 VTAIL.n379 B 0.015718f
C422 VTAIL.n380 B 0.008446f
C423 VTAIL.n381 B 0.008943f
C424 VTAIL.n382 B 0.019964f
C425 VTAIL.n383 B 0.019964f
C426 VTAIL.n384 B 0.039468f
C427 VTAIL.n385 B 0.008695f
C428 VTAIL.n386 B 0.008446f
C429 VTAIL.n387 B 0.037191f
C430 VTAIL.n388 B 0.021725f
C431 VTAIL.n389 B 0.094466f
C432 VTAIL.n390 B 0.019972f
C433 VTAIL.n391 B 0.015718f
C434 VTAIL.n392 B 0.008695f
C435 VTAIL.n393 B 0.019964f
C436 VTAIL.n394 B 0.008446f
C437 VTAIL.n395 B 0.008943f
C438 VTAIL.n396 B 0.015718f
C439 VTAIL.n397 B 0.008446f
C440 VTAIL.n398 B 0.019964f
C441 VTAIL.n399 B 0.008943f
C442 VTAIL.n400 B 0.015718f
C443 VTAIL.n401 B 0.008446f
C444 VTAIL.n402 B 0.019964f
C445 VTAIL.n403 B 0.008943f
C446 VTAIL.n404 B 0.015718f
C447 VTAIL.n405 B 0.008446f
C448 VTAIL.n406 B 0.019964f
C449 VTAIL.n407 B 0.008943f
C450 VTAIL.n408 B 0.015718f
C451 VTAIL.n409 B 0.008446f
C452 VTAIL.n410 B 0.019964f
C453 VTAIL.n411 B 0.008943f
C454 VTAIL.n412 B 0.015718f
C455 VTAIL.n413 B 0.008446f
C456 VTAIL.n414 B 0.014973f
C457 VTAIL.n415 B 0.011793f
C458 VTAIL.t4 B 0.032862f
C459 VTAIL.n416 B 0.098419f
C460 VTAIL.n417 B 0.947735f
C461 VTAIL.n418 B 0.008446f
C462 VTAIL.n419 B 0.008943f
C463 VTAIL.n420 B 0.019964f
C464 VTAIL.n421 B 0.019964f
C465 VTAIL.n422 B 0.008943f
C466 VTAIL.n423 B 0.008446f
C467 VTAIL.n424 B 0.015718f
C468 VTAIL.n425 B 0.015718f
C469 VTAIL.n426 B 0.008446f
C470 VTAIL.n427 B 0.008943f
C471 VTAIL.n428 B 0.019964f
C472 VTAIL.n429 B 0.019964f
C473 VTAIL.n430 B 0.008943f
C474 VTAIL.n431 B 0.008446f
C475 VTAIL.n432 B 0.015718f
C476 VTAIL.n433 B 0.015718f
C477 VTAIL.n434 B 0.008446f
C478 VTAIL.n435 B 0.008943f
C479 VTAIL.n436 B 0.019964f
C480 VTAIL.n437 B 0.019964f
C481 VTAIL.n438 B 0.008943f
C482 VTAIL.n439 B 0.008446f
C483 VTAIL.n440 B 0.015718f
C484 VTAIL.n441 B 0.015718f
C485 VTAIL.n442 B 0.008446f
C486 VTAIL.n443 B 0.008943f
C487 VTAIL.n444 B 0.019964f
C488 VTAIL.n445 B 0.019964f
C489 VTAIL.n446 B 0.008943f
C490 VTAIL.n447 B 0.008446f
C491 VTAIL.n448 B 0.015718f
C492 VTAIL.n449 B 0.015718f
C493 VTAIL.n450 B 0.008446f
C494 VTAIL.n451 B 0.008943f
C495 VTAIL.n452 B 0.019964f
C496 VTAIL.n453 B 0.019964f
C497 VTAIL.n454 B 0.008943f
C498 VTAIL.n455 B 0.008446f
C499 VTAIL.n456 B 0.015718f
C500 VTAIL.n457 B 0.015718f
C501 VTAIL.n458 B 0.008446f
C502 VTAIL.n459 B 0.008943f
C503 VTAIL.n460 B 0.019964f
C504 VTAIL.n461 B 0.019964f
C505 VTAIL.n462 B 0.039468f
C506 VTAIL.n463 B 0.008695f
C507 VTAIL.n464 B 0.008446f
C508 VTAIL.n465 B 0.037191f
C509 VTAIL.n466 B 0.021725f
C510 VTAIL.n467 B 0.094466f
C511 VTAIL.n468 B 0.019972f
C512 VTAIL.n469 B 0.015718f
C513 VTAIL.n470 B 0.008695f
C514 VTAIL.n471 B 0.019964f
C515 VTAIL.n472 B 0.008446f
C516 VTAIL.n473 B 0.008943f
C517 VTAIL.n474 B 0.015718f
C518 VTAIL.n475 B 0.008446f
C519 VTAIL.n476 B 0.019964f
C520 VTAIL.n477 B 0.008943f
C521 VTAIL.n478 B 0.015718f
C522 VTAIL.n479 B 0.008446f
C523 VTAIL.n480 B 0.019964f
C524 VTAIL.n481 B 0.008943f
C525 VTAIL.n482 B 0.015718f
C526 VTAIL.n483 B 0.008446f
C527 VTAIL.n484 B 0.019964f
C528 VTAIL.n485 B 0.008943f
C529 VTAIL.n486 B 0.015718f
C530 VTAIL.n487 B 0.008446f
C531 VTAIL.n488 B 0.019964f
C532 VTAIL.n489 B 0.008943f
C533 VTAIL.n490 B 0.015718f
C534 VTAIL.n491 B 0.008446f
C535 VTAIL.n492 B 0.014973f
C536 VTAIL.n493 B 0.011793f
C537 VTAIL.t5 B 0.032862f
C538 VTAIL.n494 B 0.098419f
C539 VTAIL.n495 B 0.947735f
C540 VTAIL.n496 B 0.008446f
C541 VTAIL.n497 B 0.008943f
C542 VTAIL.n498 B 0.019964f
C543 VTAIL.n499 B 0.019964f
C544 VTAIL.n500 B 0.008943f
C545 VTAIL.n501 B 0.008446f
C546 VTAIL.n502 B 0.015718f
C547 VTAIL.n503 B 0.015718f
C548 VTAIL.n504 B 0.008446f
C549 VTAIL.n505 B 0.008943f
C550 VTAIL.n506 B 0.019964f
C551 VTAIL.n507 B 0.019964f
C552 VTAIL.n508 B 0.008943f
C553 VTAIL.n509 B 0.008446f
C554 VTAIL.n510 B 0.015718f
C555 VTAIL.n511 B 0.015718f
C556 VTAIL.n512 B 0.008446f
C557 VTAIL.n513 B 0.008943f
C558 VTAIL.n514 B 0.019964f
C559 VTAIL.n515 B 0.019964f
C560 VTAIL.n516 B 0.008943f
C561 VTAIL.n517 B 0.008446f
C562 VTAIL.n518 B 0.015718f
C563 VTAIL.n519 B 0.015718f
C564 VTAIL.n520 B 0.008446f
C565 VTAIL.n521 B 0.008943f
C566 VTAIL.n522 B 0.019964f
C567 VTAIL.n523 B 0.019964f
C568 VTAIL.n524 B 0.008943f
C569 VTAIL.n525 B 0.008446f
C570 VTAIL.n526 B 0.015718f
C571 VTAIL.n527 B 0.015718f
C572 VTAIL.n528 B 0.008446f
C573 VTAIL.n529 B 0.008943f
C574 VTAIL.n530 B 0.019964f
C575 VTAIL.n531 B 0.019964f
C576 VTAIL.n532 B 0.008943f
C577 VTAIL.n533 B 0.008446f
C578 VTAIL.n534 B 0.015718f
C579 VTAIL.n535 B 0.015718f
C580 VTAIL.n536 B 0.008446f
C581 VTAIL.n537 B 0.008943f
C582 VTAIL.n538 B 0.019964f
C583 VTAIL.n539 B 0.019964f
C584 VTAIL.n540 B 0.039468f
C585 VTAIL.n541 B 0.008695f
C586 VTAIL.n542 B 0.008446f
C587 VTAIL.n543 B 0.037191f
C588 VTAIL.n544 B 0.021725f
C589 VTAIL.n545 B 0.950465f
C590 VTAIL.n546 B 0.019972f
C591 VTAIL.n547 B 0.015718f
C592 VTAIL.n548 B 0.008695f
C593 VTAIL.n549 B 0.019964f
C594 VTAIL.n550 B 0.008943f
C595 VTAIL.n551 B 0.015718f
C596 VTAIL.n552 B 0.008446f
C597 VTAIL.n553 B 0.019964f
C598 VTAIL.n554 B 0.008943f
C599 VTAIL.n555 B 0.015718f
C600 VTAIL.n556 B 0.008446f
C601 VTAIL.n557 B 0.019964f
C602 VTAIL.n558 B 0.008943f
C603 VTAIL.n559 B 0.015718f
C604 VTAIL.n560 B 0.008446f
C605 VTAIL.n561 B 0.019964f
C606 VTAIL.n562 B 0.008943f
C607 VTAIL.n563 B 0.015718f
C608 VTAIL.n564 B 0.008446f
C609 VTAIL.n565 B 0.019964f
C610 VTAIL.n566 B 0.008943f
C611 VTAIL.n567 B 0.015718f
C612 VTAIL.n568 B 0.008446f
C613 VTAIL.n569 B 0.014973f
C614 VTAIL.n570 B 0.011793f
C615 VTAIL.t2 B 0.032862f
C616 VTAIL.n571 B 0.098419f
C617 VTAIL.n572 B 0.947735f
C618 VTAIL.n573 B 0.008446f
C619 VTAIL.n574 B 0.008943f
C620 VTAIL.n575 B 0.019964f
C621 VTAIL.n576 B 0.019964f
C622 VTAIL.n577 B 0.008943f
C623 VTAIL.n578 B 0.008446f
C624 VTAIL.n579 B 0.015718f
C625 VTAIL.n580 B 0.015718f
C626 VTAIL.n581 B 0.008446f
C627 VTAIL.n582 B 0.008943f
C628 VTAIL.n583 B 0.019964f
C629 VTAIL.n584 B 0.019964f
C630 VTAIL.n585 B 0.008943f
C631 VTAIL.n586 B 0.008446f
C632 VTAIL.n587 B 0.015718f
C633 VTAIL.n588 B 0.015718f
C634 VTAIL.n589 B 0.008446f
C635 VTAIL.n590 B 0.008943f
C636 VTAIL.n591 B 0.019964f
C637 VTAIL.n592 B 0.019964f
C638 VTAIL.n593 B 0.008943f
C639 VTAIL.n594 B 0.008446f
C640 VTAIL.n595 B 0.015718f
C641 VTAIL.n596 B 0.015718f
C642 VTAIL.n597 B 0.008446f
C643 VTAIL.n598 B 0.008943f
C644 VTAIL.n599 B 0.019964f
C645 VTAIL.n600 B 0.019964f
C646 VTAIL.n601 B 0.008943f
C647 VTAIL.n602 B 0.008446f
C648 VTAIL.n603 B 0.015718f
C649 VTAIL.n604 B 0.015718f
C650 VTAIL.n605 B 0.008446f
C651 VTAIL.n606 B 0.008943f
C652 VTAIL.n607 B 0.019964f
C653 VTAIL.n608 B 0.019964f
C654 VTAIL.n609 B 0.008943f
C655 VTAIL.n610 B 0.008446f
C656 VTAIL.n611 B 0.015718f
C657 VTAIL.n612 B 0.015718f
C658 VTAIL.n613 B 0.008446f
C659 VTAIL.n614 B 0.008446f
C660 VTAIL.n615 B 0.008943f
C661 VTAIL.n616 B 0.019964f
C662 VTAIL.n617 B 0.019964f
C663 VTAIL.n618 B 0.039468f
C664 VTAIL.n619 B 0.008695f
C665 VTAIL.n620 B 0.008446f
C666 VTAIL.n621 B 0.037191f
C667 VTAIL.n622 B 0.021725f
C668 VTAIL.n623 B 0.919138f
C669 VN.t3 B 1.69577f
C670 VN.t0 B 1.69561f
C671 VN.n0 B 1.23827f
C672 VN.t1 B 1.69577f
C673 VN.t2 B 1.69561f
C674 VN.n1 B 2.39835f
.ends

