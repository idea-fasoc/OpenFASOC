* NGSPICE file created from diff_pair_sample_0377.ext - technology: sky130A

.subckt diff_pair_sample_0377 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VP.t0 VDD1.t1 B.t5 sky130_fd_pr__nfet_01v8 ad=0.73425 pd=4.78 as=0.73425 ps=4.78 w=4.45 l=2.61
X1 VTAIL.t14 VP.t1 VDD1.t2 B.t4 sky130_fd_pr__nfet_01v8 ad=0.73425 pd=4.78 as=0.73425 ps=4.78 w=4.45 l=2.61
X2 VTAIL.t7 VN.t0 VDD2.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=1.7355 pd=9.68 as=0.73425 ps=4.78 w=4.45 l=2.61
X3 B.t21 B.t19 B.t20 B.t13 sky130_fd_pr__nfet_01v8 ad=1.7355 pd=9.68 as=0 ps=0 w=4.45 l=2.61
X4 VTAIL.t5 VN.t1 VDD2.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=0.73425 pd=4.78 as=0.73425 ps=4.78 w=4.45 l=2.61
X5 VDD1.t5 VP.t2 VTAIL.t13 B.t0 sky130_fd_pr__nfet_01v8 ad=0.73425 pd=4.78 as=0.73425 ps=4.78 w=4.45 l=2.61
X6 B.t18 B.t16 B.t17 B.t9 sky130_fd_pr__nfet_01v8 ad=1.7355 pd=9.68 as=0 ps=0 w=4.45 l=2.61
X7 VDD2.t5 VN.t2 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=0.73425 pd=4.78 as=1.7355 ps=9.68 w=4.45 l=2.61
X8 VTAIL.t1 VN.t3 VDD2.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=1.7355 pd=9.68 as=0.73425 ps=4.78 w=4.45 l=2.61
X9 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=1.7355 pd=9.68 as=0 ps=0 w=4.45 l=2.61
X10 VDD2.t3 VN.t4 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.73425 pd=4.78 as=1.7355 ps=9.68 w=4.45 l=2.61
X11 VTAIL.t12 VP.t3 VDD1.t3 B.t7 sky130_fd_pr__nfet_01v8 ad=1.7355 pd=9.68 as=0.73425 ps=4.78 w=4.45 l=2.61
X12 VTAIL.t4 VN.t5 VDD2.t2 B.t4 sky130_fd_pr__nfet_01v8 ad=0.73425 pd=4.78 as=0.73425 ps=4.78 w=4.45 l=2.61
X13 VDD2.t1 VN.t6 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.73425 pd=4.78 as=0.73425 ps=4.78 w=4.45 l=2.61
X14 VDD1.t6 VP.t4 VTAIL.t11 B.t2 sky130_fd_pr__nfet_01v8 ad=0.73425 pd=4.78 as=1.7355 ps=9.68 w=4.45 l=2.61
X15 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=1.7355 pd=9.68 as=0 ps=0 w=4.45 l=2.61
X16 VTAIL.t10 VP.t5 VDD1.t7 B.t1 sky130_fd_pr__nfet_01v8 ad=1.7355 pd=9.68 as=0.73425 ps=4.78 w=4.45 l=2.61
X17 VDD1.t4 VP.t6 VTAIL.t9 B.t6 sky130_fd_pr__nfet_01v8 ad=0.73425 pd=4.78 as=1.7355 ps=9.68 w=4.45 l=2.61
X18 VDD1.t0 VP.t7 VTAIL.t8 B.t3 sky130_fd_pr__nfet_01v8 ad=0.73425 pd=4.78 as=0.73425 ps=4.78 w=4.45 l=2.61
X19 VDD2.t0 VN.t7 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.73425 pd=4.78 as=0.73425 ps=4.78 w=4.45 l=2.61
R0 VP.n19 VP.n16 161.3
R1 VP.n21 VP.n20 161.3
R2 VP.n22 VP.n15 161.3
R3 VP.n24 VP.n23 161.3
R4 VP.n25 VP.n14 161.3
R5 VP.n27 VP.n26 161.3
R6 VP.n29 VP.n28 161.3
R7 VP.n30 VP.n12 161.3
R8 VP.n32 VP.n31 161.3
R9 VP.n33 VP.n11 161.3
R10 VP.n35 VP.n34 161.3
R11 VP.n36 VP.n10 161.3
R12 VP.n68 VP.n0 161.3
R13 VP.n67 VP.n66 161.3
R14 VP.n65 VP.n1 161.3
R15 VP.n64 VP.n63 161.3
R16 VP.n62 VP.n2 161.3
R17 VP.n61 VP.n60 161.3
R18 VP.n59 VP.n58 161.3
R19 VP.n57 VP.n4 161.3
R20 VP.n56 VP.n55 161.3
R21 VP.n54 VP.n5 161.3
R22 VP.n53 VP.n52 161.3
R23 VP.n51 VP.n6 161.3
R24 VP.n49 VP.n48 161.3
R25 VP.n47 VP.n7 161.3
R26 VP.n46 VP.n45 161.3
R27 VP.n44 VP.n8 161.3
R28 VP.n43 VP.n42 161.3
R29 VP.n41 VP.n9 161.3
R30 VP.n40 VP.n39 102.927
R31 VP.n70 VP.n69 102.927
R32 VP.n38 VP.n37 102.927
R33 VP.n17 VP.t5 74.0585
R34 VP.n18 VP.n17 61.551
R35 VP.n45 VP.n44 56.5193
R36 VP.n56 VP.n5 56.5193
R37 VP.n63 VP.n1 56.5193
R38 VP.n31 VP.n11 56.5193
R39 VP.n24 VP.n15 56.5193
R40 VP.n40 VP.n38 45.2117
R41 VP.n39 VP.t3 41.0905
R42 VP.n50 VP.t2 41.0905
R43 VP.n3 VP.t1 41.0905
R44 VP.n69 VP.t4 41.0905
R45 VP.n37 VP.t6 41.0905
R46 VP.n13 VP.t0 41.0905
R47 VP.n18 VP.t7 41.0905
R48 VP.n43 VP.n9 24.4675
R49 VP.n44 VP.n43 24.4675
R50 VP.n45 VP.n7 24.4675
R51 VP.n49 VP.n7 24.4675
R52 VP.n52 VP.n51 24.4675
R53 VP.n52 VP.n5 24.4675
R54 VP.n57 VP.n56 24.4675
R55 VP.n58 VP.n57 24.4675
R56 VP.n62 VP.n61 24.4675
R57 VP.n63 VP.n62 24.4675
R58 VP.n67 VP.n1 24.4675
R59 VP.n68 VP.n67 24.4675
R60 VP.n35 VP.n11 24.4675
R61 VP.n36 VP.n35 24.4675
R62 VP.n25 VP.n24 24.4675
R63 VP.n26 VP.n25 24.4675
R64 VP.n30 VP.n29 24.4675
R65 VP.n31 VP.n30 24.4675
R66 VP.n20 VP.n19 24.4675
R67 VP.n20 VP.n15 24.4675
R68 VP.n50 VP.n49 13.702
R69 VP.n61 VP.n3 13.702
R70 VP.n29 VP.n13 13.702
R71 VP.n51 VP.n50 10.766
R72 VP.n58 VP.n3 10.766
R73 VP.n26 VP.n13 10.766
R74 VP.n19 VP.n18 10.766
R75 VP.n39 VP.n9 7.82994
R76 VP.n69 VP.n68 7.82994
R77 VP.n37 VP.n36 7.82994
R78 VP.n17 VP.n16 6.98649
R79 VP.n38 VP.n10 0.278367
R80 VP.n41 VP.n40 0.278367
R81 VP.n70 VP.n0 0.278367
R82 VP.n21 VP.n16 0.189894
R83 VP.n22 VP.n21 0.189894
R84 VP.n23 VP.n22 0.189894
R85 VP.n23 VP.n14 0.189894
R86 VP.n27 VP.n14 0.189894
R87 VP.n28 VP.n27 0.189894
R88 VP.n28 VP.n12 0.189894
R89 VP.n32 VP.n12 0.189894
R90 VP.n33 VP.n32 0.189894
R91 VP.n34 VP.n33 0.189894
R92 VP.n34 VP.n10 0.189894
R93 VP.n42 VP.n41 0.189894
R94 VP.n42 VP.n8 0.189894
R95 VP.n46 VP.n8 0.189894
R96 VP.n47 VP.n46 0.189894
R97 VP.n48 VP.n47 0.189894
R98 VP.n48 VP.n6 0.189894
R99 VP.n53 VP.n6 0.189894
R100 VP.n54 VP.n53 0.189894
R101 VP.n55 VP.n54 0.189894
R102 VP.n55 VP.n4 0.189894
R103 VP.n59 VP.n4 0.189894
R104 VP.n60 VP.n59 0.189894
R105 VP.n60 VP.n2 0.189894
R106 VP.n64 VP.n2 0.189894
R107 VP.n65 VP.n64 0.189894
R108 VP.n66 VP.n65 0.189894
R109 VP.n66 VP.n0 0.189894
R110 VP VP.n70 0.153454
R111 VDD1 VDD1.n0 69.8339
R112 VDD1.n3 VDD1.n2 69.7202
R113 VDD1.n3 VDD1.n1 69.7202
R114 VDD1.n5 VDD1.n4 68.5083
R115 VDD1.n5 VDD1.n3 39.5397
R116 VDD1.n4 VDD1.t1 4.44994
R117 VDD1.n4 VDD1.t4 4.44994
R118 VDD1.n0 VDD1.t7 4.44994
R119 VDD1.n0 VDD1.t0 4.44994
R120 VDD1.n2 VDD1.t2 4.44994
R121 VDD1.n2 VDD1.t6 4.44994
R122 VDD1.n1 VDD1.t3 4.44994
R123 VDD1.n1 VDD1.t5 4.44994
R124 VDD1 VDD1.n5 1.20955
R125 VTAIL.n194 VTAIL.n176 289.615
R126 VTAIL.n20 VTAIL.n2 289.615
R127 VTAIL.n44 VTAIL.n26 289.615
R128 VTAIL.n70 VTAIL.n52 289.615
R129 VTAIL.n170 VTAIL.n152 289.615
R130 VTAIL.n144 VTAIL.n126 289.615
R131 VTAIL.n120 VTAIL.n102 289.615
R132 VTAIL.n94 VTAIL.n76 289.615
R133 VTAIL.n185 VTAIL.n184 185
R134 VTAIL.n187 VTAIL.n186 185
R135 VTAIL.n180 VTAIL.n179 185
R136 VTAIL.n193 VTAIL.n192 185
R137 VTAIL.n195 VTAIL.n194 185
R138 VTAIL.n11 VTAIL.n10 185
R139 VTAIL.n13 VTAIL.n12 185
R140 VTAIL.n6 VTAIL.n5 185
R141 VTAIL.n19 VTAIL.n18 185
R142 VTAIL.n21 VTAIL.n20 185
R143 VTAIL.n35 VTAIL.n34 185
R144 VTAIL.n37 VTAIL.n36 185
R145 VTAIL.n30 VTAIL.n29 185
R146 VTAIL.n43 VTAIL.n42 185
R147 VTAIL.n45 VTAIL.n44 185
R148 VTAIL.n61 VTAIL.n60 185
R149 VTAIL.n63 VTAIL.n62 185
R150 VTAIL.n56 VTAIL.n55 185
R151 VTAIL.n69 VTAIL.n68 185
R152 VTAIL.n71 VTAIL.n70 185
R153 VTAIL.n171 VTAIL.n170 185
R154 VTAIL.n169 VTAIL.n168 185
R155 VTAIL.n156 VTAIL.n155 185
R156 VTAIL.n163 VTAIL.n162 185
R157 VTAIL.n161 VTAIL.n160 185
R158 VTAIL.n145 VTAIL.n144 185
R159 VTAIL.n143 VTAIL.n142 185
R160 VTAIL.n130 VTAIL.n129 185
R161 VTAIL.n137 VTAIL.n136 185
R162 VTAIL.n135 VTAIL.n134 185
R163 VTAIL.n121 VTAIL.n120 185
R164 VTAIL.n119 VTAIL.n118 185
R165 VTAIL.n106 VTAIL.n105 185
R166 VTAIL.n113 VTAIL.n112 185
R167 VTAIL.n111 VTAIL.n110 185
R168 VTAIL.n95 VTAIL.n94 185
R169 VTAIL.n93 VTAIL.n92 185
R170 VTAIL.n80 VTAIL.n79 185
R171 VTAIL.n87 VTAIL.n86 185
R172 VTAIL.n85 VTAIL.n84 185
R173 VTAIL.n183 VTAIL.t6 147.714
R174 VTAIL.n9 VTAIL.t1 147.714
R175 VTAIL.n33 VTAIL.t11 147.714
R176 VTAIL.n59 VTAIL.t12 147.714
R177 VTAIL.n159 VTAIL.t9 147.714
R178 VTAIL.n133 VTAIL.t10 147.714
R179 VTAIL.n109 VTAIL.t2 147.714
R180 VTAIL.n83 VTAIL.t7 147.714
R181 VTAIL.n186 VTAIL.n185 104.615
R182 VTAIL.n186 VTAIL.n179 104.615
R183 VTAIL.n193 VTAIL.n179 104.615
R184 VTAIL.n194 VTAIL.n193 104.615
R185 VTAIL.n12 VTAIL.n11 104.615
R186 VTAIL.n12 VTAIL.n5 104.615
R187 VTAIL.n19 VTAIL.n5 104.615
R188 VTAIL.n20 VTAIL.n19 104.615
R189 VTAIL.n36 VTAIL.n35 104.615
R190 VTAIL.n36 VTAIL.n29 104.615
R191 VTAIL.n43 VTAIL.n29 104.615
R192 VTAIL.n44 VTAIL.n43 104.615
R193 VTAIL.n62 VTAIL.n61 104.615
R194 VTAIL.n62 VTAIL.n55 104.615
R195 VTAIL.n69 VTAIL.n55 104.615
R196 VTAIL.n70 VTAIL.n69 104.615
R197 VTAIL.n170 VTAIL.n169 104.615
R198 VTAIL.n169 VTAIL.n155 104.615
R199 VTAIL.n162 VTAIL.n155 104.615
R200 VTAIL.n162 VTAIL.n161 104.615
R201 VTAIL.n144 VTAIL.n143 104.615
R202 VTAIL.n143 VTAIL.n129 104.615
R203 VTAIL.n136 VTAIL.n129 104.615
R204 VTAIL.n136 VTAIL.n135 104.615
R205 VTAIL.n120 VTAIL.n119 104.615
R206 VTAIL.n119 VTAIL.n105 104.615
R207 VTAIL.n112 VTAIL.n105 104.615
R208 VTAIL.n112 VTAIL.n111 104.615
R209 VTAIL.n94 VTAIL.n93 104.615
R210 VTAIL.n93 VTAIL.n79 104.615
R211 VTAIL.n86 VTAIL.n79 104.615
R212 VTAIL.n86 VTAIL.n85 104.615
R213 VTAIL.n185 VTAIL.t6 52.3082
R214 VTAIL.n11 VTAIL.t1 52.3082
R215 VTAIL.n35 VTAIL.t11 52.3082
R216 VTAIL.n61 VTAIL.t12 52.3082
R217 VTAIL.n161 VTAIL.t9 52.3082
R218 VTAIL.n135 VTAIL.t10 52.3082
R219 VTAIL.n111 VTAIL.t2 52.3082
R220 VTAIL.n85 VTAIL.t7 52.3082
R221 VTAIL.n151 VTAIL.n150 51.8297
R222 VTAIL.n101 VTAIL.n100 51.8297
R223 VTAIL.n1 VTAIL.n0 51.8295
R224 VTAIL.n51 VTAIL.n50 51.8295
R225 VTAIL.n199 VTAIL.n198 30.052
R226 VTAIL.n25 VTAIL.n24 30.052
R227 VTAIL.n49 VTAIL.n48 30.052
R228 VTAIL.n75 VTAIL.n74 30.052
R229 VTAIL.n175 VTAIL.n174 30.052
R230 VTAIL.n149 VTAIL.n148 30.052
R231 VTAIL.n125 VTAIL.n124 30.052
R232 VTAIL.n99 VTAIL.n98 30.052
R233 VTAIL.n199 VTAIL.n175 18.7376
R234 VTAIL.n99 VTAIL.n75 18.7376
R235 VTAIL.n184 VTAIL.n183 15.6631
R236 VTAIL.n10 VTAIL.n9 15.6631
R237 VTAIL.n34 VTAIL.n33 15.6631
R238 VTAIL.n60 VTAIL.n59 15.6631
R239 VTAIL.n160 VTAIL.n159 15.6631
R240 VTAIL.n134 VTAIL.n133 15.6631
R241 VTAIL.n110 VTAIL.n109 15.6631
R242 VTAIL.n84 VTAIL.n83 15.6631
R243 VTAIL.n187 VTAIL.n182 12.8005
R244 VTAIL.n13 VTAIL.n8 12.8005
R245 VTAIL.n37 VTAIL.n32 12.8005
R246 VTAIL.n63 VTAIL.n58 12.8005
R247 VTAIL.n163 VTAIL.n158 12.8005
R248 VTAIL.n137 VTAIL.n132 12.8005
R249 VTAIL.n113 VTAIL.n108 12.8005
R250 VTAIL.n87 VTAIL.n82 12.8005
R251 VTAIL.n188 VTAIL.n180 12.0247
R252 VTAIL.n14 VTAIL.n6 12.0247
R253 VTAIL.n38 VTAIL.n30 12.0247
R254 VTAIL.n64 VTAIL.n56 12.0247
R255 VTAIL.n164 VTAIL.n156 12.0247
R256 VTAIL.n138 VTAIL.n130 12.0247
R257 VTAIL.n114 VTAIL.n106 12.0247
R258 VTAIL.n88 VTAIL.n80 12.0247
R259 VTAIL.n192 VTAIL.n191 11.249
R260 VTAIL.n18 VTAIL.n17 11.249
R261 VTAIL.n42 VTAIL.n41 11.249
R262 VTAIL.n68 VTAIL.n67 11.249
R263 VTAIL.n168 VTAIL.n167 11.249
R264 VTAIL.n142 VTAIL.n141 11.249
R265 VTAIL.n118 VTAIL.n117 11.249
R266 VTAIL.n92 VTAIL.n91 11.249
R267 VTAIL.n195 VTAIL.n178 10.4732
R268 VTAIL.n21 VTAIL.n4 10.4732
R269 VTAIL.n45 VTAIL.n28 10.4732
R270 VTAIL.n71 VTAIL.n54 10.4732
R271 VTAIL.n171 VTAIL.n154 10.4732
R272 VTAIL.n145 VTAIL.n128 10.4732
R273 VTAIL.n121 VTAIL.n104 10.4732
R274 VTAIL.n95 VTAIL.n78 10.4732
R275 VTAIL.n196 VTAIL.n176 9.69747
R276 VTAIL.n22 VTAIL.n2 9.69747
R277 VTAIL.n46 VTAIL.n26 9.69747
R278 VTAIL.n72 VTAIL.n52 9.69747
R279 VTAIL.n172 VTAIL.n152 9.69747
R280 VTAIL.n146 VTAIL.n126 9.69747
R281 VTAIL.n122 VTAIL.n102 9.69747
R282 VTAIL.n96 VTAIL.n76 9.69747
R283 VTAIL.n198 VTAIL.n197 9.45567
R284 VTAIL.n24 VTAIL.n23 9.45567
R285 VTAIL.n48 VTAIL.n47 9.45567
R286 VTAIL.n74 VTAIL.n73 9.45567
R287 VTAIL.n174 VTAIL.n173 9.45567
R288 VTAIL.n148 VTAIL.n147 9.45567
R289 VTAIL.n124 VTAIL.n123 9.45567
R290 VTAIL.n98 VTAIL.n97 9.45567
R291 VTAIL.n197 VTAIL.n196 9.3005
R292 VTAIL.n178 VTAIL.n177 9.3005
R293 VTAIL.n191 VTAIL.n190 9.3005
R294 VTAIL.n189 VTAIL.n188 9.3005
R295 VTAIL.n182 VTAIL.n181 9.3005
R296 VTAIL.n23 VTAIL.n22 9.3005
R297 VTAIL.n4 VTAIL.n3 9.3005
R298 VTAIL.n17 VTAIL.n16 9.3005
R299 VTAIL.n15 VTAIL.n14 9.3005
R300 VTAIL.n8 VTAIL.n7 9.3005
R301 VTAIL.n47 VTAIL.n46 9.3005
R302 VTAIL.n28 VTAIL.n27 9.3005
R303 VTAIL.n41 VTAIL.n40 9.3005
R304 VTAIL.n39 VTAIL.n38 9.3005
R305 VTAIL.n32 VTAIL.n31 9.3005
R306 VTAIL.n73 VTAIL.n72 9.3005
R307 VTAIL.n54 VTAIL.n53 9.3005
R308 VTAIL.n67 VTAIL.n66 9.3005
R309 VTAIL.n65 VTAIL.n64 9.3005
R310 VTAIL.n58 VTAIL.n57 9.3005
R311 VTAIL.n173 VTAIL.n172 9.3005
R312 VTAIL.n154 VTAIL.n153 9.3005
R313 VTAIL.n167 VTAIL.n166 9.3005
R314 VTAIL.n165 VTAIL.n164 9.3005
R315 VTAIL.n158 VTAIL.n157 9.3005
R316 VTAIL.n147 VTAIL.n146 9.3005
R317 VTAIL.n128 VTAIL.n127 9.3005
R318 VTAIL.n141 VTAIL.n140 9.3005
R319 VTAIL.n139 VTAIL.n138 9.3005
R320 VTAIL.n132 VTAIL.n131 9.3005
R321 VTAIL.n123 VTAIL.n122 9.3005
R322 VTAIL.n104 VTAIL.n103 9.3005
R323 VTAIL.n117 VTAIL.n116 9.3005
R324 VTAIL.n115 VTAIL.n114 9.3005
R325 VTAIL.n108 VTAIL.n107 9.3005
R326 VTAIL.n97 VTAIL.n96 9.3005
R327 VTAIL.n78 VTAIL.n77 9.3005
R328 VTAIL.n91 VTAIL.n90 9.3005
R329 VTAIL.n89 VTAIL.n88 9.3005
R330 VTAIL.n82 VTAIL.n81 9.3005
R331 VTAIL.n0 VTAIL.t3 4.44994
R332 VTAIL.n0 VTAIL.t5 4.44994
R333 VTAIL.n50 VTAIL.t13 4.44994
R334 VTAIL.n50 VTAIL.t14 4.44994
R335 VTAIL.n150 VTAIL.t8 4.44994
R336 VTAIL.n150 VTAIL.t15 4.44994
R337 VTAIL.n100 VTAIL.t0 4.44994
R338 VTAIL.n100 VTAIL.t4 4.44994
R339 VTAIL.n183 VTAIL.n181 4.39059
R340 VTAIL.n9 VTAIL.n7 4.39059
R341 VTAIL.n33 VTAIL.n31 4.39059
R342 VTAIL.n59 VTAIL.n57 4.39059
R343 VTAIL.n159 VTAIL.n157 4.39059
R344 VTAIL.n133 VTAIL.n131 4.39059
R345 VTAIL.n109 VTAIL.n107 4.39059
R346 VTAIL.n83 VTAIL.n81 4.39059
R347 VTAIL.n198 VTAIL.n176 4.26717
R348 VTAIL.n24 VTAIL.n2 4.26717
R349 VTAIL.n48 VTAIL.n26 4.26717
R350 VTAIL.n74 VTAIL.n52 4.26717
R351 VTAIL.n174 VTAIL.n152 4.26717
R352 VTAIL.n148 VTAIL.n126 4.26717
R353 VTAIL.n124 VTAIL.n102 4.26717
R354 VTAIL.n98 VTAIL.n76 4.26717
R355 VTAIL.n196 VTAIL.n195 3.49141
R356 VTAIL.n22 VTAIL.n21 3.49141
R357 VTAIL.n46 VTAIL.n45 3.49141
R358 VTAIL.n72 VTAIL.n71 3.49141
R359 VTAIL.n172 VTAIL.n171 3.49141
R360 VTAIL.n146 VTAIL.n145 3.49141
R361 VTAIL.n122 VTAIL.n121 3.49141
R362 VTAIL.n96 VTAIL.n95 3.49141
R363 VTAIL.n192 VTAIL.n178 2.71565
R364 VTAIL.n18 VTAIL.n4 2.71565
R365 VTAIL.n42 VTAIL.n28 2.71565
R366 VTAIL.n68 VTAIL.n54 2.71565
R367 VTAIL.n168 VTAIL.n154 2.71565
R368 VTAIL.n142 VTAIL.n128 2.71565
R369 VTAIL.n118 VTAIL.n104 2.71565
R370 VTAIL.n92 VTAIL.n78 2.71565
R371 VTAIL.n101 VTAIL.n99 2.53498
R372 VTAIL.n125 VTAIL.n101 2.53498
R373 VTAIL.n151 VTAIL.n149 2.53498
R374 VTAIL.n175 VTAIL.n151 2.53498
R375 VTAIL.n75 VTAIL.n51 2.53498
R376 VTAIL.n51 VTAIL.n49 2.53498
R377 VTAIL.n25 VTAIL.n1 2.53498
R378 VTAIL VTAIL.n199 2.47679
R379 VTAIL.n191 VTAIL.n180 1.93989
R380 VTAIL.n17 VTAIL.n6 1.93989
R381 VTAIL.n41 VTAIL.n30 1.93989
R382 VTAIL.n67 VTAIL.n56 1.93989
R383 VTAIL.n167 VTAIL.n156 1.93989
R384 VTAIL.n141 VTAIL.n130 1.93989
R385 VTAIL.n117 VTAIL.n106 1.93989
R386 VTAIL.n91 VTAIL.n80 1.93989
R387 VTAIL.n188 VTAIL.n187 1.16414
R388 VTAIL.n14 VTAIL.n13 1.16414
R389 VTAIL.n38 VTAIL.n37 1.16414
R390 VTAIL.n64 VTAIL.n63 1.16414
R391 VTAIL.n164 VTAIL.n163 1.16414
R392 VTAIL.n138 VTAIL.n137 1.16414
R393 VTAIL.n114 VTAIL.n113 1.16414
R394 VTAIL.n88 VTAIL.n87 1.16414
R395 VTAIL.n149 VTAIL.n125 0.470328
R396 VTAIL.n49 VTAIL.n25 0.470328
R397 VTAIL.n184 VTAIL.n182 0.388379
R398 VTAIL.n10 VTAIL.n8 0.388379
R399 VTAIL.n34 VTAIL.n32 0.388379
R400 VTAIL.n60 VTAIL.n58 0.388379
R401 VTAIL.n160 VTAIL.n158 0.388379
R402 VTAIL.n134 VTAIL.n132 0.388379
R403 VTAIL.n110 VTAIL.n108 0.388379
R404 VTAIL.n84 VTAIL.n82 0.388379
R405 VTAIL.n189 VTAIL.n181 0.155672
R406 VTAIL.n190 VTAIL.n189 0.155672
R407 VTAIL.n190 VTAIL.n177 0.155672
R408 VTAIL.n197 VTAIL.n177 0.155672
R409 VTAIL.n15 VTAIL.n7 0.155672
R410 VTAIL.n16 VTAIL.n15 0.155672
R411 VTAIL.n16 VTAIL.n3 0.155672
R412 VTAIL.n23 VTAIL.n3 0.155672
R413 VTAIL.n39 VTAIL.n31 0.155672
R414 VTAIL.n40 VTAIL.n39 0.155672
R415 VTAIL.n40 VTAIL.n27 0.155672
R416 VTAIL.n47 VTAIL.n27 0.155672
R417 VTAIL.n65 VTAIL.n57 0.155672
R418 VTAIL.n66 VTAIL.n65 0.155672
R419 VTAIL.n66 VTAIL.n53 0.155672
R420 VTAIL.n73 VTAIL.n53 0.155672
R421 VTAIL.n173 VTAIL.n153 0.155672
R422 VTAIL.n166 VTAIL.n153 0.155672
R423 VTAIL.n166 VTAIL.n165 0.155672
R424 VTAIL.n165 VTAIL.n157 0.155672
R425 VTAIL.n147 VTAIL.n127 0.155672
R426 VTAIL.n140 VTAIL.n127 0.155672
R427 VTAIL.n140 VTAIL.n139 0.155672
R428 VTAIL.n139 VTAIL.n131 0.155672
R429 VTAIL.n123 VTAIL.n103 0.155672
R430 VTAIL.n116 VTAIL.n103 0.155672
R431 VTAIL.n116 VTAIL.n115 0.155672
R432 VTAIL.n115 VTAIL.n107 0.155672
R433 VTAIL.n97 VTAIL.n77 0.155672
R434 VTAIL.n90 VTAIL.n77 0.155672
R435 VTAIL.n90 VTAIL.n89 0.155672
R436 VTAIL.n89 VTAIL.n81 0.155672
R437 VTAIL VTAIL.n1 0.0586897
R438 B.n661 B.n660 585
R439 B.n215 B.n119 585
R440 B.n214 B.n213 585
R441 B.n212 B.n211 585
R442 B.n210 B.n209 585
R443 B.n208 B.n207 585
R444 B.n206 B.n205 585
R445 B.n204 B.n203 585
R446 B.n202 B.n201 585
R447 B.n200 B.n199 585
R448 B.n198 B.n197 585
R449 B.n196 B.n195 585
R450 B.n194 B.n193 585
R451 B.n192 B.n191 585
R452 B.n190 B.n189 585
R453 B.n188 B.n187 585
R454 B.n186 B.n185 585
R455 B.n184 B.n183 585
R456 B.n182 B.n181 585
R457 B.n179 B.n178 585
R458 B.n177 B.n176 585
R459 B.n175 B.n174 585
R460 B.n173 B.n172 585
R461 B.n171 B.n170 585
R462 B.n169 B.n168 585
R463 B.n167 B.n166 585
R464 B.n165 B.n164 585
R465 B.n163 B.n162 585
R466 B.n161 B.n160 585
R467 B.n158 B.n157 585
R468 B.n156 B.n155 585
R469 B.n154 B.n153 585
R470 B.n152 B.n151 585
R471 B.n150 B.n149 585
R472 B.n148 B.n147 585
R473 B.n146 B.n145 585
R474 B.n144 B.n143 585
R475 B.n142 B.n141 585
R476 B.n140 B.n139 585
R477 B.n138 B.n137 585
R478 B.n136 B.n135 585
R479 B.n134 B.n133 585
R480 B.n132 B.n131 585
R481 B.n130 B.n129 585
R482 B.n128 B.n127 585
R483 B.n126 B.n125 585
R484 B.n96 B.n95 585
R485 B.n666 B.n665 585
R486 B.n659 B.n120 585
R487 B.n120 B.n93 585
R488 B.n658 B.n92 585
R489 B.n670 B.n92 585
R490 B.n657 B.n91 585
R491 B.n671 B.n91 585
R492 B.n656 B.n90 585
R493 B.n672 B.n90 585
R494 B.n655 B.n654 585
R495 B.n654 B.n86 585
R496 B.n653 B.n85 585
R497 B.n678 B.n85 585
R498 B.n652 B.n84 585
R499 B.n679 B.n84 585
R500 B.n651 B.n83 585
R501 B.n680 B.n83 585
R502 B.n650 B.n649 585
R503 B.n649 B.n79 585
R504 B.n648 B.n78 585
R505 B.n686 B.n78 585
R506 B.n647 B.n77 585
R507 B.n687 B.n77 585
R508 B.n646 B.n76 585
R509 B.n688 B.n76 585
R510 B.n645 B.n644 585
R511 B.n644 B.n72 585
R512 B.n643 B.n71 585
R513 B.n694 B.n71 585
R514 B.n642 B.n70 585
R515 B.n695 B.n70 585
R516 B.n641 B.n69 585
R517 B.n696 B.n69 585
R518 B.n640 B.n639 585
R519 B.n639 B.n65 585
R520 B.n638 B.n64 585
R521 B.n702 B.n64 585
R522 B.n637 B.n63 585
R523 B.n703 B.n63 585
R524 B.n636 B.n62 585
R525 B.n704 B.n62 585
R526 B.n635 B.n634 585
R527 B.n634 B.n58 585
R528 B.n633 B.n57 585
R529 B.n710 B.n57 585
R530 B.n632 B.n56 585
R531 B.n711 B.n56 585
R532 B.n631 B.n55 585
R533 B.n712 B.n55 585
R534 B.n630 B.n629 585
R535 B.n629 B.n51 585
R536 B.n628 B.n50 585
R537 B.n718 B.n50 585
R538 B.n627 B.n49 585
R539 B.n719 B.n49 585
R540 B.n626 B.n48 585
R541 B.n720 B.n48 585
R542 B.n625 B.n624 585
R543 B.n624 B.n47 585
R544 B.n623 B.n43 585
R545 B.n726 B.n43 585
R546 B.n622 B.n42 585
R547 B.n727 B.n42 585
R548 B.n621 B.n41 585
R549 B.n728 B.n41 585
R550 B.n620 B.n619 585
R551 B.n619 B.n37 585
R552 B.n618 B.n36 585
R553 B.n734 B.n36 585
R554 B.n617 B.n35 585
R555 B.n735 B.n35 585
R556 B.n616 B.n34 585
R557 B.n736 B.n34 585
R558 B.n615 B.n614 585
R559 B.n614 B.n33 585
R560 B.n613 B.n29 585
R561 B.n742 B.n29 585
R562 B.n612 B.n28 585
R563 B.n743 B.n28 585
R564 B.n611 B.n27 585
R565 B.n744 B.n27 585
R566 B.n610 B.n609 585
R567 B.n609 B.n23 585
R568 B.n608 B.n22 585
R569 B.n750 B.n22 585
R570 B.n607 B.n21 585
R571 B.n751 B.n21 585
R572 B.n606 B.n20 585
R573 B.n752 B.n20 585
R574 B.n605 B.n604 585
R575 B.n604 B.n16 585
R576 B.n603 B.n15 585
R577 B.n758 B.n15 585
R578 B.n602 B.n14 585
R579 B.n759 B.n14 585
R580 B.n601 B.n13 585
R581 B.n760 B.n13 585
R582 B.n600 B.n599 585
R583 B.n599 B.n12 585
R584 B.n598 B.n597 585
R585 B.n598 B.n8 585
R586 B.n596 B.n7 585
R587 B.n767 B.n7 585
R588 B.n595 B.n6 585
R589 B.n768 B.n6 585
R590 B.n594 B.n5 585
R591 B.n769 B.n5 585
R592 B.n593 B.n592 585
R593 B.n592 B.n4 585
R594 B.n591 B.n216 585
R595 B.n591 B.n590 585
R596 B.n581 B.n217 585
R597 B.n218 B.n217 585
R598 B.n583 B.n582 585
R599 B.n584 B.n583 585
R600 B.n580 B.n223 585
R601 B.n223 B.n222 585
R602 B.n579 B.n578 585
R603 B.n578 B.n577 585
R604 B.n225 B.n224 585
R605 B.n226 B.n225 585
R606 B.n570 B.n569 585
R607 B.n571 B.n570 585
R608 B.n568 B.n231 585
R609 B.n231 B.n230 585
R610 B.n567 B.n566 585
R611 B.n566 B.n565 585
R612 B.n233 B.n232 585
R613 B.n234 B.n233 585
R614 B.n558 B.n557 585
R615 B.n559 B.n558 585
R616 B.n556 B.n239 585
R617 B.n239 B.n238 585
R618 B.n555 B.n554 585
R619 B.n554 B.n553 585
R620 B.n241 B.n240 585
R621 B.n546 B.n241 585
R622 B.n545 B.n544 585
R623 B.n547 B.n545 585
R624 B.n543 B.n246 585
R625 B.n246 B.n245 585
R626 B.n542 B.n541 585
R627 B.n541 B.n540 585
R628 B.n248 B.n247 585
R629 B.n249 B.n248 585
R630 B.n533 B.n532 585
R631 B.n534 B.n533 585
R632 B.n531 B.n254 585
R633 B.n254 B.n253 585
R634 B.n530 B.n529 585
R635 B.n529 B.n528 585
R636 B.n256 B.n255 585
R637 B.n521 B.n256 585
R638 B.n520 B.n519 585
R639 B.n522 B.n520 585
R640 B.n518 B.n261 585
R641 B.n261 B.n260 585
R642 B.n517 B.n516 585
R643 B.n516 B.n515 585
R644 B.n263 B.n262 585
R645 B.n264 B.n263 585
R646 B.n508 B.n507 585
R647 B.n509 B.n508 585
R648 B.n506 B.n269 585
R649 B.n269 B.n268 585
R650 B.n505 B.n504 585
R651 B.n504 B.n503 585
R652 B.n271 B.n270 585
R653 B.n272 B.n271 585
R654 B.n496 B.n495 585
R655 B.n497 B.n496 585
R656 B.n494 B.n277 585
R657 B.n277 B.n276 585
R658 B.n493 B.n492 585
R659 B.n492 B.n491 585
R660 B.n279 B.n278 585
R661 B.n280 B.n279 585
R662 B.n484 B.n483 585
R663 B.n485 B.n484 585
R664 B.n482 B.n285 585
R665 B.n285 B.n284 585
R666 B.n481 B.n480 585
R667 B.n480 B.n479 585
R668 B.n287 B.n286 585
R669 B.n288 B.n287 585
R670 B.n472 B.n471 585
R671 B.n473 B.n472 585
R672 B.n470 B.n293 585
R673 B.n293 B.n292 585
R674 B.n469 B.n468 585
R675 B.n468 B.n467 585
R676 B.n295 B.n294 585
R677 B.n296 B.n295 585
R678 B.n460 B.n459 585
R679 B.n461 B.n460 585
R680 B.n458 B.n301 585
R681 B.n301 B.n300 585
R682 B.n457 B.n456 585
R683 B.n456 B.n455 585
R684 B.n303 B.n302 585
R685 B.n304 B.n303 585
R686 B.n448 B.n447 585
R687 B.n449 B.n448 585
R688 B.n446 B.n309 585
R689 B.n309 B.n308 585
R690 B.n445 B.n444 585
R691 B.n444 B.n443 585
R692 B.n311 B.n310 585
R693 B.n312 B.n311 585
R694 B.n439 B.n438 585
R695 B.n315 B.n314 585
R696 B.n435 B.n434 585
R697 B.n436 B.n435 585
R698 B.n433 B.n339 585
R699 B.n432 B.n431 585
R700 B.n430 B.n429 585
R701 B.n428 B.n427 585
R702 B.n426 B.n425 585
R703 B.n424 B.n423 585
R704 B.n422 B.n421 585
R705 B.n420 B.n419 585
R706 B.n418 B.n417 585
R707 B.n416 B.n415 585
R708 B.n414 B.n413 585
R709 B.n412 B.n411 585
R710 B.n410 B.n409 585
R711 B.n408 B.n407 585
R712 B.n406 B.n405 585
R713 B.n404 B.n403 585
R714 B.n402 B.n401 585
R715 B.n400 B.n399 585
R716 B.n398 B.n397 585
R717 B.n396 B.n395 585
R718 B.n394 B.n393 585
R719 B.n392 B.n391 585
R720 B.n390 B.n389 585
R721 B.n388 B.n387 585
R722 B.n386 B.n385 585
R723 B.n384 B.n383 585
R724 B.n382 B.n381 585
R725 B.n380 B.n379 585
R726 B.n378 B.n377 585
R727 B.n376 B.n375 585
R728 B.n374 B.n373 585
R729 B.n372 B.n371 585
R730 B.n370 B.n369 585
R731 B.n368 B.n367 585
R732 B.n366 B.n365 585
R733 B.n364 B.n363 585
R734 B.n362 B.n361 585
R735 B.n360 B.n359 585
R736 B.n358 B.n357 585
R737 B.n356 B.n355 585
R738 B.n354 B.n353 585
R739 B.n352 B.n351 585
R740 B.n350 B.n349 585
R741 B.n348 B.n347 585
R742 B.n346 B.n338 585
R743 B.n436 B.n338 585
R744 B.n440 B.n313 585
R745 B.n313 B.n312 585
R746 B.n442 B.n441 585
R747 B.n443 B.n442 585
R748 B.n307 B.n306 585
R749 B.n308 B.n307 585
R750 B.n451 B.n450 585
R751 B.n450 B.n449 585
R752 B.n452 B.n305 585
R753 B.n305 B.n304 585
R754 B.n454 B.n453 585
R755 B.n455 B.n454 585
R756 B.n299 B.n298 585
R757 B.n300 B.n299 585
R758 B.n463 B.n462 585
R759 B.n462 B.n461 585
R760 B.n464 B.n297 585
R761 B.n297 B.n296 585
R762 B.n466 B.n465 585
R763 B.n467 B.n466 585
R764 B.n291 B.n290 585
R765 B.n292 B.n291 585
R766 B.n475 B.n474 585
R767 B.n474 B.n473 585
R768 B.n476 B.n289 585
R769 B.n289 B.n288 585
R770 B.n478 B.n477 585
R771 B.n479 B.n478 585
R772 B.n283 B.n282 585
R773 B.n284 B.n283 585
R774 B.n487 B.n486 585
R775 B.n486 B.n485 585
R776 B.n488 B.n281 585
R777 B.n281 B.n280 585
R778 B.n490 B.n489 585
R779 B.n491 B.n490 585
R780 B.n275 B.n274 585
R781 B.n276 B.n275 585
R782 B.n499 B.n498 585
R783 B.n498 B.n497 585
R784 B.n500 B.n273 585
R785 B.n273 B.n272 585
R786 B.n502 B.n501 585
R787 B.n503 B.n502 585
R788 B.n267 B.n266 585
R789 B.n268 B.n267 585
R790 B.n511 B.n510 585
R791 B.n510 B.n509 585
R792 B.n512 B.n265 585
R793 B.n265 B.n264 585
R794 B.n514 B.n513 585
R795 B.n515 B.n514 585
R796 B.n259 B.n258 585
R797 B.n260 B.n259 585
R798 B.n524 B.n523 585
R799 B.n523 B.n522 585
R800 B.n525 B.n257 585
R801 B.n521 B.n257 585
R802 B.n527 B.n526 585
R803 B.n528 B.n527 585
R804 B.n252 B.n251 585
R805 B.n253 B.n252 585
R806 B.n536 B.n535 585
R807 B.n535 B.n534 585
R808 B.n537 B.n250 585
R809 B.n250 B.n249 585
R810 B.n539 B.n538 585
R811 B.n540 B.n539 585
R812 B.n244 B.n243 585
R813 B.n245 B.n244 585
R814 B.n549 B.n548 585
R815 B.n548 B.n547 585
R816 B.n550 B.n242 585
R817 B.n546 B.n242 585
R818 B.n552 B.n551 585
R819 B.n553 B.n552 585
R820 B.n237 B.n236 585
R821 B.n238 B.n237 585
R822 B.n561 B.n560 585
R823 B.n560 B.n559 585
R824 B.n562 B.n235 585
R825 B.n235 B.n234 585
R826 B.n564 B.n563 585
R827 B.n565 B.n564 585
R828 B.n229 B.n228 585
R829 B.n230 B.n229 585
R830 B.n573 B.n572 585
R831 B.n572 B.n571 585
R832 B.n574 B.n227 585
R833 B.n227 B.n226 585
R834 B.n576 B.n575 585
R835 B.n577 B.n576 585
R836 B.n221 B.n220 585
R837 B.n222 B.n221 585
R838 B.n586 B.n585 585
R839 B.n585 B.n584 585
R840 B.n587 B.n219 585
R841 B.n219 B.n218 585
R842 B.n589 B.n588 585
R843 B.n590 B.n589 585
R844 B.n3 B.n0 585
R845 B.n4 B.n3 585
R846 B.n766 B.n1 585
R847 B.n767 B.n766 585
R848 B.n765 B.n764 585
R849 B.n765 B.n8 585
R850 B.n763 B.n9 585
R851 B.n12 B.n9 585
R852 B.n762 B.n761 585
R853 B.n761 B.n760 585
R854 B.n11 B.n10 585
R855 B.n759 B.n11 585
R856 B.n757 B.n756 585
R857 B.n758 B.n757 585
R858 B.n755 B.n17 585
R859 B.n17 B.n16 585
R860 B.n754 B.n753 585
R861 B.n753 B.n752 585
R862 B.n19 B.n18 585
R863 B.n751 B.n19 585
R864 B.n749 B.n748 585
R865 B.n750 B.n749 585
R866 B.n747 B.n24 585
R867 B.n24 B.n23 585
R868 B.n746 B.n745 585
R869 B.n745 B.n744 585
R870 B.n26 B.n25 585
R871 B.n743 B.n26 585
R872 B.n741 B.n740 585
R873 B.n742 B.n741 585
R874 B.n739 B.n30 585
R875 B.n33 B.n30 585
R876 B.n738 B.n737 585
R877 B.n737 B.n736 585
R878 B.n32 B.n31 585
R879 B.n735 B.n32 585
R880 B.n733 B.n732 585
R881 B.n734 B.n733 585
R882 B.n731 B.n38 585
R883 B.n38 B.n37 585
R884 B.n730 B.n729 585
R885 B.n729 B.n728 585
R886 B.n40 B.n39 585
R887 B.n727 B.n40 585
R888 B.n725 B.n724 585
R889 B.n726 B.n725 585
R890 B.n723 B.n44 585
R891 B.n47 B.n44 585
R892 B.n722 B.n721 585
R893 B.n721 B.n720 585
R894 B.n46 B.n45 585
R895 B.n719 B.n46 585
R896 B.n717 B.n716 585
R897 B.n718 B.n717 585
R898 B.n715 B.n52 585
R899 B.n52 B.n51 585
R900 B.n714 B.n713 585
R901 B.n713 B.n712 585
R902 B.n54 B.n53 585
R903 B.n711 B.n54 585
R904 B.n709 B.n708 585
R905 B.n710 B.n709 585
R906 B.n707 B.n59 585
R907 B.n59 B.n58 585
R908 B.n706 B.n705 585
R909 B.n705 B.n704 585
R910 B.n61 B.n60 585
R911 B.n703 B.n61 585
R912 B.n701 B.n700 585
R913 B.n702 B.n701 585
R914 B.n699 B.n66 585
R915 B.n66 B.n65 585
R916 B.n698 B.n697 585
R917 B.n697 B.n696 585
R918 B.n68 B.n67 585
R919 B.n695 B.n68 585
R920 B.n693 B.n692 585
R921 B.n694 B.n693 585
R922 B.n691 B.n73 585
R923 B.n73 B.n72 585
R924 B.n690 B.n689 585
R925 B.n689 B.n688 585
R926 B.n75 B.n74 585
R927 B.n687 B.n75 585
R928 B.n685 B.n684 585
R929 B.n686 B.n685 585
R930 B.n683 B.n80 585
R931 B.n80 B.n79 585
R932 B.n682 B.n681 585
R933 B.n681 B.n680 585
R934 B.n82 B.n81 585
R935 B.n679 B.n82 585
R936 B.n677 B.n676 585
R937 B.n678 B.n677 585
R938 B.n675 B.n87 585
R939 B.n87 B.n86 585
R940 B.n674 B.n673 585
R941 B.n673 B.n672 585
R942 B.n89 B.n88 585
R943 B.n671 B.n89 585
R944 B.n669 B.n668 585
R945 B.n670 B.n669 585
R946 B.n667 B.n94 585
R947 B.n94 B.n93 585
R948 B.n770 B.n769 585
R949 B.n768 B.n2 585
R950 B.n665 B.n94 506.916
R951 B.n661 B.n120 506.916
R952 B.n338 B.n311 506.916
R953 B.n438 B.n313 506.916
R954 B.n663 B.n662 256.663
R955 B.n663 B.n118 256.663
R956 B.n663 B.n117 256.663
R957 B.n663 B.n116 256.663
R958 B.n663 B.n115 256.663
R959 B.n663 B.n114 256.663
R960 B.n663 B.n113 256.663
R961 B.n663 B.n112 256.663
R962 B.n663 B.n111 256.663
R963 B.n663 B.n110 256.663
R964 B.n663 B.n109 256.663
R965 B.n663 B.n108 256.663
R966 B.n663 B.n107 256.663
R967 B.n663 B.n106 256.663
R968 B.n663 B.n105 256.663
R969 B.n663 B.n104 256.663
R970 B.n663 B.n103 256.663
R971 B.n663 B.n102 256.663
R972 B.n663 B.n101 256.663
R973 B.n663 B.n100 256.663
R974 B.n663 B.n99 256.663
R975 B.n663 B.n98 256.663
R976 B.n663 B.n97 256.663
R977 B.n664 B.n663 256.663
R978 B.n437 B.n436 256.663
R979 B.n436 B.n316 256.663
R980 B.n436 B.n317 256.663
R981 B.n436 B.n318 256.663
R982 B.n436 B.n319 256.663
R983 B.n436 B.n320 256.663
R984 B.n436 B.n321 256.663
R985 B.n436 B.n322 256.663
R986 B.n436 B.n323 256.663
R987 B.n436 B.n324 256.663
R988 B.n436 B.n325 256.663
R989 B.n436 B.n326 256.663
R990 B.n436 B.n327 256.663
R991 B.n436 B.n328 256.663
R992 B.n436 B.n329 256.663
R993 B.n436 B.n330 256.663
R994 B.n436 B.n331 256.663
R995 B.n436 B.n332 256.663
R996 B.n436 B.n333 256.663
R997 B.n436 B.n334 256.663
R998 B.n436 B.n335 256.663
R999 B.n436 B.n336 256.663
R1000 B.n436 B.n337 256.663
R1001 B.n772 B.n771 256.663
R1002 B.n123 B.t19 249.153
R1003 B.n121 B.t12 249.153
R1004 B.n343 B.t8 249.153
R1005 B.n340 B.t16 249.153
R1006 B.n121 B.t14 209.139
R1007 B.n343 B.t11 209.139
R1008 B.n123 B.t20 209.139
R1009 B.n340 B.t18 209.139
R1010 B.n125 B.n96 163.367
R1011 B.n129 B.n128 163.367
R1012 B.n133 B.n132 163.367
R1013 B.n137 B.n136 163.367
R1014 B.n141 B.n140 163.367
R1015 B.n145 B.n144 163.367
R1016 B.n149 B.n148 163.367
R1017 B.n153 B.n152 163.367
R1018 B.n157 B.n156 163.367
R1019 B.n162 B.n161 163.367
R1020 B.n166 B.n165 163.367
R1021 B.n170 B.n169 163.367
R1022 B.n174 B.n173 163.367
R1023 B.n178 B.n177 163.367
R1024 B.n183 B.n182 163.367
R1025 B.n187 B.n186 163.367
R1026 B.n191 B.n190 163.367
R1027 B.n195 B.n194 163.367
R1028 B.n199 B.n198 163.367
R1029 B.n203 B.n202 163.367
R1030 B.n207 B.n206 163.367
R1031 B.n211 B.n210 163.367
R1032 B.n213 B.n119 163.367
R1033 B.n444 B.n311 163.367
R1034 B.n444 B.n309 163.367
R1035 B.n448 B.n309 163.367
R1036 B.n448 B.n303 163.367
R1037 B.n456 B.n303 163.367
R1038 B.n456 B.n301 163.367
R1039 B.n460 B.n301 163.367
R1040 B.n460 B.n295 163.367
R1041 B.n468 B.n295 163.367
R1042 B.n468 B.n293 163.367
R1043 B.n472 B.n293 163.367
R1044 B.n472 B.n287 163.367
R1045 B.n480 B.n287 163.367
R1046 B.n480 B.n285 163.367
R1047 B.n484 B.n285 163.367
R1048 B.n484 B.n279 163.367
R1049 B.n492 B.n279 163.367
R1050 B.n492 B.n277 163.367
R1051 B.n496 B.n277 163.367
R1052 B.n496 B.n271 163.367
R1053 B.n504 B.n271 163.367
R1054 B.n504 B.n269 163.367
R1055 B.n508 B.n269 163.367
R1056 B.n508 B.n263 163.367
R1057 B.n516 B.n263 163.367
R1058 B.n516 B.n261 163.367
R1059 B.n520 B.n261 163.367
R1060 B.n520 B.n256 163.367
R1061 B.n529 B.n256 163.367
R1062 B.n529 B.n254 163.367
R1063 B.n533 B.n254 163.367
R1064 B.n533 B.n248 163.367
R1065 B.n541 B.n248 163.367
R1066 B.n541 B.n246 163.367
R1067 B.n545 B.n246 163.367
R1068 B.n545 B.n241 163.367
R1069 B.n554 B.n241 163.367
R1070 B.n554 B.n239 163.367
R1071 B.n558 B.n239 163.367
R1072 B.n558 B.n233 163.367
R1073 B.n566 B.n233 163.367
R1074 B.n566 B.n231 163.367
R1075 B.n570 B.n231 163.367
R1076 B.n570 B.n225 163.367
R1077 B.n578 B.n225 163.367
R1078 B.n578 B.n223 163.367
R1079 B.n583 B.n223 163.367
R1080 B.n583 B.n217 163.367
R1081 B.n591 B.n217 163.367
R1082 B.n592 B.n591 163.367
R1083 B.n592 B.n5 163.367
R1084 B.n6 B.n5 163.367
R1085 B.n7 B.n6 163.367
R1086 B.n598 B.n7 163.367
R1087 B.n599 B.n598 163.367
R1088 B.n599 B.n13 163.367
R1089 B.n14 B.n13 163.367
R1090 B.n15 B.n14 163.367
R1091 B.n604 B.n15 163.367
R1092 B.n604 B.n20 163.367
R1093 B.n21 B.n20 163.367
R1094 B.n22 B.n21 163.367
R1095 B.n609 B.n22 163.367
R1096 B.n609 B.n27 163.367
R1097 B.n28 B.n27 163.367
R1098 B.n29 B.n28 163.367
R1099 B.n614 B.n29 163.367
R1100 B.n614 B.n34 163.367
R1101 B.n35 B.n34 163.367
R1102 B.n36 B.n35 163.367
R1103 B.n619 B.n36 163.367
R1104 B.n619 B.n41 163.367
R1105 B.n42 B.n41 163.367
R1106 B.n43 B.n42 163.367
R1107 B.n624 B.n43 163.367
R1108 B.n624 B.n48 163.367
R1109 B.n49 B.n48 163.367
R1110 B.n50 B.n49 163.367
R1111 B.n629 B.n50 163.367
R1112 B.n629 B.n55 163.367
R1113 B.n56 B.n55 163.367
R1114 B.n57 B.n56 163.367
R1115 B.n634 B.n57 163.367
R1116 B.n634 B.n62 163.367
R1117 B.n63 B.n62 163.367
R1118 B.n64 B.n63 163.367
R1119 B.n639 B.n64 163.367
R1120 B.n639 B.n69 163.367
R1121 B.n70 B.n69 163.367
R1122 B.n71 B.n70 163.367
R1123 B.n644 B.n71 163.367
R1124 B.n644 B.n76 163.367
R1125 B.n77 B.n76 163.367
R1126 B.n78 B.n77 163.367
R1127 B.n649 B.n78 163.367
R1128 B.n649 B.n83 163.367
R1129 B.n84 B.n83 163.367
R1130 B.n85 B.n84 163.367
R1131 B.n654 B.n85 163.367
R1132 B.n654 B.n90 163.367
R1133 B.n91 B.n90 163.367
R1134 B.n92 B.n91 163.367
R1135 B.n120 B.n92 163.367
R1136 B.n435 B.n315 163.367
R1137 B.n435 B.n339 163.367
R1138 B.n431 B.n430 163.367
R1139 B.n427 B.n426 163.367
R1140 B.n423 B.n422 163.367
R1141 B.n419 B.n418 163.367
R1142 B.n415 B.n414 163.367
R1143 B.n411 B.n410 163.367
R1144 B.n407 B.n406 163.367
R1145 B.n403 B.n402 163.367
R1146 B.n399 B.n398 163.367
R1147 B.n395 B.n394 163.367
R1148 B.n391 B.n390 163.367
R1149 B.n387 B.n386 163.367
R1150 B.n383 B.n382 163.367
R1151 B.n379 B.n378 163.367
R1152 B.n375 B.n374 163.367
R1153 B.n371 B.n370 163.367
R1154 B.n367 B.n366 163.367
R1155 B.n363 B.n362 163.367
R1156 B.n359 B.n358 163.367
R1157 B.n355 B.n354 163.367
R1158 B.n351 B.n350 163.367
R1159 B.n347 B.n338 163.367
R1160 B.n442 B.n313 163.367
R1161 B.n442 B.n307 163.367
R1162 B.n450 B.n307 163.367
R1163 B.n450 B.n305 163.367
R1164 B.n454 B.n305 163.367
R1165 B.n454 B.n299 163.367
R1166 B.n462 B.n299 163.367
R1167 B.n462 B.n297 163.367
R1168 B.n466 B.n297 163.367
R1169 B.n466 B.n291 163.367
R1170 B.n474 B.n291 163.367
R1171 B.n474 B.n289 163.367
R1172 B.n478 B.n289 163.367
R1173 B.n478 B.n283 163.367
R1174 B.n486 B.n283 163.367
R1175 B.n486 B.n281 163.367
R1176 B.n490 B.n281 163.367
R1177 B.n490 B.n275 163.367
R1178 B.n498 B.n275 163.367
R1179 B.n498 B.n273 163.367
R1180 B.n502 B.n273 163.367
R1181 B.n502 B.n267 163.367
R1182 B.n510 B.n267 163.367
R1183 B.n510 B.n265 163.367
R1184 B.n514 B.n265 163.367
R1185 B.n514 B.n259 163.367
R1186 B.n523 B.n259 163.367
R1187 B.n523 B.n257 163.367
R1188 B.n527 B.n257 163.367
R1189 B.n527 B.n252 163.367
R1190 B.n535 B.n252 163.367
R1191 B.n535 B.n250 163.367
R1192 B.n539 B.n250 163.367
R1193 B.n539 B.n244 163.367
R1194 B.n548 B.n244 163.367
R1195 B.n548 B.n242 163.367
R1196 B.n552 B.n242 163.367
R1197 B.n552 B.n237 163.367
R1198 B.n560 B.n237 163.367
R1199 B.n560 B.n235 163.367
R1200 B.n564 B.n235 163.367
R1201 B.n564 B.n229 163.367
R1202 B.n572 B.n229 163.367
R1203 B.n572 B.n227 163.367
R1204 B.n576 B.n227 163.367
R1205 B.n576 B.n221 163.367
R1206 B.n585 B.n221 163.367
R1207 B.n585 B.n219 163.367
R1208 B.n589 B.n219 163.367
R1209 B.n589 B.n3 163.367
R1210 B.n770 B.n3 163.367
R1211 B.n766 B.n2 163.367
R1212 B.n766 B.n765 163.367
R1213 B.n765 B.n9 163.367
R1214 B.n761 B.n9 163.367
R1215 B.n761 B.n11 163.367
R1216 B.n757 B.n11 163.367
R1217 B.n757 B.n17 163.367
R1218 B.n753 B.n17 163.367
R1219 B.n753 B.n19 163.367
R1220 B.n749 B.n19 163.367
R1221 B.n749 B.n24 163.367
R1222 B.n745 B.n24 163.367
R1223 B.n745 B.n26 163.367
R1224 B.n741 B.n26 163.367
R1225 B.n741 B.n30 163.367
R1226 B.n737 B.n30 163.367
R1227 B.n737 B.n32 163.367
R1228 B.n733 B.n32 163.367
R1229 B.n733 B.n38 163.367
R1230 B.n729 B.n38 163.367
R1231 B.n729 B.n40 163.367
R1232 B.n725 B.n40 163.367
R1233 B.n725 B.n44 163.367
R1234 B.n721 B.n44 163.367
R1235 B.n721 B.n46 163.367
R1236 B.n717 B.n46 163.367
R1237 B.n717 B.n52 163.367
R1238 B.n713 B.n52 163.367
R1239 B.n713 B.n54 163.367
R1240 B.n709 B.n54 163.367
R1241 B.n709 B.n59 163.367
R1242 B.n705 B.n59 163.367
R1243 B.n705 B.n61 163.367
R1244 B.n701 B.n61 163.367
R1245 B.n701 B.n66 163.367
R1246 B.n697 B.n66 163.367
R1247 B.n697 B.n68 163.367
R1248 B.n693 B.n68 163.367
R1249 B.n693 B.n73 163.367
R1250 B.n689 B.n73 163.367
R1251 B.n689 B.n75 163.367
R1252 B.n685 B.n75 163.367
R1253 B.n685 B.n80 163.367
R1254 B.n681 B.n80 163.367
R1255 B.n681 B.n82 163.367
R1256 B.n677 B.n82 163.367
R1257 B.n677 B.n87 163.367
R1258 B.n673 B.n87 163.367
R1259 B.n673 B.n89 163.367
R1260 B.n669 B.n89 163.367
R1261 B.n669 B.n94 163.367
R1262 B.n122 B.t15 152.121
R1263 B.n344 B.t10 152.121
R1264 B.n124 B.t21 152.121
R1265 B.n341 B.t17 152.121
R1266 B.n436 B.n312 127.816
R1267 B.n663 B.n93 127.816
R1268 B.n443 B.n312 76.9157
R1269 B.n443 B.n308 76.9157
R1270 B.n449 B.n308 76.9157
R1271 B.n449 B.n304 76.9157
R1272 B.n455 B.n304 76.9157
R1273 B.n455 B.n300 76.9157
R1274 B.n461 B.n300 76.9157
R1275 B.n467 B.n296 76.9157
R1276 B.n467 B.n292 76.9157
R1277 B.n473 B.n292 76.9157
R1278 B.n473 B.n288 76.9157
R1279 B.n479 B.n288 76.9157
R1280 B.n479 B.n284 76.9157
R1281 B.n485 B.n284 76.9157
R1282 B.n485 B.n280 76.9157
R1283 B.n491 B.n280 76.9157
R1284 B.n491 B.n276 76.9157
R1285 B.n497 B.n276 76.9157
R1286 B.n503 B.n272 76.9157
R1287 B.n503 B.n268 76.9157
R1288 B.n509 B.n268 76.9157
R1289 B.n509 B.n264 76.9157
R1290 B.n515 B.n264 76.9157
R1291 B.n515 B.n260 76.9157
R1292 B.n522 B.n260 76.9157
R1293 B.n522 B.n521 76.9157
R1294 B.n528 B.n253 76.9157
R1295 B.n534 B.n253 76.9157
R1296 B.n534 B.n249 76.9157
R1297 B.n540 B.n249 76.9157
R1298 B.n540 B.n245 76.9157
R1299 B.n547 B.n245 76.9157
R1300 B.n547 B.n546 76.9157
R1301 B.n553 B.n238 76.9157
R1302 B.n559 B.n238 76.9157
R1303 B.n559 B.n234 76.9157
R1304 B.n565 B.n234 76.9157
R1305 B.n565 B.n230 76.9157
R1306 B.n571 B.n230 76.9157
R1307 B.n571 B.n226 76.9157
R1308 B.n577 B.n226 76.9157
R1309 B.n584 B.n222 76.9157
R1310 B.n584 B.n218 76.9157
R1311 B.n590 B.n218 76.9157
R1312 B.n590 B.n4 76.9157
R1313 B.n769 B.n4 76.9157
R1314 B.n769 B.n768 76.9157
R1315 B.n768 B.n767 76.9157
R1316 B.n767 B.n8 76.9157
R1317 B.n12 B.n8 76.9157
R1318 B.n760 B.n12 76.9157
R1319 B.n760 B.n759 76.9157
R1320 B.n758 B.n16 76.9157
R1321 B.n752 B.n16 76.9157
R1322 B.n752 B.n751 76.9157
R1323 B.n751 B.n750 76.9157
R1324 B.n750 B.n23 76.9157
R1325 B.n744 B.n23 76.9157
R1326 B.n744 B.n743 76.9157
R1327 B.n743 B.n742 76.9157
R1328 B.n736 B.n33 76.9157
R1329 B.n736 B.n735 76.9157
R1330 B.n735 B.n734 76.9157
R1331 B.n734 B.n37 76.9157
R1332 B.n728 B.n37 76.9157
R1333 B.n728 B.n727 76.9157
R1334 B.n727 B.n726 76.9157
R1335 B.n720 B.n47 76.9157
R1336 B.n720 B.n719 76.9157
R1337 B.n719 B.n718 76.9157
R1338 B.n718 B.n51 76.9157
R1339 B.n712 B.n51 76.9157
R1340 B.n712 B.n711 76.9157
R1341 B.n711 B.n710 76.9157
R1342 B.n710 B.n58 76.9157
R1343 B.n704 B.n703 76.9157
R1344 B.n703 B.n702 76.9157
R1345 B.n702 B.n65 76.9157
R1346 B.n696 B.n65 76.9157
R1347 B.n696 B.n695 76.9157
R1348 B.n695 B.n694 76.9157
R1349 B.n694 B.n72 76.9157
R1350 B.n688 B.n72 76.9157
R1351 B.n688 B.n687 76.9157
R1352 B.n687 B.n686 76.9157
R1353 B.n686 B.n79 76.9157
R1354 B.n680 B.n679 76.9157
R1355 B.n679 B.n678 76.9157
R1356 B.n678 B.n86 76.9157
R1357 B.n672 B.n86 76.9157
R1358 B.n672 B.n671 76.9157
R1359 B.n671 B.n670 76.9157
R1360 B.n670 B.n93 76.9157
R1361 B.n665 B.n664 71.676
R1362 B.n125 B.n97 71.676
R1363 B.n129 B.n98 71.676
R1364 B.n133 B.n99 71.676
R1365 B.n137 B.n100 71.676
R1366 B.n141 B.n101 71.676
R1367 B.n145 B.n102 71.676
R1368 B.n149 B.n103 71.676
R1369 B.n153 B.n104 71.676
R1370 B.n157 B.n105 71.676
R1371 B.n162 B.n106 71.676
R1372 B.n166 B.n107 71.676
R1373 B.n170 B.n108 71.676
R1374 B.n174 B.n109 71.676
R1375 B.n178 B.n110 71.676
R1376 B.n183 B.n111 71.676
R1377 B.n187 B.n112 71.676
R1378 B.n191 B.n113 71.676
R1379 B.n195 B.n114 71.676
R1380 B.n199 B.n115 71.676
R1381 B.n203 B.n116 71.676
R1382 B.n207 B.n117 71.676
R1383 B.n211 B.n118 71.676
R1384 B.n662 B.n119 71.676
R1385 B.n662 B.n661 71.676
R1386 B.n213 B.n118 71.676
R1387 B.n210 B.n117 71.676
R1388 B.n206 B.n116 71.676
R1389 B.n202 B.n115 71.676
R1390 B.n198 B.n114 71.676
R1391 B.n194 B.n113 71.676
R1392 B.n190 B.n112 71.676
R1393 B.n186 B.n111 71.676
R1394 B.n182 B.n110 71.676
R1395 B.n177 B.n109 71.676
R1396 B.n173 B.n108 71.676
R1397 B.n169 B.n107 71.676
R1398 B.n165 B.n106 71.676
R1399 B.n161 B.n105 71.676
R1400 B.n156 B.n104 71.676
R1401 B.n152 B.n103 71.676
R1402 B.n148 B.n102 71.676
R1403 B.n144 B.n101 71.676
R1404 B.n140 B.n100 71.676
R1405 B.n136 B.n99 71.676
R1406 B.n132 B.n98 71.676
R1407 B.n128 B.n97 71.676
R1408 B.n664 B.n96 71.676
R1409 B.n438 B.n437 71.676
R1410 B.n339 B.n316 71.676
R1411 B.n430 B.n317 71.676
R1412 B.n426 B.n318 71.676
R1413 B.n422 B.n319 71.676
R1414 B.n418 B.n320 71.676
R1415 B.n414 B.n321 71.676
R1416 B.n410 B.n322 71.676
R1417 B.n406 B.n323 71.676
R1418 B.n402 B.n324 71.676
R1419 B.n398 B.n325 71.676
R1420 B.n394 B.n326 71.676
R1421 B.n390 B.n327 71.676
R1422 B.n386 B.n328 71.676
R1423 B.n382 B.n329 71.676
R1424 B.n378 B.n330 71.676
R1425 B.n374 B.n331 71.676
R1426 B.n370 B.n332 71.676
R1427 B.n366 B.n333 71.676
R1428 B.n362 B.n334 71.676
R1429 B.n358 B.n335 71.676
R1430 B.n354 B.n336 71.676
R1431 B.n350 B.n337 71.676
R1432 B.n437 B.n315 71.676
R1433 B.n431 B.n316 71.676
R1434 B.n427 B.n317 71.676
R1435 B.n423 B.n318 71.676
R1436 B.n419 B.n319 71.676
R1437 B.n415 B.n320 71.676
R1438 B.n411 B.n321 71.676
R1439 B.n407 B.n322 71.676
R1440 B.n403 B.n323 71.676
R1441 B.n399 B.n324 71.676
R1442 B.n395 B.n325 71.676
R1443 B.n391 B.n326 71.676
R1444 B.n387 B.n327 71.676
R1445 B.n383 B.n328 71.676
R1446 B.n379 B.n329 71.676
R1447 B.n375 B.n330 71.676
R1448 B.n371 B.n331 71.676
R1449 B.n367 B.n332 71.676
R1450 B.n363 B.n333 71.676
R1451 B.n359 B.n334 71.676
R1452 B.n355 B.n335 71.676
R1453 B.n351 B.n336 71.676
R1454 B.n347 B.n337 71.676
R1455 B.n771 B.n770 71.676
R1456 B.n771 B.n2 71.676
R1457 B.n546 B.t4 71.2601
R1458 B.n33 B.t3 71.2601
R1459 B.n461 B.t9 59.9491
R1460 B.n680 B.t13 59.9491
R1461 B.n159 B.n124 59.5399
R1462 B.n180 B.n122 59.5399
R1463 B.n345 B.n344 59.5399
R1464 B.n342 B.n341 59.5399
R1465 B.n124 B.n123 57.0187
R1466 B.n122 B.n121 57.0187
R1467 B.n344 B.n343 57.0187
R1468 B.n341 B.n340 57.0187
R1469 B.n528 B.t0 55.4247
R1470 B.n726 B.t5 55.4247
R1471 B.n497 B.t7 48.638
R1472 B.n704 B.t6 48.638
R1473 B.n577 B.t2 44.1136
R1474 B.t1 B.n758 44.1136
R1475 B.n440 B.n439 32.9371
R1476 B.n346 B.n310 32.9371
R1477 B.n660 B.n659 32.9371
R1478 B.n667 B.n666 32.9371
R1479 B.t2 B.n222 32.8026
R1480 B.n759 B.t1 32.8026
R1481 B.t7 B.n272 28.2781
R1482 B.t6 B.n58 28.2781
R1483 B.n521 B.t0 21.4915
R1484 B.n47 B.t5 21.4915
R1485 B B.n772 18.0485
R1486 B.t9 B.n296 16.9671
R1487 B.t13 B.n79 16.9671
R1488 B.n441 B.n440 10.6151
R1489 B.n441 B.n306 10.6151
R1490 B.n451 B.n306 10.6151
R1491 B.n452 B.n451 10.6151
R1492 B.n453 B.n452 10.6151
R1493 B.n453 B.n298 10.6151
R1494 B.n463 B.n298 10.6151
R1495 B.n464 B.n463 10.6151
R1496 B.n465 B.n464 10.6151
R1497 B.n465 B.n290 10.6151
R1498 B.n475 B.n290 10.6151
R1499 B.n476 B.n475 10.6151
R1500 B.n477 B.n476 10.6151
R1501 B.n477 B.n282 10.6151
R1502 B.n487 B.n282 10.6151
R1503 B.n488 B.n487 10.6151
R1504 B.n489 B.n488 10.6151
R1505 B.n489 B.n274 10.6151
R1506 B.n499 B.n274 10.6151
R1507 B.n500 B.n499 10.6151
R1508 B.n501 B.n500 10.6151
R1509 B.n501 B.n266 10.6151
R1510 B.n511 B.n266 10.6151
R1511 B.n512 B.n511 10.6151
R1512 B.n513 B.n512 10.6151
R1513 B.n513 B.n258 10.6151
R1514 B.n524 B.n258 10.6151
R1515 B.n525 B.n524 10.6151
R1516 B.n526 B.n525 10.6151
R1517 B.n526 B.n251 10.6151
R1518 B.n536 B.n251 10.6151
R1519 B.n537 B.n536 10.6151
R1520 B.n538 B.n537 10.6151
R1521 B.n538 B.n243 10.6151
R1522 B.n549 B.n243 10.6151
R1523 B.n550 B.n549 10.6151
R1524 B.n551 B.n550 10.6151
R1525 B.n551 B.n236 10.6151
R1526 B.n561 B.n236 10.6151
R1527 B.n562 B.n561 10.6151
R1528 B.n563 B.n562 10.6151
R1529 B.n563 B.n228 10.6151
R1530 B.n573 B.n228 10.6151
R1531 B.n574 B.n573 10.6151
R1532 B.n575 B.n574 10.6151
R1533 B.n575 B.n220 10.6151
R1534 B.n586 B.n220 10.6151
R1535 B.n587 B.n586 10.6151
R1536 B.n588 B.n587 10.6151
R1537 B.n588 B.n0 10.6151
R1538 B.n439 B.n314 10.6151
R1539 B.n434 B.n314 10.6151
R1540 B.n434 B.n433 10.6151
R1541 B.n433 B.n432 10.6151
R1542 B.n432 B.n429 10.6151
R1543 B.n429 B.n428 10.6151
R1544 B.n428 B.n425 10.6151
R1545 B.n425 B.n424 10.6151
R1546 B.n424 B.n421 10.6151
R1547 B.n421 B.n420 10.6151
R1548 B.n420 B.n417 10.6151
R1549 B.n417 B.n416 10.6151
R1550 B.n416 B.n413 10.6151
R1551 B.n413 B.n412 10.6151
R1552 B.n412 B.n409 10.6151
R1553 B.n409 B.n408 10.6151
R1554 B.n408 B.n405 10.6151
R1555 B.n405 B.n404 10.6151
R1556 B.n401 B.n400 10.6151
R1557 B.n400 B.n397 10.6151
R1558 B.n397 B.n396 10.6151
R1559 B.n396 B.n393 10.6151
R1560 B.n393 B.n392 10.6151
R1561 B.n392 B.n389 10.6151
R1562 B.n389 B.n388 10.6151
R1563 B.n388 B.n385 10.6151
R1564 B.n385 B.n384 10.6151
R1565 B.n381 B.n380 10.6151
R1566 B.n380 B.n377 10.6151
R1567 B.n377 B.n376 10.6151
R1568 B.n376 B.n373 10.6151
R1569 B.n373 B.n372 10.6151
R1570 B.n372 B.n369 10.6151
R1571 B.n369 B.n368 10.6151
R1572 B.n368 B.n365 10.6151
R1573 B.n365 B.n364 10.6151
R1574 B.n364 B.n361 10.6151
R1575 B.n361 B.n360 10.6151
R1576 B.n360 B.n357 10.6151
R1577 B.n357 B.n356 10.6151
R1578 B.n356 B.n353 10.6151
R1579 B.n353 B.n352 10.6151
R1580 B.n352 B.n349 10.6151
R1581 B.n349 B.n348 10.6151
R1582 B.n348 B.n346 10.6151
R1583 B.n445 B.n310 10.6151
R1584 B.n446 B.n445 10.6151
R1585 B.n447 B.n446 10.6151
R1586 B.n447 B.n302 10.6151
R1587 B.n457 B.n302 10.6151
R1588 B.n458 B.n457 10.6151
R1589 B.n459 B.n458 10.6151
R1590 B.n459 B.n294 10.6151
R1591 B.n469 B.n294 10.6151
R1592 B.n470 B.n469 10.6151
R1593 B.n471 B.n470 10.6151
R1594 B.n471 B.n286 10.6151
R1595 B.n481 B.n286 10.6151
R1596 B.n482 B.n481 10.6151
R1597 B.n483 B.n482 10.6151
R1598 B.n483 B.n278 10.6151
R1599 B.n493 B.n278 10.6151
R1600 B.n494 B.n493 10.6151
R1601 B.n495 B.n494 10.6151
R1602 B.n495 B.n270 10.6151
R1603 B.n505 B.n270 10.6151
R1604 B.n506 B.n505 10.6151
R1605 B.n507 B.n506 10.6151
R1606 B.n507 B.n262 10.6151
R1607 B.n517 B.n262 10.6151
R1608 B.n518 B.n517 10.6151
R1609 B.n519 B.n518 10.6151
R1610 B.n519 B.n255 10.6151
R1611 B.n530 B.n255 10.6151
R1612 B.n531 B.n530 10.6151
R1613 B.n532 B.n531 10.6151
R1614 B.n532 B.n247 10.6151
R1615 B.n542 B.n247 10.6151
R1616 B.n543 B.n542 10.6151
R1617 B.n544 B.n543 10.6151
R1618 B.n544 B.n240 10.6151
R1619 B.n555 B.n240 10.6151
R1620 B.n556 B.n555 10.6151
R1621 B.n557 B.n556 10.6151
R1622 B.n557 B.n232 10.6151
R1623 B.n567 B.n232 10.6151
R1624 B.n568 B.n567 10.6151
R1625 B.n569 B.n568 10.6151
R1626 B.n569 B.n224 10.6151
R1627 B.n579 B.n224 10.6151
R1628 B.n580 B.n579 10.6151
R1629 B.n582 B.n580 10.6151
R1630 B.n582 B.n581 10.6151
R1631 B.n581 B.n216 10.6151
R1632 B.n593 B.n216 10.6151
R1633 B.n594 B.n593 10.6151
R1634 B.n595 B.n594 10.6151
R1635 B.n596 B.n595 10.6151
R1636 B.n597 B.n596 10.6151
R1637 B.n600 B.n597 10.6151
R1638 B.n601 B.n600 10.6151
R1639 B.n602 B.n601 10.6151
R1640 B.n603 B.n602 10.6151
R1641 B.n605 B.n603 10.6151
R1642 B.n606 B.n605 10.6151
R1643 B.n607 B.n606 10.6151
R1644 B.n608 B.n607 10.6151
R1645 B.n610 B.n608 10.6151
R1646 B.n611 B.n610 10.6151
R1647 B.n612 B.n611 10.6151
R1648 B.n613 B.n612 10.6151
R1649 B.n615 B.n613 10.6151
R1650 B.n616 B.n615 10.6151
R1651 B.n617 B.n616 10.6151
R1652 B.n618 B.n617 10.6151
R1653 B.n620 B.n618 10.6151
R1654 B.n621 B.n620 10.6151
R1655 B.n622 B.n621 10.6151
R1656 B.n623 B.n622 10.6151
R1657 B.n625 B.n623 10.6151
R1658 B.n626 B.n625 10.6151
R1659 B.n627 B.n626 10.6151
R1660 B.n628 B.n627 10.6151
R1661 B.n630 B.n628 10.6151
R1662 B.n631 B.n630 10.6151
R1663 B.n632 B.n631 10.6151
R1664 B.n633 B.n632 10.6151
R1665 B.n635 B.n633 10.6151
R1666 B.n636 B.n635 10.6151
R1667 B.n637 B.n636 10.6151
R1668 B.n638 B.n637 10.6151
R1669 B.n640 B.n638 10.6151
R1670 B.n641 B.n640 10.6151
R1671 B.n642 B.n641 10.6151
R1672 B.n643 B.n642 10.6151
R1673 B.n645 B.n643 10.6151
R1674 B.n646 B.n645 10.6151
R1675 B.n647 B.n646 10.6151
R1676 B.n648 B.n647 10.6151
R1677 B.n650 B.n648 10.6151
R1678 B.n651 B.n650 10.6151
R1679 B.n652 B.n651 10.6151
R1680 B.n653 B.n652 10.6151
R1681 B.n655 B.n653 10.6151
R1682 B.n656 B.n655 10.6151
R1683 B.n657 B.n656 10.6151
R1684 B.n658 B.n657 10.6151
R1685 B.n659 B.n658 10.6151
R1686 B.n764 B.n1 10.6151
R1687 B.n764 B.n763 10.6151
R1688 B.n763 B.n762 10.6151
R1689 B.n762 B.n10 10.6151
R1690 B.n756 B.n10 10.6151
R1691 B.n756 B.n755 10.6151
R1692 B.n755 B.n754 10.6151
R1693 B.n754 B.n18 10.6151
R1694 B.n748 B.n18 10.6151
R1695 B.n748 B.n747 10.6151
R1696 B.n747 B.n746 10.6151
R1697 B.n746 B.n25 10.6151
R1698 B.n740 B.n25 10.6151
R1699 B.n740 B.n739 10.6151
R1700 B.n739 B.n738 10.6151
R1701 B.n738 B.n31 10.6151
R1702 B.n732 B.n31 10.6151
R1703 B.n732 B.n731 10.6151
R1704 B.n731 B.n730 10.6151
R1705 B.n730 B.n39 10.6151
R1706 B.n724 B.n39 10.6151
R1707 B.n724 B.n723 10.6151
R1708 B.n723 B.n722 10.6151
R1709 B.n722 B.n45 10.6151
R1710 B.n716 B.n45 10.6151
R1711 B.n716 B.n715 10.6151
R1712 B.n715 B.n714 10.6151
R1713 B.n714 B.n53 10.6151
R1714 B.n708 B.n53 10.6151
R1715 B.n708 B.n707 10.6151
R1716 B.n707 B.n706 10.6151
R1717 B.n706 B.n60 10.6151
R1718 B.n700 B.n60 10.6151
R1719 B.n700 B.n699 10.6151
R1720 B.n699 B.n698 10.6151
R1721 B.n698 B.n67 10.6151
R1722 B.n692 B.n67 10.6151
R1723 B.n692 B.n691 10.6151
R1724 B.n691 B.n690 10.6151
R1725 B.n690 B.n74 10.6151
R1726 B.n684 B.n74 10.6151
R1727 B.n684 B.n683 10.6151
R1728 B.n683 B.n682 10.6151
R1729 B.n682 B.n81 10.6151
R1730 B.n676 B.n81 10.6151
R1731 B.n676 B.n675 10.6151
R1732 B.n675 B.n674 10.6151
R1733 B.n674 B.n88 10.6151
R1734 B.n668 B.n88 10.6151
R1735 B.n668 B.n667 10.6151
R1736 B.n666 B.n95 10.6151
R1737 B.n126 B.n95 10.6151
R1738 B.n127 B.n126 10.6151
R1739 B.n130 B.n127 10.6151
R1740 B.n131 B.n130 10.6151
R1741 B.n134 B.n131 10.6151
R1742 B.n135 B.n134 10.6151
R1743 B.n138 B.n135 10.6151
R1744 B.n139 B.n138 10.6151
R1745 B.n142 B.n139 10.6151
R1746 B.n143 B.n142 10.6151
R1747 B.n146 B.n143 10.6151
R1748 B.n147 B.n146 10.6151
R1749 B.n150 B.n147 10.6151
R1750 B.n151 B.n150 10.6151
R1751 B.n154 B.n151 10.6151
R1752 B.n155 B.n154 10.6151
R1753 B.n158 B.n155 10.6151
R1754 B.n163 B.n160 10.6151
R1755 B.n164 B.n163 10.6151
R1756 B.n167 B.n164 10.6151
R1757 B.n168 B.n167 10.6151
R1758 B.n171 B.n168 10.6151
R1759 B.n172 B.n171 10.6151
R1760 B.n175 B.n172 10.6151
R1761 B.n176 B.n175 10.6151
R1762 B.n179 B.n176 10.6151
R1763 B.n184 B.n181 10.6151
R1764 B.n185 B.n184 10.6151
R1765 B.n188 B.n185 10.6151
R1766 B.n189 B.n188 10.6151
R1767 B.n192 B.n189 10.6151
R1768 B.n193 B.n192 10.6151
R1769 B.n196 B.n193 10.6151
R1770 B.n197 B.n196 10.6151
R1771 B.n200 B.n197 10.6151
R1772 B.n201 B.n200 10.6151
R1773 B.n204 B.n201 10.6151
R1774 B.n205 B.n204 10.6151
R1775 B.n208 B.n205 10.6151
R1776 B.n209 B.n208 10.6151
R1777 B.n212 B.n209 10.6151
R1778 B.n214 B.n212 10.6151
R1779 B.n215 B.n214 10.6151
R1780 B.n660 B.n215 10.6151
R1781 B.n404 B.n342 9.36635
R1782 B.n381 B.n345 9.36635
R1783 B.n159 B.n158 9.36635
R1784 B.n181 B.n180 9.36635
R1785 B.n772 B.n0 8.11757
R1786 B.n772 B.n1 8.11757
R1787 B.n553 B.t4 5.65603
R1788 B.n742 B.t3 5.65603
R1789 B.n401 B.n342 1.24928
R1790 B.n384 B.n345 1.24928
R1791 B.n160 B.n159 1.24928
R1792 B.n180 B.n179 1.24928
R1793 VN.n55 VN.n29 161.3
R1794 VN.n54 VN.n53 161.3
R1795 VN.n52 VN.n30 161.3
R1796 VN.n51 VN.n50 161.3
R1797 VN.n49 VN.n31 161.3
R1798 VN.n48 VN.n47 161.3
R1799 VN.n46 VN.n45 161.3
R1800 VN.n44 VN.n33 161.3
R1801 VN.n43 VN.n42 161.3
R1802 VN.n41 VN.n34 161.3
R1803 VN.n40 VN.n39 161.3
R1804 VN.n38 VN.n35 161.3
R1805 VN.n26 VN.n0 161.3
R1806 VN.n25 VN.n24 161.3
R1807 VN.n23 VN.n1 161.3
R1808 VN.n22 VN.n21 161.3
R1809 VN.n20 VN.n2 161.3
R1810 VN.n19 VN.n18 161.3
R1811 VN.n17 VN.n16 161.3
R1812 VN.n15 VN.n4 161.3
R1813 VN.n14 VN.n13 161.3
R1814 VN.n12 VN.n5 161.3
R1815 VN.n11 VN.n10 161.3
R1816 VN.n9 VN.n6 161.3
R1817 VN.n28 VN.n27 102.927
R1818 VN.n57 VN.n56 102.927
R1819 VN.n7 VN.t3 74.0585
R1820 VN.n36 VN.t4 74.0585
R1821 VN.n8 VN.n7 61.551
R1822 VN.n37 VN.n36 61.551
R1823 VN.n14 VN.n5 56.5193
R1824 VN.n21 VN.n1 56.5193
R1825 VN.n43 VN.n34 56.5193
R1826 VN.n50 VN.n30 56.5193
R1827 VN VN.n57 45.4906
R1828 VN.n8 VN.t6 41.0905
R1829 VN.n3 VN.t1 41.0905
R1830 VN.n27 VN.t2 41.0905
R1831 VN.n37 VN.t5 41.0905
R1832 VN.n32 VN.t7 41.0905
R1833 VN.n56 VN.t0 41.0905
R1834 VN.n10 VN.n9 24.4675
R1835 VN.n10 VN.n5 24.4675
R1836 VN.n15 VN.n14 24.4675
R1837 VN.n16 VN.n15 24.4675
R1838 VN.n20 VN.n19 24.4675
R1839 VN.n21 VN.n20 24.4675
R1840 VN.n25 VN.n1 24.4675
R1841 VN.n26 VN.n25 24.4675
R1842 VN.n39 VN.n34 24.4675
R1843 VN.n39 VN.n38 24.4675
R1844 VN.n50 VN.n49 24.4675
R1845 VN.n49 VN.n48 24.4675
R1846 VN.n45 VN.n44 24.4675
R1847 VN.n44 VN.n43 24.4675
R1848 VN.n55 VN.n54 24.4675
R1849 VN.n54 VN.n30 24.4675
R1850 VN.n19 VN.n3 13.702
R1851 VN.n48 VN.n32 13.702
R1852 VN.n9 VN.n8 10.766
R1853 VN.n16 VN.n3 10.766
R1854 VN.n38 VN.n37 10.766
R1855 VN.n45 VN.n32 10.766
R1856 VN.n27 VN.n26 7.82994
R1857 VN.n56 VN.n55 7.82994
R1858 VN.n36 VN.n35 6.98649
R1859 VN.n7 VN.n6 6.98649
R1860 VN.n57 VN.n29 0.278367
R1861 VN.n28 VN.n0 0.278367
R1862 VN.n53 VN.n29 0.189894
R1863 VN.n53 VN.n52 0.189894
R1864 VN.n52 VN.n51 0.189894
R1865 VN.n51 VN.n31 0.189894
R1866 VN.n47 VN.n31 0.189894
R1867 VN.n47 VN.n46 0.189894
R1868 VN.n46 VN.n33 0.189894
R1869 VN.n42 VN.n33 0.189894
R1870 VN.n42 VN.n41 0.189894
R1871 VN.n41 VN.n40 0.189894
R1872 VN.n40 VN.n35 0.189894
R1873 VN.n11 VN.n6 0.189894
R1874 VN.n12 VN.n11 0.189894
R1875 VN.n13 VN.n12 0.189894
R1876 VN.n13 VN.n4 0.189894
R1877 VN.n17 VN.n4 0.189894
R1878 VN.n18 VN.n17 0.189894
R1879 VN.n18 VN.n2 0.189894
R1880 VN.n22 VN.n2 0.189894
R1881 VN.n23 VN.n22 0.189894
R1882 VN.n24 VN.n23 0.189894
R1883 VN.n24 VN.n0 0.189894
R1884 VN VN.n28 0.153454
R1885 VDD2.n2 VDD2.n1 69.7202
R1886 VDD2.n2 VDD2.n0 69.7202
R1887 VDD2 VDD2.n5 69.7174
R1888 VDD2.n4 VDD2.n3 68.5085
R1889 VDD2.n4 VDD2.n2 38.9567
R1890 VDD2.n5 VDD2.t2 4.44994
R1891 VDD2.n5 VDD2.t3 4.44994
R1892 VDD2.n3 VDD2.t7 4.44994
R1893 VDD2.n3 VDD2.t0 4.44994
R1894 VDD2.n1 VDD2.t6 4.44994
R1895 VDD2.n1 VDD2.t5 4.44994
R1896 VDD2.n0 VDD2.t4 4.44994
R1897 VDD2.n0 VDD2.t1 4.44994
R1898 VDD2 VDD2.n4 1.32593
C0 VTAIL VN 4.44046f
C1 VDD2 VP 0.52542f
C2 VDD1 VP 3.87483f
C3 VDD2 VN 3.50736f
C4 VDD1 VN 0.155905f
C5 VDD2 VTAIL 5.59987f
C6 VDD1 VTAIL 5.54539f
C7 VDD2 VDD1 1.78332f
C8 VN VP 6.2821f
C9 VTAIL VP 4.45456f
C10 VDD2 B 4.75422f
C11 VDD1 B 5.199451f
C12 VTAIL B 5.586819f
C13 VN B 14.78732f
C14 VP B 13.383692f
C15 VDD2.t4 B 0.085012f
C16 VDD2.t1 B 0.085012f
C17 VDD2.n0 B 0.688952f
C18 VDD2.t6 B 0.085012f
C19 VDD2.t5 B 0.085012f
C20 VDD2.n1 B 0.688952f
C21 VDD2.n2 B 2.71127f
C22 VDD2.t7 B 0.085012f
C23 VDD2.t0 B 0.085012f
C24 VDD2.n3 B 0.680403f
C25 VDD2.n4 B 2.28112f
C26 VDD2.t2 B 0.085012f
C27 VDD2.t3 B 0.085012f
C28 VDD2.n5 B 0.688921f
C29 VN.n0 B 0.034342f
C30 VN.t2 B 0.784334f
C31 VN.n1 B 0.042381f
C32 VN.n2 B 0.026048f
C33 VN.t1 B 0.784334f
C34 VN.n3 B 0.306582f
C35 VN.n4 B 0.026048f
C36 VN.n5 B 0.038025f
C37 VN.n6 B 0.251994f
C38 VN.t6 B 0.784334f
C39 VN.t3 B 0.992437f
C40 VN.n7 B 0.367459f
C41 VN.n8 B 0.380376f
C42 VN.n9 B 0.035125f
C43 VN.n10 B 0.048547f
C44 VN.n11 B 0.026048f
C45 VN.n12 B 0.026048f
C46 VN.n13 B 0.026048f
C47 VN.n14 B 0.038025f
C48 VN.n15 B 0.048547f
C49 VN.n16 B 0.035125f
C50 VN.n17 B 0.026048f
C51 VN.n18 B 0.026048f
C52 VN.n19 B 0.038001f
C53 VN.n20 B 0.048547f
C54 VN.n21 B 0.03367f
C55 VN.n22 B 0.026048f
C56 VN.n23 B 0.026048f
C57 VN.n24 B 0.026048f
C58 VN.n25 B 0.048547f
C59 VN.n26 B 0.032249f
C60 VN.n27 B 0.391195f
C61 VN.n28 B 0.043863f
C62 VN.n29 B 0.034342f
C63 VN.t0 B 0.784334f
C64 VN.n30 B 0.042381f
C65 VN.n31 B 0.026048f
C66 VN.t7 B 0.784334f
C67 VN.n32 B 0.306582f
C68 VN.n33 B 0.026048f
C69 VN.n34 B 0.038025f
C70 VN.n35 B 0.251994f
C71 VN.t5 B 0.784334f
C72 VN.t4 B 0.992437f
C73 VN.n36 B 0.367459f
C74 VN.n37 B 0.380376f
C75 VN.n38 B 0.035125f
C76 VN.n39 B 0.048547f
C77 VN.n40 B 0.026048f
C78 VN.n41 B 0.026048f
C79 VN.n42 B 0.026048f
C80 VN.n43 B 0.038025f
C81 VN.n44 B 0.048547f
C82 VN.n45 B 0.035125f
C83 VN.n46 B 0.026048f
C84 VN.n47 B 0.026048f
C85 VN.n48 B 0.038001f
C86 VN.n49 B 0.048547f
C87 VN.n50 B 0.03367f
C88 VN.n51 B 0.026048f
C89 VN.n52 B 0.026048f
C90 VN.n53 B 0.026048f
C91 VN.n54 B 0.048547f
C92 VN.n55 B 0.032249f
C93 VN.n56 B 0.391195f
C94 VN.n57 B 1.26092f
C95 VTAIL.t3 B 0.088603f
C96 VTAIL.t5 B 0.088603f
C97 VTAIL.n0 B 0.646946f
C98 VTAIL.n1 B 0.436483f
C99 VTAIL.n2 B 0.032186f
C100 VTAIL.n3 B 0.025196f
C101 VTAIL.n4 B 0.013539f
C102 VTAIL.n5 B 0.032002f
C103 VTAIL.n6 B 0.014336f
C104 VTAIL.n7 B 0.419838f
C105 VTAIL.n8 B 0.013539f
C106 VTAIL.t1 B 0.052291f
C107 VTAIL.n9 B 0.098476f
C108 VTAIL.n10 B 0.018886f
C109 VTAIL.n11 B 0.024001f
C110 VTAIL.n12 B 0.032002f
C111 VTAIL.n13 B 0.014336f
C112 VTAIL.n14 B 0.013539f
C113 VTAIL.n15 B 0.025196f
C114 VTAIL.n16 B 0.025196f
C115 VTAIL.n17 B 0.013539f
C116 VTAIL.n18 B 0.014336f
C117 VTAIL.n19 B 0.032002f
C118 VTAIL.n20 B 0.063567f
C119 VTAIL.n21 B 0.014336f
C120 VTAIL.n22 B 0.013539f
C121 VTAIL.n23 B 0.054453f
C122 VTAIL.n24 B 0.034861f
C123 VTAIL.n25 B 0.263299f
C124 VTAIL.n26 B 0.032186f
C125 VTAIL.n27 B 0.025196f
C126 VTAIL.n28 B 0.013539f
C127 VTAIL.n29 B 0.032002f
C128 VTAIL.n30 B 0.014336f
C129 VTAIL.n31 B 0.419838f
C130 VTAIL.n32 B 0.013539f
C131 VTAIL.t11 B 0.052291f
C132 VTAIL.n33 B 0.098476f
C133 VTAIL.n34 B 0.018886f
C134 VTAIL.n35 B 0.024001f
C135 VTAIL.n36 B 0.032002f
C136 VTAIL.n37 B 0.014336f
C137 VTAIL.n38 B 0.013539f
C138 VTAIL.n39 B 0.025196f
C139 VTAIL.n40 B 0.025196f
C140 VTAIL.n41 B 0.013539f
C141 VTAIL.n42 B 0.014336f
C142 VTAIL.n43 B 0.032002f
C143 VTAIL.n44 B 0.063567f
C144 VTAIL.n45 B 0.014336f
C145 VTAIL.n46 B 0.013539f
C146 VTAIL.n47 B 0.054453f
C147 VTAIL.n48 B 0.034861f
C148 VTAIL.n49 B 0.263299f
C149 VTAIL.t13 B 0.088603f
C150 VTAIL.t14 B 0.088603f
C151 VTAIL.n50 B 0.646946f
C152 VTAIL.n51 B 0.637527f
C153 VTAIL.n52 B 0.032186f
C154 VTAIL.n53 B 0.025196f
C155 VTAIL.n54 B 0.013539f
C156 VTAIL.n55 B 0.032002f
C157 VTAIL.n56 B 0.014336f
C158 VTAIL.n57 B 0.419838f
C159 VTAIL.n58 B 0.013539f
C160 VTAIL.t12 B 0.052291f
C161 VTAIL.n59 B 0.098476f
C162 VTAIL.n60 B 0.018886f
C163 VTAIL.n61 B 0.024001f
C164 VTAIL.n62 B 0.032002f
C165 VTAIL.n63 B 0.014336f
C166 VTAIL.n64 B 0.013539f
C167 VTAIL.n65 B 0.025196f
C168 VTAIL.n66 B 0.025196f
C169 VTAIL.n67 B 0.013539f
C170 VTAIL.n68 B 0.014336f
C171 VTAIL.n69 B 0.032002f
C172 VTAIL.n70 B 0.063567f
C173 VTAIL.n71 B 0.014336f
C174 VTAIL.n72 B 0.013539f
C175 VTAIL.n73 B 0.054453f
C176 VTAIL.n74 B 0.034861f
C177 VTAIL.n75 B 1.08464f
C178 VTAIL.n76 B 0.032186f
C179 VTAIL.n77 B 0.025196f
C180 VTAIL.n78 B 0.013539f
C181 VTAIL.n79 B 0.032002f
C182 VTAIL.n80 B 0.014336f
C183 VTAIL.n81 B 0.419838f
C184 VTAIL.n82 B 0.013539f
C185 VTAIL.t7 B 0.052291f
C186 VTAIL.n83 B 0.098476f
C187 VTAIL.n84 B 0.018886f
C188 VTAIL.n85 B 0.024001f
C189 VTAIL.n86 B 0.032002f
C190 VTAIL.n87 B 0.014336f
C191 VTAIL.n88 B 0.013539f
C192 VTAIL.n89 B 0.025196f
C193 VTAIL.n90 B 0.025196f
C194 VTAIL.n91 B 0.013539f
C195 VTAIL.n92 B 0.014336f
C196 VTAIL.n93 B 0.032002f
C197 VTAIL.n94 B 0.063567f
C198 VTAIL.n95 B 0.014336f
C199 VTAIL.n96 B 0.013539f
C200 VTAIL.n97 B 0.054453f
C201 VTAIL.n98 B 0.034861f
C202 VTAIL.n99 B 1.08464f
C203 VTAIL.t0 B 0.088603f
C204 VTAIL.t4 B 0.088603f
C205 VTAIL.n100 B 0.646951f
C206 VTAIL.n101 B 0.637522f
C207 VTAIL.n102 B 0.032186f
C208 VTAIL.n103 B 0.025196f
C209 VTAIL.n104 B 0.013539f
C210 VTAIL.n105 B 0.032002f
C211 VTAIL.n106 B 0.014336f
C212 VTAIL.n107 B 0.419838f
C213 VTAIL.n108 B 0.013539f
C214 VTAIL.t2 B 0.052291f
C215 VTAIL.n109 B 0.098476f
C216 VTAIL.n110 B 0.018886f
C217 VTAIL.n111 B 0.024001f
C218 VTAIL.n112 B 0.032002f
C219 VTAIL.n113 B 0.014336f
C220 VTAIL.n114 B 0.013539f
C221 VTAIL.n115 B 0.025196f
C222 VTAIL.n116 B 0.025196f
C223 VTAIL.n117 B 0.013539f
C224 VTAIL.n118 B 0.014336f
C225 VTAIL.n119 B 0.032002f
C226 VTAIL.n120 B 0.063567f
C227 VTAIL.n121 B 0.014336f
C228 VTAIL.n122 B 0.013539f
C229 VTAIL.n123 B 0.054453f
C230 VTAIL.n124 B 0.034861f
C231 VTAIL.n125 B 0.263299f
C232 VTAIL.n126 B 0.032186f
C233 VTAIL.n127 B 0.025196f
C234 VTAIL.n128 B 0.013539f
C235 VTAIL.n129 B 0.032002f
C236 VTAIL.n130 B 0.014336f
C237 VTAIL.n131 B 0.419838f
C238 VTAIL.n132 B 0.013539f
C239 VTAIL.t10 B 0.052291f
C240 VTAIL.n133 B 0.098476f
C241 VTAIL.n134 B 0.018886f
C242 VTAIL.n135 B 0.024001f
C243 VTAIL.n136 B 0.032002f
C244 VTAIL.n137 B 0.014336f
C245 VTAIL.n138 B 0.013539f
C246 VTAIL.n139 B 0.025196f
C247 VTAIL.n140 B 0.025196f
C248 VTAIL.n141 B 0.013539f
C249 VTAIL.n142 B 0.014336f
C250 VTAIL.n143 B 0.032002f
C251 VTAIL.n144 B 0.063567f
C252 VTAIL.n145 B 0.014336f
C253 VTAIL.n146 B 0.013539f
C254 VTAIL.n147 B 0.054453f
C255 VTAIL.n148 B 0.034861f
C256 VTAIL.n149 B 0.263299f
C257 VTAIL.t8 B 0.088603f
C258 VTAIL.t15 B 0.088603f
C259 VTAIL.n150 B 0.646951f
C260 VTAIL.n151 B 0.637522f
C261 VTAIL.n152 B 0.032186f
C262 VTAIL.n153 B 0.025196f
C263 VTAIL.n154 B 0.013539f
C264 VTAIL.n155 B 0.032002f
C265 VTAIL.n156 B 0.014336f
C266 VTAIL.n157 B 0.419838f
C267 VTAIL.n158 B 0.013539f
C268 VTAIL.t9 B 0.052291f
C269 VTAIL.n159 B 0.098476f
C270 VTAIL.n160 B 0.018886f
C271 VTAIL.n161 B 0.024001f
C272 VTAIL.n162 B 0.032002f
C273 VTAIL.n163 B 0.014336f
C274 VTAIL.n164 B 0.013539f
C275 VTAIL.n165 B 0.025196f
C276 VTAIL.n166 B 0.025196f
C277 VTAIL.n167 B 0.013539f
C278 VTAIL.n168 B 0.014336f
C279 VTAIL.n169 B 0.032002f
C280 VTAIL.n170 B 0.063567f
C281 VTAIL.n171 B 0.014336f
C282 VTAIL.n172 B 0.013539f
C283 VTAIL.n173 B 0.054453f
C284 VTAIL.n174 B 0.034861f
C285 VTAIL.n175 B 1.08464f
C286 VTAIL.n176 B 0.032186f
C287 VTAIL.n177 B 0.025196f
C288 VTAIL.n178 B 0.013539f
C289 VTAIL.n179 B 0.032002f
C290 VTAIL.n180 B 0.014336f
C291 VTAIL.n181 B 0.419838f
C292 VTAIL.n182 B 0.013539f
C293 VTAIL.t6 B 0.052291f
C294 VTAIL.n183 B 0.098476f
C295 VTAIL.n184 B 0.018886f
C296 VTAIL.n185 B 0.024001f
C297 VTAIL.n186 B 0.032002f
C298 VTAIL.n187 B 0.014336f
C299 VTAIL.n188 B 0.013539f
C300 VTAIL.n189 B 0.025196f
C301 VTAIL.n190 B 0.025196f
C302 VTAIL.n191 B 0.013539f
C303 VTAIL.n192 B 0.014336f
C304 VTAIL.n193 B 0.032002f
C305 VTAIL.n194 B 0.063567f
C306 VTAIL.n195 B 0.014336f
C307 VTAIL.n196 B 0.013539f
C308 VTAIL.n197 B 0.054453f
C309 VTAIL.n198 B 0.034861f
C310 VTAIL.n199 B 1.07991f
C311 VDD1.t7 B 0.086962f
C312 VDD1.t0 B 0.086962f
C313 VDD1.n0 B 0.70572f
C314 VDD1.t3 B 0.086962f
C315 VDD1.t5 B 0.086962f
C316 VDD1.n1 B 0.70475f
C317 VDD1.t2 B 0.086962f
C318 VDD1.t6 B 0.086962f
C319 VDD1.n2 B 0.70475f
C320 VDD1.n3 B 2.82515f
C321 VDD1.t1 B 0.086962f
C322 VDD1.t4 B 0.086962f
C323 VDD1.n4 B 0.696001f
C324 VDD1.n5 B 2.36379f
C325 VP.n0 B 0.035643f
C326 VP.t4 B 0.81405f
C327 VP.n1 B 0.043986f
C328 VP.n2 B 0.027035f
C329 VP.t1 B 0.81405f
C330 VP.n3 B 0.318198f
C331 VP.n4 B 0.027035f
C332 VP.n5 B 0.039466f
C333 VP.n6 B 0.027035f
C334 VP.t2 B 0.81405f
C335 VP.n7 B 0.050386f
C336 VP.n8 B 0.027035f
C337 VP.n9 B 0.033471f
C338 VP.n10 B 0.035643f
C339 VP.t6 B 0.81405f
C340 VP.n11 B 0.043986f
C341 VP.n12 B 0.027035f
C342 VP.t0 B 0.81405f
C343 VP.n13 B 0.318198f
C344 VP.n14 B 0.027035f
C345 VP.n15 B 0.039466f
C346 VP.n16 B 0.261541f
C347 VP.t7 B 0.81405f
C348 VP.t5 B 1.03004f
C349 VP.n17 B 0.381381f
C350 VP.n18 B 0.394787f
C351 VP.n19 B 0.036456f
C352 VP.n20 B 0.050386f
C353 VP.n21 B 0.027035f
C354 VP.n22 B 0.027035f
C355 VP.n23 B 0.027035f
C356 VP.n24 B 0.039466f
C357 VP.n25 B 0.050386f
C358 VP.n26 B 0.036456f
C359 VP.n27 B 0.027035f
C360 VP.n28 B 0.027035f
C361 VP.n29 B 0.039441f
C362 VP.n30 B 0.050386f
C363 VP.n31 B 0.034946f
C364 VP.n32 B 0.027035f
C365 VP.n33 B 0.027035f
C366 VP.n34 B 0.027035f
C367 VP.n35 B 0.050386f
C368 VP.n36 B 0.033471f
C369 VP.n37 B 0.406017f
C370 VP.n38 B 1.29392f
C371 VP.t3 B 0.81405f
C372 VP.n39 B 0.406017f
C373 VP.n40 B 1.31541f
C374 VP.n41 B 0.035643f
C375 VP.n42 B 0.027035f
C376 VP.n43 B 0.050386f
C377 VP.n44 B 0.043986f
C378 VP.n45 B 0.034946f
C379 VP.n46 B 0.027035f
C380 VP.n47 B 0.027035f
C381 VP.n48 B 0.027035f
C382 VP.n49 B 0.039441f
C383 VP.n50 B 0.318198f
C384 VP.n51 B 0.036456f
C385 VP.n52 B 0.050386f
C386 VP.n53 B 0.027035f
C387 VP.n54 B 0.027035f
C388 VP.n55 B 0.027035f
C389 VP.n56 B 0.039466f
C390 VP.n57 B 0.050386f
C391 VP.n58 B 0.036456f
C392 VP.n59 B 0.027035f
C393 VP.n60 B 0.027035f
C394 VP.n61 B 0.039441f
C395 VP.n62 B 0.050386f
C396 VP.n63 B 0.034946f
C397 VP.n64 B 0.027035f
C398 VP.n65 B 0.027035f
C399 VP.n66 B 0.027035f
C400 VP.n67 B 0.050386f
C401 VP.n68 B 0.033471f
C402 VP.n69 B 0.406017f
C403 VP.n70 B 0.045525f
.ends

