* NGSPICE file created from diff_pair_sample_0760.ext - technology: sky130A

.subckt diff_pair_sample_0760 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t10 w_n3754_n3372# sky130_fd_pr__pfet_01v8 ad=1.9833 pd=12.35 as=4.6878 ps=24.82 w=12.02 l=1.99
X1 VTAIL.t13 VP.t1 VDD1.t8 w_n3754_n3372# sky130_fd_pr__pfet_01v8 ad=1.9833 pd=12.35 as=1.9833 ps=12.35 w=12.02 l=1.99
X2 B.t11 B.t9 B.t10 w_n3754_n3372# sky130_fd_pr__pfet_01v8 ad=4.6878 pd=24.82 as=0 ps=0 w=12.02 l=1.99
X3 VTAIL.t17 VP.t2 VDD1.t7 w_n3754_n3372# sky130_fd_pr__pfet_01v8 ad=1.9833 pd=12.35 as=1.9833 ps=12.35 w=12.02 l=1.99
X4 VDD1.t6 VP.t3 VTAIL.t19 w_n3754_n3372# sky130_fd_pr__pfet_01v8 ad=4.6878 pd=24.82 as=1.9833 ps=12.35 w=12.02 l=1.99
X5 B.t8 B.t6 B.t7 w_n3754_n3372# sky130_fd_pr__pfet_01v8 ad=4.6878 pd=24.82 as=0 ps=0 w=12.02 l=1.99
X6 VDD2.t9 VN.t0 VTAIL.t8 w_n3754_n3372# sky130_fd_pr__pfet_01v8 ad=1.9833 pd=12.35 as=4.6878 ps=24.82 w=12.02 l=1.99
X7 B.t5 B.t3 B.t4 w_n3754_n3372# sky130_fd_pr__pfet_01v8 ad=4.6878 pd=24.82 as=0 ps=0 w=12.02 l=1.99
X8 VTAIL.t12 VP.t4 VDD1.t5 w_n3754_n3372# sky130_fd_pr__pfet_01v8 ad=1.9833 pd=12.35 as=1.9833 ps=12.35 w=12.02 l=1.99
X9 VTAIL.t4 VN.t1 VDD2.t8 w_n3754_n3372# sky130_fd_pr__pfet_01v8 ad=1.9833 pd=12.35 as=1.9833 ps=12.35 w=12.02 l=1.99
X10 VDD2.t7 VN.t2 VTAIL.t5 w_n3754_n3372# sky130_fd_pr__pfet_01v8 ad=1.9833 pd=12.35 as=1.9833 ps=12.35 w=12.02 l=1.99
X11 VDD1.t4 VP.t5 VTAIL.t16 w_n3754_n3372# sky130_fd_pr__pfet_01v8 ad=4.6878 pd=24.82 as=1.9833 ps=12.35 w=12.02 l=1.99
X12 VDD2.t6 VN.t3 VTAIL.t7 w_n3754_n3372# sky130_fd_pr__pfet_01v8 ad=1.9833 pd=12.35 as=4.6878 ps=24.82 w=12.02 l=1.99
X13 VDD1.t3 VP.t6 VTAIL.t18 w_n3754_n3372# sky130_fd_pr__pfet_01v8 ad=1.9833 pd=12.35 as=4.6878 ps=24.82 w=12.02 l=1.99
X14 VDD2.t5 VN.t4 VTAIL.t0 w_n3754_n3372# sky130_fd_pr__pfet_01v8 ad=4.6878 pd=24.82 as=1.9833 ps=12.35 w=12.02 l=1.99
X15 VDD2.t4 VN.t5 VTAIL.t3 w_n3754_n3372# sky130_fd_pr__pfet_01v8 ad=1.9833 pd=12.35 as=1.9833 ps=12.35 w=12.02 l=1.99
X16 VDD1.t2 VP.t7 VTAIL.t11 w_n3754_n3372# sky130_fd_pr__pfet_01v8 ad=1.9833 pd=12.35 as=1.9833 ps=12.35 w=12.02 l=1.99
X17 VTAIL.t15 VP.t8 VDD1.t1 w_n3754_n3372# sky130_fd_pr__pfet_01v8 ad=1.9833 pd=12.35 as=1.9833 ps=12.35 w=12.02 l=1.99
X18 VDD2.t3 VN.t6 VTAIL.t2 w_n3754_n3372# sky130_fd_pr__pfet_01v8 ad=4.6878 pd=24.82 as=1.9833 ps=12.35 w=12.02 l=1.99
X19 VTAIL.t1 VN.t7 VDD2.t2 w_n3754_n3372# sky130_fd_pr__pfet_01v8 ad=1.9833 pd=12.35 as=1.9833 ps=12.35 w=12.02 l=1.99
X20 VTAIL.t6 VN.t8 VDD2.t1 w_n3754_n3372# sky130_fd_pr__pfet_01v8 ad=1.9833 pd=12.35 as=1.9833 ps=12.35 w=12.02 l=1.99
X21 B.t2 B.t0 B.t1 w_n3754_n3372# sky130_fd_pr__pfet_01v8 ad=4.6878 pd=24.82 as=0 ps=0 w=12.02 l=1.99
X22 VTAIL.t9 VN.t9 VDD2.t0 w_n3754_n3372# sky130_fd_pr__pfet_01v8 ad=1.9833 pd=12.35 as=1.9833 ps=12.35 w=12.02 l=1.99
X23 VDD1.t0 VP.t9 VTAIL.t14 w_n3754_n3372# sky130_fd_pr__pfet_01v8 ad=1.9833 pd=12.35 as=1.9833 ps=12.35 w=12.02 l=1.99
R0 VP.n18 VP.t5 175.816
R1 VP.n20 VP.n19 161.3
R2 VP.n21 VP.n16 161.3
R3 VP.n23 VP.n22 161.3
R4 VP.n24 VP.n15 161.3
R5 VP.n26 VP.n25 161.3
R6 VP.n28 VP.n14 161.3
R7 VP.n30 VP.n29 161.3
R8 VP.n31 VP.n13 161.3
R9 VP.n33 VP.n32 161.3
R10 VP.n34 VP.n12 161.3
R11 VP.n37 VP.n36 161.3
R12 VP.n38 VP.n11 161.3
R13 VP.n40 VP.n39 161.3
R14 VP.n41 VP.n10 161.3
R15 VP.n74 VP.n0 161.3
R16 VP.n73 VP.n72 161.3
R17 VP.n71 VP.n1 161.3
R18 VP.n70 VP.n69 161.3
R19 VP.n67 VP.n2 161.3
R20 VP.n66 VP.n65 161.3
R21 VP.n64 VP.n3 161.3
R22 VP.n63 VP.n62 161.3
R23 VP.n61 VP.n4 161.3
R24 VP.n59 VP.n58 161.3
R25 VP.n57 VP.n5 161.3
R26 VP.n56 VP.n55 161.3
R27 VP.n54 VP.n6 161.3
R28 VP.n53 VP.n52 161.3
R29 VP.n51 VP.n50 161.3
R30 VP.n49 VP.n8 161.3
R31 VP.n48 VP.n47 161.3
R32 VP.n46 VP.n9 161.3
R33 VP.n44 VP.t3 145.57
R34 VP.n7 VP.t2 145.57
R35 VP.n60 VP.t9 145.57
R36 VP.n68 VP.t4 145.57
R37 VP.n75 VP.t0 145.57
R38 VP.n42 VP.t6 145.57
R39 VP.n35 VP.t1 145.57
R40 VP.n27 VP.t7 145.57
R41 VP.n17 VP.t8 145.57
R42 VP.n45 VP.n44 91.7266
R43 VP.n76 VP.n75 91.7266
R44 VP.n43 VP.n42 91.7266
R45 VP.n18 VP.n17 66.4483
R46 VP.n49 VP.n48 56.5617
R47 VP.n73 VP.n1 56.5617
R48 VP.n40 VP.n11 56.5617
R49 VP.n45 VP.n43 49.8254
R50 VP.n55 VP.n5 49.296
R51 VP.n62 VP.n3 49.296
R52 VP.n29 VP.n13 49.296
R53 VP.n22 VP.n15 49.296
R54 VP.n55 VP.n54 31.8581
R55 VP.n66 VP.n3 31.8581
R56 VP.n33 VP.n13 31.8581
R57 VP.n22 VP.n21 31.8581
R58 VP.n48 VP.n9 24.5923
R59 VP.n50 VP.n49 24.5923
R60 VP.n54 VP.n53 24.5923
R61 VP.n59 VP.n5 24.5923
R62 VP.n62 VP.n61 24.5923
R63 VP.n67 VP.n66 24.5923
R64 VP.n69 VP.n1 24.5923
R65 VP.n74 VP.n73 24.5923
R66 VP.n41 VP.n40 24.5923
R67 VP.n34 VP.n33 24.5923
R68 VP.n36 VP.n11 24.5923
R69 VP.n26 VP.n15 24.5923
R70 VP.n29 VP.n28 24.5923
R71 VP.n21 VP.n20 24.5923
R72 VP.n50 VP.n7 21.1495
R73 VP.n69 VP.n68 21.1495
R74 VP.n36 VP.n35 21.1495
R75 VP.n44 VP.n9 19.1821
R76 VP.n75 VP.n74 19.1821
R77 VP.n42 VP.n41 19.1821
R78 VP.n19 VP.n18 13.4112
R79 VP.n60 VP.n59 12.2964
R80 VP.n61 VP.n60 12.2964
R81 VP.n27 VP.n26 12.2964
R82 VP.n28 VP.n27 12.2964
R83 VP.n53 VP.n7 3.44336
R84 VP.n68 VP.n67 3.44336
R85 VP.n35 VP.n34 3.44336
R86 VP.n20 VP.n17 3.44336
R87 VP.n43 VP.n10 0.278335
R88 VP.n46 VP.n45 0.278335
R89 VP.n76 VP.n0 0.278335
R90 VP.n19 VP.n16 0.189894
R91 VP.n23 VP.n16 0.189894
R92 VP.n24 VP.n23 0.189894
R93 VP.n25 VP.n24 0.189894
R94 VP.n25 VP.n14 0.189894
R95 VP.n30 VP.n14 0.189894
R96 VP.n31 VP.n30 0.189894
R97 VP.n32 VP.n31 0.189894
R98 VP.n32 VP.n12 0.189894
R99 VP.n37 VP.n12 0.189894
R100 VP.n38 VP.n37 0.189894
R101 VP.n39 VP.n38 0.189894
R102 VP.n39 VP.n10 0.189894
R103 VP.n47 VP.n46 0.189894
R104 VP.n47 VP.n8 0.189894
R105 VP.n51 VP.n8 0.189894
R106 VP.n52 VP.n51 0.189894
R107 VP.n52 VP.n6 0.189894
R108 VP.n56 VP.n6 0.189894
R109 VP.n57 VP.n56 0.189894
R110 VP.n58 VP.n57 0.189894
R111 VP.n58 VP.n4 0.189894
R112 VP.n63 VP.n4 0.189894
R113 VP.n64 VP.n63 0.189894
R114 VP.n65 VP.n64 0.189894
R115 VP.n65 VP.n2 0.189894
R116 VP.n70 VP.n2 0.189894
R117 VP.n71 VP.n70 0.189894
R118 VP.n72 VP.n71 0.189894
R119 VP.n72 VP.n0 0.189894
R120 VP VP.n76 0.153485
R121 VTAIL.n272 VTAIL.n212 756.745
R122 VTAIL.n62 VTAIL.n2 756.745
R123 VTAIL.n206 VTAIL.n146 756.745
R124 VTAIL.n136 VTAIL.n76 756.745
R125 VTAIL.n232 VTAIL.n231 585
R126 VTAIL.n237 VTAIL.n236 585
R127 VTAIL.n239 VTAIL.n238 585
R128 VTAIL.n228 VTAIL.n227 585
R129 VTAIL.n245 VTAIL.n244 585
R130 VTAIL.n247 VTAIL.n246 585
R131 VTAIL.n224 VTAIL.n223 585
R132 VTAIL.n254 VTAIL.n253 585
R133 VTAIL.n255 VTAIL.n222 585
R134 VTAIL.n257 VTAIL.n256 585
R135 VTAIL.n220 VTAIL.n219 585
R136 VTAIL.n263 VTAIL.n262 585
R137 VTAIL.n265 VTAIL.n264 585
R138 VTAIL.n216 VTAIL.n215 585
R139 VTAIL.n271 VTAIL.n270 585
R140 VTAIL.n273 VTAIL.n272 585
R141 VTAIL.n22 VTAIL.n21 585
R142 VTAIL.n27 VTAIL.n26 585
R143 VTAIL.n29 VTAIL.n28 585
R144 VTAIL.n18 VTAIL.n17 585
R145 VTAIL.n35 VTAIL.n34 585
R146 VTAIL.n37 VTAIL.n36 585
R147 VTAIL.n14 VTAIL.n13 585
R148 VTAIL.n44 VTAIL.n43 585
R149 VTAIL.n45 VTAIL.n12 585
R150 VTAIL.n47 VTAIL.n46 585
R151 VTAIL.n10 VTAIL.n9 585
R152 VTAIL.n53 VTAIL.n52 585
R153 VTAIL.n55 VTAIL.n54 585
R154 VTAIL.n6 VTAIL.n5 585
R155 VTAIL.n61 VTAIL.n60 585
R156 VTAIL.n63 VTAIL.n62 585
R157 VTAIL.n207 VTAIL.n206 585
R158 VTAIL.n205 VTAIL.n204 585
R159 VTAIL.n150 VTAIL.n149 585
R160 VTAIL.n199 VTAIL.n198 585
R161 VTAIL.n197 VTAIL.n196 585
R162 VTAIL.n154 VTAIL.n153 585
R163 VTAIL.n191 VTAIL.n190 585
R164 VTAIL.n189 VTAIL.n156 585
R165 VTAIL.n188 VTAIL.n187 585
R166 VTAIL.n159 VTAIL.n157 585
R167 VTAIL.n182 VTAIL.n181 585
R168 VTAIL.n180 VTAIL.n179 585
R169 VTAIL.n163 VTAIL.n162 585
R170 VTAIL.n174 VTAIL.n173 585
R171 VTAIL.n172 VTAIL.n171 585
R172 VTAIL.n167 VTAIL.n166 585
R173 VTAIL.n137 VTAIL.n136 585
R174 VTAIL.n135 VTAIL.n134 585
R175 VTAIL.n80 VTAIL.n79 585
R176 VTAIL.n129 VTAIL.n128 585
R177 VTAIL.n127 VTAIL.n126 585
R178 VTAIL.n84 VTAIL.n83 585
R179 VTAIL.n121 VTAIL.n120 585
R180 VTAIL.n119 VTAIL.n86 585
R181 VTAIL.n118 VTAIL.n117 585
R182 VTAIL.n89 VTAIL.n87 585
R183 VTAIL.n112 VTAIL.n111 585
R184 VTAIL.n110 VTAIL.n109 585
R185 VTAIL.n93 VTAIL.n92 585
R186 VTAIL.n104 VTAIL.n103 585
R187 VTAIL.n102 VTAIL.n101 585
R188 VTAIL.n97 VTAIL.n96 585
R189 VTAIL.n233 VTAIL.t7 329.036
R190 VTAIL.n23 VTAIL.t10 329.036
R191 VTAIL.n168 VTAIL.t18 329.036
R192 VTAIL.n98 VTAIL.t8 329.036
R193 VTAIL.n237 VTAIL.n231 171.744
R194 VTAIL.n238 VTAIL.n237 171.744
R195 VTAIL.n238 VTAIL.n227 171.744
R196 VTAIL.n245 VTAIL.n227 171.744
R197 VTAIL.n246 VTAIL.n245 171.744
R198 VTAIL.n246 VTAIL.n223 171.744
R199 VTAIL.n254 VTAIL.n223 171.744
R200 VTAIL.n255 VTAIL.n254 171.744
R201 VTAIL.n256 VTAIL.n255 171.744
R202 VTAIL.n256 VTAIL.n219 171.744
R203 VTAIL.n263 VTAIL.n219 171.744
R204 VTAIL.n264 VTAIL.n263 171.744
R205 VTAIL.n264 VTAIL.n215 171.744
R206 VTAIL.n271 VTAIL.n215 171.744
R207 VTAIL.n272 VTAIL.n271 171.744
R208 VTAIL.n27 VTAIL.n21 171.744
R209 VTAIL.n28 VTAIL.n27 171.744
R210 VTAIL.n28 VTAIL.n17 171.744
R211 VTAIL.n35 VTAIL.n17 171.744
R212 VTAIL.n36 VTAIL.n35 171.744
R213 VTAIL.n36 VTAIL.n13 171.744
R214 VTAIL.n44 VTAIL.n13 171.744
R215 VTAIL.n45 VTAIL.n44 171.744
R216 VTAIL.n46 VTAIL.n45 171.744
R217 VTAIL.n46 VTAIL.n9 171.744
R218 VTAIL.n53 VTAIL.n9 171.744
R219 VTAIL.n54 VTAIL.n53 171.744
R220 VTAIL.n54 VTAIL.n5 171.744
R221 VTAIL.n61 VTAIL.n5 171.744
R222 VTAIL.n62 VTAIL.n61 171.744
R223 VTAIL.n206 VTAIL.n205 171.744
R224 VTAIL.n205 VTAIL.n149 171.744
R225 VTAIL.n198 VTAIL.n149 171.744
R226 VTAIL.n198 VTAIL.n197 171.744
R227 VTAIL.n197 VTAIL.n153 171.744
R228 VTAIL.n190 VTAIL.n153 171.744
R229 VTAIL.n190 VTAIL.n189 171.744
R230 VTAIL.n189 VTAIL.n188 171.744
R231 VTAIL.n188 VTAIL.n157 171.744
R232 VTAIL.n181 VTAIL.n157 171.744
R233 VTAIL.n181 VTAIL.n180 171.744
R234 VTAIL.n180 VTAIL.n162 171.744
R235 VTAIL.n173 VTAIL.n162 171.744
R236 VTAIL.n173 VTAIL.n172 171.744
R237 VTAIL.n172 VTAIL.n166 171.744
R238 VTAIL.n136 VTAIL.n135 171.744
R239 VTAIL.n135 VTAIL.n79 171.744
R240 VTAIL.n128 VTAIL.n79 171.744
R241 VTAIL.n128 VTAIL.n127 171.744
R242 VTAIL.n127 VTAIL.n83 171.744
R243 VTAIL.n120 VTAIL.n83 171.744
R244 VTAIL.n120 VTAIL.n119 171.744
R245 VTAIL.n119 VTAIL.n118 171.744
R246 VTAIL.n118 VTAIL.n87 171.744
R247 VTAIL.n111 VTAIL.n87 171.744
R248 VTAIL.n111 VTAIL.n110 171.744
R249 VTAIL.n110 VTAIL.n92 171.744
R250 VTAIL.n103 VTAIL.n92 171.744
R251 VTAIL.n103 VTAIL.n102 171.744
R252 VTAIL.n102 VTAIL.n96 171.744
R253 VTAIL.t7 VTAIL.n231 85.8723
R254 VTAIL.t10 VTAIL.n21 85.8723
R255 VTAIL.t18 VTAIL.n166 85.8723
R256 VTAIL.t8 VTAIL.n96 85.8723
R257 VTAIL.n145 VTAIL.n144 55.221
R258 VTAIL.n143 VTAIL.n142 55.221
R259 VTAIL.n75 VTAIL.n74 55.221
R260 VTAIL.n73 VTAIL.n72 55.221
R261 VTAIL.n279 VTAIL.n278 55.2208
R262 VTAIL.n1 VTAIL.n0 55.2208
R263 VTAIL.n69 VTAIL.n68 55.2208
R264 VTAIL.n71 VTAIL.n70 55.2208
R265 VTAIL.n277 VTAIL.n276 30.246
R266 VTAIL.n67 VTAIL.n66 30.246
R267 VTAIL.n211 VTAIL.n210 30.246
R268 VTAIL.n141 VTAIL.n140 30.246
R269 VTAIL.n73 VTAIL.n71 26.7289
R270 VTAIL.n277 VTAIL.n211 24.7289
R271 VTAIL.n257 VTAIL.n222 13.1884
R272 VTAIL.n47 VTAIL.n12 13.1884
R273 VTAIL.n191 VTAIL.n156 13.1884
R274 VTAIL.n121 VTAIL.n86 13.1884
R275 VTAIL.n253 VTAIL.n252 12.8005
R276 VTAIL.n258 VTAIL.n220 12.8005
R277 VTAIL.n43 VTAIL.n42 12.8005
R278 VTAIL.n48 VTAIL.n10 12.8005
R279 VTAIL.n192 VTAIL.n154 12.8005
R280 VTAIL.n187 VTAIL.n158 12.8005
R281 VTAIL.n122 VTAIL.n84 12.8005
R282 VTAIL.n117 VTAIL.n88 12.8005
R283 VTAIL.n251 VTAIL.n224 12.0247
R284 VTAIL.n262 VTAIL.n261 12.0247
R285 VTAIL.n41 VTAIL.n14 12.0247
R286 VTAIL.n52 VTAIL.n51 12.0247
R287 VTAIL.n196 VTAIL.n195 12.0247
R288 VTAIL.n186 VTAIL.n159 12.0247
R289 VTAIL.n126 VTAIL.n125 12.0247
R290 VTAIL.n116 VTAIL.n89 12.0247
R291 VTAIL.n248 VTAIL.n247 11.249
R292 VTAIL.n265 VTAIL.n218 11.249
R293 VTAIL.n38 VTAIL.n37 11.249
R294 VTAIL.n55 VTAIL.n8 11.249
R295 VTAIL.n199 VTAIL.n152 11.249
R296 VTAIL.n183 VTAIL.n182 11.249
R297 VTAIL.n129 VTAIL.n82 11.249
R298 VTAIL.n113 VTAIL.n112 11.249
R299 VTAIL.n233 VTAIL.n232 10.7239
R300 VTAIL.n23 VTAIL.n22 10.7239
R301 VTAIL.n168 VTAIL.n167 10.7239
R302 VTAIL.n98 VTAIL.n97 10.7239
R303 VTAIL.n244 VTAIL.n226 10.4732
R304 VTAIL.n266 VTAIL.n216 10.4732
R305 VTAIL.n34 VTAIL.n16 10.4732
R306 VTAIL.n56 VTAIL.n6 10.4732
R307 VTAIL.n200 VTAIL.n150 10.4732
R308 VTAIL.n179 VTAIL.n161 10.4732
R309 VTAIL.n130 VTAIL.n80 10.4732
R310 VTAIL.n109 VTAIL.n91 10.4732
R311 VTAIL.n243 VTAIL.n228 9.69747
R312 VTAIL.n270 VTAIL.n269 9.69747
R313 VTAIL.n33 VTAIL.n18 9.69747
R314 VTAIL.n60 VTAIL.n59 9.69747
R315 VTAIL.n204 VTAIL.n203 9.69747
R316 VTAIL.n178 VTAIL.n163 9.69747
R317 VTAIL.n134 VTAIL.n133 9.69747
R318 VTAIL.n108 VTAIL.n93 9.69747
R319 VTAIL.n276 VTAIL.n275 9.45567
R320 VTAIL.n66 VTAIL.n65 9.45567
R321 VTAIL.n210 VTAIL.n209 9.45567
R322 VTAIL.n140 VTAIL.n139 9.45567
R323 VTAIL.n275 VTAIL.n274 9.3005
R324 VTAIL.n214 VTAIL.n213 9.3005
R325 VTAIL.n269 VTAIL.n268 9.3005
R326 VTAIL.n267 VTAIL.n266 9.3005
R327 VTAIL.n218 VTAIL.n217 9.3005
R328 VTAIL.n261 VTAIL.n260 9.3005
R329 VTAIL.n259 VTAIL.n258 9.3005
R330 VTAIL.n235 VTAIL.n234 9.3005
R331 VTAIL.n230 VTAIL.n229 9.3005
R332 VTAIL.n241 VTAIL.n240 9.3005
R333 VTAIL.n243 VTAIL.n242 9.3005
R334 VTAIL.n226 VTAIL.n225 9.3005
R335 VTAIL.n249 VTAIL.n248 9.3005
R336 VTAIL.n251 VTAIL.n250 9.3005
R337 VTAIL.n252 VTAIL.n221 9.3005
R338 VTAIL.n65 VTAIL.n64 9.3005
R339 VTAIL.n4 VTAIL.n3 9.3005
R340 VTAIL.n59 VTAIL.n58 9.3005
R341 VTAIL.n57 VTAIL.n56 9.3005
R342 VTAIL.n8 VTAIL.n7 9.3005
R343 VTAIL.n51 VTAIL.n50 9.3005
R344 VTAIL.n49 VTAIL.n48 9.3005
R345 VTAIL.n25 VTAIL.n24 9.3005
R346 VTAIL.n20 VTAIL.n19 9.3005
R347 VTAIL.n31 VTAIL.n30 9.3005
R348 VTAIL.n33 VTAIL.n32 9.3005
R349 VTAIL.n16 VTAIL.n15 9.3005
R350 VTAIL.n39 VTAIL.n38 9.3005
R351 VTAIL.n41 VTAIL.n40 9.3005
R352 VTAIL.n42 VTAIL.n11 9.3005
R353 VTAIL.n170 VTAIL.n169 9.3005
R354 VTAIL.n165 VTAIL.n164 9.3005
R355 VTAIL.n176 VTAIL.n175 9.3005
R356 VTAIL.n178 VTAIL.n177 9.3005
R357 VTAIL.n161 VTAIL.n160 9.3005
R358 VTAIL.n184 VTAIL.n183 9.3005
R359 VTAIL.n186 VTAIL.n185 9.3005
R360 VTAIL.n158 VTAIL.n155 9.3005
R361 VTAIL.n209 VTAIL.n208 9.3005
R362 VTAIL.n148 VTAIL.n147 9.3005
R363 VTAIL.n203 VTAIL.n202 9.3005
R364 VTAIL.n201 VTAIL.n200 9.3005
R365 VTAIL.n152 VTAIL.n151 9.3005
R366 VTAIL.n195 VTAIL.n194 9.3005
R367 VTAIL.n193 VTAIL.n192 9.3005
R368 VTAIL.n100 VTAIL.n99 9.3005
R369 VTAIL.n95 VTAIL.n94 9.3005
R370 VTAIL.n106 VTAIL.n105 9.3005
R371 VTAIL.n108 VTAIL.n107 9.3005
R372 VTAIL.n91 VTAIL.n90 9.3005
R373 VTAIL.n114 VTAIL.n113 9.3005
R374 VTAIL.n116 VTAIL.n115 9.3005
R375 VTAIL.n88 VTAIL.n85 9.3005
R376 VTAIL.n139 VTAIL.n138 9.3005
R377 VTAIL.n78 VTAIL.n77 9.3005
R378 VTAIL.n133 VTAIL.n132 9.3005
R379 VTAIL.n131 VTAIL.n130 9.3005
R380 VTAIL.n82 VTAIL.n81 9.3005
R381 VTAIL.n125 VTAIL.n124 9.3005
R382 VTAIL.n123 VTAIL.n122 9.3005
R383 VTAIL.n240 VTAIL.n239 8.92171
R384 VTAIL.n273 VTAIL.n214 8.92171
R385 VTAIL.n30 VTAIL.n29 8.92171
R386 VTAIL.n63 VTAIL.n4 8.92171
R387 VTAIL.n207 VTAIL.n148 8.92171
R388 VTAIL.n175 VTAIL.n174 8.92171
R389 VTAIL.n137 VTAIL.n78 8.92171
R390 VTAIL.n105 VTAIL.n104 8.92171
R391 VTAIL.n236 VTAIL.n230 8.14595
R392 VTAIL.n274 VTAIL.n212 8.14595
R393 VTAIL.n26 VTAIL.n20 8.14595
R394 VTAIL.n64 VTAIL.n2 8.14595
R395 VTAIL.n208 VTAIL.n146 8.14595
R396 VTAIL.n171 VTAIL.n165 8.14595
R397 VTAIL.n138 VTAIL.n76 8.14595
R398 VTAIL.n101 VTAIL.n95 8.14595
R399 VTAIL.n235 VTAIL.n232 7.3702
R400 VTAIL.n25 VTAIL.n22 7.3702
R401 VTAIL.n170 VTAIL.n167 7.3702
R402 VTAIL.n100 VTAIL.n97 7.3702
R403 VTAIL.n236 VTAIL.n235 5.81868
R404 VTAIL.n276 VTAIL.n212 5.81868
R405 VTAIL.n26 VTAIL.n25 5.81868
R406 VTAIL.n66 VTAIL.n2 5.81868
R407 VTAIL.n210 VTAIL.n146 5.81868
R408 VTAIL.n171 VTAIL.n170 5.81868
R409 VTAIL.n140 VTAIL.n76 5.81868
R410 VTAIL.n101 VTAIL.n100 5.81868
R411 VTAIL.n239 VTAIL.n230 5.04292
R412 VTAIL.n274 VTAIL.n273 5.04292
R413 VTAIL.n29 VTAIL.n20 5.04292
R414 VTAIL.n64 VTAIL.n63 5.04292
R415 VTAIL.n208 VTAIL.n207 5.04292
R416 VTAIL.n174 VTAIL.n165 5.04292
R417 VTAIL.n138 VTAIL.n137 5.04292
R418 VTAIL.n104 VTAIL.n95 5.04292
R419 VTAIL.n240 VTAIL.n228 4.26717
R420 VTAIL.n270 VTAIL.n214 4.26717
R421 VTAIL.n30 VTAIL.n18 4.26717
R422 VTAIL.n60 VTAIL.n4 4.26717
R423 VTAIL.n204 VTAIL.n148 4.26717
R424 VTAIL.n175 VTAIL.n163 4.26717
R425 VTAIL.n134 VTAIL.n78 4.26717
R426 VTAIL.n105 VTAIL.n93 4.26717
R427 VTAIL.n244 VTAIL.n243 3.49141
R428 VTAIL.n269 VTAIL.n216 3.49141
R429 VTAIL.n34 VTAIL.n33 3.49141
R430 VTAIL.n59 VTAIL.n6 3.49141
R431 VTAIL.n203 VTAIL.n150 3.49141
R432 VTAIL.n179 VTAIL.n178 3.49141
R433 VTAIL.n133 VTAIL.n80 3.49141
R434 VTAIL.n109 VTAIL.n108 3.49141
R435 VTAIL.n247 VTAIL.n226 2.71565
R436 VTAIL.n266 VTAIL.n265 2.71565
R437 VTAIL.n37 VTAIL.n16 2.71565
R438 VTAIL.n56 VTAIL.n55 2.71565
R439 VTAIL.n200 VTAIL.n199 2.71565
R440 VTAIL.n182 VTAIL.n161 2.71565
R441 VTAIL.n130 VTAIL.n129 2.71565
R442 VTAIL.n112 VTAIL.n91 2.71565
R443 VTAIL.n278 VTAIL.t3 2.70474
R444 VTAIL.n278 VTAIL.t9 2.70474
R445 VTAIL.n0 VTAIL.t0 2.70474
R446 VTAIL.n0 VTAIL.t1 2.70474
R447 VTAIL.n68 VTAIL.t14 2.70474
R448 VTAIL.n68 VTAIL.t12 2.70474
R449 VTAIL.n70 VTAIL.t19 2.70474
R450 VTAIL.n70 VTAIL.t17 2.70474
R451 VTAIL.n144 VTAIL.t11 2.70474
R452 VTAIL.n144 VTAIL.t13 2.70474
R453 VTAIL.n142 VTAIL.t16 2.70474
R454 VTAIL.n142 VTAIL.t15 2.70474
R455 VTAIL.n74 VTAIL.t5 2.70474
R456 VTAIL.n74 VTAIL.t4 2.70474
R457 VTAIL.n72 VTAIL.t2 2.70474
R458 VTAIL.n72 VTAIL.t6 2.70474
R459 VTAIL.n169 VTAIL.n168 2.41282
R460 VTAIL.n99 VTAIL.n98 2.41282
R461 VTAIL.n234 VTAIL.n233 2.41282
R462 VTAIL.n24 VTAIL.n23 2.41282
R463 VTAIL.n75 VTAIL.n73 2.0005
R464 VTAIL.n141 VTAIL.n75 2.0005
R465 VTAIL.n145 VTAIL.n143 2.0005
R466 VTAIL.n211 VTAIL.n145 2.0005
R467 VTAIL.n71 VTAIL.n69 2.0005
R468 VTAIL.n69 VTAIL.n67 2.0005
R469 VTAIL.n279 VTAIL.n277 2.0005
R470 VTAIL.n248 VTAIL.n224 1.93989
R471 VTAIL.n262 VTAIL.n218 1.93989
R472 VTAIL.n38 VTAIL.n14 1.93989
R473 VTAIL.n52 VTAIL.n8 1.93989
R474 VTAIL.n196 VTAIL.n152 1.93989
R475 VTAIL.n183 VTAIL.n159 1.93989
R476 VTAIL.n126 VTAIL.n82 1.93989
R477 VTAIL.n113 VTAIL.n89 1.93989
R478 VTAIL VTAIL.n1 1.55869
R479 VTAIL.n143 VTAIL.n141 1.47033
R480 VTAIL.n67 VTAIL.n1 1.47033
R481 VTAIL.n253 VTAIL.n251 1.16414
R482 VTAIL.n261 VTAIL.n220 1.16414
R483 VTAIL.n43 VTAIL.n41 1.16414
R484 VTAIL.n51 VTAIL.n10 1.16414
R485 VTAIL.n195 VTAIL.n154 1.16414
R486 VTAIL.n187 VTAIL.n186 1.16414
R487 VTAIL.n125 VTAIL.n84 1.16414
R488 VTAIL.n117 VTAIL.n116 1.16414
R489 VTAIL VTAIL.n279 0.44231
R490 VTAIL.n252 VTAIL.n222 0.388379
R491 VTAIL.n258 VTAIL.n257 0.388379
R492 VTAIL.n42 VTAIL.n12 0.388379
R493 VTAIL.n48 VTAIL.n47 0.388379
R494 VTAIL.n192 VTAIL.n191 0.388379
R495 VTAIL.n158 VTAIL.n156 0.388379
R496 VTAIL.n122 VTAIL.n121 0.388379
R497 VTAIL.n88 VTAIL.n86 0.388379
R498 VTAIL.n234 VTAIL.n229 0.155672
R499 VTAIL.n241 VTAIL.n229 0.155672
R500 VTAIL.n242 VTAIL.n241 0.155672
R501 VTAIL.n242 VTAIL.n225 0.155672
R502 VTAIL.n249 VTAIL.n225 0.155672
R503 VTAIL.n250 VTAIL.n249 0.155672
R504 VTAIL.n250 VTAIL.n221 0.155672
R505 VTAIL.n259 VTAIL.n221 0.155672
R506 VTAIL.n260 VTAIL.n259 0.155672
R507 VTAIL.n260 VTAIL.n217 0.155672
R508 VTAIL.n267 VTAIL.n217 0.155672
R509 VTAIL.n268 VTAIL.n267 0.155672
R510 VTAIL.n268 VTAIL.n213 0.155672
R511 VTAIL.n275 VTAIL.n213 0.155672
R512 VTAIL.n24 VTAIL.n19 0.155672
R513 VTAIL.n31 VTAIL.n19 0.155672
R514 VTAIL.n32 VTAIL.n31 0.155672
R515 VTAIL.n32 VTAIL.n15 0.155672
R516 VTAIL.n39 VTAIL.n15 0.155672
R517 VTAIL.n40 VTAIL.n39 0.155672
R518 VTAIL.n40 VTAIL.n11 0.155672
R519 VTAIL.n49 VTAIL.n11 0.155672
R520 VTAIL.n50 VTAIL.n49 0.155672
R521 VTAIL.n50 VTAIL.n7 0.155672
R522 VTAIL.n57 VTAIL.n7 0.155672
R523 VTAIL.n58 VTAIL.n57 0.155672
R524 VTAIL.n58 VTAIL.n3 0.155672
R525 VTAIL.n65 VTAIL.n3 0.155672
R526 VTAIL.n209 VTAIL.n147 0.155672
R527 VTAIL.n202 VTAIL.n147 0.155672
R528 VTAIL.n202 VTAIL.n201 0.155672
R529 VTAIL.n201 VTAIL.n151 0.155672
R530 VTAIL.n194 VTAIL.n151 0.155672
R531 VTAIL.n194 VTAIL.n193 0.155672
R532 VTAIL.n193 VTAIL.n155 0.155672
R533 VTAIL.n185 VTAIL.n155 0.155672
R534 VTAIL.n185 VTAIL.n184 0.155672
R535 VTAIL.n184 VTAIL.n160 0.155672
R536 VTAIL.n177 VTAIL.n160 0.155672
R537 VTAIL.n177 VTAIL.n176 0.155672
R538 VTAIL.n176 VTAIL.n164 0.155672
R539 VTAIL.n169 VTAIL.n164 0.155672
R540 VTAIL.n139 VTAIL.n77 0.155672
R541 VTAIL.n132 VTAIL.n77 0.155672
R542 VTAIL.n132 VTAIL.n131 0.155672
R543 VTAIL.n131 VTAIL.n81 0.155672
R544 VTAIL.n124 VTAIL.n81 0.155672
R545 VTAIL.n124 VTAIL.n123 0.155672
R546 VTAIL.n123 VTAIL.n85 0.155672
R547 VTAIL.n115 VTAIL.n85 0.155672
R548 VTAIL.n115 VTAIL.n114 0.155672
R549 VTAIL.n114 VTAIL.n90 0.155672
R550 VTAIL.n107 VTAIL.n90 0.155672
R551 VTAIL.n107 VTAIL.n106 0.155672
R552 VTAIL.n106 VTAIL.n94 0.155672
R553 VTAIL.n99 VTAIL.n94 0.155672
R554 VDD1.n60 VDD1.n0 756.745
R555 VDD1.n127 VDD1.n67 756.745
R556 VDD1.n61 VDD1.n60 585
R557 VDD1.n59 VDD1.n58 585
R558 VDD1.n4 VDD1.n3 585
R559 VDD1.n53 VDD1.n52 585
R560 VDD1.n51 VDD1.n50 585
R561 VDD1.n8 VDD1.n7 585
R562 VDD1.n45 VDD1.n44 585
R563 VDD1.n43 VDD1.n10 585
R564 VDD1.n42 VDD1.n41 585
R565 VDD1.n13 VDD1.n11 585
R566 VDD1.n36 VDD1.n35 585
R567 VDD1.n34 VDD1.n33 585
R568 VDD1.n17 VDD1.n16 585
R569 VDD1.n28 VDD1.n27 585
R570 VDD1.n26 VDD1.n25 585
R571 VDD1.n21 VDD1.n20 585
R572 VDD1.n87 VDD1.n86 585
R573 VDD1.n92 VDD1.n91 585
R574 VDD1.n94 VDD1.n93 585
R575 VDD1.n83 VDD1.n82 585
R576 VDD1.n100 VDD1.n99 585
R577 VDD1.n102 VDD1.n101 585
R578 VDD1.n79 VDD1.n78 585
R579 VDD1.n109 VDD1.n108 585
R580 VDD1.n110 VDD1.n77 585
R581 VDD1.n112 VDD1.n111 585
R582 VDD1.n75 VDD1.n74 585
R583 VDD1.n118 VDD1.n117 585
R584 VDD1.n120 VDD1.n119 585
R585 VDD1.n71 VDD1.n70 585
R586 VDD1.n126 VDD1.n125 585
R587 VDD1.n128 VDD1.n127 585
R588 VDD1.n22 VDD1.t4 329.036
R589 VDD1.n88 VDD1.t6 329.036
R590 VDD1.n60 VDD1.n59 171.744
R591 VDD1.n59 VDD1.n3 171.744
R592 VDD1.n52 VDD1.n3 171.744
R593 VDD1.n52 VDD1.n51 171.744
R594 VDD1.n51 VDD1.n7 171.744
R595 VDD1.n44 VDD1.n7 171.744
R596 VDD1.n44 VDD1.n43 171.744
R597 VDD1.n43 VDD1.n42 171.744
R598 VDD1.n42 VDD1.n11 171.744
R599 VDD1.n35 VDD1.n11 171.744
R600 VDD1.n35 VDD1.n34 171.744
R601 VDD1.n34 VDD1.n16 171.744
R602 VDD1.n27 VDD1.n16 171.744
R603 VDD1.n27 VDD1.n26 171.744
R604 VDD1.n26 VDD1.n20 171.744
R605 VDD1.n92 VDD1.n86 171.744
R606 VDD1.n93 VDD1.n92 171.744
R607 VDD1.n93 VDD1.n82 171.744
R608 VDD1.n100 VDD1.n82 171.744
R609 VDD1.n101 VDD1.n100 171.744
R610 VDD1.n101 VDD1.n78 171.744
R611 VDD1.n109 VDD1.n78 171.744
R612 VDD1.n110 VDD1.n109 171.744
R613 VDD1.n111 VDD1.n110 171.744
R614 VDD1.n111 VDD1.n74 171.744
R615 VDD1.n118 VDD1.n74 171.744
R616 VDD1.n119 VDD1.n118 171.744
R617 VDD1.n119 VDD1.n70 171.744
R618 VDD1.n126 VDD1.n70 171.744
R619 VDD1.n127 VDD1.n126 171.744
R620 VDD1.t4 VDD1.n20 85.8723
R621 VDD1.t6 VDD1.n86 85.8723
R622 VDD1.n135 VDD1.n134 73.3443
R623 VDD1.n66 VDD1.n65 71.8998
R624 VDD1.n137 VDD1.n136 71.8996
R625 VDD1.n133 VDD1.n132 71.8996
R626 VDD1.n66 VDD1.n64 48.9247
R627 VDD1.n133 VDD1.n131 48.9247
R628 VDD1.n137 VDD1.n135 45.1604
R629 VDD1.n45 VDD1.n10 13.1884
R630 VDD1.n112 VDD1.n77 13.1884
R631 VDD1.n46 VDD1.n8 12.8005
R632 VDD1.n41 VDD1.n12 12.8005
R633 VDD1.n108 VDD1.n107 12.8005
R634 VDD1.n113 VDD1.n75 12.8005
R635 VDD1.n50 VDD1.n49 12.0247
R636 VDD1.n40 VDD1.n13 12.0247
R637 VDD1.n106 VDD1.n79 12.0247
R638 VDD1.n117 VDD1.n116 12.0247
R639 VDD1.n53 VDD1.n6 11.249
R640 VDD1.n37 VDD1.n36 11.249
R641 VDD1.n103 VDD1.n102 11.249
R642 VDD1.n120 VDD1.n73 11.249
R643 VDD1.n22 VDD1.n21 10.7239
R644 VDD1.n88 VDD1.n87 10.7239
R645 VDD1.n54 VDD1.n4 10.4732
R646 VDD1.n33 VDD1.n15 10.4732
R647 VDD1.n99 VDD1.n81 10.4732
R648 VDD1.n121 VDD1.n71 10.4732
R649 VDD1.n58 VDD1.n57 9.69747
R650 VDD1.n32 VDD1.n17 9.69747
R651 VDD1.n98 VDD1.n83 9.69747
R652 VDD1.n125 VDD1.n124 9.69747
R653 VDD1.n64 VDD1.n63 9.45567
R654 VDD1.n131 VDD1.n130 9.45567
R655 VDD1.n24 VDD1.n23 9.3005
R656 VDD1.n19 VDD1.n18 9.3005
R657 VDD1.n30 VDD1.n29 9.3005
R658 VDD1.n32 VDD1.n31 9.3005
R659 VDD1.n15 VDD1.n14 9.3005
R660 VDD1.n38 VDD1.n37 9.3005
R661 VDD1.n40 VDD1.n39 9.3005
R662 VDD1.n12 VDD1.n9 9.3005
R663 VDD1.n63 VDD1.n62 9.3005
R664 VDD1.n2 VDD1.n1 9.3005
R665 VDD1.n57 VDD1.n56 9.3005
R666 VDD1.n55 VDD1.n54 9.3005
R667 VDD1.n6 VDD1.n5 9.3005
R668 VDD1.n49 VDD1.n48 9.3005
R669 VDD1.n47 VDD1.n46 9.3005
R670 VDD1.n130 VDD1.n129 9.3005
R671 VDD1.n69 VDD1.n68 9.3005
R672 VDD1.n124 VDD1.n123 9.3005
R673 VDD1.n122 VDD1.n121 9.3005
R674 VDD1.n73 VDD1.n72 9.3005
R675 VDD1.n116 VDD1.n115 9.3005
R676 VDD1.n114 VDD1.n113 9.3005
R677 VDD1.n90 VDD1.n89 9.3005
R678 VDD1.n85 VDD1.n84 9.3005
R679 VDD1.n96 VDD1.n95 9.3005
R680 VDD1.n98 VDD1.n97 9.3005
R681 VDD1.n81 VDD1.n80 9.3005
R682 VDD1.n104 VDD1.n103 9.3005
R683 VDD1.n106 VDD1.n105 9.3005
R684 VDD1.n107 VDD1.n76 9.3005
R685 VDD1.n61 VDD1.n2 8.92171
R686 VDD1.n29 VDD1.n28 8.92171
R687 VDD1.n95 VDD1.n94 8.92171
R688 VDD1.n128 VDD1.n69 8.92171
R689 VDD1.n62 VDD1.n0 8.14595
R690 VDD1.n25 VDD1.n19 8.14595
R691 VDD1.n91 VDD1.n85 8.14595
R692 VDD1.n129 VDD1.n67 8.14595
R693 VDD1.n24 VDD1.n21 7.3702
R694 VDD1.n90 VDD1.n87 7.3702
R695 VDD1.n64 VDD1.n0 5.81868
R696 VDD1.n25 VDD1.n24 5.81868
R697 VDD1.n91 VDD1.n90 5.81868
R698 VDD1.n131 VDD1.n67 5.81868
R699 VDD1.n62 VDD1.n61 5.04292
R700 VDD1.n28 VDD1.n19 5.04292
R701 VDD1.n94 VDD1.n85 5.04292
R702 VDD1.n129 VDD1.n128 5.04292
R703 VDD1.n58 VDD1.n2 4.26717
R704 VDD1.n29 VDD1.n17 4.26717
R705 VDD1.n95 VDD1.n83 4.26717
R706 VDD1.n125 VDD1.n69 4.26717
R707 VDD1.n57 VDD1.n4 3.49141
R708 VDD1.n33 VDD1.n32 3.49141
R709 VDD1.n99 VDD1.n98 3.49141
R710 VDD1.n124 VDD1.n71 3.49141
R711 VDD1.n54 VDD1.n53 2.71565
R712 VDD1.n36 VDD1.n15 2.71565
R713 VDD1.n102 VDD1.n81 2.71565
R714 VDD1.n121 VDD1.n120 2.71565
R715 VDD1.n136 VDD1.t8 2.70474
R716 VDD1.n136 VDD1.t3 2.70474
R717 VDD1.n65 VDD1.t1 2.70474
R718 VDD1.n65 VDD1.t2 2.70474
R719 VDD1.n134 VDD1.t5 2.70474
R720 VDD1.n134 VDD1.t9 2.70474
R721 VDD1.n132 VDD1.t7 2.70474
R722 VDD1.n132 VDD1.t0 2.70474
R723 VDD1.n23 VDD1.n22 2.41282
R724 VDD1.n89 VDD1.n88 2.41282
R725 VDD1.n50 VDD1.n6 1.93989
R726 VDD1.n37 VDD1.n13 1.93989
R727 VDD1.n103 VDD1.n79 1.93989
R728 VDD1.n117 VDD1.n73 1.93989
R729 VDD1 VDD1.n137 1.44231
R730 VDD1.n49 VDD1.n8 1.16414
R731 VDD1.n41 VDD1.n40 1.16414
R732 VDD1.n108 VDD1.n106 1.16414
R733 VDD1.n116 VDD1.n75 1.16414
R734 VDD1 VDD1.n66 0.55869
R735 VDD1.n135 VDD1.n133 0.445154
R736 VDD1.n46 VDD1.n45 0.388379
R737 VDD1.n12 VDD1.n10 0.388379
R738 VDD1.n107 VDD1.n77 0.388379
R739 VDD1.n113 VDD1.n112 0.388379
R740 VDD1.n63 VDD1.n1 0.155672
R741 VDD1.n56 VDD1.n1 0.155672
R742 VDD1.n56 VDD1.n55 0.155672
R743 VDD1.n55 VDD1.n5 0.155672
R744 VDD1.n48 VDD1.n5 0.155672
R745 VDD1.n48 VDD1.n47 0.155672
R746 VDD1.n47 VDD1.n9 0.155672
R747 VDD1.n39 VDD1.n9 0.155672
R748 VDD1.n39 VDD1.n38 0.155672
R749 VDD1.n38 VDD1.n14 0.155672
R750 VDD1.n31 VDD1.n14 0.155672
R751 VDD1.n31 VDD1.n30 0.155672
R752 VDD1.n30 VDD1.n18 0.155672
R753 VDD1.n23 VDD1.n18 0.155672
R754 VDD1.n89 VDD1.n84 0.155672
R755 VDD1.n96 VDD1.n84 0.155672
R756 VDD1.n97 VDD1.n96 0.155672
R757 VDD1.n97 VDD1.n80 0.155672
R758 VDD1.n104 VDD1.n80 0.155672
R759 VDD1.n105 VDD1.n104 0.155672
R760 VDD1.n105 VDD1.n76 0.155672
R761 VDD1.n114 VDD1.n76 0.155672
R762 VDD1.n115 VDD1.n114 0.155672
R763 VDD1.n115 VDD1.n72 0.155672
R764 VDD1.n122 VDD1.n72 0.155672
R765 VDD1.n123 VDD1.n122 0.155672
R766 VDD1.n123 VDD1.n68 0.155672
R767 VDD1.n130 VDD1.n68 0.155672
R768 B.n564 B.n77 585
R769 B.n566 B.n565 585
R770 B.n567 B.n76 585
R771 B.n569 B.n568 585
R772 B.n570 B.n75 585
R773 B.n572 B.n571 585
R774 B.n573 B.n74 585
R775 B.n575 B.n574 585
R776 B.n576 B.n73 585
R777 B.n578 B.n577 585
R778 B.n579 B.n72 585
R779 B.n581 B.n580 585
R780 B.n582 B.n71 585
R781 B.n584 B.n583 585
R782 B.n585 B.n70 585
R783 B.n587 B.n586 585
R784 B.n588 B.n69 585
R785 B.n590 B.n589 585
R786 B.n591 B.n68 585
R787 B.n593 B.n592 585
R788 B.n594 B.n67 585
R789 B.n596 B.n595 585
R790 B.n597 B.n66 585
R791 B.n599 B.n598 585
R792 B.n600 B.n65 585
R793 B.n602 B.n601 585
R794 B.n603 B.n64 585
R795 B.n605 B.n604 585
R796 B.n606 B.n63 585
R797 B.n608 B.n607 585
R798 B.n609 B.n62 585
R799 B.n611 B.n610 585
R800 B.n612 B.n61 585
R801 B.n614 B.n613 585
R802 B.n615 B.n60 585
R803 B.n617 B.n616 585
R804 B.n618 B.n59 585
R805 B.n620 B.n619 585
R806 B.n621 B.n58 585
R807 B.n623 B.n622 585
R808 B.n624 B.n57 585
R809 B.n626 B.n625 585
R810 B.n628 B.n627 585
R811 B.n629 B.n53 585
R812 B.n631 B.n630 585
R813 B.n632 B.n52 585
R814 B.n634 B.n633 585
R815 B.n635 B.n51 585
R816 B.n637 B.n636 585
R817 B.n638 B.n50 585
R818 B.n640 B.n639 585
R819 B.n642 B.n47 585
R820 B.n644 B.n643 585
R821 B.n645 B.n46 585
R822 B.n647 B.n646 585
R823 B.n648 B.n45 585
R824 B.n650 B.n649 585
R825 B.n651 B.n44 585
R826 B.n653 B.n652 585
R827 B.n654 B.n43 585
R828 B.n656 B.n655 585
R829 B.n657 B.n42 585
R830 B.n659 B.n658 585
R831 B.n660 B.n41 585
R832 B.n662 B.n661 585
R833 B.n663 B.n40 585
R834 B.n665 B.n664 585
R835 B.n666 B.n39 585
R836 B.n668 B.n667 585
R837 B.n669 B.n38 585
R838 B.n671 B.n670 585
R839 B.n672 B.n37 585
R840 B.n674 B.n673 585
R841 B.n675 B.n36 585
R842 B.n677 B.n676 585
R843 B.n678 B.n35 585
R844 B.n680 B.n679 585
R845 B.n681 B.n34 585
R846 B.n683 B.n682 585
R847 B.n684 B.n33 585
R848 B.n686 B.n685 585
R849 B.n687 B.n32 585
R850 B.n689 B.n688 585
R851 B.n690 B.n31 585
R852 B.n692 B.n691 585
R853 B.n693 B.n30 585
R854 B.n695 B.n694 585
R855 B.n696 B.n29 585
R856 B.n698 B.n697 585
R857 B.n699 B.n28 585
R858 B.n701 B.n700 585
R859 B.n702 B.n27 585
R860 B.n704 B.n703 585
R861 B.n563 B.n562 585
R862 B.n561 B.n78 585
R863 B.n560 B.n559 585
R864 B.n558 B.n79 585
R865 B.n557 B.n556 585
R866 B.n555 B.n80 585
R867 B.n554 B.n553 585
R868 B.n552 B.n81 585
R869 B.n551 B.n550 585
R870 B.n549 B.n82 585
R871 B.n548 B.n547 585
R872 B.n546 B.n83 585
R873 B.n545 B.n544 585
R874 B.n543 B.n84 585
R875 B.n542 B.n541 585
R876 B.n540 B.n85 585
R877 B.n539 B.n538 585
R878 B.n537 B.n86 585
R879 B.n536 B.n535 585
R880 B.n534 B.n87 585
R881 B.n533 B.n532 585
R882 B.n531 B.n88 585
R883 B.n530 B.n529 585
R884 B.n528 B.n89 585
R885 B.n527 B.n526 585
R886 B.n525 B.n90 585
R887 B.n524 B.n523 585
R888 B.n522 B.n91 585
R889 B.n521 B.n520 585
R890 B.n519 B.n92 585
R891 B.n518 B.n517 585
R892 B.n516 B.n93 585
R893 B.n515 B.n514 585
R894 B.n513 B.n94 585
R895 B.n512 B.n511 585
R896 B.n510 B.n95 585
R897 B.n509 B.n508 585
R898 B.n507 B.n96 585
R899 B.n506 B.n505 585
R900 B.n504 B.n97 585
R901 B.n503 B.n502 585
R902 B.n501 B.n98 585
R903 B.n500 B.n499 585
R904 B.n498 B.n99 585
R905 B.n497 B.n496 585
R906 B.n495 B.n100 585
R907 B.n494 B.n493 585
R908 B.n492 B.n101 585
R909 B.n491 B.n490 585
R910 B.n489 B.n102 585
R911 B.n488 B.n487 585
R912 B.n486 B.n103 585
R913 B.n485 B.n484 585
R914 B.n483 B.n104 585
R915 B.n482 B.n481 585
R916 B.n480 B.n105 585
R917 B.n479 B.n478 585
R918 B.n477 B.n106 585
R919 B.n476 B.n475 585
R920 B.n474 B.n107 585
R921 B.n473 B.n472 585
R922 B.n471 B.n108 585
R923 B.n470 B.n469 585
R924 B.n468 B.n109 585
R925 B.n467 B.n466 585
R926 B.n465 B.n110 585
R927 B.n464 B.n463 585
R928 B.n462 B.n111 585
R929 B.n461 B.n460 585
R930 B.n459 B.n112 585
R931 B.n458 B.n457 585
R932 B.n456 B.n113 585
R933 B.n455 B.n454 585
R934 B.n453 B.n114 585
R935 B.n452 B.n451 585
R936 B.n450 B.n115 585
R937 B.n449 B.n448 585
R938 B.n447 B.n116 585
R939 B.n446 B.n445 585
R940 B.n444 B.n117 585
R941 B.n443 B.n442 585
R942 B.n441 B.n118 585
R943 B.n440 B.n439 585
R944 B.n438 B.n119 585
R945 B.n437 B.n436 585
R946 B.n435 B.n120 585
R947 B.n434 B.n433 585
R948 B.n432 B.n121 585
R949 B.n431 B.n430 585
R950 B.n429 B.n122 585
R951 B.n428 B.n427 585
R952 B.n426 B.n123 585
R953 B.n425 B.n424 585
R954 B.n423 B.n124 585
R955 B.n422 B.n421 585
R956 B.n420 B.n125 585
R957 B.n419 B.n418 585
R958 B.n417 B.n126 585
R959 B.n416 B.n415 585
R960 B.n275 B.n274 585
R961 B.n276 B.n177 585
R962 B.n278 B.n277 585
R963 B.n279 B.n176 585
R964 B.n281 B.n280 585
R965 B.n282 B.n175 585
R966 B.n284 B.n283 585
R967 B.n285 B.n174 585
R968 B.n287 B.n286 585
R969 B.n288 B.n173 585
R970 B.n290 B.n289 585
R971 B.n291 B.n172 585
R972 B.n293 B.n292 585
R973 B.n294 B.n171 585
R974 B.n296 B.n295 585
R975 B.n297 B.n170 585
R976 B.n299 B.n298 585
R977 B.n300 B.n169 585
R978 B.n302 B.n301 585
R979 B.n303 B.n168 585
R980 B.n305 B.n304 585
R981 B.n306 B.n167 585
R982 B.n308 B.n307 585
R983 B.n309 B.n166 585
R984 B.n311 B.n310 585
R985 B.n312 B.n165 585
R986 B.n314 B.n313 585
R987 B.n315 B.n164 585
R988 B.n317 B.n316 585
R989 B.n318 B.n163 585
R990 B.n320 B.n319 585
R991 B.n321 B.n162 585
R992 B.n323 B.n322 585
R993 B.n324 B.n161 585
R994 B.n326 B.n325 585
R995 B.n327 B.n160 585
R996 B.n329 B.n328 585
R997 B.n330 B.n159 585
R998 B.n332 B.n331 585
R999 B.n333 B.n158 585
R1000 B.n335 B.n334 585
R1001 B.n336 B.n155 585
R1002 B.n339 B.n338 585
R1003 B.n340 B.n154 585
R1004 B.n342 B.n341 585
R1005 B.n343 B.n153 585
R1006 B.n345 B.n344 585
R1007 B.n346 B.n152 585
R1008 B.n348 B.n347 585
R1009 B.n349 B.n151 585
R1010 B.n351 B.n350 585
R1011 B.n353 B.n352 585
R1012 B.n354 B.n147 585
R1013 B.n356 B.n355 585
R1014 B.n357 B.n146 585
R1015 B.n359 B.n358 585
R1016 B.n360 B.n145 585
R1017 B.n362 B.n361 585
R1018 B.n363 B.n144 585
R1019 B.n365 B.n364 585
R1020 B.n366 B.n143 585
R1021 B.n368 B.n367 585
R1022 B.n369 B.n142 585
R1023 B.n371 B.n370 585
R1024 B.n372 B.n141 585
R1025 B.n374 B.n373 585
R1026 B.n375 B.n140 585
R1027 B.n377 B.n376 585
R1028 B.n378 B.n139 585
R1029 B.n380 B.n379 585
R1030 B.n381 B.n138 585
R1031 B.n383 B.n382 585
R1032 B.n384 B.n137 585
R1033 B.n386 B.n385 585
R1034 B.n387 B.n136 585
R1035 B.n389 B.n388 585
R1036 B.n390 B.n135 585
R1037 B.n392 B.n391 585
R1038 B.n393 B.n134 585
R1039 B.n395 B.n394 585
R1040 B.n396 B.n133 585
R1041 B.n398 B.n397 585
R1042 B.n399 B.n132 585
R1043 B.n401 B.n400 585
R1044 B.n402 B.n131 585
R1045 B.n404 B.n403 585
R1046 B.n405 B.n130 585
R1047 B.n407 B.n406 585
R1048 B.n408 B.n129 585
R1049 B.n410 B.n409 585
R1050 B.n411 B.n128 585
R1051 B.n413 B.n412 585
R1052 B.n414 B.n127 585
R1053 B.n273 B.n178 585
R1054 B.n272 B.n271 585
R1055 B.n270 B.n179 585
R1056 B.n269 B.n268 585
R1057 B.n267 B.n180 585
R1058 B.n266 B.n265 585
R1059 B.n264 B.n181 585
R1060 B.n263 B.n262 585
R1061 B.n261 B.n182 585
R1062 B.n260 B.n259 585
R1063 B.n258 B.n183 585
R1064 B.n257 B.n256 585
R1065 B.n255 B.n184 585
R1066 B.n254 B.n253 585
R1067 B.n252 B.n185 585
R1068 B.n251 B.n250 585
R1069 B.n249 B.n186 585
R1070 B.n248 B.n247 585
R1071 B.n246 B.n187 585
R1072 B.n245 B.n244 585
R1073 B.n243 B.n188 585
R1074 B.n242 B.n241 585
R1075 B.n240 B.n189 585
R1076 B.n239 B.n238 585
R1077 B.n237 B.n190 585
R1078 B.n236 B.n235 585
R1079 B.n234 B.n191 585
R1080 B.n233 B.n232 585
R1081 B.n231 B.n192 585
R1082 B.n230 B.n229 585
R1083 B.n228 B.n193 585
R1084 B.n227 B.n226 585
R1085 B.n225 B.n194 585
R1086 B.n224 B.n223 585
R1087 B.n222 B.n195 585
R1088 B.n221 B.n220 585
R1089 B.n219 B.n196 585
R1090 B.n218 B.n217 585
R1091 B.n216 B.n197 585
R1092 B.n215 B.n214 585
R1093 B.n213 B.n198 585
R1094 B.n212 B.n211 585
R1095 B.n210 B.n199 585
R1096 B.n209 B.n208 585
R1097 B.n207 B.n200 585
R1098 B.n206 B.n205 585
R1099 B.n204 B.n201 585
R1100 B.n203 B.n202 585
R1101 B.n2 B.n0 585
R1102 B.n777 B.n1 585
R1103 B.n776 B.n775 585
R1104 B.n774 B.n3 585
R1105 B.n773 B.n772 585
R1106 B.n771 B.n4 585
R1107 B.n770 B.n769 585
R1108 B.n768 B.n5 585
R1109 B.n767 B.n766 585
R1110 B.n765 B.n6 585
R1111 B.n764 B.n763 585
R1112 B.n762 B.n7 585
R1113 B.n761 B.n760 585
R1114 B.n759 B.n8 585
R1115 B.n758 B.n757 585
R1116 B.n756 B.n9 585
R1117 B.n755 B.n754 585
R1118 B.n753 B.n10 585
R1119 B.n752 B.n751 585
R1120 B.n750 B.n11 585
R1121 B.n749 B.n748 585
R1122 B.n747 B.n12 585
R1123 B.n746 B.n745 585
R1124 B.n744 B.n13 585
R1125 B.n743 B.n742 585
R1126 B.n741 B.n14 585
R1127 B.n740 B.n739 585
R1128 B.n738 B.n15 585
R1129 B.n737 B.n736 585
R1130 B.n735 B.n16 585
R1131 B.n734 B.n733 585
R1132 B.n732 B.n17 585
R1133 B.n731 B.n730 585
R1134 B.n729 B.n18 585
R1135 B.n728 B.n727 585
R1136 B.n726 B.n19 585
R1137 B.n725 B.n724 585
R1138 B.n723 B.n20 585
R1139 B.n722 B.n721 585
R1140 B.n720 B.n21 585
R1141 B.n719 B.n718 585
R1142 B.n717 B.n22 585
R1143 B.n716 B.n715 585
R1144 B.n714 B.n23 585
R1145 B.n713 B.n712 585
R1146 B.n711 B.n24 585
R1147 B.n710 B.n709 585
R1148 B.n708 B.n25 585
R1149 B.n707 B.n706 585
R1150 B.n705 B.n26 585
R1151 B.n779 B.n778 585
R1152 B.n274 B.n273 502.111
R1153 B.n705 B.n704 502.111
R1154 B.n416 B.n127 502.111
R1155 B.n562 B.n77 502.111
R1156 B.n148 B.t11 420.911
R1157 B.n54 B.t1 420.911
R1158 B.n156 B.t5 420.911
R1159 B.n48 B.t7 420.911
R1160 B.n149 B.t10 375.918
R1161 B.n55 B.t2 375.918
R1162 B.n157 B.t4 375.918
R1163 B.n49 B.t8 375.918
R1164 B.n148 B.t9 352.464
R1165 B.n156 B.t3 352.464
R1166 B.n48 B.t6 352.464
R1167 B.n54 B.t0 352.464
R1168 B.n273 B.n272 163.367
R1169 B.n272 B.n179 163.367
R1170 B.n268 B.n179 163.367
R1171 B.n268 B.n267 163.367
R1172 B.n267 B.n266 163.367
R1173 B.n266 B.n181 163.367
R1174 B.n262 B.n181 163.367
R1175 B.n262 B.n261 163.367
R1176 B.n261 B.n260 163.367
R1177 B.n260 B.n183 163.367
R1178 B.n256 B.n183 163.367
R1179 B.n256 B.n255 163.367
R1180 B.n255 B.n254 163.367
R1181 B.n254 B.n185 163.367
R1182 B.n250 B.n185 163.367
R1183 B.n250 B.n249 163.367
R1184 B.n249 B.n248 163.367
R1185 B.n248 B.n187 163.367
R1186 B.n244 B.n187 163.367
R1187 B.n244 B.n243 163.367
R1188 B.n243 B.n242 163.367
R1189 B.n242 B.n189 163.367
R1190 B.n238 B.n189 163.367
R1191 B.n238 B.n237 163.367
R1192 B.n237 B.n236 163.367
R1193 B.n236 B.n191 163.367
R1194 B.n232 B.n191 163.367
R1195 B.n232 B.n231 163.367
R1196 B.n231 B.n230 163.367
R1197 B.n230 B.n193 163.367
R1198 B.n226 B.n193 163.367
R1199 B.n226 B.n225 163.367
R1200 B.n225 B.n224 163.367
R1201 B.n224 B.n195 163.367
R1202 B.n220 B.n195 163.367
R1203 B.n220 B.n219 163.367
R1204 B.n219 B.n218 163.367
R1205 B.n218 B.n197 163.367
R1206 B.n214 B.n197 163.367
R1207 B.n214 B.n213 163.367
R1208 B.n213 B.n212 163.367
R1209 B.n212 B.n199 163.367
R1210 B.n208 B.n199 163.367
R1211 B.n208 B.n207 163.367
R1212 B.n207 B.n206 163.367
R1213 B.n206 B.n201 163.367
R1214 B.n202 B.n201 163.367
R1215 B.n202 B.n2 163.367
R1216 B.n778 B.n2 163.367
R1217 B.n778 B.n777 163.367
R1218 B.n777 B.n776 163.367
R1219 B.n776 B.n3 163.367
R1220 B.n772 B.n3 163.367
R1221 B.n772 B.n771 163.367
R1222 B.n771 B.n770 163.367
R1223 B.n770 B.n5 163.367
R1224 B.n766 B.n5 163.367
R1225 B.n766 B.n765 163.367
R1226 B.n765 B.n764 163.367
R1227 B.n764 B.n7 163.367
R1228 B.n760 B.n7 163.367
R1229 B.n760 B.n759 163.367
R1230 B.n759 B.n758 163.367
R1231 B.n758 B.n9 163.367
R1232 B.n754 B.n9 163.367
R1233 B.n754 B.n753 163.367
R1234 B.n753 B.n752 163.367
R1235 B.n752 B.n11 163.367
R1236 B.n748 B.n11 163.367
R1237 B.n748 B.n747 163.367
R1238 B.n747 B.n746 163.367
R1239 B.n746 B.n13 163.367
R1240 B.n742 B.n13 163.367
R1241 B.n742 B.n741 163.367
R1242 B.n741 B.n740 163.367
R1243 B.n740 B.n15 163.367
R1244 B.n736 B.n15 163.367
R1245 B.n736 B.n735 163.367
R1246 B.n735 B.n734 163.367
R1247 B.n734 B.n17 163.367
R1248 B.n730 B.n17 163.367
R1249 B.n730 B.n729 163.367
R1250 B.n729 B.n728 163.367
R1251 B.n728 B.n19 163.367
R1252 B.n724 B.n19 163.367
R1253 B.n724 B.n723 163.367
R1254 B.n723 B.n722 163.367
R1255 B.n722 B.n21 163.367
R1256 B.n718 B.n21 163.367
R1257 B.n718 B.n717 163.367
R1258 B.n717 B.n716 163.367
R1259 B.n716 B.n23 163.367
R1260 B.n712 B.n23 163.367
R1261 B.n712 B.n711 163.367
R1262 B.n711 B.n710 163.367
R1263 B.n710 B.n25 163.367
R1264 B.n706 B.n25 163.367
R1265 B.n706 B.n705 163.367
R1266 B.n274 B.n177 163.367
R1267 B.n278 B.n177 163.367
R1268 B.n279 B.n278 163.367
R1269 B.n280 B.n279 163.367
R1270 B.n280 B.n175 163.367
R1271 B.n284 B.n175 163.367
R1272 B.n285 B.n284 163.367
R1273 B.n286 B.n285 163.367
R1274 B.n286 B.n173 163.367
R1275 B.n290 B.n173 163.367
R1276 B.n291 B.n290 163.367
R1277 B.n292 B.n291 163.367
R1278 B.n292 B.n171 163.367
R1279 B.n296 B.n171 163.367
R1280 B.n297 B.n296 163.367
R1281 B.n298 B.n297 163.367
R1282 B.n298 B.n169 163.367
R1283 B.n302 B.n169 163.367
R1284 B.n303 B.n302 163.367
R1285 B.n304 B.n303 163.367
R1286 B.n304 B.n167 163.367
R1287 B.n308 B.n167 163.367
R1288 B.n309 B.n308 163.367
R1289 B.n310 B.n309 163.367
R1290 B.n310 B.n165 163.367
R1291 B.n314 B.n165 163.367
R1292 B.n315 B.n314 163.367
R1293 B.n316 B.n315 163.367
R1294 B.n316 B.n163 163.367
R1295 B.n320 B.n163 163.367
R1296 B.n321 B.n320 163.367
R1297 B.n322 B.n321 163.367
R1298 B.n322 B.n161 163.367
R1299 B.n326 B.n161 163.367
R1300 B.n327 B.n326 163.367
R1301 B.n328 B.n327 163.367
R1302 B.n328 B.n159 163.367
R1303 B.n332 B.n159 163.367
R1304 B.n333 B.n332 163.367
R1305 B.n334 B.n333 163.367
R1306 B.n334 B.n155 163.367
R1307 B.n339 B.n155 163.367
R1308 B.n340 B.n339 163.367
R1309 B.n341 B.n340 163.367
R1310 B.n341 B.n153 163.367
R1311 B.n345 B.n153 163.367
R1312 B.n346 B.n345 163.367
R1313 B.n347 B.n346 163.367
R1314 B.n347 B.n151 163.367
R1315 B.n351 B.n151 163.367
R1316 B.n352 B.n351 163.367
R1317 B.n352 B.n147 163.367
R1318 B.n356 B.n147 163.367
R1319 B.n357 B.n356 163.367
R1320 B.n358 B.n357 163.367
R1321 B.n358 B.n145 163.367
R1322 B.n362 B.n145 163.367
R1323 B.n363 B.n362 163.367
R1324 B.n364 B.n363 163.367
R1325 B.n364 B.n143 163.367
R1326 B.n368 B.n143 163.367
R1327 B.n369 B.n368 163.367
R1328 B.n370 B.n369 163.367
R1329 B.n370 B.n141 163.367
R1330 B.n374 B.n141 163.367
R1331 B.n375 B.n374 163.367
R1332 B.n376 B.n375 163.367
R1333 B.n376 B.n139 163.367
R1334 B.n380 B.n139 163.367
R1335 B.n381 B.n380 163.367
R1336 B.n382 B.n381 163.367
R1337 B.n382 B.n137 163.367
R1338 B.n386 B.n137 163.367
R1339 B.n387 B.n386 163.367
R1340 B.n388 B.n387 163.367
R1341 B.n388 B.n135 163.367
R1342 B.n392 B.n135 163.367
R1343 B.n393 B.n392 163.367
R1344 B.n394 B.n393 163.367
R1345 B.n394 B.n133 163.367
R1346 B.n398 B.n133 163.367
R1347 B.n399 B.n398 163.367
R1348 B.n400 B.n399 163.367
R1349 B.n400 B.n131 163.367
R1350 B.n404 B.n131 163.367
R1351 B.n405 B.n404 163.367
R1352 B.n406 B.n405 163.367
R1353 B.n406 B.n129 163.367
R1354 B.n410 B.n129 163.367
R1355 B.n411 B.n410 163.367
R1356 B.n412 B.n411 163.367
R1357 B.n412 B.n127 163.367
R1358 B.n417 B.n416 163.367
R1359 B.n418 B.n417 163.367
R1360 B.n418 B.n125 163.367
R1361 B.n422 B.n125 163.367
R1362 B.n423 B.n422 163.367
R1363 B.n424 B.n423 163.367
R1364 B.n424 B.n123 163.367
R1365 B.n428 B.n123 163.367
R1366 B.n429 B.n428 163.367
R1367 B.n430 B.n429 163.367
R1368 B.n430 B.n121 163.367
R1369 B.n434 B.n121 163.367
R1370 B.n435 B.n434 163.367
R1371 B.n436 B.n435 163.367
R1372 B.n436 B.n119 163.367
R1373 B.n440 B.n119 163.367
R1374 B.n441 B.n440 163.367
R1375 B.n442 B.n441 163.367
R1376 B.n442 B.n117 163.367
R1377 B.n446 B.n117 163.367
R1378 B.n447 B.n446 163.367
R1379 B.n448 B.n447 163.367
R1380 B.n448 B.n115 163.367
R1381 B.n452 B.n115 163.367
R1382 B.n453 B.n452 163.367
R1383 B.n454 B.n453 163.367
R1384 B.n454 B.n113 163.367
R1385 B.n458 B.n113 163.367
R1386 B.n459 B.n458 163.367
R1387 B.n460 B.n459 163.367
R1388 B.n460 B.n111 163.367
R1389 B.n464 B.n111 163.367
R1390 B.n465 B.n464 163.367
R1391 B.n466 B.n465 163.367
R1392 B.n466 B.n109 163.367
R1393 B.n470 B.n109 163.367
R1394 B.n471 B.n470 163.367
R1395 B.n472 B.n471 163.367
R1396 B.n472 B.n107 163.367
R1397 B.n476 B.n107 163.367
R1398 B.n477 B.n476 163.367
R1399 B.n478 B.n477 163.367
R1400 B.n478 B.n105 163.367
R1401 B.n482 B.n105 163.367
R1402 B.n483 B.n482 163.367
R1403 B.n484 B.n483 163.367
R1404 B.n484 B.n103 163.367
R1405 B.n488 B.n103 163.367
R1406 B.n489 B.n488 163.367
R1407 B.n490 B.n489 163.367
R1408 B.n490 B.n101 163.367
R1409 B.n494 B.n101 163.367
R1410 B.n495 B.n494 163.367
R1411 B.n496 B.n495 163.367
R1412 B.n496 B.n99 163.367
R1413 B.n500 B.n99 163.367
R1414 B.n501 B.n500 163.367
R1415 B.n502 B.n501 163.367
R1416 B.n502 B.n97 163.367
R1417 B.n506 B.n97 163.367
R1418 B.n507 B.n506 163.367
R1419 B.n508 B.n507 163.367
R1420 B.n508 B.n95 163.367
R1421 B.n512 B.n95 163.367
R1422 B.n513 B.n512 163.367
R1423 B.n514 B.n513 163.367
R1424 B.n514 B.n93 163.367
R1425 B.n518 B.n93 163.367
R1426 B.n519 B.n518 163.367
R1427 B.n520 B.n519 163.367
R1428 B.n520 B.n91 163.367
R1429 B.n524 B.n91 163.367
R1430 B.n525 B.n524 163.367
R1431 B.n526 B.n525 163.367
R1432 B.n526 B.n89 163.367
R1433 B.n530 B.n89 163.367
R1434 B.n531 B.n530 163.367
R1435 B.n532 B.n531 163.367
R1436 B.n532 B.n87 163.367
R1437 B.n536 B.n87 163.367
R1438 B.n537 B.n536 163.367
R1439 B.n538 B.n537 163.367
R1440 B.n538 B.n85 163.367
R1441 B.n542 B.n85 163.367
R1442 B.n543 B.n542 163.367
R1443 B.n544 B.n543 163.367
R1444 B.n544 B.n83 163.367
R1445 B.n548 B.n83 163.367
R1446 B.n549 B.n548 163.367
R1447 B.n550 B.n549 163.367
R1448 B.n550 B.n81 163.367
R1449 B.n554 B.n81 163.367
R1450 B.n555 B.n554 163.367
R1451 B.n556 B.n555 163.367
R1452 B.n556 B.n79 163.367
R1453 B.n560 B.n79 163.367
R1454 B.n561 B.n560 163.367
R1455 B.n562 B.n561 163.367
R1456 B.n704 B.n27 163.367
R1457 B.n700 B.n27 163.367
R1458 B.n700 B.n699 163.367
R1459 B.n699 B.n698 163.367
R1460 B.n698 B.n29 163.367
R1461 B.n694 B.n29 163.367
R1462 B.n694 B.n693 163.367
R1463 B.n693 B.n692 163.367
R1464 B.n692 B.n31 163.367
R1465 B.n688 B.n31 163.367
R1466 B.n688 B.n687 163.367
R1467 B.n687 B.n686 163.367
R1468 B.n686 B.n33 163.367
R1469 B.n682 B.n33 163.367
R1470 B.n682 B.n681 163.367
R1471 B.n681 B.n680 163.367
R1472 B.n680 B.n35 163.367
R1473 B.n676 B.n35 163.367
R1474 B.n676 B.n675 163.367
R1475 B.n675 B.n674 163.367
R1476 B.n674 B.n37 163.367
R1477 B.n670 B.n37 163.367
R1478 B.n670 B.n669 163.367
R1479 B.n669 B.n668 163.367
R1480 B.n668 B.n39 163.367
R1481 B.n664 B.n39 163.367
R1482 B.n664 B.n663 163.367
R1483 B.n663 B.n662 163.367
R1484 B.n662 B.n41 163.367
R1485 B.n658 B.n41 163.367
R1486 B.n658 B.n657 163.367
R1487 B.n657 B.n656 163.367
R1488 B.n656 B.n43 163.367
R1489 B.n652 B.n43 163.367
R1490 B.n652 B.n651 163.367
R1491 B.n651 B.n650 163.367
R1492 B.n650 B.n45 163.367
R1493 B.n646 B.n45 163.367
R1494 B.n646 B.n645 163.367
R1495 B.n645 B.n644 163.367
R1496 B.n644 B.n47 163.367
R1497 B.n639 B.n47 163.367
R1498 B.n639 B.n638 163.367
R1499 B.n638 B.n637 163.367
R1500 B.n637 B.n51 163.367
R1501 B.n633 B.n51 163.367
R1502 B.n633 B.n632 163.367
R1503 B.n632 B.n631 163.367
R1504 B.n631 B.n53 163.367
R1505 B.n627 B.n53 163.367
R1506 B.n627 B.n626 163.367
R1507 B.n626 B.n57 163.367
R1508 B.n622 B.n57 163.367
R1509 B.n622 B.n621 163.367
R1510 B.n621 B.n620 163.367
R1511 B.n620 B.n59 163.367
R1512 B.n616 B.n59 163.367
R1513 B.n616 B.n615 163.367
R1514 B.n615 B.n614 163.367
R1515 B.n614 B.n61 163.367
R1516 B.n610 B.n61 163.367
R1517 B.n610 B.n609 163.367
R1518 B.n609 B.n608 163.367
R1519 B.n608 B.n63 163.367
R1520 B.n604 B.n63 163.367
R1521 B.n604 B.n603 163.367
R1522 B.n603 B.n602 163.367
R1523 B.n602 B.n65 163.367
R1524 B.n598 B.n65 163.367
R1525 B.n598 B.n597 163.367
R1526 B.n597 B.n596 163.367
R1527 B.n596 B.n67 163.367
R1528 B.n592 B.n67 163.367
R1529 B.n592 B.n591 163.367
R1530 B.n591 B.n590 163.367
R1531 B.n590 B.n69 163.367
R1532 B.n586 B.n69 163.367
R1533 B.n586 B.n585 163.367
R1534 B.n585 B.n584 163.367
R1535 B.n584 B.n71 163.367
R1536 B.n580 B.n71 163.367
R1537 B.n580 B.n579 163.367
R1538 B.n579 B.n578 163.367
R1539 B.n578 B.n73 163.367
R1540 B.n574 B.n73 163.367
R1541 B.n574 B.n573 163.367
R1542 B.n573 B.n572 163.367
R1543 B.n572 B.n75 163.367
R1544 B.n568 B.n75 163.367
R1545 B.n568 B.n567 163.367
R1546 B.n567 B.n566 163.367
R1547 B.n566 B.n77 163.367
R1548 B.n150 B.n149 59.5399
R1549 B.n337 B.n157 59.5399
R1550 B.n641 B.n49 59.5399
R1551 B.n56 B.n55 59.5399
R1552 B.n149 B.n148 44.9944
R1553 B.n157 B.n156 44.9944
R1554 B.n49 B.n48 44.9944
R1555 B.n55 B.n54 44.9944
R1556 B.n703 B.n26 32.6249
R1557 B.n564 B.n563 32.6249
R1558 B.n415 B.n414 32.6249
R1559 B.n275 B.n178 32.6249
R1560 B B.n779 18.0485
R1561 B.n703 B.n702 10.6151
R1562 B.n702 B.n701 10.6151
R1563 B.n701 B.n28 10.6151
R1564 B.n697 B.n28 10.6151
R1565 B.n697 B.n696 10.6151
R1566 B.n696 B.n695 10.6151
R1567 B.n695 B.n30 10.6151
R1568 B.n691 B.n30 10.6151
R1569 B.n691 B.n690 10.6151
R1570 B.n690 B.n689 10.6151
R1571 B.n689 B.n32 10.6151
R1572 B.n685 B.n32 10.6151
R1573 B.n685 B.n684 10.6151
R1574 B.n684 B.n683 10.6151
R1575 B.n683 B.n34 10.6151
R1576 B.n679 B.n34 10.6151
R1577 B.n679 B.n678 10.6151
R1578 B.n678 B.n677 10.6151
R1579 B.n677 B.n36 10.6151
R1580 B.n673 B.n36 10.6151
R1581 B.n673 B.n672 10.6151
R1582 B.n672 B.n671 10.6151
R1583 B.n671 B.n38 10.6151
R1584 B.n667 B.n38 10.6151
R1585 B.n667 B.n666 10.6151
R1586 B.n666 B.n665 10.6151
R1587 B.n665 B.n40 10.6151
R1588 B.n661 B.n40 10.6151
R1589 B.n661 B.n660 10.6151
R1590 B.n660 B.n659 10.6151
R1591 B.n659 B.n42 10.6151
R1592 B.n655 B.n42 10.6151
R1593 B.n655 B.n654 10.6151
R1594 B.n654 B.n653 10.6151
R1595 B.n653 B.n44 10.6151
R1596 B.n649 B.n44 10.6151
R1597 B.n649 B.n648 10.6151
R1598 B.n648 B.n647 10.6151
R1599 B.n647 B.n46 10.6151
R1600 B.n643 B.n46 10.6151
R1601 B.n643 B.n642 10.6151
R1602 B.n640 B.n50 10.6151
R1603 B.n636 B.n50 10.6151
R1604 B.n636 B.n635 10.6151
R1605 B.n635 B.n634 10.6151
R1606 B.n634 B.n52 10.6151
R1607 B.n630 B.n52 10.6151
R1608 B.n630 B.n629 10.6151
R1609 B.n629 B.n628 10.6151
R1610 B.n625 B.n624 10.6151
R1611 B.n624 B.n623 10.6151
R1612 B.n623 B.n58 10.6151
R1613 B.n619 B.n58 10.6151
R1614 B.n619 B.n618 10.6151
R1615 B.n618 B.n617 10.6151
R1616 B.n617 B.n60 10.6151
R1617 B.n613 B.n60 10.6151
R1618 B.n613 B.n612 10.6151
R1619 B.n612 B.n611 10.6151
R1620 B.n611 B.n62 10.6151
R1621 B.n607 B.n62 10.6151
R1622 B.n607 B.n606 10.6151
R1623 B.n606 B.n605 10.6151
R1624 B.n605 B.n64 10.6151
R1625 B.n601 B.n64 10.6151
R1626 B.n601 B.n600 10.6151
R1627 B.n600 B.n599 10.6151
R1628 B.n599 B.n66 10.6151
R1629 B.n595 B.n66 10.6151
R1630 B.n595 B.n594 10.6151
R1631 B.n594 B.n593 10.6151
R1632 B.n593 B.n68 10.6151
R1633 B.n589 B.n68 10.6151
R1634 B.n589 B.n588 10.6151
R1635 B.n588 B.n587 10.6151
R1636 B.n587 B.n70 10.6151
R1637 B.n583 B.n70 10.6151
R1638 B.n583 B.n582 10.6151
R1639 B.n582 B.n581 10.6151
R1640 B.n581 B.n72 10.6151
R1641 B.n577 B.n72 10.6151
R1642 B.n577 B.n576 10.6151
R1643 B.n576 B.n575 10.6151
R1644 B.n575 B.n74 10.6151
R1645 B.n571 B.n74 10.6151
R1646 B.n571 B.n570 10.6151
R1647 B.n570 B.n569 10.6151
R1648 B.n569 B.n76 10.6151
R1649 B.n565 B.n76 10.6151
R1650 B.n565 B.n564 10.6151
R1651 B.n415 B.n126 10.6151
R1652 B.n419 B.n126 10.6151
R1653 B.n420 B.n419 10.6151
R1654 B.n421 B.n420 10.6151
R1655 B.n421 B.n124 10.6151
R1656 B.n425 B.n124 10.6151
R1657 B.n426 B.n425 10.6151
R1658 B.n427 B.n426 10.6151
R1659 B.n427 B.n122 10.6151
R1660 B.n431 B.n122 10.6151
R1661 B.n432 B.n431 10.6151
R1662 B.n433 B.n432 10.6151
R1663 B.n433 B.n120 10.6151
R1664 B.n437 B.n120 10.6151
R1665 B.n438 B.n437 10.6151
R1666 B.n439 B.n438 10.6151
R1667 B.n439 B.n118 10.6151
R1668 B.n443 B.n118 10.6151
R1669 B.n444 B.n443 10.6151
R1670 B.n445 B.n444 10.6151
R1671 B.n445 B.n116 10.6151
R1672 B.n449 B.n116 10.6151
R1673 B.n450 B.n449 10.6151
R1674 B.n451 B.n450 10.6151
R1675 B.n451 B.n114 10.6151
R1676 B.n455 B.n114 10.6151
R1677 B.n456 B.n455 10.6151
R1678 B.n457 B.n456 10.6151
R1679 B.n457 B.n112 10.6151
R1680 B.n461 B.n112 10.6151
R1681 B.n462 B.n461 10.6151
R1682 B.n463 B.n462 10.6151
R1683 B.n463 B.n110 10.6151
R1684 B.n467 B.n110 10.6151
R1685 B.n468 B.n467 10.6151
R1686 B.n469 B.n468 10.6151
R1687 B.n469 B.n108 10.6151
R1688 B.n473 B.n108 10.6151
R1689 B.n474 B.n473 10.6151
R1690 B.n475 B.n474 10.6151
R1691 B.n475 B.n106 10.6151
R1692 B.n479 B.n106 10.6151
R1693 B.n480 B.n479 10.6151
R1694 B.n481 B.n480 10.6151
R1695 B.n481 B.n104 10.6151
R1696 B.n485 B.n104 10.6151
R1697 B.n486 B.n485 10.6151
R1698 B.n487 B.n486 10.6151
R1699 B.n487 B.n102 10.6151
R1700 B.n491 B.n102 10.6151
R1701 B.n492 B.n491 10.6151
R1702 B.n493 B.n492 10.6151
R1703 B.n493 B.n100 10.6151
R1704 B.n497 B.n100 10.6151
R1705 B.n498 B.n497 10.6151
R1706 B.n499 B.n498 10.6151
R1707 B.n499 B.n98 10.6151
R1708 B.n503 B.n98 10.6151
R1709 B.n504 B.n503 10.6151
R1710 B.n505 B.n504 10.6151
R1711 B.n505 B.n96 10.6151
R1712 B.n509 B.n96 10.6151
R1713 B.n510 B.n509 10.6151
R1714 B.n511 B.n510 10.6151
R1715 B.n511 B.n94 10.6151
R1716 B.n515 B.n94 10.6151
R1717 B.n516 B.n515 10.6151
R1718 B.n517 B.n516 10.6151
R1719 B.n517 B.n92 10.6151
R1720 B.n521 B.n92 10.6151
R1721 B.n522 B.n521 10.6151
R1722 B.n523 B.n522 10.6151
R1723 B.n523 B.n90 10.6151
R1724 B.n527 B.n90 10.6151
R1725 B.n528 B.n527 10.6151
R1726 B.n529 B.n528 10.6151
R1727 B.n529 B.n88 10.6151
R1728 B.n533 B.n88 10.6151
R1729 B.n534 B.n533 10.6151
R1730 B.n535 B.n534 10.6151
R1731 B.n535 B.n86 10.6151
R1732 B.n539 B.n86 10.6151
R1733 B.n540 B.n539 10.6151
R1734 B.n541 B.n540 10.6151
R1735 B.n541 B.n84 10.6151
R1736 B.n545 B.n84 10.6151
R1737 B.n546 B.n545 10.6151
R1738 B.n547 B.n546 10.6151
R1739 B.n547 B.n82 10.6151
R1740 B.n551 B.n82 10.6151
R1741 B.n552 B.n551 10.6151
R1742 B.n553 B.n552 10.6151
R1743 B.n553 B.n80 10.6151
R1744 B.n557 B.n80 10.6151
R1745 B.n558 B.n557 10.6151
R1746 B.n559 B.n558 10.6151
R1747 B.n559 B.n78 10.6151
R1748 B.n563 B.n78 10.6151
R1749 B.n276 B.n275 10.6151
R1750 B.n277 B.n276 10.6151
R1751 B.n277 B.n176 10.6151
R1752 B.n281 B.n176 10.6151
R1753 B.n282 B.n281 10.6151
R1754 B.n283 B.n282 10.6151
R1755 B.n283 B.n174 10.6151
R1756 B.n287 B.n174 10.6151
R1757 B.n288 B.n287 10.6151
R1758 B.n289 B.n288 10.6151
R1759 B.n289 B.n172 10.6151
R1760 B.n293 B.n172 10.6151
R1761 B.n294 B.n293 10.6151
R1762 B.n295 B.n294 10.6151
R1763 B.n295 B.n170 10.6151
R1764 B.n299 B.n170 10.6151
R1765 B.n300 B.n299 10.6151
R1766 B.n301 B.n300 10.6151
R1767 B.n301 B.n168 10.6151
R1768 B.n305 B.n168 10.6151
R1769 B.n306 B.n305 10.6151
R1770 B.n307 B.n306 10.6151
R1771 B.n307 B.n166 10.6151
R1772 B.n311 B.n166 10.6151
R1773 B.n312 B.n311 10.6151
R1774 B.n313 B.n312 10.6151
R1775 B.n313 B.n164 10.6151
R1776 B.n317 B.n164 10.6151
R1777 B.n318 B.n317 10.6151
R1778 B.n319 B.n318 10.6151
R1779 B.n319 B.n162 10.6151
R1780 B.n323 B.n162 10.6151
R1781 B.n324 B.n323 10.6151
R1782 B.n325 B.n324 10.6151
R1783 B.n325 B.n160 10.6151
R1784 B.n329 B.n160 10.6151
R1785 B.n330 B.n329 10.6151
R1786 B.n331 B.n330 10.6151
R1787 B.n331 B.n158 10.6151
R1788 B.n335 B.n158 10.6151
R1789 B.n336 B.n335 10.6151
R1790 B.n338 B.n154 10.6151
R1791 B.n342 B.n154 10.6151
R1792 B.n343 B.n342 10.6151
R1793 B.n344 B.n343 10.6151
R1794 B.n344 B.n152 10.6151
R1795 B.n348 B.n152 10.6151
R1796 B.n349 B.n348 10.6151
R1797 B.n350 B.n349 10.6151
R1798 B.n354 B.n353 10.6151
R1799 B.n355 B.n354 10.6151
R1800 B.n355 B.n146 10.6151
R1801 B.n359 B.n146 10.6151
R1802 B.n360 B.n359 10.6151
R1803 B.n361 B.n360 10.6151
R1804 B.n361 B.n144 10.6151
R1805 B.n365 B.n144 10.6151
R1806 B.n366 B.n365 10.6151
R1807 B.n367 B.n366 10.6151
R1808 B.n367 B.n142 10.6151
R1809 B.n371 B.n142 10.6151
R1810 B.n372 B.n371 10.6151
R1811 B.n373 B.n372 10.6151
R1812 B.n373 B.n140 10.6151
R1813 B.n377 B.n140 10.6151
R1814 B.n378 B.n377 10.6151
R1815 B.n379 B.n378 10.6151
R1816 B.n379 B.n138 10.6151
R1817 B.n383 B.n138 10.6151
R1818 B.n384 B.n383 10.6151
R1819 B.n385 B.n384 10.6151
R1820 B.n385 B.n136 10.6151
R1821 B.n389 B.n136 10.6151
R1822 B.n390 B.n389 10.6151
R1823 B.n391 B.n390 10.6151
R1824 B.n391 B.n134 10.6151
R1825 B.n395 B.n134 10.6151
R1826 B.n396 B.n395 10.6151
R1827 B.n397 B.n396 10.6151
R1828 B.n397 B.n132 10.6151
R1829 B.n401 B.n132 10.6151
R1830 B.n402 B.n401 10.6151
R1831 B.n403 B.n402 10.6151
R1832 B.n403 B.n130 10.6151
R1833 B.n407 B.n130 10.6151
R1834 B.n408 B.n407 10.6151
R1835 B.n409 B.n408 10.6151
R1836 B.n409 B.n128 10.6151
R1837 B.n413 B.n128 10.6151
R1838 B.n414 B.n413 10.6151
R1839 B.n271 B.n178 10.6151
R1840 B.n271 B.n270 10.6151
R1841 B.n270 B.n269 10.6151
R1842 B.n269 B.n180 10.6151
R1843 B.n265 B.n180 10.6151
R1844 B.n265 B.n264 10.6151
R1845 B.n264 B.n263 10.6151
R1846 B.n263 B.n182 10.6151
R1847 B.n259 B.n182 10.6151
R1848 B.n259 B.n258 10.6151
R1849 B.n258 B.n257 10.6151
R1850 B.n257 B.n184 10.6151
R1851 B.n253 B.n184 10.6151
R1852 B.n253 B.n252 10.6151
R1853 B.n252 B.n251 10.6151
R1854 B.n251 B.n186 10.6151
R1855 B.n247 B.n186 10.6151
R1856 B.n247 B.n246 10.6151
R1857 B.n246 B.n245 10.6151
R1858 B.n245 B.n188 10.6151
R1859 B.n241 B.n188 10.6151
R1860 B.n241 B.n240 10.6151
R1861 B.n240 B.n239 10.6151
R1862 B.n239 B.n190 10.6151
R1863 B.n235 B.n190 10.6151
R1864 B.n235 B.n234 10.6151
R1865 B.n234 B.n233 10.6151
R1866 B.n233 B.n192 10.6151
R1867 B.n229 B.n192 10.6151
R1868 B.n229 B.n228 10.6151
R1869 B.n228 B.n227 10.6151
R1870 B.n227 B.n194 10.6151
R1871 B.n223 B.n194 10.6151
R1872 B.n223 B.n222 10.6151
R1873 B.n222 B.n221 10.6151
R1874 B.n221 B.n196 10.6151
R1875 B.n217 B.n196 10.6151
R1876 B.n217 B.n216 10.6151
R1877 B.n216 B.n215 10.6151
R1878 B.n215 B.n198 10.6151
R1879 B.n211 B.n198 10.6151
R1880 B.n211 B.n210 10.6151
R1881 B.n210 B.n209 10.6151
R1882 B.n209 B.n200 10.6151
R1883 B.n205 B.n200 10.6151
R1884 B.n205 B.n204 10.6151
R1885 B.n204 B.n203 10.6151
R1886 B.n203 B.n0 10.6151
R1887 B.n775 B.n1 10.6151
R1888 B.n775 B.n774 10.6151
R1889 B.n774 B.n773 10.6151
R1890 B.n773 B.n4 10.6151
R1891 B.n769 B.n4 10.6151
R1892 B.n769 B.n768 10.6151
R1893 B.n768 B.n767 10.6151
R1894 B.n767 B.n6 10.6151
R1895 B.n763 B.n6 10.6151
R1896 B.n763 B.n762 10.6151
R1897 B.n762 B.n761 10.6151
R1898 B.n761 B.n8 10.6151
R1899 B.n757 B.n8 10.6151
R1900 B.n757 B.n756 10.6151
R1901 B.n756 B.n755 10.6151
R1902 B.n755 B.n10 10.6151
R1903 B.n751 B.n10 10.6151
R1904 B.n751 B.n750 10.6151
R1905 B.n750 B.n749 10.6151
R1906 B.n749 B.n12 10.6151
R1907 B.n745 B.n12 10.6151
R1908 B.n745 B.n744 10.6151
R1909 B.n744 B.n743 10.6151
R1910 B.n743 B.n14 10.6151
R1911 B.n739 B.n14 10.6151
R1912 B.n739 B.n738 10.6151
R1913 B.n738 B.n737 10.6151
R1914 B.n737 B.n16 10.6151
R1915 B.n733 B.n16 10.6151
R1916 B.n733 B.n732 10.6151
R1917 B.n732 B.n731 10.6151
R1918 B.n731 B.n18 10.6151
R1919 B.n727 B.n18 10.6151
R1920 B.n727 B.n726 10.6151
R1921 B.n726 B.n725 10.6151
R1922 B.n725 B.n20 10.6151
R1923 B.n721 B.n20 10.6151
R1924 B.n721 B.n720 10.6151
R1925 B.n720 B.n719 10.6151
R1926 B.n719 B.n22 10.6151
R1927 B.n715 B.n22 10.6151
R1928 B.n715 B.n714 10.6151
R1929 B.n714 B.n713 10.6151
R1930 B.n713 B.n24 10.6151
R1931 B.n709 B.n24 10.6151
R1932 B.n709 B.n708 10.6151
R1933 B.n708 B.n707 10.6151
R1934 B.n707 B.n26 10.6151
R1935 B.n641 B.n640 6.5566
R1936 B.n628 B.n56 6.5566
R1937 B.n338 B.n337 6.5566
R1938 B.n350 B.n150 6.5566
R1939 B.n642 B.n641 4.05904
R1940 B.n625 B.n56 4.05904
R1941 B.n337 B.n336 4.05904
R1942 B.n353 B.n150 4.05904
R1943 B.n779 B.n0 2.81026
R1944 B.n779 B.n1 2.81026
R1945 VN.n8 VN.t4 175.816
R1946 VN.n42 VN.t0 175.816
R1947 VN.n65 VN.n34 161.3
R1948 VN.n64 VN.n63 161.3
R1949 VN.n62 VN.n35 161.3
R1950 VN.n61 VN.n60 161.3
R1951 VN.n58 VN.n36 161.3
R1952 VN.n57 VN.n56 161.3
R1953 VN.n55 VN.n37 161.3
R1954 VN.n54 VN.n53 161.3
R1955 VN.n52 VN.n38 161.3
R1956 VN.n50 VN.n49 161.3
R1957 VN.n48 VN.n39 161.3
R1958 VN.n47 VN.n46 161.3
R1959 VN.n45 VN.n40 161.3
R1960 VN.n44 VN.n43 161.3
R1961 VN.n31 VN.n0 161.3
R1962 VN.n30 VN.n29 161.3
R1963 VN.n28 VN.n1 161.3
R1964 VN.n27 VN.n26 161.3
R1965 VN.n24 VN.n2 161.3
R1966 VN.n23 VN.n22 161.3
R1967 VN.n21 VN.n3 161.3
R1968 VN.n20 VN.n19 161.3
R1969 VN.n18 VN.n4 161.3
R1970 VN.n16 VN.n15 161.3
R1971 VN.n14 VN.n5 161.3
R1972 VN.n13 VN.n12 161.3
R1973 VN.n11 VN.n6 161.3
R1974 VN.n10 VN.n9 161.3
R1975 VN.n7 VN.t7 145.57
R1976 VN.n17 VN.t5 145.57
R1977 VN.n25 VN.t9 145.57
R1978 VN.n32 VN.t3 145.57
R1979 VN.n41 VN.t1 145.57
R1980 VN.n51 VN.t2 145.57
R1981 VN.n59 VN.t8 145.57
R1982 VN.n66 VN.t6 145.57
R1983 VN.n33 VN.n32 91.7266
R1984 VN.n67 VN.n66 91.7266
R1985 VN.n8 VN.n7 66.4483
R1986 VN.n42 VN.n41 66.4483
R1987 VN.n30 VN.n1 56.5617
R1988 VN.n64 VN.n35 56.5617
R1989 VN VN.n67 50.1042
R1990 VN.n12 VN.n5 49.296
R1991 VN.n19 VN.n3 49.296
R1992 VN.n46 VN.n39 49.296
R1993 VN.n53 VN.n37 49.296
R1994 VN.n12 VN.n11 31.8581
R1995 VN.n23 VN.n3 31.8581
R1996 VN.n46 VN.n45 31.8581
R1997 VN.n57 VN.n37 31.8581
R1998 VN.n11 VN.n10 24.5923
R1999 VN.n16 VN.n5 24.5923
R2000 VN.n19 VN.n18 24.5923
R2001 VN.n24 VN.n23 24.5923
R2002 VN.n26 VN.n1 24.5923
R2003 VN.n31 VN.n30 24.5923
R2004 VN.n45 VN.n44 24.5923
R2005 VN.n53 VN.n52 24.5923
R2006 VN.n50 VN.n39 24.5923
R2007 VN.n60 VN.n35 24.5923
R2008 VN.n58 VN.n57 24.5923
R2009 VN.n65 VN.n64 24.5923
R2010 VN.n26 VN.n25 21.1495
R2011 VN.n60 VN.n59 21.1495
R2012 VN.n32 VN.n31 19.1821
R2013 VN.n66 VN.n65 19.1821
R2014 VN.n43 VN.n42 13.4112
R2015 VN.n9 VN.n8 13.4112
R2016 VN.n17 VN.n16 12.2964
R2017 VN.n18 VN.n17 12.2964
R2018 VN.n52 VN.n51 12.2964
R2019 VN.n51 VN.n50 12.2964
R2020 VN.n10 VN.n7 3.44336
R2021 VN.n25 VN.n24 3.44336
R2022 VN.n44 VN.n41 3.44336
R2023 VN.n59 VN.n58 3.44336
R2024 VN.n67 VN.n34 0.278335
R2025 VN.n33 VN.n0 0.278335
R2026 VN.n63 VN.n34 0.189894
R2027 VN.n63 VN.n62 0.189894
R2028 VN.n62 VN.n61 0.189894
R2029 VN.n61 VN.n36 0.189894
R2030 VN.n56 VN.n36 0.189894
R2031 VN.n56 VN.n55 0.189894
R2032 VN.n55 VN.n54 0.189894
R2033 VN.n54 VN.n38 0.189894
R2034 VN.n49 VN.n38 0.189894
R2035 VN.n49 VN.n48 0.189894
R2036 VN.n48 VN.n47 0.189894
R2037 VN.n47 VN.n40 0.189894
R2038 VN.n43 VN.n40 0.189894
R2039 VN.n9 VN.n6 0.189894
R2040 VN.n13 VN.n6 0.189894
R2041 VN.n14 VN.n13 0.189894
R2042 VN.n15 VN.n14 0.189894
R2043 VN.n15 VN.n4 0.189894
R2044 VN.n20 VN.n4 0.189894
R2045 VN.n21 VN.n20 0.189894
R2046 VN.n22 VN.n21 0.189894
R2047 VN.n22 VN.n2 0.189894
R2048 VN.n27 VN.n2 0.189894
R2049 VN.n28 VN.n27 0.189894
R2050 VN.n29 VN.n28 0.189894
R2051 VN.n29 VN.n0 0.189894
R2052 VN VN.n33 0.153485
R2053 VDD2.n129 VDD2.n69 756.745
R2054 VDD2.n60 VDD2.n0 756.745
R2055 VDD2.n130 VDD2.n129 585
R2056 VDD2.n128 VDD2.n127 585
R2057 VDD2.n73 VDD2.n72 585
R2058 VDD2.n122 VDD2.n121 585
R2059 VDD2.n120 VDD2.n119 585
R2060 VDD2.n77 VDD2.n76 585
R2061 VDD2.n114 VDD2.n113 585
R2062 VDD2.n112 VDD2.n79 585
R2063 VDD2.n111 VDD2.n110 585
R2064 VDD2.n82 VDD2.n80 585
R2065 VDD2.n105 VDD2.n104 585
R2066 VDD2.n103 VDD2.n102 585
R2067 VDD2.n86 VDD2.n85 585
R2068 VDD2.n97 VDD2.n96 585
R2069 VDD2.n95 VDD2.n94 585
R2070 VDD2.n90 VDD2.n89 585
R2071 VDD2.n20 VDD2.n19 585
R2072 VDD2.n25 VDD2.n24 585
R2073 VDD2.n27 VDD2.n26 585
R2074 VDD2.n16 VDD2.n15 585
R2075 VDD2.n33 VDD2.n32 585
R2076 VDD2.n35 VDD2.n34 585
R2077 VDD2.n12 VDD2.n11 585
R2078 VDD2.n42 VDD2.n41 585
R2079 VDD2.n43 VDD2.n10 585
R2080 VDD2.n45 VDD2.n44 585
R2081 VDD2.n8 VDD2.n7 585
R2082 VDD2.n51 VDD2.n50 585
R2083 VDD2.n53 VDD2.n52 585
R2084 VDD2.n4 VDD2.n3 585
R2085 VDD2.n59 VDD2.n58 585
R2086 VDD2.n61 VDD2.n60 585
R2087 VDD2.n91 VDD2.t3 329.036
R2088 VDD2.n21 VDD2.t5 329.036
R2089 VDD2.n129 VDD2.n128 171.744
R2090 VDD2.n128 VDD2.n72 171.744
R2091 VDD2.n121 VDD2.n72 171.744
R2092 VDD2.n121 VDD2.n120 171.744
R2093 VDD2.n120 VDD2.n76 171.744
R2094 VDD2.n113 VDD2.n76 171.744
R2095 VDD2.n113 VDD2.n112 171.744
R2096 VDD2.n112 VDD2.n111 171.744
R2097 VDD2.n111 VDD2.n80 171.744
R2098 VDD2.n104 VDD2.n80 171.744
R2099 VDD2.n104 VDD2.n103 171.744
R2100 VDD2.n103 VDD2.n85 171.744
R2101 VDD2.n96 VDD2.n85 171.744
R2102 VDD2.n96 VDD2.n95 171.744
R2103 VDD2.n95 VDD2.n89 171.744
R2104 VDD2.n25 VDD2.n19 171.744
R2105 VDD2.n26 VDD2.n25 171.744
R2106 VDD2.n26 VDD2.n15 171.744
R2107 VDD2.n33 VDD2.n15 171.744
R2108 VDD2.n34 VDD2.n33 171.744
R2109 VDD2.n34 VDD2.n11 171.744
R2110 VDD2.n42 VDD2.n11 171.744
R2111 VDD2.n43 VDD2.n42 171.744
R2112 VDD2.n44 VDD2.n43 171.744
R2113 VDD2.n44 VDD2.n7 171.744
R2114 VDD2.n51 VDD2.n7 171.744
R2115 VDD2.n52 VDD2.n51 171.744
R2116 VDD2.n52 VDD2.n3 171.744
R2117 VDD2.n59 VDD2.n3 171.744
R2118 VDD2.n60 VDD2.n59 171.744
R2119 VDD2.t3 VDD2.n89 85.8723
R2120 VDD2.t5 VDD2.n19 85.8723
R2121 VDD2.n68 VDD2.n67 73.3443
R2122 VDD2 VDD2.n137 73.3414
R2123 VDD2.n136 VDD2.n135 71.8998
R2124 VDD2.n66 VDD2.n65 71.8996
R2125 VDD2.n66 VDD2.n64 48.9247
R2126 VDD2.n134 VDD2.n133 46.9247
R2127 VDD2.n134 VDD2.n68 43.5774
R2128 VDD2.n114 VDD2.n79 13.1884
R2129 VDD2.n45 VDD2.n10 13.1884
R2130 VDD2.n115 VDD2.n77 12.8005
R2131 VDD2.n110 VDD2.n81 12.8005
R2132 VDD2.n41 VDD2.n40 12.8005
R2133 VDD2.n46 VDD2.n8 12.8005
R2134 VDD2.n119 VDD2.n118 12.0247
R2135 VDD2.n109 VDD2.n82 12.0247
R2136 VDD2.n39 VDD2.n12 12.0247
R2137 VDD2.n50 VDD2.n49 12.0247
R2138 VDD2.n122 VDD2.n75 11.249
R2139 VDD2.n106 VDD2.n105 11.249
R2140 VDD2.n36 VDD2.n35 11.249
R2141 VDD2.n53 VDD2.n6 11.249
R2142 VDD2.n91 VDD2.n90 10.7239
R2143 VDD2.n21 VDD2.n20 10.7239
R2144 VDD2.n123 VDD2.n73 10.4732
R2145 VDD2.n102 VDD2.n84 10.4732
R2146 VDD2.n32 VDD2.n14 10.4732
R2147 VDD2.n54 VDD2.n4 10.4732
R2148 VDD2.n127 VDD2.n126 9.69747
R2149 VDD2.n101 VDD2.n86 9.69747
R2150 VDD2.n31 VDD2.n16 9.69747
R2151 VDD2.n58 VDD2.n57 9.69747
R2152 VDD2.n133 VDD2.n132 9.45567
R2153 VDD2.n64 VDD2.n63 9.45567
R2154 VDD2.n93 VDD2.n92 9.3005
R2155 VDD2.n88 VDD2.n87 9.3005
R2156 VDD2.n99 VDD2.n98 9.3005
R2157 VDD2.n101 VDD2.n100 9.3005
R2158 VDD2.n84 VDD2.n83 9.3005
R2159 VDD2.n107 VDD2.n106 9.3005
R2160 VDD2.n109 VDD2.n108 9.3005
R2161 VDD2.n81 VDD2.n78 9.3005
R2162 VDD2.n132 VDD2.n131 9.3005
R2163 VDD2.n71 VDD2.n70 9.3005
R2164 VDD2.n126 VDD2.n125 9.3005
R2165 VDD2.n124 VDD2.n123 9.3005
R2166 VDD2.n75 VDD2.n74 9.3005
R2167 VDD2.n118 VDD2.n117 9.3005
R2168 VDD2.n116 VDD2.n115 9.3005
R2169 VDD2.n63 VDD2.n62 9.3005
R2170 VDD2.n2 VDD2.n1 9.3005
R2171 VDD2.n57 VDD2.n56 9.3005
R2172 VDD2.n55 VDD2.n54 9.3005
R2173 VDD2.n6 VDD2.n5 9.3005
R2174 VDD2.n49 VDD2.n48 9.3005
R2175 VDD2.n47 VDD2.n46 9.3005
R2176 VDD2.n23 VDD2.n22 9.3005
R2177 VDD2.n18 VDD2.n17 9.3005
R2178 VDD2.n29 VDD2.n28 9.3005
R2179 VDD2.n31 VDD2.n30 9.3005
R2180 VDD2.n14 VDD2.n13 9.3005
R2181 VDD2.n37 VDD2.n36 9.3005
R2182 VDD2.n39 VDD2.n38 9.3005
R2183 VDD2.n40 VDD2.n9 9.3005
R2184 VDD2.n130 VDD2.n71 8.92171
R2185 VDD2.n98 VDD2.n97 8.92171
R2186 VDD2.n28 VDD2.n27 8.92171
R2187 VDD2.n61 VDD2.n2 8.92171
R2188 VDD2.n131 VDD2.n69 8.14595
R2189 VDD2.n94 VDD2.n88 8.14595
R2190 VDD2.n24 VDD2.n18 8.14595
R2191 VDD2.n62 VDD2.n0 8.14595
R2192 VDD2.n93 VDD2.n90 7.3702
R2193 VDD2.n23 VDD2.n20 7.3702
R2194 VDD2.n133 VDD2.n69 5.81868
R2195 VDD2.n94 VDD2.n93 5.81868
R2196 VDD2.n24 VDD2.n23 5.81868
R2197 VDD2.n64 VDD2.n0 5.81868
R2198 VDD2.n131 VDD2.n130 5.04292
R2199 VDD2.n97 VDD2.n88 5.04292
R2200 VDD2.n27 VDD2.n18 5.04292
R2201 VDD2.n62 VDD2.n61 5.04292
R2202 VDD2.n127 VDD2.n71 4.26717
R2203 VDD2.n98 VDD2.n86 4.26717
R2204 VDD2.n28 VDD2.n16 4.26717
R2205 VDD2.n58 VDD2.n2 4.26717
R2206 VDD2.n126 VDD2.n73 3.49141
R2207 VDD2.n102 VDD2.n101 3.49141
R2208 VDD2.n32 VDD2.n31 3.49141
R2209 VDD2.n57 VDD2.n4 3.49141
R2210 VDD2.n123 VDD2.n122 2.71565
R2211 VDD2.n105 VDD2.n84 2.71565
R2212 VDD2.n35 VDD2.n14 2.71565
R2213 VDD2.n54 VDD2.n53 2.71565
R2214 VDD2.n137 VDD2.t8 2.70474
R2215 VDD2.n137 VDD2.t9 2.70474
R2216 VDD2.n135 VDD2.t1 2.70474
R2217 VDD2.n135 VDD2.t7 2.70474
R2218 VDD2.n67 VDD2.t0 2.70474
R2219 VDD2.n67 VDD2.t6 2.70474
R2220 VDD2.n65 VDD2.t2 2.70474
R2221 VDD2.n65 VDD2.t4 2.70474
R2222 VDD2.n92 VDD2.n91 2.41282
R2223 VDD2.n22 VDD2.n21 2.41282
R2224 VDD2.n136 VDD2.n134 2.0005
R2225 VDD2.n119 VDD2.n75 1.93989
R2226 VDD2.n106 VDD2.n82 1.93989
R2227 VDD2.n36 VDD2.n12 1.93989
R2228 VDD2.n50 VDD2.n6 1.93989
R2229 VDD2.n118 VDD2.n77 1.16414
R2230 VDD2.n110 VDD2.n109 1.16414
R2231 VDD2.n41 VDD2.n39 1.16414
R2232 VDD2.n49 VDD2.n8 1.16414
R2233 VDD2 VDD2.n136 0.55869
R2234 VDD2.n68 VDD2.n66 0.445154
R2235 VDD2.n115 VDD2.n114 0.388379
R2236 VDD2.n81 VDD2.n79 0.388379
R2237 VDD2.n40 VDD2.n10 0.388379
R2238 VDD2.n46 VDD2.n45 0.388379
R2239 VDD2.n132 VDD2.n70 0.155672
R2240 VDD2.n125 VDD2.n70 0.155672
R2241 VDD2.n125 VDD2.n124 0.155672
R2242 VDD2.n124 VDD2.n74 0.155672
R2243 VDD2.n117 VDD2.n74 0.155672
R2244 VDD2.n117 VDD2.n116 0.155672
R2245 VDD2.n116 VDD2.n78 0.155672
R2246 VDD2.n108 VDD2.n78 0.155672
R2247 VDD2.n108 VDD2.n107 0.155672
R2248 VDD2.n107 VDD2.n83 0.155672
R2249 VDD2.n100 VDD2.n83 0.155672
R2250 VDD2.n100 VDD2.n99 0.155672
R2251 VDD2.n99 VDD2.n87 0.155672
R2252 VDD2.n92 VDD2.n87 0.155672
R2253 VDD2.n22 VDD2.n17 0.155672
R2254 VDD2.n29 VDD2.n17 0.155672
R2255 VDD2.n30 VDD2.n29 0.155672
R2256 VDD2.n30 VDD2.n13 0.155672
R2257 VDD2.n37 VDD2.n13 0.155672
R2258 VDD2.n38 VDD2.n37 0.155672
R2259 VDD2.n38 VDD2.n9 0.155672
R2260 VDD2.n47 VDD2.n9 0.155672
R2261 VDD2.n48 VDD2.n47 0.155672
R2262 VDD2.n48 VDD2.n5 0.155672
R2263 VDD2.n55 VDD2.n5 0.155672
R2264 VDD2.n56 VDD2.n55 0.155672
R2265 VDD2.n56 VDD2.n1 0.155672
R2266 VDD2.n63 VDD2.n1 0.155672
C0 w_n3754_n3372# VTAIL 3.13618f
C1 B VN 1.13163f
C2 VDD2 VP 0.506142f
C3 w_n3754_n3372# B 9.52682f
C4 VDD2 VN 10.0564f
C5 VP VN 7.49945f
C6 VDD2 w_n3754_n3372# 2.67018f
C7 w_n3754_n3372# VP 8.3254f
C8 VTAIL VDD1 10.4613f
C9 w_n3754_n3372# VN 7.83853f
C10 B VDD1 2.24126f
C11 B VTAIL 3.46531f
C12 VDD2 VDD1 1.77762f
C13 VP VDD1 10.4063f
C14 VN VDD1 0.152305f
C15 VDD2 VTAIL 10.507299f
C16 VP VTAIL 10.4589f
C17 w_n3754_n3372# VDD1 2.55824f
C18 VN VTAIL 10.4445f
C19 VDD2 B 2.33542f
C20 B VP 1.94696f
C21 VDD2 VSUBS 1.905747f
C22 VDD1 VSUBS 1.698979f
C23 VTAIL VSUBS 1.157344f
C24 VN VSUBS 6.69547f
C25 VP VSUBS 3.465519f
C26 B VSUBS 4.610502f
C27 w_n3754_n3372# VSUBS 0.155821p
C28 VDD2.n0 VSUBS 0.029068f
C29 VDD2.n1 VSUBS 0.027626f
C30 VDD2.n2 VSUBS 0.014845f
C31 VDD2.n3 VSUBS 0.035088f
C32 VDD2.n4 VSUBS 0.015718f
C33 VDD2.n5 VSUBS 0.027626f
C34 VDD2.n6 VSUBS 0.014845f
C35 VDD2.n7 VSUBS 0.035088f
C36 VDD2.n8 VSUBS 0.015718f
C37 VDD2.n9 VSUBS 0.027626f
C38 VDD2.n10 VSUBS 0.015282f
C39 VDD2.n11 VSUBS 0.035088f
C40 VDD2.n12 VSUBS 0.015718f
C41 VDD2.n13 VSUBS 0.027626f
C42 VDD2.n14 VSUBS 0.014845f
C43 VDD2.n15 VSUBS 0.035088f
C44 VDD2.n16 VSUBS 0.015718f
C45 VDD2.n17 VSUBS 0.027626f
C46 VDD2.n18 VSUBS 0.014845f
C47 VDD2.n19 VSUBS 0.026316f
C48 VDD2.n20 VSUBS 0.026395f
C49 VDD2.t5 VSUBS 0.075611f
C50 VDD2.n21 VSUBS 0.217818f
C51 VDD2.n22 VSUBS 1.35976f
C52 VDD2.n23 VSUBS 0.014845f
C53 VDD2.n24 VSUBS 0.015718f
C54 VDD2.n25 VSUBS 0.035088f
C55 VDD2.n26 VSUBS 0.035088f
C56 VDD2.n27 VSUBS 0.015718f
C57 VDD2.n28 VSUBS 0.014845f
C58 VDD2.n29 VSUBS 0.027626f
C59 VDD2.n30 VSUBS 0.027626f
C60 VDD2.n31 VSUBS 0.014845f
C61 VDD2.n32 VSUBS 0.015718f
C62 VDD2.n33 VSUBS 0.035088f
C63 VDD2.n34 VSUBS 0.035088f
C64 VDD2.n35 VSUBS 0.015718f
C65 VDD2.n36 VSUBS 0.014845f
C66 VDD2.n37 VSUBS 0.027626f
C67 VDD2.n38 VSUBS 0.027626f
C68 VDD2.n39 VSUBS 0.014845f
C69 VDD2.n40 VSUBS 0.014845f
C70 VDD2.n41 VSUBS 0.015718f
C71 VDD2.n42 VSUBS 0.035088f
C72 VDD2.n43 VSUBS 0.035088f
C73 VDD2.n44 VSUBS 0.035088f
C74 VDD2.n45 VSUBS 0.015282f
C75 VDD2.n46 VSUBS 0.014845f
C76 VDD2.n47 VSUBS 0.027626f
C77 VDD2.n48 VSUBS 0.027626f
C78 VDD2.n49 VSUBS 0.014845f
C79 VDD2.n50 VSUBS 0.015718f
C80 VDD2.n51 VSUBS 0.035088f
C81 VDD2.n52 VSUBS 0.035088f
C82 VDD2.n53 VSUBS 0.015718f
C83 VDD2.n54 VSUBS 0.014845f
C84 VDD2.n55 VSUBS 0.027626f
C85 VDD2.n56 VSUBS 0.027626f
C86 VDD2.n57 VSUBS 0.014845f
C87 VDD2.n58 VSUBS 0.015718f
C88 VDD2.n59 VSUBS 0.035088f
C89 VDD2.n60 VSUBS 0.080562f
C90 VDD2.n61 VSUBS 0.015718f
C91 VDD2.n62 VSUBS 0.014845f
C92 VDD2.n63 VSUBS 0.060082f
C93 VDD2.n64 VSUBS 0.068671f
C94 VDD2.t2 VSUBS 0.262405f
C95 VDD2.t4 VSUBS 0.262405f
C96 VDD2.n65 VSUBS 2.03977f
C97 VDD2.n66 VSUBS 0.966105f
C98 VDD2.t0 VSUBS 0.262405f
C99 VDD2.t6 VSUBS 0.262405f
C100 VDD2.n67 VSUBS 2.05643f
C101 VDD2.n68 VSUBS 3.15451f
C102 VDD2.n69 VSUBS 0.029068f
C103 VDD2.n70 VSUBS 0.027626f
C104 VDD2.n71 VSUBS 0.014845f
C105 VDD2.n72 VSUBS 0.035088f
C106 VDD2.n73 VSUBS 0.015718f
C107 VDD2.n74 VSUBS 0.027626f
C108 VDD2.n75 VSUBS 0.014845f
C109 VDD2.n76 VSUBS 0.035088f
C110 VDD2.n77 VSUBS 0.015718f
C111 VDD2.n78 VSUBS 0.027626f
C112 VDD2.n79 VSUBS 0.015282f
C113 VDD2.n80 VSUBS 0.035088f
C114 VDD2.n81 VSUBS 0.014845f
C115 VDD2.n82 VSUBS 0.015718f
C116 VDD2.n83 VSUBS 0.027626f
C117 VDD2.n84 VSUBS 0.014845f
C118 VDD2.n85 VSUBS 0.035088f
C119 VDD2.n86 VSUBS 0.015718f
C120 VDD2.n87 VSUBS 0.027626f
C121 VDD2.n88 VSUBS 0.014845f
C122 VDD2.n89 VSUBS 0.026316f
C123 VDD2.n90 VSUBS 0.026395f
C124 VDD2.t3 VSUBS 0.075611f
C125 VDD2.n91 VSUBS 0.217818f
C126 VDD2.n92 VSUBS 1.35976f
C127 VDD2.n93 VSUBS 0.014845f
C128 VDD2.n94 VSUBS 0.015718f
C129 VDD2.n95 VSUBS 0.035088f
C130 VDD2.n96 VSUBS 0.035088f
C131 VDD2.n97 VSUBS 0.015718f
C132 VDD2.n98 VSUBS 0.014845f
C133 VDD2.n99 VSUBS 0.027626f
C134 VDD2.n100 VSUBS 0.027626f
C135 VDD2.n101 VSUBS 0.014845f
C136 VDD2.n102 VSUBS 0.015718f
C137 VDD2.n103 VSUBS 0.035088f
C138 VDD2.n104 VSUBS 0.035088f
C139 VDD2.n105 VSUBS 0.015718f
C140 VDD2.n106 VSUBS 0.014845f
C141 VDD2.n107 VSUBS 0.027626f
C142 VDD2.n108 VSUBS 0.027626f
C143 VDD2.n109 VSUBS 0.014845f
C144 VDD2.n110 VSUBS 0.015718f
C145 VDD2.n111 VSUBS 0.035088f
C146 VDD2.n112 VSUBS 0.035088f
C147 VDD2.n113 VSUBS 0.035088f
C148 VDD2.n114 VSUBS 0.015282f
C149 VDD2.n115 VSUBS 0.014845f
C150 VDD2.n116 VSUBS 0.027626f
C151 VDD2.n117 VSUBS 0.027626f
C152 VDD2.n118 VSUBS 0.014845f
C153 VDD2.n119 VSUBS 0.015718f
C154 VDD2.n120 VSUBS 0.035088f
C155 VDD2.n121 VSUBS 0.035088f
C156 VDD2.n122 VSUBS 0.015718f
C157 VDD2.n123 VSUBS 0.014845f
C158 VDD2.n124 VSUBS 0.027626f
C159 VDD2.n125 VSUBS 0.027626f
C160 VDD2.n126 VSUBS 0.014845f
C161 VDD2.n127 VSUBS 0.015718f
C162 VDD2.n128 VSUBS 0.035088f
C163 VDD2.n129 VSUBS 0.080562f
C164 VDD2.n130 VSUBS 0.015718f
C165 VDD2.n131 VSUBS 0.014845f
C166 VDD2.n132 VSUBS 0.060082f
C167 VDD2.n133 VSUBS 0.059307f
C168 VDD2.n134 VSUBS 2.93137f
C169 VDD2.t1 VSUBS 0.262405f
C170 VDD2.t7 VSUBS 0.262405f
C171 VDD2.n135 VSUBS 2.03978f
C172 VDD2.n136 VSUBS 0.755056f
C173 VDD2.t8 VSUBS 0.262405f
C174 VDD2.t9 VSUBS 0.262405f
C175 VDD2.n137 VSUBS 2.05638f
C176 VN.n0 VSUBS 0.042737f
C177 VN.t3 VSUBS 2.11286f
C178 VN.n1 VSUBS 0.045331f
C179 VN.n2 VSUBS 0.032418f
C180 VN.t9 VSUBS 2.11286f
C181 VN.n3 VSUBS 0.029692f
C182 VN.n4 VSUBS 0.032418f
C183 VN.t5 VSUBS 2.11286f
C184 VN.n5 VSUBS 0.059819f
C185 VN.n6 VSUBS 0.032418f
C186 VN.t7 VSUBS 2.11286f
C187 VN.n7 VSUBS 0.820909f
C188 VN.t4 VSUBS 2.26944f
C189 VN.n8 VSUBS 0.8375f
C190 VN.n9 VSUBS 0.242352f
C191 VN.n10 VSUBS 0.034593f
C192 VN.n11 VSUBS 0.064854f
C193 VN.n12 VSUBS 0.029692f
C194 VN.n13 VSUBS 0.032418f
C195 VN.n14 VSUBS 0.032418f
C196 VN.n15 VSUBS 0.032418f
C197 VN.n16 VSUBS 0.045277f
C198 VN.n17 VSUBS 0.754054f
C199 VN.n18 VSUBS 0.045277f
C200 VN.n19 VSUBS 0.059819f
C201 VN.n20 VSUBS 0.032418f
C202 VN.n21 VSUBS 0.032418f
C203 VN.n22 VSUBS 0.032418f
C204 VN.n23 VSUBS 0.064854f
C205 VN.n24 VSUBS 0.034593f
C206 VN.n25 VSUBS 0.754054f
C207 VN.n26 VSUBS 0.055961f
C208 VN.n27 VSUBS 0.032418f
C209 VN.n28 VSUBS 0.032418f
C210 VN.n29 VSUBS 0.032418f
C211 VN.n30 VSUBS 0.048918f
C212 VN.n31 VSUBS 0.053587f
C213 VN.n32 VSUBS 0.851014f
C214 VN.n33 VSUBS 0.03994f
C215 VN.n34 VSUBS 0.042737f
C216 VN.t6 VSUBS 2.11286f
C217 VN.n35 VSUBS 0.045331f
C218 VN.n36 VSUBS 0.032418f
C219 VN.t8 VSUBS 2.11286f
C220 VN.n37 VSUBS 0.029692f
C221 VN.n38 VSUBS 0.032418f
C222 VN.t2 VSUBS 2.11286f
C223 VN.n39 VSUBS 0.059819f
C224 VN.n40 VSUBS 0.032418f
C225 VN.t1 VSUBS 2.11286f
C226 VN.n41 VSUBS 0.820909f
C227 VN.t0 VSUBS 2.26944f
C228 VN.n42 VSUBS 0.8375f
C229 VN.n43 VSUBS 0.242352f
C230 VN.n44 VSUBS 0.034593f
C231 VN.n45 VSUBS 0.064854f
C232 VN.n46 VSUBS 0.029692f
C233 VN.n47 VSUBS 0.032418f
C234 VN.n48 VSUBS 0.032418f
C235 VN.n49 VSUBS 0.032418f
C236 VN.n50 VSUBS 0.045277f
C237 VN.n51 VSUBS 0.754054f
C238 VN.n52 VSUBS 0.045277f
C239 VN.n53 VSUBS 0.059819f
C240 VN.n54 VSUBS 0.032418f
C241 VN.n55 VSUBS 0.032418f
C242 VN.n56 VSUBS 0.032418f
C243 VN.n57 VSUBS 0.064854f
C244 VN.n58 VSUBS 0.034593f
C245 VN.n59 VSUBS 0.754054f
C246 VN.n60 VSUBS 0.055961f
C247 VN.n61 VSUBS 0.032418f
C248 VN.n62 VSUBS 0.032418f
C249 VN.n63 VSUBS 0.032418f
C250 VN.n64 VSUBS 0.048918f
C251 VN.n65 VSUBS 0.053587f
C252 VN.n66 VSUBS 0.851014f
C253 VN.n67 VSUBS 1.79811f
C254 B.n0 VSUBS 0.005478f
C255 B.n1 VSUBS 0.005478f
C256 B.n2 VSUBS 0.008663f
C257 B.n3 VSUBS 0.008663f
C258 B.n4 VSUBS 0.008663f
C259 B.n5 VSUBS 0.008663f
C260 B.n6 VSUBS 0.008663f
C261 B.n7 VSUBS 0.008663f
C262 B.n8 VSUBS 0.008663f
C263 B.n9 VSUBS 0.008663f
C264 B.n10 VSUBS 0.008663f
C265 B.n11 VSUBS 0.008663f
C266 B.n12 VSUBS 0.008663f
C267 B.n13 VSUBS 0.008663f
C268 B.n14 VSUBS 0.008663f
C269 B.n15 VSUBS 0.008663f
C270 B.n16 VSUBS 0.008663f
C271 B.n17 VSUBS 0.008663f
C272 B.n18 VSUBS 0.008663f
C273 B.n19 VSUBS 0.008663f
C274 B.n20 VSUBS 0.008663f
C275 B.n21 VSUBS 0.008663f
C276 B.n22 VSUBS 0.008663f
C277 B.n23 VSUBS 0.008663f
C278 B.n24 VSUBS 0.008663f
C279 B.n25 VSUBS 0.008663f
C280 B.n26 VSUBS 0.019693f
C281 B.n27 VSUBS 0.008663f
C282 B.n28 VSUBS 0.008663f
C283 B.n29 VSUBS 0.008663f
C284 B.n30 VSUBS 0.008663f
C285 B.n31 VSUBS 0.008663f
C286 B.n32 VSUBS 0.008663f
C287 B.n33 VSUBS 0.008663f
C288 B.n34 VSUBS 0.008663f
C289 B.n35 VSUBS 0.008663f
C290 B.n36 VSUBS 0.008663f
C291 B.n37 VSUBS 0.008663f
C292 B.n38 VSUBS 0.008663f
C293 B.n39 VSUBS 0.008663f
C294 B.n40 VSUBS 0.008663f
C295 B.n41 VSUBS 0.008663f
C296 B.n42 VSUBS 0.008663f
C297 B.n43 VSUBS 0.008663f
C298 B.n44 VSUBS 0.008663f
C299 B.n45 VSUBS 0.008663f
C300 B.n46 VSUBS 0.008663f
C301 B.n47 VSUBS 0.008663f
C302 B.t8 VSUBS 0.26159f
C303 B.t7 VSUBS 0.293298f
C304 B.t6 VSUBS 1.32279f
C305 B.n48 VSUBS 0.459113f
C306 B.n49 VSUBS 0.308977f
C307 B.n50 VSUBS 0.008663f
C308 B.n51 VSUBS 0.008663f
C309 B.n52 VSUBS 0.008663f
C310 B.n53 VSUBS 0.008663f
C311 B.t2 VSUBS 0.261594f
C312 B.t1 VSUBS 0.293301f
C313 B.t0 VSUBS 1.32279f
C314 B.n54 VSUBS 0.459109f
C315 B.n55 VSUBS 0.308973f
C316 B.n56 VSUBS 0.02007f
C317 B.n57 VSUBS 0.008663f
C318 B.n58 VSUBS 0.008663f
C319 B.n59 VSUBS 0.008663f
C320 B.n60 VSUBS 0.008663f
C321 B.n61 VSUBS 0.008663f
C322 B.n62 VSUBS 0.008663f
C323 B.n63 VSUBS 0.008663f
C324 B.n64 VSUBS 0.008663f
C325 B.n65 VSUBS 0.008663f
C326 B.n66 VSUBS 0.008663f
C327 B.n67 VSUBS 0.008663f
C328 B.n68 VSUBS 0.008663f
C329 B.n69 VSUBS 0.008663f
C330 B.n70 VSUBS 0.008663f
C331 B.n71 VSUBS 0.008663f
C332 B.n72 VSUBS 0.008663f
C333 B.n73 VSUBS 0.008663f
C334 B.n74 VSUBS 0.008663f
C335 B.n75 VSUBS 0.008663f
C336 B.n76 VSUBS 0.008663f
C337 B.n77 VSUBS 0.020818f
C338 B.n78 VSUBS 0.008663f
C339 B.n79 VSUBS 0.008663f
C340 B.n80 VSUBS 0.008663f
C341 B.n81 VSUBS 0.008663f
C342 B.n82 VSUBS 0.008663f
C343 B.n83 VSUBS 0.008663f
C344 B.n84 VSUBS 0.008663f
C345 B.n85 VSUBS 0.008663f
C346 B.n86 VSUBS 0.008663f
C347 B.n87 VSUBS 0.008663f
C348 B.n88 VSUBS 0.008663f
C349 B.n89 VSUBS 0.008663f
C350 B.n90 VSUBS 0.008663f
C351 B.n91 VSUBS 0.008663f
C352 B.n92 VSUBS 0.008663f
C353 B.n93 VSUBS 0.008663f
C354 B.n94 VSUBS 0.008663f
C355 B.n95 VSUBS 0.008663f
C356 B.n96 VSUBS 0.008663f
C357 B.n97 VSUBS 0.008663f
C358 B.n98 VSUBS 0.008663f
C359 B.n99 VSUBS 0.008663f
C360 B.n100 VSUBS 0.008663f
C361 B.n101 VSUBS 0.008663f
C362 B.n102 VSUBS 0.008663f
C363 B.n103 VSUBS 0.008663f
C364 B.n104 VSUBS 0.008663f
C365 B.n105 VSUBS 0.008663f
C366 B.n106 VSUBS 0.008663f
C367 B.n107 VSUBS 0.008663f
C368 B.n108 VSUBS 0.008663f
C369 B.n109 VSUBS 0.008663f
C370 B.n110 VSUBS 0.008663f
C371 B.n111 VSUBS 0.008663f
C372 B.n112 VSUBS 0.008663f
C373 B.n113 VSUBS 0.008663f
C374 B.n114 VSUBS 0.008663f
C375 B.n115 VSUBS 0.008663f
C376 B.n116 VSUBS 0.008663f
C377 B.n117 VSUBS 0.008663f
C378 B.n118 VSUBS 0.008663f
C379 B.n119 VSUBS 0.008663f
C380 B.n120 VSUBS 0.008663f
C381 B.n121 VSUBS 0.008663f
C382 B.n122 VSUBS 0.008663f
C383 B.n123 VSUBS 0.008663f
C384 B.n124 VSUBS 0.008663f
C385 B.n125 VSUBS 0.008663f
C386 B.n126 VSUBS 0.008663f
C387 B.n127 VSUBS 0.020818f
C388 B.n128 VSUBS 0.008663f
C389 B.n129 VSUBS 0.008663f
C390 B.n130 VSUBS 0.008663f
C391 B.n131 VSUBS 0.008663f
C392 B.n132 VSUBS 0.008663f
C393 B.n133 VSUBS 0.008663f
C394 B.n134 VSUBS 0.008663f
C395 B.n135 VSUBS 0.008663f
C396 B.n136 VSUBS 0.008663f
C397 B.n137 VSUBS 0.008663f
C398 B.n138 VSUBS 0.008663f
C399 B.n139 VSUBS 0.008663f
C400 B.n140 VSUBS 0.008663f
C401 B.n141 VSUBS 0.008663f
C402 B.n142 VSUBS 0.008663f
C403 B.n143 VSUBS 0.008663f
C404 B.n144 VSUBS 0.008663f
C405 B.n145 VSUBS 0.008663f
C406 B.n146 VSUBS 0.008663f
C407 B.n147 VSUBS 0.008663f
C408 B.t10 VSUBS 0.261594f
C409 B.t11 VSUBS 0.293301f
C410 B.t9 VSUBS 1.32279f
C411 B.n148 VSUBS 0.459109f
C412 B.n149 VSUBS 0.308973f
C413 B.n150 VSUBS 0.02007f
C414 B.n151 VSUBS 0.008663f
C415 B.n152 VSUBS 0.008663f
C416 B.n153 VSUBS 0.008663f
C417 B.n154 VSUBS 0.008663f
C418 B.n155 VSUBS 0.008663f
C419 B.t4 VSUBS 0.26159f
C420 B.t5 VSUBS 0.293298f
C421 B.t3 VSUBS 1.32279f
C422 B.n156 VSUBS 0.459113f
C423 B.n157 VSUBS 0.308977f
C424 B.n158 VSUBS 0.008663f
C425 B.n159 VSUBS 0.008663f
C426 B.n160 VSUBS 0.008663f
C427 B.n161 VSUBS 0.008663f
C428 B.n162 VSUBS 0.008663f
C429 B.n163 VSUBS 0.008663f
C430 B.n164 VSUBS 0.008663f
C431 B.n165 VSUBS 0.008663f
C432 B.n166 VSUBS 0.008663f
C433 B.n167 VSUBS 0.008663f
C434 B.n168 VSUBS 0.008663f
C435 B.n169 VSUBS 0.008663f
C436 B.n170 VSUBS 0.008663f
C437 B.n171 VSUBS 0.008663f
C438 B.n172 VSUBS 0.008663f
C439 B.n173 VSUBS 0.008663f
C440 B.n174 VSUBS 0.008663f
C441 B.n175 VSUBS 0.008663f
C442 B.n176 VSUBS 0.008663f
C443 B.n177 VSUBS 0.008663f
C444 B.n178 VSUBS 0.019693f
C445 B.n179 VSUBS 0.008663f
C446 B.n180 VSUBS 0.008663f
C447 B.n181 VSUBS 0.008663f
C448 B.n182 VSUBS 0.008663f
C449 B.n183 VSUBS 0.008663f
C450 B.n184 VSUBS 0.008663f
C451 B.n185 VSUBS 0.008663f
C452 B.n186 VSUBS 0.008663f
C453 B.n187 VSUBS 0.008663f
C454 B.n188 VSUBS 0.008663f
C455 B.n189 VSUBS 0.008663f
C456 B.n190 VSUBS 0.008663f
C457 B.n191 VSUBS 0.008663f
C458 B.n192 VSUBS 0.008663f
C459 B.n193 VSUBS 0.008663f
C460 B.n194 VSUBS 0.008663f
C461 B.n195 VSUBS 0.008663f
C462 B.n196 VSUBS 0.008663f
C463 B.n197 VSUBS 0.008663f
C464 B.n198 VSUBS 0.008663f
C465 B.n199 VSUBS 0.008663f
C466 B.n200 VSUBS 0.008663f
C467 B.n201 VSUBS 0.008663f
C468 B.n202 VSUBS 0.008663f
C469 B.n203 VSUBS 0.008663f
C470 B.n204 VSUBS 0.008663f
C471 B.n205 VSUBS 0.008663f
C472 B.n206 VSUBS 0.008663f
C473 B.n207 VSUBS 0.008663f
C474 B.n208 VSUBS 0.008663f
C475 B.n209 VSUBS 0.008663f
C476 B.n210 VSUBS 0.008663f
C477 B.n211 VSUBS 0.008663f
C478 B.n212 VSUBS 0.008663f
C479 B.n213 VSUBS 0.008663f
C480 B.n214 VSUBS 0.008663f
C481 B.n215 VSUBS 0.008663f
C482 B.n216 VSUBS 0.008663f
C483 B.n217 VSUBS 0.008663f
C484 B.n218 VSUBS 0.008663f
C485 B.n219 VSUBS 0.008663f
C486 B.n220 VSUBS 0.008663f
C487 B.n221 VSUBS 0.008663f
C488 B.n222 VSUBS 0.008663f
C489 B.n223 VSUBS 0.008663f
C490 B.n224 VSUBS 0.008663f
C491 B.n225 VSUBS 0.008663f
C492 B.n226 VSUBS 0.008663f
C493 B.n227 VSUBS 0.008663f
C494 B.n228 VSUBS 0.008663f
C495 B.n229 VSUBS 0.008663f
C496 B.n230 VSUBS 0.008663f
C497 B.n231 VSUBS 0.008663f
C498 B.n232 VSUBS 0.008663f
C499 B.n233 VSUBS 0.008663f
C500 B.n234 VSUBS 0.008663f
C501 B.n235 VSUBS 0.008663f
C502 B.n236 VSUBS 0.008663f
C503 B.n237 VSUBS 0.008663f
C504 B.n238 VSUBS 0.008663f
C505 B.n239 VSUBS 0.008663f
C506 B.n240 VSUBS 0.008663f
C507 B.n241 VSUBS 0.008663f
C508 B.n242 VSUBS 0.008663f
C509 B.n243 VSUBS 0.008663f
C510 B.n244 VSUBS 0.008663f
C511 B.n245 VSUBS 0.008663f
C512 B.n246 VSUBS 0.008663f
C513 B.n247 VSUBS 0.008663f
C514 B.n248 VSUBS 0.008663f
C515 B.n249 VSUBS 0.008663f
C516 B.n250 VSUBS 0.008663f
C517 B.n251 VSUBS 0.008663f
C518 B.n252 VSUBS 0.008663f
C519 B.n253 VSUBS 0.008663f
C520 B.n254 VSUBS 0.008663f
C521 B.n255 VSUBS 0.008663f
C522 B.n256 VSUBS 0.008663f
C523 B.n257 VSUBS 0.008663f
C524 B.n258 VSUBS 0.008663f
C525 B.n259 VSUBS 0.008663f
C526 B.n260 VSUBS 0.008663f
C527 B.n261 VSUBS 0.008663f
C528 B.n262 VSUBS 0.008663f
C529 B.n263 VSUBS 0.008663f
C530 B.n264 VSUBS 0.008663f
C531 B.n265 VSUBS 0.008663f
C532 B.n266 VSUBS 0.008663f
C533 B.n267 VSUBS 0.008663f
C534 B.n268 VSUBS 0.008663f
C535 B.n269 VSUBS 0.008663f
C536 B.n270 VSUBS 0.008663f
C537 B.n271 VSUBS 0.008663f
C538 B.n272 VSUBS 0.008663f
C539 B.n273 VSUBS 0.019693f
C540 B.n274 VSUBS 0.020818f
C541 B.n275 VSUBS 0.020818f
C542 B.n276 VSUBS 0.008663f
C543 B.n277 VSUBS 0.008663f
C544 B.n278 VSUBS 0.008663f
C545 B.n279 VSUBS 0.008663f
C546 B.n280 VSUBS 0.008663f
C547 B.n281 VSUBS 0.008663f
C548 B.n282 VSUBS 0.008663f
C549 B.n283 VSUBS 0.008663f
C550 B.n284 VSUBS 0.008663f
C551 B.n285 VSUBS 0.008663f
C552 B.n286 VSUBS 0.008663f
C553 B.n287 VSUBS 0.008663f
C554 B.n288 VSUBS 0.008663f
C555 B.n289 VSUBS 0.008663f
C556 B.n290 VSUBS 0.008663f
C557 B.n291 VSUBS 0.008663f
C558 B.n292 VSUBS 0.008663f
C559 B.n293 VSUBS 0.008663f
C560 B.n294 VSUBS 0.008663f
C561 B.n295 VSUBS 0.008663f
C562 B.n296 VSUBS 0.008663f
C563 B.n297 VSUBS 0.008663f
C564 B.n298 VSUBS 0.008663f
C565 B.n299 VSUBS 0.008663f
C566 B.n300 VSUBS 0.008663f
C567 B.n301 VSUBS 0.008663f
C568 B.n302 VSUBS 0.008663f
C569 B.n303 VSUBS 0.008663f
C570 B.n304 VSUBS 0.008663f
C571 B.n305 VSUBS 0.008663f
C572 B.n306 VSUBS 0.008663f
C573 B.n307 VSUBS 0.008663f
C574 B.n308 VSUBS 0.008663f
C575 B.n309 VSUBS 0.008663f
C576 B.n310 VSUBS 0.008663f
C577 B.n311 VSUBS 0.008663f
C578 B.n312 VSUBS 0.008663f
C579 B.n313 VSUBS 0.008663f
C580 B.n314 VSUBS 0.008663f
C581 B.n315 VSUBS 0.008663f
C582 B.n316 VSUBS 0.008663f
C583 B.n317 VSUBS 0.008663f
C584 B.n318 VSUBS 0.008663f
C585 B.n319 VSUBS 0.008663f
C586 B.n320 VSUBS 0.008663f
C587 B.n321 VSUBS 0.008663f
C588 B.n322 VSUBS 0.008663f
C589 B.n323 VSUBS 0.008663f
C590 B.n324 VSUBS 0.008663f
C591 B.n325 VSUBS 0.008663f
C592 B.n326 VSUBS 0.008663f
C593 B.n327 VSUBS 0.008663f
C594 B.n328 VSUBS 0.008663f
C595 B.n329 VSUBS 0.008663f
C596 B.n330 VSUBS 0.008663f
C597 B.n331 VSUBS 0.008663f
C598 B.n332 VSUBS 0.008663f
C599 B.n333 VSUBS 0.008663f
C600 B.n334 VSUBS 0.008663f
C601 B.n335 VSUBS 0.008663f
C602 B.n336 VSUBS 0.005987f
C603 B.n337 VSUBS 0.02007f
C604 B.n338 VSUBS 0.007007f
C605 B.n339 VSUBS 0.008663f
C606 B.n340 VSUBS 0.008663f
C607 B.n341 VSUBS 0.008663f
C608 B.n342 VSUBS 0.008663f
C609 B.n343 VSUBS 0.008663f
C610 B.n344 VSUBS 0.008663f
C611 B.n345 VSUBS 0.008663f
C612 B.n346 VSUBS 0.008663f
C613 B.n347 VSUBS 0.008663f
C614 B.n348 VSUBS 0.008663f
C615 B.n349 VSUBS 0.008663f
C616 B.n350 VSUBS 0.007007f
C617 B.n351 VSUBS 0.008663f
C618 B.n352 VSUBS 0.008663f
C619 B.n353 VSUBS 0.005987f
C620 B.n354 VSUBS 0.008663f
C621 B.n355 VSUBS 0.008663f
C622 B.n356 VSUBS 0.008663f
C623 B.n357 VSUBS 0.008663f
C624 B.n358 VSUBS 0.008663f
C625 B.n359 VSUBS 0.008663f
C626 B.n360 VSUBS 0.008663f
C627 B.n361 VSUBS 0.008663f
C628 B.n362 VSUBS 0.008663f
C629 B.n363 VSUBS 0.008663f
C630 B.n364 VSUBS 0.008663f
C631 B.n365 VSUBS 0.008663f
C632 B.n366 VSUBS 0.008663f
C633 B.n367 VSUBS 0.008663f
C634 B.n368 VSUBS 0.008663f
C635 B.n369 VSUBS 0.008663f
C636 B.n370 VSUBS 0.008663f
C637 B.n371 VSUBS 0.008663f
C638 B.n372 VSUBS 0.008663f
C639 B.n373 VSUBS 0.008663f
C640 B.n374 VSUBS 0.008663f
C641 B.n375 VSUBS 0.008663f
C642 B.n376 VSUBS 0.008663f
C643 B.n377 VSUBS 0.008663f
C644 B.n378 VSUBS 0.008663f
C645 B.n379 VSUBS 0.008663f
C646 B.n380 VSUBS 0.008663f
C647 B.n381 VSUBS 0.008663f
C648 B.n382 VSUBS 0.008663f
C649 B.n383 VSUBS 0.008663f
C650 B.n384 VSUBS 0.008663f
C651 B.n385 VSUBS 0.008663f
C652 B.n386 VSUBS 0.008663f
C653 B.n387 VSUBS 0.008663f
C654 B.n388 VSUBS 0.008663f
C655 B.n389 VSUBS 0.008663f
C656 B.n390 VSUBS 0.008663f
C657 B.n391 VSUBS 0.008663f
C658 B.n392 VSUBS 0.008663f
C659 B.n393 VSUBS 0.008663f
C660 B.n394 VSUBS 0.008663f
C661 B.n395 VSUBS 0.008663f
C662 B.n396 VSUBS 0.008663f
C663 B.n397 VSUBS 0.008663f
C664 B.n398 VSUBS 0.008663f
C665 B.n399 VSUBS 0.008663f
C666 B.n400 VSUBS 0.008663f
C667 B.n401 VSUBS 0.008663f
C668 B.n402 VSUBS 0.008663f
C669 B.n403 VSUBS 0.008663f
C670 B.n404 VSUBS 0.008663f
C671 B.n405 VSUBS 0.008663f
C672 B.n406 VSUBS 0.008663f
C673 B.n407 VSUBS 0.008663f
C674 B.n408 VSUBS 0.008663f
C675 B.n409 VSUBS 0.008663f
C676 B.n410 VSUBS 0.008663f
C677 B.n411 VSUBS 0.008663f
C678 B.n412 VSUBS 0.008663f
C679 B.n413 VSUBS 0.008663f
C680 B.n414 VSUBS 0.020818f
C681 B.n415 VSUBS 0.019693f
C682 B.n416 VSUBS 0.019693f
C683 B.n417 VSUBS 0.008663f
C684 B.n418 VSUBS 0.008663f
C685 B.n419 VSUBS 0.008663f
C686 B.n420 VSUBS 0.008663f
C687 B.n421 VSUBS 0.008663f
C688 B.n422 VSUBS 0.008663f
C689 B.n423 VSUBS 0.008663f
C690 B.n424 VSUBS 0.008663f
C691 B.n425 VSUBS 0.008663f
C692 B.n426 VSUBS 0.008663f
C693 B.n427 VSUBS 0.008663f
C694 B.n428 VSUBS 0.008663f
C695 B.n429 VSUBS 0.008663f
C696 B.n430 VSUBS 0.008663f
C697 B.n431 VSUBS 0.008663f
C698 B.n432 VSUBS 0.008663f
C699 B.n433 VSUBS 0.008663f
C700 B.n434 VSUBS 0.008663f
C701 B.n435 VSUBS 0.008663f
C702 B.n436 VSUBS 0.008663f
C703 B.n437 VSUBS 0.008663f
C704 B.n438 VSUBS 0.008663f
C705 B.n439 VSUBS 0.008663f
C706 B.n440 VSUBS 0.008663f
C707 B.n441 VSUBS 0.008663f
C708 B.n442 VSUBS 0.008663f
C709 B.n443 VSUBS 0.008663f
C710 B.n444 VSUBS 0.008663f
C711 B.n445 VSUBS 0.008663f
C712 B.n446 VSUBS 0.008663f
C713 B.n447 VSUBS 0.008663f
C714 B.n448 VSUBS 0.008663f
C715 B.n449 VSUBS 0.008663f
C716 B.n450 VSUBS 0.008663f
C717 B.n451 VSUBS 0.008663f
C718 B.n452 VSUBS 0.008663f
C719 B.n453 VSUBS 0.008663f
C720 B.n454 VSUBS 0.008663f
C721 B.n455 VSUBS 0.008663f
C722 B.n456 VSUBS 0.008663f
C723 B.n457 VSUBS 0.008663f
C724 B.n458 VSUBS 0.008663f
C725 B.n459 VSUBS 0.008663f
C726 B.n460 VSUBS 0.008663f
C727 B.n461 VSUBS 0.008663f
C728 B.n462 VSUBS 0.008663f
C729 B.n463 VSUBS 0.008663f
C730 B.n464 VSUBS 0.008663f
C731 B.n465 VSUBS 0.008663f
C732 B.n466 VSUBS 0.008663f
C733 B.n467 VSUBS 0.008663f
C734 B.n468 VSUBS 0.008663f
C735 B.n469 VSUBS 0.008663f
C736 B.n470 VSUBS 0.008663f
C737 B.n471 VSUBS 0.008663f
C738 B.n472 VSUBS 0.008663f
C739 B.n473 VSUBS 0.008663f
C740 B.n474 VSUBS 0.008663f
C741 B.n475 VSUBS 0.008663f
C742 B.n476 VSUBS 0.008663f
C743 B.n477 VSUBS 0.008663f
C744 B.n478 VSUBS 0.008663f
C745 B.n479 VSUBS 0.008663f
C746 B.n480 VSUBS 0.008663f
C747 B.n481 VSUBS 0.008663f
C748 B.n482 VSUBS 0.008663f
C749 B.n483 VSUBS 0.008663f
C750 B.n484 VSUBS 0.008663f
C751 B.n485 VSUBS 0.008663f
C752 B.n486 VSUBS 0.008663f
C753 B.n487 VSUBS 0.008663f
C754 B.n488 VSUBS 0.008663f
C755 B.n489 VSUBS 0.008663f
C756 B.n490 VSUBS 0.008663f
C757 B.n491 VSUBS 0.008663f
C758 B.n492 VSUBS 0.008663f
C759 B.n493 VSUBS 0.008663f
C760 B.n494 VSUBS 0.008663f
C761 B.n495 VSUBS 0.008663f
C762 B.n496 VSUBS 0.008663f
C763 B.n497 VSUBS 0.008663f
C764 B.n498 VSUBS 0.008663f
C765 B.n499 VSUBS 0.008663f
C766 B.n500 VSUBS 0.008663f
C767 B.n501 VSUBS 0.008663f
C768 B.n502 VSUBS 0.008663f
C769 B.n503 VSUBS 0.008663f
C770 B.n504 VSUBS 0.008663f
C771 B.n505 VSUBS 0.008663f
C772 B.n506 VSUBS 0.008663f
C773 B.n507 VSUBS 0.008663f
C774 B.n508 VSUBS 0.008663f
C775 B.n509 VSUBS 0.008663f
C776 B.n510 VSUBS 0.008663f
C777 B.n511 VSUBS 0.008663f
C778 B.n512 VSUBS 0.008663f
C779 B.n513 VSUBS 0.008663f
C780 B.n514 VSUBS 0.008663f
C781 B.n515 VSUBS 0.008663f
C782 B.n516 VSUBS 0.008663f
C783 B.n517 VSUBS 0.008663f
C784 B.n518 VSUBS 0.008663f
C785 B.n519 VSUBS 0.008663f
C786 B.n520 VSUBS 0.008663f
C787 B.n521 VSUBS 0.008663f
C788 B.n522 VSUBS 0.008663f
C789 B.n523 VSUBS 0.008663f
C790 B.n524 VSUBS 0.008663f
C791 B.n525 VSUBS 0.008663f
C792 B.n526 VSUBS 0.008663f
C793 B.n527 VSUBS 0.008663f
C794 B.n528 VSUBS 0.008663f
C795 B.n529 VSUBS 0.008663f
C796 B.n530 VSUBS 0.008663f
C797 B.n531 VSUBS 0.008663f
C798 B.n532 VSUBS 0.008663f
C799 B.n533 VSUBS 0.008663f
C800 B.n534 VSUBS 0.008663f
C801 B.n535 VSUBS 0.008663f
C802 B.n536 VSUBS 0.008663f
C803 B.n537 VSUBS 0.008663f
C804 B.n538 VSUBS 0.008663f
C805 B.n539 VSUBS 0.008663f
C806 B.n540 VSUBS 0.008663f
C807 B.n541 VSUBS 0.008663f
C808 B.n542 VSUBS 0.008663f
C809 B.n543 VSUBS 0.008663f
C810 B.n544 VSUBS 0.008663f
C811 B.n545 VSUBS 0.008663f
C812 B.n546 VSUBS 0.008663f
C813 B.n547 VSUBS 0.008663f
C814 B.n548 VSUBS 0.008663f
C815 B.n549 VSUBS 0.008663f
C816 B.n550 VSUBS 0.008663f
C817 B.n551 VSUBS 0.008663f
C818 B.n552 VSUBS 0.008663f
C819 B.n553 VSUBS 0.008663f
C820 B.n554 VSUBS 0.008663f
C821 B.n555 VSUBS 0.008663f
C822 B.n556 VSUBS 0.008663f
C823 B.n557 VSUBS 0.008663f
C824 B.n558 VSUBS 0.008663f
C825 B.n559 VSUBS 0.008663f
C826 B.n560 VSUBS 0.008663f
C827 B.n561 VSUBS 0.008663f
C828 B.n562 VSUBS 0.019693f
C829 B.n563 VSUBS 0.020718f
C830 B.n564 VSUBS 0.019793f
C831 B.n565 VSUBS 0.008663f
C832 B.n566 VSUBS 0.008663f
C833 B.n567 VSUBS 0.008663f
C834 B.n568 VSUBS 0.008663f
C835 B.n569 VSUBS 0.008663f
C836 B.n570 VSUBS 0.008663f
C837 B.n571 VSUBS 0.008663f
C838 B.n572 VSUBS 0.008663f
C839 B.n573 VSUBS 0.008663f
C840 B.n574 VSUBS 0.008663f
C841 B.n575 VSUBS 0.008663f
C842 B.n576 VSUBS 0.008663f
C843 B.n577 VSUBS 0.008663f
C844 B.n578 VSUBS 0.008663f
C845 B.n579 VSUBS 0.008663f
C846 B.n580 VSUBS 0.008663f
C847 B.n581 VSUBS 0.008663f
C848 B.n582 VSUBS 0.008663f
C849 B.n583 VSUBS 0.008663f
C850 B.n584 VSUBS 0.008663f
C851 B.n585 VSUBS 0.008663f
C852 B.n586 VSUBS 0.008663f
C853 B.n587 VSUBS 0.008663f
C854 B.n588 VSUBS 0.008663f
C855 B.n589 VSUBS 0.008663f
C856 B.n590 VSUBS 0.008663f
C857 B.n591 VSUBS 0.008663f
C858 B.n592 VSUBS 0.008663f
C859 B.n593 VSUBS 0.008663f
C860 B.n594 VSUBS 0.008663f
C861 B.n595 VSUBS 0.008663f
C862 B.n596 VSUBS 0.008663f
C863 B.n597 VSUBS 0.008663f
C864 B.n598 VSUBS 0.008663f
C865 B.n599 VSUBS 0.008663f
C866 B.n600 VSUBS 0.008663f
C867 B.n601 VSUBS 0.008663f
C868 B.n602 VSUBS 0.008663f
C869 B.n603 VSUBS 0.008663f
C870 B.n604 VSUBS 0.008663f
C871 B.n605 VSUBS 0.008663f
C872 B.n606 VSUBS 0.008663f
C873 B.n607 VSUBS 0.008663f
C874 B.n608 VSUBS 0.008663f
C875 B.n609 VSUBS 0.008663f
C876 B.n610 VSUBS 0.008663f
C877 B.n611 VSUBS 0.008663f
C878 B.n612 VSUBS 0.008663f
C879 B.n613 VSUBS 0.008663f
C880 B.n614 VSUBS 0.008663f
C881 B.n615 VSUBS 0.008663f
C882 B.n616 VSUBS 0.008663f
C883 B.n617 VSUBS 0.008663f
C884 B.n618 VSUBS 0.008663f
C885 B.n619 VSUBS 0.008663f
C886 B.n620 VSUBS 0.008663f
C887 B.n621 VSUBS 0.008663f
C888 B.n622 VSUBS 0.008663f
C889 B.n623 VSUBS 0.008663f
C890 B.n624 VSUBS 0.008663f
C891 B.n625 VSUBS 0.005987f
C892 B.n626 VSUBS 0.008663f
C893 B.n627 VSUBS 0.008663f
C894 B.n628 VSUBS 0.007007f
C895 B.n629 VSUBS 0.008663f
C896 B.n630 VSUBS 0.008663f
C897 B.n631 VSUBS 0.008663f
C898 B.n632 VSUBS 0.008663f
C899 B.n633 VSUBS 0.008663f
C900 B.n634 VSUBS 0.008663f
C901 B.n635 VSUBS 0.008663f
C902 B.n636 VSUBS 0.008663f
C903 B.n637 VSUBS 0.008663f
C904 B.n638 VSUBS 0.008663f
C905 B.n639 VSUBS 0.008663f
C906 B.n640 VSUBS 0.007007f
C907 B.n641 VSUBS 0.02007f
C908 B.n642 VSUBS 0.005987f
C909 B.n643 VSUBS 0.008663f
C910 B.n644 VSUBS 0.008663f
C911 B.n645 VSUBS 0.008663f
C912 B.n646 VSUBS 0.008663f
C913 B.n647 VSUBS 0.008663f
C914 B.n648 VSUBS 0.008663f
C915 B.n649 VSUBS 0.008663f
C916 B.n650 VSUBS 0.008663f
C917 B.n651 VSUBS 0.008663f
C918 B.n652 VSUBS 0.008663f
C919 B.n653 VSUBS 0.008663f
C920 B.n654 VSUBS 0.008663f
C921 B.n655 VSUBS 0.008663f
C922 B.n656 VSUBS 0.008663f
C923 B.n657 VSUBS 0.008663f
C924 B.n658 VSUBS 0.008663f
C925 B.n659 VSUBS 0.008663f
C926 B.n660 VSUBS 0.008663f
C927 B.n661 VSUBS 0.008663f
C928 B.n662 VSUBS 0.008663f
C929 B.n663 VSUBS 0.008663f
C930 B.n664 VSUBS 0.008663f
C931 B.n665 VSUBS 0.008663f
C932 B.n666 VSUBS 0.008663f
C933 B.n667 VSUBS 0.008663f
C934 B.n668 VSUBS 0.008663f
C935 B.n669 VSUBS 0.008663f
C936 B.n670 VSUBS 0.008663f
C937 B.n671 VSUBS 0.008663f
C938 B.n672 VSUBS 0.008663f
C939 B.n673 VSUBS 0.008663f
C940 B.n674 VSUBS 0.008663f
C941 B.n675 VSUBS 0.008663f
C942 B.n676 VSUBS 0.008663f
C943 B.n677 VSUBS 0.008663f
C944 B.n678 VSUBS 0.008663f
C945 B.n679 VSUBS 0.008663f
C946 B.n680 VSUBS 0.008663f
C947 B.n681 VSUBS 0.008663f
C948 B.n682 VSUBS 0.008663f
C949 B.n683 VSUBS 0.008663f
C950 B.n684 VSUBS 0.008663f
C951 B.n685 VSUBS 0.008663f
C952 B.n686 VSUBS 0.008663f
C953 B.n687 VSUBS 0.008663f
C954 B.n688 VSUBS 0.008663f
C955 B.n689 VSUBS 0.008663f
C956 B.n690 VSUBS 0.008663f
C957 B.n691 VSUBS 0.008663f
C958 B.n692 VSUBS 0.008663f
C959 B.n693 VSUBS 0.008663f
C960 B.n694 VSUBS 0.008663f
C961 B.n695 VSUBS 0.008663f
C962 B.n696 VSUBS 0.008663f
C963 B.n697 VSUBS 0.008663f
C964 B.n698 VSUBS 0.008663f
C965 B.n699 VSUBS 0.008663f
C966 B.n700 VSUBS 0.008663f
C967 B.n701 VSUBS 0.008663f
C968 B.n702 VSUBS 0.008663f
C969 B.n703 VSUBS 0.020818f
C970 B.n704 VSUBS 0.020818f
C971 B.n705 VSUBS 0.019693f
C972 B.n706 VSUBS 0.008663f
C973 B.n707 VSUBS 0.008663f
C974 B.n708 VSUBS 0.008663f
C975 B.n709 VSUBS 0.008663f
C976 B.n710 VSUBS 0.008663f
C977 B.n711 VSUBS 0.008663f
C978 B.n712 VSUBS 0.008663f
C979 B.n713 VSUBS 0.008663f
C980 B.n714 VSUBS 0.008663f
C981 B.n715 VSUBS 0.008663f
C982 B.n716 VSUBS 0.008663f
C983 B.n717 VSUBS 0.008663f
C984 B.n718 VSUBS 0.008663f
C985 B.n719 VSUBS 0.008663f
C986 B.n720 VSUBS 0.008663f
C987 B.n721 VSUBS 0.008663f
C988 B.n722 VSUBS 0.008663f
C989 B.n723 VSUBS 0.008663f
C990 B.n724 VSUBS 0.008663f
C991 B.n725 VSUBS 0.008663f
C992 B.n726 VSUBS 0.008663f
C993 B.n727 VSUBS 0.008663f
C994 B.n728 VSUBS 0.008663f
C995 B.n729 VSUBS 0.008663f
C996 B.n730 VSUBS 0.008663f
C997 B.n731 VSUBS 0.008663f
C998 B.n732 VSUBS 0.008663f
C999 B.n733 VSUBS 0.008663f
C1000 B.n734 VSUBS 0.008663f
C1001 B.n735 VSUBS 0.008663f
C1002 B.n736 VSUBS 0.008663f
C1003 B.n737 VSUBS 0.008663f
C1004 B.n738 VSUBS 0.008663f
C1005 B.n739 VSUBS 0.008663f
C1006 B.n740 VSUBS 0.008663f
C1007 B.n741 VSUBS 0.008663f
C1008 B.n742 VSUBS 0.008663f
C1009 B.n743 VSUBS 0.008663f
C1010 B.n744 VSUBS 0.008663f
C1011 B.n745 VSUBS 0.008663f
C1012 B.n746 VSUBS 0.008663f
C1013 B.n747 VSUBS 0.008663f
C1014 B.n748 VSUBS 0.008663f
C1015 B.n749 VSUBS 0.008663f
C1016 B.n750 VSUBS 0.008663f
C1017 B.n751 VSUBS 0.008663f
C1018 B.n752 VSUBS 0.008663f
C1019 B.n753 VSUBS 0.008663f
C1020 B.n754 VSUBS 0.008663f
C1021 B.n755 VSUBS 0.008663f
C1022 B.n756 VSUBS 0.008663f
C1023 B.n757 VSUBS 0.008663f
C1024 B.n758 VSUBS 0.008663f
C1025 B.n759 VSUBS 0.008663f
C1026 B.n760 VSUBS 0.008663f
C1027 B.n761 VSUBS 0.008663f
C1028 B.n762 VSUBS 0.008663f
C1029 B.n763 VSUBS 0.008663f
C1030 B.n764 VSUBS 0.008663f
C1031 B.n765 VSUBS 0.008663f
C1032 B.n766 VSUBS 0.008663f
C1033 B.n767 VSUBS 0.008663f
C1034 B.n768 VSUBS 0.008663f
C1035 B.n769 VSUBS 0.008663f
C1036 B.n770 VSUBS 0.008663f
C1037 B.n771 VSUBS 0.008663f
C1038 B.n772 VSUBS 0.008663f
C1039 B.n773 VSUBS 0.008663f
C1040 B.n774 VSUBS 0.008663f
C1041 B.n775 VSUBS 0.008663f
C1042 B.n776 VSUBS 0.008663f
C1043 B.n777 VSUBS 0.008663f
C1044 B.n778 VSUBS 0.008663f
C1045 B.n779 VSUBS 0.019615f
C1046 VDD1.n0 VSUBS 0.029066f
C1047 VDD1.n1 VSUBS 0.027624f
C1048 VDD1.n2 VSUBS 0.014844f
C1049 VDD1.n3 VSUBS 0.035085f
C1050 VDD1.n4 VSUBS 0.015717f
C1051 VDD1.n5 VSUBS 0.027624f
C1052 VDD1.n6 VSUBS 0.014844f
C1053 VDD1.n7 VSUBS 0.035085f
C1054 VDD1.n8 VSUBS 0.015717f
C1055 VDD1.n9 VSUBS 0.027624f
C1056 VDD1.n10 VSUBS 0.01528f
C1057 VDD1.n11 VSUBS 0.035085f
C1058 VDD1.n12 VSUBS 0.014844f
C1059 VDD1.n13 VSUBS 0.015717f
C1060 VDD1.n14 VSUBS 0.027624f
C1061 VDD1.n15 VSUBS 0.014844f
C1062 VDD1.n16 VSUBS 0.035085f
C1063 VDD1.n17 VSUBS 0.015717f
C1064 VDD1.n18 VSUBS 0.027624f
C1065 VDD1.n19 VSUBS 0.014844f
C1066 VDD1.n20 VSUBS 0.026314f
C1067 VDD1.n21 VSUBS 0.026393f
C1068 VDD1.t4 VSUBS 0.075605f
C1069 VDD1.n22 VSUBS 0.217801f
C1070 VDD1.n23 VSUBS 1.35966f
C1071 VDD1.n24 VSUBS 0.014844f
C1072 VDD1.n25 VSUBS 0.015717f
C1073 VDD1.n26 VSUBS 0.035085f
C1074 VDD1.n27 VSUBS 0.035085f
C1075 VDD1.n28 VSUBS 0.015717f
C1076 VDD1.n29 VSUBS 0.014844f
C1077 VDD1.n30 VSUBS 0.027624f
C1078 VDD1.n31 VSUBS 0.027624f
C1079 VDD1.n32 VSUBS 0.014844f
C1080 VDD1.n33 VSUBS 0.015717f
C1081 VDD1.n34 VSUBS 0.035085f
C1082 VDD1.n35 VSUBS 0.035085f
C1083 VDD1.n36 VSUBS 0.015717f
C1084 VDD1.n37 VSUBS 0.014844f
C1085 VDD1.n38 VSUBS 0.027624f
C1086 VDD1.n39 VSUBS 0.027624f
C1087 VDD1.n40 VSUBS 0.014844f
C1088 VDD1.n41 VSUBS 0.015717f
C1089 VDD1.n42 VSUBS 0.035085f
C1090 VDD1.n43 VSUBS 0.035085f
C1091 VDD1.n44 VSUBS 0.035085f
C1092 VDD1.n45 VSUBS 0.01528f
C1093 VDD1.n46 VSUBS 0.014844f
C1094 VDD1.n47 VSUBS 0.027624f
C1095 VDD1.n48 VSUBS 0.027624f
C1096 VDD1.n49 VSUBS 0.014844f
C1097 VDD1.n50 VSUBS 0.015717f
C1098 VDD1.n51 VSUBS 0.035085f
C1099 VDD1.n52 VSUBS 0.035085f
C1100 VDD1.n53 VSUBS 0.015717f
C1101 VDD1.n54 VSUBS 0.014844f
C1102 VDD1.n55 VSUBS 0.027624f
C1103 VDD1.n56 VSUBS 0.027624f
C1104 VDD1.n57 VSUBS 0.014844f
C1105 VDD1.n58 VSUBS 0.015717f
C1106 VDD1.n59 VSUBS 0.035085f
C1107 VDD1.n60 VSUBS 0.080555f
C1108 VDD1.n61 VSUBS 0.015717f
C1109 VDD1.n62 VSUBS 0.014844f
C1110 VDD1.n63 VSUBS 0.060077f
C1111 VDD1.n64 VSUBS 0.068666f
C1112 VDD1.t1 VSUBS 0.262384f
C1113 VDD1.t2 VSUBS 0.262384f
C1114 VDD1.n65 VSUBS 2.03962f
C1115 VDD1.n66 VSUBS 0.974683f
C1116 VDD1.n67 VSUBS 0.029066f
C1117 VDD1.n68 VSUBS 0.027624f
C1118 VDD1.n69 VSUBS 0.014844f
C1119 VDD1.n70 VSUBS 0.035085f
C1120 VDD1.n71 VSUBS 0.015717f
C1121 VDD1.n72 VSUBS 0.027624f
C1122 VDD1.n73 VSUBS 0.014844f
C1123 VDD1.n74 VSUBS 0.035085f
C1124 VDD1.n75 VSUBS 0.015717f
C1125 VDD1.n76 VSUBS 0.027624f
C1126 VDD1.n77 VSUBS 0.01528f
C1127 VDD1.n78 VSUBS 0.035085f
C1128 VDD1.n79 VSUBS 0.015717f
C1129 VDD1.n80 VSUBS 0.027624f
C1130 VDD1.n81 VSUBS 0.014844f
C1131 VDD1.n82 VSUBS 0.035085f
C1132 VDD1.n83 VSUBS 0.015717f
C1133 VDD1.n84 VSUBS 0.027624f
C1134 VDD1.n85 VSUBS 0.014844f
C1135 VDD1.n86 VSUBS 0.026314f
C1136 VDD1.n87 VSUBS 0.026393f
C1137 VDD1.t6 VSUBS 0.075605f
C1138 VDD1.n88 VSUBS 0.217801f
C1139 VDD1.n89 VSUBS 1.35966f
C1140 VDD1.n90 VSUBS 0.014844f
C1141 VDD1.n91 VSUBS 0.015717f
C1142 VDD1.n92 VSUBS 0.035085f
C1143 VDD1.n93 VSUBS 0.035085f
C1144 VDD1.n94 VSUBS 0.015717f
C1145 VDD1.n95 VSUBS 0.014844f
C1146 VDD1.n96 VSUBS 0.027624f
C1147 VDD1.n97 VSUBS 0.027624f
C1148 VDD1.n98 VSUBS 0.014844f
C1149 VDD1.n99 VSUBS 0.015717f
C1150 VDD1.n100 VSUBS 0.035085f
C1151 VDD1.n101 VSUBS 0.035085f
C1152 VDD1.n102 VSUBS 0.015717f
C1153 VDD1.n103 VSUBS 0.014844f
C1154 VDD1.n104 VSUBS 0.027624f
C1155 VDD1.n105 VSUBS 0.027624f
C1156 VDD1.n106 VSUBS 0.014844f
C1157 VDD1.n107 VSUBS 0.014844f
C1158 VDD1.n108 VSUBS 0.015717f
C1159 VDD1.n109 VSUBS 0.035085f
C1160 VDD1.n110 VSUBS 0.035085f
C1161 VDD1.n111 VSUBS 0.035085f
C1162 VDD1.n112 VSUBS 0.01528f
C1163 VDD1.n113 VSUBS 0.014844f
C1164 VDD1.n114 VSUBS 0.027624f
C1165 VDD1.n115 VSUBS 0.027624f
C1166 VDD1.n116 VSUBS 0.014844f
C1167 VDD1.n117 VSUBS 0.015717f
C1168 VDD1.n118 VSUBS 0.035085f
C1169 VDD1.n119 VSUBS 0.035085f
C1170 VDD1.n120 VSUBS 0.015717f
C1171 VDD1.n121 VSUBS 0.014844f
C1172 VDD1.n122 VSUBS 0.027624f
C1173 VDD1.n123 VSUBS 0.027624f
C1174 VDD1.n124 VSUBS 0.014844f
C1175 VDD1.n125 VSUBS 0.015717f
C1176 VDD1.n126 VSUBS 0.035085f
C1177 VDD1.n127 VSUBS 0.080555f
C1178 VDD1.n128 VSUBS 0.015717f
C1179 VDD1.n129 VSUBS 0.014844f
C1180 VDD1.n130 VSUBS 0.060077f
C1181 VDD1.n131 VSUBS 0.068666f
C1182 VDD1.t7 VSUBS 0.262384f
C1183 VDD1.t0 VSUBS 0.262384f
C1184 VDD1.n132 VSUBS 2.03961f
C1185 VDD1.n133 VSUBS 0.966028f
C1186 VDD1.t5 VSUBS 0.262384f
C1187 VDD1.t9 VSUBS 0.262384f
C1188 VDD1.n134 VSUBS 2.05626f
C1189 VDD1.n135 VSUBS 3.27466f
C1190 VDD1.t8 VSUBS 0.262384f
C1191 VDD1.t3 VSUBS 0.262384f
C1192 VDD1.n136 VSUBS 2.03961f
C1193 VDD1.n137 VSUBS 3.52849f
C1194 VTAIL.t0 VSUBS 0.270511f
C1195 VTAIL.t1 VSUBS 0.270511f
C1196 VTAIL.n0 VSUBS 1.94022f
C1197 VTAIL.n1 VSUBS 0.94536f
C1198 VTAIL.n2 VSUBS 0.029966f
C1199 VTAIL.n3 VSUBS 0.028479f
C1200 VTAIL.n4 VSUBS 0.015303f
C1201 VTAIL.n5 VSUBS 0.036172f
C1202 VTAIL.n6 VSUBS 0.016204f
C1203 VTAIL.n7 VSUBS 0.028479f
C1204 VTAIL.n8 VSUBS 0.015303f
C1205 VTAIL.n9 VSUBS 0.036172f
C1206 VTAIL.n10 VSUBS 0.016204f
C1207 VTAIL.n11 VSUBS 0.028479f
C1208 VTAIL.n12 VSUBS 0.015754f
C1209 VTAIL.n13 VSUBS 0.036172f
C1210 VTAIL.n14 VSUBS 0.016204f
C1211 VTAIL.n15 VSUBS 0.028479f
C1212 VTAIL.n16 VSUBS 0.015303f
C1213 VTAIL.n17 VSUBS 0.036172f
C1214 VTAIL.n18 VSUBS 0.016204f
C1215 VTAIL.n19 VSUBS 0.028479f
C1216 VTAIL.n20 VSUBS 0.015303f
C1217 VTAIL.n21 VSUBS 0.027129f
C1218 VTAIL.n22 VSUBS 0.02721f
C1219 VTAIL.t10 VSUBS 0.077947f
C1220 VTAIL.n23 VSUBS 0.224547f
C1221 VTAIL.n24 VSUBS 1.40177f
C1222 VTAIL.n25 VSUBS 0.015303f
C1223 VTAIL.n26 VSUBS 0.016204f
C1224 VTAIL.n27 VSUBS 0.036172f
C1225 VTAIL.n28 VSUBS 0.036172f
C1226 VTAIL.n29 VSUBS 0.016204f
C1227 VTAIL.n30 VSUBS 0.015303f
C1228 VTAIL.n31 VSUBS 0.028479f
C1229 VTAIL.n32 VSUBS 0.028479f
C1230 VTAIL.n33 VSUBS 0.015303f
C1231 VTAIL.n34 VSUBS 0.016204f
C1232 VTAIL.n35 VSUBS 0.036172f
C1233 VTAIL.n36 VSUBS 0.036172f
C1234 VTAIL.n37 VSUBS 0.016204f
C1235 VTAIL.n38 VSUBS 0.015303f
C1236 VTAIL.n39 VSUBS 0.028479f
C1237 VTAIL.n40 VSUBS 0.028479f
C1238 VTAIL.n41 VSUBS 0.015303f
C1239 VTAIL.n42 VSUBS 0.015303f
C1240 VTAIL.n43 VSUBS 0.016204f
C1241 VTAIL.n44 VSUBS 0.036172f
C1242 VTAIL.n45 VSUBS 0.036172f
C1243 VTAIL.n46 VSUBS 0.036172f
C1244 VTAIL.n47 VSUBS 0.015754f
C1245 VTAIL.n48 VSUBS 0.015303f
C1246 VTAIL.n49 VSUBS 0.028479f
C1247 VTAIL.n50 VSUBS 0.028479f
C1248 VTAIL.n51 VSUBS 0.015303f
C1249 VTAIL.n52 VSUBS 0.016204f
C1250 VTAIL.n53 VSUBS 0.036172f
C1251 VTAIL.n54 VSUBS 0.036172f
C1252 VTAIL.n55 VSUBS 0.016204f
C1253 VTAIL.n56 VSUBS 0.015303f
C1254 VTAIL.n57 VSUBS 0.028479f
C1255 VTAIL.n58 VSUBS 0.028479f
C1256 VTAIL.n59 VSUBS 0.015303f
C1257 VTAIL.n60 VSUBS 0.016204f
C1258 VTAIL.n61 VSUBS 0.036172f
C1259 VTAIL.n62 VSUBS 0.08305f
C1260 VTAIL.n63 VSUBS 0.016204f
C1261 VTAIL.n64 VSUBS 0.015303f
C1262 VTAIL.n65 VSUBS 0.061938f
C1263 VTAIL.n66 VSUBS 0.041442f
C1264 VTAIL.n67 VSUBS 0.340544f
C1265 VTAIL.t14 VSUBS 0.270511f
C1266 VTAIL.t12 VSUBS 0.270511f
C1267 VTAIL.n68 VSUBS 1.94022f
C1268 VTAIL.n69 VSUBS 1.03456f
C1269 VTAIL.t19 VSUBS 0.270511f
C1270 VTAIL.t17 VSUBS 0.270511f
C1271 VTAIL.n70 VSUBS 1.94022f
C1272 VTAIL.n71 VSUBS 2.55583f
C1273 VTAIL.t2 VSUBS 0.270511f
C1274 VTAIL.t6 VSUBS 0.270511f
C1275 VTAIL.n72 VSUBS 1.94024f
C1276 VTAIL.n73 VSUBS 2.55582f
C1277 VTAIL.t5 VSUBS 0.270511f
C1278 VTAIL.t4 VSUBS 0.270511f
C1279 VTAIL.n74 VSUBS 1.94024f
C1280 VTAIL.n75 VSUBS 1.03454f
C1281 VTAIL.n76 VSUBS 0.029966f
C1282 VTAIL.n77 VSUBS 0.028479f
C1283 VTAIL.n78 VSUBS 0.015303f
C1284 VTAIL.n79 VSUBS 0.036172f
C1285 VTAIL.n80 VSUBS 0.016204f
C1286 VTAIL.n81 VSUBS 0.028479f
C1287 VTAIL.n82 VSUBS 0.015303f
C1288 VTAIL.n83 VSUBS 0.036172f
C1289 VTAIL.n84 VSUBS 0.016204f
C1290 VTAIL.n85 VSUBS 0.028479f
C1291 VTAIL.n86 VSUBS 0.015754f
C1292 VTAIL.n87 VSUBS 0.036172f
C1293 VTAIL.n88 VSUBS 0.015303f
C1294 VTAIL.n89 VSUBS 0.016204f
C1295 VTAIL.n90 VSUBS 0.028479f
C1296 VTAIL.n91 VSUBS 0.015303f
C1297 VTAIL.n92 VSUBS 0.036172f
C1298 VTAIL.n93 VSUBS 0.016204f
C1299 VTAIL.n94 VSUBS 0.028479f
C1300 VTAIL.n95 VSUBS 0.015303f
C1301 VTAIL.n96 VSUBS 0.027129f
C1302 VTAIL.n97 VSUBS 0.02721f
C1303 VTAIL.t8 VSUBS 0.077947f
C1304 VTAIL.n98 VSUBS 0.224547f
C1305 VTAIL.n99 VSUBS 1.40177f
C1306 VTAIL.n100 VSUBS 0.015303f
C1307 VTAIL.n101 VSUBS 0.016204f
C1308 VTAIL.n102 VSUBS 0.036172f
C1309 VTAIL.n103 VSUBS 0.036172f
C1310 VTAIL.n104 VSUBS 0.016204f
C1311 VTAIL.n105 VSUBS 0.015303f
C1312 VTAIL.n106 VSUBS 0.028479f
C1313 VTAIL.n107 VSUBS 0.028479f
C1314 VTAIL.n108 VSUBS 0.015303f
C1315 VTAIL.n109 VSUBS 0.016204f
C1316 VTAIL.n110 VSUBS 0.036172f
C1317 VTAIL.n111 VSUBS 0.036172f
C1318 VTAIL.n112 VSUBS 0.016204f
C1319 VTAIL.n113 VSUBS 0.015303f
C1320 VTAIL.n114 VSUBS 0.028479f
C1321 VTAIL.n115 VSUBS 0.028479f
C1322 VTAIL.n116 VSUBS 0.015303f
C1323 VTAIL.n117 VSUBS 0.016204f
C1324 VTAIL.n118 VSUBS 0.036172f
C1325 VTAIL.n119 VSUBS 0.036172f
C1326 VTAIL.n120 VSUBS 0.036172f
C1327 VTAIL.n121 VSUBS 0.015754f
C1328 VTAIL.n122 VSUBS 0.015303f
C1329 VTAIL.n123 VSUBS 0.028479f
C1330 VTAIL.n124 VSUBS 0.028479f
C1331 VTAIL.n125 VSUBS 0.015303f
C1332 VTAIL.n126 VSUBS 0.016204f
C1333 VTAIL.n127 VSUBS 0.036172f
C1334 VTAIL.n128 VSUBS 0.036172f
C1335 VTAIL.n129 VSUBS 0.016204f
C1336 VTAIL.n130 VSUBS 0.015303f
C1337 VTAIL.n131 VSUBS 0.028479f
C1338 VTAIL.n132 VSUBS 0.028479f
C1339 VTAIL.n133 VSUBS 0.015303f
C1340 VTAIL.n134 VSUBS 0.016204f
C1341 VTAIL.n135 VSUBS 0.036172f
C1342 VTAIL.n136 VSUBS 0.08305f
C1343 VTAIL.n137 VSUBS 0.016204f
C1344 VTAIL.n138 VSUBS 0.015303f
C1345 VTAIL.n139 VSUBS 0.061938f
C1346 VTAIL.n140 VSUBS 0.041442f
C1347 VTAIL.n141 VSUBS 0.340544f
C1348 VTAIL.t16 VSUBS 0.270511f
C1349 VTAIL.t15 VSUBS 0.270511f
C1350 VTAIL.n142 VSUBS 1.94024f
C1351 VTAIL.n143 VSUBS 0.985889f
C1352 VTAIL.t11 VSUBS 0.270511f
C1353 VTAIL.t13 VSUBS 0.270511f
C1354 VTAIL.n144 VSUBS 1.94024f
C1355 VTAIL.n145 VSUBS 1.03454f
C1356 VTAIL.n146 VSUBS 0.029966f
C1357 VTAIL.n147 VSUBS 0.028479f
C1358 VTAIL.n148 VSUBS 0.015303f
C1359 VTAIL.n149 VSUBS 0.036172f
C1360 VTAIL.n150 VSUBS 0.016204f
C1361 VTAIL.n151 VSUBS 0.028479f
C1362 VTAIL.n152 VSUBS 0.015303f
C1363 VTAIL.n153 VSUBS 0.036172f
C1364 VTAIL.n154 VSUBS 0.016204f
C1365 VTAIL.n155 VSUBS 0.028479f
C1366 VTAIL.n156 VSUBS 0.015754f
C1367 VTAIL.n157 VSUBS 0.036172f
C1368 VTAIL.n158 VSUBS 0.015303f
C1369 VTAIL.n159 VSUBS 0.016204f
C1370 VTAIL.n160 VSUBS 0.028479f
C1371 VTAIL.n161 VSUBS 0.015303f
C1372 VTAIL.n162 VSUBS 0.036172f
C1373 VTAIL.n163 VSUBS 0.016204f
C1374 VTAIL.n164 VSUBS 0.028479f
C1375 VTAIL.n165 VSUBS 0.015303f
C1376 VTAIL.n166 VSUBS 0.027129f
C1377 VTAIL.n167 VSUBS 0.02721f
C1378 VTAIL.t18 VSUBS 0.077947f
C1379 VTAIL.n168 VSUBS 0.224547f
C1380 VTAIL.n169 VSUBS 1.40177f
C1381 VTAIL.n170 VSUBS 0.015303f
C1382 VTAIL.n171 VSUBS 0.016204f
C1383 VTAIL.n172 VSUBS 0.036172f
C1384 VTAIL.n173 VSUBS 0.036172f
C1385 VTAIL.n174 VSUBS 0.016204f
C1386 VTAIL.n175 VSUBS 0.015303f
C1387 VTAIL.n176 VSUBS 0.028479f
C1388 VTAIL.n177 VSUBS 0.028479f
C1389 VTAIL.n178 VSUBS 0.015303f
C1390 VTAIL.n179 VSUBS 0.016204f
C1391 VTAIL.n180 VSUBS 0.036172f
C1392 VTAIL.n181 VSUBS 0.036172f
C1393 VTAIL.n182 VSUBS 0.016204f
C1394 VTAIL.n183 VSUBS 0.015303f
C1395 VTAIL.n184 VSUBS 0.028479f
C1396 VTAIL.n185 VSUBS 0.028479f
C1397 VTAIL.n186 VSUBS 0.015303f
C1398 VTAIL.n187 VSUBS 0.016204f
C1399 VTAIL.n188 VSUBS 0.036172f
C1400 VTAIL.n189 VSUBS 0.036172f
C1401 VTAIL.n190 VSUBS 0.036172f
C1402 VTAIL.n191 VSUBS 0.015754f
C1403 VTAIL.n192 VSUBS 0.015303f
C1404 VTAIL.n193 VSUBS 0.028479f
C1405 VTAIL.n194 VSUBS 0.028479f
C1406 VTAIL.n195 VSUBS 0.015303f
C1407 VTAIL.n196 VSUBS 0.016204f
C1408 VTAIL.n197 VSUBS 0.036172f
C1409 VTAIL.n198 VSUBS 0.036172f
C1410 VTAIL.n199 VSUBS 0.016204f
C1411 VTAIL.n200 VSUBS 0.015303f
C1412 VTAIL.n201 VSUBS 0.028479f
C1413 VTAIL.n202 VSUBS 0.028479f
C1414 VTAIL.n203 VSUBS 0.015303f
C1415 VTAIL.n204 VSUBS 0.016204f
C1416 VTAIL.n205 VSUBS 0.036172f
C1417 VTAIL.n206 VSUBS 0.08305f
C1418 VTAIL.n207 VSUBS 0.016204f
C1419 VTAIL.n208 VSUBS 0.015303f
C1420 VTAIL.n209 VSUBS 0.061938f
C1421 VTAIL.n210 VSUBS 0.041442f
C1422 VTAIL.n211 VSUBS 1.72694f
C1423 VTAIL.n212 VSUBS 0.029966f
C1424 VTAIL.n213 VSUBS 0.028479f
C1425 VTAIL.n214 VSUBS 0.015303f
C1426 VTAIL.n215 VSUBS 0.036172f
C1427 VTAIL.n216 VSUBS 0.016204f
C1428 VTAIL.n217 VSUBS 0.028479f
C1429 VTAIL.n218 VSUBS 0.015303f
C1430 VTAIL.n219 VSUBS 0.036172f
C1431 VTAIL.n220 VSUBS 0.016204f
C1432 VTAIL.n221 VSUBS 0.028479f
C1433 VTAIL.n222 VSUBS 0.015754f
C1434 VTAIL.n223 VSUBS 0.036172f
C1435 VTAIL.n224 VSUBS 0.016204f
C1436 VTAIL.n225 VSUBS 0.028479f
C1437 VTAIL.n226 VSUBS 0.015303f
C1438 VTAIL.n227 VSUBS 0.036172f
C1439 VTAIL.n228 VSUBS 0.016204f
C1440 VTAIL.n229 VSUBS 0.028479f
C1441 VTAIL.n230 VSUBS 0.015303f
C1442 VTAIL.n231 VSUBS 0.027129f
C1443 VTAIL.n232 VSUBS 0.02721f
C1444 VTAIL.t7 VSUBS 0.077947f
C1445 VTAIL.n233 VSUBS 0.224547f
C1446 VTAIL.n234 VSUBS 1.40177f
C1447 VTAIL.n235 VSUBS 0.015303f
C1448 VTAIL.n236 VSUBS 0.016204f
C1449 VTAIL.n237 VSUBS 0.036172f
C1450 VTAIL.n238 VSUBS 0.036172f
C1451 VTAIL.n239 VSUBS 0.016204f
C1452 VTAIL.n240 VSUBS 0.015303f
C1453 VTAIL.n241 VSUBS 0.028479f
C1454 VTAIL.n242 VSUBS 0.028479f
C1455 VTAIL.n243 VSUBS 0.015303f
C1456 VTAIL.n244 VSUBS 0.016204f
C1457 VTAIL.n245 VSUBS 0.036172f
C1458 VTAIL.n246 VSUBS 0.036172f
C1459 VTAIL.n247 VSUBS 0.016204f
C1460 VTAIL.n248 VSUBS 0.015303f
C1461 VTAIL.n249 VSUBS 0.028479f
C1462 VTAIL.n250 VSUBS 0.028479f
C1463 VTAIL.n251 VSUBS 0.015303f
C1464 VTAIL.n252 VSUBS 0.015303f
C1465 VTAIL.n253 VSUBS 0.016204f
C1466 VTAIL.n254 VSUBS 0.036172f
C1467 VTAIL.n255 VSUBS 0.036172f
C1468 VTAIL.n256 VSUBS 0.036172f
C1469 VTAIL.n257 VSUBS 0.015754f
C1470 VTAIL.n258 VSUBS 0.015303f
C1471 VTAIL.n259 VSUBS 0.028479f
C1472 VTAIL.n260 VSUBS 0.028479f
C1473 VTAIL.n261 VSUBS 0.015303f
C1474 VTAIL.n262 VSUBS 0.016204f
C1475 VTAIL.n263 VSUBS 0.036172f
C1476 VTAIL.n264 VSUBS 0.036172f
C1477 VTAIL.n265 VSUBS 0.016204f
C1478 VTAIL.n266 VSUBS 0.015303f
C1479 VTAIL.n267 VSUBS 0.028479f
C1480 VTAIL.n268 VSUBS 0.028479f
C1481 VTAIL.n269 VSUBS 0.015303f
C1482 VTAIL.n270 VSUBS 0.016204f
C1483 VTAIL.n271 VSUBS 0.036172f
C1484 VTAIL.n272 VSUBS 0.08305f
C1485 VTAIL.n273 VSUBS 0.016204f
C1486 VTAIL.n274 VSUBS 0.015303f
C1487 VTAIL.n275 VSUBS 0.061938f
C1488 VTAIL.n276 VSUBS 0.041442f
C1489 VTAIL.n277 VSUBS 1.72694f
C1490 VTAIL.t3 VSUBS 0.270511f
C1491 VTAIL.t9 VSUBS 0.270511f
C1492 VTAIL.n278 VSUBS 1.94022f
C1493 VTAIL.n279 VSUBS 0.891566f
C1494 VP.n0 VSUBS 0.043868f
C1495 VP.t0 VSUBS 2.16874f
C1496 VP.n1 VSUBS 0.04653f
C1497 VP.n2 VSUBS 0.033275f
C1498 VP.t4 VSUBS 2.16874f
C1499 VP.n3 VSUBS 0.030478f
C1500 VP.n4 VSUBS 0.033275f
C1501 VP.t9 VSUBS 2.16874f
C1502 VP.n5 VSUBS 0.061401f
C1503 VP.n6 VSUBS 0.033275f
C1504 VP.t2 VSUBS 2.16874f
C1505 VP.n7 VSUBS 0.773996f
C1506 VP.n8 VSUBS 0.033275f
C1507 VP.n9 VSUBS 0.055004f
C1508 VP.n10 VSUBS 0.043868f
C1509 VP.t6 VSUBS 2.16874f
C1510 VP.n11 VSUBS 0.04653f
C1511 VP.n12 VSUBS 0.033275f
C1512 VP.t1 VSUBS 2.16874f
C1513 VP.n13 VSUBS 0.030478f
C1514 VP.n14 VSUBS 0.033275f
C1515 VP.t7 VSUBS 2.16874f
C1516 VP.n15 VSUBS 0.061401f
C1517 VP.n16 VSUBS 0.033275f
C1518 VP.t8 VSUBS 2.16874f
C1519 VP.n17 VSUBS 0.842619f
C1520 VP.t5 VSUBS 2.32946f
C1521 VP.n18 VSUBS 0.859649f
C1522 VP.n19 VSUBS 0.248761f
C1523 VP.n20 VSUBS 0.035508f
C1524 VP.n21 VSUBS 0.06657f
C1525 VP.n22 VSUBS 0.030478f
C1526 VP.n23 VSUBS 0.033275f
C1527 VP.n24 VSUBS 0.033275f
C1528 VP.n25 VSUBS 0.033275f
C1529 VP.n26 VSUBS 0.046475f
C1530 VP.n27 VSUBS 0.773996f
C1531 VP.n28 VSUBS 0.046475f
C1532 VP.n29 VSUBS 0.061401f
C1533 VP.n30 VSUBS 0.033275f
C1534 VP.n31 VSUBS 0.033275f
C1535 VP.n32 VSUBS 0.033275f
C1536 VP.n33 VSUBS 0.06657f
C1537 VP.n34 VSUBS 0.035508f
C1538 VP.n35 VSUBS 0.773996f
C1539 VP.n36 VSUBS 0.057441f
C1540 VP.n37 VSUBS 0.033275f
C1541 VP.n38 VSUBS 0.033275f
C1542 VP.n39 VSUBS 0.033275f
C1543 VP.n40 VSUBS 0.050212f
C1544 VP.n41 VSUBS 0.055004f
C1545 VP.n42 VSUBS 0.87352f
C1546 VP.n43 VSUBS 1.82777f
C1547 VP.t3 VSUBS 2.16874f
C1548 VP.n44 VSUBS 0.87352f
C1549 VP.n45 VSUBS 1.85185f
C1550 VP.n46 VSUBS 0.043868f
C1551 VP.n47 VSUBS 0.033275f
C1552 VP.n48 VSUBS 0.050212f
C1553 VP.n49 VSUBS 0.04653f
C1554 VP.n50 VSUBS 0.057441f
C1555 VP.n51 VSUBS 0.033275f
C1556 VP.n52 VSUBS 0.033275f
C1557 VP.n53 VSUBS 0.035508f
C1558 VP.n54 VSUBS 0.06657f
C1559 VP.n55 VSUBS 0.030478f
C1560 VP.n56 VSUBS 0.033275f
C1561 VP.n57 VSUBS 0.033275f
C1562 VP.n58 VSUBS 0.033275f
C1563 VP.n59 VSUBS 0.046475f
C1564 VP.n60 VSUBS 0.773996f
C1565 VP.n61 VSUBS 0.046475f
C1566 VP.n62 VSUBS 0.061401f
C1567 VP.n63 VSUBS 0.033275f
C1568 VP.n64 VSUBS 0.033275f
C1569 VP.n65 VSUBS 0.033275f
C1570 VP.n66 VSUBS 0.06657f
C1571 VP.n67 VSUBS 0.035508f
C1572 VP.n68 VSUBS 0.773996f
C1573 VP.n69 VSUBS 0.057441f
C1574 VP.n70 VSUBS 0.033275f
C1575 VP.n71 VSUBS 0.033275f
C1576 VP.n72 VSUBS 0.033275f
C1577 VP.n73 VSUBS 0.050212f
C1578 VP.n74 VSUBS 0.055004f
C1579 VP.n75 VSUBS 0.87352f
C1580 VP.n76 VSUBS 0.040997f
.ends

