* NGSPICE file created from diff_pair_sample_0128.ext - technology: sky130A

.subckt diff_pair_sample_0128 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VP.t0 VDD1.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=3.6426 pd=19.46 as=1.5411 ps=9.67 w=9.34 l=3.69
X1 VTAIL.t2 VN.t0 VDD2.t7 B.t2 sky130_fd_pr__nfet_01v8 ad=3.6426 pd=19.46 as=1.5411 ps=9.67 w=9.34 l=3.69
X2 B.t21 B.t19 B.t20 B.t9 sky130_fd_pr__nfet_01v8 ad=3.6426 pd=19.46 as=0 ps=0 w=9.34 l=3.69
X3 B.t18 B.t16 B.t17 B.t13 sky130_fd_pr__nfet_01v8 ad=3.6426 pd=19.46 as=0 ps=0 w=9.34 l=3.69
X4 VDD1.t5 VP.t1 VTAIL.t14 B.t6 sky130_fd_pr__nfet_01v8 ad=1.5411 pd=9.67 as=1.5411 ps=9.67 w=9.34 l=3.69
X5 VDD2.t6 VN.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.5411 pd=9.67 as=1.5411 ps=9.67 w=9.34 l=3.69
X6 VTAIL.t13 VP.t2 VDD1.t4 B.t5 sky130_fd_pr__nfet_01v8 ad=3.6426 pd=19.46 as=1.5411 ps=9.67 w=9.34 l=3.69
X7 VTAIL.t12 VP.t3 VDD1.t3 B.t7 sky130_fd_pr__nfet_01v8 ad=1.5411 pd=9.67 as=1.5411 ps=9.67 w=9.34 l=3.69
X8 VDD1.t2 VP.t4 VTAIL.t11 B.t0 sky130_fd_pr__nfet_01v8 ad=1.5411 pd=9.67 as=1.5411 ps=9.67 w=9.34 l=3.69
X9 VDD1.t1 VP.t5 VTAIL.t10 B.t4 sky130_fd_pr__nfet_01v8 ad=1.5411 pd=9.67 as=3.6426 ps=19.46 w=9.34 l=3.69
X10 VTAIL.t5 VN.t2 VDD2.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=3.6426 pd=19.46 as=1.5411 ps=9.67 w=9.34 l=3.69
X11 VDD2.t4 VN.t3 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.5411 pd=9.67 as=3.6426 ps=19.46 w=9.34 l=3.69
X12 VDD1.t7 VP.t6 VTAIL.t9 B.t1 sky130_fd_pr__nfet_01v8 ad=1.5411 pd=9.67 as=3.6426 ps=19.46 w=9.34 l=3.69
X13 VDD2.t3 VN.t4 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.5411 pd=9.67 as=3.6426 ps=19.46 w=9.34 l=3.69
X14 VTAIL.t8 VP.t7 VDD1.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=1.5411 pd=9.67 as=1.5411 ps=9.67 w=9.34 l=3.69
X15 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=3.6426 pd=19.46 as=0 ps=0 w=9.34 l=3.69
X16 VTAIL.t3 VN.t5 VDD2.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=1.5411 pd=9.67 as=1.5411 ps=9.67 w=9.34 l=3.69
X17 VTAIL.t7 VN.t6 VDD2.t1 B.t7 sky130_fd_pr__nfet_01v8 ad=1.5411 pd=9.67 as=1.5411 ps=9.67 w=9.34 l=3.69
X18 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=3.6426 pd=19.46 as=0 ps=0 w=9.34 l=3.69
X19 VDD2.t0 VN.t7 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=1.5411 pd=9.67 as=1.5411 ps=9.67 w=9.34 l=3.69
R0 VP.n25 VP.n24 161.3
R1 VP.n26 VP.n21 161.3
R2 VP.n28 VP.n27 161.3
R3 VP.n29 VP.n20 161.3
R4 VP.n31 VP.n30 161.3
R5 VP.n32 VP.n19 161.3
R6 VP.n34 VP.n33 161.3
R7 VP.n35 VP.n18 161.3
R8 VP.n38 VP.n37 161.3
R9 VP.n39 VP.n17 161.3
R10 VP.n41 VP.n40 161.3
R11 VP.n42 VP.n16 161.3
R12 VP.n44 VP.n43 161.3
R13 VP.n45 VP.n15 161.3
R14 VP.n47 VP.n46 161.3
R15 VP.n48 VP.n14 161.3
R16 VP.n50 VP.n49 161.3
R17 VP.n93 VP.n92 161.3
R18 VP.n91 VP.n1 161.3
R19 VP.n90 VP.n89 161.3
R20 VP.n88 VP.n2 161.3
R21 VP.n87 VP.n86 161.3
R22 VP.n85 VP.n3 161.3
R23 VP.n84 VP.n83 161.3
R24 VP.n82 VP.n4 161.3
R25 VP.n81 VP.n80 161.3
R26 VP.n78 VP.n5 161.3
R27 VP.n77 VP.n76 161.3
R28 VP.n75 VP.n6 161.3
R29 VP.n74 VP.n73 161.3
R30 VP.n72 VP.n7 161.3
R31 VP.n71 VP.n70 161.3
R32 VP.n69 VP.n8 161.3
R33 VP.n68 VP.n67 161.3
R34 VP.n65 VP.n9 161.3
R35 VP.n64 VP.n63 161.3
R36 VP.n62 VP.n10 161.3
R37 VP.n61 VP.n60 161.3
R38 VP.n59 VP.n11 161.3
R39 VP.n58 VP.n57 161.3
R40 VP.n56 VP.n12 161.3
R41 VP.n55 VP.n54 161.3
R42 VP.n22 VP.t0 92.5413
R43 VP.n53 VP.n52 88.77
R44 VP.n94 VP.n0 88.77
R45 VP.n51 VP.n13 88.77
R46 VP.n23 VP.n22 74.7511
R47 VP.n53 VP.t2 61.0016
R48 VP.n66 VP.t4 61.0016
R49 VP.n79 VP.t7 61.0016
R50 VP.n0 VP.t6 61.0016
R51 VP.n13 VP.t5 61.0016
R52 VP.n36 VP.t3 61.0016
R53 VP.n23 VP.t1 61.0016
R54 VP.n52 VP.n51 53.9844
R55 VP.n60 VP.n59 42.5146
R56 VP.n86 VP.n2 42.5146
R57 VP.n43 VP.n15 42.5146
R58 VP.n73 VP.n72 40.577
R59 VP.n73 VP.n6 40.577
R60 VP.n30 VP.n19 40.577
R61 VP.n30 VP.n29 40.577
R62 VP.n60 VP.n10 38.6395
R63 VP.n86 VP.n85 38.6395
R64 VP.n43 VP.n42 38.6395
R65 VP.n54 VP.n12 24.5923
R66 VP.n58 VP.n12 24.5923
R67 VP.n59 VP.n58 24.5923
R68 VP.n64 VP.n10 24.5923
R69 VP.n65 VP.n64 24.5923
R70 VP.n67 VP.n8 24.5923
R71 VP.n71 VP.n8 24.5923
R72 VP.n72 VP.n71 24.5923
R73 VP.n77 VP.n6 24.5923
R74 VP.n78 VP.n77 24.5923
R75 VP.n80 VP.n78 24.5923
R76 VP.n84 VP.n4 24.5923
R77 VP.n85 VP.n84 24.5923
R78 VP.n90 VP.n2 24.5923
R79 VP.n91 VP.n90 24.5923
R80 VP.n92 VP.n91 24.5923
R81 VP.n47 VP.n15 24.5923
R82 VP.n48 VP.n47 24.5923
R83 VP.n49 VP.n48 24.5923
R84 VP.n34 VP.n19 24.5923
R85 VP.n35 VP.n34 24.5923
R86 VP.n37 VP.n35 24.5923
R87 VP.n41 VP.n17 24.5923
R88 VP.n42 VP.n41 24.5923
R89 VP.n24 VP.n21 24.5923
R90 VP.n28 VP.n21 24.5923
R91 VP.n29 VP.n28 24.5923
R92 VP.n66 VP.n65 24.1005
R93 VP.n79 VP.n4 24.1005
R94 VP.n36 VP.n17 24.1005
R95 VP.n25 VP.n22 3.41204
R96 VP.n54 VP.n53 1.47601
R97 VP.n92 VP.n0 1.47601
R98 VP.n49 VP.n13 1.47601
R99 VP.n67 VP.n66 0.492337
R100 VP.n80 VP.n79 0.492337
R101 VP.n37 VP.n36 0.492337
R102 VP.n24 VP.n23 0.492337
R103 VP.n51 VP.n50 0.354861
R104 VP.n55 VP.n52 0.354861
R105 VP.n94 VP.n93 0.354861
R106 VP VP.n94 0.267071
R107 VP.n26 VP.n25 0.189894
R108 VP.n27 VP.n26 0.189894
R109 VP.n27 VP.n20 0.189894
R110 VP.n31 VP.n20 0.189894
R111 VP.n32 VP.n31 0.189894
R112 VP.n33 VP.n32 0.189894
R113 VP.n33 VP.n18 0.189894
R114 VP.n38 VP.n18 0.189894
R115 VP.n39 VP.n38 0.189894
R116 VP.n40 VP.n39 0.189894
R117 VP.n40 VP.n16 0.189894
R118 VP.n44 VP.n16 0.189894
R119 VP.n45 VP.n44 0.189894
R120 VP.n46 VP.n45 0.189894
R121 VP.n46 VP.n14 0.189894
R122 VP.n50 VP.n14 0.189894
R123 VP.n56 VP.n55 0.189894
R124 VP.n57 VP.n56 0.189894
R125 VP.n57 VP.n11 0.189894
R126 VP.n61 VP.n11 0.189894
R127 VP.n62 VP.n61 0.189894
R128 VP.n63 VP.n62 0.189894
R129 VP.n63 VP.n9 0.189894
R130 VP.n68 VP.n9 0.189894
R131 VP.n69 VP.n68 0.189894
R132 VP.n70 VP.n69 0.189894
R133 VP.n70 VP.n7 0.189894
R134 VP.n74 VP.n7 0.189894
R135 VP.n75 VP.n74 0.189894
R136 VP.n76 VP.n75 0.189894
R137 VP.n76 VP.n5 0.189894
R138 VP.n81 VP.n5 0.189894
R139 VP.n82 VP.n81 0.189894
R140 VP.n83 VP.n82 0.189894
R141 VP.n83 VP.n3 0.189894
R142 VP.n87 VP.n3 0.189894
R143 VP.n88 VP.n87 0.189894
R144 VP.n89 VP.n88 0.189894
R145 VP.n89 VP.n1 0.189894
R146 VP.n93 VP.n1 0.189894
R147 VDD1 VDD1.n0 66.7324
R148 VDD1.n3 VDD1.n2 66.6187
R149 VDD1.n3 VDD1.n1 66.6187
R150 VDD1.n5 VDD1.n4 64.9413
R151 VDD1.n5 VDD1.n3 47.9449
R152 VDD1.n4 VDD1.t3 2.12041
R153 VDD1.n4 VDD1.t1 2.12041
R154 VDD1.n0 VDD1.t6 2.12041
R155 VDD1.n0 VDD1.t5 2.12041
R156 VDD1.n2 VDD1.t0 2.12041
R157 VDD1.n2 VDD1.t7 2.12041
R158 VDD1.n1 VDD1.t4 2.12041
R159 VDD1.n1 VDD1.t2 2.12041
R160 VDD1 VDD1.n5 1.67507
R161 VTAIL.n402 VTAIL.n358 289.615
R162 VTAIL.n46 VTAIL.n2 289.615
R163 VTAIL.n96 VTAIL.n52 289.615
R164 VTAIL.n148 VTAIL.n104 289.615
R165 VTAIL.n352 VTAIL.n308 289.615
R166 VTAIL.n300 VTAIL.n256 289.615
R167 VTAIL.n250 VTAIL.n206 289.615
R168 VTAIL.n198 VTAIL.n154 289.615
R169 VTAIL.n375 VTAIL.n374 185
R170 VTAIL.n377 VTAIL.n376 185
R171 VTAIL.n370 VTAIL.n369 185
R172 VTAIL.n383 VTAIL.n382 185
R173 VTAIL.n385 VTAIL.n384 185
R174 VTAIL.n366 VTAIL.n365 185
R175 VTAIL.n392 VTAIL.n391 185
R176 VTAIL.n393 VTAIL.n364 185
R177 VTAIL.n395 VTAIL.n394 185
R178 VTAIL.n362 VTAIL.n361 185
R179 VTAIL.n401 VTAIL.n400 185
R180 VTAIL.n403 VTAIL.n402 185
R181 VTAIL.n19 VTAIL.n18 185
R182 VTAIL.n21 VTAIL.n20 185
R183 VTAIL.n14 VTAIL.n13 185
R184 VTAIL.n27 VTAIL.n26 185
R185 VTAIL.n29 VTAIL.n28 185
R186 VTAIL.n10 VTAIL.n9 185
R187 VTAIL.n36 VTAIL.n35 185
R188 VTAIL.n37 VTAIL.n8 185
R189 VTAIL.n39 VTAIL.n38 185
R190 VTAIL.n6 VTAIL.n5 185
R191 VTAIL.n45 VTAIL.n44 185
R192 VTAIL.n47 VTAIL.n46 185
R193 VTAIL.n69 VTAIL.n68 185
R194 VTAIL.n71 VTAIL.n70 185
R195 VTAIL.n64 VTAIL.n63 185
R196 VTAIL.n77 VTAIL.n76 185
R197 VTAIL.n79 VTAIL.n78 185
R198 VTAIL.n60 VTAIL.n59 185
R199 VTAIL.n86 VTAIL.n85 185
R200 VTAIL.n87 VTAIL.n58 185
R201 VTAIL.n89 VTAIL.n88 185
R202 VTAIL.n56 VTAIL.n55 185
R203 VTAIL.n95 VTAIL.n94 185
R204 VTAIL.n97 VTAIL.n96 185
R205 VTAIL.n121 VTAIL.n120 185
R206 VTAIL.n123 VTAIL.n122 185
R207 VTAIL.n116 VTAIL.n115 185
R208 VTAIL.n129 VTAIL.n128 185
R209 VTAIL.n131 VTAIL.n130 185
R210 VTAIL.n112 VTAIL.n111 185
R211 VTAIL.n138 VTAIL.n137 185
R212 VTAIL.n139 VTAIL.n110 185
R213 VTAIL.n141 VTAIL.n140 185
R214 VTAIL.n108 VTAIL.n107 185
R215 VTAIL.n147 VTAIL.n146 185
R216 VTAIL.n149 VTAIL.n148 185
R217 VTAIL.n353 VTAIL.n352 185
R218 VTAIL.n351 VTAIL.n350 185
R219 VTAIL.n312 VTAIL.n311 185
R220 VTAIL.n316 VTAIL.n314 185
R221 VTAIL.n345 VTAIL.n344 185
R222 VTAIL.n343 VTAIL.n342 185
R223 VTAIL.n318 VTAIL.n317 185
R224 VTAIL.n337 VTAIL.n336 185
R225 VTAIL.n335 VTAIL.n334 185
R226 VTAIL.n322 VTAIL.n321 185
R227 VTAIL.n329 VTAIL.n328 185
R228 VTAIL.n327 VTAIL.n326 185
R229 VTAIL.n301 VTAIL.n300 185
R230 VTAIL.n299 VTAIL.n298 185
R231 VTAIL.n260 VTAIL.n259 185
R232 VTAIL.n264 VTAIL.n262 185
R233 VTAIL.n293 VTAIL.n292 185
R234 VTAIL.n291 VTAIL.n290 185
R235 VTAIL.n266 VTAIL.n265 185
R236 VTAIL.n285 VTAIL.n284 185
R237 VTAIL.n283 VTAIL.n282 185
R238 VTAIL.n270 VTAIL.n269 185
R239 VTAIL.n277 VTAIL.n276 185
R240 VTAIL.n275 VTAIL.n274 185
R241 VTAIL.n251 VTAIL.n250 185
R242 VTAIL.n249 VTAIL.n248 185
R243 VTAIL.n210 VTAIL.n209 185
R244 VTAIL.n214 VTAIL.n212 185
R245 VTAIL.n243 VTAIL.n242 185
R246 VTAIL.n241 VTAIL.n240 185
R247 VTAIL.n216 VTAIL.n215 185
R248 VTAIL.n235 VTAIL.n234 185
R249 VTAIL.n233 VTAIL.n232 185
R250 VTAIL.n220 VTAIL.n219 185
R251 VTAIL.n227 VTAIL.n226 185
R252 VTAIL.n225 VTAIL.n224 185
R253 VTAIL.n199 VTAIL.n198 185
R254 VTAIL.n197 VTAIL.n196 185
R255 VTAIL.n158 VTAIL.n157 185
R256 VTAIL.n162 VTAIL.n160 185
R257 VTAIL.n191 VTAIL.n190 185
R258 VTAIL.n189 VTAIL.n188 185
R259 VTAIL.n164 VTAIL.n163 185
R260 VTAIL.n183 VTAIL.n182 185
R261 VTAIL.n181 VTAIL.n180 185
R262 VTAIL.n168 VTAIL.n167 185
R263 VTAIL.n175 VTAIL.n174 185
R264 VTAIL.n173 VTAIL.n172 185
R265 VTAIL.n373 VTAIL.t4 149.524
R266 VTAIL.n17 VTAIL.t2 149.524
R267 VTAIL.n67 VTAIL.t9 149.524
R268 VTAIL.n119 VTAIL.t13 149.524
R269 VTAIL.n325 VTAIL.t10 149.524
R270 VTAIL.n273 VTAIL.t15 149.524
R271 VTAIL.n223 VTAIL.t1 149.524
R272 VTAIL.n171 VTAIL.t5 149.524
R273 VTAIL.n376 VTAIL.n375 104.615
R274 VTAIL.n376 VTAIL.n369 104.615
R275 VTAIL.n383 VTAIL.n369 104.615
R276 VTAIL.n384 VTAIL.n383 104.615
R277 VTAIL.n384 VTAIL.n365 104.615
R278 VTAIL.n392 VTAIL.n365 104.615
R279 VTAIL.n393 VTAIL.n392 104.615
R280 VTAIL.n394 VTAIL.n393 104.615
R281 VTAIL.n394 VTAIL.n361 104.615
R282 VTAIL.n401 VTAIL.n361 104.615
R283 VTAIL.n402 VTAIL.n401 104.615
R284 VTAIL.n20 VTAIL.n19 104.615
R285 VTAIL.n20 VTAIL.n13 104.615
R286 VTAIL.n27 VTAIL.n13 104.615
R287 VTAIL.n28 VTAIL.n27 104.615
R288 VTAIL.n28 VTAIL.n9 104.615
R289 VTAIL.n36 VTAIL.n9 104.615
R290 VTAIL.n37 VTAIL.n36 104.615
R291 VTAIL.n38 VTAIL.n37 104.615
R292 VTAIL.n38 VTAIL.n5 104.615
R293 VTAIL.n45 VTAIL.n5 104.615
R294 VTAIL.n46 VTAIL.n45 104.615
R295 VTAIL.n70 VTAIL.n69 104.615
R296 VTAIL.n70 VTAIL.n63 104.615
R297 VTAIL.n77 VTAIL.n63 104.615
R298 VTAIL.n78 VTAIL.n77 104.615
R299 VTAIL.n78 VTAIL.n59 104.615
R300 VTAIL.n86 VTAIL.n59 104.615
R301 VTAIL.n87 VTAIL.n86 104.615
R302 VTAIL.n88 VTAIL.n87 104.615
R303 VTAIL.n88 VTAIL.n55 104.615
R304 VTAIL.n95 VTAIL.n55 104.615
R305 VTAIL.n96 VTAIL.n95 104.615
R306 VTAIL.n122 VTAIL.n121 104.615
R307 VTAIL.n122 VTAIL.n115 104.615
R308 VTAIL.n129 VTAIL.n115 104.615
R309 VTAIL.n130 VTAIL.n129 104.615
R310 VTAIL.n130 VTAIL.n111 104.615
R311 VTAIL.n138 VTAIL.n111 104.615
R312 VTAIL.n139 VTAIL.n138 104.615
R313 VTAIL.n140 VTAIL.n139 104.615
R314 VTAIL.n140 VTAIL.n107 104.615
R315 VTAIL.n147 VTAIL.n107 104.615
R316 VTAIL.n148 VTAIL.n147 104.615
R317 VTAIL.n352 VTAIL.n351 104.615
R318 VTAIL.n351 VTAIL.n311 104.615
R319 VTAIL.n316 VTAIL.n311 104.615
R320 VTAIL.n344 VTAIL.n316 104.615
R321 VTAIL.n344 VTAIL.n343 104.615
R322 VTAIL.n343 VTAIL.n317 104.615
R323 VTAIL.n336 VTAIL.n317 104.615
R324 VTAIL.n336 VTAIL.n335 104.615
R325 VTAIL.n335 VTAIL.n321 104.615
R326 VTAIL.n328 VTAIL.n321 104.615
R327 VTAIL.n328 VTAIL.n327 104.615
R328 VTAIL.n300 VTAIL.n299 104.615
R329 VTAIL.n299 VTAIL.n259 104.615
R330 VTAIL.n264 VTAIL.n259 104.615
R331 VTAIL.n292 VTAIL.n264 104.615
R332 VTAIL.n292 VTAIL.n291 104.615
R333 VTAIL.n291 VTAIL.n265 104.615
R334 VTAIL.n284 VTAIL.n265 104.615
R335 VTAIL.n284 VTAIL.n283 104.615
R336 VTAIL.n283 VTAIL.n269 104.615
R337 VTAIL.n276 VTAIL.n269 104.615
R338 VTAIL.n276 VTAIL.n275 104.615
R339 VTAIL.n250 VTAIL.n249 104.615
R340 VTAIL.n249 VTAIL.n209 104.615
R341 VTAIL.n214 VTAIL.n209 104.615
R342 VTAIL.n242 VTAIL.n214 104.615
R343 VTAIL.n242 VTAIL.n241 104.615
R344 VTAIL.n241 VTAIL.n215 104.615
R345 VTAIL.n234 VTAIL.n215 104.615
R346 VTAIL.n234 VTAIL.n233 104.615
R347 VTAIL.n233 VTAIL.n219 104.615
R348 VTAIL.n226 VTAIL.n219 104.615
R349 VTAIL.n226 VTAIL.n225 104.615
R350 VTAIL.n198 VTAIL.n197 104.615
R351 VTAIL.n197 VTAIL.n157 104.615
R352 VTAIL.n162 VTAIL.n157 104.615
R353 VTAIL.n190 VTAIL.n162 104.615
R354 VTAIL.n190 VTAIL.n189 104.615
R355 VTAIL.n189 VTAIL.n163 104.615
R356 VTAIL.n182 VTAIL.n163 104.615
R357 VTAIL.n182 VTAIL.n181 104.615
R358 VTAIL.n181 VTAIL.n167 104.615
R359 VTAIL.n174 VTAIL.n167 104.615
R360 VTAIL.n174 VTAIL.n173 104.615
R361 VTAIL.n375 VTAIL.t4 52.3082
R362 VTAIL.n19 VTAIL.t2 52.3082
R363 VTAIL.n69 VTAIL.t9 52.3082
R364 VTAIL.n121 VTAIL.t13 52.3082
R365 VTAIL.n327 VTAIL.t10 52.3082
R366 VTAIL.n275 VTAIL.t15 52.3082
R367 VTAIL.n225 VTAIL.t1 52.3082
R368 VTAIL.n173 VTAIL.t5 52.3082
R369 VTAIL.n307 VTAIL.n306 48.2627
R370 VTAIL.n205 VTAIL.n204 48.2627
R371 VTAIL.n1 VTAIL.n0 48.2625
R372 VTAIL.n103 VTAIL.n102 48.2625
R373 VTAIL.n407 VTAIL.n406 34.1247
R374 VTAIL.n51 VTAIL.n50 34.1247
R375 VTAIL.n101 VTAIL.n100 34.1247
R376 VTAIL.n153 VTAIL.n152 34.1247
R377 VTAIL.n357 VTAIL.n356 34.1247
R378 VTAIL.n305 VTAIL.n304 34.1247
R379 VTAIL.n255 VTAIL.n254 34.1247
R380 VTAIL.n203 VTAIL.n202 34.1247
R381 VTAIL.n407 VTAIL.n357 23.8841
R382 VTAIL.n203 VTAIL.n153 23.8841
R383 VTAIL.n395 VTAIL.n362 13.1884
R384 VTAIL.n39 VTAIL.n6 13.1884
R385 VTAIL.n89 VTAIL.n56 13.1884
R386 VTAIL.n141 VTAIL.n108 13.1884
R387 VTAIL.n314 VTAIL.n312 13.1884
R388 VTAIL.n262 VTAIL.n260 13.1884
R389 VTAIL.n212 VTAIL.n210 13.1884
R390 VTAIL.n160 VTAIL.n158 13.1884
R391 VTAIL.n396 VTAIL.n364 12.8005
R392 VTAIL.n400 VTAIL.n399 12.8005
R393 VTAIL.n40 VTAIL.n8 12.8005
R394 VTAIL.n44 VTAIL.n43 12.8005
R395 VTAIL.n90 VTAIL.n58 12.8005
R396 VTAIL.n94 VTAIL.n93 12.8005
R397 VTAIL.n142 VTAIL.n110 12.8005
R398 VTAIL.n146 VTAIL.n145 12.8005
R399 VTAIL.n350 VTAIL.n349 12.8005
R400 VTAIL.n346 VTAIL.n345 12.8005
R401 VTAIL.n298 VTAIL.n297 12.8005
R402 VTAIL.n294 VTAIL.n293 12.8005
R403 VTAIL.n248 VTAIL.n247 12.8005
R404 VTAIL.n244 VTAIL.n243 12.8005
R405 VTAIL.n196 VTAIL.n195 12.8005
R406 VTAIL.n192 VTAIL.n191 12.8005
R407 VTAIL.n391 VTAIL.n390 12.0247
R408 VTAIL.n403 VTAIL.n360 12.0247
R409 VTAIL.n35 VTAIL.n34 12.0247
R410 VTAIL.n47 VTAIL.n4 12.0247
R411 VTAIL.n85 VTAIL.n84 12.0247
R412 VTAIL.n97 VTAIL.n54 12.0247
R413 VTAIL.n137 VTAIL.n136 12.0247
R414 VTAIL.n149 VTAIL.n106 12.0247
R415 VTAIL.n353 VTAIL.n310 12.0247
R416 VTAIL.n342 VTAIL.n315 12.0247
R417 VTAIL.n301 VTAIL.n258 12.0247
R418 VTAIL.n290 VTAIL.n263 12.0247
R419 VTAIL.n251 VTAIL.n208 12.0247
R420 VTAIL.n240 VTAIL.n213 12.0247
R421 VTAIL.n199 VTAIL.n156 12.0247
R422 VTAIL.n188 VTAIL.n161 12.0247
R423 VTAIL.n389 VTAIL.n366 11.249
R424 VTAIL.n404 VTAIL.n358 11.249
R425 VTAIL.n33 VTAIL.n10 11.249
R426 VTAIL.n48 VTAIL.n2 11.249
R427 VTAIL.n83 VTAIL.n60 11.249
R428 VTAIL.n98 VTAIL.n52 11.249
R429 VTAIL.n135 VTAIL.n112 11.249
R430 VTAIL.n150 VTAIL.n104 11.249
R431 VTAIL.n354 VTAIL.n308 11.249
R432 VTAIL.n341 VTAIL.n318 11.249
R433 VTAIL.n302 VTAIL.n256 11.249
R434 VTAIL.n289 VTAIL.n266 11.249
R435 VTAIL.n252 VTAIL.n206 11.249
R436 VTAIL.n239 VTAIL.n216 11.249
R437 VTAIL.n200 VTAIL.n154 11.249
R438 VTAIL.n187 VTAIL.n164 11.249
R439 VTAIL.n386 VTAIL.n385 10.4732
R440 VTAIL.n30 VTAIL.n29 10.4732
R441 VTAIL.n80 VTAIL.n79 10.4732
R442 VTAIL.n132 VTAIL.n131 10.4732
R443 VTAIL.n338 VTAIL.n337 10.4732
R444 VTAIL.n286 VTAIL.n285 10.4732
R445 VTAIL.n236 VTAIL.n235 10.4732
R446 VTAIL.n184 VTAIL.n183 10.4732
R447 VTAIL.n374 VTAIL.n373 10.2747
R448 VTAIL.n18 VTAIL.n17 10.2747
R449 VTAIL.n68 VTAIL.n67 10.2747
R450 VTAIL.n120 VTAIL.n119 10.2747
R451 VTAIL.n326 VTAIL.n325 10.2747
R452 VTAIL.n274 VTAIL.n273 10.2747
R453 VTAIL.n224 VTAIL.n223 10.2747
R454 VTAIL.n172 VTAIL.n171 10.2747
R455 VTAIL.n382 VTAIL.n368 9.69747
R456 VTAIL.n26 VTAIL.n12 9.69747
R457 VTAIL.n76 VTAIL.n62 9.69747
R458 VTAIL.n128 VTAIL.n114 9.69747
R459 VTAIL.n334 VTAIL.n320 9.69747
R460 VTAIL.n282 VTAIL.n268 9.69747
R461 VTAIL.n232 VTAIL.n218 9.69747
R462 VTAIL.n180 VTAIL.n166 9.69747
R463 VTAIL.n406 VTAIL.n405 9.45567
R464 VTAIL.n50 VTAIL.n49 9.45567
R465 VTAIL.n100 VTAIL.n99 9.45567
R466 VTAIL.n152 VTAIL.n151 9.45567
R467 VTAIL.n356 VTAIL.n355 9.45567
R468 VTAIL.n304 VTAIL.n303 9.45567
R469 VTAIL.n254 VTAIL.n253 9.45567
R470 VTAIL.n202 VTAIL.n201 9.45567
R471 VTAIL.n405 VTAIL.n404 9.3005
R472 VTAIL.n360 VTAIL.n359 9.3005
R473 VTAIL.n399 VTAIL.n398 9.3005
R474 VTAIL.n372 VTAIL.n371 9.3005
R475 VTAIL.n379 VTAIL.n378 9.3005
R476 VTAIL.n381 VTAIL.n380 9.3005
R477 VTAIL.n368 VTAIL.n367 9.3005
R478 VTAIL.n387 VTAIL.n386 9.3005
R479 VTAIL.n389 VTAIL.n388 9.3005
R480 VTAIL.n390 VTAIL.n363 9.3005
R481 VTAIL.n397 VTAIL.n396 9.3005
R482 VTAIL.n49 VTAIL.n48 9.3005
R483 VTAIL.n4 VTAIL.n3 9.3005
R484 VTAIL.n43 VTAIL.n42 9.3005
R485 VTAIL.n16 VTAIL.n15 9.3005
R486 VTAIL.n23 VTAIL.n22 9.3005
R487 VTAIL.n25 VTAIL.n24 9.3005
R488 VTAIL.n12 VTAIL.n11 9.3005
R489 VTAIL.n31 VTAIL.n30 9.3005
R490 VTAIL.n33 VTAIL.n32 9.3005
R491 VTAIL.n34 VTAIL.n7 9.3005
R492 VTAIL.n41 VTAIL.n40 9.3005
R493 VTAIL.n99 VTAIL.n98 9.3005
R494 VTAIL.n54 VTAIL.n53 9.3005
R495 VTAIL.n93 VTAIL.n92 9.3005
R496 VTAIL.n66 VTAIL.n65 9.3005
R497 VTAIL.n73 VTAIL.n72 9.3005
R498 VTAIL.n75 VTAIL.n74 9.3005
R499 VTAIL.n62 VTAIL.n61 9.3005
R500 VTAIL.n81 VTAIL.n80 9.3005
R501 VTAIL.n83 VTAIL.n82 9.3005
R502 VTAIL.n84 VTAIL.n57 9.3005
R503 VTAIL.n91 VTAIL.n90 9.3005
R504 VTAIL.n151 VTAIL.n150 9.3005
R505 VTAIL.n106 VTAIL.n105 9.3005
R506 VTAIL.n145 VTAIL.n144 9.3005
R507 VTAIL.n118 VTAIL.n117 9.3005
R508 VTAIL.n125 VTAIL.n124 9.3005
R509 VTAIL.n127 VTAIL.n126 9.3005
R510 VTAIL.n114 VTAIL.n113 9.3005
R511 VTAIL.n133 VTAIL.n132 9.3005
R512 VTAIL.n135 VTAIL.n134 9.3005
R513 VTAIL.n136 VTAIL.n109 9.3005
R514 VTAIL.n143 VTAIL.n142 9.3005
R515 VTAIL.n324 VTAIL.n323 9.3005
R516 VTAIL.n331 VTAIL.n330 9.3005
R517 VTAIL.n333 VTAIL.n332 9.3005
R518 VTAIL.n320 VTAIL.n319 9.3005
R519 VTAIL.n339 VTAIL.n338 9.3005
R520 VTAIL.n341 VTAIL.n340 9.3005
R521 VTAIL.n315 VTAIL.n313 9.3005
R522 VTAIL.n347 VTAIL.n346 9.3005
R523 VTAIL.n355 VTAIL.n354 9.3005
R524 VTAIL.n310 VTAIL.n309 9.3005
R525 VTAIL.n349 VTAIL.n348 9.3005
R526 VTAIL.n272 VTAIL.n271 9.3005
R527 VTAIL.n279 VTAIL.n278 9.3005
R528 VTAIL.n281 VTAIL.n280 9.3005
R529 VTAIL.n268 VTAIL.n267 9.3005
R530 VTAIL.n287 VTAIL.n286 9.3005
R531 VTAIL.n289 VTAIL.n288 9.3005
R532 VTAIL.n263 VTAIL.n261 9.3005
R533 VTAIL.n295 VTAIL.n294 9.3005
R534 VTAIL.n303 VTAIL.n302 9.3005
R535 VTAIL.n258 VTAIL.n257 9.3005
R536 VTAIL.n297 VTAIL.n296 9.3005
R537 VTAIL.n222 VTAIL.n221 9.3005
R538 VTAIL.n229 VTAIL.n228 9.3005
R539 VTAIL.n231 VTAIL.n230 9.3005
R540 VTAIL.n218 VTAIL.n217 9.3005
R541 VTAIL.n237 VTAIL.n236 9.3005
R542 VTAIL.n239 VTAIL.n238 9.3005
R543 VTAIL.n213 VTAIL.n211 9.3005
R544 VTAIL.n245 VTAIL.n244 9.3005
R545 VTAIL.n253 VTAIL.n252 9.3005
R546 VTAIL.n208 VTAIL.n207 9.3005
R547 VTAIL.n247 VTAIL.n246 9.3005
R548 VTAIL.n170 VTAIL.n169 9.3005
R549 VTAIL.n177 VTAIL.n176 9.3005
R550 VTAIL.n179 VTAIL.n178 9.3005
R551 VTAIL.n166 VTAIL.n165 9.3005
R552 VTAIL.n185 VTAIL.n184 9.3005
R553 VTAIL.n187 VTAIL.n186 9.3005
R554 VTAIL.n161 VTAIL.n159 9.3005
R555 VTAIL.n193 VTAIL.n192 9.3005
R556 VTAIL.n201 VTAIL.n200 9.3005
R557 VTAIL.n156 VTAIL.n155 9.3005
R558 VTAIL.n195 VTAIL.n194 9.3005
R559 VTAIL.n381 VTAIL.n370 8.92171
R560 VTAIL.n25 VTAIL.n14 8.92171
R561 VTAIL.n75 VTAIL.n64 8.92171
R562 VTAIL.n127 VTAIL.n116 8.92171
R563 VTAIL.n333 VTAIL.n322 8.92171
R564 VTAIL.n281 VTAIL.n270 8.92171
R565 VTAIL.n231 VTAIL.n220 8.92171
R566 VTAIL.n179 VTAIL.n168 8.92171
R567 VTAIL.n378 VTAIL.n377 8.14595
R568 VTAIL.n22 VTAIL.n21 8.14595
R569 VTAIL.n72 VTAIL.n71 8.14595
R570 VTAIL.n124 VTAIL.n123 8.14595
R571 VTAIL.n330 VTAIL.n329 8.14595
R572 VTAIL.n278 VTAIL.n277 8.14595
R573 VTAIL.n228 VTAIL.n227 8.14595
R574 VTAIL.n176 VTAIL.n175 8.14595
R575 VTAIL.n374 VTAIL.n372 7.3702
R576 VTAIL.n18 VTAIL.n16 7.3702
R577 VTAIL.n68 VTAIL.n66 7.3702
R578 VTAIL.n120 VTAIL.n118 7.3702
R579 VTAIL.n326 VTAIL.n324 7.3702
R580 VTAIL.n274 VTAIL.n272 7.3702
R581 VTAIL.n224 VTAIL.n222 7.3702
R582 VTAIL.n172 VTAIL.n170 7.3702
R583 VTAIL.n377 VTAIL.n372 5.81868
R584 VTAIL.n21 VTAIL.n16 5.81868
R585 VTAIL.n71 VTAIL.n66 5.81868
R586 VTAIL.n123 VTAIL.n118 5.81868
R587 VTAIL.n329 VTAIL.n324 5.81868
R588 VTAIL.n277 VTAIL.n272 5.81868
R589 VTAIL.n227 VTAIL.n222 5.81868
R590 VTAIL.n175 VTAIL.n170 5.81868
R591 VTAIL.n378 VTAIL.n370 5.04292
R592 VTAIL.n22 VTAIL.n14 5.04292
R593 VTAIL.n72 VTAIL.n64 5.04292
R594 VTAIL.n124 VTAIL.n116 5.04292
R595 VTAIL.n330 VTAIL.n322 5.04292
R596 VTAIL.n278 VTAIL.n270 5.04292
R597 VTAIL.n228 VTAIL.n220 5.04292
R598 VTAIL.n176 VTAIL.n168 5.04292
R599 VTAIL.n382 VTAIL.n381 4.26717
R600 VTAIL.n26 VTAIL.n25 4.26717
R601 VTAIL.n76 VTAIL.n75 4.26717
R602 VTAIL.n128 VTAIL.n127 4.26717
R603 VTAIL.n334 VTAIL.n333 4.26717
R604 VTAIL.n282 VTAIL.n281 4.26717
R605 VTAIL.n232 VTAIL.n231 4.26717
R606 VTAIL.n180 VTAIL.n179 4.26717
R607 VTAIL.n385 VTAIL.n368 3.49141
R608 VTAIL.n29 VTAIL.n12 3.49141
R609 VTAIL.n79 VTAIL.n62 3.49141
R610 VTAIL.n131 VTAIL.n114 3.49141
R611 VTAIL.n337 VTAIL.n320 3.49141
R612 VTAIL.n285 VTAIL.n268 3.49141
R613 VTAIL.n235 VTAIL.n218 3.49141
R614 VTAIL.n183 VTAIL.n166 3.49141
R615 VTAIL.n205 VTAIL.n203 3.46602
R616 VTAIL.n255 VTAIL.n205 3.46602
R617 VTAIL.n307 VTAIL.n305 3.46602
R618 VTAIL.n357 VTAIL.n307 3.46602
R619 VTAIL.n153 VTAIL.n103 3.46602
R620 VTAIL.n103 VTAIL.n101 3.46602
R621 VTAIL.n51 VTAIL.n1 3.46602
R622 VTAIL VTAIL.n407 3.40783
R623 VTAIL.n373 VTAIL.n371 2.84303
R624 VTAIL.n17 VTAIL.n15 2.84303
R625 VTAIL.n67 VTAIL.n65 2.84303
R626 VTAIL.n119 VTAIL.n117 2.84303
R627 VTAIL.n325 VTAIL.n323 2.84303
R628 VTAIL.n273 VTAIL.n271 2.84303
R629 VTAIL.n223 VTAIL.n221 2.84303
R630 VTAIL.n171 VTAIL.n169 2.84303
R631 VTAIL.n386 VTAIL.n366 2.71565
R632 VTAIL.n406 VTAIL.n358 2.71565
R633 VTAIL.n30 VTAIL.n10 2.71565
R634 VTAIL.n50 VTAIL.n2 2.71565
R635 VTAIL.n80 VTAIL.n60 2.71565
R636 VTAIL.n100 VTAIL.n52 2.71565
R637 VTAIL.n132 VTAIL.n112 2.71565
R638 VTAIL.n152 VTAIL.n104 2.71565
R639 VTAIL.n356 VTAIL.n308 2.71565
R640 VTAIL.n338 VTAIL.n318 2.71565
R641 VTAIL.n304 VTAIL.n256 2.71565
R642 VTAIL.n286 VTAIL.n266 2.71565
R643 VTAIL.n254 VTAIL.n206 2.71565
R644 VTAIL.n236 VTAIL.n216 2.71565
R645 VTAIL.n202 VTAIL.n154 2.71565
R646 VTAIL.n184 VTAIL.n164 2.71565
R647 VTAIL.n0 VTAIL.t6 2.12041
R648 VTAIL.n0 VTAIL.t7 2.12041
R649 VTAIL.n102 VTAIL.t11 2.12041
R650 VTAIL.n102 VTAIL.t8 2.12041
R651 VTAIL.n306 VTAIL.t14 2.12041
R652 VTAIL.n306 VTAIL.t12 2.12041
R653 VTAIL.n204 VTAIL.t0 2.12041
R654 VTAIL.n204 VTAIL.t3 2.12041
R655 VTAIL.n391 VTAIL.n389 1.93989
R656 VTAIL.n404 VTAIL.n403 1.93989
R657 VTAIL.n35 VTAIL.n33 1.93989
R658 VTAIL.n48 VTAIL.n47 1.93989
R659 VTAIL.n85 VTAIL.n83 1.93989
R660 VTAIL.n98 VTAIL.n97 1.93989
R661 VTAIL.n137 VTAIL.n135 1.93989
R662 VTAIL.n150 VTAIL.n149 1.93989
R663 VTAIL.n354 VTAIL.n353 1.93989
R664 VTAIL.n342 VTAIL.n341 1.93989
R665 VTAIL.n302 VTAIL.n301 1.93989
R666 VTAIL.n290 VTAIL.n289 1.93989
R667 VTAIL.n252 VTAIL.n251 1.93989
R668 VTAIL.n240 VTAIL.n239 1.93989
R669 VTAIL.n200 VTAIL.n199 1.93989
R670 VTAIL.n188 VTAIL.n187 1.93989
R671 VTAIL.n390 VTAIL.n364 1.16414
R672 VTAIL.n400 VTAIL.n360 1.16414
R673 VTAIL.n34 VTAIL.n8 1.16414
R674 VTAIL.n44 VTAIL.n4 1.16414
R675 VTAIL.n84 VTAIL.n58 1.16414
R676 VTAIL.n94 VTAIL.n54 1.16414
R677 VTAIL.n136 VTAIL.n110 1.16414
R678 VTAIL.n146 VTAIL.n106 1.16414
R679 VTAIL.n350 VTAIL.n310 1.16414
R680 VTAIL.n345 VTAIL.n315 1.16414
R681 VTAIL.n298 VTAIL.n258 1.16414
R682 VTAIL.n293 VTAIL.n263 1.16414
R683 VTAIL.n248 VTAIL.n208 1.16414
R684 VTAIL.n243 VTAIL.n213 1.16414
R685 VTAIL.n196 VTAIL.n156 1.16414
R686 VTAIL.n191 VTAIL.n161 1.16414
R687 VTAIL.n305 VTAIL.n255 0.470328
R688 VTAIL.n101 VTAIL.n51 0.470328
R689 VTAIL.n396 VTAIL.n395 0.388379
R690 VTAIL.n399 VTAIL.n362 0.388379
R691 VTAIL.n40 VTAIL.n39 0.388379
R692 VTAIL.n43 VTAIL.n6 0.388379
R693 VTAIL.n90 VTAIL.n89 0.388379
R694 VTAIL.n93 VTAIL.n56 0.388379
R695 VTAIL.n142 VTAIL.n141 0.388379
R696 VTAIL.n145 VTAIL.n108 0.388379
R697 VTAIL.n349 VTAIL.n312 0.388379
R698 VTAIL.n346 VTAIL.n314 0.388379
R699 VTAIL.n297 VTAIL.n260 0.388379
R700 VTAIL.n294 VTAIL.n262 0.388379
R701 VTAIL.n247 VTAIL.n210 0.388379
R702 VTAIL.n244 VTAIL.n212 0.388379
R703 VTAIL.n195 VTAIL.n158 0.388379
R704 VTAIL.n192 VTAIL.n160 0.388379
R705 VTAIL.n379 VTAIL.n371 0.155672
R706 VTAIL.n380 VTAIL.n379 0.155672
R707 VTAIL.n380 VTAIL.n367 0.155672
R708 VTAIL.n387 VTAIL.n367 0.155672
R709 VTAIL.n388 VTAIL.n387 0.155672
R710 VTAIL.n388 VTAIL.n363 0.155672
R711 VTAIL.n397 VTAIL.n363 0.155672
R712 VTAIL.n398 VTAIL.n397 0.155672
R713 VTAIL.n398 VTAIL.n359 0.155672
R714 VTAIL.n405 VTAIL.n359 0.155672
R715 VTAIL.n23 VTAIL.n15 0.155672
R716 VTAIL.n24 VTAIL.n23 0.155672
R717 VTAIL.n24 VTAIL.n11 0.155672
R718 VTAIL.n31 VTAIL.n11 0.155672
R719 VTAIL.n32 VTAIL.n31 0.155672
R720 VTAIL.n32 VTAIL.n7 0.155672
R721 VTAIL.n41 VTAIL.n7 0.155672
R722 VTAIL.n42 VTAIL.n41 0.155672
R723 VTAIL.n42 VTAIL.n3 0.155672
R724 VTAIL.n49 VTAIL.n3 0.155672
R725 VTAIL.n73 VTAIL.n65 0.155672
R726 VTAIL.n74 VTAIL.n73 0.155672
R727 VTAIL.n74 VTAIL.n61 0.155672
R728 VTAIL.n81 VTAIL.n61 0.155672
R729 VTAIL.n82 VTAIL.n81 0.155672
R730 VTAIL.n82 VTAIL.n57 0.155672
R731 VTAIL.n91 VTAIL.n57 0.155672
R732 VTAIL.n92 VTAIL.n91 0.155672
R733 VTAIL.n92 VTAIL.n53 0.155672
R734 VTAIL.n99 VTAIL.n53 0.155672
R735 VTAIL.n125 VTAIL.n117 0.155672
R736 VTAIL.n126 VTAIL.n125 0.155672
R737 VTAIL.n126 VTAIL.n113 0.155672
R738 VTAIL.n133 VTAIL.n113 0.155672
R739 VTAIL.n134 VTAIL.n133 0.155672
R740 VTAIL.n134 VTAIL.n109 0.155672
R741 VTAIL.n143 VTAIL.n109 0.155672
R742 VTAIL.n144 VTAIL.n143 0.155672
R743 VTAIL.n144 VTAIL.n105 0.155672
R744 VTAIL.n151 VTAIL.n105 0.155672
R745 VTAIL.n355 VTAIL.n309 0.155672
R746 VTAIL.n348 VTAIL.n309 0.155672
R747 VTAIL.n348 VTAIL.n347 0.155672
R748 VTAIL.n347 VTAIL.n313 0.155672
R749 VTAIL.n340 VTAIL.n313 0.155672
R750 VTAIL.n340 VTAIL.n339 0.155672
R751 VTAIL.n339 VTAIL.n319 0.155672
R752 VTAIL.n332 VTAIL.n319 0.155672
R753 VTAIL.n332 VTAIL.n331 0.155672
R754 VTAIL.n331 VTAIL.n323 0.155672
R755 VTAIL.n303 VTAIL.n257 0.155672
R756 VTAIL.n296 VTAIL.n257 0.155672
R757 VTAIL.n296 VTAIL.n295 0.155672
R758 VTAIL.n295 VTAIL.n261 0.155672
R759 VTAIL.n288 VTAIL.n261 0.155672
R760 VTAIL.n288 VTAIL.n287 0.155672
R761 VTAIL.n287 VTAIL.n267 0.155672
R762 VTAIL.n280 VTAIL.n267 0.155672
R763 VTAIL.n280 VTAIL.n279 0.155672
R764 VTAIL.n279 VTAIL.n271 0.155672
R765 VTAIL.n253 VTAIL.n207 0.155672
R766 VTAIL.n246 VTAIL.n207 0.155672
R767 VTAIL.n246 VTAIL.n245 0.155672
R768 VTAIL.n245 VTAIL.n211 0.155672
R769 VTAIL.n238 VTAIL.n211 0.155672
R770 VTAIL.n238 VTAIL.n237 0.155672
R771 VTAIL.n237 VTAIL.n217 0.155672
R772 VTAIL.n230 VTAIL.n217 0.155672
R773 VTAIL.n230 VTAIL.n229 0.155672
R774 VTAIL.n229 VTAIL.n221 0.155672
R775 VTAIL.n201 VTAIL.n155 0.155672
R776 VTAIL.n194 VTAIL.n155 0.155672
R777 VTAIL.n194 VTAIL.n193 0.155672
R778 VTAIL.n193 VTAIL.n159 0.155672
R779 VTAIL.n186 VTAIL.n159 0.155672
R780 VTAIL.n186 VTAIL.n185 0.155672
R781 VTAIL.n185 VTAIL.n165 0.155672
R782 VTAIL.n178 VTAIL.n165 0.155672
R783 VTAIL.n178 VTAIL.n177 0.155672
R784 VTAIL.n177 VTAIL.n169 0.155672
R785 VTAIL VTAIL.n1 0.0586897
R786 B.n932 B.n931 585
R787 B.n933 B.n932 585
R788 B.n315 B.n161 585
R789 B.n314 B.n313 585
R790 B.n312 B.n311 585
R791 B.n310 B.n309 585
R792 B.n308 B.n307 585
R793 B.n306 B.n305 585
R794 B.n304 B.n303 585
R795 B.n302 B.n301 585
R796 B.n300 B.n299 585
R797 B.n298 B.n297 585
R798 B.n296 B.n295 585
R799 B.n294 B.n293 585
R800 B.n292 B.n291 585
R801 B.n290 B.n289 585
R802 B.n288 B.n287 585
R803 B.n286 B.n285 585
R804 B.n284 B.n283 585
R805 B.n282 B.n281 585
R806 B.n280 B.n279 585
R807 B.n278 B.n277 585
R808 B.n276 B.n275 585
R809 B.n274 B.n273 585
R810 B.n272 B.n271 585
R811 B.n270 B.n269 585
R812 B.n268 B.n267 585
R813 B.n266 B.n265 585
R814 B.n264 B.n263 585
R815 B.n262 B.n261 585
R816 B.n260 B.n259 585
R817 B.n258 B.n257 585
R818 B.n256 B.n255 585
R819 B.n254 B.n253 585
R820 B.n252 B.n251 585
R821 B.n249 B.n248 585
R822 B.n247 B.n246 585
R823 B.n245 B.n244 585
R824 B.n243 B.n242 585
R825 B.n241 B.n240 585
R826 B.n239 B.n238 585
R827 B.n237 B.n236 585
R828 B.n235 B.n234 585
R829 B.n233 B.n232 585
R830 B.n231 B.n230 585
R831 B.n229 B.n228 585
R832 B.n227 B.n226 585
R833 B.n225 B.n224 585
R834 B.n223 B.n222 585
R835 B.n221 B.n220 585
R836 B.n219 B.n218 585
R837 B.n217 B.n216 585
R838 B.n215 B.n214 585
R839 B.n213 B.n212 585
R840 B.n211 B.n210 585
R841 B.n209 B.n208 585
R842 B.n207 B.n206 585
R843 B.n205 B.n204 585
R844 B.n203 B.n202 585
R845 B.n201 B.n200 585
R846 B.n199 B.n198 585
R847 B.n197 B.n196 585
R848 B.n195 B.n194 585
R849 B.n193 B.n192 585
R850 B.n191 B.n190 585
R851 B.n189 B.n188 585
R852 B.n187 B.n186 585
R853 B.n185 B.n184 585
R854 B.n183 B.n182 585
R855 B.n181 B.n180 585
R856 B.n179 B.n178 585
R857 B.n177 B.n176 585
R858 B.n175 B.n174 585
R859 B.n173 B.n172 585
R860 B.n171 B.n170 585
R861 B.n169 B.n168 585
R862 B.n123 B.n122 585
R863 B.n936 B.n935 585
R864 B.n930 B.n162 585
R865 B.n162 B.n120 585
R866 B.n929 B.n119 585
R867 B.n940 B.n119 585
R868 B.n928 B.n118 585
R869 B.n941 B.n118 585
R870 B.n927 B.n117 585
R871 B.n942 B.n117 585
R872 B.n926 B.n925 585
R873 B.n925 B.n113 585
R874 B.n924 B.n112 585
R875 B.n948 B.n112 585
R876 B.n923 B.n111 585
R877 B.n949 B.n111 585
R878 B.n922 B.n110 585
R879 B.n950 B.n110 585
R880 B.n921 B.n920 585
R881 B.n920 B.n109 585
R882 B.n919 B.n105 585
R883 B.n956 B.n105 585
R884 B.n918 B.n104 585
R885 B.n957 B.n104 585
R886 B.n917 B.n103 585
R887 B.n958 B.n103 585
R888 B.n916 B.n915 585
R889 B.n915 B.n99 585
R890 B.n914 B.n98 585
R891 B.n964 B.n98 585
R892 B.n913 B.n97 585
R893 B.n965 B.n97 585
R894 B.n912 B.n96 585
R895 B.n966 B.n96 585
R896 B.n911 B.n910 585
R897 B.n910 B.n92 585
R898 B.n909 B.n91 585
R899 B.n972 B.n91 585
R900 B.n908 B.n90 585
R901 B.n973 B.n90 585
R902 B.n907 B.n89 585
R903 B.n974 B.n89 585
R904 B.n906 B.n905 585
R905 B.n905 B.n85 585
R906 B.n904 B.n84 585
R907 B.n980 B.n84 585
R908 B.n903 B.n83 585
R909 B.n981 B.n83 585
R910 B.n902 B.n82 585
R911 B.n982 B.n82 585
R912 B.n901 B.n900 585
R913 B.n900 B.n81 585
R914 B.n899 B.n77 585
R915 B.n988 B.n77 585
R916 B.n898 B.n76 585
R917 B.n989 B.n76 585
R918 B.n897 B.n75 585
R919 B.n990 B.n75 585
R920 B.n896 B.n895 585
R921 B.n895 B.n71 585
R922 B.n894 B.n70 585
R923 B.n996 B.n70 585
R924 B.n893 B.n69 585
R925 B.n997 B.n69 585
R926 B.n892 B.n68 585
R927 B.n998 B.n68 585
R928 B.n891 B.n890 585
R929 B.n890 B.n64 585
R930 B.n889 B.n63 585
R931 B.n1004 B.n63 585
R932 B.n888 B.n62 585
R933 B.n1005 B.n62 585
R934 B.n887 B.n61 585
R935 B.n1006 B.n61 585
R936 B.n886 B.n885 585
R937 B.n885 B.n57 585
R938 B.n884 B.n56 585
R939 B.n1012 B.n56 585
R940 B.n883 B.n55 585
R941 B.n1013 B.n55 585
R942 B.n882 B.n54 585
R943 B.n1014 B.n54 585
R944 B.n881 B.n880 585
R945 B.n880 B.n50 585
R946 B.n879 B.n49 585
R947 B.n1020 B.n49 585
R948 B.n878 B.n48 585
R949 B.n1021 B.n48 585
R950 B.n877 B.n47 585
R951 B.n1022 B.n47 585
R952 B.n876 B.n875 585
R953 B.n875 B.n43 585
R954 B.n874 B.n42 585
R955 B.n1028 B.n42 585
R956 B.n873 B.n41 585
R957 B.n1029 B.n41 585
R958 B.n872 B.n40 585
R959 B.n1030 B.n40 585
R960 B.n871 B.n870 585
R961 B.n870 B.n36 585
R962 B.n869 B.n35 585
R963 B.n1036 B.n35 585
R964 B.n868 B.n34 585
R965 B.n1037 B.n34 585
R966 B.n867 B.n33 585
R967 B.n1038 B.n33 585
R968 B.n866 B.n865 585
R969 B.n865 B.n29 585
R970 B.n864 B.n28 585
R971 B.n1044 B.n28 585
R972 B.n863 B.n27 585
R973 B.n1045 B.n27 585
R974 B.n862 B.n26 585
R975 B.n1046 B.n26 585
R976 B.n861 B.n860 585
R977 B.n860 B.n22 585
R978 B.n859 B.n21 585
R979 B.n1052 B.n21 585
R980 B.n858 B.n20 585
R981 B.n1053 B.n20 585
R982 B.n857 B.n19 585
R983 B.n1054 B.n19 585
R984 B.n856 B.n855 585
R985 B.n855 B.n15 585
R986 B.n854 B.n14 585
R987 B.n1060 B.n14 585
R988 B.n853 B.n13 585
R989 B.n1061 B.n13 585
R990 B.n852 B.n12 585
R991 B.n1062 B.n12 585
R992 B.n851 B.n850 585
R993 B.n850 B.n8 585
R994 B.n849 B.n7 585
R995 B.n1068 B.n7 585
R996 B.n848 B.n6 585
R997 B.n1069 B.n6 585
R998 B.n847 B.n5 585
R999 B.n1070 B.n5 585
R1000 B.n846 B.n845 585
R1001 B.n845 B.n4 585
R1002 B.n844 B.n316 585
R1003 B.n844 B.n843 585
R1004 B.n834 B.n317 585
R1005 B.n318 B.n317 585
R1006 B.n836 B.n835 585
R1007 B.n837 B.n836 585
R1008 B.n833 B.n323 585
R1009 B.n323 B.n322 585
R1010 B.n832 B.n831 585
R1011 B.n831 B.n830 585
R1012 B.n325 B.n324 585
R1013 B.n326 B.n325 585
R1014 B.n823 B.n822 585
R1015 B.n824 B.n823 585
R1016 B.n821 B.n331 585
R1017 B.n331 B.n330 585
R1018 B.n820 B.n819 585
R1019 B.n819 B.n818 585
R1020 B.n333 B.n332 585
R1021 B.n334 B.n333 585
R1022 B.n811 B.n810 585
R1023 B.n812 B.n811 585
R1024 B.n809 B.n339 585
R1025 B.n339 B.n338 585
R1026 B.n808 B.n807 585
R1027 B.n807 B.n806 585
R1028 B.n341 B.n340 585
R1029 B.n342 B.n341 585
R1030 B.n799 B.n798 585
R1031 B.n800 B.n799 585
R1032 B.n797 B.n347 585
R1033 B.n347 B.n346 585
R1034 B.n796 B.n795 585
R1035 B.n795 B.n794 585
R1036 B.n349 B.n348 585
R1037 B.n350 B.n349 585
R1038 B.n787 B.n786 585
R1039 B.n788 B.n787 585
R1040 B.n785 B.n355 585
R1041 B.n355 B.n354 585
R1042 B.n784 B.n783 585
R1043 B.n783 B.n782 585
R1044 B.n357 B.n356 585
R1045 B.n358 B.n357 585
R1046 B.n775 B.n774 585
R1047 B.n776 B.n775 585
R1048 B.n773 B.n363 585
R1049 B.n363 B.n362 585
R1050 B.n772 B.n771 585
R1051 B.n771 B.n770 585
R1052 B.n365 B.n364 585
R1053 B.n366 B.n365 585
R1054 B.n763 B.n762 585
R1055 B.n764 B.n763 585
R1056 B.n761 B.n371 585
R1057 B.n371 B.n370 585
R1058 B.n760 B.n759 585
R1059 B.n759 B.n758 585
R1060 B.n373 B.n372 585
R1061 B.n374 B.n373 585
R1062 B.n751 B.n750 585
R1063 B.n752 B.n751 585
R1064 B.n749 B.n379 585
R1065 B.n379 B.n378 585
R1066 B.n748 B.n747 585
R1067 B.n747 B.n746 585
R1068 B.n381 B.n380 585
R1069 B.n382 B.n381 585
R1070 B.n739 B.n738 585
R1071 B.n740 B.n739 585
R1072 B.n737 B.n387 585
R1073 B.n387 B.n386 585
R1074 B.n736 B.n735 585
R1075 B.n735 B.n734 585
R1076 B.n389 B.n388 585
R1077 B.n390 B.n389 585
R1078 B.n727 B.n726 585
R1079 B.n728 B.n727 585
R1080 B.n725 B.n395 585
R1081 B.n395 B.n394 585
R1082 B.n724 B.n723 585
R1083 B.n723 B.n722 585
R1084 B.n397 B.n396 585
R1085 B.n715 B.n397 585
R1086 B.n714 B.n713 585
R1087 B.n716 B.n714 585
R1088 B.n712 B.n402 585
R1089 B.n402 B.n401 585
R1090 B.n711 B.n710 585
R1091 B.n710 B.n709 585
R1092 B.n404 B.n403 585
R1093 B.n405 B.n404 585
R1094 B.n702 B.n701 585
R1095 B.n703 B.n702 585
R1096 B.n700 B.n410 585
R1097 B.n410 B.n409 585
R1098 B.n699 B.n698 585
R1099 B.n698 B.n697 585
R1100 B.n412 B.n411 585
R1101 B.n413 B.n412 585
R1102 B.n690 B.n689 585
R1103 B.n691 B.n690 585
R1104 B.n688 B.n418 585
R1105 B.n418 B.n417 585
R1106 B.n687 B.n686 585
R1107 B.n686 B.n685 585
R1108 B.n420 B.n419 585
R1109 B.n421 B.n420 585
R1110 B.n678 B.n677 585
R1111 B.n679 B.n678 585
R1112 B.n676 B.n426 585
R1113 B.n426 B.n425 585
R1114 B.n675 B.n674 585
R1115 B.n674 B.n673 585
R1116 B.n428 B.n427 585
R1117 B.n666 B.n428 585
R1118 B.n665 B.n664 585
R1119 B.n667 B.n665 585
R1120 B.n663 B.n433 585
R1121 B.n433 B.n432 585
R1122 B.n662 B.n661 585
R1123 B.n661 B.n660 585
R1124 B.n435 B.n434 585
R1125 B.n436 B.n435 585
R1126 B.n653 B.n652 585
R1127 B.n654 B.n653 585
R1128 B.n651 B.n441 585
R1129 B.n441 B.n440 585
R1130 B.n650 B.n649 585
R1131 B.n649 B.n648 585
R1132 B.n443 B.n442 585
R1133 B.n444 B.n443 585
R1134 B.n644 B.n643 585
R1135 B.n447 B.n446 585
R1136 B.n640 B.n639 585
R1137 B.n641 B.n640 585
R1138 B.n638 B.n485 585
R1139 B.n637 B.n636 585
R1140 B.n635 B.n634 585
R1141 B.n633 B.n632 585
R1142 B.n631 B.n630 585
R1143 B.n629 B.n628 585
R1144 B.n627 B.n626 585
R1145 B.n625 B.n624 585
R1146 B.n623 B.n622 585
R1147 B.n621 B.n620 585
R1148 B.n619 B.n618 585
R1149 B.n617 B.n616 585
R1150 B.n615 B.n614 585
R1151 B.n613 B.n612 585
R1152 B.n611 B.n610 585
R1153 B.n609 B.n608 585
R1154 B.n607 B.n606 585
R1155 B.n605 B.n604 585
R1156 B.n603 B.n602 585
R1157 B.n601 B.n600 585
R1158 B.n599 B.n598 585
R1159 B.n597 B.n596 585
R1160 B.n595 B.n594 585
R1161 B.n593 B.n592 585
R1162 B.n591 B.n590 585
R1163 B.n589 B.n588 585
R1164 B.n587 B.n586 585
R1165 B.n585 B.n584 585
R1166 B.n583 B.n582 585
R1167 B.n581 B.n580 585
R1168 B.n579 B.n578 585
R1169 B.n576 B.n575 585
R1170 B.n574 B.n573 585
R1171 B.n572 B.n571 585
R1172 B.n570 B.n569 585
R1173 B.n568 B.n567 585
R1174 B.n566 B.n565 585
R1175 B.n564 B.n563 585
R1176 B.n562 B.n561 585
R1177 B.n560 B.n559 585
R1178 B.n558 B.n557 585
R1179 B.n556 B.n555 585
R1180 B.n554 B.n553 585
R1181 B.n552 B.n551 585
R1182 B.n550 B.n549 585
R1183 B.n548 B.n547 585
R1184 B.n546 B.n545 585
R1185 B.n544 B.n543 585
R1186 B.n542 B.n541 585
R1187 B.n540 B.n539 585
R1188 B.n538 B.n537 585
R1189 B.n536 B.n535 585
R1190 B.n534 B.n533 585
R1191 B.n532 B.n531 585
R1192 B.n530 B.n529 585
R1193 B.n528 B.n527 585
R1194 B.n526 B.n525 585
R1195 B.n524 B.n523 585
R1196 B.n522 B.n521 585
R1197 B.n520 B.n519 585
R1198 B.n518 B.n517 585
R1199 B.n516 B.n515 585
R1200 B.n514 B.n513 585
R1201 B.n512 B.n511 585
R1202 B.n510 B.n509 585
R1203 B.n508 B.n507 585
R1204 B.n506 B.n505 585
R1205 B.n504 B.n503 585
R1206 B.n502 B.n501 585
R1207 B.n500 B.n499 585
R1208 B.n498 B.n497 585
R1209 B.n496 B.n495 585
R1210 B.n494 B.n493 585
R1211 B.n492 B.n491 585
R1212 B.n645 B.n445 585
R1213 B.n445 B.n444 585
R1214 B.n647 B.n646 585
R1215 B.n648 B.n647 585
R1216 B.n439 B.n438 585
R1217 B.n440 B.n439 585
R1218 B.n656 B.n655 585
R1219 B.n655 B.n654 585
R1220 B.n657 B.n437 585
R1221 B.n437 B.n436 585
R1222 B.n659 B.n658 585
R1223 B.n660 B.n659 585
R1224 B.n431 B.n430 585
R1225 B.n432 B.n431 585
R1226 B.n669 B.n668 585
R1227 B.n668 B.n667 585
R1228 B.n670 B.n429 585
R1229 B.n666 B.n429 585
R1230 B.n672 B.n671 585
R1231 B.n673 B.n672 585
R1232 B.n424 B.n423 585
R1233 B.n425 B.n424 585
R1234 B.n681 B.n680 585
R1235 B.n680 B.n679 585
R1236 B.n682 B.n422 585
R1237 B.n422 B.n421 585
R1238 B.n684 B.n683 585
R1239 B.n685 B.n684 585
R1240 B.n416 B.n415 585
R1241 B.n417 B.n416 585
R1242 B.n693 B.n692 585
R1243 B.n692 B.n691 585
R1244 B.n694 B.n414 585
R1245 B.n414 B.n413 585
R1246 B.n696 B.n695 585
R1247 B.n697 B.n696 585
R1248 B.n408 B.n407 585
R1249 B.n409 B.n408 585
R1250 B.n705 B.n704 585
R1251 B.n704 B.n703 585
R1252 B.n706 B.n406 585
R1253 B.n406 B.n405 585
R1254 B.n708 B.n707 585
R1255 B.n709 B.n708 585
R1256 B.n400 B.n399 585
R1257 B.n401 B.n400 585
R1258 B.n718 B.n717 585
R1259 B.n717 B.n716 585
R1260 B.n719 B.n398 585
R1261 B.n715 B.n398 585
R1262 B.n721 B.n720 585
R1263 B.n722 B.n721 585
R1264 B.n393 B.n392 585
R1265 B.n394 B.n393 585
R1266 B.n730 B.n729 585
R1267 B.n729 B.n728 585
R1268 B.n731 B.n391 585
R1269 B.n391 B.n390 585
R1270 B.n733 B.n732 585
R1271 B.n734 B.n733 585
R1272 B.n385 B.n384 585
R1273 B.n386 B.n385 585
R1274 B.n742 B.n741 585
R1275 B.n741 B.n740 585
R1276 B.n743 B.n383 585
R1277 B.n383 B.n382 585
R1278 B.n745 B.n744 585
R1279 B.n746 B.n745 585
R1280 B.n377 B.n376 585
R1281 B.n378 B.n377 585
R1282 B.n754 B.n753 585
R1283 B.n753 B.n752 585
R1284 B.n755 B.n375 585
R1285 B.n375 B.n374 585
R1286 B.n757 B.n756 585
R1287 B.n758 B.n757 585
R1288 B.n369 B.n368 585
R1289 B.n370 B.n369 585
R1290 B.n766 B.n765 585
R1291 B.n765 B.n764 585
R1292 B.n767 B.n367 585
R1293 B.n367 B.n366 585
R1294 B.n769 B.n768 585
R1295 B.n770 B.n769 585
R1296 B.n361 B.n360 585
R1297 B.n362 B.n361 585
R1298 B.n778 B.n777 585
R1299 B.n777 B.n776 585
R1300 B.n779 B.n359 585
R1301 B.n359 B.n358 585
R1302 B.n781 B.n780 585
R1303 B.n782 B.n781 585
R1304 B.n353 B.n352 585
R1305 B.n354 B.n353 585
R1306 B.n790 B.n789 585
R1307 B.n789 B.n788 585
R1308 B.n791 B.n351 585
R1309 B.n351 B.n350 585
R1310 B.n793 B.n792 585
R1311 B.n794 B.n793 585
R1312 B.n345 B.n344 585
R1313 B.n346 B.n345 585
R1314 B.n802 B.n801 585
R1315 B.n801 B.n800 585
R1316 B.n803 B.n343 585
R1317 B.n343 B.n342 585
R1318 B.n805 B.n804 585
R1319 B.n806 B.n805 585
R1320 B.n337 B.n336 585
R1321 B.n338 B.n337 585
R1322 B.n814 B.n813 585
R1323 B.n813 B.n812 585
R1324 B.n815 B.n335 585
R1325 B.n335 B.n334 585
R1326 B.n817 B.n816 585
R1327 B.n818 B.n817 585
R1328 B.n329 B.n328 585
R1329 B.n330 B.n329 585
R1330 B.n826 B.n825 585
R1331 B.n825 B.n824 585
R1332 B.n827 B.n327 585
R1333 B.n327 B.n326 585
R1334 B.n829 B.n828 585
R1335 B.n830 B.n829 585
R1336 B.n321 B.n320 585
R1337 B.n322 B.n321 585
R1338 B.n839 B.n838 585
R1339 B.n838 B.n837 585
R1340 B.n840 B.n319 585
R1341 B.n319 B.n318 585
R1342 B.n842 B.n841 585
R1343 B.n843 B.n842 585
R1344 B.n2 B.n0 585
R1345 B.n4 B.n2 585
R1346 B.n3 B.n1 585
R1347 B.n1069 B.n3 585
R1348 B.n1067 B.n1066 585
R1349 B.n1068 B.n1067 585
R1350 B.n1065 B.n9 585
R1351 B.n9 B.n8 585
R1352 B.n1064 B.n1063 585
R1353 B.n1063 B.n1062 585
R1354 B.n11 B.n10 585
R1355 B.n1061 B.n11 585
R1356 B.n1059 B.n1058 585
R1357 B.n1060 B.n1059 585
R1358 B.n1057 B.n16 585
R1359 B.n16 B.n15 585
R1360 B.n1056 B.n1055 585
R1361 B.n1055 B.n1054 585
R1362 B.n18 B.n17 585
R1363 B.n1053 B.n18 585
R1364 B.n1051 B.n1050 585
R1365 B.n1052 B.n1051 585
R1366 B.n1049 B.n23 585
R1367 B.n23 B.n22 585
R1368 B.n1048 B.n1047 585
R1369 B.n1047 B.n1046 585
R1370 B.n25 B.n24 585
R1371 B.n1045 B.n25 585
R1372 B.n1043 B.n1042 585
R1373 B.n1044 B.n1043 585
R1374 B.n1041 B.n30 585
R1375 B.n30 B.n29 585
R1376 B.n1040 B.n1039 585
R1377 B.n1039 B.n1038 585
R1378 B.n32 B.n31 585
R1379 B.n1037 B.n32 585
R1380 B.n1035 B.n1034 585
R1381 B.n1036 B.n1035 585
R1382 B.n1033 B.n37 585
R1383 B.n37 B.n36 585
R1384 B.n1032 B.n1031 585
R1385 B.n1031 B.n1030 585
R1386 B.n39 B.n38 585
R1387 B.n1029 B.n39 585
R1388 B.n1027 B.n1026 585
R1389 B.n1028 B.n1027 585
R1390 B.n1025 B.n44 585
R1391 B.n44 B.n43 585
R1392 B.n1024 B.n1023 585
R1393 B.n1023 B.n1022 585
R1394 B.n46 B.n45 585
R1395 B.n1021 B.n46 585
R1396 B.n1019 B.n1018 585
R1397 B.n1020 B.n1019 585
R1398 B.n1017 B.n51 585
R1399 B.n51 B.n50 585
R1400 B.n1016 B.n1015 585
R1401 B.n1015 B.n1014 585
R1402 B.n53 B.n52 585
R1403 B.n1013 B.n53 585
R1404 B.n1011 B.n1010 585
R1405 B.n1012 B.n1011 585
R1406 B.n1009 B.n58 585
R1407 B.n58 B.n57 585
R1408 B.n1008 B.n1007 585
R1409 B.n1007 B.n1006 585
R1410 B.n60 B.n59 585
R1411 B.n1005 B.n60 585
R1412 B.n1003 B.n1002 585
R1413 B.n1004 B.n1003 585
R1414 B.n1001 B.n65 585
R1415 B.n65 B.n64 585
R1416 B.n1000 B.n999 585
R1417 B.n999 B.n998 585
R1418 B.n67 B.n66 585
R1419 B.n997 B.n67 585
R1420 B.n995 B.n994 585
R1421 B.n996 B.n995 585
R1422 B.n993 B.n72 585
R1423 B.n72 B.n71 585
R1424 B.n992 B.n991 585
R1425 B.n991 B.n990 585
R1426 B.n74 B.n73 585
R1427 B.n989 B.n74 585
R1428 B.n987 B.n986 585
R1429 B.n988 B.n987 585
R1430 B.n985 B.n78 585
R1431 B.n81 B.n78 585
R1432 B.n984 B.n983 585
R1433 B.n983 B.n982 585
R1434 B.n80 B.n79 585
R1435 B.n981 B.n80 585
R1436 B.n979 B.n978 585
R1437 B.n980 B.n979 585
R1438 B.n977 B.n86 585
R1439 B.n86 B.n85 585
R1440 B.n976 B.n975 585
R1441 B.n975 B.n974 585
R1442 B.n88 B.n87 585
R1443 B.n973 B.n88 585
R1444 B.n971 B.n970 585
R1445 B.n972 B.n971 585
R1446 B.n969 B.n93 585
R1447 B.n93 B.n92 585
R1448 B.n968 B.n967 585
R1449 B.n967 B.n966 585
R1450 B.n95 B.n94 585
R1451 B.n965 B.n95 585
R1452 B.n963 B.n962 585
R1453 B.n964 B.n963 585
R1454 B.n961 B.n100 585
R1455 B.n100 B.n99 585
R1456 B.n960 B.n959 585
R1457 B.n959 B.n958 585
R1458 B.n102 B.n101 585
R1459 B.n957 B.n102 585
R1460 B.n955 B.n954 585
R1461 B.n956 B.n955 585
R1462 B.n953 B.n106 585
R1463 B.n109 B.n106 585
R1464 B.n952 B.n951 585
R1465 B.n951 B.n950 585
R1466 B.n108 B.n107 585
R1467 B.n949 B.n108 585
R1468 B.n947 B.n946 585
R1469 B.n948 B.n947 585
R1470 B.n945 B.n114 585
R1471 B.n114 B.n113 585
R1472 B.n944 B.n943 585
R1473 B.n943 B.n942 585
R1474 B.n116 B.n115 585
R1475 B.n941 B.n116 585
R1476 B.n939 B.n938 585
R1477 B.n940 B.n939 585
R1478 B.n937 B.n121 585
R1479 B.n121 B.n120 585
R1480 B.n1072 B.n1071 585
R1481 B.n1071 B.n1070 585
R1482 B.n643 B.n445 550.159
R1483 B.n935 B.n121 550.159
R1484 B.n491 B.n443 550.159
R1485 B.n932 B.n162 550.159
R1486 B.n488 B.t21 314.286
R1487 B.n163 B.t14 314.286
R1488 B.n486 B.t11 314.286
R1489 B.n165 B.t17 314.286
R1490 B.n488 B.t19 270.257
R1491 B.n486 B.t8 270.257
R1492 B.n165 B.t16 270.257
R1493 B.n163 B.t12 270.257
R1494 B.n933 B.n160 256.663
R1495 B.n933 B.n159 256.663
R1496 B.n933 B.n158 256.663
R1497 B.n933 B.n157 256.663
R1498 B.n933 B.n156 256.663
R1499 B.n933 B.n155 256.663
R1500 B.n933 B.n154 256.663
R1501 B.n933 B.n153 256.663
R1502 B.n933 B.n152 256.663
R1503 B.n933 B.n151 256.663
R1504 B.n933 B.n150 256.663
R1505 B.n933 B.n149 256.663
R1506 B.n933 B.n148 256.663
R1507 B.n933 B.n147 256.663
R1508 B.n933 B.n146 256.663
R1509 B.n933 B.n145 256.663
R1510 B.n933 B.n144 256.663
R1511 B.n933 B.n143 256.663
R1512 B.n933 B.n142 256.663
R1513 B.n933 B.n141 256.663
R1514 B.n933 B.n140 256.663
R1515 B.n933 B.n139 256.663
R1516 B.n933 B.n138 256.663
R1517 B.n933 B.n137 256.663
R1518 B.n933 B.n136 256.663
R1519 B.n933 B.n135 256.663
R1520 B.n933 B.n134 256.663
R1521 B.n933 B.n133 256.663
R1522 B.n933 B.n132 256.663
R1523 B.n933 B.n131 256.663
R1524 B.n933 B.n130 256.663
R1525 B.n933 B.n129 256.663
R1526 B.n933 B.n128 256.663
R1527 B.n933 B.n127 256.663
R1528 B.n933 B.n126 256.663
R1529 B.n933 B.n125 256.663
R1530 B.n933 B.n124 256.663
R1531 B.n934 B.n933 256.663
R1532 B.n642 B.n641 256.663
R1533 B.n641 B.n448 256.663
R1534 B.n641 B.n449 256.663
R1535 B.n641 B.n450 256.663
R1536 B.n641 B.n451 256.663
R1537 B.n641 B.n452 256.663
R1538 B.n641 B.n453 256.663
R1539 B.n641 B.n454 256.663
R1540 B.n641 B.n455 256.663
R1541 B.n641 B.n456 256.663
R1542 B.n641 B.n457 256.663
R1543 B.n641 B.n458 256.663
R1544 B.n641 B.n459 256.663
R1545 B.n641 B.n460 256.663
R1546 B.n641 B.n461 256.663
R1547 B.n641 B.n462 256.663
R1548 B.n641 B.n463 256.663
R1549 B.n641 B.n464 256.663
R1550 B.n641 B.n465 256.663
R1551 B.n641 B.n466 256.663
R1552 B.n641 B.n467 256.663
R1553 B.n641 B.n468 256.663
R1554 B.n641 B.n469 256.663
R1555 B.n641 B.n470 256.663
R1556 B.n641 B.n471 256.663
R1557 B.n641 B.n472 256.663
R1558 B.n641 B.n473 256.663
R1559 B.n641 B.n474 256.663
R1560 B.n641 B.n475 256.663
R1561 B.n641 B.n476 256.663
R1562 B.n641 B.n477 256.663
R1563 B.n641 B.n478 256.663
R1564 B.n641 B.n479 256.663
R1565 B.n641 B.n480 256.663
R1566 B.n641 B.n481 256.663
R1567 B.n641 B.n482 256.663
R1568 B.n641 B.n483 256.663
R1569 B.n641 B.n484 256.663
R1570 B.n489 B.t20 236.323
R1571 B.n164 B.t15 236.323
R1572 B.n487 B.t10 236.323
R1573 B.n166 B.t18 236.323
R1574 B.n647 B.n445 163.367
R1575 B.n647 B.n439 163.367
R1576 B.n655 B.n439 163.367
R1577 B.n655 B.n437 163.367
R1578 B.n659 B.n437 163.367
R1579 B.n659 B.n431 163.367
R1580 B.n668 B.n431 163.367
R1581 B.n668 B.n429 163.367
R1582 B.n672 B.n429 163.367
R1583 B.n672 B.n424 163.367
R1584 B.n680 B.n424 163.367
R1585 B.n680 B.n422 163.367
R1586 B.n684 B.n422 163.367
R1587 B.n684 B.n416 163.367
R1588 B.n692 B.n416 163.367
R1589 B.n692 B.n414 163.367
R1590 B.n696 B.n414 163.367
R1591 B.n696 B.n408 163.367
R1592 B.n704 B.n408 163.367
R1593 B.n704 B.n406 163.367
R1594 B.n708 B.n406 163.367
R1595 B.n708 B.n400 163.367
R1596 B.n717 B.n400 163.367
R1597 B.n717 B.n398 163.367
R1598 B.n721 B.n398 163.367
R1599 B.n721 B.n393 163.367
R1600 B.n729 B.n393 163.367
R1601 B.n729 B.n391 163.367
R1602 B.n733 B.n391 163.367
R1603 B.n733 B.n385 163.367
R1604 B.n741 B.n385 163.367
R1605 B.n741 B.n383 163.367
R1606 B.n745 B.n383 163.367
R1607 B.n745 B.n377 163.367
R1608 B.n753 B.n377 163.367
R1609 B.n753 B.n375 163.367
R1610 B.n757 B.n375 163.367
R1611 B.n757 B.n369 163.367
R1612 B.n765 B.n369 163.367
R1613 B.n765 B.n367 163.367
R1614 B.n769 B.n367 163.367
R1615 B.n769 B.n361 163.367
R1616 B.n777 B.n361 163.367
R1617 B.n777 B.n359 163.367
R1618 B.n781 B.n359 163.367
R1619 B.n781 B.n353 163.367
R1620 B.n789 B.n353 163.367
R1621 B.n789 B.n351 163.367
R1622 B.n793 B.n351 163.367
R1623 B.n793 B.n345 163.367
R1624 B.n801 B.n345 163.367
R1625 B.n801 B.n343 163.367
R1626 B.n805 B.n343 163.367
R1627 B.n805 B.n337 163.367
R1628 B.n813 B.n337 163.367
R1629 B.n813 B.n335 163.367
R1630 B.n817 B.n335 163.367
R1631 B.n817 B.n329 163.367
R1632 B.n825 B.n329 163.367
R1633 B.n825 B.n327 163.367
R1634 B.n829 B.n327 163.367
R1635 B.n829 B.n321 163.367
R1636 B.n838 B.n321 163.367
R1637 B.n838 B.n319 163.367
R1638 B.n842 B.n319 163.367
R1639 B.n842 B.n2 163.367
R1640 B.n1071 B.n2 163.367
R1641 B.n1071 B.n3 163.367
R1642 B.n1067 B.n3 163.367
R1643 B.n1067 B.n9 163.367
R1644 B.n1063 B.n9 163.367
R1645 B.n1063 B.n11 163.367
R1646 B.n1059 B.n11 163.367
R1647 B.n1059 B.n16 163.367
R1648 B.n1055 B.n16 163.367
R1649 B.n1055 B.n18 163.367
R1650 B.n1051 B.n18 163.367
R1651 B.n1051 B.n23 163.367
R1652 B.n1047 B.n23 163.367
R1653 B.n1047 B.n25 163.367
R1654 B.n1043 B.n25 163.367
R1655 B.n1043 B.n30 163.367
R1656 B.n1039 B.n30 163.367
R1657 B.n1039 B.n32 163.367
R1658 B.n1035 B.n32 163.367
R1659 B.n1035 B.n37 163.367
R1660 B.n1031 B.n37 163.367
R1661 B.n1031 B.n39 163.367
R1662 B.n1027 B.n39 163.367
R1663 B.n1027 B.n44 163.367
R1664 B.n1023 B.n44 163.367
R1665 B.n1023 B.n46 163.367
R1666 B.n1019 B.n46 163.367
R1667 B.n1019 B.n51 163.367
R1668 B.n1015 B.n51 163.367
R1669 B.n1015 B.n53 163.367
R1670 B.n1011 B.n53 163.367
R1671 B.n1011 B.n58 163.367
R1672 B.n1007 B.n58 163.367
R1673 B.n1007 B.n60 163.367
R1674 B.n1003 B.n60 163.367
R1675 B.n1003 B.n65 163.367
R1676 B.n999 B.n65 163.367
R1677 B.n999 B.n67 163.367
R1678 B.n995 B.n67 163.367
R1679 B.n995 B.n72 163.367
R1680 B.n991 B.n72 163.367
R1681 B.n991 B.n74 163.367
R1682 B.n987 B.n74 163.367
R1683 B.n987 B.n78 163.367
R1684 B.n983 B.n78 163.367
R1685 B.n983 B.n80 163.367
R1686 B.n979 B.n80 163.367
R1687 B.n979 B.n86 163.367
R1688 B.n975 B.n86 163.367
R1689 B.n975 B.n88 163.367
R1690 B.n971 B.n88 163.367
R1691 B.n971 B.n93 163.367
R1692 B.n967 B.n93 163.367
R1693 B.n967 B.n95 163.367
R1694 B.n963 B.n95 163.367
R1695 B.n963 B.n100 163.367
R1696 B.n959 B.n100 163.367
R1697 B.n959 B.n102 163.367
R1698 B.n955 B.n102 163.367
R1699 B.n955 B.n106 163.367
R1700 B.n951 B.n106 163.367
R1701 B.n951 B.n108 163.367
R1702 B.n947 B.n108 163.367
R1703 B.n947 B.n114 163.367
R1704 B.n943 B.n114 163.367
R1705 B.n943 B.n116 163.367
R1706 B.n939 B.n116 163.367
R1707 B.n939 B.n121 163.367
R1708 B.n640 B.n447 163.367
R1709 B.n640 B.n485 163.367
R1710 B.n636 B.n635 163.367
R1711 B.n632 B.n631 163.367
R1712 B.n628 B.n627 163.367
R1713 B.n624 B.n623 163.367
R1714 B.n620 B.n619 163.367
R1715 B.n616 B.n615 163.367
R1716 B.n612 B.n611 163.367
R1717 B.n608 B.n607 163.367
R1718 B.n604 B.n603 163.367
R1719 B.n600 B.n599 163.367
R1720 B.n596 B.n595 163.367
R1721 B.n592 B.n591 163.367
R1722 B.n588 B.n587 163.367
R1723 B.n584 B.n583 163.367
R1724 B.n580 B.n579 163.367
R1725 B.n575 B.n574 163.367
R1726 B.n571 B.n570 163.367
R1727 B.n567 B.n566 163.367
R1728 B.n563 B.n562 163.367
R1729 B.n559 B.n558 163.367
R1730 B.n555 B.n554 163.367
R1731 B.n551 B.n550 163.367
R1732 B.n547 B.n546 163.367
R1733 B.n543 B.n542 163.367
R1734 B.n539 B.n538 163.367
R1735 B.n535 B.n534 163.367
R1736 B.n531 B.n530 163.367
R1737 B.n527 B.n526 163.367
R1738 B.n523 B.n522 163.367
R1739 B.n519 B.n518 163.367
R1740 B.n515 B.n514 163.367
R1741 B.n511 B.n510 163.367
R1742 B.n507 B.n506 163.367
R1743 B.n503 B.n502 163.367
R1744 B.n499 B.n498 163.367
R1745 B.n495 B.n494 163.367
R1746 B.n649 B.n443 163.367
R1747 B.n649 B.n441 163.367
R1748 B.n653 B.n441 163.367
R1749 B.n653 B.n435 163.367
R1750 B.n661 B.n435 163.367
R1751 B.n661 B.n433 163.367
R1752 B.n665 B.n433 163.367
R1753 B.n665 B.n428 163.367
R1754 B.n674 B.n428 163.367
R1755 B.n674 B.n426 163.367
R1756 B.n678 B.n426 163.367
R1757 B.n678 B.n420 163.367
R1758 B.n686 B.n420 163.367
R1759 B.n686 B.n418 163.367
R1760 B.n690 B.n418 163.367
R1761 B.n690 B.n412 163.367
R1762 B.n698 B.n412 163.367
R1763 B.n698 B.n410 163.367
R1764 B.n702 B.n410 163.367
R1765 B.n702 B.n404 163.367
R1766 B.n710 B.n404 163.367
R1767 B.n710 B.n402 163.367
R1768 B.n714 B.n402 163.367
R1769 B.n714 B.n397 163.367
R1770 B.n723 B.n397 163.367
R1771 B.n723 B.n395 163.367
R1772 B.n727 B.n395 163.367
R1773 B.n727 B.n389 163.367
R1774 B.n735 B.n389 163.367
R1775 B.n735 B.n387 163.367
R1776 B.n739 B.n387 163.367
R1777 B.n739 B.n381 163.367
R1778 B.n747 B.n381 163.367
R1779 B.n747 B.n379 163.367
R1780 B.n751 B.n379 163.367
R1781 B.n751 B.n373 163.367
R1782 B.n759 B.n373 163.367
R1783 B.n759 B.n371 163.367
R1784 B.n763 B.n371 163.367
R1785 B.n763 B.n365 163.367
R1786 B.n771 B.n365 163.367
R1787 B.n771 B.n363 163.367
R1788 B.n775 B.n363 163.367
R1789 B.n775 B.n357 163.367
R1790 B.n783 B.n357 163.367
R1791 B.n783 B.n355 163.367
R1792 B.n787 B.n355 163.367
R1793 B.n787 B.n349 163.367
R1794 B.n795 B.n349 163.367
R1795 B.n795 B.n347 163.367
R1796 B.n799 B.n347 163.367
R1797 B.n799 B.n341 163.367
R1798 B.n807 B.n341 163.367
R1799 B.n807 B.n339 163.367
R1800 B.n811 B.n339 163.367
R1801 B.n811 B.n333 163.367
R1802 B.n819 B.n333 163.367
R1803 B.n819 B.n331 163.367
R1804 B.n823 B.n331 163.367
R1805 B.n823 B.n325 163.367
R1806 B.n831 B.n325 163.367
R1807 B.n831 B.n323 163.367
R1808 B.n836 B.n323 163.367
R1809 B.n836 B.n317 163.367
R1810 B.n844 B.n317 163.367
R1811 B.n845 B.n844 163.367
R1812 B.n845 B.n5 163.367
R1813 B.n6 B.n5 163.367
R1814 B.n7 B.n6 163.367
R1815 B.n850 B.n7 163.367
R1816 B.n850 B.n12 163.367
R1817 B.n13 B.n12 163.367
R1818 B.n14 B.n13 163.367
R1819 B.n855 B.n14 163.367
R1820 B.n855 B.n19 163.367
R1821 B.n20 B.n19 163.367
R1822 B.n21 B.n20 163.367
R1823 B.n860 B.n21 163.367
R1824 B.n860 B.n26 163.367
R1825 B.n27 B.n26 163.367
R1826 B.n28 B.n27 163.367
R1827 B.n865 B.n28 163.367
R1828 B.n865 B.n33 163.367
R1829 B.n34 B.n33 163.367
R1830 B.n35 B.n34 163.367
R1831 B.n870 B.n35 163.367
R1832 B.n870 B.n40 163.367
R1833 B.n41 B.n40 163.367
R1834 B.n42 B.n41 163.367
R1835 B.n875 B.n42 163.367
R1836 B.n875 B.n47 163.367
R1837 B.n48 B.n47 163.367
R1838 B.n49 B.n48 163.367
R1839 B.n880 B.n49 163.367
R1840 B.n880 B.n54 163.367
R1841 B.n55 B.n54 163.367
R1842 B.n56 B.n55 163.367
R1843 B.n885 B.n56 163.367
R1844 B.n885 B.n61 163.367
R1845 B.n62 B.n61 163.367
R1846 B.n63 B.n62 163.367
R1847 B.n890 B.n63 163.367
R1848 B.n890 B.n68 163.367
R1849 B.n69 B.n68 163.367
R1850 B.n70 B.n69 163.367
R1851 B.n895 B.n70 163.367
R1852 B.n895 B.n75 163.367
R1853 B.n76 B.n75 163.367
R1854 B.n77 B.n76 163.367
R1855 B.n900 B.n77 163.367
R1856 B.n900 B.n82 163.367
R1857 B.n83 B.n82 163.367
R1858 B.n84 B.n83 163.367
R1859 B.n905 B.n84 163.367
R1860 B.n905 B.n89 163.367
R1861 B.n90 B.n89 163.367
R1862 B.n91 B.n90 163.367
R1863 B.n910 B.n91 163.367
R1864 B.n910 B.n96 163.367
R1865 B.n97 B.n96 163.367
R1866 B.n98 B.n97 163.367
R1867 B.n915 B.n98 163.367
R1868 B.n915 B.n103 163.367
R1869 B.n104 B.n103 163.367
R1870 B.n105 B.n104 163.367
R1871 B.n920 B.n105 163.367
R1872 B.n920 B.n110 163.367
R1873 B.n111 B.n110 163.367
R1874 B.n112 B.n111 163.367
R1875 B.n925 B.n112 163.367
R1876 B.n925 B.n117 163.367
R1877 B.n118 B.n117 163.367
R1878 B.n119 B.n118 163.367
R1879 B.n162 B.n119 163.367
R1880 B.n168 B.n123 163.367
R1881 B.n172 B.n171 163.367
R1882 B.n176 B.n175 163.367
R1883 B.n180 B.n179 163.367
R1884 B.n184 B.n183 163.367
R1885 B.n188 B.n187 163.367
R1886 B.n192 B.n191 163.367
R1887 B.n196 B.n195 163.367
R1888 B.n200 B.n199 163.367
R1889 B.n204 B.n203 163.367
R1890 B.n208 B.n207 163.367
R1891 B.n212 B.n211 163.367
R1892 B.n216 B.n215 163.367
R1893 B.n220 B.n219 163.367
R1894 B.n224 B.n223 163.367
R1895 B.n228 B.n227 163.367
R1896 B.n232 B.n231 163.367
R1897 B.n236 B.n235 163.367
R1898 B.n240 B.n239 163.367
R1899 B.n244 B.n243 163.367
R1900 B.n248 B.n247 163.367
R1901 B.n253 B.n252 163.367
R1902 B.n257 B.n256 163.367
R1903 B.n261 B.n260 163.367
R1904 B.n265 B.n264 163.367
R1905 B.n269 B.n268 163.367
R1906 B.n273 B.n272 163.367
R1907 B.n277 B.n276 163.367
R1908 B.n281 B.n280 163.367
R1909 B.n285 B.n284 163.367
R1910 B.n289 B.n288 163.367
R1911 B.n293 B.n292 163.367
R1912 B.n297 B.n296 163.367
R1913 B.n301 B.n300 163.367
R1914 B.n305 B.n304 163.367
R1915 B.n309 B.n308 163.367
R1916 B.n313 B.n312 163.367
R1917 B.n932 B.n161 163.367
R1918 B.n641 B.n444 104.62
R1919 B.n933 B.n120 104.62
R1920 B.n489 B.n488 77.9641
R1921 B.n487 B.n486 77.9641
R1922 B.n166 B.n165 77.9641
R1923 B.n164 B.n163 77.9641
R1924 B.n643 B.n642 71.676
R1925 B.n485 B.n448 71.676
R1926 B.n635 B.n449 71.676
R1927 B.n631 B.n450 71.676
R1928 B.n627 B.n451 71.676
R1929 B.n623 B.n452 71.676
R1930 B.n619 B.n453 71.676
R1931 B.n615 B.n454 71.676
R1932 B.n611 B.n455 71.676
R1933 B.n607 B.n456 71.676
R1934 B.n603 B.n457 71.676
R1935 B.n599 B.n458 71.676
R1936 B.n595 B.n459 71.676
R1937 B.n591 B.n460 71.676
R1938 B.n587 B.n461 71.676
R1939 B.n583 B.n462 71.676
R1940 B.n579 B.n463 71.676
R1941 B.n574 B.n464 71.676
R1942 B.n570 B.n465 71.676
R1943 B.n566 B.n466 71.676
R1944 B.n562 B.n467 71.676
R1945 B.n558 B.n468 71.676
R1946 B.n554 B.n469 71.676
R1947 B.n550 B.n470 71.676
R1948 B.n546 B.n471 71.676
R1949 B.n542 B.n472 71.676
R1950 B.n538 B.n473 71.676
R1951 B.n534 B.n474 71.676
R1952 B.n530 B.n475 71.676
R1953 B.n526 B.n476 71.676
R1954 B.n522 B.n477 71.676
R1955 B.n518 B.n478 71.676
R1956 B.n514 B.n479 71.676
R1957 B.n510 B.n480 71.676
R1958 B.n506 B.n481 71.676
R1959 B.n502 B.n482 71.676
R1960 B.n498 B.n483 71.676
R1961 B.n494 B.n484 71.676
R1962 B.n935 B.n934 71.676
R1963 B.n168 B.n124 71.676
R1964 B.n172 B.n125 71.676
R1965 B.n176 B.n126 71.676
R1966 B.n180 B.n127 71.676
R1967 B.n184 B.n128 71.676
R1968 B.n188 B.n129 71.676
R1969 B.n192 B.n130 71.676
R1970 B.n196 B.n131 71.676
R1971 B.n200 B.n132 71.676
R1972 B.n204 B.n133 71.676
R1973 B.n208 B.n134 71.676
R1974 B.n212 B.n135 71.676
R1975 B.n216 B.n136 71.676
R1976 B.n220 B.n137 71.676
R1977 B.n224 B.n138 71.676
R1978 B.n228 B.n139 71.676
R1979 B.n232 B.n140 71.676
R1980 B.n236 B.n141 71.676
R1981 B.n240 B.n142 71.676
R1982 B.n244 B.n143 71.676
R1983 B.n248 B.n144 71.676
R1984 B.n253 B.n145 71.676
R1985 B.n257 B.n146 71.676
R1986 B.n261 B.n147 71.676
R1987 B.n265 B.n148 71.676
R1988 B.n269 B.n149 71.676
R1989 B.n273 B.n150 71.676
R1990 B.n277 B.n151 71.676
R1991 B.n281 B.n152 71.676
R1992 B.n285 B.n153 71.676
R1993 B.n289 B.n154 71.676
R1994 B.n293 B.n155 71.676
R1995 B.n297 B.n156 71.676
R1996 B.n301 B.n157 71.676
R1997 B.n305 B.n158 71.676
R1998 B.n309 B.n159 71.676
R1999 B.n313 B.n160 71.676
R2000 B.n161 B.n160 71.676
R2001 B.n312 B.n159 71.676
R2002 B.n308 B.n158 71.676
R2003 B.n304 B.n157 71.676
R2004 B.n300 B.n156 71.676
R2005 B.n296 B.n155 71.676
R2006 B.n292 B.n154 71.676
R2007 B.n288 B.n153 71.676
R2008 B.n284 B.n152 71.676
R2009 B.n280 B.n151 71.676
R2010 B.n276 B.n150 71.676
R2011 B.n272 B.n149 71.676
R2012 B.n268 B.n148 71.676
R2013 B.n264 B.n147 71.676
R2014 B.n260 B.n146 71.676
R2015 B.n256 B.n145 71.676
R2016 B.n252 B.n144 71.676
R2017 B.n247 B.n143 71.676
R2018 B.n243 B.n142 71.676
R2019 B.n239 B.n141 71.676
R2020 B.n235 B.n140 71.676
R2021 B.n231 B.n139 71.676
R2022 B.n227 B.n138 71.676
R2023 B.n223 B.n137 71.676
R2024 B.n219 B.n136 71.676
R2025 B.n215 B.n135 71.676
R2026 B.n211 B.n134 71.676
R2027 B.n207 B.n133 71.676
R2028 B.n203 B.n132 71.676
R2029 B.n199 B.n131 71.676
R2030 B.n195 B.n130 71.676
R2031 B.n191 B.n129 71.676
R2032 B.n187 B.n128 71.676
R2033 B.n183 B.n127 71.676
R2034 B.n179 B.n126 71.676
R2035 B.n175 B.n125 71.676
R2036 B.n171 B.n124 71.676
R2037 B.n934 B.n123 71.676
R2038 B.n642 B.n447 71.676
R2039 B.n636 B.n448 71.676
R2040 B.n632 B.n449 71.676
R2041 B.n628 B.n450 71.676
R2042 B.n624 B.n451 71.676
R2043 B.n620 B.n452 71.676
R2044 B.n616 B.n453 71.676
R2045 B.n612 B.n454 71.676
R2046 B.n608 B.n455 71.676
R2047 B.n604 B.n456 71.676
R2048 B.n600 B.n457 71.676
R2049 B.n596 B.n458 71.676
R2050 B.n592 B.n459 71.676
R2051 B.n588 B.n460 71.676
R2052 B.n584 B.n461 71.676
R2053 B.n580 B.n462 71.676
R2054 B.n575 B.n463 71.676
R2055 B.n571 B.n464 71.676
R2056 B.n567 B.n465 71.676
R2057 B.n563 B.n466 71.676
R2058 B.n559 B.n467 71.676
R2059 B.n555 B.n468 71.676
R2060 B.n551 B.n469 71.676
R2061 B.n547 B.n470 71.676
R2062 B.n543 B.n471 71.676
R2063 B.n539 B.n472 71.676
R2064 B.n535 B.n473 71.676
R2065 B.n531 B.n474 71.676
R2066 B.n527 B.n475 71.676
R2067 B.n523 B.n476 71.676
R2068 B.n519 B.n477 71.676
R2069 B.n515 B.n478 71.676
R2070 B.n511 B.n479 71.676
R2071 B.n507 B.n480 71.676
R2072 B.n503 B.n481 71.676
R2073 B.n499 B.n482 71.676
R2074 B.n495 B.n483 71.676
R2075 B.n491 B.n484 71.676
R2076 B.n490 B.n489 59.5399
R2077 B.n577 B.n487 59.5399
R2078 B.n167 B.n166 59.5399
R2079 B.n250 B.n164 59.5399
R2080 B.n648 B.n444 51.1808
R2081 B.n648 B.n440 51.1808
R2082 B.n654 B.n440 51.1808
R2083 B.n654 B.n436 51.1808
R2084 B.n660 B.n436 51.1808
R2085 B.n660 B.n432 51.1808
R2086 B.n667 B.n432 51.1808
R2087 B.n667 B.n666 51.1808
R2088 B.n673 B.n425 51.1808
R2089 B.n679 B.n425 51.1808
R2090 B.n679 B.n421 51.1808
R2091 B.n685 B.n421 51.1808
R2092 B.n685 B.n417 51.1808
R2093 B.n691 B.n417 51.1808
R2094 B.n691 B.n413 51.1808
R2095 B.n697 B.n413 51.1808
R2096 B.n697 B.n409 51.1808
R2097 B.n703 B.n409 51.1808
R2098 B.n703 B.n405 51.1808
R2099 B.n709 B.n405 51.1808
R2100 B.n709 B.n401 51.1808
R2101 B.n716 B.n401 51.1808
R2102 B.n716 B.n715 51.1808
R2103 B.n722 B.n394 51.1808
R2104 B.n728 B.n394 51.1808
R2105 B.n728 B.n390 51.1808
R2106 B.n734 B.n390 51.1808
R2107 B.n734 B.n386 51.1808
R2108 B.n740 B.n386 51.1808
R2109 B.n740 B.n382 51.1808
R2110 B.n746 B.n382 51.1808
R2111 B.n746 B.n378 51.1808
R2112 B.n752 B.n378 51.1808
R2113 B.n758 B.n374 51.1808
R2114 B.n758 B.n370 51.1808
R2115 B.n764 B.n370 51.1808
R2116 B.n764 B.n366 51.1808
R2117 B.n770 B.n366 51.1808
R2118 B.n770 B.n362 51.1808
R2119 B.n776 B.n362 51.1808
R2120 B.n776 B.n358 51.1808
R2121 B.n782 B.n358 51.1808
R2122 B.n782 B.n354 51.1808
R2123 B.n788 B.n354 51.1808
R2124 B.n794 B.n350 51.1808
R2125 B.n794 B.n346 51.1808
R2126 B.n800 B.n346 51.1808
R2127 B.n800 B.n342 51.1808
R2128 B.n806 B.n342 51.1808
R2129 B.n806 B.n338 51.1808
R2130 B.n812 B.n338 51.1808
R2131 B.n812 B.n334 51.1808
R2132 B.n818 B.n334 51.1808
R2133 B.n818 B.n330 51.1808
R2134 B.n824 B.n330 51.1808
R2135 B.n830 B.n326 51.1808
R2136 B.n830 B.n322 51.1808
R2137 B.n837 B.n322 51.1808
R2138 B.n837 B.n318 51.1808
R2139 B.n843 B.n318 51.1808
R2140 B.n843 B.n4 51.1808
R2141 B.n1070 B.n4 51.1808
R2142 B.n1070 B.n1069 51.1808
R2143 B.n1069 B.n1068 51.1808
R2144 B.n1068 B.n8 51.1808
R2145 B.n1062 B.n8 51.1808
R2146 B.n1062 B.n1061 51.1808
R2147 B.n1061 B.n1060 51.1808
R2148 B.n1060 B.n15 51.1808
R2149 B.n1054 B.n1053 51.1808
R2150 B.n1053 B.n1052 51.1808
R2151 B.n1052 B.n22 51.1808
R2152 B.n1046 B.n22 51.1808
R2153 B.n1046 B.n1045 51.1808
R2154 B.n1045 B.n1044 51.1808
R2155 B.n1044 B.n29 51.1808
R2156 B.n1038 B.n29 51.1808
R2157 B.n1038 B.n1037 51.1808
R2158 B.n1037 B.n1036 51.1808
R2159 B.n1036 B.n36 51.1808
R2160 B.n1030 B.n1029 51.1808
R2161 B.n1029 B.n1028 51.1808
R2162 B.n1028 B.n43 51.1808
R2163 B.n1022 B.n43 51.1808
R2164 B.n1022 B.n1021 51.1808
R2165 B.n1021 B.n1020 51.1808
R2166 B.n1020 B.n50 51.1808
R2167 B.n1014 B.n50 51.1808
R2168 B.n1014 B.n1013 51.1808
R2169 B.n1013 B.n1012 51.1808
R2170 B.n1012 B.n57 51.1808
R2171 B.n1006 B.n1005 51.1808
R2172 B.n1005 B.n1004 51.1808
R2173 B.n1004 B.n64 51.1808
R2174 B.n998 B.n64 51.1808
R2175 B.n998 B.n997 51.1808
R2176 B.n997 B.n996 51.1808
R2177 B.n996 B.n71 51.1808
R2178 B.n990 B.n71 51.1808
R2179 B.n990 B.n989 51.1808
R2180 B.n989 B.n988 51.1808
R2181 B.n982 B.n81 51.1808
R2182 B.n982 B.n981 51.1808
R2183 B.n981 B.n980 51.1808
R2184 B.n980 B.n85 51.1808
R2185 B.n974 B.n85 51.1808
R2186 B.n974 B.n973 51.1808
R2187 B.n973 B.n972 51.1808
R2188 B.n972 B.n92 51.1808
R2189 B.n966 B.n92 51.1808
R2190 B.n966 B.n965 51.1808
R2191 B.n965 B.n964 51.1808
R2192 B.n964 B.n99 51.1808
R2193 B.n958 B.n99 51.1808
R2194 B.n958 B.n957 51.1808
R2195 B.n957 B.n956 51.1808
R2196 B.n950 B.n109 51.1808
R2197 B.n950 B.n949 51.1808
R2198 B.n949 B.n948 51.1808
R2199 B.n948 B.n113 51.1808
R2200 B.n942 B.n113 51.1808
R2201 B.n942 B.n941 51.1808
R2202 B.n941 B.n940 51.1808
R2203 B.n940 B.n120 51.1808
R2204 B.n666 B.t9 50.4281
R2205 B.n722 B.t5 50.4281
R2206 B.n988 B.t4 50.4281
R2207 B.n109 B.t13 50.4281
R2208 B.n752 B.t0 42.9016
R2209 B.n1006 B.t7 42.9016
R2210 B.n931 B.n930 35.7468
R2211 B.n937 B.n936 35.7468
R2212 B.n492 B.n442 35.7468
R2213 B.n645 B.n644 35.7468
R2214 B.n788 B.t3 33.8698
R2215 B.n1030 B.t6 33.8698
R2216 B.t1 B.n326 26.3433
R2217 B.t2 B.n15 26.3433
R2218 B.n824 B.t1 24.838
R2219 B.n1054 B.t2 24.838
R2220 B B.n1072 18.0485
R2221 B.t3 B.n350 17.3115
R2222 B.t6 B.n36 17.3115
R2223 B.n936 B.n122 10.6151
R2224 B.n169 B.n122 10.6151
R2225 B.n170 B.n169 10.6151
R2226 B.n173 B.n170 10.6151
R2227 B.n174 B.n173 10.6151
R2228 B.n177 B.n174 10.6151
R2229 B.n178 B.n177 10.6151
R2230 B.n181 B.n178 10.6151
R2231 B.n182 B.n181 10.6151
R2232 B.n185 B.n182 10.6151
R2233 B.n186 B.n185 10.6151
R2234 B.n189 B.n186 10.6151
R2235 B.n190 B.n189 10.6151
R2236 B.n193 B.n190 10.6151
R2237 B.n194 B.n193 10.6151
R2238 B.n197 B.n194 10.6151
R2239 B.n198 B.n197 10.6151
R2240 B.n201 B.n198 10.6151
R2241 B.n202 B.n201 10.6151
R2242 B.n205 B.n202 10.6151
R2243 B.n206 B.n205 10.6151
R2244 B.n209 B.n206 10.6151
R2245 B.n210 B.n209 10.6151
R2246 B.n213 B.n210 10.6151
R2247 B.n214 B.n213 10.6151
R2248 B.n217 B.n214 10.6151
R2249 B.n218 B.n217 10.6151
R2250 B.n221 B.n218 10.6151
R2251 B.n222 B.n221 10.6151
R2252 B.n225 B.n222 10.6151
R2253 B.n226 B.n225 10.6151
R2254 B.n229 B.n226 10.6151
R2255 B.n230 B.n229 10.6151
R2256 B.n234 B.n233 10.6151
R2257 B.n237 B.n234 10.6151
R2258 B.n238 B.n237 10.6151
R2259 B.n241 B.n238 10.6151
R2260 B.n242 B.n241 10.6151
R2261 B.n245 B.n242 10.6151
R2262 B.n246 B.n245 10.6151
R2263 B.n249 B.n246 10.6151
R2264 B.n254 B.n251 10.6151
R2265 B.n255 B.n254 10.6151
R2266 B.n258 B.n255 10.6151
R2267 B.n259 B.n258 10.6151
R2268 B.n262 B.n259 10.6151
R2269 B.n263 B.n262 10.6151
R2270 B.n266 B.n263 10.6151
R2271 B.n267 B.n266 10.6151
R2272 B.n270 B.n267 10.6151
R2273 B.n271 B.n270 10.6151
R2274 B.n274 B.n271 10.6151
R2275 B.n275 B.n274 10.6151
R2276 B.n278 B.n275 10.6151
R2277 B.n279 B.n278 10.6151
R2278 B.n282 B.n279 10.6151
R2279 B.n283 B.n282 10.6151
R2280 B.n286 B.n283 10.6151
R2281 B.n287 B.n286 10.6151
R2282 B.n290 B.n287 10.6151
R2283 B.n291 B.n290 10.6151
R2284 B.n294 B.n291 10.6151
R2285 B.n295 B.n294 10.6151
R2286 B.n298 B.n295 10.6151
R2287 B.n299 B.n298 10.6151
R2288 B.n302 B.n299 10.6151
R2289 B.n303 B.n302 10.6151
R2290 B.n306 B.n303 10.6151
R2291 B.n307 B.n306 10.6151
R2292 B.n310 B.n307 10.6151
R2293 B.n311 B.n310 10.6151
R2294 B.n314 B.n311 10.6151
R2295 B.n315 B.n314 10.6151
R2296 B.n931 B.n315 10.6151
R2297 B.n650 B.n442 10.6151
R2298 B.n651 B.n650 10.6151
R2299 B.n652 B.n651 10.6151
R2300 B.n652 B.n434 10.6151
R2301 B.n662 B.n434 10.6151
R2302 B.n663 B.n662 10.6151
R2303 B.n664 B.n663 10.6151
R2304 B.n664 B.n427 10.6151
R2305 B.n675 B.n427 10.6151
R2306 B.n676 B.n675 10.6151
R2307 B.n677 B.n676 10.6151
R2308 B.n677 B.n419 10.6151
R2309 B.n687 B.n419 10.6151
R2310 B.n688 B.n687 10.6151
R2311 B.n689 B.n688 10.6151
R2312 B.n689 B.n411 10.6151
R2313 B.n699 B.n411 10.6151
R2314 B.n700 B.n699 10.6151
R2315 B.n701 B.n700 10.6151
R2316 B.n701 B.n403 10.6151
R2317 B.n711 B.n403 10.6151
R2318 B.n712 B.n711 10.6151
R2319 B.n713 B.n712 10.6151
R2320 B.n713 B.n396 10.6151
R2321 B.n724 B.n396 10.6151
R2322 B.n725 B.n724 10.6151
R2323 B.n726 B.n725 10.6151
R2324 B.n726 B.n388 10.6151
R2325 B.n736 B.n388 10.6151
R2326 B.n737 B.n736 10.6151
R2327 B.n738 B.n737 10.6151
R2328 B.n738 B.n380 10.6151
R2329 B.n748 B.n380 10.6151
R2330 B.n749 B.n748 10.6151
R2331 B.n750 B.n749 10.6151
R2332 B.n750 B.n372 10.6151
R2333 B.n760 B.n372 10.6151
R2334 B.n761 B.n760 10.6151
R2335 B.n762 B.n761 10.6151
R2336 B.n762 B.n364 10.6151
R2337 B.n772 B.n364 10.6151
R2338 B.n773 B.n772 10.6151
R2339 B.n774 B.n773 10.6151
R2340 B.n774 B.n356 10.6151
R2341 B.n784 B.n356 10.6151
R2342 B.n785 B.n784 10.6151
R2343 B.n786 B.n785 10.6151
R2344 B.n786 B.n348 10.6151
R2345 B.n796 B.n348 10.6151
R2346 B.n797 B.n796 10.6151
R2347 B.n798 B.n797 10.6151
R2348 B.n798 B.n340 10.6151
R2349 B.n808 B.n340 10.6151
R2350 B.n809 B.n808 10.6151
R2351 B.n810 B.n809 10.6151
R2352 B.n810 B.n332 10.6151
R2353 B.n820 B.n332 10.6151
R2354 B.n821 B.n820 10.6151
R2355 B.n822 B.n821 10.6151
R2356 B.n822 B.n324 10.6151
R2357 B.n832 B.n324 10.6151
R2358 B.n833 B.n832 10.6151
R2359 B.n835 B.n833 10.6151
R2360 B.n835 B.n834 10.6151
R2361 B.n834 B.n316 10.6151
R2362 B.n846 B.n316 10.6151
R2363 B.n847 B.n846 10.6151
R2364 B.n848 B.n847 10.6151
R2365 B.n849 B.n848 10.6151
R2366 B.n851 B.n849 10.6151
R2367 B.n852 B.n851 10.6151
R2368 B.n853 B.n852 10.6151
R2369 B.n854 B.n853 10.6151
R2370 B.n856 B.n854 10.6151
R2371 B.n857 B.n856 10.6151
R2372 B.n858 B.n857 10.6151
R2373 B.n859 B.n858 10.6151
R2374 B.n861 B.n859 10.6151
R2375 B.n862 B.n861 10.6151
R2376 B.n863 B.n862 10.6151
R2377 B.n864 B.n863 10.6151
R2378 B.n866 B.n864 10.6151
R2379 B.n867 B.n866 10.6151
R2380 B.n868 B.n867 10.6151
R2381 B.n869 B.n868 10.6151
R2382 B.n871 B.n869 10.6151
R2383 B.n872 B.n871 10.6151
R2384 B.n873 B.n872 10.6151
R2385 B.n874 B.n873 10.6151
R2386 B.n876 B.n874 10.6151
R2387 B.n877 B.n876 10.6151
R2388 B.n878 B.n877 10.6151
R2389 B.n879 B.n878 10.6151
R2390 B.n881 B.n879 10.6151
R2391 B.n882 B.n881 10.6151
R2392 B.n883 B.n882 10.6151
R2393 B.n884 B.n883 10.6151
R2394 B.n886 B.n884 10.6151
R2395 B.n887 B.n886 10.6151
R2396 B.n888 B.n887 10.6151
R2397 B.n889 B.n888 10.6151
R2398 B.n891 B.n889 10.6151
R2399 B.n892 B.n891 10.6151
R2400 B.n893 B.n892 10.6151
R2401 B.n894 B.n893 10.6151
R2402 B.n896 B.n894 10.6151
R2403 B.n897 B.n896 10.6151
R2404 B.n898 B.n897 10.6151
R2405 B.n899 B.n898 10.6151
R2406 B.n901 B.n899 10.6151
R2407 B.n902 B.n901 10.6151
R2408 B.n903 B.n902 10.6151
R2409 B.n904 B.n903 10.6151
R2410 B.n906 B.n904 10.6151
R2411 B.n907 B.n906 10.6151
R2412 B.n908 B.n907 10.6151
R2413 B.n909 B.n908 10.6151
R2414 B.n911 B.n909 10.6151
R2415 B.n912 B.n911 10.6151
R2416 B.n913 B.n912 10.6151
R2417 B.n914 B.n913 10.6151
R2418 B.n916 B.n914 10.6151
R2419 B.n917 B.n916 10.6151
R2420 B.n918 B.n917 10.6151
R2421 B.n919 B.n918 10.6151
R2422 B.n921 B.n919 10.6151
R2423 B.n922 B.n921 10.6151
R2424 B.n923 B.n922 10.6151
R2425 B.n924 B.n923 10.6151
R2426 B.n926 B.n924 10.6151
R2427 B.n927 B.n926 10.6151
R2428 B.n928 B.n927 10.6151
R2429 B.n929 B.n928 10.6151
R2430 B.n930 B.n929 10.6151
R2431 B.n644 B.n446 10.6151
R2432 B.n639 B.n446 10.6151
R2433 B.n639 B.n638 10.6151
R2434 B.n638 B.n637 10.6151
R2435 B.n637 B.n634 10.6151
R2436 B.n634 B.n633 10.6151
R2437 B.n633 B.n630 10.6151
R2438 B.n630 B.n629 10.6151
R2439 B.n629 B.n626 10.6151
R2440 B.n626 B.n625 10.6151
R2441 B.n625 B.n622 10.6151
R2442 B.n622 B.n621 10.6151
R2443 B.n621 B.n618 10.6151
R2444 B.n618 B.n617 10.6151
R2445 B.n617 B.n614 10.6151
R2446 B.n614 B.n613 10.6151
R2447 B.n613 B.n610 10.6151
R2448 B.n610 B.n609 10.6151
R2449 B.n609 B.n606 10.6151
R2450 B.n606 B.n605 10.6151
R2451 B.n605 B.n602 10.6151
R2452 B.n602 B.n601 10.6151
R2453 B.n601 B.n598 10.6151
R2454 B.n598 B.n597 10.6151
R2455 B.n597 B.n594 10.6151
R2456 B.n594 B.n593 10.6151
R2457 B.n593 B.n590 10.6151
R2458 B.n590 B.n589 10.6151
R2459 B.n589 B.n586 10.6151
R2460 B.n586 B.n585 10.6151
R2461 B.n585 B.n582 10.6151
R2462 B.n582 B.n581 10.6151
R2463 B.n581 B.n578 10.6151
R2464 B.n576 B.n573 10.6151
R2465 B.n573 B.n572 10.6151
R2466 B.n572 B.n569 10.6151
R2467 B.n569 B.n568 10.6151
R2468 B.n568 B.n565 10.6151
R2469 B.n565 B.n564 10.6151
R2470 B.n564 B.n561 10.6151
R2471 B.n561 B.n560 10.6151
R2472 B.n557 B.n556 10.6151
R2473 B.n556 B.n553 10.6151
R2474 B.n553 B.n552 10.6151
R2475 B.n552 B.n549 10.6151
R2476 B.n549 B.n548 10.6151
R2477 B.n548 B.n545 10.6151
R2478 B.n545 B.n544 10.6151
R2479 B.n544 B.n541 10.6151
R2480 B.n541 B.n540 10.6151
R2481 B.n540 B.n537 10.6151
R2482 B.n537 B.n536 10.6151
R2483 B.n536 B.n533 10.6151
R2484 B.n533 B.n532 10.6151
R2485 B.n532 B.n529 10.6151
R2486 B.n529 B.n528 10.6151
R2487 B.n528 B.n525 10.6151
R2488 B.n525 B.n524 10.6151
R2489 B.n524 B.n521 10.6151
R2490 B.n521 B.n520 10.6151
R2491 B.n520 B.n517 10.6151
R2492 B.n517 B.n516 10.6151
R2493 B.n516 B.n513 10.6151
R2494 B.n513 B.n512 10.6151
R2495 B.n512 B.n509 10.6151
R2496 B.n509 B.n508 10.6151
R2497 B.n508 B.n505 10.6151
R2498 B.n505 B.n504 10.6151
R2499 B.n504 B.n501 10.6151
R2500 B.n501 B.n500 10.6151
R2501 B.n500 B.n497 10.6151
R2502 B.n497 B.n496 10.6151
R2503 B.n496 B.n493 10.6151
R2504 B.n493 B.n492 10.6151
R2505 B.n646 B.n645 10.6151
R2506 B.n646 B.n438 10.6151
R2507 B.n656 B.n438 10.6151
R2508 B.n657 B.n656 10.6151
R2509 B.n658 B.n657 10.6151
R2510 B.n658 B.n430 10.6151
R2511 B.n669 B.n430 10.6151
R2512 B.n670 B.n669 10.6151
R2513 B.n671 B.n670 10.6151
R2514 B.n671 B.n423 10.6151
R2515 B.n681 B.n423 10.6151
R2516 B.n682 B.n681 10.6151
R2517 B.n683 B.n682 10.6151
R2518 B.n683 B.n415 10.6151
R2519 B.n693 B.n415 10.6151
R2520 B.n694 B.n693 10.6151
R2521 B.n695 B.n694 10.6151
R2522 B.n695 B.n407 10.6151
R2523 B.n705 B.n407 10.6151
R2524 B.n706 B.n705 10.6151
R2525 B.n707 B.n706 10.6151
R2526 B.n707 B.n399 10.6151
R2527 B.n718 B.n399 10.6151
R2528 B.n719 B.n718 10.6151
R2529 B.n720 B.n719 10.6151
R2530 B.n720 B.n392 10.6151
R2531 B.n730 B.n392 10.6151
R2532 B.n731 B.n730 10.6151
R2533 B.n732 B.n731 10.6151
R2534 B.n732 B.n384 10.6151
R2535 B.n742 B.n384 10.6151
R2536 B.n743 B.n742 10.6151
R2537 B.n744 B.n743 10.6151
R2538 B.n744 B.n376 10.6151
R2539 B.n754 B.n376 10.6151
R2540 B.n755 B.n754 10.6151
R2541 B.n756 B.n755 10.6151
R2542 B.n756 B.n368 10.6151
R2543 B.n766 B.n368 10.6151
R2544 B.n767 B.n766 10.6151
R2545 B.n768 B.n767 10.6151
R2546 B.n768 B.n360 10.6151
R2547 B.n778 B.n360 10.6151
R2548 B.n779 B.n778 10.6151
R2549 B.n780 B.n779 10.6151
R2550 B.n780 B.n352 10.6151
R2551 B.n790 B.n352 10.6151
R2552 B.n791 B.n790 10.6151
R2553 B.n792 B.n791 10.6151
R2554 B.n792 B.n344 10.6151
R2555 B.n802 B.n344 10.6151
R2556 B.n803 B.n802 10.6151
R2557 B.n804 B.n803 10.6151
R2558 B.n804 B.n336 10.6151
R2559 B.n814 B.n336 10.6151
R2560 B.n815 B.n814 10.6151
R2561 B.n816 B.n815 10.6151
R2562 B.n816 B.n328 10.6151
R2563 B.n826 B.n328 10.6151
R2564 B.n827 B.n826 10.6151
R2565 B.n828 B.n827 10.6151
R2566 B.n828 B.n320 10.6151
R2567 B.n839 B.n320 10.6151
R2568 B.n840 B.n839 10.6151
R2569 B.n841 B.n840 10.6151
R2570 B.n841 B.n0 10.6151
R2571 B.n1066 B.n1 10.6151
R2572 B.n1066 B.n1065 10.6151
R2573 B.n1065 B.n1064 10.6151
R2574 B.n1064 B.n10 10.6151
R2575 B.n1058 B.n10 10.6151
R2576 B.n1058 B.n1057 10.6151
R2577 B.n1057 B.n1056 10.6151
R2578 B.n1056 B.n17 10.6151
R2579 B.n1050 B.n17 10.6151
R2580 B.n1050 B.n1049 10.6151
R2581 B.n1049 B.n1048 10.6151
R2582 B.n1048 B.n24 10.6151
R2583 B.n1042 B.n24 10.6151
R2584 B.n1042 B.n1041 10.6151
R2585 B.n1041 B.n1040 10.6151
R2586 B.n1040 B.n31 10.6151
R2587 B.n1034 B.n31 10.6151
R2588 B.n1034 B.n1033 10.6151
R2589 B.n1033 B.n1032 10.6151
R2590 B.n1032 B.n38 10.6151
R2591 B.n1026 B.n38 10.6151
R2592 B.n1026 B.n1025 10.6151
R2593 B.n1025 B.n1024 10.6151
R2594 B.n1024 B.n45 10.6151
R2595 B.n1018 B.n45 10.6151
R2596 B.n1018 B.n1017 10.6151
R2597 B.n1017 B.n1016 10.6151
R2598 B.n1016 B.n52 10.6151
R2599 B.n1010 B.n52 10.6151
R2600 B.n1010 B.n1009 10.6151
R2601 B.n1009 B.n1008 10.6151
R2602 B.n1008 B.n59 10.6151
R2603 B.n1002 B.n59 10.6151
R2604 B.n1002 B.n1001 10.6151
R2605 B.n1001 B.n1000 10.6151
R2606 B.n1000 B.n66 10.6151
R2607 B.n994 B.n66 10.6151
R2608 B.n994 B.n993 10.6151
R2609 B.n993 B.n992 10.6151
R2610 B.n992 B.n73 10.6151
R2611 B.n986 B.n73 10.6151
R2612 B.n986 B.n985 10.6151
R2613 B.n985 B.n984 10.6151
R2614 B.n984 B.n79 10.6151
R2615 B.n978 B.n79 10.6151
R2616 B.n978 B.n977 10.6151
R2617 B.n977 B.n976 10.6151
R2618 B.n976 B.n87 10.6151
R2619 B.n970 B.n87 10.6151
R2620 B.n970 B.n969 10.6151
R2621 B.n969 B.n968 10.6151
R2622 B.n968 B.n94 10.6151
R2623 B.n962 B.n94 10.6151
R2624 B.n962 B.n961 10.6151
R2625 B.n961 B.n960 10.6151
R2626 B.n960 B.n101 10.6151
R2627 B.n954 B.n101 10.6151
R2628 B.n954 B.n953 10.6151
R2629 B.n953 B.n952 10.6151
R2630 B.n952 B.n107 10.6151
R2631 B.n946 B.n107 10.6151
R2632 B.n946 B.n945 10.6151
R2633 B.n945 B.n944 10.6151
R2634 B.n944 B.n115 10.6151
R2635 B.n938 B.n115 10.6151
R2636 B.n938 B.n937 10.6151
R2637 B.t0 B.n374 8.27967
R2638 B.t7 B.n57 8.27967
R2639 B.n233 B.n167 6.5566
R2640 B.n250 B.n249 6.5566
R2641 B.n577 B.n576 6.5566
R2642 B.n560 B.n490 6.5566
R2643 B.n230 B.n167 4.05904
R2644 B.n251 B.n250 4.05904
R2645 B.n578 B.n577 4.05904
R2646 B.n557 B.n490 4.05904
R2647 B.n1072 B.n0 2.81026
R2648 B.n1072 B.n1 2.81026
R2649 B.n673 B.t9 0.753151
R2650 B.n715 B.t5 0.753151
R2651 B.n81 B.t4 0.753151
R2652 B.n956 B.t13 0.753151
R2653 VN.n76 VN.n75 161.3
R2654 VN.n74 VN.n40 161.3
R2655 VN.n73 VN.n72 161.3
R2656 VN.n71 VN.n41 161.3
R2657 VN.n70 VN.n69 161.3
R2658 VN.n68 VN.n42 161.3
R2659 VN.n67 VN.n66 161.3
R2660 VN.n65 VN.n43 161.3
R2661 VN.n64 VN.n63 161.3
R2662 VN.n62 VN.n44 161.3
R2663 VN.n61 VN.n60 161.3
R2664 VN.n59 VN.n46 161.3
R2665 VN.n58 VN.n57 161.3
R2666 VN.n56 VN.n47 161.3
R2667 VN.n55 VN.n54 161.3
R2668 VN.n53 VN.n48 161.3
R2669 VN.n52 VN.n51 161.3
R2670 VN.n37 VN.n36 161.3
R2671 VN.n35 VN.n1 161.3
R2672 VN.n34 VN.n33 161.3
R2673 VN.n32 VN.n2 161.3
R2674 VN.n31 VN.n30 161.3
R2675 VN.n29 VN.n3 161.3
R2676 VN.n28 VN.n27 161.3
R2677 VN.n26 VN.n4 161.3
R2678 VN.n25 VN.n24 161.3
R2679 VN.n22 VN.n5 161.3
R2680 VN.n21 VN.n20 161.3
R2681 VN.n19 VN.n6 161.3
R2682 VN.n18 VN.n17 161.3
R2683 VN.n16 VN.n7 161.3
R2684 VN.n15 VN.n14 161.3
R2685 VN.n13 VN.n8 161.3
R2686 VN.n12 VN.n11 161.3
R2687 VN.n49 VN.t3 92.5415
R2688 VN.n9 VN.t0 92.5415
R2689 VN.n38 VN.n0 88.77
R2690 VN.n77 VN.n39 88.77
R2691 VN.n50 VN.n49 74.7511
R2692 VN.n10 VN.n9 74.7511
R2693 VN.n10 VN.t7 61.0016
R2694 VN.n23 VN.t6 61.0016
R2695 VN.n0 VN.t4 61.0016
R2696 VN.n50 VN.t5 61.0016
R2697 VN.n45 VN.t1 61.0016
R2698 VN.n39 VN.t2 61.0016
R2699 VN VN.n77 54.1496
R2700 VN.n30 VN.n2 42.5146
R2701 VN.n69 VN.n41 42.5146
R2702 VN.n17 VN.n16 40.577
R2703 VN.n17 VN.n6 40.577
R2704 VN.n57 VN.n56 40.577
R2705 VN.n57 VN.n46 40.577
R2706 VN.n30 VN.n29 38.6395
R2707 VN.n69 VN.n68 38.6395
R2708 VN.n11 VN.n8 24.5923
R2709 VN.n15 VN.n8 24.5923
R2710 VN.n16 VN.n15 24.5923
R2711 VN.n21 VN.n6 24.5923
R2712 VN.n22 VN.n21 24.5923
R2713 VN.n24 VN.n22 24.5923
R2714 VN.n28 VN.n4 24.5923
R2715 VN.n29 VN.n28 24.5923
R2716 VN.n34 VN.n2 24.5923
R2717 VN.n35 VN.n34 24.5923
R2718 VN.n36 VN.n35 24.5923
R2719 VN.n56 VN.n55 24.5923
R2720 VN.n55 VN.n48 24.5923
R2721 VN.n51 VN.n48 24.5923
R2722 VN.n68 VN.n67 24.5923
R2723 VN.n67 VN.n43 24.5923
R2724 VN.n63 VN.n62 24.5923
R2725 VN.n62 VN.n61 24.5923
R2726 VN.n61 VN.n46 24.5923
R2727 VN.n75 VN.n74 24.5923
R2728 VN.n74 VN.n73 24.5923
R2729 VN.n73 VN.n41 24.5923
R2730 VN.n23 VN.n4 24.1005
R2731 VN.n45 VN.n43 24.1005
R2732 VN.n52 VN.n49 3.41205
R2733 VN.n12 VN.n9 3.41205
R2734 VN.n36 VN.n0 1.47601
R2735 VN.n75 VN.n39 1.47601
R2736 VN.n11 VN.n10 0.492337
R2737 VN.n24 VN.n23 0.492337
R2738 VN.n51 VN.n50 0.492337
R2739 VN.n63 VN.n45 0.492337
R2740 VN.n77 VN.n76 0.354861
R2741 VN.n38 VN.n37 0.354861
R2742 VN VN.n38 0.267071
R2743 VN.n76 VN.n40 0.189894
R2744 VN.n72 VN.n40 0.189894
R2745 VN.n72 VN.n71 0.189894
R2746 VN.n71 VN.n70 0.189894
R2747 VN.n70 VN.n42 0.189894
R2748 VN.n66 VN.n42 0.189894
R2749 VN.n66 VN.n65 0.189894
R2750 VN.n65 VN.n64 0.189894
R2751 VN.n64 VN.n44 0.189894
R2752 VN.n60 VN.n44 0.189894
R2753 VN.n60 VN.n59 0.189894
R2754 VN.n59 VN.n58 0.189894
R2755 VN.n58 VN.n47 0.189894
R2756 VN.n54 VN.n47 0.189894
R2757 VN.n54 VN.n53 0.189894
R2758 VN.n53 VN.n52 0.189894
R2759 VN.n13 VN.n12 0.189894
R2760 VN.n14 VN.n13 0.189894
R2761 VN.n14 VN.n7 0.189894
R2762 VN.n18 VN.n7 0.189894
R2763 VN.n19 VN.n18 0.189894
R2764 VN.n20 VN.n19 0.189894
R2765 VN.n20 VN.n5 0.189894
R2766 VN.n25 VN.n5 0.189894
R2767 VN.n26 VN.n25 0.189894
R2768 VN.n27 VN.n26 0.189894
R2769 VN.n27 VN.n3 0.189894
R2770 VN.n31 VN.n3 0.189894
R2771 VN.n32 VN.n31 0.189894
R2772 VN.n33 VN.n32 0.189894
R2773 VN.n33 VN.n1 0.189894
R2774 VN.n37 VN.n1 0.189894
R2775 VDD2.n2 VDD2.n1 66.6187
R2776 VDD2.n2 VDD2.n0 66.6187
R2777 VDD2 VDD2.n5 66.6158
R2778 VDD2.n4 VDD2.n3 64.9414
R2779 VDD2.n4 VDD2.n2 47.3618
R2780 VDD2.n5 VDD2.t2 2.12041
R2781 VDD2.n5 VDD2.t4 2.12041
R2782 VDD2.n3 VDD2.t5 2.12041
R2783 VDD2.n3 VDD2.t6 2.12041
R2784 VDD2.n1 VDD2.t1 2.12041
R2785 VDD2.n1 VDD2.t3 2.12041
R2786 VDD2.n0 VDD2.t7 2.12041
R2787 VDD2.n0 VDD2.t0 2.12041
R2788 VDD2 VDD2.n4 1.79145
C0 VP VTAIL 8.186589f
C1 VN VTAIL 8.17248f
C2 VTAIL VDD1 7.79018f
C3 VP VN 8.4993f
C4 VTAIL VDD2 7.85191f
C5 VP VDD1 7.76903f
C6 VN VDD1 0.153646f
C7 VP VDD2 0.635606f
C8 VN VDD2 7.28902f
C9 VDD1 VDD2 2.34017f
C10 VDD2 B 6.302482f
C11 VDD1 B 6.86072f
C12 VTAIL B 9.60561f
C13 VN B 19.528091f
C14 VP B 18.19447f
C15 VDD2.t7 B 0.205159f
C16 VDD2.t0 B 0.205159f
C17 VDD2.n0 B 1.81672f
C18 VDD2.t1 B 0.205159f
C19 VDD2.t3 B 0.205159f
C20 VDD2.n1 B 1.81672f
C21 VDD2.n2 B 4.15059f
C22 VDD2.t5 B 0.205159f
C23 VDD2.t6 B 0.205159f
C24 VDD2.n3 B 1.79921f
C25 VDD2.n4 B 3.47066f
C26 VDD2.t2 B 0.205159f
C27 VDD2.t4 B 0.205159f
C28 VDD2.n5 B 1.81668f
C29 VN.t4 B 1.72293f
C30 VN.n0 B 0.678226f
C31 VN.n1 B 0.018499f
C32 VN.n2 B 0.03616f
C33 VN.n3 B 0.018499f
C34 VN.n4 B 0.033965f
C35 VN.n5 B 0.018499f
C36 VN.n6 B 0.036572f
C37 VN.n7 B 0.018499f
C38 VN.n8 B 0.034304f
C39 VN.t0 B 1.97919f
C40 VN.n9 B 0.641856f
C41 VN.t7 B 1.72293f
C42 VN.n10 B 0.670485f
C43 VN.n11 B 0.017708f
C44 VN.n12 B 0.234941f
C45 VN.n13 B 0.018499f
C46 VN.n14 B 0.018499f
C47 VN.n15 B 0.034304f
C48 VN.n16 B 0.036572f
C49 VN.n17 B 0.014941f
C50 VN.n18 B 0.018499f
C51 VN.n19 B 0.018499f
C52 VN.n20 B 0.018499f
C53 VN.n21 B 0.034304f
C54 VN.n22 B 0.034304f
C55 VN.t6 B 1.72293f
C56 VN.n23 B 0.612499f
C57 VN.n24 B 0.017708f
C58 VN.n25 B 0.018499f
C59 VN.n26 B 0.018499f
C60 VN.n27 B 0.018499f
C61 VN.n28 B 0.034304f
C62 VN.n29 B 0.03689f
C63 VN.n30 B 0.015035f
C64 VN.n31 B 0.018499f
C65 VN.n32 B 0.018499f
C66 VN.n33 B 0.018499f
C67 VN.n34 B 0.034304f
C68 VN.n35 B 0.034304f
C69 VN.n36 B 0.018385f
C70 VN.n37 B 0.029851f
C71 VN.n38 B 0.056336f
C72 VN.t2 B 1.72293f
C73 VN.n39 B 0.678226f
C74 VN.n40 B 0.018499f
C75 VN.n41 B 0.03616f
C76 VN.n42 B 0.018499f
C77 VN.n43 B 0.033965f
C78 VN.n44 B 0.018499f
C79 VN.t1 B 1.72293f
C80 VN.n45 B 0.612499f
C81 VN.n46 B 0.036572f
C82 VN.n47 B 0.018499f
C83 VN.n48 B 0.034304f
C84 VN.t3 B 1.97919f
C85 VN.n49 B 0.641856f
C86 VN.t5 B 1.72293f
C87 VN.n50 B 0.670485f
C88 VN.n51 B 0.017708f
C89 VN.n52 B 0.234941f
C90 VN.n53 B 0.018499f
C91 VN.n54 B 0.018499f
C92 VN.n55 B 0.034304f
C93 VN.n56 B 0.036572f
C94 VN.n57 B 0.014941f
C95 VN.n58 B 0.018499f
C96 VN.n59 B 0.018499f
C97 VN.n60 B 0.018499f
C98 VN.n61 B 0.034304f
C99 VN.n62 B 0.034304f
C100 VN.n63 B 0.017708f
C101 VN.n64 B 0.018499f
C102 VN.n65 B 0.018499f
C103 VN.n66 B 0.018499f
C104 VN.n67 B 0.034304f
C105 VN.n68 B 0.03689f
C106 VN.n69 B 0.015035f
C107 VN.n70 B 0.018499f
C108 VN.n71 B 0.018499f
C109 VN.n72 B 0.018499f
C110 VN.n73 B 0.034304f
C111 VN.n74 B 0.034304f
C112 VN.n75 B 0.018385f
C113 VN.n76 B 0.029851f
C114 VN.n77 B 1.19083f
C115 VTAIL.t6 B 0.161771f
C116 VTAIL.t7 B 0.161771f
C117 VTAIL.n0 B 1.35919f
C118 VTAIL.n1 B 0.45492f
C119 VTAIL.n2 B 0.02992f
C120 VTAIL.n3 B 0.021918f
C121 VTAIL.n4 B 0.011778f
C122 VTAIL.n5 B 0.027838f
C123 VTAIL.n6 B 0.012124f
C124 VTAIL.n7 B 0.021918f
C125 VTAIL.n8 B 0.012471f
C126 VTAIL.n9 B 0.027838f
C127 VTAIL.n10 B 0.012471f
C128 VTAIL.n11 B 0.021918f
C129 VTAIL.n12 B 0.011778f
C130 VTAIL.n13 B 0.027838f
C131 VTAIL.n14 B 0.012471f
C132 VTAIL.n15 B 0.846394f
C133 VTAIL.n16 B 0.011778f
C134 VTAIL.t2 B 0.046707f
C135 VTAIL.n17 B 0.135649f
C136 VTAIL.n18 B 0.019679f
C137 VTAIL.n19 B 0.020879f
C138 VTAIL.n20 B 0.027838f
C139 VTAIL.n21 B 0.012471f
C140 VTAIL.n22 B 0.011778f
C141 VTAIL.n23 B 0.021918f
C142 VTAIL.n24 B 0.021918f
C143 VTAIL.n25 B 0.011778f
C144 VTAIL.n26 B 0.012471f
C145 VTAIL.n27 B 0.027838f
C146 VTAIL.n28 B 0.027838f
C147 VTAIL.n29 B 0.012471f
C148 VTAIL.n30 B 0.011778f
C149 VTAIL.n31 B 0.021918f
C150 VTAIL.n32 B 0.021918f
C151 VTAIL.n33 B 0.011778f
C152 VTAIL.n34 B 0.011778f
C153 VTAIL.n35 B 0.012471f
C154 VTAIL.n36 B 0.027838f
C155 VTAIL.n37 B 0.027838f
C156 VTAIL.n38 B 0.027838f
C157 VTAIL.n39 B 0.012124f
C158 VTAIL.n40 B 0.011778f
C159 VTAIL.n41 B 0.021918f
C160 VTAIL.n42 B 0.021918f
C161 VTAIL.n43 B 0.011778f
C162 VTAIL.n44 B 0.012471f
C163 VTAIL.n45 B 0.027838f
C164 VTAIL.n46 B 0.058696f
C165 VTAIL.n47 B 0.012471f
C166 VTAIL.n48 B 0.011778f
C167 VTAIL.n49 B 0.053657f
C168 VTAIL.n50 B 0.032771f
C169 VTAIL.n51 B 0.298344f
C170 VTAIL.n52 B 0.02992f
C171 VTAIL.n53 B 0.021918f
C172 VTAIL.n54 B 0.011778f
C173 VTAIL.n55 B 0.027838f
C174 VTAIL.n56 B 0.012124f
C175 VTAIL.n57 B 0.021918f
C176 VTAIL.n58 B 0.012471f
C177 VTAIL.n59 B 0.027838f
C178 VTAIL.n60 B 0.012471f
C179 VTAIL.n61 B 0.021918f
C180 VTAIL.n62 B 0.011778f
C181 VTAIL.n63 B 0.027838f
C182 VTAIL.n64 B 0.012471f
C183 VTAIL.n65 B 0.846394f
C184 VTAIL.n66 B 0.011778f
C185 VTAIL.t9 B 0.046707f
C186 VTAIL.n67 B 0.135649f
C187 VTAIL.n68 B 0.019679f
C188 VTAIL.n69 B 0.020879f
C189 VTAIL.n70 B 0.027838f
C190 VTAIL.n71 B 0.012471f
C191 VTAIL.n72 B 0.011778f
C192 VTAIL.n73 B 0.021918f
C193 VTAIL.n74 B 0.021918f
C194 VTAIL.n75 B 0.011778f
C195 VTAIL.n76 B 0.012471f
C196 VTAIL.n77 B 0.027838f
C197 VTAIL.n78 B 0.027838f
C198 VTAIL.n79 B 0.012471f
C199 VTAIL.n80 B 0.011778f
C200 VTAIL.n81 B 0.021918f
C201 VTAIL.n82 B 0.021918f
C202 VTAIL.n83 B 0.011778f
C203 VTAIL.n84 B 0.011778f
C204 VTAIL.n85 B 0.012471f
C205 VTAIL.n86 B 0.027838f
C206 VTAIL.n87 B 0.027838f
C207 VTAIL.n88 B 0.027838f
C208 VTAIL.n89 B 0.012124f
C209 VTAIL.n90 B 0.011778f
C210 VTAIL.n91 B 0.021918f
C211 VTAIL.n92 B 0.021918f
C212 VTAIL.n93 B 0.011778f
C213 VTAIL.n94 B 0.012471f
C214 VTAIL.n95 B 0.027838f
C215 VTAIL.n96 B 0.058696f
C216 VTAIL.n97 B 0.012471f
C217 VTAIL.n98 B 0.011778f
C218 VTAIL.n99 B 0.053657f
C219 VTAIL.n100 B 0.032771f
C220 VTAIL.n101 B 0.298344f
C221 VTAIL.t11 B 0.161771f
C222 VTAIL.t8 B 0.161771f
C223 VTAIL.n102 B 1.35919f
C224 VTAIL.n103 B 0.695561f
C225 VTAIL.n104 B 0.02992f
C226 VTAIL.n105 B 0.021918f
C227 VTAIL.n106 B 0.011778f
C228 VTAIL.n107 B 0.027838f
C229 VTAIL.n108 B 0.012124f
C230 VTAIL.n109 B 0.021918f
C231 VTAIL.n110 B 0.012471f
C232 VTAIL.n111 B 0.027838f
C233 VTAIL.n112 B 0.012471f
C234 VTAIL.n113 B 0.021918f
C235 VTAIL.n114 B 0.011778f
C236 VTAIL.n115 B 0.027838f
C237 VTAIL.n116 B 0.012471f
C238 VTAIL.n117 B 0.846394f
C239 VTAIL.n118 B 0.011778f
C240 VTAIL.t13 B 0.046707f
C241 VTAIL.n119 B 0.135649f
C242 VTAIL.n120 B 0.019679f
C243 VTAIL.n121 B 0.020879f
C244 VTAIL.n122 B 0.027838f
C245 VTAIL.n123 B 0.012471f
C246 VTAIL.n124 B 0.011778f
C247 VTAIL.n125 B 0.021918f
C248 VTAIL.n126 B 0.021918f
C249 VTAIL.n127 B 0.011778f
C250 VTAIL.n128 B 0.012471f
C251 VTAIL.n129 B 0.027838f
C252 VTAIL.n130 B 0.027838f
C253 VTAIL.n131 B 0.012471f
C254 VTAIL.n132 B 0.011778f
C255 VTAIL.n133 B 0.021918f
C256 VTAIL.n134 B 0.021918f
C257 VTAIL.n135 B 0.011778f
C258 VTAIL.n136 B 0.011778f
C259 VTAIL.n137 B 0.012471f
C260 VTAIL.n138 B 0.027838f
C261 VTAIL.n139 B 0.027838f
C262 VTAIL.n140 B 0.027838f
C263 VTAIL.n141 B 0.012124f
C264 VTAIL.n142 B 0.011778f
C265 VTAIL.n143 B 0.021918f
C266 VTAIL.n144 B 0.021918f
C267 VTAIL.n145 B 0.011778f
C268 VTAIL.n146 B 0.012471f
C269 VTAIL.n147 B 0.027838f
C270 VTAIL.n148 B 0.058696f
C271 VTAIL.n149 B 0.012471f
C272 VTAIL.n150 B 0.011778f
C273 VTAIL.n151 B 0.053657f
C274 VTAIL.n152 B 0.032771f
C275 VTAIL.n153 B 1.37629f
C276 VTAIL.n154 B 0.02992f
C277 VTAIL.n155 B 0.021918f
C278 VTAIL.n156 B 0.011778f
C279 VTAIL.n157 B 0.027838f
C280 VTAIL.n158 B 0.012124f
C281 VTAIL.n159 B 0.021918f
C282 VTAIL.n160 B 0.012124f
C283 VTAIL.n161 B 0.011778f
C284 VTAIL.n162 B 0.027838f
C285 VTAIL.n163 B 0.027838f
C286 VTAIL.n164 B 0.012471f
C287 VTAIL.n165 B 0.021918f
C288 VTAIL.n166 B 0.011778f
C289 VTAIL.n167 B 0.027838f
C290 VTAIL.n168 B 0.012471f
C291 VTAIL.n169 B 0.846394f
C292 VTAIL.n170 B 0.011778f
C293 VTAIL.t5 B 0.046707f
C294 VTAIL.n171 B 0.135649f
C295 VTAIL.n172 B 0.019679f
C296 VTAIL.n173 B 0.020879f
C297 VTAIL.n174 B 0.027838f
C298 VTAIL.n175 B 0.012471f
C299 VTAIL.n176 B 0.011778f
C300 VTAIL.n177 B 0.021918f
C301 VTAIL.n178 B 0.021918f
C302 VTAIL.n179 B 0.011778f
C303 VTAIL.n180 B 0.012471f
C304 VTAIL.n181 B 0.027838f
C305 VTAIL.n182 B 0.027838f
C306 VTAIL.n183 B 0.012471f
C307 VTAIL.n184 B 0.011778f
C308 VTAIL.n185 B 0.021918f
C309 VTAIL.n186 B 0.021918f
C310 VTAIL.n187 B 0.011778f
C311 VTAIL.n188 B 0.012471f
C312 VTAIL.n189 B 0.027838f
C313 VTAIL.n190 B 0.027838f
C314 VTAIL.n191 B 0.012471f
C315 VTAIL.n192 B 0.011778f
C316 VTAIL.n193 B 0.021918f
C317 VTAIL.n194 B 0.021918f
C318 VTAIL.n195 B 0.011778f
C319 VTAIL.n196 B 0.012471f
C320 VTAIL.n197 B 0.027838f
C321 VTAIL.n198 B 0.058696f
C322 VTAIL.n199 B 0.012471f
C323 VTAIL.n200 B 0.011778f
C324 VTAIL.n201 B 0.053657f
C325 VTAIL.n202 B 0.032771f
C326 VTAIL.n203 B 1.37629f
C327 VTAIL.t0 B 0.161771f
C328 VTAIL.t3 B 0.161771f
C329 VTAIL.n204 B 1.3592f
C330 VTAIL.n205 B 0.695553f
C331 VTAIL.n206 B 0.02992f
C332 VTAIL.n207 B 0.021918f
C333 VTAIL.n208 B 0.011778f
C334 VTAIL.n209 B 0.027838f
C335 VTAIL.n210 B 0.012124f
C336 VTAIL.n211 B 0.021918f
C337 VTAIL.n212 B 0.012124f
C338 VTAIL.n213 B 0.011778f
C339 VTAIL.n214 B 0.027838f
C340 VTAIL.n215 B 0.027838f
C341 VTAIL.n216 B 0.012471f
C342 VTAIL.n217 B 0.021918f
C343 VTAIL.n218 B 0.011778f
C344 VTAIL.n219 B 0.027838f
C345 VTAIL.n220 B 0.012471f
C346 VTAIL.n221 B 0.846394f
C347 VTAIL.n222 B 0.011778f
C348 VTAIL.t1 B 0.046707f
C349 VTAIL.n223 B 0.135649f
C350 VTAIL.n224 B 0.019679f
C351 VTAIL.n225 B 0.020879f
C352 VTAIL.n226 B 0.027838f
C353 VTAIL.n227 B 0.012471f
C354 VTAIL.n228 B 0.011778f
C355 VTAIL.n229 B 0.021918f
C356 VTAIL.n230 B 0.021918f
C357 VTAIL.n231 B 0.011778f
C358 VTAIL.n232 B 0.012471f
C359 VTAIL.n233 B 0.027838f
C360 VTAIL.n234 B 0.027838f
C361 VTAIL.n235 B 0.012471f
C362 VTAIL.n236 B 0.011778f
C363 VTAIL.n237 B 0.021918f
C364 VTAIL.n238 B 0.021918f
C365 VTAIL.n239 B 0.011778f
C366 VTAIL.n240 B 0.012471f
C367 VTAIL.n241 B 0.027838f
C368 VTAIL.n242 B 0.027838f
C369 VTAIL.n243 B 0.012471f
C370 VTAIL.n244 B 0.011778f
C371 VTAIL.n245 B 0.021918f
C372 VTAIL.n246 B 0.021918f
C373 VTAIL.n247 B 0.011778f
C374 VTAIL.n248 B 0.012471f
C375 VTAIL.n249 B 0.027838f
C376 VTAIL.n250 B 0.058696f
C377 VTAIL.n251 B 0.012471f
C378 VTAIL.n252 B 0.011778f
C379 VTAIL.n253 B 0.053657f
C380 VTAIL.n254 B 0.032771f
C381 VTAIL.n255 B 0.298344f
C382 VTAIL.n256 B 0.02992f
C383 VTAIL.n257 B 0.021918f
C384 VTAIL.n258 B 0.011778f
C385 VTAIL.n259 B 0.027838f
C386 VTAIL.n260 B 0.012124f
C387 VTAIL.n261 B 0.021918f
C388 VTAIL.n262 B 0.012124f
C389 VTAIL.n263 B 0.011778f
C390 VTAIL.n264 B 0.027838f
C391 VTAIL.n265 B 0.027838f
C392 VTAIL.n266 B 0.012471f
C393 VTAIL.n267 B 0.021918f
C394 VTAIL.n268 B 0.011778f
C395 VTAIL.n269 B 0.027838f
C396 VTAIL.n270 B 0.012471f
C397 VTAIL.n271 B 0.846394f
C398 VTAIL.n272 B 0.011778f
C399 VTAIL.t15 B 0.046707f
C400 VTAIL.n273 B 0.135649f
C401 VTAIL.n274 B 0.019679f
C402 VTAIL.n275 B 0.020879f
C403 VTAIL.n276 B 0.027838f
C404 VTAIL.n277 B 0.012471f
C405 VTAIL.n278 B 0.011778f
C406 VTAIL.n279 B 0.021918f
C407 VTAIL.n280 B 0.021918f
C408 VTAIL.n281 B 0.011778f
C409 VTAIL.n282 B 0.012471f
C410 VTAIL.n283 B 0.027838f
C411 VTAIL.n284 B 0.027838f
C412 VTAIL.n285 B 0.012471f
C413 VTAIL.n286 B 0.011778f
C414 VTAIL.n287 B 0.021918f
C415 VTAIL.n288 B 0.021918f
C416 VTAIL.n289 B 0.011778f
C417 VTAIL.n290 B 0.012471f
C418 VTAIL.n291 B 0.027838f
C419 VTAIL.n292 B 0.027838f
C420 VTAIL.n293 B 0.012471f
C421 VTAIL.n294 B 0.011778f
C422 VTAIL.n295 B 0.021918f
C423 VTAIL.n296 B 0.021918f
C424 VTAIL.n297 B 0.011778f
C425 VTAIL.n298 B 0.012471f
C426 VTAIL.n299 B 0.027838f
C427 VTAIL.n300 B 0.058696f
C428 VTAIL.n301 B 0.012471f
C429 VTAIL.n302 B 0.011778f
C430 VTAIL.n303 B 0.053657f
C431 VTAIL.n304 B 0.032771f
C432 VTAIL.n305 B 0.298344f
C433 VTAIL.t14 B 0.161771f
C434 VTAIL.t12 B 0.161771f
C435 VTAIL.n306 B 1.3592f
C436 VTAIL.n307 B 0.695553f
C437 VTAIL.n308 B 0.02992f
C438 VTAIL.n309 B 0.021918f
C439 VTAIL.n310 B 0.011778f
C440 VTAIL.n311 B 0.027838f
C441 VTAIL.n312 B 0.012124f
C442 VTAIL.n313 B 0.021918f
C443 VTAIL.n314 B 0.012124f
C444 VTAIL.n315 B 0.011778f
C445 VTAIL.n316 B 0.027838f
C446 VTAIL.n317 B 0.027838f
C447 VTAIL.n318 B 0.012471f
C448 VTAIL.n319 B 0.021918f
C449 VTAIL.n320 B 0.011778f
C450 VTAIL.n321 B 0.027838f
C451 VTAIL.n322 B 0.012471f
C452 VTAIL.n323 B 0.846394f
C453 VTAIL.n324 B 0.011778f
C454 VTAIL.t10 B 0.046707f
C455 VTAIL.n325 B 0.135649f
C456 VTAIL.n326 B 0.019679f
C457 VTAIL.n327 B 0.020879f
C458 VTAIL.n328 B 0.027838f
C459 VTAIL.n329 B 0.012471f
C460 VTAIL.n330 B 0.011778f
C461 VTAIL.n331 B 0.021918f
C462 VTAIL.n332 B 0.021918f
C463 VTAIL.n333 B 0.011778f
C464 VTAIL.n334 B 0.012471f
C465 VTAIL.n335 B 0.027838f
C466 VTAIL.n336 B 0.027838f
C467 VTAIL.n337 B 0.012471f
C468 VTAIL.n338 B 0.011778f
C469 VTAIL.n339 B 0.021918f
C470 VTAIL.n340 B 0.021918f
C471 VTAIL.n341 B 0.011778f
C472 VTAIL.n342 B 0.012471f
C473 VTAIL.n343 B 0.027838f
C474 VTAIL.n344 B 0.027838f
C475 VTAIL.n345 B 0.012471f
C476 VTAIL.n346 B 0.011778f
C477 VTAIL.n347 B 0.021918f
C478 VTAIL.n348 B 0.021918f
C479 VTAIL.n349 B 0.011778f
C480 VTAIL.n350 B 0.012471f
C481 VTAIL.n351 B 0.027838f
C482 VTAIL.n352 B 0.058696f
C483 VTAIL.n353 B 0.012471f
C484 VTAIL.n354 B 0.011778f
C485 VTAIL.n355 B 0.053657f
C486 VTAIL.n356 B 0.032771f
C487 VTAIL.n357 B 1.37629f
C488 VTAIL.n358 B 0.02992f
C489 VTAIL.n359 B 0.021918f
C490 VTAIL.n360 B 0.011778f
C491 VTAIL.n361 B 0.027838f
C492 VTAIL.n362 B 0.012124f
C493 VTAIL.n363 B 0.021918f
C494 VTAIL.n364 B 0.012471f
C495 VTAIL.n365 B 0.027838f
C496 VTAIL.n366 B 0.012471f
C497 VTAIL.n367 B 0.021918f
C498 VTAIL.n368 B 0.011778f
C499 VTAIL.n369 B 0.027838f
C500 VTAIL.n370 B 0.012471f
C501 VTAIL.n371 B 0.846394f
C502 VTAIL.n372 B 0.011778f
C503 VTAIL.t4 B 0.046707f
C504 VTAIL.n373 B 0.135649f
C505 VTAIL.n374 B 0.019679f
C506 VTAIL.n375 B 0.020879f
C507 VTAIL.n376 B 0.027838f
C508 VTAIL.n377 B 0.012471f
C509 VTAIL.n378 B 0.011778f
C510 VTAIL.n379 B 0.021918f
C511 VTAIL.n380 B 0.021918f
C512 VTAIL.n381 B 0.011778f
C513 VTAIL.n382 B 0.012471f
C514 VTAIL.n383 B 0.027838f
C515 VTAIL.n384 B 0.027838f
C516 VTAIL.n385 B 0.012471f
C517 VTAIL.n386 B 0.011778f
C518 VTAIL.n387 B 0.021918f
C519 VTAIL.n388 B 0.021918f
C520 VTAIL.n389 B 0.011778f
C521 VTAIL.n390 B 0.011778f
C522 VTAIL.n391 B 0.012471f
C523 VTAIL.n392 B 0.027838f
C524 VTAIL.n393 B 0.027838f
C525 VTAIL.n394 B 0.027838f
C526 VTAIL.n395 B 0.012124f
C527 VTAIL.n396 B 0.011778f
C528 VTAIL.n397 B 0.021918f
C529 VTAIL.n398 B 0.021918f
C530 VTAIL.n399 B 0.011778f
C531 VTAIL.n400 B 0.012471f
C532 VTAIL.n401 B 0.027838f
C533 VTAIL.n402 B 0.058696f
C534 VTAIL.n403 B 0.012471f
C535 VTAIL.n404 B 0.011778f
C536 VTAIL.n405 B 0.053657f
C537 VTAIL.n406 B 0.032771f
C538 VTAIL.n407 B 1.37218f
C539 VDD1.t6 B 0.208625f
C540 VDD1.t5 B 0.208625f
C541 VDD1.n0 B 1.84886f
C542 VDD1.t4 B 0.208625f
C543 VDD1.t2 B 0.208625f
C544 VDD1.n1 B 1.84741f
C545 VDD1.t0 B 0.208625f
C546 VDD1.t7 B 0.208625f
C547 VDD1.n2 B 1.84741f
C548 VDD1.n3 B 4.27902f
C549 VDD1.t3 B 0.208625f
C550 VDD1.t1 B 0.208625f
C551 VDD1.n4 B 1.82959f
C552 VDD1.n5 B 3.56476f
C553 VP.t6 B 1.76073f
C554 VP.n0 B 0.693107f
C555 VP.n1 B 0.018904f
C556 VP.n2 B 0.036953f
C557 VP.n3 B 0.018904f
C558 VP.n4 B 0.03471f
C559 VP.n5 B 0.018904f
C560 VP.n6 B 0.037374f
C561 VP.n7 B 0.018904f
C562 VP.n8 B 0.035056f
C563 VP.n9 B 0.018904f
C564 VP.t4 B 1.76073f
C565 VP.n10 B 0.037699f
C566 VP.n11 B 0.018904f
C567 VP.n12 B 0.035056f
C568 VP.t5 B 1.76073f
C569 VP.n13 B 0.693107f
C570 VP.n14 B 0.018904f
C571 VP.n15 B 0.036953f
C572 VP.n16 B 0.018904f
C573 VP.n17 B 0.03471f
C574 VP.n18 B 0.018904f
C575 VP.n19 B 0.037374f
C576 VP.n20 B 0.018904f
C577 VP.n21 B 0.035056f
C578 VP.t0 B 2.02261f
C579 VP.n22 B 0.655939f
C580 VP.t1 B 1.76073f
C581 VP.n23 B 0.685196f
C582 VP.n24 B 0.018096f
C583 VP.n25 B 0.240096f
C584 VP.n26 B 0.018904f
C585 VP.n27 B 0.018904f
C586 VP.n28 B 0.035056f
C587 VP.n29 B 0.037374f
C588 VP.n30 B 0.015268f
C589 VP.n31 B 0.018904f
C590 VP.n32 B 0.018904f
C591 VP.n33 B 0.018904f
C592 VP.n34 B 0.035056f
C593 VP.n35 B 0.035056f
C594 VP.t3 B 1.76073f
C595 VP.n36 B 0.625938f
C596 VP.n37 B 0.018096f
C597 VP.n38 B 0.018904f
C598 VP.n39 B 0.018904f
C599 VP.n40 B 0.018904f
C600 VP.n41 B 0.035056f
C601 VP.n42 B 0.037699f
C602 VP.n43 B 0.015365f
C603 VP.n44 B 0.018904f
C604 VP.n45 B 0.018904f
C605 VP.n46 B 0.018904f
C606 VP.n47 B 0.035056f
C607 VP.n48 B 0.035056f
C608 VP.n49 B 0.018788f
C609 VP.n50 B 0.030506f
C610 VP.n51 B 1.20942f
C611 VP.n52 B 1.22204f
C612 VP.t2 B 1.76073f
C613 VP.n53 B 0.693107f
C614 VP.n54 B 0.018788f
C615 VP.n55 B 0.030506f
C616 VP.n56 B 0.018904f
C617 VP.n57 B 0.018904f
C618 VP.n58 B 0.035056f
C619 VP.n59 B 0.036953f
C620 VP.n60 B 0.015365f
C621 VP.n61 B 0.018904f
C622 VP.n62 B 0.018904f
C623 VP.n63 B 0.018904f
C624 VP.n64 B 0.035056f
C625 VP.n65 B 0.03471f
C626 VP.n66 B 0.625938f
C627 VP.n67 B 0.018096f
C628 VP.n68 B 0.018904f
C629 VP.n69 B 0.018904f
C630 VP.n70 B 0.018904f
C631 VP.n71 B 0.035056f
C632 VP.n72 B 0.037374f
C633 VP.n73 B 0.015268f
C634 VP.n74 B 0.018904f
C635 VP.n75 B 0.018904f
C636 VP.n76 B 0.018904f
C637 VP.n77 B 0.035056f
C638 VP.n78 B 0.035056f
C639 VP.t7 B 1.76073f
C640 VP.n79 B 0.625938f
C641 VP.n80 B 0.018096f
C642 VP.n81 B 0.018904f
C643 VP.n82 B 0.018904f
C644 VP.n83 B 0.018904f
C645 VP.n84 B 0.035056f
C646 VP.n85 B 0.037699f
C647 VP.n86 B 0.015365f
C648 VP.n87 B 0.018904f
C649 VP.n88 B 0.018904f
C650 VP.n89 B 0.018904f
C651 VP.n90 B 0.035056f
C652 VP.n91 B 0.035056f
C653 VP.n92 B 0.018788f
C654 VP.n93 B 0.030506f
C655 VP.n94 B 0.057573f
.ends

