* NGSPICE file created from diff_pair_sample_1462.ext - technology: sky130A

.subckt diff_pair_sample_1462 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t7 VN.t0 VTAIL.t13 w_n1900_n2652# sky130_fd_pr__pfet_01v8 ad=1.3893 pd=8.75 as=3.2838 ps=17.62 w=8.42 l=0.6
X1 VDD1.t7 VP.t0 VTAIL.t6 w_n1900_n2652# sky130_fd_pr__pfet_01v8 ad=1.3893 pd=8.75 as=3.2838 ps=17.62 w=8.42 l=0.6
X2 VTAIL.t3 VP.t1 VDD1.t6 w_n1900_n2652# sky130_fd_pr__pfet_01v8 ad=3.2838 pd=17.62 as=1.3893 ps=8.75 w=8.42 l=0.6
X3 B.t11 B.t9 B.t10 w_n1900_n2652# sky130_fd_pr__pfet_01v8 ad=3.2838 pd=17.62 as=0 ps=0 w=8.42 l=0.6
X4 VTAIL.t9 VN.t1 VDD2.t6 w_n1900_n2652# sky130_fd_pr__pfet_01v8 ad=3.2838 pd=17.62 as=1.3893 ps=8.75 w=8.42 l=0.6
X5 VDD2.t5 VN.t2 VTAIL.t10 w_n1900_n2652# sky130_fd_pr__pfet_01v8 ad=1.3893 pd=8.75 as=1.3893 ps=8.75 w=8.42 l=0.6
X6 VDD2.t4 VN.t3 VTAIL.t14 w_n1900_n2652# sky130_fd_pr__pfet_01v8 ad=1.3893 pd=8.75 as=1.3893 ps=8.75 w=8.42 l=0.6
X7 B.t8 B.t6 B.t7 w_n1900_n2652# sky130_fd_pr__pfet_01v8 ad=3.2838 pd=17.62 as=0 ps=0 w=8.42 l=0.6
X8 VDD1.t5 VP.t2 VTAIL.t1 w_n1900_n2652# sky130_fd_pr__pfet_01v8 ad=1.3893 pd=8.75 as=3.2838 ps=17.62 w=8.42 l=0.6
X9 VDD2.t3 VN.t4 VTAIL.t11 w_n1900_n2652# sky130_fd_pr__pfet_01v8 ad=1.3893 pd=8.75 as=3.2838 ps=17.62 w=8.42 l=0.6
X10 VTAIL.t15 VN.t5 VDD2.t2 w_n1900_n2652# sky130_fd_pr__pfet_01v8 ad=1.3893 pd=8.75 as=1.3893 ps=8.75 w=8.42 l=0.6
X11 VTAIL.t2 VP.t3 VDD1.t4 w_n1900_n2652# sky130_fd_pr__pfet_01v8 ad=1.3893 pd=8.75 as=1.3893 ps=8.75 w=8.42 l=0.6
X12 VDD1.t3 VP.t4 VTAIL.t5 w_n1900_n2652# sky130_fd_pr__pfet_01v8 ad=1.3893 pd=8.75 as=1.3893 ps=8.75 w=8.42 l=0.6
X13 VTAIL.t4 VP.t5 VDD1.t2 w_n1900_n2652# sky130_fd_pr__pfet_01v8 ad=3.2838 pd=17.62 as=1.3893 ps=8.75 w=8.42 l=0.6
X14 VTAIL.t8 VN.t6 VDD2.t1 w_n1900_n2652# sky130_fd_pr__pfet_01v8 ad=1.3893 pd=8.75 as=1.3893 ps=8.75 w=8.42 l=0.6
X15 VTAIL.t7 VP.t6 VDD1.t1 w_n1900_n2652# sky130_fd_pr__pfet_01v8 ad=1.3893 pd=8.75 as=1.3893 ps=8.75 w=8.42 l=0.6
X16 B.t5 B.t3 B.t4 w_n1900_n2652# sky130_fd_pr__pfet_01v8 ad=3.2838 pd=17.62 as=0 ps=0 w=8.42 l=0.6
X17 VTAIL.t12 VN.t7 VDD2.t0 w_n1900_n2652# sky130_fd_pr__pfet_01v8 ad=3.2838 pd=17.62 as=1.3893 ps=8.75 w=8.42 l=0.6
X18 VDD1.t0 VP.t7 VTAIL.t0 w_n1900_n2652# sky130_fd_pr__pfet_01v8 ad=1.3893 pd=8.75 as=1.3893 ps=8.75 w=8.42 l=0.6
X19 B.t2 B.t0 B.t1 w_n1900_n2652# sky130_fd_pr__pfet_01v8 ad=3.2838 pd=17.62 as=0 ps=0 w=8.42 l=0.6
R0 VN.n1 VN.t7 430.497
R1 VN.n7 VN.t4 430.497
R2 VN.n2 VN.t2 403.675
R3 VN.n3 VN.t6 403.675
R4 VN.n4 VN.t0 403.675
R5 VN.n8 VN.t5 403.675
R6 VN.n9 VN.t3 403.675
R7 VN.n10 VN.t1 403.675
R8 VN.n5 VN.n4 161.3
R9 VN.n11 VN.n10 161.3
R10 VN.n9 VN.n6 80.6037
R11 VN.n3 VN.n0 80.6037
R12 VN.n3 VN.n2 48.2005
R13 VN.n4 VN.n3 48.2005
R14 VN.n9 VN.n8 48.2005
R15 VN.n10 VN.n9 48.2005
R16 VN.n7 VN.n6 45.2318
R17 VN.n1 VN.n0 45.2318
R18 VN VN.n11 39.2448
R19 VN.n8 VN.n7 13.3799
R20 VN.n2 VN.n1 13.3799
R21 VN.n11 VN.n6 0.285035
R22 VN.n5 VN.n0 0.285035
R23 VN VN.n5 0.0516364
R24 VTAIL.n11 VTAIL.t4 66.9415
R25 VTAIL.n10 VTAIL.t11 66.9415
R26 VTAIL.n7 VTAIL.t9 66.9415
R27 VTAIL.n14 VTAIL.t1 66.9415
R28 VTAIL.n15 VTAIL.t13 66.9413
R29 VTAIL.n2 VTAIL.t12 66.9413
R30 VTAIL.n3 VTAIL.t6 66.9413
R31 VTAIL.n6 VTAIL.t3 66.9413
R32 VTAIL.n13 VTAIL.n12 63.0811
R33 VTAIL.n9 VTAIL.n8 63.0811
R34 VTAIL.n1 VTAIL.n0 63.081
R35 VTAIL.n5 VTAIL.n4 63.081
R36 VTAIL.n15 VTAIL.n14 20.4272
R37 VTAIL.n7 VTAIL.n6 20.4272
R38 VTAIL.n0 VTAIL.t10 3.86095
R39 VTAIL.n0 VTAIL.t8 3.86095
R40 VTAIL.n4 VTAIL.t0 3.86095
R41 VTAIL.n4 VTAIL.t7 3.86095
R42 VTAIL.n12 VTAIL.t5 3.86095
R43 VTAIL.n12 VTAIL.t2 3.86095
R44 VTAIL.n8 VTAIL.t14 3.86095
R45 VTAIL.n8 VTAIL.t15 3.86095
R46 VTAIL.n9 VTAIL.n7 0.802224
R47 VTAIL.n10 VTAIL.n9 0.802224
R48 VTAIL.n13 VTAIL.n11 0.802224
R49 VTAIL.n14 VTAIL.n13 0.802224
R50 VTAIL.n6 VTAIL.n5 0.802224
R51 VTAIL.n5 VTAIL.n3 0.802224
R52 VTAIL.n2 VTAIL.n1 0.802224
R53 VTAIL VTAIL.n15 0.744035
R54 VTAIL.n11 VTAIL.n10 0.470328
R55 VTAIL.n3 VTAIL.n2 0.470328
R56 VTAIL VTAIL.n1 0.0586897
R57 VDD2.n2 VDD2.n1 80.1053
R58 VDD2.n2 VDD2.n0 80.1053
R59 VDD2 VDD2.n5 80.1025
R60 VDD2.n4 VDD2.n3 79.7598
R61 VDD2.n4 VDD2.n2 34.5817
R62 VDD2.n5 VDD2.t2 3.86095
R63 VDD2.n5 VDD2.t3 3.86095
R64 VDD2.n3 VDD2.t6 3.86095
R65 VDD2.n3 VDD2.t4 3.86095
R66 VDD2.n1 VDD2.t1 3.86095
R67 VDD2.n1 VDD2.t7 3.86095
R68 VDD2.n0 VDD2.t0 3.86095
R69 VDD2.n0 VDD2.t5 3.86095
R70 VDD2 VDD2.n4 0.459552
R71 VP.n3 VP.t5 430.497
R72 VP.n1 VP.t1 403.675
R73 VP.n10 VP.t7 403.675
R74 VP.n11 VP.t6 403.675
R75 VP.n12 VP.t0 403.675
R76 VP.n6 VP.t2 403.675
R77 VP.n5 VP.t3 403.675
R78 VP.n4 VP.t4 403.675
R79 VP.n13 VP.n12 161.3
R80 VP.n7 VP.n6 161.3
R81 VP.n8 VP.n1 161.3
R82 VP.n5 VP.n2 80.6037
R83 VP.n11 VP.n0 80.6037
R84 VP.n10 VP.n9 80.6037
R85 VP.n10 VP.n1 48.2005
R86 VP.n11 VP.n10 48.2005
R87 VP.n12 VP.n11 48.2005
R88 VP.n6 VP.n5 48.2005
R89 VP.n5 VP.n4 48.2005
R90 VP.n3 VP.n2 45.2318
R91 VP.n8 VP.n7 38.8641
R92 VP.n4 VP.n3 13.3799
R93 VP.n9 VP.n0 0.380177
R94 VP.n7 VP.n2 0.285035
R95 VP.n9 VP.n8 0.285035
R96 VP.n13 VP.n0 0.285035
R97 VP VP.n13 0.0516364
R98 VDD1 VDD1.n0 80.2189
R99 VDD1.n3 VDD1.n2 80.1053
R100 VDD1.n3 VDD1.n1 80.1053
R101 VDD1.n5 VDD1.n4 79.7598
R102 VDD1.n5 VDD1.n3 35.1647
R103 VDD1.n4 VDD1.t4 3.86095
R104 VDD1.n4 VDD1.t5 3.86095
R105 VDD1.n0 VDD1.t2 3.86095
R106 VDD1.n0 VDD1.t3 3.86095
R107 VDD1.n2 VDD1.t1 3.86095
R108 VDD1.n2 VDD1.t7 3.86095
R109 VDD1.n1 VDD1.t6 3.86095
R110 VDD1.n1 VDD1.t0 3.86095
R111 VDD1 VDD1.n5 0.343172
R112 B.n337 B.n336 585
R113 B.n338 B.n53 585
R114 B.n340 B.n339 585
R115 B.n341 B.n52 585
R116 B.n343 B.n342 585
R117 B.n344 B.n51 585
R118 B.n346 B.n345 585
R119 B.n347 B.n50 585
R120 B.n349 B.n348 585
R121 B.n350 B.n49 585
R122 B.n352 B.n351 585
R123 B.n353 B.n48 585
R124 B.n355 B.n354 585
R125 B.n356 B.n47 585
R126 B.n358 B.n357 585
R127 B.n359 B.n46 585
R128 B.n361 B.n360 585
R129 B.n362 B.n45 585
R130 B.n364 B.n363 585
R131 B.n365 B.n44 585
R132 B.n367 B.n366 585
R133 B.n368 B.n43 585
R134 B.n370 B.n369 585
R135 B.n371 B.n42 585
R136 B.n373 B.n372 585
R137 B.n374 B.n41 585
R138 B.n376 B.n375 585
R139 B.n377 B.n40 585
R140 B.n379 B.n378 585
R141 B.n380 B.n39 585
R142 B.n382 B.n381 585
R143 B.n384 B.n36 585
R144 B.n386 B.n385 585
R145 B.n387 B.n35 585
R146 B.n389 B.n388 585
R147 B.n390 B.n34 585
R148 B.n392 B.n391 585
R149 B.n393 B.n33 585
R150 B.n395 B.n394 585
R151 B.n396 B.n29 585
R152 B.n398 B.n397 585
R153 B.n399 B.n28 585
R154 B.n401 B.n400 585
R155 B.n402 B.n27 585
R156 B.n404 B.n403 585
R157 B.n405 B.n26 585
R158 B.n407 B.n406 585
R159 B.n408 B.n25 585
R160 B.n410 B.n409 585
R161 B.n411 B.n24 585
R162 B.n413 B.n412 585
R163 B.n414 B.n23 585
R164 B.n416 B.n415 585
R165 B.n417 B.n22 585
R166 B.n419 B.n418 585
R167 B.n420 B.n21 585
R168 B.n422 B.n421 585
R169 B.n423 B.n20 585
R170 B.n425 B.n424 585
R171 B.n426 B.n19 585
R172 B.n428 B.n427 585
R173 B.n429 B.n18 585
R174 B.n431 B.n430 585
R175 B.n432 B.n17 585
R176 B.n434 B.n433 585
R177 B.n435 B.n16 585
R178 B.n437 B.n436 585
R179 B.n438 B.n15 585
R180 B.n440 B.n439 585
R181 B.n441 B.n14 585
R182 B.n443 B.n442 585
R183 B.n444 B.n13 585
R184 B.n335 B.n54 585
R185 B.n334 B.n333 585
R186 B.n332 B.n55 585
R187 B.n331 B.n330 585
R188 B.n329 B.n56 585
R189 B.n328 B.n327 585
R190 B.n326 B.n57 585
R191 B.n325 B.n324 585
R192 B.n323 B.n58 585
R193 B.n322 B.n321 585
R194 B.n320 B.n59 585
R195 B.n319 B.n318 585
R196 B.n317 B.n60 585
R197 B.n316 B.n315 585
R198 B.n314 B.n61 585
R199 B.n313 B.n312 585
R200 B.n311 B.n62 585
R201 B.n310 B.n309 585
R202 B.n308 B.n63 585
R203 B.n307 B.n306 585
R204 B.n305 B.n64 585
R205 B.n304 B.n303 585
R206 B.n302 B.n65 585
R207 B.n301 B.n300 585
R208 B.n299 B.n66 585
R209 B.n298 B.n297 585
R210 B.n296 B.n67 585
R211 B.n295 B.n294 585
R212 B.n293 B.n68 585
R213 B.n292 B.n291 585
R214 B.n290 B.n69 585
R215 B.n289 B.n288 585
R216 B.n287 B.n70 585
R217 B.n286 B.n285 585
R218 B.n284 B.n71 585
R219 B.n283 B.n282 585
R220 B.n281 B.n72 585
R221 B.n280 B.n279 585
R222 B.n278 B.n73 585
R223 B.n277 B.n276 585
R224 B.n275 B.n74 585
R225 B.n274 B.n273 585
R226 B.n272 B.n75 585
R227 B.n271 B.n270 585
R228 B.n269 B.n76 585
R229 B.n160 B.n159 585
R230 B.n161 B.n116 585
R231 B.n163 B.n162 585
R232 B.n164 B.n115 585
R233 B.n166 B.n165 585
R234 B.n167 B.n114 585
R235 B.n169 B.n168 585
R236 B.n170 B.n113 585
R237 B.n172 B.n171 585
R238 B.n173 B.n112 585
R239 B.n175 B.n174 585
R240 B.n176 B.n111 585
R241 B.n178 B.n177 585
R242 B.n179 B.n110 585
R243 B.n181 B.n180 585
R244 B.n182 B.n109 585
R245 B.n184 B.n183 585
R246 B.n185 B.n108 585
R247 B.n187 B.n186 585
R248 B.n188 B.n107 585
R249 B.n190 B.n189 585
R250 B.n191 B.n106 585
R251 B.n193 B.n192 585
R252 B.n194 B.n105 585
R253 B.n196 B.n195 585
R254 B.n197 B.n104 585
R255 B.n199 B.n198 585
R256 B.n200 B.n103 585
R257 B.n202 B.n201 585
R258 B.n203 B.n102 585
R259 B.n205 B.n204 585
R260 B.n207 B.n206 585
R261 B.n208 B.n98 585
R262 B.n210 B.n209 585
R263 B.n211 B.n97 585
R264 B.n213 B.n212 585
R265 B.n214 B.n96 585
R266 B.n216 B.n215 585
R267 B.n217 B.n95 585
R268 B.n219 B.n218 585
R269 B.n220 B.n92 585
R270 B.n223 B.n222 585
R271 B.n224 B.n91 585
R272 B.n226 B.n225 585
R273 B.n227 B.n90 585
R274 B.n229 B.n228 585
R275 B.n230 B.n89 585
R276 B.n232 B.n231 585
R277 B.n233 B.n88 585
R278 B.n235 B.n234 585
R279 B.n236 B.n87 585
R280 B.n238 B.n237 585
R281 B.n239 B.n86 585
R282 B.n241 B.n240 585
R283 B.n242 B.n85 585
R284 B.n244 B.n243 585
R285 B.n245 B.n84 585
R286 B.n247 B.n246 585
R287 B.n248 B.n83 585
R288 B.n250 B.n249 585
R289 B.n251 B.n82 585
R290 B.n253 B.n252 585
R291 B.n254 B.n81 585
R292 B.n256 B.n255 585
R293 B.n257 B.n80 585
R294 B.n259 B.n258 585
R295 B.n260 B.n79 585
R296 B.n262 B.n261 585
R297 B.n263 B.n78 585
R298 B.n265 B.n264 585
R299 B.n266 B.n77 585
R300 B.n268 B.n267 585
R301 B.n158 B.n117 585
R302 B.n157 B.n156 585
R303 B.n155 B.n118 585
R304 B.n154 B.n153 585
R305 B.n152 B.n119 585
R306 B.n151 B.n150 585
R307 B.n149 B.n120 585
R308 B.n148 B.n147 585
R309 B.n146 B.n121 585
R310 B.n145 B.n144 585
R311 B.n143 B.n122 585
R312 B.n142 B.n141 585
R313 B.n140 B.n123 585
R314 B.n139 B.n138 585
R315 B.n137 B.n124 585
R316 B.n136 B.n135 585
R317 B.n134 B.n125 585
R318 B.n133 B.n132 585
R319 B.n131 B.n126 585
R320 B.n130 B.n129 585
R321 B.n128 B.n127 585
R322 B.n2 B.n0 585
R323 B.n477 B.n1 585
R324 B.n476 B.n475 585
R325 B.n474 B.n3 585
R326 B.n473 B.n472 585
R327 B.n471 B.n4 585
R328 B.n470 B.n469 585
R329 B.n468 B.n5 585
R330 B.n467 B.n466 585
R331 B.n465 B.n6 585
R332 B.n464 B.n463 585
R333 B.n462 B.n7 585
R334 B.n461 B.n460 585
R335 B.n459 B.n8 585
R336 B.n458 B.n457 585
R337 B.n456 B.n9 585
R338 B.n455 B.n454 585
R339 B.n453 B.n10 585
R340 B.n452 B.n451 585
R341 B.n450 B.n11 585
R342 B.n449 B.n448 585
R343 B.n447 B.n12 585
R344 B.n446 B.n445 585
R345 B.n479 B.n478 585
R346 B.n93 B.t6 542.604
R347 B.n99 B.t0 542.604
R348 B.n30 B.t3 542.604
R349 B.n37 B.t9 542.604
R350 B.n159 B.n158 444.452
R351 B.n446 B.n13 444.452
R352 B.n267 B.n76 444.452
R353 B.n337 B.n54 444.452
R354 B.n158 B.n157 163.367
R355 B.n157 B.n118 163.367
R356 B.n153 B.n118 163.367
R357 B.n153 B.n152 163.367
R358 B.n152 B.n151 163.367
R359 B.n151 B.n120 163.367
R360 B.n147 B.n120 163.367
R361 B.n147 B.n146 163.367
R362 B.n146 B.n145 163.367
R363 B.n145 B.n122 163.367
R364 B.n141 B.n122 163.367
R365 B.n141 B.n140 163.367
R366 B.n140 B.n139 163.367
R367 B.n139 B.n124 163.367
R368 B.n135 B.n124 163.367
R369 B.n135 B.n134 163.367
R370 B.n134 B.n133 163.367
R371 B.n133 B.n126 163.367
R372 B.n129 B.n126 163.367
R373 B.n129 B.n128 163.367
R374 B.n128 B.n2 163.367
R375 B.n478 B.n2 163.367
R376 B.n478 B.n477 163.367
R377 B.n477 B.n476 163.367
R378 B.n476 B.n3 163.367
R379 B.n472 B.n3 163.367
R380 B.n472 B.n471 163.367
R381 B.n471 B.n470 163.367
R382 B.n470 B.n5 163.367
R383 B.n466 B.n5 163.367
R384 B.n466 B.n465 163.367
R385 B.n465 B.n464 163.367
R386 B.n464 B.n7 163.367
R387 B.n460 B.n7 163.367
R388 B.n460 B.n459 163.367
R389 B.n459 B.n458 163.367
R390 B.n458 B.n9 163.367
R391 B.n454 B.n9 163.367
R392 B.n454 B.n453 163.367
R393 B.n453 B.n452 163.367
R394 B.n452 B.n11 163.367
R395 B.n448 B.n11 163.367
R396 B.n448 B.n447 163.367
R397 B.n447 B.n446 163.367
R398 B.n159 B.n116 163.367
R399 B.n163 B.n116 163.367
R400 B.n164 B.n163 163.367
R401 B.n165 B.n164 163.367
R402 B.n165 B.n114 163.367
R403 B.n169 B.n114 163.367
R404 B.n170 B.n169 163.367
R405 B.n171 B.n170 163.367
R406 B.n171 B.n112 163.367
R407 B.n175 B.n112 163.367
R408 B.n176 B.n175 163.367
R409 B.n177 B.n176 163.367
R410 B.n177 B.n110 163.367
R411 B.n181 B.n110 163.367
R412 B.n182 B.n181 163.367
R413 B.n183 B.n182 163.367
R414 B.n183 B.n108 163.367
R415 B.n187 B.n108 163.367
R416 B.n188 B.n187 163.367
R417 B.n189 B.n188 163.367
R418 B.n189 B.n106 163.367
R419 B.n193 B.n106 163.367
R420 B.n194 B.n193 163.367
R421 B.n195 B.n194 163.367
R422 B.n195 B.n104 163.367
R423 B.n199 B.n104 163.367
R424 B.n200 B.n199 163.367
R425 B.n201 B.n200 163.367
R426 B.n201 B.n102 163.367
R427 B.n205 B.n102 163.367
R428 B.n206 B.n205 163.367
R429 B.n206 B.n98 163.367
R430 B.n210 B.n98 163.367
R431 B.n211 B.n210 163.367
R432 B.n212 B.n211 163.367
R433 B.n212 B.n96 163.367
R434 B.n216 B.n96 163.367
R435 B.n217 B.n216 163.367
R436 B.n218 B.n217 163.367
R437 B.n218 B.n92 163.367
R438 B.n223 B.n92 163.367
R439 B.n224 B.n223 163.367
R440 B.n225 B.n224 163.367
R441 B.n225 B.n90 163.367
R442 B.n229 B.n90 163.367
R443 B.n230 B.n229 163.367
R444 B.n231 B.n230 163.367
R445 B.n231 B.n88 163.367
R446 B.n235 B.n88 163.367
R447 B.n236 B.n235 163.367
R448 B.n237 B.n236 163.367
R449 B.n237 B.n86 163.367
R450 B.n241 B.n86 163.367
R451 B.n242 B.n241 163.367
R452 B.n243 B.n242 163.367
R453 B.n243 B.n84 163.367
R454 B.n247 B.n84 163.367
R455 B.n248 B.n247 163.367
R456 B.n249 B.n248 163.367
R457 B.n249 B.n82 163.367
R458 B.n253 B.n82 163.367
R459 B.n254 B.n253 163.367
R460 B.n255 B.n254 163.367
R461 B.n255 B.n80 163.367
R462 B.n259 B.n80 163.367
R463 B.n260 B.n259 163.367
R464 B.n261 B.n260 163.367
R465 B.n261 B.n78 163.367
R466 B.n265 B.n78 163.367
R467 B.n266 B.n265 163.367
R468 B.n267 B.n266 163.367
R469 B.n271 B.n76 163.367
R470 B.n272 B.n271 163.367
R471 B.n273 B.n272 163.367
R472 B.n273 B.n74 163.367
R473 B.n277 B.n74 163.367
R474 B.n278 B.n277 163.367
R475 B.n279 B.n278 163.367
R476 B.n279 B.n72 163.367
R477 B.n283 B.n72 163.367
R478 B.n284 B.n283 163.367
R479 B.n285 B.n284 163.367
R480 B.n285 B.n70 163.367
R481 B.n289 B.n70 163.367
R482 B.n290 B.n289 163.367
R483 B.n291 B.n290 163.367
R484 B.n291 B.n68 163.367
R485 B.n295 B.n68 163.367
R486 B.n296 B.n295 163.367
R487 B.n297 B.n296 163.367
R488 B.n297 B.n66 163.367
R489 B.n301 B.n66 163.367
R490 B.n302 B.n301 163.367
R491 B.n303 B.n302 163.367
R492 B.n303 B.n64 163.367
R493 B.n307 B.n64 163.367
R494 B.n308 B.n307 163.367
R495 B.n309 B.n308 163.367
R496 B.n309 B.n62 163.367
R497 B.n313 B.n62 163.367
R498 B.n314 B.n313 163.367
R499 B.n315 B.n314 163.367
R500 B.n315 B.n60 163.367
R501 B.n319 B.n60 163.367
R502 B.n320 B.n319 163.367
R503 B.n321 B.n320 163.367
R504 B.n321 B.n58 163.367
R505 B.n325 B.n58 163.367
R506 B.n326 B.n325 163.367
R507 B.n327 B.n326 163.367
R508 B.n327 B.n56 163.367
R509 B.n331 B.n56 163.367
R510 B.n332 B.n331 163.367
R511 B.n333 B.n332 163.367
R512 B.n333 B.n54 163.367
R513 B.n442 B.n13 163.367
R514 B.n442 B.n441 163.367
R515 B.n441 B.n440 163.367
R516 B.n440 B.n15 163.367
R517 B.n436 B.n15 163.367
R518 B.n436 B.n435 163.367
R519 B.n435 B.n434 163.367
R520 B.n434 B.n17 163.367
R521 B.n430 B.n17 163.367
R522 B.n430 B.n429 163.367
R523 B.n429 B.n428 163.367
R524 B.n428 B.n19 163.367
R525 B.n424 B.n19 163.367
R526 B.n424 B.n423 163.367
R527 B.n423 B.n422 163.367
R528 B.n422 B.n21 163.367
R529 B.n418 B.n21 163.367
R530 B.n418 B.n417 163.367
R531 B.n417 B.n416 163.367
R532 B.n416 B.n23 163.367
R533 B.n412 B.n23 163.367
R534 B.n412 B.n411 163.367
R535 B.n411 B.n410 163.367
R536 B.n410 B.n25 163.367
R537 B.n406 B.n25 163.367
R538 B.n406 B.n405 163.367
R539 B.n405 B.n404 163.367
R540 B.n404 B.n27 163.367
R541 B.n400 B.n27 163.367
R542 B.n400 B.n399 163.367
R543 B.n399 B.n398 163.367
R544 B.n398 B.n29 163.367
R545 B.n394 B.n29 163.367
R546 B.n394 B.n393 163.367
R547 B.n393 B.n392 163.367
R548 B.n392 B.n34 163.367
R549 B.n388 B.n34 163.367
R550 B.n388 B.n387 163.367
R551 B.n387 B.n386 163.367
R552 B.n386 B.n36 163.367
R553 B.n381 B.n36 163.367
R554 B.n381 B.n380 163.367
R555 B.n380 B.n379 163.367
R556 B.n379 B.n40 163.367
R557 B.n375 B.n40 163.367
R558 B.n375 B.n374 163.367
R559 B.n374 B.n373 163.367
R560 B.n373 B.n42 163.367
R561 B.n369 B.n42 163.367
R562 B.n369 B.n368 163.367
R563 B.n368 B.n367 163.367
R564 B.n367 B.n44 163.367
R565 B.n363 B.n44 163.367
R566 B.n363 B.n362 163.367
R567 B.n362 B.n361 163.367
R568 B.n361 B.n46 163.367
R569 B.n357 B.n46 163.367
R570 B.n357 B.n356 163.367
R571 B.n356 B.n355 163.367
R572 B.n355 B.n48 163.367
R573 B.n351 B.n48 163.367
R574 B.n351 B.n350 163.367
R575 B.n350 B.n349 163.367
R576 B.n349 B.n50 163.367
R577 B.n345 B.n50 163.367
R578 B.n345 B.n344 163.367
R579 B.n344 B.n343 163.367
R580 B.n343 B.n52 163.367
R581 B.n339 B.n52 163.367
R582 B.n339 B.n338 163.367
R583 B.n338 B.n337 163.367
R584 B.n93 B.t8 131.5
R585 B.n37 B.t10 131.5
R586 B.n99 B.t2 131.492
R587 B.n30 B.t4 131.492
R588 B.n94 B.t7 113.465
R589 B.n38 B.t11 113.465
R590 B.n100 B.t1 113.456
R591 B.n31 B.t5 113.456
R592 B.n221 B.n94 59.5399
R593 B.n101 B.n100 59.5399
R594 B.n32 B.n31 59.5399
R595 B.n383 B.n38 59.5399
R596 B.n445 B.n444 28.8785
R597 B.n269 B.n268 28.8785
R598 B.n160 B.n117 28.8785
R599 B.n336 B.n335 28.8785
R600 B B.n479 18.0485
R601 B.n94 B.n93 18.0369
R602 B.n100 B.n99 18.0369
R603 B.n31 B.n30 18.0369
R604 B.n38 B.n37 18.0369
R605 B.n444 B.n443 10.6151
R606 B.n443 B.n14 10.6151
R607 B.n439 B.n14 10.6151
R608 B.n439 B.n438 10.6151
R609 B.n438 B.n437 10.6151
R610 B.n437 B.n16 10.6151
R611 B.n433 B.n16 10.6151
R612 B.n433 B.n432 10.6151
R613 B.n432 B.n431 10.6151
R614 B.n431 B.n18 10.6151
R615 B.n427 B.n18 10.6151
R616 B.n427 B.n426 10.6151
R617 B.n426 B.n425 10.6151
R618 B.n425 B.n20 10.6151
R619 B.n421 B.n20 10.6151
R620 B.n421 B.n420 10.6151
R621 B.n420 B.n419 10.6151
R622 B.n419 B.n22 10.6151
R623 B.n415 B.n22 10.6151
R624 B.n415 B.n414 10.6151
R625 B.n414 B.n413 10.6151
R626 B.n413 B.n24 10.6151
R627 B.n409 B.n24 10.6151
R628 B.n409 B.n408 10.6151
R629 B.n408 B.n407 10.6151
R630 B.n407 B.n26 10.6151
R631 B.n403 B.n26 10.6151
R632 B.n403 B.n402 10.6151
R633 B.n402 B.n401 10.6151
R634 B.n401 B.n28 10.6151
R635 B.n397 B.n396 10.6151
R636 B.n396 B.n395 10.6151
R637 B.n395 B.n33 10.6151
R638 B.n391 B.n33 10.6151
R639 B.n391 B.n390 10.6151
R640 B.n390 B.n389 10.6151
R641 B.n389 B.n35 10.6151
R642 B.n385 B.n35 10.6151
R643 B.n385 B.n384 10.6151
R644 B.n382 B.n39 10.6151
R645 B.n378 B.n39 10.6151
R646 B.n378 B.n377 10.6151
R647 B.n377 B.n376 10.6151
R648 B.n376 B.n41 10.6151
R649 B.n372 B.n41 10.6151
R650 B.n372 B.n371 10.6151
R651 B.n371 B.n370 10.6151
R652 B.n370 B.n43 10.6151
R653 B.n366 B.n43 10.6151
R654 B.n366 B.n365 10.6151
R655 B.n365 B.n364 10.6151
R656 B.n364 B.n45 10.6151
R657 B.n360 B.n45 10.6151
R658 B.n360 B.n359 10.6151
R659 B.n359 B.n358 10.6151
R660 B.n358 B.n47 10.6151
R661 B.n354 B.n47 10.6151
R662 B.n354 B.n353 10.6151
R663 B.n353 B.n352 10.6151
R664 B.n352 B.n49 10.6151
R665 B.n348 B.n49 10.6151
R666 B.n348 B.n347 10.6151
R667 B.n347 B.n346 10.6151
R668 B.n346 B.n51 10.6151
R669 B.n342 B.n51 10.6151
R670 B.n342 B.n341 10.6151
R671 B.n341 B.n340 10.6151
R672 B.n340 B.n53 10.6151
R673 B.n336 B.n53 10.6151
R674 B.n270 B.n269 10.6151
R675 B.n270 B.n75 10.6151
R676 B.n274 B.n75 10.6151
R677 B.n275 B.n274 10.6151
R678 B.n276 B.n275 10.6151
R679 B.n276 B.n73 10.6151
R680 B.n280 B.n73 10.6151
R681 B.n281 B.n280 10.6151
R682 B.n282 B.n281 10.6151
R683 B.n282 B.n71 10.6151
R684 B.n286 B.n71 10.6151
R685 B.n287 B.n286 10.6151
R686 B.n288 B.n287 10.6151
R687 B.n288 B.n69 10.6151
R688 B.n292 B.n69 10.6151
R689 B.n293 B.n292 10.6151
R690 B.n294 B.n293 10.6151
R691 B.n294 B.n67 10.6151
R692 B.n298 B.n67 10.6151
R693 B.n299 B.n298 10.6151
R694 B.n300 B.n299 10.6151
R695 B.n300 B.n65 10.6151
R696 B.n304 B.n65 10.6151
R697 B.n305 B.n304 10.6151
R698 B.n306 B.n305 10.6151
R699 B.n306 B.n63 10.6151
R700 B.n310 B.n63 10.6151
R701 B.n311 B.n310 10.6151
R702 B.n312 B.n311 10.6151
R703 B.n312 B.n61 10.6151
R704 B.n316 B.n61 10.6151
R705 B.n317 B.n316 10.6151
R706 B.n318 B.n317 10.6151
R707 B.n318 B.n59 10.6151
R708 B.n322 B.n59 10.6151
R709 B.n323 B.n322 10.6151
R710 B.n324 B.n323 10.6151
R711 B.n324 B.n57 10.6151
R712 B.n328 B.n57 10.6151
R713 B.n329 B.n328 10.6151
R714 B.n330 B.n329 10.6151
R715 B.n330 B.n55 10.6151
R716 B.n334 B.n55 10.6151
R717 B.n335 B.n334 10.6151
R718 B.n161 B.n160 10.6151
R719 B.n162 B.n161 10.6151
R720 B.n162 B.n115 10.6151
R721 B.n166 B.n115 10.6151
R722 B.n167 B.n166 10.6151
R723 B.n168 B.n167 10.6151
R724 B.n168 B.n113 10.6151
R725 B.n172 B.n113 10.6151
R726 B.n173 B.n172 10.6151
R727 B.n174 B.n173 10.6151
R728 B.n174 B.n111 10.6151
R729 B.n178 B.n111 10.6151
R730 B.n179 B.n178 10.6151
R731 B.n180 B.n179 10.6151
R732 B.n180 B.n109 10.6151
R733 B.n184 B.n109 10.6151
R734 B.n185 B.n184 10.6151
R735 B.n186 B.n185 10.6151
R736 B.n186 B.n107 10.6151
R737 B.n190 B.n107 10.6151
R738 B.n191 B.n190 10.6151
R739 B.n192 B.n191 10.6151
R740 B.n192 B.n105 10.6151
R741 B.n196 B.n105 10.6151
R742 B.n197 B.n196 10.6151
R743 B.n198 B.n197 10.6151
R744 B.n198 B.n103 10.6151
R745 B.n202 B.n103 10.6151
R746 B.n203 B.n202 10.6151
R747 B.n204 B.n203 10.6151
R748 B.n208 B.n207 10.6151
R749 B.n209 B.n208 10.6151
R750 B.n209 B.n97 10.6151
R751 B.n213 B.n97 10.6151
R752 B.n214 B.n213 10.6151
R753 B.n215 B.n214 10.6151
R754 B.n215 B.n95 10.6151
R755 B.n219 B.n95 10.6151
R756 B.n220 B.n219 10.6151
R757 B.n222 B.n91 10.6151
R758 B.n226 B.n91 10.6151
R759 B.n227 B.n226 10.6151
R760 B.n228 B.n227 10.6151
R761 B.n228 B.n89 10.6151
R762 B.n232 B.n89 10.6151
R763 B.n233 B.n232 10.6151
R764 B.n234 B.n233 10.6151
R765 B.n234 B.n87 10.6151
R766 B.n238 B.n87 10.6151
R767 B.n239 B.n238 10.6151
R768 B.n240 B.n239 10.6151
R769 B.n240 B.n85 10.6151
R770 B.n244 B.n85 10.6151
R771 B.n245 B.n244 10.6151
R772 B.n246 B.n245 10.6151
R773 B.n246 B.n83 10.6151
R774 B.n250 B.n83 10.6151
R775 B.n251 B.n250 10.6151
R776 B.n252 B.n251 10.6151
R777 B.n252 B.n81 10.6151
R778 B.n256 B.n81 10.6151
R779 B.n257 B.n256 10.6151
R780 B.n258 B.n257 10.6151
R781 B.n258 B.n79 10.6151
R782 B.n262 B.n79 10.6151
R783 B.n263 B.n262 10.6151
R784 B.n264 B.n263 10.6151
R785 B.n264 B.n77 10.6151
R786 B.n268 B.n77 10.6151
R787 B.n156 B.n117 10.6151
R788 B.n156 B.n155 10.6151
R789 B.n155 B.n154 10.6151
R790 B.n154 B.n119 10.6151
R791 B.n150 B.n119 10.6151
R792 B.n150 B.n149 10.6151
R793 B.n149 B.n148 10.6151
R794 B.n148 B.n121 10.6151
R795 B.n144 B.n121 10.6151
R796 B.n144 B.n143 10.6151
R797 B.n143 B.n142 10.6151
R798 B.n142 B.n123 10.6151
R799 B.n138 B.n123 10.6151
R800 B.n138 B.n137 10.6151
R801 B.n137 B.n136 10.6151
R802 B.n136 B.n125 10.6151
R803 B.n132 B.n125 10.6151
R804 B.n132 B.n131 10.6151
R805 B.n131 B.n130 10.6151
R806 B.n130 B.n127 10.6151
R807 B.n127 B.n0 10.6151
R808 B.n475 B.n1 10.6151
R809 B.n475 B.n474 10.6151
R810 B.n474 B.n473 10.6151
R811 B.n473 B.n4 10.6151
R812 B.n469 B.n4 10.6151
R813 B.n469 B.n468 10.6151
R814 B.n468 B.n467 10.6151
R815 B.n467 B.n6 10.6151
R816 B.n463 B.n6 10.6151
R817 B.n463 B.n462 10.6151
R818 B.n462 B.n461 10.6151
R819 B.n461 B.n8 10.6151
R820 B.n457 B.n8 10.6151
R821 B.n457 B.n456 10.6151
R822 B.n456 B.n455 10.6151
R823 B.n455 B.n10 10.6151
R824 B.n451 B.n10 10.6151
R825 B.n451 B.n450 10.6151
R826 B.n450 B.n449 10.6151
R827 B.n449 B.n12 10.6151
R828 B.n445 B.n12 10.6151
R829 B.n32 B.n28 9.36635
R830 B.n383 B.n382 9.36635
R831 B.n204 B.n101 9.36635
R832 B.n222 B.n221 9.36635
R833 B.n479 B.n0 2.81026
R834 B.n479 B.n1 2.81026
R835 B.n397 B.n32 1.24928
R836 B.n384 B.n383 1.24928
R837 B.n207 B.n101 1.24928
R838 B.n221 B.n220 1.24928
C0 VDD2 VN 3.66667f
C1 B w_n1900_n2652# 6.0521f
C2 w_n1900_n2652# VP 3.4727f
C3 VDD2 B 0.976585f
C4 VTAIL VN 3.52547f
C5 VDD2 VP 0.307222f
C6 VTAIL B 2.80883f
C7 B VN 0.71766f
C8 VTAIL VP 3.53957f
C9 VDD1 w_n1900_n2652# 1.16618f
C10 VP VN 4.5501f
C11 VDD2 VDD1 0.777234f
C12 B VP 1.1106f
C13 VDD1 VTAIL 8.940981f
C14 VDD1 VN 0.148484f
C15 VDD1 B 0.943013f
C16 VDD1 VP 3.82502f
C17 VDD2 w_n1900_n2652# 1.19688f
C18 VTAIL w_n1900_n2652# 3.31883f
C19 w_n1900_n2652# VN 3.23193f
C20 VDD2 VTAIL 8.98199f
C21 VDD2 VSUBS 1.224548f
C22 VDD1 VSUBS 1.506897f
C23 VTAIL VSUBS 0.716584f
C24 VN VSUBS 4.33961f
C25 VP VSUBS 1.415875f
C26 B VSUBS 2.465117f
C27 w_n1900_n2652# VSUBS 62.4492f
C28 B.n0 VSUBS 0.00555f
C29 B.n1 VSUBS 0.00555f
C30 B.n2 VSUBS 0.008777f
C31 B.n3 VSUBS 0.008777f
C32 B.n4 VSUBS 0.008777f
C33 B.n5 VSUBS 0.008777f
C34 B.n6 VSUBS 0.008777f
C35 B.n7 VSUBS 0.008777f
C36 B.n8 VSUBS 0.008777f
C37 B.n9 VSUBS 0.008777f
C38 B.n10 VSUBS 0.008777f
C39 B.n11 VSUBS 0.008777f
C40 B.n12 VSUBS 0.008777f
C41 B.n13 VSUBS 0.019446f
C42 B.n14 VSUBS 0.008777f
C43 B.n15 VSUBS 0.008777f
C44 B.n16 VSUBS 0.008777f
C45 B.n17 VSUBS 0.008777f
C46 B.n18 VSUBS 0.008777f
C47 B.n19 VSUBS 0.008777f
C48 B.n20 VSUBS 0.008777f
C49 B.n21 VSUBS 0.008777f
C50 B.n22 VSUBS 0.008777f
C51 B.n23 VSUBS 0.008777f
C52 B.n24 VSUBS 0.008777f
C53 B.n25 VSUBS 0.008777f
C54 B.n26 VSUBS 0.008777f
C55 B.n27 VSUBS 0.008777f
C56 B.n28 VSUBS 0.008261f
C57 B.n29 VSUBS 0.008777f
C58 B.t5 VSUBS 0.32842f
C59 B.t4 VSUBS 0.337574f
C60 B.t3 VSUBS 0.264454f
C61 B.n30 VSUBS 0.127728f
C62 B.n31 VSUBS 0.079254f
C63 B.n32 VSUBS 0.020335f
C64 B.n33 VSUBS 0.008777f
C65 B.n34 VSUBS 0.008777f
C66 B.n35 VSUBS 0.008777f
C67 B.n36 VSUBS 0.008777f
C68 B.t11 VSUBS 0.328417f
C69 B.t10 VSUBS 0.337571f
C70 B.t9 VSUBS 0.264454f
C71 B.n37 VSUBS 0.127731f
C72 B.n38 VSUBS 0.079257f
C73 B.n39 VSUBS 0.008777f
C74 B.n40 VSUBS 0.008777f
C75 B.n41 VSUBS 0.008777f
C76 B.n42 VSUBS 0.008777f
C77 B.n43 VSUBS 0.008777f
C78 B.n44 VSUBS 0.008777f
C79 B.n45 VSUBS 0.008777f
C80 B.n46 VSUBS 0.008777f
C81 B.n47 VSUBS 0.008777f
C82 B.n48 VSUBS 0.008777f
C83 B.n49 VSUBS 0.008777f
C84 B.n50 VSUBS 0.008777f
C85 B.n51 VSUBS 0.008777f
C86 B.n52 VSUBS 0.008777f
C87 B.n53 VSUBS 0.008777f
C88 B.n54 VSUBS 0.018502f
C89 B.n55 VSUBS 0.008777f
C90 B.n56 VSUBS 0.008777f
C91 B.n57 VSUBS 0.008777f
C92 B.n58 VSUBS 0.008777f
C93 B.n59 VSUBS 0.008777f
C94 B.n60 VSUBS 0.008777f
C95 B.n61 VSUBS 0.008777f
C96 B.n62 VSUBS 0.008777f
C97 B.n63 VSUBS 0.008777f
C98 B.n64 VSUBS 0.008777f
C99 B.n65 VSUBS 0.008777f
C100 B.n66 VSUBS 0.008777f
C101 B.n67 VSUBS 0.008777f
C102 B.n68 VSUBS 0.008777f
C103 B.n69 VSUBS 0.008777f
C104 B.n70 VSUBS 0.008777f
C105 B.n71 VSUBS 0.008777f
C106 B.n72 VSUBS 0.008777f
C107 B.n73 VSUBS 0.008777f
C108 B.n74 VSUBS 0.008777f
C109 B.n75 VSUBS 0.008777f
C110 B.n76 VSUBS 0.018502f
C111 B.n77 VSUBS 0.008777f
C112 B.n78 VSUBS 0.008777f
C113 B.n79 VSUBS 0.008777f
C114 B.n80 VSUBS 0.008777f
C115 B.n81 VSUBS 0.008777f
C116 B.n82 VSUBS 0.008777f
C117 B.n83 VSUBS 0.008777f
C118 B.n84 VSUBS 0.008777f
C119 B.n85 VSUBS 0.008777f
C120 B.n86 VSUBS 0.008777f
C121 B.n87 VSUBS 0.008777f
C122 B.n88 VSUBS 0.008777f
C123 B.n89 VSUBS 0.008777f
C124 B.n90 VSUBS 0.008777f
C125 B.n91 VSUBS 0.008777f
C126 B.n92 VSUBS 0.008777f
C127 B.t7 VSUBS 0.328417f
C128 B.t8 VSUBS 0.337571f
C129 B.t6 VSUBS 0.264454f
C130 B.n93 VSUBS 0.127731f
C131 B.n94 VSUBS 0.079257f
C132 B.n95 VSUBS 0.008777f
C133 B.n96 VSUBS 0.008777f
C134 B.n97 VSUBS 0.008777f
C135 B.n98 VSUBS 0.008777f
C136 B.t1 VSUBS 0.32842f
C137 B.t2 VSUBS 0.337574f
C138 B.t0 VSUBS 0.264454f
C139 B.n99 VSUBS 0.127728f
C140 B.n100 VSUBS 0.079254f
C141 B.n101 VSUBS 0.020335f
C142 B.n102 VSUBS 0.008777f
C143 B.n103 VSUBS 0.008777f
C144 B.n104 VSUBS 0.008777f
C145 B.n105 VSUBS 0.008777f
C146 B.n106 VSUBS 0.008777f
C147 B.n107 VSUBS 0.008777f
C148 B.n108 VSUBS 0.008777f
C149 B.n109 VSUBS 0.008777f
C150 B.n110 VSUBS 0.008777f
C151 B.n111 VSUBS 0.008777f
C152 B.n112 VSUBS 0.008777f
C153 B.n113 VSUBS 0.008777f
C154 B.n114 VSUBS 0.008777f
C155 B.n115 VSUBS 0.008777f
C156 B.n116 VSUBS 0.008777f
C157 B.n117 VSUBS 0.018502f
C158 B.n118 VSUBS 0.008777f
C159 B.n119 VSUBS 0.008777f
C160 B.n120 VSUBS 0.008777f
C161 B.n121 VSUBS 0.008777f
C162 B.n122 VSUBS 0.008777f
C163 B.n123 VSUBS 0.008777f
C164 B.n124 VSUBS 0.008777f
C165 B.n125 VSUBS 0.008777f
C166 B.n126 VSUBS 0.008777f
C167 B.n127 VSUBS 0.008777f
C168 B.n128 VSUBS 0.008777f
C169 B.n129 VSUBS 0.008777f
C170 B.n130 VSUBS 0.008777f
C171 B.n131 VSUBS 0.008777f
C172 B.n132 VSUBS 0.008777f
C173 B.n133 VSUBS 0.008777f
C174 B.n134 VSUBS 0.008777f
C175 B.n135 VSUBS 0.008777f
C176 B.n136 VSUBS 0.008777f
C177 B.n137 VSUBS 0.008777f
C178 B.n138 VSUBS 0.008777f
C179 B.n139 VSUBS 0.008777f
C180 B.n140 VSUBS 0.008777f
C181 B.n141 VSUBS 0.008777f
C182 B.n142 VSUBS 0.008777f
C183 B.n143 VSUBS 0.008777f
C184 B.n144 VSUBS 0.008777f
C185 B.n145 VSUBS 0.008777f
C186 B.n146 VSUBS 0.008777f
C187 B.n147 VSUBS 0.008777f
C188 B.n148 VSUBS 0.008777f
C189 B.n149 VSUBS 0.008777f
C190 B.n150 VSUBS 0.008777f
C191 B.n151 VSUBS 0.008777f
C192 B.n152 VSUBS 0.008777f
C193 B.n153 VSUBS 0.008777f
C194 B.n154 VSUBS 0.008777f
C195 B.n155 VSUBS 0.008777f
C196 B.n156 VSUBS 0.008777f
C197 B.n157 VSUBS 0.008777f
C198 B.n158 VSUBS 0.018502f
C199 B.n159 VSUBS 0.019446f
C200 B.n160 VSUBS 0.019446f
C201 B.n161 VSUBS 0.008777f
C202 B.n162 VSUBS 0.008777f
C203 B.n163 VSUBS 0.008777f
C204 B.n164 VSUBS 0.008777f
C205 B.n165 VSUBS 0.008777f
C206 B.n166 VSUBS 0.008777f
C207 B.n167 VSUBS 0.008777f
C208 B.n168 VSUBS 0.008777f
C209 B.n169 VSUBS 0.008777f
C210 B.n170 VSUBS 0.008777f
C211 B.n171 VSUBS 0.008777f
C212 B.n172 VSUBS 0.008777f
C213 B.n173 VSUBS 0.008777f
C214 B.n174 VSUBS 0.008777f
C215 B.n175 VSUBS 0.008777f
C216 B.n176 VSUBS 0.008777f
C217 B.n177 VSUBS 0.008777f
C218 B.n178 VSUBS 0.008777f
C219 B.n179 VSUBS 0.008777f
C220 B.n180 VSUBS 0.008777f
C221 B.n181 VSUBS 0.008777f
C222 B.n182 VSUBS 0.008777f
C223 B.n183 VSUBS 0.008777f
C224 B.n184 VSUBS 0.008777f
C225 B.n185 VSUBS 0.008777f
C226 B.n186 VSUBS 0.008777f
C227 B.n187 VSUBS 0.008777f
C228 B.n188 VSUBS 0.008777f
C229 B.n189 VSUBS 0.008777f
C230 B.n190 VSUBS 0.008777f
C231 B.n191 VSUBS 0.008777f
C232 B.n192 VSUBS 0.008777f
C233 B.n193 VSUBS 0.008777f
C234 B.n194 VSUBS 0.008777f
C235 B.n195 VSUBS 0.008777f
C236 B.n196 VSUBS 0.008777f
C237 B.n197 VSUBS 0.008777f
C238 B.n198 VSUBS 0.008777f
C239 B.n199 VSUBS 0.008777f
C240 B.n200 VSUBS 0.008777f
C241 B.n201 VSUBS 0.008777f
C242 B.n202 VSUBS 0.008777f
C243 B.n203 VSUBS 0.008777f
C244 B.n204 VSUBS 0.008261f
C245 B.n205 VSUBS 0.008777f
C246 B.n206 VSUBS 0.008777f
C247 B.n207 VSUBS 0.004905f
C248 B.n208 VSUBS 0.008777f
C249 B.n209 VSUBS 0.008777f
C250 B.n210 VSUBS 0.008777f
C251 B.n211 VSUBS 0.008777f
C252 B.n212 VSUBS 0.008777f
C253 B.n213 VSUBS 0.008777f
C254 B.n214 VSUBS 0.008777f
C255 B.n215 VSUBS 0.008777f
C256 B.n216 VSUBS 0.008777f
C257 B.n217 VSUBS 0.008777f
C258 B.n218 VSUBS 0.008777f
C259 B.n219 VSUBS 0.008777f
C260 B.n220 VSUBS 0.004905f
C261 B.n221 VSUBS 0.020335f
C262 B.n222 VSUBS 0.008261f
C263 B.n223 VSUBS 0.008777f
C264 B.n224 VSUBS 0.008777f
C265 B.n225 VSUBS 0.008777f
C266 B.n226 VSUBS 0.008777f
C267 B.n227 VSUBS 0.008777f
C268 B.n228 VSUBS 0.008777f
C269 B.n229 VSUBS 0.008777f
C270 B.n230 VSUBS 0.008777f
C271 B.n231 VSUBS 0.008777f
C272 B.n232 VSUBS 0.008777f
C273 B.n233 VSUBS 0.008777f
C274 B.n234 VSUBS 0.008777f
C275 B.n235 VSUBS 0.008777f
C276 B.n236 VSUBS 0.008777f
C277 B.n237 VSUBS 0.008777f
C278 B.n238 VSUBS 0.008777f
C279 B.n239 VSUBS 0.008777f
C280 B.n240 VSUBS 0.008777f
C281 B.n241 VSUBS 0.008777f
C282 B.n242 VSUBS 0.008777f
C283 B.n243 VSUBS 0.008777f
C284 B.n244 VSUBS 0.008777f
C285 B.n245 VSUBS 0.008777f
C286 B.n246 VSUBS 0.008777f
C287 B.n247 VSUBS 0.008777f
C288 B.n248 VSUBS 0.008777f
C289 B.n249 VSUBS 0.008777f
C290 B.n250 VSUBS 0.008777f
C291 B.n251 VSUBS 0.008777f
C292 B.n252 VSUBS 0.008777f
C293 B.n253 VSUBS 0.008777f
C294 B.n254 VSUBS 0.008777f
C295 B.n255 VSUBS 0.008777f
C296 B.n256 VSUBS 0.008777f
C297 B.n257 VSUBS 0.008777f
C298 B.n258 VSUBS 0.008777f
C299 B.n259 VSUBS 0.008777f
C300 B.n260 VSUBS 0.008777f
C301 B.n261 VSUBS 0.008777f
C302 B.n262 VSUBS 0.008777f
C303 B.n263 VSUBS 0.008777f
C304 B.n264 VSUBS 0.008777f
C305 B.n265 VSUBS 0.008777f
C306 B.n266 VSUBS 0.008777f
C307 B.n267 VSUBS 0.019446f
C308 B.n268 VSUBS 0.019446f
C309 B.n269 VSUBS 0.018502f
C310 B.n270 VSUBS 0.008777f
C311 B.n271 VSUBS 0.008777f
C312 B.n272 VSUBS 0.008777f
C313 B.n273 VSUBS 0.008777f
C314 B.n274 VSUBS 0.008777f
C315 B.n275 VSUBS 0.008777f
C316 B.n276 VSUBS 0.008777f
C317 B.n277 VSUBS 0.008777f
C318 B.n278 VSUBS 0.008777f
C319 B.n279 VSUBS 0.008777f
C320 B.n280 VSUBS 0.008777f
C321 B.n281 VSUBS 0.008777f
C322 B.n282 VSUBS 0.008777f
C323 B.n283 VSUBS 0.008777f
C324 B.n284 VSUBS 0.008777f
C325 B.n285 VSUBS 0.008777f
C326 B.n286 VSUBS 0.008777f
C327 B.n287 VSUBS 0.008777f
C328 B.n288 VSUBS 0.008777f
C329 B.n289 VSUBS 0.008777f
C330 B.n290 VSUBS 0.008777f
C331 B.n291 VSUBS 0.008777f
C332 B.n292 VSUBS 0.008777f
C333 B.n293 VSUBS 0.008777f
C334 B.n294 VSUBS 0.008777f
C335 B.n295 VSUBS 0.008777f
C336 B.n296 VSUBS 0.008777f
C337 B.n297 VSUBS 0.008777f
C338 B.n298 VSUBS 0.008777f
C339 B.n299 VSUBS 0.008777f
C340 B.n300 VSUBS 0.008777f
C341 B.n301 VSUBS 0.008777f
C342 B.n302 VSUBS 0.008777f
C343 B.n303 VSUBS 0.008777f
C344 B.n304 VSUBS 0.008777f
C345 B.n305 VSUBS 0.008777f
C346 B.n306 VSUBS 0.008777f
C347 B.n307 VSUBS 0.008777f
C348 B.n308 VSUBS 0.008777f
C349 B.n309 VSUBS 0.008777f
C350 B.n310 VSUBS 0.008777f
C351 B.n311 VSUBS 0.008777f
C352 B.n312 VSUBS 0.008777f
C353 B.n313 VSUBS 0.008777f
C354 B.n314 VSUBS 0.008777f
C355 B.n315 VSUBS 0.008777f
C356 B.n316 VSUBS 0.008777f
C357 B.n317 VSUBS 0.008777f
C358 B.n318 VSUBS 0.008777f
C359 B.n319 VSUBS 0.008777f
C360 B.n320 VSUBS 0.008777f
C361 B.n321 VSUBS 0.008777f
C362 B.n322 VSUBS 0.008777f
C363 B.n323 VSUBS 0.008777f
C364 B.n324 VSUBS 0.008777f
C365 B.n325 VSUBS 0.008777f
C366 B.n326 VSUBS 0.008777f
C367 B.n327 VSUBS 0.008777f
C368 B.n328 VSUBS 0.008777f
C369 B.n329 VSUBS 0.008777f
C370 B.n330 VSUBS 0.008777f
C371 B.n331 VSUBS 0.008777f
C372 B.n332 VSUBS 0.008777f
C373 B.n333 VSUBS 0.008777f
C374 B.n334 VSUBS 0.008777f
C375 B.n335 VSUBS 0.019674f
C376 B.n336 VSUBS 0.018273f
C377 B.n337 VSUBS 0.019446f
C378 B.n338 VSUBS 0.008777f
C379 B.n339 VSUBS 0.008777f
C380 B.n340 VSUBS 0.008777f
C381 B.n341 VSUBS 0.008777f
C382 B.n342 VSUBS 0.008777f
C383 B.n343 VSUBS 0.008777f
C384 B.n344 VSUBS 0.008777f
C385 B.n345 VSUBS 0.008777f
C386 B.n346 VSUBS 0.008777f
C387 B.n347 VSUBS 0.008777f
C388 B.n348 VSUBS 0.008777f
C389 B.n349 VSUBS 0.008777f
C390 B.n350 VSUBS 0.008777f
C391 B.n351 VSUBS 0.008777f
C392 B.n352 VSUBS 0.008777f
C393 B.n353 VSUBS 0.008777f
C394 B.n354 VSUBS 0.008777f
C395 B.n355 VSUBS 0.008777f
C396 B.n356 VSUBS 0.008777f
C397 B.n357 VSUBS 0.008777f
C398 B.n358 VSUBS 0.008777f
C399 B.n359 VSUBS 0.008777f
C400 B.n360 VSUBS 0.008777f
C401 B.n361 VSUBS 0.008777f
C402 B.n362 VSUBS 0.008777f
C403 B.n363 VSUBS 0.008777f
C404 B.n364 VSUBS 0.008777f
C405 B.n365 VSUBS 0.008777f
C406 B.n366 VSUBS 0.008777f
C407 B.n367 VSUBS 0.008777f
C408 B.n368 VSUBS 0.008777f
C409 B.n369 VSUBS 0.008777f
C410 B.n370 VSUBS 0.008777f
C411 B.n371 VSUBS 0.008777f
C412 B.n372 VSUBS 0.008777f
C413 B.n373 VSUBS 0.008777f
C414 B.n374 VSUBS 0.008777f
C415 B.n375 VSUBS 0.008777f
C416 B.n376 VSUBS 0.008777f
C417 B.n377 VSUBS 0.008777f
C418 B.n378 VSUBS 0.008777f
C419 B.n379 VSUBS 0.008777f
C420 B.n380 VSUBS 0.008777f
C421 B.n381 VSUBS 0.008777f
C422 B.n382 VSUBS 0.008261f
C423 B.n383 VSUBS 0.020335f
C424 B.n384 VSUBS 0.004905f
C425 B.n385 VSUBS 0.008777f
C426 B.n386 VSUBS 0.008777f
C427 B.n387 VSUBS 0.008777f
C428 B.n388 VSUBS 0.008777f
C429 B.n389 VSUBS 0.008777f
C430 B.n390 VSUBS 0.008777f
C431 B.n391 VSUBS 0.008777f
C432 B.n392 VSUBS 0.008777f
C433 B.n393 VSUBS 0.008777f
C434 B.n394 VSUBS 0.008777f
C435 B.n395 VSUBS 0.008777f
C436 B.n396 VSUBS 0.008777f
C437 B.n397 VSUBS 0.004905f
C438 B.n398 VSUBS 0.008777f
C439 B.n399 VSUBS 0.008777f
C440 B.n400 VSUBS 0.008777f
C441 B.n401 VSUBS 0.008777f
C442 B.n402 VSUBS 0.008777f
C443 B.n403 VSUBS 0.008777f
C444 B.n404 VSUBS 0.008777f
C445 B.n405 VSUBS 0.008777f
C446 B.n406 VSUBS 0.008777f
C447 B.n407 VSUBS 0.008777f
C448 B.n408 VSUBS 0.008777f
C449 B.n409 VSUBS 0.008777f
C450 B.n410 VSUBS 0.008777f
C451 B.n411 VSUBS 0.008777f
C452 B.n412 VSUBS 0.008777f
C453 B.n413 VSUBS 0.008777f
C454 B.n414 VSUBS 0.008777f
C455 B.n415 VSUBS 0.008777f
C456 B.n416 VSUBS 0.008777f
C457 B.n417 VSUBS 0.008777f
C458 B.n418 VSUBS 0.008777f
C459 B.n419 VSUBS 0.008777f
C460 B.n420 VSUBS 0.008777f
C461 B.n421 VSUBS 0.008777f
C462 B.n422 VSUBS 0.008777f
C463 B.n423 VSUBS 0.008777f
C464 B.n424 VSUBS 0.008777f
C465 B.n425 VSUBS 0.008777f
C466 B.n426 VSUBS 0.008777f
C467 B.n427 VSUBS 0.008777f
C468 B.n428 VSUBS 0.008777f
C469 B.n429 VSUBS 0.008777f
C470 B.n430 VSUBS 0.008777f
C471 B.n431 VSUBS 0.008777f
C472 B.n432 VSUBS 0.008777f
C473 B.n433 VSUBS 0.008777f
C474 B.n434 VSUBS 0.008777f
C475 B.n435 VSUBS 0.008777f
C476 B.n436 VSUBS 0.008777f
C477 B.n437 VSUBS 0.008777f
C478 B.n438 VSUBS 0.008777f
C479 B.n439 VSUBS 0.008777f
C480 B.n440 VSUBS 0.008777f
C481 B.n441 VSUBS 0.008777f
C482 B.n442 VSUBS 0.008777f
C483 B.n443 VSUBS 0.008777f
C484 B.n444 VSUBS 0.019446f
C485 B.n445 VSUBS 0.018502f
C486 B.n446 VSUBS 0.018502f
C487 B.n447 VSUBS 0.008777f
C488 B.n448 VSUBS 0.008777f
C489 B.n449 VSUBS 0.008777f
C490 B.n450 VSUBS 0.008777f
C491 B.n451 VSUBS 0.008777f
C492 B.n452 VSUBS 0.008777f
C493 B.n453 VSUBS 0.008777f
C494 B.n454 VSUBS 0.008777f
C495 B.n455 VSUBS 0.008777f
C496 B.n456 VSUBS 0.008777f
C497 B.n457 VSUBS 0.008777f
C498 B.n458 VSUBS 0.008777f
C499 B.n459 VSUBS 0.008777f
C500 B.n460 VSUBS 0.008777f
C501 B.n461 VSUBS 0.008777f
C502 B.n462 VSUBS 0.008777f
C503 B.n463 VSUBS 0.008777f
C504 B.n464 VSUBS 0.008777f
C505 B.n465 VSUBS 0.008777f
C506 B.n466 VSUBS 0.008777f
C507 B.n467 VSUBS 0.008777f
C508 B.n468 VSUBS 0.008777f
C509 B.n469 VSUBS 0.008777f
C510 B.n470 VSUBS 0.008777f
C511 B.n471 VSUBS 0.008777f
C512 B.n472 VSUBS 0.008777f
C513 B.n473 VSUBS 0.008777f
C514 B.n474 VSUBS 0.008777f
C515 B.n475 VSUBS 0.008777f
C516 B.n476 VSUBS 0.008777f
C517 B.n477 VSUBS 0.008777f
C518 B.n478 VSUBS 0.008777f
C519 B.n479 VSUBS 0.019874f
C520 VDD1.t2 VSUBS 0.184771f
C521 VDD1.t3 VSUBS 0.184771f
C522 VDD1.n0 VSUBS 1.33149f
C523 VDD1.t6 VSUBS 0.184771f
C524 VDD1.t0 VSUBS 0.184771f
C525 VDD1.n1 VSUBS 1.33057f
C526 VDD1.t1 VSUBS 0.184771f
C527 VDD1.t7 VSUBS 0.184771f
C528 VDD1.n2 VSUBS 1.33057f
C529 VDD1.n3 VSUBS 2.71027f
C530 VDD1.t4 VSUBS 0.184771f
C531 VDD1.t5 VSUBS 0.184771f
C532 VDD1.n4 VSUBS 1.32791f
C533 VDD1.n5 VSUBS 2.498f
C534 VP.n0 VSUBS 0.10239f
C535 VP.t1 VSUBS 0.892041f
C536 VP.n1 VSUBS 0.382963f
C537 VP.n2 VSUBS 0.299748f
C538 VP.t2 VSUBS 0.892041f
C539 VP.t3 VSUBS 0.892041f
C540 VP.t4 VSUBS 0.892041f
C541 VP.t5 VSUBS 0.915911f
C542 VP.n3 VSUBS 0.360934f
C543 VP.n4 VSUBS 0.396912f
C544 VP.n5 VSUBS 0.396912f
C545 VP.n6 VSUBS 0.382963f
C546 VP.n7 VSUBS 2.24199f
C547 VP.n8 VSUBS 2.29901f
C548 VP.n9 VSUBS 0.10239f
C549 VP.t7 VSUBS 0.892041f
C550 VP.n10 VSUBS 0.396912f
C551 VP.t6 VSUBS 0.892041f
C552 VP.n11 VSUBS 0.396912f
C553 VP.t0 VSUBS 0.892041f
C554 VP.n12 VSUBS 0.382963f
C555 VP.n13 VSUBS 0.068194f
C556 VDD2.t0 VSUBS 0.186275f
C557 VDD2.t5 VSUBS 0.186275f
C558 VDD2.n0 VSUBS 1.3414f
C559 VDD2.t1 VSUBS 0.186275f
C560 VDD2.t7 VSUBS 0.186275f
C561 VDD2.n1 VSUBS 1.3414f
C562 VDD2.n2 VSUBS 2.67232f
C563 VDD2.t6 VSUBS 0.186275f
C564 VDD2.t4 VSUBS 0.186275f
C565 VDD2.n3 VSUBS 1.33872f
C566 VDD2.n4 VSUBS 2.48546f
C567 VDD2.t2 VSUBS 0.186275f
C568 VDD2.t3 VSUBS 0.186275f
C569 VDD2.n5 VSUBS 1.34137f
C570 VTAIL.t10 VSUBS 0.175102f
C571 VTAIL.t8 VSUBS 0.175102f
C572 VTAIL.n0 VSUBS 1.13424f
C573 VTAIL.n1 VSUBS 0.635992f
C574 VTAIL.t12 VSUBS 1.52894f
C575 VTAIL.n2 VSUBS 0.753752f
C576 VTAIL.t6 VSUBS 1.52894f
C577 VTAIL.n3 VSUBS 0.753752f
C578 VTAIL.t0 VSUBS 0.175102f
C579 VTAIL.t7 VSUBS 0.175102f
C580 VTAIL.n4 VSUBS 1.13424f
C581 VTAIL.n5 VSUBS 0.699041f
C582 VTAIL.t3 VSUBS 1.52894f
C583 VTAIL.n6 VSUBS 1.75488f
C584 VTAIL.t9 VSUBS 1.52895f
C585 VTAIL.n7 VSUBS 1.75488f
C586 VTAIL.t14 VSUBS 0.175102f
C587 VTAIL.t15 VSUBS 0.175102f
C588 VTAIL.n8 VSUBS 1.13425f
C589 VTAIL.n9 VSUBS 0.699035f
C590 VTAIL.t11 VSUBS 1.52895f
C591 VTAIL.n10 VSUBS 0.753745f
C592 VTAIL.t4 VSUBS 1.52895f
C593 VTAIL.n11 VSUBS 0.753745f
C594 VTAIL.t5 VSUBS 0.175102f
C595 VTAIL.t2 VSUBS 0.175102f
C596 VTAIL.n12 VSUBS 1.13425f
C597 VTAIL.n13 VSUBS 0.699035f
C598 VTAIL.t1 VSUBS 1.52895f
C599 VTAIL.n14 VSUBS 1.75487f
C600 VTAIL.t13 VSUBS 1.52894f
C601 VTAIL.n15 VSUBS 1.74995f
C602 VN.n0 VSUBS 0.290334f
C603 VN.t7 VSUBS 0.887143f
C604 VN.n1 VSUBS 0.349597f
C605 VN.t2 VSUBS 0.864023f
C606 VN.n2 VSUBS 0.384446f
C607 VN.t6 VSUBS 0.864023f
C608 VN.n3 VSUBS 0.384446f
C609 VN.t0 VSUBS 0.864023f
C610 VN.n4 VSUBS 0.370934f
C611 VN.n5 VSUBS 0.066052f
C612 VN.n6 VSUBS 0.290334f
C613 VN.t5 VSUBS 0.864023f
C614 VN.t4 VSUBS 0.887143f
C615 VN.n7 VSUBS 0.349597f
C616 VN.n8 VSUBS 0.384446f
C617 VN.t3 VSUBS 0.864023f
C618 VN.n9 VSUBS 0.384446f
C619 VN.t1 VSUBS 0.864023f
C620 VN.n10 VSUBS 0.370934f
C621 VN.n11 VSUBS 2.21085f
.ends

