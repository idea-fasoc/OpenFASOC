* NGSPICE file created from diff_pair_sample_0866.ext - technology: sky130A

.subckt diff_pair_sample_0866 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t9 VN.t0 VTAIL.t6 B.t23 sky130_fd_pr__nfet_01v8 ad=3.14655 pd=19.4 as=3.14655 ps=19.4 w=19.07 l=3.94
X1 VDD1.t9 VP.t0 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=3.14655 pd=19.4 as=3.14655 ps=19.4 w=19.07 l=3.94
X2 VDD1.t8 VP.t1 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=7.4373 pd=38.92 as=3.14655 ps=19.4 w=19.07 l=3.94
X3 VTAIL.t9 VN.t1 VDD2.t8 B.t22 sky130_fd_pr__nfet_01v8 ad=3.14655 pd=19.4 as=3.14655 ps=19.4 w=19.07 l=3.94
X4 VDD2.t7 VN.t2 VTAIL.t10 B.t4 sky130_fd_pr__nfet_01v8 ad=3.14655 pd=19.4 as=3.14655 ps=19.4 w=19.07 l=3.94
X5 VDD1.t7 VP.t2 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=7.4373 pd=38.92 as=3.14655 ps=19.4 w=19.07 l=3.94
X6 B.t19 B.t17 B.t18 B.t7 sky130_fd_pr__nfet_01v8 ad=7.4373 pd=38.92 as=0 ps=0 w=19.07 l=3.94
X7 VDD1.t6 VP.t3 VTAIL.t17 B.t23 sky130_fd_pr__nfet_01v8 ad=3.14655 pd=19.4 as=3.14655 ps=19.4 w=19.07 l=3.94
X8 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=7.4373 pd=38.92 as=0 ps=0 w=19.07 l=3.94
X9 VDD2.t6 VN.t3 VTAIL.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=7.4373 pd=38.92 as=3.14655 ps=19.4 w=19.07 l=3.94
X10 VTAIL.t19 VP.t4 VDD1.t5 B.t22 sky130_fd_pr__nfet_01v8 ad=3.14655 pd=19.4 as=3.14655 ps=19.4 w=19.07 l=3.94
X11 VTAIL.t12 VN.t4 VDD2.t5 B.t21 sky130_fd_pr__nfet_01v8 ad=3.14655 pd=19.4 as=3.14655 ps=19.4 w=19.07 l=3.94
X12 VTAIL.t1 VP.t5 VDD1.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=3.14655 pd=19.4 as=3.14655 ps=19.4 w=19.07 l=3.94
X13 VDD2.t4 VN.t5 VTAIL.t15 B.t20 sky130_fd_pr__nfet_01v8 ad=3.14655 pd=19.4 as=7.4373 ps=38.92 w=19.07 l=3.94
X14 VTAIL.t13 VN.t6 VDD2.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=3.14655 pd=19.4 as=3.14655 ps=19.4 w=19.07 l=3.94
X15 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=7.4373 pd=38.92 as=0 ps=0 w=19.07 l=3.94
X16 VDD2.t2 VN.t7 VTAIL.t7 B.t0 sky130_fd_pr__nfet_01v8 ad=3.14655 pd=19.4 as=7.4373 ps=38.92 w=19.07 l=3.94
X17 VDD1.t3 VP.t6 VTAIL.t16 B.t20 sky130_fd_pr__nfet_01v8 ad=3.14655 pd=19.4 as=7.4373 ps=38.92 w=19.07 l=3.94
X18 VTAIL.t18 VP.t7 VDD1.t2 B.t21 sky130_fd_pr__nfet_01v8 ad=3.14655 pd=19.4 as=3.14655 ps=19.4 w=19.07 l=3.94
X19 VDD1.t1 VP.t8 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=3.14655 pd=19.4 as=7.4373 ps=38.92 w=19.07 l=3.94
X20 VDD2.t1 VN.t8 VTAIL.t8 B.t2 sky130_fd_pr__nfet_01v8 ad=7.4373 pd=38.92 as=3.14655 ps=19.4 w=19.07 l=3.94
X21 VTAIL.t5 VP.t9 VDD1.t0 B.t5 sky130_fd_pr__nfet_01v8 ad=3.14655 pd=19.4 as=3.14655 ps=19.4 w=19.07 l=3.94
X22 VTAIL.t14 VN.t9 VDD2.t0 B.t5 sky130_fd_pr__nfet_01v8 ad=3.14655 pd=19.4 as=3.14655 ps=19.4 w=19.07 l=3.94
X23 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=7.4373 pd=38.92 as=0 ps=0 w=19.07 l=3.94
R0 VN.n112 VN.n111 161.3
R1 VN.n110 VN.n58 161.3
R2 VN.n109 VN.n108 161.3
R3 VN.n107 VN.n59 161.3
R4 VN.n106 VN.n105 161.3
R5 VN.n104 VN.n60 161.3
R6 VN.n103 VN.n102 161.3
R7 VN.n101 VN.n61 161.3
R8 VN.n100 VN.n99 161.3
R9 VN.n97 VN.n62 161.3
R10 VN.n96 VN.n95 161.3
R11 VN.n94 VN.n63 161.3
R12 VN.n93 VN.n92 161.3
R13 VN.n91 VN.n64 161.3
R14 VN.n90 VN.n89 161.3
R15 VN.n88 VN.n65 161.3
R16 VN.n87 VN.n86 161.3
R17 VN.n85 VN.n66 161.3
R18 VN.n84 VN.n83 161.3
R19 VN.n82 VN.n67 161.3
R20 VN.n81 VN.n80 161.3
R21 VN.n79 VN.n68 161.3
R22 VN.n78 VN.n77 161.3
R23 VN.n76 VN.n69 161.3
R24 VN.n75 VN.n74 161.3
R25 VN.n73 VN.n70 161.3
R26 VN.n55 VN.n54 161.3
R27 VN.n53 VN.n1 161.3
R28 VN.n52 VN.n51 161.3
R29 VN.n50 VN.n2 161.3
R30 VN.n49 VN.n48 161.3
R31 VN.n47 VN.n3 161.3
R32 VN.n46 VN.n45 161.3
R33 VN.n44 VN.n4 161.3
R34 VN.n43 VN.n42 161.3
R35 VN.n40 VN.n5 161.3
R36 VN.n39 VN.n38 161.3
R37 VN.n37 VN.n6 161.3
R38 VN.n36 VN.n35 161.3
R39 VN.n34 VN.n7 161.3
R40 VN.n33 VN.n32 161.3
R41 VN.n31 VN.n8 161.3
R42 VN.n30 VN.n29 161.3
R43 VN.n28 VN.n9 161.3
R44 VN.n27 VN.n26 161.3
R45 VN.n25 VN.n10 161.3
R46 VN.n24 VN.n23 161.3
R47 VN.n22 VN.n11 161.3
R48 VN.n21 VN.n20 161.3
R49 VN.n19 VN.n12 161.3
R50 VN.n18 VN.n17 161.3
R51 VN.n16 VN.n13 161.3
R52 VN.n71 VN.t5 149.214
R53 VN.n14 VN.t3 149.214
R54 VN.n28 VN.t2 116.647
R55 VN.n15 VN.t9 116.647
R56 VN.n41 VN.t4 116.647
R57 VN.n0 VN.t7 116.647
R58 VN.n85 VN.t0 116.647
R59 VN.n72 VN.t6 116.647
R60 VN.n98 VN.t1 116.647
R61 VN.n57 VN.t8 116.647
R62 VN.n56 VN.n0 88.1101
R63 VN.n113 VN.n57 88.1101
R64 VN VN.n113 65.9942
R65 VN.n15 VN.n14 61.9406
R66 VN.n72 VN.n71 61.9406
R67 VN.n22 VN.n21 53.6055
R68 VN.n35 VN.n34 53.6055
R69 VN.n79 VN.n78 53.6055
R70 VN.n92 VN.n91 53.6055
R71 VN.n48 VN.n47 49.7204
R72 VN.n105 VN.n104 49.7204
R73 VN.n48 VN.n2 31.2664
R74 VN.n105 VN.n59 31.2664
R75 VN.n23 VN.n22 27.3813
R76 VN.n34 VN.n33 27.3813
R77 VN.n80 VN.n79 27.3813
R78 VN.n91 VN.n90 27.3813
R79 VN.n17 VN.n16 24.4675
R80 VN.n17 VN.n12 24.4675
R81 VN.n21 VN.n12 24.4675
R82 VN.n23 VN.n10 24.4675
R83 VN.n27 VN.n10 24.4675
R84 VN.n28 VN.n27 24.4675
R85 VN.n29 VN.n28 24.4675
R86 VN.n29 VN.n8 24.4675
R87 VN.n33 VN.n8 24.4675
R88 VN.n35 VN.n6 24.4675
R89 VN.n39 VN.n6 24.4675
R90 VN.n40 VN.n39 24.4675
R91 VN.n42 VN.n4 24.4675
R92 VN.n46 VN.n4 24.4675
R93 VN.n47 VN.n46 24.4675
R94 VN.n52 VN.n2 24.4675
R95 VN.n53 VN.n52 24.4675
R96 VN.n54 VN.n53 24.4675
R97 VN.n78 VN.n69 24.4675
R98 VN.n74 VN.n69 24.4675
R99 VN.n74 VN.n73 24.4675
R100 VN.n90 VN.n65 24.4675
R101 VN.n86 VN.n65 24.4675
R102 VN.n86 VN.n85 24.4675
R103 VN.n85 VN.n84 24.4675
R104 VN.n84 VN.n67 24.4675
R105 VN.n80 VN.n67 24.4675
R106 VN.n104 VN.n103 24.4675
R107 VN.n103 VN.n61 24.4675
R108 VN.n99 VN.n61 24.4675
R109 VN.n97 VN.n96 24.4675
R110 VN.n96 VN.n63 24.4675
R111 VN.n92 VN.n63 24.4675
R112 VN.n111 VN.n110 24.4675
R113 VN.n110 VN.n109 24.4675
R114 VN.n109 VN.n59 24.4675
R115 VN.n16 VN.n15 13.2127
R116 VN.n41 VN.n40 13.2127
R117 VN.n73 VN.n72 13.2127
R118 VN.n98 VN.n97 13.2127
R119 VN.n42 VN.n41 11.2553
R120 VN.n99 VN.n98 11.2553
R121 VN.n71 VN.n70 2.48786
R122 VN.n14 VN.n13 2.48786
R123 VN.n54 VN.n0 1.95786
R124 VN.n111 VN.n57 1.95786
R125 VN.n113 VN.n112 0.354971
R126 VN.n56 VN.n55 0.354971
R127 VN VN.n56 0.26696
R128 VN.n112 VN.n58 0.189894
R129 VN.n108 VN.n58 0.189894
R130 VN.n108 VN.n107 0.189894
R131 VN.n107 VN.n106 0.189894
R132 VN.n106 VN.n60 0.189894
R133 VN.n102 VN.n60 0.189894
R134 VN.n102 VN.n101 0.189894
R135 VN.n101 VN.n100 0.189894
R136 VN.n100 VN.n62 0.189894
R137 VN.n95 VN.n62 0.189894
R138 VN.n95 VN.n94 0.189894
R139 VN.n94 VN.n93 0.189894
R140 VN.n93 VN.n64 0.189894
R141 VN.n89 VN.n64 0.189894
R142 VN.n89 VN.n88 0.189894
R143 VN.n88 VN.n87 0.189894
R144 VN.n87 VN.n66 0.189894
R145 VN.n83 VN.n66 0.189894
R146 VN.n83 VN.n82 0.189894
R147 VN.n82 VN.n81 0.189894
R148 VN.n81 VN.n68 0.189894
R149 VN.n77 VN.n68 0.189894
R150 VN.n77 VN.n76 0.189894
R151 VN.n76 VN.n75 0.189894
R152 VN.n75 VN.n70 0.189894
R153 VN.n18 VN.n13 0.189894
R154 VN.n19 VN.n18 0.189894
R155 VN.n20 VN.n19 0.189894
R156 VN.n20 VN.n11 0.189894
R157 VN.n24 VN.n11 0.189894
R158 VN.n25 VN.n24 0.189894
R159 VN.n26 VN.n25 0.189894
R160 VN.n26 VN.n9 0.189894
R161 VN.n30 VN.n9 0.189894
R162 VN.n31 VN.n30 0.189894
R163 VN.n32 VN.n31 0.189894
R164 VN.n32 VN.n7 0.189894
R165 VN.n36 VN.n7 0.189894
R166 VN.n37 VN.n36 0.189894
R167 VN.n38 VN.n37 0.189894
R168 VN.n38 VN.n5 0.189894
R169 VN.n43 VN.n5 0.189894
R170 VN.n44 VN.n43 0.189894
R171 VN.n45 VN.n44 0.189894
R172 VN.n45 VN.n3 0.189894
R173 VN.n49 VN.n3 0.189894
R174 VN.n50 VN.n49 0.189894
R175 VN.n51 VN.n50 0.189894
R176 VN.n51 VN.n1 0.189894
R177 VN.n55 VN.n1 0.189894
R178 VTAIL.n11 VTAIL.t15 46.6923
R179 VTAIL.n17 VTAIL.t7 46.6922
R180 VTAIL.n2 VTAIL.t16 46.6922
R181 VTAIL.n16 VTAIL.t0 46.6922
R182 VTAIL.n15 VTAIL.n14 45.6541
R183 VTAIL.n13 VTAIL.n12 45.6541
R184 VTAIL.n10 VTAIL.n9 45.6541
R185 VTAIL.n8 VTAIL.n7 45.6541
R186 VTAIL.n19 VTAIL.n18 45.6529
R187 VTAIL.n1 VTAIL.n0 45.6529
R188 VTAIL.n4 VTAIL.n3 45.6529
R189 VTAIL.n6 VTAIL.n5 45.6529
R190 VTAIL.n8 VTAIL.n6 36.1686
R191 VTAIL.n17 VTAIL.n16 32.4876
R192 VTAIL.n10 VTAIL.n8 3.68153
R193 VTAIL.n11 VTAIL.n10 3.68153
R194 VTAIL.n15 VTAIL.n13 3.68153
R195 VTAIL.n16 VTAIL.n15 3.68153
R196 VTAIL.n6 VTAIL.n4 3.68153
R197 VTAIL.n4 VTAIL.n2 3.68153
R198 VTAIL.n19 VTAIL.n17 3.68153
R199 VTAIL VTAIL.n1 2.81947
R200 VTAIL.n13 VTAIL.n11 2.31084
R201 VTAIL.n2 VTAIL.n1 2.31084
R202 VTAIL.n18 VTAIL.t10 1.03878
R203 VTAIL.n18 VTAIL.t12 1.03878
R204 VTAIL.n0 VTAIL.t11 1.03878
R205 VTAIL.n0 VTAIL.t14 1.03878
R206 VTAIL.n3 VTAIL.t17 1.03878
R207 VTAIL.n3 VTAIL.t1 1.03878
R208 VTAIL.n5 VTAIL.t2 1.03878
R209 VTAIL.n5 VTAIL.t19 1.03878
R210 VTAIL.n14 VTAIL.t4 1.03878
R211 VTAIL.n14 VTAIL.t18 1.03878
R212 VTAIL.n12 VTAIL.t3 1.03878
R213 VTAIL.n12 VTAIL.t5 1.03878
R214 VTAIL.n9 VTAIL.t6 1.03878
R215 VTAIL.n9 VTAIL.t13 1.03878
R216 VTAIL.n7 VTAIL.t8 1.03878
R217 VTAIL.n7 VTAIL.t9 1.03878
R218 VTAIL VTAIL.n19 0.862569
R219 VDD2.n1 VDD2.t6 67.052
R220 VDD2.n3 VDD2.n2 65.0371
R221 VDD2 VDD2.n7 65.0353
R222 VDD2.n4 VDD2.t1 63.3711
R223 VDD2.n6 VDD2.n5 62.3329
R224 VDD2.n1 VDD2.n0 62.3317
R225 VDD2.n4 VDD2.n3 57.6399
R226 VDD2.n6 VDD2.n4 3.68153
R227 VDD2.n7 VDD2.t3 1.03878
R228 VDD2.n7 VDD2.t4 1.03878
R229 VDD2.n5 VDD2.t8 1.03878
R230 VDD2.n5 VDD2.t9 1.03878
R231 VDD2.n2 VDD2.t5 1.03878
R232 VDD2.n2 VDD2.t2 1.03878
R233 VDD2.n0 VDD2.t0 1.03878
R234 VDD2.n0 VDD2.t7 1.03878
R235 VDD2 VDD2.n6 0.978948
R236 VDD2.n3 VDD2.n1 0.865413
R237 B.n1347 B.n1346 585
R238 B.n486 B.n218 585
R239 B.n485 B.n484 585
R240 B.n483 B.n482 585
R241 B.n481 B.n480 585
R242 B.n479 B.n478 585
R243 B.n477 B.n476 585
R244 B.n475 B.n474 585
R245 B.n473 B.n472 585
R246 B.n471 B.n470 585
R247 B.n469 B.n468 585
R248 B.n467 B.n466 585
R249 B.n465 B.n464 585
R250 B.n463 B.n462 585
R251 B.n461 B.n460 585
R252 B.n459 B.n458 585
R253 B.n457 B.n456 585
R254 B.n455 B.n454 585
R255 B.n453 B.n452 585
R256 B.n451 B.n450 585
R257 B.n449 B.n448 585
R258 B.n447 B.n446 585
R259 B.n445 B.n444 585
R260 B.n443 B.n442 585
R261 B.n441 B.n440 585
R262 B.n439 B.n438 585
R263 B.n437 B.n436 585
R264 B.n435 B.n434 585
R265 B.n433 B.n432 585
R266 B.n431 B.n430 585
R267 B.n429 B.n428 585
R268 B.n427 B.n426 585
R269 B.n425 B.n424 585
R270 B.n423 B.n422 585
R271 B.n421 B.n420 585
R272 B.n419 B.n418 585
R273 B.n417 B.n416 585
R274 B.n415 B.n414 585
R275 B.n413 B.n412 585
R276 B.n411 B.n410 585
R277 B.n409 B.n408 585
R278 B.n407 B.n406 585
R279 B.n405 B.n404 585
R280 B.n403 B.n402 585
R281 B.n401 B.n400 585
R282 B.n399 B.n398 585
R283 B.n397 B.n396 585
R284 B.n395 B.n394 585
R285 B.n393 B.n392 585
R286 B.n391 B.n390 585
R287 B.n389 B.n388 585
R288 B.n387 B.n386 585
R289 B.n385 B.n384 585
R290 B.n383 B.n382 585
R291 B.n381 B.n380 585
R292 B.n379 B.n378 585
R293 B.n377 B.n376 585
R294 B.n375 B.n374 585
R295 B.n373 B.n372 585
R296 B.n371 B.n370 585
R297 B.n369 B.n368 585
R298 B.n367 B.n366 585
R299 B.n365 B.n364 585
R300 B.n363 B.n362 585
R301 B.n361 B.n360 585
R302 B.n359 B.n358 585
R303 B.n357 B.n356 585
R304 B.n355 B.n354 585
R305 B.n353 B.n352 585
R306 B.n351 B.n350 585
R307 B.n349 B.n348 585
R308 B.n347 B.n346 585
R309 B.n345 B.n344 585
R310 B.n343 B.n342 585
R311 B.n341 B.n340 585
R312 B.n339 B.n338 585
R313 B.n337 B.n336 585
R314 B.n335 B.n334 585
R315 B.n333 B.n332 585
R316 B.n331 B.n330 585
R317 B.n329 B.n328 585
R318 B.n327 B.n326 585
R319 B.n325 B.n324 585
R320 B.n323 B.n322 585
R321 B.n321 B.n320 585
R322 B.n319 B.n318 585
R323 B.n317 B.n316 585
R324 B.n315 B.n314 585
R325 B.n313 B.n312 585
R326 B.n311 B.n310 585
R327 B.n309 B.n308 585
R328 B.n307 B.n306 585
R329 B.n305 B.n304 585
R330 B.n303 B.n302 585
R331 B.n301 B.n300 585
R332 B.n299 B.n298 585
R333 B.n297 B.n296 585
R334 B.n295 B.n294 585
R335 B.n293 B.n292 585
R336 B.n291 B.n290 585
R337 B.n289 B.n288 585
R338 B.n287 B.n286 585
R339 B.n285 B.n284 585
R340 B.n283 B.n282 585
R341 B.n281 B.n280 585
R342 B.n279 B.n278 585
R343 B.n277 B.n276 585
R344 B.n275 B.n274 585
R345 B.n273 B.n272 585
R346 B.n271 B.n270 585
R347 B.n269 B.n268 585
R348 B.n267 B.n266 585
R349 B.n265 B.n264 585
R350 B.n263 B.n262 585
R351 B.n261 B.n260 585
R352 B.n259 B.n258 585
R353 B.n257 B.n256 585
R354 B.n255 B.n254 585
R355 B.n253 B.n252 585
R356 B.n251 B.n250 585
R357 B.n249 B.n248 585
R358 B.n247 B.n246 585
R359 B.n245 B.n244 585
R360 B.n243 B.n242 585
R361 B.n241 B.n240 585
R362 B.n239 B.n238 585
R363 B.n237 B.n236 585
R364 B.n235 B.n234 585
R365 B.n233 B.n232 585
R366 B.n231 B.n230 585
R367 B.n229 B.n228 585
R368 B.n227 B.n226 585
R369 B.n152 B.n151 585
R370 B.n1352 B.n1351 585
R371 B.n1345 B.n219 585
R372 B.n219 B.n149 585
R373 B.n1344 B.n148 585
R374 B.n1356 B.n148 585
R375 B.n1343 B.n147 585
R376 B.n1357 B.n147 585
R377 B.n1342 B.n146 585
R378 B.n1358 B.n146 585
R379 B.n1341 B.n1340 585
R380 B.n1340 B.n142 585
R381 B.n1339 B.n141 585
R382 B.n1364 B.n141 585
R383 B.n1338 B.n140 585
R384 B.n1365 B.n140 585
R385 B.n1337 B.n139 585
R386 B.n1366 B.n139 585
R387 B.n1336 B.n1335 585
R388 B.n1335 B.n135 585
R389 B.n1334 B.n134 585
R390 B.n1372 B.n134 585
R391 B.n1333 B.n133 585
R392 B.n1373 B.n133 585
R393 B.n1332 B.n132 585
R394 B.n1374 B.n132 585
R395 B.n1331 B.n1330 585
R396 B.n1330 B.n128 585
R397 B.n1329 B.n127 585
R398 B.n1380 B.n127 585
R399 B.n1328 B.n126 585
R400 B.n1381 B.n126 585
R401 B.n1327 B.n125 585
R402 B.n1382 B.n125 585
R403 B.n1326 B.n1325 585
R404 B.n1325 B.n121 585
R405 B.n1324 B.n120 585
R406 B.n1388 B.n120 585
R407 B.n1323 B.n119 585
R408 B.n1389 B.n119 585
R409 B.n1322 B.n118 585
R410 B.n1390 B.n118 585
R411 B.n1321 B.n1320 585
R412 B.n1320 B.n114 585
R413 B.n1319 B.n113 585
R414 B.n1396 B.n113 585
R415 B.n1318 B.n112 585
R416 B.n1397 B.n112 585
R417 B.n1317 B.n111 585
R418 B.n1398 B.n111 585
R419 B.n1316 B.n1315 585
R420 B.n1315 B.n107 585
R421 B.n1314 B.n106 585
R422 B.n1404 B.n106 585
R423 B.n1313 B.n105 585
R424 B.n1405 B.n105 585
R425 B.n1312 B.n104 585
R426 B.n1406 B.n104 585
R427 B.n1311 B.n1310 585
R428 B.n1310 B.n100 585
R429 B.n1309 B.n99 585
R430 B.n1412 B.n99 585
R431 B.n1308 B.n98 585
R432 B.n1413 B.n98 585
R433 B.n1307 B.n97 585
R434 B.n1414 B.n97 585
R435 B.n1306 B.n1305 585
R436 B.n1305 B.n93 585
R437 B.n1304 B.n92 585
R438 B.n1420 B.n92 585
R439 B.n1303 B.n91 585
R440 B.n1421 B.n91 585
R441 B.n1302 B.n90 585
R442 B.n1422 B.n90 585
R443 B.n1301 B.n1300 585
R444 B.n1300 B.n86 585
R445 B.n1299 B.n85 585
R446 B.n1428 B.n85 585
R447 B.n1298 B.n84 585
R448 B.n1429 B.n84 585
R449 B.n1297 B.n83 585
R450 B.n1430 B.n83 585
R451 B.n1296 B.n1295 585
R452 B.n1295 B.n79 585
R453 B.n1294 B.n78 585
R454 B.n1436 B.n78 585
R455 B.n1293 B.n77 585
R456 B.n1437 B.n77 585
R457 B.n1292 B.n76 585
R458 B.n1438 B.n76 585
R459 B.n1291 B.n1290 585
R460 B.n1290 B.n72 585
R461 B.n1289 B.n71 585
R462 B.n1444 B.n71 585
R463 B.n1288 B.n70 585
R464 B.n1445 B.n70 585
R465 B.n1287 B.n69 585
R466 B.n1446 B.n69 585
R467 B.n1286 B.n1285 585
R468 B.n1285 B.n65 585
R469 B.n1284 B.n64 585
R470 B.n1452 B.n64 585
R471 B.n1283 B.n63 585
R472 B.n1453 B.n63 585
R473 B.n1282 B.n62 585
R474 B.n1454 B.n62 585
R475 B.n1281 B.n1280 585
R476 B.n1280 B.n58 585
R477 B.n1279 B.n57 585
R478 B.n1460 B.n57 585
R479 B.n1278 B.n56 585
R480 B.n1461 B.n56 585
R481 B.n1277 B.n55 585
R482 B.n1462 B.n55 585
R483 B.n1276 B.n1275 585
R484 B.n1275 B.n51 585
R485 B.n1274 B.n50 585
R486 B.n1468 B.n50 585
R487 B.n1273 B.n49 585
R488 B.n1469 B.n49 585
R489 B.n1272 B.n48 585
R490 B.n1470 B.n48 585
R491 B.n1271 B.n1270 585
R492 B.n1270 B.n44 585
R493 B.n1269 B.n43 585
R494 B.n1476 B.n43 585
R495 B.n1268 B.n42 585
R496 B.n1477 B.n42 585
R497 B.n1267 B.n41 585
R498 B.n1478 B.n41 585
R499 B.n1266 B.n1265 585
R500 B.n1265 B.n37 585
R501 B.n1264 B.n36 585
R502 B.n1484 B.n36 585
R503 B.n1263 B.n35 585
R504 B.n1485 B.n35 585
R505 B.n1262 B.n34 585
R506 B.n1486 B.n34 585
R507 B.n1261 B.n1260 585
R508 B.n1260 B.n30 585
R509 B.n1259 B.n29 585
R510 B.n1492 B.n29 585
R511 B.n1258 B.n28 585
R512 B.n1493 B.n28 585
R513 B.n1257 B.n27 585
R514 B.n1494 B.n27 585
R515 B.n1256 B.n1255 585
R516 B.n1255 B.n23 585
R517 B.n1254 B.n22 585
R518 B.n1500 B.n22 585
R519 B.n1253 B.n21 585
R520 B.n1501 B.n21 585
R521 B.n1252 B.n20 585
R522 B.n1502 B.n20 585
R523 B.n1251 B.n1250 585
R524 B.n1250 B.n16 585
R525 B.n1249 B.n15 585
R526 B.n1508 B.n15 585
R527 B.n1248 B.n14 585
R528 B.n1509 B.n14 585
R529 B.n1247 B.n13 585
R530 B.n1510 B.n13 585
R531 B.n1246 B.n1245 585
R532 B.n1245 B.n12 585
R533 B.n1244 B.n1243 585
R534 B.n1244 B.n8 585
R535 B.n1242 B.n7 585
R536 B.n1517 B.n7 585
R537 B.n1241 B.n6 585
R538 B.n1518 B.n6 585
R539 B.n1240 B.n5 585
R540 B.n1519 B.n5 585
R541 B.n1239 B.n1238 585
R542 B.n1238 B.n4 585
R543 B.n1237 B.n487 585
R544 B.n1237 B.n1236 585
R545 B.n1227 B.n488 585
R546 B.n489 B.n488 585
R547 B.n1229 B.n1228 585
R548 B.n1230 B.n1229 585
R549 B.n1226 B.n494 585
R550 B.n494 B.n493 585
R551 B.n1225 B.n1224 585
R552 B.n1224 B.n1223 585
R553 B.n496 B.n495 585
R554 B.n497 B.n496 585
R555 B.n1216 B.n1215 585
R556 B.n1217 B.n1216 585
R557 B.n1214 B.n502 585
R558 B.n502 B.n501 585
R559 B.n1213 B.n1212 585
R560 B.n1212 B.n1211 585
R561 B.n504 B.n503 585
R562 B.n505 B.n504 585
R563 B.n1204 B.n1203 585
R564 B.n1205 B.n1204 585
R565 B.n1202 B.n510 585
R566 B.n510 B.n509 585
R567 B.n1201 B.n1200 585
R568 B.n1200 B.n1199 585
R569 B.n512 B.n511 585
R570 B.n513 B.n512 585
R571 B.n1192 B.n1191 585
R572 B.n1193 B.n1192 585
R573 B.n1190 B.n518 585
R574 B.n518 B.n517 585
R575 B.n1189 B.n1188 585
R576 B.n1188 B.n1187 585
R577 B.n520 B.n519 585
R578 B.n521 B.n520 585
R579 B.n1180 B.n1179 585
R580 B.n1181 B.n1180 585
R581 B.n1178 B.n526 585
R582 B.n526 B.n525 585
R583 B.n1177 B.n1176 585
R584 B.n1176 B.n1175 585
R585 B.n528 B.n527 585
R586 B.n529 B.n528 585
R587 B.n1168 B.n1167 585
R588 B.n1169 B.n1168 585
R589 B.n1166 B.n534 585
R590 B.n534 B.n533 585
R591 B.n1165 B.n1164 585
R592 B.n1164 B.n1163 585
R593 B.n536 B.n535 585
R594 B.n537 B.n536 585
R595 B.n1156 B.n1155 585
R596 B.n1157 B.n1156 585
R597 B.n1154 B.n542 585
R598 B.n542 B.n541 585
R599 B.n1153 B.n1152 585
R600 B.n1152 B.n1151 585
R601 B.n544 B.n543 585
R602 B.n545 B.n544 585
R603 B.n1144 B.n1143 585
R604 B.n1145 B.n1144 585
R605 B.n1142 B.n549 585
R606 B.n553 B.n549 585
R607 B.n1141 B.n1140 585
R608 B.n1140 B.n1139 585
R609 B.n551 B.n550 585
R610 B.n552 B.n551 585
R611 B.n1132 B.n1131 585
R612 B.n1133 B.n1132 585
R613 B.n1130 B.n558 585
R614 B.n558 B.n557 585
R615 B.n1129 B.n1128 585
R616 B.n1128 B.n1127 585
R617 B.n560 B.n559 585
R618 B.n561 B.n560 585
R619 B.n1120 B.n1119 585
R620 B.n1121 B.n1120 585
R621 B.n1118 B.n566 585
R622 B.n566 B.n565 585
R623 B.n1117 B.n1116 585
R624 B.n1116 B.n1115 585
R625 B.n568 B.n567 585
R626 B.n569 B.n568 585
R627 B.n1108 B.n1107 585
R628 B.n1109 B.n1108 585
R629 B.n1106 B.n574 585
R630 B.n574 B.n573 585
R631 B.n1105 B.n1104 585
R632 B.n1104 B.n1103 585
R633 B.n576 B.n575 585
R634 B.n577 B.n576 585
R635 B.n1096 B.n1095 585
R636 B.n1097 B.n1096 585
R637 B.n1094 B.n582 585
R638 B.n582 B.n581 585
R639 B.n1093 B.n1092 585
R640 B.n1092 B.n1091 585
R641 B.n584 B.n583 585
R642 B.n585 B.n584 585
R643 B.n1084 B.n1083 585
R644 B.n1085 B.n1084 585
R645 B.n1082 B.n590 585
R646 B.n590 B.n589 585
R647 B.n1081 B.n1080 585
R648 B.n1080 B.n1079 585
R649 B.n592 B.n591 585
R650 B.n593 B.n592 585
R651 B.n1072 B.n1071 585
R652 B.n1073 B.n1072 585
R653 B.n1070 B.n598 585
R654 B.n598 B.n597 585
R655 B.n1069 B.n1068 585
R656 B.n1068 B.n1067 585
R657 B.n600 B.n599 585
R658 B.n601 B.n600 585
R659 B.n1060 B.n1059 585
R660 B.n1061 B.n1060 585
R661 B.n1058 B.n606 585
R662 B.n606 B.n605 585
R663 B.n1057 B.n1056 585
R664 B.n1056 B.n1055 585
R665 B.n608 B.n607 585
R666 B.n609 B.n608 585
R667 B.n1048 B.n1047 585
R668 B.n1049 B.n1048 585
R669 B.n1046 B.n614 585
R670 B.n614 B.n613 585
R671 B.n1045 B.n1044 585
R672 B.n1044 B.n1043 585
R673 B.n616 B.n615 585
R674 B.n617 B.n616 585
R675 B.n1036 B.n1035 585
R676 B.n1037 B.n1036 585
R677 B.n1034 B.n622 585
R678 B.n622 B.n621 585
R679 B.n1033 B.n1032 585
R680 B.n1032 B.n1031 585
R681 B.n624 B.n623 585
R682 B.n625 B.n624 585
R683 B.n1024 B.n1023 585
R684 B.n1025 B.n1024 585
R685 B.n1022 B.n630 585
R686 B.n630 B.n629 585
R687 B.n1021 B.n1020 585
R688 B.n1020 B.n1019 585
R689 B.n632 B.n631 585
R690 B.n633 B.n632 585
R691 B.n1012 B.n1011 585
R692 B.n1013 B.n1012 585
R693 B.n1010 B.n638 585
R694 B.n638 B.n637 585
R695 B.n1009 B.n1008 585
R696 B.n1008 B.n1007 585
R697 B.n640 B.n639 585
R698 B.n641 B.n640 585
R699 B.n1000 B.n999 585
R700 B.n1001 B.n1000 585
R701 B.n998 B.n646 585
R702 B.n646 B.n645 585
R703 B.n997 B.n996 585
R704 B.n996 B.n995 585
R705 B.n648 B.n647 585
R706 B.n649 B.n648 585
R707 B.n991 B.n990 585
R708 B.n652 B.n651 585
R709 B.n987 B.n986 585
R710 B.n988 B.n987 585
R711 B.n985 B.n719 585
R712 B.n984 B.n983 585
R713 B.n982 B.n981 585
R714 B.n980 B.n979 585
R715 B.n978 B.n977 585
R716 B.n976 B.n975 585
R717 B.n974 B.n973 585
R718 B.n972 B.n971 585
R719 B.n970 B.n969 585
R720 B.n968 B.n967 585
R721 B.n966 B.n965 585
R722 B.n964 B.n963 585
R723 B.n962 B.n961 585
R724 B.n960 B.n959 585
R725 B.n958 B.n957 585
R726 B.n956 B.n955 585
R727 B.n954 B.n953 585
R728 B.n952 B.n951 585
R729 B.n950 B.n949 585
R730 B.n948 B.n947 585
R731 B.n946 B.n945 585
R732 B.n944 B.n943 585
R733 B.n942 B.n941 585
R734 B.n940 B.n939 585
R735 B.n938 B.n937 585
R736 B.n936 B.n935 585
R737 B.n934 B.n933 585
R738 B.n932 B.n931 585
R739 B.n930 B.n929 585
R740 B.n928 B.n927 585
R741 B.n926 B.n925 585
R742 B.n924 B.n923 585
R743 B.n922 B.n921 585
R744 B.n920 B.n919 585
R745 B.n918 B.n917 585
R746 B.n916 B.n915 585
R747 B.n914 B.n913 585
R748 B.n912 B.n911 585
R749 B.n910 B.n909 585
R750 B.n908 B.n907 585
R751 B.n906 B.n905 585
R752 B.n904 B.n903 585
R753 B.n902 B.n901 585
R754 B.n900 B.n899 585
R755 B.n898 B.n897 585
R756 B.n896 B.n895 585
R757 B.n894 B.n893 585
R758 B.n892 B.n891 585
R759 B.n890 B.n889 585
R760 B.n888 B.n887 585
R761 B.n886 B.n885 585
R762 B.n884 B.n883 585
R763 B.n882 B.n881 585
R764 B.n880 B.n879 585
R765 B.n878 B.n877 585
R766 B.n876 B.n875 585
R767 B.n874 B.n873 585
R768 B.n872 B.n871 585
R769 B.n870 B.n869 585
R770 B.n867 B.n866 585
R771 B.n865 B.n864 585
R772 B.n863 B.n862 585
R773 B.n861 B.n860 585
R774 B.n859 B.n858 585
R775 B.n857 B.n856 585
R776 B.n855 B.n854 585
R777 B.n853 B.n852 585
R778 B.n851 B.n850 585
R779 B.n849 B.n848 585
R780 B.n846 B.n845 585
R781 B.n844 B.n843 585
R782 B.n842 B.n841 585
R783 B.n840 B.n839 585
R784 B.n838 B.n837 585
R785 B.n836 B.n835 585
R786 B.n834 B.n833 585
R787 B.n832 B.n831 585
R788 B.n830 B.n829 585
R789 B.n828 B.n827 585
R790 B.n826 B.n825 585
R791 B.n824 B.n823 585
R792 B.n822 B.n821 585
R793 B.n820 B.n819 585
R794 B.n818 B.n817 585
R795 B.n816 B.n815 585
R796 B.n814 B.n813 585
R797 B.n812 B.n811 585
R798 B.n810 B.n809 585
R799 B.n808 B.n807 585
R800 B.n806 B.n805 585
R801 B.n804 B.n803 585
R802 B.n802 B.n801 585
R803 B.n800 B.n799 585
R804 B.n798 B.n797 585
R805 B.n796 B.n795 585
R806 B.n794 B.n793 585
R807 B.n792 B.n791 585
R808 B.n790 B.n789 585
R809 B.n788 B.n787 585
R810 B.n786 B.n785 585
R811 B.n784 B.n783 585
R812 B.n782 B.n781 585
R813 B.n780 B.n779 585
R814 B.n778 B.n777 585
R815 B.n776 B.n775 585
R816 B.n774 B.n773 585
R817 B.n772 B.n771 585
R818 B.n770 B.n769 585
R819 B.n768 B.n767 585
R820 B.n766 B.n765 585
R821 B.n764 B.n763 585
R822 B.n762 B.n761 585
R823 B.n760 B.n759 585
R824 B.n758 B.n757 585
R825 B.n756 B.n755 585
R826 B.n754 B.n753 585
R827 B.n752 B.n751 585
R828 B.n750 B.n749 585
R829 B.n748 B.n747 585
R830 B.n746 B.n745 585
R831 B.n744 B.n743 585
R832 B.n742 B.n741 585
R833 B.n740 B.n739 585
R834 B.n738 B.n737 585
R835 B.n736 B.n735 585
R836 B.n734 B.n733 585
R837 B.n732 B.n731 585
R838 B.n730 B.n729 585
R839 B.n728 B.n727 585
R840 B.n726 B.n725 585
R841 B.n724 B.n718 585
R842 B.n988 B.n718 585
R843 B.n992 B.n650 585
R844 B.n650 B.n649 585
R845 B.n994 B.n993 585
R846 B.n995 B.n994 585
R847 B.n644 B.n643 585
R848 B.n645 B.n644 585
R849 B.n1003 B.n1002 585
R850 B.n1002 B.n1001 585
R851 B.n1004 B.n642 585
R852 B.n642 B.n641 585
R853 B.n1006 B.n1005 585
R854 B.n1007 B.n1006 585
R855 B.n636 B.n635 585
R856 B.n637 B.n636 585
R857 B.n1015 B.n1014 585
R858 B.n1014 B.n1013 585
R859 B.n1016 B.n634 585
R860 B.n634 B.n633 585
R861 B.n1018 B.n1017 585
R862 B.n1019 B.n1018 585
R863 B.n628 B.n627 585
R864 B.n629 B.n628 585
R865 B.n1027 B.n1026 585
R866 B.n1026 B.n1025 585
R867 B.n1028 B.n626 585
R868 B.n626 B.n625 585
R869 B.n1030 B.n1029 585
R870 B.n1031 B.n1030 585
R871 B.n620 B.n619 585
R872 B.n621 B.n620 585
R873 B.n1039 B.n1038 585
R874 B.n1038 B.n1037 585
R875 B.n1040 B.n618 585
R876 B.n618 B.n617 585
R877 B.n1042 B.n1041 585
R878 B.n1043 B.n1042 585
R879 B.n612 B.n611 585
R880 B.n613 B.n612 585
R881 B.n1051 B.n1050 585
R882 B.n1050 B.n1049 585
R883 B.n1052 B.n610 585
R884 B.n610 B.n609 585
R885 B.n1054 B.n1053 585
R886 B.n1055 B.n1054 585
R887 B.n604 B.n603 585
R888 B.n605 B.n604 585
R889 B.n1063 B.n1062 585
R890 B.n1062 B.n1061 585
R891 B.n1064 B.n602 585
R892 B.n602 B.n601 585
R893 B.n1066 B.n1065 585
R894 B.n1067 B.n1066 585
R895 B.n596 B.n595 585
R896 B.n597 B.n596 585
R897 B.n1075 B.n1074 585
R898 B.n1074 B.n1073 585
R899 B.n1076 B.n594 585
R900 B.n594 B.n593 585
R901 B.n1078 B.n1077 585
R902 B.n1079 B.n1078 585
R903 B.n588 B.n587 585
R904 B.n589 B.n588 585
R905 B.n1087 B.n1086 585
R906 B.n1086 B.n1085 585
R907 B.n1088 B.n586 585
R908 B.n586 B.n585 585
R909 B.n1090 B.n1089 585
R910 B.n1091 B.n1090 585
R911 B.n580 B.n579 585
R912 B.n581 B.n580 585
R913 B.n1099 B.n1098 585
R914 B.n1098 B.n1097 585
R915 B.n1100 B.n578 585
R916 B.n578 B.n577 585
R917 B.n1102 B.n1101 585
R918 B.n1103 B.n1102 585
R919 B.n572 B.n571 585
R920 B.n573 B.n572 585
R921 B.n1111 B.n1110 585
R922 B.n1110 B.n1109 585
R923 B.n1112 B.n570 585
R924 B.n570 B.n569 585
R925 B.n1114 B.n1113 585
R926 B.n1115 B.n1114 585
R927 B.n564 B.n563 585
R928 B.n565 B.n564 585
R929 B.n1123 B.n1122 585
R930 B.n1122 B.n1121 585
R931 B.n1124 B.n562 585
R932 B.n562 B.n561 585
R933 B.n1126 B.n1125 585
R934 B.n1127 B.n1126 585
R935 B.n556 B.n555 585
R936 B.n557 B.n556 585
R937 B.n1135 B.n1134 585
R938 B.n1134 B.n1133 585
R939 B.n1136 B.n554 585
R940 B.n554 B.n552 585
R941 B.n1138 B.n1137 585
R942 B.n1139 B.n1138 585
R943 B.n548 B.n547 585
R944 B.n553 B.n548 585
R945 B.n1147 B.n1146 585
R946 B.n1146 B.n1145 585
R947 B.n1148 B.n546 585
R948 B.n546 B.n545 585
R949 B.n1150 B.n1149 585
R950 B.n1151 B.n1150 585
R951 B.n540 B.n539 585
R952 B.n541 B.n540 585
R953 B.n1159 B.n1158 585
R954 B.n1158 B.n1157 585
R955 B.n1160 B.n538 585
R956 B.n538 B.n537 585
R957 B.n1162 B.n1161 585
R958 B.n1163 B.n1162 585
R959 B.n532 B.n531 585
R960 B.n533 B.n532 585
R961 B.n1171 B.n1170 585
R962 B.n1170 B.n1169 585
R963 B.n1172 B.n530 585
R964 B.n530 B.n529 585
R965 B.n1174 B.n1173 585
R966 B.n1175 B.n1174 585
R967 B.n524 B.n523 585
R968 B.n525 B.n524 585
R969 B.n1183 B.n1182 585
R970 B.n1182 B.n1181 585
R971 B.n1184 B.n522 585
R972 B.n522 B.n521 585
R973 B.n1186 B.n1185 585
R974 B.n1187 B.n1186 585
R975 B.n516 B.n515 585
R976 B.n517 B.n516 585
R977 B.n1195 B.n1194 585
R978 B.n1194 B.n1193 585
R979 B.n1196 B.n514 585
R980 B.n514 B.n513 585
R981 B.n1198 B.n1197 585
R982 B.n1199 B.n1198 585
R983 B.n508 B.n507 585
R984 B.n509 B.n508 585
R985 B.n1207 B.n1206 585
R986 B.n1206 B.n1205 585
R987 B.n1208 B.n506 585
R988 B.n506 B.n505 585
R989 B.n1210 B.n1209 585
R990 B.n1211 B.n1210 585
R991 B.n500 B.n499 585
R992 B.n501 B.n500 585
R993 B.n1219 B.n1218 585
R994 B.n1218 B.n1217 585
R995 B.n1220 B.n498 585
R996 B.n498 B.n497 585
R997 B.n1222 B.n1221 585
R998 B.n1223 B.n1222 585
R999 B.n492 B.n491 585
R1000 B.n493 B.n492 585
R1001 B.n1232 B.n1231 585
R1002 B.n1231 B.n1230 585
R1003 B.n1233 B.n490 585
R1004 B.n490 B.n489 585
R1005 B.n1235 B.n1234 585
R1006 B.n1236 B.n1235 585
R1007 B.n3 B.n0 585
R1008 B.n4 B.n3 585
R1009 B.n1516 B.n1 585
R1010 B.n1517 B.n1516 585
R1011 B.n1515 B.n1514 585
R1012 B.n1515 B.n8 585
R1013 B.n1513 B.n9 585
R1014 B.n12 B.n9 585
R1015 B.n1512 B.n1511 585
R1016 B.n1511 B.n1510 585
R1017 B.n11 B.n10 585
R1018 B.n1509 B.n11 585
R1019 B.n1507 B.n1506 585
R1020 B.n1508 B.n1507 585
R1021 B.n1505 B.n17 585
R1022 B.n17 B.n16 585
R1023 B.n1504 B.n1503 585
R1024 B.n1503 B.n1502 585
R1025 B.n19 B.n18 585
R1026 B.n1501 B.n19 585
R1027 B.n1499 B.n1498 585
R1028 B.n1500 B.n1499 585
R1029 B.n1497 B.n24 585
R1030 B.n24 B.n23 585
R1031 B.n1496 B.n1495 585
R1032 B.n1495 B.n1494 585
R1033 B.n26 B.n25 585
R1034 B.n1493 B.n26 585
R1035 B.n1491 B.n1490 585
R1036 B.n1492 B.n1491 585
R1037 B.n1489 B.n31 585
R1038 B.n31 B.n30 585
R1039 B.n1488 B.n1487 585
R1040 B.n1487 B.n1486 585
R1041 B.n33 B.n32 585
R1042 B.n1485 B.n33 585
R1043 B.n1483 B.n1482 585
R1044 B.n1484 B.n1483 585
R1045 B.n1481 B.n38 585
R1046 B.n38 B.n37 585
R1047 B.n1480 B.n1479 585
R1048 B.n1479 B.n1478 585
R1049 B.n40 B.n39 585
R1050 B.n1477 B.n40 585
R1051 B.n1475 B.n1474 585
R1052 B.n1476 B.n1475 585
R1053 B.n1473 B.n45 585
R1054 B.n45 B.n44 585
R1055 B.n1472 B.n1471 585
R1056 B.n1471 B.n1470 585
R1057 B.n47 B.n46 585
R1058 B.n1469 B.n47 585
R1059 B.n1467 B.n1466 585
R1060 B.n1468 B.n1467 585
R1061 B.n1465 B.n52 585
R1062 B.n52 B.n51 585
R1063 B.n1464 B.n1463 585
R1064 B.n1463 B.n1462 585
R1065 B.n54 B.n53 585
R1066 B.n1461 B.n54 585
R1067 B.n1459 B.n1458 585
R1068 B.n1460 B.n1459 585
R1069 B.n1457 B.n59 585
R1070 B.n59 B.n58 585
R1071 B.n1456 B.n1455 585
R1072 B.n1455 B.n1454 585
R1073 B.n61 B.n60 585
R1074 B.n1453 B.n61 585
R1075 B.n1451 B.n1450 585
R1076 B.n1452 B.n1451 585
R1077 B.n1449 B.n66 585
R1078 B.n66 B.n65 585
R1079 B.n1448 B.n1447 585
R1080 B.n1447 B.n1446 585
R1081 B.n68 B.n67 585
R1082 B.n1445 B.n68 585
R1083 B.n1443 B.n1442 585
R1084 B.n1444 B.n1443 585
R1085 B.n1441 B.n73 585
R1086 B.n73 B.n72 585
R1087 B.n1440 B.n1439 585
R1088 B.n1439 B.n1438 585
R1089 B.n75 B.n74 585
R1090 B.n1437 B.n75 585
R1091 B.n1435 B.n1434 585
R1092 B.n1436 B.n1435 585
R1093 B.n1433 B.n80 585
R1094 B.n80 B.n79 585
R1095 B.n1432 B.n1431 585
R1096 B.n1431 B.n1430 585
R1097 B.n82 B.n81 585
R1098 B.n1429 B.n82 585
R1099 B.n1427 B.n1426 585
R1100 B.n1428 B.n1427 585
R1101 B.n1425 B.n87 585
R1102 B.n87 B.n86 585
R1103 B.n1424 B.n1423 585
R1104 B.n1423 B.n1422 585
R1105 B.n89 B.n88 585
R1106 B.n1421 B.n89 585
R1107 B.n1419 B.n1418 585
R1108 B.n1420 B.n1419 585
R1109 B.n1417 B.n94 585
R1110 B.n94 B.n93 585
R1111 B.n1416 B.n1415 585
R1112 B.n1415 B.n1414 585
R1113 B.n96 B.n95 585
R1114 B.n1413 B.n96 585
R1115 B.n1411 B.n1410 585
R1116 B.n1412 B.n1411 585
R1117 B.n1409 B.n101 585
R1118 B.n101 B.n100 585
R1119 B.n1408 B.n1407 585
R1120 B.n1407 B.n1406 585
R1121 B.n103 B.n102 585
R1122 B.n1405 B.n103 585
R1123 B.n1403 B.n1402 585
R1124 B.n1404 B.n1403 585
R1125 B.n1401 B.n108 585
R1126 B.n108 B.n107 585
R1127 B.n1400 B.n1399 585
R1128 B.n1399 B.n1398 585
R1129 B.n110 B.n109 585
R1130 B.n1397 B.n110 585
R1131 B.n1395 B.n1394 585
R1132 B.n1396 B.n1395 585
R1133 B.n1393 B.n115 585
R1134 B.n115 B.n114 585
R1135 B.n1392 B.n1391 585
R1136 B.n1391 B.n1390 585
R1137 B.n117 B.n116 585
R1138 B.n1389 B.n117 585
R1139 B.n1387 B.n1386 585
R1140 B.n1388 B.n1387 585
R1141 B.n1385 B.n122 585
R1142 B.n122 B.n121 585
R1143 B.n1384 B.n1383 585
R1144 B.n1383 B.n1382 585
R1145 B.n124 B.n123 585
R1146 B.n1381 B.n124 585
R1147 B.n1379 B.n1378 585
R1148 B.n1380 B.n1379 585
R1149 B.n1377 B.n129 585
R1150 B.n129 B.n128 585
R1151 B.n1376 B.n1375 585
R1152 B.n1375 B.n1374 585
R1153 B.n131 B.n130 585
R1154 B.n1373 B.n131 585
R1155 B.n1371 B.n1370 585
R1156 B.n1372 B.n1371 585
R1157 B.n1369 B.n136 585
R1158 B.n136 B.n135 585
R1159 B.n1368 B.n1367 585
R1160 B.n1367 B.n1366 585
R1161 B.n138 B.n137 585
R1162 B.n1365 B.n138 585
R1163 B.n1363 B.n1362 585
R1164 B.n1364 B.n1363 585
R1165 B.n1361 B.n143 585
R1166 B.n143 B.n142 585
R1167 B.n1360 B.n1359 585
R1168 B.n1359 B.n1358 585
R1169 B.n145 B.n144 585
R1170 B.n1357 B.n145 585
R1171 B.n1355 B.n1354 585
R1172 B.n1356 B.n1355 585
R1173 B.n1353 B.n150 585
R1174 B.n150 B.n149 585
R1175 B.n1520 B.n1519 585
R1176 B.n1518 B.n2 585
R1177 B.n1351 B.n150 526.135
R1178 B.n1347 B.n219 526.135
R1179 B.n718 B.n648 526.135
R1180 B.n990 B.n650 526.135
R1181 B.n223 B.t14 326.096
R1182 B.n220 B.t10 326.096
R1183 B.n722 B.t6 326.096
R1184 B.n720 B.t17 326.096
R1185 B.n1349 B.n1348 256.663
R1186 B.n1349 B.n217 256.663
R1187 B.n1349 B.n216 256.663
R1188 B.n1349 B.n215 256.663
R1189 B.n1349 B.n214 256.663
R1190 B.n1349 B.n213 256.663
R1191 B.n1349 B.n212 256.663
R1192 B.n1349 B.n211 256.663
R1193 B.n1349 B.n210 256.663
R1194 B.n1349 B.n209 256.663
R1195 B.n1349 B.n208 256.663
R1196 B.n1349 B.n207 256.663
R1197 B.n1349 B.n206 256.663
R1198 B.n1349 B.n205 256.663
R1199 B.n1349 B.n204 256.663
R1200 B.n1349 B.n203 256.663
R1201 B.n1349 B.n202 256.663
R1202 B.n1349 B.n201 256.663
R1203 B.n1349 B.n200 256.663
R1204 B.n1349 B.n199 256.663
R1205 B.n1349 B.n198 256.663
R1206 B.n1349 B.n197 256.663
R1207 B.n1349 B.n196 256.663
R1208 B.n1349 B.n195 256.663
R1209 B.n1349 B.n194 256.663
R1210 B.n1349 B.n193 256.663
R1211 B.n1349 B.n192 256.663
R1212 B.n1349 B.n191 256.663
R1213 B.n1349 B.n190 256.663
R1214 B.n1349 B.n189 256.663
R1215 B.n1349 B.n188 256.663
R1216 B.n1349 B.n187 256.663
R1217 B.n1349 B.n186 256.663
R1218 B.n1349 B.n185 256.663
R1219 B.n1349 B.n184 256.663
R1220 B.n1349 B.n183 256.663
R1221 B.n1349 B.n182 256.663
R1222 B.n1349 B.n181 256.663
R1223 B.n1349 B.n180 256.663
R1224 B.n1349 B.n179 256.663
R1225 B.n1349 B.n178 256.663
R1226 B.n1349 B.n177 256.663
R1227 B.n1349 B.n176 256.663
R1228 B.n1349 B.n175 256.663
R1229 B.n1349 B.n174 256.663
R1230 B.n1349 B.n173 256.663
R1231 B.n1349 B.n172 256.663
R1232 B.n1349 B.n171 256.663
R1233 B.n1349 B.n170 256.663
R1234 B.n1349 B.n169 256.663
R1235 B.n1349 B.n168 256.663
R1236 B.n1349 B.n167 256.663
R1237 B.n1349 B.n166 256.663
R1238 B.n1349 B.n165 256.663
R1239 B.n1349 B.n164 256.663
R1240 B.n1349 B.n163 256.663
R1241 B.n1349 B.n162 256.663
R1242 B.n1349 B.n161 256.663
R1243 B.n1349 B.n160 256.663
R1244 B.n1349 B.n159 256.663
R1245 B.n1349 B.n158 256.663
R1246 B.n1349 B.n157 256.663
R1247 B.n1349 B.n156 256.663
R1248 B.n1349 B.n155 256.663
R1249 B.n1349 B.n154 256.663
R1250 B.n1349 B.n153 256.663
R1251 B.n1350 B.n1349 256.663
R1252 B.n989 B.n988 256.663
R1253 B.n988 B.n653 256.663
R1254 B.n988 B.n654 256.663
R1255 B.n988 B.n655 256.663
R1256 B.n988 B.n656 256.663
R1257 B.n988 B.n657 256.663
R1258 B.n988 B.n658 256.663
R1259 B.n988 B.n659 256.663
R1260 B.n988 B.n660 256.663
R1261 B.n988 B.n661 256.663
R1262 B.n988 B.n662 256.663
R1263 B.n988 B.n663 256.663
R1264 B.n988 B.n664 256.663
R1265 B.n988 B.n665 256.663
R1266 B.n988 B.n666 256.663
R1267 B.n988 B.n667 256.663
R1268 B.n988 B.n668 256.663
R1269 B.n988 B.n669 256.663
R1270 B.n988 B.n670 256.663
R1271 B.n988 B.n671 256.663
R1272 B.n988 B.n672 256.663
R1273 B.n988 B.n673 256.663
R1274 B.n988 B.n674 256.663
R1275 B.n988 B.n675 256.663
R1276 B.n988 B.n676 256.663
R1277 B.n988 B.n677 256.663
R1278 B.n988 B.n678 256.663
R1279 B.n988 B.n679 256.663
R1280 B.n988 B.n680 256.663
R1281 B.n988 B.n681 256.663
R1282 B.n988 B.n682 256.663
R1283 B.n988 B.n683 256.663
R1284 B.n988 B.n684 256.663
R1285 B.n988 B.n685 256.663
R1286 B.n988 B.n686 256.663
R1287 B.n988 B.n687 256.663
R1288 B.n988 B.n688 256.663
R1289 B.n988 B.n689 256.663
R1290 B.n988 B.n690 256.663
R1291 B.n988 B.n691 256.663
R1292 B.n988 B.n692 256.663
R1293 B.n988 B.n693 256.663
R1294 B.n988 B.n694 256.663
R1295 B.n988 B.n695 256.663
R1296 B.n988 B.n696 256.663
R1297 B.n988 B.n697 256.663
R1298 B.n988 B.n698 256.663
R1299 B.n988 B.n699 256.663
R1300 B.n988 B.n700 256.663
R1301 B.n988 B.n701 256.663
R1302 B.n988 B.n702 256.663
R1303 B.n988 B.n703 256.663
R1304 B.n988 B.n704 256.663
R1305 B.n988 B.n705 256.663
R1306 B.n988 B.n706 256.663
R1307 B.n988 B.n707 256.663
R1308 B.n988 B.n708 256.663
R1309 B.n988 B.n709 256.663
R1310 B.n988 B.n710 256.663
R1311 B.n988 B.n711 256.663
R1312 B.n988 B.n712 256.663
R1313 B.n988 B.n713 256.663
R1314 B.n988 B.n714 256.663
R1315 B.n988 B.n715 256.663
R1316 B.n988 B.n716 256.663
R1317 B.n988 B.n717 256.663
R1318 B.n1522 B.n1521 256.663
R1319 B.n226 B.n152 163.367
R1320 B.n230 B.n229 163.367
R1321 B.n234 B.n233 163.367
R1322 B.n238 B.n237 163.367
R1323 B.n242 B.n241 163.367
R1324 B.n246 B.n245 163.367
R1325 B.n250 B.n249 163.367
R1326 B.n254 B.n253 163.367
R1327 B.n258 B.n257 163.367
R1328 B.n262 B.n261 163.367
R1329 B.n266 B.n265 163.367
R1330 B.n270 B.n269 163.367
R1331 B.n274 B.n273 163.367
R1332 B.n278 B.n277 163.367
R1333 B.n282 B.n281 163.367
R1334 B.n286 B.n285 163.367
R1335 B.n290 B.n289 163.367
R1336 B.n294 B.n293 163.367
R1337 B.n298 B.n297 163.367
R1338 B.n302 B.n301 163.367
R1339 B.n306 B.n305 163.367
R1340 B.n310 B.n309 163.367
R1341 B.n314 B.n313 163.367
R1342 B.n318 B.n317 163.367
R1343 B.n322 B.n321 163.367
R1344 B.n326 B.n325 163.367
R1345 B.n330 B.n329 163.367
R1346 B.n334 B.n333 163.367
R1347 B.n338 B.n337 163.367
R1348 B.n342 B.n341 163.367
R1349 B.n346 B.n345 163.367
R1350 B.n350 B.n349 163.367
R1351 B.n354 B.n353 163.367
R1352 B.n358 B.n357 163.367
R1353 B.n362 B.n361 163.367
R1354 B.n366 B.n365 163.367
R1355 B.n370 B.n369 163.367
R1356 B.n374 B.n373 163.367
R1357 B.n378 B.n377 163.367
R1358 B.n382 B.n381 163.367
R1359 B.n386 B.n385 163.367
R1360 B.n390 B.n389 163.367
R1361 B.n394 B.n393 163.367
R1362 B.n398 B.n397 163.367
R1363 B.n402 B.n401 163.367
R1364 B.n406 B.n405 163.367
R1365 B.n410 B.n409 163.367
R1366 B.n414 B.n413 163.367
R1367 B.n418 B.n417 163.367
R1368 B.n422 B.n421 163.367
R1369 B.n426 B.n425 163.367
R1370 B.n430 B.n429 163.367
R1371 B.n434 B.n433 163.367
R1372 B.n438 B.n437 163.367
R1373 B.n442 B.n441 163.367
R1374 B.n446 B.n445 163.367
R1375 B.n450 B.n449 163.367
R1376 B.n454 B.n453 163.367
R1377 B.n458 B.n457 163.367
R1378 B.n462 B.n461 163.367
R1379 B.n466 B.n465 163.367
R1380 B.n470 B.n469 163.367
R1381 B.n474 B.n473 163.367
R1382 B.n478 B.n477 163.367
R1383 B.n482 B.n481 163.367
R1384 B.n484 B.n218 163.367
R1385 B.n996 B.n648 163.367
R1386 B.n996 B.n646 163.367
R1387 B.n1000 B.n646 163.367
R1388 B.n1000 B.n640 163.367
R1389 B.n1008 B.n640 163.367
R1390 B.n1008 B.n638 163.367
R1391 B.n1012 B.n638 163.367
R1392 B.n1012 B.n632 163.367
R1393 B.n1020 B.n632 163.367
R1394 B.n1020 B.n630 163.367
R1395 B.n1024 B.n630 163.367
R1396 B.n1024 B.n624 163.367
R1397 B.n1032 B.n624 163.367
R1398 B.n1032 B.n622 163.367
R1399 B.n1036 B.n622 163.367
R1400 B.n1036 B.n616 163.367
R1401 B.n1044 B.n616 163.367
R1402 B.n1044 B.n614 163.367
R1403 B.n1048 B.n614 163.367
R1404 B.n1048 B.n608 163.367
R1405 B.n1056 B.n608 163.367
R1406 B.n1056 B.n606 163.367
R1407 B.n1060 B.n606 163.367
R1408 B.n1060 B.n600 163.367
R1409 B.n1068 B.n600 163.367
R1410 B.n1068 B.n598 163.367
R1411 B.n1072 B.n598 163.367
R1412 B.n1072 B.n592 163.367
R1413 B.n1080 B.n592 163.367
R1414 B.n1080 B.n590 163.367
R1415 B.n1084 B.n590 163.367
R1416 B.n1084 B.n584 163.367
R1417 B.n1092 B.n584 163.367
R1418 B.n1092 B.n582 163.367
R1419 B.n1096 B.n582 163.367
R1420 B.n1096 B.n576 163.367
R1421 B.n1104 B.n576 163.367
R1422 B.n1104 B.n574 163.367
R1423 B.n1108 B.n574 163.367
R1424 B.n1108 B.n568 163.367
R1425 B.n1116 B.n568 163.367
R1426 B.n1116 B.n566 163.367
R1427 B.n1120 B.n566 163.367
R1428 B.n1120 B.n560 163.367
R1429 B.n1128 B.n560 163.367
R1430 B.n1128 B.n558 163.367
R1431 B.n1132 B.n558 163.367
R1432 B.n1132 B.n551 163.367
R1433 B.n1140 B.n551 163.367
R1434 B.n1140 B.n549 163.367
R1435 B.n1144 B.n549 163.367
R1436 B.n1144 B.n544 163.367
R1437 B.n1152 B.n544 163.367
R1438 B.n1152 B.n542 163.367
R1439 B.n1156 B.n542 163.367
R1440 B.n1156 B.n536 163.367
R1441 B.n1164 B.n536 163.367
R1442 B.n1164 B.n534 163.367
R1443 B.n1168 B.n534 163.367
R1444 B.n1168 B.n528 163.367
R1445 B.n1176 B.n528 163.367
R1446 B.n1176 B.n526 163.367
R1447 B.n1180 B.n526 163.367
R1448 B.n1180 B.n520 163.367
R1449 B.n1188 B.n520 163.367
R1450 B.n1188 B.n518 163.367
R1451 B.n1192 B.n518 163.367
R1452 B.n1192 B.n512 163.367
R1453 B.n1200 B.n512 163.367
R1454 B.n1200 B.n510 163.367
R1455 B.n1204 B.n510 163.367
R1456 B.n1204 B.n504 163.367
R1457 B.n1212 B.n504 163.367
R1458 B.n1212 B.n502 163.367
R1459 B.n1216 B.n502 163.367
R1460 B.n1216 B.n496 163.367
R1461 B.n1224 B.n496 163.367
R1462 B.n1224 B.n494 163.367
R1463 B.n1229 B.n494 163.367
R1464 B.n1229 B.n488 163.367
R1465 B.n1237 B.n488 163.367
R1466 B.n1238 B.n1237 163.367
R1467 B.n1238 B.n5 163.367
R1468 B.n6 B.n5 163.367
R1469 B.n7 B.n6 163.367
R1470 B.n1244 B.n7 163.367
R1471 B.n1245 B.n1244 163.367
R1472 B.n1245 B.n13 163.367
R1473 B.n14 B.n13 163.367
R1474 B.n15 B.n14 163.367
R1475 B.n1250 B.n15 163.367
R1476 B.n1250 B.n20 163.367
R1477 B.n21 B.n20 163.367
R1478 B.n22 B.n21 163.367
R1479 B.n1255 B.n22 163.367
R1480 B.n1255 B.n27 163.367
R1481 B.n28 B.n27 163.367
R1482 B.n29 B.n28 163.367
R1483 B.n1260 B.n29 163.367
R1484 B.n1260 B.n34 163.367
R1485 B.n35 B.n34 163.367
R1486 B.n36 B.n35 163.367
R1487 B.n1265 B.n36 163.367
R1488 B.n1265 B.n41 163.367
R1489 B.n42 B.n41 163.367
R1490 B.n43 B.n42 163.367
R1491 B.n1270 B.n43 163.367
R1492 B.n1270 B.n48 163.367
R1493 B.n49 B.n48 163.367
R1494 B.n50 B.n49 163.367
R1495 B.n1275 B.n50 163.367
R1496 B.n1275 B.n55 163.367
R1497 B.n56 B.n55 163.367
R1498 B.n57 B.n56 163.367
R1499 B.n1280 B.n57 163.367
R1500 B.n1280 B.n62 163.367
R1501 B.n63 B.n62 163.367
R1502 B.n64 B.n63 163.367
R1503 B.n1285 B.n64 163.367
R1504 B.n1285 B.n69 163.367
R1505 B.n70 B.n69 163.367
R1506 B.n71 B.n70 163.367
R1507 B.n1290 B.n71 163.367
R1508 B.n1290 B.n76 163.367
R1509 B.n77 B.n76 163.367
R1510 B.n78 B.n77 163.367
R1511 B.n1295 B.n78 163.367
R1512 B.n1295 B.n83 163.367
R1513 B.n84 B.n83 163.367
R1514 B.n85 B.n84 163.367
R1515 B.n1300 B.n85 163.367
R1516 B.n1300 B.n90 163.367
R1517 B.n91 B.n90 163.367
R1518 B.n92 B.n91 163.367
R1519 B.n1305 B.n92 163.367
R1520 B.n1305 B.n97 163.367
R1521 B.n98 B.n97 163.367
R1522 B.n99 B.n98 163.367
R1523 B.n1310 B.n99 163.367
R1524 B.n1310 B.n104 163.367
R1525 B.n105 B.n104 163.367
R1526 B.n106 B.n105 163.367
R1527 B.n1315 B.n106 163.367
R1528 B.n1315 B.n111 163.367
R1529 B.n112 B.n111 163.367
R1530 B.n113 B.n112 163.367
R1531 B.n1320 B.n113 163.367
R1532 B.n1320 B.n118 163.367
R1533 B.n119 B.n118 163.367
R1534 B.n120 B.n119 163.367
R1535 B.n1325 B.n120 163.367
R1536 B.n1325 B.n125 163.367
R1537 B.n126 B.n125 163.367
R1538 B.n127 B.n126 163.367
R1539 B.n1330 B.n127 163.367
R1540 B.n1330 B.n132 163.367
R1541 B.n133 B.n132 163.367
R1542 B.n134 B.n133 163.367
R1543 B.n1335 B.n134 163.367
R1544 B.n1335 B.n139 163.367
R1545 B.n140 B.n139 163.367
R1546 B.n141 B.n140 163.367
R1547 B.n1340 B.n141 163.367
R1548 B.n1340 B.n146 163.367
R1549 B.n147 B.n146 163.367
R1550 B.n148 B.n147 163.367
R1551 B.n219 B.n148 163.367
R1552 B.n987 B.n652 163.367
R1553 B.n987 B.n719 163.367
R1554 B.n983 B.n982 163.367
R1555 B.n979 B.n978 163.367
R1556 B.n975 B.n974 163.367
R1557 B.n971 B.n970 163.367
R1558 B.n967 B.n966 163.367
R1559 B.n963 B.n962 163.367
R1560 B.n959 B.n958 163.367
R1561 B.n955 B.n954 163.367
R1562 B.n951 B.n950 163.367
R1563 B.n947 B.n946 163.367
R1564 B.n943 B.n942 163.367
R1565 B.n939 B.n938 163.367
R1566 B.n935 B.n934 163.367
R1567 B.n931 B.n930 163.367
R1568 B.n927 B.n926 163.367
R1569 B.n923 B.n922 163.367
R1570 B.n919 B.n918 163.367
R1571 B.n915 B.n914 163.367
R1572 B.n911 B.n910 163.367
R1573 B.n907 B.n906 163.367
R1574 B.n903 B.n902 163.367
R1575 B.n899 B.n898 163.367
R1576 B.n895 B.n894 163.367
R1577 B.n891 B.n890 163.367
R1578 B.n887 B.n886 163.367
R1579 B.n883 B.n882 163.367
R1580 B.n879 B.n878 163.367
R1581 B.n875 B.n874 163.367
R1582 B.n871 B.n870 163.367
R1583 B.n866 B.n865 163.367
R1584 B.n862 B.n861 163.367
R1585 B.n858 B.n857 163.367
R1586 B.n854 B.n853 163.367
R1587 B.n850 B.n849 163.367
R1588 B.n845 B.n844 163.367
R1589 B.n841 B.n840 163.367
R1590 B.n837 B.n836 163.367
R1591 B.n833 B.n832 163.367
R1592 B.n829 B.n828 163.367
R1593 B.n825 B.n824 163.367
R1594 B.n821 B.n820 163.367
R1595 B.n817 B.n816 163.367
R1596 B.n813 B.n812 163.367
R1597 B.n809 B.n808 163.367
R1598 B.n805 B.n804 163.367
R1599 B.n801 B.n800 163.367
R1600 B.n797 B.n796 163.367
R1601 B.n793 B.n792 163.367
R1602 B.n789 B.n788 163.367
R1603 B.n785 B.n784 163.367
R1604 B.n781 B.n780 163.367
R1605 B.n777 B.n776 163.367
R1606 B.n773 B.n772 163.367
R1607 B.n769 B.n768 163.367
R1608 B.n765 B.n764 163.367
R1609 B.n761 B.n760 163.367
R1610 B.n757 B.n756 163.367
R1611 B.n753 B.n752 163.367
R1612 B.n749 B.n748 163.367
R1613 B.n745 B.n744 163.367
R1614 B.n741 B.n740 163.367
R1615 B.n737 B.n736 163.367
R1616 B.n733 B.n732 163.367
R1617 B.n729 B.n728 163.367
R1618 B.n725 B.n718 163.367
R1619 B.n994 B.n650 163.367
R1620 B.n994 B.n644 163.367
R1621 B.n1002 B.n644 163.367
R1622 B.n1002 B.n642 163.367
R1623 B.n1006 B.n642 163.367
R1624 B.n1006 B.n636 163.367
R1625 B.n1014 B.n636 163.367
R1626 B.n1014 B.n634 163.367
R1627 B.n1018 B.n634 163.367
R1628 B.n1018 B.n628 163.367
R1629 B.n1026 B.n628 163.367
R1630 B.n1026 B.n626 163.367
R1631 B.n1030 B.n626 163.367
R1632 B.n1030 B.n620 163.367
R1633 B.n1038 B.n620 163.367
R1634 B.n1038 B.n618 163.367
R1635 B.n1042 B.n618 163.367
R1636 B.n1042 B.n612 163.367
R1637 B.n1050 B.n612 163.367
R1638 B.n1050 B.n610 163.367
R1639 B.n1054 B.n610 163.367
R1640 B.n1054 B.n604 163.367
R1641 B.n1062 B.n604 163.367
R1642 B.n1062 B.n602 163.367
R1643 B.n1066 B.n602 163.367
R1644 B.n1066 B.n596 163.367
R1645 B.n1074 B.n596 163.367
R1646 B.n1074 B.n594 163.367
R1647 B.n1078 B.n594 163.367
R1648 B.n1078 B.n588 163.367
R1649 B.n1086 B.n588 163.367
R1650 B.n1086 B.n586 163.367
R1651 B.n1090 B.n586 163.367
R1652 B.n1090 B.n580 163.367
R1653 B.n1098 B.n580 163.367
R1654 B.n1098 B.n578 163.367
R1655 B.n1102 B.n578 163.367
R1656 B.n1102 B.n572 163.367
R1657 B.n1110 B.n572 163.367
R1658 B.n1110 B.n570 163.367
R1659 B.n1114 B.n570 163.367
R1660 B.n1114 B.n564 163.367
R1661 B.n1122 B.n564 163.367
R1662 B.n1122 B.n562 163.367
R1663 B.n1126 B.n562 163.367
R1664 B.n1126 B.n556 163.367
R1665 B.n1134 B.n556 163.367
R1666 B.n1134 B.n554 163.367
R1667 B.n1138 B.n554 163.367
R1668 B.n1138 B.n548 163.367
R1669 B.n1146 B.n548 163.367
R1670 B.n1146 B.n546 163.367
R1671 B.n1150 B.n546 163.367
R1672 B.n1150 B.n540 163.367
R1673 B.n1158 B.n540 163.367
R1674 B.n1158 B.n538 163.367
R1675 B.n1162 B.n538 163.367
R1676 B.n1162 B.n532 163.367
R1677 B.n1170 B.n532 163.367
R1678 B.n1170 B.n530 163.367
R1679 B.n1174 B.n530 163.367
R1680 B.n1174 B.n524 163.367
R1681 B.n1182 B.n524 163.367
R1682 B.n1182 B.n522 163.367
R1683 B.n1186 B.n522 163.367
R1684 B.n1186 B.n516 163.367
R1685 B.n1194 B.n516 163.367
R1686 B.n1194 B.n514 163.367
R1687 B.n1198 B.n514 163.367
R1688 B.n1198 B.n508 163.367
R1689 B.n1206 B.n508 163.367
R1690 B.n1206 B.n506 163.367
R1691 B.n1210 B.n506 163.367
R1692 B.n1210 B.n500 163.367
R1693 B.n1218 B.n500 163.367
R1694 B.n1218 B.n498 163.367
R1695 B.n1222 B.n498 163.367
R1696 B.n1222 B.n492 163.367
R1697 B.n1231 B.n492 163.367
R1698 B.n1231 B.n490 163.367
R1699 B.n1235 B.n490 163.367
R1700 B.n1235 B.n3 163.367
R1701 B.n1520 B.n3 163.367
R1702 B.n1516 B.n2 163.367
R1703 B.n1516 B.n1515 163.367
R1704 B.n1515 B.n9 163.367
R1705 B.n1511 B.n9 163.367
R1706 B.n1511 B.n11 163.367
R1707 B.n1507 B.n11 163.367
R1708 B.n1507 B.n17 163.367
R1709 B.n1503 B.n17 163.367
R1710 B.n1503 B.n19 163.367
R1711 B.n1499 B.n19 163.367
R1712 B.n1499 B.n24 163.367
R1713 B.n1495 B.n24 163.367
R1714 B.n1495 B.n26 163.367
R1715 B.n1491 B.n26 163.367
R1716 B.n1491 B.n31 163.367
R1717 B.n1487 B.n31 163.367
R1718 B.n1487 B.n33 163.367
R1719 B.n1483 B.n33 163.367
R1720 B.n1483 B.n38 163.367
R1721 B.n1479 B.n38 163.367
R1722 B.n1479 B.n40 163.367
R1723 B.n1475 B.n40 163.367
R1724 B.n1475 B.n45 163.367
R1725 B.n1471 B.n45 163.367
R1726 B.n1471 B.n47 163.367
R1727 B.n1467 B.n47 163.367
R1728 B.n1467 B.n52 163.367
R1729 B.n1463 B.n52 163.367
R1730 B.n1463 B.n54 163.367
R1731 B.n1459 B.n54 163.367
R1732 B.n1459 B.n59 163.367
R1733 B.n1455 B.n59 163.367
R1734 B.n1455 B.n61 163.367
R1735 B.n1451 B.n61 163.367
R1736 B.n1451 B.n66 163.367
R1737 B.n1447 B.n66 163.367
R1738 B.n1447 B.n68 163.367
R1739 B.n1443 B.n68 163.367
R1740 B.n1443 B.n73 163.367
R1741 B.n1439 B.n73 163.367
R1742 B.n1439 B.n75 163.367
R1743 B.n1435 B.n75 163.367
R1744 B.n1435 B.n80 163.367
R1745 B.n1431 B.n80 163.367
R1746 B.n1431 B.n82 163.367
R1747 B.n1427 B.n82 163.367
R1748 B.n1427 B.n87 163.367
R1749 B.n1423 B.n87 163.367
R1750 B.n1423 B.n89 163.367
R1751 B.n1419 B.n89 163.367
R1752 B.n1419 B.n94 163.367
R1753 B.n1415 B.n94 163.367
R1754 B.n1415 B.n96 163.367
R1755 B.n1411 B.n96 163.367
R1756 B.n1411 B.n101 163.367
R1757 B.n1407 B.n101 163.367
R1758 B.n1407 B.n103 163.367
R1759 B.n1403 B.n103 163.367
R1760 B.n1403 B.n108 163.367
R1761 B.n1399 B.n108 163.367
R1762 B.n1399 B.n110 163.367
R1763 B.n1395 B.n110 163.367
R1764 B.n1395 B.n115 163.367
R1765 B.n1391 B.n115 163.367
R1766 B.n1391 B.n117 163.367
R1767 B.n1387 B.n117 163.367
R1768 B.n1387 B.n122 163.367
R1769 B.n1383 B.n122 163.367
R1770 B.n1383 B.n124 163.367
R1771 B.n1379 B.n124 163.367
R1772 B.n1379 B.n129 163.367
R1773 B.n1375 B.n129 163.367
R1774 B.n1375 B.n131 163.367
R1775 B.n1371 B.n131 163.367
R1776 B.n1371 B.n136 163.367
R1777 B.n1367 B.n136 163.367
R1778 B.n1367 B.n138 163.367
R1779 B.n1363 B.n138 163.367
R1780 B.n1363 B.n143 163.367
R1781 B.n1359 B.n143 163.367
R1782 B.n1359 B.n145 163.367
R1783 B.n1355 B.n145 163.367
R1784 B.n1355 B.n150 163.367
R1785 B.n220 B.t12 150.583
R1786 B.n722 B.t9 150.583
R1787 B.n223 B.t15 150.556
R1788 B.n720 B.t19 150.556
R1789 B.n224 B.n223 82.8126
R1790 B.n221 B.n220 82.8126
R1791 B.n723 B.n722 82.8126
R1792 B.n721 B.n720 82.8126
R1793 B.n1351 B.n1350 71.676
R1794 B.n226 B.n153 71.676
R1795 B.n230 B.n154 71.676
R1796 B.n234 B.n155 71.676
R1797 B.n238 B.n156 71.676
R1798 B.n242 B.n157 71.676
R1799 B.n246 B.n158 71.676
R1800 B.n250 B.n159 71.676
R1801 B.n254 B.n160 71.676
R1802 B.n258 B.n161 71.676
R1803 B.n262 B.n162 71.676
R1804 B.n266 B.n163 71.676
R1805 B.n270 B.n164 71.676
R1806 B.n274 B.n165 71.676
R1807 B.n278 B.n166 71.676
R1808 B.n282 B.n167 71.676
R1809 B.n286 B.n168 71.676
R1810 B.n290 B.n169 71.676
R1811 B.n294 B.n170 71.676
R1812 B.n298 B.n171 71.676
R1813 B.n302 B.n172 71.676
R1814 B.n306 B.n173 71.676
R1815 B.n310 B.n174 71.676
R1816 B.n314 B.n175 71.676
R1817 B.n318 B.n176 71.676
R1818 B.n322 B.n177 71.676
R1819 B.n326 B.n178 71.676
R1820 B.n330 B.n179 71.676
R1821 B.n334 B.n180 71.676
R1822 B.n338 B.n181 71.676
R1823 B.n342 B.n182 71.676
R1824 B.n346 B.n183 71.676
R1825 B.n350 B.n184 71.676
R1826 B.n354 B.n185 71.676
R1827 B.n358 B.n186 71.676
R1828 B.n362 B.n187 71.676
R1829 B.n366 B.n188 71.676
R1830 B.n370 B.n189 71.676
R1831 B.n374 B.n190 71.676
R1832 B.n378 B.n191 71.676
R1833 B.n382 B.n192 71.676
R1834 B.n386 B.n193 71.676
R1835 B.n390 B.n194 71.676
R1836 B.n394 B.n195 71.676
R1837 B.n398 B.n196 71.676
R1838 B.n402 B.n197 71.676
R1839 B.n406 B.n198 71.676
R1840 B.n410 B.n199 71.676
R1841 B.n414 B.n200 71.676
R1842 B.n418 B.n201 71.676
R1843 B.n422 B.n202 71.676
R1844 B.n426 B.n203 71.676
R1845 B.n430 B.n204 71.676
R1846 B.n434 B.n205 71.676
R1847 B.n438 B.n206 71.676
R1848 B.n442 B.n207 71.676
R1849 B.n446 B.n208 71.676
R1850 B.n450 B.n209 71.676
R1851 B.n454 B.n210 71.676
R1852 B.n458 B.n211 71.676
R1853 B.n462 B.n212 71.676
R1854 B.n466 B.n213 71.676
R1855 B.n470 B.n214 71.676
R1856 B.n474 B.n215 71.676
R1857 B.n478 B.n216 71.676
R1858 B.n482 B.n217 71.676
R1859 B.n1348 B.n218 71.676
R1860 B.n1348 B.n1347 71.676
R1861 B.n484 B.n217 71.676
R1862 B.n481 B.n216 71.676
R1863 B.n477 B.n215 71.676
R1864 B.n473 B.n214 71.676
R1865 B.n469 B.n213 71.676
R1866 B.n465 B.n212 71.676
R1867 B.n461 B.n211 71.676
R1868 B.n457 B.n210 71.676
R1869 B.n453 B.n209 71.676
R1870 B.n449 B.n208 71.676
R1871 B.n445 B.n207 71.676
R1872 B.n441 B.n206 71.676
R1873 B.n437 B.n205 71.676
R1874 B.n433 B.n204 71.676
R1875 B.n429 B.n203 71.676
R1876 B.n425 B.n202 71.676
R1877 B.n421 B.n201 71.676
R1878 B.n417 B.n200 71.676
R1879 B.n413 B.n199 71.676
R1880 B.n409 B.n198 71.676
R1881 B.n405 B.n197 71.676
R1882 B.n401 B.n196 71.676
R1883 B.n397 B.n195 71.676
R1884 B.n393 B.n194 71.676
R1885 B.n389 B.n193 71.676
R1886 B.n385 B.n192 71.676
R1887 B.n381 B.n191 71.676
R1888 B.n377 B.n190 71.676
R1889 B.n373 B.n189 71.676
R1890 B.n369 B.n188 71.676
R1891 B.n365 B.n187 71.676
R1892 B.n361 B.n186 71.676
R1893 B.n357 B.n185 71.676
R1894 B.n353 B.n184 71.676
R1895 B.n349 B.n183 71.676
R1896 B.n345 B.n182 71.676
R1897 B.n341 B.n181 71.676
R1898 B.n337 B.n180 71.676
R1899 B.n333 B.n179 71.676
R1900 B.n329 B.n178 71.676
R1901 B.n325 B.n177 71.676
R1902 B.n321 B.n176 71.676
R1903 B.n317 B.n175 71.676
R1904 B.n313 B.n174 71.676
R1905 B.n309 B.n173 71.676
R1906 B.n305 B.n172 71.676
R1907 B.n301 B.n171 71.676
R1908 B.n297 B.n170 71.676
R1909 B.n293 B.n169 71.676
R1910 B.n289 B.n168 71.676
R1911 B.n285 B.n167 71.676
R1912 B.n281 B.n166 71.676
R1913 B.n277 B.n165 71.676
R1914 B.n273 B.n164 71.676
R1915 B.n269 B.n163 71.676
R1916 B.n265 B.n162 71.676
R1917 B.n261 B.n161 71.676
R1918 B.n257 B.n160 71.676
R1919 B.n253 B.n159 71.676
R1920 B.n249 B.n158 71.676
R1921 B.n245 B.n157 71.676
R1922 B.n241 B.n156 71.676
R1923 B.n237 B.n155 71.676
R1924 B.n233 B.n154 71.676
R1925 B.n229 B.n153 71.676
R1926 B.n1350 B.n152 71.676
R1927 B.n990 B.n989 71.676
R1928 B.n719 B.n653 71.676
R1929 B.n982 B.n654 71.676
R1930 B.n978 B.n655 71.676
R1931 B.n974 B.n656 71.676
R1932 B.n970 B.n657 71.676
R1933 B.n966 B.n658 71.676
R1934 B.n962 B.n659 71.676
R1935 B.n958 B.n660 71.676
R1936 B.n954 B.n661 71.676
R1937 B.n950 B.n662 71.676
R1938 B.n946 B.n663 71.676
R1939 B.n942 B.n664 71.676
R1940 B.n938 B.n665 71.676
R1941 B.n934 B.n666 71.676
R1942 B.n930 B.n667 71.676
R1943 B.n926 B.n668 71.676
R1944 B.n922 B.n669 71.676
R1945 B.n918 B.n670 71.676
R1946 B.n914 B.n671 71.676
R1947 B.n910 B.n672 71.676
R1948 B.n906 B.n673 71.676
R1949 B.n902 B.n674 71.676
R1950 B.n898 B.n675 71.676
R1951 B.n894 B.n676 71.676
R1952 B.n890 B.n677 71.676
R1953 B.n886 B.n678 71.676
R1954 B.n882 B.n679 71.676
R1955 B.n878 B.n680 71.676
R1956 B.n874 B.n681 71.676
R1957 B.n870 B.n682 71.676
R1958 B.n865 B.n683 71.676
R1959 B.n861 B.n684 71.676
R1960 B.n857 B.n685 71.676
R1961 B.n853 B.n686 71.676
R1962 B.n849 B.n687 71.676
R1963 B.n844 B.n688 71.676
R1964 B.n840 B.n689 71.676
R1965 B.n836 B.n690 71.676
R1966 B.n832 B.n691 71.676
R1967 B.n828 B.n692 71.676
R1968 B.n824 B.n693 71.676
R1969 B.n820 B.n694 71.676
R1970 B.n816 B.n695 71.676
R1971 B.n812 B.n696 71.676
R1972 B.n808 B.n697 71.676
R1973 B.n804 B.n698 71.676
R1974 B.n800 B.n699 71.676
R1975 B.n796 B.n700 71.676
R1976 B.n792 B.n701 71.676
R1977 B.n788 B.n702 71.676
R1978 B.n784 B.n703 71.676
R1979 B.n780 B.n704 71.676
R1980 B.n776 B.n705 71.676
R1981 B.n772 B.n706 71.676
R1982 B.n768 B.n707 71.676
R1983 B.n764 B.n708 71.676
R1984 B.n760 B.n709 71.676
R1985 B.n756 B.n710 71.676
R1986 B.n752 B.n711 71.676
R1987 B.n748 B.n712 71.676
R1988 B.n744 B.n713 71.676
R1989 B.n740 B.n714 71.676
R1990 B.n736 B.n715 71.676
R1991 B.n732 B.n716 71.676
R1992 B.n728 B.n717 71.676
R1993 B.n989 B.n652 71.676
R1994 B.n983 B.n653 71.676
R1995 B.n979 B.n654 71.676
R1996 B.n975 B.n655 71.676
R1997 B.n971 B.n656 71.676
R1998 B.n967 B.n657 71.676
R1999 B.n963 B.n658 71.676
R2000 B.n959 B.n659 71.676
R2001 B.n955 B.n660 71.676
R2002 B.n951 B.n661 71.676
R2003 B.n947 B.n662 71.676
R2004 B.n943 B.n663 71.676
R2005 B.n939 B.n664 71.676
R2006 B.n935 B.n665 71.676
R2007 B.n931 B.n666 71.676
R2008 B.n927 B.n667 71.676
R2009 B.n923 B.n668 71.676
R2010 B.n919 B.n669 71.676
R2011 B.n915 B.n670 71.676
R2012 B.n911 B.n671 71.676
R2013 B.n907 B.n672 71.676
R2014 B.n903 B.n673 71.676
R2015 B.n899 B.n674 71.676
R2016 B.n895 B.n675 71.676
R2017 B.n891 B.n676 71.676
R2018 B.n887 B.n677 71.676
R2019 B.n883 B.n678 71.676
R2020 B.n879 B.n679 71.676
R2021 B.n875 B.n680 71.676
R2022 B.n871 B.n681 71.676
R2023 B.n866 B.n682 71.676
R2024 B.n862 B.n683 71.676
R2025 B.n858 B.n684 71.676
R2026 B.n854 B.n685 71.676
R2027 B.n850 B.n686 71.676
R2028 B.n845 B.n687 71.676
R2029 B.n841 B.n688 71.676
R2030 B.n837 B.n689 71.676
R2031 B.n833 B.n690 71.676
R2032 B.n829 B.n691 71.676
R2033 B.n825 B.n692 71.676
R2034 B.n821 B.n693 71.676
R2035 B.n817 B.n694 71.676
R2036 B.n813 B.n695 71.676
R2037 B.n809 B.n696 71.676
R2038 B.n805 B.n697 71.676
R2039 B.n801 B.n698 71.676
R2040 B.n797 B.n699 71.676
R2041 B.n793 B.n700 71.676
R2042 B.n789 B.n701 71.676
R2043 B.n785 B.n702 71.676
R2044 B.n781 B.n703 71.676
R2045 B.n777 B.n704 71.676
R2046 B.n773 B.n705 71.676
R2047 B.n769 B.n706 71.676
R2048 B.n765 B.n707 71.676
R2049 B.n761 B.n708 71.676
R2050 B.n757 B.n709 71.676
R2051 B.n753 B.n710 71.676
R2052 B.n749 B.n711 71.676
R2053 B.n745 B.n712 71.676
R2054 B.n741 B.n713 71.676
R2055 B.n737 B.n714 71.676
R2056 B.n733 B.n715 71.676
R2057 B.n729 B.n716 71.676
R2058 B.n725 B.n717 71.676
R2059 B.n1521 B.n1520 71.676
R2060 B.n1521 B.n2 71.676
R2061 B.n221 B.t13 67.7705
R2062 B.n723 B.t8 67.7705
R2063 B.n224 B.t16 67.7448
R2064 B.n721 B.t18 67.7448
R2065 B.n225 B.n224 59.5399
R2066 B.n222 B.n221 59.5399
R2067 B.n847 B.n723 59.5399
R2068 B.n868 B.n721 59.5399
R2069 B.n988 B.n649 54.6729
R2070 B.n1349 B.n149 54.6729
R2071 B.n992 B.n991 34.1859
R2072 B.n724 B.n647 34.1859
R2073 B.n1346 B.n1345 34.1859
R2074 B.n1353 B.n1352 34.1859
R2075 B.n995 B.n649 30.7255
R2076 B.n995 B.n645 30.7255
R2077 B.n1001 B.n645 30.7255
R2078 B.n1001 B.n641 30.7255
R2079 B.n1007 B.n641 30.7255
R2080 B.n1007 B.n637 30.7255
R2081 B.n1013 B.n637 30.7255
R2082 B.n1013 B.n633 30.7255
R2083 B.n1019 B.n633 30.7255
R2084 B.n1025 B.n629 30.7255
R2085 B.n1025 B.n625 30.7255
R2086 B.n1031 B.n625 30.7255
R2087 B.n1031 B.n621 30.7255
R2088 B.n1037 B.n621 30.7255
R2089 B.n1037 B.n617 30.7255
R2090 B.n1043 B.n617 30.7255
R2091 B.n1043 B.n613 30.7255
R2092 B.n1049 B.n613 30.7255
R2093 B.n1049 B.n609 30.7255
R2094 B.n1055 B.n609 30.7255
R2095 B.n1055 B.n605 30.7255
R2096 B.n1061 B.n605 30.7255
R2097 B.n1061 B.n601 30.7255
R2098 B.n1067 B.n601 30.7255
R2099 B.n1073 B.n597 30.7255
R2100 B.n1073 B.n593 30.7255
R2101 B.n1079 B.n593 30.7255
R2102 B.n1079 B.n589 30.7255
R2103 B.n1085 B.n589 30.7255
R2104 B.n1085 B.n585 30.7255
R2105 B.n1091 B.n585 30.7255
R2106 B.n1091 B.n581 30.7255
R2107 B.n1097 B.n581 30.7255
R2108 B.n1097 B.n577 30.7255
R2109 B.n1103 B.n577 30.7255
R2110 B.n1109 B.n573 30.7255
R2111 B.n1109 B.n569 30.7255
R2112 B.n1115 B.n569 30.7255
R2113 B.n1115 B.n565 30.7255
R2114 B.n1121 B.n565 30.7255
R2115 B.n1121 B.n561 30.7255
R2116 B.n1127 B.n561 30.7255
R2117 B.n1127 B.n557 30.7255
R2118 B.n1133 B.n557 30.7255
R2119 B.n1133 B.n552 30.7255
R2120 B.n1139 B.n552 30.7255
R2121 B.n1139 B.n553 30.7255
R2122 B.n1145 B.n545 30.7255
R2123 B.n1151 B.n545 30.7255
R2124 B.n1151 B.n541 30.7255
R2125 B.n1157 B.n541 30.7255
R2126 B.n1157 B.n537 30.7255
R2127 B.n1163 B.n537 30.7255
R2128 B.n1163 B.n533 30.7255
R2129 B.n1169 B.n533 30.7255
R2130 B.n1169 B.n529 30.7255
R2131 B.n1175 B.n529 30.7255
R2132 B.n1175 B.n525 30.7255
R2133 B.n1181 B.n525 30.7255
R2134 B.n1187 B.n521 30.7255
R2135 B.n1187 B.n517 30.7255
R2136 B.n1193 B.n517 30.7255
R2137 B.n1193 B.n513 30.7255
R2138 B.n1199 B.n513 30.7255
R2139 B.n1199 B.n509 30.7255
R2140 B.n1205 B.n509 30.7255
R2141 B.n1205 B.n505 30.7255
R2142 B.n1211 B.n505 30.7255
R2143 B.n1211 B.n501 30.7255
R2144 B.n1217 B.n501 30.7255
R2145 B.n1223 B.n497 30.7255
R2146 B.n1223 B.n493 30.7255
R2147 B.n1230 B.n493 30.7255
R2148 B.n1230 B.n489 30.7255
R2149 B.n1236 B.n489 30.7255
R2150 B.n1236 B.n4 30.7255
R2151 B.n1519 B.n4 30.7255
R2152 B.n1519 B.n1518 30.7255
R2153 B.n1518 B.n1517 30.7255
R2154 B.n1517 B.n8 30.7255
R2155 B.n12 B.n8 30.7255
R2156 B.n1510 B.n12 30.7255
R2157 B.n1510 B.n1509 30.7255
R2158 B.n1509 B.n1508 30.7255
R2159 B.n1508 B.n16 30.7255
R2160 B.n1502 B.n1501 30.7255
R2161 B.n1501 B.n1500 30.7255
R2162 B.n1500 B.n23 30.7255
R2163 B.n1494 B.n23 30.7255
R2164 B.n1494 B.n1493 30.7255
R2165 B.n1493 B.n1492 30.7255
R2166 B.n1492 B.n30 30.7255
R2167 B.n1486 B.n30 30.7255
R2168 B.n1486 B.n1485 30.7255
R2169 B.n1485 B.n1484 30.7255
R2170 B.n1484 B.n37 30.7255
R2171 B.n1478 B.n1477 30.7255
R2172 B.n1477 B.n1476 30.7255
R2173 B.n1476 B.n44 30.7255
R2174 B.n1470 B.n44 30.7255
R2175 B.n1470 B.n1469 30.7255
R2176 B.n1469 B.n1468 30.7255
R2177 B.n1468 B.n51 30.7255
R2178 B.n1462 B.n51 30.7255
R2179 B.n1462 B.n1461 30.7255
R2180 B.n1461 B.n1460 30.7255
R2181 B.n1460 B.n58 30.7255
R2182 B.n1454 B.n58 30.7255
R2183 B.n1453 B.n1452 30.7255
R2184 B.n1452 B.n65 30.7255
R2185 B.n1446 B.n65 30.7255
R2186 B.n1446 B.n1445 30.7255
R2187 B.n1445 B.n1444 30.7255
R2188 B.n1444 B.n72 30.7255
R2189 B.n1438 B.n72 30.7255
R2190 B.n1438 B.n1437 30.7255
R2191 B.n1437 B.n1436 30.7255
R2192 B.n1436 B.n79 30.7255
R2193 B.n1430 B.n79 30.7255
R2194 B.n1430 B.n1429 30.7255
R2195 B.n1428 B.n86 30.7255
R2196 B.n1422 B.n86 30.7255
R2197 B.n1422 B.n1421 30.7255
R2198 B.n1421 B.n1420 30.7255
R2199 B.n1420 B.n93 30.7255
R2200 B.n1414 B.n93 30.7255
R2201 B.n1414 B.n1413 30.7255
R2202 B.n1413 B.n1412 30.7255
R2203 B.n1412 B.n100 30.7255
R2204 B.n1406 B.n100 30.7255
R2205 B.n1406 B.n1405 30.7255
R2206 B.n1404 B.n107 30.7255
R2207 B.n1398 B.n107 30.7255
R2208 B.n1398 B.n1397 30.7255
R2209 B.n1397 B.n1396 30.7255
R2210 B.n1396 B.n114 30.7255
R2211 B.n1390 B.n114 30.7255
R2212 B.n1390 B.n1389 30.7255
R2213 B.n1389 B.n1388 30.7255
R2214 B.n1388 B.n121 30.7255
R2215 B.n1382 B.n121 30.7255
R2216 B.n1382 B.n1381 30.7255
R2217 B.n1381 B.n1380 30.7255
R2218 B.n1380 B.n128 30.7255
R2219 B.n1374 B.n128 30.7255
R2220 B.n1374 B.n1373 30.7255
R2221 B.n1372 B.n135 30.7255
R2222 B.n1366 B.n135 30.7255
R2223 B.n1366 B.n1365 30.7255
R2224 B.n1365 B.n1364 30.7255
R2225 B.n1364 B.n142 30.7255
R2226 B.n1358 B.n142 30.7255
R2227 B.n1358 B.n1357 30.7255
R2228 B.n1357 B.n1356 30.7255
R2229 B.n1356 B.n149 30.7255
R2230 B.n1103 B.t22 28.9181
R2231 B.t1 B.n521 28.9181
R2232 B.t5 B.n37 28.9181
R2233 B.t21 B.n1428 28.9181
R2234 B.n1019 B.t7 18.9777
R2235 B.t2 B.n597 18.9777
R2236 B.n1217 B.t20 18.9777
R2237 B.n1502 B.t3 18.9777
R2238 B.n1405 B.t0 18.9777
R2239 B.t11 B.n1372 18.9777
R2240 B B.n1522 18.0485
R2241 B.n553 B.t23 15.363
R2242 B.n1145 B.t23 15.363
R2243 B.n1454 B.t4 15.363
R2244 B.t4 B.n1453 15.363
R2245 B.t7 B.n629 11.7483
R2246 B.n1067 B.t2 11.7483
R2247 B.t20 B.n497 11.7483
R2248 B.t3 B.n16 11.7483
R2249 B.t0 B.n1404 11.7483
R2250 B.n1373 B.t11 11.7483
R2251 B.n993 B.n992 10.6151
R2252 B.n993 B.n643 10.6151
R2253 B.n1003 B.n643 10.6151
R2254 B.n1004 B.n1003 10.6151
R2255 B.n1005 B.n1004 10.6151
R2256 B.n1005 B.n635 10.6151
R2257 B.n1015 B.n635 10.6151
R2258 B.n1016 B.n1015 10.6151
R2259 B.n1017 B.n1016 10.6151
R2260 B.n1017 B.n627 10.6151
R2261 B.n1027 B.n627 10.6151
R2262 B.n1028 B.n1027 10.6151
R2263 B.n1029 B.n1028 10.6151
R2264 B.n1029 B.n619 10.6151
R2265 B.n1039 B.n619 10.6151
R2266 B.n1040 B.n1039 10.6151
R2267 B.n1041 B.n1040 10.6151
R2268 B.n1041 B.n611 10.6151
R2269 B.n1051 B.n611 10.6151
R2270 B.n1052 B.n1051 10.6151
R2271 B.n1053 B.n1052 10.6151
R2272 B.n1053 B.n603 10.6151
R2273 B.n1063 B.n603 10.6151
R2274 B.n1064 B.n1063 10.6151
R2275 B.n1065 B.n1064 10.6151
R2276 B.n1065 B.n595 10.6151
R2277 B.n1075 B.n595 10.6151
R2278 B.n1076 B.n1075 10.6151
R2279 B.n1077 B.n1076 10.6151
R2280 B.n1077 B.n587 10.6151
R2281 B.n1087 B.n587 10.6151
R2282 B.n1088 B.n1087 10.6151
R2283 B.n1089 B.n1088 10.6151
R2284 B.n1089 B.n579 10.6151
R2285 B.n1099 B.n579 10.6151
R2286 B.n1100 B.n1099 10.6151
R2287 B.n1101 B.n1100 10.6151
R2288 B.n1101 B.n571 10.6151
R2289 B.n1111 B.n571 10.6151
R2290 B.n1112 B.n1111 10.6151
R2291 B.n1113 B.n1112 10.6151
R2292 B.n1113 B.n563 10.6151
R2293 B.n1123 B.n563 10.6151
R2294 B.n1124 B.n1123 10.6151
R2295 B.n1125 B.n1124 10.6151
R2296 B.n1125 B.n555 10.6151
R2297 B.n1135 B.n555 10.6151
R2298 B.n1136 B.n1135 10.6151
R2299 B.n1137 B.n1136 10.6151
R2300 B.n1137 B.n547 10.6151
R2301 B.n1147 B.n547 10.6151
R2302 B.n1148 B.n1147 10.6151
R2303 B.n1149 B.n1148 10.6151
R2304 B.n1149 B.n539 10.6151
R2305 B.n1159 B.n539 10.6151
R2306 B.n1160 B.n1159 10.6151
R2307 B.n1161 B.n1160 10.6151
R2308 B.n1161 B.n531 10.6151
R2309 B.n1171 B.n531 10.6151
R2310 B.n1172 B.n1171 10.6151
R2311 B.n1173 B.n1172 10.6151
R2312 B.n1173 B.n523 10.6151
R2313 B.n1183 B.n523 10.6151
R2314 B.n1184 B.n1183 10.6151
R2315 B.n1185 B.n1184 10.6151
R2316 B.n1185 B.n515 10.6151
R2317 B.n1195 B.n515 10.6151
R2318 B.n1196 B.n1195 10.6151
R2319 B.n1197 B.n1196 10.6151
R2320 B.n1197 B.n507 10.6151
R2321 B.n1207 B.n507 10.6151
R2322 B.n1208 B.n1207 10.6151
R2323 B.n1209 B.n1208 10.6151
R2324 B.n1209 B.n499 10.6151
R2325 B.n1219 B.n499 10.6151
R2326 B.n1220 B.n1219 10.6151
R2327 B.n1221 B.n1220 10.6151
R2328 B.n1221 B.n491 10.6151
R2329 B.n1232 B.n491 10.6151
R2330 B.n1233 B.n1232 10.6151
R2331 B.n1234 B.n1233 10.6151
R2332 B.n1234 B.n0 10.6151
R2333 B.n991 B.n651 10.6151
R2334 B.n986 B.n651 10.6151
R2335 B.n986 B.n985 10.6151
R2336 B.n985 B.n984 10.6151
R2337 B.n984 B.n981 10.6151
R2338 B.n981 B.n980 10.6151
R2339 B.n980 B.n977 10.6151
R2340 B.n977 B.n976 10.6151
R2341 B.n976 B.n973 10.6151
R2342 B.n973 B.n972 10.6151
R2343 B.n972 B.n969 10.6151
R2344 B.n969 B.n968 10.6151
R2345 B.n968 B.n965 10.6151
R2346 B.n965 B.n964 10.6151
R2347 B.n964 B.n961 10.6151
R2348 B.n961 B.n960 10.6151
R2349 B.n960 B.n957 10.6151
R2350 B.n957 B.n956 10.6151
R2351 B.n956 B.n953 10.6151
R2352 B.n953 B.n952 10.6151
R2353 B.n952 B.n949 10.6151
R2354 B.n949 B.n948 10.6151
R2355 B.n948 B.n945 10.6151
R2356 B.n945 B.n944 10.6151
R2357 B.n944 B.n941 10.6151
R2358 B.n941 B.n940 10.6151
R2359 B.n940 B.n937 10.6151
R2360 B.n937 B.n936 10.6151
R2361 B.n936 B.n933 10.6151
R2362 B.n933 B.n932 10.6151
R2363 B.n932 B.n929 10.6151
R2364 B.n929 B.n928 10.6151
R2365 B.n928 B.n925 10.6151
R2366 B.n925 B.n924 10.6151
R2367 B.n924 B.n921 10.6151
R2368 B.n921 B.n920 10.6151
R2369 B.n920 B.n917 10.6151
R2370 B.n917 B.n916 10.6151
R2371 B.n916 B.n913 10.6151
R2372 B.n913 B.n912 10.6151
R2373 B.n912 B.n909 10.6151
R2374 B.n909 B.n908 10.6151
R2375 B.n908 B.n905 10.6151
R2376 B.n905 B.n904 10.6151
R2377 B.n904 B.n901 10.6151
R2378 B.n901 B.n900 10.6151
R2379 B.n900 B.n897 10.6151
R2380 B.n897 B.n896 10.6151
R2381 B.n896 B.n893 10.6151
R2382 B.n893 B.n892 10.6151
R2383 B.n892 B.n889 10.6151
R2384 B.n889 B.n888 10.6151
R2385 B.n888 B.n885 10.6151
R2386 B.n885 B.n884 10.6151
R2387 B.n884 B.n881 10.6151
R2388 B.n881 B.n880 10.6151
R2389 B.n880 B.n877 10.6151
R2390 B.n877 B.n876 10.6151
R2391 B.n876 B.n873 10.6151
R2392 B.n873 B.n872 10.6151
R2393 B.n872 B.n869 10.6151
R2394 B.n867 B.n864 10.6151
R2395 B.n864 B.n863 10.6151
R2396 B.n863 B.n860 10.6151
R2397 B.n860 B.n859 10.6151
R2398 B.n859 B.n856 10.6151
R2399 B.n856 B.n855 10.6151
R2400 B.n855 B.n852 10.6151
R2401 B.n852 B.n851 10.6151
R2402 B.n851 B.n848 10.6151
R2403 B.n846 B.n843 10.6151
R2404 B.n843 B.n842 10.6151
R2405 B.n842 B.n839 10.6151
R2406 B.n839 B.n838 10.6151
R2407 B.n838 B.n835 10.6151
R2408 B.n835 B.n834 10.6151
R2409 B.n834 B.n831 10.6151
R2410 B.n831 B.n830 10.6151
R2411 B.n830 B.n827 10.6151
R2412 B.n827 B.n826 10.6151
R2413 B.n826 B.n823 10.6151
R2414 B.n823 B.n822 10.6151
R2415 B.n822 B.n819 10.6151
R2416 B.n819 B.n818 10.6151
R2417 B.n818 B.n815 10.6151
R2418 B.n815 B.n814 10.6151
R2419 B.n814 B.n811 10.6151
R2420 B.n811 B.n810 10.6151
R2421 B.n810 B.n807 10.6151
R2422 B.n807 B.n806 10.6151
R2423 B.n806 B.n803 10.6151
R2424 B.n803 B.n802 10.6151
R2425 B.n802 B.n799 10.6151
R2426 B.n799 B.n798 10.6151
R2427 B.n798 B.n795 10.6151
R2428 B.n795 B.n794 10.6151
R2429 B.n794 B.n791 10.6151
R2430 B.n791 B.n790 10.6151
R2431 B.n790 B.n787 10.6151
R2432 B.n787 B.n786 10.6151
R2433 B.n786 B.n783 10.6151
R2434 B.n783 B.n782 10.6151
R2435 B.n782 B.n779 10.6151
R2436 B.n779 B.n778 10.6151
R2437 B.n778 B.n775 10.6151
R2438 B.n775 B.n774 10.6151
R2439 B.n774 B.n771 10.6151
R2440 B.n771 B.n770 10.6151
R2441 B.n770 B.n767 10.6151
R2442 B.n767 B.n766 10.6151
R2443 B.n766 B.n763 10.6151
R2444 B.n763 B.n762 10.6151
R2445 B.n762 B.n759 10.6151
R2446 B.n759 B.n758 10.6151
R2447 B.n758 B.n755 10.6151
R2448 B.n755 B.n754 10.6151
R2449 B.n754 B.n751 10.6151
R2450 B.n751 B.n750 10.6151
R2451 B.n750 B.n747 10.6151
R2452 B.n747 B.n746 10.6151
R2453 B.n746 B.n743 10.6151
R2454 B.n743 B.n742 10.6151
R2455 B.n742 B.n739 10.6151
R2456 B.n739 B.n738 10.6151
R2457 B.n738 B.n735 10.6151
R2458 B.n735 B.n734 10.6151
R2459 B.n734 B.n731 10.6151
R2460 B.n731 B.n730 10.6151
R2461 B.n730 B.n727 10.6151
R2462 B.n727 B.n726 10.6151
R2463 B.n726 B.n724 10.6151
R2464 B.n997 B.n647 10.6151
R2465 B.n998 B.n997 10.6151
R2466 B.n999 B.n998 10.6151
R2467 B.n999 B.n639 10.6151
R2468 B.n1009 B.n639 10.6151
R2469 B.n1010 B.n1009 10.6151
R2470 B.n1011 B.n1010 10.6151
R2471 B.n1011 B.n631 10.6151
R2472 B.n1021 B.n631 10.6151
R2473 B.n1022 B.n1021 10.6151
R2474 B.n1023 B.n1022 10.6151
R2475 B.n1023 B.n623 10.6151
R2476 B.n1033 B.n623 10.6151
R2477 B.n1034 B.n1033 10.6151
R2478 B.n1035 B.n1034 10.6151
R2479 B.n1035 B.n615 10.6151
R2480 B.n1045 B.n615 10.6151
R2481 B.n1046 B.n1045 10.6151
R2482 B.n1047 B.n1046 10.6151
R2483 B.n1047 B.n607 10.6151
R2484 B.n1057 B.n607 10.6151
R2485 B.n1058 B.n1057 10.6151
R2486 B.n1059 B.n1058 10.6151
R2487 B.n1059 B.n599 10.6151
R2488 B.n1069 B.n599 10.6151
R2489 B.n1070 B.n1069 10.6151
R2490 B.n1071 B.n1070 10.6151
R2491 B.n1071 B.n591 10.6151
R2492 B.n1081 B.n591 10.6151
R2493 B.n1082 B.n1081 10.6151
R2494 B.n1083 B.n1082 10.6151
R2495 B.n1083 B.n583 10.6151
R2496 B.n1093 B.n583 10.6151
R2497 B.n1094 B.n1093 10.6151
R2498 B.n1095 B.n1094 10.6151
R2499 B.n1095 B.n575 10.6151
R2500 B.n1105 B.n575 10.6151
R2501 B.n1106 B.n1105 10.6151
R2502 B.n1107 B.n1106 10.6151
R2503 B.n1107 B.n567 10.6151
R2504 B.n1117 B.n567 10.6151
R2505 B.n1118 B.n1117 10.6151
R2506 B.n1119 B.n1118 10.6151
R2507 B.n1119 B.n559 10.6151
R2508 B.n1129 B.n559 10.6151
R2509 B.n1130 B.n1129 10.6151
R2510 B.n1131 B.n1130 10.6151
R2511 B.n1131 B.n550 10.6151
R2512 B.n1141 B.n550 10.6151
R2513 B.n1142 B.n1141 10.6151
R2514 B.n1143 B.n1142 10.6151
R2515 B.n1143 B.n543 10.6151
R2516 B.n1153 B.n543 10.6151
R2517 B.n1154 B.n1153 10.6151
R2518 B.n1155 B.n1154 10.6151
R2519 B.n1155 B.n535 10.6151
R2520 B.n1165 B.n535 10.6151
R2521 B.n1166 B.n1165 10.6151
R2522 B.n1167 B.n1166 10.6151
R2523 B.n1167 B.n527 10.6151
R2524 B.n1177 B.n527 10.6151
R2525 B.n1178 B.n1177 10.6151
R2526 B.n1179 B.n1178 10.6151
R2527 B.n1179 B.n519 10.6151
R2528 B.n1189 B.n519 10.6151
R2529 B.n1190 B.n1189 10.6151
R2530 B.n1191 B.n1190 10.6151
R2531 B.n1191 B.n511 10.6151
R2532 B.n1201 B.n511 10.6151
R2533 B.n1202 B.n1201 10.6151
R2534 B.n1203 B.n1202 10.6151
R2535 B.n1203 B.n503 10.6151
R2536 B.n1213 B.n503 10.6151
R2537 B.n1214 B.n1213 10.6151
R2538 B.n1215 B.n1214 10.6151
R2539 B.n1215 B.n495 10.6151
R2540 B.n1225 B.n495 10.6151
R2541 B.n1226 B.n1225 10.6151
R2542 B.n1228 B.n1226 10.6151
R2543 B.n1228 B.n1227 10.6151
R2544 B.n1227 B.n487 10.6151
R2545 B.n1239 B.n487 10.6151
R2546 B.n1240 B.n1239 10.6151
R2547 B.n1241 B.n1240 10.6151
R2548 B.n1242 B.n1241 10.6151
R2549 B.n1243 B.n1242 10.6151
R2550 B.n1246 B.n1243 10.6151
R2551 B.n1247 B.n1246 10.6151
R2552 B.n1248 B.n1247 10.6151
R2553 B.n1249 B.n1248 10.6151
R2554 B.n1251 B.n1249 10.6151
R2555 B.n1252 B.n1251 10.6151
R2556 B.n1253 B.n1252 10.6151
R2557 B.n1254 B.n1253 10.6151
R2558 B.n1256 B.n1254 10.6151
R2559 B.n1257 B.n1256 10.6151
R2560 B.n1258 B.n1257 10.6151
R2561 B.n1259 B.n1258 10.6151
R2562 B.n1261 B.n1259 10.6151
R2563 B.n1262 B.n1261 10.6151
R2564 B.n1263 B.n1262 10.6151
R2565 B.n1264 B.n1263 10.6151
R2566 B.n1266 B.n1264 10.6151
R2567 B.n1267 B.n1266 10.6151
R2568 B.n1268 B.n1267 10.6151
R2569 B.n1269 B.n1268 10.6151
R2570 B.n1271 B.n1269 10.6151
R2571 B.n1272 B.n1271 10.6151
R2572 B.n1273 B.n1272 10.6151
R2573 B.n1274 B.n1273 10.6151
R2574 B.n1276 B.n1274 10.6151
R2575 B.n1277 B.n1276 10.6151
R2576 B.n1278 B.n1277 10.6151
R2577 B.n1279 B.n1278 10.6151
R2578 B.n1281 B.n1279 10.6151
R2579 B.n1282 B.n1281 10.6151
R2580 B.n1283 B.n1282 10.6151
R2581 B.n1284 B.n1283 10.6151
R2582 B.n1286 B.n1284 10.6151
R2583 B.n1287 B.n1286 10.6151
R2584 B.n1288 B.n1287 10.6151
R2585 B.n1289 B.n1288 10.6151
R2586 B.n1291 B.n1289 10.6151
R2587 B.n1292 B.n1291 10.6151
R2588 B.n1293 B.n1292 10.6151
R2589 B.n1294 B.n1293 10.6151
R2590 B.n1296 B.n1294 10.6151
R2591 B.n1297 B.n1296 10.6151
R2592 B.n1298 B.n1297 10.6151
R2593 B.n1299 B.n1298 10.6151
R2594 B.n1301 B.n1299 10.6151
R2595 B.n1302 B.n1301 10.6151
R2596 B.n1303 B.n1302 10.6151
R2597 B.n1304 B.n1303 10.6151
R2598 B.n1306 B.n1304 10.6151
R2599 B.n1307 B.n1306 10.6151
R2600 B.n1308 B.n1307 10.6151
R2601 B.n1309 B.n1308 10.6151
R2602 B.n1311 B.n1309 10.6151
R2603 B.n1312 B.n1311 10.6151
R2604 B.n1313 B.n1312 10.6151
R2605 B.n1314 B.n1313 10.6151
R2606 B.n1316 B.n1314 10.6151
R2607 B.n1317 B.n1316 10.6151
R2608 B.n1318 B.n1317 10.6151
R2609 B.n1319 B.n1318 10.6151
R2610 B.n1321 B.n1319 10.6151
R2611 B.n1322 B.n1321 10.6151
R2612 B.n1323 B.n1322 10.6151
R2613 B.n1324 B.n1323 10.6151
R2614 B.n1326 B.n1324 10.6151
R2615 B.n1327 B.n1326 10.6151
R2616 B.n1328 B.n1327 10.6151
R2617 B.n1329 B.n1328 10.6151
R2618 B.n1331 B.n1329 10.6151
R2619 B.n1332 B.n1331 10.6151
R2620 B.n1333 B.n1332 10.6151
R2621 B.n1334 B.n1333 10.6151
R2622 B.n1336 B.n1334 10.6151
R2623 B.n1337 B.n1336 10.6151
R2624 B.n1338 B.n1337 10.6151
R2625 B.n1339 B.n1338 10.6151
R2626 B.n1341 B.n1339 10.6151
R2627 B.n1342 B.n1341 10.6151
R2628 B.n1343 B.n1342 10.6151
R2629 B.n1344 B.n1343 10.6151
R2630 B.n1345 B.n1344 10.6151
R2631 B.n1514 B.n1 10.6151
R2632 B.n1514 B.n1513 10.6151
R2633 B.n1513 B.n1512 10.6151
R2634 B.n1512 B.n10 10.6151
R2635 B.n1506 B.n10 10.6151
R2636 B.n1506 B.n1505 10.6151
R2637 B.n1505 B.n1504 10.6151
R2638 B.n1504 B.n18 10.6151
R2639 B.n1498 B.n18 10.6151
R2640 B.n1498 B.n1497 10.6151
R2641 B.n1497 B.n1496 10.6151
R2642 B.n1496 B.n25 10.6151
R2643 B.n1490 B.n25 10.6151
R2644 B.n1490 B.n1489 10.6151
R2645 B.n1489 B.n1488 10.6151
R2646 B.n1488 B.n32 10.6151
R2647 B.n1482 B.n32 10.6151
R2648 B.n1482 B.n1481 10.6151
R2649 B.n1481 B.n1480 10.6151
R2650 B.n1480 B.n39 10.6151
R2651 B.n1474 B.n39 10.6151
R2652 B.n1474 B.n1473 10.6151
R2653 B.n1473 B.n1472 10.6151
R2654 B.n1472 B.n46 10.6151
R2655 B.n1466 B.n46 10.6151
R2656 B.n1466 B.n1465 10.6151
R2657 B.n1465 B.n1464 10.6151
R2658 B.n1464 B.n53 10.6151
R2659 B.n1458 B.n53 10.6151
R2660 B.n1458 B.n1457 10.6151
R2661 B.n1457 B.n1456 10.6151
R2662 B.n1456 B.n60 10.6151
R2663 B.n1450 B.n60 10.6151
R2664 B.n1450 B.n1449 10.6151
R2665 B.n1449 B.n1448 10.6151
R2666 B.n1448 B.n67 10.6151
R2667 B.n1442 B.n67 10.6151
R2668 B.n1442 B.n1441 10.6151
R2669 B.n1441 B.n1440 10.6151
R2670 B.n1440 B.n74 10.6151
R2671 B.n1434 B.n74 10.6151
R2672 B.n1434 B.n1433 10.6151
R2673 B.n1433 B.n1432 10.6151
R2674 B.n1432 B.n81 10.6151
R2675 B.n1426 B.n81 10.6151
R2676 B.n1426 B.n1425 10.6151
R2677 B.n1425 B.n1424 10.6151
R2678 B.n1424 B.n88 10.6151
R2679 B.n1418 B.n88 10.6151
R2680 B.n1418 B.n1417 10.6151
R2681 B.n1417 B.n1416 10.6151
R2682 B.n1416 B.n95 10.6151
R2683 B.n1410 B.n95 10.6151
R2684 B.n1410 B.n1409 10.6151
R2685 B.n1409 B.n1408 10.6151
R2686 B.n1408 B.n102 10.6151
R2687 B.n1402 B.n102 10.6151
R2688 B.n1402 B.n1401 10.6151
R2689 B.n1401 B.n1400 10.6151
R2690 B.n1400 B.n109 10.6151
R2691 B.n1394 B.n109 10.6151
R2692 B.n1394 B.n1393 10.6151
R2693 B.n1393 B.n1392 10.6151
R2694 B.n1392 B.n116 10.6151
R2695 B.n1386 B.n116 10.6151
R2696 B.n1386 B.n1385 10.6151
R2697 B.n1385 B.n1384 10.6151
R2698 B.n1384 B.n123 10.6151
R2699 B.n1378 B.n123 10.6151
R2700 B.n1378 B.n1377 10.6151
R2701 B.n1377 B.n1376 10.6151
R2702 B.n1376 B.n130 10.6151
R2703 B.n1370 B.n130 10.6151
R2704 B.n1370 B.n1369 10.6151
R2705 B.n1369 B.n1368 10.6151
R2706 B.n1368 B.n137 10.6151
R2707 B.n1362 B.n137 10.6151
R2708 B.n1362 B.n1361 10.6151
R2709 B.n1361 B.n1360 10.6151
R2710 B.n1360 B.n144 10.6151
R2711 B.n1354 B.n144 10.6151
R2712 B.n1354 B.n1353 10.6151
R2713 B.n1352 B.n151 10.6151
R2714 B.n227 B.n151 10.6151
R2715 B.n228 B.n227 10.6151
R2716 B.n231 B.n228 10.6151
R2717 B.n232 B.n231 10.6151
R2718 B.n235 B.n232 10.6151
R2719 B.n236 B.n235 10.6151
R2720 B.n239 B.n236 10.6151
R2721 B.n240 B.n239 10.6151
R2722 B.n243 B.n240 10.6151
R2723 B.n244 B.n243 10.6151
R2724 B.n247 B.n244 10.6151
R2725 B.n248 B.n247 10.6151
R2726 B.n251 B.n248 10.6151
R2727 B.n252 B.n251 10.6151
R2728 B.n255 B.n252 10.6151
R2729 B.n256 B.n255 10.6151
R2730 B.n259 B.n256 10.6151
R2731 B.n260 B.n259 10.6151
R2732 B.n263 B.n260 10.6151
R2733 B.n264 B.n263 10.6151
R2734 B.n267 B.n264 10.6151
R2735 B.n268 B.n267 10.6151
R2736 B.n271 B.n268 10.6151
R2737 B.n272 B.n271 10.6151
R2738 B.n275 B.n272 10.6151
R2739 B.n276 B.n275 10.6151
R2740 B.n279 B.n276 10.6151
R2741 B.n280 B.n279 10.6151
R2742 B.n283 B.n280 10.6151
R2743 B.n284 B.n283 10.6151
R2744 B.n287 B.n284 10.6151
R2745 B.n288 B.n287 10.6151
R2746 B.n291 B.n288 10.6151
R2747 B.n292 B.n291 10.6151
R2748 B.n295 B.n292 10.6151
R2749 B.n296 B.n295 10.6151
R2750 B.n299 B.n296 10.6151
R2751 B.n300 B.n299 10.6151
R2752 B.n303 B.n300 10.6151
R2753 B.n304 B.n303 10.6151
R2754 B.n307 B.n304 10.6151
R2755 B.n308 B.n307 10.6151
R2756 B.n311 B.n308 10.6151
R2757 B.n312 B.n311 10.6151
R2758 B.n315 B.n312 10.6151
R2759 B.n316 B.n315 10.6151
R2760 B.n319 B.n316 10.6151
R2761 B.n320 B.n319 10.6151
R2762 B.n323 B.n320 10.6151
R2763 B.n324 B.n323 10.6151
R2764 B.n327 B.n324 10.6151
R2765 B.n328 B.n327 10.6151
R2766 B.n331 B.n328 10.6151
R2767 B.n332 B.n331 10.6151
R2768 B.n335 B.n332 10.6151
R2769 B.n336 B.n335 10.6151
R2770 B.n339 B.n336 10.6151
R2771 B.n340 B.n339 10.6151
R2772 B.n343 B.n340 10.6151
R2773 B.n344 B.n343 10.6151
R2774 B.n348 B.n347 10.6151
R2775 B.n351 B.n348 10.6151
R2776 B.n352 B.n351 10.6151
R2777 B.n355 B.n352 10.6151
R2778 B.n356 B.n355 10.6151
R2779 B.n359 B.n356 10.6151
R2780 B.n360 B.n359 10.6151
R2781 B.n363 B.n360 10.6151
R2782 B.n364 B.n363 10.6151
R2783 B.n368 B.n367 10.6151
R2784 B.n371 B.n368 10.6151
R2785 B.n372 B.n371 10.6151
R2786 B.n375 B.n372 10.6151
R2787 B.n376 B.n375 10.6151
R2788 B.n379 B.n376 10.6151
R2789 B.n380 B.n379 10.6151
R2790 B.n383 B.n380 10.6151
R2791 B.n384 B.n383 10.6151
R2792 B.n387 B.n384 10.6151
R2793 B.n388 B.n387 10.6151
R2794 B.n391 B.n388 10.6151
R2795 B.n392 B.n391 10.6151
R2796 B.n395 B.n392 10.6151
R2797 B.n396 B.n395 10.6151
R2798 B.n399 B.n396 10.6151
R2799 B.n400 B.n399 10.6151
R2800 B.n403 B.n400 10.6151
R2801 B.n404 B.n403 10.6151
R2802 B.n407 B.n404 10.6151
R2803 B.n408 B.n407 10.6151
R2804 B.n411 B.n408 10.6151
R2805 B.n412 B.n411 10.6151
R2806 B.n415 B.n412 10.6151
R2807 B.n416 B.n415 10.6151
R2808 B.n419 B.n416 10.6151
R2809 B.n420 B.n419 10.6151
R2810 B.n423 B.n420 10.6151
R2811 B.n424 B.n423 10.6151
R2812 B.n427 B.n424 10.6151
R2813 B.n428 B.n427 10.6151
R2814 B.n431 B.n428 10.6151
R2815 B.n432 B.n431 10.6151
R2816 B.n435 B.n432 10.6151
R2817 B.n436 B.n435 10.6151
R2818 B.n439 B.n436 10.6151
R2819 B.n440 B.n439 10.6151
R2820 B.n443 B.n440 10.6151
R2821 B.n444 B.n443 10.6151
R2822 B.n447 B.n444 10.6151
R2823 B.n448 B.n447 10.6151
R2824 B.n451 B.n448 10.6151
R2825 B.n452 B.n451 10.6151
R2826 B.n455 B.n452 10.6151
R2827 B.n456 B.n455 10.6151
R2828 B.n459 B.n456 10.6151
R2829 B.n460 B.n459 10.6151
R2830 B.n463 B.n460 10.6151
R2831 B.n464 B.n463 10.6151
R2832 B.n467 B.n464 10.6151
R2833 B.n468 B.n467 10.6151
R2834 B.n471 B.n468 10.6151
R2835 B.n472 B.n471 10.6151
R2836 B.n475 B.n472 10.6151
R2837 B.n476 B.n475 10.6151
R2838 B.n479 B.n476 10.6151
R2839 B.n480 B.n479 10.6151
R2840 B.n483 B.n480 10.6151
R2841 B.n485 B.n483 10.6151
R2842 B.n486 B.n485 10.6151
R2843 B.n1346 B.n486 10.6151
R2844 B.n869 B.n868 9.36635
R2845 B.n847 B.n846 9.36635
R2846 B.n344 B.n225 9.36635
R2847 B.n367 B.n222 9.36635
R2848 B.n1522 B.n0 8.11757
R2849 B.n1522 B.n1 8.11757
R2850 B.t22 B.n573 1.80785
R2851 B.n1181 B.t1 1.80785
R2852 B.n1478 B.t5 1.80785
R2853 B.n1429 B.t21 1.80785
R2854 B.n868 B.n867 1.24928
R2855 B.n848 B.n847 1.24928
R2856 B.n347 B.n225 1.24928
R2857 B.n364 B.n222 1.24928
R2858 VP.n35 VP.n32 161.3
R2859 VP.n37 VP.n36 161.3
R2860 VP.n38 VP.n31 161.3
R2861 VP.n40 VP.n39 161.3
R2862 VP.n41 VP.n30 161.3
R2863 VP.n43 VP.n42 161.3
R2864 VP.n44 VP.n29 161.3
R2865 VP.n46 VP.n45 161.3
R2866 VP.n47 VP.n28 161.3
R2867 VP.n49 VP.n48 161.3
R2868 VP.n50 VP.n27 161.3
R2869 VP.n52 VP.n51 161.3
R2870 VP.n53 VP.n26 161.3
R2871 VP.n55 VP.n54 161.3
R2872 VP.n56 VP.n25 161.3
R2873 VP.n58 VP.n57 161.3
R2874 VP.n59 VP.n24 161.3
R2875 VP.n62 VP.n61 161.3
R2876 VP.n63 VP.n23 161.3
R2877 VP.n65 VP.n64 161.3
R2878 VP.n66 VP.n22 161.3
R2879 VP.n68 VP.n67 161.3
R2880 VP.n69 VP.n21 161.3
R2881 VP.n71 VP.n70 161.3
R2882 VP.n72 VP.n20 161.3
R2883 VP.n74 VP.n73 161.3
R2884 VP.n131 VP.n130 161.3
R2885 VP.n129 VP.n1 161.3
R2886 VP.n128 VP.n127 161.3
R2887 VP.n126 VP.n2 161.3
R2888 VP.n125 VP.n124 161.3
R2889 VP.n123 VP.n3 161.3
R2890 VP.n122 VP.n121 161.3
R2891 VP.n120 VP.n4 161.3
R2892 VP.n119 VP.n118 161.3
R2893 VP.n116 VP.n5 161.3
R2894 VP.n115 VP.n114 161.3
R2895 VP.n113 VP.n6 161.3
R2896 VP.n112 VP.n111 161.3
R2897 VP.n110 VP.n7 161.3
R2898 VP.n109 VP.n108 161.3
R2899 VP.n107 VP.n8 161.3
R2900 VP.n106 VP.n105 161.3
R2901 VP.n104 VP.n9 161.3
R2902 VP.n103 VP.n102 161.3
R2903 VP.n101 VP.n10 161.3
R2904 VP.n100 VP.n99 161.3
R2905 VP.n98 VP.n11 161.3
R2906 VP.n97 VP.n96 161.3
R2907 VP.n95 VP.n12 161.3
R2908 VP.n94 VP.n93 161.3
R2909 VP.n92 VP.n13 161.3
R2910 VP.n90 VP.n89 161.3
R2911 VP.n88 VP.n14 161.3
R2912 VP.n87 VP.n86 161.3
R2913 VP.n85 VP.n15 161.3
R2914 VP.n84 VP.n83 161.3
R2915 VP.n82 VP.n16 161.3
R2916 VP.n81 VP.n80 161.3
R2917 VP.n79 VP.n17 161.3
R2918 VP.n78 VP.n77 161.3
R2919 VP.n33 VP.t1 149.214
R2920 VP.n104 VP.t3 116.647
R2921 VP.n18 VP.t2 116.647
R2922 VP.n91 VP.t4 116.647
R2923 VP.n117 VP.t5 116.647
R2924 VP.n0 VP.t6 116.647
R2925 VP.n47 VP.t0 116.647
R2926 VP.n19 VP.t8 116.647
R2927 VP.n60 VP.t7 116.647
R2928 VP.n34 VP.t9 116.647
R2929 VP.n76 VP.n18 88.1101
R2930 VP.n132 VP.n0 88.1101
R2931 VP.n75 VP.n19 88.1101
R2932 VP.n76 VP.n75 65.8289
R2933 VP.n34 VP.n33 61.9406
R2934 VP.n98 VP.n97 53.6055
R2935 VP.n111 VP.n110 53.6055
R2936 VP.n54 VP.n53 53.6055
R2937 VP.n41 VP.n40 53.6055
R2938 VP.n85 VP.n84 49.7204
R2939 VP.n124 VP.n123 49.7204
R2940 VP.n67 VP.n66 49.7204
R2941 VP.n84 VP.n16 31.2664
R2942 VP.n124 VP.n2 31.2664
R2943 VP.n67 VP.n21 31.2664
R2944 VP.n99 VP.n98 27.3813
R2945 VP.n110 VP.n109 27.3813
R2946 VP.n53 VP.n52 27.3813
R2947 VP.n42 VP.n41 27.3813
R2948 VP.n79 VP.n78 24.4675
R2949 VP.n80 VP.n79 24.4675
R2950 VP.n80 VP.n16 24.4675
R2951 VP.n86 VP.n85 24.4675
R2952 VP.n86 VP.n14 24.4675
R2953 VP.n90 VP.n14 24.4675
R2954 VP.n93 VP.n92 24.4675
R2955 VP.n93 VP.n12 24.4675
R2956 VP.n97 VP.n12 24.4675
R2957 VP.n99 VP.n10 24.4675
R2958 VP.n103 VP.n10 24.4675
R2959 VP.n104 VP.n103 24.4675
R2960 VP.n105 VP.n104 24.4675
R2961 VP.n105 VP.n8 24.4675
R2962 VP.n109 VP.n8 24.4675
R2963 VP.n111 VP.n6 24.4675
R2964 VP.n115 VP.n6 24.4675
R2965 VP.n116 VP.n115 24.4675
R2966 VP.n118 VP.n4 24.4675
R2967 VP.n122 VP.n4 24.4675
R2968 VP.n123 VP.n122 24.4675
R2969 VP.n128 VP.n2 24.4675
R2970 VP.n129 VP.n128 24.4675
R2971 VP.n130 VP.n129 24.4675
R2972 VP.n71 VP.n21 24.4675
R2973 VP.n72 VP.n71 24.4675
R2974 VP.n73 VP.n72 24.4675
R2975 VP.n54 VP.n25 24.4675
R2976 VP.n58 VP.n25 24.4675
R2977 VP.n59 VP.n58 24.4675
R2978 VP.n61 VP.n23 24.4675
R2979 VP.n65 VP.n23 24.4675
R2980 VP.n66 VP.n65 24.4675
R2981 VP.n42 VP.n29 24.4675
R2982 VP.n46 VP.n29 24.4675
R2983 VP.n47 VP.n46 24.4675
R2984 VP.n48 VP.n47 24.4675
R2985 VP.n48 VP.n27 24.4675
R2986 VP.n52 VP.n27 24.4675
R2987 VP.n36 VP.n35 24.4675
R2988 VP.n36 VP.n31 24.4675
R2989 VP.n40 VP.n31 24.4675
R2990 VP.n92 VP.n91 13.2127
R2991 VP.n117 VP.n116 13.2127
R2992 VP.n60 VP.n59 13.2127
R2993 VP.n35 VP.n34 13.2127
R2994 VP.n91 VP.n90 11.2553
R2995 VP.n118 VP.n117 11.2553
R2996 VP.n61 VP.n60 11.2553
R2997 VP.n33 VP.n32 2.48785
R2998 VP.n78 VP.n18 1.95786
R2999 VP.n130 VP.n0 1.95786
R3000 VP.n73 VP.n19 1.95786
R3001 VP.n75 VP.n74 0.354971
R3002 VP.n77 VP.n76 0.354971
R3003 VP.n132 VP.n131 0.354971
R3004 VP VP.n132 0.26696
R3005 VP.n37 VP.n32 0.189894
R3006 VP.n38 VP.n37 0.189894
R3007 VP.n39 VP.n38 0.189894
R3008 VP.n39 VP.n30 0.189894
R3009 VP.n43 VP.n30 0.189894
R3010 VP.n44 VP.n43 0.189894
R3011 VP.n45 VP.n44 0.189894
R3012 VP.n45 VP.n28 0.189894
R3013 VP.n49 VP.n28 0.189894
R3014 VP.n50 VP.n49 0.189894
R3015 VP.n51 VP.n50 0.189894
R3016 VP.n51 VP.n26 0.189894
R3017 VP.n55 VP.n26 0.189894
R3018 VP.n56 VP.n55 0.189894
R3019 VP.n57 VP.n56 0.189894
R3020 VP.n57 VP.n24 0.189894
R3021 VP.n62 VP.n24 0.189894
R3022 VP.n63 VP.n62 0.189894
R3023 VP.n64 VP.n63 0.189894
R3024 VP.n64 VP.n22 0.189894
R3025 VP.n68 VP.n22 0.189894
R3026 VP.n69 VP.n68 0.189894
R3027 VP.n70 VP.n69 0.189894
R3028 VP.n70 VP.n20 0.189894
R3029 VP.n74 VP.n20 0.189894
R3030 VP.n77 VP.n17 0.189894
R3031 VP.n81 VP.n17 0.189894
R3032 VP.n82 VP.n81 0.189894
R3033 VP.n83 VP.n82 0.189894
R3034 VP.n83 VP.n15 0.189894
R3035 VP.n87 VP.n15 0.189894
R3036 VP.n88 VP.n87 0.189894
R3037 VP.n89 VP.n88 0.189894
R3038 VP.n89 VP.n13 0.189894
R3039 VP.n94 VP.n13 0.189894
R3040 VP.n95 VP.n94 0.189894
R3041 VP.n96 VP.n95 0.189894
R3042 VP.n96 VP.n11 0.189894
R3043 VP.n100 VP.n11 0.189894
R3044 VP.n101 VP.n100 0.189894
R3045 VP.n102 VP.n101 0.189894
R3046 VP.n102 VP.n9 0.189894
R3047 VP.n106 VP.n9 0.189894
R3048 VP.n107 VP.n106 0.189894
R3049 VP.n108 VP.n107 0.189894
R3050 VP.n108 VP.n7 0.189894
R3051 VP.n112 VP.n7 0.189894
R3052 VP.n113 VP.n112 0.189894
R3053 VP.n114 VP.n113 0.189894
R3054 VP.n114 VP.n5 0.189894
R3055 VP.n119 VP.n5 0.189894
R3056 VP.n120 VP.n119 0.189894
R3057 VP.n121 VP.n120 0.189894
R3058 VP.n121 VP.n3 0.189894
R3059 VP.n125 VP.n3 0.189894
R3060 VP.n126 VP.n125 0.189894
R3061 VP.n127 VP.n126 0.189894
R3062 VP.n127 VP.n1 0.189894
R3063 VP.n131 VP.n1 0.189894
R3064 VDD1.n1 VDD1.t8 67.0522
R3065 VDD1.n3 VDD1.t7 67.052
R3066 VDD1.n5 VDD1.n4 65.0371
R3067 VDD1.n1 VDD1.n0 62.3329
R3068 VDD1.n7 VDD1.n6 62.3327
R3069 VDD1.n3 VDD1.n2 62.3317
R3070 VDD1.n7 VDD1.n5 60.0634
R3071 VDD1 VDD1.n7 2.70309
R3072 VDD1.n6 VDD1.t2 1.03878
R3073 VDD1.n6 VDD1.t1 1.03878
R3074 VDD1.n0 VDD1.t0 1.03878
R3075 VDD1.n0 VDD1.t9 1.03878
R3076 VDD1.n4 VDD1.t4 1.03878
R3077 VDD1.n4 VDD1.t3 1.03878
R3078 VDD1.n2 VDD1.t5 1.03878
R3079 VDD1.n2 VDD1.t6 1.03878
R3080 VDD1 VDD1.n1 0.978948
R3081 VDD1.n5 VDD1.n3 0.865413
C0 VP VN 11.6827f
C1 VDD2 VP 0.753897f
C2 VTAIL VDD1 13.8139f
C3 VDD2 VN 17.839699f
C4 VTAIL VP 18.729599f
C5 VDD1 VP 18.433401f
C6 VTAIL VN 18.7142f
C7 VDD1 VN 0.156412f
C8 VTAIL VDD2 13.8738f
C9 VDD1 VDD2 3.04796f
C10 VDD2 B 9.982583f
C11 VDD1 B 9.991744f
C12 VTAIL B 12.091363f
C13 VN B 25.07115f
C14 VP B 23.608973f
C15 VDD1.t8 B 4.257259f
C16 VDD1.t0 B 0.361301f
C17 VDD1.t9 B 0.361301f
C18 VDD1.n0 B 3.30601f
C19 VDD1.n1 B 1.07377f
C20 VDD1.t7 B 4.25724f
C21 VDD1.t5 B 0.361301f
C22 VDD1.t6 B 0.361301f
C23 VDD1.n2 B 3.30601f
C24 VDD1.n3 B 1.06567f
C25 VDD1.t4 B 0.361301f
C26 VDD1.t3 B 0.361301f
C27 VDD1.n4 B 3.33496f
C28 VDD1.n5 B 4.03845f
C29 VDD1.t2 B 0.361301f
C30 VDD1.t1 B 0.361301f
C31 VDD1.n6 B 3.306f
C32 VDD1.n7 B 4.07984f
C33 VP.t6 B 3.19377f
C34 VP.n0 B 1.15693f
C35 VP.n1 B 0.015437f
C36 VP.n2 B 0.030995f
C37 VP.n3 B 0.015437f
C38 VP.n4 B 0.028771f
C39 VP.n5 B 0.015437f
C40 VP.t5 B 3.19377f
C41 VP.n6 B 0.028771f
C42 VP.n7 B 0.015437f
C43 VP.n8 B 0.028771f
C44 VP.n9 B 0.015437f
C45 VP.t3 B 3.19377f
C46 VP.n10 B 0.028771f
C47 VP.n11 B 0.015437f
C48 VP.n12 B 0.028771f
C49 VP.n13 B 0.015437f
C50 VP.t4 B 3.19377f
C51 VP.n14 B 0.028771f
C52 VP.n15 B 0.015437f
C53 VP.n16 B 0.030995f
C54 VP.n17 B 0.015437f
C55 VP.t2 B 3.19377f
C56 VP.n18 B 1.15693f
C57 VP.t8 B 3.19377f
C58 VP.n19 B 1.15693f
C59 VP.n20 B 0.015437f
C60 VP.n21 B 0.030995f
C61 VP.n22 B 0.015437f
C62 VP.n23 B 0.028771f
C63 VP.n24 B 0.015437f
C64 VP.t7 B 3.19377f
C65 VP.n25 B 0.028771f
C66 VP.n26 B 0.015437f
C67 VP.n27 B 0.028771f
C68 VP.n28 B 0.015437f
C69 VP.t0 B 3.19377f
C70 VP.n29 B 0.028771f
C71 VP.n30 B 0.015437f
C72 VP.n31 B 0.028771f
C73 VP.n32 B 0.201507f
C74 VP.t9 B 3.19377f
C75 VP.t1 B 3.4607f
C76 VP.n33 B 1.10389f
C77 VP.n34 B 1.15447f
C78 VP.n35 B 0.022237f
C79 VP.n36 B 0.028771f
C80 VP.n37 B 0.015437f
C81 VP.n38 B 0.015437f
C82 VP.n39 B 0.015437f
C83 VP.n40 B 0.027227f
C84 VP.n41 B 0.016517f
C85 VP.n42 B 0.030102f
C86 VP.n43 B 0.015437f
C87 VP.n44 B 0.015437f
C88 VP.n45 B 0.015437f
C89 VP.n46 B 0.028771f
C90 VP.n47 B 1.1123f
C91 VP.n48 B 0.028771f
C92 VP.n49 B 0.015437f
C93 VP.n50 B 0.015437f
C94 VP.n51 B 0.015437f
C95 VP.n52 B 0.030102f
C96 VP.n53 B 0.016517f
C97 VP.n54 B 0.027227f
C98 VP.n55 B 0.015437f
C99 VP.n56 B 0.015437f
C100 VP.n57 B 0.015437f
C101 VP.n58 B 0.028771f
C102 VP.n59 B 0.022237f
C103 VP.n60 B 1.09773f
C104 VP.n61 B 0.021101f
C105 VP.n62 B 0.015437f
C106 VP.n63 B 0.015437f
C107 VP.n64 B 0.015437f
C108 VP.n65 B 0.028771f
C109 VP.n66 B 0.028483f
C110 VP.n67 B 0.014368f
C111 VP.n68 B 0.015437f
C112 VP.n69 B 0.015437f
C113 VP.n70 B 0.015437f
C114 VP.n71 B 0.028771f
C115 VP.n72 B 0.028771f
C116 VP.n73 B 0.015703f
C117 VP.n74 B 0.024916f
C118 VP.n75 B 1.28968f
C119 VP.n76 B 1.29811f
C120 VP.n77 B 0.024916f
C121 VP.n78 B 0.015703f
C122 VP.n79 B 0.028771f
C123 VP.n80 B 0.028771f
C124 VP.n81 B 0.015437f
C125 VP.n82 B 0.015437f
C126 VP.n83 B 0.015437f
C127 VP.n84 B 0.014368f
C128 VP.n85 B 0.028483f
C129 VP.n86 B 0.028771f
C130 VP.n87 B 0.015437f
C131 VP.n88 B 0.015437f
C132 VP.n89 B 0.015437f
C133 VP.n90 B 0.021101f
C134 VP.n91 B 1.09773f
C135 VP.n92 B 0.022237f
C136 VP.n93 B 0.028771f
C137 VP.n94 B 0.015437f
C138 VP.n95 B 0.015437f
C139 VP.n96 B 0.015437f
C140 VP.n97 B 0.027227f
C141 VP.n98 B 0.016517f
C142 VP.n99 B 0.030102f
C143 VP.n100 B 0.015437f
C144 VP.n101 B 0.015437f
C145 VP.n102 B 0.015437f
C146 VP.n103 B 0.028771f
C147 VP.n104 B 1.1123f
C148 VP.n105 B 0.028771f
C149 VP.n106 B 0.015437f
C150 VP.n107 B 0.015437f
C151 VP.n108 B 0.015437f
C152 VP.n109 B 0.030102f
C153 VP.n110 B 0.016517f
C154 VP.n111 B 0.027227f
C155 VP.n112 B 0.015437f
C156 VP.n113 B 0.015437f
C157 VP.n114 B 0.015437f
C158 VP.n115 B 0.028771f
C159 VP.n116 B 0.022237f
C160 VP.n117 B 1.09773f
C161 VP.n118 B 0.021101f
C162 VP.n119 B 0.015437f
C163 VP.n120 B 0.015437f
C164 VP.n121 B 0.015437f
C165 VP.n122 B 0.028771f
C166 VP.n123 B 0.028483f
C167 VP.n124 B 0.014368f
C168 VP.n125 B 0.015437f
C169 VP.n126 B 0.015437f
C170 VP.n127 B 0.015437f
C171 VP.n128 B 0.028771f
C172 VP.n129 B 0.028771f
C173 VP.n130 B 0.015703f
C174 VP.n131 B 0.024916f
C175 VP.n132 B 0.049066f
C176 VDD2.t6 B 4.20735f
C177 VDD2.t0 B 0.357067f
C178 VDD2.t7 B 0.357067f
C179 VDD2.n0 B 3.26727f
C180 VDD2.n1 B 1.05319f
C181 VDD2.t5 B 0.357067f
C182 VDD2.t2 B 0.357067f
C183 VDD2.n2 B 3.29588f
C184 VDD2.n3 B 3.83272f
C185 VDD2.t1 B 4.17746f
C186 VDD2.n4 B 3.96021f
C187 VDD2.t8 B 0.357067f
C188 VDD2.t9 B 0.357067f
C189 VDD2.n5 B 3.26727f
C190 VDD2.n6 B 0.546313f
C191 VDD2.t3 B 0.357067f
C192 VDD2.t4 B 0.357067f
C193 VDD2.n7 B 3.29582f
C194 VTAIL.t11 B 0.363702f
C195 VTAIL.t14 B 0.363702f
C196 VTAIL.n0 B 3.25873f
C197 VTAIL.n1 B 0.629443f
C198 VTAIL.t16 B 4.1642f
C199 VTAIL.n2 B 0.782933f
C200 VTAIL.t17 B 0.363702f
C201 VTAIL.t1 B 0.363702f
C202 VTAIL.n3 B 3.25873f
C203 VTAIL.n4 B 0.803078f
C204 VTAIL.t2 B 0.363702f
C205 VTAIL.t19 B 0.363702f
C206 VTAIL.n5 B 3.25873f
C207 VTAIL.n6 B 2.69565f
C208 VTAIL.t8 B 0.363702f
C209 VTAIL.t9 B 0.363702f
C210 VTAIL.n7 B 3.25874f
C211 VTAIL.n8 B 2.69564f
C212 VTAIL.t6 B 0.363702f
C213 VTAIL.t13 B 0.363702f
C214 VTAIL.n9 B 3.25874f
C215 VTAIL.n10 B 0.803068f
C216 VTAIL.t15 B 4.16423f
C217 VTAIL.n11 B 0.782902f
C218 VTAIL.t3 B 0.363702f
C219 VTAIL.t5 B 0.363702f
C220 VTAIL.n12 B 3.25874f
C221 VTAIL.n13 B 0.696473f
C222 VTAIL.t4 B 0.363702f
C223 VTAIL.t18 B 0.363702f
C224 VTAIL.n14 B 3.25874f
C225 VTAIL.n15 B 0.803068f
C226 VTAIL.t0 B 4.1642f
C227 VTAIL.n16 B 2.49583f
C228 VTAIL.t7 B 4.1642f
C229 VTAIL.n17 B 2.49583f
C230 VTAIL.t10 B 0.363702f
C231 VTAIL.t12 B 0.363702f
C232 VTAIL.n18 B 3.25873f
C233 VTAIL.n19 B 0.583855f
C234 VN.t7 B 3.1531f
C235 VN.n0 B 1.1422f
C236 VN.n1 B 0.015241f
C237 VN.n2 B 0.030601f
C238 VN.n3 B 0.015241f
C239 VN.n4 B 0.028405f
C240 VN.n5 B 0.015241f
C241 VN.t4 B 3.1531f
C242 VN.n6 B 0.028405f
C243 VN.n7 B 0.015241f
C244 VN.n8 B 0.028405f
C245 VN.n9 B 0.015241f
C246 VN.t2 B 3.1531f
C247 VN.n10 B 0.028405f
C248 VN.n11 B 0.015241f
C249 VN.n12 B 0.028405f
C250 VN.n13 B 0.198941f
C251 VN.t9 B 3.1531f
C252 VN.t3 B 3.41663f
C253 VN.n14 B 1.08983f
C254 VN.n15 B 1.13977f
C255 VN.n16 B 0.021954f
C256 VN.n17 B 0.028405f
C257 VN.n18 B 0.015241f
C258 VN.n19 B 0.015241f
C259 VN.n20 B 0.015241f
C260 VN.n21 B 0.026881f
C261 VN.n22 B 0.016307f
C262 VN.n23 B 0.029718f
C263 VN.n24 B 0.015241f
C264 VN.n25 B 0.015241f
C265 VN.n26 B 0.015241f
C266 VN.n27 B 0.028405f
C267 VN.n28 B 1.09814f
C268 VN.n29 B 0.028405f
C269 VN.n30 B 0.015241f
C270 VN.n31 B 0.015241f
C271 VN.n32 B 0.015241f
C272 VN.n33 B 0.029718f
C273 VN.n34 B 0.016307f
C274 VN.n35 B 0.026881f
C275 VN.n36 B 0.015241f
C276 VN.n37 B 0.015241f
C277 VN.n38 B 0.015241f
C278 VN.n39 B 0.028405f
C279 VN.n40 B 0.021954f
C280 VN.n41 B 1.08376f
C281 VN.n42 B 0.020832f
C282 VN.n43 B 0.015241f
C283 VN.n44 B 0.015241f
C284 VN.n45 B 0.015241f
C285 VN.n46 B 0.028405f
C286 VN.n47 B 0.02812f
C287 VN.n48 B 0.014185f
C288 VN.n49 B 0.015241f
C289 VN.n50 B 0.015241f
C290 VN.n51 B 0.015241f
C291 VN.n52 B 0.028405f
C292 VN.n53 B 0.028405f
C293 VN.n54 B 0.015503f
C294 VN.n55 B 0.024598f
C295 VN.n56 B 0.048441f
C296 VN.t8 B 3.1531f
C297 VN.n57 B 1.1422f
C298 VN.n58 B 0.015241f
C299 VN.n59 B 0.030601f
C300 VN.n60 B 0.015241f
C301 VN.n61 B 0.028405f
C302 VN.n62 B 0.015241f
C303 VN.t1 B 3.1531f
C304 VN.n63 B 0.028405f
C305 VN.n64 B 0.015241f
C306 VN.n65 B 0.028405f
C307 VN.n66 B 0.015241f
C308 VN.t0 B 3.1531f
C309 VN.n67 B 0.028405f
C310 VN.n68 B 0.015241f
C311 VN.n69 B 0.028405f
C312 VN.n70 B 0.198941f
C313 VN.t6 B 3.1531f
C314 VN.t5 B 3.41663f
C315 VN.n71 B 1.08983f
C316 VN.n72 B 1.13977f
C317 VN.n73 B 0.021954f
C318 VN.n74 B 0.028405f
C319 VN.n75 B 0.015241f
C320 VN.n76 B 0.015241f
C321 VN.n77 B 0.015241f
C322 VN.n78 B 0.026881f
C323 VN.n79 B 0.016307f
C324 VN.n80 B 0.029718f
C325 VN.n81 B 0.015241f
C326 VN.n82 B 0.015241f
C327 VN.n83 B 0.015241f
C328 VN.n84 B 0.028405f
C329 VN.n85 B 1.09814f
C330 VN.n86 B 0.028405f
C331 VN.n87 B 0.015241f
C332 VN.n88 B 0.015241f
C333 VN.n89 B 0.015241f
C334 VN.n90 B 0.029718f
C335 VN.n91 B 0.016307f
C336 VN.n92 B 0.026881f
C337 VN.n93 B 0.015241f
C338 VN.n94 B 0.015241f
C339 VN.n95 B 0.015241f
C340 VN.n96 B 0.028405f
C341 VN.n97 B 0.021954f
C342 VN.n98 B 1.08376f
C343 VN.n99 B 0.020832f
C344 VN.n100 B 0.015241f
C345 VN.n101 B 0.015241f
C346 VN.n102 B 0.015241f
C347 VN.n103 B 0.028405f
C348 VN.n104 B 0.02812f
C349 VN.n105 B 0.014185f
C350 VN.n106 B 0.015241f
C351 VN.n107 B 0.015241f
C352 VN.n108 B 0.015241f
C353 VN.n109 B 0.028405f
C354 VN.n110 B 0.028405f
C355 VN.n111 B 0.015503f
C356 VN.n112 B 0.024598f
C357 VN.n113 B 1.27898f
.ends

