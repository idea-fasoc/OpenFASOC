* NGSPICE file created from diff_pair_sample_0326.ext - technology: sky130A

.subckt diff_pair_sample_0326 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VN.t0 VDD2.t7 B.t0 sky130_fd_pr__nfet_01v8 ad=0.83985 pd=5.42 as=0.83985 ps=5.42 w=5.09 l=3.71
X1 VTAIL.t2 VP.t0 VDD1.t7 B.t2 sky130_fd_pr__nfet_01v8 ad=0.83985 pd=5.42 as=0.83985 ps=5.42 w=5.09 l=3.71
X2 VDD2.t0 VN.t1 VTAIL.t14 B.t1 sky130_fd_pr__nfet_01v8 ad=0.83985 pd=5.42 as=0.83985 ps=5.42 w=5.09 l=3.71
X3 B.t21 B.t19 B.t20 B.t16 sky130_fd_pr__nfet_01v8 ad=1.9851 pd=10.96 as=0 ps=0 w=5.09 l=3.71
X4 VTAIL.t4 VP.t1 VDD1.t6 B.t4 sky130_fd_pr__nfet_01v8 ad=1.9851 pd=10.96 as=0.83985 ps=5.42 w=5.09 l=3.71
X5 VDD1.t5 VP.t2 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=0.83985 pd=5.42 as=1.9851 ps=10.96 w=5.09 l=3.71
X6 VTAIL.t0 VP.t3 VDD1.t4 B.t0 sky130_fd_pr__nfet_01v8 ad=0.83985 pd=5.42 as=0.83985 ps=5.42 w=5.09 l=3.71
X7 VTAIL.t13 VN.t2 VDD2.t3 B.t4 sky130_fd_pr__nfet_01v8 ad=1.9851 pd=10.96 as=0.83985 ps=5.42 w=5.09 l=3.71
X8 VTAIL.t12 VN.t3 VDD2.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.83985 pd=5.42 as=0.83985 ps=5.42 w=5.09 l=3.71
X9 VDD1.t3 VP.t4 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=0.83985 pd=5.42 as=1.9851 ps=10.96 w=5.09 l=3.71
X10 VDD2.t4 VN.t4 VTAIL.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=0.83985 pd=5.42 as=1.9851 ps=10.96 w=5.09 l=3.71
X11 VDD1.t2 VP.t5 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.83985 pd=5.42 as=0.83985 ps=5.42 w=5.09 l=3.71
X12 VTAIL.t10 VN.t5 VDD2.t5 B.t3 sky130_fd_pr__nfet_01v8 ad=1.9851 pd=10.96 as=0.83985 ps=5.42 w=5.09 l=3.71
X13 B.t18 B.t15 B.t17 B.t16 sky130_fd_pr__nfet_01v8 ad=1.9851 pd=10.96 as=0 ps=0 w=5.09 l=3.71
X14 VDD2.t1 VN.t6 VTAIL.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=0.83985 pd=5.42 as=0.83985 ps=5.42 w=5.09 l=3.71
X15 VTAIL.t3 VP.t6 VDD1.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=1.9851 pd=10.96 as=0.83985 ps=5.42 w=5.09 l=3.71
X16 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=1.9851 pd=10.96 as=0 ps=0 w=5.09 l=3.71
X17 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=1.9851 pd=10.96 as=0 ps=0 w=5.09 l=3.71
X18 VDD2.t6 VN.t7 VTAIL.t8 B.t6 sky130_fd_pr__nfet_01v8 ad=0.83985 pd=5.42 as=1.9851 ps=10.96 w=5.09 l=3.71
X19 VDD1.t0 VP.t7 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=0.83985 pd=5.42 as=0.83985 ps=5.42 w=5.09 l=3.71
R0 VN.n76 VN.n75 161.3
R1 VN.n74 VN.n40 161.3
R2 VN.n73 VN.n72 161.3
R3 VN.n71 VN.n41 161.3
R4 VN.n70 VN.n69 161.3
R5 VN.n68 VN.n42 161.3
R6 VN.n67 VN.n66 161.3
R7 VN.n65 VN.n43 161.3
R8 VN.n64 VN.n63 161.3
R9 VN.n62 VN.n44 161.3
R10 VN.n61 VN.n60 161.3
R11 VN.n59 VN.n46 161.3
R12 VN.n58 VN.n57 161.3
R13 VN.n56 VN.n47 161.3
R14 VN.n55 VN.n54 161.3
R15 VN.n53 VN.n48 161.3
R16 VN.n52 VN.n51 161.3
R17 VN.n37 VN.n36 161.3
R18 VN.n35 VN.n1 161.3
R19 VN.n34 VN.n33 161.3
R20 VN.n32 VN.n2 161.3
R21 VN.n31 VN.n30 161.3
R22 VN.n29 VN.n3 161.3
R23 VN.n28 VN.n27 161.3
R24 VN.n26 VN.n4 161.3
R25 VN.n25 VN.n24 161.3
R26 VN.n22 VN.n5 161.3
R27 VN.n21 VN.n20 161.3
R28 VN.n19 VN.n6 161.3
R29 VN.n18 VN.n17 161.3
R30 VN.n16 VN.n7 161.3
R31 VN.n15 VN.n14 161.3
R32 VN.n13 VN.n8 161.3
R33 VN.n12 VN.n11 161.3
R34 VN.n38 VN.n0 87.1314
R35 VN.n77 VN.n39 87.1314
R36 VN.n10 VN.n9 73.9973
R37 VN.n50 VN.n49 73.9973
R38 VN.n49 VN.t4 64.934
R39 VN.n9 VN.t5 64.934
R40 VN VN.n77 51.0511
R41 VN.n30 VN.n2 44.3785
R42 VN.n69 VN.n41 44.3785
R43 VN.n17 VN.n16 40.4934
R44 VN.n17 VN.n6 40.4934
R45 VN.n57 VN.n56 40.4934
R46 VN.n57 VN.n46 40.4934
R47 VN.n30 VN.n29 36.6083
R48 VN.n69 VN.n68 36.6083
R49 VN.n10 VN.t1 33.0649
R50 VN.n23 VN.t0 33.0649
R51 VN.n0 VN.t7 33.0649
R52 VN.n50 VN.t3 33.0649
R53 VN.n45 VN.t6 33.0649
R54 VN.n39 VN.t2 33.0649
R55 VN.n11 VN.n8 24.4675
R56 VN.n15 VN.n8 24.4675
R57 VN.n16 VN.n15 24.4675
R58 VN.n21 VN.n6 24.4675
R59 VN.n22 VN.n21 24.4675
R60 VN.n24 VN.n22 24.4675
R61 VN.n28 VN.n4 24.4675
R62 VN.n29 VN.n28 24.4675
R63 VN.n34 VN.n2 24.4675
R64 VN.n35 VN.n34 24.4675
R65 VN.n36 VN.n35 24.4675
R66 VN.n56 VN.n55 24.4675
R67 VN.n55 VN.n48 24.4675
R68 VN.n51 VN.n48 24.4675
R69 VN.n68 VN.n67 24.4675
R70 VN.n67 VN.n43 24.4675
R71 VN.n63 VN.n62 24.4675
R72 VN.n62 VN.n61 24.4675
R73 VN.n61 VN.n46 24.4675
R74 VN.n75 VN.n74 24.4675
R75 VN.n74 VN.n73 24.4675
R76 VN.n73 VN.n41 24.4675
R77 VN.n23 VN.n4 23.4888
R78 VN.n45 VN.n43 23.4888
R79 VN.n52 VN.n49 3.37703
R80 VN.n12 VN.n9 3.37703
R81 VN.n36 VN.n0 2.93654
R82 VN.n75 VN.n39 2.93654
R83 VN.n11 VN.n10 0.97918
R84 VN.n24 VN.n23 0.97918
R85 VN.n51 VN.n50 0.97918
R86 VN.n63 VN.n45 0.97918
R87 VN.n77 VN.n76 0.354971
R88 VN.n38 VN.n37 0.354971
R89 VN VN.n38 0.26696
R90 VN.n76 VN.n40 0.189894
R91 VN.n72 VN.n40 0.189894
R92 VN.n72 VN.n71 0.189894
R93 VN.n71 VN.n70 0.189894
R94 VN.n70 VN.n42 0.189894
R95 VN.n66 VN.n42 0.189894
R96 VN.n66 VN.n65 0.189894
R97 VN.n65 VN.n64 0.189894
R98 VN.n64 VN.n44 0.189894
R99 VN.n60 VN.n44 0.189894
R100 VN.n60 VN.n59 0.189894
R101 VN.n59 VN.n58 0.189894
R102 VN.n58 VN.n47 0.189894
R103 VN.n54 VN.n47 0.189894
R104 VN.n54 VN.n53 0.189894
R105 VN.n53 VN.n52 0.189894
R106 VN.n13 VN.n12 0.189894
R107 VN.n14 VN.n13 0.189894
R108 VN.n14 VN.n7 0.189894
R109 VN.n18 VN.n7 0.189894
R110 VN.n19 VN.n18 0.189894
R111 VN.n20 VN.n19 0.189894
R112 VN.n20 VN.n5 0.189894
R113 VN.n25 VN.n5 0.189894
R114 VN.n26 VN.n25 0.189894
R115 VN.n27 VN.n26 0.189894
R116 VN.n27 VN.n3 0.189894
R117 VN.n31 VN.n3 0.189894
R118 VN.n32 VN.n31 0.189894
R119 VN.n33 VN.n32 0.189894
R120 VN.n33 VN.n1 0.189894
R121 VN.n37 VN.n1 0.189894
R122 VDD2.n2 VDD2.n1 74.5499
R123 VDD2.n2 VDD2.n0 74.5499
R124 VDD2 VDD2.n5 74.5471
R125 VDD2.n4 VDD2.n3 72.864
R126 VDD2.n4 VDD2.n2 43.7756
R127 VDD2.n5 VDD2.t2 3.89048
R128 VDD2.n5 VDD2.t4 3.89048
R129 VDD2.n3 VDD2.t3 3.89048
R130 VDD2.n3 VDD2.t1 3.89048
R131 VDD2.n1 VDD2.t7 3.89048
R132 VDD2.n1 VDD2.t6 3.89048
R133 VDD2.n0 VDD2.t5 3.89048
R134 VDD2.n0 VDD2.t0 3.89048
R135 VDD2 VDD2.n4 1.80007
R136 VTAIL.n11 VTAIL.t3 60.0752
R137 VTAIL.n10 VTAIL.t11 60.0752
R138 VTAIL.n7 VTAIL.t13 60.0752
R139 VTAIL.n15 VTAIL.t8 60.0751
R140 VTAIL.n2 VTAIL.t10 60.0751
R141 VTAIL.n3 VTAIL.t7 60.0751
R142 VTAIL.n6 VTAIL.t4 60.0751
R143 VTAIL.n14 VTAIL.t6 60.0751
R144 VTAIL.n13 VTAIL.n12 56.1853
R145 VTAIL.n9 VTAIL.n8 56.1853
R146 VTAIL.n1 VTAIL.n0 56.185
R147 VTAIL.n5 VTAIL.n4 56.185
R148 VTAIL.n15 VTAIL.n14 20.2376
R149 VTAIL.n7 VTAIL.n6 20.2376
R150 VTAIL.n0 VTAIL.t14 3.89048
R151 VTAIL.n0 VTAIL.t15 3.89048
R152 VTAIL.n4 VTAIL.t5 3.89048
R153 VTAIL.n4 VTAIL.t2 3.89048
R154 VTAIL.n12 VTAIL.t1 3.89048
R155 VTAIL.n12 VTAIL.t0 3.89048
R156 VTAIL.n8 VTAIL.t9 3.89048
R157 VTAIL.n8 VTAIL.t12 3.89048
R158 VTAIL.n9 VTAIL.n7 3.48326
R159 VTAIL.n10 VTAIL.n9 3.48326
R160 VTAIL.n13 VTAIL.n11 3.48326
R161 VTAIL.n14 VTAIL.n13 3.48326
R162 VTAIL.n6 VTAIL.n5 3.48326
R163 VTAIL.n5 VTAIL.n3 3.48326
R164 VTAIL.n2 VTAIL.n1 3.48326
R165 VTAIL VTAIL.n15 3.42507
R166 VTAIL.n11 VTAIL.n10 0.470328
R167 VTAIL.n3 VTAIL.n2 0.470328
R168 VTAIL VTAIL.n1 0.0586897
R169 B.n809 B.n808 585
R170 B.n253 B.n149 585
R171 B.n252 B.n251 585
R172 B.n250 B.n249 585
R173 B.n248 B.n247 585
R174 B.n246 B.n245 585
R175 B.n244 B.n243 585
R176 B.n242 B.n241 585
R177 B.n240 B.n239 585
R178 B.n238 B.n237 585
R179 B.n236 B.n235 585
R180 B.n234 B.n233 585
R181 B.n232 B.n231 585
R182 B.n230 B.n229 585
R183 B.n228 B.n227 585
R184 B.n226 B.n225 585
R185 B.n224 B.n223 585
R186 B.n222 B.n221 585
R187 B.n220 B.n219 585
R188 B.n218 B.n217 585
R189 B.n216 B.n215 585
R190 B.n213 B.n212 585
R191 B.n211 B.n210 585
R192 B.n209 B.n208 585
R193 B.n207 B.n206 585
R194 B.n205 B.n204 585
R195 B.n203 B.n202 585
R196 B.n201 B.n200 585
R197 B.n199 B.n198 585
R198 B.n197 B.n196 585
R199 B.n195 B.n194 585
R200 B.n192 B.n191 585
R201 B.n190 B.n189 585
R202 B.n188 B.n187 585
R203 B.n186 B.n185 585
R204 B.n184 B.n183 585
R205 B.n182 B.n181 585
R206 B.n180 B.n179 585
R207 B.n178 B.n177 585
R208 B.n176 B.n175 585
R209 B.n174 B.n173 585
R210 B.n172 B.n171 585
R211 B.n170 B.n169 585
R212 B.n168 B.n167 585
R213 B.n166 B.n165 585
R214 B.n164 B.n163 585
R215 B.n162 B.n161 585
R216 B.n160 B.n159 585
R217 B.n158 B.n157 585
R218 B.n156 B.n155 585
R219 B.n124 B.n123 585
R220 B.n814 B.n813 585
R221 B.n807 B.n150 585
R222 B.n150 B.n121 585
R223 B.n806 B.n120 585
R224 B.n818 B.n120 585
R225 B.n805 B.n119 585
R226 B.n819 B.n119 585
R227 B.n804 B.n118 585
R228 B.n820 B.n118 585
R229 B.n803 B.n802 585
R230 B.n802 B.n114 585
R231 B.n801 B.n113 585
R232 B.n826 B.n113 585
R233 B.n800 B.n112 585
R234 B.n827 B.n112 585
R235 B.n799 B.n111 585
R236 B.n828 B.n111 585
R237 B.n798 B.n797 585
R238 B.n797 B.n107 585
R239 B.n796 B.n106 585
R240 B.n834 B.n106 585
R241 B.n795 B.n105 585
R242 B.n835 B.n105 585
R243 B.n794 B.n104 585
R244 B.n836 B.n104 585
R245 B.n793 B.n792 585
R246 B.n792 B.n100 585
R247 B.n791 B.n99 585
R248 B.n842 B.n99 585
R249 B.n790 B.n98 585
R250 B.n843 B.n98 585
R251 B.n789 B.n97 585
R252 B.n844 B.n97 585
R253 B.n788 B.n787 585
R254 B.n787 B.n93 585
R255 B.n786 B.n92 585
R256 B.n850 B.n92 585
R257 B.n785 B.n91 585
R258 B.n851 B.n91 585
R259 B.n784 B.n90 585
R260 B.n852 B.n90 585
R261 B.n783 B.n782 585
R262 B.n782 B.n86 585
R263 B.n781 B.n85 585
R264 B.n858 B.n85 585
R265 B.n780 B.n84 585
R266 B.n859 B.n84 585
R267 B.n779 B.n83 585
R268 B.n860 B.n83 585
R269 B.n778 B.n777 585
R270 B.n777 B.n82 585
R271 B.n776 B.n78 585
R272 B.n866 B.n78 585
R273 B.n775 B.n77 585
R274 B.n867 B.n77 585
R275 B.n774 B.n76 585
R276 B.n868 B.n76 585
R277 B.n773 B.n772 585
R278 B.n772 B.n72 585
R279 B.n771 B.n71 585
R280 B.n874 B.n71 585
R281 B.n770 B.n70 585
R282 B.n875 B.n70 585
R283 B.n769 B.n69 585
R284 B.n876 B.n69 585
R285 B.n768 B.n767 585
R286 B.n767 B.n65 585
R287 B.n766 B.n64 585
R288 B.n882 B.n64 585
R289 B.n765 B.n63 585
R290 B.n883 B.n63 585
R291 B.n764 B.n62 585
R292 B.n884 B.n62 585
R293 B.n763 B.n762 585
R294 B.n762 B.n61 585
R295 B.n761 B.n57 585
R296 B.n890 B.n57 585
R297 B.n760 B.n56 585
R298 B.n891 B.n56 585
R299 B.n759 B.n55 585
R300 B.n892 B.n55 585
R301 B.n758 B.n757 585
R302 B.n757 B.n51 585
R303 B.n756 B.n50 585
R304 B.n898 B.n50 585
R305 B.n755 B.n49 585
R306 B.n899 B.n49 585
R307 B.n754 B.n48 585
R308 B.n900 B.n48 585
R309 B.n753 B.n752 585
R310 B.n752 B.n44 585
R311 B.n751 B.n43 585
R312 B.n906 B.n43 585
R313 B.n750 B.n42 585
R314 B.n907 B.n42 585
R315 B.n749 B.n41 585
R316 B.n908 B.n41 585
R317 B.n748 B.n747 585
R318 B.n747 B.n40 585
R319 B.n746 B.n36 585
R320 B.n914 B.n36 585
R321 B.n745 B.n35 585
R322 B.n915 B.n35 585
R323 B.n744 B.n34 585
R324 B.n916 B.n34 585
R325 B.n743 B.n742 585
R326 B.n742 B.n30 585
R327 B.n741 B.n29 585
R328 B.n922 B.n29 585
R329 B.n740 B.n28 585
R330 B.n923 B.n28 585
R331 B.n739 B.n27 585
R332 B.n924 B.n27 585
R333 B.n738 B.n737 585
R334 B.n737 B.n23 585
R335 B.n736 B.n22 585
R336 B.n930 B.n22 585
R337 B.n735 B.n21 585
R338 B.n931 B.n21 585
R339 B.n734 B.n20 585
R340 B.n932 B.n20 585
R341 B.n733 B.n732 585
R342 B.n732 B.n16 585
R343 B.n731 B.n15 585
R344 B.n938 B.n15 585
R345 B.n730 B.n14 585
R346 B.n939 B.n14 585
R347 B.n729 B.n13 585
R348 B.n940 B.n13 585
R349 B.n728 B.n727 585
R350 B.n727 B.n12 585
R351 B.n726 B.n725 585
R352 B.n726 B.n8 585
R353 B.n724 B.n7 585
R354 B.n947 B.n7 585
R355 B.n723 B.n6 585
R356 B.n948 B.n6 585
R357 B.n722 B.n5 585
R358 B.n949 B.n5 585
R359 B.n721 B.n720 585
R360 B.n720 B.n4 585
R361 B.n719 B.n254 585
R362 B.n719 B.n718 585
R363 B.n709 B.n255 585
R364 B.n256 B.n255 585
R365 B.n711 B.n710 585
R366 B.n712 B.n711 585
R367 B.n708 B.n261 585
R368 B.n261 B.n260 585
R369 B.n707 B.n706 585
R370 B.n706 B.n705 585
R371 B.n263 B.n262 585
R372 B.n264 B.n263 585
R373 B.n698 B.n697 585
R374 B.n699 B.n698 585
R375 B.n696 B.n269 585
R376 B.n269 B.n268 585
R377 B.n695 B.n694 585
R378 B.n694 B.n693 585
R379 B.n271 B.n270 585
R380 B.n272 B.n271 585
R381 B.n686 B.n685 585
R382 B.n687 B.n686 585
R383 B.n684 B.n277 585
R384 B.n277 B.n276 585
R385 B.n683 B.n682 585
R386 B.n682 B.n681 585
R387 B.n279 B.n278 585
R388 B.n280 B.n279 585
R389 B.n674 B.n673 585
R390 B.n675 B.n674 585
R391 B.n672 B.n285 585
R392 B.n285 B.n284 585
R393 B.n671 B.n670 585
R394 B.n670 B.n669 585
R395 B.n287 B.n286 585
R396 B.n662 B.n287 585
R397 B.n661 B.n660 585
R398 B.n663 B.n661 585
R399 B.n659 B.n292 585
R400 B.n292 B.n291 585
R401 B.n658 B.n657 585
R402 B.n657 B.n656 585
R403 B.n294 B.n293 585
R404 B.n295 B.n294 585
R405 B.n649 B.n648 585
R406 B.n650 B.n649 585
R407 B.n647 B.n300 585
R408 B.n300 B.n299 585
R409 B.n646 B.n645 585
R410 B.n645 B.n644 585
R411 B.n302 B.n301 585
R412 B.n303 B.n302 585
R413 B.n637 B.n636 585
R414 B.n638 B.n637 585
R415 B.n635 B.n308 585
R416 B.n308 B.n307 585
R417 B.n634 B.n633 585
R418 B.n633 B.n632 585
R419 B.n310 B.n309 585
R420 B.n625 B.n310 585
R421 B.n624 B.n623 585
R422 B.n626 B.n624 585
R423 B.n622 B.n315 585
R424 B.n315 B.n314 585
R425 B.n621 B.n620 585
R426 B.n620 B.n619 585
R427 B.n317 B.n316 585
R428 B.n318 B.n317 585
R429 B.n612 B.n611 585
R430 B.n613 B.n612 585
R431 B.n610 B.n323 585
R432 B.n323 B.n322 585
R433 B.n609 B.n608 585
R434 B.n608 B.n607 585
R435 B.n325 B.n324 585
R436 B.n326 B.n325 585
R437 B.n600 B.n599 585
R438 B.n601 B.n600 585
R439 B.n598 B.n331 585
R440 B.n331 B.n330 585
R441 B.n597 B.n596 585
R442 B.n596 B.n595 585
R443 B.n333 B.n332 585
R444 B.n588 B.n333 585
R445 B.n587 B.n586 585
R446 B.n589 B.n587 585
R447 B.n585 B.n338 585
R448 B.n338 B.n337 585
R449 B.n584 B.n583 585
R450 B.n583 B.n582 585
R451 B.n340 B.n339 585
R452 B.n341 B.n340 585
R453 B.n575 B.n574 585
R454 B.n576 B.n575 585
R455 B.n573 B.n346 585
R456 B.n346 B.n345 585
R457 B.n572 B.n571 585
R458 B.n571 B.n570 585
R459 B.n348 B.n347 585
R460 B.n349 B.n348 585
R461 B.n563 B.n562 585
R462 B.n564 B.n563 585
R463 B.n561 B.n354 585
R464 B.n354 B.n353 585
R465 B.n560 B.n559 585
R466 B.n559 B.n558 585
R467 B.n356 B.n355 585
R468 B.n357 B.n356 585
R469 B.n551 B.n550 585
R470 B.n552 B.n551 585
R471 B.n549 B.n362 585
R472 B.n362 B.n361 585
R473 B.n548 B.n547 585
R474 B.n547 B.n546 585
R475 B.n364 B.n363 585
R476 B.n365 B.n364 585
R477 B.n539 B.n538 585
R478 B.n540 B.n539 585
R479 B.n537 B.n370 585
R480 B.n370 B.n369 585
R481 B.n536 B.n535 585
R482 B.n535 B.n534 585
R483 B.n372 B.n371 585
R484 B.n373 B.n372 585
R485 B.n527 B.n526 585
R486 B.n528 B.n527 585
R487 B.n525 B.n378 585
R488 B.n378 B.n377 585
R489 B.n524 B.n523 585
R490 B.n523 B.n522 585
R491 B.n380 B.n379 585
R492 B.n381 B.n380 585
R493 B.n518 B.n517 585
R494 B.n384 B.n383 585
R495 B.n514 B.n513 585
R496 B.n515 B.n514 585
R497 B.n512 B.n410 585
R498 B.n511 B.n510 585
R499 B.n509 B.n508 585
R500 B.n507 B.n506 585
R501 B.n505 B.n504 585
R502 B.n503 B.n502 585
R503 B.n501 B.n500 585
R504 B.n499 B.n498 585
R505 B.n497 B.n496 585
R506 B.n495 B.n494 585
R507 B.n493 B.n492 585
R508 B.n491 B.n490 585
R509 B.n489 B.n488 585
R510 B.n487 B.n486 585
R511 B.n485 B.n484 585
R512 B.n483 B.n482 585
R513 B.n481 B.n480 585
R514 B.n479 B.n478 585
R515 B.n477 B.n476 585
R516 B.n475 B.n474 585
R517 B.n473 B.n472 585
R518 B.n471 B.n470 585
R519 B.n469 B.n468 585
R520 B.n467 B.n466 585
R521 B.n465 B.n464 585
R522 B.n463 B.n462 585
R523 B.n461 B.n460 585
R524 B.n459 B.n458 585
R525 B.n457 B.n456 585
R526 B.n455 B.n454 585
R527 B.n453 B.n452 585
R528 B.n451 B.n450 585
R529 B.n449 B.n448 585
R530 B.n447 B.n446 585
R531 B.n445 B.n444 585
R532 B.n443 B.n442 585
R533 B.n441 B.n440 585
R534 B.n439 B.n438 585
R535 B.n437 B.n436 585
R536 B.n435 B.n434 585
R537 B.n433 B.n432 585
R538 B.n431 B.n430 585
R539 B.n429 B.n428 585
R540 B.n427 B.n426 585
R541 B.n425 B.n424 585
R542 B.n423 B.n422 585
R543 B.n421 B.n420 585
R544 B.n419 B.n418 585
R545 B.n417 B.n409 585
R546 B.n515 B.n409 585
R547 B.n519 B.n382 585
R548 B.n382 B.n381 585
R549 B.n521 B.n520 585
R550 B.n522 B.n521 585
R551 B.n376 B.n375 585
R552 B.n377 B.n376 585
R553 B.n530 B.n529 585
R554 B.n529 B.n528 585
R555 B.n531 B.n374 585
R556 B.n374 B.n373 585
R557 B.n533 B.n532 585
R558 B.n534 B.n533 585
R559 B.n368 B.n367 585
R560 B.n369 B.n368 585
R561 B.n542 B.n541 585
R562 B.n541 B.n540 585
R563 B.n543 B.n366 585
R564 B.n366 B.n365 585
R565 B.n545 B.n544 585
R566 B.n546 B.n545 585
R567 B.n360 B.n359 585
R568 B.n361 B.n360 585
R569 B.n554 B.n553 585
R570 B.n553 B.n552 585
R571 B.n555 B.n358 585
R572 B.n358 B.n357 585
R573 B.n557 B.n556 585
R574 B.n558 B.n557 585
R575 B.n352 B.n351 585
R576 B.n353 B.n352 585
R577 B.n566 B.n565 585
R578 B.n565 B.n564 585
R579 B.n567 B.n350 585
R580 B.n350 B.n349 585
R581 B.n569 B.n568 585
R582 B.n570 B.n569 585
R583 B.n344 B.n343 585
R584 B.n345 B.n344 585
R585 B.n578 B.n577 585
R586 B.n577 B.n576 585
R587 B.n579 B.n342 585
R588 B.n342 B.n341 585
R589 B.n581 B.n580 585
R590 B.n582 B.n581 585
R591 B.n336 B.n335 585
R592 B.n337 B.n336 585
R593 B.n591 B.n590 585
R594 B.n590 B.n589 585
R595 B.n592 B.n334 585
R596 B.n588 B.n334 585
R597 B.n594 B.n593 585
R598 B.n595 B.n594 585
R599 B.n329 B.n328 585
R600 B.n330 B.n329 585
R601 B.n603 B.n602 585
R602 B.n602 B.n601 585
R603 B.n604 B.n327 585
R604 B.n327 B.n326 585
R605 B.n606 B.n605 585
R606 B.n607 B.n606 585
R607 B.n321 B.n320 585
R608 B.n322 B.n321 585
R609 B.n615 B.n614 585
R610 B.n614 B.n613 585
R611 B.n616 B.n319 585
R612 B.n319 B.n318 585
R613 B.n618 B.n617 585
R614 B.n619 B.n618 585
R615 B.n313 B.n312 585
R616 B.n314 B.n313 585
R617 B.n628 B.n627 585
R618 B.n627 B.n626 585
R619 B.n629 B.n311 585
R620 B.n625 B.n311 585
R621 B.n631 B.n630 585
R622 B.n632 B.n631 585
R623 B.n306 B.n305 585
R624 B.n307 B.n306 585
R625 B.n640 B.n639 585
R626 B.n639 B.n638 585
R627 B.n641 B.n304 585
R628 B.n304 B.n303 585
R629 B.n643 B.n642 585
R630 B.n644 B.n643 585
R631 B.n298 B.n297 585
R632 B.n299 B.n298 585
R633 B.n652 B.n651 585
R634 B.n651 B.n650 585
R635 B.n653 B.n296 585
R636 B.n296 B.n295 585
R637 B.n655 B.n654 585
R638 B.n656 B.n655 585
R639 B.n290 B.n289 585
R640 B.n291 B.n290 585
R641 B.n665 B.n664 585
R642 B.n664 B.n663 585
R643 B.n666 B.n288 585
R644 B.n662 B.n288 585
R645 B.n668 B.n667 585
R646 B.n669 B.n668 585
R647 B.n283 B.n282 585
R648 B.n284 B.n283 585
R649 B.n677 B.n676 585
R650 B.n676 B.n675 585
R651 B.n678 B.n281 585
R652 B.n281 B.n280 585
R653 B.n680 B.n679 585
R654 B.n681 B.n680 585
R655 B.n275 B.n274 585
R656 B.n276 B.n275 585
R657 B.n689 B.n688 585
R658 B.n688 B.n687 585
R659 B.n690 B.n273 585
R660 B.n273 B.n272 585
R661 B.n692 B.n691 585
R662 B.n693 B.n692 585
R663 B.n267 B.n266 585
R664 B.n268 B.n267 585
R665 B.n701 B.n700 585
R666 B.n700 B.n699 585
R667 B.n702 B.n265 585
R668 B.n265 B.n264 585
R669 B.n704 B.n703 585
R670 B.n705 B.n704 585
R671 B.n259 B.n258 585
R672 B.n260 B.n259 585
R673 B.n714 B.n713 585
R674 B.n713 B.n712 585
R675 B.n715 B.n257 585
R676 B.n257 B.n256 585
R677 B.n717 B.n716 585
R678 B.n718 B.n717 585
R679 B.n3 B.n0 585
R680 B.n4 B.n3 585
R681 B.n946 B.n1 585
R682 B.n947 B.n946 585
R683 B.n945 B.n944 585
R684 B.n945 B.n8 585
R685 B.n943 B.n9 585
R686 B.n12 B.n9 585
R687 B.n942 B.n941 585
R688 B.n941 B.n940 585
R689 B.n11 B.n10 585
R690 B.n939 B.n11 585
R691 B.n937 B.n936 585
R692 B.n938 B.n937 585
R693 B.n935 B.n17 585
R694 B.n17 B.n16 585
R695 B.n934 B.n933 585
R696 B.n933 B.n932 585
R697 B.n19 B.n18 585
R698 B.n931 B.n19 585
R699 B.n929 B.n928 585
R700 B.n930 B.n929 585
R701 B.n927 B.n24 585
R702 B.n24 B.n23 585
R703 B.n926 B.n925 585
R704 B.n925 B.n924 585
R705 B.n26 B.n25 585
R706 B.n923 B.n26 585
R707 B.n921 B.n920 585
R708 B.n922 B.n921 585
R709 B.n919 B.n31 585
R710 B.n31 B.n30 585
R711 B.n918 B.n917 585
R712 B.n917 B.n916 585
R713 B.n33 B.n32 585
R714 B.n915 B.n33 585
R715 B.n913 B.n912 585
R716 B.n914 B.n913 585
R717 B.n911 B.n37 585
R718 B.n40 B.n37 585
R719 B.n910 B.n909 585
R720 B.n909 B.n908 585
R721 B.n39 B.n38 585
R722 B.n907 B.n39 585
R723 B.n905 B.n904 585
R724 B.n906 B.n905 585
R725 B.n903 B.n45 585
R726 B.n45 B.n44 585
R727 B.n902 B.n901 585
R728 B.n901 B.n900 585
R729 B.n47 B.n46 585
R730 B.n899 B.n47 585
R731 B.n897 B.n896 585
R732 B.n898 B.n897 585
R733 B.n895 B.n52 585
R734 B.n52 B.n51 585
R735 B.n894 B.n893 585
R736 B.n893 B.n892 585
R737 B.n54 B.n53 585
R738 B.n891 B.n54 585
R739 B.n889 B.n888 585
R740 B.n890 B.n889 585
R741 B.n887 B.n58 585
R742 B.n61 B.n58 585
R743 B.n886 B.n885 585
R744 B.n885 B.n884 585
R745 B.n60 B.n59 585
R746 B.n883 B.n60 585
R747 B.n881 B.n880 585
R748 B.n882 B.n881 585
R749 B.n879 B.n66 585
R750 B.n66 B.n65 585
R751 B.n878 B.n877 585
R752 B.n877 B.n876 585
R753 B.n68 B.n67 585
R754 B.n875 B.n68 585
R755 B.n873 B.n872 585
R756 B.n874 B.n873 585
R757 B.n871 B.n73 585
R758 B.n73 B.n72 585
R759 B.n870 B.n869 585
R760 B.n869 B.n868 585
R761 B.n75 B.n74 585
R762 B.n867 B.n75 585
R763 B.n865 B.n864 585
R764 B.n866 B.n865 585
R765 B.n863 B.n79 585
R766 B.n82 B.n79 585
R767 B.n862 B.n861 585
R768 B.n861 B.n860 585
R769 B.n81 B.n80 585
R770 B.n859 B.n81 585
R771 B.n857 B.n856 585
R772 B.n858 B.n857 585
R773 B.n855 B.n87 585
R774 B.n87 B.n86 585
R775 B.n854 B.n853 585
R776 B.n853 B.n852 585
R777 B.n89 B.n88 585
R778 B.n851 B.n89 585
R779 B.n849 B.n848 585
R780 B.n850 B.n849 585
R781 B.n847 B.n94 585
R782 B.n94 B.n93 585
R783 B.n846 B.n845 585
R784 B.n845 B.n844 585
R785 B.n96 B.n95 585
R786 B.n843 B.n96 585
R787 B.n841 B.n840 585
R788 B.n842 B.n841 585
R789 B.n839 B.n101 585
R790 B.n101 B.n100 585
R791 B.n838 B.n837 585
R792 B.n837 B.n836 585
R793 B.n103 B.n102 585
R794 B.n835 B.n103 585
R795 B.n833 B.n832 585
R796 B.n834 B.n833 585
R797 B.n831 B.n108 585
R798 B.n108 B.n107 585
R799 B.n830 B.n829 585
R800 B.n829 B.n828 585
R801 B.n110 B.n109 585
R802 B.n827 B.n110 585
R803 B.n825 B.n824 585
R804 B.n826 B.n825 585
R805 B.n823 B.n115 585
R806 B.n115 B.n114 585
R807 B.n822 B.n821 585
R808 B.n821 B.n820 585
R809 B.n117 B.n116 585
R810 B.n819 B.n117 585
R811 B.n817 B.n816 585
R812 B.n818 B.n817 585
R813 B.n815 B.n122 585
R814 B.n122 B.n121 585
R815 B.n950 B.n949 585
R816 B.n948 B.n2 585
R817 B.n813 B.n122 516.524
R818 B.n809 B.n150 516.524
R819 B.n409 B.n380 516.524
R820 B.n517 B.n382 516.524
R821 B.n811 B.n810 256.663
R822 B.n811 B.n148 256.663
R823 B.n811 B.n147 256.663
R824 B.n811 B.n146 256.663
R825 B.n811 B.n145 256.663
R826 B.n811 B.n144 256.663
R827 B.n811 B.n143 256.663
R828 B.n811 B.n142 256.663
R829 B.n811 B.n141 256.663
R830 B.n811 B.n140 256.663
R831 B.n811 B.n139 256.663
R832 B.n811 B.n138 256.663
R833 B.n811 B.n137 256.663
R834 B.n811 B.n136 256.663
R835 B.n811 B.n135 256.663
R836 B.n811 B.n134 256.663
R837 B.n811 B.n133 256.663
R838 B.n811 B.n132 256.663
R839 B.n811 B.n131 256.663
R840 B.n811 B.n130 256.663
R841 B.n811 B.n129 256.663
R842 B.n811 B.n128 256.663
R843 B.n811 B.n127 256.663
R844 B.n811 B.n126 256.663
R845 B.n811 B.n125 256.663
R846 B.n812 B.n811 256.663
R847 B.n516 B.n515 256.663
R848 B.n515 B.n385 256.663
R849 B.n515 B.n386 256.663
R850 B.n515 B.n387 256.663
R851 B.n515 B.n388 256.663
R852 B.n515 B.n389 256.663
R853 B.n515 B.n390 256.663
R854 B.n515 B.n391 256.663
R855 B.n515 B.n392 256.663
R856 B.n515 B.n393 256.663
R857 B.n515 B.n394 256.663
R858 B.n515 B.n395 256.663
R859 B.n515 B.n396 256.663
R860 B.n515 B.n397 256.663
R861 B.n515 B.n398 256.663
R862 B.n515 B.n399 256.663
R863 B.n515 B.n400 256.663
R864 B.n515 B.n401 256.663
R865 B.n515 B.n402 256.663
R866 B.n515 B.n403 256.663
R867 B.n515 B.n404 256.663
R868 B.n515 B.n405 256.663
R869 B.n515 B.n406 256.663
R870 B.n515 B.n407 256.663
R871 B.n515 B.n408 256.663
R872 B.n952 B.n951 256.663
R873 B.n153 B.t15 242.338
R874 B.n151 B.t19 242.338
R875 B.n414 B.t8 242.338
R876 B.n411 B.t12 242.338
R877 B.n155 B.n124 163.367
R878 B.n159 B.n158 163.367
R879 B.n163 B.n162 163.367
R880 B.n167 B.n166 163.367
R881 B.n171 B.n170 163.367
R882 B.n175 B.n174 163.367
R883 B.n179 B.n178 163.367
R884 B.n183 B.n182 163.367
R885 B.n187 B.n186 163.367
R886 B.n191 B.n190 163.367
R887 B.n196 B.n195 163.367
R888 B.n200 B.n199 163.367
R889 B.n204 B.n203 163.367
R890 B.n208 B.n207 163.367
R891 B.n212 B.n211 163.367
R892 B.n217 B.n216 163.367
R893 B.n221 B.n220 163.367
R894 B.n225 B.n224 163.367
R895 B.n229 B.n228 163.367
R896 B.n233 B.n232 163.367
R897 B.n237 B.n236 163.367
R898 B.n241 B.n240 163.367
R899 B.n245 B.n244 163.367
R900 B.n249 B.n248 163.367
R901 B.n251 B.n149 163.367
R902 B.n523 B.n380 163.367
R903 B.n523 B.n378 163.367
R904 B.n527 B.n378 163.367
R905 B.n527 B.n372 163.367
R906 B.n535 B.n372 163.367
R907 B.n535 B.n370 163.367
R908 B.n539 B.n370 163.367
R909 B.n539 B.n364 163.367
R910 B.n547 B.n364 163.367
R911 B.n547 B.n362 163.367
R912 B.n551 B.n362 163.367
R913 B.n551 B.n356 163.367
R914 B.n559 B.n356 163.367
R915 B.n559 B.n354 163.367
R916 B.n563 B.n354 163.367
R917 B.n563 B.n348 163.367
R918 B.n571 B.n348 163.367
R919 B.n571 B.n346 163.367
R920 B.n575 B.n346 163.367
R921 B.n575 B.n340 163.367
R922 B.n583 B.n340 163.367
R923 B.n583 B.n338 163.367
R924 B.n587 B.n338 163.367
R925 B.n587 B.n333 163.367
R926 B.n596 B.n333 163.367
R927 B.n596 B.n331 163.367
R928 B.n600 B.n331 163.367
R929 B.n600 B.n325 163.367
R930 B.n608 B.n325 163.367
R931 B.n608 B.n323 163.367
R932 B.n612 B.n323 163.367
R933 B.n612 B.n317 163.367
R934 B.n620 B.n317 163.367
R935 B.n620 B.n315 163.367
R936 B.n624 B.n315 163.367
R937 B.n624 B.n310 163.367
R938 B.n633 B.n310 163.367
R939 B.n633 B.n308 163.367
R940 B.n637 B.n308 163.367
R941 B.n637 B.n302 163.367
R942 B.n645 B.n302 163.367
R943 B.n645 B.n300 163.367
R944 B.n649 B.n300 163.367
R945 B.n649 B.n294 163.367
R946 B.n657 B.n294 163.367
R947 B.n657 B.n292 163.367
R948 B.n661 B.n292 163.367
R949 B.n661 B.n287 163.367
R950 B.n670 B.n287 163.367
R951 B.n670 B.n285 163.367
R952 B.n674 B.n285 163.367
R953 B.n674 B.n279 163.367
R954 B.n682 B.n279 163.367
R955 B.n682 B.n277 163.367
R956 B.n686 B.n277 163.367
R957 B.n686 B.n271 163.367
R958 B.n694 B.n271 163.367
R959 B.n694 B.n269 163.367
R960 B.n698 B.n269 163.367
R961 B.n698 B.n263 163.367
R962 B.n706 B.n263 163.367
R963 B.n706 B.n261 163.367
R964 B.n711 B.n261 163.367
R965 B.n711 B.n255 163.367
R966 B.n719 B.n255 163.367
R967 B.n720 B.n719 163.367
R968 B.n720 B.n5 163.367
R969 B.n6 B.n5 163.367
R970 B.n7 B.n6 163.367
R971 B.n726 B.n7 163.367
R972 B.n727 B.n726 163.367
R973 B.n727 B.n13 163.367
R974 B.n14 B.n13 163.367
R975 B.n15 B.n14 163.367
R976 B.n732 B.n15 163.367
R977 B.n732 B.n20 163.367
R978 B.n21 B.n20 163.367
R979 B.n22 B.n21 163.367
R980 B.n737 B.n22 163.367
R981 B.n737 B.n27 163.367
R982 B.n28 B.n27 163.367
R983 B.n29 B.n28 163.367
R984 B.n742 B.n29 163.367
R985 B.n742 B.n34 163.367
R986 B.n35 B.n34 163.367
R987 B.n36 B.n35 163.367
R988 B.n747 B.n36 163.367
R989 B.n747 B.n41 163.367
R990 B.n42 B.n41 163.367
R991 B.n43 B.n42 163.367
R992 B.n752 B.n43 163.367
R993 B.n752 B.n48 163.367
R994 B.n49 B.n48 163.367
R995 B.n50 B.n49 163.367
R996 B.n757 B.n50 163.367
R997 B.n757 B.n55 163.367
R998 B.n56 B.n55 163.367
R999 B.n57 B.n56 163.367
R1000 B.n762 B.n57 163.367
R1001 B.n762 B.n62 163.367
R1002 B.n63 B.n62 163.367
R1003 B.n64 B.n63 163.367
R1004 B.n767 B.n64 163.367
R1005 B.n767 B.n69 163.367
R1006 B.n70 B.n69 163.367
R1007 B.n71 B.n70 163.367
R1008 B.n772 B.n71 163.367
R1009 B.n772 B.n76 163.367
R1010 B.n77 B.n76 163.367
R1011 B.n78 B.n77 163.367
R1012 B.n777 B.n78 163.367
R1013 B.n777 B.n83 163.367
R1014 B.n84 B.n83 163.367
R1015 B.n85 B.n84 163.367
R1016 B.n782 B.n85 163.367
R1017 B.n782 B.n90 163.367
R1018 B.n91 B.n90 163.367
R1019 B.n92 B.n91 163.367
R1020 B.n787 B.n92 163.367
R1021 B.n787 B.n97 163.367
R1022 B.n98 B.n97 163.367
R1023 B.n99 B.n98 163.367
R1024 B.n792 B.n99 163.367
R1025 B.n792 B.n104 163.367
R1026 B.n105 B.n104 163.367
R1027 B.n106 B.n105 163.367
R1028 B.n797 B.n106 163.367
R1029 B.n797 B.n111 163.367
R1030 B.n112 B.n111 163.367
R1031 B.n113 B.n112 163.367
R1032 B.n802 B.n113 163.367
R1033 B.n802 B.n118 163.367
R1034 B.n119 B.n118 163.367
R1035 B.n120 B.n119 163.367
R1036 B.n150 B.n120 163.367
R1037 B.n514 B.n384 163.367
R1038 B.n514 B.n410 163.367
R1039 B.n510 B.n509 163.367
R1040 B.n506 B.n505 163.367
R1041 B.n502 B.n501 163.367
R1042 B.n498 B.n497 163.367
R1043 B.n494 B.n493 163.367
R1044 B.n490 B.n489 163.367
R1045 B.n486 B.n485 163.367
R1046 B.n482 B.n481 163.367
R1047 B.n478 B.n477 163.367
R1048 B.n474 B.n473 163.367
R1049 B.n470 B.n469 163.367
R1050 B.n466 B.n465 163.367
R1051 B.n462 B.n461 163.367
R1052 B.n458 B.n457 163.367
R1053 B.n454 B.n453 163.367
R1054 B.n450 B.n449 163.367
R1055 B.n446 B.n445 163.367
R1056 B.n442 B.n441 163.367
R1057 B.n438 B.n437 163.367
R1058 B.n434 B.n433 163.367
R1059 B.n430 B.n429 163.367
R1060 B.n426 B.n425 163.367
R1061 B.n422 B.n421 163.367
R1062 B.n418 B.n409 163.367
R1063 B.n521 B.n382 163.367
R1064 B.n521 B.n376 163.367
R1065 B.n529 B.n376 163.367
R1066 B.n529 B.n374 163.367
R1067 B.n533 B.n374 163.367
R1068 B.n533 B.n368 163.367
R1069 B.n541 B.n368 163.367
R1070 B.n541 B.n366 163.367
R1071 B.n545 B.n366 163.367
R1072 B.n545 B.n360 163.367
R1073 B.n553 B.n360 163.367
R1074 B.n553 B.n358 163.367
R1075 B.n557 B.n358 163.367
R1076 B.n557 B.n352 163.367
R1077 B.n565 B.n352 163.367
R1078 B.n565 B.n350 163.367
R1079 B.n569 B.n350 163.367
R1080 B.n569 B.n344 163.367
R1081 B.n577 B.n344 163.367
R1082 B.n577 B.n342 163.367
R1083 B.n581 B.n342 163.367
R1084 B.n581 B.n336 163.367
R1085 B.n590 B.n336 163.367
R1086 B.n590 B.n334 163.367
R1087 B.n594 B.n334 163.367
R1088 B.n594 B.n329 163.367
R1089 B.n602 B.n329 163.367
R1090 B.n602 B.n327 163.367
R1091 B.n606 B.n327 163.367
R1092 B.n606 B.n321 163.367
R1093 B.n614 B.n321 163.367
R1094 B.n614 B.n319 163.367
R1095 B.n618 B.n319 163.367
R1096 B.n618 B.n313 163.367
R1097 B.n627 B.n313 163.367
R1098 B.n627 B.n311 163.367
R1099 B.n631 B.n311 163.367
R1100 B.n631 B.n306 163.367
R1101 B.n639 B.n306 163.367
R1102 B.n639 B.n304 163.367
R1103 B.n643 B.n304 163.367
R1104 B.n643 B.n298 163.367
R1105 B.n651 B.n298 163.367
R1106 B.n651 B.n296 163.367
R1107 B.n655 B.n296 163.367
R1108 B.n655 B.n290 163.367
R1109 B.n664 B.n290 163.367
R1110 B.n664 B.n288 163.367
R1111 B.n668 B.n288 163.367
R1112 B.n668 B.n283 163.367
R1113 B.n676 B.n283 163.367
R1114 B.n676 B.n281 163.367
R1115 B.n680 B.n281 163.367
R1116 B.n680 B.n275 163.367
R1117 B.n688 B.n275 163.367
R1118 B.n688 B.n273 163.367
R1119 B.n692 B.n273 163.367
R1120 B.n692 B.n267 163.367
R1121 B.n700 B.n267 163.367
R1122 B.n700 B.n265 163.367
R1123 B.n704 B.n265 163.367
R1124 B.n704 B.n259 163.367
R1125 B.n713 B.n259 163.367
R1126 B.n713 B.n257 163.367
R1127 B.n717 B.n257 163.367
R1128 B.n717 B.n3 163.367
R1129 B.n950 B.n3 163.367
R1130 B.n946 B.n2 163.367
R1131 B.n946 B.n945 163.367
R1132 B.n945 B.n9 163.367
R1133 B.n941 B.n9 163.367
R1134 B.n941 B.n11 163.367
R1135 B.n937 B.n11 163.367
R1136 B.n937 B.n17 163.367
R1137 B.n933 B.n17 163.367
R1138 B.n933 B.n19 163.367
R1139 B.n929 B.n19 163.367
R1140 B.n929 B.n24 163.367
R1141 B.n925 B.n24 163.367
R1142 B.n925 B.n26 163.367
R1143 B.n921 B.n26 163.367
R1144 B.n921 B.n31 163.367
R1145 B.n917 B.n31 163.367
R1146 B.n917 B.n33 163.367
R1147 B.n913 B.n33 163.367
R1148 B.n913 B.n37 163.367
R1149 B.n909 B.n37 163.367
R1150 B.n909 B.n39 163.367
R1151 B.n905 B.n39 163.367
R1152 B.n905 B.n45 163.367
R1153 B.n901 B.n45 163.367
R1154 B.n901 B.n47 163.367
R1155 B.n897 B.n47 163.367
R1156 B.n897 B.n52 163.367
R1157 B.n893 B.n52 163.367
R1158 B.n893 B.n54 163.367
R1159 B.n889 B.n54 163.367
R1160 B.n889 B.n58 163.367
R1161 B.n885 B.n58 163.367
R1162 B.n885 B.n60 163.367
R1163 B.n881 B.n60 163.367
R1164 B.n881 B.n66 163.367
R1165 B.n877 B.n66 163.367
R1166 B.n877 B.n68 163.367
R1167 B.n873 B.n68 163.367
R1168 B.n873 B.n73 163.367
R1169 B.n869 B.n73 163.367
R1170 B.n869 B.n75 163.367
R1171 B.n865 B.n75 163.367
R1172 B.n865 B.n79 163.367
R1173 B.n861 B.n79 163.367
R1174 B.n861 B.n81 163.367
R1175 B.n857 B.n81 163.367
R1176 B.n857 B.n87 163.367
R1177 B.n853 B.n87 163.367
R1178 B.n853 B.n89 163.367
R1179 B.n849 B.n89 163.367
R1180 B.n849 B.n94 163.367
R1181 B.n845 B.n94 163.367
R1182 B.n845 B.n96 163.367
R1183 B.n841 B.n96 163.367
R1184 B.n841 B.n101 163.367
R1185 B.n837 B.n101 163.367
R1186 B.n837 B.n103 163.367
R1187 B.n833 B.n103 163.367
R1188 B.n833 B.n108 163.367
R1189 B.n829 B.n108 163.367
R1190 B.n829 B.n110 163.367
R1191 B.n825 B.n110 163.367
R1192 B.n825 B.n115 163.367
R1193 B.n821 B.n115 163.367
R1194 B.n821 B.n117 163.367
R1195 B.n817 B.n117 163.367
R1196 B.n817 B.n122 163.367
R1197 B.n151 B.t20 154.869
R1198 B.n414 B.t11 154.869
R1199 B.n153 B.t17 154.864
R1200 B.n411 B.t14 154.864
R1201 B.n515 B.n381 132.659
R1202 B.n811 B.n121 132.659
R1203 B.n154 B.n153 78.352
R1204 B.n152 B.n151 78.352
R1205 B.n415 B.n414 78.352
R1206 B.n412 B.n411 78.352
R1207 B.n152 B.t21 76.5179
R1208 B.n415 B.t10 76.5179
R1209 B.n154 B.t18 76.5131
R1210 B.n412 B.t13 76.5131
R1211 B.n522 B.n381 72.1664
R1212 B.n522 B.n377 72.1664
R1213 B.n528 B.n377 72.1664
R1214 B.n528 B.n373 72.1664
R1215 B.n534 B.n373 72.1664
R1216 B.n534 B.n369 72.1664
R1217 B.n540 B.n369 72.1664
R1218 B.n540 B.n365 72.1664
R1219 B.n546 B.n365 72.1664
R1220 B.n552 B.n361 72.1664
R1221 B.n552 B.n357 72.1664
R1222 B.n558 B.n357 72.1664
R1223 B.n558 B.n353 72.1664
R1224 B.n564 B.n353 72.1664
R1225 B.n564 B.n349 72.1664
R1226 B.n570 B.n349 72.1664
R1227 B.n570 B.n345 72.1664
R1228 B.n576 B.n345 72.1664
R1229 B.n576 B.n341 72.1664
R1230 B.n582 B.n341 72.1664
R1231 B.n582 B.n337 72.1664
R1232 B.n589 B.n337 72.1664
R1233 B.n589 B.n588 72.1664
R1234 B.n595 B.n330 72.1664
R1235 B.n601 B.n330 72.1664
R1236 B.n601 B.n326 72.1664
R1237 B.n607 B.n326 72.1664
R1238 B.n607 B.n322 72.1664
R1239 B.n613 B.n322 72.1664
R1240 B.n613 B.n318 72.1664
R1241 B.n619 B.n318 72.1664
R1242 B.n619 B.n314 72.1664
R1243 B.n626 B.n314 72.1664
R1244 B.n626 B.n625 72.1664
R1245 B.n632 B.n307 72.1664
R1246 B.n638 B.n307 72.1664
R1247 B.n638 B.n303 72.1664
R1248 B.n644 B.n303 72.1664
R1249 B.n644 B.n299 72.1664
R1250 B.n650 B.n299 72.1664
R1251 B.n650 B.n295 72.1664
R1252 B.n656 B.n295 72.1664
R1253 B.n656 B.n291 72.1664
R1254 B.n663 B.n291 72.1664
R1255 B.n663 B.n662 72.1664
R1256 B.n669 B.n284 72.1664
R1257 B.n675 B.n284 72.1664
R1258 B.n675 B.n280 72.1664
R1259 B.n681 B.n280 72.1664
R1260 B.n681 B.n276 72.1664
R1261 B.n687 B.n276 72.1664
R1262 B.n687 B.n272 72.1664
R1263 B.n693 B.n272 72.1664
R1264 B.n693 B.n268 72.1664
R1265 B.n699 B.n268 72.1664
R1266 B.n705 B.n264 72.1664
R1267 B.n705 B.n260 72.1664
R1268 B.n712 B.n260 72.1664
R1269 B.n712 B.n256 72.1664
R1270 B.n718 B.n256 72.1664
R1271 B.n718 B.n4 72.1664
R1272 B.n949 B.n4 72.1664
R1273 B.n949 B.n948 72.1664
R1274 B.n948 B.n947 72.1664
R1275 B.n947 B.n8 72.1664
R1276 B.n12 B.n8 72.1664
R1277 B.n940 B.n12 72.1664
R1278 B.n940 B.n939 72.1664
R1279 B.n939 B.n938 72.1664
R1280 B.n938 B.n16 72.1664
R1281 B.n932 B.n931 72.1664
R1282 B.n931 B.n930 72.1664
R1283 B.n930 B.n23 72.1664
R1284 B.n924 B.n23 72.1664
R1285 B.n924 B.n923 72.1664
R1286 B.n923 B.n922 72.1664
R1287 B.n922 B.n30 72.1664
R1288 B.n916 B.n30 72.1664
R1289 B.n916 B.n915 72.1664
R1290 B.n915 B.n914 72.1664
R1291 B.n908 B.n40 72.1664
R1292 B.n908 B.n907 72.1664
R1293 B.n907 B.n906 72.1664
R1294 B.n906 B.n44 72.1664
R1295 B.n900 B.n44 72.1664
R1296 B.n900 B.n899 72.1664
R1297 B.n899 B.n898 72.1664
R1298 B.n898 B.n51 72.1664
R1299 B.n892 B.n51 72.1664
R1300 B.n892 B.n891 72.1664
R1301 B.n891 B.n890 72.1664
R1302 B.n884 B.n61 72.1664
R1303 B.n884 B.n883 72.1664
R1304 B.n883 B.n882 72.1664
R1305 B.n882 B.n65 72.1664
R1306 B.n876 B.n65 72.1664
R1307 B.n876 B.n875 72.1664
R1308 B.n875 B.n874 72.1664
R1309 B.n874 B.n72 72.1664
R1310 B.n868 B.n72 72.1664
R1311 B.n868 B.n867 72.1664
R1312 B.n867 B.n866 72.1664
R1313 B.n860 B.n82 72.1664
R1314 B.n860 B.n859 72.1664
R1315 B.n859 B.n858 72.1664
R1316 B.n858 B.n86 72.1664
R1317 B.n852 B.n86 72.1664
R1318 B.n852 B.n851 72.1664
R1319 B.n851 B.n850 72.1664
R1320 B.n850 B.n93 72.1664
R1321 B.n844 B.n93 72.1664
R1322 B.n844 B.n843 72.1664
R1323 B.n843 B.n842 72.1664
R1324 B.n842 B.n100 72.1664
R1325 B.n836 B.n100 72.1664
R1326 B.n836 B.n835 72.1664
R1327 B.n834 B.n107 72.1664
R1328 B.n828 B.n107 72.1664
R1329 B.n828 B.n827 72.1664
R1330 B.n827 B.n826 72.1664
R1331 B.n826 B.n114 72.1664
R1332 B.n820 B.n114 72.1664
R1333 B.n820 B.n819 72.1664
R1334 B.n819 B.n818 72.1664
R1335 B.n818 B.n121 72.1664
R1336 B.n813 B.n812 71.676
R1337 B.n155 B.n125 71.676
R1338 B.n159 B.n126 71.676
R1339 B.n163 B.n127 71.676
R1340 B.n167 B.n128 71.676
R1341 B.n171 B.n129 71.676
R1342 B.n175 B.n130 71.676
R1343 B.n179 B.n131 71.676
R1344 B.n183 B.n132 71.676
R1345 B.n187 B.n133 71.676
R1346 B.n191 B.n134 71.676
R1347 B.n196 B.n135 71.676
R1348 B.n200 B.n136 71.676
R1349 B.n204 B.n137 71.676
R1350 B.n208 B.n138 71.676
R1351 B.n212 B.n139 71.676
R1352 B.n217 B.n140 71.676
R1353 B.n221 B.n141 71.676
R1354 B.n225 B.n142 71.676
R1355 B.n229 B.n143 71.676
R1356 B.n233 B.n144 71.676
R1357 B.n237 B.n145 71.676
R1358 B.n241 B.n146 71.676
R1359 B.n245 B.n147 71.676
R1360 B.n249 B.n148 71.676
R1361 B.n810 B.n149 71.676
R1362 B.n810 B.n809 71.676
R1363 B.n251 B.n148 71.676
R1364 B.n248 B.n147 71.676
R1365 B.n244 B.n146 71.676
R1366 B.n240 B.n145 71.676
R1367 B.n236 B.n144 71.676
R1368 B.n232 B.n143 71.676
R1369 B.n228 B.n142 71.676
R1370 B.n224 B.n141 71.676
R1371 B.n220 B.n140 71.676
R1372 B.n216 B.n139 71.676
R1373 B.n211 B.n138 71.676
R1374 B.n207 B.n137 71.676
R1375 B.n203 B.n136 71.676
R1376 B.n199 B.n135 71.676
R1377 B.n195 B.n134 71.676
R1378 B.n190 B.n133 71.676
R1379 B.n186 B.n132 71.676
R1380 B.n182 B.n131 71.676
R1381 B.n178 B.n130 71.676
R1382 B.n174 B.n129 71.676
R1383 B.n170 B.n128 71.676
R1384 B.n166 B.n127 71.676
R1385 B.n162 B.n126 71.676
R1386 B.n158 B.n125 71.676
R1387 B.n812 B.n124 71.676
R1388 B.n517 B.n516 71.676
R1389 B.n410 B.n385 71.676
R1390 B.n509 B.n386 71.676
R1391 B.n505 B.n387 71.676
R1392 B.n501 B.n388 71.676
R1393 B.n497 B.n389 71.676
R1394 B.n493 B.n390 71.676
R1395 B.n489 B.n391 71.676
R1396 B.n485 B.n392 71.676
R1397 B.n481 B.n393 71.676
R1398 B.n477 B.n394 71.676
R1399 B.n473 B.n395 71.676
R1400 B.n469 B.n396 71.676
R1401 B.n465 B.n397 71.676
R1402 B.n461 B.n398 71.676
R1403 B.n457 B.n399 71.676
R1404 B.n453 B.n400 71.676
R1405 B.n449 B.n401 71.676
R1406 B.n445 B.n402 71.676
R1407 B.n441 B.n403 71.676
R1408 B.n437 B.n404 71.676
R1409 B.n433 B.n405 71.676
R1410 B.n429 B.n406 71.676
R1411 B.n425 B.n407 71.676
R1412 B.n421 B.n408 71.676
R1413 B.n516 B.n384 71.676
R1414 B.n510 B.n385 71.676
R1415 B.n506 B.n386 71.676
R1416 B.n502 B.n387 71.676
R1417 B.n498 B.n388 71.676
R1418 B.n494 B.n389 71.676
R1419 B.n490 B.n390 71.676
R1420 B.n486 B.n391 71.676
R1421 B.n482 B.n392 71.676
R1422 B.n478 B.n393 71.676
R1423 B.n474 B.n394 71.676
R1424 B.n470 B.n395 71.676
R1425 B.n466 B.n396 71.676
R1426 B.n462 B.n397 71.676
R1427 B.n458 B.n398 71.676
R1428 B.n454 B.n399 71.676
R1429 B.n450 B.n400 71.676
R1430 B.n446 B.n401 71.676
R1431 B.n442 B.n402 71.676
R1432 B.n438 B.n403 71.676
R1433 B.n434 B.n404 71.676
R1434 B.n430 B.n405 71.676
R1435 B.n426 B.n406 71.676
R1436 B.n422 B.n407 71.676
R1437 B.n418 B.n408 71.676
R1438 B.n951 B.n950 71.676
R1439 B.n951 B.n2 71.676
R1440 B.n699 B.t7 68.9826
R1441 B.n932 B.t3 68.9826
R1442 B.n669 B.t2 66.8601
R1443 B.n914 B.t1 66.8601
R1444 B.n193 B.n154 59.5399
R1445 B.n214 B.n152 59.5399
R1446 B.n416 B.n415 59.5399
R1447 B.n413 B.n412 59.5399
R1448 B.n632 B.t5 58.37
R1449 B.n890 B.t0 58.37
R1450 B.t9 B.n361 56.2475
R1451 B.n835 B.t16 56.2475
R1452 B.n595 B.t4 49.8799
R1453 B.n866 B.t6 49.8799
R1454 B.n519 B.n518 33.5615
R1455 B.n417 B.n379 33.5615
R1456 B.n808 B.n807 33.5615
R1457 B.n815 B.n814 33.5615
R1458 B.n588 B.t4 22.287
R1459 B.n82 B.t6 22.287
R1460 B B.n952 18.0485
R1461 B.n546 B.t9 15.9195
R1462 B.t16 B.n834 15.9195
R1463 B.n625 B.t5 13.7969
R1464 B.n61 B.t0 13.7969
R1465 B.n520 B.n519 10.6151
R1466 B.n520 B.n375 10.6151
R1467 B.n530 B.n375 10.6151
R1468 B.n531 B.n530 10.6151
R1469 B.n532 B.n531 10.6151
R1470 B.n532 B.n367 10.6151
R1471 B.n542 B.n367 10.6151
R1472 B.n543 B.n542 10.6151
R1473 B.n544 B.n543 10.6151
R1474 B.n544 B.n359 10.6151
R1475 B.n554 B.n359 10.6151
R1476 B.n555 B.n554 10.6151
R1477 B.n556 B.n555 10.6151
R1478 B.n556 B.n351 10.6151
R1479 B.n566 B.n351 10.6151
R1480 B.n567 B.n566 10.6151
R1481 B.n568 B.n567 10.6151
R1482 B.n568 B.n343 10.6151
R1483 B.n578 B.n343 10.6151
R1484 B.n579 B.n578 10.6151
R1485 B.n580 B.n579 10.6151
R1486 B.n580 B.n335 10.6151
R1487 B.n591 B.n335 10.6151
R1488 B.n592 B.n591 10.6151
R1489 B.n593 B.n592 10.6151
R1490 B.n593 B.n328 10.6151
R1491 B.n603 B.n328 10.6151
R1492 B.n604 B.n603 10.6151
R1493 B.n605 B.n604 10.6151
R1494 B.n605 B.n320 10.6151
R1495 B.n615 B.n320 10.6151
R1496 B.n616 B.n615 10.6151
R1497 B.n617 B.n616 10.6151
R1498 B.n617 B.n312 10.6151
R1499 B.n628 B.n312 10.6151
R1500 B.n629 B.n628 10.6151
R1501 B.n630 B.n629 10.6151
R1502 B.n630 B.n305 10.6151
R1503 B.n640 B.n305 10.6151
R1504 B.n641 B.n640 10.6151
R1505 B.n642 B.n641 10.6151
R1506 B.n642 B.n297 10.6151
R1507 B.n652 B.n297 10.6151
R1508 B.n653 B.n652 10.6151
R1509 B.n654 B.n653 10.6151
R1510 B.n654 B.n289 10.6151
R1511 B.n665 B.n289 10.6151
R1512 B.n666 B.n665 10.6151
R1513 B.n667 B.n666 10.6151
R1514 B.n667 B.n282 10.6151
R1515 B.n677 B.n282 10.6151
R1516 B.n678 B.n677 10.6151
R1517 B.n679 B.n678 10.6151
R1518 B.n679 B.n274 10.6151
R1519 B.n689 B.n274 10.6151
R1520 B.n690 B.n689 10.6151
R1521 B.n691 B.n690 10.6151
R1522 B.n691 B.n266 10.6151
R1523 B.n701 B.n266 10.6151
R1524 B.n702 B.n701 10.6151
R1525 B.n703 B.n702 10.6151
R1526 B.n703 B.n258 10.6151
R1527 B.n714 B.n258 10.6151
R1528 B.n715 B.n714 10.6151
R1529 B.n716 B.n715 10.6151
R1530 B.n716 B.n0 10.6151
R1531 B.n518 B.n383 10.6151
R1532 B.n513 B.n383 10.6151
R1533 B.n513 B.n512 10.6151
R1534 B.n512 B.n511 10.6151
R1535 B.n511 B.n508 10.6151
R1536 B.n508 B.n507 10.6151
R1537 B.n507 B.n504 10.6151
R1538 B.n504 B.n503 10.6151
R1539 B.n503 B.n500 10.6151
R1540 B.n500 B.n499 10.6151
R1541 B.n499 B.n496 10.6151
R1542 B.n496 B.n495 10.6151
R1543 B.n495 B.n492 10.6151
R1544 B.n492 B.n491 10.6151
R1545 B.n491 B.n488 10.6151
R1546 B.n488 B.n487 10.6151
R1547 B.n487 B.n484 10.6151
R1548 B.n484 B.n483 10.6151
R1549 B.n483 B.n480 10.6151
R1550 B.n480 B.n479 10.6151
R1551 B.n476 B.n475 10.6151
R1552 B.n475 B.n472 10.6151
R1553 B.n472 B.n471 10.6151
R1554 B.n471 B.n468 10.6151
R1555 B.n468 B.n467 10.6151
R1556 B.n467 B.n464 10.6151
R1557 B.n464 B.n463 10.6151
R1558 B.n463 B.n460 10.6151
R1559 B.n460 B.n459 10.6151
R1560 B.n456 B.n455 10.6151
R1561 B.n455 B.n452 10.6151
R1562 B.n452 B.n451 10.6151
R1563 B.n451 B.n448 10.6151
R1564 B.n448 B.n447 10.6151
R1565 B.n447 B.n444 10.6151
R1566 B.n444 B.n443 10.6151
R1567 B.n443 B.n440 10.6151
R1568 B.n440 B.n439 10.6151
R1569 B.n439 B.n436 10.6151
R1570 B.n436 B.n435 10.6151
R1571 B.n435 B.n432 10.6151
R1572 B.n432 B.n431 10.6151
R1573 B.n431 B.n428 10.6151
R1574 B.n428 B.n427 10.6151
R1575 B.n427 B.n424 10.6151
R1576 B.n424 B.n423 10.6151
R1577 B.n423 B.n420 10.6151
R1578 B.n420 B.n419 10.6151
R1579 B.n419 B.n417 10.6151
R1580 B.n524 B.n379 10.6151
R1581 B.n525 B.n524 10.6151
R1582 B.n526 B.n525 10.6151
R1583 B.n526 B.n371 10.6151
R1584 B.n536 B.n371 10.6151
R1585 B.n537 B.n536 10.6151
R1586 B.n538 B.n537 10.6151
R1587 B.n538 B.n363 10.6151
R1588 B.n548 B.n363 10.6151
R1589 B.n549 B.n548 10.6151
R1590 B.n550 B.n549 10.6151
R1591 B.n550 B.n355 10.6151
R1592 B.n560 B.n355 10.6151
R1593 B.n561 B.n560 10.6151
R1594 B.n562 B.n561 10.6151
R1595 B.n562 B.n347 10.6151
R1596 B.n572 B.n347 10.6151
R1597 B.n573 B.n572 10.6151
R1598 B.n574 B.n573 10.6151
R1599 B.n574 B.n339 10.6151
R1600 B.n584 B.n339 10.6151
R1601 B.n585 B.n584 10.6151
R1602 B.n586 B.n585 10.6151
R1603 B.n586 B.n332 10.6151
R1604 B.n597 B.n332 10.6151
R1605 B.n598 B.n597 10.6151
R1606 B.n599 B.n598 10.6151
R1607 B.n599 B.n324 10.6151
R1608 B.n609 B.n324 10.6151
R1609 B.n610 B.n609 10.6151
R1610 B.n611 B.n610 10.6151
R1611 B.n611 B.n316 10.6151
R1612 B.n621 B.n316 10.6151
R1613 B.n622 B.n621 10.6151
R1614 B.n623 B.n622 10.6151
R1615 B.n623 B.n309 10.6151
R1616 B.n634 B.n309 10.6151
R1617 B.n635 B.n634 10.6151
R1618 B.n636 B.n635 10.6151
R1619 B.n636 B.n301 10.6151
R1620 B.n646 B.n301 10.6151
R1621 B.n647 B.n646 10.6151
R1622 B.n648 B.n647 10.6151
R1623 B.n648 B.n293 10.6151
R1624 B.n658 B.n293 10.6151
R1625 B.n659 B.n658 10.6151
R1626 B.n660 B.n659 10.6151
R1627 B.n660 B.n286 10.6151
R1628 B.n671 B.n286 10.6151
R1629 B.n672 B.n671 10.6151
R1630 B.n673 B.n672 10.6151
R1631 B.n673 B.n278 10.6151
R1632 B.n683 B.n278 10.6151
R1633 B.n684 B.n683 10.6151
R1634 B.n685 B.n684 10.6151
R1635 B.n685 B.n270 10.6151
R1636 B.n695 B.n270 10.6151
R1637 B.n696 B.n695 10.6151
R1638 B.n697 B.n696 10.6151
R1639 B.n697 B.n262 10.6151
R1640 B.n707 B.n262 10.6151
R1641 B.n708 B.n707 10.6151
R1642 B.n710 B.n708 10.6151
R1643 B.n710 B.n709 10.6151
R1644 B.n709 B.n254 10.6151
R1645 B.n721 B.n254 10.6151
R1646 B.n722 B.n721 10.6151
R1647 B.n723 B.n722 10.6151
R1648 B.n724 B.n723 10.6151
R1649 B.n725 B.n724 10.6151
R1650 B.n728 B.n725 10.6151
R1651 B.n729 B.n728 10.6151
R1652 B.n730 B.n729 10.6151
R1653 B.n731 B.n730 10.6151
R1654 B.n733 B.n731 10.6151
R1655 B.n734 B.n733 10.6151
R1656 B.n735 B.n734 10.6151
R1657 B.n736 B.n735 10.6151
R1658 B.n738 B.n736 10.6151
R1659 B.n739 B.n738 10.6151
R1660 B.n740 B.n739 10.6151
R1661 B.n741 B.n740 10.6151
R1662 B.n743 B.n741 10.6151
R1663 B.n744 B.n743 10.6151
R1664 B.n745 B.n744 10.6151
R1665 B.n746 B.n745 10.6151
R1666 B.n748 B.n746 10.6151
R1667 B.n749 B.n748 10.6151
R1668 B.n750 B.n749 10.6151
R1669 B.n751 B.n750 10.6151
R1670 B.n753 B.n751 10.6151
R1671 B.n754 B.n753 10.6151
R1672 B.n755 B.n754 10.6151
R1673 B.n756 B.n755 10.6151
R1674 B.n758 B.n756 10.6151
R1675 B.n759 B.n758 10.6151
R1676 B.n760 B.n759 10.6151
R1677 B.n761 B.n760 10.6151
R1678 B.n763 B.n761 10.6151
R1679 B.n764 B.n763 10.6151
R1680 B.n765 B.n764 10.6151
R1681 B.n766 B.n765 10.6151
R1682 B.n768 B.n766 10.6151
R1683 B.n769 B.n768 10.6151
R1684 B.n770 B.n769 10.6151
R1685 B.n771 B.n770 10.6151
R1686 B.n773 B.n771 10.6151
R1687 B.n774 B.n773 10.6151
R1688 B.n775 B.n774 10.6151
R1689 B.n776 B.n775 10.6151
R1690 B.n778 B.n776 10.6151
R1691 B.n779 B.n778 10.6151
R1692 B.n780 B.n779 10.6151
R1693 B.n781 B.n780 10.6151
R1694 B.n783 B.n781 10.6151
R1695 B.n784 B.n783 10.6151
R1696 B.n785 B.n784 10.6151
R1697 B.n786 B.n785 10.6151
R1698 B.n788 B.n786 10.6151
R1699 B.n789 B.n788 10.6151
R1700 B.n790 B.n789 10.6151
R1701 B.n791 B.n790 10.6151
R1702 B.n793 B.n791 10.6151
R1703 B.n794 B.n793 10.6151
R1704 B.n795 B.n794 10.6151
R1705 B.n796 B.n795 10.6151
R1706 B.n798 B.n796 10.6151
R1707 B.n799 B.n798 10.6151
R1708 B.n800 B.n799 10.6151
R1709 B.n801 B.n800 10.6151
R1710 B.n803 B.n801 10.6151
R1711 B.n804 B.n803 10.6151
R1712 B.n805 B.n804 10.6151
R1713 B.n806 B.n805 10.6151
R1714 B.n807 B.n806 10.6151
R1715 B.n944 B.n1 10.6151
R1716 B.n944 B.n943 10.6151
R1717 B.n943 B.n942 10.6151
R1718 B.n942 B.n10 10.6151
R1719 B.n936 B.n10 10.6151
R1720 B.n936 B.n935 10.6151
R1721 B.n935 B.n934 10.6151
R1722 B.n934 B.n18 10.6151
R1723 B.n928 B.n18 10.6151
R1724 B.n928 B.n927 10.6151
R1725 B.n927 B.n926 10.6151
R1726 B.n926 B.n25 10.6151
R1727 B.n920 B.n25 10.6151
R1728 B.n920 B.n919 10.6151
R1729 B.n919 B.n918 10.6151
R1730 B.n918 B.n32 10.6151
R1731 B.n912 B.n32 10.6151
R1732 B.n912 B.n911 10.6151
R1733 B.n911 B.n910 10.6151
R1734 B.n910 B.n38 10.6151
R1735 B.n904 B.n38 10.6151
R1736 B.n904 B.n903 10.6151
R1737 B.n903 B.n902 10.6151
R1738 B.n902 B.n46 10.6151
R1739 B.n896 B.n46 10.6151
R1740 B.n896 B.n895 10.6151
R1741 B.n895 B.n894 10.6151
R1742 B.n894 B.n53 10.6151
R1743 B.n888 B.n53 10.6151
R1744 B.n888 B.n887 10.6151
R1745 B.n887 B.n886 10.6151
R1746 B.n886 B.n59 10.6151
R1747 B.n880 B.n59 10.6151
R1748 B.n880 B.n879 10.6151
R1749 B.n879 B.n878 10.6151
R1750 B.n878 B.n67 10.6151
R1751 B.n872 B.n67 10.6151
R1752 B.n872 B.n871 10.6151
R1753 B.n871 B.n870 10.6151
R1754 B.n870 B.n74 10.6151
R1755 B.n864 B.n74 10.6151
R1756 B.n864 B.n863 10.6151
R1757 B.n863 B.n862 10.6151
R1758 B.n862 B.n80 10.6151
R1759 B.n856 B.n80 10.6151
R1760 B.n856 B.n855 10.6151
R1761 B.n855 B.n854 10.6151
R1762 B.n854 B.n88 10.6151
R1763 B.n848 B.n88 10.6151
R1764 B.n848 B.n847 10.6151
R1765 B.n847 B.n846 10.6151
R1766 B.n846 B.n95 10.6151
R1767 B.n840 B.n95 10.6151
R1768 B.n840 B.n839 10.6151
R1769 B.n839 B.n838 10.6151
R1770 B.n838 B.n102 10.6151
R1771 B.n832 B.n102 10.6151
R1772 B.n832 B.n831 10.6151
R1773 B.n831 B.n830 10.6151
R1774 B.n830 B.n109 10.6151
R1775 B.n824 B.n109 10.6151
R1776 B.n824 B.n823 10.6151
R1777 B.n823 B.n822 10.6151
R1778 B.n822 B.n116 10.6151
R1779 B.n816 B.n116 10.6151
R1780 B.n816 B.n815 10.6151
R1781 B.n814 B.n123 10.6151
R1782 B.n156 B.n123 10.6151
R1783 B.n157 B.n156 10.6151
R1784 B.n160 B.n157 10.6151
R1785 B.n161 B.n160 10.6151
R1786 B.n164 B.n161 10.6151
R1787 B.n165 B.n164 10.6151
R1788 B.n168 B.n165 10.6151
R1789 B.n169 B.n168 10.6151
R1790 B.n172 B.n169 10.6151
R1791 B.n173 B.n172 10.6151
R1792 B.n176 B.n173 10.6151
R1793 B.n177 B.n176 10.6151
R1794 B.n180 B.n177 10.6151
R1795 B.n181 B.n180 10.6151
R1796 B.n184 B.n181 10.6151
R1797 B.n185 B.n184 10.6151
R1798 B.n188 B.n185 10.6151
R1799 B.n189 B.n188 10.6151
R1800 B.n192 B.n189 10.6151
R1801 B.n197 B.n194 10.6151
R1802 B.n198 B.n197 10.6151
R1803 B.n201 B.n198 10.6151
R1804 B.n202 B.n201 10.6151
R1805 B.n205 B.n202 10.6151
R1806 B.n206 B.n205 10.6151
R1807 B.n209 B.n206 10.6151
R1808 B.n210 B.n209 10.6151
R1809 B.n213 B.n210 10.6151
R1810 B.n218 B.n215 10.6151
R1811 B.n219 B.n218 10.6151
R1812 B.n222 B.n219 10.6151
R1813 B.n223 B.n222 10.6151
R1814 B.n226 B.n223 10.6151
R1815 B.n227 B.n226 10.6151
R1816 B.n230 B.n227 10.6151
R1817 B.n231 B.n230 10.6151
R1818 B.n234 B.n231 10.6151
R1819 B.n235 B.n234 10.6151
R1820 B.n238 B.n235 10.6151
R1821 B.n239 B.n238 10.6151
R1822 B.n242 B.n239 10.6151
R1823 B.n243 B.n242 10.6151
R1824 B.n246 B.n243 10.6151
R1825 B.n247 B.n246 10.6151
R1826 B.n250 B.n247 10.6151
R1827 B.n252 B.n250 10.6151
R1828 B.n253 B.n252 10.6151
R1829 B.n808 B.n253 10.6151
R1830 B.n479 B.n413 9.36635
R1831 B.n456 B.n416 9.36635
R1832 B.n193 B.n192 9.36635
R1833 B.n215 B.n214 9.36635
R1834 B.n952 B.n0 8.11757
R1835 B.n952 B.n1 8.11757
R1836 B.n662 B.t2 5.30682
R1837 B.n40 B.t1 5.30682
R1838 B.t7 B.n264 3.18429
R1839 B.t3 B.n16 3.18429
R1840 B.n476 B.n413 1.24928
R1841 B.n459 B.n416 1.24928
R1842 B.n194 B.n193 1.24928
R1843 B.n214 B.n213 1.24928
R1844 VP.n25 VP.n24 161.3
R1845 VP.n26 VP.n21 161.3
R1846 VP.n28 VP.n27 161.3
R1847 VP.n29 VP.n20 161.3
R1848 VP.n31 VP.n30 161.3
R1849 VP.n32 VP.n19 161.3
R1850 VP.n34 VP.n33 161.3
R1851 VP.n35 VP.n18 161.3
R1852 VP.n38 VP.n37 161.3
R1853 VP.n39 VP.n17 161.3
R1854 VP.n41 VP.n40 161.3
R1855 VP.n42 VP.n16 161.3
R1856 VP.n44 VP.n43 161.3
R1857 VP.n45 VP.n15 161.3
R1858 VP.n47 VP.n46 161.3
R1859 VP.n48 VP.n14 161.3
R1860 VP.n50 VP.n49 161.3
R1861 VP.n93 VP.n92 161.3
R1862 VP.n91 VP.n1 161.3
R1863 VP.n90 VP.n89 161.3
R1864 VP.n88 VP.n2 161.3
R1865 VP.n87 VP.n86 161.3
R1866 VP.n85 VP.n3 161.3
R1867 VP.n84 VP.n83 161.3
R1868 VP.n82 VP.n4 161.3
R1869 VP.n81 VP.n80 161.3
R1870 VP.n78 VP.n5 161.3
R1871 VP.n77 VP.n76 161.3
R1872 VP.n75 VP.n6 161.3
R1873 VP.n74 VP.n73 161.3
R1874 VP.n72 VP.n7 161.3
R1875 VP.n71 VP.n70 161.3
R1876 VP.n69 VP.n8 161.3
R1877 VP.n68 VP.n67 161.3
R1878 VP.n65 VP.n9 161.3
R1879 VP.n64 VP.n63 161.3
R1880 VP.n62 VP.n10 161.3
R1881 VP.n61 VP.n60 161.3
R1882 VP.n59 VP.n11 161.3
R1883 VP.n58 VP.n57 161.3
R1884 VP.n56 VP.n12 161.3
R1885 VP.n55 VP.n54 161.3
R1886 VP.n53 VP.n52 87.1314
R1887 VP.n94 VP.n0 87.1314
R1888 VP.n51 VP.n13 87.1314
R1889 VP.n23 VP.n22 73.9973
R1890 VP.n22 VP.t6 64.9339
R1891 VP.n52 VP.n51 50.8857
R1892 VP.n60 VP.n59 44.3785
R1893 VP.n86 VP.n2 44.3785
R1894 VP.n43 VP.n15 44.3785
R1895 VP.n73 VP.n72 40.4934
R1896 VP.n73 VP.n6 40.4934
R1897 VP.n30 VP.n19 40.4934
R1898 VP.n30 VP.n29 40.4934
R1899 VP.n60 VP.n10 36.6083
R1900 VP.n86 VP.n85 36.6083
R1901 VP.n43 VP.n42 36.6083
R1902 VP.n53 VP.t1 33.0649
R1903 VP.n66 VP.t7 33.0649
R1904 VP.n79 VP.t0 33.0649
R1905 VP.n0 VP.t4 33.0649
R1906 VP.n13 VP.t2 33.0649
R1907 VP.n36 VP.t3 33.0649
R1908 VP.n23 VP.t5 33.0649
R1909 VP.n54 VP.n12 24.4675
R1910 VP.n58 VP.n12 24.4675
R1911 VP.n59 VP.n58 24.4675
R1912 VP.n64 VP.n10 24.4675
R1913 VP.n65 VP.n64 24.4675
R1914 VP.n67 VP.n8 24.4675
R1915 VP.n71 VP.n8 24.4675
R1916 VP.n72 VP.n71 24.4675
R1917 VP.n77 VP.n6 24.4675
R1918 VP.n78 VP.n77 24.4675
R1919 VP.n80 VP.n78 24.4675
R1920 VP.n84 VP.n4 24.4675
R1921 VP.n85 VP.n84 24.4675
R1922 VP.n90 VP.n2 24.4675
R1923 VP.n91 VP.n90 24.4675
R1924 VP.n92 VP.n91 24.4675
R1925 VP.n47 VP.n15 24.4675
R1926 VP.n48 VP.n47 24.4675
R1927 VP.n49 VP.n48 24.4675
R1928 VP.n34 VP.n19 24.4675
R1929 VP.n35 VP.n34 24.4675
R1930 VP.n37 VP.n35 24.4675
R1931 VP.n41 VP.n17 24.4675
R1932 VP.n42 VP.n41 24.4675
R1933 VP.n24 VP.n21 24.4675
R1934 VP.n28 VP.n21 24.4675
R1935 VP.n29 VP.n28 24.4675
R1936 VP.n66 VP.n65 23.4888
R1937 VP.n79 VP.n4 23.4888
R1938 VP.n36 VP.n17 23.4888
R1939 VP.n25 VP.n22 3.37702
R1940 VP.n54 VP.n53 2.93654
R1941 VP.n92 VP.n0 2.93654
R1942 VP.n49 VP.n13 2.93654
R1943 VP.n67 VP.n66 0.97918
R1944 VP.n80 VP.n79 0.97918
R1945 VP.n37 VP.n36 0.97918
R1946 VP.n24 VP.n23 0.97918
R1947 VP.n51 VP.n50 0.354971
R1948 VP.n55 VP.n52 0.354971
R1949 VP.n94 VP.n93 0.354971
R1950 VP VP.n94 0.26696
R1951 VP.n26 VP.n25 0.189894
R1952 VP.n27 VP.n26 0.189894
R1953 VP.n27 VP.n20 0.189894
R1954 VP.n31 VP.n20 0.189894
R1955 VP.n32 VP.n31 0.189894
R1956 VP.n33 VP.n32 0.189894
R1957 VP.n33 VP.n18 0.189894
R1958 VP.n38 VP.n18 0.189894
R1959 VP.n39 VP.n38 0.189894
R1960 VP.n40 VP.n39 0.189894
R1961 VP.n40 VP.n16 0.189894
R1962 VP.n44 VP.n16 0.189894
R1963 VP.n45 VP.n44 0.189894
R1964 VP.n46 VP.n45 0.189894
R1965 VP.n46 VP.n14 0.189894
R1966 VP.n50 VP.n14 0.189894
R1967 VP.n56 VP.n55 0.189894
R1968 VP.n57 VP.n56 0.189894
R1969 VP.n57 VP.n11 0.189894
R1970 VP.n61 VP.n11 0.189894
R1971 VP.n62 VP.n61 0.189894
R1972 VP.n63 VP.n62 0.189894
R1973 VP.n63 VP.n9 0.189894
R1974 VP.n68 VP.n9 0.189894
R1975 VP.n69 VP.n68 0.189894
R1976 VP.n70 VP.n69 0.189894
R1977 VP.n70 VP.n7 0.189894
R1978 VP.n74 VP.n7 0.189894
R1979 VP.n75 VP.n74 0.189894
R1980 VP.n76 VP.n75 0.189894
R1981 VP.n76 VP.n5 0.189894
R1982 VP.n81 VP.n5 0.189894
R1983 VP.n82 VP.n81 0.189894
R1984 VP.n83 VP.n82 0.189894
R1985 VP.n83 VP.n3 0.189894
R1986 VP.n87 VP.n3 0.189894
R1987 VP.n88 VP.n87 0.189894
R1988 VP.n89 VP.n88 0.189894
R1989 VP.n89 VP.n1 0.189894
R1990 VP.n93 VP.n1 0.189894
R1991 VDD1 VDD1.n0 74.6636
R1992 VDD1.n3 VDD1.n2 74.5499
R1993 VDD1.n3 VDD1.n1 74.5499
R1994 VDD1.n5 VDD1.n4 72.8639
R1995 VDD1.n5 VDD1.n3 44.3586
R1996 VDD1.n4 VDD1.t4 3.89048
R1997 VDD1.n4 VDD1.t5 3.89048
R1998 VDD1.n0 VDD1.t1 3.89048
R1999 VDD1.n0 VDD1.t2 3.89048
R2000 VDD1.n2 VDD1.t7 3.89048
R2001 VDD1.n2 VDD1.t3 3.89048
R2002 VDD1.n1 VDD1.t6 3.89048
R2003 VDD1.n1 VDD1.t0 3.89048
R2004 VDD1 VDD1.n5 1.68369
C0 VDD2 VDD1 2.35111f
C1 VDD1 VN 0.153419f
C2 VDD1 VP 4.67918f
C3 VDD2 VTAIL 6.67373f
C4 VTAIL VN 5.54352f
C5 VTAIL VP 5.55762f
C6 VDD2 VN 4.19725f
C7 VDD2 VP 0.641767f
C8 VP VN 7.74297f
C9 VDD1 VTAIL 6.61188f
C10 VDD2 B 6.04452f
C11 VDD1 B 6.61615f
C12 VTAIL B 6.526974f
C13 VN B 19.10563f
C14 VP B 17.714115f
C15 VDD1.t1 B 0.120884f
C16 VDD1.t2 B 0.120884f
C17 VDD1.n0 B 1.00533f
C18 VDD1.t6 B 0.120884f
C19 VDD1.t0 B 0.120884f
C20 VDD1.n1 B 1.00395f
C21 VDD1.t7 B 0.120884f
C22 VDD1.t3 B 0.120884f
C23 VDD1.n2 B 1.00395f
C24 VDD1.n3 B 4.24734f
C25 VDD1.t4 B 0.120884f
C26 VDD1.t5 B 0.120884f
C27 VDD1.n4 B 0.986924f
C28 VDD1.n5 B 3.40316f
C29 VP.t4 B 1.08397f
C30 VP.n0 B 0.487289f
C31 VP.n1 B 0.021918f
C32 VP.n2 B 0.042477f
C33 VP.n3 B 0.021918f
C34 VP.n4 B 0.040043f
C35 VP.n5 B 0.021918f
C36 VP.n6 B 0.043562f
C37 VP.n7 B 0.021918f
C38 VP.n8 B 0.040849f
C39 VP.n9 B 0.021918f
C40 VP.t7 B 1.08397f
C41 VP.n10 B 0.044192f
C42 VP.n11 B 0.021918f
C43 VP.n12 B 0.040849f
C44 VP.t2 B 1.08397f
C45 VP.n13 B 0.487289f
C46 VP.n14 B 0.021918f
C47 VP.n15 B 0.042477f
C48 VP.n16 B 0.021918f
C49 VP.n17 B 0.040043f
C50 VP.n18 B 0.021918f
C51 VP.n19 B 0.043562f
C52 VP.n20 B 0.021918f
C53 VP.n21 B 0.040849f
C54 VP.t6 B 1.3656f
C55 VP.n22 B 0.468227f
C56 VP.t5 B 1.08397f
C57 VP.n23 B 0.476388f
C58 VP.n24 B 0.021489f
C59 VP.n25 B 0.278822f
C60 VP.n26 B 0.021918f
C61 VP.n27 B 0.021918f
C62 VP.n28 B 0.040849f
C63 VP.n29 B 0.043562f
C64 VP.n30 B 0.017719f
C65 VP.n31 B 0.021918f
C66 VP.n32 B 0.021918f
C67 VP.n33 B 0.021918f
C68 VP.n34 B 0.040849f
C69 VP.n35 B 0.040849f
C70 VP.t3 B 1.08397f
C71 VP.n36 B 0.406811f
C72 VP.n37 B 0.021489f
C73 VP.n38 B 0.021918f
C74 VP.n39 B 0.021918f
C75 VP.n40 B 0.021918f
C76 VP.n41 B 0.040849f
C77 VP.n42 B 0.044192f
C78 VP.n43 B 0.018173f
C79 VP.n44 B 0.021918f
C80 VP.n45 B 0.021918f
C81 VP.n46 B 0.021918f
C82 VP.n47 B 0.040849f
C83 VP.n48 B 0.040849f
C84 VP.n49 B 0.023102f
C85 VP.n50 B 0.035375f
C86 VP.n51 B 1.29132f
C87 VP.n52 B 1.3068f
C88 VP.t1 B 1.08397f
C89 VP.n53 B 0.487289f
C90 VP.n54 B 0.023102f
C91 VP.n55 B 0.035375f
C92 VP.n56 B 0.021918f
C93 VP.n57 B 0.021918f
C94 VP.n58 B 0.040849f
C95 VP.n59 B 0.042477f
C96 VP.n60 B 0.018173f
C97 VP.n61 B 0.021918f
C98 VP.n62 B 0.021918f
C99 VP.n63 B 0.021918f
C100 VP.n64 B 0.040849f
C101 VP.n65 B 0.040043f
C102 VP.n66 B 0.406811f
C103 VP.n67 B 0.021489f
C104 VP.n68 B 0.021918f
C105 VP.n69 B 0.021918f
C106 VP.n70 B 0.021918f
C107 VP.n71 B 0.040849f
C108 VP.n72 B 0.043562f
C109 VP.n73 B 0.017719f
C110 VP.n74 B 0.021918f
C111 VP.n75 B 0.021918f
C112 VP.n76 B 0.021918f
C113 VP.n77 B 0.040849f
C114 VP.n78 B 0.040849f
C115 VP.t0 B 1.08397f
C116 VP.n79 B 0.406811f
C117 VP.n80 B 0.021489f
C118 VP.n81 B 0.021918f
C119 VP.n82 B 0.021918f
C120 VP.n83 B 0.021918f
C121 VP.n84 B 0.040849f
C122 VP.n85 B 0.044192f
C123 VP.n86 B 0.018173f
C124 VP.n87 B 0.021918f
C125 VP.n88 B 0.021918f
C126 VP.n89 B 0.021918f
C127 VP.n90 B 0.040849f
C128 VP.n91 B 0.040849f
C129 VP.n92 B 0.023102f
C130 VP.n93 B 0.035375f
C131 VP.n94 B 0.066201f
C132 VTAIL.t14 B 0.104986f
C133 VTAIL.t15 B 0.104986f
C134 VTAIL.n0 B 0.796791f
C135 VTAIL.n1 B 0.530915f
C136 VTAIL.t10 B 1.01978f
C137 VTAIL.n2 B 0.628873f
C138 VTAIL.t7 B 1.01978f
C139 VTAIL.n3 B 0.628873f
C140 VTAIL.t5 B 0.104986f
C141 VTAIL.t2 B 0.104986f
C142 VTAIL.n4 B 0.796791f
C143 VTAIL.n5 B 0.818935f
C144 VTAIL.t4 B 1.01978f
C145 VTAIL.n6 B 1.60587f
C146 VTAIL.t13 B 1.01979f
C147 VTAIL.n7 B 1.60586f
C148 VTAIL.t9 B 0.104986f
C149 VTAIL.t12 B 0.104986f
C150 VTAIL.n8 B 0.796795f
C151 VTAIL.n9 B 0.818931f
C152 VTAIL.t11 B 1.01979f
C153 VTAIL.n10 B 0.628867f
C154 VTAIL.t3 B 1.01979f
C155 VTAIL.n11 B 0.628867f
C156 VTAIL.t1 B 0.104986f
C157 VTAIL.t0 B 0.104986f
C158 VTAIL.n12 B 0.796795f
C159 VTAIL.n13 B 0.818931f
C160 VTAIL.t6 B 1.01978f
C161 VTAIL.n14 B 1.60587f
C162 VTAIL.t8 B 1.01978f
C163 VTAIL.n15 B 1.60097f
C164 VDD2.t5 B 0.118313f
C165 VDD2.t0 B 0.118313f
C166 VDD2.n0 B 0.9826f
C167 VDD2.t7 B 0.118313f
C168 VDD2.t6 B 0.118313f
C169 VDD2.n1 B 0.9826f
C170 VDD2.n2 B 4.09622f
C171 VDD2.t3 B 0.118313f
C172 VDD2.t1 B 0.118313f
C173 VDD2.n3 B 0.965939f
C174 VDD2.n4 B 3.29396f
C175 VDD2.t2 B 0.118313f
C176 VDD2.t4 B 0.118313f
C177 VDD2.n5 B 0.982556f
C178 VN.t7 B 1.04605f
C179 VN.n0 B 0.470242f
C180 VN.n1 B 0.021151f
C181 VN.n2 B 0.040991f
C182 VN.n3 B 0.021151f
C183 VN.n4 B 0.038642f
C184 VN.n5 B 0.021151f
C185 VN.n6 B 0.042038f
C186 VN.n7 B 0.021151f
C187 VN.n8 B 0.03942f
C188 VN.t5 B 1.31783f
C189 VN.n9 B 0.451846f
C190 VN.t1 B 1.04605f
C191 VN.n10 B 0.459721f
C192 VN.n11 B 0.020737f
C193 VN.n12 B 0.269067f
C194 VN.n13 B 0.021151f
C195 VN.n14 B 0.021151f
C196 VN.n15 B 0.03942f
C197 VN.n16 B 0.042038f
C198 VN.n17 B 0.017099f
C199 VN.n18 B 0.021151f
C200 VN.n19 B 0.021151f
C201 VN.n20 B 0.021151f
C202 VN.n21 B 0.03942f
C203 VN.n22 B 0.03942f
C204 VN.t0 B 1.04605f
C205 VN.n23 B 0.392579f
C206 VN.n24 B 0.020737f
C207 VN.n25 B 0.021151f
C208 VN.n26 B 0.021151f
C209 VN.n27 B 0.021151f
C210 VN.n28 B 0.03942f
C211 VN.n29 B 0.042646f
C212 VN.n30 B 0.017537f
C213 VN.n31 B 0.021151f
C214 VN.n32 B 0.021151f
C215 VN.n33 B 0.021151f
C216 VN.n34 B 0.03942f
C217 VN.n35 B 0.03942f
C218 VN.n36 B 0.022294f
C219 VN.n37 B 0.034138f
C220 VN.n38 B 0.063885f
C221 VN.t2 B 1.04605f
C222 VN.n39 B 0.470242f
C223 VN.n40 B 0.021151f
C224 VN.n41 B 0.040991f
C225 VN.n42 B 0.021151f
C226 VN.n43 B 0.038642f
C227 VN.n44 B 0.021151f
C228 VN.t6 B 1.04605f
C229 VN.n45 B 0.392579f
C230 VN.n46 B 0.042038f
C231 VN.n47 B 0.021151f
C232 VN.n48 B 0.03942f
C233 VN.t4 B 1.31783f
C234 VN.n49 B 0.451846f
C235 VN.t3 B 1.04605f
C236 VN.n50 B 0.459721f
C237 VN.n51 B 0.020737f
C238 VN.n52 B 0.269067f
C239 VN.n53 B 0.021151f
C240 VN.n54 B 0.021151f
C241 VN.n55 B 0.03942f
C242 VN.n56 B 0.042038f
C243 VN.n57 B 0.017099f
C244 VN.n58 B 0.021151f
C245 VN.n59 B 0.021151f
C246 VN.n60 B 0.021151f
C247 VN.n61 B 0.03942f
C248 VN.n62 B 0.03942f
C249 VN.n63 B 0.020737f
C250 VN.n64 B 0.021151f
C251 VN.n65 B 0.021151f
C252 VN.n66 B 0.021151f
C253 VN.n67 B 0.03942f
C254 VN.n68 B 0.042646f
C255 VN.n69 B 0.017537f
C256 VN.n70 B 0.021151f
C257 VN.n71 B 0.021151f
C258 VN.n72 B 0.021151f
C259 VN.n73 B 0.03942f
C260 VN.n74 B 0.03942f
C261 VN.n75 B 0.022294f
C262 VN.n76 B 0.034138f
C263 VN.n77 B 1.25474f
.ends

